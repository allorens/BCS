BZh91AY&SY��e��d߀@qg���#� ����bG��     o
� �I T� �(U*!B@E@P�� D@R�@�H(�P(�Q R��U$�����v�T�BUHEE%U�J%
�QH(�	P�T�(�H%TR��(�E
���T�*����JD�(�� ��$�((@UJ�UT�!UT�$�R����R���*������QJH��
UB���H�b�$��  �uE	���L� С��QB��R�)��P��dY��� �R���%@\�JRR
)R �**�   pk@ 6��P(�X4  Z0@41� +A��
kMӻ� ��` )�l�Ph���;�  ��R�J�)H��*   k8  :q�p  ��v�U�n�(��� r�p t �`��r  ��� ���8  9R
��% DU �  �t h� t Uw4t ���  ;)�� ��  6C��* �e  ���� X�JD��A$��	*C�  fqB��X0 P��� P-&� F, 440  `� ��� 
!�h( 5��� ��J*J*HEP� 7  ,�� Y&�¨ Ņ �1�R�j��0�c
 K��֌1� J`�$��UD����p  �qC@fS ����(�� hQ� �L  ���@٪ a����Pu��*ERUAIAJQD  �  s �ElK�iV �ɀ!mU
�6�((P�V��Xmm LBR�J�� !�  Zv� 6�P(jaJ ��aE3J�P �(P�( P��H�P #QB�0ЪPB R���J�   c�AƦ  ��QUXc 
� Y�@!�
� 
أ�A20 )�    �   j`�JT22�h0�4��T�aJQT�� � 4   9�d�a0L!�# <RT� 	�  4Ɇ�l��Mi��#L ��ީi��M�m&Sd��i��C'�1?������������&�<n��+&'5Қ����j�ax:��s�� �{���� *��*}@_�* *����c���������7�}?�" *��&*��@_�������ObAU}����o/���>����{0�`_��>��`f� ��:�=eN��D�
u�:aN�'�
u�:ʝdN��X,�X����
u�=�S�#�T�"u�:�Y:�=dN�X����=`�'Y�	�,��
u�:ʝ`fA� ��:�=`��d��X �(��:�>��A�"f��X�#�� ��:ʝaOL)�P�a�q����T� �0X����*zeN�'XG��:�=d�XW����
|2�YB`�
u�:�=eN�'YC���P�"u�:��X�	�P�
u�:�dN�Y�)���zʝ`�'Y���� ��}0�Y�:Ƚe��XW���U� eO����U� e^��E�
��<�a^��YW� u�}�����d��X��E� ��ze���"��z��a��Y_f���#�U� Y �*`3 ��N���U2��eAz���a���eAz����U� �UC�*�YP^���`Dz��0�=`z����*��PG��{0"dPz� ���"��A���EW���Y� �e��������"��W�" u��"��EG���XQ� ���ez�=`^���:½a^��U� a^���/XW��� <0�Y� u�z�=dO,d�XG���eN�����M>��p�VL�]�Ƨ~�����:�M]�N��l2nz�!笝�d#(tz��L��V��a�5��Y��J�ܕ�`�׬�Q!3F,L��ԫ�U���|�� 6��-_�m����,�]��Ϣ�{.=:.���B�P|+Mw7�c�[�*v��X���I�de��y��a��iU�Pº�:�g�8��nfnw7��3����R�xb�z����V��$^j�Pٶ���_��k�1J�1�]\wfSA�:�7x�-�a�CZ��e�C-��h�Yݻ�� ��"|����tW$��X����W���f�wj�n匘��љ��v�[��&jv�Fx��:��q��a�R�Q ^&����eBP����'�0��л�)\/ͦHu��{����A�)n�&�r_�Q���T+uQ�Y��e[�LzR�^�Ն���i9�jmTѫ*u��澤�(�lVf,�h�4��]�N:yjd�-�����ai��!�V5�k���e,�@�А���:n�Ǳ�ӫJUa�+O.�t���6������z�k�:v���8
�{�sA� �TB+7L�Ur�5�ɧ��4a"��E�ʳÅEQ��wW���s�P�ɖ�J���]�Y���g�����%)�������z�m��~�ӧ������AC2��(��4�wb�+S�~�ׯ�v���P�랭�׷�a"��2���؍��!��K�<����(4h��9.��D�I.���,���K5-��Pթf��"ou&����V˞�,m�w^2�
w�n�7����9�R�{��K2�e4���{��4�/g���&�%�\��y����2��\@f�	�a"�!	�a����1.�{Y�Pےm��,]��D]nb�R��V*�8kB:�V��^S�Z��b�^��O#x&�e�����7xi�yie
�Yb�-�r��Kh@	�"��)Lk���q1��f�#��&^>@����E����I�Cqm2.=���^`#c�W�xZ�ڌigAT_���XX�(7tY�:���m=��0����юe��������2���4�āϕ`����l��s�O
(�1&�:�]���Ց�B�bu��&F�[�2�b�z�����=r�^=3&6.���WelE�Y�S�	@���\7��:K�=U���cʹR��J�0c����ǆ\�P�
Ԭ�4˳:��'m�V�L�tz�T�q�L���c�ݻ�g1V:w�e4�ڤ҆�4��(�U�L\,�^{`.X�;e�V�oXx.e��*�fd�݅b��Y� �t'<Z�h��y¥-�eʺX�~R�.�sB9��S����$+�G49s��*�;l^E�e�V*�A��:�����^m�{`�5S͹M���iP��(
׹cX@�q�	��_.Zs^�e妆;
Mv��Vh0�Sa:���*�Gs|�ي�m&uqM����)'��,�R���g ��ӠE�k1��m6u,�5yX7�Zˣֶl{k�葕����k�ɛ���;�+R�*�/62�t[���W�5�ሆ"�k��{G�	�%^,���W��8w��7�/�!��/�d�Au��7�E7t��w��9�t+\�Ñh>f�+�Zu�\q���������v�b&kcJժ�f�ԗ��3GZ�sxN�\�De$��lwݩn��(�2���2��{�4�^�ɭ�у���X�9%˖�Ӥ�정�|���]l�C���J�ff�h�>ij�B���,uwAh���J�4�~ߪ�����YF꘠�]��u�,VOU&z�X��C��������^��=u��PV�iYMc��[�:*��e����T�� ���S.��o<��["f@jaN��Z��3�-�e�݄Îڍ]F��kf�x4Ւ��f���ZvBtM%BQ�q �j[�h:yFI��jDpb�]m1�[mx�ye�������v��Cj�df���՜�m�*���gNR� �i]ӵ66���$ZaXe�N]ص+��n�b�%��[���3Rg)k1���mن�Zَ�eY,7Vw��ct�G^�ҁ;y�!uA�]ޕf�<�ұaPt�;:����s%K.�Q����L�xl2м��h�6G-f�t]�9����`htܻ;��1�1�*���Y,���)�t�qi��#���,���5	nL:�{B��p��-�g+#�e`'!o%M;Ǜ��˄=EM�a�ya���J���`5n���h�U��Y�B�klҵ�rd,h{�y2�24T����co�#�X%�J��e������2��,�n�/6�u0M�`�̓)d(�T�y�4�����'��a�U[n�#r�3���, �<�71(0�/� ��T�!��]G�k��˺���7.��MA�⍨��F�U���/@����El6*���b�!Xݹt�ڀ���2,�(�Ԧ�˭������GP*�69oS�2��w�m�uK4�6���L�BY#ɔK*��z�
<Mb��K)�u���-RͰ�[k���!Wk�%��{8�B���G#����R��yzFX��K�H4n[.*�Vܺ%f��v�F�ӵTΔ5��ټ�^Z�{%���&�ĕiD��:�v�d�)k6+-ȱ�mP`֥�����7�C�6?L�7)[�`GqǹPh7R`��x���n�[8r�%�y�1-�+S�޼QC,�	�	���ҿ���%
�t�j\cx^EM���Y1�F�/Pv,�� ^��{�ө(n�xu��x�&���]��ěp�kN���̙Z�4�T����Yв��䵸kk'	
�z�g��e�����"� lkM�M���wZ*��g�{�+	i�pA�7�3sUSjm�^�m���l����f =yF5(cL�n�Bf�]eK�J=�2�M�G)��,�ݸ/Ua��7i�lٵ�nVk���*Ն��Uw��G6�l2^�b�P�V��crܚ�g.�n��Zn�ɖ�ǣ���#ț� Ǚ.����M^<[aH�lm����p�:M�7m-�|	i����:�MECl��u��:V�ā���oP;یˢ�-����T��J���A������7���`Yɗ��+J[-,�ǩ�~�4�k�ԩ&�Lc*�h*��e�0�
 ]�����ez�yY��d��u�CA��1�xr:��gAi�;R����@b�2�	���P��1��Un��5�"��:fڗX0U�P��4��UtԻ%�JJF��B�e���f+��n��)�l���eY�jj��c+X�h֭�Ե֓�/2�{-hmn�J����r�6Ţ��7H��z9�^w�b�Sy�X�)Z(`C*��"�$l�S`@��]���CzYݦ^2-,;SI�����wW5����ٱ	����ƃ�雤ۤ��դ#w&N>۫�{���b-ۦv"���JB�;\��iس�qU�[B��7�j��i~��ZP��] �o*�F��[;1�1O	6�%��M� �Ֆ%]�ɊD�.��%��hl�f
B��v�:@If.loJ�f3� ����5b/j�(�b�IM�H#�����}0+j�Ùt26�j���ZN��W'�O��&��ST��b�&d0���B,���a�62����LI"%Jɢ�,�u����i�%��T�1�Lto��^ѱ�m%�dj�|{G�$�sz�a��[�ܶ�%���.�s�2��Ŗ�W�/��Z9��V���;[���F>9��eS:���-�����g�������ڿcP���ku��8�<�;�G��4�� �+3m�c�(]�,fS'4!��Eb�1��cC9b�N����P�z�J�Z��������
� ��9I=�C���Gt��]:V1�$�ܢ�ګ��`��TY1����Ⱦƫ.�YA������W�Z�2kJX aM�l��¦M���k��Q��U�]�{QV]��X�M�#�v�2skB��*к����K�%��h��&c-"4���W[5��YIl>,[C�Q����\,Vn�X��QQ�*�d��k\��޴���d�m�2k(�pe.�<���m�1�T:ڴ�cB�H[.ݵ$'j֑�-��ǧwknG��m�IX@LlcZ��4:�y���m�D��sIӇ.�^�B���d���-��x��gN��w���Үej!d��ݣ�#t����l��4= ��("�Q@,pY���y����A�ܶ�1y���ʦFu���zqؒ*H 4C�	�d��9W�i��7-�-e�jj�H\����YxZ}owM�d:=�l:���9�����Y�d�"�L�xZ�[:�{E�օr�z𛢰��
gw�4t��h�|�����w�am���ūl*wL^'0`�6�p�̄&�h:�{cEn����)��7t�ԭ+i�V�M,u��#U�6�t�:��[j����^�ե��Bµ�V�tcJ�x�L�9u+(]2�d���r�u�fb
Չ2�d^͗LVl������:z��60���1�־��n���e�+
��fL�7�ng��tZ�oV!·��U]#~m�,<�*�o3B=+ń�W�⵲�[�1�uwJT�F�`'-��
�X�k>�(Y#O,���m*'w����O�K;��f`�)�-bȰk[f�J��چ��B�&)&�Q��2��p]�
2�^f܉Z��&�E�<C�u��������E�9�9���qV��ҭ:!�I�k}����њj�Xҋ*�c݆k�37jT�d�P̗R�鈰K��[�h�� !�K^��w[�ZՍ0e;9Z&ָ�C0!�6sOkv����G��u7�M#��v�eN��:�uұ��v���߬��Xb�W� A��
���B��y��a�(��yө]��	bC���NCYsf�f�r'�={���/V�ٙ��I���{�f]�Wd�VsojU���M�K���y!urZq6W�a���x�U*�vn�����gsT�����p�!��VSi�1Ptzc��* v􏺚���xv���J�Kj+O<�h��О��n�X�%QKR�4�����A�=��m�C���0�L%z[�{uq8��c����Ӑ�ڗ�$(�7��G��pۛ-��7��]����v/p.4;J}�L��K��'l�y���a�F��-1�v64݊�(�+vb�YJ�i�������x�ə���J�S*a���*�d�!���V)c^��ͱ��r�cfDP61�0��[Z��֞��VU�M��Q�W��a�tg�ֵ��t	���.���� �h����v0h-YG^��(eng�s���Ҷ�`��teY��hfM�1+����ha�]>��˦E^�dV�-M��-���%j�7��@st9��]�mY�
{�m��3�ujH�Fr�X�S#�U�<TZ�y(�����m�)mf3R�u��<M�6���n�v�Z�(��	j��v[�k<��]w��hmr���u�NY%�7��m�׳2<�v��@��U��f�:�7�YVi���2ʽ:�A&�v�]�b�,�KW��s>P#ʕ�м,\�0֡.
xǎ�D� kD�*���74�9nV���/I�/lX|��A�MH����]��V�=�i�I�]w�q�A��1c��
%��i�h�0��UO/D�aX��,��ה�@֨���X�db/�$m�M<�)ʺ�Jj��ǥ�SB/�nW����S�iĈW�R���Ֆ�є��;F^j��N��B�!x�^��Xe��KC�!�����)A{��O)�)ai���Y�\S#~�۱u���Zw+nãy"��nl-�,aT�}g��)� )����n����w��VY�ֵ@��������6�����]�V��H�r,�9�
f��*��؅խ�˼-��L&��)��ŕti7�F��Z���q�V�BF�u�kb��1m�Y{�����L�gL�]M!��s��2��z�k����:�X�_e�Ch��|�mY�l��նU�!�ȋ��]锖
J.U�6�5��t*��3k36CԘ#u�EU�A�-f:l$�v6E̏&[.θ��S�xX3�Zv�!Y2�^���Q,"Ԣ(ӓa�Yb��+�	���X�t��2�i�C���E;��K4E��
�{��!a`�J�[��(�(���n��L����h�������Z�aD���a�ե�8Cܤ�y =d�}�UT���u�͌}g[J��ûyGr�U�=��]c�7��Y��b�p�f�!�/-��шCɒ[��J͐nm��[y��D�ڑ��R���3��XK�R� �VZξ	�V���_5o7m5���!�Nv�P1���!��^��՗��ɻ�Iď����9�f��ú��JV;����]�D��6/�Xq���ʵ�e�2����u@a�њY!�Rf�bX�v����!�����3+�q���/�f�R.�v�L��:]�K�J՗PF�J�0����U$X�:���:td�#�o0-��%bZb�rB�*�31�V �5v�Y�$@�[:���*R�G��F1tp٬�a�ʃ@����c6�v5'@����R���t��7K,�gdH���]]�@�:R(.�J��*�{Q��ceE�+�|mq[Z�KU��tVJ�2� ���]G�Mn��B�I*���(�<�D�FQ�[շk����ךQ��t�7��ୢ�놌eDq�KKK��o��]gj�����ZΈ�"H����Uv�8����:r۽vV�+���sM�k�������$��o)��h��.�p���JCEiЁ�p�b��c��ci\�
;f�
`ي��dL�k\G0kO�+��4_^Z�Gw76����Oe[���3tGx�d�&���j�)^t�gO9��(K��Ls�[u�:-���8Qt��a�[�2��f68B��+����Ex���Y�;������gs���>�}�xa�/��7���wt�I$�I$�I$�9�9Ud�$RT�I#�I$�H$�32I&I$�U^Nw1j�Q<4��Śj�������)r��R�6[�xNj�E]<�9Y����rYw=�EN�L���*�	]%\�P;ـ��t�q�˥-D,/�*�oOY[r���!> ���O]T�p2�m�YA��O}T��`��n�<5�L7������@z����Wm��U��dT_U\!%;W9�]���MAVM�n^^t"�J��өx�ҝ�[�f���4\�S!\�|�9��Oi�x�=�Sv�E�Y2�<܁��*�[(Z�B�넌�\�oB�ʙ�!�y��td[�K�
D�J�h�����Xo�< %�jK�X`I����3���ӔHz�i���M�|�K��{lf�p���Y���[���}E��/MV!��j+cv�k�X#��;[v����� �]1�<�4;��4�P��>����F젯�6�[n�]�3��"�컬�݂K��9��(Y���T}
V^N/����V��n��&���z���t��ϱj%��7GO+FJ�*+"�C|�i��*r�arR�.ޙ�֝��Ѱ��ݗ�@�ӡ�)b,j�����ݲ_lr]CMVp��YSN'y�t�*:<�\a�Y�4��ys�d&���m�`��Vy�&o&������1��k`}To��J��]«�%�<k��{��5[�ۺAE�	�ou����X5��ΑR��\�wuU��
����a��鳺�nr�W��xwp�5�$�aIv�-�mq��w7Wr]�͹YL���f1��4�{ΰ�vCÛYY���!w-�s�����`Mos�\���#%�|�]jg\.��wM7vg8s�a�^"�y���wc��.�zjU�l�v��X�<����$\��*���]�T�����-�a|{F���rp:����6:�Ȝ-�L�ٻK)�C"�a�%p�&t|(�F򑎮�m�Rj��%]e�[���S^^<_f��ɗ�bm����Ss/ Qv�>���9zl���1Yn9�Cf�\��4�,m�E*� t=�j�r,f�b���W#0�!�Qa�)^NѴE@n�	ƅ*�k�N�a�B@k���hѵ��;��^�lbYa�]+9��Ӭ����w]���qx�nzS˿`�!�R]w��;�Nb=�|��Xvh�z��S�=�����;m�͢׎⩮�l�/�q͆؁a���z7Q+b3��s��b�%�4�>��}h�c��U-�Z2��4�&�9����tCFFiA�Ԣ����t�6�Xnv`l������N�ל��$˻��J�θ����,ϣ������1�L��p'��U��-�Ba�q�I��!%%6��Vw���ɼ1���̹�T�9�)�H��cn�lf`ǃ�1��ԧo��b��O��c��M��;J�y`��9�����u`깫�:`�	��n�t�jL��n��۰��� UŒ�����l+�RemH��J��[�-��Kr���0��H2���v賣�̹&�UwK4h�&�g!#:�b�y�t�M7'Ib_FûvK�rpt��gj�I6a�ſ��kc��Z_jC&�B��K����U�,������H9�P��T:榢�z5�5�/	�4:����nb�+��&�	��I��jc�wӘ��S2�����aY{ָ�M�aWJ���<"!4�>c��|mZ��]�L��j�V�����s�J縰����c�]3�]A�x3S�/7&������8<�b�LV��`o5;�C���k�U]�C*�>P$-��/����nII���\�����:�ш�m]]Y�T�Xav):!�Im!|���	L�k��O"B�ͷӍ嗤<R���O9�G]�U��u��9�3��Σ�尝�(t�!���wi�g6<��s�}/�����Ĵ��V�������҇��O%v���˧@��ܺ���.*h�w�ؙ���ͧ����li�cj6����9��7�kH�׸�"�g(�=J�h��rP���J�fݍx/	�j��;��	Ud{�⃰�S6���q�6u�-N����kw[4�ɵ�Kia
,��y��w-1]N�a�B]�\�w59>*݄e�x6���p����EOB�X��,NQ�齾;S��7�u�e��.;��Q
=[F���b}��V�C��u_Tu3�+:=�����y�%G�ki����|f�B��Y۩�CM��`��uBP�Â�D���1���{S�����.���f�n��b�7�YC��q�y�V�s.oe������<Lc�&R<)M���=��;:���a���=U��8o7I}9���3�^��iz٬��u&�M5\nÐ��yؚ�jE9v�j����e7t+b�,�us���*���vR��MцN�&dt��3���0�Ə'��g��I6�����U+��Q�}e���>�2ӍɚN��[�C��L�9�<��agfQ��k�e�4�Bl�U���Y·cwyy�m[�h>��������[`�+-Ʋ�<�G[WdW"�o�-#qn�iP5����vƁxF����ȶ&��qWl�ѧ�t+�P�� ���Gŝd���ʪPv�͠��&YnU�$Ԇ���Af�I�7�b���Ǜ����7��::�p���p�dxج�`f��2��GJ����W}��'6�G8��[fҒW�0(�w7;nt!�*�.��Tɹ�]�W��l���= .wbQq����o]�N�V�1�������5�*�n�a�	#�L[
���~9QI��v�I��/�ga���X�ݝ�r5u|����#��SK��X;����j�H�p�ysZtѡ��t̠����V�$�j��ண�	����1HU��wU����;�c��^]��",E�lb��`��7��G�x\�7�KvNZ(QU�s7�ű���C�<�i��m��b�����Z8�,��HA�H�7�<ԌH
�4S��׮WT���!�V�L2��ƋLT߶�>�x�{7-C��ՎҠ�6����{�&'CL�A%���y�e��95�7�V�/r�ɔx�j:�,8�,�:��h��QSO*��zӥ1Le,;6�)M��ُ^�ΉrV��/i��g�j\Aܲ���5\�j��s��R����Mӛ{N8��McU�h*�~���p9�oc��p�Gh�]˥^��Y�G+�.5h��Ц��+%ʻ��L�z�S����d�:|z�׺�;c1{Ǿ����ʏ'4�E���]h�2A2.�+D9{�U�]8�(=�Y���fM+��*uB%�ĩVz��+�GՂt�{���I�n>�n�����r������R
Z���cY���L{�2�e�l���=��$ɍ��f7ԺoBk'c�B<t��	��ɚ��,y�:��݇2S�W9�j.��6��M��6�qЍ�����뜨�M#���`UP�W���7r����ҟ\ܶyH޻�68Q0,I�ٸ{a\2���%���TҚY5Ԥ���J�iW��F���9{�U���F��f��\=OZ
�6�9��$�aCx�.ȥ��R�6nv̝�G�&M���'�c��ѼG�͠eX�@�7�uA��m.�!�`�:c��ƆhWJ�u�����v[.[g(�i
�{���	�Gz)G��w��ΒnǮ-D��o.zfvi+���_#�Xi�}�q��mw+e�	3��U�u���B��yZ�C�F.�rP���&�Z�u���ͧC�1n����<j5
�U����,e�������Պ ��D����R7ָb�gn.����j�y{����i0ڍ�����{`��|(J����¬��ژ��pm���y1�fe��s�}�͹��mL�\]���ʳ��l�֒\Z�d�#<d�:Op�:2�LרKTs�u�E�WSl3���]r�Z���:a���Vu�z�`!�5��-c.�)C^�Y��i�Ko���ufK9�ĺ<컎i5��\���n[@��v6��t���y���nt���^�c��ŵq�o�#��~����snm� �.�;wj*���
��枰#Ȧ��ZEt�7:�J�Nf�Zo�w+\��U�ڻ�8�ض.ȶ&j��cKq�{��Ys@�մ;Y�4]�n�V,\u�ݫ��.�c�[˓���l�;����v1	u�ڱw��y��rZ������؋)��G,��6e
omE��'$*�ݧg+ݗ��w�3b�ԫ޽��LǓ(!��IX����@�پ�t���oXy.��$p�擲���i�tP���t�R��$=p�3��N_ ����m2Z�¹j"��|��tE��N��X]J�dc]X�Q�VZ"�e�
�}��l��m0g5�Z]�bkr�2��o���w+�.��F&��V�RO�P�C�.��[W�P�u�̭1�ś޵ԏW,K�%wuk����88a���{��R*�&+��lL�Ҫ�����*�ڛ΅�9d:Ew]�h��aF���ng	Y9��r&4���cS�hˇ��we�lV9s3��Y���3���-_vpl���h�ɝ�mN�vW]�YoH|[�E�7)-H.B�v�Ü�}c���A�m杝Z�^^�[�3_eӥ����xA�|�u��m��b7i�]�%l�����9izѵv��k�.dT�����A�\'TU}l����E:Pcy���vbi�^Y5�sk)8���!B��eS�VY�N*�\�<�u�U�qnAA{0A��#�
�!G����i����UH축��W#��K�cI�]�;md`��E��8x�<g��B���,{�R���lyK�zsC�2��*���2mM�pZܺ��guM>ѷQqu٭D��g���;��hFݵ�T���V��^=lF{1Q��\�C�������w-�,ѭΓ]0W=��d[��2J�u���v��V�C�k�M:�z[w��i.�U�'IPR��m���!c=��Y�:����7�1��)�(=�peо��>�2��x/%,��6#�f���͢ݣ<pn�ǿU�Y�`����5�K�Fu�U;����^]Z��n��	@�b����4������3�ذr{6��x��aw��U�i6�H!�|{K�fF�NjSԱK\f+b֋�ֵK��r͡��a��7��6��vVHj��'�"�I�@��s%�f�bd�P!������j1�*ܵ�0mh��rd���F����7fQ;-+2�m�[�2�GEkם �6:���g�5%��8�3eh��8ʷ��-����t5��d-J�Zu�Yӛ�[٩�ܪ�f|�Nq�8��f�T�Wh��	w������M<�yGU��Co.V�<j��kX�IR
��fS�&��x�Z'/��u`��֌��N��.��|���cȲ삜�3�r\ƍly[BK"p9�3��[��"D:���{�JUU�����2�>�CV6z��*y��x�9�4yV��7�q��]{�](히,Ѻ�i����G�iK���f�[j�_�;�v[�6ڽ{-3�W�е�/���sh=��Ԧ
t^��׹�e����4�͛��:���1滩w���\+t�y{��mC(��8���go�Xz�Qw��l�����p�7�(������ɰ(��7~��n��a7oN�O�[Р���8{��$�Vw.2T4*e޼&LrےM]�q^X�ݱ��/�ҫ��u�<��U��TQ�.�jt�4(��a��+1���Ҟ��:�S�d���8�Mz!P���n,N��v��;>�R����*�F��r�R�s�1;i��:�6�{��:{�h��fs/v�����;���{�Ay�����e�����3Q�#�V_ �]AM��:�h�78ոƘ2�;���*h4���z�޳(,��]M�͒��ʵ�\S`R쬧��n�K;�h1vw8���|����Zvw��aU�����qꃚW~��\.�o^*$��o��[�T�I���=#7�����A��h���e�\��d�d��H�UwJ�nwd!V�<K�zA0��Z�mY��!�M�ko��^��c��;1�U��։����������-��{a�Q���d��J��a�U,e7b����1?�k�J1�\t�2��qw�=~�+�A��0lv�운�w8U����c6�5�b�	Jթ,wl!�w�G
���ir�l_b�^�R�ZǕ̈��z;�B�ک�px:�uJ�Y,���v�l �����tdu��{��tl6�"<U<�x�����4��'u+�Ϩ������A4��\F�dN��Un���O, ��%M{uI&���+.Ѩܶ7sX��f<�8��B�d\����H�n1
�7[ѬEyLm�E0*7�R&�)�!����1ֺ�L��8.�:�+�K����CX�|z��;-��s��T�.�0wg"֥SLb[{ƀ�\�OT�x\�l��9F�t�l�`��b	,�gT�{r�:�5t��ǜ��Du�[���l^�#��W_�Ê��)�Y��D)������E\�D(#:f�J��P�SbΪ׋#�mf�zC8�a�:몮�X�w!!4�2���RO�v�������J���6��X�G#7��9$�Iܧ��!m���=�;����	%� i�4�B���ˈ�l(�~CC�8�<h�eݘ<��@+4Xi0ZA �!J���(�F�&h�@�Um�E:T�:�Qz�94|�>���h ]Dh'R��� �6��5I�'�4�t�Z�(�@GMQ"��wb��F�����OÚg"mPD��ɂ�D�% �@B�t�|.��Yt-:J��$4@��l6�0�9��/Uz��������>T��|E�w��	�o����'�}TD_�������W����<�m���=�<�'ǝoP�sJ�[U!yҜdVnVq�nx����R��im�+cw����}[R������N_S��]zj�.ɬ4mm]:��Ɍ�H˳R`��h�q���4'qqt啌��vmo���0�B�ZΠ�|��.�J���5Ԛ�ːj���Sh;\�4��-I�֝,xx���Z=o���ܻ�-�B��^���%����!h̭ұ�+������(��O&��w�+�>=	e�T�̯��uQ5v�	JVn��f�	ּ�1��YR��ΕZ���<p�y1)3H|�Z+����r����s���_Iv6��7�<�������C.bL���Z�����>�7�m��WW2����T�.�wN�2�̬�W9ҩ4�\�2ee�!Y2beǢf�\i��\R��i6�g!}7������[+xkw-�2��omu`���i�N
X���Wj�l�uH
���Q�.��(;p)jɭ�w�`
έ�eʕV�.w���(+�E�J��Y�wZl�2ԙ�nA�_"�^n 9֑����wo�݄fUF��Q3��� ����G�pU��'3Eר%vp�:�B���ӓViһ��o���V�\9\�)�u�9�|�m���3���F�K8�Y��<�S���i�A
9�V�Ke2��V;�l�{Ef��j �T�s�0kJݍdac�2�%-��H�غa����Zsf�$ų�0�Kvtq!W#YU�v�l�;d&�[��"`Cɹñ��R�Pʑ�P�{�[t��Sk,�
�d�F�,!6�=�e�;����f��}}��<'k#@-���{�Vs�G��L�q��w��Y�!��.2	�f*��e�$4䕃rԀ��yBds��e`��6��}n�zm_�<���ix��F�$�D�P��׳O;� ��,�J(�����2o
ِtf�E�_f���㼤�d���vkt=eE` ��rA��Uӗ�e*
��z�,^XB��v-83���&K��*�sR-JR�(^�U�E6J���|���ܥs��-�3�Ƙ.%C7t��낌=A)�k7=Vc-𭺙�|D���������w�˗X�����,���:�6ob��������z���¥n�C�z['V�\c�Lt���fnt�n��Yh�c�K��l]�%on��V�k1�4�S�;Z[0r)2��?�XXO"�v���en���r+��#VNfc$�������5��=J'�I�'V.�eM���������n�����X����x��ɾ�2���	L�F�w�2XU���ܕ�[�ػi��
.�r���a=���7vj%�4�=]@A�h�ĞZ�\�{�V9�tr�gn��hܼX9��G���C��R{W���۲i��2���w��x�ݬ:�4pQ�o�z�(jJU��x��w)/�jr%���ƝJ�>ې�ƪH.�Y�0Ͱ�H�AZ�e�����F]��ź�tV^�T ��fά��\"z�+I�m��񵊥��:,q��md�f�Ѓ�B�5{��w<az���iJ�K�ٝ���~�Ǵ� Y
���'L�T����o����b�&:�2�r�u�!2hD;����Τ<ʇ0з�9��2��ֹX�-ܪ�y �zЛZ�T���������P������4p���R[f;it.U��L�AWX�<��F����.CAx��h�i���P�ǗP��~v�ʲ���<�)��Mnv�S����.E�\��*s�Wab��NU�W�Z;���f�ܯ�u�k���U;� ���OVIt������p�l	m�[J�z���y0������*YI^�1�����A
��qP�\����p���Qw؝�f�:!�*��s6��&5�W�(tt"P�����qa��ۙ��G:�k� &���wt��'%-�6u����̂�;�Z�`\�J�ٶ�^�J1����q,y�]ۥ-��[ۢ�ki�1��֗[��p�(G1�F�Nb�"�ٹϒVs�o78i�îh6$81*W_.����L�r����6��N�mѷL�2����SI5�uH�c�X����c�Z�t��Sn枙h�J�QUԨ�SO�R�mä�i2�Ṭb������ W���p�K k*��saݝ��w#]ݝ�d���=�r-��%�KUH-vY�<�Pssv���u;2��`I8����״M�9{L�'6�.�'}�Muv��ݻ	K:��o;{{52��N�xoiʓJ�����]����پ61�9fD�A4��ёƲ����:Z�3��&�������7�WR�06��
�3��.���&g��R��i̙�r#�(o7j�YU���� ¦T�`í�&��"��W��	�� ��ݨ���A�:p�ј�\�S�\�B����K�-5Xl�tR'�������g""�e�˸u�S���3���H����q���%��m�5����-"8�>׉ѻu����P�u�<��K�V��Fpx��yZ�$�bϹ��.7�шoS��*� nv+I�}����5���4a)�����\�/]�V(=�'jG�k:��R��r����rq�**�u���f�Eb<]_����kr����P�P8���U�!��c'9|� �����c�+vӚ�Y�R�� ���o�H`ht<�}�KkvZܪ�{���n�ѫ�(�4�[��w���L; l9�.φJ�H��ܺ��9���n�ٜ�mC��V��=�l���0���}W���:��nb�LB���ڤ�ⱝ��ն�S�3����
���uJ�l7r�D��/�η��8՛̳�]���[��5�pʊ��
h�*�іh�+OY2r��,Udy��Ҫ���N�+bM�q���8�����m����RȦ<.�l�mr�]���	v<�r�3��Zn�d�{#`�N]֝p�(s'F���*����yҶ9�r(c�`�I��d�HH_ab�vF��+�+��PB��[b��{�z�@��л�N�m�]Z��2�l���a貳y9l;}YJ��}mj#.�.�g�/BWÕ�:<�d�nm��}�goX��Vͫ-r�fcjݕu��0��u-���-���;%M�ѓ���&�
ɚ�na"Z�6�aP�/Wun0@�\����坵�ոC�����"9��nN��{�ז�{�ˉ�p�kU��լ�.<6\� oZֆ�U��w
�FŎ�Q<���rZ�q��_bF���*�먞�7��I��!�{v���0f�7��V�T-���s��XW	8�K��;h���Ǝ
�w�b�����&��R s���`���܈9-4ێ�Fkc�WvЌ\���*M�M_k(�-�-��2h��e�m!;7 ����{�H�3�RT��ۛ�G\���|ѝ�{0�բX���^J=#S��V��tm,9�_`�H�� ]w�W��=3P�� �C�Q=��#rJq�����KqBG"�E��w�ҙZ{)#hM�C�ۏ:XYƚh��8��v��tɌ�;Ѩ(I��J۷�kQ���U�B��0Vd�h4jVC"���yVd#���^F�4�w�~��oT�s
��r��;�m������U�����K+�����*x�@6KO62����}׃��PK�b�e)V�n�����yW�7p8Wd�)�0�=���K���{/k�;Zה��atMD"�\Slx�4�<A*��h-��}�]L�FZ
�o�G<'7a�H�⫼x��@n<�ѝ~�lT5w5�0Ҽ��6�ּ۾�	�Z�֪��yd��Ӎ�.
�	��>V�'N����_�[��!��.�*(!�p��љݙ>�����Ӣz);���Ms�S�1�1`Q����e&)��^Qϻ;��Ko�����st�`�{eٗ����9��d����&��Bܩ��;�,,A*Գc����l[.<<a�!�)�=��LJ���(�1B��C��N��bR����캵r��պ:��RVi��KĤ�����7	b2�YwW]�">�ti��{	��fJ���f����{u,(��S�ې:�v�w��Œ�V�E�*�+1��`�Y��b�U���)��7&,d���ClR�c�C����B3��L<&����k+5�B����65�����gh=(��Av��N��Q�B��uR�3�V7�ϙ�5�Cb��"�U
��]6$xpm�{���<�i�u���ٴ�MJcv�s-J ��V7��5��B#eIj������q�5�㭽E�����J�]>I@���\`h�X�&�ؤ�zH`����҇Hɸp�y%�0a.ۑ��P(�Ǝ<m7X4�zku������,��GN����[�������;��e���u�E��iI�ݍ��T)�K�4�.n:xe	���E�.���G#CGF����'{���%r\��ݖVPc �Ҫ@�ҕ�Tm�]�YD�꽫y�J�M<,�ݜ��J;��`�[�d��������"9��Zp�C����oL�'s�Z+��mE2��kúe�rW�5X�:�:�:Rγ�pG���-�[�&Vc&�Dk�7�����r�B`�Ka��W���)��!�Z�����B�:Di�fS2J��ΙmZ)��v�,+�wT�J��U����Vt��Y��ͪ�0*�s��2i˧��Q�tG8�����J���RS����/���4[Le��bZ��7B�ۢQkuo$�.��r>ԝ�Xz�z3�IV��W|�3�{�񝂱�ŗsBHΑ`�����d��f���강h��7g��; 
��IG%�wV�Ի7����ݗm�3m9�o;�4�iW����t��ʻT��%�ȯ�U�{.m[9�&{�6�R������~U1�!:۩�� �J���[Y]Ŧ%oJd�I6/kiH�ѷ����Iq��''os�e���sR��=n�p$rP^���N�P]n� V�6��"�(��a�w��,����:딗�K��E8�1Փ�D��٘���Fj��Ic��XUg�][�u�wQ�~��f�;;Sg(az�-2���J��K��SWaÛ��Gt�E�;�8���)�Z[��j�g-_yaQ�]Z_%b����ѵ��_p����)�N3��ե!�������UA�J9m��$��.�n�:�����Vԓt*ʭ�2���f�%=2�K��:o�h�q8ܩM#�.�Ȯ1]�6�ϫg-H`���,�޺ꪷ#�F���)�ΓI.*�t�����-�.M�[��:��y�,j�Mr�Ǻ'(��v�]����RQ:���K�c�ުJMJ���;�����_]&;6!@l�uk��%��AV2M�P:�M�d�n���Wn%�:���I�q��Wsb�u�;Ǜ��Y��Y�
�O68Sa�.��nգv(��
b��jl��cuռ�S�Z�f�s���$Ý�YOFg�٬��j9��[Wma�U*�$�v��$%�X���N��V� 9�ps����.��-伷$��7��GE�wtM>�h}7I���b�j��%�c��KQ�[�����>��-d{F�84������pMm�=�˪V��!��w�1[X^�'u>��#X�yf�ꎀ�R�})��$��"x�r5��pyW�[��a����.�f��RZRɨ��b]F����`r�fU�XC��g�����7�ֻ��ņM�����X���׹QzI+V�6��Vvs9j��}596UQ;�0����$�v�s��p`b���|�.�J&#;O�AL+ӆ�ǌ��jng,�ݦ��̞�']���p�r�ˮǱ8�BR� �8^�g�F�O�]p$�F9�Ja��ڨ��uSmr�ϷGN:5y{�;w{�A��Q��a���Ol�̵܁��{|���{^�8͇���8km�v3�t�#�������o�F��SI�7!�ڨ�|���0Zb���We=�7���m��2����������pU�R̩c�󹫺nۋ��_Z��L�o�����.�\��b%`�w�V����(y]��k�+/I2K�5����{��O8�v�Q�9*c	5x��<��)�ކ-_��;����K�'%�!5tǶ0�ma������ɯK�}S1���vފ�l�/�)�8=�oj�E�:'z^�5�ڿ$��K��;��-U�3N��]�Go�N��q�Н-�C���6K��%�;H��>�tk0��u����]:t��+/�!B�D��x�ΐY��=��۷��܊B\��v�B�3U,K&m��y�-�������7�Y��P���W�ݾ��\�{w��6����*�����K0k�d�y��컵�m>/17*��4,`A��l-�*�u9�h��U�3N�xqWqNN�	��-��m�|u��Wݎ��D��4ۡ�4uU�B����(P��dɂt�,.T�`��a�mة.�^��Wy ���k��J�D�@�iWǤuY��Ɠ�R����n9;�a��2�@��HM�6�`0�
��I�ʢ�{��_U��]���	���oFd���t2gg@7�M�򧠠�d�C�i��EG�ewS�.�s;q��m�ZYp]͓�gv��ӀA%+Z0-�}Kx��S�-��Z�؛E��	�d�g+��"��	���5���Z{`��d0��S�s��7�����o
�*.�v9rk�5뮹�e*\9��z��ºq+]^"�u<���`��O���G1�L��\�����'"骄ˁ�:����Ck��G�Ҷ �-�[�}�o��h|> ��}�x��������~�~��_��?�����~ϧ��}>�O�����|�_/�����~)(�_>�=��n��&S�B�m�H�b���#�.���Z�ߗ�?o�GL*lc��[:� ��,�*q�j%8�t�qW�+;Z��ӯ���9��w��-�rZ9�C"��,M��߯�FK��o��wsecΖ��*���L�sS�����c&Q֕�v�
y���Gh�Y�T��1�z׶L���d׉�����I���|Vf�ns�K .�������'2F�З��C'r(�9's�܈t/{uYh��}���T�o���8Tٕ���,v�����1�0�;���XP���
�*m�{��3%5xyb �؎ ^�&ܽ�-�I��w;������XA�e-�#YD<�)��mb��s�a�n�OY�)�~���w�U�7���`'�!��VT�Yk��AK�y�X�%ش�u��osy����Ԟ�*p�VI��k9��Ԝh�K�_lp�Uv��o'gL��#qii�a<�1���o_d����3�r�\���U�m�]��SW��J���m����T�os�u٢Y��݈�t�<���ݗMTn怒vmh<C+�t�"n"�r]v3ݑ�\�x��LQ-��N볘Jfo�����N��l��-w!-oL˖�о���Wg$�]�갍f��R8�n>��ػ��M5�0�j��o}0t�#�1y��Y�G��m<U+-�ٜ�VSv�v��-�1F�A2�T`"!&��t� � t�t�����4[h�����y�Od�����*M���Ӌc@kUb�Z���h�U�DPE$�F�m����F����
�f&( ��*"�(��*�ړEE�V)���f��u�)��*B����f$���`��Cj��&)v4��*���"�UQZMNÂ"*�j�a�i�����E55K[b�
���3�%E����a�i��Q�(���fv34�M{�AM-3��EkQT�5N��m�j��������cELb�B&�����bJ�f*&����1�'Fj�qQQEm��"!��+cUD2��E����Uڨ�4��"��DESDIEU1S4PkETUX�EMTARĖ�1U�M�PTT�������|d|�����U��Q�9f_-F���^���o�ٜ�0��'>ٲ����-�*�{5|�fb��v�J���i��M��,uU�%�Վڌ *����v���	�;d����g�.w�j���OݼZ���������#>�+�\1c�O�Ǥ���7ݞ��4�ܸ�Wb�2��/s{R^;�"��x����p`�,�$��� '���1�ϐ����F�m�gcu�;�����9���}ưv�x�Ś����$�tKg;n����ɋ�7�O����XݸJ�������5��̺�.�p���˄�ι����O�~Rމ6m�燁�nA�|��5y�v+�H������~x��x&�Ċ�v�'�	mc�Bڥ����Qt���"g|�F7<�|�t@Et���߶{�����6��C8��b�~�˓{�	&�F?}Aء�M[�s����#�>������Ӹ �u]@,�q���{N��9�0�Y���5p2��m�'(��翁�z���_`�ؔK
]]ws�eN7������e�lq�m�*�Ncر��{��j�ͧy� <j�����nE��1aa�\i��{&f�>����Cu)9��cgU=/s��5�m'Ԃ�k]�B�%3[�3pG{mK���t���C"MM�r8��D=�{ �īzg׈�h�Ԃϙ_zE��v{�x*�z�O˴�@�!�R\"����Sʿ�%�f^{��{�����%_{��6cˁx�Y� ��^�8�niʰ<=���"ӏ�����B�t���X;��d=i�<����VWx�u��>Y��\z}�)퇚�C��~{�؊�����3�W�2p��yfo1���ܫ�w�>��
����!��LQ�c�������n��3�=&Z�:ڷA�]�թ/6��X���=�`3Ƭ1�[�84Y�ߩ��3f���^��ȧ�I�9���l��>�`ޫ�*\	���<AC��徕���y�8���#� j�&�ɐI5A���!���� �����x���[C:ԑH�O��S<e���Ox����,{�Q���U��^�bO���J?mj�	T�j�J���gJ�����7}i,M�*5����T�kg$��G���z����O��]f�v��]O��z���/�ɍ�)��Cw"��À�dȨ�i�#G�wu��5v[�Ђ̖�����:�WJ���;:HNl���~u�F�Z�b�,��͜^�|�	;�ƽ&�z��i��sD��7�*�2��Q��zg����K/N�kϻ�����46WF��.;�ߣ~��V{���r��2�������̊d=���'Ի%¼�&�����{�C�|���WPK�߃���i����v׊�-)��Hy��g����Ǯe��d<����=��f�L�޸����D��-4m��ޞ���Z$� c��_���;y�zX�6�sg�4rx\����t���茽l ���Cι*XN��d��k3�j�my�����x����vOAz�cg����Oz�J��&g��p�K�y�Y�6�w�@lWw�f��g��+�6j	z�����݊���ap��󋇾M��QzW���ȉ{o�&gIf���ty��O^�/2�.�|y٪َ�n���׸M���b�E�y2�-�����:�y���XH��+�����}���"��TW(��,I�ѧ\�F����:^:��z���^��ژjf9JB1��\\�5ɣ
ud���=g������:M�K/�ni̖��4�4�m����+���zٟ2{�޹ü=�8d;�c.��t�-#�<ߺ��s�Cq��h�qL�۹٨�⭬`��Mv�w,;�ϼ�~z�dw���m�X���I��&�'�[$�P}�;�읝
\����P�w������+���}���t�H��'���5��P���'#��Q�>�(�0���j;�.�y�x��o	;���/��q=��^�l���>���{���b�)������1v:;aNKDQ�|���s��~���Ob�{�o�ʰ{�e���O�A��9�u���/O���S�w|�*�^X�w�zx��ܲwTP���'��GgvT�[J������p>�-ݟv4��ӴOuQ��v�y�F�m�?�]���%�ί'�$ƾ��X�I�=�ޜ=oW	-�����y���V��R>yAP1q�9�l���uw��h(3T��6���'�m���w`fDh�a����KhM�������:᪽̮�����S�MΡ��:��U��HF������W3��{MPPWq��+y�Lv������ ��y�MG����$�A);��RFy22�J�yW���V����{�l<0͓ �3��mz���v�ՙ�w6�{��˩����@�W%�o��HH��
�?6,���n�{�jƽ6���K�)�="$����hB�"g�C���қ�
(?|
�;Pu`����Ͼ�k�fps��<h�|�O	��#b���g���@�q5%ˇ5�#��7ݵ;XfL�E�G����8�M�@��ͫ�a5��rt���"��y��^劒�l�7��ڧ�I�h�M�X�Ld�.�[_=�z�^~�$7��~n��'g����gF�N�A$�l��z�q�Ϯ��{�T�s�kQ��N����V�=�w �|�A�������د��1��"�ޔ�W:oӤ�2sCU9��.����ᱶ�;X^�;Cj��̝=��L�d��&Ns��OO�p���-��O��e�O�,�S��HQ�i(>J�Ums*��*��/GvSY�,C�'`R*]Uմ����8qY]��@*R
��z%�Φ����w^�t���F�d�6�p�F��Ӈ�ΛU�rV9J����ujc�q���϶��YQ���l8�+	�d�MH�Ǭ������<u�$�;D�HKl�`�����x�Ճ_��o�~��q3����=�ۮt�6(�O_ҽ�~S�<J���Sm6������?:^ļW��c�v�P��={�^!��r�)��zė����Ѩ���<{�2�E'�d��]���u�@�^=p2�e��x��T�3gz��zg>�jSرɞ�[��#�ҁ4t�DJߴz`�Fr��C<��K�����ɝ��zT���x���I�"4>��K0^{���H~NwwOފ{2�-�������`f]��Б�8c���b��n���gt�����`{�{��V�F�����'�?���UYӖ�3�߇`�Xv��'��<�-���l�=ܚ������E��Q�'����3/+f�Z��H��r]��z�0��b@����h�6MFD��w�G���!5��w�7\h�tn�Y�}1�Pg	�RV��c^W"GcBL���uVfmV�J�4mZY����m�}����5ԫ9�+gy�,Р�j���\��,���q;�9I+�;&1۹���j�2Ռx��S85�on�\>.�oK��s���&j$dX�֜q�=}ۛ~\jǇ����*���g�\K�R�\3�.>a��c}�$��M����۷�|��*�z�|���}����۰�=�=պk�h8x�tm� ��$��oe����q��sH���"��Q��6�d��:��2�7��"��x�{�(ؐͣJ�~���z��E�z�׺>_�"����D"�p�ןC�$�?^�{��^a�BQ�}9*�p���g�9���x�<�����>��o��f���v�IS��a���ˡ����}A��X�1�}7d�ۼٲ8�vͪ�y9�ot����SR[�:f�.���=� �<'��SC�ѳ�W�K��
�����Z��ٶ1I�c�Oԃ��ӶO{b�g=w�o^�#���hoA����{��1	R[_F�'
�(���6�w��VL�I2*qܿ��3t�ۄ���r�pz�D�-v�^E�߽���P�Gs~�n'۴�@ϾV�s�uo�9�v���Ο@��,�_/�m��'B�;���o^����һ&�r�$�k��2p�N'}Q��-��Ť�]�}�ы,.��+-�T�$";OJ�*TX�5�U�Ņ���K�W=���d	��Y��t�<&k�V�����~NDIjP���2�1w������3�
=�q����U�/�$q5ס��{���x�w��6_<�:Տ��g�އ����aߏ����1�pvk8k�^1�<�'!�CZQ��z��j��T�#��'wۧ�0<�*����ޭ�'y�9}��*�}F���;n��4�B���2b���CX׭�G$�7�=���,�!����'���B	�U̑�Nf������{]����F��z���`F�ϙ;�m&G9�	�.I���o+9ļ��Xݔ�I
Ώ:��^� �p{>��N�o}���z{��Ӻ"���R���{���8�h�z�����ӆxHw�L�d���X�w:ɑ��N��u�
o 2R���<��<<����{6?������!���5g���	�}�ܸvw�V�$�L��9�y{��E���n�=vfƭ��1sEU�45�+72�F-R\�m��*q�Y���wϢ���{ί�r]�c�]�z��k�V�WK�ۮ]]�-H4�7�+{b}���o��^f	��s�>��O%�|��@�f��iƂ��mp^@�s�t4hje�"��/̹k|�v�}��?=����=�v�C���x��g��yy����a���l����'7�N�;��zN�k�B!��K)G�g��_{{��_w���$�᱒O�;dv���T��b~�M�,�^������z�������v�d{a�Y��>V��$כ2K��<*�t�sOʱ�3������꽋*�&bU��Y�І�?Ygv�ב�I�~�{�����x`~��!���o�Q<:��{֭Rʣi��nǺ�K�����x?'�_8#��~� ��ߞu�Cڲ&��-a/�.RZ�_�w΅)Rd���f��O.3�����OTU���n]g�/L���+4G^����x��=���p`H���,a��BO{~��7���_\�ֆV�YO�
��ψIS�B���d`,z~�#�>j��	����BxK5svXNXh�B3E�������6�]B9�Bgo	)������m��(ի[����f�"�Z����lє(e��+A�g�u.lC�q��ĺ�����ך�𑚔��K&���z�z��=��;�<4���pz��zn�t��&�}�g�LN5H��:���j�u������A���߰7�7��]^B��q�S�o��m>s�o�������# i{��V;����g�\�~���\�@��6�&Ns�tv0�%�A6�:�4�z�v���]���?o�y{}�/^���=�zzI����pj��n.�U#�{��xOC6>𐀷d�h�.���/�~�<K߼]s���*�oJϹx�=!*^�K�}C�y�	b�OB�^糽���#�~�����*��gL�q�'G=����ë9�X^�p#�"��3ޅ�;�w�?Z�x�E�8� Nn�{�Ќ�4T?AA�V��x�X<զl�W.V�������$׸~C �:���
������/���}ߣ������z�������|}>�W��R�o�P��Ƀ�AU�r�6�%f��l5U˕j�ʄGE���V^! M���=���ȴ����*���>��^�ʸk�;Y7�-���Ew�w�VL��8x�;ژ��(�̰ʎ�i�#Π�l[�R�7K�뱵VtG`���(<�;��!���,0�5n-�O�z­)��[�Vk�ld��.�Sn���d�W;��Y\4����tRrx��g4�.��̔��n��:v��#��7w�@�
^�����;��u���/GN����!�;E)�t2���2G�ea�eq��]���&�6F�y�ڹ�k�.���/F�]���P�߱���(wG6�Gs��+�A��c��U�re[�:��'��J�r��M�N�r�f����VG���xF�Yc��[��!S�re+�FV!�iᗵ66e�h���s��ZfU���O�eM�Ls���^Y�h�b&�5��e��ؖc$�[�_�J�8:�����Le�=�!��A�P��Iep5��s����M�gm�cu�St�ܤ�cum�4I7(�&wh�z��D�{n�s�[i��z��r��N�2��Ѯ�Z��V��Mq����F��Ě�7vn&��d�z����-�\�Qԓu˭�@ok%k9Q����!J1*������6�Sm}WFy�7���wf� �������ܧ�,tr�e[�Tf���������7f3���K��\��E�3.vX�Ȣ�Cb��B��*���ٳ���b��|���D2�����a�,Q���7�N(G��T�.�2��0������-_jtڔ��� �w/9[6�>�܊�c&�룚�j6�P��(�4�.63+���_n��rE5�ߛ��dg����*�#���%iEޑ�{"�]f]���K}�6�S�:s2#e<Y,��o��!��yk��jsʫ��45C���9}����j۝��UJ�>���x����
a�Τ�P)=��̫;��:ͨ�<�Q�G�����]](�rR�mD���G����mI��bt��s��	*ͻ�2�ǎ �ހ�P�n�,�U����QV�!��ni��tRSƫ��}��A��c����v�dP�ǇI���5�Bʳ�N��q�K1�x���8Ϋ�vn�r�0c7��wA��;�WGMb����x���,�sf;��tޠxJzb�S8�Rq���Cد�[}�'"��99��2V�Zr���C�X��ݗ��'��r"��&Md��;��PS���L�Wvᮆ��N��N�Y	)j�酬�[��G�%:��
s�Le�bRKL�V����s|�''�b��t�ڗm�8�M!z��j�2j^m�R]ʒ�؛�o-^��L���T�X0a��VZ��x$�U��s/7X�;]�������D�vj���.ǌ\l=�s�F��1��EN�TU50EP�PQT�C45TU1bf��fv��E$DAVڦ
j��"
m�ED�pf&*֒�"��ڠ��D�DET�4�T��QTPm���HQETMUUCDE[��j�h��lEE!5A�E�:����h����B)�h)��*��b����SRQV�MU�EA3�"�j�:����(�H��SMAD[�m8
����lشE11�h�)���tQ�QSUEQTD�AL�LQUShֱEN�j*)�H(*�f
(� �j64Q1��j��Q�.U��/#��T�X�8b*�Z�+�71�Fj��\܎A͠�$��m4E�ns5�sn\"X��Tx2bїZ���FcDh�5W� �nnq�-�ѬƜnc��r�6Z9Ü
��p�m���y�V�ME�ܹGbbbѭ$-h��D���x��������O�>��UOw��.d�;�gA	;>9�Lq_S*���r<�y�i�7b۽���kw'K;��k���7�s��v�	��ϲ�YrBh1�7k;Ot�H�D�&����k�����,������[9����w-l�04��s�T^=����w3Ez�KUHC}�K�y�m8�3{�;��1To�Uƪ�~�8�~�P��5L��	��Y�R?>}Ȋl����la�Z�ld�'�F i��1�Vn��3jj�"��h
Z��ȇH�x���=a�yq��
@�	p����D����e����D���n">����`	��J3�+ǣ1�ޮ=^���>
`xav"!�V�!������:�̼�[�ϝ��y�8'�Y'HĲ2�&����|j�t�On���Ivlo���'6�U,X{wT��pH�+$�A�$�O��Juat�e@$�5���6�Eê��YM���T�^��[U����w�3�G��L'���2��.�����5�|s��n�J���j&0�&��溫Z\���z���@�`B=�smmO���I��T�H!7K�1i�g�H%�w'������t�Sd�VFޖ���7��[�i�`��_�����a�kO�����&��ݪ���"�}��,֠J�~5>`��GKN٭����C��s:8���w?X�M�����:��ļ8B���-�q�6]q>Թ�v�[͝'�z�R�7.��`CeΦ�+�ỒfZ�L噪�UN;`(��=����ZKd}��v:������uѮ�3��7K�oB���I�wm|gaA�����}����\��O�1 7��d��_L0"*g������9��G���B����02Q��,b��:)WQ����U#�rL�_���?��o�}��=�N"��u����������GκR"��rV��G��߾l�(�^�������C�}�AT2|����k}����%�O����9��r��w�n�CB�	�q����*��S?�F3���צ>ǜ��-��mr��f��0�[}���D	��®���3v���/e�?Þm�X�@x{���4��M~�뮏��+W��� ��]��vigͷa�T���j����b{���}k/��B��`���F0k{d_Uϫ�v+��qZ�%s`Ц}�3f��w|3��>�1o��Ԍ�=f�2��-�<�������'�C�=7�T���WN�R�{��Gg�wޕ^����|>}ka���S$�m�|c���Qp��@vA?����K�7Q�Kv��� `�����vF1�}��\��X�	�N�؍
W�T�P��}b��V������e}C~F܈��|�ͷf�f���Z��Br��ù�'ϋ��H��sF�ۅ��]��x���<z��	v�hZ!%Z	K��}���6V+tSog5t���n�M�ԃ�M���u��۝-��c�`�h�"Ťν��m�I��Ǖ��P��h��"A�����\��=��_s�f*h��&��,�^��v��.�$vJnf�L�ɹ�Jt��H�U$����uι����;��oNnZ�i�hUӍ�>5ÔH� �S[,�}��=ԩ2�b��}�m~y��`o���\��U���/A�/N�o�=��+�!�!�k�8#�; K*�5��<��w���{�o^��zZf�X�4�->G��ٹ�����!�A��t��y/��q}���Q�9�Vv��9{:��p[�����礠�<�����D3G�!��y��l����A�����c��Y{����r��t2��i��H��bN���,(,��Ua]k	���sS��5�0	N^�R�[19Yà�M�ljg��uH������Q+\u��\����֪9�$�:�la�ɺԏ,gf���==���q�DJ��`�y�ǈ1�"�s[R��OC��j:�O�i�n�y(f�R��4�UN�W��
�a���\��v��z�{�|e������C�kz۬eK2N������9E��|�<�[EY��$g)�m�f�t	�v�P:'׺���s˸'CDay�����2;��{*�;��i���&��([�|{�Y�ۄ��e�ԩ�<3�![*�����)�Sj�6�z��l"UD��_P��)(�����1�k9��V��R�$�5�\�u�M���K���W�{ڦ폳��Eݎ�}[}�Sww��zJ��-���>��<# ��Ty�C�:"�7����m�`L�_�����hø�����|�/Z��-�l����� �r��ך@��t�P�Y�����/Q��˫��,?'"�k^e�ƕ���kj�B��1tR�PJ�g\=�N0��E�jjb��2b�D��u��(�3��	�Ɯ�G;O��2Q�͡��M�L�&P�^����rXU?2��Y}ZKN_v�~������(A`����i��s��ا�������G9�����c�M��M>7�L:JE>E����{lw�!Ŵ�� �����Cz.�Zq���N����:��ot�=Xl��/#�+�1�K$���RJ�
~���s���3d� �.pTҝ�w�3{u'��Ýۚ�7W47�9ye(x��M�L-��ye�H�̹fo�`�@���{������O6��D��VW�mLn��B���*�*���dZ~k	A`{T�~j	ĸp%�4j��aY�}�C�҃M�0Dkjh��jq�jNл%P^���uV��g����2����_���/c���l����,�n��/vǶ��2aA���PĜ�^�)Vԅ�.�K��
�tˬ��9�I�f��&78�$7��h�"� <\����o�^'��be;)�n�����k�,��%�V��{׹3==�M���Ʊ�:_r�e�zp�\8��k,:=p�_�bXZ:����*��ҹ���Ƕ�R����3�ۉ�uo~�=C���l��t(�>��	� ��;k��NT������M����C�j��zGusu��T�s��O���uɈ� ��1&,3ߜׁ�����=�ξ'���4L�:셋�6��6�a����Y(�ZQ>��f����W�lZ�X�c�� lc����ͼ�d�nM���nv`�<��{�Td�4�ݬ`�=�HrC�7��i�[�k����Bm���rS��8g{�S:���'��m��^����P�m�*�Kx*�!^�%�;z�2�.T�Y�w[u��R_�(����WK�������d?]H�ό�nڵ%L�c�ɼ���C,�]K��{vi�u_��p�	����~年�������\zxT��؝�&svv^ZӾq{�U�Gne�LP�(1kF%?zQ�aG�1��[=[�z��xA@�!�[�$8:��D�P�Me��MցzK79��&%�{H�0
�%*Mw����{gN���|��/_�&;�Ϻ^W��W{�{�Ct��U̎�V�>���3�uF�[�J�jL3�C�u�����8���~���49Y
f\:���~�z��3`�[���N ��k���+�n��Fe�P;ݦ��Rԡ��q]ewN�e�vGD�7W�f���yR]�In��&ݚ�	�ȴ$��C�zi:����]:^��"�$e�������mz�M�|Z{��La��^^"�Za)fT&c vK���vI�;��]��-:��%p[E�0��A��w������^vo=�[MhS�·���y�V)m~��H�+���Q��w'����)������LZ~O�sn.�z^���]J/l������*���0��1��
9�#Ѣz���\�7۽�����&��V�7;szg{�N���l�~��3�d��qo��D��y�H�X��]R#��IS����Z�9r/�.'7ig[rڽ�Սv���b��6�a\���6kӻ6�m!����76�=��w'^"/�g���M�r�j��[��(�����7k�>�{��]}�=���8U�C�!B����^�d���E�� �f���#�a�azچ���T#����ߓ��H�t��W��~�?C<\�R��U�	RG���p��3ň�v�&��8�f<5�ݐ���� �4]��b�:�U�WE�ȋ7Xbc��wf�r�Oȗx� K2.9��0���m�87�љf�����e)�����~����d�U�,tp�o&(�����m�xF�q�����E޻Ǹ��tei�ݬ�>#�����>C9�B�#?[�ʶ���,0�����l5�aYK]
Or<͓`�t�r�M�uu��mUu6h΃+���v��.��<��w���Ǜ>�QF��@ ����IW*�7x����c��a�l^$�·�����5K�X��+�M�����l�ت��s��u!teъ�Wڻf;W2�jdԕ�A# c=��T2���zw�H��o�@\���3�����5�lʐz�9�i��X�  ����u~Hֳ���|j*.��f�;�Ce��Gc<¬�z��,R��.:����T��#!s�~���8�bS��J��3y��\[ ]�bE
�a�4z\N<v��{]� ��A�k�0���r]��#�Ss7:d���%:��O�:=*����&��;N
��=[Ɏ�oG���	�2�[0���s�Gu*L���pI�f����jg�%�St��$���/JF��
�����ƑB~�s��,�ͼ77��zv�t���P�������d]!�̂թ4�r�}�������kϡ�n� �ڳ�6��<�%�n5�%�*����z5yo�J��\���I�(���i�Jxwf�nC�Ϝ>6���l��8�;n^��ܭ�!5�zU�`�P�^8�%Q`�:y����k���������g�%��>Oc��$
���W���uq��2)k�eҖ��5�JUG{dB+�n��l�ɘ������+��/��932��<���������sg#�_(�%�Ә�=���������k2��-����4~q��d��*�.��{e,�{NeF���x 1�  �<�����٫�!�`k`+���&p���T�m��Bը��:���}��K�_�G7�3jMEK1!��ŝѹw+�����;�8aA�3�69�@|NhmK2��m��u*���������0i#Iz��Q����3Fa������>xs끀�����yR̓��77�+�<Ϊr�r���������+1ޮ��K7k׉�v�tE��:���yw@��� ay����F��C����;���W?b�:�T� fE��C�A!���˴�l���6�ƶ3�0%������n,r��G^;��d�]Nx�E��Qx�ۯm�2W�Ar����g�o�鳦.7��6f�-!�^j_�Q��&���[��&��+</h~Z�$E��{��j뜩kjҧ�k�A�WB�ɒ��������*\(�?��&�+�+�-�9@W�K�YM����?�3V�Z'�X�>!<�`�$&M��Wc��i���};�ځ��"��u��ᦞ�� ���H|�	��ا�:����=0�j���g4*j@7D�)A`��J��l�8�����=!Ŵ'J�ї�Bz�x�1��7	C���jv�`��5Q�pM�L��u�p�\���aG0|�&74	E�=_CL!�]]aYB�����kb�2F�v�V�ZZ�ف�ǒiK(�d��dr�7b��"`MF�s��{XJ�i���d3yL���jvC���bWs?���U;{��a� ��Q������#~fИ����`cɼY`n�e)*L8Wƥ��/)�B�_ ,x%��g�Ր�5mډ��6w7s��a{9�e4�o.�0��ȩ0�B5(���gL6���y�6�/���1��Wm���cO�,�`���86,��P�ۊ�\�y�?7��\��%ߘ	�7cf�Ē���+2k��I�m���|-}c��Jt��#[�mM'Vjq�j�Ӵ.�Td������c#z+����ܛ������-����Ƿ 8!��[�C�Z�[SM�����P��n����<�1��m�b�ʩ�Z���=��9���6���GH`��E�3�A)���d;6�f��� �'w�3���;{�}M�q���k��OO��gӯD��Q�b^�;3����4B.Iʖ���E�s��{c���./�� j\��f޸<����A"�^}�i+?�H���2j�C��X@����ϛ}��6��p~�8M*)�^�� ���b����A!���2�-Ǻ�:��7�g�~=	�?���W��m-$d&�{d��Q��Ot�n�i�+��X*� ��>��Y��5�^f`R37�5�vCyzWw39�r�Ŏ��k;^���C"K��`�]%ھ�[hs��ꂍ�2���8�n�26i�tq<��;���w]�VeF�,%��enV�ⓒ�kpi�<�
	�#f�뮫����s&da�������_��J�@�ҡ@A�Ѕ"Ҵ%--U#0��7�2 �&�J��[��������̬�_����KCͯ.9[�6�W�%L�ޜ�t��S��s�G)h����NP|ش�1���N�08��ȻӏG���	?��ζ��n�̝[5��y晇r�V�-d�Z�D�^�gP=^�3��ہ�����0D���U���y���ž�����Bp:�Q���?A	� LK$���`�J�[�[�g��<�{w �&r�uDUli����ۂP��]���[ñ���~�N��s�X]"�$�57Gd� ���1�w]��6�X��Ǯ�WK�q
��A�f�>�`� Ì�i'b��R�suK]�/w}
�6�r�Տ|��<���QG�Ȅ�^��۹�^�8S,@;	����o��ۚ��S���|���lxt5&���`y��0�`d0Q��G8��ɽ�}Y4�޳"�K�;�ٶ��l7ݹ�]S�w*c�FIxWYK���C,g&%ݣc��q�n��vO���a�y9��hռY�YݵZ�[��B۬)U�{Г��M�a\�T�e�}_�E��_w��>�_O��������{���w�����z�|}�Gw��EU�3��Ɇ���{��4�ػx*[]I?���G�b*�m,3�pa�{�U�<w3�66CD�"��v̨"�0�r�_t�Z�iQ�����t����ز�t��U�8�6Eq�A�~ךc0�ܠس�����r��0ۭ��$�ek��7�+�2o��v�ҰB}�kS����CvH_�p�d���6�<Ѧn<�,��=�j��^�d��ֵu�ln���`�+&��6���j�>풯!92�6�pSJXMM�j]�v�9뛠泒�R!M��o�-5�H�E����Y@G�gC�Ѫ�A��h�GV�s�B,	_�'�t��i-k�묦cH�4,Y|z<��ٹ��%J�ZW���G��c��)lpT��m1<��hSpn'R0U<��Ĩ\Rn��':�	�9���Z)�i%w�6�n���v#ZŶ�8�Q�yމ��j�N�������;(�;W�4����7�܋�!f�~�L�G�A���i<�o���(��n�3�/�1U�ǽ�
= �[�d��ٝS���K�l��Z�rԐ��4�/{���u\[�j�M�h��1f�,fq��N��{ɵ����{8"2�\�,]���+�%�;l��%=��E޵�q�]"�tv�4�H`��N��c
�.Bn��6��ov��x\�S�jmiُ��4�
�WN�f��]C�L۫��ġ����IS�P���W`��xޫ�@��+��o�;�b�|.'N����W��\�E�nL�롵>8v(}�Y�)�:��Nq4�.IG�]�u�a5�T��Qgi�e\����1�
�ǻ����>��	hn�T&�z@��)D��K$,�}{W]�L�J��w-�R�-�q�M�tFB®��d^5�4a����Cls�Vq��f�R�Ûx����1$p3*�4�ھ��OIڕ�N�*ݐtǧ3��W���#�ur�Ԉ�'^ :���R��*�3P*YG�#��c�q�7�e�XC���w�c,:\�,�#��&�V��.p�RT;�U�NBz����ݓ���u"km昆֭���v��Tn\yH!=j�P��h�5%[bK�V�U��ő�77S8l��d�j_<��k���:�{D
�^wwA���L�	1�|�xmr�k���mme;qJ�������jcN�o*�^�Ј��7o��3���Ggm���[{������+n�(�p=Z�C3s�öS��.�,��]mЇWK8�彔��ov�E�aHT yy�%�oM~�b��Z�3�5����B�sj��x�ˆ��f��XOD�嬡]���2��	�]�\.�k]3UP��;i��VA�ް�v�z؝�+��^�?����Q�'��V �|��Q��$Idt�j���Y{�s��bt�g3�+��5�$gl$�RQ����e˨`^�,�P A8 �3M��+�`�PDf�a!�J�NĻ^I�T(�A~��Q��dֈ)�~.p�j�#��V���U���Uli�\�.1���-TsnܢӸ�35�U�m����ѱ�b�i�p�FլPf��1DX-���ES4��q9�W#q��l�f��N������Qbu�������UE����f��b9�E8�1:��5�������r5n�EDb����r��ns�CDEARb�EgkF �j���3TN!��h�N`��Y�Ac��U�1QE5�\��2\�AVڢ��TDDTm�M�EPQ5135�m�[j��MU1m�cAAQ3�E1kU��EMM-<�r9j�`�h����l�k[����k��lSED��DC\ڂ劊m�Lm��f�"��U�TV0f�(#5Elh��\Ơ�i�����nZ�s��*5�".Y(��PAMKD������m-Dr�Z�,D�5RD�5r�TUˑƫc͢
*����#�ݍrpTQs���mQKr3͆����*(���`�,�+����x����r��j$f �]Ʈ�)���f�`�n�+XAфӅs�	j�Y�ٚP�S�bY��� ��m�r,w-����^<Tn�Ϫ̨� �#J��()HP �+H��]J/t�uyN-��3;����α�*�O���E�
%0��x�X��zw��X��������%Z��+���qګ�LC�<P�ɝ�byچO��hA�v}I����|�M��B�	E�Q��*z����ye�{�<3����&c7�#Y+&�����f����'��}��Xϼ��,��pt='�x]�%� A�!�E�4��N�b�i�{zG��7K�x׆y��,�GH�˴�
��w��)ư�����}kNޡ�6�kdS�x`0&P�a =Ų.�dtAٕ5��l�.���˧�EcXa �,��*�R3���8ʲ����N��0����R��z��6w��.��E�3rߧ"��L �Z�A=P%���ю�Ƭ��r�.�\�0�Fk^;�:�f��͠��0D㌠&']�T���\�S� ��	�N���L)�6'nظ��V�͞�˅l���վ3��ހ`�5צv܀�g�%73s�I�9�N��h���y~O��d���ǮX��&�	�h4:q��`'��C+�q.�@�na,����T�g��<N�JΊ�0r�2�`��gm��|��n���cl��{ ���]��(K�.�p���'Y�e�.�|�gedZ��[��@w������S�o��V�X7L���f���w�KS�6Qa���r��u�X���~T�X�\����R��j��[�|��� �B����B�@��R-
�@O��������ѫogM���&*ۤRz	@؃8�-A�-��!��B~�&�X�y�h�wj]�{k/:���ܣ\2��JOzL� ��c؋7�iح~�w�~y�\�o&��J��ӹ�9�\Hk�@K�~�Z�k���%s�P9r�Մ������+�<;�@����:�e�Fm�i��7 ��D@L/^��6k(Y���,�%���cH+�`Z�>�����Y���r�T�#{���K�^�7K,�a�󩆜���smv������n���	:OL��,��ö�]�KV���̡�x��u=�q �����9��,�hv�a�^:��rn�)Rv���dgp��S�P�;��R��@���g2dK�p04Ba�6߬eK2N������+m�"��������_�0��լ)��^&Y�^��v�u�E���Hfr���qˁ����Ë#j⶧w�_vr���lܖ=����{2-������hi��HD[*�xc[�w�u�T�]�m�~�����B8�̕�uQx��7c1�"%�\�rU�B��ך�i�o��7��=z������r��m�Y,I-��D��\l��hP�K5󄘶�vi�`zN���.����� �[3.�+^�A����I��s僱�(hnF�U���B/"�l��-	uX�/u����S��&d���H]u�LI��^�h޼���EG�JRB�B*��H%*%R��o�+��*O�'[����3ǴF��ĸz���*���9R��5)_��ں��r�>ɶ,��5mR��uá� `��j#�X7��x�����R�3���p��nj�Jl��d���7^�gO��m\*~G�h�|6E�� �G~ΤC��c���̦���U�6����쬚�7k8�>w'��`r�9Ϥ�ENHp���w9�^��xOm���#��%�oD�rܞ������r��ۮ6|�y�p�-��9�%:�1,���2IJa�~����s	����D�l�ʕ�$���������sЗA��4�=�a�vEM�a�]ctS*��P�F9`
�-�����S����z�A�Ӈ-�����B9��n�2$��P�)�~9 Z~kJ�Z��R�
���V�nv�w�B�K��,��?�����p�n��4]q���Ӵ.�Te��l��D٬W]{�3�[�.�����Ӈ�p�=~Ba�M^F��=+c�%�c��w^|���'O��i�ἱ�_ä��Z��q�n��V(�t(ur�������o�������.�0�M{c��ޫ�j���A'A���o�V9ok��rͻw���X�21K�xFd%vTӸ���੣�p��Yv��6v��\l�y��)n��d�����Y�:C]:ږ����'��9�D�:�>�"b���#���qu�����qq�w�����x3xa�)B �	H�#>�??>�z�)NwWi���zk���I���S�ĸ�6�f@�{%�ы�d�fq��v��w�e��f���)Ї���C�ݐͳ��E���x���	�&(zN��r�a݋y�db؝�W��{s���3fc.�l �Ĉ��S轸�t�i��F�ci�t���ӷ��t��M�]��;�0ؗ󌈘z]<y斐�-"�'���{9�C[w�F���<���Q͵nԢ�Ѫ��x޲4!�<Mzꯌ�e����K�����nv�}<��Ǚ��&'���4��ͫ��jS1X�6��&Б���F=7���΢H�=F�*�?��)�iy�=��u�s)o+��8ܱ��/"<�%6����n��8��ݾzoc�=[�oF�f4K��X�MՅ�%D��#��#sP~��ĲOi�W)Rk�Dv>5s�:p;6��P�2!Ǧk�f�u����p�B���N͕0XO�u��q ���%:O�s�X]"�RJ�[��GC�U<:D��9�szsr�c �.W���3ffȯU)f�~��v
{$Î�2���_��渽J�poM>�\��1_W[����=�(a5�x����2��i	��siL�gZ�~�AΒ)�S���]֩uםIN�hIWY��3�J	�q݆e�b���+�X�%^�ev٩��X̮���:�̴��u�SS=V�5*+���m]L����^���78{����}�*�"�҃J�"�J D*0�`<�<޾��U(�}L#y��	�`��1���>�� ���Bm�Lpmь#�K�:�n�d����Y����z��_9�A���RiH�0�yz�;��B���h#��W@��j�W�v��1��蝽X���Kb�\�k@�^id�e/A(�z�,g Ļ�z5�!����K��!TX�ɒ�d_*��7�\��M̉/�Ԋc^2k�RrZ�&ޭ\�T�������`���h�쁻���
`l�P�������"��u�����t�VZ�8�m�꽪vƼ躼*�k;�'`!d0k��"SH����6����hGP;I8)�K$@:����/o��9�Q��N��n�1�\�[�w�tK<���`�ˬs�ړ��Q}�����RFgS�[v�3�#38��4���q������-�h;��4\sO�a'W���r�{���#��o4�L�.�ر�N��5L�IJ�j�Sl�W#.�[kR|�<���l�w�\E#ë4��hy���d�"��7ݙ+���e�O�<� 0�A�0�&��@A�-�g��:ʽ�-�<��;�g��z����5���3d��J�����t�=)Ŝrs�7�HM���EY~
�1�FޗY���.�܊��h�N���,k�Қ���hV�8��2�-�Bnwɤ�w_�7����R�}���j�1ϩ���|�Tµ�j�LfUWc�M��
^�����Ǫ�z�^�?U�¬H"(�@4�0 D
H�(Ģ�
D�><������ߟo^�x8��B9<����懸���M�`��mk�'�j���c9~��vj�����T��ka�0�ogwgeCk�"m�蘒�>�:�s>:���A�=�b���
O�j����a�v>U�"ӷȰ,�rq��C���x!7��f�pvѹ.�;!76��Й'�M�q�O�j����p~&�7���%RN.�#�H�h]��F3�	30q~w!�l3p`0B�Nʜȶ�r������fzK\�t�OI@��/��o$n@���3cL9	���F�LJl��܎om�9гX�S��%=X&m�u�`sH�ZF�=4��O�ѣ����;�q7����vq�����nD���u/<�^�4(��L(�.yn9r�Հ��49m<�`�ٽ�]#�$i���w{6/���`F6SLf &)�+�߁��k0bN���,)gO2��WO��|X�Lݖ�|yŸ�{��n��z`)����3�-�������&5���dR�V��/��
/]34Y\�g�5}���o,��[Q�(��3h���H�@�f!�Z`>�T6���{��c�����ؚ̃�&�L!+]Ja���������l�Æ6�&8���{�C1;;���A��2�ծD�e�R��q*:+�P�s�V)!��5�L�-YyRoW	[l�`R���?��	4����O�nR˕I�6p�<*æ(�nl�9�H2uu®U���Ǯy��	�U��E
bQ�BIhP��)P
TB��F�$�$g�~wϬD���͂;�f��f��R��Q�^�^����2%�^���y�׶��'�N*,c)zQW�ko��4k�e���,4���D�0�LC����\S9s�.���-��離#^��j�|�Y<Өy.�(��+���E�z-��Hr���F�P���\�O[�"&�'k�o�-�[��3/p0&EZ�c2t���=6�Ƒ����� �Ur��7�iv�O��5Nn]f�Fk�g�`z��1��S<�E�)��ė�{i휩kjԤ-{ѦSy�7��<A!]e�g�oJ{����V+�[Q�T~��`uYM|��LS��l�s ���\X��-���9���Y`�LW�HLjѡI�Q�g�u��z%�����ɧ�$>C���g�9�ò�����3۪���e�F@MNP���ħVRX&�IP�ػ|����o��[ ���q��w�uu�6��7���u�P��k��2��^'Ck�LRJ�
���qo�0\	s��50��G[׸c:��;p�f���7�P� ���"U�0��Ȣ酣S>�ʖ�����<���u/I���e*jH���;���)�%�Y��%�}l���b�0��m�/`�$Ԫ�wV�]�E&�M&�Y�%c{><M���o2����M�̈,����<�D,qݣ�w2un�*��1פG4%��&R�&e��ILS��=Ms��=_l�W?m�|=�����o0�)
I�B���B�(@�T) (
PB�i�<�q�����>7��6<x8zb�cp-�&n�;
6�P�U��r-?03*N����"��D��&�/o�ySbΝwMIĸ~��v ��k>����N0MKNж�ԡ�s�[zNT��[;�,���ܪ]q�Nj���s���75���ݰ ����C�Z��y�S��:�mv6*_ϑQ;xo�.mnC��ߜXK���K�=��i�Y��E�~��7p�Dqp,9em�%�%Fs�y1{e���G�l�*�OO�ǣA3<Ǯ��ņv2`3 �͊�C��=����������<��|چ��ݐͲ;'!�Ǥ��#���D[&w9OEFVޞ����]��A��ę�����x�g۵����Hz$@!��̓˕O	�F��͙�����=�I��s���KHC �2O~�����fY��a����l�<7��p�R���F�d����O��Jabq`����׸~KC�ԏϜ���q��ۇm���D�tOj�@i*���J����9A�f�'�cռ.� ;����,:/~�?�|n�<�-,n=i�0�iO��	�<wVv�T������/lH�6��`[L�r�ҾnHs�"��S�.���3�[(��Z�e�����oGf�ShV��q;z�0T��_^tw�;���J�SJ�d�z���1�]��U�Z���轼|�ޱ���-���'�$�iP�A�`�X�F�fAhR!F )H$�y�ox7�.�ȫ��~���%��cϾ�Jl�(2j��4�ģ8��z�o���9�W�97{�z�0R�,6D@<|�\�d2�<��'�bY'�3L�)M]��ٶ�X8��٦��j�]�������x�(�vl�&=� ��<���'�1)ծ�L���h՗鬵�H����b�7$��9.y���kg`�ٴ�`�����I��F�re�&�Lƿ��r����h�T���Eu�Ø����}�0�`�����M��N᫃n�sIx���ғ�D�������	��%���<�/Z�H�Fi������0Q��q7��8OS�N�iwgvb֝t.�i�i�j�QyC@�Q���PK�^3���v��gal��+��Yj�Q'��i�r��;k�LP���H�4d�5�����W>U�
��m�r�@Q3_8��gڶj�{���>��`t�@�d�=�n}�v��D�E�Yk����5͏=O�j"E,�x�嬠���z�yL�:b�!���	�pᥓ��V��㴓�a9�`��?���r����5{���0靫..����	��y�*���fb�qdhWx���ʦ��K����{�����W{�v��?sR}2a�/�������0�Hp�(c�'X����ni�z1	�?��>����;��"윦�&��Vc�	�ڕ����;��g���if)R���Be ���
@iD���@�T�T �|���޼z�����ǣ�3�-Ek&�n�K�w��#Ds;F�����d�d6�<��y�X���]w.���w�^e!�8�ɜS�jBw��|�xU�%�!��E�4�&u���?(��Uw�\�u��C2�3EwI�j*l��kL�O���=sͼz��"��P10��L���=�λ���օ�s�{�Uϫov+�p�4�t�Pj	�z�l���dgO3�mgr�Փ�ۊ��{�7��s���]|Ǧ2����U�j��^A=Z�,��#XΨdWwA9�������f+��[Qp�B�3!�.����*by�F��L��=�GJ��yN��T��Y�����!*��5.�Ʈ��so��"zf�t���ۇvJnc�wa��;��9D�aѽӋ���~�.l$hZ�T������Љa:��#a�&�T�r4�1�!��_���?3po��)���}I�0m�)=$Mb�vl���m�B1��:�M�*�E������"ߔ�C]c�e�݆������Ͳ :�09�iG��ٹ���=|>�/w��}?/����}9��}>^���������hqV3�^�ͮ�Jb��w<񲙠�Q��s�r�6���i�xJ;�����q]p�˹�sG",H��fT��G30gܕ�ŗ�@��5�k�%�����n��8qA�rO)���N�����#��Tz��.�1��V�q�8�*fA�R��)J�/k+fR��3��P�(�s0c�$��${0���U��[]�6���Z��P<R5&*�y�W���T��=&Asx�#X�w�����Lop=�*�U#9;3X�ZѳMްqc�W ]�i�̫2h�r��:�r��\�i�W�9ҥR��37{W�ߤC�!3�~E#E��x��
��tLK�
������o�x�v������i��;�%�>L��aX�v�m���YEt���a�,����#AT�\�ʡ�ˎ�X�1�Vٻ��wk*�S+1����U���~-m̼��y�����<B#[�UWn�G�Ѝ;���]*�ei�(�Ԝ�e�ÞɅR@sSv
�ic�6�N�٩�F���r��ut ����JҸ3�¡�+��ו�����4c����Ÿ1����BB�rV�įA�F�a�I�`L�S�r�K���f�8�8��#X��p�'�)��)��G��%��G�u�֞�t��&����Uyٶ���2���U�k����(Z+o�H�
{O�����zN�zA�\y{�cf�%Ȭ�)*�W�k�Gh�Os��[�!�\e�����O����3]�-g]H�>��$=B�S�[�x(uZ]7�e�*K'3B	/2�b�Vkp�ŽF:*5_e��۔��@�+����������Iy��eCy�m��А�׽�^Z<f,�A�Yma��Fe�������6\;��u�+j֓��|��N���*�LVxA 0�Yvs8�V8�/�IB�gC�sͬ��u�5���5�4���Nv�9J�:d\�R� ͪ�=���P�F㫲%0����0D=wQ�E�:v����](�5���]�5i#�k��P.׸i������ҵ�
�v1hC$֊��9p��vÐ���L갦W�Gc�\x7���Qs�N�z���^�⴮:��pG���W�)O��Z����Ț�]��u�P���ֻe��4^��E�St8�˽
�ɹZ:gFv�4��}�+N���u&E�+���k�� �sT���cQ��Ю�]�ϖ��`ѷ*o]�cx�f�们w>5�ʶ������S8�:��`��پ��̝`�lN6QZ��F;wDf��Ac(���W,ey��y��5�F<�����`���|t�t	�Zȭ����)����ʡu`�P:�����%ƹ�����ER�1[���4�k%�1_BPz�e��uɻ�N�b}�T�-�+u�\�O�(��h$������9s)eE¨r��U��ΐ��q�5w��/�W����B�	q���z儘J�}b����� ��� ��d���F����MQ1Q%PiܴI\ت���yj���(��涆��(  ���j��DU�QKT�DMN�UKDDRRCUPLU4QQ^�f�(Ӣ�jj")�I�`�&�*)��P�آZ
Y�"����1�����A&�53AW�˒EE4TT�SD�T��4���SEͦ�AA��"���h�x�A1�*)")u����J
�m��RQT�D�DQA%1U�TT$[x8�b)��b����YJH"��`��6tDU[&����<ڪf"#M�3)��T&�Ɣ�)���)�h"����B�g����a��M�d�;*M��t�(�w2�eNQ'QY�:U'}���&�<��3��­>�����{*�M�=o<�����}A�B�@�
Ы2�BĢ�"1 �����3x��y�ڮ�	�����")�	y/�:�
6v�
9�X�B/K�Ic�e�pM2ݰw�����Gz�K�2̇ǟ8t�,�L@3���:�ՃYB��I��6a������W\c��Ҟr�m�����L���Z�>�`��������ƇT�m�2)r�Z�M��J�53�;ګ'7�w&�T-Q��ߢ�O�u��*��ιP���?V��s��L�l�LE�p��SE�[��y¦�4�a?Mk���h�&���Ǡaz�/a��2%�=��x!0������iے��oj6����ǌ�t�t��W0��0�&Y��x�]��c^���C��3��c"�qnk����jAǑ)��F7��#2,���	E@A�v�tE�zġ0�K���u�]�m�lg���$=����ت�Ƕ����rC�h���\�	���I�|�՚������Ǫ|d���{���`���$��K窣��*ZڀԤ-{~��'�mk�uݭs��R��D�����=skb��t�ׂ`��q�8� 7����)���]T�{�R=��ɶD9��ERߓ�Um����2ң��y�ʨӵ�N�-X�{�vU�;��K}6<We�^�=nE3�(Ԅ]w-���;�S��W[����g�c�J��T�*�;u�v;�u��C��7t��i��W�oosꀟXPH� hP��A� bA
P
 �ߟ>��W$�����~�)��JBe^�hR�(�=����z�}�(Ɣ�P|���c	��l[b�=�ۺ�டhd��%1��%:���5zT.�9�Z��	����^+I��d�'Ou��n`�s!/�9�L9�v4;� �I�1�d�`n^�-��T�S�_8ʛ��Am�+���bTS�s@.�n�k�.Cwc@����E߱�C0�jQu��L�ոe���Ν������s:�!��<!h��D=�x�۞x��&n��B���*�*�|������U)i������|f��oBc@Yٚ�޽�a8�pd���k?�혒蚜`Z��X�a�`���˵;Q�wJ�2���uV��sז@�-.qÌ��:Xtz:�眅�b�z�^�;��#��U���&q��yJ�aDϺ�>%^��ֲy��.Y�^�?`��8y�뜖�YU[{���.�B��I�f8��bD)LO��S������3<���,ƌXgc&���Q�k��vjȊ���yO��mC'�ݐͳ�(�A�$@;@��?��#m8[W5Pk:�m5��>s�䣪���I�8U�:�c9�ks]1p(�賥F���tjÕi xY�:<\����Z��T��3�r���+&�\.���I�;"l Q|�f[����yO�����w�3f^3u$��Lo��!���U�_<}C���B�Q���f���5P�£4��������,3���_<6�5��h1��J��ɞ𲹺�����x��s�[�n�yc��C���v�_E��lEC��D���奐�-���=��{=�1��]o/Xn������ryt��Y�a�䮂�K�7�~9\]���U].̿��~�,�d�;�R%�=\�6�Ga�}^8�͵#�J��A���U�%�!�"��=[®��3�{�g=l�(���n�ӕ`�.��Rk�;��JlY4�&�bS����v�o@[�zW�W��&��inԭ��N낁��%��x<�[ ��U�OЂqDĲOi�3+��I�{�4NtO:I����Y/y�f�r���F����h�6��as����'���:O��Jt"U����t��u���B����X=k���O�W����5�?>�@Rd�q�7��fL�w��X����/\N��O�I���"�[%�1�s�������@A����?V���dnN윛ʬ�ŝ����]b�X�_I�O� e ��N��:њa>ހ�-��8O~����yy5����Q��s��J��Y��_���k\e�Y\�j|C���C��r����C{�o�����rX{x�P���xt����E�[z)��$���vc���4��c2��l� \do.[�ONs/j7��l[�z�J�6^�S�rٙ�e��ǽ�
PbZhUiE������Բ�r�N>��\ɉc���5��^U��2��X�:A�wh��v��2���j�r��/�A���y�d��U
�7�R)� V5����M�Z��l̓:�N4����΍]���]٢݃!a�_�x9o&vnu���u�K�v����`Jw[u����;�75G:*�r%��b5���@4!�1�3�r�"s;��-y}!��D�7s]	�ގ3ҭ�U��;�0\����b�-�i�;��x#��=�Ag�X�6�k%5�K��Z�����g;��%�׼ܑf��0�[���\�sͼg���w�C@�q͜��� �H��!&2�V��ʐ��ڌ�\ŷS����R�m�wI�b���F]�o�i�m�׶E;��ޅi�U�gwP��}���nB��!�-�{���6��0�q^�1j\���}���뷡�ik��)���CY��ǧx���`�^�>[�
7 ������'��0�	�Z�,�$B::r���/����2~u�-�b�����V ���Iq�1<�#T�&�FB�tP~�k����*KVs�v�ֶ�y5;�,�n�Ƭ��s���HW��I��j���H��:"��K�50xM7y
��c�Ϫ�Ո�n���(Bk������WA��cmn�['d���u�E�9�1��W���0j�����wbT3��gn�h��45p>�Эw���C���C婢  7����OŠ�B9|�qT(�Ymŷ��uB��D�(2�t$�S�nC��Q�Õ����7V��"���'�D�V4-X�I8���g��v=�9��u���ߨқ���˟�K����;�t�nVe�CG�a�i�I�!ˉ	����$��p�x;�0�q�Z�5����e�]}{�8.d!�'���ǰ�7\�OK�Ͳ.��i�ZF��zW�M��};f�u�fPϮ�p���a�7s�A~��hQ;)���J疣�)=XJK�ɤC<SR�ИYy�96�m�`�<;�AP�����D@M��:�M��lĝqvJ�âߌD$�<�9�[{HgZ��^��|����sۇ�p�� �� 0}ni�a1��#�k�д�8D�}l/�����������1�O=����Q�$�:��aߧ�0��f�69�6'8̓���os&h������:��0-KR�m?Mk�&�k�Է5�0��̙������V�����S[���9z0g}/H*Y����f�r�
&$���f<��.���5�-��޿ڿ��҆����~Y�wF��E��!������bSsy�ѱv�#  8N�ՙ���xg"U��4/0V��K|sJf�]�����b��"�ҝ�fhɢ��������mZFc�"���]ѕ�q�	�?R��,M��2�t�|)�;x�����ʫ���=�{�b��ߥ����!kȇ���b����#ِ�����Ty�C,�+����2&�Y���-��g��&|DYq"3%'�U�m���3 ����_h|t��e�.�]�k��%�fޏj4v��C&m�P�.�� `���IĈ��/2����ʖ��*/^rުjF��^ү3��7!j�V�	R�x�0���u[���cX�0ZD8�v���锖+���nX�P�Rɩ��,�	�Z4)=�9B�1��{�=[�O�흐/mۃO&��K��=kE�G7�mǤ&�#V��_�k;s�؄& �')),:JEo�l�=k�<'̴Y�*��C�.�٣}���pq��ʘ�v4_���5龙I���:����zm�y+�³��Q+'���֧�w7�7-V8Á0�����B�l���sԹ���&Pey�dQt���J.��j�nCR��y[����o+l]�P�9�-��6�{&\8y��3k>�M��7m�ݓS*��$��坶���Y��:zou\����֔4�N�A8�x�� 0�Qff4Jni� ���Ng���U9v	�7J��ӯN�B�.��K]�TZp�c��Y����	�p�����WВv�8q��cVU� �T�9y՝�q�O���ʷ��D�V鎲s��}�h�v*ސ�#z��[W�/�̩ʰ��_p��Rc$��N�q��׵Y:	ks�\���//,  �3ٮ/(�E��m�y�g��K|9#B�Q�/^YΩT���4�Y���@B5�O�t{kXx[Ac���U���yɉn�RkejUk
'�s��S��F�2Y��-��@`يFe�J�8'p�{g��)�;'-��ۏ�qM��*���Q�L�u��\=�{=R����ï<<�������p����{��|/~P����m��(�A}�m��a��%U�w��{�؇����;D[g���;1.��Xhl.,D���/z��L{��;���:!�����3��t8�	2퀾�H؊��"Y�!��2H��I�/�8�l�P1��f�on�r��T�fK^]+ܤ���{6���xmhg�G4���6����N1���Mnj���=o�1��^Y5궱��l��� ��������8�i�`��qO؂�4E��-�}{��^!���ǧkҫr�y�;���d���V��{�eP��\_���Ú���rs<��1�;���~�@��'K�DCέ�EF*�?B	��=�f�?���[�ɂI����Rc�����v�µd���7��_x�/	@���U�}�[���~
չՊ��{�b/iL��Uϑ�0/�fUZ3�M�K�zC���t�vWu���q�ɹ��ƅQ�IT�2m�"�b"�W6�a7�[��Dִk�%�K�g���q[o�ݽ�+~��ӄ�=D���祐�#q��휽5�܅%CzL`�u	�H�iH�Ϟ���;���~e��5G<�.g�i�q�MԒ�����@V���/c��/���MUu�_�R�gǦ�z�T�\c��k6�E�0�j���E'+�R�-�Ú��/A�<�!��E&��\�M�;O7�o�����j�;z�7/Y�j.�D7��/Dŧ匤��4����	�?KE�/�;sD�Rv78s��m����8�C�v��f��T�Q�\�H�R��w=X�8�;���@��X�[);�Nl_jvv)�&����ΨԊc�ɬk�L���L�z�s�! ���I*����}�϶ᭅAf�Qn��#��:� �^a�]��ϴ;MV�S�^5��4�]�A�551���ؼi�֐��?��C�N����(Bb���_�2}��h?[#��!�����-<��g��:ۢX$����h �z�{/��G<3�~gj������%��r٪\Tb��gs�����!���4 ���,ŧ�q'DYz�o��%��q��?��k�cWn�s*Z��|lvw�hu����J�g��e�)XF_n
�a���E^o]-�\����vQ%NM+^�_]�|�c}ß��Vh3��̡rKk�$�����}�!T��'��i�����8޽2c�w)�f�j�	u[��omo�6�vqfE���� ��WηL����&�A��u��szw�$�T�}'����A�܌�U��G��/U簇Du��������&�)!�6!0k{mO����u��4ᄃ��1j\��3��h�f	�I�<̾�&s-Kg/ �;Ń&��IO^��zaBf�s�VժO�`0�u-��vy(U����Ȣv�y܇���z;�ʋ�U����%�P��v�S�Ƀ�|��rqN���3f�yGh���g�CYu�j�Nq��I�5.�ơ����D�(2�u0���V��U�©��ɓ�i�;p^�%�y��a2O~u��$hZ�)8��a��$vE�.���a �5�c,�\�>V���]����6#r�CO�:a�wR���LU��E'���\ŗC�[�	��63�.j$4v^�Q�����A�eݚ.a��ِ%���7\�OS��<�6�摈���5��n_�ޘ�7���ܮ�U�/��5�xX:�Cw=	yO�&D�-)��rW<��I��^���!Q��__WeM�;i�ItH��G�G��*�;�+��_��Y/W��?��X67���3EOk3с�GCxV=ޓ+3�@. w���3U�X�Cs@����gN@0֒zm�cv+A���|3ף��� 	���Y!���I�W*=w�\���ά�OS׳�c+j�p�^���#�i��4��*k.�^oCP;�Bt���Ojo�e���a�.�Ƭ+�a ���W=�x���^`��� �cC�R9�!�m޺�*K��y��Vݨok�c�I�W=����ƽ�A�B5Ԯ2d�B��U�<�;G��C��	]�wQ�����6�y���Ռ9��R�m?Mk��њ	�nj��\�s�D��޼�6"-Sg]5���clb���́�,��{���\��Kj�2�u�2� ls�)��؜{��nDx���n�KۼB`�����e�P�l��#���#2,�Wt�C�Pg�iю�v�2�v�ɬ�N�e����Ou�6�
��\dfJOb�/�u�ِHxf��L����A#��
�!�l�7#Ek�"�m�P鋇T:)��'sE�UF5rw9�B�xd<��t�O.ne�&B���2�P}b�)8��oN0�\�C���3�鱬`�-4ϋ��]�l�s�;�P�v��ǐ�-�^~"Se�XPL��F�'��"�ǳծ�=[�S/c�W[J`٪`�U�w{�;0I�^N%?T�$H��;�V�!I�2�״���5����u�1�z}��g�������{���w����z�}~�W���b�/g(ɪ/*��^29��UݽL�U�C;&�(��D��D��YV�[r��4��b�|�k���m�z��zo ���l8�dD==®l҄��X�\t���^��B�47�ʛӄ�Sl�	�rg;7ncE�	�ֹ�"��־I}6��9`����Kq��s_	�ݾ������n#�i4k�1��Wv�d��0.7Y�S4�4st"�V#�j�K3�Y�u/wPZͥ7��v>يBY�@�Ny�WM:��d{�|�Tҡ�K|Ư�������3t�.)�uQ-YU�(��X��ٺk25'�	�Z����oϮNI�I$���$j��F�dm�Fn[� �j�OFw��4xo<�2�]�]���/m�l"ov'TPp,�EC� ��^���U#e,.���&��o�����$�h���W(�Vs�e4�������쾡u�\����0�������on�BKT"X�R-�t����:�#�N�w�YJSӺ�tz�'���������d����#��M%Ӿ	����Vڃe��3�	���>���t�ʹ�ޭ�*�B�%L�;/���xN#{�f���W�6�S��boq�}=���5�{٭Y[�s"�OM1�a!U��*s��h/�Q�Ȃ�";$n��[��U��WWd�z�HI�
d=�ӊꨦ+!ۛ++�嗢+u)n��Z����[e��ЩJ# <30K�v�) ;J3ek@�y̢vQ����ji�Z��wZ���F�AX�g&wN�b^*#d���u�F�����NR
��<����a��j��/d-FoM��B���Nm�`��n��c����;zr��.�25I��yh�o\��n)DK��]�*Ku�.�pt�玳Ss
�=XG��C�&ږ��y�j�6�P���ٷ�%�L�ʲ��VPl*���ӭ�nr�ME�e�عZs)�;��eviP{ׯ0I���g��3��!����,�!�mP�'O����7��V7�2�����%]��7o8�jJ��'g�Ǉ������j�]�T�z�����fm��Ș����/%H/r��5��&K��O�t걵�[]����SY�!�9���@�w8L)��jRY1	`��Y���C�?-�eP�o�{nS��#i�ř��#���WȰ$�\�ݜ6��vS�{I}��8C�O�E�������f��-3o4sv���_L�+��MY�6fe�&����]Z;�%鴨������y6nC3��g+	k2�L�K����-�{��1���;�v�u���K�g0����Z�i<��<�wY|�u��N��Kbbd���u=k��{����W<���0�Q�U��d��������z���ǑL�[E^Vm9��Re�̜��nRj�9��f���Ǹ�J����;+�c�0�N�����bRJxSq�Kwg �"�W{B�Z�@P0�LQ~lA�@  ����Ek�7��^��ѳ�j�
)���"cF��F��i*&H����������8�$QE�4�.�*X�
�(+M�0U�!EDQ4�QR�DESACQE1E4�AZMA�AEjf���"X`+ZX���"��("�"JfY�"i���b����)�������)���kDQUQ%351T$$D�QIRC�L����������)$����*�h"��(��(�����(
�&�)"����)�%���j�������"�
N�R��񨊨���f
	���9i*���X�t�����N�("��F�H�
�mZt�%�
�Z��	�i�&��ATEMq���B��ߦ���礠�F{j��5c\��N�/����\x�c�soy���VS��&�6���d	0��`���W���	�b�%:$��{�E�?i}�8���V�S�|w�Hqm	��0O���3��I�1�d�y�:Xab�x~[�"*�M���۾�,�"���k��N��/�~��;�*_��ϙ]�E������N����ҫW�����n.e�k�mx����#�&�7O�
'���Ä½�������8�R�/K"�G3��j��̚�ҍ�j��R�UB�ᡮ���I����Էs�.4��-���j�~%Q�����]�@������:�"�)i��']eqڮ=,okG/'��SL���Ml�)U�(ҹ�(%���sqۃ��?B���n�T�f�R�;5}�0m�׬BN����&���M�X.�1����ħ��A)����ac�֚N��y�3yn
�����_��ʀ>�_�8BO Cξ'��d�[��{%���/�Ӯ���J�r�'�Sdzw�2��Ez|�E�5u�vR:%�XG����DJ�/cj3],&�퐶�D���C��vB�n����D�&���o�؊��ȖxBKJ���s��������S<������Ҧ����><�\���/�;��%z��&=엔]��:�Kf�p���rw��3w_!�����+�J�A��[��˰����[�%U�j�w:{��X�52�u&-VԆ��q>LTB��}z�!UQr�*Jq�:���1�g6���7���N{�kH��L�^����*�!\�����O��ۯ,�b9�������s&�c�v��� !B�74ޟN��E6���/��C�-M�M^H���8�����36�aU��6������kFZ����8�.������M��&�d�1l�xF-��o��K!ٗS9طeVe)�ƚx�B���``�as>ղ��\��'�2O}2��<�J��;ӛڋ;%��Gc�P�r��� ��
$�6T�`���@!��'��OE�M��{gV�nh�Ӫ��0t���W@^�t��O���O3c�:Ώw�A�li�Y�
�'�Z�;�Ӻ��.�̉`몱R���JT�q#�WRO�9�NP��O0� ����}l)#Ҧ����L���w�6����L �+$�'�Sq�t����y��^��*���a(�~�r�����&ŷj�=��3:>��������xn����M�i�k�vQy��F��I���,gQ��K�wVRq]�[����w���#�v'7�����\������Lhɬk���M�W���;x֏��|�ȮR������h�{��;�r�TYuc2�v����p>J�'f�+���gR��6h�<���F���Xi�~���ZS*��Q�����l�9��r�q�ܲTΔ.\̐n+k��dܗ�6�K7��]���Bz��[�#�ֶꡖ��:TPs��>}\ߟ�;�>}��ܩf�,"�ٖ���;�9��伈v�\�T7>���D�gb4��1���u��Y�g"�O�cӽ3������;�?3ǈ�ŝ���mC �v�\�܍��j��S֩�P~C��@kNf�W����[E�b^ø�xg���xm	�V�!�̕�l���Q��ڀ6��� �7���'pЊ&h�P&Y�O=�x=��E<"]�繃����^-��̀�n��D�O��8�nsz}̳L�^���T� ܌;h�ִ�[��+	�g2l�����~z:� a��-P"�����u��X�1BAŗA�G���m�ۆ��{O#kQ���˙��n�L��sӼXP2}�y��L".;�ȫl��RB~b(���P��˝J��<vw�"�{L	m$ͳ�1���쨸sW����"K���v��u���-څs]��Vj�U7{����ۧ���ҊN��J�*�%~�x'�+G���/�hQ�y�����G%8�ى���S���%�D������N��:���j���ӌ$vE�*8�ow��k�l�DAG.z��;m���O4���7�%K��.n*Ϟ+�gj@n���5�Տ�p-��P���;X�vME���2��7/YM�&�5��|��7��D'�M����{�rR�i4ꖻ۽Y��-�ڕV�1u�t^wv�]*�*Xb�#��.F'P�{�Emq������7�����7Nܻpi��Z����:��e��Rz	@����8!����o,׮�4��y�ЄcOL!P� ��|�����NT��`��E�1�̖�;��u[���tuo6��b9��������^D9��/)���
6�aTJ�e[#��]��{�2����3�W=!�4�9��Њu��@^�G�4ps����T����2��ՃYB�bh��Q���J7}2��9qZvy�gO2�����[�������������@0�����%�>�G�v�m�����@�J�I�zb��z��W�=�~�tW��p�3%ڟ&R��%��-4�yz1S(��K1��Ú��@�~�ײa�v�5-�@���!�3�����i�V�9��Wn�.苀�Xt![��f)�����LIv�,�^��v���0��*��E�.��Z��������H(��C�|a�Q��wS0�ȯY��p=� o��a��ء�*�ww��y�n˱��݃�mᎸf����B,��̔�e� zlu`���<�+�4���lXn}vL����t�Yz�0�Ƶ�d���!]�z�9F�dO{�����2���W>[Y��M�Zd㥆��a/�������ڝ�s�����t�j��c����X���a�f-����̃$�+�>3<�� �O����:~şu����y��{����0G=%r�F��.6�5t�À�tS<`���I����y�lݑ�|��t�-���=�v:a��0�+U"V��뇡�8�nb��ؖx��ϭ�j���4��Xz��,b�P�1��=�v�����׾&BeV�
ObQ�~�u�3����d��G�Ь��Ɏ��,�xpQ��!>C�GvW�i�S�A�	Lm�JuiI`��R){���(;D\U����r���u�1��S����n8@}^����.s�bX��=�i�ۭ6�K�7��.����`{����� �6LBa�^W�Hk~�w��*�kn+��1����O=0@gT�W�ؖ4Ψe^8���ۖ�p���M��>|� ��L������|���Ӌm�М^�]*�*�z�ȴ��9bF�N�ԜK�v�}��=���kt0�JM��e,7Ǯ{z�Ha<�Bv�����N0,t��J�/^YΪ���z���o�p	ڀ�r�@*!�.�AwM7��N�ji��uRke~Ju��%��ς��N���w,�o?��秎�g���#Ön⎈�rHAn����%3����_X�+/L�,�Ӣ���T}�գV;�ȷ��X��a'�ϱ����Y�մl��gpBi�Rǽ�!����@�p$��6�aE'�gZi�QЭ����>ќ旝Q��~��=r~��ϖ���8AO"��H0͸�z�6�̪S�)���I�N�͍DCpI�PՙFkb����mˆm@ņvR`3?�D"�<��{j?V�m��E�����-ZU��8�u����� tE�jb<��N�{a��_6�5�վ����s���ke������$=x� �&]���k����K< ����Y�>�.;�z�-��E�]mE���]CZwqS4W���%T�4r���)>{�m�^Y�[��u.�����u�;��HM"22���})�")�K�L�#�ʭM�M^H�����v�am�R;����x��=���"^9t�w�88��,:�{GX�X�+��W�w)�ɔ5F[ԡ���g�44Q�z�����Cv3�oV�B��p1ᓂ%������+*A��\�� �)�Rg��P`�{��Z79�Z��4��*Mw��ơ�l������]�(L&
{BC�\�5��R�W��ϜM�u]'��%:��)�JSP;kGQ�h��\�|���_�������]�W������xc�!��7���b�G�c�:�GI7�yn��T�a�[J�;�]������A�2~� 
��ռ�#j�#Y�y�9DqpN��o�l#�w)�n>�u^:k��[x�P�@�+����n���9�1w����7�����Cw�%�t��'��$��)9Y���m�Laz0�g��ь&�12,��5�#qo,����y�	��&n܃�E��i9	�^��O�(�Ҥuy��۹IQs%�؛�=���>&X_���C��$<0�c�^����U�vvQyYYK�J;��&9�:F� �s�o���qe��U��:;l!��<�vOƽ�B�ՃR)��6Ճ�Rr˸��*�Ob�4������� g:�z]s�5R͕�n��}�������y�;k���ϴ;MJ�ɴ:��l۩���z�Qa�[�7k����Ȫ��a�>B�\CC�<	�L>��O�u+2�0.s-���j�ޮM�OPsKi'�s4笙�j�~���9��C*�U(��l=����.����3^
|�4�F�X;�6<�w�f��x�f-<`��Dv01`�c��9��0w�Õ��K����(�\���m�x�O��e7y������w���R�g���OCU����__�V�]y���"��d��縶E��W>���Ɛ1BA��?�|7���,�������;gz�i�)c���~�]�yɔ�~;f�ʜ�uh�ՙ��y��~�w&˙��u�V�Ҹ��+�WM�ĩ*JUK���v�7�/�
�E12�fbB�;N('��JC*��3V>'�DFz�Pp�t;a�[:��,g�kͩ�g9��B��ɪ���QX��+n���!	<�1�	��Lc�1��gr��v��������9e�/i�2ԍc9~���eEÚ����sb$�ʘ�v����j�̽���1����1e

zs2ǲb���#B��U&Ի'��g�1����k�_:}�z�B��v������c�����[���	�v/	�$hZ�zU$��GN0�ȶ�ZcKt�Q�̛ij�Uq�8o���o���$DzcCj]�4�t�Ou*L�p���6֞�G(R���U�uN�9�9�j�ӹ���dAƘr�L9�vGy������;*Jz�	�-�u����d�Y�b͚�C�i
�Ms�s?>m �]؆�|����F���L�m�Y:vg1��3��9u���r��(,ud��e�C4�2\>6�M�"n/��λY��tT�Q���7�mΆ����Ī,ts*Uޚ+�#vtp��֚&��4w��K�[fY�A��5���M����@�j�Q+\u��\��^��G0�z��W=�~�/���u?]��V���s*�k��u���c���_m�X������&�c�gM����5��G{�2Z�E�$)�nE_3��q鴡r�EΌU`pT�Tls]���=���_	�Q�h�o
�q�(6�ي��K��Nѕ-�e;k2_ ��G^�������dk]�]u��H��U ?�÷~�����}�o�5��u����a̖�@�~�װMz]�l���%ŗ�U���]���Ii�5��h����ۼ<��
�e��'W��f�;�[�.�L�t$�˶��f0���V��;ܝ���b�l��^]��:#ϡ�>0�l��#����i݌/�K놻��Qy�FqA��Ca��zeâmᎸf�^�t!\>����vf�5��ɦ�!��[���̞�}!᫟�:�W!
�j����c!4t�â��@c���$�n=F�L��)-��ݵ:�]
�M]br���&B���2"�Х~J��}�shlS=�Χ��כ�&&v�_^�mL��->���1N7+�-�O�Jl�!2�hФ�(��zw_���P�w�O���VM��ڳ^s�;@�b�0���!#��Cv(�����6ħV��7}���^���Mii�핞b���x�x�-��<$8��] �O�� ��>�I��]E�Hd#�R��U�y���j��<�)��J�
��qA����ր$f�!0\�5���~"�����Q���(��|�7-����D��,�$6�����f���E��.
���h���[��0��q�l�i�d�mzC�����\�!�ɾj���n)8�Y�W�f�o��������4_-}]4�������sՕ�y��x'OOm���?�TW:a~J�X�N����9jw�
[H���c�&�:�^j6�n.���-��У`-�(➗�i��(,j�Rw��]�8}���d'�o:ͼ�m�m�E���D&T�i9�jq�j ��`�F^�Gs��t;���ť��V������r�l�3xX������,_�����c��[%
q�;]���{W����j�Y"�b�ۻ��H\[ހ����Dq�EK��j�f�}��f�>0�1�����r։U\�O\k�u���.1q����Y��]p̷�,3���v�`�ؑ�z�+_�T2~�n�f۲!��%�����֏s�@������zm� �/>�l[�;��}9a���xQE�м�1V�/��Z�5�l�g�Pe>ݬ`}^��	�&��h����~ǆ{BKd"הGX3.ؗg���᪙ۘ�Qx������)f�����*�!\����ٴ�9��{7zL�"�?V��ά���p��ұ�4kH���V*���[�L+���m�26��&��Pw��|?/��������}>�O�������z�|�{����L�r��!z;��kK�H���*��lXa#X_����Ha�J��̊���	�i �t������cF�չ���[��W�T�����
X$�B�mH��ݼC����uL��m!��!�ї.$4G:[�����c���w���!dwu�v���嫪w��9���#yFmQj�Ȟ]�W�;"�ӚU�AҪ]�6��l������|n$�.U�ڳ��p,qv�j#\Y¥���/�(�}�wb�%�#�������4����.�V|�dm��y�:�(�kV�c2�4�l��tu�.���I_a�P-��շ�{8f�H-,���E'2���<�b�����pf���B(������77�In��M�9;�4�6r�)ZgC�_wv�N��[Z6�J�/�1��k5�fm��4h$�v�SC��y{��aq-�W�gT:�s%�K�}j��b�Wnj`�U�eK�e�=�řǄ��)�mY�f��#�K�;��:��N��ɼ����<�x��Z"�Һk7�ae!����unJ�S����\W��
b��V3E���B*)˼Ӛ���u��VX�-���;�y�޺��P�E3��,(�R<^S�Z�1[��SU�X7D�ۤK6v����i��X=��
�Wc.U��xr��v���{̋�v�'k�eG�l�xj�﯅����J��.��p�;9�b�$qS��e�ݣħC�x�"X��2F�9�2�;�o�)�Ճc���Wz��b�2	���d�U^/�p�%S�ko'-+�Z���E)���?�������W���Ӻ��X�<��Y�~�Ŧ�Of�]���QU�H�&��'l���3Z(q��Bt��v+�%:(����{�x�	�(F���Xxgr���w�_�B����5} {�h�����!�u��b)�8m�\�I"��N�e�Ĥ�kj\�wg�w:���0cɤ�oҷ���^̘m�X�*mh/x��7u�8��Z1�u��P���%���S O+���Չ�g!��\	�C_V���";u��<����\˩�ymuMڦ��XM�j�*g^�2��3�3UV�4T�cӑ�FG�g�|����q��VM<��0�/��ȳZ�m*�ݧ�Ia0bI�� ]xk.��f�gej�8� �[it�E�G+O��D{i�^����+,��r����Y�e��(d�ybeaΜ0�q�\wGP�X��z���.�x1����*��zd�R�l���N�{/{���ޛl>���5ɮ�ކ�l99՗t]R�U��*đQ*�/��f�]*2�:g�&��	ڎ��{T�=���y��w���6tT����]PfeN��K,w9^m$����c	�2�p�qkw1Ɣ�4։�U��a'���ad�d��V*�C��N]uk3�ڛ��%����X#VP�ڽt�1aJ�>���C
�a���g��\�x۞.{p�|y�PS�*�Zv�D3ST�	AJ�E�%v�)�*&�)f��b�������
i�
H���j���(�����i
H�����u��R����)h��"�)(*�����(*���*f*�������I���$Z����AVƚ)b���ii������V�TQIED�%S��(��9�LM-RD�D�LM!��K��Q0�͡(��K6ƍj���ʇ�P�R�r�%��%�bhcr3�̴h
JkM[�����"77 Ӫ	����D�r1p��4��l�ơ9b�P<+����Y�wﳸ�yF�$O])��K�X<�gT����i�o��C��{���P��Y�gTY���\�S��CS�{$�2-��߷������K��������	U��دH�"Se�eL�n��u�r��+3����Fq��ǡoV���'Kw��j�W�u ��K�&V]����ѽ���8W�,K�Fs�� ��5�aom�����{w� ���)���Ba0Y�3���"�U�7l�I��T��p�] �%:O�bUB.�~�V���� 䖧ȸs^����ק����y+.,+��]��m��s�n@L � Z�`��q=�i'�1I��7H�Am��F'����zػb���A�!��J͍��\�Wv(�8�A������w2dnO5��a�[���'�C)�{Rm�xwiۘgl����wKjߖ���T�n�}{^pq��i�@����6�i��N���)d�e/o3]tB�+ob�緍c�ݬ�Aa,���g`F��7s�d}명OB��Lhɬk�ї�,�<C�]���F�4��ںU�u�ߕ}#'�Y n�B}G�*��|]'mt^�T7>��lQ�nZ�w4�XU�[v���D��I�Y[������A~�����#a�>��r1l�����ȶ0�gܫq��_sD9�ykF��dF�c9O
�[Mq�_��N!<�����oF�V�-���=�]�XR�Ӳ�J�gs�y����M*��� �I�c�EJ�$Öe�{��;s��iN��Iu�9�5�ʬ`�y��'N�]�N�*�}�',�1���-t��n~�H:�?��$��0�D�	���1�P/a�@ΉgsJ��>��gSvF�Z�ˇE��&9��#[����s�;��P&h�Q2�Zx�w�,��*,��vF���y��'�����4�K�!��Mb&
u��Nsw���i�	��n*m�h2,���4��>e��R~�5���g^E�n�?`���Ƚ�Us����cN(H?��kuU��ն긻8GDnw�!��&�Cb��f�2��5�'��x��2pBO>��zap	�͂�.֨�{rL�vn��\ˌ�Z��q('�P%����>x����#(��^,��� �\؉.2���{�x��ɦ��Oon��e�S&|s���2�\w=7�"J�I�2�h���:�g����ܳdt�u_j���
���3j��ײ�òsk�&I�9�N��0e����]���_r3Ӳ}};Z�{�`�E!��萣a�<�2��.�}��#��&@��')2*���ԭ�w����SD��u��g�w�xa>܁ DcO��O���|�,���4�������=��5�m����I��edh�۷7���� ʝ*B3D\0������ؗq��P���ɗ��b4��� D��4a��st�ݴ߉�غ:ܬ\���ٶ�|x]���ۨ�V1t��^��&]Ǘ}Z�'����΄��woX"�.�}+�q�����l�UeYb���nB����J�s��|k����G)��ɠn���~k�t0lkA��r�ץ�?P�4(Σ"6n���ӛ�[z���)tb�˔��),kܶ���<;�@܇�`��a��~�L�^aT7�#�}W{h�Tj�~^��֢V���*�
:y�*�a���Z�=�x�8!�K��'��W�(f݇Y�g��?z����L۽����Z���W:NK�xݒ���B-�},�������-lj&{1�W܃���@u�[R�����e�j�>MW�9��7�`��]�+�Է2�MA{kX8��o���>�!6���t�wA8}�c�m�Xʖd�X�n�w(�%�l�̢��ũ�xW�q�y3o�Bf]����@�t�a�
�26�|Z/��S]����-�>��ȗ눣��xvb�x���� ��˱��˞)�lg�e��c2Ry2�~aB��������ʀ�˭�"�1����r9�W!
�k�o��:l�T\:�{���x�S�9I�j��^�;g{kB����|c���-�]�B׼0�*�t)%'?{zq���C��z=�d��id�ǃG�`�R�&gt����|� #f.�<�U�ӫ����f�psV��J���u=���L�M����ڣ��Y�ֹҵ^�>���%����u��8yՃ�]��;i��FpS3��{ŷ]�P"R�O��`�Ĩ����nRu-�fW��rN�N?ɟ��sN���<��O;b�d�NԷ5?)�ɐ�U�B���P�.& �&����fQ�t5��@��v�6-����S!�>!�݊y��	Lm�Ju�,�'�����䴋���҃��d~�m�6��y.��C�h.�|�'�_7�;z�#�ϳ����ߜN{�l�y^���3�PIR`���2k�ϭ��A�l�"�R�7DnL�*�`�R��ݾ�~b'��FVE'L-�]ye�i�n�4��6�8zd�c]���E��u�ַ2��pXܽ0j�"V��(qTqWKׁȴ�֔45Jw�L!��`>��R��ˈ��a����`�� ��Ö9�4\�58��i��3F^��;�U�t;����".���Ļ���]w��\>yn�q!0�z9�����j�[+R�Q=+����N�����REgw�[֪_��(d��6�1lH��t�#��;k��vm��nt�+2�1�I(��y�z��W�gOK�T�u��1�c�,3��g���<��}�d�y��g����	�s4퓭�����v-."��Hmܯ����#���N|Α%^]��w�{JÐvA^��)�A܋=b��]�Ji�N�Pt�A���y��%2��B�.a�{g�N����o<Q9v���;�_UUU���t����?m�۳������	�t��`D[��s�]�����ݵA�$�h�͍�K�'7�{{y]�j0�$�c�6��u���D$q4���g�R�������)�v]p�����寽���>2֘|d^�E���$cv�f����׊�P�%�=�RwyҨ�T�S����c������,���->#���FS���O>�E6jJ�����H2�S�o_[�2�
%�Un�3�c;�^�/C�����zâ�o��X�(ןw	����]���s�Gm��:�I�a^=�^��x/m��)�-E�s�/C��x$�&�{:�'�%3���m�~�	�%�t�I�de*Mn�om�L��Sۼ��ٞ�4]�V8�b�>1zz�;�ݻ�Xj����VI�?D�I�L���ʒT���y��.WG��ac����ء2���=�ۣ�7G�0�6�0��f �'��i'��'+t�T�a�D���f=v�G5��C���yЎm��ۃry�=��ip�S߉�NVR	v��zz���C��i�[��~̒v��)�G�jү�;���5�p ̣̩�1��]�ny�}���A��J��()c�ػx=0t�����)eG��g�`+�A���t�K�kM�[�VY��"����2px�{Ź2&9�����6Knv�|6�%��G����+kH�0��̵�mt�u��� ��ۑQ�����Tl�u�*9�9
n�^ޅ�L��s��$*Հ�_�Us�G��D~=��IS��R)�چy�=��[�/��?G�������C?{߭����&�LCs�����R�T+*(&���Ӭ�݈��V����\�JaşYc���}'�J>����P5�x�o�:��sm"j�hZ������j���4��N	Nf�P$@;D�sP�c�-A��#f&y�Yfwp�},�ƟD�W�z|ފw�k�7�ԙU*S����j�U��^��̠f�)��>�8���p(����d?v���� �s�����.l4�Mgx�X�7a�[�_?4B��c��+�M��X(Y���[���a�N�y�e�W{vxw^���Y�̕B��z͜eC [:~`%ެ#$�ُ,%˛Њi�5���&��:z�u�I���ב��at/��`&T�r�om�ʋ�3l ;G�#���ަ\���;�M��j�МV�^س�F+|oVڮ3�}R�N�s_!��b�0=�g�m�B�W-gQ�䕞����K���M�y�}��3���ق���T����S�Y���kf���1��T�S5"��뷋�U\�u��?Qq�	�{6*���g
�3���瘞��7�,[�y���zbq��-��y��e�d�'X��DJ���jQp�o�]�R��Sk�篻3�r��0�K���/e��d&���L�ߜħI�I.:	���#���u���&Tґ�P_��<�p����r���9�`�d��;L�H>�T�c	��%��Q[��&lLFQ��ӓ����4��/A�-��@�c0g�j�!?W�� ���,���3\+�%�h�6�CX�XN��^��zΊc�G8�CiG���ߙ��8{h���a��K�~tu>�4��]֎��Bq{:�������r�'�	Ic\�����vm�p�85�?�)ui��߀
8�o���z�j�Cj)?X5�,�1'\]�U:9�+�`Z���sۇ��q�n�z��<Ϣ�q�46�0}kg	�vuHn`�]��+Q+\u��\���[_����F�\F��J��d2����Ir] ��`��p�p�3>x��i��\��f\zq�1�drO�Z�L3N�O�GqY�6Uu�Ml���]~zm���A��"]�Z!0�=���\�ږe��wKo��ǶX��|}�i��cm3ºݔ�����Z� ��s�����Ž���n<ɱ.U���	)f襄��{��<c�V
k������}Ո��;�&��u��:6ԧ��Z>�l��'\�+$�;����4�:�7*m�f6��CGDu��:WG.$�iR?�����ͺ�	�v�tE��:���k˼ ��:�������q��S�v�p�uM1�gs��a��
���	`�4�2� �e]ok`38�`L�"˃,k�{my^@v~�t�k�e���,��f�Y?�1�/�\�(F��.6�5{�.s�=e�����تj��3s�����A��b�k^���ʖ��o_�ȏn,�k�:����t;WDT��[a�os ���[P�x!64��i�Y�H��C�s��t���%6Y2*��B��F^aV�k����Gz�2�}ځ]Ӻ��V��Ol� ��5@�����{��2%1z�L���CSG5�f���Zә�N�7��)���S��IP��l�=}Ǆ���7�����������L�ŷ��Y�ٵj��s�r��2S�e�:��T���_8���OZ����>�L;��$�a��q��wgv���8ܘu�]7��R��n�eKLC�|���6h���o�va����93C #D&���4(�iC��,U��E��%�{T�~jN%����������K��<�=�X�P�o(�I֪���5G�Y<fu1�op����i��˕�f�x
Ѹ�cw��lPw,X�SFU��ky��:�9���%��h��(c9�i_#/��m���&��L���a�5t�}G�b���G�ބ-�{N��Ӻ_���9=�ؾ�A���0t��C����-�1:v���˫}�l7"��{�q��rng��}ˢ%��î0@B5����Z��SM��U�[�
i��zW<;�6p]ʋ���8�����~�Cn9��f���ӅJ4�����|]"8�p�Ϙ�O#�UM"���Ǉ�t�n���-��>�3'\���>�,ƅņv%�7��h�^a�_���0��g0�\:so��ri~C��e#ݒ���^=%� �/>�lZ��;xw����7�a�d�buY�ಜ!^4��Tf�D�bwk;w9!�%�H"��N����u�̢K�Z{�N�r�u�=[Z����OZ��h,� $��~m{�������W�Iw3^�.�����Y����P����pc����d?\�ύ{rfڵG�vm��Peʖ�m���#�7�/��=�?*�}$\/�z��޼�0m����=a�w��uʬ`���y	a�qq�G�,#�r�V�=�g�9k��4������V�^��;�A@�K��H{�x���ۚ��&D�}�ߞ�nL��Ƃ/;�ًY C��ۇk4ukĻ7��Hr.ֻ��i����ouMc���|2�w�����V��Y���҅4�Ws�ݧ�z%�\�A,(��6v·:���f���O��Ρf�s�P}ia36���fɩ�.Y��Mց
��]���Eд��Y*��wIv��`�0Y*�5y�Z�����Nl���Ө۳R�,6BƐGd}��Jt�ħN�Će�%I���&ry�ϑp�% �;�f�7�ٷ]�s��+C��ʆ�74�W�v�2��f�8��F��F���+<�"��Xs<gDp�ġ��5i����S�������E�y�A�nD&�!�w/��-���E���׉�O����\���!�W[s�ռ�k���!R3L$��,"�`�Y؎q~��Z��W���õW5卧��	B�-v�a��Ӽ��w��r_uיc8��wm|gaA�����a�?T+�p��g�>W��l�-��m�kn�͵wA/̖�6�a\���l�l[�6�j ��$�����H�7�j��\�+�o&�t6����K��L:�Ʋװ	��u��i�����]M��
/����|����4��Gtl�M�>�M��6����j��Gi'1�a��Iy��_�9i)��ߦ����rI��]��;ʼ#;]3Ûs�ڑ���Pny�4&�L�v�L����W���������ޏw����y��====�����Uv�B*ٹ�ϲu6�b�lu���O'������0x�dȝ0wZ3jhwlB�*�Z��Iov�J-qE:H^�,]���yщ���'t
\tjN}���a�%m�b[�Z����.���1��e��Ǝ�醫'vgj��Q��19�F*��v��RK|��϶��q)CU��֍������M�|"�8�r+Q�xҲ�ͫT�|��C/x������V��TE�W+��JWݒ�4^}]��;Okh�l����b�ʄ�3d%hW���NgC �h����}�kY;5鄣B�'=5�s�%ۙQ�.�*p�����*$w�[N���ͽ����e*}��F�\������	���
�1���L�ʓ����Z&���&����B��V;�Tei�mRy�s�'��ݹAq݂^u���z�6��,��Ἆ�f��5cn�[Y':n=�-3o����f^*G��dӛ���}e�� �oo@H�b���kH\7�{��B��e⋮��l*���b�fT؎ٹ@��E/��Q���C����m�u�g��0��w�f��^��^�]��Y���3��jHh���'��2Sf�k�C�Ż��{!ye�7Am̱:�
#x�ǋ.l|/H����a�$.]�]��ڸ/h�0���^��A�%L{@E�M��$m�P�p;Y�mp�tU�R��yN:a���X�_J�T��*���c�Xr�6���
Y.̔%�#@��vY�T�6Y��֯f�pvj��A��j�͕�(N�3*u�:�>�e��>E��,��'PL嫻E��Ep�ot�m��A��Uy��H�˹׶5� Z�L՛�z��W1�9�7�-Sg��eww��J���5K��0��[���[��E�5LZ��+UQ���qZ:�M:.�s]*<�ɇ��-aCm7Z]kn�V]m^Ye�<8�Z���-�Ks�VPo]3��Ц�r�`=& �uQ�3�0�E����4��|�j]18c�8�'h��s�[1k"]g6��Km��
�g!i��%�Ν��.�N�����sGvY�����vP�v�u!վ�aAO���s�f�3P�Q���eX����taG�MA}�T�X�m��]�:�$��f�5&-V�k�m2E���S8��j�S�|E��5]^A�%zM������[{�L+st5�k��[�X�(��T�P�:�wx;�js˥Q�fhlR�z���U%V�B�x��&����xuo�zx'R�	��3��GgR6�
�ё��WV�9{iUw����w_w�F`o1�eP�Dۛ��{���,� ��̘w�f�!hB6E�|�F/�	�{��3���ͬSj�c�m�/k&�oEm�z��e��
>*#r�^^�ϸ��̹-�4�v���V.�K���:&q�ǋ�M���-L[x�>�d��R�KXg�P$I�D��
'���LH�K� �ma'A���<ǽ�׀�X1m��'6t�F"*(����Ѷ����A��X�Tb�.��������Eh���[!����SB��JMEMPE�t��I�hִ�AT�Z]�εAT:(t�T�M:WAF�R��43P;4kT4TT)����*64�EUD��N�|l���((�����Jh����)���)�EͧUT:N�U�V�R�E:Ѡ�PM�i�5F���iMӶh�4̴��SF�Z��ѠҴ��!9��jM&�ZlR���4�$�4�b �"h�2P�*���nf�J*��l�:tIF��
  >�<��:@�Wo׽���H�rjS�7�x����y�<�V�$��vjmn�{Q�	g��=��V�g`�3�2���cEV�
�PIP �P#��2�rk��Eq��k%=[�^m��"]��8��o����=S���	.+۹2��i<�9M��a����y�_)�dL�hj�v�o�i�m��k�J���7��
TmX��n/>i�r3l<M��NR+�f9k!�����!�P�jFq��gP���=;��`d��u3�47_i��uv���h�=�^�RX������^Q��a�-Ey����k?g����r��S���c#����-HRD�^c`TQv���,���ѯЃ+{�1I��4)X�I�2�n�7l��`�>�\͌�m�������
�]	��P�/e���Jn`�2�(�1I��F���?>d�,��۵�u�չ�i�]=ZŴeӍ�cL:A���S�.�s�u*L�<�3-�rv��؛��~B�Ox�t�磤�6 ��_�<[�	܁AƑ3'�/���R���qStVv�got�����T�zJ)�t���1���yٹ�_�=���¤�|�n�Oo6�?ךcjD��\��hQ[)����,�9r�Մ���N:��~(�j:]89{|�:��럟��ͯ�RdQ�w�+]J����X�"�F����vBW�����fǫл�-��2�sd��w���^�CD]���.V�Ï|	�Z�������
�Y�n�<po*��Ӯ�=�D����R��]}�uw,B�S����+��.H'k�����oG�hwĿ⨤��5�,ߌI�~%QaK:y�XWZ�A{��g�=�|��W[k�."b��;7}�P`�p}l�0t�� (�5��^�4-Z�Z���W=����Q����j�����aً�n�B�V��GC��G����i��涥�mv�a�@�T��~��rc�}�|��ё����U-��Z}�3�2%��!0���~��,�:��,�S�98m��ڸ����uf+`�f']�ԍ3rb��D[�}5���@����S�������M��WgW?a�8��a��^;�AQ��O#.�C�,�D����w����pTk?_'|�9-�u8~�<�/V��n�4�B!��/@����W~�x;[g��b?�f�;
]5�̸�a����p��0:�sI�_{g*Z۸�R���T�Z��5,�{�eS�ߝ��fR��7���~�{�G66���s��d�f�_���L���޼���&C5������\	�P�ݑ�V�����-�/�0;+�7b�e�|�L�������3�����P�q���ăg�5����XO98Yǹ�mZY�z˅��`}ӕ�V��mfq������ީRq��X�\��YM;s�m�`١Z�G��Q]fM�![��`�����V{S&�M���L̆��19�-���q�c����K߸����O�v�{_q�=[�	-�:A�g�iiG\k+���f��5�е�fRt�$�7E2��&��(��O^�֏H0͗�h���TB��sw:�΄�����ҨvQ��N��wL�E��tS*Zj���-N��gU'�%�n�Y��a;".���ʽ0t��6,�҇@⮗8����Q��S�4��eϐ�,�B���ם9������^`�����v�JtMN0-GNл%Q��,��T�:G1~���F��n{yTӸkG�4w��-���む~G�mM6���L5�
Uk���6�آ���摽ʩ��Ri�S�9��l����B��ur���.��4��f��3>U��s}�X��V7!�k�ݨq=oL�uɈ���,ƌXgc&3�04B.�w[Y��[�ǻ�A��\^��T1sY��Gd��`�zK�"�&+�C�α�z%�2o%®X��Kw�6��p~�"T�{ڌ���c;����$=D3	�i�A}��G�Ђ��L��{���fEg;)4*���y�MW�.#
��%�]_��h�7�X��T�׌C��3D{�����}ٻ�{W�E���CN��56����n���$cU<�v�r��f���J`��Q��%���"Tb��"�GJ[hU04��v��F�^������	2g����<ڼb5��2H��I�^���ui��L�W�X]'|����5*��+v�OU��]îɽzO6����@X�ii!Bi���31���ɛmIK6DU�V�ɡq�D��A�x���	9A�b��=���.�aŵ�Eޟ���J�aE�+B��f>��Fk	�������-)A�ZxO�#8=�Ac�yO~�fq�@�/r��׶=&w�W�{{�P�\`r��5���'�2.�H�2�%*^��ơ�l�魼�8VdE��������ݝ�%�vn�fAa�m�vJ��	�{�JuiH�T���\vMy��s�.��vE��z����x
���3X�V�0Y�=;�JO��&*ۤR�ba�E���Jv���ɿ���+G�՟G��a �#��"mLpm��^��OdR�	W3�.o'�ΈΣ��ʩ�n�̈́���L&9�H���7��PQ�0�9ó�����-�+Tɗut�����J����	��O��c8�������!��y�M����6s�[E�Ƥ�4i�%]�<�G��H�=]�a�p�{��_3Ye��h�SZt��{w{��^Ö�m�/���5%cֱR�r��F`wī+n°��v��j�u��ld��2�-6Y�]�eL9�LÌ�a�l��\6OwGwA\2�'��ݣ~xB��`(�'P�Ť���mU]n���1���s�k�6r�v`Kr�J�k�;�':9=s�5R͕�n�����-u�nʿFF����~����;k������T-'�ø�e�ĸ�uz8�i����B�XAf��T���ioiګ�Lx���	�;&���d��dw vP	���4����͂	��`�inl�Q��^�s�w;<�!3��V�>ʐ��Π���8hP&$����=�]��OS}݌�Ř�Όw���9�Nȗt;H��i0��1m��ty�BC���u��m�חi���v�� ��˱mjO��x5���	�"�@{�d]�U�B֚E�fBU|zߵx���E�"W���-E\��䌆�^Ͳ��l�瞝�X0,�P�ܴڻ��1l�m`Z]C���"��	ȫja'ּ0�{N!�]6�A��.b�Ϸ&=��12;�&N�W#]Y�=N��fDT�:���چ)�-^���@?A��tȋF�+�E�5P٦l�ʙGV��fT+e�Ml��kz�/�{�@'l�G�MͯЙ'�1)����s��o1_��=���ٺ�i���璍��_)�"~ݟA��@@�ń���2}���wj�~�C����`��/�K�Dw�ݗ�P�.H*ot�̨n���u2NƲ��G��,2�e���	��d�WS#��,��'����`��U�5��w�j��E�H8�rNܻpi��H6�+:2�Ըj-������mi�b��E'��4)�/�����	�!#z��_�t�"�[9R�`uWF�yx������]P��)9/,�����M����R�����-��8Z�&nN����}t��p�r!��	t�!b�H��%s��I�%�jT�'��ݛq��2��0������l�m;�Mh����������h��.�TXPY�̩T���	��"Y.��d�����R���Xd�^�,s��R5��B�xX�I�\��@{c)�*�kNھ��s�զF�yS}�u����y�
#��k�T���fYCr��c�H ��	���:Z�Zڸ��7�S��q�nj��^�^�9�!����C�e�d�2Ow�N�j�]zh�l��G)�3j�Z¼�Iv�L�z̃���l��]�Ca{[9i�)ʓ��w������7%�Ws���Ѭ� ���0i�e�N���x����@�����>S�Y�|wƪ~�-��A�,`�P�G9���0Q�5Eծ:���X��4ɧu��p��ո�׳�V�g�=�Ċ�11��W[G1�d�3+Tyss�Is�Ӯ�ƉYxW8'Ew
SO_�q�bf�jSc�b��e�]��3(hK�LHs�k���o���d��d��_�B8�"�s�U�[���cf9!᫜��i��/\m�d:�!չV�O�����/�'a�|a�>��%Ĉ��/b��{r���R���a�P���I珞!�n5Ξ�S���{X:�x)�ڈ���
��V.�?�iq?<	\�K	�����8�1��mTj��x�$G!-k��4+��$��sSO�x���ϟH��{Ȁ�	�	weL_^m�wo<�qּ݀ω�$�FUO�s��&��C���|�{��M�fY�ȢJ'���<cȚ\�1���L�%�eO����u���a1p�ޑ[f�7so0h����Ԑ�i� �猍&�z��d^��V$���..�&wO׮�ژHd7{v�8�����:�$���ͺk�/q�n�wm�Jo�3�W���c"
�l�uյ@�`mM��F��r���ӰFi�6�A�/P���8[�6gUt�G���+G����wGߕ7��8^�-i^�m�'
�����hbΥ�~5����@��ȏdBk��ǲ�bK�L��g�^*�����ڤ/ucpJ���o~6��4��أyu;CF3Py��۾�qvb��rȡ���=w��r���������_vE36�t�a�p޿�t�$MMNL����do�>�8ߜj8�;6���H�GEwT�������q��6Z�������ӄ�M�W�֤n�Yg��0��T��3@wє|�of��|_��>�3�sw��I��0f��6CĻ�J����{�:�a�)G���xX�'�ѱ<;;�{�
4�3C)w9_-zwE�q���ا��gAȮ�?��7�o�=��F���"�/�7�XU�o^�b++g��}��,t �5R1��ٮ�DCP����W�;�jDy
�>&��Gsmg�-��j��0�W[�s�K�e]�g\n����0a"����R�$�����5ĸ��2
�5�܈���xUVfm�ʱ�_�$t�����@��I(\#2��Э�Ɩ�k�!o�|�Q�� h/�EO�WH�n;H�s��P	%@/o��������Z�Y5>�gN��U�5ƻpoq���wP�#�a]Gd��F@M��$]��k$���ٜ>�J��Z�o���+�C0j������u���X��@��ǃLUdTV���G��Ng-M���)'�ѽ;�#5U
/�.���d�9����s��
d�2C�!�P'v�>wJJ�ܸ��wIj5[��b��oU��J�8Fc� �w���W�d�M����ٳ�㯻�kdޮ�Γ���hv�{��y���[r7�D-���oVϽ�V�q=yض_�,��˛pvk݉)�{�{V4�2��hf��=�&�f�ƫ�ѭ��Rjd�Ҩ�0r��.f��T2F��4;��+��c7*��@�9û���n<#����T��]E�m{���������c�uS�˧���=z}�t����[��=�:Sx�}�^$�Z�A��Wä��>{���� �sE~3*�bU���u�Iw�6j<��_�����q���Nf���pGH�#�h:(�S�g@�`����4�2��vu����4{�����@D�fS��O4[j�-��^�ޟ?��V1t�E[���1h�����y�d����wV?Moa&���w4��]�k�{�'��\ya�G�oN��Ko��Ws6�ۺ�ʪͯ�9c%�;��[9<ڦUa��ST'9�8cȳ;
0�v���Swة�[sfv��1����x�ro޾���؉�~���H����J��VR�V�GKf��h˗��]���]n��1w*����Ǜ�I��|A�QR�$q��C�=��8o^�fi��u�
���d#� �Ϡ���"�����tL{����5�߈�Ǳ��:N�|��fO�{�~��UoL�!�PE���[�6���%o|��Z�xn����6Hm�y���5^|�;��{2�pB�Q��׏�X�!�/Z��|�"�q7�)%a�T�"d��j�9���A�S4�C��n���������f��_)4�9�KJ�~mKW�S�M�AX��O�ö�Oj.���f=����h8����W�bU~�Gx�%IwH�YHPÄ;��`�v|�{[}ܳb�Y�����魙*��9�9ܹPY�r�U����7!	d��n��ї*���r`�0�_��=���iPP����z����|�����>�_N}>�O�����|�_/��>>�ӆ��Ƕ�c��E�����dU�����5�S��J��SE.�AY��'�f��+&�%��<b��KkH�n��X���h���Uv�m��c3�= N�ǌ{�ֳ�
��;�O^�x��C���[,p3��c��g�U��	Ύ�:�����nV:���љEUҨz��xsΓ�k��[��G��6�/$�Eɛ49�J��A|�d�ߎV%�כ!����vgFP�4�m��46>H\ӃJl;����9��^Mf�R����"��oY�Lu���=�5�n�f䱧�yx�q�|�p�T�v��,�Awi��
y�35�R��%�����֟�����b[è�~P����в�����-,w-��q4D�Of��u���`�w^�[�qr�٬��N�pE�|��W��E�lϮ���ͥS��R��=�,���6��gr�&�$u-��ю$/�gw=��z,��x�O��0�v��t��wtv�8$�;�J>6N.W�_���\U�u�ae^B��(j������F��)Ļ��d[�����q�d����,
�p�+	2�8��c/yQz���s�����(<�E�^p�+M���j$�01.��{�b&�h�R�`V���)lO=�+KË �3���C���ע�DT���m,&w"��Z�D��c�[�"��h��38�r�<�A�ܼ�Ҟ�v�a[3%�w:��
��x-�&�Q��j1��e�v�5����2�U��9ME��]�<�o!���%�K�����:ڮ �(B�Ӱ�!2M"�C$^��&��;���\[Y��:��x�]A ��1j��=�P���Sw�.#�LY�R���Qt�,���K�p{R��Y�&+#G\��B�0�H��=p�4�'^�E��H��O-�����ԝ+a��`���R�N-R��R�g��C1�Bq���tM���;��:n7�"�d�uI����C:�<��X�n݅[�. sv$�)�Ov\�Qo B���Gg���tP��'/zT"�wDn����(� ��w��\J��ML���TA5 �r��u�����h�#�Igm�YY�`XlTkU��k`�]0���N��yh�Z*�C���9ڥ�ͭǚ��#

alr�̃V��0�[���cH�Tc�I�����M
=ԃ����}a�P:U�ZDՊ�H�ִV��d�$�!܍��P>F���ѻy����(K\*�99�s���Zq��w;�n��Vԙ�W:}$�<�v�i��]��Ιu��D��ˮ�ְ�9��ù���W��ڂݝ.��y�ۦ)���z�9�Bs�q�'��:ІN�؆Ĕ=:����Z�vi�ڭ���e;���et&�A�)�<�7���R��MA1��L�Į�jH/U��.s�u��0=YN�����˘7V��J�O���������۶���e\{�2��n7�Qt�XkDCٰ �u�ysq���Ȗ�*�?:`
�0&��Pfi4�U�Q:����AZ�P;X)�åh"�N����M&��QT��Yi����M�F��6ukF����Tm��AT$lbq4ն�E��Q�m^9�PhѴm4+AA�lh"��h�DF�M:�����:��@j*&��TM�Uj�T:
i��`�X�X��M�Eh�ޱ�y�X�I6�E����F�4[�&�Q��EU��S�����A�m��URSIl�6]Q���h�h�EE&�(b�+l�:4k@�դ�<���Fv45���ibM:�m����$ml��D�h�N�RPh�j�m�m��l֝Dō��8֦&�����5$�6������痎z�|uԕ�f�!�7V�*T��i˰�L��L��a��H`�w���':��j̳|��u8�,�]�5G-���k�H��St�m��7��1@�
����&7[I7�/Yz�nά��m�'�'�6�ڰ�d�>`<e��5�U��jhzؘ�[}�����xtx��^&H�O�����6�z�@�b�b`��P��W.HxҨ�J�p���yw�O�\KG�
��/�
e�yAɚ���f���N�F�f���(�Тʮ��7ۑ��yǤTD�<�/��I���2;U������Q-���CTx��=ܚ%���܌��J�((e�2�[b��F�d��oMfe1��\ә�g"���?G	�,I��ݹ�Bi�*���M�n�m���)���S�5��܊�sV�BɹrD��h/M����niY�=t�r!E��z�	�UO�s�P"Xg�e��I&�y�	������u�P�!�W�,v>&u+c	W��3�IT�����>�~#	w���kXԁ�*O9խd��}�=�o���ł.�t�C|w��Z2�j�V�R�gN����Er��G��2��8�Z7٪��bu��I�oUI[��}�fZKaU��v���ݎ�,�=�T�؍]������_hm�r���Y.��ȬnqM�����+$o������<����V�O����#"�7��1f��=ݓe�g�P!�p9"5l�t�8�<mlwI�[��F��d����y������a]'�$?��*�l�v��eVmFJ��pՕ}[���{���'wM��Lq�������Z"ðͬ�w���ո����cmPE.H��$tȹ�O��o��8�E芌�fr�sV�wo^���%��U�g�Wr��LO���:C\o4��B�<�n�Ŏ���>Ѷ���Hܛ��=���3����.$��;�늶�f{��Mxw��vMf� c�U�
��f���V���^��$H8�ci��ڼ]��:����jLSﶽ��`9�?L�`FOxZ������VW��P���oD�Z�U�S��g��A8j���M������{���[��Ւ�d�ɢ�1h!�.J�y��9���7aҮ&8���:z�[�X�ڌ��Y��(�]c3%�V��KnGj�j:�"��j:�zn)�Ng+0�wG{Q�4�:���v��7�!x�b��h����<�y��J��B�|(��F��jv�{�f ��[�|$Q#<hj�#�9����P5A;[d)��k7���$���Qq�4����AM(3�z��o�z����-�Z��O/������Ϡ��j�!�h�
&'���@����F;���vt���ǎ��Ku���;��XJ��"a�%�#^����%R�gQM�oMS��d���-;}s�>_\�X���HS�Q85N�?t$�p�ܫ��ή%�_\?I�-����wr��8d6c��]9dᱷDX6����׹4�6wOS�>��(y*\�2ص͓�*Gr���PG��xFWHT��>�����������O3��9�%)wb� �����)91FË͸UZ�7�v��+h7��2fOt,\9Uܔ��3^4���k���T���L��
�k��g�{�A�W�Qa(p��==�7"�wմ=�B�z<}=� ����O�7�w��R;.k]�]��������"��r�턷��I���(�!c0b��������$*�\7���x��VIG;O�w��ї�z����$>���1����?"�E]qd�5��^S�9*�<��ک��ܑ_i1n���S���ɏgܻ���k�w�/1���g��G�l)*�%���v35?J�ϑ�:���\�Xe�g���<`NΪ��<��oe{E�o�+�o'E����vG��T���tQ�cy���z��73�Cm�LUݓUd�?dv*3,���q �3O4{�ڡ�ng����3/�5���K�A7��w��jNJ1s�Ye!����HM%��Vr�^PљF5*����ou���,�=T����#JY|A�EJ�$q��)dMz��^n����T��}�Zgu��	���գB1t���d��Ren�3s�鯰f��r�8㹪P=��/SL� �\�HEok^�=���iͻȘ۫<7�qs��k�$�HrMP|�#r�H�ȑn<�0B��7,�)�,�7����Kh�ǜ� ��JۥJD�ml�S���@��7���!��W}ߤ	�k1�0�ە�K�a<r�i�X�N%=7��9w/�V�N[Y7�*ܮi~�9o�}����gS�5't���`1��<:E�[u���5�Q��U�=���(Ghn���kL�s��>�!k�z�4��(�h�b��-��*�2��چN`\w����+<zW�O���==,1����h�o9�mݝ]����d
s�F4�Ī���nR�%�#	e���&���Kھ�Gz���]��'�7v��$Lٟ��^�\�gr��R6�NX���Tj��s�Ґ��#�X?��8���.��ڨv�U�2�s����u�������#�Vtx��Sv�ts �oC�Qp�`�v#�L�rmcӚv��v�[Ǎ�9G�$����a�����o�9!%��$-�]�񃽽�TvGt�0d��@�"I$�{M_���d��v���ҿW�4���w�J����k��H�RBs�i��S
��/n7��v�o�]u�tS�����Z/j6&��6�/x^�����-oa� z���6�=k;�eU�ˡ��Q	C�ɩ��ˊ�H�>�O���)ݮػw�M�K���i�v,>������#5���y�1�ť�އ��~ʵ)h1f�ܢ����8���	lD �3d"��l����T	�/�S�������}�D�<9^�o%jۛ�o�w"M]/��j�WS�0gA�m��(y���p��q��:���m"���ә,�PG<�$bĖ�
j�P/quM��z�"�A�%%V���#s�sSNf��p�m��~����!S�v�ovн`}r�DHX���]ݨ�IU۽�W4�Ֆi�n�&�l���I��N�y
�D�=В����d�Sus�d�YG�4%poOi�z�y>���v����Y{��#(��)�sF���H�����M��y7Z@`o�|A�O�F����hO�ıg�������3��E�N����ݨ�zG;l�,���J&�S]�߰��:O�ۧ[w�k��E�����7��1>'cX] �q����y��^���3�5C����ݭC&v@0nSܷɨ$MMO�"�e'��ɻ��n��:��n˛��0ߕ@�������b��}��M���|�Q�Ѳ���O�;J�����������vrYݶ&�8$������)��X�&�|[��vVS�c*�6���hgU����n�y�|wNk�z%�*Ε4	���u�m�LE/��-���Ec�h��4,e��M�ט�gͶ��3�s�@qC�
I�M$������;���ie�ρlV����ñ����t	1���[���U�zvo��ĨE���vr
�M����%@n���f�Oxm;;�3�A�R�m��pG�v�N
Z����t+���%]7�{b�=�5�2�p�b�(�k�z�x~���[K�]d5}�	کh�j[�{:�i�n�a�~G�~E!E�T�$q�i`�e���\`:��5��R,�fuoe`�NTȃgj.3J
���J	=KA�Z���t�nΪ�����{�7B?�������Y�M���܇*e*	T!�O%�J��1'��&��H�y~7�x�����T�En7�]!�#M�I���>]�%o������_����B�9��,[$+����85N�?PxgG��N,�����j�vh��Ƽ�&|O.�p����z��!�au����=�j܁�~�:�*���8r����˭6�^��3.����+L������$ѽ���ʻ��m`�ø�-cM����]�DsUYՐM/9����ˢ]����\�󝴆�˶�ˌp۠vۮ���i�q��ξ����R�b��	�7�gq�5Y׃%4ei�1|h��^pU*{����fN^��~�Mǧ�kW��~���l��/n��䴔�]ӫ���ȾX�{,os��}^aW�t��ޮ�F���]�HW�d������0�n�;�/{���
�8
=�7"�w���=�0{4Q)3/�N�v����e{�r@~���t"��/ޛb5,ǁ�sI0����3�R�7dq��v��1��:��0'�:��\��%�/a
4e�ɔ�1�'6�O������������rr[<tQ�վs#a�
������U\��K���kw7g�S\�䏅��=�a�d_��� 40z�o3��lzӼ��l�d�P�hצj�e����� �B|����Ԉv��ʲ�}e������=x���ꧪf�P����,�_h�Y���j��U0g��LxN���e���r����wFWϜ�Bm�,�a9�<;��O�L?ug��Z����7��Ǜ�b���OS�7֞��"�ʓ�zompWzwZ�Q	�%.��A�����gQH��OjaW�h��P�Vq���`aJ��|�r�;�2j�"��>�;���
�:�}&�#B1�q
�w�p��F��������R�{2GM<M2��Y	"���LO�g�w�����'y�b�+�%^H�$��S�n�3$ZH]�iR�1�d�Yݻ�0�6� ݎ&�ܒV�ޔ�:�[>j�23
t�-4$����`:ϟ�G}��Ш����J�s�*�ǩI�R���k�<�vis��ݪ���׮�~��d�<�t`���g�݉U��ܤ�艫1����c3�nv�%P���`}�!�oP2U�';+�r#(�?5h�r'�V_b�[$m#y;��4�L n0p�t0���l�G��=�,V�⶛?�����RS�dgxu7@�������T�"N����3��{8��u��^CI�-H�~��ђ;�{M�6�#�i�{�;-\��W���\{o]ӄ��S{%(�uN�UQp��W`��ju�V���N�;6V���lΰSmp�mY�&���{��_[�tr���Q���ā�b�첚t�f��*%j��6�s�����6���m�/L��:_h6rc�nѸ�"���y?`�i����d���	��� �nw�����{m��^\��Mr���#E=��iW�o	��;2�w�p�H�%��C&�������.�|f$�y{��L�tG���'�r�^�,Ͼ��}�
����_�X>����}k���/�:��X�&~�`���-�yj$-���֯�	ᵙ���F��*Iu6z���ӗ��R�-.|{�+&���盟�Y�ߕC�{3����Z2���S�i�|���#:�;�@Xn�ޛ�[)��8D��7 �::O%^��ګL�׭��j�:�h�nKcR0L
�Dm�P�K��2I*_Z��8���<Leonj�ܹ���F�"�D0���
[(�Yx��Z4�����=�5�)Uձ{}[�gs��	��aNA�pY1�w:�q>�G������x�}��w����{���W����z��_{�ۮ�xQ%�6{اhg��[WR�N_�wW.�8��������	��Y���m$���KVVT`[�R��;���g>7�;�Y�H�|xXW\�i��������h=�J�lj�:��P�3*S�����ܵn-�gH��5��N���fw�y`��V6����j���hR�-�ՠ��ոo9K{����q��}��_Y*�Z�7&֖m����p����6W]����6�E��O�}�����J��PPS�o*ˬ���N��ې�����C�T���;�=[���l�0l��#�k8�����{@Y�M7rIw��
*H{��*h��*�,P��>jjy8g����K��J֧���8|�v��*���Z�;��ن]��w�U+��+�p5M+YG$`������|��n�ݜ��e��V�cZ�KS-[�+n�U-Y�.vًS�4;� �t�����As�N�f�X�ʫ��nȫp0^ ��p,��-�i>y�Ss�n��+�xK��q^�p͖z�ȯ"�V-��h���0(4��u=�.43��m��5s5g6k��I]v����V/`lȐ��f<���h�#y9�+�/hJ�gI|��+�B��U�h��2*�a���;ΟN[y���r�d�P�{R�>������Γ�܅�.Q�Z�3v�{UJ�6D�S��[�V�Bm�7��ަ��O*``©�휼1����3;����:N�x',ԥ�U��i��{���V�n����$�����@���1��o#��1ďom������*�'#sD���	E�	�0�s 6�g9��9�欤�ΐ�CZ�����L�Ѳ�U[�ƭ�De|���U��Q˳G��>�sQ]��c�)\w�WL��:����C$�z���ԺǨ�ѵŮ�mi���U7c��&�טw�MQ��NaR���m��76�8��6UD,N4r��j��B�x��:���B�U;�d>1T�tJT9cӽ�L�j���;�ba��'�c������!ƙm4w_v�\���r�Sʴ�l�$�'og	e�͂�Q��JwQ�y��-�g
��O:>�!��[,��'[�%������v�/)^�k�31��iۣ�ö�����s�Mxo�Y���a.l��*�_��ֽʙ46�1<swN�.5��CE���B{!�t֠��㡨�Uȇs�\9�:l���.eZJ�76b�7*�Y)G��*��2G���ð^8�-�����l�	�y}�;��d���C\�����[#Nqn;�{_h)�ei8��<FyN�Ro�;��1��K��+]ȐڅM��v9Vw7����&j��.���~�ش�.��t؜u�۹�v5c,����"��J��:;���'Al�N�itk9����c�j�p�kOTuʄ���e�9��y�?5�DY����j�9�+�v��:�Y�.�����*�7��f
L&���������R"���M�z�N�4��\y;USE%��*�i)����J4�*�(�ZMV���hb)��(i�u��
��M:B������+ZZ��$���hb����ѪJZe��5�m�(i<O �Pjض�Fئ�F�4(�Ә&Q��h�PST�kI�m��j)"���5���"�""v�D�e��h��qf4�qfLkb��u�F���l��EAV��D�m��4�ѳ���F
�������CY�A�!�i4RPb&)i��d�UAkŭle�FH��ֆ��;b�kFɶ��i�S3F���t�[Lh��h
�;��-�5�kh"
��TUDQI�R|m�1Ux�QNɶ4:�ӬTA?_*��y�����(~X�'.�{N^CF*y����v�kv�M*�Smd��9�V��Kp�'.y���r�4����Gk�U�l7	L�A�ܽ׽�w����o+ �gړt�>�m�0���\��~5�?f�_����rE1��'j��
���wM�й;��y�q��~�

;3**�wTw��L\G/j���w%�2�be'��j�&��s��U�Ĵ.���`ʀ���*����P1)�ǨtI��v���N-gr�10�ٷ"�/Le�'�k;�3�L�1��	�>ّ�M�}�G����y�3`������}��Kݢ�A�Ϭ��;�a�Y��J�F�e���:��;1�ڥ��7{#38��fqĵ���ΰ�s d3��srK=�x��iv�m�����3Y�;a��E��y�Z�E�����s9-c�	.*�C;fVЙ7���4m����eOW�l�q�_ d��#�9��Y^�r�1�i�{�UǸ����R�a��D+�B.2}����PR)A�֨�a��=A3n�����W�m�`���¬��c!�ҳ��-�߰T��F�ݲ7�9[����o�B!b��5�ƶ�ù�����<����l�:��X�x�;ϣ��N�7v,���#gZ�7a0�8:�f�*o9���x/�'J���`�2�9�I֤*砠Ǻ=Bȃ�4ꗵ����
�#)gk6�ͣHo����z��'�(����g�*�@�	ȩ�"�ۍñvԌ���sW�4pƼ��3�M��]A$������iq ���x@�a�MH^�67�`c�W	���f��箌���6ɒyq6w�>�ϻ0[����c&���vj��@z��E״vAS@�\��Ůl�vʞ��\:3�7���b]?~���E��[�]ӫ�7�d����F���Y�}����g/:�ޡ�\�d�U{�)W�f�iE��[�T�9T�.�}��ES�1G�o@pQ�]N9����%�կ�f#�V�B��y�7���de��� o�Gy��`{N�� �ڈ��c&�5[�=���՛}oҨ���1�v��0:G4�	��u��?~Jn���� Pg�vp���,l�r���}�q�>��]xe�x�}NSe�%�k�q�r�\��vf��@���m격�뛻 ����5qf��+k3�������JI�$�M4��ڒ�j>a��D	}Ԛ��W��8Vg]�fU�t���l�ur����Z�y�g���K`:(�S�d�:��6�u@��	�s�xd��3�_�e�����AD@���گt[�5��P�`9U�8�MNrA���G�Q+ٛڒ9|H���X�A.��4v09יyw]�љq�ܭ̃,���U=S6z�#W�ˌ_xz����Q쳏���(����v�w�Q���4���_��0A����J��<�]�Ke�j7���ǝ��ѧglO,�G���=�=4�&��=
�����a=2��-�����'w���xϛ�HK�*C�j�-HܷSِ$Zh��U͕N���nj������;g�}����	+n)+ҧ�-���rM�W<oX�1K{�a��c@rL��6�������u�TzW_\%JM����Y��߇r���Β->���P����]�c�v%T.��'�{�"�VR�?���c���5�����y��/�w���u;�T{mz��������Sx��C�mʣ
����ђ���6����w5�;�����}��;Y|T�*VULs. ��K�f���Mq{�I��6�GhUd��e<�)qY�)�V\���(�<0�sO�j�o�����7�%�oW�d�M���Vf�k�g�^��7T]�����ot�ˑ�U� ��g�Lf0r7a���r{V
ƓO��M�s�-��o,�ۚ��̑g���J�u�G���`S�J��w*�Q;�iFwo�q�z�GR$'��="��N׻�����,�ަ�ݜ�փ����퍱��9�^�Ә2<6�&H�	[�f}�Z���s�����]�~���?�p�qe�Q����=ûٖ��p�ȑVY8�}������]{3՝�EШ����q�
6B`=���W]{� f]������U�"xJ�L���w&�{k�^��8;��=ܘ��c8|Wq3����'�N�%��4�N���Vn+�u~��p��F��-�r��n�����SaaD�=���$�t=H>̕rͺ���OO%�_�}?q:P���C��}�3�FgY���g�$�,9��+LC)3\:���F������r�R4�ܐ-кC����r��Ұ�*N��v<�̧��&�>��*r�� �Y�]���o�5�[�	yA�V���zQf�0��c3�wh��H��zN�V
ۺ�����nHbX���r���5aغCr
|B4	��W2�S��?A����8;����֓���
�#�'�TW#�|g�RVJ��y9f���D��d��o6���^|�/��`�1+rx(�e��n�%�2��d��ݧ{�W���Q�+&�/
z��z|ɷ�> �,�ղ7:OE��B���wvz�u�s�wA���H�ԛ�#=����0Y�z������6�V]>�'s�27M��&ѥ�h�c�B�ē�"M�2�����+����
�Ngc�Z9/8ԥL��=��k�.��5*o�2.r��P�z͠��ˉ�\vj��F�P&��@���Ԩ[<��9]�t�7�n�N�3����Nc��������S:	� �p��[!l�'��a=^/�mǻ��޽Τ_#x/F��u}v�,���g��4�8�pU��c�7Sׅ���(<�ΰ�D+�h�
�eq�}Rq"���PІ=��7�T`�a��v򾢂1��*Gh#���4�v��Ƿ��dMl�r�L�����-[
�m�4�.]+tc�R�3,rᕀ��0�z(��ȅۼ�.7�M����䜙98�����lo�g�Ҳ!�|6)�r g����$�v�G^*;u1u�Wz���;P���g��9Z�ϞEe�yz,2Yō���ɰfBh�%�S��mk�;�Z� �jf�kr.F���\��M%@$q�Vn(�a�:���/RFQ�> ��O/��k�&?M��>�wD+�@E�O���	AH��=i��j��L��9��vz�*){&�d
F�P�r.�5,�ځTL���L�|]o��ӛ��`��;w>�ndU��.�S��/�w�e��u�Mƿo���p��:����J�^I*��q�N��.!�'���dd�xK�V���΀�E�IXˍ6ɒyux�2ُ� ��Ւ��7�F��j�������26���S�.�Xe���;eO�stt�,Pu")�7ɻl�m<*������{==]�z����%4�X�?��:�}�f�AT@�Z>w�E"��<��=�P3�P�Y7��Km �/[�f�8rɰZWoW>�ו�vҘ��0�)��`08�]���wc�!@�{���'�_s�Ms#9�7�&�5K-+�*y�Ꜩ�3j$�����ˈ��1�w��}i��`�ǘ.���Ƅ����F�`�]�+�3F�֗cs�׷緒t4�
�7�fǸoC�����p��p�#;��'������y������N�m�N��.��F��Z�4�,��u�t��Vi�t����THo�c���c��h�|Ԍ�Ş��4�]���{Z��z�Ҵ��_� tH<4�%�zX���YT�8�P�Ʃ�z���N�X���lU�cٖC�ĉ(������4(K�6�����;J��)����2$R��&�j�2��#����	�;]#y����;�85��c����Y�*~���a8��y��\�><�$���"����	/צw�s��q��Ǫ%́��p,A���=j���w�g~uDY����������^�I����t���:��g��=�F�b��'�}2��Q�@�/��zBv�A������IN�V�+`�3{�U/��p8�����$Vܭ�s&vP�գe��]j��LD��юÚ6����6��}Ǜ���꛼��m)�o�f��^M�lWf>�AE,�j�w;�)�_Q<'J��㍼!�1���a�%Ięk����{ È��cN]��'�C
=�?	�3Pc1�(�H��RJζ��fS�Ե@�aDvg^�z�����sW	b��)��6�V��nWW�J�5-��H%�w!Q��η�Y=��9!�.u�:��Ĩ������H̾���[�gD����K)P���d0�,�>��ْ��l�mݻ�zP_��Y������'N�Yܤ�V�ކ2�،�m0+�J���:�+���j�^�a�4o��'�PK���] ��r�<����.�o��7��%?�}��ו�$���:��9�H�~�������d�c��D\�l^M��ڮ��b K8�HxXkd9�6��H9 �ʊ0,���� -I�p�?���~A>�,ꍌ��{�ve��p��z�(;�k$g Pfh{k�� ��d�utַ���5ya���(���F�:���v0�eP��m{�^�[�ܽ�%�ua���?���wy��Pt��hU82v�6,�q�]y����7V���-g���3)�v���E���wZ���d��)�a�i}�W�f��sv?���, �f�A�Q�.d_3�@B��z��V�U�m~�vɼJ��D���B���to��O&����0��M�1_���A\ Vkf�b�����}�;�S�x���('�'X�k�X�9��t)��K�Hc!�H�s�}��*�i��p��߻PW���hA됶�ji�CO7E��y����R��%�v�n|�� ՄOb�nAH=Ղ\rW�A�6�w6�>(~9�sk�2�Lbi�@W�Ʉ����#�RW��uѣ���1sYs�ph��곻��?_K]9�gS@El��u��u���6'��?�vtm���3�a�T����ŶS����,��|����]^N�ne>�u��G^<l�H=Xh��%�A3��W@az��m��h����㷫�Iȃ���ɐ;�F���1��WO�0n3z��js�(�Wt�7;�p�i{5��$��~�k���ktx�q��0��p�2c�9s��\˴Z���h�k�w�J煪Yz��,j\�t��lݬ��g\��%��cw%�̅7��S��]Ȫ��?������ײ�_a6Vy��fgc���O�pލ�'p��
�z�j�� ��;���D��T�C�������d�[�g�Eɟ�?�[N�L��Z;��|��iR���Õܧwt��"#�6'���4�w�2���j9����>ِ2B��o��G�ůý��'�G������@Jv��l��5��1��gc�����*鹦gsz�%�a��� �sK{�`�;���5�L��U^�DVD�j7ݱ�Mw_#�ɽ�X����hH�Z�U�S�͢;"�j�3�_��C΀�B�{�]w{jeJ��:�\��i*H�fҋ��f�-�3Qz�gV��ʆ6��y����ظ�D+�J
E(<;*�_���*a���C��/y5a�~D����<����XxF�S絲ځOqV���Ȍ�����8гH��Y��3NLa۹�n���'"������{}^�g������w����{�======��=��v�OB��P_��"]6���;Ε�Lo��<zn�;�5x��54��*����2��NY������K}}��Jg)ޕق�(�MIkNsӕ�j�܌ M�m��Y�q	j5|�ngp�!k��5�f-,�t�	t<�-y���.H�IJ��w^������^;���ΦÛ*XՃn�z:X�a%��Ȥn�K��ݺ3�&d!u��n��SQdR�,�b�(��j��d�/sH� s���Hy��1����ƹ�!��^ h����,n�2�=s��;��;���̝��h��q8��'X5�����0�C]�1G6d�W.-b��!�]!ـ5��t�8*iq��h˃kg�C�F,�up!�;)��{@L�Y��rq�a6�\���G��`L�-	�U�* �muEw�T�	ړgY��B���9�s�����
�i���Z�ʚ5Z�"ZZ0m^���/XΠ�]��騊�s�J�9�v)ɹ�(f_<��������V���hъ�:�O9-���qg��w�^�>"ړ~��EYW�3zi���z_޴h�g�H��%d��Μ��h�ƄYϯ�u]��"�0d��gn-�+(l�,xLԧ���������gP�-��QӖ��+�w�=���KY���Q� /wJ�g*!tۤ�k�"�k;��-�
��:�AS�V�+x�O!Wz��|e��+�A�� ��i�up=O�|�����}�f���DP��v�8qK�x�>����鉨�5�,�ʳ�:U��j��m�&	B"K��$љ�I��Fc���qb4
��V����,����XJw��-"�<9ޱD5֏"۫vr�zM.�o��q�E^6���nfiҙ�_Ͼ]��i�A�qP�Ӵ�-dm���\�����ʻ<�ô������H�;܉���6Q��'}�5�������)�\v�7]}��8Y��,!��S{�E�h�',.�F�������hb����*+S�Bŗk��re`Q �@��`�s�wh�J���6�*%��<N��q�W��D�J��~�F.V�H\ְ'KƉ�*��bk�k���޶#�w4P]3[�Jn������2�4S:�4nV�Y��gS�QI|�_Fvk6�2-Y+��^d��ZI:d�رN�����ݹ����T�T���e��u7���*��Ll�_!4��2�`��`�ث�(�9L��or������<pPE����w��NrG�r݈5�"��\<΂:�.�oI�Pee=2Țr�{��㑍䍨9�ފ�}݃^�X���d1��S}+:���koK�q�P��֍�sT��_9��`<�s�)2�6ti2���Kx,�"�)�[�u2fj�h�S��R�nk��^�g x�ڮ�\D �����V����Z�ʘν��&`]���+T�#���.-��;X-B^2�)`�� ��@h�Q[i��Al[h4���&�����I�N$45�L�hևA���LT�Ӷ��cthq:�PU���lhѶ��M����qTX��Xاc�i�l��JӉ6�LM�ƣXѣC�4���S͚I���ֶڶ4N�:*�5�
��������э�kE��b*(&��%���kE8���"d���
(�*�Z�j�����(��-�A��R�I�kEQIM8����`�UE4kkh'd��UT�R�me6ƃN64TPI�TQ�KA��S�1m��MKZMh�[&#[F��	��*��(��tQIQ�f���(���Ӊ�:f ��)����m�,� �(���h�
f(����1Dֱ4U���SP�l䊩����(��$����W=�(�3P�GU�<X�2jjnpE+������o����)`���WU��Ǥ���A���8�d��˒y�Y������_<L���$���$���=�N�K�"�:A�\���{�Z��t����w�v�u���t��7.4d�'�gZ���6�q�S1��Z��s���[0G@ێ�{(�ĲhK�[KZ�!v-h�V����[ݚ���~���+ʦz�����S u��i)��u`:���K=�z��6䅎���8��`0�\g�3���4h9]�C�.zh|�.񇻤�^��['iG�P��`��#6�އ�O-{�C�o��k��jr���c���o{h#�F7;hd������f�~�u*D��_�s-f���o�����-x޲�'��ʢA�&:A�2:�v�̝�w[4�j�\��v^��;x��:=f����L�Z\-W���U��p V��޵ D��8p�wl1E��F�z��N�ܲA�D��#�y��ѳ��8��a�E�ݵ��5@��lQ���y�����Cq���B��P�]!���)\�Ki箎�+��%)h���i���mes�"p_(լ���p��$��z�u� �q�t��S��SU�Q�z��N�Lj]u���a�����$���֛��&%����?:#�Q��F�j�.�#�_N�K��Q��U����5�G�+dV�.��`�J��S�y�����Ju��1�H��i�z�9���y�����4TJp���׏d\K��gA]��nm�S@U���q��ۯ��)�
�f�I�A�U�,;GM<4΁�	%�4�m2F��{&�Ĩ�xX���\���bL��ܷV��zKu���oM�������32C+�Em����Vp�J�t��E�M��w�����͡�6[���8A�+�z��2���%Q�\b��5��'p�Y����5��vc����3�AY�3�ຄ.�u���Q��&��퍷�[���;j�'���K$�7��5��V�{fJhOy���u���td�fn-��{�U�yR��*wMg{���n0Cz�`��?~��N���w0�4V�&��cڑ'11T�ԣ�F)�k7yn퇔2u��m�wu�chw֎�l�.<�;lnbV/J�`g]z*Q��H��.I]���+�+�۫[%42��ץ��t��e�oS+*�u*xwo���a��e��k�w�)�Oc��ڮ��:��V�\�a�Y��R�] ������B�2 3�~Ѹ����	����!�1p6�e�Tu"���=�ӆh�aR�-q�U<o���gts�([o� +�}���mq�d����d����Ys��{Nح�V睈9��:���ސH���7`��}�.n�xR|3�y�o-	$�����s�܌�pA����霷��#P�+V~��D�LR7�E��4���h&���/�Z�C�I��.2��L��Z*�qu�m��3&⳹,�<�u+<�[M嫉s~ݥ�`���������y9-�)>�S�F�=Q���u��Z2�B6v��`�ڥ{�����8l�@��fg���/ -���}8Gb��#Ύ�y.�����^��ڋ���d��h��S7�����2D%6C�|{�$޿E�}UU[�P��Ӷ����}nR|M�Yh)����IWW��֙uy��=2����I�30���?a�=fa��V_&@��qʈg6,�o�=�b���V)���%�p�b��}���YN�[��-:V-���ʃ�U⮻&�wFp@������cN�+�nUɧ����G�����T��pEC������E�F1ž�#i^�Om���u媹\��I�����u���l0��,v��ͬ���h�$��f��gd����kbGuIug��*��9�@au�3D̦vix]�{8��m��/��Dv�ͮ�յ@�b@W�'��ɵ�i���r�83��W�����m�����8;���]2���rZ�D�וg]�]j�C�i�w�n�D���#��#��l����s��|9�#i��(f�S��i|��������:Clo3��tm����}�4%�v��1���Z�V?��?xE%���:p�����a�Y�}N"�B�Q�=�=gl�>RGA����H�i��(���>; �(h���#t�l�3����]�+%h�qwH<��<U!��Z=X��Mkg���)���C���!�Ԉǔ��[���nl��d�C�1���v����xU7��o��b����bwBu՝�v���j'����^���w|�o��mN�ɗ��HG
gj�1�ܴ�F�u��k��i�m���ѻ��
�e.��7���V��r��̬j4�S���ᣢ(�Ua��;7"��;�N� k)#�����J4�Y��9��۰Ƃ���Q<"�$D,%��ٻ�y4MotW���$�=�^�un��P}�<7V��Z�J�Le<���3�r��ѽ��%+/$�FUz��۹�n�U�� �r*}����52�eM������i�Lt@h�d���s���T�UA�m���E����n�;Y��mnwf�nwP.FG��3���	-ˍ6ɒyux�-��ƻq����wch�W��8l�26���%Mir��`Z���1��o�Yȇ����t��l����YX��dl��v)�Q��JJA��0�/r�֮��ە�ެ>G� N�=m��]Nx�3��M{��{wjx�8�D-םߙZ�st�:zL��;L��3d��=�����1?���,�=oL��h���8{�Q�F��8d,���ձAn����a����՘5�S��=g{˪{@Vy�ba��=�[�z~�߰N\b�'*��!9܍V���v���5�����\��ȫ�;�Y�M�3��w�>��ҟ��v�q[��_t������߼�g�����lw᠟V��U5�;ll������]I���*��Nf��ulgv�7Yu[ �=^/���v|Lt����c����w���[AR:ݑ�a�c`�<�k�\��}àY�'����@$�x�5�2����Tf{�컽�l#a�"��Rzo�ܠ��JC��&�W�)��3�41�x�vr���J���1B(�P϶�"��.�#�m��s�w,fD��^��u`��+(Ϋu��PJ�z�l��C���s��W-��]�w��$@-�*Ux$q�����20��`�']p�b3�#�ݻ�%Ta�n!]�F�zK�S^;��4�4����g�3;�{�;pJAB0xEo�hґ痒*C�i��u6�O3����e���x�y�K�E�D��(m�G�� ݄��䒰�+=��ǡG�gQng-���{G�z�7h+������Ër���t>Z�� ������%�P���A,s%sg7�_tD�΂� r(H�&��R�L����{�#u�b��u/S&Y0�܂�K��ddܾ�yB��N
w�*�m��1�ut�b�^VU��D����T(P��xS�.�0�2����67��/rU�\c��k5�ݼF����9�6��������\ V7λ�����ǹ���읾�~䅿��#%$�o��P���g�C���*Ժ����_��o��Zf�{/�}ƕ,�S@*ݐoc����Fl��2T��f�>U���yZ8��L$�v�T,�ڶ����n�k��Zٲ^S]�giګ��ʂL��7#/�H�����)-���g�¯�R��w���g�i�:�l�wa�x�쀖��26���P�ş�VT�_9à��pQ�V�z�:,מ7���Ͳv��:|���u{��۬lމȉ�Z���/���@��!f<����{�n��w��5w�|���{�1�\zyQ�M7����B���ݞ����;]�%���J�z�^#�qT�zrd��v�:_>x���u�Vw#1���)w[���k͙AUR��;���.V�x������O�@f��w�tW1��OQ�':�%vN%�Qu�����2�'J�[4�7�c2�Δ�rw�ﺨ��[{&�0����M���,���-�()�JB]m>��"月gʇ���9����������wȎ���IU�~�bQ�]ʥ����̨�2i�ղu�r���"{H˄= ���>GE�\5�w^i�/�d�oj�܏s6U!���g����J��6���0w}i��h�[�5ul�R�l��I+����t�|5���dV��[Nc�ܓ��u�(��c�i�� ���i~n�+;dw_o��t�!�	�����Ҏa̭5c�dKeb�GǍ���:�%�-#RnF;[t�x{�������������`dGu��ӴJ0��'t����(��l��Vc{�� .���&{}�:��T�u��x�Gݷ��{N:�-w�R�F��Ц�u���#������T-/lt��O��1cl~� �3��/�&�«�ʻ�b����l%ߢ���]T�8���>��\�[5_�{�#{l���aK���I��SK޼��ds9�1���R΁��_�}Z���b�)^�M:���<��#��h�����x�y���-�yU�4���9���ۅ�}�.���0p�1��4����>�����d��}�`o3�G3��7�͌���S�F�]�g{k��R���ھn����gs�`��Ϯ���/9C�n������GoooU��ۣg�Ӟ�D�A�4�G`��/��68����v�W�rwp�d�`7�l�!�ۼz�U�#�h���/��N^׾��UP�4���0���Q53�ۏY�I
��i+eX8�}�u{��Mfyr�י/OS��n�����UT\+&��5��`#�rʩ��6LD<#�Yѝ�KA�ˉsb�E��φ����g�r�
-�J��'{�l@%t����ʡ���܍V�}V��'"��,#��\;�'wn�-�m���zCiF���%R��T�W�N�i3ʧ)�|�]ܻ��tp���O���8H���Cl�'�P'
���RUҘ�)��v�UI7Z�UI�]�6�˟����,�WBC>�s+�w��f��sG�o{�r���
���f:��&�a����[�t:�V�+Q������jfvēkWs�]k�y1J��u��=�|�FZ;Vô�����f���'Ӊ�G��𞰿�����c�p�m<�t�U~�K��Z���F8��'�oQ��9�z[s���%@)�|�����#��m�����3ֶ*�7cw��sոCs6�����djƂ�-� C6<.e��gU�F3��0[��f���C-��������x����<Fi���:2c���w�9��tgV�V��0WW���'��od��m�����m��3��V�0�2��i��4d�:ՄC;����8�P/���vI��u���t7y6���S>U����l�4�~��E#����f̂�#F�l3��j���hrȷF���٦3(E���b��}x*}�V���C���b�[F��B��?�n��c�*��D&��`B�y�ѩ����}�n^�
��&���� �"|tM��a�2!�q ��Ϗ�������_Ӳ9D U�Ъ�"�K����� D��*
�~����}�o�F`Y�fU�`Y�f�ed`Y�f &�FdY�f�dY�fU�Fd`Y�fE�e�fU�eY�fQ�`X`Y�f�@�`Y�f�e��eY�fE�dY�f�|lȳ(� L2�ȳ"�2�Ⱦ���aY�	�f�`Y�fE�FdY�fU�`Y�fE�e��fE�V`Y�fQ�VeY�fE�y�#"#�dY�	�fE�eY�fE�FdY��eY�fE�`Y�fQ�V`Y��2�³(�0,��"̃0,��02��3�0,�3̣23"� L0,�3(�0,��"�)2��3"̋2���"̃2�ȳ (�2,��̃0,���
̩2,ȳ(̃2,ȳ(�2'�0�$�3*��D̂�:���0�� * L�U\� *�2�ª̪����*�2��  L*�*�2 �  L���0 ª�<aT3
�0 � *�2�� L���g��� 2��
�2��  L�3� L:0,ȳ̃2�ȳ"̣22,ʳ�2ȳ�0,�0��"�2���"�2���
�����x1�g��#H
��"��L� ��T�C:�B)��*A��Q��%�Gi
�'8��~>>���}o�" *��������@U?��_������@�O؟��ܟ�W�!�� ���� ��?��8�o�������C�����~A��b��@bEaT�T
Df��!dT	XE@��P!I@%	R@�I Q�U�aUa` UY` 	��I
����"������������(P�P�P �Q������}B������}�=�/�� �������'��}�s�O�����b<������?�>� �C���'����O�T U��
�����a�1(*��>��|� *����&��G�>���)����O_ � �� �~��ϩ������  �OI���|}��c�����>=���I��`��;��� ����F#��� ���!���Ot=��/��1�`�Oۃ�?����:�'���D U��S��~)�?Xx�{���_��~\���QPW�>��
������_O/�>���S��(+$�k9�~
�}�+0
 ��d��H�o��*�b�����f�PD��(U�IJ��
�H�*���R�)T��TT�
HP��)H*mfVa&����-l�kl��v֚m�3��ׯ-�ڳ{d�a������el�۸a�j�f�4ӻ��7h���f����ju��jWmJ훷Wv�m�m�Z�j��a�m�Vkj�[M2��mZu��;����U�������S*���iݻ)m[V�a�Vf�і�.���u�铻��,�l�&��d���ẽ�vͣU�   v����s�׻{ܫ��oy@�h�����\�Ж��N�=ޮ��&�s��mu�m�;^�k[�^�=�������ez��=W�v:��v����N���7������k�T�[5b��Z�[,�U�L�&�m�   0����С��C�;�B���
��5�
(h(�=���ۅáB�
�\�o�\�ٯm�N��ֻ�s��λm���$�w�l#��Ƃ��wov���nzwiS�^��z����ޢ�������a���ܰmU��  N��I�wf�p5ƺk��u�W���W��mr�w�Wv�ۭ��ڪ{��nʹ�e�wwu����wc;�+���ǥݽ���l{��-�����/ownr���m��{��������]��Fѡ��B|  m}O�5�ںw}i��W��mN�z�[t�ܖooOu��zN��{^�ʀ��������^�p��F�E +i�tt:5:�.��ݵmlY�LU�۳S��F2��  \����5�V*���W@9�7h(���Ӯ��;#ۀrg;pPiU�5�@h�Y��֚��E+���5j�]˻s�i�Z�+j�Z>  ��=: ջ\
�ln�@*9s�+�WB��:*��Wu���`9�v�n�UmӀ��-�B��w5�v�o��n�U`�C+B�f�]�F�k�  {w�J[�����w]tURi����ոP]���zs�4=�]\  wC @`  my�KJk=��5$d�c��|  �|  6��}x� ���mp  w  �����s���s� �. �p4 ;����[U�+Yl��Se���|   >�>�v��� u��  n��  �ˀA�R�Ӡ��k�  �v�] A�U��4��Ǡ u��=���aƅi�f%�  {�}�� �[�  �K  �uwg(  wv ��S��  �V  n��t �����w  �S�)JT ����)J0  Oi�JT�L� )�CIJT   E?jR�P���R$̪�  M������o�/��k��n?��q�37h�����-� �E����xR�k-�k���}��U}_}�}���?鍶m�퍍�6?ݍ�m�ߍ�m���l� m��6<�����{�7���k��ʼ�:mKW�q9,�{l�;��@�Z�6�B�9l��)9FVZI����{�(�|+b^4��T�b����j� KjJ��V�	l �t1���؞˒i;> �۱$�eY7mA�9r��`�(޻�y�*҈���]�a�9eM���Ka�o7"є�*Գ��HW
�66&�f��D�A�+�	��D!�MŊ;���S%��V!̻��7Ie+Ϣ�ILu:�e�haʄX	�ժ��˻=M���ɚf*!Ĺ�d��w��/@�� �Ӵ�t��]����*��cV�lE����f9�C����X,,I��&S���C1�XR\+��s��J�ůD�߭&���y�������8[v�Vd�ҷt#���y���o,Z��t��u�QK75(6�2��,*f��3V-�oήVW�������8���m�mc�qr���J�Ĥ�xų�ኰ�v�$��x^[�)iBb1Tݽ�AF��qV���G(ҫ�p��͏3d?k6ն�x6�2�a��{
p��I����/T�k���M��ѩ
U�W����`%N�[J���e
ȥ���F��ͧ{e�w�$�MJS�L-0;�)��3Fq�R��%\�� �a�共Lֈ� 0a�Fzr`SK���Xs�𲆒��F�b�i79m�^<*��Ph�#�P)�7+&e(T@
���i�N��4���K�n�1�� ����ɡ��edN�駢TgB,#f�%��0- kwXӹ-2]���J��)���$�Ra�n���Zt�X�R�oM-�[�Em����Jq[�-%[�zX%�7/ ���@bM�(���J��E9�榯]h˷"�����{G-Q³&DCXY�	�$N���0p`�F�j()�KHn��:.pk��0��d�����rbaQ��
ځ�f�oqaY�a�8Cn�:��E�v��#nZ�3x6bnӠX��/z�%�#6�|�u�����+&����E�ie���.��{֗
�fjG*RW+K�D]�ٳ4��.��L�^�B�p=���� ��f��j�xma�ڍТ����V,�Z�\�?Z�F�t�⒊f	��@n9cv�5F �-L� �x�7l��Sj�ǎ|fx���YB=׮*���r�w#ԡz��&d��Fݠ/Z��J=� ��uc$H��5�+ �/X��C���ᦙ�6���t���h;����D��eh�L��4�]+���^�r��5,�֘6������Tb�X�xnK�^F���4�.İs2<̡�3ZJH�Yn���H�ݻ�W��ǁ;�Ң�,]؂�]Ҵ$�x��m�k�n��4*�����їX/r�	�k
C%k���ȁow7D����q�%�n�ݹ��]IZ�Ejˆ(�e�>w����m�2��#FX_(C/S��j�r�u�*z��ҹ��hI`�*Y�)SX�o�|���L��v6���JZ�m%n"r,v�v𫱠蒨��45-3>*Dv�]��#*Tܼ5�
k��S���� �[q[V6eY!�w".�Bђ�m�q,͕��G�B`l/h!*t���M�r����٫�ww7�i	S��Y�s[��r��n�7@��v;BL��3p�i-ԥn�TomMn�/A��D����ąmޔ�Ĩ�������Ê\�̥E轵��Y\v�9;[.�%�W��ѻ��mCz��V�oc��B0H��@��<�k6b�eB�*�Vߑ,�����$i&�b� � s� K-���:B`cF���rΨ鹕��co�o+RF���5ӭݛ��>ڀ3���#0�0aaf@t-#j:T�c,�J��,�p�s.��̗[ ��$���F��m����]ȱ�(+�����v��h躂���ߝ	�⹷J:�6��:�M�̵�L���+j���l�� Т���yr�&hV�7@ �ŉ"kZk��;u�ݙtہ�nfn0o���*Ɣ*�f9�I�oN�Y���|�ۦ�n�����e�*��ƚْae�V�۹)	�`�mڵb�"�\۰����4��$�r��*u�RӲ��k��)䢲R��S�t�N-�*ZV��óH�����Q�.��h2�i�A4`�+eAj�u��,-q-����Z�!WV��`l�^�-{q��ۦ���r�-5 �w�L����(�Δ��h��;m(ky֎Յ��v'kl�/fI���u��{V�:�d�*���A�{�kF��Z僖���0vGR�/V�:2����Gp��hȞA�*Ӻ+J5P�޵J�N�h�m^n䂅ƣyq�dl�EGXF��N#�D��[V�W.�ŦkeT�F7��U��VV�qf����MKJPj�5ì��m35�ѭ�Uh����ӫ�@���f�L�f��
"LŁob�ţt�,ٳT��h�)�7n8�NYE}���[��X���&,��:�vR�Ɉd��n%��`�或�H�PT-ɻu��v`ۉ^,U�gpe*x�Z+v � e]S��p́��&�����[�*��j۳S6ݪ�0$!�I�а��6�f(Vc�J�H��K{n]]輊��Ko�HhZն����N�&��Y&�=E�b�Z�z�XͿ�b� WJ<�Vsh��bV-Py��˨�0>ee*�����(�9 �#r&A;fm�^ɬܺ7�6XHd��&<�
�k7g7)�ā2$��P�pFJ/1){Y��/T��<�f��̼#�U�c[K�Ȅ�Klk�WpɖuB���Nm+�](��ћn�A�W[B�`�
���Սѥ\���]�B�T�w�<zUa��`�[A����&E��&��ݗ�4��mCaQ	z0�DgŨ��ۼK�Ơ��Q[�*�IԗK̽�62�1>QRQ���r��A��@F��kM
r��%�Y�MLiZ	7-V�	[J�̑�2�d+(S5���+�OU�V�'qb�z��!�����ӱ:Q�L����K7#B,1�Tl�2�6�*8�Ъ���i(7,��41i���E�!t� ���*	V�BT*$�X��62�͇Z �b�)��l3*����NFb�6h� �[�4R�omkbm�xe䅫E����lj�k��`��)�6�9���1�[Kv�IY[���MW�=R��T�1��f�zp��lP[[Aԙh���	�gjŀ�L���&��ڵ�u�+^�W�[�⧕��R�=5�f�ifSɘn1mD�b�Ѱ䲊lAk�.ʲ�֖�T�Ff
m`.! ��GJ����@ʽA�*�%m���X��0򈛶�e�fSG6��"��˔���S�Q��f��8p��*G^1�C.dZ�SV�tò]�7�gI6�̀��K�"��� �X.�����YdGr!O3��jZʨ&_l�ii9-���n� �"�$�Z#�2��X�@�&��6F�
nMr��c"���@,���WIk�����4 Mj���@H��?I+1���+X��'��b/~�H٧�,�t2�4h���Ҧ�]w�ָh�a�����Ȍ���e5Q�Fu�λr��6B2���7�!��˽q���"�ڲ��j0�3�훦6y�x��Kh͔V�Ȣ�L��w{A�4���*D�fh�wV��VF�&ࡩ�M�E=�� ��;Wm�����Z�"�d��lL�FTW�<"b�f���2i�(f:�w�a�d'i���������t̉9�M�ו
9,�2�X#96��P����ww`ۓ.[{��,�4��(��F6��N,�w����(�Rl���uwF���׎��eQ6Yʴ�BFQ�t��!�� lu�On�R�f&��*B�U�%�IV�9�v��`�7�+`X�:E�v6�L�yo"�e��n�ܻD$��m��i&O���QF�����+��N�1^_ۖV�ݹ�x�Sp�4bN�Y/F�����K�Z�����Ǧ��`��Q	SZ�4uE4ӵ�Q����mc�یL��R���UlT�.��7n�5U���XF�y����4����T&j]��B�Y��X��ef�R6)�1?��n�@-'�O������#6���әw՟���F����|K&d2�̰�
PڈeM��\O�.+P�4!�|A�P}c���a-N�,3��(�� ԙ�f�&�B�ڹz!��QT��k4P�а0E�& ��ym�jd.�b��2�(�6���Ac����B�5sչ �jP�E躛m8T�bc�Y�-k%��ظՋ���p�7�����5C%�{L住�0����V�#�92���Oq3oi<ݵ�����n�QB�E޹�Ǆ�HFѧ�����K&�h$��a�ʐ�q�َ�apIZt5�й�v�h��PJYu5Ԧf�n�,������	��ƀ��+%Ĵ��ƭ�xVR��92�f��0n�k�`/eT�)��Ĵ�E����#x��tc{Zw�J��Mfm�*�T�kRQ-��i��t���ь�W�AN#�l5��͎Σ�;�H�U�]A�X%�W����1CX���s-���Vb?\�n��l=P�8����(!1bЛ�wV�^�v�uzB�%Kv�b뾻���'�)�VJ���q���E�i��EL!t��tw>h�?\�R0xO�n2&/�r�͋[�0�i��!�q��豊\�xd�,��Ě>��ݑᕏU�֏�O* 0<TM:�)w.�5y��/f�@3�p(N�i�8�̩t�Ԧ�*ʻ����e�Y�
��Q[ԙ��t��Ə�E���S-;6��+)n/�Ɉl)ިw��R�)�å5İ���X�˭��oN����Y5�[si �㩮iM���[ˉ�"o�cr���1��@%QZ)�Ks	�`FJ0��,�ѭ�� *�u�����(V��abͰ�BX����!�3um��凫5G.l�V\0f�2���kL����N&�X���-�2��ԁb�*�m9��˭��Q��fm7o�e=��nk�N��{CA-��"���)h7nG�ci�df�Ȱ<J^�f�&��ퟒCY˦C���3pђ��@n���V�z�B���cX��2=��Y�e��B��b:�j���w���v�K6�f-ndOj}�Zo D�׉؅�2kT�+i��'ڣ�f^i�0R+U*B�TmUӢC��Vdϥ`�a#�6V�aW�S:l����Y��//fL%|Vꐽ�]l"4oB�kj�S,��p��6Pc7`()���.+�yO�i�śZ�[���+,��Y�AQ�ڕ��S�e�6�T��Nf�4������6Ҏ���mj��3u[׺�HRQ̤>��[�KkiJ�A���H2k�\��J�2��UyZ���re�
r�mٵ�<l�xM��[���%�S�/�Y�qC�S�W���M,4�%Rɱ,RZ��E�ujڭаbB��B�V�VS2��si [Ն�K����{N�։v�V�+2(Zt0� A��[gFLгX��dm]
S�6~�h�>� N�)��1�%�j�����!���[�a����Kc#7w5:�!FI�fm&�jL���+�*}�Ɩ� �X�
�}�63yIj��Ut�r�U�QvRԋN��S}�{f	|�fÍm�t�[��b���U�
`�u��Q�)G�T��E�Pۥ�B���4���#@��%�Z3#%v��̨�w�6F詠��4*�q9�P�h��T�e�jB7k�VM����Ms*Ҵ��soK!�)}`5�"�V,���*�1�*��S\	�� ׏fֹ�ˬk�m��,O��c[�s[�mD���}�)<{J�/!l�ֻq�Ռ��1F�D�T��B�ӠPhܫηH�<Ls��fcY�:�9Vea�R�j@��Yb�!b�4X	x���ST��j�X��Rb��J֕F��B`�V�Ho*��e,L�͘�����v�y5,r�뽣�a���P�7�Sj��� ��c�1alaɚ.�6	�-4��L
јj�SZnU^�Z�	�#5�ɵ*^k`�nѢ1���ȝԸ�kp)u�%L��Qyz��z�8��η
����Ҵ֛�M-�"�q��{"	Ka<�{�e'��mf�!�`LI��7[Mjܔ�-��0)����+]��Y�1-Z��jY�V�[����#6�=g-���V��ڶ�H�V*�-+̦�+2%"XV�����T�I�̩��.�i[dnHT ˀ�9�e�f)N5�FL2ȰA���DJK�EX�[+d��v����3���1�ҟ�;)�&��m%�,]mRY����F��b��4�n��0P2%�f�]:X�]0��N-�th���`�۪��e��G4\n[�:�Z(��l��I`�N�H2|�.���PS�:(��C��7RCVd*�홤�Iu/Rv�[�I�fU�Sn�_d�IK���)1sJ̷u�N7\ �t�s)[y���nZ�o\&��-���*�*f�7���-m ����1�.��mM��S���M�wrܟ,WtCڛ�h͛����7�B��K��G��[gJ����&���2���E���պjС5����m��)ag�en�'~���)i�Л�Ah�Qk�i56��7d�Ւ�;��ĂZ�J0�/taU��MA�#n�5i�C���S�����H�T������%���8�&�W�,�����i��]�n�k�R�]b�3U��髬z����r�7�+G����l�T�m3l���4S� �Ǆ��4�ݱYL��
�A,�*��)d�͐P	�1��2T������6�.���[�(�̘��Fz�W�&f\�Y�\�ɒ���:t�.�!�{ڨ�M1�^=�bǧ�82X����ӂ o�޳Yd�j�&lw�V*� 3�ݮ9@R�i�k9oX���8$���B����]���	�f�����3�1S$�I��td���h"����0u���؏_	A����W�U/QMcU�a��_g�s+.����.f�3��\�@�K�{&��,��0��u�E�Z�:�=lSL-R�0�)^���	a����Ύ�S/���
�>AZ���r��3���c�T���}
T型�E	��^�m�޺n�Q�{E�\nwW�K,:���nz�IoӴ�Iӭ��ʼs��B����TQ��c�Y�ά��*W1�v������k;�e��������uq�_4�(h:��F�[�k�.�ޔ��*\4�O�I�fVV�}�8�N΃R�c�D
ʧN�9�m������;��q�*�)���/����sT��03N[�V1�- b�j�,:9X�r�۪�=��=�\��;�NhE�QH�ܮ\n�H�/`PH��생v�VNX��K[�5Ƶ�2�PA�/��]��XIv�7�gb�h
�m%\�l���|��i͹nD�R��u�mh�p1���{v5��S5��x�R�]�
(LM�%��ի�LcF?�A�Au�mܦ�:������i�K�)J~���,VFS�{t˫��c��o�Os��A�]�ŖOb�b�wȶm*�I���й��>yX_M&�=��߉nZ��<�&�����6M�a��.\�|r�a�^�1Za�OO^t�B�KW;.�>J�&�gKy�A�ӛV�Q�־��� t�v�:�[�W��;R��wf	�]��,ؖNu7zU��0_"���µf��p��}��tO]X���[�(����A|�B�}u������yS�P�j;]�r�jon�L>|sGu_s�t�nZS�Sܜ�j�Źg����A<z��!���B�}��앩�׺������Ѝ�j�8�c�[���`21N��	Bt�b� r9Q�ĺ܀�Y��;,���y�A�j�+ 5 C��/X��c��d������Q}�EM�9��\]:Ժ-��v�'%���v�Vi��,$lϹ�E�ոo{@�9��"DΔ��}w1=U���v�gL�X��ٳ�d�N\&޶��[f$���+ΐ=�*�B����q���O���_Z�C+$ᦩ>�I��f���c憟��V]Fs���+�9Z��u��\��|�PڻxCʊ�Wlp�;F@�uq�5>Sr�3tܙv�{�u-�Fe�  K`
+��lQ��7��v�𰲥��Eǥ����^�9�
�X�oE���k4��q�*��qs��J���WVP��R������T��N�����6js6�w9m����9j,v��
�5� ��NJ�ٕ0�)��+�Ò\x �������5�z�]{�����Y�1����i� 䩬9����y��Cc�w88 ��1)�)qcH��.���]��� �:Dm�ds��M�7��+ ][i���O�D���n}w�'�CP�����\�z����s�y��M��
�rE�����a���w��E�޻�a)"W:_K�2{����/v�0�
�nf�h�kYbhH�ÖE���>�3(�k��,�����a�=�Lv������������j�wo�L�E�+��]��c�ѫV�:uJ�+�M�:���TW}�C.�T"��ٖ̭���F�d�DӀ��F�N��m���c�ڻb�����Ok��h!�f^��Z�o��V�٥V�F�-Y�X��]�e�Ҙ��Ôؐ�Q���VS��W��Y����i�:�Ge�����0_}�u;A�D�ŉL]�gr�S�#���S������ÑX��	���B,��MB�Y�{����~�#�̖	�j�j�r�ce��'Y
CzP�'l�U��2�l�'��r�7 �b\�e�����>�x���N�ҡ�KN\��Pj�4vVZ!�� ��V�^:������31�jحQ�R�l�ڍ&���;�r�eH�$6��&�n��K:�X���h*7D�o��
�҅ԈwcU�ٓ.��v�,������}��R�N��(�Q�{o:B'f��t�*(NI�o8�(m$�AE���p�=O*�G�/r��\�k�ʶ2U�a6�0C�W���O�����j�bĨ.j�]�p�����ݰ��WH������S����sb"��Z<ΕG����g8��]5�gr��ͧ�H���h[��*�T#�'�����*�
�A�5|(L��K�n��StF!a������ѻЛQ�R�� �ЁԘs�����f�$�ʏ��B{E1$^�9�r�	���ڦӹ���8)n��B����:�Ӝg��ȥ/{��pΆ�^fE�+Ʉ��������/I��ZD���[ZW7�ak�gr�xC�j̫T��j`ɒ_P�.����bXv��n��R�Sյ.j��u�����(���ZtV���7,VW���,�գ�P�Im�H�mwr����:�oTm�vĐ��!���C�EjL�
O3"q䓫S��0��R�\��!�n�q�u��EV7�I� *Yc`��PeAܷ;d,{j�w�h`�x��~�R�����l�������Aew<������n`��l�|���R�WMǂ�.��캹���x�Y0	��0�/e릃++��e�	%�8���˰��v�_Y�P��E�ͧ�����ۣ��.{&���*Xi�"���qWu)��4�<Æ�:�mW4�2���8�#+�mj+JĐ�.�[˱n�ũGjUα�v�2�1���$k`�������G(�0q�®��(*�s�Μ�[yZ8˩.#`Sҙ<�XUk5��X/o^��\��T&�ך�]�K�g��2an�f�ŐWK�2`b��i�ͣ�����@֗�[�×�][Ɓ8�})Qh�nc�;�L2�q�o�W�݁Ju:T�VL	�5�8,Wi��
�B���a絝�	R�wm��S�ۖ����U�F`ҏ��2��T�X�թe�5�)�l�*����\P|�V:"��Mu�htE+B������o0��\Y`)��\��%M��!�]�fN:t���p�s�������͒*SM1�;����1�w<� 7��q�-NfkZ�oi<�n��	]��m��wP#�P=\\�����=22�P�.sa/�i'��{��H}�W8�۷	Uu%��v$��F�3(��j�E�*�zn�S)���Rk8��
�2qZث�T���x�X�9܀/x���MNN=�������G�\����:ss:�֭o�o]>����v�cr.U���t�U������͡X)��6Y��B�UtU7J��v�$�%6V�N����ИW�x�3:Q��21���a5�,������[�v�F��L*{I��s���S>�5PMn�;�U}x,ao�� :Py�ڹ+�[���rAj�M-|�q�!fm�y�T��+��KsG\k�u�f5���R��S��d˱��_	���ҫ�1����d��LXG4Y�y0���m��i�ڦ$ჳWa�6FI���&dD\T�:�m���Ԗ[�suv�� ��2���(v�}/%�s���]=L�v�,��k8�,�Ʉ����� ���At�h�j�)���{V6	��L�Cqj��i��+�. �;�oF��K�,h��zf��8���{��=�u����W}B�G�]��%�"�,�.�z�ް���:��z��6�W˱R��n�R{�`;�m^4�9ϥ��h��%:Vą
u�r�ܷ�����:$�E^���VS���븪�}�[8q��1�٥�������D.��ˬe�V1�v�ۦ堨7s&�]�vgK���zm�h��.���EE����=6�h�M��OIXUI����t�jnZ�G
���\%���y�ұ8�;_0K�h�7eM���,d�.��Z��;���] ���w��Bj]Ag%���kr��ܹXl$8�#S�c���WCc��T3O5oo{�+pȹ�rѼЧ=θ���.��m#�-�����u�+gu�ó�̋.���Q:�A�99�zs'A�b�,���dU�6�2��ƨ6��h����觯����k�\Y�EM�y·�(����r�:?Xf1ۘ��ͥAuu��mڜ��"%��b��Q��z� (Ws]*ꔱf�@�p�qn��Ū�4���t�Ve8�n@���W	���w��ww)`8�g���=ʼ�TYi<��9v���r�]/cP9�dw��]�
h�����w.X��I��UY�\��|��۷����r�;h��/ O���{�r��̏)p}�1):�JVM�r�j��:lw�F��3�
�74P[9*9������,si��c���&�䓕�zq��M�۴�]�y ��o���0n1c,�A4^#�B��R8wuN���K-y�ӝ[F��n�pǷz.a���|���EH�o9b�,�ԓ��koUE�=8P|n#Y@<���J��_G�+:�"���+��� ���)�Xu��F����H�6�*���g��C���N��wuk<%��'iԼs�������Y��H+���Q۬��]��|��|��~�^76�����Ի\���`�IP��Ӯ�S��@c|�����=��r`�mH 4i�W(�vh���dX+P��9]%�cT��6�C�,��jo.*�\�H�R��0���ȶ���]g����d����3n1ʝ�Dt/c�y,
)�����S&uN��ܦ�6�{ٝS�\��)�o�mܢh;U2�ek�c+��6G��UJ���'�o�K3fa�%Ɏoz��$!Y���Ɓ�p��*��֔3��d���u�)л�y�5x� @5�
�L�m[]�V��[X�� z��76�o{��]}�ۭh>�#�7sBZ����� ��ٌ��Ҹ+Gb���iA�sI� ����`��8�ﳫ)sU�]b+<��q�x�c�@�\���n��Ӷ�J��#����Fw�ŝ���M��e��3G(��9���ٖ�O��w��~2��ٳ+
�Ԟ�yH��2�ʜ0�`H"�^��e����r��
K��o۷�� ;Ҋҧ�-9��Î�B���oPy� o��y��JMw���VM����Ί���vS��E.)ԜXH����T�No�X�U�=��k;�V���Ol*�ڱG)u�rWY���H��Ap�E⬮�.du�ҵ�F�+���.3��S� �.hX{�sX�-Y_zv����d�kM@���]�+���Rnǯ�����8�k3��]�¹E�X�45�Ϯ�6�F�1��2�Z����N�;$x:̎�Ԇ.��)j�)�� �J�f�k7�/����9Iް�Ȉ�i;	J!,��+Aw�]*��CzG�MV�˄�'�(��x�@�fs\ã��������������b;1�:�a4�Wr�lʒ�I1�E>�D�U�}x&�]d1+:�:��"��>�Us&�=��T1e�ҟb�κ��G0Mc����3��X��
�1X*��:�'s�]/r4﫶�,
�)�]`�E���Ø��JP��:�\�B��E��jL�n����֕-�������j��FI��dW�Ɨ��"i���/v�[Ԛtn�yf�*� {��e��Msn�b�D�v.�땡ZeuGYL�+(\κ����I�E���]b��]1�۹��OD`�,�%�Cc��/�Ї[K!�鸰��:�l5u�v��e��T6Wb�
Zī�G/���3k�wo�Ԧ<������T��!�Sp����F���Ru��7}b1���+4�5�u�w�^��ޜ�R����ůt�*D�μw�!Xn�w��wXV��&	]��[��L��|8<�S(�ے�ZJ#��4_m�V�-��
��u��C�s$5�{c`b�â㯯-t��ij��W��{�\d��.Rj�q�t��7����qz������-C��B�(�5������U̎��˻n�*�<��x#���K5��p��եhe�,�z�U��#	��E�'��Á��&�r�g=.�&��M�@q�޵Oj����dS:rT	o��U�xR�6Fu�6
&k������#��8��@�X-�I�[H�q^Lre���`��]�pNX�����0]�Ӓ���z�rb��X��榹���c�k,�Z噧�1�����������`���WcMS�5\1��s�)����e�Ic6��\ڗ�{���3"�hE��o��V͞�W5������I�`ư�.u��;���־���U�8c%�o"@w�xi��-��춒�Fk�P?�7|�^dx^�aNkm�R%o�Ie�(�u��2-�����$�&��O�5��EU� vS[�>����h%s[]��C��d!�|$R��h`
�Ү�(��f�v!�3�}Y2_l,�p��'c�mo��r_M���LX�׺.T�7�9&0�슟=7R��C�MAh�j�G������\�5!�W4�i��K�59�2�41 .NC�	p;��z�2��j#�R�]�k��@��Ԑĸn�����wP_��-wS��P��`�tFwT��֘V�����f�*qw�íԻj�o�v��Z�։ȃlE��p�pڲe�<%uX��)��vH�Az��p��o�Y��9���=�����Ϋ��s���!"e�=|fw64��x��q� ��Jػ�ۣ��4Ӻu�kp�x�U֞�'Pٕ��Eλ� ���10�Ԛ���"m��M9��V!��[��؃���@��|��ud�O.��Ѣ��Sxۉ�M�pO?�}�}��G�G�}}��_W�|�:��ڿ|Ʈ�)��E ����:�96K�T�.�)ƕ�_S�/0&3-)vZO:��ڊ�E2�]=�e�6���˥[������gh��f�*u k�tp��HoG������D_4����>�,�mx�r:�KH�z�f���A�:DL}����ff��u��6���7"mũ\��O�%�`���u��WX##̥J �܈e�0�[1a��*�9�b�W�G��85YM�Ool�����U����Z��\k�1��y�{O&R����Q��<��VT彻j�c�Y�	
츐������v���-�e���`y��)�����9؟s(՞=}u��v4�f�r��� T�T\;SrM�C0n
�+�'T�Ϊr ��>ƒ[. Uv��wwv��(�g6UbXGPZ�o��+"��+O�N�N�5��v��B�U�yf�F��y�.����\j�*�خ�هMv`����9�E�\W>�G�k=�l��f�"n�#zUԡݑd�7����JfV����&���������5�9ۉݐ��h���P���l5��<N<w�����U{�v�l��,VnC���V]EJ���{fT��
�Kcy(�g,�-�ψv�o%"�c�p]�-��V؏;XN�٢�;�:�H�l�ѨZ��KFe�|�Nm�0�:��ڻ�Gn��e�*�k��q�N,v>,x�^��0��n`>�Fn63�Y�L��`��\R�q��EmA8;4��h�Ϣܫy�su�ٜ g�ī,I{��:,);�g�F��=�5�0f_ת�.��t��1q�4��δ�ga�5휺�]>;�aȀ��'k��Qܫ�Fb���]6�����i��a��F�Fl|�
�(�ZY�(�:���l�
��w�୔3a�D�Wu&X��=���-y�@E��5��J�) ����۸��}-_2�P�<͟b�2S��W!<�q����YV'x���\���*>b�U��._]]X��7�F��A����=u�Ib\D5S��Y�n�\��>���BU:5V����w�G����Cq�╁A�Qc(���?�:�\2�X�9�J�2��ON�&ʸ����xj]���)��®<ە��S�t�c�b�/\4[R�;l`��9a�
�+�"��E,=�hu�Y�Ջ�.˱,+��r���N�Z�z�5�YMFN. ؔZ���!M�n͚�%�ϖdxT�1��Fv��p�0��@wISU�x�l*}2�L��]�'f��4;�
�A���er7��SX�ٚ$�p�r�p�)u�2k��&�Fވ�8��(8����J.��s5���4�K+���ϝҚ������sI�ԯ�	WHbtη��e���::Rd����N<�he��0�=x�.\��Y|�+q���0�ut�h�B7���@�(<z `×w{�.��{2nW
3WEF��r�+�t�m�=N�'K�L�d6�kV街v��G#��b��suw8��-0��xDjQw��J��[��p��j�������Ap���])2ƾ��"��X�)Η�ͱ2�����n�|`<�V&l֋�w��M��{y���o%Z�����(�Mk
�Fv����:�t��G����]�1�`��2w c^'Cp�$
vL� TJ��{^@ț����PМ�C0n��Ro�xR�N�F�vڌe_j�mb�r&���$=E�n:�-Q���t�r�%���@�,H�
ޓJ�i+���^Ո㴛�=��W���k�O��ط��r�vv�w�o���h ���&�Jz��K9}3�@�#Τh��Uh�n<g���\��w���s��%�Wv�G��sM
x�c#,�����ٵ��>��L����������p�u���XF�cy�����a�M�74U٣Q�ϸ�ɺ[uwYJ���B���-��ꐚj	l�un�V�%����[V;�"Z���9Ѷj��=���%ksz�4�r��8&6����S��lY�hɍ�7JU�v�T����S��r�ȝ�;��Y��k��_�f�'Y�%S�F]e;�x�aVwiE�/�\�������+n���l�X�'N��Txk{�bX�N[t�*�<��M�2��J�H��+v�+��=|�Zx_L���6��*dP��ǯ��,K����%;EK���oh�R�}�`�Y]a@f�>Ú�W���u�d�'��Zw����/��!���r�癹U�;!4�:��fC2�;|�RF�R�g,�X���[��/�;dOE�T-%=��6�;�yVhY׽�<R��Œhܔ����PT�a�E���a;]�&i6�Xp�ҧy#��u���2.����fu1LX�R�\nJ�R�\>�+0��1V��In�kx+��9���Ҩm�6�:Yrk���u�����]!5��lom��f�B����Rm�A���G&�����B��<^q(�t�=1el��`a��1G؀�]��+p������a�ܮ�ĽڮT��+3�jm(��*v,��MN��]L�����11_m�<+���]6飑�]@;�L��滒�P�G�E���x�pj���|�_êm]=y,���9h*ol�M��)vbE���M���9t4[���yG�t�O����l�Q�͡������{�N�:��V��#\����I�6����%/-���EӢ�fM�Rp�p�L��x���4����Z�i��%p�RI�)���o=�'g�03�0h�H|ɍq7�0oL� q�� *������v.�ݩX�r��]0�yo�K&�T+p��=��|�eM��H��)P:0i7E۫�a��1!�X���*TU��ve�a���ݢ�ɖ��۴2v҃^��j�'	�Y��_m�|�I�3���Щ��h�Dލ���k��������	oyKL��x�VV���v�걌ڐ_;�5�m�+��:���@��+E.AՌ.��&�4�f�$�f��}z~�mp�ը��P/�hO���v�;4����}4cI\L��4��ݰ��x:��������4�WD{��+Ŷ�zv���4��<Qа�%��.H]fھ�*�nէZ�[��Y]�R���6en�E[��9]�%u"pO���W,(�urfN�g�E��m3�y�O1�Ip�*�R43]��ĥ�l�.!�m�'�n&�7R����l���/7�m���B!d�Yu;Z�)s����oB�"��-eN�k\�Q��bn��Caաi����V,![�P��$Vq?5'[��u����q��;)L�"6p���j:�ؼ"GY"��s(].��[�z4=�6�S�z(�"r.�v�Զ��ҡ��I�/�|�[㚗s1��\�>ɢ���eҢ]�#�5���@V�
�7��܂v�m+J�n� �ݤЊv1{]�J�S%i.v+��i4K\��PޢibSkh◺e��d��a��w] �i�
����At�)j�%Hz��A[R	+�j|�)]r����Pۓ�P��������طg*�`&���9v����Z�%T�<�j���Xj����.�l��X��x��R�K8UX�@@.�P�J5y�Gt=��Gԩ.����*i���]�"���JN%�V"����r�K�zq="u�xy�Ia�YQ_$<,��A%axKz�ZJ&fU��zV���˼2�ncB�X�f0� ���c���oo��Z��f�0kH�r��4Е�Gc˳�*���� pt�Ån��[�wN���:s����hʲf�2�Ǆd�nZƞ�n:;d10��w�΃�͒'و�E�0q�	�ݐ����%S!쑩F���t^����GY��ޏ��Jg5��K9-��[�ToG\�tv�#R��B� �B�q�b���挬 �bt�\\0��賕7,y�h���g;��Q����8�ŹLV0PS��NSy�y���Z!}1�m��V�����cO��4Uң6[��[�ˮl���*Y��X	w��p=$�j��lG�	�[]�3�.��d��͞���L�YV������:�s��]���;)u*
�;[���OR���ݼ,�엎�>tꈷ�ѽ�!z�+Q���f�ݬ��#�Ǖ2i�7��\���a����k�p
�Z�gkt��� N�*)#�
Xc�z� q�&���b;Ft�㊞�f��ѫ["tS;Wr�Y��c.-��\z���݇^���n+%#|��9���12�<�^�C�w	�`�<��M����AWr�Ma	n�Tn�̾Ǡ
���S���9�Մ��7�=����r۽XG�@bm_0��e�'�u��h���g�������L���%{#�ёP���WX�f��Kl�z�^N�i8�h��>IЖ�#.�;����m��ЋI�C`[[ �dچR����RN{���۬�t_i�t�j��Թ���8J/w�	[n�
��ϡF���6�k�'�M��A��Z� [��(�Ċެ����Z�"�[P��J��B�}\�3�R׹�n�W��� ��\���KlvS�]�S�Ȼ�R�n�14R2���,�-bh�wj�oP��Ɨ�e{��VI4� z/�XK��� ��	���λ|���	��v�룎:IQ�֤i�;S�B�����įT��5��Z�T�G7X�"�_\xgrZ��K�vV>I39��{������O�Z�Հ��s��)jם:V��i��m��,��ZiS��fU�*�2�]��(���S0ڗ��vej�`��&pZ��f6�b�Y�R��i�r	�}�sP�Hd��I�=�rJ�v(�3�Mܧ[���A�W'u��8��:�|�onC��F%,��ʐ2�f�[�sGw2���/�+Rr$�*1B��b����(]���X���U �G�)gL��)��Q혉�t�z1��D`vƒ=e���ty�'�r͉��6�?c��L�i�i,�^R�pj.����S��"�ެ�ڦ-�o�j2�l.��ήWIM�n�]�un�nݴ���\�&�!�P0�h�-}��;�N�|�0������>PkZZ�H ��i�X�,�|����Zv'�r�'d9[��*�P'�Q8�S�7�C��CG]s��s#3��������OZ瀑����ڶ�ud�������S�p��ѕ�/����P�A`��M�u�e�7xg-N��A��!t��}�j�oBS�֑�WCm!e0���b�4����]W��U+/+^l6�n�"u^]��6c_DO � �a:��Vp3S��!�Wǝ��ï
�/X*�����N����Zʉ��2��K�)ڎ�lP�#V�LQص��*��Ku �V�K��kz:����k"�\��wo"Ղę�Y���&�����[1����5Z�T����k��$�{�]^���[��K�V/������4�4�:O����v6���P��b2)� �	Y�r
�u�������9�;�i�wG��
�ꎟQ��HD�uk�s�Q����t���&E���\�]B�ۗN��*�^��}�7����u�W���׉6��\�R�&b��a2��=ThE5�uuA+z����.+�������Ӯe��N���5���"_%"UѦ�r3se�;)�o(��k���\ Vw�^5{W�Õ���o*0"����W,��	5���q��e��L�%D�*��Zs�j{��wK�(hV�f�/�t��9E����5S�c*�D�:,SWb]�H�������Y�����k��$�����]�Λ�U�~]���\k���ܮ/R��`��͋����BL��y0�W�y--��������W��*�r�8&#"؂�N��F����;�i��*����S�eAm �7Js�W�W�x�����S�`i09�M�Ӡ�FZ:���<�TaN�R��eº�k9\7M���Mg�7z2��وճ�i���*��Y��h�]�r��T\�D�>K^A�H�:
��ȣ�h���6,���r�pL!�Ȫք
>S��u��1S��X�!��W{�$�|\�C3q��`�/�.
��㦰�%|{�:�t�ԡr�`�X6�����L�ȇ�K�\jP'+5�������T��K:�V.����J�j�}v�ZGV2ݚ]2���V#ïv�j]ۣF�z����$ݹ��.��P�n2�!�em�=n�pZ�TϏCmE�f�ێ#[WX��ʒ�iAKj�;t�H�
���_m��4�s�n˾n���y��7P3g5i���Y{���R�е��Qu�<�R۬���e�7���M�9�W��E|�]�ło���WQj������ې�RPΩ�\�.�+d��i���1�6	gw�"_*��M4{ �ee��U�Tęz��C�ip����}J�VtNcn�]�n��\z������2a;��4��̜�uMү.bs7tXD�e����X��vՕ�F�ņ�^h+1��[O�wV��/q�e�v/�Λ�ĥ,��m�G�:T�zF3�{'m� č���&R�pX6b�����T����<K2S	`�lE�W�ێ�F�^%��V���	��ա][��b��;��`UV
[�K�z�͢���u3��"�(K&jW�+o��F����E�_Oa��$VNB�9�+���!D�̨1��������+bb�i�W�;����'{�PU�٭����.�' �pKԶ�tJ���)���CH��N��`���5�a6�ۃ�ݡ�><ڰLI�Wj�u��.+����Jޥ�	Mr瑮�7�u��ʎN+0���_}��_W�|��gJ����8�j��ގ��C�� \��f�A�j��-W���t��}���Z3u9��R��{�o/�����V^e��l�x�E�⇆ar��hƳ�𔢯Q�q�X]��[#!��p��\��Wn�02j^&��c;U,}N��_�q��:=���O:te���}*���}t�reF9Z��p�I�H�
]� g��ט�ad�D�3��Jf��V�S^��v�C�<�����µ�����^G�]A�L��t)�ʥ)�c'E��;��A�tn�����[ehy]���H��ٻ=ʶ��S���P���S�ˀm�<�(<Ud8é�[Ep5!���ћ�8lN�)b�S�*���g.5|�	��t���P�
T��D+Z%"�9����xo3��9=�6
z����A8�Մ�2Phs�M����f�7Z�r8��KΜn��b�[�ӣuԀݤ�q�U�o�a�wB�z�zmEwj��:㬍��r@ǜ�i����z`u��hku��:��f@뺕<���5Y�֎Y�:JKz�n�����P�j��mF6�ZB��]�:�S�V/i�v+ �O+hM	q�c�o�F��ʽ����%GY��n5L1K
�f�Y]���<jظ�3�.cX��S�1���|
ܝ�N7k�==�l̈r� �94���9�L0�`Ƿ>�B�Qh3!ۻtr�C�21j_b�
����DG.̖EGT�����(��2*�'*)�G"�Q+@�"�T\*E(�Zir�.E�-�(�DQkH�"���r$�Tr��EQȢ�+�*Ď\�*�����ª��d	T�+0��G&E3�ͣ�*d%"��T�ETU�+��"�D$��BETTUs�U�(�9�"�"%B����
,�TE�IW*�H�W+�!s�՘�G)�Ҭ��"��ʢ�$�G,��"�.DG*"���I5D�p�QI%r��2���d�&r�ʹAJ!]�¹�Q]6\�8p�Eʀ�QDI��@Eʡ!#�Uː�*� �������QQA&��*L��˕2Lj�����������T*���Qt�����sP��
���Q@p�	R��UTp��?}�#�[ܗMeX�v<��D�|�sR��g]K�u,��lv(V�U�o�X�=�^r�mڜ���y��\R}�!�W�S��+����G�i�0��P�j�8�p��.�����W:2Y�z�AoP�L�g��[3��y0�|:��^P?Dr�^���H�-�ϡUp�/��ؠJ�AǞ����z�F}��#ac���i�K,�
�Q��X��Ns~9h�Gw�
���]Xe�3y��ǟJ�BN+g�'�Du��#eh�2�!�F�@�z��u�w�xZUY� p�1��3y�l9اk!�lS�`�w��`�(G^Up�B&wk�OL�w-�\���9.VP�����ɀ1]*d�b��W��v�;j��	�88)�p�4k���F!���w5���@=�}J�T:<���t�x��D[r.�O(�na^=,t��c���N���*BB���m�1�$�ڤg�<��kн5(t�ͩ����졖�:���۱��%��m����oDd��FLp�+��w2�򾹁�:۫�K[+DO�?NR F�k[=�zY��=A
���u�Wlw�G^I4�Oxک��t��w�v��7\��d=�i7�t��vk;Ӧ�Dj�4� �ȕe%���t�xc��2��ƽ��j�0�vq�~3� �/���ܸ�ї��9���扜���Qq)�f�ݍ����e��cɫx�y��B�pB���ngCurPngU�$��&�&]^�s��6;��ӓ;9	să@h(km��¿�n�`L���Ct��}ϊ���#^�FUK��i}�YQ{��mg����l7d���E�D����%�mp�m[s�UlI��w5�EE7f��2�MF��;)&�N���#!��`qȨx��iҾ��t�x�ޙp��U��D�����W�	�o�.Sq�U��������F^f��K˰s���s|�qq?/�������;��<u��C��,���ھ��.Ξy�x�1��+�8�`P-��/a���# �uN�1�.tL����.���Y3��R��Ed�C+��3���
y�F��Ďn���V�12zr��uӁ�',l�4N�b�&����|doR���d���>�O��7����_��n�3�[��[.V��=����T��=Ɩ�e�ҁ�F\v�I^�c��Ks��d��[G*0y�&;i펄ڞJA��^]NC��iU0�>��V����&ePU�5�j%���S�_#Nv�����X2�C��b�橢n0�\�'\�)s|�X�яfZ̧�ԫ�n8O;6: Q���w;���'�cH2����E�nT�9I@�G�K�V2͹�EKvQ���[���;j�?&OQ1u�*
�5�ȕ�K�����Y�R�
�_���o��6��Y����3�,�9���2 �D42S�U��'&�92�BZq֚,�2' gi��z���{�͸�G+Ҥş[�"C��5-��f���p���ڹ�]��G\Ї�.��O+r1�KFCt�[�|s�©�(��,����F�����'Ozli�0����ۦ���]���.��,imd3����&����K)<���Y��Y@b�f% '#����e�<��Lܪr{��hF��"A�����s!|./9��K����<�J�g��0jP�2b'A�t����\�A��dt�ЬY=�b���z�n��sڏUyMC��I21y|֣P��u"+a}�?��5�T��{��Ot�����U�6�Cn�e�ف_*�.� P<X��ˌ��V�>�̽����HI�%)��G���0�V�=�^���#+�+�O]x5$
�#��s��%*��59&wD6i��]�y�d]�I<1:�琅���S�@\��|����Vz�>���Z�]�2&�:�7���WSN�Xm3C�
�^��6�#�'Pi�37=D핀ߘB�n�9���S��1U��.�֘����\@u[���V���^��O�ơ��m��e�.o��;J�+D����ʻ=��*GpE�>��p��N�I�&���3Mg֖W�y�s�]@�����K�S��2c'꓊��7-����s{��$��B|�b�������9)L3�����BWnc5;�)uV�3n�ţ�{��;ө>�1��xtj½�_	r,��)�;[3��#�]�������Yd��S�����yt"�ޏmr��z���`���L
���je��C.ѕV���lC��s�[��
��8�k>9]��6nGZ\2��Q���|}0#^fF���P�ۖ�GS�Y�b�*,9n׌��oOg3S�x~���1��[�V����y��R����Ck.إ~�3��V�O;�f�[.��|�&�n̵���7�Qn&�f{	Q�nV�"f���QQ�"d;A��uQ˱S��ѕ�5u�	{;u�ԇ����Q�_�4�֮ܵFW�ǀh�*��TKgu��0f�W�
��WN���V��B�jH��f�����yamLϦ|�����/�.�+>F�3~�4&j	9v�P��<c�n��H{�[$��By�-�z�T��or�eM1j��m�k0�L+����=���[~�n�CM����f�:����it�ϣʊf�N,��ݩ�Eq��^)���M��wR�f�.�^�s�����R�F>Q>�fN�r�<����t5N�=�fL\����Q��uP���n��������|S�HK�DC�!R�:��=�*�;�uV�v�iJ�w�S���fN���b6F�46!�F�6�+]S*PB���N\�Nn)�SZ� Nk��hK��j�!b�sЃ��O��#�T�Κ���"u����*���)���gmͫ��w_v�x���}aL4���m�����y�+��`���V�nC��`�׵/i%�V��w*��U\t�`���4~�� �W��ӊ�����[�qT'�F�Ƙy�[x�2�]���F��~��!�����t��g�@����W�] �(��!]�O���d�Ԅd���o%�w�߰/�7�=�+ULƾ���Rs���\V[�F.q���=r-%�+4
	�işg�T=���^1?nъ�Q��.���
�ÆI��G_un�f�+R��wN��4�p������}N�C�ߩְu����B3��7������.9����'rR@�@����7�\�<+D>�X�ش�}!�c���x+�F����[�ܒ�h�E��1�6'>�H�>��L�eughw� ���/#Du��{I�u��uV%��˃d���vܬ����^�Z���&���&�/��g�4ǰ�,�U�\�H-T:��n�m�4u��2�����R5\�z;�Rˈ����?Z��T:<���o��#c�B��b��3=
@^�3�^��]��-�ق�ٗ$e|v�:2�J�;���G���!���Ô��eO=�qF��p9�+rd&#"��'k^�`�4��I�Ip
����iq�E��bu����9cĊ�0(>75m�dϼ���2���gT4�3�-t$���`��9���8��b���%�~��z���SL䥮��c�P�s87���I�^��v7���V �¦G�A�'�MV���1.vd˦����뎽��O*�;y-�dX��~�ػJ����8*��n&�ѱ�*���)��d��W��	��جQdw\�&^���x��y���%}3�=Y1,A�� `u	�]n�A�HԳ�6ʛ�*V�`�q�&��<D��q@?�Vdy⼒�p�Ĝ˒n:XD$�Y��s�ǰ���ڦԶB�u�׸u���Of��+���@�@�($�g���dՒUj�:�PS;#��z�{�0��ɖq�f���%I�v'�y=�^(����d��NF�tF�F�q�9�����Vߴe����"���; `^�e3��h��V	��\����-#�	ȶ(������E��g`�h	�i�X1nr$n�A�(ɿ}��Z⽺���G{R�MnK������ t��nBߊy�G1�c�;>o;�V�"&J{��11r���ŗ�i��)w������
Z��2\�O�'rD.u��;ɹ�O`#|9Y�{�S��Ϸ�p�3�g�ʍC�`)��{��g;�9�ֱZݖ#bf�jm���ж󸤱(��Z��ƻh\>'0�#�}��`uE.�3(*�����U+��XMR����i>,U�U���{�A2,F�>&�K����>�v�����机ȾTxk�mR%@��N"F����=�>r�2#{�����$֓��-g+��J��	ә��U��J�WT3�sB.;�g��܌��KF7I��[y�GL.�	���X-k�HZ��3.*��wn�ŕ5h�s�3.��è�:ᵐ���c긮;s@q�6�.qܕd����t�	R��O[���� b�9�Ȇ�����Ovv[�&.��w!c�ʆ�z2���\����Å?օ�$��P����r/>v�Ȱ�z
�85َ���&)`�W�r�z`�6n֩h�1a2k紸`6���XL�Q9�4�Kf�6VY.2�=��ހ"��و�{G���y�N���;\�0v�'�+v!s����sdܮ�9Y9�������,ٳ]A]�QK\�a��"#� �ܗ5wǍ����W��2�ת����$Ș^_&�QzKg�Y�7���2`Ǟ���'�p/���ê���:����3��f}
��*[.����UYPy�z���m�k�!G�t��&2'���H㡍�r�+���x=��J�sl2�#�'���@���f�{_�\��hA�`R�A!h0��/ 2.�$����#�BOE���z��G�-E��Mh�p�U|���5;n�؅uʏw�5�n��<G��޿ L�j�j!�)�~|v�E¦�چr&�?e����y:�����I��@6x_^�~Þ=m�="�7X�2�];���+���"ϸ/��wN֫�0R��rW�~��=�i�=�$�V�P�:5"3�\�>�*�	�4�h��g���h��:��-��D��z<x *����=��Ya��#X8�ώ|FL^ٲ�h܊�:;NaLu�qt��+}h�5�:�aN7,֎�2�z��\%E�#bݦ�tf7��B2#��I�=W���xH���u�-T�Xh�0e1���W����Ǿ�>��t��C�	rc��ee�����#��a��.ȯ�-#~�����S�9z�H:q�y|�Ww
X�Z��i�*\�q�{�xq�kQD��
m;�{}�yKcUNB�"e���EI��+Ec�����4�S���q졾v;(s��ml�s�t�;n̵9��M��A�W}�*��hC�D\��t�ؑԥ]Q#"n���6s&6�e|��9��O�+fڋC�߭�	��O~�;W���'��� 蟠��!��D�v}�w�%��5�� D
�%^�a�h�2�� �����>ؐ�����Y2�ߩ�ׄgH'�OR8EZi9���Z�|P�gp5��^
`�������	�p��N�4���*P��y��E�x�u���wn��ZF�/���3cH0�ْ��b��hl:�ً��q]�튛UA	E�܂*7�9y�cuBG��;��fW��S�����ir�b5����:�Y��Tڸ���(�D���$���J�ɪ���C�������R��V	r����V�b$r�N)��X���]�JF���dV ��DR�|N�#����鮎A�[ͧuѪ��^��=L]0��'&���n��e��p�LɖÙ��By8��ˏd#�D6��[����)z���[9c6�S��[)50������'�Y ���1���P"Ii�.�ɸ�Ҳ6Ծ��e^�$�Է��$îCbB]����U�yԀ�bH���o�J�]]�FCur����dD:�ӴJ���3XyN��zCm^*[}*�;JU;.�L,��g��F�c�˱z{R�5 F�	_.���G<���<��,-*�2��-�4��8��
�脜V�Qy�DuÀ�
V?A�S��݌�^�C\�W�ia���*���M9���7�֦o9��;�;Ycb�k~n�x�xP�RQy���;�kڝ=Ϻc���42�P�C��N��Q|��8	������;L�����DtT����6�p����M_��S���mR���<���`H��<��P�,�ۢ�W'C�=ǣ�{���qp��^pxL���6�uk�iQ'x�%�����*#Hp�o�9N7a!�*o��x��9H�S��#�
��\{n���:�윭]p���6�ZU,�.�"r
�0�����M#�+Ղ2Yʁ�˚�ߑX��j����<��@��f�����������L�*QRze˥���t��uV0^;��ӓ;8�<Hw�P��}��S	w�L���K>��7/x�� z�$b�-Wrf-s�&w�mg�s��0ݒ�}��nz���.�F�L�g��E�w���ѫ�@�f�s)B:��5����PSWMS�s��t���f#�t�ŀ_gUstvy�(��)��5�e�Ey<ͿlN��+��ƥ�f'�&��
 ��Ѯ�Օ�h���Û`_>���(s���8�[�X�]��{��Oz�]���C�B{	5*n���;[�WL:�S�%,�EDM}��.H.řB�fu]��i�6�0ⲉ��sGT����{v|����׾�aR+#�H��wz���B�jo�}�y�@���^�9M9�±�R�m��}o\��.��e<	.3U�w�[��&M�`�.��89j��/n��Ph�A���[��V5.ݏ�d�ʣ�(���l�`c��sa�1�nV��)�.�ᗨ��	h�8�2DNo�w,WSq���F�f3a�1����B��ǆ��x�w[����C���7�5<K���N��ݵ+u��/��t��B\���AƷ_(�S���Ib�cI��kye^f�C^��3���(S�8+��**�� �^Z7�i.5��tv�>x��$���J<%��� �z��zҌ>�NP�`/��n�=C�YD�h���s����t8�Hr�2��N��Kz*G>`�@I����9,W�U1W�l���I�������nr��ic�7�uMҭ���/N���*�1�;�|D���L��h��WÇd0�zh�_mnڇ������r�Lv*�>�׆[͕	�tӽ����B��ݺ�[��J�S���E+�R���]=��[�ڻ̭�����;�	9ko��ղ%M<�A�2�u��S�ۭ�M�5;�롉yQ&b�B%��[�����N���#i>�d�$W��_�oɶ��"�߭�nT�EX�ѵk���9=tO*���q��b ��U�g�=)�'{�W�K�5�b��˛k�|�Fu�T2hT����%b7{6X���q�X�)��8��p��Ͱ{������Q�S�����̅V�ss7�
�|�N7f"����SL�'B[0�!����v����mI\���'��#��oa�)P��W��J�ų�A�����bv�<���W;i55iuZ�3d`��fs���WK~���d#�]k�%�����kon��U|p-Hl� t�H��Xwr�}6=�h8��[R��1�5��˹j�%�]�5�0m=�]�j&��;�������YRjxw �cSUj�ZyʅQ�kvF��'�V�&u��M��6����f����=��)�Wl���N���*��V�.�eaYp0����/h���ܽ&X�����Pݿ�*��
�a���A|H
�뢫�t	`t*k��R�B"
���\�E����76oqȆ�fڻ��|��Æ:�v<�g^����mm�I��N��)tȧ!�ไI�A])���7/M;y|&h�Ϣ��pˬ�_!�5˪-]l � �(#�r��2B48EDZ��0
(��g*�E�1kC�̒*�+��*.�(�p�8EEQQ�$8AF�*$����-0�AȊ��TE9Qʨ� ��Fl�(�(�"9��H�"*��G
���Ȋ��I(�qZQ*UQr��jG"*
�ª����(����s�G�Ar""�QG9I2�,�DQˑ+J*�r���W("8�8E\���QFl�˕Qȃ�r�D&Q\��Q�fr.TW9TVTUȹQȈ���"
���UL.Z,
�QDTAjr"0�9ʪ
*M��\"dY�Rt��Φ
�ʨ�³�E�����p�
��eʹJ�JҢ"��EdI""��ȊI9TQZ�9˲�2
.\9��*��V*(��PQr"(��8Dr(*�EDrԈ�$���p��r"�Qh
={��ٯ��tVD�(����sy{й�l&�-w�Na�wy�d�=�o���F�,gY���'ɦ3m��!�[.I /�S���
����L*�X�(I�M�
�];��?�:~�q8�^��������C��7J���c}���;~�~����@��y��Ƿx�!��~<|�G�<����_k�Z*�`��) +�O�V���v�s�}����[������]�N7���%p)��?�G�n���ל>��=M�q7���ӼOq?!ۿ�<��®�4���ۯ�~�ݙ�����?�LF�}DG�ˏ�|N;q۽��;w�k��7���i�Bt�~���
o�$�אv��n��C���@��������'��w��t��G/�v��k����{V�+���W~�>�T��*���V?T�N���q��=�}C�aW{���Bp~��:�7�q8����������Oϯ���7i�Bv����-��M�u��0�q��t��_�� ~Hq��=�x���+�⽣q�G���l�'�?|&>����o�����7���M�v���ͧz������[�>&x����|!���}���QC��w=��{l�w��{�����q��?\w�m��o�8�^����Y�瞂��DT����DxSra�8�GJ��i�w�?;<w󴟻��:~�q8�}7��c��!>�|���9�1;�k�������&o�{��ѿ<r����x��M~�����{�>|���(��.*�r����}�5��j|q�t��qF�N8�}C�Ü�
��W��q0�;��/��ۈw�p<I���-����7�N�������$�����7�q�'\���77sK�T��~-A��}�9��*j~��|�;�i7��N{�α��j�]���O��&�F�~��x��>������C��{܏]��wa�|C���I��\���N?�]q@�'�c�͙��.�r9$R�ޣ��S^3��7������|��8�������u��:�;v��!>��}wn��8�_���ۧq]��8��q�o�_�ëN�7��vr:w��0��n����o�H}UwO>9%��?~��gwF@�@UD�C�����eӼ}��F�]��v���n���n{��y�0�z�y�~C���;�v���;t|��I�ۧ��v���x����&������ۘo!V��f�C����QOc��+�aܭ�BP��r�ZQ�o6<X�6tmƶ�F�([53��K��Bo��R���F9Bs����9&-<-Xدq7Y��(R=As�/�N>[�j�ˣ)���9ڹ,����ѕ��3`}�/79��6���*q�N�ǽ�][>'I��{��Ѻx��}��t�Sx{��޻\�{�다��������N�=q��?�~�������/�P��}�L�O��*����r����n���_����;��r���]� �C�����o��{�n?�}���n'_���� �}�$�7���yP���:<��o���������>�N��WsC�?9��q0��HI��!ﱹ�n!����� z���W8~;q7�� 8�v��q���>!�a����{�ޏ�~v�;K��t��i�|���~�x�'��d	�3���cMj5莘���5&�������N�o�~�ۼN��~P|N�q�&PPP�?;���a��t�r��7o�n'hӿ{m�#|s������~}��~C�a�;���p�>����5�n~ا�R���� }������o��?;z��\}����	����xc����'�lv���ӻ<������ v~�:v��<r�Q봘P�r<�����o�y���'�OS}_��x	^���P�ބ���Q��&~ٌ�����?t�;Ǿ�ѻ|q�v�=뛯�I���۟ǽt�����#���o��!:O����1&�x�N;q瑿!���v����$�t�&�_=�׫L���d�I��^�����~��vs��S�q�����`��!븇�}��I����;<��[�wHq��=��&����$���u��8�}O�9�v��'w��I��ۉ��ߜ1�v��p�ܳ�{�#c�>i�~����`��[�����<�ߝ;�i��9�z�������ۤ�;���<��A�#�M�s��q�n�8�^��=O�8��y���S��9��a��S�����*��q�{�I�;��� ��`����������!�����o�q0�׽��W;N���1�v��}x���,)�B��y��G��'���m�>u���޶�m��t��ϟ~s�y��#���;����'p_����k�=?~�N�v������;\���7N�8���u��&x��|.�}C�L)��=M����8�ݎy�}O�?o��|@�'}v����v�oP���o+;���r`���i8͊����%�#=n^Y\m���X@��T��ך��2{+l���wHD�b�����N�L���$�<��������O���O�yu�$�����
�Uۣ5�"�]s�9ܗ�j��N���ʕ4�ӝA-��ūR���O�1���\FI;z��'�׼'|v�8�x��p��i���|N�t�W�I�N'�����1;���'�>�I��?�v�wn��!�k�q\!&���?���y�Ϫ�4�O���LELz<v�?}�$��uκĞ���M���;L+�������_S�?�㾻I������t�;�&������	7���7#�:��N���>w���}�v�߲��=~��}�����U6>��B�}V<C����һ(����:?!�0�m�9�ӿ>������0���n~�}��;L*�S��y�����>q�ۈ!��j]U~��}�>K�Z�w�2���������߯��o���O�=(�:W����t�v�9���;��u���t�����x�Q�~_{�.��T��&��w��#���ۼO\q<w\����t�~��`�C����&������4� U߷ߟ��������~M<q���[?�I���;9c�w��s�}v�oP���N�{Nݟ{���v�瑿���A۾;H?��z���t�=���I�v������&�=N!��w��~�{�<��?0���{�@���tǨ\�t���
w���v��qۉ\HI���,�#z�:����۴wø��I�����v�
�������	��P?z���?��?.�Q�B�}[�y~���~����E]���!���E}b����|��|W��}x����:����X�����v�~��'q���®�)�Q�~C�����Ӽ|k�8}������~�~�c�e��|����ܿt{�W�*�W� ����!��������\|~���'��^?=���i�B~����j�Sy�ݸ��`��ӧj����'}@q�;Tx��޻J�����������E@���/�yə��+��Uc�|���''�Ow�=��'�����s�z�����θt��4�q�{�s�I��~��޶���N�w�`�x���'��q��8��
I����y�ϟϓ��ڙ�?��l���U!�|E|�1���߫��'��J�y� �����w����щߐ�<�޷�=C��a�y����t�]�Oy�q�	��}�v�z��>��v�������׼\�� ��ּ�8��}*�z�.�]XJ�)Lnj(��[i��t�{��R�;q�F�9O�w[�,���X�n�q�)Ɠ�iFC�]]�d�R��-#S+$��7z��cJpM�]a��Zwg:�[�+[7�S��v}U;��y��vs�}Z>�)��w�<�ht�W���:M�$�Q�o]�'N��wm�t;z����n&��oOz�֕���w~y����B�1'�=랦����8�N����K�|'25�h��"=�H}�D���G�����V�yӾ�&����N��{c�~�����8}v���w���~v⻧}�����'��=��_�i7�O��m�q\
�Vג��v^a�U��H#����;?}SG�{��7N�ڭ�>�۾rL.�v���^ܻ�ҡ���y�8�.���}q��p�7�v�]�u��;O�}C�>�c��SO���v�|�L����#��C;
�v.(�9�예S~���:ۿ��ۉ�o�{�N��i��y�oP�v�����sP���>Pz�<p�]!��M�q8��ڸ�7��8�����|�N��'���'��>=Pf2�n��$�) ��?)�3�O�~���F:WP��ϼ��0�����|~�q�����I�ӷ��HI�~[��8��7�$�P����N��4�$;}t����I�B�?u���z2��ѥ�p�~��뙟�&c�E���o�_я{��ߞ8㾧����y?G�*~�YNb2~��T�=�2!�E�� ,���
b�X������*i����?A�VN'qS�}JX�/��iU�C��\9��!���0��-�����l�^��C��*�!^��v�/�0p9�#��� =��^k��m-������3�z���K W�.����g)l�$��ހu�yΞ廵��(̌�. �4�ۧ0U;2��,Mig�8v�� ���F��br�\��:5I�P$�_�OU�V��S]I`�q[�ii�M��C�2Fr�@1˹@��M18�r����`Ve���&͹��E=��֚q���_�Gtj,�yVs%��KK�]�Nǜ��=�;�����Z�$�V(��PK��Q)/�D}	�	m��`��=˳!�IV�lD�×��>�L@j�����@�53%g�w K��m�<���S��fB�4F���@b�����+P��=A
�Y^��;�Ae�;|�g®������ʐx�^;�`�L}���Xv��0�ɝ��.x��j��5���<��aj��A�����¢$o���ZP��{c���9�tGMM�V�TW��H������}���Jy����uDp�8r����A��	h�
�V�u��yi%���n��#>b6X۾��z�*�x��|�Pl�b^ר�6��\7n�*�tv�}�	T��n;�`6��}�� ���X�o�N��~T�F/�RU�՗��~���^>ŎӬ���$�>�Չ�T�u3�CspD`����!J�,�p1,&�i(�T+�4z���}���E�T{�S��=�Do:��c�;���=՝�ĵeZ+��;��>F���ۨ�]p�k�xe<W�F�R�h\�p����rw$B˺�y�V@M3�x�W�K e*�rD[�-d��>>�-K��0��]�}�\
�w�|�	�"b�2��F�Oa��.ۺN�z/]?d���$� ��vL;n����j��h�H<��E;0jf�3ޠQ}5���r�+�BXj*��6 �id+��'����^�mkEE��~�sg'>y�Z3����f�a�b2��J���C���"�.��Ձ�k(��VX��N1*{OŔr���$UC+��v|��X쌹�Y�n��VSw �����m�zQ� L�j2}F
خIhS�E�ms��N��0a=g
�Qb*@C���gO騫!h}�����VHr��J�����'p{����-���Ź<2������#^�!'��d�]/���ϗ;�g��܌�Q,=�&�y���!��]�A�d�nV6��ӳ��BBeh8W���ʙ�q���0�O_��T̻S�D����f��\�mC�F<Q�$�y���E�+W����-)Gp*��R�z}��@�#�c�l��:{����[]����`����\,��\��&)��B���uk�✕���]`g�d~���Tw!�~�c>�'���	���#_���rG��Ɛ���{�H�r�s���a|�=�Y���&8�|f��I�C~�U���]{#>m�u傊��B=�K���hdla�R={qKq�)�%���w`xu50I�wJrc[J0kk$- LM�補��o>�pTaL�w.�;���*��Pg�p���u�6�w	Qc� J{�b����ި��۩�q'�
\$����1A�i��H�_��"" ��6�tT�L�B�<�=�I��D�p��A�\�U��!}3r�7V)��LC_�=�@yf'm���2�>�w[���Q�,:�F������2�2.�ZIࡉ�G8���rF˾���]� *84tP� �ӵ�D�)Vv�v����]s�������/���_8}���
PZڱ;T�s _�����h��U���?5�c<+�>�~�W�&���};^lr`�xz�����x�yR0����:��F&���d@�Y��2~�j\Nwh�iF��ZOR8c>�Z�ê͏q;U&}ڥ6�ۇ����U�l�a	::�������$�KJ�͛v��υ�`!��"�����Ya��#X9���ZA���b���-����qJt��q5_;�v6pZ�f�R�Y�a Xr[��غ3�E9�,��)c�K2���Z,>¤ex[i�t�𧯘����V�<���l�s l�K3+�4�t����Z���ZD\#�Hf��&*�*>�����.�N�����|߀�1^��׻<��X}ڲm"���A����|)�i��.�� �B�+E{�[̡�d�ʀ����T^�v)R���	ܪR��uѫ�[���U��a�N���;�'�X��F�\��(%DK��V�(%�<u6�t��Λ��i��uh��_U}�Ո��&移r��B�ϟX����A���1`� ����
��${B�b �gBK^��OEXsz��t���j�ϨK�_��M��LT@D�G�� g��`+�v�_%ǒV�)���}y<F�k"�0H�UOn�������)
�UR&��-Ҋ�	�|��e���ؚ�o鿸QALl!E�6d�v؇�Hަ�ê���m�W140��I�Yu�Z��ގ��۳��(BM�W��?��3�1r�Ӟ�T�g��8�Næ�1ڪDf�Ʌkf���d���3B��^q�u
�v�	Ay4tE��B�)�M�y��.M�3��Q�{sZ�Ō������r[�B�Ja��Q1��'�ʊ�}[�{*�FW+8���#Fv��r2a�Ӹ�bW�249�smә�����z>��0��p���I4��<�5fk���ee2UGNu�$�އ��ˠ�7�=�+_A�1�u��,�¨���o
B-���z.olw�_y�|25Н3�4��j�!T=�8�aqy�G\o-�3{׼��]f�Z@����g�@��ez���8h-����g}|5Jnɹ���^�ы�Z�d��v��]�I��r�|�a����y�B�ʈu��Ȝx�<���7�C�K�C�bՎ�)GZ�2m��Ί��r�bP�#��X�x���mj�"�����3^C[X�Ψ(|NM\��vW�i��s�c��ˡFcJ�"lvV��]�E����b2;6�D!;�*�Mz����/�����|P;�n�eb>�"F\^���r����i�tx���a����>&M�h�����,��f$U���+�Ǳ�ů�1��r����(�~ž�6��ºל?��hc<I�$��+�6��D����°3Z�=���GD��d(.��=0��|�!x��|��'+W_Ȱ��4�q��QP5�]N�s%��G(̸�n;.��S��Z
nj�Ec#a�2#��zr��Ǐ�;����R]�6U  �:�OcWq��[��_���xA�-v�_5C��ؾh��uo+��hf���
�A��� H� ��i!֥=�v��)�o�g���s|�u��xv�sPY�]�hd�l�1�Ȣ 1�%}���I���f�Z�=�\]o~�Nwii;�ϊ�g���,S���#>b6X�n�g�����CGP��]nð+,���^�߹`Է�֭4��@�����G��k�G���3&�kOC�2�JH�8�y��z�Oe�a�t.�	�/��Y��{���6"�[����fQ��L�6m,,�������E=��րًpr\�����h�H7u6[�uw7�c�8E�2?}U�}Gm>N�k�!Ctm���K*j7�
�`_ͻ2�1nfL���UJ�H��F'7���s�Y�j���X~p�7�.Rc �DbO��MX��I�Cw2^�w7���M4�͍�㧏+I��U+L�Q��YA����}����T{�`��Do:��x�Ď�f	y�r��pR. �´c2j'*�*a���{1\��a��g�V�ߐ�ȴt0g'I.��"n����nuf�h�@f#�t#0�u1�*�Fv�I.���m�q�oj�kz�$����ՄSn���6�u=��_2�Z[�������j++g���f��n��%�����Oz�� ]W��Hڷu!;F
دd��_�\�b4����.�2�Xug���o����Y���U�����@�q+$9`_�Qa��y󕁑��3Q�YCg����cZ���KGY�M��l��T��]R5q\Ћ\���܆"XxI_ݻٰ�e��Q��V3���45��t��4��yCA��7�*Yp�b�x��f]�������l��Z�����V��L�p[�w�r�3�B��B���n��&��g����Vu���C�������֋����	�v�]�V/w*�	Q ݡ}4k��@����V�ɱ���2�smlo9���	������W@�Z�[���%�س&�f*�r��X�m�Ә)J�6�lkn����]�| �j$.��)凭_�C�����N7
���i�A�r�Y�QލU2��>q;���Ӭ2SQV+�k�m��vm�z�vQ�'_6[9X��*��OdF��Vs�f$���6�5.���f�X�V�	H �<�s���X�Y�L�qY��Gu]ؔI]!��t�i�S͛�I4fX��eN�9��i������*i�P��d)�[���ol�Z��30���%���W;(��G��T���[��s�H�S��n���J,]aFCt�gwv�]�����=1m�Wm������CYZ9�)뻭���ܷR��V���/(��ړ�+f����	�@Sb�bNܱ��JG�`&����%=�k/2��w9EZ��:��+��Q
��\kk�;��LX����Q�ۊ#�umN��a}��P�1p���C9�i=��z�{Z,D/�.��&I�_Ln-���t��\X�x���[�n\�LR̎�����mv)u�+8I�Ytu�U�����@��!�k�Ǖ�n�u�G��m=.�<S��R�}�gq�l���.]+Nw��^l�,���j�j�h�T��uy���}Z��׶�Kz	[�����wf�N���/2��Z��}�e��KBC@��8i��XIԊ4�l����$��N�(h%��o��h[O{�>SM�Q�Mˮ��H򭤔ׂ��R�X��ش_R�U����I��v�"V���[��N�d����mKD�΂�16]�n��J��40�
��wW��R£��At}5��x�,�v	���_D�,:Y���e��5PX�]���rM���4*uޓ̉��m�	�LHYV���WV͂��ob�GkT��W�[9-�œ���P���wx �.��̴�`l�,���(Sk�)�}{5\�8zREl��
��dZp�'>�F@����A���O;E_L����y[�(\V���aW*���Z&���`�f�š{ϥn���"�Z��r�rU����x[���&)M��M?�]WN�b}�}���r��z��gC�T�U] �ĥ�����/皶]�³�E�p����B�Ӈ"�Z�ģ(�������d2M}%��2F��ܭb�T�ڃGs�tel*e�K��V�;��w)}�Fy�R*:�uw�]F(p߂Ƿf�&������y��l���'flo�s���Z��Ѵ�7,Wor;h�6`�I���S���VE��v���qZ8su:�>���ΗvY����6��]��i5��m�.D��k!��e���6����'G�>\5|;r��Ym�$���&�A�6�����P 
� >���Up��+0(�*"(��\((+�����QDDr�F�QR�f\�EE\(��PQd,9I!�Ν �����9�Q
�&�(�*�QQ�J
):���Qp����D�TZ�9PQDDA�"#���Y$��#�ʠ��ȹ�E�0��PG.S":��( �(��ra��\�eQ\ �T\((�*�j�
**9Tr ��"9Ep�QP��Er�QE'iPU�p��	6W$��WU4�� �ATEW(��ITYШ�W
(L"�QQ¹]�(��"*�raL�TADEZ��ʊ���ETA�]3�	�r	j�AE2Μ��+��}�ɓɧ70-�`��VM��j�'A�b�r�)2nZ�b��BB�V�U:Q���3Q\,�7wg�OJ�XZ%~��"">CN��""H?��C:+P��$̢�����3�R�����Y#$5ܝ{���IL���ݮ"��^U���κţ����]A|y_�$����o����ݼ{�G7YH?������Z=�,~�w�|!7��Q���O�<� 4�<��[Y'tQ���!��1�.3_rN����dco�06P���[�'M�]}�����-ȏ����YO.1��&��Dm�	t1��0�V��8��h&��W�齂{�I|�!��#z6�]:�57��M.��/"�Q��!�ĀE)h�Vo�v��N�
��
����(�U���/��>�Mtu��-[�{�
z�ϔ��Ħ�&EeN�f��|�*��$�[t�@��g��R/��i�y]��$�ca}�:����	�e��i0�ڲ�l�HH��1x�4߅_��c�v/O�i�������ڢ�T�g8��P���,�<��Zq�����_8�z��/��~���Њ��G���P�~���+��/��T�N�Bу���ntgz쫒7��x§��ٸ�wj��q	R"�m���(�[$�Osh˗�I�.��|�/��\$rs�́n�Z}���´���ڱs�B�A\�\��"sz�)����`m$q�*G�n�G�����_�">�����	o�ҫ�'B����49 G�TEg!�R�,0;�����.����6��������7�i�K�?�_GIy�_1膞�k�
t���i�b;6U��y���	���=L�
*�W�7��h`�|)}��r�؉�y+by��+���oS�kK����ٝݘd�`�2���"-�C0��������Pl�-�\��KikOy)��0�ҊΖdC�O�K�o>|\D���rq_p�u�/q.+��k�9Y���}�I�K�-̊#"m�}p�[��F���%�ϡ��w�`4 �ͥ]�\�F�gwq�{�8"��1hA!����65�r$UOn���z�X�)�+�qЉ���N;�&F�U�"`����6&���o�&ơB�Fx���b6F�47�U1t��t�m��݇��JA��j튛�UA������Q	蘿������^P}���;�	CF�u\�v�	e����đ�O_���r�p�Gn�U=t�O�tyWk��u#�����+��� (�t�ʐ�)��Gk]�_U�\w;[1Eas-V:o��h�����$��c6�\/X�:vp��/�� �è4�$��M��6u( Y����V-��2��ʌ���/K�3D��c<�a{�ζ�Ͱ{U�zY���������(s��`e��3�>�+`7!��Q&6f_�0�D����g�/�E����5��<�]T#gk��L8e�9�����^U�O����6�Z�.<����UK��>�2^W��=�{	���dW3٪��e��scrs��>r$7Ĭ�3.ܬ^v�w���DV����֭��t�q��F�Y�|C����|^d�YD}�S)0��Q�6��2FP���F��a���3�
�5����s�S����'oQQ�G:���\Fz��B}T�if�
��7p�A����<6_0<.�����Q �9/�].�h�."���C��W������ġc���q:+���S�g�,Ȧ�� J�ت�,�|�Ԗ��<+�����>���˫\I�D�ܔ�r�ؠ��]��L�51���kY�J��e�?Iv�o��^�ϲ�չ;[}'"�i<��ʃ�}-�H�N�Z�&�ٗ]�˪b��_�)��Ec#Z��-W��ٮqV�"f�T�'K<�z����tS���]ssp<��h���NҴ�L[Z@W@Sɼ�0f���˸�E��r/���l7�̧S�ޓ4t�w,�s�/z�Ɩ�w%Έ���y��դGQ�h�_���rFW��`��T�, �ua�+���������p\��(���@��a��
�?gˮ������t���B\�!H�daۜI�z��#_�!��:�0����Ѱ�DH�Wo��
u��4�V�j��m�\�j��Ɛ��@�}������+�E�:MZ�q��j��,e�:��%�������T�髷~���;���K�m�L�w�`}!⬄(�c6��zO �����m�oZϜ��ʛ�*��~mِ�ә��1�I�,�0��\��j���.���rZ������Lu���Dd$�>ϓWo&m��{]��f�nu�Ӧ��l�5P���P�3��1�c��L??���Yb_@~�MW:��Z)�g���B���>�sI`���D���!�´���L]p���GSو���p{JãÞ�8��I���zu-�d�m\�~��K�v�rgPp!�{,6+��+��Co�����R�׎ے�@	�PeʧZ�lCvX�.�w��7�����;��M<}3�:�u�|[�|�5�3ٳ5�y��M=��p�[��=��oe��iE�<E�m��a"��z�;=�=Ґ[�N���u���9Zo�b��r���5ս����-�[c���)&�q�O��ߩ���t�͕x�V�`�䦯%#��ﾊ���MaiV�h�&~^ >�V�$AY:ԓ����:FP���3�*Z�u�;�O;���Q	-t ���Ǚ���H_�_�M�\�.��=��+ 2#{ ��7�&�gJ��o{\�����=[�$��L
櫥��3Q�q\Ћ���QΜ��Xz2���z��ۻ��a�B}W�\rf�47�z�'��T��ڂZS�Q����q��L'�O_��p"ol~�l'��ճ"�u��C���Ί�>���@�c+�U@�HgUHn����q��yvQ����z�� t`��cg�hF�CA�Pdh�j�d�/���
&�	_�/��v7\����ҝ'��]����b�3>g"���9�Gt7|!7�TF�7�:�H�B �V�+;^;w�5�ST��?i�b��_��q�C�3Bޚ�|�����a����F6�̱��.��m3�_7e��tC9��!#���#�G�f�/�i�ۨ3q�k���i	����^�z�́�{��
�I&c�-�C#�Vi��Z��c����n��3K���Wv��eCt�9�7�{މ���=۞	O��w���²W�kj浉z��9���o���d�z�B���
W����Z����B�Ӆ��L�ש�0���X�mK>��軨޷�;�Ȓ�N]JF��Uլ��"��@:��*�gD���[�~����3��s:�4sq
�r�޿YO�^p�1������t����T�Y�����e�X>6�gb�����̩Ȕĺ���s \[?_������O��U^H>9�l6��S#��NqG"'�WOOo�/��~��1�)xX:_����)����D�3�+1m$N4�o�\[��@��t�l��UN-^�V/��~�
�r4&G��g>YP'��t:�����q��RRuG�lZb���
FÇl�v{�=Ҫ���m_ݣ!�uflr7����z�{��)��6�Ӱ�*����s��W ���)Io����l�Ӣ�u����8f��[�g3^�x~�Ѹ6�F˿
ϖL�٢�����kh�<����g�z�Æ�0iіP�"Lk��f��w��T|.�Rށp�(ǆQ�(����k.�"�e�3P�rX���φEet��2�
G�R��GoW�Sb���-ޜb�#ִ�<2&�W֩[ѭPb;!��|��U�� ��à+r^kk�ޥ
;v��|�-sMv�iLn����;ْ�љ��(�2����[m�/�P�
P_	Sa��q��ɷwAU�$���)�k�8َu�/z"�v�s����F������y���4��Jm�t	�gлޫ�N�c���i"j_���ꪭ��$��S����Y��wHV|�O�f�Ƭk"�0H@C����	���Nf@����
��b�z'�8��{�W�0��I_�q
aLi2U;lC����]�@i�;z%.�3��̃1�*Y��rG�#�V�6�����ν=9iџ��.jb�V���0�$��}s���M`c~�:�Y_�J��\J�@=��N�Eݮ��[���v�^ֿ-3����5S�zę0l}p���)��e
1)~�LG6��{*5#�u���[�.w��-Vo$ʃ=[�`�/q��j�hs2��s<�ד��}$0=ڱ���-aڲ��k��8z=��#�n3!UN]!��EM�ۨ�)��w��$��&/)iK�޾�³g���_�A^
��	X~��[���Bt�4��Ӌ>�
�茈I��:��w,F��Y��4����� �iFH����ύp��u�X�΂������:�kaȕ�# ���}k�2�M-��tk�}�f�����Z���چ���߅y�36��ɀxK�-�nr�d�C�����P
]!y�}E9^Խ�g�ᅑ%��S�cͽ�Jd�6�.ܤ2�O{K<�W罃�R����d�[L�A<$U�K;�ћ2�R�v�gku1F2[�x��讠,B�Y��TVQ�w����"��jSMO������i�ǋ{���;j�2��/G�G�Z}�]����53�v42�ǻ��U�=������ک��H�7d�jCT:��5F��p�����������[��;��%���Imo�¡�����|�]�ꭸIG����9�K�)HN��k>"��(dSv�P.��/>�L@j�����L����Zmh��9��0��ɯ|��&e��Q�t�T.SsW�dkTdpB���Y�Jn��RП���Z<N��q]^S Ҏ;��B�l���V���W�&vwxV�W.�G]w�N��y�4vg�����P��R2����?x�D�K��p��������n��,�����cx9����Q ��C!3���)Љ�{��>��UYx;���'~r'!��=R{�$�)�t��l�/����CבV 1�|��4���=ѽܸs�v�m�qI��ȇ��6���C*n;>*�m�2�� ����r+fØ��a��n���[����]⌟�l�)6m�/���gؚ�x�0(dCn�K���J�Q��<��ʳ��*a���Q��+k0�gV��Q]`�I��6��T����j�õ1:B�i����7�[�r�^qcjTA�S����0�L�D\�A�H�k5�6���"vq�d⮱k�dG�#���&�J���_m_,[w"��ح�+�DG�}�H�^X���i�$��N�qAO��c��~ϱ�߃ʡ/��(�J��Z(�_z�O�Qy�9���_`v���Q��6j����Z�w��^a٭\`����J������J��oJ�;+��C��H�ξ�?k͵k�L�
��$�����r���<�ӛ�zubb�t��=�t�j��O-�����J�Z�kvX��Nh���U�M��H�P�]�؆�N����v�Ҭ����T>��S%���q��F�rKB�z,ck���Y�����ѓ<�%�R��6K��C߭ݠlD4�q+"C�@��}�>r��ȍ��5��i�;��<P��b�H�/�� D˗�MWJ���8�hE��(�NAu������3ӐJ�ZJ��V��Z9��zO��|�%�(򆃧�ofT��r�;�yW�m�k��7��RA��Q,u���Z��70f�� 6)LԂ@�����5���L�/�n*��Ss�����u�#~f���:�#E�WFن���7R����s6>�ƽhP��\kK�
X/���a<�:��t� �")�/7ޯ!=��r�����oY��;��}}�����W�F�2��]^��'Mv���_l����a�M<桕�cx<C��v�O�[�k�l2�#3���Y�1ɍ�Vi����×�9���}�m���VQ@{��s_+�ȼv��*�dw|ݩ gϪ Y��.e���a�7��g&�� #^�x��m����Lg�U'�C��a��:����Y���*���t��6�s!�.
�����+�_�Q��D�$q�Ȇ�Üw�sVd��O������_��q㐑+�wO�Ag�u�cD�4g��-��;.�v�߳���Gs�G+P���pP�n���]gڽ���c��@��5����o���PI�d���et�S:���-��S�)�uV�9�?ls۩Lq;P�G�]��f�����e�Gdn���/K���Qz�=��9��~�3·;�x�ϗ���׼���)��q
�����ߞ�aW,�K�J���`������9u¸kW<v�k�
�J�3�ʙt�����)�&������J=)�����9G��WÜ^������2����0�s#X11j�p��,ɲC�:�=�E��8n��b�F͗CF�%�PK��/3��c�g�W�5ׅeU=����j����n^�M�m5}D�\�!�GS�殔͎	�>�%��t�"ލ�e�U������
}]DGl9�h(e��/�u�zme*�s����a����.S��V�ͧ�Lٚ�ÒZٔ*l);{�S�W������!��n��GWu�0}C�y���kt��kT�7��]����l΢74]!�S�I�5pP2Q���Y����?PC{+{)3n�*��pE ӍS��u�
C�˗!/clo�qJ��S&t���)�F����т�̊C8�f�ܺ��')����<�5y��B�d�i�`P��/o��³%��b�����32���@��g�`k�:�����P�Q�9�3+e����F$�'P�+1>O�A�agf��p�Vu�'R�j����=hQ���S�qjzr���� ���4�B���3�vAƯ&�_r���a-w:M�G�l�W]�܆�|�@��E�"n[����sW^ed��[/�-݈Dz!��2����j�ge:U�]j�jWF��N]eң\����E�Yg���y&��j�+c+��Mm<f˒�0]����h.�4�0R{٭�·�����Ƹ��(�F�����N��-u_1`��֩�4��yx�&S�A�N��Z���c.=n�:kX�����)���Uד����3��ksC��:3 �5_K �:nu�ln7�U�n,Uնt�t�����J��#f��q ��,[T��1��Gj�Ơ�nvq��/�4+�!j��F�]��!)G��?	Ȃ�%6�L�,��'�[��(�Rʼ�i�#=ڕ
��!��	��0��"��o�E�h���2��щ�{lk.Ү��GQ�ݵ�۔�&�JY�����"�qR?�ٙ
Yn���j���H�3Zϧp|.��%VAe�R&;q��YEu:=����.����3���%��d�c��}j�`�e	���j�T,ö���ҝX�2�S���X5�:XctMn#N��w��N[D[[�A�w��:֤{���9̱��]��?Z����,�g��Ok���WV��BEy5�g �)�g���e��� �w5��U�d�T3U�,�u����$7f��MK�y��l�r�]�t�hږL�63��C�P;e�����9u������.�L�;y7v���X���W%�CZx������ Koi��bmL�/�u��E{�Ɯ6v��Y����1IV�T� ��A%t�-��ŷ������`Sf�Ei�2]=�y;��3\�)�8�9G�����v��!R�k��Z��\���wi�s���ϥ��*��ɻ�;u�R��eގSd�)�<���m���4�}�J�+��+2�2���9��}V0�DyX���^�+��ۡ�W�=)q5�fae>��w
�\����$��:�3�2�H��mebAW1�9s�����{�"(�i�
�EY؜,���Us�e\��
((
�.!QU�AW
faPv��BgavUQ�W)�p� �.���U� ����
 �*��\�'NE
�0������9T�EEF�UE���0����
��.Uʻ*��r�U��Yra��.A��UU�8T\()��dQU\�¹���(",�"� "*8#���*.Qp���q�UUES#�G"�$�Nevt� �FG.�<TUȇ�q8��DU]�WeU�@���_��(�:d�q���.���r�rZ�u��`��F�v�`.���]+Sض���.3S"�kfԌ3���m>e�ί��}��G��z/k$"���]�[=�ߑ�QυxSyTn�у~˧1}j��Kf��@Ik�х<%@�����oeۘϛ���ve��ZD>��o�BQ���:Z�zgN����u��e,X�EP���0a7{)��k/�m�q�_����W\+���#'�G#�A]�u�7����Q�b�~;��M���+z7�1��K���N����ryB��I��ۊ[��jw���o�; y�U��u�X�Hf�E�=�Ʋ/0H�UP��؆�L���4���&���{�OUjzS��/2*����&���/��̝�o�8㊦�*�OF.,�t��5[�ª���oΖ�/7�H��~��"z&2_:���=W�I�w[V0�ٗ����z)�)a�8���_ЩTQ��o}5P^@�Ƴ�(zɧ�Ίr�}NȨ�'��)�U]�Y��.q�c넕���y.�P��~�Lp�i��ݷ�q�ToI�Xv'k��eB���0a��a5yC49�sqә���������\k��z�O��c������ҵr��{â^ep�5);MU�Z����9��moNG��v��6i˦OG�
;�;�5H�q��Р�;�k#R��m���.�]ԡ]2]�Ϟd�R`R	|�xuf�����[}��.7j�P؝�U�#��)jg��h�r�^�r�Ko����Z�EI=�����L�����h�oK=�Y�[�S�S���3�i�
`i��P��e^�mS܌�y;�<�g�˯q�2�2�����cCm�K���U���x)�E��!�LB�����"<������,�5f)}/g��R�=V��^�8�w��Kgf�p�"gv�B��z:��ac�Za���c���ğ�ڄ7r\��z��S�i<�r)�`��xg���hT���C>V��آy/�q^�y��w?n�s�)x�(_�q��τl|�܈s�)�~~����_g�m��z���S�c[M޶����&�D���!��
$!йfBؒ����/_\& 3P.R���~]]��z�B���t�k��-)�{��#�z�4ԩ|��p����nep=8󊴈�+�����c�H�:���+��M�RC�]w�;u�e�P�TRu[T���8�S"nnZ�X�h@�>�u
a\KG��D	@�$:ԧ�m��{5��Ʋ��zl�D��2�L�Ȑ�iF3;���jN�P]�g�������KRٲ7��u�z+\�{/q@���&�醃��2��ҝ�AUԚ�gM;yрAe�x+2A� �T�L��\ƭ�K���ۗ�*Τ#ꜽ
0�ED�X��E{��"#|{��T�L{��&v��9�t�d���B����q��T"�s���Tq{��;�p�Y��m��NܾJa�m�x]tuО���+�N��1,��}3�^ELK�U��83~�/����ٿk��T���C��%�9�T�vAW�mِ��s2g"����<�+�B0�םԻ�|���<0�Єظ�{f�l����i�>ϓULb�������,�Nԏ�9H�5{�s���n��x����F�֯�5����^�r���ڙ�hvٍ2b��t@��n}�|���{ڴ����� ��n��\ �q��_N���S�y��̓��B'�a����}����\�ץ�;V��L��8�����"�����l�iVG`����c����p�"U:�+[��auc���u��ͧp��)�8�V�ȓ='�b�iq��|�V�Kx��W �8'(�����5��ՙ�k�����*kPչ�Ӟ��o&�H��`ye̼��R�D42S�Y�,����cϜ����������K�c�pT�y�\)�g�ra I�)B�a�ޝ��f��u���D0�HkV�m�j�a̘��<$���;�x��bg��]�G{�J�%R�G�T�{�*L��ڨX���ʄ�ޘ�ӏ*7��E
i2D�7C0���N�Y�OW���_}����<�8 ��}q�8�5lE����T�5�MZ���H�Pq�,�{Se��ى��4�[�|rg
�#�T�u��*�|+�J9�1�,͇D��Flb#Y��֞�S".i��g���v�u�Km��tV����2�~�`HHU�&`cۻ�~��E]�mR���cԍ1κ>���#_*�l��:{��"�}Q=��v���U-�l���p(���s7"Ij���Y�o �L�n���@��v��ʑ�0�O3���y9q~��Ƭ1����H�g�}dWh���'i�6κ�G04����?� 
3-��
U@23�u�0��3�#g`���xȍ��:&2�/�0���t��q�vl\�K�U��_L����֨�tR���U.U���>M\A4�Fom�=�kr�e���@aX�.�[I࠘��a�����f�@����<t���Wk�0��nsEbu��Iu ����P����OD�*s�LK�l9�?.{u#� �N�#��.�z��z���oWd1�9eEu���ؾ�W(�0%�x����ȗE�ܿ�O$J���g{I-a˫R�U�ֆ�G킄�O!^��<o'T�V��%�Buhp6�h5���1�"r�^*���������T9着�ꪫ��d�.�h|�
��]��zsE�s�]���N�[NrG����WU05��(�~;&e�K�脐e��1���Y]qYM���1Tv��y���!z���G+�E�%�Wvb�0�SQ�~�y>���yF@;(�8��VUieO~a�U3�ע�珉_]<����Y��f���Be���ZA�b�F͗CF�ER��~��^g \���W���vzc�����S�Z���Ɇv�FŻL-���jڞ�j<
9B�)�7�(��w�[o�x��R[y���}����*���;�f�[.��Ct�;n̵�+H��v��MJ���-A��⤱`�z�o$n;9�h!��3!b̘[<�t�"��%�Cy��VWI� ����c���V�V��Ք �+�<�uŊl���Ld����+z5�Gd>�/�|��OA}-��ǿut<|j�*R���	��N����T9���$.��#~��d^
`���'G�!E��DHʓ1gn{J��"c_%�:��;e
:�H����I~��8�0�͑o���xjYv���]�l	u1F�jZ~Yj�R����.^a��%�S6·G�;\L�Q}Q��^�s�Ō�p��J�euw!��u{n;�brѶu�yv`[�Ⱥ�V�v�w��Ճ����J0���x�J��*�'����Z�t��&��K��?�����������i��ӛH�:�ً�m�W:�6�#��DW1����L^�:��=������p��o�sP:��*S��G��M`c~�:�Nk��j��)P�	T��0���u8�3�H=��'�^ʠ�r��V3j^C+��`���%lg�'�w��bS���mY
:A؉�����,��!�����s՛�
b�{�u5yC#C��6�9�P��U���*yc�CK7�Nj)e�����}��<W��� Qgh�	���W.��8bsg�#0:ޭ�\X����O[x/��f���1ᥳ�7���.)B4�l\�6��Yץ�c�h�5��M�k޿�ٷ���g��g?��uAOx����eպ%(�5�Qnv)�9��s�2�޴�Ö}~����5���b�k��O2u%{����u3�E�Ϣ�g*>[U<�=)}Y�أ|�g�.���JU�ă�]N�:�%�=MdN�7���3��/���UAD'\1���.&r�0���f���O^֛ 'tC2lxp��^+�V]�N��el.J�?b��]z���Qj^2���m��T;���z�*�D�)�FP�0h�(�1K���iX��]R^a9�SN�f���ܡP�W�U�}흨Ns�ɸF��ʠ�D�ĳԠ%��k'��}-�C�ɛ��9:�j͍&yq@#�a77(�����($� 儩Ul"�AN�)��/���,��fE�l�p��φ%q7&��bVU�p)$W����.j�?Yi��:��IL��U�r�3��p�+��G�f�]' }]91��3-�E�[����&��̜t��7�7�/��BQ�!��s �{�!ڪ�\8��*vXǕB�_j���z�idC��5����x�q�|p��A���+,��m���r5�OL�u����SeN��6ٗ�8�$<"��®�zR ����]=_H.�쮌���ZQz�!5b�6z�f��U��g���BF�$2\rϘ��z&���b^;��q�����'vw�q2��`�ugj��.!�}����ٞ@�\߭v�|<��;o�j�h��N��t%mtLŦ�̴����U��^׼����v��S�ӻ����z5 uOW�*mIc.;J�����Tt��(�^S��o:=7�<�r^�L���/p^���,f4�l����Ln���G�T%�'it�nBj�Y�jb���K��}Fc��,��f�)�(W�wg���z����/̞('֓�Z�שL��Eªgk�8���t����܃�+��^OX؆������|oonP�Ȁ�3�}��T�!����^��nLb�u��r�������ć)X:�1��ڗ��%`��ғ��'I��F��5�<�\�sq	�v�k�4v�+|�{dѩ��o��G\��@./�@��Y��.t���4����]�C�|����zJ܆�9�4����Z��_2���:L[���&���w$V�UzO��kq��m=01���4\ɨ
��l3PF����+���e���0�6����鷤m�*J*V;�$ތon�=Y���[�=9ɭ؄4��j�2r�{a��p�����AD�SW,���J�qAphNS���\�	t�pE����u&K�7�f��#DT��ݪ�,FGe-��trV +-��vL��$����G+M�*aɒ�2��]����R�HS�lo�RN\��C�M�zfgWV*�i�������dܴnZ̙*M��=N���X��.z�.���{b�u����6��}�}����v���Οj]��%	l��f�#��|g[�
��\�x.e��x�K*�8e�XƱ�㔫�t����v�5o¥NF$�7
�N�5�	�|e6h$\�=�^�z����p+��`��޹ `���*w%:���5-��Y�\B7�>)����N��۸�z'��*�ro,+�4��^V���N�n���3�_\g^<K=�W�'�s�X
�6�Pm��r��t��4�!oT�N7��g7�����^@T�q'��+v�9�ȶ��H�����S�ӻpT�U���4}''TTe�	��<�f��#NrJ��俨�8��'�Lvq�<3;������.�E#�ʂ����5�vѮEENsL�E�>1H�'����nI���G(�k��^�Vu�ek����y������z���<�؆��rRy��n��Y9Oء��oP&\�ܝY���:VMI�5(f�Ky�mC���T=�;�n�/v�p�˙kY|I�C�ҝ��]���^��[;��&	b��I��Kxr,X�������X=���4������-��7\R}s(������W*�G�}|koX���$1zGm��}v�b�k'��}-�>����|g�	��7UM�9I�˃�WH|�z�t	%�PH��R��I�R֧��p��M�v�J;�U �mi���P~f��)9�	%դ�+f��L�Ȫ��
\N,{����p5��Ft�=cm���?P�]9�zwT)��-��z�w^l��o�p��A%��k���d�5)_��>�Yu��:��9�S\���Ĥ�!񝴋NY���)�F�B�C�Ag�Z�����4Ra��EN�	�\e�ՐJw�w	��$��.5�6�*l՛�+i҃}�N�?qRfAO|;l�ݽ�+�Za�V.18b�q�\vܪbjlMf=�ݸ) u��S����'p�Sݽ����WgU�I�gd���]Zו�����\hp�������9ɨ��nwU�c�qU�zW���-�t��He�m�#�r��YQ�
�� X���)���4ɶXk6�}�h�e7.��PHHH�V!�2��pd��R�G3�SW!��Bw�T<o�yu'"Ќ(�S�Yi�}�k:U3n5��}����ù�<Vq��Wa��Y�sg�q��$�M R���;}]����[(Ա���J`�%ݲn���R�ݝ��
[7�������rgZt��:��ܦ�s��Өj��\��L�/�h��#\����N�ܺ2x�u�~�}K8���F!qJ9k�'�#�{6kT�7f2A��E��5B����ts��w'������K[�r o��b�k��aK�!�G�ƙU�@��H]�2C�Vp�l>۽C��e�H��ض7:ݒe-RD(ep����fI�U�����K�6w"�c��qϤ���:\����)���u�o��W�i�/)�J�,�^�joCrk���y������G�������5�p*a�&u��9��T�W5V��c�
�n��]mh���OR�و3p֟��1��Wf��u����x�u�y	�m�\���톧v�w�D�h�uXP���S���z����ŧBڳE_G�ƎC"[MT�飡h�lFΣx+;�b=*P��B4�v�e����,�� ��T7f�֞���­p#�����+WMI�o%��-�+
Yp<�����)�)fj[%�w+�"��	yv����qWI��R�f>�+��)P ��2���흓[�º���[!�$u�NwZaV3�l�鷎����-�1im�d��zy<ܽ.��w�p�N���'�6�yZ0����6��u�HS�`��K�d�x�Bl��p{��ؽ�TWcf]��Ĥ��S�ú��0�un-	�_ .�V��yV%��N�7``�1u�¥b����h�R��7W}b�J&`�4=G�S�{���B��q:���ޚ+lM�h D&� :��ʶ3�����([��@�KnG@3��.��mt�ŵ�i�=�8����׎���1��j-SY��]��ӳn�&h�)a�w)��K)KxY��4e�S}�nAX�y�x�i89�Z����G�En�F���C~Ò���&�����o/�oa��#߲þa^�Σ����zC�3*�Rش��`V�g�D�X�q��4�_Q��Z1�)��&�=&Y�<P��U#@�����Z�PduL� ��2[]-U�阷 b�ق�����`�ʮÔ��㮧���mG���[�dp��Vt鑤�&�x��r��⣪�k���$��5yF�g����u��z�Y��ud�嶟6ҏ��S��h��,s�.H�Zg��ud�Վ�[��ikҶ<�EE������4�]�U&�UM�2c�9h8�#�+_����'�s���ś�ǴF��*u��x.�T-R-�����Kn͌)u�8���5��~�@���
  *��DTEGq79l����0�+�UEJ�eGI�2�(�TAUE]:+!�
)��%XU��� �V����T��ʸò�9)�&A@���w9Wd�8UW)���"a� .eʪ����ʼM�.2���9�(�PW(�W�2+�Eە��ym8E�*Dr��L����AU�.�J�D�e���DwQ28\�� 5��A�TavTq$��DUr�e�"� �rex�*������D*��(�)r�L��ĕ4�	���p�r��t�A�)PG .Q(((���<`D$$�U��C��e9\9Ie��^�s��}mf���A�i��u*��yx�T1�'6:�o,ŢC؄x����-��3�{7T���}F'�������GZq���ro^�¼|�v�'Q;��+]ck(T��T���y#czS�b�Yx�<�߫�.*��YA��l�9��#ҖW����f�Z*�S�J�h�1�8�,gԋs��!����n�l�8�v,��.��x��NAônPl��K%I�_���xb��m��}L��9ȼ�� ��:�(�9`۳3���]o�@W���or!���y����SE�[8K��3f�0�S�j����4{�u-�uϚ�w�@��U�M�����R2�}�%v>������\ܚ��5@�%��ګ9��+���֍k
���6U_Ι܄�����z�s��&����j�+.�un��\��<����8�s���NC���祳���a�J���"�\KÁ���y���>[�x�j�cquB�Lr�&�0̼c\�����c�v�f�M�52��E��
�C�W�+)�x}p��~�Uu�<�6	n��<YP,��[m6�5��˩6��:bۆ�V:ɔw��厧4��ܤ6l��<�[��%�D��� ���]�/�Q��'΁�����֝*QU��K�#��}���C�z8�o�T��� �G+����H�tA)��x��lˀ�sb�Jl�*F�s�6)��
���	ܜ�w�n�5]�~�ׄ���l�)�{ܑ��{�8m�<�
�x'J�S��ߝf�Y��th���u�+UD__��~�d����Ɲ�jp�7����ї��N#q;��+���X�Vv�.�������a{Gg}��w�x�Ljq�ls�7�n�W�.5N��n|gh���tq.!U'S����i�z�ς��k|�|]�dG>$�F��d��u�{��Z���v�*%�u����rcTtA�f�e��z�:�э��R�Ģ�´����rv�ʉCz�5���:ܞ��`���^j�zb�Y'����}L�����|��t
���<Y(Ǳ]�X�ء=�,|1��TH����e���9M3�3��� 
��#�U�.�A��zE�6�҉ycWin�/[�0|[�6�j�M(�(S�4�[�v����[A�C)^�.!��1��|��&!�W����s0*�+{�s�ⱃ�J�+s�d	�r�_PtCWpgr�;]��S�h:F똞d��`�v�V�|$B�L���P�vQ�Y���e�k���.�|s\;wV�}�̵��_6���5qrK�/w:��:f�_]da�ny!����3�����I�5�ft��6�T���Ӽ��Ļ��A��нS�0���Z�8L.f�d���y��b���v7�n���
��HJ�?%n]7��
y�L,�=%եIc��8����|�l��:1P��sIGL�h�G�bJr��������~jgM�湣�����\��6*�4�lH.�NP\���kyCܹj��-r\(fS��\2�h$\���x��G<PT�DN.�O}SX���uIt'x�VXO�6��ȍ���7�>)ؼN��q=p^�<8�s����f��QҰ��H	��������������z��BT�58ak�ݫz;��9�\sj9)\u��.v0��'ug�il�T��s��^�^xp�Y�=�z�}��ZQG�{���<ݛ�w:���Us��|ѽ���ziw�
;B)�nvc�88N#JY�:�\W����+�Pݻ]-h�R�,�u%#Ӣ��_Q�>��uM���|�U�CK������qt$�<�z���'8Z6�s���E�#��K�"�{߽���>��/���^�e��ҏ!�&<e+�
���Nw�z�6�����m�s�*�G��oR 1��[U���^�H���J�w��si�4��;�	�ӣ�ܓ@X�EẺ�v�V���r:��P�p��Y��:ܭ���2�����N��[Q��)~)X>yf<�]�J�#��{���ϟK���s��	L��g�If�W$����3'b�,���Ö���B���kX_w�# ���Z�����=�"���?���(�BO�d�Qb{3��!��9ԟC��Y|�6��+1����鷬mä)	T~&\��Fzw3�n�:ʡ�xD��zX�qģ�:idC�l1�6����5)\��F؀����4��ؖ��9���-C�d1��(nGҔxE\E�p�J��t��*G�̛:��Q����erq���ᇭ:���p$�㫦�YX�jh��+���w�I��k�� �&�z���)�؅��]NשEVֆ��1|��ek��C�ɪ'���t��}I��Զ�9�������0��� 敊��j��}/*F���G�	M�,�lZI�r�YCb�ix� 
�&��I��G!=@�^̀�w6����ȼfV/�2�1�9�\��\2��^��d^���o�F1Gmi��f���sz
�Ԑ���{EWj��+�`��^;c���/F\s���?�fsW싴c����|S%2��
ǟ6F��d�F^�r�>SΜ��W�fW�2.�o8��m5>w�����v�;����8�E���;OY�ˊ���Pg��o�������ky� �����Y[q4���uEDE��[���d#���"�:�"wee����Kp�q{-\�<�)Ѹ�P�OSY���ˋ}�m5{���R`�拫i�f�� せ_>���zK�\Pf�@W	R��kgXiÎC�$�y]��ٜ�l�r)���yT07 ]Tg�sl��e�v��9���CcsfM�z)g�x�Q�e�N�=؂Ee�#=���[�/'h�%�f'���5�"���fk�.{K]mK7�er���nVf�Ui>�]E�V)����AZ;��pC3������;y���w:"�� u��D���p��%E�_�
%��B����}<����tȺ�<{"��>}/��]�1(�8~f��$����s�k0k;)��]�?�ޜ�v�\:gq.h��Λz��:J�nQ���1[]�M"�"�����5ͼ��@��t�}��t�Ȇ7�l6zn��鍧;�]g`͡m6�%V�k�u=#��WR/O�r\gy&�D0̼�5�MYٍH�n���歹Yg�H��) ��?��_�F�i��88�i��ʵo;�r�z����J�תd&�
��NW�v��e���y�ֹ�j�\�v>,Eq��r-��
ێz&��S��^0w:���؝w)z���%��r:�����jp��7��{w�Fs���yfu�T��$�$�-^��ݾ����3�%O�58���<�V,ʝ���kG4�ן����;�ؕ�;��W׬�
��޳γ{-M�lX���\,���V����Y�
�C4�W'*��u5ɍX�IPS�E�,�2�����U�7������s0Rqu1DL��;�y�NL5�9�W��kz
����|��lu^�4 �H<*��<z"ȑdܼ
�������� �FU-2*uf)ˁ+�D3\��۞JA�G^�*wl�V�VV��rruA�g�[�X-���-
�S�(�4�QN\ZӝcM�;�8�:7֡������Q�C�vv���S#%�u���A�ލ����!�˹�7�V'��d�e)�:�n���u���c���y9�{-�Ci��i��;`�S=*1��[=�T퓌�H�h�qC��+��ٺ������k_K���mtܙ�a��w�X������Bf�����y4��0��[���k�69繞׫'�RO�ɕ�'y�Gꛜq�
��Z�9�3V铐���Vbg8�4�hgO/Q�2��\:f���W�|dC*����B�TL$(�nk"�B%��ı��S�����m�<�̜4g�����\6��S��Gvs�j �	)�h�p�2��Pد�ણ��g�	w=R�{>c�JC<�w6}�]f�D����xt*�S�Uę*�����S,o'�Te㍬X���
� 雽�uЋ�l
o���sbe)����.��
mm�{o2��=G ��{�0m:��Q�]t��^sV�+�-�p��Na]!���I��Z��^�]����"��f���r/��s�6*9����"A�RZ�f�� ����v��{F7�\#x��b����N�A{}�]s�SUI�o�Es=R����D��'_Ӻn)�ٵ��z�:��d�;��PBlm Ň��'��pL6N�üzgj'��WX��-�<��sd&�����in��e2��S�?{z��}9��yS�W�el�:c�</�sG��OU�e(sYQnw�z�6�����ۂ�v�*$q���:v�^�e��gRW� \$�u�����-�E4�E#���+ӣ�-� ^s�&�g�v���;=@��+���T��n�A�e-�M3�S,��=x�=�5�u���WJ[�S�2�^P&��,���sx~����>��L�(m��d�!���c^;P�.��bV9�dz��v�=�����k[�sŕ�P���ѕÞ`t$M�IL���#���X���SB�W��>�B��n5�i�ҷ5��vZ�hh�W�=+�y�Oz�~�@\�H�b�Z�'
��m�[�kb���	F)V��(�vc�̦�ڠ�1o:37y����":KT�bM�ۋ�O_p�V�]�E�����j	w�rh����'�#$ߢ�ӕѧ��pznw]�E�7t�Q'�{[�6���HT!(�L�Kg����X{���JW{���8�Ĝ�M,�7�ߘ훆��LT!*�5)H� ��i�s�TT챯*բ�bSv���E���e�C�c�
F��31�t>���'�?��aG�VA)�2��&l_�'-ˍ{1���VYb��9��!.��D��mѝ��^э���x���B]�7I�#+���O�4n�A�[_s�5�9ꈜ2�מl����oEO���%��Js\o��HM�l��N�Lk{H��L[���"��5�����U^Y�\�'P͔�6�:˔$�Q�S�^�����)ݿ�r��������z��[�t�i��<���B�܇��w��I����Vcr���V<�cl�����d �=`�KT��X!��m9�q{B�Ji�X�d3 �3:X�¤� ̤��9����Jr ޭ-��{"��;M��b:�U�G�ɺ{rde��E��X+�{��b�O����y��c��T�H�L�{x��5I�^�S�{}��y��WO��j@c��|��Q��FS{�a�]zA�|�p6�<���tn:�%�=Md�sk�}���(wB��@+�x���d�5?U��U��o�s=@����7֠+�\�|	85�S�}Y��2QY}��>L�4�@�77&������D���N8n�̬r)�}���4U�����O���!����-�;&�y�[u��  7�%�y>E_d�9ݐ]�t�tΥ�s��X�8t��ܥ7����S#�����|-�pON}�5��ms'4�!����鷬�2��ov��	�K����Ѝ���t����ڇ+\g�&�Cˍ@rS؛|��.Wy��.�ho�0n$%s�>��Ӹ��7=�y���B|��OVb����6�U�l�+>a�<CaR����Sϧ��熑�L��o�j}l)��<}R����dv��%87:շ�$M�6��%�1'*-]qS����sP��VY��ua���4ut�����+:RG��II�9ӲV���P�I4�2�d�e�,Hu�-:�ղ�[5Ql���1�Y	�vnk%,��R�v�һ8V`td�h�a�v[�����Lwk70h@�I���I�p��b�5�훤1�'K�sb2�H�w��K9`Y�;)Y��Uݠw�i��25н墎d��+���*�A��hm{���0���Wd��K�s{\DK�ة�eԹ4�P���&�Vv��rR���</�z��6�咞���K)Y=GR6濫�� ���0G�>���I*���yj��o{��Fݰ�Q�7�ۣ�)#\�ݚ�zb�Ӎ�pk�#k{�����S�;���A�g嚽2*?��sJM5I'!�A�A��tL*y����1(xp��.�n�a�(�)�|�(�c�q���ڝes��ɷ��pM��� �T�h:��X-뮘��T+�"81����˓��N��r���hE��r:���w�b��1�ڧ��D/�N.�(�J�)h�SY�s����3X�]���\vu;�*7��5��`��t�g37Q�1+I��i��S_le������%�vNl#�\�X����(�ھ�1�P��u�6��ob���N�����k�=8*mY�ڋ2��L������tYj6-�VL�T Z�*��L�����_;���"�7
����9Lc�j����5Z�f�*1"J�vc�`(vF��X;`�������6i�*�fW7����wu���<�VVJFm��jޕ��TW�b�yZޛ�!j�ZL�ھ��oo.���B}�R��|y���7"�-1��9r� X4TZyT�՛I��V���lu����Kވx���w�4�p�s;�7��N�Y�^*�D!���
��e����}�&�ǜf�㫍�����!z �Tf`��u�6�d��9m^k'r!&7]�]9+5����c#&�Ì �7����3�o8��|��x�t�}��Wp��!���A"!�]�'`X.��d�,o�9�oi��N�_ �Ƹ_Y5������Ұ�v�PDTvR��}Re�2���j�7�sH��[V�q@D�x���g4�W���Q-��n-=6б/��h�k���cp�V��Z��"u3[��}���m�'%�q1�z9�<�{��T6/mf+Y ]:��+n�k��p&�S]�Ǥ귻���CZV�ZJ�9>�`�L ���j��u�%r�Ew�^��a>�5n={���VoV�
h�Akˮ�����l�����h�dw��Y�|��m.�
仡薅}�������ĥ��V�w�T��\�:�۰ݗ�n����f�vR��sdh��aX� ��[�����ͥw� ��_,�|��������I�\.U6U$Ӆ�¦EF�j0������!��	$Tr�EQ2r!�)D] N�$�ZI*�(L�j	A#� �ӸD4�Dr�L�QE	�'5dTI
l(�����UIӅ�QE�I�e!2�BBr��9\v��#Z�YBr�(N�C��Rt+�S!R�Z�@*(ȸiA� �v8��ȳ���8�he\��2��W"��BA�Add5�(��,�IR��TED��4H""��� �A&T(��\��a&�1����EI4����eБ�ID�Qb�W��Nr1�h����LI&�Ъ���LQ�dY'f�?P�T ۭ)����Ƅ�-fi��cB��@;�1{yɎG���.S�N��u�R�I�W$����uY��hBdɒ`��פG$Κ�^Ȓ3�>:�V/r.q�>B��9蚧�����z�l�����z<�u�K��o�do.�oN�Ƨ^7��s�g�rF��7Z(�
a�h�w�]��ŗI��Ʌ��mt�F�w�u��J�jq���oK�1/ŭj���.��y�HS3��oL��n�u]c�[;�yE^��*{9	j2�ݑ�T�e&ʲ��cK��ٷS�0s���Z�xK��J���o��wV!���-%9�+�;���-���5����'n��G���P�A�$]�B�uF�6ʦJ�!E�K��}��YL�a|�N����_H�cȬ���{M���a]Ր9�>v�y����{��s�i���P{��3���:��}|P�Z�
J�s�w�f��-��e�}/Ki�k"p
m�Hv4{��<�l��g�@�f5��,�����I�5�k�m������#V�(���������q��L"��D���̃�[��/��~u�����)�Z�*�hV��P�G�,�� (]]-����f���6Rv
���Nɼ��p����_x�Y�}Y�xSs��hK$�ڨ��쇑�S|�t�� MF7h��Hr�9�ܣ�;�_%ӑ<Z݈CM�f��L�BzI�'t��|��Y��OM��:�!HJ���T�.���"�P�7kF��.�����玒[���p�连1QJ��I\D��f�g7���wv�k�![����񝴋�2��>ڇ��@�A�'��7;o_$T�X��p��K���.�6NA�7��r��Vv`
��'��9�I�7=C�Q��oh���ѼE:18a���d��o� W�eS���:&�959�~���5�����4�^]��5ұƉ7&�zg�~�vi�V�{�?B�/m�s�wC�j���Ov�-���l�����Un��H�������>k`��{���>��*"}��+EG�F��x�\\��67� �7��@�*)�9�9��ׄ7����~:�s�MI��r_��r�.�|rj�8��J��|� ��3�}k�*>�����R|���"��mZ&`mj���)�C�w|36b��"��Rq�Ws�L��C�Y,����LB���Nu޼e��EFS��.2�l�٘���<�o�e�+{0��r:���}��8��ys�)^�3�?�'7	�>��Ȥw���_�tp;FI�{��9o�d�;;s��#qA��BY=F�q)��쥹	�r�d;�ZT���m<A���!����Y���H*��N�B�k"y��}-�S���"�K���C~MyMU��F���2=�{�ʗUU[Jb�}I��F[��J��������
�����A���/�s��%nin�<%u��^��su�֣��!=�͕V铐����鸇�m��
BU���f�j�e��5,> ��sH�%.H��W�SK!��훆��t]Wn�+�L�v�n[w׼�Vd��\���_j�3�	��-1�V1�G2�Vܯm��'��(3(r�[g�״��|Jwʗi�	',S������NdN����U��E��W@Ń�tb����{�(�����۴͗QII�P��4��T%��P���0�Ƨ����E4�fK.�X(�2ɍhb/�d�lV��_���ds�b��]C��b���=[�$���5�I���������g!7gs��KhF�,�j��u϶�cJ}ճ�m5%�C���n�h�x��K�z��(�]��m�<�B�9����Uke3���e����'6�8������p�j�u��XӾϵ8c1��}w�ˎrj'��Yn�l:R�5�i>�,<-*¶�θ���Aㄜs[�ޗ��PF�[~���A��Nn�&�wUI�}u��9�i�z����;OY�{9j�f�M���xy����
G:C���Q?U����|:U���QjA��1.�^ݹ�ݺ[9�o̯�7 ,�y��ϊϳ���͠��~��T�+���٦��R�=Ѹ���q��OgW]3�u_�i�����7�>y��Fb'1gE�S���K8���;{�os�ɜ�ޗF�0�US��z������C�Z�+V�\�������uh���Z�K�i�bW7&�̘��,�7f:�9%kR����Դ�AW��V��K�;Λ��m�H���;ȱ0ן��q�I�̻�d��]@��|[I+���ʓbz<��L�5��+��{��tT"��i��_�폭��/��76��(�<�bܽ�Ef(7<*g�i�hwX7ǰؔ��b����� d�]Mn� ��Q�hJ��јkC�G(ծD�:J���/��K}7���t�\�a��cy�}�H-��Jr-�n0�-)�[0�'�ޗAE�^,�ˡS"aeD�QsQۑ�<��\K�׷9ӆ[o��1P��%s� .uq�z�	Nfb��
���ûo��@d��!�̷.5��ڗ��3�Amы�yD�d]ἡں�-r\(nS�=p�א��bNE�?z����^�	����9����y��<���iӅVE>ݥΏ�ϭŅ;���n'z��������	�<��y'!!z�s(w,�}��r�=��1�%O�8gN���U��7�C�-�% �Ջe��y9������lA�z�&_�{��}��@=�a\���5=O؞vlL���OZ����<6�R�$�\����Ot'O�U#��4�b���6��{�<cO	��֨�����%��Y�m�u��s;:��L��γc1�|&��%v�H��]Ÿ���V�x(׽㧕v�)E��U̦11�<�v�}sd�͓1S��q@�9�m��@�vӸ���|�1f_K[}�4��R�=�DeL�/hJj;�
�RUZ܌�:۾�#©w�U�<2�-��]��7��N���N2�|�<+��G��Bo���;Y:���o[O�[5�;pv�Ĭ�Y�3��f��l��c���]�q��m�C�oq���m>��G�3+L��+� ��5=_#2h(,�@֒�Ya�}\�=ƚ�;��1W4�4���c���7�Q��ɔ0/����T�A�:��ʋ���u���g��~x�Ns׹y����G�g.%�a��A�.�I�V��I��s�����=������p�뇌R�%1�q���U�����hi2�{���ۄ����e��9��V��#&%�jC=��V^<OV�)W���5��;KP����Вsp��jr3l%kw�:/�}�*N��;
�nc�l���{O;];�'GE�����:�M����u6�X�#�5Q�ɀ�tP�R-�Kw1^'���9bA���m D��
<�VV�1wD l����#]a>r
8b����F)\z�Wԏ]NG�;p�:[��[Ȋɛ��u{s����B)�J��}Rv�x���!^_������/Ўݷ�J��8��M@y��Z�w�B�_*��U�C{�{���}^�^7�/�Ԫ�VA�\�C3�+�c]����z�z��4�oVR2BƓ��w&��޷he�c2�/TD�Q9��JLY�Q�^����f�[7\W�Qr���<�w'�yǄ7��oьX��'3^BK�	��}��ގ��x)�O�R;�	�e���B�;�.��H���aeD�����	dD��JN��M]�lg<F�+���f�R�3_X
g6u8�o��k���y���ʗ�^`�Jų"���ͧ�q���QL���|n�/Xou���4�޶�,\��w�jZ����zv�l�a�S��J��:^���`Υml��)]�f��T���R�t�s��zư��_���I;&�����4Ӛ�40mM�5R�z���u��X�ӃCĠ�[�1�h.�Z���3y�iS�ЄQ{6��H{����s	т+u,��	V.��b�ǌFu���]���^Q�r����m*��pI3#��S.�4�&��ؘ��$3$	�^Y��)�A�y���X���o�[cz1G�*�']����WZZ8��-F8��_Z/��-��[NWJlk���q��l�2��_!ï�]�OB�Y��%5�̩�+���U���z����G6�_�8�C�+�q��/%���/k ���sZ�����y�x�1+��pێy!U��F���xn)�&N��LJr�E�Iz���oo�x�!/_f�^7=m��sї�95��Tk�!��<[�}�'�V���9��v����%Oq'�:�Ǌ!U��0k5�ɭU��	)ɍ5;�-m��S�yE^��*ns���n��;�kv`)�wi�
?k���.�j��5k�K��WO�Z�!XI��G}��ח=�d�g���y�'�::�ܘUr4�:��0�D�U��۶�6�i��\��������Cu&�5�f�Y+3"3�
�{8K���2D�+:2	t"-h���`6��Aji�t�R,�+{j5�*��q��������y��RX��s�M�́r}T����ѵ[Z��i�F�d9ܵ&�F��}��n���գ]�QFdd��>�i���W�]5���+/�@ˢ|�@5Sh8�^��
%d�|��O'p�[̈m3��9:�7&��ꀢ�q0�u�Ĭ⑾�'q������S�e��콸mŴvL�����ǲ�!!��.g��*8�f53ʚiä��3��m�P��}�Q5�̵V�R�q79O�4%Ӝ[�q�����o��y�F+����N"O-G0��9!��Ak�&�@h�$c��SϢaY=����a�]�؉g*�[�C��}S=� ��� �W��v�E�U�]{��˹!"��놋�/!��NF��M=CΆ>�E4�4�|=&;��V�b�ޏ��[L��I9ێymG<T��<XHi'�����=�OxKTr���)[˭ŐS���.q=C{j�i��K��m�b~�(齽T�دxl��(�[��K�H72�))6�LXT�ԧVx�@cў������3x�>��9�-�e�̻)c}p'�{�M�B-2�3w%��ZPc0�rDåq����h�d�4�f�T�����wF-V觡U�򩦍Bz��l��J��e�M������ټ�u[H=z�5�j�D�n�Ȍ{m"�"��m�ɪ�A�ۭ�K�/CW�����~�n�����5n�����{��O~|��M�s�c����݅<5����W��"�H�!���}OY�mq�k�����f�)�9�-2���p8�NS{�m�J�q���}���si�g>���<�}ϊ�Ha]s=�[-�)�)HvzAۊ�µ��D�r�[��r"���^��S��m��ܺ�;�8��neO\��7�`�7e����Q��F��U�^�z�d����3��5�9����$�e�p��\*OmͳP���!��&���A�Fޑ��+�������8�iX�q3N��<ڧ��wNs�5�o8��:� �V��2N�}�_�g{$�W��0���W�4��OH��qqL��4��r��s����[��T��2��d��%ʖO?�磫N8�/�]��Z�M�F�)�*��u�Rɣ��Z�o`JK��F�YIh�r�
�ko"�6goZ Z\��0��p^i+�=غ]X�{�íkhȮ@�f��6�.,Uւ���-�	D��9h���t�vT��B�+ޭt�7:�$��ո879D
$HV��ߴTΥ�Nv��XZ�'QsU�#��K�ӂ��2Bq�1�誔Q%��bU�_L�}D��ɗ��ˮU�`��N�k64�����P�-��L�Z�����iDL|�=���)�8X�9��P~�(*A�]��R�'(5��+����L��yj��s����L�I���Xj��J��F�s!�ux�'��ĦjNۅ��)Q���<R[Z�fʻ�B,g8��s"s��c�T5��v�ڵ�̖�܋��{��-U���9�_5�2^��57d�����W�ښQZ�-�<zģ�;��Yϭ�ĭ�tw4�Bt7E��q���
��2����1��bU� �����r�FDu��Rw�OG\B�}yʺUى�������j���:de|f1;��E�̩zy�?m���������1����h�����`�e����[�Tۙ	Y�rև��������(ؑ����,�[�R8.�Df ]N�UJ.�A#P�e5}�E!ej���V�+i�:����٭K�Q�pr�ݹ�h��C��l��T�ٺ1��SxǙ�P�y�Ε�4&�+U��:��m�М�Oa۳WIՂ�b�b�,n��j��qe[��LR`n�N�xv�b�F�V�,��)ҵ�n��h�¢�v�:Tʶ��ڣ��$��l�P�Hۥ�W�5�<|��jPuaPU�FS��髋����'{K�l��q��2�t�[#���s\X���v�E�����o^ur�v��)*�z�Cb��GRWwYħ��e&��#Yz�R��N2O��[�+�Z�K�;R��N�Ү�Rv]�����j�(oR�طkk~aj�M7��w3��S:���w�S:�Yo/H���+ξ���Gx�Ap�]�x1j��0�=v{5pZ�d��(0�}�$�H�GO�����Ra�dY���ܗc;�*���m��1Y]��k���8�>���eD�)2l�0�T��������\*�o��Bۑ,��v4�L���y}uU��Kd��nn
7��Q[�}�B(Uim�bR⻮90�'K��ź)s�]���cS���	��_Qg�]M�4x���s�����k'��F9%�}�i��qW���w)�[���`�������M�Y)�C"ŝ��E��;�����E^�=�ol�&/v)��EL��=��A/5ӸA�J>W���8�����FܬZ�]�w�tOlq0�ݗNJ�?�Glʙ�Z�z�w\�=���:�!�+�Y� 5Zr�I��\H�2U�֢���]"�D�p��"T��M��X��]'.p�RLN\�!�3��LԐ��Qq��q��ʍ���I	�4�"��KB�UD���E'Be�'em$(��eMNԔ˅Sd�Ւ��Z%�#��*�L�Z���
i\V"r��erÉ�0ن���Yʤ��8^%RU���*.�r\�d�&I�IK�)��F�ji��� ��I\�隊�W)�`�t+�VG�S-aWJ�NQ�U��̒���$V�5���.�TU�fg.��-K$��MJ*,F��Ҋ��(B��R���h�㜸���B�+OK�Y�7os�R� �-DKc�=���u�o=j�;��YD�j�ݎ����p��{\��%eo��q~c��	4��kX훈m����!!H����M��f��k��e�v)Z��%;|go�m�i�r��j�)dbsw�����s��7�����c;�E�0��$��n9�6-�uY �΋X�H	�4�zdK��sl��N<��\���Fq�M��E�?o�<�g3����\u����s�4\��]t<ΥϏ�WTfjT�,h�T�6�	j旾�މ�����m��LV^�ukx�|j�}�,�dH�su�IB9u��*{�>kc�ɿ{zݡ�.�/C���V�Fs�D�)jU�n�+���θ:˔9�qOY�oz��^��j�OYV�iT��IN���\jy�:ۉ��N��:��$[���d#�(r}5h��]�F�IN?)�f@�m���<�d�4+yCd�,O��`�S�q�F�݈[w�&�;adf�J���-h���J��p.k��rĳu�7�Or�6��{�n�s6�Y#�
���֏v��e&�̱�t8J�h6�*�$U�b�fh�]0gc�5Ǥ���R�@�T"�s�(t�v:�4��������Da���g8�%���z�E9��]H�Pf㭅���;��{��ڡj����惛����i���nnMAS"T���/�WV�PE���*�����!�k���zqZ*nI������j&2�v���*�I��k��+f��)c:[�6��c�q��1���������%ɾ��+�G̞���}oG�����[����P��$m��ы���˜}�#n�D�OH�}W�Z/�Kzs`��C˻'�:�ROZ�zT�l��lW��2�l��xJ�Vm��S�T�)�n�${vZʺ�2���ب�s"8��H.��ۀ��Q��e�����)T�7�VD6�^&��ێy�!U��F���dvOZ�ns^�	 ���
q�����mu�I֘�ወ�����9�ˎrn��Q�p=�lS�&���o�
�o�K�s�ʠ��/��s.��շ\z�CE��H[x���+h񮥽/0vh$@ܜ{o���*�K�|6�p%i�X�N��.��*��O`�a�E���d�U컱ʗ!�r�D��Y��,=���Ώ&d�S�rv<�-�I�SH<p��kc�ɸ�z����2w|S�{�h>��n����g������gV|u��Ss��7���:X^�{
���d�;3���({c�Z�A{��gR��
Ӓ[���|57:�,�����_�[�'�
�R�<��i[�N��<��ڕ��6�"T �晸��}�[MdE3��<��6���T��	�@��Q����'���J¹�o`s�H�7oe���!��꿞t���|
�y�S��R^��n�+��Ѫ�S�fZ���᲻%�14yJ��+����ԮR^��u�t{�f�I8]�S	�K�;�3�RI@½��K�8�o^P�����"�kv�k�r�\�vNv��"�����_u�h����s�D�����r>�R���U
b�t7,=�9/ZB��u֚D1�&��9�%�&��uf/[�C޴�e:�-��1"l,T�a���u⨬+�D�Ν����jen��f\o{5�JOl�������K咀<1�/�mb�	�WX�{:��6bd�9�7�����ދ����,��cB�;˙��\P<�rK!�o�6�跌T!=NN̖ꣳj��n���E�\�n돋*��H��2��D!��N=Re����,�T�\p�>��q�3WiugĮE�0��i'!7�!�\�V�bC�}���ً��l����u@䣹�m�do.�o�\bp��n'���hi��uj�:SpR ��S��N>��7�l��w���ǟBT�#��g<�ɖ��2D2��T�{ݎ���X^���}4�w'��]r��X��~5߹tߧ��8t��ӭ�9g�~|qc�iN�Q�ܵ|N*[�=ۃzr�z�Ȁ��!���8w���v�Κ��X&�WU�j�_%f��:W4a���59�s��9��D'��N�NI���2�v2��Aó��#�1��jȞv�u�[-��!���p�5����7�Oe-MA9�f��	�cTR�J���J�p�s�����hryv�,X�u��B͌Kz���$;i����Q �R��o��/���g	39���p>k]�|��"<���� 8J�q�s�n�jy�Gz� 7%jT��K�.�ke�]씤,��iWfz�7VP'���6l��>}-�w�����o��(̒��쁜b���\ɠ�},��	��µԹĐv����bb���M%22���Wc�}oHۅrU���;�2�P��	 
�z���et��#�������N2qg���oX��!HJ?.J=����d�S\��$��JrI�Cmq'4�!���O|�p�BS�jΙ���f�6�-Q:������b%6��rE����1�S���1{P��ۖ�$���A�H�Oe@|�����%;eK�L�I9y�EVK���覹�]�JFE������MAs�!uļ��w>�/�#yr/�l�MV��W.�A�����k(m��:\��])�g�4�Okt�N��c�����N뇷�>i�dF�^;�K+yhˎRP���֕
����n*�W���2*���ښ5��N�W`�T Ы2#�2�{ Wk|�Ò�R5��N��x�A����x�v���:
}L��a{)���#X1�<K�o=��Bk���n�'���[�kvV
֏[�m�]��
�Ρ#;Th�rJ¶�θ�.�:˔tBN9���ɿ{z��p\�c���ѭ��J�9/�++nk�����
�r>?7{��s�n�ј�pn���Ѹ�1ښԆ�3�������&�3�:��:��SL����x�|���
�ԓ|T���*esⲳ��3h)��j�H�
�|6A��@;�.b�-��{���M��{|�꿩�=�Y A�������%�֬b�Y����{�L�O�<w"K{��3�M3�3��ɢ�z����N1A�=w�����׌�yrj��{�:�ۺ�E>�e�ϟK���]�1+��G�EQ[}�L՗Űt�EN��Y�h$�u��v�[�w掳:^���#�L�n
��Y[��qHΒ�'�/������ߐ�p���饐����g����0����4ZJA¦���U��_U���P�0�OH>���0�o�s�����i�6m?!g���0U1�%\8Sܳ!CO%�.�s븎��OkL9(�ܜ�+]nD��q�[t�F��om�Q���/�v��S���q��C���ĚJ݈Z�s�,TGd]��e7����	�"���9U��!,p��m�I��[��g9��=6�ZY��"�1_ ��	\OH��՛G� ���qgYux�N%ظ�2y��l�_0�B=WU2�T'��F.�]A:`�ͽ��|�]T7i�z�b�(ظ�܋��s��<��딶]$�����!9�L�xt-Ƕ���7���FD5���!?f����� �G���ϴV��������~KT�N.C���K��{�\E���x۟g�s6}:���o?\�S$(�x���|+lzn9)S�וX<�����;�>���FDw�9s2�;�=;N���U��7�A�n�������?M=�&3M�(�����̲����3p����rzv�̬^P���"��M{����	�յ���1�ݙ[�qO!�	��
{"�迅�^�C��.t�"�J�:�)1'��:3��y߀l/u��0�~Yv=ئ��9����S���l9�����x�D����Q��\׫>gג�$��#=�<=�cާ����
�����j�Q5tl�`�r���`=wK��!�%��r�t��S�,��U�0�ӝ���p;�Vi�m�2��$!2�wu���ޔ��3
�R��SYv̽�᥋qB�J���]�'�\μk�QSU�]�V7��m^��lS�

�HR�'����5L�ؗ��+@T�`����an�1���D5���ߣ�}n{Ƈ�/y�x�=�:�{�9�[{;��EKlB� �x0��^������j�\W��g���G��:w�ߘG_[�nY������e�Z�x!�.���������X�q2�4�/�j9�dZ�+�Ǧ}�z�<�$�r����E��{֤��{�u'#�nj�uA��!3-���&���#>"���a�=�i�(���}��ڛ������4�x8�����39��
` ��t��hL䨼SBF\�l.�����S~�A��xS���Sp[W�ޯ <6=U��_L�:�� ���qz&d��x�E�q�{�Uބ�������/a+dg�z��!�fP����3���I���6ĭ�����G=���z��= =s��D״E�yvt�c�|i�&�6\�~̩���UV�s��2��׽{�0IQ^ّ���ϣ��0N�3�5�!e���|��\VzL�i��N�Zh��k(���ʳ�/�����C�j��{6A��*�rg-����$5��pT.�¡�y���.�f���8r� �/�V:�jL�ڐe(cD�QXuM��l�M]]���k�jC"�%���ܟqr�W�z�NG�1��HnZ2�D^��LR�vf�2l,������r3�Q�k�5�LBև��g��m�MCV�<�l�%�$��Gݎ���w~���i� ���L��+hnr8v}T�X�t�9���5�Tv{s`.��g��D��xh��J�<����5���V��/�ڮ���:��8z5r�Ʌ�򅷛�y��J���T��ѱӂ��U<�_O<���^��E�߂ض�8��#�����,z�����R�>���y�
s�"���]W��8�X{}y/b'�~�8�}~��z߂�Ш���^˭�Ǒ�T�T��
�h�����
��p)[�!�2⒵�0�O����U�-J���g�7]���V���w��,�{������⁙�<�&=
OΣ�D���[��6��3�c�Mwwo�{���;8�ly��x؟�US�ۗ�0*��*�f�[�H<���{>����k3I��xius�{��~�ZA���`h>�w���)�`Ha(���!������=�v
��O;�>��^��)���(�ʥ%C�cb7�W���g��9��E �vLe5�J���^�!�u�bj({ʮr;^��^�g�+�6���c���}U��
w-z��^���a���!Tt�Iv���$i�E=��ԕ��Y��f?V���y{y��FLGc���(�Ej�	OD}�v��a���m�:���sy	{�N�jw�E<�q<�[;i]Z��Z�c�Cg�`o��y�!���������K�ı���|��1F�ɪ��m3~���M�J���؟K񻩣���ڽ����P��^r�o��!^�/�q�<��R/�Lq*Y���=����rW�j�,���W���{Ł��ZUt1:�tݹ��u���]H��x���ղ���'r�B��|0n�=����z��f�܇��0������\�o�'}U�9��>�WJ�~�'I�+�d��f{#�~ �Ɵ�iő�W��7����2����=6�`�9~��Jc=�Ǖ�]�)����W���C���`v�nf�=;�{}#�/��~��'��Fv����b������r�<��tF1�;�T=����9Ƚ�����o���o���N�^�HvL1��ћ4�q�}�l�!zթ�7�6�9u�� �
��A�{~�@۩���n���:���^4�Fdg����������)����(�T�e0W��W>�^B��]�i�s��՝�/�i�x�Տs#���~�����p��E�ߥoնeg�0���}_Y��x~w~U��cY'�]���gq�)5,QJ���
|��y��r��*ul�ȭ�V˼��%�+8��"�|�y3�5��M�չ7x�s�c\b������t�X%�+k �v��N`bt��@�� ��VA�!�w5up��VQ]X�/��L%�)��͛4T���������J4{���S��yڇw�T�s+��pI���׽Υ���XԸҩ������.7!�%�:�C����J����� ��=��x*h�����V:;��$5���͌o m3���nk��y�9�xh���EK��������C��V�����}Ϣ;��#h��vu���(t�j�S�Ŷ�d�w]N���qu��E@Zq�Y��N�I��"-����YnZ����������5b�G��;sZ����Ŗ��&��ڛ'�S��ԅ�c�?b�ou�sh�����W���D������Y�9���uނ���*D�QQR�M��o2�v�M��w{�L��m%:�1�qnc�Su�� �Q6Q\�r��\�s9�+V8���Y˦q��yG��	�=��Ƌ3��s�Β��oe�+B��H�,��x���	����w��$.I����d��35�B2�{�R�aѽ+1��i�2ɾ��nB����c@��z�����PZ ��*]���3�P�Ġ��ɛ����j�S/wR޻v�a5�hɕ�l����Pl����G}CM��2cڗ�{�0�	�O�>�Z0NN3K�$X�]B�,�r�v��/c��:���wH��h�{6����e������9Dt�5�^�5Of��uf|�*�̹°qǆ��Һ��z�JL��I]�㱫�9�R��@8�e�`��9t���3��ZԈ=A>�v���P�l=%ȇ���W��̗��rT�%�g6�:�8�e�ǚ�v��"�N�d��������@�Ԕ5��oE�"�����X)�����$�8���"�sZ�Ƹc���$,v�ʖp7X��ZU+�����ćh�d=9��vn�v����$wpөq�|�V�[��d���`*H;�4q79�]��!�,E�]��s.�+�v��;$�`4���u���f㗟Z�n_C����iNZi�Rm���l��y����Dhn�[��H\�j����r9w����W������l�1�o�kSz��&�����LX��7�27j�vt@�&�`�9�[C��y��¡],�����t�"�֥��u���q
F5�v�E��S����[�q`�D�F�M�]�a�\tMP����GJ�Nb{�䁻U�C�v��܉�i�6���P$ũψ��a�W�u��\�ḫ>���1rp�K�([}��ʕ� R�tҔ�r��e9ȵK�����N���fF�!C���Z��<�NYϩ�i]�|�>�J�"��j�m*T,��!%�sO�P��	(-i�f�VU���t�I\K# ̉bi4��$�x�TbI���,�UjH�*T�*Q �U��Dө�ҋԢ��Xq#YF�J(ĵ$�C��Dp��-�*S*��Q��J)
�EE3��&)�V!�%����WR�T���FJX�g�qr(ʨQM&��i#D���N��,� ��"�b"��)V!VlL)Q4���P�4C�-d��Kf��DZ�U�y���4�4Z�2B�dTyJ��Ft�%r"�*�R�����i�H6��G�8�tp��:JA��.�Iĭaea��B"�.D�(�B*p�]2H�4���.�,��h��r�N�XQ��4��@|  ��H7��ؕ�zh�}5*/�4`��7��;�OYG3Z*�,l�R���#JT�[(Wv���W�t�!��oJK	H�g����4g~[�^��M�O<G���<hx��,�dcČ��-1*���e����x�F����zf�}D��"������������_�ON�g���*����Cbv�`�;���|P�B�(h��@�*�L��lМ��/:�b��}jL�����q�I^�C3i#�ك��'�������(��[����Z�e/Y��)��棚eh�=E��:*a{�r�Z�1�-e]{��z�h�xWO����fg��`z���R��hHf�c~YMq�7��}��7�oo3gt��z+�5ѷC��zԏo��fO����<�B��L7��d@U��SY_g/O����9<\�)Vo�߻-�lo�x���~Wt1������̟9��>ʡ��;��5��z$�G�b�#vw���~�Ul�".���;�7�q�CW�?]��s�_�do�� 罝�l��w�ϙ�^���j�d���dO_K˯p��X�xӟ?�Nfϧa����~�>�8���x]��ŷԊ��H�|�t�_~L�
��$C+���W�g����]Q��L�;���ݘ5����#J�_��82�gX�ӷP���������%cnzL^��I�M���06tfl�l�6�K]�cU�N�����s�[�5d1��udo�AԹ>��{u1F�3��K�P��f�S[Գ-]�P�zf�nKy(�C�)�×�U�9+Ձ�k<�W��������4�ڜ�۩܅L�E�<�mW	��,�B��7��J�1�P=�3�i�	�T|�S���~mٕ�֧H��+�)�z.������]uUw��;����X�%z{��2����g��؋����Szk����$�iP�mb��*��o�R��e�
w�T}Q���:ϡ�^Kؓ��uh��`���<�V�Wc[������z�O�vS<���jc���(�Ԇ��.���T�x�&��zL����Ǎ�|z����|k��wQ��)�@/F�|+xG\+����4y+�6
�6[s�?�Q?��g���}�~Κ�=AH������%��G{�pY�S\:�~�����p*M쁐j���.
V��\!�U��uKOߢ��-S��9{֤����ԟU9���WL�uc�&���!�*��p{�ݮ��QH_��55G��Spr�67�\G�;�o�d{��3���u@40]6�m��=�dfob�Vj��X�DS���D{/�*C�q���ͬ�xy���]�=�_L�α�.�ߪ�WOd��OW����
�kA��tW-��Y�:�����O0o����j�ޞ�Fx;�/���. *ffk�M��^ᙆS��K#�Q�o\t�`�X벞�j]�P�\�tIl��������d��Q������d����}im,�jc��)&Ԝ�v����R��}={7�,\�\-|^�>��B1��1��}�d�fI7�y�Mb���v
���#�#i�Ξ�^�j8ۓ��f˔�wS�ocT*g�V;Գ;�Z/��^j�2��7'�U#��.'jϦ��*�v�YL�.+=&\;C�|��{:��+�����do?\�S��l�2=yU9���F����"���_^o�/�Z+c����� 1����zw�w~�5��j�ˀs�i����4�'�aU�Q��ds������c>^`!���+��<��ۯx-��A[y�C8n�t�|2�݆�7�y��X�}UӷT��=C����*���V}<��1�^���~m��7����g&�H��nң��Tߕ��\=����ND��!w,=�O�%�Oz�"_O�Ӿ�R)���C�z�����j��o´���ۖ]���&=��]y]L�_�wQ-ӺP�1_�
���q�r��:|ѩ�A3I��>��{���Q�r�� +�&�����[ƦR+���wW�-]a�J)�iƚ�5u,[�wz��[]��%�;7>oۜhɨ�>���$��7p����SfE��]��R\0V#�/j,Hf�r�7��f��|/�Aksl�'��iVCӳj�3_�G�*�W Bo�ɹ�ek!�Eh�U���D�+�}c�ȼ�[�p�:tv<lO��r���v���0���WPs/[���W�w���+)��
(/����_���Hk��G}�P�=�ʞ�U�W���>Ʌ���H�v�v�{ȣp���bj��# �L9�b��R�߱����y��Q�3��E���3�4\{���4��^|*P����lME�W9������X'���z\����������P;NR�����%H�p�\tM�{�\!N�ȉ���lS7�a��)[�g��>��ڨ{꼩i�����,��T�<]���^�>sq�=���H�T�7"����qt����m�<��MgO�I����}���S��yC#_�gՑ�g�H���^NuԄ<��|ëe
Qآ�2v�4{iF$=�%Y�Ǡ�x�!�L�7��߳�������o�'}U���V�X������+�*����ϫiΫ��p_q���ǔS��o�]���d��g��66�U��AO���y��-�B�z8��^�_�����8-_��m��gylzv)���G_��l�L޷Y}�B��+O�ȠX�~{�Agw���Kh��a�I]�P���]ҒC1���4�&�wц)���n�����D�Yo��&��I`JF-ET/eM�$������²����K�;B�,5�mh��B�VH�]^+�$�j'$[%g역�!�ͺ�!�;�T=������/j�M:��?D����\�xT��͵��������O=��o�o��O��mNr�.|DT=(�<��]����s-��ʪ��X��ߌ�^�Tl��I+纏��=n|���}+~��6��OfS P^)\:���ruo�n��v�;]���̏,�Dg��!��}~�4<=�7Ɲ�ߥmm�Q6�N@8g�G,L��&8��ԣ�S>�j�.�*s��.���㼛ƞx��ʇ�#|hx�ܲ�Z��߀�Q9��ʾ��S�U{dP�3�p(�Ԫ^�M�:�Y���z��G�ا�[>ƇG�
�>Y~���V�w'[m��;�K�w�X(���
��١8j��wCec>�*w�_�9�װ����q���+��>�����E����\C��&%����64�4<y����8�P�~A�c(�ۮ�Ł~g��x�}^��#g�{ޮ����dUê�R���hHf�cs.2�9�W)f���K�!^�~��!1�Nn;!5����zԏlG��fO���yn�\*`��97&�����J2��ܛ���H���O��ݰ�KZ�6��*���u�:6	�XG~�GOXy\�D{Յ?}qGo/1��@
�m
�ꔶ��¹���M���Vz���]�'�&ڻN�-�%�m@8�����,��mI���Y�!:3~ܶ����2��yC�̡�?A}�z�O����=�A1�p��n����縪�`U$~�[+.�����M�dg�f�=OلF���~����H>1��W�;��\�R�IpR����.�!� �Dyt�����p�ȅ��~�n}�i����^�؉m��+��9t���4��J4�גDw��'!��hϸ0;�B���p����0[���㙒�����o?^o��iX�EY�WG�g��U���vm�D�[U]�E��1�+ҋ&�׬�"jθ�����®��{��NR���q��n�J�3�s�m����U=T�dZ^̹�=�|m�-Vs�~��]��)D���k�/'�~��=���C�{���jLi���.��{-�t�*��
Ŝ�߀��0��uMTa�sN��^K���m���>����ez�^�u�S�ԧ���y �Dpz(��BA��jG�s�J׆��n�ǎ�o�zL���>�<�ʔ�s�7/=z��J�IZDx ���\~�'<G�\���~���)C`���lB�\W���3s{о�t��{}.�WY� Eu�K��JKE��A�7sU�����K��=Y#��q[z+���e��%C����{m�߫Բ�$�-^�r���d�ͭ��,��I,�԰V�VD����A��䎵8f5���,X��Jj��Ϟ7rJdg�|I���+{�Mp�n�ŀ���
�A� d���
�Y�>����=��}��'�y�-R�א�����߷�B_���$|�q {�~$,��2�n���M��܏F�h.��r	�7!�cc�i�����{�f|3¹� ��^�u��۝��7ğ*>\<=Bj��7�-�d�!O�#�M��mg�{����/�~��{����������)$�=W𪂲$���z���n;D^�l���b}��2�co�(<^��BPں��K���{bs��lz=^�@_�x!�������E�rs�6\�y'��=}�����a��]��S��7.�#ޯL���ӓ��u"�xs��MwY~��2<n3�f��Q�7����	{=>�f�����9�����;~�
�ɜ��g��õ�;�yac6}�w���tp��<tx].�Ǎ/�N,��;�p�sU���<��Y[Cpӑùn�[�ў���+Hԟq�^�= פ���	�|�ĝ��� =���wW�xP���tYY�=�'{�H�x<���q$���Xm3#�ti�[}�8Ͷ,��GY��νWܜ�7��4��^�y��<y(�5���B&�X'a�A�qˍ�\BP�w�vɆtߡ.�ў���LU�験q��
�\1�[uD��9Y��*���{�謀 ;2^�|����{�h~m:O��J���΋����YGW�롾�Hn���8�[�Z�L��آ�y��;|T��{Ｐ�ˮ�ϰx�9ۑD9Ⱥ�!�qܰ�O�%����'܌{Դ!}��y�$�g=���`��j|�ip��!�`s&�T?�� ���\Ry�xc���߮��z9�NR h�SF�}�x�{ö<lO�{���mmY9A�\
�C�ᜐr����l*�='�IJ��7�s"�ȏg�E���{����6'�g��u=�����U3>Uݶ!?'G1��*QS���dc�����+ƣ���Hl:��Dt{�8,�����[��=�Q�k��cO��*���8�n�������2��_CPϙV�:��!����U����ϰti�s#l��A�Է�\ߊ���U��k!R3�Q��5.�|pObK����PwS���y"���.�vm�h����lO<wp�:&��h��z�Xk��V��k�F S{��ӝ����	3�Y�9n��½2|��f_��BT�7"��>ʍ�f��C�x�=7;�b��1J/�3��zdI�S]��wv��n�"��:��z�ѱ>���Ծ]f)o�����fZٔʼ-�Q��&��AY�c��2��sv� �8rX�LS��Ɓ��)U�Y�d�g$
�\N����ع�DU�vc�)�7S�s��Q��a�4�w$R8��hu��^�Dy{oҟ�����d{��=��^Nuԋ�W�W6Y��G�"��a������*��{�~��#��@��ח	���7��g�2#}���ܜ!�V�f��/_�� ��+�E�X,�xO�Z"/m�b�d8���N,�m:�p�o�g��f@^���۵�X��G%��=o�`�~]�T���WK˭�ӂ����3{���;^�H���4�; ݿ`#������ד�`�(G^Up�����My9{W����؞�3�84��tQ�e5Ky!5�¦��r)�`�"ݩ�6��ϣ�]s�"��j���	��m�g�(fG�S0V�����ޙ�����d��	\u��R�;2䌮��U;a 8	,?N7��X{��"Q�����g�)D׆2�!�_�o�v����o��(eF$`�&]n�c��n�e�:O��H ٟDI��Ⱥ�z�;r�n�o���#|�x2<@����d3�(���b����D�m�r��L�q�3Q*��a�r��x(�g�M�z��zw�ϱ��y�������y$i��� �a�ɤ�On�*bρpA����<LSIg��+t��׶0+��b%|�O\I��]ºjv�e��Ă�N�����Oca������9f�o;��3�u����j�9�,6�]�&
fY���t�ó_b�yn�{l	>͢��C�[Ȯ�W�39A��e+2<4'>5Kλ��+>�}�T���-G�}Q��g2�#B��>�q�I�z�=�Ȣ2=~��b��!1-��4@��F���hxƀ���<��W�Ѭ��hO�3ͭg=�<s�z�ho���2=�Y��o�*����]��o��:���V}��͕���š{�clw�d?��sqɫ���H�ǅ�fO���yn�\*`�^Q���$'Er<w��﨏|=[7M_M�����FC^�k�̡�?C�u3��1w>���WG_�۞���=j�zB�������yK�NGc9齎6�Ƴr�~�"9�+�7�K����7����)M{bFz!,��Z���k'���׸t�t@�mϳNfϤ
݂G�`��e��������y���|}y!g{:r]�V����]�E����s���?�~;�U_R)@}3>��c���~��z��U����9�u:�w�C�>UxZ����#�5;F'�����t�l��fn5�r)Qn�Ż�f�veo�z��NǃW�?�}N�^��Bl��Z�]Z�)��d��*�f�2���Y����l���\��Ӯ�O��x�K�N&��*�f����e� �Vh���m2�LW{�Z�k�PGZ�55e�>��Ǹ�'�$-�J h�n��*��;����3�B\���bQj�����W}�H�շ��U�����$���E]�6f�dR�Y�to$\" �Kc����.���ƻ�����c.�����#����Л0�����Z�s�F���y����j�H�L�����d^Ս;zYDm���7�sTP��u>�v��5�.QB/wc�m^/��+�(s�9�a�q�q�+� ��Vh��<-(��t�炌u�2����by���8�f��X�Vs�G��OQ�(ne�u�� @���u��&�LvJC MYF��Fo7u�n:pb�\�	r�՘�N���E�m��r���%��N멂F컓�uu-�	ǕڨK+��fo]��̳���v�LTsZm���聛���]��� �
1�f�(�_1[7R:y5��F\tOT�j���08��4s:�ENк��y��D�(f}m��PكL�z�a*��^N}hv��Wc��í���̷�E�鉥�ch��o�q�V��l��'N�j^IHc�[aD�]��Q��I�\��V��v՝��Hef����>w�nۋ�b��1�4s&&jL����nK=��})k�o[�42<.Wk�ՌUڊ��wYi1̚��f���������hp����
o
]sUh����R���ƀ���S�9�����K�&��}�H=�5���vi�k���\�:Ϯ��+R
��J9K���[V%�Q��{��e�p����%PvvvL������D��W���m��K����KM	!�1����v��9�9z����v��� i����LH# �M��Z�,}˦��%rc2�r�]���b�*8�sN�/�*�����^���������մ-��w9�i]f����w�1*�m%�^��Zlͥ����;�|9�1����ĝ�F�qE�Z�xY��gOn�d�x�����*�qH�]�L]�º���S%wT�
��U�ȍZ�P�*흯.��v��+�Kv�N�X�V�(+�k�v�+���5�b�S�|R��i�B��V��-�e�c�dX�:�i��m�)1/Wܥd�{Y3�f	ei�3����1V˰��7k%�g��I
.�ԣ󐜠Z�\�W e �T�E5ك��>�T������t�-�q �>�
!�fҥ4��:Z�V�V-\�(:�1�p��VB��련^��Y� �h���ћv.} ��!?��Y�&�����SRsLӵ�p��	�or��$SS B�^Jꓫ�Ci�'W�9�`Q0sj�e�cp�{O�}�+C{'[���y� ���
���� |mf�4��1�u8J�)f�e[9B�U��9�bWBT�fHJU�4�P�T�T$S ����K
ZIE��B!���P�r�uNWH��U�)��h�KE9Õ*�i�t�h�ʨ�$���\&�$�F�)P�H�mI���H։̔L���%X�iJ"KR)S+��'2���Ρe�j�	Q$�B%R�I@�*�U:��\���,���ȣ�"�IB��G-B8aa���TYJi�ia��s:it�Y�M��U+(�9V��DMh���VUb�(�R�H��)%CJYb��Ж�F�**bq ��	�j�)�bme�H�\��4�0��H�6r$P�VZ�$��V��V��Z��QD$a�ITZ�J*tT�$�t�5h�%T��EZ�+�%���*�ef�

�(�4�ʕID�t�ص,\��|y��g%�͞�gJx"e�S]�wpp��q�[3qJ���
y+F�Q��Ա,IS���֟��ʣ�X�r�ҕ~�$�����c�-� ע^Oz�Ct�<{=����dq�v)��}1�q=��f�L��	n5C�ў����.���>˪�ώ;�u���^���FG�Ǉ�l{��k<�k�;B��'��'�i�Fz��b��}� �.��[�Lc�y6ׯ��O�-�{��]��ճ#�<z����G���y��< �	�SlD-����<�΂�'#,��^��Τ�k�7>��YӾf�����d{�Mp�v�}9A��	��&�� ���/7��F��Mn�W~���q��ȼ��j�u��{֤���4%�����'U��(�M���Ա�#�=�T���ײ1�h{��(d2���C~�������z�����g=[�Y�����OGgo���_���]w�@4$'JoV[@��)�g������PϽ���c�]�=�2�f(4$G{Iz-� ��*�6��UC�I���G��#q�"�+dd5���B%E�t��{gܷ�8��7��C�%^�/c���5�� �&�W�}y��9�[�/���ׯJ5na�X襯
� ����W��!�]L9i>���Rc�/
�����ee������X����j(������I����t��Ň�t0հ�C�`E���f����c�3e���R�wY���h���h�3: e�J���f*�p2y[iok�^�6��tu�@z�ob��p��>�y�:�S��{��q{zrO��GD�
�v�����/��1́����=���w�"��������9ss��W�k�K��͐F}�u��ͺ�Ȏ�\H�^��ۑ~5gw��'W��}�>.��p�i�g�qg�i����n㚭������eX���W�*tou�^rJ|dp^�Z. ��E�����%o�ǽ�ׇ�����wzg;�����=����y`��Fs��p�����Y�׬t�w>U<ʍw���^�\Ojswz���l�H^��8���##�]s�0)��H��C�;�ğ^KM��mq�ʫ�MR��{dI�4�}��o�l_�O��"eR����T?���E�$=sQ"Ҝv��3��;���۰}�9ۓ؟?gN��{ö<lO�}�c��[FVNPB�`"N?o�Ʃ����%r��C��+H+.��r/"�����G~�>##ܮ��ۗ�03"M���9y�|k�3Y^��.��!�7��5�E��i���
���˝�6Q���?�`��&x�:o Dj�-������zyQ��Q�5M���o��}wE�*��۲�04�����'J�ܛc�զ�m�O���Uq��w?�tAO�ϓ�q�]vp��mX�N�֜�l8S�rS�-\6x&��|�5Q�J<�/�;+-�jrUk����U#E������ё�S�s��P�U�Z��؍�W���*fd����߻�-�i��E��7�1p���4$J���.�>��{�g�j��;ۇ4�%,�w=>�W�<����m㸫�)�0/@8 �3~���ѫ7+H�0�ݧ�o9���T�V	s�+��ۿ�
������7ە"�S �H�d`��!O�bO�O��X�^�)���Vo��9^@����׻=;��F�\ϫ=���؆:�r��E���*���`x�(�ga�x���\��}���dvS!�P|3�.���F��������C}�>�1����t�,�p���UVh2�O�����^ߧ�e�Ɵ�iő툧W��7����N�P�`^�1�GI(�*.��G圇�
��!���U��q=]/.��N@���m��Fw�ǥ��?S�<{�9�R����-_x-��'��}���ۮ0;�Cۚ�r/j�M:���㞶���VW\T�*���w2�m�S�k��~��ݩ�6��Ϲu�>)�(n��9����U��{m��G+��,�X�����8[���oT2hY����*����I��C\����.�/~�������h1Ӵ��:����Uf4��5(�&ʄ�����W"\�w�^�{e�U�Å�:So{��Ki����^MY�î��JA{[1G������G�T�`�&�adD�x'Qn����?�اҶ���B;u=�L GfFz���F��G$=�xQ��G�S��3�^d=����<=�#�!�V��~��[fUu�*���\��^Py*��� uFf�%��e�7^���t�<w�x���T<��=�q��s�Q���Zʠ��+x�!P&|��Nf�%R�"�v�>��������}jL7Z4�]jiw^���p^�\V��v�<�r��2����@^u��+l����y{]\P�L��m����='ޣ�/w�(���늶(0�b[�WԽfǮR�����u5�^����Y�I�������ho�t����fg=�ȫ��z�d������nH�;�"7j{)��G5�S���������+!�g�����z���R=�3<����!�=��}�Pv�����rW�O�R�χV��R7�y�����F5����<���
��g�^��g�B��R�B}��g��e�Q��������Pլ���6��k7!�~�"
܏;񘜩��������1��1+/�b�Ko�l�)�z견��f�du�s����+�O�<�v�n�y����c�Ӕ-]%]�b%�f�D�&$�+dG���7*�\zgY�o��
%#;<A\��X{�8)�@R����u�.¹�T��Eh��PD8�ޏ{;A�Z�gjϧ���]{�NB�d�mϮ��Q�K�U���|�J�y�O�j���~�>��^H]�ٹ�u�80;��P�Mwy{~#V͆a{���a�ϖ�F���~��S3q�Y��{�^�sнy<A�R�ٷS�07dC��ayz���敢��5�_��ȁu�؞�3+��&��m��f��fVǙ�9ʶ������_^v�>�)K�:_��E�)�{/�ha�q>c`�K��x�����C�u�q�}몭��e��(���Gr@��[GE��$��_���J"r���������}~��{�x{�=U i�W|��QgԖϵ�r<�V�p��H_��xS��A�Eҵ�*�0��M�/q��jv���W��)	���2��o�6<G��<tV�#֮FT3���%1lA�ۓ���G��y.�q7��VqB{�W�Xu��G��:|������jk�C�p�'(1p���X�q,��}�KU�wZ���#�+)�=�(.�.
ϖE���J�u���Z�{�u'�Nk�PtN8�ǸvP���A~`�2��~���p׻/������_^shg��s�a��`;Ϻ�|Qy�na�]�۬���vc5$��ن�5�� e�5�i˻��ڸ�����Cn����S�Ge���2u	��3��P[�� �n�L*ή�碱��V�RG�C��or�<� ;^�5MY��RA�CT�qo���Uq�������n6wݗF LB���O�U�Ey��@�$	�f�,����S��SQ�Y��W��}���t���ㄩ� ��/�oՈ	�A�R/lI���G��m��e+dg�׬O���>��[�6r��=�^�(�c���P����'�\t\A�h�/�A�n'jȚ�����:w�߈���A��yG2}��|�O�y��J�G��*s_�}U��W�Aϗ������/�󡊽,-�]N�MNC��s�.���_���~^��x�.��rg#Nnzu����s�O�y#��{�'"g-��e��+�[x�9�7�����	�z����8l#O�M���w~�7��9�����}�n:�M�/+���&�yP�}��p슯h����mWx'C��]��V�<}�������c.H:�${����әU�нGN��x����΋�/�~�W���?�a�O/���,����x|�O�#�m�-��8�_1�]tF`�	Hs�(�4�1���-�:%w��P^�-�ve"�g�8%���LklE�M�iy!��\:𒯪�T����󏲦��v�"׆,Fy0lhL�ƝhRd�%7�}�!FյƜ�hZ�!�N]6��C��tf����4�J�)<V�^�����xx�{orԹ(s��*${e�$�R'=�����O���֧�F�� �
��b���W��f+o�پ���/2=2�#��Ʌ�/�Ν��k��6'�=�s�6�����Z �q�̎n��^�J9!�Q>\nX��ߖ�E0훋t����x؟�US�ۖb{_�.�2�c�`+9�/5;�W�
�:���f�%��)�������ȼ���\�C���f1����yܾ�ʜ�T����(���������)�9�#�Pʵ)׭�
ʟ���}��k���׻G�Q�2=�dQ�]�T�C�\+�o$ؚ����c��a�O��c�|4=�Z?]<P�'̼r���ǃ�Wx�o�\!N�ɪ�쉣�5��Ӟ��Qױ�,�6O�$E{����n^G��>�~Y�-��q�^�>�2:f߷*E¦��R�<w���TOGz�*��	�h���M�{r׻=;��Dk������L��:�O��@6|׳}>���;T��}��rU� �B��@��9����^#�qT��9�a�f��s>��o��sR�_�]�pw���{��SǸ=*�1�%u�b��4;Аwb���չ�e l�Ѧw���
�1Q��(Sobu�{.�%�ᩜ���.�+z����:�I�>�놱��Hi�������RQ��+h\>(��=A�껓Y�'u^�#�l:jJrt����ZǤ `m9Y��t���Ob�d���|�r���?1X&�w�Wn2�<HI.��"wp����3���:��K��1�G���t]��N�G�+٫bڄߴu(��z��h��ގ�W_��G_���W;���ٷ\1vD
��<�����j|/ԻՊ	9�|�s'}��37�¦���C�[�[��S�k�9�����Gz\b�jfs�Mr��GU��_��]��<W3�n�kv$����9�w�S�[�VٛGn���b}症;\{�;�� ����R)���̇�}~�4<=���C��J۵Ro�}];U��W����S���s
@35�J�>[�LdC�y6ӿp_yP�dz������}�}��#^.]p���heC�/ξ'�L'/�7O�yo��_�M���S�3�s�=�EL�d��<K�!��C���{"�#�lC��_��W�}-�@^u���*5�g����J��9肖9S����;�㞓���}�dQ���\1A��&%���;����ۚ�� o�s�ZD/ڣ���{�K��#��μܸ�k�W�aО�T�I~������k���r=%]�:����[����7գqG�-�8Wk�rk���y��"���c��d��-[�m����0���\&?.��/C�&(�4���<�+�7)��x\��='���χ���]>=�Y����"��z�/Zݩ��B��ξ$�W���!�V5e9��r�C󛃉����jG���3'�����*c��/Q�^�P�% |�Q>�T���f�o��rׁ��S#�d{Z����O�P�G�0/��g��H�q21��z<.��=�@��5�iIȟV�˥ç;�M��5���c�&2#��޳ՏW�vZ�%���H9�g`�=´dA\�C롯G��i�u��eA�/��"�ι���&��	��z#ݙ��~����������ʪ~Rժ�gPz�T2����xC;�I��N6���6�E%Y��W�;|s�3g5���~��zσ����6 �ڜ�۩��S�w=�Z|Ʈ�C��r�^�c�
�9����tX~��37��9J�t6-�k4ۮ���g��8�t2��G�p��ܒ�����.
����vF}��\��']�3�1�n�0�᩾��
k�*��Y�p������{n�b:.��1���D��Q���r��9:ϸ�������Q�V֬�^GF�z6z�P��]Y!Ew{n����E�O�uE�V�c�[��27ZE{ݶ%����\��k�,!�Z��n���X��q�u���{�ĥ�[Y���^=rq�5-Ͷ^��KH��V&w9r��!����aA���~~�<�-�ZE�tR��{�Nf'�9غV�5n�1N|����׸w����ɿCG���[����s�y;���E3�~�>Jb�#��s���s���i�)U�7k�e�,�{L����d���ʆ���u����ȉ�Z�[2'uV�l-����;<���GD�ួ!�$=���A�+�Q���;������I#��9�5J�q��P2A�/%�o^��L����5W�fFMs��A|ʛ����#��}"��\L8�����Y�R ���u���p���@4&���M��h=��3�M���z�{�k�E�ۜW��o>>����4yUs�x_L�l	�A�W���N�:>9���[#��%L܅J^j�%��v.(��Ve�7�1��}�1q�G�P0��3�^�Mvt�/^�����vW%�Iu��~�������s�'�ʜ��Ud{��s����>کx�v��͞u����f�z<�6Z�u��E���S#˾+=&r4��a����>�ג8{��U���[�}����g��%���V��@T���d#�6ؕ�uܳ��h�ZUc�I��JM��R�����Ҕ.�=J�:���1��!���E�0WlN�.����^;|�B�l���7�<�c]�����j��[.w��g��J���I�a�$T-��%:Xh�e;�ң�CDZ�ʶ�r�:���(u��q�΁��.k*�$����d}���C纡J�7�(�1φ7}�I;/"/1j����C�f�O]{�[�[��i�#3U��]7��=/\��1��J[k�Cp��X����:�I5�WJh�U�5�i7s�`[sl0�_m���N��j�k4��!2����wM;�	��3Q�r��1s�|��Wa�j���mq�ᮭ���/�Yk��A�1��c�[*��:�T���m&��#yqj|@ӫd}�Լ����&�xз��(��y�f��ż��6�h�K��͍��/�Yb֙|c{���]�Υ=�z���/R�ہ��a<���$g��z7�+�g	[n�*��2���Re�2$��Ͷpw4"����5 �X�R�^b�E�y�5��Q��7�Y��ʺֶ�>��y���n���4N��vާR�^ٵ�ISf%}�L/W� �
�f*��!��}Gɏ�[+b�e�mZ��8�zuq���և��s�A�nw>+Sui��n�渐�W���|�&8,.��VU��V�����٩�L�ї6�FQHfE�V49.۬H�-�l�kq����βԚ+I�*���R�VCH��D/yQ���p��8!;B�ǵ��׽�;K�!p�;��r��Cxt��)_;��j����Nk�M��p�����0��ͳ�pr��*�u���t����R^���ْN�h�������������vWuc�{��olP�{ˋ�VݮG�XT�T����_��+�
�X�{O#�'ף	ʁ���d����v�u��=�;i�H>!��N>.nJs.R��A׽a��|�����]�59`���G���Mq$����"��6+WvYyܱ�UI�ڇI�-a<��K�1L���Y&j4�G:�����"^ODk"RK����׈��s`�4�:��bݶk%���Ө	E`��o���}�f�a��>�a�)���7���8ǧ�nLؐK��MX��]����wA��T�+�:F]J��};0�5���.�Z]��԰�j�.�;m�,��$��A%α�O��O!�7\��F��,]���=��x��Q_f;�V:��y�Y��R՜����ډ.�A[ºh����ɷ#��Z�d̦���N2��;6�(Tr���MN�EwJԿ��cY��gB�l��W��kɫx	+*�V�S^��c��v��͵y'm��ʄzL)�-,��I0|YG��Cu�c�)u��}}��
����u�·��Pq+�j��^�S��z�4��5-�Uv\�(�����;[p�|!
�`jD&��2�a�$4D٩Ej���%Y3RS)#���J�̬�P4H�u���\4L�FuJ��:�
)#iU�V�����*��(�S�j��XhW5%N�T&�0�YJ�iB&��F�l�&I�����Yh�d��DQ�(���R(�HZDW3eʓ"T��*�*�#iԳ�EffAY�JQa�B�,+�:IeY���Iff��r��Ӫ�JD�kN�r��Ek"�EEE\���P�f\*P�,�*M���DT�J�2�-Z�Q��!0���H��2���%Tr���gJ�E�T"���T�$�*
.U�9�#�AUE�B"���(�$�A+#hTsH��QEr*%�,��r��"�$�qJ#�UD	J*���A�9�EQI�PEI	QAD�ČK�EvjU�՘��I(_��%MU��9h۷�]s�E��j�1��lw\��n)u�M� L�9jS��ȥ��Ʈ�:�Z�Q���Tv�jC����m��A��_�	�HkU}���@�s߂z�~�Y�}�l7q�V�� ���s�[;~��')H���o��Կ�ڣ8��h{j/n��K�!�����,�lE:���57�8@�c��:it� ����
�AG�:���M+�����j�+Կ9�6\���$d��O�ϰ���Jf���A���߂ض�8�_1
#�]�<Y���"�s�U�71VC���Y�����G{�f�}�<��'O����?^�,���v�� dC��o��bW�T�}���%9�>��C!�\W����b_��;�5�߼lO�G��|@�e���j����g�Z�Q�@���,S�[s"�23�y�{��u������+��@v�.j������J��*&�^��3)����}��F|E6�y%�y�y��$6Wx"E�o<>����ڍ��zyS��
�U!��PC�$7FGH~
u��1�jS�>չ�\���w��l_��1�mh���z�¦��-]Cy&����\�,v�	��r��W���_Wd�Y��8��q�L���(�#���]���f���~ .��A��{���	^�ybH����X\�(�J�y�OKs�0)��N��:���n ;��b�o鷔���Ld���u<g�&�o"��f[5� �h��I��P��
In������IX����K�+�Uw�{<whS�s骅�:#���B�O}���I�KU{�c��D���>�v'ҟ�eNCn��#�=�dt��]H��S �|�lUm�CXI�撖{�����qqI_p�íG�F5��N�󼡑��3�����${a����K��0�]g5�I���Y�H�S��F���������T��yp�~�#y��}B���c�yל������w.\���
A�I�OWK��N��d7�?6�=՛��˴�?&�x��%�=�CF+�^��������V�Cë�*�?�'����3J��Ӟ��>a��̵&��Ũ�}��;�{}#���c�z�x�_!
;6� ���P�漃����.�ē���=Ud�u%z֏ۙ��"z�2���}nG���۵<F��mN}ˮ��.��v�xfxs\��c�)\5^=s-�I��Y��x%p-�8����߯اҶ+l�eiy�E�ɐ��$׶w|�J[��=�����ؐ�=R<�9N&�ϙy�����G�vǎC��/��3ι
����E�?u
�U�r��\��д�b^��rb;#��!��*f��;Ux,=T�Mu1\/������]���*���˧J�
�=&I\u�'eq�u���JWb%�gnr;Coj]*�a*c��;5Tt1����t����@�_g����H�s1�P����t�C�y7�<�� ʞ8�7V5e��l�C4z���r�fF0̌����L�X�3Q*��a�s��Y���r�Fw��W^"��y7�vqON��cC�<�p^�\V����r�
�W��١/�8�q�7��~4��J�ٻO�xQ��>�*v=~x�c��='��D�w�(���늶(1!1-Ծ��ُW���|��*}�@�Yc�)���\��g!�<s����=���2=�Y����"�������;�����_�j��T��} К�F�cS@ޥ��3�����z���R<���3'�7�Rl��v�\�q�u���ϡe��_Έd�V��L�M��ca*dc^�k�̡��Y��5S�B��z7��(y/\�{����ؑuQW�N�.����]�E�ߎzo�>���yl)���bjf��;�;}�	��^�'�Do?E��F���{c��
фxq;P�O_K��.nT�՞��va��e.=�??_�������c~��og��*�*���j�ɜaA�$T2��j���}�'FQ𼜄��Uv���I�귓gJNҕ�!{��r����-�؞:yM5�ᕪY�[x�CS2�$zC�b��s2m�i>�%{��ql�8LT&2����B�[V��E�C���p5�n�ە�ʺQ��_ے��:��ر�X���%jV�Do��g�>����f���,��;�w�{��	�ߊ����=j&r�IV_ǉ���Xg���W5���8ȃ����mW^�bz����NE*-�طq����2��L��0ng�j|�J��O�
���2�
{"��.�^�C�9N'�h5藑=���/�P�XW{q�ۍ�4uaX�K�!z-,�;�Szkht�z����j������8�i�C>��;���#/z�x{����{dy>��O�lE��yo´���C>�BA��Nf�G�s�t�xs����>�j�mtTت�>X�O�Ǡ�^M�}�<���S��Pc�W���D�/�< W�3�L�|`zoѶծIq����'�ZMo��q^�g���}�~Ο>�0\yX�Ԧ�n���**y��nS8�^o/���xTz&�%d�T�t1pP�|�/��S�� {޵$w���{�y���Rt�=�y��5�Pڿ	�J��ME7fFDMwD1pP�T�o��߽U�{�<��ь�~�ҋ���yr������y� ��t��hMDS�A�_M�B�P߿���^(,�м�Ѫ-�jϱ��+���\����yz�j�z��Z���r;��f���͙�-5ud쭬(�]�5Ю�0et��ȩ�k��[���]�md�{���Wt�����ViZ{"�E�[�V����p�9�x7u�Se_e�\tt�^\���z�b%,����yW�o���{a�雇X��A�V*�{"M���}��}O�y-�����go
���z<U�~�~�A�z'����5���1���kx�Y��]փ�쮭����%Y��z���nKWy.S��N'R��W�A����Ϗ��E����7V�/�nm���gߢߢ&��}�W����g#Nnzv����>��� ����w����E�P�y�^�|�/e��L�Շ�BC^UE����@�F��iŞ���߸���j�2����^���VT]zy.�9쭡�zF��EWK�۲0]/ ���q6��#�*ab46������#w�;�\ߟ��j㏡{'�x���Nߒ������΋/�~��7\|����d���%@�L�ͳ#��k��6/���Y_�������K9��E���'�w'�W3�{��������:�l�^K؞��D�>�_���~3��>�(���tƸ��L��0r�vn��Q�Ď��}uG� �\RŋraC��e}�5��>�zԾ����d�yG��>�K�K� )o�7]���j� e�[�<+.\d�YtѨ<tQ�Α�)�i�+����Yq�.���xT��|�,|���'b���L��h�Rv��G����mQ��pJ�яaSm+��i�Jm�ZP����ګt7T8��P���Z�����g�|��K�t�	.=�b�andW�|�t��y��6'�]Ţy�{��BZ�hR�K�u�J�Bf|�K�1-ߤg�Sa�W<���Y��bC��j�
�@���⻫�����P�޺��)��Z�(+��������"����b��8��5^bk���o}�~�>�k��9�;�G�����G=w�Sp�
�ȓbj���Q�rۿ!z���$Eo��������;����Ǫ��=��蛇��
tD�B��v"�u�S�=��8q��.��~�cly�YJ��>�'�}8��*[u�=�g�������ʑR[��_���Ih���"�xdۋ�����j8�22�g����Q��3�����$xTX�W[=�s���ѵ �}	uԋ�u�Nψ�ղ�/��3��C��ddF�܇�߳}Ӏ@nW���c�,����m)-���P�BYp9�˞�Unr��ӕ�OWKȽ�Og�-���O��k��CjF�}�ؖ{�֜������~�>�� ,����3��xup�ѣe����;_������?`��5��,���D��J��<�+�3Z]8���_���~l�?d�wQ�wA�y�ڙ}�&���F�D��'I˭닫��X���v�d��#ĵ+�������tc��;��3�&�ĳ��ɞ١�9���ek����W5T�.uU��R�����㼺����}jf�;�c�/g�?���~��'���#�*�r�P��h�w�*e^�L��oY>V��W�b���0Z��-���3p���߭�g�l_��*t�x~6�#�]c�}��>��M��]���J}�v�Tv��E��0㹖�$��(��I]E�=�s��S�C�A�ױ�N���(�u<��w�e }�!T3+�d�Lg��̇�}~��C��B����֎vwnVoG���\jU�F�(eFF �W� n*��yT=��n�+.��n�o:;<�3�6�q��$��{���A��4<{�C;�a䌐��>W)��D�^�E6����-a���|uqBy�B�no=~�=;��4:#ʇ��dWg��!ŀ���L�b�F�z�e�T�d_���<���O�uE*��+>gإN���φ����޴@��{"��_�*�,�f��w��~8o׼�7�;�k�ESVla�H2棚���L����R�#º|{޳2�]{��K��m���%D��|��W�$T�0U�~����Ҹ~�'7Y��zԏ3��}dn�?ݹWu��(�)�;�uz0��N��5g��ұgKK�ռ�P�b�
s�����{������e���i���u��eƺC\p���fO5�*�b�SLC4@�ᗘ�vS�Ř��k�ܪT�)g�JV���0:�ݴ�����@K
w&���>@�,�߭�)��02��<�?����7-x	S#!�vG�`��"Y�&��?�����$�{�2|�{�=�B�C�B����t���s�b_�g� B��<�s�RU>�o.N�z9�/�3}^�#���g�+A\�CY����o4��oI��i�s� �>8�v8ڟdi����Cw���=�O���;�Z���0���IޝwP/���e7��_��nBe�Z���㙛���NӿgxWG�g�������$׻�9���)�Ǵy�:��`wd
�h�W/n�g������f�5�s�T[���5��%�^������������s�U�ex=�}T�H5o�h'�(��'�~ =����a6Gq��)l�F�}�!�:��>�S�e��@qT��5F^E�yTdw4�`ϻ�&���+���VqQ!��D�jF}�����O�W�ǌ��@�-� �3Q#�9��z.�K�Ϫ���Uxv��qK{�yn��{=y7�{=&|���_���{�#�FxC19A�C���Vr��mT`��5 8T�~&����L֝�Άk��7oZg]]Xg�ܑе�Y�����Ε��?	j�/3'��lb���uW	���a�z�+8U��We[�*sшw��f�d]I+��֟9���L�!x�o)��R�o��#�J*|fbQ}�߫~O.+޿a���~Ν�7�G��#�jk�C�p�z�?��]b'*rs;{�)�*��<���_�*Mz��^��.
ϖE�G��T���;ޣ<�ć�NB��q�%�4}R�n�j�Pt�f[���5Mِd4=����*j8�߱����>�Cj���f�ɢ���X<�����g=[�V�h`�l`4&��~�7���OB�7]�~�z~�}�l�>(�A\mP�{��������/�ncT�j@��<��?9��:\|� ��Փ��{����~^�FG��O��e�߰Pȇ��I󚍂=��H0h�w���]�T�װ�%�NO�DS�Ν���/c��N5���?]ԭ~��VG�^���' ���nD��}Q�GQ7�h䇨�T/d�p��j��B��\VzL�ѧ7=-�{���
{��v(1#di���z	n9)�=yU9�^�$l��u�Ƚ�!�.��Q��iŞ��w��5*��m��w�G���]>�]u��L���C��z�_WKȋ۲0]/ ��q=���<h��1�{�6T�?�Nh�i<��՘�^xA[��,����3���Kf�]#
o��09�����RM��KJ��Bb)u���P��̩b��Vr�-�7�k+rs�1��mq�>TX6�ۭ�S��|Y���,���E�u\nc��W{�X`_F����VU��Gz�����Wx-��AZ����mWN/P��T�`+n�c�ު��;��0:wgI�����ޓ�3�y�ݯH����[Yu�����������:+��N���q�r<���}uZ�<W>bO�%�Oz�"rO����[�[~�>[+H�r��n��H'��^\�`=��b�js�h��]��^ϺG��}�b|r=�s��
*hv�q~Al��W$�{�9C�� ]�������rp�ȯx�E�;y��CΏ8��*�{�ިR2�㌥�ׄ�=����ۗ�D�Z���.g%��!����IAߕŅ'b�F�Y~=�7���P���z�P��=�ʞ�U�W�C
���NSvdg�S�s¸�+!��4����fu-��}�<R�+��lC�q�1�;@1�{"�G��*m�.!]Cy&����q6��}�CĪ��c����z}�x�ͫ��q�����7�?MFķ��
ro�y���������oxנ�bRVlg۔���J��2�K������+`7!��W3�菣���������6����`�����`����6���l����1���6�1��8�`�����`�����`�����`���M����~cm�ncm�kcm�o�6�6���l����1��Sm�cm�M�����q������1����d�Mf��%��Ef�A@��̟\�����J��AT)T�IRT@��J�T����T����$%D�"UUHB�Q*�J��$��T��*J ��RT��D���E�%)B�̊�R%
�JD�U *B$�-�")RR�UBE$�*� �%%����������)�	R�IPJ�
������"��%
�@ ��J$P�%JD)!T
*
D"*))"���g� �p+!M�� i��j��)�U�Z�v�+�i۝NڨɌ`��ƪ���G@햲Z�wa�F��1%@�B�E �C�  Z�'���HP����ѡA�MF������Kq@ 
@9�p �4P 袊(���V4h袊4h��z.4z:4PthÌPth�GuQETJ���	*�*� k
��d�� �,�U��hkAZ�ccAOl�,J�u܆
EZL� A�5���, ҄ ���!U(���f)��[� �� T���(��{`c�U�Т��:��@U�1kQӫ��� �06]����Wr]�EH�� �P&���%I"�!�� 1�JҀ�������jSZ��F�t�h�A�*�f�:t4�4Hk�
���XK���U�hֺuJp6Zó v��@����l�m�� �v4Qf�X׸ ht�lM�@P�ݰ�
�Ԭ��C����Wmn�wn-J�+l(A���m5j�l�]:kP۠;�ݩ]��V�%DD��R�]`� ⽵Cжդ�5�@�Wc�SNt54j��tqv���͛j��n룦t�.��m�d�]����j�m��f�m(���b��	$)QA"� �Y� *�����]�0)��ҝ1�4�΁���J�i�sR��eV���i�L�V�)�(6�l+;��ku��U�*�4����QT��E ����K���C�3Rkm�h�L:j���gN�n�Ś����:]�E�5��c��԰�ʦ��+�R���E�� 1�)QEP��PZb��  Gt-��@�����! �]DV��ݎ��W@Y�Wwm��&�4�-FF���Ș톃Zncl )x �?!3*�� �Oh�JT�2�E=2'�4�� h�JUM ` S��f��� ɑ����SJ��)(�7���2����&`DTz*
���e ;�a=5�Jdg�_W�}_U}��?�_W�| ��D��TA_�����D�D���޿�?e��΍q�ˌ_����Fi_^ jX!ٲ���U�1�L���j'mLg7+ �1 7^K��Jc�)`VE�M��5Mkڅ��,VR��(4��$&��W�2� �&�� ����T�r��,��t������¢��nI1M4�
��T�`�U�SH[�	�2���bY������'�zc�n�8]�ke��e��e��t	� ����Z��2�0��Ѵ�7�#5J�m�ʫ;Q���Y[-�\�6��4�:�VA���Sr㽕u��fh�]�#1��)�D�����VPkF3l�6ɺi�0չ��U��g��f4������e�B�0�rE���B��a���" �
1�\RC5R�F�
�DM���@lK$Z�f��b�8#zӧ��E]차� S�������w�-l�%�ۧ^�2����%X��7�Y�5bͫ����%��3f# ��6��c��"����>���x`2�ٱN�	)eԼ1�)���e��e-Յ (̸�Y��ZƔ�6�Õ���hG1+Ytӈ��:)]�ki�[��V^�$#)�B��2�	��&��i:�R�uh��HL��]�])b3C�b���
�ˢDER��@ѱ6��B�ѽ�.4�[d!y*�:��
��@�­�[BԿ�m��em�o[�"�cK�Q �B����w4�A���m`�ɡ^�R�$�9���KQ�34����;
 �T�i�F�LYW���5�&�F4X[N����P�W$��7SMҒ��p67]��K�4�z˲)�/`��4����W,Jm�W�����.��3����Lb�6*
��g%і�^�XE7������M�$lZ-����m���R�[o�-�4������.�0���u4��_6��î��Z�%YNT�
�6�-���tT�`�+�R�vֵ�50цh�Tf��*�J�l�Y3e�:nf�b6$Y�^��a:),�.���}7	��o:Y���[S<�u��(��ٹ�����׳�4��Қ��Q����	̘�X�H`�ViRJ�6`��� �()3)R��U�R�mǃ�ə,D-bQ�kL
 6�Er��Kq�ЯM-N){yI;f��C&��E�@���a�ԃo�(Nj�ޫ
-v6�M��j�۽��f5y��n��QL��$����e\D[׆����:䣸��0H#0��Q�ʊS�[3q'urf�>SF�l$Dʛ�	W�4<��$%�Y6�C��t�K�`ڕ�Ы9�����0�0�#1]$�J��2o>��x�`t&�Ӄ�(�Pm�Y<ffE�E(��&AtXe�vM��C*�ʕ�QT1�ZO�*��٧E�
��@�̽6�kw*`t���7MW@:wX[T�R�YJ�#p6ŕ��j+�2n�7xAuxޏ�7�dnV����7,��g��(�ո-�Z ǋK�a�a���T.�I�m��Ш�3j��d�H�5�mm���!��a�Ղ6��dnc��%0�,��� �T5�l]�u�36�!HH��N9[L�<V�Z�j�V�1l�\�c�f���I\#*2�0Vn�T̓f��i��Q�v2��������-l�pƞn�P޼�F��ذ%sB؈˴Ԙ����}4P鎐�C��q]0���5��+��t.�[�۶�i�ĆH�ɂĚ�7PZ3l4vPnm��llfh�����+5ܡ�̢7--��P��!4IRY`�N�;��Vŗ"�7��Tp�����M�WHā2n�5���w�D`�Cf��L�Z�oE�h�B�9�p0h[��F�-��͸�u�4�M���$˽4n�CB-��ZU�<8��:B�2�|TٙkE�'`b��J6u��z���U�Yl�̔�[.],�v�4�x�u�8VT��)m���'�{L����&�ŵv�h��n�SVI�к.^�x���Z�<W��t)3gv�53W�m2�tc�ՈoZy�sN�bM,G"��bT����Y%�v^j�M�,�5Z�'d���)*�-�漅҃43#���Q��u�ֲE�щ����v���ǚ,�䣎��Vv�J��,�ב�OB��SF���1���x��)��qh��S.T������'{YBa�Y��Et���0;��DR��"n,.��P2�(eZ ��Y�-^�	�M�9�V��{��T^L�NȣP-ff��6˽O۵-]�㲦��H��7k0i���f�#M�¢�=lV���M&*�̆�E�&�,���WY�/�Z�e��SRJH��ϖk�%���j��w�%��e����͎����A�?&P�ɚ��`D�(EF��ʳ��٤H�0��qF&ޅH\ܖ
u��S��Yע��j�sV	���@���m��5�9`kn�]e�x�wXli%�-3X�],�5��.[Xr�vKǀ:Xe���`KSy%��(�Xwۋovb�.�k'�OY�I:��X�f�����Qy#�ٷ�35��R�m�+{��/BŴ�MI�H,&��k1�Mh���[�1i��Y5*X:ਛY-��8-LC\ٺmSk0֍��c��=(1R�q��ò�a���㤊��3qh�vl�����2RN�(�:⠰k��_�^m5���؉D�XC�Z� �� CcM�m�խa��[vb��{[B(n��
<��%ZԢ��L�b/~���8j �v�h#�
��Sp�ܕ�м�c�	Xu��CD��JO�3Kn�H��Z�iʆ�c�O�k$qZ
����� u$���-'����3���2%��7SV�2ؗI&�(�R�h�Nd�Gj\sh]d�f��L�9��S9�e���)��b��oD�e^i�	H���ITuP�b�w�lbF�����P�ظ(�c��dɩf"Zr�3w�S��Ud	�w5s$��^�n�϶I�P��h�A��+r���W�ŷO2��y[Ot[�tVac�DDY`��2j0����z.nH�:K��֥ �Gk1z�f;W���q��ե�֕ �̔��Iݬ��Y�M-�YA�n�-�H$���fv�9S4��%Elj3��VZ-�Ϙ7�T�e=h�u�+B�}n)�RP�a/(+��:9��c\�iJk7Jmo�˕3(�0i�.�"���g��Ռ�/~����>�V(��;����AQn2��kF����Y/e��Z�YY�����%�x��sxV9m���S��{�����Zg*4��7�n^Z;���a�k	
�!���-*�'��4M�!Iwm-�4�!ݐ�m��s������,�4-6�ąDT �r��T�v��4��;�n�&�,��I��E9O>ִ̽��)���4r,��WvECH|�-�6��(��ө��'4`��KL`���1�t&��#Pu�&�{o.����K�%�\�����b���%�Ѕk�C�:�A��<�����-�� �s(���-f% ��Hp��;�[����4�uWy�I'q^��&��(�C.��BunN*6�-Ҭ]�e9�4�M�l�Bժ��le72�sjL���&��P��y�q�D5n�H�Y�\��-$�� r�L۬Ѫ^��t˔j�� F������+7�8ݨ�34J"��V�PՈ2RWf�2��9�V�ˎ�17�+J'.��k6�!y�����e�(ʴ��fm:��� ΚT>hR, ��w�P���h��f�in,ՑrZ�^��Aa(N��e���Ղ����|ɫצ�]*@�q����Y�&FٲFd��2|�Ƶ�D��*�:��L��XC�!������T��>�v�g1�����Vw1*B�4�����u�2�,��3*зn���"	۵AmnJN���)-�2KtYшT$� ��hHn��1�Cej���Дy�4R�G1w6B,Vq.�a��2�1J%�'��j��W���*��W{�ѷb��<I�^�P1Pj�jMͦ)�0�Rz+h�۔�f��qȮ�\������m��!��J�����F���:�;���M�);4J�����G0��3.��ڕj���h��ʶ+�m�D���E�P�xbSbe9pŖ�J`��H�YRT�p5u)c{o3n��sE�!�Z�/jn���`��1�iV)����u{���m�J��+5Q�Cƃ�K���YX�G,��@	+&�ef���&Ս��07�f��;�ʡ���]�� �	�Z�Ḙ����x���y4ǻ)����j�^�J��q��+C%�^���q`M<�)S�t2�ޫٚ]��ߝ&��1�u#7��0;�0�t�SU�Ǜu4[��%���2��=6�6'�X�Ԫ=L�Rvk]Gb!��7�C��nF�+s�oTD��7
��mϰR���+�R7j�e�#hґ-Q�O0;�f
VTp7(^��Wm �wkp�¶>Sl�I�	�ʴ�a�w��]�6�&T��õPj;Y���~�k)1 ;tsf2��֪��B�Bb«=�teEN��9��^��k�$�����jo�p�A49�X���\��!�[GPR�n�ҹ�J}-��n?�`�oat�[�P6ݷ4R-���F�ɭH�n��8E��7/U��!B)0j@�)�!]�
�ܧJ�VQU�u�JZb����@���7V#իː��S]-pkӡ��m^`�^^9qH' 2���M��SfZGq3B��	.#v��T�����y��ȵf��Q�����U��Ed́Aл�ˎ�K�����\��X�hͨq���چ��1Gan�2R���83F]<h�wV\f��k�W4A��pR�w4�{��f�E�T[a��bt�C+%��Vo)��P��&���WV�S�Vd��Ԓڽ�e� �Rō��Xe6�8�+VV�h�%Z��Ȝc.^��୬;HPe��jj)���v�k��#0 �ܖV���׭���-;�SwxօmLzvm�ԥ��#[׍\��!��R%���wj�H=P=j�Ƀkc���`���
1�g\��6�u�uR6JGh�0*�v� 8�`�F:� �CV���*�l�
dՂг�/o>��: �	�ii�+���r��h�Xb��X7[͘���5*Jà5� ��٘��!�nLs:u�)��mh6*[��$�t�  �b��Z�5 �	���7�[�6ivw`�&H�IE@�KSUM�B�Y���[j�l����Rz�{0'Y�qiZD�j�('�F���	�
,�33c2��^ރ���]��m�R�Ae����q6�6i+��P!�3,m�C�YgoC��!���C1e�ȼ�j7�Z��a�j5V��FԗB#�,�jQM�M��@�E�J�%3E�C%�gr�݊��ap�11�mLtKÖғ�h���V,�h�wmA�k:/d�Ĩ�f�dikut5ib�`{+1�en]<��d; B�Q6�#n�.�+4�ڈq#7Dw��K�q�{U2Zۦ���wsm�.�!�'�����E3z�P,�L��5��^d$M��������z'��$\�B����B�Y�����s�{D�3�"ճ�ءFU�+.U�xQa�� �e�
p"Ќm@�ʬp=+:Ӻ%h�������l7�b�kʏ�yJ=����D�cM ��1����v�U�-�Cv�
,�[��]c1�Xh�2jK36
�ǟM7���I�����+��,��7z�1��gv ���D��܊1W[�7q�(46V�2=���,'w5+�1�*Xʁ<Up�ڨQ�Um\��Emԩ`XDR<���,�իt[$�����J���;�!��7a�`�b��l2���I\m�L��*�(d����(�
KW��A�� ��D�QM�L�gK8�r7q$!�8�e����b+�U�*89r�K.Z�
`�W-������RBcR`���v�f0�- �S��)�l��6�����
��(��$r�֔�yK)IXr�	����^d��7q�HA{E�u�
�5��v���q�5��/0�+hR�S"z�͌�ӛOsP�B�,'��B�-e����]Ksi�H�e��v����FIw��b��;C%�H�1-.����u��+F*Y�m�ɐ5[I���)��L�fVʽ�t��X�b�mzIf��Vc��K�/+��69J����æ�h����˺��J�h圤�d�B)�����Aк;+0��LReۘel,��*z�I��x�fY9�-�F%h�b����E4 �d:	�jY���b@ݽ�pM��ڗQ4�I�B;�C	�*��+��bzE�P8���YEӔK�7K��J8>�ݍ&L����y%��ś[���ؔ�%�RELm,62��I
r2t4Y�[�*w��@Gy7@�Gu��6͉xl%r��G	`=ղ$�/�,M��6��s2�ڑ�������B�9���ɦc���t%��ۻ�B��J� �A46�U���:jܷ2��5/�MV�蠎��>m��tH 1^��-9{jkj�!�D�|i�X�
Zz���(d0i���.�ո^SX�E'�%�P+q�6��-��uV�@�Y�eE�9Ql��b$L.R �T��� ���=���@�ӗcrU&�Q�ba�5%����p��x�WZ�J���IV;����MӾ�8_wW`kZ,�ՔKefI�*���XW�n��@�,��"��4�*H*m�L��U#'�z�f�̼ѫ(M��T�5z�i"�.�\Yp)[�N榋f�ͫ�$�[��!���uX��!��7ʼS^cfgI�����A���%m��}�{9T��V��L�S��y�us�Au0ݴ��;�9$Rġ��N�}�����5m��9Z�+@V��r��&-����.bı��&.̭�r��\Fh�)t=[�nX,J
fU�L{y�B�{Ɖ;5�|�����X��^��׃S���B��<������
�
R�y�9FCgJೇdS0���T�kΣm�vdv�s��h�uϪ.�hww[�V�'!����qrt�:�@��땦����J���ypQ �L[4^.wX�2��;�������lU�ӭҳ�a5E�K�ܼ��M�����,
�'9��"j`����{y�Ņ��IiԹͧt�ٮcx��k��|-(ܷ�ܭя Vxd]4��$���{��w[PjM t���J՛C4��v!���̼�.*'��Mf'u"f��r!kn�ߥ�NJ�����i���r'O4�oa�o�aC4w��S���N��t��"H��]M��s��:`f*9�z,��V�E�MU�pZ*��e���}G��PL��GS�=rg.n�=E��t8G1xm�[7A5cH�w���X����G�/����Gt�&,R�b��t��Z���4z�o �+�#�N�5գ���W� ���RZ�Љ��L[�փ�m�8)� F�B��&j�����W�.[;�b�wT��D���&GF��(�5��2���V�e�!��H�R5gA�hMt����S���*C�5X�_=Ȝ�wʦ5k�ԥ]ui�	P��ӀSו�'V��P�yŹ�?���쏧�>7��Z�F��N�|1T������gS��M�k8�}��+&dP�(gE��ސ���,'���vFk|�&vQ��k��< �d�ã'�\fW,=Q�2���݉8B;F��TKV.ܦm�v�5�e�����B}G���:��5fT��w(���OrڬBN�@����	-��qJՋ�F0����M]]Z�3���bOժ���$Ĳ�[��4o��r}t	�m���ǨNo��{�L�Պ���OPw������V�T�Z�ޤ�g�Ud	��ս�RO:\��R=�Ny&���-{�F�n�ܻ��X���c���Ł*y+��᯷�^�Ef���j�&��7�{r���B�c���_kf�[^vH�	�'��+
�:�X�b�J������EC�Ņǚe\��6�З�3����6��	��5���ĝ��.nQ��n�U�����ʰcO�`��}{BR���z�>9�jc{��[�D+C4Ԭ��o��BVE�����Ǭ䝜-�J�O���ژ:N��:��:��c�.�(tU�����1�u	ӯ�����T8��!z��5H��T��Y{�k��U�qR�P�З��۸����a�'p�qsb��l�M�4_|�=���d0%�E;���;3m!%>�ﺢ��
��Nx�ƁcoMn;o9���=d"�iN��J�<�Ň�Ր��7���(�W+\�ݐv�~����npgM�����Mϔ�r�Q�N��#���[9�+ݼk�>�`C���Y�{Y���{k5җ}n���u�Ө{����ZE�]8��i��;��M2���*{�ҝ�����܏J:����/�ˮ|�}i�\�C٤�no�eZVbu} )t�Nަ�l\��9����]�D볭b�	��v��y�C���Cv�y�4;z�w�۽��h��gmՊ�G�������B�1">]�s��hb�4	��J��[r�WScL�ֹ��"�:�H�v�d�B�
e�e�*���cE^��*��LGt%#�����8��n%+/e�e�ùN�Z��[�^�r���f"����y����]��a��E�u�$�y�<�^up�����_DM[��R"[�Xori���ȥ�V�n���0X,f�[k)R�{,��Y����a=|&�S���,��[��VfjtƬձ���Pqe���7m�q؂�{�m���_�j����uo8h3v�-��Ļ��"�Y�L�k�1=��[{��*"��e���Y��Z��rƩ&��M�Sc$mO7y�&nKg-���Mq��*�V��qְ�WV��'`p\Y�XK��6����4���靉ԌH���[����37.e��l��s�ZP�i�6eM�ܕujšJ��#�7х��C�bs*�/6dT�i7��!�|;�%��N�>ffݮ��lwer��'o�GxI�.jӸ�k4�V�lR�yJo
V"�q'j���T9�[�-�5���TV���k��7Rv����h;��*���;8A�EA�hf����FL�QӖG<"�z8
���+MaT��ow-p��n|�wȗE��k2�Hс����M�CҖ;�V&��ާ�{���׹����u>8Y���� �q[m㑗�.��@�Z�ҫ���ȼ&M��\j%��x��Q�����>�5��:�Z"�!��Zћ�m�,ט����$q��L����^�q�C�/��Db���
�2\u�nf&c�j���*oh����ko����ʝ�7Qَ����}�Rt����u��+z	��u��>�t�ʴ�3�����0E�Ka-��3��4�b�c"��du��:�1�J�jјeq��� s�Lf+\����#c]�'CK�Wu\���혓�iO���-�)d�*��}Q�<�*�{�;{��,V�(u$�èj2x&��2��o:�V$N�j�\��"����r���j�ޕ�69�+�K�0=ʉq��l�t9wXB��
;�y�y��W���X���]��ɱ��,���Д��CZ�j��lM��A��(��nm%|0�O�$9WJxMZ ��#��$e�\Z\|��A�(��=Uuk^��>�5}��N��)��۝t�ޝ���#5��N�v>�y�nypbΙ�1�ތ�J�XC����s \e�Ù)�0� /��v�]����V}j��̖Ŏ�%��;NSv�.�R�6�n��$��<Z�ZpU������ƅ�:�bZɼߕ�:t��@[�6E�u�-���E��7������|�XC��UE�y��0�u�[]W��5)Cӕ�>a� �����ޭ
t�M�h,���<<a���x�6r�2���[ᤫ�X/���(���l�Ž�dX�{���/�"6��`��.���ni����ꅄ.۹�u���i	����ݮΛ���7��I�.��X�����eԏ �+6�Yv�7$Օy�]X�\D��f#i-�3��N6r�Z�N�_�!z��w�8��C�阋Ee���-��]����kFu��}��Pp"��w='h U�c3�R����:�U2���:���w���:-�5�x�E"̂��uwW���Qu�CVíW��f:��9ef�5���`=����c�nG��Qk:O3�v�lF�N�=5"xs]���i�,�e^fgs�eiz9j;�1@����OLx��Y���]�̮x!��K[}�xV��Cn�O���h�́ܯΎ%��S��in�9�]`���J��U��Lν�� ����"g7�|����'KWX�,��Ciwv\����y��(��8�s���mʔ<��N;c�vÒWc7X��܍�-����pVrf^�;�n��,dt�?�i�S]��h�ҕ�gOL">�T��d+�t&�I��YU"�:�}0�6ub�z{��.L�8�b��V���Yv�D�f��l�)h��)���r�XN���1Vw�fEܘ�21�h�����y��o��f�`�F�}���-�K$�o��`�o���L���1�����B�c��B�é��v;U���^jd�Dn"xuE��ی�%�/�Uϖ��%���c���-��~_�`�A�OiI��k�eJ���`��#��#|�JN.
Rt:���|��z�m���p��;Gx�*:�*�ѷdRΉ���bZtS|�#��3G�dkRyug  ����U��%x�Yot�	���N)�/�(z�v���+���!�i)r��m憲��;��/L�2�s]��Ө�_�i�α���#V�	eAw�6��7]�eތ$i��V�kd��S2;�̎neEb,,�6��Uv�"\ڈ�]�ۺJp���^r���Sg�q��b��T�Mhێ�R��Z+6�ӱ6fTw��;V��5S	��ᐫ���ψ���(��A±\w1j[���'��L����۶�m��:i���V�f�0�wu� �w4\�3V�#<w��V�\�OJ�C��0�<r�������I	eA���[�{��]w���>ޖ�
}Fpe>}֔�e��Kx��p���vp��QO�v��h5,`�yN˽��#���ܼΨ)C��weA�6`Q[R�����o��>�r�����2	l4gA}�m�EKh��ɮ�N��}][�R�#�Eo]]v��[��eF�Х��c!�y��NEF�E�Ǯ��&�n��XZ�a�Or�lb��(��g���k\�u\,����G�f�DUvs>��qA��Ok���+��-<���X��@�8Wq�u�O�v����nƓ4ǩs;�:_w]3O7_Ǉ`���Ϛ/&%y�r]�3>ϔ̝c�w����#H=�Ytp�K�S�[n��$7��.�&�ݫ�����\:��Ն�������1,��Us[���\{1v����_j/����"b�)^>#OS�	�\7!ɢ�����j�rM�q
��9!�uv��zHC�:mM:���ư�L��w�����ԇY�ba�5�fw>d4bބ���#@�GT�Q�7�k���
���hm!ۘ#�秅�4����9�X��n���EI��=6��)���%�c��`��%��ڃ�+�Un;������5�-��P]]��"��:�ir�����SQҒ�����4�ê�ߩ:��y�<�@�����=&�7�7��Պf՛h��,�VG*F�R�w
+.��*� .l��7��)a}B�ngP����҇z�a�z�a �}�!ׂ��(�Ӱ!�j�8������n�,�PHj��S��i:���;MrLv�,�G�����VQ�؍\�2�}J�j��u]����F5%h����Wݎ���V�jqqV���eq��ec��o=:��.�/�;��7��24��BH������3V�Î'�jM��&/N2�EN�s4�n�(��.�a�=��9���^ڝtyR��]��,��ۂ�j3k)ǜ%�r�����/S���3z�Ӵ�vIr�K��ػj��* :�!;^*Y�$̶>K�m�y��t�u:��"��.R�S�n����,�'_�`���ةMo0LMFp+j��]:^2xa�Wv��`�TO:�v^>O7�G���Y�d�7y9h�e��fv�1k�Cn��	��N��|�^��]�9r�V�-��<G�(nQ�e�{}`pۓ��<�jl[j�d[�S�r�v�Ѵ�pZ��5q/;2�s�oa<5+f]�©2�1[Ր�*�!��UF�ַ�.u3�"�hi�җ9{�PwYO3�$���]��=���@Lݚ�3���Y7��,�7aض7tb�T���{NS��5����E�o-��)&:0�;7t��̲�N�Jp�ⷧ�����}u��g�*9=Ha�c���V��m��(�n��X�ױ6 �Cu��Cag���vZ��mL뮭/$��z�?gbi:t��M4�\l78\�wJ��fl��<��܄>��M��U��J�4���n�S�ܤ�v̷[2l���{�p��W.��ǆi�lo ��l����H��7���H��#EA�)�e��Cq����� ��T	KF%L+�� A��]k3E���e7[�jw1����<�z�T��}Z]�Q��`J�a4ͪ�-�8d�D�[��Zq��7�nS�*�7�u3�QM|P�f^xN��oFC�:����E��v���As۝5�f�孴��K@���=1q�n�Ei]C�kn��_{ݖ_{�4n�կz��h��ٲ�]���^lUb��]��\gcέ�����:�R�:�&������/Z�+<[}A,VE;
1c��Bf��mr��p�P�e7x���{%��M@b8��_t�\P�w����.�DX�A��QWy��'����Efڦ�/gs�c�.7�oj����n�od(�^*��r2��ʋu"������0���GwW5*�[���l���yƟ��<�/1�Ν#��a`�F����;��������4�^���댤��s���/�g9S�Q��M�o6���z+J�¯:�-�l
�"�Ǎ?�-�V��_!5�$�͇]s��FQ㫑U6�#��f�ɤt��[��,���$wsCW�,Q動�l���J�PҬ��]*s�>J�f�e5p�m����͵R�[��:q�
��=��%&4�z��tv̩Hh��0�7`�_u����Ы�k^�1�J��C���g2�o�y�;���c}���[�q�����+�.�f�L�w ��i"��.�Wd�����A�K���wˮ���fݺGw��X�����@B�3�/���f�Iٕ�@��s���̣����ђ�]�[YN'u�gZ�i�0���|F����{�\�J�bZ:D0���<�6�=ǋ���{Χ(�L;�j�o\�F�w ɵҹ�Z�_v�1�N�p	��L��`�en�h���{Ԁ	a�w��B�{�\zijRz�-^�8V>�˚���r�\rL��e[�����~�#�l�b����H4���,+��z=*u��2�ם��i���ass9ՠ�2�L��[ծV��(_ʜ�RKƫ;S�!o+Ѽ���Jܶ�\�:��:�R����x�2thwS+��,�n㓩1>뱯�~���"�
)�Q{�u��߽���_����IN�f�.)(�9�����;Y53�(V-D�V+�]L@Nt�7SM��,5i�v`�j<�7T�"�v�"���D�A�c�:�_9+h��X�MJ�[Y�[��{6��om?��l�S�C��Ge�.^�mn��F��{��;`k���Ln��;A}Yڍ���Թ]EKׇO9��t�/�>��B}:��`ܦ�-�+)�����a�$Q�=[��%���cn��r��7����.�Т�kwlu͔�A*�a�2��2�v�c�':`�����Ojm��]������D��d�!ɋE�pl`�Xv.S��{���]��s�V�wܷ)Y���<Iv]��-�ѷ[��B?���t�J�7X����+���'K���M�ϸna������F���2>���:g{�Y��@W;�Q�t�돛�����J6�Pt� V� ���Ʋ5�:t��B���퇹/�˙\	���ѓ@���6;4ʷN}n�IL5��]#[�9�'�ޓ*�n�Ȭ�*��jKmKPVTiw,X���f�EO��]6˦�`F��ɪĽ/�٢�[�/��9:��m�R]�+�U��o<�:����[#EYy7��J��ܗ�1k-�� 1Mxu���$�Β���݃���o��-���ÈI�KoN�*��G��%MK�q�7�ٻ�..N}aꗴ��{�W�>���Hbա�jee���d�ˠI�KK-�+%����c�Î�g��v�RPR�_r"��;�'f:�r�n��	����2�k�_B^Cy��.�X]���������42,���n��B�π�*��R�]��-��
�����tf�
�4�Y�x���0,i��o`q8.,��3oN�Y�a�Ԫyϯ���r�!ű\�ӈ�n9y��t��t���p�K�.�H|�)�S�.����1hrG���U���P�й{�P��"ćM$��Ɯ�n������s2�;٥<�%<'f\ܖd�kN�֦C'V(�z>��e��F�k!'�]��=�RղK�Ϭ��Z�ō)H����`�����C`c�R�Z���Gq�}0�/r]2����xoe���+�oD*
�ۜ�J�lH�u��j+4(��ɇ@��C:wKw�ػ�o�X�1)Ӆ�����{M��n'g\{3z�|k,���������rlk7-R�s��[�
�Y�)�Z��L�v1��B�њ��=ܖ{U=� '%=X_b��+���,+GE4�ȝWl��ێ˩�5^'l�~g�{S'g��¯��ڝ.�!}�%e5����޳8Vme�`G,�9(�vW#D#w�c��YC�55*�͖�j7�u��:6�(X�R���uו�Bq�xu�ܮ�@�{�j��uk9R�����g2:�Q�2ep*AW̋"&n�����	 ��uEr�ⵗ����(L�:�ko{��z��*��"�(,�6�#�fg_wٓ��Qujv�R��lm��M��o�#��-�\�j]��>�٧�1����t����O�����t�)@��wܮ�Y958N�,e79��uww��A��Ƀ.�Wa�@�
�ΨS�Q0k\��`٪����42��۩b�6��W�f>�U+b�)�y�z(��M�1$7�oV�v^ �����R���0�^q����@�èk�.�)�¬'ZL�G�f��olyL�guȞ�	Ū���P��^X�]���f+.�{��	�\w1�e֠��]F�5�-�oj�FX|���6���������U����_,Z����x�Ӣe
�Č�}�����Ը��b�=��Aep��أ>-Tl�3��s�+���ʬ&��RD�F>�V*�Gbs7��P��4�g����$XE��4�k{�]���;(Z[]H9�j� >�`q�������ʢ�n�a��j�ɱ(���en:S,��|����O'�w���-;��: XiC�u�p�+�ih�d�x��꼶O�l��5u�9#�	E�亮�X���M�]8ا�.'�0�2!RK�Lۻ�,A���@NB�dV
�nj�o��׹܉�pd=wJՙQ�WQq��by�;�V#�����H�pA�9�'7�M���2@V�)o>�GY�ܳ8u��<��mN��ٷ�Lf_G�}z�N�U+v�*�%С�![����:ME>��V����c`4i\��o��S�@�D�����U�ܨպ��6�$iRl5F��wO�t=��m�U6�wpڄ�
�\�5�>
�0���=Z�	��v�W���:�L]3v4C`�FT[ϔ�#.=1A5윇ԫz�t�K;���P�x���I޷�����Bmq�I���cc2���u�i�/{�	i�/��7�}�;�E�CL�mq/��H�z �����$��:����oA�U�f�V�/���
�+(X�^�UҤy<��']^���mLv����],7l����Â#��4�:�N��N]���K
�DZ$��8p��kꗉD=y���E�<�P���E+|��{K�#�M�{,V��fb�
9;lp���O�[�$�rI(�C.:xfk�D� �t ��ݥ�M�}���"��Wg���u&��זu"s�2���t�WX�E�OwW��"�1��n�G*��^h��A��G0���@T��Z���Wdok.�g!����%\�68JeS�N��!Yo�wWv8�s��,M���tu}�+i����
�a�2�dc���U$Ț�FQ��;\�X���R�k'�b��"��8k;V5I�5CW${�;����z5IN}����v;˺U�ţG�mc���8R��y�)�{�\��D�U��.���6)^����Tۃ���U�c�}*ƻq��A���RgL�ԝnކ�ס<��r�P���2Wb���°�y9�]W�^���+5��R=��+[⯚Q]�j��0H�VNc�t|cd!�������i�W�-g%ףC�|�%�TT~���)��E'��jW��x�3tn���K��d�ذ��l�g;U�-A�t��{ky)&9��g	u�P�MF{�CCM8�J�Ƭ��:ڼE��"�v�NS���s�D�g����k#<U��S[������m0c�ѬP7�����4h� NQ��Si��G��^�欎.2Q���wq��|-�⯴:?:�k�ۻ���p
=�C���L�pr�TƖơ���hr[y�\�9E��M�جL�"�w)khO��J4��X��y>�!�[��4*�z�9�J+�Z�����j���ڠWn"p:4h^nv����\K�����:����9�q�
p��7���V���Z͚7�����mn_5�R�@�$���s��ۋC�����d+ \�M!�e^�N����)}������W��9&�������t�^�#∬�r ,�&����κܫ�O���h��%�@2k�Em� ؤ����,n��e\�r[�i<<J��X��}�9j�N��LD�ES#�i	r�`�Tw�V(����܋
�:�v��Q�s��[�;{I#�b�a��^ΖaU�u<�y�VL��犝�.tʭ�Z�EZ�]|`v��6�<�hҲ^d$V�G�5[��K��3���N*��\kD&�*d�q��Y��Б�n�3/%7�pM�Ւ�
�X�}>�޺
�LɍVuc��h�}���>ݭK�8s��8B|��v�JU��+�Q�%��-��)����NHfG ޾�Av�G�`O2�)�����VpE�P������]��\�o�K��$͗zSCV���6b����@n�۴�}�
$*U΋a�Ch�\��E'��-Ҳ`Z+Q�|h�ЫE�f^���%����u!�(>v�j]k���i2�d����HIt�o5(�YK8�$gJ�WJ��\�<87ۡ�����9%[[���g-���hB�ۻ�FrØ�p�Ѓ;�{2���M�t��9V�e1'j�Kܙ�2�=�̪ɘ)��h񋭫�����A.����͞v,��2S�N��J�ҳa�Z�Ѭ}/�/6���M�I���}�����<jv%�ok� ݛ�R������鲱�o�.!}�U��U���W�M�CK�	-�&KJ��Qe������[\�5�W���̅�gv����i��Z���C�Y�Ú�qUb����
un�,]5�9��C�.�h���we�f�����g	�Ψ�&�&#}�(q�PMZv�-V���Y�hvN�ξ�_�tŔ��v��d^��KP�ǽkV޻̣��1��f`{R������E���+|p���d�ط��(���5�el偮��F��R��Np�{�b�z�ьw0[��қ�����Z�t�nAEܽ#�yU�VF�,)[�DټQ*�we�Egc����0h��<�.�&أhIm<���
��/�LY�5v�}�jko{��@1\�juӕf��;�}��'��V�Q��n�D6�"�zdx�Ơ���p�͌RL	�OoMX�[R�};�c�˖�v�������X��'$2��kܣ�7Y[q�V\���X�h6�t'X4bmp���.��(z��O^��WWP���%Ϩ�Eki�.xD�B���产KW�^�w~���؆ւ��ʅ8���n�G4[�m�Cl�V�=�hJ���]�k�-�TT{i��vއ�I�,i�g����_f�jon䋒���%�J��t=��R��A2_(���v��PDe�Z+-E��A�'f%�]/e�L��j�C19Q�VZ��K��e�O"�T�*#O��d��R�@[�����&�6#�����w 
vV�^�u[.�ݑp�Ҩ���E�[�i��h���S��D�EkvT���[4=� ;ϫZV�I����:�%�β��vG�G��#b��9�p��.uꇐ���wS]��u�Y�j8�b�k5\�e5L4�傢���z��+%�I��TYbV]���-Y�ct*GK�y��z��{���u�gd]H���"��En!E��׎�ܻ{im���tѫ3h��˩��qK��ĚX��cEnc��ۼf���$�}Oz�Yl\���ƍ���V;r�lv>����+:�fl�vtH��
�.��	��®���G887�dִ9�<Z���=�yi�<�S���L}L9)��-T�Pv°X�<��$��u���qQ�D�נ�L]���J������pD��ro��t����J�������42�̰��gKȦ�j��&�I�fR�� ���J��&�Ӆ�*�l��_U�r��\���hm<Ÿ�%��P�����շW�Kki��2d��:W�4}��|�B7��l����,�WA�rZ���q�Ɋ@� [	V�3�D��X��x�����t�|3���_&�4�		V��ZE�J��h���cr!N�T����E�C0�������"W���tU��_4:Ẑ�����lH�SB*lJ�뫩VZ����l�����W��}yF

g� ���o��bCi�\��Y�xV�,C�	����U*��C��3tD�O�����&12�GA��9,]�m�e��o;��m��:�|(�Wvɥc뾼[AM��:mKz�l�S�q"���h���h X��ĳhΜ\�u��->��9V7����]+N�>W�1���˹v�\аU�}|���������<��m:Z2�"݅]q3�h�.����u�~��7s�5֖��[苒_Bm'Vs09K�2֨&J6����K�Q�Gye��+����@k��CT�{q�tNl�'�_#�r��N��7ǁ��@���GzåD�۽:�9C�������t0#�f'�0VGۋ ���n�@|�F��q�ٝW"]k��f� ػM�%R�v�)'vZ��L9���&�{����l]����������u��q(�\��`�8Cq#����a<0g5�ݾ2�9r�C�H�'�U�]+�j�e�[���7�2�n��J����O�ּ���]M ue��v
u�M�ʷ��蕣��� %+yǴ����˴��qe>�;N�	�VEQ�Y��bc.-�.��pb�Fi36\{43v��X�yp͈F�a�!�:t
4YZ�v20q��]2�5̫����݈��vʿ�s�6*	ʚ�=wL�c&v+ۥy*ڰR!�vK��U3�lMYlqׂ�F�K�H��=}ĤiǦ����Uua�1uk j%�����w:��)��\u�M��u��ʃ��ޠ��l��K���ue�K�v͓s�7{�vC5ͬM��B��p좱�d�@s�\�nK�e�5��(@�����v&�#��j+�q�ݫ��oZJ��*[�sN`��s>3�� �j�,xދ#�3u�}(يt�T�^p�#��|���� `2�EÌ�+�]�B�z~�\�U��o.���:�U��1wH�̖J�t��� :b�׌t�wY�-kx)&�J��㺹zE�層{N�m����K�ۛw%�[f�n����ǽid�o�,�vV3��<��±HC|ws�x2
�R�ҥ񧎝)���G+2�G.=:�z��֓�+������ګ��uʶ���o������R}� �hUC�$���v���X�& �&�����r���Du���Y���Nf�0���Y��b�I�W�wu[�;�wf$z�Ae�bT
��9����W06�\���G��n�a�#���cT�
����fN�Q��FZ�(��|���]�j�n�Hr0�'r�CHyR�x%��:=�t;�t˽Pu���$�c@�ɧ��[�]b���4`{��Pf��ŵ�W	P�T���y��6��_䀧��`�.��H'���J��*�
ҷ��J�L��{nЗ��1|�g�a�,S���z+����uy�I\ۦs*V�U �.�-�B�m9u9�4�z�������߾��MJAl[���m��O��٫���Γ��{���7�[���}�#2��v�l�F��)[Nw�'e��|0=s̨�ۤ<Ӌ;є���v�',��g!����S=��=&;5����͸��s�:�.c�\v���Q:{jN�����U����e5Û� .p�G]��@�J�J=�o&�;��a��sD�n�v�.L=���+s���=U���v_L���A����0�Opp�Ӈa�4p�F,��EX������]O\�ir�j̃K8�)�]�*uҹ����N�k�W������9o.�%�Z��u�Zq���.LNv7Zk����qn �Sa7���a���u�B��W*Y�+�HG)�&�X5�!���P��V�rr���1n���K7Y���>u�����l�"*���8�%�K_W,/��H��E\Y��p#z��5eVN{���P/��D�%@��"&�kw�����If�D�9�3yQbUҮ���t8�ڒ5Y��=l10; �ki|�r�j���,	�����,`��^��Z7F�ZV�A�\��O]�<8�|��\��ժ�9۽����:�V��8��y�uꮶٸ��,�_fb������ۚn�w�vNO��eI�=VN��l��S�_;�\�Ć��,ޮ��{D�-vj��!��댽�Ԭ�-*��
���}M�C���;R�=�T�����б20�������'!��$Ȭ��3�r2V�3 ��(2�!hr(*�$2i�"
	� �!h2Zhs0k ʂ����0̋(��p���3��Ƞ��r*!�� ɬ���,���!�3
f,�3��L(�#$�b��#*�2����(���'(��"��&��*�����$�$����(0�L�� ���3(�����Jr¡ʇ$�Ȣ(�ɠ����* ������l�ȳ �����
"2L�p����#*l��ʒ� k3!i(r1�)2�32���!���Z,³1�r�L��2ɪ1�� �)ɤ³��0 ���C���3(��!2�� ����I������
",�����M�,�o�@��/�h,�_}����hR'y��E	���D�錵���8~E�ڀТSx�`��L�ۿ��*�wF����}�oX�S��<U�a���D�,�U3��o���/[��n�"��=��	��'ڃ�9pw��Wl��2��*,!=�yi!CY�I�5���>��m-��z�n�ߏ[�� ϟQy[���V^��%����J��*��ӣ�֟R�u���.*{�~��?��+U��wT���vz-���3>������u]�]����Zo���f�ytrM�ż{��i�:�6�#�0�3&z-�b����>��NN���:�S6�o�x=�N�o�csn��_+>�C�Y�������q@g�0)�^x�:����qw1cp{�4�m_&��Y1�O�-b5��-��X��ϥe��o���{���K0^�=����09vG�=���&w-�yX���4�|ˬ������7D��&P��>��W�����>�"Y���g7����n�'\=����*S����S6c��ɻ���H���)C���e@}�i���bu53K9��㯑"�kVV��(�nة%j�Z��%�p�3����W3�?���SCi��}�F^^�,0UXP'~b���:�M�Z�Y��h�ku��ŭ����}�뙯W-cw9����J���I2n�9}ϩ@�LWe��v����i��]�s9�x&�VT�r��n�G*�I���>�V\��|mi�f
��C�L!��S1+iE}7��.uC�a�M�j�ֽ}"n��F�n<�x�a�6�h�q��Ih�i
�K���_����-fױ���\��i����LP�j��a�r���֫]H�`�.,������{-���k���[fx�v�O��jt��������Z�P�$�h�(���yR�;ڢj��y.��y0�s�F��Nw��~�;�]3N�:fK�9�O[Ň�Ⱦ�y���ƫy�/��yL�C�޶�8&�M�,k���T���(o�Ϧ\;���V�;���	����ܿU�����j�H����_o�xN��g�&
6��?}�����b�"�๞�H}+�`u�����cc���"��xg���B;Pvr/�w҉#�݋��\�+��3_��(��u�-��]_Ap:����旅�Z6}�
b�&�xe]�Kw7.'�kj�6��٤�Z`��I>��9C�rW�Լ#�����/�4u���W����Y.�*:�j�"���S�YI�;2�bi��U�U1_Q�7n�5���<�v���|)�X��͎M��(";3����N۽�]0Ժ�z���L��<��]/�Y��W9V�+�՛Ɯ��X�i(��鴺��9j}\H�؃��o�ߓ;���C�L&�;�(���[���Kg�v�;�tX��\h*β��*f����U+�S��r�܆��\�~��C��{={n��qiym6����d��V���XW�I��苡f=5g����,j��;�9��٘��/|�/S\���w>�ީ{3���o��bu�a��Lt���JP�W�AB�a����&�ϝ��盵�Û�^r�]����y@cP�]D���{��Ғ���t{)���`^ q{���i�����^��3��<�a��L��oWt=��m��U���R%_</�M�̤�%��#���1��Y�U>H�8ОY6���w�`P�,9����&*#M �$�{�݉�ܽۯ���msm\�R�K�C�ܹ��T#:u�B߯yY�ḇR�e#��H�6�U�eU��ܒ��~�<	<Ӕ(t��֙����g�6��9�2���7��x_�UN��&�%�;���Y0��a�y�I�G�������x��^�(Wxߩ�߮�T��qm���+O�{q�M5}.�t�]�t0tFm��Q�����޸FS�.�A+��lY!�u����VI�o�v��N�^ي��&��m��n�g1E����jM��"��ݧS�&ӱJ��8��c\v���y�N�qݝv�2�q��1��2S#�>�D+��O
���i�I�b��Ԭ�v������:��(�*qc=]��J������Ɯ�JV�9Bj��P��ItH�^+���g<0B�����/_��k���Xp�t��/>�탎Q#A�,N��޴�<�;�x[�q/W���>\�[�ռ��e;���K=o��Ńz]o�M�:�I�҉�����3Y����y��d��OZ�H|�k{i3KO�m$���k�G�����4o�<G>�ԇ�r���l�p�~S�L�^��uc �����%�~�y�{s5��0��E���������#,�=�NfF��%5���mC�������>��ᒒᄺ�^zߨm<Z�x+*��G�1���+�}�=f�_{��6g�)�e��6YS�k����c~=�|�!��ԍ�t|��'���G:��L����9x��5z ��+��1��|�\Itv��ϗ��k�y�|T����#�MH�}6�s�O�M��,��S3e�C
4��,/fi��zT2y����I�9$�Z�)�*��ΰ����̬�2�,3�+*��f���7���3散LV��]nFV��3P=ѵ\��c�/8��ͷ��Ҙk��lO+G�9�K�#Ȼ��^� �˂p�6m��u^��{7�F���u��&;���zd�	�Py6`k{���9P��zf;�������B!c�P��7�yk������K�o��2��t��~k��#�zw+������D^�k�s�����Q�k��2xw�S=��%��r�=M�9�$�ɝw����}�a�����s�ÞU���8����_3��f��=���o&K��Ӳ�ƀ]:�*OVz\����=��Ͻ�fvv�a�ǑWn%��.l�=�k��7���__s���l�������f�|{�d�#�1n�I�o؉�f��jF{֩��q�zhxf��*:����ûfg�З�T����O<��v��n��tн��ֽ�9�au�:�̘�ݷ3�4̌n����ʷ�Z�|����;>�Y�-^چ�oЯh�G9����o�h{�0�m}ݼ9�*�u���<��:d�k0�߹k�l0�~g�G0hYKV���&�+���i�OM�C����c�g!�>Ck��
1�qn��gS�/���9�kX�IW�|�j�@�|�t��e���>�)��Nd\�xG���k�zyv�OS���߼�vk�޲�����
ݡ��[y�ʞ����r=t��՜�d�V'߂�����g�c7�M�o��V{��p���2�F���)�ꨦ�'aP{���*����z9�Rb�5S�{�{cf���_6���4�/W_�񯭅�dx�m��1�=�ۥ�������z��[Kς���7��V��~;h,S��~2<d�%�3�����Ls5�{��S��`�ܷ֬�||X���ik����Sdlt��x%�������7�����*gl�s�g�ۖu��(떇4e����`S��Z���y>�񼓶���ۏ+ws�(��g�"$e�=�ܪ�}[�Dc����~ֽ�z{���^�3���x�FS��Q[���t��"o��.��=0t��'7������Pbwf����Slo��裠���O�R��p��o����˯#�路�w��S�,R%jۿ�(,����ݛc۟�o�Ӭ����F���E��hgZ���!2���|�_k��yw1�G���>����.����迶�\B�wï\g�,y�}��l���0J�[	Ϋ��������-̎��&m�~3Jۨ�ԧ�y�{r3Z,76Z�	Z�e���L������p����!d&��]�t��k�m��z#9��qމ��3��*{6g�מv��s]��ޏ|�G��q���NF}_z�X�8�h�Jɗ|3���8���3�?W-�}D�<����K}�s�ɏN}�v��ٯ�h�d�Z1���)�vz��m��ޅ�5˃6�X�/|�7/����77Ք�S�`c�JY;���ȵ���h}�������b�{d+\�R���~��{1mL�[��m��\���3�~^�i����f1�.�h�����Ŧ�WE��M��=�����2��4ϓ�Kbc��@[�{�/EO_>[s9�>�z}��G:sQ������Gp��au17�o�10�?g]�*��|�XZ8N�]#��h�2���\R^�X�K���Qa����0e��ה̙�c�(�k�����i���w�
pYz�� ɼ�æ�Hw��Yzz�J���[���5a�N�`��eC6 ������\,���s;�5��y���V�cz�]{RL��e9� 齘<��Y�twi���kۗ�{m.�]� �B��\𮮱����z^rs3��'�W,�ԩv�T�;����z��0`<�΅�;�����!�{ޜsӆ��v.�}z��~x���w���.|C�|[϶yI篅;�"wMݮ�R�{�;^�u��Ԙ|�g�Ӫ������$罐���o5�{���P~���J����$5����d����^��X�<��9�*s}�o��F���hs������U�_s\�`A�=EfoR���������0��)����~��;�,8��Fk=�=�������7�<8�G�ا��wy-����4�}�~����e��)�ڜ�����JYKTڄO?�[uG��|����?U�M��ު�O1{|J��피�	q@fy������++�N��Ayu��/X��O5�#d�9�Ɗ׵�Q�Ddl�b��%����U�c�����Z�YT�Tڑ�O19G�s��V+%�$ف���e��}j��g�f���3s3��Rg-j���u�ǌm}�sj�~ԭ�j�[�9^o�*�A�)}�6w��L��y�Y� u/9�X�&�<��?Uv:7��X�@�G� ?�9�ִm�`�=�p������N[�Q�s�վ~f��%�Җ���E���̇�z��O�l�|;ųo�Zs�|Ԟ��+fΣ���R�Ap�g=y�S��{�;;'��uv6t=2{�)��~�����zF�<�D�v�=�}�ã�}��\���:�>x�	��qV�8d��ʫ�-^s��;�[�$/�,�:!o(�s�}Q������g��_-]쉽c}�����u�2�g]���0���t�|0�CؖUu����e��0�S���G}ί/��3�2^ܹR�n�CY�nfװK�O�3nn{Ϡ����?B����puq��Wn%��se�d�#ޟv�ubמּ�+��ց���F�k=5]�9߁�Ok�|�}�Q,�VH�4����_q+%�XG�V�t�bo�ѣu������c6A4Vv���m����+Hs�w�v�\j�0��ɝ0qs+�I}���8�3z��̏�����p�V3�+5\��>7w7O������f���;�fp�#�1����V&cV�{{o'�v۵U]u��]p���uz���l��O �J�,��DZ�j�?y��;��3����'<�Dy���RON����.��,���a���[��w�
o�ɏNϽ^��8���s�.3�C�|�H���+O�}pf�K}�q���=�4�m"��
��5��>�X�V�������'�}A���k�nK���o$�����qaw��W��R���]%��/K�<jܮ�L_{\9Z������j�5]���4�LΗ������5,/T��V�ِ{��l�s��������>Y���_p�s�{�1��-:�~�^�N�|)���6��o�Gb�������.��=G��rcS����-��gh��_��Z�����)0jE�R����f����N]��p>�t��ˆ��^��4iݠ_�U��ۼ<8[�dH��)�C�t����k7�y�C��y������c�����չx�ʸ�[h�F�	���*�p͙��Y�]��|R��g�m3�>8�{��Y[\�e���2L�a����T����;{��}�>���rS�wg3�n����c�y"V�dث�k���7��s�v�r�ɞ�7�5�v���%�;v�< VU#Ӹ�&K��^�y�v��'lT�M�ھ�úֽ���{�c�5�MΧP�����&�F�B�O__�ik7S.��#��Z���܋n�NX�\ђ�V�bY�y�h�hjИ��6w�CNs�T4z�M{.��W���i$�Hm����ʂG�]�9�:���%Xo�Y�j)B�_g	T��)���ٻ�#{3�����©j�800�+�R���;Q֨h5/�z�7���,��O���Ȋg2��5�Q\؞�G*d ʛ��z�9��t��)�
HQ�km͹�m�x�3������kg����D�5f��"�Ǣ���Yo�x�2�c�k�fv�p`������׳m��+��D�53�ެה�ޒÙA�;u|��LG1�Q�jV�B��}��a|�n�MM�5���:���=xy�7iӨ��s���:p3p��G�O5%��>��%�Ƕ���ţ� �9ّ�j�s��,�J�^㋫�`\�L���$��i؛����"8.Cؓ�r�ph�dS�ޱ�ܛ���6�|bB�Z�T��N���h+{��oc��*ΩL��7 |�M�]�]�}��ŝ�����u���w.P�ʷ���\�h9/n�U�	]��N�7�nn���oY�@/�;�ev����KF�P�n��*f�2�d33�#A޲�f�F��I.�;h����H�C+��E�۶��i�3����vᷘ�lۖ�X��#�W&}8u��Q��W�%�d�����(t�*��v0*Y��YD��1m�;�� �VIJ�fp�T@2�V�,�j����qc�����v�O�q�уjN�O�%C���GS����'بY��,ǎ��i� sf�&w*2ۑU��[=���nwV�މۦ����̀���|M�b��ǈ��)�p-��]�U����ӍJ�f�!�%ú���+�K�tz+p�p���Jf����{) ʵ	O���7�X���`��4�v�TK�yD�X��u�.&E�'�N]ƵX/�ՀS��#��K9|���>� Q�
�ڷ�R��t�]�[��H=a�Wy�W�D���fs����6��ˆ�]�Oz�!����zl��b|ui4�s7\7s�M��5���6ݚ@�ӱ��bDhw��WtP�K�l��Q
��]t������SP�I��/���:9�,���w?��f@d�0QESQQT��RP�M1Q�IUC51S��KI5)M�KK��USIDT�Lfe4DPQQY�DPUQUCCQ��1Q��%��1�Q�DEL�ELVNQ1UHEE%4�Q	2D�!@LM%��KQEE5TQHU1Y�Q$HQT�MM%E1U���Y9�4��+QUSETUIMRFYUIM�EUMU%SEPEITQMQ��E5cAUBDDEUE	M%SDUID�TQAS&A���TMS�4�a�UT�DdeJECQEfIJQ9��LIu����]_h��������|J����PÔ�2i����*kV+i���p�u�M�^�U���%�j���7����A��tBw:tc��f���q�L헀9�0ll	gi��<X��n�{k�ii�(�/���?���M����9���o{+��u�������.����ޓ�ٯY3hW��/��]gT�<�w��������hMfJ<X��`�I����On�wׂ>!�!o��}&��U�`j^�4F[�e`uXc��S׷b�ޱ<앬�rn^^.�}��7N��1)hC�n��pv�}��`�kE�6�T���g���I�����T)�o�-�/H{>~�hI"����z.3�wN�a�h�I�d:wnfzm��WT�c�o�gy����=�P���g2����s&���K���V��ض���ǭcsy��5�X�T1�7&=8Mߩɕ�Z��/]�{�{ �s�o�{Ӿ�t;6���\6�s��󌿃���	���8�ͼ���em=���*^z��G�V_(/�]x��"��I{�hkx�
_-�~߳���iw��"MF�{�#��J��t��]z x�{��"�����k����`����e��Z��me_R�%F�Vw(�o�<��8��߾�z���{�M�-�'�W�i��D��5����Տ��52��3�Z����=�"��Kktk��:⼔����N�&X�ё7Y7G{X����؜����|�����fWi�az����6��E=V�g�2;��앋�X"o�f��l�1(G:g�G����m�;��F���#]{�w�v�ɜ�=���L��KȌ~����5_M��16ĳ�p^�Cw)��7o�'`6|(��	s�]]c�?a~sӏ
~ެ�e8�-c'��yҽU>�<�ō���:��˦h/ܧ*WX���y��ͨ�Jc3d��S��y�λ��7�'�x �}���~}�#�P�(��y�|zw?V�W��y޹+��d��d�5�4�uX���ίhM���YcE�󲏷F��Ϥ�*�w�HkE�6��%;%k=�+5��#v�"���v�Y=����sz��g� F� �ö{-���X�M؛O�ڗx��5�ók~餗�3g#ڷ�)��y����r�q����ܔ3/m�!�jB^��2l-�c��Z�]� ����Wa7i�D����]��ĭķ�-SE��u%�+��������y��\:�������ζ/d����ݿT�s���Yެ��?wl�z#_=�P�����%�g�7Ry=xgx:>mGY��U�jg�e����/}s\���]������=���ӳ��89�P��_a�}���xe����[�ŢS�>Z�y�v���қ�����׾֗w��_�����Ñ�q�5z3��j���ރ��lA[:��|����[��?P�k��i�i�ڦ=.��G���;�V���Y|/���p
�-9o9G�q��\ٸ���@8�Ws�8�ڨ��������ޥ�\7�-��Zs� Ԟ��3ݟ5��s�����{����S�Y��O.�a-�Pu�ٷ�Od�)���3;
Žgw�v�~S=~���gZ;���@�d��J��l���֠��Y�0zi!w��4����M%��	Got�`��gםqC��I�ƛ:��o��~�+1��$N=M���':�^k��]�Zs�j� �/Ykk�pPLO]���:w��\���v%�="���V���#�G"��wS�h�H�建V�wso�ݦ��0��cm5�ev�<����s7�������gh:!o+�Xwel�ՇU���̉t�no�|�M�_(��ӯ'<�r]�λx]Doqs���O��㓳}�.{�3������:���&w�K��2]�0:�Y�Ι���Tb;�Y��s�]����f��Uǂ*�rV�����P�t%G{��w�.Y�(n�&l�}Owױ����Y�&G
aӯ���>f{����Bv���a�2�v_�]!�?}�|�]?�9.�?y����ܞ}���y/pv}��+��kZߚ�s�}���ߜ�����=���߸~��)szJ��d�sBP�/�}h�+�:>�K�r���-/;�?�7+��t}�Ի������x��I�O�%�����?/ރ���F��w���&A�h����{��~����4ø}����Й����+�|��.]���#�伎��W믾V��ӫ'��[���`Eo�~��Y'�<����ܛ�ν�GR�
���_ ����)`��z9.� z�{��}��|�<��}=�^��e��}��(V	^����`~���͛G�R��k�#s��P�����R�hy����V�{�{��t}�<��|������2��k����ᒾO�q��1�}߿>V�x�C�h$J�y[�� &��ǩ.�m/k҅Z3N9�k�`�gm�	G�-A�a���9[kr�N\��˖R��cw�5�'�u�M���d�+$Vɨ�U�5kl�6@�R��t&n�Wk;��}�Hp
����qR�(Ȼt���_2�U���mЏ�������#����=�K�u�y+�d������z�?K�)z~�K������t���y�z�w����G�����#ٳM^w�W�~����������J��~���ع/��p~���r�Լ����&G�`n
W^�h9/ ���49���to��y&�?e{�������۾~9�}��<��{�+�}֍���a��}#�콟�����u��=���NK�7Jy�q�ԯ�r:?`n
G��}ރr�2C�>����������s냐�ӑ�x�K��z9}�;7�<��r�_xi_/e��Z]���K��	��'%���3�K��XjW�7{׏=�{��_zy��޼��g���&��^�5��~���=�y�y���Jd������<��~�4����^��w>��δ�+�~��.C�%?A��
M}�f���<�<ּ���?~�^g�C�;��a+�;�=b}�yu��%��foA仗�`x�H{����z����o@r�=���0XE��c��������t;ϓ�����ʯ��ڸ9ϱ���)?f�y'�F�<��X�f+�����䧻փ��`ϱ�H���rܽ�쇇;��z��:����:��s�k�{��u�}�z��}���w�}�]�^���;�AJ���C�P>܇%�d�� ����#�}�z�吻���I�2�^I�0�
�����A�}����}4Wo���9m�ľ����}/�����~���i��Z�{/\�AJ�����d���rd�FK�X;��~ï؎��?�i=�K�;ߺR���3{��g{��>���:����]��l뇒:�d���w'��w���]��|� �/�SѾiNA�s��y����^�srd�]�tkr�/?a�M������Y�#]zy��߽���p�s�&�TܥV�75?�;"D�GHZ�
	�4ɸgouZ��\�YTw.�����K}t�[edngE���{����]��ue����U}�V��[K���ψG���i���uL����v^'ޮ�O<���lO>���]oz���r�_��s�R�Ry�rWQ�{��䜑�ts�z�pP�o�J���x&C�>o�?�wO��s�WwG�4����.����s?o��yֻ�\��{�þ��ݜ^�~�G�9/ҟ�������>}�=������+��7���������Bts�|�r�'o7�2!�y֟�<������?k�����~�u�=�����~��-'w��:u��^�#��:������y��w'�{�<����~�B�$��r
WQ�{��~����w&��2Os��U��ܷ���3Js�?R�UJ�o��;���ir�e�w�G��z���>�#��:�r?w���^C�~:�K�K�.�����:�z9J�5s����y����w�^}�����{����w'��{�sH{/���~�G�!��u.��X��!�rw+�d~��nG���'�w {_}��������P�����5���m��h�z���ލ˿q�9���_�a�:��Gˮw��{��������ptk�K��X�~�HDX���G�g��v��_��u�;�����s ��@s�����2z9��<��oG'�I����wy#پkp���|��.�|��Z\����=���;���y?��k7�~ֹ�\��y�W��wz����~����� �t������2C��49&��d�w�	@r�7��b��y�%��>���+��=>��>��>�(����G�W<��I'�w�޹����wl5/�z�k���kB�'������_~�n]�Ht�C�r^^A��t�K�?o�<��/G���Kܽ��J��~���ty�}^g�w���=����prW��X�'r�sI��
O�`���ykH�����믿i9.��;7���^^A�>ҙ�y�컗�;����>﫿n����!	�ߓ�M��!��E������rU<-�s ���w`�'���N�LQB�C������ݛ�:�v{ԙs<3�fS��'�&�;����N�}ON��m���J�k\�w�W�Wl�7��̙�ir���EYm�4���]Io�}��������!=��U+W������{����/[�I������������_�ܼ�%~�q�XO��OߴK��N�z 7'���P���S�g��5���g�}�v��/r��}b�9/P�s�G��.���������(��/#%�k �M��u��#���>�Ws�Ͽc�E�A������[�������>����+�;y�GR�#�oK�O =7�/#�}���w�yR�s��?o�.FB�n���{������7�L�z������ݝ|��a���|>I�x%y/�9��~���;9�GP�W}�4~��=���d���
w��y/�;�R<������a�x}�_�߯�ٛ��b�=.����#�~��|#�?}�ߣR;��{ރ��w/ ����/Rty�?+��?}�<�������
|Ġ�ড়�2�����8&{n��V��^���,��̏�}=C�~R;��wP����wy=��K�O�����^��}�=�Kܞ������O&��~�z9.�<������{(Uj�3��׷��H~��D���JO%��Z?H���z\�߸��]C�ԛ���:�����}��y/rn��GR�N�w�H�A�}���Y���u�ߘ�ܧ�}�G�Q��2�F@���=ù}���`����yּ��}ޗ;�w=}��y/QѬM��r:��w#��GR�Mü|�>���������<�g�|���	����I����)g���w9)��4����/���_�����%�,��yk��^��X�W���>����ח?s�k��p���|q5&�x{��R�
^�y�=�p�
�?{�~��oXr?J�>oO!��O|��y/���u���{w�4�/�����K��>���U��9��ʲ���C�����#X��͜�E�[�q˺X֪�:���4��n���Ҹ%X�Ö6]�#��w.*�[w������wt:+�\M6��j�����W�w����huY�6�.U���GuA���,C]�Hnw���~��������W]����5��_g#��'&��{ՠ伂���4�n^FF��w'$���r:�ܝ�kO%ߘ������C��{�����~}b�W�jQO�t�~���~�|e�C�79.��u�y����H�GRn
�ޭ��d'O�i2˸��ߚGrrN�����̯��ߐ�����"�G�:��y�?��|��K�s�/%~��C�'fby.�����!�����k5+��u��R?_��I�w9!ѿt�%���O���~��S
{?cݓ��������J�'=ր���C�s!yy/��I������{	٘�FK�)(O`�;��G�w?�9�~��&�����q׎x{?Uw�O��c�މ<����_���>ҙ�?�^�K�z��`�K�?�Gq��s�B�;�.M#׸}K�)?�{��t�|����oߗϿUяX�"u#�x{�I�w�)ۜ�y.�������#�0��=K�_�w���^��;�zG��^���������pd~�������s��aÝ����\���y��<��G4b�����,��>��w�)���^����K܏^���!��<9ޗ�Ծ��v�JrN���EU��}몊��-���5��%_v�\����{C��9�y/?a�K���惖J�>��e�{�;��;��I�]�s4���=��|��#�2?R��~�ߐC��o�����3������#�?����9Ӓ�u��}����#�c��i��^K�<��+r�G��܎G$`�P�~#�N��T?/ѭM��]y�ߛ���|����P{/�S��A���y'[�K��<�}�K�x��X;��|�]�9.�?}惻�{�r}���^��>�˯}�g�y�z�߮�l��;5����c�<�<%(���G�y�:�^�woKn*ՐO�֧�tq�ǂ��z��8�`W%Nv.�(x��Vq��y�Ѕ?�ٮ�Xs�R��Et�.�)�7Ҳ�f�X��I*Vn�X�iV��W�&\��"�g3B�v>�ʯ����n�z5������2O�����GG��Ի����4����>�	Cܾ�G�]����r�W}{���x�A�_�q��'R�~��`��EE~���,�+P�޽^C�U�p�ic�yg�k�>ɐu��r
WQ����AHt惸w��vsz!�_?y�y/��z\������?}��{��ߗ��,�]�z�X�B�y<~��M���OR�&����!�u/ ��w�|��o�9#��oG%�d\�Op���vo�C�}��K���uUڧH�C{��~G�f�>���ԾK������'�>G'�������{=K��5�/�r^A[?{�{��u���:��{<ގK��>�~������>b������O7Wp���ݞ���/;װ�_$:<���K��X���z����?��<�����~�pR����7/#'���p� `�_~#�}�������ױ��aU��g�����ٹ|���ѹw/�����/%|�u֗%�C���C��F�#������&G�`n
W^�h9/ ��>�C���G�k�>�}���g�{��o����rg�}�Wr}�n]����h�G��{�i~��ֺ���Py9/$�k�?K�����G_�! ��̋�`8��7�U���߳v�S9��K�d�;�C���#�y�2^I�{���^I����}n]��W��~9֗r?F~��}��0<��sC�1+EW���5���~ˮx�_�2�?u~=�����9�~�=��伌��~�<���ßiL��s�>��������=���#��^�֓%}�ĺ��G�G�.^��4+g��[�����!��������y/�֌Wp�?u��~�����K��N�ރ�w/<����C�_��������^�ހ�{��~U���~�`a����^51��R��<a���h�L�fnȑ�w>��.��3s�Xc��K����	ȭ���X:-@��;�K�=����_\W�,-��o�W.d=�nQ읔.)ǎR�S\�U���We���u�30��1<�P�o�6��L���꯾���;����~��;��L��O�=���({� �y'��>���8B�#ìO�������Sy�܏W�|��<����?w�����_�/꣹��x`��������w������^����]�R�
W�x����sp伌���w�ѣܾ��{�r�]�[�I�2�^I��4rW�pu����ֲ͖�����^g�>�\|��<��_���{��z�駾u�y�������o�.FH��%�2\�p���|~�w/�_m|8�>�~�7��,ܺ�������sjV��Nw��du?IӾh�NJﳙ�������&A�_`���4� �^�w���!�X���nL��)}�?}��Z=]6��ݖ��-�'� y�z�/r�7�V��&��\��d����:�y�=C�(N��IA�}���oBd>C�}i��z�қ?}����Z7kX�O����?W�}� �|���{&��S����^��??}�=������+��?�G �u~~ޞC�(Ns�ܾFI���L�����x3m����?�e�0g�~i����z\���׸���K��X����:{��]�w�G%���׺C��]�v{�������R����%�2ZS�x���oj��ܲtG��ퟪ��Jר�8}����}��+���ޗ.��]�H�y��X��y��M���G�y!�׺_��^Av{��{���G߿��m���bDrH�0����+�8}��q����7/�����e�_��H�!�>Y/�w#��O��r�FG�NI���5���7�Q���2��ou�3���.�i��o��OP�A���r]���y����{�b��z�.K���~�_�n��u/#�c�_##�Uk��A��e��
H?��>�wle�R�n`�X{�S �hW=u�:̵W2���&R�oIΈ9yD qJ:cԪ�4h
�SiX�
7�k���*ws��@��ݝgZ��p#r�{�BR�̛���R"Tt��;e�:��t��oi�Z��-N�T{i8��0��t�xv8i��\+���{��b*��o�KRԧ���h�v��  ���Z�d��q����u�O�N���CL�����4���Vt�Aիf�Ŕ�,J���˻,+�C'Wujڵ���AYRR�̾zq���Y����{�E���b�	��tz��à`�n�o��-J�R��Ο<U�b�k�U�K����J��G��]�ɓO;3�q��"��_4����p$rF�um���m7�c���I�%�\W�iC&C�p�$��_�U�1R�a��f$&*�Z��k�%�<ҩV+�1�,RvM)͉}}L�f���9�L}�p��[}\��SC���G�&��q��ՃN^7Wim�!v&[!os�lܵT�C�ۃ�ՠp#/�� r���խ��==ȹ�y�	"��ǔ���6�6v��#���:�K�W[l�����mһ���cq�l�VƵf6��Θ�� �i��9P��c�/�5�|�ݐ�.�5E
������MN�!���m:c��F�{�pusPJJ���mve忨t�Hc�L�q-��5�3�a����Ι��]���-��YI��*M̷H�����s�x���]r.�,hX�mK����Ƹ&2��s6�u���`uwZT�q�w��Γ(۔rŘ�@�:,�����:��)P`��g�rmVg<ں|�g�Ё����ʸ�5��w(#yVn�]Hvjq���������m��5���3Ƚ�ac�s����e�9�',��O&�2U�g�KC��Z�̡q���j2X9F�	9s%���`�h�b>�WՃ4o���=��h�@�~�A�T�����"���H�k]������^�8M�p�YU2���E��P	�G�^K���PE��:��̓9W8q�ݝZ��ʐ��ݦʁ����v�ŏw�ȷ{O�8�zqI'j�ۥ�2R�"���p����>g�R�R����,v-yX���'-|���"�'��b�&Y�"���=k9YN6띩b�[[u0g&�Ŏ[Ě�����}�(��%pp���,K��Mp�skt,��,V��4�k;�6*����F��Z�;\��(/��9ܹ�s(�/n�Z�4V�ӻ���ҹ"�N���#�2��0�������*�xGn]l�Q�Ǜ���W���8�(A3>=��^4�4�.N#�v��Gg�Hes2�
q�j]w��.YKyD�g��F�Rw�Y�􂙶�*��;�Ѭ3if�{�V�u�,�J���k�kqڱ�=�T��'�}2�!�J���1��$��g�]!G�͇�m�(t]rm��}����o3K�%m��*�0  P����J
̈�(�����"&�i���0�Jb������0��!+"*
&��d�hb�������"f �b�����"Y����Z`���"�j �I"�$�*"���b���)�()���j�b�����&%��� �*����*"�"����b��*�f�&�
����&*�j"����&�$��"h���`��j�(��"���b(�(���*JBh&��f"��j*������h���J�� ���(�"��f"f"������!���"��������*"����i
�*����R&<������#c^.P�y���/5�L��g�����ws�GFs�쪽�T�ˉ־k���Ϻ�߿���~���ߖ��͟��(_�k �;����L�r�2zߺp��oG'�I����wy#پkp���|��.�|�5֗%��{.��_ֿw�[��*z�I dħW����Կ�,����AB�޵�r]�Ht}�$ܻ�����(A��ϱ^I�Ò�w���W��z�Z]��jz=�y�9�[�޺��î������p�FK�<��`�A�^GF��/�rz`r?J�}�M˸�M���9// ��L��o�y�#�_~���_��s�pX�Ư=�y~~��c��}���3C���k$�S��7&C�)?9�{%�u�5#�;�A���Ͽi9.��;w���^^AϱL��ǝ{���"�ij~�ܷ���z�z?߼���gN�GR�oyѭ�OWi�H��m�H��Յ�K&ͩ�n�)�9�d�2�g[���7�4����7xGV�+�oq�G&�(����ҧ�U���z䭾%ؘd����v=7�"�s���=���>���V9�^�����̕q���pHkE�6��sMٵ��!�;ff������zM��w~؍}�G�S�{���]2�zX�s�m�h��]v��P�es�J<����=w��uw��*���u~u��w�ᜰA0�X�B�;�tI��@r��E�m5vmx�s���Vv�_a7�/��|��p�Ȕz����7�eb>�	d^>�ڵA��ط�ל���R��x�0�ޭ�V��W��@,�ٮstv��&6��W�}���0�Jw�8y���u�V���`��o���n>R_�_��ܸv��^Uv3�7�)y���>aP����Lzs��_��;;���O%��!�ᾛ{�JMtyt������3��O�z�]��>�P�%o����P.[��o3��e��^cL~����ϸ��qk�oF�_��rI�w������:1���tgݥ�q�/K3����1�����w��y�?`q��jޯs��{nۛ,�r�����o���KS�[�Ώųo�X	Ζ["����r��״foD��1����4w��S��b���l�2g��>��ї�Ai�=ͬ�Q�q�[݁�r��tv��b����ة]k{
띘�y�s���3��a�fw����7����σ���gi�o(�����UL���~��}gvO���MNf����}:�NyR��3��xZ�+���:��0�=ٱ�Y�qu��&mٮ��˯��^1r/r��×�!�_��r��X��\ʭG���z���wm5�j��u+��z���R�_LR�Nr���$g'V���drʂq�w���7���OQ��˲�$���`���\0ѝ��k�s&�W^��}߾��|�o}�.>�Ϗ�:�BJ�/��������I�.W���.hR��}���ImƷ�r�S�n�7}yBt��xׯ�*r�nu�V�>j�g�mt��(e֟'�]K2��g�jd۱T��ʡf�<������K�ڞ;Ƭ�$a�F{ڽ���m�櫅��z,	&�S�	�8vPO}V*:�Y���ş8=���g��ӓ�3�G-�p?��t�Ϳh�I�p�,����fک�7��\�V���G�i�;�n9�Ę��s}~��q�eJTt�F��6˓:�Uc�����s���Ƽ�`�q���\��U��p�_�މ��& �|���v����[���r՝@�uA[���/���e��1y�W���;$�w��߶�y��=�R�˴�nN���;����kT>�'~�s�]��}�t^Q��\�4j��;^�i�l!�d^`0�Y���d��G\�5�*���:�v�Er�xwU�S��� ��eI���,�r�ӷ3q�f|�M9�[(�kq�W�W�L�p������u�y�I�nܧ���S�jh+��u;9�w�m���.��1V��߬��ǋ5�ݏw��� U�<��FK���:pjOg�{r�����3�����g!��`�O�~���K�}��s�59���K|h���z�U*i뤽�3�}�8���tu>K%��Tf��I��q����ns���坻!x�l���m]�DNύ�
>l�~��_ڽ�_z����}����q������5S9ת����Cx�@|GE���g���By���4�Uϓ���yr��ͮ��A�׶�C��k0�\��{[��~g���y�M{��l�ï�z��_�N���%͖��u�%ή�S�z�[��2�v�M�����/daݍ�K�̏"��֋M�2����v��z�+u[f��{kzu%��C�:�UO����i��$�-��_џS�b�e���q/[�۽`��W�q�]�US3��ݷ3���*��q�1���c|�L���d����n�]�.����f<���r����[t��T��\L��az7xn���z�W�y�S�j᱆����GjV/>����ޔ���{$ժlTe�)%ê��3F��ۊ+��ݻAr7E��%�4��\�Ĵw�ﾪ����ݗz�y�6���	�*_���w��}{�c5�X�[���n�4�KjF��'f���v����׋=vٔ�;6���\	P�`챘o�wA�='k?R�״|y�^�6�kj���ۿ'�q�>�e������a���m��l�0V�aԼ��=��'o�{����/T���G��ӑt��}����[��p�SG(��9�X�U��3�1������'#�qz%�1�e�}�ٿ����ޞ?p�(�~��b}^��)i�����ׯ�U������S'_��]ɳ���4�����q$��}uY9�~��p��e���MlJ����w{o�^��	^2�)�;o<�\�{��R%�?C���v�;�腼_������Z�[����ܺ����ٹ��Sm�yX&I��L뷁�mЧ/�s�X��>;F�y���4�-$R�����d��+.ɨ���&Y���N>������S�P���gV�lTJA\��U,�0M�PD�>-���/�oT��!�;v+�\M�;G�>8WB�e��o�����������{��������O៽�����_�k2�����	W�ƥ�9/�>�.Xn�>�.������}�w��ύ��:����;�k}��	W}v���aɵ�_y�k��^u��Fz���{,)��۬����؍r<�*cѕ��r�4���0���ז��5g�s�ܭ)=�(��-�ûfg�П���.��S'�v=��-׫�\�g�vl��GۜV��%{{��ԣ;I�k;���y���l>�c�tI�N}�{����q؅m����:�MW��Ax�}�'��"3;��[��Np{G�f�gn�7�vl�.�{��Fߔ=���ŭwpm{��n�f��{d[ѩW��3y$���n����Y�o�ׄ�8�5�W�^wi�жٌw�½����쥇7��'�Ϳ��N�˷j�t6�k��㚭��l�o�[6����Cѭ�]�a��k��i��Y&�ǧ7��f���e�17�"��К�p��L�Az�s�$��|#��ȷ�J�+}�t�'wz�T���Q(�Z{���9�U��A5�(RT썩�m>.��.:��uǱ��//5��L���*v��,�u^�͆WL�}�}������x��3W�c�5I����gh��.�N�|*��cg�:��>t��`{�q�����M��o�m�,�|��||X���\Û��xV{��Y�Ōg�
�6�>�'���T��r������;N�Cx��6���r��WoD�s��S9t{�2l��o�D������Bdyy3��x_���W�E���;��
��9D��Y�@'%��J�/������_����%�?H ��	ift�οk潕 ������>����]��-�kپ����@^.j���zNy��� �m��65�4�ʿ��o�c���!��y�lX�C�F���iOv�и~j���$��.����;�W�����f�}22�N^�c���3;�>r-[��PwO���-�=���I��<	;OWL�jω<d�=�y���X����W��ЬU��ҽ��N�L��#��:���*A�Z�t{Evkg )������+U޼���;����-�!=�����ս����Û��)�b�7��P�K	p�ID�FI�p��	�Si�}W�;yeͭ�}��
Y.�mH��L�,^T\ƽWc����}�� >�:���6+ϧ�]�vl��z��g�>���Ƽ�`���_x���nIp���X}������1�(?^�����@vm��W�A�V�r��&C���{On�^ti�ϻ�����^�xӵ��'�@\��i��k�o�����_Dc��^J]�U�o^f������<h��v�R�O�aw���)n^��2��t�|�����/��LI�����+;@��az�nY��IS\�^�X������:����!�<e|�適����b[�Vt��y����0y�R��фhC�u����rl���M�eL헁�y�?n�	�)al��[�Ls��xo��r�������x�t�o{+É]��<��2CٗP�n̈�q��}!҅�u��p5���*������la���{��佼�g[���5�k�ψ{����S�¶"�r�|��w �6��ƒ.�ֽ,n긭�1kX,� �vWn����f�Eڥ!��^��F3&�;n}{�_>Oy���-�p]�Q�� �+�*��Sd��Юf�@���}S�vs��q�Vv�4YǙ[���$�D��nլ���=���U_U}_S��/j��q~�wk����Isn`t�g��VR������(k�1���p{8�ɣ���-̎�@�֋rm̩�מ�{j�{��e�v�O>�Ǟ����ͪ�)�G�k���܊�,8��}����B�V�ܽ!5���zR���Vf{��ۛ�`\�f{���m����[6�1����`��ʗ�G���}%�u�˶0k����Sm�e�&�u<��P{z^�vj��z��F��Պ�s���ϡ{�fU՜�r�ܦ��&Ó�o��:�M3g{Y�����ͯ��l-mRW�o؇+bm�_TkVM�����Z����^���+\�R�9ǹ�'o��z�Õ�i���g�S���w��:��榺��,�p��/���r���ՏX>��8U�`߭�$��jZ�;�%��0��p��g�~2���6���c���j�m�QW�.��Τ)��S}�[�Rk��]HՖj��k������h����� 9�g�Y��u�u�i�K�N'52�LZQ,�mG}\6�V�aP�<w�C��R���Tw8�[�խu��T�S,r���gnE�8����e�����͗�g��{�_��j��>1�L�|*WXM��L�4��x�OW'�x�O���]O�ӳ �nY������d�\�yڃ��p'�j
�w�I�ϳ�N*���<���8���v���b��,!�Ár������k�����Q����������s�ɒe�λ��t셼aG��PI6��}�]/r���TC%<��>��IW�fW��}r�KU�D��s�(�t�O�l�䫩��^����N�f���Fk޼uG�}��^q�/�˩�:��%k=��ʱMn_�����������+��Y�N�e���x'���oӭev�M����2�g��[�G�ӳ�M�0Ww4�׾���
��ؿ�����=_;�c�㱣�.�{)��+ق���r��o��Y�}^�sd�a�
��6$ǧ>�=C��vv;=s���E������ ��r���h�T@�6.�nQ:���R��y(t��m,��o1�)����h&�E^XY�7�4;m>p���rn΃K2�+��)(L�p����Ӷ�Ok����N�:J.G�wS� ���K��$��g�fͣ.﷡�S� l�f�C�PV�/����'fu\ͩYPh��]�q=��3W�杆X�x�s8�T[":�g̕هg>t��[ʚ�;�*u3^m>�d�]j�7xv@���ٍ֚r�5�Y
���q:���}΋?kw&�e����Z��t���,��py�^��:�K�#�j�Ż�c6ὼ+d�f�P⛙�1�����.h�t�Ĥ �c�W����'��.�HGg_ķX�NenV��u�v��t�%� �9�!`��Y��ϴq�9�ǰ.�B��Woh�M�F�|�_!6Q\bmꇐ��k4Ӝ�d����v�.�+��B�:�*Z���-b)ls�,����*�%�]ӅJ�w	��4nj��ggu�����+���׵+(�4�s��N�ؔ���c���r=ǎ݃����v��;]���a���DL�ot�3�F���'�gLq�H3x|gXw�K�8B��뮨
����/_�DP�t�gt/0�J��B�r�o	ʋ���y� �72��k:7DS���t���&\-�h�X�E�Ūۺ3����Z�y�֤4���m"�&��9���1�nb��P�в��3���d��#��`��7
�t�F��k$��&^vQJ;��pzgjN��"�۶�U��_x(���n;�_v������YC���;�rM��7fa��g=���(���ns��,�Q��Ԗ��<}��*:G�ެJ݅څ�W9u�dّ�T��Vp=,�X������Ӗrer�h]Ym��lx2
&���h�iuW%]�������P��p5Ƭ�WQ�B��Q��Yڒ�3x!�]ySHpK�y���Z����\yv��LD��;��e�fQ#��g��ͤ��"�x�z���V6�������aw���V�VW�uLC�I�#�L���ms������i;�kQb���B���iU��άk4�#h�"'l:b��p<���B�u��]���,��c����..+�V\Nnj�vg��S����׮P��,�"&�1]w0��چ�hR}��]�w��r�T j��6�nb��5�(��$��ל������o�̱�dw%������hnml�K�^�cѽH����A!��η3��đN�;�|6�f�� ����2���wyХ�� ZOof�&�t�v�*ڻBJ�ªs�u$KC�IPP�g��O4�I]ghU��'<F�%�qU���ƹ�9p��[IV찜�}f=�Uv2�Z�VZ*�iV�|�q�"�5*���Y7M���Z�(\B� �l�z�聃�'5y���Eb���u���E���c�p͆�]�Y���m�G�ۼ�u1�o�z��d ����j���(�)���Zh����i��"�"�JX�Z"��("��bH���j�����*(���
"*B�������&�*�)j�B�Jf)���h
�%"�������
���
������b������bJJb��")Jj� ���
��
���
����j��"j�	���Rf���*
a*��Ja��(��&���
��((��(()�b(�")

j�h(�&!��`��h*���*!��� (�����I�H���B��h���h(������	j��J����)���*J��>�+� RfL�A¦g4�<ە�)w�]"\F�˗�r��L�L�����%��ұ�յ�ql�Q�\tq��t�t�{�^>z�������ˁ��俪���+\_V�����jw���\>1��s~���n�&SXg��{=���s��d��Osóm��:ޖK��62I�1c#3�n�y�����޷�9��k��'�B�[f1}�p�ծXN[�c�9��V�9�q�;�~���M�����{�6�XS�[l�o�[9��nq���2{�Q�S�\�ɝ�3�:��;���au;Ke�����pd���r�y�N��_�i��l���`zf��Y֎��ln�|�)Lz�X{wU��z�}R���l����8ʙ��.oc��������`Fa��P���ǱIշ�ﭙu�z����������vNw]����g^2*W�R�	{K��7�$�Fߩ�����zJ�S�/�C<�_x���x˳y$��&�jm����ۻ�nm�����x���b���`w����V�����W�c���Ө4Q�)S�+Ę<�;&;Ua.��۩��=O�<4�4�z����Hx�����,�xWZ�Հ:'%"�=t4��e.�B�n\���6��o��AgEp������%���؁E\sٍ�?}��}��|j��<�p7^��V��r�J��'Q,k<i=���_��y�(�׫=�p�����&G
a��	&ؗR�xL�ׁ6���U�߫|�t)m��Ԏ��Uz>2B{�En[��A���a��<6G���g�d��n{�u��o,h���G�/���-����W.w�K5,�����Ϳ^t�<����3��}lk��>�|�>�~q�^�
�[S侙�;~���.j(> ����w��^��?xenL��hڝY}�O�Վ��Ϲ�rI��~�y��=�N�˴�j��)�C�Me���Η�7�c<����	�����v��rz�Vn��;^�a>>�5�k�r���ŵ۰>����{�XNt�Ԟ����������c*�/��L��:�w��e�	d�+�쐿�2��3�7�m�o�:�e�(�������w@x��2��	�'���9�ʘ�9*�m;�`X�W���H#kb~
�ڬ{G5^�Fߖ�w�4��oLԝy�C�%J���U99H��u��^n�Ԡ�a���^��;���˾P��-umAk�X�]{�U!{��}_UW��^�3�[q��0��!;:�u���{�{�W;eg�s�:`�j�zC�!��s�޷�Q3r���5�+7���N]|����%��R^�^�*ڞpn=��>�V	�3�J!o�>��t��볦�W��9D�j�@߅I�[����(��n<�r�r����z�4���������d7��QF���N�\U}�K�r_�6�N��x�y���w�^��˝��}Y�=������-̏�S�	h���*K����J�[�O����>�>�[)�n_��b]�lF�nEIlXp=
+�g2�{�U��Of��h�ɿCg���9C��O{(��*��9�Lnt=U�:�pw�ϸ�1��T���l�On�����}���Оz��t3=1��1rw�G��R��<��{z>aP�|lI�Ntݽ͗�9��Y{4G��MT�nͧ�8O�� ���_���GZO���O��[nL͛�U�R���&sku��	j�δ���Y˪倆���u+�T��ݯ%yk�"��<�B�9��(T��3���S�+��*;K�l2_1�e�A7��(bG;,k�]�V�1�s��?}�W�W�w�F���X��wm��^�f�Lm��9�[�W���W��w-��%
������V�ԫ�8�=$���K7p+����\����j}�����R��am�Ŏ�p��-9s>��8��|z>v)�=�]�|X�Ux3t�%�<9����x����V��~�fw��u�f9z���O��aY��K]L�j.�Sf�a0��yL���Q���7�ל���f16Q�:8�h�C=�N�Z�z����w؂Y��Wd;�r��{��
~�X�v^8���E�(�%0��U=�^�wc��zT��=��?w�M���.K�:�<s`�[�)��G��g� Ǩ����:������=*y��K�cR�䭾�({z��,S��Vgu��t��T�]X��7л��6�{�̕q»�S�f�[��J�u���t9�m���Ay���4��y-��d��|sL��Mg����z ����9���(8��X׎ك�IO�C�^v߻���Q�oJz�s��ү�_i��]IN��Ч���U��K0L̗�@�g
.�����Ƞ�Y�ԓ���_}��F����ϥx��ݻ���u���Ror�'��I�_5��f�;}�������~c%wV�e{��5�`�+��g�ۏ�<����=�˦�_f�o�^�}�&�{�q��t�u:ͽs��ڙ�oם���-[�P^��U�o�y��OP�=�~��=K�M��d�¼u¨�1oPog���V��k��^�mN��q�3�|��!�TN�����ז���%�ӽz�)�_\}�L,�ލJ�s�]H��Sֶ�zu��y}]��~>���R���	���c��
�2=^M���ff�NS�#��sf�P�4�ꖧ��eã�d�**��?K�ϴ�k�����v�Fd��=c���6�}j��/�~k�r:w԰�n3��.����zd�	�Sɳ>k{�=>{^�|-��}@�]J�=j�F6Rx�ma�-/[��q䫱'vw�r3ʔ�e���{�	յ/�4*�JLU�ľo��+PͭWr�Q�\����bv�NsԄ��&@���u�e�l�cfǳ��v�5�{�X׺(ڻeΠ�T.���u���UUUR�~���n�������_Tfǟ��	�W�7���7�>�,뺳w�S�?�Us����D��� |����;��~|��M>�p���ք�}�+2���E�aH�����i6;��+4p�w�ѭ�z9C<�_x���Wn��'�9v���9���oK����Ƃ��b���B�}?e�z�[W��G׳��ߕ�~���O�J���0J�!}��Rz���ݩ��{/��B��|��[��b��wLȮ ��_�
��J캣�mH����\>�Ja�����K}��i�f��Z�?��W��
�s1��QkV9�鹗p�^������=��w�G}�
�G]�����|sz_%�7��K�%cZ�g��!�j&�^)�c�>�^	�������>TP��D�>lǧ����������~׸��gk�Ռc3�\�S$�&����$̯Jk^	�&	�m;�7���u	N��z���B���;�F�+֔fGS��}s0�^F�4gF��S^Tp�6�[�%�HXw�����XL�&�t<�KI[X!K�{&���Ь`Ր�kӍ��o�Ηj�
���+�}���ۛ\.�Aͦ�6�vᵐ�N$�M������<�/[ޯO;�q�yf�)�E��mF�+|f�t�Ֆ�E{Rƫb��c�aɞ������o�<��^�3>�s��B�`�wڕeY��V^U������}���3��~���P8(L(0}ޤ�X��Nu��Թ���=������zr�{���W'��<ى?x^�w�̆`�d��?\$��i
ɴ�fr�[ˠ�,o ��>�T��y��l����@⠖����Ţ���v^;�8'm���N�e�����g,y]����Iث�f�Y�,�<4:�
��O$�ĵ��P�.��v��˚�ۄ{�&/t����fsxwrV�#�������ے����-#=.�"�����:^_$���AVK͋*��ӷأ���्"���i�=/9g���re�4OD��WR�i+Z�� E4�������.Q��?	W�A�EB�`r�.��h��^�#�&����;V(8ѡ����l�JUx���;��|c�����eE�z`~��xȕ/X���Y����}~X:�-A���9z�[�j�`2���{�)���z��p<��}�PS *��w`�"����5m���T���vycنu�rUՌ�T2F:��e�=J��V
I�3�m�4:��;jA	wۯ�k{]�w"�,��V��\Ew諭���Y�M�? v��I�Y���)yh���Z�����Ň7��A�Iw��x'v�)a�_N;?]�(�u/+�c��6|&���KʥϹׂ��\3N�+T��}��aE9|�7�u�IOd�bT#��N���ýk�<+ڦT���sƝ�:�}�7���h4�j�y����ǭ��hߜx���K>�zE�m׬�k]��L�g\�U;o��/�s��=KxW��k�}�!I���]��^ޖ}uɼ�Չ�f+Uw%]�Y�Ցq긝K��y���P�W����n�9��� ��,����q=^���W=C�bf��ҵ��zϤ��Fr�x*�o�}N��tOYR"��Fm�32���K��&9���΃����*�ٷ2Z���������Q�#l���Қ`�a�8��,�h��*�9*���g��~�cg*�i�o)j²�B�G+P���Uu{�:hw��3�q��Drc���w���s�4Ѹ}��jy�@�uP���T�*��.��*�=>;k��0�}����cpR���˚x��a����nj�C�3�����/�]�2��y�2�E�Y��D R�nF�YeE���1�D��$m�.�l�6Ө3��}ۗ;pp��n�Y���;�([�ag��O3]7A�U�o���}�}�Ӎ���S��||«z���Y�ᬳ��XU-��=h�,�49҈�1��^x�GΝ��8g�!�,.�:�}�W�u�kAOP�瞵�=P�����g���+�2�[��\������B̥�X�fD��{s����}�%T>iK��(����YENW\Ǫ�ӔQ{v�2^�}�>��	<��t�ZI�[ϛ���@v���t���8�; (	Cw��.�Gسg>��9KA��zR�>��K8-�)r���U�ژk���!�h�[[�~�6�P}��K��l������>G�O����A��*yX��{|.�_�gA,V+�S�M=����I+����� 4l5Â����N�Vh�r8����T��Ӹś�u1��=��|��g�A2������[�un!�P�\�c�cK�ή��}��&�*��M�W��);*>��B.ua�+�E��L���2���@}�^"�8,o���Ҽ�r�/o�FV�����Ń�p��?m��r�_�υL+��v�{�[���ͱR�qu��xSJfLHeꔓ�N��0.��U]��m�r�K��3��Ŝ��=���*��|}. &C8�F�����\7�]�|3�ʥ�R�ǖ�0m��w=�w������4�%��>�W�>���Šfs`i��Xz���W� \�=4���+������8'�0�����v�T.�;�B���]�Yk���=���^�)�Wg�of�?!��s���p��G�f�$v���P�t#bb���|�j^nw-�ΚO��<�q�+řS�� �X��
�oe�x+-6��eS�b�g-�~S����ܱWk�h2'���bV��S|�F&�--�8=4&��GK���L��?{yԚo4��@T]Ոh��i����m���榩�E3z�+#ڮ�F8���yf��+iߪӞ�;���.}��H�eqq Y��a݇��}����c'<����XS6i+v�ܳ���W�b��v�4H��@֮J%u���̼����di�R�� ��{F��Uup����na�|}��;�똅�@�7�f�+��Eחl�mD��	꣪ p�>�;�n���'{l7�+2�\\a��u����H���b��/E/��6��W_�ڌl�c�b�f�r�:1gt��+"�]�\	�(C��>��3�*���U�{ȓ�����G��p����-0��ʼ�eS�M���EӶ�S�Ih�e��,3|����D�����c��簶�^o�Q���b�7�5�E�]�����"��~l�GL.�L���@z���T܂uq�RM�YP���xcQH�u�P� ��y��zZ����,0Uz�x���ݳor�"m�h��M;=�qW�dɵ��ٵ˃ʛ%F��p;5!�3Tw&+�B�K�u}�ȇ��j˭�wi��c������V��]��'̮�"��u}�K�yCy	YZ͓�fu�&�����ޛ��
��pee����f�5�=m��Zz*7Θ��e�U܀�{�Ić��c�p]�旂�;�46�F�Z+��쒮�y�޺��@�Y9��t��-9��=}�i��;i]�a�qdn �������}]��ӫV='�V��
���8�����dIX��8�)<Yt�J�$mF�vc��Mnj�iJ�k���#\1Ů������޲�[��,1\/����W��`����CT��f������:M/t����}�\�TZ��eqO
]J�	b	��Jٚ�Y ��O�K�<5��{�t(��,��פ̺Jj ]���M�<Ku5+�r�DF^��]�sV;���=�[�jU�\�Z,�j ����t�u]�)Q��`��,��a6���q�*=ݳAʍ`p���Lk.V�݉8] ���î=�����Z�N��aI�bP��%�rC��ꇁ��c�Wf���Q͙�$jK{�+3LJ���q� 1j;��S�Yu���BdGd(|{�D
���������̂�����']��ý�|��-��X�Q����̙Kx�U�m5��R�^�Y]]�v�"G����� _WM�|��ڋ��1vP��d�_cp#D>�/:�!c�&�EWY6�2�y�oKj���ALy)���AB�˛E�Sw��܊P%��y\29il�9t2������c�>)��U3I�o)X[|���Ӽ՝��0O
j��6S�yVut��k:��3)��o0�!ή��]1un�TdS09K2;�8�Ћ�������vq�����L�w2l���h�7݅E\��jJ[C zUb��"r����8��,�`�tKhU�Jt0_ EDؾ��.�]�Yrv�7v���(4_!��jRp�0�}.�a�|�%��ɖf[n��jjt�*�X�x\�5Jw>E��}��Z�]!Z���+�)��gP��9Xo{��7�鍄�T2��񞾋���ڎ�G��9\!w�ew�=޻��̈́%y��'Pǆ��}�ӻ�y�[h�ـJ�:�(�4E��ǧ0�����GX�0 �Z��] c+x�8��;Ȯ�i����[�Ū��e���Q��A�\I�iv�P�Y;�^gosٝ���v��U]�6�q����~ ����R�-4���QE%P�Q@PQTQJ��UAQLMSEP�KCC�IDI�D�4�U�APPU��U-��J�KICH�QETP�R�CT�%�T$@RSUJ�U	LT4UTQ	MRS% D%,I@-4Q�IT5E��B1)@R��HU!E4����	UBU	TDR�P�JTAJEE��5D���UE-$@PU4�5IAKMP5KI���R�HEU!@RRU%U]�]�]U��N/���θ�Tu�C/jR�x(h��sY�y�ٌJ�͋�s�*.�,^�=�\5���ީ��N
Ӡ�������� ���]��������r��6���ر�0$�eB�lQkS�O�8��*��!�ͧڽ�AM��=*�P!���p�����K�ڇ��l�X����O�=�V����'d����0�u�8�uм�Y]�ș��h��x��\~�j2c��Ӫe������GK��Z��QM��\�8
綝��l�Bn|�y#�:��>�~=�xO����Πbį��Ћ��`���b%f�JU�C��!��X��ѷ:o���i��3�w1x��^�z;�myS�z�	��4�-�|�W�^Bu�=�݊�ªh\+p�`��\�ϝ�⿩ˇ:��!9�}v8��A���]�bu�&��&���-SV�kUq�rɮʄ��R-�������&5-��#n�;�������{��4;P�BX��U�^Ji�����r��D��P�X�F~�ƯpZ���c-T�6c�5I�e.Ή�QԦ2�Qj`0*��)�����i�w.j��<�q�{a=X��[�_8dl�]°]-�ܽW)�����,��-t��=�:Ue���ww�����)�$NM�E�V- �$��9�{V�q�B�P/�஀9�,������Z�;�ġڷ§WA��
-%y�إ@���գ�A�;3��|.�]�����N�oռ���&xߥj��H�uHGH`��o)�(t�5�����S���F���[����	��/�q��\��&W��L70�5�"I6v5���_���d��������\ft�5�J���*�����ˇ�	�P��F�Z�8��]����Z.�䰯�~Е]ު廒�XC0�2`p�;%+Z:�oD��yz���-��Q�]��$��#��墓J�Qȟ�ًoK���z�f�6�R�Nop|͚��%��mL�ۺ��S��3�A�̬��i�"���F��|�̿��r�h���պ�m�d��/�U��]�K�/:�-��}��S>�c��T�ye�>2�\����B<�'+|�V�ׄ�l[��I^l9�yt�1����.?U������$q�׵ؠ�ܱ��9M.���ݿT�r�tkRF�Rރ7���R�~�}U�(u-�P�U@_���:'R����״}���	ȝ�$�&�$���.N��
n���^K����U��n��t������e�T-�,��&(�'T딬�������/lpp6�f�#_���zIG��rN��;�-^�|Ү/��,q�WV�zV���ۗX'K�:����޻u�1"x/Z=����:�dk}�uߌ�L�=�x�6��5"8��$�LΧ/"����|:*˾���m�S�mq�x�{>����W+�jg�Ze��aN$t=5"MG��p�LO��BމM����8�I�����L�o�t�x�g�q$�w���W�,[� ��ꭵo��iO�Mi{�b2�i�o�>*j�H�}���(z�+�M�zR�4�kc�R���oώ�3=�؈��b���z��2�R<eJ8�l�Y��+�����X�4��i�6�M^	ִϏM�`9�=jb�]����"7o�_� g�o^��M�V�Z@���Jꙍg��צ�`�6���p�J]x�p� u'�;6����Yjg�Z8�1�!�t��[Ȏ%����S~��ݯr�(��z���{�j잮�r[���=�B��nT"XBy夅f���y�7�^�exo[��[ؔ��8^�t�_�E�V�6�������W<��-Ӈ���W�7��н(�4nZ��v*�Ѽ\{�}<��?w>���ҠNd���렗vp��V�&�]��9���JP�x$������`c����x'����k�z�[|_k�3VΛ1*�T��&���j��
������ma���jRsYè�΅>�<���LN��)#�X�ݒ�<h�g�E�X:�.�O��f��F��ۇ�y_��H��
��Z/������<����C>�,jO��X����],��J��wnAz�����c�0�k��q\r-��L��wy�f�+�_8,o���:��}yѭ��Yܸ�g�Irͫ�d��]�Q�m��O>0�#�2#����n;c��}M���ud��C��e�grђ��OR���$t�<F-p�/W{��t{�>�Y�[�z�3˵(/��`�aΔ���깓�H��#�zH�'|�bL�*��e�������M��M4�Y�if];��jP�ޕ��uū�t��Pʏ�	���߯���}�óR�!hB{j�Ԣ�Ԍ3���8귐Ϟ�s�4��x]ջ�.h�7m�J����+L�U	b���w�V|x�)�өEO;��x�i�F6P[�Ej]�/^��ﱅ[�3QN���3�G��ӛR����Y/�%���畼5�F�nڎ�];M�P?^ۯ�m�Ӣ�ؙ�����m�����܎���|k���hg㺏¨BYo],ݳ�wU�	�ݜ��݂���v�Xc!�x5�%�إÇ�mD�SZ1ޥۜ�ܳ�*�sx���z\����$xf;�8���q�P�֭�C�v��5rP�L��L�M(�L��f�w�,;�V�+���Q�S�N�V>�3�xO]�@�#�E�S�Q#���OԮ53IY��=�︝�h�$��y|�G�+0s*E�kQ�L�w��(�$/um(����ss-��1S�Զ�@�U�P�Ro[�r-[�0#a�ȃ���
g�	B�Taχ�W!F�r+�xJ��N"/��uKW�	-A�x-�ΔIw/����ok���b�~��ǼHލ����ڀ�>!�������g�F3�>���*��r	Fi�����ip��F�}��u�x:�>���3ʥϓ[��<2n9�D�T~\����{W�h}�����7���$\�~���w.�U눌��FY�y��/N��G��]��5�+��X���i�/m��4p����D��>�+�Z2�0&:|���=̙��ظ�"7	��:���묮7w���5�[L��Z�Ş���r���y�]/��K��n
��?(F+j �{h�j��q���<��y^Zij�/��$E�y��s8ǌ�x#J�u-W�^wo��8xf�~Wo�œi���d8o��+,Z)��Iٱd��Ϋh����G+��(�ޠ��D5�nK���Z=�A���/]�f=T$�m�>ĹD���N\9�-�	�g����Ǔ��礲,�Y���O���bKG��l^ m�;�߃�Q_�NBoj�ws��~ڶ�K�?(�ܥR���ֺJ�M���^A��N]���ȑ��'�tUשFZ6�H�����=I7�=�(y�9�V��hjZ�`8T�ze��j�X����'���_Y�[a��x�Om��	�*߯yY��&x߄��\�F�RW�H`�A��ar�%q��v�{��(�~ﶳ|���sW��c��v<E���-��O[92��G��	�M���l~U��$���!r�o��x������*�A��P�X�L]�2������!�j�-�a�[�[��Dy����B�~��GP���_�Yk3�3�,>�+��W�����io�fz��J�X�A��r��ZIg�)�T�"�U<��O��Ň7��P�%ꄪ�}~ې��Z`�]�8�4R���<�Z,�2׀�U.k�
�E.�.��=�c��_�	�$z�;�ma�R�r;��xyםK�[����z�5u�&�Ϸ�/]����ta����w�'7�;^���O����{��܎���$�ǘV-�
���B�;xM��H��0�엓f���7�a�xl�O���=S�tU��MXt#D��'c�}a�X�޵�p�2��c<�{���g�ז�:�	��c^��be�3�\��ǈ��az�t������/����n��ٜ7_m�U�Y87�>5��׆�Ű�cC"M��ig�������~9*C�u��b�>��ȓij�+�U�c%C`?]�^�"[c���f{����<�eb75�~����mؚ}S���Avl��;�.X��[��������l�wۗ[�n��v��x6Rޯqq��c�Yj+#H�V)z�KL߲�5�a�4gO�!rY��^��2m�Q��C���5Rm3�t��eCj�1Z�u����e?oX��w�rH�e��yؚSJ�{���˞��_�6���O3�w�N����|AЄ�k�'���}1��X)x�W�޷^�k��Y3:v#Nv(�+{���2�z��V��ݯ���e��m\�tO��K��P��iv��.yo�ִρ�-�y�S"�(=��j:�3�h�7��"
�\Ey[`
G��Y��i�2�ͼ����6��Əg�c�$W?[����ݚ��J���Aʷ[��T����s6.S~pNڻ�X�)�3ϵ8�	���m��한�'@��<��5Q
ܣe��]|�����jh򝗔��v�<ɡ7��-.�>T~��V��C�ԕP��*e郗����ϕﺕnF��n)����K[���ѡΑ�].^�~� � /ǨKD̺�Vi�<�yV��/O{���(Q�\P�`�/疒���:�/>���9{���v��\Ζ^�g�QyX=������U�M�=G �����Y(?h���v��9��zۮ�u�`�����5�����O�>j�)�](�ϋU��"�mz���{)��X����.�F�^g�O'��v���gy�+���;�Nzn����`m��u�����{�1��
�Uabz�~3�e3~��C7:��v,#G8,k�ą��R����ͦ�)��ˏ�k�M��\9����<��_)����-�������j���ݺ%��X��՘o�q��ʋ,+�I�)5\Ur��M�p��`�cz�x���E�*�fw��a�҃���unN�{�W��|n��k Ң���/��'����1�R�����f��/�O�?T�~�5e+X)}��o1�Z@�[&�5���T,D���@\�x��i�7s�� �WĻȅ�̔{�%����ھ}|�v��p�{ۑ��VY��ɪ&a�^<�^���״'6�"f+�ԍ�Tޜ�}��_�@C�)�v�e��<<�?i���V%�Asc��FF��.b�OR�}՝y���=gG�C�APP���ҷ���i{���8K懆�C�gq[�m�v3rr[a��շ�o��Q��.,��I����>�j�J)�R՚�+�+��^�&/��l2/����wh�$X�+��>���ꏺ�l46-���?	��r�þ���oN���<o�휥��֬4Ht��5����ξ?eg_��=�&4릆6D���|︋3�Ue���OIXt̗zreQ`�!˘P��jx*$|:����ߧ�����n��޶�8�M�9c_���̩��(o��&\;�OY"��H���2e��m�^bX��,�|�a��inm��'Qk2t����dA�+�p8)�^U�L�E����w�f�qy���#��P�������Y{�p�t��廊B��cE���)��
�d��xo|3��e�9�����'Z6}>�@T
��t6[7���/W���ElRޢs�ߴ�7×��I�bb�=�r_�w��Y5��["�m�'/G�IQ�e�J�jv�H�b�u�|n�Q�l�lm �Kk)i�q�D5;(�]d�S������g�PhG6;���ù��Yw+n�f;�k�����3�����ga��Ko��Z�:���J��v.8M�Ì�_Da��P��U.Rb�]�ș�W�q����Ϳ\Y�H�}����0:=`>�M�:��re���z����2R���櫭�7*g�v�O��W�?S�:�j{����W��ܼ�*���~U�g��c'^�0f�z �o��V�.���r���PT��ya�_n��G{ļs��P�^��w,a�����9�铃��"��m����2�m<P�B�_nˑ�z6��*w����m�6eu؛bu�y=��ִ���p�i�Yd��K�+䖏/ .�/ �h��ev#⟩�rv\��BvL��{�MN����,{V|o����T�P�j���Uû�#y�3���ܮ�s;L����E��;�߂��Ã`�7,��
��.�[ʮ.2�r;���wY�ў�
��}�-��p�zu��{�ϱɞ7t�e#_:��t�	�S�����5S�����r��2�e�����:�KC���K|����d��V�q]y�7"Ϸ�y�rxifZθ+�8e��<���t��G�>-q¡֚�e�"��Ab ���V�]����[r�m�g,P��9�M�ݎ�¨ի�ҹ��:Ļ5�ugEX�qد7��GaK����K������ee]��q���q�t��vcT�V���&ȸ��b*]�{�A�駒��e[�>o/��c�z�]Daa��O�[9S�Ov�T�w_K�{�j�8�/�E�)���œJ�����t�"�ˣ��eV�m ���+R&�CN��C\�r3K���i�=g8u�Bmm$�Oe�Y�sga�����u�&��}����ifot��}F]^���,����6�x�/��������/�Sj�w+�@��n��YVJ�3*ԋ~˷�1��lR�W�e�jY�t�Cr��c�)�_.Y�T��偻�s4hKB�z��fK��@��V�vYa�"R;�J�ޝMV�5�m`v�������f����Q,v���]�r�.q<�bUt�3�}� H��8x�z��\ʕ�k��6��U1��6J�=ٙ75�Vֆ��5HY�wݹ��l�s��������}t���m�R�Z&����@�{)E֚ߗ+T��R��#P�d�;�ٛOw(
An�QAiI�
���:���97��I���esn��X_cD�u�<�j��d�3�C���p�"�:��{��j���L�!|�B���ն�-�Wd����)��tT��v��c�^t�_\0����P���-ep�VRV/V�.Gr$�	j�Q�6'Gf�%�eCV2��*�1�1�-�rn	���;od��x��A�u�+o��mp��f��wc��I��ӂF��{�G�ְ�*������뎉|�u�E�.���h�p��y;'$�E<�~{VA%F�t�9Ж����ÇK��و��j��ZB�z��h,�q�f�]��;Y9.]�o&P�P�2Mٝ�{n[���Ei�f����.��rV�|V��;V����&򋝭��+Z��hpĤ��z��:)�b08	�k�R��9wr��4��(;�&P�=0cj��F=���T�	��v�W�m�ۓK��el��2���FŦ�Y�����iM��R���e�A;�Ith�Z���fv�vy5��d4�5Y=����܂JT�q�R�^f�|��+��,v��|�ŷ���MV���Mb�f��Ǳ��eo)/D��Gkm�N����3��
�,�W�F����u:��u��;�Vk�X�l�r��ut�T�$
Ȯ��&�B��4�V����jcK;��ݯ0�޽Iк1�S�<���P�Ʃ#��![G]˥W]Xw�.���/���o,�sF))p�C��6/9�$�N(ލ���tvFu��t��O7DEn���\J���
=�C��}��}~�ޯ|����H�JU DSAT���CT��P�����RPECT�1UU)@�P�1%UD�IAAKB�PE!4R�-P�!D�1T445C@D�ST4��)TĴBQKIEPQCT��+L}���%ER�T	@R�%�P�4)FJ&0S�� PR@�QKJ�Ҕ-%CE@3%1SE
S�%UE5AQ)B�JRdENFCUIB)KIT"P�K@�E@9䴹�HQ�"AA׶3_Q��=��;���E�A74�*f���fM�wE�u��sX�2z��R�����V����K�3�ź�X1N˻'�ډ'�dϐ������1������P�^Z��g��}����L�F^K��Q�����.��	�EʿC���Z�Pf.Xp=����}�� �����3��Zэ؜�����IW�)傥quA}�G"~�]���úà��Ѧ�*��]�[�)@�L�W�r��K��]���h���^�\}�A��M�9a�ugLx=�nښɯyЂ/|7��V�a5n�h�S$؎���QhB��J�~��.�5}3"��G���n@�5���5�kا�L����hߜx���K�}��X�����3������O�K���f
�2�U�9=�땯!I���o���pyo\��[;��O�D�ws �{���)�Ғ�2%�	uS��������J�s0zU�M<�(�^ٔ볙l+1㶇��ˈ+�j��4�x�v7��T��{bN����u~0x{z���+���ʞO�qq�x�{+-EuB�R�E��K�]B�y~�X4}�Kݕ4[C0�a|-5��yw�ŋc�uNL��]�EA���۬�i���5n<,h��7�i[�犑Z�Ww�~>�y��U�gF'v-�Ĝ�egS���������K"K���t�}^EĬ
rB!׸��AF��i�9:�7���cw�eo��Ul�û+��~���d�g�^��T7�Z���A�#iu�(�ӂ��B��*ݐjp]��dQ-zj�����GOV�c�Ƨ,�e#�%�<F��K��h)�����{�۲}t	>#I#��T6����&g�Z0���
92��^S/.�,,i(uOj�n��鹚����4Ml����A=`-�;j\�НkL��B�s�z�\FJ�zVe�M�g���ڭ"��|�i��(��3Ϩ/��צ�gP�=�K�Z9�ϡ�iv���W��Oo���+���bs�1L=yh�:E�b�z�s=q�{Wk���8�������>�i���M����]�ޔ(�7��0P�ZHW��q��q�
I��_�����J^�esG �_�}�\��H�N(^EV�9�#�J���f��&���'kRy�(
.fo{�Z}H��Q���y �q��V�4o�`ۂ��҉�O�;UKFLW���z�B��3Z����r������mn!�\��gϠ�V<�2�F�έ���Έz��H�3X�"wR��NC2����=�η�;o+,����ڝR˨�3�x}#��j'p�)�`^6�/�U��R{�b#��zɺx���c��������(�="��,�U1�g0,��:ts��8�i�C�Vkj�Zc$�ˆb޸q�C3y��׼��Vt�&=AP,,OJ+��Ϯ.뼓��R0��Fj�ؽ#s&f��Ӫe�>���
�.�x+w�������#��<2[6j��b��rb���v��޹�[F}{c�˲3�FP~�grܕ��u�e}e�p,Q65]O�D��D��������#�)�jm*�f'.δ;�;��sju�G��aTY�o�VɈ{v�u[����B(yX��l�g;M2�
�̿���R���>������=|7�p���{d�1C\fUQ���`����$�(�}6ц�sj�sBt��w�Ի}~���X,;��e��̓�_!���3_Lʌɖщ�㰹Ԣʫ�ꦈ%z�<�F|�#ok��@ЍfHl2.Y���ԋ\\Y���T|U����g�Nq
���᳘�V>�<ld�7���B��4Hn�j�<�{�
f\�=Ǽ�y{-�gF=c�*������t�8IXt̗zs��ٰl�:�{��U8�R������n��5��x���߲�4k:�k��ɬ���Zf�N�e�Ǳk�̡���bH ���
�2�<\Ԁ��f��a��=p�]��/uw_���~���8p=�b"Yi�wK��RDTs*�*5]G�rW�m�ۇ9o�<^�Zd�Z���W����Y���C#�5�V`�j�\}7���.��$d�w.,=ח�B}�,�D��U�[�a�޹�Qk0N��+"�]��
g���ݎ�I��ew{�/;���FƉ[a����GE�KǆU���/�M��'� 6����O���u=O/�V��*MQ�}��(�ܒ��s.���^SQ#F�S>��x��چ��5Vu���3X�w��L�{�����I^kR��GU�T6R�9����E�n�3����{FIS��x+�y��1��q�IL�Ҝ[��{�Lo��)g�d�uM5w�m��x�c�|�46��`�������;E�=(o���q����9�M/5.l=�|���r�R��Єo�p��89�`��f
w1x��z;�nj��MO��g|ι�G��k���t&=>K�U	5pP��h0lo�r�>w��9p��˫�F�M;�/��=�4�i�y�2�#�Y�[�Q<��M���4\�k�����{��v�Y4��q�֥�xȏۂ�����]Ӎ���[r������m�R�si�\,�Q72ʃ��:;�h���ؒ���)[\7t�,gÓm�tғVo�v�����j"��/4û�ӄ�E��.���$R���un�R��=-����o��;oV.S��#2���,{V|o��՟%䡰��h�/n]��Ab:1�#����9A�����0/ҏz/��k�����Dx�KR�m-�Mۜ8��Euv�~c�W]��sjZ�u˚��p�zu��[��+6�6Ġ�KH��!e�7Ӹ����|����b���,?;����:̡������W����73tf`i�C����=�.'����9J#K��
�Ϛ�6;�%^y�^����lo��1���g�}�wbͺӧ�&]��t��t��O�.}w�<:�X�&���S7��K��'��g;��a���t�0s�kF,NY��l	������ʕ�U��t��Pu�۫wWA5�M�Y�p��֘=:�+2(^Ev��(���R�a��P���T��y;���zjl��X�3}Y=Zu�/��+�L&�ЍnR��r"���M�l�vfݸ�����E7�7e���nq�Wx�x�<W���s�ѱ�#�az�t�E��e��޿��ٺc�^Ѭ��u���M��5i��X�^q::w�X�6S[�0p�'0��R*>��t!���;M�8aU�5ଙ��{.p�g@��A̙�Pmu�dN�sq�����޲���C�^�G�ٜ�q���-;�����4��gb��Z�1e��o���;���w�4���^I�]k^B:���/\O����r���+[}}}3��q�\0hu���8})-�%%�	u<�;�P��@��[�U��սr���콜�^���q4�J�upǷǼ��e.����e.X��U�/x��ޕ��Y�q���[9��3��3��9x�j_aq���{Q��Q��A��%��KB�L�\J]�	<��k���:����#�M5"Y6��s�O�M�t��L��xl�顀�_OMY��؝̵�������5н�����m��{1kaUJ����q���e��J��c���h�<g�Wiq�#���]��u�i`;���N�a���
92��Z���U��}���^���V9�����%'�¸C\����6�u��.��Xw=2��8`���Ls�<{ݭ�4{�h���%l2�����Ao#�_�p���dnq���si����h][�3��5�qwt�7�
�~8zJ�^�z�!g>�S	�A��-�"��:��}wg2y~���y�F�F�C�k2�"�a�*'-��:�S�YX_��[O$��~�t�Di�-[���z����3��{+Y����9ir�-�P�@5�(����}���u<#������a��Ԅ;������
�����6��M:h�'Lr�����Q�ԏGEjv�;�j5���~]������ʄKGt�ejI��˺c��Z|�_R���Ga�7c]v;�\/�;�K�tf)�
���>G%v�Q�I33��vE?5���fP�1JZ��S�k�vz-��;���"��Ee��@L�k���t�U���'�k{׻w��-ߪ"�^\X�۞����ߒ^+���0oK��X�K�P��i�]��B��˛M�0�-:�����ۇ>8F�0���LG:�&O�Ψ�dz��rm��,���z����7���ō�^��e�_'��x\6�wQ�[N�b�w�)��{�����:K��`Fۇ�>��f9vG��C��ܴd��Ou֬թ\YK���Ђ��⽛��O1Db�>P?����ڜK�0S������g���[����EX�;���Y�	��T~~�jA�п����@B�2�8;M2�|+K2�;��jPÓk�U���%��̂���f��e��kMC3ꭵ0R��&��bW��QE6ч��P�D$+lgt˶�6>�E������/��b��.'�v������G����^K�I:�ұVC��+��Q1V��Mޗ�x�W�lj�,��at{�E�Q��\r�'N]�]l+�u�
��Y����R��w�8pcgf�������^_~�~���u�C�b��>y���Xk�Ԛ �1U\e$G{��(3�O+͡���X�L�i��Zk=��)�C��ƃ#��CmݭG�,x�.,�c�sc��G��y�o��y��2����<o�������Z�ڸ���!N:|9ժklSK�?O���)�'�}�דI���4�^��q����%׭�2��\�P�[�g\z��^xc2����AK<�P�z��҆l��b9c\W~=�T���(o��2������"����'�1�k�g��$��&Uґu�˽��PN��ds6��z��A�E�39o?X����!��a�p����<�x�1e�Rm�'� ,��0K� ReM�]��>��赣�t�˸^�PpBJ�?Ww���+��sBs�]o9Lc�4�kL��IX��*ܰ��c^KzQ�n]ß?R��C~O(��w��;ܶv-a����B����ɝ�x��0����j��D�O�tM��mx�ք'����d�q�?4���(���e[V� Ѓ�̒]Z�-بv�ywλ�!��4>�=s/���;��f�SU�\nW2����e�+����92�k�9���<�)�"�:�[y�0�,s�8��-��F�1��]�ӹ-�s#u�.�5�J�c�ř�`b�/m��~�s��^�Zk��sM�����^۳T��E����aUGZy7͓���`[�����.�ف�<������W�;�!�A[Lͥ������U[���O�T�1.:��-����o��bu�aބ����Ĭd;
w�5|��ͺ�Vx�G��w�/5��[���{�,2<������\y%��������&>�=]��k��q��M_�NB`j[��D�ᰫHЅ��ø�����Z��;��Uz[ܾ�����n�H��ByMH��y�0�V^�]�&*#M
�z����TGH|b��c�27�R��]u�p;�5�gN�h~��f�w�ؔ��H��_���d��u[����G��$�B�K�/�3���^M�u�4�s���OK~Y~ɀ�8��'��w��7���v��u^��H'�/��(8�}��ϗ��S�
��	W�Wg�5����0�9�=�2S#ϲ��<*#C�&�L�����C�;�,_���D��JQ�
�D��&�@���ġ�e2&a�F��>����CPt�gU>�.�{&����^uv�^���v�给`��"�$��)&�V�P��a�49P� Gt��R�k���̥����DCwo��u���)��a�yC3x9�wL}ړ}�����͌7�}O7y���R���',�\O*��?>�m�D����՘�s�u����t��t��Xw�R\\P�j�."G�IK��]��I&x��tN>
g�n��}�/ �k2�ިtr��f��*���B4K�q%�҉���b�R�`�[�=ww��=��j����[�����^D/���j�P��T�Fǜx�E��YmPz��R��8S�n�M�d
�z����x���%�~��i�ɮ��!Or����Pv1G���L��.��H�����|{�T:x����j�*�V`���J��P�u��k��S�x���"kz:�>/�!\��fy6hW���fG�)�e��1e�:���u`.s��qg��ddd՞�[�3����4s��$��fg���~K��-�b_:ȣ>.�h�����鞩Yrw���m>��T~`��v�#���P���p5Rm3����-C��j�}Վ��v������x��P�G]R*�g�l64ҷ����،��akk�O�^z��:�=>=:������H�X{�Z35czy5�k,���#<:C�͇�Y�m���Z5^�9~�u6X�3X����Q�T���خll.}�x2�����I܆WtX�_e�M�7�p�o�\��}�RT�
���J2X��M�+K��3��,��L�x!�X���zk1{�
.<��Y4�w����i��Q�^�*[�i��f=�p�UӸCB�B����
#���ΨXC!՜�Go �+g�b��C�:���n��Tb�8)c��"��6va�o<(�`�X�v9ut�U�ν( �#�9\W�.����4J��w��t�����%:7��K�YXP}��8�[n,�o��ײLբ^�<j���c�*�gMt�R��y� �8u����m����D:oP��J�`<c�i�Y�7�����3+F�x�|(���-���I��kD��\��a��&&��u#��7��㦑���F�ºZ�Z�F��<�{�TI���kw��I��=��0��Λ�1���-����M?�p��٫��x��b�-wI����M6Ueώ��3+�t���;�n�N=2ݼ��dZMj��vK�z�r��Zg`_N�6�m�o1b#��J\��C7y�����`ޥc_b�"�Ihޙ3r�/`���f>�Ф�Δ0�,�����z����mtQ9�u����0�#]�X]o��`&�(@"Y�y�Ŕ�Y��ˉ�ܵZ�7Ζn�����E�y�ozR�,�j:V�Z��>*����Yz�r�\B�����%K�E\pB��5t���IMN�d7�]�:!{u��Ywt��Q�:jZ'^Θ�7e���im��m���.ewj�Sw���gQ������9�+c���N&U���W�����F��p���܂�Pu�{��{�[=��R��G��<���UL�����NU�ʩ�E]u!�U8N��٫�릀�ح�J��[!��իo�
�(Z�b�ŗL��u^�7m���e'$R�*��}թ5ˉ�!�6�N�ڛ����1Df�㎻V�����V�F�M�9C #N�n;��|�;��X�EQ07+��Ky��a+oW[|xZ��Q밚
��e��gT}��Z&��x�6��;p����j�|�1u�]���5��X`v�"M&6���7�d�V͌�-k�6Wl�9/lh���z��Ҩ�����u�P�,��J5lr����m�.�+k
��jV���#���\�u�K�e�l7��_K�8����u�fI�9{
�Y�e�C�\�t�huN�=;��?=�����bc����C3i�Y���m��}j�nW��l����Rң�|F�_Y��΄'O���ˣ]�r����XwP���ԯ�+��9wN�K� oiP�����-R��5桅L�,.�k���WԎ(�Ķ�TXy��&�Н��}��Xw�>�c�
��Q�R�)���P�X�U�9%%%#Y��哐9&@d&T�FK��M �KBPĔ�D�!B��d�@�� Pd�S�RdE�K�d�D���Pd�!T�	��H4�.C�A��4����)BdRP�P��Ҕ�Ѕ	��Д#��DC�����1R�,JPP6bE
a6a�ĀP- ӒdP��@4R�4-4�`�CU	T�ABfb�� ��D|�������m��U���#_P��ۇ��c��GTBo�.ڿ���{rbVd��pi��\��Z���4���ΝsL�S����m�>6�`�K�v#���c���H2:����ߏ��y�ٮ��EtOu�Nl��mߧ5>�P�����?=��Eq��8�ԃ��1���ִ�<��tS�h�������e4���Y룾�i�L����҉_�LƲ�dnq�����;�T�B�ÍN�)��&;P�&�f�	ꘅ�*bτ���:E�t�gG�ۼbi}Y�GW���a�龰K��'Z�ڍd��_��히JZ2�0P���C��l������?n��� (� ���5��5�u]�tS�wF`
b���U�K�=F!��E��쾼Zˤ��N�� xMh��b�巗r �:�.���3�XK�����A���Y[j{o{c2��Q>��zD5�X��d�k����<z���R�
a�#�3��Tg��օ
�m�013�:a:lnmÀ�]�P_�^�}qp���=itǌ�+qnξ\��vq�5�Ε�[�,o���E���}�c<^U���G�m?�+�i/^�%�e{n��3=n�O ��O�6��!�;��kZ��
=����ʣ�����Qce$2] w\���'�^#�{;̙]�MY���L	�1q[}	�}��Z�L�L�V�d&�k�Σw��Z/�m�N��1`zS�1q|��+�����{$ޥ�u��M[G�������`r�cی��%��	�ՃV�ql3����z5��q>P�T.�V;Ƭ�p�S�V�3�������=M�y:���'^ 	��u�:�v�xD�	��48֛��̸}�i���gS��|�X�I��v6�dw-������ss�~�����P�ʭ�2�"�1C�u3������"�|H��=<~a'v���Jf+�N�C`C=.��b���4|W}U\fuDu��eg��}�&U���0���ORjO>ɋ�!�f}8�dX�hm����]H�`�.,���g�{��;gR���X�=`�;�C��ɵ�E9��%�^��.Ո����rP�E;��~�K�ug��h��E���|+���2��h�;ܠ�~�I�_��9��CR*3ݹ�l����9dD�t֥RqL*�TJ�-429c_���=�b�衾E���]����>���k�wχ�d�f�!��t�]yv+�nE�:�Y����VD*ή����^Ղ��Kt��!�UF_jj��k}D�3ݽYK`���P�N�c/��q�GH�7J����g�� R��&S�5�m��t���j�9�70]�
�b|]u�wm��цR-1lN{{�P�p�ǈq�������=�;��ڇb�5�D�ε�|��(:
�����{
Dqi>�^x�:1A׺ǌ��Ν(����R/w���	)���*����(���'�~�o�Uu�g�P�|�8U������=��WY���YG,}25�TM,0lI^kR�J:�r�Լ��}�]C+8;��^�]~�c#����+�q�gm�Gèx����jǝ�H��;�©���^�y�� �&��&i�Izxsg�ҡ��w�iteVCgN�#�����.�t;1+���S�s�����Ҩ�^���@���7l��^�1:���[!��>��Ϙ�������[>�5�do�_���0]�Lt���O���\�*�u�m&�>�7_{��w���&�}\��'�ϰ��ێ�U�L?��<N
k~��3.Y>P�m���7��z�t�{I3:��V}6�P�BsRޮ�({S ֑�3	��.ii�P��NAS�ɵ�V�kco�K�g�u܉�	�y#/���C�a��WrɆ�F�gE���+s�V�Ϧ�X�K�a�34�RI�4�-IO�[�wqM�c�r����҈;��q����XW�c7�7I�Tl�����V_S�.0��E���}S:���Ϲ1�T����7����V����Pz�1���T�2�8X��s�e���@Co����~���*f`���g˚��B3��hз��VU�z��]�kM��Rg���GE��@�aK��B�;��L���^
mïT��Xs����#[�]��-׶	�$�\Z���o" �Gm�TⱾ�a�^k�O
����}ѕ�!�Λ�Q��=�l�B�6����¡�R8:RiX�du+�����罷g��y�j���%�{W��J��<f����%+Z�5L
2�U�JG�5��u���}�j���N�^{n;1Tf+3���쵇zU%���y���^׽����p��%f�k�s�y�����ł�ۭ
E.��8=�7��V�a5aЍn
d�(�w�)$=��fV����6	�^Bp[�T��ʸ����5���)J������'���3��/K흜l���z�Z���g�}��'3�x�>�2k�V��u=�>�Q�L���W�0��C��c�a�ۭM��bp�\����Φ����B}W�9+�y��g2��V#��k�0Y[�Me6��Y�p���*��VE�Jň'�L��u�G}�u����6��u�43,��ɼ��M� ��gK�޸r�w4gwZ�R�ũ���R�]B�9���1��������oPu�96s6oN�u�-��e����|�M,���]�o��aU�-t��zK���������ٵ�k�`(���o�$୦fS����sW�.�s���zו�8�c���mVN��?F��ORdo��k��=�H�ߞ��,na9�'��6�ߧ��=s��6$���y�죋��D�Dmj(hCԝҡ�.�<o�4��f�v#,OX�[}�r}�g�< �Y��˻�.�;P<�]�v�M@I�$s\.]�Ϻ�4��L���F�,�mnW��K#>��#���F<��^��/&Z<o�f��t�6
���]�ԃ���V]
���m+�yN�7�ɵ��,��ֽ=P��v:ֿe�@�J%©��
	�Żȝۮ��i��=xQ�z��W'L������z�z�!g&T�z�WsF��Dq;J�+�{ٖ�"rޏ7���+p�˿sl��N�)�	yp�j�ޔ%�ʄ\�Bx?6fe?Udn+����y$'q�J�(g����� ϟQy^�TcS/Um��N��|<����#(����{�Ʊ&�����J��ciwyl�0G0{��[�	����Ն�js
���Ν�4F$c����I_}^��^]LќՆ�(�(��Ju�u��=�e>�u�.�e��j��!k9l�f	�
�,�V��z�<�f=�s1�3H/}���h;+���巗r!=�g��뮌������̋�E��v����y4�&l��:'��,��qchŏYa��u�$�W���E!�]���۵uV7�����b����(T����f&ugL'N��:��ë�P���L׽��k��y�Ƶ�Y�}u�(B�?��Te�V��M�×����O.rH�C��+lo��Tޞ�L~��׫��������o]�O�͊�����^���|/1��[���^I�ǫ�l��/AZ��Qd�o���^W�īi���a��KP�Gs��;�f�հVOu��\�=Y{�l��'�*���V(0Bf\��Zu��t��z؉_fa��šJFNΥ��me֞����C7ꭵC��1C�u3���QD�-����6��xo2�7��#�H�9P���C`C=�1�9Xi�2M!���AC&�6ɥ~�x���xV���O�=^�Esϲb��k'��Y���j��E�qqX�N��=/|�/�����RW�Y�Ox��O�Ze����VV���d�gvRL�3ݒzf�-���i���6"��Ǭ�"ɶ22�?>>X�L{�R�0f��+*I)rS�+I�9�3�T]�-pw���.�2k���X�w�!�M'5]3fK�d�ɯ�s������uGg�v�ϓ����(x��׆���/Z�fZ��U gv���[����ʽ|Ǳ/qa�>�P��iG�dx�YV}��!ϋ���𞙜re;^���UB��:���b�{����6�-�M+�R��oz�P��e���~�����U1q7N��G{�3G����z��Mخ�����.T�%����z�5���y��ݽP+�ڒ)��*�{v���@9]�RGG;L�0��C#����5>x�U��v�v�72��i��ǽ�%aʄS�lQkF,�7�˸q���χQ#f�1���٩���j��F��;Z%�O� ߟVT�+ݛfƊɹ�U��WL�&Ｑ�<���:����5G��g�����h���,>�My�$�L��{����M�	�颮t��������`L��/~#xl�{�4ߩC����6t�q�"��枝���*��I|��OO�ܰl���`����J�a�9dWa�`�^�1\d�J��Z����}b�ǙX)]'���\�v�ƈ��kr�5����;�O�Drh�@^�Ø[(�a�r��v�uw�wXKx�E׆T�M�Kz�U�+���\0�v�*��[2�����a�����!n9����8��1l/q�e�}կ2��cP�Y���F�\��a�*��U��UC�^AB�Ղr�\����|$�X�I�.��T�d>���>�Xdz����7�J�Ϫ��2�Z<�"�/!�ya�^oML�gP�=�jg�-����)�Lj[���Acx�ʴ���XHXwkrn2�����yν�y��ǳ�)W���3]܉�	���F_��y��ð.��a����U��b=���sD�1+K��K�<�qyt�3�r�)����F�������oյ�$�m����lfEِ��UJ�G�;���0h���P�����L�sW�
mïT��Yǣ)=���Id��Z��������Sy�{*���o�0�5�:D���/��(8�o��y����M����w�o��ⱕx�ƨ^�����¡�R8:Ri_�L��d3�y�P��z��f�/'K(�=$�r�N�L�Ev<p	)ZюX��O
��RJ��H�/Q�ٜtb!ח��-��u��0�}�m1��J��/Wl#���R��v����T0AW����s�C�N;�;�����ݶe뻡� �߅�ۨt<R�І.�Y�4��{������n��S��fΑk�k�W�4.F3��R�Nl���n{��l�nvk�{�N���Ls���� �R�}����v]�uAi-t]�@2���Z�^_�ׄ��\2���2�7�a��j��6��${�՜�g�bO_�S�2{��/	��C �^C�p�C�V�i2��RO+xMx���w���t�G�
��d�nB�m��w�`��R�y�J�ۯ�,�^).�nxӴɮ����u���t�-Rt_���[9f����և���6r���1r��Z�]����J��P��8kp�Ƚ�gu����]�g׵�m�Ի�����lO�=�WJ����U���G�q�b��1)<�ܼp.�S��OH���V�g
r�?��^�8�W�ɳz�kʰ�˲��d������l�";�
^��Wi�ðӉzjD��#�s�O�M�w�:�[�)}�1�^���:�Ys��^B��B���Cg����i���g��2OX��mYPw���u�wU����s59d�G�R<|����?�����m!�L�}5	��8�ޣ87�Q�;u࣏+{��2�H�Υ)O�d�W�k�A5��nͼ�����u���-���"a��Wۺ�ix\ţ�uu�-3�(��=��ߨ[Ln��L�0�����G=�=5�L�7��eٷ�cݑN�]B2��l��ڻ;fd��v���|��\]h��N�Z�K�%�듬���W��5\���{�Q�]���|�w����i��,d瞵離��fŏƙt�;���K����$6�u&�+�?\�]����g��3�9�Ԩ|��^_�ܬ��ꘅ��SO
�Z����M�^7�	��p�O�Ec�o���tm�3ǁmF�K˅�Ev�xJ��*oh��z��F�mL=�q��!�nZH{J�"�=�p���� π}E�g���b�����e�ϕ�S%���ˇ��3-�PӶ:��o�З»��'�o܈X}��ZE�;��oC��������K��F�*��ҕ�JV�5׈z�Jk��xg�w�~&����:k����o)�{g�:ƥ��*��0p��Y�	�{�p��0����T���[����fo7���w�;������׸�>+H��X�sX=+�r^�E�ojb� ���H�ʍ�N���4��j����#���"�z�zWz�g�n2�}�&w-�[�ƻ�Vʱ7�.ϵ�[�PE�[YK��
�Wr+��j��8�}{l���>�,=A������4WE�\"3�Y���tr�ܡ��O��t2-�3r�df�w�ԗC���5\���=''I�V�%	�N\��p��sU������?7�֚��Q1�_ P��ö%'g-�ASÉ�F����0,ɰ��j��1�w�끰�������A3��菚���)vUΰ�fM`_#A7-��=����yi�|I�qYb��V�T�����×J��$�3rufAb8�M�`�U�*µ�����V��u�}���9-n�S�5�7���ve�ٺ��vq�<�3�:���$�	�-�Η\�:�u��M���ͽ\�Kc�(
��7�H%��v���zھ}�g<V��_�y]��,���+b�BܤpT��|�d�]2kP������]K�n[��-�Z���$=��h�O��{������jv��2`���M�9'Z�Fk�H���{3"isLb�t��UNU�]�C����f�S��Zc�Z���+]�1k��:"k�fk5�P4�ki�`�{ �绔��0^\N��\�iK��������H�I��k�[�"�@R����2�����n����CѦ|��m��j�<��GY�>�:��ZU��� 2��4Fbƨ�}���[�d���W3ލ��rlA�'��d}[S~qA��̃P�*oH�M�Vj��L��كU�.u����/[��0����&IЌ=��E\�
<�lu�������sKB֌Kj
Y�T�-���j�lZz��q;q h!�#�%JÖ��F�snQ���Hf�ަ�h����y�9�_qφ4��KZ����ֶ���m��[YwRtQ�]%$�m!X-v�x�F ���h*U���x�L�����͈�V,�����9�pf�:�x0Gaq!�Vx<�V�eJ�C��^N9f�����*4q=��*X�I].NK\/�p�KU��X��NȬ�x(<ϓ5��P�.	wZB�w��5+Y�]��V��j�U8��s��u}MNPv
C9� +��u����1Ӛ0�Ϣ�j�nr��5���T�Y�Pv����]�M����Y`b]��kv�z���ͦI�+W�p�j���t������[��'5�՜!X�� r�i��@5�Ɂ�Ôy�7�����H,ū7U�0̝ʹoOj�J�k�E�M����#����y���c0L��%	�B�hГ������5:1�]�0>oJ���¡ɛ�.��S �&���iM�S��t�YJ�R�y#fM�Hb���̭�6��5��"��NS� *��f`�R"��[at7� xt�Y�p�F�OdT������l!���q+���=W�Wd}kVY�:һ��t�Y�&vfD(d���5g��\�-���<E���ٷ�2���.����˷Т�z/�$N�;g������Aݶ[gQ�q�bQYF�E����X�i�7Wj����z:�i)ZB��'%��ZihL�j����l�$B����iJA(((R�i2L��2�C3�i�J���R�)22C!��$�2Ji"�,��
@(
rV���\�V����2B�W&�(Z�2�L�2@�(+#JS''%�Zh�,��r0����B���rJ��)�,���hJhC$ʂ �)����%L�2��'��Fp�P��BfM�]\Y�rÒS�d T��d����X��	S�l<��N�������9K+P�P��oYӌ�y��~�>�늱h�z zj�ϩm�a:�`��2�9�i�����j���Pl�:����=
Њ��_k���GO�FF���{�}*�U��R�U�xx��1��W��~��u��]��4�r�=�x��Ψp:��lW��'@�?�#�P�����%Y���a��Ŗ���p+#�m�e`0�)��N��<�&/�5�8�dX�hm����E�U�']�2�v���}jPZf:�5݇�1?[�[<ld�7�2_5�^0�V"$K�	D�{v��GF�0rĴ�:�`�L�)�,?[#N'�ë���q�>�3�ph�UvX�y���~�νWjH�l)��5�.:���&�M�������m8�ϳ��~���:��a���q�ù���ȢH�t�����˰�X��r)ȵukI��ujٞ�t#>��;������Vx`�C˪0�?F�,�ċ;-+<��-��e���z�^�����!���%aʄU�38��`r��.��Fϴ�LO}��2������xi5r���tp�$M�b�^��B����罪^vl���mR�bg> ���G����ݾ�Zۈ��ԋ7a�_T�ǒjw���a��n���f�$<���%�̏����^U�6E	��| 镫G7B$�-�}:��[%%�6�=�Ok���L������\��<(S�8$�5�xt��n���Sν����zx�I�D�P-���0�g�y3�;o>�1��k~�I&[Ҽ�\�٧�c�X=S���R+G�JmBք'�ϗ�hp�/Mc>�k��u���,N%P)[���"�o���=b������5�c+0&:%~2/:�����T��=�kV�B7���G���;V���Xgܙz��\#}r�|rx׍��5e��[j`��R�2
˼լ�o\&��v��q�ޮ�NΥ��_8��̇�Rޯ�;���]Y�{R���'蒯F�w����!�}��
��V_�,���&�z�l��yъ�S��Է������m���u>�o���^��X3��\���K�Ա1ґZ=>~lw*�#Ӎ	�ic��l��Yc`����t?���n&=O�G��|2�^��Z�ϩW���g˚��B2m
_������wz�f�'�g�s�v�<�vû@�<C�jz�v2��<�zΟc��m��E�n��ޑ�����o;F�:g�$��kߺ��~������^x��z`�0[�'�2�*�c��0: H*�9u(5W7,��N�2j�R�S���`�.�8��y3�@�w�v[�<[�,ңC.u�TD�`M�}g������GFN��*]@�_�e䧋���=d�`L4M}Α&�#��qxo��s}k���M���g�y���ֽ)�~�<��P�X���e�g��e��}ғJ��du.�(ew5�||���5�O���g!�	�Z���3�eL�5C�J֌X���� _�b:�K�z�׫Oq�u����U�CZ����ZÀoK����y��H�nJ^]��ݷ���֬��~���[$�{G����ۮ
�Sަtr�1f��)��k]�2�nu�|s%�xӫ^y��)%�%�c;�z�5+�e֟
�I�^"<�tZSx�v�2=��pI�����4}��G��a3��0)U�u�+l[�֕ᒪ��OU�4{ۘy��loӉ�����^��hۡ��0�`�����g�ji����>�nO$$��wsz�'�콖ǯ\
كu�0|/k�c>���c��=��i_�%�ܷ���xՖT�<�du��R�����������M|;H���r���ʰ�5.j�A�ڽ�ɳp5�:�(�+r��.�
X0>�����Y(�w��[6��Ź(�,-�r�AH��5O�o��������tW��ϞXqMb���s���*��]8��fV�.�Ia���9�gi� �,��Pr�L��ݜ+'vN��Sĸ��x�f�a��qtvhK�̰�|��^�'V(D"��K֞T�+�vq"��sni��Rz��l�}�ѣ���D������q�_:9Ml���R��>���4Ұ��3|�Fs�+�Z��O������ ��l֎èlȱt��P5������l�Ӊ�ۻ��r�cy��WX����f��Q�&V���8i��-6%�&�҈��q��8��N3�L�&��Ó���+?Wo�����0�~�Z}8�ׄ�B2��;�t��t�T��a5������]�z�~;j
���Ca�����.jU�ܫ�'�bpL�� ��[Xb��)ge��]���@��G�]:�^�{��/���O�[Q�������%�8��d$)[��yw�ᅊT*���4�8-%�.Z<�~����ڇEy�3�^^Ǵ���w�GSyL��{lK��Kb�l�,��h�l<&���WI���w"�{��D�w[�Np��g��P����=�Y`ۂ���t�v���lr8���<�U��=_t5qJ��_�f�=P�;1^�k��+��Y�s�)N�+��+�G��Lo4���gj��v.�fg��P���@��^�B������M�r]khɭWgdܥ'� Ѻڶ��&h��q|�H����+;��l>c&��\��R�˓�����b����c�,U��1�#<,������ib���M� ���y��fnu.gձpwy&�z����i��-��+�r^x鿷7}}�jv�&5�z坕��,���ʩ]^3��sU�kզDX���]��{q�3�I3�hg�wZ���˗��1m�oa�x�S��
�MD�Q�g���5e��ڜJ���Nfv�Jf>݇v8y�j��uh��xW��=5qe-�-:�
�ٗ�;M3�,s\]���Ȼ�����+K�����V%_����ǣ��24?���3芭�u*ݤ�P���z��Zٽ�ƒ�/.S鸌!ΨZ����({p	��P-	�.������ܷ�YĹn�<���׷r�ȧ�}:�W<�&(G5sM"},��T��3.l���>٤�LW��p��x}J�9͎�su�C����C����<n�sYi��ޡ�3�l��96r'�յ��}���m��D�6T/ �L��)�,?[#N�x2��`�;ܠ��M�5�SQ�F�N0�X��mTEB�n�n�uJ�i,���r]O1Q6�[��W:��oi�'^���n �.^�`L�Rw�k�[a�N���[��7��oges'��퀻�g y/�x����l���dfp��no��j��(��X��&w����������~�[ŀ�"P�!��Ik�P�z���&�M����j�-�K#��q���:��d��c!��!�F]C��K6�B�K��N.���t��x<��8��Y�����m�P����Y~]�^pU�0��2���
�
�Z<3�0����y��;Z���3<`rV��-f�%9P���c�Z�r��.�ϟ�yFs�ѯ�X����o�V*�ﳞ�wy<a��P����V�a�W�ԽҎ��w�	��������ހ�x��F�M@^i��Ɏ
K~��*n9�]WP�L&�;����[z���3�NU-��d�����wd��Sk�5�	��'Լ�C��֚�}�s5�꿶;�Ax�L?g�{�d]0�Z���N�g��uF�w��vQӺU�Uz,ʖ5X���탴t��,�T��j���oӻ##��Y\v|������χ��F�\v,OXV/AC�,gҒ��U��c�^��fmn���bn����N�qu9��T���ơ���a�����=�Rb����?g�s��d`�Gv�J߽���E](�]9�)o��X��;�)�߶ڐzJ.����3���K�b��͐�k�׹���`��uuG5��JO��s�v��x�eE�V�{��Q�N�^rC�S�5}xð��Yk*����j��$Y�ò;�m��v#?�%c˨�v���E��ΌV"���Է��
�������#~~>w�]��3cDQ(�ł������r�U"G��jFp�;�߂�����|��xi��[����]�v��BZ�4�	4�6آ+��t�3�ܹ��m�=�:��
�7;�އ��	���#~=�*�{�be#��0!�_%�L�C����p;w52���ͭ5��?k[9����X�/�9��}������`�L6&&��$��q}hPq����xMg۾�lU�vQ�qlOSRX��Ձʘ�<'�8'�CL4�t���v��X�J	2-����n�f]���e������^L��IJև(M]<*�����O�vw���+�fIO�Qf-^�%�V/�׾c��7�P����$xk�^Y�w�zV�;y�ɶݦ�@��<֒�����p��낑K��E�3�f��_ݾ�+{�6���Oڹ��3�|�Xy[^1hB�Pd{=�WU->�$���>5��ŮV�h�逸�J��f�o��(N��}e>n�L�u��Qu����M�=���U��a[�6�X�\~ӄ��!"]@81S�v:�û8���� ���O,�����&�[WǱ�Ⱥq[��(9
[���%��t�]��L�{��:�x:�a�k^_�wB%x��L�0)U�u�E���^�\/ҭ��~g�����];wF/XS��֘��Ƨ������Ͻ=l�o�������,xƥm����b1��{�icZc�f0}{\D[c�ϝ���'J�K��n=�<p�43����sװ��o�]N
��E�o����G��	8+i��S��rv�8��PW���d5'����ٚk�X�!�R�ER���q[����N$sΤK&�"�s�N����T^�~�Y����$���{�-r��f��M6z���ƚW��P�e߸p��co�>7�G��؅�������e#���G�Ҡ>�+x���M}G�|�_��}{N��A�q��_^�s~�	�������_r-t��,��͜�/8��U�;���f�D:���N���A��2s���OT#/���m� X����e�hq_=Tx�ucf\P��<h=��O�.k�	y~!�W�����1=����g;Tj��6)9��M?`>,p<sI2�v�Q���;���Z�L�[�0��-������7l���ݗx+S@ˁ�u�θyqصv޶�X��#��N3ڋ�r��¬銯s9P���u�����a��yM�͜�ӷ����!F�.���[�r�}t�����]:���{��/G��'b�ڍg���~�힪����(�x��gZ��vl�e
�
=�"c5K%��h�K�r��]�tW���k)�ȕ�y�w�����)�}�K���!ؑ��З�
�$_-����בd����٢�;K������H���Y`ۂ���,����f�A��>X�}�֘����[5<\=���uXW���r��v!��ƥ��+�[���Ճ����ۇ���M�t��n����1������9��f1�{��x�}��9�,��(p��%�5�A�ڼ	�n8����=��F����+3�L��V��~�2#�}~3�#��v*�x>����,��#�B�g�q&�aѶ�p�a�\zF��QeOqn��سV�� k^��}��k��G���nLs3y��������'\<���禮,�����WA��2�6�Zg.�x�LO+ެ�wӫ#'Y� �z�;�����V%_���q��J243�xz%���`ʗ\�V� j�;ENnx`��C8]jR4�7[L�^��Y< ����c�7@��կ�DPV7%�K4�QK��UdUkOr���
�e\��c�2�M��zs��ǚ���������u��/ө�:�����vuL6U�m�S�w��<L靝a�˺%�����꺱���i\�QE�ql��R��Ვ^OI�DP-��<D_M������Y��y�\�i�R��f]Q��2��覯	Ԣ���1B9��hq��ǅ7�����W���H�O��"�A3,c�/ wa���p�7��x߲_5�/"���B�wx���a#� W����rL�.�^P�e��������~�9t���a��ڼ��wq�բǶ�3�<�k��C��_k5�\� ��-��^~��b�mq�{�U���y��%fx����.>�(o�ɗ̢YI��t�]yv/%��W��̞��1x�YF��#��`�`F�r� ��WoS�Q�a���=�#dv+�e�D����}�[�KNU��~��gt����B*K��E�Q>;2�]�d�jJ��Վ��}�ƕ-��
�P��}������tc>��4Oo�
�,0o�+�jY�a^����;2���)��H݌��٨�L�T����L���Ə�P�L&�@Փf��:�Y�ץ�H����V�B�������]؝�zj��-�4h�m$�����̵���ʖ�t�W\�N�*�Qu�U�힓5��t(M�{T��d4L�XGi:������K]��9��?�ƒ!
ȏn=j��; ɫщD���뎟<Õkh�	F�V���:[@0Q�k���-5Kz`IdbH#��r�n�'Pī��67�g�b�LӼ�/�7���q�6�U� ��2�[U�Q�(j
�UmL���5*W<"Vm�A@F��L�z:��8,dhT�!���de�P �Ύ5���V��L6�ŬǏ�>ӊ.�l���+��h��z[L�Am�˩��`�^Q{��p���=�˧ՁΊ��P���j
�sp:B��i&�m ��,�/A���F�\s��$eފgv��ET��s5��
f���jV��Ϸ�`hIG&�a���tG^�\�AU���ب_V�{B�'��U�i�w���[5�B������NW�K���9Q`{{x�u�48��k'Q�c"\4.[*�r��擫r���[�X癨�_C��%�S�ׂ�j�M�S��M�M>��]����[+(w7�[��n�+-ż�����

|��8����w
X�^�	�����-e���d�e���7ۺ��8�4Q4V1ʭ��Z��o6�w�u�55����ᅨ����.nZ5	ɥ�9<.H�U�C��U-����� ���j���_av�̙vF歎�tє�vs��~�i�$���mp��x+)���IR�єm��wos�)�ϱ��V)}��a�D9��p�8m9z�ͣ*r�"�"� 6��{n��iͣGkY��4�1��] 0U�wk�d9�o�9n����X���Ϲ��u��s�u����Ĉ�Pd�G�:[������r�̂z�m�TN b��u�q��+�dk�� s.��[Q�-Pwl��ٖ�VK�����n*R�LQt���VC��.����V�����ㄺ;y��q��/Zj��Dtՙ�Du��n؎�pwU�s�Ϸ�����Jk�k�[B�9����%,�r*�VH)�k�s:P2��U��Orȳ�]���5�ӒŢ�i	t��u�7�pJ�Q���]˕��#�Y�b͋&��@�԰�,Ǳ�/��7Z/z���������laU�c:�����9�����W����c$-ʻ��]]s|��sOl��U�*<�kD(ѧ�	�5��!�WFb��3F�o&�#�쭏'�eKv���g/�S�W4�,��%�i��Gc�Q��u��m'�� ;���������{�}�~y1��Ξ��އfұ�ę��P<��8�y��z���Ct��ar����|�I��gs"��[au��c�(��!�]��^v+Wܲ����5�U������b$�r�㯶I���]}�\�ɍ΢TYx͇Q^�!�.S0!:N��	\�K�U�j����@��I�e�VXCB���"PҎY9%	f+Y
�f&@��4+T��E!���4�A�&I��Ed��䔅�BRP�.N@R%9�4�-PaR)��P�I�@�&@��!��E.KBd%�9CA�RR@Rf`.K�d� d�.CT���K����d�S��Y�
d�C���4���9 d�fHيRdP�44���>�
����9[��T&m�9e�s@7�ta��n�:�ܨb����t����;f4��cM�t��nrT3;n�����)�2��vw뻯��u���n��tX����z����|�=�UE�7��wQ*f��'z�I�znzg^۳��Y���_{��1C���0&:RW�"�.:�^�j�ݣD�s��h}}<M���=LW�����^>���e_��+�g�+�И��XϜ��뀼�mR��÷o�j8�
xh0o��&�ϝ��NfC�S�`ơ��G\*�a�m+�y![����qfg{NXZ�;�k�]IK�I;��{+��r��v�7��9I���g|};y�����O�P�'����O�Z9yQz��H�(L\&�2��;����L����Vxp�����^���bm�~���l$���%��d՟muvvT#�\&�ٹW�y¯ޢ�oSF}���V}�<�}(;W2��wh��%�L��T�;4u�r�>�<#��w6u󵰏��^�,i�?zϾ�����O[9�zɆ�&��H�Dq}ҏ1���c	�mi�������A�͉�/Eڧ�L��}Ձʘ�==��ϧ�Cba�Fr�1hU�Z�^��
nf�|��o�N�b�ڸb���؏�Mη5����t�ͷ
}��.q7f�+L^j��Glݭ�:'Z�J���eKy�q+�.HVA���V3�fv��s�s�2l�[�s���8~~��6���1Bҵ�Y�$��]�������|cR��Vԯ��}�8��Z��Pg��y08j���)Z��	�ke
�	��Xq�z����m�}�Uf�:�^Z):T�j��J-Yc��t����]�L��!TG<�ףtg~l
T6ɇ�����d���Yt��^_��U"�k��Zf,�z]��W�4u]��~�zt�_m�Shw"c	�w�O��X�;ּ�X��{(����[T��<<����k�c������o���>�s�<`�&o�j�x]m�x:Ҽ2R\/�
��~���(��O��lꋉ���;ܱ谸������g�j<o�Wh���t,(L��\�w�ZL�)�J�߻2��� �[c��s0{��Ҽ���[�o�l�싻�0��������H`�+�V:�`.s}[H�|���NV�3)���Թ��}Xܕ5ٓ�Ƹ�a��=G���Z<��SV)z�υK�)��S�MH�M�E+�����k�����ݗ�6U�=��i����Zh3ԝ����o�4?������Lg�5��+�t�v�hd=q�z���Ej�]
�V��z�]��l��j�-��*I5]�^�	fn�Ag+WeJGdU���t8�}��]m��
x�-Y����gz��-
ۍ��T�]pm���Y�GY>H[��͑K�)��Lqf��c�T�h�|:�%���N�e��a��o�y��&R=b]����Px����N�mm_��H�m���r�_�v҃W�3}�ӱo'<reoz����H�w�JR��p�r���i��������;ӆ񖺐��u�z�^i�3Ө^Ny�^��F^L�ذ?f=���vzPǛ�z�Y{���؎S2$#���a�΃�O¥íxK��ʡ��4߭z`}��ح�s��y��~���
� pt�ZV)�.�������wŵ�yp�s�3���S�u��'�7:��`�P��`�,<�����"�\�y��7qM5�{P��IB��9�����sސf��:ç��������ܪ"��4%��V)>[uR!���B׎φ��SY>�>S�+�����$VpEe�n
z�t�v՚,�#�;�3ջ�uC87�n�gfwK�>�탙x���{ޙ浺�C7��K>}����� f&udx���ۆ�����sS�B�X��s���i����$�C7:��t�!�=��cJjƵ+��ʿ8�$�QӸ�mok�2�Y����djo&��f�J��]PBI ��Q�:M&�5FLm�QߟR�{/��V�|Uݷ�Vp���6��6�n^���k�J���e�R+�n�񈮶,��~	qT�����D�$�\�֎=�!j�C:���Q3e����[�/��f��V��~�2#]Xg|���9�nL�����K��$/��	���Z2V3�n�X��D�5E�=��%l'ڜK���C㷗�	�p��MD�U���ofxs����u\ڇVR8Xzi��G�G�it��V^aBħz��ʮ�Ŷ�`�3\b���N�(Z�0���㾼�/>��x��PĶ��M�y�)}劦�A�AC�mC����&�0�ΨqԾhxl=�&c<r�Z
�zu��j�;z��G���eUW������+>hz)��N��>Ɋ�[q�Ⱥf�����^�=�(\�^V�#><\Hc��x����9��㓝��/,��v�6[=�b�P�v�$O	v������]L���p��.'�k�X����rj^�i^,��a�����ç��fqɔ�6
�S�_H�d���r�[�=�C_G���|���PdA^��i���>�+����s����͛$�iqX)8��|�F�`X��}��n���� -��*�G��o�¹��7|Tf`� [@.T�aU.���Bݩ\�R�<��H�X�d|<�*�Vf肛�9���f��>�����gg�3��t�+Si̶�E��s��[pw+8�{��.K��諗Q}�̝C�_d�s'R���mzu�#�q\A�WoW�g�(a�eه�F��˔ʵw���T���Jx�U�LvV�2}�0$�IP�rf0p9E�%���W�k�![��l^l��0�^O �$a�a��*���|��poK��AB�9a���ueN{Fx���%t��ybQ�_��:ѳ��O�ʥϓ��g��O��U�E/8G7)���Ay}�ѻ����JT�>}-��c�e�c��=離��ZS#(�+~Oe��2�k|�ק����^P�ӟ}�#���l/���C7-[��;?f/=��<��I��0��˝B���ur�A+ծ٘��/5՟zK�o�_��}<k���SKo8*i-����1ǫB�l��*�idu� =ޤ�X��)��yJ~L�;�A��}�#/D�����t���HM�#d��>�J�ʭ6�UWR��a�I�ޤ[+��E9	�Kz�q���]��-�<�J>�v���U�@�Q���/*��\�/܉�j�����¥�Fʲo-b�� �C��.#ew$�تc��C�s	�}1&*�T�KQ'�ٖ�,a��ڛfl/;[��ǻ'O��f�H�������me��V�v�X���¬�W�E4�tdr�6��/b���an�T鈻��V�0NWW�gf�+���F�c�����klܰ	��XTF�K�`�	lS>�\^];L�sS���:~�<Y8��xI���t��[��+>�x߾��be#���?qy��P��ćb����T�W#V�c�1b�>���ͅ,i�?zτ�����d���&&�:D����� �\ݧ��s��r�Bڏ��y��]�),y�*��8P�-�ʘ�^G�l�Vz�V�FR���yOi-;�y+��J_3��}q~}e�Ϻ�=	y08j���%+Z��^f��~x�w����3�\tD��Du���R��hj�觇K-a��t��\P�bmˮ9%��RWꕼu�N�:Q#A�t�_���m�O����K�E�U�>�K����[��̜�kWhR��{{�/%[�j��7�pS$�J'��L�Z�>�Yg�ʦe��J4��"�H�uM}~9\�N�X~P^ױO"ҭ��h����;	�o��ۯ	�ط����3F!�$�%��9{*^{.q�퀳�^4=�z��t2 �^0y�i`���ݢ����i��ޓ�Ayx�"4߷o�n��~N���3S�]�qmF���t$*���_dݵt� ����ORr��a����|���5v�2Rʖ���| ;~��Dv4v@no]�/�3e($��z���a�ղ�{K�B��o1L,�ocN������[)D�Lw��^�g��xz���̀���� �+ltX�fx'K$�[8�'��l.�y��D�~눛�7Dz͖�U%c��\�9��`^��G�,
�fe9x���׫��X�ޮ�7�b�̳�ݝ�w7E�5���t���C�Ӊ�������
�CM�u�}�ÍT�L��+ydʇ���!kMl:��J�̻��W�&{)ie]Ύ�X��SJg���v#'�i��m�kGa����KЬ��o��v�:��[��M�|��d�}8�p�蝈�`d炎	���p�y�2��bY�k1t�*V��Vm�\¶c�wAz�W!���}Rߑk�w�ٴ �����z���5��yhkkB!�7_=���>ۤl�����eȯ�8�x����p�^��ㅹY����Z���1{�j�íf��m�V�*�:@�:E�b�B��=c��/�D�A򜱾��s���i�;�W@�oq��gOJ�eB,L%���B��䮝q��]���~��[��*m�6<�޺��(�^�*�/�A:�-���IM�ږD�f*��YN�pY�D|���;%��^�����K�[���������.��R��&M��'�m���ɩ<7�|$�J�:��el6,Y���h�s;(9���{�ٹ���y��Kڞn�V^EV�8��;"<&���>[x�e]��:�W�uF*�����r��q�,%�|�$Vr+,pSԳ�N�Vh��k�`�K��[Y����{pAZ�UnK\�佤����G�=��=<,U��`�3:�<GO��r*�w��n�;9��[�0�f�>z��j�e3�m�1�^��t�"�}�����]��ɡ�O(f��}\��e�U����=�q�t&�J�o�O����&��sI]<�L}Y/u��n�(`��;���3����Z�ł�c�YK�;[a1�4q�������[���c-v������>��a���v��{_�����'��i��Ztu��&͞��{�|A|e�p	��iif'SS0:�<sӯ�}y|^VZ<o妡�OR�9����Q���Fuq#}X2�Д+ܡ�0��Q`���eΨs�R���!��3��r�n��o�<��Z`]&
������Q�"��9��W�C��N�,������v��Եv^%�����O�����L,��Z�έPt�N�A�΄�� K���hD;^�9>]�$�fL�� 9B�v�k���W]FTwg�&�npV�/z�\��/*�v�\|��S��_
z�q=S�dڊ���8�IJ�����$�^��3݋n�.���+Ռ*�wkU��X�WPL�uE���?!���چ2�p��>ԭ����6�v����r/Z����BH���W%<�h&e�JO����|�Ϗ��TΕ��{�g�W��Xt�wzs���Ä:�� �5��_Թ�A3ǃ��z�*�n̬�mh�ҎRVwΗ!>�,k��Vg�{�b�衾F]C��K"�"ƺ\W� �2�M�˨�1c~ޮ�-���/٦�^�u�9a�ȃ�WoW����ς��2�Ù�y�;׫t�;^�=C\/�p{��<^�su�ǌ��J���
��1��Qk���ܙX9���]���2�C�7�m�g��L]N�����z��sz]$�P�]��o�,��{�'����T-g��臲�u��	]h���@^i�C�T��g��SG@�Y;4��^��>�0x����T��v+�a����Z�h���XZK��w/�Xt/��}��Q��L�x`�e��u�9�#������x���e�;xl������̉b=�l�+rk���� �.c9�)��F)��Ѿu�F{έ�������D���}��L��e��l��}W�Q�:ɋ�Wd�9�.7�&�7��Q�����}u�_Vݸ>Q%	�	Ok{m�Po4�i(+���٫�~���(XdS�w���^�3�Cb����e_��+-�ر>��aR\�Z�.3��e������9�R�'T:�����A��I��;��b�̇�Rޯ�{҃��[*o]�GdQU��4�}���Z=>~`-�x �m�yъ✄J�9Q~]o�5���S�i���Gz׿ō���P:�%�K���عv^w"G�By!���ﳳ�纴u��"�����|����+�g����5�\��آ+�߮��o]j���m�N��,���׊���N�i�{U��8�����i���(!�IsQj�6�f����Y�3y�b�z�pu����p�Х�"���Y����O[9�zɆ�'=���2v\])_�Z�;ׯ���V�0�8�CZ��A��T�0k��� �"�z�ʘ�=��C����Nr��'����Z��iԚWT��_3��}qo��o�3�g��`~]�6H��g;1�gμ�+]��¡�����JE�eJ�)&s�V}�E�/z]$@\M��׊vgƑ7q�ƺ+�z;��3��T[@����qn�	��³j�Y����SFv�_"�b[���r0�y�Qo�=�1ƅ�xh���إ5&�[�z�v�B�+�4�Y�z�]t#�&�Ty�C�㦸V�%����D1�y��IW�6K��\�d6wn�|i^l��:N6�n�w�a�O�D�t��K)���edTqLlAmf;�M^��f���-VƩ.�:g�e�6�-2h�*̝��S$���S+���v~��FF�,�5��VU���{wu���vQ��j�������j^ҽ���	*Q�b���m�Ym�l�av��U,��t��Y�:�)�������v�S(Ȟ8�'����4h����=\��:��v�E7���n��`���-�Ǎ'>{S8��{�����<��^�7$�JL��nlpv��+w�N���޷sjkM���\1'gn1YS5'Pڊ�d.W�a�Q2�.��������Ǡ��v�a=Z8�UHt��ﷹ�s��t@t�ۦ�>��b-��ʚ�fE�z�u�b�eCq>���h�PIt�R�qe�u.�׸5�t�">o%�7���좧	n��/ikM��vRU�����0�W���jgEFz�Z��2�U���٘����qZ6���I;�f�� � �P�ַ����ʂ[G�mq�Q�2��{��l�aJd��+9\����mbݗ�����6���oza7!�qt��5W1���޻���-��N�.�y���-�.��&�ݚ��K�B�q�s����2���ƻ��ؖ5P�����:�9������X�eM쌩�v��M�I�yС��;/ܓ�^�ȗz��x�dի�}b��VM�xλj�l�j��2���X>�~%�I���;��LM0f��v3F����^<��2�Ԝo���D�F���qm�t�fnR�
�Bf�{bV�|�s���;�E��b�TԨmeYr]f�O(A�CO�wF0/��B���z�����ʙ�q�^T`So;&:عu�k�YO*��{ȇ���u٨⋖���}�Em'�Y�t�X��t��ɋ睙�0s�y.e&�m=�u�ƅ)�]�p�t�LKD�$�s�$���\ָ�љٔ��m$��I�p'�q��'y��h��w�jv->᫕9�gڦZ�����Gn��9w&��x�˫wx� �6ɾ}
�w��5:�\ڝ�%��@��J=F7�םFi�Rݻ|Nk�Ll�r�f�%�.:���A�wvŴEo[o�G�o�u��Ί�����zN�ƍ��c긮��q
@a;|�Whu���U�̒�Z��
y�C�+�F��T�j�a5�jX&��L�ڡGx$���t����ݫ� ��	Vm���%Ď|�kE�93;OVv��˥Fm��li���5;��W5��kz.%�`���B�Jd.M�9d�EHR-T�5A�9`5fd�NKT�F&FA�4%1 VY.f4J�4�يdB�4aaAKf PU9@SFf9ђ9A�BR�@VNNNE��Ee��4��Y�� eIIC��� 乘�ffFFCda��d�	T�.T9eEN@d�-�!5ANMQYAA�N@d8FJe�d�e�T��4�DC��VFNJRR�@D�eRd9�E�@R�e��d�
QU@�e��d�A9�-U�V�fd�YC�FcY7����u��s�=)��ƴ�+�C���U�[���Y6+���\c�:y�q�l�`�[ppֱ#��SBﰞ�Cf�*w�~�l��Zw��w��tH�lIK��Ѻ��<6���^Z/-��E.�ŧ���[:�T���{f�/�:�}0��B4M��I��O��bgzאy��[�3�=�� {s{ݙ'I��Z�:���7�B�O�k؟�qiV��4o�9Љ�������u�E��7^���i��,����k��mRL���ם��nX�X�i��-����
�O��k�"��I��z�_0��̌U�y*~����q-��:�c"pp �S���έ���l�1+0{���mѱV,YK�IX�2�,�`*��R#�=�0��3�~u�����8�>����zRޯ���x�0r�Xn�h���#l��h9P_l�HĮ-��i����u{���ɧ�O��a9�'��6���?�ʇ���!ai��ܓ�Cf�g��;�Ov[��`����sMC7�	،���u�ܟ59��X�h��,�1��]W�Tsv�m�1ZEO�#�WU	,����N�a���3y}��O�,3�㇄���rg�n�I��:b���j���p�39�p���d��Z�v�n�1��	�U�\b�kM]�X]f.���P�G�|]�uLdӓ3�'cbTam����p03��Z�x6�N���]����գk��}e�>�����ҽ9̠�ov<M�TS��J���0UũB�Y�W�u�=C��d瞵��:Z��=���x����=����W���K�s���cHF�����R�ֽ//�p5��ȼO�U͔�㏫z��w��9�yS	�A��4�K��-�o�^�9���N���U�{W���74�Mc�U�yz{�]��
k�τʄ\�BXyi!Z�rV)�ywW�Lv�:W���z��xA�:Y}hq�Q�Y����2V\*�'C��#�J�Tk׿q����+"
�Sv���b��!�pY��|.�P��x��[����Ee�n
z��N�(���{��.�~�Ó��I�vF,���δ�G={I/E��b7��K�,U��1�%�|�<�v�(A�y_����!�ǂ*j��>��/��;����U���X)����$p���^��7�>���1A�80<��'�k�����+��e	��9~�2"ǫCv�h-���Gs��2Lˣ�{�Q^����c��M��2.����T.�]cL�OhKsH�Yۻ���lUgՓ�=���0��j�9}��A	��	�q����_�/:�̻06{*s:�GL>[����;�:^���V9n*�ǃ����9��rÙ|X���Hg��OoAD��=M�}��F�+��l��)����X}\�J������f`�3�:Xz����ܝp��֏����,��������{�-_Hs�ߠ:9 �E� �4�X+K2�����c�>����}y|:(���)gpR��;mC�.{�H�'���O)P�w���_�iE	��7�s��Ծhlg�֨�'�ĩ��5]���o���*��>[J#eqq`U�`��:�]�V����'R�y��Y��dBwYK�y�[���^m�/�M"f��wkQ�+��̼we�wa�	��ڹ��o�b�����C�z�1�<`�מ7�w�z׌.��H�%��aШs�}������q������͙V�z{��>Oׅ�Ty�q�>���s�z�,�A5��X��r>�{�'��z���-��n���s޶�/e&�%�~����j�.0�Z�	����ȢH�V=7�3�u�`���-��yYR���˱9v�u�>�`FÕ������<0�W��Ɣ�0��͝���BV�D!��H�g��.ea~�wK	)!O��`��^��7��t8�z+�BPЧc{��̏��z�4c�E�_�����Щb�̤��fi�<�,K]N��^�P�T���F���ϑk;�:��w报��I݇�k^oS���<�GV��Zm�����v��[�)�[�3���k7t�2�[�mlo�K�������h2��v�0kK���FϦ�*
���������;*��g�}��^��9r�e�cZ���{��kt��un�=�;���,zV�/:<�YC�qz}n���m�"��>��y�1���}0�����H�2��S� 1M��Є�_}�0M}�ڗOp��'W���f{��?Ǫ󂺘$��o�(u_�]���f�w��+�i��ݎᨤC`(rۿJ�ֹJ�@b�<��v�W*X�ya�C�ݰx��/m�ꥬ:�/VIp���/��U��er�3V�$D�1�3>[iઇR��P����5;��t�d<�?$r�S&$��U�[������*4��V�Zi�U�e�&�BM����<��w4���G{�[�]ߤ-�T�K�Lv�|�*1�:F��0����=.io��Zx.]���D�J���=Z=�۝�gf��2pv��_=�7 P�Xs`��a��� K�`�	lS)W�{-��r�ng��R��8-r�>>��Wu�d'�{�Ͼ�x߄��\�GmݠE!���J��?[F��'Ӷ� u�0�ͯ��Fb�T�=���pAb��`@��pw�QB��Vv�c�.�;6�ܾ�7��7�v�SGosI��M|C]}T*���{� ��Y���O_R��i:�f�0v�̢X�L�ǁWD�r'[�]�Wf=��T�\(l��i���^�M�u�4��~����,s��`��a�����G���b�]뢳�%d��$�Ÿ�⿷�l<^k�OT�5�J���EB�8����[mxBS�Yۏۛ����
��xi�4�T��Vgw���>��r�R���7|��~ݔ6m�Tᏺu=_%K�7brϧ�Cs)%C�"��T�"�U3T�����{o��N� ���7|����Cܼv��."G��,L<�;��pu�=-^_�Q����ݸ��	;M=�߼댋LŃz]o�V�7�'�'<U���^A�[�zyʯ+G��=������w����m�k׵�P��W>�8��԰t�Ez�b��V�E1�͛]�vt�+t����U���"�݆x^�bcۖ=|\M�9m,����vT�ª���Ɯ4g�15Wra���`���m�t'��z�ʞ���4��<�.��!G'i���@�R���츨+�yH!���C,�`/��;� �Q�� �u{O��=�Y9�8̀>��z�4't�cZkQr�*��&��j�vN��z��U0q,��؟[��i��43��쳶�P؅.U��v��{;0��kw~�/ct�)۶�J��kX1jG|�Q(�>�W%[��J����g��_�X�o�Z}��r�^	��W��</ݝ�w7E����*K��=Ms��[V/b���g���9��Yv%ۄXNv	�M�tt��eC�+(dQ�cW�7����,9b%d��<K΃P�p6r(�ҡ��،�=cL-mv��MPL�z��<i��]kE��9��ъ7`Ĵ��"Eb����x���ř��rs�G����x8i�����S�-n�h���3Q�>�4M}��F����au �c�Z�O�l�d瞴k�PC��wM��/��^�v����Z�ơ�t��t�I3�A2(nq���si��íS��ŕ����W��u���՜��S�-KZ'�`<�s�ZI�]軇���/s}��f�����^���^(�w)WP�j��
k�ɕ��
�$�}��$��,�=�a����&ƺ�<�{+90	�^Vn�Fd�0����s�>G%v��DCo	�����r9�$9���^�:�>�����h_��=��q�,%��H���ˠ�Ի	��`g^��!We�Eh�gK�W]�
��]�튥�OFP������R�/�~�c��i�$��2���[������$��
�:���ݕ�2,g9�ƏrA�c�8:M��.�`���A���� �[�scΥ���]J͊��K�V-��]�=\D5α���k��qpww�~Z��0oK��X���	Z�s=�
�r.��WK���OS��676�O�:���xe\\�I�쩯!��I�s�cS�\׊��W��^��x�W9��{���۽�^��X�W����c��
vWV�a����}X���m���5���˲=�n2�I3�h�[��]jөTH�Y�JW<}˜�꧳��_��rj�VX8}����ٙ�9�}�Xz����Ld뇼z��zUE��=�p���5eSا�� R���B6̦�M2�}ZY�N�(|��J�/MV�i�}mg3�-�u�C����O��YZ\��mL�C�L!��f%oiEM�a��T-J憝U�s>��SnL��ٞR�s��p�R�hg�2,U�e��:�懢��:�V)�� �d��a�q����Q�͂�#��hm����]H�`�.,���1ݖ�����oy��u����z��c�C��Ny�~�%�^�!t�"D�.�45rP]L��L�:uRom��YL����V��ˣy�u]�12��}h�l�-B+e����t6��GN���,�ZC�^�t�p��m8�d��g6��v�8�6�nư&�S� ����5�v�*�n�r����g7�`�3$��^J��� �Wd-b���i��j����^�e��c�*�v�#N=xwºf��Xt̗zreu�:���e�s�t�=s}y:_��B�e�\J��Cc��J���|�L\|"���p��%�����|����h���d�&�,*���;�v+�nE��Z̎`E�q�Ev�x8*������[�m�˹��C�64l	��\)3��/i�ٵ��wY�0wL	+T!���.7b��N�ꏓ�|�ˆ-6&]ß�^S>�$aՓ�����L��%����)��z^�A;}�C�����>���y�]	�٨�N�*�>Lp��g���5��v�+m�3��#��K&��$�&[ҽ�J�X;�bnR��#�W_b����g%�v�9�Q�vѵxǫ�=��.i�R�W���mw��^9I���9n��O���]F���w��1x�5nX�v�����uR��5Ճ�\#QD׭��]=!̻��_�=�ڶ�]�9Gz&y`{��H���܍E�;��S�����*]�}y����He���f)�����G���yx��k+.��~{o�{�u�������|�2��@��`_`[�X~�?Oz�Ku,�JT+��:5�zd�~�N3$��Sq'K	���㩽�(QdAm��M�z�oZ��33��K�b|q=���78w;�]�E美�U�L?��=>K�Z<�����m����{���7*m�bf�c���yO��q	�5-��3mu@��R,�������T^��-�U���w7��0޴������o;�Vrzyg@�}�0�	Q�~������I��c��#&U�����Ð]K\s�\���#ޝhտ^��q��Pv�e#��@��R�!.m�_d�0����P�&WRg~v�j��M�u�RƑ`9�޳痢�,�Lܱ<�]�*޽���Y�n��?)J~}"K��
-��^k�OT�5�W�>���1�-<�4K�.u���wb̀w��~�4�t�Һ�GR���s������Pg���Vf����~�����n��9]�9Ε���>�̤�ґ�1yh��K����=
)<EN|z/'�)f�C��Zs��(dP��+�|�R��Q�%�S1��U�����,&�
������<`�VOV�ix���tU��MXt#D�$�J'�N�6ٳ]uT!��fYw����Z�� �{�������8h�x�z`3�xSq�3�����9zO@,KE�ތ��S+��oM_f$3Ijt�K0�Qnc�vep���So���gd=��23z떅J!+�u��i<z���b�`���a�̙Zȩ���Ҝ�Ui��اp��=u}-�4�����'�a��hߜx�6_����s[�~�*�}���i�x����V��90m�Bǽ�����LxnX�X�i����H�C��߻f�(�g��n�=88:��p�|�ᒒᄺ����f@}��qgն:%i^��;N�o���z�z^���N&�����[�o�yx�^WOW�ł�iV;&�a�k;�Jg�ɭ��w�/I����x� �S=�S���5.j�8�Ɍ�0w�ּ��H�(�i\�����-{��N��5�@��>H�4ԉgҡ���r�����V�UKP��A���n�Xw�Is73�޵S�T2`|6Dҷ����;�=cL8�o�x>59`)��� }F�\����g�?��#Ĳ��\D�������x��^,���F���lBe���	�6u�^��~���r�_s����a8���-�0�i�6� /|��<�[[��+j�T�v��x�V���Z�lC�֍Z~�����ӣ=�~���{�z��* ���TA_�(* ���TA\Q�
�+�PTA_�QЊ�+��W��TA_������D؊�+�* �b
�+�TA_�
��W������D��@O��
 �����1AY&SYu�t��ـpP��3'� bG����Q@�UP��QT �B�J����R��T��)"�DJT(%EB��*�RIQR�)"�U*U(R*���zd��0�*���T��UET��
�*��
*�D�a(�%*(�$�P�!(	%I(%
���˻��R�QBJ@�P������
�2�(��"R�UJ�*�JlaADH�QA�	!*B*R �YMd��T)p  �]
5Bhb�`e�6F
�XJƆ�U�i�(�0�� ���-��PZ���V����DR
R���DC�  � �Bk,�U�Ij���&UhR�jMSR �Z�ֵ#ZFY@ ��CV�3��l�X�P�j�T���)UDJT��b� �U�B�n(t4@(Xsp�(P�B�
Η
   � ��(t4(P
��(P 4����B�
(�껅
 �*�P
4��� ��DR��H�	(�EUp  ��[` m&
!U�h ցb��*��X�[`R��5��hh�*�(Z�SYZlh��`��U�0�$P�JV�� �  [�e��V�)�jiE �`�4i0)�R�m&���Q,�F����� ҭ�	l(j�,S5*P6�"$J��UU �T�  -r�m���F��m@���U+mI&0��4U�f�DP�MPګ( 4+a6�Z!�`ef֒)U��@P$R�  ��(�i��m����(�iT�)m[*`�5��3T �,QT4�����mCM�aZF�P��T�SARR���JTTD��   ���h�ն��ɕ�dؘ �V URd�B���i�6�`SF�i[@ 3A)�*H *"$�   -p Ʀ( ���Z mE� 	��+lU��20 
�E+[XD (�
�ERDQ(R���p  ��V����ZS
��+A��e e� bƆ�V�,���Pf��V����RT� S�0��(�h4 ���hɦS�A)R h �z���=@  �IfU*��C #�"� c)�d����I�p'��H@�#;�y�㉶{����kmW�{� IO7���$ I7!���`IO��$ I?�	!H�B!!�����.i���?� �+.�,���?�y��MVGn
%L�QÎ��x��7@w��Peh�G+mL�nŦ��\v$gh�K�v�^�.�T@c��Պ8+T�2�i��Ͷ	8��VZ�"�F���6�l��O� j�8<�Z��SVR�&r�����V�ZU��Z�$mq�^�y��A
���e��f�)�GJ��aZ�"�z�r�,(�(e��{K^p�R���Ol,������`���T䩰���v䂣�Ѭ����Ƣ%R���bF=ѥ�˃v�NpPm��6'y*��̹	���"WNͪ�Y�,y���mb����E8�P���@Ƨ�Tӌ=bPR	�fӭ�0���T�oq����q@"ҩ�6��ݵJ�ǚ��v�>w�E,�A�ߦ2ެV�S'#��4J�5/޵Oi����ׅN�cgYKq2kN�5Z�c"��'I"�}���l�R^��V;l=%Sb�XJ��*%%��ө	W��2�Q� ���V^K��t�A`z��S	��2�hm���z ��j�������!�[)+A�+/``�6�;��v4򑣮j�n�ɢf�Ĳ�B)���Bn���ܩ1U���wV����²�ao�V�6m��+Sb�;�SU�lK��]=��桷Z3d�E+��y�b�q�x��Y�	�Y@+ʙ]֫(,Ք9.�Yݬ�C[h�F��a-�S$�T�k2�Z�uf�ˁ;2S�e�c�ڈ]�qn�l����w
��r��%�NT�Z�hfD�ͧE�i�@�j钨�@;�k�Ԅ�~�T�T�Vn٨�h�ՠ���;i�%��`ͲhE+pR܃�Zr�L��@�����I9��	#)��]�+c8�-;nD��[h�{FF�C%܍�RDE�In�x��1�y�����ul)A�$6�ǥL��ӥ�=x�]2!��cwohl,��M��W��G,��.XQ����]���ffV�N�L�R���@���6����C�V+[g.�Msyu.�F�K
wD!O e��VՊz�D�)mn@�-e�H|l��b]jc�ӡkq8n�R��*A�̲�q�;��cݼ�j4�&�+X4�!�-���E����F��kuҁ=V2�!���[����Ffc�F�!ڽ�U��cc������˥�0�fܽ�,x#�q$h)I5�RE�곺Ң�y#F]l�Z:Ջs�(6�z��f��DOq��bxE��)Z�-[Xtm�v�GVK-��U�c8);`�9C���oa��N�̔�l[5��^P8�Ӻ �.�Ѧ7i�Y��=z�)E�v�l������i�x΄���FS8r��ܓw)�t�	��!X��f ���8�W�Ǆ�hb��& ��rSJ�Vn�(�-�Ҩ(��Sp�ׄPuqF��f�ܹ�0��0]F�^5�1[w(�ܐ"���%mL�d�z�`"�F��&��O^��hnڔ&�u1NӵM�8Vf֫����!�^�� r��WbSN��x3,m��/)�-����:Be�۸�ڼ��
�MM
TY��>��LMkx���q�˔�\7x鏜�+�_��E�|/��T^S��M8�)Xt����*�]�V+F�CF������÷�ҧ�u�ȕcĥҶ�����F
�
E�݄X8�5�c�eZEK��:�Tj�m��Ƕ�ehkY��ِl���'7m��r�f6��M�f,nP��{���M8��A��Ԇ�ol����/n�50iҫ�d�Õ�0�B��{�t���nF�K�F1�/��M���息>d��os�wjӭ�.<X2n+�ƒ1VܠumTԳfƝl%���h��ދͳ0āD�" 5	6|�a�Mܭ�B��.J�-�4�2n<n�8ĉ]��C#(��Z�ǻ(9"�wP�5k6�͔$l8]+IW�F���E�g�ncʆ�L��ւ�,+`;�Un)�~G1l����tU��B̙[��4բ�f%v��;�wP��m�1�" `P&F7#�v�#�e�n���#���̴��E1B��G�	Ot(�����'rԉ\kd��k�z�;�bY�(,fCX-�-�ĔZ*Q�]kP|�Q-���
��#kn�u���fl���j��j�e)�饶�|36�J%�5H����;*6mZ&�0�;�Y����.�-0p୛��;6u�$z-�C.�S�˲Bt&��(���,�ae�Tkn�����\�5��z~G���U�����b������TlV\Rԛ��":��M��A�m�� (g*��5��3S;_��,�03���Ҽ�Zw�p�q ��4F6��J�j�'�Dʹqi�����fh�f��!��� ���̭d���Y�xh�X6�к�R��l��Z��M��(MA�U�k,}};8�g�͵�O�
܇)^���`���ZY[zC��j�&��"�]��4<5��¶'�F���R�m곩-u����=��@6K�k�m�E���Ci�em;w��®����(��¤E:��7Lwh]�U���V�T�ДZ!�C�Y�Y Lҳv�bN�T`�eK b&�Gov�n���n�t�bX��צ#� 4��VY��*�@rLP-׵���� �Y���N���t�P�s,�q����[ٷe7{���mjQa��. U��!|�eU���*�Z�!8�He'ys$�B�9ݑ�*X'kT8iQ��S2���q����3i��#����s0���
jv�ڤܺ��[{	Y�`��������j��(�bH݃��m�o+����0/]�m���z�+,j0���b��Y&ef�Ȥ˽�u�;C�H���qE�T�VXC%CNAz-Ѧ��9cWNcAo�[|���ft�%]W�z@p[n��5Ņ-�o#[z������t ةV�[&{g!����'/��(�v���E\��H�82/��s�Q����m��D�HR*,�S]@����m��l,	ѽKu��J�aH�u�QV��V���u���l+�N��ERa�������SZn��n����Y
e�i�uh=j�.f �U�î\շv��BU��������	�*�-cdj�R;V��Z�S :2�d�EZya�E�fh�F�r���.�Z��W�#�N�A���5R4�8��EKQE+�X5Z�M���*��=�ZKa���fd۹)K�H�(g�c�bcxs:R1�N�.�aڄ9O`d5x5eb�ע��U+*Q��H=�"�]�-��k0�����7�@ڵ�R�	�Z��ׁ�KsuU����L��T�!Tee��A�0�n��a2diT�4qH��Z�)�+l��9�Zߦ�
m$�j�m�#��T�p�e�ºl]��M�sSS&��Yv��E�v��K1��(^�FV]�p�%հʐ���NnI�#��ZV�;���a��m�IYk1Òd/lc�$��Q��TC�_]�6��T&�nѮ8-���x셀K�2�cy����B�-�c�r���B�4��k.���F�5�uH�M��������d��Gk�KqB�������2���u(�u�����y2^���V]-;X�Q1��A*J��j���u��,v90���B�R���v�+)�
���f֙g^J�16Y�6f�ؽ1C*�b��ɤ����DȖ��o "�J�dCn�����K%���St
�]w��SqQF��wݷi�VN^U�� V�R8�����t,��Xp
�s�2�(�6 !��鋪�~0��X+*�[��a�4�;2�ʀE�NZG�w�,VLd�9V{7^�;IB:г����!_ua>_nb�T�*.a,Ej�cG���l�
�8%`
��ဤ����ݲ�YNXϜB�LU���Jř�Q!DhȂ��YW@�V�fZ�ּv��Z�W����A/
��tx��
����6�s/m�ȃ�h����Ҹ�̤	y���/5ɭ��v����ɴ���=�u��#0@]ĭV��Β�v�72��L�F�K�v�J��r�;-ū;X�����]���;.
��15�kr�%���n�bie�B�3�9OQ?+��32[¯ �"[���b�2�7��[��dݽDdz�[���N@<�(-c;��dU軚i�uc��F��@�t�
�S������1�hs%��M�
��PI[��w��ڷ�t`
�u&�9u#:��RA�Q�q��R%F|����2��Iɷ3V�L��Oz���[˙�w��Ń6\�*�ޚ�W���	i-*��I t��b,�P;b�p���6��CyD)N��X1V)��Mj+F�]#�k;y�\��X�ڦ�Zܭ{2�`@M��逨OC�LQ͆��ܣO�J�شl�Z bÂ��	�(6�����WrJس!�5��@�. ���R����D�DF2��9(�_5`�Sl���8�X��1@�V�mh�����=��G"���q���Jv�6�D0�Q+���[Y�����¢ɲf�Û`:��(�@��U����� ɵ,ة@Mn��ʺ��W�g�Gu�B�f;�[�57: �/H��1T�6��!j����qF^Z�A�F�b��f�-�(a�AF�Lv�m�������V��~��GX�]�R����r�He\J�bճPM%7f,����Hd+ ��̢��[j���#I��)\ۣS�p�J�Q:�7m��	&�f�d�R��[y	"19��M[GTf�ha�v�6�+�[t�	�U����Ɏ3/x��-дb����SU��ұHh�7��+�ƻ`�-Rf�"t}��!��Z�h���ƃ�޵h�� 1�[������}<�-���Ք�%�AJ�`�]�L2���!����G��$14+�/R7��[6�R���V��֔����(*c+AEm;���^d#-�Zo-P�YY"Ӧ�vXY�q^T���S �\{E��&��ʥ�������.����X����4,�`R�n-Rl�u���B���JB�D�`4D����aj�h#{��Q�xt�U�c�;Y7�@���[u��4�*HA�`��Df�o2��ݹI����|o���Q�����04'�bݶ�75�*��ݵxΚti�48�"���q ��v��m�5+&Sgj6n�5 ��B�!��]�Q:�XF��IY�ON�4�a�N����L2n��N�Jbl���5�#a:��1�MMb�_m�@F^�P�VwP���ѣ��4
�
XN�ˠ�h�gv7wk�i�]�V���$h�RU�6G5ZH問�l�*��l�V�4
��ݲܢh��K4��v ��!Zu�m�+TM�j��H�ݧS+V��Z^K���AK96����RB�Ȕ��tն��ֵ̈@7��l�p�a)J�>���b��nƻmicc2e�W[yuok1*5�/��K@�7����9�RdS��ܽn#��X��,%�E2�SiaF0Mo�x�қ3�/lA��-�kt�p�*'J�n�ufǮYB��̡���Dm��\d�@^�F�jQ�pZ:2��L��l�i�or��d� �p`���%m�],T���x���{4hw�
ۏbz��v����b˳uL��%��U�n�G��r�QP6�)'����F�����z(���=V��Z6
d�bҘH�r��ս� r��A��ӎV�7C� ��lf�}�ƙI�&%#3%#Q}�^7��B����%�u��z����5<66���oV Z�Y��S���*#�Xͧ�K�K*��!P��� �Lb��Y"�m2�{��`��V)�%^�ra����Qr\��rQ
�J0�qL��ؔʓ�̓6��˨������Q1x�m�m�����.�{��tV:�V��l�����kmSK2�+e��	�P���JP�J��q������hf�Ѐ7�pAd�y3^+�ə�8��0)�)�ʆ�	/>��`�je0��7MB���
����o[�vZ�R�BK�u�w!X$5��jn'�!sdVb�eXj�H��iŐc��ͭCi��D�M�i˵wv�ї��;�)X�2�ѻ$�&�D&�W�"�Rl��T�����c0,I0�f��%ݻ�HD��r�����ˡ�#���p�/�x6�f�Dc$DZw��	r�2f�WXjM�B�ҋɂi�.e2��2�(Z.e���x�G����dߞS�f��ێ�=��[$I\�k�z�G(=���2Rw`�f8C��ų1�Bӣ��lk'Y1��XCan����7W�,A�擙��U((�bN����Y�KkT�.
��Z��+6+E�m7R�y��S"�������4x^��Mm�8X��MT��.1�%Y�f��8�K)ەyp�P�*�÷^dq���8�U�P�K�cF&1��V�KF��Of�����zMMYX��_LA][��PtV��J���2�̰.��̂�:u�����WQǡK�X��N�E�;�mT���l6�V��-4��S8.^�1�� �P&���Բ*��D��N^��ߠõ�XQڒ^dv�ۘ3dpl.��mZ�ڽ����W�Ru�$Rޚ;��SEգ�PH�h!!���%��1K��$l>�H4�H2f]+�Q7��Z�T"�����@j*8��
nnƥ �P0i<�&��AA�kq�l��\KU�1j�e�A9�+��K��a�U�(����M���֬*����%�=	l:�c�sMGb�JѨ�ަ)5*h��R�C,+4iB��f���S�N�!��O��Q6�ռ;x4JǤt�8��ޑ>�sObݸ��9��U�J��A���oz#�=�K��	�� T�m�:�gj�wV�\Q;��}rB�Е��xо�
3��Lf��r��B6�����l�L�}�v�֭�EL���!�ˑ�o6B��Y�����yNQ�Gq��_��]�Sl�=��	R�T�v�ޕR��_4/^t=q�N�����۶w���L8���=���e4���c0`���q�-�}��pXir���e����&i��|�j��TVV�X�D����U���T/l��r��1CW�|^�R�o�+2�������m	�W�����j���n���(s���VPfj�i����xE��N8��vb�n-�nfǒ�pU��u��{;0�t��A�J �V%D�Q\&� ��ս��j�v��`F,Rq72�����屸�!	Zk��X�5�T��Ԃ�Ċj�ld�������2�L�x.��'�\	\�]L��q��G�	�I�:n�u���w0s���;=�D��5����Dշ�k��7G��z�tY��<�g�����X9�� TK^��B�T�L�%�R�%lf���N���:�󻰀c�H*:)\��T�|M�`�t�l\۳�F&v�����t�>ۯw�%�����7�N�%��a��.��i7ѕ*�z�f�}f�����-Z)����ګ�`S�,;h�=2��%ؖ؄��s�C�8ڙ�e�3QE����T���ZζP7hR��e����tL�,�(B�A�>H�E�BdjJm=D�R��On#la��:�uݷԔ�N��c�6{��lC��ʻ˖�P;Y�������ofm���\�T�[:v�V;�������o!x�Pטѝ	/P�e����6��4�;%ث��v{���T�Wm�W�JnlO�r�#x��5,�NK��Vֱ&P�SJ=���4��}�)�3�t��V_S� ���{�iN���Q���Ws��죳"J�;V��T�}���3�Ek�5C�;5�ظ�r�	�ѫ;';�N��0�쿡ʂ=��>m�7�>���u��;u�j{��1r�ڏ:J��*�Lv�l��ά���R�s�p�l�ჇC\J�i��>��M��F�8��VꈘԲo-1�$��
�2��k���U��/P9����k
��n��4��7]p��{��cы+)�j���8إ�)v��-Ea�*��7z��gN���I�U��֯��5z�v]�ֆq�;�W��1�(��VGm�mM��+N����Ʉ�{ȉ��@X��Lj�q�;��GΤ��2ͤz�F�Z���~�O
]ۼ��\S��k���Xy�#�}���B�P���t���wt�Y@�;��.����)�}����β�*�=`���VEr�m����*�m�>9p��]1u]�&����-�}q_rw� ��qY��/��3^]^�]Mٚf������m��mfI�u�B��û�ݤ��yNs����^i�ѽX]0�=T��=��"{<���j�9����Y]]�d>���
Υs�i��f��Y���8����2��԰�M��^Lg�c�k���y6��J�%��fv|��l�=]EN����\zn^�{�L<����ѫ\0WGm��)N��m��j�J�x�k�O*�g8x�:΍<å�ë��>W�D�ŀٷ2��Xh��=��
;��#�;֮)�
�]m_j�L��f�R�b�3��n��72I��^����ά�*-��W�j�2���6�ם�/��
{}�K�f�B����������javst�v�ވ�Ǆ�{F��L6:.Y�Q�D��ƻ��S'r�6���Syr���_i�;Qe��/��J�8���â����qa�EX̺]����<"ZL�������NԂ)�1��P��wf1a/>[%m3j}3j=c�ĖNwH���}�1���h��tEE����Z��q�+bX;,qt�|�j�:j��Mn�T}���p�7x�ڳ,-�3eVrkUrҮ��� ����07�C��o��4�"�-hfZ*6��loW�iy�&0��割��e��,�Pp��l/�c�'u@W9�T��f	x�
Ow:�]����Vn������%Y��Q$.�Vn_F�WM7}��jY@�Q1��]N/d�����J�Խ�ݳ������T�!�k#�g6#˟m�e&>R �L<��i�W]Q�
��{cn����I�:LfaW�%���U���c����$me�⩇�8E�ۧ>"�u_X�ut(���d+�m��\������T۱�r��&�tC��$Q�/*���oq�� ��i����;E
Zԡ0�Y/K���KMu�Ɔ
:2�� �]u>�a�+]q�wO������%���q��}�O˩X�Pq �}�D���3EG(�dő�>H\��֖n��[�	�y�'r'7$%l}��:C4ڭa�7м���x�e��q��8^-6���ݱ��Cț����y�ǃ��ԅB�^�0-y+U�ej�lT��5�2�4:Ε�\���(K��i�];�`��q��u���N�[�0�.���hDͷ6N5m)A��rn�#Ήlᷛ�G�m�|l�J�%wSw���I\�.���Kz_G:l��XO<��2�C�
���Cf4�^�m�[�D���]��ݬ�0))�
�eC�9��λ�ϯ��Rv13y]�՝#�opҙi��<�yk��e5FGҝk�G�a�s�"s��@���!�3ij��l���`[wk�4#��z��;v�����ܥ���æ���ZҔz���LB�aƮ��Үۢnnor��f8��Ԣ�\͗ �ma\4��[ْ\�e'{�c
�+�[�����R��Ԇ�̻5����aˇ��������^phg �a٠{y�1}���P:y���.ش�y�+�k�a��˚�M�ʙim/a��EkŜYY�c��O."A4�<����ҝs�[d�8��,�R�Vom����.�8o��Y)��FnJ��S���3�t�v7���]�ڛ]Aj�n��Ws�v�]1]	�5�S�uG�ؚ3�����NMn�vg5�&1Xi���Ҁ�����	m�����m��P��ˊM��WDd�p��b�ɗ;*1MԒ��3±P�U�t!��o�Ү �g�7�	,����E�a� ݣ�8��=�D����3�Z�-pνJ�HТs/-:���.��L� �[�uո�hݩR�X��G55h�| � �E�U��٩�F�U�4������ �ڝb]���s�Y��s�P(w��P��	���ݫz�U{}a��]�-�6k];|_��4�d������tk�\���c�:��iB,�]s��D]]Χ3M�ke������lO�R��6Z9ٔvݿ�q��l��a]kO8v8:��Z�D�x��B��Y®�(���+(K��q��i�H��j�b��l��ܺ��1�GRb5F�8\��޼�̹+�l���B<�]�J�V�L�1ܘ7�aˁrd*u�r\�nі�V�v����7u��S�>�د���9]9��,J�DǷ��/7{s��V�Cn��d1T|��7��W�lF��ۡJ3�Q��*� R��ǳU��Ƴ�z��޾��o����*�E�aD�O5�[oB�K�kO7R �>���s� �ec��owe-g�!z�}N����"��w�m�U2�3��^хcu�L鸦��.���S�F��Q��564]%(TkqjwHJd��ƍ�N����L�u�Q��]c��u�e��0�;��H���������(F苾�7�	y��\��<0���+NPt�b	A	ܷ�8����1�F�ky��9�WsK�=e�[V+B�/,�Ô�n1�m�v�p��V+�)�p�s�Es�t��q�U��4�;LٻW������BF����hu��S��;54o_v��¯s��PN�9���,\4���6au��:�m����opf��N�ΫK�9s0��s,��<ڸ��UljVrږt*𷳞���:�����V��"U�⃋�����P�6S��LW���^�{~R!�5I�T��M낙ۙ�ޅ͋�v6�̝}/bY� ��L����������`��΢�d�F7x_9H�ŭ.hEf{,T-3\����j��er�D�r�K�ֳ�"]R��B8�\�lc[;�C)��Xn,ô�����Ra8�r�l�%H��2�zz@����EeJa3�r����\J�1�L���C.��4��]�4!�AXC{�[m�R[�'k�<{Y}�������n���1�|6����O���c̴� ͝�H�Wl�r�T�yf�� vDo�P����d[�]���m�ғa�-:&��V����L1��,v_]P���+�$�wK�*+�cc�f��;���p�o]��xK��T��N��1���`�����=��7��:rx�(��;n���33]m��;��봳#�D9Ja�dƮ�dgVR�l�q� b�2�ՙl�#FQ�mN�+[�,�%���43�kO痮\�<��<zvfK>W��.y(�A6w�& ���oR�j�<kL�T9R]�f+�ǻ]�s����\�	���i�*�+�4P�K�����.'�q�ren�o	�X�wX�������A�N�t�:$�;*C3�M�WK��]�erW�� /�Ws��^:��}oM�����ͬcy�ܫ�<���(ՠ�0��
m�.��Z��o:M������İ^ՌI��U��K��V9E_�̇�Vm�Ǒfت#;�T�������7�r�>W�f� ���t��V�O+��y��!7��[�82AQWP�{&R��T }Jd�Zpa�z��e�C�֮wD��k�N���.xr�z����P흍:3+2ļ�蓱��<�̈́*�l]WUλn�ծ�5��X���,Cx�L�W3]�N�}+��f��8j]�.��z�;��ko�Z&���]��+V�3����%1B2�Du
[�~��89��k��ųr�2ދ�D��W$0J�oVuS�[�*�;�o#�΢��;��o��t=�k�
�'ޣ�)8��1{7����p����m�s� o���r����I�f�� ̶El��wV�N�\~nVu��+���ݓ�\���l���0�<��.S'V���=�dƣ[Sn��V�j����H����k�*��l��}¥�\�Ӿ��F���.��d���Cka�0r�K�uy����q�/iob�4ej������= ���͠�g^n�\ V�/��\�uu
N=��+!�fmtϫFe���K,��5� �Q��d�p�N��Ȥ��Э�+���5�N
��K$^�s��ꮰ�(��ĥ����F�_M��bHq�����wm��]��G��uo�i�H�Wl��|;�����4b��ad�;[�gp��ڍ�\V�T�[��6��esg�r�c��%�n��T�p,U�]ը�cWj(J�Y��_ͷ)���Z�G��ݛP̷.�`�ou�<�R�����sVur�NQ�P�s�qY�]Y�3�v���50˕��Rg�J7��\��L�we����왜.���1p�uۥ�����QN�ДVr��4��a���h�Li̍^�L���+��oa���)q��^��±�+@�E4A��Ǚ̔��a��֊�ʀP`�˵s�8��/�!�k��eXu�J[�X�Xn�=��Q.�����Gtu���@yҮ������.�k��7E쒹x��8�X*��>�2��`�z�U��,<)u���.:qRj7]��7�0�si�{�-�O�ޅE�;��salZ�>�|$�Vm��[w��VmF�[W��l��J������ϳ+�O���8�ޗ���ď�q�:`��[�GZ�=���ֺ�b����G��u���/�.;��8(����";ӡY�Δ@��+.�:�4)]ɘ�`aiӫT�kM�	GjuYC	�h*MNB���δ��\���9v�]x:�� �A���r����E�]Y|ټ���ݳE� {��@�f��V��1�A@�v���5s#W8�4O[�s�k����[�#f���q ;6�Y�d2�J}�a�oj�5���\�vH��� k�PV��LEC�+��W���n�<��
̨=t�<kh�0�\*V]��w��t�����.Z���K���Z�k�j�=q���
�(M�wk�:����#��Iյ��$��@vC�^��r��i�pJ�CO5�s�h���yGmTu܁�(^`�ȟH�W�n����r�lc7�F�
���ܘ�!N��7�K�j�-�:R̮�7��1S��w�Vk��iff!t;o�7d���t�n���- ��p3 �R�؍�˞LR���ךR�Y��{��Ϸ)Śi� a�b=�]��3�(�[�EW���SY�"���}y�b��n�l
0��^�;�Qv۶B�cɭS��4��nh�1۸��oM����uݔ$�Z�_.��w���OIkv���S\P4F���k5�pB�b�WZ�*�%�q���J�N�3�'�wGq=OUeg�*��kQ kqbF]6��#1l�F:U��X��ۖ�:dw`h��\"���H�6'c8P�%M�_h�缥�*�X�d
f[�|j���Oh*��u���hw-ӎ�Y6�Xt��bS��5��]����>���G���m?{p�4v������{o+^�S�)��Һ��-��u=[p�v4!)B:�L��0�Q�R��JX�r�K�]���%iwj��)3ۖ���an�Z��х��
)��?���ꪐ��@�$��}���۞w���{�w�	EO����[���N�uI����~wFa��;A�QJ�`d�
�{�!��oP��A�P2c�s�J�Ds 5k4�)�|�5ǃ9��eԷ��
G�����
�P�욺�ͧF���às5ft1I,v]C%�hk��\�R��-nU���]��͑f�g���:�����*�(Kث;����q�q�xfyP��}�燪���ɻ��\����[]8�Z�B�V
��T�p��c�o[�O���ċ��;x�Ҷ���*w,��e:�3J��I:��@�iFQ���8��o���F�Ut@��كWs�[Nj�9���3���&Ӥ�2�J��R�w�h�M*�q��t+�r���P�F�*��ݩ�t�oZ���L����w�fV�t���$l�]zh��6�e� n�Z/�7M��K�ՁB��2��4�u!���v�2��ko��Ѻ��<�ĉ2R|!�ٚ�/*J���]�v�mX��Y�e��U�ɡ�����Ƈ*���'`�*K���]�h�z�8�2*�;��,�b���/^"�U�(�{�`n��Ӽ�Y�C�;�x�S[qˁ�u.=�{�-ѽ	M�uW�0�l�˷��ټ�@�j�9w�]��6J���,�)���XVB��82���栴l��1�pӉ���|�H�6d�̾8v�`�й'����v�
ްNϴ���lhcC�]S�S�(��p]�G��JU0���\�\�g�}��x�*���|����w_7X��zF�6��^u�&J7�1,��Շ�ƿ��e��i�f�L%dૅ��^>[��=ע@�� �v�
��YkkH���{����wmtU/��T��(� ����^���7OJ�e�ah�AB�^�,����c�MF�jK	T-!�s���մ��OLow/cʛ��*��(�۸=�RZ�j���Fz��q��Zk���j��#��wݶC�%-�����	٘���t��)]ǣp�T�'֖c�ѣ{繭�5e�_u�e<��`((o-�t#���:ke��\�߄��m�B�����<���دj��h�A��E������F�Afݽ�F&t*w+�J[��Xj}� #�y��v���IϾ���C��猥k�5���Fbc����y��փ�,j�mMJ��,j��1^c-���'Sx'oVG]*Cz5X��6e�xe���V��c�N��]���f����nr����|8�L���51�+����n����42V� R�2dWGKH�j�:�Y]9N��m� �=��yK��OA}Y�����\;F�̸��=�)m�ݳZm�m�@����򺁸�J��ﹽ\���Y�c˻8��1��?mhA��sef� O]n�Υ�Uy�&��U`rܵ�Z[iQ�.�p���g���ဧ&�W;Ӆl�O��xB8>k�<u:]��"Y��J�u������JF�0�\�#P���WE�fV��)��|�n��i�]����e��w�Q�
����S�)bc&p��>�^K��뢫v�a�\mGt�����p]��� W�QC��c�6�CU[�w,��	P��̄4/�h���A_
��Fk����ѣ����YV�L�nl1�V�(��ɌN�7��fd��{��|iA �tU��.N�V�5;4|N��85�c��Gi^))���-Mj�ٔ7�RMg����k�Yy��-uh�u����)����ž�Pf�O��
�Gc��v�7A��!��iCݵ���S����c���V��5�%��s
6�1���H�@��W	���#4o*u��-d��k,�g	��7��r�(2� �	���f>������m���������O4
���� �z���Yk�>�4��@�؂�=�J [���6��C�p_E�	�%˾��Ǔ�R͎�I\�v��C�9�NR��.U�����U��ʍj�I=Ĳ�j��Յ{���v��`�A���g`���5�<��v.J[���j�:�sK��k�^Ʃ�@R��tK8� ސ��.\�,���y��w�RYKCu�$�X>_l;� YV�'�u�݇Y�]j���ZV������gm�=�r�o���2V�7yҭ�D��C�E#�o l��X�S: +�qGښ���q�֗;e`�ʠ.�M�i��&��RM���^�j>Ƀ�[�]ی���U%*7Y����JU�'�	L�f�j�CA�d�G�.��\���b�z�s�jh�VfY��n�f�N]�8R�7�-�6!:/�R�^t�J��S����^lZ8����ݮg&�zz�d�z�-�}�[��λ�X:��*=�s��K����%�c�qR!��A���x��ïdޗf>�(�,���S�#�s���&V�,��I�ע��e*T���s�YU�2�N����'6Q
��գ�U��A��2�ʻVo�-�p���w)�&m\+U
�&��K�h:;j2�m����#�R��Tz������f�2���Ӑ���#���M��ڸQ$�qa���a�@��Uu"Ǖ��.T�K�Mm�}�����Y ]�o+��[�N)�R��ev�Y�'XϩpZ�_7&"VVf�>��t�6x�*T�d��B�eT��7���J���j�lbB��L��>�ѵ+��Fp]Ғ.Q���ŕcbb��(=�q�&�w=;�;�3m���yÆ�E�W�5a�a��$�X�],e�4yh���:���B�����vo+�hfR�ҹ`��ԧ�*��+��ĵ�v7hQ�)��I;95�I��]�J�g3��v���)5
+��e���P˫H�+�QR����͊����r�	�@�G���N�ɉˎ� ��fl�i��S���l5���8��-��s'FҸ*Ӑ��Ƶ������RJ�#n�u[��pd7�qK��V��o���3d�R�Mg*�XF�rr@�����Zt(u�O��~���F���)��A�agl�Cwa�Il>�k��ml�P�E�@�D����4�5��;��m輰s^��β ���;�d�{ۉ�6��H�o��U۠ʱ��wWM�4\}X�*.tq9��r��o���ŏ��a`���\�dWX9=S��Z��Sݓ���;9�2��,:L�(CԱ<�f^���f�4�t�B��:���x.��Ny�H��>knc�7�sc{7�<�_]0�9�]e��V�aq�(
�W�)f�`D\ʻDfJ�d��/�0�������ۮ�zcv$�V�W �V��/��l���,r���`֘vF��ܬ�I�E�v�56� �U�e&F�D@�ָ�j����d�v��w���$��Nd�yt���BĈ�y����=���	�ݨ3 �S���/�Ҳ��|��C��0
�\C�˸�t�\OD�x����sm��T��[v�5�7Y��H�-�;������uG���d�gx.lì��u�b�NJ7�%��)�`�Ηf��I�������&��r�����M��pVn��n.�̨wUO�r��8%zj�J�]LKi[##�͙�,���u�ò��:N`��#%�-��c[�|�MJ�����o��On����s�%56ŹY�mV�9�m=����^j{)��yi"�K��+;-�����b8U�&_�9@Ɏ��w����]]�A�Eu.��� �S��틕y��#"��6���<�
B�-Eɾ�8;.��{u;��I1gl�+����R�y��:b�[�u��� �	,�o2�W[U%4�w#��Y7�1|��M;��F16�bʊ�l�f����@7,�pպ.)B�ݎt�8��n*�+���)KWJ�M�,�O�Q�"saV_g]2�Jk��TT:�䄬�n�e���SIO�J�:;in��j�--����NU��5�t�m[�g3�+�˘���j@� ��ճ����2�t��U��뚙����U�y΍5�vVVS�y5V�O1d#j2 ����Z���p�#�H]�/!t����<c@��cE�3u�mU���Zc(ѽK١M�*D2i�#V�b	��t£|yvu��J���ԣ���yW��>�ʔ�bg-���J����u��Aκ�iv�I4E�m=B}""3��%�l�Z
P�-`Ꞟk�&��m`�ښ(��4
��A4�ҋ7z���u� �5D�9�tq�mG��s���>���`�t��-}�m�4��pf���5Q�21Yg��܉ѹGTQ�mРN�r��6���;��an�FNrjQ5B�̽�̟rG��_&0	Av�ꣃA�Q}�����C;v��4�_Swq���cZ'�x7v��+3Q��VՍ�C+z�Š��q5��P`�(:}+���Z)A�ڂ����
"LV��g,<�%�����$��j�[H�/��k��:�&���(�n �6wh��P�M���ܺ�ۮUô��b���u2�!�*;
�e#*�_f#aY���o�s�E�C\��@W:�� �)�В��%�l�g�L� 5����_b2���.Nm1�]u�g�
Ao�RS����hu�s�ߠ]�e۱�$�X���C: :aI��q��䇡��մG�
=;�Z��wu��B4-ӏ&�9�Q�9[R<ډWFd��XT�{��+��On<=��fխI%��i�l�6�}8��e)�X���n�h�}���͹�@=�p��XmPCP��TvGX͎�ke��^�	�!]��*�k/�B�ɔ��S����Au@�ő������i+.]=����e7o.K�}�}�#ݖ�t�*��s�+k'1��	����nGۄ^a8����s�bl��o���c0��c8,Ie�I(w���g$xo���b�$�O�6�8F5�nD��=%� ��,[��nj�z�FT�"��(ֲi��̾��fO������k�q[����]JV^�;�6���j1�������W���o�z�7�m��['2��<Jɧ[t�+��0�;u&G"�kY�-���>�����Z�Z����幈�U��'FW���{��g��\c�%���3��j�l��َAx*؛k2��3��1�u��;�-a���W�G`w���o�����ʶ�wR�Ԋ^��2�'57j��{��̭��Er�ם:�D�n��uА�Ri��"w�YjH���j�/FM���N`�уe�l��k+*-.��UǥfeM���,!G(4B�7�O~�v�cu����D0��l��ݨ�f�p>���NS#B���N�p����5בP��Z++�Za�ƘZ*�*�f��7M��C#�@�E����1ps���?+�7VDFښ�Y�57]]wMRe�42�풢��Q�o�"���1s;�
M!�9��}R�AH��<��v���������`VO�˲�g_'�/���&�^��P�b�0��ɂC ۙ�A������׽�l�:O�K yL�Ǯ���w����L���w4����O�W�΂�.��ᖴs[�y�p��v�+etn����T�{}�v/�"�K�J�O���|XhwA�0ֹ�x�>�[�5j��.�De�k��Ԧʾ�ػ7�G�qL�֥!:�T����|��g!u+������@�6��4�v�.Vr����]\�v�>q
��s�	\����;�wA�+����U֔.��	+S��]"�#�.U���6:���)f�2Ŏu�e��e*�v���$G5��h�b����}+n�$�h|8k��d�Qӛfl��<���6Ҭ9*눂�����-������-�Z���:�s&1K��4h,��e�e1��k���&s��G�>��6��Q]>��Jc��u���$	 �����=2�JXdۏn��tJ\W�V��5L$��w��%����ŀ�=����TX����h��RU�ʊ��^�f���
}��0\F�XF�*|�싅%�Y6���ll6�Ċ�\���S�k6��t���T G��iv�Sҝl�i��cgMX*�4۾=5;�n�I"�)�V�)ֻ���*����6��f�<�v��w��;�z�����֊+W�7���*���ǥ��o���ʈ�m�(�'uy�t��W�}�.��J�*PΔz����J��F�"��V�����-��Ņnh׹�[����,Ҕk;�h�.X�Fl��p�^S�̏��g�i�dD��Ψ+:oD��+-Tg��|����w�E�В�ہr�+J��>{�`Ӡ��yU�{Kf���۶��i:�[�=��%�o�f+E���$q\+��)��rj�K��j����\�����Z�sN��;o�pb�q䭥��v��Kܜ�k�0�&!��p�jP��*�jD�f  _1�}Bgvb�m5C�]��a<rp8����k�&l�1�@��M�����������
mŎ����+��+��s�:�_305�[�Y/7.}-���ۄ�Z�:�|���ƻ{/ ��$����0/��/��#x�l�:xV�hmK&�e��bN
7�W`�L#����*�1��YG0iXc�G�A�,Ш5AX�kݠ��/�ٮ��m��+��;�C� y�f��o<4L�!X�q�
op ������=/%*�5��%��Q��k�ТGj�������s�E�Qi���
�fN_-LV��Z�/0���4�D�<1)J�'.M�Tw/0Lt��qrWK���j�\�]v���yLF��ܴn�Np&]Z&���)GL��)ˮܲ'V����Rcڱ��� �0Q���mǁ;�I�AJ�;�}U�����<\Z���i��!ѳ�qeDK:��NA>�5kqS5_�7�Q��k{��v-sO,eb2
�u2�;�^i&��+<%i�OyVn�T�Q6�pL��v����d��IE�gw4��ȴK��.ʲ~�W 8�t{�`�0��w4^�X����;d)逯p�j6ʡB�
������ꝎW9���Mu-�
��ٓ@X���6�.\�;ξJ2:��s��6$�z#��i�U����[�u���ՙ���r�`t��P�K+;X�}vu���6���&Ȣ�YR���)Qt�L�j�-Rݑvf�q5�囩�.^(�U<�T��w.5�K Q
�t,9%ܡu�T��X�pL�-��Z>��NQ�m�(���u˳i�#�5��⬊]���*mJ��W���ɮP�����oqu��q�]mO�>s8n��{{'�Vۊ�\�Í���^�69�,�wx�'��yN�]g�j.�s�Wu��KoC�!�]�*%S�u�����l�$|�v�+tE�J�j����ڸ�1���+n] �U�JdMޓ��� !��ut�����:��jY��#:zɶ(�������{�q��sql,�o-_�-�IG���$��ܰ6k�r��.L���/5��'��
��ڈ����y�/����H�?�}�7oiή���[����>�*���b��E����*�ʬm��EU�
��%kPi�D��`Udb5�ődj�""LJőB�(őJʎRU�T���E+	[h�e��m���R,"�V�ʬ�Z���D*E�ʒ,��
 �"Ŋ(�,RҹJ
,�h��+b����%j�Ơ,UXDQ��D����A
�X���UA��P��"��DTUR*���Y"�(V"(֢"KB�,�P1��DE�Z�E�AUXT*��Ģ,E�XŴ���A�(,��,��Q`��"�R"#m�TR,EaA`,b������H�DH�AH��2V`��1��
�QTU[ZFڂ�PZ�(QU�QamU��
�`��F��b(1��PP1�PU��F
�&YDUb�UQEdQA`(�P��@��%Q���[D��庶�tOxZξG5�ɝ�
��w`auZwZZm���[�QS�W,�ۙ�(
<Z��p��r�s������T��g$������R�N�]��{����,�}.sp8�P���e��Zo��k��햫c�p�m,ҹ�SՋ7/j{1:�+DV�itf��XEs�PG�䤍j�#k߆���G4�j��\D��UW*�Ƨ�)NkΨ���7�$� �G-#q?�y��>��q�xYV�������)��ԈhS�g�I��7>3ظs��:��wr�FڵR�XY֦�;w�q/��2��١�L��M���U���sx��NϦ��Gƫ
ͪK�aj��X�ٗ�2k�m>Ra^,m�����j!��K��K���.e�����x����t�Чq���,�Oy=����Zf�T$`nNe+��n�^r���jy��+m����Z�:�wS�Y��צh]A��W�qұ91^�E�U�q�L���nZ����;m_��P�Qt��;�3�$���w������qB�T�C�/BJд;�n�*2M�)[f�SoU�g��O#�\���;,jfL]IZ�o�Z}�7�����Թփ��F��ߴ��ٷ/��`� Ś6I]Q�_%e_d�� �c�������N�-����Շ{6$;��T��۞����"�M�VU��(��W���-�M[�:N�����̓�YB�z���\�_+%����~��+SU�.kة����z�*M4ʷ�3�v��u����ab�QP���݂P��{mM��<5�W�WV>��-���"i�k����*�`�:]�e�Q{|�e��T�pG�� X�3ױ��,�˶�.��+ˇy��U3���P�ܖL�L�3qy�Ew��ک��/u'��k�4�w��*�����:H{���������z��WW�|����s`�N�
�%\pRȳ�]��;�K��R�!V�ޝN���ָ:�MU Z�á9I�mi��fg�UT`{��o�=�eb�֣={j�pt����䦅��G`�g'���5u���.NV�"�"�`���н����yj�����|�v�]����r
�чN����M��_O[ވ�8�v�-��=��X�VkUd��Ty�^��;��I��+?>�ä��Q¨a�{��ٯ�V�8`j�]:�ʿ}�ŢY�����@�nhfu��j��s��x����]U3��5�e�!�O�{T���R����4����n�4,�wa�gGTge9��+��Ͳ�v��3@uA���l7'2��N>���J����9�S�y�M�s��a���V����YOk��0<�R���.����$����éRԎ�scoS�:v<����u�S����%x��=.1�����ѧq�7/�Ѩ%~�-����:�f�j�-p��uur둠�Za���L%Gd���E��J��[{��b�uejɉ�������t��gc=��tHܿ���.��jh_Ro�Ml��L��;���vlhmq�L=��;�V��p�Ѓ�)(Ubo:�YXrq&�C���e��St���֣�Y���2�����95���;#�-Ӭ�`�=|�*�h��9��}�k3-�$�4����ܚ�	V�������D����ᱛ�g���[������q7r�VB�#�W[���K��H�u��9���:������9�ќME#���x�I:����Y�i;[mU�}�o����]��ג�%1d���d�7�.f���)c7�鞐Z�����|�SJ����͑N��]�2/������a��� �H��X���v��j�k)��zt���_��W�c�KN���\����_��"�<^�`$9�@��)���N�{�x�?CB��v"u�����/�7����US�Ⱥ����,5UWɳ��_����b�FBhc�sf��U�䶯�QS�w7 ��i��ӻ#n����=��r�i�|����<�ʶ������M�jpQ��>�&{��~�j�����{y����a�f!I�{=u��2������/f�.���W�Ib�ֲ^NL�M�� ��k��M�f\���d��F�I�4��;ݍ=C4ۮ&����V�����}]����!����M+�����4�U����Mm�h��n�>Pi�����2cш��8�@�'q��L�'+��μgE/�����\��]m�Y�T��ݲ��!�6,���M���3��F��6�v�Qf��)\t��bq���9^�|/T�}��v�:E���d��'g�Ȉ��u^���i�g��G	
&Il�OP]�T:����Y7W�
�z�@�5lq�\�9��T�d����g$���u�3��Iu������� 百z�V�x̭Sl��"�W�b���aB�T���FA@�#"�(Έ�=i�(��s��z2H�T�*&7�֯��)�^ %C]�GX�BѲ��W'\��r�֯j�"9.9<�}d]h�����so�W_ř�p���űVq���a�h�y@���cD+�)�;���E�Eo�ioǅ/�)X���EF��QcT���
�v*�QA�i�ɔ��k^-ң[��+�"����Q#�R&#���#L�s�+�p)�c{/.k�{;�`�-������;<�h� (F���Cq��v����4��o�M��㝵�up�AQZӿU�.,8	�SQ4�F�eŇ��zI}
�"��ʬ
{����L3#1;~Z�#�k��94_g���A9b6�q6f��Κ���ي���o"�Hw�������~�t8�˫	���`���]����ĨӢ���1nPد�(�~�Gw6c�M+�].\���vNׇ�����'G�bn�SwWL��˥�*�%[���w9�Ů��0�_:N9:t}���^@:���z�	wN�-�����I�Q�2rLf;V+T�>�rmׂٴ�υnoܛ)�{�q����PȪ��##!��W�'ۘ�`l�qK۴�;N� ț��G*�ef���M��uKf�<�X��ݴ@u#J��&2�2�^���;�f�#g�!���Z̫����}!a����3������`X�!E�9Fg4w\�	�mQ�Q�F*�<jk��ztB�\�e��K^v�b�}Cc��Oa�;��+�)O�w���Y�<i�����!�!�WdӅ�b66f�x�zې�(i���y9�֎�J��&L�C�K�5.j���O�nT
�LP�n�1 ���BՀ����F3v!=���<Eol�-��WdL��(l�A�=$!�����Bb���ߵ�2����(����ryq�W$�]č~�W�-���pF��Lq��(B��%�����9nP��[r,��Q�j���G'Ӿ�e���YzLv9�Њ�����ᮒ��M����y|¨�S�=�����8>�귰���[�P��c՘��`v�SPw@&'��n@����Ѻ!iߟ��Q��n�����9���J�!�.6q������8��|�/�\�R+k�=X&���.��T���9������cc��"Q��`jiE�w9N"*,S��uN�ܝn��a�H��
��)��z��I��GrG��Qڰ-E�s�]�t�.1��MJ�ub��;�p���V	6�BA�ׅ�b{;�h�{�6��-h�a��\:���du�AY�-e�9���oZފѩ݋�yҪ�/*F��$d,ki��vnZ���͍rb����rX��n���$���E������:&�>�'�4�V&n2(F7>��k���\27.^��uK���;.����z�b��dM �^�l��<�]X����7N�\]�޻ʖ� �ݳF�m��t*!��Q��u-˃]t
�5^�g��N��jN�S�m%G�p�q�b���W\��.vr^u�f8�t1�+Ԭ'k��E,��{�K�_WK���H��vR5�=���6�*�pQأn�낄8Ū��ȗ���ޫ�:Ƚ"nk��j�ҋKB��#��G�:hNM2�T�#�\(�z|�_��2�:Ql�NB�mV
��|��-V	���a^u��xetա�TF�۵7�ݦ�ΏY;� sU�-r�4Y3��ʟҔ��ٔ󯬨%}�㼊U�,}��je��\��%�
��gr�vS5��1㡤���i��üZ�������heGQ*�R�����q��}�$3�~�i�H�@��{eZ�5N�i�716�F��锆���qDj)t�1:qS=�`_��}�0�َꠄZ>��v��dH��yk�&�2af�ؾ�|f�(��O�}f:�t���1ђ�#`�	��!�Ib�A9k�r���H�h1�rq�v�q�G z;�!㞋�~JjJ�o*|=}7�"[%�Qˍ��xmT��"Q:T��d`��*�s�]g����IQ����DLB�6�y�LjY��9�C�ˊ�TS>�C��=]
3ܱ[gE����r9��pr0gl$��oq����a�D�1�8JF�ƹRb�Y*=CK��p=G{�(x�fTj褹���S�mw-�ьN���؃^�pDO�)}�\��UfE�:�[%����3� ���+���ho�/[�1\{t�(EC�rF�2xB���R�/�_�
�#,��.7����0�6��֤�ئ3hZ3�\[!�0�]S9CK�L\
��xK�����Q{q���S��Sί����1=������+�D�W;��h��T����p<=~��寻�!�"�Ek{��6�>ʐ�E!�o���ق�X2bF�����[I������[%�ڛ��~g��ie��Ň�Y%�)r�]��J+��ץ`h�';1C���f�{wUPݻh�}a�Á/&��7�SR���H�m���,�x������ӻa_�"9n+����Zp��I3�~�V6�]��5=V+�����Bݓ�5j̻�fޔ�Ρ?xX�Gx�j��M�UM�q��o!Nyu ��8�dI�W��C���x߾l�p?�Yc/IL�r2<Q�9.-��£r�0����\3)�w۲i�{G�Nt^�z>�+�����c�7X���OB=��B�Il�OP[H�Պ2���;�k8,LVN�|D�O4Ц�7Yʗ��<.�k�v떂�u������X��إ���54�|�V�p��vtw��l��S*ƱBֺ
��[�\N�Zy���رzşow�B�Ըdj��N\:ʉ��U�xr�e�RU��#�]F#:h؊����u�6놶�)D�����(#�ꚇS!G��ӎ~ϭ���|~����	Bٚ����;�2�{����b�b��FU��"{�@�c╁UO>MKG	�r�q�^�/,�\�2P�u-��șem]�zѐx�VsY� y�گ,=e�U�ήʭ��Q}��k��٩>Z�m^H��J��}��T^l8��nr�Zr�. �os�����y�-�"�o|���O �{�v�N��.�jJ��<���4JXz���{r��Ek��Dk�2��ȸ"$ Tw�"b8��"4ȬT-8oz�[���9�����H�9
-g��}y�ֈ1P�.�Ъf4�=b��ݑ�#�,Ѹ��,-���<��8{TK���w�\!e�3`��5	�~�^E�2��ڵH&w���<�����4��n���y���9ɢ�<�Ԛ9b6É�3�!���(�7Q���r���m>1V<���MAn�!D�f<X+*�}c��0ܸ��y��hv�Ӵ���w30�+ܾeV1�M�	
FCs>���W�����^�1m��6����0��{�y�]�L�f��%h>��	l����q���`DS�v���x��]!gXs��ٕp�'C������3y6L�r6��j|��Ӗ�a�6���j�$��D�a�6J��T�e�r�S�;Y��M+w+�)�,v2��ִo{Qv��'^t�y�Ң#�C�\E�!îɧ�6o�3L��u�v�&C9�24rU�+}���A�۲�n���R�$W#A�N��֐�9b���J��'���=��4)�q'Y?B�]��on��������f��N'9XR�K{�b�u�����:���As�^K�R�%B���p3�-���X].d详�w[E��9�A��Wa��/��ةu���J�����r��1�*�x�"z�/��݀�u���:Y��]j���Ʊy��%Ewi�vkYi��m3`�����W��i������k	�C���+��a�=��v��;:��Z]w�la�](�.�U����h����\��VgQ5��[�79-Y�DLM ���frm���NT|Ed�����p�_p\$0�]һiZ�!y��Os�rX$��c$r]ѥ�2�Y�Ce>I#�t�f�y1�fX���n��)�M0��V5ʳb���1vl���h��t8PA^�k���P�q*u��R�D����v��w���_vq�� ���8
����Ǝix8^��Mwò�k�"0�Ƴ1�����JU.�"3�
qgZء�H]ʺi<݇��k���Q���큖q�lR���#i�/��|�Ć�۽;5E#����ӗ�i ��w��s3��֌܃���͂+���X6��t�Q=��&��#�.�#k*��6eL	c��H�:U�ʕ�*��4.>{�ϩ�Xz2)9�[嗸:{��>�xqd7��]5LT4eӑ�c�V�Ok��]��Bwz3{�`�����+u_Tk�P7��e�b��N^�����r�oI�u�A_4�R���+v/���a6�H�$�7��)Ry]�f)� ����պ��t���n(e�p�������w=g��-�i�6�4�m�vuj��=tP���SKKhJ��:� �P�B��8h��T��>i�k�P�Fݮ�:���핎>�D�stN.����ӹݭ��VUs�����4N_r����U�&�]����%;�6�U��)�9�'rͺg!�5_\@I�5PΡ�z����u�3���r��Rƣ�K�v�Βn����Q���<P�^�w�R�WK��*�fKS#YY�b��t�ٗ�k�D<UN5�.�W�g� n�8Ԡ�S*3&q����	9m�紷�ΓXn��_+���q��#1m���ݰ�D�n����B�.�|~\C/�"=�zd/1l��X!9�ۘU�M��vk��X��f���ɻxIyN�vZ��*�2��E�b��c߹��ZJW7il����۸񼨫�2���RgZ7O��W*�ۺv�A�G7���';St�}�W;Cw�PeNw׺{���dй�0��L^�5�k7�D����5L]Sn�61Z�ޖeu��\m��v:��n�ݑ�J��c���[F���N͞o>61:�������j�3ڳ��WO���K��Du��7��Ҕpw1;�V�gv��SAR����]^Ω��HOoo�?k[ED6�A��B���PT
����)YX*�0**,�U��+UDA@U,Eb"QQbŊ
)����X#(((��E#��QQ�EX�DU �V*�"�dX��*V*�b��V
��
�V1Pq�bQQA*UDDT"�TX(��b1��DQEUF"E)�B���D�aY�"����EH�U��H(�jTUUAE��ETUc��E ������AUTTU��8�ER�DcX����&$* ��Uq,X(��`�EQEV*��,E�*"֌PQUE�*�H((�Eb��`6ʑ�RW(X�[�����?]�{�q�Jk�h��E-n�t�h����f��̜ne6V	��`���p�\��?eOU��_<楢��\uYw�G_�w�f(��c�"��P+�B���n�=D����;q��4�<ƣTFU��bb켙�lut���!�zHAU�b�	��3�m�u��_��Zan,�j�fDEqk�(+m�@��xC�#I�1ƽ%QBH�JR��*'EŸqB��9�6�TS��o�'J���V:왿"���<����%�KEP�1p���$d���3=^ƏV��N2*.�WC����PN�
��b�RDH@�� (M��*��S�{����]M3S�B�9R�~]1��h�HS��~�[���ؓ�9�gy;oo��S�������b�OeLq�^J��t�E�W��a���������,���̙��R�HA��Z�D.0MH�Vj�i��A���6�����!���z�g�P�����eb�k�<a���d1���B��@�d�ГL�bf�"����Jiᣂ�=�:�3�7�c$�v5��Dh�U0����j���qRhpr*��� �[9G  ޢ��BQW��$��tю������27K����^����YƵ�KY�Yq�E�ʊ���l���kwr�y��-�E([v��i�|o����4`zq:�K���U��.�'��t8�ܰx2U��:t���ވE}��GC�S��HةN����zmCҢ��52��a9pbCˮ�W��L�M��Nٯz��:�y�q��j�e�%�V�ku�*���_w�?����`��S뎈X~N�EJ��>���7������3aҵ������z׆P��X���E;w}�7����{0�
J����Ӵ{�S�K�\��i�p�594�ʝ�C�Qg����_ �(�R�c{휸9!ܚB�z�̪���޽��J�(�`h�p�g$��+��Et��Ӆ֦�+�prĖ���N*Kr4>]�Lv�E��8�:qOi�
0��V
��{�ln�����3�{
�N�*�+p^���X��/Q��������c�7K�c�%LF��@�!qî�AxNt��\�!�Y@��P4z�m����"�bT+�H�@c�D�3'�(1��8F���*&�mQ����5�d �.\���F�r�K=���tWya<%�]�[W��Y <��$g��j�l�J�� �
�}��^��У9b����H�]9��)5xn���m�变a��i֑�����m�*֍[\�Y]v=���Oh�zَ�\�a{%{��Yާ����$\�;q��ci�s[�]:��<�#R�%	[k9�7L�Ü)U��*�1b���*S�G�
�]���V+��s+{�0�xo`��Y�-;��6J�g��+�z�)�V���k%G�i|\Z�<D�8|oB~)=��}����z�y�K���sbGA��H&t��Uf�A���G��z3�q��T�ѥk��tR�5يg�:q@�"�ߡ��jMA��Ԛg`.����X�;K#n���,�ث�-�S�g �a�m��e/����^�>3�\P������T����$���>�f͜hLoԛߙ���]al�p���5�_��yf���y�f?d���&jcYý;U��V����׵��q_�|F��v`�!�ml ��#K�}[,#�^oo`mh�^)�9Z�����t}�`dJ�*�*�۷��8XPl�E�^oش7����Ĭ�6c�{��ÃD�������a�~K�7��壳�	=0^YF�Eަ��y���z���+qe�^�hn�G=�����!D��-�2Sɋ5��rzs,��jQ�ݦvD��i�M�77J�[��F=['�)�4:F�*��,�a(��C��R��P��}�j����t��瓤g��.�X�̛:l�g��B��`��;�H$��J�t���h��j��W!���	�V-s~3��Ou���N����{"�ڟZ��naX���҇��4N�k���|��#��P���̪9��p6�؄��T:9�T��22
Ձ_��맔7��m�������<G0*@�TYQ1}J���y� %C]�Gnq�U=���^��K4и6�{�Ϡ�l�G����]MC$(��:p���[����A�Ź���g�����"�]<g4k���k�`�{�Q�b&�*��e+n�:>| ��h���wX��}�d@�i��,m~;��u��>���>Ћ�!Q~��I�.���@�O\!N�H�b�u�4yH�#a��h�9
-`�
*���v7Z �z B�����I!N
lR^Z|�{���28��>3[���L	�ڢ\_`N�T�,���5�j$�BV����Y�5B�Դ*�g�\��SC
���)NΖ>R�}+Ù2^�wRh',Fǔ�R:E3c�g60ҽ�[���O�X�EzkP[��aD�c�b�r�g��C�C�=3=S=M���"c3���ޙ��Q����MP�cޟ7��Yw��1�x?��Z�
V���)��`���Ѭ�à"�N3Y�]W�� (n=( U�w�wReiL����[�6���[7�\��(�JyW�vf`	˷���ƈ�wl*�?o��K���z���P�ov3g�M6�"�57��@���-���&�o�k`
mV���Ⱦ�Ҝ��P��Q��]/x�F�>��ǂq"iX�7�L:Ѷ��r�{U������ve\,	��|B��Vi��6L��{�ۡc �mC0o��`B���&3�i�xGC����.9j�7��T�j�2��vg�;�O�^],�wyt[s�T�� ��{�4�d�6ll�2�'^�n�dS��r��ݚ���Gs-Jy�:�ڥ�S�\��!�åZ���"�ʁ^쐢b�+v��%�cX�9����l�P]��v�ۇD��%��r�F|�������u)�A���5��
++��J
g�	�=�Sb"����C��y�w�#I�1Ƥ�
*H�kҕ�̛DI�sAƛ��oyEwUC�,���ϟ�'J��&;�̨Q2B�(>��L�	E��]�N
��S͹�m�kA��n}T���x.�dT_��t:��wn���3��*1#Tl˙ꫢX��N|c0ˍ�<pN��@ZcK�ڕ��;�w.����n�~�4	Fn����c1�J�Ν�!֓K(i'r\M^�66�׌�7q*�'(���e%8Q��Û4"ȹ�ӂ�C\�1��-PLhSM@8�I�}'^m�8�M}`ϭ���{��}�0�.Hm��nn���ad6�b=헴i�tvK��9^����>��8s֮���.����{Qrc�aQZN�ȵê�j%����0�᪻S�]'8D�o�7��=8 ҟI�A��#!a��q1C�r���@�U=ͧ�$���������Ь����B���>�8�&�
�&n2(F6� *w�&�Me��پ3w�~��8�Ԉ�!�3��"i��3����E v!�j�f��^��JMo�3u9�W�z-�{�P�8�Pb�r�ć�]�5^�S�	��ٵ9��|��}#����v�%�p,I�&ˁy�v��;��b{m��Wzv���>����n�L̵���m�9��������A�Z��3���n�삄8��LC���v��=J;es�&2��x������8��&�AΘgӀ�594��S��ri��	3L��Y4X�y��r�{(!�NOFZ��{�S�����V	��"C��,�g��Ev���mg�V��@�<ü����3�Z�"��T����p)��0-&D���t�Bv�縌lL�I!�J���yo	�:f���#{O&��jQ_n�%0!��Ʊ�P��u�R�{����'%�J&�����H��R>(�6�dR�.����_QUk,B&,���v�U��ճ|+�W]�Y��,6gk�}��g���g��WtWku���v���ۖ��X�*��c�����*lv�9l�@x�+-Xhg��{�롡�溂�_0b��/���9jq�~LJ��Q#��E�H̕����sٞ�\�or���㐨	�6x�fG��A�ξDg�mʁ~�=��n�E':J�s�WN�xR�z�F�Ic��"P����`�\S>��p��z�g,V��!#q�Lƹl��a��[��Ź���5WU\�~	�"B��A�	H��r�T�Y*=Z_9����w���_1��5�������	}`;�9��T�H<�~&t��5�)PO7wz�v���(0��ը�g�)߆�1L�'N(�"��@��sRk�
�:'QS�mLm���l�-����s��@�M�j󕊰7h_�l.��C�0���PNP��A���<a�ƽ�f�sQ�{/5��GD�;
����sMf�{ou�P&�7n�1��Xbˇ�7�I�z���.+4N��2�/P��*��ʂ���,Dr�W��w>p��E&���ۏV�<�?g��D��a0&�`�R�ϕ6F��Q"gc�y�{ٓ�.yY7��A�P��7���G �S��{~n��'�rvڎ��ս
�A6(�YC�6�Y]C�9bB���Z�[��hc�c�rd�����-���<<,��/���wd~�o���{�P�_p�t=�hՇ�ꬊ6��Fr�r�8����(r��G'�@�R�E�N�t�4��b�a7[^Un�ˊ�k�y/���m���z��͚�zt#�9�Áa�;�����c�7X���x���
�'a��;��E�o�F�%��E�Ժ}�N�H�[ؑ-��d*\s��B=9'evK���m.,/!��t�:�.0���B�ɥF���p0q��$R�ƺ���޵�s��(w`$����;��h9���`u��^�/��x(���W�q)�Z $jVL�.�R�8+g9%��Hֺ��e�ľ��:`i�%z�MC�2z}���/��8��Å�N���2����΢����dd{��&Z��D��� �e)�;�J.�0ܡ:�(���J\��F�iǘf�����n�"��C�#<�Q#�R&#��g�Bɼ{�u7�N��%����6��EPq�C��!E��
*�%��v7Z �C�
����4��`��1z�KC���\�d.�ų�[+pq����q�R�>�N�(o�Z�f�4���0N͖P��,I��̼��vf*pQ-�ܻ�<*aS��x��/�^����뫤�Tճ�h��&�s�����z�1'���]s���:Cl��ޟ��{�>���Vu�>���	�e#1kO��ݴ�r�������T8B��f�#�B�=�9�Gp:�BJj�%�� �qqS]Y ��3�݉���=7��Í�(�7ލc�ܧ-�E�����h��ez�Κ{O�X�h׬�.�Վ;�_];�y��'/�S��%/){���3]J&𜣭����PȮ(�FFCv*��>��{���3����v�����C��l^*ؿ=����>��4�Q9��'�%�BN@��Ŀ0�SQ>��,eC�����~5Q��3�O�f�2�x'C����Vi��ɲdpr5:���P]�b�n�U9p/`2w��1�L$cM��t-R)��9p)�5���F��q���۸�!q��V	K����E���*vi�rGB�ɧ=1�3L���܎D����X��QU��������1�OV?�Ha��yx=B��\)������`�eF_T�z�#��c�K���_G��9Q�ߜ�@;j�M�@���u)�A�����ȉ�ޡa1�kM�Os��4cu���K�&�a��+��S�pw�S��0u^;��J�C^o�Vm��ځXw�R��a��+ ��tp���oNq�NԹ��36�T!p�A�n�[�z��Z���ǜu��Hu@�҂z�Pۍ*V�������]��p�3��k8��Eq�}:�w�/̇�;F� pَ&��"Y��[6wjoa�*�]�7�z�Ӣ�>iև>|���>�>(�	��m)ǃF�yA����f���!�odc�g(Gk�R4'�հ��Zm�P��t:�^�	���|�r4(�xk����R^��Y�P� \d�����5��Y�@\c�Қ���N��u�|�uʭ�G�dvo1%���N�@��#�ˠ*c���Qq[#���cT�G:�Q��L�w=����O;U�NF��*�����A��҃$d,}[N&(vn_Z
g�W����,�|�sWg���y��/�όJhVC؃��B���:'�4�D�daF&�����o��
h�	����y�|k��^"!��ک��s�ܜ+�Gv���������0�C|D�}��NvwA�{B�ȗi�Y��l0�5��.O�]t
��{I��z3��>:k�	x5��O�����6�T�f����:�v:�C��Jӵ��i��+�\tL?P���K�p[���G"LX�D��u�JShf�H�u��]{�I�����z�g�-e�զފP+J�^�Q��GE@��Ý�����.ӝ�mm�p�DWO��Vݡ��=/%�a|-bAU��s�W:���&�NJ��k^�LV�ƕ��`�X,M)�3�,�|�,�wf)m�<��BF�0R��%4{a�0X p�/WΝ�S3Kg�4�پv�
uH*��ɢ�@�Q�[�r����.�D�+��.�m]<�i0�6�Cz[r��WgJ}�]�< K�o����e|��y���u��$'3nM��Vq��"���*�È��0��b�+�*}��� �ٓ�Z�,G�h�V�YͧoH�{�V}�v����E��9�=��8漴�O��XX ͫVN
���@ w����^�ɭQ8]��8B�ƴ;F�2i�W�zi�\�ƥ!��+M���M/��smj�qٓ�2)�3-p��V3U�-��ٽB�ʘ�����[[�%ǵ})<�EG\tM�Kܣ}5�yDn�=K8s���YD�s�5t�.gwEt�%����Q���S;+�����MP�N����u��-XE�	Ҳ��h���v�šs���=���
g]�@N@�t&���պhS�A��K���b*�X:��±pr���5��[+�K�嵔�5v6�#k%�x&��h��E�!.�d��o4�|�kkV�"]oE�ð����8��dW�7���sV�ձj��\(��gWIj)�΍��H��k�n�q�����-�y����n�=HN�\�I�$��� �o�oV`͇�n�e[�ʦotW] P��g�	`��"Hl�WXP���j.K�۰&�,�\��� (c��򜽪���y��1Lɔ�'j`+P����Nv>���V__.N���y�6�3���t`�c�r�vDrB��Iv�ۊʕ�h5PwqU��Y���SV,�"ޫ�h�8r����KMy�]dͲF�Ҹs��k�]4Q#�U��E�Q�r�pM�|��)k*�P����D 坵#�I���<�V������][b�e�ݤH�N�U�*��(���Qm`�o��>�����g{ ������N����+��m��)��8�Ӓ�.�z)>�&C��>�˩��$��q۶;�WM�cs9�z��|�>I�0]h��v�D��w�5v��	�YN^u�ώ��(�Ī.뺱�����K����{�\��sb�%�N�l�};c/+:������n��X�g��`��݄C��K���5B1�*�J��e�j;�]�R��;�{j�v�Z�[��o`���k�����)��۳%l��@���I6J���ޕ�{���X�7�1qѽWPX���j��xx��ZB�*����fy�n��������S+���P�i�/=�Ӽ���ss�k�t֐���.F�����О߾�W�|z1E ��ԋ ��A��X��R�`*�0(*�,lD\CcB��UdFAb�E�Ŋ�EE`�h�����%�B�)2�YXV��1̂т��aiE���UH����PZʊD�VE�.2�*̶T��"�R)m�*�,-�l�(����E����"$2ؤm$�+
$X1�Ȉ�#"
H��PQ`�XȊ�H�DR�@d1�QEV
)e�D
"�E�F0�2"��c�


�(��E"�¤PU���>@��k/��G\�2�욳F��y�Z^ʺOy��7c}�5t�*w������94�նi��i����7.�~ z���ù���!r�����h3�ҵ�����)�U��7=���`�"���ީ�tn�N��v�lL}�ٚr�ja��V����e�Yz*v	ɧ
0��B��Tf����,vR<|VQMu8�s�)9ν���H�>�$9ȡ��5$L!B]tWv�����E�_z������
���|�븋F�T�Ft�(��0��f��%�Ҋ��W^ll���A>Z;� Y��Y1��~߸M�a�1��l���NjÈw��@�*C���M (�������I��٤�'�v���>a_̚�4�&Y1��W!Uj��x��Ӆ����Ȉ z##��e�VT8��vn��U
�w!��Af3fy�����4��b|�����_�:�O9�Xi�P�<��6�1���C��V0� �Wo3�#��3u���|��Mg�m�0��d�Q��!Y�O�� ����VE&3�0�_d5�B��l���<a�8��_��u4���]�c�O��u7��t$���]Ȍ�{�ܣ\"���]#�c�`įg��8���VLCÔ1a\V9E�N!X����|¦�H�=d����1E��ɝ½`T�Cg���'̼�+?O����֐��/�}��7����Z�����>�M8�Խ7�$�q��p4��H?P��p<O~Ն%CÔ�m ���t�J�Ak��Ri�!�oT�l�����y�4�R�0��jq�� D��Z3_]}YbrmN�}4���c���b���O�����a^�~�5���8�]��w!��PR/X=��6��b���HV�WG�Xq4�Y�����u�E&�PƠ�	���详��s�}�s��Y�b�r
+)���f'�Y&c���"���j�xz�r!k���<��t�V:��FǞL��A�豳!�~�[��{�U�Խ���Z�Vvegh-�Nf�o�a�\S�w�VPٯv�`mpޔ'Uz�mui�,����k4s�]��/�����5���t�c���txJ9�=aP1*��x�d�G���W]�?wxLB�L��p�;�m�XV32qI�+:��1UIP���u���f�fϨ��R�>s�{f��^y.�NN\_˔��@��Q�0 �T�m��
��~f!�?sG� ������,�:�4�ϳi:�g��1?���L+�f���$��s�ɮQd��a�\0%|g��a�oٸFcͽ_d�K���� ��w�����o�Y?2���!��I��c=��c?$�ě���h��}�m��
�ux{�I�xü�ĩ�hz�H,곆w%z�QaFF3��U����߰~�c��>�X���^Y�&�a��T�d׶9gY*�>�+'��+7Y�'�O��0�½d���͟�>d��߼ԝ�
E�>�ɤ�VT:��/I���bߚ��Dx�Q�G�C�Ă�_p�>CL�¢���p�|C��Co��6�|��1QgT�S�)+��&0�՘��W|��ݛI�
Ͳo^w��B���g㟯v�m�]�����[�}���)6�g��~��������oX'���`|�R��M���S}~��񇩈i
�yq ��c1>E:�$�?C,X�I�ɏ�ĝB�}�g���SdA-MM�:���"<x��}֤��N!Xy���N���~��mįY*>w�N2mE�wVM�`T���=ݓ�/�{��~a̤�q1�=�1�$�Ѻ)����k��w�9���|����5�ؿ0_P���@�c~���ް�M�u���h�z�Qd��ȺgRc�C���wgY;�~>�N���<;��7gY*s0S�Ox��C��>Ci�&���^���Y��̿�"�v-Oܧ�z��G��������8�z���̢��~�k i'U����B������gm1����qgXTS�@]!��3�����O=�OgT&�L�ù�1/.�W��R�c~�x�����'Ou��(~I\�����OP����u��=a]��uRu
�xo$���|��&3��wU�]Rߟ`x�'�>f��9�&���S�x�{�>�8�胅�X����j�9�Z�K 3���!ud�;Ƙ�=uxAOp@z�u�dwN�o�2����̄�O��J'��g��v:��(���+-;�z�ea\�����X5�ڶ���g�Ϻ��ٴQ�ֱ�E�WL��̚�`N���|��Cp��q�ޓ'����a5�v�3���C����r��1 ����LY��a��d�m'�+5���H,+>�Ud�ğ!Y�Y3�Y8��7��ҽd޵��2T����'SoX����4�ݞ��f�,�a$�~�x��6G��ǆǇ�I�x�w<H,�N����z�H/��;`��d�/(La��p�IRq1 ����ǌ
°�gRc�t�$Y�&BMk�~z_{�Ѯ������k�va<a�x��N~�!�O��>I�&�?�~I�7>�������2m���8�*����$�؈�yG�� ��Fm_'71=;������Hc>d�a�|�S~�z���{�jE�aP9�LC��|ɜ�wD4�W�S��'��6��~����w�m�m&!U:�X��#�HoG����ػ�k���D�,
�?X��l/�M]0��cY�by7@�VLC�i1 ���~���N����$�Y����y����B�ϩ��m ��/i_��n$���q����T-�3�;{&�[��x~��&8��N��Һa���8�P2{Lk'ɏ�C�Y?2򇻤�
�ܤ������ �I<{�x�� �|9�I���*O���P6�"1{��f&�<nT���������̜T�����d��<I����H:�L?Q݇T�v[�����Փ���z����O�����R��W�߻�?r��6��9���?*��Iۛ�s|���G��& ���t�O�
��O�6�R]R6wܟ*g�6�ý��m���ig�i �Ck��P��wf���H��+��P���N����
�U6���P߾�dMDu|9�=�x�� ����O��!Xm��p6��m'Y��sl���w;̇����}��|����'~�L6�Si�~]�x�G�RbA!��i�P�O}�}wF2)��q�U�*;}��S����G�0颁�T�B�Z���O>�z�ޫ'\I�{��Rh�u�~���h%z��܆�g̕&�������P?w��O�{�M2��a��[Jj�CX�u� ��~��v���cBή��i��hsF�̽�3v鎷Mr�D�t�B�w}@U��1�n�kΩ��]j�0�L�-�[����1�9�oV.���֮{��Hcs9!�b�V�{�#b�����70D���7j�gf �DℲzJ����<=�{7"|�9���4�Y�?���&Ң��fz��/P���?P6��/{�bT�& z~�g%x�S�y�]��1�w,� �γ�}���XT�P<8�t{�/EB�U_nG���E���~>���E=d���)4��T�57b��B�����k&�M$��Lt�ܢ�ZE��Rq�����IyH~�d:�Vu�S��3l�Χ�ߗ�P�b�����r�v, ^{�~�ChbA���Xm~aY��!��$������(�P�T�}�1'�+�TY;��
��}a�#i6y�3��w��iI�+�M����:�ì/hf����79潺�y�ý��H��La����Si�0�<;�4B��^>N�!�T?'P��C_Y+bz�9M�|�&!]M��ɤh�,1�uğy�$Qd�y���TJ�_��;�o�ם3_�xw�yύ{�>E�d�}�E���c����&�~C�d�~�崅a�e?v��SI�'��_~J�'���z����<��h�ϑ����1��V�*J��������Y�+����~���k��t�At�$ǳ_d?!���o��jN~��
�Þ��6��ٴ����u��}9�@�N!S�{a�HV'߻�o̟�M0<��q��d�QM�E"�X~��ύ����y�wr��y���Y�8���t՚a�B��>O7� �l�f�w!�R�=�d4�!�1�}��Xu�"Ͱ����|�C��o���>M�{O��q����ǽ�R<U���r�k�<}ޯ�����z�1C�P����v�U'�W�������0����a�z��z�'i�0�}�Ѵ8�E!ϳ*O��u>C�w�&�d�Y�m�M�����}�}��w����3��^o߽�N3߬������a��i�<S�i �5�L8 c�]5���2T�i_Y:���I�*e��?d�)
��L�n���bAO9�)>v�Ĩ��?~oo=6���}�vs�����<qn0_�����h&y���a�T�Lg��I�~T��9M"�]3�4�C_Qd�8¡��m4��l�<�
�u�~�=`T�B��~�>w��.�o�sf��r�7g~N�*�q.8"�h���������u��n��t�:�O��*gm2n��3�^5�]Ϝq�ur.�7L��Kͤ�JV)�B���`���"����|tC�"D�לqR���>�[,�=z���U�P��5f�V:�no������g٥7�3k���ϩ
����
�ɾSL�{ܚf2Wl��xs��)4��C�K�׹0��Vc�w�m�C6s"�H.�^�a���ě����xL�8�Β��+j���ۯ�j �*$��p�&�P����o��1&���d�<d�w ~�aXT�i���m�d�7��ҪO�WI7;̛I�?8�L<�]�
�l�c>E�I���w�
h���]�:��;��֬}�1���t�cԜf!���|�V,��0���?%I���}�b��sL6½VN��;̇�m ��y;��Z�VM��&ߙ*,�O�AU@P>�
A��P��d�ylv�i��}���tx�e�Oh�=�+���:��8����d�'�$�*,�VL u�ך�����y���%I�b�`VuRW������]������@ʁ�L}�T�x0�5�����vm��Xm�{�ܓ�m!��;��H
)Xa����
�����d�s$*oV~a���r�a�݆3�J�f�����٭�ʇR_l��MG���}�w:<���L��kԻ��bAf��w�0�0��s��A�'�|�!�s�a�E�vyCH���4]5:Ɉ
)����!��f�;��=7f�z q6ڻ� 1��\��*�c�ͶMl]����'��4�v�C���M��q��5�B��:��y3���͆w���x��TR~;�<I�bN'�)�%b��@������l��z�"�L+�d��(���z�y��w�����6�H>��s$���T=�M<d���t�2iE�'S������<C�O9܇����?jj��q1�5���O�I����!����$Dt `xF����T�5��YO��.�>���8ßXbT��:H,⤯g��E ����omd���5�d�:�-��Hrӓ��ɤ�6����
��ýɴ�'�;H~�g�G���z��+����x�/�-�d�i���O�:���zɩ�R|��|��v�4ê�g���i ����gXTX<�4��b|�������a��y���HJ���rm�c& /���Ӽݧ�Z���`&����r��i)e����&�נ�Xx%��L�Cʣ'�MW���o�Z�>��Z-�L5��i-yi��A�Wζ�e=�ۯV��Z�/��\����t�tw�k%��a�9�A��r]X
�.�k	������nX.լ��9!Uy�*��{��U��M�~p�+�X���CL�&��-�0��d��G):�g6kX���W�Y�θ��}��)
������Ă����:�C�TY���i�'��>�}�a�Sq
oo����Ż��咧gy�gb�~�C�6�ڲbr�"�L+��A�.�q
����E��0��M�R)�Y*,�lՆ�_Y53�W�
�hl�>���<Y<�W
�����[����>n�����v��$�ěK��F��|5�>!R�<�p<O~Ն%C��:�H,�a���Y*)�O����C٪L�z��Xq<��T �+�A�o�χM��N�z�<���;8�PS�ϵ'�<`V�4�2x�����l8½d��k�.Y�J�6k�����z�����O�Cg��)
�
��,8�H,�G�P�:¢�ٛ��~s�t���u�_��m�;�3��Hm�'��t�m��1:y�>aP1*��tM�N�c'�̨�ĕ�l{扈Vm����L:°ᙓ��M�Y�^�U%B���I6�8Ǿj�3��0������ݞs���tXy�B�ǡ��Y����3l:���T\`Wi?3ߝÈm �����Y�q� i��ٴ�B��l���p�a^�7��u�&����rk�Y=q�Xw�y����z�go�<��nbn6��aG�`D{�=�4���9b�z��6�>��'�^Rިm���u:������=q'�}�H����Ͱ^!R�}�<Ow��?}��ĂΫ/ν��������+[۽��c>����$��C������Mj���!P6���6βT<>�+'�4e�!��r���4��
��{�6~H,������I�(��Y���3�{�|����������_{��Iⲡ�t����>Vy;��:��Ă��L�3�=;�L=aSӳ�6�|��5���0�����Rc��&0ެ�P���I�Ğ!Y�O�{����s���*&����U���Ӫ��=��O��'P��?s��*�:�����
M��>s�0�ԅC��gSl?3�ğ_�+<a�bB�<��Y+*|�uH>P�e�i8�<����ʧ�S���.�os��"h��$՛M���b��}��4>��a��|뷦]��ޕ��H�q���}�.�gt-���Dp�N�����X�r=����/��{ʥH2�[$�f�]ٳD�E�z�v�(�w��Y�s1lbἬ��  ��wzM1}����m
Ͼ�� Qa�5w�㤟!Xy���N8��~>�@�+�J��}��&�^����q<H)7�����'��P=��a��2�I���q�P=10��E$M	[1=��N��tS�R
N��q��
�կ(La����OSI�}>�Z&�2TY<�2(u%zèx{��vu������@����w����%@�O�{b`xFu�C~vby͜����ᮟ����&��Ν�i�XWm����X~�4�Ne�X'���K�!Xq��`i�0�c�~�3�ugXTS��`���o������v�m�{�[�S�Ќ�'���_��m�@�;>��I_��&3��E�+�o�I���G�u��=a]���GT�B��o$���7�$����X|�ꐯ�=��'���z�L&�����.�n;��s�!�w�����k�shq1H>�ý�m�<N0�wY:�I�
�v��٤��²z�O���K�,�q���!��zɹ�`��� #᫟Wp���Ğ��7����P9 ��4��Y>e�'g`m���N���w<H,�N���z����w!��VM�Y�P6��_P��%I�bAM}UI�Y*,+
�RW�8��:��u�1Uʶn�.�Z��i�̗�d<aP6���NnβVs�E:��</p�>B�̝sw�;�6���9�~���g�At��QAa�ˉ%VT��)3�B��y��ۭ��_��������߰�i�0����j�egP�u�L����<����H>Xy�wP�,�
��ό4��+��&}�C�+���*O���3�>ߘB����4��I�W�����@���|{c~�Wܒ��Ǽ`
�O�PĂ���"釬/�8³�c����tea��4y��H,����Shu:�$=�\��f��O����u
�>��w!�����c�����ѦxD���]c����=�~�Ɏ3S�4����o(��2T'�cY:��]e���vO~���&�V�M~��O4�Þ�^$�������L�T?c�u�
����~��X�=��=�X�dU�gY�p`��b���2Xb�T�-�,��7��	˃�����pG�*�*�:��l���U�q�ҦO�^��5�!WBc�Ψ�-�ba��C,�q��|�s͙�������z�Fw&������m!��?���x��A/��߯�&0��?�~��m&���:�+�%E��%Cĕ�5=�Civi����0�J����d���'�b&���O5�^�c£����lTt|���UI���;�zst�Af��}���'2�<��4�RuS��C�.�
��w'ʆ���0��i�3�1�C���)�a��
�Pă�>E�"�0�?[?%A�<c�G�QY��R���\�#=ٱ����8���~����c�ܓ���6��CHF�q�9��=d�
���!�6��w����~y��s[hݸh>��1y��iP�߮��*�n�$��FF��ۿv̦u{��3^�ʸi���>���{7�b�#f�E�� ��iN�/C��4M@�z����a�l��j��ۗ���؝r��K����'����z4z��a0X7[K�ޠ�S[4�1�ni�d�$ofi�f2\��&�����>[�~�v��m��v'����^>���'�
͵\*k�RD��X����g{F��~�ii�Y�u:Rv���mL����bhl�|Al��� +󞬲��w��w����A�9W��i��qH���C�ͻ�ȸ@�Ζ[�f�}l7�n�jk�T��$�X�s�TZܮ��U��2� Z&:���&l"�����Y'��}��eq�u���@(��o0ʲ��bQwZ�A�6�+j`�(D^%s�i�+��u���H��b��و�Hei�w��W7zv:���l��C.jȻ����#�q��W���V��ʝ%M�y�t���t����y�ՈqA]~��7>�{^x}�7
�xF+��	S����s˧O���z�������r7�+��.њ��%/N�r	��D?D�
&��5�����@�j���5*�7[;�Pլ+PW��m��s��}a���i�"|��2�#�̉1�E\�]�Yl�)Ǵc��w�J�.��a�
���gs�
>�0�24:QBjr���Sp�y8�j$5�V�Q�s�����Q�8C�7�LS6��)�W!�5΅IB=z#n��������Ogb��o�mNϒ�Q:3�2�H�b'ͪ������:\L���M�Nn��ϗ{P����Q����0iqh��P���Pb�ׁ�\z)�E젡*��M�N/w�����Z�h<Ή;��q�T�vَ;C��^Y{����o��D�������&?W�Bu��~�U�ǃV�NW�8�=*���<0ۯ)[��p7�
籒#�8��a��y�7�Y�M�����bA�l���Q�S�,(���nE�nM��1K8Zd��;Er�r{��V,�e��N��M]
�Ȝ����Y�����a�}�D�6�_w'pٝRÊ�b�V�W07�Y�.ΑMB��ڦ�7�	�x�OC_h�p� �
"��&�2�Gj�C�H���s��w�����d�<+8,n+/b��z|��_ �(�p��Qyװ1��=s�d9ȭ����g^3�g(��S4�|�@��*��.�/t�8 �>n�شl&�ň9ӈ��q�
"9�r)����Ju�0�}�,H��m�"��mJ���i��f�E�b|�X�n����OǱV�`��ѩ%q�Ӳ�=F� �!��J _u@�._J����#��-Ua��:�d��]9��;%E�򜒄lgx�D��� �t��m���*_Y��u�B���mM�)`-��^nt��}Y&�P��0��T϶Ap'���;|�J���X+Ssi(�|�[gE����rPNn_���1i�"B����hI�r�]h&�i����0�U��`u�G�$F���{*P����QT%��A����#8)���;+������`�Q<;���Ҫ,�I��EP�F=�N�P%�w�r@�Վ��aj��h��-KJt��:%3BM3�,IȚ��U�������L6�L`�O7�����<�nUe��m����Z��]Z��1�5�VkH=Ө=��JI�r,huO�k6�N���!�
��T^e*'z�o;��hڽ��I9�d' 
`�G�Z:�06�{�V�s�l]]\}�eY�����\��.�s�d��Y�G��
��������Gq���+��t%��3�!a.u�8�ͮO�p���mn5v���^�:Q���.tS��$C炒q��]!]onK�.eL��i2��\��04u�i���aǂ��}3YR�;v�e�	�P�v2]p�JPPok�G�=�K ��/�ux檾�\�YulT�6&��e&2�.4Ḇ[T��ג�Yv��H�*RP��X�b��QKŸ��t[��c;u��O�W��y��Uў���H�K��gR�T��J*h�.�&�X�������5��]^�s �M��:�I�V���p�W�)���n̊���+4���i=p�(���a"!��<�s[5s����W]��,���9�Q�u6sW���dW�jd�v��D�۪����%m���M�SbȄ[�A܎�����
=75'oY��g���W�����Q6�H�<#I��x�M�
�l޲ĕ���)2�uu��:ޙi��]�!g@��!���{���N�%����]!qg�V��m��I�B�d��#�R�e�C+G]���ŝ�7��:VU�������\�=9@j��
;y���K&��j����1�l��ӛ�q�¥,��sS.�s��2�7����qv5��O	;��:���{�M�w���m�%��3�}!�y�����Y�8�+�}>�+-���dG,t���C鐑�V\�Q���u�CQDq���lދ�.Q��m�6\�g
�\��� pe�K���}h�ʛZk�>]�wt��UHw�I�T�6^�W��E�"`���v����-
F*���B՚���IW�j�Zi'�C�Z.�+l��@[�8�����	cr��l�л=*�����M�it�'v���jf�^n������2���leg-��� �L��%��R���r醷6V�M�nΣ��YΔ\�brC_u�L�� ��Xs\�p
�4���V-m�O��d��ru
䎇Gd��3V�[����V�R��A3��p{:�D2=�㥰��uF�;���ͻv�W�qIv+lvW\�*�K��3t�imZ-r����w�XO#�U�.���;����t+.Mv+����\8��g�����#��r86n	I����#�8IYgn�^����S�`w���qA�����'/s�{ƺ�hf�Ax�`���m��(s\�\M@Wc�9ũfC�M�1���[���t��4�]��[YF�,����<삞0����k5mΦAyik�G3
c8(�Y�{5n�v�}ֳ�=���
�x�U!C#�p�e�ϧ=�_:�)? (| U�m��b�
*�QcX5
$*�ъ"E����0�*�DT"��
F�("���1UDDd��EAd�(���EH*+�b�XcLlƪ*(��`��\IX"���TE �,EDD@EX",��mPb
���Z�Ta���rʫQ���QUd+DT�FEQTD�֫1*AU�PH��Ub�TQ"�S�1�V
(#����rЈ1E�E+Q`��������,PX��2�X��U�֢ŌH�EX�UQU`��UFe���EV
A`��Am�X���T-)YEb��hUP � �|D<M�ح�yw/�4drVK,�}�K�j�_vރ�h�l�����NW��VR���,Qg;r�B�T�rD!|���������N��&��}c��D����|xkD�tP�t��И�M���^��+��{����Z̾�b�gjٞ�P%��e�jofC��u~���VA���#|�[���6���U�h��k�*���]l ��#��X�_{���R���t}�ѫ��瑴DγAqy7�,��Z��g\��A�
F���7n���E阸�Ȼ|{7���C��}N\{p�;=�U�IOF�rPG�Up�[�^v+޽����H0T����c'R��'y�#c�KG*v�_lӁ~�7zhSr����t��-�E��lk���m�p�!��['�OA�Cjf|	B���ܚ�;ƙp�;{#��;���iv����X�W�T��22)�28N��J�]H
R"FK����Y9-rE��"-1��lw+���x�ӎ�#l�Z7�.�%��Θ��BJ����S��bU��]5;x�q�£ݻ�����^<���y���ʍ�S�8q�3�"c���b��͗T�j�FЁۮ�R���t��}Md��7E���Q��_o�Vݶ*�^�+u���6�����sqxkCd�I줈�k��e�*�]������]}�f�p��ڗ�}�4ۂ��V���h���u�68�R{6_d�t�z)�tc2�v-�4���+�*7U~��=�{�ld�j3�3U�U
Tz�\q=���C��f��l;>�H�>����<�:Q�Y���9o�C��BL#�BHجR+4�
/˄�4s��~�q��	�*痔�2rI��� ���˫� (`��^��-�g/g��ݦ�{T��T������b�Α�Oylw���+.#��s��h�@#L2$���eL3��	е^G��t�Tr�nT�yI]�1��aa2w[wRS,F@�.�68R��d(�$<5&��޶8k�6!��#��`m��11W��)�g�9So����^�T��8��7[J�*]i�)5*��G�L���Fľ�(*w.��1ӭ�(4�S��ȼ�U|f�*I��J'�����>�����VH�pn�{mRg��>a��Wt:+Ϥ,,VX��q=*�vt��ɺ�1Lr����X���
�DF#��}V��qz�8v����h�7�§7_*��=Y��F����_��*�����Z��E��m�8���Xp,5juUNNw�ʵ�65Ң"$rwe "r���z6�����g�s]��:�M��i�'_�>L��g���un1%<�6��K�u�5aa�ֳ�\0F��j�"ae��Z���ĭ��bs��f�!w:��l��J}��J��xxx{ލ�Z�(rh�QＺ��9	�^j�V�sл������kPuS˅,��˚�WE(t�7��?vWZ���]�b���ǹ��F�o������g�;}��
r�]�T��x0hz����T&*�Cf�Ͳ��}:�n��.�#	���7q%@Ĝ�uGm�*�/�P�$lSr{s�T-�y񰜨P�1��u�2�Ơ���qԶf�MUdt���t2P���K�N�W"��"�
}]����O+gFD�y�g�OP�]�ˢ�9�"D`@�� �u����]�t�X�=2�8�ݦ�qt+�����E�c����v�\��>��VIL�4!*��
 �oԈZ'��(�2�M�+<9�[���\C�Wƹp:Ӡ�ܾˆs��(�/�}�҃$d"o�v��;�If�k<5��bz�_@�
\��LS)��5#b�T�#��B��v����s��.Mq~��ȡ��3��w:�/��Kj�('>ȯ55fX�;Ul��5�~��j��r��w�O%���O���{e�A�/7K�]�YYݭܶ�����u,�:��m������z�^���&{'mrt&�ж��	�>fn�j��cV;�/[�%^e��9�r��OX�"���֩wl�x:NwU,���=��Y�6��|�lT��"�D�����@��W����a��]A�r���M����V3邳~_lW\S�x��t"e���R���G0�R��Y�����qC:f1�6,�n����ݕ��+�j܃�����.a��Z��_�Q��53T�櫮zqi���t�Ŵ:Q�K��&�w)g�1F�
�����!���)�B�N�@�^��q;^�-��T�</�~�4�=�ʜ[9����yװ07=���D�8:�Z6�I�c�w�
���#L\)0;]����瑟7z�Z6��:q�J�SPm���w����T�=���
��$Oi��FZ�H�t��ΛN^�p�u��ϻW�����&�*={*�'��#�R��Um*�+�<1�*oP4��U���65N2CP��䝊�8�w<]�1Bm�$b=	���z, (�3BvzͶ�ڇ�4�E�K��<!LF�<��٨�z:o�;��*/VI���(�A�r>�tx����\ ��J�4	��2:�=��v�V�Mwa�o�}V��5&�e��%��#M��C�C�J�}j0�R��9���KF:��w�U5>|��It>լ�&o)m\��[\��o�V,�m;�Wtڪ�������m�\cg�g�Gk#c5c�΋!#q,������I�	�"B��p��ǆ���A������'����MG���=�P���)P�M@�%��١:U����c��S�	�KK���~���C�J
TO�M��P���k�hSQ����T>�3���Yʧ%95�y��dp����x��L���>�n�vȤg��q��8s�T"�[�u3{i�Փ1vxaB���O��&}�n:+�i�fb������A@�Z�4W\.�ɸیK�i�����XBˇ^,��)�A��/���-"�*���`c�����j2YE#�����y������`_�e�w�u�����#k� [ŀ����|��aU���`��vm��Y�u����F�Ht'靆o��Fs��U��t����ޞ��(h�PC@b{gyU�Rܱ=�w��m?�)b�oW�'�M�E���=������W���5�9����)�A�-��#j}+�L֙���&E����[9S�:�f���Ὁ��n�wu��YQ7�1�&�G��/�Co����U��%{fA-��U�v��3$�eN*��E#W�M��u:Ia{�w]���`�K��^[�5+��"�򔲑}����*ݻ���xp
o3��:��[tl�5])��Ӻ�Z���W��ͮ�ܮ�n������w"+y��*�>2;k�$�Z
u���CƩQ=A�V��f���HJD*�t�m�+R��}��픩�s�z-H�,)�3���BP�
H*]���(32Y~��`C��2*8S��
@��H����Z6�Y���ؖpup���yK��"۫آ<{��MBbd\zU�b�߭ڋ������W�x`�*����:���CMi��bD�̳%ƕj�.]P��N./�zX]!�p㣙�s��'ہ�"��na��O�9���� �Ub?X./��LG�#b@�T/a�Q˄�4s���~g���G��p>��c������k�1P���0N�P��-�f���n�g5I�ZpT�0�����q�;Zܘ�����¢�|���5@�@:a�TV86�⾻��"��ov{�̶[{i�s�G��PQ`k�E�'u%2�d�U�tӭ���B�pH׬�R�`7s�א�W�#n�*㟋��c3�خ������)�Q1^O�m�szg��L2'
��q�)�D����/z�`+5���]�hY�݈r���bA�w[�৚��r��|�w�J��	f	���<�߷	V�{l�9�t{�B��
,�>�5nR�xv
�9�ʝ\R{^ kq_���t�y������v)P|@�Lk��X����G�?�����ᅌyw�m;�	���Bv*��;�Y#��,CA:��T(<���jkL�HSY��Qˠ�v�/���^�,F��
W#!��ڿ_mSg���v�j�t:2����r:�>��I�;��<�2��d���m{D�	%�QBMѯIlƛ2U��
���{e����+Zx�)��a���o�ݮ�h�j�%�`��^�P|����jR?r���o�m�]�6���`���C���,l�iX�y�r!��Ү�[>�1�.+�vP�u�V��u�3yp�r��0;dlR��PD��X�j����E�p��1"�ϛ���Rm���������7頻�S���b�1W�65Ͳ���E#��Gsn��ȸ
̅�[Ёt�C�]��	o,$��0�'�tPC���������)W�	ʅ`��ݶ�=vFtn�譺�K�7�_���"�� o����#��3@K�m��<��EE���uN7oj#{+(�A%����>�
ʎ�1^JH�@��A�;u5��-P��\)t�v�a��t�N̾�d�<T�oe���T��)�;#���!Z�!�u�<�M\�*q�����X3D\�]yGz�v8��oU��]FT�z����[��@�e����MGs��}W3���|���4��h�c��
��;z���P�}� ��G3M,V�Flf��p.e�B.rϐn�$�r���3� (�G��cMnq'Oflm�+}q���ODX|:��R�u�:
���g�k�}�0�24:P�J1�p��]&�;�/��
5���co8�!ӛ�&)�	�hU��s�{�
���a:2���ذ�ou-��3BM2��dTcS��gU��u6^"!�����_XxE����yS~��މn����aM+��E�ySu,��=�/1^�ÊD-٨l�k�1*�F9�Q�n�K˳w�#�#�Oھ�s�,�WG�����Z9�
���C¤���0�Ld���I����9=��ݚ��[�����>������|Ҩ�<R����ث���k��xpļ��w ��:!F��LC���n���U�\
�&��Ѳ<~�*�GL~3���/=�$Ӿ�S���Q�=>Q@b�e�N�[9�����^�K�|��d?s�]=ղ�WO�
o��Pǐ4��co��>ҩB�p{L��t)MS��h츣�k{b�#�� k�n��\��~r���F�������~��8�"���ݝ~j�ȫ�+��sEc5�c� �J�|�v1P�������|9��8�Xju�ۙp�o�����R���@@�J�\���������(ؖ����{����;��5�o����A��r$N�~�"}j} m�TlgM�/Q���X>Q:8j�-�w���5�hsu=+1ђ��;�� !6����tD�𬚸j9�ZԢ*�W�G��u��J�~�H�X���S�U�;��p�d dN�A����*	�	M�q]]�?G_J�t�ä́�t&t���$߂"`��x�G���\�k�Q�Ssw��rў��(�P�=���5#P�NB�9�m�䘴��G�q�Yd�vC<.�r��ĘnzL@�Y=�/����:�r�Աd(����76 �-ۇY���V�=��U5C5QU��R�p_%C��d��+�~�F=�'NB2�X}Ug���|�]�P	/(�*�{��_�
��Z}�Zj=��M��x���CV>�8Lj��X� LZΩ��)�A��|W�J��)A����f��9o�=׳Zݨu&�[gy
�;�Z�j�0�
^��ٕ�S���YG´5(�<z�vW;����|E<����Xѷ#����������D�e�\J���y�H��Y��<ұl������{�c���j��ٖk�<�V��Z�{T�34�ǅKiRm��X�/�vZ���q�3.y8�[�(-ޅ�xp��;��Um�Ρ��U��� GQ�:��-���$�F�:n���B����C�=�N�]B~�c���5��g]ҭN��KB��3q��n63y
p��u ��(R)��pn���zf��Ol�k�<��aȺҌ�Nż�W�&)9賒�=��\8�W��V
{&l4y�EA�U[��u.��V#(�q<((�@�-��N���N�!�w�4)����f���;�ݻ��U��~s#����Og��#I�@�OPT<0vYZ�+�����m��h]��=#�P�(Z���	̨�Y"���=[KK�xtj�{��z���˛�z���}=jݺ8�e炐:}��#o�дl9u�/"}tƞ�*0�Tj�+z�t�^�`48��&B�m�S��o+>?^��̈́v=6�����=�][ޝ��v���;�`H%F���y��jZ8J��^�>��|\�x<�e�Eʬ���]�w.��|��@�#b������$lO��it_�	�h�RX]1�3P����m
S#���{�zgHQI޾�Ԭ�)cZfm㺺锚�W,jJp3�'"U�P�d$�>�݈Mt�H�Ј����y�5�k��i1M���K�2֍6н��rف� ;7��.�@\�A�46-�}oݷ��ۡ�Ckg���t�w���ǲ��o3t:j����2ܠ�ZTb�C�hsfN֯2�#�Z���g{,�a���oTTv�v�9��L�G�����z�}Vs�vqn��fg7RžI֬u�Rv����5iTˬ�rgȰ��Q�;{nƤ�I`.ѷ��qI`衱�=�[v�7��*�xa��i�@_��`�o�.nX��+a�.S����;�sL�}1��u�5V����q�e�-*��l�փ��wx����q��A��z�`���Q��mvѣ��TT��ק�Z��	Fs��
�"ZƓ�/\��u�p�,쾺�hB�ԚÌ0�@h%��T_68u�L��
e��Qn���[�N��HRK]v~��z�]\ ���,>�r���$j=2��{��кȰ7Y��5���77!i6�#���)n�sl�h� �X��qe�[ْ�R��A���N�5l�qX,کQM���u��L +�e��,)��l�A8J�C��*��Q��S/N�k�YkDũ��W�΄W!\s�A��,v$n_n�N�v�f��ʅ͝�Jл̦�ҵظi�dw�:Tm�p�L�a�R]Vv���f��hJ9y��G�P�oF���7���wue�uU��T{q-:�1hWV���O~��^&�Sk��t�S�ŋ�|���졜�e4�厝cj��&����ϴ�:X�D�j��gJ�u�����#V}&��>���*Л٭�{/�$�_I�ˢ��S"D�Z�7�̻�r�Aw<2IV��L�Yh�v�.�E8ơ7��Wy��t���fȯ�;c��ZQއI�|��p=0��n�E6,���(��G�pq�U�34m��T4�@�����za������k���>�wP�)@��e��c�)C��A=�Bgt�����W�)=�Vh^Ҷ �s{�9���:šQK�N���ի�Ufs��&����@����%M
��,c�T�x�4e��x�Wm��U�`��̛m�?-�L��
	d�8�[��v����ed"��D�W�H�~O��z�x
{�,��nN�id:�;�+�%�V�'mYc����uf.�֥۴m�@���Bh<y����.�Q�m�V�
�pun��!m
�bK%��^޼t�`�[w��t
oml�b]gr�����U�cM�ds��F(E.����J4v_n�t��q�y���y��G���o-�%n�n;겜����g</t�!���10��穬��a����vV��;8�O��٧j�p}u���{ԫzێ��Եo~�{��\���i��Gp�Vϧt��;ڠ
P�*"(�b�QADQ�����TTU��"����QQQ`��(��#DFe�V6�Eb��
�( ��H����Ub,Qm��(*��b�b1ATEV1DTPX�Tq��W�UET( �ED1E-*�EEUTF#b��*&Z�DX���5U(UX����"�E�Z�b�(�*�dAcTEUEF1c�%���"��(V��+*�PUUb��H�TX1"1��TQbc�dE`�Q�cX� ��`�B*QAH�((��J���
 �-kŊ*�"�DR*���{��ؕ�9�Z�c�#��.\��M1�R�5��F�b��:�]���������22���r��*�F�S�vO��x Vt�m4�c�?�;ב��h� (�q1����37���M����[16�����vE�#�y�u��ޟ6|:|��{Ʉ>�X�O]��T�7n��-�rL����prtK�������qc\�/���r�lX��i-���V8yf��p����g5>��$Z:�M�cs;
�ʭ�X��<�(����[5�w��i]�`�T|��=�����p��)���##��{"F�+���\U��Ӝ��@<�����s�p�����#Ĭ����_.MвX���$�
V$d87j���M���0�{�*����[�f;ə�m�}t*̑�j��i���dhr7A���<k��F�#��Z]C�Ek
S*WD����i�H��T
��6/����я�i3W9G	q�bT��L�!u����c	YQI���flX��9홦^���:	�Ns�l6�b{'м&a��*\SQ�K���C����/���$8Q�]8j�]�-'N=���rZ(�z~�.�׼�\��.�l�ǡn=�c�k&��{����<��F�s�u��4��l�m�DH�G<��}�
��NFBP�����.����ݖ��g5b}5M훣�?4�|'&:g#C�	f��ZҊ�zt(�\"���媶_]~���'ns�7����AH�4e��1C�P��}!2��f�X\DR4>�۫�3����u��T�1�ұ�F�K���D�� ����������J���	�P��ٴ惗eV�GxE<�O���`vRɛ⢤��d7���%�B��*}6��]1xVڹ��cvt礓��*ޝ�F�����i*�q�f))"$
�::4�yS9��:6�ꖏ��Ｍg@�5���=�Uls���>nf�NA�B���c�ʝ�7t.J���Z�liad��'�D_���z��)�VK�f�)�L"	-F-��/��4���jB�d5��1]���B���ͧ>Q^�W!�1˒�����f�lR�J�S�&K�}3`I�C�3q�1���uZ7�U</��HmT�9Y�\N��1�0j��>�#S�M^�W�R�K�T>�B
�����Ţ7L�`�+h�U���;j�׮֣�cR�ć�]����C�ܚ������7G�huҬ�0��ʇ�t���5����ʠY2�f�KE��jlxw1n�̗�`�dպ����[t[Ղ��m ��wGQ��{��K�p��z��,����vYܝIX6��R�WV$l��X�o-+�0Uw�|�D���K�`{>>=���Ҙ���eZ����Ef�]�O�9Y�?��u�^B����Ȯɨ��@��O���Ted�.|��w+�X�}ЅG�j[�F3(c:�����;8ȧn����^i�Ƚ"h\��L3���U���=��=��/
9��KÖ�j���ꎯ�m�e�}J-��NE�`cs|g��l��F����/]򔏲�*+A�4$���Q���vʵ:j��g�޻q~7���y���N�5"��nv��5���eq��}�2�Kf:�PB&���Tt���Fn�P�86d���cy�]�+��]�а:���1ђ��;xH>!q�*P�JA�e@�lF����j8����w���8��bT+]"Es�h�*rJ�b{�¯L���o�A�9�H挼��L��WȌ��@�S���vW9�Tc�<<��+�D�"��Go\�Y�<��;8Y��V�V�ϔ������r�m��7�r5�s��wy&�C��/A�Y����o����U�&˺��Ed���⣂�<�N\;SP:%�_X�y�{XI;W ���Vrv�F�w
;�K��n(q,�)����O��Qp�0��\I�*k��"$�8�M�]�x�6 �#��Jn��JZ��9�n;�P际\�z����fcWz���18����v�t�YR`��B]F���:�v�M�fN+�{�6�s��6�7��\A�p�I�8�D3�T��l�(
+�Va�뤐ʴ�[�ꎦ�tOC��l�:�ׇ�ΉlГH��nۡ:;hZ3�W��S���(��j��W�d���xaLA�ό����'!E	�Z�Q�,B��X.5�P�A�3���^���`k�1����a����*�p,q�*"w9Q��Ζ�k������g�ۊ�����=�n��ݦ!�:�bۧ�X�Ӑ/�f��X�DuEۥ���;v;'\���jHȥb�!ק2�lf��g�P��-	�Qa�w�A�u���=��óto��q�J��V����9.-eW�6'�A�A�5z�φf�H/fIr�M�Y��7��-j�G�&@�}s�{	l��
��4�l!��[�:1��؝�x4�(])c�V@��S�H�9%]%`��3C�mL� O�JBt$w��#k�<hV%E��E��"YW�P��	T��9��v�t'cb�	p��E�^$k����WgR�ܙh�>4�}Օ-73Xp�z)?ne�X�K��Ba��E�BV�H�mK�ݥJ��� k[�떑�sY�N܂E|U�"8nL�̵�K�Á蹇z��0v-˂˹Q��ۜ1>8�5s�gaMv�vrٓ]v;�����{�S��4�\� +����zLU��tq��^yH��v�mжmˬ�x'ƅ�d��Q��������Ò�*�MGP�=>��u߱ڋ����6��W���(��3��ժr������o����H�	]7O��Դp����Ϗ���r����F��qQ�g����En�k���c�VP⠈�
���	0ʊD�N*X��Y��d�p��9�pR�[�Se��u욦�A�=K�X�����V��U],� ;���ӵ�>�*�ˮ���N�7�R���I�Zlq./��ߪ*���/���t~�G�#ǃO]��A]�Q}��I�<�����޻kU�z���8�L����`',F��,A�"fm>p��'D��Q�&g���ǾF�I��8����T;�ʭ�_90�y�Q1A4+h�noL���6��1��IL=�s�}XŚn�W,X�O�����bP�r���N� �ҩ����p���W���Z[[�loU�*L�A�͉l���FC�v���T�=�>a��c���сۻ��M�&�>�%��3o��g7��K�M��;�����
�����B*��L�zm�!������Эf_���a���!��׀�tw�b
Yj>�Ua��/*b/&��.��1�,S���f�b�3xv����u\�ϷS�u�J�E�����P�Y^U�E
���m��>�6�x�4lZ9�'E�Ԕv�a���\
w�}��P���>�����#��c�*8W�n��Ѩ�����ׯ�(di�9��4ofi��'^��&Gx9α���]�k�&�g������Q�m�V�ul9�B*�\�(�.�'K/X�K����s�#�g�=�rh7�F�[+8v.�pa�>�p=`T�$Z����L_�hq�eaqH�>���Ҵ����{��۠�v�hn�{��7�I�8��!���JR�sʳ�mK�����3)HI��Z�y�+�v�`�	���u��&l"����{ %�;�7OŮ_Y6ow{�����]��oH�u��*�[�u�IV|6���U�x*\5|���ѧ�	ڭR�l�WZ����A�;�h�z���ѦT
�u��K���n�$NAG��\��>���/6��Xr�iץu0���ظ�y�ˇU��S̅��d���x8 �
}OZF���S���21خK���+��9u����5�n�4JS]�7x��Qw���d��w�����o��<O	��ܢ��o$٥W[;��+e`ʺ�$�-��$�?�ͯ<�r�\����ʹS<�Xt�{κԥ��'[R����\N�;yQ�u�E�_G����$�2�W��du�@u��b�ٮ�d!
�ߵɊe3�B�&�[g��<�vVI�������P�48A'8Ԛd+7��󦑼R��"!��:�]���y����\�=Y���N+eEI�Ȕ@�f�fb�ff+��.-��^�f�6!�m��)�]�h8�G�1>yu�*گi<�I��W	�hI�&����M��M .���:��T���0�;C�;+�W�������yrN�G`�C&p�5��soc��s3$��;ΖjR�����賂q����;�;��W��y�Y�Mz� ���+S"1�ɴ�w�Ha��]EB�.��aМ�p�8�Fv��^y�(�pE'"udC.���*s�GC���]=|fߧ��98f��0݊5�iT�{���y�|���bw��2��G��]͵�yp���,��08#��6H�-�鐄`�>u�4��ΛN]tKv"3F��a���=�}jT����m���UV+�xm��'r��k��%@vt)�Y����5c;�[w1�o��J�����3�P� %{�>��.�����*1Z�mYBh�-�#��5�9��q�Fuo�%7ĭ�؉���+����gM0��܍������}��[�&�-H�}%e���!-߇�En������iTs���J�c]"Es�h�S�U���C���Gt�=�Y'�4N:&Kk9򵾴L����i��6ܨ)��u��Q��*;VI�"&
�@��8Ü1(<��lv�ؙ�Ip�:zw���jF�Yń� +��LZ(eaNm�Н�\sJ�LG���^��X���G��_��y���v��d(�E��Q3Mz�<�z�7њ��Z�D���*�cN)��'�{M��EsP��s��*��ar{��+��
��U@,��{G�YK�.�|pT��E�v%�����q��x�7�i��ؾ.	�͚��'(iy�"b�P�><+iX��?<�A��ĖJ����7.6�3���5^���ޫ��5�E��kh[3�r��R�>�z��<X���ȉ�=�˃,p�vi�Ɲ����v��|�a�n�~����a�֙�8]����QJ�A6�7ʨab}��8#^�2)X��g2�do���P���<;ݒą��N_'r����ɝg6��]u¸�Iy3��8����z�6��rW=q7K�;�Ȅ�}Xoe�j־���e=�Z�cd�ipL�]PG�#��s'lYR���!I�T��T�2V�eY�%��/xVrH��r�)9ٯ����}T�I�X�����#b��|�D�#(J3��qk*�1")�=�w�*�p;��L^o��29�aߣǪ�9��ڸgU�IN��}����V��g�k��+��)���
�|�@�OM
�8u��q�dv��%]%`��2(u�3�P���T$r�-̼�s��tLk�[FƩ�\�%�~�(ZN���z-�j���AN��YfЮ���3��ܬpތ����zLP��n��y� WP�h�֝fܺؗw>�$?Tm��d��7�w<>�1@�1'���SP�d(����n�ZyY�W����{��r=O+�2ɭg_���B�LM�.
C�T	%�J�m�E���B�]!�V]˞K/<�o�n�c��j,oz�G˛
5�[�qgڊ�"BD��F��eE	"tМT.ƗAF�ɢQ��lBE��v��;�0-����qub\t:������C]C�e-�!��1�����9�]��L�y���8���p��d��<5D��N�<�`��\�&�MDǔH��x�q�s ��of;�{;��>��}ױ�#�U�g)V�nfWdiy�Ω@/{�3�3m�(�&}�);'E�dN�8e��]���S"4i.[��N�.���-+�P�����n7��S[����n��Y���%Ž���ņL��Aѱ�j���a�g�W����>��
(�1ҹɮQ�z����M�j��X\5ɢ�:�<���ň:�L�QGq��i����$�sw��a�
����aV*n2�2�b�gb�\����a����O�x�W6,a0b��2��X3J�r�CƔ�iW�cލ�ae�^��R��1ӭ� �3N][���4y4������eΘ%�{�Ҝ�u	_eL�ĶjN@�~���Dݫ������z'�Lx���{���ʸ����:˕�w�5BVW�fQB�~5���~���7s�C�,nk����
,k��;r�S�O�b��P����4���� p�[1JG'�et]S���K�sY'�w9��!�##jniGd�$ofi���[�Ȅohd0ڮ�Y�B�Ms�vh�⺵F�
�5!R��%O�nT�(��v��%�z�W��Ǩy��K���u��5�����׎���l�s��!S�cc�1W�/=�m�����A��gNDu��(��k��F�گ [#�� i9�f8פ�"�w:9{��\U���n�aMa{�Z��y+����F����6m�1��Z}��p���*�@�gH�\�H��4n�p�5�%�K��TnP�e>��7�lOM� �厙Mm7`K'��.=m��ڰk�u&��j#o�$u��]79=޻�R��$��4J�n�_ЛI݉���]+M���j��ۢ󄡫����<�SC�d�UwV,&*�B�\y��i�N��v%AS� ���Q��N�/z����:2�!?	��t�������8�՗n�A\D��_�!�(�M5��)M����Z1�E���.�^`�UuZ���	�z����@��=�R���B��FWQ�do:�"+����V�q����A₅hd�=��{�w�ܻ@^�J��ڻw*]��0Pz�8�����F�;;e���J�e�Mu��1�
2��t��PH|}��ׯ=zi��ӮĈ��bdCu���p<��*��K�vk���S)�塉��7LAƆ�o6���;�f�CU\�j��T!�e�=�Q�^4�E�)��:�����o����]oX�A�'Y��h���a����Iwl�ٜj�^J �v����Y�U�Z� ��:�Z�zް��G��5�_8��S�޳�X3�; �56 ��\F�&֔\aGǯnG�����u�R��엶+z�.��.�n�v��hT�)�v��AAFvjvnu�Uf���L���lK��sd�>Ǩ�[t��`�����GrC����-ep��[kZY/n�|��q��k��bkf��Y7~���`�>ǥ��5v�G��(��t��J<\YÖ��v�Z���/�����_>��B��X�cgϤ��3������'�.���x4���-�b.�c6���Gg%+t�ܱ}�^�WF��!�֨4S�{2&
U����s�i�V�.�$;�_��o��23���< ��)�3���bų��_��U+�R؋x��9Q\����u�v�1�.P�������;�IJ;�8_T���a�����W9)/�eB�=�j�Eq<�D33���]YKb%]mӳ�`��%a�L	�os,��=u�u����`����[WHg�s�u
ñoSH	jh�9���a���IL��]}��^�01��ު�	v�
�9�,���`ƍ�
W#��],.� v���Rh0��ō_>Ogt�g�:V̜�`�e�G 3�ܓlS��+�5�"�,��e;reM֯���Vi]P��˼��_v&��gOgK7�����9����Y8�E\��b��3�u՘�U��:�F�[�](��E,K4�m�c�:U��9G�wfSJ�eKY��:�N��M�mXڷ�3_(V6��]�1��νc������Nťg5A;7@��b�ݨ�Tԯ��G�7�:�C�ݔ�=��ڕ�õ)W]��{���6j=�֌�����t��6t]�yϲ$1��Eb��TX�1"?!W(UA`�AEE(*�XTA��(�PX
E���)RQ�(�*Ȱ����`�0�E,PPX��QFPR*�\�VEH���d[J �3,��`�����ed����U��Ŋ���*�Q\j,`�E&5dQX�,E&�Tb�
�X�1DET��UQTQE� ��AEQb���,PU�X��(�E(�UŋWV�*1�1TX*�V �EPcE1�0+UQ�b�*�QDH�eQDPDR*�H�UX �Q�熅M'��U�90�U��v��Z�p���s���j�u�PNۖn�k��l��n��7�z����Y���TLO�������'�}(�D�VZ&:��d��$T{ �2�%b�S%F����zޙ�h�#`o��2H
��x�S�ܜ�+�\u��	I(
:���K�}���Dz��Y�t��W>���eӁ���r�\ا}
����s7 �r����gF2n�����z�H�p��6zLq�y=d�̋\:��d,�:
��_e�8\���;Sa=��j<RҪ��D:�(MH�V@f��LW�f�q��*sc\��l'>Q3�q隵��k1'�b�,a��t*J�+)_��Aa����^��g/C�t�r�
��PK�k`DX��3��C�͗'�"P9I�-���$fb��[�,j�zQ�����Dv�@����1/.�5>�ts��^�\U{��5't��Ҩ7w\Ʊ)b�Hͣ�r?fݦc���b�����"�&�ǚ��S>�C�*��B6���J�#�wW�lyyt�t�����z����۴�;8ȧn���y���"U���&
DZ"����*5�d4�U��j����>-�������N��zA�������~�����s.��s�Zk|d��<���VۜY�mu#{� ��������gd����S�.�s<��˵���Ҝ�З�4�j�u��|Yјkx�
�������&����|0f�9=e��F̸�>�Ū���TS/�I�N��
67������w��n��W��Y��
*��:�/�F���Z)v]���y�|�d�(s}s7G�z��ő��j�_���s�g���:L�$H��u�T��>u�4�˵��d@�6aLv��/�����QcX�*�֡`uKK�	���18H$!:Ja4݄M\�z�P��Sՠ��+֦��9�q�|ĨW�t��s�h�S�U�؟�p�N�cB���ٹ"�"�Z4D�(��;�I��mʁ,֗I��|�IQ~�Ւl"&
��[٤Uo�S��_F,垅a�e�H*'�~*V�OB��,v��Y	��#Q���+�]&���=�M�w`ר�o�^@x��F���*�S���|Tr�<�����0��	3������.�:1�����`���#r�A1��fE��yL���v��aI=5��wu�O*1�u����T;�9"uMI���24Kf��;��H�ك=Q3Y���{JKv�B���ѐ����5��x`�Q^��F5����!�i��p�wYfǚN��9S����6�_;�Nm=�V�8uI+o.�v���s��h;�,��`�-p.���x���e�V�F�uko��UC��n�����؟�mFl>��p=l��#�
���Vx�oipoiX��Jx4�[���\�ݬ,Q�sv};��(z��1�l�T���Kֶ��=�bPx1B!^�۴�������z��=a�n+{Su����n���b��[[t������u�t��5xо�㯽��e���	A4�'�20G3�Hȥb�!М�q���S���A�dZ.�Ʒa��mf��D��Ϯ��ݵ{�Dt^����Dϸ9@�Q�NK�S>1�)�=�v6�^��4%���1�lvE@���?:W�~o��-j�G=�����	
$%�u=A/RN��{;UM��m�y^��v�V@���B��M�@r��9��v3������"�P�fz��X&7���r���V\�Eh��F�ɧF�M��`D��X�jǓ��[�Q��l*�-�����W7��/#
����*@4���P�b�}j��S��@��du��["�T�F������>I^ډ�O�Lh..J�����
=#o��w�t����Ï�m{�
E����2Z��F��j2�^U�e���Z��ƨ��Ul�H�/�q�t�B�@.�u�Ϣ��	Qw[�֒�S�UK�66�\�Qע+�P�vh�Ꮡ6��2��e�p���WN����������v�d�F��	��k���Ӏ��z�EG���++��2�D�"}�?@�K���[@J./�zX�4k.����. �U��mTtN�w����������"$ TO��#BL2���:jqP�U�r�ݘډcN�W6����z-����O���;<�h��p�����$0����j��X�=�����{���H�0+M�q}�;�P.�ģ�tK�L'T~�[�^	DԂw{ʔ#��ӥ ��dfs�6�����8C\�/���NX��bX�;3rZ^+]��ٯ��T���¬x]g�Ԍ������V+�*�}c��b�t�a�T�Jm�Ee�o��y]�<�0���XǍ7���,{қ��˾�.�z/`n�� �.��w��A���r`;y��x�OrxS��%e���/x�l
Dd8�&�_��hQU7�2�z*�y�]+[� �̫����|B�Z��Jj����u���D����9�>�xZ~��1��%8�vFOP����n\
v�b�}Cc��L��3�\j���;뫓&���HU���t%W��p�n��x�D��1���0�8v�F$�9g��Y�=��9j�TK�*������W_.^�z�x#�WWJZvht��d�®�_dZx�37f�79��q����v�*4#���K���";uB����)��C��f�2��F䃆t��sJ; �����2�:�;�dPs�ca�;�)8fo��G*�㞇���D����U�P(�
J��<=�|H^>���S����Q� �{3�$����ݟWؗ
;9�!:���=$!��t��Bb��&^3l�Q�mc��C[��.̈��۱#�n��;V �&xl���8�!��J��j�[c�7��[J�'u=u��s�� z:���&T(�>�.:�2�%b�S/�{F���\�Hu��ďW��w^��ӌ����S�w�IV��1A)"�
:�oψ�ۉ��Q��*$��*i���P��*#Z_-ʁs~�X�[��uY �rS����2	�:d���xT@U�C�a󦆕-z.�K<�\:jj�d,�AY�%�\3Ӽ�D�{I��[�ܲ_O��}���	�
 y[J&/�ӄ!O�Vy��(U�}�脹��W�y�h�d?B��b�RP�F�h�L�s0XuB����O���{}��wN��t ��]'uVe�h�e@Ǵ]��Ը���
%�E�᾵i��]�7Fi2
Ve-�X����,!�UƲ��*=٥K��w)�\z���Ddqq����9v���17��z�A(*bm�s�7 ���'�s�[��,MO���3���ފ����ݧ�kN��"#�Kj�('>�w
j���qRk��T�� 6[7�6(����g���+/X�[N�]�V��ƕ��7f��Z�'.Kˮ�W��M{�ܚ���u��`ȚQ��v��R�jrV� �#�Ty�m�㾎�!�ey
	��a�]�Qa�W������7A���L�o�n%��v+ӳ��cbM:�:������ȗ�w}��+�3��23�xNŊ�]�Ei�C�}~�e��e�N©ɧ
0��Fު�^>���ӯ���>��R��wl����ڦ�+�Ai"��A}�Ykf���
�q�4�*�(kRn�V{�O�e�Kv�ň9ӈ�{L����>��2D�l�L�"��S��N�N�i�b�����O���b}�-m�<�Z^c�%L'[J����3�ה���z���z
�e@ޕ��=G�C�1*�D�gb���$�v!�L��ʜY�G.\���
:�Ypws���*�7�� ��9Β���Ւ^�R���Z2,|�a+��#��!\,tk���1�7-�-̖^2m��1r9]��-�ˎ�轕o���̠�O
��M�+^p
g��&ms����y1�
e��ػs��c��\̹�)��;݃�[M�;a�n黸�O*c<Hն��t:}ݮ��﮳�F���D�l
+c��GX�BF����E��ͥb$ː��Mtf�Ln�䘴�!LG���I�r�T�+%G��O2��e4�\�]J]O�[�J/6X�U	}`u�7X Җ]^Tv�
 a����P�"^�B�o�܈�j�y>���Eh{3ЏC��:q@�T;� DO�MI�
�1(��T1��ls��O#mZ��,7������]N1��z٩�G� ��/�������%�}�d��������ur8(�ݟN��a@�U�f1���|<)z�жg�LI_Qx�'6�НNq�|�"�h�������^z�#hv��уz݁[��5ζ���ug>�l���l]<�w%�C��T�#+>�Q8f�$dR�U��	̷��)��mW��U�D: /0�������W%J,5n����3,�&G#+��Q�9.-g��1")�=6�-���
G'��w0�o��@����ҽ�o��-V#(�q<(\��� d��i�r��}JQ��Q�H<�[^� �5 <�Ǧv�6���L�S<�%��CJq�v�*����)�*��<s�ɭ�|h���p��gt2�:zCڌ�,q̴'m�ownOL:���KuP�`�͍	�T��s�����(�����ʘ�W��;�v�yJ<9�t�@�Chi�M�&� Xt�Ź��v3�����Si֔�كVݹ��̄���p}�1�FC��vM:7�m�8�ek)w���9��9��t�ST_'1�jΓj��>�p^��Q@J�]HR��[.LW���tp58���
�\��f 
���,�ͨv"k9�:�ac%VĬ>�=�A��3���o��w�t���ϊ��6�e��8�o'inX\_�����(Rg�L"'�\	%�J�l9QQ�t�B���ڀP7��j!Ў�<��F�95v룓��EA�(�w�F�&QRD���k���ٝ���}q��R5�z�E��z9�ԅV��u�yy���* BA�z`�wY[�[������`3�|�⦯��3����7�%��y;�C�@���5��j'l�u�/Cj��R��,�TҬ�&��V&֫�����q��/y;�4�#`l�&s���}3[1����駴�0�U��k�zSP[�~>��ł�ܪ�90�Ʌ�r������؋k��F�H���Z���_�����Z7�_��8�PS��b��������a�J��6��\;���T��<��3Ji�\�0���.37�{�!�O��SJB)dt�hU���K%V��e�:��M�ï�����j�9wӻ�[ҷ2oN�+���<|N�2'�	
'ё���{"F�t�c=�كhO-Ad�u���X=���'k{[ PmT����y���)N�>�-���)X���	ܞ�D�2�j�T���^a�W0{GO�f�2�r6;Ϥ,5a�f���D�#t�o_=R&�Ok�-�N�\��OQ1��2�8�j��6\	|�l[}Cc��H�f�A����!CΊn�9�w�E��9%Mq'!��ӎ�!H߶f�y���܄�f��F�z�u��Ǽ"�ڔ:��	t�lM�*�3r8Iq�N�V�@��
^�;p���$R;�V���z�J{�u�ǟ���g��*�1 P��[�T�&�t�v:�&^��f�(r�c�Rz	4w�;��5z^�4ۼ�l������L!0ID�\���N]�� �^S���6=}n�8)ן�P��c�vL�EEI"����(BT�QR�lݸ��ܗk��-/�s萭ZgN2*,S��u���A:�z||6���]G�� ��/��*��\�-�uwTd7/9�Ǹ�)B�����Eƥ��u&���=^vL���Z��6��@�Q�~k�Kt%;��l�x����j@�NQ۽�뫈�Lt��y�����-���ݔ�^mD/���]�PK�`��&n��tq�7D�|3�]1�˯7_YL�b^�/���䇏�Ji�t�Τ�υL�4��O.�飥/<���y�Td�
.����[�l��]v�t�F��c�>�<�T���̎p��S̅��g�8�jѴ"v�%ћ�e�zpA�)�L"��TԌ�`�m(��_k�B�1]#TlE�FR�Os[��+�}!�Ы�����D����DĲ	����Ϸf&(65�L�r�5S[ɫ����J��H�b%�S����)�3{.*Mpr*��$6[8ᥢrL���6鳷��d?i�F�l�[�%�z)�s�	{�yG���iߐ�&�l�Ri;���F=X=�n�`,kY�S%3GC�ey
	��~dWd�[ܠbI�&d[]�O+2�u���ϕg���$.�X�b��v����)�W늤�U���E;w}n�M`��$V	5ښ誛�զ�N+j?]�R��}5�����(���g'��\�-�YKA�W��l���
V`�o+�<�wK��E���"C��#BH�n��@W�*��t�/_���Օu���{Ùv�2q�4��{��ʰ@7�4�Il�*����D�6�:	�+3w��k;7�'�9��Z�梜̱��B��(x��)՞G_�L�hT��.�A���&�`%��A>����V��x�R�*A�KE\��Yn��W}Z��{w���Ьfvtz�R�cV1f�+��zRx,��ǽ��ğ*W��>9�ϊ�J�gR�����2���[����D��ܗrv���Ȝ�Y��J&���nZ�1Y V�ǇN�����n=�\<U*T���J@��C�C�7ʯ���!Hr��sWfQ����}[�@�D̒�"ԘW�6ũ��'p8㛛6̻��r6v���l�A��e�v��N{}`PX@��R�)`��� =�C�j��:M��U��]i��_�;��w����U����)���/guz�;����'	�:��h0��ow�v&X��ڵ��YF����89*��{96���S��4Ib���zXvXǲp�4�w ��<�=w�@w�$=���Ҟ�A�h��"7����N롘|'����z��W����rP��ү���9-n<he2y�]X�c�e`:L�M1��qW,w�[���y)�'�η̌*�z�ǷZӮ��V�����o���TDk��a㦱�׫���l��Z�.��{�J}R�D]�d�3+��V4�1[5�{��[!�9}�<�`ݾ(���Eh�[�Y��:ا��r\�7.<�{-g�+'Ur��6S�3�wSV;�2���-P��q��V7��+�RԻ3�5��5Sݩw}���*��L��9�^Ѕ�*յ+k��69����7g:0��W9�+t�x0ؒ�qJʛ	���7��.�}�!��b�YG�dԺjm�;;NC۩{�o1��5��cZh}7n���xCx�<�G���:����b�[i��������󦸧���d5)�3yR�,��16@`?[\"/xL��اZ�9G��ӡ��%�Y�L����6��+u JX�����d㫳.�V�P��Up�*]�2`�:��i��@�=�U��Nu�v̥v���x�i�k%�l[���l�w|��4پ=���]��A�t��4��d�����v�P�o̮���]5�ʻy3's;)W\��P���O+)�Aŏ���9�V[9Ü��ILtL��hѱ���-�*!�Ѹ��i�Ƃ�/�k�3o��*V�.�Х%��×��!҃ׄ��-fV䥥R��cu��TE�Po�0�p3����w@����﫠�.}/.��u�ӱ�-@�m����5���
���R
��umK�P�e	�.��&�կu+�ʷZ)V�`��/U�\��k�k�񭗆A���I�� n����^@'e�{�N�*pS��Օm�o�
]��٩Ջiᖗl����ih��5:�YxK���Ϯ9� P�P W��H��*�"�����1��UQ�����QR"�AUE#@QET`��AX*EV0b�5X���E��

�U�ł����QX(�X��� "�UH�[b�*娣#"*��UAUE�(0U�DQ�ʔEHŊDQ��b��-lU�UDQEDF� ���L�R*
��PDX#""�*+��J�V��V+TTDJ���*��J*
"��U+b"�ڢ�A������U���\��\r
*��J�U���T�"�Em�UiiDQQX(��b�*)eT���b�\Cr�*��b2�"�U+AX6�X1��Xւ��[JT��X�kYmj�61e�Q��`�\�Z�YXR�T�JH���4eQ���kJ�&A\�Z�ѢũU"DE�(���y��~�z�ߌ�n������;A��Q��n�E�壝nb�/u[/�ǎ���*�gt|'5����d�75��N��Β�6%n��Kx��ϹX�n1��8�9ӈ��3��g�X*�*^�)��	�/33]ta=��uWЯy�O��Mm�6ܽFn���>X��$R����Sd��>����Eu�r�
p�3�_�GE:�"}x� ����=G=�q���!��Z8T��[f�����[���os����@������6}��:sz]`�J��|��3�=Dp���4'NG{����; ���8�G��p	�l�\(�OWB�V�섍��na��'�����jŻaia��
�]䘴�!LG�ø�Dg�Jh
.���}��R�n�%�O���w�h�Íu8x�(������4�"'�9G	P$�ӊ�P�FV��*pV�+�������xW��ã��8�JP� Dg�MI�
��<��bB����u�ňK�`���+}�-�����p&Xnna2��D���|f���Lm�D.�a�%b�]���68y?<�Baʼ��w~��Γ��5�����2�X�L���7f�K4��&?F8��4^��Y�}֜���7�M���ڮ ��ۗ����U��h5�L��Bi¹y�r�s4CCւ�O�bl�HqT�B����v���ޙ5 8��n�Y)0�Σ�2�YI���|�[�p����ޤ�;����qY���c/���*�>��<*rq�&�tv��ћ���cv��~�[٧������w�L����$����W^aYOU3�K�]x������Ws�o!N��-��l��o�@޹��-�J�Y��t^���(����FU�	�M���ai,\;�~l�W��O2��zt#�ή��^v+�O�lr��2������!C��ϸÛƓ�p���DQ\]K�ݦ\���M
nsɺ��S�s#��`䫤�=����y�&�:�-��h�c����Bt:�iQ��m�8�ek)pNÅn�F3��M���X�Ω�5T���P����\+�H�A�l�Q1r�����^)���Wb]��)�:�K����S��yy�^��~�2���W�1�p��;g��x��2]���iή�{o�xE(�~}a�h�{�X1H�2��0��;���n�.;�M������ %�R��	�0{��[���|\�z6w�p>"l��*�@���)L2��6�*������K��l��C�����N�V�ЬY��=���;�{kM�,�]i�hJ]���*�o�mp�M���]�����ř�ݬ�t��N�f�ݤ�tU�2�xʆ�7\Z�=���}GuL%�V�<����BY���y�t��VR�����mz�J�jB���������D� >@�;m�7}����pxl7�'�|�'�H2��F8ޟM�ݤ�R`V�P\V�^�Q�
���2����re�͈��f�Z;�8���Q�4�+U�Ƈ����JS�U�z���8�rh������ݹ�O���c=H����]Xtr����>��`+<�M�Q�\LP��X+*�F�y�L�`�e�yյ�L`~}J&(6��3�S
���Uc4��J�/�X��F�W�..�A�⣔;�<�'���ۦ��C��l ҙ����ؼj��ՅBɟ�6%�^��)H|��LT�EK�wI�p�����t�`������ʸX��/}2�5穌�50��{�P�3����s��\��'(ׄ��q��BX�!�v��;�ذ�P��^�L��D�@�gpjǾt�-� �SX��J�lq�xn]C�ϲf�iϥ���7Kn��n�D��ˆ�Z=��B��C�í����OJ��B�eӄɉe���\q[95���N>��WQ����v"!���iw7qXn�<�r�m�,��s�H���Ⱥ��:VrK%*�wӹ�3yb8���C���*bsa8oz���ϝ��J(3�C�|��2��w&.�;�o���錥���Lj��Wm4{��ym�ʤS�5B��q��ׂ�p�z�
�H����=$!����v:ͷ3��X�0�/W-�F�i�\DR41�P��n��Ga@�s��q�(C�CeX�;qs�I���ۉ��\�*܎��R�>)�� D�P�]�7ǃF��>>��X��7�lLZ�����J2�v�
�H�>��W��N2*%��:V�ܜ�+�\u����I����6G5�8��z�8�O�a�u5��)лU(�S|Z4ʁR��B�.�����7	XW1�ٷ��GOH/��'�J�>SH�k*�c��QXK<Ȱ�u\�<�u_9}�D}G��,����yڨǫ"ˆp8 �
} ��t:Pd�����x� �秇��:xL@q�s9��=���-옮6܅К����:&�@���LK!Qp\�C��%�x�ɣ�4��Ϙ�ڴo\�-�Cjf?A��§ؼ/kʛ�����v���gN/�^t2�����C��$�v����n���A��Źpb@yu�*گi49��C�P����7��=K7�1C��fr�r3�ʞ�7�`C�2�G�1Bmg�?\��炍�s�y� ��t��2�%o�w�;kܬ�D	ԚH��kD=��Oni�N���ɋ�&�].9�cn��Uۊ�[�`|�[��dwo�\�d�hGZ�7�f�_5�;o�����}�����6�6��|5���>ͻl���>���-.��E���s5�
d�F�k��x����X��b����ڞ�\���<6�_�x["[���n}���TN��u�G�̮�Ӿ��i8��x���+�V����ᰏO�l���4�hQ�F7�sn�(6�����S�g"��:�����d�`Hs�\#RD�v(�@UyǢ��)4�ձ��Vo\0��@x��w��c8�p#:m
g��N��"D�c�+lMgN_jb�i�\�p�k�wa�GFt�r�#7E�b|�c�P�:���1ђ��N�Ӝb&`�\)�u�
漽,�(ک�܃��P+��H�F�s�X�H�X�ѻL5wR^�M��'������u2���fzT��l��m�P.�ޗI�QFh������LEb{Ϣ��VIP���8�G���\S>��p���z�`��=�Iɉ��S]�'��T��Rv&��-��]8���J����H���ME���ϳ�y�XZbx�*�=��n�Lz�n��#MA���ڵa��n�11F�4����T#�Y%[������ޱ�A:*]Z��cͣa�R��G�Ρܑb�҆�}�K��Qޗ�=ce��v�j�k����_F�*�����".քQ�te�:N����d�˝8x�(�__���GA|%@��8�m�qwٗ��u������z;�h�(
+�U���`N�Q(EC�@���jOPF���l)�ˋ{�}}Eɤz�1�@�J��mfl.���H{g�����������0�ǁ�Xt�uS�9>:D���ҭFb��v�5��a@�UM�C�Xb8����n�lf�K.�=��k3��<���8�''y꜍�۫F�w��bc�Y�mr[F2�jl+牮�1��O��F�N@�=��5}B�ϔdO��F�>Jǳ�w<0�2��˼s׈��V�j��o�A�dZ)��A�w�F�e��*�������+^���p�1�ܚ�⛚��'��K�)�pt�?:W�a>Wе��2�<M���>����oF�MsP������V�t��8�1ޚ��M�@�*qa̎��N�;�����՝�c�<��N��/PT&aO�K^��ʣ�T�.�K*����8^�7���/q�P�ΤF�EnDu'�� ��*5���&�"��wL��B0����n౨mc䋽�x��c^��Nܢ��J��X R�W[�3�'(��i�e�gݚ��ܩ�� wq�n�,�g;��Y�R����]/�h-.mdw}�>�om!�y��9���k���%¿T�H�.Lw��6s�N2�A��D(�����v�0
����:�.r%���q��Ĕ#jeC$(��o��3(܇��������z������A#�Gc�^��PEQ�~��D��p>��)�y�K̼ݙ���ԧ�Oz�4z�28����CF��S���'ہ���W�PDJD��)����	��1��w����Ğ�$J'vEf�����=�QT��C�K���n�A��	&a�+���ȩK�w�Ax'!T�3��B5�ӠF�6s�T��ƨ�؝��
�pǫk:���w&{�k��j�d}.�!lu�ٯU�[��)��U*:����NL0h:4�}�1B���1�,F�� �X�J*(@�P`<+>jf�|��ҝ^�C���=�W��bf���kc/Hod�
҉��hVѶ��́��26��\Q�FFCw�dl$�r�u����=X�yu��>�gE�߷i�v�l^iT�<���ƪ��)N��fĶk'�A�M��j��p[�[�:�[��Z�V;��3�5�7X1�4a���m�m����
gĪ,y�rή�ְT�.��&�ܮ�'���a7һTh������ۑV()��j�=0�d�8���yo�K����3,�1w@����O�.lII���zS��Yʱ@VǤl87n�}2�:�����pu��h~�]e����P�cE�U[�S��RO"q%��К�>&�d����q��BX�!�l����6,7�6:5P�ǽf�]A��顤�
P+)hǈ?*k񨍎0����q�fi��N�N��q۹lgmJgTEf�vXtC�����iWD����g"�
�;(Er�Wd�
/f��v�tuÅ8�;�9��O�\��h�}mۏS9��3�Z���>�Al��U�b{�@�������6:ж���0���_A�R.")�(u���dv�z�xi�8$�Vh'qT沶-*�:��C�����*܎��U����_��F���K��g¬"����g��z!��˾����)F�v��\hK�F�W#�t�"��O���[�u'ZJ�F`�͔�^�z�����wE�MV�!�����d�=�kInE`U(�o�GE�룙��ʱߢ����u^��ޗ�03j�AL�5	PeL@Q"=����2䨻%�d_�����3%]p�]V�<5!}�bT�j�=��"�:x&/n*��ސ-є�,��+p�16�EI��qsʋ�NS���7�Ȳ�0n��Z�7�wj��<iSx��ݺ�����8l�Y��O9�.�"%v�֯x=�׍u���6�7�{7s(�p_�L]RI��l����#~���.�\��AO���#C�Ԍ� <��\�E��}�62��i�w)_C�:�ߵɊF�rCBj���C�
�^��tN#Ri���_5�ڒ���K<�2+g{�7/����R�h�T�
DC>mT�y9�C�SVf��E�yS��9�=���={��@`�����	�fm�`Ң��a�S]A�r��ʞ�X�i=�0�����9�<yr�̒����u���wے�m�ݶc���b{���y:Zu����y��cV���U�P�3r���:}�%Fa�\h���8�6�׃:�����<�.M��&��bK���쳻kS�"����ST�4�"􉫜�#���\Z��}m`�?�d����3��6�a7�|[�QL���Qyװ1��3�>�Ⱦ�078н]�`DFN���e�.R��n���c���y�|ݍv�x/�Y��.
��$u��wN�'�(]qѻ|�g���"�}�;&��i��f�(�b|�}jT����.V�;�-#�����Ag^1+۹��#gki�z��r�}uJ�ʶ� ��|D#\�����M*Q��r�"*�y9@��_�y-usvJ�-����mX�%ǹ�{�o~��=MB3�2��1�{�W�Q8�u��b���:z��\uY|�NT6ģ�~5�4kk�*�΋�ÅM+������P��H�۝q�5`)_E��K>���a��v$�p�L���,ϧ�A��l�)�@t������CF��u��x��֗b�С��D��]Y&�"`�����T|+�_b>ïG�������>�[0��y�xj�P��#Q���c]�I���b=ބ�ɍr�T�
:�e\�}�Яv�=�<�=����O2��Ӈ�tY
*����7X ҟC�ƌ�\+:�64�Y�A˷���T!��bF��g=
���f���x2z��<���)g���z{n�{�8"Ěg`X�f�}�-].-��Zۛ��'(i{Yˎ �R%+v�w�`�^�_�R��m+�u���C7k�C1�P&�]�c>���D9��5%w.�霔�]qpd�-�^�1(81J���hxg�����ݺ�t`���hh`�vc(V���{b5�����X����of��t�8'�2$`-�FE+Y�1,I��j�E%���=Ɲ�.���ڠ��.�WB�m��I��wTU�k�|Q#v�u]�;z�lI�R�ʝ�N��������u�;_e�r��R��69Q�Kc�Ya� �o���]��y6����0��(�%J�-c�TG*^���<���!0�4�V;��e%+6�KW+Q����n�sw���+��F`ʉa -����r9Ņ�p�y�&��kt���6��0X5-�^Ν�Q<*Z̭{ل�=ݦ�A�%J<��%�`�ީ�a�Zk�컆�A3��T���0ɑw�|������i��³[�΅,Wbk��v�Zȳ�fr�-Y��R�L\y�U�z�\�lj#oJ�����Y�7W*�he:�m��5�%�z2�s״��AP�%)��]_z�v}��\1�j�xK�֧�)em�oq�7A�X�đJZO�����%��L��yV�י�wF�+����|��R���ضg��YK��v#һ#}o���rQ�vM�=�˵�
/��\�Mr�ƕ����ڜ���W��C��C�W�#�>G_Z�7l�mJ����!�.��ގ�>�[��w-f<ShU�n�;J�c���p��*Kk6��0���!�d}��_6�1��1�zP������Oedz�]aM�1�gڱ�"Z�K��mN*�A�2K��3���+��$4����bRM껻���oM@�Y��hR��]S.�Sh�ǟc�+�ښk�m��X9�Z[)�f�^ru�X��.�q�q��o�*_J�i�ɥ^C4�:NՉj�7.���5���ڔ��ݾ�5e�V	��4����}7-]t���NY[ ��"��Dm�Yn�4ݫ:��ACZ)��o��2WX4qR �:g��=V���Iز�>�J�<���Rws%ӻ���]�j1czMmgL�Bn�Z�JgR�:Ł���ۨX4�Cuc��7��J�˅��嚶a':�yu�j�!���𬺶��j�]�PVj��:t�y7ܕ�ɍ�;�uf��p�ˮ;�Su�hb��LM#��Oz�vn�1\�J�x��27W�&ke��*N#��J����;{��0�9M�2��Mo)��������e_Vm�V5��=EL6�1 O���������9�*��wS�U���t��y��yi�÷�2l�8w%�tO�_3���\@�(���F�Ŏ��x�f�tm��>�3�^R�eԮ��PR�G�{�R*��{ŗ��!�#Ԗ����:빰��i�k�u�dWr��|��Ҍ,j�ݫ������J��'s�\k���@�å:�xՖ/n��>w�9*��!��^:�����[o.u��б�8tt��0<)FB��2�epx�lv#�zt��9l��u�`(�e"���52)�r�O�5��8����͘)���zi@.Zy��8^$�fƸgM�n������Ϻ>�� ¨T)D�A�Ekm�X��/�Q�QQm��j*ڢ��jT�m�F1Em`�6�[j*2���Qe�*�[DA�X�J��
T��Q��I\amV*"�dEJ�(��ZR������iq�1��,YKR��$m-�X�Fҥh�������1�*���)�V�Ѳ֢(�J�6�b�#���%h�������ƉU`�+d�mK[X���TTJ#�TGڰ��
*��e�E[h�*JإlF�,�V�"�b��1E(�TV,b���V��U��eB��"V��H��Y+Z#�UԲ����*R�V"	s(�X�h֠�YUETDV!D��ڊ�����֋K[B��-�4�%���P��V�c��"���V҉�WZѣV$o��J�Se��cy����,(Gi��X\���:���=�GL���8��G����:����9b�-����,��t�ZU]�|!N.�<��GT��j���t^��E<��'��s;�
��%;<������|a��ODaA�5��^nUd'�[�ݪ���S�5���*�����g7��SHQ0�f�OPw��4��CkM
nsɺ�*p�g#C�ېze��P�M�&߼���CI�}P��
�&�F�p,���Bъ��B�wor;�����^6�]��`uR��4���\�N���v5T��3�+�֭����e��3�G5;E7 WV;D���lۗY�'�GLh=$��_�MC�2{2��[���z�Wv�=�:�_�7�V���f���W���
�Z"aއ�b�x�u�.��R�_t5��s�"���T8��5`���j��w�p<"���*�1yqUU�Y:*ާ �Ɇ\P�'�xNu��(��OCど
.�\t2�;Cu�i|0�{3Q:1.��N�BO�� �e-H��8��0���~��E<38/	�ޟ1��V$.��		g�X'f�{�Vqm'lbp���{M%\����F�����gV�d���vݎ�G:n��+��+\GC����t�m"���(��gv*����QH�+2��#e6[��u\E����S9�,�Y������k����^2��]�E�fQ>�L!�
��x�+U�Ƈ���Y�i����^��r#v�:�d@qyY2o}u%��d�8�}��O	Q1뎱u�;��6�xz��y�z��=��5˛9ʐ���h��&nTL'�r�~S
��E}�x�{J�U��Ӥ���=ebm�og���9�W�Þ�4���ƻհ4�b�y{{�j��ґD��}5n%��{��f,#��kyW�t�.;26&n������3�sP�:�VkC��3�	t��Ut�X����N�8�M@��!�����َ8J㽪C��\
v�l8�f��Z�"�D���δh�՜�	N+h�e��>Tp�"�74�B7�4����dN���_#�ϗm߫���E9α��mWD��נ��6�^b���
�5Äy�gz·��Qʉż�;r�1<U�X�j����s�#�L��t�>�-��R,aQ���[�w���,_��me����V�c��w��A�JypZo%���x�^�y���AU���|���__�
g�/�����&)�tn�
;��vtĺ�@G�n�
G�Nh�/.��v��͓�^��I왪gб�q�3K
�듛��b��ز��M��q�wm��V�w��Q5�Fr��.an)԰����"k[����ܡ�WJ���LJ�e�no��a�{��],׾�ꐩq���<n	���2Q�mur)t�"��{^�7���w���5%�}�ԛNA��m�v��P�n�Au
�WI=��[�Y�R�~�7ţ�ܨ4��!�Wf��v5�rz0��?5U��9J�ϔ� k*Lq�*+�,�"�3!]֊ۻ�ںy{mW���X)�VlK�gs�
>�}0�3��TԌ�d�j�m�{�I�*�mG9D���g�T�ƹ1H�B�|&��pA�rf��5�|D�R�r����gg���5�η65;w���3��c�B�45�9�3E�u�{=Z�W�}�Ü�7���Ff-�n�Scv�浊m�+�lu�^ŝ=�F�Ĭ��g��h��2��%�k��2�����lK��5X.���I�������yV�zf���0|���R�NL��y~�A�*���E�9�j�r�����l�ޱ/Q��8+U�lfT�Jqx��nM���<�D�
�qr�
�΁��Xe���j�_f�3;�"iV#W��J6�-mN9i,=�g]��;�m����!#�&txtZ��M=���=�e�]v�|�<=���b3�~t��Q~�po�F��G|;+u�^n�n>�3B���F	Rq�8��b�y
Qvf�ڊ�;�ͦ#�-�-��L:N��f�Zv�8Hy<%8޹<$_oMQ��i���Ew1%��jƙm�n��v'^g;�ë"��C�:��Բ��k�)��K!!�=:>T;%M�I��jƱK$��g�۹�LT�p\Ҽ�GA7$�P RQ>�ԺuSK��W3z&j�S�n�l��t�f�V�
ʠ#�ϡ�&\r����-�������Z3��ue�C��ҥ�J�9�*�� ��P��.�ҩ���@�z$�Q]"&Eh�Iͮ�7����J�=T�Z�����% �j�4u�m"�'g�����~�׵@"���s\Ү���/��7�'��(8Fq���´�R����Vw��n@]�k�ku>�V�;�50�o�_�Y?<�M
�P $q���ҩű��s�k��Z�hc�K������q����5��eb<��KR�\�1i�E�G����3�ow��8��uړu�u
ܹ{{u�"��~<뗔�-�+�k4l��i�Sy��N�2����b��+Ӷ�-M�IM���p'�� ]�k��M�.v�K�nH����"r�v�$���E�����৆,2�̼�5��M�U6'���%�����ޙ��#!挚�U���3�g�(�of�F�-��xbb�J�+R��f�'�USx:��SKi�vU��3@uA��qw(p7�I.���E��z�:������g ����̥i�}*��a���8<�8��"�����{JT�w�.rd�C�1��nުv���|�B�@������^��zvw�s�vNKV�U�-\k�e��}����F&׮�b�y����A��7 7`�)�vJ��*m��-^^��U�Z�q�K�{�T���W���p��Y��>�J�D����$����熣B86c���R�m��WcQ�V�2���݉N��t_f{����{��h"��<��}7k�S}��ڟt6���A��Y�Ӹ�+:��]>;8�4���U��!���h{�mi�����������7��y����(�r�ɝ�}׽-^a�Xۡ ���} ��	�>��M�������d�4�s��1ر��6�]#ͮ�v��w�U��w�CY���^��*���]1��dʙ|]���*/}���<{���}�l
}��se�#�4#���Ŝ�Ɂ������gdU@F�V�ϯ�%ut��//�ON�!�!oC�7����k�P�>����8�*��[]S}~�=���G˼��~s��4!�!�<I��~������[�,����e���Ww�h��1��ܔз��D�>�ŀ��bo7+�Q���G8&�vK�}:��p�h�|2h5Xhk����.*�_.G^��qj��s���6�vb�u۝��Pi��MN�N�7�]cIi���z��p퓙J�8�ݼ��lws�e+Muy�,�FtR��^��<]�p��~
����z��H��M��aA�L:����][핾�wz�n�Nuk7P���d�Ts�&�w�{�k��#F�36,>cgS����g�-ֵ�����
T�S;�{"�|���&�f�Σp=5-dQg#�[m�*̢oD���ߺ۩8��»;���lݖk�IW�˖X㊷9Μ��)����4/ ����y8��������I�LN�L�|������M�u涸���Hy<%��&�.�&o/�d�=�k�<HVm1�y<e�X�I��:ҍét�lp�3e��6�X���{�cq��w���薖�J��uջg������6�5}{����V�,��y`����4�N�9��ޥo��0�{Z���sE��ElM�q^�ܰ�U�p[�s��T&\��'o�-��^�)�7�0�B�ũ�0����}	�+49@!Gyt��W�vG�uZ{��Wϭ�>喭�9
ś%�.{��O|<�-�A8(�pJ|֨	k���=��^K�T�ZNi.cxuu�|�e5T�:��pPt5 �❋엑�$�>���{�9g���+H*v5Į���
w�k'��=��cj�Nm��>��+�<(��o��ke1 7T&aǧa�j�@v*���ħPò�=:j;��dֲ��Ey��QŊ����g&�7;1/8u��n�\BT�`�D����|�q��-��G�9i����&����	oU��}&���Ao�>���Ԩ���η:�=p���{
l���«�(�9GR˞��`�Jy��z����$���v�v[�kd�k\��S��?�*��'�����Ḁbm��-��M��a�98U�)n���Z��:�מ�e=�3�Pp,��d�rdo	!9�쳛QV���<��������kr���ypy#�8��(�UeB��d�aNiM9|���������z�ۤ�μ����̓!��i^�9�N���p;Y�Yc�[��-X�-���ݷ)���H����X�cf�,�w�������:��rf���XއP�Y�ٚy�S�ϫ"�D�i>��c����r}҅%���Ӫ����u�
�f��n��\�l*�ՈVUF�}%Ļ�H��э�Z��Do^��%�V����嗵]n����9.[.8�nu�;�'5���wԊ�O-�g�-F׬��Ǧ*�����C���N36��sL�}Bڳ5���68A:�����	k��eZ���xΠ�9v9�-�+��B��_ ����um��z���Q��v�:���V�&�wmO;T1���RW����K=3����\�t�|��g�:75�U���R�ꠞ��6F��y!,E�-���$���<܂��B"�j���~\9�敬�Q}}~o'�Ѡ����F�\��t���C5���}�m�]~MH��>=�g ��ג=x"���r�p��s��X��]�{:���;w�q/�fB���ÛwS;֟.�7\-4X��F�P^<RԻ���ӖG��v�	)r�|�+t7�l�4d�6s�]�Rs�&�i��PjK�t:���g�_N�����lkKh=�ʷ��huA��{�w9�d�.�)ڰ�o��8���ͻ�a��a�̥i����k��<.�������&D����9���ua��|qfP��_�[cU7a�n��OV��sRn�+Q]=>�˨�:��7��)VZ�*he�D��_W�hиw�������Q#��	`/3�w�s�z��5s+�d���_V�*+�=��i��G�
닋Ւ��u�pq�v]�*��e��г�kM��oX��)��'���A�*swyh��zWwMi���G_��c���Z��v4�{���;���+}�)��I�����e�=;٭-<�bF�܃�M>U��SX��+8^E"�	�CF���5����jÕ���a�Ѳ7$P��є!gwm8ܽɺ�E�f�ąwKuj����uj:�jݲ𻍃�GH(.XGK.r.!��4�f�Z�)��������p��	�]��c�:����m���5����J;� �����n��{������9�}����+ec�YeF�#MB�Yq\J��m�Gr�L�b��|�p��J�_:nX\eN��g8Em�o�5^X�P8t=�ky#�ޝn��������r/\]Y�[ܨ���Ρ�D;>�'������b!�k.��]��1enm���m3|�4l�|%����hc�v"F�3�
g�1Ax��;�-vvjy(#'�6����������Z�	��X%}�S���h+��y�]@�4��lC�'<z*�AI�={6A�yM��;�컏F�_b4��P]�;�]�Tl�K� ����iZl՗Z�9��h�ugf�V�c�徹��՚�Ί���{ܖu
VP�[�;D��t�YV31�n�G�s��Y<����内��ˀ�i�P�E�\q��<���o�}i�V�I�F�y
-f+٫�B6E�YAt�龠si+�����$����B��s�8�!.�Փ;�fu�[���7���y���Z�lC�s�u�jQ�R�(;$����m|�_Z�B�����n�6�ֹf.���d�2���fI[��Z�m�Ҿ�[نe#�	˾���ŗ��5S��*Wi�8!Tz��*�iڀZ�A�i��ώ^��2\i��$��%�D"��z�+�-�Ɜ*��PԆ.웑4f/t2H��`㊂�ԱՃ���;�~��Ϭ�aEZ�kh�IX�kI�C_N!^�BJ즗e�2�k���8�4!�f�O�Sc���	�	X4�'�'.7V�w>Uܷ$e�Q����������(��:�w�ӻ�xRg�g7%{DU�}M�"�uƔ����بx��Ow�8�n-l��C:��7��F���-.�p	즕8�.Z�IV����Z���C�����?�';#��q�����6!��l�P�JYX�"�v��R�V����SN�݁j��^ٗwi,F5O�K�n���j t͜��T�(��g$1^�g�+�\�v;����P}w�����i�M����O0��:�ƮM;ʦuch]K����������
S����um^���1���^ň&:�y��vj�g��E��kA���b��7�5x������E��f)�@W˅B�\��*a�p.�Gu�4�L�QKG��$��lǹ&h�H�uNu���՜%�v��р�o����p[���ٺd��)X�RP��������)^d}4!�J0��cf�qڸ��>C�٧1ej7\�s�.�E��*�qy,)'kcr�B�x>w�\= TkM&F	�)���8�eS��B�u5S2�+�2ɠ�U���T�=�:�������ܽ�(�k���I�2br��I�����-�y��]|ht�hZxBt������i��`����g!Rk��	���: �P�=u,:ڷ���][[Y���I�(a�ړ���9/
��e��FU��]�5�na���P�sr�[�]Cm�����:Ȉ=˵j�ʸ�]���Sc�ĭ�o�1�l�7_Rև]���b���r@�̪쥎�>�S.cY��v��$�]��Ĳh�Sm�*�MS%�>�5�����c5��ָo1�X��0����6��u��Z,�r�rd�Y�L���҆p��eE����8�9�S�u�P��ͭ���A����1W:CRv)u$He�foP4@�5w���e�"�ڙok���xV��UVB�![R�VFYF1m)Phڡmm����֫YV)Z5[iKmKiU������Ҫ���m�U�R�**�j
�+*F�֭H��akT�˖
��E����(�ڵm�+
-lkIFm�(��E����@��b5"%T���bQZŭ�j��b,aD�VF����ƌm%K�fJ�d�*T�G39J���Q�ZR*�)Kb����j�DK#l�-AaF,��
�`�l���*�ę�J��eb��eH�T�X�Z�X�Ī�U�*ր�V�����dK�	QQ�4���Z%D`�E#K!m��B�T�¤Z�AIU�q�-B��*��ib�,TH����H��F�,!QeJ*�Qj��1�(�b�md�aY(�m��h�QH��H�Y�QT�R��U*�B+[
�*#
��E�iX�b��������
�o>��S%r3���N<+o�$u��'�^k�Ǳ��7|�JP'ehwzUr��
޸}8��A�w�-�:�':M�.3i�V^,��H֥��3:����Kh�|2i��C\�C���ZrL��M��w�k����ZN�7��������{�1M"�v� j�ɹK�Lt�<-l<(�{��MC��"�)�̥~�r�Y~����a���V��ȴ(ޝ���[�=���3oL׺��y#��+�&�xP{a����&rペ��p��~�0�x�E٭���x<���bqI�}1$�l�峐���ɡ�{�±4�8Ϋ�j��N�����c6���\�B��̫�ܩ�Y����u��ڕ:�l��-�4�w�R�Ӡ�v,����dnu^\�ɤ֑A�����w,�h�(X�o�ﯩ7�i��)P����ջ��:���u3��w缰L<��,ID���]]J�_�	W���W�7jLO6.�Z)�c�ѼXޒ�^�t�XJ�2�mw$���?n�-	ǳ{[>낹�Cs*l����h�>��𩦦k�u]�tgi�2V-=Q�#�ӭ�7�����N����K�f涙�o���Y�hy�NN�4;�[�T��q�ꊷ���}Ŭ�y�Bqu�<��+�',�zh�Kz�o��,��n���Jb�4���>T&v|u�ܬ��y8��f�Z��x�[��S�+��!y8(��(�H�M�e�bv�t�J�;Fl�����>5�Sa}<yV�T_XaЌ�
��X���RwJ8�6W94��F���jv�T�q+�ɩЧb��M��<"��K�ՑB��Է�0Zf^#Y��NgR����8a�q>�]�s�X�&e��O15Ŭ�(9�<f۰&�}��ouڛ��ks��	QqS��W.ge���e��ʰ�����xc��J��r71m��c�a]&�E@�������-IObƿ������*���5�>��F��W9<��y���wF`Z.�N��,зq��Ӱ�=�{y5�X͢�W��VtUu�ε��wI��*��bwg��u��ުnުv�:�������s����d��&���Z�1�ǒ]��K%��m�=1Yjr��%�t��;�m9u�4���Î�=�S����yG�
<�K+�r������\H���a������<��/y
h�,St�	F�)+}+�l8��.Z���=\���κ>��o.��]햄�GY�{evAi1�[�n݇I�9؎,�~���|ι.tOe��u_~�F�c�ҁ��d���M��M_����e2Bs�@�s@��t��	�霡��q�w)�:�Q������.<��s��0.\vS�ЕkQ�>�p��,��{GWm�^�'`W�)�uޥ݌o_*�S�r�K��>��=�@w�H!��U�+�T>մF�ܝ����Fs�	>�m,ҹ�S�^Oqk�#S�P]@� �2L���ŝi� u�K\�"��a��.ՎiZ���__Xom�Z�,���-QH$�T�F�!�X�n���
�T9�	��J����
&؉w�>�N6�O)3�A�زF]�hvu���ۻv�x�g�}b�b&�����hc�C�45ɞ��K���°��sP��b�Ӱ�z�-)C,L�������C%7U�:��dSR����]����dpm�kz�k,��+fc]W(E�:+���uo��������ΰؙ��6�lr�/�#���v|��Ƣ�ӳUY�_ۭ&���:ps����������FKSg\���@�A�lgF�,��Nw�����&��7�S�g�����C�1M-{=u�kL���Y���e�2�L��:\�ۏŪv'6A�yy�>��à�)Zk��,�}zf�������B��INC`*�u;���Am��=T��ۓ��&cB�B&�Ժ:��޽=y�D�s�T��݁'��j�kߴ�{�3o
�j�w��T�����r\Vlo�nH!���)���*W.z�-�`�.�m��;j��<�k�4չX�ë�D�����J�Tvk���O\�U�w���?v��z�7/���WV5A�n����F�4t���D䕾rc&E�x(u12�^�)��[Un��	�@w�CY�%%\Q}N���Y�0n�����z�(k�	���lw.���r{�M�5��g�1�f!�T4�b5�9b�钏+��ۥ�v��V+�d�~���4tJ�%�3p
t�fK84
j�&�� �ȣԯ���-�]l�E�ٹJ]�|F�>B�c�eM��/�ȯd��e����z�ݔ^8o�!n�Ka�-�N��!��ҍ���to�5���C�^��P�|�p���WS��7��Ѻ���.�������������פq�UCN�..�U��}{�Y}u���wm�*�mUx�aߡ؎D��g�\���Ȟ��Р͓B�j���^��X|7�����Mw�H�&x)ы�P���V�j7N�ֱk��Z�ڜ�F�:�ߵSv8bCh�	�ɯ5Xk\��	(͆���d�N�<���Jy��4����s{�:�#!�nP�W��%Ɍ�l)�:�x؜W���侕�k�_��-M��I��''�0&��"��0�����5LfWe_�ޙ��#�_��GKc{
q�{�_zv+7Bj
���G1ة[����}Xf�;���	RKw����t+�[>�uTR��8��~��2��5Nä�g^h�+6w�%����nc7G���sۜ;�����}Ѐ���j���,N�?���6�K��W�7�ۅVZ�w�(�]�G�	�e�o�t��#��v��w�Yc�����eط]s��օ���=ӓ�v>/#�0��̭*���Ѣ���s�Los�>���d�~e��e��{�ޕ��\#��+2�@���l��V��{�����>��Jh_Roj��U����n�%S�Z��;X9��8��z4)(>,X�N�9��]6)[��a'޶iI�Sцآ��.����,r��0�IA*.A�6�����C�D]���:�
M)�ٛ�a�����yGyt��T��n�ou֪�j˛jV�G�sE5�mv��䲚W7O���۬"���	H#Z��3��n]Mł�M��z>?/C7xwq�Sc\����øv"}��
 J�33sy�5W%�Yz��rw1#�oڝ� �낷��	y�k5j�����L�)Q\�zRS���A1�2�؛ɼnhfu��NݎpĀ�5��%A�qzqB��V�-�LF͚�9289������y>��f���4����/+���i0=��Dս"���u�! �*@�8�]p�Vh 6'J�躖j㵵�N�-�:�S�X�7Jl�4��"�uF:����4�m��P�	D��}�^�	^�"p�j�t0�:!���R����H�{á6�4c��+�I����-nv�����y]�~j���Ft9�p���=��*��bm���b�5�8�k�uوP	����V���{����̕N OR�����v�6��ܰ3�}}�:7=���f�}zf��py+tc1[��؊�-�Ҡn0w�-7+��������S��:�������&�VO���E+f6S�)�0%:'�����]���m����v�<z���Jn"�;��n!S���y��u��$n@lvJ�:�5�I��M'o2Ea����%&1���s���~r���+�l�����|)(�V�qn���qmЄ�1��lwT��|�s	P֣��.�+*����p�V�[�6.y�N]�ѻ����awoX[mUӽsa4�s�X��D�Ӫ}�#��Z튶�
����Y�Tj�W;��-*�y�=�c]a�z�m�)J�~.n�D������7tK�X�����V�Ӭ�|Y#�����s-q���GW;�n�.%#pޫ�����d�����9t�S���k��=[�W�zb�S�����5�1�v'1�T�c1����Ӊ�B�gK.Iǹ�[��{x�.�em���k]�����O���!k#l
�T4�W�9�ҵ��P/��o.0j:����������BC5���|9B��P��*�e�r����1
v#lF�x8���X$a�l�u)�T���ˁjOS��hmn����ܙ	���͝d�৆(.�	�3uݶ%�۷MB�
�1�L��^V��c��A�d�2Z�:����&X�p�*'v]����u�Oݘ�v[���s�(4������=�
*a(�ƅ�=������=*,	o^��*uzX�a�̥a5��Գf�lL��
����Go���<e���rpOI�J�91M�����M��M�:�c���\�P��Ry��㞚�*�W��ƨ,��	�y\k����&8�X����&�����<�9ٹ��qW�ؑ�d7>8���}�*(fR��p0���k%i���$�@���C�B���	F���*&#�:�k��FQy}���Pc1��*p��7�\���#9��aV��и+qd���
��ʆ������5mt�N�ǛK��P��N�]X�ն���e 9W0��8��ro�ɚ�r��lݩoZ��V���O8�ZĮM4ʷ��öA�����a�9��"�|� �8��sW�ܹ}�X�����T�2��l^\�n<�ע�j��Ļ�-x��L씢F�9��[Un��	��lw}g�ޫ��P���ܠ�*�8�#�N@,$N�j�;�yq�i���þ�nA���P����V=�}�rl�PU�JH|�L�b���\9��¨��ٺ�����ڛ�+QY}a���
4r���H�X������T��54����׮u��P��;<����jb�i�kN:�p��2���x������ܸjƾ�����_Zrd&�;�b$rx"�����]��7=Z��|��b{�Q2I���s�C|��E�Շ��n���߫$J�����*�,3���7bo's��7�á��4��v#�U.�9��޺wɉ��x�7Ɠ:V�/W�gCK�U����`PN̂.���)�u*<�3"��=�v����z�E���̃dur���!jV����a0؍n�vݢ1}#��w�����gZKf�������f�ΙiV�����<��5������R�8�������Ö�o��V����ԗI�i.}*�@{zg�/�`*�mҹɓM����@ö�`�ge���Qby���������oc��5��<H�*@9-�Q���C}vNml�JJk�����n�T�I�9ٸ\U��"C˭������v6���������\4�o4�w�b�&�3��Ga�f�_m��(�j�F-�mW#p��#�qb�tm�;}I�i��_�ic�q�Mg���A<����z�垱���X}R�%\�}k��[쁛�fr�l2�3K�#V�<]�.�OY�������(%S.9E�o�a1W(��f���Lm�S�)�}Ԟ¬}f��@Aw�Y�L���������uh��q�Z�s^�沚W2�qy}a����#�jӣ*�;�a�1�2�5;���0/��l5�y�[o5�a��p�����ٗ-���k�	M_q��l�3�]��[\�ݦ�}j�l�q&�����پ�������Q���#�8T59"ev��f��sz�MŔ�uJ�;���]ʀ����̔��n���M��ǌ�L����q�-Lk�����dLn`��,wu*�Ñ�9M.��f��k.��zf��t��J��#�Cw�}�5�N������8;�w�u"2Z���w
r��wBpI���	L��lN�.o;hq�C^n�Va�Q%����F!}Q���3;n�T��TT݉�⻭6n��WU�p;��dɠ�h�+�H.yCQ�V.�b�Oynl���Ws��٠�cv%+x�o}�Pq��)r�/l])Y/y�Zflg�����D�;�햕d����xlV�O��%��/"Mt��+��wR��,��ʺ���Z�u���w&�9B���]���QJ�t���ܨ�Z�7���p�rF����'|&<㌼rR<���� �&e��90Sk{v4d[��3r����+�V�Qft����v�J�i<��ܟg>��<���vv��"lW^��=��>�Xl���!٧:�j�`
�R�p��wo[������ev���D�!���i�
��e�.��j�u2-�"�^8>�X�<��('���dx�γw���Pm%&f\�.%�0 A��WktVJ��(��f&uݞ7�喻l=��6(�����"�Ӕ�G�m��xޭ1 ����qj�H��k|�T�w>�҇@ձ�Lq���v�/�B�-œ��n�F�j�)���#w��}Υ�3wz �!)A�����;F�R�x���2��r���UއD-΁���� �wl��/��·.��f��Z-��S�=�p}��8�MT9\�X炌Ϋ�e=�k
|�����^�C`b|h�m&���9Z��,��o+�`�Z%�j�@)�i�x뱜�P�y�WG]�V����),Q�Bd��vW5�]tRz�io�Nj�o[��]"�1(�'�0!{����&��+ic %d:U�u�y�(�W<ۜ�>+�,��գ@7^d��53��JwγS�؍�C�����v.�"$!�(
N���P@�]7U�Xl�ә�1em�z�Nbu���+2��Z�I��0^�D����p��4������AQx_w��3����	]Y�켐R�T�Ǳ���pixu����/���Q���K�������-�_�]��_Ib_���ɻW��X�cf��9=�	��ʎ�f3�h�Q�#u�TQB@�ˎ��&5�ckxo}yV�S�e��j�_��d*�.����M�b�j�:Ik;Q�%��tB�Z{��b��q!�֩독�u�2pK��ݻ�|�>�`��h}�H�w�{�y{3Ц���í9(�7Z��g3ǁn��X���
1�"�-@�QA
��0H��B�T�
0*�(�R�AE"��(-aP�dP�D�bTr�
�b������[eH�V�P�²*$�,+
���AAGmmFT�E�!R�*�PR[AKKD�Q@Z�F�E�J�E)RŬV&$ReZ$P(��J�2P�
�*�`��*EQJ�	YDJ�
���mb-V��eq��R"��"�eB�aZ�4����ز,P�FJ���4��R�*�6�����±T��j��Rѥ�����*(��V)
�Ұ��Z1AH-am��X
,��ĩ���,D����[eT��U��d�X
��D`6��b���m��)lb�--B��*K�Z�(�b�Qk*�0UPU��őLJŊ
,X(���*�QQVF�TPEbT(��Y#iQ�#��
Kop�����er�o�l����=�.F�oy*t�>�4YS�%�N��N})N&Q�AM�]�h9�z27�}��r�f9�Y�T���+��Ӽ5s�-L=���D�P]Xp�:���r�o��}��߾tf�{+Y�Wki-xk�]~MO��O+�ے�K��ngs���\�:ѝ ��i"��ԡ�5O�|~��P`�>l�>�o3�eRM.�/وc�6u����\ru�g�+\�}�;mOv��"��+�b�C��6���V�rphs#�8̕�n;Y�����"�z2�L�rok���s�1
	����)�a����`o�ڬ��(�ec�sk#[��?OLW;�g0��Xt�Nî�n�n ���z�$����S{f)]����-	�:�؜s�r��P[�[A�a�u;7	���Qx:�
���kMwC;8g%���K`�״�z�0����z��Efjkr��;���=alHܲ^�)��"�ͥ7��B,]`�F�3l���5��V�e�BيZ[��5(�u��`ﭵ�5�
gl��=�YBl��VRM��l*B:��K��lM�ْ���S3]��w��v��s�V�pq,��T5V_ao�k�u�i�^I�gWR�p�)Fw�z�W%s�Őp�\zSEuc�9X�{
��<7$���~��]O5p��6�MV���Q�-uj�t��J��^�֬VUþ}%��]b��KsW+Z-?ȕi5��/S�sa4��.����,�}���E?bl]��W��ʀX�o*ggź�=�ƫiKJ�S�I�-sg���ȗzt5r�`�7���^3��Tk;�ʰ�*�|�j�j�4�KSQ�#{��V��5�kDR�Ժ3S�"|�Pq�����w��f�[�P�i�u���:;i�m�LM��|�á�L���47>3د�0���t�8V]
M���m#��^�Z�q/�%>�9�C\��xb�x�ͭ,�9��{������ۤ�o-R�g[����m�2k�V]�Z�K�����	�x�2�N����5�I��u�\�����*�֙C.\�[�N��CAڭ�g�e���Gt�]�}��#~:Н7��w�w���op�	9g:U(��Qs�{I���Xn'^��V�Rh+�żF�5�2R��N�H+8��Kd��F�A�Oj���WK�%H��*��tʋ`�Nf�"il��;U�RJ�Y9Ϋ��O���� �)Zk����	���U�vj[]�z��]G�
�㎑À�c�ш-�����#!���hL�M�{�ޓ�M�j��8���
w��(s-ܞT;%���
�c�J���Z��OL갚��>g;7%�X͂$nI��K�	@����m��;���ON����-�8�ZĮM5nV;g��#p�V��k3�.V8m�(X�v�Mz����b{�>��ڷl�-�+�']S�r�Cr�9ʲ��ײ��7��e��c��}mUӿ�l&�w�k.��u*�b��Ժ7�ޒ�@����a"v�j��{�����O�����O�m�;��������4��=�>X&vN*����';͢Ѧz�Vy����w�U:|輾��D� ���n�#���<��������ۺ;v`�}o����.`�mP�K[Ͷu�`~*��
����-x�RiuM�	+�E�õ��˅������L������m<�7L[�gf9Fi�������K�����X�GX5��p��ʺ�-'ݮ�ukm�ۉ��>Rڞ���ƨu֚�j��C�9I�
���M�۠¸�U��:S�R�ɥ�HG����>��>����з��F�MҚ02x�IQ�0�1�������s�e�M��74gZ�U7�o�	�ɘ�U}�x�1�6ә݋Y��E��%��xb���fݬ��nou�\�z��Me���|��e�ʿ>�3^�2,7 �R�Ǖ@�F��z��`.�P��n#MJ��9<�,o]�0����YOk���$`\���J�MJ�{��#���h�y��[;���<t�:�ޭ��Lм����=F��\��3��'nks���ɹ]q�%ze�	�v'L�f�\U�����`WU3�׆r��O��ЕE��^씬i��i��X�A4�gZ��f��zI^I��k#=]�4�����e5$sP�єԡ}I��ik����;��H���T20�k�ɘ�����7L���E��4\���E$���g=鴈����������Y.�&�=�I��K��Z�\WN��U�wá��:c �Z���!nQ�2 �<(��۽]ӨPk��X��jT��˷n�`nwt&߾����:[�)Ծ�A�{�x�sB��MTM$c)��2/j�����%Z�uc�)���(%Be�<��kug���ALV�.�>��v���{.�uy=�X��P1�]`��r5�M�sׯ�9h�f���U�RҩB�*//���)8(�{3���_&*��O����IO��%��8�Ϊҹ�����\�KS���b�+b��w��]Epi*��:�w=Z��ki-{\J��h�yة(�1�������X�B93�Aъ@2�X�ɼnkٝjoS�Q�R�N�J	Ա�E���A<�3��̎��f���FN���Np��ʓ]ڙ�U/����Z�l�y]�`5Zk��rs)c*&)M���+��6i>�ݿ{6���a׻1�h{]�a��L�\wk�^�X���c��(�U��0n�HuZf��L;�c��i%}K��P���Af�>阋��Jn�P���ɳO G\�عE��B�UA�s��6�\��ɭ�A�sFg}.<�jv_"�C����W.Tٷ�\�V�.�hYWu���n0Z�8p�yy�>��ç�����,��L��je����ǔ ��瑸~H�*Nu;��r�j1KM��9����~�°EW.�Rk���ج�,�Y�{�������-�n��ˉ��./xj���^sU�L�b�{O-�����%O�xvJ��6�k�n5
]
�U%.���Vƚ�z�,|���=��zA�zPNJ�a��ʪ�{�z��p�j�M궹���k��ւ��F��ieۈn�d�.=��P�'�8�v�;m��N�̈́Ү{
�>�A)+SH�5����]��<��[�B�N�J�;�VҖ�J����@�n/P��El#�].�1r��#T�8������t/��Q�_4�s��u�Ss*¶�[=��z��X"S�PpF�R�D;���x��Ek�n�>��֊f���εx��ݖ�[N<5��|N�:Gz\=���u,������y�u��!�퍃|�j��m�l
WwGmz�P������aҳtM.$��|�P:��ݵ�i�J<��i�vV��;�������=��e�)V�؆u)!���uf���g;�O���z�S�hS�C�5I�
47f{�FQ�h���fIbn�J	A�9�]-�~��ۓ!41�9�Z��28b�AQ��i��?eN�Ft��r�z���^�|��m�y�%���]�������E�+p��ܻ�/�8��M��{�-��>v�]�=�ʕS`�Uۚ�8��.G"��UNrs)X�s�v��r�]{��U�u�h�k�6�{�t;��+��u{���*N:W�ɓM��F �%쫮[��;^�{<�j�n���7����lh��}�T����O)�C�Y�{j+xЬ���AI�ջ�t9ٹ�K���>����tn�v����n�os�7��.qKm�Z�b�i��w�},��������N�}��\��t}��S���j��+�c��mQ���a�H�y�X���#w�93-ҭ��o�vt�[��ղu�`�ĺ�_e�)
�F�M[���}˷�Y�M*+�K���
\�&�����*��r�ͮ�{ZLr�����ڛ�Z���ucśK����p'�;1-o$|M4�J���,.D欼���o$��Ѱ�ѡ�(.�2�(��s�SU��`&�|];�q��Ǔ���o.��~X��}%W�#�����	���m1't�v���J�VŹ��gtɛ,
���oqk�)@A�J�|�L�b�0"��JṇF�M�\��KX������u�7�%8(���k}M�xotV�uoF��������%ap��T:�MUx�a�;<�ϸ(9=Nz;��ͻ|Z���]��/�=Ev񭷜Ul��;�������hc�v#6�n��9EC��ʚ���,hS�X�	��ntfu��T��%�ee��Q�q'bv`�rObGK���ɑ���� �7`M��g3M��7���e�M7X!y�%C�{�������ܫj��xuAϬ7'2�Ǡݬ���)L�d��Y3�B�]�k|��ٔ�&��Rʿ=�3^Pp<T8����lF�ʙ�r�m��Re���(V�=KI}1��V݃�l]��񉐿��Xw�}��ldܴ��9�w�uiˆ�\E���M٤���oe$-��xO��+������ma�3)���#��q��P�M���ګ2����k52zeG;�ͧ���o������ަ<t�λ[՛ϯL��~��+c+n����M���	��k�D1i�]b5�|T��t���6���V8��Q.�a��#���D�M>U��J��o`���J��imQ+]j�ޛ��Os��y�b����T�ΡK�vښԛ�4�ٸ�;�G9Q�
��kz�0W5�
�m[�{
��>ᣤ���,ID��s8��fG"(n�o$�+j_�/y0�֣�c�4��Fo�X(%��������z�Rڞo��9~[mT��(z�u'����P";˔����:�h�ݥ�˭N�ȽY���i�w���iT�O����a�F�C륂j7���\���^H!k�kP���\:��������/�16�7���v�̭����\Q�����ϫQ�u�i-q/��p���յ�^3B��;WvcQ��1�ʞ�hz�+.����Z��B�(���L7Z�ʌv���|�m����E��V0����y�2˕{]+-�Z�H�`1K��Ҵ�E�ƧDxc�M�
�{N����,A��������墑è��p��e���9�Ζ�%gz٫�s}+����W���������]�* 3㾕�wm�V��p��2|1؅6hk������o&+/����cE
���J`f�S{���p��v�U��џhs#�9��n[��V�ʶi���o[n{1���c����ho�[^{]�a���x��4��{�N$��Z��N�925�����0�Z���S��u��ɌW�r.ӸwbxW����Ut�Q�N�8����-�T��.n�Q��V�N��<��=��_{����yJ��ryP씯L���wwP�����p�q.����\�;U�����b��i�l#rHlu	@��T>�t��b�Q�%[��ޗ�\�{�5�JᏒ�+�{
�rAA�xZ�¶�QQft7�����O�ћ�>1�I)t��R�x���ڏ�����$��B��B��`IKH@�xB��@�$��H@�xB����$���$ I?���$��$�	' IKH@�x@�$����$��	!I�HIO�H@�xB��@�$��IO�����)���D���/�),����������00���q$����$�q��J,�m�6�!�Q@�J�H�d�ݓU�-j�Y�	���\���j&fU��m��\cZٴV��w
�q��ն��Z�6̢�(m��7'6�j��fųjҴ���,�6�3)�bUg9�5�kdc6ٴ�V�6�n[�hv	�\�v���3�+ZͶVԖnmͱm�����8    S�mIR��d��F4B)��%A2i� 0�M@�12dф�14�&����R���     4�ɓF�� �0F`j DP&�0&�'��LO��I���Og����W��I��D�ꐒ��d�`�B��BH	�HH$k����A�A��fm$T�		)�H� �J�H�8�$!������f�}����l!!  k;*�R����Ͻ�麤������~]�_���m���9y�+r5�+ou���w��H`��X�Α�)��5`���p��N8��X�unKP�-V�"b���;�4�q߹��e�����ҚS+@Н5�ڼD��̆7`��Toh�S@��aTan8SW��L�1M�W���u�Kڴ�����0Tv�i(��/%�݁��CpSĵ=*�@hQ�v�Y{�lGa5r[�4d�!j o��^�Ŷ��`��<@e�+ї% �
���ݝ,b�x��lb��ݡt��B�І�mh���0���]�� �V��rY������/V?XЭ.áGE=�C�˺�v�I�2�������K^����H;���b4�.]Q԰�t�N Ct0���NR�7I)�A:��t����@C�	��4�w�-{Hݸ�y���w�%J�{��Xr
�Ncn��D�䗻l��벵b��ƝT���k�{��b�e�.³�������Z
jj�X4�Xt˖A�̫�g�E6�T� �a2j�rW����d���קF�*ԏcx��KʀQ�,Z���'z�]��,�!
�3h얱�)����%��-�T�����6���4j�i{ �e�1f�-�Lkŋj����Y2�a&n[�))Cp�Z��VU(�Ȕs(���vf�84�&���tΆ���&l�ϑV��Ŋ�`�"�n;CU����� a7��

�܏ĵj�7	���Ҏ�0[�J�o�η>�5j[(k�CU��B�4EG��s.��(f�͛Z2����C�5Ġ�CRA��z���	b�a�Q��T��"����"��LGe$cA�B�sj-������bn0�U!P�']���t�h�Y��)W�����~w��Gr��[��s��tN�dyJ��Y���0�Z���$�.�*�P�J��h�xZz��(Q�Z(�X+j����yX,6e9���o)֩I+�	��.�ᵫ�E�� ^8z⼩vNl����q=N^� �I��7RY>�ʲ3�+\�w�������MST� +6�2�RS�(˘U�>�^P��[E��e=X���é!�ʺ9Z1�w-�"��O������9��ZhH�ç} ��๯Qm���5^nf~����u�� C�\��0b�,�AŮ���D�̂���Ck��6�gV�{������r�\�hU�4��V�
OL�4�L�ҳ:�J��Fqβ�.T�&�Qޠ��\�A��r�!�+{�}wn;��)�7��LÐR�-�y�\�J�"N�PS�^�
ƚ�;9T݊�R��Bҝ'��-b��P��\- {�=V_�D�83ĦꚻF�_r�w����$�+�V��ہW]���ڱ{ȣ,5��v�����i��gE�����˴�x�l� e�{}Hk閠nBj�eh���@1Y��ގ�y]�n����0�7ۺ���S�Cr�	�>���@k61� /9d�V�*�"�u����d�8j����<�A�s{Z��]�L��3�aǴ�f�9x��8�􉬸�-�9:�$n�H/�`ј�X�]����83��w��tp�n�Y�p��;�fƇv�Mޕ���v8�WP)E^�kf�,%k���$��ڶ9>ݽ�Vַs.[zYE]�N�v��!����h�����Y`�wL�9�s�C�
����L�����+��՘�3VS\�1�K���%��vyP�oI�nPLml�]�gـ��]�$lՂ
�c*������N���+x��mt΋3��9��7�b3����#�y2.�&����mlT��&��1ab}�N���,������Z�e���u�t�Z�۽;HѝB�Q5�o���b�T�ŀ�|�V��T��bh�n`�� �3P5I�����|ʍ�)�[NN�s���;/ �=ժtQ��ܹV�T_+��ĩ9O���uCM���xW�D���(��bY��>M�v��M��&T
� �u������ŉ���P䪋��$�ݷwP��Տ�j��]^�=(4�#��R�J�%ᎅ+ѽ�{��C@|���v��l�5��hU���P�2Z/ �7k{�,mE,��X�)Dd��rMx�O�x݄/��$��F� �u��;���ې�ղfj33�����ž���za��ys�t[;6��G�QDZ�]t|γe^�z�=��o�o9�Ys��x������z��C��ߟE��	! y�	x�d���XH�8|��䄄������]>�ϡ���V˦��֜W��m� �Y��T��Du���B��&���e�^g\�MSKzRf���5��v>�ū�4�+�L]��4�H+����Ty��J�r��#o��N���߅�\�K��WE��Mˬcf��`]&�=ǿh����;E���K�[YB�(��Z�+��Q��K4��?1ln
5�"	�����Y��٬�F� �ʒ�RW*�P!v1�{.T�u�+�N����y�킯 �'�K	�vl���ǀi���"'xM�	ȃ��b�WWeޱٴkN�h��i��}2�	
c���*T6N���QT)�n>U�%�lT� Z��v�A6&���9)�HQN�ID7`P�b ���,Nn��>����c�+����N�Hf�5]�b�+�����cؤ���m��u�@*�R���^h���ZL:�s,���;(��(�u��bó���/6�������)��C��Xmm��<X��|8Xz."��ܔ���ؑXu҅�Ii�H_PQ�����w�ӵre�h�5C�Z���)*Û,u9�)*rhR��h�#(���͔�:�y����S^�&��5��sb�Რ�>�Ux.�N�Z��f�P"qPo��*�e↭�PJ7H��zSۭ�x�O/�B��Q)��C@|
�3��-���U"{t=8���@��E��kKp�WZ�3F}��Qr<%,Gf��H�SZ{���Un�9�n^ܴH�wo0(��a��F4��\��ڬ�V	���ڽʴ�OoWi��PٽW"v��%��7KkN��8r�ov�]3��;�1�kN\+�\�++T6��s��@��h�z���%��nS&;&�d��"��c��[(v����{���U�.��rU���XMM˒� ���)��_wm��N�;��$̎�%!�]��t���}�37��K6�l���b� 1C�_�MGu�$օ4���2#yQa�csP��V����^�Cq���DDB0�*K�t�f�Uxl�����f
X�u��
8�4�F�O����&�f>������iv�MَuBt�ʟu��9���y_� HH+"�������-��>o�՗^ɨ��GH�c�d�/j>6�i
X�Γ7��eJ�.f�{Xٳ���x}�!�#�_��r��EC3��x����6.��Z�V'K��mܫ�@5�D�n[Ƭ)���ãy�g�뇅���EURS))��r��4�T��r��@��&H,���
JE#������\����o�5κ��f�o���;b{y��ƥ��m�$<Q�k�S:6�����n�h�qg����i02��o%�{D�i_�}í�
�}ޫ��w�~�jgl���<�P�*6�@gYu���|���{��ny�mtݬ�âL�!�G�n���Yt0E*��[���W�^&�sGI�� ۭ�Qn��0*I�Nǣ�1�����ūc�o��j�
��ư�6,�<�T�=�g���S��z-�׍wqՆ�(N3^n'��Q�ݗU�7>Aj��l�V\WF��8(��@�������s$h{T��1R{.�d	C�]p��"�j�lqJ��ȸ��ד-���u�kR�jyk݄՝,����PV ֦��@Q�M���_#zwa�]��SX���C^�%�I�����)���~��G?���Ş�ƴ;4?:�2�5Vݐm��S�i�nNZ�O���$o���S��&IB~Z��J�y�*�$7�T�r��Xw�T0����{�ܩ;��?,��V�^X���o8*�B�f��ju�6%R) ;�U�p����2�wm��0-�К_�����]HA ��
�����#��ٹF�xc��ѕ<�<*|&�\ͩ3�+(�T�!ȣX���	�'w�W��+���\X��o�n 2�;勑j�����~wM�;;���� l����1�X�J�8�;k����7}&�/!f��Mjg��z���n��vu�ن��U�θ#�o�KB�/'u�����k��X��_'�]_�S9���=CƠ�@R���8wrӋ��9��5��^��@�˪l�i易2�I�;U��,�V�[�Z�S�W
�n��ߒݔ�ɻ��>�ҍߥ:�-��EF�g�����3�����~�N�/��w�W��;�N;�u�a����>y����]YX(��L��q����Q)į:��8�>xW�1x[BΌ7�F��LR�rnǳ�>C���gJ&�l�g�����렏N�oQ-���(ēb�~?��}��魞�L�p���e5@�C��T�nР�ؘK�D�í�5��A>5�C6��{�9�5��%��M�WN�d��o-��tmK��t|�֓s�WU�	ɓ��0u����]s�����Y�j�"���`��<� �U��"*$UX�ň2��R�R)��*�I���H��b����*�L)�`�׎�{�|��*k^$sOu~��z��.�	�m�Ѯ#r�S�[w_z����5�w����>ݰ��F��fbV�<����⋈5HVbz��Ke�*��p���]ۧ*]d����F��{�SԊH���gc�q���F��f�c�/�w���`#P��y�K2���޶.a�,�� c4X��S]����%��؝�Tc��WI����Qb�O�#.�x�y�Q;�ݵhO]X� k���H�d
xe�g�.;Pj�b ��i2��q��pą�K�B�ZB�������?wm��V���3�ʠJw�r���)K�T3JW�X�ff��ڇ��}n+>:��>f��	����ګ�~���+�I{������:!�MhՅ��_�uD���l����)>�n�z|������]�Q�ֳZʏ?�$��+Rx��b�P-ڝ�\)u��l��~>Y�=���_����O��uC�Ϻ�g�KC�ѿ��TV]�⦴��K&c��Z�	��L�v� �+�l��(	�c4�m�y�/1�N���ƴ�Q��-���iB�v�)_S�!K-��(q���D�z/a�Ӫ��[�L(�m���z����$������1����C)��,��b�z�E���� �����u���;�L.~C}�hnDL�����2^	��0A�)zY�Ot���cQ~ts��n�v���#k�V�һc�-�ّG$�����ܸ|�K{�{��²\�^������^Y��v�Ԫ|���{Y�U,�.����-n��ܞ��_'�ly~��{޴A��*Y�E�e�d�ʋ8@]~�s����5��Pٱ���қ�C��G�vv,T<�p5tC�n�ƭ)Q�� �ԧT\^;OFL�G�R�o�P;��#CyJQxMO6��eZ�����3�G�Y������\l[̴����cyCK�NE�7����l����M�w�o�����c������w��N������q5J�Q���c$�]l�W�#%�팽5�
Z����A������/��S[�ҥ9�F�=u����?�o�c&�St>�6dT0X�,�A�+��}�8����Œ�&ʲjۤ�]�����ɜ�KI�ǯk8Ы���^^��^hMN���u"d�4EN��9:urŗE�XS�ڷ}ݑ5�v3�]w5��2C��&��X�"(�*�"
�1J�������EDEH�Db�R�%4���#���J*�Ab��F*"��E�ª��EU�,V(ʪ�לg�3�u�>z��fb�.l����Ym���i�-���O��8?�'�2����������	=�?g�\�"��퍜�/�u�lU2kޔ�[l_ˠE�܎�4�77sw{QA����v�hx���2b7�K�VMw�<�)��l<��nu5��'>��-�=~�֗�>�;�)�xW���s���@g~�U�ۯG���s��}�;���������u��A8{h�@� ��o͋F�P��������w��4�%�Yso+V�0^��mdi��fL>]Sg-Ԍ������{��ػ���jGZ�XLc]7A��[9&�3�x!v)W���������3�	�׊�tI���YMу��I}�R�Ff�IAIy��w4Vp��z�i���6������5?fӘ���S���峰In�] �1x;�kJ�y�{�W�œلޜ�o�#f����L�7wEO���F��e79?�֜�e�:+����٠����~H�hF��Xs�SѰ&^N�ճӤ��`�}��9k۟"M�S�p�ɽ��ۚ�>����[f�	
�}�s��~'y+?�s8Z'�+hFd�~N��u�*�Tu���N���l�.�ze���:�^����NT�2I,�cX+����c>8�f"�o=���^���֮�V#��}�ǽ���W�����:��ox�^,�+̝���Z7�.@0�����$�a2�@�$�[$�0�JH``i$�PY4�!�Hq�& ������@)�l< 8r��,�4����� d!���E$�ᒱD�L��Bi���獀�$�[$-Ĥ�m���& �{q0�A�S�L���xB��t��1��q$5���CL XR@;`[2�<2z����U��WU�1SҌY�ɽ2�ϙ���>f����'H�y��e !i&3���HɆBI4���2�v�2CHB�!��O,0�L0��ZH2�,��U � i��n�&�[e$6�BL]��<��)J@������a#���鴃�^�Tm�>�m�Q|�P��`
g��� Um���\5����N bU"��|������R�yڱ�۳yQ��Ū��6@n	LқyB�Rg�
��}�b��'V��rʗ��Ճ!j���U�뒖l�gP����l�����j���Z�܌�� �VX�S)Vv�ge
�2J���)�N\��ϲ��y��w���pA�P�]��!(�K5�GGƖv>	�����]8�eS�[vug��u4�.�2D�ǹ�!�w�N������u�+
g�z�.ǻs-��A�d���S�]bQe�Zj�E�k[`bǈH��񃭆0R;Gv�I�Cl��&��A�jD������Ԅ0��_!��ZET���(�4ݚ���E�
�ETQ����Qi%Dj�$Qi�Zi�TS
�i�MUS�RS
X�ޯy�{�Gfa�L�������x~�����M��ѭ�	���sϳ8@FZ�%m���}��2�<���jv`l�6�{-ث�*?[֎����'�2�f���g��|kbj�+4��qh{�fo��y<�+�L=gi�pٴ*��s?g�B���%��٠k��m�	R�e��b��Uv��LD��u��hQ9���+w�ZX��.����]/ׅ�8n0��0����yf�#�|�7��ވ!�q�{�A�������/�늲���b(�$.��P8��6�y4l��]�/�G�G�W�'u�[��\�5�45��[u��SZf`y����w1M�zt�^J�џ�3�z�� ��Wq"xb88V�����؛K1T�YL������j��������nQC���)�2 6�,)0�Y�D�b�j�z���HK�7���μ�k�	�<���]�������8�nP��GF��P�uލ�P�O�\���0�]���nbV�u��W!���R�bJ�vS΍Ǎ7*#
ٓv�F1E���f������O�io�3*v��wߎ^E;��T]�mN �{u���u�n*��8<e`�Q���]�`!��ov؏h���r/
�v�o�վ�E�՘�:
c���V��I5i�t<������kS�x��V[�GSD��?7Ϯ��UŎ,W�@��C�]i�t��|����E���I���ŗ�W�k�5~f.��6�ܽh~�����\V��Vib<�}�}��z�K7Du??���V�CjuF�LN��F/!U�}hۧ�(���z��\2%݈ut�l�w.�0�7U��j~�W?C�A�mv���1V;�m��o��3H��y����;�ڶgn=�=u*6��ډͯ)xN{��*�jz������Z4�Aͺp�-j�<�[֙��y��U.����C�?L�طV�����_U{��P�H��(��$�3�]PKɀ����~}�N�<� �Űm��ʶ�$C�ّ��������qg���.�hoQ������
��fBJ�R�q���x�I])��i"������N�ڻ������M�X�5F奔�Z_P�Fê�ދu����d�f"�vtn����z!��ɧ�rv��^��x��[�_(sN1%Ѵ�f�wxRFe���v&
��8,�l֛����s���V���Te��r.��CL\���s�\��:�]�_gl/����>�������UdcU@�#"L�(��UK
����R*ĦP�,J�Eb�1��(�1TF��TTAw�R�3M�TX��y����'��W��ïO~c���ˡ�e��ߣ��B�<��/ �����f��{�b����!п俷�{��(�黛m艗��z�T�o+A`���}����ǹG��g(V��fZsv'h�Ҹ��s��~���C1�� ��2���Z7Ji�DX�GE�")=�-э뢦�׆���P&W�$�p�R�࢖��)${f���ά�`��Yd*���
��.���GM��'���~ď.���b��'B0�x�ϙH�&���u����n,ӗ�T��t�D��}���A4,����f��{va����O�>�ly3�M^-�s�K�4�>ܚ�E�>�T�W��I�p��5�@�G����j4��u��.{�OTE���kL	
�|�w_]M_���~��<�����6a�c��]sR���eW��5��82��޼�=^��������M�j��h
���#{h�	\۩��ө@:Cӿ_W���P3ν�~���ʹ��@!�!	ܷ�.7ob����"%��<��M<R��,b�itl�\�k�����h��Z��r�Z��|�z�2pVf��諾��Ȝ��<f��ݕ���{I�t���q�!Y��痚���MI�޵=��wr��Oڃ�{n$��Y�Ahv�/U�x�ל�T�H=�3|�ݶ��հ<�n��)n����Ƣ�0�h����J�:R��=�D[dN�cLvC~��VW��v+��=�$\����*�({ٱ]�{���;���=��C������JE�d��/eoaۻ�W㊻��N��O�O�{�A�Ay[�H�ټ��a���B��A�O�/Fg�u�9n��f���4�����ob��WJa#Z}�aR�Xe�Dh���o��"m�褝��ޚ�Fm�:]�~q�;qV<��ׅ��=��~l�oiш �Geڻѿ��sK�D����9��Vgw喙)���yT�{(��e��3-=�Zy���m��u��Yl��?#A��AHMc�'wR��4�/.#�}r�[5(	rmiHV�iwT���
5�(kɼ���M 4���g5qWVg%�-�A$4.��N�6����;3ȡ|�+9M-����s��0k.�*�'*�-@>U� C<T�ɢ�iN]��"Q����Y���ZQ)���TJ��E`��NT���*��i�tUT��
eBъ�R���K�ED�ԥR�(`��DJJDDc�U��DQPDV"�҈T�ʊ,Il(T����ERꚢR�Ԥ��V�Ny�{��Ʋ�V#�33wt~�l4�t���ФI��������m��d��y��YDH��)�ܫ>G��']\���l؃����ІO1����<[4��w���0UC{�Uo�S���Y3d��o�Hjp8Q���I�
��ȴZ>ϲ\�+� ���,%Q���Z���Jg�Ȏ��wH������aE*B�ff��'�wj���yU,;#
~ˆ�ڴ_���&߱&7* W�欿m5eSz �Mo�p�6��̽Ԉ�?���^ێ��9�VNfڑ�Qb�����]�L�%�١��w���K�n�,+�+��H��j��s��L�b��d�Uߵ�rQ�.�U��	�E��.�b�u��=�m�y*򖀯V�C�}���s����&o�e�E��e`J�_�V��WK���� ��k�Hq�&�����wh.fٙ��7�v^�/*��V(�!��{t�[b��Q�ݩ��=D�ϋ��U��\���/_��]�w͘��۹���:�[/<�Qm���LQ�A���]m�eK���>��x=|��[�ܕ�G	NMXc��M��I�]�w������W���|&;���?�ZO�X�������̩Hҳ����9s��/U2�g���ƻ�K�oǣk;��xJ���:_ozkBq��/ٝ�(�m����}���bgϯV���*�՛��m/*�'\�	V���eA�k�~�9�ܳ�N��|� �#jQ>���pϰE|�F������ʺex��_�+�^���/��L]3 ���ˈ���6)q����o<㻪P�}1x�~��P�j�x�z/I�G��w������ �5El���g�ʡX%�E�,��\g�g��~!�(�ޟǈ�90Ż��&!��E�9J�������ϊ���9���������΍�ó���/�2��a��Q�[�g:0�j|68�"\w}����>s��ں��+BÂd
��VL�O`�%�q`�kqhif�A�Wʳ��Lv�6����P��ھ�̈́��E��2����7��^;�`�0Xfα5Y�2$�gw���Y�]L�ЩJ����l�C]�)�A*��PqK���[�i+u��������{���[C/A�Zs��+�q�<@]RI�K	D�ue��iX���	��r�f�BId��C�����ݘ�"���UX�����)Ywe�JB�b��]�V-����AR"v��ER҅����e]�j��R���1i(ZJ�@�)E4�U%ZJTDТP Ѣ�H?跰��ޮz����{ߠ�}�v.Ǎ[mO��Z��N.�Qj�ߒ,U&O���"�.d�zn�t�qez��V��l��1y����ٹK�8�r��!Lг�]�����p{#N��g\��*�&sm+���$�6�́vf�id罙\�����j�-qRo�����g5�=�#��n�`�gm���u*s޼R�ԛJ���A C�/M[ԅw*�bm
{�j��T�cΥlT�6�rxR�w��^�U�`��Ѵ�`�a�(�Y�:Cӻ��$5���bw��כ�S��52������~���gp�טC{�E���[���������U�D�[厪_��.GH}}����n����R1��b]�gm4�=m�d��h�m8�{,�AH�(2Xr"�����o^�V.��2]�/[����4��Ǽk��,��L�=f�1%"� w>�td�<�C(���Ȩ����͝p�|ǈ4��VTP��Z��e�0�X���~������ݮdm�[gC2�C������&�������p~yXT,��,8�oҺ��f`��y�ly���m,�u��ޘ=�V����N�*��fz��n�}�$�b̊���Q�;�R�D�]����
7V�:��d�6�r�z��ݽ�j������ G,�iqw�f�w����Ջ�k����r*.�Ò�&׻�(y�9���+"�a�kۣU���yV�^��^�E]�]jyoe��n˜�7�����w�g��YZ�-�[~z4kvM�M�y����V�J;��ݦ�e��7�^ SRJ#j��'^e�_sW]<.��`a�1 6��m�8�,�\���F����Ǭ�V
��%�ٚ붽����ɚR)��%]���G0T����/3�GxI���nT�ëdcl�7��rbۧ�ĮN��p�O��a�=j�&=�B�n�Rk��Mc���ѓ*��0ɗ���&�&���ow,���-]Z���+^r4 7��kN��nI��}��{�Y����=@�pXML���8r�y�\����g'o��V�XX�k4 B]:�Y�a Ay��yV�2j�� ����t�2.��}7YS��O���j�����IJR�MUQMUՖUR%U#T!KBơESt]�IB4�l�TQcJU5UeUƊ*���˱���K�YWCV�%QTū�)�TSiIZ,R���MTJ�^C2��%R) ��Ҝ��Z{��X=���2кz����-�NnCZT��\��n�;�sY�}B��>��h��v��*�i�Y~m<���+�@R�}ۉ���҉��=��D	�#CF�Qû����K,*|n�����'���Z�|�Z�h%`}ضuz�Ů��O����K��Y��n�#�`sn.WC$�"��gn���9��`BV�"��d�U\��4��c8�iiL�ti1��YU4�2�a5�W14�,ޫ.��.������Lh���X�<��x��m��O*fr�Z)CU�X��_�۝��';�CL�i ��Y��m�3X�[M9ë��m&�6�L�C�o��C<�i��2�'5�:z���N'�Q�QL+��VgN��
�6�m5���3�	�2Һ��;����m�u:a��MYf�/L�P��9���]ެP�{l�+tp$'��C�t����}ۆ�8�2�F�`e�yEr���PM���r��IhkTe�.�v�H,�V^&]4�I�Ґ)Vs۞�&sS[(�$�&��ۮ��;��@޹�go1@� [�]�C�X�&9AG+(cU����-���fi�P��u���ڡ��r�]�i�*F� |fw�fwf��'Y���n��Kgl�N��zރ��:x�x�3��ko]V���ɤ�ы�[;��1l�m
zKgH[�=��M e%�I|������z@��V(���;��8��Af�u���^���i����re;�)��abf4��h�\�^��V����F�=�����N;L�M"�����!L4��X�{p�L�[&�S3)ۇo{1�94ɆC-�ӝg�f�oI02ٖӳ�f�:L��c#4]i��	�%�.q��ᗾsN��8�ɔ���tu��*x�@��֚:r�:fa�(96��J�{�:kБP�N�Ί7��8;��M��%#���&ӎ�f;���3��P���7�i6��k�)���GNS��y�W1&��B�'[��$�Aa�Pg����KH��f��X2��0�3wZ�uS)L�u0�L�(u�-F>#�!U��h��z�<0?s{�.��Ok"�!�+4� G��6?��K�N�E��n�eON�+��f3GHS)�al�{���oL�	c+�_7��"uR�Xa�q�����m�%�nS+��9��5tZ�Y�Z��6�U�S-�MVv��hRJu�l����G���3��Z�S7ѹ�P�C<��X�� &h31	7����ˣ����x��M�nn��c��V�8��S)��<�����6��v̲�i��̳m0:i2�=&�R��:f��V-C(�GI��2��]��d�Mr��S��;fl4�o�DAPUQ�
�K2�W��I�bSF�7+%)p9��Tv�1C�����/pk%[��@�ñ��XR8�oVb���]�Z*__W`=��u�2��w[�P�[9d<����⨺w�vm���s�ې�o:�$��l`�b����Y6���e��m3nR�n�N̼A��r��mL2���M%��5�i��-����U����*9�0�/@�R�����jmh �3sq�������E�L'�r0��;˫���R4UU3L�X�iU�J���*��+��+H�"*�y���s|���QA��}��7��4;C��g=6U�M�Öm!��Zb��Mj�i�HSw�2Ʉ��NwGa��I��S��ۤΨY�r��2!�X��p�{ۀ���a�a3�o�t뎓L�����8ɚ����ZS�|�y/u4Պ"�E4~�߰��	y^����7EMs�q�l[` �s=�òxv�v>����Ƙa6��6"ä����܋������{Ã���0�ah�뮪�3�Yi�e�3l��[��6�i��fuN(��sF��V�=����fSUD)���u�汉�q���]�c�^���5c����u�T�떆?����Yr�.��Y�[����}.����Rj��p��e&XZ�-��z�c���a��7Y�L"�͍�HVjct�޷�m�Jن
kM8t�gm�K����B�L�4�U�t�n^2�l�U2���fRVji�p�um����#�(ՊC�{=��G�� �-�r�:h�1J��@��������Rt��˻0�n�SL(�����2RhAJ�lf7�5�M�@���V>�������W���h��&ʁh3L�,�]�R��:t����]R�0vc���?LeF%n�#f���7��v^	d��EL���cB�n��.�ݞ4�e�|�iV���4y�^xj��ڰ����w��XT�;u�ܪͧ�+��;�_rRγM	
� ~5�r�����%=�9P�kx�x�"��qz����B� � ����|�h�N>������ᆬ0��<K�Q��NѶ-*Zj��b �Ʌ��/�(\�`v,!�[+!�S���Q���nސ^����ó^�ȭ�S��C��^d;�aMG��y
���{�r�Hv�8,3@#��w�[[o�T<�0*�1���\�!^j߭�7�d[���O�-oj�|��LX<�y�� R���0�&'��h�ģ�{�1*�Z�hȇ}_�Z}Ȇ~�W;TӸ�Jg�^�2ǂR�+1EH�^o���f�ܩ�������E�&t�lg{y^��b��,��ر]� s�k�{�i0Km۹/�Z�����Ԥ^_���m�#��i�$}���7�G�Ym.��xN�*MS�{���R�yW"e���J�ƾ��1���q�լcAw2��S��J�jX���◱�U�Y��~c��V��o%9��Ƌ����؀�#ժ��LSf1�)�;�����Vѹ}��a�5J��	u���o$�҉���5c7�4�f"	k�᧐}�u��%u�e�AvbG �*�Ie��y��1�j~��x���Z	�P E� 4�sj(D!U�m� a�r^�'^wNƫd���p���4� W̚�E4QH����bT��U[��Q��(�-#E(��H[�x RVn- }Z���V��K�1�V|kz�vU�]�U�s`�1+�U缕��ﭰ������o3�O^l����ב��Q���k���VqjsQ�ib ��WWT��H�o!��#b���-�/�x9\���t�pxh�kUd�-[\������c�A��
�C�:��z<<v����$���K����y��1�;g��纺a';Ǟr��mKN&��CX�'��wg�����Y�]�5��T�o���.���|vŏ�a�L� x��:�K�O���Nٽ����������X�I�ģ�k=y��zTBziJ��\�L)��@U�)u��J��	s�ĸ6N6��&~w����m�����+�@Yx=^ ,�Z��ȣ�*[�/�eK�u��N<k<�������2&E�w�Yov�D����[�2W���{��=��X��4k�o�B����]]�W�<�&�w��-�D��5s���������e[�%����S�PȦ�fy�t^�w���c�꓅m����rijx��Y��4�
u�VN���^�mx���;�jo�y��y��L�.�g����U�棷�PV|(]�@���ا�x�=����S�$��;n�(��f�����#��Cv�y|L/ئ2���6)�0�w\݉��J�xQ�o��x흝(j�sw�Ջ/�j�aK�E��9]��.>����/�ķV�����-�^���{{�����%+���56�Z�lU�=�f_������3P�x0r9�sh/z�C׺�-�<��:�-�/�3*V���m���'v�v���*Լ͚��m��:U���OL�/�;��*�=!��*�]��7i~�c��#v꽔��_�ܯ����~����M"���*�		�>��!! }�l�:HH?D]�+veJ|�Qyg��d�r�50���6�#�
�K�p@+��l犒`0%uA�0��		��P_	6��_�����������x�?J�P�}�=���7��slޱ�f��\8:����o�BB@�Rw���y�|'�Pj���? d���?�2�,*K>s���>�|�0���Ib>�_�������{|� Q���?0>���?��@�^������-(��z{$̏$�ej��ŅW�z�z���=g�v����e�����"��=0�.�>뚰�h!! ~��\!�8U��$��Ϛ���[ɰ�̓�a�0x>�����h��W��Ğ��=%��������g�\��!��!��?,I?����������߬2�}�ʄ$$�3��O�u�3��E.�c��S��(4I���_A����'D?�|�o�W�>F������Q�HH�{؃ϳ�E��<|	�C�?�	�jDD @����BB@���ĉ�s���4'���G�W��3
!=`~�	 jh�Z�ǰ.X�������ɚ�&��|�A�1ã�&sM%D��Hj2\��P2�P�6`�9P��?��!! vX|}�������H�!�A����ܓ�?���ǳ������}�������T}��e������>���!���_��y9��f�		�|�z}2~����B�O��g��?��O�����ӄ�'g�%��rg�3$lO�|(��B�o���$���u��H}?�����tjs���|�BB@����=��z�po�{����I��=D?gj�u�vk��2�P}��A�dB@��$�/������?I����$$t���OH�A�w����GARpI��O���yI?T�e u܇^�G���"�(Hw�L� 