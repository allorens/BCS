BZh91AY&SY=%��_�`q���b� ?���bB�� �֫@�[1�*USi$���DJZ�*EHV�)MiA6j��t����ԋZ�QKn�*ݣ����ɶ� ik`�a(�i]���u�>p��I�=9�6ʭm���:P��uP��ږ�RD���0��X��Cm�l(�%�+NGW6�UM����ʶ�j���&�f	d���n-�3U��ak�;2�۳]�3Y�RfY$)�4R%b��5KF���[j��Y�fm��m�ݳj�I,au��m��-f�+���l�S���j(Ֆ��Ju�4ͭ�\   ���j���;�.��{���e�=�U�a6�n4Q�E]�t�D�+�Uh��ungUhWm]�Y�b��.���3�qMm�k5m�ʦ�^��U���  ��ꔐu]ԩJ������EH���*�L)�F:T�JR�K�)tԪ'��Ŵ��ޛ{ǏR�#���A���^���)UU=��	�����e"���   {'_R�EJ�yê
U)��s�f�*K��y�R��{�7"��B��*W�����R)W��
R�c��Ru�*�w�z�L�@[�jصB+j� �6�&���   =���P�ٯ����J�(+X:�R��mފ���5;���
����)S�t�
P����RQE*�w�Ξ� R��m�@�mJR�'�6e�U)�(�E���   �ϑ%*T����JT�`��{�J�5)JǮ�)\=�{ҺjR��Ѻ��%*Sr��EW��Ҫ�mRB��iw���+��)n��zR� ^݂=���V�B�kY%e��  6�ϕ)U6���d�9*R����v2���u�J�w����*�磺�J�i��y^zT�j]��T�J��8�v�Is�wJ�Hn��el�4jT�ҘF��o�  {��PU��z�a���*��B�){���"T�N����%JRu	�4�J�*n���
Lt�iK�����爒�*Ǟ{��ow�ؖ�#��%(�������  �| hu}p� �Y�k�� �v� W���\+@�7B�@{K� 	
�F�{��s�MbM�* l��3m�>   �� >�tpP�s��^�����]�h���U�V��n����zE{�+��Mv1C� �N���6�4��Vl|   �  گ_x 4��n� W�V:(h<��Ǡ�����Q�U��� ���p�T��T��
W�    �*J�� h� F�"��F)J*� hb  ���%*���      �~%*��@     ��������  ��  �IJLԄڌ�E<��Кi��4LO�������?��A���?�k��*������*�j�w�}�/�����������~?Xm����lm���6��61���������A���d��������������]����w��W��clm��w���d?�;�D��`�cm��7�}W�a;��`��!���Glo�X�m��`�����C�!��m��o��m�86� �lBlo�M�8��}	� }0B�Л`���	�lxv�xC B`�dq��}�B�����&60}0>����0c�v 1� ~c�1��1������lm�; }�m��l Bl`�0�;c}�81�86���Bo��І7���И����p�v��m��lv?�o����ǝ�|O����������x�yw��r|�5��i?.³�*h
�뽣/�?Q�Y��@-�o�H�l�vmL��>������#�|ZT��]��UEaVV�3FJ*PQ�xi��L`$�n��z�]�mjyy��)��7CHڌ<��9���o4s�{f�)�4ݾ�%��F��|�Nn�Hn��"��,2��Ұ��(�Ȼ�qk�~ыj�Ǔ1iԣ٫$M�P�vq��7����,������q��D������sv��cmk8Q/�J�J;n��.í͍�[d=��l�s5�ѷe'U�koH�$Y���q�Q�pdr}��ǹO2�����P����n�4���?C�t�9�Y6R�MV#N�����ڙDo[�� 2��ݝi��u�)���ˡQJ$S�e��MH1P��2��A:82�'Eɕj�KlP{.�H�Q�k �p�]��6鼚�Qؐ4�'p/��h�óM��"�j^6DĚرn-S+xe��`5��2��d�Y�Ro4+������(`ޮj�+��=�t[K� �V-8 _m����
���GCf���+*;�2/����քSÔ����-x/(3��_
a��U�$�NVImcˉ�W��1Q��/��u�m�唨���)%謭K-%�σ4	�ى����-Xc^�"�r�B�lr]�ߛ�Ŧl��Ano(�GK��[i�BlRTk\D��E{SF��x3K�M�ì�6ޣWV�����m���U��m]^%��k�b$m3���@�V�<K�O	o4��1���i�/q�����͠���L[I�i�z�
H�SS�G�hXNR�Y�a�wY����'�Ś��ec�R*7��%�{/��/6���l&��S*jF")Vr�A��t��Ji��
���FLѰ:��XN�s ���)f�^����p�1��j��C�X�]�/+e����4/4q\*��]�g�N�ᶱ�H�ݯ�`Fĩ͡`��;�S-M�������U�l�3)�m�q�(y�P푺e+[M�e٨��Ä
�-Z�CY�n�����û�uvB��w(7�R�MH�)�e�#f�r5��'���tX�R�V���$�3 ���ŵ.�@I+M�֪�=m���6�j��ְ8�-:Lj�o,S�9�u��(CT�]���F��BS���{���8�kY�7H��V�!�T��q_m�Au	`%��E��vs�ۉ!���	DRz�rgۥL"R�3qJФR�c�[�����ӊ�b�����"���D�ݰ�� �DJ�,����0�"�r�h��:� �)!\l#���D�	����S��2��+^�h�Sp�S�B��e�X�əX��ZL�����ӂ[�v�}�r��J�P���;�޵lr�b����wl�j�K90��K'�,���5���I�a����X G:oݦ�I�ɕ�mV�8��=y܈42���;�-VLB�ҟ<�W�]I�p:n��5�-�(<���W�M����ա���`�e��B��me	Y,$�ԃ\�W��yb���Ȩ�F�P�a����*���j�"�y��=���]����/6�iU�r
�X6��`۫3p�e,׫*�)�+��U��[�[� �+8��mJ�̦sPO�5ى��ңZA�����S�[���#6�ZW�͔,�Z��Ěϵ��5���w�!�si)gqm�;����q0�׫Y�ڳ��n�����^�t7�c���Q��g"y��j��RGOr�ŰE��C�����@���J���$��s+/�&�v���	�E��N���
Su��jz��Ւ�!�\Z��B���h������ޫ��U�t�Q�V������6Kx��-�!OY�,#~��r̙6*,�j�i�Hu� ��f��,�q�wneia]�P���1kJ��:ȴ���P`&C��KiZ@;j{`�a0�sq,����h�^d3
��B�N�t�v�V֋�nܸ�ܿ�.9z��m۰�n;.],ģ�u�$�ʺQ�T5������NpQk&mX$h7&�{�#��R��Q��ǭٸְ����[H�v�I���P�3`ub���r!���j&�7ϗ�t�eg��Y(�.�#3	hVL�v=[nܱXT#{��]�N��NҬ/r�����0"Dv�!��'u�k,i�[�؈@,҅�I
8R�0��-b{%+۬�4r��F��U�@I�؃	�a���#���l0֛J���n@U̬�Tл����CSu��-��Xi�Jɡv��2��ԴC�0� a�,G����Y�f5s��!�;nm�q�͡�V�eج��Dl�OA
Z�\!����ܧ��eZ{,^�V%R�ۆ��^���6�me���`����V%sl�$�Y�����wm��3U鲵#X�El

�6�^�R�Ji	Y���SB�����2�S>�j���"��AjT�ɖS]���'�!��"ir�Ͳ��R���f���<YKv�(��M��*�L�,�sT,�b�ڛc)c�4�Ģ��:o6�(1"O�.�kw�j+������ċ21s�"�5Ah���:P`:� M4%^���" �i�X�:���=�i���J�5vO�0iS�0v*[7blQ0��M�2h��읚�3x1U�;2��e@&�[ur;5�X/Q���]f	IMŰ��Yu�Q��b~g-,����P{>6U��`�����J��T̚�tqA�EM^d�&�f-goF����
f��
�%5+$����f���b:����c1K�L%��J;���:(��qL��xwX��1�~M��M.;/���v����)�T0A0j�^9c&.�؛�"W �22�j!	��hcǢ:vIל�%J�6�+�e�#�śԲ�R�m-t��&��B@��Ay��z�;�CbMTKB�@q�f�v��0RC��g�	���=İ*�QZp�Ś3� mU����Gr�S�Q��N�I!�q)����yXrl$̛xv�VV��Q��̓u#�&#�1�4�fH8u!�S�-�����-�v\�]͠��]�N�J�én�!�6�)���U]m�H��=�4\I^�� (9$MH�W}5uj%e�EP��:��"�P���%4�-f��jb��O���ڃ)6�����hZ0ڲ7E�a�_X�v��]������U˭��tc3	�����CF]rYgpǱd���V�v�V�k^nG��L9`)j�lj�V�w�LfT�7���y�6K$�."�6�B�e�	�$��2$ؔq9&E7,��2��e꺒FEiy�pV�K1�A��d����5�;�ub���c}�z�t�����{��ʦ�:�7�Z�bٶ13(��$�P�;f^�
FV���yu�%�Ѵ.�h�c=�"�z��*�`dI+�!���S����Wb�|�T歨��C��Uؔ+�a��n��P�To#�g&�S]�Xo��̻�.;4&5�,����
�5n�w��ޔۤ�3RЦ�4X��a1[�����XQP�]f�VE�.�q2m�N+��B�P8�SD,p��[sUeg�ҕ�@�p�,HrbYO3F��gу�֑lc�mhʵW"ڽ��G3���m(���x�n��B.�l`�r�I��婁
f��,{��'Aծ���!n�2�|���x	������@�ڹ+���c6;�]eEt�՝�LEn��2�z���.�m��وM$�Z�Jwu*�J��k�'�n�c3�V��¸Q&�7\�Tt���	�Vjۭ���2hMs^��"���^<� 5�:�ѕD�]]%��<ۉ�%�]#[��u{��0��u�J�R���>$&��K��q+!��0���I]e'J�S������Ƭ��i�#�$�(��I؎&�'6�l(m�#�*{e��p(wXU%G[��x�ڳud�Hl�Z�o����
�X�A���k*n�xH.���t����k~�c� �ȳ��
������
���bI��p*13`fc:�JՊ��K1]���[B�k@I,�m�`$.�,�U��5����Ff���UL�,5Iˋh�YB���E�+""#z����@`y{pm��-b��&r)Q�Vf�Yk+1#�e�r�kw,j1���&5.a���6^5V��
�,n�Dʛ����RKh�7� �P)��
3F��j�[Wq�n�aM�
#'��h_�MW��J��U��
��[(j�k5C�ӌEm��V�gf�1bmI86�7�.�#9W�� 9I�À�vwYI�dإU�|�5E��yz#e�.ι���5"��e�f���5�Km�fږY*��]&V�B��P�q���m�/���;JFF�AU����d@㛬Q�L���l@�;Wx��R�[Z��a��S\�sy�-4�>��?i4��{*H7e�Ӓ���
0��
��NY4�rr��Scf�]�
�\ɸ�NM�zf9�#{r,I14Kr坫�FPH8�t��!u���ܙ���Z�En$�ϥ(qh�E?�H 54j�j���[	M�4�ll�F�ڼ�65[�2�:�����1
�;�JsFJ�+&���)[N�5j��ܖ(��^n�"Xv�Q\2�k,lw3,��1�5���ڬ %Sr,����ܓjR3��B�2q6��8�a:���d��'*���"�w�10����)��H�I�k��wt-���B�w�;����KV��Y��4��Z��.ܻ��p�(G�5�j&��c/7��$�����/���D�<�����nU>o*�$��cwI,V��&���Č��ř��k��ݒ���#Y5f�v@x%F�BX]ix�m��b#hI�GZt�Ç_�� xf�8�I���Ђ�n�X���!��d��^����L�H� :�Zq��Y�����6um,W4K,^�f�HY �7t�E%z\N�����X�*�LP����#���t���<6\� [�u�i9�v�f�����k�ǀ5�2�bEm��2����h���9�ݦ�����nEBZ/k)>w7��?զE���Z�A�ɒ�
;6����K��ڻ�3aۦ��d�C!�V#�S���s�|j����*�yZx�Ma�Wuo:��Ёܵ�谳�$��:*˲uc�^���Hڊ�Se�ot��a�f��%�M�-8��!-Q���3a[sp\Ů�i@�i���F�R���z�6va��f�Y���N!+6�#�D�ն,�
�T�`tv�N�뤲�+E
�K��l�U0(a9xUlqTwQ1�hU�X�W�{O6m:�j�y�mZ��P*'(��f;q ڐ�q�ϐޕ!b���;t[��Ҩe�]3�K��U��^��@'���e@���(�����lC-�M�����,͊���u�H"+BVD���q� VL)o�mC�]ݭ#�b�v���j�2�K�j�,h66U��sF���T�	-X�D�.\�%����.��wiP�I�#{���Z��B����J4�x��;��2MփH�>����Q�ze�ǔZ��c�,AY�[�3ˡ�&j��q�ʚ*;Wz.�����)�Id|X�ʚ�d
ỡ��+l���q��G�xV�;G�u-Z;��M�&hT�$�A�Ʀ(����X��,�e�v���Le����p��y���Xce�n�fV]8 ��ըA`��i0�o4I�s�N��!m��DU�B�S	 ���^�U�^m�Ϡ�a[V[X�I��G�ˡ�N�Y$j�f��8��i�`1t�çn����VN<ss]���N�lZ�n��2����AR�[F=�Ӓ����H�7����U�1�2f3B2�d�2����e,�K*�	�����֭�{��-Ҁ�L�Q�V���I��!���m;�a�iD�᫵/S�V)m?�c��K�3���:�TVB�
�M-ML�%eb:Ve����_R���7��ݻ
I��%�H��֓*
��Zn���()@)B7���#1��6�А�.���D��L���5&��6 ���0Ve��mRxw�Z#ͭ�X�(m���ǳ����Fŭ�`��&,��`�nk��'!ڼ��h�9&z�+R�R�L�]�X]��.�)*���v�"ʢ�d����R5Zm�w�[�[�͗�P4b����[2�027Qot��#���p� �Yf=$+�fK���/&'(��u�uk�#	�D^�%�u]��k"Q`�jՓUh����6���`�ۦ]�%����XHIϲ����/D�U�J�8V�Z���!*��9b�:hf;ٴ�Z�Q�;OvT�t2K�QR�ȭ�ݱm�R�A֋�&o�&7-���v�E�-��Y��bzLz�è�E�^�qS��-����YX,��nP�0*ۖ&�xj�J�繽I�_��V��:^"��#:�3yN����FS��@$ّ^�$���nZX١Ĭ��Q��mL,;ӹ�KYG+LU�/iJ��cX{�%GB�6��)	�)H ��ee2�(�v/1�1�֫q�2�%Z�:Ux $V��n��#T��U��(M��ƞ,O�Ӭ�d�,�I�C#"�B�
8�"(�n���+�3!{q�2��S>�F�<�`�N@(��ʹR-ŀf�JpqG����(�[�#Ȇ���X���%���7ٌ[Eh촳
H&U4�<Y�ir�n�R�mԆ�Sh@�1z���ni�m��ъ��sIj����J��2T�����/��^=ĳMn�r��M̙�nS�$�r�؃�2/��N�eE������;MF�QQݴ�n�R��1�ۛz����$p˷O%{5�C�����Z�uB�d�;��0�^hj���܉�9R?��~��,+�����(��ѯ�}{�gsV�`���[ӑ���̌�܄Ms�<~��:��	\Z��k���OJ[�rܵG7z0)�d�gU�{t�+ɜ;�Mה���� �>9�8��07{�k�9���jd��):�b�`�(qP����i��eN��Y��SjR`32�CC,����wnv`�E�A���<�N�����+-�Pz��ȣܕ|�虴oҩ[�(F�����R���g��../z�˫�>�/�:M2�S�\Ný����%��3G��t�V�-�A�lp[�r�f`<��X�|�]�t��ˬF\����{�)���mJ�F<1J(���Ÿ����u	��;)��3�AQ%]�����eXT�P��ԭ�=r��hk�䎭E�ŗ�v�m:
���Y+
�� �o5>ʵ9�s�Pޫ9.\�(b��[@ �Tb�9�9�V6ٕ��� rf�L�Wn�e��3 ��.8T�Zi��":ټj!&�����g8���J�)�ܧp�G ՗)�jt�!��q�a%�m�?���6c�oFKɨ��Z��#[8]�{{}�9X�I��cͬvp��AHΈ��f:�u�旛��������8�����W��0P���a ��r�e7=*�V�����k��8���g��H��<:P��#�Fhy�r�����i]ػ����(9̹s(:�=�<zlbu;��v�œ�q�Їv��!�r�}faJ�WD�E��P��u1fр�*i�:ی�K�[I��u$4�s��Œ3�b$9
Ġհ�u)<�b1,c&L��Ń�zV��L�����oq�uѺ��2%��ޔ�Q����bp=����3�F&��M꡸�m${��3�y�ru�F�KV���,��	�	8� �-I�j���[l�kG���;�R&���Nܛ�gj5F���.������D3��f�)b}w|�Jua���.�ɸ��}Ժ��Qh�7^Lǳ�C���6v��v�ciЃP��U+��ӱ��wn���em���0Nޥv!*t9�5��q�����i�-�W�����!�\�M�:˔�ބb%c�3[腸<�����H��1�j�v�v�e97x!�eO���:�7�(�E]�����5�fl��l�n�lW�V��[��+掋��q�#*�I5�Z.��w�	u� =�E
�Y;�W�[u{k^��roP���n�cE����`b�SS�M�=�V��#~��,�S=w�|)������ŷ��\��B3����[]��ai���z�(�H����!��(�f����8����s��?
���{�c»V�]?KpW�G�X�C&wT���<�<U;��)��+}�gt�����i�rH��!;���^]`㸷�uװ��863)���Y��鼡��ڈ��d>ȷ{N�ʺE=8XW��U�#�҇|��g�`�Z��ʑ����u�V[��wWT�`Q���B��Y7ɋ���5@g�:�����%�b����m�/�X@��ٵ�sL�Sr���g5�0)��v+Uk*�
'6g%]Y��(��Y��:P�?u�i������]�<
���Q�+�U�*VϜ�^�^��	�Ý�ӝbD_|:�YL��麩^b0w�W-�{J�9�]�j��7]5����̮���"�.CÓ9� V�[[�ή�F��5L�<� �D�!���<�V+�!�.�
.P��æ�����IdN��f���J���V��0�ɳ�k��͊��P	Z�]+���Jj·F����+��]++fj�Fc�5,Z&�%n靮�n�D�@��2oP��]�j�0lq�6��-��Tu��)5h�S�ꪨ��n t���Ypֶr�Q�k]� �V�
�[<��Qe��R��o,���H�~ˤ�iݵ8Wj��-��.4���=Gj�cTͺϹR�2NY͝�U�]�Y �7yV��&w�Ь�]#�
�ѕk����N�hi]����BU�3 }М�s���
:��h�~\�s5q�gy:�>�N�h�2V����l�t҄��	�̛n
w�SpE�c�f�L��dò3Θ�엃�h�'�BM�nG˝�퇪��_-������Dz�5Y��q����Ij��J���n�a����c�og%Qłț�S�N����]]3:���'OT��?��!F""[/�ޔ�ӫM��e�\��54��H�̼�Zޠ�u�]y���l'f\ؒ�wl�`��)΋���Wt͒�-M"�Z�=����ΰ_�Ѷ�<�f�y8���5gix*a�y�pt�'{m�t(���a
D7�mc�S̺��z��
�#���-ޑ��۟p����cO�9΍�֍U�b7�h���s4y�x��
�8X�EWk��M��#�h�eGy΋�.mM�6aXV�����L�a�bsY�7B��ǷN\:���V4�*t�ʽE\��}6-$����?�F�.&��j���ca�(nVp{R�.yw�[��e�仴!\��#I=��C�oE�C�o��@Mެ�l�ҫi��1�Q��<�9�_#�=�ާ���u����u-����8��M�Nѹ�N��1�R���#�O{v�*AMۧ���QfE�k)gcE�a��;
y����7AA;����Ss�b����W?�2t�(]5��@�X��ZOkA�J��0_iyܾ;�U��ܝ9	��U.�ڳ4\�ӍuR@��q5���y�eGs���nvК���|��S��wpv�	ٵ�t|qᤣ�n���yZh��ƺ��h�5��|u�K�V^����b�X��A���W5��ogl����K+���N���5���)�o�����{`.���OX����̻��x��u�t�u���0�c����I�Q��ˬD
v�f�.B\�� Zɮy��2�i��\*�ÓE!�3��Ȩ�K��n�X��1u�7�/�Х3�%�(�hM+�:=�;�����+�M���D��+��F1uw���Ѥy��&��:h^=234��s�g��CV���gp�L�E�x;�ᛉ�����%���2c�zf3��'��Թ����"�W7u�vRGW�J}w������{�-�	'[�t�7�ے_3�l�=g �\�:r��!���g3�i�s���y�ZEi�6w��V�%�/$��Ҟ2�\��a��_i�����e&J ��"Н���w�c�׭V�P���L\�VV��W���)Y9�����J��U��\7N�X��+�2�۝v�I�B�x%r�z_P\�R�%@m�#��bY:�-tq0D�L�uf������rHC&
���� R�iI��웒�`���gk�;͗�[l�1>��H\w�>�ut��VM�]�w�<�;��J��F�	.���j&E�rݮ��tOhP uāVั����w(w��J�mDRV��A,7u�4'�U���
<��uz�MAN�*,%۽T��V�ܠM�(9C��A��3G��I۶�դV`�
�F�n�����ޝZ�Os�״��;m:�n���ș}rnn�����Zjf4��M��p7 �Li��*����I����^L�m*#�J�]X��G��|3H���U��"�h�D�Al �$�fp���Ϋ6hM�Hr���dچ�l�Y��NH4fL�ٻXA5XvtAw��E+����X�v��������!]y�_J�)�o�փ]������H�����)�0Z�W��S
���Ә+jfN�,��ø@��F�Y�Gfr]хY�1�5��1u��������������v-����W�kYnVL�ۑ���rԠ�A�L<80�&u�o�U��4.�,�.�� ʤ��l�Ykޮ�ׯ$��r���Ϫ��Z�yس&�݋�=�^|��;;*b��'�MJT@{!��\��@�D%]��NC�mf͕����)�E���SV����2D#&�Ⱦ��0�}�bzr��WS�J�s]էL<�(+'5c�J��������w��v�J�qkE��)u�H�y�}���@��J=�h*.���鳺�^��9�|j�TF�1�0^5��FU��i�sP0�Yz�~<&cW��R����.����
6�o*79��i�[.�%��sU0�4����n��/�����(Kb[-�Z`��B��y�%p��
�芳����h�.�r	bYڷWT�z��&�:�m��lUyDR�Ē�vY���ؐ���>��u�D���A��f�6��r��p�y3s3U+�y�&񡸫o�=K���ub�v���1�e�|�m8�[Qh2"�L�{�v觭|���Q��S�>� R���&�I3�p̼}h�]����Eq��qpO��{�zK.�tΨ4<�.�j|2��E]#n��-��62�]y��:�L莺J8o��`�k�gp�n� 	���渧@�m�pfp=I�V9d
����q�i/�&�u7]f��R��eW[A�Ȝ��5m]ra( +��הO����Ds:�tj�3}�À�o��@�s�&�,l��5�(NvJ�M}�����]���6#%��>�:����f�n�=N�4��Sn��(��i���&�s�����8/i�Ӯ�Cw,ܨ.�t�"�2�H�=��I[�^;�I���K�wr`i}������m��H�'[�����6�5o:�RW�Q���<�_nW��b�
�^>&�pX�I\�gi�t�̛�j÷�b-��<�"����G(1*ȶ�#.�:����͔͋6n	3-H�nV�[Pe�4V5�u3Ur�V"�L:��uդV��i)���o�:���O�t����%�h�� �sp�b���R䶲��6qbuk�n�nǮ�b�9���.6��j\y���Tt�^<�[�;=�f=�\b���e[�v�e��6Mv�
��'[���R�S��C=�G�Ǖ!�vŔ��#7س���y+c�YIA�s,\�5�$'����˻�-CY�4���[�]-����1���35��h��c�6[�ѹ�Eܒ�lG7K�/�J���0���m����]2�P��|tn�.u�CjB�l�,\��V�d�M�6��c��-�N���)�X����Հιү9�yb=K��8��f���Q[�f�J'6��#J������2Ӱ�Wn.2)[�[�B��Muim	�E���z��~�p*�jJ��;�����3���&��F0:��(�@�����C-T�rv��g��M�-���b���;mUq/,�<���\��֜�\�VK�ee�,HN$��b��V-=Ԙf�nK���4�lsXy#ע�(;2��:تh��ݳY.�t��r��.����������]�Uy�����V�[�;:I;�+oS�>hwh�B�ۊ�{�Bc���\2�#u������Z������7I�a�J��,v��k����E�fa���-&��+2k�s�4:��BM���O.���n�K�����-D�S��ܺ��m�}sV�iu�P��Jӛ%ê�n��9k��i�n�8�	��2&M��A��)��Ę�4�WV,7ưY�k�����<��D�����	J�B�Y��6��ճ|��o���=���RWSF��R�Ʊƪ�I��62��gu�2�=�z��sVk����f��*��1o1��hǊmK������L��!|�;��MMK� ��RyX�mxX�;[�J��%�hMx;s2����3.�GY6�\ZH˩�3d��w��U�5��*+��Ч�l�2��|�4Y���o\|-�Ʈ�\�t{w���CС�������eYY��-z-�׃��ܹs�=�+e��{\���mu0*֌�s��ms[����Mn�¶��E��=�b���ɐu�4mGG��*8VL�3,��d����%��["ꊚ��1[�c9m���x�6��>���w�8n�s�ׇ���S�t��∌i<��e�
��BF���:�M�N�6�H'}��m���pLP.&5u�4��%7�I��:��3t#ס���n��r����t�p�qJ6'dP5ӨZ�p�kM��&������bWk��5�¯ ��WV�.��+���wQU9ǣ�v�Ԫ<��J���X�8�VٙS�����p��b�F�d��fD����?Nu�%%�4���*n^���ى��)y��������9ua�j2G3)�b��2�M���twr���٦�Ew݋Jdjm��͊"��#ͼqX�Vf\���(�!};�w6�k�gwLt1u�te��=��O��W4�L���*f����b�׊�t����j���5����l��R�V�2Q[�-փ��h#Z�Wc0��h�q���h�o&f���iФa�1AÅ�Ўu>@
2�o*;���eH��]7g*eHju���dY��qt�r3>�V��h�)�m"�;��8(�����qgLZr��b+�+��.�)$�ӈ��7�
�4�u�s��#�ɮ�/d		��.Q���hunꖥf;���̙o{�֚ފP�ALP��!����iH�d3t�tyry�V�WY�
W[��Pc�U�.(x�9.�t�ҧ �j���x�E���yL����� ,���n�ɻr�����j�sVcB֌fEc!�̶>�Φy�5�U�@,��F�`qVƠ����:�B�L��ޮy�:�݇xg�(.�SQ���᫘����YJ�c�a(_J��`]	+u$g�QTz�\Q�ä�w�e���v���#�A�^�$����6���|�H �ǒܽ?K !��E�R7���u5[')���;u�2P�pWp��r�j�@z-�2�Q'�o
�N��J��4��w��W'��wݠ��w���\��P���G"(������^7�;b���=Q䭟[�*����X\"�%ju%�+��T�٦�i�˽�����9���-�з�O�b钕�Ť�T*�f���p���f��T�J��+�2� �n�� �r�+%��\��c�~��_���m���W������O�~��cm���������������q�o����}����3��-�����2����O�sgge֜�v���r���q��κ�!E�L�O.VL�҄I�1�/eK�J*�:Wͨ�x�0�K:���`V�9���L�Q�J���En�A���r��5!o����Z+����:�@��9��(A���0"ݒ��m�b�¼Z��4�P�m�#��N�U���w1�wQ�a)]�c
f7`�`��-+��,,(+�Y�PJ�\˳;�[y�rtI� :2�Gu�Q6[�M�] N��-�]l6v���i�2�L�WV1�H�ՙ�U��7��@�Go�9�d�6�L�	D�gr�w��`X6r X"�0�e�R����.�f+���Ïx�Z���^�VrV�	�3����T�U-���0w��U����1[��!k�V�)d-I�ٵ-!H�SN��t8:m�8����� �#�7�(f��;�1o]p����i�8Xu�L�+R��lEM������56U�1.�3y҇u���󚯅V�����p;jfv���uYz�o޼oS�� 7�8͘$�K�]ni�-���S�df�*yk�]� 9$��zݍgU�ީ�3�UE�3�5,:�{�G6tc ��D�̒-�%ST��l9SVu�EuԕI|�j�kM&L9R����Y���Y��-`f�<Z�.�W��moA�酷K%�ۓ*m��2er��v��G�]s�j+�vrVI:�VX�U��C]Oj�[ג����'i�����D�ݡ�4�:��-�9��ugN���㘎s�m:nc��W��Q��uPe9�:��VJʐ�<-Y�*��݋�x��\p5�W>�ME�[���U9:�!wVAm*�W�B���` �g �syX�f|�X� �]��5{�]2��o-�e��1ݒRR�V��v^�{��s�[��h�i��5�&�kҌ�NoF�K6��ȴ�E7���:�dꝅ���{z$.6�,���)��ڬ0Jb�16;�)�s���v��o��}�UЈ�k��3v�T[*��e�p�et:�֤Х��aT�[%�2+mwJ*�3vw�b�mD̲E`S�ʐ��E`�:�*��u�*;�t����)fL/�����Ӳ���h��+��k�D���Y/���{��
�U�iQ�j`�cV����F���&��8�1tDdI�A��o:Pߘ�a�h���x��w-B�d��F�K��M�{�
�1�c[e�@���@�鲰?-�e�Ԫ(;A�N�&L��v�.�,5q+��Y�{�|8�k*C��9a"�.�pf��J}g�xt*"�8���`&�O�v�w�'O�t"��!n��2hb�Ŷ�q>��մ�/�����\j�W�>7M�c���=}�Jh�j��d*�kev�]��gltA�**N�u9�^�O3�h����ԋ����^Y�:����݅�2J��y%�X0i8gn3�� @�K���m�R�)L�Gs[�J��)cMe�4�"�_5��خ�YB3J�uZ�na�&e�[Q	M5ք�b��U ���]:�gg5��k�b�?0y���[IM-����D��C��ֹ�7�'��g�(�����#�r�S]�S˰�@���v+�
ѸeÔ.bɵtT<K�N{lgIsjE�M�4��c=�vYcN����6�w91�w0S{�I�u�r��T�@����94�vĚ��ˌ�y+���gf��If��V���mWj����nC���k:v�������gj+}��}�_r40�j�d���Bc{�Qv1��x�����*djYW��d��sΉY��*t� ĲP��&]Ⱥ��B�Ù)P�5�`�,�J�:�m+/�h�ͮ��wBjF���8�*X�|;G9��G���r�͝%f��hR���ބ�����T�"�:�����W2�5X�ù�y�$�J�Fi�=���Fj�Ƶ���;�2e8Jt��#�!�Lnl��vP�+�ܩ��l������u������� 
]��?��qE���
P+;Uw�<�h���K��a�a�Z6����2�V�ȝj|����>�B^�u�&6���x�5�M�I'���/Q�3jR�.GD[<Qi�TI�(]�=r����y8èV���|�%�s����g���Yz7.:�T���A�$��ú�Z������KѴ�r��K@�}a�:f��a�B(0��Ƌ����6��2����򛦵��>Tq��C%!hY�}.[�hޑ��˺���c��&|V1�rg�ũ�5#d�=D!�4r�� �q�R��(�Z�N8ZV1ol�J��s[ZwS�y.��
��."�Cy_۬rt�l�d"�i���\�7;�5�ƇKغZ�n^���y��D����$Fvë3z`=FnlW�.}� cE���Q-�M�Rʝ'J$T�:����=	X��[#:�<� F��5z��k��/I���33LL.:���VR��`�iT==OX��!Q�b��\ʿ���N���z4��t���o22�����!�-�2�7do���{�u7�̢Y/a�|:j���t�����[Xh*���//�7a�^d�P�TZ�ݓ�[i��j���n�����f�ұpq������1N�Y��*��ƀ��g0��^�sxsDx��e�'R�ʴ.R {l�)R�\�`��쿆bd�#��UhQ�J���Pº����s�6���-s�DV�0����K������H���dw}G�'��f2 7@��A���Fs�^A�K!<�zĥkl�wXW��+�".˨���	f���Օ�9�6��\�=O�ma�Ow;\T����1\�o+��u���CLXP;��`���M��Nw)&�,�ݤ���ƙ���x�de3@�F��%� Vͩ�J��(�5�C�Vj�o:p�c!�
�v�4]Ĵ`��9�Զ�Q/�ǌ�­2�eԫ9�ݽQ:̲;�wĔ��r�7*@��ô���UiJ���	q7�ž�Y��Y��(@��w
��c�R'�*'d嗥��x�L�S�glWk���Eh�c8�����+OQ��,栳2��LVr�%l�� �D9��f��i���ͱ�.�(��ڹ:����˙�/-gq_�(�,���9J�3Cʷ5ڤ�s67��I�6�8XK�(%[�\]��UoV��.j��mH4d�`Z�[%�M�c���K�����خjѦ8�!�)����Er�&%���W,��I��j�
 ��
�etGu8۳�yEM�]��p��i_;H*\�yW>��%ۤONA�t{-�F��H-������rp���3qu1[Y�m�ړTs8��Zd��sCD|
Ü�p�϶�c(8΄�Tq��H�{�N��֩��6j[�T�������i�ܥ���'��
�D���L�������Q����trb9@K��Q6n-��P�͹���Vc�ݭ�2�[��H��`�1ۃv��Z]G!�6G(��B�5����b���;��;c��Ӫ��R�E��vw���*	SN,$%n��R9{�mN�mռ�ˏ��+�w����1O��i9ՔY���1��.�!�o�X�F� ��,�
����<:��n�ܧ.��Zz��u־t��d�'VG�h|B�:��5�btoD�����Vj�#ߕi���w9k/���A���f��i�M�E���ը��L�2�qod7��pj�5/vk7�hV�F��mD�!�j_\�_U�՜���`Z�w�����Ve��Ө������HD��t϶e.�+_>}�a80�2〩�q_f=�H1��׶͋�)�O&�˺�d9��5ϣ��lsuC�VX8J�}7I2�8��sk9��f��x����7AF®6rSǳEc|�֍k욶��%��]A9s�贊��Fh��[4S��C���|j=��]��Ѥ&twr�Y��@k�mE[Wg�Q��os�j��o�81����[�5Պ��,�ܫK
['�Í�7V�F ���+����]7A� y�8�k����9(A]�곒���S����.�jy3��{����(�ʊ�ث�\��D͏{��ţ��b�l���ՖRM�����q�{�e�ϖM����9|6�L�a=�� {*�/�lкj�q��56��6u����F�r����pV���|�82�j�Pu�W(Ho'j��cQ�H}�ޮ�3��p��I�P�;B�t��o�a���:�(����]ZS�t��|��t��$�����n�Dڼ�@'�+ܧZ�l�Rԩ����A���.��Wd��u�	����ڕy,`�AΈ�J�*���K��~�CSX1��6!Xj�95Z؜�F�2�i��맖L=X�^�)Q[)d��o"��Y��$i}���JB�f=w{2V !���*�:�8�og'B�|�����GbMy�e^�f��y�(!���Zb42����"�n4s�W!�f1ҧǦj.��إ���c���EsѦ�k&�b��"��*pٻ� �K��.��z����X�䋳��ٖ>���lӜ5Ɋ�%���rh�$��tjA���\��bl U�S0���ξ���d��V���U�7;o���0�v�򠳺(�Va��+���W�����@n�ɩ�-;�&���
'zs�:�j���en*�6������7y�3D�+D�7�nF+�X��VH8�4W�R�5V�����{&�ܷuX%�3+�՘�]%L(Ye^%�h꽬cao/%���>�K�N����3���B��5w�s���=�Uw�PZĥ���ڋHX�%�1 �:Ke��B�Вmŕ�(�J�� �K�R�>3J��,w�vnc��H�"�|V$��K�t�l�\Tr�����5�5/)�^K�m+��2J%��j�s�ě��}���D�wg6�Ucf��ͻ-�r�<�*��/KR�����Vj�4ŭ�M=��gA2�e�l���N3���C<���`�T0�HR�H��Sx��U�q"^�;�V������K{j<�ӂ�z�l%�X*�&Fe�U�Ay,K�A��m�5�E�Neu6*�%�0�mXٔ� F�T�ެO�Ͱ!���r#S�A�j���U�8�颥Ѕ�;##A��`������4:�u+���@�����F����;ܚ#
�qMeǑ [��`�)�-e>�QjY�7hM�m���!�A��� ڋ+�t��",v���J��%5.%�heќ+	�F���/j4��-,�Q�d�Σ��Ͱ y%��kX�)Û��%��Di&�Ө�Z�)8�����¾�H�%�!Ǩ���B��&��,b�aΨ�ՀT&��-�#P�]˅m����kG��n�bd�`�i�|�j��,��I�4˩l���U��;uvٝ��*��p�f���)��7d�[ct��b����H�_:�؁sR�̓��mJ��9-B�7�<���$f��D�2��xX��t7u;'���1�n#jN��{�S{Uvb��u:���n:/�3D�^�e=�5;�U�ȭ۲��Wd�l���-��3C/b�o�R@8����v�vV<´��pDq��1�a�$]�2��Ζ��4�#����N�kr�rW3n��M��D>��<{*�����S�����a�95k�� �W3��ku���ii��ښjL���њJ��1��/u0+�a)̝�wU�*dx*n���b��G���wY 9)�%_D�ˊ�8�]y�m��uy�_K�I�|�i�����c��pEr9C���h�c�v�$�(z����ΠD�x�R���j�d3���m褂ȷNĭV�|r�PY�7ve��)ћʐ�z����\i2�D�,*��N�
��s��s5��Y����_e>�ܹy�W2���举��&��= .ՁZ:�j�����b)ci��ר͛%t��xr3n�S����9�{(��0�i\+q�Lfob\ƨ-TZ�S�"]f�)f���W}�Xy�ǃ���Wu��?�b��X�4��{��}�2�E"�d��r�w5�r�6S�%�Y�'��xP�69�.v���e�sk��f,���� ύ
��S/6�pK�+��VRU�y���7v���|,���9�뗅SCS5���&�t\۫��i���Ʀ�\���Õ�Lk�ܼ��g��]v����K�]1��a�]A�{�T��@ZwWM�N�Z��`tkVV���VufJ饱�.��;'�!hܵg �c�2+�AY,�\ K�|��X�wN����I�r�b���+Saj\[����������7Dq�2�-���3�p�5�-˸!/�Q��y�A}�7z':�*�m[�*��ˎ���O8f�,��r�9uO��LІa0�S�mgΆ����m��!��&�0֋L�}��=�������W3��m>��(�1wâx#e��= J�n%��]�If�Щ��*�Ý%4���)Jͱy�P�EBXꕍ�9��BӃ��i"�8p�Q�oq��:����T��賂��j�DT� V�#�@�����R�7`�y����V�*��ۙ6��D��`���K(0t��^vev�z z���|ՠ��ܫNy�=��\/n��̓��6�ݪ�!k+]#l������,V���bLR�D��<��u�8yf��k�bB�>�G�uv�;��lX�&!{Gpve*®ւO�����Zp�0��Һ���]X�|���[�*`���Jwu�E�W*�j��*�m�����c�����ɔjb�e�N*VL�fFY� ^��LI���\Ѡ*��]��i&5cam��S�]ƦS�X�:��=̴�����G�wC�Aќq��f�LR{��.V����6t�bⓖ�xSa�Zme�����H�N*�-���RV^�ݲ���})$��[#��I���8����'���o�?�����_��/��������������L���Ϧ����	��6PY�Kx�� d�c8s��d����b�j%\�*�t�k���F@��+2T��|.��Ѩd�יhm#�P��8)�v
�b����ʻ�K\=�����=���eq�9�QIË2�gJ�z	5�����wv��q������F�M�w�9K�N��f�`|/�:D!܊'�������ƞ�=�xyߖ�̳��}���N�s�����Y�:Tv+��3��j�2	�Ћf'���
�Y1oia��p�Z��C�ʖ�]�x� ;�E�d�j,ݨt���}H�ܘ\"�6u�U�yҷbۑv�;�G2pWt�8�:�W�/V ccò�"�|E��6z��4�BH�r�f�v��O�-���fZ.���=*7ۍ@u\��\�o��Cc&�Mn�r���P �כX�e��j��Ͷ���'[ZZ�F���J8�̔/yͬu:	K���z��tls(aC8^���sT��˻Z�A��o\��rv[r�������G:�7kw�2 ����E��Qmiܰ�x������2�mj����8��|�e��2���PW|��]��|�V�ͩ���oPg��{u+9u"�  �ӳ�![�dwR��uއg�-B�=.���u�#Q��@hQwJ��)�n@FH�6w�¦ǁ�T9C��7�}�_gB\\2��L-����������CEw���0}t�YT�N� n��xZ.��u�㪂�E|����s'6h瓚���%p�<>;�%����˗����uG#�9����u[�
��n9㎙N���M�9~0�G�8/�Ut�s�-]g�y�$=��By��{�'"�4�9%Z*R�D�a����O����J%>0��#�yT��z���{�0���T�����m-�P�Z���[�;����rGwW)c��_����Jse��qc�I�b�Hn�w��+���Z���r �5�q<�)K�+���~W��z�{�-�I�wtG���]y��Ih�����8m3����[�����NN���#��xd丫r-��p�H�	vyT�wKa)��MD�rz�<�B�v�{#���>�q���xED��>:ݴ"���	��s�[�ɑr��R�-z/>��;��r�%c����}��ӭ�\��O9o��S�|��	����Jn�_1�'���%H��B*�?'����p�G]�2B�J�˞hb-_(���TE
�����Q?!�G*�H��H�Y@+�#�ک͌q�轖\��
��ǧ��x�Q�.�Zr��iN�!s;s8��q�A#��.�7%%u�R�&6N���v��j��ԟv���Hs��~�*�^�9��ܭ�!����Bc�������`����D��xMFFι���Ȣd��ʺ�|g�����`7�J4�\��i�>���U爑��Gh��A<K�9O��ͭ��Uy�qn�e�t����;�2�`��5q���p��ۮI��$�0�;y�ͣ6����{��5l�W�!�Rʕ�=��T_N����+gە=@����q�g�[Y�}y:N��Ͳ;g��PaNA�y��#�ob��]n9{�/b���GYؚ�;D�H;ϳ�q�o��a����]?s�]�ߪ��~O˳����3|߲{[>�fm������<�}���d����t�(������5#�y�t� h��ݍ���'�1ʭ^�ޣ���4�x�����Z�.���{���y���ٴ=���7��rL	QJA��6D@��mm�:bth�|͝W9u;	u�Q�c��h�5u;����w�6X( �+��W+�x��U��{��PiCi��.v$m�7;,�c��+�^�-�`��.��<�d�̣�-��ݶM�ў=�v�`�n�$�.19�}��G�W2�Uөj�6�
S��C�T����$�)!��GO�N�eb�oT�#�c��Oj�<��WL�����oI���]��#�hL�0LX�.�}ĐH#=���Mc�싆� �����}��o��f�r.}�z��̶�@��y׽=O��*���T+/_d}^��a��I�5��Qa���[�Ƣ�-�Է������}�)��U ������z�m�'+��5�~CM�F���j2 n������Ο�9U��<I����.^.O�3��k�Q��/ޥ�:�����W�yd8�ۢ4�vz��=��?O?z��2O�I_7� '���죠��*�޴u���9z_)����}s=���yW{�l��#>[F����VB��B�(�����evI3z,��� ���I�����=۵��| ���L,s���4�=!�*�*��ZA�����Qٜif�yp$��	s���ڲ�ٻW[Ja�2�@������D�*���5�.;�-��!6M��q�u�n�R�7u.�6×Թ�ߧ���f�&}ow����3�N�8_/���ky�s��r�Tk�Y���S4���Y�ޓ�X�H�ßOC���ċ>��Mm3=��E��|��./3��5�Qza�r���o(�5F�F�_Sܐrt��Ϡ�-��If�9�M�yΦK�̊�d����������K��f�+�&Ekug�f}7i3t���r��9�����i���*�@\l�n)��nw�����*C�'n�0jF|E�+G������N^���6*r�篎Ȝ&��N�����*��c�b§w��k^K����l4���t������(�"|H1�����cNE���ܜ��f�z��v1F��v+g�t�e��;�	�S��4o��e �8�"��{sB��`��C�����Ȼ$��8w���*�h�Gn�xa̯VN�ULz��z�PqC��`dfQ����1[�ɩ�x�~7y�w0�����Y�D�I�x����w&��T?N���0+��81|�jQ�Z�j��� "���)n��g�9�ʾ�2��`�yJ�-]����P�s���-��t1unS��P�k�)r�]�S����5ogtގ�hlN]�1Wk���Ḅ߾�R��S�\g{�:&׫�md�ڲea�Y$�~YU3wǥ��k#�5��I�=&���:��L�8�]���a�!9�C4s��'��$��lI�"6��i&����{��{Gbۇ�i"q�z3�d���8Tx?`�dp�m� ���$�q�M�{�ݒ�)�{$���-y�]�0m�#����e	^o%EQg�Ӽ1���ԛ��$��4ǲ������g����ﭘ��A�ʺ�R��Jl���ڇ���j�V�<9�|���Z�j�Ml���]gM=� ���[WI�Uמ|<�x���4/g^�e={����~X��S�����4�d�H�ۥ�T��O�ؾ�ck=}^F%nXk�.st�0shs�Ӷ	����Xp�����r�����>ձEޣ[묂���5�zEN?<S�ޢ���<Ϸ5�-�&mw�W�W	���%gm@�>��4x����w��µP�7� CX�-E�t�Y1X7���w��m��yD���..ɋ5�3oz����]l�}���#��21�t�y|1u�����2�6�2�^ ����pf�@���:���2�Ud���y���&a��?������	5�Ѱ;/�0F��r���#k�2���2�p�I���|��J���yQü�^����A��J\�L��sfw����G]{�%�G����	�t�9��q:�\�E�wםO��I�n��"�8=��"Op��2h�luA��vE����v]r�s��E�nut�M�
����c8��|A71�wf���<�ܽ㲎T/FON�U�b+F���Q���A��q3G�ў��p�g�0F>ݜӵW�n���j ��a�\4��H=��I<s:�8��s�����.玸��!�N��ާ����m���G�`��j�������X��1$�S�v[d�$df������ MJYCކ��x�y�.%�{;��u2��=�������>=�l�fa�R�r�^��ן��jCz�K�*[Mv���ARJ�(�*��A��9�W^�SF�Q�5�9�{��߉�ۚ���f]Cu�SJb��K[�=]ӕ��9# Д���}��Z��*l����t��,ҷӵܔ�)�d���˳�X��b��s���Lڒ�_74j�i}���9�GYؑ]GI�9��a��^a�K���/\�ى�+7���x�L1TQn�醷��7������ۡP..~k­����q�^�������"W��e��wi��TѣƯ��ך����CS�T��p�q�z�0�//d�	��ez[Ǿ�ʖ�Sƺ����T��k�m\�WN��U��R��zJ��!g|j&�X�ai�2��ʸ���}x�����G\�D�]#h7k�x/�\I�s&�ɢ*�	��U�ˮ��q���x��љe�w'Ă4�_`�Ǘٸg#��a�+�ؘ�r���C���6�uo�?6ר?�{Ɵ��F� �վ?<��C�������x	:f��Dh̗��31��B��#h��F��x���FAwϟ�����)��ޭ:8���Ѵ�Uv\�A�hFD{t�}���ܲ�EUֿz��6t�ʾ�gi��:;��bx0�q�u�*l뭎�c2K�]�����<yF2y?q8.�vг��˯o�{�@C"%f����Z��l3D[�$qeÆI(]di����jFǮ���	�)uԙK��~j��mԫ���xa*z�誻\_4ϓ������~�}ꕳ:���Ą��6)!ú�<�5��M\a�q�4�T�W>�ci�qΡ���x=�G�gE"�Ǽ����˭-�I����3�$� �[-t�F�R�[�"�^v�ۉ!�p5��)�������O��|�&l���ٜ81�.���aM�-��5�*�/e6�<�/�����}~��K`������_XP�评���U�L���Jx�<����絾�u��3ֲN�����U=��${e���u�X��}t�ל�J���۽�a��nƑn����0�R�� уT3e���k��0��nkP��lf�����z�:z�kƪ���N2�&3��h�3V���ӧbW���[��#w���o:����F~��^�������8蓝A�k�~�UZk�~�t��A���m��6���{����}��YN �	���3SV��z����n�v�r�cס�.S�x��r��V�l#��m�W�-��#��b�Q>Y�Kd�zb��J��8�{9ɫ*�Q+BY�f��GTس����{�.�w8N�f4�ڻ��Z���hn�����h�������Mm���*�*��o���Z �nX�P+z��7�{]~�1�d?q ��Y��-�Gz���J��1��D;��:�u�~�l��$ֽˊ����~,����+��_wc��U8���������κX�N>d��$�η��>��\���f����]É�3Ǳ�f��4�"����>+��e}f9�1>Q{�*�r�;����&���`��s�Nf��$�U����U!�o>��>���������Y[gd�M�&��&	���Ws9sBD�v��c�c��yC������v|$�%{�`꽜o���z|;��5z��P��c0<~g���kw�+2x{|j��*�R��2̨j,�������W=&��f�q9|	��:KQc���׫�(Jl�'�f�$�A��݋�������)��^��=�s��jt�(�|�V������d���_	O�[�ƣ�^��Z�s��̝r�J�:��Y&���o�NhT�P�y�+��
�;͏����6/9i�v����JD�2�s�ĝA���w�l������\2l�}��Zx~����zC��ײ�SM���:�x�5t�1�o���8Y��G�߾�&J�쓻��|��鋤�{g˩8}������#�N �B�C��jo��g����������kө�W�
���|�
3�3�m�����*�
I��-q>�~�eN�z�3�<4sI�BR�Y3;ؔ;=��<�����W�B���� ��7Ge�&���m�yvh�PkA4�.;��یӷ�gi�{!�� etώv��^��[��^�#���*s;���l�5y�A$@y�ì`�C��>�]rU^�ɫ�y�=�box&^�5s	���a!�$�w�{G�_,���f��K��[�ײ:��|��}���ԧ������OGf�ܭ�#�����thӢP���v��������ȟS�FG�Ci����zM=u�Qo����� `���EQ�����J��[,B����0�V=W.��n�g�������i��nyݟ��S����U��7��D�{&��Z�؃��rN�Y�'r}#�s�G8V� 3��5��	r�˭:�p]9�P�9�6����9fƥ��	�h��sgi{N��c$��|0m�A��tӸ���k|�3wWR�����Bg��1�ϳ!�[8�o�3E;m�=�Ѯb"λt6�;�^��f��Ϊ-���m�>�L��_�C畇�]V��۫��$�؇�Pׇ('OHy�?q�~��}�L�������jC0�B��W�Ԗ�C�Jӈҥ��Ey�u�������3����?zI���.��Z���MLZ�h��͑��}t^IE�~�a�������[��o�=�U�6_"��si�~���T�^���&�ɜ5��K��wi��=�11�@�gq/0WivW�˔Q{��]�=;ᵠ����t`ȫ&�q��M��`����۫���[~�2�^{^3j�R��W�v�U3^��ӽ��P̝��N���5u��tp�]�݃�����a��`�� ����8W�-ظp��ـQ�:�)!�>�P�ju�+ܤɜѺG�L]&9�k���/��ٸt(���Rh7ws{"�̭�]�����ˊ
��ݘ2h���֍*���[�
`�9n�#H�SGP�]�C��{s_;4x:}K���闝A:��J�trQ�D��`-1�6�A%*�%���П��j�g���g����Ь�i�--�q�rm)݉ڵ�u�L�������*m:Qs7JR�noa]3����MWN�\�د:;��⦥��*>фN�T̎�*�\�
 �v�fLKq��s-�sR�u|�vң��̺C۵'��X(ϻ�ȭ������&�BC��VP�[�m�7ci޸*cYɵ.��QڴV#�I��\k���DPF%W��[�bQ�@���l$�QV�<�&�g��痷o��F�
�|{$T :�m��ɝ���Y����7�()��Ṵ�g�_��,��;%^���TZ�~)	��R5bK��N!�6(+��bS��h�<=�n�����%K�1P���bsݷ�(���TwIU�q�^�7R����o�Y��=�>L���.�Ӱ������<��y* �t�����f�|§�y��6{����1Ю2�Lt�c�g6I�T{�	��AS�Z��Oi`��]�C��g�^���/D+�g3F�:����w�dr��Ņ�Y�C��lS���K�ݚRv���'ê]#�c�v���S�;� �����JWV+��o�y
�OV����Q��qoS˘3��MY�N�ە�g}���h����Ԯa�i2�jވg3w��:h�.�����*����*�/7Rs"��u���}��E�y˕8-.G��J
of�!���H�	#]x��eEC�����t�-���L�8\�sZ����x�J�6
ݧ�����/�p(�]YH`+5�Z�Ŏ�),�L��v�.I��੣g p�5�Y7�ϔ��S����Cfշ�%sj��{���7��n�^���z r�Ǡ�n�Z���zcsEoL�Ma�!��l�٨�6(�V���Wo�,�22K{q9|0ҕ�ײ���ʻ[j�B��W����ce���Wײ<}�`ށ�XT�u#)�t���/�������6��9���1E�\�F4:����I���Z���4L���	i�d��et�$�=N
�§N��C�ӃU���R�ݪ`|v���C4-E���m\��i�ڴ��jU�Q��Y2�=o��"[�l�,-F�g^��M�P���%��sʬ$z]��hwuf
��/z�����<;WR�XKHCW�˻��A{h��&����V��WI�:���v�_�t�0Z�ECVy]$��W.Twq:듒���sj�
�ԗ�/E$yv�TLs�řk7Rop����}����%0��n7���bN��\���+�y�����2Ds�7�T$c�ђ4mAڝ����(��Ģ�(�s��>3�ZN�n�x�f���"Js_:8R�nȓ41#=�sW�W�u�^9�
�|yr�.�*f�r�DU��D$�EI:E�:^�*��-��^�+�*����H�p�M
��NR��\�I]N���7�^R�t8��f����$D�d�jN��?(G�B:����<����H���:�Uʤ�s�.���ˎ󔒛��J���|v��B�w;�t��yҼ�VS7v%貔�"�S:tSXP���U$*�K7����3��Gv�9�d���9�й����=hID���9y]�\���͕�*��'>K�H�IC�ZN_^�z��S��WL��W�|��W�UA�	��,��0�ܗVV�JX��I�{����y>��|a7 �4]B)�9�Ft?:`�a^y9��)��>H��z!'g��Gr+u����TSOt�i<%�ˍ*T,V���sd���8O'v���YI�����?>�o��߯}�_�uJ�L�43����w�kyp@W=�K.��8iZ���@wvN�wBA��C���vZ��t�n��_S���P�3���WA��mF'+ &��ݬ`��H=x$ ! r4�[E?�b)�7W�%��s�1����1��d�VŬs�!Sڞ���잔��wj�haVa0T�#>�ͧ�ʃ�9���>��kl�S��,�
�=����&..��T�>S��&ڇrTͶ0������w��f�lD,±�;�:;৽��R{`l	I��h�輌��W�Z�+����!�6n�á�Qj]c^�s�T�s��Ҡh��]��Y�uj~���ip�+E��(�	���Z.d�G3-��d�]�s^q�^|��ĲOa#4�J�����fF�+�J��>9-Ǒ6�no���Eˉ�j�*�}���_�``���Vħ�O�bS��%��5��\�W��\:��)��qR�mm��|{b��ne辖l�L'�;.�O�J��JO��Rr���)b�Û��/��+C��o̀�2��s<����8?�����<�b�K�:���}���R�Y�/y��dڗ9}��'!�4bXBJC��0�`g�sL9�vbYs�VM7_�Us]�� ��������˒:2���|�Z�Ҳ>J�w�D�_���e�Bg �{m�1��J��V�'��z��ӹ�r%F�g��|^a�M�s���ˌ�v�ms��dΧ���+a��t��ٚ���mDyH����6�c�ڇ����?=�i/nD�K�^�O@'�|;�	�^C5�@!n�h��N̉��`K:uc�KF��f�֮c}��yl(߇�����'$)#2
�9��G�F[��2�Ei����F�y���S�����O�l��_p?�u���Yҳܫ������ej��������cu.��%r��W'���0V���QE�?t��w9V���l�=�����������1�2j{\��#�+����w&�	M�j)fM>��n��MS<�46"iv�89�%�u�z$� �OLLLw.�����S����;͓6��M��{g�kP�X�ħ�VŮ����#G���?[� ��d8u{���Gӵ����-jJ8Zj��3��
�d��Pb�YUnOh�(�Za)�P�aw+!�*#�3b��s�<�F'1S]�.�l�����'���'+ K"��>��|jʋ�5p	\9�޺����gs˸"�DJ��9�<�Q�
)��0����_֨{�yu�H����$��tsT��lDi6g�I�ـRH��B��s ��`�b�y��7��ޅu���Vc���u�u��)��r�;�+AD�\�M�_^q�ܮ���:�
h�/�J)��9w�yG+�Mf�8�8�rg�w�+�!Zz.e�`���nʯUTy{ܧ������?2��p5�7O��p���=��N�#BҙI�X��w[���\.���9|˘/WE�m���p�A�m�g����3�{A�}��JkZ͹#�1�N�>W�)p�.}�:�fl�;�0�h���>�!?t� ���,����1n�ֹ|h��.i�ﳕmj6��fۓ��sN"�6�vk�k������GjƼ��Q�Ϊ�}[^Ւv��јrFEkU�gFR�z����-�.Rz�������da9BD���X�8v�\uM�+v��y5��|�\"���5"ՀbN���*�
�y��T�/vZ���Ƹ`Ћ���h�5ع��X{d+iL3�~n��#�hv���%k���+�҂^���qA̢]��Ȯ標4��+͑h�zU��h�c�D��Գ-��E�5J���5�R�i�Z�2z�b�-Q*=5أ��d���V)��0S��,��qkr=˻v	�̢�WoCa-��r1M���j��f�1מ�h?m+�P��_�ʛ�Y��S��S�Qh��C���w��?�(��a��L����I�n{�\E^����n��6ч�;@�0?��u��SD�`5���,�	�y��QK�Mm.��,E�t��@���5��B�����M���Gn�w�#�1�(�Z�8�2v6��ixF�����LYf]�8C���C�Pi��O���\�O�cx�+�b ����_z_��GJw	�R�9o2��Lq�:݄��W��A=y+��&|�.6�5t�îyg�u}��f ��EV�
�*��D,ʴ�E��Z��jl�Ҥ-{�2���Q*�p�L)��Z�se��S'{+s�C� ��r�4,C�)�cEy��F�ʌ�:N�|k2*�hRyq�f����1G��2��s�N�eyծ��1*�,��!
��	��֣X�!)����}��f�-�럖R����,PR��7�Z���H����:�������m�<&{�����W���r�������J���.��OH�t���¼�|��ґ�ab�7 7�v����	T@NjU���]v�6���'iey�dRt��F�Y��U�ӷP0i̽p��۶�+�d�2�M��۞�N�^f�z͆`k�
6҇@⮗�1i����]N��1=٦/��]�2�W���6���Ƅ��tf)�m:v���2���ԕt;��E�cv�6�����5U�^5����3*W�v�^�%[��'�,���C趘U&f�|����T�{E
��x�a�=6�Q�kX&�:+�D��Ƣ�of_P7��^tv�m�2�����D[9����{� 6�5�_#O���.g����vOr#���z��<x�@?02ã�������j��E���J�`OBר�	6&"��Ʒ<�{�s]�Ӭ�<�r����D/y����ʚ8��v��z�6��A<�����k���w�+��,x�}IO�_��K.�fZb�;0�h�	���!�y{��i����W�e5>�-�ͲI/�����D��9� �G�F�h�5�Lp^!��[�;�B�Bb�9�U^����q1��/z�A��v����	�$ !>�i��nZݾ��qJ�!��;�Fl���J�&��Tw���zǶx�Wv�f�e0T��A�#:ًg]�����v�-wRf��>0`h�暜��+E�z��;3mܔ�e�A�s`d\�	��yڻ�H�Z�Yn��������q;���I`P]�>���t>�`��^W�e?D͸,�3 :0ݴ�o��� �M�f�Mhǥ?x*3�(�Ƕ�O���i>�Ō$vQ��`��E@�����s���&�z_н�Z��	�x��I���V�Rk�":�����S�H��z�Mnw
3t}WYN�m��PŘ#f��S�\�iTsEa��)(�ێ~�F�9Dٯw�S����WZn� ���������][kR������M��q��CcZ��^��$�>߯I[�=����eݨoZ�ݮWP��s���q��֨�VV�֭����&Gf���=;5|��(,iOd�P~�N�㘔��H�TJ�Q��i���k����P#�MD�<��]����#�Y�mIh�>9*Hԩ'b�t�X���T�`f��+�f�*�M�s�������!����&��ڞ��8ޢ������z�=�-?#�3n�(�F�����B�׳H�&d��c�����zQ��(d8=��n���𘘕{�u��M��߆H����П	�}
G��6�ϼ�#�
"~�z[�<���̉�ՙ����:�
�u��)�d�c]�a)9lF<�+5�r�',k����Y}�i�C�k�7��87j�D���剝��zr_V��:�ë�cYc߸����5�[l?�uv�� �W`�t
��:���y�#�]!����=�����M�i'�df�+�Bd����-��W<s�N�TSࠑbEu��\-���3�革
��T���v�G2W���w��)��@%,ɔ�x�i�e��g��f���R�$��~.S������/�����O%�6b�������f_I,����#��^RGK"��*�,�5���ǧlf�X�����M�9�������za�,t��5��ԟyL�~�L��U�!��]�l��2>��f�w��ګ�$4ݚ�M �J\��0���E%Q��IVo�����oWE����s��nHĲ�v��d0o�`7� �[��ܥ:�����3�z�Xk��OӐ%'c�DȺW�~����V��N��.3(�7?Sǚ��.C&��E�z�l� [:y�x����l��dB���}tf�l�Hҧb��wB	��a��q�߼���p:�w,��{�k�������D�|(8����.uq���ڱl �ɊN�F�+UI�5�8�7��c�!�-�!G����5�k;������	�>&���p��ێ:d-|{��	��#B�����2�&�����\���=�"��{;~���k�!!�܇b��1ԩ2<��K5˲�t�*��@6Ȣ�h�zwȸ�4d|gb�����S��/fF���6�.��/�lҘ����_�.��Ƙ�0>��D���+T��;T��kD��"�R���*�{jLk���j�,'�J疠r�'�JK^ش��Y *�GK4tv{�g--�iI:�-�
ZЈǞ���uf��� ĝqvJ�­h�vS~WZ�A{����{p����/l�h�O&bj�)7O,uN��  �4=��<�v�,:��t�љIo�,/f����(�ܭw��m�y��^��ډD8�μ�)�]�'�@sNbGo����	t��ۊ���V�5sNA׼����N���T�����5/d��s�����`�Ť@��]09��Ȥ^8�_�s�PK�Z��.;r&�!��T�Va��*d-�;��B���=0¾^�d�e���2=�P6���˱�<;j�NZk�[�\�iq9�6��+����~�	?�y��>!�qko&	�][�NͤL���Xy".&��\��^<�0�q�S0�����-���;Є�����1I�T��t4U����Z�V����0�3"�x���)����c��<S���π��a�l~J�h�=�Y��'�T��� ��׶��:���xn��A=�B���O%q���S�f�G�FT�*L��썰�r+���(,� ;����*����v���iR�A��ˡFʣ�V�6JO=%ν:��$���s�f*((�x �-�#���jn��J2a���Jl�d&O%��`6��n��C����8�]Ʊ;�\����x�ĦjU_��iN$��0��{�Y<�w(mש�if�mpTԃdN����MAJT)c�V,��H�i8u�{�� ��ތ��}S�eD�iA4�u�@��8n�vq�9��R%��
��L�[1��gA���^���Eג��>λ��^IE4r1��L�A	(iyp� ��G�e��WՏB͎�B��u�F��GkLg*F�5��r�ޭ�9.�O������_�}U���$��k�&��>���2��c�:�7E2)Ja�k�BB���F���&я^�����
��5i��6���ܑ6�:�%Q�P���0FaI�)�#.����2��ql��he"|���#����h��Q�9�uHLN܉:҇qOK����PX��%ߛ0�x̡⛙���v�5�\:�:��<`0r�� ������u`����h]��F^�Gs��t��tµ��3� ���t�A=�x���zG���]�g&$�lG���ь:"W�N�z��_'h��&�yQt3`��{�%�fK7P1lɐ���@xB8���.0����ʌ��7�a�5��|�� ��2�����*�s׊�,�����ă��8!Cj�FIq���;U�n7vZ2�]uC'47d3o�_�G�:�1^�lZ�X�c>�ys�| ��K�M~����+�iy>x_:�9��h1�n�0P��a �o�xӴ���i��㫕x��Y{xn��E��pS�����s�r��X����x죻�$���;�`x��m�T��N�gN���귊��k��� �{�&�O��L���mj�ӍyQ>�f/���?%�}^�r���)�ٕ��� �����Iȯ�e�ˆ�쭭�&�،.m�Zv��l����׻��=����O���D�8�(��um܂g�� g��d��a��)M��/6��5�,Aii!Bi99nUT�K�ٛn䥙g^�	t�w	�����_���^�z�)���6���Rb�_�yE�����V�JU�>ё*�↼�W��k�^Y�'�8���؞i=�3�(�^=z����V���]���ݗs����{+��w��7/7:���5H�B1W3�B	����I�y#4���Rk����9�<�������/j�C{�<qܺ&hJ��<��C����!=�y۞��^��E2����F��i��k��si�#1�e���=���ki���6׆��e^;.�H9*Ou*I��b����)�u��&�Lqsc8E�H�﫝r�o�tH/��@D&�ڞݱm%��i!7K׭Ph��]����;�&�eUq�	=j-#���0�=!�XF03�
9��q!��U��ĝ��o:=}Ӕ��j�7�+�b�7�'��cz�1���۴�;���(����R'�������#u�����r�|AT�m���5�BO�q6���~��PNH�Z����k ��- �EHс�W,��V�.5���y�y^VP]I�h��Oj���JQmZ���h�O	6�����5�"�¸����eM�ye�l��y�:lX��W�����9L�G[���A��N�\M�ȺH��	<�\��˺�z��r���3:W/�^��#Ya�;!�ܦ�KN���."���;�)�ʳ-���l��jQ u޹C7իUylY�Eo��_!��V&H�L�:49�芺9���P/�����^p\�5������i��ӭ���K6`������ʺ�Q���V���a�"1��j�^ǡ����9RtJ
�x4������駑��̡�4XT���{���vd�h�P�h�Q��9[K�5�%Jk��d��h>Q-��dۏ7�J�Æˬ1�T��o$�Ly3LYX�nY�0j�a���״�+�m�#�#X(`�v3k�j�#��Q7��Y�Z�Q��v�N�Փ�h�Y�ӈ]�"��ݼ�/�l�U����/{����Y��'��wSL�;wh�u�S����-
i��k���i>ߏ!�n�UƮ+�ElqG�.N|I��l�	����s�[�ٱY&9%v�M�*��u�m?�gVܤ��¢:��ܢ��:�;dѫv�
�cWm�X�ϱt	�HTӶ_=-I2�㒕b���kl9�īp�Y�0櫹5����:�ɼ,�l��Ӊ�0L���J��m�3��1aM��:SU�F���}�Z�`
�٣S�U������'(��F7���]�æT녕�*nS�{GhtÑ�������k��N��u^.@���|2��z��t���h�2��6�t�P����*�2;Gm8�pN��k�4�i�u�|/M���,H�&��ޛ�Ҍy���o�kE�й�!�1L�L�D�라'N�u���s��ib�M�7r% ��k����:������ң�kyC�����M�b��
��k�&�cWr�	�S����5��ռŪ�.^�,^����J*
�!i*s�<�	]d;,�#�xΨ7A$�#38�C��R����Jf	�@���S7�Y���>�'F��o�[U�m&���(�m��+�� �Z�82�LVC��b��(7��@'lZ�n��5�4�\��c/�3��e��b�ܢ�k��f.7�p|�̓�b-��^E�)�X���,��Q[�.�4 KŻS�P��x�Zƚ�:LyB,�2\�^��)�]oAkd�M �r�k8�t��U��7R��`({
W
}kQ)�ܾ�6轗D�E:����y��dL��y��W���AX�0�N��h�4��3jn��R6鋐��R[Q�Ŕ$�o_"�E���Y���Ů��D��qt��l�65]����9�Qzh8�KwQ�*�$'��IT=|��w[0Q�s��V�(��s�s^���_���.Mn��z��ݜ�t8Y7� ®$��ʙ�e�D�M|e`-Dn�@�^��v�@��KC�EL�jT�3�v��A����ۢ��I���ա�I������I&#���[����t�S�^�:��G+��*Ȉ���yϴ�q$�>㞵w�y2��$]�\��>��~%8&u�qȳ�rNRH�]N<��=�]\G	��X�8m�V��f�����mCE
i����C�PԊ�1I3W�N+y$~1�a�R5R�T�y���N}\�޻9_�B���uEbr�N=�"�����TehU��]ZJ�4IaA=J.�'NS��<�N�Fz��"VB����{��ANDgA]s�����|�*I밨�;��*ME燔�(�T��%UH�E��EY_w�Ih���a*Z�+�4i e�<�i=�C��Y$*dD���*�S�v�V���d��\�MB�ΊAI'*��E�R�$����Fd���*�Ek,�
,	T2�z�����eV&���z�*dW���T�����2�z��1E�]�ii���C ��֡߾�쫛��8������z��f]_m9QS4�d�T$q�[�Sy�6�}Y���V����N��6�{�4-������ī[�įޑC��h����j����ψ� ���U��c��"�xd���$l~��c���~����>�~; �Y]���j���-�=���vRpK#4�_�׊�,���6����v�m�<ƪ=J�A�2���,`0["ak��̕��� �M)E'kڭ��9�L+�=�X�'\�f�U�]ā�0Er��->�U�``��\>��S���w*���j�vTg	̪�Ku�lq/����dwEF�����ir��d	Jǐs��E�ٟ/:]v���=1g�H-�ơ�	]M�+���E`��="آ�Gڧ���['�r�w�����m�-	��L-{a�U��ثj�t �Z�A=�%��k9~��̨�sG��U�!7_�����������Zr��>FF�a�.�j:���{Γ��#B����M�H4�՞ۗ���Ӿ�#v��t�Ҳ�����M���2��t��ǹP^q˫|X� �V��-��Ӕ���GN0�zh=�����ׁ��ݿC?]�u�Lwç�mn�&-�&ڸ�*�^AD�~��v��}��=�ӭ�*@��
��ټ92Nn�A� ���7��KVs�z��.�]�sډ#�qO�ȅG���%Z�>߳�m(�wU���f"d��l`�+B��Ҩ4[�?f_����z����n�;�k�6��JۤRz �h�����N����~�!?TuP ��Z�;Ѣgp��exz�n�Ɇ�%�x��E��9�b-#$dN���ҵ@AYc������y��KN��TW>�U�)Xi0�'�A�]Gr���<}=�DM"rҴ�N���3#*�Gd�^lb�9��9�]j�Y�u��%QaV�y��WZ�A{���9Ff,���/6l�Eép��卆[�	���#�{L�I�c�^�W=�������*4�<Mki�����}A��T��h_����|�?d�=���,9�� �n��jZ�X��ط]��F�WO�oK5qS[W@����
�}��<�c���FZ܆Or�rͺ���I��d6�zL܇fV���]����R7����BJ���;
�G�YG��0��1���coH�F_X/lܖ��a��C����T�0�8��3�@���$I�`LAV"k/�`Qy�ԑ�e>���{k;�[��xja�W!
Dך�e�o�abA�$m��
�e~�13��f6���$m�xK�_�j�<{�N/�Y�{Q#�\��tє/��qn[�DT��?m�����&����p��>���̗;���8,�,�[ʔ��]���R�C�p�iaEwwW�#!�����u"��o2���`�2� >������8?"Q��v�����g��¬?'��E�TkQ"v����ˠ�,�p;�,�q+q/��:�b��������Jz��kƮ�G9�����:N�|h|*���ԙZ���rT����a<��?��c�:��,�?W\
�iu�5�[���w�	���i�����k�R����s��LR��]�ټz��	��؀�Z����#T��<=���-F�ռ��p�^�h+z{�Ru��K$�tI�wG�\���W�a.=@�k����9%Q�=�BS7(�`q�Tpc^:�%���0@#R��n�eC�n�`Ӗ���p������r��9���:��G��	���l�*�*�z���҂��l'��SY�$���������xR�c�ag��B��Cò#f��56��x��`�F^8T�Ae͑�pTº���\uԎ�=l^�T�n0����=_�ض@ɉ9��'��.LvXy6�Q�1�ȰW�u��	{��+RZ�̖n�����8yB8��b��;F��ء�!�ymE<�;�U�e��S5o:і� �m����R�Ջν��]��0v\Q��Ӷ�v;�[ 9F/���dTw��<��zsǩC�KF�húNQ�:���#�虅Ԭ8�SΓ4����$vV���d9����LƓ��ҕ�Qe3���n���i������{ws��7�j��,3m��Lm<u>�3�N�3<�T��Q��&~��6=����u�}����RsΥع;���~��=$=D�LW�l[�;���L�Z�b�㨍����ص�HzaS�5Յ�^��D�c>ݬ`��H=$ !�˲�]vND�7[W��ט��	nZ�pS��K�[ ��d��T^��қ[w�Be0AH�'Ek%�����o3>�{��1�|0v�y���ȭS�)3Aig�.1Nz�}<��Ժh����M����t���l���SlQG(=ٴ��V�t�w�-������ᴲ�}��BS5�M.x��xz]c�'"�$�)��A�Fi=�Q�aG�����o�����>�Ŏ"�zō��;
�d^6B#sW���1,��bY)2Z��:�̍TW(]���u-�^L��Ue^�Wb]#_��n1a��f�mǵHZ�:O�bS�]"�P�J�[`�-��y�(��w��}U�:	�-_y���M�?t�ڞ��`�B�ҥNb����ۣ��p{A������ ��l�iD��gw����2��z�V��t�C`�5�r8��ޒ���=���G�cD�]ώ�X��]O2���i�-��a��w�mt�����n�=;N�޳�lgU��Ԭ��:���h@��{�hv�"����e&��ŗ�o�tC�����|rFLh;#r,ϗ��%���,�}wo1t���ޜ��\/"��
/���������#`��@�#�N�2�2H�y��h�<�}أ)kr���;(������(�z>;�u)XQ5|w���G9'7|�u��zj����heP�}SY`2k��s��}��(��?��`����D�c ��b����W��T������:��Q�GWs����]���u)�S�X�8�����p��G�M��>-�C���s��r3��$!�������ma�,�g��=���N���0VBB�ݖ�;4��<JwY�ޅ�L�	Vxr��je<Jh�������s�G2W�A�����,�%�Q���9;m.�;&�{�)N�/^K1i>~H@���uE'�|e��
:f��']1m���K&��`�+Lb�4�h^^��L�@�Iڒ�d�#.�o�i�m��ȧ|� �Æ_�}F' �7/h�q��M����o�b��:A�0�&��G��eH��=hI\�j��*Pך�҆ -F�u���b��8,�\���*���R�]��;1Vb�*i���v[�x��0���
�X�Ԩ֕�:&x�D����k��S��f��� A�	iuN9�/�sS/�m̙��l˺����9��k�SdL+n�a
�QJo~�����z�l���j|#�����1��ðUm�ӱV�;���]�,�,�kY��:��8�n���*�7�x���f ��"S��j�.�;'Y5z2;s���@&)y��4'��2��jm9�WpR��W����,�ˣ��魟��N�����a�##.� m�2���WW{��c���-]E�l����*Q��q�jĪI��t�	n��~�ଣ���{n�:�̰�;����5�l�=�(e�5���	���"��(�����|��1���kÖéii`��+^ʫ���щn@��CH�I��&m�u��i�B����r��xCC�ޯz�+ ����M����^���uf��i0�9+�Z�\��~	IcA�a!<;�6�:��.y���ۺ���ɮAq�|BӮ㛓����Vj�Y�bN���%Qjf���=�]kZC���׾q%���
�4�U�B�O}J�^ �hXv>!a҇.>��#�{L�\J�[�k�w�WsZ���Z�d�n:�}e��P��ca�C�,���(pǦ
�z~Ƀ�v�L��?B,ؼ�fm����9/��oF=IE:\P�/vc�J�l��0�NB�(�F����h�rJˉ5'��_�f���^�y*y6����#��ٕ��9Ɣ���xx��(�҉Z�=�$|��;l��71aT�G�j�Ec���Y����]7�}�华�����cE��Gm�]�c�ֺĥ���UK\���g&;��h����p�K�o�ᄿ/�nL�\�>��_�z��K7Jܢ����f:��f|tE���l��k˼ `N7U������Ft�P�L9��P��ݻ��u����!��r2� �eC�mኛ�6�tb�廹�w]��E�l�%���!L�V��U�m��1���	Ҩ#���Fq��Y��v�N�����\�ӆ'�g��t���."E�B��yvUF��ɃFF{�v*�>������(�3V����ˍ�آ"��]8�8>6`�b��s��FL;�6��1��j],�˦��*�x*lC6G2�F����T=�x�Z�L��E�Ώ�1�C��f�U5/�q�z����.���fIjP�����Ғ�5)J�ߣb�HŖ�)�i@#�:���1:	m�V���rm=�`�K�k�;�Ru�1�d�g���QJ�
��W8k���"S�^�@��˪�ۡ�="�5�#9H�d1��"U�=�I�F�X�ʱGH������'�"�*Wp:��B�f�M�j�YGyErNdة�X����K�A�`40�$��P��P�<y2�s;jV�c�:"9+�0:�rε���!7��};ES�+�<}�7J�Tw)�ݏw�*9Q����
aq��Ӗ64�j/*�AZ!mk� > Ɨ\�Ke�������4��F�64�(p��c�Bl��B���*��]/B�Z~iFo�d���+�G��.�}w��!��|������~��'f��1Lh:v���n�L�2�~��K{6tr�t7a�t7T����*A=�ഏP#_��b����jL������{�W+y�+gkXP+�sߊ�^��+RYe�7�����S֮B�ҟn輳�|]�\;n=�m��*��x�}�gӯ\fy���1���1���e�k��Xu{yquw����^��A����=����f޸\�9��D��LW�lZ�>���,Pٚ�s´r7	�Â�>'�J����t��ā�X�C�&A!m�j3�X��h�w���G��#�W
_G���m�OC�8[�G�ߺ��잟&�=ک�&�a�e�!m���۾�ݔ��/^]+�dÇ�ٴ�<Rf(*����ßv�W�L�Ѫg�?�%����u�_�����Mͻ|1J�Z�`��rFl�zǫxU�)�0!E�]��h�64��fQ S�e�Q�{�"5S5%<LwH5f3�������7���+e���Af
G_U�=����X�4&��f����N,�� n�-���v�'��w9�#{n��X�JF�>h��3b��	}0j�5��۵��q҅Mӫ�W�_{�s�b.2��r�:>�Xr�دw!	�A2�&�h�'Rb�i�z�o�������b�)�s���(B��U�A��;�,p�U�A�N+�ĲOa#4���Rk����7��U;P�KU��'��Re.�?��j&�����0��<��S��^��%�͆�~rf�9Ȼ����Ĥx�&Ե�5��c̚0t��H�Dt�l1�*RvRNC�U���"7zao
�T�h6ȣXh��^�#ϲE���G��M����λV��:�e�����:Kgu�=���2��m��b���R	z�H�\��l��s�xj�n����˳]֝����z���vQy�cB߻���ҳ�<�"Ƽ(�8kTƤr`��yƚ�z��E�8ۡ��Ȟu�5"�׌�ƻ��FM�ߕϠ�K6W�Ż�m�YU$@�{OF��m���0��4,��ռ�L�-YCtеa̦A�k,{����/<�c3b{��YE��}Y�Z��о����+�qP�&->ɍm/}P���t�~�z�p��IA�����5�X��T0�>�¦t�h>AU��	j�X7��橦�*�O�xiӹs:I��D⮪����Wh�	ͩ�dN����Υ�]���@�_�h�U�Q�[;+/I��]�|�so>;g��o+�P�i��;u*�������:3�������ȭj�[�>��4#�L���F�/���^��{�wPn|蜗�/e�����ϵ֯B��Z��������^S�)?N@���:.9��5):�!���F���6�W�Wתec^�$g�3-S4P�]��M���":'���oΫU2n��t�@���|�!�S+�Ξ�]��S�S��zN�جja �ˠɒ�!��3���6ʲ���`*B�m��d��Fh�1��ѳ�.��}�T�<�Du���$����Z��	�� K"��>H�.�ʺ�m(5��l�׶�9b��T�k$S��@yq��˟#;q�9'o�J��������6�\:̱wz�]�qP�4i\��t+UdmE��tצ��x�?s�S�܍f�;p����E��������]�ki�v��sǤQR�'b:q��E�*�N7���i�:A��������0��'�_ˋ��C|d�O���y�1����%>�Mb�vl���-�a�2�4�r�t�c��ʐF�-�,��CO�*Rz�6Ⱥ��9���"u�CzV� X�#�&�=$����2������4R�BuA��^���P����nmgʎ2�8W>�i�W��p]�<�pC�R�
��*�nQq�s�Z\��d]��i �|1���^1.VV'#'��n�����y��Hkgn�V#��+��X�f�3V.H��N��L�Zb��*�{я���ke�Ysf<�C�z��9ع���"�C�{7&��9��ȴ`(����˗�|N���skWSb�[���kj5�S"�{β4�@��o5�#/�)�x�� i�t{
�Py����$Oz��q���p�s���.���m�L�z�L�#:v�6�eiI-�A�ֱ��p�5T�w�K���I*e8�X�����L�2V�F�=��n5A��u#h��T�X��XkT��������5�yp���%�MvvZ�T���Ȇv���:�a���M�+zc��Q-ڬ���%5ټ;.�Z�lyY>�R�E�sq]\@T�.���m�uewm�����n/����9[��	%"��6��b����z'8���Q<�T�AR�ht)�+fS���t�o	2�y�a�iuv�2�%��F'Vq���Ӕ�M�	�ܩ��h����I��%��Y�`,�(3;�en_;&�ΩT�k5�سj)Ɏ����鋷����i��\�|-clT�/q����|*;nqw�]�L���l�����]F�,����4��<�Qu���a+Ln!��Ю����]��˫�n�����U�Pz��ad׺�|��{]��%�#�҆u�e�d;w��,Σuq��=�\�c\�!g-���K�3s���6
��*8��h��T��x8^*��C�ch��]h+ZTnq�9Yj�κ&�gv�E���΀i*2_k���	n\�,t�V.j����p�oz�\#D�!aWber�"���cQ୷P�"��7���w8�qE�G���a �G*V�L���|�����Q�X;;+A�&e�휍��1�
�iD{w],�*�t�� �Yy.� ��"gl��a��=���@.��!�s��9Q��V|�bia�:O]�.��Rɠ�;�����̢jj���B{�d��z{�0`�VL��ኢP]Ԙ]z�w[;tWq؁L�l��J���d������k�t�jA�t�j��/1g0P�F��=�M���[%f��.��_l]���ou�	��ޭM'��l�ﯶQynݠ>}��h9���n�>_9@.���A9�3�[�����XG���b���7���Z�Tc.ݦ�*0K�b�U֭�� �1�`n��n�f�������r_q��R��������t�Z1����ج��%C)��We��Z2��ٹrp�#,va`��鵃���
�����D�P�e��gy����U쮜� ��¶���^�����އ��	جzO44���AI��t�Ef���s����@�D)�P�t��-,$�&$dR�T�U�Ҍ���&�r�5��Iʂ"�>A���L�8�.RE!(�$�J(�PYϺ��b�p�S:UvQHr��
#��%J�T��[S�	+�Kwb䏏 (v��Dt�C��6Y�h���G�L���D��E�,��<�np��#����8\�ԬP4�T&JlN��'��0$���H�LJ��%3V�[�D��ªi�.R��W$�Q'�AI$ө�XU�*�
�J(�����w#�G.�(58bVϻ�����9 EUu�M̌6Tt�T(�qd�*�G���SKW���(�P����(\uB������$��H�����B���P�a˴�24b"��(�j�=���]�g*�e\#�>̋�9�J�Tjp����H�jFG�i��d�H�,�V�Q�{�t|���̊P�"(��º�S5Þ?,��i��ѣr�Vޑ
]�����B��-J/�� ����e�o&�\W71�iw$>ѝ�� q[�nk߽� ��Kn�=�n��߽Aŗ���=����5�(��L*�J疣�)=_��Ƽ��0;7vu�*C^T�<d����ݑh��)HL;ˇL����7�=ά�K����,(Z��R�O	��\T+�U����t�#�?X^29R	��q���Bæ|}#f���B��D�q�]nC1�"d���]�w,��E�lq{k
��<Ũ;�0?�G��L����&	��;ße"`��S�ʇ����0,��PI�'rR�]^*��R���/a�ό�w�\=�V��<2���uX�dNv7vW)�+�Y�uc;����s��&Y��{��4�r���Q^Q��i���9�ĭ�)Ǣ��zA�$=�-F�"�Ȩ�޽�$1v��=���D(4�2� �d�mKd)�v�x��ܡjK�j��Ѱ&Ae�Fd��*����n�A�Y��Pμ?���y�b|�xu+^�~��	���zrS�X~!�Aw!�漻Ti�Td����:ҟi�2'Fû��V�EeR��2�.�2u��ޛa"�*��3�A�!���F����܄�}-��52ă\��1]J�]فVcM�����ws�ɥ��SO���N��>ZL�2�V��f���ݎu�5�W�4���~��4����O-�W�U�r�6�,�%��u�⎚E%�.,w��-�+�m.Rl��\g�)i5?�Rz{%��{P����5_���uW
���<���ߟ0N�2"ѡI�Q�`��{��S�; ^�B<�uq����Fva�uu}[T�hY�� ,S�A�	Ll1�N�),O��)c�W�->SJҘ�{��)-�k�]q�N����4��^�a�H�I�1,��n�dR�ß�����O{:J�W��w<�u��s&�7�.~�!���"Ux�
N�;"���J.�����٘ք��6�4�G�)��2AId�Z�c��=�B��P�x⮗�(�.�l�1�9	F���5�*�^>=9����!�[!�{��6�����EՃSlP2�!�&r������iܮ�
;�a�Z��S]R7T��z�yR	��ഏP#_� �_����z���Uut.����PՈ*���aJ�a@���~*	{���Ij2Y��b�9���@s���9՜^�U����}t!�ܴmǯn�7Rca<u>�}��j��c@ņv/y׺/�(no�f�߁<�z�\9Ś�e�sCvC6��_�1�I^$@9D�xs�����_�F��冰u���p�x�PL�X�F}�D�w�ޅ6���Kh���k/:;EA$���/�c*��� ��-O�7�&�$�WV&2�@�+��N=�x/�c�AE�6�.D˩��,f6'v�n`6�v�f�c������< ��8=A�$�E8�����>1.�89a�����J��K�:HA���X�C�&
�aL�L9��@Ф�=��p����N�_E���a��"Y��-- !�Zjb�'�uE����t�E)��.��,6�0�31�בҙ���
�WA
FL8y��O\�o#��\nb��za��p���x��;�+�z�{e��)���m�2"��g�됤^Er�ji>�!*�;l�\��l�j����뫕>���>�^�w!)��A�Fi=�3�+Ǣ��
SI�>{��8dhST������%�2�!ò�� ��ٲ�F*�?B	��?�#4�¥I�yӌ��,\�a�����\�����2d�\%RO����6SL&
�cH"{$���)�|s�]�l:���&���.yg��4h=��*�5�_Pc̚0t��O��Dtd�q\�`ߛ+��mU��^�Ѽs?E�:�S�5�&,�c��<�-� �z��cjx4�!�3]H1���]��cO:�wL4�����Z~X�A/^�ZG#�0���F02(�%3�쿲K�v��=�@��1|��.r��;���c���ٵ���S��`XV1�햦_��(k�W��f�N�U�_k�%-,r�up|y��/�%n�*Lg���څ6��'+v��)���ޖ�n�H��:�E���W�UUUzC/kq���[��sݏj�i���k���c��z�=*s�\m*;�r�Յ��b�%��5jDM��f�ȴ%�����uP�u`Ԋc@ɬk��I�X�d��ҟ@52͏��-��4�;�r�ٽ�H��d����(h��)�kVW�i�j�Ja��5�=���o5����s���P������OI�����Տ�c%g�YG)A�ǭ���}��v����ͧ}ܛ��Gg9SC4H�s��R��
�BƦS�_�9�ȘZ�GT�d�x�cr�^����i���E��[���J�Nܔ�&�r��'�`u��~�Y�pRҦso��t1̭�.7��g~Zg�ְzew/�O&m�;$�j ��A�܌�M����y��["����5O&5؉���R(�^��1sm��U\�v�Se�H8�jd��A�g�fͲ��p��˸l_#Xo�+	R��l\Xy�C�TGX����lU�{�O�xa����oA��pכ	S�y�Ⱥ}�J��=r魤	��sA?.9�s�g���]��!k�z��;*�?�.��[ɗWRRj��em�v�����L�{(;�<7����{��QWLX*�3+,ý�r�85�AڍMٓ!�,��Q��/+�%����rv��-��74q��Cz�Ƿ�򷐰#ԭ�ԥ՞���*��{5�W?0�h�����߽����dǊ��d���=��?T�S.���z�\.1�$Ao1��MO�r3��Py���>j���E��׈������^�Hеr�'q�dG�n��س@��G��w5I&n�4=%myV�z-ؽ�.�|��7t�L���[t�OE@�f˳e<0�� wj�����+��gz�5�ؐ�����
�p/G`K*CH�I�ɛd]ax�"�6�ٮy�ǥ��z�tf�⵱��D=�Ԏ���r��7"}^�L(�.ycu� ��&ݞ�����
.��S�|��)�K�u�Q�
�AN�� &��'��њ�GA�:������n;�x�*y
�����I��91�;ʨ,2�A?�
zW����	\}cf6����k�i���U6���D�Տ�������P��G�P/a�ό�����4�|Nr.)\�Eb��Wݲ��YE�5-X�p'3\�=�Y��RŨ�-=��d�B��N�8�ES4%D�	��|3��Bbf���f�������r�
ėj�1נ8��I��u�P��^������W��6m���u��m�ej�л�)�j�w�	5n宜�,;e��F�K���K����u���c��<�JwC^��Y���M[�#I3c�K�GO���x^ܬ} ����"�xvU�.u)�Cn��`�$��=��Ú+W��o�.f��.k���uLi7F�N~��*�~O��+�^�β8;��G�"�x�;�������#�̫3n��{2�:C�nS������x:�1w=��ˬThn>Ř��gkχ&*c{l��G�k8ڿ�ߧ�K!i��5ڠ�����B�U�Z.���v�����7�
h%#7���;<�c��A��B�Ru��ޛa"��^�rS��ً�`\1�t��f����kf�����&]c^��b��(Jl�d&UhФ��G(]��ס�V������Bu�m�y�O�oV����a�4�:+�+�4�S�A�	Ll1�N���1�R����*���O��P�,�8��FUe_z�k�y�|��$0/C��=��=�):�ĲN��)��0�KQ�7��	�����}Ug�9-����ɹ�,=�!��"U���ݑI�Ԣ�)�KI�j��:�K�j��j����H6�%��M�z��M�B��P�\ꆓ,�1��Օ}��x�.���/���}9���!&� ���0��g&'ˈW�������o_�e��o��n�~��� �jκ��vTT�>F��t�]\�l���F�����c*p���|���z.��Q��s����A�����8��R��Q�ʻ��.T�������¥�+�X�x�{�$�=�NR�+u�]&M�1WS<�m]��ػ�{���=�xs��=f"����a��om�J�Adw:�WC��d��(-�ఏ}���v��Ά�2e^l'���4۶�-l�)��OJ�T�.�Aew�@1lɐ���%����뱗�7�����'���G�ZV;����3l�AT�ߓ�S�1����g��}��-�{��:��9�]�Q��	��<�����}/�P����>�_�1a$<x ���A��r-��w�9��Z��!���vS�w�r�Caqy4���󤉠�}�X�C�\�v�i�y�=7��r��t��D�i�|_E!��ɹkf��x�#���t{�l�׳,�|lt!��Q���]z[��md3t�4P�)����B��E��z�ob��-,��Ϗ�fw��X(��3�3��B�{US�O^Y3mZ��m�2�*��&�Q�C6m>4���t�w����LWdXy����d��yS���sլ�y�xw!)�ɔ5Fi:��G�ը�Ϩ�C�tyeׯ�n}����i?`d��`r�d$�f�"�b�jЂqDĲO~H�2aJl�/.�mc�e;���s�#��D,H,�f=���yRà&�r�xY=3.�kX��¿��´����A������t��*=��^߫fd����[IiV�gs�(]��k,R�Y��pɍk4�![j�\��jK��WYz̻��r>����y����E�����6����Ϫ�J.8��&�|GH�0<#n=�|��'�3O���
��g2�4�
�m�`I��t�^�JZ��cȚ3��rrcA��B#�Oй �	��b�G,���&/z�eo>y�Rr���)W�Qa�Dŗ���찋`!#��"mʶ9^}���壓uOg:��gvza��&�zb���R	z�ZG#�3Ǥ?Hh�����S��q�J��:![({��LKj{�ɦ��U�ga�H�R���߹ZVvG��u�%�"�{�������P��zB�e��<���������,L��ғ��FM�ʏ[٦nM49&��9�#'�~+!�d?���Ż�$��}!�<�@h��)�kVH�����&5��m[�d�n٬�2'Z�ǥ��쨭j �`HFĻ���ƈLZ}���l��g��KT:��ٛ��;b���є�8�ٳLB�EM6����T��E�����t/�SA�SX�-������B�p��AnM)E':;��1������+ʆ���# BO��"r�#
Y7`���+|��)�X�N�hy'ץ�8 :;(91�ټ���'i��[�2�]'���9��`hdcfV;~�f�u�*�Z�fV���+��4-�8��;�jV�9�h�Mt��t&X)s����L�J��Idk\"F���(��=�Y�k�������ݛXd�o������7[��@̳L�C�Iv�6�7#�-��={�m��Rᑿ���cv��wOU���EM���I�v�ς�������^�	]L�A�3���M��u����������p-��򔘡�\X~�f)#�L��sG��O�e�/@�n�b���Ao?lB��_�
��Tn��]H@p�*(8��yی<U�������jȘ5U'�Y�V6�|�y�Quc�IL�ں���鮥eX��~`s�S�0���Q��]G?d��۰�6��y��{bS���DJ��]�N0��Ы�� ����9�;xU�l�|M�ُ��Pp�s6PY.�4����J�,c1V�"��D�6 ͗�;�0�"I�~Mu�)�jem�d�"E��^�Ѯ��A��,����ݕ)=Ⱥ@�i�H���qyJ*�+#;���B���+� ��w<Ð��^�NL܉:�aTrW<��)=*9��i4v��ٞ.�����*̲;�H���R
�A��8����zn��1'\[	�����*����ݼ7[��)���s���G�ה2�OIΤNs-ڧ�\V��v�����R�>�Rxdd�NWu���:�'`���Uܤx���2c�D��WQ4:u?�Dރ�EuK�@!��G*��Yժ ƾH�rG��E���/�}�U}��]�\Nl�����<�UN���a����;����,:P���04�ߝ���]a^Y���+����w}��w=2
��pK�r�����gC`�^Z0TSA�yv�p'��,ݴ�L9��T
n��]䥚��
�b���-=x��s&D���p�K�w��Y]��!�u�� ���;<%ا��f��LIv�,�^�8��HD[qm�ݪ`h����:+����Ç1�1�^�β9�L�dY� ��Z�
��V�Ǆ�o��܄W���8�6=����G^B]�w-.�Q����>���e�nu��ͬ�Suf;�)H�^��H�z~0)�3�鮝rSX~ :�	��e���y���Η17�����6����n�E�����~�2�]
VO�9�DG�Z�(+��F�^5֍o��f�ܡ������f�nQ�͡�	M�2*�
OaQɡo�Ӛ�1��1��(�=�Y��%T Rs�u=�"9����y��vW�i�b�j~BSbS�	I`���B�b�׼�(`�C�	r�EG+��G$Cf=�x4����/@�9��?r�8�Z��Q�fwmn�Jw��\p�gs�7Ι�b�Jz��A�&ۅ�xT�֭�w3&/pU��p2�����pF���`H���v�JJ���r�vۥ:�r�ae� ����π�ƨv�4\B�]��t�����si0+�}펵����r���I�V�����M���/�c��͡|Vۦ��~n�ܵ�p�vY�K`���v���t*l�XD���ܮ<̔�b��\A���ϴ�btyBR꾽�ݭ�(^��:���N=���V�ޔ2�[r�/3'0�$d�|梐�f'�h����l��P6F���;��]�I={Y٘�pqe�N�}�Y�ܓi��I�a�����.n�Ï,��˷�6���|s��1�]�]=�Y{C;<�ʢ���i]sT*�0�g���ϵ�`^�ɿ�ա3��b��m���w�'u'ܬ�{.���7�S@a��5�n�[�R�l,�6L͘;=x�XBS��Uκ�W��f�A��I5*�����S&�έ�š����1lb����Eʖ�ȡd���u�FCF��x�꩒�6�Ƕ`���J�Y���΅D�^�ԅ��c88C��[�Ct;f��`>S\5b]�n֜�P�����e�0.)�떍����>��tn�>߅��y5���g:Ut-ͷk�W�Nsr�7���`)2ws��Wt1n�����K�Պ�9ԕt���-^�Ӎ��]����v�tg8��q���ͭ\���H+�`���)e)���}�U����;]�o�Ͷn�ї��gl�J|�J<�=f< ǐ���[q�����\�Q���[x�oP���ʻ���ڀ���>�'l6�n�ܫ56�u*\��#v�b�c�eL�Y�����W�E��M��qP����V9��P��%�"�ꗼ�%���R�˸�Vs��u��"��6NT!�%�p�pZ?39���s̐�.�8���c^��t�4	5�J�%�"VP�h���Ko�Z7����ٛPnWmԎ!�H�)vf��M�7$���YE�Z�PGf;5�J[nG�j#H5�}�ڵ�J�Oy�I�C>2�Y�j�y&����Ǹ�����u����ʹ�Ҿ*c�gӟ>�gd�&Um���Skm`��Brg���	�ϏR�7�қ���S��^�������B�Kn���e���F��;�}��/M-�S}q3%.�;tE4���e�?�e�$��̭�5+�8��9w���j��]Sb��@��Ed���ѕht�R����V�ے�8)r)�ǥo��6gt-���N���@u�h\Cz�j��֦�yt"���7��F<ȅ�9Y�"����9�n�[����]��n�bFDS�/O=͖�_ox�%��TsyQZ��*#�YN�����:���/���J4��ǅc)��ni]��ѻ�C�[�v�~�Dujo��,Xx�Pi�S�`uU�Ml0����V�<o��e�������{��i��M&�*7@2@�ʭJ�fW0Ī �I�̪�b���s��(�ڛ�9gf!j'HB�&ZV��Xh2�
�R̒J3HR�¡*J�*Q0ɥXmP����Uq9q!9utp��_n��\��(�dQ|�nT��s�鮏��:��}�ۇJ�sʒ	��8sͲ���C4�9r���p�+):Bwu�S�C��u�zrs�
T#�B�̜�'&��E2�2�N�����x�+�K��*wZ�M\���!M3�r�;|HTaL�B×2��Ֆo������	s�^�y,���|(\���0�V\�Ӊ_t�r�baGg��T��܍i\/��#JAn�d�:1�wnNF���Щ�Fi�t�:��=CB�	�	�����ۥ�=�>�_�ԺE�Nh�8�z�_��L�8�w�}��S�I�R��!7!p��~{�?�őHd.��r�s���~>��y�ﯽzϦ�Ȝb�ĵ)�G8��X��S�PuGX�̕���>162Xǘ�Us���/d|��y1P���S~��=���t�a�D�k���y;�!�Z`��;zGt�N��K$�k��z+�]꓾�l_x�t�8�P�U�XX�������?l����`GP9J{"��%�7GRjz��]�/�c����lS�N�F9f`�������li�u{�BcGr�p:�eJ�6��]SJ�sr��hoV��)�:妇s����KL��{�,�C�X!q��n�X_
9�xͻq[6�����N0֥�h]�Ta������w:�ϣʐLn0���I��J}3�^�nֻ�u�>N��*�m]2Z�(S���{A/r��-AfK7W��`�`mc�������������A�9��<����1���7:m��
���x�|�gӯC�F�S{exz=Yҷ��h8�k=Z̬�k��(�s��9���V�b�,,��!�dvJ/���=$>��Y�&�&.EK%�ynR�J>�
�}�=�(A���\dJ�/�Q��a4�nf�ԓ{.4����ϴ�
�W��=y!	ޔc�,����kd[����`��-��ãܾ���u�+���;�G,�
�D
�o%I(������r k��	�<ގQ����t�[^�������K�ǤO= �:2����=��&��z��G��d��ՃuNɍ���Ԩ29����fҭƷ"U�0��{8s��lM\�_u��F��{���0��`���&���1����۸e�>e0TuH�=��AV9�cTRf1ALPz`�e�~�9p��l�T[_ub�������*�}%�")�JTͷ�PeB������5�mM'�L�����{n�6��%��~!��rr}H_�ְJ�b�=�Jl�(2j�f��TgP����)�u����m���۫�)��Oԭ&0kXpG\�;���P�U�^~��&%�t�[���p�40v�n�cL�{JΙ+��RL@���ya�>!_�f����8U压�΀�e�e,�WKKݺ}��]�A��4k�d+t�j�"d��Fv��?~��ߢr��}q�{��Q����r99	�)?9�NP��b�Ú�1e�Ϲ�l  ��%��n��uk�6v^?u�Vؽ�$6ז�5':�ۦ�u�-?,�P%�yH�Fi�O�H~��Y�KFVsVsUs>�Tsp܅�% ����(���}5���e�}^g�����)~	GtM��ݓm��q�i�J��5h_�ݡ�;���\�����\����׌�ƾ�I��#&�Xj&��d�� �`�Հ%~s�~�����y�d�ܻ���L흃��g+f�I;c�:�Z�N�3�r^oN@Z�`�#�멎v�B0��E˞��Ɋ���yJL4zv ��v���c0����]�����k��R^'���__]!�{cc���~��{��g���fY��>��2
��ix-�.�ֵd��hZ��t���1�P�no�u���Z�����Q������h�k ��-)���.�7��-E�"�-��]Ƭz�%�rrs\�Fi�����TQj�KE.2<�$�S�lr�>��d��|N�Q�k
j���3���&��|��i���vJ�r~w�/\�o`C��ˋ�z�����EP �kH���u��NO���3,�4W�t��TS ܺ��ִ�p�fB�!k(غ�c6{��RS�b�c��E��nn9�i�:� ɩ+��Cz��D���8�1�|>»��Qɶ(�Q��I�C�\X}��RGd�Hѝ�Ö��3��`�^�NN�f��21�d	c\Mk=x��f@�tפS��sA?.9�\�q���e�T�gs�*EC�f���J^|���LRux�
T-]���8�:�5�)�L@~??��	�<*��bF*=�?e^WMv�5m�ㇾZ��*y�%~Hе	�����Шt�xu�����f=�̛R��j�[&�䣶��Ǚf�	�Q��c��P��z��v;�Png����P��)�E����+k��h�>����������������3,U�R��|t��a���0rt��x�7cy�>=s[�>�1s��D���wO�7s��n��xxi����tP��gk���81�d{�H�I�y��Xn�I�h���i.���q��,LgV��e��z��B�p�.�T����m�)=#ȺE�sj��F`�2�FJ5���%�+֦�̆��D7��4���[�痫�MȟP�O3��;TmU�M��=^�*Q�jx^G��K"&�/-�PVr>!qԇ7��u`�гz�����GR�'N�"\r����,���XH/vZ�= �؁x,;�æ����fߑ��J������]�E6%������X/ҹ�(%픺.8#�y���g��f�j']�̧Q3����V�h��0��z=��Xk�P)�'pJY���b����A^�ό8�oD��~s�r�ss�����,"E8���2`���7`����	�.��1���f���4�]e�pP.tks���nP�5��j<�&4y������d^EF���$?��x'#v���T#E�X��;P���1��ʴ˴�`tv~���`�,y����	���X��0N���}�
��j��^c�u��v�O�fYo�4�hh�Q��3��$�q���Մ�φp�腾0}�RH�G6��VVAo2��좐��ԉ��A�Zir�^�Q걘v�ۄ�	1�a�f3�5c��x]�/dQ�7)�e��뾆�\o�l�������[�\��Ƭw9�����}�׎�uDVq0��ƃ�|3az\�3��S�\ga�]:����܄ws^]�Rv$Q~��J��T/n����G���xaTˡJ�Ty����	��c[΂�̋��]��S�o)v�=��CNԶu��;R�������2+FD��{I^�p&lk~�/�9���{?K͵��P��iN'��4�HW�+�4��O5 ���6�%:�%%�jR�^��z]�Z"8��s=Y9S�ً�-��J��O C�bp/��#o��7fIs��K�{&-'�A�/�ڼ�K�xi�杻��u	UP����M�|Gj�^�u�J�����C�=*uKV���Gy1��q��׶Q�~�� $&Rxr&����ف��[�y�2�,L�ۡpu�2��)��](➗�Y�O�~J<} gG��#���,�}�\p�uW����i�r2��U�Vֲ�����q�j ��c��Adw:�
�w=�3��ۇ��-��ui�E�woh/&�Oa��Dp"��ŕ�s�lύ��DzV��^��Z�Գ%��R�jX�gU�Y��+��?��;( Gc��ǅ=k�Ou�Gwmn�B�졯<Air-�2A��	��ެ;i���c'o��ș2�d#�6�;��K��r��;�u��K��tHw6S��J��w0���]7�T�݅fڬv[zpWq��ɮ�V6�K��G�xx{:�/p��/���`0o�5��?yG�\a�G-N^����OS���dϧ]��1��E���޾�YU�,��S�g�ɾ�}���(!�����uC';�(;���.L�[�Y�q?��!��H��R�eԝer���������k���c�!n:0��Fs��oMos<�(��;D�e^N��P̬`a�	�����F����H�孟��O��-��f�e��ż�B�ٻ9�\���.]j����ws��"�GOuH�#�h*�<�j�L�()FV��2iŽ3���jB�,��*rr�Lǡ>�L�P��m��Pe^�6�5�PW�yun�r�e��P��W����5=�!-)����윟W���	_�b�܄&��2�&�Fi=��y�7G��`�f"�Xus�S�4��6������?���`�1W3s��5���b�o칽Wעc�j��D����ƒ�TlTW(K��G�I�v>#�l��嘆�3*"��N_?M\R�-x��cžj��r�� ��wO4�i6����<΀�Ȏ�'Hv�>!�~np�FAC\�R��$�ő;.��kUwPӵx0�9L�lV5:\��hެ7�s��{MH�ͺoǸ�2�:��H�/p�2�pLB;�t��k��\ʖQ�[�A��!��e��ѷ:q��O�U��US���z迸6}�.�d,�'��$�^S���R�/��i���b��ϕ��~(�p˯2��9w|�;����f06�;g��:�A�M��8ŧ匤�7��������1=AՌ5ȍ���-�]��5�Ha�
:5i�ՑNh���T=��Q#�������޽�覉Tn�E�[5�ާ|��R�#�J#�5�Au"yo�fEs�0%��6�}�)9n�y�V�ˋ@�&��rz2�|�}u� 1��	W�b�д���P���S֬����o�
�^N�G�v�;��)��5���M��:d}��6CGug�J~�������� ��-=^��*]?�^�;)��ya���RpK#4�$ ,⢋H増TS+ҏY�p.,g�K�a����k��Δ�wPns�e4�Jm;RR̚yAwC�|�o1Ꭷ]b�s�MO�3���2�k� LL�:Ω��s��f���t��^*m�j��"��;)�S�������Ry^2;�H|abb���Us���lV4������x��1��lV]w@5a&�Օ��%*wZ�޺�@e��ݭ��i%�O�᚜��
�Bvs�7z�#�֩cy���3߻�5B�z=�����8
b��4 vh�!CX���| �&�Y�u�(�˛�,.��n��������&V�b{��q��W��}P�N��[>��n�z͛n�2��愦������}���&rGu�4U��}�rQL�=A��;(�|k� � I��N>{J�ܺk�)�Wb�'��5�(�d5��b�v�br��ack "��2�V=�b���
V��
juE�.��� ?�	p7��X^f���ʞ75�>�1��mp��Ǚ��"��bS���P���t�Ǧ�˯�ͳ��6�qԵ�=t���"�|!·�1��.�4����J�,c1V<�"�׊&��f������{���[Ug�%������hvQ�巳��}��������'�b�S�����\��2��쑏s��<*����D�oY��8|h�<���z�Nl�l�7��wL58Yig��$�s��̡54"�Wtq��C#&�/춭l������WmM�T-P�u?m�}�j�Wϔ��؝�`qTXP��̦E/(�u�7��P��O�>�Z�;��&���+kC*F��2)r�Z�t-~J	{e.��n��=oa��}�B��5}3�K��Rj���\�k�F��\_��	��`�5�׵/6u�gDTx4�w]���z�A5�)��߽�훘U>w�ú���EőoI;�c�&R��\VԎ�6��[�K5�����My;�m�#i=�`�9��,rxڿ��Q^
w�R��p��}�}C��_V�Ç��𱐙Ću�{jY���Ú��@߂~��X��W0ŵtO�p'=LznMh�]ݻ���
�	1��'���M孱��.�d�e�`K�v�L�x@�'��p�������������<�$Ǉ����*Sʈ�/{۲Hwt �' ����P�uŶ<�l��]�HN�B� �.�����qI�H�	V<�G^B]�w-�i��^�w3-~���Jop�{�Ü��]x%r�"k�7N���s�,��C���.o34���_S��n�zn%e���-j6a��ǔ��c ʂˡ=^����f�pB�K]z��*2�H�雛Ol��1�Y����F##60�\�KsP~BSa0#�F�'��v��r��-sr	����T��x[�;G�i�.$���C�|Cob�j~BSc�_���18�yI�'�37���3ݑU¸<��>Yi�H�i?�!�H�a�!?{��#�פwL����q�ڮZ��­�RKU���TR����y��,,@�&��;U���9��/\���Lsf/c��i�q��� �<"�fn�n�	w�^�DJ�+�T��T���hH	�p�����+q	sw�� ���+w)�;�E�G���&�)��q%�-w)�&5����a��X;{�Ƒ�燮bw$��<���jo*����_}�Uy�>�N驿�?�b����E��U�ӷQ�J�Lɳ�|uvS�R����/���➝?]�i�C��e
�hÊ�*�z����J ��R]��'��� ���ѬVڈ���^�v;7GA�QbuS\��[�H��Q�X�Ψ�����s�/n���Uj"��j�5A��~��������rbNul�keaJ�a@���~*	{��jKh��]�fQCЪ��լ��&z��>�<5�ǰ�)\a�GmN_����T�6�:���̩��3��C���^�]��p������:ytyxyE\�b�+�g��'0����k���2��UM�v^�e#��6G��P�� �b�:�;�D��Ņ���Ҭ/"v�DFƞxM?����~����~gv���%��O#N��􍈨~��,���Q�R��;d��5�M�Rʦ-����z\z�sP�v�f�e0IT�4#%���+��)��X=x��T�B�c��y���J��um�_5�!�m|���Ġ��K6vA�jm�b��w Ƅ8X��<U��Ju�'.�m��fTe��s_C�t�O+��,g&�d�P �m��cE�0����C8�+j���h�3��s���W��-�p)Z�U�.�A9F-�v�W\.��;z��4� Q#�)�ݤk�n��(rCj]є.l�`�.���sv����e�{-}'�g��-��7���8�o%��vV0�{�M�;x��*�Ζ�W0ŏ��A�T�&%�z���ÆU���J��[��̵���݇u٭�6٫D�Su�1�:�%Y�����j�L|�t�;�3E�T2bhS�2蹿`Sw��PG�&Y��s�����5#����}s8�) ��\
h}�^m�ӫ���b0��j�<5I%`�����%�d4&^�ʸOL��::�N���W>x��Ą�/���Lu� ��D�|����Q�:�/*7Gn����]G�Be�F��tky��d��
�v��#�)���h�x"����PZZ�����qY��k]twX죗��L;E�'�iVԼ�RӲ��WQ[������]��SoU�Q�j����}��=�ѻ�w��ܩ�Ji��"2&n+�'K���.U�mT�4R)�Y\�r��K�4�N��c���z��ڋ(���5GE��_��y��F<1���W�Yӥ��i��o�;Or:�2�Y�L�ɹCd܁�ͫKc ����L�M빔��L���<❯��6��)�K�]6�w�R��c���Z���x���/��c���%V��"���dR�R����G�;|#���"Y��I������W%��|;��f_p�g ��F�3&�� K��,�gPm��ɬ�[S\A[����;0S��x�.x����+�Z��j\���}j\�B�-��"n��
*��"{Q�s)f�ǻn-�u�nD\E�踷�ι����H	��[��*���U�R�=s-n�[��LX����x��B��Zm�� yE���|�a��i�v0�;品ۀE�
�T���M�4�![��=�0_k�	}ыW=���֚W�կ����x%��9ȪŴ��[�O
}1��×�^�M�y�թs�<Eb�!iY��-�Mය��uF:�I�p\נ1�z�>��<Q<�z��a�kn����D@�6����q��}��ݠ��޼}�B�X{F�6f��s���՝v��H���W+�v�u�&z��VIZhX����㼶Ҕ�0��ݓ3�n]�t��wn�[���K2��Z4N�_����]]sss.Xp�S����a�Rn�悺��t����Zz�����P"�^�G��dA�:*�WSņ��FeJ�`A�|�Q��k�yu���H۲�)�i���
��*�#��Z��9ld�U.,F�we�%R�!�=�WV�x�U�;^�8�<+�Cn��K��������`uK؁�YG�ۖ�w���vH�����.>�Y(X��!#a]�*��v �D�"�ҷYB��ޥ��܉�R5*4.='����U�ϺyR�]��x}4�SQRwǇ��y[(���$i�����g���S�wɑ=i������w��D��rיOT�>w#���}�a}���t	$�"8�����۾h�Hfl�[�(�<��W�ܛ��_���Of`Y�p���SQK��ʷr��r|�䟜O2�{�5�:�'�|��/|�T��)Z|۠���>S־]����"㛏�a�'�K�^�z8A\�y�/ȏ��w<9ȭ,rC�F;���5�k����U�� �+�r)-�t��"j��DS|l�¨*�����B����"?;���u���v��չ]̊�{��_;KH�	�H2�)N`�y�"�UQq��qBʲ��D��B7W�:�IGIZ_���b�?`Y���'��Ү������c�5���E]��^��M�Nh����Wˬ���+T��Im\�i^���Z�&H3���UU@Ƣ|���,~hm���N�ŵ���2r}\!N�H�;��@Jl�eL�X��F����DKP���Z]V�\�,����"��|�R��rV� ������.�t��]<��>o}M�kMl�)¼�mOe�V�Rkw�z65Q\��T y��n<��0��YTb	�{��)k�L�f��!�r/� �%:O�bS��%��&��s�O�p�� b�ڲq�C�P�.ZN��n�u(�o���k�e�)��P�Gu*I��Rr��E*�E�5]���Ѵe�˥b��L�p�� H_r���C�;�r,�*�t3
\u?���y�{Qi�W�Fh#p��5�;�iw�q���}�M5�cL���VM7v�֮ ��K$k)|�	/�.$�Z�ƁSv<�9R����P���
!�k�ꏚ<��6dN��L	>���W˃����Ρ�l�k5�Z�:���r�n�6�*=��f�zwf�v�?5g�O����`���P9����b��KS9�j�=Ϝ�:'X*�k-rz=9���|�?7����{����xߎF>��n�G~oӿf^���?+bS70�ۯ�T�����*���gm��}~>�o!�/y��}b�U��񛊖`n���ΧX�6��r���Zpr��R��Jn�����P��Ia�uabv�����H����M�K.�v�I޷����:�����ꯩ��E�:�����|�n}9�~;I86���`��	�F(��-�Q{�=��$"��[x)�����f!;;)�f���uH�J�u�w&����y)fM>��I�]��5���`��P�f�]�(�P^1�.�!����SRS��n�8;��3,�/u���(�%������Q{�j��\j��<�������D}������*�}]c�+�:n5�i�Y9y0�^Gwe)��yrCq1l��6ʆ@�t�a*B���rb�:# wDՅ~��@#Mo�60<�Y#��s,��ϭx��g��w�
��Tn��^�`�Ø�yq�ko7��?UP��{uy}Uو��ssTd.z�� �ɊN��J�RaMK�,�)k���Q�n�B��N���ܩΙ'�F"z�9�d�G�m�2�=�a�Jui�	T���GN0l�my�ѵ!v�p���'}��\Y�����^�C�C.�v!�͘i�I�y��_��R{%��ֽ�X�S�[���A�Qt���F���DcL9	��T��q��m�}�H�uY%ub�q�<`G���M�YX< %]x��	W9)Ä�+Gou^�~\�)�1ר�2��M!�T�pw�䩈�N��M�{��]���8V4����7; :�v����Sݼ���k��IAݰ���YlS�Ȼ��XڼO�XZ���;�8
x�������˶�٘<Z��j�����Z���Z�zU(�e���5�wT�����
%q���I���y�.������"Õlf�5�}�4wG����ȁɤK�j� �� �;-�;�v�5�x*� j)𽺵\�c�5t/l(��,�%��y�+��#�*���ک��ô�px��nC�2���3��szW�h4����ͽ�E.�Q+\u��\��%���E�x#�y���;��_�j����F��A���2ё�0u��Գ-�;h��:��|�bqws&3}�Ů*21|s�����s��p�]J�]tI�s	�|E'�ٵ,�:�wK7�,4]��P��m��ƅ>�[�����m�3����%v���&	b#�(�s���/{۲Hrx�+�y�yӖU���q���;��b�9.e�˱���D����d!\MNe$��t0�h+�r�"�oW0�Yo���k�݄��PfPO~J�!A^i��t�uC���� ��T0��NV����my=�{B}p��է�kW;R���yHZ�0��,���<����e�v|){�pb,��Zذ�N=���~خ��҅Jd~���nw��e��龻M.�Fȗ<{�_����S 'sj/'rP�o h+w���{g�s*E��,��N��R�r��}W�U�P{��D3y7�<K�YR⛼�oe;�"�I��2Zw�UTυ�^�z{��g��ŸC���
�m1��d�k�%62"ѡI�*9B�c>�M&ͮRb��'v=���\6��E�W\�4��ex���<��Bc�bS��#[vs�H��4(nv�\ȳ/v�"�Oز��J�p�P�pW&��?m�P<+�׭U>�ը�nsܵ*8M]b6��b[yu��OH� �@̷�>̶H�L?K��ȴ̨�]p�8�"L���w\2ݓ��o%��jQu��)�{�v|�+Đq`�Ç2l��������+'ko_Ffe��[m�*G6�[�)�$ڝ�Vb��ZPX֩.����\?k��
ثw~�΢a�R'NO^���Lp�nى.�Ű,|t��ß,��T�Gs��l^���m�_�^ɮ� �9���G?�Av-�ps��
&�WGN>'�s�PK��:[M�M��q�F�ȳ'��	��G�W�5�������m�?e�Q��<|�4U�Yt�W�Su��Dӕ��������,Ľv8g��h�^FLV���uC',-�82^1DA�Fm#[d��kK����*^��s����Z���K�
���,bvW�G6�����#Ji��t�}Na*}u'��tWJ��t%�1^�W�Y����pa5�jkb`��}M����e�]�í�rK�v ��MmOT�6u�dN��sM|<�M�M��xRz���/�c�C�"���DS�:�G�5�O���`W����fEs���g3�WA���j19D�bF�c@�H:A���ӷ���H؊��Ȗy����5��؇γ�F��,��{mO��/^����;�S4W��L����p�{6������v�3·�X*��"��r�x�ϲ�>=�A�)f��2�*�6�5Oi�!��g�R���t���V+1)��	I�a
.���윟W���	_�b�>�BSd�
x'l� ����Ȼ�z�!Hjd/:h���Y�ujiM'�4�.���� �A�vl��o+��=�D+}�ث���,�#��q�d��3L�R��qo�@r��I���I�q�GZ�*3a�CUs{�zp��h�\��Jt� s�����wO+e�ϕ�k�_�G'69�y-jj�wlP��̄_K6R��Ǝ˰RJ�;�RN��9C`I@b�Ú�1e�'�ӱ�uڱ�x��y�s?��D�S���gh��a���=q�O�|�{Ȁ�3��ro�T�O�5���T��WŎ(�n���f��{��<��e�d�z5]2	���M@�wd����
ώBxϦ�p0w+J=��.�V�n]�
r��z��Wt�h�Ѩ5a��qƊz�q� K�oy�]��9־�|���}��߫sd�/��@cF)�|���a�Ϙ(於����7v��N��=��P����Ѣ���6w=��.�a'������^C�z[�G��vdN���L_�Yzi=i�T������7A�_"j��=���Ԣ������x�"r�W�~a ���!�]����.qU�����aE������5���z}[~�q^4)m������8��[����S��4f}Z����t�Tw�|�����i'Ǔ��	!o TQj�~�H! ���G]�0�����(��Y�z�_<��R��5l��罛�o�f-<�£��Y�/Y"�,�'^-��]J);AyW�e০&&;�Xً;Kʤ?eR]���7���� �SdS*��%>�]��9���?j�O����<�@��!�Q�+f����q�6Vde��#wkFU�Eo��h8B�d�W(5g�b�n@�t�9���q��yf7^�%n��4���3d�G��L��B_Z�� �ȣ8Ͼ1��g�Mz@�	��Q
ﮢN�oLXP�-n[� ��J�+�x���7+_2ݞ]�5�Vh�"JցxQ��2L��GSγ��<��8�)����5���fI��^��-i�]����u��
p�;=LWJ�P۝�/Zo��P��J�2��Mt�깒���
E�J!��o���xz�z��'B~{k��+��'Y5xFB��A�9/)��
V��
j�,�)k�oϭƢ�I)�]�mW����f��L�^ܗnd��?Bd��ħW�V%RN.����b�f��t^Ҹ��:��Qm^q���1���a�e���CH�3#��&X�LR�l-*ԹO/�¶��-� ��1*
������}� G�B=�>�!?W��^���޾�VY��l����f����m��+Q���ٶ��x�1��vk�]����
�;U5�wT���s�x}q�q��!EkU�ጤ7��s
�����$�i��d� ri�ڵ+9���gB�Tqq��GlՌ��F�p�s�+]@ĝqvJ���G2��u�$��}j���M
��X��~����uk]������|-�  tsu��^���Q+\u��\��^��U���	����������S��^c���P��L����Գ-�Û��@�~��X�j�x`�m��8����^f,��]FO}\�b�ʁ^�@���G�O��S��[y0JN�����Q`�^��+�|Kdf��Ϭ94ۑ�KZ�罃W�+
�m��-�՛6v&���LR���13�R�ip�Q
	�(u?ǺR���7MN��;X�-�1kp��߂Us���'M��;� 敥��W#jV�.f%���$^_L<�_گ�dʹ齲w+��o��Y��q���tE���Q^Q�|<�F~Q0畑Y{���␙h��r���Zf
�/��R	@�4�F]�l���m�`L���w��-o4�,���x7G�T>�]�˭Thv>�?f>������~J�!^DךE�Ӫ~��u]�(�m7S��Tx����0=D@9Hs빮^ʨ�]s�-ly@X��0�*�t)X*��z�l��u6צ��]Cv*��/��Z���li�	�����cY#�ږ�����&BeV�
N��%�ϙ9�T��|����w�/��O���fMhh�F=�O��Ю��#�O5y�	Li�:�#��܆��m����s���q��,R��]�V�b�O��)ZL@C�@k�+�x'�ƀ@�仕���l9���Yy��9}�Z�����]g\������:�P3-��#�K���ժr�_�<�ּh�7����k�b�i�$���N�#0��^�l#�<�+L�"�tW�Ë�����Z����t��l�����ʎ�
6҇qOK�����9buIw�#�����-�G�����N&��R��������y�y�Y����Tv��wV�����;��2���C�%��r�i�jֆ�PA��������+����C�n�>2(���Y\M�n5* �O�[�ɨY��{o�ա�:br�yH�v[P=9p��"�.��g�|�2&��oK\A'Ga��<|G��֑#X���y
��0,t���Q�������w:�yF�]���]�^n��ԩh.= ǃ�= �4c����~���Z������f\���q&,T8���Ws�7�K!T��޻�vG��z���ᯊ��Z��z��?X�"���<�X��XV��	�N�q��z嘸�6�όg��`<�yɊ���9�]m�[��o]\�ci5����f�Y$�Xc�C�"����:"���Ǟ��9a֬��3l9\�v�z�>6˄M]v�*��K	��F�cD�A�$ !�˶x��O��n���Q�[D>�ܹ�������J��h��&�_l��^��:g���&*̦
��PFL8~y&w<��XoS��k�E&`yATg�|bb��z�U>�C�fچ���o�ˢL7CB�̨h��TN�F����<t��_�B�/"�O֦��`JV�"��(���t>�!#;�,��ָ�ڇW��g��ś$2j��4����0<��#q��k��Â:���cH��)y+|J�ܦ(
oF��J�▩�U
4�O������j��D��*�&�9&�����M����o��2�z�^Ҁkr��2�������.G�gu�(����])�)b��	�ldy���ݫ�:X���x��=ZjT�Xw\�y��b�}�Uo�U�<��&|������MNa���I���=<j�{J̍TW)4�\lSwѦ]i�8k�,�g)D�zE��8m?b�\r�V��Wl	=>�4i�F�V餲�Z.U,��c����Ջ������ji�,ʶ��4v]������R���'(t	\1Qa�#lI�n�&��)�eйk�z"��}+���1��ȳ%�S>�M���'�c�y���;Fw�+�@������#�zQ��(d8=��ٸ���Ӧ�:���Y6�$Ud3�<��Wu�ײ�<���\�����gd9H�xQp�=��T<��Ȟu(��+�fC��z�j��O�c'+,;X�)9k�d�̨�x��6Pؤ���AC�i|�b說D�X�X�֙�-М���ZhZO	�s�Z���/G�Ι[a}l��� ���ޫ|Ή��Q����U��Et�G�C��W����rC�R�S��	!o��&�N��/oP�걶���w
^�	���	�f�s���+4���i4ߒ�N�R̛��XA�0N��V�ښ}���A���L���4 ����59�z4�;��ftT�+ ��u
��/Kq�Wh��kL��
<��/��� �T��}�]����k����3�5.�4���4�����jp��C�ΪWY�����5ؘ��P��a]�/Mj�댌��e���\�`m��{��tn«TU(>���V^�|�s��WS�V�̕fR7źhM�e!���Xk	�8���8�gD�����>���7����R�o2��*U�rj���81[ �(-�[�4�NV,wy[�9��ٜ���|욁���C�n��i��4���p�0��j�Ð�:\t7�hy�s��t���t5�T{\�J���h�#��ʋ�����$�b���p�1ă��_Q+5�4�ެ�B�����suw8X\T�̭w��p��cybu����ڋ ��U�غ]�R�D�˂��  �;�u��oi���Z�k��c�V�vtz�˕�m�t�p�vH/������z���*N].��],,>��չgo�7(�У�ڻ���T���5ܻ���j�ܚ�p����&re�sNYKo.��5Ko�чt�!r��~�L�Jyp`3q�q�D�-��:���ݚ��GL�R)v�7L
��_c�V*��m�\8ږ�v#�d[���2����ԑm�w��GVf[��5�eΫZOng!�)�j��ǖe>ǎ=�]৪�c���9�su��U*S�����D��ܡ4�uh��rWټ���z2hէ���%=�^71(�cEw@{lX��,2\+e�tk��H۶:K`�6���V�Qa��F�G�ܫ�Ϟ�F������*08Ą�aV�z�Q!�_2uuy+���&ť�����9�k\�U�ƞu�h�}��W�;���8:�*y�D��ң�o!oU��d�IB��.ɮ�nq����V��s�\���/��k�����9�sk9��\z�ӓY�.��1f6_]H�>n�bM�����v�B���}Ev�;k:V��r�pl�н/�;g�k��q9 ��3�РsZ�ʮ���ϸ<��n
z�b���isU���p:��a���}�>�e;�G���͏�o�hg$gf���F��p��
��;,�r�IF"����m���x�p7�G1<���O)-j�Q�5q��կ74� |�9��n�A�LVav!	"��c�1a��]Y�P��=���ɘ�ou�5�x�V�VWy�'\Kr��4�dY�0�^�p���拑���u���^�t��
�Λ��ޚ�k�`�U��.�r���:��
�z�/��x2C-����X���R��T��ʤ�
8Ǳ�L綉��Թ��,�C9��T�`Xv�e�|�F^���z6�ڿ���;���h�����*J�>��"DZ`��}�ۛ���0�������l!�ڃ�9æ��x����u^���s��#0I���ɢM��J �y|����Xy��OȆ�*P�E(i��:�^㜺(�!�(�=��ԮaԢ�D��)E6/�B+�hy'�t�	5D�׮EC���$���r3�{����XU	%��磝"�L�3A9$%,����J{�ԫ3�s�K#C�%�ҝ����N�Q˻2*�T�G�9x�W��V|��QK�M������>�z��S9(�]��L�B�ӑg.kT��wv��Y��qz�f���L�a�P�"�#�rȢ�ξ<'�]��˄zUQ!Z���!r��t5$���Nl�"%wiTI��h,�2��X�J�"�D��q(�I���B5]s�K�Tf�wO$µ/q�=.�\O=י|��j����%��Ћ��[����;�Կ<O�up�-Q*<����z)\�����Κf����&�;�A%�(��/�$~2�q�D�%��TC���zDEQ���>�����<h�+~�qf��<�v�kI/�o^�r���
��2q;�p[a�L�3�&V.���.�L���߇���;��k�.��"��q����$� ��O�&&=ˬlŝ��������H�d��k��T��ۏ��?LPx{����#TR~��);b#��9ǯ����?l��ri~���e��P%�̦ys!�C��MA+���yݶ��L%4<�����l핧}�]A-y��k0�])���Thr�;m��'��a���ʁF�����ƯeEÚ��Fc�-4槼�fE!
�M���5Es�dk&��\��2ǰLRux�
VRaMAu�3�l~�}3բ��OGw4�U�k-Q\ =??��ԃ�.Ѷ��h~��=�1)Մ�\�mb�s47CO67���tB�=�"��{�����vH8��!�{�]�i�b]��J�*��֎�Cv���9��B�H6Ȣ�8�@�����N��AƐ!�O�:�_�d&f��2�=��lj�����׫f�X���Z�;5�5J�+��ڑ�;J7Åm���T������k*CV�[E�P%s�W�ܤ���O{%� ri�ڵg�w��)�F6�s�����]�����)�J��ڷ2�t��`ذr�k�0ڕ����]�Uñ��&U����A����:�f�^|i�Ka���t��Sg
�8�ɵ�#���]��"�:ʑ��4����Sq�4�x%r�أ�2�6I�W�9v���U�Bf#�|������ЕίƮ��$닰	TXU��e6ְ����N�-m���s�Cۛ^aq�!a�CV���`smv���%k�-е�(%�ʡ�З*>WD���pن�Щ����3?�����mK2��Ú��@�~��X]tc<�)�.`^W�`#%����ܨf�{X�R<���z%��)���2���0Or�݂wL~��X9^4��3=�L]r�ؔ�IK1סŴ��V=>�V���_~�*oig��O�]Fu+�7��u��N;S���s�������0�3"�x����� ��˱��˞)�xlg�`NY
�4�f�۴v���<�U+(��zצ�s�wa ��]��PDך@��t�u�m뽓4���ݹϨ�������|��k]m��Y��jl=�P\�]�-]
EI�DXNf�4i����{3ۛ���0��T>'�{"cH�0�}�yڷ��J��KsP�Jl�!2Pׯ`�5��u�4�^��a?���X�����o�.	���S�^�C��	����[�{���	�:YY��C�#CVM�
�\��w�Y�x)ʖ(��W,��!���f��(.�,{����U�s#4���uj���(��2�)���:
��l�r]�0�t�kydS#����r��z�ĳ+�/X�� �����ȳC�O9�j#���R�/�Br��UW��;ml^����֯��']_���5)J��l�=k�<'�|w��c؇H>pBz��*v�I�X�=�z]���nW�2��^'K��L�����Πj[�xDߝf�d���Zz�[�٦�0�u�6�֑*��P�;"���jQu��L�؍;qs.[]�k�k�ŷ�8��j�o�#���)��-e�Rr�;JQ�=/E�>�J��Iw��}v�Y���),k �x.���Z`���SI՚�`Z�t��qTa�dw:��*������fF���muy��ʐO��`x=#�>#_�2��ښm]2Z�(S�*�@G7����t��=g��=�<��݂^��Z�Գ%��:!z�PѬ'��'�G-[ht��̫�2�U��������|�>�z��j�Y�z�p��p�4B.Ŧܽ����~P�6:��9h��u�d潻!�g�Q~��=$= H�o|�������jiH����k*���Yk�'`���q ��/��3�, �gv����a �r�v ���y){\��1����"�F؃-&nT~>k���O��u~3�$�T��P;��}2b�Ȟ�oa�-ow4��1[�syt�wb���8@�e��B�J�S�%��W0��ۮ���)^}~C��
���f��m���.u�� ��z����UL\��G�>�[���ĳ�F��度-�s�Q|��J8|7s��?W�����p�8�6)�*�:�Z�˸y1V���N���r��B�X�ck�ǲ��߿07ޅ炭�醨ɓ�{�(�l^��`Z����ٴ����F������c��xl\���&��j'�gu,�H��n���}�v#�R�&��i=�Fu��|������|w���%���Z;�^yTsś�λCt:�G
�U�^~��&%�t�K"��U��P%RQ���d5���/�*wbDzN$����E�ۏj���t��.��t�e@�
�[X��澾��3�`��=�7^]�[��ֲW�ɢ��6�S���`��%C��u*I�9�NP��gʞ":��X��
skp��#�|�˂���!�G�������A��.4ϕgC1�|vZ��������k5Ow>ǐK�h����L"A��|#��Cg�n�ĝ��:��ߩ�"�:�糺w+�b������^�vԧ��g|�#Z��5�@!n�O-�ۄ�Ⱦ�Om�f�TM�+AN�TrR��Ja�����y��ݾU�GM��m��;�n��`��i�h��ۢ�;Ā���.u�X$,)�ԛl�;�Q�z�̷Q��H��$c�QB/�u�D����у]�W�vb���9Ij�.�)�D/*���;�X����v�M���q���z�*�M��ƻғ��FM�ߩO��f��ͺ���;MBl�j��P��������Q��;[����k�д��Ʋײz~���s�~[a}!��
�xR&'^��WCuU'ٛ|A��;:`\<9��a�������Nf�+�BB�*(���>ܽ���TQ�q�ff�s�j��gg�坯%�&�k���/wPnyp�i��Ӷ�Kaщ�S[^sl`d2����.'Zԇ}��H��O�c�०�&;�^�Y�^���3jn�I�����Tl��hW��ڂSl�W�v��y^���9R����`C���F0��$ZE�V��U������جl�H8��1d��Pj�Fq���6�S:|�x<��ϡ��fqV������t��TF�T�`��ثn�A>7{ ��YYP(ֳю�ơ�s�Gbz�{��xc.��<	������Zr���;o�sן�X伧Db4)XUI�6����ɨԻG#R��V�i���̽u�q����篠���˄tm�:p-|{�/8��9��\e�Ɏ�K�D:�0O�4�ܰ#8ݨ8<+%��r�T�"��ojۃT�,9��*����,9����Q��PïD�iɻH�y@Q�T	�DB��ȲMiu1�^�ɫB}.֒u�ɇ'5r��p^��Tg��^�)��=�oR�	j��~�Y�`����9�).΋��*�őm�~�g�<w#!����#�v���ץ����d���=�szG��%a�����&��3e�8|��� @AƐ!�O�:�\��p�L:�+e�)gtQܼwj|r�'�Ͳ.�8��E�d�"uD��j���ԇ����<o�S������8kǹy�ī(R���U��-B��O)Ab�&$8-��jwļ;��.F���s}����|B���Ӻ���FjE�u��%QaV�y���a�/vY����ʮ�k�A�ݛ�h�u.3�����sH�a1�ͺ;MV�V��[��{�LG�YZ��q.�]\3�6*:�	���PK�����J�z��-��,9�J��A�fl�jg�^�V�m��\��!��f��
�b�����@�y�����$S��[y0Or�3#��Փ)�՝/I���q��]��f,l�$�y�u�
�	��^�=��h/qƶǶEw`��힆S;�_����dܖ��,ÆdY�����F]��tzu�&}8�6>+uX�Ga۞w���i*�7���ǃʻ���Ӡ�nVo�{�<u>����T��7rإD�L��{ޤpoe�^�pbe��J��V�hȖu��<u��]�a���̇��wX��Tw�6(�t<��##�sn6�$��m��)���7�R�p�wZ�EK��d��C`��0���ڄ���[2���f.���^|�J�!H��M�Ӧk�Ζ�c���yo~W�^go�+{%k[��0<!�Ao!3*˭���Y�ږ�<�/c�A�WB��\dT��Ɉ^J�����F ��(�j�䧡�X����s������Y��EФV�l�|��J�EǄ���cj�ؼR-M&`J��[HN$�p���^!�"�R���Y'�̋�%�9K ��y��뼔�	�!)P��iXŗa�*�$�!ء��ҔSX��lL���QYs{=ш���0/,5�脝pc�:���W�T�S�W8��P�`8H�p�k�{�za]�O��2����L6܃Q��������O9���:����4�4�sw �����~�?4{��miD5�!1;sA��5JQ�=/޳���PXܼ���7(K��(�ix��!'���� ���0r�����6����:rEo��0���-�_�ؘhP�X�������^�T�Z8-#�F��Av-��bNu}�>4x�loY����#�4b&�Y1��� �FU�)wCLt)/ڡ�m��##�Üf[�Dt��jx����5���lIu�:�/Wv�gr�l��>(t�Wfh�f�f��ۭ�xΛ"��:Gt�D90٘����Z���Z���=�y��i���'+�,>���s��K�1̼�%���8`V��&8=�8��f-���f�ko]ܬލNՎ��6�b��3���3�ׯq���,Ƽb�;�������՟��?hT_"Q
I�/�W��Ec�|�b��m��E��Ǥ������9�=������LbQ��q�v]�7u$�j�u!�p}N'�5Յ�3�,�4��^�xz&Ir2�XoX1����o^_'\Ư�(j�2�C��r�S�9�s�g�Rnn�R�a0:��_3%��]��N=���.���dV�.�6()�L�p��]���'��D��[�²T0��2*y���óҙ�f��֦�&�Q�Y�i���N���Fh.򋋏�C�ܟ#펈��g/w�0�S�^�P��d������E��M<�[�D@A@�kK���()R���S�g�"&{�=aO^@�B1W3s��i0�]'���+T�5ߢ:.1�{gO�Q����)�U�y��j]#_��n1a���l���6�ڎ�Γ��ħV�ʊT��҇M�45���~���P��Vc�Z���6�=���hl=kYE�TB��?^T#C����^�l���-���5�ǿ{U��b�k'���=Q�t�29���qĳ�f�j�N
��]�U���iR�J+;�ɐ��0=��H���"��]\R�d����>�"��c�� Ʋh����C�{ �B#�z�7g��Z�^�[i+ڎ��Q8*���B܃�fR`Z�1e�ϸ�-��1�nc�l�ry����g�{J
v�u�'V>�Q��մ�T��d^�)��j-#��$��am�C�=�L5�cL���}����Лj<񚼽w>ý������:�a�S��T��$hkc�@2���8�Irƍ��YWÎ&w���8�f�FMc_t$��b2m��)��&��t�9,WzϨSK��9S�����;�!_$N��ce�Y#s�+�s�a�Ʋ�'�Ӝj+����8B�UJ�dw����D�V�F{�d�➇Ĵ�����:���������%�H@:��M.+J��f}�ór����g����`zQ����>��ف����7<��I���j�3G��Aٳ:w)N�+�f->&���,�4S���%�p�)鉉���6b���
�i��G��;"jz��E�+��f���j*m�j����)����)1c�D����V!S߷��i��ϭ���p:�.�r˥�ѽS�?��α���[��k��w�[,���qN�>/rS��������-��%X��2��a���s�x�e�7�� Moj)^�imp)�muL�!͋GQ�8RO_7�C	��m\�6�{�H�ǘ;�_��7�������$U�A�PJ�(ų�l�,qL��Ô�wz,F2=1�BW�f���YK���L6g$�b���O�c ��YYW�5�������j�b�,���2*��3����.���:9��H6����tL�VzK�I�=����Oۥ�.+W�f��U��]
�		�n��[JH?m�~ʜ���{��i��V���ޣ^�MS���|;2A~t���
@�~���Z�Iu���ƕ�'G(<Y壒)7J������]9��!��!t4����:�+�(�]i���ꞥ���)MԸ�:��"�v:[=R�@��o���1�]z��6��ʙ�b���*�qtMJ���S�Q�e�[e��#��4���nӮ�^��Tf��;*��+]��L���T��d��{w�"�D̰#�7��N3�{hv�T,�ڲ~1����o�,�ؙ�"n�0mrX*mV�.�ޤ�mm�Ɩ<6L�����5$֎�oQ'�.���O���`����:�,�!3��;�m�W�Id�]��<�.MoT*�3�������b�u͚�(�3
 b	Z�*��9�3l���Z(F3k��B�:�o�7R06��f�%���@�t�����*�����:\�zgm�3z�j�'*،�6�*�g7�̍�}�l��N�в�W[AS�f&��η���fgAN1��OqD��=}:�����R�ك"Y�Y{��B6�^���Y�	8j�xr9X����հ�19g${-�#ZEX�N)-�5�R4WL���ct�!��"�u��wZ%-��x�e$�)����W�Aa�j��={շ���}�i�����u���^��I}��jXy�"bt�_hZ� �o>�,���Q��2�V��� �L���N�D{N�9C˴i#���x�j���W	pT���巡H$P-X�T�̣f�������`t��̨��������}i��X�sYdT�>=��o�jzl)�_y�[6-�y{2kƹJJ��e��jN�恈�gv���,d�>�������:h8���^�v���"��F�e�h�L3`sH�d��V�mhFT���Ei��(fZ]B��v��	4�]��Õ��u[|�&�2���.k��������7rqQ�Ύ���G�6����Ë�%w%`f9:���ifҏ��O̻���dE���_zk*�0E6�@�m����N�\�£u��0��qvᜃ��겹\.�γ���s�k)� T��6�,u�*�X�u�͈��9|y`��6�E�2�N�gH��u�Vm�b��>X�0����-μ`}�/�]b�JP�ճS�s\��[�����Ĝݑw8�_|�5V�"�z�t��;���|��A��J�2��D:�l9�b�����R��mv����C��g*|z����3Pq�>��W"��!��뼻U�0�'rl^���.1�ܮ������;���u�;��4r�kUB[��Eoc|�qwv&-���+�u\�	�Oj`чrӪ��}�o��W8�^��3k�	Md6LZS��p�V݂u淛�SE�
jMyCc�L$:��_=����" 7�m�P̋�M�6Ü�$U��+��P$nV��B�� ����s���{�Y[��7�.빘n�%F7bؕ�$�}�헂�cm�'CBp�a��p�b�k�Y]R�i����C��8,w;�dy)�����C�Bb�4�w�������|�bxa�g��9S+l*�9[d�V5Y��gd��7CW����U.�`ɨO�$N�
@��0c���B���ONR���˩�=���E�NWvM�+B�p��S���+�0�Ժo6ྠ���z�2��[R�ERiʒ+{k�z{��K���r���P��q(�����<�|�TJ<�p܇�N?4����_]ĵBN�QDzow<�y^5#/R(绎=B>�V=�y	V��/wp�L���^�U\��8�У���(�%Z�B���q*u�"��0����#���%�d�ژ�^K����=]Јs{�'�e9�wWs��q�:ޮ�<��y�w�s9��QO$<��B�<�������ʨ�冹 �a!���y�^`\�J���2J5��NF�w"��_V�9J�����I#]�D���E���뻽D�"���ǎ��B.L���I���U�L��������DSף��+��fC��K�q��*����U=G�a���*���BUaʲH�\��盯(�Z���OG�X��#�,�=r.U\M%:�MbW��)�E���:�/wry�{�y�]��y뮡|�B���[��%�������l���*�ƶ�-�yN�n�w\�۔paf���^')l��l����]������vu�#9ZŐm��;l\6��9��������M��c��!��{e}��x\����[C�d��rn�gb���>�8l�;#�t�V�`n����Ψ�+2Xm6�2�utl�Ȝ���r�h$���O^�s�ԁ�"\�����6��gOXh���b��;�Fe��;�
HO"�tR��r��>
j��5��ȩ�3���@��E1w��3Y]�s���y���&Ƞ+�7v>p��n�ؙ����,�S����* �Ty�2�ʭ�@FEH�Im�AZ��<��c���u��>^e���TJ�fG�(?:{';;��ڹ
q|n<Nxj4�׼gg����H*u� ;yq.f����$��А���{&�k�z�3i��z�����f��tw��J�ɭ�庑V��[�h��Bl�Qƚ����=m2�F�6�`��#�RV�W��<I\�]>k�X5�)��a�:.#F-����pݛ�`9$�-T�*�+mgSzv�QX�ڕ�ݨ��k9��N���ea�v��V�(�����Ik��� �Ξ0M;���н���o�t�";s����O�ٚ����]n�	���m����ެ��P(J}Z���'��PJAE���6���̄��w�5�w�-�d�
}2�[#g��w$���&��������8WN�;3��0��R�V����n�+X#���ߺ�Œw�%U4�b�c��U�]o,�@�/^R�wB��i�k4�8�zF��jʈ�jAl��Љ�j�V_:��f*+�QD�W���ޔ��p�!�M���L�fN�7v��[nJ�J�����w)��'�4��Ryh��Qu�3uPf"E��ðp�M�؏S�(�rG�I	�4(֌�E�ފ�|��T!�2%a��ԯ�à�J(���nj���|��~��U�Z����)��!���,���������dn���1�v`���A�ʅ�זD�Y�VR�6)����A+�������*m�ۥ[����Ӄ~�)*�a�hҍم5��nd�.��w����Kcc� c$͠'�S�\�ui���d,��b�\�t�]BH�Љ@PR�����Ү���w 3�\ER[��|EG����j���+F�7$����t^�N�rYN��%ϣ�u���[z����
��tmn�7h��9��*��"�$|��䮹�S��`����Z\[��m���&���Y�	�ʣ#g����}&���y���g����2�K��wP����t�C�(4�	z����ځTL�IU�>�����2�'ס�̤���e�/@ӓ�-��b v��H�ts��nꕚQ����Lu�Ⱥn�N����t!��*A��;�$�ٺ�f�vZFnLa"�f��O_r�&���e���ל����8w�mL@Ⱦ��=Y������m�9uf�ir���}��d�<ݞa�˩���5Q�ު�3B2����5�r�dt����=�kTג�]�}�X?kljq6�kZ�L�UM��sp�8"��; �4J�\��r]V��+�T��6�mЍ~�S��x̒	Ӟ!�Q�K�}#�}�iQ������=��<j:���"�+U^�6����O��������K��V�no�,8�\걈t�
ʚ�]L�`_T
�w�R�UtH��n�#_f:]Jۊ�)l����ɚ[���H�Oh�:��z���2�� ܧ��F�&��X�]��h:
����+���|a�2�������j}	
��z@!3��1pwM��.���N#�_�*�~��g)�V`�ps�m��;q�;EA�;H����.%a�l�J�p�j���q�E�b����7��@$ȶy���2�E�	�Iv�ª�̰i�u��=d��f��3-��H�U>y��ڡ�nv�`�[���ǜj�˶����zaaV&k(߻c0�YAJT�+��^j�m�ZGZCU�yakt6n��v"w��̤��Z�F�Oj/�&�
:�i��!k�eCl���֛]�hN�E=I��:����#o��r
���<�,4t�5�DCP��Kc�ٹ�G��tӚ�� �\�:A�ۄm��W���w��K����z���A�5QF�A&����v[����t���!J2쯤E6k�x�������o�m�"��T�OS�t��s#F?�d��"i~��<J�����O�^l�Ӽ{�we͙�S�Ε-]��S`_d������>��8#�8�z�x�$���v�t8E �l��+�7�6�o�; ���t�uO��%uXp�C��n^O�*���H���+j��Y���N�8esV�1�])� ��H9n:�W{���q<u�SK�q�]��[d��K�kn,�眦��lT�W��t0�!Y��9OL�b��Ī�qtH�IB]������KF�E��<cC9�Ê����0&�.4#���4c��w.Uk�D�y)V�&�8�g�#�U0�a�{������v�T,וw��d�f*m�ee�7���^oR��F�I��=��Zއ���.��c�#����zy�An򠟧�'g�c��Z�03�,���f����j��V?
����Ѽ}�Ѻ;/�$I �0���]#M��6-�g΃�^�8ȶ~ڷ�Mg����<ѱ�:=�d<�
Hh�Z�\�Eac��(&�Ɯ�yQ������h�ǅz�-��eu���ԃ��^�P��g���+���j����'����+c`�@�Ǭ%�VUmǛ�Ij�ve��js�i�(~�xv�9��#G�E�\.�X���	8
���$/D����:���^��#�@��3�Z힋�JpX4N�/w �odx�vBw̼rTܤ��Os3{5�Ք1�2����ɲ��eX����������WK���wn+���[݁Vk�-J��Ú<+ڵ*��8�ؠ�j1.vy����Iv2���J�T��Q�ˉsb��7^Y$ck�i3���ФC*���ͼ9�.��Z%b��r�t"O$T�T��r��3���� P5�y�G�N�-^|������{�$��Gow$�`��x�8D��?آ^Y60�?q�Rb�3��hRm>��#H�n�{"�\Yx�pLd���9-ƌ��hO���P#��<� w$���&��{�ь�BCa��<�s6�	^�[�#.#ݭ���-�ά`�n䪍�q�(�ۢ�N������>7�f�n�W��~��a�<�of"�OuGct=��U􌭻��쇛������]@�j�5C;�9��p�5�*���]�Ӫ<>�O�6��u(�ٺ�S�_�Ǩ�ܛ�V8ˍ��;�!��R���Π���\dŮS)�}������.��ъ�|�'wf�%e��z.,�	��4�W1B�Ï��BK踋/�A��`�Y�4�5>5�C*o{�m-�y8����{H��y�r�
<��lb�n#P�p��qr6�d�K3V.�;�'h����(٪t�v���%f��G��zH�H9<c�,��1!aA���sm�C'� ��W���~b�u��+��;2ҍ�Y!+*�UU\���E��i~�q�/X�
S�s���G��Ұ:oh�Ya��#_76���:Ll�"�R���#�f�YJ@ا2�X��s�U>�5\�6��3�BsUY�P�PY'�W�i*(�Nm+�uY
��e�uo����j��]y���U��;�Tdor
�����3ثޜ�q��L�'��S3���+��^����0�B��P��7��l�ځT	��0�I5>�nsr�Z�8ѳ[�|ۧԭ�E[<�c:m��c�{ m���$�\fND�h�Bo[_��tv�A��C]9����Hl��S��I��9I��U=��,v�;��:��N�`6ɳ˸fCf>��.��c�+a�'��͎�i]�y�7z�M>f��R.�p;2Ů��"5� ��8�fX\O#N4���>��~��Bӱ��Y��삹:����=�\��g�ݿ��*%A��$B��/�����D=��gI�K�l�+T6i�3]B�v�-r÷��s���m>�'qOͱ��~���5�ݑ��el����� �r��$�H�aye�v�z�J���f���bگv.�֩���˱�`㵷��Fu@�X�p�n�U+3�ȸ,/�n��Κ�J�\��r]k�c��5#9���r��b]�2�vm�<9A��z^��iP
��}[@�]}-C��v:��穻7���6���ͣ��F.����l����7��ݶDs��u�Y;�ҵf��TZ)OPe�mӁ�Ĭ7�y&���P������kK���1#Mp��
�ȴg��r����|�E�����ٹ��ǭ_�֌�e�%��@�+*{e(�w�8CL�~Ƴ#i���{��#/3��ÎR".�DNJ�}� hYAO�T����/)��w`�P��=Y�ع�T��F\X� >fW)�H�أ�+�#�����i�k�E��T�n����.3s:���v�X���Y�q�2�}�k�d�{s���ZpGg_��[{nd�Y+M?�)�Wu���ڋ�g�� ��6C��Q�:�q�r�ev�k�Yq`��fŷ�:4kec�g��f�B��t�l�k1pj�o��ݷr	��3��ƍ]ľ�l�g:�2D�o8&|]�?W���T���0g2k(8þ���d��3�'�4�j��NE�hHH�n��@WV�T�6�������L��ߔ�a$��=�_mH�R;2�2<�(F=�l�Sq-WV�t_�k��$�rEXn� OW���5ә��Y���$E>Kcv���$i���::�BӉ�R��q�u�1�g�0�e��:0Tn՝�3�8��tW��wD#�nz� $�.��IE���N�|xwOg<eC�Pù��a����~\k��������˕L`��������S"y��12�S�n���v6z�n0����
3�{v?o�׳����۠����Ų-�K�}�ֱRRM��h1���Y�q��K��[˅kk$U��{ѭ6|o�PZ�����'x�`:�Q��3�,�]�90xwM�uNjf+�&�i9~7�닫��Nu��]1��N���y����]����
��a{�[�!��"�ꋧn�N5)r�p��[�x�)�aX�NK/��}}�	�����7��2�:��9��m���j}O���q�0h[�#�j������9���ك`v_*��y�`��6�fv�X3Clj�'v;V��+��:~#~_3���љd<�$��"��!v�/\]��4'SY���P�Wo,sc¼��U�_D�WX�dn�EW��{��t�Ƕ���M>����x]-`�����+*��FE\�2.	�8^�l���U�f��L,v4�Ґ.i��e�q�`\tO傡�e5 �oDTʲz^�^�Hn �rH�2��M�x��Ĺ�V΁�z�)
i�4�w^��wjz��x��.�܂4��T�*��u��|����������x���td����#o�wJJ�c	+m�#�)��ۚ�F���y�}�Xq��q��)���gh� �B�i�m�)E6G<���p��p�B�x�}�v[�GپaH!�����#@�4���h�E���l>b|	�;�yb��Ћ�c>�Ă4Z�/:>h�b!2�A}���ƍEN�ܵ�q�)���"��ݭҁ�Kx�t�@�RA��K%�r�滾[ls� s�D�s*�\�B��=e�9;��I��8掠��Vy^���N��UXeX��k�a/���^Nqzv� �޼�GI��-�#�o���U�i��Tj�䛜�%E���nofv\��F�����
��-�J�:�wI}�v䪋6����dՑX3���Ʈdb��7�3'd�z̉��݉�|���gPK �T�� �F�ˬy&�l�9-P�����-g��ĲLm���r{���r�<2�}���-f�r�3 �S��ol�EPMpN)�]b܊һ�((l[�D����XL5{L-b��LYgQr��{o9�R��F�:�s�ϐ@�䫄�R�I+p�p�g�QY6
�f.��h&�4pj�[��#.�sJ�n ����t�Ye�HU��e�>$g>�Գ)��)Y܍G��I�yA�G��i���Ȏ]v ���qS��9L[��׀g�[|/0,����3Ue^ �绬�e_K��M�d�nL�����X��P�6�s�%t�����:P9b�Ϗ�ە�Y�xyB�7	uԛ�j�gb��hJ
`ܝg�@;A3V	Y֟tr�Ci���q�s���}��t̆s�w}�rq��Eǆ�͎	|Z�h��[\"�q����xNe�:�/�9.ÍK���YVΌmФ�>�̼�_nlJ\{!3F�/\I�K��vyE:%�ׁ_h�h^�;ڹ�mV;k;R�7��V�:�W��sG�+�2�%S�Mk�o\���8=Q��9ݽ��|1*��zI��u��n�J�܃�p�v����V��.��qe��f���6TVծ0�h��F5!1�Ɂf�U�֕���2�<�2�ͭ�ND�%Z�}ֻ-��6�l��\���V��eͭ ;�5����^����˦D�gR�=�'R��a�/j�& ��WD1��0�"8��YY�T\��\	�{:�u����UƔ�]��l�+9�|p�'�Ǌ,�1I��O9e��Y���èT��*�U���jX9A��~|o��j*
T# EbÊ��p�|�{9�Ռ���4����t8Trvv�)M���2n�]��,�7�eK��le�zr�Z�����h1pv#P���"gT<�II�����Q���-��LXqV�m��1K�����j�,%�v��d!�\Y09�oW�8�ђ�իub4Q�$9(u-J�q�l�����g��K��z-��Z�MU�$ʁ��\�P���+륛�a�!V�� uu�Js�qm	�%n��P�[YC'BvP����,��X�����
�����x�m �qiU�QQﬖ��\:�B��C�j,GE����	����>�q:���q��X����_b��)��ˮ�K��إv�3r�W52e�n;ǟ���SnV�Ι��lN��]����������{�_����J�]���#~Mʞ�֖�g�\�<���E+�(�Z��������<�� ���t'���"���R1Iз=ҽ����9Y���4rw3̃�^{ǹ}x�Ԓ����Ot���O���J���ܓ��A̓u���/:����
�.<�9Y�������Я+�GR��Z�y�k�9;�V�������K7w����;]�]2���~�ԾdsYF&�%���S���s��Z�y-%��ژn����	�Q[�����P�\��=W]�{��?t=�r�0��WVG��z��'�#�=�N�z��W�W����U��G\���s���wg���yE.�;��Z�o����P׸�G<$#���ҝwB����y�^g�I֖;�VIz���Yw2�1�t���0�0���(!��w��~T��:aAF'ի���Q依T:�|* ݭ;ɪ���D7,c��y��!`�3#©Z�S�꠸K�=�1�"�9&�3Z���N<�`�gQnFX�m��-��;2VrztV��^`y�j��1��f��qF�3�0��Me�~��8ǃrU[�{lx��SX��s�����u��?:��T	��
&�����oJrA�q�Ş�qE�}kU��ݲ)�W8�O����4�9G���n�r��8�O�P1�7P�7݄�^���7��\/�I��L�#o�=�O�l�#���"䃒�Uc�]v��]�:���*B�B��:��0�D�7�z���fZP����1l��
/��w�*0/U����%_�)�FC?�0���6��t��f7hs�UfD�yt�O`���<�kp�g�Q)RV���b���u��,�Ga���K��SL���u3tfT�"�ڒW��IP(�fʨ�ِnGm�<��+�~�͖9p2�;��~ڕ���,%�_I��T]�Y�����n�����7E�,M���Pb*�N�i��:%�I��wU�x�.��J\͕R�T&L��ϳm�(iH���2�h
Zm��8��Kot�K�E��QI��UlTVB=�)Ҹ�<�ɜ3#�Ԩ+mη���$�s���������v^L�N�q��J�}�mDX�r�Ґ�פHkd6�Q0� ���:���C]�]o3��~=��q_����5��%c:,A+������H���g��zg�27����"�U�e%Tі�}��@:Cdl�R;���~�^�"C+��?�T0�}W���rf�.�l���V�r�ɧ�zt�)Խ>m�]oeh×s�<s�:��q����N.m���A��a�Z��r���EE6�����)�jAL�t��{�mv.�6�J]�<�:��OS�'
&��s[DD���i�!!a��r�{fuW�MUܗZ��Yf	������O�o�fXr�8o�q����vN�^
����$�7R���W�Vs�=��/#�Cg�7@�0�̂4��=w-���ﷺ�n�շpygj,����o���H�?@�� �k(P�ޤ���y%F�;��X��{E�ٓZ86���|Vp����5��)�Y�CWml%e�oΏIVs�қ9�l�X�z^C�q�ޡ�Si6,nLn�+
�L#��K������S�/V�[9y�T�lf����f�=&2SHˠ�w��7iv����y`�.�m�l��K�,��Q�$
�E��6:)�#�ˮ��r�l�(Dvy�F�/���������C�q �#N�R�\��9�!���!�=�������*_���u����8����HI]ml�t�b6]���1�6{a���"��O���W�P��\�
�J�lT�aAe_\S���ݖ�a���vs���ZOUϮi���:
�9Y�i�'o|\*�U=(筦ʼ�[(�����g�׌�K��%�z��@=��	pcFr')g����ڈ���e���ݙnI+a*	NI��\;-�fd�0���/�Y����z�BW$d��	�/��C<�C�h����r����-7�%]L�^���(KX��Ѥ_)T'��Jk˩q�]��[T�{e�۸�zr�Qm�fK��/B�#�ze ��P�J�]F��5� "nle�� �6�p ◴<Ѯ�ǚ�W���D�� ݬ��B��q��lv9���� $)$�,��.�:��㐲�Yӵ<�y�1����ki���D�x�T��Y{����̸�3yi��x{_b�]�*�M��N<̻��y��W�ח@��f�x��oo�>}�y����(�8�P����~����͞���<��U�&�oK
ь��7�8(���⊜�7{�rڮw��O��E��{�_�#>F�{٠����]h����E]�偳H�mÅwx�F�~�V���1��Tl1��M���L�?-�5w����R׍�Cd�F�e�$H�������h�o��M\���q�"�{B��O$Y��Vv+Q w��d<�$��������y�#wgWA�g��kT/P�*�7¼��U��\n��3�$��n�S;�g.�{b�z�^we@�W\'{�^�Ίu��,���������k[n~�'�o����)�\��"�m�
iT���ג����8A]�+q��~�[���"6.�:��n��y>?cj
�%h�Q�'�o&�Ϫ���Բ����ߙ� ��{e����b!"�Zm>�	�(.�����������P���Y\8��ɾ'sd�K;OfmX�_���Ԯ=��0Ή�Yu�-��[�J�#~0�R�e�ns�	sٕ�e��q�Ml��N�M_Y�ώ4���B+*��ܭҝ�o�K�S�Ph�׈H�]-�#A��O%AJU^}�ւi���#n�o�ݝ�.+����@K%Ɇ�)�b �2;�%la%m�j-�c����c�*��1q	y�����g�F@�t�� �8ФO m�)������]��؉����B�f��OH�����`0���vy���xW���g���5�?��óN��>�[�q��<��<�ly�o]|5�:����ےsވ��)�]~�ktJ0�t�ݟYƘv�Ї���SXb���8�� R�
gU{��.mi<��f9Q��oJs"��6�wb4�6��yy�m�n��m���5�(�ٺ�v��sr}!�eI{�t���j}EPbS�4#�od.�-�k��Ǥ�/Y�rX�GB�~�q�F�#�V�� �g@���8��M�W�:^�:�:R�xV���%�K�P�_
�ԯ*���r�Ei�g(<<�k�������Y[Y]��.\+-�h�o�󛥣)YW{�X��J�]tgp��l�`5+yM:Fj��Ҹ����C���U>�P�b��&}�.��;����k�u{���N�Ww���az�HH!�[�`�#b��!����.m#����Kl��b*�/zf�4�ݳ��=qK�V��,�+)iQ��9�)wa�;9׻��q����L�F
�J�v.y2��3F�(�_�rmԌzÂ�j�%��/hJ���~����IԱ*BĝJ�#d�P%>W�h�P��em�{H����_������ް��U�K(4�'�H�=���
�e%m1�g��+MۦҊ�F��ɨ�:����Ya���Њ���Ga�3j��ɓV^y�mfi�y�d��uJ⒦��t�t�-�cg�{Q]�i��oFH�o�bv��T2�c�2��m�g�q>�A�Y �C�
�{��uϔU+�ywk:�M�h�\��ax�Z]4	���O�8�3�a���;��c�`����׸��}������Gb�Z�.��u��δRxΧ̶�=uz�%��a#����3�ZUĳׁ�%�7;M��Xѧ��6.���i[�.�e��eu]�hcC���RMMpWk����t��Γk�A��]a���c�+IԚ����[kV��Q!òQ^n]�a��_o�7���'�Ⱦ`�������Ϊ&�9Tr]B�u@��cb�{}�����������U01���#� �Q���#pҠ`����Q�0���X�=WwU��g����]aTt��7�7X�6�g!s�w�.��-�֮���}��~z������Ӆ�R���*��'���Y��>�����yM[��D��oe8��#e"��à�<�$��8$��22�3L?@�����v��[O{�z���@�v�齣�{2�y�$ITF�l���x�j���Ǘv�%nܑqχ�,�Dp�b�����������H;#cWQ�{|�%�����ƺ�m[�����%o���=U�>��Ûk(i���F;�bf��f����v��� �\��s4Y�W �^�#b�2��Z��rcoxt�H�K�I�=$�S�u䎚u5l�@PE��='y��������q�{�	�����n^�0��5~�u���yJ�#��e�r�H��?2o:w6��u���.T�-7�8Gq%<6m2T��v�x_%k��F��|�-�`0g:r�:�Xʐ�U�:���@���f��weoTt���nƹN��W�x� �ѩ%��%A#J��T�K��`��J�@Ս.�)�mm�3B��(�s݌�u�݄H並�RQ<�<���I�8�3�us[��7����<8[\H�#��*���:�)�Ը�.��v.1���B�����%�����9m��.�9�� f��8����Yq(Il�/˝�f���=���>�dy�l0[~\j:yQ��o�=;���dUe�n����}��Z�QAV웱��[��`�q�Ìy�F_vczwg)��۹8{%V�C�(Y���{�)<����V���H��[Rk�MF�=��o���'r����u#I�qZ"vG㪖�a�3
w�]�-Pj3�t��%�F(���u�d$�F��TL� �r}��$1�����fm�(d�z��e4Y��Vof���Cϻ����ǲU�;���>W媆D��2ď�Ev&vmL뻑򉁋(�B>�"3��n����2�gd�����Vjn����7��Ź��i�:�}O�y�Z�H)����&ٚS�	jQ
X�\��M���n���nop:+(�R��8�̯�U��pE��~�_�*��a�E9�,�B`
��J�k+�VV;r��O�=]����=�Lf]I���ܒ��R:Yłl%`dfQN�l?u=�3UoQ%�*����6L\T����0���J��6V\ә��:
λk������՛~��T)�Ku'��*<��=&������}sNVeZEXk%�*q�E�V�9x�H�Tp�	�^=�� ���F�O$�)�mWM/�	����7��/�t�[��xd�9C%��=lD��{���>�x�#h(yg�7�unh��3���p�sz1� ��:+���'����b�v��g���/�٦���!�\���V���4�C(?��ȑ�xz�򫪬L`Uu���Vc��lo��x���86G� ����`��y'ep촻nT�˥��l*�#,�ͥC;&{�D��S^5� �Π�q��SMMЎ���}s���A|��6.��N*Ֆ�7����`S�ц٬�g[��:��ˋ0��v?�a,S�<�� J{�W�u&T��BN���c��M�=��Ѻ�u8���QBQ��/EJ̒�N�c��][��Z���q�����t���
p0�K�ۺ�¶�;7�Eǫ�n��ή�+LTO.�Q5
Oi�j�ᧇ��;��7{vl�����,��KF�cnH�J���C=�����������!�i�s���h�!��ɟ�gЌx\Nὐ�@�-���yԂ�O�̩�޽;8�B��1��FGPc��'FxVO�oR�~k%�򨙖�ڸ�^�.�(����L506��{b��C�7�����ي�ߴ1�ة}ڣ��1FRɾ���g۸���⮂V�"͞��#b���cV���9KlC��>�����W�1wF�T��r5$2��@Y���i���4;v|���{Ua���ن����23+��:���r
�%!_I�2FS0q�6��㻘���.�q�W�.i�E[pWa�X��zD���Cj?����񨆘���ľns�F��ђj�}��Vꭜl�W4HE_k�$HCh�͋��i�ǒ E�p٦��7�PT
d8��Y��]�Jsd�b�D^m
���}�4/��?9��:�Ԉ����D������KK� w5`
\�H.L+u +"�������z���*��^�V��m j1�A1@{U�$9�Ӝ�_]��;�끭s��X��ī��\+������f�ļ�㽠%�m,#u '��5�-��ǧA�sx�\��=�p4+��5'W&�8�sY�R�ř4 �7r��x�d!�;�(\����ؙ��BK�1j�&g}z�MLݣ�����Tm������AI�V�������͑�LM )b��C�G��'���.\��tL͉:Z6kL0z��z���2,c!��됁J�� �"�Q͕����"b�+�/m�ijL�+$��	�婤{Ml�J�!��l4��`;9��Vs�҃��:��&�Y1,�Q��eO�%d��Q'����4���|��Mnց5�\�v�;��H�@��V��ϣyb}A-B^���@7h�\'.�i�@9�&9Ju8n.WCNw�ux���=�����)���=y>����V�jU7��q@�sF��j:�9��rW�5�y��=2r�����Wt�+��y��+ٹ� �bs���Xnʅf��`��E��7�>:0_y{"��B��^X�i�J�g#��AR�NV��nZ���׭G��)�:�`�d3U�<+W���`cv:�&_[QK��.��;j�����:98�i���m�i��?:o�<�v��X��ɶtҢ�uf̹������o&(�����.�Q�ܖ.����3b���.���
�;^8;B�{*X�ܨ��ci��nf>Ւ��[ .���3��Ȧ^)���MX�W�k)�tÉ����OiCAt}�l��s��u�)�{V
WI�h���ۖu&cv��ogl\v]I�� l^m�vF�p�Dd5�<DSX���Sx\���lփy�zuT�s��%
�JS�7(�4��X��ט ˾�}�x!�񍓖ug:�i�d�1(���N�;��f�N����ҷ)qhr�1��Y���2��Ks�1'� 8Q�T+D�R:eMK-�\`n����NG,s�DYgxc���"��4���F���}>�u]hP��b8:��b��ڝ��n`J�\K0�&kT�q]>����o��V,�{6o�§���A5�o��v�r�X�Z�i��˾G�qT�f\Gh3Q��v��T�*�rlF;t	�x�h���F[e���Vr�K��V�s}���DY��vu�WjҤf�J$A�o��l����[z����Y��AE�Ϯl��&ݴ�e�ڷ3z�N�j:�i�6���E`��O3J���T7V���o��LE�%W�]���\�3����0[}�vZ4\�Do�4�>�˒闡	K�>I�77�c�$��ce�eJ��3��8C;�����C��H[�;����S9�-��QAU�(qYiIw��.�IՎ��޼=�>�z��qҊ���V`t�4~�^}�v��)�����n�ҫ���>����QW�D���G$��Ţb��e�dV�4(����-����̪�]iU�NF��'�c��������P1��ݐ�Uh���7wc��������z:e�'��Ps��t�v;��ȕ'�;�Ek^t>l*�ż�hOz����!E�D��z�NI!VH�ǽ�'�i^%9y��-rs�y��9��x�<����0�\P�Ƚ͸~z��	�=ܐ��6�;׳Ԥ�y���'�9����8^�<�X�<�L7G|�s\uҢ�E��9���i�	�>�޽��V��t+�����5
��������f���'rp�Gqu��Qd���<�6�o3��U�$��t\r�wjV}D�w/��:|��vGGG���8�{��G������ݜۚԩ"T�r+d)�����q5���ő⻬Fdغ�bJZ�ڗ��fsN���.㝥�����L�~�����dS�y޸q�ߪ��T�9�W��y�)����&�w�T
J���K�=�\Hh^v�̗�L(�扣W��/���[>X^t���W�l�<���!�}f��'xv[qUk�$%�rT���=��u��D��~O݈��ʈ�n��{C��#���Aa�7[F�ٕ��s�;�b��mj�	w]OH�1�..mi�x�֮X9-�q���q}�Y�h�7B�ǒ �a廽�U,E�z��m�� ͨꑛ,6����oB�G�u��<��3u=O&�p�>W,V��D�W_�G��!�}�G1�t�I�؛�����o{dM�o�g�	��R���A��R��á�G2��d�.oy�OXh>��ܳ+���:<rʊ"A �K��FG�)�,�yR�E�{�誣Y[�x����=1=��M��9�C������������������Ʀ]X�ا2C��ӥ)VKǝS�P�>�V��WzƝ�q8�Y�Ά��Â[%�C�8s�w�Ge:�k|)L��l:m���㈓�Vc]Z���qJ�=�\J(�e����]�՛�f'��t�َ�ia}���2@���s6�:��S�����¼�:�lL�Wv��P5e�U�6�ҥ�澦��/��'rպ��X7�M���EV�@\�ٻ74��z��=1�&��ڃ�(�O�U�K���+�V������K^#[17}�/|��(+&�=&��T^tK��h����Ю��Es槫�m:�$���&؈ge�$�t��(�5^}�E�PǞ���^�-ɮ{�����K���E�t�":��7ia�%_��ID�]�\�{9�
{wʼ��7x���IÆPrH�#��-8���]K��5�-Lx_
#]���!�b�M�c���ՠWO����h��P�_���%��a���%{��Mf�]ڦo��Ǳ֨`�q��k�.5<�fd@鈠�q����*��fV��mtr�
� U���!xf�3v�[�������p�@���7L2ua��p"�u�����ཞ���?//x����d��͙�U�R�'�B�v�G�lMDTї[M[r�4�!hC���q��\���W��wV�C�+ъ\����By��2����N�݃�)[-;v��V��5�aE�����@��Tv��+���@���{�Z�d#c�cޚ���*q�ܼس9;9{�Ǿ�\��+n����<�����c��Ww��ڞ/n=R�ؤ/�I�8
����	3m�Z	�	���(�a��Sm����Z��Y<��;Q����Vl��lw��/����<��3�}�*0V��Ih��Q�y~�_3�bbbť~����ts���QkOvs!�	���]��8!i)	R��H��#��6�u ��%L�L�{�X�V�볨�D�aRd�T�Җ��+]m"��ӝ��S���ū]�f�}�=ZL�c(��ؓ۞���IP�ePRnN��V[���-�1��3s��]/�p냒p:C^#�t��'��Bgj6xL�f��Nqvf���k`�D��c�p�&lF��t���;�sjfl,��s<�	��~��khTV�R�/3���{���o�9�gD��{j�{���N^�ZZ�u��rt�\�`!�G�T�ju�<���5o��jhh����f��&䇝3�S����ʶ7.�ٴ%$����^-�<v�s=ѽ|*z��9ğ���|�N�C8"�:+kk��d�r�)n�}:�L9�1�t��9�x��"�7J�k�}�],[>�(q��iޟE�
��F�U�vJ�]�;^X^<mlO��괉���#c���ȵ0�����tf��i��\��t��ͮ�ڶ�ģ��;�$ڍ����k��o)�{�6�Q�=���ꑳ:��T���^�K��j)Qfl����ƻ�p�w{��Ḑ(/0#��0�E��3s�S���h���}��l�P4���k[�vF��:Cn�h�A.7S5������E�7�|�Q{��I�e�jU$O��I�FGPg��w`F�%aF�9�x�maÝ6��w[����Z6<r�PJC�Aj��)N�?H�g�"Y[X���1�7f�f�Xh"a_S{JΨ̴GqJ�V��-����γ��yy���-�#�{���v���ml�Y�5�XC+�@�����U��)!�MC[Xn
�f*�pu*���D�U�|��n�ٴ%u��=$t������M���F�5E��Sݙ��_i����ē)G��;93��7�w92���&��Sڍ���{�W���0H��o�bxz��������!��&��Qƀt�d쾥S/�3�7N�\�Q�g��,q��ݳ���Ќ��w �����K��"���Y���NWw��D��A����r�����>{[,�P��2#���i��[<%!y:��Jg���YV� �g"��P����ZF��w/�DL���K`|u��Ě�tJ��)*n��]:���-b4j�@姊k՘����G�h;)�/�	-n\F��<��&���L�jbE	ɽ�&�e2,(}��$t��
GZx��IMK�m��6�S��Fϯ(����ͳKy��(a�;�9v!v���ئ}ֶ$u��Hf�0����Vk/�3���緛��k�8�l��z.e��5p�`h׌�S�۫������خ�9��U��FQRnF���_�f�#zg���S3pg�驷�>ف�i+����콗��'f����e���� ���3XͳR�\��W�\b.oD Δ8^M��ǝ��)e.���	{33�e-�6��:N.T��V�����j�ܶ�Ƃ��G5���%Ur��ʹ�b�W�>��^�I��,t{�7U� P��,_���5��O='�l�����.5�U�ӕO����i�QCy�zV�G��J���2Ҟ�˝�katY�1��]N�g.���p9��$RÎYH�	H(���i(FnG56�i�|b�_5�0�B�$0�bJ��X���uz���Oҁ�8vD�X�'��Ό�\�!)^Q�u:,'�(���F��eV��I;8Y�����30r��we@�W\'{�dT�YŃA*{��YT��D��Q�	�ڌ�l;��t�i��^�A�mI�u����3���+�� ��g��z���j�0��Q���tJ3Dė�UG�:%�i���(�DQ���	|�=T%+�
|Ѽ6����|�R �\�S��d��n'�5�(���Κ�|�JB�$^���b u��D�˻��t�O�e[�"HfQ̌Ft�]�,���qmφU?N�M��8ESE�+�����r���zE^vL�Ť0�������U�UJ���^ڬ��nF#�[�pz�p��w2��vV��W>���-g��`[U;yϗ$-�����J��s:�ts1;�(�e�J$~��	^��=�}RE�G�딃���|�`ꌽq�wj�����o3Tqќ%�A��8�T+T7�:Q9Q���_�g�sNM������_oDѤ����
8�l��`���$Ƈ���p֮�z�!���G�)�^ǕZ�QJ�XH7{>�`�����8��w���	w��C	�ej�v�T,=�4��W�H�6:|i���j��c��GY"S�zN{=y8/eƩ���:����1��1���_(��\�lx������zu֮�(@��0#�}�[�cd%#0����#��((��m�i�dG��nyڂ�Y��g<z���A��':�7�V�X��5ݩ�l�9��	HO����^_��tc�yÞ�J�-����V\�g��l:�K˻wR��2M �&�����6�n��\mj3}"��c�,�M۴p��B�)Y*�3�?x���P���4�5�mz{S� ����z�Z�'���/����3Ռl��4J�%ź�q���E�H�zV���0*a�p��Q�.ћr�泝r��L�w�X�M��ĥm���uҰ>�p��+:{Ca�9Gr�L��;�-��"�)�+��^R��s$?I|�U[yc��ko{����s�͋�(W��U;PWܒ6���@���n���z�d�n�SN�������;��غ|܂�Ѝ��h�aMlÇ��0�n��5A��F��g��%�+lDm�ܮy�������n����h��J���5ө��������V\��R̥Q�[&'f��Ci뷎�%Z4���Sk��{�aHpl)���Fw��R:kj׶����~�������;�uX	��#Gkk�@,j��[�O�ov�HP�
�ѴDq����9:(ī��wdY�푽��1/&�>�Ϋ�|�,� �`S�{3��xtu��K��j;y?C9���lU��8�#zS��#�!�<���ܝΥ~����Pu���2�oa�Z����Y�w�2zz<ꊴЊ>b̩�3`�ҭ�fe�B o���U�+]A����ջ[/��TI�P�7eV]��pP��Υ��7��Ws�lp��&n���\�ԑ0+xw���9DYyR�a�����&c_ݹ!oo:H5˦/���g�/�O�?=��jۗ���!��5퐶Z6Zm���7��0��xRz��]���O��H:(Ϻ�k7ú�SK����m�6�������;'����e��H:\�=�)Hا�͡.'cϷ�_��{q�#}m�}���xQ�h<���	�@���k��U璨�)����ʟI�K����b/T�GGu�pԐ���Ivj��*EC�}zt:vzvnI��A��4;���6�J�#g��)�d�<EV>T��U���2 Q���7�����2( �d=��Y�Rd�����ژ��Y�f�k���%�T�̝��V꭯�
ED�)�̾fܭݓq{���z�f��X�jG[��T�%T�G]:�+r_����'o���#����L��r;�%~n\i�L���	���U7q]ݞ�y��;"�ח9����~JY0�t���)ֺb��[���*�%n��+-Q�s��b\��ܙ��
̉�������u+�}�L��Z���t�NM
���p��qq���3��R�R9��/w���n���;Lu���X_3ݳ4dJ�U�9�\hC?Ơ���W�3*D�Zxi)�ir���w��3wK`�����9�Q��t���$A26g�\����6���-_���cƥ�n��S���K�����ކ�����I�"��a-Om"#n��N��b9]�o����TxԌ�m0|��oC��=ҖMv���_�6�]�f�L�7մ`��յ�Ou<v�w�Pn�w����W��ڃ�;j�/�z�i�Xz������n#��i�T[JG��(e������U0NvcY��)�/l�R���,�Q�;�)������&T���_on7(d�L��c�8:#���q�8���s,���F�k�OaltH����f��a�ߢ�9�|s�=�o���ΠρDz�ê�TD��_����cg����[P�{��}W��0�Mɜ6�D5q'����}��a����/�����(ű��6���`�6���a�k1���wQ�-�IN`�l&�``ɀ7� 8@؄�1��#��o��cG�m�!��=m�8!m�  D�m�1�țm�&�l���'�Gm���dq��m�D�m���dCm�;m�Gcm�6�n��hCm�&�l�6�#���� �Ȁ "cm��Ȁ $��Gm���dCm�;l��m��țm�!��m�D6�twm6�#��țm�;l���#��țm�!��m�D	[��ll� �l�G�̞� ��``6 �w�>����?��w�6���?ܟ����������w�������G�PV�����߯����[cm�?q�'���������lm���}��o��?�7���~a�.?�?��~��cclm�����}��o�}�������v�xg�����6�����m�!��q�� p�`�m����l3���lclF�@�d�09� � ����?w����m�ce��g�C�c����������{���~��G���lm������/�?_|���c�~����'����տ�����q���o��������m��6ߞ����~������A�6�����7�ݶ��o��[��h[����c{'o����w�����w罎7�퍍���B~��~����}�������(�o����>�����/�����[�&�Y߿�}����o����O����o�7��ͻ(9������������?���������!��o�����|�r}���~�����7��~����߳cclm����v�[��cclm���ߟ������o�?�1AY&SY	�8��ـpP��3'� bF~��     >�       � @     4 h (   
 �   �  �lՍ�ح��T�mm��aj��V��V�&Z�kbe�1�}�WYlʅ�jm ��LVYw;&�$�TSjV�cj�R[K �f�j���m�C�p�mj�ZɌ�iB�Ehkk�����-HQm+m��!���2��kM-�Fekm�ijA-��I+f��T�mUU�m��mFY	�-m��-�m��m���   0�ѷ�˻T�y��Pބ�ۡ��:r޻�l�v��w��mHzr
v��r���Zn�׳�+�k����7[Wg���=�mΚ�ݯa�m�R�,쭶��µ�SkYJ3QV{�  w^��>��
(P��;��B���>|:(z h�Сo��_�CCB��Э��ܵ�OMm�Ɔ�vw[i�T��Y�ziZu�-�Y�-�;�.M��Wn�����x�ݺ
Ξɒ��m�ݜ�)���   =Р�M�ǽשiTV�U��wq�Zt��z�k�wu�r��{m5B�T�j�S�[�]��Gw�+v����U;J�Ք���ݵm6��:s&u��n�ێW�Ք�6IFٴflU��  ���]�S[]��iOC�[p�N�=ۧV�痯:����oft��2�e�==C����u�s���YT�RwKJW��K׏myF�Kos�(��V�ml�l��klŪ[H�k�  ��Ѡk��t���hI��,�Tj�iT�cU��!m�M��w'J����"и��cn���5U(ҶZN�;`կ�  7<T�^�eB��� 'e�h
����U!3��������t��)r�"�q���Pl�s������MV��ժ�S50�RM��   ;�
P)��9�$U9:���Ө�GwZpU�V���9F�+�:�]���Z�ڀ�m]��-�ƶ�m�T��٥Yk+5�   <  �F} 
��� F� ���  #�8@�  �Y@�w�7 z�޼=�  �/m��jjCm��L�m�U��   x �]������� 
�� �^�g� ;��p  7]\4 7q�4�� ,�  ��Q���abm���fb���  珠 h�{ �=�Y�  w)� eˏ@���L  �ۆ�� ��p@4�  ��y��  E? 2��F�di�M��0�%J@&�S�2jR�=Q�� �0�~jR��� =��(6�  I��L*�� ��=�W�_����a�O�Ϳ�6��V4d�mT�+����מ���<ޒo^�������cm�ߏ/��0l�6���i�`�����o��6m���m�����>���ք?�+t�QE�O�^=�aM��T�j۷7��`�f�;�G��D�ݮ^�.&���@ط�u��vr�gk��aӽ�}{��������U��ý,74�A�E�lM���;�n�6�d�T���Bɩ���d��y- m�xv��A�pg;�<nHn=es<�w�T�U34��j�~�s�{�%��NV�`����l��z��w��͗���E���>3[]���A��:��N�-]��[^�1j7z�>���w9�bѼ�1,�N)��`�e���U-V�]�ѷE�:�4���ai���=;4ݷ��Vh�Ƨ	��lV�����f�si�f%-�ט�qu�J��`�VY��)T04�;$��v����+����x�?��,��*�E�|;O�I�Ƕ��r(�6���?��\�q�bo�8p��>��p!�8�M��:���񮃭a�/s�%u�t9V�v.�{��.�]Ԥ�L�I�g-N��"�ޠ��Gr��ݒ��^�<�Q�����+{m��7�k
&^͙�of���up��#w9^Q�,�F���$L��<[�5�%��Ix'^��̕W�,������d�!0��(x�ԔI���껯O��L�#�w��Ԝsr���~ck1�t�3vm2�J�-���^�j�A�Φ��޷n�2����8�{�y��ʲb��u�Wl�DɃ4<� z�3�KÜ��wl�f>�����A�LLU���VK:\ #I�� x��A���i�Ԓ���/��Z[�4�<��&�Mj_,�N�dO4u�43^k��gb����]���&�}V�&&� ���W~������{��x4'A���;����i�Xl��;��"��T-�FnC��O�����8zu&�17�Zaqv���E�I�Bz5`��k9���C��8m�k���c\�鷟d%3���N�#՝�Eʌ�v�^�aV��'91����9�H���U����1M���L=�������R���J�Dǎ����QhMA;5=�`�`l�y�F%]X�'1r��s;*�<鮅�w^�I0�������87��;4-#������e���^H�.�L=(qn���UCy�Q ����t��d�C�Pw{}n�&fד�F�c�̬�ag7���vu�8�	(�CT�k�V�{:朙�Ƕ	w�lܜ�����D�:\�h��J�dȵs@��'�y�3�b�x`���{��{�n1{9	����Q�,n�磱���M�rhg)����$8ɕ�uӑ��;�"��\͹u��ϳw�����ے۱�����;�ge�#���+�!؞���hX�*��-�rRٻ��x�ѻr**p4wG�m/�`OBc+r�f�N/�z�VM*���P�Z 
��,f����ϥ�G�B5�l�-W�g�c������;2�飮ӽ۫�b]� ���k�.v���;flk�x��݈#�N͒%�(x�P؄}��y�ً��K�
u�5���oBs�-�y��b᳉\;�ap1�:��[Ӡp�Y+`�r����Hc�ݘ�КȄ@����򥚔%����^�t�,�9Y�"C��s(�$�5Ãt-׏tU��v�5�2kʱ^���i�J��yɜ׫n�%-K�!v;���՝^0�`:(ys`�8�Ha͢�F����H��!�	�K�t��Q'���%�����"8�(���5d�/;Sߩ�;�v|��qvz��Iѫ/���䛨�Kؖ�-���ӂ1���i�&)+���2KdK5�u̽۝Ɂ�o\�9cӶ����s���c�q���s�!��x���A�s�d���=�^���7]ӻ]���BЮp�i/Qt������3#��3}%١v��XzI��jAk�X� &��t�K�,����.�ߧumn�A���Z���{�0���ƾi^�q�(JVg[��&�<���I*ܛ�9�}��oR�
ٺm�ۜ[C#ŝ;��v�{C!�B	����gik�h՛ݧHټ��\4�F�c(xVƐJ�oE�8�r}�}ĭ���	�,¹�=ՙ5i�� �b��97N�x+�ro8.@�47�͖��z��+��k��ל�z,Ӽx����ע�8R�EU�����1c�č�ܴ��9�&i9�=y6�35a*,��';������x���֞Z�;/E�j�ǫ;�w
�ݖ;xU��;�0L����;��v�lz�<�/܄R��V�+�|6k�f����Sðgi�\�8��kgs=^�J��;���|�kR��d�9SЌ��7�tp=�q�����H��"�U�+����6�t��v�n��ͭ�����^/�n�Gu�iY�0�E��8;��z�b�n�{�� 2��xu�.��}������w�ZnK{pi�4��^gn���|qvU�h��ǋ���ox��T}��%٫*�9�������/j�~��%��y�zv��
�aXgxMy��g^(6�q	}YV������	I��F�ɝ���$�5��[D�n��Z�	�s�[ij�F��n���m���N�:^�y�\�Ǽ���ζԯq;i�Q'e�Mg`��GT������k':|ts#؞StrLp���Iݫn�w�+�B#�� �Xc:
U��=n�����d���,�����}�m���w8^L�\q�Z+�����%f!r	e%��c�_g����ʶ��I�w��Y��۹�bc_>�ӓ���j��.��t(���cr^��G�A�H.v	kGx���L]&�wYtZ����w{@��0�i]{��ǒt�%��`@W
B'�D��6�Ǻ������ф�A�������`�FA��Ò�f�,��%b��������wN,���������e��{�����dX���#ڣ}�q�1���M�	0� �C�n�
�5��3'+���#j�e��Nj�n֋Ś4F��q*oo�7"|�P�5b{��)\�?��E�U��{NQ��9��v�7��"`a���{gX��d��:w�������{�-�� c�o��r�v���.����e�7%�oT�{�˪ʛ�*	��[�)[OJ��e��9�ʠ��iͻ�>��M�w��[��da��o^�sN���<B�8�Es�h�<�j�W-�BK�^u i�Lh�I[���k��X�{ĉ���N.������D�ᜯZ�+�:���C*�C�l�f�Y�E�gL'����H�^jo���FZc�CT���&��:��ueJcZT�=K�T�R�yoGz�y���^Owx�y(�O7�u��4�ۓ�<�����-ζ8�8tD�q1�p7˓�X[��zl!<�f!g�3�����{��<��ɫ�S�#S��Z�k�j�:ΊV�0���/��ƦD�a�MG�9j�"��'Wy���n-���e}��p���p/���Ls���ˮe�nʰ�X/�2z=Ou���r��rM7p�st��\�́D!C.�E��U�a��17Q�DhO�vG,:��j�P8�;��z�b�������1}ˍO�@�MqG+������E�P5��js��$w��⻆�b��ʒ��݃r�mS6v�f�݌j	����obX1f�<��!�r��.���5W�\��Yq�j <�DX%��F>�2�X�dN)�SdeIM`��ٶ���ڴ'�U����:�����ΎEЋ�g^��NX�:[jj��)�M��>?�o��zx�L\�������p�No �EXj���|�����*ᩬ�����	ޯG0vv	�J�Gl�����^0��-]���vtG����h\x�YՁ���G1r��㻐�S9���_*f����*��*�p�:40��};.O� ��
g;�;A�tX��`vl�M�;q��V�i�T�Y��vC�Z��
ana��h6d�/z�FS܍.@%9�+�w�)<�"Ý*�ާ�Lb�R�Њ{L�d�V8�v�8��6�k�V�}�do=��S#��ط�.��v��So5�U�q�U���E�/RZ�V�;���n7�s�$9; c�vŖ�|w�����!�2O�@�'2h��3���n]�tx쏲�k8���U��	� �3tD��E�NwɴR���!ÐX
�6�81�{i���*sb-̊������&Q��l#��R{��ȰM����t�i�1�$�+L�۸�����k�|jx�㓝Z�c�rdp�ٹ3��K��e鸗��c��֣�����5��j<q'�4<]@�q3�{iȓ�Ŗ�͛���$����7Q*�ݒ��ݨ�c���M��&I{J�P�Ђ�2,�j���t��O4��������F�n�/��Ly�oɊ;6Gk�I�'i�/s�K[��߷���I[z���v�ӛ�3��`�b-d$��u[��b�Z^ռծ0�m+i6ׂ<j��w�uv��Sx�K�j���J`�Ķ�@]�����q|����l�pb�Ɋh��܃���:���C�E���m�Eۥv��,�9�8�d�5��68]�5�L�aӲ�!9ю@�:E3N
1)N\1h��uE��f<sm{�3�Qs| gK�8���*A��rn�7\[��o9��+��]�	+���.U��p�+����b�f�%�w�ݶa*��s�F�p���c����kȆ�p!�)��6�~c2s�g>چ澸��>헞8����9pE\	�`�*�᝱.G��v���-��]��� �2��e$��Ux��~��^�f{��R$ �s2��v���%�eȦ�2��A�YQh��}"����^�+;���p�9�nn%ݑk����oQj����Ź`f�(�4�-E�k�x��Y-}���t}�����u�ܗ:�'FT���Ǉ:4{��&F�EθK�$1����+��7�hC7;Kz��4���gV�ޘ3{�|�it���*a�m���R�f>�s÷w��8�c����P�m.��{/מD m�1�LV��-m�;�����H����휖傉5f��]{�Id�^D4�n�}˚J��.�����p̨]���Nٚ;x]:._����o�n�ŎD�
�����K��:^8x��Q�T��]�a�n�2�ۖ"�e4��;�h����*���\`���q�=!���\=�v�I4k�a܅�V�21�-ƺ�<��ӻ;���2˪E2@y����Ӯˉ.�C�s�d�������t�a>ܺ� �Ӽ¢��ݚscܚ4C�wl��x�x2׹�^%��[�a���gr${s[Mh�8�4�ce�=�)�{qt90��}����c�I�ZQ15@qw\v��Y�ZF� +m9���No�}�͉�+����v-wL<��q��vp9XR��w)���(gn9�E#�+��@,����Gd�x�j�9f=X2�%��Dr��Ё]#�'`�����Qq`v��!Fs�,�|�:j�{B�5�s�۝�_����g����Y8��Łd'+ve�n[�~O�᣺�������]��^�a���)r�{M�Op����C�[������r��5�Wy\X�qp�Z� ���j�Z������a;t�GO�C*.j�>�vt�!-נŇ�����9��4��\mΫӋ� r�q\!Y�w;V�WoC4oM�,��`��o}�g�^��VrK]9�`Ĩ�[�س�#j(��*)5Ⓡ��Ƣy����a��;5�Ʈhn<�p�w�!��VXΙ8Lcr���h<���5w�f�ֻL  ��2NE-�f���58cL�;��:�����7*�BG��S4��O�v�ݸ�Rz��D�'8��M���qvt,�����dx���� ���4&W���1��t���x�^3�W#w+Ѧ���Lj�e��r�)�o����uL�=����kq�-��
{r�(leq�q��yװ��`��{�롌Q�t�F��V���5�;o@���s(���{m7"׳g�V��Wܱ��L����y���\�^���� Y�{[�Y��l%���-+wN��0'�wK����v���Q/Y�
�m���I�b���"O�[c8�Ѿ7��=2n9�.�ILj���,�?i��Gm���]xt���\|��p\�SI�a��:	%i��}�������7��{��:(Z�g�q��b�sPR�S���f���݆�d�5�]7o�idg3]ʵ3�^:m��u X�<c9�	��hi�@�9�5�3Pp��ex8��Zػ��[�8�����̏f�������a�r�X�U��-�Yѷfn�Wv��r��_YųA��v�W;Yn�TE��7"4�;]M;z]�uph<�xB����{Y����\�y�A'�Ɓrv��:�N끲�D˛K�Mί5c.r�0�o������D5��Uן(�����.�69�>���p'�+��P��ѫ)�cl���ExkY��'�ӿg] �y���̊�,�CD��v��!���G�E6��\,V��K��]�awC�XN̓q�#�q�QN�s{!d��,�����8�^�'���4��g<�ҩ�K�����J�F������=b94%Iv�nq��$��W����s��箶!�zJue-�}��Х�l��\�W���'\j�"�u�X�#��X����^�yug=՛�Y��Bp��g|+y2�W]`���8�pzsޛ�P�M�3���9Ab��׉ѱ�6c-��91��9*��R��[�M�6�dԁ\��谧E
3�^��Toeo��K�c��s��U#!�n�V��L��^Z��ndn����S3�g��L[bG}ۅ@���=z,"\x�a�{�뎓��}�T.�DŊ��&.;�)�ޕ�F-59Oy_;m�tӭ7�`s,&�� ����
�lژ 4Q	J�ܗ�1&��[S��@Z��CD*	n����^ѭxk/cH������X�'bu�;i�6͸�./2�P�0s�Q�ڰ�M�<��ls�"|3rm�=�5'Ip	�׉I������hCkw7���ץ�@�N�g���ڤc�X�y�յ����-,w5���d�n@��;	 �p��c��6f�]�qg���yF�+��p��5q��0�n����׻���n館�V�U��%�f�Q��s;��8i�4�w�44{��٧���+[83b5���B(e+ �'|�X�v�}�2�]%x	��$��e�Z��Ɯ��G+O!>Zd�݄ u[&�̃�)�l�]�|�M��oLW�p���ߞ,ۓ���1���<��b��u��n��;���Gn�4�c�8f���X�:��`���2s[��T棘i:v�U�M#�kR9�i����x35�fJ{�nQ��-�)��Ԅ�We�a���ܘ֚��Hy�V�O_u-���\��E�,��捥�����R�P�qf�i���(�^�X��$����1{8h�Nv����p۬tu���L+�I�tmd���f���[ 1��.����zx��c(^7�.�؄��M^zN��Rʉs�jġ�S���hs���n)���c����z��\��
�Y�V�%\��NaZ�^� �� �܍P�E�0�b���p��c+��Ds�dwn���ܮ8����[[]�C���Qݪ2j��W-�z^�ǝJ=m8��m��v3f=�oWt���A�=�[泰1�g7qYu�Q���JVÉ�G;��i�������*zU��gk�=ڧ�G��$���gswN��pa��gXb��k�c<�I9��/�vu侃l�z`�po<����|y�?5|[��9�^�|ҽK
=tݢ̋r�n�X7!f�[[-Ė}�)�t�gd,��	w�6xd}�G�By�c�c-�9�V_�u�xg<�w�6�C��(N���lX�E[�v�cY.;"�F�C# ������P�;vgt��UA�wb o/:L��z�z�m�Mc�K��ܽ����O��8S}"�T�^E�L�ϧ���5��k�7$���V��#Yz�n����[��!Y�5#���7ۂ�cm�̇uiG�;6����:�;�e�v D����<�2<9��V�d AI&/Ql��/�-&�x�R���e����М ���rewmѢ�W���+|�9�{�f�݊��f����f:T)}���]Y��z-s�ں�`��qr�P����7z��j�����{�vv��'ȏ8�Uh��� �0�I*O�Y#)�ˆ<�G�o�r�1�փÚ��J�L*,�s�_>-�I�m]
O~/Gl]��`ݾ�9qQ"v�Z%TvkRPm��ROO��7xh��%Yo0'�bZ����
Ҽ�Z� 1u3�;�a�d���r��ق��XN�FX��0���ĉ����;�pE�@#�^��t��u�΄(�n��##�_r+1�yA��+ޖ�r/��)�)�T eq]k�3j)�n__:�W�y+E�MX��}pM����0QVM�\�/Qi�ړ�gy���h���Vy7�,|,�c�i5͔4�S��΍�+���Q[J	�zK��b�\�nO@��y���%B�4]����h���@ ��-wm�����{Tv/>�E�qf\�����ȶ�"-z=Fr�F&6�g�>����*��n�3s�/w�����������-B�gȋ(H|��k���+v,ة��q��50+��/l�=݃��m}|{Ɋ��О�+.O�܊��i�"�e��ޜ���Tw�oy@En�)o]aͦ�fc�Lj�j�%�v�Ġ�c9iH)�#���޻�����z�B62���>>@����6�����T�6���h���R� �*�m+�W����[a�*T�[䌆�^��n+r����'MDu�\c�!E'�{�kw�w=���T�{���y]l�jrZ�54���t���dKV�>j��6���d�J%�J���*%��1-�y�j*U�9T��\�m��Kb�N%e<�V3���ɮq�_�ȖD�w7�.y���j�|�U��z��;hs�#۽[qZ��Qж�^>����S��0�[����M��P{���כYV,�M^��EHM��Y�-Gbf٦���}ޙt�ꋧK����fU�G��D�3p�qR-}A�:�ʥf�!5����h���!e��Լ�*�ÔoK�j@�B0�C���Kιh��ԗ9n[�)�[u��ȸ3�ҳ���Cs}�L\W�k�����ʿ]0���7&�����cLS��`m�.>�{`��ZU��� �S�H�%�oHx���ʭ��x�(J��ķ���#��p��:�J�|/�&X�:���5�w��I�t�&��3g(�W����R�W�&8+nCXGs͘�u�uiW
:M��-;wl�Lt�8�:�]{zʺk���h�����"�@�'Ms����B7P���Ţ���6��@EE�O�I�Ω�����%��_nz���74we^�A����d�N��j���.͙��BD&G�+*D&�����(y���.�Aq��a��ވa���p��nnp�h�D߶�Zdˬ;�-"ߌ�[MZ��f�5%��MF_<*�X^��hٵ�����2���u�ȪJ�|���	�u�k�m����֚����Y�I��Nh����p�h���������p>\FCF�>��¥I�n�w�*Q�AV�Q�I�W-�x�-�ene���h]x'S���Ov�:�o0ei#ZB��U�=��St��}��sZr�����&2��[J������v9�<�����^ng+y�%f�r����Uw���Eѷ�hm���4.l�@���f��/�ݪf���!J/?/.��#U@ (�_Q������^��O����v�jXi�=Ej��5j���v��P-�EJϟ`��mA�̚<+��铻Y��\ٱ"py�޾���)Pf��YR�9�c���U����`X�V$�1�����@{�9�j#}&zC�S�������y�3��*~�}�za��$�C��
��[;R�^90v/yQ���p��H��M�ȚC9�ah�Mu�c̃�N�����`M�Cz�ň��mˠ4�OP{s_R��mJ����g9-7��7�9[�)��@����*|@{|���i��ռ@�j�,ڹY(���!M0;��o2���/2A��;���Lk�yۙ��̤/���z�-/��7:!5��xt:�7$Gy�J�2j�۠0�Ґ�o��/�9E���\ �ɗ丩���n=Io(,f-��3�vk XuR���z��4�k�.�j���/
�����J�&�ΝO��9����j�U�4zh���U�E�;�J���*�\�-�a�Ӣ��Z���`�s�;Gp�z�')R	k�x��%*{[��^6��R��"+h���y���P��6��[����[�|�ݻ-���5��;�j��nE&�M�W�0	z�qSxӶ{d��v�[���d�t�͔9Вqb���2Bd�|{8���j�AΌ;���31�X+I�)C�Y�i�M#����AFS�6����v�˾�|�m�tM]v��2��|�#�i쀢y�a�v짹|��?t�����_}��q�cܺ4����i�T���b�w�>��m3;K3F�կ4F��:.��-���& ���s*wR�SÙN�/�r�������a��t��fit����L��@7R�J�9B���+�x�6#R�U�/a�;4�:�\kI��Z$N��o��������GC[�*�W69�ܞ~V�]�"���<�t�9�
����7�Wͯ�]h���Yt��b�[gTMt�봪O��2K���E�&�%؛м�Q�$�+m�=6�(ol���.��5[��pRm��B�6�&����.ȉ�[

���;Du���B�q�Z�!��j�m���۸������u΀�r��N�Y������wk�X�g��0�)˫�J��Aro���pvѾoSh��Z]�y�Ѝq���Z�5`�����ǷPu�{fޜ5ġy|�s}��Q��M�YF��Z�:v�A���#�Y��ܵt�䄀N��\Z�+��
ax�H��;,�# Z΋�s��,Lsͤ���������|+'q��y�]]v��S�#=���B�u+�6�V��twy,�t�y�d�.�R��!�R/�B��\�B\�V�����synuIGc���I,D�s�S4��,���c=:t�#%�$̬ga)���^}�XbD���jMF���G�臗�^�(]ܫpW/U��_U~�u��'�_-,����Q��4*ػ`yJWH�fTw.�g,:��r��B麊�J�ʛ�-=uSr*��q�s�:�7�%�,(������s�N._kAZiP��k:YY�'!a�]}���n��t�458��B���ۧ�A���>8�T�6��>T�%v
��;�����O����!�b�.���wΰ賴**}����P���N��W���;8��i��W��w���U���j/��9��ol�{]�8�k����4m�J���"�ʝ�MmLu�*Xr�b��'Y��8�m-T-�P�����fY���(��$1�/��bW��r������_!$Y�����g�7]\EX���"�u�șxs}�)��ż���GF�WB�������%q�64�*��Yl��)U�y�#�	��$�}݆�����w8\�kA��d�zsd����	�&Sځ����#���&d��>����A@�mR'�tY��7{G��-�+e˥{[ǁ.���df�E�R%��Llʕ��*�D�K�h��473TF&��/qk��I�jVaV�E�}�U��5�pQ��@0����9�&�.�WwL���Z�����覆H�f)���F�}G-١�Oo)��v���+�0�'s�;�-����W�2=V�M4�D�6��t�D�+�X�%ƒ��ƣ���gte�l�	V��Wn�9��OSgueM�gm�F�o����yd�}{��THOr��y�}a]�������%���Տ)���E�����ۺ��7�,�����gl��د1�7��Y�+��C"=z�N�<�» (0��J�í	MX�ˊ��\������ji���%Z:�������Ң�x����U[r�����t�+���m#n��<�!G]u�t��˛� #�e�G/��#Kav2&�C��֜�닶�ݵ��U��J���>��y��[ ��K\�yeR�la�-1zn�ξ�l��;���Dg��uJ�f�6�e��p
�t��-�;�j�l�ZѺ�]��3�A�;N��X}O��E��6g���J�K���	I
L�`�D�h��}�r�6�۹�d��[T���v�5�ƪ�<��xW ����w>h���qR�l�|1`�t�C�0���b:V[�e�=���vUoo6��j�i[3�vK�&�#��ɼ�ll��й�`��M[�DG�}���-��Ӣ�'^�T�x90���u(��~��j�я2$�Z��F�/�M�|���m	�i�ל/�r�v=�P*g^�t�Of>�X�%Ķ�3uϛ��d�����x�őÁ��Nw<��<˪�g^|&V����qn��Ih�n�h�s�eqV6�>����ͧ.n4D�|ŵ�x���B+4����	��w�j���JgX�61����&�~�ٳRŧ��ˮ��|���/f&�k�R��M��	n#.��&+��,p��
��� �K��i�:��K*2�H�*�dR)������>����M5EjgQ�6���.��{p�R�a�f7Z�ϲr�zJQ�ww�ޱ&����u!|�x���BY[.�ENV󣹛Y��}�PWQ�CE��Y'���p�[�V�UdZ�űnĄ�:�Oo:�!.aڲ��N�n��v�;���B�ECh�˓vb���U�G���ܒ��y�q6}��\����jo�-��lbL�At��.[G\��/+�i-xЮ��c�{Q��y���&�j�i����[�X����4T��[���j�l�S	��eh����x�E�j�C�����G�FWQEJ�x��]�N9  �J�R�[vi���܏��#�l���|-�Goy�;S�Ev�Nvw�!|���:���A�)<:�q��f)�F�:��f�Yw#���z��X�H`[b��ɮ��Ѯw�p�%�}:�j{���c��(�Y^Ŵ/cT?�2�u6mA��
�#o�Z{�6GV�t�xmt;R� Ie����n�d�j�
���k;�*�ҎΤw�T�n�CR�6�8���[J����1��r������d�Ӗ2Lݑ.�rʴGoY�D����];�=��H�5�F���=�3�W ��Zz�V��j��N��&2;j�́S���ή���s^	��rI����^=��w�ǃOG��㲕=�Z���\�x)\�}P%��	��O�}|��M��m���0l�{���{�����m#8)�5�	�������9���y�����|�{d�r��Z��I���=4wI�k��P���{�vBV��G,F�H�g+5��X۩���V���1��pK�DG��@M��9>֓;[-�Q�/��fE�(Ĭ)c�\(�ŉ��Q�q��	�"��K1#��y�C��Bc���Pu&#�ɬSٝ�r�����	5�����o���4a��>J��"� M���t��wCtK��mM��SS���_r�gr�5��B:j����Mjj̭�&b�h�9�]�&�:/z7���"�$�Hu�!٢,eޚ�ݚB�&.��9Va��T�ُ}X|7K�8ꦬՇ�D9���SY�bM�18��+t����@ۺ$�nu�5H�WV���q�:�	��(h���C���]��rGo88::�v����Xn�r��J�ӗu���ݰ�L�����Z�)q"��L޻�ʴ#������d셵�UL�`e���ⲝ�[BAr�y���訙}�F���;@��܏VR��}�.S�U淼{�h��,"��f�4�B����r	_<���Kerbc���k��Ы����Ar�4�l�]�y�3���{K'?���OE��J ��)X�]Ի�i�E��R�B]����b���ɮ��gn�9eҨǯ��¼yo�o(닧1s�o�:��K�2h�=7L���]@/v�{R��4WEn�^�<�Y�+ٵ�M�i�wBWy�=��+����:w���z8���7�O��ל?�p7��S�dx��*=��M��d+,����`�2�;�:X����3�f*3���d��C-�]������ǲcIlZ�5yD.��4|bFq$a�@U��,��:�T����\���S��s�ٻZ���Q����1��;�r����`��+{ ��6q��m�d�p^b��2S�1PO�G��+0�ح�C)�K'Ӳi��i��`Ui�%w�fCcm�g�V�w�m�X��载R!���7�ֱ� !��\xt��*��"�v+�����)W؀=vL���^�o�=��6��
KxQ��3.e�qϔQ��a4N�ͩX5�O:=�JN��S��s���q��c��Kuv��Y6�R��V���4eKƇ>�n[�j�U�+Wy?O�bB�n������i�� @֩5��|6]��y�|���6uoN�?35,݌jz{�p�/��Q��Z9@�b����ys<E|����2��ڢ��4δj[}ZӷcgFR]EП�-1�v`7��:��n��wX�X���Z[���{:e�k����..����P����L�j��8=7�ّyJ7l�y��t��<��$�Ӂ�������g';�B����l�����>iH�]E�0z[*�I��vv��u�o��bq�o��0W:|����ff��E>�ՊT�=��\��S��vÑ��������Vl��)�9��UUw��'�H��*a��*`$yؕ��:��%�l�A�pě���8���$��B�c��m��W��q#��펻B��WP:�� �G���fl��^�D�սHn79���҂ձ��%�0�2����5ye����B]�g���I��޾��R����8�0�c]�}9E��f���nlf�͍�*HU������Oz�f>�0�PC�.)����vK�q�����N��/2T�EK��.��t����q�9-7s�<�͔F7{��]n�I�aWqP�ճ��E�!i�u�6R�E$�X�Q(3)�P!�oTX��M����"�}Z3qMwz��h(D�G�]G7�=�cJ���e�0�����gc�X�F�e�]�j���.N�@js>ޱ������T)�� ј��Y*��u�
���g?n=8��<t���� �~�0�K7b֧XT1�fHI}�pQ�nԝ�xN�JSag�uh�ϊtL|�|m��fK7T�b}���a���z�b��4k�/���X���|Ұ�Mr�s�n50����ҘLPu��Z|$� �g�������9:��*Y��V�^�E�2�����C*Z�� ��ې�<��H�`�1Q	�@9Jⴙ���ܟ{=��{z\h�=>-��gzz!���<�9�0UG���P'\����Qvh�~"�[y��Q�܍(��sz��7�IGG�@�2Af��xÔA��d3�؉�Q�vU���<��-9�s����=�$C�yv=AE���J�޺�]��^,X/��{�=��ކm]����pgAh<P�\�C��`n�$���3ܥ�)Ggvҥ�a=���챏��������g���9=�G��l��kN��YMMq9+E�Mq/��k�'�Q���(trO�ί��4l8eX�^��|ƍ��W�[��z$-N��"�=��+ц����v��H�e� Q��n��oD�K��hs�����~}�7��5�������/3V\�n����*Rh:�Z	X\F���P)���፵�ұS���hfidꭡJ�D_�Nټ����۽cN6s�sa��� �w�Cu�#�w��.Ca�2��C�����,�Ծ�.V�an��lW heu��~�1� ������ј�+rWU�Mu*�]ݤ���*@&����sź�o5��Sy�&XGy��t����-����%�E����㒅��"n��X���>�%7ݞڀ�����+��,������t�o��n^C�z�c{�i�zI��?Lc^ɼ��
-�}��]�,K�Y�@\��f�Cݓ�2u���d'7�����%``����5:��/��c���P��;�/~]F�f�b?1�E����J��A��9�q �Sz'	��d�T+�z�d�^į�F�qY��Ǻu��ZF�S��w �X�d��P��^�=%#(a7�������ћ�v�}����K��9t���6���sֻ�.O���)��4=�3�{i�-�y9�D/4���|�)0>�_7���$r����mk��w�}��8�2C��f��'���hk��ԱNT���m�\]�f��؇D��V�T��_^�|L%N�E�X���X!�Z���s���F���7rm8�tk�p�2�߱S��0��� :w+]kC��#���G7E�V/��ɪ���󰓐Ȕ�a/�jW�Զq4 �	�U<���CP�_?62�s3ä� ϶��"R�ң�o�}���b��p�,żCZ�cɮ���0���Nȇ^�Gi��4�-�-l�Cz�Q3v+��1��!�yv�p�nb�ķ&�ޗ;��ez��#�K�����	�#�����x��('�8�>_v��v6��Dkz�s:$��i�
^-˥���m�6�.
���{�����jzS&f�{"�wR�]]�&��_cy��>5�(�3� �ЌB[���*���Tbl��SS�d��(��E�r&�<�e����lwt����~�ʷ�Ĥ�5���j����c�[۳E.��hs�w�s+��G'����e�>v�Ȳ�p�fC\sd��F�Xh��v�N���L���紬�G
��][���&?V0��n%,c�xS���Yk�"��i���r��3K�s8v{J�Cy3�����Z���S�l���YfO<��J:.��/z�����X�;�@�%h
�$�4:��a�:�5����,�lm�ٵ���3L��%8_�љ2%�%2`�k~;��#��U���M��j�nL�g &�U�_}ɯuv�w}�_&���s"{B�l-MC�>/Zi�r�%ۀˁۛX�:�9/���k��7'cv�r�L	�u2�LU�E��M�Ţ� 8�U�& �;}f��L-3�Un�ʆU�/��䖌�L90]�"�HOR*r�`����;��j�6�\=T6�9^�k���7���5{)�"�K7��FzOL2��/`�qn��W�Շ�&��$�X��9�4����T{�93~�������M����pd����}�Fo��捫o(-Q3�6�*�fl�����gu��y�	i�Y�]�e ɕ2Rt-Kt�'�0ٷ�X��ܻ.x�k8�j�:��7�Ӯ��FհH�6�p����O3��7�s��q�v�_7r>�[3F��[���y'�,��Q�����q^�{��7x�lĻf<�����C}Έ��ѕ)9J���0���ۆT�Nr���ӽ6��f.�
�A�5�E6�7/)˻�ma��v@P��Gv�oM�v����eJ�:��TUv�۷������>?c�
�$]��P�^�VI��ϻs� -�\��f���������b�u�����7�<6�g�t�[���+Z�ḛt�W����|�o��$�7��7S�ei�ܮM����jnv�En�g�2��ĻV���Xc�s�Z�c�A�) ��wQ�k'6uǸQˁ(�
Ȩ3xm�\1ŕ�3ni��H�a�1�oU$g�U�RYq��m�?��9����bu�S�=��5k��}�S�^���ܠ�ц�a��;q�:矷`]�a{�ʋf��\)���Y�vvZ%.�u���AV����[yK��f��[�6g��ط�~��_
��(��5<]3܂�� �sJ��{�y�zC!кK=YQ�t3���<���Q�@�ӵu+x��r�)0.:
��Lu`8Dʷ��z��N־֑q]�|^,J-	[�W�eC���}[L}>�{��q��Z���$@�&"����Q���0�1��@��}��yώ3���Y��ĵ}�)�&�$�(�����@B5v� ���v� �^Sꨤ�u�QW7:bِ ���]y�ú�ۋA]t�ȳr!9�ޒ��/#�/{L,�k*S�]oucg:�,�6�m���t�P�_I���a<<҄s���+���/`�)�Q�c^Ȁ��Z��pw�w	igd��r��mI/h��'8|΁q��m���*�w�ӏץ�/<Ã��M3�n��Aבd{����4���7~U�w2��y�7����)"�l�4),�՜�vq�%�m0��\:ڋ����s�5��C0$��)���F��b�{�`���bMT�z�UA���N�9]޼qN龔8Q��&.ɋJ�Pwj�_ishw9�����ޛ=����"�Q��J�=7xk������7pl�Yp�Kn-ʈ���9�ܭ�bCR^VV���j����ԭ�uǫhÊ-��d#8�O뺗|u���M$Ԫ�Jެl�L[���_�*^�F��`�Ԇmt�+��ò�+�bx�w�
���ƌ�������f�3���r��@'F��_g �i�{b��u}�����W]B���ԓ���AǦ<�)m��+���#�@�Ԯ�ΧX�mZ�����'J��iZ��®U�@�v��Sѝ�y�V�¹�A#��'U��4~O�¸L�NJΞ�v�l�"9�ov�ZX���tϟG*:F^ͷzc^m�ﱦoB�*�}��������w���惔7(���D�c�����@��Jx��{7i�,�\�*�r6ٓ�R�0�ʽ	ʋ8^�u��%���f=��ڻ[}NY��R'��m��V<���b��$��D;[���˝	�� a���+w�Vf�r�8u��hїώ41���9�m����;'J��ݳ�Y�G�j؎ƫ����ܠ��c.���l�:�4椙β������L;�����eC��k1�5<�_!T\�7}��h<[����w��f�T0Mu1�3���2#����K��l�T�A 0Q�(\^�(��D���z���Q�.Y��XNP���o q��]|��^�8�����H=�� ��;��Kjw:a�b�
���w�0�U��[6�;D����ٳ	B��x;��ޏwE�Ϙ��۹��������0< ��%�g��U�By���6E��Sdh�VC��p�:��0��]��tM"���I#f�WW��Z�&u(�p��f1î�45����n�f%wƝm
�#y���M����E��ZE�οp�,\�\�Go��w𭛙���X�)4�#�Ǔ�1�t���/)�_[(r�׆&¨,�ܜv#�]���@�]⸣�rQ���h���^osЮV�G�&`���H��[3 V0�䶝��oJ׫jk{��7�}+$��,������X����좿��	�)��s�1X�xr�KQkz)�:yn����#ׄs���+$`���Bh7�v�34-�[��1i�Z�|�]Y)�Ԇ�fՂoVM�]�I�!�]ы�mGp��^u�YF,�;�n��JZ�N�ũU'h	Qu�ǲ��1R\:���d��k[4d�2��2nc���X���
�tn�t�c-��r�ٵ�姂�a�w�U
��җ�5�W�r��OB��k)�̓K�F��P����&��e�o>=�^"7�)IO��w�c�ks/��"�X��b�K�����HUN��L55�J�����}�EKL?��X���)��z�SF��f�HKה�����{��2u��-�����ĉJ0k�}S��v�����ܺ������F�ĺ���`��}ޯ(y}�h]�0�=��pm|m`����X�9S�����20PV�2��f�<��(��z�#
������c��w<F��7��o'�˗�s�Z�\�l����Z�/ͥ}ң��/��s(�[δ2jMmM��o3/U)�;u&mpX���\&zea�R�j*G	Ck6<-k�W�����X��x����YMߏU�s�OEb:4�KAAΘ;u$�����ʬ�q|����꯫�Ͼ�h��z�����5ǎH��d��ZduL��*כM��a�a��J����%㘋�8��Ҝ3vr|z��N�n_7�Q�%2z�#��e&ɕ�:mbH���5�,U�&ŧ5��ܶ�[��%]���C)��}Ù�����5vrq�`2;3��T�[�?)���K���F�a�nM�;���1�T���9���&x�>Z|5���/���mܔ1�kԽ�C6UL4��q=���V��8M�x,�4�rr�	�fkz�{4bs0v.퍝�����h�"�C�q�[��y?OtS�G�;��^y�,E��y$�:��k49��&���c���gx/�|�t��m���3����9o��)��2E֢������$�9�֞���;�
ޫ���E�_}�`�<�7�b�w�T������Y���uI����˅���`�7Wa<*�MY8��tܒX��+t��T,�u�y��x�*d���rcbc:�,oa����;�F��4z�{��	]�Bp̏���Kц%k��bˏ^p�7%�!&]Dm!jp�hwl�u�;9f�ج�1@&�s��-o+�n��c�����+ct�e�zûxlT�[��dN��|؍�eU�]�Yٞ���ɢ^��h�X�R�a�;�8�����#�Q�[��6'�V $���扮�o*���e���s5�(m�6S�V�͉iK��3/&KɄ K#�%r:�9�)����TNg�9�y��3c��T�u��rg��Z���TEDU��n��s��)8��u(��ܜ�쪨��A�=�/q�]���
V��0�u�ʬ8�%.ah��m9��[�yb
�QT7q&�T:Y��(�AU�
�9.�9VBu5���n�54��J�� ����좈;�^�w7E��rԹT9%DU��w]�rIXEաN���9̄*��«����A�:r%ZIۮ�a4�	��*=��\":�Ԉ���M�I�=L����U��9L�vZ�N��z*\�LԳR"�SUBB��%iY�:����QH���$�s�$*�B��*�DE¼��ww	�����J�EAr��eI�r�΅r���TAs�"���矞�>jI�Y��o"K��.���Z]%_J�Q^_chʹ�=�F��H�§Py3t�F�#nVŧ
�p��oW�s$�	�B������yY�� ���1:���O�e��'4,@w=�85���{�i^ɛ-����Od���8�u���|�>��kx�V�:A�?`���H��+��/,�c�~���1,�PW��ڃ����+o��xe��\̬��<�5�4���N4(���_��vX�n�Gf�pV��ߑ���4�m\��n4]./��\��X�ܖ���x����{L֭��P�\D��w"��ռb��N���3[�P.�I�����׽�tPq+K��L� 1�01i�fGE$��q.�=�Kf��Z�j��Jk��֣�����0���Ϫ��2Y_XD�3�-Oc,���1�"�O7=��b�6j��D�^����k�Y��>��rΈ @Y��}�C=�pl��	�9�-����e۝f�+�,��]/��t�\&b�:69e4���dP3���ԥ�vF�9t�1��f0坷�=����:��}��jy܌����;
�ܮ==�ڤ#M�J0��䖨��ó��݁�4�wu
۳m6�3w��mWԁ�r��ۺ�=�VE@���w���0֖�F{��@�I���	�[��m�����Q�*1꽫ђ�}!�n;���f�Mͳ	K��fi��i729�;�����N��md'������B�s���WwB�ɉ��ު>�^w��,p�5��;�5'J��[0�v@�<iA�T;��{�s���٫�{��q$��"���v�����/J��q6�A�_	f ^��!Y��{.��r��`�����������z��I5hdC�H�b,2V�w�3�{6�`�C����@�v@?y�������JG�*�����S��ޙ��V�G]+Q��螤6i�8[4��q��<�B��v���;g�)��g��y#��D!}�{B��r�2m�@s�{v*8Œf#��P�~���w_'ɇ�C�*��y�h���V-����˅����s�%^:�v�eҰ��0�s�1��_1��OZ-��J64c2��x��(1�h ڧ���:���u��ʱB��T�4��N�Z�RZM�ﰕo�?)0�ZvGA�δ ��u\�#7ֳ�ixOwh�/^k�C���^߻�a��[�]��B�S>T5�gw��a�&�O$gԦ$�y�9����5��:��Aj��"��Ŗ廽\���3@��@3-12�:v��ѯ�PVI&X�t��]��C�8�]W\r�n|��r�EQ�Nc��gdѱĉ1B�l���6���ٴL�'xK2������(�+��*��pg_Lz�1z��|*��ZU��i�	�ˤ�V���m|���G|�����ľ�-�����K�d�=g����r����s���i��)F�2X�<��l֭�fKN��}���;�s[�Չ������]0Y�ʳ�Cr�X���f+L�x�qu� ��̵���Ӽ�u�r� ��[E�yE�S
�L}σ�3�gjW�ͳ"8j|r��fI猳*�x�:f6��%�7�$\*�0[[M�}'\9�p�E ������5d�8̶O}}����T3�	��ZM��̀���TO:w.�y���S�}���3��Ʀi6@�W}�Q� ��fBZ��r��{CY�u1�c�o݄�J] �}���ol�3�)��)��6��,�9�W��<ʓ�sґѯ*�H�6��c��ۋ���gh���W���7�p�.�2Z�j�q$ ��(�]���<��ַL�.��go-J�B����i�Έw_�'fJf#|� ���fI� ��I���kӼ���b�v�����Ctgi���v��O�3��n��Yyyw8,g�*.k�d5_[�-��&5�dߕe=�����k�Qj��.��z�)��>,A��˲���xnڵ��OiX�9����Q����4]u�d-AЦ�M��)qql88䴎�)g\ڭ��U�'قڨ�qK�j6a���!rwr/�	��y��G
qa�T�Qө���r��9^}��CꈙU�g��}�lh�4X�j����}\����<4N�3�+ݏE�{²�m�N��8�����uԺo/ТkE`�)��m�b�!�6/blV؉�:�(��9!vL�J�h�s�����Q�.�1�4.�ُ���DT͔���i����j&YY\�R�0LC���`<�'@���wl�%����n��Cg9E����Kw#��"��Q&���p���� ��F�<�\�yD��SK�u�6��]y�G�ʖ���Ŏ��ε�������"��t��.�,��(Cg���5�f����
�ŷٰ*�^\���.�K���0)��f~3ԅ��t�Ϭ��T*Wbn�c�0�=�f�� �µ=p�tcy�,.&V4�À�7�J��7M�ɖ~&(�?T)T���\�k��|Ƌ��O7d��6��d@\{]%��Ϯ�SF�H��Ucx��wD�H8��Wp���w�4�Dۄ�v���"��a��]��r#)S��Ս�*������J���&����u���y�`����a�9N�_g	����1y��x�Ef��h�4Jm9n��}�����tٲjO�5�L%�]��g���Ju+.��l���uG�s�񉖛Q�,R���Y0�a�nH�nH�sH�GL�"e|��R?�V/-`���U���n��}��g��E����gʝ�~��_4�:�Tq�n8��[�k�����Ǳ�=��Y�f��|��d����A�����k]l!��,�#*���aJ�*�td�3f�:e�oJ�IN L��������W}��o�g��M*d�]GaE�]����Iw���L��B���:���rs��e(�ێK�[��?hȬ����]V�v�1�xO CR���=��v~<߬}�s���s`ּ�{�S�J�^~��=��'c�P�
��@����C�؇uCB���0(���?*�f���D�t�P\������Q<^��o:��pT���|�V��9��WY��h�D��A���s��m�{ۮ����*�Y���D���L
���`�����w�>���^�+h�� k��{D�ۤ�֞	v� .�#�B{&��EK����NS2%s��R��
��ӏ�q���]�"h}�PL�gW>�nf%G���U�u�ZʡL��.>ؠ���#�9;�(k����ur�ry���
ݜ'kmi6B��q�w����&��W�0qo�'w�E�� k�a�zWd����Lt&U�!�);�4&�DY������Cp�:�ٝ\n�7'0�u���Ow���/��Q���{`�]��nH���b�9��j��ꧮ�'�/L�#ҩ�8���v�H��.Y'M|�x������^&]^IwS�}v�=��z̥"{��ڄ�*�ò�[���K��t�s�]u��땡Ќ��`�o{{�+�Ip�I�|r������: �EU�]߭��m9LH�k{g��[��C����G�uZ�;u��9c��k]�Z'(,}s���Rx�q��z�q�HL��]������[��\�5�
�춧v�X�pю����(cs�JS�@��\�	�w,��;����0@�ai4z.g*���}��5H(r�<���VV`!�W7u�e�yjN�oIC\�P7&�^�$��Ͳ���ґ�į�*!Q�1*��3<�0B�
8�s|�s0���@����UQ���	�x�?w��ދƫ�u���X�`e�\i/H�^�R߽=6��R�2[r��۱Q�,���Ò�T,&a_s�]��51���˜T�.� �񖖬5k{j�.���`ԥ�b��po5���n0�վ���	e?Ng�ڨV��+s%�g2(� Xs��z�5���ת��8N�+��k��v�]�7R��Z�a��L!SW�v� 5;�lZt�[[�n� �a�ŷ�J���ՒN���+��Ǫs�85_?�6Z�!=3Y�=�2]��`̒t����WKYYSU��	�����l��Ѱ�R��\�B�?�ʱCB�i��u��5�U[7�8{��f�슡�Z"�e����'RUz���g����� ���gh��Z��z��{Fi�{W�� �x��*��j����q2�+� Zi܇�=dL��v�K�цc5���:��������z�l�|0�dU�|�2����0x��)"���˽�'��u�-��+��ͷQ�of�ี$�����L�La���M�!x��Ŋg��TDWщ��5�����r�X���+,+��@,-b��Y��7�ܐ��"�@0lF���w;(�qJb������Hf9���Bj���~�1mb99�Vռ<"�I�g���|�E�L�F�m�K�%��h�>�����@�Qw�X\l�WB���*��rY�C�2�*�@�e__p�O�%˨�9�6�E��y�vyn�\��,^�P�,��+֡��ܖ�P$�F�Xoa	6�\0`��N`�{o�s�D��}��;R������Օ���8���Z�#��j4N[˚�U����؜x��-�'�%��`�_���e�M�5%�s���++"Lv���]璁]rG��x}�FG���T��о�3�*��w�j��	&����[���f縤O�b��%�g�}�X!�Oc��5]ܡ^}xb䎹���1;������o�Ӓ����3����Q8�QJ���]{G�+wa�}�8���B����V��s��|jLT4��7'1��X����?N�놂�]����x����;�0r�ڈن5�W�$�0�g��	����dHsg`��s�c�]H5,���� N����u�g��6��bh��j��@I}G�xQ���֠��x���G��}0顚�
�"Vp�ݷ=S���WJ�������@	1�|et5=VI���8�|ѾwPw�Z6;�]s�(h]#����h����qML�ʴ���=�c[��zQ8B15l�\�'�.{�}���g��Y�QR���n��F�X�����ڌ��5�H�����L�MO2��t�Y��m��8�a�p��Be����ݱ}*w�:�(Y~[͍&�W�w9��}��3�n��nJ�.v�YѣK�7��mmSޡ�FRѾWo�ˡ��+�)T,ִqG�����<�����"¸�<�p�ܗ��qB����F2v��\I|#���7jmC�.�T~��]D(�qd!:����k��x�ܦ{����&8ry8��Yt��Y�{��n�������Թyw�l}+�J�B��ތ|&�r-@d���{2����`xd������75::�\�<c��]��1�mnL��-Y�I�}	+֯��*��o��������i�r#:7�t'�}��O�
�U�B�3�2R3�z���4S~����N�Ζy�Á�e��&��Ly8S��י�y�W��R�T�kw��Vc���_�S�X��1�k�]\;;l��)LX��J��'�u$��K�t�Jo��}=���a�SByL1��������a�-Yg�V��b��GE>��ykr�Ǳ�hya<�	W���i��h�6�Hi�l���d1l��R�eD��\�b�8WQ���ft5$��v>d:�'�㵸c��ו�[�u;��ǽi�`9��'�@޽LJ̉5�_�X���"k�Ǭ�/΁�ig�[��z�)�=s���3vr���E���YXk��f:��ߍev��<������c�g4!Ѣd�'�>�Y�^��/�3���S�z�_��ɮ�*�G�jNB�4n`�>u�C�5L���<���r��9r���V�����擇f��%��Ŵ�r!@�[�����V��.tP�6�
�lD���t1}5�r:��}��oW���4�+�t��x�oJg:�|�e�V�G��|���WX�H@(�E��xbY����K�T������?]#���j@u�X���P�\K�gq����[�(8�=��-pY�y��}jϾ�3U�U\X��ʽ9*�b�`bbӤ̌�I���l��8j�fƥ{(��V}��~7�Y�L�W�������oc,���1�#pm�주b��%��N�?a��(+�Z �,.�heڄ�.��EG�Z��ˣ��z)���	T�{��_q ��5ON�ǵ	�s�-`�d����i@s�I�M��s���"���<�aR#C�S����+�=<Ԗ_!������*��x�A�X�v������k��t����?\F*�g!ۯ���0[Z�"�8y>��0�qܨ\:J�D�t��Ӆ@1��������AN���놇-W�^��$}��d�f8��췴7^�B��7�Z{�n<��[�[���q�Wx��E�ڹh%Nt���j7���]���5�]���xY��*��i����C��^��9��މg�WN�M�V.��Z@'%o
�u��N��n���ז�$��r�)4����쎥���m��^^�% {���Ӱ�i�����f_hQj���Z�e^�=��ɉ���dѬ��nyJ<,/+��@0{pS;".lm�FYR�łMV�{sm�C{���\Z�w-P��Wz2��)� ��rń.�����1Yj�����?%wE{S}=��,vM��L��嗢M�*։�pjq�n�9cVjb����0��g,��r�;�ڕ&г�� ���5q����!���<̱�w8_T�z��$�]CG@�j[��b��Zަ�ڄ���y@����Ǌ.�i��d�E;љ������~��c;;L(Z�;)/4��*�2}e�\�Ap��t���γ/aL�%�s��9�t���E۵Ӆΰ���4Oe���/E�57{7�M.<�X܆�.Fk��2��0���1��3�]��xs��j����=iVU�9��̜tR�����X�7b��c7��9`��چ{����lm�]��A��Cu�ipr�S���lٹa"%����v���C֕�����E�٭��v��ݾ�;3{|| �}>����k����_t2g58�e��6U���An�p	����儍JW�@ov
�u��~|:ޝ���Ե��X7���'���Yv�Hc]�T��;��)7�FW=}Ռ���=���w*���ےh&V/�a�:h�=8��5}��:uf����I�5�ۖ���t�V|'p{.��3�P������KC�����n��h��ț��S�f���R�e
����ƞ��M�_��pW����������u��*ܹ�A�/|}��8�p �P�˨����l�nB�p�ؑ��\����!�[E�Α�J��o�qe��H)|�{���R\���mἾ��|b#�e�ۙ���qGLx�W:�ԍ�����:	� ]@�ҵ�F�F��bs&���`����AWF.۱W��0Y�Ōy�h���	t��i�;����%�e���>�T�N)����؜�F)Xh-�W����	)i�n���J���\���|7�^�N��.j�ئ,��e{��$�ȑ�ny��	�&��h�}����MEZ@�4V��ޜRB�����m;��C4��,[C�T5���"�;3m�$�r�����e=C�-�4���3��f_.��q��vuћpTk�N�B�s9��g��Qn�R#Z]�+3��}�Z���4\����{����wc@�SW�uȥ6��A��^H���n2�����(�H��ڼp�a%%{�LS���W}��&m:��,d�QU��k6**Z.䚽m��vf^^L��0��U�-J�jv^�Pp�&Eȋ�*����)]��yDZ	��C�*#��r��*sUQeI�=܎블't,�G'v�̈�AW+�g��Qz�L���SE��䞴���wqN�!�t���DQ�	#�P���:[*2B삂��G����^I!C�Ax`UQ'E�\ �j*�UD�:Р�"*��s�+!e:�UJY�J�tU)UA��\�(��
�"��Q]2�C�z$EÕ�*�w6r���'R	RL$��H�]����'YU�YkNT9�r�Ӊ˻�"�".G���K2/V�!+�T�HT�SX�#�IШ��#�l�|�]�������m�,]J\=F��໻^'��4rP�����}��dl�k}��G�|��T����A6����t�g�
����E/�X��C�
����"�����:������۷'&��?[y����y��������	��}v�{����v�?�O!���}};봇~m�T�Vx��yR�v,q������H�
o�;���	����~��cÿ���w�=?S�N�p���]���G+�M���:=�x����}�{q��7��޼������'�=;����&w��/�ۿ�_=C�}Uu��ϼ�f��e���ߟ_�����>������������)�!:v�S��&�Bq��_cxC�����<�p����S�s������w������^�	����U�/3#C��վ��}��nC�)����|C�޿}��|C�aW����)�	��z��>���'>����m�<��I���~��������}[rrnw���0����xO=;x@b��\��b�峞�����;��\�<yt��oo���o?m�;���<{�o���M�կvӿ&�y��~{zO)��}�x=8��C���x�����~���1;����/���w;����h��
�ޗ�F1>J�Tmr��Ϟ��zT���)�L>��������w�����;��OG��P��v��C�{�xM�	��{��y�N��{߾����!�4�g��|m�7�r��� }|x��K�Υ�{Ѫ�����������|~<;������?��ǔ��9G����9=����	�]�ǂ��q��&��y�ǔ��=�r�����n�[���v����k����>\
o�H������P�xO]����wy���ţ5���_�b"01#��y�P����=�o}�n<+�w�V����^�z�xw�9܇�=�Ʌ�P���?;�S
�����yM�	7�ǎc~C������8�H��������yy�U�����L����"=~��������ݤ�����<z>~�y@��������ݧOW�<[xw+���ro��~B��,�7��������aw�z<���zq���8=����Ӈ;��{+^]���;�l��@#�G?����4bw�����������O�{xw����7�y�yL*�����~���	0�G�z?A�]��v�^��zv�󿝯^��P��'*x�mɾ!?��o֤�����(ֳf��'G�c���1@��;�qh%�!������28��pe6<��r,�wk�ϳ��۞�EBG�;5vh�ɫ�<�?g7���;���vn{�y�ʡ�J]\��M���v���b�̃N"��ym�P����U�ٴ�B xE�go+�+:����8c�#�>�E�����(G�>&����<�yM���w���6�S}����~v�����]'��S'?�X9�S�O����?!�0��ގ��q�px�w�$���ۑ��|�����޼n~�z{���_A���|��S|�]� ����݃�&�����׍��M���Í'�{o����bO��&��} D1��#�9�>��"8B6�w���c���>>���]����|BC���F�99������N'.���7��oI������s�G�}�)�������zw�i�_|]��N��;�y��"/���D|����U\���0}oug���ߟw�������������x��ɿ�~!�ߓ�aw����㟨reE����x~�*1'�����_nܜ�������n����o)����돐��@��3w3&C�u���vV{���x��߶�Wyv�~?x���S۷��ǿ߸���ۓ��1ɤ'�?8�>�'xw��-������9Ӵ��9|Q��L(v���.��toTyU1��A�!_�}�h_ғ[����߿�=��L.�r~?���C�aC���o�P�o��v��	2�O���~��i����G�����ohN���cǨě���<8&����ې>�^w��:�%�{�o�WɥɃXh�ً���������}q8?x��|O��{M{������P��A��NL.���yw�xC��~�	�!&����x�<F��'?��>���'}w'��o��9��A}�$|*+��˴)���V�2�nl���LЛ̬���{SJ��xL�'��#��N��>�����}���w�{o	���ɽ~~�z1;�k����90���}q�=8�������R8G�3��D~��[��?����o#��x~&�÷''��;����5�����hyջ�oHra����U��ӽ���c�yO���w��=��)�!>ݼ�����0����>���oI��bw����m������v���n�}d��2�Q�]�����&�O߮w�i0�=���.��tɹ�S�r}q���]�>8�^8���90�����y�!�?���x��'���q��N��z�ןA��g���G�}��?ˁ��E�q���t_I�?�'�ƶm�{���3O��}���y^{����V�<xv8���x����r�u�8�D����|SL,lMy\�����Sj�`�]˺�{Ӈ'@�WMौ��P6oe3�R�B�����̷#cY�2��V������y�w~���8߷ϟ|����w���@����~��.��!��~OI�Ǉ���&�����F'|C�=�h{O)��_[Ϟ�������;|v�=�&���y;��~��ӕV��q����.1����r��X�� ���xğ��ߟ	�'���S
�����|��ސ�z���<;��M�����;s�zq��}B�o�r���ɾ���"�ǄEi�����%lnqq����=�/�g������'8?|w�~q�9�?�������(}����<��m����]�����ܝ����~��q����zL*��|���7�9��������%�ٛ�Й׽iׯ���ȥ�$}?W�ǯ�����M�O��<'�p)�;Ϗ�����;�b������ߟ��������v�~}�ǌ��O�{�o���~v�?����~O�9>���=�'&��2��h�B"D}���G�f�k�{�{�����;��}M<���ճ��~'���< ~Iޜy�w�{v��P�s����ݾ�����F�{��˽;H_���\.N����ؓ�yq�Į��߸�}O��|s���������<w��߿}_��|�?oщ�P�I�<��90���|C��]��P��X�q!&���)��o�w����v��'z��.<���oχ���a_��O�~�=&�~������'�{v���o����{��5�D�����M���^�{�٥7����}�yW��~x����>�ǧÎw��o?-��㓜s��Ʌ]�S�G���?\c���c˾�M�\��f�jM�K���><�?_�UWS^�9����y�I�k��ztoZfto������ܮ�����P9$�������>;yM�O�z>��<��M��0s�ۓ�X<�/�����<'��Sxt�!����r��Ҧ���Ä����L8��v���N�|},�H��z7ח��?8��<����S�aw���c������<+�&��=�߿q��$��>�v�P9'zw��<��&�w����S�~�P��<����/�ޭ�M=���X�p���">�Q�8yp�]&�_��o��9�������'��<�}���~F'|C�������~NL?�ݿ�����r�p���?��xL=�<��)������Ǽn˘�!u: M��c>��=8Ln�̲�Ž�d��RD$F3ل�N��[7v��7����f��>b >Nizɤdw)Fiu��^x�ܦ-���[a]̝�ȕ�=J�s�.�)麱˘���>�Wn�6��X�s$ܔ4��� �����JfM�����9���ߺ�P�W�>'&�$G���o���]����m�<�ߝ;���ɿ!~���|�p)����<zM��bO�~M����9������>�t\u�y,�=ޫ��;��{�L*�����=����y��;�ɹ�����aw��=x��L/��<ݯѼ��������>�r�˽{����I����|zw;I�!?�����~�!Lld/8qW2o�u�[�[�}D?]�;����xw�j���|*�N�����×s��x�c�}�9���[�F'}On;��?&�O)��O�|zO�|C�{<��xW~M>�yO_����U�T.����V?c�����O$�?D!}>;}@�I߷�|m�ռ;roG�~��k� y���&����߯��hyw�i%����<�xM�99��<�+�M�=�'����=F'|OG�s`�B!��҃�p���oG����_�;�]��w�;�|��ǅq�	�}{��)��oG߿����v�q���Oτ�_�c�a_�~����o'�;����<;�7�t�}Hv��E}'�P���(�
�3T��|*�\��>w�{W�����c���|o��<��9?�8���s�G��^?!�0����|x?'��p_���|���o���O{��Ǥ��]�m���{C�nL$�W�8ޔ�������.�ǿ��W����9ە�_ۣ(�O�.�y���o�����v�?�w�'�'{���|o.��V�}{���!�4���Ǐ����ߝ�{�&��w�{?~�����G�!�e痭�9{bb}
;����>&���������xC��_��]&����A ��O�܁�'�����}[۷!�����];_�ǭpI�!8<���y����o�nc�<0} } |DT���Uy�Aξ�^�_�}�������o��9�����o*�S&��^�f�ތ�&�^\�'�>Җ����Ţ���;�c�DY�'��?L�NAZ#�1N����¥�>��U2���)���cpn�-�KW0;+s�j�	eisվ�(����B<T������ί��ƯD"�<QPՊL����RC5E��
���}4tOȡKw�׻.�H�����Y-��1YG�({n:�ɋk,Ƕ�A�!�ǣ)��x`���M>X��^�e�ڜ�g����枩��|�� ��F]J�/��x�$���`!'�����9xP�<��Ư�?�oG_��4���t�U,v%c�n�*��:i;:!�`3����9Ie��u��B��E_���|��I�L�![|�?CRZ��ӱs����[?\Bڭg!ۯ�����Z�#�ԝ*�,}|v`�1���J�8��.��Ψ��������p�Ebs����g4���Z�=K��R���u�����Y	����d��2{T�ϙ��ʸ{r�u�c�,]�]-����}J2A��ܰݐv�?��Dų/�`��@
��C�Q�B�f�3o����γ�ү$i8�o�]��_���cn�d�n�İ�,t��*:Q?O���A���`��Zm]<Z��W!n*c��7�W�'���j��S&O6��W��>5d�\�I�����Z�m�yUK�8,u}N���'W[�C�O�.G'w�3\��X�A�7'�<r*��Ǔw9��-8xΖ��.a������&:3egh�b�j�c�tS�<�ۡ'[�y�\�W`�H��k5p�{J^0]�i�57��l�'��ҲA��U�[` �s�;]O�����GRt$S�uZi��ʛSd�s%%ϴJक़q�w��� ��Y+��*o��-nS��RӉ��{��.�q��(��<��
�ܩ�v`]��tU��J4�\��'RS~���Q�*P�k�{�ߕ�>�ja����W�82���Y�W{�/��.P�}�v=��&^^�r�
�.���5�T��0@"�y����d�Ab-j�E���W���3	��Ja��2���()�iO-	�븼�T��] �	e�MO2��|�(s�3m�p�ٴp]�I�z�Q9�z���s��dO|���Je���TDTbu򱮘6�+�r�X���pb��ǵU]�����}��Li�����Ĺ�ɵ�q9.i�Jb���;c����`3�판�2��ۘ���(�y��?1C��d�uE@=�H_%R��n���|�׆
�I�s}��^]jGKN4f�a��8z�ˁ��8�X�a���TT ##�@�e_|}æ�Ư�d�˛כ����NtK���b��>;��!��09�&�Q�(`��H���GgU�y��ɋyvo�Gu����ƾ��t�d���s����V�P�����R�v�k\�"y1��%�jB���a�����3qs�U��J�n��J���G�3W��II�<ҹ���LZ��,R�r�mo+�F��\�>[ku^����n��c���<��9N�_W����uq&��͐1��K�X��*nA]˴�#k�����.�pE˞GF�)�7��k��lƄ��Kȏ@_D�H#K�'Cc8�;�R�}�a�W�ERοV��o��B��Q��v_��vd�Bs�>�6�x�y��������J�KL������fGI��]q�ꗆ���}w�	:�����On.��q汪xO�q�U@���I��`������oٞ�Aג�Ч�h�\��v�%l��۞��8-�����X�t�3&5�H�����:�[S��Oz=���ʡ6�7����z(�Ft�n3m[���Cu�F[:a��LR{�aM���6M[K	�ЇH���W=IZ�\-�S�G>���G ��Jƭ�T�,�F-������Ni��`��*G��t��y��K��0�R\2	����vtdT�H� 5���!�̰3� ~��QP�p	����هd�ɨ8}B�*s�*`�0 G�b����J����yU����J�X�Ĳ��7���]0��1P�*Q� nA�3%s��z�/,�6>�F�O8_ ��
/}���[�V��Y(�x;��Z������u�+�������Q�M�v�K�yfԱ���l��(�v�mk��v����c��)��&�zh;�Զ��X���[(^�nYut����uʛ/oq��-���A�����-]Z�6$�;��w.|�%"n�y�c.�S����b����(��K���nص��ؼ�o�k48�:����ÐԖc^�c�#T����@eD�p�s���붧�-�;��P�p�Ҟ:��r�W=ǡ���=�Es����)��)	{+(�N���l���z7뭂z�d%��j�`��kgF�T� ��E�5�����4]�����ؒ{���K-��W��u��ᨅ_#ӓO���W�����^�l!��,�`�Q�J��ʺsg����Uy�GTh\�N�	Wz�.�N�N�F�%#z�o�����t	(Ŧ&(�.\�Q���JȆe��"�F���m��؝Ȼ��Q/tn*���;��j��IOF(
w^��<�Uro 0�cY4v~���~Zh����a��(����-s��z�˥)��)�{up��Ӛ� �Ίc���\͈�e��ޱ��s8j��V��PN�Φl1�]O��ҙ��w��0��k+y��W��LM�#�{��#�E{�	�qY������k4>C0Ϋ��]��TC�PVL;�Y�.��˞^���6�C�/7z��\��Y�h��j�6��C��];O>���q�ϲ��w�q�Y��V��࠭��ؤ�I"�����E��:��TͶ"OǸ�j��c����舩=,�.�v��Z� -L1
%ͳ��fWP��:.��+�e{�j�0�!�TvN�P*�0?��;ӟ50x*��s�X��>[E�Jt���3��{<;%��M�-hy�֛��	����������mܕ��[��S[	RO�D�4���*O7=��W.�1�����:���,q^a�=1M������M-���u�BAf�Z��`�OLh��u�o-ѱ�)�-d�$�@[F�#�Y��~4��V_V^����d|�:�^)��D�	�|���jK/�E��Z��>�}��Q���@ֳ鴷 �l�p@@�FwL�~��Z�C�_MC�8`K.+��YV9��v(Mn>�Oi���[������a��먁�<��������ދtE��O><��7e;�YPgL7!�B3ԯ�߫����n�b�8����In�{>tdю���et��t���!���$�§�d�X�Τ�]"bٌ��� �����jn�G�E`�����_1\��UY7�[����c�Jd��۸�Ow��+Ua�א���j���1�b��:�
���Z�h.��w��{�����kXy�5"^Tݧ>�ü.�ƶ�dS_N��/�I�;\� ��C4s�E=�vGF��a�s�l��.ծ�O\�x(�}}x�Zz�8�_�޿���!Q��<ۮ�4�/�pJ�Rf�Q1 &BG
���ۮ�{�D��WVu0��7��\n}Zj���)�%� kP��W�b�=b�Cyw-,��{>Ӌ�.�C��;=��}lX���ϯ.}���s�%c�.�ՉJ�ު;�s���ᗆp�q�:`\���L`Td<8'��1xPc$�A��>����N`ų֞��6�D���n�O	�t��mf���s�Cl�D7Y>dQ�v���@J���8��m�=���>��1�_���c'��S~Ͳ�����[B�'v誘]Q�ŠU��_`m؎ݼ����vQ8�� M��HϩLw�ɧm���� �K�phr���.8��mX줹ZP��Ek��t�!#t��Yd�y��-��+s�3o�u&�nN�yQ��Ѳ���޷jI0�'F�	���)�2�Q��ˠk�����m�ec�r���#�������ld�f��k�I��Dk��o�0B;�Y��(�S
�L}σ�1�Aw��dVc�ޫU�lS*Je5n���&��2ڏtT�ԟ�����|�.TR���c�V����H������&��o.SE;F�r����MLkO��`�2�����V�e��2��O-�3e�f�ğ�凞,�6�<�'_`	�*��*��]uE=-Dx�t���(&�2��c�����^�6���9���<|����%=�Hg�'����~:�}���7�5��X���}�AL�n��y˨ƥ�:5U�lc
��NM����񾻷���:�����"�AQ�B����{y�κ����K�r�g�y�F�I�� �0b���X2왏u�H�����D.�|+}��i�rh�δ���z�e8�_Kco�}�����\�
={�R�k���t�z6p�����{�.�����¡DQ�����Fi��4;L*�n���Ȱ��]l�'{�n9���/{c��s#�>�r���|W0�M���L�|y�%�|UҖ-[�X/p��ȑ��1�;�7�*��_ou���b1R�����-%E���mV�o@:���te24�E���o��6�鹊�D��\n�z�/.�X�P	�!@�E�4�Z�+���yO���D;���n]q�k�f̦�cM0VfL�� �8��o��k���3F���՛W��M�|�8 ����m~В«�OFyvU��=���\�oӻM�,��:��^�V+��9o�۬���ۀ��0��H ���ejծn��լ]OV��)����r����9i2���մ�«q������#�6W�Ӌ�v�f_ëZF�in��r���OC/$�mUј��t9��+ӓ �lܼn�M�<O�@��	�V��D�%T��݉J����C�'$���4��X����b;�V�m��$��]^Ѧe;�i���ҍ�����pn�pc.L��<�WTW(GlK�hݽ�v��0h�5��g�O<}kg=�������!��5g|�T�X�\Y�DĞ��j�M��ݣ�X���gK{�)j��ւb���l�}�
�5�;�s[�W�;y�Oʃm/7Nr��_��N�� N��ִS�k-�<��i��j��n�@�+��,��b�5K͕4qL�	ئ������N&��w���s�����c�Vqck�+�:�5���N��Q�X�]k�>�;��>�ܸ!�ph�^�� �3\�uB�ww\�ۑ����um���V���*��4[���K��wWX�Ѱo���\�QfMuv���nћ6�G9�7u�w��:����:����n*A�`t�8�����B ��k��Wt`��=�G���ZWʗrד��<#Q����l���m��n��ՊqG�<w��*��0x7�ov�n�M�>j�ͼ�ʜ[#�����9��@��MJ-��l��5�ԙ����u��r����3�� )�%\�U�7�N���EF�����r�(�ds�"��1L��"�e4&W*.EfF)PEG �Q��*G$�v�br�%IURBUEª�L�I%ʂ�Z�(wwVAh�E˖e\�(����=DU\(=e�p�"dI��M(�d�BHUAp�e',.�QUD�TTE�NH��Õ�U�AQ���&Xb
Q��"�W.P�����ABABQQr�h���Qˑ��9*U�3�V!e�ETAp��"9r�tÕG.\��*����:Bejs%�FfHTr*�Er�"�(Y�N�IL��AE��.�"�rE���$�R�F�
+�Q�B���EV�˗ Ζ�Qu�\�#R
��QQ�Ҫ�̮��"Ki�SC��D�i%TʵT�I".U*���^o)ۘythSr�r�\�I)a�L�CVWq���V�Lc�M�����(�)A[���S��;�5#w��J.FegXK���X�Υ����{q݅_�R����̨�{���J�7��q.���]4�žW
�"iH647�\�c�8z��8iR�V.J5�}&P`�ZM���s�m| ;��3su8Z}!�k��t�83r��Ct�x�����$yK)��y��qɝ��p�mJ�j������D��k��t��3�9���o�gv���w��ϳ`�ej�W�����@��������a�f��iI71�d�%�f���殍�"-Os���l��d���Ղ�qT1B�"��ƩZn:!�|jLSIٓ*h=Y���X.{w�u&#m�� ��fI���՜�mU�p��R��o��+�_�w�1��o)����.�I�Ʋ�\Cm��l|�[@�P�1��X[�旞a�|��Iw�W���ކ�6n���F�1bh�Ӫb/�̬��,5ĉ�]Ԉ�" v�[��	mL��b�XI_U��	9�\�EjH���b4=)��j��<s7��u0sc�^����],1�����]쥱Rkc�ٶ��ʳ��'[?sc;s�d[����^E��P覎�ـ&ϗ��Zn����O"n�1P&ޱ]���i�������aW�6��2R6y�ߗ�b��x�:X#��pb�콾1�	�H������>Im���v̉G�nX��EL�^�|�Ҽ[�;mv�%O��pT�v�W�_NizF�հ]^E���*b������.���/�uFt#�)G] �L���X*�6T�/3Q��ᖸmݬ���4���<6*
�ʂ���0]2��:���fV�;�� ��v:����Cqs%K�aM�q�S2���+�������[�����u�].r͏��ٿؠ�I�أo�-<z��(E���|1i��ӿ���<=��.ah��I�W ���mn)�����������?WХS»\�z�]ev8�6#�DF:K����[<��7j3����=1�*!��U��![WfY�7f�8ܑ_7D]9�gs�d��Yy3K)7�^�7{�TQn)}��k7�M�Z��nF,��N�?�H�3#yS�o�qQ�jy"�Q�W�⃮H�+-}�BG�ɋ���caz~��[)�u��p�s�dm�=�2V�ӎ��3�T1 r��)���@�~ЫNH+z�M��UL�͗w�o����6B1]��%�0k癡l�!���M�6���ظm�Y
��U;h�;�V�4o19K������ҷϫ�ӌܷW��u��:hѯ�ע&�C� 5�Wl��*�%�q7ٝ�	T����Wa�$<j7���#KN�_�����p�+�`�0h�?~MS%�3,s �N`����M#֫VN�����[�[g�C��tgBN3�8EC��&���Da�.㒣�n%B�<���2�1��߇� 8�n��,M��Ubz��)�&�Yb��t�YсY�>�\��FF�L	�O_42[ɋ��
����6������)�g[�������q��U�F9��C͕�G[�[�Z�9�iD��hl\��l�DEI�b�s�P
/Z� �j��ep��0f9��ѝrc�K�'&3}�xӬ��A@6A�����w�)���^Z�+�|�c��֊]7�d8�J��خ��%�^�U�=��hv�Ф-6ǭ�C��^c퉑z{��}��Gp+���	ݏ�7$T<�n{m���u��Ȝ����Fwd  -�*��ͻ1T����珵�)���*cI�����@�ON@�<���	�r����� �16�^��}O.h�fDyGp_�,P�p��¼.�(�lК|��Ƥ���`�2���p�^�����xMHh��˾1o>yIL�r��;�^O���+�v9����Ƃ�+�2�)�'�䫞L���wK�t��U�ݹ�c:�їu>��h��@-T��
�l�R�/��s�IN�m����f�@�Bӌ�\�Mt$TOD���"-�h}.���W�lk�K~<�ޙH�p��Y�v�騇,;7�/t�7��{΍�;N���V9��ά+H�J�1zlnM���=�%�����Qz?LK깊�~�=�ՙ�����F61C�m4f�A����X����&��,�OǟXly	n�`�ϝ�c��2,1n��R��.�u�r.�n��6�T�0ٌ����T��BՏ�A`�U�{��{�k҂�h�w�����&1��-��Z�i�8_��
7\a?J���n�5v�ˌ���G"�O�m�輊��v�Ʃ\R{_wɪ�-ɒڐ57�b;�ꎪ2\m�f[�Ut��W�@㿥��֭h}Պd�f-u��5-��cW��']����O�=���^��Z>�0�:(	L��1a(2\�����A��6�r�"h������B�����T���dz�T,�w��л��슡�b!��EV^���{m���kp�� w�P�3�t|n��8u4[]��za��c�]�����|:IZa)����5QO�1�����h��{ೀ�޾���n�uJ@�H!!֙O0L\)\8���޺�Z%e#m=A�9f��2UW��ͮ����xS͌��p�}��1�I��,4��K��"Oh��x��q0�Vݮ��0�ǝ�U��_M�v���o�.�8zf[%�@�`	����&��n9���:*/g$�}E�4�lʘ��rkp�.��t�ܛ��h�t�Yd�y����·<#6[��RU4*���b��_��rWzu�g��KDZ�����dS�'�ҷ�������7)��ƺ�Nى�E����Rgýe�0��q�JY�ɵC=�K���E�1@�˝���C�鉨q��*�����m�v�5p�>3l�P(G��TTP=�H_%R�n����<3w)��_i �	6���Z0���p��p8]GK�Z0��{��FG��dR�iIΖ1]��o�xdn�||�F'���p�9O��Ct�l�0ꐚ��OJ�!]�0����҇�P�󂶴e2�D	�8�.5�NR)���}u�7���V(�Y�\;�z�0���vY=C�F���I�g�|M�g��-]��͍�c*!��%�!�M�R�y���|�i;����6x�X�q$QJ9��8�����a_B�D;/�#Hn��G�c�˒��+�S�QI%lo��-q}�H�YD��c;����ܝ�4���sjT	���(������Fv
$j낱b�!Ǔ���=9�<7rt��>�Ů^�*�[-���Xܬ�G#�����"yN	�
Y��ذCo�kMI����ͽ���:'�>��#U��&6]�!�����j�{�mV���3�tY^����ؚ��Bum\�P��߬<]wB�dy.�y�C�6>_d��x�>U:���f{Iؙ��n.Z�?[gκK��S��qj�L���g��Ń����r�H������/I��-nZ�J7f5�T�Qȩ��;Jefڶ0�̷?4u����/Ew����a�3��j~ڒ��pt��=,�DT͔��T��Xհ
�e��ų���f�:NV��;]�#���4���c��6l�/B_s����MF=��ZUxS�ḚQ�b��m�t�㾷Z'9�MslVJEy�jn�a�K"�T�:�[�m�!���.ytpv{�_bd��et����:!�)��w\a��;�������Es�j\����6=�hn�W��f��Q���­��n�<Cr��u�G��x{Y,��#`7�Ee���]����7�x%ߧkcƵ��f���*]����p��zq���n�6ƀ�i4����8���\���C�(�촎^���Ю?I�������w�F�ۥ1�F9d�[e�+��~\�������5�h<����2,Y|�tq���W�1)q����I}Gj��5'd�f�r�`�s:T\����v��\�䧶n�Ͱ�����y��B���~�Im�B_3�72�Mҡ[W=ǜ�1�s�����j�Q����mvK�"�����Η��R?���� �99pިݶ~��n/�!%g�7J�ݗ���$T�F���C�=���j!R=�L_ϣ�6a���������+�� b���NQ�Xj[��l����0�T�Q҉�����i�,Z<��!��y{[8�����]���k���8�VB��U����Y��jI��gf�B�l��(�)��k#]Ѧץ	#��Z�*�R��&��� b����j�@v~
�x����1��k�6��r�l#qM_qȮ��g����jI���N�r�>�c���P���!�u�=�ec*R\2���j��E����#ͻ�M3���y���*a�c!��e\^˾��vz�%���n[�\��6�(���W?�,�yg�����w�@:�}3��)7�vJ~;���50�F��X��m��=�N��֛�1�U�0.����P7DW��O��LK�X-!Yl���9w2��'B9U�\�Ĵ�Z�ssr+n"�Ǐk����D��:fq*3�(����c���(WT��n�q��&V#Z�N�%���na�+3�V��[]oR���RXubSu�������KQ9yD�Ֆ��}_}U���j�=�=W���ϩ��%�g�[�4��և�n5���'��EMk���OV+W�6�Mm�&{��UP��nH�����o��W.�1���}=��˫P���*E�?e�ͷ�/��}Fr����D�<$j��Q�^�+on1p�Sjtw �i�_X�n����-�Vk���IU(	��=(C�44&�+|r���D1�6Չ�z�����K��x~����X4� 1�J8�3��~Kj���n��X�`e�~֖����d*I�,)�J�i! g3�/�v��
�5�� ��l��a�׮Ѽ�0�G�(ם�JW{#:}>��t���-�Y	���Ê�X'I��z���Y�rsmN+�o;�no�C26b��pF
I�C"�DķK����ge҆a�7?����,a[�� ��|�o.��I�9FY�v�+����|�5��^D3L�>U�-"i�&&#-���Ϊ[��B�!���ݽ�MT�Y��q���_�=�Jdɶ��'�sʧM���:/��+*
���l	-�S��f]}���Hż���
)'BŲNih�ͦ�SV�%eTJ~�~��^���sW,�����x,m�<VX�Aj�@�u�!�^��N��wD�=��N�
�эeM�P�11c5^��;�x�^�����u6���꯾�;ǭR>>��~f,�;1ǤaB2DV�i��W[B�!��Ǫs��W��n��Mn^�oS�{�N?���v�e
���0��u�X#({�q5x`�R��̝�����N�8`����̵Oۮ�f��;w�+8!9�W�@��*����dK��v�'�}�8M�D�z��ȩ��g>n����43NDn���_6*pW��$��^P�v"�~�*	��*�2�+ L0�i䌥0�!��q?Mw]��W��
=
�	^�bY�U�([�� ���\���t�4l��Z:������p�f��m�ל��	�5h����}V=^���_"M"xy�KD�zߒ�.6E<�K���oʇ��x^3W���Ď5�V��G����1ZW�tQ���A�� T�@�k�^9W�E�1@�p����zF�q����R`���u1�`3���}�fو�82M��`6�H:�{Ơ�D�k�[z��������,.�\a��8z��8T��J=>��e  �)nAľ���
m�\��C����f�zɥ�My_T��Tl`���qu��\�/�LrP0��}�� z=��3�7�����hs΍P^�Z2���-W.�c�Q��p:������5���Yω�;+N�t�ie.ʇ�-HO����>����[�w����&;�̀����Ĺu:�>:���TC0K��O(��n�v-����� �^���v�76{���q�\k�I�E��ش����w��w��tOZXa���k��{��4�!�IHQ���Y��K��o�c]NOCs!�<j-��,6���N�Z=�O���`�O� ᡥQJ��C��W�C!�j�)����Cx�-&��|9cڨ�`�-��OH��{�9�3Wk�Z��#�a����p�p���R��x�U�7Տà��bK�Z`�	w�hi�P��S:ẠEq��䶁x�>t1T��-�񻫕yV������u�>�j'�,����lh�5e����"�:�,P8v��dE�D���S�7����]7��شY�P�ꬶ��#aL��V�9�n�h�UW��+?~8����+?)yt�a8n{E$1�K��*fʇ|�Ӑvb%cV�ȉU̲dE3�D;[p�#s��w[��KZ	�~�,�uB��`Wy9%:	}�k���c�e^�����PW�fy����a�ior��<������v�������͸�]�/v�5��F��,��k�Ҭ��
2a��z��{h�R��S`D`*��Um�thv�.V7�+(�a��A�GC��d_3�[�U����X�_<�=���]���*Q�u��*Pv(�qͺ�����򁺀Ʉ�R��{� �;�j����3�SS�F�}(h�cdW+vW�5���T7�-����	Xmx2w����v�v���(s���/�w��_n=4�r����[Nd�ís{C9m�rw'{w8�����C���>�H.�sʺ�G'ت�(e(�]�k-�y��K%��Cu���=��a�w�y�D6�c�������BF���>Y�ݪ�����4�j�������p�㫱�y�Y���mM��n��c�\뤺�(#�Hc#�ڒ�-���h^J/���z��9��
�*r��u��q~K8J5�!�������_���[���]g�R�
����v�tC�*�/U�R�#�U�ʮ�=����c����ƭvk��;�����fC� �A����ڴ��ǗN�$c�Is&�T�n)Vr�3HXxiIϫ����4��C[O{;�*�Ȏ[����Եn�f���>iݲ�<9w%MƱ���C<q�x'�Vxo1+����Z�VUΗf;V^�t�x��(���Hq��V�����EO9fXįd� ��Q�*wWo"�)�r�f���of��euF��i,f�d[Z�zN��5݁�u�%��%�:��]ؖ=�+��p���9�N�i5�8�Bo�MC՝Mhmv=���0tϖ���y��z������!�������E�R3T�S�k.mm8�U�$R���8�lI��^�6�F�dc�r��l�^�Æΐ������[���l܈�1,��̡��p�-�E�X7"<2�To�l��6��ڬy�����&:Uhq�W0�'%}Zv�is�j����m�om��7"!}��	E�5��q��|ok���놘.�4������sz�o�Bkp��+�s2�7{�Y��5n�Y�~KT�3��ޫ:���OxFV��Is�u�u�͚ۧ��ۜmDm�K'�$�M��p�әF�b�ʋ��u�\��-�B ��c� �)���I��2���mt,�ƖwOr,MP�O\ *�8πLAʚ�n#X���<�o��U{n��2�]v�Q��;��R*�ˠ��*0v3������2:��ۛ��3�=���=����5{��5x�[�H������R�,�J���We>Z�𰨲�����Ws�����ہ�h㋺=ۋ��eh�Nă��ٚ���gR����D��<5��(\e\�gqb�V��er�,�Y�x���2Y')lc��l94�/^
�Q԰]t��d���������o�2a���2�k�N�z��G�N�D�2�UB��@| '�e*,�����$�)e"	�Et�#�m6r*9�:	��S,���jr�*��PQ�p�Q�p�Y��
(��öTr(���fsZ�i$��DQ�"�UV�QA'�W(�����)3+��]�*$QT�!3�GeUP\(��tӴ�\�֚�A��PE�� �Q�
�����(�E'I�jp��C�Q�
'(�R�2	���+�����e4CHI
���)AM0�gNEQ
��0�92���R�9��b��g
�h]g
T��J�Ԋ�U�G"�(�Aˑ'i�E�(H4"�g"��� j	�\)%0�
�Qt��B�0ʓP���Z!iV�E�.�H���F���&"�D����=���n>���x��K���A��b�4�ԓ������9��6|�M�G�ALs��u+�J����}�}I�5��O#������/7��``��PW���V�-�<)�ٷ�RL�{�W`����L�@��|9W�W��:B.��dE:�����I��kv=�?���DMz A��{ܩ�q�S��͏�*wbsu��0��{D=������5���h�|a&G�\�,��w)_Fcz�N ��s+>�w�����|�SÐԖcm���я��S?,����u9�_]uJ��:���'\9 -�����0�V�H�SC8�({�9�c��H�T�:�[H8��������35	 E/����y����Ʃ��_��sv�{}�X ��TyNf����/�� �\�4��V
r*8����=�tZ�V���BuL1�)a�;7+K��4�q|�;ǈ�~���7-Yf �J�_Q�4��	�A*�]�i�ţ̥;0ȅ;B�+��SX����}��_ϕ���=G���L����W�0DpD�c. o��zʵ�q�I^�}ͅ[�mf�p���-��5W' 1�7,>����?V�����e�0y�^�2�;f�h{�%�����8jQWua����W�Z��B�
��8umNr
$�������(��f��-u��bc*�7�{&�ۧ�����4�FR]�]���(]iWd�"��<mڨ���4�h�r�╺�w ����������3������\��V
�Y_V��9��l�r��Q{6#�wzr5:˜�M��J�,�U����	>sw6=��Ĳ�xWF�cѥc�/��q<szS7���*a�b$����`��{պ��V�D�j:ۻ����HŃf�4�kƠ�a�V�؏�]����1��uz�ƹ��źm���s�8C�sl�D7V7����J�0��|e�V�����,��wY�둹M؜��vݦdJN�
]6{>W_f��W:3ngMK�~��<EJs}�4�w5b)���I�J�J9��nHp�y�툷LB�u��Ȝ���۩�-�{�wk��岽��� �3�b-�,�큲Ǆ��D-Wp�:zph�=�LJ�oh���C���j�=��ѹW�W�	;S,	���\WR��b��lК���`�`��u�o�É�>�����BmS�ιlS��6Q(�%�-I��2�L�~���k8�����R(��k�ȗ�c��8��2��}j��
�T<\�s>d*�ji!��ދlg�ꈞw����7&�wJ�C	jmL9�29�p�ǃ�J����o��Qz8�gw\B}�����y��[�#f�<�'wϱ��=s�Y}�g?��L��q�֢k#]A�T����U�C�r�ل�����;,T����������R�|�t�B.�P��M_��9�Ȇ븛�n���� qY ��@�'��y9U7{{6���7���R���Lp{�F-UX؄��r��"�%q�:��\BX�͉�:Ԑ��k�W�Z/��A	G"�Z=y	_�>Bc9L2[o]���]۾�݆�է�|�
f*����A�d-�a�'nmM4;g��7�O���UTZ�ɓ.�Yc7g-io�8�W�k �qn��Og��JP��+k��uu1k�鯡���40[��Ľ�4����yq�	O̕y�����^��a�4��S�*�=��}�k������z"�*;�����]�ࡒh ӧ���Y���4$[gT=�*�s�*��~a�bY+�ow�j譎��X;om +��P�"�ٞ�뙎fE����m�H�(��S]��L�ջ������+�z���:�|��%g�a�&�O$e)�ɲ�Zپj�GQ��z-;��Âm��'�QE�,�S�w�n�Q�2��1ٻI�}	j\p\5<��0��]��\i�ˮ�������5�ƖX��f����������N�Γ(�E9���RJ��ںUbV��N��h�=�4���B�c�,N�����s�1��o��X�Rh\�X����ǳW6��g��TtqnX{ٲ����/Vսsx�T�����oLE�?n��q3���kSd9J��$�'��tL���*�ёO'�ҷ�����O�G���-�P=.��F�ҙN�}�'q��E) �@@b�b��ᯰA�Va��݅j}ǣ^l0�cV���:C��rj��|f�����#Re���y���v� 3��mg���3��E��!�#LG9�5u9[1X���>�����Dh�(���W�T�m�5�. ?��� �g�)�B�O�&�t�8\9�|u�ᤱ [��!/w{G��=!�.��f�c{��p�"G�N��+��?_]��|���|�tCg�`8����e�Pt*#�N��k3����v��%�!F���_t+K�<);ʽ{,��Z��s|8]�Wd�+Aꂴz�Y�g��D�H8hiTR���x,����W[Ӹ�v�v*軛�Z��a��c�9���&��7��k��X� TqD���_�Wa��Z��e$��¯}��W�7ѝ��ل6����\$��Bd9��h��WRKѓ�7��aF�ݑ]υ��73-Nʛ���[�uv4�^�̤wuhɖۡ�* .2ER��αg*f�>͊-�ү��-���i�I<��Ol���g�
��=D�
m�����d	N��9�ba5������j�s��\ु��������m�m��梳ޏ�z�E)b�޶4_�j��ULE���fVD�`�bB���(�*h��cS������bL��f���;��h��*;e3y���;s<�|ѿ��Aـ"�(�P�;���_}N��40l�|��}S6T;�Ģ4�lBƭ����d��=�����SZ�c�yZR8�w�q�;��\��˄��T����:1�Ǣ�:�<��3+���u�=Or949ԕ1^��S����^lyƝa�p�PW���V�-��:ki��p�W[[K�v��QN8��� k�����Br��u��7�5vT�B ��?&[���6^�R�Z���:y�T��l|�+�
9����c/��;��|���YK��J*K�z�('{����޺5)k��6�fX�Z���B�O|Ԗcn�M��#\P�m��6�3��nE���Y1��4|$��"��0�W��oV��Y�{���a�w���	�+8�E�E���7�q ��Qy��!)��CT񂲨A�^N|;���&�ѩu�nן�����("H6����\}u���RC�E��c�����Q��*���Y��a���U�
�[h��\����T��U�ܘ��;Ђ8��T�7�76-R��ha�cl�d�������X�dI+�
ٽ�	��;�oy��.�VV���h�k���y*�O�Q��F�C�=奯��#�Ɍ}xo_gxdO��[����I�/O��i�-Yg ��~Q��@>P�a*�X]���f�ufj��uEӞF*�] �>|��-���CJ�/�<��N`������L�� 3��-S��c�"�=�8����L1�y�"�<�15W' 0���]��U��6�c�L���{���%s݁����'�������}�"�R-���1���lGZN�Njt�8�`�x����y=[3���޶í3�5@�^����$��m�Ri��W�+���t�u�!~�$uvz�Ê���m�2�Ϯ*�oh҉"��W:���7v3��h�O%Fr�dj́o�zO�R�0n@�͸A�UEĹ�w��ռb�T�`���;�Χa�&�r�ݣ��E��=  �ŧi�I;�\K��*��¹�Q��:n�%��p4��%�,��W�����q���	�:��;����䊇���m�bĺ��gӕ���Wt]1mJ9�s2�_5�u��͋B���[�ֶf�7#���,��������'�ǝ��C�h��S���U_0 ��O(X9��T�@aV���JtV��0�c���c��허�������=��ʒ^���zR�jQ��^��`�vT�9���b�� �P��fo{ޙ�{����u�G�/�`.Ҽ>ǋ�V!km��,��φ�a彸L��y�aZi�qŦr���1��!��X$�L�$>�WԄ1q�`3A�B_*z^h���X�2Es�<6�9���m}o��i�Ȕala.N��6��X����W��_^��P��k��(Р��'G��H�Rt��Վa�Rx�J w3�BF����q�	ޜg�5��f�͕���q������(ks�OCuM|%��8��*Hu�sS��Υq��A5��{#ף��^���-v��0W�5h2��c&��˗I������W�)��gi�`�=�?oG�	�����z�K������ttɨm�ؖ �2j%���Us�Y�Ca��W�B~@���/��z/i���q�WI��&��ˠ*S�v���hFBQ����5d�\�N�ₘ���~��l��:=��%�O��kUͧ�ƹ]��?2U�o�u�aXtP��u�X #�l4ռ���Q�쿹���u�;jjųq����la\:��p0	��"qX���~�e��k��p����޼f�Ǟ�� ǡ��8`lÞ^�޵Tڨ��3�����Ղ[}f����DeѮ�'z�f95]�ze-F*}���+J%�	a�F�E���QK�_������ަ����s���t��ѰŵO�=��/g֝��ߩ��� J�g�ۘ�<Nm�5�n�^K��I�O3)�� w���]C��g�f.#���;���|_CԤFOv�)2�,�|y���Q���+�L0����0�7X�[7�W��-UR�M���gG��b4�g������u�O�v��U^��:�d��h�/Xs��6k�7+Qͷr��|��R�fڨ�1�rp]�$����%�]=o�U���d��Kз���ݔ��=FWH��\B�{�')�����H�c�i�!�\E�R�drmP�r̾M��e˲b�i�yܣ��E�)�7L}��:C1�u5P��ͳ�+����O:*����r����L���{���2Цc��{u�)��"�K.�h�>�����J�Z.J*ꎴ��σ�Gr�^t^O���+@
�k����ef_p��O�&�t�83r��D?88��2�RX�oh~˧�$��wltȖ�N�G�|JU���\^蟳�Db�_RN�,�٨}#w>Fr���O$b�����b�Qt���*U/�C_�k@�l�o��ț�i�q�����CP���wv<�S���;�f��
�Mڵ6	)wt���,޼�%��j�C�r��b�g��{����7i>k3�د���k��.]�"�X�?}^�y��L��伾w<�B>�J1�1��6M j��\*�)��O��f�z����Wjl���a����*�Y�}�8�W�*�W+��8b+L1�j�r�w���n�K���7�$s/�I���'�Nb5��26]�%���b�X>��F9Â��S���v�^�]�AI[�Z{W����Z��MZp�ClmG\�ج��|ۙ�g�73{Z����N�S+0��ٯ^ջ��{x�xC��++�W,��-f�"�ރX/�O���b��m��ѵ�v�W���x�7�8ؙ@��DL��uN��5�L���n~��7�x]�b���˓�@��Ɯ9��i)�8��NUv�-S��9�z���ηg*9�ʂ���뭹*}HmOm�[��l�4�αI�`��J�>��p9/�	�jY��o,���uIl]�r�7it����_ɧ�/����=�RL\6ē@d�S�|f�s8�e�[U��%�H��6@kD�'\��׬���<�4{H�s����9^Z��I��hO�Uf�!Vw�w��u]K��/8@��@�=��ԗ-�Vy�������ibRXz��u��E����%TP��:ю���꯾�I�b��<�� �T���éJ����ކ���{_&�٭�3����ˋ��{��j�p�'���+i%q��-�ߡJyp�kn!�z'(�\&X��i�;�.���NF'��2K�����*�/���_P��m�ɎkdJMƌ��q���c�g���v|X0R�CSY�ud�B�.���^� ��,S�^I�66?)F~�9Д��y�F���)G^V�}X�x_-�;�>6־p����q�p��Q�����ѻ��UW�p�-�d��h.t������=�vˍj�:"�L���T�$����@���owt�YK7��s�p��i�=���+�$�O�å��e.�k?{�Y縼�Q������������K���we�1�xN�8���[�9�\{d����q�⧟Ԯ���h���M�ny��� �s���{滲]�(�Gs�*]ai5:���z��RL�u���F�֨wb�9r�-�C��U�'�h�>ڏj��x�z�R:���Yœc@�V����5�;���jTXP$�<Qҳ�}^uzp�|�'ky�?O�#?4�J���:e�= �}1ݽ�em�z�Z*A��6���knͧՌ�E��Ѯ�������?=��҈b��i��(�2�v�ֆnsp��}ܥr���8�I�b� ͅ+�����Ѭ�s��{�n��;�.��g�B﹋x��$�2[24x��Uz:�v�sx�Y�ˀW�=���U��O�]I����0��������836��-G�ֻ�D��s+�,���1���`,�f�]/1q�jvm-�U@H!�sml�ooc�ǁ �����ֻ YT2�
u����:�=b�[����pp�ؙ��C�k�S��:�y��)eJۜ���j���mWK%��;]��8���d�{m-�6l�]WAE:����n# �
�՚�h$�-Y2�{$�����k郇elW�J��'g11�D�G��x��{�zG�b��@�wE1�7inluf��sqA��s�D�w��G�o}_�B��(��%���y��Q/P"���G�-* ����n�ZW��w��QG�%],76Ć7���DZ��o��;d��
����h�=kPK0�H���
|�f�W�mm�=K酚�-�n�K���\������8J|s��.r�7�75���f�)h�q����v��ҹ+Y'�*cU��<�r���s���t8D��\�;Jr�־4^�8\�Z�\�GW8qv#�m��O��G�/���ۛխ�o,��U%�w�`�ն~ǎ7���-k����'VS��w� �\�q#	[Hl��*2p��i�y&�<
�u4/�K�r�Ga9�.p9o�CSS	x�H�f�.����,Q^K&��y���z.���Jgx&|�l�M,�B���v�c�2�Ö��g(�횊�v_`����Mΰp��M�>�s:�nw+#��D�<�nNλnP�Xc�--mˬX��,���Ir{��Y,�w�l�Y�/�Ύ#�}K�����q�t1_/��S�|�C�����L�ʡ��:N�Ir�T.�VZ{�Y*g|Q����|d���)ˆR��%�۵��N����ݱ��G��K��p�f���4�k�Y�+��ѻy����th+��K<��m�}�<Wx���F�j����2^W!GݨYfܮ��@q�:��\5��V��ģ\1,�L�٠�$ۮc����dno9�#�Ǖ�r�+��rS��2諜���8����v�z��c��#)�n�^�,V�&3֖w.5�a���5���09�è���a��9[�u��-�+��r�u;.|#�Y���2�����t�`˩@�reTWؖ��B�;y����cs���VxN��YZkm�lI�G��  ƍ��ڕd��2��Ft2�U�p���P\���PA�*�eAF��Ԋ
�NQW*����h&�iK,ȉ��uk;B��!�a�͔�l)"�,��)9����!0��ɪTPU	�Qag,(,��!��KB�D�l�8��NTI*Õ�.�bf'�a�\��,�D�乪\�Rj�MՔ:�r��jEB	&ʊ�+�Y!�N��eҐ�U�b'��\�9����5dEQAr"�&TDat�#9uRjYDE�Ք]�G*�Y�"��Er��daQ&*]�ܰ��P�J�&��*�
�M!5H�$�#V�r�.D̐"3
���E��vh	�9I��u��(�1��B�$绔�8	 �̇�G��ۻ��٣ڊ/�u���[g0����	+��c�%dBl��$Z�d@#vv	�yֲt!wY=���}U_}��mN�}P���E��^��{m�ǎS��R��=D�3u��^�9�t�z���D�9�8�i�\ظ�o[���ٷg+�̢�qV��US1��P7�5IB�;ӮOBWZi��\عm�ߕ����V9(ͽ=��o}r���G�;j���~i��T�C]+�����/���%��i}{r2�[g�r���j�����1 ��e\WHUU(���̴2yl�8v�`�"<�8}57�5:�}T�ڹ[~p�O�[��Hu����C���܌Ґo���n��o�٤�P����s7RAu�\{TeC�V��������Y}z����gT6.a��C���Xh;a8yQ�z��c���A�s�w��'�nZW���ED61�o��	y.zl�<㡒yH߮���NlMow���q�I�l������@3UQծΤ]�
Hm�-�cJyyt>���1�dz��J�Y�sO΄��V�g(��}��W/(\�OR�EFBۑl�}���7������E�+k�lV��f���~֨s!m�H
�S�[@s.����>�9[}�������
�2��*KJ�K�"��G�D,�{�q�{�P�������䶮'_>Cj9s4��曢�܁��8�
�æ�Lf�ye�ֲ�OSޡ�-�/�z��j?/o ޤ�W��m�9c����,0K�$�c����-�E^�
%�b�ڎ�o�=5<����֘9.��o���NX��G�1Y�Y��ՙ�N��Uꕜ��9���Ϣ{(���5:�ڷpԽ�OZ�t:��yٺ�3.�ܵ&�SбU�.��̧��f�ܗ�{TM�n
���7�_��6�5���vU#�T��mQ�7�љPv���Oem�L+�m4�\�R�h4�5�吲�]�z�m�I�n��휨�P7�']�uCW\,�Ȕst�nw/b�ɾYn+�V�n!�O׶r����v5�ŭ�=ͽ���ia�a�.^Mū��U����<e��[���l��� �)�t�<�8��X|L��)�o�ВV�O��s��vwCn��76�^��m~���o~6�<��6�������>K���p9;6z����1�͖m��jLz�зyJSo�������`����pݢ�J�,�u%Z-��t���`�]��.�J�>�ꪯ����p��e����:+��|���kg��碽��v��}�7ztÛ�$�g���]D���Zֻ>|3�
�R���3�OjA�9��p��8K�ٓ`�OEi� -�����_s�;��EՁ�Y��?�Y!�q��1�\�Re���^ڏ��������	�u�r��&iҎ�R�R/}7�dJ�xpRi>��Kw $�A�;����=i�,�yyŦ�;g���5QBW�����־77���tnt�(�[�$��W�r�|�[����������k��u������<���^U�i�|���z�������/<ؤu5i�5��Gs[�p�QC�Wk��B�.�L#�6�>~����fx����.{W�nڗ��2�1����n#�hV>�Q��|�]�vn���36�~��m�ju���T�dm�A�24yk�$�[\z�a}W�Edo#Iu��lT���iU�fz���X�)U�m��0��b�b.�R��*�CX�$��pJk94�0l����请�e�f�+��1j32�n�ms��%�JYi�w#��1ly֖j9&�x�l%ʤ���_UDN��c�����D5Ck�לѬ�3*�*��Y���?���TM�(��Z-�[�6���?�$��.޶�{�f-�ʎ`��NϬ'�b���	x1�I�����
���M��[saD��O^o��~��9(>�*���|�)��m�-��M5]�GZ:p��(KC�����_ɧ����o{h���M�|yȳې�h	pw c��⮺¨��X���j��Op�>����;�Ŭo��r.�Hw�@"��?�+��I^*�[�JSˆ�Z�m�p=)M���|
���g��C����}rz�	'Q���<�mТ�Z�b�<37�P7N�{��ί��sQϘ��O��^��U��zAJ���O5�S������l楐�ਆ�"��ſP�ի�5[�z�'v��-��L�J�{��F>9MsW�����(������Z�[&�^2����ڼ��,矱w�B�-�6s+^��q�{����E�˚-m<��lq���#[��o������k�n�#9�]��GY�uա�48S�^�t�b��Լ|�Τ��4+�Q=��!{��4R�n�whԑ���8N�#K��ﾪ��,�[�}�zV׍���q���I�A�'�i�ö\k��lW��]�7�*��/���ǰx����a��âH�~[�5������� V�x��5]�7h9�Ke�ɸ�p��/$y��[Ug�^EV(�񜷞v���U��y����%n�y㱴�gU������1n�yp��*��l��%ΦK�"�f�>�3���3-J<q��Y7:���n���\��%�����K~�-��z�b��q�\�.�77�76��,���{W~,�ʢ��=W��d:���m��+�
[}p��o�{ `}��KaY:��bt%�F�`��A�[N��T%c]+بy��SM�������7͇,>�f�O��{��j񋈛P��Ʈ�e�kA)�����=f�]?�'���[���� 6`�0*�ԝ�����7+���>���{r#��w���Lu��u�C9`���Hܓ2�ۏR� <�'�Uϝ��˱@=;,�uʎw��i��t���>���������[ou�Ov>0���?�1$�ޘ��t��
l�V[NI�wo'K�����ꪠ����/v�
6��σ[p�=�|��%P(t�Ϥ�?�c�� ���*��g���9��V8����S�/�,kW�>͊�+�G\/���I�\��[�Orn�7^�����Y�v'��ZW���EC���x&������kip�~R��۽��S٩��s�V.8�I��?��-}�cU��c�ĎA/�]��\8u�y��|��R�V}<�ծN��_r�g�%�k"�m�k�g,gD��eƫ�B(��6w�~6�h�<��K@�'!ܪ
�],WM�Xd���F�`�6�]�ʚ^�y���趯�h��v���\���j�ʎ�������z9�.��xC�e;��Vn��Z�b�]l��|�����2�.Wp���&���'�dk��F㝛UsBoZ28k��mn s�U�NS3}3kn$�qڢb��eK�r֯�����}�aj�ֈ�dT#v,���otfp��{]OW����_���M�:|��:Ἳ4\��6믅(���q��}��Q�z�����1� �5#C�����t�uЁ(��Ӕ��vc7]�uټ�ŷe�\q�0���qY-��*�[��U}��x�&�&�������fQ럃�{'vJa\@��d�h54����9�'N{���V2!^��~���H<
�ި�tjuCQ�t\�rrO,֝��K�f�����Sm\:�������7 �G���v5��g{i
y*���λ�v����N�)�k/���I������H���s@��^��u���JJ�=t�*���o�ְ,&�٦����r)^�Nq=��r���ۈ�imZ�.��(�{�Z�c�_>F�`�H���r[�{k��}"�G��{��_u�������L������jo��^����[�e��#��R%%{V��5p�1�[h��h��s��r�jf����sLe��k"~�H��t���E�s=&`[��J�zW|^kY8�gn>櫉�^����m�w�\b�L�!��<�u�GC��X�Un_��ΜgL76jS��K�u�L�5����܇}uzo]�c�Ab�5M����Jiu�m�R�����x�o_j��+6�m�4Q&�"�)F�#�A��IG��z��j��'��[�V�웱�?}U�UWG�t���J�^�|��Z��>�>�M&&�]���"c���i��d�3�)�JK.�S�����D�{W����Z�I�է�6��8��8i�۬��hCht�-��_L��˟(�{W�n�{q��)��"wg���5�d��tcw�T����_9�U�73���ZjzW-���������
تj�9��Ds���3���s��{57�'�:5��;�޷�`�qW���l\K����L���j���������x�_"jF������ĕ�ư65�l\Ko�q]9�.ke��nR��ti��cđ���Lʉ�F�\5�ʋl+���\�{սA�������S�.YH�����<�vx���¨��X����k/��ç{ys�r�
y�bW�s�9WxTe���.�1��������o/d*l7B�*��2�M�5z��<[n����2T�h�ˮ�\����;+e�7�j���h��c��*Jzu-:��ʍeGK�*/�jf�=z�1V�h�F:�z��W
·N3a;!�xRpX�'�9Q���Ð���ﾋ1�BS���]����}ݘ$W���w�'�P�w�jjOx��{+m���X�Fכ�R����2���b��3�t���K▀
(��;��-{MvoŘ�<u�>�E���s�wB�J3�s��9uN��ni�i�3V�A��%���&��������x\��_L��ٔpQ��v��)�{�	��_�{�F����� �>��a�\k���V`�`�jQ�c:E��n�7B�KYV"��`�5��oQM)���@}τ��;�T��w����~��s������趬�Ȫ�Q�'⍷T��7�6撅����oV�7��v6�v�l�y�\�C2:J��8��f��>�P����v�7:�Dk��Y΍tj�SNoZ�*N�@�-�MGnӮN����kasaK���f��ͻ9G��d�b���y�R���U�!���H3�AP��������������}�7�Yi{9`ǔ$ʡ�Hy��3#�z+5�L77g-��_-1��DY�GZP^�`o�;Cge�6Iu��Ec_YZ��^iM.=B�t	<}v��Wnt�F~
�d{�ﾻg15*��S�.�sU=����_�LZi�����֫�vB�Nw-L�@Ł<�p՝����U�:�#iԝP�t�9����V�*Y�Wn���Yr��,q)����������*��j񋈛Sc����:1�N�{�JD�=���}:O���H���0T�Ԟ���gL�M�W�U˖w(�Ĺ[F�6���k^�]w�\6M����<� �3`�Z�2z^r��c�����p���9}�����gSb����P�}�ypVWOp�-�;�s��'5���̀��1>ۇ-+g5n|�h�ld���r!�3��;^[�v����]���G�j�c~��w��y�)v٩u.�b�3b�z���=���|ß�J�h&����Kj�\�>Cl�����w4�VfsW9�r���\kW�O!�
q�[�q���Φ-��z���f�Q�f�S��<�	�W+t���c��GdWkQP���Ć@�Pq@� [����=��L��=�h w�y��*w>U�Z���1�4�B!%;�a��׳����'v�l�D��K���h9b&�q�`,n��sZ���:S�����1����!�i�'��0�js
�;d�l=4��Q�%7�j�:��4%�F�7�$P���.�S�<�T����(fw��'r�	 �hx.)VA��N:�"��[] =�"�k��5И1�W9Ĳ����<¥�NWM�:.�����Msކ��$���O���	�XY	byۙt�#�b�reƅ��B�n�K�`SHS ש,�`��-�JڝM!.dk;r��n�d�tˌ���|A�������rr����}��h���W��X�w$[s�%������o�k%�:������8�{��W�z�>��I���*Ǔʃ�j������Ӣ���A�YLuh�f
?'�H+Oc{3����wTMo�lL��Wv��m�P�c��]�V�0�4�s }NvI��Z��:�l���"��G`ӭ�[Ohc����f��Cn@M`?W��~�J@��{b�_j�ѧ"��Vp��uE[$TWf����[K��������eJ�+jӏ���&[
��і�h�bo=��H��\��h;��(�,�Gr/�YKu���67H�M��"�RS����p<1^�_c)�|U`�:m�&�e���O�t����w����ޮme��#�/�rӗ��Yl��SqX�ܱ9���s�A�L�nl�x�vM�rW�q��V��U��n
J��]E��e�wWV%�VN������!�w��N���݆�ɹ+���{�d�{����ˈ6r{��6c����"��)Ig&�e��H��\���l"�:��� �72����k�*�0f�g���!��<E�	�D����6bٟ��4��.p��[�����)�#��!o=� gvHa��f��E��DG���\m�������;6
#N��	J*R7�rg�wR�/h���J^�|GD�Y�#6m���c���N7hj��(_;�lE���u4��,	1�>u��W�w\A����w5LFWi:�L���.,�ɽz�4��-�V��͖֍�pк.82�᝔M����<�;!��*g>PW"��QnT*��Ǽۊ���g��W���θ�t�I�*��7�h��kB�p��ls���6ifB�w�4q�%J�6�����mӛ���D��t54U�8<�u�
[��� OF1��`$>��w	�]����]"�����JT�V���R��� �'6q(=����Y}�����i;|R~��r���+ؖ,wM�� ��a����M��U��P����wI���x�����T.!2�d�Y.]�w-��,#*��v:��uˏ���{w���{�y�w����ן�>�4��p_�&��H���ar�2�I$Q31I#B�PPiy8y��A��wT�YI"T�	�!�

�NRAA�dʳ��^�5��*�P]�lT"i��9M2�*�*�YӈC�S�t�fV�+**#�<�j%EY2����*�
ID�\Ŗgs��2�*�X\l(N$,���8PEq�K*b�QD��F���4�$h��6�\���0�ɅIXev�"�;������顑�t���WRM.q"�f.��u'(���2*�ΓDˊ�!"���'��9�G:IZ��TT��˅0���L��y���(J�`��*$Ȣ,���{��BAfd+X���+�aYAF�Ͽ�����׋�%��t�M���r�v!�k/���x4wsȗ!n�;�,�G	�v��%.L�Y�r%��-CǷe��K?�W�}G�R]����:k77�ɪ5��q��T��Ș�:`Zڀ�n�ʍ��Y�w���Q=��RN�3^�>�W���p�(�r6�w3��� ���z��v�]$ʪ��kd���F�ju�m�����]�˘y[��pk��T��`�}ޠ�Y3s;��qڢ~�i�]��7�H�fn���d�>r��t�>�?Y;Bv_��gUĔ±�&-4�}��
nw��٣��3���7���w�M�\��e�蝕V�r'T4:#�-�35}n��قb��b���)��vmþ��l�DRG;�uLq���3��Իl^��2��௔󁭊x�m>�t�Y���l��6����y�ќ��vt��u�R����|��=M<�4�w�-�I=�Vx[h�=�t$�mRޚR�\5�v>�&��[�b{�Z�=W�[Oү<����ٹ�=�̀#n$uMJ��f�B�]m`�CRw4�m�{�qo;u�\}r�a�+X�`����J���c>�΂�յ���}�n%��5Ձ֒��k�6���kx�d��6͘��w||r�xv!ן��;[�g��T�+�J�3^��"�Â�G7ub��u
��r�ȯj�~��l�1���N�<E��
,����Е�ƌպ��P�ɇ(��GLB�������j�p
_k�,A��m-�z0�e�jl^���dLG
�#����`<ڗ���z�5����Uc��5��OxeC\�6�;�O��PЙ Ϝ���l��Vf��h8����%�g}X}�B���y�^��I��k �0���fL6S��5W�^�m�窯�o��m �㲨�-�:�i:��N�m�r�X�4�N1]��Rԧ2�QX���fu}2�/���gѼ��j�E�]��,��kfŔ��s�r�Xڇs?k�u�b"���U���V�u5=�vf�j�[�:q�B4u�9z_��W�mG���#u�fTAw#تf���=�v�`Z�uS�+Z��%
p9���s`�X�[�{�n�W1�n�,�y�E/Tyt󝭭�¡�5�o}�w�ώ�S5�*��z��E�G�W^	cx�G��3O1Hz�v�C��U�ج�;��$]������l��'Ν��=��c�<�坧� �⛂�T�0���5Ƒ���
��3[�m_t�/���I�a�OM��ϢuW_�z��F�5͋�m����]��s*��1`Cv��)M�֪¡��N�e��	^�J�cb���O�_=0����d�3]��,�]5=nYUH��t�{�D�J9�硬*b����LNfd˻�c1����V�罢w��aP~�l��Hn[�1�%�=3W�1=jM)����yOE�)D����U&+�),"�q�(#'9�\�{�-��mk��/��}�����r��:~_wIcB�|J�Hi�M>���u���5�;��ݷ
ZV�jY�;�����f8�a�0)�o���*Wyj4ޗ<���F>8�4�e�l[�Glؽ��'�e.׷8�-��!���mɵ��q-�ԝ|�I�i0�92����f�X�#�W�E)����YV"�o�#��oU֩���yWl�&K6����.��F�+���J*�Pa��&WQ��#�Y�%q����y�)��)�;�9����6�J��(�6dp�ܣz�a�Ĭ��>�v�d�ڎ�)ɚU�5�Sn�Ѽ�i�܏u%6̾���۴�ēJ�ӲZ�7KT�# B�o9O���X;Ӻ3<\n�e��eLk�'�赹2���iv(���;����O��RD(�-���o�NW�k�j�x��[�1m�R�	Ӛ��1즺+�ܦ�\f�Q{I��Kǟ7:�k�՗��;7Z�b�Q<�ajz�n��K�J{�~�I[˪G�6�e*Ɲ�W6���u�{��E ��D���s��7Ɩ�n~����V�IPՌqi�z>�͂��|j{��{O�'n$���齳��x.�*�j�����t�6)omh�c{f)ċ\�JY7�-�&��|�����ʊ@l�r#��<B�o�Ll�ow;Wq�U����=O���a�U�FQ���u�M9u~�]�p��aZ�Pu��|��>m���_�m�\�1�����M����W[�9ݨ(p/t��r��r��/�,iO��z��-����e�^�l�Юv�ks?
7R8$�`���!DT1�G/*w�fi|+ >���L!��()�9���:�-��Z�`�C��Y�a��^�B��c{k�9����w�q\��H�%{-j��\�_���վ)yN!tܼy;:V��~fL
z(o5�ub}��3��!����a5�[�@�0��f�[���P��E{5:��@X�q���{q4Y���u	��Q�R��S���Q«��	/��s|�I���<��M뿳�]�����w�B�$[�����.5�,�Q5���@�kv��̃�y�[TVg8����\��SMmy�z5'��`�n5�ʝvD�"��9f-!CW_�g�cq�DGՋ�i^>Y�?N<NW�9N�qY��uC*�,�"�����LY�$8�q��-�w�yq�^��i^���5�θ�-�����7X�eA�#1ovJѷ�'�Ɲ�/ד%��]=��b�V�k5Y�����!w�\>Y�[rS
�8�l��zS����Fg��Đ.�o�-�������tNϬ'����wӞ]�$#�qM�[���0�MfBw��]F�k�8�M�ŀR&��;>�?F�d����D����1���5I+7��<´���l`��]ʨ�q���Ɨ���67��Ke�P��7��F��j�@	�E�֮ĭ�`�ĩ��!��8&�d�W�OT��[�&�7bV}m���ֹ��m�=x�k(ܠ0k��if�9t�q��5MnJ}=X������[�5���yk5��m�JP��"�,��x�q��7�d:x������#/�\����[���M=0�Q�����<�jx����t�pbs:]��.�[Ҋw�ֵ�v5Sj�{*w��+���V���}P(t����Z+O5��[Չ�<��z�ۘ�8�'1p���iW�[f佁�h:o.X�6�~��8^�r���(�8�5���OI�q��i/��o�\gʑ�#�@���E,�{q{)�N�MF6Ӗ�����=�y;;^��m�l[�d"��CrٽQ78d�3�y��Fz��P�=��a�oR�l~��4�`�&�]�����e*1m壘�����u��γ+��+�~�ޜ����#-�MP���x������-=#���`���<Y8���\(v8�o�Xy5��*��mK��gJw��Q�O.��=�Kh#�^ʵݭ�����O���E��-����av�B+�)�pgK��M�ܱa+2yZ���ᛥmtZ(Vv��Nwmiib�Ԡ��K��SV����݊h�.:�趬��fx��mdo=��btQ���d�c5�1R��Z��*��tn5ٺ�2/�|3L���DV���s���XךJy�@竖�p�x���\�g����7_s�]��/���HĻgn͈ͧ�nS���%��+|�͋�o[Y�y���}�f #(=B��%�����*	�=�+�n"K��5X[�6ozvm¾�I7�[�Z��v�	r��X;���UN�5:�+��X��<bi�l��e
5��l�A�l9~7ʷl�p_Q�TF�q���
R�sy��uF�|���5�1k�N^t������P��IPc��F�Q����E��+�&o>mx�v���Ba������e)J$u�Ϥ��I��7
`�!�����)���%[�u��T�i��ې�Ψ���9Fx���s5Q}�a�<T�^�MF����ܭzAZ��ʛ�l>��]b�s���G>��y�f𭋢�+՗]ob�A!QE�����}-	&�ՙ�>۽�5
u̼���е��s�!����9ط��T��A�gEۻ��l�E�Q��!���)���+@:�h$�Y��j�8?���Q�� ,��ݷ
ZV�jLe���LB�H���C��5wr�^�
Pw#@�w�c	��|r��j�|��-����1u侀u�|�T7:bu����CnM�us�m_ړ�|������_�YOMe�C�[0+�-�t_��Oh�r�\]~��$��I4�y2����wv�+&O_f�qm�-�ƮTF�"b9��khe�D��cdV�ى�Og{�yn{�9Z�Y轫��'[x�2��v6��)�L�:��Q��.�*q}���7����2�.Wp���/i;*^<nu��m���ʧ������S�W��\;���'�aS-LΩ���<��ݪ+|W6.]��n�X��m�X.�8Ό��н���Bc2�.����!C\1��i�nW6���u3����YZ-*y�R���P{z����k�O岤��s4��XY�N��h���K�s[���C��6R�y�6�z�n�����ʑ�;Zݤ��;��\�n;L-���.�̭M��C�k-����*�mJ�qZB��W	nˬ��%��[�Дt����Ij-+k����
p^w-y|ggD��́X���"^m�i�V�y\K�·>���<��Q���X�T���=�j���q�
��S�n��������N�������C��r׷��.��C�9]���e�8�=������{o�q��P힮����;B�哺��.�Z���֖խ�w-�e��Z�ey�{�_iUΡ�׼�q�9�'�mO}�%�R��_|ub}��p�j�HU���wW�nq������'�3���Z��oأ�7ߌ`��b�;�&�ݐv�2�W�dL*F~���+���ȷ ��rV�	�M��ڮ'e��2�>f�|�.5��*Q3�����Ij����쮧]���Pu*r��^��������4ۍw*b5��u'Xć�׽8�O.�S��ŭ��us��ׯ���u���*�������������+����ˊ�Q�̡��g8��XlU��5���1#^j?]�{}�M[�{:�h\_w�ޜQ9�WnŹQ�(����הއi7C���t�ё�|�l�4��q7�i�ޞA��-����D�Ǽ|ONjZ,&Ix5�Js9�_L(�l���k�%�#���0-�@�u2�."yp��N�j��Խ�OZ�_�j�	r����p�v���=Mp�.�߃�d���.����YZ}=~�O�Z\/��Wg���/a��l��u�{�1n��r�U�ʢ{+n$��j�d�n��yn�=�Ê��K��E�
t��\K�;,'9��7ܯ�j�����.R��k�Q���7��j��+���h'e�62���+]yG��i{l�1�OJ'X{�+������m=_:O��ZX�t�r���N�k{q�R;<8+�������¨������j��C�Sn�_^>�
nLlby��|����#��Ғ���u������g0N�ܱ/��U��RcE�f8hgT>����y��.Ejߧ?��y�q�\�q�y�ݯ�p��u;gnC}��l��o}*EC�ѓG��(��s�q7�9z�xoZXӧ�~O	=L�����Ui�����W�e�>�`��%B��ƶ�����Й�BA�No�"���;k�v%;�A�p�CE_<��CV�v;��!8�"6M!��V�ָ���t��]�Ӝ��k�6�s�^G"yՔC�����ƇW�+/�)z�#:M��w�OsA�&�f�b
׮��Y���P�n��6�>�5�{�n�$���`V���.g{�i��̻�K:5� ������	��
�]�f6�N0J�U�%�;�ZF-CK� Y����g^o˘��u0�k����u5(��w�>5�(4
N5qU��>]�}���mG�dSN�����3�r�v��t���oU4�s�d���S��/gh�A����v���k�ZM� ]\M��o&ʙ�-+��4^샋<a�}S��i9Sp{毷JW;6�B�W���_-}�w&U�e�����޷B��)�a��o�yxK�&�J�KD'yVp��ǁ�-�b��}��|����4���#�B���P%X���*���x�|Sc�2���w��ҭp�7��=sƺ/nsu���;SD4(��7Q�R\�2p�"�vX& �;f�=^��� ����3�.݋�~�仩9j厄�YI�J��Y݋�^m��<�0�wn�_�-�MN��N��!�	j��@r���x�개��,��4�{Oŧ�&.gZ\�b��<
��8]��S)�J��P���hN�s3����k������د�V���q;��C�_Y��N-��g9�	��P�O_��9�t2���_u��]���e�9O�����i�6��m��ǫ��h�)Ҥ���$�oy����
!Z��NvC�/xŌMNmDws!׻�3�[<2�����Po>ɤә��;�/h���Mn�1f_-�t���5HS�-�q��F�rso�E�vy%��u�;��N|e�!��c��wD��G�.���Ǽ#���}c�n�^]������p�h~�ݞ/��̰"���xVsT�r�����sz���I�"O��{Ɓ]3F���kO�9���+��W�����5=�������y�&!V��u��j�W4��Sw��S����+rq��գw���O����|�U_4�9Ri��<t�:��l��]��kkGZT�6�2KҟQ�Yp1(ƯO��5����D�UrZ����vnCwx���u5����4�T�-�ډwvV[���t���y^�u�;aC\�5�,,�df*�|�Ԛof+;vӤ����rM�*�r� ]���X�})C�I�F����-���\��y}�c`�q��j^��X�ki$�U.e������ȹk����y�{A�2q�C�WNm�/]��l�{6�5)0Neh��	��mV��M�\���I�}�]���Lan3�\����� 2d��/ �Ԅ-P�4"�*�eF�I�A���܎\r�2����V�)3V�������92���\�"�q�vNwt�"�q�Zt����'BiP���Qʍ��L�3"#Ju�P����t�B(�Մf�QY��aQI���Р�̒.Ңs�%����Q\L�+�B������
�-E�jӅ+Xmij�c���eZ�8V�$At���u���d;��Uf��P�j۝�Ls���t���s��!��8FIӚJ�5,�nI®GZ�����	3�tj ��E��D�!B�"9ܜ�����r����ND�������K9AA�s�eQ[B.S����	�I�V'r]"��e�uK)�^xh��A
d�YʒK�jӖ�(�:�.��L��V�I�N���9�Ԫ�®�Urb^��d�)��	������N!:�V��^+���aKN>��3Օ��T���o���tFk㿜��2�ד��7����<|obi[9��3�*ȟ�#�s��T�
����m�b��A��ʹ|�rN���k��m�w��A�J'���9t�q&�v�^�M���	���$���z�H�?_���4�`�n5ށ�WfPѭ��Y���5Dj���v1v���{W����Z���+9>���1�*��)��KS�=���ج����[P38���˚��{aR���;I�\�P���-����c��󹘍vn��Πf*�f�1��蒬fm$�p�P眝^�al���W�o�2;��1w��w>&x������{���2��N��1�Ɯq\���yw��Y]����_�Uo4��9��j�)gn~�WWӮ��K���V�5͂��;yXjA���Q�Ѩk�)��{��~����j�-�%���X��<b�-�\�7��.Qnc{f.�8R�4$h3�
���vj�6�W*������Q�p���Sw�E޸�Pc���=���Mnb8��"��U�vu��ӕ!t�+��M�];'-���`��k,�� �ܓ��F+B8�tM)1e�y���u*���I:�@{��[<���<�����g���j�3ʁ�֮>��#�H�DR�r�xެ��"
�����{I����;��WϔZ�$��R�<}�JFO&�QX��UbL�9oc��žJR�:~����I���_i��t����{�	�s�9�^����gn63�.Q�:ڣ�K�BU�٣՛W�^9���Oc����������L���x'����,����δ;��G*��_�M��簛_c��5p���gOs�Q�&rz�f�'7�5���1<��<������q-�R{|��7Z�w{\��J?A0�b\����N���Cd��[��N�-i��5���𦏲sI'����E���I�ۍw����1��/�6,. L����%��D�S���[�^��Ns�8ec���g�Vn�1�d�}s`XX.�ymz���2Y�u���<n�)=@�6����z�t/�j�/+S����5���Ĺ�=�����`uz6W��9��@]�����Nv2z��
)�2\�Rsv��r��1����u�Tէ+i_V�:���̸)����M�)��7%t~����8�N�S���nu���C�2�otM(�$�kQ���9��zY;�N������_j����esb��oiҁT����$�qo�_���t�>_���Nϯ�q,*���L�e�*�k��"�5F<s؍���>���.Z	���uZ��ہJH�!�*����CJw���m�%[�<��}�E��Y�v���)�y�<�O7*�jk���39���:�Ht�ұ���ݧ����>��oD��7�9U����K����-�nԭj��TKti�{q�Z�<��l�FUM]R&�RM�b����`�����[X�|Y{o䵮|/uUỖ@�]OE��nSwX-�]�}�������`YՉ��Қ܍Tع�+���-��1x�����H�h4{ڝR��ܪ&ϕ�x%kV�Ug�REj��@��f��qeax�ܶ�`�����ilQyJ�SC��ȣ%�n�kl�}�V����\z�è�*���W�w]��#���r�\���^~�ih{�GLІ�Qrc1�񳹖@ka;�w�r̝6�j�urr�����n���S�#�Gk��>�VL;�ۜ�a$Ӎ�M�����+�k"U#?S��R���{H�� ��K٧ɋŔ���P���\�o�L��p�Х?r ���r����%8;kh�y]�m}�������4ۍj�>�d�5����O_=6��N�C�T�n�|�Fk���Z��N��8e\c����&gf�+�k����]F�k"�T�Q��{v���Y�^�䰒K�j��x��-F��խ��n>�f���󑘫�{q%hۈ�_sk0�%�-�j̮�q���X3�ө�J�Eew�s��D���d��*z7�~���:%p���3r��r����͘�����fX�p��|��cT�#��^�k�Q+�+�`l5�d�������^��r��x�1f��y��j����)�(��
��p5�OX�z��|���=� �L˛w��S�81�,�bY�_Gls0W��m=�&+쌯+��ȼ�[1�25Ƅ�7nM|�*bX��,�&���0sd֖�-Vⱷot╤�c��w*�bb
�4��p=�/�u�*�(��S.������\{e^ل�l�G�\5��vg ��L}�쪈������T��w]aTJTW7��Y��h<��kn��9���������5B�s�
���f�4��mQ-颞�v*r��ǫR�JA�Y����P�Z+�P���*�-y�w�������>��)OTV7;��g���7�+��K�g��	dn��K�g6ER�O�ȩ��]�~��^&����ړ�[9���5��(�q���ά�6�泻Ԫ��hpi�W<��$�=�s-�3�;���;�]1��ns�-��\;0��0mk��Kj�Rڈ\ï��/�x^Q�6\���n� 0Z�k��4��Ƃ�-�Ѿ���@Ƒ�S�J�u�V��WA�m0k�6%�	=.#u�4��qQ�9�kjgT�̸�\�)ǆz[�]�[2�wSZ`�ڷBr��8e^;Q�c]����|�1_m���C̩S�����[YS�o�lX���Ra��{�-LݳS2�D�}�3c���(��*�z�Jg�������Vlƒ�n�Tx�����p����{�r�͹dsU�P7�n�|~��&{Q�u��k��"v���2�}�Y�n��3方ko�=�]QOr��.�m�WΆ�G�&;��s�uh���|u�v9c���������=��W�1D�Ɯ_�sb��om��vl���Vv�d���K��M�̢�`gT�
(�al5ͅ-�H�}Ž�'F�������%\z���	�;c�Z�Z�R\it��L�E[e:�"o���ᰮ�����l��ݶz���N`U���s���{c�^u7����=]Ă�����D=jOnoP��� :~+���iw��F^=i�/��%k�A�{N��m�j-�ʅ)P������������җr�v�;�p;41�Z�ޗ����b�g|�Ψl\������7^K�]�����?�$�	豩����wgB����jX��=WR_9j�'/nd�N�g�<g�}_	J��Ϧ�ys܀��|r��W�הX�-4�t�z%�w�s2K�<�|t;�n���1�7-��b>�
�w��ڢd5��vTb�n(:-K�mw��N
m�{�^��s��kkP���=�\�(q��CWoVk��R�[iM��)�e�uX&����R|ɉe+Yw��j+j�����u�^ՆE���Y�	9{e�>W�1�mM0�q��XS�'��n�kQ��N�)�׏n�؉�ɘ�w�5Q�r�5|�����啮��;�Zնm�&ᚴ�Rהz㭋��]��CI�r�jOj��xN>�[������)�4"�پM���l'7C1�ͬ��\:��N�������>nu��t9UP<��E��0[^�����;L�v��Y0�k1��+}sc�>V��\N3{x]v��v��9�&�[�$^f_j�y�`����į{I�QrN򽎳��Ko�Wf�+����U �*�V˙s	��&�.�D��͕�;�Q*5Jp1����4���\��+����9���m�H�{�_.���+�yE�����#[���oS�t�	��8䌌|jbs+��=q�qJ���u��\��>�5uco48h��F�'�S��4܎=�}k`�X���Ξ���!��P�jZ5�<V�j�����Y�h�^m[$l�(f]�G��96����Ir3�{�D���;}�-�籯N�P�=$aUbk��Y�*U %����gZv�2���=���ztE�ZnG����ˮs�1A/�������Kk�|Y}z���g�m�J��:�j��4:֊q�����t�`%�����`Y��l��Y��"J�u����r�9�r���,�ʣ�	H�~��f��\�1�y�!�f�3�ww*�5.34�m%����R�G ��h�i�?��gS�����J�K�kN�!�˙�����.5��!Mrj[���q���o+��O��&�m\D�=�K;��]�j����q�\�0/R�.gws)��o��w�m\�n&�V(��TW���N��j�3��ۗUN�ULMĂ����s�pkw3���s/�ڲ`<V��í<�����em�]��2/Sqz��ޞ�~�n����!�%~���i����M���3�o���mY�K�;8On0=�{q�p�'WދI��(�
�[7�#���[Z�ݹb��1x�[-��y��.��dU���~�Rr��qe����dF$ػ���k7ud�j��;Y)����\��^�f�ӌ.΅��q�@W�J~��x�ʮ�ͺ���.��e�譙��<[9�kg�tU�9-�qL,i���͂���K{�v��J�`v��2��]o;�RuJ�5:��k�Q���7��j�vk�]$U�5Ҭe�ע�R��b\�jxe�UD�Q:���tl<[|�lK�jj�ʋl�
����5q[3�۶y������>��#�#.���Q����C�h*�s��X�u��y��M=��MP���0:J�;��)+[E���M��pGn�^hp+�S�Ѿ���r�tH�_>���K@��#�	�'�^�����>5_u��>����P��r���$w���؛���;�����08��E@i����1q�I���j�d)E�!w��Ә��o	Ps\��K1|ox^��3M�����K�Wv9�b���S�*��y�J�n�pk=�uM��2���m���D��֏��sŰN�'
5D�������ԅ����E_ӣ�?���!�%r�q�u�ZF����H��\�%��кv�w �p��Lf`�@rT�#�β�0F
��Y$��r��2H[�yq+|5�c���kڽKW0��*��׉C�j]h�u����x���K�-�F���m������5�w���Ng7��y�Xd������7�P�����Y45��9��'� �|n>;�
�{��T��-{�*��r��/ɜgQz}�y~��W��k��s��=qˡ]��9���~9(zf�l���Q����?җ�k����201���w�s^��;�Ox���=�&��?��>�n�<�tc�t^~태��ś�φPs�L�QѱR��9e���� /�Lsl��w�vB��*�����/��#�,��x�'v��e} �.+�U��5k���}^_�����[;�Y�����-3އu�r*��ʝ7e��pf�=LOL�N�\���:��N*^��n�ӽ���~!`;��K�o�c��v5�Y�'��}�����.*#���)d�Z޾�G`6���>���ޯi�t���=�ߝxvM�p��`�;%�+埼;����W�ܹ��d�첝Ӗ���;V,��	��V��L�L��Ix��O\�+���n��+�'^Ż'g��>���&�W��2�_H��GA�bgqs�Jg燣T÷@��%�Q�`厇��(�D�d��Ltb]j+�s]Z�U.Y��|C��&p'�GRէ���\�v�Y�uv��VM�x�_>\�G�A���W��(ރ4�n[#7H{<4s�̚��>Ժ�i��z�t2��!1�긜�r�S�]��p�������'�R�w����|�FŪ�����EE�:���%7]��q�o�ǺC��C�N(�p>Yy_
Z�;�/$���B��vz�V�?y�D��Ȗ����\��h���:�cc!}��\�x �w���5%tP��znNte��egN����Z�J:m�FYBB
�G�#V]�:����|^ѝ�dJu� �Nn�گ��X���|a����$��ygGS���c7cR�9��vr%!�]lGzqb��ӞU��P{8�y,�K����V+,��;,<&iW�������OR�1��LV)|��;��A��]�a�� �5ؕM�p����z�Fv�W)IP�lu�1f��4╈!J�}�Z\�f��ڦ���5�9��}�S�wGoQ<�D�"VG�
*���r��l�b��=�iø{�T8�C�L�Â��	���4�GN�����L�V!��,F�7�vi������������Er�7xX��U��c�����w���9��wA�upAS�"��XI����*�
+��U!���UoA� ��T�,cq-�9��ad�h#ԨG�3���+�nc"O��<�8�V���,hX^ŧ<y�a�2�F� h�=�z���ie
�$|�@k������"�����$�����쬽Y
�������j��r��G���JP���a� �Q��F;�.��>8�'�Y����#L�����u������S/,�A���&��D�q�s~T*�h�ȴ����y�z�Ӈ�G��*ޣ����&�xo�� �&���m�=��X4<j\�;���TGB�jΥ7�t�h��~����n�J�$��n��{���V/�����j�AkdSu�bʐfwKI�F>Vc@�۲0�Q7�t�&�5�Һ��*��
P�:A�@бj��[�&1&��,r�K��+p�f���߰��q�̲m��B����5��t(���t1��D��FU�!tbT�e����ٹ)�f�e��"99*u-ŀ�7�|&��0w�̭�Ku-:�O5��6��z���ڣ��U�������,�y���#ݸ��������>C�>�����p��ޫ�7r�O �z�ks��n�MJ���f�gD���`{D뒗�a����fm�ff	]X�y�v�a]j�.�F�t��%�/c=�m�z�u��(����{��2��D��:ܒS݉�MR�y,u�w,�s�K--�2nA�L�s��.�t�̙j�%b���@�㜰�Ք�)��J�%R�v��b��s+)f�d�)$���$�"�A�9��d�C�'��
r!-+T��J�Ei8'%B���f�Q\�J��L�3�P�*�9
�YsYd%G3��`;���i��l�TQi��h�n��vU\�)P��βL8UrT�*���uaxhmQT�T]Q��h��)�L�4s��{���EH���9��MQ	$աX��y�p�JOR����z�U\NhD��	��*]0�s'9�QjY��L(s�̜�$�M-Nr�[,�K ���z�"<�z�ykN�we7'w�Mm#�r�룅蘕�RUqZ4��r4(�09f�D�z��.h&�pF.�lǛ�'��g��y��Z)�n3v��(i��4t�������,�N�\�B*җa5�
0����n�>k���[I	�K5Vj��C����#�o����^�\M�w�9�'��Ͻ�|{<����.��lW�(�a��F_:��h��&�9FUG�}��	��L�3�3]�"�҅/W�#��Z�����Prw��FYħ'��𽇒���L�zd��������Iyי�gZա�>u�lx�Sf~۸�B��X�6��g����O����U�(��T�w'���W�Q�Z>�s���W#Eϣ����1^��{��tA�X�ޟS%�xΏ9:çrB�OT!x�ʃ���ggnpF�uz �N��{��K��B���B��~Uro�7^�5�{!։~��Qd�ߌ��qӂ���w��=�ڼ{�\�r���K��=�iM{�=���M���>���{v+��d�)�(������ɓ�d��*���t�W�|xesW�w����^\,�o�|c5�+�^o���ǫ(��}������W���:XD��i��f�p/�:D��z���u���^��؏z��^����>3X�W����t+���}��<a�������f��/ꬫӕ*�b�`
���u�~:k֩_�)ޡ��;�޾����4x��+rs�h�C�
Q��3��<���"v%�y)%��	��yb�YSr�\�/�R�GNG2��g�����Pqd!Wk��{�%�*c�o>+��1�:��Tޗ�����>�Zܶ��c*O�s�]�g�c��4����֘-c���;�uA�ꡕ�6���ػ�1R�44�u"A�������r�0} ^r�H���zNW������V��y\*3�����Is��0��2h�ί���-��)>�r�{�z�o�įl�uz����~&�}�$�rI����M�Z��u�c�851���T�|3�UG��� w��}�����/�g��yg�o���'�*�w��=�V��|��� �`L�X��n�3�wG���>N�4/������I��=Q�꾺۬����Ȭ�=��fхJ9
U��)zd-�_>���zБq������ur�FkZw�{�t����K�Z.J,	�c���l����j5�%LW���������i'=c�us��ӵ���ԇ[�W�>�}_��K�X
|��d�}7@�����yvo�3�1��#|�F�~�Ϗ�����x���3_)d�T�ʹ`�Lܫ6���'�z"r��^Ez�=g#���&*6�5~�{��O������̅���'ν��D����8F=�7��Xw3V�r�*J�d��z�V'�_���pUn�Ȱq�Z�)��=��Ǵ��2_k�N�L�R�6�.M�:f��k��`�kokp���e��䇜�V�[^�LO1Y�z�-IF/&V]�wպ�	N!	��z|fp+�t��s���Ȋ�O��:|n�\{�ܘ���fO�}|�T��>���,Ns�G�/�_qD��0���˯���oz�:���1����3��^�� 7&�w1�k��g}�TzlH�yS�C'��Ɇ���a�W�t�ԝ Vo[_c�U껭}�ݾ�P���`���"7ޮ�{ޫܚ�2/K'3��/�0��/�MߌV�N3��x�p{�>�J>��������zgޘ֧��Z;#��g�ɴX8p�d�^���\
��;�^%r�ը��Rw|r�S%����=�Iȣ�,��>�����r�[�8ܝ�7Jb�}�w���+<Y�D��XY�uz�b��<� ��q���oΗ����}��֮7� ���;s�w��1��3��ya�G�T�$�(z����uW��W:,���Vw�����z��~/h��{���{Ff[8�I�?���\6g���P�KI�b9%'ʘ���S�ȵ��wBFo�d��,�i�~��Ύ��rԃ~C��+�r=�G�������C�%GĔ8)���˿ý����L�<�g�˄��b���E��-�ZBP�A����+l��H{B�0���@X����!�T�\�[���l.�A<;	��!�JO6c��6��%�Z䦒��{uJ��3�u��IG�U���x�^N`�7��� ���,�'e�F��cM��F8�>��\M��~ӑ���V�Q��IP�V�4��K L{��޻�b��S���� �(���|=Q��F�+��W�#�s�iQ�*�o�����M34�AFw��~��O.n��+��l�W�F��}�#��7��o�ه�޿x�ޙ�&�<�@��W�{�����FG�2S�&<�Q7��62):|{`9c��VF�y�����������y��z�Mei�ۛ��=�Tl�3&��=Bf��0q�z�}Z��rƾ�ǌ/G�S���]䃜�
�w:�����'z ��ԃP���2a����j���K��o4$^�`U1��g{u��5��P��ח�<�WG�O�L>Y4*#^T������	mJ��U���?�1Gz��=?7ͨ����9l��G�^u��dy�{�k�������}S>%ɯ[�,6.��q���Nz�{��z������V_�Ϫg�O����:�ǳ�s^��>���z�~��s�n����Ǜ�3s����3�Fp�=�t�</ 9�몬��*Ux�ò��{� dK^�����
�xG�;���WS������S���Gu�t�͗���s����R_?�����C�w���	���Q�^���g��Մ;n��8m�c�|���4^�-J[b�q
�bz�C%�EQ��ɷr�o5����+;V{���}#�`�5F�.J'jD�/=���ŕ:n�;��2��(]w���T��"׃��>�+�n���M̼q��;��3ҙ�C�Cx��Q_FvT�,�+3�b몽&���rw�-S�;r���f�[���#=���"��|��?SY^�<8����R��e�x��_�UW�1tȁq^�[�ђ��2���+�,��~���z��=�|^���#�_��j�n�+�H�J��pw�`eo��맑���lU�[�^,f���>�TO:w�9�'��Ͻ�|{<���4���ٙ�4��h�����<���AmA�$�W����e��]�#��HU��i�N��x�=�i],���Yp�<w'|���sުfB$�� $=$8��I��^gv�
�֭��ؚ�~3�8T�Q���ᘚ����i6�A�N�D�J>�0�&�R�(�}��{9eS�{��y��Zp��=����҉���tx���7�t�@E�� �^#�c"q��ȫ~9ʳި˭�^=sX���Y���}��x[�q����#Ƽ �d:�1�R)d�̺L�nH*Qaq��>Z�xmF,}��̱��[��R�k��)8 2�uE��=��3^]N�:~�q^�:�RQ����8kS���wge�SKk���o�y�7$sw�����}��%����؎��c[q�X��Yk���9lʴ9.3)�q�~���R�ϼz�Gt�6׺��������+���yT68�&N�_���7�,�7^{�q���Gxl�W�u{���+�;��o�μ�Y�~����)��˃�Q��\���\1�k�uP{�9����p��|J��K
�l�wU�:2��J��c���<2]{s�9\����c#�c�y�:����3����[7��f�����N�b�w�>j?�����>�Ck�=ξ��׃�:հr�Y��{�cx�l��\ΝE������C��\o��Gk�&*�����;{�w���� �y��*r��3����Z;>y\+���;E��zK�F�rs�s:�J���=�G_��]�7N\�}�w7��T{ex����?�j�M�
]9'F]@Jz~��0�����k�L������S,e����4�w��s�'��r=��VG��y. 7r�+.����li� �|g�H-'��������U��'~<�����j��O�l��>�OB�^,�=����v.J5
Te� ��g��9��z}�BG�4VH�.>��|��8��ٷVӒД�JЭ��۞��;N႘-�K����]�u��ML˧�sK�R}O�鳳G$�*�WpX�R�^D�\���H���R��v���X��{c&�z�;§*�:J6� T먡Lv�A��زY�s�5��7��r�a2�f8̱ߝ�vy���*�ꃆ�=N�\��C"@������W�ƣf+��H�"�ԅ,V�����}Gѻ޾��3ӵ����RO�H�O�%B�*]� ��H�pc.R�1��;^��o�� �����>���oZ5p߭���� |sӵ�oδ
sl�,��ax���o�+E��$�m��N�=��
��^�J��Y�_��&*6�W�7�O�>>>�7��Z���L2�����W��8�=�%3!�=>3,+��D��c"�W��9z_{j��ܘ�o�d�K�M^G1֎��a�n�������ْq����˯���n7�î<��0��m��41�ۂO%����%o���s+��z�X(Tkʜ7��ꁓX��gոv):@�AF	H��ɋ�Y��ֻLh��μ���q������Q�ɡK�R2��d�٘^5v�ݖ���y�6ϰ㵋k��V�#}�x�{�{�^
]W��>���K���vv�
��䜿��t���z�D�?yge�,
}L��j�]{n��L��|v}��ߤ��J�>�����rS�f>Y��{�k3	?bsVdQs��~�&f�Z_��cS�{n:�\��p��� p�r���I�V�@�O�%��]�f3� ������>�Y����U�or0z�����E/���0ޠ�e��0����xd7�:�[�̥vԦ�9��X�\`��:o�,��~�6?U^��^P&xzz]L��s��8{����>s�/M2�[�Ǫ�*�]�d��P��O�����4�;�� �����[��"�ȳѯ�a��W�fC�z�O��0���O��^�~�*~+��=����R��e��e�&�1u�J}9k*���\}�=GwWwZ�v��A�=�n�y�s�$=�?[�~�w�(��J�0�L��g7P��ŏv�s�|�VK=�u�O��{�q6�ߴ��}^eo����RFTC�a@�� yN申Gd��6n�1{P��+k����W�����tǔG�֑�����>�N��I���2v�y����u���@�p;O��'�~��t�|7C�F�֍F�C~��dzw��>'@���=�e7��������/�<��@�}��W6�DO*Zq=�#m�nL~�j~}�"�����>�&x����錁���ɤY=Bf��0q�z�}Z�񼏹�QH>m�ͭ�M-{nօ�O���w"ߝx�����C� Oz�A���z�L>6}��_q^�^Q��D%U�[tJ���{6-�U�Ɵz���)�}mK�7��+�oj�x���:G`�� �Xl�m����!��R�_�-J�2ӵ�����J}$���eR��\���qF��E`	��*��M�l�����*��=�r�˓w�oTN�V�&t�1��<~�N���N�c�]~�=+޿�Y����d�����KMgu�7�x/,]\�fz7�ER��,�����g^_�G�W����@z\�F�*z�Fw�$�x�g[U�o���ص��}�����ѧG��-�$�'O}���g[��f}��TG�=��!z�yA�s⽕��Α��?~\G����t��2�Tӡ�UVYѕ*�9e���� /�L������Whο<����#��l�m����w���.��i���g�8eK�<�׃��f�>�����\���K�g��֭�>�x���!�r!⨬��qe������1q]U�=��*�]��_�{i��W���U~�Y��w��)�!�'+�|�*Q��<H~4�lH��U�}ս܇_��3�{�~˂��7w>��9���=�G��9��S��@fZ��i�L=L�`]^�>�r��@��L����wG��+�뉸t��r>�>;
���j�dWW��c'%��g�r]�fGe�z|��D`�P���>�n�����u�B��֑���qY0�vZ��we��\�����V�� np^�^���H3�kf�Nljd�7v�7Kjd!ۼa��{C\�t�+����O8aDƂ�%�)�q��Ɔ����k���O��eݭSU���kM���lWGxq�d�3��o�ː`�1��
�?�M�����]�#�0��@��wc�XΏ3��s�_�ա�9��l��f����f�A�X��z�����o�:��˘��d��S�	�bez��R��7��W��sE>ʔ���r����U��p��lx�Q>�8S���%ӹOl!x�ʊ�㍰���{�]{5wkPuyٖy�Gz���G������y��>�����C�L�p���f+wކÜ���W����g�T௧<���WJ��9�+��׺��ΪJ�~�=&��P�A�k�c�y��;ә�nǊ�>���F������뮧Ǆ�U�_)��:��d7�1���.��%��|'�{�.����srt+3g�Y.�d��l�s3�86):D��c״�<�9��o۬T_�S��ܮhy���}�{&���{*p�qd��wKU�zr*Ux��f(�S��۩n�[����~>^�>��ޏz�o���Y��B,�ۃ0���{]�Ґ�8(���]o�.���K�=쏆׀���#)����W����C�Z;!�p���$��g���Ֆ׌� wS4���<w��_skJ�w(v�5xk,:�r�R����^t@(.���U�;�5��s
+������V�e]�*
FD�R�r�k�&C�qr'�����f�ܗH����-�Ź���ׁG8\�E��LC�֌�W��¾�����5փ��tx����g��`�Q�<���+*�[�:%���3���d%�N��p5f����{��8����l�M*�TI��}m_}���Y��%���v�*(.�g|��F���Y�0�&S���t��%Z�E�w%�a��̒�GG�6l2��`]�_]<h�~�F�G����f#gQ�����8��-�FM���rF��:v�%�{nl_c/5�*jܮ�O�j���01-Z�M�k;����=��;r:V���j���ʎ�"��z��gWA�iW����=P��XA�S(Uޣ����uĬ�6E�}H�T���Tl	b���[�V�[�(�;�	)65V؃(-��m"�
���x4hEݛ�����q��v�dm5�zy���s�x&��-u��e�c�|�Ɲ�'�-�"�7��Cv�lᆣs:�u�j\��@�P���m�Y�i�7]�snٻ��ͭ[��]��b��wO���0��L���b��!NI�"���æ��E�hu"1�#�iǐ�Q�R��?�]�uTφ�.Z��}���b�����پr�y`ݿ���,�1$q�9���r�W�#�,~@)�Y��yw���c���/��w¢Kw�v1R�����e�L��]�"2U���!���J������[�\��kxPd���]��8f��)�4l��;e�u�&��Ц��� �[���ꋅ�bc�b���rO��$�.�0T�"�sQcY�龼��i�6�u"�_3�f#��i�.T�R$(���V�������5��og�RV�e��i+zw`C¡����"^�9c�o��?����^�\�DH���}��P��%��8�ڱݕ!ω�]�Rw��SR9u�D^S�"�t�O���0�>{����2E]@j��0����/������`����V���z^�Ĺe��1��n,�1d�6�3^[�G��M������ܳ]7GZ�E��i�nϜ�v��x<;���K*�IkD��$_�׎̺�����;�=���41$V?n��zU�x�̉�6ݟi[�����g-�����5������=h�eN
/��B���]_`��7���u�;V[�\���L�л���-M]ɠ�G�\�u�j���@n���1S��x!��*����S������o#�ح�2���%,sTw1s�)'&c,ʕԝkܲ�gA���#h�8�Ē(��!}���en����`��{�TnW��W[���,�����N�Ow�w��O���>z�|2,��qNp�W.���Z!uݤ���h�EI��u�sbI�s��Rey�.�r�܋� S,<㇣�C��I�E�@�\�c�)"*��r ��ܖE
��<��Ν��e��u����8�8���Q��ȣ���G�N��(稚�2�l)(䥕Y%sZ˹,�=wc��.��*�T�W"�b	G<���H��ʼ�6D�T�*.�H�\��	�XS���P�+��
�#��d�� ��U%{��
#t�]�Ύy�Vj���NNn��g��:l�6k�u��8绸�N�G���G9�U�]C�IĈ;S�H�x��ȯT�7M73��^N�E���rr"�n�F���;�U=J��r�Gv�E9�9WT���rtq�A���$�aQw3�`����z9�����.;p���	:r9����������׿=y�M����(����br�d����Y�F�:�E���7*m�.�Ҏ,��o���.���EJm�,�})O���.�KURv�}���]����G�W���P�W�����p�����A��M���Y���W����$�O��*��WUze��TY��:���ޯi��I����K�W�����b}�Ś�q�@g+��C�A�g�P(�/I�� y2����R|W��U��'~O�TED��Co���0��)>=g���i�}�_( y���R�ȸ=-�}S�ܣ|Y�x��F�f�W���v����W�>~��+|��^�����P�\�i�*3�bb%��g}|fkLqg,e&�ϟ^�K9������Z=>T��;\�{��I����z�iL�. �#s�\ātUvM�xk���j���z_���Y֌�s~�Ϗ�����x��sl������-Nr�i���K ��⤃}ԅ�R�3�r9��&*6�W�7�O�>>>�7�vuj��I�2��$m��'A�L����`k<����{��}Ο�����w&7}l�ǽgܐ�3<&�ԇ9�)x������նj8���%hɇ�'�X�]Z:���ޯ�#U?x�r�-�Cu7wY�ԅ��:�e��p�C�3�.Qk2t޻ʜ�I�2���;m�g���;���=��Fz���\ӽ��3c�%�z�?f���\��וF�Xl�:o��ݾgx��v �=�w��x�*��v��L%wM�#�;�^�Ⱦ�r�<�C�}���L����=X(k��9��O�L5p'tø��yh���Q]�}j�&�6��ݏ�����lxgUׇG�W����]���V
7�B�^ʑ���ݳ0�{C�������w�����3�2��9�@TE��3��ʏz���!~�V�5���À�Qmn�CՄF:8�[�Y�Dϰ��z��ڮ=���r}�zJ�+���EzsǼ�F�_�xp�KZ��{�v�J�qhܝ�G=,e	�
��3\�y�A�P�������oݞ��U�&��εr��L��w��u��z�����d0���>�ё8��q]��O��nW�VUP1�w�|9j2�D�����~��=n�� ��]�(��Y'�� L*b몔�}5�x@[s���y�������м���Ͻ�G�߭�q5���H���Áy����ח���{��nJ'��{��|n"�.���ϫ̭�*#Q��)#*S
������G ��������]�X���r'	��݀�9���q7���s�;�Ｋ����#N���*v�aU����n:2�UhB>-�cmq�œ8���r2��.�.���Հ�l�\x�d ��l�������)�Q�ܗ�9G���S5�4�j���W5[�Md��΃A�hv�e=Ϋm�%H��
j{��G#�[>X>{!��!����vgT*�������x��Dx�q-�����s�޴j6�[f3ӽ~�ۭ���{�����]��U�h�G�hi
d�6ja�Ds�llRt���2ǯ�r�8��p���|s8�o$��[�����r=3�'�c 9s2T"��0�Y��q���V�|n7A󓕥]�R��n��#�W������~n�fn��w�!ހ'�u ҖOW�&똹��g�^������)7��^��ב�~<����]~�=+޿��M
�^T���ꎂtuB�n3��s�IO{*�c���C�u�v��|�#�/������������7�Pz��t62Lyu��4��3VU�ה������Ot>���92��9���u��g�潧�w�z{���� n�/A�so��N��A�G���6w��N����ʈ�C�����*U~*F�=�� ����C/#6/�aJ����+�f�����u8f�+h�5:n�;��2�Ew���r�V�1A�v������>�~���C��x�z��!�!�]�����qY>W�xA��z=�֋�)�_��6/�nP�W�@!_�W�g���ѝ�A�8�1��YV��l�?���uy.�+՛ئq�ܤ�G�x@=\�GkU�+�R�S	��7�RK�Q{�W7dл��KiS� g�~�
ll=�?������[��َ;����R0� �]�K퉦��G�������.�)?�����3ޢ�'(5�����9\+��R*�$��tL�;u���u�ͻ�;CşA���F\�tZ�5��w��T{����T{J~u��O��m�s���jϑ9���I�P�m�E�u'�}^�A�iߴ真�#�'ǲ}$�Ts���P�э�U�3�G��P(T FX�*|i��������O���ܭ<J��1׻"RJ4f��O����^����S1P�J5	Q�2[�"�����c�u�>t-�{�ݫ�^��~�zw�������:���:��d��a��<LL�WQg�huB2���;x���=��~L��*�Tg��`����c=>�O�#�tx��~T�@��Q>�d/�;�Vz>����;�tO�]me�g���;��q��B}>��n��<k��C��H+ч�+j���K��,��v$��1�C�d⧷�.Jkr��C^�c󻓌�zJ����W�i�e��@zkӂ�s���:+�>��g�r��Nq]^��"���������^\,��]���isHg�#�?t�XNᩐ��B�+��[�ddr����p�+�c����u꫿Z���5u8d��K԰�uo֗�m3;��)(�8��/�qn�+l�2m7���WH��	v�Q!fw۷�#��oI\�_,�˪A�]�]�竄�ͼ-T��LP�5O	����:���Y>�1�'�����NQ=�,y�	{��]u��B����E�|��q~��ޚ7��~�x&�����{��_�FoЛ�1q뵾32��oT-��
�������2%��ǽY���U��Gl��R)N`0��l#�o[�P>�\�(S�E'w�"�Po mxQ���"Y^��^�|myV�ȇ�³�$�����ίy`*�=%��j��;�;]>��s�=�q���|���ת+�z��O��8����=Yt���z#�rO�$���C�L;����}TQ��ޫ w����������3�^φ]�r�/L�3�����f��@�� �A�"�}\��Ig���7�9��Ӗ�-���)�z:XxK9��6�;%�<��`�2/��۝���T���K�����~���_���W�z2��+|��W���t�:(�(Hτ'�/!Uy�E������sy��2����G#z��.=>V��O���RM������+�<�?ݏܶ��LyW�aԧ���#˶4����>� T#�ӧJV�>�de��b����f�X�F���>��͵�t��9�A_�h}� 66w��������t�~.�5�t#G�fZ�����7�����z]�&�7�����}r17�p�kfNt��b6_S���5w7/��4��oS�G�c8�֍F�~��Dzg��|r|�����;�O��r��h0Yo��׏c��ސ�3�l�3m߅�*l��r�o܅F��j�&���'���L�c������䪽#y���3!�31�6*mV����^�y�񸆽Q�Ԛ���-*����ì����N��ˁ�N���E���ɇ�'�b�w��gժ��r6�f��V}����Ii����1{�qq��=2�=�z�Ղ�F�������HvN>呹���+�}|�O{l��(~Y�lxgUׇG�W��k�x=��:z#�4+��{,��Zrc�7�5C}��\�g��)�A�Tz���"�}�����^�߁s>�L�z���!z�:�7+A�G��!��'���eM�'}��t����.c�=�z@^%r\
{�~.W����ݶ椮Hsn���u ����|k����Yۙc(L�W��1D��#} 5���i����1xW	q6���ŷ�~L�)��z��{>u��u��ز����g�]U�7\�=�^���6��4��Ƴ������ r���և��q���F^���{�-W����	R*Xh�9�Xi�وA1����]\����T;a�Xҹ�h�T�@�L�-ƻ�ZNC2wn;V�])��딠�P���V��S�'A��p.+gNb�ν�]���3Õxq��7#ާ��Q�3Zc��x�YD��3|���v��"�}7+����禕���,E��^��p�x�{��u����&�-!��< nr�XT��vж��.g�g�c��z*�z�x�}w�q^�\K�^��s�{=�G���2�Sљ� �����Wݒ��<�`�'H/������y������\Mǫ֑�L���V�]�ߓ��o��G3W�1�F}
dPP���H���A�+��w��Q�j�m�[f'��V]��<�s�׳�F�����9��n��sl�D���50ݎ�&&��h]r����^��=+��qV��u��������y��ώG�wļ�Tl	�N�R,��0�p'��D����fc�����[��Y���׻k����dx[�~n�M�O��:��L��K'��ǣg7}^tV��^�m��d�_���saV���>Ϸ�4T>�[�~��x�@z}����&�F���I����4k}��qatK�,j#L-�{׺r��3��}��o.-�W������}sW�25��}����w��[u�^�v_�I��c�9d�ݱ��^U�nI��E"�m��l�mUM^���[�%���F�&F'��j	9kpf�q����}J��J�7��F�:k1�*.��2*&1ٲ�����Աɫ��ݱ��o6�YSD�7.м6t7�~�<l���x�A�C�6t;����/��.��y��=�K�����QH_ضw��^�ޥ���gZ����Y���3��Daʙc���:��R��+K7#[�r��}��z��Fg}��R�^���eꞔ+~���!�ǀK�evUX��ޫ�1�����V�Q�
`Vx:������5��9^�x�wHof6/n�O���,53n2lzs��5���Jk�]�G_�띓�n�o8��C����q�3��ǜ����s�.ʑ�k$Fڟ/juY��
��e�?p
����7�я%Ҙ�uP�^�i��I�{��q��^
�Y֓Ӌ�e�^в�=��d�r�&~'�H}Hۤ��F���q^�A���N}�'���ֻ}2�����uv���Y�B�\m���]�6
5���T��L�P�S�*���n3~-{�5����&�A���z��}�:U��=2�b�(ӂU}DO�[�"�O����2��]o٫�N���޿��3ӽld{��M��.\��2Q�o`OA�w�����l}��B��I�����kmI�oRØ@.�v���=���i�h��������]�q���ȇ����0�u ��k&��{un_ �8A�{,C���kosgw7gg�!�:�Ł �!���F�k{��r�ja��:�6�b��]���єs��s�>�/��c#��D����>T�@��Q>��e�3Q�c�;h���V�c>*`[u�;J|6�U���*)>�I�7^��^ w���uܽ�ji�ɛ^9��lw�>��<(̮7\����"vW���r��5��|�W�3��=���<�w;�4���{n�G�&�L2nP�p+��q��_�F��M�]ԧ_������`��ā��%�1��/#}P:��]������@Ɏ���]U{�FRt�Y�����(�Ɓ����{�˴�����g]ǅ��^��߽��}�y}���f�����3�sL1[�_���f��EkH�*}^���
���2_���{՞=��U�`������^��	����͈ ���y�h���Et�{����ʙ�����c��H�r��9^�|myV�ϞWG��S�q/ѩLX����{�M�������&V+�7[=��0��M�Ԧv\�g��4�B�����Z��\T�/�z�
���$��(?0�y�o�P>H��?;�������S�)���F����P\��j�~x&R5���&��,=��ϝ��Q�t�i��4�K$�m�4�d�sF^V�K�ײ�tc���T_^&�����A�֜W4Й����@&�7�g:qp=%5
1�Z�a�
���r�|��*����}�/�dz�ǐ5�b�Q�NH=_`@�,g�ʼ.1]U�U3�P�)6���o�I�O�|��=L\{d����}�m�v.J5���K�!����*|D9��ԫxc���u�z���H�S��og���\z`Y��J��� ��\�������f�P����o�+���u������>V�G�k��ǽHq7�IQ�1^�fum�s�
��{���9n#r��|T�2�\��@u�ƴj6���r=3��9���7�l�;]���G���k?`��h� pό��l�3k��^E*l��r�o܅Fߚ�I}��"�����4KL�>�χ<�V�.i�ȤY�31��B�mV�؝S�6��>+�p�4"�e>�����O�=��������7��{h�>�$�"���d���1S���57	d�Ǿ�Qݝ��<7�(o���	��.1���V}�U��*5�H�,�P��ӬZZ
����1����Q���w�s�s�,��c��3�/�>��~���O��4){*FlDW� :�"���"�?<'y�+�+.�؏�9�Ғ��md��S/�E׍��
��kjG%a#5�7����c�7G���;V�
�_gf��&\}'��d{�L(hdm5+^v��B;�����he�Z[��T��x�
�x�mz9N�J�ӌdur]�)V���T��Tg*�rC�u$��:�G�ɻ�򺳍u��T�����-����[� ��R�7Y�Yc��H�JѲ�u�h�S�0n�k�yN��ޙ��S��@�q;yi�iWn��.B�qy�]Π�ϴ�.�9&�֭���Y4��m�"��ATQ;�GլU�7m)>Mg�ӱow�ʡN%ׇ�|�V�Z��ֆ�mmp����'K�4.�	YX<����͞��[��Q<��˼�x�9��Ύڛ���%v�If����sN�LtB�wD��	L�A�@&�R%�\��wt���)#��Nڵ[GwF��j̜t^쳀�wv͝��0�5S�F/5'CYÃ���,;��n{`yGD�;�|pZt�X3ۚ&�}i�'q��ү.�`�q�rPS����!5u#�(�f=��Y�Y�$�2�r� ���{n��Ks�οn��J�sO�����hs�R����m��n���$�U�������˴�@���S�϶�w��oHf��ɍ�T �[��uc*���-��nSVښ�HY�`fa�29v%� M�)����St.5vq��W6��`��ej���o!iu�/1��X����
Y���o��X��ˠ��={Hn/R>�}��ل�|h`�����v�FPK:J�Wfٝ�k�b���)~܏=&�98�U���2:���Fi{���[;�DZ���d�d����};����o�Sw� ��2%��,��[tH���`V΁�Tsgg�.d��ם�Z�V��D�y����7Wk��E�K�P-�	b�(;KvB��X��p�>�k��@nK��VLe	�Q��cfXʲ2]�Ă��-��Y5���n�R��b-���h]
�uhgs��A+�#I8�RΚ�]���	��R.Y���TGV1��S��:��Y���L�3�T:��S��p�	���4`�I|S.�Ӣ��Fo4���{���z_w����昏�^ͭX�&�\މP���k�i�hv��l�{�sE# ��P�u��eQ�V��tI����u�-��m�-VRaiRܟ�<���7���U�П�kgR����{:��
`cv��k�3ٽhւ��i����t[��ݤw���NX�O���#��rЂ��B�N�]�[F��q����^}bD6uYK#�?�O��M8��j:;�Tѣ溭j���y#�;�y����b�E�*v���1V\�Ѥԧo,��6��$�EΠ��gZؖ���F�9�:�{+ ��r�f����v��D��gm��q|���OR�o�>�K��]Ȋ������ʗs��)�D�*���pR���E��9�tʜ�\t琻���d���" k�z�H���㻺����Es�q	S�Ȥ�$̯W:Ts<�*�ɚ�wuѹ슊s��Va�\閦�EVheVe\"���/ZQQ�L�.�
5#D�(��T�K�e���R���B#�jznN��u���砑T��E�*�Z���y���!;�8�'��+:�.9��*<�"�Ur@�fE���nc�L�09R��yJ�!D]ۺk������]�fi�*��痩p�!qc��6QJ��Z���Tt�T�=wh]72��Ӗuݸy�H�\t4KRn�"�����WP.ʯ't����\鎈Gu�sEK��"9�p���<��G�����&e\*�FQ�EJ��WM�
�(�V*%����.�훰��~������9�ܚ�r��N��6z�vd��k���:�iʹ{]2��M�"%H	�.*��� s�W�%�<�ĄwYo�EL�'�B�b�|��"]W��;�Tw��/]Go���h\ǣ޾�9�c;S��p��Sӕ-o�,�6�>v�gʙ��~5����߆}.W��U�Kڴ�>����V��g}~��*�8(����2�P�১�`��."��~G|�} ��^�;oE.��X>{M2+���;��6�tgeN����(z���Ϥی�O�c��|�5]�;A^���φ���h�1���q��p3�3�*x�YD���ǇG���aR�x�c�Z�v�1��=�T׮`��o,C^�`Q��ϣ�D{���qț�T*OUחM����Ǥ�g�U�I�c x��G�-C븟��.������{��#qRFeWOd�&t{#�{<9�~ɟ� wI��T��W��1�\k��z�9��\Um��3Z)QM��{�~���FF�O�N$5�����1)V�W��/��GZ�ǜ{���3R߻W���>�1���3���'�c5ͳ"��^�50���&n}ƅƹ��uϿ~�MN�Px���9�����G�UۊM�D��]ː�kH��|T��k�a�y���*k/����ƍ>�����?vC��v���͜�9��PJeJ�DR�vS���W<�m5W�qo)�ys����:���.[��F,'v^T�,��2�nMv?;�g+#���G��G�Ǧwļ�Tl	�ө�'��3���E�\t��΂�Օ����D���K�[�A���dx[���ħ����ހ&��R��c��a��qg����R�˿G3��P}�]���W�^o\h���c�]����W���d�i��:ʂ(�ڵ���{�;�����_��o�����E��_)����^G_�J��6q�(ʫ�7O���=�=��]
�l���
5%p6t;���K�x�/��u��n�.�������έ�5�����#��}޻����M#���h�9Q,~����Ό��W�_v�����^�m��ق�
��`D�z�Ez�ǲ>��r*Ư���l8.�v��>�UB�u�j�a{!��::�t]�#%H�K����"��z�W��+��L^����'ݙ��{���<wg�}�,�3�,�ʨ�����w�<����<�o�d\{g��C�1�^�<;"r�.qO�yG��Uw�P�T���,����$�_I�5�W]5�>ȋU�������z��=�|^���N�{F�>k?9ec�!b�W�5Q�PU��X�H뺲�>��KM���M��xv?��v�k�f��z��F�(�ci��{��s��=�ޅװ]]�˲S�ox8Ά��߳��n�e"��Nu���%'Lާ ���Zr(��Xk+y�B�I�˪�}�-�I�{4J��o�n�W �*�S�I�%�#�Hۤ��k�>3�M	ߚw�#ԥi�l�tnNA�R�-6�9��yI���<�d�]�6
5��A�&
��7�[,f���Ӟ��'n�����]���>B�]hh����v#�N�{�=2�-�\�i�*�������C�Vw?Tg�o�e��ភ��������C�z����[��.'ޘ8}>����]�o};vkm��V�׬zɏ}-WQ��K�}��k�k$h������>�8<Oy΁N����e�3����7�{\�q/�#�Hɾ�Vr)O��Ϲ�?&&3�5~�{ޤ�Ƽ �jQ��m֍s}<4�^o#nǣ�.L��,�f_��S��_���u��w�������D�pt_yY����\7��|�2}���9�*���L��0ʚ���X��w]K��j�/>ޯqP�<$Ev❍���4�,4wў���do��/}2�ެ�Z^á���'uU�:�f�\)�*�����s�J��c��V<;�:�g��w����z�q���B�T�,�����?sN����r�oF���״�u���4��󻅳�,�'.��K@�䢐%A��}Y�`�����"�N$ntױf��d}�3m����pnD;6tq~�1��\��q�]ˏ�.�w*Xʊ�u�CPQ;��N���5>�KGC%��6IM���2�#芕\d.� /|��D�V��{վ+������Q�ʑ��3�c�4Əi>y�<������a{�[w�*e���k�
�~~������Tc�^s����f�cXaڀ����phܝ��C=2���
{�Rz�\3�� �4��O�^>��9�Swv_�{�s�ܽ3�L��߮7�Z������z�P�@���,R�,�k�Xk�+�M�{����i�2�D��=���ȇ�~+>���,���{�v��e� �.�Q�zh��2Wfygr��m�2�hJn�����7#�Gǭ��{�ߌ;���F�GĕPe���#��"j]�ҕ�N� �9���/N{��}q^�p�z��FG�W�^Rp�J:u
�\�F�`md/Bᛴ�^�4��@� f�$il��u��*�_z����y؏z��o�zH׽�fw��n����ý"}�=*��P}$L�\����~�Q�h�m��l�zgx��2+���T���ώo�.�l������Zt�3J@L�-�=$L���yJ�<;C��~�*6Z��JR��Qos(xb��J��X��� �6��ߟ�|�wD1��2�n���m�ʽ�/n�dXj

nwB3X�k���C'	�
�ױݥ�4�sK�� V�\�G2�h���5�5g_;ɋx|����H`�>jT.��B��@8K��Ӑ�E������Gޙ��u�O��̊�zk�3�V
��]�bu��~��ڜ�^�[���g�wS]$yQ��ʈW��L\y�Y�o���负��H��5�~O���}.����}շ�wg���z+ޯq�ޯ�+�b~��q��=2��z���`�Q���d��U<���{k8/eUz9�OxǮ����R����~.#:��2<��5��%�o���2=�H�v������H�Q9�#gv��EV_�ʙ|O]/��:��3�����;�K�sZu8�ˣ0��.�HL���{/����O�Ӷ^��t;����$��;.D=� ��������#<]�?���w�􎷿T{����h���ӷIxc��	t��g�DT�r)��?O����m�.{f	�ce��~���r�^�Y���F:3*���l����+b�cfl���M�;�kKc-�>�������a��x~��c}�~<�t��A������=[0a�ey�zi{61��D��;Z.�W�ӑ���ݼ� /z�{���8�Q�~�=�>���\��d�=3�1^�d��27�5^H��<�H�ЛvbMgJ���%]��f酉�YО[N�͙h):�m���YYOjZ�z��O{n&������a�UᣩS�����J�0��24�gIeJ|A�
�α��"�n���
��u����f՞g���0�I�T�[ڨ�oj'Ν�NG��9�t��4��v*:8m���x+���U ��l�P� ��K�&u�n#��^}��#/ʢTz�i��0�.{�N��ў�{O����W�������2
.g�Dķ\�:_��=�z##{�.�ϻu�}�����c�:�.=3�MǝA�uLȥ2W����w����^SCw+B�!����3���{��Ϗz�ǹYq����O�������z�`L:u "��&��+�^��>�[��_s��3��}g"+e>��,y�;#�ߕ܏7>'�<g�w��_�����1)�i�n��o�.�ǲ��s����l����k�~�q���������`E��Cf}Cc)�)���y�H5��U��n�u޾�WKG��>����c~�Dyߪz��j+}��/gp�<'v}���t+�/&r��`�������7"�4J9�/��27|'��Nv{u_�,4{ў����(l?Uw��UA��xP����>;;q3���·q[��������w�¾�]Z&�Yʙ'΂.j�5�(c�ҫ��t��{8����9�KeCu/v�QcV�A�����W��9V�v�		74ްc|�������~-`x�y��cyg.����xҹ�]�A�QGV�uM��Xj��
)u�Z=��x��^�^���< Ȗ�~+՞=�Mގ���҃'1D��
[�ʛyW��w��(�C�Iգ�T�������dK�S�^�x�wHu3?EF�W������Yz�����~3��2�����w��z�C�����+ޝ��z�hxw�<>߼$�{�Ȣ����Υ�.���,q��}��j�Iy���Y�n�@�W��O�ԛٯ�����8�[��gОϡ�R��]�6J�,z�X<��q�M��t|n��,+>(o��:�u�y�&���G�����>=y�p� Ͳ�P@����9e����xn����(Zz��l�^�z�ў}�h�yIҮ=ꃕ�aE��J���O�R����3�߱�or-�.R�����Z�Hh^�;c#�N�������ި:j=^���(��`�ע��{��J��[�	�`�K��ґ�hu������2#��D����>g �f�Nt���Dgoz�5c����N��dy=$LM��Y�R��Ʈ��К�I���H*z��q�C}[���S�uND���g�C�[G=kٹV��n�5���!�Z���67h8�^�E�9C��ƚ�� ���O&�Re�8�7e��)���]:�.e.�v�lw�8l�2�B�.�D$���f�eN]����]��{}jm��z��U����r ��z�t�&n!O��	~9N����J��.9��m{�={�ə=��.�|Vv�>̐|��;���>���ʠ���(�*t��=8�u.<2+���p���f��&�w|��>�;�u��]���/#}T_ެ��ٛ9��ꁓ_�6�?��ƽ�0?v�ū���>\l{�~�JϷ��gUX���vxw�w�?���F��(Q�T=�8.�)��[5�X�Y��j�>�pm�~����"������μK�k3��o�^���g�M��=�y�����F\�zF�������E��\R۾92�K�^ Tc��H�W�&}1kfv�wNA}���Z��;ѷ���~��_�DgNI����,m�L�5z�_�߮��Et�gz�w��W�jrw�q^ z���;ǖW�[ɿ&w=j����Z��Ͻ��X����$�J΂\=o����\tYN7f4�_#�����nv��A��	W��m��/ǽJ�����G��7��X�>E�/28�G{/��u_���P����'�|n����C^��=Ln{������d�v.J5����S�!���]�(�����h��$C+����-�w��K;�g=��߼��d�)5n�#(��;
��<{�eiQ����z�S���Z�-43@��8'��#��һ�]�Z6�ހ�FS� �40�qh���i��\�H���Պl:��j4����޻�`��|?d�}u�����#��X:#ϫ̭�*:Uǥ��:�*��}r&r��+ۃ�l�<D��� &�q6zW�݀�5��q>�+AG�k���ԇ/	�}Q�UH�T���k<F{�LMD)��V�>�&%��lt�}��Q��kF�[�6ggy��3�q��r�=j4s/���h6�h�ٚ�R�5-���D�oօ�ԩ�ô9~2�\'�\׷S��^��W�B�$8�Dv��7���㞙��82�d$Y�3�V
�q�x��>��v����ޚ�]��B�\|�$yC�o�d���{h��2M"�ꁓ�M�(;�������=ˣ������Wz���#z�:���1���F?H��(����X(TkʐW���G��į��;����c]��0�}[�b��=���p���/�<��>��𗾫N|�b�"���Ivz+��]��<�d_�Y;@�^6wj�V_��_��K��w�.��霟���5��ѝ���}wPz�ܽ�NT��e��?���O�*g
�}�4�^��T�r�����Ǒ���"�]M}����T�1��{.�������s��M����'1ܞg�h�����!{�c-6����j��K�Ov�����w��{�o)�H�����gQ�.���L�(�(=��V-���2��.+����&����^���K��^�
�Eɾ��g}�zv�L�zsǳ�y�r�[ư�&t\/Iӷ2�T	�
⺽g����ss���m��r��S�P�>�~t�|W��+�����#��:n�'�̱�܈�n24Vx������ܺ�Ǣ)Ut�nXk������"�������?�~��U�S��y���P��X!����+l�^3����R�-eAv��p�����'�;��#�?[��m@��`�>�z������?|.K5�,���z �G]0�k���{�&�ӿi�'�w-)��zs0�t�a��wa���=�Ftς����<���[���Z�uc��~W��Na������]E�zg8��ǽ'J�����g>�2
4ࠪ}DL�\�:_�[}�
�sZ�K7��;'�G۽^��6a��޶��zg��9���fEG�d�M��n:H�t��f17u�������������lxχ��r�:���1��+>9����Tl	�ө:b"�=�.��xv|5*�E�'��DJT��d��yʡ�ϕ��s$kJ�-��ޅ^������M����у`�����cm�c�����`��0l����cm���cm���o�l6��0l��`�1��M�`���`��0l�z��o��6m��`�1��=�`���6�o��6m����cm��l���d�Mf#3Pp;~�Ad����vB������x{l{�l�J�����Z�5Zl�j�Ҋ�Q )�[b�,�Y!B��:�5Sj*�Ƭ[U��L����B͖I�jR��TcF�3 ,�7pEL��Ml�R�6�&�cF����l�&����T�Y�T!-���{۽ڭ�� �z�Sض��a�.���;dX�Kj��2��Z��Yv�ȸ�&��妞 ���$�8�m�)�������eB�)��{�  ���Р)�}��}��v�@��;�����DMi�� eqҔ����u�u��:�]03� (́�n� ;GU��6թ#� ��h��`4��SF&M2�� D����c���l��uҼĶ-����� ��KE�MztP{m�{��^�]�M^Ƿni�Y�w֞��s��{ޗe^�(+sZM�f4ӻ� on��Iy�QE;���s������Sb��{�at�<�4�Nv4V�z��]:5�Q6֖�%5^ w�Qg�@��pP�L�͖
wa�tBN�z�oT5��)�`6�0�M���J� ^�CY{� 6� c�����N��Ǝծ�9nc���.���*�Xk@׀���H�ӥ��5k�\����t��v�����6�
x �)Zs����hR��@��4g]p�8+cv�g�� �   �  ���IQSQ�@��	��4����I(���i�A�F "���J�h       T� JR��Q�M��@ �4�D��d����eS�SD��7�O5 �?%(RP�0�   0�����[�<�~���y��x�_���y�\q�
������*��!�H
�OZ����/���%C�ꪊ����N8�������k�������Wp��'� ���"����� ����QE_����C���A61�%A
 ���QM|>f����&~1xo?�忿٣����ַΦ��v
� ��&� �b��+���� �^��
�����
n}�DG�}��Dfc��m$T��I"�������_���?guO�����!�P���c�$#�s����QCN�?���s���dTlc�٤�
�d��aNo
;aVҳa�ܠ`�f��$��swtd�[;k�Kkt�wB�"��A�P��mn�U���\�L�T���356��+070��<�o)hK>D��5��uսI���,S@"Y�B��Ul�&-�p�ջU�6���&��:ŀ�8cAٱǫ�Hcx�X���l�3p`�v��]�ρ)����\�(�L���@��]�,] %ZU�y��Q��]3b9��� f��
ѹ	���n1���1!��73FU��>�\t�z�������:���k�A��b�{���锱ز+������NrM�W77v�-I�PaNޤ�l�Ňd;-K���a���շ��6���73/�80����ˤQ�D�\635���m�Kw�"�ҋPŗ�w*���t���n_mM�+B�f�;��.���)��Ĳ�kdf��pjЧ��շ�g����N�������}k%�
ʀ�.�ǣ_�ؙuO^�̇e�ıɏc��wsUe�`�&�{��fn�v�C�K%��0�g1��=Hh�4miͺh�{Ef@�@����V���#�4KSd��TX�y/"����f�N����'Ul;((���B�f��AM'T�+ǕR�][(
��n�ȫ������ΰ�o>�,��&k�k�b��*5F*Ijksh૚ݝ!T�i�V�%ӣ����#G1�_:{G4e�MH�uR��1S����J&��R����X"�(�2����i;��V�u��oh-7J��+HO����(���mS�"��9E<��4r�n+�OE�ۛf��ٱy����K��s�A)3��0${xz�ibݕT���-�m�G��{�,!</a�4�"j�A��B�1(IW���g���p�S[2S�W���&)-�Z�z�N'YtR��J㸚�嫲�SEW;�]��{���o��oPDР~.'N)��&�a5a�`6�3]�NQ�tq�sf��cQ5�9y�A���]�������[K��ٲ0b�YaF�0�i0�X5���\"��<�-�r�6���W���=)�M��V�*`*���-ڱ��֭����[Z�0��+�`Rx��
�<u�5�>O���F�s���z6��:Z���4�x��oY{P�ʟ\���F4���T܈e��1d�5��C�4UeeP7���j��)Pj�QU)w�wL�[�3|��\]���������M�z�k	�X�+gEn���Q�hf\Ow2����
ÝCb��g�}���'�Y��z�H�^Jn�-ǐ�yڦ�v6���E�H����s=Xi�;��v��y��B���m��Š�,���#`�n�[jP��!���C�T�U���(ih�/w^��ė�i�0R6l=t�-�D��V�VW5i޺����(�$�u��	���>ٶ�ݺkl��l}�Zڰ�Z�}�M���a��,d��YE�[F!��6�(����8��[��j��d�e�o�]e�9C��&�e"e�e��m�Yf� F��1��3]i�Z/r%�m�w��F�_
��� 4�u���Cyy�p5��#5��+m0��3�r�*O�s�J��v�� +�x+�,��>�n�'W��3G�[�eV:�smSǑ�S�B��1���U6EE�u�#]�E����Y:qv���t0�=Zur�f�����da�&ж35e��y�s�%�/8�y�i�K���V[�Y{32�Cmա�s$9�
5W��U�!����:�;l*����gR�aLBB��ۨ���TNeYj͍�+��KIY�^�eX8E�xj\ݷU�!�T#��X��[��R�$4⡚��x`���v�����CݷV��:wt�<�g2�Z����qX��-{٩:&bڐ6w�%d�����l2aQ�k3d"f�Ӄ7j�Ͱ�P�����%a�s4�ۯ-�I��+����G�<6Y������Abȹ���XF����+o^P��M�۫�UFcm6�]���`xK���L�(��$b��6�/z�Քsem�Tš�$P!+xwV�7F�E1��V|lǯB�\�h�I���<.������B�kr|N�30��\��^i"�4�c�K4�-fT״r����`�Bd%ޖt���k���Gh�i«U�����ӽ�56�����L�s,�`6��-�$�{ ���{��5�k�*�9Zά�ᬰ�ům		���̭��<���\����ͭ4�*���UKʦ.X2�e�3X30��e����ݓ�P�1Łj����.TcM�h�h`�r��6f<F�isC�`�H�V&��%X7�l�N���Y|�^-Uck�e���<5��	He���Q��{��n�[��{CrF�"�8NeX9���⚕��	m�j�娮^6٩AZ"�
n�?;8�PT�*���69q��Tfom`�ݛ4͕-Fe\�n:���*�R�!ś!����Vmi�BVm�n��N�m�����Ң�<՛,�W/,�ۏ��/��أK�*��t���c�j�L��p*�5���AP"���ס�N�7�u���a	"��jG+��h�8�8�
�����\N�)�PS775Fe��
���ڲ�N;�#)�Mc�*���^�߬IC.�]��Y.��C�M���f�L�j���b�
t}c���_r(�\-��sEԉ
�n�+�s]m�ܐ��U�^�cVS��'��,[h��]��z%�nҲ9�X�Q+0�1ۛ���=��Q�$��
��Z�)m�S�4�5op�K�hƮ޷K���9CnZD�n��-T��m�q@B�P�0�b#���V����s�z�y����c]:rj��Vm��,GajW7��ur��[���ZlD�U#W�a��n��u����c���8H{Kh�ڱ)VUG[q(,�;aW��q�8�hW.�p�������~+Slf�nS��.(���Y�O,o��̺ �쳮�ʴ���,��<!�ݼ8�ui�ocyv�ٯ�VmS;T*�4�̻ߴ�ׅ6+7�-���J�>�VCy���xuC3�t�	�(���(���Y8����Xg:C3��fb�|��O�W`S��F�A���(aOU�V�����p:z�����-5��7J�U�;v��m����X�4����D
D��c^�;�|X��\^��`��&w�K��r�-	ՠ4�u�mU�B�,�y[:,qJ.�*3+t��E�H�,��Ǘ��[�.C\񭴑��Քq�]<QF�����+w���u5vo�Y\�����C;��Z���-�IQ�yR4�=z%O%��AM�;�UPVl��kt��[�]$�m��È�Y��E&,����hњ�tF���H��187k��ry��>\���j�L�!U
��kY�R��f�4E��ä0kl�[o-Ͷ�B��9�	%)�Ya,s+qИ�l�P1Z����,c̵����b�xͳ�;Tt<�U�����W�Zϑ�g*�-�u��7����~91���R��� �8Դ(Z5���~p=�O������*y����H��=�w��wbj�)-
9)����^��|oу�čr�I+ �9'Xb�.ιvfI�2�kꎥqP��p>	����S��wFr�8mf��wRq�������<O	�N�#�8M�|�{+������R�\�kA*w%�p�"������5�6�����XWЪ��/)@ޓ���2��2�iP�͸�`�xHH2��k$�E��l�壡�r�bԤ�iw�g|�:�8�۵fx�zdBХ}�L��|���6Z�W�2��jCu�w�Z�1���e,�1����]�Qwhʗ�y���xgQ�xv�E��f
�c��(ۅ�;N��u��3j�<g8'32Y�M6$d+���j��U��)u!�o6�!"{ELܮ������J\�޵k>�wGRѦ��vdd�A��u>��&��J���\��q���e��od#�7Y|�`�am�3��.���Bw���J�7�����o��nE�pۉ����gg�ا�qü��SSڹ|~��&P@�cXZ8��)ܷ���Ǯ���:����S͘���W�*L��ކpr��#�T/m�c����ȏ$�tt�Jw.M��+�m�ZR�3�Yu���o)��(���.,۝X���g^S��������c"��L+'V9BkEï�p,���J�_d��G��G�E�0P\m[u��p��=��:,u������kT�zT)���I9;5���V^f+�ӂJpg��
��z�γ��Ҏ�lJՒ�U2�,H�g�n�y���x-��׊Z�'l�5=Goun>�`E.�Vw��h��7��S�x;Y90�a���X�2Q�t����z �9�&�yC]`:�A��r��MnV'���w��#���ܾ�Tı����^=����tBd4�7Yp�}V�4�yc�ǵ�v��d�k��ԦK/�C��l�5�>���D���پ�鷛��G��q�<�bS+��Е���S	��]�
M��g2�^S�����'gg��#O7ҳ��.�!_=LJ�LL�W8N�=���7������q7�IY�/g�fD�#+�D��]�WvQ�й�h�(�dd��X��i���9���[%a�Y+��S�Q�s�n֥�g]Wd�ռT����v6H�C��x7��a|�
I72ᡅ�&r��c%��.�����&��H$bZ.Vnh���W-��}e"r���2���B�B<�gٴjQ��Z���|+� J��r�*.��n*�k�_@����k�+wX	��Q}�c�������&b�':Yu�����ժXm��M�@^'jL�d�-2j�V�\�i���B��p���u��^�ͼ����3U�S���	��͒2�pr���ήC��'G^��g$���AL�:�]X�CB`qx�Ǜ�nZ�$�̢,D]��6�R��f����]��]�G6��Y�A�@��etpEƐ �j��q	�:�����a\��B�5k��>F����:��f���b��7��29��evuv��DYSe�n��;�uk��j�kw`��`m�8FW˵u��+�x�O8Z��;�� �
���VZ�W8��r��j��!)N�w֌)2�BJ�����KgQ����c��v,��Wen&Q���E	/Q��
v�է�����J���A�\2�fjf��g:I�ݐ�GϪ�Y��O͗j��ԖsiT��l�Q�w�)�ja�����^����V����76�]轡>*��O�3��;騍���JИ���;v��q�Zkٻg:ևZ�uԤ��j�v-���z����w`B�F�GҎ�g.&������\���u�9>�{4઄���E�@��g�\���F�2�˅Y�v	�0A���N�k�&s��V��B�j!�Z��z0�F�p\�8Ih�4�3��LhΣ��n�����{+j�	�1-A�0S�i�=]ܖ��,޺��#f�ݪ&����RoQ��M�F��S�p1�5É�_k����Uq�r�P_F�_9hqYJfI&�����3���W���֦��ח���a���i���{�f��V�LUӝϪ�#�AN����f���v �Ԃ���fT��Ԧ�e^�]����ʳ��)۱\v�h.1��to,�^�U����1V���#K�3-�V2�d3@��A����[�Y֯����X�U�L����;ZN�֞��mi�Sl���Aw �:ʊ��*��OZ����_j�έ����x�"�U��FT��{��vF5 6D�t�%m\h���g3f�M��kt����5]�³� ��ݣy���b�R�IՎ-y�[��ݚ*�Ʉ��
a�7��j��1��+JզJ�ܪ�%��K�zFiƘ�E�ȜjgZ�M�r
�|U�t�ojJ��Yʖ�����+~:콹{�8&�m&�3&܄c��c�HwA����a��D2�=�ëV�ve���.9ܕ�F
|��R�w%8nlh\��CN�;h�)V(�襎�QY��,�k�ŧ/v������⚾�bs��=��e��w!|������@���ﺓn�Vv�r�{�@���0,�]����t�;9d`뚒���EcFm�6е�z	���a�
Yxc9��
C
�K+�%���gq��$eK=f�ϥ��!F�{�^����e{�XPSz���m����)f��s�n`�WY�]J�q��9|�ܗB�mN����L��j�^�3ro��$��B�&��e�#h��v5[��]�`�Z����H�e���b���)�%��7 $�+�b�km"�`�v/����)�bޒ�	w3:�+�br$mhOe�1&��箼�h����u�<h�a1UmX�^��z`�Q4_�{-d��tb���S������(M0��L&�lT���PLN�⎪GzTe.:9E(9ul�ռ �uI����ޕ�䇠1fG`��g��w�#x-��wz
7�4�L(m�q;%=}t8S�8�m�;\��XU�&=�Wkr�&����H
��^�[}Q�l::����nK�*C��Sb��7���E.�Yӑ�;��ɚxV������
k�ov��)�R	x���
a�s!�fi��yE@���Q�����r�g����sV6k���è��.EWX�m7��en�`B3!��9nfp��w�p1���e˕\�o���4ј���mR;��m�+#���IDf�Βu�`k�T�Y�w��}�:�$3Vv��ε.	�6�x�*t�����4����1�l���1t�a��ۋ��ᛈ�fJ�Xk&(C|R9r>���ɂ:�0{l�}�����r�iǤPWr��`�2���	WIZ��r�ǐto���2��Z����2����W)'(�J��g���gjX(�eû�ۧ�Je��&ꥊ��uh��j�Ÿ�lҾ.<]�$��m��ࡈҮ�{��ڕu���������(HsF%��4j]���<�	p8�]G�P�V�̼%'�]�Ê�8�Y�88>Lmp��`�f>�ft�T�l�}a�uy�KC�����z�r��3��S�k9��wOOS�|;�����ݽ�����nv$�%g>\k�B��g[3�*���omIQ����
�
�Ǚ���`����m�]����e3O�����/�b�U��?8L8UvJiR�]d!񴲎#�1gMfr����������Y}X�	n�-X�X�t���3�����H�p�*3d��Ӻܗ%)Lw��%��.�[.��+'�7��r^ ,(P���� ��i!�/ tp���X8�L�V`�,�H���;�����2����ygK̋>�V�:�#&�٭[���4�yd����5y��G._cX�J�ջC���@�\���ɥK��:ǂ���=��Q*t�:Kie��c�Q�.��]��J�ٺ4�[w
��!a��]sy�%NMvg�g{v0"�a&��zԚf�%^�e�0���f˗�֍��mDUM!LW¾<ovE��V�e�f�d�s�I�MAQo[-o��8z����ԝ��ꅌ�.����c��l��VE����V�ぬ���
\.j�깄7R�*
gڄ�g	Zx+<{9;E�i˚��Ԣ-IrB:����2MwB���J9r���1���}���/�]M�p�G����Җ���n�D�����^-��ro)��K!щ�g+�d��<(�A�lo*o�V�G���t���u��>����]FT�7��m�#|t��QK���2�]����^�Mn(�QHE��0N���f�>�e�z+%�u�%o8��oeh}�0�G���6i��� ��m3|/�tu�1ڃ��D�U��f�a��'7���Y���_��7�z�M��w��2��&"��E�3� �KV�-�&�X���W�s��0�\er�:��L@]�*'j�P5-�n�C������VP:�0����S����ǧ���mM�F�H��nXH��\�Ht �e"!V��׳[�ǐT�$��2�0k�`�m��ܣw�5*,RT��r��O,��l�c.U�7�����w���r�9��u�C2���q��e�����p��k#��q��Y�,v�;c�^%r�V,��]jT�b��ń��M�9w������I[偘�:rH<�6��m���5��k���Ȅ]Y��.�Xհ>�0�	;�����W��-�$v�z,�Y�Q֙9A��[*�j#tE�M���3�����44)y���|�p`��R��`ޟ;)V���Җ�l��p��|��
�+�9gMi�4 �;�E�6�?@;G꺼Y��QG$���d�tc�&u'���ͤ�r;��c���\c�kJ�SN^��[f>J#>�ͼz�]��*��O���
Ïc{�x\÷�L�At�m1�%�d�'��tb�;컷�m7̶�u�+AB�k�=���}r����~c��C3���s]�[�K�[�'�O�m�"�&�d�*^�I�z7{N�D��%qۤ��T=u��dKfз��7d��b$�X���������۔%�\rʾW�a���,�1�� �b�,�~]�]��j�x�9l('����\��`�^i9c�̺Wi{]�-�m�g!W�Gg�B��Gwhk;`�qD�WU��K�>�ן�(��Q�Sw�J��gFn;��Aɴ9W�d*U��4a��{R_o|��WZ�'-((2೔���|�[�7:�L��1Vmf��̻�{��ji��$:ۀ�[q�ٜ>F��[6��9�5:��]��hn�yȒº�쬹�&���	��R��d��j6�TJ�ԇ�����b�ݰ����V���5`*�(G��Θ�=����G�o�Zt��N���er�Fh��)LP���N��yi���ĕ���m��OG�+%wW��+�W���u�gTYڭ&.��	g�����JV�����h�_%]��M�Ll�C2�����D���-%N	;V1�,n	�a&[U���b�UR�hL?M:sso�/��V3�7%�Rn����U��ɝ���ʔ��Gh��=k8W7׃�@��܋�5�
�(�b��K��,�ٷ���[4뺥���wp�.�<$�R��d"9V����v�ۂ\���ѝ�C7Xz;G+q�ͼ=Ms���.���es�;�RK�����.�GA���VM�-��FH��x���И��j��P�WWV��.)g� Ѕ-}�>�E"�nn��ի�n��7w�Ո]e�謢��H�7A��d^��o[�éS
�8����C�yg]2��
�e��7�_��φQK�U�`�CQ��rҌ]��3aփu}�҅3��xSmc�A�YC)�U�_c�R]\r����豺�8IP>�m�+s���]�x�2�ikn�W]�جQ܆��8=jގ�)�ܙ:6뀻�����}ϔ�%�y�>�D�%dΡP� �Ί��9h�)RY:��pU��V�IY�9��֥��vm�P�������1rCA�8�-���im��,���d���U�*��re�晤���[D�a�}�ro9\�ӘW�+���C�h�7��29�z-�{�d��
�=[�%c��Yt�W���E�R�n��Y�ӽ�x�"�4���y�5H#Φv|�����'�e�Sn���V���k��q�K�v�#�Ѥ��>X�쥙+N�V"XY����V�Fri����!��$,{*�D�)���i�&�::V�d���]("#��E���Vm�ݺXm�7rGY�2]�$e��n*�D}��d�J6L�i	g��n�y�<!�WG��|^p���JÂ�q��Ҷ�tԽq��;�ϊ�lW=�:����& o�R��͗�;�#¤u}c��%e_&�$�v�)̴t/\�*��G)�����k��f���͊���6�8��&-'�����u�Xc9��XФrA.��v�ۤ��h:�a�Os��CW�u�%Vz8�)�y���ԗ��73���ZO�|Cмv��K���+�u{��/i,r�>�l�mˇ3�S�4�\���PF\e��l�֕��F��ݺ�2�:�Į8rc�S�L���m����Rŋyƥ,Q���2�YS���R�H���0�����B�f	r��+��\�m�z�L=V_a�p�*�nƴC��H�'��gX7���[�x�.u�
���n�E1H��;���X�'�
}�@c̆��b�uKLCǴ���t��Õ�~#�r^�W��K޿�6��D	pP����D/��Z�{b����t��B�_E�pSM�1e��)f�v㿦��G4�MMT1j)q�ffvq�4��1�]��Y�O \���	6�r4�)����wn֤ۼ'-�Kx'��ٷ�]9Ń&/ ����W8���ι�a�7xk`-_-�+F0ӍU�E-���n�"z�_$aR-r͔�b�Kd˾��vc����ެp�PkTy�ӸpJ���Kwj}�4�Z�R�]t�5�vK:@��Ųf9�_�2K*��ӷo%�3X��-_G�J���|J��F���u��e�܋�V���.�e�6�88m�q�jS�.�ò�`V�6%u�2rcl\j���u�+�yt�8����S�67�%c�6dö��X#&���o���>���\ꇩV��`�4N�HnԂ�E��k�����G��0��?${A��Y�]v�^H�����p�YB�!�.3� ~��1�a��|�<p
���Ad�栣o��foU�}1n�Y��5��-�<�Q1�YMYy�-�2Bc�H�Upv+��=�YΨs)�L���ő*2=�5u��`�9rowT�\vf�2P](�:�.MD�tB�1fF	���<���]��~݋
9NN�u/�iaCԴ��.s�q���}0ac(�V�"ۧ��^6�ٮ�raCHd��㦖��λ��X��\E�1ӛi�u�]��X���Z�c6-��1��W���;(=H��jٝ�Yu����<G>[�n�L��b�K�؜b��+f^��l��%Ds����Q,�o6Y������o��;����8�>��<�-�rƸ.���\�9+j]�d��%~��]s��4�}v�����X+��ez�EUͮD��6.n���L�'[,4+�Tg��Az��[�&��:���V��MAL.a]�E��x�{.���k���q�{ ���S�@�c��f�4Gv2�qw�5�l,���1�����l�j:�y��2&r�s/[	��N�#v����
���N�siG�[�O!�P�eTL�x\TDW�G\���tle�s�۝r
ukR+m��g���.��p���3�**��\1�|������1�WF73A��#r����Yi\�;�Vt��h�rA��}�)M+?����}H+��f ��Lh�����e���z+X쩍E�h5�t��U�4�ޱ{�w[)w=��Ӿx��ɽ�n.36���p7	���aNn5��� /	d���AB�}7ٮ�)׫�8N�,����(g*�7�����=#]FNnr���P�"#<�Az���0�)�5�Μ� Α'�w�EUJ�q��qJ��C��ѯ,a�1qI�{�4R��(ZK1z�jI�� ������%�6���q��?hf�;�xAg���\�5�Ӥ� ���j8]5t3��Ei��e�c)dnE70��M�b�� ZM������۾���f�:sFrz�� 5�u����E�X�h�eB3����}a;���q��<'\kk����e�I1M��{M�P�-�IC=�[W=����IY\`陻(6
��s���Z6F��°iwS:������+S9���ڀ�gV�����|�>��J��yjf��s�e*�j���q�d>�k�y��D� �rˍ����pIΦ����]FbRPv�%aJ��ő]�h8Nm"�G�oG^��Lu��V�`;����[��7�g*)�ZR^�Q'QAn��Z��tc ��I��go�46;V'�C-���T7c'�<�:;ˣ󋥈�hsW����`{������u�­#R���4�i�Z^�vb�0S�s-��|�'��{�S�[�e�֚�遹<gb@0��/o+$�ݔ8��.C�
{]tȫ�e���k�"�ّ)6��d-
`_C�y�"���읍�<*PX��:3�L%�NSݛ�h�+��VU���˥��E�~��6َV�Z1ת@A�b始$Xg)mF����,e��^��̭�e�12�Eث�	kX�Y��&n�	�o�'s8�IǍF�\J�8��p�Z�s^�r7�I�� �����N�4՝�͔!`"DN�A�o����mGMU��f^"ap��[�3��Cyˆ�U��4��(�3Q���� �0L^�ǕD|�x��A����P�~���E>��jC"�[q/FE�B�uwk��BȌ�^d��!=���[�{6��7'�/{G�%g���ft�5c<%�˼}�����pW�جS�|j-��\kk�R�H�����=�.�d�e�6�&B�4nVr`�EދJ��w���z�NT��F�j�� R�k/K�D����%��H�e��tO��9n&����ܦ��r<οJ�㲌]uE�i��6�o���U�/;����O�:8��&����{,s��o\�,d�v�0� -�"�U��W#�0$wz�x+s��F�8V�0����\0��.s�y�y����3d����/�PP5/N���h@���i��S���&�.~����{p]����E-�x �Q�����M�B��
�����;��&�:�ej(*�s�*ܗ82�j�A��m�ቹ}M�ΔH�Ȥ< E��};d"Ȕ�"�m��\�JH���ykď���V�9�������S��3�y���5'�U�qh�)�G[�7 ��5�_ܤ��C��.�nLT�e��}�&�$�d�6��{�����������!�+Ĩ���˲���I�Պ��0��$�����f��o���{e�N97��Z2��@{��S/i�j�.;��ڿWV��x���]I/��F��&ش�sYu��2������Yb���g8~2za�Rno��B�f�v��b�v��Jf��;`�q�Rir�<���w齝렘��z��r�7��3��CS��^�oy��b�9���nV�U�m֢�;^O%N�yܲ'1�u�'H��*��$g:O&�[��סzѸ9w���F0ȭ7Y/7X0_��%�f��ka��Ol֠�.��ZV�t��x���y�b�m���5�+��ո�SZFB\Ț��ҩ���Q�խ��˿H�"/��!�	kF=����{rz�i���<1�QǮ9<�&J��WF�{��z�:��#%i���ލ�<�s#�Nk%�c�:�qGE��{�qjP�($&�J�j9�Ũ)��$�N����޺.z&�=�˖�����T���D�H���L���n�:���Xs�c{�CJ�F H����	FUA�'��L�[W7�M�*�T9��$�yr��j-#z�R3D�eNB`C7��{X$�Gd-���wo��Sx�׷�-��X�	�l�S�]߶2�"i��x`$Aۊ��B�+w�8΢Y��7��J���nu���|��R���r��!:�"��b�*���'M�7>GUK�h����"n�I������O��\<�M�w#�Ʈb0nf-�5j�����XZR�EB�fC8�����9f��c9�?0Sc��d�k�u��i�J񹈕��8��l�'I�Y�]����s�+�����	mW��޺��a^o�S��b�$[X�M��ٗuV�y��U�EK</��i�bgX�)�2ݜ9�:D�KUAR��Β��M7�¦��g�Z-\?.���4�᧽W�o9f3Wj�? u�[Gn��:{����<�G��/37���_�}��7��E�4�':*�s�]��ޗ�����a�0�ɝ��E���r_X"Ǖ�LO�خ������t��i�~�ty �����X�}w��繊U:�V�F;��~�5��ٌ��|�d���7Y�.ݬj3ӱ;�&k��WR0�+ڭ��c �Nq΀�O"��,�C//����BЈ�o�����fi�U�o;�|�@9<T�1����)P���a�R<��xvxt��[��~�Tke��΍V�U>c��)�K�I�Q�nQ}Q��U��Ý;��h�/��ܑ߯�S�i0M:���UB7�=��]}�ʿ�����J_��E����N�fjl�v�����%=�{:��fe�0�ӽX�vĕٲ�ّlֱ;��c�yu��	(���^>�XfV�*�̶h���R��/ j�ԡN�ԞH�8�3��
�sjX���]�V�y�i�z�a��‱	1w���TٲM�V�=��f��W=��c/k�;�ѹxh�2:���LVJ����9�2Gz��g�G7��+W+� ��<T���30K)�qnХ�v;mҗ4�{��;�/-��\�\���7�T��0�S`��[4��dj.7E��Ȯ����jE���}���
���w��4m2$�m���6� �C�n��v�6����fv�Le<�sL�l'!�n�}_D���n���0+���{��r�����,�rQ�끉s�zU���K��v����*,�t�$�E�I����u��oS��s�1�n�2�q�(-��0�J���s�7�hc�r��o���B'-!Z�q���B�j�IS/n�m���w Y�̥� �v+
�����8�ٻ8�2���x�	>}v���|õ�:��b��	\/�7(�Wnf�����(��A�
��MS�%����V�.��ŀk�<5�1<��-�d'�����Lqx��>%k����7cM���,��b��;��ec1��2IF�!g�n4�ݎ�²)��f=܊���A릵tq�n��4�o�t�'���	����dGR������䔟���x+RL&���Qz�v�{r;p�,S&m�Qjx�)=��	�՜:YF&�1I�y�"�2+B��g�J�F������Q�(����@�s���sqr5�޽����T�\ց�]�w�W0��&I���C�B6�WDd��n���s=�(�<̈��h����i�u�(b��^gw���L�KE�㵙�ݱ��C�cILcm�;�Z�ĺcd�۳���'�3Mm�����s-�]W{�=�s�0�L���� ?W�R�>��?1Ն?�>��銮��d8/���%�-x�ɳ$NOV҂�>/#�3�wˮ0���1�N��b�����t�M����O9����;�}�e���0�����e}z�9��99�_b:RWԼO��״m�?+��BE��G����t�5 9��)�@E�)�M�-��EE������Z�u�%jbz�LB�d}�9�4)��t��:�юf�N2�1}'�i�O�4�idM<ڴ�]�q��N�\|��*�y�'�������ō9�Ъ�ٽ}�����/�޷�YN�?���Cx,�w���m7�����F}���@\>�E����A���o2�&�=����w�n&ҒV��u�eӮ�K �,��kV	+�sGǑ;��%js��d��B3o��f|
?OY�z���U�וoUs �w�g\>Ɣ��$Nl����vgvh���Ӄr.b�.w���m�=�ӭk��$�u˩3@����=��~P����M.��.S�&���u�w��z�j-�N,��j���`�ME�#٨25��\%D5ј�L}��e�ߖ��fw�z�*G��f�������'�� ���f*d�l�u���'h愛}C�󰵻��l��Hd�ӌB�hg���ڼ���q崭�I��f��e::��LL��N8����*����;�W3A�<}�_cOpW�b/&��q-��Ǝ��&��u�����Ur���U;Q��q��{?s?7ݐ�.:��}�:��;��]$B�i�0a7�?i��������P���/��
iIV�}�2|��lI���}�~�6���el6��oRE�Rb�_צ�Wov�˅�L���l9C�蒯�^�����*�z�[6�@;]b���n6��?�	]'F����Y����DW����j��z�ɬj��7��]�N�!�jp�;|оܽ5�I2���|\�یN�9??X������
�x9�>����߾�p3�▌�Xz�h�@0�����1V�]E�qz#s���]�<E�;��ϟ߿i`R���*u�=vT^�]���C&0
V1�����	���ŬEʾ��b�����3�T�pk��n�t�ms��p�]���f�M����0`�3��f� 8?��[��LGP8�Q0�"c�oq	�q��s�=���~߷�|����=�^1\G�&�6�#h!��♝b���\�1����ۚCQ�����gO�~�v�����ms�.�s΍�uA��8�i�ֽ��s:�J��cC��,�,Q�-�ֵ�*�^n�Iҷc�%'����]}��R�<íP��$�7P��mzKE9���@�C����V�*�=1T�>���P��=����ʏ{QqCԨ��@��^�����^�p���ǀ��s�s���/���8h�#���G��}�*}�P&=�+x��z��*W���)�^!' ����� �}x���~�^�x|w��~�9�9��Ӂ������|x{xAo��\�q�F��\9��)��9���>O�}����ϧ8~z��BD3�S�L�w��b�Dy�6 �Q�5����L����Z�5k�;�:�{B�1���Z��TE���{��*qj1�[�@i���D�<������>����;�7��}��7�QLD�P�D!�0�*T��n) s���7���D��9��{�~���|���ϧ9�3�}p<!wﮜ>!�o8�>'=<qi�&�Au1Ju� s8�PNb9�7��z�X�y��懘�
�. j+�����Q	ۡw�b=��?9�p_/8;�ω���?�����ߧ����NHs��R�n7�j�1	��1* [�\�z����^Y���2�o{iTl��w�ӽ��AXf��}�FB	x��r
e����=�{9q�;�-na|�CcA��9�q�������(��ȕ�R�������~�^�L�y�x�����s�����
"������6�*V�d^��ˣY���:��xq�Se���hb����*'1K�PN`�D7��:�b51�y֭�7�y�������y�tUZ^�z�Z�<��C�R��Ķhu�[�7,�Ax��H��z�:���s��N"�M�z8�y�D/T@B�R���#�83JZ)��X\@�K�J���&+�:���o:��3�L��LAvD/��aK^�As:�y��H!�73Bs�J�7K��jۙ�q��޹ڇ03����h�tsHb.�Pq��J�f�;� ,^��!j�1\B����N���]o�o��q���SP@s��PC'n.��=N`�D]�Aw��;/Jb7�Z�泾�1��u�=t	h� ��05:�bs���7B��CsQ:�w3�s +�T��y�\��y�Z�w�+h����/09���E8��9�H���p�9�uw@�D1�0_��*cֺ��}�[���詇TG��-T�+X�8��BCQC�TZ��T�PB�����E9��z:��)���R�g���(�h��	B^jU�s��f��;r9��!�[5�jKB�z�]��0�\%h���M��;(�
�agf��HH���3����D�����J��w���":�H�s�Kh j/SqIPI�����o���w�J��7�D:����EɚS��S�
���Nb�\8|L~��Ǟn�ޔ���~����8O�I8��������'GT���:���P/�T�Y�m����u�5ŵ��Z���I��9�1�)�+���Nu�CR��=���o8�����}�%��||����Iʀf��/дG��1I�Wp5����P3���*"_�IPMF�Qw�:��/���`�BDy�"�s �=Aw�B��R�^``�)��Z��jQR�(�SPNkX��7�S���\��H���!"%��N�B�bը��S������B����� qƞ7�j�뎳��\�j�Q��D$KA9�����x���qH�!j��V�p�T��q�s�s��y����Ͽ��x��翡�����"_�`�OQ	�mqqy���.b�/0���"�D�q�ٍ�<������8Ou=&N���>�o�4!�Kn�/qN�)��7sp\As�T�J��r�6멌o�fg��9�Y�(CyD��"�_eC����{��XWu��Q�^4��q��#�|	������E:�g:DI�Lv�)�|�ms���8�H��5�)R�5�.5@q���)��%�����迪:c�r�=��z��⣟-ȥ��O﫜Pr�����緀)��h��l��)�BB��"j%�B�l��#}��ֻ/���ช�8����TP5�����:�!�-�I���^&`�)�(Cq,�+<�x�{����W���5��s0WD�������?��������rz�[��T�[�L��*L�^�U�8�m-gt�v���Ψ��aic�yz*�t��`��'�ne=\��O>����5�E�\���V&ч=:�*8����B2�;k��Sual4�k}U+��9zu��e���>�j�zi�r�����e�_-ڹ[�k`x�^垚g5�Y�ٯ��'TV<,lvԾ��XMT"���J����.,�ȟCӥ�}��QWRl�{��ҳ9e�ԙ+1G9b����`�$sh�`!ZV"LjY�DGn����J���K�{��Z��^l ��۽C-k��.fa��]���S�F��=]��e:G��#��]����r�\�Q�'Y��	� ��3���pCk�#�~Yw<Q4�g�fc�|�\`���1n���T�8��M�/�׵��P5|�������u��By�[/ƙ�B��4�͟��,x�L&��q�4�nZIs4w�;%�F��<.OUm��G<y�\�^���]�<�lFi�%	6V-�ȯ�" ��"�DL��.O��M4���U��ڇ<d@k*��8���'ƍ|qnm��]��y�3�¾��xM醶E��c�v
�|�H��5Jʡ��>B���<�mÛԲ���n�&����kj�n��a�V����N&���Bj"�'�O U�Yl;�[v+�~�QΒ�T�j�����^�l싵Q"�Io�W�W�g�]n!&�[�87�"�����%щR�q� ?��^�3!�����-]u�6DQO]/)ege\\�d�+�c�(Кi�ڱ��Y�)�g�E)���70���{/7+���]����o"u�HfwG�4��O���t2��݅b/�$ga��>K��}��F�V�6�
��:�u8*�?]��,�����˭ȋ@�=[�2q��S�;�e�Z��[�-��#RbY|']bK*��.��EnJ�{�v�QF%YJ"���m�OM������M�b=v'T� �6qge����u��ufF��c5* f�n=8�[
�����V��e[��ZuTpA��t#$y�.�����/��Y��xY��n����&b�ƍ&9�ڝXv9ǩ��X˃��?e:k
yy��)'�e2�r�;�BWky�[/Y��g����yy/���S_�uD�A��S��T��2��H&*q2A�:F�"k��1.yY�#��S%�
o	Xi=4́�;^�jݪiD7���B�Y���CTM�q��I���SZscN�bg��-�AxpX�zkD�Ft��$���gb�o��wI# v�M�h�K�� ���,;Ww��/,u뛳iԘ5TМ�J�$�.�9FkC�BP4��K� ��Gv�ܻ/�]�'"����:�γ�i2��w�bۗ˖�X�jӏ%k^�g�s#Ğ`���?�dH���}�Zx'a�v�9�>�IF��ܧs�r�7��&=Q�����97�q��HҌ���P2/l(�x~��{�d��	\��o��\�f.Nj.���2l�2�;���=S���b��w^Ьt�D�j�#v�Y��C�D�#�vjz������ۺ��-�{�{�.j��piY��ǱvTUE��	�Q���B+�U5��g<.j⎭�m��W]q�n*���Rd�*Qx�ۮf9x��2��۫�uz�\��[=�؍�$�ݺ-��ˊT�EG��焩ظ��{�U;l�{�(�wX�'YtSݺ�<H��U;��Q�M�ܴg#�S]֭�$�	v�����u�N�����	��������积����������q�|gtGgr�2�7�=�n3{��7�+�Q��o��<��y߷���$���9�]����g~k�ӗ�ཬ�#4�z6�Pu����z�]9��.W���ݛt���:��>h"g���Ө�2��_��o6�:_�\Vzؾ9^�,c�f�	��3LG��7�w��{WC^�;�~��=kk�1�l;?:1�E(��;�gc\r������x:+wIn�`��vp�hC[sT �Wѕ��u�ʉ47��������_�^�¯�C���Z;A�ͽ���2�7l�a5�&�)���g;'��D�A�!���+�Mg�ۍT�<�s�W�D+M���*�c\i٬�*��nTY���
�D(�Fv�u>#e��s4��yJ�b��}�j�S�9���/f�ۥ��/w��N�4�{�W��d����	M=�;'��]�:�jK�_3�yU�yVj |uVs�}H*�.}|u�+��7���9 �U�1Wɩ����-	�ZN�ͮW �L�Ze��7���J��VxQ���ϟX�"�/ҽG-�4���W���&�6b���YÝ1;��Ge��בJD�}E���G�k��/a�J3���y�+z�K�j���$I�f-��Z�ț��d���/A��jh��
��z#��(O�ژH-��f3^Ү����B�(��z�~K�F3�kn*c?}ҧa���xT�ٍ
��,�a1(kE�K��-[u�"TO��_\�=�	p�5G9#(����^8U6�����d��[L��]y�wP�E�j#��s���{|i��O<�9S��Ea�X������`ߣ7�EU�������y�)[�,�I[����*t�-�R6�*i�da�:g/t�~�q;��I���zWj�ҫ�SW�Ⱦ�!v)�兩�V�'��x�	}n��gs��ǯ��4Lf�%�H�P�g�%[��{��)�M9��ߚ�����g��������wg�¢��<�y��`�3X�rn�)���6-E'}��0��=���ᵀ���2�Z�z�τ;�Ұ_�c�M&w��WVz���:wA�S�κ���!���V��&S(��.N����s�YM�6[%Zd�=�@��^&���[���C�eW�D��/�!'Fa昺ڶ�dkf� ���`o)��w�W �S�3�'k?x������9Q���\r��gT��]Ȭ��#��mGr���{q]e62��űyXW^��Û�����cw�GߣޏBI�%��/��MY4���w���"��M�8�k�6�!Z�o�F�亮u�srcT�ܾC(�:�_<hd�ŧ���/KU|�o#���Z��M��1�R8�� t���ڴ���˷�q�U�Q�V�_f���k��i��(�xEDŪ>34��E�d�س���0���a��E�W�K��N����G?4�>`\��rw��"�z�+�9�z�;k� ��*�
j�_������f���<��
�ai�X��g5 �f��--���vʼw����B%eۥ�{d�<�329�3��=���B���DG��8�E������\���"bd�1Vo�k����y�if�!4�*x���֘Tc�p
���ōm�%Y���^{B$�2�	ᙎ�4�h�aׁ�L��{5�u�����H-�"b��h�x�;�����7�=��t&o��WO���Z�8I4��ص���α���1�B�w����ۯϔ�!d���ot�8F֟��xS��ҡ�N�Cn�C�^�}�ȯ?f~�{)�*qhRө�\ӓ7�Fʙ�ʹ��Zm6�"����S��(ơt��j�Fd�}z^�f�	_���D%����1�d�� ��`�Kww�[��X	�.	D>»"����	[�4�r�q��-=�u�lwkc�'65�3yT;�e-�����e�"�I4�'w�il�:T�J��0PR�c��p��IǱ����7.��=�E��̢�;�n�p��U��bT�􋳥�:8D�(��
'y���q�m3����u�u_
$?<}ӆTP�k�@�
���!��Y�O�?%��߾��g�:5���U3�ɘ�8�l�ܣG\ڵ��}�47^�����-g��Ku׵�p�)�t�+x�����j	~�DG��E��H���x~�H��\u:1W��rOF��:u�h�1<r�Zf������b�i^�g��s�ž�WAj|��xv�=Ŏ�Dw�gh�Fc���7g\��a���E�>�id>anN�R���^g0���f�E������ʨE�PZ�U/6�t��X�7��u>#�`ߣL�}*���Q�:�C-f���X�n#��Q��dOTƋsE��.{e�l�(Ӂ�霜������r~��ʕ���7"��/ei�]y����N֍�����7�v�k_�k�O��j�ɏ�0���=��8�u�B�=%�fI?���ꪆ��T���ߍ�fI�=��;9:�E�5�3���.QFa2��M���}xpC��P�m$�[���5�('8�7a]f'Vfh\�7R���s��,In9�ݣVú�[	FW[�����[�#`�U����̉<6Y���׆Mco��z�cb�:��xx�=�o8�/+qv0j�#W$�2R�,t��Oq�T��u�k_�ixGI<}3���1_�p�:�`v�%�aU��+�����T������V��y�>fQ:���H��\��^\ƩU�O+ҭ}�l��*�h��(q�:ʘʝ��/��)9�=�D�6�o>�����0�=U�Wн�H��J���)9�SW}l�������mBbˊɷ\]<`�_ȁ���z2����"O<�����K'\�V��
�F��ϑɒJ���H����j܉U�̌!��n���3��7t��Dƹ��j�c6ckZ�4j���gDd13@Bz�����o���qB*�3z�F�^�w��m�ӽ�{
9�j�b�7�Ok��f��2�~��5t��۷�ǭ���1���'V��f�K'�_��u.�J�&�#��<;�+5�-!�P�jL	����Zf����(��3y�r��n�.�]�N��MΌK2w8~�g ���G����9�n�Hʳ0�G��q4�*)[��s��)3����
�>�&n+�N�m^jj�h�Di����DPy�y���6u<9x��{F��� f��z�Jd�o�T")g|Lf��J�\���n�nA��Es�{��8��q_<r��Q�/u�7\ ��-JJ�T�YW�5a皑u�=��@��j�=�L�3iLwz��^\�hD�u+O)k�݀�.��Ҧe^N�����h�B�:�K	����\�k���Z_J�m�.t��K��eKCGi�I�F����x�|
{ާR��X�&������kC�9�o��MB8��d�,�:�1�O�Gwb�V��������#RV�Uḷo��U�=��L��dn3�q��C��W׬P1Sj[���������%�=0�Gjki6�OJ�)���1���Vm9Iv�I�'��JHB��b�*��s��KJ�՛#@�0e$x��qr�yY�$sV�qen�/4�+��1�Dyz��뾩ͳ+e������a��2�	�)y��O\���/{��	����]�D�v�X!7{�2��+6K��V�Ԭ8��Z��%�xksT]���u�I]V\O��fV)h�W�MQ�m���յ�3{�ŗz[86P�]x�gϼ��ٽ���p ���L�W�2(���)2v��D��ݻ�Y1F���1Kv:&[Cc��D�5:%N��䕱�9�ג��Φ)D��,����y�Z&h빌���Wm�T�#�⑚���י^���ӱn�h�.�`�Ǵ���%Fjs����=@�:{�	,�ɰ��ȸy$=Lm�.��RR�[v��Շ!u��w�u�:�c����^C-ABȩW��Vyu�qN�/e-g�b�c'&�+����9��ٽ��:�`��BJD���֔��N�1@YnO�������.z���C|*��#�KB=]���z�(�Uz�9�i�U�.��!/��VaDd��+Me�Y4�����,WZfmw!&�n�,�:�s�F_�B����c^F�c~���u�t\|�&6J��F���g
�R�Z�������b+�Zz-��M;Uw/#e��rM'~��5
�_<ي:(��:���dGY[�%��/j~����V��L��X��s���礕&�j|��{ ��ۚ;�>�T�ux2��,�������7���睫043���-rl�ɗ�M���Gۥv!��N�&ܖ�wp��PK���D&��/���ݘUP�fi)�Ѭs)D�>���\!Fk�BuUVs����^��ͣf���xq-�c��&�]�6���q��F�GE��MF�у�Vcn��vɋ�hq� ؉G �D^ޡv�����*�@��ˎUbzˌy��:�UH������7�2E[���5H��]b��e`�pTg>�֖>wd��I���oac�un�E����m�����oԏ�v��m��Mk�X=]6v��+�5�'1]Iw	�F�J�e�
�ᬦn��ד{�7�����8��o�z=�z �PJ���=�#��b)*��mr��F�2�
-����Qe7�FqHSMvg"�p4\i�3(Ȏ��%�\���͂{Q*��dv�7�����_�h.2�ٹ�罷5B�F{�'�5;e�>�q�z2�導:��:1�5� �]�.��7sU� ��W����R(Ll�Ax��J9`�U'��b�����&�6���́�ֺ��
iJ0��Fߤ5ޏ��5�ߦ�>w��杬�:�juK j��̮���:��u��R!=�[W�����)ɗ�)����	�;l,q1�R�eW�G��2X��q��p�G,��d
'�UgC�Ng��	�U3�+}c*�rGFD��6�s��z*NM�LV���q�ē垃�6�	�9ͥ[���Oj�^�`��a�^|9(����s� ��Q��b�e��i�x�NwS?
�SWg��{��=�Į��y�L�Yb+9V�SH���Vyln�i���zUcy�Q�G�4�ו�$�A�j���*u�pZЬc�K�l���!��?��v��)������*�kJ����m]~�O�Ny���;��}8���۶����pBBۺ�gqL9�Bݡ�iS��H%~�����i�F��2at�q���c7��vr�b��Y.h:�{�iמ���t蔚 ���-+�Q��@����j�gF�!n����]f��s�l�@&�I���+bf�5\,���2H���H�`�T�>���nj)�xj�+,uA}�z��W'�p6c6h�Z�4
����t#/U8j�WT2R�Ao*�v %9맚���/��kc�����`�N�7���^4ټ���e�����OT*�9�ڿS�����ގ��,xO"�7cqnV��d��(t��Lq���U��,J��r zdV�+W#�g h�_����Ěed]���P�vՈxX�v�w7HF�HۓF����g[5Ҙ�c1��p��j"�Y/�B��Ĵ"�/W�S�J&9�ǐ��g��F� �� \n�R.�vU�Fc����j�`S�6������94ٺڶ���ƪ6��8{\ձ���Z6�#]�
�tS�0"�����
���ew���4��^Z�w��M��� �"� ���g�+kD��?:^�I9-b�ZsvQ����ve�*.I7��a�7*Y�:���J��)� �#iɵgA�@՜��7NZ���u��R���G�ڂ��[4?@�"(�q�T����Ʋ��O�Z��r7*�X����"�8ڇ�R�	3��jI�
ƶ+x�Q�i��s�:Txzk��_��%�.�J��ap��Ԉh^�F�WM9V�6��]B"C����(���⋂�M�3>B]u-��ka�}��y](����*v%���Z��q��[t5�.VI�9�36�c��ʉu�if���@��%�??�ez׆d.���#�s����VK��EQ�i�{WV&jK�Z�a���wFW`ĸ�M�r�7P��c��(�Yò���Fs����D�úU��,A�T�m^<���j��`z��:�2�����\R	�'��꾄o�v�u��@�b0ld9S�ǂ$�<���MS�-�TOq���i�{6j�B� ��^~����kɷ��{ރU����P�N�F���BX�m��qV��������E���t�ӏn���3'nGS#YW\t���.�J�,s�Tq�}˻��.Ά��Q7u�	�f����:���gi��}21���$�t��j�7�Y�ղ%˺��ke##�c)�"�:Vl<�iI{�'?��ވ�KS,��`�F�sۃ=sF6�FAo���Y�)y{P�2�N
'ᾓk���E,��q0H�z')��O�R }��+{�DT�I�Xl$9����Ny"���W���ق����ij��Ş>m��^!�4��!�m��z�x!g�2,��CH����q'��q7�{;ٲf�j�D��:^�ł4�!���R�JR�����^�4t�Cئ�+�%�W@0�gަ��~��B4���3�A�l�cdBȞ�/��)�z����ot{^�$��ZC_<.S�y;)�c�O�������4Oh7L�劏Ved���ǐ�H�H]3R��P���b����ATP�[N�n��;�aX��%�B�� ������%��S�C8E5��?]@�Ӈ�q���ˬ�!����O<�������W��=�r7	���S����t}�w
\Ý� ߺ&��Rg�7
a���Gx��9��Ƶx�C־�������ow,FG���k�8�E��y�=i��W�y�+�]�����n��ҀZ��y�W��F���J6��{�������(�W��������~~�t��5�~�ݶEj���ؑ�Ȣ4Ƶ7u�.8��r�yԏj�
>:F�O�P��Q*L����ޮl&�a�������!<��Zx����E��r�=�2��xڎYwQ�^;W�|��9�m�I��\�0E�c���c��k<�����Y[�/k�!9��Y,TC:G����☵ֳ�f-;};st3�����4p�3_ob�U�Gy�U�!��:�x�%k��u-��UC�;�eb�pb��E
Jb��\8�)R�j���F�/c�h�٭q�g,�u�"�ejj��6���[������c.�7i=�
� ��M��֖]�MW���}�Sԕ��qz�!���Q=��v��f�;K�*�v�C!���b�F2��U�w9��f����]��?jNJ��� ��պ��\��c̛P��`(=���P[NJl�ng �a���Dt�$:0���:�����α�/�%��7�(Kv�D�i�I���Tc{sޗB��&����n,��]�v4`+�Y1-��!��仔�d�%	%�.w�Y�efRFR��͎泹P���FiǺ����NR�}�����.Ṷ��:�D�.�Վ�ҏ<olҦ���X��
�^eEX�f�p6��5�V�@�}�)�9p���r=s�ogM	^ks�r��M��5i5�?�S�Vgjk�MZ6��WV�l�K��,�'Ӷ�F鬌�
�u��,BN��������ioo[1_dx�m*!�v3��4��,,$�\���]k	����ԝ�BT'>���mwm`6�m��ݗ�d���@fZ��jv��ux$YY%7J;�J�c���"R�Mɠ�����g�I?�M�����T��n۵Jqx*�4U�܅�4.1�^v�g ��8�d3�'�ȡs�$�<x����q�����jH��<5g��M��R��ʦH�0��zB��s�aF�¡ۘ��Ʉ֍�G.t)0ll���q4�N����N)̛E����]��6Kss!vkr^<��<u�H��93��6�Ѹ������$wF�DJ#�<���e։3I1��S�{G����k�-{�U���Z�!�i/���	2��7Ie�N7�UW�M.�{xt���%1�k�] |��([cI�@�+zd�JE���8ty$�0�ְϤ���bk%���'��!R����A����k\�XǋH9���fz�50d�����W�$�5��rT����H\��_�r�'��y�=�n]��5�tv}���'H�_X!O�B�{m����M�9TC�[0�!ǈ�_q�|P1����۔Id�G�1g�ʈ��W����>�:nr�����I�NE��g����2�4�G��^��A5Ծ
�H?�a`,xz�a4��_ۃ�ߒ*�(���5F��]p��I$=�=�A!�H���g��ut�s��P�Gr?�s�F;gS��sBI?�L	�Q�	���Od����P�Kw$p��f�JΩ�mnH;�r/����{�;ݞ�E��Ӧ�z}Ǝ��1�2gj�B-Y��8����ȭ�pm}~�1�;���Vt��v������o�ᦸ�!u�m-7Hm��Y����#N�)k,.zo���&!��������t*R椑�𷫈B����Π.���T�Cʄz��n_{Y��{�b$x�0J���Z��XM8��ԑ`D��3�SO��reLQ0�M���s3}��^��`h�y�
��W0ǖ�ƿ�#MB
TfY7{�����݈��N�a�L��(U�sێ�z:���@�FY��	��]�,F�#.����"x�}��]<���W�eP��r�w ��zy`3Q8	�{*x݂yJW�R>&��9�<q�m;��n��h��j��RІX�8E�[�/��D@->K2��jҢ0�X��3�h~c�ҳ�b`�&�G�z�s���#���?_"FjÓ�-$t~�ɕ����Ȭ^�0�,W�vo�"b�f8b�8�\Te�N"oV�R�x�>.����e���{ƞ:V��כDB��lQ����O!�԰�8a��K�z����$�Ci�H6�x���B�ޛ����:��~r��G�>�4l�$��Ƈji|pޡ~��{�߿>�/>�oљ>���U���=���j�7&C�I�[�	%�jWs.}A?1�X���ɥ��+��s��w������O��{}�o<�����������^?��������`�רO�TȽ�'=m�8�+��Q�{O#rK��ⱀ�d.C5�&Iӷ1D�͹(X)��J����I�e�~�͝��e�_�:t4F��B/���:U������"6}9ᜫ��	x�U�$���8�S��O��zРl�ZB�i�#}�+�;G�3�����_$��b${��p��8�9���ݙ}�-��?a@j�Xx�g��b�����v�	
��#U/j!�^�ʁ7�A��_+`ƽ�X���m������e�s�S����70+$E�֋�>Ha�Q��*����8֯Hz�.��x��S/R��.h�B�X�F�_��O�����	]\0�4 �B�u�����|���*}_}����~���戮Kh+�=�������KB�|�*q�V-�e�3���81��8wI(��u�jF��˙Idx����Q|��쉻1f��{� +��ޏ@Q�6��~�U�$�HNXH6v��<G�٥��=���_{��?Ŝ��~c�G�hQ��$l�ݨ��{^=��6F]�(��F�,�Aabi����u]�uQ�����q�|[�ϯ;��~~?<�ߚ�9����[O�^l���!���k �g �'V��^w���F��"F~�o�a�r�,���.XYd2��5�⪁��[X�B�?��/>����7A�d�,ۗ*`�9���3
Nձ��
Ĥl\�Ǘ�.-���m��5�� J������eg^����\�l	��|�gk<GX_q�����V�"�!U�[��)*�^��B�����iyp%'7�*��%�͟L�1m9�ao:6��)5G�E&���$�.	~�G��H��Nn2zfD���eGO�=y����)A ~ܯv�곝���N��P��>za��2������Uޘ�^�?Q�奬xv�a4ff�y����N�u�/�2cf/���j�d�G�j$g$l��ҙ7���y�"�)�|p�st�f%��͸׽$���߆,lu	��>�0���P���ՔW;�emf��П����4��O��n�XwL����n�׫�x� �tb����IV��]��ƪ.�>"���	s�����Mܫ��V�߈F���b��lØ��ZЋjUT��.L���z�b��5�mD�VmG�۽�����润���kڏ�=�O��4%z2�{j�sj�]�ZG����g.A&^�]ĺAq&�q�]�*�S8p�JV�%/��DzxSJ&~&�hTg����ŝ<�V�FK~$�3���<h�?p�������~daPc�^�����3����x�E�������z~�вVT�������^�a!����c��Lq~B ��o�m;�n���B=� ג~C�⢫� ���x�Vw��au^����,���=.��<.�0��wV�3���SB��>DU.�3�VE��ꢬ��"�B�e�\gr��3��s<)NL7P�6\�P4��K!CO�=R�����/�@�x��\�'��^���<��K���oT�O���<�����z�{��ny��g�ڃ3,����d�#7�4�51F�Z5���:W箁���M��Ŧ���n��zЋ5�p2U�c��j؎�5��� �=��E�ۯ�&o���*�3��Q��Td�:3�<�_��������}�̫���Sߟx\�_j����o�N��B=�:l�l�� �/��bΟ6������,���E�}b�*n��aP�N��Z�q����I�6~�@���:t4F�E���LM��ݟ]+��x�B�O*�	������R�uoQ,��_�^3U ��ٍ�"{X��+��^�]�3��	��I4~ؚC�yᔙ�!�k8���]��7����#9
�� �%fjOS��_z��7k�x�b�Ku}WLa�Djy�M��������e\
�.N�}qp��%^(ՙOb��Wţ3��M�)3��.���k��:�\�t=;A*q�&g���s���Ç�����￷E�����ׇ׻��?1���Z��_�0:��n����*�>Ha��f*.�V�)��)�4�fE�Y��!{�XZ�Z��6��$0ЋA�3f{ރ�����ݭ\;�A�Q&���������im�����5�s:��EUP��W��F��>b��Ϳ^�#�q�g��\��G�a
>/�5z�����P[�כ�8�^>���hu�(��7��Ht��؁2qz*����㜆�M>_S��ˏE��7��=�ٻH'�w�y�Mx�\EJb�=.�<��*����۷�������$�1�H�ő���a���>*ك����s���Z�
��IN��|�5=Z���[wwsO�fۻ�*���QB�,s����\���R-��`z��?�������l��W&~���bt];���T��R�an
Y;/|��#{^�-x�5����D��)_u�B��[{����m
:}>����N��EV?�"����������"�=#�6��-�f�/ˈ���xs7�ˡ���6i.$����2�LF��:�]5_Z��e����'����=<��H�_y�b/l�0�[��\�f��}��)Q��:��?Q!��,xu�Mi&�l�W�?p��3X�(��?Uc�I!�Y����Ѭ��(x��#b�Y�x�_$��e߬��0_l�UC���E�.�������deҝ4U������ݙ�=?}IxX�O��a5��L�+��k%���N��ficcfV���b�I�B4����ʗ�p�Y�����F�24/��컼�����o�N1�^���U�/JJ�`�.�F��Yg^����i�:�.��3w�#�xd ��:���t��{wQ��}2�dN�_���n�;�;�Ǩ�7H��*[��Os�3{���9�59OAѤU���ѵ��Y-4�{A=�zxj:�*r#[�n}�6�V0ƃ�U�C��\;z�c��ޭ�bhD�D���Q�&��B-�����W��peX�w|�Ƴ` ����9�;&ǙK^��]_diR���$ �k77^�i�a��j�Vj�=[+	���4�e���;(#X���9o�'�o
/z�8�v1n�����"R��RoX����n3KYh�3B0Hr%}uoC7�+��)G1���;s�ww	��Dt�]��3��g�(w�i�-�Ɓ�ˢPW5����N�%�T���ssO(+,j8�9g�]������E宰8�L�$�ݮ���.�5y��䴨m���Xw�-r
����sx�:+p�D]�Gz��"�h;�?s�;cq��,s�b���dK}�����C̺�����~38�#�M�yj�k���ӹ��,˻X %���z3x:C5��Gn�˳�>���nHfV]�K.Q�r��Q�ƒZ���R��҇KȚ
4��>v�r��o/-��I0�-�$���u[F�L+�BQ\bk�s�^"��J����FV�		���LU�2:����/%M��h�s�̊�h��(�NE5��ѭ�v�<���(&mrW��yL��� aM��S�!���˅�hf��n9r<F��x�x)�;C�IZu�]
O��*����r�e�vL���$�Q-�t-��v�y��jD^B��x�!e�A�;��dSqh�:�³��*�&��Ud�x�I[�����3��u����\�f�Frqɷe��"�gY-Οê��������Wwϯ�����>G���������|nc�\�}cٲL�����ʍ�d�X�@�7�C���.C��c/���vX����K�$���t�M�G�b>B��m_�OU{��G�H{#H��Z��.��=���'�*N�J�ǩeu�W.Z�w��~#����7FKzG�µ��f�UF�33��UD����dK�g�_ι�!�R'�aͺ�Uo�k{C>:Fz��$q���<a��B7+�W$�=1Ӓ�=�3.�C���Y�qr��Ýe��\��\Y���#���ȑ�ׇ�^��s�����i��zj=�ǃ3bJ���%�c9���&m��	�u��H5���({ݑk'��f�BX� R��x�|�n�G���Dq�!�Λ:~uE����0�ah�;W3`Y���V��K��eWըY��v'�T_�]���|G��0�.
\���c�����E9sXc�g�I�P�E$�����t��ޓO�Z�]�ς����bF�$�FR�H�C:��v{﷘z�ˍP#V�Q�32����53\�	�O6�b*~uӜ�h_�;���"�ٶX���c��Uy}�,��C�㶨��x�2��il`B-@��Q=����xxz��K&�3��Q~ɉz���Rdĩ�U���ѽͽ�#����wIF�,3�q~S�'q�����~Q�?1���/�F<v��1���m՗���3��R�����Vʴ�6�[�
V�ѹKq[3y�{c� T��oW���[-7�3�	sm4��V�q���D2��dξ�پ�3P�S�C�o�$��=��0ʷ.���Jj񔧲�����*��t'��Y��>�rob��6�2nzP�S��=� t[��E�k�0��^�r�/*`�U�q�lGg�}|�C��g�~��}���l����_x�j�Qo���Z�w�L��.��`���KH��0��1��b��h�!��c����/��ق̵��>�kI�U�$�䍤s�fG�j�oo����F2c��XA#N�/����%����X�P�$�k�_.C8$~���?��@}������Tt����N}�]�q;f��q��cz�lݼ�yL���yOu̠�*�2�J��}%���el�E�'n��-&��Dx�M2������u֧z����GM,����]s��~�%
R��S�����Ү�[-�{X1se|i�6��������<ǋ�[���_����=���LJ���H�α9n�K�ww��Mj-�L�ꉡp���0jdV%�qBk�ո�e��o����E��xG����H�.��-nm��rz�@��Q���,�K�5��=c��k��`\)�$V��"$�qc͘ekˈ�ν�K�&Կ__�92�Yať����:Cyq�Y�tv_�;}��=ܾ�*D��	#k����_C��R����� ��,�d��^����/d�����1V=���-�d�ڛ�XN^�1��J��x�U�Ȓ�{����[Mz��X�}�m�h ~�|N,;�1�+
���{�2�W��O7q�1W�&_ǳ	$����hʄ������=m�1�t��#�g�A����)J��P�m�����L����:W���#"�I�����ã��i��9,�ϔ����c\w�m���ů��v�.��k�8����>�b$�0P�8ч/֦#��ff2��LKv/������!$9�j����fy�6|j��������"���Ѧ��h�nS�+��`��6t�(V������wM�'+�VH���o�1�,�c�I������/�wYd5���拏�Z:�R8��1!GNj���9^<r��0<��2�{L�ء�f�e-Q���p+��=-5����:��g5|���,��	H���9�\~���<<�C���y<j֗�Cƈ�C�s�����s��=�ǹP��ԔÙ�B�ʒ7��o��wf�g��/�t�#"�>�$�O�2�U��t>�ȣ�n?���Oq9Yf/��.́�eݳ��4BHM}氓���;9��q�������e��gBA
XC��B�1C�u\��A�ص!9Ӿ�1R�n��(�$��0P�d�0�凍�I]YR��k��|&�A����t�
�)`�1��Y��:������Q��z�||q�O~�ʫ���S����6�/Ȼ���ڪ[���Zvh�X]����o-�%_U���-���a/��٩�#<�@8��Dܛ�Z��oW�Dz=re�q3�0�z�c����l��a~���k��C����Q��=K�g)8�����G��#p!g+����5��k6�l�5?2��:`и��Tݱ]���ʂE���Ĉ���+��qn���Q3ƢvE����8F���'�_����>S��=��|�%�=|=l���\7@l\�
�Ѹ3j����Rfgg�*꡺In*�m����R�6�Z��oA�QgG�Z�~��7�~���k�����H� ����Ҿ����(y��uHX���go����h�F�Y"ͮnZw�Pne���_�"5|�ԇ=�N?����#�BU�Ŝ��?1b��43�
ϚHq�Xn�ЦՎ7��K(�˘EqVE��ѡj]�7,Z���o��������on�����dՉ	����ٺ˩s
dT�ۮ�co�3/��aۖ]ť�Su��Pt��l�$e�f��{*�`�}j�������՘�H-Z��kk7�O%���e �g�q�`�ː�O�D"Br���nxh���H���q�=xE3�(p��&�
ۧ����F��������=F�������O���3r�ᆏ���J CG�NBR�4�&%���ޣ|;Q		]u�=	Qv��F:��rz���*-��{Ȟ�����]�������޵���>�[��.��{�z&t˧�^;k�y����d��/�X/�]0:?���*~
3�V�]��L	]���g�;V��>��Z[a��Oj�NV\��N�YΒ۸��Q�t�G�ނ�i�#k��Ld�*�?��:>�?�̗�q�.��%�����ڳ�
�s� �P�[��0V��)ݾ�̗]���<]���8I�+8;w/.���18��XhTt>�_Q&�Ό1!���x��6Ϫ�_�x�p��?]/���Ha���xgJ�{�z�$����kE�a�+��t;|/�Ϳ�xO�� Z�=u7�Mxᗽ>�@�N��=���*��E��3E��ݥ[J���3����r��>�}}�TW���$���j��~A����6��L�_���$>w�KϘ�D�9����Ňʏ����"5�S�㷕cq7f-r-��u�"�3�.�>[X��n���Ԯ]���P��x��;J�Y1K�H�6V�!����r%/ވ�z8�{ZmOOΡB�*jz`��$Ϻ�"ΐ��X�����w�� �aW,�F���t���:�1׭�s�1Y�sN!��"�0�-8g����ʬ�T��zqϚ����ѿ��~����F�
ZM׺������X�vf\��Qz���U�LZ��M�㬒��m�<G|E�rs�D�:ZC�xt�ޥo���p�͑Gr�Ԇ���ƽf�α�D~�?GׄR�p6��0R�GO�����r���I��zJkH�ZO]ϓB�m!�VX6p���앗�����I�d��'qq�C����^��*���f��r3��
��
�9��񑑥��3N;I��JB�ɻQ�V�Z���yRdɆ+[W���'|;eGػkw����n���tmVe�玕��`�*�];zQ�u����ñ=I�W�D�G�q<t�%e8�ld���$�srb|X�b�Y�Ũdk�N&�R	ܘQw����]�Ӂ�a�Y��)�l�h�l���jʽ/�dėo�WT�)v���f�C�aas�c���̸���cW�sk�9i�ӣ��_=�!�c�<9mj�,����^;\U��A�x�رG�Fg:|ĮWpD�oP�G+h! y�f<�KV��)-J����Tڌ�a���B�T�Yˮմ��a�wQk�2�����ɷsK�~{���+@���)G��fm�
�8���|ӄ�����Wq=-�=�D���CmV�둊���n��GE��x_Y��RI�c%%��d+o .��N�B�+rf�54�y/!����u��CY��̇����{eMXV�n�K!T�#�}iLo���f�����ah{l��i���K�g9ڧsn�.u��h&��)�;A��A;;<����odR�v�1�p��^�q�Sv�	��VC��C·`-g�ݨ�|#�w�t�:J�:=A&�9�b���q^t�O�ܰ;��A����_#���f0�˓����vE8���V�:�e5�G)\�k�����"!;뾚�l�K�E<���6%.�Jy$�`ǡ�-��=z��3s�j*<���FB��Fr�Fї��ٱ<�s�h�&�2O!E昈NJ�TZ�W(�ʇB�&u�/3�5a5�KǊq5<s�]snapIW1W��;�ɸ��9��UEUq"6&W�F�q�)�����;B<$$�3�3�\�
��3�9]�1�3b����H[e��̛�����rJ�WT��*�4*�����Z �
��֛-�AC�(�3!qRD?'������~���|�{���ϝ@9p��W��lJi�J�6Q�COd���}����P��CAl�t�(�|��K]j`c��so�o�-5��NML9�`�CW�DA�a�s���ٷ��ϋ?x���4kq��4��<�}��E؛��4\^..����9q��Y$�=o��Uٷ�}�!z�%|��0+�my�:B�0���6�{��Q�C)�0��iB8�0G��#.��}�,Tt��B*+i��~�]�	?��1,���g��Z��,_9W�L4��D*_{��A�GN���<�s�&��}U�����z�&�,�7Hy���ʀ��^���a�L	���:�U��%LR��W��W�G�d����xXd���n%�J��5SWF�X�m�ᧅ^Sܧ$��V�/���ۇal5��y�d��p����~��R��b��͑�"�y�kA��,��q+#�;���*�w��?d�ӆ�ߌ��l�@/S�_lR���BXA�H�1��A�3��z��\)*��7�,��b;�c�������Xg�f�B8����<�����&^�>���ٜ��0�B����PK�����"Λ�=k�N�E�*D�6t��:��L�f����� �
�ު?�ZE����Z�/�̅��^��������ψ�$u������>cbE~XtR:�2��Ƒ���D���q�^.��(J\t�(��HY�}��˯]�*����R����՚�D:��Au<�Lf�	�k������)!{�5ms�47�73u�fKS	�I\�&'��z����);1a݉t���m��N��'?�W�T��c����I�~53S�����Gs��U\�۽����ka�<��i&��4�0����3RJڒ�{���g鬝 �c����X���cǕ�M�y����s����S�
C_=6x�����#7�>�6����$u+����D�.6����X���ٯT-��ʆ���5��[�i
�sq�&�E�6au����w��Y�;��5qw��>4�O1�\l�PXG���o�}�!���]�x��Q&�bC_=79#J�}}��q�ֿ�\�8~�\`�jZ�!J$0�"i�+�����}gI3ɪ,w�E�a�Eb���|�?�5Z�{W<+>l,���:N��IT�����dl۳��,^�p�w/P�]=��[�G})S��e@�AY[�Ob/���Z@����k؉�8���u�a�4/z}��ӿ
��m���{��Ĵ�����?9�^Ts�Qc�1qU��ח�rɲ(� �0�!�ߋ�}��۳�{��Y����t��0�o������4\��w�X$ԥ]*p�u˵.j|ULH���S�f)�H`�H�����.r�� �/<h[a�E��:EL`H�k�/}~�S�1x�)�Dx���QӇ�0eqấ:�1μ\+3���ύA�x�b�
����:����F��a&ϵ}��M413|���;^���Q>��aG<B�N={�,Z��c�!���&�����@`��u���ucF�G�1}���\���- ��;-�9�[��f�G�0	�]��B72�y��/r���q�JV������nL���8��C��k�r�H-A�JC�⢳������s܇E�l
V}10����b�?�T����{=��։���\E��\.B�n!�G�B��\��z�?�J��"H�A������J�s��U��P���s�D��鎘�Aj��∻`cˏ��Zu|��y��h��X�p���P�
l�/Ez��ɶZ���i�~�C���D| ���Du�˧wW�#����6����ј���9��F��+D�B~��ە�����<��l�C㜑���d?���������W��L(x;�񇈽F��y�4�(�;�Q����~��e�f�ݎW�����<��l�	:����n��B�[Yb���kԳ� #�j�v�].�q�H�9Y���0 �.;1��xk��A���]��I��,H���ET�O�Qʶ�8_��S���q�R����	�@���i&��6F)��5H����1�����1|��<V�U��6,�}���}U���񔙫C��-�!�?�x���Q���g�gև�e@�5��l�Ď
@/S�D���W�4�l���[�s�	�����a�Ls6���C��V���3��CdyYW.��M	V/8W���P뾨�]!�_i���#��Ƥ,�<�Շ]Um�������Z�S��Ț���
���?~r�}/�U&<����?{�nݻy]Ѡ�q��-.�.�)�����gsY��ա�[ۥ��B���#���:�5���	��ՎF���G2� ���T~D_-"�jx�#��g8�T���{Rh�x�!渎$�TzY�C��Tt�K�-�_����]+��P�HHCuy.7KŋCl�G���Jp9*�0Y���:C��@�ZZC��j4���iބ�����}ط��t
�)K�r�+�I@�ʊ���[�>�{+ev�G����x<�|_�=��Ϙ��zp��~�^�9M�U�r	ks�/�BΝ"����#���ezv����/�%��u8gc�K��5ߊ��=��%I���P<-�,��J��@~B9=���'�!��mvx`����V�$��sq�Ț�B�s�������j*��6��^m��Q[jo�|H�T���������(���/^�{;�L���'^9��]�Y�&�b3c����N��)���܄^]���:/�.,_^$�H�A�T5�����*�ڭb��y�E�&���I~z߷ܳ��6�6t}.'ݴgA����l�T1T s'�M��,4�G�>_&��{�B��x��AV�fz�ؽ��G[j|��9��?0���L&�p���˽���!�z��!���$ᤅzl��܏!�_L�O�c���La6aG�4p��5�t�+���� ����=t��R��0���I^`",���e߼�
8z����l��<�(F�dQ%u�~Wa!o׽��P���|�A�Z|x�CI0dɟo��~J�6G�΃ǯ"x�Sͯ������TV?(�+)�J��d���=��9�똷I5&��d,m��&S��,����/t��i(�a��@�1�M#�Ċ�y�:p��\w�HŞ�f�/�m���Bz�~⼀�[Ҏ������{U�~dYBcMUҰߪ���q�e����Ŋ�q��ƴ�Q��N={�$<]�5�ݦ���ޖ,��Ɨ�C�Y�ܴRCkR�<c��M?o{�a^���kX�gp�B��GM�a��U�/{~�.	v��ZD:K_g��Oq	�e]�w����������3�_$/9�O/���c�x��8��mv�ûO���"�[�>v�:��9R��2���'��cy=K�r,4"l��F�#����c=1Aw���_��Z��������9S�/j��D]"	�iњ��m�JYr:�WyI3Q{��<�lbmR�����&H9��rg��y�\������c>��:��
w�"��e�u!�Z$C�y圸�h�Z��Ʋ�Iy��I=v�Ć����4�V�B���y��*�K�%�_^,~�_�{nM.��z�'�CM��g���:�VGy(hC�p��?�nL<~�>�q��^���}�x�F�~�ح�E�����h^����������@���$������~^�Cn����xF��Dz(F�
�<_!@�[ώ��~^e����-wy��P�Y,����=~b;zy�2��ͳ�s��DC�Y�>y�k��|e��.�?2��L���{���Aד��N�)��/c������ �ۢw9�i�rA׷*��ل�h����7Z���y�,�˃���}Y��\VV���#?l�s�6w^��m����n��q��������A���	����+3���'�r&�|0|)^�K���\�y�C����=�sŀ��J��7�����ҥ��"�����-kU� 
E�o-j�z�z��䧓�EbR�w+t�����Ig1[��n��������Lxmi��:�-함Í�Υ�κ�3s��Uq/bnQhڝCs5M�M�7j���N��R�u��V8��0�����Fu� ���t����70wrR�^SD\���؟"��]O�����e�Jx�cv]��d���6�Ǘ�;׌b�[e#z�Le�7tc����8� 0[|�M��,�#��xn�.��u1I���l�Sh�2������\��u�Un>q�'�*�j�+�!4fMY��f}t��MS!Ҡf^U��v���NC��V%a��m��J.�\�ud"�sO!�K���0�Q���նk�!��§�&��%u�D��[4��[�aSe�)���ɣ�I�y�I*E��� E^cS8�95̘���{&��_�I���d�{djٵ�jE8���b�3	2��X�v�*���p��]�VM�NMMڝ��z7)4��0�$�`EM�4��Ӳ\���U��[M���t%�rU�s'}WSs���0����v8J\�x��t)�!�����������y�rj*�i��U:�r��\ٍ�D��x�2Y�A���D��#7Tm�I9�r�(5�f(T���t�Jj�UsI&��܆j��(�'�ё�KlZ�s�2���-�"�sY�4J��ǈ,���n*W�	��m�n\��͕DxNy.�D�ӫ*��- ��vH�+�
�S5H�m2l֡�v�rL��gw���8��|S���4�T�ç��1�9�#!N^�f�%~)ۊ�u�&2`�D�]a�����U�NXK���f�ݷ���P��C��j�ń1�͖C�3�ef4�۶9�WOơI*ԙs�]����]M�T)���PA4��؟)���N��ڀv�"!�!H�5��e?g��/�a�H���Z@.Ǻ�-��4ՄC��S�_{1!�VH6wPG�q${���;���o��v<��3q��"��a�\Ly ����n��MC�w�C�覣G�It�"� oV�F�a�F�L�P�D��;�>
M���*L����d컭U"�[�<��)NLH�]��64�_i&"�0���U����:!��/�������je��4�y���Z'��[�=.�n5:��*�\�:D�m�d͹��::��LL[�����|��ޱF�x����,yq�Eꊊ�w����%�{�HQ|N�7��7�M#�h9ws_UM�?3�z�"��<���D�/�����{|v^�y��I���8~�Q_��b)��H�[�C���E���3/���kf��Ťx�Ǎ�^-,$�AOk�W=7��͜ U�#�Ϲ{���t��*,��7gf�v��������������VE��=��s��֐�+&֝h#��?#��J�[ά�Uuy�aj��"E�H�������:��׎�B_V^�ϸ�<�"�:I�c��G���+i���#�����v��T�R�#-��4�&�������$*gb��;ֻX��r�i۰A��ܒN9��X=shu��Ϯ�W�LQ�B_!���O{7}�t�Ҹ�Z�y_/��էH�'ʏԵJH/c�ۛ�0��åF����.5������M��h�m���":��`qٌ�)x����a�$i_�R�����`5��~c�S@q����8}����g`X|p����_ޖ������ӓ���R}I{}���>�a��'ᅌCL7�Vz����K�2���}{7�>�&�+������Ɓ�,����$<S{��/׽��bC�QHx��k�r�CHGRΫ.�����Q��=*[	�;1��+;��0�:Y|��jμ�d����'���!�
V4�k/ӱ�k]�J�d�1cPЬr�<���;�/Y"�L�->��o>����c�]�>��D�����R�@�l�*~s7���(��_/����0$/�ϓ�Ob��Y���oV�w��Yl�[��P��AH�	�51�n�Q5�6��pq�b�Ծ�e�țeQ���:�?�_�}�ë���=;0�ٓ��a���Ή����7��I쫬�5{3�ǵv�zW�؋�`����{^��f�aq.ٽy%�O;����5v1���ζ3:���!wzc������ro�ۣ��1��!�ۂ��j�/;/t��ڎ�}��z���/�� �>=���J�NKT�A��k@`Y��&��yӰ�oH���$�7r�z�=5Ƶ�T
mw���������#\�ڵ�h���WA�����ށ�/+
�`��cf�
e����Zzp^�!oU��4t�A{XN�o�Zv�&�l�QV��A� �������xQ��\w
�u�m1���"���[c"�����|�z7�����=5���p\�����Q��U����]�{��T!`��sq�_���T����I�}(ā;H����mQCF�Y�l��fK]	$)�z����*!��
<C�X�]L��x`(f2�J�O���y��d�s
�b�f��J(�Pܭp�������Lԩ/N�0�O'Z#(2�.�e������(�u;8.�S�A"��4�C+g`A9Z
���`QYQ�Qv���'��
�(N.��k�[�Ōw�jnf�>��	^�T̮�]���V-b�Z��P�!�2���Q�N=Ꜧ��H�,�Oן}6��򜿪'�ֵ�;Z,rK��㵥��L]�aƓYj:��<�:{�1P��w�k2�t�?����]4����=l�9o�^U4�[���Љ;E:������h��Nuf����#]�.�T��?	���~����H^�{ Yj����s�S��d�-5�ΙŻO8>d>��a	�9:��q8�Zw�O�l��U�n���q0N\<Ȱ�<=Ȟ��Am�~K7zei�	��֙���V�.H4�8ݴ�W�v�����P�m$C����n��D߄�]�be˷j��eƷ�@��m�Bf]m|S{�?r�	��ώ�[vi愆yq�u�v��7$�&@�V0֮ːY�ŜuXKW��\�lK�[RM�­	ʁ�1�wNǶIrо�JBR(.`�8�+�*y��il�Vb�Kǒ�z�Y1�,���r�;�H��yA���J$&�=gm���r�z���Ei掞�^��1��wmR��w��0��]�;��OWS��R���@��9��rx[�P��d����=ui&@8]p,�D��� �Tf�P���I��D��"����u*��ys�^�'�J{��9	���Ʒ��ߚ�{��;8�i���ΐ��*پ�=�fī��߇��C+G���u��zRD���xQ�P]oT��sJ�B:���<�<آ�s
��f�ozj�q�}�]�Ex9�����j��������r2WO[1��l^`��s��Y1!�<骾�ܧ1O�!�0hN6�?~W�	�(��-{��=�Ȣ��|]��骬�Z���q��ry�F�S��1��<�w5��ܪB�.��ֈ�ӛ�a�_4	yNu(�#f�Z�A��(.5P�r�lU�����c�s�m7����US�p(���H�5�Zǀ�[��-n�1\c盨V��Z����h������Q���v�(><�iI{�'
��K�t�8b�7�O#�i3���}Ud�y(�b����S�GÎƺ1Hےf ���3��x<��;f�Tƻ�E��Q�U)��5�:�qW�*�yV߭��77���J	=�s�;��GFԠ���^�F��<�uL���^�
Y��56E������5Z�nI�
����<o�����z&	�<��f�{5���_g
�����dae}H/�K(.?��1��G�J�yhu)�Y
�q뫃$7@o��Z3u-�iot�]9��o-��s����R�vyL�Y�����NξL<փ52�3��֥�6�y�$HY�uc����.���ӵ�K[���.��&��\Л`��7;�o���{O+�dۣM�\́��4��:T�v��௦6Ү׻�6��88p�rg,<�*9��a���ʖr57�j�fvQ�\֗�����E��rg��,u�U�B�����sO^�k2d�K/����^�ۗ���4>G6X͘y�F��E��2�����N�<��"�����4/w�c�A��ჸ�IbG|�zT�D�ES� :��ڶ������)_c8͏M˫�!�x�ըm7�)L6\W-`��!rr���yOh���Y��,����1l�:�R�����&���Y&R��m����/�bc�*��F��43�W66w!/�[hJ�ֲh�B�+�XC�/�`�̢�U,'�"���S{���rZZo7tփ�kt�p�.��2�K�W�V3��QR�GG�G�E�ұ�)�;p.�9�cK�1�E��4�\픗kC3pn!j�]�[�2R@��&�9|ZZ��-�V��z�͏Z�Sɧ7wN�Z�����y�R�"nG��U] �Zi���o�r���~W|�v����Ã�����փV_X'��$ۚ��v���S�̲ox�]������E���t$h��͖��3�gY2cR����n�`˿�[�%-&ԫ��Y�,H�M�y�Q��Rb�Z�R(���W&�d�j5�%1� �m��&K��������-h��acm�ʺK�j�3ckQ&�*]*����F�r�,M�$�ܩ�l����QJyQft
4�ZȪ�a�kVg#�a�NyHd֋FTh؉�X^'1K\�v�;r��.�Y����Q�3Ȋv�i�lF�btNU�0e1eyY���-�Vd�`�!����z��Y��h���*�-;�����Xu�P��Nۑ��ǒN[{q�6��=L���gy{L�!��á�5YZ28.�w��鸶�8 qw*��$�Z�z�d����T=�	dQ���RO��7.��-�L�8��2UV����}ѧ�:j����:��e��R�ˡ��F]\Ӄ���-����.��V�x<��R�H��<<�"�D��5ȍ��㭎/X%eE��"�7D-�Ca�mNC�_��Fu��c��?ʸ���z�V��T0txV�r����NXs�MU��Yb����&��~��&Aa��
APh�l�y�2�|��t�_$�棉����?-�E�'����$��;7�M\E���kS�ڑe]7E�</�cM�c"��ر2{�ɲk�Ȳ��+�:���o���L듙��Tɠ&�Z0v�@����1b(�%�}g����4�5��u����5Nj�Ìk�{A�bw��š+�����������|L���r�� ���SZ���EY����֑�~�p7'�留��3����D�Ѱ�ꍎ��pwdq�G;U�|vZu�Zwp�k�1����&����TN�;��dd
�n�+:�M@�rA����� 󁹇��U�r��K��z��募q�<.��xv�����^�u.>���-9ǋ���19>n������i|�+��yա*.s=]�r�)�u�9�"@��i��r������h�[����qm���'���W�L.}�-�rW��ZY��U�4g�:�2:��-o�;~Vj��sB����=�U�WW��-��z��C�"�ߙ��N׳��Y*a�%&+n,G`3�N,�kXR���c���zJG�՞�v�k�uZqB��Z�D]\�!Q�o^��/��W� iMω�è�ɚ�����M@[v璋f4\����^�X1�GM?Q�z�i��w�ciS��.�̭� �g�i=b���YT�+oN��8f�Ga��o��HB�,�/�����\����:�%w�N���=)���s�J�Hi`��3������E��/]�g�6��a��1���`�=��[T2����2�oy�wM�d�TCIܷ;��hZ�eB�z W.�l�b�6�G��Ï2�脥���x;�onV�[��˷KF�G�"�Fg,�-0v�j�7'�G��V�k��e��q�+��W-���!�d:��lA6S6Egc`�؍7M��yp�Y��B��T3�8
�2����痊��S,�a��
V���F�HW�X�L.ѹŶ��Xfy�@�w��q�-�jVL���ų}y~����crGFL�8���v�o"�rppn3�N��֘cش��V�t8�A���/��]v��l�S<�j&�2�zc����_;m��4����2q�Кᧂ�b�$�����Y�`[����Mk�G�܆�a
Fm����5�'w�vd$�L'�N7�7!>K���uuʶ�ͻ~��#���$��I�o1�\_����=�=e�r֗��^khLEE���*#��Z��oG<�����sx��������mĢga�a5G�*|o;����[b��1��i\�Y��P#�͞��q��'o#w���,���TG�0v����6ћ�h+�:9Φc�;n���S��xķ��7r�:D��$�¦�ݵ{��L_eѺ]3ku�ɓlL��R�2n8v�j��wwH��ؓ%ō�"�zi�{;����@4�ҷ��y�öK;�H�.6��ZNZ�F����
�td��,�D�[��qr�W���^S)=��nzV_�u]��:�	��w�`�Gb�W5��
-ߖ���<fi�׽0�J��(���{�W��~|/,C��E��b�i����Pƣo�Nvn2���T��Z͚:2�a���Ϲ�d5����j-(��:Q�&�S`��TL���|rMARn1�<.h���s��;�M�V![��O�ߧZ��l{�:��qu�s	�͎��N0$D�$um�@�ƚ��o+�BW;�����R�C�7N��4vK�͹�\n�j�/�$�R��||<3x�z�£�9�C��NTf'{���AJ�M?��[^�M����h������ki�u��k�dc+0�1}�q�Y�A�e���<�� ��G2K�j/oP��Oa���;dg`�:	U����a���gظV�)(�^k���5��&�i��{У���D��I%j�������Flv+Q`�>el|�����:m��x�un��{���,SB��8�mHq��8�ԇ,����>�ૼ����׳+���f�}U3blȻ�&���v���]���4��8�5z�YR��Z�;aǏ����:JNQ9�=�<*�Q{d0r���߳�&�}�w�����2�����h�*��}3}�{YZ'x���}�$P�j{/4�m�W7f�ɺ�2@Tud�t'��e�f�at���@�Gӽx�L(_f�5͚9A��I`� ��I/Op����;�{5=�vv��{�_'���5�%�v�E���~�8��ou��!F���*߰��N~�j���k1)ERmr�){H�l/<�󝆖|��i;;9������n�í��sݚ�rR���17]���WQu��z*��vy̗�m�9K�g���r�qE;9��3O�3�&��+G��޲�|m��ݞe�0>RC�� "Mñ��"z���0�.x*�'��dQ-�˞�uR˚�s��Z;`k�Ai2���׵�P�\�3��"�M&9�5h���`C�7U,O\��]�������O���7���<.ZZl�J]p�x}��z�Oˇ��b� \�Z�>�J�PsK+�C�ڔO>s:��"%�b�t�uC��==�<�֭����Bt���������'�*�<|�Й�2���~����RK�w��IN0>��Iھp��³���Hq�e�B˦)ɚ��mTɘ���Զ��R�����ǋ��Cv��q&'.���2ڷ�so�|��TA�+��e�[DS7;�E�k��I`%�G2��	xn��j�FAz�<?w�ٝD��m��+V����j-�kph��۝k��������d+����[�pߌ.��қ��l��1��/j�Zɨ��JX�	�M��f�Vc�휴y���O������9:�q��1����ƞ.ywn�}\u��a��3gmq�t,�nEw�HU)�3f�v�*��d�L!�'fPq���+\u,Q����k�*����J��c������q辈הb�5�E�z|ޔ�:/uͳ7�������IbAa��ގ��Klw���'��:)2vj�U�'Ȏ�׹���C�sH�2짵u�G\�ݎ�H�Q���|!�'���
�S�@T�$J��>b�q�z�N{�����nԵ�cW5��q�ؗZ�[,0�f�
�2l��D�}�E�ii]o����Gs�sVs��ȪP#g�n���Ԥ'-�
�;8\B^��j�]�L^�z;�LWSu���j�ӭR֠�a�-ɎQ��s�h��=�-\wi��ô�5rb=��e7��F�V#V��uMĮ�v�/'ˤ}t#���MGi)۽���)�T���Ec��y��J�Wn(Uc�iϸ-K���X���#5�:��4.n��[�&y+��͙2�m�g+���+���ֱ;r�\��Z,;�"�[&�V��&YsJ�x��9�G����S
���AZ�(��Y�;����sD���ܪ�[m�Ӡ�գ�7'�:���u*P�c��MTf�[aY^�s���O++ge���ݹݨtb��XV�8�=�N�˻VBIi����d�aX͸�1��Ţ�rV�#��y�"'ʩ$%5C3�aԎe��{�����ۦ�˛5[�d�%#�Y�<Y���>��V ��wn,���O�i=Ʈ&C�t�fd���H�Z����3!����E�m��I��fE�wx��&���|�`���9�+��k�f;�o��p��E��m[���U�KD:J���j�f�lsadh��Z�����a+������׺��n�m�-�2�ͬ��r�P�q�蚷s�Eq̡t��I�yk�D�w0���0>���_lKyW�Z���/&�vV����y� N�3'���&�i�u�x��5Rj3.{��p=��Y��E�8�^����9�5yiTp�7j�בh&h�0VQۀ��\bi���
�u��zx�����64�H���-q�X�sӒ��,iS]}����=(�r礮j��{8ť�{�4:���ɢ����A,υ�3�q>wN�&�ᘣ�׆>�:E�au�T4����*ɀ\�w�u�h�n����Z��a:�3
�� ^晽uA�ǆ4D�7�g�ɻ�\V�އV�1}��v�l'��{� �ȌG.$�k+�t��2Yi�a���a��3Ր�l�z�z�g/�x�����5��dM3x��6�3�Fkг-�wVzt�L6�胂��ft8��fH�������%r�35��z���h��h���T�
M��L&�I�|��< �]�#�\�|"�lsx�ܬ��gH��ei����k���PU��y��/j]1���t}|Ay��i"��z��W�w����ʄL�����������yM�ey�F��v�D�Z���Z��W��(�4F�eOUs�܆�M���l"�q\�vå�cmB�ɸ�j��rY��G	ʶ�m^׵pĒ�*p�)F�3_��|�tyg��9³�?.%Y��B��$C�]��y9��acK����]��%ȥ�f1�0M�v�bu�33�U[(��/b��G15wձ~��G�x�U�@�Q�#`a�O{l����D
w������qq�!��^wF��s ��|�xftI�/��?K���0��B������`)!���y�2Jt1��:�hہ�/�J�xW�G�����%�e�$�V�4�r΍��OSsaL��"���5�We��o�M��S��5"�VL��n���w����uһ:�}�_W�g���0�I�[y���EO�}�Wfc�|P<��,5���.@{\�����Sf鉄�B��Q,<��t�rAXsY��<�\��aR5m\��j#v�0uҦB末{1�� .�F�jgE�ϋ�l�9���U�͂�k|�s�x6(�o�Z8D����Tf�1�w# ��gh�~U:�ZP��{������{�G��/"�]���I�+���	)m=��F�T��i*���)uˑ8J��M�Al.���˷�gru@�Yb�-�p5��.C}6og�B�3���,������{a�ly��=�yi
�"w֞�NaN��:A��ō���_Y��n*�K�j .�%"�1TE/��[��"s%�X�>>O�eW�y"[N���C����8�`�p6��_=��0��;��u2_���yʕ�}�fО�^�pS���@c�V�N�P���;�rS-v��v����&Z�3�N!�9�m���!5��W�Ru�Us9����$׋��)�<�H23D�f�u�nt��t^�tGP=v��k�vWFZz�D��
��w	A*�%��t�����"#�C|^y2���j
W~�$���4*�,����1?�J�.�9�e�;�4�=r�d��^	��ZOء�g
��c�%8(�#-%�S2�Jfzg��Ҭ$U�/�������fF��y�We����U��<
�ng���5{n^�l
|�h���z��^�Aa���v(�x�8�����CƦR�c2���՝2������+b�'8&3�v���/a[T�G��+"Y����6/>}�?a_����l���䁒����4��֏j+̓�V����4Y�,ۋk&�=żc^��j�&tYwU�;u���{�ٞGn��$Ԓ���9toV�EZ��I��#�_m5Q��m�}�WRR�%�N|єMn�`�8�Ӡ*#|�h=L����	�fb�3��Y�[�&�hۡZM�d�.�u�-��1^�$�xFV�e�6���Xg��P��x,C�x�l�9ׁkE#�޵�`�X��Gۍ��o�L�w><��9��F�q)f���Y��VC��"c`W���>GN��M��N3���f�D�F�wc;t��{�'G
�8��5�Q7�1�8����si��AM>���&�s#���YFS^ܲgmL��Ffgi=�{gY������65���VJCق��F�`9�#.雈a���%5�|s�����"k"rs�bk���i�^r�ۻ]��O4yI�p��e�U���Y�O��{Z�#o���=��d��y��U�B�5��������E+R{�5idN��KT��K��:(��"o]�����.u�fځ�B�O\n�-,��pnd7qޘ|�@r�p���ñ"����Pq)��4��V͊���C|�F���IS�i�&�A'v:&#t��X��^�[ӌ��Nף�D/�I��~�[&��6R�mX���p��8��iL��U��s��y��������ҽz�XM��6TpVN�-$뵃ҔbM��Z|������Tm�(�9���xn�\�d��� ������d��պ7̵����t��T�I��r��k�ޭ���t���i^�"�89�E��\��M �����o8o�j���k��1�%+�A>ȗJ��^����/#��|�Cl�ekyW��4�u��i��iI����3�����%^��uGhw���տ?MXK�D��yiuų�$�q�-fƳV�?���>��,P'��>��iAR���,�B ��-E��AW���h"
��~�Dy�?h�<B�1��1�<�N���qv�[P���6@�[ڂ����) T
��UX�T� 8s��8���{�>7�z�(�ʢ�
��E�/����^"q�(�QEP|n�B�;�We��L��%v�uB��i)?�{�T�"!
� ���l����1�o�6[�	IP'�\)p~��B��i�.Pr\L��ٮC�(9rm��-Q?z�z=<�8G��ύ��AZPTU�Bo���s�y7'���� ����\�x�QEXT"��R6p�����{
���p!�$�pe��{K����?�y����!���U�{�QE^C���KI�,A�"B0����B)���=�b`�r�;���PhI�x���П��j�\�x�FZ�@��Q����k���zp���O��Xׂ�Da�������b�c��������t�4K�%�h(�j ��H��J��b��Q��X*����y���8C�������^�)
�$C�	RE*	R��$�d����z!���ѣ�z�=��|��U�W����?i��S!��W���,���L���?��VO0��Q�{�**�����!�5�G���	���{�?����tw}TX�첖�b�S�Q��=����d��B	�C��B|ü,w�|\�x|?��x�b���6�����2�G���? ���F��X�? h�g��(#T���EX�y*�*���	C0}b��S%	�X����i�u���R���?2v�P_�@29C�Z$H�{ �V
=E��k*
 ���pR�~���`Y�E���[��B&KB��	���C�[���]7i�<��`矼x:t�|A~��@�y TU�E>ɾ�>ø�N�x���*�~'�_�V]��hS˽�.y_��=C�� �;���'���{��{�����K��Gpy/qz3�'�zΠP>���=�>�>a�nz%��A�x?���is���(TQW�}ώ<��$��)�������G�U�~���i����C���W`w����v� �;����v&x�ā��!�}��B,�.-��;������b�}���)���SZpX>G���q����]��<'u���
�*�󇘞�1�K�;ǉ�w(.���CD�!D'��y��{��A��P؁b��#��F��e��?� 3�����

��@��~ X��'[�S�C�����پ��� ���i�����wS���1�p�t�so������I~4��'��v�½��/��ܑN$9
߾ 