BZh91AY&SY3=���߀@q����� ����bB��      <u�$�֔A��-�*lY*�QAJPPi�٢��am����
֔Zh�JE"Ql�ZhF�6��m*#L�*�QU�I+[k�t�+cXҢ5Zk$�KiSK[A�� ��ѡZ��km�kIA�EFm�Ц�j�l͋V�[T6F���Ţ���m���A�� �n��l��S[�,v�-�k6-�1�m���!���[-�͛F�kZ�UkKe��֭������lŦȱI��Bժm*5���TԵSmZ��kKV󛐴P�ұ    7]_Sf�-�����9�7Z���iڳ:cUsiGJ�۫J::յ�ns\&�	Hs��K��bӪ����]���ֶ��̭l�ڦ�,ٵd*k*��   ���  Û��
P�Z�+l:,��  �:S�V�S:2��*�Ν]@�mͽ�z��B�=^�A@W=��@�u�A�L�l����mU�x  ��z���� �h�s����`
��@���k�p((PN���z ^m�hB��s{������htz .��  	��vV�e�6)A-Y�< �x@ �ŀ�En�{� ��]ނ�oa��X R�7+�8�� ��� =�� �l;r�P �m�ꂔ(9���Тf�[,��6څ��x O��pow��� wv�ձ� Yˀt($�9�P sv�h4q�9
��@Et��SN��-\�uT�k�6lٶm��#h�[-�� ����I��  i��P��� 6����@:`����K� �A]sK�t f�uT yV����6��F�X����ٌ̦x cxC��G@+�� �K]�:��˷P ��C0��f;� �p j��\Z���Y6U@Se6��x  �
 {8  �, �(QA:� r��뭸t V�k�
æt
���� v���6�٬��)�*�Qk�  �� Z�(W�N�8 0 P읮 *�0@Z�
��Ҹ Ѩi0 (���5@��a���Q�S�H���   �t��i� ��  .:࣭
s�\� �t1� cu�h gg  .� wg >�     @ ��2���h �� ��i�R��1b `@�&��~&BR�       ��@��J=@�`  `D	��6�4�LFQ�1�����BRA�QJ�F�    �=�|{v�&��V�m�����~ala��+e���~Rj@��.���:�Q�3���_*�� aL� ^7��PAU�6�A�:����������
���b""#V¨���oq!�!RaAP��M��6�,	,!��fS0���&`3�fS2��̦e3)�ØfS2���`s������G2���e3	�L�	2��&a3	��f0�a3	�L�f2��&a3ɘL�f0��̦a3!�L�e��f0���e3	���fS0���&e3)�L���0���&a3!�L�f0��2L&`s	�L�fS2���bd3�Ù&S2���a3���̆d3�	�	�L�f0�̦d3!�L�3��f2�̆a3�L�f&2�̆`3!��f0��&d3��fC2��&e3fʃ�s"e3*$�#�s"`̢9�G0��A�#��Ps*�dQ̊9�G2 �ȋ�s � e̈9�2 �\ȃ�s"e̂�@f\�#�Ps(�`̪9�G2��E�$¡�As
aQ�"9�G2 �P��Ps*�	�G2 ����s�d� ��3�� fC2��@̠��2��U�ȣ�s"�`Üe3"�Qs(L�9�2 �G0�E� fD\ȣ�a̈��W2"�A0
�\���P3 �*�eT3"�s*�fV`̪��s#�\���&g2̦a3!�L�fC0���&`�3!�L�f2��a3!��!��f2��&`3)��f��f0��̎e3	�L�3��fC2���&a3	�L˙��f0���.e3	�L�0�0���&e3	��f�2���&a3��f2��V�SO�^��1�U�����V���m�TN�[�k0:�rӤ�i���c2�lj�kn} ���s*��X���j0�%�V�v�j͵�뷟¤��Z!��Ck	`TX�ٛK4k�-Hȧ�e���x�F������i���M��"%� ���ʎ�fۣj;�9�5=L��Ƽ	nQRj��N\r`ܺye�(�>��F*��c �q��h%n抳��Zc �a��/D"��њr<R�w�2m��33`�M2����M��-4��
�:�Y#P�J�7!��
��Ÿf��h8��F�f`��Y��%��r���<//�f^�֕��7���F�YHMڔ6�&�]�ܛInM�Ŭ���q(�;����s�)�[[f�E��.�����ֵ�o��Tod�bb�̆�&���*U��)Vb\74��[��SCEh6���뱴�:a�Km)#��- ���>-
�l(0b�"�v�S�jR"�n2̼ݺz������a�;*�I��2�ɸ7k7N�)Ӵ�Ь��U����m-�������$L��R�أd���0J����HeG��4H�b9o膵ELPr
��A�ȼb:�V��T3Ec���K�֦�w�����j։J+]��\Ʃ`cNT���t�{�4�ơ���j�nl�I�1��[-�B����3�":b�������_M���N�+u���&0�486Q��h��(c�[Z�owx0*wn�U�T�2\��`q��ֱNͦf�{2��Y�v��.�S��0�re�'��b[tI��˽f$�;�>J�`	���'�J�[��񱆛�V��c�U9H�3���.�K���}�.�*��MG���T)U�씯P3j[ĵ��Z����	�,4Ӗ(KR�����xU��
�Ɛy,]Ǫ�pfS�DYc7kt_��n:oU
���x�U/q6v0�6k$(qL���X����tM�����~�,!���F�=�Su���W���1Ób�������M�.���z�k�R�S�R��� �#�Q�x���+(ho���Y�������KLGC�5�����m=�B��D�rbЕ��e�dL�*bY#*[�v��tql�E=;g!6)2�Q�R�uX�zw�ɶ����h�rAR�VZܤ�R;As���D�0�ov�d���v�	#S����R��d�5�^�I#��ĪU��m@5�VjIf��cR�eI[E�Z̈&�T��8��VLHA���Op-2�U�w��hff'��Eޚ� AŪř���J�/0�k&��l6��l2��j�F��F�m�kM�0������E�6���L��&hU���,�jQ�vʎ�w�e��6Yb����b��RĚ6-�y�+Y�b��z��5A�(ٱ�qT���1��xLs%f��a,���\,�]��w�� v���N�Z!�����mi�B��96��w[��%C�q���@�R�w �����c��h�&��Հ\�K�Յ]h�):�ՅrM��zr�n�^���l2��Õ�T��U���AKRn�2��(d:w�uP��Rդ-M,a<��v�[=F�=\ؼ�YN�v�$'yt�w�;f�c}�t|�Xg���[q��5��x"�+&m\��q�X�=����3oS��7JN����p�4��n��J�z�<ʙ���*0�n'����6���V�I�	�]���zB̃]�%��e�ܭW��c^�ɑ�ڽ(��,�%鳡�4��
<eHۼ���w��k1@��̰ 2 u��
o^nЫ.]���d��4 VT��u�G�2��J]ʵV���
Jk4�T[u\�%��E-�Y�%=�x��열@̤��#XjB��4n�@�B�bAuZ,����ʘ�%dBi���?�Ų���)-#� ���4�L��D��,�c-n��n�2�[J�gC�/K*cV&��V�Y��u�4�`*8(U
%�#s6������R�͂fRd��
��0�ʕ���t�H�\:t��lG,�9���i<�F�4��5�+YZS-C�n��n��Gu0a8���n�䕗�n^���'t�]/:�laۭ�
�ٛ��GeX�Gmg�^�+ELu"����j�[����(2�DnҖ6�8�a�.bd,�.`���#n�mbv����ݭlۣn�&�;�ѸL6��Q�mV
Р,I�X@��mc�kp�2���z�i�a�2�7�A:/^���-��I����n��f�n�Vj^Tr4a�M�"��u��c"�9z��b���XE�A�&�1X�h@��t�7���M��*`7���ڙ�V�bk��B��Ja̰��{fY��ۻ�z+i2�<���)�XW�����rc��Z��o3wf]�4ޭ(hڽ��t�0WQA�wS��t�Yp�5Ȳ�Sـ��Yr��f�<�cݻ��d�
�C)�KL*�&)y�T��R��P�M�2:r�x��f'�L�$�ٚ��8�Z+"����J�]�+,c�;����`���r�*�F���+�e���}�]mw���i�J�g��ū:�b5�[����9o֕5�����T���9�v�]�M�G!0%��n�n
FԱ_E4=1��nX����q��:����N�BÏ���)S(�t��җ����wM��+���R��Y�+_%R����L�Q��#v���p�*�ش&D��D�SSVN;��{yA�ZB�-skH.*��<�?!Xrf�	't˘��ɂ�vUdR���pAɕV�+)��Q���E�m�OtX�e��-��t,�,��䥚�L9laH;��BR�.r�l���^��(\�9�XW�%mO�E�0Mo�-4���1�[ct�\jҭ���/�j���?#<��A�2GHB�Vc+��[48���.��r�B�Ї�C{v���x�7I$j�XjY�&�B��3M��k�!�Y*��;-*X񺼨30=��&b�܁�r1Kn���>[����m�pmT�Ӂ<�c&A0b��6����F0�[`n���wQ���,L�ߣ�q�wbmc�n:Ŵȷ��o�L7gd�P��ǅ}coRe`d{�Q���%��p`��X�BS#e\�EK��v��=W���	��t���46�GF�nݻj�u����M�:+,A{gej6z����Ż�WAa�wkC�6j"�E����9�6V��A���=L�Ă�����8EdӗPm���`�㥙�d�L�5,Åmkb��  ���շQ�:�X�y���aG������'���9eMŢ	��׻W�����%����
j����3rA��B�7u6��|c�.��Su�6�kM�����B���ϛ�{]�;{��B&
7�����\�GZ��1,3�A�$�b�֣vB#�\����-�#,�5�Z�-W�z*e���)��.b��{�Q�˺àE��c� /�T7V;z&P�OS��o�)�é7�
fM��9�:l����y���=ܒ`4���Y�i�c�c�b�;�+v^E�jnK�ת�F��I�*-аУ�����gQg&GR�h%>��%�1��Z[V��dI�$Ұ|j������M֐�jZS�ː&t\Ǔr��6�搭��ƙ�'3p��P$-��V���bz�KdF�`��O^���Ր[Xv��A��{��u�O+��Zrʱ�����M����ȫH�7JڍKGkG���/U�V�z��7^�vBY6jO �ee�� &7�C�u�
J�[j�8SZ�J�-��v��i�ux�AHݰ3�A��o�y���I�9�H�Z�����U��*�LQź)�\��A��b3��ÁMy��������	K������Bc�N����+օ����mj����!�6Ԓ�:q���Ңuy�G7%�:��{�k��Z�meɂ^	0\�Y��6�­��[E���5��ky1�:u�f�r��tEĶU�*����"�x.���H��,�J:8��k�7Z��o�*fc�9�@�T��he����t�Gj�Ʋ	"�e��m��+8��=q\4	��慶�ˆ��r���`hj��I�x��곥��֚�f4i (��;'r14]hM^%�BIܭ�v��и�b[o,o��Q̹�H�&���V%�L1u��EA�u����"�h1}Kr��5�6�&%��5d9k^H-&�N�n"읗!a\�kDwG%�R��F�\�L�X���{�Yy �wV7d�����:ӷ)ޔ� � ��)��:j@k!�˽4��'q�9�ei��(AGTy1[-�=XM(�i�c�:�h�̛n�MYa����Y�mY�G	ܐc�1m����V��Vc�#"����!K5��_��Gn�Ӂ##�#�������:Ã
}�M�;�$n��s�J��VS��0VS�"�lfPq�� A^D`���4��V��V�iRU�	#0�A�bb���b9JƓ�U{lJ�9�
�/&���\�Xl���5�i�S�!�J]6Xׇ	ctZ�rm[ofQ�ӳZkFBA�tD�� 4-+��C>x����WYq dT�SB�F�H&6R���5��ol�Bei�V�� ��z�]�[�-�T0�&RU�P�b�n
�l:D;�q��I�����K&b�Il=yO��X�R�mѕ>ӻ�ݼr��l�n^MǸ$ӻ�5z7�՗>����(��ȑ���ʸ�u!��p�w�
Ɉ���܀�r�́��[1�Ѭ2�ʻѭ���� ʳ��Oe�A�7(��-�v�ݭ7v�e��*�L�H[����L9y^���X{&a�*�r���[Ov\ݚ4cD�<������E�Jα���75�3d��l���	4^�JgVьoe�1Y���k gkPAeW{`�׸��S ��Z]P`ע���[��Y#�����śQ`�h�F��9�Vf��)Sc�*	$q^�4:U@��sd�ba�L�XWN=�6�e F���n]�7�d�Դo&�q��VIy-#��V��J8a�I�;Hb�k�c4:a�6�V�Nզ��V^����LS&=�2����0�ܕ��C�ADZ,;Y�f홬��O30�fs���B�&��E���)�Lw�Vmbʺ`Z�lkx�q'.�B�ʷX�ـ�^�ؐ�+u�D�SZ����bO�rd[��rR�R��q^��X!���Z�.�{[m��\���HJa��������p����L�2̖+S�,d�,&�.���̬�oiV���4�-R�I[���)���#/��:�X�턗$l]s��ad�J����Y@�2 -�ۛbv����j:���S��,�e����`y���@�,m�ʁfǛ-D�KKf��XQ�vd_	*�[�VIJ�"�)-���F�˗Q6���r�n��#��^XG82�u;�-�����[-�0U$���U�v-Q���y��|]qx]����TS�
٢�иE]=���upc���bII�N�)�����EA[Fʫ�e�A��tsnk�-l{s,c?a^	���W9�c�2��ٶ����9Z���7/A�M"(3�[��F��w�7��0� �Wm��(�9���DV�,ҍ�/��>`Z��C����/&�y�T��0�Z�^��`�Ǩ���\Z�hHW��s%^ܵj��``㢘�Z�lJĄ��4T8 /�Nfʰ�,G�;�i��3v�wh*�1��Qc8�["ǴM֪D�ݫ�1���4��x��̽Wdk[q�IT6�B$eP�k�%}+Q&�HmVe4�S��@��6��a�ܐ(��L�����a��f�Y3F�q����v�d��
h��QTɐ1Z���fS��X�+b��A��@�d`؋{Wv5X�n6��œ)��h A�A����7H�Z9����]�2oR���vDAv�-tt�u��f=�[7,ce�:ډm�1�קd�Ve:#r,�[Am4�;�x�ńڤ-�B�l&h�;>�*��@h��y�U��rd�*̚/U�ٍ'l-n�P�j��aT�3@i9��MF�6��kT�c(���L�f<n�bNQ81�.]dV�7p��մ_զ,h��K��W>��V�ЌY�<;;(]��S	�lM�1�Л��-��T�Qie�{׳o���0fH��3Mgm���Z(�@�/r��;V����b�"�х���c����0�q��sV���+F5xm��h��<z^I��6��:&\�;���b��+t-7�T�F�2��`��s� �`�[Y��$A[.C�i�@ݧ�DĹ��r�Z��
k!ܡPb^X���l�����]�L��t'Rnk�A���ާ��0����r��[i��A�e�J�`f��*�<�pU
�#�l�
��Wg�<�^e˺!��f��q��S�I�����BD�[�7�a��-6+a<��Wh8<,�N���E��j��-f#�4Mx�-m�lWK!f��z
W�7��Z�`(�Jr��\�x�v�qBbu��D-u�G'�W�\���e�4BK���^G���P<0�����/�}N���2��b�<�l�5&��w��ZHI��"7),��� �y�ⵁ�e�=���5���`U*�9���T�)������y�胻'C�r$�җ�k�i�QP,��YshܳGN��$SI;8H�^
�Ö[�0ٓ�S�ר�2g:X �*��"�Ǯ;�w�n�:u�6�-LؒG2��Jp�N+ ���.�!*���i�%��Ɔe�3@k����⫐��G�����m]�{��q�d;c�Id�����m��cb��%:S-�aH�F�(%4t�*��{k\.���J$ì�f3.=��V)�f��w�Yv-q����#�	W���N�Ѻs������M�8����K��h^�	�Ï���B����S����}�0OB��!:A���%H�c�,:r���.K���`f+�HQ}LTŋ8�x5\�88R��]{�!"��;��jQ�{�Y��p��^�[%�X��녕c7���g;lk�i娝�*�VԷ:�%���&���
}�6Ŋ
��ĒuZ\خ'÷�̋}=c����O���w�.�Ղ_(���:�Ku&�IL��۫B���Mc��1m��$ɋ�nJ1�ԓˊh�aw�[u��6LBLy�ϖ����*9�(�n!݇o"c��4�u���q΅f�Ư��lev��c�o��aw<�qv	f���5*3����[�}�6ơ�j����L���s���E�f�q����l�ZL/IJ�2º�+��vjԙg�ܦ;���9����ȶY�z1H.KK�Y�e��M�p�G��X�P��9]�L��sk�r tn[H��c�H�W���k;OeeV\��-]�Y�	}��M���+)��-�öL1բ�J�B҂�˾��a��r<Ь�KlWm�Yy��,P�"����p�pn;i��Y�,��5G�TCv�CE�� L����Oޏ�e�پ��k�-���,_0�h����=�}Q\ �R$���9>�V1�M��A&D�=o_p��BU��G�4=7GV`*9F�_Y�S�C��>�6�	��y�����t��h����]íc�9&�-�T��@�=+����7J���!E�Y��+����囹�:p
�yLh�:�f�C�v�w@>��{�i��t�$�#B��M�O
�s�����ӽ`��(������Go��U�1����w�Qۛ'6k�ok�r���&�.�i�J��/	�;�&�S�c�U�'ت�!��U���V$��!CgžsZ=9��y���x�4ީZ��C&%]��iD�]>�t���F���
'ӌ����^�����M���]u�͙J�<v˕���D#�p��xa�8�-���� <�Dn�Υ"��2WgQ�i��DP�՚��vcY�q��:od�Yـu�4�R���5ju%�<Gwu]��XbCB6	�%<�aݙ���
�T@� :�j<��괏mv-IӜ��D��M��o�(��ثQ���z��Z�TژYI�*�Q@�iG&r��{:\��2�Ɨp�8��\�[���rAf4K߭r�6`��s�4��gYE��%�ƗEǫ]cv��TF�)�5Y��2�az���9ZS��W[��3e�4�eJS��ڇrR��R{	�ڮ��[KW2���"�	2%��M����C���p�܊���z�.�+�d�p����a#4^,=��/A2��av9�ذ��KSDZvE%��G�0(�3.ي�;,�[��b�^n�Xj���b���(�vn�Y�Y`����⺵{����0Zr�u��G�`�z�<�s9�0s̻VT9���e�z4��[3mm-G)�D[��曘��N�[���{�X�w�u��0%H���[�DvB���7{�SJ��hX�g+3�Ʀ�]:�����[���ج��R�A�&'��,�o���*�Î<{���i�x���;�]�u��]���k�I\�����,"�va&���6�կ�b���7���ӰV%���ᔬ�یG"�Wg@�'G�!���r	�ݙl<Wo���ngk�.oj]ǃ�u���`��3cp�����HC1f���Z�n��+���h���KY|��o
kZ��f�n����XZ{��ԓinl¶��)��	Ƣ�6��D YC2�Z��µ��x7�uځ�nS�n��V"7Xz�G	y�e�GZ��ŹKHR�ÇV��o��EV��W1F�X��67,ܩv
���g9��(�Z)[�f���RnA:�+k�Xkjsb�_CN��P�u�o�r��o�N
8�:qws��EZn#,Up�v�j^��.��i�7�+j7Mm(��1n�ꅠޚ���M����W[�QW��{���/��d�%�5v�
�ZB�=V�������GJ����2v�on��%��G�YD��P����Y�W�C�������Q��BƮf-��3CP����7�}����cWf]��(��3D�*dLXm:{6��Ꮴ_�gjݧ��DE���^��U��f�e�$#K��"¹�.R�ܔ�9��t����ޅD���I�s�vrpp��;�ܰOP���&ہ"�M���"����\��+��@]g�aVi�N�+�1C!�Y�7b�<��DQ��d`ͮ�;X���<�ۙ�����j�`�3,�-�5w�UY3�e�T=Zt�ȹ�R�ig��(<�=B�^6���e����۽������p\���9\�)����̬���1��ک%傟Vk����Eɪ�X��|�	i;sH66M��/d6�K1)����w�SX)�/��O�L%ӗu�+��N�8�V��o:%�_IzghنZ��J�� �U7.��*J�����5�ldL���G�Q���w�]�d"媹����q黛Z��R�>�.jb#j����ӳ�[S��k�]ш;�����J>�j����*�p�+��٦�T�z�VZK#�6/��y����aX>�=�K�)��\]�NjG�ݧ�K�5h�:�^�-1x��E'��Id/׎�ۊ<g_�nh����x�o"���.���Sl.9p�9ގ.��&��u,]��y>��|6�XA�*�ù(w���=4��4%�|�$��;�q�v��u�K��F�uM g+��,8���ܚ�J�*�����y �ŏ��7`�s�fZ#�N
�X�O�;��K�bD&
T�X��jw;:����9���к�L�����N��y>%�>n���nc�LS`�7YOA��7��[|0y�um�H��ٳK]]�mM-^����:��.]�)Igtf��B��Y/Hv�n�3�`N��%=3{�jS��X�A��I�2��8�
cz�,�XL����ȝ+��e��q�e��N+V�[�Ȏ]�ö5_f���}(9�zW;x�b���@����[��B�1�w(�:NSҊ��I&�GF�f!�`_-�Ѓ���̿���t�=١�
�"������7}��{5Z���B����|�m^���{ݩ+�2 *|�$�2��q���9�t�gS�['Z���b��3 �C��ow)6����J�b�Ƭ�.��Ҁ�6�u��vgQ��6op╚A�+�Y��ܽ=w�����j��;[�yǴ��D��p��2C�E��Rv�:;f ��^s]S��)������;��G1+�v�f��/.�oC�ɜORǒ�#��V�]��C�6��Fu(ގ�+�۱-nl�S�A�#��m
�'l<���!7h����}��������n�-=�n�Z�=x��WI�Γ��MzF���A�Թ�@�KtUʷ�E	��0�u�4z�^�iY�YQ8�JӉ��"�`�a��1�ˮ��3�#wLFW5;�˧ȿ��6�pG��R��VOB�Cr�iCm�`M�:�qVۘI^����˖���k~x�b���+L���A�i���G����1J��D)8}	�v��J�M=�ªG�KF!��ݥ�Ƈ�3,e�B
՗���:�X����`A=;���`��c���*��:�]�&��2�@��� -tZ�sB�{�5]�Vn�3yt+������Jܹ0���x���k_b��:�ɢ�P�������ܷfD^i�4yusVehF�����u��Ş�'ӍI��f������0�*��x��e��c���4��2=��^]����Μ�t(��wm0z7|��y����QG��W����F�����_q9�l��N�Z!���sr�q����Q�Ѓ��b�e�D:�Kg7u%Dn�k�r��b��Yq����u2�N�(�4��8�t����݊]�˝1��o-
�G{�>t1� ��xQ�g��ȧη*�_oS�-�Y�=�vAm�4pbpMΝ%Y�;�۝�v�v%B�a;�t�ni�0��U�8�V�q�+^�Ԥ\垎�k��	���J������1RY��)��D�3�cWydEݪ×�9!�{��*�!�c~������f78�n�Xd�w����),�׻$eS<�U�{qY�����nG�
�ܧ�6>�hT�q�򸌰�)��c��p��T�0����)����\�����'��QQh<�c�~z%ߟF۸͸8�Gl��-4�\��h޻��n͏Z�s/kؐ�z7�9��[|ł�d���GU&)�G�	*�xЎ��AH��Y}��}�JfD�1l���CE�3da��l[M�G�3�z����*ӇiGB^ݼ}+�=�m��^\�-3Q�B�RP�m�ή���S�p�媍�q����z�N�%��{�+�jR�	�9�2ͥZ��̺{��k:oLe���&�c�OWV-ދ[��`���-���S��7�ξ"vP}�6^���f����VR��a�b$ˎv։g���u���=D������~��(�v��[{s��Qm>w�Z]H���|������Y���0l"��q�3�ק�IB�TT-�Ȝ���*DS�ܢ���d��Xf��N��N�$	����D��^�l����+�`�!�ǹmeARP����X�xS���Ԥ�j���6_KU�DS��[��y�msx2�T���L��n:�ڱ޵��m�}h��L`�tO9���������E�59��A����Y�co0�n��Kw3:����׶6UE��;v��jKqaھf�.>T�2���]�e�g8���[U��V�ME ��:sE2t�Hґf8gX=	s�H����qt�����d��R��kyDrƙ{�X��u�٤��\k��v-,θ���7So�z�ư�"n�23�z���W�8�Ɣ^�婙��'q�uj���B3IC��kTx���o~_iU�M��E�Y�FJγp�P(vЎ��e���v�,�B����.�f����^h�33��v�
B�A����=��;�ؕ^:kFͰ��).���3��z�
�o`ڊ��::�Nr�\GwB̜��]|��Y��hzݹ��$;y]��8E�B�����=X�A��!��}T�o:�3�<�*�{J
c��I��r�Q_e�q86'���J�eB��7.�QFU���^ʀ���͟erlݮw���n�c�^�Q؛�E����
��&�35]irʅ�z�!`�l�Y���Y�4�O)c����z�Ğn*кK�*1��S����F�a��=L�n� 1-�㾫5kjc�����=Hkڻ��atä8p��,AA��U\���t����2Lʃg0䮻��۝IǶ�y���&��q�m���U�}��P��o*Qu��r�n�d���x9�F�&�n�z��j6��4��0����ƶI\meBc6+���a��7���w�����_Z6����m�E0��Ҏ����]]��8��n
:���M�)���g�f����bVŅW~���~���u���L3f�D�6�t�Vq	ɬ�N�H�7m٠�[�tUn��b��F�\�\55�gK�.]��5�̓�����ux��Oޯm��s�=�fU:;���2�F�d��~�w�Y�f���ݷ,�	�f8R���t��`Z�,vdk4����j�N���+��ŝFf����5�}����$�ȩOC�7N���|/��w��M{&�"{f�Όռ$b[`�g�v���Y� @Xۥ��l�+�cz��i+1��:EdB��!��X���I �'lv,��w��&l�nBQBe��3�5w�zU�2n₄M�hen�-ӭ�X�4�d�L�'���ȫ��<�V7!�A�"��s6�<iQy.@�l�N��R�9���4���C�]�f���|�"D0�HX�bs��9՝t�7�J��3��)8q;5�l��j�Q��A�\�Yl3�b����|)�j%Yc����-ݮN�n�����3�5��Z�.]a�70+<y�u*�S���i��C���hWU�-B5�K;;��<�.=+)�+y��i��͉���T�Xf�F�[�}d�z}�wOiL��7��ɞ�T�4��#�`���r�
��B��<��yc\nސ9M�;�Jk��Q���FO|�Y(5IM��8W!�<�eZ�n��N�R^���u��wC)�N�N�p���m(lJ��Bq�S��jq�ʼ����ےNfqGP��y�:�Nz�L��z��֢ɤ rl�j\=]�s�1�6��z.��39_͋���x�A
���FS�n�{y�q�*9v��7��D���}Ҋ�mɎ���f�ÖA�IV>�lȜ���G'�<��=��I�!��rs��%%A�R��Sx��&Zm�����r�w���,�sr<i˟n�Ke�]�+95d�4Y�+��;���G�'$��WNb�x�a�-9)���.Ja�똭,�&�dB�0SwAc�)PB��~*�)5j�A
h�����U��)�A+�a�b����P��(���X�]���$���9~�$6�,W�ء��Y;�ݢ	����M�P0���	�2�ª�F�K��c�ꆃ
��`)eJ4̂ZN�B\��WЦ�mwB�j�(D��JpB(�(>9�$�0�٨�O��5�!Fi�(�ԤH&�h3�RD2�!�%6"�b�n�OF��������(#q�����	_*�:4�ȸ���
0���L�l4z�ٽ,�0頄��k;egD$O�0�0.�yV�E�Li�m�W)I��ב�TQ�5A��h'�C��" ��-�&��3�(�Mq�k����U%��ۨ�ׯ�s(>�8L!:�^e���c.�����%��}I9Y{�Ġ/p��c|�:�^��Z�:] ����5Æ�� d��, 7Z8�D�Z@i}��b����J�2wo �7'C`���[�wVN��tE�̍�V���x�V�*W��T_(��%�����_.r��W!|weE�-=�Jٯ�c��Q��U=�S��uMo��H'�1�W�B����d�/��#�	W�us���QC���R�k,��>%[�Y��bkj�}4�SPU�ugEX�XfWf�
C����6�m�;�I��=-d0��4�H�g�A���j����S�@�6u9P�
�]��%֫���Q�[�x��m,�I��$3M8�N��`C���[y�-�z�}���1ڶ+n�eu.JS�܎�j�w�����ꠘ�N�`�7���{��w|��pZOt�ĉ��"�a$�����i.���8-�f�Z˧4��q�w�q 3Ek2ٸ5n�Y!���'iPO=��Pͳjl*�0��.R�*� ��ʀ�8T: ��
Zɨ]vE��@�%�ڸNo��8Wc�h�V4�x�a@*5�k{��+lڝ���K�ݷ�\���X�b���u�����D�}��n��F��qpm0��n�>�-��wp7t�&��4����B����߯����?w���}>�u���ׯ^=z��ׯ��^�|z��׏^�z����׮z��ׯ^��g�׬��ׯ^�g�^�z��ׯ׬��ׯ^�z�~?��������ׯ��^�x��ׯ^�޽z�^�z������ׯ^�z�����z����ׯ^�=z��ǯ^�z����ׯ�z����׬��ׯ^�>�?�}>�O���-��L_bk���4�2B
gB8��ͥh;����\ʁ�yW�#w�-f�6��*L=�:4����V�� 	-C-�ǻ0����.��L���oJ��At=#�0+���a����4qe������qՓ4��J���0u.�BX�킓&ٔ&�r�LY�-�Ӏ�_v<�mV:;Q 6��{Mݿ�Ea=wP�N�EK�h�bI�'YV���B�x��5�´lyq%+7g�:�9�S;��n�ʿ��DO���j�5�{��
���ML�{mf�JLꙬ|gZ7�+���W��i�k���N�=[p,��n�Zj؂y�yf��Vn11�K5�;w�R����/�O|�`̵$�w�`��>{��m�L�R۶��{��\L;Vl5�u(�$T&c�q���M=������{V���Ɇ�����/Yp_[9(2.�'Xt�U���䳤ބ�NtoV��N�i�G-r��� u���սf;�C���Iyԑ�jyXJH��Vhw;Ip[A'yY��s�K�+�[V��hE7m��ɑ\L�f��I�E��,א��+��Ϋ�k��Z��vȒ���,�e�ȠW5���9v�4���˲���}-������O����~�O���^�z������ׯ^�z��ףׯ^�z�����=z��ׯ_o^�x��ׯ_�z����ׯ^=z��ׯ��^�x��ׯ_����~?�ǯ^�z=z��ׯ^�~�g�^�z����ׯ�z���ׯ^�}=z�^�z��ׯ^�ׯ^�z�����=z��ׯ^��sׯ^�z���}�w��������1,@n�U��r#����'�de���H����f�c;�]u�P�۹@���EI���۩mj��Vku�/j�g$��`yb�6k����N��-��2u���r�3�w�,n\�m�f�ܛ�K�Õp>��Y�[I9��"-���D���Y#3��v�m�uԺ�2�q7\���9^+���e� �Cm�dR�I@:�9�AY�e�;Z+j�s�6�9X�^3��s��We�_:�)�ѽ�9,�;��{$:P�\l��l �\:�r�9���-���*����Oi_>uhk������
E��3([��:^�HMu�2��� H�5�:�;6�E6�F��H�q�`�a�h ��mSfu�'p��Z�i;7F�����ƁkD9"额!�e�h�'E���G���|*�s�nά�k�;�r*h9�*�GQ����Y��Ô���!�\.���e�&6�ԞNJ�u��6��#��.۾F�ی�pJ��67Id�D���x���U��d�N�@�N}�����rU����9k����
s��j�c�}>GVQX���U�|>W�
A�m^���*�{�h�X�ʉ�}+
Ln��LY��\���
#�D��}���D�5Q8�Z����PS2���^[n�̋R�	�W�ʚ�J�9���i]��f�Pd4z��ݘL�x�W��afm/�bY�f[�Q�gz+�/'fΒ[��m�c�������G[�n���q��0��n�o�*T�ŗ�ojH�G�)����x����,9��f+v:�-(�&i�@X��,��ols���Mw��*�P����S���4���,$
���	��C�E��]���L�"��z��TǷ������f
}}��%1d^f�U��M2T}�5��T��_>n�8�b�ZI���ӳ��6�fK��˦vP˱q���0sHZ;�62c�2h��J$s��o�D+0��o��k1,��ކ,K��yq�kP��v'%E������
UېR�Bj�R8�ѱu<�����h�1�or
P�)ݡ�5'ܐ��>�DIU�iT"%���Ÿ�;/�C����c�ճ$:��.�v�`�ky[�p,���M��R_c�`�Z,�eV���w9�b�E�t�q*&�]Y]�wu�*%a�)���X���@�b�B[ �Gbw�ҵYBv�J��闱7�R���By�.�c�#|�/bz��4	R��z�\{��a7���qZ�YV]����q�"fk�g"Ռ��i%�����0:�t��_s�H�B��N�b�\��ww�=�#Q��cuJ�\�
����䬺� ��t�
5ա`ԙ�'Rp�{���>K����8�l U��p�m��ЎH�	��P�y�[����l����%�,��T�y�sj���woQ�gK�]����7��;����4��O ª=��2�d�r�%3&��7T8����]�J��1T1T�%oA�#y�Sm
��8�&�i�yE�Ӌe[X��ŗ�z�^�s�������f9��5<���frv:�E����_4%^.�oU����Υ �o[�bHRy�9;0|�=�w�a��'f�u0͜�� !�"�P��NP}�f�w�H��*�I��B�o+oD(��J}�-�h�vQ��Z�kV�X�xմo��D�/&º�n�'��3_)[��ͦ��f��ڲ��B�D�#*n��yѸ�}���(gm�,��([�[4�PP�yTh�{�s�*o[;��`u{�Sl�η����r�j�'ga+Q����C�!��m#�/�:dCB��4'�4�k�g�{�g%���@�avEc��R`Y�ٽ`	\�h���OI����q��ʙ�/w����yn����U�/d=݀���%��5J.���'tc:PF"��;�T)U"-[�v>�l���N�v���o�P��a��+�9�6�^:�t�q�H�W����)F�-]� �ǲ����w]NʑM�XS�]z���6�L�zt��j����9���x,!1��c�P�fը�"�[ך�.�-:׮�l�(`�xamǵ��J�]n�:1�t����Mk�g��#1dO��EG��l{.$ZP^Nؔ�9WX�2�T�O�̛b:��RZD84R��Ֆo�GOvC#��a�y�z�A�����h�Uo�)Q3����+���e��kP&���rغY0�G5X�-��iC��ɝU��7ݔɈ1[�⓼z�W!����¥�C em=�",�����`o��M�Е.����T�0�\���-5l�}� Q���^�<+sQ�KU�˜]��Jk�9�7ր��M��6l�B��b�eI��M�Q��C�ZI�����kWXV9M��z!�Bv�3-��N��Nͭ�h�s�e:�Dx��vg!�"x�M�.�R�j3m�&��Ҥ�����0"J&�F��Ul�9���]�UgR�:�X�חݟ,{��ҕ��6�[�{���.�F�����pf	;��$����Ρa� �QQ1Y
[S3^���_q�R��������Ҳ��Y�4-PfF�79�	I��_Y7/*
��];0J��Q'.=�̲�f�<�e�o����WNsc� GD�N����Qd���M�f}}RL������E
f�s#�BA���Z#��I2R��+/#�֩q"��[��+�]�y}CjsB��d��������G1�b9ܮ,����w/y�D
����zl��F�V�y�J��	�Ы��,L����vݑ6mYu�0��c�H��.�E`���E�K+V�͒������;w� ,7;��B���n�[:�ޫ�^5g�,-!��HE�7�S�ѽy[.W:���W6�h��K����}��@��ו9�574�P&9���Q��<w���ϯ@�('FW��d�m����鍭��c&�[aw����RsF��jL=�G�[�}��Caq��j��p�(�V��e�Fo�i��؟'fк_N(]�X+k/��.1@]�$����t�ټUN�s5!zh�[ӵ��.X�;$D1h$5ї!����[��m9�mbu�^�is N=N�.��}m&�������s��Ϻ���r�- �A��G�7A:�*PϮ�-C�J���l,ۈ�-�{]
�\��|i�rV��J�Wqh��s�މ�*�q���`��&��V�!�5�vu�B[륐�[f�}��W{b�ٖ��f�Q|�*�n>�Y�Hǧ��P�%41m��Tv��iޛ���b��tP�q>u�;�v�5��d8����~Pm���ȝI����Pu�x]�N.wV2Ya��]: rF)unJ����s�����QL�F��u�Q�qe�{e��Gt��;�J�vw78^ttӂ�%"��Y�6��m6uTB'����]sGٸ˵�)ϭSr��hVm���`ʾμ1+�V&EÅr�p�K�z&���M���w��=OEb��@Fځ��٧ C��/��q�Χ�����ۡ�E�N:��(�����_mcP��
���/��WY���e�{XSe�ƺ��f}�)J4[m^k��Z�x�\
�5�
ňP��p<O]_vU�6Aū,� ���Ŧs�w���Ц$Ŝv���MԟF���Uz��1*��F��:�e9�~����*��X�;�ٵH��}%�\�mn�Gbr�b��^�+ o��6�ToND�����ڧwM���4�Gi�E��d�����O��9O�n�ؕ Ԏ���5-]if=��];�
�����ٗ�
��8H���T,��6��\�̬L9��].Ŝ�\l��͛g������ɥ�SP���>v��Gӎ�?�d{7:�ئ����5���y\�>�}���q;�[��w��ة.0k�����U������	.�W	��-'S}��I3v��{�wZ�-�=iգ`Cs�NІ��]}#������W�¤�ʕ���-gK�q�?�X�6�b���h���T��P�Spl�{���݋5�^Ȑ1��0�*����������Ż��uf�3/sr�6��<�CUdX��H�/-�ˬ��Z.q���%�"��Sy��P�㈚p[tj�)�l�;0����8����LŪ�΢�;OxE@�#7��|����o�,ov�ǒt"������Vϭm���v�M��핌+���/0����vm�oȃh���;M�L���e�ƺ��T��^'qd�I^ʼƣ�*�ѝƞ-c�F=�ҟ4�Z+k-�63^��J��e�#7���z���"��{u�~P�&�w7�%#��du��i�V&�48�W�`Y� V+�e*�)�+���1�`�3�8-<�~�&�g<m������_4�kD�e��z���N��>X�����9�^n�a�)����U�ʳM��Z���p���1X�jn�:��q��qLo"4Xf�Gi�����Q�H��],��CTv3���vv��+�yۑrR��y��<.�m��AP:����S���[Za�5��i���Djn�W)u�y�j��L�%fu2~���*Z.�M�w[�0�bKS��+��g]F4uL|2ʐnGU��yf<���ʛ�7��\����kiK/�ʘ��D�F*�V�m*��l0�栆]�L��Wel�G�<9-`��m��;~.��l�(�9�a� ��ڰP�,y܅n���g��yA���dZ�a�ח#���6>d���i�v�3A���R$u�u��o��T���������|��Q޲�m٘��:+kU/B��.v��&���-pF��]گb/]�d��u�;Z�^|�̡�n�Ne��{uz6��j'B���e�&ƶ��eB�,�PjT]t�sR���Ȭu�g
bU%�v�h�8n"S	gb'�Ls�aK�n�&�Hn�řĆ���d���a�YJ�V[�SSm�Y��WA���v�Q�":��;w��I]w$��T�f��::]H>'B�2�X�}�q��w��9�E�e �86�ȷGe�4��H�E��j��r�ނq3!�wv���;���M}��W�m;U4�ֻ�� �csk��M\ĩ|8�EgM��ą =�Wf��OF�׆E�[�ت��G��B��٬�i��Xʇ���r��*X��Z!�n�ݹ�I�R[R�5��r���ڭ�� �kG_W	(8e�J$���c�ޕ��ܲ�Q���7�9�tXvl�\S1m]b�[�K�����l5)��'6x;Ɏ���=��.pc�{��o�ďP���ew=�dX%=��a�t�owt�S��!�mX�u�5RY�Ɖ�\�ӛ�P�qtd5��e�0��ﯲ�jR�m����
��׈�؀���b�f�����^�����l��D��hT�3�&��J��4P��(�k1c���	A ӯ��,��ʡ�]o�;Ջ���N�)���X�F;Mv]���}�&��؇etY4.��H�Ꙉ��О^��#���ώksL%F�A�:v��P��*M���4�
��ۋ�Md>36�)��"{Dc����i��r�v ���3b2����*�k���yq�{�Ef�
k�9���_a�m���Eڒ���n�'e
�S����J/ ���b�Q�*JC�SfFLy�e�[4�����U��T��=v����Mu,�amٴ`�S�ڒ��X�⺰8�֍4:q��d}�(s�Y��3Ca]c��oºD�fA�;�BV)�"G7o�p��Vt4�8qg�p؂��փY�k�Ǜ�$-g t�H�vۦV�YB���*D��󝵑:���Z �Ŵ� �Mp�a��>1�W`8�ז��(��6�5tT��[krG�d�Mw�e���f��e�g22����rK}���͒�Hf�)���:�y"������BL��X��]8����9��
�r���j�Ej���p��/FΨ�vsFa8T˓w+��#d$�c:|��V&�!#Pk)��]�]=Q�t*6������V

��*+U�X��VY����ב��+J"N���,���Ê�"Gk�JX{�NG1����y���W�2AjKP"�H3�M"hC C1�[�$i��,��M��h�dQ�B`����T�2(ĠqB�7t�G�ZI5�z�pōƩ�m�i�TG9�Ǘ*uTcQSQTC��ܒ�Ts�&�ys\������z�~?������z=�	@PSS���6�;q�(���h�˭�"�c�(�h���������~?���ף��IICTvi*���)k��9<�4��CAHRUD��1$��ji���iH�����Vت����l!)���
����"j��Ӣ�i��"��)�f)�`��5MT�$�$�TD$TD����i(��`�UQ@[:��hh*��m��
hh"
�&���5��A�bh4�*��F!����y8�
�:B�)
(�a���� ������I�7�����������y5F��(k�a�̛�!�ʊ=6�<ْb�^���Ŷv�c#%5�!"��4bX�79�r�Jy��95��N6��U��eb�Z9`��H��G*���M1l���Z�jG�r8���˓F ����x0TrW�k���2sb�nar�h���-�l�n�6��F��`���|܎I�
�������~9�ˇF��矺>6/id��)>x-�YG�(.�Y)�r�ҁC�
ǽ}�4j��8�Y�n��l�f��&�|�(�: ���0���>��ރ;����$Ik��Ũ��M��+L��e������:���=�ì�J�w_o[�gڳ��h�m��fk*�o.%���$��Rك��(u{�x~�x:���^���x� �:��F[tY�ۧ(��\Ց[o�>��W��.a��ȭ V�{�	�\�O<x�ƴ����;{��yz{jٛ�Y"jB��vP�������p|=H
�F0U���{��Ў�^���s���k��gl�F/�^�Z=�|���^��v[�V�l{&��{Z@�l�Hh�q�y���b���ں�G�/b�c�"{�W����f{��:N�s�{��<[��8ȟe�~�14�=�k������o�����'���>"Nq����zN�[�㔝iy��ժP�I~P�%(��V�C�;�C<�W[=�-��}����}F��c'k��@�	�s��6vۛ��7,V�+Z�ʛ��w.���n���?@�"7�O^�ς5��}�"�]�3��2܂}�'V�v��}��Zr�hX&m�Ī��ݝB��7�M�Es�c���F��J���������53��[Jm[t�ԱJ�0b�r���׽�z4�׽W�T�l?y�ǻż�T�����Q��q�_z���=�h��Ϯ�{�q<1�)�g;���=�J�.S�l�XZ���]�#ŋ���=S����� ���|bh��d���ޭ���N?]jeV!���{q��^�������|Ex=����L���(l�6��A�n̂{�]<Dd6G<�`����9��0�E?�i���6NC�o�O�����ǕfC�W�����tĚ�3ޭ[8@���g� ��ﳷeJ]*������p����gdk�jM]�Se�.	��]��odS���{g���~�62�g�Wn{��t�����);u_c��y�ڜ�6L��ax=Xg��4�Z*\�:�9�#�`��ׇy͆{MT|c��{Ϊ��}<�����\f����{�\`��%��8�+��v�.r�t'���hc�Z�}�y�i_���k�ʻ=�.���@,]�uM��5�k���fZ{�\���pv'�S�vk�f^vu�r�A��J����t�h�S�z0�	�����`�n�4��/GBFͅp���y�Ӎ&Jsz�~����S�zz���y��|��o�p=�Ь��n�ag�j�Z6zǙަW�"}�>#��O��l��$Sz��ɼ�wf'v؝��|�95c[�Oxi�<3
��5�Y#v!���mM׵A�%?y�,�z՚����/x�9gf�����Q���^�!����*q{Z��C�*���')�y�4��_���:�Fkʈ�Sڷ��N�W����8�[���כ^��O8�����~CW�w�.v�I�:ڊ��Ŋ�N�Æ�xP����7|��E>�;�@/1o�k�+\�n
c�����,"e�5c�/u4�N�6�W�T��a��9
<^jq���w��[�n���S�s&�{�G5�����-��ݦ�TMN�^Y�+��2Ê)����gb����*-���tޣ簡C���]«����Ó42��M��H�0���=ӌ�.��~b�2˻L�z��c��=#��]6�ΧN<��kf�5��}�UX@	�Mս�������y���N�뜼򳲃��qw�w�v��>b�Vf>��d���;�u��i*��}����*G+�y�>}�>�����H�F���l�N��n���o�A��o�&og�����$���L�r�{���{��*j�����Z-��*f}�� Vq���g=�z��M��t�H�kR5Y;��S�٨e�/he�Ѫu��>O}�u�Ocf׽$;kR�L�/�]��g�{�����2�z�u��b9������f�Gd��G�1wF��̋���p��j���	a�����A��n�%�|���؆���@Vjmg�.zv�	r'M��H��4���/ 0; ly��MK�p�moCcL����.���=s����M�74������K�I�]'�w��<��Z~��uZ˟�܅J�?.�{����y��f���乐+���1����W�>��^�{Q�-o������x���8[9�����&2���1FD,́m���]c��͚�b'�vot���T���������i��"Ъ`_�L>u�B:��BK��/EsƆG�0ʢ��orX�N�XʒB�U�wG�pV�쥕r�7i} WW�l��:���&�t�"ᔚ$Тn�$���cq�.���Bu^e��ӿQ��7���A^s�Y�h}7���6��2��$ե�:��^����`��y�=1���T�W��~�0ňz��mgq3�Fw��+�*��N��xDT+�g��C��9��3ի��;�o*�
�����n��}u�S��L��D��"��F�-�F�8��	��'�siȆ�w����_�7���s����{^ߏ�|}�i>#5Ko�+R�=f��^u�&D\}s��vc'_��I�3�f|���<*�u��{��8��Ch$���+1ϫY�mG����"���ӳ�A49��{�2���L�q���pژ�ڵ>쵳�b��x\�>b�pb��n�{ȍ���p�A}�#rdy��?*��o_���I����U9��.����]g�����n���͝Ǿ�<*_����Lsz�d�>�l���\y����7!kx���]>򫡩�|�������JS��ᄿ������t�JM�����R#��?���
u�U����)]���Q��+�K�������
(ڑvcRj��ڦ��ݣ}�w�T��Mg�����cb-�e�C 3��AR���̝ӫ�޴:bsq����ޝ�&��f�3=&�����X��|�[g���}[�(ǽxxy����w��@ܛ�I�Ӟ�k�����{�s.��	��^6W���]{+�.��L�u��
v���{���V�X�Y޷���y�n��o5�oPq���t�h�}&p�ᵂ!�=~�\O�7���!�k���!�`������1Vn���hN�
��|C���2|�W�{��d̊���<����ü h�+�z��S�ꭍ<���7�vt�y�/-���w�������4=���e�G=پ�O[��b[�4��"&��fG�/�N�t�F���=�],fp�B��ٳ0��]#�q���/ѻ{�����#��$�5i�-vkl�{*���QF_��g���_V�1�6|fɠ2bo�4�nvc��852���;sZ�P��9�|�NG��n(���od��I���c~̶&{w���r��d�[����wB���m�V��uw�^�X��� �侨�t�p�t�L6�r��J��ȮX(�l��`nv��eLaލ)D���/VH��o;h��=c�����@;�$=�"cǮ]ϳX�m��۲f�>ތ��&���,*����@��rop��Gq�o�u�tstp �l��ls��a��x�en �N[��*w�B}������{S��xU{����us}=���k�=��WZ �2�Z�⼮��b�X�)�
𼏆Ry��ו;�5����$߼�h�lO{xz���/zy9,��}��U�X%<�<��k��?t��3`��n��o����lکg�̅�W�kn����y�6E��{��c�{֞�Z����e5z��;�?ux�߉�X��NT=��)s�[�+��k����9�~K˳�TƢ5�=�y�/�;��zG������ض��꬯q^	|׽_��p�s�Fo���5��gOf=2�.�.�ֹ��f>y�,�4F]���M�.�_��C
�1�`+ �鈛yNų������G}�܆[L�s�}�"�:`�Hfq��fYӋ�H�Ç(_omwZA"��N�P�aB�p�U��*,��
ܭ*��p����_#2b�r�T/Օ�(d��{s���銜�Z��q�TTd�Ӈt�F2g����
�r��+�}�2{����U*rj���u�OQ��E���;�7�W(V����l�Ue�\o�T!��S���Iܻ��Q�x��$͜���ׂ}��e������C��c�_7wZ0�G%bW�w�����g�3��ޔ��h�`�N�P\���oX �r,d[�Me{Q��dLp���^��ڦ 9�	7���L��ؗ7V����N��Wѹ��4=��:WQU+(�:~��=2z{'�>x��v$FmYĽ�񅐽�����y����f�lG���G0�~탘�MbKԖ_{�����g�FVE�����>`_�o�;�_a�'�c�����X_��Uݷo.����AUc��s�9���|J<r=�,5Jy'o$��v��VGmZ���oC�y�4P��f�% �Y�Vg��{�k�3��.���˝�2����9�U�U���,Z�Q�;��gVŝ�T�yksry[�n���N
=}�\��,ڝ Ոj�W�d]DP�q.R��Y�on�z�V�e+��a�^W�<��l��xxO��;c���U�>�=$�݉��@Cl�^2=����x!��}xT(�ڼ���S���∓���P�77ڽ��n���&���˷a�ɒfU�cps�,=�8�gѷ Vm��^��{��!5^מf��V���t�ub����:�טx��a^���9[����;7����+�ޡ}�{3��޲��e ������W�<�Y[U>��4뽾�y�/Ҷ�9⧹��#��tG꜆�_�k�>�K*s����~�S�,Sv�<�\ݽ�ӻ��9�A$i��IѱO��e���NTd���zi��{o�a�ӛY��r*���|7Iql0�s�{~{b���,?Z���:���d�9�D����j�.}���d�q>���쯎h��k��K\6q��72z�p4F�w1��'!�+a��I�lϨznS�x��Ϸ�>�d��.w�g��gc��NZ�V5s����fák�#3��"K��z���[ǯ����%�:����F���t큜>J�z��7(����$NZ,x3uC7�35���0Q�8�r�+�cOv��Z�Q�l=$8�ѨJѸ`���ˠ��������&����MG� ђ\��	�,V��Lz��Pg��eQ����2��ȹ�=���➮]����8%*g��K]^{]S����@g�{{����=�f(a^������$�fz�]9���4\9;1�t��!�Q��w��zN�tf�>�A�&��Ow�T��[;g9�]����C�]Q�v<�5�<��Vx�3���¼���>���<�~"?�dv�nf4k��q����| �^Ȉ%�C!�N�3ȹ��[��>B��򽞐)އk�ٻ�`9�x?�_���Ўz��W}�'o�?#U�Hw�뫈[�{��k=�6j.�����z<�t_�Q��|D2��پ�|s>�=��q��{�����A�=G���y}�X��Y��=�T�lf����\�q��(��W�[*�̨������,z�}��M������<<��}S�ɚ'��wj���B�ݗ�8e�Y8�F�U\�MZ�LB�u�������sAͻ���obHiPxOw5��1�1!��,�͗�l���t�L���z��Q����Ge?����z�k�_3:;��d[��Jx�\���b���!�F��Ja�,��+�Vq��鵙٘�Iө\|��)2�9O��}��(̎u�Y�i�Ϊ;��y��N�=�/5���4���P��hڦ�c}y3��P�ړ�^ݜ�Ϣ�,E8��NVǬv��{��ʆ��-�6�\OX֜]���UwGK7��S���s!��f1(�΋;�22�6��N�nB�8�V��Yݴ�*���P�1Ψй�E욁P�!@d|x	���c8��T��N�� S���i-e�s���0���r얔�fTg �x3s��M��\ޅ|uΚuM�.�yM%����n��c��M�U�zz��3��Ub�E`X�<)���<0@n�&n�c�Gz�zb9Qu�y���*�ĺ參xnԴEjѬ����ݵ8��\�V����1�sUf�P�G����5�u�:N�0S6�.��kgX�;;���/5@�X���\ �� 1b�}9F�����f�Nu��K�SG�f'���.ʦ��w%�d�`�B�;"���c(
��T�rL�Y��U�f�R����d�P�6��8NcI����u����¬��1����RW�
㭖��:����=��e�u��k"&��-k��Q��6U�A�Zm�̄b'^u��m�Y?{�ub���^�r���ԥ<jP2�Ā�.����Yh�`|�֘*b�nS�<g\ߡ�pmܵ�y�؎�M-�o��L,=MdcNނ=7�E���^e��om�PR�n��q��Ճ�����(�5�K�UZLdE�{G{v���:�v�:���ld`Z���Yx�,@9תp������W�g�p�jr����e�xӛݶ-��y@�iדi�6Q��n�%f�
�Z�U,�؊Μ+^&��$��#��h�<�HJ:�eb6u��Z"Wh����e��&.���۵UK����λ� �Ӥ)-8ڛ���SIի�yV!Z��ٳ��fe6E�:uҺz��
����b�k�$�'�*hi}���C>�v�-�!��mֹ�7/���w�nZ=��/�[h�;�6�B��	���yp�j^�>Z2�W3IIqI'�z=�1���V/��](0Vj�ƚ�+���*�59�"��;�[�۠A2��)h;��v!㔻'"���Y.���o�d�QiA����	�/���͋d��dFq��gwq/<7�t;x��BF�ńMF�˾��m�ץ<V���\O��6��{7n�(%�t���Ic`��5mp&�p;��oMD�T�B���7X�g7��Im&W�ϊN8k�:�v����{�|��G�s�?���F-N�66"#:Ɉą-kCF���N���((��ᱝ��δ��rb<��)yh�S��K�9N9��}>ߏ_������~?���ٔ�"�?�Q��+8�4�בX��-�/X�\ˡ�I�~Ɠ��<�y�޸�ȭk˓���Z5�x��'�����?������~�_�����F����7$ѧ����l�o.1�i��UT�E���co7 ��w�~܊�lEUD;f�=Γ��<�o�9{6
MkI��Z�,��11�MP���qk�b���7$�"����C������gm:M���@R��X��4�����A&�l;i�H����6Ʒ.<J
��Z"
CA�]TIAE4R�45HP:�D�)CIHP;ӹ%R�sb���bt:
ii�(����%$K��R�-P4��)CI�ꚡ()(y. "
j���h4:�h"
"��������b�4%!E@QEQUUZAQM篷�e���ɶ��ۂf��H�>�����)�v	ұ�f�3!��Et�,å��EY�k�=�\l�}'{���}�VK���T��������?9�$L����Y0C׸�8��q}���z*��$�W�9w��r��Z�3a��ť��[���2���`��H�d���P�%�=�Rpe5���g�拋�ُyj�!�l׆T��#ZP�-1�S���s��cHԕ3kz��A�,�`�i��ۀ�;�|�ut�W���1��x�.��-�â�"�zz�V0J����o)�����-B�4�Ҧ#-��ng�C!�~q 0jm����!�e{�3��^<c�c�{B���%�τG�!�.�eX-�%��mGM�i��]7r����@(�5�ONQ�b�Mn�Om�L��Sۼ	<2@Q%ٳv�7	࡭^��J�ES[��#�3��s�I��"S��SH�kg���6�ȸu]Ń����wh.����`�4���;�e�,�t>�U���.�L���)9o,�<
T�a�y���AZB��(T��rG���h�G�B=�G6�����S�.�7K��S��ѯ �{�\����\;T�1��WSǁB��	�~��-��h0Q�Ñn&=.��N��vr�j.�����}N紏hlچ�;�oX�� �^�v�
�����㽛wZ�p\�Z2�%K�%��LVQ��W	��	<����n�U��)R,Ye�,�{^Q��؁���h'�Os��bRr�DX�@m&�>����ҎDv��������/+����G�U��=����as�/��A�/�ߦ���/�ܭ��w�A4~?C�Q���h��hɇԵ4�E~���q����ܴ��>�+������a�f"�4p}�v� ��)�f5�����
����!�`�m���L;�ƲǾ]>զ��A~��#ƃ��`�89`Y�{=���I"|s_���t�jϼ�Du�oM����bXnqp�ߍ�sQ~�-E�;��50�B2���^���)�����u")��s��������w�;�#�ѧ:D��4]�ð�q�w��!w��߶���
�*.������������'Y1lS�`���43d�l�;z����:�m��\ܔ=�ލo{�/mt�H�ߗI�6
?"�������[�ߋ��z���7k[�%���b�2fV�C��h8�|�M�1<�Z#6q�8�t������4F��|Ǧ���)�&;9����s��ATV5x�A?1�A9�ƒ��z;���ǃ3���t���F[l3Stbf\d=����18�=��5{&?;��yEw����@�U�J§�L?�5�ܢ?���o�{�:�E	�������d{)��*;��-���� ��[/�o`��ַ��*�Hٛw�R-��h/ �X��Wwb���5��Y�-;b��S�.�����`��yn�{�W	�\��}�&ڎ�l�@���ܥoN+*���ӎ��_ٖ�i&I�����3�uOX�/�b��򛜫�U���O��vnЛ���	�{�1������N(�Эޞ�Qس�Fބ=���WE�'��ށ#�D9AĈr4���^�;w�^�&@�LP_q����Ǎ�=����r�q�� ��@2,v1�x,6����c���|�`�4�3������з'N�_Jt9���*���2����>z` K
������=ʀ�~\~������wl�]b�<z�YA,*�J熠������,i�a>O^��2���Ӈ[�0|n%³�͍^��C,6�-܇����yNW�z��0m�hUt�O�h��3�>�(x�o����7���y��|�$檘�;��^�̜q�ǥk�J	{kU s	]bu�q�l�Ʀ�_nJx�yB�0{<����i���2ɽ��>`�����l2�{�Ӗnu74؜�콢��yߜ"_8��1�T5X+�}�"@1��'��L!�6ߡْuٲ����,�ʟ@(�Wj���#ǜ�B	C�k���+ֽ�Y^[�$���DЯ��F~XG:vn>��k��'��T�#�5ģ4ۍ�l�䀩�w�`\��N����,��˼`_Ͷ1�^��ms�3Q��6a�ӯ�������*PS(^\�#�h�f��-k�E[ُM�hϮ���;Fn3NQ�E�֬�̇9�]O��Z�VUh���k��. �=�����ӽA�p�샏4L�C���].�H8"�P�xc��`1�2�..cVU>�Έ͓����؍�SQi�_��r-]�G:W�&��E�7��WL\:��gy)�*�8���V��P�,����{��x������=oM~Ԥ&�k[2�YB����u��ޜo���N�m��*����Hz��������"cH�0�`�ֽ�Y3��Jm�S��,R%;�q�Lu2h!jy<�]�C�z�i흠
-�ҠI|�1���/��4�)��B)�ٽ�{J�걎�v���e���S�f�IT.�����P��ꉇ�p1�$8���?���	�_G���]1�f��sNu>��.�EL�~	�C��}���P���_8�=��p5��H0͒"	L:3��6#mdl�(����r��9B�s��EL,#R���s�2�������4��^�6�w8돆1��Gt�����(Bn���g��)�I�;.����� �+���PN%Ϣ�[7�j�r��@���\< ��9ni����`�����r��@u���O���լ6U<Ke]�cYyd�XK��,@~ ��Zv�v;�5<����eP9�+�2�LPT��7]�kR6w�[�Vkv��@�u7	�sf�؜@��3a<�����i�DWYq���ئͨ^�}3RO��WZ��`��P�l�N9g��g�����+�x�)=��`c|-���t>��6ã���?TĶ*�Z�[Aq>-�,q�\�zY���Id��x�����ط���}�tWK����w;!w0A��s����C��i�f�y��]�/e�Id�7-�'���0��2x4��z1�q��P�=^v
>�	���-���sV;�d=3k��J��hјv8�k79Zd;e�rp8�s�-���`:"ط7�=��������gH�r[x'��~���5���kx�
'$���ޠ� f���~�]�������^�����2�E{��W��K6�!�j+���8~~05g�&@�n���2���L�^���YA
�%�=4�טUlm̟�m�Wڎ��?T7
��R��b�A�ώK���O=^�4�IS6ߎ�o3k�<�	��k;jk���N�!��L5�� Y��K�_�*��s�D�`B����"�������J��W���<�`��W.b��b����ڒ�Z�X��߄��oO�P�9�������I��~c ���\ ����ТO+,E���9���r��%�{�)H��Mw����Ο$�7^5���W�fx�H���U��ᾅ�-!W����L˭�
�Y]��6�"�;"��k�@ͱ�}c���X�F�d�ͭZ�n\̸7;�E)=!J�����|������V�X��<�NSq"t>U�����/?����<�1rd=���Xm`���}'�w��?�Nu@�<��T*��r�?�(���~�|���m��r�7�63��m�1����f�S}%�H�I;���])-�Ùk\���R���sM��.�����lU�zq���E�����x9�j`�m�{<�_
�cn�e�(��n[z����j2Uv�Y�|���Uژ���(�=����B�e#Ёgi��ޚm�S�S�O���%x�c��ɔ=le���F6���篿,Hw��c��C�1�^�1~�����"�!3	S���+zH��b�z���IO�`-2m��O�Tφj����+��x;�z��}V?VSfa���3;��$^�_�\�����+��?��W ����=5�{z�d���1�uے���:����!�m�	vO��R#kݴ���a�Z���m/�ܵe�ajxEoR��٤�l�斆׬G3��\Lv9���K�mם��ߎ
óE� �Z�QR�2�e&[/�:�pC�ώ�V��z/6����yѢ�ba'M���pl{o/�I&~㿭�a(3�m��U�X�`�Ù�Zz0����\:gi6��~������z�b��e�A�F��v�E�J�N�,��D�+E=wPZ�����b�,8;ejC�Uehu�$2M;�I��9�~ܑSڬG�+�����.-r�{4WD�-�	��9Q���4Si�������þ�>@�����	��ڣ6�[m������m �Tà��hѳ_�P�e��
I��-�B�,���7�D�zy<�΅���;lpw���3Vޤ=�闰�hpq�!��~Ke���<\l��2�"��=;�.1�x'9�\a<���˨�1[��P����NHͼ��1�t���vO@Z�,[ԗN3ю���z�8.<���@
Ɗ6����X���q�0�.W��X�C�}���uϞ7 RukU
O�.XKh[s��v!��kL�^NR���_Z���p�\��8����ȁz��]����2O`�JrQ�Kz�s@⃲��4�k2HC�oM�ahGM���mь= ���A��9�ղ4�z��v�}J�.��1+���:���ks����ij���+^�$�78\
�ao'r�gb���#���2{6��Ū�٧	��Ev'�}���L;"�{^��oyK�1�~�Pm{er�� ���AjG��):
�އ���r���|��F~�����쇬�~�2'*,��<7,�E�,J;P�Bxw��|y��ӝ��zȾ���[���!��D
d����F������~⨰u�:y�������q��M�̠�o{�ǯq����� ˵L�g.�&kJ_�H�fX��Z&Z�s]aV˽��3����1Z{�Q�vpk{��ac�Hz0�_l��6� ��v��{��w[�*�^k���Ȕf#ӬS���gw]8�>�>~yp����ߟ7�Q��\�g9DBmҐx)[��鏙2k���j`kd��д������iA/mj��륃�\��6V&��=\�F��V��8aHG����"�s@L3,�{E��g%^��l��א�����ή�$�TP�s�] 8�ל�����~�"]��d���(����#���oY�~�4[�N�I�tOd���~p�N+Ҍ��{ͣ�{C���,�(>��<����y�T�j��l^;lL�#M��<���7�}�#������ ����`vP�-3��X'�ow��g潒�Ub��ü>�TC�u�ڬJw���c6%��D<��#��Y!k0E��Or�s�Z��Ue��h�)�/��:h>p��h?����h��-��m`}+����!s�;2�k(R���ƫ�M;%�+5[=y�}�����Ol>1P�^��r�ׂ=2��#�~��Kfa��t)��)	����R�ŝN��Y��d��ف:����w)�k��`!z�����F�!�_W�k����Zl��QwV.�[n�&���xE7?<F>�.�Xs�E!9����E�;Ǥ8�oB����&	��2�m���6����v��mA�[.(rJ��P�`�ۨ��&a�
�+���)A�Ӧ�޻�-�����ހP?|��qIOz̭��(/��PP���y	yƮ�7m���ta='`��๦�r��[�`�}��E5ڦ�������s�D��~�����z�|�z8 �H�7��R��1,��g�\��]��������2w����0s�H���({Y�_:�A���"U�N��%�f9^�eKMCq~�,�0lv�cZ���go_n�H�Ekk@�f,�>6�2U���v�*��]/B�i���AcAt�~i�E��xlO��'4�!�#�~s !��^:W�vS������'(_&o��Q�Z��IZ.�����3�v7_9Ʋ�~���-�|�ǡ��TĶ*�Z�\X��6t."k��ɫP��LV:�PK�=�Q��YP��b�901��C�s�v�M0��o��j"I6���[;:���WDs��n^eO�9O���;0�p���z7���!�����5Cc���i��t%�>���%�]��1�/C�@�>S�`T|@�BG���J�ǿt5�:];��ݘ�x6�({CCx��M*�{��t�{z��l�m�<�hO�p�/���a5�;�l�;3lLFv�����>��J.L3����g��EV�۰a���f����s~d!�]���а˼�����p�|䥰ĮL�ն��S-�)�g)�f�w9�
��U(\�z&��+T۫�\䁓O:w\=x����k0�͈fw2*��cL�}���ۭ�2v�q�B�Cp�F��-�z�xz���/;������AO������ D���$����f��E<5�yg��-�(M�����S��^�6���75�rT:��[z{����CǞ�J�8�Z�'h={6q=z��C�S�{�h��E��q��U@c���Nt����ս3�^C�[�<�Bu���T�MAb�U��)zq��`�V��ZĿ�fȡ{)�?Pڞs'mN�=�=�0�VL��<��'9D�O~)M2���I���	�|k���=���\r�&��y.�m6��㐨����z�HBo���DJt�����H^�V%Mm~�����c'�׸x�yJx�W=��?��Gt�l?	󬎖8S}%�H�H�9��(*}Ͼ�m�L7��F��Y[3q�*U�<d�!5s������뇏>�E�8� G�"m	��{<�^��\*���-�]%�l��LV]s��Hx���4΂��:�M0��at!�0��Lxr4��O|���˴��V��MsI�g��|߰��윜�0�U����x�d~��_�,y�Dp�=d.�G��_�.L��l��F���ȫr��E6P�X�~�S�-0kz��������G�{ھ��z?�vIK�Px�r��1��~YV�66)�c���=��n�s+1&�F��̅�$o%�E����vI\�&���{��@1e��ձѧ�n����:Ε��.)yOY��Ȝ8R�P�[[�^%��x;�%,����u�rd5�`1ja��+��l>G3N;&��.�7��o�����N�,&r5twa�g������y|a�ovdҰM�ʾguv�Z��6tW9��wYRr��U���[uX�R��vY�,ж��ps�2� ;��Cm�Q.�{3P�e򂳃4,e�*m�ҝ]V$��%���g[4�.�R=+�FhԸ�.�.�*VAl�OiMiJ=م�Sѣ	�«��걕��uh�� ���4��u�gY�e�.�r�fV��K�B���cse��Aha�Kʋ.�P�}T�h�
O9^�C^ޜu�%n	��Bܽ�%z#	��]Ӹ2������r�R�{�1Y3fs6	�[v(�s:����B
ˢZ�U�)��ɓثI����w�Y�െ�<�H��솵kzn��b�;Y��,�s�[���s�^��s��faz�!��Gw�$����D!!%��oЈ7L�7n�M �K#W;�n�md�b�A�$�e���}р�$e�ݕ��y���l>��o&����A\�u�"�<O-�]*��'j�pG�T��WR�p�ˣ�E���$+(�ħqwT*�wa���:��T�ۭ����s�Q],�Ri��q	���оx���|ty/�6pw��a���j���Ħ���ꨎ�>n��=��@�J����ܓ�u�{
�:N�{T�J��h�㎏,/��^���%]K̠�.bm�W$-��|5��WwE�m��dI+�t�����ҵEoW	:�����h��@�5 �.#E��S6�.]>��ށG�Yx�_3�5�,A�b��md�zê$B��v
�OV��A����dcU�s\�F����e���N";u������:*����6d���Y�1�xƝ����)��ݦ����kk,\Da���Ew��-�!T�^�k@��GF�y�@6�X��p�Jv:�z��䋭	��kR�W7�5�%��fp��Y��^�ل\RR"k�;NB��ܖf��zV�V�H�yy�
,m���f�i��M�s[�hdn��&�4wҢ�o3S�T�4	���릍:Ə��׮e�]ma��(Txe�=��ʔ�"*z��PJʊ��!Z;Ak~�ݭ�̓�4�8+�:��X�}�+]ۄ@N�ΐ��Jm�j��k�ˍc9k���,�B��A�7�Q�j���d�&ŭzC�+�ɼ�t�1k�t"��=[WI\�:f�FnZ�לv�m(��(\z�`ڀB��t�j���[�ovmC�6�&T���i��(W,3�>��<t�+�`��ɍq��3{y�JR2<˵�Aˮ�**����LE" �Q�r&\��^�K8�M[�L{����SJ6��<�<9y����~{�"��j�)hh���* �����)<�L��E�g>>=~=z�z�~�_������~���
J ����(�*����

#��$O�>?�O�������~�_������?)�$@MD�ER�ŗ]��}�CKIIAM��@��
�:T���QCM@RR�J���f��V�Z����4��W�45@P#JPRPrt��#H�y�E+A�P5�,kM�A^�`(b����I�*��$1EE-KAMCKG��< ��HQCCT%%D4�EQ�æ�A�H��hH�(���*�����B��B��*��t4�P�P�T1)T4RD%%4�X�!E	M	IDM��5������]������\�t�m��/˺��R��Zӷ��<sZVkUcJ�_�K��^d�|�n��g�vvW!R�M/%lg�*������k��^^z��_�}�����Ǉ������_1�{9�(����B]���ȥ�d��_Y[�.�V٪�-��!ݸ������in�Gu&��r������d�צ�myŧplFi�Š�1\У"��4���Le�A�Z;92�߃�E����8�b��1��^��瑧:�����ZGD���;���Čo�fs��|?A��d��6���,C ύ>,8�~_�;_,�o4	��� )1]t��+9�{3�w��J�:]�%8�5r2�"���<���6E;ǆe���*:�ز��]ƕg[j7�ix�F��:AƜ��%��RFiY����,��r���1������3.�#��y�]_�~>?�E�b��uޘ��z}'�:�B��K����c�d�C��67����3#��g!}��JB�ps��xN��;!�8Ʌ�]�-{�(��֪��a~�r��Cj�,�ո��]����s-��}�q����R.�0����f�7ҏ���9�Ԟ����$��~��]{Q=�AU$��FͰ�;"�t��yၯ߂�������Dmg����@k�As�,�[���C�s�ti�}�I76�l����߅Ѽ��u����p�\y��k���t`����A
"�\�,q�Y¾B�,s��N�Ȥ��Af�����<j-���.� �j2�&���c�) kH��s�fV��i/�X������\�s��~���}�s���9߾w�m�09��y^�&��8^����qŠ�cL9	���#�N�<a-pb��,X�jf���;b�)=���m.��9�o:���	���Y˰kj+��9VY�D�օOO`��v��^m0����&@Y��Ae�/E@��`�xwd>=fU���4�5��7����	��)�
Kǥ�]t�t9>��|U��4Uְ�ݾ��m�ɍ�z.�=�n����K��Ö>bŮ�Ƅ������s2Xd�ǥs�]����SP�IuO{��������^����]0B��%xk�Y�y�f���?~��VT���]��T-�'�;�0��T���6�U-�D��r�Ɂ�8���B&N��0���d�0^
f�,�����w:u��Q%���[�"3��_ŗ墔K����fyVXFA0��柄p�je킊�n�=�n� ͋O5�2	��yt�L��m�lg�*�!`�E[�;�NI��E�d�'b���L�~�P�?��/߱��y��]6��S�\�׺S�Z��]0���q��)k}ܮk�Sz���D�N����i�T�V�z�_R�D�P��|&̈Ğn���4�=�V�;kB1z%����6�P�jW#�U�pxӢn�=b���6�_X��92_�Ȝ��-�<Ոu�Ɔ�`� o�Ȉg9P-������?�=�����{�>f��8+��{ƭIo�U����n��H\�]F�P�!#g�\��\FnV
���};��-��T>׶)�8Bli�	��#�k�%�j�����M�z}hO�y���Gu�%��Ͼ�k`0����XQE��Ͼ�C�W��c+_|Am)z�	�31������'B���I~�	�g\dR2s[m�g�Ӡ;�
1�:A�m3<Ӕ��::+����	���B^��ú݇]��؎.G<1�+��L�R�s�_<y��w0�[��e.ڪ
�)�͇Lܢ)��}��>�_Qw�y.�#0���L�i�n�NX��OU�pª�vu��]H3�w֎�>���	�������%yf�K����YPX�ޞ�����Gp\F�\���B$��-���^:W���"$������r(�*�=賡� cn��R�So�5t���.z �b���8�#Xt����\:�0�ۙ2Z�M]g+��2�m���V���Wk�*=�����w���@A@p��}��hV��uc���Γ��fCu7�P��ӌJ�W�N��9oS�o�D��� �v����f�iL���qm.��J��}D|�tw3��/�|Ҩ�fz�^ͱ�%�8LL� �z{wc?0rVϖ��jEq����&�l5�o_{����xT@�����EU;�ϺQV�Zf��LSg�8�ca�u>]�q_V����ڄ�ʁG��A��azm��h/�5��-�	�Ї�r^��_gג�oe�c�^��x��q^:�ϟ:;[�2��7#�e�r��t{-�;1�u�� �H���Վ�oP~������$?pF�=N���U����2ܲi��)�^������hG4��2H��IP�!�+��C��5����d�S�xf`:�X�M�v��%�<�y;�<�楦f�S����??��)z�O�#��~����=��c�����n�-9�f��h!�'&��Pz6q=cռ*"���[?�}�X�^����VGwn-��Oݕ��Z�V�V�4e������MK�{�Ms��ǯ[ռ��������uS��.3^\��x��F�XP�T@XGn��B0�5tB	�Q,���%Ѫ�<�	).���U���Yv���|�v�m��F��\�u<k�fL
E�E�}�N��1�ީƼ4�٧r4J�pn�ʵ��nmK ��ǜ@���*Y��82�},�O�����2�����������;���%��lǷ�5����/�ii�R��W���&[��"��Wyf�c��a!<�Ȣw��o-u�+M�.�X�Х�:�H�W���0��Y>/��n�GL��(�;,u�-d7��̬[��Lrk'\
�p���vQ}lLltqrU�q��UH2C����� }�|����Ǽ=�xN{(�+�#Wcy�k�����F��}��l!#��Bm�����Q{T�F��O��1^Ԣr/���s�X�PO ����ux.�a'�?���1������3-t�!�Ll�A:�u���)\�~�<��nrF���ߟr�,K�&8�c^C��;�܊�[���
��5�M�w�P���`K��ƽ�I���&ޮ��������!�k�>��-�/"��[oܚ#�����y�_KԻk��K\�a�Ʋ�����3�|_l?�7?S'1�ۯYK+/n�������P���<���Μ�؏��Dn���pǒ�
��r����sz��^�Z��V���S�"��s��@i`���#���X����w�k���Ȝm�.���qRiީ���Q�gd	�mb�C ��~U�Z~��$��M�Ϝi:��l��HAM\�d��*�=�����0fm�L˗P�й�(��`ˑ�i��5���6�hl�w����B1�*"���TV��Qۊ)צ�}]{��8���rb�Y(5 ���<XٜeC [:~1.Ϳg�����LU�{��.��^���>�@E���in�'U�S�80�c��}s�vu�sv )�6+%�m�RX��i]3�M�i�ޜ���i���iC��S�u//3���$ؙ��EAC4ɕh��on����0��t�>�ϟ9�S��r�g8A���������R��g�z�ُ,*+��m����vo&�P%�y.�c�g�{l��1������8��T
b�r�6qt,D�S��N�l�\�:!Z��):�buB��x7ղ-=�kX�q�ma���q��\?P��x!7��s	;^�7�^�ԙؘ�d�'�Y�v����ʙ=���*mU��6=6½�Шt�z$� k�����O�3�:�+0xF�4<��_eF������&�q�y��s@���4�Nf�xa��B1���?uS�zp5�u��s9A9н�}O�2�;vL���6Ⱥ,�f�'f��ߙ������a�7�O���ׄev��S����2�y�8�>�oyԘU�\���= T�4چý��J�zĢZ�1ij����à��`鋸��Q-<��F����8�qTXPY��jº�u8�6%�e�Z�jx��!�k�+{p���HA��ͭ��:�9ꁭW�E-s'u��J�'*5&�6&`E��z������V��踏�{�M5��]�\���ᯊ?-˿�y�];تOL�EZ�媵��'�[��t*bn��7���Ϥ����mřI�e�-2���T�?)�M�P������knM#}SU��YSP�B��u=X�{t6��v`�v�����+�&���X:̀�\��Bo�>���篾s������*{�TL�*�+:��ގއ��7oiC��5-�܅yx�+��$�0��M���j`��ߪTڎ[�cN&m/KL�l�;)0��$�0����;a�h�c~�t�g/\��d	-c�2��7P�a��O�<ۦT[j͜�3c�lC���Ӱ��U�6���%�8uq�,u��f�4�2*ϴB.25>���{k͍`$^A!�vA��HB�5�����A�Y��]��0�9es�:)��>%0���q1w5�bj1��xeT�6�k�t���Q�Wg<N�f�������"\t����~8}�4D��h>_����R�ί�9Q=tm�Vh=��@#��X�R{��`��z���S�; ^�0���!�eN�{X�OqnW�7Uy�o#YO2��)�P�&uނ�<��N����~v�)A9sߗ��󦃈�wT?sY�P���XhWƽ ��N���K"�=�ʒT�S�_8���N�����Ʃ/�~3s�)�����d���^�!�}|$J�����]0HԨ񅁺-�ơ�`%���e[|�{ϝ�L�tc��sr�;u�᝕a���xA�S��[m��7 #h;�PzL�VR�{M
��a'��1eWCR�vW,�*��W^�ݶjN�H@젋[�L�!hI�iA�����P�gA���}�7Ͼ�O�����o�?�
��D��Y%�sו��p���L�;65�M��7g��
60�wGt�Qi���m�E�����J�T�kг=�EĻǎ�}�����֟GZ��SE�OIa�C	���O��f�/,��<�m�r]xR�^�oX�z��$sP�������􎀎j��~�gB�qR5Y�-'�k��5CsՌ(���ް����.�;_ܠ�ܨPur��=����A�{���d3�����ƝX�ۯ�ʓeO��S�ǡ�9��3g;�����|w3�+7YߖA�=c��I�^Ļ'ټ��={(�[������q��LZ��q�Ű�e]�ײv�������%�[�a>A�8��7�r����P~�3kCO���H{���c��l�meM]�*7G��eO�����dK< ������{d���[ѽ�����f��N��m8
����6rwU0�둁d����O��o#^Y��sKO�P�qb#۷�dd?��}!��,��'�ے͈�זN0L��e�����V��	�y��M"â�%>Ic����&9c,4^���s��ˇz1�}7� C{i�t(ͱ�Jף=�q��릡�{�s�"�L*�~��t���g��ls$��ke�m�-U��[{�ѝ]��Nm�3v�1
�)R9������˶3-.8�V�fNw�r�V`�v�("K��9���9�3���O�c�)kK)�62����7ۊ��x�M�9J���4�F0�z3�i�p�Wj~B�t��[�0'7�2���N�)3���EF*��'��9J%��4��#m�ɭ^�e3WFLe.����L��]�F����f���`�_	�"�d��'I��JscT�c���=�7�V��w+�	������8���8�`[>�)f�L�l�0��]��Q���ť�"�\=��UnnDZ�7/|�Ȯ��XsQ����}��l#�!�"mNJ���Y��Oݎ�l��r�L��2ty����/IE�������i����l�
5��q�/Ɩu�:�v�yKO:�SM��F����(�R��^��w?z�k�4���61����p�rںuz�|u��P����E7P��ƻޔ���kL�z��S#+�b��{�~�Ƨ�}�Ji<	�<ia�l��g�M�ä���=K��M�jÙ,|�;޺ǐ�O�j��1���T�ɃJqq�3�M�4?���dd0g9g!�vֲ�̞���Ѝ픜��0�g�B�ջٺ(����_���pjf�_�$�_���ȿ��ئ4�2k��צc�W����ڟi���L�&����K�O4��&�d���uo]¨����n���j��l�+�����N�8��������R~����?���������:Vo2��[����	���Z�o��C�*�,`��c��#~���d>�	���ü��ö�w�	\f��	f-<c����_9���%�q.9��0����/5LK]�7�Y�����i|\dz �j��{ҭ�(�A�
�i�Z��E<�$T<�-�c��H�xɥT�?!��h|n�^�����kW��0?RA�k�ɻ�d����=xf�2�ΞԼ��h˺6/Z]+V�$T�����,*:TV5.��X;'�P%�y.�g���|�*�on������}�p��B�Iq���ֺu�d:��tc��):y���.�Vfg�+�E>�tXg�1Ī��ŵ�78�j.P�ށ!�z�"��v�{,�/�73Ȁm@ݑt3�*&C�]�7Y-\���}�d[�'��]�6m��E�*K8k���yk�H8�rN���/<�fk��O��1;�%J��ֱ����Ȣ�䉫���/A�m����D�$F1��lZ�!v���Xn͸�N5�΅�	eB�L9[�l�O\��"�x���mx�T�o�xA�r/G�㊞=�Q���Œ;/1j N�[*ӮZ����=�r�6��쾤h�P}tQ�(�ώN���X���iV<L`�T�B��L|�=�G2!1��26~�
�$�6�ιe�σ�Y
��=�QP
�o{��t��rʇ)���΍F�2��ob�ga"����b/�9�雊�-�J�E��gM�Hl.PՄ{u��Y�&h�꣝2�r�g:Yǭ����@1���X��o�z�3V;J�p�|V��Dr8�6��ɼll%����Vwڳ�ͪ:��p��ջC�'��u�n���!�B�M홂J�S�m��;]�K��jn����n����˨������'�<��9�B�tAf�q���1�#fɏs&�"�����v�K��ne��
�+�c���hz���y�Cg]���U�7����FF"�7 ��k��R�%��Ɵě�VK���ݑ��N���CT�%ԣ�m>�ݳ�=�^�q����T�"��llS�9�衭��틼��[s��Fr���C.�-4M�nM����e�	|���{\X�]��,�d���Y�{�꧷��W��De��.��qy�0�X��^�Ka���0\�|�oX/� �s��[��YqKLr�%��v>�*i�WG
��ޜ�T� D���U�����Q�(�R�˖O��FFK�b
��{�g��T"lШ��ga�&��iܵ�;����8A#���CH[ڲ�#�xE�v
2�yKRyn�kh�^��~�΂k��k�_���R�lw8c�ޟKkeN���:��m.y�&`����ۧ
X�a1��ϱ�hM��Mn�-�����dӹ�;\w������%�u�.C���	�V�3&J��a�6]�䝑���M�ss���[(|��^�	ga�q(�,
��L0�Ҳ�i!Z�}����D�c�Pܵs4j�wI�G�хC4��6wMԂ�Y02�4��Σ�2-����dE�^�Z�^R��8G��(o�O�ǎOm��:��&�HDVJ�-�|��ɚ��Պ�g%h��AvX��H�8�5V�_�#v����Xf��$�\1���q������b�Fej�Hk�ZuA{�^k\m�g]9�ީ�l$���;��	��
k����M�fЕr�z����@M����:��5,�nn�uMi�)�	�g�d��x�](���4�/$�;WwA�Yx^Y�Ȏ�KT�S²�3����was�[6�2�ۭ������ ��HY� ��p;nT;Hƹ�6��K�t�L���F�:2���+* \{Z*�* ��=!.R��S��M1r�RȪ�*mP��k�1�3j__#*�,�V��n����fN�%!��u��:[e'#&����'k��R����)�k�=�Z䜌՜�������כ��_}�6�ׯ?��=AM>��>��4�%*QQP@4�����z�z�~=~�_���������J)((iiJ�*��������$'=z��ׯ�����~�_�������b*��������!��Zi)��bo�2�II�!�AM6���P]���Fa����[� ��h���:Z)�����(*�@i���B�)J
�䇨�R1%$HPQT�2�c�14Д>Z ��8�:�i�v�����BhZh�Gա)4�yh�� D|�d(����{����ģ�)��t�jfui��I��	�t������Vx[��p��t����{�׾|?�)���D�r*��?�?�Ͽ�ܬ/������/)���
/��	�U�\��\��T'��ܰ���w��a�y�Q���H��'}1�Aæ^d����y�U�B��̝qw�QaAgO1����ST�@��fuS)��5'��:��mnk��a1����zhZ�9��:*�h%��>Ub˃W�c[�c�T�E�~�V�9�8/�~��~F��fY)_Z3��wqɌӽ>�P��gua�Mc�wh�jXc�(�x��0v��w��!0��
�*��HL�R捖�Sop���l�l�e8¥���ג�v��-�8�r��yw����f�c�eft[�c�	�����>0���&�m;Ǿyހx8(4��K��l��1�}y�syR�r�xj^���"E�8�W�vR{��Ƕ��ּ~!�vA��HA2��Mm=�NN#�=|'e�2�z�m���\9/,��'�`d�d]����O���UKcP�B�b�g��6_�5ѻ�R;U��:�����/}Sr��E3��pL&v�����w(s=����^��@�zwp<�Cr�;�i"�ǃ��u��a�~.m�B��f薪���r��m�}��E���މS&=Nk�ݱKţnWd3)s���4�+Ӳ�}�~����NK-یӾi�Ԃ�e���,�Ty$/%}^������q���
�z�)���E��N��R%�D��*�v��z�o>��vA>6c�/�����Wkc6Y����[Իͤ!����ђ�Є�E��*S�!E�63y�ׅ�;͕�(&�,&m�4�*#�fkw똵5�}S��C8@BE�H�I�1�d]g<S*IRaO�|��!�Yl���*��:�z�k�nZ$(f$D��.Ct��H���$����LL��#^X��+��,�˧��X��W�2�5 �^=�zh3dy���uz`&�4(��$ڝ��n�k{QP�Z���F�ղ}��E1]���"O�kg�?��B�t����y~�'I`[p-Q�J�<�E�k{3�^	�1k`�U}t7�α�6���@B5�K&`g���_��3|�����}�9T��~�MeJ���^�I7�8�X�Tx��t�W��~���vB�:
��0�܆�f�R�������0��C�n=i�d�>4��(�|�S�ǡƽ<�ܳ��qONHi�&�.-f�4�2�	����H�Y�D-��r���}�}>���-���,ji�z���2���ٙ�{�PyW1f�p��Ȼ�N% �VN�aVu�c�-����2{�\����6�ƩP)��Z�����%X�!��ȕbi��f'}$��ֻ��Zt`�dK���ᦥ�ċy8VfB9��&���g���Xd4p+�	����
�������]+Q����ك���	�����&%��L$�����{����X8�s#:���^�$9O8&B�/��[vS���CB���i/��ӱ ?VD��" --(d�C�$�%�ލ����b�y�	U�}O�3�w�3JgXK(!\����ɴ��6����a���	�%�4R�i��j���E��F�j�@�ƒ��m������	�$v��l�|i������gw[���y���GXN]	�>ja�:*�q���N��lr�5,SI�Һu��ǯ[ռjj�:)�j��W��Z4��xŠDK�D���Ed����D �/YxY�R�e~Ti5�vJdT �����S��`>7L�W�\�8��ʴ�+� ����~w��?x�Js' 3��uv��I�@�����[��S'ȸuC���j��mLpe"�Y���a�J�o!�dN��OfX3n�,�Nb���yim�F��}��`���"Su�����Gz#eO_vT�2��`^K��|�t��.B�R�%���bX�^h�h��2�F��c��t.����0h��3U�y���^���M+o8�t�����|4��:9幇��9�l�X��pa��ۼP*ؕ��;`:���ܫ{��R�����7F��2�wW<��xa�gC�2��G3i岕卂ٰD��#M�� ��Fv3%���O�s���Ͽ�wO��?����>����X�9�Lo8ֵ�^
��^�����:|<�E�xQ��ֳz��h����{]�NB�=��TK�n�J~1-�6ⅳ�t�VoIO�~Zd��Җ�U21���"e��f����uݚUCqa�9/0�Իk�ޚ��a������O��u7/>�hd�!�o|9���F�>���z�E�1�^��~<`h+؆-p+:�?��l�aƗ�]y�n��ץ�}<6�ܷDK�h
v,*�X/̢ac�(�q�Xtu��s�/{��Hr��e5]��eش�^������f�|e���g���TQ��&�2�Gv������UZ���j�r�������ؔ�`j]�����o��)�R�U䛉�|�;���(Ћa{�lObj�ʆ��M�H8u�!-�-���γ׳gE��8f�RɊ���̾��+��_����)���O��@Qr	�yo[�]'��׭@�;��)���F�.C�l��\ή;�T\>ۆk�\��Iq�1<� .�d�2as�D �\�t�*Wu���[��3�^a��5|��iM(�pt�2�eoV�w��Y2JP�[b�����Oy]�8F������#�'�jIӣ��Jt𱢠G5wL"���z�K(����1��-��!�φn8���si�����3m���������i=c��u،�i2'�
����������z��9oR�"��v��n�Q6�:k�ɼ���0n�u�^
 ���(�Nl�B��U��ѳl'�-�tc{���p��[����gSEewA��_K6�#�K4�Q��u��r��I}�Dׁ�8^���N�˜�݇������6.d!�'��8�X/�;vL�S.r�^4�iyv'�]K88�2��OM�c`��jY�ל?4XpKȇ���	�=<hQ�4�Uz̮xj.S���$㣟v�[�Ջ��o�;�����&�}�b���nn�qz�u�ul9��/���������Z�����T�h�D�v��+Aiߊ�������U�z&�{L�o)6Bz~�������F�^�1��B�zcBxH��r]o�ծ�@I�,��38���0��Mۼ�U	}�j���6�����j�qT�]5��ݢ�q�nj=ˁE�3�I�4����m�}Y���r�}�� ��óau�6#�gex��9�C���^�h�;>�(���_��/��c�*��5�7z�Ү����Sx�_W��K�[{=m��8�x-VvU�RS؎�!Gp�+��{X���Z�)es�ծ��Ff��[��ڠږ�9۷Wk������az��ՠ�"S��������0�����r� +߼�����x���&S
�;����G�!�TT[#c5�L���poH$=%�A�L;?v3��d�.�m��r&����ܴ����E���}�<��3+,��U��2���Cؼ9hSo �'����o�	��z+A �h��!ZU�q����<��r��t?~�gv�ЯcD�җ%���<U�)��ۙ���N:�5k(RJN8~ޘD�㦽@Uj@�.��:`���`��{b�߂� 	���ޝ'h=;���fa���˄*�|��Ƥ&��T)=�]�.���z�oMl�zdss�n��.�`�5����.���>����D�V^%9�
��5zT.�d�=k�<'zf�����&jj�[����
5���*` ^�8#�Ot�N�1�d]s<��$�0��ϊ�A�}���5Ke�nz�K�}hz�ܰ\��r��H�^���讈���~F�]t݊�|T��0�D�^�v�^"؆.�nNe�k�w؀�M(fƘ�	��0t�o�i;���FCb�˩�Kv�ٞ=�}5��WN���a�`�,k�t�~jN%�<v찎���t�O4��_ɧ�,F���2�R�Vt�� \��d �٤;f�V������d���*�zi��܇�#5�~���zv�jT�cU�=��l]����d�6�4�X'K��mTʰ\v%�*.6�K�
gt[x��v&����}�ؕ���w.��=���pۖ����� �������7�Ec3�Ǖ�-�'h]�r�^Y�s�+�K׻ sIzp�7 8�#Xt�y���%�� ї׹��Y���XO��bYdl��[�0�=+^҂^��
Q̮a�s��?OH`�6���g�z���Y��}c?�@��O���>KmPb��ȩLHeO�9O�����1���_6\�ޙZ!���<9`�< ԅ�Hv���-��Ն�����}y9z�yw����-��lV �5-T�ܞg�qkՁ�;b���w� ��ā�ˁ`K�:W�>��:�L��9מb��kڜ���:�L�8HK��K����?_�D�ǐ��҆A>z�ʞ��ޏO:A3�d�1�k���έ�-�Ӵ�4�,%��R]����z�m�{^Y��sKJ
y��������S�;�q�	���н�mEK6����	�$v�����z��]"��l�kg�=��|d�t���3c�5����^���*U�������o��ɪ[� *��%\�xP�1���rr�rMeB콕Ku�7;��m��h�a��d:;��1�����N4Q,��)M21]�ݑ\���H0k]�\���s��^�	��2����ev��:�CqZ�_�����EV����/[��&և>Prh�I�����t�{5S�x���
�a�i�Q�����]�v��!r]XR{�;F;����<��˩ٽtC�C��[�ɽh7ޯ}��� P(�
R���i�/l��On�!@�Q%ٲ�| ��y��9�S��gu��Qw�9�1egd��b2���Mԑ���nO3c�:�tzq�)K6��eF�죌ԨN�<;ͫٝű���A*����)9\�$��a�A�������G��M��l��4Q��Q����/�W����1v8�_��}('�K������I���l�j��ng$�^2g6�3a�2���H����;�M�3�k]�^+�d�c/A(�zO��Ā��]PXeފJ���71��"R�v?1�B��<�� ��WTz�}Ն��'�Y���)�e��A�m��(��<.�5(M�;�r��s	O�GW�&N���P������O쐒	΍g�MSL�����ٸG�Ѫ-%������5�V��~����.��k����6|	|������)��4M �q��_��j�{�9�|������LL,s��Z\.U�;O�t��p�Ɨ����"x��Þ2�ZG.�Gh�/C�m�׶D�����Q��㬯���L�s9��#I?��n8a�ޭk�j �x6U΢�k����b�N�i����1S����+���f���mˡ �@n���er��ow�׋U�3+-�ir�-k�kUl���ѫr�4�^�n����!N�(����q���[�k���7�� Ee�%a�7�&,��Q���c6}��Bk��y�(�A���i1��]�=��<7��a�s��\�&~�����΢���0vy��Wp�i��D8���Y*�BFu��"Nw.���޽dc�C$c9y�zw�
H!s�f<��r	�y���O�ga�j^��#sY���[=��6�d�3�@tv>5��uW����Iq���ֺu�PɅΔ�
v���0*^ c��1�htpf�CQ~/<��%Tc�)�nM�uEê�D�(3�u0��c�bz8�nv�S1"�Y�'.�dQJ��b6m��ȶ�C����8ܱ#��DM��P���(rf�X����.ӽJ�,`&+��Б4���*	e�A���Ӯ����ck�fx1ac e�0��pG>_Gy���m�%=Z3l��/�B��6�C�x휖ũTvp��sO5J2��ώ�=�y^D9��.���*D��0���\�Ҳ=l�ӛ��w��KMKǋ�ŧ�O`�����W^) ��k,_-�����Ǽ�|�>�O����,֐��|^Vj��h�ۦ��qQD�m�ǹ�m!��{Z�)�ޫ�cs�'8.ݙf��Кd�W,.�j�� mh�κ��*�\�uN�݀tچ�wV8�O�������C�E��4��*n4���,������j3��U7�'>^o���?��4t�j�F�*a�# sU:�5S�q,'Ӓ�9�}ai�Zx�����N~��U?�u����9
�zs]+ϓ����X���͏����A��V���@G�,xs��y���ۼgc8gU/��ח��knrT�]5�|��r�Է5�,���d����vL5P�C��0t$E���6��0̓��v���,+�I~.���L˴�lS0*Ʀ��wn����T�}�iX�i~�=���������Ӳ��Ӱ�Ⱦy�oH$=%�WF\TlqR�tH���Z"ؙ�M<�̀��A��|����!d��X����ze�����y�zP$�o��Uq[u�6�wU	t8�L���)�WL\ �)�, Xt�?���&��Q�F���bWil.���Ov���E��#>ε�y�WB��GPU�0�q�^�����Oذ5��I�SEqɂF�Z2-.��n7�R���Bl�U�	��"S�J;B�t�{�ᦞ��ui�٩pq���m�Aղ��k�H�PοӅIb�Be�/�PJ�`��*��d�:����n���K��^1��l�hapYZj=�e��YMs: ��1/��K��:�:m�F�P����qr���c����t�]Aa��:�R�t$�t*��y*�rt�:XZ%�1��S,��I:�Krm�(oL�V�{�����׮)��7�d�"�|��]�*��Y�n>�sofD��w����7�T�uN�u��V��ʾD�ՇE��F��-Ϡ��::��3aX�J��k���
�+ٺ� M%�x9���L�|O�o��BWP�<��41�/���E
4��h���G�$�87"���;G����z�nU�f�,#�a��T��MI�d����82�����k[}r��k}!�2��Yܧ�Kټ�2��9_ٴ����(�Z�u�f�k��x�e�M�
�ְ��R�EP�v�1S	��2l�.���Ӌ��mA���`�o�����6���gc�;+<��i4��B������	�!��n`�v6�v:C�1o�I�V��elo
�PȷՙqJ����ɚ��m8�Jk^&o6(������Z\z^v�T{l�}"�Ҥ�xZ�w�λ��Kr���K�ui&��Z��3d�m�1@����OK�ek�s�2D���7xѢ����&����N��۰�W{��9�+�UmN��m����C�E��ca �Z��+���w\��*�橉Z����MS=����F
�u��M@!�����=����;~��D846-{2�"���5���8��mln�;a�iV�wf��o���vQ�sV�&̥64���xi��S�h�x�j5W�6"D2n��̖����N���)����]-�
����7r�Hn���$8��r�`.ٸt�6������i�l��m,��� J8U!�@_P�$��vgGg��u�mora�AV�="�ط��V�젞���T:�[3%��Y�UXj;�$2l�Wv�n����V.0���q�"g1^�����嫕\�M�vu`�d��m��*�8֋�]���SVqʚPȁ�N��0�冺�
>�٤9A�e]i�����HkTOs8��=40pI�.����*���u�"u2b!y;,�i��vp�rWtjŌ���n�9�M�nQ�y)�1�dM.����En!�bt8`�eзY�%�.�Mʹ�����gׅt���خ�V�� I3�-�Oz�Ԅ֙�˳Paғ{;�maz�<r"�f�n�L�&�R�U�_F���J���-]^|�vIO:��s{�]��)է����䮹�]ʝ�ԫq���u��Wv��VA����70�"[��Y�87�
�չ-uBvS�3��"��y_xn��SS�@ʟ_�^��+�Wv�h�4��iՕ����AM�������;|\y�#��`ڗ�:�b&U��!�㕙�lm�}2wHn��%a��A��`L�{��N{ԙ`D��_$)E��q`즬�ZqDj�m���zÙc���6�Ջ:�-�g�*��ϐCRCy2�\"m�7߯���s���<�����I��~O#���4%%)TL�}>�O�������_������?�?E#���w��g�ǯ��^�_������~�_�翆�)(JZD�JB���Wl4~����<$䜆��F�F�M5�G��4b�CG!/3Ƞh����AT4��
Z9)������1Wa"
V��ILAQ!Q��`�T׭�F����H�ESMU�!�M%!EE�@z�J� �^�=G!҇��}^H'$��H'��#��\An�%� �(�vx�	޼�v+�5�s\ӯ~�G�Tmv=9��\Χ�ï]Bٴ7��[���7�wYڴ�|�h8����?_����p<쵞Ջ1��u��g��^)�c�x���t��z`�o�$_��L���E�s�2��}�Qj��g�:D�)`�`.)��7���3k�a���A�/��U}E�AȢ����nF>����0�R�~A�Su w��W��x������~d�>��&>8bD�`茈���^v��.�QF�^�b	���౥�a��㩄D������1g���Wg�A
*��eV�Z�S��L9�+�[�	Q���;�ի����4����8��k��hH�5��h��h2�p��C�cx�얰93l8������I/t�J9��3n�`�0����hl�h��5Q@P��ٵ��d��mǽ�]Rc�GS��N��g��0�3�]�]]\�3b�}5�W��H3��/Uyg��o ;fz�Q~��=%�Esklt̐�[a�~�����f;�|?Q_���I�[&���z%�r�����E��{�J��?1����^���v�s:wQa���MH���>/���6"���M4JZZ|��i��I�b�g��0���ȫ��'�m�v5L�\����.��k"�Ϸ*�A���^��Z%]���^���A7Bim�ˮ��v�j�&b_S��LN���i��.QŒv��1+��L�VG��9Ԕ<ʻ��ˊk$����>�u1̏)up������ٷ�'��3��w�����������\���֟��f����K(!�<�Un�.�r����O��?�����;.T	��͕��A�Ȳ����j}%�^�4�y*f�;(1�,�`����Y���LR0��CY��{.�Z���\��Vj��V6���D&��(2e�7��������*����c�� oH�u�|w��W�f����vA2Uss�	ƎQ,���d!�j���3y�^������U���"[���AK���S�eLs7�A�y�(��\6G>���s�c�Q{�F"y��Lk�L�����kz�\:<�@0-�(f�~��v��tɐ���=�y\N0�fÄ�b�).�BTi��)9Y�0�c�h��х��<�>�<��;�y��gac��L ��<�� ¥�NBc/^����	z���.�`y@��[�uٖA)�v�{C���!0�M"q0��^��M7g)Ʈe�d�c/IGsד��튈-��n��;��E"��L|�� �fHT\��v.v�����R)�������'浦M�i���Bb]ud�z�]��s�Ə��!�!��I5fzJ�%W�&kn��K�q\�����_r5[C.��]&8@}�R����M�U����6�<�t��c[d\e-Ձ�3I����b�iuJzk_=��Ln���v��Q������π�|*��lrt��U�����y�v���v�tw�'�B�]����GV^�
��/O�k�Bf�e�sj_F�-V�iO>�����]a}Ph��AZ������k�����'~�ò���8�7����=PU��pS7�,8���7����/�ܱj���C�;V�l9<�bn�ˇR��
O�1
���t���8�<��(�w�˟;ϒ����r���`�_���5�-G�eo,�y����X2���3îu��:�fϯ/��ՃzM�W�^�g^�[��"���#�-��F�+�Y�<9f�R�ȧx6��!:��cYx��Ogw8�jt+:Y+�sՉ�铡��n�1����3���42���=;�.2�BOޡ1������ﲢ��t��WY�5e�e��sX7z�z�T�tL	mI?��g�_[%�eǃ3�P.��q��ώ�1�ˬf�U5	�+oTt��j<�(�@�I�:!j�J���
j[s�]Qo�W�D�s�7#	�[�܀ў]u�P��L�.��e�����rȺ1��J��UE8��l�1׶�c��ӧ;+-9���5h��l50V]vP�w(��S|��)Wb����¢
���w?	{}��������`u�a�DW��6�� ��qֽ�m�o\࠷�t�uӖ��D�)�·6�c4��F���\�;���jl�3ѐϽ����y>�}��y�fY���n�A�gi!���H�̃H��v��J� \&){�E�h	9�n:p�n{7�eP��2o�/'��6��[���c;_�`�7�%��m�%=XFm�tY�3U�l��k�B�Djp��0���.��?<�{h!י����z�����"M�L$ٔ<1ď(�خ��ѹٸfސ�)�v��i��(�ð�O�P�~=�@E1�q�F(A˝�
�u=�y�]y�xM��4XRΞcV���k����n5�r[��[�`LU�q�s�L�-'�8zEb;.6��8��+������q��M<h%�+�!���J��g�7N�����2�B�s@L ͵��,5�g%@�e�X�9C������e���3����g��*�������w^�P4G0�<o�����fI��v��E��Q)�wn�A)�m���*�N��ӗ������9�ز�N�5�LI��y@������ް3i��R�����Z���ժ9��.n����ge��zc�&���π��B,�|�I�U�����}m�����:�t�M_��G���0�ȷm.n50t�!�3��++^t�xރ;�H���?x���B�z���7ƇW�w���"H0oІ�"�y׍�[�q.�
�i��a'�rK��ɺ�lŲ����6��w#ǚW�3G#DBZ:82��h��{MSy{�v�A6�G��3�����33���SV(����m�*��$ ��5=˦��d¿TS;��X_�!ܯ+c�\Y�P�s�=ݭ��^����4���Ƣ���`� ��ȕ�J��E�'�X�!��lK<!g�Z���}@ⷰ�=��h��(q�dcq٘nm�BS��BeK
Or�h\�^�u���iž�.�:��[��ZŔ��r5k�8(h�^��|	殄%2��)�ʔ�5EP����K�ܜ�ؿL�/���{
��%U
`���F�v*G�Ä�O�vd�8�%��/Ku<�j�3:��N�-�b�,)�/�Pw0�[Zvk�D&��%�n�_	������v�Ë鼛�V�5Q{a�1�W�bX�ΨkL,ɷ,��ýg�|P�f֨"-��&nɓ�r檦6�T�ېwͅU���t�Z�O�eAc@.��IĻ�p���``鵘ч-/,Ý1���!��֕1)������'(]�&0�Gs��t;�����z�<xn@q���1�"��إ�V<F��!0��8s���m;=Z���3�'��ς��O)��y]K6�i�Y���<1�����ף"XX�b�-��{'��i�6�]]_,����[N��o[�if��t�a��"Y�:�P�uP���뒧{[���55�u��%G�u��n����L�7���Xv�,ݒ������~�����C���]����-'U��C�0y�T�����D�!�]4óm��t�+ʓeO�)��h8�k�2�s��$�sƬd+nY������	\<�пy���<�?�輁��~���,YKQ���o6n�t�e�Y�Z&+��Ũu�v<��H9a�����6^��-�ݯsI������ݻ��zC�v�i*Ŝ�z����[�}��2'<�!-,��19��ԋ�k;�Y���TZ{�ݡ�#73M	���rw�|�������R�Gx�b��w%���SH��Q���sS�Oz���IS6ߎ�h,�`�#�sg��b��H��T�NFY����f �<H�x�!ŵ�<�"���V0J��W�o)��J���M'��ne;%�&��[�e�0���\µ]���Zz�X�?1�`p���x)���W�UsP��x�Q;�b�{�5
̮4�݈�۟ ��6��k����9�<���z��1D�f�t�e�BHu�q��[��`���<�(�/���UD��Y�"��F�[X���lz�Y��ŵz�mKT�.u�4�gY;2g+(v_;vR�=���y�f�#K�m�sE6ؕո�Q�� 3��x�$හT=ix+���p|�YL�d�پ��3
�Z!�.��+UY�2=�.����q��I��x*Xb[=��F;k5��<��l�/7���ƚ'��U���3��Ƿ��O��z)9X9�Q[2�\���>j󮆯��Ѩ���mzxj����&01�{<�^��K�ل���?"�%�o)^]4��ꙶZ�����ӣa�� ���9� �`�����xe�Bw���g*ֻe�Y#Xˤ��Ov��U;���[�m�M��z$3�����z5�Ǿ=�}��%~��������V5�ғ�v�Z��h�ŴMQ�1o��3w*�)��^طvm�����7�v�E�K��^��O��pw�p��*�V���%��ɔ�{�}Zfx�X_N��鬂�л����c\w��ڮc��x�x�z��s��B ��)�#̌�,�ށ�+��fǦ���3��#�ڨ�#s��Ң�������X@�+6C����BxėbZ���y�B}���r���S���@rU�1yT�������ήb�)͌��^_P�ޓ��-'��[�4��QAJ��8����GgwkO�o��nX��M�0( �-�{��ϫ�6����>h����Q�K�T�b6<5�`j�y��=oY�H��j���8qh��Sis��w�c{�Ң���2� PS3YB���kS���V*�	R@�l���{�L� ���c�7��=���]��Vҕ�rokT���f�[�{E���]�����;���ߪ������,a�l-��gY�6q�dgO���R�:��LFB�?�˯t�i��f��'�!�r�ȋ�ڌ��J8�j������v8���s���`�.|�/%�i�7M�-�k��ޯ�լYs�@� �^�(L�b�IL�xK���p*Z���Ao0�G3�=a����y��Bas���&�KsWD&I��"S����2��)��]�ٶ;"�u����u�Я�=��j�����C�G�����!�t3`l��Hޅ)� �b��E��4���Ml�.k���j��޾=���u:��H���#ZD:Nj` ^o�K��i�%=�Ⱥ-<Q���xV{AӨ��Q�����1���部
mxp��p����E�ޗ���_85m$�aK9^h�g�;}��*v��W;�`��0�|��{�C�o6�`���e~�Ѿ�����T�K��ο7Szg�P)t�8� �(���<�=W��A�Y�9R	�@���XtZEN�~[��]4M�w~���L� ^��̜qC�Jװ��֪9�������ᅌ~�	�A��@cB�Rh-��p�鋶�B��nS�dج�gf�`���V<=K�ʆ=q^v��p�b�
�m�E0.ߴ|ˎ�].}/��lA��a���e�F�-��6$yWZd�b��]�;�mb���>���R��{��3EoU�����IG=����9�]���>>vB�G4���C�+��\����3Ց��Em��mj;����pҼ�P�Ϸ�K���<��̬s�x�M宸���KƎ^��?�|��÷c��y�F<�{i����XW;�;h*��F����.�046�yOl*���k"�LP.d��.J\��/�yx�l�v�R`hl�^4�>��sż6����@�������|=7�����nf���������y�אy�%��My�\e:j�L\<��<z�s'C��	t5-/=Q;6��nB�u5@��-�As���A�z�PT��؂�vFq�^�tS9�Fg��w��˻��[�����/l�#�B��*��K	�"Sm�,S>`<-�ј�7�rO;U�9�������[�<4�����mI��g�������9<�Є��r�Nl�Lf6m�B$Ep�#�fIV��[�j*s��?=5��[AtC�&O"�@"o�z{�Rt�^#{�\-ʹ�G^'��i�EE7PIRaO�|��a=k�ٮ��AT�7�B��g��k�AX!�Zw��X�{$=�y<��o�¥Y��Cۻ��(`<��h�=���Iz%?n����U���FF������S)�,Lb����1� OjVz��0��5t��q,�:��"������[��r�{������͜*ebؼ%ߋξ0���]ctS%�Gw�r����;�B
��	���XLr�};�q��sT�-��P������O�)�z����,V�C� XC#�g�#��1��Lɀh�#zh(lg��<c����3�T�0g��ì~e<U�h39�����W�u�-��#z�BD&��A��W�%�W�hS*�����{�3�E�2wv��&���4���������J�ü��-�2b�;s�O�ٲ�k:m����'�bL�fX
lcՑُ�Guz��0ZNܳH���:�(h���䎜�d�W�^��xZZ|僮��yO���{�	���=-"�@۠;�}�9�Xh�ߛu�*!�_��s����؋�g)e��_�����WÍ�3�����]�ǧ{����[���8S� C_5q�h��㪕�v#O��>2�/V����j����W,��R]ļw�P�-2k����y=�L���gR"�ZF��^��5>�{׶��*f8�7rS�$rC��z���Qx��n߅GHaF2��c.���zvM�X�!�b��i��kx��:���${6�>�z�Ls��@tUD��Z��`D��4�H��_Yrr���Q�c�L5��Vb���&ʭ]B���_1�:٤�N[Y[�t��7�KiW\��eG+Ytw[FT�Gs�ZB=�����t�&Aej�R�s�)����Q�z���J�l�d�Xo�Z;yh����n�RUw9.��h�K�,�MOi�W)���AQW˪�ɜ�֧�i,��Y�6��b<��e3sJHTy���!o^�7R��cH�\%���N�';�XUs����{�>�r��j�����d�ʶ�"�5��zKW�.�U)�u��L�9\r���n�ckkB���P�Lښ�=�}�q���4J�E�f��MΓ�έ��ۋ#O�"�`5kT4FHTĎ�s�N�D�m�u��aX�Z�阈;$&�Z��{*�a{��&]PV7&d]֚�]�F˟P8.]	`A[CI��4n��������'�$&�������m��2��OE�ut0@�C#��f�YN�su�6���5fih'�.�-��'<�Q�7��E��Fghb�0�Zit�]��$N�G�L�竨.�2WZ�{rН|u�(�d�^��G��doa���ԭmp��Su����_'���S#zf]`K^M��t�讚;��D��M�ŉ���9�K퍱.�����2Hх*7�R�R�+T�k}����o��,��Ͻ��ݴi3�	�h�e�X���Y�;S�d����!�[�:j�;5\At�����]$��&���}h1$��EV���>%�V�z��e*��`0�z����צO)��Iͺ�B��/u���R�Pɼ�(��γ���0�]�_f�v73v��U1RPmΙ��C-]vN}���I%�X\7�9t��G1
�^�8�q\�%����T�!���	���̹\�(o�\0�bdgׂ�k�Uc3�2���ڍ�c ��wW.��!CkE�*j36�DLe���n����+���>Щg�(��8
f\�^�Z���M��U��˙4��	ٯLr�b�Y.[`���S1����u�������,�q�U��	�hB[��.�m�Y#��Kƚw�nVA[�{Ky��aůc+/��%�/�)ˣ�չ��\� �>��:_kI����:yeu��7�Añ�d�D��7��N�Mm=�7.������l�����K�´����u-h��z��M�d�G�1OLĀ����>�5݈��9J��;yS4���r�#T���c�����{��6�sL��%�5���)����������w��E�z-��I�fWM�L��Z�;{ m���^���al*ٱ�to�ҍ4�g�|� ~G�R�JR?gl��8�|~>�o�����~=~�_�����~�]���9��h��Fx���ׯ_������~�_����JO��J�A�=�<��t��U6�A�)����G����BPQ�=#h4iNA���9���M�h��%�i)�['�s5l���nq��:CJQC�8�(R4�I��9y	l�T�R%�(iv��j� ��r(�.�Ѥ��B~��:�iB�(
\X�(�md�M|Ȣ��_�O��`�Ө�`ڪ���y��v7+"�(��{�Z��,31�u�#��^����ws�b���9Q���E�w_S���y��d�9�ZE���{g��S���a����()�`M�Eyq�7��ɲ�n9�>t]\*�{uF�L���`�V��_Z ?�\"�͏py�B�����}��2y����ɫ���Gv"%����e)�V�Ъ��Z���l����	���s	�y��sO�����Wk��f�@�����!2O`�JrT	c�Mm~���5��d�:��@.-�ږ��"��U=����W���3/C��>��a�{%�N�*I��a1V9�Q�����/O������\��\wFsK��>�P���F�C�ۂ�D���.�nY'����O#�o<R��d.WC�of�j�X*�a��<��^�i�ڨM�G�;�{�y��HLe�hSw>L�c�@<�(�t�����~� ��H���5���uo C��BdN����Q�X�y�ߦ�!�N�[7����n#O��(���N+���eл�"^�
�B���S�5�Eᩲ�wp���D<�)�K'k������<�����|�O��δ��a� m�� �Ё\���Ʒ�oP�(��!�h��/*����P��`��䩰��n;��R,&ڪv��_]@��=�'t鋠���DW�ܯ}%v�=�,�1h���U��j]�o�ż�w:]�N7u��Z�A;�ˊLI.��ʕ�,}�.P�;��.W�#�!�O��w��W��3��	���2�*�6]z>�d�7���t���'�KL�l���nZ�{�>�^mnl�ʹ����1�(gd$dm���Vm���#@�]�÷6�c�ĝe�p�[�u*M-�ͪ��Y�T�w�!��L���nb��͟E��o�
��<�$�<�T���6�f5u�T��W!;i�
}k��o
���(E��=�Ƚ�\��^N4�dGK<֐ⷮv\�6rwU�C�N��L���e��[:s�-�0T��<�Cݽ0x��'n��@�λ��U�]�m�0y��l ��@�4�V3�1�����ߤ;B
H�\X�5�s��mڋ�����efy��&;�� �Z��=)��T+/ʫ�SW�ۜj�.r^��M$� ���ݖTh(o)�#*c����(gJb����(�b)9����2S�|�`�oe��<�C�#���۲�uj��B��$=���,!z�f�ս6�(1������Yu�t>��蹚��}�HN� �b�ם��H́��ƿC��^�s�8�Y;̎�^�M�=�����I���XS��\�;��Vo.�IG��=�}L�ȧWN���v��i�]�\�%���zrm.�z;t���9�Ӝ)V>�S:���/��^o=�����ȃil����ks�t�a�e5�@�S͔5�����C�*���ւJ��vs^S��DHl��0 K�y�y��a�	��K����Ʃ��w��͘��x���n����k�jiP�����cץ�t�M��`��U3�U�ѥ���&;^ye�/`�5�ʡ��<;����w`�u���6���~�]�a��Vps��T�zJ���N?��⨰�,��5j�XH	��, �~�ӱ����W��t/�a;��a#X�κ��s'W���%�����P�k�ܞ��R+���p���=�4��3��2Z�>�3+��,VqU>bEc��MKsd�,�0z_e�hҮ�n��̍���@�x�~��^bm��L0���;dު,+�Iy�ku�V�Ʃ륝w]����a�'hvP�,�(9D�!ZyF��d(�����<K̓�Xs�Ї)C����8�� ��i׊xn����(E�"�#�5�]�k�3yLV���z$l�	��!�5�א�yj��2��B��m�S����y����#�ffa�2K���w�p6�Et�=�M@�޽�kl�B糰�*���J`ۇћ8D5��_���jtE���6���ٕk�p��-�hg��t�+���EWm��զT��ǚJ�[^��h��dm]��x{"�;8	;02�xr���3�v9®�[S��.���9�v��Tm����Һ�2rtnH�n����ɸ��y�����f��gR [@У�a�'�����j����i��̖)����A��s��C�QqW9�2_l��za�U��`!z�A���$H]^!�_)�t!)�<'6��oE�Kc�t�֞�m�]���3�t�Q����l����Hqm	��0y��|k�=E�ɉ��aX���-���Fߐc�~1�5E��$�@qQ�|����5���Q	�׆�˒Ķ�fFҺ[�tu�n
JK���0�jQu�7E2�-4:�`㖠�^<�M�7�q�R�nL^�p[=��C�ܯM
W���y�ꚗ�r�O�S�%t�~j	Ĵ��y��M7n5ST���}�Ws3��+���[=��vt�29��g,��_&���f���s�����'!���<���;7H��:�>L�Q���zb[�qA�?t��V���ӧ�f_� �z}�O۪�P^��fT[��1�~�_�h��+:Y�>�C�f����J�}��;�����[���|ܳO=v������&H�^�>���vO�����ׂ��'F��O45����2�uY���.:#ܧ��Doo��<�P
d��1b�v�9s�ҋ��*�n��oE8�z�3��t�/�Y.<��tC5���s��dV����O�����'�.�*�vs���>�2�4�o',�ח9]����o0��.���5����w+����'2�w:�v�e�ʇ@�c_}1�vL/C��.��g(h@��Wn���׳h>�N0�����- ��b�)�cb*�"Y�2_6d�L�D��s����0!,�
�i鴽Kս�
���}L�^ޒ��K(!\����-:�fP9[�s���g�J~Le�#l:
����\�ǣ�E�cHԕ3P97RS�Q��l�ۦ72�2��+��:��ٜ���eut��0����� S6����`\D��	�5��t�ت���z�T��^��OF0�ј�oV�A{fk��f
FV�" !��Ys�c�3����Sw=������Y���_����9�<�ۼ	�]����?rg�J�r���XD��2y�ܲO��Js~*E1����Ϸ ��L.G[�P�l�h�ݦ1��d"��H���}[,�O�g���R��<�b���(�H�ه5�.`�X�S��7x,�s<��c�G�B�a�9��1��E�O|��m�$�9E���s0�eH�M�Yy��5��#�T��ɼ`���m=)[���Ȍ��\:�
n:�����*�`˰?�?V�qd�m�>�����`��b4��D�vvA�xX�~T�f�l�L�D�mv�V�c�@g�ڦ;��������0�$'e�?SM�>�~��,F��r3s.{�3Mל�Uz̮x�M�������;������H��u�=�q/~����� !�2X:�}Ba4�dN��մn(�J��;�gW_�<KS�2�Zp�r���Y����-�zB����n�Ѯ��ഇ�o(�����J嘁�H�e{E�M�۬8�xj4/l�,:��X��O����ܑ��A���5�
Ol⨎>�:�Ъֹ݁;k({b^��k�鑻�)?��]4¹4���E�ܵ����ݓ����C�� ,���n��ɺ)�>��|+�1�o9��4t������-�Bn��K5b۔!��t-�9j���!��~�Z,O��6�T�c�l���Iv��LԴ�Ք��"���k�s���b3�,7���~���P{aoql��@W��͋m�z̤a���ɕ��@F�������pdFCH�l�tgO<��`��a�y��zab�\GvF�{�]��sH5^J��t�[��^>71K���;H��D��b��]X��t��u��c���Vv�7�˧ݽS�ø+v��8�j3�x�����;�	����UV�`���������^��hfrJ=Is�:�S��++]��̻ض�×݊X�s� �5�$m���bgiY��e����h�oW>��,ЋAH�}���o�޺��[E�0 �g��`�q�<c��{8��y��e�|�2�,T)XU\���Pꋇ����Wbl��1��Mֹ�H��/�.�
v�����掇�'�)��)PJ �Л���/p�N�ͫ�7�*�Qm�f��������Y�4�{��ҥ2,�s����"���q������Z�Ц��|���#�E�~����ʹ�2��N�2G*eP�*�ʓ�q}5�M��(����n���^m;�>w��8{d-{��Ժn�wȼ2�|�jp��m_Gl�e{���
���\��9b��_����A�ƭD�����Uq�j��b�m�B^S�k���'\]�TXW�t��{�f���}j�=�x�LM����,w�!�=��'ք<�pchLc7ƅ�̜q\zV������Q�$.�:ԲL�����f+��:��pC>$��J�(/��ˏ�Y�h��]s����.�ǿq�9��K�x�Ε�кь���ݖ(�,Չ���w+�Ƀ��aS���sջ���ò��~�~��ʸ�}QCB!M����򞭻Zݛ��MA�},�6e��9u-]6`U��uJ��
ʴk�W>�h�u(�q*jM�1���%��4m��$j�O�#r%&͛O�>�ͱNP���c�hܕ����{���h!3��a3�Q�r�c�x~?���f�0l�\���n���wC����92$lkݞ�����q�ȇ��¢���:�sT���3���Y�"��5� L��}u��2�p=5�x���p�aP{.!2b��+ǣ���������z����V������+���k�"�)�P鋇�k�<Edښ��`�����X@h�zi��{��*�b��ڔ��veR�,+	N�͋h�-���k��[1]���U�a�<��p�mc�5È�:��d�0�D��P"�P����oٯ0��w�5��	����b�)3b��X���f!����4�)�Є����%w
+A���i�!�soh<��B*��E���<�{w���2!�D�I�_<��t�E��eP���v����L�s�2�d^ƨ�TT�6�s��*S߹��M�v���\���t�& 2ae�L�]C/D��fz��(wE�L,.�E��M�L��8噃kϝݢT��Pdu�nչ�a�0h[��2/z��I���z�yF'-~垒��3p���c��ԅ
��tzX'~�2��9���Ip̵�V0����"�M���kO�j�$�ZS^�6=�}y8ڞ���,����b�V����[�}Y��v�	F�$�s]4�9�>'P�X9����鳭ܦ�Y�]���p�|��}����(���)6���*�����4ƈ֑	�	��՜���Ra�Y>��ubS��Ӊ�<�!ȡo�x3�m-.����B<�a�����Bm
?��U���c�,��2v�Z���WK�:�:�'+�vB�`�^��{���D������X۸�-f�ԼK7���\w�w��Wb�y��~����p�ʁG�ho��ǈ�^}���+q�f2y�K�Zm��e�����5Hv�����c���@ۮ�Oh�nn���5z&}!��ڻ��s)]�M���DԢ�/�Vl���>�ս�����q4�:�-�#�P��\V�O8#2��s�QoK���-~����/V�wg�u��=�%���PB�).⠽�se)M>��N^���.���G ��!4�Ň���&=�/gӍ^ԕ3Q�A����У	��Jܬ��;'�Se�'h={6p��{gV0�P�[fE�EǦqS���ڊ�M���}M	��3>��L^ {x)m�0� �$��u�x�f=zޭ�fC4 �|�CDSw��n�$k)���#S�f�zS]\/j8S
��=o6�D��)�>�ɦ�V���cP�_MҺ[��]�5��6{P��Ѯ���较�K�ʦ+7p��jq����+�㸨=�s�{8�8����je(�`)t��ݜNk��t8/�U�N�9XU�6Z��򟪇���|>��0f��`�xxr�ǹ����~��N�j�q\�Y!0Q,�ThR~���s�:y��x�[� ���j��J���@���Ԅ�aע�O<xPҙ'�)�ʑL��Ml�ہ��.	S�.�"g��^j^~�M��o���,sc���Ϡ�z�f�󸑽J�|�&*�<�)Ia��R٨����A׽{(�w>��~\�Lk�c��0��|�e�^���[I��Z~Y�m���2�̈́;.�&�w��Ga|�-�yv%�w@~������^��j�7�����d����W[�b�UǢ��mx�e�J;��㸂����gad�.{w��@�p�O�/-uEy�B���~�]9�sՀ5�RS�Y���T�j����wf�v���9��A���'�㴲��(��}�L���]6M�id*LO���tv='�g��h?�C�n;x4ݳ�eI�
���u�2���L9mOR�ϓ��Ck:Rpm�M0�ɠvW��sW���hV�FG=���l��݊C�q��Y؎p�#����L�{�͠��3�Яq�.�;�>5m0y3���}t���q|���NJ��Hя.M.�aP=��䩉u��h�d[D9Pý.&�j�B��h4��@�:vs�9nw ���K^�;�t$��,��E�2_F��U����9���6�ofS�a�}]��N�,d��NcKc�P[�ʺhH�8�$�VW"o]E{�.s� $�%�14�gn��Qe6R�D6��f\V�34�λo4tZ�g��Vl9�����aӬ�4`c/�n�J��3�9���δ�R����2�"��J��.�u}�d��ei�t��%ݔ��a����5a��!�ۓ0��%��Ա�m�l����%��R�17��]ǲ;���c�s-�QZ�.�(�U�Qv¥��:]��>�p*������iw�b�	׃*1�_M�JIj��.�̋�^����2�M��B:��p	�U�"����z�K*X���]%���Ѫ��A��2_n�M�G*t�f��~�*d�|f^Wfش��*�a<�����qM3+o���NU�TG�I�`�^��^&Ȕ�v��w-��,ú'���1��&�t����e�q;�ݢ�Uw-��`��*exjr4��V��s�y��"�̊Yp����Y[;�k�h����?.0�Tv)gd/����zum{:�p�緔���d�y��G���&�ʹ�;w)r걜��$��tf
j�*�V���q��*�;���(ƈD�BAf6J�虊�۷��r��(��в1��n����C���1D�с���Jj� )�|�˪��Ͱ��)�o���a��N�wՐs^4�����t���rw�L֜����ΐ������ct���pu8�����PTls������78c��,{5�����۹RY��Z��e6�Nb}G���'�S�9�K��
�l��y2�$���ٲ^�hߤ.U�HSk/hH�
����5[�;6���p`ǊtԂU��W:N�/"�w���tA��6���7�����Y�*wM�Ĵ�¡�vj����͢�h��\�q�k^�gt5�^sB�j i���u;��F�f��Ƭv��H�3���U�b×"U�[�I��:m�]LΘ]��_G���-�n޹3�*P\�}�ۥ������I�&��ju��v��m��� �����ߎf1rl����q#��k5ْ��_	Dʳ�F����g����7��}Q�{B��b�{&^lX�2mu�uq��f���=;Fv���0Ī�W]3��yaZ���C�K���'x��e����cOoo�Ve���Q�T}&�4BQ��nS��^ںX��|�+k�3X���_ ���y����Gk5�/�l�.F-x�ke�Tqٺ���+�qpN@�d��
��q������4�C����԰&��$�ݮV�ZGpfm�b����t�"O�(��q�˒ˁ".&�-D%&�l��d�c�O���g�y랸��E���t�Fڳ��I�NAɤ�Ϸ�����~�_����~�_�����4U%?��Hѱ��`[cGH3T�<>>=z�����~�����������Gm$ABUtM�r��RUE�QT��Ssh���F(���b�jb-�IZUQF�E�/9�jƵ���h�1� /\����E��TPQE1-�5SQr4ҚsUTy�Q-s>���jK�*�J*Fe��b�)�(�"��k>>nPV�*�ѩ-�Fڂ��""��劋���(F���<��4[V(��mA �I.Қ�&F��u��1-�c���qCB�e��F����M�n��t���qN�.y�[+�Ɯ}�'�8�HL�����}�uc�ժh�T��y�4z������85UC8����A\��p�~�P��-L������-��$I�C�Zsc6A�H��BE����%�v�Q�7=���dhbz���=sͼ��~���Ψ]���'���T�2��9)����v���z��2;�� rnjK$�����y6ʇ@�t��N�`��Xt����޴y������#�e���ǅ�ʀ+��)��� |�� KK�Y����shh���w_z�X3��5�����'ꔞ��T"����-q0���\��i�	��"Wx*��ۜf�;�R/=&�3)WV-�T���sy9�w�Iڽ�#���M�^��=��Nl�As[���bwGL�ڑ=�vN�6�R�1�J"c���a��Hv��] �D9�WK7�^�ޕI����Yd�����Ŝ�����Z�$�Ur&�20f0��5����W�C*-�$�f��F:�l�;�ל��*�΋�"�x	�iy@��=8^���,y�?\�c�o�U��M��3e��2��_*�*,*�.xnYr��A`2�
��y<;��ǐ�ƾ33��4E{��N�����jr3�[;�Fdʐ[�qս��w �u�=+���E^&��2�y���m-��z�ڇi���c�$2�lT_WWc�!rXHA����z5���'B��&�5�̬�X��b�,�W�k]+�-��%�L�g��ax���?*��y��������a�AE7
�v�� S$�Es�Oq[�Qa^Y��jº�	���sӇ����X�ܶV��T�P1��@q�����S��B�6���^J	{k
��N^�KU>�4�����g�;!on�aHG����p؟!ٕ�]sݭ��K.��l�ղkh�^i���.�]�����s/�i���3�C3��t)�������$c�c���K���������,�zF���D[��_G<��� hlov���k��BHu�L�pE�Ɯ��qq�ax��y��K};�H�����3؁7�y��^'lF�@tA�����`P`&�3���Pu�N���^lkH��C�v9���HB�5��;n�̷���0f�E��n��M�S��:�[:��C-q`E��{P'�r���jp���� �^Y�%'\=F��/U�A��,����g�a0���g��h&�q��1^��d�fg����|�&K���<˻�᪶�5����݄&��{�C�]���0R����>��7 ��$J��|��i�,�U�z&_%�g�QG�fi�P������.�f�a��X��"�gJ��D��N�\��K��а������~�}=dg�}��!��.��=ϩ_X�f;*��i�'X�tWG�mCـ�@�"��sԂ�yY^}:��j��JC/bw	'5���3ho����w�f:�vh4�����zT.�d�={gO"���C�h�BA�Jxr�d�\�ʱY=:�8=�f� ���^�r�I� �u4�^ƨ�TT�P�|��� ����]��	��.��1,ӵ�O�F��;
�!�z�HS��N�;��e�6��i?ye�M�8噃k��M�FH�!c���qkl��`�����@�zޑ(�'q)k�K�����,J�0��+�5�N=4J�5 ����i�`�d+�>�����}mi�9�xN�vKj�(_&��c7��<��v��\��oM�`Y�r��:|ã�:��xlY�+�?�Ձ�0�B�i�2nb諓wѹƭ׊�UҰ+��HNj���(xs����M0��o2	#*kL��ޤ�f:Iީ�\�Πḳ_�2�O�ܗ�9P���ۤlg����5ft ��%�\ӒڭC]��&�C�M��a�zZw��o:�v�G�."���U��ғܹ�t�Jk��8�j���5���O���t�6���V0��rC���������,��`9^<b,4�eEa����;���3���:�j�I�t���{�����b�Z2�'����S��02n��ku�ٵ���\B5��u���}1V���.��8`�GtV��m��e��?|���A'�i��7;�u����������a�z��4͙4GY�{��g���t�ŔyA�oGv}���u3MoI`R�7�qo-2�!�U\6�V�M��ծ�x�L�({�0Hax~b�S�ؚ�O=�Ƒ�*f���m��>_B8f��g�� ��ά~���u�4��^͜OC����S���#΋�?�B�����#6���X�͵�ȹ�����H�l&b�dIz	t�
���~Z�/���f`�6"X]j��Ȫ��ʄ��֛Cud�����-`�!N+�K"���%&D�Q����ηѶ��vF�B{h���v�����#7��;���$Y�^���N]�9*�x����~��2��u���5'���4dΫ���<����[�N͐�WC0Y{%�oJ����b�sυ�ȗ�����D)�"u[��1;c�����	��86�o�(��K�zE�L���hv��WX�q�����s�9�n��a>���%�C���<�4����=}��{�y{aqD��WR���5����t���[��wv��v!�3��P�����bI��)25�S�d2�-��|��6[3r����J�����ה�Xywp���%q&�]��{���*���pmGP��+�r���}XH7"=�M��K]�J��S�R����ujh�&�b�C~�r���L�X�}����'tj��t8\s�|~ �@O����z����7�A+H�sS[P�5�v7�':8�J|�"|sU�NR �എ�!⫯s����7�>:�n�Ծ�H�5�jÙ,:�ƲǱ��P1����2R��e-�t��8�`�@p��b�!�z]��ޚYғ�l�i�&�@������$�i�LH��k�����5����;��xB9��`0�б��L�6C��v8ėbC�h�F<���P�twS�2��'�E��s�dK�C`�渘I��,"���O�x�í��՗�Gsn��:c9� ��@��� ƴ�9���f�\BL9�-�}��t%����^3�՛K�S�+! � �����!�$d5�g�֎���������^����I�2�C{���?F�qaAO}5Q7�!뽀�;C��&Ԕ�O\TK��]3u��כ���{�N�!T��vZ9�s����f	�[Q���fn�䳮���M\ļKhć @��"P��u�g\��:8�i�	liC�f^��؏cg�g���2[����ˬL�Va��bud�:�J���8���B���&5�\j�������������o`�y�S�Ɯ�Éԁ��]�[�,�d.R3��3qs2J���:�ǋ�cf�AQ5��}_�U_'����Ỉ�ݘ�;����-�B��P�YE�B�U�`�O��T���9�?�6z�j�+�k�"FN����s F2]pF�����C��W�N��fⲂE���t��S�H�J��>[=�Ie�����l'�};�3O��Vl��*���t���.�C?ce*���Қ�m�!���qt��!)�ȳ�U��,�2B��
�]�J�h�f�"^�����B����łc|���P�� ^�o*	�ӫ(��Z5PmX����6�n�ލ���R�e&�`�� ��b�
����]%�\v�����'�o~�F�~��w��c"Kɘ������P���U��֮k+����[��*L�n���'�M��� _�,��,׭�U��q�F7I�o�f�}����xH�8�`8*5�������?K�g��ܛ��x�!�v>�d�E�u�x�R��H�e򘌤�n挲��BҔ��Û�,_u�ۖV)���3�)u2�"�kz�eE�cw2�aWAR�5�� n�P�ˮ#0���g����g/��؛e�W�gp��̃>o7����L�q��'J+����m]7��7`V"GY�h���S^Z*���{u���ڼȼ���5Шm��{�5#..@Ċ����ݪi��3]�3]���m�}��9�\���P�`�������>]�PɈ��l���[c$kK���������=�=����2*������H��DKXw�P�-���6��*�aG]��hmq�@/�g���%*�U6Ul�٦xi�sf[���;\*�{�yV���S�%+c��&I��o���H�
�Ç�Г���m٠�(���'y�di4�<l���܏n�\3	K&�ma�[\�z�:m~8l��ս����S mli�� Q-u����T(��{�e��Ry������ʘ���p��J.�laѝ��K�x8���9�;���������zb1>��Ѣ�j���#����h��� ��v��g9���i
~����3�eF��̼d_%b�*�*�Ŗ���7�{��V'!'�xa��6%7lr�X��yd%��L�loJ�=g٥�<��x�9QK�UDV5�Л0���:U���  ~?y���f���P⻶�(��Vfϲ���Aq��Q�^�z�}����o��g+=Y^���j�t�8Oh;C�6�6 ��򳭕k��A��6��$p+�N��Ki������=���6$ss��f7w�Lu;T{4q��r��J�[s��iDH��=�Zu��M��b���O�iqiTS���^w��|ؒ�rw2��Fi&W95R��bgV�������gc@l2��-�쵂�.��OQ�ghI�f�4�Mv�53�ϛ�=�I��#�>͵7L�s��,���]c0�����|u�;�ڭn�OC��'�4�Pˎ'mi��4�h �3��Eӱ�M�}Os �#y�:���:}C�T9J4R�AOIɫ���YN/�|~�ث,e4i�b ��T�%"�O�H�\9%�𻊕�"���b�4����%��ϖ����}SfP9�+(�y87�eS�÷"�{���ɚv͈'9�4(M�/�>w�r��j�Vf�^&x��<�*��P �6���Q��u�$�:��
��u���y[�M���N^,�q��$��ܺ�T�������v͵),��L6f C����x\4�rT�-�S#h3�3�_S��'���@Q85M�4{zRVܸ��v����Ð�ٝg�^�����aƋb߄g�5k��L�MF^;=D]�n�Z��jNq^O��]{h������Z��7�D*��E�{�~�\{c���l��3�'^A��ג�c�a#-�<�l0@t�~���ĸ����g��0��d�4�*��R�ޚ4�ʨ���������:�%�D��xӃ��L�6���Ǩ1Ք��;:�[b�2!@N]�.Փ{�$u����7W���
��?%��.M�|4в��9r�_ָ�V�x���/^�W�*e���`^����T��kl}d0�:U�k];��������W��Io��K����S�g@���CS�"�Θ�iǨ���U��ݽ�{��I'��&"4�G,�^�247������c�CЩe[��� �cWC�V�mu��H�?������l��&���]|V�H`�(��	~���
!�^t�~E�n�v�p�_o.�A�����w6J�! ���_	�X�)$V.�2n�x��;R�����B�b�[ r��;���7�������/Nc�Dҫ�����;�JȐ���:����3ӏ��w�F�k��p��9ʽ�!r[A�4�5�ZOY�R�a��f�n�vY�Y��Rg:��(w�-+�s���2wo2<p�3���'�]�y�:F�,B��A�x��?��qԋ��@�Z��I�޼5v�!�S{M}�}S;{Դ��iy�g�ζ�[�$.}(.�Eg�Y��M���x��.~�)m��2�#'D˜�p�t�5@a|�n
����ub'}ݽ�hI�x��I�|Z\�K�q�K���;=,1��]4��Vj�8���7�OAs�x�V�*��V��h�d���;Xs���I�n駑MC?����;��fR��6z���^Y�f���P�{"�Mp��Ӽ�!���6}����S��J������ �3n(�w+��/�;���O$L�zi����y�r��zҽ��[.�������
V�)T�4��I��v8&��N���k2��,J�%�����:���cܺsԶiC�oU��a���P+�mlޮ��n��禋:XX�3�yǥ#��Z���Õ`o�tӹ&�"Z�l�L����ߐ´e?[~����w*i�ks�:f�C�������=
�P��m���֔�� Nd�/r鉛Zӝ��f��nJ���
�e���k�B���7[KRmnM�m�c��3����ph8<�3�W�k�8Oaa_X�S;�ooCm��e!
e�^hǲ�{��l�|���ӻ�BҺ�3._4[B��2h��RӘˇC��BM���١C��M����5΢����rX�^.�	��7Mj|�V������$��c.�u�P�6�=
��8�L��n�=r���`V��.������O|),��,q������m�����x�J.�-i��m����qa�a>�hG�}�|�M\��W]5a#�O��y��[�3�N� h��.��)U�_j�.j3�m�i��S��#��,�;�t9c1臃d��۾a1�Х�֒t:N��M��ɝ�%��M=���ov��*[&c� ��Wjytr������*dM����բ�**�}��TH�n����t.�����l�du�OWNx8���f��:?��kX�ZaX0�Nl�U YD�^��X�"���rx��O��r��
b׵P�@����[1w�D,�	�1�b�r�dLո�m���\�ɱ��ׯD��
X��7Kh��S�6se��L͊|/ZZ��9)����9\ʄR*���2F���`X�S������q��WP�qڅ�[@�c������m���FD��Q)l*�ai�A�¨����3�0�Y��L��uT�~��:O��Zx�O��N,�6�T+�ُ'.����yN�w#�����#��:�}����х$�]��L��A�.���̵��IB^&������P���[�V��{��q�#�|<�:
��:F�܏N�G�S�Л�uϗ:�:>;��Ff-Ʈ(H*�6�:��-�'�v�J����-/U����z�+��13N��p��NR�u���L̩�}Wɭ�pv��
�W�<��k��q�E�Uk����!�ܺɖ����W,�t����x�yx*wm��ۼ�Qʶ"�#U��#T#F9o�nCd���/W�𷚴y���t���mEG��5*�¸%�1��>��Z�ff��+%zG�}��)�K6��[�i�M��`]U�9�D�7h�˷9�}���.巖.*�:��*�vJ�1��͉x`C������x�<�4�4��Kp�?ϟR���$�*���J��ESh11D�UUTL�����������~�^�_�����~�jd��9�D�M�SDUtQ^Y��?O}<}>�O^�~�_������~�����ESD���Z�5TLQG�4EU��!sbj"��+lP@UU51METS��U͢*(H.8�$E$�E�5���s� ��"������(�����)����娯t��*
b(���4E�q3-�L5QUZ�E����3�,EPUDUI\�PQ͊�y<�Zh���j����f� ��(� �G*�	���� �����d�EDDz�0DU5E��UA10DMI�0�M͋ժ)*����*
g�|oD��+ynv�{���|7_3:J�x+!vA���\��	(�j�X��WS��=�w�U��u�X���lU01��o7�=�Mq�z9�~4`���������1A��YCp�"���+pI]��;b�&.@ލ�Q�a���Y�=]}���q)���������{9�R�
~�=���\����� j)���+��������y�[�����%u�q-����yI�Mr�_����3l�}���װDG�J<��cj�sC�8$Oa�Fȑ��p��K:w���}}{�/�|�)�a�D�p^�۹��+�@�Է{旝Zj�K��wl��i��74�F�8B�
ǟ��n%Y0��\�B�E�=Q����ݼ#;��B�;U 	�s�l��&��UnEv�i	�h�cu}��^]� �
|5B��R�B*���F�)�[ߤvQ���w*�T�"�a���Ŀd��9�v	#����$����)�sV�S��lI���J�啚TH�&�j�wK�.�C�>���N(S�n�;��VIb�i}�E�p�Im,]yYkn���lc�;��`���'%�z��sl:�}�)�W�f �&U�յ�8P=�0Tpe�sR.����{&��y��������.�?,����
+�@ݞJ��"�Bг���8v3wk�W|s�^��&�(8?��ɍ[{�v�h6�4��Q��
a��SR�6���Y�e���}�S[a�GO�,�?f*�	����GD��Ԣ��A×&v�_:�	;���<������o{��-��b��,�F�F��Z�'zww�|�E�䉩�Jpf/%>��7��q��)8�9|��lH@W-�����d7n��8��	r��s��XΙa�-��b���; V_�Gapr�j�FW�R4���ې���aǅnvƺg�e���%l���C��� T<O���H�l����D���5Ϗ�Un�ˢD���^\c!�!]�%Q���=��u�(���yӚ^�I��7;�� Nh�KE]w���V=ϪY�tG�O�F��ǒ�� 1�y�z|�6��;,2u��0��/���O�F�ƭR��xR�C��-����9����d/DcWev�ܽ�L�t�cf�C�[ͧ*���^�b:��6�_kR�"�V�nT���0+�����u-j��Y\W֣��n�����BQ��w����ֽ�z'o���GɎ6��R�(�g�q��Ed�����k	~Z���O'GC^�ŵ>���E�u�R�:@'pG�&��	�Lk��a�9���1SѠ�}"Ȍ��ۭ�t
��)J5�eV��y������Q��q�g�������T��ۧ=�����Ԏ���qT���)�f7K5���u	ي >\�}�O �y��T��&��T�W�T���׺��\�",�<��w.��Fc��t��I�О�v�;S+؈���xVv/9��nA2{�O��_'�T�7@an[ 9Ҫ�T�\V��Y�5KƘ�9B�H�_|m#4Wt�ǀ]�m�����g���	۶#���w�2@y&}�Fʮn���*B�ޓ(UY>�a!���vc�/�C�5��!(��"6��a�8� �V�G���u�+$]������%���.��s$��ʽ�;��:��1������2�B�r	���`:Q]��=�6�Q
���)�aV�O��y�gb)^��G6-���c�1�\�f�5�\;���}'u�a��gR"���pY���6�ާa�^o7�{M7Ou!�UA� �0��?b4 ,�ZrE�]LvU�n�J��O��v�����֩;��o�O��f�@�n�[B������n�غ�/���ɮ��s�n-ng�ɾ��{��J�ҡ~s#a���N�	&69�V�Q��_{+:Ϸ��}��'� �4�p��=9��E�CHwQ6"{5���%�:�77y�1��A;C�+"!.�Jq[�zz�{�a&�q�Y��N�5Y�z�b�r[C�� Rk�v�1����"����Wen^��H���Ma�\�S�s@F����+�{95vd��r�-my�%��^�?Q�֛�L��ezaC5o
ҘwN���_b3y�w �c�]�n��ȼoQIO�q�t�)�̑tB�X����-ER�߹!u'4��[�I��W�*R&[+_��Ng�q����6��٘%���ג*�G%���hpҰ*�Nټ���⯟i�Iyf0w	��d��{����0PvSt�߅��
�XV1����	���g%�w	s��mH�lu������s7������۟B���;�']��%/�|~#���{��5�:�B����%R�\lk�+K섘ua���Sv�GC�� ,S�Cy�]q�W_������t�%�>:]Z�~�M��cu�ݍ���\�~�^�l��; :���e1�ȳ�T��@,�3�en�kk�:9~��J�(a#-��!����WW�qH�4�96�J�����ӎ�C[O��5f0��V�r�H�MѾmO ��5@�
��Eat!���*��;�zv�{��/i����2p�cp-��.z(�g��/�fsZ�u�U( 
���ˌ��s�#�Oi�8:G4[,f�Wo2�1�F�D
��7O6N�5�/-�f�	D�<y���������٫1;ïO�6y����F��X� ^"GY�Fό�2�L;c:z����������F�P�zJ�K����xbEd�)��Z+:�e�`�{)4j��i<[W�D��p{�;��xYmj��"T�u��3I]�k�H2��-NaP-*���rx�p�9�G)��3Q���4��q��D�XRc��/-�g���cO_*÷�4-�S���xh*��s� ��M�v�f��������K�Uٮ���'���ז�F0pz��PJ��#��F�"�L%�v�9����g:�x�������)�^x��D��k�,���Ϣb��^e�Z���Z�u��	�E���!`�R��'EK]V���i����u�M�/=�M��)�5�_���s�RV��RI%w��W��🦗@��uȼ���ЯT ��h	�pR/��W��%+F�V9�\�hl���bi�_�"v���:��y��/pYQ�f��в���Uv��������u�k�r7�r).(���(� u�<»�'�6�0hu1�ݕڶ6���̧��W�F��3�	;��7�N�����p�����j���q��_"Aʜ�wW4�`͠�յ�VЄ�ubS�f.F�}��ҷ������O'0n���'Y��"3����:��݊��ޜ�^_����omz0�N�$ih��%�"E��Nt�b��]a�m`J�D��ހ;A�p���3V�jѱo���(}:��$�⢈�S��"��sd������xc�bAɜBj�)�Q���O2E��>��_SZ�Ҁ�'[]�)����SG_n��I	X�q��(ĐKK�L ��o
�M<�8�܆ae�����̈	�qX_'٨�=͕�z7�F��t�*$݅�f8;��*�8�g���	��e�o���ב o*r���nd��~��������j��D/��!]�*��;��4�s�5��e��ٝ�0}���$��P�-��<����9��j�b��/ �.�S����6�Tof�(�$3��M�Ii͵7L�En�7p7�.�.x�~~
�q*g�7^�yQRy��S���Ob�ٓsN[hs4��SէKt�oX�Q�%HƊBr�4�-�t	E�)JQ�P����_$N�Viͺ��5f���U����T��Å��ԍ����U<CL����j���&7"z5f8GOi��Pn��^�Hs�y�������/.ס��,�;�Ŭ�{�P��Ɓ�	<��{�c�{Xz��p�,��� �_�z��`��z8�C��O�!}pq��й��_��j�x��,���ٔ9c�X�Z�(a1mp�ÿ�S�s&d'x ]������v$Ɠ����
�T!<g%�rF:�u��zĻGT�\c��֘�tJ/�]�������;|jL����`��(M�<���Y*{������Ì�z�+�m�tc�DA�|q���8W-y�2Ww��F�]��j�L���29��݃0�sW�L�:n����9ἔ����N��L��b����ʋ���7X�P�A6���=�z�i��Pue{��l�E��A�ǉ�k~�w�o)�
}�`g�� B��:����9"�.j�����l�o���ޔ�n�GH;FGPc���>����:�ZJw���64Ʀ����&j��^e�OM���M�;ϧ���xI�w/���@�|��/��7����y{��D�1 i�O��4{NYnjs�	��ٹ����wm�<��9�'�)@���P����Ä���:R�$�o�h�=��%����N��ܿΐ5�<�x
���2b�.Kh��jN���~�������yeߓ�2�P	��h�c���G�pz*����?�b���.Tސ��2�mX��^��9�z\��N��cw�=Y}^u�u	^`B�B	dN0?�w��Ty]�� �*�|�Heg�t�d3C��E�f;�I�{rNP�0��nH�sqn��
\�:J��"s{����{�{����d>δ�/TK�Lゾ�,���]<�r�l,;��$qJs��G��&�������4�i� y9����Q�SfM��N�Y&�L���#��ҙс,D��Ot�)�{�"E�H^t��US�eh����c�h^�6z=��)Xn(����D�el�Ns.��U��'Z=���	� iz=1�֨8/�G\�K�q�K���`�MZO��{?.�1�J[�p����u��_Gs��\g��*�qtR�:
�m}�Ն�yG�)�}����2�N25y}���Ƣ ]1�Ȳ|r�Ĳ;�YΝ���x�-��}9�$u&�Kl�o��دL�3u;�,˞��p���dq����W�+�ˤoKv��g�s;igf~����*"m`z�o��g�<��qF�˦������4h�c��c��X���Im>ϬU�k��t�g�t�UJ3`R�W2-���pV�v�:[10�٭�a�4��^�:X��>R��]eV���k�9�9��g]D�Z&�R7��tȓ����YǄ�v�Q����Z	���_	Ari�n�^o7���9�W�)ub��b&�3�-�#�@��=���P�ǲ��k��S���$����V�f���{7�HD�<y���lq�dnm���M����a��ɴ�'���֕D��^7���͝����'�Y�������V���ܚE����=�� ��ܚ1�2�/�goB.�/\����e����X���*��32J1�fڸ�7�K8B�#��=�##���w)�~mM���Ηqó1o�I*��*�vI۹��3�qHi�峃;=�P��j%<�,÷xH�=#�#T.�ĥBUO�{,��h��8n\Cs=�f5�qь\�d��f�b�W
�/xϯ�%a��o�Fp��B"%�j�#��  �kp�f�������}�uC�[Bx(��)y�ivXEzآ���GF9����n�9�f�ư:���hm�� ���d�m[{�r�l���&�ʷ���O�ng���y�aDF��o��yJ�/�W��㻍�s �*$�ݧ�*���z�q]l��
[�������p���тж��u�x]�ϕ�՘��`��Uȁ5�hg1�]�iF*"$z�<�H��^�uBb6xl|�=����J�9�^��7������,LϏm�[Lk����ss��\[���ٴ�}����l��6�u�Ҩi6m�-���	�b�BQ�5L�[J��`��q�z鷉��m�S����ބ��5X���\܇�p޹	�N�Q��#�cہȩ���±<�Y=� [�GJ��H䠯1bۨ���Tx,V��������p�����A��cO��y|��ii���m�-�ł��lc3vR�d��dn��̔��7dh�2�!�k��`ֽ��05X9�ᖠ��=�u̹}{ym�.Itd�{���1d=��bT�\�ҫ��C�j���� �h�V����g�w�K�ř�]��/��ʊ��,g����@J)g�Gĉ�M�dV��sm�rdV��f��t���N��d�1KXǀ���C�x��⡜�L[
�։{{��E�ԅ���	�'}gk�e�V�-�8��yhh���v�c�\�P�o%�=�x��xh4�J��%���n���Ϭl��	�#h�^�z����T)k���W;6�r�%]��F,S��Jy��T���A��p�Q���
���)�u�����.5E�f���֋0Y�U���e`�7�.d,N����ԇ�V5�ܰ���BU�j�߱TO��	�:d�r�v���5�.�˨⋵Ϟ.C�?ȍ��I�
���3���m�i=6_��Nͥ�X�{��50�9�TXF��Y-5��Q}[ ͨ�(6��i�2E��'�9�r�W����X��`�g
��L�nBg��b�"�v^�H�k�/�Ci ��[z��)؊�%l����4!N�<T��2��X�"���ي�X�F-S]b��e哼�R�̱9�+/b�V�p�D1@��@�P@���\����˩w����25N'+���ͩ,�����	��;������z�V@9�[d�)������
7�7��5a�ce�s�p�cv�31:�sz|.���w�]B�n^S�Y��bΠ�T��/�ٲ�VV�:N뾮KmA÷;�IΛ"�ù{}X��J:�h���j�cF�.ԥ6����1XBX�i��ϧg0Ԛj�Z�WF� �U�;6\���m�U���cN��kJ(֭f��=(�k��lWLI35g=)\�:�g'|��3�����u%sr�"�Vs�v�r-�J�}jO��AM�ml����_R#*ȸ��T��b��	�Z�6��Ġ7h�-z��]�f����l\$Wx3>�O'\@��at��&jp�O5o)�qE�
2vm�w�;X����`!�%_o���/X�z�4M�ļ�Cv���1����,�rbz�4��b�"	��0�4�t�1Z#�ϔ��PU�@?5j���G>"|Uҳm�{��s�yy������5��EE�gL�USh�p}�r�S3$珏���~���������������TMUQRU3�`����Z����jv7ۜ󚝰O�����}�~?������z�{�>�Fڊ�mm�b�(�(���$���bR�����"v�O�4W�"+N�|�bh�b�#AD���UTSETQc̙�����&���b婣����f��F�1UIE%L�5\����*J*9�ALC�CI2DPT�EM!�QÖ(f���
���O1��h)"��`������/1�f����CDRS$�ETQM>O�"��mT�IAM1̺&(� ����J(m�ULD�QIAD�ALQIE4Aԕ@LA1$AQ0L�x�,�DAL�%�UD1U>cAT1�f
�� ~��4�l0���[��}�|k�'ۃnt͕�r06�,�r��$�û,-��v�_��팖.�z�<�[����Vflu��A��E,3�{����ۼ����w�4�H-:H=k��եZ$�\_�������������<e2�h��ټ�픒�ɠR/*�|N�k��~����^�����RR@֦�E�7�@ ܌���mW���	o���N�.v��w�ْ4�٫���l�{��h�la5�bq�~��T��Cv+�iS�O�sf�x��4��Ovl�#�4�	��N>ّ\VɽG��<*-�0{?}��u�
����v�6եZ+d�mf�Gt-`�c�
���)�knu���.&�o*�U6n�f�Y��^:*,m�n:]�kWC����b�
h��5��ݽ�[Q���K�[])ا9B�B
%�ݙ=�h[s�Bj�/���p��������7B�F�B@�@���Z<��ͥR�vXc����kz�����	פV@{����P���LB��Jߟ�	�TfYc��ɥ��;t3�O/�m��	%S-��s���կm�0RQt}r�GL�������QJ�T��ͅј�o>;2��׌���.�;���9U1:	8-]VI���G�d�YG��"f��M
{т%��u&U�Y�m
�z�7c��~��o}&�_I�>�+�8uP|�3¼k�����C��E)Uv�W}δu�ݘ<6�ȭ����9����ԈE^��C��~�����8�V�W��"�kv{���Q�՗.�i@7����/q}w[�'�o2&w8��Z���'����f=�m�B؇��ݼHZ�]�"����H�t�Y-RQ�W"}��J���\��x'�;���q��?��8��T��2#z�]q�f�k�6��w.Õ�!��]F��Q��M�w� �~��1�	w���Z&&�d���ʯo$�w���}��s�˝5V�x�=��-z����y��Kc�"�w��J��Ǩ1�6�K��
����^��n+@Ƀ�2v���y�����Zs8��\ٻƸӓ�����$Sy�'�t����C8���������N��ݩx3	%�5�J�w��,U�z�eZJ�������]e��Ŗ;^����7(O	���gHSW��� ��І�O�~~g@��޲mm���u��tlEV����N�t:��."�:�3���3����u��8�+����Z�ǔW�,�zT�?/7��s�KgN:i��/�i~���$�o��^0��(i�e=7�}����TS��16�x�/5��^Y�Ǆ���:��-WE�Rӕ3�6j�mR��ʹh0��P�M]P��	]�rTFÝv����:����}��m��6����`�⚪:}�`XM������C˛+�n�E�����[F �S�ݍ�HS
p�
�X�~�Z5��#f�S9ܵ�YûxG�xك�uU{�w7�^��:���$,q7/SW[/"�a��w5�M���|r�yҔ�:4
JLq��X7-��dH�71�3Z�yk��k5��i	z�p�/զ3a"9"����&[+EK�"*���\�؇G0���Ϣ5�֨Y|[�
��Ҹ޽�*\_�Lt�R����N��5OG���e���W���Tqtu*G/oPWS��ˎ�_:}�����&�;�<�[}҉�C�U*�������l��Q)�=2�m8�=�Փ�f4Z�Z�F�&�rA��%{p�Z�M<��{�=v�۫2ޥ��Xcp�e<<-��u@�eL�]�&��Kb
j=��s�3�&w�h��z�d��=.c.�]���v6Cv!�oTAO�,���c�Ě��h�=}&��o�.G�ҭ�{�t�y�P#@�w�vGbhe]��SA����¥�,lj�Q��r�G���WB�=M��������^��c9���k��Y�Ѡ�\����IPl�����ol�]F��ŝ����wuZ;������J6$�p�*�����>����7�v禮m�3��9�Ö?{U���g��eC��B*Ѡ3[b�q9�bQ0���6	�/VKe�"vٽ$��.dL��Jc�iLu]m���Dd�,Q.��nC���oE��&z�����?��0�y`P�A+w&�c���x��q�gM�j���ޚ�,�t���%�ה�\ә,�B=P("��uۅ�b9���aZ��7��Y��Ɉ�!ei�$��\!vw�̛�e�8��y������k�j?�;U�\˩��d[4�鮥���'{���oC�p�S$F;����LM�@�h�M��ϷE��1{7���J� z�U{����*3۹�\�}�3�Ō�JH��^r��kd1��bG���U07X�z����b�!��ae�}|���uaMڍ������g�L��C�f�M�j�1��.�'�˧��.�R�K�������Un���4��\�׺�떲'�+��2a(�Eo�)8c�ۓ��@j��߃�"v�/>ٟk�kz���:+k��G���\Z=�<�T6��m�x��ߔ8_�ױi������Ο2n�ԁ�ɍ[{�Z��ٹLfa�<�6vo9����h�
%q�Gr�:���+nˡU�C�l��o/Y��[MLq4��b9U��y� �� ��,���z�L�d	���0�x8?'���3����=���H���e��O�(tĤ���-���࿸ 8��
���޿Iܭ��W�l��;f����3��k���!����13�
��@�;�\Y��Oi��v,mZb�<��;��7g}&~���چ�մy���;�kJ�b1�q�0ڱ��/NWa��֣��<;�0����D!�j�)��+RjW������3{3�H�{/6�i<����EZuࡈ��n�����ל�K0[�yYl�TܼZ;�m��e�6�[���,82m��F�!I����]��M�~�|>��=	�;�a8D��Ɲh���S��3���+���#�F����͵ϫ+:�M]tO�J4�!>�Z*�k˛/���c����̸ˍ���Xbы�nj�н��HH�Cd�J�:��;n�ELpǧV�hoK��r$,���	`f��>g����4���Eٺki���X�We�i�ǫ ��|�F�xP�r ��.�n�5�*�)F3��'9ط,~����Grc��ʽT�=V��9��"��p�|�3��N���&��SS�eЫ��+��������ԍ/��!��˸NG6_M+8m�Nn�PH�%)+n\hk�˸�-��6� ��M���W6���������1X�y�µ�G��o>Hܕ~�����l&�g`^n@����Y�o�Z����=�@�l��|�Erדi���c�%{��YQ+�p�����׸G�*1Oݷn�ӫ����{�� G�%�bJ��k�Gڏ'�oE�)yM�3f�T��[Iᮩۋ%�T�Ok�ׅ�'�}&���]A���;,7���9��MDn��v�B�i�z��qdWpBdFh�~����{$su,��ު�<���W�K��bT����h�	O����eh=����s_LΨ�)S�y��F�y�FDm�X<�ǲ��
2����]�˃Vcs�χU^S�v�f�����?���*Y�繟���{���~sq��sp��ʮM�d�1�џu0:#ϣ��cB�"�[�S�wt������f��҆kl_Z��:F�i�O4zX߱���mP��k�MY����8 $^Ǟ��B���'x�H�8��Y>��Y3_D��N��Y��:��83}T��0�M]^^,Du�9*"�i�
[�֣cl����#�>��B���U:�r��Gy���%���HW��߹1޻�����Q�Y�i=t�������!\`~����VH��=�tӓ׹�:sk�����$�̚�U@��:i�ڠ�?ké��,0٥+q)3p����7�pԌ�5h37�[7��FV7MRu	�����:�GPS�S+m�Vw����P��̊B��9���lU$�W��ɋN��)H/_v�\����X5鄼d�ʨ5���j�Ox��p�c}W#��]��u>���Xi�p{����f����R�C��h���=� �u>�ʍNbmؽ5��e6�P׎��B�ލ�Hߛ�*��JD�l��G�����yݞ~��n�z%��t4d<x��#b�ʫ���%.���YJ��Ktc����)��WI���%��H�Eq�����t�g=� �F�ܷ�.7rd�;Γ�{��l��]��}[��?�v���k�����gV{�,�3J�e^�,e�p͆�8�]�̏X`���Rs�ͫ(j5���:��=ԮW@��k�gP#Gj���v�I�p:�5����^V�/�#A�M�_)���� �@�l�6�wB���Ngc���6ɠ\C`�ϕٲ������*�&x��Ͽ!�u��t��l�$}��R[��=��΁}a�QȬG����#����5RqP���3~��_롎c�4W-���C����V-�U���d�td{���1�Df��ې���ow��Ҳ�rn-��*��7n�g`TO�Uۣ	R��Z�,�d)I�ާ�VL����S���>�șu-��W�n=B�iڝ��1�>����:e���#f!
��f�6�Z�c-�[	�/���Ҩu��}�W'0���Hh]������_6b<�ILm]?��v��t��y|��9yOۖ�w����t�dN�MyK:;�K��'F��=ܠ�6=��ΖΆl����a�� ��q)e�u��Uڤ�o-O�i��z�_.J�1YF�=9���q����4LG��YE#&�����.��T���+���,�R�в��~�e�{3@7�.ܡ������AH��gT8�UT-�z^�7�z�E�\�i�h
�y�J�u�g�RK�L���W�j�y��t��I���w�ut���@Q�%u�
(��\[iޢ���w9����ӛ=I<o���)gn��Hb�NB��k������b���^�;v5�oD�d�[ë���b@ެUǺN��f��+�[�֞�k՗=οc!�|r�5ea����&�D�,=�&�a��0fmڙ��D.�ۭ�JH�.�?`B��Z��4��7�? �jxȅe�.,Ϊռa�҆VV����x���_���b��V�9��pm��u�Ƿ�h�k�mLN�B�a�-���ȫ�WX�~�Oz�#��b5��1���&���}黀>�y�}e���G���psdh�ٕ >��{y-�$ML#>���oK�w��u����#�<ϧ{�;�/@&jS�ˑ8h�~[!��_)�xe�?�ދ��2T��d�)x���ռ��҂0�e»��}z��:[���93Ҿ8�s�����Io�{u�T5a��t`F³Qn�x;R.+��r7/�qw=�q��PR#G0'K�y�g��g��Ю���?J8wb�i��;��+�FM��](�f���E��wM���mR��*
j��b��1֢���ubݪ�^,��!�hl�iPH�O�mS[k�oh�;��e�+��C����5��q;Ay �
Q��5��o����W�dN֤�d��dPa�TP��xB�V�pk�Vо�̘l�
�ˮΉ#I��g����SG���p��Њ�z�#���W,����l���
6--�n�v^R��F���+b��F��mqP��ъVf�c0�S,N�[o;����J���-�=�d�G���x>ڗ��ml�t�|�:�[�!p��yY�j�okN^����a����s�x��/8��Kـ��+��YWEZ\&�&���I��5f�6�ͬ�&���� �ϊ��S����H�k8y���Q�V��t7�Ht,�� �`��)�*���ڭ�MZ���3�-)m��j���AzT3"N�}uF��wx̖�Hd���c�9q+��\�%lpͱj�Oi��׭3:�6�t}����}�^Ma��6s.XQ��,��cv�@�67{�{�c����-���Su��cgN$��Z�l�sF��u:�ZYsR6���[f�#o01��]��3p�+`}��l76ޮ��T��6��s���5%B
���N��������!j�	�M�6���o��5�!r��m��au�1.�x3�)���G|OT����B���"Us�0*���p��'z{'�eҜ�́}w4B����5C�d`޸���k0��.+�l�����ީ%�M�7�#<�/��Y�c듑ض�d�e�Q�Œ���ı)ƺ��)bG}iá�N�t|i�z��L4��]N_'�SJ´l�������4����1�y�(��u�s��
�o��P�(�֑�-֎�;�3�"5�mP��J/r��[-}*�X��6~���Hi��z3��ˋ��T��;D���;ͱ*�4#��6���i9�+�$Dgd��t����=}X*k�[88�xn� ���KGa���!+�wW������JP{��\(���Ey(o,JԘ',Q
G� ���2�A��u}�F>K�C���ޓ���ۚ(ޢ�Pܩ>\:��I5�>\x���U/F��.��f�D�S�w�+;�3���ƏJ��[^�3��� ք�&����cL�/݊�3� �k���4��[m�h����b͆�G�@�M_#�
��M�{Z�̎��m�
�j�;.���Z�3�N�Z��V���[�$��+���v[�\����Mhx(m��8s;)#wwpS�*��6��5K���>k.7&B�v���4I.�����Uͮ�^���P	q27��q�h�y��'���	ﴨ� �N�'q�<�D8�AG��KX�=Wϑ��/��m]<�رJ�kn�kJ�w����,�������q�DD��q�sf4�Q���nk�(e���T6C/^�[�nr�s�v ���<nj�h��u9 �6��db������]���b؊�Z�ߖ(��\a=�6�fM*R�)�L�:;��I�-�X����r`�#/6��;����RT�$���-TL_#0DDESTEE0QS�d������#��"��(�g�_O�����~?�����?����E$}�4�TQL�T�TQD5ED�>?�������~?�������ED4=�TPR�=��U��U4qQU�Q256�����҅i1QMEA1��R�i����)yh�(j�6�QT1��D�450�S1DM���E!DQAAMsb�(�*�����@PNش�J
���Ji��֙�
<���RVؠ�r)
v1V6��@�"B�ՠ��(#m�%R�s�c���r�U$I�i��"���� �'6ib�[3�8se�<l@QI@Sr�ɣV#R�M,M<�M4�Sȭ<�\ڊ#��s^`�d����G�ר��Q�Ѧ%�X�e�l��h9h�f&�9���5IksՃ�y�\��msb� �ѫmPh��,�t�m�1�U�[bI.mQ�D�3Y�EN͍Z9瞻���������w"Bq�r��UɽBA��iͅ����������0�oiB���jC :ֽ�˒*��޲�yy�����t���������=�[H���}��]:�. �H=9G*b��Cs�����4z0t�V��h����7W���O.�{�����K=�Y��Y�y_�[kSG�I�+��h���Y��;%ugA�(%����7�9��L���w{�ÿ@�l��O_(�W-y6|�� WtM���x�����vO ��8�B��ۍ�͆��\v��{�0|$D����!A |ٗˇ&=Ö������;�eT%m3t�U�8 `��8(��ᔙ�X�w�r�V�X:���w�/Gr��.�1�$^��۾���؏3&��\��`OCwmoXo_�o'&��Pc��rn���h�<����FƆ�����^�=��Gi���kN��c��N�y��ji��n�5���w���*���?�@�^w֍昽�}<���!��Vv��HJ�A���ε��/Qx�,C�1{�	�F�E 7�{3v��;���A���5$��h�&,z�s�E7�Ͻ��R>��+d�:�8���b�mo2��Gy�0�wD�-ܛdt���ǥs�Y唪�����coz�,�߼�o�{E½qo��XQ	0kR��^&���B�Gv�"S�~����wv�Ce��{x@���N���`�PJ^�`���^��ў�	���9:�/���}:���|i�I�%�Ǫ�D��,��[�@�y���W���z���w9 �8�
�&�uU��:i�­��\�t�r�aT]�ѩ��O��Vh�V��$�g\�JA�5A�u=�uȵ�|�z��5!#���:b�8�ս���䊾yR�<��N�"�����v�VAm�R72��lV�T/�@n�U�����N6���{ͯO�:�7kvb��:�>;=!�8ipAX�d.�1�/���e�����q�nE��t�l���`./r����|�C�ި���cv�z#k��=7�{g�;�U��
���ʝ�W���S�Fo��8]`q\��~-���X���⎄�׽�^���ݼ�2\�d�@_5�V�y�*ұH4p�(�/{�H�л�v��[V`n
� ��1�˵�7F�3z,ǽ��db��q�Ea�V������H�{E���T�m�Lu�av�Vm�N��X��!�������[d�͇s����~j�s|��Th97>ӫ({�l���6z��}uQxt��kf��o��8�L��C�Qu��U����f��f��g�ٹY��o+Z�2���Z�bxu��$7�j�ǈ3>�"r��%mu���<[�@��g���ZoB��m�"pNH��C3���k>,�/p���ؼ�l���)d6[�d+�U8n�f�O��y��Ǘ�́yB�x�`-;���*����Hs��[V{W_Wuu�h�N�"}��^R��O��C�=�.�b�Eff��ܚ�Gr.H�����0�YgP2�Ԅ���s���t�	�}��������]���zEdy��U{& g���$�B��NݰkSFjd̑N����g/���ݼ���+�~pMϝ��˧�> j��8����Fd�W=�z/fu	ًl�#��צ��+(��2��4��E_��Ig���Ci��̫�&.vV>It�L�l�Z��,�(my;]���Q�j�?��TV�u�-��k!���X���w]]��BgVt7ho4���V�jݬ�i�[Ep� �X��C����l�(��+�5�������8��DM�wY1w=;I�WK��oGt�{"$�tW��~�&Jl���N�k ��:+hO�g�,�v���\&˪�����d�VS�*G<�Y�>�-�RO���i�s��eE�h�8z{ʊ���E��ؑ����+��f<��]gr�[ػCg��8�+5�t�o��;�O�5vr���W�	�6M�����]Len!�����DwT1�z���;⽙R\{o�y-����Fi�͇3���A���{��8'��u�~�^nF{�S�<2�:V ��@n�c'Go�>�!	͍���_��V��^f�m[��p�9�a�˅s�{qd[z�ܼHhٗ�N���FoL�P�-�;ѳ�+�upQg0����0Ys3	�`��b)����;�P�l�����qc�EG�h�K,U~��~�F���(<��H�g>ukhE\ʽ�Uь��n��(�#�k�W�r�3�L����א�ޫ��˗��r�.�j� ��\���ʬ��^^��ź��hO_��	>;ޑ���9�ת�mn�M�]�=x)}g�]���u�O�ZHޱY�no \��*)�Ǫ���V
�N���Y�� �$�yB���2h�SZF���(���ϗ��7�ڹ+����c�T@�n�XhD���=�RC��%Ť�֛�:t�<����cUa1��f�p�;���B��辕�k���7���-��;.GD���޳ƞ�Nk���ݻW4�GS[fg�����Ey��Y�w)��������wn��o]��^���	q��.
zd�\�U��V� �yA��hIm�$mKU7������m��p ���M����^(��>��N�ߠ|wc02��wf��GƐ_�M��zZ7�%a�q�y�'�Q�3��wd�kvGb��[�:�>�a�aC�f���:o��µ4�T�*\�>�Y�3��{���٘*�74�T�^����@�9�2XJy�og�����g�W=�)9:TP^�^��C�8��?�Uq�	�Ϳ0]�Ȉ�;+�͹;M9i�F��Y�ɳtcs��1�ޣ+B���`��#6��1�ɠF�=�4k%ST,e��|�ӆK9LQ�)̥�Pw���(��G:��͂�r<�#g#�Ba���e��v��˒�$�����ٺ�r�h��X���Խ�4e�4@(�[��+_f�b�X�D��wַ��Z ��l�S�`�`����g����;�}�ޣA��G�x�hd�����p]�����y���-�J2Ѐ�=Z�E�]LvW&���1�v��0:�!����Y�\�s,��P|^}��%B���K�����28����d������`H5���]�gUp���}P����Hy�h^t����BDcf�xv����.������S��B�>b��T�2:�v�v�:_�*(쮛��@���C�\㄁WF}��j���j�뉳�SU���'/��,���'�O��2�4�i���0l�t��f�dϠ����z{]wƹ�d�s�$dٓFuU����Mo��R]2Ӑ2s�4d�#�-�h:Bac�դMmymk���xF�RRc���� �s^ɍ��7Z�Ue�5��^ݰ��*E�$\�Ph��������c��J�<�wx��a;���t��s�J���X}��z�7�뤏J-��X��S;Ew�����+��zʎK�/*�����	��|z���n�I���adB "i��`�BƃaOyk���@.P�ylc�4�{�LRT��u8��&���re�
���FM�K���F�Z�ۨfouS�I��i�o��������$��h4Dl�ɤU:�����:C���*���%n�̺�3����]�QO=�~�U���3��f�%�P?�[�3�vb�0A�{zp�˶�]�͢k�Os�Qؼ����H�+�|w�HP����5�,������ħ\�q\�f�:�&y����˿�ʂ��4h![���,2�O��M��f��eL6u���A��I3�Xf�ҧ&�:���Gi84Ba�6z���Q�8]�1A�2�h��3�L8͇
�]w,�e�y��9׵�3��MU�1�5�w�����Wa��g|`ȳ���@J*��C���c�5ˏN�;�s}��$vDn	:��;jƋ0V�f���=��Q����rrڰ�t�3ss;33�i|���#�6��^_�_;�� Dy-I=F~!��6`f�n��f��՛{�ټHD�����:y5�,�E �6��κ*l�P;��岸�Ε7��]
̡9���[�t�>���Ճ�2�u�ѩ�h�q��0̋M�,'u�s_���*�t2�X08Vn�u+��QW���D�U�����k�E��B����Uo�k��.&�y��|${:�uΔ�����5�;��sFF/��˸�'�X��/$.�i�ԋ�s��?����7͓��,`S�; :�J�-IVKC�!U�$�B�B��K��[|��m�ȫ54�@�gu�d�lH��D��t���8d�B�a�Y�v9�n=��/b��^�MP|Y�;�����]�#2�
�D
�;Mc�o����b��;;k�H���=$�Døc����H��M�lpN���9��*����� �O76H�+}�*Vvϻo�1m(!��ꌼ��T�)��P�������	.�B�OP�����N�(�\_�����j��eT;��U���t��!��;ɪ��4�s���1K4��N�\f�o�����}�7H�`DX&���f�I�+��y-H����˦y��Ln��>�� �I�}�o!��6كq�%*�����]O�vGn������j��� ��J��7sib�=CN3O�`���W]�d��4�D�f-����*d[��ɹ,���F��_AW�$�|!��>3E�ҏ���m�MA*^�{�Qۢ��SYCf�zQx�K��`"^Ty���v%EU�^nN�u��z&ɽףVcs���)�K��!�sh�!�a�h@Ynϗ8MHm��]gƣ~��>{]Ƽ˧y���7�>����g��÷t'͉I�z�[aޞ�}c�oԷ:��?,�y*�O�a���h�`��/��y[q�|�	�' �r���M�KM��^������V���h/-GV�={6@��b�{�א�ܦ�@ȏ!¨��^�����	�'X�����Z���k�1�C�k��M�5��

��:a�6�(�u|7�Z�9�R�M�8;���n��;�'�mW�fHܫsVUA�X����c1u�	j���點��n�R��ԏ�+��-���u5l��@
Ymy͔[:&�_C�O]�٦��&),��1>nZk�WJ�QF�G\y��U��bw�)��l�Tݣ��m���^�D1���:���7�$9q#^zI�Ǭ��O;S��ծ�lFU94^����Ùa�WM�dGG�m�d�����[JŘ�	�Ͷ�u�NVQ�L]��YbK'C t����a�B�z��ngs/�jƛ�f�'%p���å�d���F�n{�z7����i��	�s<]IpP�ö@���Z�=�J�S���n�lktonf�ނD�2�B-��1]��oOU��rכ���n�1{�{o9�h����j*P�|{�C�[\3a����>��#d���
�z�DG��G�W��X��7���Ҁ��}��=f��V��34+�7�o�|p�e>��c�)�; ���۾��7��vMЮ�o`l!Ւ��v�,�ղܶ�&9�'h�Pcq��J��_�?�"b�~$�%���)߬�GqW�33D�.���ʆkm���ka�;��3�V��&���[!��rD8��v����@,�x�!摡x@3��;�W��G-�Z���v���*���=�k�f�bc�v���j��6}�yH�As��grb�v;�4��C�jL�a��^ S��,��N�t��������(*��� DA{�נ�D�'�aÆ�
z�G����e �!�a@�U�U�!�d@!�a�dXaVP� !�a!�eXdBV �!�eVP!�eVV� !�`��a�a�eV@�@!�eXeVP�!�a�dB �!�aP!�e��P!�`<eL00�#���L20,220�0,#����# �"� � � �(�(� �(�����C C C� �a� !� !� !� !� !� !� =dr�2�0 2�2 2 2 2�0 2 9�x��� 4�  C" M0 2�2��f`@	� �A �Q � �U ��Db`ees�ņQ �& @�d`	�`a�edfffa��LL �*L�C
�$0��CL C"��� a�a�a �!�eXe^`p��C*�ʰ��0�aVV����n���8� (�(�*����v^������B���`��3d�׻��p���j<�N	2�}7W;x�:��+�t�O���((
�z@��+����Āaå9!|��d�� ���� ո�m�@�[ڗ��K���Î$�����
@� Ъ  �� P�  I ����� (� " � �P � �� !$ 
P � �� %� !� !$@	@ �% UV @URA�	U�@�  �	$�		@�%�` B%�	%�B�7�J�g
'�"��D@�1�f7�N�m8���ՠT �.��� AU�z�7�ZW�g�^V�:�J�%�~n`���,5�B
��!�ɿ���UEq@UEr:�@�|>�� E[3�MA
��� @�:�Cҫ�-�4� =�9X�2�,
P( ���G��lC�e6*���Й�^B��9��B�^X�'�;��TV��s��AU�-
��B��M���zP�H^����v�kx���%��UElKb!����(�P5�@�ܺ�S�V+���+���HeeEY��YX��Pܟ��
�2��֬&��&�����9�>�����
�%EID%R@��H�*���	T�R���EU$����Cf������$����ET����"�mQ���mj��mem	*4��d��d�� Q6M�&1���ؒ������i�U�PI���kE��V�[M	lԊ�UFj]�uJ+V�V6F��S6[�ٵ�Y����
��Kdh��l��DШ�MY#V!�M�E*Z�T�&Ś�UKm4hƳM�Q��6�`kU��cM����  6��m�vwu�gEn�۫nm�m&��Yh�;]7r٦�en�	�[e�nn�k�m+4�ݛ���٭�:]��r�E���֛����ַc��wZq��3��JRV�PmJ� ��@<�B����燢�
(P
r�
(P�B���xhy ��fۮ��ݺ�5rv�R���qvݵ��5��wviҶ�n�+�g]]�j�j��KV�]�9۲wv�H�j�F�Q[f+jV�j�XA� lOW���w[kv
ˮ��[T���%-v�;�v�MnۖݬS�[��J�v����v�����2vn����ٲ�S�ܵwv�tW6n�[wv�m�V�쥝m�BvٳMe�2�&֚�ͬ�G�L��b�ki�ݶݭ�5Kj]�9��v�u�l)�RY������pc:���.���5k��u�ͮ�j����gWU��v�Uݩ�]�l��LM+kj�! u�J몹˻XS�wv;N�VWN�����f�hꕥ�5�n����m����ƫ7c]j�[Uڝ��Jurm�]�Em�Ƥ�V�ZjhѦŕ��L�  �{FSj��݉\8���]j�����vثX�ۖ�[�MY�kY�Vwem��UZ�Ms4����t1��P��v��:�����őkU���m�  9�T�K�w;�������v�:���9��:�  ��� ����  봻�  v�  ���m�5��kf�%�P�5^  j��Y�p  ;%` p 
�ɸ  u�� r� ��� At�� 	ݜ  �v��Z����ilCk2Tc�  x  /A�  ^���i9�� �k�( �+  5[(�  �N���fL 4��`  a�#�m&��iZ5Yil�   gw�� ݎ� 7T� ���(;� ��� �]@ �kN@���  [�x)�	�*T� S�0���4d���ؚ��� �JR�  �~@�TR�h0�R!6�I  H@j�b)�RKk�@Sz��L�(F,,~�uؾ�\GR��|P���� �|>��{�?�@��
����"�ܠ��5 DVTS�������b���a%��P���#�@����T׮�P�nȈ+�s0����UaY{�3�*�ʷFV^�σN�
ð�*Me�%î��eRK�w5���v��P��Z�@�uh���nQ��u&��h�x
u�B�<` l��m�x��J�ؚE�/�o-9�\˹.�RB�<�+������i���#ue� 3d��;r�ʇp��RÓj�2 ÅE�gCz�PoK��3@�R�Qf��:����_ ��5���Aitq�iA�(藠�oŬ,ש˚�%�_�YJzE	�N��JQ��C��v�!�,T��-t�YP��@6��� #yVوMCT��km�R�#�tm"�,����[�kn,�[1��H���60Q{�xEOu`*T�v�<��KHa
: С�Z���/$]�݅�g(:̵�l�aC��>y	*�Cu��w����uZ鴬jI[gh�Q6���[���J�����dK��*j���թ����v��Z�U��س�C�*2�)HY�Sx�f�m��;����a퍨CO#��&�ю��ɱ^��ĩ@)\�B�|�i����{�vI%�!�\ c�L37��?�.�iR�ٺ�B�� �2]	v�ޡ0,�ͩ[�%棍�lPP1L%�h��Z���?+���SxQ����dKy�3R��=�����q���[�@�U��ĘlT�U���N;s[��髟*�Y�%G�}yCh4XJ���f*VBWR�ؙm��Dl�p(�B�ڬ�Yqk�r�����QQHt��6�e�T���V��ۺ,XZAI)��ŉ<���:*=�,KtI��vH�mj:���ιĳ��V�G�5Z�"�V�M��$�ݭ���Ԥ�@�I��������YmM�,`N
��)�t#�A=;[����j�a�!ect�h�&6��O횞���GE���Xsv�ն�IUo/>ZU�ϥ�X5��X�,x�+1ҹ���n��#iJ�$�z�ה�/B.]YG�yD�0hOFnmb�$���qCt�����nହu��bV䙮'/��l��N�f��s+u pk��M�hR���|�2�Z�ާx��wo룴�Q��b�Rqܘ@0�4����:8�dr�Vy�%�N��	F���zr������z�X�U�Z��"X����>}C��b��~��`��M��,�(�qV���"��*�w6�L��[t��҆�3*	����?�zU+�2C�p���J2�`%c�.�н�V��{���:�K�H�"��tNet�
b�m�M��K
8���D��2�J��1���;M�O/
��c�����jjي,�P��Kx�ҫn�ۍ/ 7/j�V�ATmcV�^,�1k��d@���ȉIn�;��FPɥ�3 ��c�ޚD$�.�ԫh�6&2(�Um��	���x�@ �ׇ���F�[̼�A�F�9nV��^��w3-eIqn�M[�E͙��&�%�.�Su	�F�Z#�Nf^[�^�`ʷ+�v��M�R���C��jIT�q	������A4��u�[Y�7{5�^$�"�u��d5���̈́����D�j���N[o�P��,qWǹ�Ţ�-Q�3q%�'�
/�w"ע�Q-��C3e�
�[����hI��ov��2�����Gj�R�b�!��uV�-TV�Z�U�y@?�+:\�XZV���Cc�5Q#(��o䶳@�*����)m
��ӂ�d��śI-t��s��-=���]�&mk	�!��*�V��e�$RtƔ�I^����N �LO�KsV05�;2a��ˡD�1��n;����Q:�2��\��������Z��G��E�w@�(�]�.���+:=X�Cv�v�]eF��$��f$:����b�KѰ@�� &afU؎�6�f��(�"J`4⛴���n�^3�@�-mB&сI5�ԭfc[%E��*/(-[�ٚr&�������w��OdQC��^��*9J���J{�\kkj����@r�c���ֹPzF�/^�[�mE5�QU��4I�3m�Uz�B�D��슁ݛ��C�6ZR�N��gH��fQYw�� [M��׈F@l�J�bz����F�RZ���Ɏ6Un�����#.��c5�Zy�%Aы3	�!�%�C&ܫ��l�Ԍ7�8t���T�1	O
y�Y���T��d�xң�#Z���h�����zy��y�͗����5"3^�����e��f�J�j�ÁTu� k��Kњ�d��H4ږHcd�>�j�@F֭��2j����r=�r:fY��)��ݫu"h����"�&T�ҵE%Gr�b$�Y���էj'.�������@���u�땇E�������ט1�V'�^,(h�4�A�f�i���n�V�pQ���5�/3�+%�N����ݲhݴ��ವ�,��1nDA��taYAnSx�;�����m�;W��d��:R׺�"���Qbw�ʃed���ⴓNPʏ%�+L�-J܎���oe`]}���X
e�}d��X�M��#C�3K�0��AtZN^CA���!�A|�%}w�E��/��d��t����ݱ�5m���G2��@��4'�w�B�g"��kJ����H���z��Ɇ��&4�Gc�z��Sv��2˕����+�)훎�Y5�ĺ�MA�2ѧP
L�ziCYu�(���ZQ��Yz�fU��p[�V�F��$2�!���U�Z)<��8��XkE�ˤRx��o+B�����l���J�X3>ے��%��x�D���w��Xy��N*�����bEu�d��ر��QU�
n�"���Ǚ����YmT�ə�T���,�TX0Ճ,��U�ݠZGC���Y�A��)��{bW�U���L*aAm��j��R�-�HnmD�cfNYk�^�F�1�����HEoj�Q��0\q��T:�/bKîhaYRӤte�J�J6&ͺ��É@R4Q8e�Yr�ܭ�0�^m
n�,3�[j����;*�u�ֱ�a��Z����.���E��+mKmFE䥱<�K.nn���5��d�J]����k$�2���l$��"�La�t/��
�1��kâ�
��u�d���K��/):M=fVXi�a�f9�N���2�Ln�l5�v]�C5�y��
�*n=��ya*ND���C%XTu��.;e)����2V�i#r�	A��ӔW���H.�`WY7cB���kU�����2i� aGW��+5*ȦItHM%�F�vL97�jU���^�ܳx�YX����nmN��9:��9�y�� �4�e�+b�SS7j$r�l�Fl�I@�`u�Q���c҅��N^(��I��j ��n=QՂ��f��i�I�e��mՓqn!�r�|Z�J�P/`8+ �jR"P{h��p���M��74��x`�ص��w���ڍ�N�0#�� �ط��Kt�@�,2��F�3�6CGj�jX�a�6\L���cƒ�veG�0�/��d,_m��J��`�j�R�VS�ڂU̚��@��U�`��֚o1�`�lR�QڅE�P��W��Gy�F �M1�$լZ�EY>��si��U[�"V�d-�z4����ۥ�1$�-sf��	X	�K��P�m1jAUcV��ke�V��8�N�]M�N����ܱ�^Zt!,�17J�Jg^A�w][�pav��a�6�Um��mn���7�,fᔯY
A6�"�q�oJ[$v+
t�B���r��`�4�L9+���[l��ݽ�I��2f#���Uf�"c�ҩv(:�tp=���-���Ǥ5b�x^#A|Bx��h�0��6���j �S&�H�&qTZ[�c7p�M���%4TXŢi�yE 3!dm�������I�CvK��hۃsnM���W�%.V�b'@5"����T�ۭPaǉ;��νb8�d����wN�!��eC{*𧗺�UL-���ȅڇ5qf�L��4�/a`!���Cd�&�Hٗ�b���Yv����&�֛	�F��w����5�q+J��(JZ�"��j��H�v�R�j��k\`D��A�ڄTG�()j��
�U�Z_�H�NӇe��t��I��۸bB��,*�RAݵu��
�
fRoiY�N 		�J�؎,y�������KU(����w1;�f1vD�e��hV�a��ֹ�'�����څFqV��YQ����
��L&f��lT����)�<4n���V(�f�wʹNLՠ�{�lڒ$�b����&J��J�fB_��坠ј�47�OcwpbU��Gn|P��-v(�IG�Y�k3�Ʊ�(�b��`4�W�a�mFF��"u��BP`��HTӉ��<��J�śG
��[%�ff՛I͍�XԭJ���+Ǚ��I5���)����,1���R�`ԟ@QɲS��0Cx�(��;HF�1�+uvAi RcAi�&�� �f��yz�^��7���;���S$U�uw��!͕{_שe�μJ����q�5`ܽe��i
��0��S�˴����)�%]&��A=b�h���$���ivhc%[z�pk]��<
ZwE�Z� =�bV.�׵�X� q�����²*�7i��� XZj}@���<����]�+i�LL$˔�t�h�U�.E�*z��T�mܔ6�j�6�WVм�3`�y��:l
K^�̘�׆]���*ѹD���Z	{b��t�X�XF�X�8^`��D�b��:�pL��]f%N��Vt�&����gb���պƴ2ⷩG�@}�pꭻ�4Nv�+��I��T �]���nR���4��-��(�"�he�ي����â���,K3!4�N�:�t�(���s&�Ɏ�.�M�]�YM vKJT��I��T���Z����;��JC$v�5�u"kb�W���W[yKr��*�[{�6��Żj|P��u�� �����3A+)-fma���7wI��n*Gi�m���5�Ȅ�r)J�ƅ�X�Q4�V�]M�4X�&���i���Y�PX���
/4f���k�Tۆf��8է����Xh)���Yo0P�Ǎڣ[���0+ /MVV��	�]֛��������t.���RɱKumBD�i�7v��\�h�c�b�/�kx�dݻd^�m��O3�%�I�6X{�Z�2][�wk2���,L�&֋5������Z��TbN�1Jܫ�mb�!�[�
��x��(��8�ա�UL�K��n�i��(�N���<�H�3K���B�o����p��h�,��?&�@̫�,&��6f
��䴱+�S6����	e^$V�0ݵ噡l�&E�E��\R3���H�y[Q�n�KB�Ds�Kn��6((Ǻ��Z	U��ݘ�,A����ņX�)[xSx����թzU�ɖ^M��v�km�Y�f�(`T$�!G3N��#�ea���In�!7���	�m������9�h��T��K�+ ,lG,�t��n���.d�Ɋ�V�ۂV��M�1zI�R�U�EPM�� �B����M1M`^����H�ܻ���<6�K��ih������M����u�Ť����%��v͌j�ÆA��f��*�K�f��(Œkt�@�n�k冑�I�BK;�e|��z��u�إ2!�Y3]
I��P������Ӛn]GR�e�+b��N[�m�T��A��<v�N��P�tpYԢ�y{a��L���[� x���b�[Y��ͺ�r���Ɲ�#Vp���9F

�����w��F����]m����J�I [�֧�F�j��y.�X�҅��B4&��{�D�M�N��*��$��*Ui-����9H�2^n�t2ѣ�7@�̓"ɸ@�[�m�-����AE�hn���-��
�KWJ�3 �����aL8,j��21m�Y2��Ni�檮�
*�Z��w�6���3�zch�iJ{�E]<N��Y	�fhP&p�&�u�Mm=���l�,���{nk�+r�y��*ز�$e�t��Y�;wrn�i�c˼ۙV�f
�m�z�f��I��Wj}�C`عKE��)�p�pem�Ƅo$*��w{z�Q���e�F�<f��O\x[�
���j��B<�d�Q����΂U���'**�&;�Y#��EvG)���+�$hr��{�e���Ed��i�Y�R���u�	nQ�opY�"+tK�C,J*�.��#�P�&�+צ�{���*b� X.�|�C*`Y@BJ�.���8Y���`�qT�]:Uq��/�*�`�*Э�Lx6�5ctԏ�w�.Vax�^"�ɏ"آl��a�
baR�Yin���ۍ^b�	��� V�T*:�
"Ɍ��Y���M�	�c�kb�eӨ�&y����:Nrq5u`s�yyx���M�gS7kUEja��v�Nާ��6f���^�u5���8�f�k!�����T�e!�/iS�㼛�D�BZ���)�)%���R|��v֌��L9�iR�Yn���~x�u�q��r|�eb��6��;��%;q+���(�ٚ��R�/u������Jl����:���Q��ő�T��J�\���"�]d���b'J�kB��W���G�x���T����y[�^և�h�)�4;lhyj� �ח�Su�x\�bP�5�/(�06lf�	�*#y!�zl�*P{4+Җ!˩b�^"�T&����,����B�3k��YyZn�E3-o�-��̸�6���w��"�eX�W�̘l� j���h�^Sn
�[CN��m�	�H'�fC���pR�q<SO��V��XNjXԕ�r0o�z�w=�(�U�̀ z���&�sy��f��2���T.q�j�[נ�f�T�ݷ��|���*׋lmC;+{�[	�$7 ��RwS��*e�'@k����N��rAS��LR�'���6�P�Mt[��V6�z����ڵKV����ݧ���:=>p�i�%au2����Œ�t.�gwIѹ�P�t5sI$؃�O \Vw#�������;�Vm�jмU�11M
�8���VϞu�������D|�7��e�i� �����襎�Ƭ"l��Dl�w�Nm�Ε�piӎIkR��R����ʁ�ڴT����^N�ˁ�SVU�v�V\tQ�.�����]���6�n�wlJ�n�՘���&l�w]YИ8���uɽq�E�s�8^v�����l^�_7d�.8���u-Vl�i�H o*���lvow%(�9gɴ�*��U��/�g,��T"Q�����eۭcP��uxC�^�6g>����TWIc2��Yj�
w�R*ޢ�a	�wRܕpS�Nn���6U�y�z��"i\�V�zԀM�//f��I����䝸7�FH�E���Gj����TNw:Wk��7�.#A'��y�,J�ب�;Z8 �b�M$��)�ٖ�>H�IL��H��-��MuR��E(��=�p�Am��j*)���};"5�4��P{�.���:Ǒ�ߐ�E��畊�����g<��q�aCȨ��D<�ˌ�7�,�k��-b�O,]�wI
Q6.5�Q"nb�%�$;��A�'�;���]� ����n�
:��w�)JQ��������Ɏ�yqy�F�ДuMJFvo��CJ�o�?�Gʬ��ۄ�֋�����xh�=��'y�ov�q5�i�ـ��O��*�b����q��e���!a�%��̍�/[��悘�l�f}�͔{�i�3�����>���qn���׷jԸ�� 6(|��F���qY����X�8�IԒ�3����)��X� �v#-�b�z��8T�m��b�8M��.{��cYY��r.MW����N=u�NM`{�Xgt|����B���2f:=��l�yM,JHZ���®�]��4v2,�!`r��U��n��B��}�Gz]��]@�����˷�KwE��gP��1�� �LJ8\i����N�&�Eh\��o
{ٙ�0t��t���Mkz�w��Q�+��>��A�tlн�M,cG'N�.��@�:2[��r˨�'è�g��k��;j�\y�:��v8%K�����{j�f�W��ڕ	�n����kqWsT.5��)_���鲯M6��ڢ�A>�޾ɧ�� hrc�f]�_؜ݿ���݇��ٹ�Pɘ�ܜ�r�CG��:���ɚH�N�>;p�qu�1�vi��Y�C��p��c���(�=xpTx�w8������ռ�:;��$��K�V;5;xHف�'���m���pIWnʡ��ʹq��5�1*�C��D�����2�uF~�Br���dkV;�@<�1]�@��"�ʻ1u�S}q>�`����IxU���B��\�����[��Y�ӳv���x�Y8�U�5���NS��!����}z2V�E�}���t�A&���)��#S�z1����2+�WV�	��ft3�\h����r��N�`�HV#��Y����C�:�e��s�᎚|�
5q�rn�k6þ0Jnfk�K�y"tk��d����κ��)QUȶMwT��\����6\�@�.i��j�uP������o#����뺚�㑢�V
����T��R)Y�S|��r���Օ�k)G��]E|.grB>���V�eZq1���U���~۶c���ZJ�p�}GV��	PV�!C\�N�2uK\L�9P9����%!���m�)��R�����h���DY�)��aJ�m�0˒�S�O�v�bfN��mkkh9
믯��ތ�S�;����"qV��+J�ehdH8M�˦����GLW/X��ȜڹA��$���	�)c���XT���ʳ}���v	y�	kM:���+��(�k��µFAN�l���3o:�K��3vȋ!��c#��*��s]�T�+DQ�SK�p��:ejy��]�N����v�*䒬0�uƍ��;
鯳��fs�J��hB����Y3l⫭b�� 9��(:�uq�thN�mNjG�گlL��sv7i��MѧX�Mm� ��W��V�3��E��F�ӇH��gqj5��®4^_9�#�!/�����]]��Eٜ·/s��%O�v��'����Hf���QbL��"��E�YWyf	R����eJX�m�Z���/�upZ�A�0�Q�����G[��s/q$�]�P�o���VVlҺW<˦�=o�b۵��:��[�[��X�k�i����u�k ������X�I����u��ËEt[�m
���G@���l�|������u��'�O���R�Y��'H��n��fV7`��a�jwZ�<����iyn�#����)8�:;x��d���Fv�fHQך�=��Ws7LΡ�+��,�5�lw����w|H�����~֩cv�c�ԥ(2�����eA�^R]57q�_m=� ��e �v7��l)ᥠLnJVI'n�֖"�iug^�~r�@��C���ˎ0x6PI'Ш����\{q��m���q���2]n"u";�y��*"����%-h���-j����Pm���d�)�d�������j�yF���Mu�� Vgd�i����,������	+��ywC"�}ݏ�C8|;w�R!2.Vr=.G�6Vܼ�����j�L`��/.�l�G�/��e��n�	�B�%5�U3l���l���b�֪�n��[g��:��i]�t���`�5Y>]�0��Em�x�3q����nA s�,:��к�v^<�&����gs,X*ؽH�sh�5�6�������ҷ�
̻�Z�[�PS�j�j�PiO���d�\��7��`mm_Yˁ`�����xʲ�"��G1^jN�-�#{:2�oGm��+��z�;t�Bvv6�N����µ����Zk���\3H˓D7�T�AW����"��S�֖IV(��.ؖ	�J��pk���O����%^�����Mt�;�U�C��U��+-�ŝ�L�(��n��3rPF�Bw�W����z��a��r��u�0�n���Ø__#���$�Oմxih�%�\�{�N�W^;Y|�>i�2�
X7�^�Y�B���f[p)*��!{�q��t�=��E)���,WL�����e:�;A�]��J��`r�
��M3�fjﳅF-^<6������k���"\Dm6��e3�=���ٮwD
Z]M[���wYxq�J��VT&]�C.�6��GM�2[2���4;k�V�nܽ�i�I��TK�s�fੂ�lI8g�8�����*�L���7e��R���i^��;6�vQ����i�az�|^�����ڑ��i�搧^gN�SGWi�c��$�`p2셽����\���&���$���-���i�ky(Ԏ�Q�ܫ�w�V���-����C�:�qe��G
ݭ�[Ƙ�ι>�(�Q(-��Jv�Xp�ξ<��א\�|��҂�2 �E�v�oض�R�Cr�:(!�E���-`-�N��,GD�<K�&�l���C%�%i�����8�" ��c��q9���1���pMb�$'[�5x*F�/$��f�N����&�Ϋ6�qR���D����&Ds;��9[���ۦEGʖ��{ rf�16;R�m� �N�e8#�dv \���!�*�V�k�g�W��y|��V�����j`�l�L]����dE���V%c�eʔ�:t�Ejl�m����aie�=0��µaSd��Wdu0^�T��Ɣ�-ܽ5��=��LT��Ww.l ÆE��EP�w=������u6
S,)"6H˝'ݹ�j��	bW��9�|&�՝P5�-q�wQ�M�$�U�*k��Pf^��ͷzw��3E?�~�IWBW���Y�Q��v�1�x�Y�BӁj3nP[��r��G$���U����C�>ڟmG��Um8�`��0���؄�77����jn�E}W��(k0A�i'��V�1�k�9�c_��tmۿvx3(l����Xɏz�n�y��*��^=O�>�c�n	x�{Q�"+��с0Nܛ.�`��B�<�����6���u̪��!F�t~��o�٣����'�+�3�d�X��,V�d�8���.#W,U������y֓[]�C`ȯ.#����sC�5Q9iۉ��C۳.`1һ����z�9I�\���x��ع�&f�֯�
��2����O,��m�p�"�O6�A�B��QGZ[\^Щ�݂�7�q�B�8oi�B�����^�)C&���t[�@6��22���o�gI��NB������2����y���ԋnI��{c:��ȣ�n��i��4$���T�[W�.���|pfX���aZ����8�,�f,jS�J��3��Ϭ^���@ĭ'��j��=�̼h�BOPU�pn���>�؂��.��N�䜐���i�­μ��X�;ӂ��7\��I����J��}�t5����g�ֆ]ui
Q|j7;2��Cy�K���{V삘�Ur���1Xp1�ZEV��o,�z:�⧙dD����eky�b(�l��p	ݡ䣧��\�0G3��x��jZ!�#���2�%����R�p�������-����9=AW6q��Κr��tC4�w,��F+����bu�wn��u����gQ-i$ؑ�t�-���@�ܟZ�)W�m��3ȃ�,���|�*�t)U��/�B�P�Ʈ���;N��7�-��5�j
��u���A���J��r7��
���s�����[ kJ�=��r�S
���N�^]:�q�>M�����x<GIG���mE��o��Źj�v��䋧�&TҶ8wGKz�n��}��M&����iQ�ݸ����F��*��sz�tD�����)ѧ�e��(��U��=�ovy'����p�^����Έ����U�A�gY�g)��2s�T��c�"����ܙ�ˢ*�09�mY�T�`n���:�6��\.��`�ݐ�q��f p�D�'�ܓ9�SR��;��@J'&�V������Ie+��Etd����e�N���V٫��}g�ǹ��gq���dms��}e���>J�b
��MԻ���aK�U�c���Y�;��&J�J�j2�Qnê�t��B(�X����~���H�k��Y,N�c��δF���:]�m������V��r��H5�E�-EO{�f쇃��9���[E$C�q̓o��ʩΌ�ݫ�r|��#-�d�2�h'":(*�Y}��l�W��&5���6çssn�[��OeQ�ʀ褫l�I�=g+\�G,w������2�jI�f�G����zU�P���	��n�̀pj�M}A�}�h���1l�e��B"���bN��*)��)}X)^K�����WO���|s��h�յz�e�B�J�c/0$l�(�гQ9�,VuQj�����]nP�9b������H�����t�P�-q�ՏQ���k�$���'ws��(;	��\e�}��,��UZo��w�w�+Q��-�a�#�ݲ%��]����lz(�W�ef:�\�Gm_T�(�c�[�n�e[�|BY�z�ư@�C��Z	l�i���g�2ي])��g���^w�ןg.�G#>��u�-��BǅU�}|���~}۰���9��ڬ}�p�E��.3f�lSA�R���ҩFC1I���8˜����,�ur�X�uv0c�9�u.o��rwb�X��\�N �r� �Jͭ7�`�dܫ:�gܜ�"j�ŭc��j�S�����R�ubfڇ���u�}K1�n��)f�di������
��=�bs��)��nR�=݃ �
Y�k8�&�E��<̖��`�f���lTy�eL`��n����)m�!I�VLӇ�ˣz����8�r.�Q������k"�5%�51w٢�f� �١�T ���wQ�p'Z�-���M�f��6WL�H9�P�I\�{{Lg�Z=W�IW�v�2���Mi�`��4�����WQЂt�Ե�.Cr�M�7t�;Z���٤�ٍD���ԥY�$+�=ˊ Y�cY���_ǘȣ|��\-ڬI:خ9q�<H������3�<�\�.ýOa�c�3u=Cp\�+�5��0nd���CE��)�Z�u]�:L��}!�[�E.n���sE�"SyP;��:��+��i�,3Ժ`� �ػ���y�E�Qw|7]r>�[9�U�囯��7*ZӇ�˞�(��-\�6�HӅ��@�T:d{�n���lL�Y�����=G����x��+��}����;����Fu�Nr�n�S���;�(9��]cDw�-㜎�:z�.zW�tTdpҸ�ب88�\�����.ܑ�n����/�<�ݨ67Gh�5<��p��۔=�o�`M��|�^�#�j^��:�Gp�V۝��B���^�oMj�\:̽U�"�<��A��S���%AX�[��T��G���es�C�3��;��{�ݫL�Q&j�6�t�m�,�t�u���ќ�(�J��/��֎gMR��R��zvk,�vт�s���E��vYܒ��ܝ���».qH[{����S���iV�:��\����/w7Bi����[Ѧn2�[	�S�Ї]��0�"H]2���x�ɑ��	��f��Cs�;��lf��nvp+^�s�~�� ���rPU��@DW���ߥ�:;��~p�yo ��ٸ��f�g�8ցoL�'`Ɣ��f�x��SF��-<�
r�Tthrnt�&Gm泃�ԕ���{��Ǹ�%{s���Z��4L]i���ةjq��	p��р�L*�ős�h�����#�V����SOK�q®�у0�Nm�@$�	B;يpnf	�D�9��d�j)�8ϓ0 +I�R.���G�ֈn7Ug�g@0��w\�D��tְS��I���_>wԲ]Am���b:WN��J�
*�|�Dg�M�R��;=�
I�(i�#>*�֊b0Y5y��PI��SP�i8̡�Y����ӷb�PO���2�/��w��Q��]�F#�/S� &8�1�p�ԅ���K���9'qm�S-n��J�IIMPS7-v�`UwE�n�jK�݃��;K���h20��:ԃ���:�x�d���H��{��v�s���́�rX]2"��)l�%�GH���X���c	h�:��a I����=�I1c�[�f-͇�=}[���b7��M�IE�yP��GH��r�����A�f�� �i咭�:1W{�Y89��;s\��K�c��o�0�a��\`�V��Vf��m�d��u���VW _@vQ�o{T���!��C�Ή�s>�; ��oQ#��nѝʑ�f����b��}�\�l,B���9�r�-�n�eF��
|�$�WϾ�#Һs^��g	�
h�[zy_p�KPӫ*����B~cAI0�ԧX'��܂��xn���f�5"c8�Ա$O˴v�@V��o�S��ҕ.��`sb����!N�~��x�;����B(2� QZ]p *��@3�ୢfT�>[�i�Ǯ�1�V�}F`�'f�Eu�k;��;@o+��|�}{J딡��:�M�fp\yY��AT1��W;a�`mgmR\f4�cC������M�,���}q�B�bX�p��-�׳#�5+F�T�o+�{(fbƋ!8+��WS
�}����.�3j&��hT,�wt)����N.F�ck��+���.�o����S1�1�4(T�.I6R�Ogu��4>��a"q�0dʅ2�ۻ*�qn�VPw� �e�N����ST�u�K���T�\]n��6&jb�M�i��[W�|��2�J�|E��Nѯ�k颤���hu��]��j�˒�;S2\s��
�t��[�l&�%���r��g�j�J�=�F�:�1.��$��	An"h�w�~9 � cK˳�Af�*��S*��>�г�07oa��x���#�,m}][�eųWX����c���s)��jY,#͕dʗ���IV!����v7X�Ӊ��<�ҏM˃�t�N�+F`�{$�P�πvI�Nʩs��F�K=�8�>#r��tZYIu�EN��O��e��O���1��ݏ�*���O_%}w�*�@���x�Tjr5-/�WY����޾����Q�I3��S��+M��\yO㬫.aT��Bƭ4Y�a\��\����wݖ
.�!O%0O��|& ���Y�6�J����+�3�_lCW�-eF,��ֳ�y�v땻����I����R�����<���	�u_:ߥ����Mץ���ҽ�kR�گ:�D����ِF�7Hk�N��pF�+D�z��F�B$r�a����T��7�h)-OQW	Yn���m��K�LzRK��7�֚���ѷ��9���mjY���3bw���� TJu����^s牴�iYSm}�Nѵ�Ggp��E�Z�c.�INo�ea4��ƭ,��	��2,�8�-of�I;�|��z,jT��}Y{|`��@ s�l�ѐ4+f�b	������|sM�&�A�q�e�/e�D%�Zz���z���n��9VTM�J�Rܭ{�&x[�Y�;�V�B�����hpl|�a����N�)hY��@8of�`,�xp��lˋN�ju���ˣ�:P��aF�q�1�~)��w%�*�mQ`�u�4�kp����̾���l];��Κ	t`�Jre�ã���T��Ŭ�86���K���;���̑��Z(efφ�x0ElJ�̼	��Dc��%�x����5hJ�����ۆ�����' F����m�F�����,�}Z,'���^���4u�V"Q�SO�J��rV�-Z��1v��e�ޜ�Q�����W�cpm.Lu���ǲ��k�+tЧ��K����w,4�<��j�6�r0e_	�"�WANƞt�،�p4�����U��
����}u��XD�}���>�hn{�[BUY-,��K��4-)in��;�i��δ3v��rl�L�x^�������g`�17�%��a�ҡ�0L8%�\[�6�L���S� �J!Ωu�ж�]�g�ӷˉy��G:N���L*%j`ʼ�R����W,�ҹ�{K�� �ș֕oj��p��t;����* �,q�a]��!>���WMUҶU戩���ī�8^]��˟m���!]aN
{p�!
�m�ڄ�����zX��K �0i�gki���cN!�#!����z:*�ܷ���}�>tt��c^�����Mk@Jw
��ø±�L�v�K`[��Z��K�y`��Qn���8Z�ٛ%e�$�:�W�v
/%�r������ߢ4�����E�Y���o�L��V�PJ�Y� ��3�]��O��d�1�7�(���3Tk���)��mfBcTlT��P��u[�x��ogK���ݮ\�5��>�Qɔ7!#��cJ�oS�DT�n����eK�;m�b�*�3��6v�����g�7��w�os��w];�*s�I΀��d�%2%�\fB�T��;69�x�\��V����l遈���J�9̢z���a�#z�!x�����٫g��f�r��Է��J�4KB�Tb����-:=ݗ�.���:v�T>���U��t��`ʑ� f���������ףN�Hvn�ĳ�:�=ܲ���8�|եYű����^�%�ݚ4i5��XO�U]�gjijn},���1��&�+fZ*S�*b8C�%=wJ�j}څHnĻA&:��p 
{��'����ӌ9���[� ����C~<�T(�k}ZЛgi�����0L��Q�Sj���Ӵ���6զ좪��@��������n����l��̹�ka���8m���13!垕j<la�J����YU�y�l�pi����H��ꋢR!����W��9��n1V�m!mq^�hn���k'�2�g����jz��J�2�Z�%@r�H�<$�;�2�t��T��r���(�+ib�iu]��*+Ywv��%;�#E3o	�	T���PS�=�2޲����oq�xM�o�L�M&�]W��1R��ʙ�fWY���W�y�=�N��U���۷f�ڔ,�տB~j$�e�Fn�mVSW2��S7gw:k�N�
*X`��ۻv���oKۭ� �ZiV�ٝԊ,�1WC��}��t���鼂*���Z�S(�G~"�#ݼ��i۔ڨմ�B���t���7��x�UAND��]kԳJ��;@h���E/��F]=���N7�l�d��Et<Y�n�X.�Ie�X�v3ҧƅ��K/]�5�;	�ª�+.b��s"���:;�����r�� �h(&�\l�M�Iژ(���X�t�իkE���'2�6���pس7T� ��#�gϻ0�g��v�9g��N�Q���c�w�i%��i���z��,��W��)����aYR�JWP�˗�l�~':(n'r�����<��S�r�����O��w]>�Xj�"*.W���.Ӗ�Ҭ%�.Ƨ�*>&�^Վ��V���t��l|ð9���Z��')2�eNX��#�����&�Jq/n��(�Ig;��:*�9�5��blM�MQBfJ[���mr��E�a��U9�}�MK�h�^��p�{�Ծf�E���>
�l=w�����z���"�c�"���p6�f��P<��������^;j̘�H ����/0����崎տ��Wt5-���vKJ��,bھ-�l�f�αG}�c6��ϭ�r5��]9�ܦ���Է.M�O�H
����V�v:8gg�NU�s��uX���Z5�,6o:4�(>��P�.�B���cT$"���@"�7>V���Ŵt9s9���{y��y+ȩ8-ʬ�Z�0�"��{g�2'Z+xa���Ѭ�b8^*V�9 |�JدPc�Y�4�U�&��:R�ӈw",��ãSqia��Ƀ����t�f_�`��E71��ĭ�Cou����2���wn��dX)h\�`qFYkAcs������vMZ'V^�5ي�%$� �mV��Wz�_Am ϕ�"��5�H=d�{f@6%�Q�0F� J;�!;�';w8�⦮������#V��.�P>��~�h�cV֨����}��.9q�/�-�F��������u��LmŝC39RRwϩ�[�F9�U����P�Y��d[@�Ii�feS�!9IU��t�l�1�Y��y2���i
tC�TY.�*�9����=0�mM�xwvk�z�j��佑�C���H�UyVn����7��`���&��
΅��)j���r��Poo) ��XI���n���j}�1�OY����ѵ%�X�qc�U]�J���U.\�Y�;D��T��F�2��y���̋��i�t�M���p����,��x6J�h
b���Ф��*oܱV�GB�]�i���Wx,L��K�+(v6��Y��v�J��i.@���ۄ�֥�<�3OV�z��ҹ�����V�.�W���w�*���u���a/�Oi캅n�Y6è�ծ'� �m��˥� ɏ�t+���ٺ�S�*h���Df����[J�d�[�����«fn���7j��������K%[oW�zk�ѩ 폶_�ȫ'�P�Ky�*�i��P�YEc�bʎT�yG���T�+PL[N� i������j+��E�t+o]�A��+l�.���2mr߯+8�eit�������̹S7�e8zU���)�w�0�'��v�;�� ��,��vj�tҫ*��]΁����xv��9�rm��;1B
�*r�э��`U��:Ee݋����9�U�]|zQ��4kAeL<��Yϖ`e��<6�a�yNIH��k��i��v�i
j�Vl҆�{܊��*Ԕf���`I4]m�ؔl4����8�X2:�O�6����ɜܽ[V&V�T{�ȑK��ۥ26�I+7�m���s���T�e04�%��c��aA�HR�Vmf�N��5�
Z� ����-
\	�uмބ�����>[����/����s�� �nG&Q(��o�{oF��di��m�앱*k]�ۉ8;/xr<�Wh}�>G�w#ui�r[��ss�Y%T��H�)�p�^�w$����4�`p��@�/�efaz����KZ��`�c-�.��'-��X�Y����� ]�Q��±�=]�e��L�r׬�®�6U<�)���x3k�'8�~��y\$�p�W�<�
�Q�yM�{0;���Ȟ[��&5����I
�a͂���54;fD���w:��45����z�n�N��÷#�$q5mvPv�l�:Px�K�:��Gp�)Wpc(�[��F��Ŝ�;h��k^��*}Yڍ�y;��d;�6f1ڙGM���U�Ŋ��i��t��r틧����rܔy�=n��\���TB�pp�*����47�k-,�9O�E)�S�ޮ��[0�޺�ᯏh�:�Tڕ���S�ST�����xUj�v%��.WV�kO;Jm�w�Qc����v�VN�&*6��93K�3Q��8��u��P��ao>"�ow���ry�6�-m�jrhpaS^�b6�'`���ola(G�R$����s('�
��|�)�cC��qA��$�V�'P]����H�cz�yb%�c���[��q�Y(ɝ[��Eh����qTr��s�ib�0��X�V�=�gV��1�s�7�T���!8t�*��eַ�21ßG�ˎf�7�2|B��,��.�Fv���GΌ��#� T˫��s���7����zk9ٮ�N�40t�[�R�βfS�Թs��p�V��U��(��w83e_q؎\��7ɴv�8y������o(46^�Y[�0E�rF�*J5��t
Q�P�����\����4��F�ܬU}���nhBabX����0]�p1��U�KE���J�t����=�[O�P�q�"s�s��/~��c��lͭ�vC�T�i
ι(iW�ǩM�6�\�����5p���F��h���WvP�H٦���ʻ���aokƘ���P|]l���!F��9�$%�N%L��n����Gk)��-������j��@�g������L���Do2]���` ���{|{�R̊�*T�z��-��1��y�X8���d�'k�����Q0)�`��첑���U�ť�.�}���[��9MrA�e\y�Smо�k.�p=ʋL}��59��řO1qՋD��"Ŷ�Bj,,\�b�]
�5H;��Efe���C7��÷�J}`���)-�Ƨ�,88n�'Y�Us����n4AT2���(B� �V�;�����v��/,�g�З�J�<0�A2�gnNlY�&UJxz̽��2�<j�K������B��A���;pGFR��ǟ@t�܄�oqN��fȨ\���J���>�����Phnj���H,�%_e��a�;���G8������:�����m��o]vl�^k���"���D����.bώ?�`����/;86h�(�6��yJ�d�,`j�*5ZO>oTT��7�f�zi�&dV�p��CVⳖ��BVNf8s��]�dX�n�Θ�J�y���;�:�`�Oj\�Y)m�F�a�.�,��k��h��&'�_�%޾�0:To�^�ҭ�R�"9v�%#{ͮV.������R.T��r�ɳR6���TM�Jn4�oN�؃�E5+���R.7�`�t��x1ƫN�$[����	��fS���,�5V8�ޝ��u�1�sl�CBM4�����i٠^�і�Dz+=uWFqy��mi�7�a�F������1�L�M�mZ�0�s���e롴Ĳ�"�P=��n�
=� �z��|��2�׽��z�*�mY�j��6��&��� 7%��݌ʎ��ھ=���D�^�>���I9h%�i�
��Kj���3mso쮹Igm�&�b��Z�d��L�ш��߲�Ē�}��YoiuԼ������h(�H��l���=Y�e�T������:�_:��뺃Hf�`��Lf��ҊEuo����,��K�z�����:���M��L��"��lq�ڵ{x6EsV����R�ڠ�O6a\��v�Ͷ��U�:�n`�$��=�e��y�2�a��2���]G�^���_�
룷�[A���q����b����Jfc�Rfb�I�4TД-4�@���H�-)ETAJUQ�L@4�FJTMM��Й	��9E��4T��B�fQAE%%)ITY��ED��!�PQBPUfU#KB�!@D%QEIALQ4йeM�R�!HR5@��#BSQUQKFY)@S@ѐd�)��$Ee�B��ESM-#Td9 S�eM4D5�dQAH�HSIД� R�!H4D�@P�%e��D@AR�R����H-4�@UTJ�4P��P�M%IJҔ�!@Ҵ!IAI@U-AAEP!K% R�IJ�J1���.����?z���N� Ҩ�F4��_�wu��}��6(�/k9�j=�ɓ�+��vU^���R��eG�sW�J�Y�js]$�1�1	�������wf��j�p2,77#�7�ȉ��4I]R�b�,�m`WV�5�a�������=���݅�F��a�i���XvX�W��Bߗ�z���Υ5צH��w����C¯+���ZS(ׅhF/����n����KI�^���<n�����E��a��]�^b�Oz�\]<k!{I��F�V9D��BW�kL[�؇GC���b�a�ɳ�(�}q�g��1�uN�-L����U8�Y[�u��;ʟ���(���ֽޮU�§
f��	C��1z�A��O�D:����ن���Z>vB*��E���x�#S3�ŖN+U�	q�����d��Q��H�ʞ�G����>�ͯ>{�ֱ�ӝ�J��d��ݶ�J�	8]#�.���F������������{�:��ג���㤴�J�}��`q�^:�[3>+��Iv�\�]\~8hi=��p
I2�J�'�v��xMꥅƩ�>�?!��b=U�^ʋ�D�IBh�epۊ�������"�V��2jR��q�S.���+�D��2�+�S�n_ɫ��t�=�$�v�^��ޱ2�;T��A{�q�FN�&�ʣ�B��������s������A�z�ݕb�H`����w����2�b����o2D���>��{*���v�߮:��l��x�#��F��~�}��a����DՇ�4�N|=����=^�@L�Hd������F���a�J��t�x�'Ѧ~&��|\��%��v3��P‡s��i|��YB�zB9t��p���}�f$���W|1]�h�mS�tz��^�󸚃�����,�!R�~fU3�q�͟x:����� H������駞)��o]۳Ƭ��.�NJ���T{��`ә�o���Kfr�\9l�6'�7������S&���~f�z�cęلu3k�?��mm��rS~�����Ӏ�=�׭��t=��y�$��� �Kڠ5��gb�׹V�A,Z�z�B$QXjey�ݛx:�Y�G£-���ұ1c�}���W]�c�Ob���t��V�X��z�_*Н��3�V��]	��^:V��I}���
�Ҹ9�����Ļ��RXm&o�I�
I�Mw޷U�'2]e�}�梫 ��;�R0��;Eרz%f�,:ܪ[���Vo���{�}yCۃ���r�-Z�i+e6�ʞS�R����BbIV�6��뗋J�GX��Q�	��Uv�� ���xz���A���+e�@K����N��@�Λ�V��G;�ȡ���R��2��I��t]k�����r��-Z��n�/���&�����v|�'6]�[,��n�-��,<������ت��b^��׏��c�Լ�#5o�D��9L�ȇ����s�3-��+��h��&���%��4����/z���S����ν{7M!Ჾ��T�V G|n���m���H肌� �B`;�Is�r�Tx��|*����[*U��9N��9B�9P��{�U����ʱ�ytû��~�Q%��� wćGU{J֨�+�^�"��b{���_��,�*�l����U�^�{{��Ox�&��J
��\����!?h��_��Ƌ*��ɰkJ���{inl���OLK�N��ؕf�)[�D��|@#�_�9{w�H���f��s|ΉW����z������XD�͂�w�\����%�VN� �gDT����ӳ�t�R�8t�q���� c��kmѸNcD1p\�%���q!�Tp��o�v3��tB۫~.%b�����!��T{%a��UHl�1�]-���#QqQ/�I�(�*}���~���kگ�!�d�dPX��ru�ڷi�0,ڏ�9���#�t��v�|�fW<4-���P5a+F�F_C}���w8�Yڰac��=ڣJq���8	4�N�&f�"iKn��j���.���I�h跜�J�Q�y�-<��	|��u�=@�4�f��(�5�|ʍۿ���'wA��傕��M�:TI�WOk�ǳ�m�Z����}�+u`yP�>w�G�Yb��T�,r�xI��>��u*�j�������؃�,�Hz�ƅX�2��<�u	Y^j|���� �S� �Ǟ/`����m���Y�	��.Լ>�~"E�S���h�s]l�>?:#����"N�QSZ�{��O�!ζB�^������W<����s�>x��_U��C�-[��]���ɱ��x�T��xę���u�x�9XҜP�.D�+hw`�Έg-+����c��|u�h߁+	M,���q��_Շ���y���xE����B�[��N�a�;A�:e�֯@����yWʝ��M��ݯ0	�0�����t����ɜ�]|���}�>�^G�y>���1�kzހv����R¯��	b�H���0/A�/�ǹ����3ttߺ<~Gp�vwg<��ҟ1玀XmfԌn��IP	D�u`R��2�ͮ���[܋ͥY��_H&^S��f¤͞IY��MTH]/),ܺW��u��ƌ|�i�6�9˪^r��sއ]c~��kw�����S�}O����JL�Wj���u�m��2��v1�z�L�NbaFtq��cy�^˛�BΗO%�Z��ÉǬRPƋB��=D��o���^EX�(���y;���Q��4=��n���N�cQ���!��͝�)�f=�7���ۘ�S�fE���*�#M�.�m�yWeF�ڞ�ޫ6G�����W���¸S��V���ŵe��V�}
R��b�Ң�Ōy�t���ӑꠐ��i���-�Z�
�w�K��=�_{�j�/��1�����[�ut�ª�;�q�X���+>'(m�}n�˵��k�Է\+7}s�����^^X���fc�ZQC���#4=��N���Aa�;�ls��]�N�^X��8g"���uTw=���{�İ������!�²}�d�i�%s�^�Q��e_sQ��M�g�2�6�����6 �>���Z���<1q��k)���_eG��1�b��$6���w=tk���j�� �V�뭵��i�������<}U,W X]S�ܓ�p��������:~~�{3�%�� ��V�+p�uN'fQ|�bǂb�^�6Zw�N����u�a6�+v��"�V���)���B�G^��L��5 �4X��Q����؝j�8'�V�o+�ųh�F��0��A����޹Mu1�w����^��=�']���v��k>&�I���$�8'P�����Nr�t�d\T�t�3yp��c�6�ި#��˭ou�����%!_Y��,/j�%�&����<ܑ^R���UU�W�3������9�3Ս�їK�|��"�N�������o!QN�bP�L԰���ü��U������-SW�BQ�>&�Iˤ�
���iq�W�k�sW��O����SX`aЄ�k]�:�e�q��1�jd�)�6
* <J������٬5sk��̀�������}�uO�|Ώ�׎�9�F��~�D��!_¤����ݧ����������r��6���CU��z�gkޙ�|}�P���m��Җ�k�F]\���1\��LS}����:�ȃ�$0S��`�nbL�'K��޸���=��UWH�o���;������׀Nw���kWR*uz֋Q��w���hg��[���6���p�pJWҡR��>�i*��֩�|�w����ج;����}vo�t�����[9�vA���?{�bF���M܁���of<I��a�>\)�=�2�6�tG]�[dj4"u2wz�@���Ne�� ȣ�協���/3F�ܕ��:2�Q"r�E��p��r��,����fIlTιGS�1��*�����R=�v�s�J7+N��ج��k~ī�o�p=s�ƍ>c�X�����{	�֦ۆ�p�d��Sv��2aa��넓����ygU�5�A��bꂮᗾ6�x�3�ܱs�o�?[�3<2К���|���P�>곧�>r��h��b���V�t�߻v]����W����{��0�l���i
�ܯ1�֬(���|׶�@��uK�1�hzr�6��e�d��Y�����0�w��hIU���]�/�5��������k n�:g��^�p,N�<�{ݲ��<�Y�Lx+tx>K�����~o�����J��{��;����u��q�ɨ��xz:�?z��K�ϸ�^���^ + ���ǲ��RbS֜�kg^V��N�zܲ�־|�p�P�����yM�g����
+Ԋ�w.��O �J5���b�g+�K�:�1B|�3��\;�/OK���/��l���-߼�l���Q}�RR¦M�Fת�����+�@�Ň�^��c"�X8��y���x�1x���]a�U.0�_Y���2��\����_���<�����U��I+S�F�ʏ��X-�N!`�J�r%�FM�o��޵B�u6��`���V?�������g�����v���oo�%�E���*p��������ʆ�=7\�9&���x��;Cc٫%:Z�:�­��4r�Vh�k:�o���r2n8���M���x{�#��\�R�$#�Ҝ�X_�$B�-�_���ro,��u>��������!��9�6����
�RP�wJ:$'�#�ϴ/GW�m�V�Hu�p[fu����Tj�tS1��%?�� �"G��4fc\�N��s͞WhE�z�����X�a�K�y��;s���jN��G�
1z�'Ǐ��|+28\
b���_BW�_[a�K��ĥ��.1��'�'w�bq�I�^���P����K�5n�L�m�h��?��H5�NP���9����o*磞x��5^/]�����J���xͱ�2,@�+^�*a�
��a�X��L^ߢ4���@�S�ɸ�m�z7hlf����/��ک�h�殢r���-�����̞�u��;6�:��@���EߔW+�F�y�X��{~�W<��g�y=3�׭a�i��Z�(sM��_{���S��qOUm�4�鎪���`P�N(V����`�����S�a�f-�7G4z��A:��_��l������� ��6��o�.޺�x#b���+Y�_]����O�n�\k��z��*�;%�y�q�[*�Ya<g�Nꛮ��6�-���)�t* >#]�ٛ����^�q���[\l�>9��sOg���I�e���ϩ�]�G@�8%4�+!�n��_�P��N[:�t<��{���̚�����Vw��F��>h�Z�F��υt��
��~�\ d���ק�S8����+��w${�C�g��7㴢�IB���BQR'n�/!Qg��V�8-e��\���~��~^�y�#.!������3f�J�!���j�=��h�9�7k���:��\��#o��re?;��sH�$���#���;گ>=����O���U�|
ؙ�Ι�*{=�5+�����xCnbo)ݳ"�L�v����B�K�m_��r�QQD�wкsz�,+S��Wڶ�C�Ֆ}ŢU����0����E��y���P�G%���OP�K��]�Ы�p���>0�u���%�cŚ�˓�z;��y��xZ#	�,
����ա{l]G}�m��EF���Փ�7�Ht��(ŋS��XL��7,-"� ����'j�auF���ͳ�}��N�2>��`�v��zW�����ZD�����rsI��׏[�4�ܱ�u+�T�#�����%Os��,�W���"�J\F��e�8�j�@E���N�c�wc�c���a��`�2P�ihys��G���^��|T���>�����\�;�5Ρ�z�9+C>�֐�}'�9G�!�~4�������Ϭ��Ycb����Xw�g#�&��N�4��� c�gx�<~=�^b��ޭ���Md?=���`����F����(�ѬM_N��+`��_X5ɥ�����<t]�%V���-�s: \��c6�Sq��]J��r������^�
��B~�W���i����6wrq�\[��9��={[����R=�g���ʝ7x������`��Z���j�c��	Qޛ~�����h�S�à��Hr]?W��ᇣ�+��>�	8]R;��:Hy�� *+����2r�]�o�;�8�Kjz���
����W�{½���>�F\�V�(E�%�U	��bU�k��A�\�w��isr��ޮ�b��5I�g�k��������l9�2��6
5
+�y궟�PL<��o����m���mRg�M�Ơ�tx\k�i�uto�ڽB*��]A.���j���WC
.�����A���5�ނ�o���R���y,bs�H�������=����edč)Zzw((���v�T��Љ���Tͬ�f���X8gQ۾#j���jle�쵕sR��[vl�F,t�Q��~��T��n����zs7��K=��3�r1�r����w�4�k7��4h�&�;��;>/����w��T$]U��V_iV�C#v"�q'�2�a�~�bU/zREH7��z�V
¬Gt��,���
�9������`��k�^�	\;,�%�Ǝo��WX=;��e>ަs0We�)�˛���wc�����s5r'_;�bf�He�������[��ǀ/�s��B6���<�;��5ta0}�"p^�B���ܱ��9Qmq��ۺ�7qo]����ƚ4�N�`��ޫ��#�V�!��xM��6���M���:��I��f���W��]�xwG=��W���C [���y"Y���m�6��]�Q3V�\8練(��� ��,[���<�fS�&�N�NH��0'{n�n|�*ź�{��9l�<#���5�,A�TΛL�!]h�N���R�5�^��:,��h�����ĕp��hi�j���X/k�!�q2�+R��R�M��軈n�;T;lZ��9&�
�̱v��/4��rX[[���D��SHhR�Z�S����×���ݸ�ݠp�6�<��g.o~��ԯT��FOSz��&0e$���x�U�+�a���;3��t��{�Æ�N�Fb橆��d�t�{���J#����ݢ�E7oE�A�-�2j:��9�m;7{��l���)lcA�Zx�	��5ÇE�Mr�vY��\�aL
�������&��eś�8+J�/���_�{Љ�}�|ON�#ma[�]�ؗ�R�4�=�f�%�S��)˕�n�06�]�׶�ZI@�pP�Ii�◊�fX�y{�&V��ݡEHy�����֖�}���� ��Gw�S�4�'GPs���S��ۻ����/|���v�_1�I�\�����[uH�~ssC,��.��z_-�\�r����b.�}[�m��uP[AWr8�p՘�*�0����&����I�x�Eo;��=7_;ӃY ��©Lcٽ���)1�aIU�.��;�[���[Q���|���ffi��U7�Y���Qeu@�4�v�`��fwr�yp�����1%��N�%��>�e�C1���Ў��wWf�����Պ�Y��QJ�t�Gqi�q~T�'�K��8'���X
��\g��
�.���#5t�`�&6�S��_l�#Q�dNjpZ�w�I����uh=]�F�cIw�M����a�	s��S�}I���h�0��ܾ;n��7 ���F�"�!J/ę��W��g � /�ay�f��C6�Ns}sx������N��9U';+q��6�JKN�W�3��
�� P�C�A�f��$���}�k,�Sfk�´�:�9��r.��Y�緶���:�����R�%#AAT D%5JU% P%�+H�0�P)(2)���������KM-(�Hk0*��S�4�:�ʔZ��
�NER���G	(
j��h
�BeB:�$b��� QU4)ABR��k���)B�� ɪR������GR�jS"��h��B`B�ZJ
)�.KKAKJ��
QMP�Jd�y�w���߳�{���`�K��rr�G����DI�M훸#P��t--�1ٝ�q�쮩r�!�br�x^:����*"�n<juv���S�;�Y���BU�5A�}�3���`��7~�Q�J�{�.���A���?K�`��{��������r\��2:=}_|Ǉ�}�=W��wl���k%Z����pu{.�U�9Pe�]F�=���K��o�h<��!)�;5�k�S@m�T�=��ְ�.��d�|��N��z�C�X�G�j?A��j�� ��6�NT#f���l{�o/=����ɐr�����#r�^s9����?k]C�9.~̻y�C�;�W\�2u���[�%%厥�yF��a웩
M��
�PU`��5U%�.��pQS�)ְ���<�^���s�'P~������Cs�=�Oo9��`��;~����!��5�`��WR��9����L�#����hz��2'��w^b�5�o��K��}��^K�Fh�_�߹����k������-�jru.C���w�/��HZ�C�]C�3�|�-<��Rs������I��}��;��P����kEѸ5=y��1i���;>�A��^�������?|���U!G����������W]~���w�Td��� �%�?IF�|� =�#�{�=ˑ��>�����T�bjA���?o���	����{κ_�c�J|9��^�������@Y'�	W!���{i~��_�ܒ\=���?|��?�!�q�aG�F������jMG�?v��n�����A�K�vu�ᯣ����ִ��%�c��{��yNK���{����Nk{_�~�2u�}o5�d��3s���G���xh���F�7=K��ƿ}��Mԅ=����:���s��A���F�)�N��a���*�Gpj �|����j5{�2��d�ּ��r�����7�0'X����H�"#)�;�b�5������g%�7�϶�^�=�#�~�y=O�䝾g�o�.�U.�!�uj`�����C��XnGP��=�a�u'W ԇ:���<�_��X��/�	�ό�~�O�	�d
�?oHo����vk_lu}.�R��u<�_`��?y��*���p�X����y?����g���]ڟ��}�A�R�5Q�b�`��1G޿w�p�
��4���Lî��+�-�{R�//TM�.i`��S�*m��~���|Kxo��>���p�B�	`܁*��H�צ/9�u�:fʃ���4�s]v�mi�R������yN�__T���a��tޑ���kͮ3��,R�������6��>�^��]�	�����0L���:�{���7	]��0uji󘺄����sa��\�!ٮk'#�j=����ϴ����MG#���}p��f��.��Ht�5�C	��H�G�U}q����k#;�:>ԙ.O��b�C�1� ������G�ߝmC��}� Ԏ�ÿy����4�ra�{y�P{/���&��٫2Yg�����~�^��~��>��J>3�2��7�_�u�W�tk�r2L�y��˨uFG���Ƥ�׺��-g�������\��3\�/ӓܹ?��i����H��q4r���m;�����{j#�w��	��|�t�����;��ꃨԚ��P��
�����n�-9�r�=_��j�'߱u��^kOP��.ts��;������5G��Cл�W�В��@�}�k�=�Q��Z��~��:��2�]F�>��7����_i:�s����{����^��s0yjky�P���S�\�f`jy��}�o�kag���2%���+7��.�@X�D����P�s�lz�' Ծ�N���k��]xk��u>K�ó������������!�u�7�V��e�n]F�����)�rw�O;����)ҥ^P�c/��H�,}}��P��A�9�~�CS�N�៽�dj��t��v�?OPjC�f����28k���~�Q����u�d�s�w%�:�:9��ڗ�H��j��f4qw�:sUo|DE���>s#��\���4K���\��NA���:�b�O���{����d�g��y'S��%u�4rO��5u���@QA�}{�i����?ty��ߟys���~s�|����:�.�Q�O����O�� �%?��3{������=���%���'#q��Z���^i2A��}��BP��ϴ�G]`�}���?}P��\%G'%��̾�u�^��<���`��|{�	BV�q>��ܹ�!���Q�OٞF�)�=�����(���wy'�jN�{�o�}���tw�d��=�����p�#�Z.�9^#�d]wvH�؇{�{�Q�[ɧ�5^�룞����"t	�Չ��|��a_ں�P}�z[�|�Kɐ޾C}��i�x<v"��w������+QHa���d�(�&(*�jmu�9��[m��ep�&�H���d-�j`Tw��i�=�Sd�<}�T!��!�RNU����H� ��jꃨ�yk��_h��\�C���������:����Mɕ'G�����I�fk�'�}:����?GP���|�������ZwRyC��3c����]��;Ә����1�?{�����$���i���]C��ߴu��}��׏���P���w�'����!����u9=������_'Uִ����j���o�'�_�V�z\3�jd�U�v�o������#���Z��'ѩ5{���������`���u��O/�����~n�&O�b��;}���U�g�i:��5�au�r��s���j^ď��{zMF��	�jq�]��#��R}�n7R?��y����˷���f//cp~���s0yq���Е@m��ny��乬<�z��rMG�᮴����~�}�Q��T}s�6��^,�#Dz��дnt���G�jO ���}�����tkp�Ortf�?��?A�gXn]��!OG���%�`��N���\��o�))�r��i(�:��eOg>�Џ��"!�{:�����_�����2{���[�p{���s�<��s�5'gx��2���XЗ0~�Y��e�#'q�5�˩?ֺ�P}W1y�4uPd%������G��>�����7�P�UU�����{��/s�������r��v��wR?O�V������阞[�S�Խ1��&�Rj��J������5	s��N�!������ ���������h��Q���o˼��{�z�p�F{�.��������K���vy���229/�Wgߴ{/P��O�`uT�ޅ���u�!�3s��b���Ơ2y.fa�1C�#� ��/!C�뮮[��;�����_����'�䚍��#�Jw��L��~�Pk�7S�9{'�5ϴ&�!�#��>�����{z�A�x�]C����˚̐���PH�>�D���
�^���>���]�����0���JJr�5��jO�ʻ=ր��{��~�c׸&O�y�}��>���%����S��G��@n�������u	o���<#Ç�H��e����U��b;���G*YJֽ���u��o[9B>���
Y��m��-n�|-���#��C����i]�������`@R�O`1U-��|;��ݔD�����Y�w������f�L��Q͖D�Ԥ��n�Vv�_L��wO��~� ��g����s���:�\�S��A�r������:� 7�5����r�^F�~��+�C��_y�v�HP�={�w�?A��2<u����rj~�>�I}@}c��>�<!�<���p��r�:����}����%R�|}��9P����O�����c��%?s�0߸>A�J�a�\�pj|:��0�]T�z|�A�##�{O����ː�G�*��@� �5M���!�o��2����nռ����>?}�O�>C���}yֵ���.fy���ЕA�q55���Fc���<�$�n�}��%:�ɸ��jO�X�����qߘu	s!����﻾�7��_~����w�{�ܽ�r2~�϶�w�R��϶��>̀�kp�FK�����i�R�y���RRS�o�wѨԞ�ә����~�FG��9�E�n�s�c�`G�z2�8��|����oL`��=P�:������{!���>Į����=Ig�����ع�`�s��]p�]y�Ɇ��XdϲUr��O��Wx���D0�V��]�#�9�E����0]m����
<�׹W�}��5G�N�rdu燣��^b��Bw��gt��ƭİ�$�U��i�t�ve�,p
oMO��{~'A�z$�3)��3�9kp��9w��~l�yl��܀�G��#>7���<�Y9��u�����z]��IWu�� �}9Y����$?��7;��LF��{~��>}����XI�����H״����L;ትE�Έ{Gya/g3{�lΘCY��=���^o����|�[W����e�ʙ�&�cQ��ndW�Ej����N�ҳ��t֜��Z���5��,<�@�|�^(�\WGv����Ȝ�+jK��.e�XVk��Wo&�y� ��������|z��o�K���;^w�r��J�F_+
�v k�λ����;��Y�u��ʞix��*/N������!����o�p�&�{�6
4f�<��l�˽���ɳ䰐׊�W�ڤϝ��k����q��r5�ã��v��;�/_��ZGmܽ��r�E�t�`�ӾTL��䍤��YP�'z�g~�{���^z�X�?y������/]�S�W�/|�`�Yj�����1�5�
��v��hq��BI�	�'��rfdEa��[z��ݔL8XD�6� �u��d!���G�*uz��n9gZ���a]�>n2ҕ���G��j�ɤ�h>��_�'�9.j��Ψ�,������.t�0ط���=�-e�﩯x�͗��{\6�E/JdѴ����^�x������{S�we�nu*�V!�j��w9����O+���Q�]�&
U�_y�]Ad��CL�Bɼ�˓�/��*�N�C�Ɔ�aj�a�H`�}��Ο+݁��1s�V�y�{��c��%ֻ&�x��%6X�!]/,��/1Ǭ,�<��W&�#����q��Q�B��:�3�𽽩2�3��7�<�v�<o��QT��/��o5�s�]��׋��.|���� 9ϻ3�\��Z]�	Um����סޙY7:I�� �����꯾��!���xg���Mf�̭��Ϻ�!]�{Q0�Y�p�o�x�]�}D9�ʚ(�޾Q�)jҷ�s��J������ۍ	*�x��Uu�T}���(�:)w��	��i�xƿW�@���E�m:���9��jpF;�
=��b��'B�_{Rw�t���
:G����]��ۘ���ɗ\A,�u����<�Vd�J����h����I��,<��;	<�� �g<j��T��,�/Ჾv5K�`
Փ��)�����P�D���{fo��s��!b��"�^'Z+��Z-�~\��L'}����=^|.Ϯ�:>�v����*~`y�~�+{)�u_4.I2�8
m"|�k���GҺu�b|�xXJ��au�h:;�E���{MY�1��8�ƃ�Pݻ��\�h�:
��R_%�'�7b���3�?[Ha����zzE�iyw�p�z?i���K=���P�IJmb@���^=����	��<��9"5��f��S��f�$B��RU����)�Pz��](s�Ӌŕ�T�卺�+4Kǳ2.��yMd�-A�ʞΔ�`���Rp,�Go���ƻ�\z���'�;P�+����RP�f�L\S�t�6��@S���)���m����4l[��p]kv&z�c6qɐ�0Ϋ.��Uv���+F�M��������\��lή�1W��;����e�p3A��[n�f40�J#^�,�ݏ�d�2�u�w�����<1T�T1�kUx �xm�u����#��M���k=���FAP-�-[-[sW�v8xz�U%|������B�GcNgg��T��ܛ�u���N�1��jӽ��5ng3-c�H�6e��� ��s8��Y�!RPH|�=�uף��VXUk{�����v�Us�툇ffu׹����OyS�\hS�<M���u�[^���"#��\�Z��},��ǲ���/�ުb>j�'/�0>�����L����ݢ!�z���R�K�+��a��}O�>-o���Q���˫�^K�������ϟ�Z�/�6�9��X���w��߼��;d����O�䵛湏j�K���*�[ǁU�{�C`���k�OY��?S����I�U��V�����<>c�8��L{�<�j���TY�!N/<ے��ދ�����K��(�]gP�������U4�L�6|+��:A]^�K�_�m+�a�����i��5P�C�2�����V�;���'.��d^�n*�c5Q��~����r��&�[�^�iv�D\1��D�ͤe�Ä=�I.�2��ل_msP-�����Xz�aKUv�\��ck^u�:;i�Ҵ���#v�F�NI���>��3�`y������&���.���u�{��(�M%,*y�0Z����+���_b6-��h�����bt�MO�u���k��eǝ ��ͩ7w��U
@�B��*�:��9Î��{�TfՇ�SU���7M�T��2{_����:�f�S ��:��5ܫ�Kx�Ɩ����[����&F ЍX�헲��c�M�h���m�M�����߶�G��M�.��괎��Z��T��8.P��׌r��mǞ0�ޘ��k̷�dɔߌ��9�W����/�U\��2�.�P~	��.>�b�hU�w��J�1Mǵ(��ԙ�\�Λ�M��)���Ja����&��҉�/꭬魅_h�Zͷ�w�['��+|yl�>S�!������]�y��NX}|S��j�:��6�쫖��񹧎��j��(S���5T_���Ħ�9���������}���֔�<C&S:R7S��L&�i�[�������fns�Rgx��vey�3ާ�=��)l�W�O�Y~a]��P<�V=;�r�=�� �+�p�81�o��B����7��7�Y鯜��wXF���V����-�NGD�ȯ����ٲ�n+���L�/}�Blᒔft�bqR�\CZ����.�y{��=S<冄�+G���}_Wռ����zz]�T_�V�4�>ӵ�R�_i����Ϯ`v�h��]��ָG�d�2]o��1~>�*54�����vm�(A9��
����ϋ��87��|�����)y���-ϯ�۳�U�6�oD��kL�|Ot���k����wbZ���M_��p!�:z%v�Um�#Ȧ����m�:�g�z��[ꑗ�� `\�_��}N��g��������4|!@:^㻅�����a���:��'R�zV[0HH�����L��p��`[O��ܢE��k�
�+i�5c�cӬ�^~C��M���͜���"���u�������4�&�tʰW���fS;�_MAl��x�#��F����T:�e��c�ɍ�����b��[e�D�|��ߚ�E�;��:{�>g�]ʽ�M��{�Fzv��o�=�%�w�W*5���T�;�!B���?V�w�~������m�B��wQk����Fk��@#�ݰ�O�P�\6�+��t�����Y�B]���"az{q|(i�;�J�� ���D��}�!��vY�YtLf�B7������'�;�J��TwtN�2�9�@���h^�yH)֦l�]kӾ�	ى���Ex���{����Co�J�e�[Z�ů$�c��̜�,y[	UF$=�]�}��Gٹ����Eץx�tc�����Q��*�&�u��3L���0��56�~�Bf}Jז�p�+ &��S�����^�u8�Q��zm'����C��w�fw���x$&V��N��'�(�{�[�=2��^ƈ5�[g�J�'����mt(�.�/�3�`߫�:�X�I�i�ȕ�^����a�� l�.G�CL�=�M���!�z��*6|x9~j�{�M�q�+��{9o����"��>*͘V��	X�Ҭ$+�nW���Ef;����w�^��α��\��!ҢҼ����Ymo�m�����d*���/��V>�Yq�ܤ}=��~����o��! &��m:��g�,��;���
�h�Ѭ�@1���7Amk���붺�]w�7�>ت��V%�
�%�Mj������cY��U{g�p<�2f1!aC�I��#��d��>^�R��ӫ���<�x;fw��9W����	� �+/}��dO���c����� ����>��Z-�~\���0�_zx}>�W��UZ����]�����f�:��]���K���Rc��Ff���Q��1L���ڬ���;���s:�`}G�8��;�[$)����McK�u��p�7�t�V��pUw�ˑ�;���W��0�G]X0�j"���i���7�ָ��v�LxSS�r#������m��{��<rAoa�WN8�S[�\��������][�>�|��F���^Q�we�(����Ly���Q���z�I]Ǔ\鑣oql��g�h�x�\0r�ذa��Wn	RZǵ�uf"E��S�J��״+��)�e�Kj���#���xa������4�X��]>�z�sW=�T�u@�+	=��
�R7�M�Ԟ�۫�md#H]o�˔�=|q9��u+8�5��r���c�)�kqM�K�y!{�,�2ɍ���j��L�Im�Z�^���4��WZ&eť��۪��Zx'^��y�wӸ�*+���peA9��WFtJ�(�}�ϳM�q�]��A��Cy b�S\7�*����y]YGs��\������r�"��:s�'x�PQ�\b_e�U�oe���{�{&Q�0��)�s�ޫ�{�'b��,����Ucl��k+1��F����b��^��S������,�:�+�ϸ>˟kʼ˹��M�-����M;�����:4C�
�'.�&�����J���{�BRpd��Ǳ�VgP���(ԧi�wr�������4����SO�庅�5�ݎ$U�y|r�u*�
n�f��;n.������y���Ԯ�b�u�lL����U�>�=��9��{�V��ө��6�B�e��r�z6{�
^��r�{ãeb]8�bCd��u^
�He�0�]����)B39Kם�;��:�v^����i���TF��.���T�r���KFwn�AB�@ޟZ�:w7�����ȵe;Y�o=�i��0n��G�v&\��k0��%eMͶ2fԎ�K7z餩�8���Y!��{:<�5p6�9�Oh��U��o��%��}�
}L�#���;t�s��P�0������<��Q�t��n�FJ�25	�M����wU��y6�IY����S��.u[M���Im@H�tW���f���U1]ӵ�4����zkY��(wKV���|���OYo3:�W|��ʏS+5�L� [��ws
�r:2��Qwӵ��쵭vČԥXA��찦�Y���}~WwQ,�n����s��gr�2n�	}ź��Q�</t)�:���rs '{�|���L�A�A��,�?fn�4�}�E�鳰�D���SہU�ml�u�n�[����[ƙ�֋ul�'0N�����h��܎aU�B憪�����C9�˳fr��}��7�PS�d�@�F#N ^l��f`O�]n��}%�δf�Q*�}��tu�r����P�Pnۻ�й�ݐ��rwb%/hѦ��,��%Y�܏����Z�����
Z�(i"j��)�))�LCTT�4�PT�R�QAICM�M)IHR��J4�P�U EBe�RSIKBSIB+E*SQ�d�E,DC@̥@U�	MRQIT-%R4�R�	M%-,@��!@�BPД�Jd9UH�ER�JD)BPSKKB�#ABP5JP�4��B��T��!ER咀��nK�w�f�l�M�^�c�q�gm�ݭ��#�#�;9�+[�3�4��K���9�vd��-��<�|M����}���}��zz[�L�aE��=W�@Q�\�w�M|Si^��o,/g�&�fh�Y��4r�{|=�E���ُDc���4n����՟�:�P��+�ԟ���y�Ӹ�|�w���EW��Wq)�h������F�=���G��\I�z@~�T^{v:><4���C�Uex�'�)��~��t�lBD+��n��^j!L�׹�.��J,��ڬ	���������ZwyT��y�9�~�������|����v��C�Ո����2w8�#�*6_�*�����,xm�{����2=+�CF��̲���i�J����y.��5c�^�IXD���i^��PZ��.U�Ꮇd����IQ���u�א���V�Z�ݡa�-9`Z�#�XC�*"������=��9�^�aC�e���J��졧�E�S��x���1��yS�q�N�l;�Pok�5gpM��� ��z;���1�,<��}�����MF�b-T��c��R��9B��]��R5�a�Uk��F�ar�aƤ�c�t�Ps�|p@�eP��{��p�鲱�lN��"�粘;�e+L�;�*\���D��U�1�P�n<�3�;.*�t��\�V��t�Y?;*]n%����kҰ$��aC9�K걄�9�����}��_.�ՆK�x>�~�[��8�����%��/%���}=3���:��Ħ�^����mz³K��.|�t���s6#\ǵa<XUW�4�=]qۣ�P�}�9�K�Z/v�)�w����-LW��a��u#�gY߬c(I,G��W��j1��'Bd�z�ߴ!��+���øRr���'���~�`ƅ��Ed8�<��p຦���%�co���r�=F?o3iuި;�ڧ�C�p��; �Ͻ�>���Ӵ��H�3=0� me��[����ݾ=�L�}���f��?W�*~>�r��:a��Hd�����Y<� 3W�����7��qɩ��)Ǫ@���Uc�O�)>��^�U�o���u��Bד�=o��OX|�#������A�sԐCU�3�/L-4�kF�S��z	�.-�4�u�ݿw��Yw��D�Y��<P��D���H�1*�CW�τ�~�8��n��"Н�ܛ��S���&���\_�˕)ZW#�%[��X��ԬQ�V5�>�u�֎��޺F�f;[�;}'��;d/�|wY�ݾ����E3t��l��u=��:L��]��Ғ�[�%�I���vj	LJ���T����9�q:M�]�׽ʸ��C���Ҟg'*���33"ԑ�9��tdۙN�.���;��>��荼��`��Y�#Dj���J�>�����["���Zx��Y����H˴��	X�[~�w0�������Q����ͪ�7�� 1_',/Ќ���_��vY;�DE�p�O�����^���!��`��ն���v,�ذ�c�H'ۜ��g�n������ٛ�moW��H��Պ B������Q�O/�&�7S���J��C���)�v+�!���V]���U6�Tq��QqK>�>&����T-X�ճ�O�������<w�s �5��G���󏗢w�����~Έ`���&�Uh�i�Vo����*���]n�8O���"�����ޫ@������:����o��+޷�Vn5�}��}'s���z��t��$o3|fp�u.}�b˴����\7$W���q�����V�3�+���-�``�vLƏ{�י�R��<j�q&7M@����UP�9~/�?y�6a|�S�^���4��"j��;M�j��p��n�\T�?T��ӣD�U���T�_������y���ބ+�pI�nwy�`�c��yD���n�ڏb�,�pA�FQ��]��'��)P�c��ob�8���MՅű;i�o�7�,�`Q��aS����t�7)�?��/��ngz�l�z���)�2���%&�6u	Ԥ��=�`T��_�����շs�ڷ��V�a�K4�~:|J~�ڤ˧?N�l��׌��9Ñ���Mqy��yԭ�Z��_mԱ�҉�O>�Q>�P�������U�;��.�3�'��Tǵ���J}����|�ܱ�N�I���p�Q�/�-h��k�O��gևn������),��S8�J�ƶ�
I�@7(�P����u�\K��H��{O�H�o<c��I���s�l�:=�������P��SN��A~�i�0\#~Wp�u����
gjD�u>�|�x��/��}Tb��aϚ�8��5v��w�}�tč^�ɣp��5��j�n+"FU�~�T��l��=�RK�C�����p�M�.g�U<�c���}�&
�{�J���������BJ���Y��������CL#ڰ�%�C7�^MT�;9GCQgwq\7f�|�톖ƍ{�=��|�*͘V��f���]������<,Bhc9��l��*vm�NwI@�C���޺{�W^��鿳��[�	5x��EWYg���Pߨg�zg�t�ؖ����F=�4�74�����\f����#[�������e�V<jG⌠���.N����-��v]e�si��b��_q�����P�9^��yh:֩V�!�U<=�]�]����Ӧ�ѐq�o�M��)mE2�?Ͼ ַ�lU�a�5:��s�C M��#e�?%����	�l��X�]HX��۳GFֆ{���J���xN�^
��R�����$n2e�W�ɭR�{���p�Dc5�5�jf fƯ�}�]{�ۯp+�ŢM/���T��M/j���au|��(����9l�pNԱ�v�y���7�&�PW����Ѣ9Y$���Ab�:����?.W]j�W�~>�Sv@���u뵯$b�Ƹ,r�5p��k���!ع$�*��M�O��w����y�d�ՕD;�J���Aʖ<.5z�1�r<v�s�Cv��\�h}��@iI|�P��~�!j���}�2�����ll��Kް�
e����e���z���ҙ*t �� �y��.UW�� 
�@�'�����s7���DY��_���n��]xAS�Rv�*���R��:��(|2�s��$	G�2.��tr��eq߭1=A��z��{@\k�V���<�\����>�Eo�{��a��^:f���3w̏@=L�!�iV(fp���]VT��^������4[�R�52�j!�j��M����X4"�X���Z���g^�k�� ��-K=\mn�e�W�;#��M���c���.��a�2C�����kd�	Tm�a�z2�J��Nv���o���� ���}U�Ԕ�{�y��珐�X�]��m�y�0�m�����=���\�eϭW�+��S�Ff~��^��K����дXf��`Q�R�F�Z�9Vkw*��?:^WgX����#<lǾ���`����x`�����o§ݞc����,^�3�q�N�o�� ��Wc���]��͆	g ���1�=�-�em1 ;%�!��h�c5���g�(Y���U�#~��������אk�p���Gm���x�%Q1z��2�d�Cۄ�����R>S��y��_�]B���97*��A/��Iy��cگ�:auK��x�}���x�L�Sީ�5��6g��E�+��������P�^#G\��ʨ5M����fs
��xcU���Ǯ�z���e��P����,$u
?w�+_	M-�SͶ��t���!�7^�?"|#�[������8�c��@,N���.��Ҋ�i)*kڙ�.v�z��#�����ev�af����;u�%&n,���O��k��eǝ ���6�e�O�64}��Y3��u'�7n��	� /n�Z���B�Iaaq��!�{|i{������}Nw��F-%μ�{��,<�@M�7��|6<�� �/q�X�� ���㽈�AA���sc�:��)Ԗ������s��.�d݅��V�\��SNՉ�Vq�tna��������w]�}�\_��*��
�9���:��)D�7L<��p�w�����1jc^�8L�K�U�;X}zf�C�`�*�@S�J�:G|ЍX���T�{�hK9z/w�n���n�l%����#�e�ܹ��F$��4Ek��_#���|����W�NZ>MRrz��Z8 �Q�^�(z�۝���zN���*�Γҹ�*�@��:G�t�i��wШ[���#��9��ܧ^TBڟ�5�d�@r��行���U �걗��ym4�ŹP|y�=nj$K�t������h�Z��#]u'-��j���� 0�`x�Fhx;?}���If0S���r3�z��e�M�R��ּך�IC��V�09��Z~�}k�8V{���*zZ�������^or�Iw�+�xzᵟ{~þ�~�z��=Q�?̯1F�{ճÒ���L����^�ܸ��+����]i�/�<M[5�����)m/�k�kꄾ�M#x�����rڞ��uL��wi����8��4�*�*�^���8���|���&�ou;��eޟ$j>y�[����T�O���n<�(��/zì��d�ܼϡհ�Sq̏>�Ov)�f
jI56��Ņ֮Q���wV&\у2�d�E�l/��`�hhU�ڙ�����Wl�Z*R�sub��@�}~�*U^�cFt}��G�+��Ek�x��Zw���i�uM���0�C~���:o�,�����8!1�^ef�)h�+�f�8EYq���i�E�7$W���?-��5��~�8�ϢܶN0G���`�avN�m��YO�G�|!@:_��/Dit����j<�0�K�^�	V}gm?>>�Y$�w��"k�luҖ�ݨwS(�_NL5tP��<;�C�}L}����@L��SM{�m�h+���Mx@�d�M��`�+�w<o���ϼtX�cբ�Ws���Y�=�gw'��"�xߏ�םp��<^�O;TO�'$o䟝k*@�]<r��+=5͊���W����~/:��lig��+�W������h��\��O�4D�{�[���.��0�����_Z��kn �MZ��"b�4۬�^�])F��-?v��T����`��o.1�&��y۵�Z�]y�>�ᱹC�P����`�x	UH�	��_��N���\z��}�zˣ��}�ø�l��6V����ͩ����MMй��o�X^mٱ����an��`�����$�f-|�u��UXلT����^,Fl��X]�Gwz�M���vb���S���o��Ph�@~�F�~���[h@�g��v��݀�����{6ʈ���P�}U�|��Bw�x0m�}� �y\&hY��:kl���O	u���+����E��z�1�+s%�������b������j�\�����CL���iڇ��G���㾕~��]���\﹕f��v�*��+����Vl�+qƓ�
��7f�SU�>�ړF�1�^�7�(S;����h��u_��8맮c��͹����KN�3�6FW ��/J��*�J�8s�������
��'����3�~��x����]��tg��*c�1���Y^��2�G/s��OU�9P�L���1��p�K,��)���y�s�]$5ׅt��99㛫��Z����p;$�����������#S���K�`
�©ۧS�coۣݩ��µ}�і��V�0AEVI�/���סc^\�An:���Ͷ�+�N1%�>q���`#���w��}��dCQrIڨM�H���O!'�s��6W��z�?q�����M�F99ncA���?@�,����B�ӵr�õ�.h�3x1��o���+ˬ�X�Qfl�ˈ"*̮�K=vQh:WK��r̃2.�%'*Ed��-�s�3����5�+o��5��9�����ˌ��^J;�%��2��uɧa���pلڥd|4b�no,Fu�����Z/�}_|>5�wy��:x�2)���qα_����e]=9��h�m����5�*v<���RyNB����>q[���^�I��,�_Wڝ$|\�Cg���n����a��U�w����(�I���KΉ�>�dX�9i��ya�P��Ӟ���]Cً���N��5���k���Q=&{���C���E ��zo�<h�>/P�T偿Z>�/��[b���^���J�R�k�ޡY��R��M֞'X��0}5����T�E�5'��7zR��;���'wB�`9���M}�b&1�H>,��1�}x��?w�� ��-���w���6���f�<&����"�:��b�,^�54�A�͔$�=2�=T�_{�\C���5�{���J�Y�;��ac���kU1}]D�������2��hE�1j��w�l���lӢvuX��0��'���U)��^��x����|&k۔ȿ1M{��0�d^y\�c���}Y���N���ٹIp�T�Z^fĪk���ĸ�]P���R�֔��֪��Gǋ5�l�a�;�m(�2a�V��>Rih�M���=�Y�b���>��&'p����;��J�W����z�O_n�ǫ]<Dff3s�����m^�"F�:�o!N�%^���pB�dK�]3��!��J�W)�]g�BT^ke��mG�;�Ƞ�#�uz��:��n,:��˵��VS��R��{L�{O$��xM�i����)��v�a�pAU&`��f�r�.m��8d���`�����}{�9���Q�C�r�u��}�5Ku3i�l�8s���M�o��uv�`�w�i��P{â�כ-��
��8��6
*.��{u�/��w�\�����H�q�CN�q��7��e٧�b���1^3�*��7bL�j��ż�V�>�7���rs���R���4Mݚ�j�����ؒã�49d���o��}�sB3��tu�����p�.3^���K��bCR��҃Xv���KfgUĕܦ���]�u�,���p]ҳkG:\��YVdްIXv�uQ6���
ԡ"��𠂲Po{_�Be4wf�}0��vյۇ�Z2,��J�v��� �vz�*��nW?��c��W!��ֵ��DU�l��̏��;�N>r��,��[��d��6i8˧qm��IIj=W��%�>!�l��.��G�7�4��{�lt��<���A� �����w#-ŕ�x�btf�[J�y#[��k_m������T�o���m�/�/{2=��s�'�^�gG���9�7�2%���e�M�$�!�j����0�lok�"8���Ď��'@��o9J�tE�&�v�\�oh�T�77��ꕭ¯��Wr6�y�r���p�`7Rf�L��sT�K�F�T����]RA�`�y���=��������1����k����˰d�;������{u7ж��S5�P�.�/�n],���:��lC�D'�{�슙�ә�[5�����0�R���-���a�ڏw�cX�NU��+�?hM��v���a�!�v�!�P�X��L��́^͎�����*�����m�����7�;���0�S��)���u*�U��s]�\v{��
�wuo�qa�;����]H.�u8'>X;u�_��:f��WL�-~�A����·����B���ۘ_�0�u�@ҙ�x�az^��op9�6ZR�X�*��Bt�_
�2֜s�3f#��X�6�勲�"坅����x���N����
t���˶��$sz��X��%�٘
G�ո��׊���a�!����7��㎐?F�L+J��L�M�ξ��
TC!�b��>�˳�V2E�B���p���	�6�\.Cx \o�����w��A%��}R��e]]Nw�ʟ
�BP�4�́���Q����.G�v]脠s	�J9l�E^��r�S9� � '�H��%�j�5JD�aY&f9#M#T�b�.AAB�%	K���E@P(d �d9Vf#��d�VIH�%%"VC��R���% 1Y�F@dP�&f%M"4�6bd�A�4bd)@�%OȀ P)I��Qx3�\�osVV�r�K�&Ab^v�td����\�2���Vl;�Q�JʺAl�r��=�����=����W_��_W�O�9�
��mF�+�帞�m�Έgܴ�VG�l���/
u����ds9w�^w��[ǥ���N>��+�!�r��S��>T1�b=�� �	~�X;���D��HX�pj��Cnυt���W{w��c��=� /jw��UN���QCI)����Ĳ�0�~���QFR/n�%��~	K���c�΀X^l���s�X��y+��r^��c 	��#�є|Ck��f4�z`���mb�<_(��0\�tĔB�X�-���u�mV �"�G��TO��%�l�����B59�<��D	�u˪�$���۝n�X���)��x�+�<_4Ek��#B��8.P��׌��^�az����cWY�����x����b�*���s�I��r9U��m�t�#ԧ�}��{sObv�TU{�K���Cٟ��S�X�DE���^�NT!x��:���zI��ޕ�Q(C�V��X�C�����6���2	��B2��>��3.�{��3swO���`K�_^_���`���ƺ���b�!] 7�5Ln�����ح�����&5h��	�YZsU���������u�Q\A�,��Ө��f�t��p-�u�:G�˪�IZ���o{T���Wo	�LшfL��T�@���}E?���r����~~6�����.��PIC���ZDs�z�-t�q�Aɳ7^�g+J�Ĭ����.Ҟ�^��mY����͏���S�ϲg�*��	���C��A#�"�1�����!�b�Q!���V��]m���My-���=ia���X<�v��޽��>����ֻ~^��3�;6��;��C@�5b��S45��.��k��o�0�~�w���i���T��;��w:77�!�=Ҋ�:�
Z���L/������Y�R[����_���E?,�o¶Uy�k�|�m���M}�н�}i��v��)�O�����U}Ra鯰ÀQ�X��z4�x}����0�*����a]Yw�MyA�<y�݊v��+��]S$yД�_-@��L٫�ޝd2���~��#gُNJ�˱�Z��2J�����z�<���-(HgA�ZS���&}�_M{�th9p��(KV�;h�#����uB�J+��O2��'$m'�ZXvBlW�Z�i	eU���Q��Y)����0Q�>��w��F��d*ѹF0RSr��m�¨�ʻ�QnU�1���Xn��y��u�$k�q�u��Mh��ں�(ު����kweJ�Cw$GC�6��#n#�mC�^Tq�M�9��O��r�m{�舏�Y�8����^���t��Jj���P�'[��u�"Y�B48��(v���9M_�X���h���n-�s�2׭^��ؓ>�:m�L��(�P����`��p`�H���͏`0��4�S8�x}�\�&s)Ѹ�/NU����-B�-*�&�7Z�5� 7�of�!��'d��lE-/�#t�:�T{��x�9Y����i��쬹\���Si�0��!�s雇�]	��WgrPԕB'GT#A����nD>�\Ϭ���mt(��d2��xupu���[���I~*�!��7^�.�P�!�rզ�y/�pv�y,��y�=�%,Q:����а�R���f!�_,�xl��n�`������_����vm�d��� �����0x�V�_�,v�0�-+�������-��c�ոГW��$�y��8�-;����{����(i)8��GĚ�x,��׼�˞w�;���LM�w�B]mZ��}/�֍y���%�]��>m���h�L�
�e�Z�2�>~���}��O�+`]�u�)�Y�9 o&A��QW�����)��4��A�g�����HKw��]Դ�l�Miֶ��iVBrQ(�΃����ۃ��b����6W7ţX�fd=��f'����va	�U��[���.w�j��R2��(�Y�S��7�'�g���K?_�Z�p<$�G��X:SKڪl��|���2���q�ޮ��L�y�"'W5�8����55D�QXx�8�|�pik�G��EYԵ�I�o��x�nr�AwV����������mT<�5��p(B�v��h�D����ˠ_���[�^�-�렺ɬ��B̿�\hg�(��(qX�I��r�oy�MN-�Oz�yi�7U�X�H@��'�%ܧ���vyا��q�*��ڝh�o�z��(Kg��8l1��S�{2���"O!��K�9{w�DF�����E ^�#�Z���xo�%�#,���;���ƕ�?�ׄ$�6I���B�b�0�f�2�_�<��ء��y٪�}�n�E+�1��i>��q!��Q��U����a��W�xm�n.���lާ��ɱ�Y�?N{�&L4��FṈ�h�������ڳx=۶�EK^�L��=���y;��V�!'SK��6���Of|�E�����~~'ٽ�K\��k��R���7�Gwu}t�
�D��5��v%ZUl����������H�7��@�0�rτ����^
��։�ث�b�%6���
� �@�f��;�So2Wi!�k��{Q(�z�ե�:�W(u�;�/9Flԓ�Y�"��[�f?꯾��H��g_��}?c�i�~���/7Χg������}��y�� ʁ�#C��{^<.w���Em��J�����/+Z%���k�j�k�L.��]��<��}��_Z[��ʿ˷
�Ao��R����K���ua��6�i�w3�1�ߪ���7�-��KG+���j0y���4��/�7�����8=�r�\��[���5��̺���Y�F�� �aή~��1R��+o���yC^���u�.
������0'OkL�� r��=cƩ�ݯ��e���,���~�8YP�xj�aH�����e�U�SY��@�o�{ru���J�MAI���e����6�AN�z^?y�Gu=�ʝ��������Qo��q��{͉~{��^�M���{��\�|�mԸ�#(?���N6��I�F��k�M��?fj/���lQ�Py�}Ot�Ϗee�yl{����+����ϋsn���' �N��>��x�2�IJ����i+��=Zn�C���nIb��Ǆ�mH�����T���\^�I�h�'jQ̏v��pv�k}]�ʾ��|�~� %�%���ǵ�m��
m�T�f����� ��+��J\�ژ�w{�(�[j1ʝ��Z��v���n&#���`e����%�3��s�,��.Y��>���M��֘p�[�F�:��2���53댬B7���Oo[�Y6�"qȗ=����yT�8s�	��hͫ�S��r߽KѠԢߜ�ϰ_��E���6��ռ�I̼<�w���{ �Y�9�Zm���J��,?Tog���r����k���l�}�����T�c�U�K�in�f�Ԟ����:�����(���R�=�w��0vT�a-����B���ۗ�3:k���múe���dd�D������ot3F���Yq./V��i��_{cg�SiD�K����n���6��p�0s��+)BWe����G�o=�ۇZ��*�x�S��Y�����u�J�zK�;���!��&�^��-t�6��h'
��v�wsQ!S�PR���E���`CO�[�#�RbA�.m2�%��Gv���iW&t[��k�85�v��YVT��3_/��u%Wr7� lZz?}}H,��^:�76q�0��K��)@�}�i�y������ދK/��]���}����_�6��+ ɂ����Os�X����O�w{�_�^�4b���u$b��1�ʵ�-ͷb���hQCtCKz��p���%^��^��tzLo#�(�?���D�J�?oٲa���-�5L�[ڗNH7�׏<r�<�|��0x�О`��}R����
�f⑪�I�=wl{��"&�k��$�9����އ�m�H�5@=���Y��՘�4dU�	X�Vzj35�B�1-r�8�`ɛ�l�_�3+5Ҹ�U�S��R,�(�.rS��{VTn�w���ظ�����6��.|��^z���k����Cf���D�|���b�h��5V����>��6�9[�;��c=��ݧ���Ug��]��I�1a�ќ�K�܏g{#5�λVն���vt\�yYY�[h{��+)�1Q��hN�~/�\�56���g�o�]�����kJ-7��]�:�2v�O �]�it�5�־����t]=�AT~[�OY�V��tŏG$2F[��u� ��5�}�Gѻ��M֦���t,n����k��xמ�yn� ꖖМ.�ݯz�E��^bo�{]b�U�R�秏fyٞ��/v�_��ZA��W�ޫԐ�ߒ|wr[x�Tˏ�*���
&/V����u�o����Fb�>ǯ0��j�Gg���y.�����o�T5ap��7�lz��N��̘������\5�=��=A�k�yT'���zkޡ��섗G2 L5.�W+�m�B��pכo��*܅�*� ���=UwN�`��f�X�'ܧ�߹��w�5���z���i��w���l�����U�빨q �]����=��l쇊�M}'���_��O����A�RF9�hC
6�հ�5�Иp7e�Ά_H��h��?_F�����x$�_�(;�oJ�$��)ז�m������=��
���ƕ��FV���x�0��]$����[�.����/�E(���#�G��m:m#�U�dE8�p5�2@���I��u������������|�y�Q����k�Gͻw'�rS{��bv�2�>)��v�p�<�g.'�&�i�lӁ>wc��Vz>uw�U���b�������W�}ɼ�08�>�:��E[5�!i|0��D�H�1��-~{b��G��O6,x�c�ʵK�L8t�ߑ��HN�9_�6��sb���F����}K*�����Y��6mG�ԭ�hkojj#Rbk��c�n'�;P9:ϳ��P�G�;�38m����zj���o�v��$�j!yÚ������E��nוɭיU�'Kf�d�k�=�Q���x�њ��i�j���Ûr�~��n��)�<��ԟwnޤ��Zu�F��Ҽ=[��ו��djz�\���^��{�����P��N�Z���w�.�w�MϠ�����'�
���Z��:�r�(�^�{��{KH[���
ǹ�V�(<ӤM��uw9�`iaN���i���-RY*�˄�?^Cn��f3�P8����-S�Wt����q[o�lZ{nOnk�(ͪ�b�^��sרẸg�е����y����w^l9�H�+ s�I�Iӵd��D@5�JW%/�k
��9���mJ��nF��w��vݣ��8N|�����5x�U��K��e������%�8��g�K�l/���Zk':��8�fjX�WfjS$%�o�q����쐔��烺OϩfW�L��V��~p߮#�e&�_�^�aL�0��{y�OS��,���\�m�\՟m�t��~�p�_�,���d�5�����'���.f�{}�]���e[i{'�w���e�*�RO=��3ܪ���Ǳy�ȗIH^��6L3,UFɸ��/�N�=Y����y��݇x�>O��y.���B����0�'Pɜ9;5,/K���u����}�����7����A��B�f4����
3}v����E=��r_����}�WNmX����3	c��Za������Qo�!�������Lk��L/P/�_�j�/=E���Օ��6�k���M�9����a�R�9�K�O���t�b5~=�䶫?�o=P��k[�;��=x���7���:��j[ڞ[�? u��}e�1}�������}T���})������vwJb 9%��wF�WP[��(�uNk=W:3��Ą�|���R�����U�]G�&"N��p�v�0��X�XP;�=�_�0��$��՟(��� ��3i�N���&(珞i�'ALl���qC1�R��=.��uk���<�l��lY���7g.i�$��1n���F���]�Z"]w��i�Oy&4E�)�a�5y�
�+K�݉�d��я��x^[�ۭs��gs��z�D�[��֕�wؕ9JNY������z����K��t�(�S��{A)%�YTY%nS���(�1j}\��J<|��ƦSg�Xx��H4�[N�O*8^�y�r�㉸�[a�k������@ITx>jb+s>�C�b�3��e펴%%k��L��dף���:s;I#�"��b�(�V��6�Ra�2Z��I�ʝ�;�]uGAq�U('��qlH���N��N!��{�\���c ���6w+��v�ZE#���%��ݡ�nN�w�1�����Ä�����5Ԡ���U�%)�WVD"S2�NFS��1�F��K,���)��u���Ove�ʎ�TpA���?j��)"[�a�z��&�\���M�m��[��^�Yo=Ke�æ���+2H�r�,n��CY��M�҇K[�uTXwHT;�J{�(�3��=x�+��+������C:�ou���2����@�-�ھ�C�{���Fd*dv�	���d[�oB�� ��0<� 7���*��+���Om�<)m�?us�B�}Ю2��sNd�i�t��r�<��)�;v��:��yh�kr݃N�&��</X��.aָP��p��4V5p�dhײM��z����pT�����j�й|;E����%u�&X�k'OG�5(�[�i��J�}�tS�U-'�=Pe;�ih�9�pc������n�FX�/i�؃�w��]6f��b,F]p`��v��&+��������6U�;Ӟ_D���L�w�;NKڶ�èjyE��w��0���Y���٩ޫY�&���*b`���J30?��@�����n�1J��u0L�Ɋ��k������An���_u�hĢR�8�6YTY׵:�w3#�s/rl�PѪ{S8cr�˗b�SK{rfL�V:�plF+M�6��dG�ǯ��e_�����맷���@�[˷�q7�w�5�J*�]ӱO\�b'l7�/(>�W��f�iKڏ%��Am6��ST�z�͜�ڲ�1�2�P"���i�d�IDt���f���7��;�v� T�4��i�1�;������a*<�&vnZ��srܮ��m��X#���z�F/b#(�
�a��r^2y�Yhy���������[�W9r�,�խP�!.��ѷv(&Z=�*9��p�� Gf���i�A	��~��J!�?"�JL��%(2ZZ\�" ɣ',�%��p�"����[02ZJ2�02��1��p̥ʜ�L�0�Ɯ��������r���#+0��h�"l̜�����jd���C&������i��",�� �(�J���(22��Ȫ)h��ʜ��b(b'3!*ji)hs+0Ƃ�̠��3	�"��Ȫ����X�L�rk3'	���*�c$��	G��H@�I?�)Ҧ��.�M3��5�b��ݖ^r�.by�z�����-�^wM9��{��P+��:��z�Kz���y������(rr+a�o������q�=��v�Ѫ�Oe���sN��p�����r#�㐫�s�ϑ����N1NĻ��m-#'Y:8�8:+{e�K¹1�9*�^w;�>�W�Z��EF�M�|�e'��߶���� *8ܶ���A�4����5@ک�ʌ���Q��jM��{C��م�h�S��O_��wz����_�����;Q��\an��v�v��	UE^�A�X}�ǔ�n��aJ�2J�������5c���u�X[�ЪWJ��Ɨ�S�8j���D'�-ͷq���9�,�h�G��jQ���!k����c��V��
Z���~�~kq��~��s�t�M�9��R��\s����2��Y���4��������n���By����uyɑih{]t�=��w/�=W�(n ��jĳG�54�<nô*!��D�5�ҥzf��fZ-Ÿẝo�fv	����Z�bS�M"׻<A�:0��Y���� �cj��D��+��������b76���v:�w,�L��\�wj�d2p���Z�޽���nkc���8PT���u��ٷ�ܹ��w�
���<-�J��yUG�����%�����s��[������e�2b�i��]S���U��W��|q��C���{�)�Ox=��c�+>�<�w����[LKn<��nc�:�H����˳z�yxܺb$)��y;�|�}���i:��jP1��vw�cf,�������
������}A.fyV��o(��[���<�^߼�q�SH:��c��H��q1���p.��or��������^�5�i������kE%�
.iZU�f����.���i��}�����=�{_M��v��l=���sg���߷��{)��\���Pڃ�>���x��G.K�{�Y���p�'&����k����t�0o�9�k�}\��i%���7��Kuׯ���*��6�C��	�[�N��<}`��G�at�9����K;�I荭�f�i�˦��b�����z�mA�����;�t΍;Yk��rw�����^њ��r�*d��%�v�*�е��9Y}�],F�+rY��i�v�&WN��Gsƞ\�0��&+[�A'��He�i�VT��X�u�H�EԻ��g{��{�z�y�ʆ���d
?o���-��9~��+k<B�Ӯ ���V�t�d�I��[Yy���7��bf@�o*6f�W�Jt�����!k�׻����_�aS�;��u^`���Mc�r�<EL�c���?�@�zo�����v���[ϳ���R�u�RE��җ��%s�.����FPtc��/r�O}�g�I��c )�cZ�f�����M�����
ᛉ�Jv����P2�
�:rrϵ�i\�7�VfH�NYU��ױV��ڝI���y�X+��F����f�'������2�>�	e{=s��~��u4���Cn2��3�����E��H��92�x��綦UN��~�����=�k��٧����� >�j��0J�[S�mX�c=�.x}�3����E����L�wYY�jǚ�1��̻<T;vRR]�2��֘y�msČ륹}��:ً��7i4�:9�A�8�����D���p�!ٯdw�a=ֲ;lU�ڕ'.h��;|�r�����V�s��o&�
�zMŻT��G�k�����e��l.E�����I%U�y�]���Y�|�K}�5Y�6�Ww��#{Wt����'x^��r�����M�^Qz��d�����};�/j�-!k�KF��Y�J����-���-�U'�:��'Ӻ�s���=̟w�c6�.ƶ6x�P:��J���1��O�i��J�2��<ب�kpOO<��v1�z�˨YT��Y��r謾��-�w�u��K�����SCv��y�l6�B�W�xk�J�5�����#!�mI�wt]|�I�k���%����5��}o�ze5ꋖ��^���̡�O�K��5��;���}��n�ѻ��ro�����gW�J1������;ڿ=E�0�x;$=x/gyC�+�yn[� ;�p��*g��D-����q���xӯA������ص5.|����o{�bN2g�{�(K��Qv�!�Ƶ��^��Qw�.>ԅp��Z�ӀiCF�<&�u�Џ:��"���髹�(�����\���K �LY;����3kL���p��]&���X���Z�ա�Kn��!��7�Z�)V݉�N���4A(�Y�Gm+VzV������gf>vq����v��f��\���{5�$g��kL;ǝ�78��1߽Yس��p��i�V�MC���^��~{����f���z�C��x���~ç�:[��<E��U�[~=�g���7�y�gw[j�%�f���W��wuny�p������^c@��{Q-��y�ڪ�P�.c�ٯ��Bz�xg�rV� ����u��_J�w���M��5!|�Ժ;�dy�3'_�%�S~�zzvg�g(�T�l�SV����<{�xO�7+���w�rK����H���;�KM��	�e��}%̵w�=��讓�V
�u��lz^�y�_jM睧�W 3S[�[s�~�jy�6�A�k�=�c���ߖ�g�����o8^�A����~
%��Ǟ��e�����]'_-�ٹy�s�v��}��xq���s�J���I=<S��l����s��U{+��u��t�1d2����*�;��=d[-y��D��x�7)s�_Wh�(���}��#\�����6� s��I��Z��Bٗ0BF�WJ��J���`���c]ǎ�K<��3O����g����{� �(l���v�bՆ��{�����R��y!'y��5���~0�%p()��4e�Q�X؟PF^Bn0��]�Cu��[^Oa��
��|�`~f�ɍ��DQƽ���h���S���%�d[P�G�SJ����w����y�8�:^�b���
�xF_�mX��k9�n{��9�)y�������o������Ӿh\)C~�G(5|�sz�9���o��El�t��{\y:��$��&��#x�C�-:������D��޻�]����(����7�'K��6�eC~��~3�lR�<%�*A�(���=�>Z�y�O�ߚ��U;=Ի�������vi�l���4��h����8���N��^�r�|��z�L���^�j�ĚJ��7+�yKHc�
�r��o.��
�÷�v���@�=xxZUH���Ͱ�ٛ/qR���]p<q�t�lɨ�,n��%^��t������HZ!���He�3o�VF�\�#��=M�&�jT6)���;�nt�AntX��P,�%���䜩�yiiKKG�u�&�'��������ݛt`���VU��"��wf7��yM�F�UO\[�9V߳؏W�,�o��>s�5�*�+�ʍ��5o��i��M����l{|rc3�u�Ŕ��,���n�#r.�:��F�l���CtetF����y:�5�hM�]��k�����bc啻�e�#���O��9������~���i��Q��N=��u��W�-J�)�n�7^�m�d��/#=�ez��@X}�ef=�媽{��ߦ�r�b�}���n�����j׼�|fy��)=�ش��/eu�6�����lT��1���oN _��Q����Le*�y(<�"���W��m�wc~>�-#)ьq���=�5{����]2���q���k�׮�z�l+f�.Pw����g,��]+=}a�Û z�������]�i�ӏ4�"(8�ml�$�=�[d���zHK`�/+�����0�Hi
�ޟW���:z�SO������죴Q���o{���KZJ��E��?��îSZ��4*�p0j�S�@l��=��YxʬfZ��ma�g���ԝ~߼��Ra��y�#q0��:�M勞�E��=iM�gZ�U�i����
��O/��ܛ������Jx�w�r_U�N����JG����֌�[���\^�3����{�K2
.7�o��-z�����K�W��~��}6������l�}�z���`�+q.��g�ZqHKk3�3\j^{G;����3�J����Z\J�'�FZ�{HSq�G�[	mx(Zx�)��bۅ�m�ȴ��:���/ӟ��[Q�g������:�j�rt�2������)� �����ҔZ/\{����z��[�T�J��0�V<د��y����1��.�E���:^}.�g��%�r��K��PU,T�0��8o�m�Tyo�l��˞sm�zq7�lx�0�
*�Q%'{tU|�T�$���
 ��Y��6�btm��{�i��lW:�J��������p%]��4g�5d��xkN��,�j�S���_T#ŰP��*���K�w�Nû�I��s`�R��㑮���D�w�R�a�q�M�������;�oRY�u��̳<䧕6M�%���	�\�=[�
3g��(l�o��s�t砱�� �rn��ئeu����$�G��7���z�����y'�����/;Vf{0��/k������aW����
���TK�i�~[Y�*ʫ�kk���FJ�R�VnI�n%K4z�4�7��6�oѐ�/Q��5��^�2?{��K*��c��&�-;�u�$}_%�k�އq��%��ћX�ow�7]���o*�v�l�5��Y�-Y���U&�@H��=��=��t�}y��?u�T��θ��߯��"�?k|�  +���d�(z��������b�T[P2�?U}���1�-m|=�Q�Kjs��Փh�z�$j�˽�kW�N�C��=��Cߗ��ij�ZZ'����+�%���	�;»�`�Ӹ�
����ns�~魚��j�
�װ��gĠ�>Hš��up���JwO��v��V����ެĩ��du%�ͨB����S�;�!�MU�%X��_��r��Z�.f������J�T����Jƨ�.��t�hN��M��H��C�q�[����,�Ơ�
]e�Zkv6���ss�]�q��?|79�����Ã��^����y��n8���+YgU{�8��Z��A�W��,9��ɯ`��^o�\~���R��:����mcK�T���=��v�x�VnG�)7���wZ�\}Tf�����~p׮o\��U�|��U`Pz�$���4��[~9bS��1oݾ����2xzn}��OOvJ�xQ�'� �u��'��D,�4�a�0�Kn"����Rɯ�O��X��O�}Q�w��w咖�[���=^��~V/����c`l�V���}����������y�+$]}^����()8�3���V�,��M$�x�=)���2��+���m��5谦y_�_:���̕LOs��f��A�D�^>���./S��
Pݤr��Ac�����bY��N{-�}Npn�]��Gtt��&<�8o6�y\B�Po'����u(�^���v��nSut�R��n���BGB�����fs}���)p�@ٴ2�=�7������R4��%�N:vg;炌Y�5�aR�|/���l�~���+e��Cj]����t�MY`�.϶A9�t�>=��9�n}w��G�c�S��XXM�8�YEL�@p�B���f]wq�(:*�,r<U,���ݡ�Ed�����:b4�������P0-�K�[u����jE�pU���1�)�0�$��cpܳHݭ|��:ه�������,�+�p�`�.R⧫�)�w�Xt����u����b[}��k��,RL��^��X%��e��ګ�3;z˵N�\
��u�]|����L����M5m5V�'R*�e���1f�U��Da�yTP�⳵��ѹ��w&�I2�쨵O��bεV.�\UC}�G$��\!N��"k�}%����Ab@CYH��M��w^�5�0N�sׇ�G�JD��2��\YW���`J�����l��FNJ����J���ݙ�ptI�T�⊰�x�x
�3E�&�,0G�َ�~�g�X���s~�n��� ��6eu��1��}}��Ou:�Z��ř:�����hQ����� �[�3/����sO	7e�ڻ��;Q�ka�S9��ը9O/�X��y�ٶKX�Mi�M�2�,��X"ݝ������V�h��	����Ev��GPm	�U����� �ɫyt\�Ǵ՜J���p�,Ӥ�A5v=�� �2+��$���c�-i����bh�2��]Na6�]@�l������ʝ�KZ{]�)��E�Z�3ub���r�0�v�g��y�J��Ӌ$��4���
��ięф�
��r�o6p�:e������b2C�tz��#�ƃ|��	[��2�i���0{B��s�.�}ʵ]��.`3DkzM��']�H��W�{����;���#��]u�Br�՜���-U��afe�{%��!ܩV^�:x(2�]� k|�GO�{��s��ap�v�`�P�3K��	�V�y�e���S̭M�g����;3���g3��.'�k�4��p���ՙՋcu�Ӿ��O��s���q4h�4f7����l��ɱ��4�N�0�xz6ݶ�.�v���SM���5�U��+g7g:�fZ���Z���u΍މ�z-:���f�i�����Kq��j�ܖ.�@C5>�����y���J���컌,��s�ysO�Sۮ�t�d�ٶ�=� J��Y]#ҮP��+��v#���}H���}x�::���pW�3���YX)k��cn�Z���^<�+>P��e<)�:���W�f�O�k�V�¶�Z]-�w��92���i��&a�ۥ��[N����qփ�� "L@L���4aE��QQ4�P9�S�D��R��adDAY95FFLFfM�d�dQIERU�a%e�K�c��JY��YY��PEACCT�E��$@P�R��aEPTY�ĵU�afdULFa�UAMD�DMP�f�f`AU1fTdE1��M�E2Ff11c�RS��EM���ED�b�A�Q�a94�Mc�ĕ�VfSDQ��Q%fUVc�Nff8TU�S33�FREYTEdaDUQD3UP�AT�EE�a`S3CDf`�D��EQb:���ܓv�nV�I*Ul,d)}K^�Tz�)��neH��|�we:>�y����F ��2Vl��r]�i��q�An�l��Kҗ����|�¨oju�'[�g�Y�F�����<\l^���(�}�47�T�7�q�ͤ�˅�[p=��U��LcE�U�!�������q��6�U\]�+ި�x�ٯ*3�n�T�iw��j��/q�r˵Y�~���d�n�J�����>�W��)��x�)���5�j$����o�N��%i��|ғ4i~����y���O\4�VQ���'FC�F����9,�.b��7���7�]�3g���P]^߆��SF�%��3J���k�lSI��)�y|��{l�~��E@�f�Jx��������V��6��ڲ������6�μүn=R��=��~ɺj�@�z���Ux�W�s*')�j�+�߯�8o�p��O,�8�4�r�V�!�.�g�RW}�Q���J[u�*Y5�I��5�Y��F7���s$��we���7L���ՉD�K���9�Aק�/��EhH���c]�|��ö��a9��Vvn���Õ�pS-��q��d{��F�ܜ�]4�WE[RI�.	Rt+Ov!�3�'V	����Τ��ʚ�"$ԅ�N��y��/;^H�qw�[y�+��:S�<pڍ��V���)3�PR_:	�;t���Oyx!��A�΂zN6g�`j??n.�'��R�o�>x��W�$�x�;���>�t�}�?l���ν��z��U�5��S��J�^�CS��2�֬7�æ
#:Q����^*J�kɚ"[�䋝P�a,�d�W>���|�M�MkL;�7��R��!A��]^�~ܞA�����ꁷ%�K~�����~m���yÚ��c�ѳ�3����Pm�)��^$^/[Ϭ��Z3k<������9�zx������V�?Z�������~�{��~�G�}iv���~��٤�ȉ���2/s���x5z�����N1����r�-c���U7>����)��z�O�ù������u��u�o���~SV��Y(qK�yw��ұ(i��N���B��T�d�p�7b!���c��&1F�c<��.J��V�I���[^��// .^�'�{��.vc+��W�9l���ڔv���{ng6[8��I}�#�O�bh>�N�����FR|J�����XpN.xV��(#�PV9NBĹ;;cf��o� ��M�d��;�6�+��M�J���n����e(J��W��b�]��_x����6��˩��㩨�k_�;S����^�����u�����{���!ٯOM�VǋL��^o~�FhyH,ɤ�(�)I�-K�\�~b�Rga=+�g�&�6��7�p��ڱ�oA�(O��P f�o�ږ�}��5��T#ez%�k�g{��C����?R�_��^}҃�~�UF�iԽ#ڊ�6Z�q��ɠ�j�KՏsKi\x����o"]3H��dY���+���WyXp�@��5��ƥQ4{SI@oC�fШm�+G6���e)�T�L�|}@�,�sR��_{5�bG�k�����/x�K�j��/u����J�_��=_<:�N�O�Z5ΰ߻Պ�)K���8��r�gÖr+�sk�1�4o�P��-�w�LtR��;��ۑI�y��>���)Ҩr���ptsG������Z9�����QE
����l�-@�R�+7
o�3X�m�5�6�i�6��y�����9Ƨ�{.Utid�����ӌ�%{#����~5���\��_���%�X��@�s�����Z��'Z�c~�m�����վ��讳���xj���Z�zJ�Iռ;ֆ��-y��kW�����~������{4i�֕��티��Q�S���{�&n��+F>�G�������kf�)�0+oy��'��h�/ZZ&��Ч��PP{����;��3c��zCՇ��&zX�]�g�{|r���*�Ã�/��{��߾��\le��Y�/s�S��0\��t5���E{Z��P��|k����t��	����qG;rǽ�q�1_Z��p�z�<ߊ��[⪲���~�������t�6���JR���?�r���U5�M��8k��)4�~2q/�>A�鐃^i]V��zC�V�';!⥒w�����q�~����ޞ�i֍��њ��q�pCz9�le^���U<S$e7�C&�ĥt6�
�a���y��
ˋn�&�{yyR���5�{W0���f�-ݚ���Bsb���}���G���^R��]��)\��㔈���j0�=6-��L'mi�E����v���՝8��~���`�q��5��j�^�x�>���t��d۟g�nW��cI����kS�-��)`���V����xrߤy
Z\�/=�����m����DF5�U��3s�F�byN�N��4:�,�Ľy����z��}�	�G;�Cb��y����8��ǹrܼ�[���ofsZbjq�
�F;#P��u;��xDvu��ԏ<;����h�|��R�j��fN^�f�{ޫ{<�_�%�+��f�'��D����W���JmdKf��Ny�5�Ӈ��w��|�,�]�Mɰ9��=p�ΫW�h��ݖg��ji��=}���U{��o�M��[72�����4=^O{H:�ih�@�bźi���*LPv���ֺ��>�%�R����y=�����k��к sZ��]s�/��^3hT�[�y�W�d��ޗ�A���9��k�3|���v��u�(a��u�) ƍ���(z0�]p���Y�Twk�R7[�Ma&�n�N�Ͱ���Y-d&�m[�ڳ��0^��9n+�zɔ9ە|aД���}��7g�W;�R~c�m"�ԛ
7��s-?*�o�U1�PU�g�oJ��߶*q��+
�Ij�2�5xi�)��G�'���~�/�ꓵ�y�A�ՍV�<���is��eZ�J��^�+��~��ϛsG+!L�~29�ja�����0������B��FOk�����+r�\l��m��|�-��y�lʟs���x��n<<��^�-�e�e3�a���{�|{���dZ�5��}�@!�w�ʷ�ȹ�e�y+�EW�n5��M+��k����o%�5�!N�[_�l�6�F/x2�g���SR��}q��Y�+䵨oC��<g��\T�]v{��6�uE�v�ƫFTU89�j%料��Q��������^<<`���03/%�qi-��/�[ʫ����HO�ɿwL�W/W���k���=�����M�A=a6;`�\#���W�U�^���f�U��Sh��(�yH8:��u��[�~�w��\���(&����1���ޓyKȦ�7tg�[Ò}wp#w���峭�M뀮����!=֏��� d=����������O,t��A����=o,Ƕ�E-���.9V�^I�ƴ�p=Yr��Pҭ�<�
t�x3�=�����>��K���v�|��^g�4iU��L��}}��ݎxk^����eC�n��z�/�����ܡ+2E�%�}��0���'���R��<~����عϻ��~Qf���i�:�'��G�����M�G~8��Y[t���
�69�5�}�=��3AR���lΕt���zXO(��+�����ʽ0y�_y&���ىp����o�Ǖ_��9��v6�w_ԟ��,R��*1��9����C۫~���g���]�n>�z{�������JO`yjb����`/T��6��^��&���e��:��v}��xQ��m@�-�����fs�zZ;���=�{8�w���F�/G��~�-���&fS��7,��WE�\ �ô��0_Kq�|��d<��l:�����obm����Y �1�[L^Lߺۏ R�5��wW��n$=���������2>N��9*^h��YgW�����;t�VPjV�i�}S�l�Q��b����T�w5��m�r���o�vsUʓ�P��O����+j<��Ҹ��{��?3�L��_���Ǧ_��Zq�}�!Z�+p.K��s�`>�>�吗����P%�f�l]N���7!kD��ד�q3}��sY��m>����D>G�ӳVu�ɱ��ul7�Lo���\.ҧ���[O�Z�eY�X�P��ֹ˹�<6z���I��h��5�^Aۨ��{�{^;I<��ޟj���{+�vR��Iʕ�����}㊩���?\��l>o4-�H*�m���\�m����睧M��֯��k��{�ޚ�K�w��ZF�����OQ�%Z��
ʴ��t<���w��W�>�1.�_Ǆ?6y	�ܽ���>��c��]�=+��J+޸~C�"�p{��$ �k޷�!�]��6So��m(��\(q�mg�m=��c�ى����T�X�>te��\,}Zi9ê�.�"ΰ~���mYU5�����K$�3"���quf���(�;7ܻr��ϖ����L���X����r����ͪ7x�-`]�#k��\��Jƛ��~��CM�s�ӆ�1��
��B�
�k�s���4�z���s.�o�U`0u���nK�>؛��^�I�s�*ܽ��c~���om�{{Q��U�d��RQ��9����V�����9��5	7��8k���,���i��Ax{#�{�׆�����Q6l{��h����K�Z;����D�I��P-��s��沽6��>�r�~ �o�q�����g��������u	��Y��j���<�r�!�ض��r�De?���Rq�|\w��wO�u��Y��b�h��wv��V��Ik���M�El�"��ڈ{7���͋��I�=�Cuü�襍c_5�k�އl���L*B~�G* ��_[�g�w�5yqbz�Þ�������D7�:����h�O���3sk�O���u�������5��U�bʅ�䓙V�K��p2�����7yYb2J%x�P�R��IT��&W@t��Lu�'Y����lX�C}Hݩ �E�,v+��38I�m���X�ŝ��<�`ڑ�ϮE[:/�M�l)Zѐ�,�4m�����(�4Vt��y�7*�=
���M���r�L����X�X�z�ΑB�'��\meYo~���r[Sy�9��i���>�ޯ
8Y+�L��}��j��fr�&��_���د����u�N�~r>�)�t�y�GX	)�x8�z�R}�~��8fxIg��0���lw� S�iz<��CY^
֞;�L�ǝb�Mn޿k��6�|.�誁���^t2<'���gƱ������k�1Z�b��x�}��,k��/Ŷ�ݧ�.<�ſxI������)BW��	���M�s�z�s��Ǟa�Hf��I����v��$���2��W��\y�~�8Yg4Z�Җ��B���)������l߲��f>r�H���K�V����&sɮ��--�4�+1ㅔ����7b���l�����o�j�k�]�Y�L<:y{�]������os�ǲ���(���*~�v��u{��"��oM���2� �t�S�}��K�������e`-�P�\5*���'�7}�w����jV�Ɏ����u�Jb�	av+T#�{�z��?Xl��a�����T�SK����+:��p��ݒ�����Ȉ�f��a�Y�5�e9Ze�s7��]:�h��T;յn���\Y��+v:j�䕅و�s��/$v�]v�:��K�yt���`����Ğ,��?>ф��0�ɒ�y���w�p�����.Ê����*��-J�
��,�/���k�]�8������KTj��s���c{�R�ϣޡ[�ܜY�٫�fSBr�(�v�V:>����S����^x�WՓX�3SVJ�Y��9�����3�6s��fG�$�J���nmM<�[��v2F�qmG�o{�:���B�F�JX��m���� A�D�㉖.*z`wݤ�Ւ�����e�l��z�4��})�GNm�XR�&7QE���6�d ���Sj�x�mX�HmQne��JxsQh�c�v.��M�
r�Y]V�i��I,����H����� ��u��8����vi�si:������pN�֠�[��1����̦�ʺ��i\��O�3)��V�ؚ*h���rO]�ˁ�vM=�3D��d&����X&�j���И�Ca�ˮ������;˕!���晙\D,V�;�
c����-�m.�ըQ�ڲ�*�FE�����l�v岫{p��J�F��!B��r�w����
3�
���hPG��	u�T���;/����o��eKnj��2��u�/+5保�V����bR��;Zj�;B��ˊ1o3�y0�1]�	y��_I�gf䤇V4�k�a5s^��B�u�p��d{U��iA`�-�Up_bɮ];kvI�h�b����v��R)Df�]�ڛo���-�J9�ԉ��L3i���X�=Tet�@ps�T��'�]�>��eLh�6m�L�uGh_JNl6B�d��0�p�|�iG��#�M��Dn��*�pN+Y�]d���V!����o���km]Y9qf��|�N���e}Su9W�w�;�:�co4I�n`�����(p�v(wV.-���k�S���RA^�׌bL�bZ�I����˾H��]��}����W"�F-��ywp�!��1�%���
Yb�$꘺�n6�WM��G�]�ܞ�y��v�_�Q�0a��f&03��p��1CK�㲲��8�`�p�uD���X:�s;�D�o`A\��s��M�+��kjl��Qn���!���>-@�eպ*����z��	����wt'O%�&��ͣ�b0,d�q�����ܗ�\��w�NVEzԺ�u@�;��C��=Nu��̔;[�ƴ�
"���N��Q�.�I�f�h�;0�������2�S�6/%7�&<��NlVc]j��=[�U��r��dq��h�]N�a7�,ru�vo<�5����������Ե�3E3o2��bj�1���*�',(�b**+2��**(""���� ����&����(���� �����
�32�"�
Z�"i��h���d�(��"���� �����H����j�+3
�(���*�"�����J)������h"������(��)�	����$��"�b*
h,�*���i�&���(�r, �h���*"b��h&(��#j&� �*Z**�&h����� &X�J���d�`���*K,(�
��"h"���
J��*� ��)��b*(���
�fJ(b����*,��*�'*��0�� �L�&*�)����?l��z��������Q��@��H�g��)�q��p�V�I��.�V��q����55���	!��^��=/��G],�КP��a]��l���5�я3J�Y�['ݶ�d�A��^m]n�\F��f��Z��oC��V�]��k��x�"�ӷ��*�+6�=���ҷ�Q���H��g5��n<�zl�,#I&ߦ.��YH�CwdLy��r�����d����sU��2�y��y��w���.S���?h�=n�k�Fmg�Y��9�δy?V�饭[%�ަ�u��iO���t�[yU�n��6E����~���&�j�d�:y�r�����n��V�S/5�Ǫ>{G+����.����A�/l�*�5��ٶ'P���VR>�5]����>�$��-!zf+n�0^��9K՝����s�x�_�j+�j<�8�]�\�)�����=	.~���o}��8ލ��(��/-e(J��W͊��M�+}�U�0�D�!ϵc�6���4
�P�걙�Q��dj9ГWl�m��QU�,�"��1VFy�����65�a�KUt'���'.L�78���_T���q�V�b��ȹ8;��l��:0�7��vn;�:�݌_W2V�����yD�^9��M��28��]�=_'���/�KϪ;d��9�5��ǐ�̍��׷���pׯͽ�i�W�~�����!ꨉ)<��6U�S�d�Y��Ҽ�Ʃ�����5��,��Yn|�HK�n��9అ/�{����#h8m}�Iܷ��{������Q����\��ίy�>k��~;�R�����34Pշ�m���x���
��>��R=Ϯ�c�e�e��<���y��VM����,��M%�oC�U����3K]�l�}5��/'`��`s�o��f�=�O�/��R�1n:��
>5j�RSZ�M�w�%R[�(w���Z-���bN�h;�{���l��n�牵3�ɉMǞ�3u�K����g��|wC}/_W��1���Ӭ�텵�p���X��E�*�W�Ꮃ�uyyc�'VSΛi}R;�x�n&��������n'W�ful�5�l��Q���o�q#�O�{.Q��I����Qp�;�E����m\�)Ֆ�wp�w5_�C��C���Y�B�jv����۬4��*J��K��\,�z�����b}nv�'�ZPr*��[�5��vz����W����o���)���LD��=۠w����������r�TG�ƻ3��.|���+a0]�CA�7^��z�ޱw��ŋt��x5@�3r���z�>���@�/�����I�%(���}q_i��mDK���5!��u$^z��2=�f�*���8l4��X���\5�^����2`끊�q�;.�-L����Vf�FV�U��x[n��m�ä��*�m��X=��f=�	oэ!�����NPڈ�ښ�����^�8YP�yp��>!K���\_���5�i2�a [#ӣٷ����h��3��������{�#]����Až�6}B}��8��}�Q���{����mT�^��y������^`����:�4�S���C,���C�A�1�[:<�����"Q�.
�1wI6f.v��]�\�_V�5��в��k3���L�/�z���b;1mՏx��K�o��i^l��9����:B�3X�{a��Ԉ:�ԟ;�#�l[�(�5�V��f,�f�SY�9����AHr���$<���u����۸ϋ�i�el`	�}�Q�b��yX�Ӱv�L����庈ծi7��L=�}�	�i��u��d�9��G�Gs�^� z�'���j�{[�6�g5�&�q�
�tF�K�������3��;c�{�SH�H�K}煾o��N�4���y?{�3�C�Z�ՠ��d\:{y!x�s,��6��mM��s�~kO�N�E�߫�+*w���}��kmm?-ߞ�v���g�.a���V�)�̻�n��X;"j���w�%N@r�N��{�(��f�/֕���.-�Ӄg����t��/W�[�YFzx�ٝ�_�s�FޯU�zҾ��%|��'6����y��<+ko�PG��w�1Z�b�t�\*��O��g*|ڲ�0Ht���Z�P�gnA�T��*�9�e!Q{}i����qz�L�]�n(b�0�ڽ��Z�R��Z��r�F�2�鲻�gR�Je��L\��eKڽo.e����t�h�$νy�⤍�ʼ��7�NYNظ y��|�2l�ܥo�ns}7�'`�ۦ;��-�W��%�/��1b�.`��1Ͱ�\]����h{~�v�{���&��r��W[��7c1B���{3~Z1ż���� ��`8d�^�>r�H�ݗJ�M����53�x�G<Mϡ{#RY����8^w��7M��()_f��L`K}��8�+|Az��{Gf�:�aS�jq�~f�%�5�;�l�`_��O5�I᪯u��s�ρ��Qؙ���Ұ��~�m�ȉt�B!`��Z|q����/o)^!S�`��5/�4��ٸ������l�c�&�j���r�[�U2]@j2���������1"齩�i��1s:r&P[�kwQq�<�H������������=�Q�n����!q�l{.���������'�8�{H[W׺��FӐwu�{����x���i�9>
zs�>˗��F\NY����M�VC�;<c=/�	����}�,Nlwo�\|�dϯg�F������ϐ����r�;1뼭ha�BMVSe��i�Ƿ�UF�J�t*n���y|0�Ѡ�?à��<� �Gv���m͖���f��|�0����2�s�<ڔ��7���B�vN�.��c&�d�j���$:����s&Bu��c���{G���;&��C����*�;��W�u5�c��)qy��v����<)�����̾��~��O}�P0LMߡ�G;E�O���Q��D�0+��/G2���Z�}437z�<�F������6+l]ߧ�ߑ��G��faz�JE��Ma�4�^�0+��Z���t�ݲ��o��U�G�xZ9��=����x���?3�몑��� ߾�T8?@��#�=��M�a�U-�U��Ei�j��ԃ]T�R�h[YR6��I:jJ�FUC��<��ܸ��/IYs��W�q�����.����/=�qܧ�θo��yh?�[:	;�,	������b<�o�x$��x~^������q���F�/Oi,��p��5�{���8 jڹ�]�OL�x=q�"����b���EwRs�h`�'�m�zF���ˊ�a�i;�tܙ���m]Y� b� t��d��W)��FXW��=��;c�����t��a�t<�Q�^ΆcOD���oL�5���1q+�h����P��dxj|����mX�;���K B��V��(���9�����7�<n0�#]���B;�R9p�&��c��D!�_V��uD���ӯ[o<���b��e����V�ʧ.�9���p�.��k�����ާ7yr�5Aqe�r�v�z�Rn݆V�hgW-S�p������?�g�.��/���镀�l��&%�u����f�.97�z�t($�y��`�~�=�_Q��z8� 3��`�JY:/����T��5I	�`����1����yx�#�z7�������Y=��}�rf�{Ozd�eMA���M/T�q�jw��g���9��n��/
j������Lz�WQ�t�v�}yf��������1��CɅt2����g�d��X���!_V����g��8j����.��hN?l��w�ݽU�Hen�'HgH�����'��3М���Wi�N���`
�r�u]z	����nO꽿{&А{Phe�g72�A��]e�k���3�׆ʲ� w9�S5���䑳љ�^�.#�+�wI���S�ΐ^�vZ�)�;qsġ�2�h��+��ED��c4�^�{�l�Iis{�4�̰�uq6��=���u*�͎y�.���I��e��g::܁f2g���l\���}��OM��������P��{�q���9x��6��,��y�I��۵��[�j��G.���X�s�D����INC�:��\��v}���3i"��	�u�ߝ�=㑉(���S}���r�@'��Iwm&m�f5�s�Q�\8&�h짘͋�������w�I�;J��X�[J^�-{�����b���:�1�iljT�s��	��Sԅ��mZ�qϯ��}�Lg�:�:��v{Ξ|���x���u�/�b�g�Ӥ��H�G��4�`��~�B�[������efe_{�f�������9�)���]Q��rx�2 j�0�LAn���W�#PѼ|�'��4"c�i�e�Q�ts^��ܶs�}Z4���ꑗ�v�\9�� 55����A�^�򭜑�&\�\x�=��s���<��F�}m�D�i�9������."z��m̒�|�Z#Ip���z��i���P��.z�w�8���eq���Q���)��'��:g�Oz��sl�J��Ω�BK�"����Htm����p��9Xj�SҗI����\����j=�=��,$�y�u*\��o9ђ{�IT=0��J�嗃�n�Mz7i����1�o��\<�S������o=�Wl{����`�q�� ������0�"������j�.7/��횿Z��l]t��%zw�톕on�!�~���~�8'�-�r�q8���2�eC��W#���	?�����S;f'��ϴ�����F�o�K�g[�>v�y�:��Ά���D�Il�!C�m�P���� R�֝w��m����T>u�<���
��X�\Y;�ֱe
��J� 2�p��$����6�ur��;���\mGY��NeΛL�l� ���{��f{��.����㵐��5,�x���L�a�k3�h���WW�3m��P�5ue-l���R�:}3�+ɫ��Φ�'��:��K�*�����N����4&W�&���������*O�t�FL�
��n�ǁ�]w�q��׌�Wyn�=}���z�<[�,sS���g��C�����o�A���4����Hg�WqN=�1�;���~�������;^F-,�f��w��
�=�L�on�?C���z;���Xr'b�<��U�ڳ�#~/�����}����zK5�%TA�p& �wF[+֮��ɍ(�؛��o�~�]4��t�{��s��u ��b�}�|;��.��T�I`Hn�U��Tݟf�u�X��_Cڰ��S�q7�iAs�+N>��n;:�d��3�dT�u����%J�[]�&}^�p6
G���E�4���t��3��0�mu��%g�Ѹ؜���<�C,��RFm�tA���;�=�3���djj�0�=��A��%�����uWT�r�t����`��)����fbf<�ӳ#��9���`�H]}�Om����`ѧ�6���?yi��\0J#x��r��c�A���v3:��L5`<��V>sE�=O����֑�fNB�f�+Pmܡt��&��(�+�)�uF��Nmo�{�oF@�Q4����3������tZɬR�(��G��]н��ȡ��gk|�m_d�2o�)@gz����)d�} �zG\�{>��+�U�ˇ���.���<�^^����i�UK���}WF�u�o����fhToz�S���>9>
⺳,�����0�O��t��B�{ۇ|z��q�\?|�]��=���{����v����dϯ��>�	}l�J����&���á�
rP�F�v��ѻ=��-\w�u5�awD��]����4�f|z���Vg���k�n���a�ޙ�ځ���O�࿍uq9��L�+�	�>��uֲ��걻�ɛ?��y����֌~��N���̳0�By.�5��Ӡ9`����-Rv�y�)�^�F]@��1+����^������H_ز�M��R�0�j�C������@7����P˅��41NȜ�q�V��:3��N��ަ9{�C��t���#n"�I:j$�5UC���#�{��b�t;�,�{�O˲������vDgH��ѝqܦy�R��~�|KgA'Ib���������%�M��@<z�nMJ�h��|�g�KJ`h�e�1�ͣ7�ъoq7\��`��;��^�o@��ea���;�X���"8PX��hp�����*ޗb��|,��A�DI�"��ya����C��7�s�X#��{�u�u"�d��1��W
=r�OF�T��1Lkr�,��X�	f�5���Up8�_f���r���˲�ͽ���)��M�=������f� �S3���n,�¢ԍ��٭����vp5-�̹��0_A�^2���٠�=�a�}�K���lwe����6tاwLk7YH$vnՅc;!ob�PaK�<�l�V��	L,e=�)t��nX���m��d�VY TM[�9� �Zk+,Ϊ,�Y}�!���8����ǁ��>�| j�Ϯ��F�P�`��\��F�u<�.��0�Jӑ�7p�!K!�n���I�SB���k.\�8m�)"�%̱Y���&���w?�Gp�a`�׊�}Z.�����b�=*��qV��B�P��2��b�����[y9�J����r"�L�wי���3��f�L��e��e��L�+�Ͱ�j�j<r4�u9��z������5��ܕbo��I��WSe�[xA�BT����FNn��oog��ѷ�h�`��u
O3{��oZu�(���ӢP�t�%U�+�Y�pb�M�ܭ�ocIJ���3V�Yi9�
�Ѝ���j}�/rˏ>���]�7� v�\mU�]�����V�a��,�M�ׂ���t����Y��
<d�|@�vlj�eЭS6I�b�V��RE�ޠ���Tԉb��s����S��YiF��Mg��h[�st��S]���,�F�B+��K�mRqG��ň�|��Z����Wx��6����̺�n�=�Vu,�u���BT�ั%R-�1�/k�z��,.#2�C׬ۤ���9��=��U��G��ļ���^Z�AT)�7e���\ز�C{ԡ�٪̝Zj�5ZX��N��uI�{;a&��:�*��O������X�%Q�Vo\�Q��Iu6CC:��� :j�G��(JS�K��>w�(V����%��U��f�W�����dF�kX�̮ÖF<i�N�=9���x;��w2[�X�����3oK�õn��J����&�ue�2>�꽖��U\ѓ��	�ZJ�i��=�1�[*�73h�ン��V�h�[Ԭ
�}R�vr�8
��7yh��V!fG��6(�H�d#dTEv�q�ly�w����L�ɖ�+�Id��]�fYF!�f��=�����)[����@u-����{�o͈���K��Ql<���y��G8��CuTGz�����ȹ�Woi�뙸��v����#�K��n݌pV�&����]]�mi<�4����,t�S��0��kP5̤�����d�Wm0g�9���������ޝu;�߷�u����(�������������h�"i���is1���
��*
R�

("hi��)��R�*�(���("��*I�j�&��)��Ɉ"L�$�# (������+%�(
#3"����1h�����	 ��h2
�)�&
(�(�"�*�h
�
,���������br2*�&����*���()�������
`��
����,����*�������
�)��Fb�
��"�&���0��*F��h(��H�"��J2�32��h"�	&i ���r��(���� ����!��2��ƨ��Jh"i���Ȫi(�$������̬j��bik �(���#�Q��7y�BO
����{g#�����dμ�����w�F��t@Ɣ�ʃi�pU]�+����*�g>|bc�%���eN�cQ�����C��S��v��^�}���8�>���b�y�}��6>�|7���3*-Ur�Q�U�A�!OP��q����BTOu��Оu�s��v㳮'8]��v��%_�\o��Z쥇��%P@�F@s ��@������Zz'���i�t����5���]9j1:�z�=��N�����2Y�D��12����^��P��=^#Q�u���z�ޒM�ZP���c�uĿG�d���Z�{�&���]C�0�!R���ʦ}��75�`������iOCG��q�ˎj���>�@��� 3��N�P��΀K�T�{�Tܙ�����q�ĵl�3���T��q�/M������/���}��������(�*z}v�mX����׳�.���:���O�Ix|2���_�v����[�0��z���K�v�^YV�ƀ�ީ�w�����,�'hza(������n���۴�nUxp�뗡�Hޔ�����H�|nL�B��/����x,^��@��6~]���x֭����]��[lY�W�T�xO�ȡ���������h�O���Lb���Ž��*�)N�ڃʷ�ʬ�J�y��v�jL��I�2d�U���Y��.0��R`W3v���@��	d1��}�&Pa�Uǔ�Z3p�B��g��Ap�چ���=�]r:I�;��pK��Urr��ua#��.2�R<��a�~5�C��Ua�R����#�G2��X��>�š���C��"�U����]F�|����п�䝣ġ�]�ra`��V�"j"�M���G�ǯ�h���g�;���|��=�u���q��瘼S�t_ײIܛq�'�x�~��sX�JP�:����ӑ.^t�N4�p>�{�wOq^��q��^F�A�(SRr,�c��s���}tgǢ�H*��
G�ԪB��ϟ�X�����F�t��A�^��#|�]�gs޶�����w�k�����ƒV`H)* ����j�:w���}xv`�
K�=&g�u��iMw��D.��m�!8n;��;�.Od@�Fa���u��Į+������V���^���N'�Ww����w!�h�o��F_�wlU��� 5#��h1�l҉Zb���^oG�cx_��\^�1��[gǧ�{���n;���z��Y$���KS�Q=zz��;cױ�x���u-���=�����/�"x��g�O1>>sl���ែ�ґ~U������4���06�¿.o�U�f�V��;'1k@�)��jo����V��{��<��������7쉻�W]�6�a*�ly�����ʝ,�u2&n��砮S�aw� 	3�X���G6<��C}��e��'�w�3���qיִ�ˏa�i�M{�6�*%N�q]+^*zR�#�r�����7�=y�X�~��(�`Wj�U����B�����Q����pOx�KYx=N{^e1���<�]Й��!&�9K�1\�;�T�nJ ���R}<J�釷��
�+�0ڹzyf��jR9Ooz.��`շ�z;W#�}C�ߺ�9��ɡ��R=y,��|��P�\��Q�;z=l�wQ����&ϑl������}���<�bqFv{D�V�����K�Gz���{�q�	O8����g�I�N���p*>��q�Œ���+���%�׈�a�L�}�(�O�orJ:��U��GI�}���"�Q�%��;�d�`u��'O���;�j�uA=ϕtH�yߧ6�:ߐ�^����J4)i���gK�T�#��2��f�?F�c��=ކ�hx.Vd�\��C�iލ�A �эk*Y��������FU1u2�ک�Oa���9��(K�s������ C��oX��g3��;���藔��If��J��Á?U��W�{lhY��*Ӳw=��.�l��K)u3�T�0���uc 0��gaM�+�^�!�Y�{�rMUs1ǚpS�Rz�����7Z[���vH;Y2dMSh^ö��i��,���/�r0uoK�9�����y��J�7f�WҊ�-�M��[K^�ri[������_Һ��t�s�����R2��x%��@���"��,���UH1fԸ�ڽ�|/g��{���c��>WD�ZG�\��Ӑ�F��툮�fm̂��P^[J�t�����'���1v�0;���FުA{�}m����3�zs	����r�	�Gl\u�kU�����N�_�(~�H�uZ��W�Y	jhK;���3���dm����ܬ����8w�cV��1ǔ�Z&�L\�1=˓�f_�'|b��u��M^*c����T��
#oW6=�.��	J]C��\OzO��n<�N@!�G�QR�����U}��w��/����^�����${����w:�6�����i�C3C��r|��U �=#����8�4���4�=ᇪ���zsJ���\?|�]�{�Qq��;ݗCaɟ_�<
7������s�����=>�"�He�����n��q�j���L{�]�K��Wq;�^i׊,߽8_~����ĕ���m_�KG�Ã��V�_?������W�}��q��weɡN.)x�-��e҇_t�|�[�w'��fmN�*9�,������:���I��;��r'���r��G)'GN(��3]�D��W2{�܂���ĲF[�{AY���z��b8���]��T\�G���76��o1h�c&���ﻬtVg��G�V������~�<��8s�N����L
�'h/�e=���|�+����r��&W�����.1eN��<JWa��ڇWU#qn�n}�����͝���������1��9�(=uZ®�sYR6�t����5�P�XD(�<g*�+�����U������.����vDgH��:��e�s�_���!΂NŅ�6W��u�;���B�@�}Q�S-�|�u<o�n�U���i�oH������b�x�k8�U2/�L{������p������!�<ܡ�����HM�u���'�m�<q{Ϭ�3De�.�{7��=�۽1�D���:Y$8%r�z���AOs�dڊ�g~S�"������U}�k��{�q8n���n��" 5Bt��][F�=���=�����N�ݜ�����0wػ���=ԉ�G�d�t�}Q.>s=2��;$L���������>v��oQU���w�����F_�ھ����8� 3��`�5�s:,̾/z3������h�e���wjE�,K����$v�[vvd5��uȺ�p�w���t��}�����<U0�!�,��x�<��n��S�g7N�G�����X�U���'x[wV�{��y���&��y]d�{�i��Q�z�y�Yu}})�9,P��8#�Q��%N�?e�������g(�ا��]���wto���7��7�����2R�ȡpz�3���}9���fg����
|Ԭ8.+�ݗ��z�%�Xac�tz=�� ��S���w�uU:���3�zx�P=1��X���ZN���c�r�Bu����SKK�֡lno�F�^��j����c*�-�2����Uw�Af�v�i�i��[l �v��[磍�G`n���dˬ�:����ua#��C�s"Ҟ'2��?�a�z��obyϮ&��ݹ]o{	��LK9Y
��t������H/.�B�NI۹�P˙~7)��ލ�[U3���c���>���mˁ��6g�;��\Je��}��u*�͎y�/��}��K���j��0�kU#Ĝ�chL��'��m���{�a�OW~�{��{���n�s�]�����z�"�:z5�i��<n/d��e �,_�*�����sX����G�����������^B������;��o�k8�E�IJ�$�z[S�WPz����|���a�C�"�7�����X,q�H尾�B�ŤYx�qۡ{`����%0V�T�8�Q����6����V¨3�uS^�۷z�����gc&�Q^�2�F��we�e���P���m�+���x-��e�vV���6��\(���	:��*�I�u|S�H�?i��;+��ޡ�o���7�}q��\�4ȁ��Á?�IqW;�J�Ѻ\xﯵ��z|������z �W#��F�}�R2��ئIr���@��xj�wfM�ˬ��^OX0<��#P�z��l'����i�9������2�%�����������m�^U�A��1;�®����F�|n�Q��j����y��3�'����ȯ%#�i
�ܾ�����G���31���*�s�h]t�5x����#�w+�1.}f�<�7VT� ε�e��w=�=z&.:!Ox�(2w�؞񊖲�z)�a��̦6һ��ܨ���o(.��Z��nu���M����.��oeH5<J�釷��
⺳¹zyW1<��{�������kl�g{w����U���e��Ý��Lo���1x�cߌ�����v�*�:��Mo^��J�����D�����\n=������;���9�;������.Ϥ��g�Ú�2F���������Nfhgm��>�u�6ju��g�yr���D�w<���p��]x�DG�g	��c��Εf�hЈ\6'�mR�-�e����vC(��m+K�]�O���A��H�^��<ʾ�X�Sb��O^�&v)oRt���y¤�L��p�;�U��Qym��J綠�/"�\��ꝼ�t��(�����k�wHT�o��:���i�G:׬A�����/ͥ��M����t��My�yܷ�I���.����\u�q�=���5p5�r��.�7'�)v��1x��M��R�,z�����#{n�/�i�����ܩ�H�e�^޽e#���L�u��]y������m�Ơʦ/�H�m�p�p�A��j7F3�֝e��{c����/�8=���gw[��/)K9�%Q�p'�ʡӹ������U��=�^/,�x��WpY�}�r��.��wѝ@==�d{{��t
%��@�����s��=3���HW,�R<�h4W��QǺ�(���!�;q��#/��fD���1�]R��%w�j �����A�/��Ќ�m����ُ��3�zp����ߑ�m_iɹ�ګư�)Z����H�Z���#����f���Y�G�R��~{���t���n�s���ZSk����/���
v�%��@���v�z%�u��Mb�9O[K<Ϙ���R�W�B���\6���;��ǀ�޹��v�H�/g�;�풻��Jl:�6~�G�[�������	@}��&hy���|���nZ��yr�\n����}��d�:�NȎ\�����k�f��7:�Lv�&[;E�D���J����$9��#(�E���]�o��T2Q����M�\ͧ'.���1�C��K�>��:�YyD{ln�������-6�e��s������<��y�� Ҟ%T���b���B�iϮ�!��t�謭�p�H=��N�@~P�^U�~&��n�h5K��N�;��/�{&}4rd�|�>��8�����v$x��x�gW��U=���/��ܵqއS]�=�)qy��'x>�U�u�\7r�j����
�88�}�g��8���4��9�X��/GC�}�G��E�lK��,�;ٵcwz��z�g�G�83�'�b|g|i����7Պ�y��Gm��w��#�Ӷu�q]R�a���bʝ7g�J����C��N������G�����Q��\�����F�����/��܎�1���hp�DK��5�#n�I:jJ�4�O�ϣ��ޡ3�
1�]�e#q�*������=]��gH���g\w)�W:ᾉyh8K��=ʜ"��Y5x7�.�IΙ��WS+������NhV�]��ޑ�������WZ��<A]f}5�[��.Ѿ�l5te�!J7(+�|e��=�h`���[G�>t���3<z���c.h�G*��ld.��oBj�EM�{R:V��Ծl~o-��w��<Y3{}��m=�Ȓ�ˢؾu<��^r�i�*�b�}�K�̕slc�S��Z�Y˦��7
w}�LQ$m�qs�S����3d�4]n,�+����mz�V���u]pG9g\N];�a�ʀ%d����W)��FXW��CU��6��L�a=�ޱǽ��q�n����]}q7�f���:LOҺ�������W�a�UG����f�9R��ox���O{��2o��@��u���g�U�!�gd��e�@�hl���&=���q��څ�4�F\6����@�5��'�c�`�NgF��+pz��к�d�����skIL���xT%�q����Ѹ����6���&E�,��\g�L]t�~��k9���L"澃�Cn�u+	ǵ���=7�W���ޘ�|����w��ۼW����퀪׋����7��g��O�za�����T��֓���=˼+s����<yu᚜Ѫ�J�=�ѫ�'/>�V's�C�T��d��fT	�0�+��lӬ��!��U�ڗ/Pյ�m�0�]`<�r�y��G�oe!y~��<N`0�S�}����Ʈ*���G�O���}��Q�Ƭ��]O�Nu�o)|�F��8O��#�/���U@_�9C��x&>e	@۾����`��L�^9d��7_$Ds���w��=._;����_!��ع�o��w���fQ�sh�P�d9Qf�
���v�*�NN���t\X�Ag_u���i�\���f󒓳�T�ތHfɼ�m)����0����@�%ͣ�&�DkږGC�N�eL���$	zs�h4��V���cz�K��P>:݆],r�
��S��y���ۏS��9�j���j��a}�#��W`WpN�V�GnU��Ma'�ruCƲ�Z� �����hb�`�V�q�M�-lV �s���d�A\���ڛu��I�o�v����E��}�+��V��`�>x��	=�N��	�"�l�aM؞��T^�9��xUY�Q��̽h����"y�b��sQLR�`����WWΓ��n#0S�v��g�+QU����^��bAU ����f]KWv����s	�#�a���+md�׹��f�:�*�ꮜ�u�*�nNh0�����wO}��l� w��n�����0�2>u'��`m�ۥ]��K�Qg�����q[)�'j��CDKu<U��릲�&�\�-b�ؾ�x�sv�:�̹�^Z(V�ʱH����L������^[�w\�+B��/���o6��db��I˾��S��ACx�ܶ���aC�U0.��ⶸfe�2���b٥�:
�����,e�3t�I����֎��tq�g������]cJ�u�3`ti�q̸j8��@�5V�i�,xޝ���]}8���h���aU�U\�sT�)6�z���^n����ۛ̌����%9�����iuA<CeP������VN�Q����'F;R/1C][WHn��ycYhc"�GVU�2�+��ܒ�6ޘ+��R�+i���U�;ǒ�y;�cj���5���\[B�Ɍ��aT�6Vn�hu<`r4g/�7���F��y���w�GIQ'yJ�Oo�lvk��MH�q�yA%���+����"�;��)�����ލ<JN����vud����Me�EJ����UN��5kU��U�]��s�Vj�
Yvݮh`ꪌ�!�ʺ���vڷ4s��S�a�-��ʐݓ����� *QZ�EEz��v|��VKs�B�W*��9ppY=�\�3E�v(0kUH���M��}�r��M��ɃYYQ[�+��Z�zE�%�Q��|]�*�V
Go��ȣ�i�pК�`7�՘��Pz��l��Ժ�+ġ����j�׵�g�M:��b��F��T���ũ]���w^�M��N�VI�I�,6i�}��s����Hv.r���V�٢LF��'���l���G*Z�}g8X�G� �}�'2ߵ��-�6/�qJ3�_H�$c�~�Wֳv(U��\0�+�|�ی�ݱ̋���)kx���8Nn��<8D�.(9�z�,����] *Kzt\�姓�73E� ���3�(&bh*�"�Ĥ�h)j��""�Z
"*,��+0r"*�����*�	������$���b
()�
B�3����"$����0�
�"���������J����$��2��*
br�$)��1���1
,*���)���)���r��A��&((� "� ��JZ�B��00����#%�����)hhh))�!)hj���32(r���"f�(JH�� ʚbi�)���k!2i)"���J
2 ��H )((J����JZZs1s3%�B��2+1��"�����(&2hʚ��1��3	��2�
r(���2 (���20�L'3
ZC"�����`�����&���$))�31�������7�&���Ҷ�۵���Q������y�`ф@�bi�U���+D�i�V�:Ӿ%v$��-=�8�N�/	�>w�� �iή��?�d�y��9�϶g�<<N�/�nw�;��u���G<���W��kBEff�\΋�ؿF�U]R|;��$�����EL򘸍�B\�F>��z�t�/�wOqGi��m��,ׂB���;^f�Xg���h�A�X���R�].|���_���h���͕Wۗ�R���T��~�7�qۈ�w���P.K,i%a��)(���֮��՘�����~�#�w�b�D����򹕟oPý����u��x\�5��Á0[�&�D�X�{4�r�1(�w⽢cQ�{Q=��/!��\���J�ꑗ�]��.qRs|I;-�U��J=���~��)�&/4LcO��8ޞ��e`7�׀\�{��o��;��N+�ʢ���f̭�%���>����HUԽ83�e�z�F�&���<���g�OL{6as1�=�F�g=�ΫG{ �d��\��c�^�xО+Ƴ=:�dr��]тFm�.|�{3r�d�f�yJ����ƞ�$�Y;0� Ox�D���Y��ϛ�\�g�_��_H�h�
�Ö&�%��C��[gH&��ۃ�[������r��u](�ˮގ<����ma#��]�o�w�iRF:��{��j�{9:�D�D9�i,Εe�6��QK�؉��^]E]M��㊂��cq%�J�q�ȷ�̸	w�:�������!b*�������uOq�j�`�q�RF������
�0���5�h���UOM���lV���t5|4^���'3�|�C3�{�Ý����#ג��������۪��&�_0�о��Emv��S�NDb��~�W��:��'�B���G;�����؇s�>8`ۙ�o�����Om�u�'zg<h���U���{�F��.�:�P�i��z�3��I����#��������~��G��L�rp�</�&t+��8,ӡ�p�X]�)���چ����G��5J���Ѩ����6���^3�*t�Y�R��3����F��t~�3C���f���k��6�����stgGSﻫ��}�Hr�^F.ʖo�:I���>5U1EL�{�h�e-fe�����Ϳ���Y����X�ވ�����gD�ΐwR	^����L�%T��@��7����t&����]�Q���֮�񿝽�����H�;�Π���U#.;��w��kKU��U�lyUr�� U�I�'᪐7 �U��E>Ws�i>���w��G�d���g�hUu��X��p�N��P��4[�T�D�dw���|/.�׽�7w�S������xvb �Z�f8���;.�fQS�N��'"�[ �������X��ɵ�;R�B�8k���	K&�s�2dޒ[f�{jwb���ۃ�����/f�w���U����L�<3�fX���Q2��A�/�@�S�H/K�lǠ����ɹ,���s�ޛ�d�*��DS��"�̖iT����"d�SB����<�VF�D�"�':�d.W�Ŏ)��|z|�~�Q��D�2�퉘]bw�*%�u�-d�;��/z�Qt<����jy��_r�����t�ކeX߮ ]r�:�=���a�Z��w�&�6�hg���Q�9W�zny|;��:��}\L�^�\���w;��gV]v:Źm�s����u�r�i�*5K�q�\?C}w��=������ב}��F��<���D��+L}�yL���p�Oc'��W�WOI��ݗ��-\s�=�tN��۬b�Y��v=�Y�ɾ�Ώ�y�Ѷg��G�N\L��P2p9>�� ү��0+��/G���5�37y���*P��@��W�������ma�|N`5������xe�N��z��)*6te�	N��<��p��{�����Hn��J�L�Vx���U�/�+]{��t~�̊�j@���wM� ��$:�N_���D����Ix�ʹM�6�V�x��/���]�׫�A�hz^��ٗ"�.xy��5e�2�XO����`(a=9 vq�>�\g�;vS9���&��7�΄���]2�P��H!}�L�/�]�	N����Z�9{MP��3�ȼr��z�ު��w��h[YR6��I:L[�uUN@3l��wG��Tu�Q��q�=Y�n�����}�t�/3�;�g���/-�i��7]��Ww����I���'{��J���熯]K7�V+[�ÜG���3�ج��;�9����{^���[�5��} �,� jό�!�7({�WO����	���C������\Q��䭫�IU_f�dx�|�'.��qD���A�:Aod�)�FXW�m��x��=dye<����gX�һ���{m�ϟV�7��������fK4���&.WV�_��oל�Ss9�Q�X���u�^#|��t���|7�wV�w��i��ʸCg��N譙j�'�y[� ����S9Y��4�F[j�������\ ��5�W��J��$���+�{��4:�a���
��'���Gإ鴻n;�����_F�u���������e^܍���s�o��G���SP},m�����O�WQ�OM���ú��I������h�袞kj[�@�l'�2�p���9�H��Rg��6��r�
��YH(�|$b���VUNz�-��WX� �+�i��q�}"�U�.����^K�ˌb��E�|z�qJ�b�����(m�\UU�����y9^j�'��ܮ�u�i��3D;��Tz=��N�.��z{��F�%P��V2�;��ÁS�'67i��~����./�w�Ut,���:3����z��yʬN�~.͚�[�<dew���x���?o�h;��1W¹ۅS����}�W���`)�k����Gѽ���e��z��9�a���'8��g;��<��+*���įF`
�cVE��}�s��yO�|���h^)�:y�qU�F�h�GW�ɡ��3���T��p9�'�'��&��Ƿ����V�fE%��T�w��my�WhＧ$�w�Iڙ����S<�.6�	sc��z��u/v����5u�(���~��,>�ӽ��\$:m7�Yq{$�,	�b��T��OK�nhVg<����b��>�+��{9�p�tgPgm��fo�r%��t��`@H����3�ۀ��;�K۽=>W��[g��;�1B�%w^|�+�Y�0���HN��_�ƙ5Q�p%,���{"���51{=d�|O2��F������n'�yA~�G_N%vuH��b�̟,�=?d��"�����Sɿ�Pͭ6wߠ�����y|=ޮqLm�#:�cM�"��h�+�����KE>�D�O,羅��
�j�}9�w:�)Lѥ��6�k�C�>b �5�u� �����Bj���1�m�i����-���.���lY���&Ɉv�� �$~Ki�`�����h�Bc�H�ǧ�{���{���주<}:��S����=�'EmI�7d��'����zpg�L�7P���u���Ofd3�-6���g׳��]h��5�)M�"�˝�30���
�;ƅ�J�W�*zo�]R9.��U/<	�]G3ٸ9Jn�w���h�wO@��5���%N���lOx�k+�"��Hw9�u�=>�ݓ���ݗx�}wA�H���9л�,\oeH5�Ī�{p'0VXk�h�׷�5~z��<��ڭ��u�~N���>��}�A�N�mX�W�돲Y9�s;����G�z�ڑ�ax��2��z�7��8}�_�m���uU�O�up\�#��N�gg�d����'x`6\ʻY+��L����p��2�j ����8p�ģq�p+˝�{�SO��s����vf�\Q����G�T��4�Y��w�3�g�oי-\EOQ�%��;�,��B1W��^��
����A�?C��U��{�~��:v����=_:X�y��tu��zU��[Ҥ'�^K�oh�F���ф�n��Ps�� �դ���MNC:M�hkBgh��}x�L�l0|�g!-��"�N4�/G�ʲ�\�暐WN����S�k7��I安{���/qc�Ѡ�!���-0�bW�Q��6%�תq�nn�ɯ�v���1�"�㥏.��+�t�/|]y�k*Y�����0�����M9��^�+ӫ���.��m�p����5���gA�>q�@=��c��%� ��YcI(k	~��B�j�_D��n����{�j�v��u�:�G9���QتF\w]��-�/q�g��)Ү�}��)�(	���U���򸛞�H� ���>}#��LY;�̚�;Z�g;1��/�j����,�Jɐ:Cu�����B2Ѹz���ف<�4����]��^-UWه�Na6��'.��2YRHk�%r�����S�����(�y\�:.ǖxcWY�#;_�ܬ����%��G�:s�rsD�.���W������* ]h7}!���՜��]�HuƷr8\Gr��k�q=�<w�f��T>��(�w K����Q��w�t�9E��W�<db>��e�i��/���]�y�U���4�����:��J�
�P�s˕!�}�������R�<r2���r5K�{o���]���z��7�;��������;sJ<����*���W��&�Ң��V�ީ�E�y��� ���j�q�N��S�$VQ"�JG�å���F��a.q���{���U;�!n�O,����޽E���<^&ޱ�Bvjp���W�W�<���q��F��@�uXk�̛|)�RJ������L��g�Dx��Nq^�p�����n��q�j㜙�1=�Ϲ�U��Ǵj��C�;ڮ�w������#�'	��<|����ү���LѮ2�H�9��J����6�w�y�b;��i�O̭�p��^[y����^�½k�g�Pv^^�|����ld�:<��"�r�p9�]�{���>��C�t�% a�ꮝ�^޽����CP�B�L��n���5C���/��޹c���7�K��צF���
��U��VV���ޒN�/MA�P��3���,����?i��>Α��uGv�������\R�̛w�x%5~�	���Y/��Z	:�.U��ѥ�*����t�\G7}���8�>ڏx�0Uȕ�2�΋[<4�|��-�Mg���,����,	
P47(z���=҄�Sq��l���kM�*��|�RY�xvvu�9�#�vu���u�0�.K4����2L���+�����?*5ӽ�犊~غ�C���=�7>}[��g\N����m�,�"T'I�DG�}r�~!������N��)�ܸ�������o�����?6r%��*�w8hV%��m�����vA�ݺD�|��N�6�����x2Y�P�W�s��;�)��itZ��O>�]����7�����w��︁ǜ��f�i�ȕ;���t}GY����`���=ԉ�q�M�wV����g�k��������=�S�j����B���D��u����\SBc�����}ԁ�}Ƹ��f�
���/���o��n��U�H4k�> ���O�D��u/�Q�R��%�q����7%�4OF�Fy����mc�54�|���2/K����*h�Xہ���+�{|/ѻOKU���f�&cL�̇��:P�����)Ѹ�v��,�i�3㣉[�\�⧰�n��,<���϶��g�`}wx8y����ޠ�}ژY/���fV�����+�^�������.zo$(���t�����5|=��A���.����G��He\ȿB�'3�[|.���
k�[Ь��Ρ�z���L��5�
XՐ���Iqu�}� �z�舨;f����z~��.�|_�z��K �[)��7r�1��[���M��y�CgSv�[�ya��y�$�`�E.�w<��)�:.j$�K���KG�K�*�<��Lv&���r�x
͍ٙ�Z�͚�Z7$�}�>�ݗS���J�]��t��6�pf������l�꜍a����d��KL;�f�"-wx`�GJ�S�U���MW$�b�@�7�>B���2q���@ ��5�"�@�(���̐h��ՙ[�y�,�0C����R/��#�Jez:��/D^F�Xe���і�ȱ%J[u��g�	���̹���{W�[���^n��Ѯ:��}�A��|�;}k�c��PΒP,"D�	=�g���y��/�.��LЯ����-����eg��0�d�>;���rx� j،ܑS�׃�n<�{�:&z���u������q'�Z
 �W#���Ѥ�vuHΪ�*6,�~�k>�]qӳ+c5U�\� g���s�����j6�
�����>=>��Gz|^��h�ޞ��z�?V��{ *m��I��T��l�?K�HU�T�83Ѧ_z�F����׌��{�j��y�g�*|��3^��$*.vs�3�*�s�h]t�5q��qY�j�{,���{{0���t�я��Ŷ����3���z*6{�I�E��=0����TKYx��^���8��\^�<w{�k�pۄ��p�}wB�u��� ��P���R'b�,��������z{ �z*�.�����Zydj�7*��u\�>��\G��9��vՃ�nZu����k���y���5}2�5Aw��b�&�e����vK�[��,��m:���oPlp �f��kSH�iP^6wt<�=׈K��d֖a�:t[���*�T��7Z�X-�{�U�{[�n#$���\2vG:-M��Q�5���zep�e��\�"�����6�=�e{���t}�1wW�i@�є����WHc��o7&k�&:Gwr�3�4b�CO1喊rg9���!��nNH�7ڨ�.�e[�����X�#%E���^��f.[#�W;�Y�t)j���և���4�-��[���(���L���P�(R�mC�1�6l�����T5��ܨ�Nץ�쭰u�Lm�n���*�1V�d�)m�l��4Dq����4sW���r��oYU���L���(�����<�qE*t�SI��Tz�mm�'�f��t��-Bl0WXU�c�Hh�¦��{�g�ݹ��(1L,���u�K�:ZV���s�ww��y��-��EXICc$��`���B-��u͗a�v�WZ� ��v&iް�J��N]���Q�L��N�d�D��lOk�8�Z�E�u��#�U�.�*�)�ܳr<�U�w�[��w*�^�b%<QJ{׸i�NƦ끱�νYm-��	޲��m�:�L�b���4e�宝��k><�0gnRo�	c��u�	�o�tdY���a\��-����f�;��A&d�7�n^���Rv��2�r�b-.���`�Pٷϩd���o���˥W!��аo;�3s��}�*��k��ݴ�����6���]Ѩ�P�煴j	v�c��t ��"*(^���ҵ�M$-�7FM��V�4B�;�.�#t7]��gt���|�+�3���98f�<��z���ڈ�D%�8��ބ--afF�l`�ɒ��+5���֔��ޮŧ�st�w�VS�9u]i	/�^��S�i�L{v��ݴ[�Lnі���r�smr\�V�E����KZ�ۭ�����8`�hs�Zį"�i��7v��pU�5��KE�WVL;�Sm�3K\���ѕµ%�&f�w�UI�z-U��Z�,y�V�r;�D�vҨ�B���۲���v�|�qP�ug�z���"�#v�欑����Ȳa����Y�HT,�M��u�ZU���s���[Č��*X#p�+��|���-�8���Ou�4�J��w �V���ĥ�W\���O{�����x
஋�Q��wٳ�#P^����X3�;t�Dof���ݸ�Nܸ��D&�^�� Uo��ݜ"�6s�ط�O����raG��ܟA�&���3)�6�l�M�� �:��.{�X�'���D�hL�R�n�I2*t��j�ԵN�!r�E�K�2h��a���e3v�N��2p��x�����##s~4��f9}J���K�!��kٖ��$�xw������/Wd<K�YB�iF�{۝I�3�A f?Ow�?{ٞ��=d
JiB��0r2��0©� �Ji��3�h�h�"����i"L�"�
�����
+3�2��0���
bih�i(��(*���B���r�0�$�3
K,S$���B��,"��3$����(i���V3&&�������R�r �2��2��(Jj��h��J�J����2����L$)�$�ʐɢ���$2r20J0�������)H�B�,�L����ih�2�$��
(J�2�����2ȥrC*JF��(�!J���i�H�bZ�
rJL�� �����i�H�h��)rS 2�Ƃ�L� *�)ZJF���������2ri��V���(j������Q����2�I����������;�����YDM�\t*���Mǂ�(�{�e���Z���E��(�%!ol,xB�v�jJ�E�v�eڛ]���m=�6��ﻗ�?�ô���LY�n~`0�}���\���}����G;����^DTX�Z���r����g�XA1�/�w�kM��ģ�p*<�\w�����殈��Lo��
���>HbSէ{5\%�L�+��J����Ix[	h��_�����;2�W{�@lT	�֏��܌��]�ԙ`��g}���^3�*t��Rߌ��gKS<�ͯt���FaE�7�.�{��3A�F�c��<�}]�{�����ב�k*Y�:I�3�Tu���'w?U�MW���x�X�H�m�!\��j#Ou��tOq�Fu ����%�t&=%�xG?˹�-l-��iޥ�I��1�uB�2��Z�����ۊ�n��]#�ﳨ��H�Ze��T�|%�N=~��d�Dl�5�I`L�|
Goz�4}O���D�ZD3|Vuo�v�����!�F�Os�u�˧V�ۙ� iY2Hn��C�FZ7U ��q�q���|Q1�%h�j�������rNa7�w\N_��|d_�d�J���d�DI\��ӝ㏫����fz=���{d0B�9�a&����|n\ѧ�\�J[����՘�U+wCL��#m�D՛��w����ȍ����xv��gD�r�U���+��_v��+�*Z����i���W��s��/�A����}9�2�瘴M���cɣNױ(�*y�����毃�=����-G�@�����e�ہ3���1]�cn	�7
{��yzz��y5f��Ԏ�]�\������7��B���6T�b���Sg�����[[���}E3�qˇ�.�pQ����<�����y�"�ͣ�}v*n�iϱ��b��  O�a\��7��HJg=��g�?{o���£�@u(^WNs��>�̉ۮ>��w�n���/&}q���G��X���+��.��t���|n7-\v騙� �pD�U��l��c�1��u���'o�߯4�f|o�x���3������iW�s��vw5�D�R���s�ˆ9�>�:�GS������T�E��fa���,c�t�����퓹otq�ק�m ��+��'hp��{�κ�+��Hn�we!F,��qx��Ǟ����'w���.���A���s:sm����d^9}ӽr�k�����_�}SN����|7s����}s��jN�*��(�#q�.�x��?F����Α��θ�SQT�
��֮(���><-
��z�n�"���}�f#�1��3�u�RfwK!8j���J���+y@������{VF=�:6��W̘u�We��w0�n�2arh`�;J�����R�<f��x:�S�p��k�;ӏ(%"9��'	����T�qxv�33}[��J�sԆ��z�s���2���*�qS-�\m�J7
�X��n�I��ݻN���od�������ۇ����x�p@�FX��nP���ǽX�����9���=�O��]zs�OJ�ၿu=.7�aێθ���a��|������{$s@�<����u3�<�G�g_����eq��==����m���t�����q]}q7�f���/���?B��mʝS�~�¶h:;��T7p�x��;cǺ�=�3�ɾ���%��[qӵ98!�b�=�73�fG���&%�uO�3ni��MWIP�����p9v�f:Z���d�v�n&��Ns�R��Ng��Fǥ�`��|r�◦�.ێ�uTDU~w�{�%ز���d��%@o{�j��g�dҘeMA����ä�>V=��ݧ�^}se�۞���Q��R�t>��zc�z+��vK�;}זoOa�Jߠza��e`wS�pa�uՆtʨÏ��s^���a7�,>�˼=�r�{�At��hN\y�%t���<Nd���?�/߽#�Ĉ7��e��Fk�Fu!����y���"���F�dY�ݹMz'Ͻ����~�=�Z���"��&�+�i�gGk��C��a�'�K
�)�aA���:Α�G��Z�rAg�.��ͮ�Y�c+��r�^���{(��q�Ǉ�ΧB�"n��+���[]�K��)�{�����S�ޔ�Մ���Ű��*	����?M�曕���&���g�[0�U�����i�)cVE�*�}�s��yK�:79�.��fD���ўv���!��X�Ϣ�xdK��Ek���|el^����ٞ�������r���*���.W�Fz���n<�G��V�fwОy��S�t\^�']%��	h��i~�R�y��3Ɏ�����ѭ��Ѭ,����gP����{��[���.���Y�$�,	�b�U!S�X�Bq^���2w����kzvz��U���z:X���w�s^��h��i'�������N�������C�#��[S�WPzݿh�K}x=��ef�;vR��������s��HR/7�چޞ��`�@肕"l�������Or���r;��F�}�R1e�(��.ڨ��ܼ�l�v��L�5�����Z�/O{��4m�i��G��i�{#Ƣ{�ob������{:1ϫ�=��x�.��o�2K�KSgd��_Ru/N��e�Tl{-��C�O͏G����[�3�.��w�sV��%�m��n���aW^L��1)O7���n�]ގ9ԁ����2��T�/J������9E��N���ٹ�ԯ�p�W����+�s��R#�s6vMF-N�y�����1��j��$�ߥ �.t{�_����Oy��m�;9f\@U�Q.w���V"���@�B����ƹW$m�����wF.>�G����z+��jd�@����0���6�o��s'm��o���WOa�̤6�J�7�tt��]���ފީ�x�����NO�<h��X��¹V.��}st��W=��}���ܿ_'U��P�7�v{�h^����yJ���%RzC���r���7�̨w��D����إ��ھ�U]��W�s�s�fL̾�SY�3la�%d�D�}��b�Ϥ�O��������V�%q(�L�\�;}w�w�$�������s��t�zβ���w_~��Vi`��9>K���tk�8."���3��ܪ�w�`��S���<�0� �@�J�,;������C��c�t��x��b��c�W�-N>�9Sۆ�����X]x���+A��}����:��>���Hv����ŵ�,ݝ$�h� �V���^���ފ��g����齻����b���x=��sѝ@=�}lv�D�Rq�y]ݾ}�}>���n�j�2�>A�������b��x��QrѴ�Z9,�X������=�������ĸ��i�u�H�o9ִ6�;d�\;_}5����u p::OJ��T,v�kUe�B���B3��`z��������-��Z24�����
�'z �(�J��(�eR���b����ﰮ#����66��P$ٝWo��i�]#{���� j���@�v���G��\M�u�A�-�������j�3���ת��sO.��^uH��U�,�Y�PF�H΃�⇽�Eţτ�q���S�
�z��`N��gJ��1����p��q���]w�EÙ,�h�t�H��L=�V�)��L��b^��Ui�>:�z���M_=�Y��=>d�}ƣ�)ۨ��e��0��kf&��ߍ
y���ȹn5FtɎ�y[F觓W��\kw#��+��q=�<s>��sy���vM�~��W7=��u�=�2;�^�=��9G��{*�.��ﻝ]� u>�(��8�m�IO"�G���ٗ �l�*���#��WVa�/Oi_%/O��P��'���9"b�#���5��#��ѹt��v������Q���ᓁ�z�e�����ѻ/�ʋ~�~$lw���g�tVB���ˡ�L�1��R��9]����y���3�W�~�CF��ͮ��g΅u��m�jL%so*hw�OګF�~k��y���G��L�1]�8Ӻ�.���̬�^6(����E�N��^c3qa%�.H�8C�ڻ��tt⪚H΅78�]�)I_g*�ަ&|�P��pG�6�(��z��C�̹�;dE4L��
�o�����=���Ω��zV#w�܊x�j�[��2��۷]>�d���2e�c\,�Y5��u ׆S���E����r:븯u���҂ŕ:ow9���23��bU�d��0�h�Tu�J��m��{���r��z��v���ݖ�Z��Y9뮺K��z�GD{r�+��N��O2
�~�<���.���CZz��:G����0��_����B�OFn����h?�[:	;�,	��S-�_�uR��4)M��q%��<|ǡB���,�v{��^�}�!����\=�t�q�. ��X�hnP��wZ����y�&q^򼕴z��S�bn%���w����#�g\NOU3E�f�P@�F@�q}1��B����ߣ��W$w��s�#<�>��Os�<{�ln>��o�θ�3���̖T^���of��f}�zt���� M�l�>��i�0�Ͳ<5r�8�R'�:|7�ՀxM:RcWmh��}u��L�O\���}�G3gd����7E��ͨ\^�1�	��7��= i�>����75�.w�9�����o��,4pcʸ��^��8Fi��_�iྫྷ��AAh�eϚ�KD+�k�
Oy+Ӻ�˷Q�wk��S��7*���$��]Hf��u�y�$���o��4Mt�� 'R��/��Y('�sg��]�9������� \�������y-◿TyXk��8׿fg/i�����R�e_��'����s��r��7�@oz!����g�d��a�4},lq��R��Ƿ��7s	���tmW�>�'V��=�yp��}w��OQ}��N�W��i�3㣉Z=0��������� :<=>�e�WPֆ9�C�ۦN���.�pN{nt�sݳBr��-_�P?1�7�>��;��Я󭬋�N�|'�0�+Դ٥Xz!m�}��|=��A���.��s�	�Jgϱ�^�.q_ej٣�7�x��3ƊU��Xo�R���4��.u>�=S�#�s��F�{����^����s����ܶ1Iݹ�JL�3�
���F�ۗ��F��xz��s�@)�Ä�3��}^KYX{�R����U��<�✓���w&P�3��T�)��t%Ϊ���:
�=ޜ�y��~/�`R������}=�z:�� ��ߙXe���іE�n��7��mRՃ�ܽ���fz�V�t���������C�r·���k�c����$���0���S�H'�
�MR���p.��S��w�eƺ�5�|���������& U>�Ŵ�\�����C:��.���zVݺQ2]���	�҇vg^W+��<SrG��i��qw,��ż8,���vNS���B��aoS�c��p�%gw�Ӟ�[�՚E���R�l�G���E��<�ފ-��]��u��;q�HN�F�����c='�.w�;��qg��1Q�p$�&���{�#P��ʢTOr���W#��G1vD�d�z�k�NN�5="�.�E^̗5� �� �u��zz��h�Bc6�l�� ����W��.��ꮼ9���Vp�� =7�q̒�*���� ��*K����/�1����#��P�olf'w�غ���t�'��|O&k�S�d��W.vl���
�*\��{Ū�ʣ΍��d��s���1��z��u�r���Q����oy��E}��2MB,��釳�������xn�.�j�s&:"^m��l�5q�LjU^l7�t/�y�:���7�ފ��}Gg��{~��y���o	�0�a���0�/Oj�U��q�~�	�����q��uXs�W�}?(�`VK�������+�H�����@>���P�\����R��{m_:��&=y@ӫ���Ua��h��ݜژ�ﳳ�/�w>����p�vG73�`Ԯ%dˁ��r3���s]�dlT�{�&p&-�{>�Y����ҙ�bp��X�k�hU����;�AtR�2�X��:�ޥ����j�s��MA|���#�S�����"M�M�[\�u��o�N�I���Ʃ]�T�tT��ٽSFP'.f�i���z6:ׇ�%>u��>��j�f�>������S�Q��ߦq�e��Uw�p��/a-��]|=|:q�b>���(X�����`+����e��wM�t�3W��o�p�<JVe�v�,h5�cs�AJ�
���J;�Y��3�o�C��dsXz�q�:��D>���]!������YR�l�w}s��m�����ջ�|�8v�y��g�ک�O~~~�ѧ��{:'��Π��;
�h;w�ȬSV��3��/���:Itf	�<��cn"��6���\�}��B��u ��M	���tZ�`n�c�q��z�[ S�X�n�T���z�4}O���e���P�:��F��m����#�:;:�e��l͹�Y���W� t���|P�hV���l�Ow��TW{�7���ف׵̿�Na=�Q>���!��K5
���ᬇ���S��ʱ��^�n��	��&?<�G=O�Q���c�{��#��Z�Q���M}�Q�����I"�^u-Ό�n��ts�-d��u�\�.��������k��7_"+�J ���* ����"����P@DW�("����P@DW��_�PE�@�� ��\PE{T_���U DW��"��@�� ���"�"��b��L����@l� � ���{ϻ ��� �Ǘ��%%(���i�62��� �h�Z�E
(&�i�*� ��E���[#[YI3Ѹ��kjՆ�R�3+Mh5�km���UZ�S"� n�Q����u6�f���ef��Mh­�(����6���Ym���mZ�O 3����eu00;��wcK��Tn���p�0(����%��f�C�6�[�Y�]w`�x u�  ��   ou�  � �a-*�5i���dB���k�d�<��s��3(:�0�̐V�
�Y�U��i�@�D��֚�mY�KE� ���oqLL�@���'F���n�eԍk����e�ۆ�R�e.���He�KY6F�<�h=�m���֋�uͫf���4R���G�n��۸2�Y�V
k�u�sTh�Emۺ�R��0h����=K�u����i�;�mkNm�m��w[)l]��U�an���g+�+S7v��uk���E�im[m���A� ��[�����U�5w+�n�]�\�ƌ��mm�7w,�v�ҚWW�ݍ�lWf�ڷ-Ŷ�3��lkm�-�Rڼ  �޻�gj�4�����TѪ��j0f(�p�)N���C�m�2���k`^ s����4�vt.��ws@�WX�&֔]ۂF�p$�`��]i��a�����݋�\��$���k���Y evuԕjM �M�^      �4�JEP ɠ  �@ S�R��z� �     "���IR�i20�## �M4�4L5O��J	�F#&&�#ML 9�&L�0�&&��!�0# �$H�	�'���G���h�F�O�������>�>�?Gݷ[u�Y�7[��{c8��E<�?��a����a�Xp@�~�Q@���dh@�R�����H�6�3��?��;C� �!I��M�D	0���=�4��RҢ(��'�������`�����~?���D7���A��փ_�Q���?n��8�}��1*��D���}�<���M]c�Œ��n�G�Fc���*;W��������Z�jޛ��ݿ��L����4�L>�lP�	�ޕ�䩌d�[	�$QB�6�����ٰ(�m���4�S,�z��n��"�1�&k)e�����B���I��]��{���e%��ڸ�6�wXRj�Â��˓�Y�X1��c��\��YL�Z%��( Co&��v�'I˰�p,�q�ЍPm�h�ֵh�4ss%eӴi��&��B��/n*s#n��5T*�`�2��'V��	�l���d(F"f�]V�FV�h]�U���d��\���&��M�woX�fK ;��U2�͙)�Cx2�(����L��ǎa��	�5��(�嬍B��sA.ĕ%jl��e��ǖ/OҶ�f�7�m�J�Kѡ��BJ�EN�#:De���)�2j��sn�٦okK��"��0�z�,UH�Q�[��Y�[d'��
R��r�3h|+ ��coC�m�G�2��̓B[s�<ɨ��W���tJ�[:r7,�E]^Y�z���ޡ��܊��۳aH;�cN�T�L�Tf�n�f��d$i�ef�
kf��.��h���T����j*�/1��ʋ�W��C��ɘV<��)��)�����F�4u�����$f��wR�Q1'R4FO���,RUo^Z�sh
���=��XZr4�Ɯ�ߵ�5�G����4[8L)�+�(�X�^�W��X�o�V7)���l.ŋ��HS��`�;��J��#�bc4GZ\�2�Em��Z�5BR�n0��&ْűTko1�d�,f9�����*ںlI��	${S
�z�\��{���d���3B�����B*4��0E[��m����j+�:Y`�1$�j�G�BH�b�]�Ҧ��V�����$
���1��ST.
��"Õa+P�4��I6JHm�UAd�vj�H��5dbq��85��31�	�B�R�.\��I��,���Nf�4��*���m�ۖ�i7�h!me[Hd�H7�=��$���\�f�K�t��]��C4,×*򮜠��
�/Ps(���&��.Fm��;�~��b����Q��ҋX˼T��R'3r�]��ѕ����a��{��%�#�`�U���x�w���v�Ğ�y4I�vr���f�y�Kuz��p��1�v�3E����T$A����N=�[lQ���u��۵�ڷ6�V�Wr�]���
�1 �;�
�82�7�d���9c,����YBɛ4�YE:�����طl���A�������t���)٭y�J�unl6ڔX�4�=ʬ���}�+���E�tX̍h���v��V���+��hV^^�\�[.�N�r�4bݔ"���,8)���w+`ېK� F춲�Sc��XZI�l0E���j�<d�*�E)me�*���,��)��>B��;����["��2�K4V2���RY�C��2a��^;�Z�,^�1]��K&�����}n��B�b;���t�A��^�-m�>�H�����.�|�2�0�1eL�ׁʳX����d��nS"�݊�{{k(�,&*A�r^D���C'Ԏ���t��n@崫	�EE-�g"N�����sH���6�̦�ǭ�{�=Z��	�+V�A[�j�wA^����6������c�x�2�t'�ҷ�%FI���9��ͷ�C�b*A�X��,%W�[��;��+0������@���w�+�n�܅�jU��7*���Q�#*��3l����@[On��/p�L�7.�D,V8�2��q�45ٺѸ��5T@��	�$�l2p�כ�פ�zS���J�����ic�	���������f�Z��Ҵ
��fZ�ap۬fG��^TuQ�@�t��R��q�̼x���֖�U	.�X��h-�$E9i�.�z3j�����Qv�$�@�8mm��b���Zu�V�/�Za�^رiܺ��86������`��r����u�IXm'55Ql�K*��e&Zx�QbѠ]�q�F�p�d�f�a9Zjf�.�I�+�ˬ#]#{�(MܷD$0��k(�㖭��U|�cMnP	 Thl�+\Gs�mh{���RJKxѭ����w�jz��n���J˥J��-j�j��a�mjH��&n;�`"m%���n�����B�;��X��K��2����rGn�tݓ30�8��f�X�
d�iS$m 4�����m���:d)�h�7Kx�S^]k�J8��&՗��RU/v�XNEL4+p�ko�����+
�(nM��tv����8�Y��qf�v$-PS[Ʀjղ
#ܨh=�֡�RAK���!��$e�Ӳ�ٴ�d�m��d��EV;����RV�E�]���Q9�нi�,��#ݻ&m�hY�w�d�t��N�;�]�jV#6��6j�ʻ�vbv�,�~���[ʓ%������
y>Ow/r�# �$�d(ّ1���z���~JM��`���'*M���&R��'�*{y>Ӂbse��^MD�����|��h�Q10+��;�m��)a���Z��/&,ͅZ�f&�Ṡ<n����a�viv��7p�ae�٭#���VEb^!�M���P��,d��s&i{h��� vsn+X%2��@�j�K��Ҕ�����C^�cF�3�Bw#��$2�P[4ඬ��U�w�c�m�ڕf�+J�.���A/2,�B�bP���[��<F�K���c
[�I�Y��x�N�ʑ���=���{tp�u����l-M4�]0�U�mV���r8q���vn�U���Ԡu�ܹ�޼��D����ڑÙwW��`!��0l�.�n�p���Z�w2�GF��l��&��e4�Z�/E$�l4��P�"pAL�+b���Ԛ
����wd�;X��d��0�"�vR9Ol��cͭ`:����Y�*(�ݲlWV�e��1V;��p+pb	��:%ͼ�]b��ӷh�R��Q�nb�0i�SrU �T7��sX���g�S���V�Z"� ;�Z��]�gS��ѡ*�z��^�ѵ��Q�^�Խ��٣i���D�([D^}	,T�=��(��j�dܖ��ޜodj�f��d�u�o2����dV�q��;���-���� CNT�JX���[qZ�sPE-ͽy#���VU�e����nَbIŖ�:�f�]����c+/,\�jU��b.17^�Цi�ڹ1Ò�.��L���ي-��2�V�b��-�B��\� �w�����#��������E���Ɩmn�����u�4$��4���Q_Gءx�PL�h���q;���Ӑ� Q*�9TY�E�BZ�쬲���ǻI����2ӫИ,ѹ5�nL��-�UE�F�eU��(:{�h�X��i�}��dp�H���+��s
%-��I��m�h�ȍ��QK�>W2��]�Z�Ե-j�Uw#�"7��4/5WCd�6�|��*D颓&J6�S��55������Ԗ�ާCN����Xp�M�I=�%^3C2H*0o3�P�Ե�k^f�{R��zB�r�3�B��T3#�٪u��	���;0�5���Ro�e���<�6ED����-��c�#VVd/t�QX���m:fAW�&`�bZ!�{WX���f[�Rm��n��(ɕ��y�t���i �h��Ҷ�Sǩ�Tةz���?��-j�a�Y���R̷�KZ�n5�f(����z��l`���\����8T�wn&�GR�u6���StީY��2�)�d�J��nm؈��Ȅ����ā�CP(X�N���T�$�V���,�W6��a+C�@��b��Xt)+b���oC�x���bglV ��B�!�m�d��[���Z�o}�O�?�c�~f��}��N�3������_Q�'�����N����ѱ��7o���̭�z�3鷣w��4	P�5̓p���s�8��{��%.�w�T���	��QT��h�۹W,sfJZv�D�"��^j����3=`l
oO�u6�V9v,	+�e;�o��v��RH����������Xs�/m�{�ŷ��˔4Զ$߷ w�Q�����R�T����4U^�3f<t�(��ި���.Lΰ뒵x%%}#	�#k��3�߀1��P��;��}[��y>�Wg���S�!�f8h�@H5e�FV��`�<�O�����oN��y�.�[�>���v�w�l��"�m�ǲ���8�أw����U��=��Y[	�H�-wn\�Qw2+�d�`�A`*4+L�	�r�4y�1\���J��Ֆ��}R+Z��*�9z�·v7:��"z��q���w�3�DZ 5c$=���8Cm�r�7�����MH�Ja�XS����s���"M^^��S�7�R�2�`��.�j�zU�=P�OP�.c��6�z�;ݒĔs0=�!�oZ2'�nWwC��ʼB������cE�B�mDK'������/T��{sf�;$���)�S\ݘT���i����{6�Z��/P��gls��4���V�M̆�������`�ڝ��.��� f& ���ѓs�'S�x[�(�������7��):}�.U#�M8XC30j���,��r�%Z�f�e
+	t���D^�<U�1�K�W	Ky%�������]�*Uؐ�۪�,[�n3��� �'����,X.���$n���dRb���K�#�jE�X���&�����Y��t�K,�z���Q<X�I��Jƒ9:�Cك�*�L������ւ*L��z�l���=��:x��3X�j=����)j����+u��J�R��R��&<�б����j@���70������٘Q�i�n�e��
�A�%�5�fV�ճ��od�)R)�>�"j�t[t-�>����:E9l��qa�j�(��>XQ�qސ���B�h��(�EK���<�2���ih�s���}��sr��if�m*L�6��`��+rb�|u�x�
}�;�[o����c�b9�j�p�^�f;�U��˓:ăV���9�[tˤ:��G���Ȥ]�v�\�Ă-뻶�kmud���b[eL`�[
�sq��,V�m��n���cF�5�aN�*�Pm�,+]:�7e�}ɓ�Em��gE۾fdn��cpf���H	)��>@�HgF�į'q��'��۔s�nRN��a�.�s.��:>ҰS��:x p8*M"��/�c����d4�A-��5�����]�sx�N�q����#�E�W�yj&�L<�,��ԛ[y2�w��7�V�[���+�Z�NtF-���7O�_`c�u��wI���$��
8�m�#hf�9��w���;M+�i�ԂY��s�i#5�o��o@u�[��h]"�g��pe�F����.�)� �KAʇ!���*����w_2�`d��3(Wb��2�&�ޥ��ĮRtA���7&�-b�f��q����8NYD:_t=�Qܖ2�P�;%j�߃�sM�6�b�H��W��|��9�tN�v�	řt�-x�v��Z�B���D�u�fV�E�wȶ�����j�0r$4�> �C��&��@�ɳS]b#��7X�ᆲײ�S�G:��L�n���%�v�sF�j�����l��[%�vۙ�M���ңJ��2�-�˼ǣZ���V[�V��P��]�>���|�N��]��)gƈ��v�A���i]���
��\���$��a{���W����W�G��X7�W+[��ȗpS��r)��X(v恡h�r�ں䜆�%w�k4|S�6�<ii�G��A��;��͐���qs|^�t@�+Vf�cUS-f,�����EϹ�c:B�oJ���_J[��a�;�y�h	1�V�7-P튚`��뷺�לX�U�Žzskm��˨yJ���Zᕽ�j�S���40���,�����p�ɭ�Qv#��l2��A�_�/1m�_`b����W|���8���x�w�<R�[��3U�s%-���A4�c�# �ʲ�6h���,I/��J�᷑�p���.sЈ�4D&,�+��MU�S� V<�F89N��P �̳�^�u)�!*���ݜ!� �>��zV�����d�yM�cv��ѥ.�I�jg4w:�D`]��:�qŃB�vҘ��bv�ڻ�E��E���a��A?��_]<!u�B)�ﴡh4�J���Rf����z��܆Z����o��Fܽ�tK��2Yh��\7�e����ƜC��׵QIw�`D+aWƞ$)���0r]�F�̆���ʜ��K�w+�A(�eȬ��+/����aN���0r�Km�zRX�1DvQr�"捙J��:���R���,�}]�e%�v~��Lg1�,�fU	�#���+p�ʎZ�[�N��Y�%���&Z�1]y�<���^*��Ê�rn�i��"�1>�u#e���8�HT�Pk��ȡ��{�����8.�]բ��2�C������w&�)�rj�܊��,�ɪF��S���U��X��lv�U&]�PAE�Nt� �/�`Ζ�ڒ��4�m���n�`��"v`�b��p������s������ X��ء0���&�Y�V2�f�m��,=��]�������s���鳄/\�W�r����WVf���+�.��oGU�#����Ԧ�Uv�N�	o��1"�Vړ ��%�*�D���t�N�HO��|$��B쮝�Z�ҵ}e��m��p3ٮ�8X�טh��+AN�����^�e��Wp���}��R�s�[6Lu�!���}D��9-+��rT��BvRu��-���z�֦۩J�:���2���j�ŕh��A���NQ��餕���L��+�v1�NZ��1ƺ�v�oc�d�s-���6�c1]�'P��"f9�v6h��Ѣ���V��!�ظL|�J�C��7�g'*�[<���q�Hw��S�� [:����Gu*ތ�~�h��怬��M,i �2�:A���.o�Ѱ�u�k��e�]*ЖQ����rմ�.=����Z�s5��vYu¹��t�keTih
5ڑ���B:J&6	��6�Y�[v3��:O�+��AQm�ȒbLM{��z�缠�j�t��j���L-�مD0f_,��*J�u)%�׻��At���6gt#h��{NI��ѻ֦ed��[_m�(;(�9�3�	x�J�}X�-h<��\�5�: y�����3
ƶ/oh#�f��D��{o��{��Γ�5PΛX�l��[��M����MF��dȖ�tFI��٪1���h�u�H'w�����\��Z�od��!RQ��Ff@�1(��6)�(��'&�RfP��I$�I$�I$�I$�I$�I$�I$���$qI�qcI�5��KN�����ʜ�:#�e֓�2����gU��F�a��u�*��(�h1#b�>�y:�l��)u��m��u�q�FE��P��3Nk��qۇ"YJe5}��g]P�fjS�]�ָ�f��h����N������b�����
�#���vs9I�88�9w�e�J8���:U��tn�ep�_m�`��h(�e�n�c��%Cǫz�!t�]�M�2�% s3;�ڪ�!���fv���v�t�G�Gn.����J^Y���w.��\h�E[���:���tl�e�Ύ�3�����	6#{��[�UK�;$9�[6"6�;:�o�m�f���m���D��Q��Rm츫��We����֔��bn˷9f��J��c�u��C%L�ǴA��M�u�nG�l�E��ȋx�����Q�K�Y��w՗xg��E��H�.I}bZT����5n���w{�\Vh��_��������>G>~S��j((����7כ�
(><Ш��{�Ȍ��&� ��?i=�?�u��;�o�6�i���="TE�L�{��!H�a\k��͔7�N�V6_m�N�pteabY)�ΰ�P�v��R��vYz�k�����U�D߫G,���5d(�P��f�1�1�D����Y���c͂�3	��iU	�j	��l�sd���X�kz���=j�����f� �	e;�/X��C,r�2��hoQ��`�$;�AqبX��	�D�j�3�Y�����z��rv�����n��}E��r��#wF�7j'Ӷ�diG��v�
Zol���J�Rʎ6DP�bTÜs!Tl1�8�6^Ch�Us%G���OR�o37�y�ȫ���٩����^�6)j7E���b������霰b.Ҏ8�Ϫs���ꎠ��ha�=�#��i@���)xbR���U�p&�@ƬD� �AJ��m��,]2��?ve1�׳��Ud5ӝ�'�Y�Y���t&��W�%e�u@���W3+��%�Q,"�����c�������U�Z�M��@��X�X�s̊��F�|�)z������9:u��*�H]N����tMf�'2����f8�8�Z�a�hܺxC�#,@YH0�|@�C��OfVXx}�Y�$"��X��R�2�|�(��ՈY%����y��\�H4�����#�U���*j3��#g.��-�B���O%���]�A3�W���][�z��hE�&iʬHbyF�]ʑ��
��:����[�b�����	��^�I���n�����9����"�N#X�����@Xc,U�pAFN{P�=<���SbO^̱�GJ�}������BkL���X渘k"��nr�1��� /5-j9aC�$F� \�u�/��ֽ#{{��.^`&�ػ?44�)��RH%]�w[ām���#�tJ�^�M<�Ұ��U���WdA�������4�.a��Y�C�B\�ʙ���߇
%�&6�o�,�9��cn�H|�v�L�CQ\]��WM�h�x�ڰゝ�
�NZ�6�Eґ�R�A�?Ej)۷KIf�P��lJ^Y�%�R
�U/�r��g��T*[��c�z�R�r|ve�x��N�-�N]m��K���t����Z������Jn�T��
�Hu�pdG2�u?���7.a`�(�P5�V��h`�b��F���2��Z��0z���/me`�Q	��W����V�[�����K����j��j��p
{T�\���Wk�(��S�|�63F\��󒯈��ƙ&:s���]�m�.@r�A�b�3�V�#�V��x%�AU�rh��'Q�m3}y��x�L��.�s.`����5����]�����7GZ
��DW	����$�|�fXbrmD-���B��Q��a��5������Lv%ݢ����=�����/S;b;a��O]M:w9k/l3QK�@帨���C,oH��$�]#L.V��W���d���0�<]8'��N/mH�]<��T��8E���
��1vŖ�a(�cѡ����Uˏl-/3_Е�6��E�4�eƞ*8+M��E}
�ޠD4ze[�S�ʰ�bx��l�'f�NT�Y�T�y�"�v���?s#\�2��n�$?�:p�g�RyX�e9�j��p�6�i�M^�(Bir<���ȼ�Y+p:��`�Y����0)��\�ND�ms�%R��c��n>��������8�ʢx n��z�M�5]!Ԯ;F����@���	��_�-f�U
N?���B# U�J�p���b�ʻep�� ql9&�2�a�<٠HPN7��\��^�]���Q �r��#���m�Uݜ#�w�k�pl܍hE �pO��J���M:���3/�N^��J��>ë%��ޅCXq"���.�{���l�֬:o0Pf�̼U�&�B���L��[$ nr�J�G&HڽE�0�_��XvÇ+Tq�I9-��sUjFPn�WT�9S�^���a�iʜm]��+q�l�¦MA.�d��Ӊ�p�DBpUA�K#�ުt �OEՊ����1�1�x�!�HP�u)�tBm��RPA��_
��J�i�D6J�Wa��vA�ge��L��ʕ�
����2����+5UYW�:���GN�D�����2����v!�\13R�>�$3���H�ݗQ�˲a��C�Z�1`�����$��otSʂ�x���߮�Q��i`q�ҫi�]�e#��oP���N�\��k
i2VI@N�az�t�x0ld�>�g.d���/.\��9VF��N#]���0��F��4B� o���F�o.�un$,˻���J:8�Gz�|v�)s�J�q)��`zq#��(��{1$�0�~o[X�1�r\U;<-m<@�[aLq�f���m<Ye�f��VcKM�Ñ��a�N4k���ƽ����1�9i��U�z3�Y�a]{CKc��m����]E��$ݜ��q�:˴��Q+PL%�Dq`_b��0���TH�8IJ�T���}ue%����oS3�3W7E��u��m���=��w�6���ˍ-�μp|���T����}
cp�Ө�}��,��H�zs�
ݍ��->��g!�0�-�QXl����Q9��F<	r�)���Gk���fL.a�NU�b �I.��q;��R��t�Pr�8u�n��ܨ:��(�bPF.��]��lE�N2Ȇ��7�-�%�l�!�u1Xn�`�b��Yg�⏮��r��憹V]ѫO��J����W6�nfRDX2�i�v)+�HҪ��P��I��]pعx\
Ҋ���jiͪn�m���PVe�n(�Jv�3w���̎}ťu�u�B͋�G.���>g*��ꐷ�c}bކ�\Bb�ܪ���Ze��#$�l�	μ/�VU�j�q���c!X��6���0�xEM
���^c��[��2���v�)T�`��T�i!��g2��tK�`;���h0GÆ�����U���y�b{g�����N��
��(WK2�Y�c���v��yP��I�\�.Kx6���wv�����Xl���HF��N�ݽbe��	�J!�&jkE&��Jl���{}H�it�g)t�k�u�1����yB�����6j_U�2X1]o[.ī����F�b���y���Н�Ũ��HXJ�$ۜ�t��3�i�80�6h8˼35��J�[ى��J.���BJ!P���=��CS�[�5��v3�5�mӴ�o��2��.��k z��^ �:kL䘲br�i����mnXDT�M�OXy�����אu/J�P ��lD�#�z2ug_�T�p���H�2��.��6��L���wtS6�� b�6��2tU{�0�Y-��28�,��R��J��	6bs*�k�v7�GJT�	�Wo�T�j�9{3{^���d�TP�Zm�,���J��:��e廵B�� u��$�Or��za����k���F�����&`��J�)�F۰�iWN�:ڪ��g��5s����vT��k{�Et�]<�`��&uxrK����&�>he�Y�O��]�ʴ/JP�b<��d۳��9Q��m<;�l���#q��[���m�(�ٽ�$�ʏ^�@��OpP��a����{p��ɩf�93-a���`��b��>	,�6��R���ݫ�]��3g�;)8�W�o`T:�I}��eِ�,���ǁ3+U�A�pG/�4bPV��vc�e�]���uIf�nt4�	̛7�{��gm1K*ԬV���B�!�mȏ]��&d!f��b��M�3�̓�����a*�4#�:��U˷�>��> Q�k�����p��9����D��>�ڹ�m���G�~f��5+t��(�Y�:�o���wu��fX�Rr�	ݽ��`��';܎|Cy��g)��Sw䉦�ҪEi�vl�9y�Ū��6�gwt����Md��>�"��\F{xB��u��d[�ŗ��S�M�qx%i�O�ʊ��i��H�e��:���7���Ef5xv4.����6�3M��c�nt��
�Zb�����>��ռ��q���
[]u�9�oAw;JS��,Q'�*,|�huj���p�O�	����)��,ӊ�lfV슭�P����$��8S�w��2;�� �QR��&K��d0�6�u�Į�/����ᴧou��a-�j6[\c�=��հ�h�M�3�kz�XQ�Ī˾�,�ݥk��-��+r O�?=S�����ĺ��� ʆ��iF���ue��AA��䡑�2�"
(R�(F�����w���)F�(i솑&hv� �
L�22A�҅m��4��T�%	M%� �	@m���A��jĪ(�Drj�h5�KIH6��hrv�
����z��?3��c�)�zko֞'r�T�n���i�2�
�}���Q�;TRM����r����Zk�Ⱥ���޹P�]�kM�����6y�E��n�r�MfX�yy�`���r9	�="p����%��
�P��˟]`&ᴣhل�-9xu��
ssWMc[:zh��y��"^��/���1�;WPj��>Gk�^�/��S��=PUQ|�
W�Vd��g�~�u}�<"�<�B�@�5�<���,�kI�G��x��K���ޗ�����3�5��1Q�ԓ��e�M=�
��ؼ�6��{��Z�|&Okܯ{�FFb|��=z͌�+Ӡ�惚U�~q��q�'*;��N���ؒo�66H�IZ�z�%����[�0�VH�F��\�8l���io3i�)���Ŋ��j�*{r�X�̔����9�=p��u��zP��kWp��� ��7L� C�ĵ�� 鞇�P͕ݔ��S;���ej���/pR��]����<�]��/I9ɱ1~
�{o��e�jQD(= �����|l�.���J��f�C�E*:��tE'��I{��ڎ�zӬ�ޏZ��jq�/���:����.�4kƬc
�r��-��G�W���C{�/�u���\9Su�ŉ-�(b�m:~�p�j����88��G;ٗ�*�7�7�nk��$��$�c��(�s�KNM��}�F�ɷ�@�yb���($�)���'?x=w4�O=�x�?N=-<5��c<��t��ZX`�(��ߎVdպ��j��W��7��G���=����JH;pu���ᒞ�2�Ŕ��*4sV66xNOqW���C��~����i��N��0zuҼ���z���rv��M���@�*�p�gPIonʍ��fPCBFoe��T��m(�}���䈵�υ���D��ܳ�5��)s��V&]��m��D�4rR��Yhhֵa��5�彻k�芢�ʙ�YwX�i;�*�8�ٛ#�їp@ӒF�^��Ì�߭V�+S����¼G��O�ӫ�c��2��e�s��u���ΐ��O��Si�Y^[�'y)	w�3�`�w3cu9S��Ui��]�Z�P!9�[�oh3�ٌ���Ù>�"V�B�S�8ꫳp�lێjE���Pś�jWʳ�r����T�:O ��y@Ƃ�Ҳ�MƸ�Yy�!�a����Ұ%ו�j���W:0M��m�,qXBw_�lc��^j���;-5J�hm���7�D�i�(R�L�9.}���Y�_K%��W�Y��u�i�ת�B76R7:����N�f¤��"��*8�b��U��⽕��9����
�٨�W(�Ⱦ�i�'��ub�n����،�rt)�����_v-�֎�[�[�[�9�`d�bxjg4���ăq�CU�jY<=�ѷ�ɻ��qA�;%^"�:���������M��vS�/�n2�hD�K�-��ow��b�t.�s�md��NM�v�\R�u;P��;6z���x`6�P��\0��t:�=�I��>��K�G���z�u����H� U���C<x�9�Ql��2U�6kQd�e--U����♍����u��ݼN1�&��ǔnYD�h���ڋ�E"gc� ��W��������@?�>��tqb�fOI����
�S�N�H����]'ww�ૠ���̪)��Uv�Х����<�f,֢һ;׎p4���Ţ�'�6Sz0���A���Q=�"�_@�ܖ�4!�Ը��(�v��q��=�>:Ǽ�˵'N�/S�o��]EZg^��xM����o�m���Z�i�o�m�1��Ewkd6"[0�7�۵tt�/�|)��׫ҬH�"{P�Y���m���ӽx��5��㭴&f����N1��u�T�Ɂ�׽�>�$�G&�H_){#��8N���{�a�S��j�n��څcz0���N��g1�Yu{�;R����1����px�b9_�]���}E��GX-�R~���j���5WR�z���׃/���'d6�c�v+��:O���f!A_k-��m��$Eb"z�2:*:ȋ�}y;lj��IOU��-�W�
���W=gwe�Z3��miA��o3&���S��,��t��\˭{T�K�*��{/.�ǜM2�n���w��#C.��k�9d����q&C�h���+u����� ��̓9���C��^���0o�����s�c�]��U����%��2���W9���<�F2j��$ގAK(���1J {����io.�������K��f@�P�ZM������SB��DémNT��O<�#7�q����Yʓ�۸K��N��f���W٫�kep���P�yuM+R=1�G.Y��p���k���+a�uC��1�lX�rm�!�]���7'�7�}��!�Sp5��SW�^��8����_�E^4R��y���.���P歫U����Y���FBY��h���;ː���?�e������!�`"�Sa1ε��-C�����,�-���P�l荑�\
xT���O{'j7	���嘆W���!��`ޛ���2HnoG�STL��T��{�����h��{AN��o�pAi�1w&��l��f_'��VN��諾����V�zTs�ӗ9cY��ظ~]`�gE�z $��qmɽXY|�NY���سa\bm�śd�������Ⱥ<5�M`1�@��I��%:'bU\����,�i"��
���[�]l���D'�t7�k\N�
.�|[��xB��z�5CT�M�3G�z�Eq��]��ɣmͧ�at�!��b[�#�V?�YB�U���d5z�f_ez�>�����ƻ�L�'H(_eM�{j�.�dd4th���d��q����\�͉v�%��m̱Q��N`#�V�>��g#��%)%o(���r�/	��Y���1]s-�J�8��[���z���$̃�c��}	>1��kݧ�(5|��u�ٻ�K��v9�j9l����Mg=NƒS���*�#��P�j�C7uk��ћ��7�.�����xvI7y�bmէ�G*klf���
�C���ayǧ}&�)�o�X�_�G��V:-� 7U[<KAƍ->�����Ʒ`����b���s���g���:f'.�Aϖ�;'�a#צz�6Q�t����z042�F�ԃ"�P�]��4�u��M�jy6�X��mY(�/<7�)V��f�H�8�c�ʕR���hʱ�T�i��X�Bkڕ�E�)�븵y�>ZUI�j�WT�[y��w�Z�5u&����h�%�kY�]�ά`unK�
d��KѠ��y�ؘ�s��p���ʑgM�{}��G����3�:9KojY�;8���9��9p�B��g7�s�:UZMA���W4Ws�q�Gm8����o��h8a��7{F�A�r&[�eԂ��e����w+^��0�:�b��Y}8:"k�h�o�K*��b�����dE���eG�]��-1��M��l+f�E�7I��fj�y����s��7	��
����z
ز��ԩZd�ɡ�P���e�l��Vlv=_�>�+��}g�.�掸먵�E�YS\�<�V]Y���4)�C�u���D��SA��]N��k�̨&��,6y�q4p T���C{�d�xwXX-��M��)��:��D^���<����L*��q�X���hͪ�r�t�����֎΁�����,�כ9�[��`�f| �j����k# Ҭ�^�y�����\�R����Q8#W��)�f�V�awkt꠽��K#��f�d�G!�SsC���`95fi��+@�:�Y�V���L��!�����]՚Y�q'\[�n�x;`@�-�e5a��#�rm�i��6gk��'��%d'4�t��mq�5�ĝ�]jsb"�Mpں��!7s�3�=Rq�G5!Em����y)��B�_�`ʪ��P�KMDP��fE&NB�STQ���y��E%%+Hд�CE+���jG%�R�P䚔���
iiL�$�p�5�)))B�2r��
h�i����Z�i����jP�������Z)h
 ��)Wجg����k4�����s]%àܕ��ي�K�Ny9I'7�ڍ��9��3��� ����
���/�q� �zkxbG�yT�w�n����ښ{9�w�u粏��l�쯗l��b�x)p�lS��^8\���^�ui3�x�r��fcD�4*�/_eh�^�k�ۚ1B��֞R	8~��]'=yo�4
:�YwOz�R�{7�0;#!���n���Bi�po/Ϫ��tc�	��v�2�te˥�t��9����WY��N�q��1ihNc����)�dO�n`t\qǵHk�[��)9Du�wrU5�U��v�E�OR�5G� ��ao��S�J�n�T{O��t�Ա�f^7r���Ÿ�e(2I�) 8d�vvO�LL:�O
�^2�;ed���.t���j-On��,����x-r�zO�k-��,���yw=F\a�p� &��-x���;rB�{'��{ݽ�k��X|�����n9��X�un)Wk㘦�qBVBMf�q�Y��A�B�;d���+zv`3�Zȓ�$�3U��b|S�)�Ȳms�⮘�}��lu����ЯP��b�Y��������ō�ɉg�Ǟ��&�P�fLOɎ��!��c;6$}D*�e��}n��q�X�1g�a/�p��������ٕ�Ҋ��t8�r�wKWڶ�۴�U$�u��9��p�͎9�~b�,dnKbo���Q m����D(�o�SU}����8��LZ8�nK<O5�+�Mb�<��(br���.|ZLps��͞��k_gT����4�}����Wʠ�dʳ�q.���K���e�pO�t���GNq��ǂ�N]g,�vHM��(>ӣ�V��Ж����\�`M�3���@�X7�/J$��9�1OU�MM�������q�R�&�t��&��2�c[7�4*/��i��"�ž����v�NK���e:v�;�J-9!#�ۂ��fU�|�6':�9޶k��vh��Z;�"��s�����	t�d)��/��E�I{{����[E�^�գI���kWpټ�i�f�x��ޙp���i�@u#�xi�(#R�=[�b�%�E����na`�G���싨�up�{�\;{�\��]�򇲧���9!K��G���G�#op=�5�	[�m=J�'����9��Ny��̸5�s��Ͼ!�N�ް��]����B��Z �e�_m�M�Sh2�G�7��S[�ɭw��u�~s�^���FJw!��%��� =�Q��ɮ�S�ii}��X�2�:�z�Ѷװ�rq��z�7뾽��8�JqsPu"Q�y)ԇp�HPs	Cԋ�X�]���:Z_d5����o<��y��v��}�㮽�S�5�=Hm��h<��z�8�$O'P�!A�X亼��]u��ּ29�~��}�[�Ro+��w�u���v�8��S�h]���py�8u!@�C�u�m/2�wϞw�{U�r��f��8��m�^���TR�6{4��d\-_J�:�Ys����,x'v�a*:�o����]��t���i�=�G�`i���z?:��5>�n�^�(Cx�wx�:��L��]��� v�:��2WS�w"k㍎{�l��7�޻��]��`e���C]`�d���w�d)���S���;�s��
7��$ך:�m��[u��y�~
{�K�Ԏ�xs/��.瘾B�m�*g8�Pk�Sx�Cl�`�6<�;��!ok����8�޻�|�Rzs����Ԝ�P���+�Ļu�̯R<�o�N@��CY�R�A�u��׻kY߼w�}{׾�w{����=Jo�)̼ɷxwy(lu�qs#��h�x�8��x���ZSy6�~}�5���ﾡ��R&���.�}�%���_e��9��Ѷ��/P^H���y.�����՛w�[o��߻z)��Jw%��B�Qԩ�w/wr�fr�/�n��H�qs"d��=���Y�U��ζ���x���P�u�wԴ�0�!�	�h���v��}��@ռ	ԏ&�qy�׼s�]y�܏C��G�XԺ`�W�;�68Ù2B�^`�Hk1��6�=�@�إo)��������}��n��|6�;�Ӭ�${���ԧ��X�py.�*w!B�s&@q�̽���o�s?��w��9�ڷ��ov�眷ߝ���!�0T�W�S^�Wr����L��.�s�e�Q̅g�Z	�0�牲���UԖڝ:S���M��o��x�\u�>y�w�b�Ԧ��Խ��9u%r�O0R/��*o/�pk�|�ί8�c^��}��~z��̽Ǻ�z����osܧgr�'R%m�=�u	��!�/P�=ü�	�w�֮v�wߏ}��5�Ĵ=�xfj�9��S�l$z���R�����k��r8� M���N�)9�q�|km��Ӱ���\�.^��s��q!����Ǹ���x�G�y��N��v��:�6���j�{�<�9��O$)N ԝB�!��Kߘ)�Z\��:���C��#����5{.�y)�;r]�Ϟ��~���ɐ��ް��C�|�����^��w�Ѿ�@B�!�c̮񑷘��\��;����ߝ��Bm��)��<��s��C\a�r>\�u��
j�R�H�=�o;HqƷߌ�zמ{ߞz	���/�gpym�2{!N���ph�9�Os/�r;���s��� k�T�sn���ֵǻ�ߞ��H�<B䇦a�/Pw:�7u�ԅ!��d�c|S�|�oq������m�һ�Cq�>y��Z�=�ΏQ2=��S�1i]�:��
<�:�u��^l��CqO%��%;��6�a|��9�o3�w�+�������&�ݦ���,qD��7%b�GF%�&2���ެ��Ju�o��o&��/)ZcWʤ,h���+1$�
�%�įȈ�{�)�m�� NH��ĺ��^#mb��	�;�#܆�1^!�=� �0;����a�N�Ü��~���:��M��!x�RH�{�#��.�`�r�@�=����ԇXb'q�	����u���\���K�xOs6��$9�ߌ<�;���G��l Ժ��_ �T����Ì�<�ێ�3��y���<�~|��E�^��7��K���cԮ��o�T�V@�!��!�s��r���R>s�o���~�ߟ}�����7��]�G�b>��q'p��ɾ	\@�|�>�J�FH�u�A�'s�ܾ�����[kY��z��@�Oq
G�h�6x���}�����-�z�s�S�o����}�M��N�:��4u�}o��ߩA��)=��2D��|Z_.�2մw)̧F؞�Hj=���<�(=瓾�ίw��|�=]�r=�$N�<��߬��S�v�.w�<���!IԮ�c1SQ�{�=yχ]y߻��>w�9)���I����q�B��u�����/w��K�}�r�ۼ{�
D�:��}���>��^�&H���І�Xu	ݿ!���'�
S�q ;�g�x��T�*=�S�o��c�цE� ��'������3*K���6���q5P������E	�e����{��+�h̘���n��)lb�(��$	{i�w$%se^.��=�89�O���DL��^g#�w��k�Oe�� �e8��N���:��M�ļ���=[q�V��wػ߮�﮼G�yŠ�)�o	�c�F��:����<�7��B�6�x��6�9�O8y/�b>��}��֯6�q������~�{����3�Nc }�n�]HPP{Hyɶ'r��s��BI������q�þK���{g��0�o=b2���`��U���I��^|v���EӬ!�	��좱MB����:!��tekYq�'KE�˄,�'�Ƒ�B5%�듖/s�!���D���`aX1��1|zl�GVy��o��\27
����msJ�����7˳�)Rk�س�z>�z�h��r�V��n+�힮\F�����GC{��ft�U�ss6�l�V�=/8���۟mi5��[�(�}�6>og&�w8w��z=�{ֱ���O��q��հ���W
!��jL�Ŝ�q�J����1��׼��`��ǥ��R�t���ft*v���Hp�%�������z,ݞ�*����q �����zC��f���?WVP�� �����`�u�]s���B��s���҈��J��k֚�J�l�ꁗr�\��~}h���q��m����s�M�*'7�����	��q�O;��p7]g�����[��z���o��{���T�%��M.�`VIe��~~k�z��W%��ô=����*7��X/v���ޙ�o����М��nU���z�Z.��iƯ�ᒴ������{ޏG��2�p�&[�����Py�=�k'��V�{O#M����;���n���(*��k��|�'돕�Ğ��Om�ӷ�RyK��\TK��a�t��'ւ����2�ii��Gd<Of���ŕ�b���
���Έ37'�ݪ�=mWA���a�i����]o�]�0g5LN[���;p�5`I��s��V2'�ֈ�;/7]����ͳ�P.�I�Զe_{(��
n���kb�$�U��^5w�a$�YQ�5��2z>�3�~X�3�f�*��s�K�+v����)M�N6�ga��ݛ�냩�3��DҤ���v^SQ��]��R�dѭ�G��}�����
.�j��hd�P���É���o�R��F��j;�b�;����#�2���9Z/[�][��/�TS+*���]��Z�˅!���u��3-�v���Iq�|[j�A ��7s&d���Z�8e�.�<
�+{j	���Է_�)*�,�4Ƀ7���n.�A��J=v����fD-���@�Ցō���� �Zg^o42�b��:���� �Kaֹi<h�/zKT9ѧq��0������Tz��X\WZ�fS�tiP�TD���+���C�K*�)��=*����S��p�a���n�3��D��1Z���3\O'�v��u�C�)h�t��z)����X�+t��.]&��k*m�����:1�>�#>�_[���]�¦�o;+b�g�{Y��r� 8R�o��|,�=]e'�Tۻ�0��s�J	���}��m�����D�+	1���P�F������v�z�;g�۽�4$1Y*6q�˃��Wɰr�eڛ���RS�r�C��ȼ�]h#0m��/�`���]Ho]L����{�����Pm��$e�8sL8q^����7�P�nηnf��Πћ)��y{v��1����'2�v[63o�,U䉋b�E��[t���L]��Ws������Y�l�-�WF���j�Lj���K�j@r�A��Y�.���d/��{dB�b���@�zk2	�����%\�](��+-Bµ�Imr�8v@�S��"OgGut�^� X�V�r��ƖӐ܄:HN�,V<�T����^�b����(�3��"�rr"f)�iʮth��TUd�gŋ��c3,�"(rJ
ṿ5�Y�X�6YNI9c�TY��VY�4PY�5�`QM�SX��f�0�
c0ʜ�2�c �J��0h��)"�,�0rr2	�Ȫ�ȉ���0�
��)�#*
��� ����3*��-�Q������0�8FTY�fffa�cTQUM��Xf�i4mfS3�Y�e�eE�e�9�T.�������s�y�S�����@eg<�0���xT��S�ڝ8N��������8���f�5��Q�Lqe]{,GZ�ܴe����3�mu�c�����Ў<��s��d�lؘ��E �с6���Y�&��-<�:�\<���F�k4���܎�XM�9�w���S|0H�����ӧC���v\�V�)=@�h눘$x���&���H�1{�W��t~D:��@V�|���u)v6�V)ݔm�6S�݂ ��1�':���G�6��5�=�G"9EEm�+8X"[��$�sI^��v2�u���C���*� k/g]KK��z��8�]��i_�I���,�|P�_c�Y�7�Sx��,T�#yl��!p�C���""=�x3�m���=3� ���m�M� 5�5̲�0��,�1]�b6�zڬ��GAn�3Un���Hr�)\(މ�5�䉍�u.h�j��J�5
��G�q��v;s��FiƸ;;�z֫��Zr��i5�csX97;Q4�B��b+9�zo^��˷�7�ɵ�������7w�
l�N�<I���o����!��El�1�W��k�#H��Q ��T]N\U�a��\������#8�3ޓW������R*��cB�D_��z�/(�!^kbm	�@M9R�r�mܫ�V�颦׵���^�y��h��:���;�S[!�B#y����l2O߾����[xi����ʓfxi��5(lhB�\�������gT�.0�R�`x�%G�������r�H+;����� �X�K��P=|_dح�.n�^a<BH�.6{<a2+������.,&;��o-�c��e�.�^�==a���\k��̃\� e�{�TC��1�8'X�▯ =F������9x#m+�GӶ��/z����3β�떡�O��h��.I�ip���S����3�uY��	�[=u���V>��c\Fnsf�7�S�W�
���)��$/H��.��/�M�1x���6�օ#�wd\�L�-''��}��#�Km�`�Yx�y	e���Pʑ�ҋ�*�E�o�#��+�l��#�%I�k\�܋5f
��W��y��7m���l7��N�ɣB�"��p��殱Vʿ��7��}@-O���^�,FjE{���.�Z=�m���e�m�9ÓC�4͞�$�:&��PTk�\��f��RM�R�(�F	 �`��ɦ4�e�/ �������4�� =�3�?y�NA��q�=[Y7ݖ���1M`ҭ=�V���]_�Y�mu��3�������AV��2=�d�)K�:��/�fSR���̕OZ��5�1+,��+"W�!ڌbJ��HÏz"=|K�lcϽ��7k��Z˼`�۶Y���(�����d"nޫR^y���`嫸3��WNP����ƫx�e����랜Yi�<u�W�`$�鵙��之�+V��W:⹒�'=��1���lgD̔�IB~ݸ�Ń��aC4"�n,���[�<$��Ǯ�-��6�+��5v���B��W'�D�i���޼d	r"O��)�����[�>����΢�Z��ٽH��rx���g��7N�	'oن��ܫBY9���I�b'hi�BCl#��=.����r�:�RG�Pxv]G��۱��aĺ�2�s��U�Z��K@)}���ѬhI�����7�ڃ�]4���NR� Xa��C<�n�s�%t8�p6�����!n&�iuw�Y������A�; a�q\������ʩ������HO�AкL�
�}~���ؽ�1k���fN*����:�M�ɮk=��c�$�+��ֈtA�T(Z�s�dZG���#��]�
�s�1�X�鵙�'��և!h|{ysOoJ�{7�_n<њ��1���Q���4��U՜��5���{���j��C����x��y�1���9���vD�4�RU�귎X�V�'�gvT-�yՕf����=qat%�QVWy%�z#�w��n����
�G=ӓ����S����ⱻ���' �3є�L&\"��δ̬8�,�\-�A�v���a����uq���e.r��T�D$&�v�dq���Y��4[ջ-��
���phj�����^���{A��a�����n�w��2T�<�L9Cm:��ꆣj*����ݗ�O�.�1;�]�{1���yȷ>lmy���N�Ő��do�%�):��;�:0�`G�Wb��F��v�g_��[/�a�jxl)Ԅr�ղ��z\Bm>bNVK3�8��q����s���1�.������W`mH��\�rz���*+;�WޏDDNv&��{�C�7�iv�����D��vM�Q����E��b����7v��n C)C�iY�N�2Q�W��営tna��3��m��J�R�윋�R5���n��j��VcKZ�i^lv�f��-&��%�͵�c�aŔ��oxlp]4��ʲ�%���N��*/�,��]���̍��$��ײ9@S�_���\�.�s��ooqa�3nELo<��I�6& 86�^��#�}����h'�*Jי�*e�ȼ�.���9��ƣ��A�<�0��4c7a�;��杽w���#:�WH���3����;eڙ�XYd�Y!�&r����E/����+����_]
ԗV�p�h�h��n�-+��f`V��Qr��&�ᰚ�qY:;mŊ��p�;]񶶯#^�#�jn7�)�j�-:�v>Uz��Ӻ�G��G^q<��W��V�]�ٱa_&��qƺ�r� I��Ьd��$�6�u�:�@���Ov;�zM��1��%&X�٭�k	$t��ɚ�0��6�(K5��zvN�lr5���&"v�8�g���˹T�±��P��˦"l����W��̝]�f�@U�)VM�5����'@�J��6rj�T�2�bn�ΈaS2����R=ܪ�Vt$��z=��ey�e~����Q`UΏ%��w�r~�^��̈́D*�T߭� �y)� ڶ_7=ey��#�\��+�{|EcR,�W�gﾛ���l�ޢAnOP3{�
�}u�$Y�&0��b�Gi�˪iW���ߛR��:���n�����q�r�Z\�n�ѮC5�|/Q��ǐ��Ory�Lv�Q�)�C��8�C�S|��qC��� QEO;�S�ʙT�ڊƵ���gl�rya��P�2�1
T�E����i�>�s�jbH�=C$���z�R����һ��|-b"��ͻ	D!�l]G5�ӰӮ��Cz�˱�G�:��\l:0H��	���1���j؜�RA�&cyD��zv�j�*�;\����T����k7z=�����G�]��$��kT���m��γu\f���"ҩr�Qv�͒V�Ԧ.e,,_�c�P�O�Q�ޮs#�7(��IZ߭��j�kg9{c����YF�8nգ ֐�F��;�k��@L�2i�p�@6��ֺl#c
�=�x�ֶ"N��F��@���e¨e�Gp(�u*snZiDV���\���Onk1�Y9��P�5�-N�\$�Yӷxĕ7.g�f<�m����G��bN�:�3H�8AJ,c��ClZ�s�<q�I�u�h�4�;���w89[m�{�&��3A�����y/�n{L����Tuϐމ%{�hY�:nIj]�b�V����b�2 ����¦`�F��»n�ct���Ӕ�N�+�L�/G,�fnPS��֚���7U3���d�:��"Ҋ�¢��f���-ZGnwvj��-u���[9��݊�Ч%L���x��0h}JoJ�nu�I��x�q}[R,��U�ԕ��oJ����K}Ϡ��eb���I�ܔ������=XoV:!�ݖ�oK�����
�-M �%n��ӷ�!�vidX���V6�畊hE^��[�Iّ��'`�T)��vR��7��O}#� ve\�k�,ڕܓ�i�Ĺ�$��|�٥ ]��
ԑ,��c�y�TH��t5tC��{v
@���vi:�v�b���J]WFeRTE٘I�cQ͕K��H������*���Rd3-K�5h�i�(��)���5�UPQE)T���MeHUSma$PTT:�����o��5��繬��{���;%,FRt;4�8�IsKj������DG����r��֥��Wg$W��P9+��<��)�+��Lѐ�v��Lg�3S!�|�9���;'$��4	�2Ds�Oh)
g^mX��P �i��7���*C�;��{�6�mn�	��a�:ani�jo^>h�xoR�B2p(���6�e�u�j;���m��J�Nim�|�\%uB�D5��{l׻MË�ζ�FbR�����5��whUn�����
�N�:|=���P\�����b��P��j�:1F.M#�p���&{���*�O�j��3���ݹ�1�W�+@�+��;M]�-�&�V(f�R>�&N���ޏz'���b�����1�gs�%\�1+9�%��1p��*�8�ƌw�.p�\���p��nC��k��W�h^f�5�� �쪥�َ�=�W���ԡ��K�zB�k)���q���j<ss�l�.l	ʸ͵��1>��[��r=�D���
��q�qUȲ��|UVk5w��K	Uq�6�CP/��_%
��3�sǪ01�"�x��`�K�:�qvZ�������_��gd:��Mq���ogP�jƹ4c��L�Gم99�`�3U�5����f\G8����ʈ��p�-YW�!	f�V�<x��{��u�)�����?=���J�/Sk�c4�3��ܙc�o�K�F��I�⯦�կ�gZ4�	�c:�c������:���m7���ݷf{�D�s���е��Zp�n��Q�hﺪ�c�í��ĭ��Vn�Ӫ=�E>�Nz�����{�6>���h���M������V*&���]��R�h̩��{1��Z�%O5lr�A���6-�A�=z�2Vb@��'���&��&����9M�2�gq#�ՕbR�����^,�D��jN��:���2�f�#�Fq����3�s)%i��.a���M��% ⾈���w�n�t�/��DQ�����\ĭ}��,�R�
ҫ�PI	�"�L�����~񽞷�t5'V���z
���M5�ƥ�D�)�7�F�-g�n��V�D��p�S��q���[l��Z��w��C��5�����;�iX��{�Fv��dt�-�0�Ůq�R�k���YY��#Ԗ$������������)Q25�A��J�g��0g��CȒUc�&�4�� ��K�G���+i�+j���)�A,����*v7'4��U��b�����_�x�"4��:>I��*V��h5Q�Utwvo�K�+��\W��,6�y�G�CO�e
���I� ��!4��iN���4��e��sW0'������11~ب�\)��Wy�*v��< T�5��/B��$�֣>ƈ��qb����~�ު>�a�y�X�
�@4v��LV��/�kK�����#Z��"d{�C��!z��<uI�V�j��	����%8x�;����B���ۓ�;}��Q~VC-+/½S�W�t�!R&�u�ev&O?o�>��{�v5!0 ����i 
ܭ�4"��}ā�W�x��k�x���
�^�7�'*��Z����\����yU!��ޜky���˕�I}-˥����k�<�m>�J��ܒ�Z(�mZ�m{f���lsB�	���5�[�ob�ɛ�m�wb�\�c�r	��m�2rN~}UU@j��w���\�$:�z#�_5v���1U�=�)
B7Ǻ�z�7f
$�f�"@,�U������㺈{�h���/�Xi:����l�s�I�짧1a�,���"�,}�YI�|�<���G�\ TR�O��j������xS�F6E|�ư�"� hj��k����E�;��2ʃ2��y����)YPg��I(2J�U�G�o{ن�?DҘ��®xW�wpr� 7�����z�BH��EK�	=��鬗��1��.!�ϻ��N��g�w����$� #����5��z�ڙ���r�=q�0r��ՙ�R�X�cPƐ��c�>��h
�i`��K{��\a(����h�P�L-��K�.\h���mQ�r%c�6�L���]��JV��}�����8�3M����u�{����?��%��Zgs_��1�$W�t��8���%��#�\�}w99�����4�g2�/QMUw��˯ieL�ꊳpg�ȉ�U~�V�l>�/]�.6��v��I7�)���Pz��eqb+8��pU�>!ڷ�U��{=ۛ�����Ը���a�$�/�T{��8��u��{x2*/j��$��L����2��=u.r��e�'��*�>���E����!'LHVA��H������8�nV�_�E�K�kf���h�E>.�K��r~���,٭�pz�����C�Fw��J��a'��/KK�,r�C��
��w�2���^����Р�	�Зb)�R��9,μ���0�˕{W��Ո��@ʭ�ƥ���E&�wV�1<����	Z�f�d�+�z#�9����O�z�!��lSC���
>5�ŋl-vW�좼fgv�$a�^?\��ږ�>��M8�����{d��=۾�!�1x��㤟0�{A���s���>��Pۨ��ښ��qn�ɯA��L�d��Y��1OI��ޜ�B�lX�O  �d����l#1#���֝����:D�t�i0��i����r�qڞ�w�k;6DԮ�]u�{8�9�|v�Ǎ;c����(VX�K���=hF)�������ŤKwks�@�ʙ!QO]�,�j�6��GA�/&Ϟ"wm7�����w0�>5&`�90(U�+�EA�ͮY����G۠�{� ���2n���v�+��Sԝ׾��}���6y�I�G'Z.[�~A���	��6�^�Jl�&[Rb��%9?+�MsMB�ݹ��{�ȍwtP�P���� ����Ш0^2��!�]M�V�G�c|+�*I_$߶��ٍ<��F�sߒh��<s�f�{������Z�-J�zbC�`j��:g�!�sݮ�^�wk��XG��e
:y�r[��.��v|^���PT��tvm��%**)W
{�cy]9gWs|tOO�TK7�&LJ��uA��@����`�̅��)|��'A�r���%�
���&��N���,׺^�{����'������1�E91����W�L�ܧ�����4%�=֋��C�K�[�C��N�O1YY:��v4���f�kfe�5�B�+gMg�߀˛6s<�皤�89�u����֬8�G�l��B�*�I�K�(�y�vq����"I%���;5�ܨ��+�5��;����3�~�D����1�e������W��d��Y�x9!�X���,`��EoP�M�IavI�2�����B�����_{�k�,�B����g�E��<Bj���4���㼼vЗ��XhM�%�ɾڗ�P�ⅩWQ�F'�`�M��1K����u�\�J4x� A�Hc�Ā����|~*���fU��Ɵ_��D(�/_0�
�%D�$;��2�ɮ���l�ç�<2�WW��3[c�N�]5B����瀖e)�L�u�}hL�<.�#
4t��/�Ɓ~\G�NCdל�����A����~WC�9����*3����ʢ��R�ݟg1��f!m`[#'���-�$p�Ǆl������]Χ.R��$����s
x:�]�L��Z�1������ժwl�6F�?ZOp#52��pZ���=DJQ]���[ϰ<��GR�S� в�*��*�[��T`�-�5f���Q�Q�:=�0��\A�ᇱ�H
�r�bZ�ei��*!r���Z��Q�����
`��:�me��UTuT��*�����M�������N�o��,�jݣ�v��}���b�1&���ټ�"9t��&��L��үa��R�^�A��5,�o3��c�tm J��oe�BvQ�G�#F��]�F�X�"�J�+�b%֩�o ����ܣOY]�=�a�7��a�}[>$��]�h�W5�1hNw@c�\���G�*�%vb���>T��eK)OZ��f�3g/�<�E�b�>�p�=+��4���]_�2��l��� ���ih;7k+gF�o#�>�l�
k�>B�X�f��|����[�!����-k:��,ҳ|�n��k��S�����p͊��S	cD,z�s��Q��-*bgh�����i���|cڣ0<�|&��R�3�E��ͻ�����Ю��gr�#�����@z)@ֺ�:�ۥ-��}�����O�N>n��e��ݫ�:���]G�-ot�̤��-dc�:?6	XǺq��v�����9Pi��Id�o(��b!���]frr֮�E.��D����F�J�B��4�a�B�<���L����W+b����1+���JMtQ�jo̮��\۲z�dΟ|�Ƞ�hj�3(!��*k�2��+̱+8�Օ�I��[�UAT�2�2302��#J�"���Z"(��M�����5&�
�Z5�X8ffed��X6�Rjs����:ۋo}۫�:��\�sa&�۝I������������t��9/�{�V�O�D�����@��>TA�^��O.��q�iE�{�u=��D�,��ޘ��C��O�*�R�V�h��[w���A�w/!��^8}0��fY�uҼ�v���ZF5�����fE�a�������ص�]\����[����3̗���C�6}@��{����I~�tDxs`KYtǟ�0ߐ��wtt�T]QcW>�6���Ha�ꆍ��|�wt�%O�Kn������w��},T��]`Hs�b�iq�\�K�a��l�7ƌ=���0 C;z:� ��BUf:ź���!�9��v�l*�|���W����I:���'?vAL�����}��K!
K%ڵ��/��������Ȟk����$7v�*eD�<����g���,�	��$�l�\�s?~�G�/Ot�[]�����-5�"�:Ibk^��S�c3=�n�7$���\u�V�sjb0� Ն�#	��w;�M�ok���-�su��Q�+�hj�}�8���7�颼������W�-3ʃB�����Y�ɪ���"�w�X�W���$��u��Ǽ��_p��;=ۣ�Q#�Ǐ׈��K���M^Q�9�6]5X4���O$EMuA�*Y��O2��W��?jD:��G��;�T�S{��}�ٯ
�#!��Pf�b��4Y^�U�sG��>A�N5������d�G��<z��`e��������qN^Hi����#"|C: B	Հ���U�v���T���g��'��?j�5@�o�����Z�Q>I��9چ�ऺQ�{��f-4�YG9�2}sYd����#}l�1Ͻ5�ʁ�.c�eeQ�
dК*I�b\ஒf�f��<9�l8�.��u������uax�����LL�{�� M��8څ~v���u�s*�� t*A&�u����������ԍz����`�)�(]Z:>�z+�Z�m�}��9ЗkǺ�3�v����!JzjbWq�'e&KNfm�9q0E��>[kܰ�)�g��j���YĐ	�P�fۺ�f'�1��ݏUR��e;��~�����kz�?=/$��đ�9�u����.�����'��7�JC�[C�qD��e�e،�=�-�l_1���}5Zj9�x�D?�x���CO,-e�HWzr؃AV̯(C��G�+QU�/iZ��3`պd��
�3#��yW*�����a���[-M]ӢU���s�ba�Q�Ij�b���F�qi߾W�%ϬD�O�:t8F�l�qvy������F��4(�5qrt�yJ�	z��|�� x���bkd�]��1<@t48��~CqF��J�c�����<�̯z���<��^5��`��kX�zX�y8*���uv�͖�[��LYL=S�*KL�G��S(�>U�V�M�{�\ϭc�2
`m��|F����5�q�f���������iӆr�����w
X�,�S���0T��P�t��㴼C�a�!5x��8��|po?hK�?I�*d�ݬ�G�4^�fM9b2㲌O��N�6���mج�Bޠ=�v�$��đy����ڻ�y���̈́;y^=B��v�fh�ȋ^Ǵ<��+F��u���]o�)�0l{� Yϒ]$�*M!i���m5������+1"��H��E�SLt/��:�s�_0�HY䨓��
��
k���|�z\H�{������_y��s��v�X꥚���]"�1�Qs�9$��x{����K+�Z��,�6-:t���G���NmOg��C�R�(_�N���}Lz|Q�i�����軳3"��l�(�q�qe |��)��٬�/����{��Nb
�#��gm�1�|F	�$����g���{����=��$a�[�<I
!������&k���^�w
�ץ>~!�|`����!2�VQ�)�̂s Q��d��FX��d�_Aj�]5��!�P^�n���!v�#ѰȚ�����2��<GX�GL�D�NK4��2����o����Y*�^Mҕ���8����ud�ۻ73:]z#c�<��K y��ӄ�9�6�8�{[�9��ԟ�@r�{��4(����Pb�la���z���ҦiK�&tºYt,�v�q�)�M�r'�:0�2������XtK�?X<U��,Q�oO=[�!]��Մp
͋�;z%�V`�~¥��{�:p��+�*�OyP�1�zZD�KyE�l��p���BQ�}ɬ��1�]%�mʒ:���M$	:`)N�:I^��:��FC�y�^z}X�ʷ���Ӟp��r{}������i�B^!��s܉�3>�AQܸ��L[Ͷ�z[��u35oO��wŊQ��<�9q �BM��},y��9P� �)i�D���3H:^#֮.��%^�n�Ӟ-��"F�ł/"��V���B�qi=���b��6���b�޼�<8�y����&��R�Ϛ�VHwnV�7�˞>��Z��hÕv���ݓs-��o�4��Z��-��}�^vim8������K���ƢxƯ��A�ThJgy!X��������� �ҎW���kY iu�`\���sf�7�D�.k�V>>�ˈO(x��O��x���zu^������έD����ʐA��̥u�¯ 
]����yX�uW��<�xP(���3�ǆS:!2��~�w���<��I�?���l�Nu��u��d�u2������v<l�#1��v^E|�ͦ	��q�Qu�m�㮜�|���Nx+ޭ��a4P�;��v���}\G��E�=:�T�iR�#]��	�X-ON��ڹ��W���Xt)� �z�g�ei�N�x~"��
��7���b.�^:�e�|�d���l��C����e<��x�NU%�����<N�V}B�׳�I�%ڂ��o���<|㟞����eG@�����9��lT���Sj~{.�npw�!�;��m/B�{�]D��9��K�I7��$;�'Z��U^t����o�o1�kȄkH�&���&}kO�i��v򳽓k3�t�G�ǈ�v�x�-<FP#�29F�2ܼ��v�zO�u<p�q���Ӡ�4�<՟1�x�^�|���=����^1���9p�9��	9y��y���N� �7h��W���-����!#kf-���YN�:h��52��'h�ֈ
(��O=2�6G��c�sw���Bf�L�[z�8�Ei������ ��O����+�"����U8I1�փ9�
�*������%x�W&���B�f�m<�s; ��Sb�EWx�]ݞn<���9��m��t�	2�s��N!�{�z]��j���ޅ/��O84�[�DMs�;��v�P�_�5�W�����e;�_��Xl羥Qd�d{<���F�/��㼼h�[�oI&g��Ѱ����Ƌ�<X^zz��f&������^��:β�e?w0�+��I��VtĆrG������ac��=ۍ�WΣr��TT
IQ�,$;�0���������Y:��,"R�j��Py!�,Q�U]�j�9vo�p�k��kˎb�zX��ƴEA��XWe�nG��{:Oc4}kI#֨gF�j�����<��������W�ZNw�3N���J ��z:�)Lf#�`R���1m�������݅��c���9H���6}�ĕ��֒��4u�6\T�`ehҠ/-	5�\�6���.�f�kΈ��Kz��r><%k΂�*�r!w�0�MF�?�W%�n��+���Ǹ��讹��{��1�>#	�$f+յ���r���9��y�0巄�
Yw"`86��x�5���őٍr��E��+}�Ǫ��/��P�����~���Ʀp���+'s_���!ځ"�w7}�����פ\l2'��c͘o���v(p���X���ܼ=�XEe��K��la��
���5RU|餬����O��{y6*g\ta�09�sK�)q��:O��G;�%�ҪZrK���N�tCqQtfdq�u�Ŷ��V����	�A�.�����D�z�絾���[�� 8k�`�F	��p�n�����"̒v.dH�����$����s��Te���v�22��]6+�#߫��*>?�*�����ײm�`b�!��C@;�,g'�q�����V�H��h��?JGY��y�k%m��0t�m�I��,�Vs��𭓟��8eh��%7Wת�Ӆ��o±��3�^��R��L�;J�#�Es�eeF�4ڲq�јfdW���� J�T��o^чU���I�f��a���P��J��1���>ds��كb9���A7	z�dW�V��ȩ$o�|��N�WN��E;x>J���1	l��Mb7���k���E��]ew>�2�[μ�h�����3Wل�R��2T�St���%N���[�C��`�(X�'o4��X�c�V�孓�[j���6A���xD��8�i�J�v9|z^eԭ�Ⱥ�����օV `�<�xh8mS��n�����h9���ի��y��*^�i>RڛvuV������#����D��3�ӣ��ǵ�;U0u���G:���ʠd��n�Ώ�=3�wK�.�0����$KS.ӑŧH�]�ك�m�Tu��H�x��MM��_�;N�*h��K���S=q�*yJ��J�WӦ�|i4�_��E^r����A��"+47Rg��%y�Ysx�MZ�4�5D�� ^�vصM�ϠGy�GD��XZ�x�t�
_s;c�yw�m:�S
�VU�Ն���Թ�jf�|�J�jٮ�zu��&:��ԕ�WMWxN�=����M���'M�NU2X)�)i�P)*֒�R�v���S�k;�׌��7d��V��m��ڤҦ.l\��#!���ż���(ܛl���6�K��RďX�‥�=r�g�nK�*t��s�Y�u�U��`Q�aZ��Vj��(�sֱ�e���5�aafYe�kXLDd��֒�њ�*��0(������j�k��e�e�ae���I&ٛf���°�)�01���)�*r�1��ͧ-e��amdZ�2�w���e�A�j�,�,��jh4�RdVe�������o���pL��}X�=�l�J�5�@Г�y\8���V�w�������@��q8�!�5�s܉�=!�_/+�[�D9~�v�xyQx��+^�}�.�.��|UY�)kͩ��w�:d�f�"��J��.!%���<u�ib��q��nw���`�� W��>y�*
�z<��%�맩>�~�[�	�� ��Lи�D�(i� ��a%�p�"�~�M�k����*]_����W� ���U�4��ї���� ����U�
,�ˁ�׌�5����˙w�|h�c���]Z$q�Fsn���vT)0�3XL�����4�̰��R�yb]hx��]�-�x�y��5��qg��vx���q�)3�*��n�g���6��xk$�of��öd�Z��M�=��7�+,���Vې���͠���iT}Yέ=f�D_DV_oR��J�Խ�BZ����ٱ����[ַ�)/��d2��>�3�&6:�
-\9}1Ү���O�v������׳��g[�ڄ���NPW�W�Z��mh�����:�υXb��ж&BX���o��8j�Su���9�\w����g�j��B�DZ�â)�Qz,ɾ-x� ]{&-�Jᄰ���6F�,!��5���
%Ze�zO}�Yg||,�k����z����@�tv6��3��,�8�H��wf��^��?&A�Ó�\y:�U��!�TG����8�6
"Ǘŧ�A���,�p����(ph�w묾<~d�N!�t����㥞^�������?o��h�hZ�Ğ����	`1V:l����`�/5��9�h�
&��e�/u��3�����Cے�c��b	ҧyr^�u8�:3d���1#xv-��5 r��v-�$)A�J�}�;���~�����ꎕ�.e�ќ�R��Q�"_��m����a✉��o>3u��-c�Zo�n<qe�v����hFR�=�S��F�
�1o!t�-3�=�ۺ�ةp��Jgf��1��$�.����[�/,v!v���E�����*���I�Ϸ��8Ͻoe�S�������"�m��C��n.\���3�c��������bj���ag�ib�¶����O\c"�h�!5v�6z�S9����P{�@+�)
c]�&�Vt�2�6r6���Y����
��]�i�U�:�%F%����5�.�Z0��`�P��)Lf׺-\.�CH�&<N���3�r�(So�5��7���H�=+749�-��;�z�<����loRԎ޲�
���\�R]��K*������u��{������Zec�!.'��6p��ش�춌���S�}�</��#Q}�� E)_���u��G9]�SM���� 1�#�L���kt�<}ꋝ��O'�ܰ��P��&�C�SqKP�H�=�1C���)X�Ϡqx���]_�ezջ�v����s*n�/*�q'WUq[+N&�|�e���^*����0j���!1U�&P�Qg�RZ��V ��[�vu�=ƦM׈�������E�G;��O�e��!}������3�w��0��ے<��Ь��*,U!�Ia�� ���r�#Mw��Y� ��%��oSO32������r��	|��\n������U�`3��/��>ÇU��]�G`�( �*3v����������QO����mL}�.t;�	*�Ŷ�8�o�/%d�zI�܎~U1�۱1�X�o�F�a7>�]"jw���w..� 2��3.8_�(����L	��<xS޸ ��o��?oN�ZIx>c�����㷌:"�I}�r��]�{�oO!X ���ݲ(C�0���]~�цnT�Bm :���E��3�p���,�=�|Fܹ�D�v����{ؽ����xFZ�j
�%��&:Isqs��Fyԕǅ�I���I�t��w��I�H�<B��#�k~�z����R��^7a�ȑ��"��f��K5<�@����	�^WO�_�z������h���DP}���k�	S�D?q^VU�(�������Y�3QH{�[�Ǭ���O2��:��(S���d�v^	�����T�ov<���������ױP�7�0�ݷ����RtrP�16���W�U?g��
�ߪ�q�,�E��t�.!9"�(o����\�w��4G�����鮭<l��L?����8�����P�������7�GG��8O3^��;�&@���2M�]�~���EZ�T5
v�4���[9E�5���{��*#԰���!v���yada���v^X����M��pg�U�����N?hzxHq�+��m`V�_�v	�4��Ŵ2c&�q�U�<�A���$��f���K��p"����slQ���+ dz�{��s�jy�g�oV�P�i�:/e��@��t3	�]4/T!�y��:zT��҂_h��ԁ����VK�*�{^��#��<3�����s+<%�:'�bz*�E3Fi-�$%wm�U���@М�5�~ܕu%�gHo\��z�ww$����m��F�T�.pV]F�QW^� �~)��Ґ�Uݻ�3{�:�&����c��v
d1�ǠX�m
v�Ə�c8�/5B�СP"�|�xo�_B���N�и���i�^�(����T�s�
.����^R��_Ƣ]�Tsəbf�Z[��53��0M�['�Ze.!yю�.����}����5ND�Ʒ���Du_��x$� ��͕\��	緲�\m�Y���up朩�V�&�?�>�y��|{Q�췦Z��̔�]o��D#�{��v��5�8�4=F��pp�ac�x�p��2ѽ0 ��\�M�U+.�`L4o�b�uHۅ-�R��<rKFf+_�)�z�8�G��Y2�e,9k�n+6�F��p8�v��}nC�5���x��|�׻��{vH�Sq��I_zji��g���_L]7.��G���c�Adq����{{ޮřlq�S��vI&�*Θ�^Z[E(�U�-������ۨ3ʵTB�%D�#/7x��^�o��~�k�a�ף��
L����B��j
me㶸�8�B���ut��K�=f�:vn\6p��Cx�c��μ�� ���p�ڃ|X�Қ����?�=4M��T=�9Y���"ϼǑ(�����l��R�&%�q�&
����h�3w2h�cť���D�/�ϣz\�^7;|*���Vww"=z�\A��ç���#��U �s.n�/���Zq�&�O��p�C��ſ���G,ȹR},9m����I>��Gn��/Sj`�7f�[���A*�Y��J��H�x�;�{;�>��up�bJR*
�Yȥ�ً�E\��d�{3ZI}��沾��Y����s�*�6�V;���9~�Y$�<���J:/�EG�V�zE��`��e1�y����L����~�K�����H]]a�B]Ô�`�TX{�{�[ſ[�� ��ܾ~��6Iʎ�3䆱�K�c� �{5=^�v��^O7�q��C�!�a�L�������U�ɶ�g�=�1$�/�"���A�Y	��\Fg=-"D������.�q
I>|���:
zvS�㷌aa�H�[�~�>w�y��L��԰][�Bc�!��]�ˁ��'mL�xJ9� ť޴X"�|G#]?r$:О�R\��{{�ݿa�X�G×"D�X~�a׾01��b�9q&U����u��D�\���6ӥu�����c�����\�p	�����Gaђ�aY�N�gNT��vY;r��c����[�Q��#���/um�o������7��r%}x�x��}#�u>wox\��ꋍ�7FDPP:��H�Ba�+}A�n����o�Y��*/#���Ls
�&%H52�&��1݊%�t����Ӭ	X�E���^P�֔`�a���G�]���p�G���a�Z���^�;�ӥC�8��r��<������dz`�8�5���Rդ<l�*A����h��#%���S2'�:[FL*���B+�lu�r�qONa����uy?o�N6{�ja�0�k�P�*�0�/�v�N�w����JM|D�K��$ʟx+˥s&|vB�uF�oa�!�'�sY3�9�1�f�/�bc���Ҫ�sO��|n^cV/[���7.}๰x�)x����,�Z0����b�m�v��B��-N\ ��ȵ�+�s�}��}X�^��$��L�E�G(K7�y�C��f;S���N9Re�I��{Y:�]��]M�8��h�ns���1)�k�T�����&UՆp�n��P���,/�v�vt֓bADśl8�]�B4TO���u;�%�����´��L����ycpkU��؇�n�Q.V,˭((���FO�kPf�q:Zص���nF��y��5��8 �7�9�[V��hd�/uq���:�{ʲNu.wLWyK$�w1t�3b�[(�t��:|d� �Y����Sw��'C:��ٷ� �;5��Ǒ��{��6B����N��zF�&l \��y%l�3G�zc�w)f�Q����W4x�,|�0ed܈�m�㊓���\��t�^�k�΂��w!8���We�^GE�˗����[��R�!wm剴�*�V��]��4xS�&s�7;|G�^�]�����r�ɝH7W�o*pt�O*WX�b��wf�fFe5eɬ�+��Jp�p�G)�7�j�J�c��_2x�lv��V�7jF �`��;�i���M�μ��M'r3z��[IQ�)׻V�iYZ��кJ�7oR�[��o`�Qڱ�BC]ba��QV�Ot<�ӛ6':w8Ƭ���|e�y�KD<є!\6���"8��X�Pfݞ\�-:&��.nV�$�]�ȋQ���"\����u& �s����U�OnT����f�n��D��5Y�k�e]�*����R�55ݭc����U&MKj	�56&du���d�VafE�dTDm���#VTVF1a�dfY�f$Mk}%d�̊w���2�̤�A���YF��-�ūaFQ�FA��m�U��ִj&����SUIm�F�6��FѫQf&N�m��D�F�a��̈�)r*5�Ɛ�l\�ƓQ�Ik�;Q��C0Q�X[Zܸ�G���8�a%6V��Q���_���o�����-!��i4-�2��JZъT�k��%��&,д� 2�c��
#"h<���D%�1嶼�30F�\й5>Ν��WTj��n,yI�"�࠮�t��$�k�_�Hk�CK���/:�r��4<�>z^"IW����k'_�x���	�#K�����D#ZC�4���Mt�f��F�~��%�!��'5�@����ش��#�;��^�|��Q�^��q�ó�ݩ���4t�f$/�(,�\9'Hּ��E����U�\�$ǥ�IX/�]{=�`���������d�h�v����Gơ�+���oܻg��0�3P�0��"`#�ό�h���^�9-��x�ͨ<(`V{�_`ooe-������둳I�ڣ{��fQm�B�#+*�O�t���2�]��\�۝���qBH͔��\I}�zt�x�!��1���x�i�*q��b�B��]��U�{����?dצ�g��~0Z�6e =K��rԲ�o�r��,CV� p 
��hr�]<=|`�c(�ow�E��m��x}�B��;THav����^#)�:����s���OP����[�b�0!
��\f���AJ�Toҫ{�	�ԥ>�� �x�5MW-�$`� �&�������ś����b����Vr����B����Tž�˞�~�B_A]X%Լ2�s<4&~�멒�
�q%H����c�z�>�H!�<����d:+N���,̺[�y=��,�؂�4Fҿ�Ň���x�Fߞ�	#�'0�J��W�4���
A�H=�]�VY�w�����^g����ISA`��1r�O���F�
�]���@S�C-��3�\x��G�路Km�2f�
b�*���bv[�G���񥵌���=:�C4�&�ZD=pd育���H�.̇}�v3�����&c���h#Z8p�ZD7�5���`xR�����X�Bσ\x�L�!�cҘ��y����WSqv)Mv�r^���;�h<���0*fƣ��~p�&_�6���K71o�o�n��d��A��D���Hq�1Qʎ�w99s���禃��i%��v}Ώd(3�a,4��v�9q�Ӄ|�����R�6s�*�|}C�����L��������=��7�����BtK���{W������K�du�B�urk��..\��u��M�dd/�=�C��Za�GdA���������BZ�&�O;�wwu�Hw�&���j�hnq�)�F�+������HrG���N�f�����LL��MԊ�.�zr�×0����&e2��_�ƹ�@�ۧ��>�ˮ�[	
�=k�#�O��*杞�
�����g�Qd��G�9�!��mK�ꙋ}o��/K.��Ϛ���EI�=�� ���h���|&D&����#ԏ�BE7C���B�58��������������z#HU/9x�-��������d�5�g!��e^{��/<zr�4��Dx�H��.:`и�%]�7J\�t?:�T��1���O� ���E��x�h�T]^�o�4���i�'֬���=]>Aߦ�S,D'-���Jt뽝Џn2q�41#�RY��9D׃,Y�ӓ"�f��6�}�<�����t�>����!N�����υu�w�hz�&O'�_ma�t���X�_J�ZZ4���ח��6�h��7	��x��	����Ki�C�
c�#^$��q�U�������xY����6{���PX�(hA��a�qq1���1�W#���N.�@ޑS>��1�R�\vCBݾ�b����J��a Beg{D�J������☸�`]f�+��� �| J��Ŋzw+Մa|��G�p�EϦBx��e�*O<�v-��%��Z� ��)OML	����E$��3�:�^���{����9V������	�3Z.���XE��M���eN������3a,���H������$����;w�^o��D�	�GgL<e�Er�y�iEU��p7o|�Ӧ��z,���5Ӿ�"�^W����u�<�=S���V�M���Mz5������;3��/�](���y��v-12�L�fS��lI�}�Լ�I�A=��p��!|�������*Ș3�(�9w팽Ε>��|�L&�� �Q]��)M�g�r�8@�)��]�1��3ʗ	��ow�}�h(I|<* kl,V��q�����Բ�xn�>���{�k��~b�
�9��|f�E�~qC^���m��ŹP�x/$L)}��3z�LPf���l�n�^��RUW;>s����R�Df�fAL�}�����������y^�b�,`��zk�Q����Y��$�X��BM��ˎV�k�j��0!���Fچ��&���8_Y	�Qj�K��NH���:b����xEK��[��౅�=؜�ʿ�3������x�V�!Lk�I5
���v���C��
;b��>��n&gU�+]jN=喇�d�8�z��#�+#W���>�`���*�s�G(q�.2oL��v$*�[���{яt$�0cf�`_/{��!�S�Bb�R��E[�"���wZT|����k��ua|-Lh�lZ�&��v������zQ��,������k���X�f!.'��/��µ[���Y�jώ�/�D�fxxB6���j;2��<>�Ux`�ψ��_i%?Q����qn�\U���iJ�6��a�a���t�8��jR$ig�h��X�_{۴=�A,"rIQ�/���L$0���\O�V��{��g� �qgO���ZV�S�D�Rr�f.�k�$�Kהj�X����E����j$�<��خ�(�@)��
�ys�Pz����݆a�����;-�B���dK�;ݝ������urS�����\*�R�C�rL9��^��v�]��ҳy�G]��6D��3��N������5�s�����߽��|��˛���9��γk��jB�>:�K��la��V������ ]�Hz��ʽ�������d��b5
��2�O�����P�>�#�t>e=�z�PhS���8o���c>�ݱF�#�&���A�z���!<{ʇ!�6TZ[Ʒ3���$�<+��Ѷp�!C��t���xͼ���snS�i���=���w񡢐�`�U2�}�*������0HL��q���+�Ȁ?j���E�g!<FЗ=��뽕X�]$K\َ.*�ź�uGr��ɝ�h� =z>�Z&�6����gOhUꇍ9��ד8F��.D�x�v积���oO���!����li$iç�[�ʾv���.��m�Y"6�Ƥ!��a�%���hX��I��ձΑx��w����4UnI�7��ms�&��i�2J#�I�������G�s@VP�'K�뺰p��p�H>4�J \��E�~���>X��	Pt�!�r~P�֔Fx�ڈ���nowA�kI~d�F+Af�8_oO��M5��Z��[��w{�e/#y6>3��;��)<h��l�ﳷ�A�5i)��C��-q�U����d�R�p�:�� (��M
��<�ؗ3�XvL;�k�iŸ_4^�V�w����O(��ž.c�%-&+"�p-%q��H�yP�h�\��PzmNLl���Y6�!]�^5�MtX�7��>�u�CPC��¢å��#ME���JZ��"�[ͧ�L�T7Z+��o�Fe��(Yȑ�6x�o����x���y���(:|oEl-f�^�
�1C4��wZ�ÅN:�
ʼ�T��,/�ˏn;Y}k�GH���S�lIG!��)$U�=`�Y����J�K�'E��6��Z�aDN5L>�S����2�uʔ�S/�s�^y�4�	����d�1i$e�N�;>0�W1�Xж��-f]����z1��QD�=��NK~!�i15�AP�\��hJ��4�L��
�A�&1�gس>5��B��4=��s����4���0����3�h�4-a��=z�
��+ۦ:�f�D�>3#�d���Zj�v�1o"z�v�uF�j�a�W!�)Ș㼸�owT]��:[)?VS���]#��T99{+����qf���"+5��C[��d肾�k4`#B�|���f+������XW(��Je��Ȼ�8]����f�jX�+��e6��mp5�V3K�r�ü<LV<��%E}�8���d��띦gc��ս�m�Fx��>�G@��j���[\�ӿ�>��HBPT����(�'��d�k�ɽ�B��
�6(٥��\m�!p�n��a�Cu�bCxp\�l�����l�c�Lt�4�i�yD��j���ADKefu�J�tͣHp����U�� ʶ7��_D�gKʜ���XmQ��rm&�t%Xf�Y��)0y4��
\a9ɬD����Aιmꊗ��z�u�գm�c5�+,}������;��A��N�1of!Dl� v�T�)�A��"ܡD,��ANvȎ�)2�J��:��@_LT(-2i�����E�8g^m�c������;ORҜB���GvMpӬ�\���O�q9;�lDu$��p�P��s�Z��Uf����s6ٶLM�0�b��`�9/�tsjj��VڝDHM��\��.�&�q�@�ɶw3o;Qk�υt@I�1�.F�ox����n�h��T_f��S5���"@�o��M�
X;)w�c���&��SmG /yuA-)!Œ�l8�<�։`�lȾ�ۃr�}'D�ci(�ގ�nM͠�]r�|�S�.fmr�$f�2��2e�����xҗZ��y@<�2�&"��X�6(`!]a�;��1o7{&�于�a,��I��Ԟ#��y�;M9�A��r���˽)VC�����)�5Hx��hx宮�Dt݌,�D�]Dt�%�_E�m�%�R�7B�Q�˪���6�}�.Q9�L�'QM�)������i�I��k�r�P�	���ͫ�Ҏ��
�E�~��[�̮-kQ� ��X�o��JM�p)��Ԇ���+Z��Q�-Q���[��Mma�MS��2�s1��7�&6�$٩��*�m��
"�VI�V�`�e�2�S�Y�Vf�+A�f�Z�f9��`VI��QYAM��E:̪�6�m�mDlFLŬ2I`afXffe�E���*�Օ��ri��$�Y�QTF�kS��cQ�0H՚���Vf6YU15��JM�T�%VY3%��#�����	* ,�*�kYS:�'{(����|�a�:̦��VAAKC0Z����q�"����bbJ(�X�T�9%9a���)��N1N����&�j�ՕN[ΪI�ʈ�eT�V��(��h¨��0*7�
h��lƭMm�j�ͳA���5j5[FV��S��kT�噘��A0�	��	$��KGP�;"u}u��J���/!��:�r��w-�#)A�Lr73������!@��^�]��-
�
*d��^�����c�}=�{-�0m�=\�կ���P$0�;Xr�5���8����º����)���Z����[E�XZ����yvq^󊟖u^UҺ	���鉍3*�W�ŒU���΍���w��&�$y]�t>��G��g��P�s��G�y�Q< aU,L�uc�pTe���_�����CS��g1�(�;�@R�Q9�|��c����z���qI9�ǨA`��<8\4��8Q�X*����_��z��}��}�Ȩ2��f`O�D��s����$�,�~�u:@�1�Ť&�˦�ť�H�L���=j�az�o�'���83��y�G�b�e6���^�3���8ܲ+)n�Ŗz�:���}���njU&���@�N�3���g98	2sN�9���g}�xX�����5���!�.!�GSHLO�yr��[���W���HR<W�xឧ׏J��y�����M����Z��LUj/?��A<��L�m�w��KI-%�/��p�$�~І��y/דHq�'-��ygL���'��a�C��P����/�UJ`mHp
�M�,�Qr�Q���`]�鶩�R�z��H��ܽ��Y����z�#����tz���}�c3O�st�����w{�'���e�}�V �}b+=�z"�x��7��+ܒ�|\��H�,��66�����:
zvS��{�eNV+;73��>�MF�G�Q'L	
�=k�*s����A���9wU�d��W���v.�}�,^ͥy~��g���x�S��t=
� u����g��&�31>ںOJ��RV�r(�7�Eo���yNVy_NLVC��G�o ��S�'�߫����s���y<"��U�ւ5�|g ��fj���j�Yo�͔�\�ɸy[7�gySB���&^!���$�g�J��~�v�H�R�^7Hq��.><n�n����0Ye�QǾo��)w�
>�X���4��@�5���
�-�jI�9�:����>�*�BEZ�3�}��@x�Y3�,�s�g���>�a�\K�H@���h���z|��i�h��[��\[=1}N%LPw2��ﺣ�<x����R�#�]�xK�&����4|;d��S,y��J��.��9b]X'���헙��!-Y^�jqc�Y� 4�]]
L�,jv���ќZϹ�f,���ͱJD��s�&��╮{G��%,Ƹ�9��Ŏ%�Q���7�*��"F��F�h/��]�dɺ�t:6�nqd����`�*�����:M�dq@[��h�ʼN/s����oh�jd�36o=^��k��g�w=v)�95�
�x����j�H����`[ؓ��pY�^^����rg�h^o����n�G�
��=���gᓷX,��A�,�,�"v��[A��gw%dhW����brL`aX1��˱�������n�Ӯ`3[|/U�e�hp���,�m�)�W�bv&4j�����֣�����P��5�����V?lT��z#jĵ��"F���ݩ��Kr��u��_JŻ��Nr��3e��)�ů295n�@(Eq���M���%��#$�,>�R��o#����i�F�����/K��Ęw7j��X�r���弎��E��� ����p�W�:8�F�:���lTfI������q�&�[f�g2K[�ss�A�^;��IF)�X;V��ɴ]k�i�@��l�ꁗr��յ����.-v~�\������ޝ�Ӵ�����>O4��#�E�i���t��9ܴ�n.��	y��LV�(�Mn֫ל�8O�0��ʩ��Y'�^�ӊ���F.ƹ�nXx��E�=�(��ᦸŧL���N�ܺe�������{)�N;
.���-m�{�[�쵛$��� K�1$�'ᶛ=ѣ�`�'p;����O9�`7ձJ�:&5����9}&瑋`��8[�+��0����MG^�0��Ck�xWM�q�}+�8rK��	�Ԫ��3=x5Q�[�+���S����5w�m�����gPW�B�r,\jh	83n'���D�f$1��Bm���X����F"u�����d�ЏsUW��]렒�*�3&���8�^�����a���UF�����'B��yU���^�\-u��7Z���u�����&�7P^���f�2��GQ�8�t�8��w�ks�0���o>��,9QLy���:���M��NJJ ��޽�p�*�*����<D�r�gk/i�3�[����V��U[�)���Y�ͪ���P{��\Q���h�/(^�R��p�aٸޝ�I�
`���������4Y�Y�,�)�״u�S�'%ri���P�5�59+S���g������f�+)�E���gH�o5�0���w��)��+jLI������3���E��4���=q��{��X��D���A8�~��LmR�z![ ��c���bҹTç,5�P�-��)��V/5��U5�Ą����Yo�kɰ]mi4�Y�Mc�̝�������I(ƌP�7��J�w��Q�C���~��pM���:�j�x�L�sl�w7j��SE��˸�+#M+��Y����j)�uղ�L�=pvsf(��4u�V�zd�/��C�:p*��kb�ꡯܵwv��>��P�`	��8�Y�	�\�Q\B�5�a��'ڰbB2l�i���h�9���n�\OrykHޑ6# ��Aqy��SMp�.�oD�odY��l�89=�Y|J{8\��[��+�N�tXŖz�.�sڎ�:�F�u�4w��%{��
r�{(�;oF����J�RS$GNiF` �Oc�b��AD�����N��ǌ�J@\�0��I�Arp1`ȭG(��h��r�s���`U�Ѯ�2/�<�u����v%��X��1��]������ofZ�=��L�Ger�h=�U�1^º�y�f����1�tO��f:v��Ɯ#�{f^o�xrY�q�9�U�v��
��ps�{����*�"yߡ�����i���o_m���YI�Y��E�ꐱ-�*�6�f�iI~B�"Ѝ��/ȅu��D�Q`�<�sS��`�Lޤ��mV��J���x<kq@/
�b,�s�%k{�7�[���� A�n�6��1L�m��yOptk�9V�$���R�蠔ԋnuƒNAq4b@]!4���I;51<&������$a�8�=�N�bUb�܍ֲ�e�x��ۓF��E7���]wq�B�鼉�&KPCӼ\���'s|l��O�h����0K�a����E�U�O<��*�M�w��JZ�n�Q	3,¬O�d�T�8�1�P7:�����RxOWƦ�ڐp
�O��6���!����N腔3=�1��%8n˘M�;��N�4A���ms���� �y�+{w,�"ݬ{��V>����IV�z�C0o���S�F�h�s6Иt˻Tp�T����}�e	�	J�������K�1�N�cu�y*�L8ɩ��h�
�5��P��[Z��iky�.�m���#����n�δt������}��bq��P\�>�Vꙻ���:�qa�@����=�f�p9T%R4zVk��"�e2��];̢��㬳u!u���e=�vf�VBj H�)���s&�t�%	&�F��³2��ۃ%s;.-�Ԯ	Ÿ2�m���зv.FP|�����V�*�a��E����C�A�L�9��
�U.�A)�6��MRٛ��w�[V��O'>)��Db�h)�����.�V����m� ]�p��0LF����6U����.oV�S�h�q�-X޻/��!r�}��>��&<���i��.�u�u�F�ɣ.�wAG�缸hΓ�:o��$��D�-g[�:w�ή��TT=;N.�if^���x�<	'@Ak��*홸�@,[i&���xNz�
Hp��K��WT,����{�-)�j]2�;�*��� ܜ�9M긡p�-����"������x�|{�"���-j5���T	�u�H���3�!,s�/\��gv���b�Z7Kqi$��m��i=����2n����˂���${��ޕ�u��X]�-��z�s�VwE�eZn�l����R�T],𻎱u#Y��k0I;""m�.͡�\�(v_�3c�w�]�[��&��l�6��X�1�h�$r"Ru�����+�����qN}�;T��0`�`_v�(X:��e mX['Z�����(��3�k�#V��DDUI:���S��beT���$Y��K�(u4Ph��llU&�`�4Q\N����ڠ2�X:*�AT�d�CN�o	��2hf(��ͱL��������
Z����X;F��;ڵ&�䴖��AB��
JiMf4�C�jrB�!��!�&���ɨ)����Hd�6bN�)�L�iL$ZslDP4BҶ�ȡ�r@�  �	 aG��R�hk��μ�Vi���tڙG0�3���d�ÎErv�I8*��4M�w�HF3��m;�/��9����TTu�g}ƫi�:��P�<��q�/�$V�S�Id*��"܌ł^�T���W:�°Q�,����[�r$UU�Z9�N������X��.e>��{+�E�.�d���Zq�M����5��L,6��a��[�x����6������k���$ 7�÷1�;q&4mx9KxWN��������iz���#;L��j4qȬ�g�����m��J�x�p
���؎��1󺔼�]�7Nz��|L������sVZ,R�R�q��Tґ�_ԛB�~%v_�ON���[�)���Hrff.���H�}�C;��#<��F�T"��kw7y��(Y/�]W�f����ݚ����N+�p&Ld#q\z�*���3�F/�F��qкp��2�ߪ�	����2�l^>�v�������&n��o�K�뎫����k�H�2��b�F��V9��yw��>]�'���Ɩ׫v-�$�9_\F�N(��ע7+zt�~��E��	� �܁��
o�:�T�u���O��Z-��U<��~[�qK��i��/yvCQ�A��P��L9�#hE��%j�cw�U���eO��7)ʺfN�gSu󧺶+�b��%3�IH	�̒Q3џ�9���&���;��0s^'˖�Q紛�uٷ�n4����N���5ve��T�B]k7��i�2M�l��'SX�B�؉�9�HEE��P}��,���oB�a$�a`�o�(���b�ߣ�}E����8�����^����y7e����qW�6/F���*����(�!����l®0/�a�}�#5�-.�vE��K0#�]��t���7���:��y�4�]nagBt��S4�LHw��۩�x=��h���e�p��[9�J���1y֫6b��b��i�3��p�O���R��OK�Ҿr7���1��=�H�/{�v�W��������q:�\��G6����u�=aT��غ�Z��`�+m��[ڻ*����
j�Ȋ�����
��i0��^�&4��h�(�+&�eWZC&���Ua��M�/�ol�"�&��Nj����K�S����%V���^q��z�;ֹĸj�29d�T.�2��[�0g�ߢ.u���W Mq��"����獞9}'���,��M�۶I���&��=&��RlS�}t+R��~�D�K� �{�y�/v�A�5��xh����keg]eK��v@�r�,��2�g,s��ǈ��^l_:��bn;a��5̀Q�\������9���3�q���yҾ*�J���F��&��p8�ȹ�^,U�z
��U�/��;�xrn7�$��-:�35ч���5wr�!*�p��
&�#V��db�JM������=J9�lf�4+�pl���AjlXd8��V0��5�]εm�{՗7������T0v�5Ѭ$�*���S���zKM㉾�5��zvN�����9���桭�"U�f�Y��P�Ycws�r\����=l�ZPZ��fiQP��>흗���Ĝ�8��S��b��N�h7e\XOK	��|�t�����AP*KM@�+i���۬��I���N9!�#rC�ۄ)w�9\��E*S-Sɥ#�Cď1k�r��Zt�˛��s�A�;�yw�^a%{ݻ��}~��֤�j��T1�`��F{F�`�$�ߛ�U`�SW���VԢ�&\��X3^�q����\�j�qq���6�m�GU;��h�ڡ=�pYS}��>�3e�)���jyST���ڊ�sN�_���ҽ$}c8WB�'zN�oV윺�˒W��:M@f<�@UxMQ�t��Pe]���GƬ+�=����7��i���>J���R��g�4M�6�a���v�.����9�p�<�=���kjK"#�ǻ}S����lu�b�I\���fn�ki���ɸ��)6�˓פ��ɓ'��5����]
P �w:1�hJ3���Su�KM��jBm$��'�u�W&w�~���|���q��#'4cI�k9�m�#��:�ێ�Ns�u!���	Q�%q� .F}:�J�b�9נ�H�ߩ���5�L�f�b'p�FFmK��|rӋ���P��0K�с�`m�/'k���i��B���kD��lk�tl��"%��wω}g�#1c���k.��#h�Ξt��P��f-�9|z_g����ަ׹J�֝,��;1��b�	�vLF���sT�U���<��MqK�TlN�v7"�Y��MU�C솞I�UƤwb�O&٫e�P��WI[��8M�f��k��o�=y�b�X˿f�B����I����&j:��k׷~�����S.�>���|�Xq1�h��CΛV&�//@7��eo�3$�[c=F���'
i��|�z+��-��K7 G]V]�ݺv�ι�]�j�E����6��]glW$Z�^�'`��/��Xں���8N�(��u�8�Pt�H���`2��or�f�]^����o@�(�йD�#--'U�{t'��΋J/	�M둮R�G������\�HP2�5�Sz��EY������,�B��F�ˑ��%���P'Y�*�k%�-�͞���5;&�t�\�BQŵ�������GDÑ�������@��\eF#~[R���TnV�cy���Wb�o\���DmM��;�w�I��UlR�R�h1��S���U�Ds��	�#�פ�N���DjT�y}��ϴ",�n%� %=����G"3J��(�GW_����E����;���z^{5�.�є�K!���gb��d;�0�b�Ukt�0]��f�3�BݘnC\o:t;p�]r��ˢ׻�q���֙.f�M���.8��îo!Pftd���T��w��%��r�i����|\)�}��q�O�PUtyw!u0t^4��V��6�&�]���!��Tw�����R�{ϙk�w�͵�T��+�I�3y'��m4�wҮ1�������U�@c�����C<n���m9j�u��lk�W����������4�����Uh�h#�3����QĹ�����DV�#{�]/o;�$B�k##j1�>�dw�\��s����%t��u������r��Z��x(Uf�oe�2�f�o�%W�7�Ge�;eI�����ܐ�v�:�C#+��KS��������֛���t�W87���+6���,B�6`�	Ywګ�k��2q�\�	o�ܪ7����+�m��gH1��·�]�jJd�c�.K�Xë�S�W ��,R�;Έ��pT��iC-�:�\��0�4�SZa�y��2.�g���-��$̾ӗ���;/jZ3��:���d85w'��VQUF��Xy�
\P\_q�͍`��9�tB�s�Ֆ'�ϔ
�&vY8�m�Mޑ	F����W�㭥\DD�+��wl��U7�o���z�v�N�g�4��6��qA�I3�
��U�M1���=�j�e+:
͜�E�(d�:�y�t,c6��s�	�áu��l�z���I[ҷ���O:�v�I,��M�����`=��6�Z����Sc���:B�����\�e��i������+Q�kuEgV;���m�����i�3�Z�U�q�㸂��u&���3]�蘺���{c뚆i�H���Z+�'\(�>��~����]�x�G)��pfgo�(��SZ_��z �=�ۚ�)C�+6�֎�ҝv�ǁ�U�s.�/�E�;I��5�tI��d��T�xGV�۱��꧶4B-��N��X�\����]�����kH��K�n��a��W1s�����x�K���3�Z�1O�и�����[Q:
[ڹƆ�M��L�I-�f9w��:;�S�S)P3��ܚ�h��&q=�88���.�]?Ew���!�Zz�ȵ���"R�"D�)CC�&@��CK@P:��4�HHЅ-(�0��hG$��r�(�6�U�()�Z�( �B�(
i�2�i����)�iZv��)������Q��ȉriԅ��J�4�� �B��iȡu�%% QH�R�)H�Q�	 ��3���y�����͸�P�R|��9q�w�f�K�3T�5��!�����5W�F�^�*��v�����37�^g����4�c9`в���r��Yܛ+�]��*��u�t3�$��c<�0�q��oƷ�MR�F;W�]1�lrZ)&�f��꼻Z�S��V����;W�"*^�C)
3o�'����۩�����t�1g�7�4�/�Q�Y�i�a�0�u�x�Z8����O.r@�-�����m28�Ճ�
�ɄLG�%��r�](M���ߖ�RO9��m'~�7ԅ2��m��r+q����Vr�h���UY��M�g�۸�\�/o����`�\�0�w����J�&�&�P]܍)�N�㢷�M��.rt�*�A+
A��?v�q ׸Y��<��H\.��|f�>��iwo�ͬ:�s@�wT��ǧA�4\��{[s�F$�qv9��F�E�'D�.��nf����"�0\Z|DJIG�7b��x�X���<
� �%�L!Ƥ@��<�kd�l'qCn)�۸x���a,ũQSoos8s�8��0���w�nZP1�hv�-mt?#I��6��4lYy[;"�x���r��@�wma������ʅ��8�f���ef Rk)OL�&w[��;7�8�n9A}{��QU�������whܜ ���ݚ�xP�]�-򀝸���t�.j���$t������.����y*]�W�� V#�mC��8�
��K-+fuvh�sP��ܓq��E���P�<^V�Yma	%�l�j��l_F5`l6��.���G$1 �7Pȉ��rB�'YM��Jq=E��� _��!iٝ3�"�7���!�'�ŕ�޹!kz�Z<�����a�����?Q9o�Q���t~C��sv��i�O$�a�z�]��{R����|�����sP�^$�"�f�C܇MTmu{f�J�}RY�7�ؔx��{�A�"�uR�!{srܼ㌪��\r���ۙ{��⮄K�8��y&�E��mK
\����Ż$�(2A��}�PFWz��G�hx6x㻮���'��s|=�����2�%�"�m�ْ��A�rI� ʚ�N�\q� I�ϴg 4w�q�}_^g�`讲,���:k_n4��G"�dd���s��ޠ�8Tʾ��1��M��{��4�}$G�.��;ՙ����lq��nGz��su�Tz�d��w��-s�ֲ�i=�
�Ǐh�+_��К�/�$d��+��	;���kiaqYPy,�n1+���8*w�����}�d��=�ۜک��P'�1�:�V�U�u��<Ǳ̇ X�_���-Kl�$䵛�p�ѫ�T�V�u#]�Ͱ�lJL!��O�o��'5*���',e��3��vRaי�ֲ&��K���5i�-��`�?hQ̩�X�6�7����*|_I�GZ��hU�u���}���i��Q"94'�r���]���\�M���s'0�q����oR⸵���b�g53��\�,��
f;ΩD/;��E�`{^�V�&@)��J���MG,�ʳ�r�������N�㰻�zR��0�b�p��N��z֩1�kD���x��EG0�[�y�*�hnJ�;�
,,�5Lg@酏:� ������T:���Ļ3q#	�܀��b�'FT)K�q�����<����y"*j�jS��������|*i�]eH��}�P�"���1Ũ���qw�-BЬ&v���	~®A��}�}�߱�f�qܲ�Qy0�_\*u>q�<nt)�δ�f�F��ʴ�bm�ZiG;�0�^��p��x*7@�K��A���h�xzcA�\����r,�)��u��k��3�b�u���-������fXE�iqC��H]S^��l�}�o=su���ҍ�fR��q��;n/���q����=M�!�XedW8�>:&v�w�X�[�-��5�gE��Q3��Y̎s���	u(��d�UH�F��N�u�O;�KP)��u-<�C�}��Ƽ-�Ρ�pf:]}���1?j^����������횽���gjM�펶r�n�kS�-UC��\�#-���I%��;&��H�Ry��θ�ȨU��1��Ԗ�^%��`��ŉ�r)���nٷC��o���zD�u�)0H���i@{
�	w���=$:1<f�H��"EyP����AT�^�-�iSں�>QJ�Х��:ǽ��~3��K�r;um-%�uݗ:�w!\��vC�t��լ�ӱ�@��iL���z����Zzޫ����1���eˊ_�I��&I��^��E�6v�'�	�ڽ���N��eA������[t�j���jq���v+/���(�:ZLX�sS}M���a���n������:�V YdAM���������f�9��z���ڦ�
�����d}v�=�	��~Ft���t��S���$	;y�r�I�8�ݟ1����ˢ�Rǟi�=�<�q]=�t�X��uz�$�L����\���>@�=nOr���{3-�id;۳�#r^+�wi7}S�4B(xl��
��b�~`��n���#Gq<͔#3zw3N�zӾ�rd�7��hė VYK�q[7�$�]��uu���`��ڞ�ݶ��i6��M6��l�� ZOs��,��RJ�8�����8�޾NjniaW1ͼ�t�K	�{5AUvr8L\ԡ�����9U#�`�=P3z�\���.��yw�C5�El��g*wN�.ym��s�#�zx�scp�&���a�\U��d�|cD��z�^�w��peM����e���$�"8ׄ�FC3���XM�_4�X}ne[�t��/�����s��$7�Pa��Ÿ#5Ε�u�W}�X=2����n��Qz�F�u�
��T�pI���#���y�#��BF�+�7�Ax�k*Ca��&�y�X�;Q��F�f:��{� ���P��q�"�)�}ӱvZ�h�Ӏ�~��n��T�#���+�u�Q:��?$������y��-u��hmf���������ngV���4'0����z��kI��rԁ=����52V?Na�V�&���ޤ��Vl��l��c�4@����d$�i8��p�::�s����Q!\�5��U�yͬa���d�*<��F��u�}��i��>�Ĩ���*
��&b (����������� (��m��Y"x�lh�N�σd16������v�6���|4¢�@��[b�(@��R�)�pM�rp;n��&$o��|,q	�')�C᝸r�b�	�b��'�T�D�C_+���ϯ�>|z�OP��A�z��0����nf�~�`��F�r�u�8`s�iצ�����y�&h�{�n�˰s�(����3��5�>��?���@�P��DQ��}����?�?�����0>������'����~4�4�q�w�w�>A��}��@�?���?�����"���r��Щ����6!9t�����v'�nj��m�f~&�V��������X9�?w��<p�M���sD���c���4o�~��'촟}��aoT!�����Ù�h7����&�}�z?�6>Ԉ
 |��8&�p���C��Y�6��~���n����_�=�����~Jo��O�n�����!�������j������Q�qg�H}a������'������86?�0�醇�1LA?��3�}ߙ��������]������>A��7����?�9>��>`}İ]}���~�������n��� ����ИNb�|�D#A�QD���������ưO��v���^��GF逧���	���"(��pը��|N���`�c��5����.�.����}����˳ͯ��e���.D|�M+�?�u`������N���[��
�:�}��~��O�O�@�����V��|�?C�?���>>����>�������??�Z�`��~��E�>�G��>~r�:���)��}	�m���` (�������>����&a���?�'I~�@Q�n~!t�����P;�z���x?1>������s���D�N�?���W߁�"���??��������?����δ��g��7�m��ˀ@Q_w�'�'	�����bZ�}�nI����>a�|������d��~�3���M�0?��)���T�
 �_���@h����
}��g�>���>� ��i���!�v��>����v�0^������Z��O�S@��G�)��|��y�rE8P��F�