BZh91AY&SY����8M_�py����������  `�~�W��(�� C�o`t $z5@{�    z=4   �        ����Р	�� ��^��v��s���5[���z�Ә��� m�΃_}�s�`zt���۠��#�(�� 8@  }��[ϥ����C{z���`֏CN���� t��;�CZ7����^�t�7����/G��  ހ |wx>�[�uJ��p���ݨ���w��m��N|o*�����eEnn�����׮�� � = ��Ƿ��n��i�{ޭ��z�v�a�[��}�s�}�룰ew,�(p6>�q���^  ��}�o��Zӭ��p�+l��tA�_p}|q����;p��cZ��X1�zt�km        q����T��#�*�P�M0 & ���$�PM �2bh� ��6�&�
h5�&� ��@)� �T���# `& M0  � �B�F)�L'��CF�A��h�
�&�����j0��� �A�h4~��$j�!�C������� )������$:Ȓ ���� )��i�B����������g�����O��Z��	�~���t :UD�p6��u�̶���: 6��#�U\$�I$�����.
��Ivu�z}��#���ߏ~j�;�qO��U�4�O�geG�����g���;E�C-�D�&d��Ϗ���]m�A�ظV<�Ⱥ&�|���'H�d��Z��zK�0Z�o�Y8c*�5u�Q�֙x�B�⾱RK���w-v�y��؋i�l^�L�n��/$.ܤOI|!�w�Ԋ��P�8[��$U�a���;�zI�pW�\ݬ����M���*㘲�B��D�	n||������o�86�ò_"�7g�]$�#��U 㘊�-ȋM�]E���2�cN�F1�3a3�b��9��$�G-z�u߆ؼ4�m�i�m�/$/�R'��"�>�!�ߗd���P�8[��$���EI���Ş�a�!x�.n�m�cn<o��ιH���CB�ݩ�r�.N��,�Ҥ��{$���q�a�0zI}�Z.�.ܤKqS4|������T�Pm��%�r,�<x|��G�/ �v��d�"-6.�V��0�U�j�5(�F0Fl&t�PI~��I8�z9����:�y��~�1O��_�ݚ�;;�^zת��o���-"ҺJ�!c��78���k����Z�&.�.��b��u;�,:��L]�	��]���q�<Mx5���_(����I~[��iy��G�g�b�b��t	էO���l\S}s���������v�WNZ���[���Y��I��}K=$îI��zI}�Z.�.ܤK����O��!*i�6��6��b���9�+>b�#����U�r܈��_>"zB}Hj��>��E��\�Tg�:��N�rש��:�yߺ&}Q�)�3�������Ӎ�/��7����H����HX�������11D7�����	��R���>���b��D�^�	��O+ߑ�}�=��}k~���	�lO6��g����/s������؜]Et�Q�x|{��Ӛ��x���Ą<N#�3�	ߓU�^]�?'�R��$*bb�	��&*�q,�D"א.�+�pL^>�5H�h�X!y	�g�4||,E�<�{�ho��1\N��b����~Z��L���"��U7Մy�#���3����9�g�N�w�'��̷��ʓ���:���<�&0s>��ǒIo��RC��@=%?	�
��\����o�����{ᎅ��|�|}��v���k&��o}5������p�:�n��	m��5����	���6gD��>>1�����ৄЄ6y1�߾�Ս�B���^1��L�s͖���~�6��o+����OȞl��t���������xl��q�m�ck�Z�t�6��ۻ�y�o�q��CG1כ�������}�C���=���@�>�M�~ry�/6�L����+�R>�o�U��[;�̧,n�Y'=M��IY$��[e��d�'��O>�t�)��ll}���<��F9�})���M3�͞�s����pq������w�v�[��1�y':����8����м�;c�n������g_�l�X۱�$�r�V3������N���9�0�}x���N��n�8�h�`��0}��z�c�f6��y�m�cLry�u�n4c)�m�6[<�4���E���I��f�>�7Fyw�}���G��Іg�@�Q�:��W��6��Hp��9�'���:9c�8܃��6��V�V�Cl�����Ώ�9޼���L;'OI�歼��A�rH�l���X�І�4&�yF���n�dp�<��`�T��ߋ�����G���T�9!H�IH�FN�K��-�Q��n��C[���^�_xt}~]y;$�6��.�<���m���V�03�qi>
k������񼧘��Uܕg-��?}�|u������,o��O?[a&�u�d��U#�6��[1��fS�?z㮒W;����K�%��M�����t�� �M�����>9<�-Ɏ�s��S�ldm����C���\r��!��!�e�v���-ю;`�%�ι)��Ls�׹�Ƹ4�9���̎��cgY�����$�r�V3�ⷎ���q��7 o#9���6��3����q6&�מ��������y��9F?sc}i�O>N�-��f>�o��7wM���y�|����[�s1юn[�S��7����[�c�k�Q��;���!�Hs�s�������r��&���N���Q��������������.�އ[�:�3��7���$�G���;:�>OOO
|)�8�yKk������`�T�$���#�8G���T�9!�z¤�I9��I�I�8S�R$Q��1�wn���[�n�r��<c/��˭[�vJ��-f��:=[��������;Η`?�A.�ʉ�ה�N����2Bޔ��U��ү�G2�+Lf��#�-։r!T�h���K�����d��MҨ�6S�e:e����[�*�W-�,OH�����UX�1c0�Qڙm�*�ŊHܵ_��ƞ7X�3%}�u=ե3�ܺ�~�j}��4��/L����[od��ϘٓY�4�HY�E((p�ye�J�,N��9{�PX܍{�f��(��詎����Ĝ������iRoC+yZfŻ���䝍G�{׋q�/w�H��\`K��z������e�\�u�T}���&�zew�O�B�֏�����z>�/�f���w!��}�2^����|���=�}�;�!c���\��ʾ7Vf�(��V�Y$g��o��2T?}�}�mX"Y1��+T�����I�A-�7_��&5(���Z�)��Y������v�m�dq�W��)T�#�X�RI@g�3ݚsu��l�,�y��ܛ �H��J?�:�D7`��7�*˶&E<+��b�7.-�Ҿ�G5�]֜~�駑�&�:�zE�����nȠ�����Ug�/�k;��}x�Hؤ,�8��ͳ������<��b�95�3a�,��Q#�g���Dl�e�,2�	��r�����00p%{��������x�dߢ�7޵�f�&��d�Lц��QS����d�{�F1��$U6�/$~�5��fϧp�Z��z�s������{���9���ÿ���~k��خ���.
"�)@1��B�s�a�z����Z���3ݕV����bg!ߺ��(l�&+�CZ8��h������sB�2������]�t��o7�|x�ҹޓB���sު���_LFb"�-ڊϺ�յ��P��t���e;���_z�_{�t�/Z@\��+p��7���=9K�T���siZ�j�]k��\�$㩫aa%X��/�ey�0��m��G�
�lJC�G�R�N@�?<�����X7^�F�>����Xs�追��篱k��g��*�����G�{&�16�_Eu����y�b�^G��q>�n��8(�YS����d�����fT�ǃ�O����0�������ӻndy>ˏ{v�z~���~�7�'Sos��}���w�\�I�eܐ��ED��0�w8n�hcLz;,܋8-«
�NɌ����ޘ@��R໯,���K(����"�|����]�*�kW���~���z|aJ�?b���3�c���lL����$�+K/�ŏ��#;�r8�wn~�G����|���P=�����~���|�	"��������[˞c9$ ����1�4L�"g��>��dt�	��U��_�خ��&�!��,BkJ<�*���k��s0�9���̖�RV�*��*�B�͜��O��G�S�gs?�����v}�30͉l��Yp?�=_;'��Vt��BD��[����,@��ٳ�V�_>k7;s,��Dk���PM�fZ�am��
ݰ���-�	.B�E^x6𑼗Þl��/�F���*��^d�ڲ&-��n�N�w�MٝQef[gwk��`l�BSO<2�s���I�3q�z� ��-?<tT�_�ǝ4n��ز}63�zс<���:u�]d̢�	}n��:_�N��jx�:gr~������:� �g�z�ϟ�����ݍ�MX�w�b�lQ��k5����}������/��h2B�E7;�.�Y��;�;�}�n?��H#>0��vν��7ٌ���ztY���ulᅦ,�~:t�D6�<z/������t�&�/y����_v}�x�gžy�	���A]sf����[��nO{7v��0�x㼺�m����_���f<�~�м�GЍ0&����̵�mj����vW\U�Mx�[�9浬�['��M������ ��lx��)�m��+�j����}7M�oѦBc	�)?e���^�~=���˸���f&zu�]���Tȧ�#&e�;7����]���dY�!�m�=�v���>�Z>�{/���sϥ���#G���˟�����4e�c�o�UZE+/��,��߽d�Y��E�g�� ��d=q:�MA�Ǆ�r���];sI����h�KQlQӕ|i��C�w|` .�Ʊ
�唲�1u��-���w�ƻZi�(�R!Q7���U��
��W��b�v.��J�22:�]�����Er�U7��')��L���w��B�#у���2'Tm]��V愫 +V>�47tM�m���5)$!-ܽ�7rۏg޵km�W]S#[���{��1�|�U]���SMv���^���)ॷ{���jmc��A^��l���7jSb���*�e�rc$S���phRh��R�Nc��-d��U�4��"b��///+�Ҥך��%R�*(߿��W�I�M/y��V�h��8��ըX(�n?Sְ�)!��l�XDӉ�^Um�Q2���r�b���\��%|�_��*��nf)bl9ms��B����M�s($ ?Qk�Ҥdh9?7��.�I�j%�*�����$�����ģd�yH�0���6�˪�鲋R�C����AوU��&��Śb"���g���8w�:*��m
��0Ȯ+���� �@",L�E�z���bQѷjo�@�B�1���_�T'���.�4��r6ݒ�,�Ӟ��q9��A�PE�b��&�QX��կ�����o��f���7�c'\P�d�Q��Z�	/q��*ų�����2�M�B�Z�]>�o��7��ު�y	c�j8W	j*x�d��ƛ�r����D��F�%�e���պ����'q;���!����ynU>~���ST)�#�J�6ʫS&�9,>7yX5d�eP�HԖ���m�|�� s1g �_$j6D�-Mn+�������)\�&��h?.3�I�{{:��S�㥉5SQ������j_f)�	"l��|��"l�)��;���I|����dP�"���:�b�&�H�:�U7 ��ɐ�L�r� �8�~��xe�1��}��Ů-_��/>)41P�L�#|��BT���c��&6_V ����j����yn]�2b�'��5R6�r���93{����4�1c�rW���bQ(��C��E�5W���I+z�Ț��	��+Q����ʄ����b�4Ԁ�ʢ��� pS� U;�����%Rڢm�F���c�L�������ء��r�
,~i��ξV�Mo^"�aP�+�PM��Z�Cy$�~i?j�RiL4�%PF��zz~;D��!��������S����Y���$^��5�M�=�o��,Y����3 @� ������ x@ `t]� �( ����@  � : ��B �P@�p 0 �|��$��M��o�����)    ����~��� , ��1��p ,�8  � �  x`�� t  X  X �|��wH�Ķ�"�!����s�s� � `� : /��'��x��@@ ]�Ո  �� �8 @  �  6   <0 �  � g��v��Ȁ��?0{���{��{�Pb  <0 �{���� �;wwV �  <0 0  X � x� `0   �� : �zmC��Dw����c O��( D �|��{�t @w|� t@    �  �@�p 0( �   ��  @�|��p�O� 0 p 0�w������]w� P`A D    �@ �
  �l,�
 , A� x@ ��M��_p�I	 6AO��?P��UTH�I �o�?�����X���?#������ٓ��4~f��駮4��N�q�o^8��z�������m�q�Ӈ8��i��xۍ��N1\8p�Ǉ�M8�==;v�OM'���8p�Î+�:q��8��q���⫇8�;;N�ͻWv�n8�q�q�p�Ç�(�v��K�Z�
N���4��EDGn�A��B�#26B7k�EeP�
R�r�J�<���Ƭ~�Q��YH��+Pq�܎/���'�
�ՎU
������p��̊��-B��VK�4��R�9���FX2ȃ��,Y(��c�N s��c�B&�$q� ��Uhc�n����A���ei���~�������L֡$A`�;p."��(\C�[+QEK
�M1ZԵīLY!�LQ��Vd�(4�i�\'ћt�A����H�!���MJ��6����~�1pW7�UU�ZA�ƄI9*h�'%
�����Vr\`�Ȕ""cȫLN�U���S��x�0"%��$j�O�Ō�붓_���{>��l�f��| �J�ؤ噍P
c���D8Q�8�G�-bp�h�nX�j�qj9AzV�$N_F^���٢7ʚmV���! ��G�(�?��{�9��{7�kY@Pf,3���Z�UEUa�b�1��޵�`f,3���Z� Uf,Ә�foZֺX�f,Ә�foZֻUA_Q[8"p�d���Fh��wE��]m���!���"��ح��ӎ�q��"nGj��%U��/�A�(�[�8q�
�PR�P-"*�14U@��N>!�TMy.N.UD��w�nBZ%X���tsi��0G���P�NF�|�Ms�%S��\��D�ˣ)8�0���Òq4愺t�Jf<a��l$%�P�;W\���!�-$��j>�Wob���c����C-�M�['@���l��f��b4�F��F9&�S(�~�e9���j��~h&�ɜ�	��d�dŒ��i����Gd���u8�GocSv�[�n+��]:i�a��l����ZoIr˻
�0�5RB�y%Q$lL$vil�*]�uQ���
C����+�6�4�2�8�kZ=5��S��m�k����F^�3ي���1ٳl0�~[oD��#�����≳�J=_�C��X����7v�-ը��Ka B&�
�R{�G)2u RZ[4�a��[���&��Է��i���"SIް�P�;�5��];i�c�f�a���Y6�6Գm�j{}j)z��#��9�ݝA{^�E9�-h^��b�����f<��F�wkV��es�c�^������n8�6i���H����Q%�)Hƭ�q�����[��Z��cT�&�vtL���HS��f��=�2�z�������T����s=��O��ҝԁI	���W����j������Y� [E#�p��f:��<�9�nk�_��Ƙ�:;� CVtӪ�˪�k<�5�	�&�8��5���R��8�N���S�v�z��v�JI$�M$��k�rT�v�%b ě��r����V��H&������Ep���s.GQክ4�Ǉf�a�繊GLB����] /����q2��J�R����v[n]���\��x��S��O���I��*�%8�ô��M5y�;R��2Ia���ٓ���9xI��l82�*���W�&�]�z���i�͛aAM�\*��^#�"Q[#%9�mW�V`m�d�|gF�o���ܒ0��X�Đ���O%��p�q3�����HN��gn�m8y+ؕU1l�z��u�5�`Y���Ye�����<o��3%�둺�N+A�U���<r�X�J<8O3ERe<�+���£�C��;Ry㬴�(���:g^�׶����$-��5o�d�Ȣ�O�0v8P>�R�%������<�&(��;"PP�0b�)cLU6�Tr	k�]ݓC��/SӤ�)�M��>�35X9�BLI��ϓ���SIIך-8��yBe}Gt�VBQ�N�}+��"�@(m&���i�ԤR�R땕�i����p!�e�Ye�9����^n8�2�$�!'�������Չ�tq�x���.t���~���;�U]S��/���H묪F���F�J��[��CN}G՚Q��n��.�-"u��&"g�3��'�I'�d�����	��>0�{�I���Y�c�}�	��Y����礓�d��Ś2:!���V��ά���3�I��������p!�ࡄل0p
*#�'b�a�A�E0�8x���Ĥ��"~�O�+��M�	�I�\0�	���k���pQ�LLpL'A��=ZDz"t�<�L`����&И?�CÃ��G���xDpQ��h��C�}�+>~������1��f_���Oz���m�w{f��g�Yߡ[	�4W?����{1�k�=�f{v_O@��;�}%\�>���9�1��2�7nfL����t0�1Ը�d���Z�L4�����ۺ��ڴ��'��wn�V�#1əy���Z��6Ye�Y��v��X%խ�m����(�Q=����voI�0	�%��1���4��%RN%9m�l8�(���:�����r;�X�j��R�Řd�d�{�I$�B�葜->j�p�L�OnHϜ��*4���P(��L�L�1�D�v��:�'
d`9�ĉY&4�KK������O��&b��%Zm<2|Ye�Y��z��X%ծm�����(�	�S���)�6�3F�H�ȭ�<�ygU�qk:�euKjHD;d)��U�(�!9.�T�r�B?;J9��":q�0�V�u,N�b�#�5���(ϛ�R��-,�����
,���QxզS��}#&�=�J	�1��%%���*���(<�lCI�;toꃊ�(�C!���Ye�h:�,,D�����&�{$O��8�37�[s�za���-QZ�� ���p�}�ci<b�N�����ڗz�EO&#u��mV��q�{Շn������"U��Fc�^M����3�U+h�'�ˋ�m��j�3��� �X�+���H�,�q^59#��B52�&�͡����s�ã�H'��s���R#y�ɞʅUN��5����SY]D� ����*���k�3�5$ț��i�m+	E���[��'��n�Qd0�J��aZvy�5DXכO�$���$Lf�¨����E5��G���F�|I!-����CɌ?$K����Æϋ,��2:$ ��!�n7�E�EQEC,[��'b䢀�����rY	*�����J�~�z������k荑q�Re���4�H��"04���4Rf%1*����V��.�8�����ux=�3��a�d����D~?U�@Gu����&�.�$��C5G��@_�)p2ψ�Bi6�n<���q��i�G��j�LV���_.�U�V�Z���:�7�e0e0��(
b�"y6R�#���������ҵ�x�ʩ󊸱�h�C�\��r5Bij˩��$6�"u�r.l�`^)g���i]�2ܛn��Go��j>B�5�NpC8���'>'*J�Q&R�)���t��J�qa��~�g���M4�M�;Vb����3ּ-�(��^�D���$��$Ne�}�P �pQQ:�K����"E߬��!UP�IIqVb��%8c��J<���<Ú��3�MzI�'�����M�5I��@=p)���i�7���{���Gqr�
H�o� �$����{�&�䥨�#��Nt����#Z�6��M4�N��;VM
&��64����η� �Ưk�Cd#&UkɔƩ3�jȁ��|����Wz��g1��W��H��4��(j�1�XWPȥ�#6��pȅ��J8<��4��S�jE	i�\X���!jA��`M�nSvl�'�v�N'$d��L�	ԉ_'l�
ϻ�ʻ����Zba9Bh�x�^�6�ۃii��UJ�����"VR���D�t)�nI;Q��{;�{������8����M���I�و���uvd���J��N�"n��/9i���0@�VR�{(�A���,��4��d�t�jsZ��l����IzƊ5_Q+ć��2��1�&,9��e(�Ny)$G$)8�r�T6��Ŧb�"���J��L����iĆ��M�H4[G�Ug'�%��j�"܍�.D���
*4�D�eJ%4x�D�Ԥq�Nr��^a蒩u�l��r첬"`OA&�'R��\$���q"�����Q2\���j:�dd}�.ώ=cӣÎՆ��(�tNGP�&2D�"s�H�2Aa	P悇��I�7چ�84T�4QIܸK5IiJ����I	%�r��9�\ĩ��})���q�5dn4�&�yFQ�.r���r�J��,��n�W�!<�L@!�Icl]���O��%�ERc��
D�G֕1������H�G����\�d�]�cӣ��	�%�����n���!Tm�O�ʔIS[kt����4��b���0�~�[���3EVo3$�j��NsX+S$��;z�Q�L�u��-���}%�.����Q�n�a(J2�THCq*C��.q�[�6�(��F�[�[��#��Å�
MRq��K�%�I=�B�0O%���(�D�)�A��\:L����<<?���~/߆~��kѓ��px~'���a>��>�3Ç�ϣ'	�͌ИY+$0��}���3����pscC$�pp���'C��	�Q0D�QJ�Q�G�&
5���Q������V�&%tpv6a:L�p��	���M���A��0Q��B��	�D�Q�UQ�D�+�'F�!��Çı����|'�d ࣀ�Lpk��y\ɿ��t�l������2��;�*�����x1�i�H�'j2�e2#���m��yySB�#1���fz'��µcw����k�S7�&,���p���R-��W0�m�7�c�rgf��[���}��/���i׋�7вu�z,岹�,��g&
���Q����b���Ϝ��[Tb�Ҟ�q�|�r�D'[�w�y�������<�o�}�=�۹�X�����t똤>!.N�x"���7g�<X6ζ!ѿ����u��1W~d`�0��k�Zݝ�j6�,�%djs��;�u�0�Ż�Z��F�S?]�,m ���J\���0Q��>T[�3D�?9l�9�뫷}�ͨ+���a��m�%���Ź��;��`/��؜�)\��2b���M7��j<�˭m�,ڪ�4����w�,�ݖ��M�zr�N<dx���;�z��W.@����K�a:�~E�k	�e_�3O�K��9�P�1�q���.���dS��HЩ,�4�,(D�_�E��������?<�Ƣf(�8(D�m��`X�9����_�LU��<Q:�hƇ�G\n�YqIuFg0B`G2 r	>4�ԃ����RN9�U�?l�6��+,v�WZ�9� px�j�R|���Cr7*˲ݡ\��/���wZ��~9<N�<oWw�v69�ww����W�M�S�����e���c��wy��̻�[�$������eޭݒy�̼����Z�6B�A��� Zj!>N|qW�2�	\M��WA�5R+	]���c��R+I`D[g!AH;$�A:����e���
��$
��qZ-��i�Wq."�������H0�m�"����/ZI,DR�aZC<I$%�/��u�i�e����>�ȷ	!���y3��+qcUKs	c��Ɩ9)*�&Ҕ���"k���QF@�RD�e"c�<��$h�tӈޣq�Y��F�kێO�"j��P��u>��iB4�Yh֧�Ő�Q|,�J�`�5��E�R���M��1�G��j´���ZTFI��
��5��(�A��R���3�<��a7l�ER|��+�/ +��ͦ�ك. ������n�]�ħiW �ȃ�����r���N^Ux�$����KT�8Ni6�tD�F��JHN��p�Z|��d�M$d�
J ���~M��2�$���%%|6��ƛ==v�+M1�uI.�Ȓq ϛ�~N�1���dN���ô������
g)"QM%�)k�����S�Ĩ�Hq���E��,�*�4\�UJ.���O7��[��g�	������Z1*��S�V$ ���I�9J��U9t�KO8h��D�$�����Ӎ�Ԥݺ��N�G�[cӣ��j´��Ү1�b�Vd�%'r�SEb8�R^�I��2�jnMѝ]�\���Qq�b�ƫ�L���ݎ2�0�6�k�JL��������\qԻ{��ܑ���③^���Ş$���"�N�&S%&�n4D��R��$�Tj'pHI_Y$�Z4��`B: �n�jR@8�)1�(�1hD��0��So�<QEh:8$��g9W�5b�]�57ɟI>F�����&I�dI�)1��r�m�)������둺��t��uo���O�^��>]qw����U��:dfs9�OE�N�b�]�q��
�^!-B�j�NH%ŉ��[blx@V�R�G���U�]]D�l�Jh�Z��D��8���]&�Y�h�v�UU(�G\�t4�J�ޛL`.Ҹ�/I��Y�ˌ��B5�"R|G9�KF�f	$%=q�$��(�*QX�a�L7JN%e.��*&ʧ�Q �g��))�F�6h�h�ɡ��lbKI�Q�Z:�qGQ�K�ۣU����}cӣӷj´�o�d���Wq��~�)	ǻ�P��SI��\@ĕ�"e8��>H��"'�I�S�1���!��>M��S���Nǐ��e��Ř�����C��(�6실�����P��Y"����D���fR	(��f	Idz��������G&LN��l��WM:;<v�+M1❂}9��*��6z� ���|�q4�~�B�)"D���z���
S��H�H��11u*T����4��A���LZ*��D [��9���=-L�	�$�O��6Ә�����&i0�7����N��������)�=�RUG(䧩T�,���I�	(5O��x��Um�F�]�
�Lsst���F���G��Z���ۓ	�Za)���N@&�sS��p�yy/sz#D"� ���R�4z�IT{Q��|��	�%:b1*�$L�G�i�I$��I�@7�A��9Ëؔ^9D�	�#�۪H@8�JL�$t�JH�+i@TMx�֚�G#���OU[iѳ�j@HY
�7iw�}���B*}��FG|�g\��t���k$[��J�fa���ޭ�7�]꽪	�U���nf�v�Z��t���	T�*��cS���1s"����\NpU4�Y݄��He#$O�����3�Xz�-E4})�R��t�JG� �A��4�S�kHݥ��I�F[~{a �Jb�H�㚒IR��H���4b��|��#q����b��N���>H�MD��Zy=JP�z��F�p<`�:Y��p��	fjο�Ԛ'n��_���[c�$���H�J��ϛG5gہQ#�*&M���QM�g�*cС.<�X�d��`C�Y��"k�!`s�-Nr��9�KOl���ޱ��ȡ���J�Zi�u2Ru6z�I�@g�K �&%&S��~JR��LJ F�QOz>��ۑ�?��|CÇ���;'ä������_�������t���	�L��p��d��l��Ǆ���hL��p�L$0�88Y0H8~'�
84��GG�D���
68"'�W#�IP�V�'�C�0v8::LÄ0pp`�&�̊#��h�#�#�/�2��m�^�.=d���_W�~ñ�0�0Q��<LÃ��Gࣂ��X:7���{Mx�~a�-,o��+��|����ϙ��Q9؋��9r[�����Xi�G=("R�h#�SH��%<����6�Ͽ	�׳�E�#��+G�|�������M�����������'�����9���������̽[�$������f^�ݒy���m�3/V����wv�����I�V��N��
�i�)�̏��-��m��4�[���G����Iz�g!wWup�ä�p�o�I�JJ��&�KF��D7H�b�8�P�n'�ZO$qI4��D٢i��m(B��&e�X���J4�CL�g+�e�]�J�né�/�"S���qV}_jHKdM$M�_]��i��۵aX�9�ڱ��`I7nO� Ha��y��m����_��@�ye���j�tto$��.�a�!	���b���N��ˤ�R:O���g���5RͧS�Sn ǒ�v���M_�x�}���r��Ⱥ�#��jqU������@H'���}��5�^���h��(��6�
6�QUj?��l����Y�qEUBp�{ۻ��&8�L�&48�!�]�m=|�����[ʱ0���+��Y�J�%�-I�����79Yl�i�I�H�� ��i��d�丮\��A�[T��B�Zț��kf$"��a����a��p�Ri sob`	�=�%�p������SKi��"q�,H�Za0~r�S h��B��$5�(R}�յ�>�Y��6�㢱꫷N�G	 ���m�W�Ԫ(Zj�h���|�7Mjd��TZZF�`}sD4QV?o��^i��	e˽�b��}�2d�w����Uaзdku�L2��S��I��ai���7YPW��he�p��4�f���A��6�E�6'L��_&���&���FI�3`e6�~��I�i�o�x��0��x��hڰ�W2Κ��0w�x����Ν&�ҭâ��#6U�-☒��El{r�Ym�i������n�E��Gk�~S 鶥r���U�������G����[�r����y2�`:��׮@c2I'����𭶪��Յbϛ��ֱ�q�,Y�m�������U����Н'��#�P�$��y-6�2�`q��οv���+.����	F�L/��k��$<Fhbm4�O&����Kp8�'�c��ҫ�j�4l��aX��}��tCo��H�������}���D;i�ݲ(/��o��x�iuȷ-oPѵ�̻�x�=�ު!��Y7�^6�b-5���{ZN�K���%pHY�v�A]�<��`�J���U^��q-Q�M�H�v'ID�	%�V�L:������h�WMz���,���I�ñ��d��QRUaϯY�@�N'
�V>�]�����YWi�	�$��O����__U^�l��aX���PB�FhC4Z��!$L'�9�V���������T�I$/=uRHé��2��
U��v�M�I�	����9���0��:6�^�hK�$��֥ѣ(���2�T�(ۤ� i�d:��x���:CDŇ�� $n�y����{k���s�G���Tf_Ԣ��D6KL�R��p��)������]�E*û�{��[�D�f��]��W�R�7uwve�����>��r����!���g�s�6�.B�9�JZF�RE�`|�ԛO�����O�(�E�[V�2֤�F�����C3��%Կ���%,�T9.ZV�����-9��nX�S�@5�J�.˞����7���=��~���l����HBP�|�5�0�-�㆒�,�o����t�����M�/���a��x�/��:j;���I���0�,��8OO	������8:0�?C�k ��?���:C�����||~���8:?C�be����&��0�888h���#�W����A��~M�W"��t�Z��'á���\!�c�0L5%xp~$]�2*&
9Jࣂ�&`�
~!�W�Q��z-�œ�?��k����`�\}!�:d]�̊����]�8(��	����K�RS+Z�U��Y��,N}S��0n\�N����%�f�}]�n��:]K���$� �RL]yqa�㌘���I"�0Ӳq6�ll��(��v�f�l�a�K�/f�v�Z�&�ae��1��|�\Ǐ�"u�N�[1��g�,��T啸*�$G>=��z����s>��?�(�&�[�,�(���?�E�F�3�-r)o"�� ƾ�E
���D�a�_�G�,�^��;�ipM<�8���)]+�s��&��2X�5�YJ*L�V☝�Ϻ�ּ�y�vY���ų��MK�"b}j�e�Ud�Îc�<m͓YuO���#�X�[��vG�>w�L�V1FtR'� �U���Q�Q;�ۦ��:��yi��y���R�cQ=��MR(�m����N�}���l]�퉍
B��h��T�|u�_f[\�Hp/���Sd�,�!Q@v���
�1�:pnʔEQ ��%�g�k�8��y=�c�Fީ����SVs�<�k�X��m��B��)b��5j��N염N�m�=vx+o��z�^�绻���̽[�c������f^�ױ������33V����wwn﹙�u�}{���w�̤�Z����M� �o�I����݌�KϜ-$�R(^I8Ƭi�	I	X���E�Q�]b ����$�+J�NE+�؊Un;S�A"nT��r4�U9k�T�	`(�NU�u��9丢֓�l΂HIER�]R�q"y>�`�M�zd�46�;�	$fƒ�9)������P<ry6h�@��|^�CI���hgC�ƞ�9�5
��wx/U���Ry'��8bk�&Λz�1���Յb��[p	�	i`q�GY�F`J�q6e���JŶ�Jw�IEQTU|�N�����wF ����/�RK���m��s[�iS�~���>gMN��BLq>M~�e56�C�䲪j_ѧoX�>�p�]�m�aLVh�W�NWJ���&�#��I�����ޒ��R�T�$�r����n�7f��n�}��Lk�cf�f��i�<�'G{<����j<���O���>�M��������TBTU;�>�^S<66`!� B��)ʪ=Ghί�!I��vIo�'L����Ve6$C����d7reoz5�V蹉�fa�p�1�K���{�Sn��#n��y=��'�O!��K�%{��BR�T�}E��:��@���p�މ��d��+�����x�}����|��=�1<{i]Gi�2b�v؄?6@�&�w���^�伯fb3� ����W�;�k�g%�,�j���:eB���]6��4X��ؔ G���F��ؽ�;u�u��̺߱=]QE`4uV�`�D&�U�"�L�(�?$�*ef&��E�f8xJ���QfN+�Ēө����R�`�a	!�ѐ�l�RCn��Mxvq"|��`m�`C�Nu��d�&C�v�����úѸ;�k9α�ߺ�]�'�]���٤�M�k(��K1��s��f�gݮU�gv�1�$�hDD�Y���> B�j�L�U}ɓl� �n��x�X|&�$��;KrP넬��Pd�m)��I=��O2�7#'�H[Y���R�u��?6[�ys1�s1c�f&�fL[P�Ą�m#xH�K>��RUT�&ӁU�Vgk�����i>�D��UmӦ1�)��l1��_��w�-�q�8+�&�C�Z�F�|d
�6n6d�|��X��?m,���V0��R�"�*"/vm<�J��U\��jI�;��7x�
*Vo�O���~�!ǆ�%L��O�� ��טe�2��N���N�B�86@�1��I%��T�4��U�Q�������}��\	�IBT��G�v��U2���iϔS��!�ȫ{�:s),9�Hi2�v�9$!	2d4m<e3�tO'	�FG��;��^���Ų��F��㧌c���hHB�s0W��l���uw�N�����V����']�Tg�����k_ue	���o�*|7ۑ2�"���%0�d�u
2��!�$|�P�.��1����'��H��1dCP"�-T��Ӫ(�mVܢλ�2l>t�o��I��7F�-0G�\������E=F��a4�wgN���o'�]ļL�bb�
��s���~)���H�>�Ob�z���\b�SӶ�aGk��@N�u4�^��2M��_3�^��������<��_��_{��D�#VٙG��u��5Vɣ����b��#���jԀmƃ�y�`/$ C�{&Ε��-L���|~=l&&	���}7�ä���<L��Ç�t�<&��	����&d&��Dp��'D��tp�<r.�&��&ia"8
8~�������t'�'��Ү-WkW���*�j��Y�vȸ(����+&	��v8&�%`��|CC�]���
&
8(ࣂtk���~_�����^��>��v�W�;��||C������E�	�#�GB�
&`��s�]{>��w�Z�I5]����n�I�|�Ş��I����SS60v���&��f76���y���!W{�-B��Ɔ�s�}��s��w��պޮ���ۻ�fj�oW^�����35n���wwv�����[޽��ۻ��j�oq�ffo{�y�8pD�pC��dC���'*� Ru�e)�e�u6m�S�����>�ɰ�7�M�1��Wu��%���+u��T�x�>6p��Ez�1�1<�l�)�h=�f�{�Y��j�FQ�Љg�� �8d���b��M�m�:�Pi4�+3���c�2�e˘���6 B�M5��}�p�і�]H���.�7��$k�h>�J�*���?O�#$2��e#n�:����$�lLi����e<�h�<h�4l��!t����ڗ٦���ǜ��Ǣ������tқս��Ir\�4��eKcƲ��32�����jڭT���&nI��%	���k"��LuӒ��"�(n;Ɓ����J��I)5`�(G�2�G�ꀙ�����O �Ï�k��YKJLr��ZL&C	�a3�!��N�2KKN���'ϓ?0w꯮]��]��=Qv�=HPn��7���<t��D.�����r�F�Q���jt�%u7�m��x;;m�2m}���]�д�@�e4�m �=�<kNS�M4��I��ӈ�С�~�������"[�B��ԍ��7R���*ꌻiF]j�7�:Ko!�����C�$"l�p����p8l�~���4޺oZܖf������Xm8|��f�&���n��K:���{/(�\�	
&1p�Xh�	,�G�ݻKx�O��3AtI[��k$c�a�%�mˢYn��]]����!e�GHf9���_Uq���J�sKYUԒ��ȓ999x�]گ�yC��f`fUE�lc��$U:$D���/���M�M�����K��L�}�$�iu�$��ǵ��>�ʾ�J=���6\e-2�-5���z���r_254�U�^�;;R���aIR����q�B�ITuE'��$y� \�1Z��ǅ%Vt���>����n3,�j�e�,����h��؎��$��T�*� F��I�7[`
cMg18LHU�iY�䒊fcV+KZu�!�H�N �D ���E��I�}�Zeמ�5�q6���HS�q�x�`:Ӥ�D0bi�o�=��:e���y�%�,H2@c��rDH��@�4���QU��m;�9V*�z�����J۾[n@-0�Kf$��L��	�8OG���������g&��ȪI"a<��)0e6�'�.��	j��+e�*���]	ƚhV�&bɖ6i�R�-�a0�M'���jX�V�Uq��ڕ�u�'�n�3Hn�z4��;_DD��!�˕|�&D6Zd�3�ߛ�,m�q�UJ)q.Wn�&��� �%h�,��R�=��a#U��g�LL��'�r�L�e:��L�}Ԍ��XekTJ4lD���ǃ��+k��35�U���6,�|��J=��o��J�aĄ�JKÑ-4x�q6��4Ogu:�M�l�4&h�EQ��h����,(}d��c�!��S�m9��8y2�u4�L�G�L�+�jp��g�O��,�+��t�zL;�����0|�0�O'��x8r.�&��D��8=!����d�����"��hplr�E��G�G	�>`���������ñQ��ׅ�'�?��	�E_¯�|0	��p�C�����0�	�`�x��<5����"�"8(�(ૄ�t���
�Gᯉ������'į���&�!ᮎ��̵G]�(ૄ�b��N�8k���Z+Sj��5�t���j��;u�Gˏ3+x�5R=�#w�7-�U.6R�(�FھiZ�-lȡ���+�G�W�ǘF���m����3(EҪ��y���g�T��	���`�,O2��d�.[2���h��^��4:f�*ǝ�k�;X�����j㲲,���]qgV	��2*��+"}��6�Wc�:�n�H�phr�LvU2�UWr9���R�}�2<�i��Vr�:B�x�b��R8�Sу���%G��>Gx�q�,Sm�A�n,�����<m�"�T6���X�Z&�(Q$i�D�z�%\��Z rr�G�kyg%��a��f!З�'����H�Ya&�b�N�š��-h��A�)6^;m&O(B�x�\�r�&Q�W�� �2��B0�0Qf�T���o�Q[�6�i9�80yP�a�67"�4!�v�ͪآhnהx�]��h}.dM�k����U8,M��+d��']�1e��Tm��T'�/E9Y�`�5�՜k�@�QR��2*��j�P�U�T`�E�~"��౸i�թw����^~s��f�����1s�fn���s5n���wwn����u�ǻ��UYz�n���wv��/un���wv���qZD��� �pA6M��rJV�T�����Q�EX87#��]���R:"�F�6Y\���E@T�������9�%�E�!�Pa�^	��bb�`�"�:���8��T�U[+i�Ҽ�,L�B_v����g9��)0�i��W_&%$&Ms !��������땀��9p�dD��ȭv)��mH0]ⱑ��ө���|i�*�lxv�Y��y5�&��o%�G�2rK�Pw������S�ن��q0�I�n��_aF�9CB槣���0�ki�Z��Uc	x���*���)�gC�>Ӏ,"|�J�g�$�'�Ǌ�}Ux����'�C,3��L��vO�!(�7�#f2�����)�֪�M���(�h��u���T����A"E�U�.��R��q2�U��&ߴ�}#��e8������,��ߓ9[�&2���,��UX�U�c��+׺��U&�˓kVq�i%�����1.�܄T�����7���z��?u�Hl�(�*�nGi�G�d���ک��i6��<&py(m,�~�!/�ΞG�����1����K4����F�h++�L3�w�,��2��k��Y�Mo�or�V8����=u�Of9�^�Ƙ�R��Q�V��9	HݣR<ˍ�W�@w����RDv�qb�w,	�v��&�i.Ւ9G(k�e�V�&mό�^��-�ļ|�4_R�xQe0�ݢ���d�Z�P�%O�%`�-���IE��m0�I)Y[�;����FFA��#K���2�zJ!�����qV�?��(��6 G盨]UWlйH�2�R}�2kgZ3N[rTM&a,�0I!�?d��'��*�Դ�m��	|��?�؉���WI:���ٳVBGP�a����=FQ�wh���B`�0�Si�eǉn�XG���z�1���ڕ���I�u4��$�=���l��Io ������3�qjՙ��d��Ԍ�aEb�7UuI� m)!���q����x��s�Jֿز��/E���m#?L�u�~t�^6*��a�e���-��z�9:�_��Ne2�YB0d��m0O��bt��'2QeQ��gjV��.{r�U-�#T���8��d\<�ga*UF��9M����h�1��"V�a��fe�1u0LZT�?i6�JJ)6��C�N�,�S)����%i0��I�ϘCI�����W���=p�>L�:ն�}mlx��,�o]��4�M5��K�j���n�;�U��L��}4;��P]�\YE*r'k��ڬ7���q�P̽�����2�H���XUe�"�>J����M"@�U#F��`H��-)
#�$yF҃&'��72<τEZ�P֨��>?k��7G?d���&
tD��ɖ�aI���Ǵ%EUg��j��2�ꮻ����qgȳ���9'�ԩ�c�ǏC�	��V�H��{�Y�
¾<��!Ш�K<G��.7u%T��8Jr�N�%�8^_^��*��&�D��q2�;�I{�o���ʢB�$O&�8�̜6l���>8�ƚvۦ�q�n<qǮ=q�����m�q��Ç���;q��x�N4��N8rr�;c�8���Ӷ+��G��z|�afl�4a�0p��x���J�Æ�8q�gggo���>4����Ǜ^8���n4�=W��!�?���m��g}��{�����7�r�u�O�p��Ȼ��LH�����N����|6I�G;w��\}�Ui)V����bm�Û���(��w�����e�i��r�����P�:ǵ��I{[��Ͼ�kZֹ���s33Z���[���ݪ���[�֭�ݪ��[�u�ջ��UU��u�ջ��UU�R��Elcm;Uv�wگD�uGr��^�M랒I$��3!+Ĥ�A�}�_��X�U<��QH��0k������7E���)�P�g�\��wܫ��t��s��7Q-�3F�i��ĭ'�BON���[kq��1�x�<Uv�N�*T�0�$���&�Oe��~�m��kܪQ*�(�
J�TtH�H��##��H���Lq
/�$�H��x~��)�i��I��t48˴�h磌�Q��:p�a�0���N�}�lnZ�eL>�)��>{6w�;�ex�g^����u�p,��.6����Hn�CY,U��@pG["��^5���ӶM����[S�$�J"���AǑb*�%ɋ��/Z����8�I����Oe8��oX�ѩ�M���i�G��z�U�W��+Ë8�U��� �IÅ�Mq�'�݃q�IP|Iu%�iu��7=I�����>=N�]�&�'�d�i�ME���������������o����97�{�7����ڶ6�pcb�k�r_�ėwf(�.B�p��q4���b^�'�%���*�:4*�"x���8x��M�����>�z��J�y�a,�Wx�p���VWћ�+��qѫ4�՗uz�B���!��I�ɠ"u1��y�%�0�����Hi&\lܐ�t""t��Bt��N&q&�rQ�Q�s����lx@���Y�����>��5��И1�$�'��8�=���lbm��r���&��t�,�i�͟'HCe(��,\��	3�������fO�y�na�<ٶʜ������Y#6�&&/?ӽf��M]�+���J7�kq�;��߲yuc���l�|٩���HDi���3y���c/xD�O�.������)�$��ʢ�4*�
�-p�z�������$"A �A�-<�NjB�ӗ�q��3ͥ@��@}�˷�+�ZY�ͦ��C�D��=׻3�1U�ǜ:N��R�P#q�.X�QB��WK��#���ϳ��1�m�z���~�hTOe�Mp�Qa(kP�?<�!�(��ې��u#k�n%S�֒&�!2�H�0�z�>�z&*��d*���u7O��Zy�m���#�^?Qu��6wtҭD�:�Q�,D�!p�\�;��wT}Fw츱��nBZB��⾧\	CG��air
)����v�Q(�42�0˗�Wl[Y%J����(�f�"���+M0Ɲ8'өi�SIn���ڻ���;�i>�U�v�1뇊"p������M�|��w�G{����tV��s�I��'pk�E�1dH޵�sRI��>�эj�$�0a<�;J|����!	Z˓�z%��9~1�*J��%B�4���ɤ�ʋ�ݯQ
�t��44��8㍸���<}q�v�N�q�8�ۏ\z����ۆ�m�q��Ç+m�ێ޼q�M��N1\8t�Ó���q�|=m]��zS���+���Î�c�8���N8��|||8��|>���b������F0N�x�ǭ�Ҹz�N'Wu�.o&1��|����^@��螦ǄH&"��إ�
k�c��~�73��܂3���$Q9J������32�S��٦(_n���IhvM��=�kr�V�J��=�,S"�Z��i�KR�1a��y_�rG�2]���V3u�8ٗ�;V9[���v*W�wZ�S�Z[95�*���G&�X1fO��4�{/1�*0M������樽�9�l�UDp�n�E�M��hn�B�imfE,vduܴFe�1\�Q��b���Oe�ʇ�:˰��w�8���w��T��k��sS��&����LR����b�U$��,>�XY3;$Q�\���h�Y��q���(�RYJc�1�ʑ�S�Z���Ld��N�5�so���|�!^0"���qcS#�QRs��^(��Qk߶]�+N Њ���}>ǻ6�--[|����ai��J�U�H��m6*!4�!1��h#�5�B�V5��4��1*�a1"#D�q���,��X�mUj�U]�X����}����=����k�a���335�Uoun��[��UU[�[��V���UV�V�����kZ�ᘷ�ffkZ֬Љ�!h�pDN�6qXf�F�R+T�J�n�j*��K�rX��GU�(	�ڼr؅	l�+x:��b��+Ul�jQV����&YQ����iEU@�K�ݓm�F5�Qn�K�֚�S@�.�R�.%��RF��B�f^�}�r�'d��N�>$�	��4m?��	���?t@��w�����4Fl��4�c����u-H.D�.�:��S������֍�b�L|c�Ӵ!�u\����Ҵ��L�Io�$$�v�Q5��g�|5�!(�~�#$�h��$��K��׎�.�j�g~���H� S�bKT���u���UR��IvY�n�I{N:L��NBh�舖CD!�!W�%��Ӧ�)�	5��BO�)�.p9��R꺤gl؇`�ۅ]T�D!*���ɖ�&Wɽ'�m��=�8�>2i�'ɂf>Σ�G�Uz��1�ޞ*�c7���䪢]�d8cIB�9���Ζ	�1 �r�&�hRSPRR���s�]��������B�m�c�bꪍ<N&��6�z�t�i=��N�@�	���)�&I$$JM���'���*�c�1�ݝ��c;ά���p���u��A��F�����|�^�9�N'��j/��;7�1����k�-uμvbs�fZ�2���^5jUbG"u�r��Q��T��Z�)-CM���^��i`�����yQwFv��pH�&c!	���[M��v8O�P"q8��$<��=�&@��L&4�t��D�Ĕ��r��Wk�z��ʄ>!�����7�+�a�w���p��_�'ɤ�q�~����섐br�Q�b)s�;E�x�̩��mU����R�����%��e���4�8=�����K��.˽^W~�C@9GhD�!x�p8@���Ϸ��!e}�S������*Jt��h܉ǯ\������ϰ^��d��fX�X2'E(��B1����_��=���|�v,�F�N�����}���1��a�O=)}v��dq�Lv�1�ӳ�Qt�!`��yԐ�M��]:/疟��v�Imi��·SwUI��HKK�f�m'�<L�a�&$�t�<�>!<���Rk�M��7�֡�m�z�0��E�QF����i5����[�����f���%䶢�o%n�;U���G+��,w
��s'2�ҹ\����u9v�phDQJUYʓt\堈�^K�[�B��`�U�mBQE"m0�M�'��"e2��kn���UU
(����"q��I�s��#���;!'���:�ۣD�����)��1��b�ҪȐ�B�]���ƕ_�c�öb������WwFAۤ������N�u着��%4�ru��2���;��u��SŮ��"DE����ZL�v��c4��I2�v�Li'JV�b�]X���/!E��!X��8�\z�������m�q�1ÇV�i��xۍ�N1�+�p�㦜q�M�==4�����|8p����񎸼q�8���Çq]�:�C�D��`�'�|���i\8q8q\c�}Y�fyr��{w����n��6����{�wݻ1^���"ߣ�=�8�~1�����{����h�O}��7�ƳT��F�}5|�ڹ��K�)���գCj��{���ջ��UU���mj��ڪ���z��n��UUov=[Z�wv���}&��׻�uU\T�j�Z!h�p8@�+��E���G+�U���Q$"u>0�Kt�!!�l���7j����յP�MIO���ϭ����B����N�s�+�i��'ٓ5U(��ɹ�bi����=p���DާN�f+|S�qw��9�j��ɰTvJJ� \PV2)t�����U�.Բ�e)\L��&��I��$dЙL��B%2����m>���[���Β��#׳Qc�kJ���Ǯ�͡!!o��Z���oI�� �ٕ}M����s��r^[��%�d�2.븶�M�����'Z����`�q7_$G�&GbCP*$�n4����$���%��dA$D�v�Q]�4��40U}��f��ӄ�޻N&��$!�N|�x�I	!i�<ri��Q�8>�U�e3���9�����nA�ƚ�Q+�j7�'���n�VO���W�;c���h���ܒ���VL#����;):�+�$v�NO%�CFݳ�Uz��̆��'��2ex��O�\'�\�R�BIcҘ5��Q�8g��}��nD�s)�fHCeQLxzm����y�f����&�Ɔ�d��yO'R�>r�WC�L������$�r���NG��';�	�賈��{M���I!	���c^��o��t&^�&KK���8B�p6@��a�U����QB�����X��dmin�1��]]�{�g�$�9����f������x2�dZM4f=����z��i��i���L�SgDK!���d6�L�;z�E��I��ƥ��ZZi��쯙!�5�L�eOq��̃N�k3������cqv&�,ZLڵ��]ۙc��X��-$jJ(���Z"�lQS�rȝƉ!AÈ��D�a�WtUA�7�ɴ��0[	!#�Ͷ��8�KLd��I���z�|��0�q4�&L��		>�'�+5KU�۸1��\����!.BHA�����r�l���U+�M�����l�9ޖ݌�/d��y[V�W�KUq��c���g#J�k����]���U��Q�[�"&��WGO���l&�d�#$�첮�i-"t�$$8ᨴɛ5Z��R���eq:�D�4��<� �vnC�٧�[�C������C�����S25\�U��]ILCYue6��HM�SD�\K-<p���e8���aĒL'�B+d�x8(((�J+׻�3`�e�Ӏq6�JL&�%��O2B�awW!	iN$�J9��ki�����D�y2�)/�m-:��!!LN:̤6�%�_�����$HD��I-��m%�1�៖~����]?�K?����e��AWfhF��0�[�M�odD�(������*R,��Q��FDX	 $E��Z��T�D�,IRQ*J%%�E�QaE���#
(�Q(�QR(��XJ,��kДQ(�%J*IE��%(��*F$QD��QD�ĔQ(��Q(�%J1H�(��X��"QaE��Ģ�E"�k�E�Qd(��X��!E�(�QB�*FAE�J(�Y�%J,�E�(�Qd�`�#H�Q(�%J*(�QbQ`��QR,2�d%"��d&!E�(�QdJ,���#�f��p�j����:�Qb(�%"�%�*X(�(�,2�a(�QR�QIE�E���QP��Q�FDQd(�Qd(�QIE�E���E%�bXQbQd�RQQ(�Q(�Y%$�TJ(�*EK��E�Qd�X(�)%�%
(�X(�Qd(�J,�"�X�,�IE��E���QD��E���B�%"��E�(�Qb(��X(�RK!E�!E�(�X�,�J,(�RJ�H��QQ(�R(��TJ,�EH����IED��Q`��QQ(�QB�$��)%L.
�03#�(ZB��b�-!b��b��K��,P��eKD�R�E%�P���KB�!hX�YE�YHYB�(X�eQ-*Q,RP���,RYAb��K���K���Qe$��YE�,��Z,Qi,PX��Qb�YKKR���X�i,���(��YF)#"�(�E���S�YE���(��YI,Qe,��,��E�YE��)%�X����YAb�(�E���,R�,Qe)%�X��,Qe�YK(��(�BYE�,Qb�)%�,��X��,��RX���KK�K,�X����U��e,RʱVR�%�YK,��"�X�)b��K*�X���Q:��Y
�XFHR)�H��$�T*�%D�,E"�DX�E�b)$�XJED�RR(����Y
"���H�JE"�d����H0��b'�k���~�~]>hJE	���?)��AD		UD� D$! ��+�I�?�_����μ�}���K��U�_5�z־��~}���?޾�|�~�����qy�jڿNyn��;?���K��	����i6�*���z\��_��|�T�%���ˬ���T�I"?�?'����������?0��d/�`��'�!D������?��ܟ������?��)��/�A?���	��>?w����4~��C���p��UTI���#������$%ihniC����n�c[���������S��Q���٭o����b~i�����X?��)�fB!�o����ފb� ��h��
 U�)Ej*
�� dP@> �o�F֙�¹�����?��'��u�������>�����T�-@���'�$�*��2(����7��?[�i��w���H?Ry���)�y�������[�`G�����?��?�*��Z#@r�k��Կѽ��x��u����Wd�7�3���JC�+�?�?������������@�i��?K�����_��#�������P��UTK��`u��VC��+����zl�����:�C��DL�?���'����E������+��W`%�P��~#���N���m %����P�Z�RB�$���~�ETJ ������l�lb�'�6�K�����|#;�ç�����7��{��1�^	�� R��5��B�����>���.�1UTO��P�I�П���?��b�?`�����o��?2�ҟ�I���>����O�?�O��~�����xg��R"~��#�'�G�����L  
~E���(�?������W�/�UD�?�d?qݟ��9��O���������t�2��c� @�$�,Z������KH?��|'�� <���t%��i��p�A��}��"���O���?��4B5I���?�?����1🕏��߫�6�>�H�������̆�(x�����N"~_���П�AJ>��a_����??�v��� �����{�~�]�z�)?7\����W�!�	T�i���7�����]��BC��h