BZh91AY&SY�ѡ��o߀`p���"� ����bI>�     /��R��h��I���6ƢH�
�M��)kI%+alT�[lm�ژT4Ҥ4ڱ,+Z�m��H�E*��Y,$��㮅"V�kjc&��aI.����"��m�mB���h�0�e�Dma���ؠV�Ԗ�̊�T�P�Zj��IKCZ h`�붪�Y`ܰ.�Vֵ�R��T�*�l��˳-�m��Urwi[f�Y��+KeY�(�I*H���iE)6�[
ԕ��a�B�̄�Z��;XekiV�p   �����T�=��wn��ӣ��Ƭjlu�ٛEvS��cn�֝P)Z�U](�_` �Oe�R�����jWT}�<��Z�Ȣ�eZ��+&o    ���M�ޥ���
�{��=���׽�����ڞ���s֪[i�Ws���^��&�zo{l���m��}�_[��E��J��Z5�s��ٔU'���_4��dֶ���*k	����  �}���kfk��^��/��x}�|�6ڒ�����֫m�����ת*�C��ﾏ�_mN�����k66�^}U���	}e]���U^��_>=��ؾ�U/�{6��l
�LYTm�T���   ��|�z�t�������N����|�ﾺ����l��������f�j޾�>��jU��S�\�x׷ܤ�N�^{��Z�����|�ҕ�R�������UM]�ǟ<��a�wk����R�j�KTj�H��$_   �7��6��;���>{ꗪԔ����ﯦ�k�]�w>>��K�Y3^����Ol5�5��ݭ��,km��}�jk�s��������u�T�<}�ϴ�F���罯:�Gr���Y+lŶ���V��*U|   ;�ΟJ�'���W��o_m����kmh�s�T�]me��Kn�Ͼ�/��N�+�G�x�d�6޵�Oo����YR�����*W��y��ԵV�뽺ދt	�kIV�M�b�UTUV� ʅJl3>   wv�ޏ��V�����'ֲ��ɳ|��=�j���r�����d��u�=�[oJ�My�7<�)���zZ��h4'zq�Tzr<�N�(�]�H����J6ֵJ��),��յ���  |�i�UoW�ïTWkގ�������E
���ǥH-C�uTn�ztp=
W��\ 6��Â��j��m�={*�ɪ�TM��h�   �x֏�U�u@(s� i�]^��tQ�v�z�8<B����M[PY��tV���Хa��������5;��٤��DV�Ԙ$��[�  <��H&�� n�Wޭ�Ox;�����P���:0Qv	n��@u��ދ�U�5s�p�]V�ޯN/d�wk�      50T�T CA��M4�O�1JQR�@`� #O`��I@     T�UJ��@� @ O U)��     M"$�)	����#�Ph��Sjz"_/���ј���_�&��>N[6>g�y��;zv�=ϝƝ���w�BI!$���( �NBIH~�H I'�	$�O��������$��@�I	"��*��I	'ȇ�A���!$	'?����\d?�HTBv!62M�&��l@60�M�&��$؀ld�&�b@��,H!��2$�b@؄6!������@ؐ6$�!� ld��@��6 �M�c l`&�c ��6$�2l@6$�F@��6 ��� ؁b���2 �c lHcM�c$��6 ����6 �M� ���60��bI��l@621���l`b��b@ؐ���� l`&�b� ��6 062ā��6$�b� lH�c ��aCb؁62I�$62�c6!c$�#M��Cc!$6 �� Cb���!60$�Đ!��%� �!�!dd���B@��60��Đ	�$0	��Cc !�	 l@l`HCc !�!$6$!���� 1	$60��$!��I�Cc$�6!$�$!���6$�����ld�� ��!�؄lH@��M� �c c!&�ؒB	!��lH6$@���� ��$�60 M��#6 @60 @�B�$��	ld�6$�&�c&D��b�ld�M�&�I����lIc&ēbI����6$�&�I�$ؐ60�&�1$��6$�c ؁6 �c$؄��c$��62M��bI��ld�M��c$��!6$�&�&�&�Cb��|�z���������/���\��N�+%�����\U7ssol]�L�T	�5A,�cN�!d0(A,��v��8lh�w)+��o]�rGrM���=u"�@����Ңv�(.J�e|�(�ҙ���c2a��X)cT�3F�����`��C��hڼ���oE�@��m�ӥ7Qi���4�sU�64nQ���s*�Q�)N�p0&��4��˗y�įK�i�.�&e��oF� �k+j�#N�U+h�6�0J�ϴe�!�ț�P	����n۰�[D�ޭǁ�2�17�]Q&n̙��N���I�Q�%��ѩ�ث����j�Le >��Z+�J����t,ɫEV����(�Z�)#.��@Pu��m���)Xe������h0�ٕ��T�Fn�T�:�L��㵧^�L.LHf㰶���깯^c#֒-1*�E��7u�ЎQ��w	���㡅k�lR�l����1w5�R���Ӆ�Q%�6��m%[C6��o+`�Hu���l�`�7@u�&��bL���j�`e�eէr�-��=+�ᔺ�h���-ܤ��y�0��%�!��9S&m��צ;µ��"`�eU�D�rıR�0v�+7Kv��Z�MhY�F.��b����c�2�[Zv�k�ݶqn'H�f\��J���,�Իų4e#J�jؚ�<T5Mԣ[M�[��MZ\��V�y�u�iQ̮D��}���BҮ�[<�*9�ڐ�]$ِލ������D4t֌l8f6�ùJ���������#rX]nG�U�N�V�spu��e���#�B$�"LC"P��*ܫ��p2�:Kwr1cj;���.��):�V��U�u�wG!�I����H@��3���џ�����`ؤy�E�r�W���3vR��%�ތ��,�*��%��i� �Wղ��EU�8�.P���t�;=nJZT��Ć��Vk��Cpu�5�[��뭐������k%)�
W)�pJۏQ�n�Ge��1� a�W��o~�s1��5��4Skpˈ�����p�;�.����� \�����Z8�����C���ݴv�J�i����4��Xvm�ݧ�V�O¶�	9E^�[��e*4ݐ��j�RvF��vʢ�G��Z����%M֝�z��°��� ۧxh�B%]kB�ǘ�g�̰x'ݩ��}h��[ٸ~Y\�7B,1�����	ةN�֖��乪f���@�&�9�6��7[�JR����
�5�"ۙ#�S
)I0JA�я%��b�7Z�-)Z��<��-�Dq3�Mv���%C���2���9#�@��Ch�n�S���]�mF��1R	:�t�e+V�ѥ�tA��9�����%�mP`�y��[�=�-�֝��EqX�m: =�9v�:��[�V[���lP�7mS(�ye���}��pb��q;_[����Q�@�t�\IC�V[�7ICi���эb��.�QE��,�F��ZS�����ڭ�r�o�ǚ*���!�9��a���KZib��5��v�!f��V�2��V�q�[�8�7G�e&�h�v��n�ћe+^���Q��+c�NP�ò*:0кu�Z�X��-;��&WR�YѬL��`6�;�n��$���gP �ܭ&h�j���uf�F���Ŏ��tl�[F�?+ܴa��N��Bf�D!4
�h�MǠÉ�Q�]L��%�p��
�9���`�X��e�.��v�ai&�A@�K
�;V�����Y	�a�M���ʹ�f�+.��-�:�.R.<�	�0ֹZwH3hS���U��f�-�cX�^�1�`նͥ!b̹%��խ�~����]�!�08�m�E����N]G*]ep�u f,��ڽ�v�(�YA:6��8�-�tY��kf:�6Y72�=��Q(�>Y� ���� 7U��{l�dӧY
cl�"ێ��L6^������kC�n=ɲ�Ь�Ƶd-Y!i��!�������d��R�r�	d�t�E��#�.�;	�m���2�N�̑͒�a�n��fP/E���X�uxfJ{Z��a�cq;��-��̹A�4fށh��(e���x��p��&����e��+C����ږ2}�2�I�si�!VF��kp�u�y���2*k���#v���t-j��!['���b�"�k���ORɒ�H4>(|*�!V�A��%���3��]�Ȓ��n�ϤݨB�'(�͢�̧rnЦfՃ7��y��%e�I��&�K��fġ��̂i��W�hRX�̵0��[A`h��M�v���s1e�Z�tt[���4���^Y�Øn�#��x� ��!��OYj�=/+�"-a,�s��%"*�G1��L�N�_��l⬗N:FTQ���߳>������*��ٙt�Ty���V�3j�ûw �Ʋ�Ņj��ݺw�C7��Z�=YH�FɌd۳I4�ֳgA�2v;��B�,0C��7T�޻��ҁ����2�S�'d�+��y,��4�<o�W\��I�v1�ULY��,ƌ�ʸ�vj��,�ʎ^"g#���+ֲ�+i�����KoY�A��V%�d�!
�2قS�tP��h�h�$�th1J�#����b�e��~��f��ͭ�U��m�P�H�5g��"t/E�+R*eu�ըb3a6��-T�6�9�-��4ރR�Gpİhɘ��b�c��gt@۽ڱl@�Q�E�S5ػ{��B�0D���L�YkE�N��z��cv
6�y0XoN��0u��1��7���G/�XU �/�Q���fK�)�{�S+!�3woFI�c8��9�����TthVXܺF��n"�w��36B憨���$Po�j�RJw/���e��4q�F���ieT0=,*dƄ�W6�OopZ���94������eL6���yW��c�li m V�Pe�bɔM���P�ȷKu�T[�0^�	�C�/.G6�X�FÆ�٦���#����D�f��QY@�Wz�<�ɓn*���0�aB��8��F�T�ALm�ӏ-��m�cJ�uz7J�E�ǀ��>�ڙi�݅��`����۫�3^,�8�: ��KYF��q���GTni8�*�1Z�Y�tn�VK^mI��;���P�-fƦ��[�3+$�B�-�kCztި�vJ��5ow&�N�����;,�[;�)�%�l֙���n��h{��Β�- v�ݍ�Ф
���+U�5��H�xP�����F�k6�e#��҇W��C�Q�镯/3]��0�H��WS$o/"�n}�����U�Y�SU y	0��S��3 K%X�k��u���d��q��5<����G4Qͮ@[wx(�OuZh.-�=ᶒ���d±n��R3Zc��F8�/!���b:�ͼ�aq��1���.���0�{"�{U���Q�p�Ʈ�m�J�o�t	E|���4U)�1и��2�tU�U=S8���ʌ�n��
��NU�e�9Mt�n��Ѻ�
t{Iܽ��+Xx��`��sƐ��l�'NCa��Y�7{��+kv�K�K����x�A��l6wZ��u�L��e�ڮY�-��^i�e�B�dEA�`uu)1��ddãN�.�f e�h�d�mf5���9RD�������� åw�ă�ͺfJ�Y��TIR#s�Q�}z��rL8�*�1]��x7U
�_�h>�����viХ��6R}W���-	0%��f��u%����k"J�7�r�6�q�耓8qhեƠ�n�!4����/�8����;,<�_e���iAV�F�O(`2����t��hCam��0�b�]�#�b��t�wvl�^��ia4���Sk*�D�m`Ee%0`�7*�r]�	dÉL@Qn�F�h5�;9j!_&+�j�;K4�e�{{Q|V�T��zX:kif\�F%WCR�	��IkE��Ԩ�ΌԆ���Igh�Jy�M�FЧV��AU���+/!eH�94���w�\�'-^�	�{�٣�h�+5���h��ݰtK���(ef�� 	hק3kv�U��V�v�����=��>Bе�t�	��h����Y�M��j�`3[.�A&���z�͏T{�)YOLڐ�܉��-��)���q.c�D�=�����pe���]�olh[R0�,k��kc�S�K+o���|�m�T�z	C���,/��C���B�KWqܭ�Cf9�HTmd5�!��7n���tV��6�^#Ե�M����(C��0ͣ��ՖY�UA�r�ܳ��JȲ�n@�Ʋ��5� �����4[8�B��]=�oMJ��F���Y��d�J:h�%�{[�Ӂ��oZ���l��N'�'�
�	��F
�ki�b��{��	B�&��Zl%�+3�8�2Z���l�4�tj��-T��ʊ�BA�͈c)Y[�tF��5,�Iw��,����`������Wcu�� �U��ֶ���mFiͩ���L�sl:`Q8C7Y��L�`��T��	;1uJ���j�Bd��$�uB�]%��i��M�qe���iҿ�^�t�]�2L��Ć�6��2Qj��0Fv�V��÷��n,�HM!�tdM�T�mԑ�С�a���u2�XY+"�����A���M$��l�TZ�Y&n�#NVۇM�ٛ���P;�.J7B�%^}��12���M"Qp杸n�/T��!���`Ŷ��Ռ`C���(��z]�	������*����]�\l�Ӵ�9Z��
֞�M��4]>��m��Yʵ�,���N��i�y���p�\�̸�MMEB�7�@	^�i9ZnPzIV��GL��I��
j!Xʕ7"��-t�ep7µ#چbP���m��]�"�8�9yD-��)��C��R[O�瘈L�X%���N5�T5�6�e��ۙd��%X��օ��r��&�b`:1(nR�\��e�����V���*9�(��(����;�n��vp��/�݁V�ǋ0�E^���3@ۑ:6�&�f7�c�܋#�\wI37��q�'N�W��護��i{R���0he�F^��YUP[��h�/�i�bG�.E	�%��D[{D11��h$+^m�q�9��d�z���F)�SN��4��~�?)�ħ�e��5�L��ːf����Q��i<ikXƗ�����T_2�Z�oL�*�w��$���1;�e�B;'lU���tLي������lgFm�6��i��5l�4��U��3�Q�,��(!��˒-����;�,nӳAYX�+DŴP����AI�ɻ��{�Y�:Vf�TL���"b���;�KnA�F��1�V��dv$n�pX�� 37f&/x'[Su����j%h��� ��k/X]��u=���	!�F^pb�<}��,Gm�<���������"����M�o.ƍf�e�n���F�X&My�m�ޥ�tX��aI�x���sl��V2���ز�B!��7�ɤ���bT�&��-
�kY���I�f���ВKv��[oE6�N�����-
%��/ڙ@-���1�A䙻%���_	K@֛�Ҳ!X[���j#�qr5A�6
�X��kKW�W#M
!q�tqqEf�<�^:�sh���q*�[�\�6�P��GPj��.�W�@����L�;F�
G�8w��G�0D��D\�I��-�(�55n
������X
�e��Ǵ+`֋U�Q�Y�%�{�� m����n�e��'t4^,�qCQ4b�NeIn������bP�)�t���4:.���!̪ܼ̠MZ$^��-j#�/Sɠ�.�ҟ�J��6n��x�hɧ3$�WqKA��[zw��D�9�F刋��t�
kl\�BL�ۭ����j�D�+BŔUQA�\-��-V[ۚ5�-y$a���m��/cݱEإ���0�vʂ���hY���z����{f��Rur��b�c�sdP��Z�]F�a�D<9��ʧ��v��/l��u1���O%3IzE�I���U۱{�á#�)Em��
�L���m�֕�R1�D��%X�Q�ƪP�z7�L���%�����7W�$��P8�S�:l�hbz�H��^�r-��uT�x�����[d��f,��7+yr�=��l�.ܧ�V���g2δn��gF�����[���*ًp�D�e���
�M�f����"�����lH��y�e=��J��l�B�ʘuñ4�XݹFVe��m�(X�A�S5n�qbGx5�2�b�3� F��5b(�[�ҕYDY"=:1��W�P��ؓ�U��p��Yd�����`���A�cT͑Ħn��"rm*����q���ʣPH7���j�҄c�H�R]j̬�ҚoFj�b�h�hXfX5jf<�� ���.\tX"�Jf,ݱ���L�6�[0]`�c'U���9��D�@v��9��x`i$�n���� ��l��ۮb����s��V	�)�괘�N���])�M���f��ď6�n���ǧ��x3sU�V�n�8l����?8���2���9,+iQ\B~K��2r�yW߄�:Y�!Z�޺�&N�=��D���hc���e��ׁ�l.f���؛/��wp�y;Sdպ5���'��l&c|�W��P�:r�r�ruk��N��L�M�2m�eWb�ﾕs�l��M���D &9ݮ�֐���p��f4�S���E�)t�X0㣹�!+��xU�
I�7��/��z'�t֜Z.���Y�O���l�.��:�M/��� �[6Z�4�;�u\7JC(�M�	�G�����v���E2�;Fk�{��g*�J�'�H�q��Ѣt����7G[ Q'v<��3*J�٧�9��$���e�T���|��S�G����>U��>�}P
������3�?I$����^��,M�t=�oe��yN]�t%rT��I��:�'/t�I�\6��F]�ڋ����M2x��y�q�ͼPb�K����-n+W�ݦ���k�H��1O�Qu��f�:iPMC���Eԛz���5)2��5�smV��\j5	:�!�4���eqn�[b�)�����1|��Y_[a#��Yv�����M���=�-�+�v���@,K�ӽZ��I�MqF�-��ǽE\U���8���C�q>f�${%�p�ҪRR.�&>PN��,pǚ3��2� ������l�x�d�w2��5��]k|:��d��yD�ʇF��A'��r���z{(�]�Ԏ�n�䶲S`=�)����)B��YN���f�q�Hi�pT:�]�l\����b��z�{��k(�� �T5̀	�n^�4�wh%"�]�9��N��C�m_J0��1�^l��-V6�˜�0;].�$�;B�.�L8j����=�N�zP[�$Y������*mu�QV��Ō�Ì�
��s�R�N�E�ѳ�`���(�q��0M�ن��}שK�N�1��gW��WT��4b�,#�{˥�P�,nZ��{������8��{kS��d�J�Y�شda*S	b��]X��c�x�v���f�.����BLo�R*��WJ���:�EV�WQ�A�n�u�C���.���0�;\�cXa��e������fוs5�V�eav�7��9�Ip�Z�����j<�h+ă��рs�f��i,�Dn�n�j9��t�lL!�>����뵃^4�b�oBV�:�pP�n#w����f
㺾��*tBu�{.��BK���n�5;�k=پt;E00#6n��qie�<x�ڡ[9�l�tf�+I��2���Pn���`R���U��˳~�fSM��r!Zy�[��
V�f	4U����Һe�O��7Ƒ���{��q�[�V���%P'*NWZXZs�L�8�r�����<2c}pY}��ak��xuے�7/���9��	ڠ�s�z��Jd�5n*e����ZrI{�}:`��< 6��'j��%t#*�Y�����ؓ}��.CI�S�X��4��#f�eܬRR�V,�����NVl��9���q7g]�d\��R���[i�?����s�˜a[�FcǦU��^�$�Cmm����&��ԚpU���h�Y���:�r�5o-噣��P�&hkm�#c��dM�Z��:�X���:J�\�8��Ţ��y�������7����_�u��+��;L���J�,�ɫ&�6�f$�A�V�9�p�h��*c�t��J����a��P䎓��̾�i�˨������88�fe�C���*���X�ڝ�Wɮ��p��YEA��5c3��$��J�vR}vv���_�hK�}4<C���ۥ����+�k����(ȃ�.��v�8�h`Vk�X��� �����:�ng���J�Ϫl'6(Q�쮮�9֝e�����C7�[�8S4�AE8n�+dfu��k9=�yr��� H&��1T�,�������[�u+��9q�-'M�9z!Q��;��Ũ��b�-�B��Tֶ�`�ӛ���N��9��3P�UfgE
X�I�F�U˄{��Z�k6����6'R�7N�K�C�:�3Nd��P6-I��{]�.%��&�՗k^�e�q�2�+s�հ��f��oAB��M7�:��f
4E���cea�E��������I8���^V�����]<�IҪ�A������-�n4��O�s"WAGz�����aJ�l�7��=��b�Ywi5q�2n��w��n�p�V��.��X������1�i�G��z�����' �[u��%)���ZDѥ;�=�j_}�:��|�F�6��OzJ儣��󅈖�2��8r���+B����:Xͣ΋Ίha�3�ߛG�{Z�:+���B�#"3j�Tņ�kB��,Kb�Em��c.�<�����ˤ{P\�G��b˻�����e�s���ts-�V�kά�Z��=��r�R�³�;��4�F��N�1Nل�&3�l�
Gٵ��{F�Ny�ؚұKY�XQ-j����6D�vx��)O3�Re%�f�G��dG ���R�q�\�v��}�k�q�9QƝ:���c�M�[c:#�V�L���ۭ�=;:M:�;ovvR�'c,J����P(l�,�_t�yi%4]+rf�����JTܗL]XɌ�]!���E�B�ʭ�Rp�Hq�2��]�k��5�=��]�&��9�������k�4G6	h�-'H���7���X�x*��`�]m��z��
VAα#����ּlar�Mi.p=�WB{%n1���l"m`#ުU�Au�u�I8N3\#x�Kܡ���f�U�"4(>}��m��"���+��:m�l�%T�:��(�� ���uԆ��YV?��ǥ�Ҟ򕨮���h�*� U��8;W�B8AWhz%�]�ٲPn��I�a�އ�[��B����-T:�ԩ�>Vp+ ���Uړ�sa{���f��ȄV��_a�}6�v�k�z�,(f�KWv�U#R��+����5Æ6�}ף0! +�{#R�p/7-���R�����n�>N�����
�\�l;��+ �C;��G4�aKX��,����,�v��h�9�3)��xEa���;c{� ��4.n�![��z��r�TA�tWX�����+X�(e��0tC'91�X��/�n���'jDƻ�̐��!�Y����m��ǧ��P��� o6��a�W�����yb}��$��J�y� :��}��#X�]j�\�u�U�;��օ�H0�@8gA*��u�Zr��2Z�v��0�ݗ��'���%cY 1f�}�ս+kg�r�G���zv5\e�s\�w��d�
F��t��(	@aۺ)�?*K]��U��P�y�$��>[����h�{ȪWgh.�j�nu�u�D�*�K���{�Z�N��//;52m�Ԝ9,<�g@�XDv�t�t��vP/1܄m�G�p갠�4�>*��%&M���iJ��"<(^�(��	Ys�s+zG+U�n����h�j�\΀�kUU�$6���}�����=�ܤvҏ*v��a�����F]l���2����[(̎�,:��B�\�Av���M��M4�$}�b���d;ֲ�m��<4y�Tr)�{�*��]�����͎�y{�a�U׮`�t�Rh5�һg"�ݾ��� �q�8li�A��ݫ�N�v_U��z�\�5%�t�#��ܱ���O�r@k���ph[�,{j�}������r��0	2�E��u��n�7U���N�I�*F���Kr-�����0��M�|ƭ���=j.Sj���i�t����&+s� u�V�)Sjv��NW&�%��,1�fӓ��i��r�3��M�*q�|evl\�q�xFtA2�	b��}��\�H��gZٖ��r,�]�Y�����n]� ���<A2���r��7A��/�E�[�PK��;��oGq8$�r��w݀smbx�2�ɬj�G+��{ө�{��c:K7)�ߓ���ϕ���,�gJ� N*��杸��~��*ZZ�{V��)�����[uܵ�3gwMA�6�G>�v�D/�<�m�e�|��e��Fmo;&TfB0�ҍ�J1��s��:�8m�ա�J̾m3�x��GN�Xx!28��tԭB�����I]��]��j�e�{y%�H�e9������ں�Ղd�{h�J�[c_ô�y�n�M�	�,t��Vw.�t�������r$�ъpo�����*7�nٮb���W` Y�U�Zo`�a��U�n�Ǜ�.����.ţ�&� �T�j�B�/r��,$v�|�>���\Yb<�&��kp�E֥�X��h%ء�e�E+p�a�[�u֦��f+b!��B�ǅ)]�E��ͥ�CCc�hj��C���Eq2�3d��A�����K�o>��o���� �VuZ\9�b]�����������f�Vպj>�|�U�=�\աJX�p��Wjo�!�=��ѥ[�κj�PGe�p�H���a=W�y�U
��i>�r���qИ�D��!�w8M{�7�-����oM��u��֥��C'�lm�Ks�@�d�iU`w]�ٝD�wkt�ⱟ.W��+�`��Ge`B�oWj��V61'6D��J+��g�-��d��8���'c��H��2
R�;�nl�j��v:�����B�;h��N^��
����詵tk�.:�U�NZ�"��9׬m>�P�V�4�Sc�{3_{:��(Tk�6�݂
�Of�pl�D>��͘��#�6���������=Ŕ3-j�h[o��߳u��ᕤ�שX�����@;�N��w�Ym9"���^^ËF�$��1c�a�gQ��\��u���SrXW�\�Jݮ��m^qw��D��M,1�m��3#խ�8-˖�_tӪ��i�Ϋ��۸�6
�6�0FmV;��;8%�L3F���Vc4nřtO�E�Pb��j�5&�b�f��4�fmo2�j��l�sܾ�$t@P\Bf(m��Y�&E�Qf��B��2��Ac1Q����^�ܥ���"��`���U�cYYr��Wk�7U�V�ć��/MC�$���i��A���:�v
hCn��ξ���Vl���W���2>wԕ]�-WQ��\��!ٴ�BS�2��|)#�z�;��O�W��U�����h�!l��n�Ղ�"���.��z�ȷ\r���������i���/jN��A�����U8 �cF�c{+_t�М��US���=H����w7^3ײf�q�V:f�����V��)�m����+U�k�]ze�ky���}��k�(�ìKC�^�{�E������UJ�o����)5@��]���(�dy�s���n�q�	|zQ��U凯���ޙz���'b8�fMÑ��2ﻮ�Xz(1�k�A�6��
��f[���)MH���U%Ksr���Vz���Z����u�/o�T�:Lr��w�<;�Yصz�(xu�<�[�v��Ok��-��r�	��pp���өË�����|ۼ��]�_^Lԇ5�wd��i��`��-Z$��e�ĪA4>3b/3����4u�Jq#<����a�pdO�<���mD���B���ܦ9�ya��!"$3�{2���9�����v��<31:��Df����������DPr܃�s��Mݳ�3/9k�i�=��Ѫb�J�*���"�<�\��A�Xȋ�]l�H}��WU�p�Iu�6.���evU��!�I[
7�^��ou�Z�
Oq����T�q���.W��|t�y�\���l;��/o�l��2^"Q*���Fu<�k|{D��ó',;���N��5��ƻ��oCW\p\;�Si�tf���R�l��9ٽP�B�ƻ�ݕ�6��.u-q\�B�����^��=V��}�*x��ݠwq����َ��W� �r������e��A�ٸ��S]ebB�}�v��c�����W��"��n���t9L��޸��v��Ud	d4��8v��IU  �⭧�+�)��ÅmҎ 3H5�����;�9 .�k�0�m]��m
jBM`�ͥ��]Lkݺ�L+��oކ8M�oǨ۴$��C�+[�{�l-��ڮ���*Kw��"wj1ϕv��*�7nG�>f��K@e��3�nr3g��<-U�ZZ�I��ײ`yϴ�y`
���!=�he�Ss_)u��el=3;��Nq[�,Z��%��F�k��/��T�]ތ!��/9�lc7�ɱU4�2�.��g��ip��G���Z%ld-��;1ī-�b��+�N�yrg,�,���{+�Z���f<�/��&Mb�l�71��Z����e�\9����jB����h�tِ��i�;{o3�����={�-���))�)�L�ȅv�%��M;n��Naj�O�ˈg<�k]�Ftд�z�+�K]c��qM@Z�܇u�ډ��RZ��G��Q�P9M����(�=V�p�:��03!#*����*0z��#:�+��vI6 `��ipX�r�٤���r�s�'rW��������ȉ�/mփ�k�T�0��u�-��d_+D��w�v��S �H:�g&�c�mh=�ԑ��o&�Rȭ����F*��t���Jx�Zr�Yݝ��xӸq޸\���弰c�ce���Ֆ�c�ے�S�db�%� zIC��b�3�|�љ����[�O�-�k�ÕJ�j6_^b�t��e�w�K���"��%�l֋�v�;�i$[&��J�Vk���K��F,2=;y&t�+e��E�d��J들qV�5��0�bN��cr�ޮR��㈞�,͍��t2�.���$�v�VK����]�rJej���JP
�S8ݪ�Qν�d��%�
�[���KB�b�9�i�5�u�B�9s����Q�����J���j��9��a�NrZ
T�ƚ���u�dj.ّ'*�ꅦ��d�9$���I$NI&�I'nwwR�܅&��#���Xh�H��U:��k%�ʁ���#��j�Q���m���LD�,��=UP�0�$e�R�LQ�B{�<EX�VB�T��C!����X��K-7K��$*����"�40�	�b��@D�s�HY��	h!$	6r	���
�%E0LIIɊ���r�T�!�a%� P��UHU1L�� �
>J+.�Ϊ��{�U`�.�����bCƉ	~�+7���!I��i��밐���~�g�O�H@����!�?���������}/w�w�`�_׌�!��*d6�F^C�ޅ�7''�[%�3�e����7\�'e�B�Yf1�f���h%��7����2��]w��_��ě7J��4v�]6�i��vv	S ��/�ːP��zuu�ӴZ�R*�4-�8`ނ8"ީ�]Ӛ�:���"�<��J��f�3�5Ar��}�^�3dLe�NR���8�lV�gm�
����֬�����t���Ɖ+q��㰮�\�Ԧxe(�����Ũ�-�F��~ͤF�j�N}"Y1���G�[��fG�t�2�j��2�96�
g���1��\�Vc|E��k�o����{MQ��v���-��Q��Y���f�62�t��Z��;\�0ӽ����뇭Lx6k��l�i5��g{����șS����@Ed�3�����fֻ
M���urYR*������8(��_bV6(�	nu`��γ
)�!�XS}�/�(_L��3$G@X{L�;I�r�̍�@�X�)]2^��VZ�
&u���fA��δ#�:8�#�0�2�cJ�!�y�M�����6YeodA5e��\p�أ��3A��]�6�C� ��_,��\��]��V�����T���KFj���M�t^B�+`�ڽk.B����JԲ0'\��fp���r:jp���O_��������_O���=���g�ٓ���{=��Og������{=�=�6l���{=��g'����l�{=��g�������}>�O����Еf�]�y���8��y9շ�e�3��X��E�{hs}R��M��]�Kb����YA$7kRb����o>D���9Ռq���4P���kb �q��ZLV���5�fΚ{Vc�6�P={hI������v��
�J�t0V�0�U���Hu�ǖR�<�����g s��<�uĊ���P�MۡQ����KdδX�K"�	pB��������4e�N�&"��k��P!�I�J� v�Y3Ruut]䤴Żzk^�:y��m�81�(�kl�����Sǲ�*�S�v�4��ڒf����������GU��;H����zS�G�T�����b�"&Tz�#���Oݎ�lUWex3�kI؉�4�V־4�������'^����p����V�HJ��,^��[xtp����Ɗ�8�0����R�\�w��mcϗ�s�5!�Рq�7��GK�����	�J yo�H�9�)�����V��4n%�s��A!��KZdJ�/(F�єL%���˾�B�oI���pjgt�4<�Hՙ�ШJ����'^��-�泀�[YXд��v��h7�X�i�35�5}�J�>�fއ;���Ck+O�e:������%!f�J��n��r�ڒG].��/����wBr�u;�NW��u����i(��x�V�2n@��z�]���&�ϓ��|�'����{=�'���g����{;=��fOg���ɓ'�c=��g����{<�}>?O�����}>�/�����}>�O�4�5�Vr�4�0��Z�n��Ӡ�r%��-��+2��[��A�7n]��3ueV�����>*��R!:�N��\i�Htgl;]x�uk�%iL�&��j)�t�t�Q�n;�s��te��j�%�}SNM(� ����c�(<���3�wZ�ꕲ�ʙ��:VK�al�!TR� z4�6L����WR�pVS��d��.��m>.��i����^�v�D*�Vi&	�R\��JL-����>D }W�ģG�mJ+�@vp��yϰҾ���7d�r�;�>�A���)u�7.<Q���xh��-Q��k��U�١� �@�
����	�
2VN]��9��]Z�� ��ڹ�U��c�`��A����{��2�k�Sw����ZJ��ϯ14dܩ�۷���W0 f�m-�u�ݘ.�[m���l���p�2a����U�;�n_S��o�s���v,���ɥZڳ;�[�oA̬��!��I� C0��?
q1�X���5�0�#W�������t�o�r9N�dj��wgjeÀ5�2և]�"�ro:#)�K�+z��Gq�)�}��/��g�&{���g0�Ϲ�M��u��f��w[W����䗠_p�CyS�X*��?Iٓg'��3��{=��g���zOg����{=��g��{=��fL�2zOg����{=��g�����}>�O�����W����}��]�*v�k���j��]Y˳a֋�:�.�a�i#6P��鉝�e%��i��j�׍]���o���j�9�d �ث�y�l�T��s#�x�B��Op֡D_=T��+�z��]��a۝���`�V�Q�c�b��-D��!{��iǚ���HW����;0���!����Ż��z�Q�{����*i����]��o���t/�'{��Q�e�C���Y*u�ʜ��;*	��Hi߰J=�Ҕ,v .�Z��>+dp��1�������Y�5!��7zc�y���r��I��9���P���-'jv���[�Xul4��↬�Pgw��wyuvj����ӏ6q�s&�i��c-�I���dC��k��莲S�+5�,�*�,&����י֟ �m���C'��ou�s`9������(�s�����2�S�+��}�Jpv��V'̢C��j��묥٫@�g`�y�X��Bvʂ8k�����RL�o��,���}dނ@vwZ��>:\��
��ۇ#S@�p�K�u�h|!t8v��>�Kr:r���)q��&��4y�*��\������c~��v�^ۥ0�n&�Ei���$h�%ԇ�c�C�|�2{��Wr8F\����v@�;���� ͪig\j�,�{;��5��>����|��O����{=��Og��g����{=��'���g�ٳ&L��g��g����{=�Og��g����{��|��O������*
vô�3w�����dW	˃�.��X�Zغ]� 2��9J�����!*Y/h^=��
�U�U���y0��m�Xy!�u�ʗ,��i'	ζb�j����G�
t/8�d��i6��������n�f�ПL��M�-l⹰VK@+Z���r�z�=i����Z�b��':0pMY���{��^Uݑw~���d`��]�^�x/X*ܧT0�*�q�Kpli�c�N4\���jɹyٙ-��,ˮ3�H��#J��#Oe-C���{s���O���cm$��;��#���y@��4��[��F�էOQ΃�AR�L�(�KGF��GÕm%�N�����b�uS ����ʴ����ʃR:��W�b�$�4����O��uՐ֓Nۂ�.!����j�9Tw��n���Q͜��Z��],xl0TF�w���{�N6���U@^G{��#AR-iג��G%��[�f����*���C�+��Xq�S"e@�X���ק�7�{�ʹ1_�x���O��A�V5`ḭh�ܩ�7Mu��q�Љs�����\���i��R�*x��ݏc��̘� �����?U�%����V��p�������:qIeʹ�ph���fP�1T�\������Ҥ6���э�A�B��4�4�ћճ)>Λrs�0��@aɱ���݃Z9c۹�)���f�|�it�إV���ɵZ���8[\��{��phЗ�fk�
-df�.�ճ��b��jԢ2"T�9$�V+�oP��w��ڞ�H����z�3+��!���ת���Z.��qسT�F�V�f�0Ѯ�����6�ѥ�fe����\T���y�Y��.�l�`�]��e�ye㸘��fB�ͬ�-V;81� ����
��GQ@p_k;h��9�U�Ţ2��c�%@�`��)�y��U���U�NC���Ui���v�*�]/����nk|�"�ty��BB���h�:Ӑ���j�d����H�;"3�r���,�0�E���wX�!�o�:�52��D�J�ws�s���7�clu��U�5���^Ђ1�JY��L.;xr�Z�7�XӴ;;%0T��s7���u���ƊE�yR^U̲w&��R1�Be�q�L�EAѿ��K�k�B�}&*�����X���|�-���&m�iK��4vu�6vh}��-�Ju:��X����ɳ^<��1!�]\B�]���wc.��ˑ�n�x���˕Ǖ�e���Q�)��Gz�}(��X��eZ@�6�:����i�0.�&ݑA��8�5g$A9K+�r4&T�0�6��g3u��tJG��U�q`uGW\��V����{�-�v����*�u��"-�n<�-� \x������T0Y��/F�aO��{8�'��؂��>و�μ�tG-�[����	v�gb��G�M���j[7�9v��C�^��r�6�oV��!�j8�V�}u6�J}���
��2���w�,��S#P*ff�K���S��ŴӃ6Zt��X���A�:������v��v���Ǚ/a�0i�:�x5f��-sI@���9l%�9�)1��Q�Y�#�ݣ����_a���h^�j�|�G
Ol��n�� ��ۛؕ����='���Fq�����53rօg:7.��z�7;�b���b���l�*���mv�se�u����M���ب�����*c�Ի��Ԙ�*�8Vn����3MԷ/���@���v9E�d�m���jL�"Xy��%6�6[�g$���!�FSH����3�̎ڎ��7g4���e���B�7
�L��;��!�
�e��]M�E�9�K���_k�V�x�������I!v����T�����*�a��]�-���41nh��g0�[�3������N��%-ۖӒ�f�`f�f�>�����K����v���x6�?B������ik�a�K�q�T�.�d+��N��r���'aR�Y[|���#0��Cͱ�q���9e��vi]z��s%lüd��܂ݕ����HO��{\�L�]�m� )�#Y��VtTB6�0�zછ\�`�77�]��@��e�1Y�4+7�h�}]N�J�YƱ9�7ai�@f,1��J$�Vɏq�z�T�f^���vֻ=�a�(My�TN��2v�����n��<v`�&���J����㭤�*�:�]�\H�7������3E�se��BH�e�T�v0YF���o)GL�x�r���n��(�>�-��ud���&��������qkW;�d�su9\�J0ڧ���o-"lG���GW���M�����q�h�k��i�H���<&�45ݱ�L��y�+(����Z�ܝ5N`�Ad��:��`0���]#���l-�u��c���dVS�w1�`��g��Y NE�Ρ|v�@�i�8��<�W�������/�k�ov?�B��m�)�7�u�,���<T��.�U�35�tu�5K��ͮ:
K���z}+7�X��=��iv��ږs*.`e��u��;�P�_^sTF��GV�X&�PJ��\r+�X��h�]�)�0�j�7���}G`�o'���-���6���ΚF���@P��v;��e��BP7��C�q��l�"��|Ȏ�gN�u�	�Zj�����-�W�Gn�h��j�[B��щC,K�&u,���9�Nx�\��Fhs;�뼝|�Mt�
�,�!�pd�he)b���=�z���n7Lp�(b��t�=��ogF�3���]�Kʜ6���j�Z0U�vB���HgG	I+Z��&�;s�	G����W�Ṳ�y���)J[(�F���G+m�X�f�ϟWڄcP����V:��/��?��73�N�����9s␲q�sQ���,�.λ����:�%�t�DLaɭYˬ��;>�n����XҪ+4���>D��h�&����gf�o=f�鹁��C]�Gp���^:6�HOï@��ٜ�.�(v&�b�L������^,�_Vp�/-8M�	�5=}���13�[4��2��*�ʎ��p5Кv���l�q)�r(H��άŦmu��{4��4V-�*�(���C������ȩSD�h��vuu�I��<}v�ٿC1CG���ԛ�P'��?�B��Ք���o]С%$�,	ݔW�D��av0A��f�w=�������ݨz>�8P�*�8�N����,K�������^��&�b)NG�6���A᫓��&c�����y�i�t�����pV\�$���z%E��5�-�V,/o$���N�8�8빸^��t�l��Z��7��1�l����4�%�b��B��L��N�dM��9�2\j�Ζ�;�J�[��J<uZo7p��y#��鈁E��:2d]X��)c��V�G{�&����fo:Y9�^��Kͤ��j�������͙ٮO�*�Ǥ�":tF��u�6���x�kn�;O�u�h�@��5vI�rf�t�MV4�a��֘��<6�7Ӯ2��e���cu��s%Ι�Rq�.�ͥ.]e��,�$Dŵ���z��ۣ֜��39��,G�N��C5�֞��DI��.v�(��T��r��Ŭg=u��;J�6����n�c2�+�����	`m����l�Pb�g(>�tN�_��崘
�S�C2M9+hGN��6Cu�%�D��姽�b-����6�x㳉Y��]��a�í�`2��1��KlI�)�C�e�Ea�kr��&�2P"�F��i�{q�[+�kT��&T�f�;7�Շ���Q�b�0�
�jN����N�ݝ��RĹ�/gA�n��Ð�j<뫒|p��af�I[�2��^�p���yދ�[J���
�CҰ�0�zZHše"�����L���l�u!��kە)�60�҅�gpu]��&.ٖis[J�KY1Y	?�8�y&��7.�p��*�O��x�2�b�:�;���V���X����KQ{t�_8�ܑ����\��[�h��BȏO6���tPb��հK�U��-���[:*�W��ɱɚ̧�4�.ɬJB+7��[��vȝpN�:�R���@M��R�
�#+�;؋�
���>x�+������$�O�Y�?^������~����~��2��ҋ���ҙw�W1hMTA~����\���H�l�Xc�r���ݽ��ǽj0T�"Hq�R�s����1��$��֚����(y��S��q���Y`�ɪj����<x+�u��uEXg�H`{�X3O�AX�����pZ�kTaT7k�]����]8�l,�F@5��\y�{	Ѯ�4*P�Lvn��3 �ǐe�t�-����˔ݨh��\F��RX�[V�.+��)�$�������eK[S�������}��l�N��v��d�����N�f޽ҩ.�Xq���Z�RH�&�����X���*������P��`�P����D�]Y��D�9������-�p2:_Kek��pk��D��+5��w��/)����n��۷��.+�:�\�[���v�^�t/�o#-Ԭ�rP.��v�Î�;�n��Υ������dU�]av�!4�$�J�6�W[�ϥ�v���H����"�{H�G�L���&s]m.�}k3�'ϴ�;ȹ���Ռ��n;��*8�������зۃLr��>�*�(.��kw8�|�=�n)R��m�wM��q�0�6�F���)��ΓӉ)���xQ�S�ɔ6�o�m��d1�Ze��2 �����y�a���7z�nnl[I�5�{C�&�\۹���v�+\��8��1��p��nU���ܹ��Af2�4�1`���*���G��1;B��H"�j6���̙9>N΂����KX/Y��a����yM���C�9q�\`R�vاj1����N��w�SQbֵ�R*̵TV�i��*TֱI�ͦ%d��ۙRT=L�NaYg'g���vصT �Zʪ�>eƢ�,�3*ζ�LE�O(�*�¹h��Jl��vt-����%b%�!�p��z��X��(���py��S��Ϗ��[L�V�g�5���#[hWLa_b1�������bʎ&�0QE��
-��k���N!�J�8�ec���8�;���YFG)v�8�:������Q4Aj6�Jŕ�n��+k(V��[Fq���J��T���V�ƹe��Z��ULj.0�KKeT7sh�YYPn��TY�K�.+�3M�Z��ګ�U>�$׮
�yj�yJ�Ƣ2�i[�g6�w,� ڽ`���	��y�2��~����|O��qѬ�N6	�p#z^q�N��l�w���/^��Ș},�n���.�%$�/�(�T�q��8�����Ź+����UG�I�]���5�3��ε������=C��r�}��㔻�~��zm�p7S"!}���������3��z�ڭ����&}��^y�l��^����=o����z�b.$�{�ɡ]��z�J��*��~����d����Wq��]���!��ؽ^�4�ƞg;���l�u�w��O(f��f�1	{�/�{�N~���?/n�����G&esF��#�x�׵OkC>�E��Lx�M_D^�g�^��2x�_�y)^����a��e��N��ί�i�G¼��yl�x
��������!2y�}^2zue��cQ G:��z��9Z���{%�SOH߸�k�j�);������<��w�>�������ny+-b��z��Wpf�_W�&+�u��+U��߽}����}
�jy`����g1���ub�[sM3yW`J�W�̴�^b�t���S�*��өH��e�n=8S�V$
��#z�ah�ɝd}N���;��{��yKR$9N�ju�$�r�4�!�Ch��ݹ�^>�;��}���.��Ǟ�:���tgegP�Sc��=:G1W~��{����.���/COgvx.CR�,�&�̭��Oz��L�=>���l�wP=?o���}�,�po�Q:Zn9���1�G�'��A�3�J�¯G�ʙA"9ᮯC�~�,��=v7NR�rt^��o�O]sn��RE ڿ���>�v�=��NV< t�l�v���oχ�����y�x�d+��^����������6ħ�����6;�1�=�t&���U�Λ�/]�7+��ugyFpd3�{۫�p��ѫ|=L��ާ��m���J��Ty�Fk�ϳ\���|9s����[��oE�����>�k��_(��~�~SvS��,l�"�o�pvڛ��߱{]Wb����8s�����^Y�:�Nb��U磏/�ҟ����}��&��{״^Γo��N¬�ƽ�kt��f�hc���I=5�"�M���.���k`ɮ8��:��]w#�GV��Y�`��c�;#ͦ�ݽ�bun!&�Xs���uo�����`
LYk��c4�ך�fu�&6���jLZ��N�1����(���:���Km��0��Ӱv�2@l��Uo�dώ��t�x�c'2��I�;�A��l��&;���ܤ��ZR�`�7�|��Sz}u���\�g*OOoʽg�h�ɟ0:�d��{c
Ww���U_ G1u)K��~�T��J�w���)[;	6V_�9Y���]���ჳ��+�_F=9Y�q;�y���_�k�D��g�z���|���>Ԇ*sC|�N��
�������&Dw���(�ଛǠG��>�_�����:<������������T�As�	qٛ촎��N�8�{~?�b|�����ɟ3�^T��>=�3	��W��q\_�R�@9��]]���Ss�ߙ���]�o���иM�3=��c݉o����oɇ��'[�ƻ��!#T����1 &f���B4������=��cݴ�̥�Fy�O����r�Z��Cm*�7^W�v�� �X`�q	\T}Y@>�0�鞏C�z����.�$��^gN���G,�xF��G������E�C���v��y=NX�>�Y��x�i���X�B'pf��t�T����vq�ٗc੖"�Ac���]��Y���5R�Lճ/���9|=�2��~��/�o����s��s��:Z��3�S.o{s}lF=u�+ݓ��//s��X��D��Ɣ=��C|�˽��6H�_K�/���Vb�Uu�>�z��|�������;@����fͼ
��F
��LkF�͞�g;c�������ao(;��T��߼���v��t��p�o�z���;*�?f���y����_�?R^������6�w0�yᏵ?zм�'b�G㾪o�(�>�2�]~���}E����_:��U�{�9W��PX߻�}ݘ%��0�~l��z�^Ї;#��Ӄ�W���.�`c�~�>�n�=����������˪�}�u���)��c�Fk�4VM/э)Oo'�Ɨ'��`bs(湟Q���q����ly���.9. �=\�3�;AW�tЙ0���������ｶ��sz���N�*E���:�+�`���(%W�O�S�K�z��/�n�K�����R��]ݞ>�9u��`�Qm"�V�ݱ�Wvy=��G�Îs��3k{5c6��i]7�%AdU���2>�����q�+_/}B�ٓ��x�F�a� �R�z��B�,M���ٯ���g�H��xR�չ#�5P��}��<����T�זt��Y�*��߇��h�40w(���:f���g*��Ҳ����ҁ܃Ԧ��6�ms�gUO�"n�>�o������[�,J��=�:#��w��7�G�A2�c������ڱ��O1��7Ǟ������Qa���ed��Og�@�FH<�rvݏKW�����[�y޶����b�z��(�-�{�M��^���G�\^�aꜗ9�%�+]�V����3�{�J/�� ��.;5�^��̝�^[<6�ޠQ����N
N`*�q󖩪�[�S~�_<�O�޵ʹ6^��ڮ�eF�{��K�[���� ���z8��޼��~�,q����kbҙެA�N�#Ml�� 1�h�;�f�mg궸�+�A�x�cG�ϻ޻\h^7@�nA��i����i��h��.Kݹ����5�֎�W�V��n�Qq�ˬ�ySj�� ��(�-Hٝ�O[^C!̲+�/spA�YN�u��!��ggq9}��}[��(��D⏌�����:�Vn1/�0{���n�ֳoZs�F.�]B^�<�9 ?m����\loF��t�6�N���I�r�1�vY��a��!�gPً���~��O:��ǵ�N}8��<�op���\�P[�ɭމ��$ε���c���U.�ݨ��Ͻ��Oo���a���R�n��b�u��FzWx*ϸ������U��vb	�S~�}��=��e
̾�>^1�6�ឦ���V�d����A�az}���Յ�%�T�����:�<.VvwM�H�elc$t�t��}�q���D
�l�:kD�r���E]y�\�e:��>~�t%���q�ʗ�(M�"9���.�j����O�MJ4N�q��͋��{��m�'�+���ϥ��;	����w����|��g���^@h��QS���,Vdp^׽J��K�="��� �c9��)�����s`Wd�K.PWܘ~����ek��=�A�^�Y��w��N���ӌ�X���2������x�n`	6�� �,�M\�����n��V�+�|��s�T�[6Ɯ��Svy��׈���ocՉ=�uca�u�jEn�nC�<Te)n��ͺ�,�B�ۑ;���ݝ7+CWӻfeL�R��gw<S~��g�6�>���	������k�9��F*��Y�Z��Auw����E�ޘ��u�6�s����{�Ǟ�B��b��[�x������'�����y��3gKP1@�wM"ܣ1������6u﷠�S����=���9��I�}QgO<��b�v�zx���!����C��F�=A�����]S�e{���^�Eb�7=�W�/��)��{��yr��i���|��$�gjz{<W�������Ъ��iN���=D��ِvt�vb�{�OvA��]�����y����v�E�l�t�}���F�{E��� V�|<���W��n�1nsc�32c6^���ڳ�Ϳ�㙣�Zcg��w��4'�ך�گJ�����hÄc��is�`v�z�Q�����c��{�Z��㑵\�rj�Q���x��UeiWQe���k�}�yK������pS\*M��M�ngV���{�V�v!t�
@�a�Ec�,#ݥ� ��er�O5��N`N}��%':c����XN�0x��z�ە��Y[n�D��RN�`�ZKi�JZXv�s,�]��M˒��wg�S�w;I�4$��9>�V��ʣ2d9FEK'-���k3u�Ы���[����g��I�m���'A��߁k}
�����v���	OzB�����������U���~�k���$��n�d��<#i���%J�c��y�OH�����(Y�cf�=�TJ��+l֩]��?g�l~����	�O�Eϰ�4�x�k�bZ$>s9��3��nc��8}�yYX�kP�R�����ޯ��z,{�{%�7�%�\��Atxj�7��j�_�'�Wg����'j̝��Y^&�6��C�����B���{�x�~����3�ߜ�Q��xU��߼���I�[�t&�vT��7�'���z��xc������\3f���F����3���A��ug{�H:�ɫ���;�LNls��-����W�1�u����J7�DQ�/v���� ���v���v�X'i�+����Ҏ��nEY�}�v֩�貭����n�7\^�Gz
����s���'{BH�r�"���d��i�y<�+�ͼ�!�)�V��9�����C	"����5Ye�+:>�L��-�{��<G��g�>�9���;���W��;�T��<[�ٿ>��ROT~ყҪ��WC��2��P@����>]���o����<_9��V�3��{<�^Cʩ�l��b��{�ْӯ�ʩ�v�ߖﰸ>��I<����d�g��u��蟠�Dﾟ/_Ƒ��ikϷ=1�UC9l�EyJ��pq�^�w+O��=�1�����"=	]:���ut�ߞn]7�퍩v��z��nV[�i�<���=���<��sj�}9;�
��Km�|{�V��g�'�lIK*A�=��Ω�^�j�F.6(}�^�Ko�e�UyK~+$t��1���2��{��/���/�E�7��y=�e����^��
�;��G�������{�M]׋����Ok
mcV�=�Τ/�/Rd���Hu��j+=S|a�P�mz��w8��.�TI�)�Α��F���	M���-lr�
ۈ�Ԇ�{���Q�2��s�zVu��0�F\&E+��e��v�І��-S����sL�m��i���|����ǁ����>�8X�W[_5W9};���~�)�I��j���y��3�U�9ez��:��i��'���Y�fS|j{�W���&������p��q�靫���K=���.O:�T���b��r��N����s=�W�J6���b�=羿�n�����Mp�j��*3�VQ�̖���ז�m��SA?n62������T&D~����^BE���l���}y�߶����ԏ�����x���y�Bv����o�z#���Z+|�p���k�9e�i�����D=x�9������M�{׿yO%��Ώgq����1z�-,w�3�4k8;�#���n�����̿k~޴�;k�Վ��YSʲ���X"�9eఽ2����,���C�g�`z�H�g�����W�����O��p�->�i��~�B�M�JV�M�x��BN=������ڨņ�L�L+4�i�*����{�[�ʹR��7Y�]ć=w��W��J�n��Zԇkr�t�)�O���vN��|*pq�J��3vֵ\�xfE��Q�2�b�fn����B^hTgǡ�.��v7hk�Q��q�ŧ2�rZ\.��zp���gw0�C�Ϻ(.z�e���Wz�x�PN��\ټ*D�ܳz=�9�x�Rf�rZ/���a^αʸ���mn������B	�2�\RVO���Xl����4�P�����w>�
8��e\����,&6hL*�ouAL��a�d|÷3���U�QVf18�.>*4iзʥݥ:���f�W�8�����w�����d<I�(�Wq��r�A�� � մ��*�7oN���'M �T�NO�x-�N*eg&;��(R���<�����Ś����`r@����C#��s�����Ԙz�g.��:��9������[�gΛ<����S�{��S��uܱ����9Ս���*+6B�W�fĞT�L��c��ɜ�pT���he�<�3N:Q�mn�κ9�n�-ʋ�ظ�w�H�N��B:������t(-c��w�c��r����d�@jK��E˞�P�t�YW57;�)��Њ� 8o;#ո;"�緼�:<K�=��4k�8�����A���l���+����KU�y�A6.���R�y��1��#e45S\�;��;}�u�c�Z�Z"��$_R���ao%*Uu�� &�t{���y��9L
ҷ�eȷK:�\�r�Ee<w�)�sX��I�;z	��뾑Ѡ�ļ���!G�^�#�s��{)�v�F�n�x�j���˹]�fRL[!vaW�f��m�W]"k!�9�%�Lh�MD�hR�*� hs���f�L���se� ��X�pCI(������K�\I��.X�X���`h�`�f��V�MXZ�$������u��13\ßH��v�W���]Hv�tl���_��巡�r{�љƥ�[�\�����4j�v�A0k�:G{P.�ۯt�:�J��@���$t<�h�ΉQ�L_	�KF��p
��Yk\�c���M�ś�Nj���l1�,��o�x��&��ũk�C
ʲ�e>�hoL�zz�`�`I�x��2c/r�X'�锱W)��Ы�*P��oYwE�-�wZ�x^�n&n�䵉��s a��|�(��s�s�B��P�zm�1�r_�΃(&e�oC38��2ުR�����-�Li÷SM˵9;ͺ2WK39�ǈ���-��P�8����N���ѝ��K�·Z�z�L���Fw�qU��Y�jmЖ2�u���X/N�2��\	���&zf�'�<�r��d;D^�;E#F|��.GYi͡�;%[���>2bӻJ��l�i`X4jUz��>շ֖%�kV*�6K����7:��6�Y����sS�۟x�@�G�M�� �F���d�X��<q��h�X��T��Ȝi��B�L�<���K���Y�e�k6�JZ[Z'ndke�X��nf��-o�`�0++.5Ls�bgݥ������9;��ǉ���+<LMJ�]t�[40̥�,���Xњ�r�Ȇn�+32�^Y�:�''�ggAb�,��b_)v�)v����$LuƓn&�|��Z�e��k\k:�91�J�JfZ3�Y�7����������Vm�A����(�,A�LC3��#e��i/2WU�9f��aA���ae���3-�Y��Ki��2�-ȓ+��w��p�0������S ��fJ�z��ڒ����U��C0�0�%��*�u�̆,�<��KmC0m�,�3�]k5ɋf:�#��xh�l[���s���r��e�e/vM�2�a�T�5;y����T^<J�;i�9�9�����9��1-�블F|��83�v����̠8b�-��㙎#Z�|M�eJ��{�{�`��y�F��v�q�n�(�ܻ��-�U5-��֪
��5�,完���e3L%j6��|�̴۬AL�
r�moy��2PX"x�i���/.'�Ϳϛr���efB����}+||�n]��>���E����N�Uy(
Q���u�b����W�H͓�C��+bYq�ꯥ}�����u��9f.��W���s1{5��u�V����D���s�'�r~��ZgU�z���U���44oG7�_�>Q�͋wy�`����Ŝ4��m~��@��'���<�/2�7`�t�G4�~�}o����׆��<�F1̏so�fU^��N�^)A���N�^�WSF�1�Ng������/����\
���a�k� ��9P�W<�?'�e�_�ݝ ��{jT`��r�6Ѝ��_�����B���0���`OF`CߕGG����MWW�w�S`\�o�R[2�GR��+��>���M�̶�%�«آܸ�u�v+�I�q��ו���]�߲ji�DJ[�ʢ~߂c���x6�tW��>j�N[�\/S�x*��U�-��B��x����P	ྨ��n��?[��v���G���k	���yŇ�4������Y4�[I��x�M��w�7�SZ�!/�~�w��	��i����'�~f�}<�����]1`���M_�l>��f�1�ur <�v��xd}�g��z~�����n>�%��z�!��x�V�~��0����0H۽�uf���{r�e�KF~{�|���It��~��wtH�yZ�E�g�J�v�	.���NN��ORF�u ��6�m���iK�+ڱ<�I����)���T�_Fv�V}/�nL��e�T�EU��Ф36�s5��d��eo__)�Xf��n�D��mo�Ա%�dj�mG޹�L��y���|a� :���%�?�O8;5P�#��|����s&-�m��l}H����⼗O7����Yq+����1�����G缀�y�-#�WB%�TI͌TFHk�)�H������-l���+�
;@��O��ð�5��o!����ʬ��Zϲ-����^݋��G)E����j�Զ��MV�q��`���R�gצ��3koiWO�3pm�vn0���X�=�*=c������۹1�l�3e��y���L�aU�=b>�}�'�~��6�P������c�d�c�n��1��A�	w-L�ĿA��U��5��'�v��~�W5�m	���ߺ�Ǆ���w�|OCQ�ۗo��Kz�\�p��K8W�K3{��E�O�WP�(͟D}c���h�T����*�� Z�Gᕷ�ˣ%��l��B�L�о���^���`CT۸(ͻ�=v�c؈��M��x���~jUZ���U��F�ȳSl(��E�k�`�f(��+(V�*�Ի���ظu���}�v�!4
2༬զ���?�G��5�=�`��C��{>�G��>�C�o���[��%ͩRM�JE���q]��`����FMםv�Y�t����:�AkB��N���	p��0���� ��f�A����Z�>����2��4P$�H���O̙���U�3)m�������U���O1�;5����2�Z�O�nEaR��u<�w��^)�|�u��a�Pg�Y�3��� Zڏ <���E��6u�<BO��.V++�����e�(=U�M�N������׷}oci�dC��˳� ��p�CuI��yi.�y�V�~������ѕk���<S.~�qT=�,�#��.9j�&�ƾ?r��/ܨc�)楉�	UZu�ZZ��{J���9��[�v4jP��yӾ$^=9,,3o��Bn�^��q�\=71e0��"��.+�-W0�Q�ɼ�L��ұ�c���dZ����Wm��Êc���M�tO�vx��?������Jm���j�=�"��xR�Ph�=4(.�MY�K���DJ�	kd1�`̘�o9�ze�!�}���n�[cq)1q^��\@�j�0n!.��9�4Ի��('��xܱ�����Cϛa0� >��ĲcҧX`�k�XŻmQ�C��SC�St`6_a�Q����~_zٞT"?-"z��][�:��2����>d1�^dk��H`LN��%���c^�u��,�X融��~����3�+R������h2IuL6{=|8#.�9�X]=�L�m��8�َ6���������h=]yK�4�95,*9e�($����_��-��2�������p;z���n- b�B��T�p�^��k9��y
E���n�_��8�`*���Z=v�>c�'1�!��i� ��(ͳ��t�몈���籛GS�;���ꉶ�\��2h��ob�����l��<ܝ0�\!��l�?��F��t�lÑ׬Hڹ���:]��~����ʒ�F4�Hfٵ*�`�q�$R���*�V<�O�v�uL�jm��k�MYD&��G�0u�M
R�j�L�A@*FD����U�}�Y9Tŷp�OGx���\^׻Mk/08�]7������ �����;���x\u�70z�!���|�����1%F�m1��6b�VL�;��2o8�m��]c��;]\�;ω��NE�C�NM��w��b�32�� Pe��<��v��S�W�Uk��'�I��Ƣ��f�|�RO��V�{��|5ry ���Ulm{#�4Z2GgR��))��R~k��Ე+:��B_)�F5�3����ʰ�/�wL�D�5���^ڗ��/^D���ܗ\���v�%��ÔOW�;�I���珑|�����@O8�pLx�V��8�䌫޾<����_*�5P�&H�����n��^�m��V����e�$nDx^�lfb6��{�6d�d=YyP���k�^��W��ܖ�d����^|��t+��Z�����:�=/�Y��ͦi�=x����%%[�:{A��X��u���65�y�u�Q��%h��V0N�CA=�,���_/�,��lgMQ�}s� mF�3�E+��9�Ӗ����V5��n���ja�9ކ-�i�#M���%���ݩ��!7���*F�lj�Ϻ{��h���v�y�t�'���C3���n+k�z�(�����m�Ca��HPSײ����Hv��������8�ƪ��S�"}�B�d��jN�u���5�C^��z|Y��'+՝������M���1��i��%M��[/��!�3��57�����}+L�	qq��qΑ���c����˹kx˶� �l^�nX�F��F�<���K �v�C�ݺ<i�U�i�,ч����.���Jk˺����H�V������RY�ΥsC-���E��w��W*��P�#%�"��L/��ޑbSͨe\�k�M٦�=�y���!H�B�̌��pU6�1�ߖr���S�0c{�7��"��I�=z�
{������&ƶ�Ɵw6�|�[RYZ+���I�p�E�p�w���;�RW���4��ocmYC�v���d�ǱÝdݪw�[�1��Թ>�rγiv�M�d�� ��N�	$Ż4�`!�����m�>s��V>�4>����0UkûG�kށ��蓏����lO(��h���߯�X�;��J�݉U�t^6D`����<���{juK�׀�!��k	�������TZp	����ɦ���.�m�0���ȋ��ͶW�6����԰,�4� �T�6����Cn�<)�;.OLS�9�Z��`jy�3��6�?5V������$�$��-������-3���������jCjj�j�uW����K����B9�\�.YM�`i%����;u�@}��-	��痾��a.kjeh���k\2�m�\e�r�Sߊ2Yn3�X�Nn}�d����f��Οx��vF.��}�M�\1T�^ˋN��Nx�0����1�}��sz'Ga2��`�˽�a�aE��c�uk-����vt3T�y����I���e��q�41�t�j����Bs�Q���O��XD�o�q#�WBU�6�����T������<_��ގ�
G&ghT%�}8�x��y(�ܢ[�&���i�b�)��7Cnd�w�	��p���C1��Xv(^��T�5��qn�5���C{`�|[��yOJ��N�`9�33����n��#�=E���{�5�F;�S��P\K�ͭK�hp��j�c�e;Ιw܋3�Ah��+;f%�3f�x^!ҷ!���ű}�����=7��ڗ���&�b��y���$]���gS4��Uq?j�"�n��s��GC���X��Y��&���`��{u���LF��
��<��:9 �^@u��g�s���˃�h�\e�D���>q�s,�$������F<��G*���U��0�8�C.H��p/]0�T �A
��� ��� 6��<};8	�)[Yt:<�s����?S��9��Fv��J��΃(zO%րVW�m�U�)����'0}��}:v~	?��h;�TV���-M)��y|2= u�|p�����R~��"�4���۵V���X�]����E^�l��/��,�5�(K<҂8_��4K�(cm@�F#fZ)�FM<��hoX�z��7��K��]舭�3�E���?v1�k��/���_pp�E��ݨ���M�.ҙ�?�$z�yN�(�*�6g���#�:tE.���PZ\s�R2�l��4���ܞ�消�������,,��r�����X_F���c�:@��8A66� l����^�56;!��&�#�)�y��kuR�^�V��BX��2�`����Xo�� ��t#_�E߫�]��˽\�Df�vZ�������E�@�`�Yd9sG��(���b�G��՘i���nv����6V�'L�؟��-�آ�n�R�$�u�^�{�������Ï���nt�m?���s�=���@���1�����%q,��o��7W�!9jf8����ٜpf*e{�6�=Q��/�Iaö�L�Ca=u��Z�4#�q-Av�2`�.cyz&_���S.��,<O{UB�kۃJop{C�����j�w��ƬW�&F�1נ��s��FCA;Ō�tz�_U���d����X�eB�zX^����M#�1��V�M��Uy��եr�=SI�`�	���~h�?y���zGR�[����)Da��aK�@��:�t@��qe���}#��RjnA?��ϟ���uJ����pϟ��.s��!s�e���i��,�wpD{1����!��-"ĕ6�������J_�����]f�92ӱ�Wu��0���|��J``��W��]Cv���^��=��.Ylۖ7�iN��y���@�����|�D|24sk��$�1zԈp�q)�b���B-J���ɾI���L������i�r��=;�K� �6��L�ܢ�=�=�
lo-#
M;U���Ρ�z���P��MO�W�\���d�2�&�Ļ�BoW��d�Cx��C���P�m��wh��ڗ�tv<��C������ �Nƻw2/�֍���J�!��S���>
��L��o)�*��n���V��r�y�X���4�7b1�p��ֻ�'b�e�f�������8����6��6v�w�x'�����/pH~D213������c��M�֠[�z:d���MIe��UL��ƿvy�m��
��B���$�|�-���z�cEJV�
���D�k�s��vߣM.{~�'�f�R�v(���Q�q��T�uUr9/h�l��h�s��mk �^K��(An��@L��wE�RS�����/?7JQ�Y�y�D�x�����ѷ�[�qi��Ly�v|�C���>�q�e��(��rެ'+�(�\�;���wqU��e�ʈ��r�NM5�%$���N��[Yθ5/�DD&޺�`6|7���T���fx�uZ�ʣ�z�0aP�-�Lxϴ�Ghy�w����_������@W���J���6+r��8�?>�S��#lq׻�l�uQNy�u�j��SƫZ�"�w���O͍-w�CW�@Ȱ�n���֋��Z�ֽ���(sv��7���{���t��=�P	�>���ʹ,X{�\��ʥ�P��j�C��
az�g����25���:LA=#�.��3�l��|j�����Zx��������=,���E�g�t1��;lCO���7X��%�`�H��o�ErlCvE� I���Ȭɛ��,�ck.��"������x�S]"�dg�j��Wd�[�g>ݽ��Y�4�3�H�T1�%����7���ۉ�Y���{��1oH�Ʊƪ�}2c�fv�#1��8[V�W{�]�p��ߞ�_��I0�������E6�d����T�N ����0S��kfX��sNdKCN�q�iy�DzXE��"O�[.�4�[�y��'�ʒߩ15B��N/�,[�G��U�GU)<���{wB@�y ��ؠiy�
R�+A�֞��4�5�\���*EЌ�Mz�_�K��t���ŝm@3�]���A�M>�X��VU6�d�pUb�r�(�Z��&��L3,��﫺�G�#B�v���]���;z�t�t��E'+`KF0*l�߽V6���́���4̬�]�y��mܚ7�#ϡ�Q6+ѽ\���Q��,S����-A5��/k�3Wȩ��ђ���4���$�.�?��L��z��9^��3E�W3�
�p���p�D�]$"�y�fm�cz�Tu��@@"��e����h��%� ���h�Qp��U�dR��z����^���f�;�v�ڞ�����`�La��`�r^S�#sֵ[��4ePڭ3���r3T4��=��������6�X��$�k�k����Q!�J_���N�{��l��0N�雖�3����sV��n��q\�'�N.��X��{*MT�k���4��t�&��핹ԬY$W��\��/l�&�9ue֫+�e�QX 馱32�04H��.d�I쾓lL��3�>z;,3����&8�2�n¦˴6Ȯ�U��HD��yU�Yn�tHӒ�+6��_N�J��׳7������ �f��hR�V#���Cމ�3�����ƙ�V�\��执@(�Κ��sd�zjj_bqk�++*k�*��f菠��3��2�V�ܘやV2%�Z![Ԕ���M�5S5p�����=�k��I���V>�U�����8 V�� `� ��.��r�z����$�j�
ë�ulC!��tP[��e�*hT'R]4�����*CyA��!�4^V�MJ�>�s���7%ྒ��9м����j
���r,,Z��v�*�]pD��C����^��^T�\�Io/�Q����6غ�Pf��D���s	ȪE-e�I»N�i��2l�Jɼe�YU�s0����l��<�XK�Α!�u_:p��� �^9�s����4��W
Ӧ�yR:�@���A���a��*1ȵ�ԩ��@e��a�8���z����{ԟ:pF%ik��ށ��nF���鿉�f����V�s���%`��c���IvK
�&�K���R�#9��͹X�ȮrH�B���A�َ37�
���m�0"V_v	����Y��`Xl�4�o���5���J%J��0��tW�����N�be6��0�(X��-PW��Է�=��h"V�`�\f��)z^�����Y#���ۡ�.M����)^G���!\�f*|���R�f�e�,�f�ⱔ�p�����G�5*z���U4����^ML�E�܂
�;_����]��4�Z�CI;'"��&���g^iU���h�:����Ɲp�e���COg����6���\Lt�E��?�K����pɒ�4���o�M�u	;Daս�u�7������syà�e���x��[؊@c�.>�B�A�Z )�\����E�o��k6�\:��NY@N�2��06�R8^s�!U��#L�Lf<c-U��w[�u��'�dl�olŷ��Ӧ����t���XIK����WR��h[��8h����l3��@ѫ���e����vyA���ƲC���S��q��v�^+(Ut�O`��Ҳ��&��V�;�b�gf�S6h�@6!�pyM����<�v�K3Q���б���Mi�E7���Ī��u�;�K��k\Mr���l�8�p���s&âFEo9�X��5��gq�	�)K��˻���o ٹ]z)�tn�(��i΋�k���Nƫ�9)϶��1�7y�ujoYW�^	64���4{���R��C�[�
�-X7#�ձ���7|����\�i<Dy xr�D��w5�����Ri�z&�0ѮH�?�$�"*�@�e�_m/�Q�aM�A��?'�Pr��æRWsMN���o���!�)���y��(|N��i�l��"7�wm��|s��PL��nw��'kk�ٳ��rt�
c�Y��gob�,3��V�Ĩ�C;n�h���E*jT2++#�+:8��r�fN�'����kr�Dm���QQ�ZUkm��E�X�,��R���|�1�U�Z�2�O'����|/���rs�Z�U�8�ݦb�VR�iuر�Q����)w.[j2�Ҧ���g�����3���з�1���X��Lr�m,jV�U���8��*�Էr��ݛʍ����rߛ�chӗ��V��Ң6��*
���V���	[KJX��Q��S2���E����=�`��l���Lk���b�3YDTEʶ��JՂe.k�Tw0-
��� �T�.2�qV��[m�~���CQE���i��Z�B���҂�2��[F�%�iLWmr\�.jֵ�-�*J�R�-%E�DB��Qb�n�2*���J�8���EU���bD�B?�IP��J�cQ�/+�~��&��T�Π���9m��&fpܧ؋�{ż8��u�d]�u�:�]ܵRCf�s�ܼd�`�=�h�J8���B}��HH6䬖�m>]p��/6��zO>3��a��(6R���ϩdx�oD���s@����2};=.੻�ޑ4��������aY`�;Ǆ�n�y�(�����%�U~�v��E��C�I��u}Q;�%4:��ҋ]�@@v�ȃ��X�O���E���e`s#�{Ub���ﱡ`r	�ˏm �h�)�Xdx���,,��;8Lѯ|]�r�����X��YZ��&4�Ȼ��9ܘv���>5�迕Q-�~LMP��9���OCQ�͍n%��FI�x�	����sÊ��œ2N�¸ҩpa�E�_�H��y�ّa�e��
�}��h�#eu<4�ewNgMCP����ҥ����K!�_tę�K�P;u+�	(;Jk��ī��{̔����,T*y1A�֔,4׮�'9i�R��ڦ�H�{������Tկ��l�#�|Ű�>�)���OȘl�#cK�B[u�Zi�<��|�EO+U�ȱ�V�r{��� Yq�+6��e[��C�o;gP��<�h��<�����/�xo��V|�*���a��uLCw�hw\4�s�8 �[�S;;��!fXm�ͬ�<�gf=��/F53�Gi	/��|�{��pAr��ພO9���-R���V�rT����v�o�kʹ�x.�|98��V�F|r�����k���*�JYEh�ݮ��Ns�Ͼ�����$�F2��`��}����׊cj�/�S�M��/e\���+e�c�B�V��}*���؇�5�u̙���W�省q�g����F��K���jw"���d*��h談Ѣ��w���7��>�-��x��lT�0�w����c�҃J�9��Z�ƍL�Yht��6���ٰ'�L!:�Yr�[%h��5��b^�石TH��:�Z�aeqJ�z44-s@�z7'l�z���Z��P	�c�S�~:&#��k��|U(���1�/����ԫ�>��U�ϳ4��ř��!0Q�b�� F��C�:͒�>�W��{�������S�Tɪ�����z!��0��<U�������@ ��&���(v	�־�sL��C����U]��0Ӧ�@GR-M��*����31�X��h�ͥ���������έ~�ճyQPw�s n�̓�Ŧ��
��S��Z+�%��Ý���- _)�$�@%:�h������}�F?FȎ/w����Ԅ����zd5d�oeΖ�2+ېS�=�!��
E0nFm�>�Cgohr���+w�k���pK{�)J�/z��)���@�[�a��tWhs��Oe�ՙH6۽��ѧ��-Y���v��_#hCv��%+�H!z�Z��o��H�ԯ�K���#��́ u���#LVlRe�̽z���=�_�@���1}�x 7��#�4�O�c��"g�C�Xg�?x�L�a�����n�j��^�!+��W��H��mȌji���n�)GZ���!�^J���$^Yx`W��3�L4��Y�dh��t1���]-J�\㋱��mxo��n	��hA���-7Hv[kkfm�zO�0�s)S�Ia.�e��=m�����y�\S��H{9MKM*�s��s�u��� H�Nw��`��������h�E�vj�;q; 煂���F�s
�D&Y~J��9��m����'�S۵3{P�#�!9݌v$����������0-�=t��y�{H��PnP�3�V�Gf:(tM�f[���"ë惲�E��Δ�c��5����p|��S�p��"p�� �C�=�v*�X{��F�Yz9���O,Y��pN��a��s�qT7��� ����(��%LQy�pF*��z���9I��,3��4p�M�vƀV���J��32��f��h���̬�D���f_�dMr��p@��䣛��߾�Q�0N�	��àS�����F��O#�<*�ôSX϶/�G5^:މbbRY\f�1����X�Cep��3�����oPG��2�V����� k^�� ?+G֕N��!�iث��_�ƃ��9�6-a�U�_s���x�ϴu�4m:�nZ��AJnw`��~p���=o�B}�	�� �{���o7�UZ�!KS|e��䨷b�-B�z���fu��r�����C`v;��q�ئ��y�[�1�I^��e��1���'_bѻ��k����+��.>��h�[��Փ2�B�9ws�#G��k8���e��l�)N����s#���w��,Hf����ޜ,�T�Z�T�V�=�v6ER.����$䖡.0��fö��~|�;N�c����f�ͱFĳ�xUA,`�=�>����僔KI(�|�/|�S�9y>恙�P�+i���B�N�\D�n�{s�oABmb��0�ޙ#0ihC;w቟�`���k��f�T���MkZ�g�5��SL<+��/J�W�䆋ON�	�7�7f�}��xAĻk%V�l�BZa���L�=�M'��w+���0L���.$[���Yݡw�
��R�޽Pؘ�5ϝ��p��B���Y�0�ø�Q�Y#'��*�V�S���O/������'f�S��^vmQD�zNFc[��b~��v:V����6,c��1Mb� �n�������ՂI$J���2��,Y`q�G 
��+T<�:�ϵ��nB������%�ba�Ff'��'�h�[δĒ�z��V�#�)xy��&�(�ہ>`�N_j�]c\[K-���r��vmr5�Z��n=��1p�[�$'�H�$��@!��F;�I�n1�_!���U�-^&�0�-�=��)��d�Bצ��2Y�p�WLK1�������ڄJ�u�!Ɓ.�\��R!�\V�����s�a�(�@f㼡��7;'$�k��i��V��8�KV��]g�G��GF��r���iO�Ǚ]�dZǳ�[޻���^7.J��szE6�z9r�S�^�x���?}�D���H��.�=����W�pq�1��`��Z��<�/)�yi�1�2n��*��-�hOB�Ϟ�O�@�=3��L���Xb�9u�K�hx�a#<��dm��U�z�_�"��Ȧ�Kdl�!��1f��G�)��}�P�A���t�>��c�Y��X��C�����q��a�]^�Kq��~�[B��5�s�����N�?��ϡ������]u��/��p�/m����4:��߾�6>'$k֓��KJ�g�7C�te��;���}�;�j\K�N4��i�aC�\��}�뛺"p���;�_t=�k�Y(�oq�J{M�M,�/ϧV!�~Îe>K�;���Cv��yDⴝ䵔���#�ٛP>���tM	��7��:L��,݉�n���7@����yV�0 �Ig=�2�;�5g(���5��k���{eۚ^D0L8F�N�Ra1��_U}��}�#$�B Ē�!>�w��~���""b���S}w��3�����A��0��Βwޖ�7�+�t����j���+79�u>�B#��ETE���Q��.b�O�)Z���A�=������[�6F�9 Ph\v8.�Cbjv����o�.�m��`�����86�^�^�t˞�εe~x�1��Ku./k�P���-Tخ\5Y#2=}/@���j<�J�+\#x'x�R׶�ifUȈ�5�Y�9�ğ�u\��L��[+U�A���
,��~H9���d��yKΝd	��|�C!!��f�1���I�s�>��W�+b�����T%vǛ�������M;ѾVs_�����)�AL+��F-=��f�:�L�?O7%h���:x���ĭ��sɍ���N��-��И�-��[�8��I�&\uҝaǣ���k�B��Lw�o��W��{ɫ>6�$Y?xx
�\jG��׷=��D�Jm���T��㔲�h�����W���'��Z�ȃ�w�耮>`��3��z~����jJ���x���9�#,`\��X�.���\��;}<)��]��$w{F���������E�Q�u%����g����?z���g�磯&{��,��L13�yuvq�S��+#��nA�h�G���:��M ��Xϟ*[s�hMV�T��|������D�$1�@c	x3 =���]��!7|���2�"�j9����F	m��W����a�rv7ᯠ t�dl���`�Z���_n���2+*zp��˹�IދӐc��C9��;�:����_��WK���ȗ�;���S���� �����5͎õ��^�׷����!����@%Kk�>��H�mN��V/o���5��90�C.�]"�蛎F��a�6@,ٗ�O���;�<3��,������������7���B�k��]�`8�!���j,�X����n�SCVd ��)��B���K* Χ�ײ�\�wM�cͩ!�aȵ>/�F���o�[D��Hٵ*�`��pM�LZ���A{e�����]
ſYbh�r�S�%�����S\8�{� ��O`<�	�iqZ�+�(�������;SnM�d�*�j�P�r����vm��C�F<�P��݁)U�"��˼��Z�9`��S-�Tȹ]��.��ৼ�#5���®H��ʺ�<ٛ���a6+�.Z&<���E�������It��U)���
~Y�aT:g���)���)j�C�Py�%F��vU-��et*�4�{ �c��^�ADҽ���=[��"jܵF��IR�c����W4�i�g,����t�W}w]�-z��ciCq�f�\�&7�N{���vu#�:M�a�)î���r8���u]�HhlН	�a~q�L|w}��|����HH ��bB��HI'�>}���}�~��7�x�o�M?����.��'�&��@ML���J\w�))��R~c=�!�*�Tf�	��IF���X�î�+�+wy8�Ѯuu~��'��#;�P8�o�?�v#0ʁ���m��6���8��.ۆ-=5�i$�k+�C�"|BK㽂�:�Lgmj�U�DR�r�,���m��%0ҩ��<�}�Ӟ�L���f�v�wax<�~�q9mc�:� u�
��յM+ �P`!qY�b�w�Q��}��O��lS8'˅A�����T��x���d��{�.�
c�^=X���Fƽ'�d�֮��O�Ƕ߬��55���F�9�����r�Y��#t��l%��k2��Ys��G���i�2{�`Y�����A�ּN�M�V&F@zuUs��x%��r��b��Վ�:�\@/��@��ZD��������iۧq��J%fSv���Ёk�h7b�àf��\�� [
���	B�:��=e7B|k�yw3ӳZ�u<p�����f]�$6�Fj�������~W&Lz̓j[^\Ǭ!E���k[���BߏoŘ�������>��G�LGxM��(��v򶐁Dle`�
�s:��>��Os���oγt}�L���������g\�J���m���ܙQ �郅�5�3e�X��O�WK�f���t������:-���=���`;��U�s�_����� Ą�`�7���UW9��[��H�����a��'�^lP~N����E�he�VI�zwy�{/B1�Ul^XQ�ŐA����@�-W�u湨e;oz��'Ԟ`��m�����NC�Y���:v�7T�c�Z��±�42Nk���-v뎉8��^P��R�Nl#�-�\���<(��u4j��2�!º�����Dv�|�@���@����*�Cb�a'"I:�w����M�c"�Mհ�=QyPu�Xό2Ji���O�o�wӢe��l�NǺfzΟ��y�^YW˙�	�]6��R	uj�l���o�o�D��Qx-z��ËT�U-r-t��0��R�v�b�u�.�c�h���㯘R��0���d7@攜Xnwt�stC��Pb�l;:;I���GA��B���Zc��`�7Z�I��̪�U]�=�dOn�?E ��hda0�	<4k�����0&�T�j؟F���<jw�B�O�jX��[a�Qp|��[�w��tx���Am�y6�)=t�ź18�#CK�^�b]>������r��_�Z��3W5��-%g<��4�'�A{�V���"qf�W������b�8M���c����n� u�*��t�ntս��l�AZn	*�ٻ��θܐ��s,�0��$�_,��b����`�օ%",c�]�
o}|�~z��$�2I����I )$ )$���~��_w������c?�:%�^�:< W�sImAh�Ϳ���倶tj��U<�;�Z�;��W������4\Q��5%�ܢW�	���_0�>y��_
��EY������(Rn�>���hs�]荃�\��(_ˋK=ɉ�,�sc���1Uz���X/D�6�V�!�.7�j�(0���J����D�����&�l]3����ǁor�lb4FS��P����&��ۻ2�ì9Σ��d_����q��-m���^��� o�~�a9��5}�N��:�L��C?��*��J`�ħ�*ޞ��=�:Y�j_��.4v4����{�����r����}^	�O����W��:lg�wQ1x���2/ok^v��)6��zl���"���..�V\0��[���cϝQbY� |�8��s�q �qƫ
�_²���}�Z����˸��/�]\�j��\�Y�ZD1�g��Φ�D�g1.�.�Y$k��8��4]��f?<AN��c�p���5Ct�Y���A������މ��APZ8]ڛ.�m��h4�Pu1ַ�]+�3[!�]yۣ$�>ƺ0h��O�U�t9�Os:��/-6�<٠ml�T�E��`�@˩E���i�n'nBέ��ţs#U�a�M����7	�a/iŐ>0Â{:���ts�R�Ǔ���ۄ����2ou�k��;�D�1�8Hf�Kk��_j��3�,�9b֌ހ�����j�\8`�V�6�O3���������vE������/�Rl�.�'Q�{h,�·����X0�lt��-^���d��HΟv�4��hP��͖�u_�p|����k �@�z�ɵ8EĸP� �[�&�e�CP�@֫�1��tu���4����yV�
�}7]�o ;-�
�V������=�\�s����^�;እK�f�Q��瓥�r�JV�n'�Aŉ�V ��q�oYZ������tZ2�� ��_[��o�f�x�ٵ����2n�6���IA+v�U�����Xv8�E��Q�f룻
ܝ��A�(�΄5f�ӣJ�9��|#��8��of�\5Ӑ�)�9*�2�2�v_,��+xQ`�O��3�=��6�k���J������mWx�n�ʆTt��L9�t����R�*�����&qΕ��a�;�據:q��=W����9˘|������������T0N��D�Pcq1KHg���墻Nҗej�2��Z2�4p;���Y|K@�������6_/qЙsn���gO��8������l����Rѓ��;���V�������G��i��ח�Vj�в��{_;7��P�w�3@/���Ό�X%#�J��X
���;^�9&ӌۧD��Ś�2�s\�;�%���I���1�:�T�f��b
��˓ct�*j�����ڬ���vX9J��E5�.�0��f��� ��l!�4��M�1X��j����㹃�H�J��F�G��iVg9o�ڥW��C��p�(ͭ����,,j5�&����w��|T%fC7r��Ecj���ם��O1�����¯Egmp.��;dLD�0)і�k�jf[��۴��%��\b䧆��a��o�@�r ��V�AR�+W��)�:�y䮘� n\�o+xQkj���oJ'g<��vڬTo.�`����;�|����{�4w6��M�U�3V�V\�l��*��Mv!+��X�-[�����Qtγ��`�B�������
��J�f��������+��Y�Qd�w�z���� yȮK��Z��<MN"�:uyW����/�si�8�����%;�.�v�TN�����fu��z�VS��of�F`� {Ƕ�:��f˩��5�3A9�FSΧ�Ʊ����:�fZ)1�"E6�wb=����l�N�75<qv���i�MZ�i<��b��D� ��s��[FT�Z
(��җ�MX��6კW-L���7-Fљ;<�<�s�0DX�c�()ݱ�)`;Ks"��i��1��%Q2������̤Ub|-Qvl�|����^�r��Z1Z���Q�h����UX4��m�YR�k(����Y������J��	[F6��V-�b��&7���(���l���֊EQ�V(Z4��;6|�&�O��Ī=���ꪈ,���ڧ�U�ּ�����+.!Mh������ۗPTUEF*��TJ7c��ADDN5
<J�kUk6�ZR��b�b��\���QPmhҋU�H�֪�j���x�5�UX�DT������`�����EA*������Λ1X�(3m���Q��3mN%�ډ�V1��ܶ��JŊ!�Q�j4�Y��EETg-Dۂ�J��j��0�L��U���X��-^�x��M��J�u�Z��U�%bjqȈ�;k����g-d�s\�Tb&Z�D�iJZ}s6�T>>f����/s�X�Z��	p�m�,*Ϯfl�-\owb;v�Fr���r[L@ll�4��<ͅo���<�c*�G7/� '�HB1$�b@# A|��0���\�u�ߡ��K���<��d�y�^L:b���Jc�����XZ���'��R��F+���9#LaL]�)�Ce���-f4��0�>ӆ�8�Jy�]�f�7�"�&_��8�,}�*x�>��6� J�&�m�I�?�{8ػ�Jj���'n�X�;xOW/��qh�,$-ji֠]�o3���]{�Ǽ���˿Ї�W�E~2��_p*箦g~w���&�X�#O~��t'����;/ʼ�=�����w�b����B��p����-C^-�bʺ�sPL渰Lc[��};�{s�h�k�Ժ��~m�2z���|C�p�)�:�%�>��X{n�S������Y�f���S��wK(��,�)D�6��
;���uŚ���~BLɿ-'P�̈����yZ��;@��a�y��/*vC�j�GN��P����ej��j��Ï�@�{�*S�c�6632d8�<9�C+��)<˩v4��ޣ�Oa�_x��	����Q���Ǝz�'B��A�O�q����p��r��1����<�v�W3'[�L��]2�ލEvl�	�J+|!�FS<����p��R�����a7�|�&�]ҧ/^r�>}s;.4#X��e=���랋�Z��ȵ��CY�S1�뜣 �c�������}_U~P� 1� Ē "I )!�w�\�-�Z���h��PM�H�����
���&��%��6mw��#��~[�G�$;\w�q_z�Y���ĉ�P�Ob����d�骭\��JӌA�6� �X��Q�uG��MշkN@�,9�&���=vC#��5�� �
�)�s���VT���`?1�~�FT8��M�h��<�A>�n��0��}s��?4L8����U[l��j���dn��i3XYt�LТ�A���%���C��pt�rh�d<�E�RS�1�͕r"�21ɱ�V��!�e1��[�'�y��Bl�I��m��������=��[�V�T��d�g�j�_A�/5ڄ&�R��w�+����8��H.q�<Wڇ�D� m�w�we�߶��
0u�v��o��j]��[_jU-C� l(������g��Gk��	�a?_�n2��LU�*��r�Jh0��������Ac�j��SƫZ��v5�h�[��uȎ�$d��w����0����2�N�6m}�G/���6zC�S^�-%�r�;霛�i�
��Z�l��Sަ=(,}�q�Te]
7�	m;:'&p,A�2���3��tb[�iUU�Oι��cjT�P&�l� Mf��oC��,�5x�?��;nQ<�B��e�b�'M��An�ٽ����+(L�m��n��U3��f���x�iiL�PB�I$�#BF2Bb����uk���}���7���9�'c�@�a0��zB�/^�ls=ܬ`khw�+��~@*���F�m42n�W�U��DRH�&����?	�O�<3��2�ے��5h��!,\!��8�����bAn�rs��ASi�ћ�F[L�-�iq�Q��K���>u
�r���]3n�L��N��j��3i��Y$7	[F#��te��9��4�!����ǽ�~9����Oi��۩��]{X�F�5�2}*69R�G�\�Ә��"�fl�i��au*��6[_FE��FE��	����L��f�8��&�
Q,�,YT�eek}dr�De���kI潵���Ꮈ�s�ۃ)��#u�>?L�=?>�^ō�ZmG:O[ϥH;�u>aȭ��ٝF56	�y� �Q����f�$ٓ�Dv�c�]��?r}/i��N%�O��#}W��Qi���a��&��v?���j�B<x��}�y\�S��Bʍ�w�eȧ�U�R�����@EE�QI�s�P%�+^�O�n�4��a�%��x-3�>l�9� �e���Mp��W_B0����󆏞x�J��Byam��,&`��勔��2�Z��'Q�4�Z�:�Wz])��f7�v��3��wuL�#��B���جEG�J�n�ŚEd|��=�a�{o�S�<�|��7��?#$@# ���H�� )!����=F���d47��ŧՙ.ݜ�X���g�������mH��-�� 3�l���"��T��ub���Ҋg5NT���P%��/@��iOe,����Mª�[L��d�O�T���4L�$�&�'�}%��J84'��O\�gU��Ra��4'�[#�~���RT�=Uٶ�i��ü�h��B8�J���w�!|����A�yߐ�	���g��6�G��?���uV*��;q�"�8�9��!?�g���oeZK9���}~}�%��V�غ1=��s�3E�t#��K|P8�|�,=wʐ�P��59�CMo+�� �P.׮�
s#���Ni�'yȖ�B��m0Nt�h�B�5�O��ۆf�GR|�/N�a <=ƭ���ai �������!��q�t����ǻ<��[�A��m|A�~9���lBd��3�wlt�g�������PC*Ȗ�]�7����D�ݰU_>��^RrJJ(�͡���|����7,Tu���0�bR��:e�(�1J�C�Rw��Mݜ�X��aK�w٫��`�G$J��|���1�'f�ݧٔ%�[�MN��Y�%-�bU��hs�ϝ1Z�Ll��ǯK�hp�;��Qn�j�Wv�rӘ���9����)����څ�\����qJ��P{�������ߟ;�n=��]?	 ���@�I��B@ �ؕ����\^��l_`3A�C+�.r	҉�V��C�e��;�������?{��S�OM����W��s����%7������G�܅���y�,O�� Z.�wѯiYy囹9!H�(p����Gb9iG�u,��2���F6���>���4�}CC��|y�6�_��EAL3&�j�k�1YJ�?C�觊e��G����v6��������Ң��o4��VN�Fa�n�y/6L���I�3	�r�29����[gm��0������5�n�[�e�w��Ǌy�>.�:Z���;!�b���+� 냔�����]�Zk��l	��Y�Z6��A�	�������_��h����_������ޕo��#h8NS�����'z^�w��f	Wh�i-u�8W���Pd��v���	a|��k~z�"��e�[��/$�:Րd��4����	����&����3��"x�uP]��>�QW���{yDd�@|d��4�ƀ�p�1��1�`?�|}�����4%��ΐ���~}�����6*:bKف>C�B�^�:�Q��f�;Na�Aں�c��a��n�T����y-�}�:�u˶�v������Ub��N��ڍ��l�N~�	h��c�\^��WC��A,�y��x0'W����QJ"�^��ϫ���T�1$#"�A��XI�IH � �!�G�y�f{�<��{>��^�.����{o�ݶi��q\τ��i*��m>Da2�.K�,�-�>s�w�K>�Ј��P"aq�W�~*85).[ci��a�>�P\��Cd�Y��Fh�Ɓ.��y�PB���ً�j$��Z]��]���i����0e����,d�6�9��i��מ�-ү��n�r��0�������nX�j�p��9��i�|�S�P��oR㚴�ZK K�����|�.*�6 �r�mk�D��N�^r�i�X�CL��.a�^�q&��Z-�P���Cq�)�f��s����q�q>֝2��ܥ���'��Rp^η������r���8N٨����D����X��$&g=�T����Y�Ts�aD��-ª)�s@�ⱺ���0l�_���P�Mt���3)��f��y�|��w��«v�>)�4u�\���y#f���3��z��>Q�ח4�?�ˇ{�������vA���J�R�l������coH���K�?E�Y��u�(VtT'nrt�k�r�a:F�㝰�i�i1=�����m�UG��P�4z����K���u:y�o���c��Wj�Wh�ﳱ}�«�<Y��������N�'���~����	u�4Ԗ>�T��{rr�j;��0���z����ݷ�%��>��Wu�+z�苊�yk��V䛄�L{Q���n�Y��f�k���0�1 �HA�@�,F�d�z�ϛ�����٘<)O�<����/"?{Ȫ���	tpz�P�{Om����!�P�+���~^~�ν?�1�)Õ�iKQ��c{��ĪX㍅
}�����TS�v6�c�9n=sn�'ۓΰ��kfZb�o
h0�	�6FlЦ�Q������>�>�oL��h����L�Vm�J��[�;�ϋ��C�?A,4�	����|e��=��9���u��3�o^��6+`��vӹUv9E��^IT:5�±����<��w
a|f��G��05��f6��,
�4�Tp��\���f��z��5�s�2q���0O�{ߕ�Ԇϝ֎߻%�����ש�:>��%:��-3�3�;k_��i�X��:6�`� s�kK�G����y�2w�Z���s	�J����qM��Ht�0�]5��0�5T�2�d�R]�	K�.)0��ݪ�}"��b����k`A����3�ʚ����}�B/ܡ ��u�䆆����+QZ����[�y|b|W�֘z��
7Q��K�f���j��B�K&�eSW��sl�AF�r�Ȉ׾X�X9Z��UQdu�\�eH�y�h�����s[��b��#��XjK��NN�'QY�rK�jUwN�U����ଢ଼�f�f��﹞`�"���4����}������|�)1.%}ﾹs��������`	��H�I� , bI3 ����y�+Bk��_�@(��^E5�
C*���"i; �hCp��g"tRu�u�a�ĭ�Kd���o�#_���/k�dSm3x��
��z���G���B��2m��#���i�u��+b�*�=�5��j%�d8��K�^�ʶ�M�K���]�aJi���O�kE:�³�\��ֵ Z|> +���9�eE'��@���#�:U�0��/X�-͈Q���u.�j��*��Cb�=�!\h���&�0��H����X�j�s�#�d��tIx ��m�6A�QK�d||���W�dS�z0�g�)P���<ɷ������e�ώ�CbQm�lk�W�̴S���d�I
C{C�~a^�^�%��S�?Fq�z�L2�k:~�:������3]a�s�W�/f΍�`W�Y�9� ��]ˤ��\n�zO=<ht�d��c����|�y􈹵�ŤgɆ5�����U�\^�?��$�H�p֧�CG��*j�+2�ll�;z�9���;U���D;hzq/�����+��Гl��,Yơz_,\֘�,�.m��k���VP9B]��"Z��O1�X۫��Si�E�c�"p�ys��	���_Mz��7������
�v���K�%p��:j�O�4q�N���@V���m��ܬ�pr�i����|���^�^|�}���C�0�X�db
��H�@Y�xx�4�3+KY�k�!���f���>�ތ'i�=�3�S�P��F[L����1��b�6s�9��r�@t���7�[F�]�͘���G@���;&}�ʪ�+r�[��K��ثVۭZ�7��.�����s��S�\ǿ(�c�j����D
�z��a��Х�x$��V_)��ݲ����ފ$漒���h����M��r2����)��R���D��=�Uz�z%��5���3.�5NH���cKS?�ۗ�GT;)�.<%��Ci�eF�zۮ��}7����ET���	x��צ.x����?`K6�v ���V�q�,(fò�h��i��O�����G�\���ng�(}�W�b�csTl��n�)���^I`�o>W{Clr��z��L��������.��!{VK�ЗA��d�=f4�'�ߦJu�?M�.t(o0�Tn�n�a�m�9]S��:,�/_e��g�q��	�P��ǔ�/	���S	�ީM��9�\�]��(F�i�*��V�:nr�į%���\�&-u��M���z��r��1:�=��;:p5��<.��f���8��w��~�"��fk̊u�^	��J}�6�X�V_�V��!i��_���^�x?<^:�������;��ܑ��u^��7kd�k��ej�16+�\�v0o W�^q.O�,�8S� c�d��]�f����5���������@a0�
� � d`��;����>�{��Ѳupo�JJ��hhX��pq�l}5&XC�:%�������AR��P��ݴ��]J��0�zy=Q��/�O>�Qj�"�CE W���y���^O[��� }M�3[�l�vB���t���	<�v�1pmG3����b���v�C�n�A��ȡ��mVݨ��#`�టz��^4ŏu*-�c5�`���|}�KPsb]�WH�t[uF�^���<I���E�8��=��GE047-F�v�;C�����j������&��R���W%pLU@'$p�_%�l��g��+'�SQ�4b�.�Y<L:�^�0�n�0i
�u~�:s��������d(8��Y�gOC�֯��v~"5�|Ê�M~���Ίk�bы��4�DTN��d�v�r���g��ٷ,cڪ\W�����\0<�g��Ox�����ձ�)�2S(���ꦶ�r�&��ƼUЬ{��i�Yr\�l"E�X�X���m�[“��Snٱw��� G���P4��Ul��ojThW{gV�C�������!��.��M<���M4}��曖��@�f�@m���;R�cGfAf4�^nWK����p[<���x#_�X�yeI��۬۷R��p�77���'��S3���v-�G)�����WllǧBu6ն�8m��YoK�[I��oQ�c8%c�ͦ���̚�!N�]��'S���&{�w��VF���n�ʺ�P���]�`�͚n�4���f���0D�B���D8�N��ӂ�d�:kr�*��,s
��5��(�(�X�Ujg��Vd��؎i&�E��>��@nR��Q�lϳE*,�+��c���[�۽���~�&�X��{�r˼7,V:�7i�&-�Y����(�`����z�Ea2̇t]�[u�H��>ݻúNk�%���:��L5��I���"x�\Z�=8�'J�qV�V�f3����D��5V��n����k&���%�	k-sX3�j�1#�"yS��Wj���c����$ҩ,֞iR��Y]����.I�)ڭ�vU�j,.�\�DF��j��1o�'A�n5}�Fq��4��;Mv#A�
��T�tu}��އ5H)��ӷ.Ckw��l�eΥ+9.��rq��6X�QՔ�\�.z�#���x�]�T��8;]mZ6��L28�|p�z�������X�%RT�Yz�iުZ�`8�%�+��@��5��M5c/�<��չc+�dz{��ik�j�@h^�:��/)Ǐ̼�4�1H�^�2c��|�&�:}�Ծ�2_=܈R�(_u�-��`b���ps$^���D��h���v��Ai�S�����:n���])C
l�D�����9��j��K�ɖ;��_v^уh9�C�6J��%t�x��XƉQF�e��t�EMk������}gC%MV��f�u�#��N%cu��Y�u���2����`�|7y^U�{7n�=���%�Tw�1�P;������we�^C�Q{�2*�7C/�	��xd"�n���}R�J_uؘ��E�saf7�0:F�M��Ԍ:رJ_'�Ε|+����he,C��:��}�f�D/�N\�_n�*2�
�4�NU�ɝ,y����)Nb�'vN�X�g<�fEza�m�p�G��c�����%��7v�B�u�r�%�Qo
�7���>*��mLc
f�2�f8n��.�БQ��a��l.�����%]�-�tW5��à^�z'%/I��`]���ެ�֝5H\7����c̬ѧ���Y`�_rj`���vu����a�c���̊�\z��9�&���3~'&��Z��fd\�]�K���tN�59��P��J�B���};�^��f�+�"�n������ՙ�+S��j�3�!�4����&�zr�3��ͳ��dғ�s�>xYݕ�|d8c�4�ޫ���*�b&*�B�)rw�ڮ��{E�W^)#��Cw5=�ĺF6���VVл�=�n�]�4l��ˤ���m7[�3�zuಥ��Z,M���(���U)m��EjU�*Q�LDYiW�1��Uv��������'������JQcr��֬�r����.Av�%>�8#Z��W���X��g.�ڪ*�\j��gg����ƋiDxљ�X�ښ�F?�J��e6�)m+am�����h6��vy<���U�o��$�*�+F��mm�"e�.�� �R�1�O0��%�8d�,�>NN͵;eG<��
m.%UY3r�*V������b%J�n����5TAƬ1�U2��;�25�j�J(�Du�*�ص�8������<۬����0�׶���o)�J&R����Q��Y���;J�h��˄U�\)iC�`%�E�*AĖ�n`7�U�1q���mnS<i��8��"��J�R�TS˙j�e;���9j��J",x�ZQ�ͦ�R�,�����K��R�l�����m�����\
Օ��Cw��k\j۶��(�/�c�x�e�v�Ɠ�u�-�4������u	���5R};`ݩ��Ϋp+ɋ�7���0v����N$3���u��B����٪�6t�2���E"0�a$#�1��B}y�����79;>_.{B�9O�Q� i��.�|ǁ`]���?��U2.qt�l����V�p�Y���*��#�;�y�ƾ�N�Ƈ��юC]������w��u���!Q�;��;�B6֊��顓�gv:(\`����E4�K�5<!7c��=�ɠa�,QdS�0�kU����,�Ƽ|�3�8+9�d�gC�����vX����w�Q������+RO�Y�l�|0�J���W��*4�Qϧ��z����o�H��i��GP��6=Z����e��7_�b���B>�9��� }�OI�{��n���ܟo�V�(zYz�*%G��(��͜K�&_z��ط�qAÌ��#[uF���c�ܵ)��3��T�VE�&� [��u��,�si8a��ϐ�<&P�1�q�o���F66�zF��=�i�9w�nMFޮ�]��-|Ɨ�b}�.�z�aQ��9a@C�$(��͎w�U�|���'v�:�x����m���o�%��x��/=�;�O���><����H��.�BCJ�-,���kVߓ��m�B1�zʻ�5�o�~�F<7ilƊk�*����h�c
���p(��Ε�V�1���b8�G��C�������4(��N�h�y\�[Eʒ ��'1�
Wֱ��sղ��S�U��
�p���ڋ���]=�>`��U~�a$RF $a�$Rd`
B����>��Ͽ�����>?�U�i㆙���-��
E'�*]��'3���ip����	�WJx����t&�r��
��>���`��D>%	�q��9mc������OT�q�s&G��.��[��=�k�e
z��yU\�kTP�o^�d�EqT���S�����~���<(-�}�������d��Mf(���3F،w��2���?��k�KRxf�ew�E=*k����u����w�1�`����G��`o�!H�K!��~�UdP�q�)Sҟ+a�8�#�ߖȦ�)Vk�`Y>��1��<�BZ9A6��(6k�V�<hm�Ն��ჯ�Tu���F�_I���8�Nx�� 5��l5����:��6��3�����k2�wz��(��ӕ��(A�:��n�y�rzf)����P0$��&X����l2��U���e�f���VZW���	���i��"�=�t=��O�\�NĻ)��U$�:`0���K��5�lwp��923�xhOĊ�<�ؤSWa�/G.SJr�_U��񢚾�S��F���r������+o����Ò���K/�'���h����B6���
�;ޏ��q��(�A�z؆���Okt*R��6 ��tu�ĸ��-�}��vS��o��9x����\r����N5V^]s���}�����{��?�H F$#,X 1 �,$��$�����ڇ���{�����t6;1w�%���(��W�S֙}�i���H6�V4#B��2��m��&W1/�Ǟ��z���j��8#�cxK_?���I�kU�P��jc%�oc��!k�N���-t��4ު׮1a��7�C��4��p��[�]F#���cn�?h�b��G����kshu�����_���S�H�?� 7��6n��hV�E�=�Z�P�Q���!�Jnd�
[s}>�d�{�u��S�*�������1= �EV;���6]��~LLGu�s�O�;=�����H��[wa&,����0�`-�V���q�и�yZm�J �d������x��6d]�IOޗ�qmqP3/�5�~y�w��Bbx\��Cas	�vqKv(��� =�u� G�P���Q��dg�����{gBҮn��>r}���Y]:�j)>�+(V�5�)�-�xyP캃ظ�=G��u������:U5�x3Wݶf�h��C���tX�(-3�O(�eCNh*�\]Ƭ�a[���c�	@�Zս:�FU	����[�V������W.&��,%P�"�Q��m	:�^	LLi�3{�v_t"�W>G�},I�l�(�����+ٶi�.}cBX�Z�	����]M��Oo�"MN}5�k��rCR�^ާ[�t���u���
� +�$�`AUb���Q� 8ֺ1RCPxV���-�5�N2j���n�)�S�M��|�σo%��Ee)|�pF�.��OF`��8�'�9){.5��[�0z�`ي;M��RÛ�Q�q�M�"����~������o����;��}�|�m�� -0�9�������y&	�LS��Փ�O�yW�U����L�6ƿM��O�Ƀ��I66`1t7a�
�6cLm�+�St�R�u��"��Z2��I��#%����A��kM_��~N�Hq,���/4�%ftNM_b�g�u[	W^��Ĭ]���.;�T'�j;��T�5|�E���z~Lheq���;�A�}�w���Й��V*)����ޢN��I��1��E��s�:g�a�]����ʮ��WuKj65 x���1�?�}󆾠.i�u~7<��&o^�:���gǓU%�B�`��=����	8{�3�$o��	�S�w����z'M��H�+h�M3�Ŷy��F��>�~Mׯup�n4_S@����^����g=�O���<����:��y��i��F�p�o� ���$�k9�;N�F&�h��o���<K�{;��	�Q$��8z;�W�zz��f>���y�v����X����bcPނ���O�0et$��h���-�W�6�C}���7Jc��7��]"�+6We;�˝�Ϗq�瞾WF���1���Ă�1��d$��g�u�F�
d�9��]yIw��� �K�E���g����Ü*]�cY��_'n��Y����vk�>Ĩ=]z��C���������:�T���i�������w�ѣ�n�*2�T����F��k19�J�\����	����۝20S^�)������;<em���o$U�O sӾ5��¹�IU��C[ L[O��t�n�x��Um}�Y9�3��u��omy+�����w)��t;o:g{7ޯ�^��!�T	]�E��_zP�:��'vd��f[[El���%���io�4���l6闧k�r�嘛��.}�-6:�-]�Ɵ���V�JxE'{�zm���J���MI�?`�4�G'���Po�P��w�~PF	h�t6ZݓtK�67�T����B��^��R�������5G7P	J��*�~q=`��ѷ��_]��6.W�#�ф�4�O���W7�a9B+Ī���	tqԈοք��n���u��y�!��%�=_��>�B�� m�{�gss�7bSY9>�{�~�L����魯���B�˲���ME��um�8%��C�o��kY�w<�LnV8q�M�d����̂�:�m��f�ujΌH� �l���S�WW�&l�&#(_Fb ��t ����(.�1�E$Gj�6Vu
��G�0�#Ny��6�x��=��y����PF20I��$R�~�ǻ�s�{� �04y��4���g��5z^[�@�ު{�R��êiO��n�weLҥ�n���6,ź��%�ŮxKW��򠯏�����?�v>to�O��'wg*jKsh�"����; > :����4.83�)zΰ~~"~ks�W�A/<�aR�.���b�Z$�T2$��%C�uny`^v
"~��Ο��p|�CW���Ǖ�=��a��׌k�a���#2�f*s�pKW-�n��-���,H*_�/:�坮�fP��k�c�4���zǋ�T�O�(��aN\yk��q-��$<�	�J�!�G.�,g�0Q~CҞ�V	z���S�&�&�a�yy��#!�4����&��usl:F%5��Y<Sr�nU.՚e����ɺZ��Gȏ��vۂ��OU�K;��A�Q���=���՜�_60�];�ϲ/P�z�{����³j Zޯ]`�iQn\CQa��)�9��(79t>c�k�Ы���\�TO&˴i�ؤ�͂�T@j��B2�:V�Y�J,d�㐪[y�9��=�_~�/C�\���ui��O:��FKi02��.��`a�_�{.��ϕr���6AU̦]R�g�+(�Im�r�ʍ����"������=X<m�s�����Z�kO*�A��:aeL�'i�\L���I��]�\��gD�6��̴��b�'[it���>�/n�#�? ~D��@��`� �7(�J�6*�a�lw8�?J����~�P���l5��"-�K�m��[�̞�^����72t�x�����:,�3��$v`"��u�w
�K�Z��~W"�H��ע�[9�?u:��jq��4H!�r6�D�u����6��QѣuHz�0"��f�Y������`Q%���A��f���`�;��i�6��ms��t!�C�K\R2�K-�qn�;n��\:u�j}Ϥ������ ~}�QN_yC9gN���ް��A���B�]Ax�E�/�О�l��w��	�j��8#�`,���u�P��Ū\n(��[L���k��OSN�m+�e�e��-�Z��5:��1a�� �@ U�9��c��m.:�w��+Z&2��]VG�ϻU�b���qx�w�2Z��OW��|p@o����GEܡ�ŗ��q�q�^}���=!����D`��ln�E��������}��e�-�@�P�`.%>�ϳ�������J7�Pz�|��'�� p�v{�c�ۘ�������x'��_R�����*|���koGsB�t�6�h�R�4�m<�,t:����֫�7�Y�O)su��81�q)rj���%��-)j:V_e���.���%�LȟFڻ�ޓu:����h:�+�fB�Ok����}�a|P__D��̧�s� �� �b��,"@�j3�L�Р����;m�ሪ!hByT,^� �T��v}G3�~9������6"pxZ����ʇ.[Q,�s�.+e͞'�C�4�].�u�8��^A�{���UN�)�Yò ��4T�wl�{�2��QI����Ͱ����MN���@� z���:m���w��]/�i9說ż�T7�!�Ze�x��J:�-q�m*�qg��nH�r7̚D��U����DM*��-b��<�TX�q>|���b9~�]��EY�wr٪�%�y�]I��\�{ƥ/�/HC�`���bg����0֮v�1OI�m��RӐU����Nu��d�Mr���s`��Ȟ~n�	�Nx,��4�a�e��1P���6� )���4��M��-}�XmA,K��,H:3R�e�B�L{��cg�]�T�!�f�i57ڇEX� 'j���M���R�ڭac���1�`�ޟ���� �e���w��������ᴦ��Tyng+�1R��͸�]<Ҏ�L/'5�__�g������s<�<B[��jo-l�RdM�����t����j��,e9,Ps�%E�qJ^f��)�ǙosyL}���h∏+zJ:�t��W�UKH'dJv���0���(�sk�z��N>;P浩�u�b�9y]mi��Ko&1C��Y�zR+&T���әdE�C���n.��y�?1���@�������[�T�M 0-�1��z��]K��OQoQ'U��%&2(Q��BMSkQ1l�۱�ŧ ����gsFς`�aw�P��@龧���޴p��Ά��ę�:1�)�%�k�,�xtN�	S����G�:W�Q&<<ă^yO��,+=;>�5͏j��М�衖2U����ͮy�(����Ot������������b%�Fqi�NG#XF\�
ͤ'#�g��!l�q~{��pm%�P�*��^Y��zb1�32<�0�1S�w16;����$¥����'�{.�����o�듦>��r�m�mU/�^v�$j��6�	����Ǟ����> "��A~�5U%7R�T��3���V��]
Ǳ�EPYr\��X��քWg*�VM� XӅ�a��!@*E����Smܡ����3)�~z��} ��r�� ��~���!re�5�˗sl��|M�E
g:�����Z��y��abze2�T���e
謼����S���K}F)�|n�QQy0*�<�.l>uA�Zr�0Wd1� ��at0-��#���Ƚ�G�޾�[�B��5n>ƹ��Ůq[���쩗̋�R�h��y�H`�|D��"�������^oG6� |���̭��#h�`"�.՚U]� YS��ڷ]����(��_;OU�ҷZ�>�����P��y����7����xq��2D�O�h��bS����m�����m��
j~-��:hN���?��{q�P����w[�,��P|�L8�4���<瓑M��l�
ΊhNǈ�Ѵ����?WTQ�7�C(�E�ɧ�OsR�~h�l}��*Ԗ���"�U���D��b���{'��z�q�k��$	�t��Z[�I�x��ddڎ%��*�a���83�҇����ļ-.SK�Z�4D�`+�v�V��<q�Ɣ%��c)��O����������]���}�۾/۳:%�EA
y�K`�;��<1��ˍ7�[���H��{�B�탚�m�1vgL�=vk���G?w�������FΦ�~!g��6B��V[��M�A��u9՗��+Pi�#�&�ź�us����z�W�>X������Π�8���'w����)�l��uwb�{���Ω���]���@n�v�Ӵ���c����P ��'�s˜�`jʉ�*X��E����5��p��<�5��d�y�{2e�wxӴRRCm}舳>�P$ k���5�}�����R�m?��h��J��'H���������|���0�OM���N��Xg��$v!�m�*>���7�Eϣz���[���ŕ��ޗZ���,d;s����3n��u��,�N�g(V�qf��f�0�|R��*Pk���XE5@�*Qv
���& 6���)	��|�QpV�� ����`Vu}@�SV�bRø��u�8P
�θ&��W�y���gX��Cf��L}:��YX���Ƕܜ }�t��n��5j��Ɵe�ք<�!\�-o�����^�/M��)qسޱ�(ӦJ�/��.�Z�xN�km�XZ7NM{�K�عtWY4�@]�F�`,��8<��OS�M.�@�m:*ٯ9�\���*O��}�Ebyn$zȦ�W0Z�v'PC�w&�JuB�bm"nRu�ctL胃���>�a�0���6�ݛ����t�=�pM�*�K�r��Q]vT��s���ʲ$3v��C�vBV7+h��YSt����C�;���ٯ3�RS-�J�yk�>@<LGML����,fb�]n�G$���w:��XH���R/��]��j]ˑ�y#;����h�΢曧�R�������g6�:|ך1ސ�꾣�Ɗ��6�l������4D᳣W�^ڶ���\���S���$/N�q�CU��f��]qʍ6{"�=��_IV���p�9�Vj]7�Û���ҝ�ky,a����TR�������+����mq�豆��b�1 �wh��*�<��v���9����#���u�:���;��oj��#L��!���f����_d\M��)�O���#)��Ě�wϙ�Wqn��A_3qn�.�!��_H�$�©}�����/Y-��ٚҎZ��N&��@�ރ]���և[*�-������Ǫ,$u�ɆȒRk��ZtI�V�DwC�Qᝓ5�m� (�z�E)}�qU2݁*=��w[ቾR� �����%���;U�&��Z��
�A(q4��!ջ�6Eh�y�ޕM	����l��x+�u���e*+R�8�=v���<'������k�UtG<�E�Ru�s��J��xz�y��
�m�����(=��٥��1:9�ͨW]rD�Ͳ{ru�(Gn,F�>���.׹�%�鲦 {)bE㼮c�v>��}��ɸh��%�p��87+�y:�q9[��7���q��z�M��cm�oCɭ�n��a�3$�9Hw���ҏwmvs��T����v����'�{����WUK��(�x0U�so������W�fl��1.������o5.��;�[/.���c��^�<R=�F.hn��o���ۨ�͌�*�����8�,�GIR�Wͩ���c����LBw���N�Nnwe��3'q���[���1:��o�{s8����:�J�V���X�Z�h�qp�0��kJ|fr���lՕ�ܔ˳�v|�O'c�*VW���Uw,s�\����&V�P̗�Wւc)U�j��lVe1�Z"̞��g���`��aU+D���`ϙfZ��2�\±��mˮ��1�Q#�-�m�<�O'gIыX�7tƎ2�J��6�9�eJQ�}Z�-�-W�"�)̹��W�ɭE��L�>O����N%b���/Z[���U�V��Iu�n��ܹ�M��M���
��U��]V��R��%gmN�YEb�ī*�Z�UEF�w3ȶ�*#R�Vۙ��+�k�bDU*T�^��"AM�1Ԩ����TA�L�EQSm��QU^[Z����+���Թ��
�ʦ*)���"�,�.%�(�3Uĕ�U
�Ci`���aQF%�\�0��Z��ܔm(#F�m�n1C��j�e-U��8ܱ�EV"	YP�[JƸ�(�8Z�8��"������E\��k�A�_R�@"	$)������ua�:T�m�����ָ�������	��d���XwD���Ƌ�%������_�1��"�;��{�>�_���?/-��Dk�8���5�\����_�L2x��3'����s�+ť>p5�*���e" �vۀr���Mf(��A�m�����]`s��z.���W��TF�w�D1dt���[R�:�!t	�yoR��&�@ꆲv	^N�"��e���(˼H��'Zbo�Ü�����#��;�Y#'���h����B�����<��B6֘�|g2w[
݊<z�o��t�.��yň�(�gQ���E��u7���ʋq�\��K�ty��R�7�*���-�إA���:q�����{�ejV[�*('���@���(t1�ږi1в孂�u���y�qІCL��A~�>��4P!
��"r�T���	��bze�{3;kX�uk�]�����M5����>��PE<��A0�چ�>���� ���)\N�g4l��SbP��c����M�k�$d;��O�����Hk�W��y�}2���k���y��Ŋ����ϽK#ƧT��2���Y�����A~p�ʕ������3�����=F����>��4K�XA-�{�V]�V]�ө��=vfʕ�C�;�%/n
.�� Λul��ݦ3t�4M�I�;��T�=�nT��h��ua�v�WvD:�lwr�[���}�>gy���<y�|�Ϟ������b1$
֬�A����\����e��q����4��GD���ǀa��6w9=�I�R�NK쬨~~k[$����0;ntd{������mߌsxf��.(�	�����2����f^������3��l�����`�zY����^��} mq{�g��E��
k��ـY�������d��8�6W��8��F6��!F�Pb��C�mUA����;z�L�h��1c֝ii����z;�H1�J�k�bx�9�0k�������*�=��%rzu�d�NN��BN�.s�O�1��Y	��;8�O$�f[A��2����L	�j�����/�M����nm���J��Q�k�n���}I����+˦�H�YP\�N��p��w��E�����޾`M�0�qra[�k����^��PXz�3�;^YrՉ*�q{p�B�6v�b�o��J{�Y��Dn�0{�Ob���-G���8S�l�wL$�Ty!m��י�w(��%��
��z��)������e�2A��<�uI�钝D��# �|J��HJ��ׯ(M��i$��ɗ�[�)����x�YK@V�v��K����t�����q�}|�%��'�f�Բ|0��h��M�sή�����W/�7:7�T={��A�����sY��o0Ѽ�����2�x��u<�����u�ȃA;p&���!���,����b��?"X�����߫���貶�fn�.c��G���u����#M���r���n�����7K:jU�T�0���V��Ḫ��0�i���8�}����|Z����PM���Ǭz`&����N����Ѷ����*vxb�t�yV4ч�U�/��%��`^�"��Xk��ИHa,���N�"�͜���i��31���ό��B���Z��zy=j;�e�%���M<�]�wT���c`4n9Y&����z����ϰ��?:E2��-�N*�5�����7?OU.f���2F���}E�s�E6��4�p�Jǆ:X`���L{�Ֆ��3\P�d����1k^��l��+[MՀ�ȇ���SA
[]�ߔ?��@��3ʢ? ��p�3���Q�Z�b��d���M�k�sE�m�jʆ�������xO��R,��w�8��x�(�-17���\��,�j����=�������c�Y�ǾG��x�{�6�'�E��9¥�@��|3mW;�'�;v�sV�zaSә�ԙ��+�U��M�x厽���-"r���p����_L;AC,6�&�y��n;+�����n9���8(n�?g�\T�/��R�ڪy%AI<�k(K;xY#Dw�d�����x�n��h��Yy��iЮg~k^s���fQ��(!�:vEks������[�)����C�zd��&%KoO���U>C�������k6r;U%	���xK:�-R�4ȩ�boW]75�H��@Z�[h%R�f��i�l�z k��7D�]|<5�Z~D-:t�0�C)]~���.=��6�U�mN�O]��ߝ7h�IU9�Z0X�j�ԼM�|ۨ�oo���Uk`� +(5�J�}�c�?�P�K�m=���jdfvp��1�h��ʤ.=~n]66��(7#;�V�S�c:\�Ƈd���$���]�p2���G1�Aףv/�*�7v��igQ���X=Ҡa����t����U�k�5li!Cb������H��4����k��_��l�+�hN��<��׃+�����@��'���|3p���DF�5J�.p��%���^��n
�OaD��u#��Tc7�Ыȋ�D����JщV��9��Cb�P`�;�ޯ
�l��E���U-Ad�⣛�B4	%�F����z��ST�* ��	������/��b���8`�kz��|���ϯŸ��>�N��m	��Z

|�07���Mr���7�wlw��a���|e��8�=�C�C����:Ţ�u�[�Hm�T�<����{!�y�p:�;W�UyG�u�w5dܴi,y�3Ea*����՜�8 �¶-&�0ݬ�txs+�08��s]\����L�ݚ*a��As��F�wn+�Cla�Hsk��K��}�篷�ߞ�ϟ8~�#�c >�<�c���DW���S��1S�ǰ����+����Z�^��l�|��"7�~��J�=ƙ���/Q:�}Z���ջ_28�����хއ���f���,F��v��ꏙu���W�>�g�7��g�t"s�;l3w���>`���(`*m8s0�o�e�R�n��녢#�6..�.#ѯ�f%�u�\{D��wzL�D���T�amY2�Zm��fT,Ff��i�l�r�r��4c��#y�KBiڣ~3�GU�埿'���#wa�*m8�E���6�(�S���E��$��!�F`�~4����`qy̫��=�q���sjWOr����&��C�d��^6׊ʦ)\�V�Ӊ3d��Vn\�D�e��=?a��R�c���Eb܆܃"4�
8伧�<؞Q叾3yE᥯Nn|r��T��SIr�7������z0d�w�BWK�VA֣X[�N7�&V�����+9e[j&�%��^̭�3}��ϡ��	�>��O�=lh"7R���Ȩ��}�*�.��=CQp��]�Hky�m�l� ����4����[��乱B��/R��ûko9�"޹{��`��ý$���t��I��zMl��x�%�%�7DE��f]��'r=w�"ΩY���"±r�t�xKruw��Z�����t!��"��'<���v��{����� 1#��(Z��1V�����;���	x\��rM?2l���C9N5n@E����:[;bS��##R�m��^N�u1����8x�����i;�iyG��a�N�v���\u,��ܼ՗F���ӎC��-+��U!d�8,��X]%��$w7��ψ���U����QQ9�I��.�TF)�])P���i�`�Ѩ�,�SΩ��L�`(�40��\F���R��3�_9uWt�2h(-z��'�Ggd�'`$hcV�H}�UZ��1b�i� pN��t��8ٚ��Sg�<
�H�?��x��Z�ǿS�l;��ɱ���n>�F�(/�i&��յ�����[�C�b��mx%�?���9c\c�r�;τ��&�.��`YQS���i��	�j,Iǲ�P�t����%�y�'���g�@_��3��푲���͖�L.'%�x&Z���{f�T�b�>�������TB�sƜ��ߗ����R�)�8��u�S4.�{6�Bk]�e̵k�@�A����w��ۼ4�}r��?�HCR�wI���2��K��-:9x{�Ov�b����^ӳ���q8�0:z����j�:+���5�mڥu�+3��o�=�f�TW�u�Xeũ�4t�|$���瓱�L;ٜc���m��0^:�I;.��wZ]^l�ݜ惕}S+Mh��9�~1�F2�y�Ͽ~��>�\י��@��E���S	;ҵ�gB���f9\�Zr�M��+*��s�1���i�-h�eК`"�t�����)A}�&}���84�t(n렴է�ueCM�%Y�,��v�F��%���na�z푑c��ذ�,�G�P�4C>FΊ���O���T��5\ݦenu�]7��O7*�nI��:�t��(��-�f`�˨d�,�f�����lʬ���aʲ�&��o���D�^/˟�>�f�n�K���Y�&�ϣG�Y�ADkmD�z�Њ���VFVϐ�㪐�@1���)z��˞8j=%�:|Ly�	������n����<��Q�ؐ���/���vH�ƌ8�r�s�Vh�Y��Y0lp�7�k �=1�rP�jT��H�\����矐�s��6.��P�moT'�Z��`%����_^��Ҳ��70i5*�ꬳ�!��yA��聢9`�u���isu�GN����WPģ�����4�o3�N*�e�5�æ*�C���ZH;���{�!��0�}W4ɏJ�mɜ���m��`o�n��u�^O;�&<Wf�ۥB�b���bx�9[����ଐJ�Y��+ �����gH�a�'�6�����
Δ�������/ꗚ�f�]��o#�ʍY�gg,ʺ�L�[xʝ(;yܥg;X�j8r��d���gx���k��y�y�����*�7pT�M���S��Y�������C@?VC7��ё|fGEX{����bO�j��3�",˴�|v���-�_)���*��=.�ƾv}�J����1� �G�*,m�#v��`*�#��vj��ُȝ4y��Op����G�E��9¨DKlݮ<Հ���ڇѺSx({ށBj-dX��S�v���r�APC$Z^[6厩��;�鷉m�Jɘ�F�b�6�4%��Qp�"�"Fϭ)������P�f���uT�Y�ǩdi@�[�c���4Ԑ�{��M�hG���Ĺm�S���2�|�먡;�:��\N��~�ΩDc��jp߭����N���U�UZ�w1�6N"Eٶ&E;���CG�l�L���pk�v�V���-�h��,p��<��M��ˬa^*/&z�\Kca�:��r�-$�-{�gi�����$b�ܽ�"f��=��tU)��Ҏw�{X���E�-�	V���랒&� ,��Z%��E����]�4&iW'ǣ6_�~n�����|�k*���I���%�_�3uY!]�]:�DsbU��1��z�ʒ�g�T��a�ʓ����l4���>���ot�b�E�1�̴��.U�qR�ٮ�l���0ɚ���rv8�j�f�i
}�k�nj��
�7�9���������Ef��h����󻣂c��{"Y\)-��y$���4ˉ.��Pۅf��y��b��T���̍�]���
���>!%���R�����؏���aO��ݸ�|}EL���Ʌ:�#��������-5��]�h���U�ƄP�f�Y��h����e����cgQJ��ntD����}�Z��ц�dD�<�ޖ2k��a�*�%���cq�����	�� 4�t��{�A����3=#b���G��E�E^��{K�)�UR�x�؇y��\u���BE�O���c��Ō<x/<�T{�`�I^T���ȭ-�Ql�	u�{�%����9�ɻ<��Ō�2����vl�C��4��������8��p�͔�^��Yy�;z9�Ұ�6!���S�`pH�E���k�h�ɘm�3>�����k:ê8J�`��o�X�|�����P(7n�*�-��b-�(�h�߃L�����Y��<\��J��ҧ3Dgp}�L^]%�_�D��6+�=i����5ċ��/^K@�i���m�|b�j#�eJ�[�m�h��r��P� ,s

҃�[.�t�*�:I�J�Q:�rJ�Ձ�.�P	��)_<��la�jhEd쏙md��_VW/��vV�O�V�ts����9� �Y	ю
u�oOn��.e{�k�������)���+j�@�蓯x`�MB�K&���n�Q�='Ŗ=����
��fV6	q�N�YQy��f(�v��-g`vGD�{�):���6�`�o4�H*���(�دE^Cۡ�g��4���DE�&����k �����Bt�7VA Z�a#��O8�?I��ѣ�[	��h��հ�m�n:$"A���ݴѠ��Cz=�>a�8?���94��^΂'ͩG	��e���9�H܁�n�v?=��k��m���!s�*�<�s��/���#ӻe�ݰN�h�t�kE���)�<I���m�����w�~��l��U߈g��
�n��r��Q��7E*�]�)d+qQ����\��1���Mϵ�2ٱ����!G���X!LYfU/�w�����j�z.�����V�Ra���	��kk�5F��c��ͬg��%��@t����Yp���<׊M�j�	�Aei�̣����c�e���5Z��fu��~0�Ҕ��#XYB�;zDkj4"@��ݛ&�!�9���=��s�3�C���)*�O� �POa���N��.I�S��ǋ5����j\��"`�8�pe�8;+�������iY�Hʱ5S��bښt��0��إG�r����t4�a�112�w�:��XfI���;+%uI��v���(�.,T^�l�"�Y�_Oo��;���}�<���aV���}@ɢw(��u�)�E�W�$b.�&��I��H����Ԉ_ �Y�-����t]��\�;x�im!���ⶴ�oS�2�L}�6TԀ� ��݌���)��1v�a��0M��>t��ZgKV6����	�ha�>�Ylo�X�V�&���P�� >u�lV��)�	�:HT(rٟ��t��+�=��Cr3����;+�5����X���Ɲ��Z�,�x��9��u�##d�����T���\o����%Yލ?	��f�c�tǐv�H�ʾJ]�j;���pp���k޽�{����:�.Al���Ӄ:��xԩ��:�8���99��Y��7~���Q�2[][�e�sD tӲƁ�@y��mF������ĝǝف�Q��
�\tG�J�d]ބ�x~ i�k���6@.�"'���N]:Ŗf<V��K�%`�;�Z9|�Y])d;i�wYvO�_N@��3*��^�t�ܳ���K��* qT����&�=��2ء$����	�����ೞ�-�6���W���O��<����q0v������B�gl�
ep�J��Lh�M=���)�9�n�o�n��h,�t�ʏ��b�:D�.G!�)�X=�eC.W\ݿ�����%�vb�)oY��:���aUC.0_�#_�椠�Iaۇ7�g\�HD�����0��+.�QX2���љ�G�{V�(��zռ�ړf�twk^�K�����`A�Zb����,�t���{�=;�IO)j�Bm��V,�KU��V�Q�&�l���=鼵�e�Y�*�j�9�E�f@X2s�Kq.U/O[ͫ�)�G �vwf�V]�4�s����9�VL��ʼ�V�:���u�9$�4zv��'�\�-�Jk�[���η��](�T���)h�:Ճ���9�5�Vྕ��E�n�G_��{�xױ,�[��:g�F��3tⷷ�e�}���*�=w�gT�-ǩ�ڣ&*w�y�9kN�ف`{�vF���mؙ*6D+�s�T}��)#���,Z���W1��Zݽ�ah����NvMui�.��M�41͢#�F��K�|@8�5�%���f�(�e�qm��ޢ�Lc��L�䩉�i[O�s�[+�[e��U�. \X4ȺdT4<���MK\G>y���{,���)h��Enp��oB�T9��9�)�p޳g��`��i�{7�PRGC0��.���5WwT�ne��y؜��j|4�Ӎ�QVL�z䋶�v�w�����CgF<��7eI\�W+:mra���v���s6t��ۖ�ྋaI��.����z��F�J�Rk�m%]��v9���[c)d�\LBw���N�Nwod	b��8�۹�ب����w@�f�A��J~�q!E�q�EBiZt�����JMң$�]�,�D��
�Q+Fضzʯq��U3�O2�M\��,���������Җ�J�bkPY*�ep�U-i`���Q<jR�R�Q��[B�DfO'���ثևS24�®R��r�\h�5A�*��g��D���"�����N���N�~R�O�~i͘���*�"��,m�#~�X��X��r�
�J�R��RyK���ϓ���أ�P�R֋�b"&+Gs&*�Ucm̸T-���(�Ŋ1�l1�R�
"��qƬ�+]�՗iU���q�,F3(5���kr���E\m��Dk*֨Z�6�Dh�TJT�,������b7L���)�S<�4PR-J���H��D�5f�n�,�`�Kh�r�b�Z֔m��c��2���[\q0R��2;��cRĘ����hV���-t��lZ6�WX��wu�-���ڳn�U���m�
¸�B��̼j����<�^e0�X|j.Q�q�Z6��J����7nV����4R�f'�Sk���F�)@����
R��L�D��2�&[l�b6�)�\�Q�4^���U�����t�P+��d,���΢p��+!Zwm��9;^ǻ}�hx�����2�w�ǂu!=]�r�@�4�Cnb�����b�A`w�7���Ϯ�S_�/�G�Ѐ�X���'L����ͧmc^ݟ@��5���t�U���z��1u66��z4��{&�Q�q�R��%�����垁���a�g�V0/ӃL����=*$K��C���t��(��X��,�fHF>U�A�e�D�����>񮆩h��K��#e�nxt�
X{�$�l�Ժ�e�;��?�yA��At�;��~��5눒�9\=��/r�Ox���T��uj��V���{P�(z�l�b��⸴�j	m�����F�S����#.Z�LR���F0�>^:�L���U�`�g.�ڇt&)���QI����4�&��jz��ްoS�jZ�\4U�d=gSط<�hj<�ʛ)��gEP�e؞�P���vN�ƚ^굽b��ݗ�6�^�$��ᮋ_'6k�y�ٸn`���f2�����W߮�]�
�B�b��J����G�uSez:*��N��%��-7�n��ݦx��d�*�nG5�������`a� S�T�s��9��V�FϢh�����_n�t���h^="t�4Mo�OeҲXǪ����p�y��V�j��3+!��&7�����:��N���.��%���K���@=彋b�n�:{��F�=��x2=�TfC��	|e�L+��޿?]`�I�>��*a69ʼ�GK�]�>�P�Z⎬�ׯ��<���~���1��"|�>��H�u-߄���|hO�8�[�U��FW��N����r3ӡ�Ȋ9>2�l�����!zt�1�x��i6 ��r��D?'$T{�8ЬU(q�za9��2�RX?`l�#Xm?,��������D�k�>d�W���[��P�c�׏��	py`�Pb��U,�-Aҡ�7���8�}X�ّ�[5�{�K|f.��ƺa�����=sL���Uͻ�)�_$3��;���.�f-�b��? ">�:wʚ:���r�ϖ�ݽ�lYm��aSZ�U�C�'������v�!�L�,z���8x�^0^ʿO�G��~t񗿚oe�!d@�[A�=��q��FwW�K�~?��ާjnO!���Q�'
�T����N�L\�R�&1;Z�m�a#��.���Ʈ�ږv�{�=*Pn��'MÇ�8rw�	EB���j,����,�"�K��8З��2�[=���͋�J X��hAп�����S���~v�T8�+>�i��Xg���m�O�G�mĹiw��;�[O��z��K���@*�<Z���Ƈ�fw��W��$��m�2{\[�fE0{��5�E�o���'9���s`��w�ą=J�칒��!O�S�����+#���nXʾ���|�=3��k��݉���e��2�kjT��`�����ZC�zF����)e+}w��ڨ�S��<>�x7�`ivb�T�W&/ �hv�E^2J���.��d�2M�E
aŞ�@!���C-֢��US`��«*禋 ��*��s�.�mYSx��y�x����XX�\G6R�XKk!^�z��Z�E��H�+O0v��c�+Mx��t���۽�^7^t�s`L[r��<����׼���U���b�%-�2h�&��\w�ҮO��R~k��^J��l�ց�J�c��E�h�`���
���Zh	��?Zg�+�������uN�Or�D����֍���x]/��x||O#�� +�{�l�"�L��uM՛"ZE�#rͭ�fT�ԣ[����&P�aj��l`ScD<yg M�B���Aϼ�|�8"�M�Q�C=�T9��\&���nd�eܥ6��A]�S�'z#�
�#�Cwks`<���_:��Z;"[�UX��lCkp�L�/�W���8�W���f]�,���C6m@s�[k�� s��za�N��UK���,=���
0�zr1�xr�Ō:o��٭p�A�ny yP(��Q5���]�u`9��~���>���p��hů���LW�+0�������j+�v���HS:�🩥�n��̨�VK�Mt�$)�����}AG�r����^�����-�yPW�2���T6PXхv�s� n�9��hB6)Z���kѝ7�`����Я��Dd�R4A{pQ�=նG{c߮F��D@�xeJ�=<3rwfe���F�zT\�?I���	ql+���s#Wz�}���f�f��Y
x�PT����d��5�Z@�7�� ����e��T_)��_ �PVŘ���J��ܵ��]�&��N�;/�Ȩm{�RY��\U�!�w}L��4�g�i�?oóB��Ww_��P��8���8�g���Á0C�<.���FW�\��.�w���-DM=���ռ�L�B<g{z7����ء��!P��X���Ai�aK!�g��XqkD�?2.�Ps;�	�v'�}�`�x�*:�Q�v���T��p)��bl-�y��g'ӷSYJ�{����z䄸Ə%s��6v|l���2�+��f��f��+]�����v��N�aR��V6��(��W����t6��i�;�\(\�.CsO��B�v��G%�ɒ(��U���Zn�y�d�G��'�\�N�K��C�$�a�G�k�����i̍��·u�,4L�v�Q-�����j��H��K��R\1����$-�YY�\٢�,��s�P����l,�kp��1\��C*"�%�5��Q}`���Wl�W�Zc5��!����1K�N����R"z�,L�(�J[��s=rŭ���{��F\��9 6P=Vn�����}�X��*Y�6���}܁-���K�9r�5���U�v��M�@�&�9O��n޲�uE�U3�VR���r���wM{�.��8Ь�0ձ�	ȵ���y��!�F�s��Fn�3d��U�ϋ@C 73�[�L[Jsz�L�q��w�t^g�Qx�-;�V�o�1�=b�!���ĉ񾆆v*�ݿ�n*��	|�}�s�-8��7����r�+�ұP7��D��<�AOU/�E��ǀɕ;57h�U�S���욌�:�=�r`�E�O]댌 ����1e|���o��Ɩz'�MY��ϑF���]n�Q4���/#6��Pq���q����*��Q;:��<�0�ّ
 ��{��\�]���z�Kָ��2B��f���ΙC�*m��Kg"�n%����k�:�z�š�|&�^���S/w��K����.����P*=��|�<��J�muc
m��wӦ��ۂ#
.Sl��@6���yw�0S���$ĦưLs.{R~��Vg���jp��+vK%r�M�� �&��GjT0M���"��o�?�ޮ!�mZ�K�������*�����Zn��[�<�ub��$}g���ƭL�������`!�v��`[� �w��gF1��uؾ�\+)�E�m��o_��U}u�RWV�[O�\�DX|/ �n���{k��8���@�8ū�;]c��{r.
$.ˋ�����bi4��ܹ���9�5r��U}F�i�N�z�ٖ���-��OM;I]�e��:���7��e��']�pbJ{�QLy� *}��ݍ�$ͷ�_�T�����t�_`C�����g#b�y���N���[4��e0�MJnN�a��Ѹ�[HJV8�	�90�(����jڛK�>6�t��e!J1�&�{hOnH9�L8�4ڮa`d�X�0�[6��n6�/C5u�۷l��+�:�
��1:�ŉ�C4T{cqy�Z����Q��گ��(���A�Kvkp�ǜn�� ��t�
'z&40WI�o+��ɖ~������Z�e�1�;or�C�-јp��`����Q�_y�^[�A^�ƕL��GZ�pUϪ$$j��n;D۠��N,�4x�BlOH��sأ+�A�����h ��Kϡ�^<����X)o]�f0���	�%�4=�BÖ[���cl��Q��P�bɝ��
W���f?��t�Qu}ZV�q��p;�v3ٻ�c-NN��{'�6����Nl}0�'�c�	�ir�M�s��؜"�M����6<ts��+u��V�%�yqn�����gZ�:r�M�S9|m�BL��t���x��p�mLt`�J����w�.�>y��E�!z���;���U����5v3Ĳ!�{�T��(0�.�[V5���J����!��Y�b�&v u��]�0�[��s�fU45�,a�A���I�i�.��aҘ�e1������i�p諨a>쩆���L�����Y���:�֐��s,�j�f�m�t�ە]��r��l�w j��JޓZչCf02Dfs@�����Ǎ���Β;�/׃������n�Ah�j�w���F��~̢76�_?Y=�4�:F_C�j��Km)]Ad܎5j�V�7��|� �l�^�"�]ltV��ۉk�Y��g�5����ߌ�/xn�bd�K�6Ba�_<��_V|V�?��vM]�4�y�q��N"�s47��'����2v�1G'�5WHg�0�d�Neo`��� ��M,�Y9�ӹ2۽��mnYn7����aa�C�LBއ�mJ�U� r���ǃ�3X���T�_���W�b�GX:^�o9S��EzMu�����Q^���º=�m�[H�n�mR�oM��M�=���2s�1�.�󱋒���LZb��h�����u�P��Ĳ�=��Mk.ZV���%��4�2�[�CGme�x����R����F	=�q�Ӈ���7t�e�����r�����]�3�Hl�lQ7y�]V{=<���o	��v#�df���rHS_]Y<3+����0���7ca�{_��6V��.ӛC�$�Лؿ&��֪�Y���ƌ-v�ѩO�3��8��B�
�t�%y9�z�\������j=�"o\2C��%�?�3�����UC̏X�2�M�Ꜻ��h:�Vw��/��c���a�O��C_8@x�T,����K��#���ܭ�o����w�\�n�*u<1@x�j5"/������#&D*�ۆ�"���^���
)����!Cj�u�u#��T�k���5%��K��VȻ����Q0٪�N&�@ZUAĮd���ڄ���f��x�b�u�����!��(��� ?B��Kh2v�qV�J�º�#;U�%�f����nT(�x�=!��}k緸�j��ܹ�I�T�Ӯj��27nA�e�%wX�F�'��̹�����6���&s�y��q՜ܠܣZtu�fO�yG��X��}�+_S3�Z�s�>�<9$q�s,�쵐������P���G������ p��,�>p��^�Œ���Ms5p[L/�dj3Fe�vV��Z��D�VKc�8cL�Wd�iN>��c^�pB���U�17��n�Ɖ�^�؋��f'Hͫ|Dm"Jn�=�5OU�u(�ut3�:Y"ޟ\#��U3���gëtu��Zǉ�����jEu���f%�Mπ8��
�����Aj�*yl�Ox�r�Ug91>2��[����.�,�Ex����{(�ʸ�0dAtn�WĄ^l���S��U^���̌����4睟8nX:j1K:���ײ	�>�vaX�����T��UM-�A�w���'���3�x���7̠dO�4s8��8U���dv������Ub��ݠ��O�c��j:�����c�@;���J���Z�f�D�|��1{/��]V[���67�ŎV�GCi�>�B��h��{n�Z���a/Yr��4�3W-��82*<����gwC�]�wQE��g���<S��������S3����3
z���`wT>8��77����n�L�}|�B�%Yі������]�c�E�����݁��;s$�{�0i���t�����Ѷ3�#|�>�]}��l�M��Dl��#�P���u6�b�z��sq3�����ܝ8�^&!z�ǳ�a/���<�+ˬh��׎��y����;��g].^�Z��tǦ'dbKj����'�k3���ON���&�sUTH�����B�˨�	�&]�[`Lyrz}�*k3�ٝ`���|�s*Gomӛ�z�7�����*�T����bE�6�v�r�Z�;�%�v�LF��� ��r�ҒX6n U[ r���[Yɱ}G��@'�Ƕ��bR�"��v����H9|�F�n��B���l�7�����S?en.p��Y����=�����?���J�4��n�RzŻ!�B;n� Ԙ����/5�3� �:م�ջ&�]�z�Z�ݞ+�(�c�i��<���택]��y��2�2�e�0�̗Gn�#@qI�+�$�y����	��t���{k,M�:LU���m;�>�E�8��u�HȦ��6���<����<�|�,��w�i3Ԅ庻�܅vG�]�&��$'�rbw�R��&�O���ӾE9"��W&�̎�F��׮��ё����l��i-ݼ�9�����A��g�蓴We�l�8�(wct���l�I:��������!ȼn���A�6������8�I��+:��[S��i�:���fKy�L���F������@�]^Fi���3Ne���%{�K �t��s�s4�����/�L9os��A�2�,�F����Xn8
�)#mUz��''&5"�V!fD��8=�3mI�R��P�%ײ�]�V	6���8�nC��-^�t	����|�`bɷk,�1��;;G��L�;�X��:�i�m�t���At�YO ��c�W_1'\��A	.i�A�+��#�[x�[��n�k�4/����4�:����C��ޮ�7�v�i²��w_S��0��p�Nt��s��.In�VS�u�rP���,q�U�݈b�<���iH�Wx���'
6Ź�xie�X���qc]�wV�'W�Zê�V��+���B��L�Wp�i�bsok���n�K�tv���=k��YYz�&3�����z��J f�����4:�;x3iٟ.�����z�cKb��5�U�� �!�1G��@a���(GR�c��#Omwv\�M�J���f4xa��Dq�k�d�	���c��,�9��.�G7Ҟ�8b���w�0��q��RZJT,���F;S��@{^������Ql�1<�ƅ��ݵR�ZO��n��L��4�,K�w�A��Rn�����[R��`��,&�]�ҵ� C�.W9�� UЖ-�h��h
A�y�����o^܇-K{)�'vvY�y��%{�?��R�L˚2��X���&�%Jo.�ܜs0*���Ck/��#�Y�5�/>ܞj�][>9(gIμ*�W׼�����D�Gv�C�d�i�2�(I4�:Jj5N|�jX��S��5S.�����Y"��Ա��\���PSY��wr��;hmf�;d: ��ݦoCBG��v�AY�i��Fr[�n�)�zi��C��Z�h<jq!�p�1R�̉@���k�0�iXT3 ����0eN��|���Ʌ��
b��Z�)��E�M��p���]Z�X����b�p�'v��i��]u'32���}�����;,�b�ȋ̊��RaI�fp :%^l���H�+5�k)��o%w0�q��[Y���f���\�+2-���J�̷)�E�{�Xްa�F���%�lU*��c4&�7"��N��n��"}W}j>�f�F$x��E��tN��WK�RP��#Fѵ�j�6c�.�Z�[p`����L0�b�����׈b\F�oX����I�Y�����I8Nv�Y;�;��	3z���%���u����u�e�"��)�X��T�YVԥ��be���Qu�rl�~�����/(����
�1R��\B��-3(�E�-*%lE[j�U4F�`�V��κ���ٳ�������Cb����^��!-�k*8�r<j�T�OZ�P�N�Eg�'��vvv��
(����Q1
�%�C�X�PU�2�s3
L`QK;;;;;:
�gYr�2�i�i�QC-DR�p��mTD�TD�5�e+E��-�\��Q1+��al�\Ph�5��g�2��)JȊ[�l�E�eu�%�(��-f���m
ݸ�s.��EH�`(�X�ږ�%e��k��]R�ZX��Q��ը�c'�k���ekh\�j�Q�G�2�
�b�S*�)R�j�Q�.��Z�����i��5YjТQ�B�qr���D��I�ܕ��F1B����Ҷ[akEDQQ{`UTu�VQb��S�UD�"�(P�>4o8�ػ��1���櫮����RN��J��>͜���:��or���[a�}�8��a��W[VĻdnh�/a�<x7���q�C�[<�l8��5���a�fӾ(guf�vLӹ݋%��F��a���N���L{zr{���}���6%06����i��z0%,��׎4F���gv+�9M#�c�z=A�F��>q��D1��5#K�j��/fZ��O܂�y�T*'���f��d5k��A˻��4wm�Q=
fV�G>��O�X�3w�`n�m��}��J{kt��#�`�y��h�#9�ŻO�<��"��U���L����o��ɩݳc9���v��%Cd@ܰ�����f=*+�؞���FV)`����.w��m1��W��lV.ԓ^x����<j&�y�1���=���m5H�7 6�Q���k��RL2��ѳOtpv_���I^��4F�<4��sm��އH�R��vo[��{*�ÔT���W�����T�=z��դWf��H�����v^f�:�T��^Vi�]pSI-�y��8u�i�V�N������"��#tOi��Y��35�}Y`�\��վy��Y��b�K���]
�.�1�� ��ze�4�g2T�t�}�̳��|>��;�ga7�i��j�0R��������%p�t�7�]gm�w뷋��G�h�`���R�WR��M�ej��h\��ˈ0i�+xS���;��3�����P��ΤЯ0~�b����^��t��?����j�[7��wq��F� U��i�qz�m!�g9��u�-��=Zp�_6Up�DQ�v}�@1=iB���'�m z��lpœaM����;������&))��\oU�e s\�M9�v�ũ�w���#��{s\*ilL�v��z�R�d.~��~ń�p���:g7�?\�NZȕ2�����E�=d5�X�Ȼ1ض@��<Z�o�e�qyI���"v�S���-�B>-ex�v*��{�_����h֏��3�9�+n��u�n�W*1Ũ/o�Z]�v/:���d�����\
`l���'m\Sy�6�-���yU�`=��uK�Y���'7�G�,k�zw:�'#���s\r��!���UJh�Jq55���m��)��C�L�Tt�oV�m��BRc� �u����ژ���"Wn�I�;Z�T��.�����Ű����^�B�(�+����� �%�Ds�^�<K�2;�GF׺��	Q��j@�GA�N�^9�ܾNS�>m���cWW��V�\�/
��N)�+w k֯o���ꄼyb�	�oq<�AzUt'6*&�%�z�UjV�W9C�ʡ�:j���yd�tw���/+9����k���m�oL��-��e�Y"��qNM\�n$׮F�j�׭6+.�akl�:E@��pyW��)�u��Kk:�c�"��Z/f����r�G1'v���G�_N��V~�⩼�C��>�Q��>�l�j�n�+#ʺ��J$w_�t�D�_�ŊF�\e������$ND��m����إ��nݐ��-�Ȱ��7}�b0D��F)}U;��!�Oy��y-�ʽ,q�r���x���M���O�F�i��ϛQ~�������b���
S肍OG��zoyr��z[sl9w�۶U�>������n��QCHy�wI�X鵐��{���m,��8�G����w������s˫$�o������`퐍r��Z�E/VҪǪ��NPH�S7�y4�o;�⦓ǔ���&o]=뗒4����^��dZ��\l[<wGc}�xd�'N�f9�����>yW�C�#�md�~�4u��N�.�M�w��B���K[�cI���XS�P��:Cb��WU�����HSe���T�&��l�𛛾 _v�W�V9�`s�}>�k�b�|'++��E��F��k
�ޜ��5CU*=���[_7�L�**u�tx��/l/&�4`���3�[d�B'4��l�.��oGs`��
Ϛ�i�َ곡Z��Ba\w�UlWmo@��Mݶ"j|�����l����$�oE�-��I.�;��{�(w^k_�D� �!�g��@nT��~����%�4��)�^&�}Mb�3{tռl��U[݌�6i��Mǫ��Ԋ�q�7`kn�D�9{Y�_)it��V���4UՋ��aw�b�N.a9�[fG4F�Qr���#l����>���/�D�[X�f�T��K�狲���Y���*��/�g�ʢǦU��Sw�u��Z:\:�U[wM�ਖ਼�z�x���ݛ��́-��p�v��n�>��Y��sP�������r�����&��CS�nH���%nkd�N�V:�0�q��od�es�},T��E����������)�-h{Z?V�l��0�Ghn��S۷�l�f���������YlNْ���ݷ�VC��B�X�Z�%^&�AB�Ż+���¨X���9�Ӻ..�Cc!�nv�ޛ�i���Z�IN�����M���Y��g3�c��i�H#}�#�oH�܍��Z��W��&�!�5��1UVN�1����dKsf��qe�Q�J��쳵�b3D��!g���Ĩj����q.u��l�9w)3n,Y^����ޛ��o��}�GHѶR(T�εln��9´EA���>�K�C�ݴ�-�f`��-�|�VCWu6���悉=2DgvA{̐�����}ql������8Z}Ǭ'<ƃ\S2��Wq%�G��:�4Ta�\MvS:�粮��ڱ���T���,mh� w`�z�`v�7�u��P^eT21�84��L�Ƚt׫Owaϒ~�����*���I��{Qg��d��r1/�M`�ǜ(���p:�
�-��u�n:��|"���b�����tِ�Ӹ�~${t<]Z�K;�rwx���W�=�z�]�5I4^>1Kg�㑁�鼻��ڊ>��]�C�Ԃ�!�2�F�+bk����U��*X;�S\fӴoS� l���zE���5��A���L����:���Y岖o�\m�z���H-w!��)��������Nd����W}�`L����.�A��r	�Ҟ��kQ���n��`5K��=#�FЊ��9�U���j���@��qH���Ε�a�L/�R��Z�U�A�\[5=���W�֞��� 6�j��k��)l ؎�m�H�[�UdS��Y�X�i��c%�j�|��]�ɣ��d��y��G-9[�v���jb�����c�f�\W�� �\�{ �-~��a}K�4Yiyq��6��(\�v�K�
/�.�{����u�x���-�J�r��~���JG<�ٜ��4�.K�����EN!g��X-kCn���NWh$~�w��'w[�34��7��W>7��E5r��ũ�_y��ѱ�~Õ~�A|}3�e��/��t�S�T����)/��^�0{��!EˊU��-��%�/7;:Q@޾ˊ�s�G-�Q���o֏o�񉫘-� JƢ������	�j�{}�p������c{T䐕s�6f���v�yvs�Џ��\s,��@Ջ�O��������Y����,'L��L�����ʓ�?zk�0�v���L����L�7}�Ȼ�^6��[�Ổ�0��3w7����[x�J�⻨��Q;�^�Gd�>����e���g�DB���U���g��+�)���f4���k 1Gk�Z�K<^�H�lR����* x�L�a��[���7Hc=���t���Pb�S%�W�G���IQ�Y�Op�\�52�&������O5�3�c�HJ/zv���!Y��2�V�-gm��m4#4պY�Kٌ��!�����]	J.'W���Bª,���Tz6GNo5�����h��R�&�z'N%�����~�T;R�0q�MD���F�q�y��s��V=R�A+ʯ�z�Z�M5��+�hU����y�Z�I:�l����s���Y�{��*�����ݩ�[����[�W�/eE�|�k�ɶ�o:�Q�i�Z�{�e���E��A7�W6a�gL�mf�*�B��18��!��ٗۖ�Ĩ�v�؜(�U"vx�E��º�z2�ְ����^��ݹ���cJ�nhu�ǯ���=:yh"�-��-��՜��Z�d��w���,����9����Am����y[��"vnchĭ��|d����1#w(Ȟ��Ά���
�h��)��Iq}�#r��6Nc!��,���bٸ�״D>k���Tϳ�����⫸�vX��(՗�-f�s��ފB�af��a@��*�w��ly��M��"�f��Rݴ�v^�ݝ=5<��حse���6	�خ��ײT?q��k#��ب��~#D��p{�D���Dt�4�>�i��6�G�]b�]�mAr�5\>��z.v9��ņ�8�壷!h�e�a�8��M���
D�P�$B}c˅nϗpX+�l��{�
��L��Ʀ���v��*�׈*8�L�3g�Onr�)�R"mu�^f4��l� �%�@*��ex"�rЫ�tĘ���)����ǽ�yӷ�$a�8�{� �Ҥ���ͩ���kz��4r���P���y�9���?�����(xA�}���e:2���>}��R��Ǭ�w�dW�h�O�d����`�]!웧f�/n����S��W����@��b��k�v۴8pC/"Pĉ����}M�]=o}�mû/Mޞ��fן��SzZ�I��k��VH��l�z�(�4o`��m:ރy;�67�U�g���*���8R+I��5��c2�˖�\�W�GbG�b��*Қ���u"�HwWŮ�RM�ޟ��u���[�)����X�������R��R��m�Pz���iO�dH��y��cdH�{̏W1��#�n��ڶ��[
��7���v|�ST<��o�C=��`�7	�uI6�Z	������z�d	ɎA�*��#k�(�v�S��s�&5oP���r�}\y�t�L�t��gy��j�pȍ})>�WŬC_ Xb������7�k�o�:�e^�ok�O=-���#�Q`N��<B֖�#5�O�y�2ޑ��T^{�L�0}a�Zzgd��;��K�"�)z]q����?|<�W�n�_�ԎuG�@�H��݌>+e�2�C˕��r�2p�X����}��m�%��mn3�ρC����z�O�G�pL�d�-s����4VoT5����[���)A�c���cښ�"��	6�wih`\���J��}� +���}������	t�t�r�9>w�h�;m���F��ݥ����]{BT�s{����`u��h�n�?^��l���gTc�����|{7�� ���lɸOt@8^��l�}������ٖ�c l8`b%e�܃�\,x^��6�g3����5� �G��L�˻�ƋN,H���M�܎��-q�����Vʤ�Β������j�=SVa���L����(�U=��f}]������Y[`u_zq[�t�܇���UY�� �j ���y�Rm�E�)�}^�PR+��4�RX����P�7&&[kDE�7�U�aU �EȄb��ҖޕT�x��\��?<�֡��bs.k1&]n��{c��\�Yc\���lrW�wmBcp��&��'pT���䜞 wS�*��r�<�Mj�_sGrG���㧚.a�A�?�ã��5�I�|�X*J�Q��	�Ou�����JO�Y��@]ҝ�q�'Gg����N��*[д4qcZ�.�6��7{Q�
��`��3����y;.�v��P��o	y�[|�=V%>�V!K���,hyB�w0�R�3�]����M���F�X�ɑv����+IfNh�jI1jY���M���ǳ�Bc���-�gKo����i��Fj�%��QV�EcZD�%ǑŹ[���6�/�]S�*����D�0A�z3�ڷ���&ɽлH�?[�����c�3�mLq���K5R�2��eg-���7�wV�JT���;x��6w3��+�m�]�ǎ�>�Cw����$��vB6������v�ݕ��a�n�b���%Y2�#�#�Dl���Au�t�p���kb�9���FR�EAѽ۝·j�r.��M$w1)fU�\2�9��J�<��t�6�ϱ��h���k �䰥ϕ^�M}7'k�y�U��@,[�V*�2�[��^�-U��{:J�Ę�F�GC:>Ǝ1n�el��]I��6��W�mb;?.a�z��{�\��b,���5����Y���數�F��Ŵ���l��
SjQ�0�3&�r-kNq#��֓�o���N�X�t\�#}ϙ��ᙵ.�^�q0�^�u1�k4�g��������'�:"��HL
�q��b�KB��͌��Vv��1֗՚��؛\��b)G]Ysz���X��i/��i�4�C7w�"�mx�S��so"�.m�w=��y.���x����7��2��pl�kq��W鎡���|UꋤnDU����B��:;寻�z��i�qQ���q�ή�3���|��C�3k���K�r�l�ׄj6��N9Y�O�fQ��A]1�MB$�Y����!2W+�Z:*%U��o�AĨ�S�Ʒ�<�,���v�E5ю���,vY�sTr�R��q:�2L��
N�1K�h���k��O�X��{���b�Ӵ�a����/���e���7�Q	ױ�x�$�Zqʰ��So�7�N�A�뤘7cݥ��7F�"�S�S9�)�7&P�Ps��քҼۻ7$w\���~�[֭�6�-[��b����z6�>�eL�p3(�`8�@�8-���5��Ju��g�-���i"��Ρ�t��:�� Ei�w)k�r:��j��x��H젎-�/�鼓�E�Fq3��u�G�ڋp]��3��+���깓��٫���Y�Ժ')�;��W4k��hD�g���9Ӟ�7K!�8�ŀq�g��}����ܾ�-\��h����w�^��W�/�Cɧ�C�X����aT8��M)�w�L�h��'v�x��W��1f��cJc�)�D0gv��gv[���ܳgn�������4��vѰ[E�h j�,��l�T���T�c%]&/��i�0���Q�r�!�+��5(�G�,���[�dƫib1Q�UCm�P�6d��������q���E"5�u��m�)�1q��a[J#��bF$A���QS��ƪ(5ܩg'����ؼz��*�n>�R&%D��1�(�w-�ZkB�G��h�֨�8��ƅ��'���;mE:�eC-Q/��`�(���)G/�b����
�����M�Q�ɳ�����^��;�l����v�fa�Ɖ��Z4��U��-��̣*UDD�F�G���Ym2�J�]lnY���9h(
�EC��(��H�����¬m�J،Y�EW-���ֶ�*��LJ���Q��D^R�����#�`�i]w+�W�����U+��ĩE��+����V[UQ���ŏmN����imH����6ә*�V+��b�7���(ܸ`'�v�TyB�]޸���vna,�G��冸���neLLʭ�S+\\̭n\\�=ʫ��{��)�Q�[S-q�婖�1��r�-(�
���q�-O2�N�Y�
	,�x��$Κ���u���Nw��'�)��@oՔO`W��Z)�X����3F�36��f�/�X:�p��׼wW��Be���P�2t;��<]��q���B.zz��Ϣ}hGxoz}pnc�M�n��%i��X6���7����J|�O�ۉM���Kn�?:�</[�{L~1~Z�{��0r�,m�D�֔*+�buLힽts`Z �M>��|cU���n��=��!�5���3�63z7�g�ST�����S8jkva�a��w���p���Au�KPdL�Y�V64�7,��9/���<��NQ-�Y�ݲ!m��%&d���o�����	�d@Zg٘db���;�9��[3���������غ��;�s��!�z|�!�������ê��V�$�b�Ѩj&h�dgOGl�v�'[m@v�%�AT��:���|T*��BWq2��T�Zo�T�q.��j���:�p9�C%Dj����9{����W5��D�fνp�P��&&��kx�(��'�Y%b�I�ǖ ��4�����N�O]2�rIO�w�&KŰ!yg�#�n�ؼ�*��3\/o>{�'

Z��Jv�o0 뾡��;�!� �}�v�BJ}כ������ٛ�����*p�ƺ��N6�aL
�|�����{&gZ��ޖ���VҚHԲ}o��悮Nc��e0��3x�2õ�������wH/�ey�.�)+�R���+ܑ�mg,4Q=�4�}���7�/6jTb΁P�3��>"Ԙ��fc�� Z�ʼ���lz��ɲN*���mW�wg<��
k�����c�S(����d3�����d����+#J�WVVO[�������/!�'��t�<�:b�)
qh|�wJ�a�H�P{�#p*;SHk����Y}�y}����Pa+Pm&}��B�"�cm*��LO��H��ͫ�:������v�n�E�h"6@�(2llPٴR��o�~�Ej�u�B��9��#��R�P���-���k`����ڍ{%C�Q;���MSu�뼒d=U�Wo+C�8/���4�>�,2[G4�2�l�����@�q3��*T��!H����^d�b9.�/��Ll�d������x�go=˽�(7�[��v��	>�L�79;v��뫙�k�N�v��mI��t� p�,�1e���Mt��L������ڜ�)���W^�ͬK�9Z���]Ypl��&�Mg3�F�W�j��^�m�9��FX�b4���g�b��O-t������3����_@�]/��n�V���,,@�FCr��P�o�����-{�}[�0z�ӟF�17Ɔ�a����Cy>��
����1t�E��Gg�5���m�x�kMi\Mu׮�p���9����M``�"�n'V��vCz�:ԇ9��f�����Ih�4�F�����/���8@{V̬]���\�����`���շˤ?KR+�>tC�TŪ��(���Zd�H�Ԝ򵹩MM�տ^2��r2� �l�1y��EnF�]�	6?���V�y��>B�t�G��׷c�lM[O�.jS�c(�����V��Eߗ�v_�ʲU�i�zCt^�+v���ގ�r�3�|�+�q���x��4j�#���#�y�i5��i))҈�)[�ue�rp�O%M�ӫo/t��_,Ƹ�H%�ӯp��m������!Ӣf��F���!���"��OlO�;kn٧IA*���t��F�{urً���\���*�mwnVY�(�m�c\��,=ʱ`�ꍊCa�V��]��xxU��p����vW�z9�Cl�� �Djޯnɑj��;���z�Zsc�>fof���Hg"U��v*ӌ�قgO��'ߦ�G�Z K�O���i����VPf�^;�{��9�8����������-���Fu��tp����阼��:��\�4������3�=��/R��&�]yp�W���~2����8Vr�ǶJݒp����f �ܡ2����hn��'p��l�c�v�9�>����Y������׭��:9�J8]��`}�<w���ɭu�w����O�lL�3��R"���v�cN�n��ݱ��Z��,���M�j��w���d?�;���|��X�|l��߸�y�O$�O1�Ks��Q��qp��4� _s�N��j�5�32�E����堮G������h�V�"���?�`��m��4>PL�"X	9Ih�c�}��P:���H�T���v݋ֲU���a�%q�Q�O��)����H��6�wJ���8u�`$�@#����ܱo��xo>M�k���=�y�j,���a��3���I���s|K�v�sd��]z�r�z�;II��f�G��=o0��N����&F�Ǫ/�.���)O��ֵY3�V�R�ӡ]ݝs��Q��bF��,��l֫J���q��J�+��&��u�h_ccf���lӼ6.^��^Y:�1�������k�Z���"�^¨�J����V.�&�"��Sp۳O���<��es��t�>�b`�����Ʀ�=����|�VWt�%}^�^<z�0�i�3h�Jڜ�ymJ3;�<:���y%r���vQ*����tE߻����By��;u���i)��w�7��t�*x��t��PqX�����f�>���v���v�!��C�Vzgcc:���W���4Ty�G�2\l�F��UC3oe��݆޺6�A�3�,`l���V8H8���}���M�y�U�	��c��W��b�_ED�4��*_vê�o�<�zfXb5�L������\O��<�)��.ue�n�r|h({i�L.v��q���]䕹P�KHkm�MC@�ֻUo+�^A���������}�D��ӝr���}��A�1����F �����/9�f����D�w���bm�I�A������F���|�i��.g�7Hc#a���0|�깽1ȧ4�Y��f�g��8��*��dl�܏W�T��zu;�C�G����6�Gv�-�4_�[A�[Ie���fo���w�'TC���r1C��y�-�Zd�׃����ڪ}	l���5�@��n��W�XH\����n1Y+gk��U��DI�vY��L�*�����$��P*�Jَ~�0UBd�je[�:�C�Ds3w�vg��m�N�:]���Z��l1��~��gh�[g:4É]�E��P�U���W����QY>k�Ty���X�\u�br�ѺI�!�5�h�"�Y�L`���qɠ3��7����)��4'6����g�D�{&�^�k0��6Da��@|3��mE+�nߊ�
����D�vEC�����l!
���$m�w�r���-�W�׷�Gt�4Ò]Gs!.�j�N��ښx�+/�k�wy2�V�Z�  \�enQ&;��S8.Тq��@9�F�&��h[uu��%r��oSπ;�p�fN�:�糋{�����`GQ���U�o`�Z_��\i���|-�����c��+!��z��,�:?�����������3��<Uz]t�\g�m��&)�)P+4�Du�������z��w����L�`���z@�H���ޛ�9��=)�Ϳ���"x��'������Ǡil��p��}��C�F`�5��ѓ�rBz�+����/[D6n����dy�doI��g��Ţgm��h��e�'7xP�`Ӓ|5>9�ɏVa즑}�k�h�g���;CeȈ�b�V�?$Z(FnȀ�=B�2ё��:�@��-���U8�jM���h���=�l��L�)8v�qwm��@"kW������^ɒ/s��ۙ�ٝ4��M����F�=��QP"���pfPV{����&q���P�|;N���E�z���>���~��\�|�sT�7�4��������S��N�r(��8�T����2�\`���v\5���%6=��?s�?U�*H��zez`̃39�XQ���Ȥ�\���p�qW�=��|n��z-���U3������g� 7
�;�U�X�ɺ�b��b��]&�"�ݡY��QS6��m&�QPnړ&�'v>��G$�W���O?-OG�5M^�ߒ8�ҷ���]WUf�гYP��S�Px�&�&8^�k\R;Ag5OZv�,�8�M�����yU�3S]5�3�MK�H���S!�1����/�v(���3���US۶7��-v6��Њm�gE���F'�S��:GhG��WD�{+R������6o*��l����^ð8�T��j|����oh<:���!.m8�;���A�4U[����A-%!��Jn;@"흂��8�O-W����/5dOWT��i]�����]���-im�Ft>m�\Y�Y�6M��Yv�g����^Ȉ���]�p	���ޜ��nO���v�_E�	�W{y�G���hm�"_H����3�/#Q��'[��Җ�Y&�̙�s�OsFs��96��L�v�"ŝ����M���
��"�R�֞��Y� ���~\5�8؛����(֏��Q��m�ֵ�A�[c�p�G�b�rV̖���sR��v,b'�$�EE�:�J$�X<��p<�Vyuɬ�vgns���hf�w;�7��ɫ �A�)Z��Z�Y������+J>����O֍�$�K��tN���k��~�K�ñe]5���imJ��7��{�N�h��j!�{y�_M<���6� �+�����a��V>��9t]�k�U�v{��8���am;i�V6[���J�[C<�]�����֖���ԁW6�1����%��Qӆ��t�ᔊ�}��M��P�;J/v��wI����*-�Һw ��vP���+�x��]�����ͫ�O[m��pU��+�~=�&�Q��j-��nko,6����j�u=�e2��4�b%�0������>�j�{^��ۅ�j���z;V"w�n:��ou�Q���P�4?���/E�$ܛ!O]GH�ѵ�m�ڜF7Ӄ�;lڮ;�I�r_<WK=�lf���hk��8���q��b��O^�s�Ts�ʄ��ifg�kPy����+0y_�vE�P�m=�̙o�9��:��Dg����ǖ��.�vC���3o�5]�w;D[�*�w��ʒ��yK��wc�r�	t{�\�{/�	g)Y�cz�kKq{7[v���we��Ҝcb��N��Lk.�v�����^�MI"�T=�1v���ٙm��\S��[��������O	��e��{n/���d����a� :&b5(6�7��R�����Mk�a�VeN���"vl�;�ũ�<�I�h��`Fّr����Gb���4�S�]�*����UK��l�l�N���<�-�.��j3a�v��sG���ͩ�~�/s�7�i?��U�:�=��j$t��S�� l��p�z�V�2Ͷ���� �j�Š����h7��-bT��:����g��x�p���0��2��ޞ5�1J���[��_U%wni�3xB\��RREj��Cð4A�2�]
[D﩯x��i
b�;=T�Ml{0�5ם`���2AQ{-���m�+ñ[�u���D����'�tC1���FtTLIe^�U�]�f��溮���E+s��dmEω9U��)�Hwh7���{�U��b-�M��3�M���F+���c�rJބ\��f�VL��(,�V� �(J缹,��f�aI������d��6���:�聩új���5m��Q�fGw0<��`]B��Y�	�抩��P����7ڸ����(e��;�v�	��]AN�A9��.����8�n̚��՝�
B0��N5�h��Y2g�ׂ�q�.�SI�!�4�%��B�*�p���,�[���r�Iu������G2i_uZ���n�9�5>$;V�'+�"-FWS5�=��N�ح���.�1���ED:�f(*"l-�T�*�l����ݗb���v�\E�Ql���m�)KWR�t�B�)X3L�-#�NDٮi��3/r��N���Mp�����ꚄT�[�,�j��u
�ģ�Hǣ1�XҌ{fN�B�WƝ��q<�f����F1bb��`A���nZj�N��U���8iׯ3ŋv2�D�i8�Ǟ��w$�9���zkh�yϻP,T�|ăR���fM�;�7d�W7d���|��LCGwy��.d�t����q����>|2��Ϻ��"��56�&5hԱsN��nNΎ��^;���/4��%=vi5Υ٬�ftD7��^��~��颴��PK��km�üW)�E�/�32�U�t;W��rYx��kDjK &�Mns!R���$�Z{0uݷ'�a���(G��8p�g�n�C�e��Z�_h׃�ZV�;/X��&��į7�F�̶{��ٮG;b%�ɖм�]m�D��<÷�G�}��'%�f�P֢7A��^��v��|��k�B+�{�3��賸[A��ޞ�jXX8���R�q
�U; ���'�(�㓕��m�"��-D�L��δz�Q<�իb����R��/*�6[��Ŏ�ڂ��*F�=�V��q�3j1AnS�@w�D�NɄK�tg��V��Z�rC3,�b����ML�и9�gO�'G�6�}נ]�������*�j�m����9
N�q�ڋ�f��xE4%3Sf�Ϟ����������WFͣl�Q����n��`�:P��6B�ŝ&�F�*F�^��y��Vf˭�m��b����읍�,���<�Bv�ީ�Z@b�=\:�@��U3.��-��$����.�ꔢ��7�W����P�]������ie���zU���BsK��b��ռ�z��na�S�y���vIi侾�Flդ�1�N��m��3jJ����l	����n�pȊ4��˥��&�#ڝV����i*�K="R-�P���u .�up+�:���f���r��33�$ �.ͪ�ӷ�]�[5�uB�wh��}
�t���]e�)�si��i��U�{㘮�vs�.7�y$���v-��:gq��ٻ���ߞ��}���{�#�EAW-��UU�*ĩ�A:�֣1Q�2�H���32幙ͨ��,T�7La����<�v^�r�����x���Q�����(i���̳0*/n�L��E��V\�f�G&���'ggP�)^\;M�\Ţss1ZqU6��3i��wi�Mۘ�ֵZ��9<�NN���ㆲ���r�̱I����..WƮ2�����/02Ƣ-�0������=*��m��%��U�b1T��`+Zڶ�UKV��l���'�s2�8�T�B�
�jb�*���Q�ylZ�L�֫
�p�YYYP�� ��1(W��������!��b����*k<��b�d�Z=����00�Z�*yI���)qG�t��7����*��Y0Q�(�j�i`b�+kF���E�*��<q&��QC�
����J���G�����e��!Z��RcFT�PbCB�Z���iFӭ����J�W��PE�3�-%A5D�"F��7z'j�R��2Z��wn��b]E:�23�K�&:.+T׻�omGurr��ˡ�[��z�k[����d��
����v��4{?E�]$o��:�j}4�>��8ʨ�q��ߦ�9���Q�4�{�7BX���r���+|��2���8�k��`�ai���y�%�c2}hQ��Ӿ�%,�O+��X��2:�t���h[ۛ�Ω��>C���T�*�k��x���(�~۱<�-�bC�ˀ�t�����zHu���rC���=>�ȹ�썔���LCuJUY�\<v�i]s{e���D��:��@V�|<����`��߽q>O���7;{C"��%lt�i��y�V�ڜ�ݭ���-���l>m��Gj4D�io0a;^���7}�;(lI}&sḬ	�t�ט&Xg���Ԏ��q�y���"% �&��u38���A�#Z��>1����u<�6�����K�Z�~�n%�K]�O�1:eLT)�1�������ЎRw0ٶ��c#�;����_eke5��8	C��2���{�e�8 ����]?7gÌF�ZD�%4sOd��e}dЏ�S���k3� ��X���*W�[떯/�އ�aZ8�+�������7�Xj５�U��/y�~ Nu�:c;�?~�!��Zx�f|"o�{^f5��m�"A�4�����M+�C���z�ײ�p3��k�\��Vs}#R;���A�&���3�8ނ&����>]n˥��Y��R�g#�g�W7!�&�������oSP��!fQ@�G��ѻ�UKm�=��U˫;�L����י��>����3ho[{cmϸN$�҅��s��nUs>6���YDn��}[4��Lg#|j�/eT{a�є�2nz��Y^�%�zՙ����ʽ����귨>�j�Ų��E��ћh�b�F޹�m�/"s�ꈾӬ3��4ݪIm����,�q<VX��Zz�ѻ�@�fgqQy��lC�H����wux�R!k������u����sozht�hF�㷄WH��5��Γ��%u�#��k�^0�3��6<��Ua������tX0���л��.�125��D���^�d|��Wo�L���;�ޞe�k�;6��7̔e4R�ETWAQ;�3Aq���c�촥nX�/"�w|������zW[�z��k�� &ui\��XV̇����{`�Z5[I�R���Ы �L| �{��|E�Q<��w;�)D�x�x
0�����òq�%�9��c�L���^��^�;����R/R�oNOr�=�ӱQ���Y�ݞ�On�9��q��.V�����9M>�/�w-�(���%�����(6�m[�	�>٘
̋Ѹ�G?f�s�5ԩ�<�8n��T_��z}�P}��@hy�c�����T��`	&�;���C�'��t7G6q�]�]t�W�w־�ΰU�[���-�l����ɺVw�깮��f$b�B1���d��n���G}{N�'u쮘�eV�&�����Ã��>z��[T�>��J$��Im�.}���R�Fڋ����ֽ��;�6-5jn5 =�H�T��-t�6�Ti�J���)I�j��=�)1�1=��%�L�58�B'�}�z|۰�6�	"MD�`���5�;`�N6�͙�����P�p#�Yjrҧp���8�=���g�z���Y�n�/%�j�Y휞X�\����6������wٙ�ʁ����r�2����*�J�Ao��ڗ{��5tk�WwNk��]=�a��'k���:��o�*�3�5�i�����ЍJ�.߳.̓F�{_#L^�
���4����u��Q|n���)��r�̚�sz^�:l�8GS}��I4<ܸ�d�WrJ�}�����ȱ˸A��YX6n�wp����[dR����P�\Sg�%gQ�e�t��=�6��#��M�i�7[;]��D/7S���螲�W��X�Ul�s[�*O1y8ov�4�Z��Xv���q'|�{ͪԢ����Kt	�jxנ �{[�Ȗ���X�'�fI-,}{��#ͼ���8.T�:�m��m\Ns������<��ָ�y�:��{m���Q���~i�-֭�y�d��;<ã�k-OHs���c��l��`g�@^v5�E����ӟ�q渍B>�U��י��$k���� ?\e[�+�/
ߚ�.t����a%�r�bʋ��ˑ�Y�������tʞX�h��ԅ�#л7Y��YyfYi�9$L�nH32��Z�Gs���`��3�]׏t:��}���"��09�����ζsL��+^<��5(�]z�d�?�Mn�K����B������fׯ�z��3*Zw�@K���W#�Z�;�oP���yȢ����/x��R��%��V��f�}��dRC)d�Ä�kW�r؜���w�&��'u�A�Q�U����t�DǘbK5m�e��gEK�U�����{�����,��Q
��D]߃��+���4խ<.��O�rt���whU�W�EG�$Vc�ίGR��@��V:�9�;���Y���˫���e�{��U�9k9U���O�V��\�K^#����>ζN�m!����כIJ���*�yWVM{��wS7��Ñ���Us��/����
�ö��U����EwR�--I`�O}u�E�O��rN�G�Bm&�7e{�\�Vf�`�p��:�/";�_��NdA�q6�2N_u�wQԬ@�f� ��!fς�ޗ(��gt�7M��?e��{ �wy[���M�K7�)�0\�v�yj�t���zy�yWK�ѣun�ًL9@�@�2`Z�] �
P#�j�V��5D]�Ad��'[���5w`,����q��0w�}�ǯ�v6�.8��ۛ�s*S�<=��8.Z0UT��_���u4�n��q^�:��T�����߰G�|Qjշx^���܋���]�5Eb�e�Ǐw,�a/��\��6�~���q���G[Oz2���=��`�d85�)>�] ���yh�q��g�P�P�x[�.ê~!��j��n�C�p؜��"QB�3 #`t���i��N�d���zwZ*�p뱴�|�}�mZ]�<VdD�*��;I�s��vJ������bp�ֱ�hW�Y�0�4n�����/ϔ/���14�v���U�ՄQf~h��C��/-���B&M�쌵��.r-�t�k��kU��1GN�iͦ�Hz��Vr	��q��Z�*��?Cey���!��uY�0�f�w611����-�S`gU~�K%�G)WW	ML������J��T�C�s�^�N	��I�i�sEB�qK���݄��]�-���YL�m�/.LlH�*���:k��n�]X��1$s7^�Q�M�j�9wTvSY��Fv6��I���w{Bz-��v�!T����3r�ƴm��'_�ÍNB㪚�wG�)�a�:�]5���%�U�r*xU�Nǳ�j�PY�;gd���P4+��g�i��`����U�ꖷ�M�l��Mo
l]�5�CX;�AMfh^���i�ڳ��l����i���X��_���;�Ot�d�A�1�Ϟ���D-��ź���.v��;!��u�#V�����<Lcb�݂1��y��"��+�.�U��f	�,�g͝K��km�l{��*�U��<Đ�[�)@��l���V�N�(��-��JY��w�c(���k�������_�O��F�x�;�qՔ�=�!1�r�k�ўi����{ӗ�759���C $ZP��[	�*̔t��x���b���ь�9zɃ��gש���a���fDf��n-Lϱꨦ�zxH�F�^n�k�wE�9L4� �ӶˉW��h�E<S�u���?�i_'��C}���� ��F�qn���	[��n�]��<�g]!�
���uUך8�0�]sH]޿,~lv#Y3יw�����+���͗,�U� �c���nv;]Z�l���#(BÒ1�Ѭ���zk���G��\�ʏ�z��+w���������K�{������@��H�Z+�-��8�p��$��u�wnd]�����Q��^��w/9�Ce�[N�4ө�9��dˍ���-�
SZ���N5�vX�)L�QG+TV����R���mQt��9W8��̇����I{!���i�i���Ū�хu܂��d��V��Ű�P^�\8M�s'�����{-&(v�T�MA�	J��}�x7���9�bb�l���M�wbJQ��r
�T
������������]TK.}�	C�h=|;U���઴û �ڹ���e���5I����ټ�;y�DX�#�Ǭ���7.4�h��t$oh<�uPk:�Yz�Bn�gl��6T�|�C�
uV��P�[˗���>Y*�k�$�V~ʬ�m�joF�O�Ca�q�r��z=M��V���ϔ�vZ�XXw�K�bnl��u�ob�|7B�O��߉٧y��߰��RK�3޴�d�+6��T#ۚh��ImvG���
�
��c�Y[F���s}ة�֧_67��1���q�_d�������$%}�R�U؜N�rs���:�3+:��\���6ue���L\�Yu���-�N�6_��Y�}�.��ޝ�954w�a�#�^�iQsyw+j�'�'|�24�e���P״��]Q'g�r}�a�����2��틷Ul8�O��Bϫ?uwq#�V�������=�Ϊ�(�)�S"4g�d�|���7�c��0�5�c��}�Ci��m�l�.P���E`w���f�jˍ��$���e�}�gz�\�32_�!�� �+�*�	zy��-�;ߧc�/��"���r+M��|g�*���������-F�f*���k�m:��Y�U~Uހ�U\���|�^����Z�k*�s�_I�#�Z��ʢ/�D+�q�3c��5�j�N��.{;��Wer|�뱩e'N*�J�~���������5�1]6�9��W
�ƛ��=j���(�G��u�\���~�~�LH0�U�&�0uS:JC�'&mbjW'��:}�`��(U��9�Ԡ�+ݪ�	د��%tYGa|v��lD�b��;k��Z�5�2d�A�����N����L�7b��o^���H�̤j,i�m.%T��>�7z�D�7��;_��S��+Շ����#�I�}��+��w�J��R�^N�Vñ�.�$����"�oFA���Y��F��QQ�ռ�ái��~�3��v{[���������Oye+�"�i�W��l:ޣ�줦儙�l���t�=��I��w{x?(�$v3<; ,C,�W�"
9E!�38�e����$�̮�k����B̛m�veb�o�=�=r"�M<>�r�$�c����w���M���Y`�YB�6���O����g�-\���Ҏ�.���["�H�z��lW���WB��t�~�ч��Q�0i>�w�3���}T+��g�y�^� �B�Uc���h�z�lyTOF1�u煪;:�:<F\_Ϋ�֪j���ow��ʲV�f^d:��7n�[�A���#|z2�0��}��39?/����,��9>i`I$�����$������2(	?���Bƅ0aC��ۡc� �@�B2��HB�	�� �"�� !H@B!!���	���J��#^&��X��	� �X f�&$!&`JI$�F  �I "I$�R# E� � -�P #  $D�@�	 �0�"ā b	1 1,X�@,A��R2 �A��� H��� �"F2H �A�� c,X� D�� ) � 	�@"� 2Db�� � � !I$B! #  1`2I$B2 �I"  !"@ B$ # !I$B$ #  $m%� �BD# FI#$�H"���?��އz�:�?� �$ �� ��|�?���?��������?��������_�O���ٿ�}�'��`I$���C����HHO��$�BH�̟�>�"��?��>���$�O��A����ِI~���������_��?cE��XBHH�	!H�   � I� � � 1$�F   � ��I�  I$�$@ H	$�2H� $�FH  � $� �`O�$�   �  H�$�� �  X 0�I@ R �$�d �  3�O��_��	B(E
d ���������?C��hl���뿐$�BI��t?���8C��������'��l7���$�BI�}@����?s|>0�I!$��I$���`~�'���?F II�?�3��I$��� Y��HP�]'	���B��B�w!�L�>���hI!$�������$�BI�x{����!���w���� �����x~��$�BI�����$�BI���������?x��P�G�����@��������I$$��?���hh����O��~����$�����͒HHJ���=�������a���
�2��S��P�� ���9�>�F��o!QO�R) ABUT"��*��B�$�	B�D%dm�4hR�$����fQ %��PR�JU"*�!)�$HQU&��R*�Q($����PF�B����[e}��(�a�IQ
v;jJ�5Jm�eQT��!M�uU%BE��UT�� �I(B)EE���T�HEQI=�E
������*�l҄
�HT����QQ�ȕI!�  ���B���kb���ݹ�ji����{���\�S��6��R��aL	$i]��֚����%�u]��������w%@���R��UT�Iu�   �0�((��B�
�E
=
(n+�Q!CCB�
9�w(P�������k���f5��;��ݺU;VF��(tk�;5��Ql��U��}ܺ���T�$�U�A   }�m�F�vu�giUCz�t�ǹ�V�l�l��:���1�ej���^��1��XM��:]���u(��mMڵv�a���ӭ.Ԥ�RJ%EU�)A>   Z�zwXwB0�iJ+7gm��w:L��ۅ)�e4�v�a[���Т��GZ�V����R�Z��*����P���R��R��������P �^��X4U>�����3U`�4�)H�2�V0�֮��r��A�%���(�T*�FT����QJ
�UT�A+�   �uU=j���1TSm��� (5�XT^�r�AAvΕ�!B���	Y��
�]���k��kEkJLTW����BB���   :��)rJ޺�QͤkTH]rp�j���k���M��hɊ(e`  v�8 jX ��RH)D(�B�H�    n=@( ����F  	�5  �` +ۀ 8  �  ��@iXP � 	EA)(������   vw�� �o�B���((ڀ  ث� Ұ 
�a0(j0  �� ��0� 2�!"!
=��R�0�  m��Ұ� р �( ��  	�`  j�� hlP�SA��@�`H ���R� 2 S�0���4  5SٓF��1��E?�� �S�R�� ɑ�L�"T�����=���������o������py���j�ެ�`������K,,-�}�������꯫�Ľ|��m�cm�1������6���m��l�!���6?����|��}���,�V	� ��c8���;5����aҰ^H��u��LPf=���RFH�7�S��K�Yݱ�R�U��3i�wM�M�VV
ob��ŻIQd���XE;�x�
j�����N�l-,� ���ƺ��JݵI�ͥ���i��
�� f������1
���#N�
�!{*���â����+,�"�h�D#��%�;��@cC�7f�����R+ʸ"�x���*l5��#�4���M�v�=��ڭ����
��(�WFE&����f٭2�i�����hm���J�dФ��כ���gD�%��a����pfFn��%5�B�+uؖڹ
�)U�K��%2�dհ�����46.�$���T��ly�����c5�;nS��<fm,�t�M2`X������ޱE+��(Lɪ�R�h�' ɩ��o~w-Ԡӓ�kKy�R�m9����q
�36�1�!LGX���i���k+��,�8�kV]�ҵu�W�HRK�fָ[�{Lr��83��oc��_XuK�b��r�Q�B�8���k{P=�̫�l^
�ޫd�(�1��91�r�d���`:]�����*ƶwyx�]�a����srmYJ��ORBb9z�ov*;F�e�ƒ�,MH`UJZk:��6��F�Q��!��v�X��F�kUb��vd&&�I�1�^�R��p�36c��nT��_��ܚE6�Mܓ�`�ԄՈ�1 ���!��&��[i+��!:�%�,2�ǷZʸ�y5��ԒI�s�c�@��� [Pݡ��2K��7Z[��.���7�l� W/m��!�w��˱n�߁�2�IU�'Sd�ϱ�����tc����p�I[���4��B:�͙��0M�ZN$5�`� j�ʕ�F�"��V��]��٘F�' ��-BWx�j�]��(�Kq���Õ�+ڻ��"�䩤�0�l���,���nD���4�h�uc*�Ҹ��Q��42�8#���{�4���AG\WYBK2B�8�8�)j4�@�5���Q��1f���!@��Sc�u-�#+NM8�Ab��8n�Q����<NRů�+�G*ՇRS�W�n�?d_��E�jz�ޜ���`9`ܼ�wh}��x�n��G�\�t��RcLd�m͋U�2("1L��+ݭ���[5���rP��  �U�����s���ȕ�w��;�
حn87u6�b����XT�쫢��o�%����a�t�j�k4D�1%�pi&+������*�n��Y���ю�%R�i��tfJ�vm�-�
f�TF�%�vvZ��[����� �6�U�5Цd��K"<a�m�%la�Y��;`�Y2�U��0
w7B�84`���:ô�8ZD������5
��f2�[Z`v�SXFj�5����0�ѫUCEKܙɂ�yp}t�IP� k�I�R�M+
f�PC0ثgD�Y�:X4f�e�Z��a���»�p#-�#v��A�E�&3X-X�U�;�	�i��h��'㛌�$�� I�g$̽�4e��4��%SV���L2�&;酘d�m62��r�ʰ�N˦��tضk����t(�n��H��^�Bu���RB�Ơ�.G>�,ݓnVZ������"ِR�
,���!�5���Z0�4��&�O1[R�[Zq\�(�'�e32L[�,�A̘,\�ꌱ1kY�(���T�t
�9j��ڇF�X0ep*ı
 �֭�H�N�w��)���YA@�m�б�ín�TSm��������-5��z�+���5�mŶ��Wj�U�h�A�õ��0���ƙ4���w-��FMŲzv�
7VV�l�Ѐ;�y	f[0*�˧�Ӎ Qst���)�m����`��O(06�:+o)X���i��L!��R�Kت�*bܲ�ݎD8U�º�n�F���Vm�d鹖͋���;N�9>�X�����J��&�El!
�'����*Yf���yb�jLB����s6�4�q=lY�VVӈ�5�	T��P�ɗD�v�j9VV'x �#��1e���MRCPY*���Q�)]M�m�Fa*{l�yOF�/Avǩ;�ʀ�;�t[��φ��ïV����2�1!�b!�pa;�KTUî�x��	U�V4���̺+.Z"��G ���C Z�ӻ��9Y��Ǒa ���A#�۔*֧&Jij�[l��.�V��Q�%��YC!R��-0R�3H���k$�m�v�s����DvR# f�-���+\VPe�x�j��EӡM�����{uwzƲ��.1�W� %e4�D�Gh�-�$�F�x�(���WD3gY��++&�
B���1�"��5qS��,�Iʂ��)#�F�1�paJ�#>���ut���1�X��j"��梘Ʈ��^��Հ�J-K����T8��"
��u����ZW�KR�+	&��P�����ͥ�ֻ�ov
�(�n��S�B0�/u�oZ�x�Sҕ���p�Mi�hX��
�5��snS*�֬5XM)[j�I��^m27f�y��q��nح�wZ�Ql��:��%�W6n��^U�=�d�u��)��lQ��1���;�blR���ݨ�;o`���+�Q�ұB�c���R1Z�nʫ3n��
Hl�cum'�_
�1�80a����b�Ȑ�Z�OŊB�Ƭk�w�GSv�7���[Єo^��K��\��Ly� &�Ѩ�x�%�[�L�.�g N]��������4��j�Zɫ��Z���TCp1��m��J�26l��-WZEL�)�zƫ�T�w�Ea�K����#)����)۬ú�Bėun��a�ۤ��Y�5��Ou�5xZWWJC���S0j�{�J'E*6,f�,���B���kvkTKY0���Ҕ�]L���7��v$�I�`'tZ�:^�p�-T�.ȗ�ݨ��@%!G\���0ƣ�MI�w��h�{�!V0��ܱY/U��B�;F���4��"}�04qTjqSgX1\X��w��5Kv�U�A���U6���t��7�c�n�+p� n}�͢.J�^�2Kr���J��1���N^�eJ**cm}h,�-�nb��e���:2ݱ2��//VE*��7Rmڊm-הq$�gI6�4�\	���/5��x�)zh���EY�#;�&h�|{���r�Yi��CL髼�k��"m�
!Ә�Z��wRݬ�M��(mI����Х��<е`�i��F�ǏC�K��[V���S���ثI��>dh̶�sN�Y��a'GsR
�J�`����,nc�!x [g(��F,��� .C����(��N�p�Z#V�^Rb:B�UZ���֗�2,���+t*)H'����8Ef4��a�eȚz��ecs��1�:Պ'��`�f��
V�5F�aϷ1Z���ku�]��d�^��l�T����vL_  �����f^1N\Dgȗ{V"E�y:/t�TSW+C�)����RnV�I�(]�x�<��4+��~�u�]'$�U��B˪����ye��BP-v2*X�V�5�����9ej��e�6�o�*���f��&]�A�@nޖ�Cj[cED�[Z.�{l�yO���";�yg+���:ʷ�vǰ���ؠN�^\x��ʗQc1Xneo�O^���:#�GA�D�!IZf�J���)ܫi2j����5�+n�JTe����S"�*[��F;xE"V;tZ$��q]J�h���F\��O��4��X:nX�
A�Ԛ��0�uRL��u��^��
O;��;Xr�9r�S���z7[�+Z�����;�F��C�%�WW
8���tѨיt�32P1�8�wN](���)�{���͑/�ԚyR(���.�vJWi	��fH3]��zn�#���!�[�q*�`�
Onee �5n�W�D+�� �M8�aki^։�f�РXUmp�)u��kB/O.�A���y����&ef^��L�:v&�z(AX$�^����[��!5�/(B`U	C���Y�-$6cQ����E#ϞC�E��V!��'
͒�Tt�Ÿ�:wKa�Q�T��1�I�ȽC����0R+�oM�`5h	�ލ�k^ѓ@V�.1�0=�b����d����7���~��ަ�ے�n���
�O�K݉�Wb�f,���
� 7k3A{��M֣7�4Xxvʫ�?��yu�X�M�4���ۺof�l���I��u�S�.���u&�cqĪ�8�[J�f��2n((����Cs5:)e�E�v���c,�J����@���Q��[$�[F��L��X0�����V�a(�a36`��P)X�^=X�u���VѺ����kMm�9Fa�v7I	��x�m���r�!sv�r����m����OZ[��l�H������e���k5	앺򂱔��t],���헗�2Z�����iktC"�-��^�YSn�ʬ�nh�ڎ=�I-��ݧq�I�*�EeVm�U,�72�7/.�f��(V4�R�d9{�hِm�)+.�`����nk��u�f�c�X���[o(iB�%��0-���k6U+��1]����إ��d�Z�
�S�Ш��J=w0:�t��a,Ҩ�j�t-��r���u���VU=y�� �;`�ݖe��" &M�uv�hЖM�fa4�S���M�C�EL�
�`+�^:o!�o��z�a��5�jǥ�O,Q�Ѳ<*�)b�P���X#�Jec�ysr�-I4���ӥ5���O�������X�b��dUm���yAv^�uoLt�F�Q)�2�$��0�z�Ye1���W�1�);֯A�D0�(�j\�Ď'���y
찟��!���]�h���2J,�nѽ���kb���Z�%�3iԖp&�R��c��jmER�&�rR�4�	ٖ���T�9�֠,U��׸�i�MTYZ��y� R0^V���9pǻu3J��A蕚M���u�!vټ1���pe+��[)���t��o*�u�fR��V��rcW�֫�wBƕ��9 fڕ�z``�U��b8�5�6C�0��Wv��wt��
�i5Q�t՜�SD�FlTBy�u}��KE˭:��-f��4 �%=j�G/t�i����ݹ��Z��@��,Q�m����r ~�7vT��z+j*yx��=(M��V*׋c�T��rTR�Sm��^��.Z�]A{Hˣ�ث��n����a h&n���
86VˈSs#Ȧ���IB�-�cqlRb��m��=�1�i��Vj��E+KVBE=c�ڄ�^�c�a�D*7�@�ն*�o �/[�[�-i6�W!f���A�V씋��0C.�=����Ff�؞�٥�wX��Q;�����̷K,����5$
xF%�4����քi�Sa4��9m�m��I��́^��چ���t3f�¸ld��rM0B0fj2�:��*1jbW���;K��sY��&�ri
���x"� �m1��:�b<7��|Mi�q .�؎�ZW�5��Ѧ�K�t+P!�Z���te�N9��u27xeJ؍1{��B���ࣇ�^��|rf��, �L��V��Wcpm�/
��K����b�֒T!�j�{��:���x1�r�9�m+6Pw�R)j�dT��Ydǖ��f�AicM�7L &���١'��é��Zln��KJ�mh��5lI��բ�Ȍ �i�b@�]	�Y8���q��GsU<���g�N:_m��nU�P+���6�1���I�`�i�}��N
ZJ��t<�n_LKP,6�RJ�p\)Y4�KQ+Z��\�b�QïB����P�a�Ƭ*uv2$U�Y��kn���J@\�����p�uh]f�-'d�ݗ�-���Up	)����ׅa���N�!*8�VLn��E���݀ʤ� jl���t$ 1�	mE �B�8�ƌҳlY��〙�^�`���e�y��t��M����.P��˼;B�]����۠F����X�)6�qfPBTd�y�v�
�b�t#�eb�%�Ze�
�ʛ%Ǚw/m����7��2���1�ͨwFK��-L�n5X�J̪!4�С%�kz�����23!D\��-�������u��1��(SVH�z�����փV�	��(�TW�2�L8�N���pm)s�Đ����b�ͩ���_-(��ff*
�n�4]��/WyNr=�cA'N��\�����aŌ*5��c׷E�$D�R*�7l��S>�,��@ֺc�۱�6ŨQ_Ɠ��sS�pL ]���2�rnI�b���36XgT�i��Tƌٻt%��ʗHJ��c�@bN�(��lL�(�u`ү)лM���k�wL-m�Zr�Ct�[u�R��ݝv�Qj�E�"�5pQ��+��A#1�NI&fQtF�TE.a�&��7y���"%���ն�Q�YZ���,��2��
�:���O\b���oNhQ���I����r
������ޅ��C(�6�Ti��N�-b)l�J��5%��1�6
�6]���)a��YVAIA�{�f�R�Xr)W��$�$�(�w@�!d��e$��nJ.�+͹.$F�ͷ�L8�oac8h�6�N�j�2i=��˗����0[�h2UG5�ٺU��Ƥ��q��ҎU�[tuL�zURCJ��*A���n��f %���{D�k�!��򔙔��7��r����me�%	���n��Ӛ+%�"%��d���y��壏pD�s�.�E�֞�YX&��஛��T�P��톳���=����yz5 ��6�d�Ϛ��;���Vm�V��7�K9.Vm	�³Oi����������C���r)�ɻ���2��u���{!!]Sn�f�������ѭ�n��#�]�M� 鍎�(WZ�'�k2��c8�J3tC��}w�PSKZ+ݞ�!ؾ�]�.�����!��U��W]�E-��f��S0v.Q�ۂ��	�*�<���K��pΫ�#�.�r�k�0.W܆��{ݙ�r.�F����c��\����΋=x"N�)n�+�i
T8&1���k7��H�a�]cE��̙.��3�L����;\3�F �d-n���M[�%�~�E�]T�t�*aS��n����B>��J��[��[��e���u{ȧ��Qul�d���nm9�>��u�N�``�<�K{kum�|�j5 �N�JVuK���@=U���.=��t2m^���L�[ɥ2�e��V��fi�ͤ�:�z�*�&�U�%�O,J]~�d�J7����
������~�����S\�V��)��k�QKD��ml���r0�\Е��\.^RRb�9&t:���}	�r�Q/:�T��<�D 7v�F3��[�r�`4,9�Wp>{�����Ȋ�1} ed
��C�L]�JHȋ�A�j��L�^WX�5 gVֈ����eeu��~JV)JX:�X�#�9�� :�nw-g�����>x�&��V�AS��t���+a����z#p�n6�����1){����M]f�)���՛��6B�,�4oP�u��w�.�'oJ��#��L<]]]6�ط��t��U���v�ي������q���3+,'Yn�w	���W:kqJ��kj�68XU���n�-Wf�_v̿�����.Y��\�-[*�u��u[��_�m�/z=#�>����V��Â���
a]�Q[��裦�"���w�b��n���(��Q�Ȃ�5��r������i��K���T���{y5͵]�CwWy6��1˜*G��T��;o���4��Ƣ�̝_6��,R���1��"k��y����E��f�q��]8L���bt�{��4Ш/�]�3���&�D�(ΫWh��՟�����j�j5̡@�8�1�Y��ڰg��f]�<4�\����z~0wf j��Pb��V�k�����(S͇�EbXŹ]���T��Ȯ=����U��\���˥����[���d<F�N�
�X�^	K_"]���oY6��V:J�c�֭��ef04)�+_гe9�`���|pm�|0�/�S�����aέۮ�^�ĳ{��w��鴶�K���-1��
�E���pP%Z����Gf����wU�~�2����B<�h�fbb�����`w�	W�;x��JB0��қ�M���kXCG3�,<�⳥�ʙm	�K.��Ά�F��IKwn���u�	Q4��j�[ڴ�Dw�VlCs����.�f�=m$M���6��Α*�C�E�3�߱+��=��6��u��1��H�4$J«���GY�%�]�]bv�m���)^N�:�����6��ю��'��]l�M|�e�9�'R#hJ�����pu�:bʼ�����$V��z��s"��x��
ŽX;UjT�K�2I����\�d�w�S��X�w�[{r��z )`Ow��h�UjTcB�gX7\k8�M�9��:}��LGَZ����5�м��e�U��>M��P��v? y���}m�Y���T{�y}tD���d��dc�(����3,휝[�*iΣ�sGJ�D������1!kc�kҳ�gpm.�����l�]��#��Mo�� ��у.����Y��v�.�N�W��}yX�g����2v��vw�~�BΛ��5���=��]sӫ�����@���v�Z�o�v^�kn�k� �a� ���g^��!ᦇmb�Π:�KL螪ɝ�AAýX�(̉�4�4_:Ǌ�u��mw�][�A?_Y��5��,:Xo�,lI��H�H�����0�Z�;t���Iܮph��{�u��.g�[H��R�|F-}�7�ó���[��������*�6�v�ۑ����
pɑE�hy;�-g���ͭ	\�9ES
��� �B����:���9�\�݋6`cyr�'V׀^Q�]��T%�>SDz��9�Ő&U����7�;����KB��N�^���*�<��on�ޫtޤi��T�{&�ɔ��듵�.�b��x`�# �f�t!D�[v�=C���hX�&+��%�:<�gv��+������v�-]Bl��R����A����*�LN�i����k�o 4�3I�)[�|�c+*ʘ3/MǙK��Wq���Y�&V*=f����jG�s]�Vr���ʳ�oNȥ�c8Ll�J����4�y��C��`[K��ΧY�6�]�`��c�lk^=��V-����)lH6s[��+���9�Ǽ�tþ�9���!�(�>�%�2fa�ua��gpi^o��:e��Z%<ͤV�5t��nQ��mm��씢��C����n�v��Wwîgl؇Kh��N��bj�V^ʻ*.W[�^Zo2Z�D�m��']���r#��y�(�_s�к.ѐ�/�tFvĥ�w�ZU�W6���Ĳ��`X�5�'qPZ�ҹ`Ɲ������y�C�-�ޫY�o�nb�(a�_Pw��Fw���;G٥3�8��;�8yU�7B%`����)�3#AR�]@���<��qW
Z	�|����AT�ꝛ��Л8Χ�ۚ!,U��gr�'ɂk�nM̉(�mӭ��p}���t���+i�3O�6�q.�y�yM�D(�`�'U&�b8d��e�˜� �z2�Q�ˬ��6�ry��.��0�WUʰ2,2]O���He���_���v7��1�#/��s\UيN|���`��o
[{�=�W���s�Pu�|�2ۛ�����FU�\�-сҪ��2��7��k0W��/!��B�����fE�w.�Wdu�Dv�ǵ��>��/���x�m:��;���B��`@QS#�M�TYi��R�c�f��cD21�V
 ���9u���]$z���z�$f�sk��Hc�̰���H�ڢ�)�r�m�kX��ث2f"�tC+�9�)�#�W�#>�]ђ��Z={��Cvr����ңuu�#�T��\Y�X�E.����󵂲�	b�kͨe��n��ê�a��g���3����R�ϟ|���t�4&m� !Yfة:�/���)���R�s��������-�wXn��YV3�h9P�#�6��<[�0�-�wb��}٠�ĥXG:ݺ��vƯ ��s�f��R����u��=J��R�8�I�ψ캓�G+�[��ә:��\�]3$��e���N�Y�r��%�P[|'n˻6���P�ð@�R�l�i�TV��z %���g;�cv�xbcE�ԫ��˱tN�86�����}��Š�L]٢^М�[ooY�����B�Z�\�~9�YI��Msq+ۛ�q��a%��nV�C/���-�D�d��0,&�ݧ���tRے֨(mp��&�a�R%� ��g�It:v����R�4 u��%<�@e�q�5 ����c����i���'Uǭ^ړ�[���H�G�ǚ�2��B�/�]G�U�t��)�qh�W�˙�sѮN�_����oƐ8*�9l��+h�א�����Y��:+4��+f?��K�V��Z��ZFW���wi��D�73:_���YJ�[`��%ʤU��x���M�OTâu0��Q b,�>�Ǌ�%'���u�E��1��R��t�3
64��sQ]��m��f��8��MKF<��zJ�ـ��o�n�'PX4)�d�y�A]	J�۝�c���'t����w�2Ԗ�+=��yZ�Ύծ�X8 {���Ѫ��΋56
j��s�%71��on��Vq� ���;h�і*�7B>�{O`�������moI�pŧ%�[�M�<��]4�	�klMc��Nv�u�io 0j]��9̬�S����j���ӎ�VsP�R!�BV1}��gK�}(B1��F��1�����Պ4뮅��u����l��F= ҟ,A���Um4��ć.�š#z%#Y��3�")�p�L�t�Ae������Ul�&��!**B�ؽ�o�v�*�_'_ �V�'�F���94��2�`�6+{�X�b���}u�co��P�J�Z�W	��Zl��wP�NeLf�sn�pTh� ��C(�Ũ�;��y�tw{9W:q^)�Poۚ_ٽ�L���K܇���I�(�+�ZAr(`kySC&LȂ�׎w��ٻN�䬰[y$�����Z��B��.Mo��2�윷�v[f��]�[�X��"���;��)��)�T+d��FI���M��[�����1�4^�FOZXoӮ}	�]�ylrn��/��ݫ<9�6�wa�n�w@�]г��ua�A�eF����ka\�hF�glf�T�G�e�i��fN�)��B�6����w�I�s/�T��O�֪UREfw��KX�K���u_ma�A'�}wf�wn��98�1��2\�z��L��������G�̏�Đʕ�fj��m�N�q��c�;jś��%:2���'3��+���ć>��Yʭ�h3�������VF@��l���2��@cd˩�(Zب�ݙ-�b�v����(���;�ƹ)�n� �H>�G��,aQ�,l֑*�e!�:����=�8�������:R3�������k-���{sbt�5|1�q��4j_�9LXo�l�� *����%q���k��;jRi��c�ri^�+�]8�oz���4�{��";|a��ʺ})��cCe)��v��ڛP��ӝ�y��.��^ɰS�/��8��J��.��^p�ʉܔ
�}��5�p���5c�R�T���qS�e�k�n�n�a����m�)��w�,�z�����ok��Ώ�D�0��W�7����u�I@sGf �<y�F�ז5�M���%��m�nW%2�upW,K�:�\Xw��4Wk��S�]�h\�W��i�6���v��jW�#�Y�ɮ����]�N�q�0q����muq$�7�W�u��[ie��#p.���z+f�����s�\ܜnf�PU�£��HE�K(�r�j�E>o!	=ڝ +�Q�O
��C@�W��z�*;�n����D����n_ �E��C8��β�n�j�M��z�և��#���Ube�\�=�����tFOD3�/eC|�}&��*�)�`v$^Ŭv��:O3�@fr���.^K�a�H��kt�}�-D*-Z�^�N7nLS���z�X�K���iw��V��U��w>�q���˺7j��"泣I*�(Ot��AC�}�����U�=Ohe��5�j<����oh��yw��dݤ�ʊ�+\�+���W�r��5��h��)nu��tg 8�Kp$�|&
.Am�t�t��J@�f+�G4wب��-��N��rh'���L�} ����XO�7i�M�/~�A�4���V�9��&3z�ܕ]�n�\MHn<�zW=}t��n�u"p��B����jDO\���R��Ót���ێŢp�R�h(����W�fK|���s2WD��#!$!ǣ6����f�3xL`k�p.��	��û�7n�"`\/B#Ţ����ЕZ;Bn��Ֆ�d�BE�mS�v���v��v�(��H0	�w�iu�*��V�Y�4U�"�0v�E^{M��I����R�p�����v�D��P�%�%Bt(L����7���}�ʂ�@��g	k/���/E�bnMem��ӣۂtHpg��Mv���eb�O���8v�;:p�/�ӢP}0I�,���:�0^���D��/�rܴ������܌����KW�9o;Q'����x��j���,Ĵ�#�4�e4g&�U��$2�3�������f��{�:���&ڮ�Z��0꿳!n�;��j���	�Ë�.�S��rq��_lu2�󘆺�8Y�,-j�vo��98��Z���X���j�$^�JoPWG;RD�K��M�r���S�;��,�+���_�Jr7V������S�W�C�5��w�℮7-����r�5�f*[�7*3����5�O��WX���]j��[��k�9!]����n�ض�]���k��Ȱ�E������h��˙�)G��̖dGcߗ-R�1�(Ef�Ψ�-�2W\LX�gc�9��.o���p׆�.=���͉��!�)�3�$��++mS�̳��*�O]��K���{����h���o�L�̡ö�쬜P�uiu	�.������*)�B����T�5��嶏FƁ�R�d��,��^`գ6�4r��tY���/��Nqa�f��aN���t$��z*�3�bB�Ƈ�F���t}���s�2�2�/RX�;(.��f6:��׷B�<U�B:���a�*k��B�H��y�RR��ݘ��t��k��a�]��M����1qӮܙ����'J�SH�Vr�qp������*��"�A��/5����0��0��L�y�Ihɪ$9�uˈ��}R�u��n4;��);2��e!�mR"���&�;�u�G��\:z�b��	�c��YԳ!�{���s�hVf��;�k�5��pǸ����D_U�ed�OW:����y��Ֆ��_�fꘛ�]å.���$]�ת��^-�s�#���<í��tv���N�5����"��Ӹ�!��v�ۻx�s��v�����.K2oq��l\�7�̾���
� �O(��$���[�_R����1������m�oGz����x������d��IUvT�j��q�R���z�O2�񡳸^�+΋&9A&\@��̸6_wY	T��Xt|� 7����SV�Q
ۂH;/]5�qq������5,=*Z�&�f�=�E-�ۆ��H@u�ә��P;uoq��q"�A�^̀DZi;��9e��;	C��%jq7{��D��^M�X�[.�e�yݵz��q���<n�\A�o���	{EŁ�өιr��U��okl������r󨝗�X�N�"�5��&�
Ц�et9uɍ�Iz��ǽ�*)�v=9d��α��OLit���Sh�\�U���]H��R��:��مe�@���`H��h4��\����4gR�p�o�]G	��Da��%PD�n���S���0��^Mk6�7�d���LA�&��K!9[�{��w@�R�hǴ;���Ph��P8���:⩹�k"�=BI��Q�t���lN��kq�j�����8먫���TN��EnR�Iue�F�����6R��chD*���q��5(8A�Kp�C5� �Z]��Z	!W�����Q9�U�.�n/P4��w`�]�N�@�ևbU���&Ҵq���y��5��sHf�u�y��XSK5Wԩ��w4���}������Y<�^S�[�w&<lx��]c�����������t+{�[����;�Z�/x"��Wg �ɹ�.+]�`JF]�)�����2��Uyْ�[�����n�$P6j�*^;���sw�M��T,t[�W��j�Ư ���r���n�q��أ*i��l��4�%��C��cظF1b���K��s����Y�Z�\�aW:ֺ��͚�#��[۝;	��U�y�F1`���%�+,�o\���"�_f�" ��c0�f:in��s���Gy�c/�cG��`�\9
R�K��r��P`�4v�q��ܔot	�'GXw��_E�w�X�E�ؒ'E�"ࡕ�n2������w*���.�@�*^�9u�R[�J��.��×XN�]�
�>�R6�'�a\�|hرM�k�n����L��%�
�F"��6�l�&,��6�<�n����t�V@�1rN̖$���F#�{ð��M�i�Q�/2�c�#5
-8eI��s���j�Zi���ҍѮ��q���lN<�Sx�YX�u�C�nX��8os�E��r("05�[C�S�Y��uj�NWL�<��ZAx,2�U�&�]rA^u�N%�"=�Հ�㍼@8�u���nN���j��9ksv9��jƾǅMȩ)�P���W-|�Q˸"����N��t/)P\�A
����u�4֚�9κݧe:���(��,�dvȘ�o��pᵈ�b�ȹƖ��ݺT�������]:��$��%�Yo�%��2@pv�:�4ؙ �#�_d}غV��fo.O��_}5�+M'[�f��J�C����L,��O[`03z�����ա�d �9kY�R]�!�����Lg=��9���.b�I��X��9𤫚����\�M�#����+�:/H
=�SƮ�bܝT�7/�#���S��Y�'h�%��{ss���6���M�]:Cs��b����ٙ԰���}�)����O8J|��:��yWX6��b�h�r��p7X�r-�q�ȑ% �AW�g'L=���a� �V�8�G���ت��0�V����\�m.1%�n�U���|2�蹃�Y��b���(��0���\m�{\��y)�Nd�ɛ���d�yhP��,ir���^�'R�d;\��z&S8�:�zH�]:�cB�S�)pia؀�a�vE���T
� ��v�p�����iMr��Noz�9�1����RX�@�5d�Z�9�Q�e�=��X�;���ʓ��7�r�����F�4�
�֜e{e���@ވa�<6��<��v�lb�,�;��2�u���]I�pzF��N���xV�f���QQ��ڵ��ȅ�}Y�vs蠬
����r�)�L�=�Rr�m��@��Ί���Pܮ�y��ee��dY\��1��Y�˴��U��j�h�"V�L�Z:v,J����Q�ٵ�)�t�!�Ɋ痝����L�IA'w�A�D�]�{��R�����<��{(r;n�&��beAyW�{f���eNC2���~eiQ���s���
Z�ꮋ�Ǯ�a����901=Ӻ]��&��j����!듶[W
�\���#n�j:�.�+��XԲ[,k���q�<�&:?m���w7�>Bi���e:���X���yJ7�S]���ö�8��1҇ ���\�0U����\����v�
�5�4Y�Z	Bx�t�I�pٗ}}�}��i5*3/'s�Mun�[Sj�
���.+�;��Vc�{[��G�S��7��6�kTzȲf���w;Ou��-���t6O[]`gm����<�}�ܖN�t�(�&��5[�3�uu��;�0�K�M��Zɡ$GY���΅8�j��!H_iYI�-���J�UwD�2�����j\;��O�I:\9ڕ{�Yi(١v�fB����0�nD\u�j��s�'q|�p�]8�|ug&w%�M\�{�!��/nwb�1�]2�tnG �hk���:gJq4F��C�����X��y��ڀ[�b�]Z���ݐ��Wfh��{&��vN/y	����7/�7����핻 �zu
b���Cj�ܓ�O<�>E�]��(K�wt#�[n&3(�ř�N�ke_/oN��oJΥ�1������q�ﷷ���+�o-��ZÑR�>�it�R��֪��@�t�+�ަ�(�lݳct��$J�"Y�r��ds�̤i�\��tH�������y�ɤx���
����gM�y!�K��É��b�����3�����<���i�ۭ�v����M�n<pD�����F�����'.��Jˊ��}x-m��w�ut��R�:�b��N{�b.����҂w��u���+���+�Q�����-Y|u��J!���m��:��"�޵V��^�	Gm	+j�����b&3Uq��q�2T�!p�]|�Γ��}xuVk�]B(��ӱ^X3յ^S����<1*ө�P�ܵi!])��h������{ua36���p�S\cPKTA賀�}m���tK��:��غ�Vُ["uIZ�ҹ���,Ip./���	{o����Uϰ��9�������0ĕ ���[-Vŵ���cm�9�+�^��[�����F����#@Ь��㝝�Q�N�jHį{4s}��K�ҷݑ��nXZKk�e:@ ����u��3Yg{i��VGM���v�]9	Z��r�N.��f�Fˮ֘��#.��'7�d�����3�t�%oL��*W:�{n����"�t'�-²u��m6+7��ݭ�'h���+���}Ɖ�]�ISC��k�@�}�Sy��t7T���6��f
�86.K�ƴ�9���M��=����J��OD0��>u��t���H!𫗛�FNn�-U��:�j���5�l+�w-���3" g-����\�E�=멂�tX�hmuu5-]�Z��KB�t�9�ʘI�B���3����nrE�:�r� �WR�IXB����:-���"f%��6��v�\�"Z��+�׋ޕ�q�u0]�����ӎl�7���}K�Wٰќa���;E�f��`HghW�v�"_]%:fu��p)�G׫����2r���Y��4��|6!����<��>�ȼ���	�M���z��`�M�i��
��	ZXmPaӳco���b��H�����K/ #�r�k���t�]6+yp����٣p�8�?�N3]�p�3���|�.��`ǽW�l��on�QX�1��-��em��Yh�d7+L�<�N4����6{'C�7���[z��j�4;Uu��c3:����X�Qc5:gt���u�O�Y�;�]e7v��Nﲛ<ļ�P��$�F�tBE�V���p<I�M�Y�L&%Z���v�_G�/��P��Sn��EL9��ɇ,9|�;A�<�k�/۴U�9�ʻ\�4��@C0���:�
�&T����|�x`l��KF��\I*6؅h�x���@����0�3[�ȬIm��ƻxDo6Y*����%�s6`&n���-����so��i��Kt�,���a�;(ҧ�/��.���c��/�,=���:T��+tH�)]�c�F`�|�_0l7��L��>�u�{�6w�<��f8�u�wo�(����@���u�=����4�Es{x��8��J�3=r��^#�&���;Wv���74�b��e���9��ړ0d�,rݚU� w
Ū�6�
E��²�;6�,��UVL�9k��1F����dd�݋zt�Lu"�|���v�J��8��3�)K8�$Zenh�lgR�Y��U��a4y?���.0�7���{�"�u��G�����Q�n���T���RY�\�+�+�j����{'U�r�������YA�5���s��Mj��e�d�wosV���o���H�:����m�`7��e�ũD�s���j]_"�*	�v�G��8�R�fsB�:�T8^1cND� �լ$�L,����A�9N�����*�n�G:�Sg23Ô��a����1R���γ5_�M����^ o� ZΠwbt�KD����!���x�Ҧ_VJ����,iZ{��ԁ�ZmꚆ� 0�|����-�ZA��f�n��<�ft��K^>���sz�zڀ��K�g^I�=����(���V����H��!��E�n�J���U�烮���'�" ��"{��/�Y�˅�*���m��"d6VD*f�wR�f�wu�[%�:�v�sųp�ĩ�[bs��c��3^�c�z����(N�f�i��g^�m�+q�Δ��x��q�j�.o��Ht����E�C�5�!7�S9L�wG[�Q��(�c
���]�ݺ@���4,�����fkf�]�r������"��:�I���-�zi@�^�E��u�	5�L�l`����+:�0�`�
�,r�0�b��"��{���fN���9�:�L=��yݣ����"d����-��6E�f�TP�M�I��>ё�["���ua�PP��qǒ"�v��r�3��B�n��x��i�I\�Э�B���Rr��mVeZ�+�#ţyc��"S5���y�$�*� �� uOf���0~pV@�L��Cu��Q�a�Kg�*�3Z	\���Թ\e޷}]��Jݡ)�K�ob�j�;&�=�n^�Y ��͵��Fe����@�:�g������ɕ��<�����V�[3*�	;V���'a��1e*;I�4jC)��'u�0o�r�SSOPe10@�����<�*��N��V涢���R
�rD+*�^�K���2�oUh�(�D�����b�WêfA��Z)kާ�x�����c�c�;��٧�BvV��6O�<s��AU�q4�)��F���k,����;g��5��6���z��a���e�����N6w�����6��]�HV�8oM�WV�7Ki��~&�=W��8)��cl<��V�)嬕4��O�1I,}�����%<)����/�Z���t¬�:�"�WAx�P_h�a����Myɨ%���-Q��T�VƭZ>�KD�Eu�'6�m-N�9pj��[��`���^��^��� ��*�K,�29"��z���\ǆf���vf^A�)v��3lH(� 2�u�U)ݼB�<�2�}�tO�lZ���%����\V���ѳ�di��uvIԺ���>�C�E��)ѦmgSY΃����Wv���S%}�U7N��f�pu����J�G�c���W��Q���z�y�N;hI����"�^,�(4<@J�lm&���}�_����
�u�W$�dT9�sڊ�wv���m��h��㮘�3e�V��q4w�Sb�T=�;\F]��ɓ#�������M6�m����#�ٗ�����ζ/�Ɏ����� �����{���H仔��d���|��^i�ޮ_Q���]�ʂ�E��ë�R�~�06�*ɕ�l�O-�S��'�C��z��3��Y��t*\��jb�F���2��Q;�Dw����m:o1+[�˗�Ãw��kT@�'i�`-�=�\�����Yn����Ng,Ww�,3�h}z�aE��=6�M��w/�Ǖ4������E�����A�>k޻a��I3��bi�o�>�u��uY�jH�gV�V9=��V_u�Ya9����U�t-۝��)��Ji�������1�K:�0Gۛ��*&ͨ��j�Z;�1)��Cj`mZ�V̋x�mXzZ�{i���s>�6jT�x�p�����06��a���i��%M��Cl�8bb�XF�!v��S��ЊGV��G)�]o2"�q\�Fa4����n�p�M�6�J�[�VL�*�$��#,�e`�\��ŋ886��%ſ_s��db�ʆ�,�i'S`j���Q/*-��e��jXt���%N3Pǔ�ee��b���h��y]QiR�Y���>Jn=�+E��7A\�6k�:�����:7���������諵U���r}���܊���ʶج�e:gJ��+#F�#1P퓺�V^-��P��-�WvA��t��R���k�_cx ��bT�������}V8��$b(b�g�@��r������o(˭��]��9��ɫ}lr��4�<�V��>�dʱn=�Z.�&%ǆڹ���w��Y����	yΞ���+]\[n�+���9�4�e��K;۫t�ms7�b�C�C ����ﾪ����U[�j5
�	�U��I�O;x�����Pf�,�oe]M�S��_V�V^�Ż=���
@�s�#�YKah"3U�ie�`\�����ԍt�im�޾�zݰ"��J�-"vT|�r-U�����[��+o�j�=�+��rb�R.�;U]ʼX�zE���rV���tԝV�C��m#�T�z&q����H�w9�ԭ
�VN����m1�9�KO#�K��U�֮�_J
p�Nح;Ϟ��m]vL���\���D�a���������N�L�M�iD�lҸS����Qz�5ik�u}O_��T�f\��@es'�A��L
vu�G���Jq�����s��gh�}f��4�Y1�O��n!����m��Cjq�ʦ����j��Ջ<
R����4��� �_R�/Q@V���n�)νwGc\u���
�B��"�%��2�A�=���:Ԓ�i�9u}�B��K�Y��Ƕ��|���؛�g�f���;�y�G|ѷ��2�e^S[[Z����{D4� ��+r�Ų:��>��Ф#-KrvS�63i*�WɳY7]޴�p�V�-�El�/��[��6,�}�gn'�&�;������D��i�q��1y*vo�V�����)0m�յD�9�|b�|-md�Z����nA���ew)�)Xw�i��]a'[�]B�o9V��
\ګV�Z�hjs}O�=��^����n�Yu�tĴˈ�DA��u��9�b�J��HQ�N{�)��!���StSd�r�.QZhE!J�蕘s6r,�I	2�)RT.S)R+	$$���s�k�C8��%��]MʶPUiI�Kt��Al�D�BF*,4J�aDjUD�e[Dm,��N�����K��36����d\��r�P�(Ј��waԮ�QEUQC��¤�"]܎z A�[�]Ӯ��j��ʨ��+�lt�j�=ܜ��bp�diH��j��AE�

閤K�\B%f-�������K9A9-���a�̰E�)E5EEB�gG2=T��H�I�R�h��Td����j�M(�ZT�ԓD��I���bfd�N�!���E(�r
겭R-�t�"+X���������>�=�{�ҩ�wfY����������>�t�0�pJ+�eo^v�k�K���kFԋ�}�[\�ve��]UGoR�����Dr]����3U}�/��x�;� �Z)��t��Tr����Yu����X5�q��ȸ����3�_]�6yb9X{��]ʰ:�KT4JڼQ�@��6�.I�0�:$�7�@�.]?��I+ܼN��\+!�\_vE~)��g�L\M��Ɋ�zi�Ի;g��kw>l�fb��O���ȇ�p�������m<�s#1��Λ{w�#�
��q�(�����G:ێ�I���[��{!�S�pp�Z%$��ǒ��N�Wgi��B���	�Q�@�Q{H
��䋊Om�h��z��_'�/A��N��W&��,@M�87t�=g:����S�!� _>��Φs�:��o7��\��PF��W__���U":n|���R������8ixo�g����
[���K]w%nK{��l/�P��ȡ�4�8�8$L�n�z���0��3+rg��Qk�� �|yݎ�N֌d�Xm9L�]���^��Y·��Z],@W�\��|�m�cd`d�3�7�d�%���t*������Ž��kp��VpzfP�fʜmnB�{r���й��H��}-as�.�&�;��J�3{w���e��ﯾ��R��SyP�����;�ˤ��	K\9>�j8�jj�|#s\YVm�wp1^�m��޿��q��8G��r��#V���B5ARt쁽�r��첎vY��͠���Љ�Ӝ��DJ�Z(_6����w!��ݵ^�1x���BG�����ߢ�	W�3�c"t����=�.8H�V�#�e*"܀���}�5J��Q[�*�&����2�@H��΍)��Y�Q܈F�a��+�uP�1��U�~�G-�7���`��ݘ �S�d:����b\8�(}K��Ǹ�
�[�>(�I�):�V�g��3O�f�s�$�������qZ]{� sʀ�ʮ�qG�#�������)�e�7S��gxw-GX,c2L,J�����OD��º$�5,�����f�t�	��,��(�:��m�^��b&�LLGl��Y,Xr�|ڡ&*���@��E>{�}��p��a<Ȟ���x������8��++�o����ܸ@��
f�I�0�u$Gd������˨`_ID�~�.Ӓ�:���}_^���3��Hц����(��3ӁKs�M�j��=�?�Ţ1�����T�6=�Q8=����j�%)ǺrIQ��n��Ȫbl+��-@ofHE�|*%gn�����ұ�l�K�g{L��Y]�ԉՌA�t�Uvh{۬.%�i�����c�C^�˗CY���&wl}eb<�a�׶�0���[:�X�G�(e����[8j�,ϕ�>���}k��*���L�[kl"h�1{ms��@2I|b��s���♱7�yDn���TI��.k
�ɝst>i���[5�R��o4I��ޯ��l���(X�5�O����A[��P�� o��uம�9��L*7��9���T�%�L��u�i��s��9�Ƨ��-=���8H��������F�s6m�T� K��|@�uL� ��Q2�����ܽ*jx!�"��F�ɪΖ�
�1o��$��9+���S s�����\<�9����gy݀����]�2���L ��U�M|J,�a#�6��A櫡��~�2g���w�&��)��&�6a�n�+x��+��D=䨎���
V�-G�B��+8VLc:���ҭ�Zi%ڋ���E[��F��8��ޣ�`��%��&�q;���#m��<�Vm{ʌ-�ŝ}�۔���v�f�I���[��p'3q�#����r~GI�G���xu?7ҽ���ͅQw׺��i���<X�W�#'L頣��
OK��rYC���WC#1�Ur�-��aP�#�����{<��խ)X�� _�|��O����� �p�����(�}Хŋ����:QΌ̱q��u'���
ʭ鵗��=m���
�ul�r�OM�ap�%xV�OT1m;�=1M�2��(�Kt�n��?>6���^N�g�	�������`{w�����p��7��r�ذ���1PJ�f�3��
�^�zcD��L�%�lSU
��+U�;v��Y�G�	]TN}�G/	�2�XXH�+>��vrvwJ镎r;܈ތ�{-0��ܺC��?�+.55��u�(��6�~n��h�b�@c�T�!�4#�fS�9Q�.K�藵�x��P2)�7��+��ت�w6���=�QUC�8(�hn]H��K5c���VhH4'�E�i�/왎��s�������3�s�n�����F;.L`Orde��X�Ǎ�xH���\jQb��v#&~��q��U--�n��;�+�����k-7��ߔ�����h��믂{���Nʡ�K�Wݥ��2R�m��{�7ɕH�P���>%y͜/��+' �+ �(� �:���ʘ:}�8�D�F
��C�9&���S����F�u��m�w�&��mo,���5��K�ׂ�X�˺��w���^V�-��R�[cx�g��4�~ٵ�U�ʦ�J��uh����,H����1�X�S�����zeY��r]����#0�3���k;7"X���-.��&�������c�O�y�nJ* �A�z]H¥�9�e�N-T�=��X[���0`�熉�N�1�s�\�F��S(B�f��C �H�?!I��{{�e�[��טh��\wA�-l��=W�Ә�x_��qS���5�TFR�Lr�D��r�c�2�O?f�cA����9 �Z��2�R"5�����hEe��ހ�*�>˷�K��IF�<��� ]A���^�{Mϒ���>׌��^�����rb�\7�l���ka|\�����P��,X���ȴ��3�QyDu��8E|�ƅM��CKۼ�l�@�"9�޳f�H��~χ2I_w��ܺ+�`8k���Q_����U��:z����w�`�2������\G9��W�TT�on��yG�8@d��2JF�>��2�ҷ�mν1���e
_c���`O�����9Q�#Κi�0���gC�ؓ��n�3�.�A=K�pp�	B²��
u���<)9"��B�Z6��_��l�,T�V���}:2�T�/w�ӻ9Mn<�
As=�:��J_&v__7�
�8���ڟ��V,A���c��>�6���>
��wϫ����7�in��9�e�ہ���m����tGWK�un�M��LQ�:V,Y���5!vmv��JA�n��>��꿛��6+���ea�t�և��>&�Q��y��d��/��k�P�n��׾�oF��оz�ixY����������p9�*�a�T�A�tM��S����XlW\^�o͍�ηf��h�o/��O��T�J�'�xg��ϴ �GVf����-��҃�l�W����M���Zit�^t� ZL�e���m5�5<��n�����ʩ�;�2����;�ۗ��U���خ�G��#e��
ԅ^��r�\���2C�cÑX����8(8�m��tv��#7n�]�����ڗ��m3����da}����\�ɂ���A|pwqnRˎ��<�RmU#&�[ܾ�]{�EM�?�R��:f�`!�ڃ��2�v{�H�o�~ba��Ha��VR�Z�(=e��hu��$pƣ֬7"�P���q�,§�`kwQ�]{|xn�HJ�]��M����c���\��Y@u�y`T[��]�⏅9�Gn�%�^H�'��Vc�)ߨ�KRC��@G��Y|�d�_{ъ�����d��ә
~�yfn�|`�3�'P�5�X���
�Ea�#};>��P�j���e,����5�E'Q�bc���ᡟ&�� �Jם�]v �uck��Y��j�39^r(�C�����=��c��_W-9�`ѱ�~q�)\u��"b�%L�ŷ?>'T�����%Y�Ǝ�Y�/x����Э��qx�*0+,l�b��(;�Ud�p�1Pڡ&)����WD@�%b�{|�^N� �\I�:v~��0��zk\�3s�r���%�9�$+c[NW����{�}Qm�e������V�:ǵ��o�e+W�ԙ�	D�10A�.y��d�6
@(�Kݨ8i��"��0SYGL\��8P�Z�CK=��	#�g{ue�t	��Cru�*��$> ��p�����CZkӂ4T%�F���rpG�5�j�5ڌ���2�u�79S�q��~���l���\b�an��_>�<nX��_J�F^?W���fq�v�5�z��5����
�Kg�mSGu��'�^7�Y�Ȃ"V�݉�ך�yx�2,}8n]<SY�P֍yrR��8i>e���ŷ,n�sG��*vm.Ps��Z2��ǐ�fS��}A�r>K ��Sq��GOc�o�|�b��M�IK^�Ã�]�t�0�hSJIx}��,��"��{�V�@౳�1�2�q~��s}Hz��!`�hK�}�g�.5g��k1�UyG�ew;HP���*��f<��~�;�WJ�L�ݮ麨��K'�N��s�c.�}����oY8gK���|��|�^_Y�q[G:5������c<����E���w�;I ���q8*��ȿ����	l��W1 "���ϲ4��$C�i�ݑ���ήF��wft�C1�8sr0��ydTZ�R@�c��1�$B �B��z	ݺ�$��j�!��j}��ĞP�����r�gY�����5k7�8���:g���Q^~�i\�1���t����܎4��T~�I:�s���$ŀ�X�2`�;��v�N�����FPz����^Ӓ�u�-����5��9����_r�L_Ȫ0ĩ��ЎOd6n���8�q�i�۱"ƈ �$���3ٻP���|xF�;�eBf��cm���ӽ��n1\=���QdY����@죆ׄ�s,,7&���us���%6����F)���]��3:�'#��<jg_��n��p��_8e}9Ha�-��7X[���{���t�7�-L�R��p�5����Aϛ��ժ���:a����Χ(��A5O�W_I7������,��oK�W�~z(	~��1��i&�z9��2�W�%��ϢUݣ
�x����ӏFz�C{�ޓ�v��u�{}uָmA�]VZo�����B�S8���Gn��)YÚ��L1h�k��q�i�ުhċ���L,����n���_(�ZV0�7�&�Q�`W��d��Ϧ�sE#�>|��6k9M��R�;z���#U�>���hˢp�#�ܢQY�]>$o�1�������-Mk6���Ű4U�Vv��[u�~"�|'+dV���Eh�����y@s�M��׋9�8��v���y�U	�.�9~ctʿ.���������\�l~�S�8�,��Fm�޽k�����K���av̎6���#�N���,F�.xE�r뼨Wmwn6�>V
��}�8�� b=gK�b��	ꯧ�ƣ����#\�.�lDvͥkT�d�ZҠzɊb�5�t���:�	\c/�������E���f��E9�m>����}v�R%B���
�G�$�m���][F��n�G�"���wB�L���Fv�)��]��`���/�� �o�V����~Cj[#_��a�>dY���3f�cv���$Z%,-���˩�jX�sûƅ�)�9]o�j��5�c�e��J�����Cz�"S����6+b�T_kS��F�X)ܨ�S{P�{&�T���5w;b8�����bb�"�c�O[�YȍS�]�'����8�	���J0Y����V�]{��J(��$FVky8q��[:�#��;yEp��5�wf^������<K�}]:�c=O���:��Ϯ9�aꉜ;��<(�Q�W�̔RP���w����G ̳�YgEa�uz��X�n�]x^���]Oy4&��:cu�o��{��Ğl�@��5b�+u���p�AaYto��6P��I��i��hۑuϵv.c#�ǇT������7��*��b�����s�ypv}����ĝ0��VW!�.k���yw?������꼺M3�^?�H��'�8���u}'�E/��U���ü:��s�S�a8I[�F�a�ï���(h��+�i �%n�z�셫�n��B�����aq���VA(�-��r��4�U�e�b�D�K#�]9D#A�iL��}�s��n2XB+�R���)l��nwOB/J�u�Di�#KuS� ���^�gs�Z\ARl� CN�<�܅�DL+u���6��p{3 A�Wґ8L��0)I)6�7j���������T�P����5b��\.���l����"��Aj�}u�|�v��+�ݧ�$N]��JZZ{+N��{'=��l#�oq�|�e�-nDN[���;c�ʱ��:Y;Z|�76}t�X]f�b�C'.��C�8�ݒ�Nv���VZz)�j���74u�m�e��P�-E�]�������vf&��x&��T �N�!s�o*N�Uy+�o:�!e�;�1�@T��6�>v�x<��0�����#�m�\y�`ބ��t[��9GO`�R��ىf�X(��b�F����&V.sn�)!�:q�"x�5�v�e��p.���-<y4s�#Z.Ì�ت�BЙչ��	��헥Z��Yį�[r�Y����3ni�䩥d\���Ec�U�龠�%Z�1�8�����g3��v�M{VvC��nŁJ�@!i�;��pB٫k!]�������3��J�rܲ�h�}�Z*�rj�G��r��k��Nyu��E��e8��4��UN������Zʙt��H*�EiH�h�upĦ�?�{���3�pt���4��y��.:���r�K4jui ��V���|έ�ߏK*�<���u˾A��u$[�S6)��c�M]�f��x��oP̏+h�/&#Q�9\�8O������p��EQg:�B�cDΒ�<�t��ɶ"��f,x3.WEv��V���{�tf�9E�o�:C�6:�e���QQu�r0���}�M��Q�.�?lʑ@��o~0�����'y{9�G�gL��A�}�2qǫ�ʗ�#���Uou�*4(A�����-OX��}��v��!Bw��`.Mopەӄy�H�l<'�ۭ[���W�b��y�.�cFr<�)ܭu<}f�N��vD���j�E[aȔz��Zu���xěw�\1��m�y"�^�V��J�jא��T��.�G�Ԡ*�Bp��d��|��C�`�8^C�IխV�7������Pᜁ�dgLF�0!���t���O��nC.����P�n;�i]���v��ݎ���H|�+�e�]5��(�c#�j�U�O=3._G��,)�p�h��T{_dw���i؏^��ِ&+��Q��Td]�)��Ƞ%5R�u�O��P�5w�fm*҃b۫��7EW��R�oi�q�c��/l�L�ve=��d��Z�R��4�{p�֓bV_8�b{v���B������7��gr�cjiu��O*q��_`D�5l��i5[c��a�Xr�Ňc%��hv�kp)�JR����	��מ}�Fx�q�P���/)"�Ǜ�n!���yk�c������-]v�Xṓ�.7����}\�+�Y�C�!ݕ8I��1Y3A��b��"v��wKM�V�c3�"��yI�L�ɉ
�9�i	3Q��(�H���WY�vXa��뻲i_gi����Af�2�[2�]�PJfԓGf��:�2`M�����f�vH�x˻��"�*Z[�ǿg�c�ΙGT,�eHJҊ�5˝$�
�9�b�I,6�����&�3bWB
��]�L
�QIҳ�(�r��l.�TUVt�6Y'5L��E˝��#�I��t��H�3�q%f�D��(�	Zl��J�j����i�	$9E�%B���Zq*��B�+�(�.Y���E�%�*)6f�[g-BLP�$$�ZRI��'SJ�)mYʴ#�f
�EӖQ��R��2*E����u�b��Q;���jPFJ���P��:&,(�(ք�)�G#���u�uJ���!W-���.fkJ�� ��G"
�dd,�QT�Q��r�Sb���AU�F+Bt#����F��
�dJ�%:�w��a3�aA��EO�)�@��
9:,�]͕K�D���[�[��&7���d�D�zk��7��p��7��R�گ��{�w�ټ�Gg^̬��$�w�neEm������f���]�*��*]}WG�������0�z+dM���M��9�@Y��=����������w�='�?�?z7*�$����<L?�?P�|��j����'���>���>�DF��MuL�=�%;W�BC�|=���99S?��zBw�k��ן\���_~��^}�|EĒ]ʛ�?wB�7������>����㏮������|C���w�9�� }��>=��^�Ѹw3��ٷ�Ͽ�/�~{��=!�0����= ���7;{;�~'�ߨI��oϿ{�o�'NҾ�}��܄��_<�����<C����?��?��v�������q+�q������ߎ�����w����>�Ƕ�����">�"G�ϫ�xG��~[���\c�<M�	���� >�!���?�����=;N���_}�oI�'oG�r�M|���u�a~&���1�Q���"!" ���\�ex��l�N{e����>���G�='�#��p���o�<|C������x������睽traw�[��=}�Ϸx�_~��M��w;ߟ;oh!�=�=���99������C���r}����>�z����fs|n�z"$��"4G��",GпP�O����M '������<v��A�	��R߽�|B~�w�/W89���|ޜO��aw��;oC�ܩ�����zW����w��~{���!<�9!�d�qď�}�>�#���I㏮�NCߑ��P�w!���?x=&M�=ow�~'��_���<Aw��nC��S�ߨIψ{��o�N'����?P$�P����ޜz{��x�=���dэ�d�f�z?��"�����x�&���ߛN�\���;(y�~��ێC�����߉ߑ�aw��������U޽���&�BM�? �㏨r��{���hv�'���z8	��}���!H���"#Զ���S_����ޓ'�n���܁��z���[L��iǳ�����߯+���M�	�����<��!�4�'�~X������~A���n��x�?�|�>���8}}*vu{ D�>��~���!�����=��Nv��i���O�?]�}���
���O[��~�����+�SN߿>w�zC�O�~�w����Mu'�-�7����wڞg�{�e�;-.uiK�{�ٴe܆oHc�����h��mJK^Ҷs?D^��v��QΝ�<��K)Eݪb�5��p�K�H6y���U�ִ�{����^͑��/u�-.1Y��;TJ�u��܄$�c52*dw5���#� ����6Q�~ŧ�����Q�{C�~G�@}~�&����㷤��ܮ��o�x�S~|���zq�������!����7�s�{��w���=�Ͽ�P��]���r!��_��#�>���dЯH��=]�>��4�����P���m����c�{�m�ǿ������z;�����OZ���o��ϖ?�����n�>{폎?]���m鏥�d�cng���H�������NM�	(��������=z���;N���o��7&��׸C�5�c�{�!�0�������_ ���<K��㝾���z?>�P�>;<�?��������~{Zz9F��0G�"����f���1!�4�^�o>G��߯���&��w&�&7��=o%0�N<���N�q��~&���w�ߏ����aq�����~��0�V��~���&绡P�>� }�>#��t�P���S������BC�5���F=&���x��ߛz�c����:q�������;I!�ܯ��P�0���s���=�����9��~-������q9�}M�c��f��7���X>B�f �C�aC���כ뽡�>!�߿m���������)�o�$�{��ώ��x��=�������z�s����m��>����>$�OG�"����_�JϬӌ��S~K��m�N���=� F�B���w>��?|���>�����}O��0����?^M����w���$��I��������ߟ<ǴI��=�����4����?�_������Nק��j�t�ؚ��Jo3}�G���{���M�c��<E��;��g��v��O������Ϝ}Oo���߇�]�����x�Z���۾F����y�S>߿�oi��?��0��щ8����}��r�+�"4E�c�NO�@s�������&��{��#r�}_�q��ӿ�������?��+&�����|���|B}|���o^�w�}:q��(G�ۙ(y�3W훓���P^S�7����=x�������ԓӏ���o#x��?��~�>����;����~�Ʌ=���C�<C�~��9��A~��=c���>������X#�
�>����O�^�6�(��p~Oiĥ��`\��Y�>�;��7]��'GO���'^�������,U�P���v�NGi�唲NJ�\y7�N�f���l�� ��V�6rN%��̝j�25�&<���">��p��J�=>� `��#��1>���~��﾿=�HR;�m�.��>���o�r���|B����ϧ��'�?�<L.�}��|M��v�������nA��?��߿}�z�)xS�$�����"D{�ƍF�b����{~���w�aW~&��=�7�=��~�瘓����Io�w����~�{y����`��G�X��AF<��}2���]�Y�tz!
}���=�G�}�񏐡�Og������ޓ�7���>��O�s�8��߿|1����~��?P�0��߿�c�r�r���<��*��Y���ɧ�<��������nk�5�ws��J��>��#�Dh�}�=S�M�ޏw��v�_�}��������������;I!�����7�%@�|��&��S�8�~�r������ߩ�0���܇'��~�����axc.o�<��_����T���s�����Aw������$��x{����ɾ�>��8�_��~[�8�O��?��{C�i����ޟ��.�������������w����o�/���y���� �Y�Y��;�/}���㏻���=�����Sٿ/���o� ��,r�{I7������w�`�}8��;׸�ǎ�~&���x���]��������L/���������;�������qݎ�^fR#�Ab ����������������\
o�'��}��?�	�����;y�;z�[������s�aW'!��w�����t�'�9�{��Ǥ���}C�#<�.M�b�ֺw����'т#DF�
�����ğ�C�{���������C���H~&���~���|BC����'�p)�}�:v���=n�C�4�����<@���I?�|w�}�@�ezɨ�.��W���^{��'��?\}����ۂC�>''�-����0��|
>��>'�9��x*��?S��>}�ǌ�Aw�����ohRM�߼'?�ܛ�{��;J� O�~�"(}}r?R��dg4�y;����߿NC�i4���봋��Ow��P��|q�����܅�η���!�|���7����?����I�����~� ���N<ǯ��I�������
����
����R����8�����]�tɈ��bU˼���i��`�۬������L&W:#�ΔiR��X��p�m<LH��*=�@����KsF�0��w]�m�{ ��c����Q��+�;�[7��֜��8�4y�f �����<#DG�fH�1y���W�oVo&z�:�}�X��I���w���?czC�=�O����n7[|Ov����>~�&���|�����\
o�}����s��'���7�},�����|t��i���.�ͱ�<���}}��{����aWe����;�a~��2����;�=��)�aw󾧠����&��p~����s���?�q�������Đ���߽����7�'���z�N?�����|&W�N�-P��>���O�t�b#D|]8�~��<�L.�i=���]��*�X���9��{��3�C��޷���I�aw������zC�{��ʛ�?S�?��0�H-�޾?߯�]zo*�,����s�F�#����߿<�����nL�x9��W�����o�I O�����[I�M!��Sǝ�]!�YM����=^+�M��=��o:1!��C��o��9���y�Z+'~�=佰������>B>�">��~~�Woĝ��������q��?�����{q�������t�����{���Uދ�����}����9ۿ��q�u�đv�d_���!
v��7�S�ș����h�o�� }���?#���^F=o��^�M?���x!�#��>?���}s�1��Zz!���*���cE���{}�:��=4/������Y:/ƮϜV����)ұ�n�J����Z*�܎�dL?\��̂n�����lÌ���I�Q�U���l� C�
�:i9"�=� ,��6/ꋶ9��j�h"%{[���y��`[�#�=���/���U<�8iuH�����n�q���Z�l�.0ų�uޚ+�֋^��":n|�8�3��T������ԢS��mz��<n��m��ɻ��}Ĭ@�:�ce��2�=}�2r�R��a"c�˺W��ќw؏3biJ�}�m:�;K��,�;�0*"ūV�� pub�+@�GV�y�+I=���VoâGi��$Y�3Y�����
���~�u�'O���j]�,Cn~�:�nN�bD��r7�o���mG�͞��s����,�*Y�*p�}���.�g��.Lh�F��_ڪ=q��(�:�X7�K1;�ݭ4��K�&����,���w��-\)�9�5�;������r���gS�|��Y�g�9J��N�h�8�U�v�����Cc�m_��{N�04����j��f)���Ș8����6�}�>H������	��R�y�	>�j^XbN�7�6�/;�)Dn^����ܑ�
4t���3F!#1]4(���"	H�;e���8x���ayտhwq��a3�]����-Ԑ21sTp�}�q�g�޸��=V�,v�uU��6���rD$�}M�1q�"��J����*���I�ļ�;��������u'��z��~�]��Ŕ��q�7��1����p�͚�7�ld�F�(Q�l�N~�.u(�|H�������T`U\��agl��98O�x�U�j��"iЫ&��Zݦ՜q�>U%y��2�F�e6��ֳ� 'V�ק�T�T�W�[�:0Ф�uV�m�$�ҭ��K\�}��ʀ��f�h�5D1�\ߞ5�n��$�@�������ʾ�e�O/������3���F�ީ�ݝ���}��W/o{�A�vί��q�C�x�b=�'��uٮ���_�倧��� �S+�U��̞εs��J���㵁�����瞤pȗi��,u�b�߷�^��x<J���c�W�E�z�4lY�	��5�f8aߗ\5��A�܀���l�D�K3�k�ϭ�Å�/o��N�9�{�ʧ��-O x;^:�?;�򆰇t�'�C�V,�AY��I�NJ�eMR���i����1q�#]}�����eq�ct�j���G��Bz��*��u�9��K��T�K>�E�M��L�-ƴt�J����g�Դs�\L]M�
v�З�Dy�����+�ݮ�P��u�&o��	����k��t>}���^6��(fR=f�{�B���7e��W|!ρVc��	�_@T���]�5h�������s��=��ftb��8;���,u7�	'��B�% �W����$x��fB��f*�A��v�\b{kh�q���?l)u�r�#����n�ȶꠅ �L�gz� !�*{����<�p��;�mJ��Z���D��d���ۢ�q{���xz��}MKC$3���d�߱6�ڶ�!��]
$���gWt{��vwvR�ozZ�ig*�`����b�Io;�u��CV*V����꯫���qV�i����b��;Nf�f��W���8 �+��?R�R@Hls�e��f�O_�k/=�\�'�*�q�)��,��1����!�eS�PN�n}�R��Ί)ֆ��ԥw��ЯSZ��[R-T���[�A��A���3{�����~Iճ����t�F���8�p�H;^^U`l�Π��x-�i��G]��t�_[��Q�r����L�/��6��X�&84� � ��a6 	���L�p�7�}y���{7o��JU�T�ֲ�s;ձ��ʄ��}��k�>!ѱ��WV�a���%�l�F�L�2���mGl�ĴԬ��C�r�ӡ��=�7��fq%|ܔj����kB� �n�����W8���B�Y��\�\��y�^̫��*�p��§��W	a�{��kj�`��������G�_P�t׫1�1{)W�Q<(\d�1_F)��;T� ;�Zb������׺�aK�,�B�r�u�ZY�aw�A�*���xBo�}i}��cY���xVd&.5b����Y��;�l�)�ǻr�/�ܴ��Flm�}f��������F�RT^ݜ���5r�R[���*K[}:@�� 0խ�eΠ�7��=��mw`g����[�jm��J�,�)ʬVd6��O����`�B�;���m����_}_|�lk�{�j�;�c�y۰6�]}���wZ�#ùJ����κ7�I��7,z�V\S��u˧�j*'K�U����<�s�cB��B�U�����tV�ƎU:�om�cO-nء,�*��ơ'�-�~ct�9B+��P�ɤT !7I�{v2n^��{��\����{tuh�������uʐ�W��i�-�Xȥ�$<��f �[WLU-�J���l?��|`��U 9���)B�a\=W���cQ�m�qR�B�ˣp�\�X��F@X�j��$:�
r�a����`R��V��q�Pwݪ(\�p��yi�Fr�ҁ�b��V� �����f�ؙi�gԺ���7C�sI�<�IV��������֊�aX��\���pP�Sx,�����3�k�\�����aw��,��w���D0�!bW�'���FO�"���#)�=;�L�)�afĚ�X���w F����\�3Q���5҃��3��0�z��M�{w <��A�) �����A5ƸD��3lŭ��� �#.)�D�u������v���7 n�(��t�U-)�ܸ*veׇ���7�.�N
����n��l*�»2�ݍ����*�]h�i�(Ǽu�Bh�SQ8�[T8a]�r1GP�J�w��W���>��+�wV7vT O}&�ӣk�a�c��1N�x���7_�1Чj��5G��Im]e����:�t�X�`�m�Zخ6�R������. `�8������$dSD3G�MjKT%݂ݭp�/�pV�Oi�/���U�[���7�!!2�N�r�;uɂ�|�úQ7�q�炻������7>K��Hh�����+Y�1�-��{Cf��@)`���ܗF2�s��!��s�_n���������$Ē����:���������TO�~Jf�g�z�!S�q���@pxn:,�Z1��_j���N�&��׼D��[ N��eL��N�q����UHm:��/��#�[/IU�R��V�ŹK޻�~�S�����g2ꍠ3e6��	��=�]�hS�X4_�ڿ��`Љ�x���-�t����e6�-��`s3-*	P���1G�,
��y�����U�8��5��U�!�VRG�@��r
�Ȩn��Xf4D$r�hQ[Oy���!��a�v��Ȍ�W���c-�'�a�x3�+� �!@��Y�ĲU�
��lM31�D�be&�6X���Z���9���4�������J+P���b��Gǃ����y7v���$�g>MK���GN��"�}<�]Q=A�9s%�I+i_�>�����m��9gs���
���Ȣa2N���T[�"*zN�L��* �A�KrE��5෯�V��};�3�R;�BLW��0�\���\7�E��8�y�]���wgkcK�t�~�;����*!�|������F���J�Ɍ�~zj"T�E⋤)<즙1�#����̀|V09��
ю�u�-Վu�"�p�B����y�X�B�3Dp�z���ju��Q�%	1�[�n���D��{���
���:�� ��O6��t��&��p�y2V�p�:�s��W��K���3X���B�]�t����B��f�����/}��/%f�ᇵч8�(>���pԪ'�Y��2�L}3��ח�4;!��T��2Q���t�C���Cw�
�U��[ʍ	f�l|.����m��{̎e-����5�~�\.
�'��9���O0�����W�泚q�&�{���'��T�Z���|��Ã��_y]cZ�TPV2[?\6����.g��8B�Ŭ�.�]�9wSô�5m�u�qg.�!wY��sBd���M��D\�X$�K��\��"��ć\�f��)��F4�����:��YpM��
���g,�I��:'���o�����͋�  ��U7�M�
�. 0����w[��S��l�M��e��"�w�8�;�lTJ����d����)��oE�oKK�̫���\Z��O��v��	*��(h��u»CFI�X`}��mq-ѫW:��Xq�]wO��@S�5�{�&s����y��49�i�l���[�6�)\[\�N;�N��%X4��Դ{@�r���MQͲ�/9;[��q�f՛E
�2Z�N�f�\���H�
�Ww�eJ�0��ng+c�c�i�x5���|ꄡ[lQ���X�E�`��˜C��%�y��b���FS���vk�Y�d�aF��z���S���Ql�v;�S�Qҥv1#�V�g!������oU��_<]��ͣZq�̨-��X����ӏyV�	9��]&;j�Κ�y��/{��=*��N޾̎�be�J�V�/�ce��yz8T�=X9�;�l���;����RL��M�+��_1������wJ{�;��*���yϧ���v�dْ�2�r��^Me$N�Ю팫t;��;��k����w؃Ɂ�(�����K�W�dAV�N������	9S�G-+����`Vw+QC���(�,�T�6�&��cmLw�a�3���G��g��� M��%�z9���Κ���`����5^���Q�8u�z�:�[qE[ajR�
:-C�@�5��3��vd��u��yEs`B�Ù��M'�`
��&�5����J�B�U����	D����Mh����9Pzhmn�Wc�Vy��M�b�ݪa�;fV�̤�[m:���r)o�ث�a�l���t�.���STDRSp�y��^fӢ�6�59����<�fo'�3�&���p(��m+!of�M��]z�(��e-�f��i�w(��������ݭ�;�(��4��-u���څ��rA��]�E�M6D�Z�v��DV�t$�9��J��8�u�k�E]w�o��c]����΅;`L��d��kV���9�)3#��@��Tb��*�Ƀ��]ګ-)�s���0�]u��5n��o-���=Ø媣	�q����d��ILՙR��������mh*]��f�R��@�S�6T��j�f�mFsjI�kl(�t��|GW4D3w|D}�u�cn�[�1��V_G�ӗ4�WW�C���$d�De2uޏ���]�f�;�N�]LV7�j����.���x�.J��#��]2ފl��\�:���� �o�q5	wA\�:���-�Sx�扸4�uĳ�\-"�]oq5�_�蚈��;�� �K�Y
�)fJj�G���D�{-ʆ�EXݘ, ŒގU�ҫ�G���"�yTE�r�S(��d��V(��!\��PUNX�I��2��a�{u�+Գ5�R�:�TRTTFB��\��]a��|�vC�Es�e�E:�]�G5*�����y�(�3�Wȇ+���Yj��5dr���Be$%EI�Q"�Z"�RSηdE�w���\�
-͜����"��5�E���9Us�AR)ʤ��Q����Q�-eI��r"�
��D�)ʂ(�g�A2&Eqč0���
�PDZ��U*�T�2���$u��4�rs�U"���S�Aa9�;�
��Y)�TDUr�3*J�\�J9ȹ��Qp��E��W���|�NT�A+�"��;��9+�a�U$�G'"��]wU��ğ�!�Y)F4�wU���j��)`��էM�B�ᏅgI:,Ѽ)�G�_K��9)�u��&Jg4ip����B�9:��$6}_W�W�1�8���-�	���ڋ����.uU UMf�C[��F�:Q��<Gss��s�u)=Ζ�����e>1��J��!����RH�~PJU���R`�ki促�/�qj�5_��E(k�u^8�7u�:!��bo��*������D��溸Q!;k�wJ�f�,����F��O�ʝ�w���ne`KRU�n�� oZ�P�<|.��&�j��خ�bD�S���!��w�I���qVgJd3#�Cr0�ǖB��TGML��߹w&OtDU�эR�鬋��0_�\������G[��1eN35K�X��j�#ۇ��������A�^J�^�?��$N��d~ո8�pP�6�}��&e�d���;��ڻ���!t�1`:�� �a�+�����n��t+[��u�s{;9ob�^$��r0<׆��fD1PԀݖ�0P�P���L�p�7�}y����������n�a�Իľ��w�X8Fʴ�-�N��/�`���G\�+�1��c��"&x�k!�Y�M�.֤e�B���[�����Vǫw>֣R_5����i��hw����^-�������r�꒬/|p`�^R����s��8�J�Wv�w՘�AlwL�'�(`�K��O[���_d���WP���j�Z�O���꩛�S��6䂅��j�~X��'	���Xf�׳��\ ��qm}M=���U�T`�o��x^�M���bC��T�h̙�m���Δ\j�bG���u���{=�\���av��pÄ��q%�κU�*���-*�fs;|н���@q�܃��U:ے�|�) vч��d'����E��%#rb�mL�f�u*"W�Z_h���ed�Ӈ}�f�#0�q����s1C�co�W`���W���H��Q?�g�w].�˹յ�Ջh���#*�q�<�~�R���瑎ϝ�'���غ���d�@-�g�k�ٷw�d�L��,��D}��W�|��LP<k�\<�M��O�n��(EC�v�t�U�ܨcpg�=ܟ3;����Hn��Qr�
�A���#��<4Mo'��O��+�����rr��7=�{ҭ+�����$�_GϩPK���x���Ƽ�����_	��.|�1�od4��� g?��DR(���A\v�bc�E�&'�:%q��2��� ���a�J;뫁)�:����c6�r���2�[g1Ԝr�]�����K�We_F �ݡA����*[`��eY}p�	���o+*�C@�&��6�|*��)l�]�d��^=� !��g��b�s�1ܑ1��L��q��/��Z;�着�����G�~�ݞ����Xײ�X� UmdQfY�pJ㤀��%lȼ<�:�۪�3f�Ji���;�cDL4�1q�[8[�#��`���dU�D@�vT���-���>��X�� _QX�m!ZN��L:�DU�$/�X��7���\NV!��o���,�7����/nЫ�	�o�u��k��޾�������mґ�"h�u�z�����ټ�P.��0@
�I�00����T\��X3Q��Nፈ�[q�mp�KF�GS�<�����'6��Ѕ{��a��[�a�(XVo���
}��Fs��W�u $8/�����9ײ��?�,;��t�>��t��(n붏������rܮP���v�|��t��F-�U�9��1������gZh�������A��~U���0���s=I�����m���>7����Q��@!���7�TZ�����S�[qZ���wy��5������4�(�6ܦxg��c	��[��A�m~J�b����V�Nj�*e�{N������Θ�%�M�*w@��N^oe�����FZ���5m�2�P}�H�~�>��=�1'r��B����OcŦ1������lq:t�C���g,`At�#��A�M��.M9�"�J�ޥ����7?�������;����]B�q�ʴ�k���o�����rRw�_��Gc2��<vc�PS�@Aێ�4C{�TB omT�&8i,sS��������C!��*��m���z5�m=y�%՟=ؕ�q��ݼ�3���|��'`%3�c �"	���zpj�[ݻL�m�[�Zˍ�I��([ `��u2g�hN!�	W:-��E��"*R�F�"�V�J�V�7����2%qW�6^V��ހ"��QIS�g\�n�T=�s$|q��6�A��'�p�@<���,5	1_Tkj����5&�)�7���۽mDI��<w����v	K�&;V[��_$f�ؾb�gs���
h��J�������f��(�qI��Y�N�z���;<0�Kn�u�-Վu�"���i����>"rs-M��W@�S1;bὯ��M/��BV���y�HW����+Q.ȥç��QK����|��F�ʀ�^�u^�瞤pȗig� izo�$�;�
|�b�5��l��pڌ799��������8����X��/w`%�IF:B��]��x	�B}%̘z��˦���)Z��#z�F� i���ρ�}ut2�uh�,.�+���$2U�l��F*%Q�|$����ᷳȵ�I�x�S"�"�7M�g���着���lp��I@�_� �<+2x(. -�Z4��0����,'�h�D�M>�6@�V%�"h�J5۞&R��n6�ÿ�R��1�.�o��l�j������kO��t�x�{k�Y<���K�l��,V/k��5Y��^��A�_e��]�r�V�3�d�<���n�N��_.��-��u �� �\�^!7�[�h���x�x
Ux[�We��yI��a�'��@m=Us��|~�]Ѕ{N��|9��T����9�H��9k�Ӿ:��Á�̡��5�.1��§��()�JB�����~P/�J���,WF��Y��jV�b���rv�~���ۆ��AF8�7r5�)��c�IEt�8`h��W`��ј!��?;Ͻ}�C���hq�}��)u�r!�9��h�Sc[��9&h�f�T����zf����(Kzr��΂���8{�t��f�;�|��h�{�Y�-�K��50k�d���+2i�yL�)��`�,�뉟�L1�˞����'hs�T�.�^�ۧ�+�Lw�^U�֧V1�L���^H鵼�<2���;���옧L��9N���wS�'Eq�����2_i�Ƶ�7_cx,D�@ݭ/�Օv2�b�'rX���˓�;����s����p�IV��Ԑ��+<�x�����2��}��_}�f����� q/�,Fą.��[U�뺵G�!\�k�_/�����T�����kCp�٪.HnnLX�[LWs�����t4�����<u�.��֩��ɫm�ٜ#%��.�LB&o�� ��a6 	��'� ��49����Jò}����3ҏ������eBf�%��l9�d3F�a�\�.�0�lI8򭣃d�m���}{�Cp��k����6�fԥ�S_�z�����#Ʊ��I�yQ�z������w}Y��VѢ�+|.U�+]}��~�߲_]�K�z�s���cj��&���ﻊsXz ���LMf��܁�Hb/�!Tf�L0�� b�\��q���KbnH��/]�3�� �>1��tm��_�kl��%"DP�ș��}��Ts�f�㈾����N��gB�~JlGo:z^��2���j��:�tu��ɛU��v�߫����шx!��z���o�PB�jp�����y{'�wLh�Wւ7$Fj�'�G�R�;���$z][1��2���&ʉX���[gP�u-�5x�±���n�r��Xl6;NSSe��,������)l&j:F|w�9�Ĩz�������ŕt���A�o�Yg*�G��S����v��|s9ԙs_�W�UW��JI��^)1�i���5�K���ï�1@�}p�.[/fa�ӌ�東/�/0b�響��z��#��t(@ϮPhŭ�:�S�D�'i�
u�k6;ZF)��u�]��q�(C�n��8R*��Jo�PK��k�<s>��<��^74g����su���`����w[.t��ןDЈ2�p �v�C�Q �->�a)�b���53���Țf��5�Y�ßwZc�V>vP=�ހ�d*.X�_���2�_[n%{ԮV��n�(�d�!s�n���v�L�[9�8r6 ]�3ydZrD	�w[���+��0��l'u����Q}[&�J����Lh������ٸmP�uX>TI9p�5�v\M�ֹk��9ԛ%���X<5�-��+fj2P�3]҃��w~�`#�EJ?^��JØ�3<���:����l�
�hjr8}a�([�DVG���NᎽ�v��,T��W���)@�5�^s�ޟy��OU���R�Y\.����e�|������`ة�ڻ��-O���Q�j�t��J������'^W����=�NV���g�w&fiL�^�����yGa�� ���JeZۥ�pÐ*��Ӛ�O괱E�EMEP�7�A��'%'	��puo[����������oNUk�t;�˗s�20R�#��W��}U!����p8+�u�mp[�l��e�c�an�G�s���P؅|��9[9ͬ�U���ؚ�/����u�b.3�2m��wq;����E}_H���8�/z�`��fq�߷	�f]�_Y��QTD�&-s�����:b;����{�x�xK0D��m��gf)�0?������@��p�#&Q�;L{T�VJ/�)���6nf�A������'���f����x����@Q�rl�B�*�;����8�G�����X��톥0���7�0������b��G�È��iW%�;��t"�3v\�8|��c{',|�����,8��8������\1�8���2N�J꺌Q�K�������Kw�`��ʞ̊�3n
��$R�]�!���r
�:S"�n��Y����BC!�o��L�w���/�#� ��Uƾb��7q��3e�h+ LS�"�`��̱�����Й�I٥rLh�`��t|bzw`-�ӟ������b��E��Y@p]73%m֗;1W&���V��6ciV��J�mᮥW~�'��k�e)c@p}�XOe���.b}�]�,p+k�>�&��CqN���6���6+�F�ۛ�]�����Q��+�]�әo�JY<u\{菾������91��.�>���Br�N�_�>��b���[��T9B�|����ROSouEg���]�].���y��U���SV��P���W�z�W֬^G�~�1U΍���ff�ԞJG��GL6�b�����]��w�X:}�q!\iey�Ǧv�5��c�[x��_.��S7��yP�Y�LX�����#�D�NJX됝��U�1��=�(�)��b��0�;9������ZOCUM3zdU{���l���AAW�����ؘ�j+6����h�f�~Y�8~b�xmt�oO;d���C���MgdV��a���T��x�%\!˒���y��aW�:�.5HF+�:����6��+�m���ܕ�[�+Cl2��3:���e2�A[��(F�xpuQ+�+ƴq�Y}=�*��Z���u{:U�G�}.�:�='vb��(��p����Rb�x�l���E����WOCՓ�Z3+��X�x�V��nXۅW|�Ґ�h��u?(�����Eb/8�*j��31�cO��;�#"�&}]�ڲ��'�31�ԅ�#�;�wH����w
��p��9;�73q��Mm^�U)��ʓ�y��Px]�^Թ���ƥ���}-u���j�ɖ3��vӮ��5ǯT�������T�<��ꪯ��LE����2#�� �^�J��ojc�b�zw5�#�㺆,�U�]/tT�c�B�����]a-�����<�-�,m�k�̙�)u�r�#�����*�]��M��3�w �f��=G%��k�*<9�E/�`�;�v�f���(�x���N�4��3'hrotHG3.��o�'�8�w��I�c��>�/�!���8��בF��4�3J(��Âl{�����׽%�����#�vR��qrɉ�]Q"�������"⫛y���2�`�?X���T��D �@L>�zK�rR��g�o0�:�g�Ot�
� ���uq-��u3�zպ�o}g����WTb h�0�7&��[�o���y��)#��=K�Ӹͧ��ƈ3�eBf�̶�,����h�����p��·{(����ۋ5GSs̓��b����W5��Y��W��-=�*8��w#8����YYv^�}�ݡGu��eɲےL`�����He�g=z���oؠ�*�����n���[��Ak!��:���Wq!�6������!�Z:iw/f_.D�B�By�ps��x����L�:4ӽ�<�z,��~�;\ԯ*�9c-�'�Kv]Gv�����oX&}b��fdv��<�p!�z@i�"��9��������|�7SzVZ%7����5��NR�#U�f�"儖u�B,��tK��-^KR�c��|;tNߘ3w�y{4]��Fe��3��DŽu#�tVo,z�uI/nP��id�j�Ԑ]6�e70�+��.��}y}�k8՞G_4�5���U�	����[�݊wpoV3GJY��O�6�h��ɘ�^Ǖvu��.ܛ��t�@� &'�;-hC��6�Z�]mE��i	�K�/Veh��M�ڲ�r�M����m-�uÃǘ`E
}yYjI�nۭ��!�Ղ:�*�U(`�&R��l��ˋ��®���33y���9�@�r�1pXȦ.3�HV-h�ծ�gGIMrg�t{�s��V�d���;5�E����N�y���k��n�HR���-~=�c���OPU)-<�d������%=��r҂�+nLn�R�<<n�.v=�2���crAm�{ܣJn}� ��*�w�lW=D!���4�
w�H�Y&P�^ꕼ�f=@�ޜ�i$ ��P��uo{Vo6;��e.���)I���7��v��Fv���jpmNX p��ôN9�t�[�dotGJ{�'�ɂۚ��߸Y���xB��o����O�6���C�k8x|��ӖC�ingV=�H��4�v_HwS֔���:4v�a�m<�.��[OjdE�ɈQ�Χw�h�8�i���-j<k y �Ze��;��m���_��v���q��*�� ���v��5l�\�D��v�WΊWy���C�P`j��)˩o��o���eh{�5W5K;�;O0ryLFr�i�-""
��R���͟$��΢��[��z:tK]k���S���儨�<vQ�P�}�u���2M� z���&�Y}G("47u7vx[w�l�&����3,�:�F��)�9BU���)���h@�o�k�j�����g\�$ZU�����i�]Y�Ҳ(ѧ�B����W��2`��u��kf��Wn�H�M�vw�*��n`����ŭ�f��n�,���@�8��g��wF���u��Y-7����F�l���ؓ�½
;@�֍{��X7e�a0�J}
�&oa��_|�z��\����J���fmf��U��J'ᰃF�ڵˠP�7��[⁨㷴�Z �6�J�� L�7�b�/g�-�n���/4���G)KvAuV�oݠPffi[N�h\�?��u��gC�Ҩ�1f�D��/�v.�P� o,Jr(EYq�[C�D�	W��*�S��_ P$�"��;��JVӡ�DQ�Dr��p�.b��r�/D��������x�J���9A@�U\ ���e\�U"+V�����I���2"�Ӭ�v���Ԃ$����̊��]"5�(��wR좋D��CD�<ꉩwTD��Ǽ��W9�*EE�
��!\�3ѕ�F��G5#4��B�s3:�t��sL2�%B8r�*�2���k3*���j���FQ��NȢ�.�d<IQ��ts�򻨅�"42k�TUJ�]����e:%¹�TUEEG��DB�l3,�d�UUQ|�y
�r
�"��VN����:��Q�8j&]��@��r�Iԣ4�|qs�YĢ��\Չ�)�R(�(����=B+�)u½B(�U:�U�:��Rl�]���^|	�q���pTZ�L��M��N�����n�X�R���yo�+Fe��y���t{��]J�puŹ���W�#��#*^��0R����7�}}u.��xk�@�9�>{>U�(��&a��R&�Nm�KB:�U�/9��tg{�7L@�3
�n���m�c,�|в6�byQ�P���9Tp^u�HOuڑ�k���͓�9��m�����B����U��-�óbg�IA)�U�(3w	vM�÷�[H}nc�A!�W�Q���˯��Ƚ8�S1�R���-LZ.��
��}��}���vת�p�#��UE}g�V�(4�뇐���F���7�P���pg3�VUJ�����t����\ !d�wB�� Te��WXpk�-�_q�Or�o4�od5N�dR Q�\l�`�P�L�9(`.�����R��yv,�F<nk�M� ���v�i�ޜ����\:�y���qz}������c�n$3�Zꨛّ�*�i�[��1�u��RP|dF���X������Y� Ƕd�R���q��t���w{:2�X1um�L!��a����h����>��|x@���B'y@��ȚT�/�fv�V�I:��y�z�X�6Y�)�V}����Xۗ��ݭ�}ܧ)}��W@��󊫼� ��ݙ�e�k��.�Y�# �ڄ=m� �0��Lv�� ������8�[���zn�w]�3�do5#]�6�G����zU��ޭ;Ζ�
�t�2�S@g_s�YG�p�Sx�пUW�UW�OLa��ȧ�E���W�yDu}j�MF���H��J����N͛} 6n$�8#�����J0��5wH$:��V��e���l\�3�3;�t��<����Ff�䦉]�+�yK8$�i��� ~� ��A��W�>�3���qx�������TЊ|�a��u��o[U.����ٶ���
\�#�K[X��������or;6@{�NꇽV��q�H
(SrE�	�!ڭo����\�������<��[�}�ƻl��dS��K����#r����wR��tɸF-��yZ!;��+��ʢ.U�gf���k]懚i�Cs���WTY�f���ĕF2�s��L0��ه~�(h�a�����vaR36_:iP4W�	����Rb��,%c����Ubt���r�H�l����VL�˫�a�zyN5�ʯ��@-.� !�L�&*w���'��fC֝��TK�O��1�eVoaz�P+,茄sN_�9���0W
�]K�g��<�*��Y�V��ծW*�v�f���M6���
�\��n�'�B��~Ř���%m#֩�N��� ��� ���|�ͷ�#/N��n|��S}.[�\�}�i𶖃S�C��ppj'u��W����f��JK��������L*�/�W�W��f�8��w�Dz�)
ͼ���f ����Y�W�}@�L%��b���ﺜ���0���	�
��~�4&�#PH�T븷���d��L�n��Y �
a}$Z}^m���ݚ���x���+iaωh�����6�EwΪ!��uW� )?k"���Y��^*ޥ{�}�:k�7��R�P\~@8�bFyn��V������b�.q'��cq�e�XB��_r�;��ߪDnϷ(\et9>Q�Sȏ:5�~U���+�J�ɫ���Io�,��Sw��m.�j�Ux���=�`>R^��v(����b���#\,S�5�<�����u#�vlԔ6�+��LT5�󿂺 ���?`�y��HWZ���qO�7�ηl�f�����f���&#�Pb�9��r�1�P�M`���:kbeqљ��OM��j�����O���YJ�
gg6����㓨a���i��!�������NWt�泦��f*�;F�Z�r��LU/���j�vɸ-����ǧ
�\����:]@�s���dV���%-�cQ��73��΁S+rHZ�Mn�q�{����`�V�m̟,lEP�皘f������Ky��:ﬓX�Vk���ց�'�:�͜����lP���۾(z�[����}_}U�n8�����v������[#0ڵ`���8�����R��~���531����ĹW'@uʒ(��.ƚU�=�:o�+t���pQW�M���5����ǸTm���ith�gQ��5Mה��	꫕�d>?K�Z>��V� �k4�>�Π�zo�歔K�VZ�ݠ��[�K䡳�9�BDN����ìf����Z��ZhV2])oW�{~=Oq����L���+{p��E�!q�%�܍v�n��RQQ�')�4�u�IA�FK�;%��a����Cg���\^�낍DIWɔ�dH�q6�	�$l�\�)�z��}z��tV����T�<�����7v�f��wft�Rr!��0_��w�G���۲0��{,��UJH�֌*U�q�/�x@<v�5��M�q�s;���T�<z��w.f{�b:CwpP.H�+������&2�THY��>�!%��������={t�i'V�|Z��䘰DP�1<�L�9u�+�a�!&4�9W�-�R�ѪΩVi�k�
VbU�H��)�I^�\�%�5����DϢy���Ax����m�®e�0���ޥ��m���F�m�
M�[ɢ�闽LN즕R��5*���Nކ'o�a�[��L�Wh�����8k��z��)i�G[�.���RN�u����������gz��ݭG��sS��c*Ǝ�T7��h<�8h��wS�oU�h�Ows�Ԣ̴���q��T���;�90��K2���TY�F�o.���U��Z������y��.2�X�#?_�����#_�u?;�k)��)K:�8����oK�;�����s)���p����f���s��9�(1�ڷ��Zb��^����z��^2#��ʔ�[����2m�"��mb��;�銆��rX���a��vxJ���ES�B�8 ٸ}��׮^��תi�ڗ�.�n��[j!�T��F����1�{0 ڝ�L�w췾��.��{���W�F�)s��!�C]Kʮ��m��l��C�%=��gj5���%����e������@etFUG3O.��J��������P�c�!����X��`_[�]�7��&�C�y�H�4�뇈�l柘�4�Begf��1B�Z�{�V��@��6?FQ�<=Ʒ��F�сf:�_
m�牢��)�X��aa,8w��9�����:r�i���k��Q��QQhX�v�V#�R̗���{l�ӝ�ܭ�(���i�f�����,���l���s��#�w2<��Kދ����t��+�������]�R�M�.���#S1�:,�}�W�}Y�F�Z�Ҡ�1��u��b0PB93�䡈) ��%7ԫ�˱b�x�����9�0�Y�ytC�B������|%�ok��� k��E$&;D�o鉎u\Mv�ݔ��e��ر	�po=ݔ�E��˄e7I3�J�E�xP=7z�wlY�c�Y+�����9J��ڳ\��⨯P��,�Оm�;�Qɋቪ�6Ԁ�
����e�X;�z}kT���^_�J�U���8��w-�J�R�j�P�7Jo��2�6�*Rv��'S.�>��Ux���f;S���cً�T6�k�3��g��d�Q"f�k���R�P���
���h]�2�.�����ΎHr����u'����+jqpƇK۩������A]�q][չ"�Z�75�ZPi?�(��]I�叇Mچ���E�|7l��3��.���7�	�n�g=T�ݿ�~��K��l<����uCW�>�ҧO}�ʺ�G;a/k=���q��J ޖ�mvz;��Y�xy>V��"M��hsD��v�E���d���9��BiW�8}`뼗�ե��bc}[��^ڂɼ,�8�a]����ܽ&�vh՗� ͅ�VB�B�=�M �Q�ސU�ւ{��}�W��(��3�u��V���)WK�8�-�*=��7���o-�>�!��fKX�ew����NR�|��O�ʄ������DN��d���hw��s��k��1��T�3X���9��V�d��ƺ�'y���ItSp4����t��z_=�׏�>o'�Um�e8S
7���ݡ.y:p�XH����{�����k��٨�Ҹ��p�d�M�W@��k�O?H�i�|�Ƅ��^z��&�s�7zU�MB��p��m^�F[�z+�y3٫���ޙ�CM?P�����ƻ��8�Q�,�|h�o!N#7q�w9f��8,|�f@�H ۃ�W��̿�y�ǖ�3~oiȜ�wˊ������Q|�ud,��TJ�xQ[��ձ�>RC������p��G;��抯�P�ે
@�i��/��.�K���H��d�9�ʈ��7u���vgi�SnΑ]��+z�� @�(�u����Y�k�)�����X9u]/�]_�ҕ����Ķ��\���Fp72L\8�R�WW5�&�p��p����P&N����G����5��ֹެ�}x�<v��j���*�PV�A�x+k���4�����.4���e��9�� ؇h�ы�z5�]g�ds�7<��zm�{<��B�#��v���.���2�Q��p�q�!���W}K��oc:hĵ�J�^u_^�%~w4�����5ԝB���疷LʱP����ڢ�\���E��F��[g�M���x�����9���۱O^�u���ơOt�&s^��=���r�rm6�Q�~�k��jUr�cHV���u�	ޯ�{�i�'oiMvKp���=?A{ƥD�/wz���T��>��1~��~�Ҥ5K'���WW��-ۆ��%V���m�S��7o�e���I�t�4w�;������}!4�8}���Ɇ�<����!A�oh��i�p
���a��s1.��}��q�7���z����ad�j���m��u��ɵ��2�p���^�Ssm�
1�lѿzq�/�wT����0o����ęE�;$`J�vxQ��|�!���y��`�Eu��bX��1���u˷r������{G[�i���yZY��][f�����a:��I���U��D}W��9+f�P�u<}�p!)�	L.�	��]�ښתe�ڰ<#���ʎw���Q�2�����"��G�gʻq�Ʒ��+��^�^/GU�Sg4����ν���;�;L�Aw�ϩ1 t[Cy���:V��d�~q��y�.��Ң�5'u=Pչ�3@-1즽'<��s�^ٿ{Y���%NO�/�V�.{Qʃ���mC�*]@T
�Bv1%4��(,5��H������Qx޾v3���]	���ߪzxE���GA��U�/j�!Ji�6�?SW�,�"��JŴ��_V��,��S�	��@[l���5���j���@nב��vs�-�V(�S�\�D�7o��a�a=;�_���;Sϳ��ll��hn�y�|�gg��*�͍�� ��/-0�������:5\[�x�}÷#��ۅ���3���m�wN0_w��8���qK 87�҇�����α�����:L��`Ĳ�kƋtM���A�hT˫[�C�k̖Df�
�_6)��Q��u|���w�������)ب�v𧳇i�&u]Y��۩2U}�UT9h�ów���Z��OI\��\�(k�Z��=�M��x�b�����p^EvR^���B��i���Ύ�WS��˻���{ɴ���\�D�P[��fӃ�#]J�)1W�%�)=O�/���&Ɔk�]e�)�qw�7Tm[��B]���F�}L��YkG��3���3K���μΗS�.3u-qؗ��&�%pͲ�KDjU����C���.�y��6����ߢXߔ�P��#W6�s��݉�(��]�9���e�G_�,�Z��^�1>7~��4�����Ky�S��n�t[�H��Q��q�U:wܻ�����pa��h?OnMc{����͍m[�;�q���R6���w�����U��^[x;~��qc��[_BTr�1W<���p��M�:�Gb�"b������I��_m}Qy���ŀ�v�?|S��g+d�
.G�m\#�#
���U�2kN[�m�(������-;C�b �p�%>�VEL��9���^��@��(���1���t��$F$2w=�뒌_H��00�k���f*=�5��eC���]Tu1]�Ǵ1`�=�1�b��-e���݇���@_Iy��̝��.}}ж+��� us�2�oJħ]���V`b�۶,<F� OMb�T�133�Ў��t�S������	�+�^�uL��n,k�l��j.�j��廇���g�|>�Ў�lw
W��M2Z�l^�3H�Rf�]3���AW6p����Q	�,j"�!��ܡ�oa�*�Ѕ>7r��u�\�o{T=�d��8��]��SP��D������/��j�����u:w��C����M�]]�Zڈ��+�t��L!a8�f�+JΘ�?��9>\��ذ��Z(��1�۬)�)��EWK��눎�X�Ú��\���sv�&u�i�cuӸn�n����!2�%���8_�/��5ݒ.��Ӻ�%��&e�AK��G�<��=�쮾��00PR���&vq��ll�Ӱ㬝��r���\Gdy�;v�D9��ad�E9tU����,�͐���=��c96��x��¦H��
*�A]E�1�
����WgN�l;�����}0ڍI�����1.�׽CYr;���a�t���iN�����^J����ݻ��f�n�iԯSt/0����۶�	b�������m�u�E��K]�\�;S�1�@#y��YZ��e���/;��4唭���v��򷅍��ʔ�ND���r��R���!X ������x�.*@|�Զ/�>}�g[�+���tGj�|�Hv��BԺe��'6�U��Pj`�Z�u�Ν��L��J��jٴ7��T���H�,b�T#�w��;�*�Եr`�L�#pf���\�:�ֳ�<9�����K&n-��t�^14y�uϴ�y����'��<���mL:j��e̝Pg|���0�Dgf5���9er�Q��9*`�<fs;m�W�ʑu0&�H	����gE��f�i	B�N��=�u,>/=����e	�e�`�'8U���O�ЧCG#��]�,Ӱ[g��
�$��$m���9�:��e���/��X�<����t���ۃ4�N��a*S0�nf���oS��l��9�V2a��ڮ�^���ї)�Ȓ�*.t����X�יB�����k����5)4r���m]�[/z��KlheL�鷜� M����yH'�\��]8��ؒ��(x��M�K	rfk�#��Y�����3t��2�������,*\�lx�ŷ#�����Yx)���K&MNݙ,c8�Z4�5�-��Rj[��WL� 텕�ZD���;(�b���C�ٻ�e�P���uC�Wϊ�V��W�3�WGNT=xЬO��%�R-�CV�o)rf_qBA%�G�~1 A�hU�(xJ1B�o"NW+R��^��*��]ܠ�Uԏ\ݨI�ʇ$�w�w��	�QZ��U�uC�,������N8�T^�U��-u��y�x�nU�r�Ȥ��$>5�l�*����4Zm��4�
�,�W$Ą��ȸ_<G��C��rJ��J/)2-d�d��xZȎ���4C��".sn��eNI�s�z�E�Bx�J-KZjY��e���<�����	�"�����s�☔��{�22 �02IE�U�n�=bd�ȍup��.���y+��TȎ�<�xG��(�9���'��-̈���YȮ��s,���-j��p�A\
u5	�p���g������aAQ|��Ǳ�%VHNNp��(���ؑH_U�7H'�I-�A
�����tH�T�0�bMTv�!�6�A�J��ȇH>�Ӓ���Pz�e��w�9���^�i����9���!������5'�ƹ@]��%��;��\+�X��/1^���Z�Y��xV�/z��zCC��MCx2��ܨ+�b�fv�l�v�	��X5����ԝ.�/�ޭ�c��F��!�k�[�V��ZW�\�����A����8��y����ogS��lT]7���j�v�2E|�K;���qae|z�Է7Ԫ�:�����s{p�5��P�])�B�RF3U�\�P�=-�u~�"w����-��T�y١rx�ʰ�U��5���P�f��t��ՎQ�r{Tf)Q\���mw.�<�7y���-������)���u�����>��ܶ�ƕ��������W�c��of�6�|�-�ǻJS��l���9�f���+pd"�H�������3�n~�'������Wg����n-���lN�ȋj�� <<r��V�{C,Έ /hb�N�T����lZr�v��&>i�-�H
)q�n����l�o4�V�K�P��r�R#Y�[�w3aS�T��9�T��8Mf�����O��0s�]F��n��1�'>���o9v,/4��DDG�wJ��]�z+��C{F�鐵݅ٗǓ֍�=N�y�p�Y�u��9To�Z�Ũǆ���%�!5�ĭ̸	�_�VW�1�=�����@���֩Eu[��Ѳ�:����L��JS���V�/(f�nN����N��D.YG;������Ϻ�)��f��������:��;}oVsa]iqy���u�:�!Rj�CYN�+_�_A[�՝�.55t���z{���~*=|����wW���8���u��.�d+�i�{��w��[Ax���*1=5�&��W'��47x�Mnw�X孥�\wP[/wT7�v�.�b�7�)���9�&�O[Dy:r2��r��r6�`���wgu���f���ݳf��O�|B�ꜰQ˗CS|o�G�X�@���S��r��v��`��R�7����@g���t�p)�-F��S��/����F�p�ﱬ�s��e�e�ջ\����ү�)�^��*�x�	�o�~2�}Q�:8(Uw���&b�˹ɉ1w�Z�v���K��B`=�w�]�ÌUދ�UyH�U�]fq�n����	(>��u�B(ۏy�b �����T���>���º�빸Ĳ�Mn;z��͇x��2L�vq]P�$`z�\ʛ��^��c�y<��U�O.1��m�|��_vh]Ϊ�q�$��s��ak�b���U�Y-0��R�ȍ׻�/'�cuL���[���Nw@Y��ن�BS��J��3.��?#&h�I�n#�xks|�RZ[��t�e�����L�O�]ojkf�l��[�v����\�T�����pJ⨋v'�R�Tt.ڃ�+��Z���[��]���S=W=���}�����p_S��3q�؟�K<.
�-|�w����jю��b��iw6j�	Q�IӰ�>��!��hL4�� ��/;k����N�o8��\y���9��g>�!�\�i��*])��yP`n��z�P(v��
ܣM��*�{Q�A��N��w�B�j� �.j��%=d�+{��/}�M{s�t� ~,e{��Ӱf�X�F���68❚�\�5�i�m���gQ�2���­��A�b��Dݭ��o��l\����gϬ��K�n/S؆��{�ŋ1;	n�.]��$S���g$Dg~����u�����L��䖳Un��/�,W���E��b����ʸ�ŧt�ɝ�^gpICF�b�U��ZGj{[9�x2�r�쨃���m�Š>1�b�)D��tTm��WP���mg&)��oϯ����k�y��<T+������j3��R���(��L[�O��G|ѯ{�k���ɹ%���$�0�zZ+4֛�aY���!{H����[q�ۇ���oj�f囒�#�sV��q�Ap<'28��ƥA�u��<���u�UF���Zi=Nv�Vj�75=|��b.귘���nA��R�Rc/�Y'�!'�1����1=�{i�ec݇�x�Ӛn��J�%�L�5vHkhƈYUe�n���c�z�&���v\e)�5XU9H�J���.�-m=�v���.ݩWT�$�޵O�uw|���~��=�ˎ�]�+���o�zo�<�\9.��y��̵ޥը��Ȗ����r�C[��7ݑ(����VK��@޶�f�(�ĺ�N�Niƞ�/��{d>s;�s�Ϋ�(�M����7
�t��T���v�K8cCm�\u�-?t�Ncu䇅ٔ�d}q��������%{��:��c9�?_�Ft�]qR�MG8��Y��6-�=J�&y>�saY��f)�&�ݾ+*91���}V�kR]���ˉ�^b�z1��q1I���+r�u<(�~�9gv���%��=���ֽ^���:'E���.p�>��Yp_m}W���ŀ�}i�E(��<�����*�a��P+�o����K�w��h]�O��A�n����ˬ�etN'�jb�\Tt�_s�Hd49�����ݸ��:/M�K=�[�2��M�:8����iz����[8�}}����s��5���v�d����6O�*	���{U�(ĸ��<طOr����\t�ɹN���Ԁ>�_<��Uȉ�1}J�=�qʾ:�.y��<쮱s���7������t�a�댃�T��gP�~�"w���j���5�Ş�:=m���OkIAV�}J����DA�����.��ͧ�G2����Z-�Yث �{�q�;1�ٝ�5�1�v��)z��l�7Xr�e��m�����g֩�k��yז��(�!��ev�G�Z�ȘJ\9�@t͉Y�L������o0���_������E�<����	�?nu
�щ� v��J�8�Z����$���Zˈ�v�z���l-�
dlom�Z�<K�g���ō+0Yf��w�;�O%�ͥz�n��[�㬮5X���ci椻�����S0밹�\;����w�����ԯp � �y����4^k��0üaІ�BY]0��ٗ�6Ҟ�Χ]��D�]��=IX�����܎����(�.�	��V�XO2����n�$����u ��p�H��ީ�i3_q��M*g�]�VS�a�Ի�U���Z9ҁd�ݫZ�O`*�����>�*�co��K�n��P��uW�S��O�x��\��q�q\Bn��K���	z�zf�8K��H,B����X��`��}C��{m�F�b�Gt���B���殦�]��zG���ꄛ�dU�n�6zv��٢\���wDn�Ch�����[�e�5��y�u�b�e���� ���)�̝Y;Y&� ����r�W-��M)Ya�,]�0����4��ֺO�ιt�u:��[�uh���:DS��K#O-�VvV�ꪪ�vB1�S��}W�죊�-�7�1=7�u(���j���&UF�L�Y��
�n<�z��[dx�]��G�WQ���~ӨJ�dc���n�f[��O���׶1�X̆A��Q_A~�����}d|f���:�'Y|�r56*��N��I��OI�6�q���Y�)d;�A�$�7�r���r��Ug]�끉ci�'ow�b5�+�Uq�5���e��(W4�jm�u-����=��̽��>A��x�"��YU��򭘼���;=o��`�^�����@_v�����?m��8�SJ��tL.��Y],WV��v�x����a+�l$YЗ
�3=�ޕ}0Hg2�5OR]+�u��S~�OS%�8�7,���S�]3>���/OƄ��C��The'����������ü��U��IϺe|c��\;76(5]Nχg.�K##�ބ K1zxzz�;!{.�AO:9;KJ�Ba�Z�+�Qw�l��i�Ծ�ú����T����u:c�P�%����6=�8��X��Q�)w}±�c����]@����f��gr��f����I$���Ndߓ�QL��U}��y�=��7t����̶ym��=��@vپ�����g���'�"�J��CL��{�4�Of��5�+�q<�
�BTr�t�P�ેPl��X;vzwZ3j&D�s2��mE�uZӋ�.{QiYw��Cu�|#�քj����[E��
��nQ�uy���,��:J�땏1������՗���y��P0T;�v��v�����\,��;����/'+���+)N����$%�q��1�!ra�V+�j�pq��7�)�7(�����nBQb�v��S]
�o��gz�R�_��)޽����Ҳ�t5�v������mԤg�O��o�XG�W�{k�-���yN�q��{^r�L����rK$Rpn�<����U�.UꝨ\���S[�޽ ���O������'!�}�r��T&P� �5�ݴD�?,����c��񂶞)��4K�++�t˨N������I�I}���`d`P��hg1�OY�
��q���o�`tx*��N��ئ�F�t�	
�\��-wMvovG4\��|�W
����2���O�t�5���W�1t�a'3��04ܷ���:�a�Ҕ�%\�[ͺ�PwI��>����ϛ*��=oZ��p�3]B[����׿ݿW-�Z���חղgg���򒚙����J�>ʷ�Ni;�a+�	H�ި�`whz]����z�r��zC�7s<cͨ�ҿ��j���+��e_�������۩�nİ�.�o+���P�Q��|��7�_��B�O;���}�F�sҹߝv�
*z��]�|U_D���K��po!k�0.k����nчA�6#sG���r�2�&�=ހ��y�tZ��;�xۛj��&�d�mB�1-���Kj/M<3��rߝWf,���ҳ3�20��T���T۸
���Ye��}�y����1���Ļ3:u4w�0o[�T��QϜ��N����l+���8���ԑ�'8����o^�Y�n���q1���9��/n��oV����a=c��f�����n�����J����Ź����s��,�/=Q���hݰ*�Wy��*�Ջ�YI�-��W�c��3a_Vw l���]'|{��ՌcӨG��]{�;�OG]JC9`z�A�9�ݛΝ��r��Ѩ���ꯉ�ӞB���qߌ~ұo�Խ�_VT��;o��K�����lŭ�fz�6�¤�M�����(�����]3�Oz��yov�@X"d_�ݝb���HX�/Y���W��m���7����>��j����y7q:���Ύ��s�k3�.���Y�po\d�+���kV97V�M�ɱ�DJ�ᩩt�[듬�S��6�k��gn\j���F��Q��\%.�&���=|c�<�&5V������ޞ�/�<Έm�ڦ���=m ��ܲ]���D��ص���;�;����si\F������n�D�84WV�
xm-u���i��zf>�\�`Ԗ.�=&�ޗ׭ά;�[̭	z���B�	��5�YV!��	Mt��k��/�)��ӑE`7)^f�f���(=V�f1�	�*�biJ1_r��}\�̄��DƎR�c���A���[�sY�M[=����R��[��%i5pa��{����'c6Z=J�ޣwԱ�� �s+m�Z�a��&v�;�c/*�N��P���w:��Q���b����%z(x%DE�߹��F�i����QZ���b��H�iR`j#9ҭ��
*�B\�u�m'��Y�,��(��Ȏi�M���n�#��ʮ����#^=��V�X�	@�5#Θ77���1�ݜ+V�l�[�Li���=����x���.�*��chX3[�,w%��c/o���hM\�h:;z����&�,�:�1�Ws{;��n�bfr6���Amr�uլ���)'��E�޺�q&u��Ҽ��>��)#����q�0�\�n��j��/[��]]Ah'�����k]we�Â�\�M!A<LgF�8��Ӹ�ǋ��������Ju���ө@u���Y�WR���{z���ed���_��ꮵ��]s9И��}�|�E��5����k��c܏f���]5[k Ǚ��I�=Q�wp�2����ƅ�}W}e�n�T\�G�hJa*��#A�[2Rݪ\r��D��b7�:����,,u�[]q
&�����S�v�pM])�o\&wP��(CLt,�h�7:�Y��]neF# L��[�jȌi����L��Z�9o�+�c��Qc��5��+�#/o�Pj['�@=����Gv�yq���.��Sa�w�]¤̕�vc�@_nT�k��j���.��9�J�s�c%e����]qNj����:8Ôkw��pӢ��Ӷ2��jQ�V�٧Mg����\fr��� :���-����6��V�/�PBeGya�ե�k�w��j7�_p��ۤ\ͱ���p&���I�k3��-Z�hX-��z�d�4�j��:+�W�*=ux�|5�N���sV���+&]������6��i��k/ )#�J7�p��ˎ��C�:���}���9w�N=�/i��X BG��n��<'i�+v]"�%d5&%�rޣ<���y;
<�؆楉B�|{��v�6��'M�y�R�8x��	��\�,�v�9-�HS�Ư�P�¶Ʊ��$�y���=���%E�w9N1
�VZ���V�]_kd��E�ՠ
9�
E�إ��<Ї|�X�vF��y}�1�쇩�T�,����s���f�K�4�-S�>�
�,��qU�X-VB�q���F茧�gk1ӝo{�b�j#k"D�Cif^��$NQ�c�]������^Q�+v�Vj蒮РӞ}ąe+���H���r��.�)���[$��"]����8ͨ���\�]�3t�!�)��ې��02�$N-Μ�����У�Ց.06S�u[����ޥ��a���?+�*j��=��f�3�@ӻk�BC���-Vv,(��(iwe����V��L����v��[(� ηD����v\ݝ"�r��bO$�b�I8'�y����ݢIrF%8��J<:kf���HO<�i��F�I�\��rGwdyK���P�9FH#˗��V��;��,��^���9�RAfr����Q����󫮦�N�y�H�TO.s��!Fe�z����h���F!܍�q�v8��Z�t���\�t<�mD�Ρ��Z�U�����^ty=%�[�E(���Rsʽn��(�<,J*
B�B���ܨ��uef����Uy-<�)�-r��hd`I�Y��8UT��bE��/;���yx���-�/<qA!��U��w=Q�#S���N��랊2�2��n<�IbUk�h�z��*B�G#�$�uܲ:��D��$Q��D�dDT����K�Z%AA�[����[�9D�yz9��j-2.���-�yגX�#�K�����D�1MUuT�L4$P�IK"!J��/']�"M�*��C�f����

Ğm��l6&��ϲqoz��:��t��oR=X�m��8QS25��,���]������]�;n�����7�v����;�#i{�x��n�ڍi[����Q��	��
+���=���qt�r�KQ�尹^�25��YQ	Q�I���>���t-1�e�����ֳ�b�ֺ�]#Ӯr�\�c1ڟ)�������ѓ�L,N�q�l�=�B�K�}Awm�j��؁�A����oQ:!��s�)U�!&~wJ�Уn��y�2�j�A}�q]G�>+/Ύ�O����4�;q]�V\�J@b�pن�:�!�e|�����B��n���CAߴ4w��<m`k�>wq})L\�'��U�Y6��������۽�k��죋�a3�}Y����~�*�Q�w��GUe�lS��s�W�M���W4��Gm������(gSwݾ%�~*�@T��:��9�Ν��jkU�����
��ܘ�׀7h�ŋ��>QyD[�\��{>|��(71��W�#���3VF��$���%��`�1s�ƀ�b�7��y�e�]��ϥ5���{8-<t�ܹ-SN��=��:q@ѽ̺\� �%�:��hKb`��&������V �97'��;'��y=�����OEƶ-u{�S�����G�Uk�jg����tY���sᑮ��R�Q����O�޻*ZS���.;I����Z�/�*���QOc����	_��Qk�-5�d�X�`YX{�0���vb9��q��G��˔W��*�BS�]2�VcBڷi<7��"�};��^}����*�q���]}ǌO�u�9�@a�.�ս�sU��s!+���&�ྦྷq�f໎��R,����ú�����W&��Uc$Y�K�n_O��g:����|��I���峂_,\�n�jƇ�}��[y}OF,sP��%E�J3Ҍ���KR��s��T��mc`/��ٸ��l����%����=���p��׷�y�\�.��A�lg5.�ع_ɾ����/���pœ�<�ة ��y�[ո��Et��������j�[�kG�и���ZӞ��&��'&+�erYyՕ�〣���|�|.]�@�.���)��DU�q�,�^f9�z9q P6I�GXt�Y	� ]n(�p6�>��Krf6���3*�Q*uL�����Jy)!���x�M�W�)�a�KX��]���[���^gY������0E�s�:��]>�y�v�}U�<�w��5)���*N-n������ކ�3~�x�Fhن��0k�鉭��M�2i����)a;���i�K�w@Q}׼�F��{^�1r�T�Rzo��\�*P�am��-�_R�8�>]�_sv�y��N1�����6{uRrA�S[��y�y���R�u���n�P�L"w8�v<��W��#u>�oQ�\(,��ƺ�%&*>�J��I��Ν��N�+�Qگ(��7y�-����1�f[����r��Nn��+������!p����:�8�K-��W�5ɥk��q�2���3�BOv�
�O�:z�JO�/r�6'�����V�ִ��S_9����m⯭؎�RxEVŎSϻ��i���Q񄦸J�y��۸�o�_�z���r͸�kl`Op�/;lz�U�2�x�{q�[L_ҷ&���o�++��BW!fv��=�8�:C�2y䍑y��x�[��h($�q�S�R��}���ה(`y&Z�Z4ꭙ��j��������v�L�ܠ��7J��e�m#5�,���f�Ü{�a˧��7eq\����Ldr��}uq�V�'����1���!_΢S2ܨ5�x;i�ŎSq���d�ҝ�{Ņ��	ʧ�5����>��
���Y�_A������a��LS�ڬ]o'��f�\���9
��;M�;��]C�:���-:�ì�jf�#�7��� �����*}���hdGj{S6�1��絻�������uy�-�~1�Jĺ��Q}Xf�lW�fq�`�3r��E~�Mx�8�.gp��^�����P��p������<�y��c�-�w����P��Oݕ��5>���P����`ݍ��?_R�����rl���>��O�z�;����n��oj��3^��ѩ3����P�~�{��w��S��x9���9�Ӓ�gD�H��qmV��p[_\����V\LM��C�xb��2��p���O�vS�M�-�ㅻp��ef����9T�K�Bñ�w�I��T:�f^�*:���©;P��x\^+a�b�U��h4oU̥|��p2h+9�ۙ��;@u��C�7#l
ѐG�7��*v����]C��5���*J����x|��5�FWR�U+����5w��_}�Vo&gs�������%��_5�GrX��&��o+���nvmi�&L�������,�,��u%�xT��=<O1�
�����i��³Uj�r���U�ȷN�����[29������r�rX�����¦���:ֲ =୵1EبG�L%�F�{����-5usܙ����r�{M�;�7�wS~���xK��o.�Be<ۑ-I�7�v��f��v@W)QU	:��CY^@�z�i�㧓{rOL	;ٽ��j�x%]]눵�-�O����BmF5R�+c1.J�{ˆ(��]�����E��ՠ��ޖ�#���n�K��M�΅�3��z�y"g�Snk�za���U�:)腉�q�DmEp���\�.{���|�����b��ʂ�-v�8��e�;�\������]Fǥc*�k�m&O�o�zy#Oj�,�@Ua]���{��gP��e���X�q��-v�{�L[!�)V�s�E�n�y�Ⱥ!�2q�w���R�m��QD�=��	=Q���Vo��
z�ǳ���?�}[�2?W��Kg(��m7��^�-��X��W��Oov{��XWVŇR�/jR�g�#ݿ)k�\�<O�>W�M�W�lm�ݣt�Z|q�n�R��2��]��������~!�
l]�W�����+�EN�� xV��]{o}Th<��d���};��탫U�O/ݔ0ܭ��u��q�4��.k��am�($dc����+�KJOY��*��}�5�ڄw�eb�v��ZR�c��q��T���^������ǹ��(���5�au6����z���e9E�9@��K���F2&MI�U}�s*e�]�p�:x��9�P�h�n1T[�4�����y���&���ս�����.��i�7���i	n��x����4]�('���2pr��g���h��@ĭɨ�Ov��s��BN���Ώ�N��s�e�r�C-p����nUON}��������k���λ��C�H��z+�d��0-�wWw�k\��ٯ9=X=2����R6����)��}�KO�꺝be�t0<N'�O,����]��}L�a��]<��ޘ���mM�e�>x�`�恦�ri.�M)ΐT������U#'�}��Xv�����{�@��}����*�u�mI�~}���� ��-���=��[����?P{U��w�)������+ː'0�@楹�25��Z�\^]�jB�z��7��P��X:�/W��m��7x�U�˟]� ���q�P�pb;�;�֫Z
��<EL>2���"_N��&pOI�-���N/W�Ә��b����������fo5m_[�^3scs}Ӕ��f��Eq��(��/5Ի{&�I�^������3(��V������*�݇F_���{>����|� ꬵ��z�iK˼����2R �󍼔����y��EN>����'��%AU2��܉�q�����t�ҫ���v(��Y�W�����z<�Wq���4��G��>w��f6��sM�
�BSa��<�O�=�f��԰�:�h�E���楌��.��Az��X�]My8�r��'�U�=�S(:���k��ցۊ��޼���U�9�ʾ��H�
J�8<�މ��"�|�n3D��4g扼��b��v�軠�v����lo5��ﾋ9�.�*�_W��^r��͟���&�����wl�b��k��H�X2.�R�Qz�A�~�5��f�}�_)k��
�1��l3#^V����m�́B[�>���)�2�݅ٗy;��?3��wcEc����3Fӯ{����ɶ����;\-��Щ���2�1;��Հ{c86j��y�n��W��FfҸ>�*㩻���
�;s�ʶ:iᳫ��w�����se�rg{�6����ۄķ��AV�*�:��ڃZ�ATKɮz{Xݥ�uױ#9�c�ޯ�S��!T6��w/`+������J�c|�t�-����+���Z|V6�(��n��t�d8��j��%��1ʯ)�����{�{�J"�Ҳ����>�Q1Ԣ��}������)�Q����R:�_��q���;t���Vtc�\�`�4���TLaȫSkHـ�Ҭ�n�������-�yݑ'��_���^��Pj��z��^�{�w:�[�7��z#+<�:9�N��{�:��g�I7gn�f+����ܒ�I�m^N�������GpC�UXN����l귶N�S��fy;{ܯ��M��싘��~��UɅ��Yܑ9�Ӭ�3�Fl�6�n�'ي�k��m�����t��jTr�o��W?eP��'��sC����
l5k�����o�ɦ5^+��P�Kmt���S}2���@\�`4�ܥP�h�o/���mmGM1��w��yx7f�vy!@���d)���Q(ĥ¯��Z:~V��J�,ɩ"s�ɸɪ�SuO.��lu@�����s������&F��]��m�|�,��׽�]#M�.���;��g��݅�=����m7���罺�w��Χph���U�D�I�אa��F�a�4W'jf���j����`Rn�s	7Qں�}����C�R���ޥim�݄���WT�ԟ&]���/���8����Nw��>���t6�M>৚��Ϸ�#��QZ��[@T��m1
���B���k�7�p�)��r�W[{!���kK��5n�=%f���<��h�UΎ_3y��o����fK7�:TVk�zQ쮖�gzi���f�e�����b��\`��+�7�X9i��tỦ2g>5��S�[�_l.].���W��]1����ՙy��%y��4�H�du�w	Qt��֜p#k���h��ŏ�����a�d��NNu/��Ǒ�M��Pԭ���)@�P��d��M�WK�v�E�q���4���I��w����H\��F=��I�C�t7��p�\������1��2�.��Hr[_�}���YɊykm�ڏB�j��{��[gᥙ������Y}��5Kv�伱�c5�o6��9����z��2�3Z��]�{�z]�bXls��O,⨋;�:��Ĳ�m5��������̝��z�C|�=�9O(�x91S�bu�S䯶��իBv�H�'N(k�H��q�6��򿆅�t[��B�$���W=E߹��9Y6>�������4�W���n��6�	H������H����,�5`Jpf@�5r��r��;Fwi\^t�#��1���Q��b�qJZ@�Dy"U�+��O5��h�+�k�V��sY�4�GYw�n>�an�	&�����b��ۨ恗��A�XZ�q-a�|�P�Ӝ��yg:E��7��m:�zг��
[e>���U�	��YY��*�VҢ12�	:Hӕ�.�E���3GS�y��wWs��c[/��Stji����J�;T��Y��%����!�W,Q����A�n�:JF��K�W,e�v��_pi�c;�7�V�.���P�m.�U��[�� �k��v��R�OG��B8���h�@빨���ʙ#U�v_t�W'���g�ëI8͚b�V��v�b�r�8i��hT���]�P��,��]�Vf_u��X��;i�HQ
X��'�uo�=����F����eZ��7T�"l���Mk��j��Z�c�$�
g
��fC�8�C[ۂ�g:�~�w6�4�y��9�u);t8 aU�e3u�sxo�ɽ|TFf���:����e�:�{Kg��m�yGF7Y�]ov���|�,�;\-RU��d��VZG���U�>{2��;b���lb{e��K�c e�2�]� r֞�K�v�l��C���}a�X�ڴ)���/A$30�I� ��T�3M��4��뻉O+mլ���;�\�Tд�X�}�σsQ]2���7%lܻ�S��Y6��w�Aț�[]|M�;���	�+K�H�[].՗W1"_C�<�:q�q=W�3�!GS,�ǩ*y���s9�s��41Z��Ք656���ñq�ZqD72+�7N\��3��Y�a��Ңk+J��է7_&�I�tԫAb��$�d���T�ڵ[�Jz&Ԝ񘻊�����7:ގ����hc�
t㔀GT �}�n\y��Ή����MgK�����iT5at�/evcz�~~����F�z�+zU��(���]��n
�`\Օs�+�CF9`jOZ��y%ͥÊ�pP�e��Ս�SX�0O��\;�Y[��n:�WhжU�<H�F$-�_�vP�)�ƃ���V�%�{7��{;��e���)�p��ݦ�V�Mv�w8���v�>ޡЛ[I���-"��g���������&�^�G�
�-hiשd�_+��opto��6�m��݉�#x4�[<ʢ�o�HpM4i&N.}�ɾB��ۻBњB��X�M��y�CA��10�n��mJ���b���L�H<����8N�k1��>[Y�b�]|g��,:��S�7QT��/�]�73�n-;|s�Wj�,QE^/�
����f,���9K��ea�d �2*��NYsia���LmKNa���(���a�P7N=���I�6l�n5%�v4*j*_L��X�#�&:�w��t�錮Q�G�on@ٵn��lz��W2ܚQ=V��C_Y�h���0��u�U�Tt݂b<N�I]C>:�E���w�x�����<�:�S�Io��x �{��D".�W�z��˔�y�*�LT����Y%h����8_���G��$E�%n�R���ꓙ9PR���f��B.�{��y#��
��i.��D�.PQEF�����"$s�H�f�F�Qk6�W���%�H�K#�2"Z�t��B#�"��ue�J�\S��rq�)h[��̊4����b�V���̒�D;�������B�^Z+���u^Z��֙E�`TRV{����%�i^�^c��4��1WW"�RI�y�us��(�-)֮<�8�o"�fK�A�^GVja\�#RJLˤ�1¦�I\�L�wR�ܒ7v�/v{��:���GH�*!O7�燄>yܞPي�r��V�f��d�������'\vU��K��d�%	Y&)�bWM1@��]�*![7^qw���$�0� ���iܺH������ǨFu.W<�ˡ��$����$�\u�(�"R(EjJ**IVRR븚���y�z��w,ə��w�t1��M돂I���,���WֵuĒ�z��n���6D�T�w0�O94��&�\����r�}{��γb�r���6�{��qB�5�v�j�dӥ_7l���\$�~v%������'���Z;��1���SP�U7�9���n�"���R��	����l�*���~�k����d��Rk��V�P��8��s�������n��\��y[���j�6j�x*��;w�(����u\�����/�"&*�ˉ�])1 ��4���xf-c��9�$�4}V�Y&C�=8ou��%_'��\,��ߏnQ�uy��U���K��o{�L�Y=�]`/�J[�w�C����CyN
��Yg�M�m�s��@�P���~q<���6��;����j��2��g�t�]����&������O5�7l���qչ��c�z��90�ߛ[O��T�\V�{�X������c�U��#~F�)��qf�yuu�}�:�/������n�FG�81�x��%�e�ƅ������$��சں��.���ut��O�����镫)qٛ��_ޏ�9�x�2��){E~��}[�A�Zt��u�Q�f� ����W�͖�\s��'��u�L����M�3��`��y|�6c5�cc1n��Tǯ�oΧ��r��r{ө���ԫ��=Y��c��ucx;����XP ��_Z��/��X��<�ׯfq��XZ���wc��
k�j���&|?nu������������Ae�w�^N:��|���z�f[kj'Ωʈ�5�t��b�~�KyM�� ��g
��_v����Qɥz㶢�Zr�r�=����P�O��R����Ϯ��v�*��8��e��'DD�XY��,��`��/j�Eh��Pc��\ek��/�u6����=�&�˞�K5�Ԡ���ci�*�v'�R4Tܯ�s���+9��$�0-[�"�����K���MC����Nc%1�����[��oo�L��^iu>Y_%G)&*�P��t-1�e���ZP1�ڿ���\0��@��f�.������\ʗ�Y�g
���ѠJ��
Z�*f7��S�K������7��='�9Jލ/$b
�]��1S��!v�-���{]y��� ݄��Ԝ��wo�K�#�{����I��}���^@�ݩ򗱜�+���j\7a��vn3���}2�yRn��sr���ʷv�3j7e��p��M��ݛiv���m�K�]ط�w�b���::��rպ�ꍮ�ce����WN�"�
�n�W�<`��g=��#�mܭ��?���<놕*�W3�f�=V;�<�F�K6��6��g���[do~��8��o<ML�V��Qָ�������sb]�{��u�K^��n��{���.n�p�y�g5_ѓʠ�cˆ�[���d*��~�C�ɻog'�mOuh����9����C�r8�q�����4�ݶ��Y���BL1\��v�CV佘{P�Ldk�P~��U�Yp�r���޸�/(EK)���#�E^<э�{��_%	)s!.k�Z����u��$;�X��^�[�7+)�����6��. �'�&�]Z��<����F�f,[��[�$�W�{^�n:}�&7�-�qf��0��FIS/oA��aBqV�\�$�[�X�����lv=7��6�J�T���{�+�4��{�u��5���2{������o��|ܲ�B[F�7>��{m��7qۛ�4����{��K�騅:��y���T�/�J1Q˶�s��;<Ul��ŵ� ����	f_��]9�p�3�y�q�����,�"���Yͻ
(_$��6���pi�^�ݓ��oݲ��Pڄ��p�O\)��>�11�Eh2���q5#�7~�Ү^�E�7�F:>c/f���~�A�s��R.��ŮW�iS�U0�Pu;��`�W���[/|��:��y��'���'�=�"�skXR+������Xw��T{mѾ�����v�W�$PI�,�Y���Qj[ߛ�\2!����y�3֌�z+]�8�dus[�C"?nj]�g5)�D'K���{I����K?w����k����m�Z��Ao9vPĽ�dy����#����Իz{Y��lT<O�Vcu����Ŝ�L��l��m�/)�����m2�x�����y:f���S\\�,�&=s`�ʝ��,#U����:\nh��M�6X�W�V��R�_Z����x��0\\ԏ�.U�����ȉį���uk��������k���:�B�R�x7-��jq���n瑾w6ڬ����!v�M`��>�~~��E�_�d�>Fn�ٞ�ǂ��Zo��)�;j�+s�U��2y�Z���7���f�Ҭ����s9n����5�㍅���v5��s���k�����G�//I�~����������}ҕD��._8�fv�R���u�]���{����֦���;U㌘�I[6ʱ	%�Y�C�3a�݆��6;o���p;�Z�CĦ��%����:�6�rx��L��QTz����0��\D�yave��:�҆���ߏ\��W'`���w$�6w:��v�ҖxY]�al��'>�O����sW��^�ʝ�M8�\���W]8���Y^B�|�8d��-���O���1��rz�m�+��q�Q�l��6���.�*a�;,�ڃK�/1:
��}��{h�p�tS��E��wU@�E�֏����Ŝ�ʻ�A�i��Z�7Z�ܬW�����}�(�θMa��74w�jR��U����q.}\��p��֙��U�iQW�Wd��b��=q
x�wy�x�+��f0�y���]�ӯX%����?Wn�~���!냵^���2�֖\����2g��&�c�����+�bS�:�՟I���\2��n��2+x�Z�77t��ʥ���>����h��+�K�z��Q7�i�KG}�,�����0�7gu�ԥ����niw�UdE�*�{U�.��HQ����r�d���� R�'��o���W�(q��=�oo�/mQ�N�V����0���!�:�}�'��Kkr�����;z2I\4���h�w�.s=�U��_T�M7~�]��}>��.O�!�څ5�j�� p���*Fe���5�c��D��^~x��L�
z�(��|�8���8[�ۍ�M��t-x�)=n�c��ÝmLv?�tnT�����������p�U�wn1F2��N2��
�biN�k�+���y,*�	H�J��b�7���dͪ������gz9w��J���~�;q3y��g��f�n>}95<��J��,:qWX���Ժ�����n4۰�m��ע� {3�ۮi�'(v����GV|@�2��U�yr�N�rP��8���}0��^G*t�&���By%�d�D��5W��2P�.�{������Y���酮��ˎ)���0L���Q{�%�[r�uM5����Qn�"���z+��,}��x6���y��)��c6ʠ���Iȗ�����s�Q�3���c���T��7
ޞZVv�x���q���;��p���vs�,��~�	�X�|�&�����oGa{��꧟s��K�j/����������g�`~:��c֝Y>�G��NϖM���Ù]������A�^�+���G�y[���^�p{����0�W��I�)3�˃g/�Q6Y�e��E�G@�Hɼ����#�k�+�k�'�����{H ��
}=�4�r��� ����v�x�ϼ��u�P��V�<��z&|3M�N�q��
�2|�{s�֙r.&�¯���t{:��>�m*c�����e�Dy�#��W������#����TP�k�梣l���vߖ^t{,׾���R��V7���=��W���}�u��Q�Ä�|ٵ�5sGI��p��π�>WU��}��<�[5x~�}3���v`�TW�v����'$c�f��v%����:w���/�ĩ��su�t��.�Oh�� _V|{�5�#��_:���U�>�Xd^�b�=����X-r��(N��#5Q�Гo�!Π���G��7������o U�<%���+�iy��z���c���=G�+�z�dzt|��-�\��W�f�;��(_�1�ؙf��T�U0(� g�ykn�<���>�O�z2#}���O�r-�W�u�a��5\��p;�p\�'��_�P�O��"ovW�펨�j!���ٜ�����U�s�O9z�P3ק��Q^	w�F�O��)�,�'5�<sq^��@�ђ���1��k�ɞ������7���W�#��S9��'EE����{��]� 7�LDZ��=l��{��~��5��7�~�PZs!�㑭�o������x�|�#O���e��h��I�����p�^�{����fǡ��+���<Ό��i��cm�["=T���O�9>����{.WN�U!/���V����T\nկt�'�'�=qu�2�LM5[F��>��4������^7���L���j����N�M���D���H��;su�2�L+�WI���>�j�8Zv+*/Z�g���/�ȕ�7��x�.ǆ|^
#�����f��ݨy��=��V���0X��{T�uOP�_-,�(J����PV�1]<�lutn����Z��w���m����u�&�A��.�N���R
�����(	zE�˶X2CӨ�1�k �m_�J�q�ub���U���
�9�ܖ���ל@�^�;��R�Z�6a�N���~���'�leyݖFDz`a�5w ,��hIG.e���e���V�>ك�� v�=��rUgH�k�F�n3��TF+y���<J�9(�{��*���ǆf��m�X=�ypv*̳���7�����:Xq���ͳ����_q��*�{�x���;<��H��/R�A�DI�:������Dw:�B��یU�.��<���q��ʆp����GY�Ϫ�E}���(��`��ğa=qP�k�3��d�r�;J�j�OI��r��5{�}3U7����@>�9���;�c��6�Y�%I%;5	��ü2�y��B�����Q�E���+J{��z{����L���[-U���9E�� J���ޛ�������4��Y���Q�^�=�4'����=���9����w���ש�7%���,���"o
������z���K��w!��5��)?W�c�;���20�W��<��'�3�3�X�fs�s=Y�Q��1�_*� {�Y�.W�c��w�v�\z��C#��E�o�b=WQ�����e����*ȵ��>��8q#aܧL�XL���v��a��:�uZЀ*vaCh�L٢Ʒw��*��pX�~XTT7*a`u���u6��;�8	�	���fP�y+7d�ǻ}�#��Qo���y�m΂�ԝ�%>vv`r�Ѽ/J]0�p>(ݫ���;����Tz�A�;s	�E�&&�W��̴{����$|1ם坊ދ4��<�W���s����\y\?S��Il� =*�&'�}[F���F��W�ו\=�[���=��U���4����]`_��`�-�J'�|ٛvl���['�{2!3��ٶ�޶��}�U�s��B�m��?X�s��X��3�V�D�c�6��M��/�y;���w�_��LMl�i��],z����|�T\���T����=��p�{�%��������Yrk+ٿ�S��u�?K��N������޹�3{L���lx?Nz���~YV*Q�C��Rn����������'�o�)����\e{��p�}�L�Uo�F?m4OQ�{�����~����Ka�����|(Z��ٯ�w�X? �}�^Ac���~�C�CWB7�4tz�/�=Ǝp[�
�@�d�5�o�\�l+N��q��\2�G6e�=7EWخ��L寮ٞ����d�b�tf�۲�G{���'��+�܏?_��_���\w�u���8��Uc�늦��ԇ~��a(L���m����C��>�Lڡ�*k^:x�jGQ^�Ի2��g�ֱSw)��s�k-�Bn��4�������-�
篅-<�0��S��q�x�;�#�$6�ƺ��#*8��To�_.��jgp-��v(�+S�,Ү��k�Y�{�^G�<��N�S�v�#;KxhgK*��'v`�X����:��.tޔ�XJ_-`U��� $.q�_NPIS�xT���2�
���]s\O�;���E������n��sz�`F� 꺃{�ї�AX="��O����z�v�s~�ys�*�R��kx�B���}f�f���)�fer��҅�+F�5.J���|@w�EuN��3!O �j��s��wx�n<������}]lu���JM���3��Msh�}�s�8�7[�6v�B��C���u�w0)3�ع��Y���L�t_%4l����5}�w^kmFEwL/�{�S�w-P�'+M("R9��j�L	���9u�WRgu.�P�j�[i�m݀��2��J��1��]������*��gZֲKd�N���S��c=�|;R2�	�z��m)385�5h��m	t���|��9����M�:���;��[��C��S��x�'2��H̢Msd�fX�m����E�:����U�������W;��&|{Dp��d�4kk]�њU�uٙ�9-�+���5K�&Д`�����������\�vlU��[DSMuwjYv�I�,�,�.7�����/�6R�W���ú>ۇ0^�� �c*�`��>{i�:�?j�τ���%��$m�`T���`�*h�Q��*T��S/*�C9KVE�{9"%�ǜ(���p����91V�^�ȰU�#F�W��Q��]k�՛7hf/���(��'&������p�K17,�N�\��kɄ�]#��jU����m�s��R�\,MӔ�7X��W
�t�(;�̝�@�x֛�O�]a'�]��0A|U�rak�撽�J���Ԝ�"�n>ޫ�|�8m�����è_.��'g����H��-�W;Y��Ÿ�e�X���M�oZL�N��q\jᢄ1P��=�I<B����l�}��jJ�@�V�.�_#}��3r�N{x;�t];�1��_<%����sXn���_*���o&V[�Sᙶ�ݑ <�L��J=y�ػX4u�ΕoR�כ�>���W	�̣�um�y��	�J����[��J�i�]�.�a������Sn)����q���4�+9�����9�*�,��;�d$�	lgg�N�]esC���D�gd2,�S������V��6��ζ�wfh7�P�;i��~D0����1�hK�4S�ޚػ�g����#����x�U���,L����%�����XV\q=n����������P��W_]>�mi� ~(����,��d�G7t���8nj�wO��㻥y��yq�1:bh�R�#����\]�s�)�qӬݗ�(sJ�ws	(DZ�륛�����uwy���'��G�Ȯ���n�z���r���u���U_5L�Gg��]�R2	LS���yw\;�t���"��F&�z�5<<�5̩V�E���Т�6�J!Vt$'W�B�M4ʂI�v���:W���{s"#ի�t���/#%�ܩP�t�>2=5�dw<�u��D��B�I&H�� �
Op��܉�3;�9�R����<��u���J�����黺�t�LE	&TRΒ"z�N9�yw�<t�,�-Gw'KL�:"K��R��^#�]۞NUܖA"�̯P�s�1w]H�Z�^)f�\�ˤXp�]0��Mi���*�B��Hd��d��Z�Y���yȧ�(��Rz�=9p��w**-g,K�
B&v�'�rH֛���a����E�+K��Ы$��6�aa��r�dUb$Zbu5u����ʼ�,� |(  �H�����ge��^���'�2Ut���V��:A�ކ�κ�@f���*��j��6�Dʖz��t̺fҷ�L�d��\�G����<;je�s�C�a����.܍6��7���.�a5�o���u�?�1NI�>��U�MO��y(y��2=�~�<��83Чt�����W�d���e��r����N��и�f�Q=F����LA)&�W�܇�Bx�hX_?:b��<�_�
�~Q���˕c!���G�9��� �j ���ʓ�^����>�*�ZF��}�*�V_Fv��F�����7���:��O�Bp󞸙�Qjh��:G�7���2�:��X����r��A���qW�yZ��g�W�� ��D��L�7��M�=Qj����{"�N�}������a�a���L�7�Tw���Q��>���^����I��h���T�l�/��H���㾅�o�:��Eϴ�׳��������/��c�H����&3����ϳ+gUKK��~�i�I�=q7P�m`}>&��u��K�����C��;7|+���r��w�j����z�z nQT&�7%�۝�^���L;�6������^� T%~��y+�w�x���˺f̫ݮ�S�M�;���^-���5(T��˿]�����T��\Y;B_<kE�Is	�vMc�L��Y�94)��^;�'q��d�Ƭb;��GL��� kS��$f9���F]��|�ˠ��(vn��i��^w^H@�[���5d}`G�v���tvu�>4�����}��2=�Z.;�'�\L�v�j�uC͙ñ����/O��w���.�����\�W�v���x�(�>�:j=;f���ٯ�z ��3��<��KY���y���>Ἔz���P�����:����7�g�}넍�⸫�m�-�::rp�ԊႺhՎ�w��j�o�W�k�o&uL^�B��Oz�n5>���~/���j=�W<��70'A��Jz�{'ט��Ni�NN�*�	��|/���ͩA�uA�����yϑ�\�;v֥6\8ۺۻ��wJ�(;��u�A��x�O�����O"a�R������Ō����{[�և�O�U�q�y�\{0^T��|��X�:�8��C�M�'p������?���ߕ�"'���"A�З���6s��O�w�������1NQe��'�no��Т� xN#5�>��{^�Q�u�h��F��O��j5oԑ��Oe{�tU��z<K���0w���=��g��6�$vUVZ��o�z��*{Nd�i̅���kwq��~9�����F��e�Qn��lXr�&�~�Aح�W�����q��&0S�):���7�=j/6��,t�k^-���uҙ��N��O{b�8R�{9�*Mn%*�<h)�P⍵ �:o�SM,�����C�a�ձn�i�tz���.�hT[˱�C�[ �hv��ei��A5�\/q[��J��1?ees9 _od�v��Zw�����=�U;���雗��.U!����x-�\�;E�{���Q7%��u�+���5[F�χv#Lm�W'E��p��gxeƼ;k�֨�p�O���vp���o$�ߦ�d�]���Z^�U���ps����I����9����j�>�~�=p����
#aܔr�X�6���C͟i��%
MY�{�ޯv�7�	{ٗ��E�{����.���e7	(�,,;�N��Y��R/L��-5>΍�T�|v|L�����s[��s�o��qW�G}�$���E�z��&���h���x0��~ɭ>��
�o�o�8�7��mc<}�Wq���\R�|;½�ٓ7��yݸ#��h+ƌ{�E{��.����kK3�7�v�{0vx�^�^�⷟��xZ�4V�.]�c}[�õej1q�%#q%�=uP�j1]1y3��1ˎҳ��a�gEY�^���B��7ק�μ�z��S��4d{�)�=%���jި{Hgx{h�	犫x�q~�e~�F쓌�Rg�
3�2n�����I��oo�7�kŬB��-P����Uv��>�۴7�������-v�v�r��/RM(�۾7R�����Μ��^�4s*d��L]KY�!L�XUȜ��ذn�8i�2�Nc��Jm�*	��Q���2cH�;��?V���_�����ew��<�R�Uz܁(�;�->�u���[��6��i�RSu݈�4#�ѓ���ՉE�*�4}M��}#Ǹ��_Mz�:�^d�����:��~dvz5�->w�EmУ��8|<�(��Bx��'�HǾ�x;^;wM��C����1T'�����I���0�5t ^*�+��>�ح
�u]�{�H����K�|"{�W������>��̂*�3p��Z=q10�_]"bb�W��ĵ�����z[<�I����X*��~��*�'ׇ���)?^��q��׍�r&Z=s >5�1O�h�����P��#({զky=��r>�!{��l���>*� ���Qo�Q7>l͆:�6�]+;G��8Q2oos�߶M��Q|V�7f�Z�M�y�G>�uQ��;�Myϊ�ϦX\i|/����(d�"g���C�gw/H�b���ft�I���X��{��������U��8J0b�,�׾�^ron�G��M�G#������ٵ���N��q�5��*�dx/N;�W�R�E����Ѐ�ӴF�p������[��Q\�����ڼ�3h9$Z���V�S��<�;=�ʋ'}��o��X��e�y�*<�� I��)|��e�0r�d�0��X���L�7���zh�T��Gl��33�=�OvM�j�n[��k_TH�Vs؞H�=����2�������ӳ�}���8V�}�L�V�$y0Tl�	L�}��^�O��C��!��h�����9��aՑU}����WY�r�[|�������������C��D���=�	�
����Z)��(���zn"���w�����rj�b�������v�����{�1�z��";ʟ��_�;�����9H�
˼�3�����ʳ�关~eI�.���{Q��&|��6�x��ά<�.��"=�~)Y���W���),���L{L�������=[x��n�ɝ�S��o%����G�<���*|��+M���4r�d���"�(3�/{�oPY���U�q�F���d��R<M�����!S�_
�v¿ip����8�y�5�z��	"=xw�oQP�~��ȅ;�p���=���F+�+԰�A-f}�
Ep3�=K�[ns���}5�C������v�/=@xS���o���\<�����SB����/gJɘ��y�ϵ�ݾ�=��5ϼ�E/�]o� �k�Y��z w��"�˕'�&X\L=����ؙR�i�h[�?���{�V*5�mz�����l�\���Q�de����8��fU�ؚ�:��&��;���B�5w��u�'|���y$���*����u�we��hIZ;NY��SIE���*�	��p´f�ǝ��=Lj�x;\Ɉڍ�Z���~�=�t��PO��7�Q�y]���W3�;��ߕ?S�� �m��L��z����^��v���uᷝD:�ZdTo�|{��۳Q�ύLtG��yND���w>�}�3~��/��q�2���>��Q/ND�#�7Q�y[��O�I��:��c���K���vyJ�]�W\S�X���	s��_u�ZV����N�/ten�w�^�q��f�������}�jk��G�ު>R|���{.�<�c�x��L�v�j�uC�ڭ-lOS*X�_w�������������{ �f��o���>�v~���?Z`��Z'P�=2/ُ�:^�Ρ���}�^�q�����n/W��{g��z�#y⸫�m�7��x�D�s����َˠ�����EW�ɭ*�g}1k����ޫ�z�ǟY�\u���7Q����љQ�o�-	@�Q�F%q�S���T����b�g_�6�s��<�l��F}�:�=�J�����t�_{�R�����s[Q��1ލ��j$�7T���D���S���aS�D��V+�zА���m����=v$7�[ٻ�d�ig7�H��s���Ƕ6A�CmF'.�*������|:�pE�L�S�B�����e�3.��49�yx�1�nb�"�f��F�}47��ڤ
;|�a��:��m�ݪ�I7���U�z.V�����P.����>��ޠ5;��S��v9��'��_�P�LSt��+��z�!�TZ�ڪ����㾉G�os��|=)�q>���C�z�+�Pe�@!�@nv+�@�yzdFT�sk��|�<s*�`�2[/}��+��^��G�!���[��UzK�{3�6w�-t٤����9�͏!�ު�3�<�]O�߻�Ȭ�+�Ģ�ޑ��{,��ם� W��s9���4J���|�\��ujȦ{��Jӹ�p߭��G���c>���9ɘ^���`�w`V.���wfA�s^��ȉ-���}q��b~��h޹��FX���u)����QM�C����7�gЧ�'f��@z�z�*<�)�s>Gnn���n�Y��=������h\�����I(F�fئ/Ψ�{΀����xax(��<Ĕr��c���^7��}��[�Q*�{��o�J%�>;<ɛڅ�M�_�$�ψ��Q�n<��&�u4В�\�N��t�X8*��.�����8v��H�gV����ٽ)��q�,U�w�5��w�|�G�:���:TDZ��*�>��M_v~���V�A:r败�@����!K��Ԇ���v��v��\Ҝ+�	V9|=\%���a��h��}�ӗfm.=���.��l89ãpY�t�Xiլ��֮X���u%m���NK��7�u��T���]Z4�K�������Q�yk���ǐ��i#���d��}9L=W� H�X��5�e��Z]�O�i��#}7��������d�,�W��^r�n}A{+=Y;�#��ގ�G=�F2=�{M����2�ɭ,^L7޺��^�"��9�
��;ۜ�;���>�W��o�hvym�b��n$�;f��b�&u����W�vj��ܣ{�������?|����3����G�y�xo��(vzw�,57�MCb���V{`�|�o���܍�j5�U�mT4n{�p�8����L�8��~-իc>S�Y�@(}6�Ӿ�%[������컽}����ov�ϲ6hj6ߕǲ!z�:�#��w��n%z�/�9E�w����g��L�wr��S��|T��=R0�|��ǙǲG7��U��l�w�W3���6"��Cja��D�����p��zc��GM2X�0a*���PO3bʞf֪a�1��<&D����W{ݽ���}���K�ߨy��0[�j���W10�Qt��}>ä�wr�=p�ϒ����s��{'s��k5~�(z"{����
Ͻ��� ��^6�ȉ���^:"�Vџ���*���qJ8���tխ�
Gu)�j���g�,�}]�e�͗:��	8�T"_!dݙ�V��~ꎌ���;4;�(f3�w��(s2��$ax6fQZ�.��o+ht
���rVN��#��ZV��:����5�p|�{� +�{�_[�M�ςۈ3a��Cu��n��}���]��P����Ӳ}�ito�J_���m�׮l�{΀�9.�=a�|ωX��ׯ�ۃ9�h����h��fօd���fit�O2���v\�G�I�^�l��=>�>�f=�W��G�I��NIl���~��Y�8{�s����U���|	��j`P�B�Q��6�[��"<t��ЯUŎ(�_��#����4����k7�@�\g[3|�������v��P<�$�ܗĵu�}�$T=�Z.<�Wqȓ�:���ڇg���}��e����K�o�� ��R#*�߉�[8�v�������Z)�Q�X���Enq��1Qr�>͹�M����C3�^�>f���y���^�q��K�}���7
��8l{'QY����)T����y^���ٍVn�`5��&��
�ez|3jW��'x';��~/�{%�V�4��)[�؁�pH=���i�P3Ŝ�l�>5�OH���1S��o%����G�<�h{�3�}wH��c������p~'��w2P^�t�g03l���:�:@xj,��jP�Oq����[�ꖋ����8�N)���p���hM��V`��P� A��U!�z]�l�$�ݷAթ)��Z��F�܀���wϪ7ˆ�y�s�]�W��}.�ޠ���qĢ�e�I��Q�zQ�U��b9E��q.�A���UH�%#��/9���O�օ��n@WM-�;;�7�B�@�{G���|{c�LC��#�>��f���!��'�7qT��^�g~�?#�;Ϡf7z'����6Խ��I{e���ED_�܁q�x\8�p�5�@Ǭ;�.���yu�7�]�sW���g�c�0�}�+�N�zϞ��� ;�'�uNzNL����~���
����fǰo�:��{No�
��(�����y]����>��K�{�@]�߭u�3�k��mX�D��|v���TC��V��wǲM1�Q��s����b����M�j<U�7�k.��`>��7XM��^�>�L5���]��t��s��.�=p�Y>do� ����X�2���{��P�����rA��$>9���[��׸����f���H��9�d�\s�)�� �o���b=��':t*��n`��<���'N�͝�xn#=����|^�S���^W �Ax�Gg�Fu�Q�݁i�#�>���}�t.�Z/�=�ǲ&|3L�X���ZL�Dkss�9Eۗ]*[�00�S	BTәeh�n��&;v���ϧo3"�ɉ5+���;j�1��C������1��I:��˭y�w���k��p�2�
[f�>�W�=]W�-��^�H��]A��
��%ýݝ:�۴��n�����u��K�#��)�T�n�L�Z���;G��\�����ډ�k�J�����d������[���ռ>7ql�U1�د.-�5�\z���۫(�li��2�s���vR� �e��,p���n�+�5l����-��IV��h"��2v��Y��wx��h�rp;��h���PV�y+4����:xL$�]|� �	\������
���n�d�|�
X;��a3mKO-K.���3p�5�hӭ�!����"���9|k����Gk/wGض� �*? -�w�t:-��� ��Υ�x�7�l'�,l	�y4h���$�J�c���
�����]�uN�܍M��q�8,�;��@��Q�M`0H�0Wr�!3$�'w�n�$�(IaJ�/]�J_,��:)�B�6����&SS��j4k�l���k%��5nv�@�U��Izc�a�|�TUh�\݄:��J.��#ދ{l���"�2xXb�ʻ�Aq�p�j��R6��R�j�����ފCc�l��]"ɴV��q�T�5�u�OhW]w��D
K%pʚ]gm�skz���h�;��R	U��S�}n�(�<�l�8-�õ,�[�BSg�׹���&��cvʙ��4�ڕn9N���#xr��0
�c�]��c(=Dn��~^^`��r��1󲂅Kl��w���lK&�һ&S*����e�X)�mJde
��V�a��j7�(Ac7a_Z���U`���:���N8��3j���5�5�g���.�@�v�T%*�׮��O���ɰ��rV���1ug������Y�;���MP�<7V ��Hp�k3Wdoyqc��Hi���9?��c9��C�Zͫ=rB͚�0���;TDڢ��b�Y�-��拕}���4�Xvҗ[Ze���,��n�Z��^
�9��r䏫/�R�8��V0��@���[���'��ɂY�����{xl���g,�-a�����;j�h�UȒ�gY��R�\�5���{e@���Q�Sc�)�ęV����x�l��m�c�U|]��KK�uN��cu�u;k2���t2��Ow�3Om%�"B���C�i����Yu+iȹ��j[]2��	#u�VŬӷ9������hd&V#6L5!<aR���pI:Ia�fn�����ˈ�SJ �'��`--
��軺4Y�7,㽃b��iR�\%e�e���B(�feVQ	� �0٤(��[�H��f���h���4Ei$%-YI�RXF�N��:��"������Q,�wrH��qIUj<�!���!"*`��A�SL�����Eՙ*`a�bШ�����Gq����eQd�*��IT�5ICB�K$Y�ҺK�Q�I�Gċ��6b��)Ȕ35�RâJi�	ky[�b*H�Vk:�M�$�,��UJ�$뮸P��N��a�<�J2naC�VθGS�����%����u�Z����%��B����V�)C	]K�Q�a�a��_-p�$�"���$]���$�(�!uIKbh���a�H��LP52)�ܤ��J�.b�PD�L � �	�B+4�{�c�?Mpl˰�����X�����q����U�GzP�<���>�ܷ�آ����wN�ak���\��u�q�z��w�g��u�JW7��@�j}�5z�O{��^��E51�˰�7�*�=z��-�F��ӓ������ɝ����BsOz�n5��7�⸻;��ϝL�w۷V߰��7J�CK(��8JF�}8]S�x�d����R�s��ϼt���Ś[�O�ɤ}x_���X�p���ʏ�[*�--�<�7��oC�zU�\��ۃ/�C��sc{]��I�ӣ����do�_����n!��b��d|���i�D�[���7�ʚ�y\W�J�w\j#�|�+!��;�>V����W����pnh���T���grw��ӑ�ƳsH|= oN�y���Q���u�H�{�L��'E��H����%�o�{�]5��y�� �'����P�oAai���_���*�ֱ��9ģ{�<_Vhڷ��Um8��+āQ��v�ba:��D�9�Ҵ�B2��7�adG���a��yם��	93�jlyvE��~���ӳ�u�fA��5�(�����n���W����h�>�K|w$a'����O����@�8���.�9�N�c5�7�
�˻uw3�$�a���{��i�����JNZ�V���ڼ�hC�l���ǻ��7AmݷJb��ij�X	ݐ*a���l>��-j��-�WV�g(�D�ӆ*�C;AZ8����<,����1��\��'3w25!�s���~�=����C�\���d��(��u4-7-��3�v�Ҵ ŋ^��.���ޯE=��ﺐ�^v+�������c�;Fǘ��\D����r<WV/]3��W����R���>�f�����7�~��Qd_��鯽�s!���0�4$��:�GS���A�׋˴R����QB���z�2v�n#K�ʗ��^����Y>�t�vu�md�v�xmP��gV?0Еx��}�$�i(��;Lfһ'´�#==�,�O<�m��\޻.�}5}]���(��ޟGnu�\.�<b��Wq�>ë*���&����k�5�^�k�.�ݬ�~�&*~��*��@�Դw�s�W����ym�b�3�nK�zf��+�/&u�U�+�Yyy9[}�N'�{n�n{�o�G�י폽�������AC�Fȕ5X�75y�ڼhW=ȓ�����G���|9Sݮ�d�5������������a������rs����Io���i�n���%޹�aҔ�{4%��Џ���#�t���W��G;W��>��� �g؜����
��t�v��LΆ���c#��eN�����$K	��Zw�,�U�;�q�05��
eF�i:P ���oSc���;A!�98w���ڝ�)�d9�s��SǷ�c�wwR�u��k���Y�|�= r�wB�.Z&�X�:کs��/JF1���:�xv�[{c7�şGe��gç�X�0Z5%N�%x�9�r�s!�x?k�)�y�����˼r���u(>�<=����7���3ِE�f�t-�����D��O��p�������t�s����w�����$��=.j��9`��{נ<��'�~A�{�%$���Ե��~�����2}�-��5�=�p4w}5�q	�W���_��=�̀;���~��'�c\:jN�R��~�Cw]��4w�U�U�k�/O��%/��ݚ��ֽ��!���s1��o|�r�!T2�g�K�U��%��X7LQ~/J���x�0���^��2<�2\s��8��L�VfOcǕy��K$�л*�o�vQ�k����3�;^������Zn6]~�X	W�<6B�^� �b�x�f{ϒY������Չ�u1Q@N�!��;P��ŋ�٭7����A��c
<7շ�w� <��n��3���:��喅��+E���h���t�z˫x�����,l��A-�^�F���u`�`�s�n�����$��A���;L�.幀]��4���8,�p��ʍͱ�;_L���^���G>߷*�n�o3��bqF��L�4{{G)A�T��rf��Y�Y�	-�����V�]���L�y8���;Az]�:=�H^`�6��cH��*wd�e!>���u���7�}���wy3�o����w�ׯ�s�t����6���g��Ev�ux�<f◻�]���/�{�lh.�|�=d�sᑵ+��'�Xy�������=���G�p��*���Tj�����X�Z@(��޸�`Q��;��e�L�w��b3�t8׬�Z|��q�u	C���i�wK�q��ǲ�,�g�%�@�U"IH�>���B�|s�����>���ź��̍�YF}���������M�0����S�7 nx����R�W�aSO=
}Q>�����Q^�=����Q촍>�����/}@`�[��W���y�_�2e��r���Y9��s�C�=*� r9��G�n=��*����p�k�Y����6�}n�ʓ��8���=��]�Ş�}�L���&)Oi��;��|y�Lw�g��Nx�N}��][ݾ����G\j�b�3v�^N�������;~�Q��ZdV���FX���7p�x��4aG��G���0��d��g�*�����\���}4؏?A-D���[�:�waz�3Fb�ZU3Xf鮰:����VY�|��8l��Xj)��U�x��u��Օ� Ӽh1�����+�n���i�W���S�׏=�~z�1���{��u��I��^�rݹ�"[�FV�֌���P�O�}'����D���ĭ$y50�en�y>&�\�3P���uU�3�fc����w3<��q8=�;�21�y�X��A��7%�۝�^����6��>Lh�{��˪�H��oV�A���T�/U������b��碴^��t��/q���^�uq�@q+Q4�c_�#9L~����`��0�}w{I��"%ͮ���5�բ��Z/�h��Itח��뽫Im���fD���V�z�|�oO��M�>�׫��o�8�v��\$|�TW�)�|H��_�(��!������VMixN�c��З7顷ׯ��F����l�W�q{�~�w2�.^����>�p��k�(����p��`M�x�y3�ӛR���y݇]�9��Bw����9]�gG��י��W���Q���񅑱2�D�"���`Q�@ȳȭy18� $��ۼ�-y>��|w݌H��z�g��v���}�b�ڧP��!��:x�89���c}��3�Z�=��}�Y{��(�<�\{"�6r#}�=��0w����2!NQe�����$�L~�wy*u֎;ь��|�c���2s�3[I�I�V��S���w�Ƥ�)�#�޵���Q͎���v�k�����[�8�Z�d���N�v^h�쇉��k��D��ON�5"�G����w��Γ���Q�r�o�ǎ�Z�et�3?0;fx����d�n>�(�J��׭"�3Ȧw�pLE?g�C�D��*M
���@���7��n"`���P����@,-8�_��kwq��~9};Ģ��c��W�D�{g�
od�˹a��%�EE��$:`��D�S��ѧҴ�-/W�K�{���߸?R����2c�u���;>��y\�5�(�;�u�2�LM5[GY�ݾ�um�p��⓴��g�o�j��/U����9.p\@��Ty�R�g����>���q�yL�t�r���u�a#��j��t'�zd�����[�<6 �vȷrQ�X캼�[S��0�b�}�ӹ��U����������m{��q�5���̿^�,���Ptמ]��(�����"�;��4��(����K�ᔱx\��<�U�x�a���H������xg�Q�%�uϠEy�[����e��oꑐ���~�`�~ζj��q�ZU�>����M�t�:�<�'��kp�PgNg�$�����V�)�Q��Ew��:�*��3���c����������^��r9�s�y�T��q�HQ-�SG�M�"2��Ủ1.��2k#/d�Od=nU�ɴ��n3۹b�]�ٻ)�M�J���V��>��H+��q{F7(Eeq�ծ����;8_�擖of�����[�E�x��c}�*^$\y�#��Q�;C��l��`���xO\UC��R��Z��]�*�g�:�[G�Gѓ0��ӳ�����G�י�\�j���3�{E �6&Q!���s�y\��}��=y���(ڨ^7Ϯ>·ҙK~�{ �p�S���޼O��|9�RM�M��evz��%�y� ����y)�m��r��ǰzR8���=�}�[ޕvt	�wwF��A��=��T<}p������B��h��c��>�|�_
O�ي�}���I���Ty"+�ϣ�F��_�G�W���-�0a�t���V.W�d>�Y�ٻ��Jgo=���{{���2=�E�����c��+��G/��0��t��}>C���>��yR�-'������������ަ���U����d{נ;�fA���9-����I`�A\ɪ��FV��}��}��ݐ�G��˟���ί�#��v� ~�De�Qd�޹��f�wx���H����!T[��Z}��n!)|n�Q�׮l���<�}-�����/�߅��zf�/Y}��b�W;}�<�R�t��(�;	*>�������mK��T�J}��&[
���4�;�}3j�I|����U#\�D}�9g������lي��ڸٝ�+:��(�'�l�^f�Y�o-Il�4���^���y���N��wSfo������N��b]����G�%�d�����3��*8j!���ӑ'���Nׇ���>���Y��׶������������x*�w��z�؁��{��Uǽ�t��=��v�v���{��5�c��#t߰�Wy;�z����u[�5���F{%2n��"������|2��7'�RȪ����=�W��;�*��n<u�ѓ���t}�@�\CWB6�9�&�{8�y9��<���Z)̒����I���,�]�ۛ�����EX���d��o�&O:�Ə��}ޗ�g������39�B�b}'�k����g��3�l�=QP@��So�p��N|2#jW��4}�״�{��R2xE1��߳|�@W�$zx��ۍ�^�,���%���uL
<�'b7i�mN�\y�����yў�~E2��$�yY��j=i�)��^��%�]�th��d��R<MǊ�{��+�彟�v����o�vءk�v�z
Ӿ�#��#�qW�C���A;��Tcc����;ߒ�^�������Il�X���5�<#4�N��μ�(�F��u{�b����f�)�}c��R���t@/`�U�gH�t׹������'�˗=�J�4�F�gxC�����V��|��#Z�p'�ٺnW�w��
���_�veK!R�dCw�\���g�-��j�[�H�s�H����/#}�#�z�X;��P��.�T�Lw������"h�r�7�.>��E�< x]�G��6�q^����k�Y�^�z���;�1k]�U���ez���e��s�ժ"i�i���r��q��\,���ų�5�tϤ�go/�oq������,
�>%a��t�^z�ur�ȭs�=��Cvn7=�/ו޿VM��(\gb}�&=��yNO� z���5�>%iϤ��������'äֹ�g}��Ǹl���j6�|
�ٵd�o����A��7V=��EG����X��^���L6������:c��E�58�1RT=��7e7�����3��Ԝ�:��/�Eh�A<o�Z;��2�[=>�Y�˷����>��B��ڭ7����u�b�`Zs���k2'M��P�����(���~���B�U��A�e���/�kvP�+�2jN3��n�K����9�u�i�aw���g��m�mZ�u.����_ZY�T�!�R��pe����9k�ͅ��rNVQ��,��0�<�֨�k�����v�\�P��RW/�x6d��},N�_:Ri�w���F������7�>xI��!Tt�`��f���7�tFHJ�olv�@�k�1+9Q��)+c�O���p7B;4/��{zL��VV�D�鲑��=��{Gl{+Q�8JF���,���b�g_�d��hW.��8Ս�
��
�GG����G���U��~�>5���?q�߀Mo/��|�q32�!�h�ӹ=�ڨj���XϺ_�F�Ӫ=���Wh1�)��;K�Q���5���V璧����0=�V�a�>���|�=��>�x�l�xwl:�_�Í�G��a��&��Ͻmkfw1O����[7]4(�ԁ���/�\i�Wn�i���"���D�3�^��m��vK\��3��k���ٸ�,:�T(��9��X\w~�~>Ī):�����3g\ŀ�g��վ��f���Ҳ#��꜐/�g�baz��D�=�x�8�FX۟AP� ��^�v{g'�W���giLz���r'Ӑǽ�ٟID�Ih���>��MV��^mM�����\���w���n�Ln��tz��mK����������`�ϸ���}�j)�+����r��9vn����k�'C��	П^�,��@�/���^
#���D{o�xG=�ܯ�P�;u��Ժ<�@S����b�Gc6iu��U�'F��7�Z"p^>W�xE
=���E�ӛot�+:�^3��^�"CrR�F�����jp���f%�M�[�����%˭����v:�ӝ�xh=f�L�
��V�E1tqm��u�;l�������ͺʍ�5b]�}B�	�0.k.s9
��m6�0��Yo7���E�S�/V�٭��a0w�+V��U�jo,�P1���B�k-Ν�XKD�
R��*'8�t�ef��"9��Ĩ��f�~E+z{�ҡ�k�.s
#�C"�A��N��k f�Wu]Y6E��>΄�'.S�G��M8yx2�޻�^Und�XA�����:�]�p �r�}Ȃ8�oU��'h�x��J����0�$0������vuMw�[�rV�,$�r`���n�g�U�R��JX���u��]�un�ι����$_N��ov)�TE&vK5�X�'fmur/0X�d�;0��M��J�[H��B����:��lN�4�H�,�bD��G�!nq�������8�e_t��G�ݓx]�9�iK(_k�w N{�V�����3x�o�{6��gVnɼ6TzFM]�+��bNIӺ�0�j��0m�ɹ��dXp(x���o(է]%
ڃ��v_Z�x��uoz#�I�6�;zi>�ة����ə�U��6����>���vlTY�b#�2�k�d�Wu9��k���c"�.���T鐀�"�w�����I6�&��Ó_)p&���LŜ��t����=�`|�3��yݬ���2s'z�S��p��r��������U�IbJ���ф��9(Ji�a6�Y��-q3h4-=�"���q�2��v�ݓw�-(�8:�AfP�cT}+�jg0�F��7��([<�c-�/�pv:�Pew�sK�vޣf�����B3����nE�Ն����RJ*��x��r.��<M٘��X9��n\�9�q��Pc+fk�]E�x Ĭ������E�VV��W�����ַ�[�ΫN���K��څ�)�+��|��%ى���]�}A����|��a ����ʭQ�YY��Q򠫑mwg^ ���+vK�<nj|��[�K)[]L�'Lk�-C��1DcV�u��q&w^��3P�/Nv]s{�(���7��-�>��l$'SZm��d��h�I�u,/6��ɲ�9�
q��^WU�M�ϲI�v�f��v��]+�v�i-[�$r�'+��S���t��ge��Bj��t�C�f�.�V���=�7U�l�l#���K�@�Es,�jδ5N:%Y�|�ӓk�t�
�A�n���%���*�Ǚ����.^5�wk�l����*�U��2r0,]��G)�7��'����c����{�Y��d���k�����H3B�[�1�О�R�'�vZ�j`p�����1SzG	qTo-�6��k�~'���u�R�r���$Jt9�t99�ݚYr:�{�u���� �D}ȁ� ��Er�+@�$DJM%K��:E�4�m32����k1QD�f�QgN�a	iZ�*e�ӑe��Eؖ�PI
��E��:���ʢ��J�"&��E8����T�Г��4��2IL�qu%HEI���q\�<��QkS
��=F� �l�V�z�N|{/�e�;��BL�rw�!ȹ�(��S��Y	g4�3.y⮇IS(V�|묛��+�N�VS4�Ce<�:�N��$5�(4B�Ȅ�I4-�Ĳ-L�3�L�䕑�����Ȃ/!g��Ӫ�� ���Z��D�Jah�\�i�tGv��+R�#K!(��Ez���+��"����I��)W~����t�Xq�؁�HC�����N�u;z�L���wn,h�][�Iu�]z�gZ��å�����3���a�P=�[��R;�J/춿��Rok�{�Pz7�Ž̿?U�/����2+ݙ�=�~z#�r���.2���n�>9L���Nφx�{s��zX�L������W�g�/<x�$�#����>٫6,��t�W`C�������C�{ ��~h,���X�>�u��M�gK���r��"��o�K�`��^��v���rUo˰��='�Rʦ2������L�9ȸ�<zTS�}�Uo��^x��X�s��ב�y\:��;<��1f	H�D����C��~��u�N|��]粛�����ɟ3�3��Tcms��>�:�=�{=`u��lp���ZS�s�9��y��w7�^]�nϾ�������f��}p�i���R�e�p�V��j����������ly�����o�,	���y)�ojģp��ȥ�l����A��'��Њ���DzQ�z��AY�Z�5�W^�\�M��Ǚ�}D*���S랩�»p�]�f�`{����ǣ�s9��F��[�y9^��-����*5�+�a��x�~��"7�ꌭ��Y��Zf�N��,t6��Ŧ�j\��J�y�6Ĕ;�ʶ�3�vu�W�7��ɷ�/J�bQr]v��edc7]ܻ�o�vv7M]����ra��pTv�w,��n��J������u:qM�U�b֓�l��W{�z>��B����e�aE��Hy�06�
�Ah��(�Wo[:ve�Q�>�U�-̫��q��3Lz�ަ���U��m0VG�z��dn|i���FP���/ߢ]��4��v����f�ע��{���?	�����@y?��W���V�3q��3��;�ѕbgƉ�L�ݳ6��!u��5�/������٨v׮l߼�"o��>[Hx�T�y�x9+�T�E�Ԓ}�ĭ�,.77,,���3k�j#e�35��\By�9Ce֫��Q���a�e��{��z3}<n{�#��0߿Ie�#��};^�2wO��;����,����|����ѽ}��G�U�|����Ч죆=@Oi���ۈ��ye{���+Գ�h���o��tϵ��:�)��#��i�r<�_�YhP�����y��}�R��2��M���&�۾���T<��=��7��WB7:d�s��ߝhu����-��B�"��5S�n��ӽ�5�=80��,,UQ�'==�@L�O;�ֽ^��)���\w���i�̸��g�tL��]��G��\jc}u��)�q,�`s�R�f��,��v�y�^���9B�W��a�i_:{�͜d$)Er�u^	p(���-���y"���n_NX[�$;+�^��S:q��^SɮQ��OG+��OY+u��;�-��[E�l�(=�T���\;��N|6J�Sά<����}��r�����+<�T�gi�9�7�F�s�,��Q���qT����^�����ԏ�e+V���c�U�i�W�t�z7A�pz7���>�p��q�G(��%�@�U"IH�9t�5���6�;�Bͩ���%_���C��}h!��:b��P����DmE����y��X�Ѣ\����.����&­��՛��-V��v�����h[�RG#��@��}`h����Eǽ^7C��ɜ�����y��g_�l� vE�Т��%����?^���Y�W�7s�����f-�&��Qޜ>b�qs�+�E�x�M�ς�q0|=jH�s�v��=
e��*;�U^;��0"�t�7����������'.@I��>*M��4v�鎿��C����׵���2Ƽ�X��˹�.>��k��y��'��e�����,x�d�i�u\fއq���WvuAu�̋�Uջ+��ǠϾͶ��d�\/Pw�;={V=��EDy]� k�g�~Rߡ�k3��(�ot�~j�h�T��ښ��;�diպ����YOo�|h����]�&6�E��wo<r���j��U!u���Pj�Ʋ��o�E�C���+��WPU]�Wf�A|'R�Sl8��
�0��b-Q��=�V�- ��u�!�ܺ�I;�g�o/���������5��;���O�	+��g:��'>�w!?eP��C�8+��IӝM�,)����=뱞�%�NNz���<7����mV���zo:���������ck�C�6f�873'��b�R=o[��\=Cѻ�Y쉔3M�;,e�m¸�����M��W�v/W��d�/�%�H����¼<G����ۋ�y��8�O���T��2kK�w��Bsq=걳�%"�_~��Hk삇t���)���d����vym�pY)�\�=qT����c	����s�ʮy5"+X��
^��mϤo�'��{>��xo�s�w=��uj�k#ޱ�
�&Q���*n*�Ρ���>�qI�ԗV���ì��*��r���_�FF�%��z�9�Rt)��;!�u*�·o�w����P��j:�[ԉ�{���P��q�g���^��K~�ѣޯW��]9�Q��ms��_�7�7 ps��_�q�Mv�Tr5�Į*�׭#��3&w��u�jѣ�!���w"�z��^@ 7�s�Qj�Qs�s ��]O���kwN��I��{�I~�Z��@m�?;�����L�?{ݭ�<�/\.K]���|zr��Q:�$~��[v�<�#E�a۬��^w���KQ�O)0n�;�8�%E^�/!��Hɂ���]y)f�;FR�7����n�P�(�ձ%O���NT|�tޡ??���~����X*-�9 _ȴz�&��1N{�FA��:ezsm��ӝ5��i�ىaW����U!\zz�0=s�L��pq�fA��^%rZ;su�+���q<�}�r�z�,9��r�vG�1����m��� ���s�zǮ�#��P$��8�0�ҴUf)�^��K+����}KL{���K��j�8'�k�C�Q�9�ꇀV$�~�xB��U�we@4_�gGh4<���P�6����f����y���E�{��dב���:/e��]�(ˠ�ў�p�ɉ(���-7�Ӳ�x�{yU��K��:X������Mw�;L��k�)��d��9j5uF������I=��҆�Ӵ�^MiW��Zo\���e"�x�f��ǒ������=�g�Ͻ��7��+���g�_���$z�.��2�&��T5g�݋8�zGe;ʮ�˦� }�}�����x��s�2��!�����IFE�)�/	��C��^���+�e�V��d�Dn�h�ɝ�y3�ʣ��o�{�y���W�9�C��h�}��<�ȫ}X��Ә)�����ŝ�]����H�dcb�f@�Q=�&;��01�m,�া&�+tz�i��������nL=|�Q���-5]����l�tS+�h�t�"2���Ã�}<�}7�f:���4
���o���j.�tD.��v�͘���Fൗ�|7g�lv��G1\�=xe2�f��Rk"���~Ӟ)����q�;�5f�]�����{�-�
�l�*� J�:zn(�&)��7��wjĢߕG�zR57�R�Mߜx��r�wZT�s����U��2�\ <z@�u�P\�M��Ǚ�}D/�{�p�k�Mmu,�-]��rY��<��ߣ�a�~�d{E˓�fF�0a*���A+�a���׵�\U�y��������}��w�v�zg�A{�H�ȍ��=�[�jD-0az��BϏ�Ǟ����c�k�t�l�.�߁��{ԑ���*����`��z�~WLS��R
tl*Ƅ�<
ƫ��Ң�M�Y����di��1?S��7��=�L<<��p���_�D:� �����+��尧o�Yc�z/6�&�X[fl1ٲB�Vɨ�����T�rf��*�8L���e�o�ФO��}>�X�3�.&XH�M�
�6�;��񚍗�ɯ�K9�컅6,�
B���~�F��ry@]��F�Q��ǹ�O��۸��p߿Ie��>gN/�����k�o�%�b��7�b*QzBW;b�����᳛K�k��!�V_���6zӫG�薔�������ea�3Kk�`�}Z��y�wU�T	��Y�>�#��yؑw�L����\���;2�fV�R2�����k��!��0S�q�[$�ђbK�)U��ѕ�r�Eߴ��ր��<�ǆ�q�#ʋ5��*�_��tǐ��Ih���C��~73�x�&���һ�%v�i��U��l
�V�$?d�'�to���'��Wq��S�.��H\���k3Շ/�Q�rvcێ���5�5t#s�2W�uk)9���Ϸ#}���^���}��u(yF�t�,��Q��F+�xN�{�>����wq�z��>�K�}�JZ7X`���}#�i��۸��5�QY�$����@��Sb���e9��ڕ�y��c����������o�O��_�G}���ݪ��j�+#d	F����T���^�d�ٴ3=M7�=}=~�Ύ�++�6wk��>G8�9�u~��d)��l�/2� 7�Shw�� �N�+���޴�f|��>���#�d*�y��B�{����J������~�dxd)�� 78�o��F�P<���%�m_Lɂ�	7��'��1��T��fßKg��*���uH�hU�wCӜ���t��}�G��́�j"�Ш/��r	h��5���n����p�k�^�U����Ȓ����A�ݺ���'�xK"U;7���/���N�]V2H���.��K�)����'�~~>��m���#E���UՔ����C�ѱ��j4þ͝t0`������$�ʶ�|�e;[�y����G�&�N�ӑq�u>`�we�Vꜩ92��s�TZ�&���ρ~;�!L�7��\.��蒙C6;(�Ej����]�|�sƤߔ��#����,�h���q��E��#~~��Dh��2�^B�4W��G�1�7l�m�W��_��yIf�{��$ל����#�ud���:����!vMz����W�t�}��`��!���I��Ǿ�:	O��Bz����	Xn$�:��k��"���[=��b8Ю�I�@~��fj/m�)+��b�QjNG����
���љudFP�f=��[�[�h�ޙ�,����^�_�{�=�LBo��S��vi�E���~��Ld�ڲ����!?��O8e��<0?Y������x�X�h��F�_�/�q�s8ˁ�Uu��6�YR���i�wTw���ݶx�?c#t�+V�o��V�KK?*��C��anI�T'���%���	J���~/�G�{��=�(�Qe���s���"�X�p�@0�����v:;�5umt�#�Xw=��O�p(��y���W��:�q��m�Y�2�I�*c�w��5�VFѡ�Tm���YR�����+л'O���}Ϭ��B�6��t��ω��[�����=��(C�i[�b^�zn	p��崬]�X{�	�qL��|%%�j����2���L��z�%Yɮ�05�n�Q:u����P�}[]O���z*7\$�c[�2i]?��f�w씷*z���3���f���+�|4��A�G�F��s"}�o}��)�܌�^g�A(�a@ȯz�8����P��q�g����D�wf������w��@��׾��B����U\��t���B�t���h�q��,�S���r��ǯQS^���<�DxY�}���߯FG�}%� 4��`��L�ϑ�Nd.���	:}�8{����q^����A���{�4������$��\���Z�&����v��tn+�[�����TR~\�%��O?g�ؙU�������{ِj�פ�s�-����po)ϲ�?O�Ǳ\��Lz�iQ�r��G��p�\�ߪ�G��t��������w��γ�yn���þ�n�ۓ�a[����O�����	���s�@�Yn�xmg��mj���������C�{��%���X�3c�7���k�n8�&j/n��y���E�S^򩀄�F�U�oGo��8,�s.�{(�h����T챗���뜮����Q�z���W�W�::���?а���57��t��V�,��Fj7����(2�tFQ����u�e
����^,�MG�SOv�����	���:���Ԃ*-�L����-9�<����꾐Vp��f�/l-W+��kt�s�YY����T��֖��lʏ����ў���yR���'}�gM��$��s�CN��U�^O�iG�ޙ+�]-��[г�_���,�~�p��ǁ�z���b��}�x����}�VESc�=�� (�/����VgG��FL���R��k�c�U{ċ���<�to}��b���W��^���F��(܈~m����LmR��YY��+2�!�*?����j�x�{)��Whh�f��'}�̜�K��ځ��g�dK���Rf]�q�PW��x��뇟qu�9�L�
����'g�c=N�]=�Hr8\�Ss�Y�r��<zn(�&)��7��v��J7�;~Y��ĸ�E�QKЏ"sק������N�7�� ��= r��]
��h���<�ؗ�����	�������o���B��M�}�U����k����Y��,_�d@��R�6h�~����ɾK��[�v}�W�w��~�hU�v�X�~�g�4���������`�ƿ����!ŒjӍ��c��]i11���%����:����&Y��=�ށn���cm���m���l���m��l�A������6�덶m��l��m�cm��m�cm���`���������m�o�����l�{������cm�o���6�鍶m��l��6�1�� �`���6�1����
�2��LB���~�������>�������s�UEP�� ( %  J�@	T�J � @J��@QUB�(�� �
U	�:(P*��H�J�QBP� *$J��QR��RhjI ���!F�URH*�H!6�(` 78uDUT*�R)R��PURIEDP����*��@*J�Uvb!)ED� �REQ/��P$
�� h����HcU�)�kjjD��*@U�kb���md Z��j�T�0Ɋ��H��1EP(G    �8�@)Ud`PЍMP,��J)E�QnM�(Q@t�����8�E�R���E(��ݎ
(G�R��T$@�  ӹ DF���ɪ�ն��Uf2�
��b��l0IM( �`(�mU6�Y*�(��i*�� 8R���)�R���@Pԑ1�hTʛM�f�m��ڱ3mmSmU�`f*�hҦZ��5Um,�D$H�Q)C�  �]U�m�P��eRUC2�j&���l�L��lf�k3j��df��Ŋ���2��cjZ��քf�j�U���%*�LdAH�H)J����  �]��Umm���j�f�U�MZ5���Ͳ�F�Y�b34����	Lض��JڬkR�ѱR�[-l�+R6�U2	$���($(�p  !ʝ�k5�hUiQ��j-�l�ZM[[[e��h	�F��ʥ
�@��V�MZ������F�0k 6��KP1) � P�p ��f[D�m)���)Y���ڵYZ �ٍU2�Re�LT+XZZ5T�V��e�����%U��e�UQ��ZB�APP(��  w%�m-m�����Ucm��KKf�m+m�l�Z�R�m�ҭ�	m�F�S�ij�&��fih��kVkY��P��ER)���p  ]���Z�bV�UMh1�թ
Vڛ#fm[*�ʕF�R�SV�ZZV���MF�l,���&�j1��  � Lh2��(a4b` 0F�S�R��CF�b�4F���M �ddL�z&���F1O5!�J���&0	��i�L!�0	����L&i��M$D�UI       N�������/}�8\��+l������L2�D�z�Z�(���EDQ�~�2#P@A7�"�4S�B
��Abq�?͏��R~�C��A����b� ���p� �B1VE�r�}ӝ�U��.�N��(�7��KK:a��b`;�O;�e�A@~������_�R�X9W�U�ibͬB��qj�;B�w�$:��,�RB&��Ӿ��J����Vu�V��@�)6�,�]�mʚ��@n�����a�mn7L{�Th�u�v����^ø�S�J��UAJ�f�/]�0����9��<81��fG�2c�67y���u1�P�i�a41{Cֻ�.�ɚ���w���J�i�PA��j��#C^סU"�[E�sS��!�`U���4�3��T#	
�uBH�O	D�!�k*��|��V��*|mCWg6<fm7gtG��B:,�eÎ�$�EjT�'ţ56�&fa@㠖�YD����j�������vŀ֗���!��m��F?��P���x$�@֫��A7����9�h+��[��s1�mr�u��>B�o
0�� ��ky������WX����p�Ո~�5
��-�� O���vɆ�6v�wiO��+4�j*�<�kqU�'�t�S��ޭĖV C����1�O4����`RO�ռ
�.�ȃ���g�����%A	h�e,:Ue
�O4}3h�.�C�%�ó+X���MY���-��nb�Ƙ��T�-!����=���v\&���E�q\8�u���,��f䖩���u���=o�V��u�|ic�=53�Y��`�k,lvwFPr
�ZZ>�[*E{@���	��^-����#sy�x�����ݶyPӸs�M��ӻ�si������i��Z6�v.��)�p�N�%F��p;�2 ��e�T
�e[i�xYDY�Qws6�uAn峃�
���6����m`���t���{e7L�2�j{��;(/����GK_�m(D��ۧI�h���ߝ�>.���E2V]A�h| ��J8��w�&S��U��������Ҽ�����+h��.e�l����L:�q�^TZ�;;C32��%�M!V=�:����#�Ԃ�gc[ذ��J��E�ݺi`Wb���S76@��\x�'U	yN���KZ�en]�U�� �n 渲�a¢�VN���\�'qi�SK�b�.7�9%˘�^��C[�^K�Z���f)���9�p&ef\�-d��KZ���j�(o�Ĕ���N�tQ��8JK{yn�y�6��HkԞ,� \��JI �ӷ�ި����WM�[`)w�@(�O7C�=�Wsh@%C���7P]5�;�Z�~�Nm�,�1��w��.�JDm��34�S
V�W%ٸvQ�2��M8���񶐬54�����u`*���q4ј�0e޳��q�i�Kpv��kCK�0�r{���D���m$6�&�]�oQ��&oX,n�l٧Nd;�.�k[��1elz��kGDM�2e�dͼ;`�	�!��C0�i-
���ʱWP�ăW�
�d������pvb���M��W� he�?�Kw������69Q�z�V����z+Z_����;�s¹��7�	^5X�z����wsO�K¸�Sc�f�J�HU��:�Ԧ2��ض,n���2���V0ƭYw���fX����N����@J�
���^E�Nfk�6�7���y$��ه&�ϑ4۱��W�A5w�z�E�KB�3n�	pkߤ���op�1ʽʼ��aq�v)ۊࣂ�ۢQ曶�t�p�a�ٖ*�J(`�R�mmZ���)��*ܠ��iX��2�P�@��5	��r��
���<r�Ĕ��2�ܠ���K��	�᫉*������Ht�N�3+v�Ŏ��/jd�w�XU1�!c\l�6t�{s̺)�[����gp�
�Ȯ�*]�BYl�حFq��b��i�c[ab��iWa�v#�?r���B:�Z!J�P�`S�S��n���e����2-e�j�u�E`O-�N����\N��WN�1��D�p�Z�pY0����,G��޶3>1T�K�R����N�c9�"Gy�+y��U���8Y�E����L ]���F@����J�Fe�J�H��a"C�VGSE�2Φ�����fO���oRy�$ͬ����af��z��{��j����?<���� ���Oϕ�ʶu� M��Ȇ�e�H�`X���p��GVN���g�uk,M5OMm&s2M���xw���0�n�#M�!eҙ�*�h�a���V��r�ЊW��k-قl+EH5�߮��Ki�8�[�75(�Hj]�%]���d��XLiƲ��v̺����R�k�H/�r�,��Z�N�Gs/%9�eb��^P����v%��`�]�$�PZM���-��d�{�Ǝ&��zC���ެ:Q��MM��6hb��m;p�oH�o.����+q�ӓ1�'c`�����A�L\Ī�X��@*�a��XN���u�2*�0���*�V�.DQ���Aߵ��.Q��?���yr��ywIc�U��Y3�����5�+J��ݝ�m�E��]�W�H,,4�7�1�_"u��ѻ7�Y������Kov=��Zp��5�G���t�Ee֞��nƮ�_:�6Ooo+1�f��$jY�07���Z)�5aPG�����ɣ�6�}ڎ�Hu�P-]X�m��Vì��Cjc��w�2l�@u֛�
�D�I-jJ�6ԑ;wa�ݬ:棶�%a#���+;a��O��[Z�IRm5XC4ZI�/tř�,7S]�����j��DgV<9��Op+H66�}�)�KJxRK{E,�h%���]��tN�#�5�/8il�C��]�7���,�Yjǌ����M�YGT��f%[t�@d`��Q�oe��^5��*%2��w�v�:����E�=�;���;6�}�E*�#�@��
��wϒ�ƒ�f�U����F]5��cԲ��
�f��x�Sn]]ӕ[ݠb�7*!�*�$]��nf�J�?+{���X�:��l�j�ąiV�-5���1���<�f���w `�-���I�iFn���	�R(���J��6a@dJ�ټw���6J�V-��ڦC �y����,-�W|��h��Y*����K)a��Ʀ�(��FJ�c&Juu,��7��C��f���^dʧ��x�$�/*[G�D-���ɚM7z34n�7j�Xr�$�p�j�Ҕ����y&�D�˔%Ѵ,�X/��ł�Z!�vI���ur���+fn�÷�T��y��[��aج͔eۃ.�kC��"f�;��j��57!�8Z�X�=��*fI��I�m�aci�j�9�hPzDrVr!lD/p��Z�5��q�i�kXj�f8h�.�R{�鎥�Օ�&-*�GQ�X��u����GN��)��ѽ8^�!db���xi-��������T��K�*�F�ܨ�.�=���*f��s%c�YH� �'qI
e�ŗt&�����e*Fn�ESqm�b�K%L��V��7v,�ݭ�n�	UlH���b�5&��.�������0�����ҧգo�@ �y�Cz�b�]��6)����K�TnT��Վ5�MhyVԚF^Zb�p�����|��)�Q�A+%�7w��M[kVә�6�D��靎�a�$9�H-��+v�c��Ľ���Skb��Ɔ�.�U��;6�ԕ�RQ�T.��e���r�scm�j�*� Y�Y�t4fhj���I���	�6DB��6�n'n�5�,�iDXώ����V0�+"��Q�Y�"lI�:[�єc��=�-@��������g��Cᨴ�l�{����n�ٵB��Sf�ŀ�ɛY�,,)Ҳo$�-��V!ű�P�vK`]��� �6��;�M�Vgh)��e#Ɗ��P*��#Xf�r��X�m��3gוj
�:�<n���y��OcX�5��Wx�ˡ���6��D7,�����&����U��)U�J�Q��V���ب�϶��l������K��&�݉m�&�.�ę��ګG�RG)��=�򍬢�#W��dkV\� �si�ac���۳4�fMVihۤ�Z�׎Y�OF�hڭy��P��	�*��F+�ChT\7�c�����yt�� �K`/T91CwD��mz~%K�nj�+غHɢnT�VZ�$'\�4
��x�/�л��ԋ�}OR���p-Y��ĭ�3E���W���jPM�wO?�M�D�[l�����7n l]�R�8h`Tkl��1��!�ۄ�F�p�jt��`-�f�M�����Ј�4���^�cM��h��f:nh�S�O�6��֖"�F*x�
�J;�S
쾻���
��={o��$û����2�XKr��o6���.�i�9�[��<�5Qyt�\t�Bi)�N�n	�rJ�n^���Ʌ��۩VY݂������P͙�f)KӄX�Y�N��P�:e���-.|���	�Z��Cj��iD����Ԣ`8r�B2�l�۷��Y+/.�Y76HD�[��"��;5�h��e�����oe�WM|/�gt�.�M;x��h�3j�T�tf�X�:�ͬ�uп�*n"�ѵ�f����s�uW���5<��n����� _,J4��1��q[�c�/p���U>�!�)�q�y��h6.��`�젎_A�
&�W�<ۍ� ��`\���m]�����f��U���DP;����)�:�fe�輡yT�7J,zƣ��?��Z����S1q7��&��Fho2�cum��l�(5o,զ�'r�vȀ!���)2�)��f�oi|�r$���q/�:}�P���It�o3>-�
B�{v�+�	4���y{�[�b��Qfl�W3q��$�Ar�2�Ӕ�'�*Ւ�9t�;1!���( �lǿ��+v���e:��Wme�A���\�pF �N�� �Ab�.�F�J�o�����^� �ʬXM�Oj�6��C.dB^�Uy*[��n֫�B�����Ȣ�h6�q��hnlъ�!�U�:K��Z&�r8�m�$;X �n���l=�`K�&�ڰՉ����N�c��U�����=��+h���.�4��C���M� ��LH�������8V�Vu5�1��B�V=߅����̬�����5��1��-]�Cv��Z�ऍ=�A'Gα)�̻8$��o(\Ym�Ə�=���]�4���6�kY���(�g��Aܬ���HC�e��1�{Y��VPF2Tyyc)L�U,�,�مſ	�)��)�Cu{�����U���-�	�p�0��,Q�^�b)���t�`�1ʂ�����ԫ�F�yoF4n@�"�Zb��ڒ��C5�٭���x5��7���oaTq��.� ���E�u�
����H�=J�nʺ[��zb�	�Y-��P�;�<��q����M�\Wu��m�^m4dǃw`�f$J���a���J9���/U[����S�Bb���$�;0l	`���ӱ�:Q���dZ�̨�gE0+�
��b"��2��U�ih6���3�G8�e�����kh�/1�F�YG5���5���zu��;��_%�l��r��;B��[x��FӇ)Q°#�n���Tt47b��+$�`(LJRC��Y�(!�Dݩ��v�%]�.3�`�̣xj�oְ-���ޙ1
	���1�s0Z:NloRP[�Y�����ncɘ�i଺Su�I����i��̩Rʢ֒�#��u�
C ���Xs	o(jw�i�n���1W��р�й-�G6��c-:/��'�����\�*��Z���zk����H_`Zx[�q�k,�ǙY,�"X�4�Dk;��+x5�%�Xi��o����q�D�D��nl�k7A�&��.VU��n袠�h-Ӓ2m��mD���d;Ws��K�4CW����0�[�ɣ��w^V�
@�n�ŀM�4�o�^�ݦ�A1WY���^bIe��ы�V�z���i4g�֥�B�ڽɯS-m��r54j�Q�,l��6��L)Ze/�:�ܬ�(��ef��
��b�!�%V�%��M�\o,7�l�'����]@�7������̺225�2���c"��8���ڗ�˗M �N��y�u�UL`���2�"+2l��l6j�l2���,�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�JI$�K�͍H7�d��*|�׸)��jHwu��gP��mkܼ�$��kN"J��V"R��j=�Uw�x6i=p급b�-D�:��T^v�$����EQ�@=o:q��H�fV,YZ͛d@��ĵ���	����i\��И�Sw��ݼw7��F.�m��_E���CinR�o�pT;�\�k]c�K�-��.����f��&t�K�Ն��=���^��{�}�w�.k�s<wWH>���,j������1��aT+*۠�`I]{�n�9��#Ek��CV;d��E8�����u���2�k�f��ѫ|��r��,�IU�'m�Ǥ|��ك���{7e�5)�ώ+�w�!����P�L�7�>�u��_r'k���"��Y�7�s᎚��F�ؘ6�?��ϸ��ձlq�|6�;�">��i��+ۚ����<���8򒸪V�5��L��mdy#�YGfQ˂�"�m����*�b���bC��k���T�ݩ]�Q�8S=�/1os仅#�h��]��(�Ѯ��y/c\�mc�VmITft���N� �5�$jӮ�	$�#³�M���B�\��q��w\���2��x:��ȁtәt�`�4����`ţ����K�o|f.C��,�]yGm���YfF>��-�.�et��j�2{jnšحα����&�d���nu�������ir��.?L�k��.���c��koR+"}P�%�=k
2�N��:i�G{�����KkC|)KVo�[�f�j��V�TJn�W\u�3c����ʵ�:�ǥ*$f�����ڛp�Xjj��e��(	� �հ���÷ʱX�T3ۍMӪS�9U��ܰ��U�hJʄL�9�W4�@X���$�Xܳ4����]v6�(��}ֺ�(P�N��w#�MH��UmXI������F:h��~�nXz�ɼ��8�Ƿ���-D\l|3l�1.F��YY���<㽑�X�� ����b�8k�*.����b�fF�C���'ՇJ�V�h��x���5t�mf�J	��4��L���J�}�A�r��`+�6u'�b.�XY�3B�����9��MĲP��]��NR��p�3;  '����R�≻�:����с3W(c)�7FFy���X�U,�%��ؘ���Ģ1�t!�뛶*V�#��E��`op�h��N��\Kuۓ:�,:��;J ;���;�99�3Y�+u��3��ǭ�Z���X�*��՛\o@�_*��f��Z��4uu�0��P:�D�Wcc��c�u����p��簋�G�,����.Nw	�Wd�\��RJ}o�I��uj.��Y���:�R���R&fھ�i�5WG.��[�/KD]�X�;<�L.�Z��9�\�����s3���x뺬�A�PۭnZ�µ3�J��^T�`���=�0��%�]>��T�R���5y3QJ�<��3`��$��$�,>a:�P�9�B�{Wv*�	Ւ\߶�u:f��#��!��"+bΘ�K�h�܈YU9ʱ�;V���Y�\ނ�8l\�8�6z�᫝u�뺘�`솭t݌}�)՞�@:�6�Σ�Zw�� �O{`��ْ���c�s���k���r`����J�-u�I�޻.�"չ�Ysf�Ʊ�4�\�����
�Z+Ŕ�7���כ�����kjw+$v�
��D�N�*�J��w_I�7�x�sv��>Ń��i�D�Y��W\�ږ:/���t���g��^�C��М�v����ߥ�R�����]�\/�7�+s�Y6Z��ok�io�rb�;��C�����D� ;;�Xdqz��ǹc]����`v��vk|�&����N���S����Gpk����K�v��֗J�:�h�vE#y�X��:�JJ�,Jy�"��]X�3y���2R����}]&t�ƕ
�'E����>�}p�W��ՙ�W_WE�)�ni�ݲ��f�ky����,�kmj����eh����f�s��*=���ࠂ*��O��&�J{���A�.Wd�:���LS�L�3"5��"f�o:g�C�VK�䡰Hӹ+��w����R�L,�A�qP��&ƞ\�4-�[ّd�fǬL�y�,��dP�єX̗ye��9�SF����^�b��ت1Gmuj�N9ԫH�o��;@f�Wڈ�&7�����M�A�����"�KX �4fA��:�N�QC��[��r9��Y�t����۩�s��[뇰	tL�t��'��#p"bx�O�Wf��G't���a���hr���:�uj���3.���۟e�b���X��ٖ�u>Bm�=�h�����VE�9��Ĳ�ݘ�5�C9Z] ���F��j�Qn�p f������+�5	����ڎk�]�{�.�l��VF��űyd�Q��y�b{w0��vNv:����D��S+����ԑ�Fov�T�J�K�ˎ���X�H�5�⠾۩0a2�V��@�3�N�e�#�n,躽葹��W��E�ʑJ�pY:H�m<{�[�HAUڥ	�+(卢�ʮ��ӰrD='�����b�v�+1A���@.	��}��)ќ�&t�2�{3d���[��1����8u���,YeZg��\�I��Y{�;�t&�{{�p�=��v3��֯�RP��Ũ틼Ĕu���S��=z�du�9�M�Wݯ�#��6��QG)*�+��uʾކ!�ϛ�i5�hǺ�U��Z˸��Ti�\M�Tb����a"�b�W����Jo�q��*��kZ�԰�@��G�{*RSf,$ܡu��F�L�����j;\�L;����Ԯ��[�f�i�Q�wիa����J˝d�:������y6х���f4;f��s��*��[��]���z��`�uz1�w�������<m,d������սA�&��;�D;���aa���BX��w"��2�v�;i�xNh�\M�l�ٓ��〵�;s�F�o���R�Jg�}�A759����s��0h������B��Z&+92#þ���Uz�w��*7%o�nQYFM:q��cU;>wX%5���M��Sv������V㺅���*S �k�x�r�5m�E]�#|�Jo+��T9�<y�ٝHL�}�^D��e�Y֨�a:-���m2�f�Uh�V��	:�1{P˓n��V(�8���DU�v^溁V��h�ɸ��F��ͅ�k�T�t8�l'7Z��*���=�:���*�ݱ��V��Q�㌮�Ǭ�4�tM���v��oM��H����QJ��^VYє�Y����h���3n��CJ��6$r)�ݬtm�n �s���5�l,k(A[�:-���8���f�޲q����8(�y{@���$�t�Pu��ܼm��)ݢ�͈=w�E���}w��ѻ\��Y�l���M��tjei���y� S��]��Iv�]��]�K^Z��oV���&U��`Fʶ��jHFH���#�;&�a�j�ȞD��F���v��h̐����ئ�l�)C�!����ٖ��C��l�۾�䉝�$K��y�BmݮP���7Y1�>2P�.��>�ty�im��3%����:�n���a�t��>f�jsF3igTɔ�#��t��[7�7G$`��م�j t�	V�N�"�pO�ߍ�1���9.���
��2��Ή܎���1j�KV�7:h�׷r�.�0�Shn����a(,�%�Lgѽ̡}��G����u�D��_:ܴܽ��[9UI%d�n*�>�C��N��U�gF���؟b��T�zw��m�%[(�ؾ6�W{pf�3z���Y�h�h�������J�'�S�w��F�P�^����p�
��Yx���3eZ6� *h��Z�Ž��:R�g9��kR�4��l:/k
-�s�C�����ҥ���a�<�b4��FHZź7X�ǅ����:���㕵�KH��i�o-����=ү~���'N#��]��M#�F��cc���'�7�C�D�8s��B�"�g^;�ub��PK�b5H"���*�DِhL�9U�ĬF�;BT������R���W�W�:��m�-d*ڏ�e<�d��)� x�d�5M���{-��/e���ZW��Z�YЀ`�/0�S� ��(4j�����{и@��R���b�� �ZY�9�}uee+�d<��ؠ�.-�O������z�v��ft�˚�hʕ��0��z�t�=��ۃ��m��*�qդ^�gZt�.j﷛���skr�v��ڨ�B�!0��gn�7r�K�3�]�Ԭ�t�R�T��K/���RN�R8Z�w��l��q1-v��-��9��p�+���)¦fH{:�&M�����&��r���o�A�i�m���%Gm��<���z�.���ŧ�H��Ln�K|Lt���BU�\�+ԥ�N��t����ޱ�X���m����d��m \�{pZ�G/�q�a5��جH�䙿K�YH��W5�r�X7���`:�4��x��s;s!�sw1l�f��نkq��D�Z�k(t30�-��v�ҁԠ��1��O�[��,f�^N��ʼpig���,M�bR�u�أʢ��8��s�8{�����)R�f�[��xb.�seaP��L���T��Ք�s��� ����Vi��	���طp�>֞5�b߆V>���+�Ж���k5ޱ�
뮾rW
Tk�6:>����4JC����γ|<��i�����a�t��Ս����R�����ΧEƷN�<jS�}-)�S&�z��n�uy�S(8�+2T�y�D�����5�7�����SK�u#�R8�&���T����l�b3�Νf*��Y�p���0J�Vf��t�sySK������8�j�s�v�_D#�ѽcfl�P}�����2�U\�Ow7��K x��DR������9O;�Y��in�We�Xq���&��`TF��s-�\]^G�d���s���o |�"6��:;>p�O����p�]��K�n�w$׼9,.޵�n�uf�8p���L=>�2J�Ԯ��[5j:���7Zu���|ݻ��ʽ)ֹ���� �YsAF]��ࣹ$ݖ�d �xWv�2�C��飬��~�f��V��q#,ލ��e��8��Y�3[aج���aO�����ke^̜�����t���e���p��t���r��ZzJ��I�V��+�)v-���&޲w��~{c^��Ev<�ʜ�v��a��yC&�f���_
�9=��,l���(n�s(<ϥ$�J2�Yw��x]�.te��α\.�&dy����NʂWbi��z�5��Q�n��#��U�&jΙo�b�jH�)�b�_���<ܘ��ν׳>�L�f��;ђٛ�>���Rmf������VT��B�E�[ݛ�7�1"\�Vv��G��0���cZ�]��J1��z Ś�`�n�=	33i!X�"� ŭ���u7v��(�im�;����]�E�N�$7z ̨�*�q���lS��S�1T)��<Ea�Y*�gNTr�g=�	��.α�E�r%-�J�9oc�}�$T��v��|�r�r��]���xf�jE|��#�p�6��Nأ1G�u���skpv\ӓX��S���4JHj$JH���:P�w;TYʑ���t�]��s�?�v8=�5k�KR�.j�,�g>��t��S;
zY��Z�W�v���&0�rwr��_M���N%Fl�+b{܃c%q�N��G�UK�/�}/o��#.I ���+�O#�rE&�p��!�{c��gM��\���0�J�L;x���j��:��#��5*SQ��Q�ՎE$�ēR�����bގA�<9ħ(^i�\����9kf�'&���$�I$�I$�I$�I$�w��c�[�p��`��r8�Mʹ�ζ��u69	�Դ���ّ'��Ƭ�ҹB�SޣQl��WS��twO=Ms���u����S�]uD�gnq}�.1�-E����jI$�I$�I%�o��O����?��?H�������$�SU�^�DEua����2;����(�;�q8e�_
�mRֶ�+��
Ӹ�O�z{�*9f�cz�s�>�2F]�32�M�`˶D,,�/C�,;Χ+��6T��}�|f�-X��V�w���-ѠDo5��1)K�����.t�Ya��.��\�&��K�Z���G�;ݫ�p�.7�sD��a"ki�Y9.Z乑��L�-�:��q�*ˌbv�|麎���=91n��]�yb�C3�Ed��ye:m��N��n�ye�O�	��u����
{Y�P؈��G)�X5���<��[�4A6���Gkm�]�������g6tH�U��A���.9��{�셭6�n��]�j��'��@n'�]��s|���xV���(\r��1����菹�7tչZ������V�w��"n�����+{{�2M�o�t1J]b�}8���&v��W�w��"�"���P�L��GJ[X�=@[��s��r�_�oׄ��:xF�`w0#��w��mSKhGW8���v�8Q�����:��E��&��t�1v[�Leb���Vi'7w��4rR��*�s���,��L�\Oa�G�ܑ�ÎP���Tu���/U�|��̣�B���\U����^p���A
���z�<�ڴ`X��_;5�ק"T�N��YM�VAx���a��X�os�(D�zԣ��;�j`%�����%��t�Vա�K��n��7w>:��m��)�}����L�q*6+Vй��L����]ۭ��V��r\6E� 5r�wԺ�-�w�V��:<~�݋Q��8y�^X2�z�̷%����8%5yh��)]C)p;�5V�pHF\�����l��6��{����(6Ӿ��Z�����dr��z��T����P�
���p춍$����,;N�C3�N>����5N��m"Uor�M��"��N�7C�u{nv��N`$��s�^Iۢ��+&tK>\NJ�����˩y�Zvɑ����j��H.�"���p��	/��]\�`kC��*Ӣ�9��(jJ.�f�\������P�����ܬlm+C��\�P�nu;W�gL�-��l�զ͎��U��Z�L�%5�5��w^&=W&d	��\I��\�-�xn��q��S
�X�4ػ'7-�=�檀�/5Q:X0�*t+M힕��q��3a��zѬF%(E��C}Y�:�y�k:�w�j��k�k��֛)����p�N�%]��J28<��;ò[���`��l�2��ӽpӮ)�+f�Y�{4i�McH��pq<΃�Z�7y6���5�M����]�b�(RW,\�۹�zgn��T1+=��^�ܒV�I��HǄ)9�,�/��t����U�}b�Z����Е�eV�Kf��[��Σ�M*-3.���,����ï1[���y��Ø����[Q�*��Z�㸐��{��m�4c_L���EMq��8Um�J�ɉ������oG����x�6�&]���f�Õ�Ğša[�M���͵}���y�saa.w�.����[4\E�8]�\1d�FM饾��7��Qf���L�j���&��0���=��X�X�j����ʷL��]Q=N�;.�p���W�
�AJ�6��j聰�;َ�&��s�����v��(�/�x5Xk/��Y�c뽨2��Er�x[X�*#6��4`ߒ��ڭ
���y��aμ��vm�b<$2u�,�Գ�:̎�n�v�ΙJ]I.%zx�Ȫ"m����Ϸ
jΗK������D-�oz7R�Wjk�7b��vLy���:��RPS��z�d���r�Z(�r����rԵ(�W5ʻ���R6����iq���T����:�{d�'O��(v�0X��y	»��}fnm�x@=�7�4;t��B�Gl'[�(4��Nxi]q7���2"���œ0U؛[��{���`J��D��fʋ��h�C��w'*���9�ͬ�L�"$n���|"2�Q�j{�eg<">�Q^�)�4���e���M��-�a��6��m����꾬L��0P�%YZ�M%=���7�I@�kη���\ ����{J�{h�7ki�c���&�w�ي� ]�]9��\����DZ1��f�U�*�J�;���u����>f�v� +��j��^�F�-ҪDU�ء�w�;�.�@�T���#1<V��;��.ӆl��H��Qp��8%��a}|F������&�8Un��J��k6��)6�,z������,���92j��I�>�utCWĝ��|_+PT/;n��j.Wg.�6� �/�­�qu�t��Yrt�^�&���^�C�WlK���:����1��-T��Wr��zN�
�;C�.�؈�R�nf���r�3�1��4��Z����^�w��5����w��`���I6���9\�y������y�������dJu^[X4*��U�n1[�tN��>��@Z� �:I'������,���H��"sS?+�Z�C��@�s@r�x��DT�;�W�ﲐ��Ɍ��p�|�q��f��ݠ���}�Y�:ob�N��g�6w :�-5�A43E�YVj[�o��s�ْ�f�P9�+R1��7�ܹ{{]PV�8V�����#�)�����T�h�)-��n�kX D�-F��}΀�Eh���!G�)�>�4��"6v�rŦM�cd�c��1f<z��8���.��.���C��:����tk/�Ѿ`�nZŊ6'��-3TR����ii֥�9}������kd੺V;6ws��XzX��e5���[צ�V�5���=2Z���Y�L���@�d��=
�Օ��TjT�Et�Z;V�HS]R�����j�ۼ߬�~�;\���h�w�<q�gi���
�W��S���e�6�=8:"n a[�T�ii�\���Q���[���z_�D��1��尦�X���w����k�н�WAmn�s;$�C��h��T�0��J��@5�;�ۘ^;8c3��3eŌ�:���ά�`��7�OX$�C��4��R��N�iS�](��R�����EI��ZZ�[i�o�Ȇ�����2�Q����=��l��+�`hS�q��	2�B�7�S@�M��|E�D��-���A���qJ�jd��3����W>���m�n�̺ӱ>��ބ���-�x��Q�+j���)Q�_	�l����/�lm
I�_.�}Z�WpH,C)�VWHl�L���vw��w�v-,䁼�It-�ܧ.6넼'���U�\T�[�s�QdNi��+$�I�E]6�b�)h��J�6�\�N�ց����島���Mb���:*[����Z����e^Q;vp��n�f��#;�η>���=���(EG�fZ&C�F�%(�ὔ�]�I�f��V^��u2�"�[]�w7(�$ô^���=kY֘w]V�]�g��G�ǀ��N�5t �	K{C�4�H^Ś*ރ��|�M҆���+��3 ��=�/k�I갬��3)݄K[4n��ok8���
Oh��Ԏ��D]�(��V[άJ���9>?qʾۧ�(����t�.G՗J�=q1|����1e��a���F�v�=�N��x��Նkkεq�qi�hC���}��M����� ���4.{}|s)�ҢOlTPn��D�G9�B���;�F�6���:�3y�*YSTƹ^�6�[v�hũ�}��Y��뎷	N	S�<+(n�3�6N����
E�r�N������r�ro�)j-
#ZD�:�:�Yu���h̵�-s�{� �-I�&t��F�t�맊���4"�_ש����o#��7WMB��d뚶�{D0���v���Wj���D6�N�|r��F7;*�䬋��(Ӯ��n�v�9�����tOH�[b7��s�t�&e������בu�ӹ3�n��M�yƚ�L�F�����j�\�)pI�<B)��;�!H��W��]�6I'e 6��ݩ,Zŏ!�L=ѝ��y��W/%>s@Z�Nr��ט��{`*kt�죔��v�'bc����L%������n�p� ��-���Y*�	��r!�������%a:�Ι��u
nM*��&�z�ŀ�\ͳ{��ٖ���&���;O&q�ٷq*ua��ox�m��QzN�u��X��Jȉѥ�.�DW3Ckp�`�Ku���y@ov��������:B�Yk���|�6
t�Dp"fH��+
���5�h�[w#μ�j���G����ū6��v��3!�߻"��D�_�ڵ�`�j��Sh���Y���n��.փF�]��y���'�n-�:����Y�YB[���`H�B�5�D��@�m��ה8bl�Qs)�w���˳Yz��k�'Y[[kv¡G#]B��.�v4F)L�ʺ�<e�=5���ݭ;ͻ��Q����b��9�2�[��F{X����.��vukU��ǥEIZ=wRۗ�.Z�
�tk1��|ӡ�|�q���wmM�L*��o����:�&UPT{4!J��+iU�Pa�,���6vt,R���v3L�+ �t(�3K���u���ܦ�;uQ�����]q�= �P�E]nN�!�#oj�z�k}�����I����2�����3�!�ft�R��ƆE��2�lu��O3*1�k	U�9[u��ٰ�J�bE;�l�hI�[�'x�fS������.��P�qړjdy���5�裳�vfP�5E��pr����xE�(�i��|�Z�>��"��t�]��geJQt��H=�	�XN��ܷR��1e9����n�Ⱦ�x2k���ዩ��"V3�
�zD�����ܽ����r(8��tVYǹjt�C�z�ij��#���=��'P�_nDէ�[�D�i��{�
�r[Ɗ��	��(�kE��Ђ:���;z�kͩ��#�-l���<TZ�O;��\�լɝ�bRm���p�L.i��"1N]�:���\�FRI& �"'�7�R+u�됍Fd�mUܳo!����vr���`Vn
�?��l��(6�#Rr4�,b��� �rK���
�0aD6�i��2���T��E�
�sq��Æ��6�%rÊ���1a�7�Ԉ�%f��W��w]0S�W'���U��ʂ8�=���2
�clm� �2ږ��?]5�l �F��Վ�1:��̽������ob����ѥ�ΝV�t��K3n<��ds�i��F�@o\�nS�҉}tB�E6�T3��"h���M��4b�W�A�2�2R��L�ݑ;sN˲ke9�w�t�M�u��tY��{�ݪlj����)�F�k�Ҩ�w� �����O�^"�����Y]��2Q��݂�,��>��Cq��ΗʅL3��C��﫻��N����Hi��j��:��&T3�ԍ��K����=p�5eK*W}x!n�wfm�V�Vs�j�u׋1�2�udt�6�p�$��]G$E����@];dq�y�?f�]a}�{���[��ҾM�DL�L$��"8-���JV#���]����{�8vy�pm�H��L؍=�2�8'/(U�Hf�h�ƣ�M����]�g��L���eᗭt��jr.��x�ug&)�׌][�U��֒3k*A���t_Vڬ"�W�݃��v�Ҩ�4[��n�4t��$=/"�+)�[e]����ѝ���d=�uf��IR��r\^���3t�����F.�F�R���Q�)���ٔ� .%^6����X6t�ptB��R���)�x�nm&��"��l���ˢJ�E.M��H�;0�V�tF�ujt�5w���؅]��M���:�5��ɚL-�ZТc����S����Um^t��]m�|ga�V���Hǀgb2�rP�bĂ�c�q�Vv�oR��{1Ӭ��]��g�6����v��t�8�e����܎ұū�J<�nl�$�OJ�\�c�.���	�P�Ql�˻��Z��
���ceDp�ffu��-JSU�
)dbm
@���[�v�`��G.�6��Z������fn8>F~���m�~��xh}ו|��'���"���I���ޤ ،�*�S�zI$�I$�I$�ڮD�cE�����f�흈Vb�sLʜ�z�<�q�b�K7���e=�Ej<Mr�ĝ+g���	��W,ֽřw���Ր� �-���T��(w5rC6���˸��ʭ�SU@��p5Wt��48�B�7H碞�Ky����ip�+$���u['�nN�N�vM�t���۳F�gP�f�ԭ��3�R�˭����-lǙ���Cr��z�gf֓;5Ү���mqVTo�@�_R	��qC�H�ڕ�U�F�������5ЛR�n�����^eY<�B�?�]�.QE˴C͹2�d�oa��̶6�K�Wgr��na��hK�u�PR�><������n$F��7�9������@��s���q��,�� q�fP�J�vj�S-�ӺH��%W����	s�+��5|��W8(�_]��������,��8�v�:�M�j�4~��`�`�wQӹ��Yt��Y;&�Gl��Ph�̾�ڂ�_lv�;#P�G�����J��zŁ]�h��i}�nvn��L<*$�;F-�UueK�N<Y���At�rN.t���cOeQ+��F$��֜�pEP\�ߐ���A7���`V����u�إ[�r8N�.����1��h�f��Kz��}�yG$N5e��F沜�Ne��M�$ro��x}�-�2�Z�iJY[hq.�r���TP�I���ֵ�W-Y�bQm�c��f6T�\t�Le.�)���[r���堸�*#+
�t6��ZPU��.Y���9����J�H�5�˧=�K���Q�
��q11)��j��1)�C1�."���\p��fSK�`(�4�J��U����\
�6&5���Ī&�i�nd����h�t�T�30ȱ�s\q*�,�R���R�p��ծ�Դ��1���K�
��*Y�ႅ�B�ťkTUG�m�f�ZF�&0(I�y	�!-�>d4�,Q�YH�6}u��6�V	R�ku��t�\,)]emTh�\��n�Z-�����-�a�R�1�.S-1�nd�/��"eq[h[�0�պLu�`�%s0�i���w��j+��[e-Ԧ5��[J,EPX�+mUB�X���r�Qh�I_2��M6�D*���#[Qj����h����JcY����6�����������
�.ᭁnM*#���B���ܛI��'���um�����R� )k���_\s�I�����*���}��cU(쉵�	��Q������a��]���xMd�� �λ�8/�mYH�)���'�c����0�Xt��۵*��q�����0�v<�QE�v�M�HJ06)�<걛ԏ$���C��'ѼE����&u�~�V
o%'���b[��!�NA�U��n�(U��u�g�%W���Ş��3z�rgNf��n���3�0�r8V#�7Cg��T�m���}dӜؓ���&oVq��1|'ؕ�]1@&!���5W���~,�=\�oV�7_.�c��v3D$�&_Dw�S]x���r�̸���|�c؅m���x��}܉�o�[um]�*�����uT�.�ҍV�]T_PP�m��y��z�-n�������1�q�7y�夘:]�����A$療��^�v��â�m�5�������Ӎ�CR�;�.l0�\��+���d�.nf�Ea��;�<�u7��J�+�R�Z�.�Y�x�rCAn&cS7������_��l�k}+�xta�쥇����}�a{/�7��v��=��]9L��P�8�1(�[)���츆ww���4����K�yP�>2�����L�/�R���h��$��k�_���]p�]�߼�NbDn�gx��nu�ؼ�SV�0�\Fk��z�Q���k��H�0�O����`��>�9�/�w-�`�[y%�ta�:�k���.��8�y���SuN�f$�>�Tϗ�p��|6�̠�V���NU�������j-'9
�L�jE����;���؅��)i0�ʥ\�3Qٛ��B�us���dJp��r�!ʉ;�檄�ڋ殚�vr1e�k�U�E���0���Pi�J�VvQ�GG����~$SuʛoTɘ!�VU�-lM��a��m�5�����;D7���U�4/[7oy�fX�}kFj)`�Mͥr�_Z�-�f^M�4�,r�*��o�1 �R�Zx��\q�P�Ch�B�o#(���WQ.�Zk��+�y��B��8ud�:��2c弖X���r���c*��"T�L ���ɂ���\���dՊ�[�>*L��R�#���� x>�6��!���0=�,+x�F�T�|=\�߯fS�]6FJ�-����]a��{Cf�W˞��\���Ž>�H�@�p��|g��z��bW2�����]�nqowd��^���T��zZ/� �TTO-��֙�F�Ե�un����jm{����e���a�j�y���z�L�a�^�y�W��d{�$��B�b8h��託9*��L�euwk:�﷫QۉU�]���w��y6;bZy�mU�U�B���$!X3�+kH���(��*uK��"=����<c~��=�}�״o�8�G#��NS�8�cc)84���<0Ɍ^�\��*�ܙ�XhJ1��3lˋli˼�u�cjm��f���Udڼ��=�S�8�-Hn�o%�/xn���ң*SdH���7��R����y/�U{�(��O9<��K>�Փs��<�9+��cFd9���}c���ӝ[0U�7�lL��%iNlk��+���Wa����9������msm��H!�Ф}�!Ul>�.{n�3l�L��/q��3&X�ZM�XU^o"���d`i�Ħ��/�L���]<�s��}��F���$U�y�Fĺ	�o0�g�����n�;0�{�^>�u�2 `&��f�Ŋu΍7�B�6.��w{5�;-��}�5���W�vj"M��-�2�e�'���Ѳ����I-��/ݜh�ף~���0�P{���R�w��]KўT����'0��u�1�V���P��9��c۠�A�V*�m�]��딓�q���<�T�1^��>�j��z�_;צ9HT��y38����׮�&��.����2.㔪�HbV_�����x��je�9.uƢ�[f�$Te�k����I����R����/�]q����A��� �]�Jɬ��N s7q��=�}��1��
��p�jHo�|J�b�y�Ǩg��)K9�g���ͻ-9t�:E����wuq��POE�J���ħ��/����]z.�>�g��=m3/�j-��T2�Ң���!�Q�.�(��n�b�\��z�h{��dh|8w�T�����u�����\��G�˝�^S�q*���F�g�FU��&׺�g�X�s[�x0k�9�5�1O}43Y�l_jڰ[w"ۋ~>:"���������@����F��G���f�y �P^�˔1�`�\���^���dL�:��a֥���"Xf�f^wf����޷�#�qM��=��D�9�=|q%Sb1Q%y�g1��z�i|眤[�T^�CfN(J�V#�7C:&��e��/��(i�'>�t�ׁ�7r�{$��k�U��P*6_!0�{��6`���3cmˆc�
�aoMňn�4���9&GZs�� �@��G�Q�295+�p��t��� �Z���k�e�&��KVȜ���[MɚjmzR�����0�����c�k9|SY��E�T��������3�����@�]���O`���h�s���}ۜ��9^�`K��P~���s�m�=?k�53��������>J��z���B.�]eQ�FX3m�(.u��]�V��hGu������Knu\�av24T���b����*Ӌ�¦����[���Ǚ�z9MN[�2�ư~�[S���6�qؔVY�mU�q��0�oRH��k�Q}~��!�2�S;t{*�:
g���ϲ����jR:���d{��P�{�v)��{ms�)u��m$�t�Ӎ���N[ۋIΧle�Yv{�ط�vV���Y�BC�R��tv��Z�Wmb8{�Or���D��>���Tg)P���2��0��k����%�ړ@<�ӽ��w\��8���SV<����[�c��O(��pr�7Bd��M��rL�S7��7Ѷ~��e,.mr ;�a�j&wk���KY�2�N9 ����B���O�o�c�ݫ�Q��"RF�3ڒ�/���h����H][,o�fPO+p�AXM��L�^|�U[ț�)-|�\�HwT��QA��1�OYֻ4��{��������}�;Sa�b>�X
O$I�J�T'G� ��k���G�&��{)�l���][�6�?ul� Or�α����2�F�˲��E�8v�1�em<�	h;���'p���Hd>0�0\[D��q+�FRbK���t�����햓�j	�����TfZ}�#���"OW[�t��J,�ڡ��L@��J�ǻm�nq���˫�$�&m�-��!�ƅxZqE���;�������^u�w��;d��YDO��WYT^�-|4w�q��Z��Yw[���()μy~m��Ւ��BL\�;8ә���aNhC�$�A�&j��� �V��!�m<���ã3���*v��
I�0�{(ӏ��Ҷ�S��7�!�}ݤ�G5a��Ҝ))���Z�r��v�Y%�k)(�e.]6���i9t;2B�6u����oy�$U5�XT(�kE�]��N���ǘT\ms������ ��NE�q��Zg�8�g�G�^i���\ntʗ��9��F�u��Â�0Lw8 D�=!���=�+��Z��z"g'ݏ��ka�j2}����ˊ��؅�9���v.��,�ŗ������So��	V�)�~k��42!^��4_yk��z��瓕%����
�^�h�΋�HU�#�!W��X�϶�뙣+�|�j1h>W���L[�
�7�^�k�;	���turB�ׇMiz�V*������:X.Zq��	�q)�vʤ�>K%n�L?wlP��G�+D��)!�7��#4�w�j�^����A�]si��07��T�E[���_�=e"��)��pb^�k�2���m��_���~��1͇�u��}h���.�Ub����!���k�dhF��`{�\j&m�Bbj�d�M�)#��G��ʽθ�rS�G\5p�Q�t:�m�e�.���BW��0Q	8wo$a��]79����'�D6��6�����p���c�p��.�m������XKv�����9K���;�j��e��U�2�[q�6FrPF,e����{q^�}!�u��޸4�r
�Йbn�X��Z2�Lns��ʺ��ڟUq�{��!kv��,2:��n����
Jq��\�|�㕈��Q��rݜ@G�ݒ�Zdl���]q�-�@ʑ�վ�t�?=�"����':_��ʎ�ۥW��g�yW�W7$���c��^=&�]�s0���vJ�zg�:�I�
�玘��q�8���f�幯+_8ܳ/Z.�裔%,=�B��Ք������q;i�C���H���M�W4n�
��9��:�񥪅����M�@N�+�e�f�̪6m�Y��R�n햲yF�%�uގ;}W�6JW��}=)J�M�&��n9�)bT֫��C4n#�:�>u:2��@� sjH��z��'�	�5�#��r�#E�.��i�I�r�<��0��Iƽ����Wh�CFDli����}jm���m��K���:��Cs��0��H�QR�.�D�:��}`����	��0����_.��fA�b_;��i� ��b I�蜪.N���;}��Y�V��~����Pf3��H�Y��Bhȉ��O��[ōW0��"���4���N�5�މ�s�0.>�7�b����?]�׹<�vȺ�Fmp9m�x=ڍ�6�ݺ�YӵD:
� qjo]�4���2�eW�f�m/7�X/�J/�gX�^�)4'�"M�3e���Y�[)c�R��
�����'�X�پ�w�s�+��<*�%��뢆����:�~��)l܏�F��wʖЌ霗9�SM/�j5��u�����>��ӥ��JO�-�j��-����Y�	�u��*���[T;1$(�4k@��{]�:����/i�z����}��;	1�$*	Q�m��-��9R�2�j�jW]a����J��77��u�N��̢�(35"86;�X8�Me�J��ae�,ua���X�wn�tˬma���| �J�Љ.�i��i̳r�[���ྻ�V�����9	��I�ڂ0c���rf� �F��ǥn�v���p�[=Re�Nl�6ӆ��s+�]������=7�=Y��9f!k����y�AJ/+��9��2��9�FX9C� �"q�;"�WH�{�H�kN�[[�n�D�|��4���^������9i�lr��ݙ��J�n��-��ݪ�삮ޕ{o��`�QX)�k�_���JT��{ۊ�#S��O"4v'�r�VE�_t;����a��Y�+b-s)�[�$x�:wu4���r��TΖ�j5"咲��s��hncmQŗk�D��K��3b�����<�*�!��2R���0R9�����4oG!]��2�XƥІ��g
Yk!�Xr���(6I�l��3,62��4�R���R���i�!�.#L�O4tv�q@+�Pi	ÑIT;�p�8k:�� U�x��1�v�2�ռ�\��[g���^�f����?G�֒o�I$�I$�Ko�c'S��׏��l��	-&�,��a�yYXd�9�@�)ݽS2rc6�B"ͺkm�ら�P�h5������ED�^l�� u*u��ZT�%�ƈg�jz������W�i�@�P�)���l�{��9�e�jE.�`�`ӃSd˩���j����aۂ�h�"�u/.���^*��H��%�����ю5+x�ӫ�V�Y1��E��]�D#Xt���I�v���'�� bڳ�tev�lC[*]!z�^��Eq7���^ )Q�>wL�. +t0�bzH�8Cpڊ!��wA�D]�����H��u۫�A'C�`[/!�ȝ�a<�F1n��IB^�j�B�(���6��)U2�0����aE<�a������\:�1�{�� ��e�tE	��U�Fn@ְRʋ�B�/���.ƣ���w�ih��c��쀊�h!�@h����8���b�$�tôy*�9��G��Y잛�ha*TԠ۠��$ޭ�IF�E��j8NkV}���.���bdN�� �-�x�a�v�ԥ��y���D��(T�;1C�5]�KcĞ1 �RsxwJQȤN�r>�ͅ�$��}#��N8����~ϋ����g�c�)��V��MY��UT1�m�AIY�kZ��I�*Q��T�]S-)Z(�*����t%Ǝk1��L�YQq�YR�V[��2�Qs0���V���(At���=u�AqEm���QT��b�-��FEZ��D�Z�\..��e�r�gP�[R�J��+s+�����\���u��k��uB嶔mK�1պ�Y]�pR���jiZ,EИ麳YT޵�C-��T�1e��U�26�J���*ۉ���h\�+T�����7���7��	�YU�ara���V�����L������*��S�+s+nc���0SMwO2<�՚��31a�#�Ҷ�uJ�i�
��̸��L¢f��ݕ��Q�ppZe[�*�d��.ci�����2)��̶��+L.�� �-�33�i5�.T��-�4�H�eұT�w�\�GZ��Z��S,̣�̘��02T�(��\[�mˣ*�.9L�.y�ɦe��\W�Z*oz�GMM5SX�4c����&�]SZ�.�7m\��*[]T��Z�QkL�-˅�eʷ)G.�ɬ,VҰ��kF�]e���uL�&��ʛ�(�mƩ��2բU��zu�V\2�V���o& .�{����B��f?Lq*�,����k�E���Üq��j��-Eֽ��}���v��F4���RnS5���kt�-J=�0��n�s��yZ8�r����nG�UaB\��O�����o����`���ȣ�oo֧��\��U��5��6������[>�����9o+R�z�t���@�C�Ϝq���N���s���ᛄ|'���/��~W�^���^��O��!H�};�דD�n�'ow�w��$E���W��M}+�l�6{bA�WV�I�e\�a�VJ�|�w��󟁟x�J@B�ف<Ӿ��r��N�V��]z���w�K�*����J'�
,J���ZC�@�U����ٵ[�X�:Yi�w����t�����<����hz��Տ@6�j����J���دO0��'`�q���%��qpu1(�͓���宝�+霚H�x#�pד
�'p|�.b��X�Y��-@����/�V�U߷鯩����8>�);��#�&��9&ƞ�1��	n�E���5�%&�1���t8�j�'�Ux�7yԮJ��m�,�OR��vky�'2Nm��ƺ6�u+���ϩ�H=q)#���Y:_�A�{���o�S��{;EYl!V��~���qN vR����^^��חY��t;DH��U���z� ��8��Aڹ7S[e��D���V�5|r�߳mn�g<�Aݥ��^´f)@�NE���UG2��_���'8�f��s��Uy	57MP�&"n�S<��r���3�ݣ>QY�Z�%6���I9t�!�,��F������e���x������&��\��;񷷦Q�Om�1���5�bCT���*������;x�,��6�۳g_Z�m�]��R�gR��J��?��r�߭;9�͑%{3�]u�E�}�u{+f�u5���7����Nb��2ߏ�W*��w(�8{ �D�ӿ|{��bGj�U�J)�:A�X[������wծ<��nU�F�η�yc��t߫s�Mw�jK��'>��cۓ1ͅ��lc�����UḕΒjh�	S7�mŶ�N�!����^#���%tqo-������:W�73��:��$3��� >�\��[�3j�j/Kʪ/%.nk;���] ��P��LW%�R���T+�x�Q�a�y�ֈ��4�`VS��J��ܝIC�^�W�r6�+�j�9G�[1��1���GNs�|�޺淧&9F	W��Nte#�t�+�����µ�{�%O+YC�.5e��<�\�}����DI���m��R**�����Y�A���x����7u��E}�ќc㾬�fx�8�-��Y�+X�oP��wZ��J�ya-۫op��2��RΎ�<��x��BI��H�r�_iL^'�5(>V����p����]��<:��x�ؒ�.���3LeIhm�q7�rT:��8Љ�Em�s�[1�w��J8����N�(O�'o�*o����3g�T�WJ��*�nv�}ݸ JC^� ��ޡo�b���*ʬ��x��h�K��R7N#�b��pvV��<�u,Òm(�q7zV�;gxV7���X9��0��������)�9�ծ��ŏK�3�脩I�)#��<�r�;��2��Tۼ�mC�u,,@Ϊ.�B7�9ʓ��v�n>Sx�kl��Y�k�ӝR�=6F}9�J��>ڷ#�f�:������/��U��;:��s��O�:� �M�K����_��Z���+t��ے�|�z+�Zd��H^�aH�wv��y�'ҭ���a����:�E4�)1;� z��Zw¹�oLV_H��`w
d!��z�|XT�ɭR|��ݙ��O��m�20���I׬��/���o&����~��8�br}CL�����a:�Ԙ�s\�@�4g0ud�a��}I9�2��&�d���O�} DyǼc���zE��O�v��]W��D��N�L���uS�������2e���$:�Xk9��u�G�,4���ٙ	�xɯl>d���&\�����ޘ����SuPǼ>Tx|��8�6�d��i"����d:��9��O-	��z��&Zv�Y+'�y��$�&��Y?2O�}���?��������۫�O\`t�a�	��h|���<CL�`o�'��I�]�I�L�܇wd�f�̇R~k!�Y��* ߕx	�1�����s~�vt���	U���+�lLt�dJ��o^n�1nP���Z	� �6��r��f~��-����H���y�H���z��ݏwk+fuL�	/4�"�����\�:�C�ϻ���uwL�Jki�/R�$ިܑ���I֩��E���}U����'�r�q����I�y����~��i��,���ԝI�x��S>�!��&��l:���';���{���]W�W.�����
�����" ���M��M3��j��2k}�� ky�qY&���'d�'�>`v������j�ϰ��|s������ c��<>��q���!�߰��z�a���=d����BT=a�'Y�<Ր�2h.��d��o�N"�d�';l7��o�~�n����j��w�� �̏�׼xyg�ROP�����!���I<f0�7�x�z���4��
��1���X�{��"#��@����'	�gW?�*��>�I���:���4yI>a��o�!���5��x�	Ğِ?3�C��`���g̓���OY�CYg�4��"<?�=%�i�uD��g�1i�xlz�O��O�57��N[$��6�!��08�oS���o���>Bq�@�6Ɍ���0��+w�8�)����ֻ�k}�￸��k8,��E��i��Xve�Y57��$�����	�x��N�9�0�3�n}�V7�q����q��Ty���F<��33�}5��I��g�`��:��Y?"�yl9l���2jo��	�fs	��'5d���!�I��?~�+	��U�/��������;���� �{� �����:�d����8��E���fS�����1<�������� �g���_7Xt|�F��fOw�����ɶ�w�p6�2M��5�~f�5���&"���d�*��u&�X�$�=a�̞j��䛋�{�������g�/��\�.3q�19,�]�7�nG�V�z��׼�)z���2p3�ʌ<���Ȓ�0J+�⌨�Z�Tه{x��j\���fd�Hw(Y��cnL��7}�M����&6�,��TI!֙,L�8܄��ܼ�J����{ ��xd{c޸��d��g�>C�'�{��'���,:��LE���� T8��'|�&G��uO���@�Tc��i�_۷5��g�s^y�;&�LgNP�����&�q��h��$�
�L���Y'�d:��,ü�-���a�T:�����e|��]�if��-
���\��$��d>I�,>d���0'̇SL:�Hq���
���H�u?~�Qd��9N�<�CGy�P<I�A7����M{�מ��H�~����ɹ��M?��M��<d��Ì=�u&��I����O��?$�'�>�{��@����z�z
���k��ϓ����:d����@񇎘n}�@�����5y>��8��	��}�N2OP�,�C�OǶLd�h�ɴ���}73����;'�ޤ�ؼ?xz`I��rn�i�{����2NSim4�~�+	���BT�,���Al��:ɩ�ru�z��d�)'����~�6,��t��=��7;�:<��ğZw�	����2݄�����:���ß����Ɉo��=d�=�E	XC�Ri3�P���L�:�y�kW��v�}����= �O�{����ԟ�;l��~a���u?v�S�'�;�I��''~���~q'��x�d�Lg���f�|��>�o3��C�d�>gMR�i�}��?$�Ԝd���l�d�4{��Xz��C�koR��~g�O��I:�Cݾ���˯��Ï}�}��i�}��<d�N��x���:�4e!�Ơ����r�'�ܓ��`x�a��~;ܐ8�g�� ��!�93}1V-D��dfՊ��.��d��MŎ��J��!rn7��κ��sʺ�X1D@+|NvI�̫�����?ʖK�eaes��E��c�k�K�Z)u5���st�mL̼�6 ���Ю�# �	|%dՕ�����1�]�z�u��3G��Q���2�+s�,�$���E��(E�I�''�XN0v��̟����{IԞ=`o�0>d�>��ۿr�g�~��~s�����ē�׬��N['Xx����a'�+Oy��qr�'�P�>I�'m��h q&���I�xQ��/���/7��j/3�: ǌ3��l�w���a07�`m���Y>a�Lg��su%a�{��$�4r�'�-���[&�@���q
�3?`��zK;�Բ�>��W��g��g'��o���I��ܺ�~CH��U��`N!Y;�(��I��O��<�9�魗/��4�1��1�t{�=�G�����	���Y��h��|�X�$�S��g&���~E!���O1������r�w�_5y��������Ώ�I�N�X�	��d�+�M�q���[�$>d6���|��w܀��M��I�=���M߲I���<v�ʬӂO}�ܶ޿	���Z��~@�a��ua���~a>�dRW����IY�P�$=퓬�gl<�ćS�XJ��.���������cw����>���{ ZU�@�-��su���zԓ������$�hM3l���&3��Ϙ{� T{�@G�N�Lm�����r�g>�ٯ:I�M�Ӟa%I��!�XM����-������2cw�HT8�+	�O���8��Bmk�@��8������k�����c�?3�'S�4��OP6���G��8�����4͟s!�O��o����=t����+%I���d+�6��N�����������F��~#^�~���r����䧴��-�ҟ<��F�u4�:vם�IB��oT�G��|
-�(�Eb������=Ed�zu�"�Cl�X�h��ٱ�*��Ů�]jr���WW<��Hļ�fI:���jHo����UT��:�s��{ Tx�s�>�{� ^]�O���$�,���z�������������u���Cg9�������t{�؋��P�:���b����	P;7`m�L�Ր�4oܜa?$��N��k�p8��Cg��8��M��� u5�r~z�~a�~��OϼV.Л����\���Ͻ�8�Ǉ����d�w?Qd�<HV���!�{����,�Ԛ7ܓ������$�����O�:��k�C�7��k��|�y�,0�I�WK��m	|q�!��	�
饓S�����N3i2��4��,6e!�'Y57�!��I�d����O�yL�#L��9��;w�/����lBq����d>d8���zͲ��a?0�>��P�$��`~I�'�8��H~I�M�$�<�y���_:׺���<��I�Y'Y:�i���<���<z�NX	g���~B|����+8����B~aP��,����,�� Dy@��޴���;�����IӼĚ`w��O��w!�䓉���i���x�|�+	�o�3��3HNs$�d�8�>� (g�ȫ$���خJY���о[rh�u��#ި:[��?ZE�Y=��!8���d6�a8�j�m��4g'�l�_h��}�N0=f�7�d�!�LE�����a-2����<`z���@� DI夝���O�ɲ�q�ԛw3;�N06~�z�q���6��0���:� ���PLM�����߭����Ǽ��}���Ԙ�6k�	�+&��Y'Xq�O�a=��?2jj���6��>d=7Ag���5��&�����^�>��p۠��#.��v�TxM�ف)kk��̙B�ޣtz'��|�	�+�w@�|;p5�!��ζ5*���%�sY��P|�V�r��s`;��Uܘ�W��R�鞊Ӈ6.�ÉDbQũ.�=��{�Dz �/���������L�l*��z�0��ϳ��~E�ĝI������:�X_��|��������'�}�"=>��<���bΜC�<�>~��Z�o�������/��N��1����8�
~�Ê�8���d����xɖ��̐�%a�9��u��,1=a9�	�x�߿{�k�~�����Vy�Hs�i���gx{`)�"�$Ru<?s!�`��Y<�&���b��ho��
�;���'Y9��a��՝�]٭D��?�z��§��gY5��'�5��M��&���!�N06y�I�'RuI��OO��wvI�o�ì�d7�d��<LC~}��������~s�~���`,
Þ�5	���x�P�j�'��'Y'�6k$�:����>E���u'Y��O:�~�Ͻ�#=�¾"Rz�r��U��vtNga�x���=`z�n��{���Bm���'���l�<5Bz�`jo;�� n��d�򓬜E��i? |�ّ�n���?�q�=Q���Ǉ�<{���Cÿ���z�a��<d���"�,�Xz��u&���i�|��:���y���}lno�9��}Yw�>��>@���N�Y�f��O^������:�����y�'��Փl'�������c'Y>2���ԝ�c�՗���j�ȏ�G���g��g��8������N'����������',Y�C�s>d��_k�d�U����>�_W�71���v�r�!Zw��T�&�aܤ=I�MM�$�@���}l��~�:�ǉ����6�<;�$�ܿ�����3 �=d�|��0��&z�o��u%�_vY��*<-9�Wi�	��FL�#(�εud;dl�g}2X��H��e�d��"�΄�Zg�pz`ͭ�Ք�#�O�T���Lf��e��t��j>ُ���o8��-����eÛMQ�%�rƎ_/����߿}���C� P��(�(
E�E���Qb��

~����8w�Ί0`iP�<I�O�a��|��&��Z�|ɼ�I�	�o��0�:��0�g����B�zԸ�xW܋�3������;�*��2c?*I��CϰQd�CS�(E��`x��dP?$����kP�07��m�I��Փ�O�ӌ�l�[�/�����0w��<&<<�k�@����d�Cl��yBu���h��8�9E����e8��O��as :¦���o�&ޡ8�=��~5p���k���|�睐��`w7�����3��Gy�Hz� y�d:�l��7��Rd�nv�$�L�Om$̼@��*=�3�8�����H�g�~������!���:��d:�2i1�$�
�ߵ��8�o��i��Hn�C�=d�Y��:�����$���Y=a8�۴��T��w��̚��lxL
�{��>�4��L��y7`,>d�k����+4}��E�i��myd6�m��y�:�P�|�������7�}��_o�9l'̝��m�$�?2z���$��k�	�!�Si���=�1�����d�~���8��`u�ɟxR9�t#�9��y��On��@�D�r�	��hN���r+�G���d����ku~���>I�)&��B���сa������箛9(%x1 ���]��'mXc��u��Z����kDX�B-�w����QY�j ��D]������	��Y�o���Z<u�������f���Q���,/3,�
�R�C^ uW,n][]�	�N����mubҧ<�29�ۖ�<��s��$;_P{�#7Ւ���{ ��9.jV�t7�z�l�����[B�����i��Fzm�N�y�m#E�����[�Cq2���v',��y��	XH�h��p�����ȳ�`�����u���U�f1��:�k;�X��;'Wj�Ok��m����4���Ttu�(ᣙ=X��*�l�I'�ī7�������B71�u�]	��I�ŖS�c���e�h��Ebʻ���s���lo�C��񓡫w��N���X��Ɖ�a�i�0���n����\�]��E�S;3�u.��32K�5�p�BMt�
0�0V��ub��n<C�,|@gF�����"����LW�����u�Bp׻��q���%�2ԙ;�]v4�Ϝy��VFS4�p�7K��J�m1E��4U��:wɕ�%�Ғ�������r��P���)y-��'2���IJ����i����ok��oh^�ocг�F�B��+�t�����豆��2tv�k;�	��eV��s�Dg/��]�P�q��߻�%'�I$�I$�I$���KW�>�-�лƜLߵ�%��d�umK4/d��b�1S=�N�$켹�͚�7.�b�ʊH SҲV!u�M�H���\�x�\oQ�:;-�4�[��t:pGҬN�yf]��i�\AùQ��œˬ���{�1mր�����h}�w�՚j񻊬Um%��EYT�9Yt�!tthan,ѹxiܳ;�Fj�f�Z\K���X��8Z��P+TQ�S
wrDY�j�F�
��;T�B6yq7��#x�	�Go���f�ԏ���Hwk1�\9�y��G�0=Wד�k"�C!��C-�v�uһh�4���+�q�BFĄ/�K�Sbx�j%��2ִ�R'�9e\���C>'��^�.�N�ȩa��`r�^�]��iWbª�C28��2��F˴�p���Mu��#ek	;i+�>�nI5�9�/㸣���l��F5�]�8��0*�f7C��33��a,Z땥v*��h�R�J��NQ%�3t���cp�Zn�@WNʄh�I�2�"����S�X7+r�gS�:�!
k8�0��z�4��F\�{�6��2	MR��	$�ZLn4�P�$��k.G$����H�q��ݬ����2�`��f	�f\K�-KZ�)����%F�YW5s+������]3
�V�6��r��34ZⱣ��ZJ��S.*�\1;|�M�r�j�L�p�kW�3tZ��+g���E��1[�&%mŹ��7�E2���(�d̲��:���j�.%.F�\��Z�K2���&��q��0mpȹs1rw�"9��nU�S��k)��)��31��V*��t�-�i���]����1r�+�r��q��֛h �R����ec2�b�-VMR娢���[E�U��n7*�-Q��i*/��h+�T���kR�Qb*e\��e�3*.R��K-e�b�£�}�1�eӒ1TQ�J�X�mMYX�V�F�m�k+|�Z�h�G�+sD`�J�l�B��mcq�ݸ�b�1TjT!��	!l?�.���j��J���-��¶�N7ZnK��pr��ոҍ�����uff��Wz�1"�U� ʋ�9��]8���8ٵ+jA-j�J�37#7��t�n�ĺSV��T���v���|R��2Lm�弖 ��N�$��Tp�3����ԏZכ�`"��O�"��,�u`�Gt��;GfgW?¯����^<m���d�n%���ה��Xyq<z�L�7X��)��f�X�)�Z�Z��g��Gsr�_��dmЙ�BqЂ���j���m�#�=Y.�&�;獍�I����lW�H��X��SN��Ў�@��bEUMoN��/��Z������"u�6F|UL���3��y2>�u�\��L6��3��^ǔ_���e�m�޿濫�,<1R��<��罳nQG�n繞�G;T�@�%ߛs.x+��y��jz�L16x�d�:Z������H��E�I䋠g֔t75q<�/u�5�������U����_W�*��Dk_O����ʱG�zZ�;
���;Z�lܓ7Fw5�C�3��Y��ͭ٬f��ӥ���ֳ�K�����'&%q'��s1*��C�8�R�	��h(Gk ��g4��2�T��v�֚S��4rJH�������G����Ύ�5���ɉJ#��Vsx��w���N�㹫ā k�ŝ51ֆ���.a�%d3��"�t]#��&l�N��^���Y�Vԡ\�bRwA��$5p���}&�^uB.�ÇuU;�+�x�)ַ�`�lSݮ��X�t������5V�����g{�_\�Q���Ux�#-8#�׻Q+倖��Y+��Og=T�V��|�1%2_���r������]cw�B��uV�o/)=�L��]���JK������%���/�
�V |��;���9Y�i�Me��ұ9!����d��@�9<�װ�_����(z��[��'��jrK��]���S���ʵ��7�&����g�^���,g��p�ƅ*ͅ�[΍eu|�Ǟ����0p���s��b�IFU��4m&X��D�@��ո�Y�3���N��;HKZ��9�Mv�j�R]��ȐU��yc&u*7��7S<��=uE�L��x���c5�ח��#&tt��B��;�g���=������7u�����>�/(�xo��RM��ސ�s�>�s����C����򣥩��KV�4�����{�4�773X͋Mvi����'&A�������\+��J�U����=�/WW<JN�,�T�Sb�lL�l�P}�_o���C��oS�՘�ˆ:�v!���4�B�p8��:�1�nU17i�֧j�X��Hx)7�W��`���</��X�E�LY�7�6ͿnDҐ�7~�(PA���$�Qs�8�,�:v���w.[���j��W�h��e��u�9m����$���(�(뼾g��h*�"�|Ϫ�8}�Rӣ��������c3��ɉN>�+�j���¬VU�B�6���>��h�^)�c�S���2	��U��Px��<`N):�;,f��U���w�%� ���,a�Rw4JȎ�s��QD۷Ju�Ļz�(,��N7�/qa�ʚn�Iùk�3�Qu���軩��hMQ���CN�[�s������I���'��:�Ry�ͬ۝k����ՔP��W�"`sxVJ�t��n�&�{Ҍ���ym�>x�HF󄛜�b�K�ͱȥ�F�(���j�U�iD�o�޺yYdEL���*F��v�>��v��,�J�'V���E�M?;�jQO-�����P�V':�;��>�Ȍ��쌉���ݫ(�A:6�w��6�Z�����l{�[���z�:���.��&�Rڝ��~T���΂!�����)��|��Fn�c��qE�v�:���Sa�������1nU�.�Y�������ӕ��"�E�݇8(4�A�‖).���l�'�9S�BiɅ=U�1�4���u�D'`��#�����*ɳ1	ڡ�\�+\������,�zv���℺(\���^&|���"�PT�m�-
���g�|��J��`�)�X#��Uͻ����ύY=�V�����'�[�2��V�K)$f+�\�v6�$? ��wV�֝�Ԕ~��gl�P��}J�����AΦ<$j���~���(��y�����1��b�uY�Du�v7)�K�S�V]�!�u���y%t|�"CW:�.����o^����wo#�w�*�=����)=ǱS=�O}C���\W��Ը �� B�W��G�	ﲔ�b�Q%$����2�lF���j���5�/nz��*�/H�'�Ӄ��i�x�۽����&�)ٱ8�>����c���-�ڢ�׋|q(�eh\�ʭ�H�����k�{�ܽ4'��]��}t�*g�zq�Ckƹ�[S�p��̞\h�T�>m��;�ؚ4g23΢ۥV!B�u�{c�@�0ڒM���j//e5�DS�>��V�S%*��>9�c�8��$K��z��d�Uؕ�B+����ON�����̔��̊��^����ڌQ�+E�����t�m���-�w�{ڦ�Ֆ!Ŵ-78Ʀt'�S�v��޽�JS�����6v^�D����MV����_W��}B.z������Y;}h�vD�Fy�e{���-�.Zʹ���ۨ�Cd��W��D�ק�wiVR*�P�(�f7�{/���x{�.Q@���p��m��镱s"�Ի�#�=�۱r촲�Eև�W����0�����T�Fh�5Y&��o�%L^
ukpع�j�f|�9�U��b�}MҟB9�j�]�ܺ�Z؉�4Đ��Qs8�J�g�+j(�tD����}N�)�&8�/�t�����ܬU/�Q����-E��\<��m�y�������n��2�r�����-�!�E�X�"g�Yo�0u��o⡶���׮��v�Ws�v�B�y��c��D��K��޹릻p��r��]�n�P�l�+}��.�a�əo3 ���]�������w�8�4�p��|L3�\���#Z���m����0>7\��5��_�u�*I�I�-�Y8a᭻a���孾	;a�o��VT�`���gf	w�B�޽���,�Iw�� ������&���O������>Wԅmzr����Qhi���k$sһn�m�f������+�Y�Cn�9\����ی"�x��Ȫ��~Ǳi��yW#Uw�j-�U��z��[vdc�i��{�/��k<���D�����dd��/v�ȁ���ôy�z���qDN�=\eS���r�"A�WVFS+�j{,�</�/sQ��&�����4j�,mP�yg�l5g$JW�.D6l���7yi�|��+���T�Ns�1�{���F��ηk�2V����q����X.HV�;t�H>���b��9U�H��]X#Wa*�z�e��`���k��
�$��8BP�G��vRΚ+e�h�t��fP~յc)bz���0������W��wxs��ш՜�1cU�;}:�S��ýAQ���x{vU���* c!���Q��gVkB[7+�K5���f��wuޭ�r�8&�@ӡ�O��ȅ֚o��L�Uҏ�d{Eu^l��EI6�F�#8�]s`d_:6h۾%J��󶶃9u>�ȗ%\�F��ҁ]��!���_}UD��yľ�G�+#���o	B��i�����&b�!dNb�s���}ք?k��4b��C��e�g-�x)�f�����O������ֱ��N��/��(v0�"��cg���楳U�����y��=�����F�Im�G^���*�*�n��3�n�M��,���e����պ���7�n�5���n�e)��uV%=��2K���T� K����#Ew=�w�S}��B=��]�v	x��7�m�[��LN*,mQ�bQV�#��m���!%V�i��A��w���<d�O�.�	�b7���8�v��V���НT���CJ�ݴ[�cU8()�bcu��z��G4��W�Jd�HT^���Y��&!��sc�ԭ���)}���XǗ�N.��#x�)iʎ?p[�tV�[j�>��I�-�.���fsco:G���53\m�8)u��4@M'����8�|J.���Kʆ��V�l2����]�����1f$ڌ�ԕ/�t�s4J�$�+�!�>�����1§��n{_��5�%��ƍԷK�!�v�̃�J+͇Hl��&��d�mQ�b�!H�yK"��#�:26��PLfJ�od����1���gP��T�j��2�*�W�XA2#Z)��.~o�D�m�U��s�{!�Ժ<���+n���mDjw]H��G+�Jna�WD��7���#���#�b��ZoN��^�#qKN�QwE�D������E�gGF���"97�,����ΊZm��f��=!�ˮj/����IV4:
���7��N����Ή7���z��Rqc�[�:�t�O���Fs��Y|����hEY�`VU�E1W���A	μym��t����]���Ȩ��E�N�U��xv�%�2�s7 ��s�lp�M�W��*���L�ID��#[�>��r����Y��Ը��4�O��}���5"1ޘ��y���Z���t���:�}f���D*�j�o��0����K������ۅ�&��VZ���$�ά�mP<6�'���VrLC�q�Ng<�Lv���E����zdm���`����;�#i�2m�$��N)��DR<�ǹQhd���!bT��h�[044����GGl����T"�*L��.��ϥO���$r�'\*���M���?k�>�S���vă��K���.1�f˚���$����4��/��O���_N��B��:�'1����{iI������m�*�h�Y}�j���?�8�٭�Cq<'v�:�)
G�B��r�Vu!O�C5���ZvUD�f�(�I<�4�W�U|�Y�6�9��z��t5�y'4��<#^���N�Qs8�J�g�h�����/�8~�6lW����{յ�9N��'19�&�¯V���a$6����˳��#Tm�J�v*s�Z�3�y��%���g$��9���mCq��u�
�R7g:	r{[WK�i\��&�0��;]����K����qCqR�������}tۈG�$`�)J��:LB|)gݧ&��K:��P�a�Y�ͻ���m��`�+���7���hN�[�>ZEl��|^r�lM2�Ыb�]�1���r���+�s6Nˣ!���,3#S�j�)��{�n�lm5}�%�H���;���5��7�k!t�vtK�jyN� �lbn��\imѺU�����f�T�#JKOw�0����Ug���M�����.�`�GT��eEQ��s'X�>�䵭�2-e^�6o@ʽ�(Fdve�n�Ğ)/r�.wG	�m��5b�Z�	��m�)488{�Ƈ@-�f��4��]q�fE�ƚ�Y�Z�3yZ1��jٺ5F䓥;]Hi����9�����A��ty�C��qb��fh'h���])7-�]�J#����V�+�O^��x�_	tI��_��%J���3�SD�h�w52��]�	�-flC.�5@��R��|ѻ�7�m[5V�;Q]�ɕ���l\�6�y�{]Ǩ�rK}�%F6���"x�t'��ܳ���˔b푆$L��<'�n��m$�RI$�I$D�ޗ�+w,:��:�������w_8��w2;����Y��{�5gL��6�I��-��,�h�E�A!�z@��+9��\�LRe��qk����w�ۆRwh]�ǈQ��9��Z���`u���(�f�@����n,]�A>)`�Le#���0I�l�$�\ �h���)L�������e
��eY�Ԍ,Tޭ�CDz��V����c6z�������:�-.��ށ�+Kd�M��x�Vd%� Wω���q�55��vmd���]�;�sl�K�D�R�̸h8F.�I�ƫ�1\詺ٻ���G�k-#vJRh<ۼF7`�y��L<�Xr[��(�u����ӈhCi�Y7�:/����t�ܔ�D�]#��M�=�8�?5% jr�)��[-eM� sn���Xtl�] �)��� ={��x�Zek�
����u�V��Q��1g_�J���i@t�v7y�����
7$Kb�O��m
ɪ���>֢�f�5w%7%�ݹ��*'2]!���E
��T��&>�8�F�.1�e�����rH[29$�F�z�V
��VYU�-���
%���ml�\/��b���)Bʊ"%�NS2��jPU� ��QRҋ*�V�-�A��Q����� �B��֣ƕiq���J�KB�kU�,��)�T1*�ѵҕ�[j��V2���Eˬ�P�Q���-�Z��,��F%��6ck-m���Ց�Z�Do/�"j"�TD��mQ�����
�6�ؤ���-�kU�[�00����f�r�-�QT�����9�-��f��+�ŮZ�(�-��.[.U0�k12ڮkEJ��0ij�k+L)R�ܲ��F��r���)/��e����#kG2�
�Q�Tˉ�T-���k��*���aE�kQ��,i[eK��-�Ɵ�nyp������ar�1�#�����Ŝ*�@m2��B�v$Tjdi�Qn�T�9�y^��++8a��y,~��<1nv�Ac�Q���l���pr11;��+2�!�bͽ�J��s�]riE&0�o2]!����>���'�Z��홭˳�n>S�22$V�W�ކ����Ͷ�y�ŗ=�Ɏ�u�ٝZ����`w.�m�DH=Jnl���^6sdu�pf�s|��t_��s~��ۊ�|P���n�dR@����B��q��;�*̽�a-W��m���'$3��6�ӕ��u��Vy��He�nug^�oL�p���z���AW#Ӗ��x"����9�����I�8��S"WE��o<��'�Cξ�%�Y���2j���a�*�H�>��D�G��Ӎ���_VX?S����b�ӷ~:�s���k�X�/}��=���ʎ����,�93�ֆ�;�کm��;�����5���>�cs]��~�j8,���O��m�w�^�}�,l��g.q�F�u,8���k�
s���W�C�^E㪙��pj��U���}��;�
2j��|�Fs%��u����,�d6�H��u)�S�υ�Və��u��RX�R��RG�����j��o]B(��˷����_��~#�D�z�s$CT�G�|I
hen��)�*(��n���g�������ͦ2�×�9d�K��_U5�[M���N�\�%P�q[b.FDL5������Y���	ϘU��%�x� �dpj.b�n&�c��a���k^-NW�s�V��u�+�M��(RSw��Me)���$�6�ǾN�����I]{-ڰ����Uo5E��/�Ri���Q�pһ�b3�����e�F�t��V:1�Y슙\��~���y�Ħ��y�n�4u莼������]�0�j}��ky�WUQ��V�5��.u�������4����(Pyu�}�d��J�ٙc�E��n+׋�����x��x�HNZ�h���T���[HV'����5ebR��EL�ٵ����6i���i��L�AW]�^��ݑ�\C�p ]vn���&)`#�%���85��i�Q�K�������O;�uƄ��u�N�<4�2�}ӓw�eZ;⫦$mWc������܇"��^T��D��WGc�q"��8�N�ʼ圆�$��y={;
�#m���ʳ����m<#�q��P�K�f�=��Ollm��J�w�PO5cꔆ�{q��d�CUQ�Ο#���I]X+��q@c�6&VtM==l��D�Nw21�hˍ�#��(�[��iԉJ
��A�Wrw���Иbl�>�Ɏ���$Rȯ����H�5��P�H7��L�=��iC��1T�)pj��d�����"'���2�%t���C�8�(S<(���
��2ʱ�_DLg3z�+�5��ɑ6l[�s�)E�W��Y���yt�=�f�:���?x�괔����*.�o(�[Xsj��̺Ղ��.��9�GSWM������E��>�z�|���7��o�����պ�k�P�����݆&��4��,�ʖ�pFj��C����B	�8%L�q�ﾯ���P����S�_���;I�cQwI��Wmg���[*�/_$�r��˕���ö�~y��VS{��p���yu`>���GY���a�|٭�{a�b�/�oCu+G��0�{��9<���kGy���Pֱ�^B1��W61K0��{EX�{i�Dv�#�Rc�d�(EA��'�xmx����v�M��Ǻ��%�ZԷO�wv�N]�B��q�(mq�V�8 �y�l2�,��ݫ)�;�J�j��_�[r
�����6ϫ��q�[����#؅��O���V��R�r������x����t���nGN��r����
�d��U�p]�\>S���x�9W������9�s�܈�dÜ�O�/<Z���0rSn9���EZ���5�/�(�ک�}��+ʛ�4�w=�N����5���wUr��w�:
*��	�3l������O^��o��������\x4x�1۪2rN��%��Iw�� w��}��;��!�:ĭ&e������k<W�ӄ�6�����5�+5�s$R�W�!P���΢/��MU��U3.|��,�'�>���d?�w��/�4X���������jv�%γ�.y����Jyk.a��Y��+�HN��*L�ȥ]a]7{(pv514��j�}�#��Z�SY�����n9�oI��I���1�j:٢5=�¡��'I���M���̮�c�;Du��mY���h���[�l�A��d��<�J<���q����/:R U�xoc���|�,Ԕ�n�|k�wٽ���zc���*�%���!�h˼s>{��\���s0:΄x���u[���,N]f6�r�u-�21��^���u��*�ͽ�N���EMb����=��οdw�4��LԾ�K���}�4�3R��)m"s��w_`�o+�uݒm��ܸ_U��B�]�::ٴě����7u��Zb�k(v�J�VN�3/�Xzl*⭽r��� �}�8��T�%v�I�ﾯ��i���.�V\�sb�\��G�t�;�w<�vJ!nC)�lz�f��aR4%Ɣ!;z��}�}<����]���oN0m�/"]6��w����{#�Z���xϧ�������=ns6����Zu��2K����[>z�Ն|)��y�z�0j����w��<�}J{��Jw?f�{�
�r���P�[D�LQ:=+ʸ_3��u+�G�7I~oǻhz_;�����svyXU���O��%R4+��f���ʓ��6[�-��hep��#+��6F̟q��2pE�Of��S�����*��:���{wFo��E*D
c�<�ʴ���Cw�R���X��U1u:�H�v�m�4���O����(�=�e�Yʊ����x�5x%l�=��C�����[̴������@�Ou�^�0�y��qQRzlˀa���}D��E�DI�'���Ԭq�ہ"&���OK:Q��e��!����\�̬Є�p�������\��C�`��c�(�y�?�U_W�,��/�Lׇ���X�<0����0
���u��x,�#/	�ʓ�E�9�3�S�{�����dH�U�Uɋ;Ӟs��qa���,c8���qV�X�r5u�����"T�(1yC���Tߑ��s�^��8�V:�P�
���;Q�9����N�=藷=f0J�[�mSFK���!tNGCU���-��R���w`Rw^��s����|~P�GY𔲺�]T�U��d��#ձ�X\G7FL�,��=�M	� Ǿ]�����*U�V��#�"yh����+��ukKl��ʎRw�{V[:V��P��F��]A����:�K�GD�XF�g�ᓏu%��J_�P�o�`Z|Cn�)>��:�8��^�Ȉ�&v:WYׇ3��Kc�ژ��Y�9Ɲ�l"��Q�Y^��Fg�\��7q\�K����Y��1�Ͼ�,[::5��p�\����O�U�|�R���8�id�Lg�Q�wJ��7�{�i[*d�yyPm<g�D��p�0�1X�=�n���B��T�1Lq��i�\U�pX��[��ݗ=�NWF;/�H�`ouk�wt�86Ky�Ӫyч��)
���y'WrK�����/n��Y��L}�rf�V�9�]q>��z�e�c����V:|=h�i3����t=�/1Vm{�c[�s��^8T(����.��kn�vl��o{���Q)�P���,�49�pK������Bb��nyR��R��*||l��с�Q\��D)/ʄF��3Ҽ��
�/���d��`��Z�lu�N{����)���R�$8��2���;�HWx�w�pV-�l �^0|��+���M��#y��\l�G�f�%;��"�W�
���m6�Ƹ�/j$�8�虋�˾^��#�N�Zb��S�d(�8^r��ר;��ꘫ���<H����h��{�4Z�����9g\�3�}Cl�̤EÂ�����`u<��t�s9����g�^nA�w����o�K�}gG���~�������\-e��K6o��K� ��!�Ժ4���&*P�d�x�Ӑ��ȥ�
��>��E���S�U�c�uۜ���(����{+!�<��sM�To��	���^�7�L�e�˛\��5#��(���Ϋ�ҧ%���0� ���35���GS2��eY���riTg��k(�r�%sU�h�qt�Ԑ�<zZ��	i=&\�����W�U_�G<o01u�0��%6�Y�}�O��lۏ�ۨs�hN��*z�ީ�W�.)gj�|X����)��藱A�n�.��蠸�O
=�au������g�B����y�mr���Z89��`����ҍp�5cB��E�Ƶ���V�ե����ש�U���X]�����S7*�$G����"Pa�գ�ܠ�]��0�؝�� ���cm��]�D��﮼f.�,b屬{<6���C����)9��;�zo����3�3ѽ�4��"ӭ�DPt*�d�Gƶ]n��A]:���d��B��6
�W��t�(�Jg_�'94���F�1q�꬙r���ըɼ���M(�|�F�ӝ1R+�Й���Bg"ܹ��<��]a�&t���������톍��u�1^;eE��/���`�);ٛT��R�Il(ʻ7�R�oy�"���ﲍ��IT��S��;
p��pŀ�:I�B3�k6eou�FIWY�[�fЕ��k��TC��7�����V��y�D���GΉ�9��"�����ި��n�m9�<��v
m�0�_VF&�g�U��o�ѝ|�&���Y�G*�����	S:��n����3��m����j$w]f���/h��Y��pR9Uļ���&Z�s���>��O-�{�j������BŎ�WϽ�'��B����m�<+2=t+޻������8Ԙ{q[��SHeP�;���~{Wʮ;@Urm,��d��8����G���o�s�@�X�L@P�O�����\�^tl8[$<dj�WIXz��x�ъy����yd[l:�X89�T�|��qn�cG����ܷ`4���)�ź�s5zc�2���*V��KG	�e/.%ѵLhѨ��>[MݓG |���C�؅��Y�V��\�T��g��᳛����xh�F�u��,���b���7����zUiT/�U����P�~��V�3�ם��(��ݰ�o5�9=%c��X���h)g-�e��Hu��@��ј���v	l�hͷ�^�eLa�L����4�l�EH�һ��S;,��a�L��'ft ��ۺ̀R9[�\ɗ]d��[񒯶�8�����mb!��_z���;H�7��{;:��![��ba���`��:02��3����͗�H�ڢ�j)p���8Et�Ԗ)?��{i����j*�l��.��5��7*=�Ǘ'H��ԙfΒ���¯30�{�����$��Z8P���)�JYJ���z�w,��]	fu� 6���VHW={����}�����U̥����г�������Yܭ�7.��uٌm�:�n���loS���ski��L�ѭ���"ቬB(��WԾ�-�����!��
��@%���V�F��.��u:���[��/�	v���OI�r��c�q��h,i�vq�_!��#�k4JH��E�ԩ���{dV�\�sl���%�ޫxu�+�`9Gh!C׻��';�`W��U��^�����-=t9'@�����8��mպ�	�"�M��<`6��Ȼ&R�ea3�rL�%�\�]�1aݤFnr��:�j�<�����A�e��Cf�N�⻰�O]��E	R�w�:��x2J���ÊRb��r�ۆ�m�����h����;k�]�9�.v٨#
�F��������r����4>!��iS��+悺�yϥ.�m\B.t��2�,�J�f�%wJ�5��wn֋= j敘gn���Jt7���$�I$�I$�r��'IWbW%R�:ݵr�e�&��ժ�p��}�Ҭ�K�w"�0�X�;1������}(:枑H����A���=8�U�5�Q���"@/�֠�2�j�u:D#x�h�r&��73.�KWq�p�;攬Bһ�Z%gƲL��7�3p����C��#�r��\!a(j�ɰ��Eo�mj�r����h�A�6`!+�'�F�o9�؆�y)M�7��܌�yJ�h��u?�iLGp�kF�q��9);{�2ɥ����z��z)���0p�
A ����ue��6��ؘ�S8�d����$��κ	ܓ��2F+l��K�j���/z��R�7�r�U0���VLw��h�f�QT�pln������ͥ�c�۾̤gsj��f�Fږnrw���]K7Wqz���w�u옟V���wp�`��,r�=���>@B(Yl	��6h�0-�_v50�`1n������*�E�',D
�JvG�! �`��sxXҧT�Kj�R���V���Թ�-	u$�S��Z�[Q�3�ƍ�>�W72ό��H57.�k�Ȝ���-����\�UǳQo�N5�I$�Ls����|�n9
fE$��|%Հ> > ���)KmUl��QU,YU�Z��7�\*T--�X��Q�Z��X��f2�ʨ(ڍ5��Z���V89}ɎD���V�i�-(�[J�e���K�Z5kcFԬ�El�iR��ֶ���P���[jVTA�V��c)E����UR֬AKkh-Q����[�R���jT��F�Z�RŎZ�YXZ6U�J�2���Z��j�kF��)��1�����/�U��F�ʂ�j0m��{p�b�IK[�S�R��
�ZڕW��E��(Q��m
2��F֥�Pr�Q�E�,�(2�nT�b-J�b�%Rj���Pm���J&YW-r���&-
]S��b`��.b҈ѕe��Z*��Z�Tkm�eťV,KhҕkkUH�[h�c*.2�B�P
h�8�pI(�,����-eޜ'��U�Qӵ�70����3�t����ֳ�8�"�TN�Ig� ۺ��Mh��S�U"��r�PHl��>⋁6���Sٮپ��>��b�.M�f�F�U|�D�K�@4ж�1��@./�T7�N������4�,�۶������/\�0}�ZK���Qx}�xW6��zɼ���b�y<��t*�N@d-�@=�w������|��T���t�3F�oW6��;p�����̱u�ᄺ�*��� �[!��p�q[l�w�eN]Q�t�B��n�>�-l���{S�^� �]0�t�_m���'tկ=�v��C�zV+5,r� �����nN�8T-��s�����F����"�ޒ���)R��s������:2yz������h2�������P]zC�'Z���_��[�-�b�'R����Z��.��Cv����6��..�����SSOA~�J��q!s�ur�*��'h�ryh�x�Y�~7���mɩӺ�p⼸O�aE,yN�][�.̩����ʰ�/�r��4X6K�P����7x���Չd���9�_k�	�Y�QQ�������t�ML�W�5m�R#��[��+८��vv�73rGbQ��<��������t[}Ϟ�������_���@���.w���t ˫��h!�QtGe`�Ԇ�in��f�2�=$b����B����dS]'�O��<"#"!H�:�iL�6�)��t�ԸU!A�}a�wI�^�W0*�"�l�VM`T�b�?S���rc��X�G3G{�Z�D���8��h�vӌgG��ʟ�d�%>^�P[�o����,2�
PG	隥[��u� ?�4V�F�|�U����9ί)��_1����W@�ȣS%
��
���>7My�s�\ i���Z�^�z{1�C�2A����r�t8S _���(�|*�B�U�'ԨI�P���l�;[��,ޅr��J=Q��bJg&g�+�����l�	���%��fy��U���E�`�7��q�:e��P+�9��+%׸+���2�`�{te�Ü;�)��'&*��tdh��`��z��������D��،�D�(��R�.L}�{�֊����*��`I��ή�z���g>`�57��٫����Ɲ�ue"z���&���;�9�
�e�̓����GD#-`|��SQJ�K���m`͟�j)@#L���aɮ��� <#��i������<n~f�`�Gc*P�å���&�-\y�;so ��q��˚3�9{�F��?]"2�ʡV����)CJ�=w�燮�u�a��R)�8����ۯ�t_����Ǩj+n����
[3��%��>W���7���f^��~X�F���&��cӑ��qL��������co\q�W#囻�-�@Ѱ�ĆF2���̨p|�+q�:�ٽU�%�z,P�i:=9���d�o�i�j��*�W���Q�LW�����r��lK�*�W���(�By����=S��lz�Y��o���xx9�ӢP����|+����7�F�b;T�y�Q����V��U꘢)H�j\M�ƻ>�ZX8���� ���=v+h`�c�%���V\͊Fd+�%trNșÐ�7�<�6$J���U�w�������o,��Y$����Jjfs�؄�ƈNr(iDC�09L\HZl�&Tt�(! ��ƫk��{���'$�{i���.�Iw��]��������Ծ����b�����0+Ju��x�"q�øuձH��bR���6�Ko��j��}_�%�{)aOq�7и�d'f��\NC�{�xF.ξj^T��ht���	P¾8�8C�wB����s�'�F��0h0y����c�Ժ��F���)�7]�.r"dbt&gy�D&r,7�S�Y�����˞��|0�Q��YB��蘠U��	p��B����bA���\6�̮�ܞm�Km�|cE(���A��'��!~YR�h���6FD���iF�u(��{���k�H>�D{���F
�ʠ#å��x��v���-i+��Bs��v�${���G�[���\%՗'Cg�l4�'Ⅳp�VX�"���d���iWA��̈́r
��ط���bw���B0],O�Ӄ][CeOV��=�<���	���NRq'�5�SУ@��9ˇ����>wc"�DW��QDK|�UƂ��eBg���(QH����=<������5,�1g��
����[i�Ey���X�\�%vco2TX�Jd��c��W\�q���΍��&�}�	0���f�hZ��az�s.�6�;qۯgx	^���/Vvh:xVɺ���ܜ�:y��*u����
y��P�IK�@*���U@2��I�"X�BY��ե�q�3iGD�h����,�Iw�{��W��679���iV�ޓh�J��TN���qQj�D�*^�]���S�5��G]�������j"J���`wMT��B(b�g�B�?��]�_;�<��kU�g��Խ��i	xt.3O�*�+�R���1���WT���+�XtF̗�t%��S��uS�
�B�{J�o$�T6L�r1"z/�3�B�ED�q.,/"�S.�ޕ��^�ՑP$���V4Jt`�k�w:�u���]���P������c��Nl=�*݁P�q�c*��1�B�S�윊RCt"�1aթ���9���}Iv�8n���ܕ�*�˿
��ٲ�I�T8nl`��%������=��~��^xR���"h5�aߐ��
�ry��t
�1::��ɣrm�|�[�����������q�%q��_���X2�@Uw\!T�!;3�[1`�/�ݞR���	+d��Fi(E�� ��dŧY�Ò��u�yVXW�d��l�p�ڂ܈�E��f�����E\�]͗Y�0�$��j֑y��^N�A+�a��EA��a�2������sf+����;��u��m9�I�/T��Tu�uh�i�Gf�c(�=G�ιp]�*��a�Ԑ�>�直�8��~}z�m��Q�]�b���읎qb�r|�d���.�����O_e�-f-%"`t��V;m�9Դ9��π
���S�=�M^4���Y��c֧,ȕ��&@��Z���[���
F��p�d�Z.�9��\9���0��,������}pY��B�#j�wc��=YY\2�<�A�9�x��ˉ��x�$��Sw��w�%v;�G�p貜X��{V\.�����`�S��c��f`����ٸ�b����R.^�8��������)7{�EtMb0!�K�{����{}�����r������=��o�kC�[:W#�v�9T���ܩ�o�¥{�� �Nׯ��7�.�l��Ճ����-�)�,���(.4��% vZ�Y�rli���>�w��Ϫ]ΣઽG	_/.���=
|~
�+x�;0�s���/�wgq8��q�9�ؖu( ҧ(M��l( WT��[k���l+�	Rm
�6�������m�j�tf9��_JrpS�:�+1{���]�u���s��A�Z���΁ӹ�7zd(�N.	ۻ�d���J�cuǹl�:_H��E����kd�=�0��˂(��A,!���W!Hm�K�.��xxF�\�xЭ&�r��v2&�˶ ڧ �ȸ�j\N ���J�&*��k����������ix�B:��=C���e{���4���0�����bsn�q麙v�
|\�[R�v(�*E�����P��!�5�������8Aޯ>�a�9D{A��X�X�+�����3��g`C��|;�d�"�1�6v�`�'}s�>�{�)�
%��o���62�n����j��A�ؼ4�fӆ/h8��t�{��;3z��Y筥��p��{Ձ�GGT�W�T�R"��O�h���.���O;�-���.3}V�%���Ӆ���z0��S5q�15r�	
.�L�79J��G�zv7�����w{I��2��9׵p�S�a�.:꣧ �����}��D6��/j.�bF�j(q�T1R�x5ڇr.,:�ٱ�]Cf����0��*^Z��hU`⃨����`=�V�Ǿ�ô�Щq�:8�z�*Pג�1\�4��%R7X�
�:����]A��cT��� ���*vm���3݂	!�z��œ77��$M��KF�F�סǰo.X��xX��*�q�Vw/K�-�3ۻF+�Y@��^<�n�Jud�
��ĵ%��ᝅ��٭�;�Th��X<`\<'%@�0n�g��-�27֜�>!VV��[Cmm��T��S��|ks�Rо<�q0����&�( ^��W��>��$,h��9��T�K��&�A�+fE
Zz.�t]ç���;<[�R�����G���_P]&4E����*.�@�1�!h�]O��fɔ��5��IY���^��� &�#$���E�gX��"��n$�0dM��"�#��O-�=t6*ə��5�PFOE蹱�#�Щ��a3�a�����
,Օϖ�BN^�����A���)
A�Š��_�?^�^��� Q��:V;+�Vz��h+�#�7�S�լ_��,�	�"p�uw��U,�����7P��g������
������p�K"A�H�jf�i���>��K(x]��A�h�y�۞7�T^�{s�t=1/�����kت�Y~��{���D¼P��:�<�S���@䫞�����6�f�N$�0V�YS ��\�6����}����\S�|V��X=�f�ű{�c2	�����&�.݉��;��:��8���qݶ!z2tWcQ��qޝ��k�f�ry�uk��}^��[���%�B�_"X�DVmtX�p�R��c���;�6LO*Q��Pg"Z��ഋ���V��{wm��5I��`�\�ryD�k���GU����]6�1B���T�z�z�А�.LuD�("ؠ\��u�2:�	#֣"�ӽ�f���-��cx�t�j���]CM��������\�uf���j޿v���i���O�Z�=�N�]P�Lİ�^5����e 6ρ��~���=�/٩
�7̔<]o�#��#x90�a����������:hF/P��CM�N����'4yɯn�O���Ԩ��6n��X�H��9m��8�u���-�C���6��TKll�<�C���J�0�ʰ=I���8'[	e��@�cMK�ۋ�/r#$�UѲH�<�h�G�r���VK���^��4�ork2���y�)q^|��m7�+��>'A"�1�D*��eEJ��{�bS1R�e1�H}}�:��]֖�J�aۜ�mE��rCq
�|Vmݮj���-Aj��o2U�y���o�X��"�v�Z~K���w���/y�&���d�Ũ��I����"�UѬ��;��[:��Em �񅛩.��ŝ�>cs�� ������R�kԅ8����^N��^:Ez*7*/D:���㭾j���qմ�j�D�U�I�"h5�a���g��C/��mM��ꐬ��1�A����n/2��\|0��U{���D�r�{�/�zo_��?����}c2�(/I�E�⟶E�ݤg"�&w���A�j���k9���y�}K��T#����Y5��өj�����qa�L79]^L�DMu�^����U��"������6�hjy����fq�f�
5l�^�P'�r�;Vf���"2���۟U�yg�,^�R��r�=*�xx�{g��U)To��f
-�P���b��ر��k���@�j;@��u<�yv{�]��f�Zɪ���9Ӟr���5ib;}�.*��� %]mZʔ%�yЎ�	���k�n�fX�H��B�R\��q�<��
��a�Y�+bV���f#u�诲�=�{$�.�mSv
����[m\oJ�]���77����[8YCe�;���o�k;�[S��<�cGp^�W�8�yH�\:ժ�����oYU�5ؐJ�r�"����)��a�3@�U����[�fm�*��2��>�+v�N7�Y1V�x�\*5�2^�v�Xn�4i��Yz�ahTN�6^�K�W�¼�)e#��}�f��F����|rANe��
`=��&U�MhZ�
ћq]Ah@H�>K"\��åf���pI�h�B�i�c39o`�x�}sF�?� ���dZڈaZc�
��pzs��)Rܳ�D��"R2��	{���pŋ�r��X-���C4'��!�w��u܆��)&�r�2ԇg8��F��X{�%qz��r2#���V�{$�p����=��_]k�-�$���a�Â�J]�fE^�]���� Ŗ���@6�+U�Jͫ�'*5���H^�ӝr���=ɫ����&Yq�o+I�����e
v»�f����Pt��N�X+np3Z�Q��qL��<���6��2�폶�\�с���p�/4�Ir
�Z�^ԱG�;e�&��ڶgQavb�(LX�TI,��Ͼ@�ԯx%�ia�y��0��bb��G)�y(�f�ќ�h��c��`�ֳ�V�NV^Y9+���I$�I$�I$��K��Fd���
u�6����+�uq:��Kv�l�r�o�WM伆����i$����eN�z �p��Q׸�΂�eU��g�s�YQ�u�����<�ζ6�`�R�E!e�T-�=16� x�1p�ìT�0JTVI�kVY&�'��\a�!�l��	�+0�=tX��/z3W_�'	�Xp��/q�����l������d��er5-:��,��u�_*�NQ�Ʌ��澎�pt���Z]���f�ʗ
M��k>���RUY���ɔ��/K�j�����k����E5�����P��qZC��GQ�U�Zٺ���Q�5�r�+]�7H�̣j�d�P����g��_c/��V%��4K��o�8ba���Ů�Ed�=��Sn�jiNt���v�N��{%���c���ufI����YW�f��P������nFZ�����Xa^U�Ě�	c{c��g,��,ћ}r>��ϱ�mI�)��&�����2*$[Nv�n��$�ٷ��ߦtTb�hUթAbv��Gt�w�pU����-)P,u0d�,�ұM���ӵr����ѧ���OK0�����6�=�ɣ�[�^�P�G:�q�����r�Un��\�i�9/��Ȫ'�f§D�i4��2C��䈧�F��&dRIee���T(V(�̣�-V�[F���������e�g�*(*�Kj?�Ϛ���KwCb�0��o��"�*J,YR�"�[*T���=��{Ѡ̣�a��V��Z��V,ۙQbŭB�EE��J�T-�YmQJ�Y�UPM�T�X�h�Z�h�kV(��QFڊ-e|�` �k)��g�SF�+Zy�b��=eM��X�-V���*����Eլ���-PGypVT�U�*"�­���Kj[j�J������hZ-��%e�e�J�ۍʎ�U	�R��clQj,����CV�o��2�)KC��X"
##h����g����8��e�FE�ԨeJ(�--�Z�Kh����֕�����mue���T����V��L[UYDd3�_�צx�ϬӨ�����P<�s���&+��دH8��ub&�msQ5SY�J��g	Ӛl��kb�I�U_}�1�~��{���w���<��7�S!�E��
TM��ni�&4�����Ob[��o��ha'�;A|���C�l�t��7l@k��evN�l�2����k�,[��C=]sB�x�2Cb����
u�Jg��D �c]�̃�P�T���۫n%�,��pKR�H�R�e���'#�z����EzTX�5��,���F�Me/ǅ�qmW	C|j �xI���E�b��o��5a���B�,s*�d[��]J *�t%C��'{3�k"�ӏ5�0�J���d_�;:E�!9��F;�A��?���q�u(t�r�k5��!���9�6���Ŕ7���F���}qX���׶�2,ae����7�ۢoci\�͘��g��=�L�l�5��[c>,�`�yX�����ꕊ� ��{io�8��9k���)�H���<?y�.�<�e�3.vS���`�t�oJc��^ީ.J�ik��sD�A�G5<A��2�VX����͍4� �d�lІ��k$�١��-���[��Fm_h�{�Ýѩ�u��Ef71��@.�SpY3�eRN��͵�t����M	q�������K�vXՙ�F�L�t�͌w�yN.�/'�3�W�g �5ra!E�靜Av�r�4g^g3� RUР�:����7Jd�x�zrT�Y�X����z�-�b�ku[�j��\
BGC�Q#�ʌR��]-�P�3�'lJ�j��&gk^b���X,��t��J��+�w�=��n画YU,�b%��ln����s1��:�HS9�To��BUl9����st�0l���ҍp�,�����X�n�{�6�fZ���T�Q����Uζ�y`�a�� ��4�Si�Ou7�x���Θ�)pܘq�]��A�.���Pd*���Zz/ԫ����2�U��'�/Cv/wr�򲭋�{ƻJC_y�U==(3DW-BQ�cV��Y�L2�Z2jvj����..8d�
�;v&N�
�pE�s�S���%:�BÙ�(S��NG��0�O#��;Zy?d#K��J��:��(*%�zy١���V�'d�g-]�S�e���eU�������T�A�����ح��]O2ܦh�I-�L}k���<麛�&K��gG����d����Hů�<�KY��*���s�T&�J'��tL֢?.�v已������௬Da�} ��(�*X_oM=ohK��ԗ| � ��I��V�b���tlLU,��m*� �ִ���gЯLHz���%i26y�=\��g�c��IJ��=��t=�u�oJJ��)������ �.D]�m^铍��%Gs!F�U�sw�!���Z�LM��(����b�F6Hk%h�aM�٘���q�.9U�ߗs|����+.M�TkU1��������޹|��l��j\l��r��T)H�5#\�h�������	��K�3z����aXu,�#`ܱs��茍r��GQg�9p�Yz,�R=�kieέ�੒W	�Q:<6z�'�c��Avw��~���g���0�V�S�Q������)��\�y`�'G3��<J�LhuzI-���~��oM�ش�twø�´W7@�Ö�s|8Ι/����cJ�{���Ef�0i��>�1�m��g?Yb�qh�Ҩ*��ֳ�Тu_��h�\2�I�F޾�yB��ꎅbrVE$�V�
�h�"�C�>�N�7��4I�2ʠ����-;�y}r�s9��o;�h��(�W��gO-Ig���n�mjN7����,ʗ�:H�^X�v)�gCTb�
���f�G�V��o\t����1�`�xzV��ɸ�L3	�X.�'Ƨ��`��������2���::���F��k��g�D�c}k��yV���N˳WL��c��7��7ɜ+��ԗ�Uu��-RD
cC�h�;- ���8��jp�ٹ=�I��ʕ�r�C���7�^%��^Aa�6%�P�:GLgwc�:6�ri���[��;y
�5�f��%."����<����C!Tl����ƙ��=8�`�¾�l�A��H{�б+���4��� ��B�[���3�i��}�����5��U�R��OW�A����o������\p��I8&u��(����/��ȃ��D/�1d;t�꧟���7d!	�P�*5���]�p����Xٍ�4��\z8�#`a)�^�ż�0.��o{=C~+< !	߽K�T/~�X{󸞗���E�f�����zT"4��[�sE(�n��nt�w+nlT�^�祻�S��'tг{��}�_~�����*�/���[#x�L%Y����Y�݅�ȋ�W>v���g��ŭ��2�u%߇����6ڌˣ�)`�T��VT2��DlzL�eKS��h��X��t�]��S�W'\�(�nY7���,)��}X\>S])u,����(\PJju�&͉�ޘ�ԓOv-;�a�2�ƺ�65Ӌ���PUi���y�=gQ�_�G���Q�^�5�9����8l��L(��r��Tn�c����� qy�с�;�t���z,�'�Kz�j�r�:	�'�b �xs��5��M����|jgv�)T�u����k��,��r�x��,���0��ƟP\)��:x<k�Қ�Z<9�N
s�U�q���h]��~\H� �+�Q2C~��隧[��]tw�6�	������~xM1:��2$���Nҩ��ԩĚB�\'f�k������.�Je�cz׽1fC����!���?P�7��P�� J�̡T�9Ac���4ͷ��ɹ���/ŗ���&Zu11��t9L�͵�RiÀ|69ڎ�l��n�l��®sЭ2��(�l�ݞԯ�xh==�M]�G����B�B7p]l�lCZ�	��^s��{{k�y�2��ː�i�EG��#����$lv��.,ǳ���j�)���2�*�M���G^���ʼ���S��
��#���f܋XHqy��(@�;���	����s;`��of�{�&�´G�xZ`��`���a�F��e�ܱ��`��p������z�k����4�e�R�q#�,B�bٞЈ�]��B��iX�g/�C8燨��vo������b ����O����/�m�; ��*h�F!WH�G����M���:�t��S�7�r����y=����g![rAڠ���e�Ҕ�Q�̩by�e wl���S�&���p�g���*7/���<�S�.s=��U��a��tS�5��x�|��W˅��*�n0:��QD]�t���M�;ys<�,���U��΢B�5�+��;Up���['L��kg�)Zwެ��0{�裷�U��������<R�Z%E��
���|F��z8�Q�t�p10]ᘫ���
�(C��K����;B����Ϗ/	>��F]��y�n�R���*�+�%\*Τȇ�s��W�iY͜W\�9�*cM)��\._n�[��Yi[9�W}U�ui/���O8��Wh�n�fnfc=�H����+GQ؍�NW5GN�5ʸ\��F�*xԋ3�2���VId����ԧ��5���X$*��b�.<�r���P-ƚ���n�;�X"����d�W��Tc�
u�yr/�k�w/�1`�:��yhU9<&������]����FT�f�{�䓼sa)��p��[?SP�C��b�[R�pud
J��V_�v{ŏ#(`�����V^aI�6�r�;�TK�0eE�1����g�4�b����n���LT��L��y�0�_xh�����M��}I>�t=�2�].��%m+�b*���N��=i��H�K��8�Ox�ܱ�S���@
��d�t�f�h7�,�]{�!�|mYW.�M���w�Z�]D�5��s/a���@�Q�I�E��$5u�V{�{lD8^G%�Z}P>�fq�]8�!p�&���0�_�)ÛG!�.>����!	�-F��`�y��@��vEkx��]ri���w=��P�c��J�*��T1ʋ���NEe8��#�t�B����ޒ���E��\_[ءѾ�B��}�T�=
w�rM�Y�=c��SR&�(>h/�}�E�5{Mw�k6���5}+��t��%K�Jm�� ��8O+L91Xݒc�ѹ{�J�vv=���iI�\�&O%��v�b��Iw���^���f7����r�6�+���I� Vф,Ut0;Ռ/�`S�Y6ǌ̯+�$e�ps����ł�M^��V��R�t�Da���(uoԖ�y�yq=Հέ�n�|d��<����u�Q�<����W'I��^4r�'l��Z��wR�_.���x��\+>�3��kHP���qH�}�i/��s��P����4��df���6��L嘗锤�%D��.)M�ːs��1ig�n(_���#@�B{�O8<�S6�LG�>UP{Po>]���
@���u�u���q<�[�l�g'q�nE��<=�x��Q�p�_�˄�c��xݖF̋��(�7�;��K.��ެ�éJ�l�Z��^��%u���"��x�ຍ�����E��ݦ__�Ͼ�FbO�3�t,CS0j'6jd�
���>�%���|��]#ƥ�����w}�r�.��0ੱ�j8�!WPb8�����9�L�l�T��;X�B�W�,ވ�0�b������JH���\4%��f�qQ�=]N���G7�x��W�>��w���'z
�(�����2��.A���ZA�Xi�9�Ґ��Nr���$���b!�
�Ig��wU�kEɞڟ���N4���|0!�j�ۻ=f�xY+�@��R���u 8����7���qz�`ؔ�y~u��n�*�.��f�X�H�}�������o����+���Q:ܤB�Y���?���>ä!j�%�b�5� ���j;WR�;���6�P0���v�p0�u-yz���y�L���ɯȔ顬������H�W�_+�)�����Œ-q�z�N��_�5��r���[����z��2�K�q�'w��Qй��z2>�R�
��6<�P�o��7�7�)�Qf�f�>���>\O�����:������jˇ�xŉAGȖ��L�HT붚�H�D���� l:=Du�G�Tj�s�\g0�]@{��{P��%N��G�y"��w��"�[�P�{Gh#�N�t�\<�W#��ҙE�G�(��Nu�j>+���Vө~�\�b��`�_���9�N��R�a�\�|=)�.�Jk�������xMҠ]��Ȩp{�T�|��{#7��V�������sp�O�)��t�v
G痁n�G�owClg*�����2�˭=��x�٢��[os-Z�yQ�Y��,	�fhz%DA� øJ}3��t�(��K���6mo2��Ɋ3�e�v�����J���ߩAOLש��)�<6�A[�����cq�(Ɯ��@`���UdN�V	��D1J�L�4	���>'�\.~,��3<��ݞA{��>ɍ���\%�D����#�u�<���ʦ��
融�{k�Ń��J�%ƌv�W�����E�J�GQ�Jg&Z���뗪}U��H杽N���P�Y�ؽ�Ɍ�:�M͹���b�P�usC��P�n��䗙�&v��B�v���Ŋ�^v��,�V�`>>x�����G�:^H���~1H�+�`�Ry����;��:�;7��*c
��Z*�n:�ц���lB�Kou:�4v80dtDt�3��lj�y��WGa���0�b�vS�����s�<!��t{go�u+b]�~��
�}n;���OYڛ��LM\�h2}���ۗ1v<�c�koG�R�רGE�2w��<�*���|v�qY_R��i��5`(3�����sd�\���=O��mpa4,����ڣq�y �,�uǝ��������V�q��]"3���1��� o�Gp��-WQ�=_cڟ;voKC��PT�n,�]��:gE��Y����F�+�k��Nb|s	��#��֧'��!�q:
�{y�����������Դ��+��l#��j�O�)��c�Tv�ퟬ���v0-܍��7��ü�ٲ�\˲�ΈWʖ
��9������2@���{}����g	rg�r����S!����%a-�FL��:�d
�N-ӛ�խ{��v�Ƭ��\��Z1c/�:媹�e��6��'�uݴ�\���LQ�"����Sr|�]��=���wW��,��).��K�tWjF:]�dԮ��OAqN��i;|�ͽ�6A�Qh��B�T��QZ*��<��2�஥^�Fҭ�\��rgq�D�V
�x^<9d��W��D���$�?+��+8�nm˝�01��n�تԾ{nw4�;ƻnbyF��@Gs�L��97��)JJ�����Ыۙȅ��j�\*r�c�*�P�zڔ:�@b�YO1���MJ����u��7-t��rV�f֊�Xx���A�ѾW�R}Jf�-�⃵��n�8��ջ]���g�ǗF�n�m���I$�I$�I$��nM��%�n>D& !+�����2���b�5E������r��i9�ލ[F��#��U=�ɠ�8ɘ��A��1�h�����.P\�W�mH��p�t�!�c��(���}d�Ҽ���7��Oq��Ir��m��K������)q#]��R
� �]��aV��.���5�k�C9��h\�#�wwۀf���A75��l�T*�JV��G�Ai��*�D�����Dl˫�,�
�rQ2�Q݁����!� 3	H��X��'yS�!ހ�gP�wЄ��RZzŗ������)QY��0v�{[��+����:�	4DK�Y��)��Xx��vٹ3]�Y����:�����?��^�2�;Z�%q/�
�P�ø�F�֓�]�e��h�'k�I��!<W|4s����4t���gl}�pԥrݲO�
��o�W�+�e۠0���HnVk$�ۧ�n$����MNO�r��q�W7$��:����Xӹ(f��m��6��Y�/gpF祉Z��)�2��J�Ᾱ�pH��aՏ��G�Rn�k���"Y�ʔ����t����bn4�jHr!-�䈭jF�P�2F�:�6�'���t��Tb,Z�����(Q�je*�Y�EJ�DE��DA��[b���%��8&F���@WMuB�b%��m�V�UDDU�*��U�ƈ�-ոZ���\f5Z��"�Z�b�Yq+党��\���1(�T*-E��֕��Ƴ%l*�[��r�ƕjm�E4��Z�Aq
�J[jAĳN�b���H�~ִ�mRƻ�*���AE��X)��E��&�٫�ȡU(��feD��Ŷ���L����Ee����ӡQ�ib��N����>�QŎ[�����,L����*V��V�"��ڵ(���+L�����j����Q������6-,Es.U��Rۗ1��1��U��L��ڦQ���kVcs��/���M*ۖ�j6�s��n�VU���^�˃��]m��*�ٙ��y.GG�f1�u�Wth�nn��k�9d�o-�4��bq�j�Z�{������{0%t��q�]����Gi�Mx�
�_�VFA�E���:�8��H��
T[�ʇ\�	I1�T�����hO���G���Ý�%��;L�>U��]+=�6��9��Hla����{��Z�P7d;�*�F�,b�*��z��\<'%��Ǝ��^�Ů�Ǚ���⚎��~u>��3���!Ş%��~���r�B��J��1+C�(Ld6��<��0ƺ�b��A�J6�UJ�I*����c􇊣bF��q�7�{��j	����k$Y����:�0�L7�*v��t�`��YED��ҦfMڍ���)Xe�DWx��{��ٵ�]�ҠJ2"�dd��r㥓�9����9�vt#�=�^�u|0S<N��#��W���w�QM����މy��o(��9P��e��<,ed��6��F����z��zOK�u��;��j��b_��	�@�i��|L(��pD!����xz%Rˡ���~���cǙ�h�ǻu�e��LI�9�^�╬0�A]wul�W���K�8�)W�����k�-�G4��`�(ȝqE�Mzt���i��.����nl��'!���|?{�?x���VLv)�<�/4�8c�:ZL
>�^ċ���Z�fkϲB��q�&���k�`h��e�F�9�a�nR�6�C+��/h\djZw$�=9.�w"�%=�Ի^&�nqCʇ�lK�>�X�6�)�W��k����<:`��yC�N�sonud����>�����Rѭ�b�#��!��8� '*Ut(;(��'N���_�\�j�9p�~��l=dmJ��0u���Q:<2��h� V��w3�rq֕�;�Fl%��8uj���X+Ur�4n\�ꔖ��(H��wҬE�T����j�R��$ءj��}Sg�Z�{4� ꮙ.B��N����b��'X�k{���n��3R�x�=�AWŌ�DmM�X�ܝJQ=���q��'A��I�[m���|hW�����s�j\����9�3Ƣ�:�t{�v��4e>�$|5U�u5�pY�H{���>�z'��u�͙8 ��.U��O�s��,4Y�B�������y�r�M��f��X�'�B�w[(�r9t���%�{@�I�`sL���`,��^���g������9����������V.o3J���6�ؐ_��B���{���7Ns	��#��b�u%߇���<�m��t����
�||��?���\�� p�o�
����0���m[���ŗ*�^J��B&�_���B�8��)�\Z0��U��B��nM��x��s=��b�aTE)#�tI�ņ�#<�L]A~��_Ժ���fD�^��֯���]~y�YBw��V�0��F��f 븆"HT� Pj*�$�u4�ņe�qᎼޞ�����,l���u䎛2���P�Q�����̖����t:���J��b%�w1Pw+aߪ�I��#la!�8v���,]1�kg^��ǁ�������೟�L@���{(�W�d=t�2�yx`�a`��A9;	�뛐�S`��w ~�5s��������:����ް�����h���^��`�hWA��b,��7��XR�;�	\��dA쪚|k��=1O��ҵ�j����6ϸ��®P�GlG^�ur�e�@ʇʜ˰6�9��B�Z��B9n)������GP�B��d;�P=��t�p��w�>���$u�2��p|R�2��&�*�ԽSCƒ�n�!�D�:]�o�r�`�itc.���ˮ����L�M�]���[�N{ȗ������:���}XH�h�c坍�1��
�@��Ԑ���]���nu4#��b�(S=���S ��� m$�j�g�x���-/S�{v���!����z�ez��L.��zeE�U�uˌH5s��Z�ڴ�����KM'�Iq$j0!�O �<� �'x�������:�?�9U�&����s
����z��kv`1������V�x�g�\=CI�僌�0ή߇�[�)�KL�r~��b]�%�:�H�Q��w4)PS-�\0���S�/��c�	/�������<�o�E�E!�Ꮥl�o�
��>�0$AK��*��ºeG\�q�b�X_se�B����|��c�����:P��4:�~�3���y	�v�'᳑���U�~��ڧ"l*�w@������A\�C��(Ij��%�f���f	�[�E/��m5���Ji\�����b�P��=�weά��<|��$�R�ज़����?G�,ez�W��X=���V��&Z~�i��Ze6�l����ue�j#H�bdkܚ��+�Wݵ���O�^G����V� �N�kׅ�h3�/�7�[桤T��QБ���6��NM��U��n�6�+;:�K8����'J�����N�����Ʈ�=�%^u&�����r]���$��Ր,l�����^{Y�.�q�l�A"vR#���/���	{�&��RY�]U��K�VÈ�Gj67�O�cl�y"ފ�1�+�u���uNR��l쉙c�.,a��.�l�r���z\nsV�To:Ȣ�V;E�v\9���X�A�U!��B�����k�#��6�S6:\[�P�D��}Y�Z{�e]�z�Ys�o8/WJx:|��`�]F��O�֋�k]_>%���~���ཡ����Na�z.x��D��j���|ݸ�5z�:"�c ����=K����:P/7�|��D��Ֆ�.���K��"T��E�jZ(��.�����iQ������&dl&��̑3���8s0��V��7{L�_'xg<�#!E��s$c�|�p����S&����O���N2�/ԏ�	^,W��1\�g$��Gdݢ��K��n?Pr/6�"m�ز�%,����ؠ@וǤ�>*�x)���Xo	�ܓ���X���*w�D,R#���݈�i��ES���L*oR"1��y��[yIe=�
Y��`PV��AS9�-C�ۗ}w}{P�	��I��;��.:�t���;�M���^�[Ďaef5�T��("�xl!|�v�]�պ��f�+���
����k��a���c�N��JR_{΍����^��-����W+0��ٔ�gV��n����.a�!c��}��(��4�FLT�s���wM��j�Z�Y�{L�2� F����VEI�ą���h!]����\T�=��y��E�������ތZ�AbA�cSR��*��5�Б�|m��ӳ6:�K�8�Y�\=���l�0��Æ9TC���G"�$5u�kk܈*��"�0��{��a��#¨��~�NO�h��*�9��go�H�ذӹ'U�fB���<�����9��\c4H�w�o��2|.\6Jc� �҅*���b=�7��'�Vm�����Z�6��m��Z&��S���N��L+E4/�]��C��<<;�ʭet�0J�e��4J�c�w���L�̇CS-{�r��wꖂ/�=3�@�cW�.
p���;s*jꮅ<��Kb���x�Ty�<�97P���q����}u܆v�:Nv-2�7Hc(�T�y�2�D��|$�/Ȋ�"��v��^P��&3sw�D�H۬�۷�\@��}�C�:�I_t�}�Aٮ'!�����y�֡�M��&z��X��A�Q�~zf(Gl�k����ٗ3A����IZ�(̵Z�m��iA�K��:�>��AN��A�օ7��b�qh�ҴӬL��]��.�r�X����}D���k|%-S���+�)g�^�0H��!=8��%���đ�WV����\�B��@���2���*j�
�̜0j��D^{�w�;����Q͗^�{��o��p*�??��|Q�R�Dn�@����mu]EW@1����吖��6eS�w̜@j��W��	�f����":����,n�Ez{�F"+��n ]�-���N��DD�\K�Ip{F�W���rVR��6�S�;��XhM\
��0MB <��W�v�^ WB�;[��f.t�al�+u�Ɍ����X����t0�����rj=Q����٘���.�[�>�h�Z3�����5��9.v�ᄇ ��P���,\��VDUǞRw��mg" �qn��L	�5�k�ݗ�弑�zTA֡$���]y�n���H.�����9�g�����]\�4%q=��ld�wb�}m�Vj���+)"�ee3X,����(AٶPT"֪�J�ވR�?�i����@�w��~�������U,�^U������6ˍ����@T F�e�ޞ�[���䉾��p�B�j9�Q`=gt�n����L�^
b�=m�a�:�����:��Ǥ�73:+< �h{���ʱ���.�XQSj���>���NjF�v�DfKX�y��mY�s����̜t.��St�tNFC��Բ;�}sO��fM_>�&�B��KC�\O	�W�+<� ����,z 53ڲ�d��Þ�ȧ�ZHXT8l�`��PB=Щ��Gfz�r}��o��f�]ז����[jR�tC�0��|���8���F�5�]}G��Qpؤ�4Lev�q"��_B)M�Q�l+o����/���'ք�2
��|�`b\�:��j�6b4��JL+t�uب�ٛ��)��.1�s5N�)J�zV��z��� �I�rx�s%T`��ț�>��L�"HҭC��w�S�"
4�!D)�|����QI|z+�/M.y�,"ŭY�=T��w8��\��u���ʏ���K��"�Q�v\a�n�l������MfX����Mك�]T76�ח8tc$sw��wIi�� �zwR箶GX�Ҁ(vb���Z���Z��,~)�x����ᰋ<.���3Ă�u	�&x ��ҷ�މ��T�`���;;�>���!1W��EE��*o�1Rө��P�(5��n�w5lK��t+�u�J�[#�m5���K/O�z_�\J��g�d�[��ʲ1G���F�>�3(��0���[��A+�u����3�!�}�M<��z�T��Ėv�r���9�p�k2����:ϴ'e"6�T�����,$zk>��s�Zr.P�[��dx���S6��|�z���s���/��c��P$;A*����:�+�E� ��J���r��1�K�������إ{f�Ni�ƯwS1m)�cE�Eq#����&��e��T�O�x�״�����)���KF��_$cu�p��|�/i:,O�ʤtR}T:�8��؊�>�J1�F�R��s�ƛ^nR%p��k����_U)6��h��t�#�v��v`�.1�7Y�F��wj��s�Uǣ\��VL��*�b��>ֵ�a�J�|Wo�uJ��lY�畻���w�Q�=����otu�k�6�fw(��]�K$\̇]oe�j����p������m)��[JXzF��8��Aǐ��Z���m�	w\J���є�ʷ@KC�~���y<.�MF�=�iD�C�����x1��ț�q�
�kG�s8�!!:"fŸP�-i�S��s �8���^��+�$Ńǆf�8=�.�J�Bx}!��:��^�ȺSO;���G�+&D��3���ܸ�,�"�j�d;��!���/8q������̸�*�����HW����a���2�T�����
���WK�V݇q��������~�'_�%�RQq5H�� �G�[2ύ(�9*1E��Xq�yW�ϗQ�0�?l���B��L���n<<;��m+��&{�R���P{]%����⡎�;/:�)	!L@�N�']���r6Q,{�!u��������9���%�_��a�h�0pZn��0��Æ1TC~ڨʞD��XwMg�����a+�[鹞r:��W���j��*��DdL7;��0�_�)C�WWrl5�B����}&��+/h�Z�;��`YR��h��j�mL�/�Ka��4��sQ�bN_�xR�\��8�o�}N{���z�-k�U^�ݠ�k2ܧ�͌wT�Vǡmp0��- -S�|��K�ОZ&�	l�i��p��i��V��Y�.�[0��/p�2��mXI]s�I�_=Ņ��>xvf�Z!�a��%���8ޕ��YӸ�Ȼ%d��C���EZ�!:�Od��`���ޚ�ܷDIԶ��gs�oW]sw>��qo<�7J�^�����F�N5ݪ�F�:�?[M���T���
�rjUz�e,8D;��/+��>��Sgr�J�7v��)�QV��n��ԏ"�p%��op�ss�"�u�̥�U�+�qU�hz�����M�.�	CX��]tӖ����:��K��Zf=�I�w�[��.���Z�7@��	b��u)p�4�͇�ERݼ7��[Q�گ�+����j�^u"\hU�۳�&8�cO6�3"Z���3۱�?K���I����/�fm��*<���T�w��[r��r��ut;��f���P�\ǉuw�k	�F�}�uepR�YY{���%[|��5a;}����k.�ne��U�f�
t�Sx�W!(�3�-�0K��n�%��BsNv_.�Z)��4���N�5Ύ�W�j'H��S�\T�I$�I$�I'GDG��(v\fv����.k��wW˥ՙ�%�[��� �@�-վ��1�`�5���p[�;�Ś�Zr�]�A�DG�N���@-�הESo���]Gw4��d�L�l:���0�=�m�'W��y%�6!�̫Zʵe>�:�Z#H� M7F������@�m�i7.���-IL+��J����٣��w����A��@#7UX�
��v;3��8�!�T�=9�`�!ٶ��{����׍`��,`�FP��%��^��%�;o&hStxQ5S,�6�;�hƴ���A�o���	ʮ�V�%�.�PP�0Z��1�ɔOPԎ���`��h_'C��mB���H�H�w2oܳpi����į�dг3E6p�;WYf��dt��xo@�(�T�dmsx."�7��ZقȒږ��N���Uv�J,�I�:�񹼧5[�@�k�1���U7Y]}P��՛F닾x4U�V2�ٳ����b<�8���A^�¸��K(29Zq�1\�w\��)�U���|/[���)$7K��RWv\Z#��VE�>����v �V��K��	ā�br�m�ԊdRNM��0���������߫�	V#s�h�,��dGY�������%;�4 1ә�T�MZf�Rڛ��5�љ�5�ж�Q�j�����W,�Z�ֻM&(�%��W{����Y�,��2�ް��U6SzP��MRQ.Q�"��3Ifڨ9j(����4e�q��}��~�f�3��.�8�O5�ˉ�H�)��0��
��]R�괠���Z��fQ=�"�0EPE\����I6�M�2]�
��-� ��.����ED��F��E��暍��ϻҪ�M&[X��u�a�t�(�}�M"~�M��(�V�T��_�.YV.!PC-X��ӎ[*\Mr�B��8ɧPQUeE�d3*25�J"�e(*:�#����4	  hV�|#���x^B�+GRww����1.w��e���:TL�@�/����V�ji���g:�[ �N�������z�,��4z6�0U/�g�·>1��N��A�.�*�Ų������IGj�sp��PS��ao+�#��}�7=N�:��S�9<,/�������B����A��@���/m,�w�T��{X�D���pE�]!vR��SO{a�
C	�
u턇�Q��B��8"8�ﲲܙ�V"O*�^׆O_'�l�=�oD�yq=1T_.��^�B��t+SOf��U�%�P��T����íj�P�����	�p>/����:�|���������-x�~�OO�wl��Qf���V��W��B�ռ��R}|J��u[�UgMӡ{i\��[����f'��ӗq�]�7,*'@�@������']p�����5%�ISo���IwH�c0�R3��n�7Q��G�'èY8�Q��e�./ej>.;����]OV��#�XKָU�Ʃ�аQq0@�	qa	��3�b�me���P�+,������1�O����/U�%�fn�v7v[��T쮭�`�YN��ګ�}����8�u�hpۄ[��m�>�"��sN{"��V�|��|T��*��Iq���l��$� ��Sv1Pi<�w;��\NC���I=�L���)k��xAz'�NT� ']}I��!20E�M��Ij�ɤ	q�t��q;]Xm��6����6]	;J0A���� UD>���L���v���3��b�?B9���|��_T�*o$�t	S�j[����y���}s���!x�ϛp�Zߩ�{DgS�/$=b��B]��,dm�$8eRnm��ۊ�mU�hΗ��� }���X��z',A�$1�ELP����n�do��C���=�;i=j��h�Hމ��UW��8#z�u{(��5���ku
+8%�����t�fI�C��}��T̀�:��ܗ���R�ׄT݅
q��K�z���g=,�6�tT�^Ӈ6�ֈ�17�9^���.�6|߼�����%B�&(P��a����6�l<Tʌ\[��	V��G$��+0�B�О�y~s</j���H�OPB<��L��\vg���9�t��g�4��p���Ĺ���Սf����ݪOF��]�_�
��j��zZ�sV��g�Dp+ΙYMͭ�q�jo4J��m��=���ev�hH[��Ru���j+'gL�G���x&#P��)=�$���F{��KYb�OP{�H���c�h�z��� �&�[��>����4m#��Z�B�z�(���*[�m���g���K<������ネ����ʑ��c���׷ֈ�xs>#�.�P�ʭ"EF��ă�݇2����� �����K�0M���~t`�Z-�ةC�bQT�H�R'qRKnbu�&�˫ڿUe,'�z����sP�<�E�"\dM
��.,B���"�:��g9�Tq��ǈ^�*ͭV4�;�q.4w�'�Jx�d#��d����W�,o���ל��w�0|�/�k²���2X����k�*�Ud�̤�l�Y-�H&�X~t#���;��{�����B���Ғ���\J��WK[�Uٻ�i�:%�?vO'O(����]�f{B!v�!
r�x[����K3�K۞��Z���9�x�0U��t�� ���Sz�,�X~������j*I��y�b�yi�\��wt�Y�:����fe�R�ھYt��\kN�n��/%Yt���o���,wT��Ȗ��'FN���2U�cn�~�$̳ŝᲠ�s���;%�4s�$5 �ս�U:��tk/��$ިܑ��������	��ϩI.��#�xi�͕8f�p�\	�<.���D��4g6�Z�vO�TK�!�zD�Pq�5@��eؽ�s'z�7*�':�՘����(r;U:��P�1����4U�}G��5�5�4Cgx�^��:�;����h� �͂w����ς�C�Fң�x��ZZ<�$+F�gC9.���Y5Qр*�b�B�Y��Uw���oh��Tt�ʷ@KC�ƀ��m�￉�Tn0�x���7X��=��~b*�d)y�x�P�F�<H��d�}�F����<X�x��8�eMPW��\�d�PR����τU$i�LFU<��z�Aԅ@a�TfD���xL���%/SV�/�rM�J´h����v۾Cq��z�>>�+ϐ�h�8�ю��S�tu���SW�����*���Z��.p�:%(gül&����xJŎ'	��@QhX��MΎ"ĭ�s�5������σs0����e���͕thw�v�=�Z��q,��9m'uBѽD[
�wq�t�R��7�R�wtb���#�Z�ٍB�+i�ĥ�+��6�ID�i`8iq���c/�[9t:���LT��B#9
�g7a��AC�m+��i� z=Nd��R���0��l�̝R�be���P}����Q9�B����?z�>*Y�����;�S�Jx�����J�c�Ū�t�]�7��L��fU\�ф����s�X�Tķ�.�c6\L{���w$���a�Eg����}׼��=y؋��pL�Ag^���`=
���Yk�°� �#6����V^���-ǩ���`�ۻ邯-@����3C9zl-�:�B�r�n�2��o.�a<Pw~��׬xm=^�<<u�6�t�!C:�b���<;ωu'�J��qs�)�r����~/��H<{o`U�7�� D���P��/-�f�Ur�{u�ӆ���S[
,9qEҙW�U�J���x���86V��+��R�s�<��X���[]7�A^��@��ǌoM�/��� �ZfpMe��k7X��Cq�M]�=�e���Wh'��=�Wy�J��uM��A���]|�)�4�a�_ו%�wI�D=ew�x�$rn�N#76�rGEV�n�m���%���jn뉇sz��5�l⎵uzJ���� $s]r�o,JH�Uj����ƣS�;�=���DO�@��fwK�0��x�G���Ԏq�P�u����}Ԣ̞tb�zN:�
3�D�^�	�7Chu2zp�*k�t�4�xu+��]^����[EH�һ�%:1B�8�."PBvf�J��	
4�m�I;�u���4\��oJrH,��#M(�����ХN&0R��'a�3���������+��p�^�l�s�Ku�$Rbøt,Aj��KR�A��=�+�Qi��q�<���߳B�u6 T8�9�(ð&���B B�+��1�^om�=���;�5�4۶%t����#,��*L�������u:���wPQ9�z��ua�]n�P'Y�U�Em��O7�W�W�U�!V62E��{��'s�`e�ɶA����G���VF5���r�\lQ����r���|�j������-�J����+��+���*��b�񨞤J���1[�Z@S��j�I����)��u��L��Ш�ށ�聛��.���ߋ'�>F�J��6�"�xP�y}ʹjs�b單@���OU;�i�r-������*Er]�=˙�-�Be�rI2L.kԖ����_T�[(���ToOD�\#��"�s��O@}/n��=T2���TF�;��o��{�ڛ2�s�у|+��t�l�s=��
�t"�q�z2.8�CWG�bg��umʩj��R�>h:F�Σ�>��O	X��'����b���Sr��obcq����n��5�8a#���]C��W��:����˻-U�����Yu�F=�0;�_����u��.���v�<� ��Fz��X�w:���|�73N�m*܌@�U2��]n�����\S�^�d�	ܞU���W�ֵ��o�X���3�EI�5=�qT-"EB�TbAh�2[�8�b��-�p���S,
��D\�$�k�S�
�h��g�����DR�DDi���v���F���[�Q�{):锰�I�o�C3%���ݿ/>ž�y;]��$�>�_v�C�q�`T�q.�Su�+U����ʊv�S����N�_ݾO�1�z��v^o�r�0�|AN��;؛�d»�0f��Ѷ�@L�W�)��M��s5��hZF���"K
���n�uK}�3�˩,��ɒ́���L*����9�3�*��kA�h����v��m��6�[�"�V�.`�=���?���������ņ%?*ž�:��yׅ#����K�-�|it����3ww�<cR^Տ=KU}�h1�%������09�el+W�v��MM\־���{����=�&��@`�yWc6��M&z�f�q�iÀU��܏����Ϯ�.]��x�@U�z�� 
��e{{8�tvKt��*��놑&����
��T���kh;���cz�9�rs��Lqj�
OS������f̜xo��v;�T4q*��E :�e�HF�Χ2uS�4r&o�(�t������f,܋b���#�NŭE�[�F��;"�䫰�-��S��]|�J�P�%w�Lz9�%���ht�z�Sf�l�סN�q�
����,�X>�Wb����T�G�>���3��hU8�O�T.�=����;Cs����-���{1��hs��DX���>����d/�oKf��3\4�$�bT𳫘����C�^�R��!��L̢lv���NG�:8k~-���T=��O7\�6��d�xQ΢M�:)�B�ٓ/7:�������[�n֐���D^d���_xӇ5�A�*�����G����8�eMPW��Å�)M��[��I�t�1-�/<5wL���>��p�7���5)m�&Q��%/5`��W���b�
�iܝ�fw(7l`������.��
��0_#g'ckP,d�Q��kj4�jo�Vb�nd�^���<��c�l.~h���1c��}mP�W��.�������$"����������VEL�q1��8<$�J��eГ�ie�jS�xy]X>Հ���)q��z��H~�LX���jf�q����s���yӾ���(Ad�g���8�({+�1B�`Q"�$L�Np�+Ky=�/Wr ���x|�.T���x�p��pʥ�t.|���m��uw%�J��F,��6�C�1^y���3�H�p(� E�B�n2�u^^�ָ�M��ڸ��d����*�y������z��ݮ�m0��R�%m2�<�`0u{[:����0&�y!��%{���&���\'v���ͫ\n3}׀���I�H��Ԉ6���o��� �|�f��?��ٛ�a���abZ��o^rz8C�!}��q9�爛9�
�o�_
.�o�b��������Գ3��+Չ�M��v|�q�
K����؜{}J��ONH/h�{�p�=��j�P�F�oaOu��Xm�H�5R�[F��-J���S*�иQ�Q��`!ڐ_����y<ɘy??)"�Mq���j�#F�*'��b��3��<<���qUƭ���f;$��[��h��k���Ҵ���t~�h��@�6/I�)չq�WD���7�q�3�>���Sא����l��O��P��D���&d2@�#��Y�@�������VFn�	�R����ԯ{��ns7,��H����T&;�k��7�*�z��f	��bU
M�t�ݖF̟q�����;4���*�h������͜7���<v*�,G	`�'����s�5I��P�	�3���=�Eso;�yݜI�JǾ�3�ciP�
� Â��	�jbu!?�`=�Sw�P�UjBk·<�zuF�4Bќv�N�9:TZ�� ��Y�b��hɨ|^$VO�u.n��wY�*����;5%o·R�Y���b�6l�u�]ђa�-Y�;��3��y	֩�t0�ww(f����8�ĺ��n)զ���[6�w7�Λ�����aR�$l�
����&<�V����{��=�WJ[���Ô��9�N�:ƍ������ZAc|�xy᫤�=m��N��y$�"���e�i�����s���O_;#6�2�++����z�����̉C�TB�g�l��Rs�BwB��k�{�Vk8Ի�&a�c�m`�\��a�F7,��uҲF��2��QM�U�r���D�*��"{B��-�����`�jz*2�o[���RR�.V@�-��dK{��j��ᶳ��u1h�U �(�����l%6�K�cU=t�ML �;�\��M\�ˮc��4�ǉ��(�S4)i%��,��_Y����6�Cqį������o8Up"��V�AF�i�w�������q�F��`�͙q�6-t&��{�-;t�`�ǀ�Wq�xc��s-��̊v'�pι��GȖ�2��m��:ki7)�a喻x�Y��S���黬侬9l�Ȑ�:���>�;b��{��i�Y�0a����q4$I��=�����ryn�Ǚ���I$�I$�I$�$tU�p����R:�6��^�/>*�fk:k7hЮ.R��b@�C�`L9;�f��F���+�2�
}�d��j,�����=��xx�1�4#���CJ�i�4/�:�h*�d����3%������1	$��#��X��[{S/��QS$U�|���
hЬ9� �Fu}hl�J��j��r�(vBa��T.��Kjn���erh����[�RŌ�hۚ� �(�J�:��4�C7t�M��e��4�V9Hnsc��˥��l��Bt'LV��e*M�R,��y�s"�wD�2�+b�E[(�S��5}�'u82���������]�<SC�9)��އXU�T�z-��.�yu��"剳Fr���vƙl�Z'n_)�\���e�ԓ�J�x�n�x���g=!���;XEl-P��ܽ��/M7puM��e�t����������2��d��{�ưm@*��Qr=�K6�~^����h��ض�Ֆ�o!�Z���ۂ��r������-�"y�r99��H�q�ԊI����eeWt.�.�kEc��r�e���iM���Sn���IZ�`��S32fR���a��;��Leb��T�P�L���2��2���r��4:\LV��V�Wz�Z\��J�MsVU�Q��[ur��4��U��e34�t�i�C��*-��2b.�WH\h�-¸ �
 )#�\is��V�>B
�1��ZbUF�[U�]3l�Z��]�f� ����W5��eMm�kI��5ui������3YL��k[�ė.1���s�k��!�M�Y�f�D���ģ�]�c��Sl,��c������K��m�޵�n��Dѳ�W`�mj�&~�4�P�+�QQ\--��(*ʆ8��Vi�n9�5�E�Y\�0�h��:ʊ[bԢf��*Bڪ(��h��j���ՑTE���liQTщ�(�cF�ն�ailZ�D6���O5Lݡk(��k0AՃjʕK�ȹh�Į� ��E�MZ��4�R���Q��L�ʁZ����e���y����*�����Q�Z��G%|(�Bn�7a���M]X\^$j팷e j�@�b%����`2��ih�
p��I$����4�1���"�諨�#0V��+iƊ��!S ����-���)��
�:s�Ǐz{���{���&��
�^�A��u�)����)��ΗQݯ
u���*q��$�pq{.'�pp�z�A�q�,K�=@���DA�QVX�k_}Yd{y�]sP_��Z/�!���N�nF�NF�ٵ��^5;�e2=($���=����=d�1nz6�16�Ddl%�C��h��͇���ࢼ��{��b�S6�Ŕ�3�V2�u-���J��<L�4Ė�_==���Ti-;ޝ�R����84z�#ιVb�P!Dm�7��Ul_K�Q�]8 c���.m�g^��Cy7������-�w(@�0*��P�Er�U�V�Z�y^b�#t��7}��7���zǏ�
�����j��9��PN��*�DDt/@a�'n���-dC��γ�5�T�U{;a8�&Wr�k�9.&�S���p�qq�P�0c����!�񬏽{�1�v{�o�����ݏ�6�A[��gYu���M��/�����K>n�������a3r>��u�j�-�������|�n0$k�|�Dfֹz���7'Of��j5o� ����j�9�j���X��<Ӽ�s#r�إ�2h�a*:v5$?Ϫ�<�T�K�R|��[Co�C�/����4��T����S��6��$H�>*�H!��wH�@+�<�$��k��w�X��-P5�:0s�Z-������ᆯG��"Y��/x��"����U�V��F��Q�t��:��8ѳ�}�g��[	�q�5�o�J����ƀ?._�N�U+�v�bX|�1��OƗ�x��n�ͨ��� K�r����C�w��`Gʼ(lDp��M`	+���
~�]ԶbE�_fR��3�^^:E��L����nk"���&\���S���un�Z㬹���cz�A��*/r�~���*��<�ٞ�+��&{B"�YlΕv/|0�}���"<+:��a#0���tVxz����xG�UB�y�զ�k�?�m�oL꽨�+Շt�m.���1�z`�Gh*��X�N�9��}����R��w!گUŴ������d��!15r2����MEBHF�t���Ҡ�e�N2Qfg,�͌����zb�f!F֙��n|P������+sj���z��\���\�sw�Ո��L��qfݮFv� d���!�J[�w��grԵ�c��_�R�S�����"�7X���+h�7S�(�^|�	�mn�8��MQ���ٚ�J1�p�Qqj�rl4���;0��OE %�������snӅ|��V�t��O���.z:�dc+*ZwN��>F�#��	�ؚ����kkۛ��Z��,i88z�7�"��C��}u���:�9�l˩�PC^�ճ �t^�^&���j�T2�!.Ŀ�r�X�ϒbåˆJ�:��S)SL�V��Gh��t��4�8�6 �Z�(�~
yxM8<2��7
z&��q}��G~.�������S�w ]�ȡ���Ht*Bvdg�rv�:4硕��H���LI����[:��pc���=��g��;��o��k�g�Ŏ%��-��>&���r�գ�'��$'"#3X"�g7�RiC���)����X Y�R�}r'  ¡��0pа�QĐ� N�I���j�&�`)"M%cZ��-��IvcaZ�E�!?r��7�&`*;n9�*�����]l����gA$h.bp�B�7�ё'�%�P�œ�lU-��f�tc��w�8\��c��o_iV��2����GR�F�jV���$��|_���%�0Y�UhK�ξ������05�+!̷�ǣnn�a�`��͖/���7s=&]ߡ�׍����:�⇼]�chL����On���c	�m��!C��W����,+�.xΙ>�p�)�.J����J��l���H�)ʸt
�r}�!q��� �#k||�f�uΰ�緲<�
u��/�+*�������<��C<�����FU�w��|$�։$GU���? �cy�F��`w��
[q���s�)�Ν<į�\CB�e{��GE��P��"��!b��A��PmҙW�8@eͿ?=�[Y�I�N�|�sF�=�i�x�W�J����z�X�?����T8QP4Uq�G�%K��P����������Oز�ŪS�������]LoD��<| 8�������36�6�[��b�id�F���U_����(���^N�\���\��m��W��.��3W�6����}.�4q����̳Ycdy�&�k ���@����U��j��ǎ�G��`K"Tۛ�y����!�:&����u�ZQ2N��W�7$ye쥜�� ��ys��V�����]��syS��q��6K�H�u!�'L���P�:q4%�C�!L�ic�6�
:�����1O�28�]
�p�yI�C&v�@M����B�8�x�b�r�-wn�j4a��Z�>\�T ж�0����y�]w�םP�WPioa���k�y�"N����.��/]Fa��-�s���,x>3룃���r�u}��Z0�ߩ&�(/�N�t(�{ʊ�`��!j��e��T���S�j[�F�$��<��|�*9p�ǹ�=���<!*��@���{���[
d�������*5M��άm�uD΅���.�]ɋ�&z�"�ڈ���[�!q��������p���N6,a�A����u�BF�/ڻ��kͯeA\ۡu�8��7���
|v�L?�ȵU�Q����LAå�)	�u��:����,<�I~#�5�/z�θ���KPD��qǉ�6��S��~�p�w�Z��U�������,�l�9]lff�b��%q\n�.C��6U]��)�i�j��-��cps��׵�Ʒ����c�T��d9����@��u�H���ĺ9_&w+Sf�5[,s�qN5��*cfKӗ�V{7�d]��kD���\Y�U�E�oFlL�0�녻�.��w���c�����N6�N��H�(P��G T�Bv6��ʋ�Nn�3���'ݨ��A��K8���./c%՚ԡ��ٴ���@���Q���R�����S{,k�
��0�*9�;�t��0<=Ch]X ��y�B������#�;�W��u�]u@��	W\�烒�`��8�z�-GMwK'v5#Ƈ !cM�â� ��Z7����bD��*�Hq1Cb�&������Z�'���p{GI<pp��@k�d8h�x4C�`�{؀ZxQ-Z���*4u5y{GէE�����K	�ꞣ���h�xd"�Ut|�C��&6[s��t�	k�p��xx@.^��DrGL��U	�*m�;���w�3��s�V
::�{�į{��F
�*�Ët������{k:��"�K�odm�p��SQ��l�p0+�����'p���+k���GXxq5�ViTf�aw�����Rg���S΂�`�4���xǛ���O>��b�\,��q+Y'2���&I�+h��pV�s����b�Ԑ���ْ(|w}[v�9�D��g r���(�Q�z�/�x����M&�Ų8y�S�()��ɘA����`y|�9p/��WR�< �|=��ޮ~O���.��#�E*c�tv�da������%{��S���	g�űp���k���rz;v+ό�y�;��~�'��h�Uᨠ�P�OϨ`�褐�o�<t{��U�zze���Z��rE��g/ޔ���a�O�ϩ4^
�\ֽݵJ���n$",�S6:\[t�®�ɓ�)J�Aه;!�bw�&)L��Y�M��V������ :�ζ{ь����=7�nދ�9����I�7yut�U7A�(6;ԗ�����!�l>�
b�b ���l��7ƣ��r�:���q�������7BQգ�¹�J����]$Ń�Fv	�&������-ҶI���
�_�T��"����(��yx9��[������7�h��O�ҽP�Y7Y�쮴~��D��;�ioZr�����r ��ʽ�d�|� pjԎ�fN�v{y��0,�r�bE��ڙ"&ul:Nf�ֈ����ƚ��p�YՑ�d���nG��t�'�'yL��Jj
���S;)R��B�3��0_#ggFGji{��i[��J�ʛ0
���Kh��'Kr�U��Nr��ms�)�D��sy�|�[2j�f�DC�NsJw&*Ey��P���r�|�������D���')`s����z���bĘ�.���b�Y��p��X�S'ژ �*y9�N��
jaqz#m,�yw�c"��V���)��?)�V�c�`��q�D}�����z�r@�yg��!u��ԳK"������7��R?[�L��Lm���&/ɥ#���v���{������-P��i�8�.\
g;ifdA�N�w2�έ7f3	�#6�9Up�Pq�^���\V�v�����r�i
j0�i�T�N�!�����j�����qu��8q��H���ĳq�8�y��uƂ����0�Ut8�V��`��w½� �S���<Ư>����3�3�x�|0_ڎ$�cƗ�۾eK�t�8J/B����O&�D.��Hm�ُ��"cJ�HU�JMė�4f�&��+0Ӈ-	�����+���=6Q�w�uDxY��\�7�����>��ʳ��J�obJH�|=ۅ�M�[p�B��+2eMG	���B�ʙP*o��W/��/�7��w}X�|��td�]��W5��92�#F�"r�-����L\ �sɬ����BKDuw-��ô�;��9�N���(Q&xNi����qgd��ù���=��
�&�ֳö�Gz1��� ڕ`UЀ�mv*;H�~>;��5m��\�8tw֣���*�tґ�4���L�P�\I�5��q�f�����8gT�gڠI��*#!C�="Aq�<���V*d��@n������A�Un�*s��ۨ�Z*���KA|Ht Ѵ-U��:	�:���V�I��z��}I>�t=WX��Y�]M�u��౵K�]����]=�P�L=c�@&;��6�5R��U�
@�����>�OM?�p��J��v|x��bR��*���E�a�%\7�BZ@���Cx�Y/�@���W��S����~;ا�yޖ������uau�K�����4d3
�&�k>W&��ڂ�t�GV#�Հ��/*������'�մ��EV�|�C�>�����3�:���c$�C����qu\\bt#������E�Aa�t��K? �̞iF=�Hg��6�JqnX26{���;S��1ڈ��R f#�C�������=�l�ؼ,�!ܐ��[� �p�������ޱ�I�u��<��ٌiH��h3��ؾ�vj�-�|Vx�q	��~>5���QX,���vos�>����Z��T�|l�c>�t�16���r�����c��\wjRy��1�wp[.�%=!)u%�F�Ѧ>h]#~3��ʚ�O��#�t7��^���W0ա��M����A�y�35h,��F��]B���V7������0�^L�j�˂5V9�*ژ�OC�ا�'�H�b1"/�]A��⟒ս| ��z���m7[�r�ʯg���Sy�&}�Y[>�~a�kkx^�S�/t��XYʽ["�U�揅!\�`>1	Ѽoᓕ?��J��il�u6����>�.��wm�pJO��僄^Z%
�1�F�������7����ո��*���\��:�Ik�]�ᴠ�Vb�K��&Z �|��''V��9]��v��}��s+�l�-�K,�k_`�rj����˾�B��\
�VP�#)n�Bw�e�Z���aյ�����Kl^����s�M�o$N�rɷ[G��ө��l]E��yC���΀ꊭ�b��4;�����wU(�l�့<�.�WL((��*�	���noQ���,s���x�b�ymڛ{J�3�"=0�jt7rti�]�u��@D���0�Q'����W�};c�A��9���Nb���ftc#SL)��Ʈ�f����ۓ�,"~�}1���(حQ.��b��%o;�2�Uv�Z�)�P��~ҲT$���E��7�<�����6�cÇZ��e:�����I�+�#.��V�e 蜥��ξ�2S�\��F]�������r�2�J���K��;"Wk�ɏ��(eD�Y��t�s���!��HN��LΝݞ;v�Qv�����=�����fŅШ�j��&�\�*J��O�ck���x7e	a�+(0zg\ܭ�n�G:��J3���Yc�z���R�+�K�]���h��a]�(U���9�y�&��L�K�� �$i�mG����oCx%5��欹RB뮸a�Z�Y��a�����U��1O�d�޺���g.ug5�;��_rh�ܒI$�I$�I'9m d:��Sab����Uҋd���n�8��a�.�ce�wE�嗉T.�dQ�9����Z^�+���A��0��f�\t�� T��Y�+�c�R�,N�w�Jq)�Y��y8a�x�eK8�m��#�7H��<�4�7l����n�/����`�]�OV�c:�Ba��Iu���tK��<�׽�W*���'wň�yW�ʾ��C&�Hq�=�pv������ݬr�+�e����\0PV��q3C��S��`���;�q4:Y�7[\���s38���X�ҋ|��j
"Ù�F��K|�����6����]%�,X��ĒLq
O��{p4��ͱF���VZp��-�E�����o{����Y��FSvQ)�6�����^�B��'�^^[U��2��������3Jt�O2�>�4�c�Fd�P)�-�٣t-e��{ʁ��#I;;z&���e��bj6�W١I�n��\��+u���ܨ�e�����o��IK1�,��/�����㵃�!�}�G�=��nu��Ȕǡ�|�s��A���KD��If�ݜ�JڎL9��oۓ����M!����i��7�r8㌶ԉ�NlI���V�$nD�r9>��V~quaZ��ʿ:b��EY�n&9[�D�V��qX��w���1�3UF�,FE��La�WYr٦.�Z�Aq���,�Tr�WwF����ZcK��څ��b��aq2���ˉ�L�*��k*[i�a\ݘ:�ʹ�2��f����"[�e2��U��X��2f\eAW-�]�ۆ	�T�oVf��k�1Ff\*
T��X�!��2˔mZܻ�5n�5�T�̯���.,�bar˻R�d���n���ycu�v������-�1
3�L3ޮ-�QQZ�iQ�YJ�(fU[]��4��.�+�/���;1����Xk�&��ͳ��ITvܵЖ���,`�,P�Yq��j�+Wz�����cQE�q�CM2�)3(UE�㉴����8����ch9L�х����wn�����(�LB��FҦ��d�*��a0b���f2�0�-h�X�U���լ�cs1�����C/rf��I+��лu�3[i5w��wp]U�9���Ÿ�`��)=���.�ޫ֞�x���򞃢o�#0Ɓ��I�J�ZO���L<3�A�:)W�6�F��j��^c�=�/�>�������Ru�+U��&���R���9ڻUK���d�U�"��s�t����v=���w�K���-�͒���+-��C6�l�߽��6j"��r����'92�M�`|f&,eC&�7v𴘭w�p:ձ�Uq�v�m2�n��ȸwW��l{�ܷSV2���ݓ���[}v�m����H�B�>iX�u����V�C�4z�q�N���7����=�t#t�t���C�_1q�Sb��-�-�Eg��l��\G:�n�q�9~B�*�/ZTny�y=VD��Bbj�N�*j(B2��Àz���,���a��7ҡ�P�q9#SGaT�3<���(Jx삹�����T���1�W��}|zd�R�x<ʇ2���̪�s�z1���Ev^��6�^'�ǹJ6�L^y�#"������"�	M�z�O-t�h�4�룠-ǋil[�_aљ�I�V������IM�-SB�Q��֧(xu�޾u���V^� ����)$�]0lW��^�d�
֜��/�s+�����{;+0~��]JEp���Z�/�Ό�]�k���Ϊ�"#�]N�1HU��X^�_������\C�[���Yl����n�J�>ZS��Փ�sY�Z�h���m������e^�~K�䘂��Y�^{=�zz����*2	T�З�<~��2d_���͉�qaˍ������1�,��J2S}&���.tBRcb�gb��TK�0*��J���`�w���z�o+�Ďxr�N�a�G�@l��'r�"Y���U*`�����;WY-��~��V�+�U" ���sJw�1R(7B#y�a7t'��x�CF�'~�o{�=�7F]+�!%Z�Bws>�����~���eGvc �>/��)��_���Q3��X>��iS��?��n�;Y��b˚*��75�/�{��m�N����r�J{�W�b!���m#���:��x��\���vx�2� �����V�tkږ�y��ѶwU�}���';_ѽ��+G���8�UǌL���z`�ܖU����(�׺������۱(��nq��{wf!\�V�c;u�x� �6.T����~�IB�S�{s�tZ��j�����26-�;�p&�m�DdPY����K�#X4b�[�Y*,@���ͧ
l#�ʠ�!뫀�*⹣��uA��F[Ŭ8���e��D���L�4��[t\1 �q>�;+�C��W�:�������gټ��)��L��j�O|����hq��[(����>�Un���ߦ����4��hOJv�^����*We��1�+�x:�\��zb���˗\��5uw����nv����#��
ӔN��ƴR4z�'!��.�l�)҆ͻ�<I���Ԛ��Ԡ�`l�D,3|��<��J]5�'ڼB3�F���9��֋��Po�,�����͈��/�����*�+���s�n����\<��Pຈz�p��w{����)WU��d��A�ϕ��A�0�ޙ�i��.$f�=s'#6����뽰�F�*#´b#ƕ3[�E�d|�	�xU׼���BQF�{9�(m�3����W��,%#/
 ������˲%�Ud�s�yn1Ow^b%��3�[�����6��,��&�ض��1���.�ml�*ܰ{7j�7V��CEwB�d$� �ۋ/��5gv��sybRG��>���?�I�W���C��߇P��pG����;U�%���1m���ú|� n@�ӱ��F���X����I�T�H�	qb����Ih�xю��|c�}�Ty'�&JHs��LYR���3�
��,���W��qW��,��t{~�7��Լ������S���&�J׀F��s<�C��<�Ś�=b��"o����G��N|v��ɑ��� ���A6��/��b_y��b/ڈ���ʵa�w=}����u�P�LWF�:��`�,Fm �PN,P.BU]fȅE��ﻞ�O2�E0$d^�b�y[�[��n����qFN�S6��5r�=��zx�"q�jr�]�',�eZ;��1�e#�x�tf���öׇ���e�h���}���?1��D�c�)Ǝu���S�v"A�&8Ez��Z�$iN��|�j�zd�렌t��{ ����j�Rر(0�fWY��]C٫k�+ѻ�������oG���j�8BY˳^>��s,�V��^�5m9`͍Cʼ�'۶/�0�3%�TWXzꡭ4�k-f�+4��3��e�	Tk�)�ݖ��X�%C&�&�b�n�S�(K�XːMWi���)n�OjA���H٦veG)�$c�u�+$��_���|�P�S@�Bj��ˆ����r�B�W	��D�?*��%m��<fr��]��S�2_r�x��\s#<���Q�=Q����ˋ�\)�upc�&��F�φ�T֜biV�m�i��t��1!���7�p�9�s���:�E0�GF\��Y�d���ӈ�'��N�O�6
�D�	hM��lʂz��9��L\&�܉*�W��s���P�{�8�V-c��Е��`�?4��� YC��[.�H�'���v�������E7\+G�o�C��(/��_�p*V�v 37�D���N%u��1�ִ��5=mׄS�C�a�QA�����ax
T}���K��={�G��°<���%������
�VP�S��g�ս����aA����Mޓ�ضwA#;i�8y�c�/����׋��>�c����#�M+V纞eaG[����N�u��D��	���~C�˱��kQ�լdR,g)X��j�p���a@fYs���l�9ض�����AV,7�c u��ܵ*2�;��ϳS�o��Dd���)=�Z�?ԑԽ=�9k������=�x��F�q���"���~��-�95a�v�wy�Yº7*�T
�ƾ�s��VD��B���Ei!Ŋ�M��kyno?.}�py4Ws@P�o �k�2w��r��' d[|vr.���,+@�D�X&|nBzn��-
�u�MD����'ۼ\k�<Tt���M��|��IVf�����GN��Z9ąh.�����~[�p�<=+{B�\��go3�1��_I
d���D�Q�
�,'�����������B�yB���.kpM.mܕ���y�lW#X=� �|�v�P���|2�r�u�8T0�T.� �,劉%b�=��s9EEЛC�C�tFD��vo���&����O�7b�yl�7f��CUE������TK�0y�s,8c�ml���)y�%\c)�>�l����ܸ�UbsqH\N�^�4��@����$�+6Wu0q<�Y�̬@Sc���lڣ��U��W
�V��ڬǊ���v����Q=�GvwR�5�t��9Jr���lv����i�����3#�^��-�@�r�Y����U�oTnH�V��^�Y�h7��0~1c]%���@�[]EM��C�{��:���WDƈ��	n�{},��G,����,W?�1u��1@�|��*X�R�[Br�ն���n�PC�UĴ�rjd��!�|���*p��x��_���.��}ǒi�L�H�׌�&��\CN�d[U�Ui�1$<���6\p���N��-4�aU�.��z$��>���Е�N�����7�dlXiܓ�h�>z�!W^9����9���<����/֩>ͮ�6�CJ���r`p4����"�m���L{�e׬�;���PM�#���j�ϱON�=��1ˍ�)�Y�{��\�p��Z�ys�/���,p��]��1�-�td����8�(@��-�2m���p���O���Tj�V:��-�t��ih��Sˉ銠����R�%w������=���g�=ea�p�x�
F��D�=C�1���S�c�_Q�^�,Ω��Wf�Ϻ�a[]�X:fj�F�*�kEd:�@ ���Zv�h)��ʻ\��.��ղ8����.���RĜ�ۤ���v�OӐpL�����V�oLJ;��6�zzZB��wr�q��P��7�1��xp�}��1{]J��5=wʹ��'<ɳܫn��'Dcj�N7N3�=��u�@k8WA�f��2|ӊ��doXݹָ���M��!�F��֊9^�T9�v��S2;b��46hC�]�m-5�X9���~;g_���>I�{ͮ��w	��
�8���Ԍ�t��Lz�d�FeU���/9�ΎmI{���U��k�\Ɉ6-�7��KN*P�C���5}#���<���l��X�r���L"!;����q-d3µE\�OFe��m�.�mܒϾ=�}H�׋>�I�6���W���Togi��o�{�)nJ�vز�U�zS��c�X���w�$cS��32�oh���*�w�
��}���ǱM��4Oj��8sh���hؤ�j�S�����u����@΍���y}b�e�'��{g�����q&{�4�g��Zn�3K��d��Ok)��@���*VX�o�6��w����`�Fp���)$��-s��oaK�rݒ{�/<wJ�9�C|��*���� L�Z'�qx=��Q{�V���z����$��Y[Tz�l�v2���>~�yE���T���,I9�2�#n��
�|�^�`*g<շ-\@ݔ�6��m2�7�2��C�dh��Yy�o+�oqf��N4��=�4����G�Qp���43��L�rZ�G ��)z�w��p�=J��lo'�fV�/9��.7�<���l��8�򰂑::��,�����[������~�Q��oVc��7�lBι����^L�l\����+{Rk�3��f:��Sl�O$��<������!�/����W�^w:ʨ�45B�SY�ւd`i����=K(��T�G�;��x92R<�nN�Nk�Y������Ǭ+�f����7v���['x^�4J[C���|a�j}[�_�}�:�Eqf�m,%n�q.��hͭ�J��-�4vJݫ�E��2��-8�X���mI�IA�Z�&r'�WSP�.���LN ��E�SN]�o�ֹ�z��s��YQF�8�L�
���89���O!M��f�^�^����sH;HS\&��3��kn��m��-[��m�V�sn7{�S��,#wE�D�������\�m���Y�r9]�E�湢z��}���7�Kv����| �3`��G^Rǋ�q��ަ��}y��.]�!j��v^���>��u���=��yo�����
CO�8�֊��n�7�B����C�����ub&��h:F��u�κ ��r���|���G.�`�6�1���i��8��$l� D�.x��>�z�i�ؠ	����Ȉ>Z��ha�w��a�2�'�WF���I�bŷ5;y<OQ����"�LLDDDDG�L�(�4�9��E�!G6�zAwșa����J�<���k���� $�@R�
��"���£a�1h!��y�.�kmTF�fVtH{���E#L8A�l�N쯮��0��<�I����R(oXiYq�a���$0��B�g�a�%b�=�-�\2Q~	��t�Mxqc� ��x�(�?�@�EDQ�Cz1	+C�����M���/�p{��ğƚc��:��B�^��I��ADQ������r�";<�F���Ѐ����d; l��{I� Y��P��І�7 <v�"cUy�����r�
"�eh�\�;*yR�aP�(%��PC&+�V(M�N�JwzX�7MY�Ҧgx������ ���&�ۍ�t��RC��.)P��@f%r5mW�h+��?���w�0�o�I��!�F݌�%�.��&��O�����.VO�w�4t,�. �yON�e��$E�j���׈xj��:���{�4G[�@C���1��i�c�g�I4];�z�u�6b�h���� `�+��bWm������`X$2��\��@n5�" ��4hF�����Q�č�q�.s�9�>ejX'��H��@��T�&S,X�4	yUG&�ټ�;�ro@Qb�g >�	��`o��=�G��Ѵ���n�v�9��k,|N@P���'�8����C�lJ|wi0
�>�PE������#�&IW����w (�2���1�C�螆[s?���BkM.�hj�V����D���J�AE�q�z�m�<���-~`dC��n���{�h`�6������ˬ�X2�oޑMSƥ��H5������:dî��Qd<���f HTQ��6 �7���`R����;�)� .�p��F���\HB�S�t�����xE��J9�p���)�Q�>�