BZh91AY&SYFxj\׺_�`q���b� ����bH^�      ��
�� _m 
T�P�@�T($$I-�Х((P� U$ �Q  �R�I(E)JJ ��l�2����H�����������@�h%�h+l,�Te�ح�4�4�
���FV[l�!�[$"@�@Y[f�d��m����ݨh�ִ
Т�j��IQAR��Z�[kXQJ�(�ѐ��"�V��)%�AlʩVک*R�Z�1R�TA6n u��R�l 8 �{4�بP(nn���څ*���4�v�e��NttV�5�F�6�n�-�wZ�-L ��7k����{��*�ZڲԪ*���� �m�ݮ�t�Λ�4�[43�� Р:�
F����]
m�wn[���jJ��r�.��.�N]��T�\�gT.�S:��m`6���h��5F�i$%���Pm���� �wx�������Gkm��{���I�=�b��s���Q^�һt�{E[aL��T==�mW^<z�²��/S֖��U��z�(w��Tٕe�YA
$)��( 1�ݍ6�j���A^��]��Z�hv����6ʢכ��A��wt�+�: u7l�h�L���h��Riێ�B�F�7
5���z�{X�mT
��UR&�JY� � ��tUP�Ks-ʫ���+jA:kZWts�4�f�s�U;��
sv\�U����ptn�M�����@WTië�KU�
�t�i�:�{䴣Y4�5l�!c�   ��Kj��V޶����u�kKcmL�e�m��v��j���Q֦��f��]:�f���n��ܻ]�YM����-��^�-��ME2��-�eK8   `��{�k���lڝvu���ճ�3lh���ܫ��UBwgm�����UU��Rd�T:�9��N�(��JQUkT��m01m\  �=V��6��!��Z��J��G:�A��u�Hn�g �0�TPJ�e��%Vܜ�@4{:��i��ԥ+CEK+b6p  ݍ�٪Wc�*��Wus��F��u
�P�t��UUP��TU7�����)@Kj�(+��jZ2ER#f�j[T��D�p  [��E[]�
���㪀 ���%�+mۡU]\qʊ�ι������*�[�EE����     �   j`�*T4�  @ "��bJJ�� h� F�"y1
J��L��	��L�L���R�       ����%Q13P�i���!�%$'�&��S�SG�=F�i�4z�4OD��z�v��e��=��.�X�6LOTN��ޛ���2�c��߾����E U�:��_B��*~�QW�?D��*�g�z��������?�<T��
 ���U_<:@�#�'��Ѕ�'�"�������?���0�c ��?��}���eOl���G�2���>0����S��<e�
x��2��+� �ʞ0�e|eOS��=0��)�"x2'���+��D�<eO�xȞ2��	�xʞ0��	�}7���
q�<`O� <dS�T�~>8�Q�zeG�P<eC�Q��x�>2�#� ��>��A�|dx�x�>2/��� ��>0����ʞ2����eO�A�|a�A�~�S��3	�*xʞ0����
xʞ2���"xȞ2��<aOS��|aO��<a	��D�<`_�T�<d�T�<d&�|dG�T�|aOS���s�ʞ0�� ��>2�����A�|`^���|d�_L!�(��>2����*{`S��0����*xʞ0�� �ʟL��Ȟ2����"x��0���� �ʾ0=�>0�eO��<eO�T��+�"x2�L��
x0�0�)�x�p'�	�x��2��<dO��S�D�|d�A�~0�#�.`OG��|`_W�<d{e|`�����>0����ʞ�<dG��}2���"�Ⱦ2��#�{d<a�Q�}0�����>0/�� ��>0��#���>��@<`�)�
��>0!����*�@�C� +�P<dza|aD|a|a|eP|e|a|eD|e~�OD0��2 >0 >0��0 �0 >0�>0���/��'l��ʈ�W�EP�E���A�|e_��A�x���x�>0��#� ���<aG��}2���(�������<eG��}0/��� ��>1>A�(G�v�h�S���F���c�o+$z.R1%��,zh!ĝf�T,�
��[��L# �,$��{��ؔw�j��&{cp�o k+��H�WSb�� a�L��ֳ�!�4*��P%W!51�3&�.�Dd���3r��XW��;�ܭL�S�Fwu����m�ՠe�y��I��hbn̦L2�o��C)a�T.���a^���� xV��� �Oe��r�@7�pر��!g�e�]h���*�ֶN�-���h�6¿)/*Y�2��wX��-5�*�!�tͭ�6k�hO)z.��yT�����Wo����D�	@�q'_kѪ��p]�+�m��ʵ�/,ń�H��e�۹6n��l�j�S�$lb0�Ƀyr�a�ݶ�	r(�׷���^MLT4���	�x�+_�Q����M�5x.L�2lN����z��uL�4.���j�0�ۈ�ZN��D�Vy�q���� 7���P�x��!��`{���{�Kxw���b�����##ɕhkK�ݷ�̳n���ӛ�bOX�bGz�p�2�JTLٕ�J��9��(:lk�	�kmnkP�+W��.�e7N*�`�Ln���<���5�O�Ɇi˩cf�*��m5���ֽZr:��{�lm8�����B"��Բ�:�v�͂h�V�� kt\y�d��v��k�rL#[�������Y%��n�w4nfh����Y��Z�;�B�+J6黦��ГU̱&���N��Ͱ#���i#X#e䣛����j\#I�:�0p����rs�e�rӨ]�ާXL�~�����Cۣ����M<u	�%�,�(B��1X��Ř����A���Tb�&D�U�d��W��MdG��a���#��t���4B��$�`��N��ЛA�ʗ!28���KqJp�2��5�T"Ӧ���U��B��0AԻׅXӌťװӔkl�4��n���f:��t"8�ӍV��ZM�HD�5�x�-;Z��+
�sw�`�l*�K�ݻ8ޖ���lW/%�ٱr��C3K+]p���wV�bԻ�b\Q��H� {2V��V�;&k�hL+]��1������*�f�Rbl�0T[��7vb�t�CAI����X�T6��xv�C��d�jW�!�X*��37s;��4F���!Q�v�i�v'5	4Aw��r�ұ�������7xDE�%m�į��wZw��5�Ia�ص2�la�6�#T�K�+3l�ɔ�N�ۓn.��]���۔��6��tG,y�XPZ�x��J�0V����-�8N��f��3-G�h
�)ޛ����s�5�-*�s�e`��
#U7B�V7�CFe��UZ�4k���[cU�)� Z&+��Y�t���V�&��A�bXvd0e�zDf���I���#�rD�z70fL JFQ3N6���V3���S��e�����I���ŭa\t&$kL�;�f+��%J���p:K��ز�� ��w�"�؝�A#t��H��33s&�˺"�{��F����.&ɗFaY���r\0�H���:�k7�*�K�V̥�w+n�N*�E���x���)�*[�Xpl/Nc�vyI�ƅ,�Y(��,�&\}���n5j����)Z3���g��9�*�W$Un���wXoY����5���2���c��q˂�n�)��L�bVf���%�:�8��I��Ă�a&D�o��FI��aW�-��U�ѠfX�wn� ^	�Daˢ7]�ga���S	��ԛ���5�ىVSN����4������v�e��G/jn���[�Q�6/$�B'(�n�0Pr1{�^��nJ(�ia�H�ba��5��7��ov�.V1�jk�+n��
E����z&��&�kkM�/:�H6^Ib¥a@Ӥ�{�]6��t` ��yAiƷ*�)���M�i�f4��	هn�˵��9O���1�l�P��J�:�.���mF�I2�%��
�!!H3�S�2Ko�ɭYsj�e-n��0 ��5X١��If��N�q�3Pv�8�)A1F,��tr�z�m��-�*nZW�&+P���pej�r��y�n1(��j���Ӧ�����uo1�lR��Zv�-y�� h���V"XM�1�u�T^�IL�Hn���̠�͋�ƮS�ۉM�0���X�C5+kL��B���z��ɖ��	���۷cp%1��3p�گ�u�����cܱI5�)�!ّ�X1[�}�����u`���l�`"%U-ͬ��\m�I����J��j�R_����9!b�c�dP�����ͬ�3�
b�/p�g[[Z��e	-��En����z��ֺǎ��L��2D��wO^�5t��������R'b9�u[x�DӼݎ-�؎M�t�x���2f���-�ɇNEf�S�	f�U�F�%M�lb������Hb�e�j�髛�JC�Di1��J�n�2��g��\
��;���KD��֎;CNb���n"�*�1k	���2�ݠ�4(%��u���`�]i�mR']��H!v"��sE�5��9a���G[��&?k�z.݄�8����@lݙA?[OsX�l7.�%k&��/Mf��2�����!�!˓C�|o@^4F�2�1�1eύ�={��ͤ�F��[��â�F���"1K+��tz�DS�Cq�с-��(�X�u�50�H\�W�i���ͅ�	�.�����M@�K�s�w��{(���U�U�l2�uiQ"f��Zj�+,Q�^J�Ϫ�-�7��+RYO#4CǑ��hٗ+wFl˶6������W(փpB�2�a�����zHl�Nj,����'�u��+^Kڴ�#��f��©��-
Zͺx�˷I�0�{B�P��2�Zq0�ق��:M�,�cW��r����c&��m0��2����{[Z���	
�suẲJt����j��ɠ5�m�ɘ�M:�u�1WI\���;�ؕm`qe)����mff�����C��{e����q<W��aVf�6�ml�N�31����Ұvl$LM,�FV�b��mJơ�Ř�݋B�jV$���=�<X�
jS���R0oA��iFe݃�Q�]�����m[E��V���#�HEk����Q�U��wt�C�ވɏ(�tD�F��C���/R�ĂH^������[��m)��kze�Ӥ��[�U�bn�;�Zh#�k���p4��m���a�.���CRH�(� ʇp�f�Bn�gRB�;�0��$���m�#ń+��F-
����W���ܡWtaa�#W#ĭ��-���wW�M�U��8k�s6�ƃB&���,��5�L�-҆^y��n�N���z�-���{-lB)�����Ԁ)tԘ��
�I����	4p,��=�b�d��*�m��B��l�E�Wr��¦5��ƕ�i�V��N��h�܌��X��uU�]PsN�1cC�wK���Cv��u���ǔ���&��*K��m�B�ҭ^-LF3��ۓF�u�i��i��Qn�j��$*��Ŋ�V<O�bh�Y�At�K�L��mʴ2��1PN�f�{L^��������kEɹ�n-�m�@�W�k#)l���� eiYN�&-��&H)�"��AE��@�/)���iJjU�E޻�hL��m��R����#9�v�(��5:3��-r��O3v�U�Y����kd�ݲ^��pc7�4+,���.�#cV�yn?=/ �AZ�GUL������X �0��ŭ5
��]g�`��{�ICzE���*�-+ԡA��U�w��E�h)x �
���問t)�v��$KշW���F��w�	�­��Y<t �+X^�6�^�I�:��T�u���57�*B�c���D�*����;J\z]*Gr�rPJ�Z�P���9���ɻ���K+��7w.�.���X;t��z�e�aǺ2��f�+pÚ��yK"T��X�-�0`+i7��d/75W����]��cW�f᭽t��湌-��Ok2J��=�Hḍ���]�s!�3,˰�*��/X6u�i�n�V`�ћ��md:r��F&L�H�/	�o 5�]�h���e\�&hytZ��z(┐ys*n=�`�02tf9%�M��q7�!"�e��쪘da
�H��I�̱VRY���F-RMVֳ(��˕�(45���rRpm�M�%�,4�32V����Y��[U�
���h��\�Vz�ll�4�W��Nk,�'��mǗ+��c���J�U�e�m�����-�[�
vk �X ����)V�ء��$�GgFe�)�OZ7���Ri9n*��k`��Zj�
�;m?����-&1���û��ٕDhaɹ�n���#�����RcX����+wf�%��z��Y״\�-�屔MMrŐuk����reY��d;t\3fk;H1f�Vnf���D�K�t��eO-v�[v�����1�5[�t*WE��Z�h[�T����afM(���4�$m�J$\j<�A�ܓQt��+meK�*z���~�!�%��+7)�YvKM[�1�M�W���0�����m�Td7��b�/q[��X��a�����lQ˺��6�Q�kww�+s]��F����J�a�]އ��L"P�Z΄Nm��ʧ�c�fA܌���ܒk9�	��a3�X�+.�=V��&��N����!��.1�U�7��l㥦�xd��n�;����� ��ev���9����׎hM`��^H�n�Ņ����\ŔUi�i8i�ohnbh�1ߒ��k��k7Uʖt��u�#fi���6��6�6݌�d�d��7��m5�@k [�n���<v�K�6�ׅ
Bd�����X[u{�6���<nE0n�@!<��4*	f�Y�ȕ��?C�n��
F�ӽDy�sn�����ALȤ�l��Di��L��fݗ���LY� wTJ��.�fdc*;i�q��	�hV��g��B�f=��\:�h&��'r��l�ۆ�������E� �l�Yan%6��Ř�A%�f�SX��#;{��ƻ�/
J�^M�Jˢ�]���1�[�Mx�cm��5CM�6ƃ��(���*f\��t;�	�'n��h]`�m�b&m�#O�	��F�j�Y��\�m�'3t�Y��˳y��N�YA�u�M��X7�0�[�{V2ܫe�NY��I^�Dke�j��m� ĥ]Ht��D7�UY��/Z�*t2�����O������2��"��D��s|�aˤƌ�"u�B<�� ����9�-��
���ڲ�a���#a�i���.�mf��wz�kZ�t�=�%���H^�1휛{{E,ЫM��M���D35m��6��	q[���Em��
mnPu����V��Ɓg.��D�a�Y4LJ�R�0�mK��*h�
�@J��w���4I(GZ^i�vo2^MǤ7�Ǘ,f��yZ.`ɹ{�hVu�0�Gm�hHާW��Y��6��aǧt�bh��ٗM�
�cĪ]����`��LnY���ѱ��[���Y�T���K�3H�Z7����,��A*�͉GA�j=g
�WH`��1�عy$�b�,*Zaڣl���i�E�GAYZ���Y��V�$��ܔ������ܩ�+����1��1RYQkJn��)o�7emY�n��u���c�t�C&�+�͢��M���5j�ӯѵ�X�eS��*��nj��H'�lLȭ��\{�x����Z�����l�(VT:�H��̙��⦒+u�����m��&�۫�P9HJ��Jm�^�d/h�37�[8�ܳt���;���#�1卆;��\{�sU�&�W"�6���E-��/&��n��M��ܽ�{�]e��p�G/A�[[��mK #s(���B���7V�4i��W�Ȃ&sO`���
#o6�ƳV`kr�-�!yyy�����V��T�Nˋ@��T��-u�]�ɢ,�.��(j�ݳ�xJ���Xŭ���R�<j,�1�{E����u�R���;ї �^��B9�1L��V����+�A�Ɗ���j�7��)nY$���T�ҫv��b [�&+z�n�T��!ŁT�{��ҀǪZ���j/r*�j�׵*+��Ԩɬ#�{�٩Q7rD��^Q�&P���{�K�	밲ʰ0Ɉ�������s*+�bű<�z|��M	[{��U�)^]>O60��&	�i�p���g/,�3L�^K��P�'S"�;��C���j�{O5b�2F�v�+#�Z[@:O�-�������,`n��͑���&k�2�T�nJ�ܶF�z�P�@yR�k%�Ʋ��y���{�*옝� �j��s �o(T�l��h�i�cK1�n\�&���U�g:�,�3K	�PQ-��=��g0ȑ(�h�Eil�Fe,�V�i�d�;�޶���N�ϖ;<#p�4]�p+�(�ک�h&y�x+8�J]��ˎ/7��:F�)%�H����H�e��q���	��P�%�Ŷt#�)9ÜFG&�KJ�� &�T"N�줩)
�]T	��+����,%N1?M��3�T ��a��I�+5��&*�)���Ep�x�� �v�֜��aH�!�4,4��Z�G�Cpy1F�E1����x���AAK9�#C,�5�d��|�Ш vwEa*�KA�xr� tH�2K����Y6�2*�dP3�
�D�aV�,���*�I�Z]��SK���Ȳ*9F�'6���*�쎤�"ID`�mE�xL�Yh�.��4b�K,��bte	�Ùk"�TU�ꖬ��ǲ�����bX�5��_�
C&�Ēt���+�������a֗7�� ���a��~����]�5J�O��?�a��F����5�u9-��<��i�X�xʋ5���Z�Zn�ky��A���+�a�ZH<=wv��B���I�T��({p��v�Ipy:Ŗ՗̼�H(��o]*�:�V{nܓW�YE9eL��y��g������l��l=��0sQmt:���ě��R�P}���J��P�w�yf�'wtwVx'^n)�� �
+�3���e��Η����ΔOc�f�9�U�c��epڼ��&u����pO�v��R��0mr��C÷7D�V�V&���]���l�&N2�٩ڻ�˭��cv����qrW��$�:f�.���(W���춹�ܒ���HZ�$�Yv�[a���f�scK�蓦�Fb
/MF��&�x��2�.�⩊�p9[g�>z������ܽu6�ݷ�o��-g$d��:m:��x���d<�D��f���ƹ-�m�����������0��O��̚հ+\�T�~q�CX�k��f6�%.{:�<��5r�`�1}/Z�5��\X;��e^��չ;�n;D�h#�������)]cj�^�%c��9�q�E��}�0�u)���.z0%�R�+�����[}&������4���w]�xp������W5MK�^^dch'�B�s .:�">����)I���3r���v$�(���n4�W"ɥ ,+��-��i^�걃��;�;W kG��8���Z]r���C�{���q��@���X2�e�[�wR�ƥh�\�� �@��*�air�{8�'f�X멞��'�V���b�:���f�e�5{2������)ve�M[z�fir^*�
c�l˳���bN<�9s��ݪ�H��t�Ɇc�/bre�K_�F�#i��rk�T-C7�V�K���{gEҞ"/���듥Ygc8��d����IȐP&QK%�f��P�:V����k�t�d-{+�K8�A��3qq1���wa��d�����S׮�X�G(��pZM�0�Pݮ�9�r<��D�ҥݼ\����SE��Mr���sW���ξ�S��N�^gD+���Y3`�y�:4��h������S1e�����Ł2s6�:QQ�E���h�����YH����dŶK0�)�}�7����wa&8`��8(���&:��2�B$��br��D:[��4�Ys_)a���6���Xʹ��ý��,��}�U<�g')� ǹ��Q�XmJ��.��\��v��#�|�+#)�<q>m��D��{��[Q��sQ�V��h��^a
<B]��:8Mf�nv֔3X��mD����n������Y4�زl�{��ۦn�2���4��z[Xt��2D`Ԭݲ7�\�k��sS�[�2�(��^���'{3����
���u��7X�Kzf���;���'��/I�D��j��[h�O�̓C��Na��Y�3ΚEx�.jy>��:f�׽.�!ʩ�\�c)�o�a���]��i��Y1��(�NSH����tKH.Vc�CGc3(	@�a����>c�mpL�ଡ଼qG
���������������U�˔�6�A��}�A�tqr�j�GX�������C�#<�w�S�y��]�
�ѭ{Xul�b��iՂ����{%�S�Ī��3��<p���Z47�����@�I�S1m�b9c*7:ƽ�9KXC�7^���jQK}���4l�ɶv��S���T#��f�����܏��BZp�:8Ys-.F*ɖ4<�����q��{V�D`rӷ�n����$�K�+3�S8��y�z��;ŷݚ6�cw5�P�t��!}�7��=$7|�Vk
o4���[Q��
ؓ�[�f��NRYJ	#�9c)�,õ,rn5���R̊�#D��g�\��q��佻HtXi�W�F��G���\KFB��Ð��˼�N���̀�],��Zy��\.���2WV�|ଓ�j�x��㫰�5ʣ[��j�K#ON��z���ڲ���eu�7:#��\H���B���:}8���3t �b�����lֶ�|����G���D��5��n�;-&o7'ZF�ncq���i��7i�i���j��6h�!8W���=A�[M�0H�(�Nu�{��7��=�n���nuKfE�36�U��:�Y��κ؞P����_&���l��d���!�����������O n���x�/N�n&�)����á��E��:��q��F��.�v�x����J�v��9)����,r���Lp.��t���Fv��>}w�W�[�КZQ�����ٲ,u�3�Wfۅ�&�M���p^�6�MM^T�UCV�=����lK9n��b^.�38�-�BU4�c:q�z4t����;��0>���ьւy�}t*�K2^;���)��Va�E�O-�+�G�%oB�*����2���_p������<CjJQ���2hWW�j=��KB����ő�ca�+�E�՛lYْff��v��ou,Q0���r�Z��:(*�´v�Dd�l3�9y�QL|�^\��i��å�����\����S�0�]���P�b�W�w�.���"k;2�:�ܮ�u�r�pv��3��-��+~��+Qk�w�3}rJƈ���Y
{J��ؾ[�ka��n���B�S8a<��\j�_*��'��h�9�*�3vwdo=��mv�{ݽb���a4��L�N<���d�Z��5v�u�A�1`���@��0�]�̼`�ӗ��P�h��nv;�Ѯ��;�U"	�[��v��4�&#vGnǄ�U�L�.	���ʍ@Ud���i���{wt�NU��'Q��L-tKoL�0	{�����5�鲭r6��y�D�t�3-ANF��t��N�,xK{�Bu�3��D�쎖�\�9A�W}�iXVlyD�-圖/EvQ��jQ[ �+7q�J'�����7U��t���#�*И�������t�@���_3y�1t���>Շ��Dh�T����-�H��PT����[�[��� ��离�7TI�W�9��l�]��i�x0载,[vH�i�r�Eby�kL�9c��iӗ��3}.��Wc#���5B����"�˕���B�.eY}r�
ظ�]��\{���S=��u��P`�/����q&� �[r���QI@�S9�yݤi���@�UInp��k����ac��,�ɛ+�Z���ő��)Mnkt]Aon�B����Z݌���� g��R��ך�{|��p٦S������}�˯nHn�wk�Vа!�]$�ܰ��-VV��nn�:�GR�s[ⴗ�c��X�iF���uL��͗ ��kZvj;�2*�y���%ͦ��z��!4*n���s�k�&��]������QHq���޻�i����g '��	[�r�e��!kT�$��'�|�ܻW�1^��k!�I�iq̭�"#n-3w�J�\p���3m��u����.�3A��G�)���g�3��.���9q�+��{�r�s�]M���C+n��ʩ�z޾�_*��	lXD;֑�I�]��+4L|��D�u���˕�3&�Uv�&�:�#��!9�+�T�M�o��B�v��q��B��v��j	0�q��T��yY��5>�ye%���p&�38лap�͛�9�
_IZ�˲��(#OeM�h��4�����w���&ˋ!!���3�V���Ϣ��$�T�A�[oj�9�öh]���ʕ۬�
Ŗ֪��I�^N�jiY���3)>�XDbi�w��o�tɹ����a�VGC��:�*-�������NY�5�pҷ�k�ˬ;�`�S�^a�iA����K�P���i[�hQC�R��2�!�իU����(�m��Z�<��!<���-X�/s���fv�:ۭi� �J1��#��S<�+i�]u�O�̱���ŗ���e�Av#m�ʾ�R� �c��k5d2(,q�iV�ԩ��O����m!K�u�v5�
�1�W�j�*�t&��Nv5'a�D�,�|�%`�o.ۥ����cW�q[ �=�\��
9ga��>�t4Pb�ő�
^; �w�R�J�vt�Ȫ�"�#��|z��L,l�q�/r�$*竚1�,���I���ӷ-W^�6F��Ш�r��x�T@�b�=ԁȲ��bU���1eg���MHI	�ۥjq$�@"�	��V	QX�s4��3`��پ��ӽ�U�jTul���7��"+�T��A�.��wJ��C����Nd:&��.d�싲!׷;]�a��C5(����9�6�F!���[����M<d_Vv���9�.�9#EA�Zi�� �a��]0���3j`�v�z�3���4g���&��k�א�@�<x�M:�f�[ߜ���tFJ0���eO�3m�|N��ޒ2���b�A�5]a��h-U���m�Y ھ멮Sf��%H7�k��U�F=	>�E�U��y��H�\��+7T�oZȤ�Td���F�ޥn�4sql��#�'>uR�>)�1�_ ��.��.���qK����ն�����a�N�a���g�u+��y{u�����o�:��-b�F��(Q��M��Ҋ�`+�j���˼�:���#���M��v4,�S�H7e�j���we���U+��!4��h��vT��;��T�Rٽ�Y�Q�TQ����L�X�T�Dʟ\�4�z����{1�,�\��J�gc:x1:Ж䰨P����:W^�h�-�t��x��g>�^Z����lj��H@x0�Rݾ7�Y|�UԬ=��[�PK��>��ʎb̨��Y�H�㴃��M����Uɍ�o�J��e�}�g*=�ypgJ9�bUr�t�C�g�;�a��8��ZDlLӭQ;׌fyJ=�ʹه]�N��:�ڕ�YjÃe�m��'�Q�t�6���|�18��t�6v�_E�3)�d�� +R�w�D�[�	��k*����rK9�U�1wn#g��7�!�&^N�����ݝ��7�OB�S��e+�/�[�d� �ު��wc��e�f�S��I)�wi��8�xȻ��5:���+8�N!�U��Fm↏g��t�'� ����-^����)����e�,�����Vc�2���L���ە�6J�j�^F���5���j1�ar�f1���;o���a��.F�v�I�HT���\�=�}���X
�`x�{%WfU��.�D�[���ɠD�0ؼфd�+`;���JAV�Js���	|��fkcr�X@V����Pa����ưV!L�(��|<��]D��pw8�n\8w9�_`b]����饫lTT�Ҋz�dX��Y}�)N�[/O^(�rƑQWk;X��gN��K�4j����U�3��{��kv��	�c���U׎M�x ����6#��"3H�o*4��׽ K�����p�wU�N��@��5k���%��21U�%�#���W��H]6-<�ӏ��o%�!�7�{gl�5]C�l�G܆T��bL\��/n�>6��Z��X�GnN�ж���֣L�ӦG�-1ۘ��+\�}7�VF<�Dr8 $��j�1т��Ҹ�d�V��F�2����0�L��?�*Qp��ރ��^��d��<Zz�.�tr:=��ڦ.�je�mt����$F���l�M@��"���W�����異v�K6�MISTǆ`���XiKljͲ&�nP��ˤ9 ��%v�ºÐX�se�O; W��3zf�|r_�����t���,<�5´�.�깪?=b��eV�v6סtV����-�ݕ�Em:mWV�*n����+�dI'��[NV���{Ϥ�8���������nMˮ���Nx��npUyPF����5:6�U��\��Nq'en��V�S9.H�@�|��'#�ۥ��[kq�Qh���]Q��%�[�'V��;1[i��ꕣ*���eBe���dl�e�7;k$߸G[�ݔ�=;��r�%�nlv͜yp���uX��qb��
�U
�l/*oq��z�҇]�:�٢���$�|���mio���a�x҆ӏs��3yw͐�\���h��b�ڭ/w�TDGQhd����2�):���:�������u5e��#�
�[/��@�L�/�ф��؏�RYsL=l�o���9{�`�)��Lm �-����2�.]Ai���:�����p�@��hҧXGv���9O��ϸx+��n���#��ϊ��v�����;j��h�mRq��'��3�̛:�N//A:��[�慭����󂼛�����Z��z����*�]\���63v�ە��8�[��C)͖�4�I�F���f]�u�c/��m��i�F��������g4�ͼ�ImY�
�mґ4v���e�\� �4����q�;�"R.�ݝҢY�t��/061��:���m���ʚy�0gi��3a��p��
I»"�i-�U� {M���փ�Iv��M��m�ڃI%�n��۰6֔�2�X�[�23gd҂��4��j�-����w����u3"�f�%߫����Z�N|����}G���G�� ����4>�>C�>^�=���' ���t?$�S�}�4���Y��O�;�C�>�<����R��כּ��\N�I���G��}���h�y<�6CH�S缜��/W~�P�JN�����ri;��׼Gw�Yz
��?��o��
 }��������'��#������ ��H����������������O�{�׿��wgt&+�:�˥��]輦L%ava��)s&�����]�H�-�f�
�"1Q����[�����N�əK �X�\	a�������T�
a���%�2�
\��)�k':�]�p��i�6��At���}Z��O�|�W{M����G�K��3{e^V6�7lAb��+0�ɂ��:�O���
��K,V�;P���Bt�:;�F9G���<�/(_**؈�-���i�Ɩ�\�}YR� ���Huv<=�_
�e�3��w�7�o3���� �Χ��f[R��W��8�W2$����ѹ�l]��i��SŮ4H\`�}���2�Y˯ovN��Z��)��0]|��12I�9��Y@��@�;F&�e�.���>�/7�c��t���th�R�y�+p؎����<v˩͛��[{Dl ]��:�����Q�� �J���)�u�h�,��Tp�A���T�s�v�Xx+�C��+2�	u�2�Lc�Ǻ�"���V�s��#�n��t�=D�y\N`��V���R��A��,Q��R~ůQAn�u7��t���$�s�7�]i�7;Ac�� KJn�����ogt"mIy'X�pVh��B�Ȫ���0��gn$gL|�^���άź�,�F%��=�t��dk�:�E�8�ո^���4�c���n!+fsm�S;0^oP��ېf�(b��$	��#{_^��|uil�ͧ�m�wJ�4艁߷-`����d���':a���7�2�0]��T�D��F�,��Z�e�����7+�"�����K+���DFA��R<[,>)�w^2�Y\�Ճ���-:q����v7Q��-^�\͌z�ʽ횂;�f,���1,pe��-"�ë2������s꾗qB�Cc�|������i{j�WjS��6]\�Reeţ)�4�43IN�՝"�2����ǧ쉬l��D
̔�A���7��Tt��i��	⼙�ry�n��*��|�y�L���:��'X��\2�R���y�t��uaU] sѐh��k)k��ŗ[��}���e�2��$����8A5�(Y�B*��<�I��;��@n�`S�0p�][&-84���/0ot�b���,�
������nl���oe��.n��J<�OF�o�m��4��$��ns�+�]�ĕ�\�Mf�+5Y(��[�2h�cZ�wt:�owT���j��pL�Z�N��v���gd,i+��}(�j��&�P�d��wѡ��x����#Z��U���ږ���̰�t���I�i��عip}��m]q��Lܒ.Cd7k$�؎�;�j:2���2��T�"3��`��^ˮ��5S@2R�%���o]�zvFw�I�l��3�TǵѤ��-�O7f��JJ�b��i��;�H���̈]�ǌ�|��Ķ��[s�7N�
����%#2ېY�n���pʾ�NT��`��L;�D�o��{knk�J�oJ�Q�;�0m�)whD�h�C��Q���/j�I̱ç�T�
��9or\�x���N�L&X҉�}ÇS/���wE�����ٗy�O�hTO4��^[�9�ռ��Q+�m�Cy,�/�%��N�1E��u���M��â���h4�>p����ނ:ڪ��o�E���l��j�09�b�e��Ov�c�<�s����G�A=�Q�ۤv��|N=�w����"��#�^,���ri
��i��׭k{�%C�F�Ͷ����Y���ܒL�%��֭[�¹�R����� �u�Vm�G�8Vi`�x(a����$2ՓDon�Q��S��B�Y5[�[yTL3$Z���p�;���SU��n�N��u�7���dc�$D�b�5�n�M'��[�e�
J����%���(���/Dعy����\�N���+�nc����j[�9^t��V����p;���9>+���jAG�6�/�v�
�p@��޼�>q����f��䡎�.a���T��[����[�V��d���ݍ�V�E�6p��'��G�f��bap�{3Vn��p[�n��ǵ����;�oU��V�v��؞�Dn�� Ykr᭜�1ji�Ў5�|@P�������r:/�^�����F;6�ɼ:����o�mw.� A�<�8d˼�Q�z�s�w��D�:Q� H��f��bnSym���a�C2a��˷�.��\ �2�K��������R�Fvd�9+�F�4E`�X���s�����U��+q[%���n�A�P�n�{0�o6��R�:2��ӻ��Wa�ܤ5��gc�ot`I��R�fU��1t�Y�.L#%�kk#�++f�yƃt>�J��A�>��`��4ޱ��Y�)\�ι*n�\"�I�-=9���Vf�2iB2�^�z�Q�D^��C'#����C�3�
S:3l�3��ЗVT(�{�eԐ�K���KIn\��neu��Z��u���-f��'�7:G���bLbr�C��K�E%� ��3�^�����K}��dH-�,mtj�9�Iۜ�o)�1Q+R,K'e�noA�)���j��T���[�k�T�`���y�#�����k7�n9q�E��"&]�W;Sn��
�fc�Sdy�h���ut6�ث����y�+�pxo1�n��OI�;�:�k��k_$e����D�������{\VYj[-V��t�(��Sٴ% �n!�&�9a$��*!�Ŭ��4;���H�uó^�̵dW@7ɛ�0i�\�*��X�A�0�r�ӭ��
v�e�X~�ְR�)f�qS&=���^,��}'e]`�H���ېog8 �6���K��r&$��T�ڊ��x��Mn�d�?fn�8���z�:��OM�y[�.�K-&��Z��^]g��
4��i�ZS��b���].�9��ÄJ䩵�_Y8���d������^=�C{D�j� Z<6��R\�䛰2��x��\[+7r������(jn�r)󼔎��<�;W�Pg���V��X�mR*���f+	�^�+���M��!�8�m;�մ⫗n�;[�ݫ�%;�[;U@�2�o�a��� �S-�Op��nA�{�f��WC�c��5\yQ:�PƷWm�'W�L���dY�F�f�8�r\�NU�6����I�yk.��*^�l���4o0TQ�W��u��΀-�b
1-���}�V�Hg4l��^��+j����n;�tD��9f�R������Y�疖i2��#�%w	B(�Cs���l�a�Ш.�N"L�oW�լz$�z���˗L��M�����lodڊ�Y�gX�zR�kv�$�֌�vc�oro��倸�U�{&�M�z�4�_g+��к�pp^d�Kۭ�.�;��[�S!�Y��)JE��?LU9�*j0NJ�=y�Ǥ����.��̌L��r���`{{yv���'f��u1�p�JS��:v�)(�GR��D�2\�m��TZ��-��5�q��.��O��ܯ(,	o�̚XA��V
Y�T��`�v�W��icͤ����4�epl��{j�ؒ���Ƅ@u�d=PV6��妧F�,;Y٠�dm��Gj�f>�6'~ h�{��,9n4�rR�b�ޑ�L��֊��(����9�z���5�=j/]�6�	1dt2!VQF`-��νN阬V7+\}�9�`��V���u�:���L]h�r��J֯sn�NL�RYb���%��}���mf��u���� ��=ր�Y��3G���5�������c�/:���v�rU��򔼙�|���7�y(r��`IW/oh�T0	�Y�	�*Y�])p@�����Ma.*uAa*10�ٜ�`�L���MǸС1_a(ج�c
�Ӳ˚�Q�z����7�t3oxg1P�\�w�&�i����]Ԉxэfu����f��/2�����l��i~[�<���Jw��7y��|8E7�F��B�+f�"�i!R+�Ԧ��H^���Õ$U��8�ϪE��)���[�~@��ͥU�>}��� ��k�]�S�ue��k�fV�r��w�]�tӹ� Sy��}v�[���톣U9[4��ws2�F(X*�Y��S`uMg*0�m����,�inO��D0�0XU*�v��NZ$q���@v�K1��n:^�����u�vOJ��z�w^��6�h���C�!���i�,��6cJH4��X�r�U�C#Cjep�Q��*���ӫ��9�x�VD��}Pƞ�͙m��iP!m�o����Zq���Q1dF�u��aÒc܇����z���Qm�Yٹ�O�Ha��;�w����G��}��bƈu-o`��fAk�fUh��Ә�w&��#sn������+�gNۂWP��cmr�6&ή/&�4�X�홡��Xp3[h���8$���s�wTh�l|Z�U�#Ś�y��cT��ɴhdU�������{�#˧���&����8�IX��m*src�-ܔ����ˡ��%m"@��$ ��	5����3�c9��H��e�,nN�v.ը@I뭆p�|V��Y�]��e����>�vz*�)r�K��Bӑ黽1_"%�Ӄ�si�Ǝ�l�}۹V�ό�f3�7`p\�4�Ȥw�S]�x3�d����<]��vd�S�M݆Цmus�����G��\�t�Fě��r��������CN7�d�hWo`k�W2��ʻ�#0�vt�u� ����c�+���.	�����kF�
���n����˂��
��G$�o��4�9��8��YnŶHդP�,uRv�|vќ!������GG�T-��ث(�z�ŀ�iS�L죎�,�S��U�|�q��l;܆��K���:�+7�G�T�{kt[�+�W�^��@N��23̱]��Cz�C3M��7u3.�Ę�a����K�t���2Ό�\b;t�v��;Nr�F�Wͺ���f{�os����:w_[���ne+���z4�өR�r�EU��c��St�Ҕr��!�Qx9�D͹u���b�� e\��r�S4��O/j�թ��c���Ioeh�;ym�1�:X�P��l�;+_
uZo�v��~u؁�mU0�;� �����w�Gf�h1zж��ۡ�C�����8$@OI�1)4��X��g�jr�Y���7��	�꽝�\n��Ռ1Ц=�y�^ZE�æ��u�2嫨$��y�N�Ձ&�n�^!e���ʍ�CTxN#���/�Y�t{�VlS��pV�f��x�5Ӭ6U`�C��j0�"���\�ۛ�X�	�y%�)x�3s5e��̗y�Y)8�j�-^p%�{g/�'0dޚa��j�޷g;;^��8�ڽ��%��Q���,#!�]��U�_K��r��p�Nһ5�RX9����������������ᝮ7a01�X��K��v�d�E�۪��nev���7�f�\��%k�M���;���M�0A�7��KV1�eفnek�03w/�"�qػuS��W;��,(�CmV���[>�*��j[DA{�h|�3'[b������������2�l��m�����"�X���݈$�34f⺷�f�_.زV��#/��p���3�%uf�;�x�ɺ(��_:����W��pntg$�R�F*�i�_�Q��b����v��/��E���}���WR�ӆ�C]�����ա���:�ݵ��u�%r�.d2�p���77M�6x�����<ܺQ�V;�t�m#G����X��N���]�J뗳y
���tv�=��_!8����_���,
�LN�i�λ�YV�⥶�qd�a�عk�m��V;�'�L�Nܔ8�(�ӤNj�X�y[&�S6�'����亨�i���C�.�8R�r�X�x$��ֲ;gm�J������`�G��M�F�Q�ʬ��6岲���&�<�4�!#Kr�PV���nV�Ꝼ,YB�{��*ʽQ�xo�
���
�yM�K�D\���"���0����1&���̭���1��FR���G%3�nH���y��t�a�]ufv���tp{�e��qhtq��޾5�1�ڙ�%��Oiv������\�_{���㰶��
���:��+m�.=&Jǌs�­�3�𳙺k23e��뺤zj2��'����MՇ��f%آE�=��p��g���lc�[��M���j��wB��$:�Y�WoGׯ��Қ�]65�J�p�֢Z�;�I��`���(ku�E3���D�NH��t�7��ګ!���(9o�W^�9��mJv��rƩM3(S��%Z�i��r�w��q��Z��x�&e�4�U�۰\7U�w
L�k��Go��kZ4�b	L���P.]=�a�~�Wh��7*l�5ցx+��s�6�M{����p�P�m_vw��Lۇ���vN
���W��ݻ�	�V�	�,*S�������d�#vv�±�k1fN�	Y�C3���a��f��`A��P�4V����[{qU݈p�6��yX�D�q���gaª�|&��Wu�v�-W�Y0��SR�����K��mC��RC�v ;��ǚ�[īy*��W��U��,4aXvS^3���{��M^��Szd`4�������.&�ftզ���i��uV�T�6S��_<��<Ps�aQ�6C�m��u�\�{;�\T9]��C
�w.ľ�X���J؛��P��+��ݳB���/mQ|�Of���(Ña
�MO���yJP%T�i��h�U�y�,�oiA�`wXn�������9�vs���� U����~_�����ҿ��������W�G�{~=������������=�����=====�O��4��۲��[_[���?7�(��$���	I��YBBE5#jF��ʩZ� (D�؀�2�F@�D�XI)�P��ʅ�
$��P��I�F��
&:	�TÆ}��5)��}L��F���h_
�����D~<>5�.��/�Z�x'^��;�$\���b+_dLghNwlgH��vS7��Z������-6tT����hSZ����Yb���iRi�nq��v��4\'.�X����O2ˡK[������b��$�^兜xڠ;.��2�YSLu&�����:��$=r���l��Nl��dʘ+V�9�u���uLUm	���Wj.����fڏa����C�y�7�b��	v�lN;�L�����GӋ3���3��q�#� 6�av�wZ����{t���9wJ�ݬ��O�d�c]��yǝ��RY)�÷E9V��<�K��q�v>ZOt��Y}T���Ԣ���N��̰��� �FbMZs�R&�:<LC;���-l�9TĠ�XmVvv�%3M^k'���We��<�j��3M47������v�R"c9��Mֈa*���l���ת�\�]�ԁ��ا��Bv�tL�à�6��H=Xm6�������f��qXw��UMِK�ɶ���՛�y��R|��ҷb��t0#�C���c|�*UڱΞ��U�{{t������̀Xc*���F�#]2��a
`��>�D�E������M��yk	%k*2U
5O�
B���7�H(
HQq$ㄨ�4�q`(�Q1�HHj"Z2����1Ķ���t�"?�PH�A�P! D��!9PO�	���7�I/�D��n4ԥB)$��fc�8�? ï�&6�1�e$q'��$C�Ěd�фB) ��Zh�r�@d ���eE��m�A��Q}"d��'�(��!�26ن@�A!U-S�@\��\��Q&!�2�G'�aQ��[�mTw)��6���:�:���]Z�-c�(y�|��E%'#EEui(b{�qʂ"�G0:��:��I2h5C��kN���I��փ���`�ss���W"��U-�h:��s\�ɧ��M$9rB��Zy�DJ:/�CG%:������f��Tui(44����kTR�����W-��c�C͂��4U-6m��A[b����4TQu�����5����κ�
fZj�QÙъ��g��A�"^AN*()j���m���+s	w͍z���1Mz��^���т
%o�w��<lE�	 ��.2PF6�-2�`���u�!�5���5����}eo#x��ž��]���v�u�u���p;W����.���������d��G .���10�m�PhE���0\!HX%HT$���'�|�o��6��e����V	I���	���E��6��g@/y��؜����7�]}�s}����<�'��E���*�Djq��5�3c>�/O�7�B�"7�W:>�|쑮x���x�&.�7^�ϫ:��V@�����-.���^q�@v�j7vo(s���Qa��:����Ϯ��a�Z�����wswѼ]��]���$!�sw#�37���L^��'L뮗x��#B{�h�wo��lwb��ee<ڷ�_H��>�r;_v*�^Sowd[���曵?O}�w^C�}���$T>�0B�r"ǳN�M��OI���
jw�J�������<�=�ؖ}ښ��_<YO5��W�>���~��4���'>�������{���*�K���\g$�mK�V������m� k>�{�Ӎ��$߷sԃr��y8ˉ;�v]Um�"�vL#��^��*��{�j��5��=��:��]L,��}��'pо,keU�����}��+q^v�or��t�/j����u�/M6lӥ��e7:7u�4�Фtc[A�'�:�`��n�n��a[�OX���ֽxN�۶^��ss�m}_'p'7+��B׵� �F+��]t�]˅ә+sv�.��7���%\B���q<�wQ�홉=T����z$u���-��Sd�^�-^����t�A/����*9����g���Q�U\�,f��͆�JnV�v�lT>�φC�j�W�6�lN5��V�2e�6]a�۝�83���;o�v����/�ϡ:�=�+�viuD�f�k��*�d�¶�|�q�p�k�=Uz\p��t���L}����sw������I�5���F�[��wۄ{s�=�*t��.$Ũ'�#��@�j��>�9̜#��9=_f��s�^}ݜXQ�b�<grwtjr�m���o[Y���n�|���3�]�]>�Չ��i�l����È�`';t15�{8�lј�����ReQk�ﱕ�Y�d�b��}�֛T.p��n�u��co/Jn6b�$w�+��'Y����L�M9Ӻ`}d���|�}��Ew�z[�pH�!&�9�tN-����k��غW��d��h{��W.�K����~�x�i%I��7J��������>~EX���z�����A��e�I��G�k�z:�L&���m��:7i��u�׶|�5�^bn�Y�J�w�˖|9P�ZR Ot����	��
��20!]�L%C��s:�-$.�We�+a�&,�ߒ͵
��>��!lX;������>��� �w�������^,��g�����ڦg&�}��V`���D��msޞ�)��J[����ɼs۽s�w<���?��S���B&4?)�t��#l��oG9�s	������=P�Q^�wP�Z,S���&g`<�.��imR�:6�M̾w��d*��i��C��!��b�@����r�ʇ{���P�^m�����i=�it��(���V.Ϸ%V�%9�]�j�\�V�}��9�����l1�u"�'��>�^О�����˪�b�
�/�s�}�����4��0��`6�wn�2�Yw%��[L���gX��|#�4�Uj���`���(��k8����h?�GJ:��4%Bd��ө}��r���!�����8����bhn7}y��uj�fe�"��@�T�L��Ȕ�ۂ=��}�w �Y3}I_�t
�=�@�J��.�`>:�M�&�m��y�G�bmwN8@�<h����&E�w�c��u���<��|=�u���4�$�f��k��uW�I�̝�'$^�ȳO��m6��El<XB]ظ��ws7�7�/:Y�`�6A'���ɣw�-nξ��1Y���o^]v���sS�ا�\pO5>p铡�]�YN�{2�y�-p���#j�qN��ܭ����m��SMf ���b}mRf�
/�,�hI[�7��A�`9Xm����[�pv�Z�p;ڊ��\�Y�Kt������*�6Q����=���SF��:�B���Y�&�xkDV�'�]�@P�����2�� O0�7�����*�~�ty�WL�n^�rc�p�W>Ϯ�D��I>G�T�r9M�rQz�����_e�M|l�\�����+�u���3ug���V�g(ip�mcQ]��[��^����][��V�8�_t�Qhӕ�D D^�}h���][0��&E���:�,U��0�mg�|/o=,Y���N� ݡ�����5��.�9���c����ǻs:����"V����F��i�S_����_�y��V�S����ۚ~��|�}X���v�[�WlwS����gl\pZ=/"M���@�����8��Vx$�5X;iP�XUq�ʷ���;بo�N�|��+���K���ޯ�d�l�7���F�:�Kh�GBEJ��co�ѱP�"�v������Cy���3x��]���$�7��UI����ɕ�W�l{r�s%�� q��TͲ��"�h��=�1= ᜯ^�/"�d��;�&�7�
=9KCp�p���rI�d�M�5r���VS(vl%��#z�f����:�pu�{�`����Ӈ�L�S�v&$��R�1t�s����ʩ�U��P�*1X��H��3���0���ɟwϕ?�C�v�3��gQ��n[������}V��̠�lv��UQ;��wP$��v�5���_U���l+�'/G��?jǜ#��"��!�+�)�z�U�����ug�����WR*�df��n��y����ig�VU׬����8RЄ�@w��(�wȝ��qپxOnsZI�훭$	Kө7�ڛ��3�X�s��4�
ʏ7,�	�fel��7��%�fe�d�餹�uϜ����3�䕾�+�ԫ7}�.־���f�Z�0x�h푸���I��a�:k�{���_ܵ53���}� ,�ڸ%lL���E�U���1sH��\w[�z�����̅�{��M�d%&.yg�!!ǧ�נo��3����<��#��q�W�����h�<����2��������[ײ�{�������Ħn��r�ځ�wi��/���O:�o��wK;Kw�*z_f?z����O�l����77 ��?�DO19��Hk�k�WzN��s&~��o]�/�;��/ ��,��l>��U����b��^�=�k�N!QE.�>�7���4H�S��s���;�G�e��쒦�q��`�AmN�5b�n�6)]�����\pOcg��E�D�� t�얩͕�nbݴ:���R�[��m���4L⢉L���>ܔ�;��:\������D[�<I���E�}����j%�#�LvN��w�f�L�p%3;E�٤�ֲ���#ת��I��]��n��ns획XB��W|��&����uG�_e�?��F$�n�0�j7�l�j�.�Ԟ}<�"쏡�9�x�Y�3%�ʩ����co�����1�Pw�r���rέ��ݪ����p���kxk��_��ɞ;|l�j��/ހ�3N�lq� �=�0��77�[�1z�����f<E�d<m�a��r���Z+u�ۤ�74�̿�"�ͩ��s�z��UU����&�٬���g��>�y��_��7�P�w�Ǐvt��g+�==�ne�>M���
�g�{|�v�z�z�y} Y����u����{˷5��Ӎ�[���#���^s>��^ލ纄��GOu���.�Wq�U��NnY����ϡ�3��3�Q�3�/��>���[�����ؠ�WɃ���jLT��7�H'�M�����G�gx�g��e;���*�}N��O4�m|���
�����c���f�F�*���޽�zS�aAێ�yn�ӂ#@1���alਬ�w@B�ۃx_�A.�少�4ڗ��H�ε�v���hk[�*ii��ʚ��S%�:��v�f*������$S�����5�Mp��D�ˊ�޽�P�(����n[:�c�������Cv��ljj�����l$[9���ؾ�JZ�&5�q�R���n.˗nw�D���M���劦t+�!V9��AUo�뭒��}\%��M�c9�|&iI���Xg�7�{E�I�/����۪����cH`��a��-6���!q�����o�&6�<�򒺬�}W��n�;�g��
���F��S����ݶWm���W<��ݪXg���z����ݚ:j�� zz�n:
�U]��sϷ��on}��<E����SP���슘��e���}:+�m�r#���T�J��ws{׶���B+:�E���N�Ȳk�B���pDjs��#�c�y�*�ul��҅,ܭw�����g��>��B̭��ٝχr;]_cs��6�Ak������-Y�:��*zU��p.a�ւ�tf'fm%��"ns1]`�����{�^'�¹�z�=�X��S��x����>H�5�:]@wS���޻������]��,��@ܖ�qf�V
[��4�2��4�X�еS����	`b1�+=�7���	S�ؙ�8	�Vo���ߩ�W��T����t�o)�w�{��+�B���/�v0|9w��'�@���y[��6������z������fm��WD1��:�R܇θ�ɵ�Gv+�)�5�Ogk�T�GDM@�5��T�˾�]-X��m����̋|V��=��g�1S��= ��=0m�w\k�8�ɮ���k(qw�y3�s�E�z�ꞎ�ە���W�!Bb�|�Ȩ�_FF:�E+��&5*��]��sؖ��b|�sp��\vcsp;UIw�"u���]����3�IL�x�+er7��Y����c���a�ޠ�Խ���<`�O��Du���U/�8�+&�^;���8��ٖna\3�6�t_���]�����L�	�Uϵ�N"��Ŋ���kUN�c����������Í-��%�廙�g�5s5��\:ȮMb�S��QHGF�k�+�s�Ռ�h�Y�#sf�W�=���+>�şcve�O5g�V'>@��_vlR�8��c)[��H�|ĸ��-��9lZ�l�Qj]�֍':/[�����Y��N��$�y7Dg�[z����{W�4�����۝��2�]A��-��fɻA٣<j����+�Kt_�ZnM�7���$���ؚ��Z��Q�f�{g��Ɉ8K��W��a��q��Or����T_csٗ������v�\k�ch��UmjUۃo����*�>�x����YYO%��������s������L�;�"/9��&�����I\wqY�EF��Ll���v�3IRK��
�/���4𽅚݌�ˣ�e��ՑW�Dc܆�wvV՟O����5�eP7ά�T�{����Ç�'���{�/��Q�^�=>����3�����\;��`���.琢)^
�p��X�YAZ�.��GWN˿���"S��<�g��rޫ��ff�'�I\_p%o���sZ�0��<��|]|j'��ր�z=�ߧ����=�>>�����������>�������z=>�o�����kE�o�9����#5ݝV��;[O/kn��:��B�ex$=�V8���$�9Ɔ��tm\{޲G�}X�.���1֥�0tŮV�<V]���b���c"A�#ɺ.��Ś�V l�x�ÄV�]��2>-�Xhi�+oaO�m���ur^	��+l���ޣ�ٻ��m=J��6���n�zN/s�.�<�o���'R7o{mPuuɨƿo'e��j��#���WGI��.lW�]X����Ʉ{%��E�[��g`��X���6!%OP�D����s��z���j2��仪�݅��o%[O��9]��A㨞��@���n�Q7P �����1�p\��k�W`����(=<h�tג_OJ<8o8�"sʔ���j.7�tj�5n��k�{�� ���ͻ�x��t9�8EW���<爻�0�#�ҡ�sn��V���<m�Na�ǃ;/c��������cۋT�[�S��F��ofB\�y��ܬ�K�����k�r�w��Yn�M��A�"]7��d��)vL�gV��9��Ź��mb:�N:���I��1�]�
5ޝ��e������,��e����R�l�z[̠S�@Ҷ�B�
����Q����.�<�B��6��:�r9�T�\9�av]��v��w;��Ճإ;�v1Z%����\�)�x�~���Ƌ��E�ЇZ�7���D��1��+xa-]R"7M�`10 ���TB�6*�Ðqۅ�Q��ܻ��ǅ���F���Q"k��v��m�Wv������-h���=x+�
3��+�D�ܼ�ݮӬ�gQ��g<���{�=Ǹo� �m�]-�2�>�xu/z�U��ę�]c7؎�>�<nlen�5�T5�mɜ{UJv�;ۺ̀pJhuͼ�����m�t�O\��Q���R�\�
�7��*̌�8ň�ٔ�Jd��O�]�$�`ɖ�/E�\��G�^V� (b�y���L�9���5��\��=#8��F�k��O!t����p�Jv^�� z�ǹ���|W.u�2;�y��e�]s/���gZᘟ&��z�Gɚ�� �=��j��
�gd{���Ҵ����cC>H��f�p\c�I���1ﳎ�d2��k����	������9e��i�w�a�woM%��S�b���������gF6j���ֻ ���OtmYX�'Cd�Y�臙��r�������}�lfU;�f��{9�d^Yé�I$\���ά�l*>� ��H�� �΀�R�˙�8�6�1m�n��Wd`�����ε��=��p:CY�g[}zy2�������b�p�[]��v	�O��6�O���>Jn�k.�lb`�-��	�)�Xv����D,9i��Jw�a�fQE��W�{�����!��K���&e��tJ��vV���L↉ȓW���Z���7������z���IKd�S"�������{�U�F�-���F �8�*&Zjte�ӭ���\���rŷ\G�4Q�����
����h�v	�M�⹹4p�j6�p��ֈ�X��9;8���-z�ͲF,��]n��b�S��j:�䙫��q��`�ۑ��j�W�r(����g�ryȭQ�mĊ�m�Q�h��󛞣*�t��w=pMs�x��(��q�d�[���z������:�s���f������7Y܍���'�-��A�H��!��L�� ��\���5k��5�U����c�G\�b�ۄ�s�`�h�Am��9����b�lX.u�Q�:�Û��ss���tu�9�O�;�U�N8�� dM]����J�Â���}`������{��N��nh�Vb���ۄf�����8ۼ��Vy�n_� �''T�,`ck�ܞ��L�x�*�z�9����J�:o�sY~���-MZ�.�t�T֪٩�n�D��ihv�;.�Y�0G#��Ӈ1S	��TFn(�^�1>
�+����G�3 }0��w�ყ�^�uY���2�Oo��U{T��@,��Q����j��{���e=�3��۔F|�h�E�pF3��|���l�oM^�d�޹��UQ�lI�j�fkt�'�ð�1q<�t��_G�����]=����cߔ���9�������n�+���Aq��HǺP�&�Q-ͽ�s-�\���a�[�]��a��cs��� Y��3M_���
�������b��y�����Ѿu���"�R��ȽW;�C6�?�q�}M/3���gT*[�ծ!S�e%K�P�!��k	}RyŇ�4��%���B���xkh��f}���۞�wYt3>�^h,"V4�}
���6��v��G�-�'TW�@�w�K���ؼxy�Ň�;`�⑏t��T�h�p��s焹�>��M"��i��CEeH �o?�콆i��+|��[���Y����NGL�!&r�_^�o����>�o&E��iAnc��>�W��9o+2��Ֆujq{�ivn��J�m�ۍ��ٳ{1�[�|ook1YilE�t�.���Ҝz�+rI@mR�l�Z�\(�ݴ+]�=��Ϻ�����y^��ߛl�8�w����d����П�ԉ��P%� ޵�p��O
�oh��=K;[�<�ӏ�>O�YM)dc ��`.�},�| ��ׄ�� Ƅ�Z���#;�W_:�t!t��ܨ���;<�Bz6}w�nx��>n���Ԫr'�^��N�,�f���L�� %���8^Dj����S�(ȶ�{"�����Z�v� ���h��UlГ�ڿbt�zf!��wf��e!�9�d{�z�4�7�:���s:�#x}	���H��1�+<�g�U�=E����~��z�MP�$Xt�VK61���`�������#��ݣ�kN��,}�.'�!�fq�l�Z[�STg��ϧ�G���(��fM��ƪ��g��S3olʲ�[%��K��T���nP��h
$CλY��k�X�#f )�d5c��!;�G3q�3e=��HoB�g�{N�l�,hS��#��<4��|r��@�S���9i�å֡����B�;�h�;���Tu��U6��y�Q{�s׬��n%�+�ZE�m+�M~#�����k�^s��7�]��ם�t<�,�<&�X���zf�˧�f�SVي�s������A*��9��"~���a'_��q{ ����V�u��W5�x_Q��2Nْ��q��Z94��0��PDZ�gj^IܡOT$�Y.�ڏ};L���:��v-1�h4 6�����n*������q1��;*h��{�2/V����P��%[�-��>t�1
�e-��Vl�i�͇c�����ơ�8�,��1i�]|��<BO�G���e�s��޺˾���ut�$ip4��();s�~���2ʦb���K��t�l���p�޾�U��=��:�β�g*���,%w?QLt�IW�Y���of+����g����1�X�?9Ϡ���E��ߖ��+#oJ���٦d:J�
Ԧ)�:�,����J��Q��� T����d��kV��e�¢�T��!�ߓ�y�d���ɗr�sH�d������ߚ�_����3?mW��ȓ���٥�r�S��+�0����@�4+yHa͘Nm�\Z �������[��2V+��m���	�<(�D5�0f���<�}Ne�z������g�����r�ȞҚC죝�=�㞡�1,쒍h�������|[a0����\�&0�X�����5n�״�d������TW*lt�Y��U<@/X��}�	�)�GS��rl�*�XXkd\z��ǨKeٙ��zj���#=r�3vl�5R	��1��F�2�oV@��u��{�CUV�5s��%�g,���w�	��c}(gy�[֚7�l�݋ym��^0��[쥕1r�y���KV;P�3F9V���q����I���%��U��S)�2�<�t@�p4������f�
�,^���(p%�\��l2"}*p��5��L�I�[��{n8�fC��)�_��l�8��6�N0iM�k�?��eUʟ��
2=ڡƒ�f7IƱ1����2,U�fE��)�ڦ��&0�T �m�H���=l�@�u�iw*I�N�]���)����t^���>K�sUDKu���mmD&��$�Dہ&Fu�z�����EṈu�M�li���)��C������7�V5�)d�r��{]M2���ݕ+������~����U����@b	V~���H!��>v��&�
�����~��O5�,-;)�ݸ�S"�TSoZ�ecF����uqA�h�r�&e��|�Uź�8�bԽ置�q>��p.�cbߢS��]Kw`J���Pq���9�5��C���HO��rZu]@�����aޙN��P��C Z`�N!�ga�N,RS�u_��G4�`T�~k��
��rt�ܩU��l�B�<G�}	��zL6�c�������J�On������i�����z��K��۫h�uzߞ�t��4��٨7���;�3"�W��2]�OiG���V qX1�T�fl����A].��ä��}B��2V�8�!����'mKO��Y0��c�M�'�P��e��]�l�#x������fK���_��圷2q�S�@cmm���c��u�E�s ��]ʿ��t��?Ez��s�j(1	a�(�b�LeE(k΅�Q�'Z�;C�'zƂ�]�(>����ȣl�Κ`���K�t�T�#���̽}�2���Q%�/�|�0MV7�v���`��b� �d<��E�K��N��9)��J�&{�\B�t!@֑}*�p7@0=���`��S��\-q��^��t~^?�$�6�ʨ���{��3 )

zʇ� �Y�a��H��b/�������z�H������>�����P�<My�}�կ���dܞ4"�α��ۀ����C��^6�#�N�TU��q<5�ݛ���~����&p���%BOSQ�r�O��Nf]�_��ŝ����󺚙�qfuƙ׊S/i��M~�����'���)��,�����J~�}i�~�����'jj����b��(�)�9�;�o$��1��[UW�*J��5���ߠ��CW����Y�,a�i�mT�M��r�o2�x8�:d֞�hK*�l��v��xi���"@�����������v>~�l!Wm�a�H#+�76lhicz,�:��XݭƚU�`�=����.f�<	+^��6>)T�7x�:f�`�W��'Rvsc�,�X�)���Q���x���
�\3,�T&�����{�ӪM�=��5����Ιg�����u4�x/$H��@-}�;#�N=�E'\��)9��E6ג���:�/Y����YɈ��.�U�;�b]���E���jذ�-F�mPy�tX�(����B�ԁl5��=�QC�J���Y������1����O�f�AvO�Q�����v�䨵�*/΢|ަ�m��	�{Y��U�N�womS_�P��i�`�s�@ʦ����sԹ�l��wK���U�fvL�s=bV�m��磧韵�u9��;~�� �+H�kȃ�A~]����g��4�{[�5vOݚB��G.KJ{H�e�cڱ���
���;�Ј���9���w�s����[I���1ك���c���h��;<О�l�.���i;r>��	! fg�q�����j���W#ß��|*$�SS�x��T#;�Y�j�Α@�V�{�`h.\��l�cI��ͅ������1�3�p� �MD��|z�7��� �78W`��޷��0_�KU�U�~zW��X�׮{{D�< M�J����zb;ƦL�ig��Z�}�_���*�vA��h�dl8��=ӛ�[�M�=��=��+�w_]#a�$��36�8�u�:�e\KௐY����ޓfм�S��EZ�������j��pn��jF�"�X�����"r��m�?��/{�s��Vb{��q\'|k�M���&D��e;���͖^}A,�Ԣ-�_�����y���X<=7'�2�=\��%E3�U�,�	�Ӳ�2w�>O�����r��8�,�T�=�Sp�G�T;F�=�@NINju~��]��N��qM��������c@�A��)��Qn��7��s���=������j���|t�/Do\����D�M��>�[�̃(r)EV�P��ʵ�6+�����N�3�E�^jH�^��>���r��ë<;�|n��B�;%������g��㑸��a�D4�Z�&8f�f�T�W-�f�H}������)wش?Y�OA������n�)��Cv�ٵQ�F%d��s5T��>}��f���a��k�R ��j(�ǯ	ru{� ��Y���'��*/��tb�v�������.�p%�����^㰶/������bn���dX!��\���݂�R=ݛ�SZ�*.�FC�aVXX3 &)�Lrt5���+{�!�eX���������ck� Q�Q���쥹LǞ�Fz�\i4.��&�A�U�,7�e�g,YO�\a����?���n+�7�E��9��Ӑő�0Q�1�����񳗓o�����ĕ��v��LiA�����!G� �s���n�O�)�(��ou���<biF��K��)s�-�0�.���dy�j%��z�Q�3�۩���`-քR�Si:XN�Ec	��������6aݺe����c`��K��1	�P���n�{��ЮPaşڄ�r;�e�������PS�3+��V�q�,�蹯�1-ϾLh`��אz~��{�z(`6�}�T����d{۶&dڛ�����jb���7v��1�	�.��u�>#��DKl&[;�2c@J�`95�E�:RPnE��fUs�/�N��h�3 Alsb@G���Q�����8&�����+N�9by=�׵�z��7��e���
�,�Lf*�0\�:��4�h^Ϛ ޻ЖW'J�/Wmem�"o'ޣ�?�2#����+o���޿�T��Sm	�t���I���T&���^<����������o�G{X�N�\^>5u{v����r���p}"V��VإX��
���*m7X�P�\ò���^�����
�k�*�b������=�D���!6���Z��ˈ�G73��9����<?{�/n�c 3`l��׳���S��
��a^-B:UccXͬkx��w�����c�c��7u�U���b��jX��_Q)f)M�f�.�!�@7��!"W=6f�\��x���7YD�ʊ��%�o n�����C�� �Y�TtǍ1�PB�n��(z�B�H���%��/��d�(������4�ٲPx�\�ͮ�|u�����Z�B�gpue�iP�yS��-ݦ3_�7V�S��۫��_ϫ���bp�F��K�U�~�L�]�*�E�jU�~,���T_L�uQ�wƍ7/&~���:�F.=����cS��= �ge���ҹ��$�	����1:�����d-�fM���#a�q�T�^h/1����͚�?�Bu�Z��X;z��\[�TS�қ/͞OͽER��1�g��[Mz�qwHT�B�D3�\D'�����`��z��u����;'���-�U>d䯠�Y\�x<���*������/�`?D��y��$��ᲔsK�j�v�Ї�fX�k&�/�v�����l`��k\�O?�6w;���ށCO��E9~4"�H]�^��O	��c�U�sy�;��R��TS��)eyڤ��5��['}l�-n�Z�`Ũ �lB0ǻ��cn�UF����MOr��]ˋk[3���2!�����1>�P���ヶ���moZ�V�_.��y�-n�R|f=AQ���I~��`���nj �z�"��z�'��.:f2�(�"}�:dL�U)��J�-R��5c�a�}aBuf�/ ��#{���Md8�'�Uk��,�v�k(X�%�bn��ʹ]Z�,�Ƭ�� ĥ�V����q����c�wV��fks�[�Vwe\�>o>��S�,t���R�u�L�oa/�˷���c{tYN��6S|��)A\������V#6s�\J�xƽv[? >a��ھ�H��MoF���f�1�s˾��9W���y����V�~^�쯸�7S���S�w��#$O�ǫc�CI� A��,�W[Hyn�=�N�j��5Bv�yP��}H�G�����o�e��_M��V�_��_��r�nx���mz�W4٫%����Dp稈��!�^�U�"����..�fQ+w��; ��.�P�3G9�d�J%��V�U6ߊ�ֻ�kL�h��J�}�wUMy~�2��Ӟ��Z�?U{ ��P�u��QB�8��N�緔�u�`<��Jl�ٕZ�N4��7.�O2e��Wa;Y�S��QMmB�]�hdph�S��k�y�tI��O�ӓ���l���g���]s�:4ݖlRÛ�ˠ�[�a���\00������]:��/����� 5vn�ηy��Q��7�2�i����9PI쬑�U߷5�*�ա����\^�Zg�����sPoz��xc�{y�6/q���|�7��lceV�7���Xc2�4"X���!\�oj���j
z/Gr�-5ҫ��uBhN�G[�����[����~�ؾ�G�?O���������Ooooo������ool�����zzz|}$eF���w�s(���g�K��p`YZ[w�	�SzָfU�K�`��O�n�f�kTo2���a�������(�E�\���Q:�f�g+�.�=���-m.NVѷ�6.��;�kp�`��Z�VΙ�4��θ�o(�5"��[ٍw���m��E F!�h�!�k�� b(�n
���S�h�d�l.{�m���hY�6�Sh�֢��%�_�¸�nVj}�U���n^�V�V,��LI<�y��7�����b��{X�Z3�9jY�,.#�)�0��\���mr:y�
�K/J������Ws�ʷb�A�p�1��޼���w�❄�sF���@�-VNl��쾨��ֹV��^��ä�vwu@�i�ŔN��u���bg�\Y��a����2�u��\o&�L�ċӊ�..ki��=�j�)�# %��%uu���˫��:0�mXM.3)��j���j�Fm�����3w���[8�'{�����8�ihnu-��+�a��ݢ�3��8d�ϵŕ�ӶŶ ���q�h�R�vTy�n5��4��s3��Gc}�r�[���B"�ݍ��L�{��q�2���UD��q�!��Sb�r�%��p,�!|�'�[��\[[u�$c��/jq\�(�^�vjz��D��f����W:v��:�k���s����0��`��Yj�z����:�"��I�@h���F
��*|��J"o�(�<�^%%����]��8����]�N��gִT.kQe[��H��T<r�!�T�on:�HV�!+wsu54bh"x�K��i-۩{5Y�3NY�k�j�$T]r�,�vs��Wd��c����Mя�l�0J|�p�/tn��C��1�Bc;!�{a�ӗ�sWV�;c9�v���9ʝs���Ҭ��9�����y���\�Ho0�IXH5A^1g\��z���Ukc7T3D���a�$\9lDM�+�G|�v�a������1{�s"�(�K�W�y9��Z��/k����*���/���lpj;��/l给��������d�W.�o.w�HN/�S��;n'�f&`��v6HpnY6�q�BD����ʌqQkeӏ�}�c`/�'�v�R��Nu*O:n��u����>v;���N�8ɻ�E���Qt~Y ��4U=r۬�1����ˮ=^�w.]1�smH�N�󤖊�d��w�s��rk�9;P-;���J�`x{��n�&��7i[���L)κ��;;b�AG�-����l�w
�hE�&��Ӣ�3�5�˅����J�����ƍ��-Tͺ��u��Ys�C��Yl�vԨ���Xcll
���@��b���2&���ܦ{���S�:����ڊ'�We���H�dY��}|��˼���@�c�l��"��+Y��fY�XWU���;E�f��-��i�o[Y�I)3[�s2+�71��s����1�tX���s�l^z1�lUuWk�u��[���O]\��p2ng��'-�ˍ�(�Ǝow8H���'�@%6�) ��O�������HTA�}�%�@��S�������k��.s�ܰF�F-��,oS뮈�D�Mr���GF���"b��_jE�B�Bd0
�:���4{ɚ�깎FO�q���6\���.s9<Ï[td�յ�|�C�Y��	V��(�>(�,�H |�C�D�$a���Hb$�ӕ�����ÉA,�JZ����A H`��@bo�cd�I!T���t�^���s�y\��6��m��H���'Q5U�_)�!B(��-������Zh�c�Π�D�1�ns�d����E׮z��=\�W6�e�m��ڳj�#�����[��8��O5��%O8�m�[r)M�uՠ���u��F�գN�G�`�����%G�r����Ǩ�­�s{�Zط���[E5�.X�cFg�}��6�[(����끭s��nEQ����嶶1�����sS�:*�h6�v���~%W���}�9Y?_"1a���B4T-ژe��jٱ1�d�Cv�`cZgi=,��y#�S¢�m����9��/%��5 SW�����bz��V�d1���ʚjZe".H��6�"$1����nO�G��עϸ�i�(�z<����j��տ��cK�
�p?�TC���#���]/\f7��~�m�=yfϡ�tL�I�{g�l}o4��-Q)N�}��3���k2�)�|���塁ۍ��cL�o7AN3����K:Di�����b���ۮN����NvD�BCcFD3<(d�;ey��W��� f���W��p��O޻h(U!��ܻ�S�e�V�+�fӊؿ	�C��x��ô��f�� :��d�cl�ݡ�)��ʲr����զ�xwm�D3Z���'��|��wŲ́���-1О�<���'_��k�����Z�]wQ}�R]��t��vm�ۜe�-�!��y;s�B5�F+�g��ty�ڦ�8��������{�3�H����F֯6��zN-���fl�5^�P�Q������׫@״*o��?{�y��T�<�k�]鏭y��UDmd�P��\�0�0�Z���A���(��+�;C�c
`&�3w���7I��-L����*}!�Q�z�����
�_L����#��d���n[����/����l)*W��^2����z�m�������0��v=A��7��N�C�gnY�F1l���soP]69p��E��h��XtC���RԜ%R
`z��GY��[T�0���i֥�i-�\j��f��wy���M���+T�%� �S�)�*���ZP3t)�//ӕh����gkAt3\8�-�W���$��'3s�C���|��a��� ����7�xţȫ]U�N���"lb�m�j��Co������qM/p *_��	��^�R���鳪�Y�H3!]ʕ8S��)�?`	O�}H危'�[�)��ރ�c �s��5�ny=��X���ukk33*o3g:��6����)�%S�S�T�G���-q0���,��p0�v�{���;i6a�a�KŶԟHL���z瑺��2y����X	,X�\�|{`*��d͕</��M�Vա~T��K�-^9'����1{�[ʌ?����
d��7�u��vY���9�;�\R�qj�OE�6�D~`�cy�f59�QL�6Kvwc[ՙK3�:U~ⷭ�W1�z;iMo]ܣ�V_���=��u�Z��o�ľ��;���?h����"�����I���s/S��s�V�S��j��9�.�C��@�����מ@6Z�����I�̍Y�*&`�N���::t9�B��6ZW�`;��ŜϠ���g]�\�?���C���?I��a��^���C\���6��BnV8�4I/cj\H�m��]���-�n�R0H*m�O�M�'�7�����pۅ�j�MS�k���zڼ@��]�Puz�<�rk\�����	�"�dۄ��F;�*��:��H�~�O1T\��|.'��A�E��0�@ܛ�_��s&ٖ�N�wn#y��V�U�o4���,���zH%�rcҵ�5�;&^����~,B	@4�B�-
�F�"�wWtD<v��/?DKX������}�ñ;Q���56fl�0�����Sy���7�	���7V]�D��(�RAgTd~���(r�_�+4���㚛��8Ƽ3�Sk_��&��7�:��Es�#6n�d�|�r0���(�i{@�� h�`-����AP�j_�����}�R�t�lO\s��{K�vp���̒�O���y}I��̱v1mD8��\��wĳ��	�������l����BAu��l�s
�e�T��f�U�o{�Pº��ǵ1���5(j�tuL�WW[>�n Ld���,쇟�G���It��M܊�n# ��I�c.�sp�g!�$v�����ּ��6�3����͒D��Lx=�EŇ4���`�#����ˣ���Jp�ĩ%Qת����lUō�#%H�`�A�8����w�9�Kx昑D���]n<&m��Y�t��y�tk8֧�����z��+�4<���`�����>��i~;�*e�E�-~� �ΐ��2r'�W"3]�c/j���@��Z�
-j�m���z�A� �� S�}�R��;���p[�����0�O0~���Zq���aQ�=���W}� ڵ5{(�����[�+a%�SeB���F25I��%�p�6ͺ�B�ni��Q˶2�Օ���PH���,�s���qM�,�oVI���	v7�����,&�껾Q���}|��׺����!��
�B4*R� ���������{��J׵"O43��o�r4�]�����\�/͠�\�6�w����c��L�ئ@�;��Ng��}b|;����Pf�+|	�v/O������\-q��^?%^!O�-;�zsHo)��������0*z0�3c�Ǩt��F75���.�zF���9G3E�����U�
Cq�)���<̡4K��-0��wl'v��7��b�zT�Y���)�y}3��.�^��~~���|�O���	3��&_��˾���/'�s1��SW�]m���v�Y�{fk��"����f٪�A^���������(�N.��a\��m����2��T�4�曭^���-�T���k�����J�̞�I{*�s�i�L��>�L7~P|���T��,�ya;��&�Z'�ׅ�)���&�os�ּ�A�W�D�mIeSo-��=V)�xk`ܠ	0M�x�5Y�JT���Y2�L������y�f��/H5�����|���o�k�%9�m�3;=?\�R8����֕mR�,�v6���-M��m���dk}RyŇ�4���
�NK�|ޟSp��]q�z+vYY��3[7B��	��ކ�`F>?>�33i\K8MbX�����:\�J]���S2���e?R� �-��:�\�K�rN(j���!��V�V�X��nV��z����[&[dݝ��u������%(-(�*1%
�T�B�$J4H�- "�0�IH��ԞV~{,����w�\!)A8���*��`�oW�&}�X��ǲ��q��)��]��\h��giܕ� b�aQ׮��.��U{N�6���R���^����Pf{����!�'��>�9l���Rsp��u��P���J��w\�K�e�b�tkmv��	�����C��j^;�	���
x��:4d������s4�s5��|)�_Gk�T&��3��qz|�atr�׉#������ ����k�KM�s`
(�Z���LK�=s�k"���@�hOK6}D�4�S .��q��/]&��O2o6��4���%�~ (��ƾ�vy��_������'Vxж�t�/�9l�ۙ��sVV_{ITZQ�~��HdCO�1.hl��͊@enNG�χf���shsy���M�g#�u���5�V��:����%�>>A/-�~�Q����I�^�銡�͔彷���D*J��a�z���hs\�@z\�?HȾ����`3�:��=�yw�Oy���H��)������9�5�]��OgV�o���Y'D� �D_z���Q���H���:<Σu����yrF�E=>���}u��r-V�t언<����VnP/�s�Jsp���F��gy/�R���6C|���[5�]�[mS�i�]�xƘ���}#��˲�I;t�L�89v�2g�X͢�$黢�%9{p-�ה�ͬ���N<��� 	|A ��
@Z !�("EF�(��$�ZA`�R	P	eJ	�����\�z����v}r�5���7����Nf�r��A�?��ߠ�+��1%;���/֍����a/s��{����R|}B#��	��W.����)�}�2����M��^P�\�{rd�۵��9۲�JXS/b�m/�)�Kɥ:� ���,��u[Z���ۻ�2.�b&Z�F����M�~�=j N�8�����[P��ݵkŷ�M�5xC�H�,ԣ��Zq�eP��c>Lds���z�嬝L���ywq�ơ���n;��!7 ����hOO�>c��)y��{��O׫h���hdP�v)�{~�)�2�e���t�^�s�:����&��s�-���>K��W��H�B��{G��/�"Ґ�������Id[�`4�}'\(PZWl��P�k_e���r�;��A�9�C:n`[��[�<�ёTpї�Z�a~H�d��g��n�ܙ�r'1{K.3�WՓ�H����.����f
s~�����/L����Í��P��A�z�Ӫ��H���X�\Y��?{ME��"�Lh`� ��07�}#���N���x�����{��.(豬{�i��z�����:<մ���ޏcD�2=Ѡyr�Tw��n�0EK�;�HO©�km�9SM��ޖ�2�tS�E�߻��P���u�%q��1�4��rקp&��=�vV�7��ePw\L���6�j$�dг�bsQ��}�z��� �P�$�R�B1"R"��	B� L�  4(��(R� R���{����`�ζ�$��jg_�P��)1�����*�mn/m�0`4��u0��!�C�F�\s��ޮ�G�TmZ6)�����C�:涜�8�Ο�)�?�zqبz�Ƃ���P�	�$N��`�	o:h�}|�sB_2��żn��S)x�aY�����j�P�+�'�WD�b����Y��z����*~���r{�LK��A��DW�t���E�� �Y�D����K��ϻ��K �i�	�~n-t�5g]i�g��[Qt:aym�ዏ���ߘq_��,=��k��Ig������l��[�J�#��q��,!�*���ɩ��<��:���>5��z㚦���F%v��d�r�j�MSf^"������W���q��b�;���7��G*�� ��;6���t�_�x���|eh󰉳��Al�ɥ���f��/�ئ�u�����Y������<G�"x�@A���kZ�j꧒Mټ��k:�Ӯت��.	�4��HA��t�k��wD&X��&�7-Sm�k+P*3&z񢓀F�[R�!EP�+��k-lۇlS|��5�� Y�1��=��酄�Sw`J����:���?}��~��Wΐn����p��\��1�����B_3�����Dag�?�X����;�r�Ѯ=������`s��f�P��Nϴr�^����N;��n�[�I`��V�����.�CT�1����� i�!�&��7,-(>Ȩ��0�kqk�ܮS'�~��
Ј�%��R 0�BP�HPҠP	J�P"Ģ4�@"�ϼ ��`��u����x��j��qmA����.��'�&��	��~��j�X4����(�0�݇[_\݆�̼յ\v�ЁY�qq�'�^S��V�O�F��R�e�μ2ؼ���^7�Z��Nc���c����#���zD4y��9�~?4�|ƆV��"|E6��!�����(3��S[|q��mY��\��H7!@Lsr��
Jֹv��O�;oS���7t	�p�OI����۰��r3���{c/,�}R�[~��)�s=���Ȼ��L񸏪��R��9�@�On��.��X/q!�3�
��'��=1qJ��
���W�GGqK;/7��SA�G����CM��|F��`�:t@�"�b_�XH�X�T�^��ls>��W�����˾��47�m'ܪ��p���ՇE���a����0в!��M-!d兕��w�;��w���u���:'2f�M��]ϵ�1� X�u�/ޗO��%� 9
�L�ߟ�T�n�}<�7^�&>͜�t�ʚ���̆���`�b;�ϼ$�0ƟjX��˧��E��c[�١�4[��_��څ�ȿ���Q�쾭mGjQ��Cu��:x��}r/��0o�u�\of����tK
��w�`�߹�t�{{C{�YUc�_	��ݾ�!�F��9f�nѹ'w����;�d��6�/2�"����4Y�	��Gߥ�"@B�F���Z P��% &U���QX$~��뗾ϣ�=|���xQ�"���7d�"k���
��a1>�^�d�T&l}J�/VӰ�QqUp��2("{�y�F��d�[ݝ�S:���Ԅ��y5#�.�Z��2kO[7�K(
m����Ʃ�xb������W7=����{�j�0�8���ݩ4Z���o��I�|��߽��6Y��G��k;gJ��s�=Z��v� �v7A��4�5���Aʗm���XK��,?I��W���c1\�689�����W��yדKf͈��9ULa'�O~/����o�d�ӊ'�1N{���Q��嬃���>���(��G(m�'(CJ�վ���] ̼$���W��#J����=˳��y�0�z���j�$���=ܢ��n�v��WC��������{��ݑ�?ߞ����u��%�M�2)�����r�4�H�e�̈`�)���;�i�N�&pڨ�K�25;0D3;�ѐ�Լ� ��z��"��ܬðlsrzY��&�<�Fk&�J��=cw;0�O�V��DF3C(L�r�d��1x��>��#k�����l��^��1�\q���O|��w�\�!6;��w.`�a���)Rج󋥱��/��+°q�yk�"y�V����+2uѱ����s0���>��e���R��=�^	���t�HEd�a��T�Xy�o4]	�hwz��ZQ<��u۲�n��b��e��ͼ{�h���n���<������  � 	2"� ��D)@)IH(� �40B-;���N��y��P���ֵ����ɨ`�����v�>���ƺ�5��ߌt�Y˱aݚhY{��Ͷ�ڼ
/n��g�=%�*�`���_�E���8$:b�Gt�`h��M[$�����3�3�jj^�_���hu��ށ2́��\��b-�����޽�㑾����g<�i5?���;�M�\�f�!s�L��;�>��v��E��5:f���`J��EC��mP���Gu�n�k7-b,�����X�r�-����W�f+'}681�����P!���w��uͩ�=�[��o��F����.���~k}SvnX��w��hf�R��A�9�]e��˲rV��[���MW�hC{S�(�nF����`+�~_O�8j�?~S�ʝn�!���K���O8j)����1}��1��3i��V�6\Vƭ�aC�u2��zyd�;-g�,ȋ܌��S_�5k�ɾO�@?L�� J|��V/^�k2��嵲�ck���y�
�MF�Tۑ�&lK	v��l�4�2h�2�V��{x��[��s�H�H�r�ƙ̮}swo{�x�s����~�o�����������w�����{�}��/}���＼�Q�U�#��c/�镲e����v�F�hFv�9Q���JSv+�wXy�ߴ��|0&cdq�R�s�c�d��#�%�o�ͽT٫��r��͵�qN��G϶�j�5��t�����i��z�61/M���K�{�a�s�/�Sg9���x�1��%_-2��u8ހР�V�r�Y�ʏAd.��ĥ�Ds������A~#{5�n��yt��v%l=LEP�b������;5��]9��}e ͺ��޼��P�u
�f��0�P�������$�F$M�xT�^>/�`�BhF�7�d'�ѫ��+Yc1��8����y
��s0��WcWpe����O*���g���slM�f�3&����]�R��t�pu�mZ�lԘ�{y���t�0�����lu�_Q�L�/69BTD0����v�*�Lۅ�D͇a�wS.J����3:�ֵ�d�	�y��f���4�ξ銥�^��I/@�%<��T��W��#{�PLq��tέ߫x���(���ע��b%/��W�(mň���$6v퉵�]ØS���;L=Y��E�4��vX�	�n��w��5{2�����>Kn�3�Z���E�{�-5)�f'f`�x�`��apHflD�V���xV�'`�b��{5�Lz�
���~�]���l��n��e�n�sTKS��U���*���b��/�3l�w��0�n�p���7#q�7"�[;�(K[�ݖ�4����fwRF�n�
�X�}��+2ʺ��e���L�RY5U�\��WR�/L0lc�l����Jj�gv�Cg�Axxݷ��^�`{�F��s�
�b�.�]���N��p��݃�Q��ټ�p��jejy�Q����u9ywQwl�i����;�I�T��+[����W�@�ɘ��������[o6ә;���W���7�1R�W`��[�sVY����scGp�6�PY)��u����H׫�Au�o`{���5�.f+�
�^֊sa��X��:��a������[�3T�g{����x$.�b��oJvz���Ҡ۷P���ۙ��n����P.���_l�Rd	��Ӵ_Ԭ�?㫌�<!�Ϸ̞bИ->�C���+�����j�t���r�Z����G�n�]��1T�.(.�^_1W��h������*�aٸ��J.v��t���.����כ�7e�(�p.�|J]�e�z�w�!���w#�.2���)ͩ)����v����9�yս���#���J�C!�*^��O��OY�� w��a�3CPn.����ӻ5l�h�0���;l���*u��gj/��u����[Ҫ�:G ��^�4�{��V�*��Gơ�yy$]��^CVw�u��q'#[#N5.]ӭ�Ͳ�$7�I-i���IM�E��8b5�yRp��v��S�����:��4j�b��b��d*-�P� ������6u����bы�W7������6��8Q_9��[ܹ��l���f�H�cm�
uD�3kM����[���S-��66���m�W˅G�r��
GPUdd�20$JD�O�������ڍ��םp�њ׮?Qʫ�T[ov9[[i(9�"�qb�j��;j5�F1cN""��Ũ�Z=p����(֦�&�b�b/W.Q�["���:�9X�l�V�X�/�1���Ӷ�"�Ź�r�fbh ѝc�W9µ�b#[�h���M[&���Z��3٘���U-i�n�s��smm�kSU��SW�GV���6�k�Zƴmc��������
�*(c���`����w��~��u���=>Ʀ�np�3�l�p�(�S{��2����e�(X�����L]��˘k���2�cͳ��c��	·��!Vd��@�%@&�$�����bT)F������_]^�M���x���Կ��|hO�ɐ��|s֘g�BkN�c�oy�y�(Y^���E��%w���
V��^iמ#�T�&��Rqz�y�ֺEsa�N8ҞaA.�n*���y��c
��Y�v��e )��L�����W��	j�����;������:�-�&.ܟU�Ŝ��{�׫B&98 ��M:�����<�~`��y�	�S��V��mM�O�*#;�#�{����C{��P�5��+MU6��w��Cȃ�������'��!{hn˴aV��u����l�2i�mzT�H��:��ƭ�4k׍T���Ā���W2��Y�a�=��m����z(DIS��_��H���vz������&0��&<1�|V�,��-�TP�N��F��OSTc���U�ԨW~��(���j:���wt�G��6���0F�ZzqL�m�Z��[�h�@�>�T;��W����1BS�c�g�wj� P���´U���|j7I�ig������R��<&�|Պ���ϙ�1���k�F�!셏��zx�����}��M;i����*�O�*p�{�u+�9���8���
�Vs��T�;"�fdΑn�j���|�;�:s�Dh��U|{�㸉?{�Gu�aD	N�OX�ԝӇw�	�u_h�E��?��wMT��w �P4�n����uz��ll���%*@��T��D�ҩHҁB�ʞ���O���E��D�����n�R'U�����_N  ����uf�����A�^�	q����j�@�uϋ#6��>��4ˬb�om�b��Cȷ�u�@?z5���-��6Y�j�n�k0Tŗ��;����]���&bK
�L�<�S"�TSm+�`J�ɁUySٹ"�[	�%%et52�#н�$��zy��k;�\�O~��zR�MݩU�e�e
2m��<3�P�t��N6K׋�j�{h�2�R��ɻ&�`?oEŀ��:���T������8�"�Ը�vr
�5��k�i�6�g7�N�"�J �������c"��R���ͩx��]�B��=�PK��k�������|��`�~�=B'�@��w�տ�e�f^�R&z5��KR�S�M|��q��y(��P��-��Z��y�6�����?t�u�i�	�bz�u��T�4�B_�N�"0́N��
)Ύ�vW�W���k`��.Ɓ���L��-�z1�/o��[ �R'���v/����zc�66y ����c���jhz��Gw5�]���7�c~yG�{tE��7��ǒ�����zM�&m��=aE����0 ip#�y�9T�Ue��GRy��I���:ͺ�8E���;Ub��u	$s76�eWe�.x��;|'\�nD�T���c����sRUf��iK��������y��>}��J�(̪� �B�(P4�� z����WN��/K�R0�W���v2bw!�Ħ�����>H�f��ҘP��0+�bp+�펤oq�Aq��� �t��=,��g�����}N�|��]�'���GC�6ǘƴ4��-��C��v�@v���n]uEw_��inU� (w��Pμ��f�*m8zn�=s˾��;�d��8�%AO��'�)��+[��wrL�d�g���e�QM>Wf��5�f�SC���]Bz�}T��:� SLi�b��Ev6�ø`��S�j�m�^�3^��0��eM�k�J��j�m�����Te'�Vm���������$�u�6�t��0{���k��>��&�W�D�6_���o�mk_4�6���xƶ�l�7kQ�xe�p�ay���)�(m�m;��X=A4ǳd)��M|���%�X<� -�8�����u?5L��h%9�mj{b��^�����-��
�m!Ę�R���z�9�Ĝ����^��\N,�@����c���j�re��{,>0��<��>�f�*/,�U����� Փ[�GVlҶ�䨵����u�u)��[C�O����#a��]xy��������wc�X�i���H�*w:kMF7Z�NN�"+4k9�d5����ڶ���=wZk�|�y���iM�?y���}O�MD������D+���9k��tv(s\�Sw*ln��5M�j.���K;���ܝ|�� �%% �
�Ei�@�i�ZA�篝��{�o=_k���Z��j<f��s��=���)]�8���0HSk����1پK|�;�\��s���V�B�"K�qb��C�e�iOa#%���+g��MU<+cq֏~�t�8��{��N�	��m*��^ސ��KG:/B���F]ʋg�OD�'>Y���me)���곮��l̨oՕ���8�VH��@���_D/�Ǝ����
�B��J��>���kuc�UU�\�+�1�~.���;�͡��w�l�RZ��9��bM,���u��tѷ\{��@¾���Oc���L9�,y؏��(���ih_�E�w˥E�2E�=��͞U��2ϛ�>�į��3~�.�L�Xi ����l'�9��K8��i;*��ko{:Μk�+�{n`P��x���i�Dc�9�2#��1�AWN�<����ك8C@�3�uRI��]^�x,q���*l����n������PC&�r�-� ��Um�7��WHI�wCL�<6K�>�=p%"���\���|��S	ĥk�΄7��oO�Ҍy���{]��Ъ��W��M�AS��z�N��HP0��_�7|�=�!Z�u}�ř��䝖0cհR����$ʧ��
[�J���Kmg�$�JȔ5�S�խ�&�Y1�[u��)ʻ�ǋFݩ�����*��b"��bE5m�ep�1}�> ��x3xxo{�.�r��m�]��x���1�6ڹ�y�T?:w������H�

yͩv�W�]\ə���P����O��e�xb����(^�V닽Q�aW�캚-���5C��[U�i��w�O}��uL�)�Lb#����2Vz;J�$�f�j������u���܁�\����oud�'��L��	zU����1��{�M?C��QL��(�����b�k���(s��sJ�߰�J+X�"'�4Bx�i閽K��w=yO6L��_L(R����ꤲ9��<��ǯ��cU3qU�aa��T�Q�0b���� [��4��~�F�ხ8�\����v��Ѻ�Zq��`����W>���"~���a��\[^������"C���Ct@5��q�oCm�ۧޗB���qK�򹇯,��eI`��\�0!F}!�L�Rc.�xr��e}3�TQΎ����+�Z�)��Ԋ��{��߱�� g}����*D�@�<`=�V���+�]en���q������1e�f��8�p-����s3�͉v������_������k�WUʖ��Պ�;����H�ٵ�Dr���b��z���MP��5V���z���F��g0;O�H��9��n�T9[U��OD�$^�)5��b�Ad�"wT�A�{i
D����N[i<��Ι�o�������J������C�K���#�H�³�z��� NCغ��|�C�f*��O>�F-Wc��[��0����D{a�H��8\P��ew�z- y7r��9{�\�y�+���T�����wP�H@r�`�vm����?�����f}���;�e���ۺر�g&�V�=�f�C�!sd:�6� E��Չ~�dO�4s�3�
�����K�jXFD�;4��YXq=[�nZUScX��%��ؕH�r5kH�����
��"k�5��|��u�T{U�aK��[�6'���[z�n�d�f$��Y�f��wB�d�>�|�Dj{x/�����k4�`��f�2w�֑u��=kd1%�wL�\��.~:�۪�V0l���g��:ɼW� �n�*���a�� ��M�l���r/�C�j��bc����M�ٺS=d���5V�꙯.k\�s�ɜ�Ư���J�ml����l�d>�\w�z9�
�M�W-���m����Ec�.�]�~��s��'�y��z��|�]������<�����x��sn�l<&]�SB�^ƉxqR�I=��ؼ9E�l
d��e}0=��7}+fo�!HJ�b��*�T�u�X,lo�4�pl'*yr���y0���4+NL��+[x����e���6Վ�=�;MI���a�:n�2��V	�	x�voI���ђm$P�uZ��hc>�&AќsR��b��DG�|������p7�[���׌�V���������_�m���*���PK����s�O�� �w�#|�(3�qU�x�w��j�˾m��W�Z6Z���P�[/��c�6pJ9�lg�(,���@fޗ���Q�x✼�������֡�/ç"�ʛ��%/W'ձ�n|�(�֟qk�cL�Ku�kl�e�5�&-* SC��G�v�������H���z&��߯`d�p�����ι//7'��|�G)[~���е�����'Y����?��yn#��~�*E̍nnSFo�_;�}N�f�/�Q?KK�{hh�I~^J�dX����&N0T��Y%�	q�E�v�;����^�%Uk�vf�Ӕ��^g�}�H"ASi��˯4�I��M����,��+�u,���)�ҷ�D$+�(���6&�F� ݏFz*J���iU���WP����W�<�Fyr�m4[���������4��p�6����PV��ߜ�a�����̞���/VӰ��."5�}���U�*����W�*w�t!�]��O�%����.jGR����Ѓ&�^ıe��̕?���H��n�\c�\�(�x�(M��LY�ZV/����څ{�O'a�d��n�*+X��k�Ʌܛ�%Z���)�@x^��O���z�rj��^cd��vpмp�c��R\�����ۙ���Ɂ��Wd�̮��x{�𫉮.M�s��a����n�O��@er2����Jh�4�r;An���:�]�����>��;H��*E6�oM������N�#�4�5�BR͵���Q�q��I�kTT�ɋk�u��:�(���U���kQ8�[Ok��t5�J�|�����nwk�Z��z���Gj5��5N����t��TW�����H<�֖����������n5-���ľVh��Xئ�%�2i��昮�v�o)��nW9cܺ>��G�p����wmjŒ��ݵEav߂��*'��}�|��.	�<����SҜ��/9�o�^��(��mN�犛���>I��,/�H�?>�$^Zy��M�u%�_�k:}#[�1]�Ӛ����N��`�=��)��>�K)n"N��'������M���xg��dtӗ�������������-�X`{�I������A��H�`��Y�y�zC�sӗ�/Lh,�[�{�:�BU�OaN�,�.�L�Ff��1��Ti�F��F��_/��ޤ�LE'���J��e}��v0�9�V��Sq���U'����V�>7d�#4n��-�(_�⩢�Ω��Ox�ꔟ�^�B����w+��
��&�`�R���������C�w3��� 𭼀EQn R�҅F��y(:��f����xx��܃Gp�n���p�������q�n��.��5��U�j1О���M-����a�Z��^!\�=����,����2�cu���ϙ�됌f��ᜌ����Kx�u�u���<�bDtS��s섞1Ϛ� ̀s[�3��681��V�Pn�*�$�͋odKNN����/��s�P��.��}�*ETE���lqQ��s���O�t�O/՘Sw�&�`��A�1r�o)��1d�<���>6P����<�O���ZK���c�v��쬊8ǡ൷k�u�QI���m��
w\UYP�E�;#^h�摧&��XZ,o'�N�ʇ<nD{�
f�ٕ9�x�~&�v.U�{hV�Ҿ���ke�]�E�AY�r��nZچ���.�.��k.�uI��&Ju�mSl���
�g���T�[s0�BP�����[��X���ʨ���'F
�7=>c,tKc1�<�A�a�����nO�jT��XŚ��[�"Q�m�'�1��d�u�#)�b,*�$.�z]��6i�u�3��#�?���+1/{��G�Y�(����q�m69��l��&�J��ze��c�`E>w�9�Ci-	젛���T��}��hG�^���ꐓ�5��
r��j�1;-=���@����ZS�0����R�{mf
�;����d-�$�p4�����"#�k{��f��0�#%��3�$-��֡Ϯ��1�YF7W�#_��[�S���0����R;f詈Yǲh�N�+8�P�zy:��q|��i��`�Aމ�4?���E/�yg�|���Yݫ*x��!��׵QLf�z{�+�I��Y�tU6����]�qg���NR/-QVv*�.7ӭv��5�a"��q-�rT�6���-tL�F��-^sb]�똀��6CR�ȼ�E���L���&��~��TG�H�XVz�Z��_�����01���<[�H�B�1:�뷧':کk b��%�]TG�b�*p��	>��O[p��}��3U���z�m���U�z�aC,X�9�B=6����Bz�L>��-�����������ٝ�yVs�N��B\Փ��F[p�����!�y	��� �ʘt��S�$w��#���Y�.�.a�ZIT�tzs�Y;qGݻ&JBDҐY%R&�=�X	�5P��G= fggd�[{} \����q��'U��\+|���E�׹�t)��P��ʭ�x��zJ��D��0�y�������O�Ƿ�����������������������y�{�]P�q�f�]�K�7u��4_�FX2�X��pg|m�\���`���o���D�`�b��I���5�'O�f��x�g��j�bWO
m��Ei�N��7$��ު˥�r�L�%r�e�\q81��;x�].��9�Żx՚ˏ�N)�{�]�g�ÿ��Ñ,p�9���hSo'�k,���:l1�X�I���W�K0��n��&�paɆ�(g:Nc}����xՍy�lD�HJ�T�����i���9�bT�@��9w�F��"s�t�7�Z���vj�y~�c7������ʝ�\���8+6�a�2e��d��3�1�����v��U1<]�2��w^��Ig���{�$W��tW,^P9����Ӂ���2i���njΧ�FNC%�y6�vJ:X���x\m��ڎ*tٕ|�5Wv&>ڭ몘�>0<:o�:)�wz��4p@�q�\�se8��$V�Ӂ0����H.�0�q�n��8*��2&�SZm����hA%m,w�`f�����(�u�拏@
�RW:�ɴ�̆a��Iՙ&�p:���?\;^݂�L�z��#��ݘe�<Z)�J^��Yq�"�Gx⳹�{���ϴ#'�ܮ�/0=xfV��]A41a7;�'�klV�5����͡Y�2�磷��9���6v��r��U���R��D9',���˫Ŕ�>&P�(	1�W��7��sVi;UhA�6Hp�E*����
�oK�ԇƜ���f�TT�Ӊ3qS�6N
�yLCu��m���w�����x��jYYۜu��qp��PS��;��7.W
5G7k�=��ګ��6�\,<�n-�+{�XƆQ9E�
��]k^7��6��ݵ6h�bd��gi(���s���:�������-I�<�(^GH_+/lϺ��C+P��A��6��@]+U��J�����7��M�6.�1n��ͮ�Y�$q�]�/s���;W��*k��Es_C��m���N�3ze�՝5��������ڡ�͕�+3;�y��p4���x��h�H��]U�	sw\��Xqj�T�S���Y��Η��/��r��������s#㮣Ы5Q��W�Czb�^܌���S���niH5	��q7�UԚ$Φ�V-��G^��`��s3�Wd�\㩬�c��7��C��9ر��m���6�I.���m�;����m����|�W8�6��=V.�qP�a;�78c�
����a�z.%iM˹���wq�fcc�f�����ݫ��������:�ݎ�ն䙓w��YQ�*�`}�
YNv�j�9�����E�P�Cʶޕ�w^�T�uU�8�:����E��]J{#W9{nx,��-�bo!b"t�]�fJ�dSc����p*��b��dfdf������I*٠q˅�X�E���c	���"p��I���%8ͫ[*��1$I�p�"*�� -��y#ZC��Z)�.y��:�5�OS�c�7$*�m�d�9���Q71��7�s��qW�/'��kTQ�棑�\ɺژ�kSAZ�֌F�ضDUi))�Eժ�����7*�14:��{�U��p�cr�1�W�5��mZ���F#lz��u���j4Ӡ��ճ��r���1�U���klm;�ʮZ�(�6�kf���cO#���É��h��s�1��l2aY�'��4�L�A�rU������W�u�^�z��Q��tk����b��kLrª�5Xڈ�[�]p�"$�OV�Umlj�&��;�.b�ָlb��f��������5�����9c���1����S��*���s��(�F�\�i:���E��ۑ���4ujne�ɪ�lhb���:���;s��Z�u�<*CI����3|�pӓu��64i��[�qꢋ�E%kA��r�l'6b}��Ap�"�"(���ljJ�=[�����-?#�Z*b*��`)}C��b٤����a�8z9���H���$�\e@X-�"D��S�ÙU^��@�*�n��v#y��X�)ʹǵY�S<
1��{�"�v�=�o	��\.�Ҡ�e�ͽ8�⸱��SXLq��R�3?@�!�D���T���O�% Ԓ���f'B'���������>��SM�J�k��I7p�����h�� 6���=�5R�����e28��{��=od�t�f}�53HVc+�C�B�u�N�4'�dΧ�$ЏO���gh=z-Q�����Y8;�mȖ�X��k��mx�Um�,���xֶӻ��53�R�S�u��=d�xY��TZS��Lnl/$x47=�G����o�g���)Z�М}�t
�g��D'֯�;��:I���'b�<h����{�6�&���3b,��Q�����Atct���:�xJϷ�7�eN��r���s1�
"1�ߪe�}}%����n9aEy(�屐��֨v�p͜r��4;R��<���=��/)�T����D�ꂟP]%�O���Ʒ�p�a�6o���j��ۢ�+�7��O����5��L'�yi/����k��1Zz:O>g��v=�eT͈t��U�ڽY�ݯ�H�C�V|k�P?�h������6N���@��BDyN�k���Z�u�P��w�&�X[E�{"eb��#9ޑ�+���z����qD����>���D/ߘ��>H�J�;@��"4�:<��Y�x��Q�W�6Rѐ�.>�TJY�; P{C.���=,uawqoY3���%0/�C�L�n��μ���z�[o������Eډ��Ҧ.�3sQ2��o X�w<����P�tKiJ�[��}G�(�|�">���Dg�aV��4��<]���$@�T�{�E�YP���ߚC�6�xdI��Z:��&}rm��t��r<�z򌓦�sXH�6�4�]D7�ک�?WP���N��t����#8�kK�왏F��j6n)Fk��yU�`�j�Kz��'�)Rf�T�:~^8&=q�u��f]����V�7�U[1+�������Q��w��������^��5Z�d�M�ñ�Gl^g)~����d�_���̴��v������7A@M�A�x6��e�5vKx�Y����T_u�	M�Y�"�RS��ڶ6o!�]4y��)��
�m����t1;"�]�˽�e�&R�
zU*q~�2��%j	�"�E����rr^�ǲ�����z�%�WB��;�8�}�=)����
���L��T�9�����"���
�[I�$,��82T-���:��9��?k�Ő�ŤU�S�g)ƠH���e�b`ƶi[�]�v3DrW������wL�4��
��.z�_�ԉ�Z�-[���;.SJ{	8�|�����'�k�o9Y�v��0f��K�)�"w*e�(��bi4��s!��P������
v2�4��r{{���Tծ�V�[>���}� �#E�Ӓ�d�ךFgr��s]���H��rMXf�U%���o��X�a^�[F2q�r:�,��m�V��)����U{����'�F�T/��SD��6;7���u�<M>b����\R����0���K�Z���e��r��9=�^F����8���jPyJf2"{åDX�z���]t��tR�ʿoK�*�Vgҽ�ל�841y��F׍Uk׸�������6@���ؠ���Q��S��j|�B�.��y)ܰc[#��w�g�m�/>c"��}4k�7YV�k`0����cEgmA��F[А鉡�N�Ƣ����)ʢ�qՒbo��Ҿ��5��<.M������x�D
��a+���� q��+�/��f}���X��N�}�)H�o.D�ML�W^�u�pcm��xH�>��P�S�Bп�����o�2"�w�5�䋫�5�c�{����Q�ͪ,��.V_�'}�'δR���W��H����}���ט˧Ԡ������n#��X�B9�J�;U19�Ǣ8pd���R}�%�+o�z����[1 ���>�
uH����M��՘�����Ϟo7���`tg��91�T�=>�ϵVp�r���*�qo�*n�c)��a��y���C}3B1{~�4Y�P���^��;Z�B���Tڜ;e��O&m�}ʕ��^��:U.��+�Տˋ���Lu)�]h�J�$�k'A�Fi�ջ�u7K�OI��Ԗ��7�t�Q��t=��D'^�0���5l�n��������n����#��Y�K�o�ճ���h��bղ%�W5�L���'�dbFI�Y�:��*Zo�ߦTŪ�k��
��e��0�|z�@�W�e�6ꃯ��%:��)�?`J}ٝ�|�jB�xV�"5�p��O#:��3"'�a7KЀ��z�{��=��9�#�2=��d�a^Ԧ)���4d!��")f�͚�m؃��&�)\���憘��z�Dcuz^uL�^�0y�`LJr-�ѱ�뷣7��o$�p�Y���2Y,g�O�������!��ȼ=E\`�������F7;5��݄s�zQ]B���q�w����|kJ	�ֹ}z�zC��h�3�D��y�v!k��E'&Ĉ���u���Sk�&��qV7<�3�i����ln/m�]�qUpiр�ʼ5Ѽmt�P+%i��G�����z_>��,w�8d��+�6�?A�����>ɟ�X����$N/�~��l�*#�i�^�֣��q��Ŗx��,�!f*�Ɏ�BY�T�.����Ϯ]��a�������I���{H�Y�d�������z̬��;7l�K�� b�Q/S���P�a���"��HR�2�	o-�xl��,55v��u�Kg���/�m�b�F�M���ڴ�4)\�/�g_p�L< ���W��\}�|6m ��[:�}������hu2z�S'��g�w`��X7���NV��z���\D���K��6���!�*V�&���
��qx7��H�}����U��Y{�q��6�U�C^�1����T!"r�V;��r��:a���ɹ��5e;і�-W�U�i�saK�j�O���lm�"SERmVX�J"�0�>;v2!�eㅍN�]�e�Ҿ��4��[�m C�/tdٯ��8����+d�xf�v)��h+2ő�=�w�]��V"�x�~���Wt'�e��KO�K1(���C���?�>"�}<�]ʕdL]�+��Ϛ��{��4�YX���\��5��j�@�	�>1G >�s��9*�'�9��Zۏ0w���z��>0A*�m�f�l�c��8�/@��S⬹��59���?/�<����@dL�:{�5��v���H��9�E>:�/̹������'���3ǌ�	��ۡ�Ar���7Sy���z�[�
%�0�on�"�@W'�PK��u#��.�n5��'�:�Q�_�a�b��~�'��\5�C�R�l&".�S-��-MB����u�[N�A���˶��������Ϛ/:�����f��r|�ؖn�$E���ϫ4i[
2�U���7��%�gZ�Ud�y4�݄ܢ{f*T
N�� u�h�'��=H����ۏݖ�R�cnl��.��rȕ�����,k�K��i¯]��PS���Ŷ�w������sz�'��O�x����O����t�/-���-��Rn���Aez��[o5xn����&��׭��~��t�9�S��T)�ށ@u��
�G�yWث�6`�}�e�T�6qJ#�GT��	��[��#�J�{�]+�����a�ks�1�a}펖�A���r��c'9�I4/��i�^n�*���4P����E�5�l�xf�e��dw�ǋ�S1B%ͥ�r������H���ڹl�C��>�[o���qo���9P����nZ�5�X/<W�T�I�;������s�h����r�|�32]�w�;APCf��Y�4���;(xlo��" e�Ą�����`���yu�"৩��]�5y� ��Pzi�D�	�_74��g�G0jc=�����G��U�IY>v�Ճ$߿2��)�}08����Ⱥ�k�A�l!��l�"r]�x��{*g˛mSrY8գT�L�@���p\M�D�~c��ǯGS��WC2��eZ���-7��0S�t_�~8�Smy)�{�T�l�fò�ן1<ѳ�4p����ǀ/(�`�ꭥ���H����[�������Ae�9-�׏9���U�3�FZ��"V�ӓ\(]X���1��x����ki��*���������'^wg�u�աԍ��޹N���n��ޭ��M�7��¥X�ьn��҄�ņ��}����|M�Hc�1�#`�sך�u*X�Qi�����Z�a�@��ǣ���i�4Lbz/�Vwk�^|v�*㙠_O3����,��*u�w J�/@Z[C�,�mZ�).��n�Y6�t�g��'�g�<W�*1���܈U;�8�=����Ę�����0k�y���8�����w�3�̶�/�B^S�)z��q~���z�M)�W`x�f(M�aQޤ��^S��
�v�\�A� �a����;�e��墕r�}/�q�Kʂ��܅�T���*KAz�W�nGp�r9P�[�$ � ���1ha�aq��P�������խx�׶WP�e8�K�[P9�6h�N���_K�K���rd�q�>��������b�\��||�d)a��]���nadt��<�7僔K}�d�O^E��)��y�n+�>�{��cLz!ÖKE��v¯�/��2o�g�o����ظ�\o3 �g�m�WP�Ά<���v&���}�P�L���~Xݣ3)7c�8�
�ͮ���4qF��e��ˋ�ۨc��͚qvN��m���9	�Nk{���6�d\���Cq�\�=W����&{N7��b' �S�c&7YSMi�x�<a�d��2p��VXYv�Y�!n�fR+P�.ҥljç@�n]��R<4�'ќ��X����wk/������3��}�WN�Wj�y�_����V�E|�5����/F�q�vj���񋹕��U�:�'���Cl?��"�B�o�S���*�������U������]Ii�=�V�����r�}��F�D0���5�P���R}���7��8�aM��bGT;"03�5IC8��W4��5�[Z�O ^Իw3���t�t>(��`b��
���&h��m[�z�K4D���5��q��eM�ד�P�-�4R�b���q]|��Rs�ϑ8�����k2��6(�0Aw�O)Ә�E���+a�~�>�o�Ae�5z�U~�)�x���.~�pf���;���s=����ю7D��r�`�ƟC��{�9���)���|�)��º݊��֯�Cݱ�O|3ێ}��I��J]����#�K��>תn/@c�>����Ȋ�y7]���*j����É��U�	0Y�3�%����X��)�0�<=Q�\Sh�x�(r.��{�#�����Q�i\���9�.6��t��댿#%��Z����3�������H���E�O�~��O:�m�t]����<g"w��v��w]opV���+7�}q7ڱ��k+a�笓:t�ld��Ý�h]�xy3z��\���q�dy�ә���I(��	�ywBmn���v,��W����[����-,&����S%��3G.���l���O��"+L�g��{;�:�
�B�Iƹ�H$��3s���1x�^[������XԠ��G�9�븋�&Q��B9{\d�׺o�`�(<����y��O�>��Ĳc
1�����adƵQ3Ͳ��/����S�οn�-~S��%cWG��|<<ă^yA����gݟ�M}͏j���5��F�I��)��轑�����x�S-~Ϲµz�k=0��o��[;�Ꙕ.qX'ޗ�����V�͔h7��xfPˌqw/~؂hq0JJ���t��뀎��x����aP�9�+h|6��v��ۉ��#m��MW�X��P�mBD�j�^Ç�YP�A�v�aRv��Ǫ�m�^�\M��i�ώ(��z�Z�TS�"�]���m֤&ԪD��Ɓ=�*!ߖ��%��z�Wfu�![�2�64�l�j����T���i�*��w)d��)�]~�X�׉p�իՓ}�a&���n��uC'@hxE��ƨsN�JAk`�ˑ�!N���{�Z���}҈|.U��1����aB��cM˶W�e�^��"a+�ξ�?���g��L@�>h&�{�(�0�+kE����]��׮eG�]���/�F�}�#|�<��>�a��$x�S�^9�Y�3Ԗ�e����G	����!KS��n����ys�=���dh_h�cQ��E��}��ë���(��l���*�qy��~��q�k��^��:�Q%�Z���:���]�=�O��E�j����DhuS�sȪrR����<�*9��]k�=q�\1�<������{����*V�5�&�pF(��{~���屶nc,��%ٓS�)�b�^���R[݄Ĉ%N�cކ�oc#u�]��_���T�Y����pA��t�� ����m�8��39���7T$�ܲ(-c ��Jt�\9��U8f�^x<t����y�M@K�kLgM5n�)�<�KFK���p�ζȅ7�1�sk�҇)��j�d]�a�li����_�*�#�<�?�<;�A���Ÿv��;�7[�zC����gH��jk���)��_�v�Ɉmx�,'����\�g����6[�i����ky�21�u�5��ܘ�0����U��D�kh�Rd� �~,��{��`=��.��0��;�g� �՟BW��;@�����l�"AT�p���O^�ﭗ,���I�zb�MN���=�fN�8����'Ӕ���z�~���R�1�U��x�=�O����������緷��������������������ֽ�[�pZά�9WN�.k�Ǭ#<��/I`��K�űk8^�?�V�I�3�Q�̾�ݩ:kqcӚR�B�{Kk������7,����L�&�i�v�3�1��^R�[^�2g+F�!j�hU�������[��zzb�E��Ii�d��;(_�*��k�P��ݧ"!qq2�e�74�3�m������VZ�6ЕҜ��A�d�p��l�뛣%�d�b�x�
�n��~u;:��7Iԃ�1ճ�n�vȧ�r�u,� &����Q߈�Y���6�fvخݽ"s2��B3o3�C���/�����7|������lqj�b Cq`Ǖ��S{ ����{y�8�L�,��,���+k��K˼�qՋ��U��z��6�
B��S����9��v���'B٫���{	��Y.�,q��A�c[XM�3jJ�iо�^��b�̡�9��w�"���;~S.hU�شg�<��X�&�xêf~�����h���|rX��gQz��ݛ8���"��7RV��d���{��|F�ոQܷ��Nc-�#h�+k����-���-w]��N���pY����x�����$�I�ۓmoon=�o�`��(b7+2��e���V kdR��IXr�v�H���=�\av��l���_S���Y���;_="�o`yl��Ņ�ϺK�D�i�0�Yt��!:J�݆N�2khA�V�v��eҥ�q
����8÷�:���R��C,+O��b�U����/�$��f�f����m��Э�sl����L���كVf��ə�V��S���㐎-�EС���UP�;�����O���o�#���u�)Ӑ��:�@{`�����>����̀�̛�i�y��|�Nɘ���qQ��0+,U�s�::���e-��G�7�mh�[�.$�S��q��j�z�r:�h�Q�a3O7���Н�M����mh�ݦ����¯ou�����mU����<Yv�R&�r� ���I#��_!��7�q�M콨�=�Tm9'7&)w�3ä.Z��b�r�,3V����e�˥໼�r�u��1
UܪF�Xɡr�B��0Ws�d�1���x�P��w�|���1*����^��{O�f7j�K�Ys��r��8��,9�ȶ�\
NF�[�r�����-�j��E�n9[s,h���`��4���U��Ռ��=bn�/f��ٙ�o
�ks�f�y��ٜ󌙙R�wh�#�후e+��i�ohڐ��'�ԋU�\�Ӵj呸��SYԄT�:���R�y��%A�:Hv��+u��wR§q���A7J.�=�ԭ���ON-e���L��RF���M&ڦSoZ�9����:�(#s�_oC�����A%DZUF��:�A�����sj��ƵU�գI81�X5O*�T�"bbh�:����bglr�Q��]>�jJ(b�E�^��'%��QQ͉�`��e��cl�cP�TDS[j&#��)��T�:��"
.Y�j�ZngE4r0T6��9�u��QY�\���f
A������LCQR���3�kQZ�5UC��[f����b���"
�Ij*`�x�O'MD����`�:)*�(��v(�#�����s��*�r��[m����AD�U�I�V�-͡���X��)��a(��s��AA�\�m�Z(��Z�!ETb���Ω"*���5�9Pp.W���~A�+��.�)�4�7%@Q�nm��s�
+cO�q%�R[D��*H�,F��A͂��C�,I���������
H�����A�Ӡыsr��"������H�)f))��_OoN}wy�{�u]���
�hl�Uч[%��{:92���o�G;��q�k��f���}��u�ʬ"b���?���υE�!�4�.>/SQ���6æ1*�^ߌ�y�T�2x�61}���Qeq�6z9�b�a��������pr����b�{�@<���	����煮cT;S�5�]�$73� qU�n��e���-w��bf�"�s�+7���tHՏ�~>T����y�����q�=$v�y��xz���~#�m��n�`Q�����G��5ʽ��b]�9[�@@�?exK�A��9�z�s�������Y~Y���Z��Sύ� ��73P��0Ҩɺ|O�	����ƟL(d�B�f�/���z�+-�w�M '��*�Z[C��JN\
ɪ��#l�e��y�1u�Csp��M"���os��Y�EՆQ��
6�4�mBr�)V�i������q�����Դ�v�A�=_\��O˽b�����CIӡY���͢*���.K!�sD{��e�ϡcE6k㻶�F��:�a"q}�gx�����<��>we�S0D��0�[<О�͟E�<�v��#�8���Ƈ�?����|�_Lu���>{|v�+�\ɫp:��QTj�8r�j�R�Ͱ����.����Q��O�O�h��S
��b$�yt�剙e-�mc��i�eh��`B׊6�*��,D����u�Qx';�3��Z0�5A7��T��MD�a]lkQbf[M��(�I6�D���e�.Y$�®#�zNΈ�m�)� ���ֱ�=�ꕦ�y�/ʼ�<ZD��R�3�en�3����>D	�l�D��(5���c��`���/n��0�E��⸓�|2��C{��&�v�G�EC���^�(:b�d�cl��ק���}�s&'~�����t��u�nM�l�-e�m��.��<	ok6(~�:�Du��6�}�iS�A����ڈ��H2�M]�3:=�3y�	���״=]mQ"u�=�	>��8��pKR�1H���]�eݒ�����$}H1��3��ZJ�-��S��Po���S��P.�9�rT�5������=�[[|�����
so��C(z���W"sG*��1d�<��v]A�2%M�oj>��7]�Gc���^�Z�#9�\Ʊ������	�{ĩ�5[���[c:��}�3l�C���M&s��SUv�ofm0l.���q���8�[�h�8ųfz�ޘI�ҟ"qP�u1�XMDB���J�����n^ml�}w��/�B\�� ��f4�'�� �=>]�ۥ�=_Y��pζ��v��}Bʧ�#��懕s�	�P��[����U�͞<B,v'[hmi��I!�Y�x���-�$��:bJ+5>��f{wP�D.i�j��alࢹWo���y�T���]k�i�blܷ�l��<��귭B귻�2~� �uB�	D/���Wޠ/��:�w�Ϲ	�6�Ϛ�jg� 9�#КE�P��̔>��+S�p�P�U<ܟ sR��˧���Z�(��\���M��4��#���ޕ���IZrn{w`��ێe6��l��\h&�s#%��3�$-�mj��y�3d�u7ʔ���ZI*'h��؏EUo��T{��Ъ��fX͍OIGs�����ٚh�<��:ҫ�������u��H0A�X36:׿L��ye"2y�#ucR3��<�j�YмX��M�U5�:K"t	�,/ߠP��BM���Ӑ���\@�#�9�c���.�6�F��=�h�S��gX�e^�ڝٵ�(c"}^��>0�r�m�5N�XU���NT��sKm����vL��Q|��ΘY9�z�Ƽ���L�]A�����8'�#,�x/�Q*�\,�Iq�D,��xQl�c��vnl<D�%)��%�8�A	�''i�fL����q8{&˟W#���o@SQ��c*�!��דM�{k��\�T �C������9\���v���o��C��'�x`@��?۔MȜ�|*��ST{����ZoT2"!��S�Y^~�{����q\�V���͘Ja��Tֳ��Y�k^�$A[
nn�2e��o�q	��`��We�Y�����r�Å×U	: ��5h����e�U⒩�ҩ�������v���w�N��0@��V�H���E�w��?M��?	�Rm#u�k��Z�5��7�W��L���W���Ar�ڳ��%f�=,��`qk�s].�x��<҉n��6�%��Z���� @@��?�~͋�Jǲ+.�Y�iY�e���+��~.�l��x����/CD��ԍ�]�̱ۤ�@b3m�N0���`U�>�d�w8ԻeLۯC�DA����Pvf�Uz�ky�/,U�=)E۞��Sw`K�x�^����c!�h�"-�&�`�
�wq�|�ͤ��d�@V�n1��!��E�]:�/���iPq������6뚄�K��$	�&�$��*P��� �g��b�o����QB	S�ϝG2�̄�Dw�ː
����=�y�ߚ��#��*q���̬�G��uЩ���KO�WT7c�
}m�gX"���)����wF�UJ�T�*0���"aG�ycӑb�X��%/W�ٵ5�υ�y7���YG:��sN�>f�]8ܚ���.���D@Ƈސ��"�﮽�����*���>���NP�L��/
u�=F�> Um	 ��w�,��>������'������f#i\�j���[�Luw�}3�W/�zB5Mʕ�/����2��*1�+��d��A���j1��Vv�Q��L5����.(���Jq�D�I��5uWrn�c�9c��b}m^;�z��#z���3k�ס�~l�Cj05�R�;/�U#�f���~��n�̷��.dck{.�OP�z�2w��ÇD;i��l2_d��j闔��}�5�e�m[P��fþ������x��0ISi����P̜�|�[�7`)w�A���c�H�	�&-����>���v�&Y���Ƹ�0�7�J����>\v��۫�~���YLg�L�p*'^_}�-��蚏T�S��}[���'|k��HԩE���K�mJ�ju�TN=Ȉ�*m�W��e���Ur���o���7#-�m(����^��0rc��Ғ���L�K*��+hUS���9�y������X��r;��>����f�-�'�	b�� �x�~�L��(��x�SiQv�Td8��v]A��"�KT�N�5ҽ����a���a)v�-�4]�@��]N/�J簔&&����Z�a���lY�a>[3W��^�6F�9�=��!�Ν��?3h���u*�?@)E�����T9��oW���������`�N��Y�9 �F����1��E<���
��E-��7�{9�;����_�v��jc5.�bn�āDn�	+�eSb�>�n-g�́�Y���x�ؖ���[��ۍcJ�ֈH�	9��:&.0E�5.�3��[��	�y��+��J�����D����P��	rG���M_u;P�R$R��ێ1� ��EIX�a�%f�~�/hp-��X�q���[K����x\�ɟϔ�`�EH�^xB�u�8ʯy�M���Ő�d�X�}cE6V�;�G����Q�&o<4E͊��fZ���uggM�1�@��U�{��͎nN�cԌi��Ƭ��Ў-�7����C���}�}ӎ������C
���j���S���A��.�{3|6�I�10>����^�004��{�]q�a�<ˀ��p,���_>ed	-����n �)�����G�f��ݥ���~�lm;��=�=��v`������}l�=+s��]秨�_;�:����<����B��Ȑ��k�n��_g:I�X'<��Y���(:jy��Ỷ%f��V��NϳՌjI��XY�BfנH�f����׊���6����o�,^���в�P��w��W���[����kR��UCе^�c/`�A��@��T��)�q=�0}0��kI�[x�~5;�����W�r��s�ҕ�	�t2�E�l����@� �=ȭF5������&�f�(ZW1���}o13��Pe���s;�[�S�5Ҳ���t�޸�@&S�K��l�6���Xϴ�6-�x��TZ�Y�%��J�B�ؐ;��:w�{�$��\����2�N�]1�E����'��ڬgA��:l�%t+�V��ṓ����/k"gD�M�+O���2��?c�C��T:yɁӽ��;�2/��<{{ئ��*s\�U�yb��R�R�ݝ���J!�ǵ�W��;Y�nfJ�[�b:E�L���H�$ՅJ^��=eu���۪Ciѻ��q����%��p �/�^�S�j:$��Q3Iz��,�@�b�G�ko*�빕�伷k��S�R9cnL�LW�2n�*�����������V<���/���B�٪A�CyRa@���>:�-�*,S�p����l�پvw~�M�f���_�3-U�D�5���t1�с��L��	�\�¤h�L�ÀY���H?3Y	y��[�.zUC����g�	�L�������hU*�8�3f���/�R[<�࡮__.����ډ��]?Y#4d��Z������K����cK���nr��^ԕ����rE��x߽nr���}�N[�Mϣ���U�"z&4�z>_�|V��(�i��66I�y��/)֥��C��8�bbqÇ�̍�k�-�m3������,���R�k ͙�uY+�ڵ���9Yn����*���إ��Y�����
�������<fn��}y���Yl{��سZoF���>�L�/�-�h�4<Cz�]%;
i�h�T��)�8�E�t�O��N��������Ju�\���M�v��@v�����Y!��K�|a>�h�E
1�˩׽���6�����2�3ᭁ�|`s4�5�e�v�������������z�q�&�F<�����[Vo�0|4y	��dؙ�S�=���\D�E%8��4ѯC�� T��Q#<��;y��rʌ�ޘ�D=��y��0�X�
7wn���yA�����m�<���0jl�*`a�t<�m���Bӷ%�l�~ji�\$�Ún���aUL(^�)��Rm��c���P�Y�K���������6�o���N8�͵%�|8`fisb}l�E�w)d+��>���*���S�d��Q=�/Fm����fJ�?k�+Ё���!TK/Y����jBh��;1��1u)�8UN�P^�N��=�,�L�=�U2/x��R��
�7Q�����]�'hG��7X4�;�[�{����2�Ǯ��]O~��R��<�[uz��m9�^.-�Y���ٍs`��EaY�XD'`��p9���>R��T�{}3e��?7�[})H��#U6Ol��<�|iw��]ՙ�IN;�
Ï�r�r��*������_C�0�)�jk��A�*���U}�k'r�UбNbm�]����&�鼵��<]=W�׏���Z��R�4lNM<(�ݐ��$�Ь����������$����vp�>?x�O�!>4m|��cB-U��y<��J�.����K`k9���5u�����r}�1��W���O�I~;ѳ��A/�!#�'QӒVh�˚z��R͹��o����Q�a�6
��?ϼ�"��zy��h.��| �Q���]X�;OeN�-h��<Y^v��jZBF�3�����z�_��.9�=���T;�L�m�4���G�+�m׭~^�t/O��^���S��޸Z�K16xG0�(3��vx�/v�o��
FAOX��{M��F�5��aw��6�͗�7`� ��κ���ʮ�����r��l�[���_���N��P���b�ٶ���~��r���p sm�H� �X���xex�|�w<��6h>��דO�W>T6�>�����7{ԍ~~eN��D�)��^l�􊪸��X[.\�.ڏ�9��UlQV��q}2���O��;2�$g'�۬ҭ����k�*K6�b[(YN�}�."'���{h��*�5�K��?���
DBQC\���S���0d���T6(F�}��i�t�Kg��,��k��K(�ƅƍ�0J��VԂ�N9ӢVGq�NPr��r����ߧ&��*��KD�bִ9}�&�w��C�y��q;���%\���2en�CXjV�<�u(p��fζ�����j7�7�e]�iC��+^��I��j%�m����["dZ�����`w��crL��\�=�ԕ��̪]����Y����L���Siθ�� �X�2�,ʵ��r],��E�;r�螥[��L=�yyxdE�5	K4�~���
�S\����\�&%�+f�[iCm��:T�l��x�T��͏TY���?���j�xo�Ӎ�y(b��>d��\]��v��)��4�O\���{(�a�ⷚ#O���r�dO�b1�z��'[3K������{�]���2;�����0���-��� �l��yb��}c���ͱj�z&����k�rV�İ����&�LZ�>4Z�yk���<>0�B����J)�r�;�E�(ټ#�̽�r�-)��%�p;=���lz��s/Z�}g��v���v裐���-����!�>��C�4c�y�\�X%�8�.��s�(���1��s�0�'�'��n8ң�>	�o�'�1a�ֺ���zv����gv�x��w&��O�������{|}=�����������=�����====>>3M.i��bN�)�i����!���%`�k�0ēf1Y[����:q��6�N�r��*J8A�+u:�]�[�ax��"��D*���3�-�o��{�᭨5ּ���*Ѻ��mF�&�JJcdw�n�fs�w�.�-���n��jX��|s��_'W��;��ܔr�ǘ�ō:��!Q� ��ڛ]���B�w"b��b��ؘ\�$u�&n��b[��51�q�B�X5-��X�t�@�.T�'g�G7P3n6,l�P�d��`t��[Yew(��	s����8�wzKkh��#6囕���&�
!��q��Ȼ/fts�Q��{s���꤆OFˠ��ie�����*��қv�\k�2��U�(Y)^�Dj�|H������&U�hS���1RnX�aA) )���7��ky�ʉ:o[�_UD�è��euc�˹A�DD����:��oY�4�5�P�g�J�3D�d��NJyj�	-�'k�k^ѧ�]漾��b�)6y1i^�>Tƻq{�٪���w(n���*"��=���4���)��o�u͵�.��;I����	�nu�����V(0��{}Y�c;���DJ��8F�xv��M�5W�����F�l��뽥z^�m���Zǆ\��k����f�u��}7
ߥ��Ծ�s��`�2�aW��l(8��a��<*�����ZN0�y@���qY9UE�����3�ӫ�;�7Mmmu�)��q���f�{�׋r$<�z���uV�0�G<2e���l�K7F�F⓼��ō91b}�s�;���7/a�9���.�5\��4�ٮ,s�d���93�݄vbs��1	ײ�d��;�陌��	��v�'SeWk;g30Z�m�+Dzs
�#�+��1d������W:²�(\�3i��gCHo<��THFry��lcJ��E�.�E����=�n��l��/zN�V(��MD�B,�Ee�Lfbٛn�)�\������6������1�F�Jѥ)��+׼�j��&O�։qn�e,�2���s����$8@���mf��.�٥�r��*�Û��q/3��PV����#uj8*72�<-���ug=[޾���J��zI����GdТ�3�aNx�*�*t�=�Y�\�?�"f����=ZsL������7��.����*KH0�&S�.�hI�N𧜽�9ڦr����wʱ���nB�ǃj���0Ri���Z�Ӑ��}�ek��5���nث���u��V;�uάW6w�l���c[�GyXe��'I�./c#s6�e�n�1v�/�ٙ27��ؼ
��'�����8�k�]L`�447MF�6�墸l8n����Ѓ�Syi����ڗ���^Crf���M�/.1����t��G�7�j��nM��[�e�REV��e��ΎT�A�m��&�"�J
�I����ִ4m`+��R�]QM�b4i��t��TQ�sm��f��֌h��<��QI7$ЕI2[j�*6]@lo\�r�h�U5[��F�UIK1�K�1-s����j4�S0PQE1���f((JV�����M!PQKP��E� )���h�5�Z�h"J)q�K�Th�MQ�9m%hv�6*�9	�mi5mC�ͳ�������y�q46�Bj�4PQUMm��9\7-z�G:�"+���IE#AAEU��"$������h5K��j���h(��mC�MSAMՃ�k@b(��q�剋IF���������EAS5�U\�(���B�F�h�"(4�詪�ađ&�$E4�MP�U�py'LM�Z�mMTW,P��HQKE?6�y�R����>����J�BJ�EI���FHO�	��_�g��c���<�Hl5f���{8gIyJJћl�Nx��5�#�.�WDT��ó�m�����k��R6���	�K�D�-6�1�H�,3�|cr(Z8B
H  �Q?���œ�Z7}��⺥·\[��N�4s�!�Ԇ���M��_�LMy�_���^P�-|}S/�K�o:�{2�L�Օ��������G�{=�Z�b1�=x���PLik=�~�Dq�������~���`����y}2X�"=�̡���4���y����6�Խs��P�[Ew
��M�W��Oe��1��p�5�yA�@���8��9MÉ��4G�.b!��Dmd��5���ک@Df�
�O4�m�0���eW�Kr�y���5g-����6艛X�{�����L�������^PS�eH���J�;6��O�4����m�[�
BY��ۮ@�ӆ��b�q��v���yǃ�z���a�3�Ś�&�c��=S��P�>�w+� �:�O�^� ;[{��}��dk'!���UI"��/� |׬!�=)����T��heد7��d��s� '�4��e�R�oR9clI�Ɋ�O/m"2ש~��*�8x�����sj�3�vU�2�E>7��3	�{�{]s�o%+\Tj���ظy������&DCVH#3_�3f
�� �����t�Vgu�|��<j�M2Vqs�b��O,+��aݻ!!�y�R�|s��\Lp��z��'2�[�f)$��r�N��S{��qd7�旨9죛v���p�f�wAIow1)�;b�L��NM�5�R�=�� =���xK~�?�&1�y/"ɑ=�L��mW0���K<2_0MM;/�Ϛ53t.Qy�1��/q��d�	���'����h��V?2�(ٯJ�	Gc��{���k�o��N�1ky�`*f��K�"{�~�%?"A;Aw�k�&Y�;�oJ�cR�����/7�B���X�V���/��2T�6k�p���*�d<��	�־�sL�aF38�3�OE��od̚�_�Fy�\���M�v��@f��!�]�0+��J{`�re�E�>��f�`��~�w�NGUA�c�']�a0w��Z�S+Po���B��-s�s��*$�Ksf��Qj���"2lM�^�oS����/�����?^�xc�l.�����o���_H~�߁��@��0����ANY�
i�XÔ��03�]M��xW#N�q
m�ƃ�o����?�2?dh��k(�6�2=K�j�]ͷPJe�֑)��HM�ԛ��ި�s:�6��������v�����4*^Ί��D�<L#�(�A�qˉ�2�Sl�y��0t�8��a�56�me����0wayl�$.��]9��{���:���*��wm�i��H颽��]:����v%I���@y��m���۴�}��분���A��9���E�{1��}��q����kٱ����>���O�q5�s�����\�ٳ�]�$`�����g�62 $X�����(	��A<FXj�UT�i&�z�
�3I���,�%T�>'��K+QQ�0(^C��w��T68�9�԰��KC�m��_���t-�4Y�o4��es�<L8%R��W�o:u��k�le���KV���|�mn�&�]��Bm\h���"��O'�1I���G7����b�9]�`���;o8�,��>�������o���U-���'�	U�p���𓳨K����>�iF�����w�ƾ�<���
���>"6��w*��7�����"����~h���GvB�PX���Ʃv��5h�q��κD��%�446�ֶ��-��KڌY��{vb��-��y�R��O��3�n#;~h.60�� |�yz{ֲO8�]�����ck�^����#[lDrW� ����;�_A�p����M"v�r��t6*/.R��W��8r|f=A���'=�|9H�̌mk6w����"Kو�������3㖋�u����6v�k�ne�	�������Y� �/ug�{���$ټ6�A̝U����G�D�4g
X��(�3������"���Tv����v:�Vz�N��`����wt��+�xd�6"Pnj9��\�^�je>�yE��t�q?���y��lh�+��%�*+*��mGga�n9�I�y���+ٌ��<l������n�s@) T�����	�W~����<��� �˿��u�����-M3-偡-�>q�^	-z^
���@�v��5�d�K�8TS�۬�)��_�.ꅛ�۵�Ⱥ�{��P�
�0�pL\?V�U���mʑT"�S\�Jd��@�jβOUf5k�i����v��}>v�S�kZ�SjY"tf��xmaJ#=��vW(��W?f����xX��S�T7B���Bd_�}�P���Q��T[CY5��?Vj���P�y�V�ԋkMMTH�C����ѳA�Dn�\_�M���.y�P���B��ČƉ�S�ur��2Փ��v=�� ���i���/d3n�<�� �V��I��ϓ;m�>SQ�H=�V���sO����'(COW�to���P���_|��o�h�_c���1Ә�<��s� 9T��G�.��k߽�)��'�XE�?3�u|B��Y7�z<���1�3S�iȗ�Ws�֪1�u�/��*O��i���(����%j�g4�!��/on�u	r<��i���*׵#�����x����l-0�[̧Q��9��e��k
AD�ѷ�vf�iٻ*7%�Jwpg-}A
��CMJ�s���ۼ���}�@�W�h���g����a�8�qD#j�p߅�2��b�]�)�_�2K���2.N��H���L����B��*9н؉8��1>��CCc��������5�*�܏u��46G�
���[@l�R<T�q<k��\.fA���-�˖��M�'�dOwIN7�C�������y6��>{N����"b\�?��2N��`lV�yG���4�=�	|��9�d�-�'�V�uU�E�����0��]���^k��;Dd_=!�)��5�N�b,Jxn�d�;)[Y��3K��^0��FF��KPJ\N4��<���5��m��4�XP��lO*-�n�$�����]��'-�9����AWA�ܦ��ty�D�μ��d,���,���;��{� �sc�c���ڏY͚��~e�B�)�CT���t�\�^�f�U᭿o1+������Uu�*]Kȫ��L-z}$2�,���]
7���2��=J8�]#9VwFLm4|�v�������Mx�N���k����;�2/cR�G7����K��4:qX�E�'�62
;u���o����T\�on�
�S�F���cj��&\;q��5���V�Q+kr`n޹�h�� �G�2mw�ƳK��y�b�&n�`N�EC����`�����;�J�ԁ�E��a��M��R�Q�^��q2�/r�����y���l�������qy�i�.��iف��
�������Ҿ�����>=�p���{Jd��]�bJ|Q�V/^�fP�Y9/m��Y��g)|�]'>7�#36�k���u__Y�4��k��&y1�i;�	]"������S����i�ǅ�a��Y�}'�Z�{�p���E��G���lek�q����dRb�9��n��D��W�NI�.^t;�O�$k ��O���twJ��"R�9�%k�RyJ��r�5y�k���̻����~]S��Ƚ�^�1I;��n�����+��[�lErs���u@0>����)�R�����L��tθjhܬ�\��@�ǂ8��g$iY�0c�Z�ؔ�}7)E͈Z�������wvkǹP]�#�>I��z�l�m2�����癔##�N�����-[�f�������i��8ٟ��Z3��^��y���KY��i�eT��<ڋ�,�E����mc�:�Jy2��j����I\T��&]M�p�^]!��V�Р���0g>8>E����,��+g5�mI���{C�6��2�jY���]k��$
���눴�P�֨���Ԗ�x�Y���mv�#��Q��[�~��{s7x����b9Ri�n�M�R;b��v�i����|�"Ａ)�7��$A�I��w���w��i�]�����*Cӳ!�����Ϲ��EW%���k�a���"��R���e&l*��z��k2�[-E��4{���Ԯ5Z��'hN%~�62j���W�<��zI��牵��*���-�K���\imO<c��5i�[�
���P/d7im��]j/7j�V>^2�~nX/}�Y�_�$��'�\�'y��4������yz�|6��%l�ΏÝfߡ��s�6����v�; N��恼���i%ܰ[��ʥp�B����3}C^4�)��hn�,���#���'�����~��++.��x6c�^p���ʉv��3�,�s����"Q��	��^N������
�h;�G���6rA��R.��슚�4�ʖ�v��lG�.^L�r����B%�s=aV������Y"޹)$	�k�@xK��g�3�)�V�V�$7���)A��92�Y��pjMC�.T���Ő7�=��*�k��������r9�����3����3ѝ�G|�>[�����7n��t��1����Yc�%ۉb�}��3���q�:�}�qܪNMC�T������ι s\���+�L�|�"�;=�/ms�[iW�y�9>޸��;p���{.	YՃ�+5�sw�,�K@�uO�3U��3tF�&f��C&�J�틨e%�9�خ��l����R���"%H��S��}S%�2��@�e�w=V2{�/�u h�
����`w��X���$��[sWvc�ٮ_��)>q�2¹����x
�h�*u����O|�&�-X!�e�R+rv����{[zd{GB)��\�\���KYj����X2Tv��m�9�г�yV�H%e6�We+�U�G�ɺ�F�hj=n�E+�.��e��p����tFye�䍨Y�ҭ��+<��?�`��Ym��C[�ۦf�T+��������C�_2�"J4�օ?j��6�
��]C�"t]>���.�KT}bݢGT���ӴZ��w,�Y/�ۍԮ�y]��-��\L��s)��ԯ9�q����`����;TeЉNb��K	���Ƶ�:�i��6�6����2icq}�9��۱- =7
w1��Z��٦���O���k~qy�h�pU}b�WMt%�Q��x*_[�N�q���>m$m�<wf@kq�5��p>�p}�l������ڗ`��f]�2�+ͪ�Z𶮼#��W@i�Z�C��#zn�v�f��6%�K4�EM/&�+wb6K}��ɘ������v�@l��2�v]=�q:[�ƌU�;	۷��j���zR�wWX~Ksl3`�4��l��V��
�z���������a��\��2�+ݽD���m�Ti���������"j��K��$�i{�b;��<Z���ؗę�t�u��n���e!��9�K�]"���\�3Ln`��z]���dۉ�0qm6KHs|0���ߣ/�%"Q���P���"�{<��=��q��״W��y�Î��d������l�Ąj�ީ��_��a�.4��ΫK�Յq��7�M]���=]�H�fk]�;�]j=��֭��+ٴ�IU��:����<+sz3X=Pz��5)��{5�[q�������zvp�];6��{^�}qN 8�DM�-��T,P
�/qH1;�x���飔E3����C��fql�K�qB�����u#Sj����/�'Bi|��[�SN��y14��ݘy�_W�1xm���,��J2����\�v`	�4C����}`w�4��өf��e���n!8:��s�.���o���h��UC%��4���ٰ��a���F�'����H���5=z��d�vY5�xٻ�e�mWꇸ�ؑvKCTO!ʎ�@,*"���9�^�H&;��H�흉U�9]Ċ�5-yɳ=	kU�LޔŶ�M>ָ��2�H� VG2}7�q.���`��H��{���Nn�6���Ӻw:�Vޝ`�qxAH�D�f�TM"�̤�yn��8�B�l3��y������g}!��;�tw� �H���+R]�'=�y�S�]�EM��&�K���ᕈ�e�>���u	�Fdo"���_�>�O�������{{{{{{{{~=�������������{�{�Ǘ\��?.e�^}d�9`��&R����-
y�0��t���" (��`�c7�6�.	-}��o]A����v
X��t��֢�f�nFV�@f�1p�D�t�����<�R+��'N��9�Q���pm^�a� �0q�Ǵ��$0�m��x�;�k͚h{��5���fҰ+�H�6"�|���-�����nA�[�ɻo�1=X�ir��i�	ͼl�8�U�q���][���P{T����-+,�]���|���D�j����w:�5�/`��.��}���x���r�7����w;+�e�Z�7,"�L0]�E[J]�h�Z��.�lST�@�{ʶ3����HNh�6	�t����˦L�U�Ȝ���d�l���ӎ�x��hWk(ݹS�����0�h��TDy]���+Vo+Y0r�ԕ=іw��6T���s3O0͠L��8�l��ã����,_M�l:n��7��F�.�X�=j�c����F�NU9KI�G������mF���n��a�-��]��@Ƴ��)����L�z)�-0{b}��U�+[��DNC�T��ˍ(`�T���S���,,̤:�1[4��aM�i�er���V
�ܗ�n�xb_��c�z��l��0��Z+[�!�W�e�p��}�qE ^r�~�~�IM��%:#�[��D}�;�P}}Zx��1�7;uȍ�����&�wj���6n�Oޝ�;%����QI�V���l4��t��̇�G[�b<����˳^��
���^t|��u�d�nxj�fE�y˝�ֻ��.<�t��%��[V�9����Rn�k����bފ�:��I�o��߲e�3��z�ͼG�l��M�C��C&��wǶhK%2p6��gIZ1�k/���DvE7:��ʻP�7w��x;tѬ$Hwj��Gu�e�^�.��)��o4GY@�꜋s�2g�N�s�xћ����ì��p��G)�LM�כk�����<�(n��v��.d��6�R-zO_H\*t�o��r�v'��f�&����tJB�n �\�×����|����Nց(��5��k*�en����`���.��F�^4	{�H'w!����3���Qڛ�[sB��{��n�@\�Zʁ�4,:�a���.D�mi{��%.gi�Ha��>9�|�Z��v�vZ����GZMF6깇�ؽk�ޣ�r�([��(>1e�u�4>���c�X��\�}*o��qT��@��ų��mo�ڋ��_t��+9�i�����1����}�:^�j0Vfv�n��/=9�_�I�;�*��:&%b��v3d	O7��l���bN��<7�E\S�,$N'�w�멵��.��YH�oh�rc��'r�<;h� T����++g6�KH�Hk��m�5��wl����J��2vCx�Kr3+-�ƚ	���wwf�.�]���e����U��m�)(����)j��@DX�h���JJR傶3PM$AH�T11UkSD
�������U���U� �A�D%)��Қ4UQV�IS&��*�����I����VH��k�&(��*���E1/%4��DO �SIm�������

)N�S��RQHU�Z�����*���*F�).j5�5u�<*�@���ph��0sᪧ�yp�
Z*��X�J"H�����1�J����塪j�+M�4V�\�r�W$�� 1�f��v1KG��V����Z4�4�h�{Ɩ咪�:夢�����N&�cT%	I:�!I@��QK�Ҕ��@��Ph��\"����JL-\#F�Ei�C��9�M%]�O��n��}[����~k�-2KxNn�N��J��c{��JmŴ�E"{���m;��ZV�F�`˴E50�����K�{�#@����G�|��oAT��~���^گTekz�r�uR�oO���j��B:�m��t��yd�`>ϡ��Ĝu�ڑw|'�دw��Rp+��;~]��&�{"A�=!��X�^qN�֔-�>b8�#�t$SB�Tj�����3L��N]�Խ�O�|]�'9�$!R���)���=Zvj:]�6y��x��b�Z�d��ø��/�#H��I�!�1=ٜ��uwTވ��.�=�QR!%16n�33)�4���Q�������s+7�?LX��f;��}�L���`=r���ϵB��R&��YJV���vh	��s��;
�5SW*��F^�r��{��\dt$w�+����=���9�i�{:��g��+2=U�R���UM�fj�S�A���q�M{��4sT7|⫳j�9WBF�Rv��9(ݪ0�&�-���4bE�͗���c����Ib�z����۩���Ng��TR���dU�0��o2����:	p.8�`�>��5�	�gl�d��󪠪�_l�=RfL�L����V
i̍:��� Ь�ÍQ���.���qc%��z��t'U�G[�x�L+{:��y����|X��̝���]Y�N#��%IR�~J�@�y���5:v����oꕗU!�8��kT_s@����c;i�L�0�xc�<�w�0E�D�	��x(oӽA�_`��w��s�!��f5g�+l����,�|�w��3�%�O�]��t�K��f�D.���J�r]�oQ�\
bg,:o:���M�����9-T:6V�eʞ�I	����uԞQ;Z��yo�$7[V4b�x��Y�v	�g��u��vbܟ�~;���n��{��;����3���F�=��P����ʐ��͋��g���k-��Gbx�u���-��`X{�2�ԟ_��� ut�9ޱ�`�=�۝�a�i%�����{z��e�X �%�ԁ�ؤ���x��كT�����G���H,f�k���(�mNi�u�L�v�`f�V:G��M�u���\�t�Q�4�v�`О�KEK+�P�]�ʳB2jH�zܸ8��7�ɼ�ՁǍ���V!Vis��yI���M ގ	a�t�yb���Ro����j"-s"�3�ޭ-~���֯����'��nR���.�*�0 k��4�����IV��ԍ�� 5���g-�M���i�{��כw�D3�Q�y�n^�_�(��������k3�=<Sl�!����=}��g��dU�nQ0���^�U�9�\�x��ۿn5���➿B�Ɏ�'�z�^��v�T6�J���ԭ���8Q�6T�m)�	Ѣ��+@����	��wٲTy?������T��ᐻ���	k�h��L�����ѩ�p��j�k�q[9�[B��
k>�r�8�ಐ���f����y�,Wr�2�l%�+��F��g�IlWB�|�*��Oj�Z�^�i�h�Zzʷ�}��<l1G��n�(�-�d܆Y�
B�����t�	m�g�F����S7��j[�l?(3�o;����1���ckb�JΓC��Ƒ�����J}����a��\���t�v��_���:�ȗ�(��L�wx��	E�h`���<�5.��d����9�L��e��"����ϰ�o2��M�)��p�H֐���[�O폝]H5���v�f2�\T��R4l���t�1�;W�ZaBh�{5B��Zv�TX���u[y�N�go���|��~�w%c�Ҭ�Vu���gj҄\��G��+�/�ݛ�-�^0 �N�/���ל]�^~�����2�YGZ��̦j���ݶ:�L�-!��:c�I�ѕ��=�x�ˍ�ak-W&M�����\@,�h'�Ty�BΆ��A����f���r�۱cr{f�?3�@Dݪ�`2=7w b-�.;��JP&Y]�gB�ig)���;-=8'��{�D�����i��p���л�W�e\�����sEm��_��GM|����ˋ�����C1��,�j��K���CU\3a�#g3{`��U��UC7�}�O�gy�*�T'�W����E�S:7���{���s^�֕櫩�6�E�.��ڻ��ϑ�xt�M�JW7�+zky���D;v�)clһ�Wq!����8E�3�������~���|m�f/�gr�r���"�Ȥ�{[�M�w��\��+RT:�ȇcVyo�;5��Vg�-�j��������}ru%;1���!�b�Bɉ���c��V���-�T�:i�:(NI[0�k����!�mb%������f���Y��\Y��(�h����~�d��%t�G4
n�GEU!�9�0-Ua~��2�ׄ:���o�&������(��Rv�[�#��:�t�T�.�D�Q9�vz��˗3S�p`09v���
F�� wRoj��%6����Ds5U�zbw��RmI�-����v�[�O�Qv4EL��u&�m�lg��,$akSl�3l�ᷚvޑ~�R"z�c��NNki�5����脼J��񜰄93u���Լu�qa�U[��V�no��em���C���Rc�n�diTN\�Kሣ�gKi�����ƽ��q"2�kAc�'8n��Go�67��<�ec��m��:�����8���zLa8��;B����S����n���G���,!�b9��ʾ{T�r����5�<�f�_ .�(37�o��>_|a�����H��=?d�,M�d합kWGz�(+�uݰ�z�t���(h����n^fD��F�	։t��;�nk���h�M��r^�b3~+a�g��/���F�M
�s��aN�О�f��rMk��Bq�g7n�?}��o+f�4�;-�@x�e0��Gt�ݒ˱cTy���+|��b�������`���7U�?���P��e�{������D��7�}�4���LG+��t;�R)Ga4���8��=Aly��^]���� YPcs;��)���ޮ�O����t�t����v���X�+�ϵ�S<��t�f�>�{>g�ن��m���b;@6�%iRbo.�L��Km<B[ڲ�dn�"�к�qh~$V�����%A�wlR�]n������|{��"t�L����Y�Y���w���� �%o-��ڌ��V�Jށ�yv�|�b��[�s}�<�`d����dJ5������[��)��B;����V_lU����sZ��¶���ٲ��.O5b�DH��қ�g�w�5C��Bd�F*ԫG^:������u�l�W���4�[0�W�ʕ���e���a�5�x���C��3������Q��#��~#��s���~먷��]�kgE��_U�q�Uc����ʋV�S�%!xb�$�u��o�Z�:c�e7��3�T�՝�*l-��MY����}��v,�괟���ɒ}�;o��̓+B��qw�Q}���G��tv-�97:�7ym�&��� ���(�
r]y��ʦ]�ٵ�R�z��,�фȀ����xl�y�x�݈�����5}���GE�N仙�g �����U`�j�n�*֍���s����r���{����p��U'��
1�x����r��Kx:^�V�-��PҚ�p�௕3/r�W���P+�[�Z��a�qe=tlt��c͘}��[������J.@�l�S�CQ�R={T���Ɏ������*a�)[o�Ҳ�P*��'i+���������l�V�,���*u�w�f�\���1
�����w@c��>��&��\H�{��&Fl�K�e�h���d.�QR�9>)g.�PoI��QۘI=�,�M[\�"Aݩku�����!{���y��.�nC�x��Z�1� #�Ht���>�U`uxgA4���Fg�[{+�q���^�?Y�	���WJ��ո�b�"o-�dc!h��]���so7_#���2T��\4��H�b���+��l7升�N=�2�%'�e�`ُ�vvq=�;3g��}�'F�H�R�o�����=S�9����B���:��4me��ڭ�;��憁J�שsV��\`4�Q������	��ޕ&�ʪ~u'�Ӹ�U�(gS�";M��[-��:�*
Wq8���Ƭ��ƅ�r툜4s"ȶb�թ��(������(�Rov�-�
A -l�,��H�X�NO�ǨJ��r�ڍxd���ۥcS17<Z32c.*�f����S o*~�����6�G��K�wW�,=��k����#����ݶ�>�=��-ؑ�=��;�0��d�e���ʬ54�Y����j�X�����K��Ѯn@\���R]�AůV�P��#�e���Ӎ�W�u��ocLA$����>����,AT j�Smu8TC�Z��٥bK�һ²���𫟞f%��]a/<����8��_��44�1�c5ݿE����J�po��N�a�`���˖�(�W����Y�hN��I���`+����Y��:���d��/��^4��坔�z�uG�v��u����OM����� �P�k��}Z�UZwN�"Q���g$��N��I5?��;ݾ5u�l��TO�6�<d����[a�f��(�46q	�n�4�s-e�B쵍f T;�S�R��<�x�=��`ډp�~T֮��Ո��i�hⅼ-^IWuB�:��]>k����I�wz��1#���n�T>z�T�ֹ9\QF�V�+�T�4�3�c���r�ź
㶗gv53	��#x͐��)����)gOn�] J��&�a�������^�y���ݢ4��y�.��N&�i����Ϝ���$��{y���l��
��z��I����xrf~�@n)y<�]OH����j����a��ٷ���%J����X�gP�w0��'Ǳ(O���\�3�]ٴW�Q��*�D��n]v�,�Ny3Ko�|y����#PudּZ%0�[�]m� ��/\7���{�\+��{�2}���������NҔ��L�����&��������]c\v��hT��=*�F'�ݸ�G�t7)�n���k�6v�!�w��s�#���.N���r�b1����B�&7"��*h&�8���];u��h�ݧ�	B��v�Í�J�i�jL��Vmk�X�}�")�����͟}�e\*~�d�����;rO>I���dim4ύ�9>N�U��}H|zn�uY��w�*�a�sjL&�7�n���TllM?f��5|1�k�t�Q ,0"=DR/�vcF�x��ل8�|$�+��=��~�x*��)\������+�!"&��󋻗�eJٸ��lWW�'�2evBH�$\b�h�N�j��F�x�N�E_����|��hڜl�ʺ7ɭ����"��~)f������;��j2�]���Q��T���ؚ�����|��
����b��4��km���10Yu5��w�k��-�ͅ<�»�,2�k�U�n*��������?~qvJ��Y��Wt�J{,�j�"�8-�1�����wR��O}�H����&�b�g��2z����������=}�y# X G���������������������=��������������]]���C�\�_l��$m�0��͠A�Lho���¯F(�{'Gŗo�M���%�!ٹ�:������-%�p�Vs]���L9����;���CX55�ԫ�T��0�|�v�ڙƕ�L%�h߶��ńv[�[]���(�Gv+��v��u�%ku����̭�y�����K��j�hj�A��.�ӗȨS�VyA�l�"ٵ�mJ�`2��XY\�a�E�"1'3c�����7o����Z�8����MC� M!Zn+}��j�d�m\�h�ݧ��z<�j���7�"l�d��PV��3u�1gf슬R+q:�����'CRэ��"��Z������V��������mB���䮙���t}B�w��,��y����q��#Zb�wv� �z�>�̲t�!��A�J-��)lL�\�qN�|���=I�L���a��H�2���d���*P)+�9Pږ����l˄���aЈ�2�o��v���ˤѼ��<��
�n�+b��<܃�
�5��ˊwg�Ɩm��7(k�㕵ֈ�4P'���)�Yj�twݼ62)�}������\5

���cӗY��of�vAI	zc��,e��e��ѻ�9����1��%�v���7���E,��&��	��m��*b2�a��T�bt��R6�������aڥ���s;�ӁRBi�n����r��C�:w.����U*�Ss}:���[R���Y2�<M��7�lw,`�39}�!�齲;,�O+}����\]X�eP�Kb���$Y��iP݅�n`�á�C���������K�<ﮔ�9Ӳc�R��e��U��ݼ����c���.��d�f^ڣ�N&��)T��7rro����_��W�Z�1�l�;G;_ʓ�.��'EG�W�^���1[F�9׻XZrM� 9��5y�󻗫�`���S�vR�8��E:g\���a©m�9ǲS��:��s�U�*hӛ���Ƈ�-䕠:�z�d��5vE��ζ6[0צI���Cj�fǶ���K�������	-��vֻ����6:�f��f�m�|<������.Wʝk306�Y%��mU�`'g&�f�K m5q�I�(�X-�X"�ɷ�!��Ãi�������v�VLvlk{@��N�uD���tVQ��4ݦL��Y�vy2�b�6�ދy�^M�j����3QpSӂe�Lk���v*��F�-o<�ヸ��*�W�wR˚�=�v�Z�b��U\e݅���4��%��î�"�AL5�Jb�ET�!�b�@�Ʉ!���ڪ{�a���Ci�U�K N�W<3Jؾ4�B����{ͻ�J�����_ݽ%�T0
�L}'�'^6s�˞��s9]ۇ�"�/�s���f�.��w_���xM4%	IT�D!AE%#��D�P�Z�ը�"�ű��
~X咄z�>�R�|x4R>�ESDAu�LA�F�p��)j��:bhh"Z�����"����\�lD���S�%4PUT�F�J|6*b�Q���-!@�JB�Jh��4i(�)"�"��F�Mb�h��*y*���(�:������{�8:*���Q5!R��L�S��t<�4�k����f��5hJ�bZ��Z��uIKlj&��M9���k��Zҝ�#��N�v��NlQ�G8��àiiV��{�F�Ŷj��񒹵& ��O]u�TD�u�rM-TUm�Ic�7���[b��A��AA$_wӜ���޹%��c�@��_DG$rD�1Ϗeᜒѩ�W���2i=�ۯ��v��oS�X8]f��u�=��.���(�� 9*��)�l�@͝,�R�۳�^���~��E".�qp(ڌB	���!��P��RC��A$G
l��%�
���/0}��y����~��R��f5���G+u��v.6���=�E-����l��v[b8l`옳=ޗ����VV��My����+�W�@~̞+:�y��ہa�!��8M�z���SWYZD3��> (�V�m%
���Yn��[,V�>�?y6�A���n W��}�Ò:f��M{.�F�x�؞��{�Ⱦ�����C�Yu��kw��M��h2Kd����,���������@5��	�uQ�Ȕ��Sʈs�7sˉ�ݨ��$N�k���wt�#0�(�T5N�8^>?)�[G�[�y�'�OU�Et��u;�.1�&p�}��`�-����`^&V�-�*�m�t�K�2�}*�zu��}Z4azh\v�&HS4l�u�`n�W�ln����t���⭦��y��D=~�k�VCuY�wN6eb�͚�wj֌Q����0�=�W��	^�O|ϕ���6�˝�ʞ*��(�7*aeA�Y�q������.Dr[��V�eиʯ��szBH�@,�:�����D@�p㷤I�H�01M�.�h���+�]���㛶fv��)E��܋	�k���lh�GSj��d�c�u��a���1�=}W��箵-�O�..s]+�7�屧j_h�U��Y���n�K]ǙTy�er��x������:��*	�g-�'�=�hSY3-��fϪ����D�ۍg��7�vsO��:עCk��{Փ�6�����Q��@[rr9�eӃ(e	����3zH��͟2H��Vm����|녝O�8�Rj*�߲�Gs�3ž�T��w4z����\m�(�.�G!Bq��S��]�{в�-�.����A�������I%�x�+��P3Ě;��i�W�;�z��(�0�>@��\7�����1C5q���t�y�Į�[��⍽��}ξ�g$�� ��P>d�Dv�^�M�ݢ
�����n�깞����sŅ}v���o�:DP��ǧ�߳��`�~쬌�5��n�~��8��c�W�[��Vr�M���f\d۬R�����Uv�TXW�S͑갅
 x�� :�c�D�{�ڷ|���dJ��a
�s��i��d��+\�	c��i�֔�Ƽr�D��,��-9�&��Kvݵ��Z�}}�5��x�o|�����c��e4����LY���xa�c�NZF������ᱳS���0���7^k;���ޢ���1���OB�T���]��3m��ml잫��)�1!}�23�a�f�mq$u�P��z�Z�T1�v�x\��tJm�}�����uк��g�s=�~��X���V�i�<�T��ck%���Dr�h�㡭1����٧�13�.�y'�X�Z�������{$��S?����ʨ��&���y~�i�5Bp��e�-��vÈ�',dW_�2����wT�u7��C/fO^`��L�N�l�N���ޘd��z��wW�i)wZ5�;]��ZYU��h0v�?M�3�u[_��pƴ]�����=_&�������l.�vf�QO���b�G��%��I3�`3� �~�]��Q- f�TM"�����zU��u�Tž��v�6�&f�ղ�RSK<x�@���,���Υw�DV�]�i$t�C5�rK��B��4��E#��K1���L�2���|Z�V���K~�dn��geEs��}O#���";�V�S�D�Y�ޥj��T� �k�a~�&�i�݊�V'�K=�̺�f�C�<n��#�{�5�t�s�%�Ku@Ίw���=o���)�7Z����`��,J?�����}���9�\�gJ;�m�k-��J�ot��[�+[�f�	m��z<R�Ӵ4��[�|b���(�#�TU�Ⲓ��c�N}��*����������f(�u����m���v��q���9�ex���A��/��8r��Z�r#��q���{|#��mλ^T�2��s�j��ٞ�g�<�d#�vO�de���2!;�<j%�Uߗ|nL�vK-�������m��{�z6%dq��3R}�X�޴����A	?ky�m�^�dm2Z�$��n�k��ܮc˻h"F�!q���˫-�|�����V왔��TM�u�p�/u\Ni��ϸ����PՍx��M9�V�}Oʩe]��n}�A�F�'���ߙ0HHL��x��E���1$��	ʛ�Cl#b�B��M9�A}U��q���Z�A��Jڶ��)Թ󬸺���u{�4Z;m=	��w�heԑ3�C�	�d���Γ[��[��	�u�؅��Uks�ـ���:�܉�*����������B�Y@w ��vQ'Z̙��w�T����.��Z��%?��{j'ٶ
���<zPg=�)m�(���[�H����T-֪��p�̑�)Y�׍ў��s5@��].����	[�}ŵp�]���_�'�&j��]y#��$r������/ɫ|~�����{&c�)n^y�r~mt�>:֥�:R�~�/=ZY�c�6���\Ab$<5����M�ӽ�_�$�Am��vc�W���m���w�.��z���i`ДF�����Rؑ��ܱ����}%N}��8/�j�<h'=7�c���R=3^و��J��!SI8-�`�
.%L��3)g�>� �Y�h���2ʀ�ru��Y=s��nb.�WwsO]l�s��S�a����{�1]�G˾O�f����l�=�G��V�.q[n�>�K{ɖ5�vo9�;�5kɳ|�	V���Ƚ�&nӖ�n^N(�y1EN �ymi��eF�p���@`n媝�B)�Ќ&���9���E�d��^��Ru9�6�����o=V�������I���u3?a��9��/=���]��}?��>�~�w�Z$�9��7\�I�]+�8�7�v�n�κ�Ii�ө�R}p(�N�<�H��1!�}k���μC���^��)̖���H+�O���l���l8>���y��>EbK��RԪDf�s EQ��}�*��zHdq�>�y�ՠ�����<���9���2�%�gF=*��-�|I]�
�jR��"}�]j��w��5�q���'�ѫ@�51�wa�@g�3J���2���=��m��󑫹(�C�O_��������n1�S�r�}}�`�����f <E+�3����'�os��9Y��H�Y>�kk�dH;�.��Sh�A���+;[��s@�7��_�:5�������'�q꿛dy_��64�to���pF��|��� ��1��h�o)�p����m�{��KW���u��M�5�9�t�r��Z�:��Wk�1�4f�ԑ6���V���(��o hV�B�6�[ Ƿٰ�sr�V��x��L��̧i�[���N���$�^z����Vn��1�9�`cel���ٲ��Ӯ�e9����LA���F�[]Ư/pD����3ϴY]��v�r˟�C>��OY�a^�`f�k�0��ˀ6))�^�tP�JR�&���0Ι�����L+7�����ϟρ�ö��w��5@j�Xg+vVĖ�Nx�v������H8��>�`�l���b����Ri����so�F�r��;wϓ��ߗ������6w�t��o�C�x�w��'n.dՊX���{��p3�yDb� �݆~<���\��z�@�fx����3x(/��b�{tѽ�+!w"���OrO�����ߡ�h�~��\T��ѩ�LUw����x|��lǏA�>��T0c��� ��\���b�CJt�(�^����6��U�ͧ�3S?N����
*f=��POX��1��Í��F�I�w;�n���`͂�T�q� *��z��U����l1�uj� ßWT������}ظ�^Z�{<�@���*����S��۬n���w������J�C��:�o�^�;��)#�j�t=<Z(a�˻�܇3�
Լ:�0%sT;���Z�m�G�4�]��uک��͛~����=�o{h�w��5�:D�{����wl���aZqf�Yor�J_����N�ϊʖd%������W���㩼e��|d�����Jr.�#�G䲝����;ۮ�i)c,�f���Li����Y;�պJ�]vٶ ����$��!�qn�{|�P�'vƒ�i�2�F�n������}g�`�����r8.�ZQ-7��	�S�
��&��΍��ד����֪
w}Ƞ�@wY>�[�2
G�ST���(��Ȍm�i���|$�,D��ܲsy�D������
��w�����En4�g�<�Y]U���RN�	Z��<3��)��h�D�|�;���m�NPO�F�{�>�Em�$c�m���z+y��x�����f�.z+o��k����8�}��T��L���e�.��ӕuɈ����rcee"�gOT�Nv�R���`���3�
͋9�Ų9�6��o����g��x%��v�ٛ��?r��Y�8fT����f���{Z�c��h4�^�8EZjE�{��D�	/���.wP굃��.�t#T���N�48��Gn[Z2h��\�g�g7&�],ᤵ��bNOR�;{����[�169��at+xf �Y3�$`f@�ed���H_��ŕ"��n�0Rmɖ�zȝ��ki��l�8�nT�:C\�wL"�&�FL��y�1�V�2�=��>}O����^)f�4�a��x��ڦ}ق�v�Gj=���ж����DM�	�:��~Y]{�;�}���o|�99����S�&6�H��j视˝f��ঔvQ6��Y�G���n�G��T��l݂��U�u�r��6.6d.:�*Oy\�D��w��	�T���A7j�c���̏5y����*J��3�Ke��}�جHΛ�9��ꮝĂ�d�S���{�&����
h�ej�1Ũn�Kf�W�v#e�6�SFg�rV�����D�lP.���R;�]����J��39&��ȿC�Y���*�� ��%gP:�^�y��[��b��p���2�Y��I�רּƒھ�vL�eI���-�FMg7 �nc�B7�m+�)&�{8eXuS�7���0il�y�Lm�e/'��e�}��+���iv�-1ua�����}	�25c���������D�o��D�S���B]Bc`Q��T-��N���ܿ����o���7��r�l��-!���wԲg`>tϷa,��F��j؞�Ba�{�X�p��=�Ml�Zg8��>*����X�a6��1aY==wӺm�VM��3������ᅸe�"1��|.�p���=r`�Q�JJ��B�t��?3A���c��[���0gx
��a+L8�ɼÝ��v�Q̎Ս�������[0z׾���H3�eV1Y�t���E@f��g��KFf/<��Vp��d�����4�l��z"��mDe^�"7w��^& �eSg�.�l_)ڽ�^AHd��R_tyg�{̈́�"�g�K%�����Ӳ2��Q�ED�J�P+;�Ү�Bn^�/�/��v7���;9Qޔ��v7��8�\����}��O�����������������{����ޞ�������gy1�N��8����\��Y��ѕ� �Y�UN�m�f��N	t�h��9yl�{{:i�Ҩ�e�}�"�'V�S<�7��c_0靡��x:rk�v�� ��Y��Y�ѝ�:6���6�p)���uś}ۯ,�`G���cU|��AӍC{`�hun��,�y]��Z��|�t����L�Q	��b�K���X��Nk4ud��ػ��N�Bv��mn	|��1�w��kp<&���=���GyP~�z$n���v�/=�5a,d�lp���ᐺz%�XY���4b=-nn�6�t8Ƚ��,+���Ei(+w�;e���Q�m�g�#K�״J�ۮ���P�]�1��X�L�;C81�.W6Cd<5�_K���9gz4sun�kw�L�:���n����k�NV��]�3ɦ]�,<	���>oy#:��5m���ں=�2�p���B��0��n���quk]h��+�̣n��j�Di�{A���[��:��l�5���9�AlǟM�X�.p����(B�ݻy�-��ޕ�B�9�s�L�iV/u�,�(,7�=׬+a��g5�A�+ehI��z�8��X�W4 "���!}�;r����K�{F.bP&�er�g
a�䰯�q.����CV������m�6�-gp�9��n� ��)�J�di4��F`Z�i�W����ͼ$ũ��3��gZu���X�G�K��74&�Fny�!�gN]�Y�c#y�g+=�v���f�ę\5ᢡ��;b�c��˛�R���9zV+$�2�ը�+����-@���9��]�fc9�d�:��![�q+���z�ͷE�v:��E>����T�'���|Dr}[st[O��*n���ڻ����3"�t�̱|���\�N�Q�;��T"��V�Y;�6i�v_l]�V�����+Wb�L�r"[slj�2g^�w^m�B�MJ��{��ۖܜ϶P5Pҫ�#�F:[N���)��ۺl�y�t��	�jb���ёD�n�]�Q%|�9�^��mgXKˍ��J
�R����~�ؖZpa3S��\�6��F
ؑ+s#S=W��t%���$� �]umO=5ga}9[	'ۺ�0�m@��c�Z�s:�I��maǦnM�\�]X�մ�(L�+2Ib
N�U��	R�j"��֯�Z��s�ML-�g^;������58h��/d$8R✐/^V��Qd^�G�释-,����L��A����t<��Q�a��OB{_P͋�����d<��0vd�kuz2�wN���@q���;�_bش+v��7,��n�ˮ:�@skA[$�mޜb�N�e��
x�nʒF��;9�:�Ø,X�P���h�.*�����-��棞�.G*N}P��{�j\�*��[�������3^�΄\�,�e����Cz�j��4,�-�-��s{�����PX,����P�� U6`���sF*��
�ZJ)�W�a�I���ǩ��DD�CH��T�{�E]Y��|��DHP�PQM-?#E%!ETA�b����&��m�@{�\���i-��Sؘ��q>�9O��
�b���N���RP��\M{�*��"�A���d���n��))(��RASc��M�M��ABTAA�~K���i�ܚ)(9��4LD{������W��5s�PZ��7�#H�(��P��u��lF޸i>���kI2שm�>gQ�U3C�֚�1����G'��
&�~u��5����sb���sa��� �����WX�U4�^��uT@TF�CF�EC�zgמy�^�	-������R�C����E��Yo�ۭ"9֥F�C��$���/��t���6����2�N�j�}b�������Rm�pM�����=B����~��U���⭖�b�j�u7)�6y����Ovl���@��e#Ot��K,���ɥ��X�wc_]�0�������=Y�D��G)¸H�+kͤ�l�Ԝ��%v�����z��.�N��͗|���Ȃ9[���{ɽ��+�/ۯy	�j���+�jU#�w��L:9�uK�L+3q�))oy��I�!L��A����RWCp�W��;{Pϼ�����ot������l�̴���A�+ܹ�B��.��;�m���m����wM{����-�q�����8�4��8�\���?n��]Aoϴ;.�7��~�w�}T3k ��/��1i��o���Pz	����v�� �3�
�ޛ�<M��b�����>]7�QD�������w���Ƈr�^�a�Y:���f��J�/`3'X�\queo�����*�gj�H�U�ݑ
 Sf�Y7���i���Fv��p��N��D�4@[���iv#o�̼�,`�y��o�[�Y��2:.��=��X�#[�  ԩ�
l0��ɉ�2�a��n��}��<���������>N��k��z�a|�&Vϳ�yP*"�O�Bv���u7S؀���O��M�|����+�����˼f��%���m�j�:vg���
��j�h���Y�9 1U/f�:B���eL�Wqǫ|�K��|Bz��Fc�ڞŎJ���_�B{ L�`l�����Z�͏U���sRH�ԗ�г9>J���n�>H�X�x�UҜ���[���*�"���K�V��t��u���S�e��Y���Λ��0E���g�����Šmj=l�O����3\541�q�1�����r���܏dR{G~ѓ1��l�кm8�-7�H2�wrG*��({&��:GK�V��ݡ�{��MU��A�==^wn�uR#��d$Y��H˗��*�]�d��L?q����]Ҷ�Gk3�O� !��ߟ�]�%�\+����q;���3�ؙ�E����Sj����[�~�VY>;�]�5e�.�����nMFGW�b��:�l�,�ekt��vi�`�b��o!+���b�nc2
L���!�
ɉ��٧"M����6�T̤�V�oY7znd+J�Ò��3�!�X�m�mq��7
s'���7�����y��K�7��wVXH�[9*�_g��,��ǳ(���Oofo
lL.��f#���QX�E�U���p��r�xGU�~�;7�x�˃��0[I�5��&<��c�&�;R=��ӭֺ=d�����gw��l�I��Pl��'�^qO�%���Vl_`�[�ٶ���.���e��x֮�X�aV�x;_H~���w��ŕ6.{n��3�9u+J8;���������'�$���\.v�����U%���:��x[םyDk7�r�ʸ��<Fb&,�4��U�T��N�s�>�5��M�+�a����n�=�ٚ,������y7�JdV�@�Ko�d��-P�ƚ����^�vv^�ӻ�鍦=R�P*/�ֺV�
�mj�]f��m�T�ki4.x\ő��h��ʮ_SZV)a_c�{�R����id?,�
��t6<f<�6��բ�N{�~ӅMo���wRw��=D�$��O-�u�
u�:���g�*j�q7���Ҟ������)s�����ƖNj���M^Z�ԎMy��t���3�q�y�b����D@ü޺�%[,��������o7="ѫ{�|�k���_D�ƕ!��S��r[Y��Xɠ�[3�����Sx=cT���S{�#K�ҭ�W��븞�qu4?���v��E��#w�s�� Qh���ˍ1�ũ8<��������f�nK4����Fr�Z�@��p�0:�Kħ�?���>/��}�]�eUG�y�B.|�v|��)��-=r!ʟD7��TlR���ן{o�*H{�{��Qu�ͺɻ�� B����ˣ�þ��.3��+��Q�k�v=�í�Y��E�^��%��`3Q)�HȎ�>��)�C��Χ]��!st;Q=�3;GL+[{��5#z�����ao�����{{��gMh��>歖	8�=��Yh�$�1FG=26:}c�&�k��G����+j�T���7�_���_��ܗ���%O"f#�}*.���i�z�Y�蝈�6ư���!�<��2������M��.�/[9�i oe��D��x�Rpi���M��ם�R�����}{؞Iw,��N,K]�>����/��}�;2s:��x2-�*�%��qFHRZ46t��Z��D��wu��fo�)&�����G�C���w]ȧ���*)��X^o��&��b��IV�%Qժ���>V�Mr�������-J�,����U�&ѭ��IHc+�ѼO�y77:�g����T]��m��wR�/]WBt���D��V�^ς�(�� "o�	�Y�V�ȏR�x���k�j�t4����#9��/R�0��i7M�W�=ǦP<{�Y��,��fU��/D��Ǥ����/��R��:�
���)����.�G���cQ����ݩl���s�`ӵKe4J���~���6���Al�
ᘖki)3|M�]X�5�휪뉬8Y�jȝP�^�g�$�2._4�.�}��z�zt�\TX^�ũ�CctDf:�A�h��7-���aq�������6��^]��X��=�kQTl"�7ݰ�BƜ����;+ل7��Q����[��x�`z�+�ڗ9�A�@m��D�A\����UxԮ:.�ك��+m��l�.���9���ski��.TP��vޗ͒%���}�ǝ��Q�{Ѹy���z���//��ʾkhF/C��ƒc�GZiy�?���p-Z~QV��	�N�n�Ixș����\��աI�/�ao9�+ݴx�K_o�a�;o���x�R�|�Yvs*w�2W�&�n��	唳�5����o���0����xңk���ĊN6I����y��ʘ|y��\����;~��;[��j�y������v���=�
�/1��ún;��f]E��`�l��͞��=ή2���H}p��Q0��M��vُ���}��Լ�2���1�s4$�#�k�=�NdjmS�h=�^�5T՞��4Mչ��^^�}G�j���D�N6�&��f�9S��k2�1U>�cH�n+P*0�v���>�GP�s��Pי�/��}K�����b�|�Kh��6�>��_v���!�R��d�܀*��ޓ���J]V���VVz�a�J����x̘�uu�wj�� ?�o)��d\ Zې6#�n�[d�N)��{9Fh�MLb��ݱ|l����aN��[����p����h՜|�����<���տ���{gM���@���y�c�rj+)�sd�.�)���,�[��ۛW�ܫ�ݧV��Ak�F�s�e�:T�Ww�f�C��Y�2;�Q;qܨ����Íef����ۗe�5N�Nj뛙ٯ���\U��e5�R�g�C��5�G��pU`��*:�Q�8hp螺����9��5q=��-��@��Wt��l�N��/s����cq��ʶRun��8�B��9 3�;�}[ڦ�2�������E�wV��"������H.�og������t��3"*���R������;�eJ�3��x���n����-jm�_إu.n�=������	�G���LB�1yڊ�צ�� yt�ļ�}.)��q�3��tZ���v�d��}>�T���3��svVߍ�
q�Ib+�z����s��q=~}�>�Z�(�Y� +3�ۋj���&T��[8;w�����Z��}�pO�+2^���k���x��b��,B_ق�.n1��[�j�,��#}���dq ��9[�Ζx�j�g��Xh��U'����U߉��hK��P"�f�{���KvU��D�\���<��Ͱ��\QL��Yn�����;�{�zmss>m�\����|�� �s.�o��N@o�t0�-	S�Y�L�N���ѭr��^Y޷��w{�Pɜ:`y6�QyZq�"���i� ������n��}�(�6}�\T� i��*��aU��e���U�t���ûM����Ʉ�ER2DV�|�@���5c6)�Ϊ���N�^Q��б���`���������� #
�w �
Q���p��9ç9����R��2�m�(vǚ���KU��R�aS��*������A{�&�#ϻ에,�I7j�Y��H�eS�`�]�@��^�[ٌx�����Ƨ�8A��{���U�[���'�Ԇ�S;���8~�G:��{��1��<��1�ju�x���ܸ׃i���Q����tj;�3�`:�3����N��	���z:a�ĝ����\�,�!�#��۲�&�s�F�<rzh�f>c0�4סʑ������[�Hu�R���v#��Y���ѵ�S��ݩ��C�vz}��<��xu�i{�|~[�懖ЃoP6V
[��ٿo���8 B��}[2M���b0�M�� JyN�:���b0���85�A�"�1{QGc+ 
��KOB�l��ص�1pL�z*`��Ԉř�+�v�V��K7����d=X��K��k���������/�?M�|��,�rg����o�n��6��]k�u��jߗ��{�������vS�����>n⏺Q�۷B�k���y�?���[�����������d��R]�̳yym3aʿ����!��a"h`�{wh�l{����#J|^�U�����Ѷ�F�������ļ�pn�J��F�$�]�{��*�*D^$�n��X�L�oS��͇���S�bn��U��sS����Q[�)�U�����dQ��L��m����l=;2�=q��}[sa�:�.�k�q���<H*��[I\�W�w�]-w�G�t4��S�Y8�k=�z���T��g\��yNiY�rǁV�e�`׾���2��k�O[�h~>~-�=Ml*��n����y%�gbUfV�ݔ �w���mʡ-�,+�?��z��Q��e���[1�0��W�WʯERk �������aD��ۗ����hh�5�"�J�|�t�@Z�Zm�3�;��ԛ�m<][J��X[�+���P����Fmc��,����:�ק˷��cĹvld�>b�k���*�jZ4�W�ȎK�7���~�Ѱ	lp�q� ���hkbq�g!p�=w4��S�t-�5S����3n֨n�ٵY�Ϡ{�����􉨬����t�\m��IL��~gz���e��,p��4O>K���}�6n�;��D-� ^d-�M0Z���͎��8���<��"f].�8��#q�l{<�}U���KV_wS�n�%���VU�׫�x|w��g�
����x���M���W���L���;U4��[H�ۻ�����m�y���L>5�ejz�tfp��xe���(�e�@J�O��v�M�ޝ�U��w�p��u���`��}��;���뵗�V^/��˻n %$�SM��]QI߷�e��G�xd� 5�iLv�>z�?��z*�������'�{�����WUU�7���_�%E�T�p�c��>�n�S! � L�0,���0,ȳ(�B�̫2,ʳ(̋2,�3�@�"� L2�³̣2,��2����̫2,�3"̫!�0,����+0��3(�@� *̃2,��"�0,����3 ̣2,ȳ̣2,12,³̋0,���2,����3"̫0,��"��2,ȳ(�L2,��*�2�³*�2,;�C�t2L�2�ʳ"̫0,��"̣2,30,ʳ*̋0,��̣0����L�=`0��3�0,ȳ��ʳ"̣2,���2,�3*�*̋2,���+2���̫2,2#0,�3"� L�0,���̋�L�0,ȳ̫0,ʳ"�2�0)2,ȳ(̫2,ȳ(̫2,�0�ȳ �C
CՓ�
����!�!���0�aT1   U^��*���0 2 2�2��� Ȫ�" C*��  C
� *�0 2��ʪ�*���2 0�
� 
�0��� �!#����"�� �(�"�"�(�*�!�,0,0,0,0,0,2,0,0,0,:�2,���2,��(�0��^���z�=���eE&Eh�����~3�������3|�� ��o�$�~�����3u���v���Bl���?�_�>��@y��������D}}$  *����b@�4�����>��C�@(��?_�~���������������������_��PX�REX�P"U@�	A � BE@��P%YUD`	T�P R �	B@$A	�P!E�P$aT	�P(A�!P���XO��8~)�h��-
�H�_�~��w�~?�����!�=��ϟ�� �
�?����:�����u�'�������"=����ڟ�
 ��~�?�~�g��>H��� U�H~D?G�����ã�� ���~���E@{'�����}/�=�A?OA��C}�'G�z4���p��
 �}��~G�??����
 ������N`>���>��������������C��ĀP^ϯ������*��={����C�Re���p���}'�p����z��_A'��� U��¡��?D��:�|�������g'~/�PD������ �+��������2��b��L���uf@ނ� � ���fO� ď3紽�j�"�[b�`�U�����thֺkj�(�]���DQHh)Q�j��R���P-�V�;w5E2�*�a���D�3���U
���%ARUJ!)Hn����뀀I!);uң�UّA)*TV�J��aH"-��N�V�v.fT5����q�T���EUt��.�J6֙-iJ�I!R��E�vҐ���]`�j*�T����B��WFB�
UP�쬉	$-�mT�S^   q��ť{�\��u;{���b��Kwk��Sit�ٵ��M���:�L��d(�i%���]�Uխ����:ql�(nîWD,�*��V[(I{d�)QJ��E�  �4(}���]��
r8B�
(P����o�
(P�۬�:(i��U���#T�m�-���Ʃ��Wm���-�*�����N��5�5��.�:�7mNRR��U@D"*��� w}��}
n�n[R���[s��k55�kh��`�.��w��WSzݝ���릻5�ֶ�Q�H4F�Z�B�[dj�*��	�[���iD���iT�fB�@���  �SY})�i���*�u�[Yw[�f��Ҭm)m�jmd��� ��0 PY2����� W[���I*� ���C݇OM��  ύ�T��2�
��KE����@m��[d	c`�PS�r�� z�v�hcd���Ք�4Wl�AMh�kl����   ,�R�j*�{\��Ph[J��u�����8�UYwg`�Ew���
V� h�E /C	Pv�i(#Z�w/lR�I! _   ��h�Zik%l�5��@Zi� ՚  C�(�` �4� h  o����w��UH��R���Z�  |�  -��� ����m�� [vp
t �n��F�v�4 �� ��� �� t�=d�"zj(�Ԅ�   7��4j�h� }��  ��h � sp hh�0( )h�T h6U�(��`4 ݥ�	�BwaĊR��   >  S P��ܠ �h�E(�d�� �ZS  ��: JF�  j,  > E=�b�� h2Oh�JJT � 6�PUPɵ  S�A)J@  SޣA*��� $ʑeT���������} �����?��ΰ�ga8�]p�p����̫�-9�M�>������o�痟�01��l�cc���m��`cm�� �6ɰm����a���L�迪0���ؠ2O�ӎ��*�D��v1ϖ�/d[v�4!�
�	�9�1�ԁb�����I�O'fҸ�v���U�i5�n�v����<[�;�%�}���T5�\â*^i�R�Ǡ�K�c�"cs.��q梄��)��Y)Q�-1Y�7h챧�U��$���Ü����P��3G-��ʻl���B�M�2�A1���!�1Qʿ�-�>������aK���Ә xUI[-�4�8��V�c���˩]`T��Pܵ�nт��1!�5I�ۚű��i�tq:�N����*���v�SN*�)1�U굍��,�7����x4V���i���G`h�l|�i�+m���8����[p�̸K�&eE1k�h��'2�B��Y�[#1���Y�[*����݄F�?Xv~�`���m�7(�&�M����eD1ltE�dP�u,x#�͸����L�Ε+O ��{@��ζ*`��+�fҚ�liK�������x�� x=,�ݩ�TB��[�r�0�	���[�wu���Y���1�4g%��J���y��J�H�,��!�Q{�+[�XyI�,��PY�N�b��Ď��`�V�jv�V��1�d�ܵ��CP��@��ډ���[F�����7�k62�osi*Y���M!��]M��A�Iw�r��v��zZ�a��ů]�J�o�Pwh���+T��Ԋ��@|�+�*�0L�rdYN��2���m�[�$ՇL�
�R]�{�����-݂�G��&��Bձ�3X!����f��JJ�Uӭ�L��F�3C��ԣ&�Ye��݅Jv�[L�W��8FD�l�ʰFj�R|X0�� A%o1����&�/FU;F��O_����+�{m�(D�l�a�ŵ�q�$�ʫ(�d��b	 �
��n��44F�����/R�lۧCK+.��ove���$��YK4��r�i:T0�96�Q%� ]�p\�BX�����n����V�LGӔ���kn��'x��6B�[�4��+NV�j�Xn�PS�PͶ0LrG;7�d:�Ȕ��ƠH�V��D<�@tR�h���[��E��2Tб[�^�r m�;��X�I�g��(�mCl5Mͦ�i���hKi�g�7s6��[�`��k�+R.R7i��76��VKW��u�b���5v@��M�6�0��ȑ�l'V�IX� �+l|KȚ�m寳���y��="�%���`��b��C�2��r��6�.
R#Q�he�(�am0�c]�&�uy4K-޼�`�ՊB����HS*����AeKXR�ϕkO�iaɛI��%��T�Gv���Ik{�;�%�Z���zb����<�#B��P�1#ݱ�u�J���EB�mkWF�(2�*Y���̂޹����AV�X�i+�37lP��j�X��@�)���!amab���w�P�N��Zak(!��������uc�,�V��d	N�(��j]��� �rԚ� ��ս��љ��F$�ɮ�n�+V��R�\ڂ,w�Y�Ǩ����/Sf�K�",���Q�WPeJ"�n�@ktm,{{���u�C�݃H��6Թ��Yّjk]ݰ,�E}�G6��P��hNwL%6�fR�+Uj.���RR�s-��P;����x '1�۲��s)��!e-���*2��s!Ӈj�=�A�O+Ơ7� �]m��A�:?XR�i������r��M{.z-˂ ��tɠ��]fu��u�ă-3:�kj�D�����2��ԕ�h[C���֮	�^d�cF�2��֡!���Zo3�U
׶�;'B�I$�kL�#���[k�#ks�$H
9A�{f�WVBt�ZN݋��mS�y-����M*D�ʺj�+l��z؄�y�*j���mȀ�m��z���1SQ���u��3EQfb���1$����Lиr��M0�x�.h��c���njn������乘�>r�[n�޼"�cdnP
�r�VA��kq�یVf�j1%�3&3�[�=��ӭ�.��� i�f���x�\4�u���`�	������KqVGr��r�H�y��&���D�a/�U�	Z�dZ�E鎝��f��лv�A+��[���� �v�%�%{{�2�]�xT�����\A#N��S�����M�v-R[�[2�ĆBʝ+cmXR��n�\�-QmB#ݰMh�7k>F�k����x�b[�j^��J��UOmR��h��%����QOnm�SZP�l��n,Ɣ܆�5+a1�t �����建))��6I�5-+�HF�V�A���]m����>1��X�9�����^J�S6��ɴ2�dR���,DıV.n�:u�y'�B�T5+AI�k2Paia��ⱸ���$���Cn�5W���U�Ҩ�G�t�Њ���J(�ȱU��k�$�W�i�v)M�qZ�@�6��b��ܦ�G4�4_�U�Y�v�ȷR�ҥ32�H��(����5�7Z�p��8n�,ܺP�J��ȇ�Iłi�*��p���n�ެ�b�]�L,�#/m�Zf��j�pZ�uzi�ei��{)ު���KE�/V�CZ��b$J�� *0�{�M������&�Ϟ��n9ʬi����:f���t�� j�1k^�Y%�zQGA�\!�֊x`����r�nbaͦƵ�܍�kP�w%��%�-��]��-JQ߆aMm��.�L�i���)��v&R�*D�k1��qRv�ڀ�Z��\	�*��j��l���sLâ3cL�$�-��z�7�-	@�w��6:�`�%t���e$B �:鉋1Q�r^�5�ccv��r��^s��,�vu��F��ntf��i�f^e�u�aT�Ѩ���Dt�Vc8��z,��EHbU�we����'ۆ����S1P�ˬ�wF�31��JV��	��kw$֊�h�Su��V��-��6�������ą˕W"��M&��J�e�!�q:�tZ4�kKj�묱z��c1�`�sl� ��r�F�e,m\���^9XM;q,����5�j���q\#*x� �*[�-�
��`ݫ���UDKu�d�/M@�jgHN;ڼ�tb���ش@�ٿZ]�jR�ͱݫx��q*�Tৗ��N��VKyp�K]Z�*"6}  �Y�G%��Nֈ� �6C�K���Ú�j.kva��FӁe�o�=Ҵ����nku����e��`u46P���v&�Ŭ9���-AMR�ӥ#Z�;i�B��Z�"�lkm�&�Q&�:aZ�
�͡�fl,JV,�Nj�� ;��aSM�4��(`�t�ڗmL�n�h�5���ia}��� #� �;��hՊ��ɥ�5������V[����q��3)R4L�2���qM�+i]Nn��eT�K�i4�C2��"L��e4={
1`�QУ�6"
M��х�oNm2)��h�Ll9l��=�V�壑J.h�$�l7�,�v¨1�SL�5dـM֧U��R�x�������h�-k��mL��e��ud[+6���Ļ��*��A���,��\�� ���n�(}lܤf���F��Sw��V����q�ql�-l�u��35 ��+/D�Z�/E��,�If4��YZ�� ]k�1ӽz�ck` ��1� "�#��'Mk��*�{k!zN�AԬ��K�y����ѷ��u5g���Pc�f�&�HMm@&��"06��nn3����uG0P���]*;�l�vrh���KӴhP��(�5�1�Iz��߀ѲV��VL�#Z��[B��(��f�TsG�r�S�+4�=�1#mfP��~в�� {K��!�,DIj�F��jh�-C��YWP�H�:`hU���VևuY{�Z(�eܫõ{��L���b���S�¢ZMA�;AC�v��6Ӕ�����Վ4-������UM�c��]ŵz���Xw�T�J��%ZFe�?[�p�v���5Ķ�lŠ�%,J=��K��,�w�0`Ŗ.��CU�cu��#�R��I��B��a��R�G��ˬƾ͍գtU
�ᕭk��>$���N�fE(�7wi��Q4/�D?��Q9)��w)�͆T�;�(U�Ê����e;u-
�74헅n��A�+P�q�iL�ӓI�B��*ѳ��Z� f��ޘ���3)*T6�����@�e-߶=R�H�CTPMvi��ۡ,�X-��7I!\N���,s�m��x����̭n[V�ed�4���ƽ[+N���q]e�Ut���^����n桇+�e�x�U� ܚ�����-e�M}���r]4sD������ !i\T���i��]�0۴�D4��j�f^��8��]�;� o)E�?bK6��]�u*���}�0�{�C,-+E*���t�1��{r�
��DN8�e���� �DV�����	��n:v��5�hZ���Ӏ6�m"	^� lk.������"ɻ2`�
˸���%H�b9WdN���Y��3[���x��p��p�|~�@��je��9Pz%��%�]������E��4-ŕ"ו����&���c�n�U�U�Whi����٩!J۵"��{�qǸi����NIYQdP,�L�G/`okww~k>V�F�a��W�j+�"A�]K29d���.;c�f�]+G&*�3Q��{��$�*el��Ol]aJ�j������w�ªh���wZ,"6ީ�u�Ҷ�]7st-����ڽ��]Ga-�f<;)�`6�sl�9�c�xb�*�4TX��/�����Ս:YlCF=���-���P�[z-�����E�h;hU��g��"�#�9��́�0K��w��0m1u+]0�q��RI�)�V3H:۶�qf��L[��2���L�!0��{�a׆ly�8Ե��+t�Y�#���c "���N�D%��d��i�G�Rw2;:�{��ܷug�[�.��-XPؑ2-[񅗨�3��)j�P�5e9��ȱi�o�ޤ;%��}"��L�n��,�Qi�f�[ ������%53����z�n�!��4�ê�ç�w��Y��mAi��x18؎�т��^�u,�����M����6�bM���K��ӕ>����ȥ�drҌ�'c~ǘ�[7��JS�i�͓YՑ��b�4-WL}����a�YM�+3���Q/T�e
 ����mh��IG�q�X*<{���1uuqLh�DL��[b�J��

�wy+(�*l5T��D�h^���T�N�!�MnVI绬l&Yvo�:�{�NL�<�f#(6a�ai.ZI�����F����A�N�}���ږBH�yk�U��i�:�S77nU�07-dʙz���ZU��.�Ǖ�Ռz�*�)Bّ�N��ŵ���Mb}snPCC)Ƙ0a%��jy��A�h[�lZ�	Qh@�a˸��T5v�a��c7�"�yp�l�p�&U:�����)�Լ%Ė�C/.�h1�mf�j�`�����<��/w($�
2�xQud�n@^Մ�EL���%hYQ�͂�]Ì����R	��C���vm osX.ç�\Ԭ�y,�HZ��n2�SRe%�KQSEI���׎^��Yuroh�TP��ʻ�9��T	yJ�����#�Wxk0�%�{L�)
ED�cik�ÇF��%�]�R�I����/tc�1�3l���[M����n�����C������F��M2��&E���sr �&��4qӌ�cS��M �<�uv�����5���e�0����b������z!r��^�fD.���A2'��7*%����i�T�o�h��lU3+-��5�Jaf�e�,]�сFY�p�D2�x���v�Ҙ.�mn��C#AVQ�v���MY�[[2j-܈5,�"�KB�P��;Р4r:OsRK7hOt��V��IX��d6?U��]F���2�.ar�86 
BΈ�7�l��n�j����o��t#���Y�FԽ���&�x.�f�s�M��Al�Q9y��])���
��(����0��4��1���9�\[u��O1ٌJ7hY���K;u1�ŠۉJ�%c:ew���\9���cƎ�2��w��ҭ�(��+R�ˇV��t�Ͳ�'��T��խ�[k!N�db���B�Fmb�s.XT��+.��\�sH[[�q��{��T�, ���o6�j��/"կQ�����6�°a$&�x����ݙz�uub�9>�����Ш��ӈ!{�_�!�؊�b�U%�3<��3C-��[cFM��)������ga�KV����W�o�����/Jdj$�*�\ˀn�r�0m��Mf6Ԏ����pPX�!�"
��ȭۘ1n<̳�>�4ku��a�T)�T��GC/�v�����)M�ܨLD�V��)		Y(9�%��+3l��ILȚݙ{����F�cc7M�̥�,ͫ�~���Y����4(��2^0�m�:�����S��hU�2lFAW�)Һ4�]�JP3��|�H{1����2�iP�ahJ�wBf�8�֌�k*-�=Rab�ԝ�5h���ӡ�����Q�.�h�c����c;,Pʅ��]˚6f�黕4���63E(�����zq�w�T��U��Ty{.ecHA�M��5�Q���1���eٓp��kn�Q�s[
�w4B��&[�"R�ѻ�z���nZF�2�v�@%�6�\7�Iٸ
[�MX��jF.:W�8�kZ��2��׶)�W�oVX8��ƶ�<5�Q�VӋUH�-�]��yX�b+2����i�����;.-��ڶ��;��U{%�IL�	�ct���Ӧ�Jo�X���\�*IMh�ʬ�<1B���R����%y|�d�Mc�X�6/�.��JW`�L]v\���L�F�+���_e��1_-��;
J�it���b����4m��{ffV�Eс��K���M�`zl�a�{��7�+C :�ݹ�]��V�'^��u�VL��u�JO:���hdzt��I.�O�&�KRN���-)���Lh�T���M���W����\�\�ElS5|V񭸡</^rSF)���=#Mү0t�1f��K}caSU��u̺Rrޫk�Vb�6��U,�ݒOX��1Y�QZ�r��)Ϧ=���X�oHX����JJ���a���YYlqm�-�VC	�n�S�ys9fpq�X��Y� F_"��q����7�SG��KA��]֤�\���D#��%4u�v�q̨Fr���r
����ra�޷kI��Ժ����:�Z�[aY���Ӱ�@V]bg�"�ԭj����.��µԋ��������3��J�pu���xD���ٯ�q7Z˒��IF��,:��=1�bq5ig	��]����Z�Gr����x)�\�8i�����]�:ƌ<�J�����2���I]E hRw�ݔ��y��ƗMqY�/�6�J�����m���W�n��vS;�J�g![Z]�SsFa-���u ��9`8���l�+�>z0�zh����V~Yl8gKP�H5��W#h:�t-u�e���N���[p�'���IRg)��ec�Rld�}�@�d��2��晝݋�bϳt5�I+� ���g�Q�c�5vH���;JR�)5b
���l�Jw)9�^=���!�@�^�S�m1��&��N''��7���³��w̭	a�쳯�ܡ���r��±5ה�}��"U��Dځt3&(���ԓL͟s`B�]+�X�:�\�[w�:��ӗ��Z�s��[ω'3 �\����r��D�S8f8�Uj��͋y|{;����:L%�e�t&<g��`#��=ݚ��eN<_^����kU�s_P�-l��\�t�J[{��]�섶�> �ګu���ز,\�[��&L�|ȶ��E�X\�Rqx1�F�4[kz�:2�I��aбճ:j��{4V�,�8�mZ���ˣM��T¯`��0�xm9���a+�ʬ���ȝ۾\���h��,4���S��b�*VR�L��wz�ѧ�=��u�u��z��[|���z���#.���Xς�C���z�=γ��$���d#^C�Y�������]�tjo�|�RG�y7ms��W��R��R����H����V���X�N_`c�q5�5���YL�u�융�*��U�Zi���|�K���h�>��ّvΐZ�%���`Wk��|؞�)� ˗Ք�;�A�Ӓ�X��yz�PV��kb���<�/�CJCzP��Q.�����v耑s4q��zȕO�[���*r�͛�3������
�ݠ8�	�a8�"z#�W�uq���g����+&1٭-{��C���y|���weoW:�s���հkYF�u�����Y\{��h�KAX�˔ҏ8��K{0�as�k |��9ۻ����}B�P���咥`}c>�� �m�2m\o���|��9��ʂ��q#g#-��V�#�{��r7����%v���P��%��<IS�(��ιJf�t�tF&�]�'UA���4Rk(�l����rv��{d���+��CY-��k�۽d
og�K�e��������oR|�Q�n�'}�0�w%P�=DV�ѽ5ى<��w�j%���� �C���֜(�u�������4;���=҂����Vyv�9�f���ô�*#���so�����So���*S���vɑU�9V�o���ݠ�m&U���D����X֡��LւU�lʍ�����9ο1%���B�S�vU�1�0e����f�[��w�.���Ɛ���_$;��m����wy�P���rTw�:���m�������+F���7m(o4��*��u,`�@�*ۧ��r�仱�-m� �����l���Ýӊv�v�ެ�� ��]hcu�����y�t�M�@ݘd�iw�b�?����䮞Ѱ��5VjWQ�\��T�I�5�2/{�-�[]�y��yF��U�8���XU&�Է6�ul=�;���шكW�摒�A�ۛ�
��I��L��+�T�;�*�vA���R�H�ٶ[N�t�1M��UAfdr�5$t�h�wٝY`Y�`a�؞͛}�2���˞#uT�C��.�p��h!�b�����gv�?_gdC�'Ykn�S�W��]��*VƠ�����h����}c':���"����G%u�]N�|�����/Ƴ]��� ׽6g��3j��u�-�C4+�wM[�xLnG�S�����n���C�r�[|��y�5�Mg��ر9T���1�6l��KqL}�֝����1U�R������bI��x1�S�V�Y	J�vpѹ�"}�Ҵ����بm����+-�KM=�34]C����v�����b�OM�f�2^Pz*��b���o��������w���;��F�!��!�ar���"��jg�b��(�[�7��I�㉾��G6\ж�oQ;ɀ�S;����c@�3%�=ѐ��=ۣ6��yV���૽�@8:�
�o[�zi�JSn�1<9|�*W$�]]�_qo58��`���.*v]����u��q�v�5�WCSk{�-{/��enW3EV�r_b|��.�T貯��boN�눺�3(��'Q���n32�aw;5L�rc�Y��Flr��-e��Y�3,�˻hƇp]����y`U��sO,[π �vN	Z�8\�J��ϻ讑]e��l�[�;���\��r�ٷܬ���6�4���c+�����\͊37{yFI[4��0r��i�,y��.��	��3x%���k�K�꽲9���>X)^����,U&uNF���r֒��;q�"����8x���ϛ�r*9K��i�ɷ�2�8��72�j��t����l�G7*&1�`�֜v���q��5nھ�y�*Q����:2*�uf�f���BZ2�4Óy��=�o{dB#��ë�E��z^��闭#�q��iFs-��{}�������z�tP�R��W*����P%v]���2�;�A�N1��dd�L��n��@�(ֆ �K�.�M�+sX��@�櫪�%�����xxs	������G�V8�j	�[��r9m
J�c讞��	"�1bX.R�U����2i9����:V�:K�����Ֆ�&	�`�WKY�JUβ�������U�P���T����2:��(��vp�r�EoTu�T���'�z��y9��N�:]�(��M}��L;4vJK�J�����Mhw&Q�V	��E����˵�0T�/qق|Uc�i�ţvU�ҨF8���#{���ޥ��k�<N��{N�����X�Q}P����N�	i�2�m��uc����f�^9e�U؎Y9d��Q��jX��ˣQ�O-T��Ü�����ׯ���;,�:wjRiV��[�%��T�غ�#��P���e�f0+{�#���YJ�GJ��{2��Az�p���.w[��T��r��N���t32q��Y���6"�����og�e�/��p�QGqz�5o�V�Y:�,	q�w$�d���:����d�#ʱ�����.�Z�@0i^��_:�ݷ��~L���%f�،�����o�gf����9�x��Ҭ��칓�Kʀ�V#��q���#��W�fD�*�����3j��=c
"��l��1�;��̫�(js���[
��+S\��Zf��g"p�@<
�<\�k�^q��.�	���l�I����:��i�V�t�ʞ�
Y�gbɏh*��7N��Q��j�;
y|��擘w��.�%��oV�:f�lD�4o39��t�˽�NM�Q���|��v͕x� vvZ����K^݇Z�t$m㕝�Zy�:Y�r�u�f�s��U���m%�j^+�뗭�Q]�ø����õ�:WdJV�5�5}2���-�������&�q-v�O7+n�Qx6�5Zծ8�ɼe��X��SVws��㒶3\�uZ[�â���bd4�-81��I��,�*sM�We	�a���jU��bt;��S�\�]��g{讼Ŵx%��6��C��0�;�]b�3���W8��6t��j�u<��l5]�Q.V��3yC��gP�yn��;��S⩗��&�G���KWa]�6��!P��%��崣�:��ߣ�;rFy�	p��]�rv�ћ6�U��r���/m�J1\_:e�`�ƺK7���/8G��{ ԹT�E�k��/j�|U �U7DU�7��f̥���(x���]�!�tOa�FC�AXU����h7Āi!Bct�TWT��p�P���f�L�ɜ������`P�	����܀�R�����?noӧ�V�ۧ�~�Y���tY�gܭ^l8�#�M5���]�|M���[\�t�{ ��+v�{�b7M&l#}��U��c`%_>�dor�by�\Y���������Q�X�779��g��c��0*O5G�́T�X荾:8�*�4T���O��>t�	��SJ��hY�:A��}zZ���f�Ȅ�h�x][�;X�ԋ�����*���è7�3�l竊�ò�n��Ơ9#�R�+z�.��&��o��Zg�o+E���-�q��P�st�A��gvf��˗Ԁ�*g�k��6��r �t^�"�1u���dɺZ�u�k�}lo��Wi*u�(6�`�Y9�d���.�v-�%G��6�6�3P$LԄڶ�ٺi����l�����Y���ܲ���7Z\ҥ�1�j��V�'g��o���ϕ�M쫴�����������l������Y�q�5x�ݽQJ�V���fպy>��W��#{*��Z��(�3����y���M;v����t���o��*���Pmm�Wp -D=\OQ�7]�W�
�m>�W�j=�P��{&�X��^�
闥����`3�ܼ�O��Ty��7�ړ9�-��c��n��A����Ռ�"�)Q�\9P�`-� e#Y�֝�}��wC���
��r�)]J1��j�V�����BD�K��Y�v� �|�9VB����
�F��T��;l��R�O*`|��G���ɺp�����H�X_ȯevֈ+~سk�[�Vr�YFӁ�!C0&�]u"NA:oNo��]5�C����C�s���ٺe`�]sC��N�j�����b���uD^�s��;���l����fɵΗwF�H���) C�zby��K�%u�nQfB't��
|�t��޸Rm������r���)�^2�v\[{�ov�$��Y-�M�0�e,�Zy��A�3cZ�hcE�v���fwt�d$��.�m�VA��ձ ��>�}�-̂�լWZ�o(I�V���w:l�:_r�g|i)���Im��֜ˊ�v^�����o��n�sv��uЪ�'�e���G&�B��z�Z�m�w��f����y��K;�/t���B�Xz�4Iu�=�;i�	ña+�+�p�M#��W�(�P�-��E��@����kpb�.)�����{F�%��od��pS�[3n�;�[7��*����P�po�+#wU����3u�i�<�P�G\R���g]L����<�p+\��6]��Z
�eC�^����˥���%m�VGA���������Ip�9o9R�6.��d�W�hwպ^v����q�$_qX�+ZoJ +읍�%R#Ֆ��g�-�jg;��.
n��{���!~�n|���㜥8�B�0��[���'��%��n�S4�iIC#b�1���;��y�q��栾���t�[{��:$;����`�Xz��0��v���e[�^f>]�:j���$�Jα��*�o^2���PK��e�/�;�I�R�{�f�uw���F+jeǎ�哕������i^H�w(d�9�tamu츳�j��R���>e-)����OeTJ b�뼾��"��F�O�RJ���	��oo�#�g@��np�e���jC-!ս���ʳCpȯ�s���y�D������nL�c��kܛY���wKZ���ł��&լ�fӡs���Q�j��񱑵zeV��}1�)jW<,� �1?riXê7']B�٬Dk���V��@8�n�[T�n�o9��"����޻����-���u$���+��G]^�.�q�)wm�e�PS�;�([ht��\��\���V����jiV�A���]-�Ռ�ͼ�!
�:�sMY��|��	��cs
2#fm#;!k��Z��ᕲw>��N �%:��v-��%�|��AtU�ՋML�~|�^�۴;���]���"V�g��Uw��V�~�z���*o:�@�<�r��9��f�`T��On�X�;N^;�+����"�j�}�-�{aR��1�,�ڲ�,�f�|4�y.��n#c�>���3:�A������Qɏ ܬl���[dQR�k�H�E�	�[ky�r�pV?�����oM���6��d�-��w\�j0��5�T���'SS�fv]ww�)�t*�X`N)��I��_e�rX��a��O�U��IU���0�Ts�8��]>�$,�}��Yv*Eͧ�R�:����˓/���4��̔2uI�V�/;6��':_�*�k{]ҥe3ݡ�취�9�v;q�YZ�PUg��0w(���C_<�������6�\}:�����:��,�
f���;�9�j9�=��,�>�P�OR��d�D��|�*]��eΩ���.�Z�7�g���cވ�{��{��01������'�y���������R������ʤge���ڶ�A���78Q�uv�\b��؜9(u�0�����0��<m�_Ҷ��g),\���ŕ�$DA��y��k"� ^-N��fn;�����h�����vbX���A�c!�j�y�1����6o��fNr�=o���1T-��[��ʕ��.ǻV�;-�F���l7G�bl�B�<<���V]�2ѫ	�
ۃ���:�$�ptͩ�D2�N�E�f^oC�.s����%^�����I�4�D���h�f�tq����]>��E*̬-��t{)v��Y"���Ԝ�i׏�nX�g""?wuؖ�b�T�me��p1�BH�(�b�W��ZTA�Ҽ ����SEͶc陫X*���^Z�e,5t9o�}��yw�iҿ�ZYɑ�juծ�orh{�����������/������u|�r�۾[k��B��9���1'Y�2�t#�.�$��Kx����A�{���.un�-���� A��X�7��9*�_h��^:Y�L_y��F�ˤ����\b]р�j��X��Y�P3C���*���,������k�C=u���9
锕�wS��t���i�K��ɳ�oPZ���7:1�u<=M���5��; �mɢ��^�\�W#�뀋i#�|�g(^�EM;I�/-6}j�d�*R=�kF�TR�OoP��t6�M6k&�?Y�-�� �i�ͮ	�4��uph��`��ӎ�WO. 4t��R�]���x�z��V��:Ke��м%ޕ�Z@tٵ(jO���u�����ݱ��� Φh�I45�7�e�a�ay�t
�-	J�Va{Fv��P�ۜ6�҉�KB�t�6»�NC2p2�,�]+CA��ɠ�EdF��
ݼ�ֶ�v��W)�	"!���SŲ�q<83vGS{I_;��E;T�@��l��<{�'�$�Y�2�e��D�˪��
Յ��\������w�&��)�Wn�
Τ~	�Fv��vL.�#%�ŕv
%�������`��t/B+r��W��u�M$�-k�Ȳ�����JX]YHX���H�M �[XZ$�ɑ�Y]͉/9�1;�S�j6�ǔ��wE�U1��<��޹����d�E���^���V��,k���Ll)!��֠]�8�ϴ�f^b�l].7b��q#.*�K紞]�;P��2�i��s�4F�r:Ӛ9�`�uK;ǅ���nPF&3pf�׊�	(��j�z���ز}��6�t��G�!YI�Ύ�J&��1�6!KA�[l�.gO�-����%h��V�!�U�©a�!��b�4~Ҡ�l.�K9fivX}Wl�ʿ�&�	�S�;03�rQJY��hƚ9���U�/P�wT=���"q>Ȭ��'o�y)�9aY
n��d��8k�Ҝ�8T��ի�Q����gR�|��ǻt�h�϶��N<|�n�b���OZ��]��n���O.����i�\Cz�jMA�◢��7;v��n��F�b�vbˁ��X3_�]Z� �[)a��.o~C;�:��`�(7 ���t�{jė���j�O=6��7����{��o�%X�8�)��JX�9�8M��I����.���=�ܸ`���Z��Qc^5& �Z݋�`$�_\2ىW8&b�{���)W|���@�V*L�LB�QV��uA�rњ;_�/ ��}xz�mjmv�u6��t+������ӎ�vcKZ��l�Û'*%��=��V��+إ���yαǋ�k/K�>pIff���3��p��h���o8
�w��P������m���yb���'b�8�>=�e!uiv��X��p'S�+7��X����6�Y��඙� +��k{���l5>�Mvg/��O���D����x5b0���W:�ʵ���	FoS~�F����=z_�U���O�^냋oJWs)1AP�L����q��ʞ����W	}��(:��O2!�݊X�v2���)]M��S0^�gl���[�}�@�XwD���6(�����F��M��[��ycN2o�Gw�5Ѻ���*2��o�g$j�����C2���>��L�S�{�E��MD�PǑ��4�,Z� ��ݼ���G}X��'��U`���F�[�=2_��fTy\���\3n��n;�y��3��-�ԃ��r���w�]$��&!fuu�B�i���W����:��RT۱���nQ�Y���mYQ7�0ؑ*��va�ǻ��l�ǝ)h��2�0�t��CA�Z�Fef�����G^��t�\񙷩����+uz);�!���{�+�
ȶ,؟#��lb��jJ�@���qsJդ�s��eS7`�2�+��S�\=W��u�n�f�� Z��ѫ�f�Vs���վdDz�:��p2nM؝vu���
�P<tk�D��H��YkL�d$��i3B|��Ut��+�g]ʾ��[���ͣ7.Y��Fc��n�<�s't���+��<�Z�HX�Sn���HۻOi	�u־����x�(�w� ³"b��ۡ��9�v�x�F�,�e)���&pWZ*��Q��D�;Kn�S��\:��-���X��ub`8	��b�[��X䐵B]��B2��\ip�@��J�S]N���i��F�鷃s��H�%uй�H �1��"�؋Z�uIQZѡY�ዪ 9�eD�|%f<�l��S���+f�)cI���aa�N!7
6�tx�H��[���j�З�_8��ǯ\c6��)���6�z�2���N�H��ݺ=\(䊟EHZejwƍ�0^�m�Z�·@v
̬{��qqU�	̆V��}V6_(Z2�7hX-S���t�X�vr
��\_U)�\V���d;X#��;ݗ�@+��ެY �#��g<���ðk��wz��ڥ]E�o��u#YMQ˝d>Sj�w�(�x·���W%.�
���֪ö9�G�KM���K7��F��h�/��!�[�ۂ�������б����Q�m�9���)V���qJI��N���T5:�4��=#+����F�u����e��y�i�F��S��5j|+{�k�����H�;Yh<.�Z��J�3`��J�_ewa�`SkkS�Y׷+vQ�c:��ҹ9���K��;���+v�IP�����Ψ;ZtC3 w6S54oJ�;8v�8@�˼����O{;�6���+������4�\�	X^��o&�5�y*88 �^]:�͡9���(=YK	8Z��
�7���"0Z]q�)! 5�r���eo�5<α�J���0>�g�P����+p�4�i�n��f�CZ8e���)�mڜ���ec�p�-@�9-�G�^�3\$�r�Y�zly����
Ky�����r�����y�]a��\����:�5DWL�1gv9 D�������oY�7Mۏ�Q�Rv�&��gR�,�%��7�u���5�oY/]rN�N�æ�oN�+f.���u_�ﴎ����Zt�$,j��t1ib�-u��jCQi��[�ޛ5���;��6z��##�zdUn\u+�Lt�/L�Pր�j���-�=D_g5��x��6�V��l�d�9V,ǫ&pķ|�ݙ�X�x�Iܕ+�fpU�׍:��\ ;�v "����YU�ֶ��uBK?rͤ�wegr��XX\5���5s;;�iU�:Oo&�N��]{k���0r8�殳��#���W�R�����91+���=�c�o0j����Nl��3�����;��@^������E8�I�u�,5��ۋ.�v��~ѕ���"��O�6���W�ef��ݫ�ЇQ<̇n�C+�z�-3"&��������k���e�I��ʴ&G��6ok��J@vslGL�{����p7J���vg�	�o
�;��"&����ff����ɢ����&�ok#�#���f�Z�m�O�X���}:��y7R;�Q�eDM	��>=,ʾ��]A4v�,�̻X���r�B�.�� 9�a���&p.};���:,��yf����+���ր��#f���UϵC3��ҳ��gG�Qu��x�V��y�RM�p/�ҕԈ��7������ZƮ�K}W8j����Z�5.o�߅��CB��۫I@��q������/�
v��V�W�TkL��9H3�IJ�a�)ڰ*g�u�����P�/1�� �0��[.g9�m�4�0�ܾ�2�r��{]
��.]����%u��a�1����+��}F�dܫ�P���m^�R@y3(Y�V�d�	2�@q�@}.�w��{��%z�XE�_ue��]JN�_;��⤾NwL��2B�����ŝ�l
��48SH�o;��YzV՟� �vc���P�J5�Md8b��\�!�1-כ.�,Ds�5��Y�o��õ�o�&A��M�͵�WqV�v��u��S�3h6��o�*<R3�8t>J���ai�ńw_fgc�j�(������Ϋǧ;q5�(>O��5V�;@�壈Ӣ���F[����Z@C"�A�����<��H^���9,�`�Y����:��=��9KOÑ�;��f�(Zb�cȖw+F��v]r���X�3�dC�d��f�q����P�Ɩ���m�wI(f�u#'a��T�&����[V����ڕ����`�����u2��Q02��v�-p��A����8�P���[� �:�	��N��#U7����ru`*b55���e���D�����֤닔+-�u�y�=մ�z�2�WHqo�6ĺ�.��c����D9)����34}�D�x1j��EP�3��=�6o�J�^Pz����)E/ksF��FT��T��8N���������;�����rew/�M�S�G,	Ͳ��Q�y)�I��m�s;۸��>6cX5���t�ŊT�A)V-�Ēڇ�ݾ�����㕝�����9�(-��P	?������z���Pɢ�to�V�[�i,��v�ifn��Xr�@w�D�N���Nѥ�tKٽ�n��4����	k���k2�=�UglV��cN�Q�'e�X���\ӎVwi�khZ�W[}���\3��c0��^꺔�ptEC|���4�!Z{��!Y��i]ղm���;����H+,t��6��GmJ�����7_T�_w!@�{�l�T�������+|۶�S��C��Fn*�xw����S���V�fY�,�k�=�S�d[�֖��M�ö��j!ޝO:��Y����ꊍ��g-`^Y��h!���T���/r*��^0uO�2��edJ��mIK'a�2�Ɉ�#�Gu��(!�l��.�U��e�{���5��5Ǖ�
k�������r�е7t^��һ��E��T�{��{��S f�U��J���;@y� s����RK�졵G�U�٭u�Ft�zz��ˆ�6؁�2=--pe�p&"u�@aڮ݂�e�s)ws��.���tt��b��zI����k�l}�[�%�6����M��^b� �K)��r�eJߟP7�1Ax*��̚qX����'V�ŧ��xR��o�+�o�bA��_nޅ���y���ni�eZO��h�0��1x�wr��D��˭�`���n뉔w���qk�̥8�'�}L�n�NKkN���\�]��)�'��t���є�s�Q��6�:�o�*�hQwtͭ��U.ٗD�vR,���{71Hf���E6�+��.�ؘ_Zt�{]]
�6�]t���3W�޶���u��JV��$n�T-R�I�F�Ip=�Ĳs@� qn�{���PP��(;��J��;e)��P;���|��ݝ��/5+���.�����Q���ԇXi�x�k}6�φ���Lj��x��xP��7��I[U,�$��쾅�2��*a�%�����MN���b���c�Po��J�+1��l�O{A��>�XE(���Wҹ^.����#�k*������.���}7��y����Yԑ�H�lMϝ��;:�4�7��^��Nr s�iřL9�����}G�X��e��q^������/�x�ɧ��d,U�.�ux�X6KȀ|/I����|UgsM����R���XB��˚��5<�l�썱�uhع)KmЭ&B�����5�Ob3�K%lb�Y}�%���> 
���x�y�����nНؖFe���&o��s���-咹d��G7,�٫4l�QKMn�]±E��v�z�b�����π��e�-��Z��{�Z&�b�&��+BH�������l��R�!*[|6`vwT׽eQFu��Mf����ݜt�>\�R]K�-�}�ݬY�i��b���+�	B��Y�٘����T�p����K�7c8 ��>J�nL�kskv]g]�M�V�2�e�[���D���fFfN�79��[�ˊT�ɺm��R�Yv��ڳ���1��5������7��Dz@���f�;P�N�ݺ�J��FS�h���(%2
�t�5SnN����OyR���f��Nu='����6F���7�5�ւ
G6NWs��.��65�
}8��1ge8Φ�R{Y'n���w�/H�*<�X�vr�e*۵�N�t�K���&�[�����B�=6(Giw�ξ�.<��;��g�:���2�����]���Z�Yz�kȧ%�L	f��ED���!�Q(�h.w2%���ɬqצFskn|�O��մWV Jj�&mݑ�	����iiڐ嵇��b�ˆk$19uy`��}�[yVv`?u����Gk8������ܻ!X*q�4��8��z����n��4��vfJZ�2<|��EZɱp��W(vu��7"T3�(�]��,�4Q�S�TcZ"�}��Am>�*��¶���I
f`[һ���-�*C�/�K����%Y�^ٞM\dʌ��kU׫OLp���>KB�Nn���������NΎ�mX�����h�ͬ��g��:$����Y�u�hg��ݕ!gr]*�����q8�C|ww]1����2��F�o�F�XS�Z�)@����V��t�q��S%Գx�G���݋K,>���S�})�M���}���x��Z����E�A���h�5��>F1��炉�Ay�H�V�k҅���F�M����c뼼�q^+�+,�±8��#��+���Q�k��o��6M�M(훥��ً�����)�ג$��Kf���v8���^o��GH8��W]�!fo�<OMv�I�m�:�}&����y}��;�L=k�oz�X;�h/��u�:�v*��)�z�6i>����܄N�q��6ܒ�5����@N���z�¸�w��+1X8=�a2eҿ/m��y_�y���6��q���A�;e���=��Nj���kxm�R�V{�`�
�F��s=wjŧ����Ev����?^&^֭��5��.j��q��V�s��Kd�qZ�!��p̷��vʷ`G+2Ga���{�<y���fgp���tŪ�;*>��p�q��l=�,Sr�ɭ���"*Ci��c����4f���J� A\6�a�(7� ��rQt�V�k����M�±�vvw.9i�����d�b�3b�����ao��]�ţ�����R�*)�'�J
.PQY/�(�r(r�9QUª�VB� �UW.."%PuYW
�9#���K�EQjʻ�5���#�Up�&�
��r��sWT*�#�Qd��QPL�J���r"��L��*��.(���dT�)2�TJ�F�J��R# NPWe�#ZUE7r˵Y��Er���,�s$"�UUp��0"�D�0�*r���D�PI),����d r*"(���p�N���EEr��H�8TEʪ�Uzt��DAG8Q\�.uY�%��T�n+.r֕J� �L�UE9C��" �T��r��fe��T�9ʹEG�p�G9AȯV��QUE;�Q\�TV�^D��s@J��\��+���L˔8s��DQ«�B����?|������W�b�+���V\#_@sR.5C����\Q�lmrKc[�����;Y%��[.�XU�ut��C6UU����S�X�+?�䥐 �<+�lW����E:���Z��. U��}{^Nl��w^����b`�4��DP_��2�[#g�#�a�>fw*���R��t�������L]e��c�G���Ca��
�lUo��첼+xk�[��E~+ig[��+�<�E	H%��X�q#����"��l���Y}cE�G�'�DE��/>�ֻ���i����X��ɘqƔ����3D��r]m�Ls�F���Ow�����RԱ�����>���+��v�W�`��w���XV]U�^s 4.k���V���\?9�+�^���_���}�Z�gq�Ƽ������?*���}��y �u��W�~&P�9��x˫VFyW�����NRT��ꝥ}_z�03&cc���Rb��\�&��J���@����L[���������³O�|,^���`a���p3�6�s�h���u(DB%tR2���Νq!Kэ�a!��ܬ5�A�^��)j���/��#<J�$9s����j<���r�8�r�k��_JO!������>%;!�`􋡸P�v>�!�Hھ��8�T�\MT������e��������:Dn���O�T�aV�ƶ��xv)�6����Bb��>�K�p�{�S�(���qv�
�s��꩞��|"�FD��Iʅ1�����3������Mb['�R7�̧h��wcT󮲸�\��4�}�34H�fv�OÙ:�����3���NgwJ'U���]�%҇	���v��Zy�Ӹ�p!���I�qі�����.+��!�e��ޱ|+����U�QGez��;��}��̥\�� I.%m�}fo�i�W{��$|T%�z��@��v�|P�C���E
=f_³�����!,_!`�:֓�+��L��{o9���?���9��C��d�~�?]�CL*�NE
u<��5�~��'2�7�	=G�+����eT�Z���4����k�mG���B��}'aH�2��wmt���-�nb��L��
i�T."T�Zi�*�&]I����q�����������ʞ����w�38������Լ��Q]�����.�<����� �W��8���T�g[~�~�����IF�~q�AȊ�Geu�њ��媱c�mK| �/��θi�.�#lPD�j\�g�ݗZ�@�����Z��������L�:�|Zc�sp��q�V��Q��_S�^h��*T
ip.�l��ŗ}t�V�n.�J�PǷ��ݍr�5�p`Z��S�Gǖq��iT�Jk�̕��=4��HqF�T9`� <�9��QM4�{7�Y�(���pj�ԑk�N�*��l�A�ya��ma�<7J��o%B��p�T�:U�FeZ�_ a�%���Ӯ�(u�%3�~���a�y
w��H�6�X!���蝞�ig�M~����V'��;v[���͈c����r2#]��Bvb]���K=�:5�r����޻����%Z�y���I�P�~9��}�]/>���9��5��!�2.��G�y������u�ׂ���Z�y��Δ-% �]���>��}>���ӝ���H��N� ����SW�m�§�$7{U�eF8J��g�D���H�������Qϔ��pԺ�+hS�ګ���*6�zs�&L�r���3"V�D�i�/��:��O�w�7Wؕ��6���٘��ˠvU�.��Z*[�=�Xu^�ю�T�P��<9�*SQS"2aIљj�3e�G�D�H�������E���;�t��T�-ybB��6�p��[�U���,k���5�޶�T�p��)ԝ��N�:����um=ȥ����	"{&��&��IR�I�*�{%F��l��(29�۲�e<L��gűG�Z]�"�@X�촸udM�ʕ�tḅG8(���m�'Lj��:aIWn��=|/���Qd���7
�ѻ�)���	a���������#��K�=ם��b�iS�t����̿��>U1�z��c�7rdL)�L<����w2������Sw���|���Q�l��~�q�¼�ݳ�ށ�J�pi��g6�N���uVc]���0��3�B���)0T��-�K���e.��a��t����1in��0u�6]�SyĐD��p���q|���EB�Ұub:����)Xx~Ժ�k�O{�fI����cfk�輈q�g!jU|���B����[Veo�&�1�ڷ��[�vC�n+��I�q����o����J�s�b
F�|F|m�ح��OL���`�R�;�m
;��x�!#֟����^�}+�1����������l�]�e�=p�H�6BԤl�gt��J��F��uIV�����į���s r1؁x��n�N�RӝE�9z]^����v%���ziI�f��	�*���u@��϶� �q��&�a�5�n>}�Ou��ٓ9ONp��cB�w���n(� �W�1�{�V_@tI�cX��t��u6Ɗ����~���7#Ɔ�лd�2�j�w��|׺4)t$�M�'���93:�}j��W�;4��(N:�4�7��Gqv�f1`�<��m���]j��Sy,����Lu����*��;c��^�o9�&
�cVS'��Q�_llO!Q�1A��v��*EpgPi� M-˽U��{}�}�^��Ҥ؆A�����$#b�i���q>sй���^����P���;�t�v���+�iZ�������F�P�49+:������B�,�%��F���Bё�� w7�yy&b���+�T��u������h��ٮ�^{��K"�;�2\��'�2�,[�愑z�m�r�jb<n�Pv���T��#�9��.��No�"7�C�JA�u�X�΢�*��-�3�=ɛ�k���2�q����=�����f�g�q���t��陎d���#S-��݊�i�I^��=�W�`�<5��eElTV8�Q���.�ԭ�e���O��2��߲��"�Z�2��nv���ށ|�u�~����)�d)��5�Jnb�Uu��O{M�܃1���zj�[ۭ�����:r�y�J�S=���μ=�D�|��:���������+9�ɝ��������:A��޽�Q��tu��v�s���'e����L��-Hb�\'�a/-�T�x�05��&�
�eu�O%m�L�`�`�Ь�	\/���D�3: G�]}����fF����PEP��<h�i��B�X�Լ�S��l�L�s�'Z3:N\�k����ms�J���i�}g9/����s�y����\����"y`��g��#�6�^fL^��C�W�6?�о]8>L��Tlz�����q�Ʃ:�g#~u���gL�3yՅ����G*�+����u�\0L�5�o���%�%7�)���O�[�*K^oy�_g��R���͛�N_���n�K�QӍW0�@p���T�y	�9Z�8W��WH�B\mt���T��ɼ���2GhP�22"���$�1���WB/o�a��駔���CU����-=jb�c����؃�����P���r*
JŦD݌��������6>��Eٱ �Z&`˳��܃57��/��z��Q<�DI嘆��JQ��nd�"�T�J���u��HTE����|��;�t>��7��'V4��Sm;�]����	_c��]�����	�(r!��������.Yf���*vԂ�:�sw�(} �=�4�|�
7rW���<`oz�>��#K�*�M�
�>�~�>�+��|���4�rfb�Ї1��}B��wiζ�.c2�o�B�ԧ�*�5N`�9̾t��[լ��k�]FM9�O��^s�����-�t�c�қ�LM�ԃԔj[���w�.f*t�;� �;#��Q��`d vJZ�Sw:9z�l��v��⹜o���ď�n�ff��wz����\*�s��+������ϓ���/�^���3�FE2a>=a�țw5������.��X�F�X"��p���	�<��}�`�{�zWh���*e=}~ˮ��Y��0���l]�\�`��N�:����<<I�4��X�5GD�Z��Mc��a��-��'3�a�q�>�e+�C��=w{HZ0`��Ei;�����e!���5Ck���ȋ}ma�O��)Z�v���f�G�cE�=$��ӎ-r��&Z�w���e_��_lJ�v�-#�,����mZ�C�ty���^����ܦ$�1%�M�u��.J�C�UKp9�ۈ�r25�a�#x_��ϳ�]
ra b��GC.�v������4�����b�D������:ce^���մ9c�!N��c�
TNFI�����=6��v�
��'M�
��ъ�J�ّO9a�9�4�g>}4Ȍ���g��b2�zv�d%�S��${�O}�/+" �:>Q9�%d����_�ic�쮽4���K�|�L��z�f}�؁�J�hedh�EG��..�@��gs��-޾F��Ee}��%�v��eU ���uY��<���5���QuMv�pd�;������VS<�3Ӡ��٦k���(ݹ�E{��^�m��I��ğ-.l���L����v2�w��<x�:Fh,��$�"�ՠ�"D�@hj�y|�w��}�X븧�N�L�=�O��,�����F�fa���l�������!����4xw"^�G&u�Y^�og�����u�5���=K"�pl0#��N���r�������*[*{���b��i*��lH���������tF|D9�\�ԝU����ۺ��b �'�-�v�I�� >��w�K�\-�YnlZ77��f����L}a�y�Cڸ!`{df�'q��'y(*��jFU;+.��??F��,\ �ap�(WG�z��c����y����ޡ,�W&�X���&
#c��|;̥����B'轸LZ����uV�v9�sI͍��Z��\r�NuB�鿓��jv��⊯J�&߅�9[}\az��!h���W.���Qwzm�=b���Q$sÿ?��[��׮Y_b޴�a�����渭"a<�7�#MO*��Jd�,�1�Z!:�
�Y�V��T�p�T��	�Mj�˲zJY�m	zon���w|�^[L����-�W����0(��=+ �z�8*4�`@P���qw%,������b��GHd��v���v�M�nR�8\�;m���,nT]Y[W�98uvj]!�蠧��U�B��]ZU����}��B��;6�Qce$���g�*��i�q�'%S6��u�{��B�ZpoH�,�.6���*���s>�ҬGgȼdo7p��T�����7�o�5+#j�:;�l�\,���U\5#��M|��R��sWT��Q��q�=��{F�[Z�[Ib(i���,ӓ#����\��u3JGL񮈰�j"�Ø��P\]t/w�B��R(?���[��6za���)�<s.��Ǧp@�t���b��rk�w��g����:�
�G��5B[�I�B5*��c���9��i�S����{�7�k��06�<���u[be��K��m96��ԄsO����Y�C��"H:�b_i+�+�T"��e��R���O�dz��v�ޓ�����Þ�Us�� ��n��fs��ɳ=�s@�Wn] �E��T��i�I�\�T�}��a�ɥ�
��V�^�\wn��v�O"�#B����ٙ)����@W�K���[#g�#�{�͡Zv����ܼ��΋��[�h�h�V��6���5d&�@�/"��ݸ=۵��� ��!�(;�O�-��<��6cI����9wL͍�b�� :���r�q���f I}u!+�C��&��k�$��cNfYv^�e ��Ӱ;T�[�p{�r=��nY��-�i�EwuJ��]�RqOv]�^m�T�d������V01���)=ڞ�W�9���e����S��R�=����c1CB�O�!��u֌#铂�t9f�Mll��d�(]��#�Tq^�^�R(l��'Ý�.� �lw$dC��}����WYy&e�/��P�����Ǫ��XV]�zV.���|(J��c:��ob��6�^冴�O�Z:/g"�F������5��s�y �u��{��[�/#������S�]�ގVfYfvy�Zݰ���6=I_7�&+�L�⺽}�WV���%H�}Ұ�)y�>�U1^�#��a~���az6��`0�4���!Pn�D̓���k��V�p���;�[!Kщ�a!lGI���q��e{��j�g�y�5���g��޶�	����r�;*������P�µW��*��78��~��K�S�����>��m>|��#�e�<�|�+� ߫awR�V�f��Mg���#���gg菷���}Km��¢�P����F�#��+ 5��C;�>&�UÔvK`l��mv��S|	�T�d3PQ��|�qZ'�\��M��:�3L�n��:SWȍ����M:̬����|���́i��/�Wt��������1
m�e��i�ۓ;���p\c�Ӻ���[L,��uҁ�:�Τ*{+&�F�و�^W7�k�޼zD�ݸf=c6�p�>
��+��w�h��hfΑ��:�.�}�n��w�v�s�n[���hTw�ҭ%ƹv]:"�h���O�2����ك�E�V��щ�+'��K�niA�����.�G%����fJ���֦���!��7g�unu{cI��y��b��ٔ������.�B�;Mi
����+6������t�@ͷY����Ҥ�go"/Qɔo[pn�;HfN��氡z5��H9TL��������k��t�1�q[՚���#���aѴ(5�B�Ք����.�mat���=�M.����Z�k��bZ�ͥC+�e��t��"�zm`���]�5�!ܻi;s�*S��V]��zi�頡�9Fn�����f��&�Au! O7X�j�	d�oQ�Z.��c��Z�Ǫ�B,�4e��m�� ����·zA7E$�͔�Ό���u���ޕb��1W=L��))�Xd��,��v�-�t��<��vz�}�%��S`XXwr�7o<I��Ok�Gr36wm^ҙy@R�l�ŦMysQu7�raW�ຝx�� oj�!z���z���YY������ ��]EWv�F�R��X�D�t�g�s�#n-C �dB�
`GA�	#�Q��F9um0r�ʖ%a�V.�o�R��5�'sє_n�_5&J����	\⋻��*U�e٘(A��un�9c�t��	�v�*޳giD%8ڲl]�L�����n��os�rܺ;�7$b���Y���-.1���S����/4�-�O,U�edޮo��`�o�sR9#jb�:ͺ��VWv>B�ä�d�����Eb��7��h^��XA��)�d�)Cr�B��n�g�j�����8�	I�FVa&�;/5�8����N�ȽB�<�&f�q���b��]�-�jd��s��PO��u�f�D�JA}����Z��0t�mۓy%W8����	�6Vթ�*jm�ʬ��Z�F[��(�3���釆���T�԰ PKH�z��o���^N����r�d;�)��R�����N��Au`.�����>8j��5#m(A����$7M#W9�1��g*D\�v�\f������h]�>Yt�ީ��;�}HX�wf10�2x�I��{t����Mak�
��������1!^���Zp���e���r*;�$�fMꄇhvn�n�N�;Y�Wt�.�BzW���їN���6o9�;)#�I[c)$���
!
 �%W�k��ȯu�p੦HAvZK����Ȝ�u�6{�NJ�צ�wI���P�q�S��:���L���*��p�UT�q�\�*���Er��^�(��Q8�u�̎�D�9�"<�HDNU�j�.y���q�Ã���w:�a���㜊�R�뫃�eU˲9ETEQ2�h��p�f�UP��*���p���Ň��7I��"΁TE�vE:s��D�*��թ%���������2.8�"*"�����E,*'Tr������	Tx�w]K*8U�'KD�8�T��N0��E%j�x�#�S�L��"��ʂɕ�:Nu���E˦�.EUU^u�e���,�ਝ$L�QR��*��ZUDG�s��R�r�9t�'TL(���"���H���h�NUʤ�G�gJL�	DG*����r9(4H+�q�u�pE� R&� UH�w2͍��Wn,[�S7xCۖ�h�m��@ouM��R���N�N��s�n�k3�u��}j�u��w�7��"�`|��R�>�����aw���῞;�©�
�z��&�9�!�x��~q�q0��?;�;O�������z�χ�i����ϼ����@�*zy��_X��B�*Oe:���;�������?������i7hN��{���8;wNӻ���ǯO����c�!븩��E\
o����?8���;�^!�����S��'x���E`��%�����>#
r�����G��eg?}��߻�}C���z��]����އ�s�v��	8�M���|M�	Ӵ��~p�t����u������ x���F��&��}�~q+�qV�Y}��OO�(�n��xz�1{I�Z���oo�b�����}��R����W�����oh;L*���N&�	������S�v�������v�:w���������Wq5�n;���a|O���)V�|n��t.���K�z���b�ȥ?|�����v�t�r�;~x�����O�����O���!�i�C�<��&}qߞp���~;����޺���;����t�@YS��z�ӎ'�*~��sSb:b*c�������y�?�_{���<��?��$�=��;L/�>��t���@�O�����:v�(x����)�s&�	�����:/�C����zݸ����|��$���f>O�q3?DL��1n�VVlw�ܱ��}��{��P|����D~��|QN?��8���n;��?��u���0�oS���S�L/��� ���n!�����7�q��w̦�	�������P$ޡ'���v㷞X8���D�n-�9���ǣ�q���@�������v�&��>u�Ҹyer����q<M�9�:L.������A�aWv|��t��n��|q�C�����|@�'i�{�\��C�>�ں�,���1�L|& LFu�7�W~MF���|L/�nv���M��'���[t���8�<���q���I&�	���q���`�O������0��}��cx�wN����Lۻ𢫶-��������11�?T��>�,�������޸�q����e��O�?���y�0��I��~����^���~��+��N݇�s�v�O�;s�������'gV�M�	ް>���UG�r�������`3��(��.�b�[�:����i|�(������#쉶ӞN��N`��¥<�ޕ�s�u����6go��<���*�[�ΣP��.���&��\'"*T;�e�c2s�N��pp$�ϩQ��w����VBͥ���=�����x��� ?�������I��w�C��7Ͼ~��>8�����y�!�q<M�8����������G�|L.���7Hq?!�e�'��|M�pn��=|�����{u�gWߧ�>xn�>&�������ݏ���twc��~�v|��}w��� ���N�?;~M��s�������lx��qYPg�ُ����x��k�b�[��o�wN�&����N�~BC�2���8���t�<I�w\���7HI�|��C�ז>n��0���9��G� �7;K��v����w�֐�x������9N:x����=�d�	n��;�������6���0���8�קq7��q0�����u)��d��x�!ۿ8�q�cqߝ��7����0����ϝ�������y�[���Q����;�l�3?l�ӏ~�擤=M?������>&�ɮ�=�َ�z����}y�C��A�N<|z@�w�i$<w�X��
x�'~q<q��N����=?������]�U9�O%��>���`�w��x��0������;�'�q����8�]��7>�t�&������^;|M����'$�'�GN'�,{9e7<I�?8�.�1�:����n`ױٵ巼����Gum��pzR���o���탈~q��?y����|L.��:���7����޹��I�!'��q���?����> t���z���=��i��.��>}Y���Z�� ^��ʮ�K{�b>���{���q7:��p�oY�]���P�?;}x��se7�O��y�������7���v�����0��p���#z����@QM���9�L/S�^�7�~%g��7۷�u��1
c$8��N'�Pw�!���_�0��N��u�n!���|��;Wt�w{��c��SO���Վ�x���;<��bM�ߞp�ۿ��;���x���?G���}���M�^8g^^�]a��N�v�C�z~�})���^���?'��O��C�?'}O�aw�~w��|��C��;�,z��N�㏮'��C���> z�o�/�r�#�
�>T�Z�}������ݹ���I&Wxl�l�?i��I>�C�q@$�xv��_s(ۺ�c�eޛ�<�$�8���ͽ���-����#��~���`��{uIr����li6�7:j:C���44Z�q���,����3��������"��������~��u�}C���?9�t��i�aC���w���8������˧�C�^'ϰ'�v�]���������1��Wo�q���9�^�w���^jJ*ף�S����5Q����Ԝ}��N��_Sq4�܅��J﩯�=�پ!�0����?���>��|=�8���w�N&�	?;|x��s��!?��S��C�𽏾�v:�\�	�;ⓈS��Ɉ��#ЅO�;^������� �\�G��;}w�����c�H}O�8�s���ӼC��s�A��
���߽c���q��xuX�T>��`=Iɧ�=	?�w��%a�w�x��|�>�i��:�
o]�˧z�w}pq���r��������x�$���y��Sz��}�I�'���'��`:C��;���[�|L.���}�Hq?��_P�&s���������������+�8�wV��Aw�ǎRM�v�N���M����t�����8�q?<�����i����v��"��~yc�ym��+���t����}��7�y���ﴪ�J9{�&~����~��n���aO��7&��8��V8��M��un���;?=���;��t�}|M�>�!ӷ���!��/#v�����ݞ�}��;q��Y��{+^�o��(��LL�?	�gzy���o�I�����v�7�'��zۉ��������v���ێ�۵�7����0���?�]�a|C� �!�<C�����|;L.��P�{��N�;ю�07��vt�����t�\�d�G�8�x��8���8�!����{���h�����>�~v���$>��ڸ��7�����w�]!�4�����>w�x�$�w;�c�L@����N�w齦{���ُ�`�T�|q�����$?!�q>w�7����O���<O������M�?��}=��<q �����{|@�$�q��I��z�>�N�� O|��s�	��Z�s��}7u����7h&�{�����"�7n�x��q_�o�A�ι�:�;�#״�'����u��=���8�o�+�Ԝ{�����{���={~�������0~�7��٩U�/���ډ�o*�*��"n�p�xm��i}_�j�Y*�*��&�~���[�N�^Y��5e��r&�ZQ���R/Y}j�6�+�n^J��T���{��ʀ\�(�)��b�`[���폸+�\y�w�}��������_!��8��һ�w�F� I?��n~��n3���]�gv��7I�BO�;<�����p)�w�:��v�8�����z���<��{��c�t�}���?�"h����ک�������/|&>����Q���Ѿ<wi��>Q��~O㿓�Ք�0��N�Gi�C���w��=C�wÖ�|C�+�����t��Hz�����<v�o�z�����D�Gg�bJ�gPQ����Jɔ��@���r�7�����M:q���������;I���t���*X�o�q��|:�L�����g�c�I�awG~p?;�?��8��ĩ�t������Td��2��3}:�gb��j�w�zɿ�?�wϾsx�i��ۉ��=�'�_�n��M�H��o�`�	4���=N�;H�C��Sz��m���]+�M��v|����bC���={��b���Y���M����5~�J�T�����w��x���9���8��Rw������q��x����s�y�/�_z믬9� i�z���:nn\�4+2��h�Z����ڝo�������$Ud���{��r��#y����s"��h�#铂'{:�tM���#�y�OX{��!�^>5vy�a�w��S�X�7_�xeo�J�S��>9���Wۼ��w�E�7�q�{���g�֋t�׃��xJ�W�
�pS���}N���9q�f'����_3͗j�^n�>��t��*����3�8}����4�@�ܵ0WE��� =Unσjq�O���/=�����IX������~��>~��LJ�]lB�r����� X���o`e(����G����L��+���|�����F���YVJ�:�����I�f��2����>-��)r+E�T��{a�n���;1�8��,+��Y�������ǅ%�Kޥ�h�Ư�Lg7#A�7�ʽ��=b6v�&!�ܧ1�[T��9���� \��]��2w}��*��oq��E�?���ق��W��B����C����5U��tx�c���Zn	8��ū3=�� )� �[�C�EdKGJ���&�,����h����\w6:��W�޶�i1����>�Od]԰!I~�X]�jb�c���i���$t�K<�3e�r��;�=Q��wv��J���V}��Bg�R�4#�v�he�m�6��y~_C���2��ެ�ӠEDy�-��s&`!��۬��%���D$*,�̮���!��.�W�-o���
����w�/��
�1:��S�31ov�f�T &�)3 )w �Gi��H�N��=Q�v�.w��*�.CC�o�%h��s[f��ΫPt7�}s'"왷�qD !� �h���wI���K3)���!h��׶紊S�+��[P����u�/۠1�3Н?�u,)�r{|�b9��֌uI��n�y�^��p�B�\=7�'¼F��j��!a�J�O�$�n�ZT��9�z�����uh����5�Ѷ�b���HںTz^e��r��4%R�t`�K�/1:�5�HƔ�*֜����;��5�yW��V�h��k=�E�I�^�}�����F��Үn�w�^�^��/T�����ک꼈�ϖ?��+�]-W����S�� �������$nn�+z�D��X�"���7�}X'3�a�q�>�b�}�N����\�c�v.��x���e;�����w�p�u[�CK���DX{�k=eX���ԥ�D�Xf�=�ѥ�#x?�Q;z^025Tk�cό�'6R+�Q�c����5���6<�r�L���,(W�ZY�R���L�ۈ�r3]�1�:՟g>�! ���l�b^̜�;ŵ)Y����UE^J�ϭ,w]0�������r�߱�2%��-�e�	Uk#��v5Q�������(�T+0�m�
�� 9�\:V��sԈR�s��;��
'q �H}zyUFV��T���2���TvCw/+��OܠS�ZY�;-e}��(s!����ݟ��|T�G�18׭����19.~���Oj�;f���R�J]�XDp�n����7�S؈�;0�]�PPq8M}q�d��:��[6�1+��!�;��G�a�L�:�m�����zt2[̩Us��nk���j�����@��o��kVh�YK��O7�lw��3�t2�Xٴ��i"s>'r�/-啕Dw����w+��f�l��.�V#��A���wY}�v�ܦ*Z/���+�#�(7d	��م�љB6���V��L\��?�����Z�ő\]�h�g�0����]�@��h�2çM����g�dP�Oδ+���<k�!h�Iړ��c���uG�uj2\�S���Z�[I����PhvV_�yL��n*oU9��k�S5�N�%�j����8�(;S���\���w?\Bah.�������V���ʳ¼�ݳ��E[qP+]Oa�w�����Ӫ_
����m�lxJg�4�'F\��灤��O}^�B)֮��l�]<ή�R3�9�k]����aM��J��j���kDR^d���c�a��X���^�9��n�X��TȊ�6��W� 9:�/�p��ۭ]H5b�ʞ�m{�w�ݩ���Թ�ڹ���sz5	�GM)�����z���p<�ȫv%nd�7��Wwb�cL����#¦�D��k�*��ݭ��PU;_i����a��ܯ4�&��J8t��.�$��B2pB�=uP�t5�%|e��\0r5t�g��/'�6�+
�e�aL�)����T���<�o���ڲ�G��Wr��mn'<.xfSY^��V	�j�(���.0aC�m*v��j[7S�T��4�nv
wDs�;Gz	�B�Hn�ܾ֖���v���=���-urz�'_:���X�IOD�������%;ːq�\)��cʓ���;�V���)H�ܧ��Eg�t�����L�&��hQc]-�����q\sw�<��v-ۓ9KN)��Lo'd>��n)�< ��U���{8��qꎘ|	
`K#�&r'M�=0��ȇԦ.={����[¦aK7݁p'N��Ŭ��s@v���xv��Y�o�I�T�!8$ӳ4��=���<�w�o����雜΁C4�+�$ �;
��g�NM�9�\*�`�|�Y
�֜T����$*����j7D�6�A�hGz�1�*V��u��Q���[�z=���tPiLZ��[���ggmz+���=+�νwt�yW�B{NO�����V�ǡ��n���7���|�I��Gy(ێ�q�M��F�t�fB�ٙ)����@W�K+��[#ffw��7k9��-��٦���F�D
��֍e\�cf�lŞ�7N�pcg0��M��t�;\��[P�������+��\&���3�.�P��j,pOn�:�C8mU�['�pǖ����Gp�R�¼��.&"���/�D�Vm�!��)د`�V��ݭ�-J�W\raY`�v�hs���b�n��]����#�cc���2�e���D����/#�9j���Es{�FH���M��.{��gQ�Nw7�@���ձ�oY�����s}���{���GY��m`�lX��V�U|�
k0�6z��땺�Y�#�5+,�f�7p��w޽����q��˯0��rϑ�mW=g��
˫�y���::1�v׳�6��c�8�j̗W�}��|������f���@��y�T��*�����`��ٷ]�Cu�=�I��WJ�s�S#�k󾘨����оU]9�9iX��3�ί��aå�5�ʈc�|�㽙�stx���$y�]��C��Ncx[T��9��~F��_F��A�U�ڒ��u��g��y>ڦ!N�r�����'t�C�j�M�"6�MdSt�;�NΣ��9�Z%�*z��5�!�X4U�Ux�Ϝ��s$v�	� r���;{�8�{�3�����Oiuo�?�q�m:�������>�<�X�{���oY��۸tY���[�84�g���rAb�����
%*�B7�]� A���]6�O=2��_��Ht^_���5�jD�vy�B�:up�e��!"��`v/CW�iC�5(㥪�sY�2d^պ3G����`�m��r�j���_(���{��v�:�tY����#{f9gS���FH �"pp��L�u�����0�s���ix:V���n�����*���P��mk��;R�����e�M������_U�y��^a�����k�4�Kc6�*���fb�{�ShT�B�1�
\3N������T9��mn�����k�ݑ�w�/E�No��90�Ca_\�ϗ���%���^����2����T���K��I������ߦ�e����0j��OU~?{溇�� �j�yI����T�:��hA����sn6U�9��dN�/
��1&�*cx���񷏊��@�쯓cn�M�s���O@�Ͻ$+�� �~�c4�u���YY��R{��{�Yj8t�q����@쬱s�g��3=5�k�?/M�J�-; �bY��6���q�GWP�S2�[7��$q<��L	���� z��gZ>��t芭o�z3��5�䬄�����wЍ8��퀢4F!ݩ��l������M��'�m)p4��~
�{����3���{�tk����S�)��1¤��?�����\�a1wOV}fŠ�^͢�o��4�`r�f��Q@q/uxpu�6O��|��մ9DG\(���WVj�t��zV4l ��Ӏ�,���H��"�nU�D�B����ۧ:�����-�]���7�λ|�Ұ���]�ЖIB,d�:��?=�nn�F���]Z�uWSc6%Y}HU���Ɍf�|��E��I�ݾ�����
`:,@.���]ւ	����]|N�нե�`�Zg_fs�8�%UA����Q�x��η��{�����>}64��o�b9&�J��!�H�J�^�*�t��V��N��l!kj�;��ND��nd�{�ZD7p	��8��1��^ͫ�Hc��E�l_j����#iKR���uv�F8&Փ�Ѧ��#9Z��|�����w�WW�0+[���u��˩�]�������ix#Rj�R�u)Ѣ���L,W�j�5U��P�u��f�رCs�M��j�%E��|9ՋF���l�A+.P��g ���$�8E��sW�p灾wj�������s�mK�J\��{u���qw��8rm�����,`��Hi�r/	�ذP%�Y�\z_
6잔��$f�̖�ېk�}��2b�w�]�Ff^u����[R��#Νw�*�b\�w%փ0R |�� *ȱ�W3�Qk%U�6���=�igj���r�N��Ѣ���oU_�t���s��!g]a��Ø2��agT���kVk:�)��+�xlnp��m��J�Y�BB.kpLW��4EY�� �I��S�0nX�F� d�H�0�.(�On��)g8X��)�Im]���}o�Y4	�ȚɈ�{C��O4�"���m*�[#n�����4*�^��B��aи�\����yB��M�h4"b�F1�Lt��l o���rj)�)��x$��� ���f����ڭ��c�U9^՚<Re�ֽ�ȰM�񳔗_C7)�W��`�s�r#�&�`V��mgnt�%Dp���J�\��~�AK���~�u&G��-f�ˮ��+v'f�h���5�]+��}��W�(ܨ�j�!��Bd�tr�x�^���j�6�`F��WY��C2p2��Wt�Y+����n�m�A�4�[Bc�&w/�h�\/39�B���.p��N�%s�Z�^]J�8��f`�1�]m�)1����t�c	%��s�s�@��\G�5+t�\���\ M>s㣈fZ[Xi�2_�	
�+Mϵ��uzU�hM���m��|I1�fɣ��5g)TS[��+��6"9�a6��*2���l��,���r���wV*�9܏E�!p �S��ß3�`:5ŏ-oM@�,��CS2�>ӷ�6b9X�#hT�3Hc�z)�p�9ݨ�Մt����SϏ�a[����1:W��%�i���)\�cM(fU�*�A=K�Eœ��	��f��`�]�N��*��"�3r�,��Jh�P�r���Mb��u����1,�,S��s����q�צ��Z�wS�>]�:���m��X)�@P�~���XS�IR�":�
8p��IdZ�E�P���u�s�e ^��"��B(�uc�qW.p�2��ܥ� ��������,N갩S�����:�x"�:�(�W\�ԹȏQ�B�#�WuB�:r�
(�"�zByXV�Ǐ�e]�*tȈ��6�
�8�OOH��G)�C$����)*��8�����J�"�+"�.T�����9��B�P�2�)�B��TUM�r�㋸�.��;H�2YUʪǌ��bG����2���QE�UJY"�!Wr4�dt�N0���t��Dks��9AuCR�+�ȇ�ypr�ZF�S��%�8�EC���\:�2��J�n�rs����N�UI��h��@]6�tE�p5i��}c�3���d���e2�|�.6�^.��z��_f><���).o5 ��SR#9����5o+�z�n��Fa��wd^?_��,8��9���C(G4:�
P����Q����6Qݲe�#�Ї.p+��+�4�Ȇ�^V@n�Q4�2Koe]�����o#{�SWG@�(���\_7��S�R�C���'e'�l#"R���P���|�/"���̞�DS6��͞�?�֐�c�8M}pU�Hst&�Y:����t��x���[v�ۛc�*D_��AQ��j|+�ٓ�]�믺S�+�a�0d�'C�ϟnT���1���J�:N�!��T��v��Z*w�"�{+����m��n��;������Ҙ�H|mm��"�8m�3���j4�'2��p?��㊟����]��*�}�Z"��*���<D��;2Bܚ�2o[��l�<S�J��ٗp�����,�ʦGdV\#���>�:�hS��ƹ��ݗļi!ҥ���g�1So�je���.���/yI��m�5y���8G[�<;��Z��A�f�Bc���:��bf�N��!�ڬ�~�T)�K��#y���&U�i��n��:X��7fz\�E�#o��-3�V�!��2��TF��=�b
r���Z���<�N��2φ��&i=����Byrv���P�	�l��Dm5��(L�V:�;��:�Ez���S���{�i�᪶�kR�����U�U��W��Q76�6v:k��e����	C#MDW�m�=x�9�"P�����o��P�Es]a�9A�z�gwp
wNՐs��k�_�pve��*�W�:W�9�8�7����/U𪍥��n�+�Ep�C����#�W��;���Mxefs;Q��V9���NJhT��CK:+{IHp����W�v�RJ���dɎ��L����u�2���:5�����d���Q�����do7p��-ۓ��>�;�^������#r�'�Y�]ް�n��0oU��+�y'<����{�<�}�ʞ��QB۷&AZ���f�`���f�����K���(�Q�����9��o�z�L��1��FT�fᨔ�0�Ԧ,<x�N� ��5�,�j2u��g����\mt��P������&��䞶!r�É鍛��/m?/��Z�['r◺�;���=x:��(FB��gh��l�t�Cj�Ѽ��������rتҠ��?۫�zAl���Щ�]	/+pDW�)P��إJ�Ru��2<��[ZOG�%�Fe�z��@��uL��%�u�����WH�z�X�!f-���ܐ�[,�z�F�y�_l�(W!��+2���4I��X���Ζ+{���v�&U�ޒ.y�57.�ƅϤZ�n�L�]L���7���P��m��:d�����V�E�Z�Ou�����t_c��ʼ�~��B�������g��}�M�ޣ2�9iY!P�Èw��Pf*sns���:��?B�ٙ6�����ys0��
�O(�p[���)���k��<�5
�M�M���ٗ����7ͼ(@�����9�&�V$�ڒ�c1�:��.�o�^߭��FsH��iO
��z��_��#[�9>̇��T���7�-:�Ҕq�!��z�;���!����x�X��{v ��0wG�{#����>滔e>�z�
V�E���cEh�*�C�<%
˪�@W�.;1mƔ������o�_&�?u1�'뫁_E�~��e؝�t�#�9�|��6+���{J�m#Lk��]�j/P�����.#�\���큒��n�`��g�y�Zݰ�_f+A��/ݢ����7޵S���[o��?8����D�2%P���qzЃ0��}����޽��Q����EL=�zڵ}hz<��`穼};�z��^_Y�b��W���
^��c�E���7����e�U���j�tٜ~�蹐_ڈVU'����w;(���Y}ܴn��&1!}h8UŮKu�ס���>C�%:�7%�ʂ��s3v�7����V��*��o�+��t8Ԝ%ֿ�i���˾�{e}xҍn%m����S���V�o�\w����_}��U\�<���r����Ws�-@U����Hq��S������<���(:�*�a���-�%�v2}�Ѓ�]?�u�V�z�B8���ߒ�K�wܳ
1�ܞ�sĽ��&��]��8�4��
fv�ǰ�A�Y�D����蔲�؋�]�yF:/���q}֟"�#	8�[nr)�Hkt�MĽvmٺ�m��,F/�D$+�5r+�w7n�����!R��Y;xdb�0�����֚���2���;uޚ �U붇9�q�Ue�P%��fN� Vũ��+��ݐ��"V����ٸr��kBw 5�y\��m��H������{h�y�iK��_?I��}w�~2��=*�FjV�Tbu�"�2�sȾ�V{]��lJpF� XT�B���#�m�ʿ����<tG,���p�v���K�괹��=P�<�!���u	�$v�Gg�����!v�>�V�{Vu_�� �Q�i7H��F���<��ݘ8\��pew�TK}e}Y�&��i�J�?<��;�k/Ge=#�v�ASt �s�P�6w�肥o%㫹ӖuVmFc�L�G\�1��q
��Qw��?;��v�y�L,�q��s��Vt����h�C]�9A����.G�����E��?�ۗw�#�<5�h����Zg��2$u�ڑ��}}]Vjƫ1sHt)�AC�>��g&�������7��$�!骜n�zr�� 9�"Grr��޲��V��y6��Cͦ�����\#N'��`/�F!ݰ�|f�ӑX��4WK}oʭS�'�<��z�1{�رX��]�^��UΣ"9T�9���r��aK�]f���sJv7�O�|R̃��K,K�ʊ�8Bo�U��<uV_O��>����<����7�g��j�w�/�_���ON�T� �� :�Uí*�R��}uJ)�3ϸy^Q���;9�ͤ#Xz."��*,,�X��9i[u?r�{�B���}���5w��.����f>���}p�:�-�^��`}���Q�k�X#�:�t4��՛b���!K�煿����;���	�&�A� ��	��fkg)V�N�*U�E79���<oa<��� gu*bN�h�F��2���△#�<
�Kw�1�n<,�xfqm->��.�Y�ר֋j�o8����^%-�YB���)!ҷQ��fbk{nN@��(��2A����n�VP�����z�QE=}K	�-�}�g.��p�U׼jV|T[��q����HOq���Ё
K�bb�.���&l��^�����,c��{��I��s���f�\�}\gV4���.ޗ�e�-��2~����>����TSIBC�W��!\'�p���h\�Ƶ.��x�m)��_O�2��z�V������7���Oa�};��w].	w�1�����.�[d �i���Y�'�#��=X���Oʃ:$�G3VYJci����5�nq
�Si��g���
�7|��R���q�+=�8�#�V��E��Ÿ�l�1�����%ݮzV�8��������m֌��s�ߒ����������Z�w��>F�#��r6�����j�#MDa�p���A����{��q�z/j>���JQ�&����f�	ui����(�1�W����
s�ߎ�8T��~l�������<��1�1���� �3�:��4�G�vxJ�J�/��ğhf���u��Ѻ��o}-�V�w��T�+���;H��䫼X�x:�_N@���P+�9�JGLs�,d�߸�do�ʡ��[�RC��lt�e!Q�J�_W��z�%�N>fB��f��~����
7�A�|
�ݹ3����,hVw��_s�����)��y^93!�(�����^�
��UJ���&����ط�����8Q1�E����B���ar��ܬ1��h��tioVҤ��N[�"x�krt�y�qf��{h3�j+�+��䣴��1�Ɏ[��5,����dy�aT��:��(v?}�����e�"��SОnL�W�,9��p�.0�D$��R��:��T���3�6ξmL9%��ӽOI���X6[hy��<=�hRmQ����x���W1��UЋ����엎�c�$�
v���f�`�Ъ�m9+M�]��}�y�.[�KIdla.7��t]%�E\�u�,j�`����O�dz��v��ǡ;��ttI|�{p.J4�.>��ʗJj���5��Ds^̵1��-�_iy�T��q�j VVJX��Z|���d�{��Ր����հ�T�f|U�L��2�n;���rO>�o82��'O-�H�O��9�ޞׁߘ�����U3|�	��d:�ه!� B�[���`��{��ȫF��xVTѷ����V:*�4��j}�� ��ń2�7U��k/
��ME���1�Z1��]#�4ͮ���8�1N�xՎu�W����p��؍;��=�����^�<��W��R����p�kE�U�����e���=���oT�o2���^i������H��}�`�^�;-��q����X$ӛ���
� �&��c��iW�״��~糳]��W�+C��0�ݠ��r��$��U��>�V�s�\�s �_1�j����w�D]�J۔Ҭ�vŀ���5����
��wܾ�dǖ��r������H*~������V�����t����E�)�.�N�	�ע�q��$o��T�b�]}x��P�k��g5��;ݝ�" ��j�3K�9�7z�1e��UO�o��^��U���`�(]�텧�͛�8O�E.D��`��{|�7P�r�1�

vn#Y� �1'J�8�-ݓ�U�|�ǉb�h<�:!˃��B�tD�/FBt�Hv:�$l�l������8��Ϻ�fS�Rx /�f�4jf6�͎"w)��4,���&�9]�2��s���%��G#�|��톸U����u�C�*�^���S���s��f�ׯ��`f���i����l��	��s���"~HL�J[vlE��h��P���_�r���8q��\���7�=�3R�A�>���F������u�<k���u��u�p����YX�y(��Q��lw@��B�FE�P�A�����˪�������-.Eз�S���ٟ��"[�&N����p�"V��*ڙ;u-�E���aEu�+��|��/<�Ќ+��	ֹ��-#�i>��4p��,y�$u�Ivb|5[=ף�R7�>��
n�����;��J\
�}{����]�
o���gPe:R_=Vx�ɮ�l�S�%;
��_}�}����盋��Y3^�M��$B#6����.�Tf��}!N�r!_Ȭcj�&��{w��.��Y*'>�����*���{�#Z1��U����b�$I=JX%�-]�98:�GZ�����r���[��Wh��ٟ);LNWޤ�݋������y>�v� �Y���q)�NC��!K���	�����:c�-���'�{NUЏ�GX޹F񝵮$�]����:|��nY�fe�&Ru�0]đ��u:�\K<���rP�f3}�x$>Z�]��'i���ţN'�x�`9�ct��Mrzv)���cZ����6� ���Y�ի?����ҭ,򩜇g<��E㑑�������A��5���Dﻪi����:�ӣ���3�#|����ʭC"6�����ʅ��=�e�aU^(���Jt�>�-��C!Q7��o���5�P�ө�|�k4��yWś󹁷�]v!��\6/�@/���s��B����e-�+ �B7�����A�K�[�b�4l;�e��_i�<�8w�ߐ�{V߽[��sx+���C�*�띎j�u�%-W���'+%3>��M���O���;��S��a&�1S&n8]��Ňg��wS��L�n괉�W��WW?�h��:ݻ!x�L���6m��������B�k����H�d���9�}P�:���i��Z�&r5�Ü�h �"D�UX��:/�%�os����A/n&�z������n2���!�_%N�	И(c魛��,��s��\3�Y����4���&3J�zDC:}�jF���=����/"���:`��Sm�v<���Y�F��ݑ�����@�WQ��T�|��U>���4=�
?A]k~��넓��xL�v�˙40��03U�� �{��Z~gI�{�����4�k����t���=.ϏRS�IK^������T�P%L��.�E�fFU2;"��Z��+=���5���7VSu��g�	��}�
����y63��5w�OV+h�����ݬ>�+N�W0����=�S�A.��z����ܑ���]�'B�����x��Ѽ��
�r;���w�w�S���m��h���cҭc� u)��"Y���*�a�ԡ�(=��g�@.�U���x|{*�rd��ԭ�(V�E��ʾC<�׫�ٝ+¥}L���ʷ�X�wm�D��0��3��:�	Ʊ(%bݠ5��U�b�&R4*V��N"���;Mu�a� ͹�W���˜i�F�z�뫾��}����I�W��#1m�Hql�XR�c�2fc�\&���f�µS�]��G�������kS������]X�4VJj���<����p�g�]Zf���iP|��r���s9o%M\yj���7�Sᲇ��Z\!ǉ�O�貦�N�R�ô�
ӳ����*���}��x)n�{V��A����B��}�W�7N]�U�Ogi�0ۏ�GZ+�����s��8����A,��&�J���(\�+�wm<3��u�[ԚN��--�v�4f��|]��IR3�)��bv
�ʸ���������IԨк"M�;���|�l����VQ�xW�������c���b��{���j�r�Z���z��9>T�YiN�A�1R�U9��t�{/Cs�ש	�ͬ75+�Jl����Sޞ9�L�AG�B���$��B�.5����oj̬�f��s��x-���M񱷠�V��VJ��j�T���Wk	N�R.�1�9'o����tBU��*T%�9�N���5k�u��=�f�3�.�r�k�,�M��/�Ҍ�&-��>�r�ե��I�w��3|������G��\�,�ñܻ�cx�םG�O���y� �]+i�g㯖�����ƥͣ�{�,&��U�p�#M��(۬ˣ g�K��~��\Gu^p�rv��o��:��k��K��L�ιm>xQ�*$ٻuj�s���u#�j�\n�'�@�Uj囄���1s*�3@gTX����C����U�C�F{2t���ۍ�[�є� ��M�R�c"��LͶr�r��K����S�\h�{�Je�j6�1�c����QP�
��.��M^7v�):WZ�X���:����s��K�HYW)"gmr*�ξ����z�N���lp��6���� �0�ա2��jE*��D�]�Y6Q�59ݬ�:�JCGn�BX�{��0TѪ�e�����yIL�P,�����]�ݪђ%���\�
�z���Ml�'_4���h�nYZS�,����6w���+GS�jcG7��*Y�G �1��Wdb��{��S��s�ɭ�6�����˛aM�L"���pIV$`ᠤ�Cϐ��u@z&9
Z�CZ��'-�-�!��"�݇k�]=�ki�N�`��V�M혌��r>k���\������T��(���hH��?x�zy��U��Ox�����̂ꋣY�l̦�w>?-��b�u�q�y՝SX���\d:aK-'dP46�y�J�#�6�闱����^�tWϕu��M��Z(�  �%���]rF��"�s���8�2J�edDt�Q ��p�ܹ�[�B\�������M$��=r��̱,�b��\�QQ37\.s�ۓ�u�qb.:�YjS���kD���mu�4\su�'N��4u��J�	Ra19�UjV�&X�T �f(ujej&Ҭ��Jb�$'���%b�'N�]\���V���E�ȱ#)IN@�N]2͐j�a�]��*j�db�f�JuhHdXA�9ƺ�.N��R�^<^3I$�9bU�,@�n�9EE3�D�0�V�Y���YG�9,���!
�L3�����ӑDQ�H���)K%-�rsf
˚(�u1"DT�F�dB�L���\�B�C$���
�RE
��T!��r8�H�"�^�y1~�|���)-EuѺh�pu�u;�x2:����?W�#�(p��Z�.�S{���#�Wf�fuN3t��_}U_W����S�z{��ı�����|�&�r0ϩ
����Q;<,���]�k��G�;���\mΕ���z�e�lE0g{�������ے(F
ƕw����V�pW�٣�6���ܬ<�%[H`0X�v#����n�O]??����'{ѷ�M���;a�j��d���������;w���}�P|7�& �R��,�S��S��*��K�='���ϐ�exb��̾�V�����(�I���)�b:a�hvtR�=�l'|�;Γ=ս��z����
�3���<�P��{�J��Z�=5pV=HD���)&�ձ81�t�&(vx���Zl/R�:��o�lB�����F�C�ͧ&+��\ڼ�'2;��'
�lhߩ��8�Y
��&�e�.gH�#����[�u��Q��;z�,w3ӫ�b�gf�-op��Z����8�\Š�9[�2�wr6rC뫾bw�r�b�'+���-HO.ީ���X�;�j�)���f�u�o��Fuߣ1,�뫞ʌ{Z|773s�(�8�dkI��b��򭵡X���F�f��{���5�W`�}K���،жz�5�G�O ��@����e���4��윎S��]A�s�ƻ��)�c(��a�aͷ+���Buh���]�3�WL�/n�`����<�iP*;y'[Y"Z2�}��G�.�&�����D
�$�l�s�x}�����7�����C!��l9�0h@��UEa�D���sn��q�#��V
C��Ks���;\0U\J^}	����J�NR[4������]<��Ǘ2k������X{M:6�zU�<�+S���S�c����Q����%%���ST�SQ�u�:_ڪ�q6vȍ[4xdE3��
v��f��
O�??fVlKF��乂�[��m��I�)��.�NG>τ�k�{9�]6Hؠ�r���[�U[�Em��ڟ���g}��4%�tav�ȕ8��c�1��ڞ��3_W��;]����m��&�5��x�Y=���{3�����Ĕ2"�����s�r�9���ݝn��&þ�3���<��s�KJo�)�����^�o���f��R�Zt�H&i1	Դ�)"ûԣj��t�v�W��d b��`��r눛�d)��j���^|��Ԩ's^ZW8IDww/��xd7L���A�
cU�cHو�j�c����Ф����w�%[  )n��v�=�ڳVڡ�"��ܶ��tZ8���rx7����Etsڱ(k3�iP�H���j��wm��'v58� ���'fb��w1&(��Bލ�l�o%�.ήY{�EoUF�l�a��#VV�L�1�}�G���U��'��k�Lz3�����ߎ��Hs3���x;�,_��B�U}ٓ�)Þ����������^mC%nA���N�	��#>}Bzm���w�����G�d>�m��x'E�hi�}ʪ���v�q�;�t>���9�7^��A���/Nh&�V7ٓ	�=ם[�_T'D�ن w ���U�7@��p�X;���ٸs��B2-��w�����ǹ�f@Vݵ1�D�i��uЩ'�#жϟ������8�7�D��*������G��%��yP���O��.E����c�Eሿ�1���[Bv{{�GW�W����3�	���$a��-܁���8��"��'ljN��}�[.s<��yoZ��qG[�c�J��|�H��.��N\��݄'�_��\��/E�q�(p��h̷���q<���-iPl8]�����x◓��T���7Z�����DX��e�m�?y�n<N���f���7>�j��;�w������4F!ݰ�|g#� ���;�o;��F�����P��SB��+`kj����C8��9���a�d���p������ϔy��w[ �qx��P�y����	�qj�lN�����q_QX̧	Y�]s�tD�#��Z��菾�Xs�������tWU�[#0�+Vt��B��ZY�Y�p�9�ې��r.�Gs+q�6�#V��bzP�L�.W��ۮ*va!)E�M�
*���W�U��<��_��4�e�BS[�ӑ���մ:�==H�5r�����J�1ON�T� ������^Md��8}'E%�79�К���~:ը9���]L
�
��=ջ{TS4�N�"����9�l���
�|{�g%��������b%;�8�i��aw��	Tv�����m��F]<R絥�WL�b�"���j	p���t��&a�n�^��e֚�Y�y�|Σ�����Dsx��Ѿ=>j�G���ྍ��Ԯ.F�� kW[����g���>�T8,�=ە7��X��TkF:T�8����^'�|��M5���5��vV�\�u�ܰ7�2�C����V�
!�؀��U9�<�fE���B	�?��E�i>�Ht�}��ݣ��g�<�a�PS��Ju����Iհ��f�Mμ]����b^ӑG]�Дѭ�x�\b�ͫRcМ�@��X��vׅ4U�+��\>m�@Mv�ؚ��+���.b/C�����b|,<词���bos0��Y�Tzl�����U2���oZ����m��Dw8�{j�vFG^WV+}��^��<mL�^pz��q*=7��~F&��������}2��^�g��!���J��u�Z� �ށ�M(W����@=�^M�fTI��. "8;�2a�nI,�]=]���h�a�@S{\Sނ];��Y]��Z�ۣ��<��w�w�5���X<� ����eo[�R�"����=U�ZǦ�={/6���#�����q�p�����RY3SM�5N�������s��Y����r�����S~>Ŵ�����k���_�YG�1�w��������elWꜞ�(7��=�ܭ�T<T��.��F�)y�x^�֟-(;[�'�S<�N��}��w���|��K>��I�X�*wr���|�IZ<�Qdr��[�֚���6OA�XӔ���cp����o*�8��H����.�.Y��{̄y6h"V�cs�L>|��cJ���TҰ`��S���)��I�������j`NH��w���h�sNJ��}!+�n"��	����j5���J��[t����x�U�'c+���պ<��ǝ����l*�(yI~v֓��y6t����\�i�IG`x��K\�':�J�]
}�'��!"��JV���*�|EZμ`Qo{�i.�OAʙ|�ι�fi'�:�3mЊu8�ct2ؠ�2w�1�q��#����\�ɬ���|���:��J�%�K&����5RỶE�阴U��lVΞ58Ԯhn�\��LB{ҲO+{�)b�&��AvfT��9<Kv�H����t��Gvca;m#���s�I��WtT,�Qe�ܬ5r1Ѯ�v��q�k���]�Vwħ'"V.!�n�VA�Ob�cV!��#ٕ�����a���6_D[�Z���+�
��Nk�P��N;���v[��iE��PZr=bټ�Y�v��G�)f:�$!5$]e0DfY�Πf��\%N��%]�6{�)v�X�w�FX�3�w<v���o�҉�R{8�݋��Sʣ�qS궴t[Aq����vRܵD�O;ӱ:R3���͸��K�-��ޜ���d�gy#��$�J�NԎ;HX{M�b��������Ǐ�a�%�ގ|y��u����_�����':⚾��X��2vQ�R�C^��uWr����5���e����ڱ�O�Ju~�o��!�ĵ�+d~+��[�6Am+㋝�\��ݗ��bU�fR�[!�{w��]Ӫ��{�u�j�x���oh
(����q�G�������P�>��=tUa�`�xીJ��޿�����oZ�J��U���*��r{��=������W��g'J٧J�f���h��jo1>x���qh��,:���E+�`�ҁ\b��Rͤ�\\dX�&�W������^N���E�1�7�;'o�p���o��Fsml+eKËh���ʢ>���Y�=��6���N�Y0�D�%�z�u�}ؑ��_su<�N�dJK25��@L���){�������q� �=����g���f=5_K���D�IW
������κ�&iJ��yF��wR�E����{fiv�ħ��M.�����A�a�ǔ(	�h��-��.!��#W0f�&Ů�/�Ί�V����n	�e�������#K�)C�2�E�w>��-��W���������x�vf̣��=6���5����O@x&�銃��u�k��5�e.DX�7y���`i� �F��^oWa[��t|2�b�N��RgZ?jǋM��x���n"�J�WCc9���	ҎZ�}���}�X��T���2=��w�5��!�I���];�0M}�'���-�:W�����Z��x��<u渽��cWF�6�Au*.5��Ol\�y����ɩ�5]�4���3Wun '���ͭ�o��r��j.'��C�1���HGE���|���JPOS�9�+h.;G��n�F�\oDinq���	PS���co3���S=���~^A�r��m��<����~���,��;)�\�����C�wZj�c�jp��^�J<�u��T�_5x5A��H�W^V�:>�<ҹ��>m5���',������R��s3��MT�y��Z2#���F�w�,�^܈}(�&��4�^A�L��W���[g�K���t��l�Ox�u�")�7�-�JZ�`M,��;ogj��ni��/�X�s�i��3���D�qB	�Ϛ/sQ��ժd�'$�\k���h���,D{qb��~��z�1��ۆ���G�r�(�Tgc��k��Yօ�s��q��gL�k\RfŹ�X,��^�E�u6�x'[%w��%P�#KU�meJa{���v�,���r-���A��$�cx��%��k&K�{�;���}�����ﾉX�y�����&�� �T�a*�䮍Bf�Q��N�i"��������ĺ'8��	T&�q;�VB�����(]�Au��K�䳺�3�OF�Y�U��V�!����8���dr��E,`�����̋�B8]���M-+/+��s�yPUʴ���>P�C���2`͆t�5Ź��Pz{)��qO*��q��}�]Z/��|]J��3��^B'm�L�	�`�����D�J�p/�����_\r���#��ێ�i�h�]Z��uۗ�����$󗛹�{e��vc=�4f���QXm��"���f>/XT��pj5g��m�q=��o�V`��c���F���P��K���輋s�b�*����jZk�y�;��9�ʌ�H�E�ƺ���6�+	��ivF���g�-�\'���|�ݔ�f[�S����H����fXe��~�4��;eF��M��bH�G=Q2���^��%m�5�o1�WFe��u�.	N��<�o��H�}�Z�v�n{���cV`����S]ՒH��|�_mL�;�p5����s]X�*��[��pާ�	y��ﾯ�����OHs�����޳`�q	X9_d"�da��m\q�S�e���
ֳRZ�y�+X�B��s[���m@��'�����'����"*���;�Uw9;����;qJ)(�$��9�s̙��M��o�C	-������=o'�+��Ҡ藁#7���D\�MqUj�v�,�mS���|̞Z�9�#	T�%qj����%YEb۹Zqg;Z�.Gm�ujW<�k��}<��
YJ�L#����z�Sy��ͻ;y�>�.q܉Kt�m��u'j���+{��g��3㡝�O��A�����)���3�����XS�|��
�c�r��3V�b�ŏ��P,�2�;p-���*�ލZ�]pU��'7��XE��Y�*��kcSڭnpIlP�w7Vk�A=�U�O��Q��z�tM�퓔�H�zx)��Z�,k�O.���8y�G�t�m^D8�l::o�_h��K7s��$f͂��Z:~v%M(�ud"#�N���:�&ʳ0d��5U\�w���J�Vسvz�� ����5C��N�.��!W�!���5�R�ʖڠ�	e�!PdZ&)MRM�]���f�y]��d��G/o1lT��9
�{Q�y�ع��������I�B�9��!�ٻX��[trS&lZ�����]׫�Wj ��n1OM8#�\ڵ:]w*�'�;F�{�]�����%�eG��]c ��t�۠n]lSh.��r�Q2���ei��B𕪉����
m2ӱY�m��7����6^_T�tB��"E��,։>Z���np#E\��Ĭq�(���!��J�W��;g9�W&c�k�T��ؽk��ĥM&���Τ��[*t�q����i��#kj�ۏ��:�����e�eg �d)m��[i`�v_s�F�ΩF��Q�gqD�a���Ho�qT�R�
&�p�����[	����;X2N����$�b��Z����Z�r�t�
���i&�c��{1��r����v,�~�CI�D�S2eYyLb�[�,j�&s7�ܗݡ��8�Z��Mb[��vh9��;lrX�`ɔv�к��+y����Kr�m=��}
Q�[�4�G5���B�F�'���훦p���R�AG\9��fw�إ`j�I�
��9�q���)�D;UQ��@��F�[l��M�%s3l'S{�|1�3��څ�W�-9O*�����c�s�kS�2�K������;3aM�XC��Y���W2�H��8�wٙO�.U��u��f��A��j��V�.=��d�HMY��Z8� �7kN�R����ZW�3���/�Xw����u�R��[ұq�1ͺ��s��+�}(�d�@�Wghѭ 1΃��lnM����� �֋�j%p��ٷ�+��-gOB0
]α����)t̳�Ot�6�E�v*�DM*���mM�$��ٿŷ&�Q���0tm��&u��N�<�)H�_:�^GWx����ϱ
lZݶ�z/�.J�]�5ȅ2��^"��gTc.��5�1m((��|�U@p��R��=����r���.#5 V��S	a6�t�
�Qc���^:�vy���ki$�����ے���=�����gx�����ݜ���(�7�9Yh\}�x��̹�Atmt�&�:�xƳd�M:�>v�]����
�7��t���W��+��禅������=nj]IPź���Gk�
�딍��&�8��Y#�ͭ�l�g%G�2�]��.�u1[;w�fs�f�7#p*M*;J�� u��z24`���}���ٙ-Z6�yYts��%���z�cЬU�i���^��~��h]�\b���6yHG6�N�U�<�9j�����6ޅ��6���Ąy�)��������n�*b������Zs	�ö��v�����C(�j�>��EV�p��q��E$f*�,в�XEE���0��h�I$Q�'��*i�54I9EjTP^W8�q�ErI%�0�ub9	*ըQ� �Z ��F�Jz���VA�u+RCfX���t������dd�i.�b*R)E�-i�:�&�IQdd�!�aRJ�)YԵ#��YhjYFDZm��)Z�\e@��TW9��-=s��Z�Y*�SY�ԣ�:����HYij�隦t�D�U�J�̭Yr"�2K9&V�*��4RK@�6��]ĺs3�˜ʔ�8U�+��*�4���tܦY��
-.��el��R;���4��P+�iHU�R��e\��"8���QR���'H�-PB�!�!A�UVJVȃ�.܊j�%$�1�-�ÂZX�Z�T���ĭ�+:��s��M|v��mϗw�����1׷����e�L�}���tj����p���A�i�6o��<��(�:�M= I���}��D�$���Z��F��q��I�{MI��NJ9�5;�՚2U[��9�9�.�:�<���d2�oc�k���b��˪޳n��e��b��"����j�{�G>Rq������v�}YFoV�OQ���7�S�2��[=��o�����w�j�q;�Ր�������]��|�-�����6����̙���3TID�d~�����&��Oa����G�;`r�E�_kMuh�0��\ި�Y׊���nyr������;~-�gP�~�"v����0�k�|�WkYFZ�ݐ���L�ie&�&`+��GE+�E(�1�[)8궢�Mp��<a7��)�6�$����G�7ҭ�ת���v�8﹬�0rc���;�X�q�w5����i(��.ϡ�uä�$㣟L���� %p�;¬�۵+.���e��/3QXMt@L���O��R���~�;k2&�wi�#��q\���ҦmＰ������=y�ûm�R�#�^/U�ea� ��g41�sP�C�w��Q§��mǘҧ�W�u]��{ɞ��V���4�o�5կ���.˥�X��v3�Hl��k��T�(��\����}�Dp���8�kzyV�c{��\�~�wzS1���sw�{؝��!��2��$��[�nBs��AJ�	ՙ�v�2�$�[K=��A8�䳸��Ѭ��[3]��w>�4}~͈e.^mv�wBԑ�6�%�����y�'�sO��� 3�!��g� Z7��'��I�4�W���1qF�?����ʩe�+��O\N�Q�{,�:�ܣ�i]n��������њ��H��Em�Qw*1�:�j��}\N�����e*����;w�ҫ�=���Ο>�+��1�E��J�'���pq뒬L�`3t�wn����tAO�V�\v�)��u�����#=�]�{Ė��q5+|�{�޶���g�.4�RJ{��{b���W5�j��b͑��N���G$c:�o'7�=�kz�=]�A8�%����)E�Z�x@}�s��yQ=�BWf1�n��7Tx�B%X�Vr�F��c��x�:�{ϙ��G�|�*�k�K۠02��{xr�KV�10/`��8�2�W��Y�����xx�Xk"��&��4��T�����I�Z�=�Ж��V>wK�ܢvdO��.���U�}�g3�������^��9��m5�ْ�o}���$�s�u\H�#2�v[M�^�� �E}e���]���"y=�ң?w��q�~��s��K��K�M����U���Zgԙ����&>y%6����|�C��mL3Ŀu>k|�����J��I鿚/r5��|����� �6�ک%o"��\�B�T�t�ELrW���죹���Mi�P��GH��ZƐ��E,��=�k���]+Ȍ���#� �3�K�Å=�L
�l-�w��i�
;�NW�2�3o"��|�`�z*S�2��٘�IQ����1�T&R����O
iz[�������C�W��&��N�1�����u]�=.���͸�޼|5�ZY�*���b�-�(�3#@��w�ϓ~O���W��ŗq���__.�_^�if<.�@��*>Ϭz�� �<}�9e�a�7�բ��C2���Q��]���,�{]G���[��4��R�mr�9I�`��/:�5]��`�KC����Ce��|�qlzwI]�f���J�`#˛rgu�=���۝����j�}�q�}G�������ҽv�1�/��+��[���:����j���.gRo���tʧ�0�Bz��&�8�k��~��j�
�
:>�;���Y��� ��I����8������O-"�V���{���NE,�*儓�<떵8�W�5Z4�#Ins�P��6��G��z�W�T��{�_7��֚�p�z�{k��O?�}��N���Ϡr��[�֚�ͅ�z��9&kf�kD���� �5�B�	E+f�8�gc�z����H��2�N��G�d������!t����Pt(Ϣ�
�댮W[.��1OlY�ݭ��b+_�e��$�]��'B�	GGa���	�g�u�f�n�@䮗�t��3���M,���5��6�_N�tk�ve�90��v�o_�%��'K���4�OL���P>:sT.�k����ې�m0�](0�ֽw��0S̳���Ԉ��&2 �&���E��8t����b7B�a%�:�(�cy�BN�����=t���{��_as��kG�,�V-�]Inoit�Uuj������=�\'	�u��R��;��L��b�����>����1v�Sؑ���o,Ȕwp��9�Ob^�Y�p��ʹ�&w�s`eH�B�m��m�tfe⿄r��")vާ���';�ٷ�&a�݀+N�S-�a��&�b��3=��Q�R�ފ�\�
�*�AZgb�Tj��n̎�眜%��39[r=b��Ͷ�bW��^���3Kε.��R{7�U[�B����uC�w��|�Ȼ�Ipb��L��in��r�d?��Śn˥[KԔ㣸�!��}GP�K:��:�f��}ډo��x��QX�����������g~,ּ�p��U����{�w�_k��`��v1lb�1��N�����m���Q�t4z�[�棎���
ὕ�2z��Uc�(�p9��o+����̪5%�Ȧ���Z޿����a+g�)E�[�QcJ�}�)?=Z�wh[n�G�.�������FP��Y���loh�N�K\L�uҦ�V��I��R�
�pd�� �7}٫�l��^GnGX�G}z5�[����J�R}��i�C�^�P���/\����`{�����Yu���=�r��S�(ّ
��諭���gezzVog����sa�o���/�9�iX'B���1rk\����]d���u*�>Y��|�Q�M��X�'�Ϛ�p`�V)sf�x�������U����ˌin}��}�4�����u���AP1Aj�f�+[c����5�O�T�UX�̃�_��GZd�}�!��5r�C$-�9���W��<�(�}ԍ����ѩ�$M\*�ӄ.�e��*���2%)l��n����.#���]7Ey��F�OW��s	ܽ�iJ�î5���v.L1pw���f:3�������v`C�a�B�٥���{m\��N�P�B��q`�-�r�ص�8eL��앛��������(�e+�*Ս��A��7�$��I�P�����}�Z{x��IV����k�T^�i���T\kS�	��rgjět��tf6iA�2'mf��D�+"�l�+�f3�.^{���L�鬉���-��y�\�r��uMWc���(��]+���l�^f��u�\�ͣ��AK��ۘ =��p��Y]����=*&�v���v,�¬�Zk�]S=k�b��l�Ijү:�D}}�Rײ3	ׯV�������k�Ư��dq�f�������j�f�s躃x�(��#�\38\�o���W�Zq���(�72Q���.ύ��mo���삷�9�6� ����?/k'�������P��R��zCݞ7���x��F�Sg%�i��:ݾ{��nI7�9=t��f(�XtK5<�9^��V������Uй�m3�"�6ϓ�ֶ(�Y��D����\r{3��������R5l���\��H)��g��_Y�&�f��A���K���p�UJ�˧>�T�х�����<�M,��������-$=����Ӝ�i����5�	T}=�ݲ�y��B�9K�1�Ckmpwgo�QdvzHi���S�G"`��-��TK뿤���;�,�dsM�ѽ��祪�U��ޒ��/pEB�#������WB�3�h�c�B�*��a��ǅ�`�YLQ��3��P��s��bnQJ�ALs�[�,���s���WG����&����7털q���EZ{.�Y�t�t��$�Y��k2N��TgRp�$U�w�K��U�J�q-!�q��Պ����n�ﾯ��s�}^O}ϲ?�l�0Zg����!�n}>cv��D�t`�-���lj��'�;���z,�OZ�3{\�N��3�*ؤ�6K3v����'~Ё�5�6=+���2��WJ�:�m9U	�o��x eb���K��mE��\���f�،�W��V�:�%��oJ����Śzr��F���_�m�CF~�%��r�/\g��mmƯLL9�ャ�2�(�N3y3��޲�*���F55	����Om�v�m�����`5�t9eVi�Zu�|�s�7�g8�3�ݐڜ���A���q���O{vU��)U%��t~��]�c>�ן_�V$�>����{���oY���l�����Tؚq7rn"��γq�U�k
�V�-�}�5�o�۱
u�]f�洪�j�cҮ>T%�P�X�7���A�?�_zP��Ν�2��ݺ���3�f��Kn�7n��#��aުh�t�q�*5�p����	?I=mc��95Y�(N��[�*�am�WS���n���H{%�V���d�8�rw�	�>T4�9��/L�y��oxR�ww�L�x_��ff�g�.W�_U��S�����[&��>;��9�`�ۥ��{���g_�S�U₏�b�;Ain���(]��g�<O"N�x�+�0v�����������YX���m�,{�N;UB��q4���1�T'idK�K&��U�P�zp)әu���䚜q�fD��7�ޚ��_KΕ���:4��֥�Ӹ���%z��>
�o��[g>'�Gt�fJ���Rr�X�������4�DC�0��[�]���YP��m���^�(f���v�mL���L���­�p��v� �w��z*5k�V��u�=c>n��$��w�e(gk���5�w>������x��4���da\2��N��!��O>JښZ�pDs�y/7�Uh]�������EWT��=ֲ��^�cW��}z���o �Qz�j�V�����d������}\4f6��'��ԑX�&�^��BU���������E�3FR�[S|��<M�Xnp,R��/�{T�;+l���{-r����kg�zz�%a�={�ܮ".t�,zz�u���[N�6�f��/�-Mpɲ<��]�ۓ6_1*h�_}_F�{��S�ѧ��z9ٮ�ū�������=�^�x��,����q��%�p����|�,�+��hWQu�Wi�v����㵻��]�����i�s���k�=�^A�r�dok'��s��i?w�P�qP,ᨦ�ikN�n��S��t�w~O��4�K�&6��3�J��_�7�m�Cu��{��<�G8��өn&�ϩ��s�� �F��+�q��)D1�e������u���;��c�+�Os���ƘŪ6M�5
��O��:�����lo,4�"�֏��8Rè����KK=��j>N��#�w�s�3��=�LP/U]�j��uQ%��E�j5	jW��'�fq{p��/�k��x�Z���={E�H�0DL_��-�}(��t�5����B�Eo:���;	q5�oQ{��e*�0�_���u�J{�>7PTeZ�V��w�n��;J�jD1��ɴ��k���3*�@�Ӊܑ۫�C V�&�
To,�s2�w}�\��V�nf�&��O�9];n�p;3g*}����ݹ�,�U���$fٔZ����&�s�g��H�6�-=*��u�=�Ϯ��a�f봆dt���wu�r��%�\w�{!�ox���m;fnՔ��V��9��D�v�7�!-��]������u��h�a�VdQ�폨�D�o��X��.�*�VT����;8j�̕87x��&\"����s���D����lvۏ��E,Y�݀�N�8��}��@��xB����S��j�@1>�O��lm�FeX�ܹcGn`�|"�,U�u�ے�E*����;��ɵg.�u�1&�ԟ5�����K*�w-�����q�wh�:��]�pf���\�r��pD�o���������@dryk�����,�|�s+�]`�qbע]KJ�ʱ�f�����#`�z�}wo�M��Q�|f�2�A��Kͼ�ښE� �Ұ��lY=� �*�0��8�W(�wZ�7�I���hU��i�sgRQ�����;V^L�%n#�5�-�����Õ�(��o|��d���O��[�F�<�X����`�Ǎ*u�rص�����yr��Wj�p= �=����m����O%d��k��O��`���u�&�W|�[���|Z���tw�VX��'S��.̷{�Z9�;&��R��]v9��\QO��{��ɬ�d���:��A�$��kJ�o�jY��|�V�+�
ͳ���kݯ���fe*��Y+��k���B����.-��G�Ltͻ��;��_=�<��oV�s�v��F�����)���Wvo�4�t���.�w ���@L��0�6ۨ	�E�	�
E�L���nۂ���H#���l�I�ۿ��]�﨑�����!v�wR��֭v�c���>:Q��Ǫ޻��\��[X�.+��炱�DR���3[��N�2��38T��	|ﺳEN��b��v����Ѓ���Oz[�t�҄ի$��S`H8q�W)�+��S��Qs6��0��.uՂ�o�<�:]���𩺚Ĺ�Ѵqk1�oy���V�y]���L)u��>�S,u����7�d���op8H�NM�	b�L�鹹�ekG��4�<�u��D�V1��QVQ�5ݦ]��V)ѾS���u�Y���n�@a�!�Ve�3���;�Pur��m��i��Uvf3�/�2g kl��x��':�h��71o7$'Z�M	w��V��V:4���
�-��iuN�ǺkgGF>3�U�q=}y��V��b֡��Ғ^����>W�pi�;��g��i�3:�rƍ-��mJ0x�u>�	�RN�/w�b+���t�457���%�x0kW����F^0@����B]6s+7P�{�>��T4A� U��sD��1(��*�\��$e�#�����#ǎ�9�W-EE"p�AX�EJJ��T�@�y���R���I�Z��jG/Q�$�C9(XY�J��%��Q�\���P���Z-:�V��KP�"�j��uJ�jS-VbUEF����IZy�S��Ǜ;���g�VUE��D���B5i��0$�:eV*�u	H��#4�UR�e�b���D�*�Q\�֕IȔ���%0�w0��j��YTa!����"�BB��Z�%�L-������(�I�RK+��Y�a�jr�[��Q�9�A�R��ӨiFi]U@�K�0��KA%�$��Q$�˙D�e�B-"#	:�T��f\�r騪U0�IFftP����e�l4��iY��\V��F�
UIhp�Ѯ;�⢪L*8fGYPz�0�ٹUan�N���kE5Fi�4&T�3����fY!s��k6�� o���#�j@����Y���A�G�N����Q�����Ic؛L\:Po��,`̮�-u���r�.ڢη/I]�.]�0�૝�����[͉Ȃ�7,��ԍ)�}���ʛt�G�5�'����eR<2>��:��U�jCI9�s֊�xé�S��}�9^[��}qˤ\F��y��V��['aTz���	�/�����c��t��t��I?t�r�>��lV{W���
~{|���Q��\r��G�^)mO[[��Z����a�><)c��F^�s����K��c�s��es�cir~�+l�4���{.�C�k��v|�JD���i{��Q��h���}�y�!%�۴u���Ҵ���;H˼n�i���r�Kz���m�_n�0���%����wѥ�^>��d]1x���yh���9rȞOr#ƻނ
ʵ�כ��2�W��������W��Sڏ�^`�����RVYQ}nm3�ږ^>�DU��fY�a}�ʹޯVߥo,�HwY!�=C��7:qЗP�9��\F7lm�2�����̰��)��P�E���e,U�Ug�"2���ΚF��|������v;.(��\���'�%4����W�4�Λ�=2�UM�imB)����)�5�'�f�or#Q9W9��a�_-sen�{�6䕟>�����K�"��_����}��5�b,�Ba��[H���:�\������່���@�	�B��/"���ag1�֑S�l_�grNgK\�E�L����7�z)e:3�[�!�3&�ך;t�[lf�Z��j�������.{"v.!�nӽ�S`g�ذ�cFD���ꭌK��h�=����Tb�W�+�������ۨ:U�Q75�槏������Z�P\���lZw��J�R�c>��t;��%=A�/֎�-GO�r�6�N�����?���{j�ť�R!f`Q��~������o���g`�5���i�ێq=�[�\pN�|�f�b�}x�G�f�36�o�:໵t�ϸB*xYbWA@��S<Ǡ���Xo|�GL��)G*��r�C�t���2�0=n.�jZ.�4����)�`�Y�5|�����;p�����DU�n垤7c��V�u��Ӣ�g�qcz����tcԳ1��1�r`j;�q*��fܿ꯾�M��|��x���}�~�)q��
��ղv~�ɟ��f�g�-�,�J��'>�u��K��H�ylQ^:���Tj�F�dF����o����p��M��Q�cI�S��}�\f�6������W�]��
�4Vv�[��1�����HGs��o;�Ӿj7���Z{~��Kc�)&ڪΡ�ݤN��ToM��7�8�ܲ;02���.5&�Ŷl,:���\�h��8�k��^iܳ�ׯ����ͬ����G�zB�� ]z�\t��Сή��W��$8�G���I{��,}V[I�;�\m|��/�6k��3ݢ�	F⩭2RR���ز�=�˵��B�j�2reK߻y�*r�uY㙨L�'��<�iU�c{��!k�(��Jt�5p��Ϙޓ3Svfyc���<�L'�TB�U�z����]��)���-�I�T`m>��fv�M���nm��pK@�,��`��/���X�z��Y1{PI��ڗȧ�ō���
��oKf���=�v�7V���K,����a��Zc��w%=�I�R!w��TJ�}�U�aa|�:O�F�0��Y B�tfQ����؂�\��Ֆ�������e�IN���:�_�m��U��؜���;�ѼK��Dl[����o5��C�;��;*��u*�Q=e�CD�8���Lݑ7�#�̣w�y��6���|�gں�I����8�[�9`ǘ��A�zg���<��&�g��fz�kj��O�
�O�r�4�$����&��S3[�m�M���͏�S�g�l��v��c5ڣ]������r�w(�l=�(���wn��nON�iy�m�@�{Y=��_�5�j���7:t�X���o.����{mo_О��|
ܔ��t�R�|�5W7H�&v�-}�����5ѹԷ>\�g�I����}x捋DZ]��1�KZ�W����VoZY0��EYmg�E�×,�O_J�)�����:^���a�\�Ĵi�铥�g�ݱ�;E&��@YRk��_c�oTxC|x�I�v��59՘ҙ�c1iZ��2�c�Hݸyn��7��c_A�B��5���e�����f�P�Y!�8fQ��W�����EI\ܽ�{hRKUf���o^����v*�9n(�&gc[���%��$᝸��:�)���5s��s�([t�����a-��T�f�{���Մ�{��Е7 f�ĮZH����As���Zt�dL%Q0�|�Wҙ�G/�SX�k"G9�r�;ݦR�ݬ�H�8��S�ʸ��P���AudE.{�$%����+�/��(�2�M��cd�=��ς=��+{�w��V�I5������'3k7�;+*
�W$���P�����w�w$���X�������o���|;�z��}e\����q	�e �o��G�!�|��=��^������'��y�vV��5۾ڞ��TSi��U�x�:�}ϙ*7�5���K��ro�;:�h�v�V-��ch���o��Bĩ(ϟ(��i�FJ�1��z6พ��3�T8��b�t���஡+��Γ��,@�`W�c`n392�O,��UyN�x՗�֎�l��,�veP-03�p��E�i�������7]��O�-���` �{�S0^����Zg�Ձl�yh��FV�s7���kY��Ξ��ŚNue�}�q��{��=�k��'J�����v�n�|�\��r���P��}�}�*����w��8ۛi�u/tU�zztj����(�g���{�	'���c)W�L��we�f�yW<≬V���T�Q���k��̢r��yI��l� �&��E��(�p,�S��W5q���E�\�y=��#r\+=osa\��5I��Y�>n0���s�#�R6��¾�Wޛ�V{���^�я�e�K��Ӡ{[ݕm	�P*O+6���W��==�"gn�P�����To$q4�Oq��t�<��[�L%���u ����M=��G���A�Z�'��8ɛ�̧�S���ਅ�������݌�S&�7gl��obCΑ�i{�J;�Bv�ml@j�*IOa[� -]n{�G^�Mb�����<WEG���f����Y�9���o!��j��ۀ�aI���dΰ/*�*s#�5�d���ƶ�����~���5�=�*}n��ٖ(\�R�� j�j=����0��}ճiuYN�-���S�A�u�.�k�����u7WGU0jm�����.r���P��g]�ܣ�'��wʛ��S�w���r���Oh�mQ	��udzf�>ہk�3dս��|J�%d�'5Q�|.vT@����f��'��І	-��독�f��b�l��Ǘ�U�w�t��>9�!(Ƶ�	�4e�~�%��t~���uڧ<�i�׸��Ũ�\��R5Ɠm�U���^��Ol[����)`��1=Fr~G^%��N��������ۏ�ƻ����ZXzMS���W ��/��e�ر�<Z�x&��՟S���wڣU�6�`����m���ɺ�F᲻���(5��r�ܗ�;'��.����1�V9^����lLJ:۠'kA���o>-��y=������W:�߆�{Y�+_�h��Dm����P���f�|
}�2�;iе�vJ��4n��JW�Dʑ"긬�I�]g__[��$˂�}(�D&�����[�j�w��:�һ�;�Բm(	�ǫ��t1��1�5���:�L�a)��.�SA�3[6pl�6bTn*��-��:k�,���Vԙ�����$�)G��v�Y�ۮ�#R�k1�\�Z��%�ZX�+�܍_�"6|1(Ͻ	$��L��� #��$[[c�_sc����F4�Q+Qm%�h"v>d�æ�$�z�*���]*}F����>��7��RY̔^f�Q	�T����ϡ��]�F��iZ�v����������������;��=p��̀��֪��yiW4���S�,Í�R�r�P!:�3K�7�Ow[񥼕��d�w�p��E(ޞz]�CS�`�'�_,�Fr=q����Y� ũ��4�Ji�h�䷺Vj7:T��j���h��;4�Ks�u1��G�w&K�U�҅j�{��*��R�Q=�����r�Q�zl�m�,���H������3���i��*�Em�r�>q��c3B�0k��н�G=JU\�P�Z��Gϊ}���Qf�(I�3�/��sТ���ϰ��Tt'g���iX;z͝W�Zq����q�\�w]R���������hy/Ev����R�oQ��iL۳-���(;iثDn�x�y��N�"�K�,,�ꄳ��e��1X� �믑Ĩ�Շz��L�5��҂��J��;�sT֊܇����z!:�$W�_W���ܽ�m��E�6�s���>>�����5@�byQ��׆����W��g+r�V�W����["��O�ŭ�OWdG>�n�X3'��%s�V�H��F5�1f���#���?o�M��Kq4�m�l���y�}��<�B.�Y�+w��\*Êp"(��R1�]�%χ'������uL��v4�K-��J�>}Sw��g�;���Z܍Ec�e4�K=�R����]e4�q�c��83	TD�%t�R3��:�B�"��9�;��	�[A�t�恷�|�`wj���SɄ�鄩���d����z��:����Z�s�F���1�'!9�opE}��0�؂���b���f��ԧ{�]͆��VRL������1���2!]:���5R���&.��
�9�=�O�������+8��I��aC9
��b͘�{�]̉#@�Y3�{.(�vǗhhA�,�ܫ�!�T%x�vQH��U��@1�6d+�\�[��n7�ԩ���-���JT��Y� )A��XlAy1=W+��舟�/1u��M\#��;*�9N��}���Z=sJ�T-z����)]ewb���DD��u�c.����p,��n��\5k��YĬ;C�Zq$n�[Fm'�������Ur�땗��4U�.��}qˤ^���=*��-�GzD����c��^=�{ܷǂ~~��G����|��U.��yt�M��ҷ����J7y���n��7Z����.���T�ZW�6{]QJ1��<`�f�>WX޴����ƛ�9G_�[��x�q=�zE��G_�l�d�aH.�$@EhC�:��o;]a�5x5�F�Ԉ͌��9J<��\i}F�D�K�F����o>*�kX̒߰ڼ�02�+�[�ev٘Q�448��{��+Ӊ�bQʺ��ҍ��)X� (��0���{~|�m����YsL���$�s��i}��zTt��n(�Pv�����)\FR$�RK�z�8���E�ͫN��K�0�u�����Ȩ��7B	�؊��l{c�-��&��O�T��]w��T��<Vy۴T"��o�b7}kANV�;�w���jУ61M�ɰ�T���+�﯁1Fr^��~�/hY��a\%O\���n�O뉣OQr�\s��
yn�Vv���{ÔaoZ�������xt�5�۸Fei��8ز�:�p����x��(�ڗ&n�<����3�Pu�X��L\�I�*�o� ~���3qW[�s��r��V�Tۍ!tX���W+z��ܫn���;܍A�l�״>QNnw@���c�a�b�e�$��ac�G�Q�;��ֽUn�Uq�Az�-.���TlH �+�P���I5�o3:1]5:���r�W�)R�Zc9çCtKf�%N������m��x���y7{������[��y�nJ5�B�kyQ�v1t��c(;���'7Z1�ֆ�D����%2��\33g��K�һ��� ����7�3Ju�n-�D����`���LWt�8����%)ǻ3p긂N�����m5�(������wo�%���A#*5�������g&��4�.����K�'U���4v�iJ�:h@��/�}��RZm<\�^\l���pҴ(�X���+S�d�3"aS&q޻ј��A,���#�Qn8����j]��̻�� ����D�`˦��gv�֌�N�VtTFP��Q�d]ơ�.�|<�+q�Z�X����m̗�DRB�qjܡ���W��u���[��ie>�,Gd�L^��*�v�G{�F����[�\)ڬ��y�l���X�A`�e�I]���t��z��i[�u��	29��F�Y�X���a�E�S�"�^�611Z���E��+��x<�+VY�/q_m7��c^mƼ�ͦ�'8�.�R�P��ѵ�d�wv �&	Uu3_�J�:[���c��{�.�Aj�8˜�A|fS�t�i�� f!��+�G%^T]��q�jng�읮�ff7�+8�Z�˓��i@��&m�b�����b?hq,6KOn��N���V��/Ei
�.����u)EWc�#)�2��N����QBm��nu�u#i�S4k���3�sӷ�38s�c��.ʾG#o�u�A��e���QhD���ʴ�nLi�w�vP}����T:��t����Ս-�(WX�e�bj�W�j��7�S��r�/��u";5�Af�+/jt�h$FX5���f��Z��)�>�w�%�6�^��KDJS-BD������xo�M��ux��6{{�i�rr���2�x/�2Y]<��)d�j�� �ǰ�y��im^��nl��<{ǆ���޿�b%�`��8��C�Nڨpd�[6c���t��J���\�B(jN��ž�Z�ýft������J횵
�l��Ü�.�����ß$&����v�ӔaOb��yt�&��L�+N���C���\g{wZ���oB�[�n���ԮM�uàV�]O �����rO%��!<�N����;���j����y��u}�������"�\��I�ͪҶEhj ��(×B5�q$6U�"�r��F�*�D�R��ʊ(*g
-@�U���5Z�Tf\ͤ]
�4I��#�r�#g$��L�%�Q8�r�0��#�:e*��t�2�$�UQR�H�.\�$&hX@��QfFZ�IirdR�HJ(�G�8Lʨ�R5�I��N����dZR�L�(8w+�΄��V�fUu�p*�DVZf�s�s�r���R����YBH�TQγR�3�l$�զ��U(�.��$Ȭ0�#��Z�f�0�)�-3�	�
8Xg$RJ���MUq�NM:`�CB�H�R2�jQQfG9�CR�:U�"*�Ȕ)"���
2.k��T&I%1(�Ў�%Ix�ÚQQ��:fQUv�WD �+Q$��L�29RV���Va�M�D ��>1�58�j�{�s2�m����b��ʱ����"�ظ<|�Y΃���n�e��&�]�ݥ����d��c�%d�+���yyM~h��K���M+���gϧjZY/](+�
����{�s��vw�ʹ���f�_B�j�W3�񕏧����1a��jfL��w�����y�-�#v����-ȔwL�a��|]�{8��n{]7�a��4�-EF�O7�}�niv����al�<٦�1U����q"��j}[�Ob�0f�>���6ME�������bZj���X�Q�<�����Pց��&�anz��.Ҽ>)x��Ӗ�oOT��~T��-���ʥ�Q;О��CF_��z�=�B��c��R����C9~̈�}Z����|��\���=����i���P��J��n�//ͭ�q��+�^�P����b9i�Vy��]����:A'$��qO++U�>��T�zg�S޽�����#���{^���x,`�[J�fm̝#���ټ��tʡ��)�'�G��.[����-V���+#(]�U8,�;�=���/nW[��2������d.eb<�0{�M gB{Y�g%ݯ�+��_*�3f��9�v��I�ק��}�F��̶�+�Z���an�쁙=qE��m^w�
�����#j��n3/!s[�'�K�$�l^�������]��fz�E�[
w;��hʪשbR5�Wѥ��4�߭�aa��e�sJ�:�k;��Yk�^S�"�K�)v���6^} ���]��u�)�D��j�a9���G�/��W)JgT��h���p[K!�=ٮ6�����>UO1��z�����N�N�L˞��_Ov�-������6d�����4�md��Y��_4�BU������Gw"S����x����|h.%��K�F�m���q�������?g4�_y#�f�c&�ºr�([�F�fq�q	��'{īc�R�-u㗜������k�jS��ס�r��=��v�I��&���VøC�l��M�7u�ٺ����׻��eô�*�욯V�Tﱨ�Bp�қ���WQۧ��bU&���v���B�2P�B�wS5757[ZN�6U+t��x�H���E�jӕ�$�b���[��u}٨a��5p���7$���$O�V[���{����di��
�w]������jZ�a;�9Tk7�ܭ��L��cy^n�����>�Qz���o"�Qz�X�M�ʙ]�Y��R�:B:6ˉ찊߂�ϴ�[k���ճ:�,��W3P���=��C39K�Pn�.��,��C�o�qӊL.��)��.�..�=��)$އ9�U�Nz��Ǜ_w�ߧ�K�=��[g�����rw/Wf�ɊoQ9�rT��@%�inj�o�-o\*z���rR�s�7d󸕹B(��άqi�gv��;������t��ks��]�m����|�v�b��WwT����p�d�Ȭ�������mp9r�
}�܏d&�k]��l���a�Tr��6{��wq=o�P)#7���F�>p�L_B���DE6�"��:sKj6���N��&���)�JFq��4Ú\��k���"e��N�+�.ɩ,_ 2�v^�MoQ�_Iۂ���3���6;o�7�e���k�9���oM*�YQ{rN�H���m]��V���=�+s�Q�����9���井��|���{�]�i���nt���$>��gsk��e������L.o�i媸N�,���&�j7}��%V��<fx���u9�?eW�����Ϙޒ��/p,
�`�=b9QqDTVM�e�kvsy-����n}<wr{i4r6�Lg�_BǺ�:2�;ٜ�z�Yo�wt;�X��.�N��y���A��5��r�kE��ɀ�)���n�((K��7�v����8�wڵբ�ʹw�u(�̵C�N:LԬ@Z/Vp��j���'nN�^n.��ܺG^�9�}1�Ú�b�.r�,U=v�4_ѧU���ї�NXggU��skLVPq[d�ׇoY:�v���O���g`�5�8_���糾��Պ�-�u��CC�x�j|^IO�u�c]�}OS��?R���{�~r-\��r�ܣ�F�2ۖ���o�o<�(�����b/����Ok�����e���ɺ0eQ��A��T�YP#{6[���NE=�!�����O!
J�y~bo,C��/)[�^wm��kl��^��q���6�t�����~�/��s��l�l��m���S�^E�/�kU�]�h�O�c�P�� �����LQ�{F�[�h��Ev�DKԻ����Ƒ~��J����'Xm\FW��rЋ}�k)�ԩ���D�r�x��w�	����9��[lZ (ϫ��-�˒nbz���W�8��r�	$g�KԚ;ٸ
Ϥ�\�A���(RNo
\��T��<���\^jT��8gm�G"�(��`��v8�Pյ�u+L����m�%/��k5U���fIY��ה�D�t�a-������Ȓ�Ύf�]�l��b����>�e�k4���VZ�4��9ˣ�6&M9�R.�ES�ǭ����1��j�	�Y��.{�w�'m�s�F�1�Np�m��w|Q��9�9��	����σ=0�b܈��W�����-\���$m&8od%ƚp���V����p���6M�����A�X�e��+jIQ�������n	Sw	�g!UkS�vanz�[7��'-)7a�ѹ�����!��̸�����$3������E��+�'�#tx}z��,9�PM��8����C����=}�k%����-s19�3zZ�i�V�lbZ�cɟ\�R�6!1��H�x*�\��F��E.��p@�������>���Xڽ�R��dT<��]���U�q=z�cؗ���܀�у�����_k����G��X��:�E�&���Q�.F��'��`�kMz��O�ϖM�f��=*�[U1>�=�P\;"���׈r�z��s����s$��bga�.�l��l�3[�0j�x���5(譖�k�z(=����o�o����S<ں�O����o�:��z�hng��Zw�)�Y4yWI���)3�|E���a�NU*|�fCͪ�V}��)��X��VN,{Hz�s�َ�1�ލ�O<F�����\qmᝃ�-J�f�mକ �]���>�oN�9�b�k֫����)xi��|n��E^K��~�����!��dv���L�
�L���:���t�'�~��\�1{#������+��6���b�oҫ�t�x˴F��z��%� �r��\����Gc)���G����싺�\U&��q����*w�y۟�w3���۲#s<��C�cWzWp�D����]�az։���u�V�8�֐q�ݸ�eG���:��
�1QE$(��i�&E�]�I�!u@�䶚�wu-�3�u��u�9٩�SB�+� V2+�Z}�
�����d�h�r�S�dF�{�着NլV���g>�t�}�:�-���z��um�Bu@�o�:;���&����d�y���O�?r�n{.q��Yb$O������*��k�8�v�C�wN�]v�P�[�zXb��ў��g�6����e绲��ݻ���2�9���������S_\k��]���hLpBNj;�3v�:�1���V?vL�ݿXC`T4V[�{�]O�}�j����R��~�82�U9��U�=l�t{;K���{� �0��n���F(ރG۞깆I��{�RS�}����=Yq����Fפи�]"��>�� ��T���R:��^O�������G�t�}�/�)W���~ǵߊ��x�����>�"��3)_���[̯	N��,�/��eg#ڻ�O�S��2jzny@&Q�GR���T���[�/z�������c�buǝ铽�y(ᾙ��a�<�B��iʜ�����н�D=9����;���זQ�a-��׽�0^���e*����N���1����1��dv�(<N�l�T��Z��ɕS0#}�����]ڷ��Â�mRU�W�>������g�f�߂"�����>9Hd>��Qq@��]�{�<���%sQ������D�H;�:��[2�t��DJ���=��eA��p�[��
�B�X�e'��Y4Js�=չ���zӎ���O��Ζ^
ɨ^�z-U���gN� �k�3�!9y��EeM�[��;�h��r�t����� ��i-�C��}����x�j����2���(ɦ�K>w�e?�b��W��·l�����ڣ�b3�E�1�Y�ߦj�3�	���^��t��߼f��B:$+��{���9��:�(�\�}Gp˝����E�|�]�UÉ�n�+���2C��)s:3��⚸���e�sݣI�G�3��_�ۦ�"S� ̷Y깿�v�dm4=��dGO���1"�o>���|��{O�E�'����3]>�ws<�~���-����jG�I7U7����W��W߉��jW����z��'�y���`:*%�^Fg�ܵ� �[&n�sʽC?}KXZ�~�����t�~�+kֳ���~��]tJ~ۊ����ʳ�p���Y�%��a����8!�����m_X�==�iβ�hv��2=J�ާI)���x����І�H�>BԌ���g՗��}�o���|=e���N�$��mFE�{3�خ���f¬'��{_�e-uw>��֋g�@�ʥ'�VJ���y������(�W6�+�䦗��f뛵;�>�;4��wCebζN�U���������^gr�-�a�k�,oV/��0�>���}m�l�$N/y�yg]?����s���L|
��A-W��_vK�B�9�n��Q�D��1�²NPfr�3z39%���[�曻J�9-��G��c���E4J��WS���_K��a%(�/[�5=��`�Iz˯����5雈՞���+X /��P����ȇ��ᐇ����R���O(�s}f��A�������Mh��Oz�4ә<�zB���Fſg��qW���Dx+U�D�Q>�J�!.���=��ݹۍ���6��0�s%�+�ی6���[@�;�%����<�x\d��9���h[�J��HG��6��軇�q�-�mW1�U�OA���^�ޯ)x��nf��󲇻��;R�"��rg�Ԥ�nm�E��*��՟d<��}U�Y,�I��.|���W,���{��GZ^9�ߘЮ�J�|�~���V����Uw��y'����c!�,�lJ��6<hx"7�ddW���к�2� ��[�������rg��q�t�ռ+�WS��,S����q��cُ!�O�ݏK����n�\_^�����F=�< d�g�f���X%��:�*ެSy��)�~6��'�����4sݏ�ӎn�O
�ɀ�T9��:Uڵ�Z�t��|ʱ� n�'-n�]�f��Û����D�B9��8r�e5�z�Rg\�onF�r���U�J��[�ϖ^h*�T|����8R�z����^�w�V�k�#Bo(mi|�{T�{|�y˔o5v��J5z*'�˅ǲ&C�**��T[7��Mz&����Hz}^w�7\g����U�W�ήi$$���C�����(��?�h7I{�e$����(�f��G�N�p��%v���V���*�8�Q�>3�z�L��W�2�!��e敖*�'�\�=�%_���=�`8殖~�Ə>�c�x�~A;��?/_`^~��B.�϶'�|C�J@�ezTl�@f�4�Y}{�W��+-��r�5q��U�^�b{�^��Gył1��#��]h�?	a���1���t/mL�~�M�u�K�9>�k�,����s���%�����}�R;�\�?m��\s�[���|��`�!��\2��;+�=����
��s����s'U�-�.�q7ۉ]M�Yۋ���~�������h��o��C��[p�muC��Y��Φy�5�>�i��jM�z}v�n��)��﷍��E���OI��X��4�TgA��
}z�!�mWz�.����u[�ǣ�w.j&�����g�߻����dq�y��9�XAg��ͼ�Y&AȻs*"'x�	Ջy_�6S�O�;�L����e0B8cU5p�u:�w7�.K�&1�ǰpVNɣ�L\M�T,��ܛ��C��e}�8���a1�t�E��e�ᾆ�K��E��y[�J�n��4A@/�̉�;�:.��x8]���L�����)n�-"�WM�ܮ��y[��{��g,[O�$�&fܼ��
�W	V��r��8F}�@�q���AB�2�J��\��N2sW,��ȣ���9�iY��3U+����0��׃p��i��t��lq�_0�ٺ����;u��X)f�,�T4CW4T����2�f�k:�;�)�;#I����2���n�j
.�c'�r.�{�mh�3�|�U�헆8�5(>O��C��x{F�s2h皢��VZ��@^
F���|�3�=�qd�煮5�yR9�E:��2,!�m��Ģ�=�j3d-\wB�ۥW���`�յ<0u�+��ˑͻ���:�)�0:�_d�R�iރgw7ϩu�r�/%��s�y]���6������eC���%�*j��� m_��
�9���q�Z�vi|x�m�R����"�5��|f�pbp�ٝvE��]�ץh
qXc�y�r�"锩<��Np����&8�E7+xƔ�vsq�"��+8�Zu^t������ �$�(]�G8��	c72�y!��:ݾ�u݂�ݦ���"s��aul�'�;$;�ʗ�M�Y+>�,QIgi>��&����P���x�S�%���R8�]�c�;�rƮ�������S�[�&����5�EJB��ǃ��z�Vm�qhAs2�|���y�w��6�s��2��� �+�r� ���$*f�M�����&	PR��4���]�1��XchV+��|sCB��%���u�F :�<��O�h�I:e��d��//��v��;aC5�v)^�ζ�c��	u���8��iX��.�:�e�n�MT�>��#�+w��Ս��lA�;��������<2|����'��Y���k>��*ӏyX���Ò�_r�
}-Q�1]�s��72����g7��j��췍���/�dG#x�� m^C�)�*fю�_b�=³^9ztwa��wg"��]ώ��F$鷡n��>�y�
ύ�1�I����L���%M<��K]�u;\�ҽ��n��8��ae�v�e:;\Q��_E�P��u���وs/[u�U(�{���N���ls#��*�9��+C��H����)�i�pB��N�1!�C/���~���{0bp�7���[3����+gE��s��;DP��f*�OS|y�z�����т��Zh�k�K�U����,�&�ݵ��ڧA-�}�2�:�oM+U�K��}���û�`�:�������f���*빣��g�K��K4a�����r�y��f�\��7;kk�v�Q}>�b`Pf8-,���h���O�x�ȹ���9J!(����eW�J,�T�9���Q��J�ZJBr�9ª�EC�U���'��R�*��I)EGr�AdI��5(�E@ŅJ�E\ -B��Iw9�1�*��a�:(���IJ��Փ9V��Vy2��*PN�T�GN�E�MI�"�Er33*"�F��3�L�3�D��*g�24�NQ�(�KQT^T%�h�Q��E%9�G'E%rI*�G�")�����G-B9��EF�9\�""*��U��8W#JA!+�QW9QȪ�r�E2��r��qR(�""�"HЉD*��"FQ�s��J��GE"�DQ*V*ҩ�\��Xr��9x��EDPd��"�\���G*�Q��� ͤRȨ���+uWWW��u����]�\�uA��j+7\ފ��kA�N�*�y�-�q[Yz�_47ݧ�³z�sf��L�\t��m�:�<c3�X�*��$�;��]\���~�����Hk�q��c���mpW������c6���? �V��!���*����ߧЇ��^2����2��#�����_�X��v�@���iu�5(�bH�;T%�������S���j����ns�h�,Ĝ;��w�=ܼ�����,�;󬇳� b[˵b%z�����Oq!s����������'�nyh����G�<pI��ۏ._��p�H�: L�:1U̳^��4;��ծ���p�Y�����,�=��"� �Z�:ѐ���2��u2�	!����}q��٤C��;���[�{����{����Hhw ��7#�Y��c�7�}s+�&m�߭Pت��1��oX�X�ſM�쩍��>�˶�y��8ؓyK�O{����)�'sq���eC�;�*P�\0����%�ሽ>��QX�hi���}Yq�����@��Ȭ�n}p���.��Τuz����w���K�ѽ�J��ԟCu"mz&��>#z��{>���7��dQ�W��e+��	�����նgS��a��WP��f��v��v�R^�T-�)��v���֧snk�_v�u�	��i���c�n��oG�����ol@}%���+��\�,A���K{��*�ui���o*�l�)�4��k�7�^j�q��G7;�'E�7�Z;��b�_֖����9<8_���i^Z�z� �1T�쮸z7ơ��/ëD�;�ˠ�.�~��>�؃�`�W���֠ƟdI�ӕ>����� �Uzw���:6�!2~W�ŻM{؛XW���T��y�q'���(�V�K��}��w�(���&+kd�'����}4�����/��^���mWz�#�Ju�Gד�-{=#Ɵ���1oڲ�]!پ�s��~�+^n���xR�`�o�_E����K<l�(�,�[=M��~w�g��w�s�ޡh�C=���ؔr�A�q��,��.�d*��͂���0��4�r�_�����cj��h��o���١5F{�R�>�C�[�\�*eL�����t��^\u�C=�x_�Ռ�QW��*>1�^��O+����zQ���=/������q2��2�W�N��R	:�)��[~���k�8��;<�C���\�H'� ���]7��gNǪ�d���� )Q�h������=M^���/'�|2�؉_���,��g=�z��o��y�ʗ�N�ˏf
��N꾕�"�����H\���
w�ce�i����_?�\��x��]F�������Y��!�eT&�AN��I�Oj�fʽ�]ԹX��4ˮ�E'�e�� ��<�웻t���yRhF����7�&hmo.`.�k�d<i�S+J�o����z��n�:=K�l!O�CO��}�z�UFG�?Ug���.���*�b�X����g6�5�#Ѫ��"(&;"���#o�E[W�3�u�%M9ҝ�9߯<	�bC������\Tsν�]#����:�ߋ�eR_��Q׶U��]*�f��|=x�zL�i��Ɗ�{˵�d�Y�R���o,�ƿz�A�u>��S��9��b\7c�r�z^?�E�	ͷ{uE�y���0+ܲ��e�L/]�'#�nA�ّ�c��dE7>�����Ndpw�J��&��N������gU9F�`�3_b�l{~��Z� ��⏕��@��6�]���CFoڹӽ���'=N��F��:=5�X��-4�Nr{�������2�dQ�x��m����x�=��OOOJS�R+���~C��v�o���@�bgZ�u�l	��m�S&�2cn�����Q���u��I^6X��4�Ƞ��p�.5e��ڮc>����&�����0_��YV�/�|�S��G������������a��R��nm�P�J�*������Ra��/*�xsS�^�7��t�Dk��F�w<˚_g�1y:�_F��i��׌�2j�㈋�\��o;º�pP�9"��r�`���u�c�ի�{��V��b���n�\��]�ۊ�v�;|����V��uʐ���+1�αlg`2C{je4F]��j\=@�����&��c�Hx���a������fWVXs>������uA绘�����I��s�1�,�l�[cb<hx"6<i��^�g�~���2�����H�+}��\��P�Q�z|Ʈ�*���7���yx<~Gp�۸}�6/.�1
��b=�Xw��O�<��_�-e���X;��xn�zU�X���v|��<��Ucb����^Q���݊����_O��QP�yh�������!Ͻ�H��&(��5�0*-�4��M!H�ǟ�L�c�#��߫��h&Y���f��G�O��Q^1Vlz9x#�����3�ϝz�|v_L��{�f��뉔���x��o
C������sU�����c>j�FBy7�_�`ϟ���ww������^�S�گJ C�[/���v����yvR�U��.�f�_Jͮ����ӟdj}�Ǫ3�W1�ݙ�:�@�:�/�fn��n�����>?��rW�����-`xg���?�O ��#�az��нr������:�۔�K����z�~S�҉���2�F�2��-7o(��`n3�P��R�oj�Q�0�n==r���s��AΠ���&���wY�.y#җ&��%���f����B�0��FԮ�b�Gw�!���:^L���\�����;��ހ��cs����:-�+��4xg��W\=Ϳ�xV���S=�ӎf�yf�3�^- �>��ó�����%�5�@z!�r�
�=9�ӑ��d�>���]�ѵ�=]`�Φy��S=Uꮩg���'��3�L�)����?{�e/m��?jru��V΃Y��>�w_-��
2�ol�ܹ't�ϩD��q�׳�lGy[��1��(d{��ӰU>۽�C�Ĥ&����P�����3���{��}�K�(��{<��6��4:3���q�u�� Ec���!z���y��_�%�ԭ�S|���C�Gq��J}�5�k��W�:}-	��C�dg��M+�'3��G�wﯳ�k���S)d]��⩰�����[�o}�ns��眚:#�������1���R>��w3������ެ��"[� ķT�F��Z4��c��ɚ�Z6����t"�c�>�'{à{�H{���{=�ܝt�ǳ�O�<�������o���Cə����5��ًۆ�y!��MA��J����{��h�I�̼�vT�=�v'!S��hx~TϿ\U�����˯�-o0MY;�4q>��� �7
� �kV��杤38�wG')�'�^X�ţ����Oi�ƀ�t�N.�
�y
���Z��o:��*f�V�Eh��ڲ���=�=�8�ul�WK�p��ˮ��53N1��:��Yq.Ԗ�K��'��P��EG�ߦ���,���Ǩz��Z�y��j^Ἧ}��7�|����Ee��F��)p���w��)��O&㱻�ʌ��s�[�|:[/��=��i�栯P�^��o�]G�}��}��49��]���ë�/\��s��<�~��!ן3�>��rŚ�y���ǵߊ��x���3�Ky��ef+�J���(�G�UC��@_�������M�#��%�9:z3|n�V�tx��n�����hD�܂�����������ki�D�}�9S��/�!{�� zsG}]Nwѓl���Kʭ����d�����V5^�9��>�V�OC�AC�dVG{���o�I!��E1���7�A�߶A�E�ʽ���ڮUΥ:�s�{=#!w��q��yU�Y�9��->ž�=u�&7�j��M�E������'Gjΐu�^c�_�����]/m��ۘgn^���q���W�-��c(b
�.��E�Bf��Rn��/(�m��N�b�=7;�Y�����Y2�ݥ����j�i�'m�:���p��(��l�
��b��
�.��Z�9r�[d�{엨*VgE��ft7΋�p�od.ZM�0��k��v���10�������dԵ.Է�wc��7�usk2S3��:��R�����iRK|�T�G��R�!��޹�Tʙ[�p�k�n�+��c���c'���0�+.oz[����EX�{!�O�!���$�bv}����h �e*�2�e��r5a=��z5��ݞ圕�l�uyv��B��Y�E?bC_� X������˜~���2��Sc݊|��`K��oS���]~!~��l:��|n���O����3i��K  ��py�ܩ�S%ɝ�'�ZF�v��q�3��9��,_[��ӱԸr��L7�r��_�z�ߪ�p��J���	���F52�nEymZ��ߨy�Yp�׀����ds�u
s�����>/ß���H������Buԍ�B
e�xfT��^�#*��g՗�m�Y��B����6Z����nt{ލ�)FyOO���s�7v��s>[���&�>�h
Nȹ^
#{����S�;bh+8��������H
�G\?�/�ż�����d^5cA� �tUzW��3 {���{�~�˶�z|f����#k��>��42#M9��՞��ǽW� :��7��ZDV������VP9K?$:��f0=*��g��7�=�F�!gR���T`Ic!Mi��[�n�t���hq�Ӥ]do\�2�6�9�%γ~��z�����@wC���܆W1ѥ\C;O4�%|����Wϧ$��s\K�m�uř��Ĝ���e9�;����\�Rµn��f�5%S���*�숮�N���z֎�u=�ͳnd��=�Ða���/;.�~=��B��e�z��8|#}�G�P������{���S<���4�`JP]d�6��b��š����IOmO��R�k�m���̛��q�-΁�`����ݪ����A>1��#�By�;�߼�>U�n�s��ѧ2Z����Y�Cw.v�O��0W�����/��F��/����.���&y����0]0w��o>�WVFzE�s5�9Xq�+����d��H�m{��h7�p��m��u��>��Ϡ-�a�����>���}ܹ��oG�eL�˺��:�#���v�9WV��m�~R�1��Bz"����;�B�s����s�pb�x~�G��ѱ�)�d�s(�+>4g�W0d�kw��þ5bpXw�{���%~؞̎��F&!dEEB��Z*ٿp��ݨ[��}s�^���_6�=��udy�[����3/=ݱSooՊF�T�9S,���f��z����SYU��#FK0��M��a^���y/��^^�l��3��J*���oR�����`޼�}jmwT�ub��:��@Msڙ��Mu}�F�Z��<N����N_9�t
V��}m��UގWP��vW-#Ԯܻ��`�Q��ػ��!p�cOӊw�*��S��{b_L��~외{�UzOg²\�h�:�5gǢL,���>]�^�6�_���V2�FBy7�A~��!��ϐ�ww��;TD/W�>��w����3Y����Է=��=Y^����sk���sªѧ���y_�è^q@����G���"�P&�dV_s:�k����0�{��ǿ���C�X�X??g���,����lzuz����Lt6'��͊�gfx�$q@\o��F���On�GAq4xe�dW\=ȍ��#z��s���Di�2��� #}����~�W���}�m�6,��;�57о��>�$mh�p�\m���������g���q���8<C��R���}=���5����K�jz{�(ʇ�a��U���E�>�S�ޘ�Qo	���?F�^�D���#�潞#c�O���=��g���=4PZ����FF{�L�5+/����H>�35��{6�:��࢒y�z������g���KVG!��Ov���a7���c�>���f�ȥS+���6
`�Amҗ���>�U�p]~���e�%�紋*��.��R�-اL|`��u�]6�3�c��=	�/���Z�>4����sك��u*��J�-<^�(�����E���۩'ۻR��M>#IaΧYVG������K��Z�7��!�;�ދr�w��3�:�iH�z�M�]v mt�����'���J7ր�ۃ��^w�qo@U2�".�|a��v�S�l��NI~��x�ΈZ�0/O����T����<:���"[���]�p�h��s��M��u�T��\ָ�i���T� ��ڐ�lOI�ۏ.e��ᯤO�p-�B�q�DY�<&�w7��>�<�� P�ؚ��i\Y��[���!���f^yX���۱9�,�0w��9�;�vrO���Gd.�<�p؅T�7�����߽U�z���O�s%\N�v�����ǳ+4���c���謵'7�'��R�Sqλ���չ:^NA�u�ʌ^~�
��������o�]g4�|bv��FDPh!utm��^�B��H��G�:�=,5��1����6����ޏF�\�Y���a���7�4�dPdvDW\/mv�gz�FQ�N���H��[>��79�홟wZ矮��r:�R^�ɩ[#$���M�P�v��?n�H��2���V[�*�t��ŏX5�s�3j�d�C~�a��B�;�r��_N|��D=9������?.*Nyu;J�4~ ��O7f�[2���B'e:��i��4^X.�+�IƱ>�
:ݬ��4���uȀ�̽Ə�ov�w�?z[=���y�h�'��8+���c&^K�[��ISN��#�K	Fڬ���&��d�pJ�6[jts0vSo������\X��#��'l���J��1g9��E%
���g(�����]������j�Ս^R�o�-*�1��#փ�9�\����ɫy^;�W�n�<at[}u���Z�C���g+��G���ҷ��+H��V@� 8/A�Y@�ݒV%��-�K�RU�R��w�wX���	Eg��\��=Fv�hԻ<�xo�{@s`86t�h�r���{��@�`�\�����fNJ����/L�����M�*i:�+h����Wo�����K�j��@�:������:1+�_#Ӻ���\m�Źٜ��T靈r��͕zSCWX&�M�cY8�����fah����6�E�ҴXp|������M�M5�:�n�;����z�^��ݰ�#ޭOi}�ua�np����&�&9&l�S��v�j&c�Vm;��L��涆���9�̻���lt|��V�(M�	3b&�ؽ��V�[�D)�wO�K�D�W���7{��қlq��O�1��%���Z�ՙgW5)���ntj��(Nڶ-쭮���{2��R���;��%�8�x�D���99����N�S+4_e�\�{	�yJ�ὒ�z�R��s=ff�:*�0O`�b�b]\�m�So6��������ōV`��Qq�]HҋI�y����S���:nwvh�-��Q���fE� i�Fފ��%}���Z[t)�tQ%�^��A�Su�Yu�����5��]ҵ�^pm<&��Sp�A��u��5����YS^D�4
@�n�dӬ�yq��Z���W���n]uɬ�Cy�Z���Զ�)Y�ޥu����
��ESW�_��n�p⋫v:��ɸ�w:�=��K-��C.6]u[7�}g�Zy-9ͱ��!J��g-)��R}/+S'��2���Lc�w;���y���r�_O*µ���B���9 �t�J\2�qF�K��)�RӯZ�����zVep�P�*RXǡ�њN7%c�d,�a1�IY��{,�	� 㮾@�/2K�3x�J�@��wYnQ%�^��gD՝�F�˪6y�����Z7]]g2�㢮B��\9ҋ9�N@;����봾���wM�NYC����{�V�w_���jTdը��1O��en�Z�,��wwq�W.|���璜Z���oQ�VIv"����]�Ԝ�]��p�N'�e�s���# ��������ͻ��3�T秚���V��ڻ�R�
�("(�#�I�uJ�*(*��Y���⨣�."�г�I˜�*�**�
�ȦUD^����"*�K�U�.T)�Q>s�rg��ÔTQ\�/#���N<z�uNEG9G ��.�̹�-��ReTDATQ�$zHD�V]T�*9�:��S�EA��.�kJ�,���Es����H���� �Ӵ���.\.^�T�)JCR4H�Ar(���Ux���Q".D]��W��TEr�N)�y��Ur���(�:re\�Dx���f� �(�9r8\��U)ȕ0���C�Y!U� ����TW�)�ÔT\ΰ���*��
3����� �ADQAΜӕUDA'H�(�TW� � ����S���1"/)C�DUE��D+�zB9UP][��L���
��I"I\9Qp��E�E�
���∊�\�s��!Ap�˸��\.U\��WH��
 
 ������]��b��U�oSo΋�NS�t�G��ܫy��t���Mj����4���:;�A�ķ��Q}��-��濕��M�kٵ啑��=�5^�9�/g��>�a#�d15q��v��s"{��7���̽��|}s�6ǫkd<����j�<�j��Υ:ȣ���k�������7�����@7�3҆����9W��8��3�\f�V�K�_�o��d���hvrC�b�<��h���%e���{�u2Gz ��C#��w�ǄtU b�0�.��E�Bf�=I��w���0���s����`���1��>����fi�u��FS�R�B����>��L�ʸq6� ���=��ytU���M&�N��:��Fg��b��-���lg��5�G|pOK���&�ċ��@�~�\�^,��|��%�c *z���]fF}��}�pиz�E�S�$7��7�����˗�X}=��.�h��><�����'�#���^Cb\�c��\=K"�[��?��؏��]��ؚ&ުM#��[Bg������;��[��ӣԸv��9�o��R�T=�͎�ٚ�>ˌ�E�^&R�U]CfO��b��~����Yp�m�����g���xY�y_�2J�"�>��`9����ʌP}S5+F5�N]w����i!�zg�w� ���Y0AL:Ăjz�ۦa��c7��1����y�O�b&je��5x��0@lX�O!#�uuBp����ٝYz.Q�#��"g45��>��5m>�hH�3�# y�1��'�.U��q�I+��<��Q���� I����}Ĥ|������6�|�R8���@�]��|K��J:��y�F��	Ys���>�^ɉ��R�$���_��zo�<���wc����l:��NC�&Ϣ��T��@�����Ѵ�+P���o{�q~�����D
���~��zv!z�19�z܂3�~;�ч�A��Փws<�X�%[ɼ�^�Ϸ�Ҵumtp���'�ҽ���A��}RG{�{l��Օ�{1x��(ƟR���	k�=����c�Գ����-��T��>���_�~:
�g���OF	Qe��Z��zǣ�{"���DFC}6H��ʩ�v��s�w���L�Ʋ磴�:�tǋ�����9��J'|t	�i���+��?n{�)�|-��Ct�p�/�Yntc:&�SUJ1mz=/�gh5����6�����%���yߘ=�������l?M)Y�ۡ7%P�s*���y�}j��v��q6dzH��u�/��C�]�Р��t|iɕI_�VU0����ow�̒O�բj-s��C�3{^�3~W��\�3���=�+�����ƙ^�g����kp5��1T`�'�b�p��\��=�er�{|]x�n6w]i�K�c�A[����a�$}���(��.w-��PD�����r#�sZ�2���v�tu�cxf���]pƶ��k�T�J���\�
:5]�[h}�l�W;:�͆�'�CΊ�d1���kO�A�H��.>�KϮ�e@��9����yyb��M��P��7sVr�����W%r�G�vB�*���弻V. ^F�t�7��(z�MՀ`joΫk�b���7چή�{�^G�v*n۬���s訨^��U�~�2���W�Wg�9�}��G;%�Q�2}�r��r<��x� �����{��<��#>�lvUL�/=5y�Qʵ�v�k/̣<�-9�c�C@��|1?M�Ͻ�y���g�:������3o}t�ʯI��ͶqmN����n�`>�s~��o��p��	S!;���/�4{ީ��C�s�=�`]th5U��}�9��u^cJ��r�J XR�z�}�]�W��U�4���dx�]�Q�w�X!�w�>���5���ޭ��ԔY�Gz��T�>1�k���wdmt�	�_�Q��2��#�w[����w�j:�ns0����d���u��G��p}]�Kcz+��m��;´ts�����r<��������}��	��� `��9�)�碶z<�l�'�5UC��o���UDK�����<*~���rBh�5�]�s���n��8�v�3��m7�S�wԢ̆��������Kh��(e�T��˖M����e5�:��ܢ�:κ�3}C�y
Y�3M���YP@����]���q>��^��)rW�C����Y�������o��{�e*�➓�c��٧=�TgA�u�����V��y �o&JL����3!dF�s��B�LdQy��{<F���3�g�8���O�����+��B΢}>|w���F�M�
����iw�����.�\����dlg��qmS+0�v{̒F����}�s6�"eoEۙ�P�Rn���Z�8�^c��!9���7s(mL����{�鑕��G�%u�w�[��T��>��Z��*Ϫ}��}Ӄ3��z7Ի��79�[�yx[at������]��q2� ķ�v�E��Z�؟d�ׁ����j7J<�C�����B����JC�\�O����!��YbD��Ȫ�lm␘6�H.��m�iO�}��_�L�7`G�id[�~�^��!k~�3>߻����۱>ϳ��R��5k͝޷����E@2n1X��txv���pJ��P_��x�xU���je��J5�����sqrQ��5�Vh1"՗�9�����)p����x�
s؞NGcw�r����tK\ն���y������Bw�LvuX��;��h\�ZK<,!|�ɹ�4Q���ƻ+����z����g$�]�w���hNd<*���o\ڟ��X�ّ�ڷ�ۢnY'v�}ݠ�5{��������"���;��VbPL��,�Ndu(_;xTv^�;�9��~���/�xm���z��C��ˆ�o�<��I��t��qφj�繫�z�zs;<|��|U��Ȇ�y�/u��a���7�4�	doW\/dm�y��7�g5���Ė}*��'WkR+�G,��ߖ{=;�g�L����w�!7�^	��t�K�r,p�?l`�cʷ&�uW��E�C�}������:q���-{3��z�z����{���/u���g�[���oFsX�s��)��o��+�����!��IϹ{<o�X'��
ܲ)׍#�sT������G����]bQ[[ ��j}q�|F�w�	u4�U�d5���7��CT�{�mMn��gw3NW�B}�x�Y`�=­��s�3Q�|��s�FP�w*��y�c���>��y4�|x)�����~��������|b�6����s5tP���&g{�w���ۣ�x=k��χo��h���薆�~8�o�������d=��>���Rʸq/q�+�mtN�}��!�<�W�A ��<�{���lx�������C�{=2����Ku#�E��~�T�%����x7R�N�8��"�Yp�DS4����u��N�����H��0v�iUʱ[���*���ˣ##��N!���2k/'`���h�ܕ��5�ׯoq*�Yΐ�m���$�;m[�܇W;ҫS���:��٭��\�X
%e�s���!�޸h[Բ,��6G���D��̗ٞ�Y��U��w]���·zD�"�@S�����Hr�n���.��y�{��i_.q������;�ӽ�~o����M�۷bg r**�-l���ֈ=!������b�\��U��)u=*���g�WG��e�@�yW�-�P�m�����ds�I>�=��B�Q�Y](�gu��;�*���_��;�*�w]3��ܩk��eW����ᝮ�
��㫧�ǖqC=��P�D+��徕;�7�a�^���ly������(�);~ظp�������8�'��2�����=�)���f�f��7����^�NGz܂1��#�v��̎��ݹ�5K�0G���+�WR���������|j�49�����
��,z����ʳ��5��oz+н�\2����O�ϖ?�����}�C?)������<sg}�6���`y�o'w`�PR<]�긣��"<�h�4=���]��ھsj��9��=�qo��o��O��y���H��7�"G���)W�7���*�o�����ӗ��Y/ut�/�^;E���fR'���]ϕ��z�R�����'-b������.4l�;]���(��3��(��+N�,dVp�]�g#�oe,l��Q�ڎ�%)��I7����g�9���ѥʹ:�6��I�㔄dk�m������ڲܳ躬�K�����笽W&�W��mWJ��~�a�g���0z>�_���e��*��3�)R=W�L���Z�k���L�;���u�/ Y�qν���I���jT�=V�Q�c��N�G?p�;��I����xYV�,������􎍤��ג��~YߧԐϟP�$2=�8��/w���G3��\�pu�L��S%g�u4"}�>c��)�6a�cb3v��U��:����Y��h�q^�����{�Xs�b�-�*�Z6���W�z�ݳ����@��NmSaϽ�A�D{�pX�r*o�n���h��^��[5�
V��3�s�����7�mw�}���{��S�z����܅���e绶*n߫����r*�Y��:^�o��F���/�����6�dp(���B/ӊW�_���\��JfQ�{rf���h�v��DMg)���iOo�p��a�l�����o�~c�2!*dd'�q�_�`~u3����}S*,{�f��	����o��D�{9��׭�)�e����v.nD���|�_��d�Ό�~��6l�ziu���r^=����>5-r�;���L����zz�(l�O��z\�x�k�99��F���'�O���L���ô�Qxt�������u��4�*��~'��킞`�@f��6��=�I��D�4ǣ��E�G���T��m1����4���x������m}w�G��v��x|����Q�=
}�+�GBw(_���x}��b��W��X=���{^F���֘��X�?ybR�=�q��L����L�+�	��yI�ے��)��x�3�f����	l]��9L��W�g��]D��nQ��\�A���`�&wŬ����^����>�t���b�;�Z��A��xg����$�F�E�gQ�z��XR��ǰu����w��G�?{.;����=���x*����C���O]e��Ϯs�5s6�d�.�3Q}��6�:��਻�{���a���A:�mOdcu7�������J7�Ǩ���l�x-���m����)� ���Z;����z{����#�����:.�)}�O�1�hw�x���~��}4�-�\❋�J˺�\U6�x>՞���b��õ�;�{˼$�;srSV���4�;��~�l{�/�-��-�Eڱ�F��ީ��߹�/iA�^�$��j��<�Op�pӻL��Ŗ��g-n��+;H�(��R�z�vfu������T�V�:*M�K��[Ǟq��|�@`?Xg�YN<���x`�d��W+C	p��|�����^��������� ۗ��ҧh�x~$~���q�H�n�i��ڐ��̩�_�����q3�O(���o��Ҏ�CN#Y����dP�oU��e�a���q	d^;9��WY���̼�vT��J��榻��j�g�O�DdT.�������/�tT�g�?NB����Ǩrޅ��{>��G}2���d��ݵa�T4V[���>9K�M��:�9��n4/w�&d/���D���0s�j=��ʶ�D�۠-z�Ap�@�G^�o0�}k��^y`+������-����s�,춊��*�8[�{�R:�y�O����6}K@�9�����+w�6; s~�R��d���ŏBt�U�g���~���~l��Y����6��}���ܪhu����ϯ�p�3��c�;�f����Y��s3����7����C"=��_����G�x����Ez�39]�۰��%R�V�!�]���U���\NL�X�N㈵=��>w�ʷ ���sQǽ��Hz=�$�������x}-,��g��(��.�ߧ�n?���-[�T)>�Jq[WJ�L�������X�s=�RX�w�<�<pW��eE��fa�q>�)j��/h�ؽ��H���r(��������0�]̍z�&*��-�|"��Rq�]75�������������&���U�@�$�eoEw)�D����=���e}\ckkd�s5�e:0v��ӳL���&v���7��o���yט��>a����r�!lw�팡�*Ϯ�͂��y�{0Q����Y�s��z����o���x��;�/�ӿx�4�zx<�*d�W��`πS+7kDG[��/1�ߏ�4?}��I���>�놃=��ǯ�]~�y���D{����=t����^���J}��n�o�zok�L�US�zԌ��h{��놅�K"�"�� �Ï��g���^����ݛ���3�Vh<�>bb\�J�e�!����(z�E�;k}@4x������J�י���@C��p����v&p�l�-Qn��L�-�9�re��0�mvJ����Fw�H4�Tzm�Uz�ģ��oj�a %��+.���m_X�+��wk� �h���^s��<���� 3��Wឧ�k�tϣ�y"[�ӑq^AdV\39~��٦%Q��U�[�b/ܭп�.��I�O&�9�a�~w3宮�ӟC�&Ϣ���7[Z�w4w�������Jk՟MoT�0�yF�6�hCS�<�sз��#`��v��-e�Z�a��I)M:����s�uoG�[IZ���S�M����W�7�{��.����z����]�f[�*8��ŕ̛�n۪�K39�Sr��^V�Ԉ	�����f��mót���'gq�+��u�_
9ζ���'�v�˷�m^�qE[p��Ţ!��v����w9�.hc[׸�����jٵ�Pzb��R>�9b:����L���]Bt�@'}�d^�'^�y��h=ə��KI�ux$jt�o^cm]��s�
����5��"�Ԏ�*f8�e��"��]��c糙΂��*�(Z����/��n�X�)^q���%��;���`u���(Վ�*���SC8��߻O]L�V�,e^�uc'ro-ͷ����X]�nX��֥.�t������m-$��>=n���\Q����p���]4���I��OR���N��ݭ�a��T8����vb���Q�^�Z�n�1�[�ŋ]�z��z�5r��oshmq�|c-���ҭ�4��Ԝ������X���g�b�
ȱk|Fv"���T�\.�řz��ͮ����ē�
��Y��8{�+I��Z��l�Qۋ�_g7�R�^��zv�^���C3��5���U9���8�rUՀ�\�t�Ü����q45�������Q�B�<g�l�c�I�H
�5E��]����<��[&��_ujwY��>N���F��,s�ջ�y��&�ɅJ����wYxI(��/{;�ͥp��le �+9��?t��nG��o@ZlFNny8�𬼂��ݲiۚ�v�s�	��!�Y|-�+�s2�sj㪹8�ٓ�E��8XF�4g6DՋ������9cFm+���M|<«w���'U��R�3")`�å2Ʈ{lwun_s�`w�KŇX�Ȼ�,���CV��V��F�g#'F�#@º�iYq.5��,�Ҹ&Toe�ηok��\�]����%w$�[L�LM�����m�8�:D�9|���):�؞�[��f�اTY�i�;˹�1,��ա��-S�Fz�cXn��J8�IL2�ˌ�\ƛ늭!|n���P�`4œԻ�R�fL�+f v�{r�\C��P��u��i$��V��J�LH,�ֱ�5��rˠ"�}ڶ�"�-��z�f�Mm�Pu�0�j`!{�Π��pb���%b����[GCV�55`��E�XKYy�����G9ݬ�"�Ĩ5с�X���>r\W�G�PCl$����FiY�L����A��s�x���r��g%�����hr���G\&�;���}WV�9N-��]z  �KZ*��|�7uPwT�������:��-
')-6.�E�1�
���Y���i�g�YY2­9R�_;9q��%T��a]*�L赾�^d���Μ�?�y�?"9�\(B�J"���Tx���G�UUE\*Q	�U�8�D�>X�EQyJ9s�PE*QÄˇ%H��\,.0��QEp�Ȉ�*�ʢ4.,�A뫎�A(�0�TE��D\畅�reȪ����p�R�YTr���"(�(�QgH�dG*���UQZ�QQQ˅��8TE7�PI�*��4�W"+�h�\�M!(�&s�9S ���+�DEȪ�H젠�x��Q�\��Q�V'
(���eQ]D��U�
*�0��r ��*���(���hNX�zH@jUW#$��
��*���PUp��""T���G#ӥˑp�Qr����*(.N$
*� �*�N�p��Ar������P\���"UWE�R+�\*����TD�2�AAʪ8E�QQʯ\����"��A*EO<�{��|�_\��:���9Y���,kpp��{ë+3:WWGV\3�t��v�f,�;�&.�����ˉ���t�4eՌS��2�o��lm���M�ry�;�7n�������w^�u)�1�س��4n���׼w����F�PCr*�>�8zs�%���5���TcM9�W�������U7i���}���\�F�X�b�dT��� u`��.?����+9X�{՚i̓��g�m� =�;�ɵ�27z�#���aJ�;�;hF��h��Ж�۝����6��/���D���v��}Ϗ�R�r˞��m�9մ���݊I�]!
5���� �C�7Ͼ�V���{��V�����]��t#�C^���~`�=�T������)�%�M*���F;F,�qq�׫N��޷��̯}W3m\{�Ra�u�/��Cؒ��6<i0���&C�j^J�3�wS
���7^*+��ΣBiz)�Ֆ=3V�zFDm&m\�2~{�M�4<	�/�M*�ź��k������~bD�bH�+��@ȏS�1�NU�=Xf�����Ld>�����R��<tF�tX�x��q�ǐ�'�~��D���e��C`�lK�q<��苀=¯*���2�f+r2n:'tF�N�mc��i���\d���uo��0V.����o����bVr��|c�6[��G�7�([f,U��R�y�7�ǠVnnQ��7NAXq�F��j���c�-�R�"s7�PWa�&���^��qixWVs�[w� i�u/l�ix�ʻ^\G��u�|�{�b�o�\,�ʊ��v�g\X��>1�EL�x�ȏ|C�|-Ͻ�lQ�W���r���_{�b��z�H1T�5Ͻ�	�s����g����L��SQe�X�`��.O�fr=�y��N�|����p��g���Lւ��/Y>�����V�諾'�VJ��BY����dz�����p�`���g�^�������~��)E�)�|�] ��='���Jޭ�~޿M\u9�T�s��Ǽ��щ�����t��������E�9�̏)���	a�T<��O��=���|3�~�U,+���0d��W��$���I����]��Ҕ1Z�Χ�����Y�vWϏ�h�Ƞ��뇹���SZ=�[�l�zһz�%~,z>>��Zo�'U��C{h��]��/�MN}υ��y��#h{G*[VɬJNK#ٝw�x��FP�u����829��<����v"y{<�������ns��Z��̧W\ �?Z;���lxX~�����"ǧ��!��w�4z%1�Qy��׳�oz��7���{#���c5C,V&�W!�,:4�Y�u�S
�K�j�t������) A
�sE�r���<�jG�;��=�V���(x��Ά�
Mbٴ��5ݛ\Q8�0]��vq�d3HOqC1�Y�Up�m�+e���폴;����^a�[Nc]��?h�ĸ����~�EA��o�*��W�֒u�؎�^�y.w��R�(d?w� �/�����RW���L=���O:� ��!�Z;����{\�3^���]�<�n����ixt�.���2"��#�+�������*�]�E�O�����Abk#�Q������fz
�,��OJ���ϽDY �{�3���Ù,TyL���n�r=��mN@c�X�R�J�"$����Oq!s��֐�~6�=�dɛ�n<�ȇ��d5N�����R=g�w������UL�B�`3oF���ߦ��\4��͊k=C#Ό��ǳ�e��ZU���Z��o<�&&}����D�|�1X��txv�~�bS�ߦ�缳</�����ze�諼~�(�̅C��O�s=v�j��T4EG��2?:��������3���ui'��O|R���o,�ڍ��\�Y8�9�]���<
��Y�f�t�����:���g�r���0O.�)�'�άJ�I�o��^ڹ�c��M�D�ёA���:�Տk�T�T@�5ۦ૵{�Zܩ�b�,�?d��_��yL��Hկ��2wF���`	�^��N���5�t2��O����u���=\~K ��}����>���5ث�����uj����.�WY�Tko9J���S7
�ٵ9k�x�Z��������X^")f��g���F�d`.̊�s3�%��Ii�^~`g��d�	U��U��pߟ�����Ov��T$A�{X{�챞��Ǵdo��ު��p���6�g��m���9{"P�����ܪ���Y}|=�/͑:G���c^;i~�R��\���}k�E0����~�;��/��k��ʱ��q�c<WauG�W�/F����=���5�:b�`�o�����ҭ,��}�C��-���x �"<̫P�v���ꞿt�j�����\F?s�;�)�@l(���r.��FQ�s�s�\�^飙�9Z�x�S���'`�k��}�^C�=o�"������xB��ݱ�CU�nf��ḭߴ�έ{��
�Ͼ�D��P��m��K�쯼f�a��'"��;pyީ��_vs0����'��g0T8�j�%�놃��)~�����Z5Ӳ_��鞀�x�t����{L�{�U������`��>�U͆�Hͦ��z�p�,��~Ć����I�l{=�����ˍ�J6|��ge�B�۰�f[@r����:��h��S�dZ�!k��5Y��N"�՜U����'��{�����ݗ|��QŖ�f���(�v��������'a@��G�uq��ˇ4@�t6�N�q��O w�J{��l�Cx�I9��
�o���b96�Jj`l� ��+Q��:�:1I�QUw�Sڊ#��GUw��^�<�/��ݻ9
@�EB�Rm�����\;���\>߲n;)?;���j����z�V:7ꌇ[~�V��V?v�E��P@����kЭ�?~��V텗͜��ҧǊ���.����~�ϓ�����z�ϕk��dxnT����-HϪ��u���x���
�p���9�о��Ϛ�I��S��N������{!���+��A���x�~_�m���7m97�4/}U�="���q��z�FA�W��!����/]�';��{�rG�ǟ�o���5{�ކ:�F/E4+GDWS��V˸ͻ##���!̟����є�k,����T����m�� ���PB���~��R�<�Eu�܈ھG��w:��t53�Nו�lY]�|��~��q[���ռrȮ{tD�>�$	�F.���_/<�Os콼������5�_��{�s%o��v��~`NF����WI_C��la��6�7@&3�]�
��;W~��ՙ�ڟz2��㖧#j��ڥ)�6�Aߚ�x��;��=~��OqOK�
Ro<�|L��S��(�Qۣ���N:z1ʳQ�Ӵeк��zP��5ݸF*�2��bv�2Y.t
T��C�d�GvQ�u����!�ƟMPCgm�ټ.L�׺�m�R�9٨�I�����f���]<z�[һ��NMV�%�-��ܵEW���j}'M�o��2u�U�>�{!0�}�p�2�kb���p��L3~8����y3��O{�,���7�u��S4�WL�Ya����zF}��z*Z�,�lJ��b2�~�������Hs9�����=;�]t�߸T�c���wSP"z���ާ+=�X��nכ*3}s{�q��Ebc��tW���=�OS����b��]N��Z6������j�8�yp�*3�j�6���~6���%�{�b��{n���!{g�l
�~���ۙ��wz��6�oU6h�D�O�޴��Ԫ�Y�!ǫfZ���_<�V]��+�>w�wN�G2������x]N
�?k�fx���?'�9���S��-�_L�w�����Ǭ��7�ŻQ��>��t��ށY>��oX�g��_�X�������;�EJv�hW>̴�+��L�<�f}/������$��7���mw�\u>��N}�g�]��^���xv��:���TG�9��F|�ّ�c��g߿T��m1�]~������#k��?�|3�/�������L��0���{>n�X��|��]�^�k9�7ʒ�U9���٩J�8G(M��ʅ����p�z<O�aO�s���nDo�]�A8��K�-�ج��--	{�Hzs������榌��]��)���s��fInt��[sdS+�wOx<�ͣ�aϽZ��>�aG{o&����FD���]p��O���ޕ�{
���c'Ѿ��Ʀy�s7��� `��8_b��z+g�Ϧ��7��{#��&��7���׎�X=��\�Y��Φy�Ys�;���25z��#��p|�I�2�/]�.��|[��'����]a�[:g���fCͪ�Vh�Jc(���~���S�d��eLX;�������Q��ƭ7����Y���*�T��nf��F�'^����y/�<�!���ـ�%;��=��4:��z�;"YL-���m��U2�����E	��2�x��GM��z���Wf�4:�rk��^��6r!�����x�����hV��s�x2���u>oނףc���-�6��@� �}�~�o}�nr<���ǔ�@�w�g��=��лՐ���Q�韒/2'�|��
��Ț�E�X��y_�l�=�P҆�[!��ޥ!��&zn=������U�0��5�w]��iU�13�]益_�!S������v�C��ȼvs���!�U���d\���w`-[f��S���]�˔�fM�^�/+�����w���$��!(���]��VOx!ۉ�2X�W���G8묓��%�Hظ�p�YS;�N�
�����[�/��35�Vn6tt��c�1����ʪu}�)̸击�rQ�S2��eKڧbzzQϱP��G�lH~�aU>�M��e��'�I�V1j� .>���t	'���ͽ���4T4�rz7�'�K�M��5h�t!���H�N{�wSQ�:8��o��2�!���V��'���p�^��lP�+.ȍ���W���
�  �fwxc⏲z���v�VA�>�N�N�}���w%V��דxՉP}KFEG8�M{=��]W,�[�p����g�,���]y��f�K=��^�NGz�y{.�`�҉���-\{���Ҷ�4�Sp^�\8uA���p�z�p~�i�39�L�?V�������)K���_n�~['��н��C�vES�C+����d,�Z���w�b�D�^����ފAn�	��Z�7]��j{��O+�#�|�*V~ȴʯ{�իc|?;O�֖~Q�Jt#�wR9��g������}%<�~��0ߵ�y#a���t�X;����`W.�1Ў�ؒ���ݩ!�#�T���w�%lOSc�b����g����_����j��P�O�����~�v#[C�����ǎ��Xؙ�z��;����*�<	g�/Q9�oeӴ@Ww�R��MX�ֵ"����]����+*+Y��^+ή����9,�mB�Lx'Br�^�c����C���Mwm����p����w��A�ND6�gB�I�XԷ��{�	�7�Ͼ�^󭎺���d9�_���M4�<��r��s�ϫ�ױ��Y^�뽋�{�x��7��2e�U����+��놅���l�[c|f�(�	�۬`@׹v|�r��WXA�H�:�:e��
�n�����j9�ԮC�bC���dF-������xz8��8�=�v=U�&e���m]��^Cb\�z��V���O�3-�k��{�PC�7�~��yu\@A�{�*o�n�ʉhq���z�`�`�l����4kgӖ��ܭ"���"��CO��}T���z��Uo��ed?v�\=��� ��ˆ`읚C���`��/w��#��X�4�;S��N����y���|iC��g��H��{�ԏ+Ɨ�uzqE+�]ݞk�z+.5�m�{�4p��5��8�M�yz�0�Φ|q���t]�u̽��͋';�W=棐�j�nU=�+%xf�\<�z�F|C U�d?ow=;���bu?��)f��ש�⣼d1�]���V�>�\�/ðŋ��ߕ�CkU�~8�}z���P��魐=s�+T�>{fo�T�J��Z<)�����
*�gRъd�r�}�����tk$�@��З��ai��5Q�*�m')�]ؕ��.�94�K�miā�����i��q���lۨ��Wt��w��x먤�qU�fڝy��b�n�n�[JA~���o�'e���Mt������w_���ϭ�-zo����O-C�<G�J�5�1�ҕz!�L��g��{�dk����,�Ȏ}�Dy���h{G-��;Ն;�����g���!N�z9��{˞�M�*5�hu��߻T��f��/L	��\���Vs�{=x�E�$5�z{j��Қ�RǢ|W��o*~~�<in)����'�~����}���=��n��	�J�G�LY�C��k�^
(������I�������R��9Y|�k�s�:q·�^_�M��WVXs5m�g�I��m\��,�g먽�����ܽE6����>^Ǟ�;T��D�A�L�Ϯ�h*D>cc��W����o�wl,����xI�i�zo!?cb6#�U�7Ƈ���y���p@lLOK}�ڱ�������T]��\g(�Y�H����S�=X���^{�Vǫ~[<��@��e��;�8���uk6��2�n}�D�zT^�� $;��pݤ�;�c9�������/[ϟ;8��llo���66��01��0����� �6р1������1���L�m������� �6��01��3 co���x`cm�|�m��`cm�� co�����1���l�m������1����PVI��L�@5+�` �������n���UDHA*���A"B�EUQJ�J
���!%B�$H�(�B���R�*�UW�EE*�)!Q%@��k���2���l��m�5֊J%kjͨ��EH[d�U�ΨOm^ڑF�U/a�jWm$�P�;f(�i
�+C��͡4F>��T%V�ͥ�2Z])B�	T�JTu���ԩ*��V̠*��$�Z�e!#U�R��PD
Z�+�T���a�Md�i�*��Z�ȼ   �w��,4z;��Ws��{�mws�q�wu����{��C���{׭^��ޱ�{k�ۋ��W=�V������v��;ޕ�s=z�z����s�=w��=$OF.ڤR���l��_   ���J}���g����z�ѻ��9�ݽk���W|袍3�j�G�������� � ;�w  � �>o�� tz:4ts�X�GG�@h ��ѣ�@E ���e%�h��3m�.   G`}���{��n�uW{�WW������Z��kƩ�+��{�EU���[�bi�^���n�Wy�x{ل�^���l��ֆj��[oI�B�EٕSv8;-�[D�   6�ϳ�M�׶��n��Uֹ^y�S{vZ��3���d�޶���ڗ��3T��wJ������zt[k��.<��{��{�ە��S�����W=;޻�Eu��z؂u�k���-�E�%־   ��)�;w�{����N��S]�t��y������U��י�����=���Ҵ��9ꗳ���O{�w���׻���������ڏu�F��͛b�r�랃����US��l�lj�m�*�6�   ���w_c�n�[�vm^���.������u�m�bov��ƴ%��^����ӻ��痛˷\��z��o�7o@������z����n��W���]���u��ۮ��mW�*T	D���(�i����  ���_ṇ�[��׻r�*x=��]�n������[�v���omӯx�ݻ{pw�wW�t��������n�S�{�u���Z�v)ӽ�g=�w�nٱ��E�{�3����zl��сY�	ڱ)O�  ��w���n����ox=�=�{��W�wuk��{nz��u�y݊��½�����^z���of�z���Ww�{ۊnz޼�ǫcIor��{jK�Gw+�m��C�Q ;b��:��"Z��   ���/�5��뺝�s*��l�l��n�G.����w��qv�m뮜�=�m�������@�S�^�붻�������{z�;�^�t�{6�ٹ禔h��{���/Z��zB�P�Y���a#�  z��}nƧ�[��m���Q��o=�أ���g^��۶�s�So6۽����^��y���ۣ���S��/{rY��z��S��{��`v[�닸��=��.��)�4��JT @��a%)Q�  ����R�'� �)� ���d ��ѥJ����d�a&�)���*FM����_��]��UK�����{������zk���}��}�:�	!I��	!I���HH$$�	'�BH@�?���$���HH?'�������_ח�o���Xu�T��W2�Q1�Q�`b�C�VY��in�e�&�ܨ��"��4*`: .V�"��W�$�{eS�-�����H�w�Z�'++7�Z�w%�ُ%��tܦ�m2�`R��Jĭ�i֙�=_kɯp�Z�kq
X�i�z`*�F�B�ӬK��3s/3ӹ�LS�B��^fP8�4��͔lY3eG�u%�u�4��yv��ɀQ��T/B�[+�+�uQ���X������+d�A�*�2+#5�֚w��q�:2����5z�i4�Xа�!j�7�f�&����Hi��47
:�Z��P�&�� b�٫9+f����(,�vhGCJ%K� d�X>)�<��ѐ4T?f9�g77O`5�I/vX����V�B2;�5r��v�`l���V!P൪�\��2��Lj����ت;!;!�ݻӋ2å�)�3)҈,e昶�8�в�،P�xpҒ�F�!�&�ԐZJː�/saF��b�Mc�t��'�+��7�L�[� *��K�VK�X��T���4�'P�.v^�زÈ�#v�p�ř�ME��L ʹ �'�SƊ�3�u������֝��n�H�E�˄�V�\�+Ğ���4R��ֆ��<�+i)�@����˙�ѦU٭�2ɶ�`<��,݆7y�O&e\��:pDZ��T������Ҳ���n�cŒ 0�4e=��nhs&�R)�͑8h�;/q8M�[�d�V�QOsV�.[��g^Ч������vDR�n`�ٹ��-�V���;V/A��Z�J0i'��1�U	����jX���eZL�!akp���xJ�r�(��.aT�$r�G72�V��x(U�g)�u����ŀ�ׄ���a2^5]�� Xt�uy$��eV��(�:W��5�r�����0�6���7ܼ�L���R�рQ�+�5$n�SF�����P�	k��r�7���Lц���K1\���h�mH`r�{���ִn��,��=��FIZ��-�-aݵ�;Y�^��%(ݬ�lJ���D�:�r\�2e�َ�9�����i'���/lP;.�qn�u�70����b��h2�i�kI58!x)���X�bؗ&��@t�j�|���1���0��ͼ��]&@j���{R��P�5���j��ЬKc3c��a5a}��`ʻ�����v��*u��t� �Q���d`=x/tn�רkX��E:��Z#j=�ml�U�юhL�.H�z�cĪ�#d�r�5�YB����e�Vɷi�u-�{��!f�Z]��sE� \_	V���ͥNZB@Ej�.�,͉̑e]K,�zIB��q�0��%5�E���U3�R�Ÿ�Xq,�v�߮���<�M��`�V�1g�\׌<Ncj�ucJ����Ց���0;L�kɺ�x�Au�d̏v�b�#U�i1���.�d0��e���Ȭ�SFVe�/l+��ٛp̖�T��ی���{`�̥S�z(+R:oBuw�nYu�|��ӫB
�ܰL�cЕmع���ڶ�����ygmn`"T��;�`&��
-TZV��֧E(��tԬ[EF�MZ�Ĭo&�{p��yr��m��>C0H*���9�v���Ԫ�HGX��(��2���L��YoYk5���ېأ��tmS�&f+ҮEOT�q�V�7u�,SgMԾ*����a`,w0���P���_`ʸ���[�6h�o��\9KRvc��n�Rh"�J���Fô��[���cVR;+n��9j��Z#�lG;Ik�z����YK���d)�]:�����B��f���j��w4M��$�yk�+Oۏ�F�c:��y�[ӗe*X�p�T�xʗ���B8 ��CbP��X�Y,M��5��{ �aeZ���I�h�
Af�[�N-̱X���d-�ݡaI4��U2��O5n�-�f��̇��n�Xؒ���/d����-j�"�n��iN�L2@Ē�ṻ�C�Am�oB�tS������L�X׺���Je�m�.���J.R̆�{�SY�n"����0�
��FՊ�4p�	�.���)�J�+�9��v��̽��^��?,jIR�Q��M��^�@�L��l3��:�2S�2��oaW�4Y��j��ҍ�8�PƳU�f�Vc��B��Ů�ڐɢ� &�v�t��ʒ�U���.U�)�X��.�2�MZ�Q&�^�U���!�\N{v�8�%�o�����$i��v�]��1����du�-2���5��L�X[0�4�z@�ZeF(�"�YJ�+n��-�F�FkS�J�`�DfLua'�V}�a�w���j���E)f(dW��n�l�Y��ZHn-�C���-^,�i�.���[���L9��S�hJe���b�H��i���̚�j���\BE��nV�/-o�BV��(G��cQDm�W��	TZ��wb��	�r�YnQ�ź��	��ւdSh��c�KB��K���kYYs�9��q�o�-���B��z�]�jK�HӃoZU1Ad3�1�>j�]�jou7Lv�Kr�[n��;t�rKq4�E�cwt�Y��Wq�M���<�ި�Vk�ԢZY&ҫ%�B�g*^�)x^��WH�2����[r�C(�맭Xw��W��w Öo[@ޓ�X��n.�bވA10�\t`�1���B��#ow~!���Xܠ>b-�nd�f�V�%P�;E�p1tT�&eE)2��9X
b��6;�=�D�A��� iR�sMZ@��L�`�Z�M�ffe�l�[��������Qb>M�2���"MQ��Koɘ	���@�ˢ�m8f�v��b�fK��.�����À��-�z�H�X����s6��o˫���WD|�r��4*@A�9[d�@���5�^�s����ы��v�D�PK/��]
U�2�̀+-V6Ҵ��m���jWOP�&CK�VKr�`ǖ����5Ry�5�A���x��0fk	H��k/mJҲ]��)�@ 7-��@��6�Ɋ���p�S�CtĭN��
��3Y�����7^F�!���d
7z�W&L4�7*�I�Or�S��n���T�b�J��V^e$��e�XV^�v2�4�0U��i$�IЬRf̓X4q�"*��f*	��]�VT�����1e��jȡ��Z��x�ǘC��vӊ-B��U Lf�?,I��%��*��{Hط�����m֭�6ۤ�e�Z�n�@8�{�0Z��U��d�n�x�ZCʃJIJS���ᛉ۱,�uw���w�0%Z�K1	K��,˰��*kn�8Ϭ:�PR�b�\�X�%bL�R��G���}�eiW��Tv�)f��`7��fV*�ɡđp��WxBv�f;ɺ��m�"A�+Q����e=�k�>�/^��q{H�,��v��+71�#<��vJX�9�Me�A(�;v�e�-i�)���x�a�X�{�0� Z��S6�ic `($��u('X�:�X�����䧏ṿqܷ!#3!���(X�ALӋN�1����VM��6�餦< ;{�譡�sX03�T�(c�Z���Ҥ5�6'�k��iޫ���]�Z-���Ϙ썏�u"�#JѡwKn@6�1u�[�*���#+)�e�F;Kf]��-˸�fd����A�r�]m[r���ٻ�)яi0�Zރ��zPŐ�f�6��e7R�VD%Ab� ,d�(�0������!
���BM�e�oo��V� 1�"e�Y�Q���̹Q�4T!�Y�Ʋ6p��ª4$Fe�̱��l��@�H�Z�N9]�qK����9���FJ�n�G9�J��\��A �G`!u�Z[����*&��C&�ș���OhnbH[ziR��"�[ۥL:�L��/m'JdX�4Y��,]�+\;�ٻɷ�]1��N��G盱q�]n-��(ڂ^J��`C����lC����2�jj�E�Mh0�Ĥ͊�M���G	Y�QRX�B�;���J����a�%Z���0Y�[Wb��D��]�d�z]���D�R�,�B�1�,P�F"�ݱ N��)!p��Kl��C���CX�N�zJ��ot�B�Oq��n�y�E�y�5-��GU�V������ʋ.�Ub�"�J͎�]��cM
��Z���%PW����Aɘ�%WK�v��;Ѐ-Xb�Ո���n�T�.<���!��Tl����Em�A�Y�Il<n�ƶU����3"wPX�z��j�AJ��t77�2��jT,hެ����U�t��ǂɟ`.1!-��C�)�k�@"�@)�����tC$�b��i�go]fVj6��q ��1����'3@�zT���]kY��e�Ǣ�С�+Y���K8�*Yt��	b=�,k*ږqƶ�1�؞U�,��k�lPұ��X`��Vj��fȑȠa�z��ݵ�m�bkj��[%i��r���W�Lǵ !��d�Sl7�U�j�H��7w1kx�'e&���Yqht�j{��$&� &�)'4e���m�wՕ`��:�}�`�YnL�odAfad�N�JhkeH�[
ӎܺ���e]ele�E6p�e�(�0�O>��Q��>h�N�e�)�%=��Kܫ�db�ڧ1��btS����H
je�p�l	�-LP���u��ҌHN\z"�jyg����5}�xuQшS��팆��z�LK~�� �g)��0�)��EB�^
�T�U�Ï.�/T� E�0���M�%A7m��Һ��/6��?b��%!a�FK���x7��sU͊QL�tӗ"u��B��t�L�/*Vb` B����mP��������՘z@ue���b�r\r�I��0�mY��kr'�b���cb��*)���ٮ�b�7r�&մմh��J�+�^m0X�[��ˎDV���f�@�f�ܕ�ac�:��G��A�.�%��7	IOiP��1z�6E<1VnI�NVF؟+Qϕ�Ԝ�J��Y�ګN��;�ok6��^����j���}������X���hf��.�	�ک��Wv��������0ַw�[L��[!������ѪV�8�6���Z�@	)�8Z��Vki5�+]�h5���L�6�fP+4K�4N�.�Z��`�b�n-ۊ�c�t�5/E�nkh���ФV��ǹ/&];��^(E�w`� ���b���V˫v�+�u�����1HiB�ˤ�܏,a%��e�r�&�m���jg�{t�QT]è\9�ݠ&ne�TBX�]��z�h �ĉV�V5�H֡�TCi�:N�D�=���8��ڳ�Uq
;��
�]��EI��:��4�L��$sB�pMf°J�J�G�:uq��-6�P�dR5r��,���Tr�%A���ܴ
��֓Z-	��Z��D�T^Ө�+X�]0��#�h��cp�m�aŨa�`C���G4r��xㆩbj��FY��֜�"ӛyv(�-��l1�* �q,M]Y�F�f[XmV@ �m�2��İ�4)2���s���Y��wfJ�C��t �E͹���	i�(��cŸ�p�fj�v�e^-��b��ͰU֓�@�7�GH^y���ܔ�h8��Od6ʹn �jo0m�5�f��jVۖ6V��[�o!��7Z鲱��t"Q1oj�4�E���B8�5V*�ǦK�.ɕ&0��*.�a�M�ܴk��0����6d���� �DP�Tq�t��]�`K +&��t��F4Qw�+��U�U`�*VŚU�Gh�+7B��Yە�k ��Fgk�/�j��2�ڤ�ࣴ�*�A��� 7�w(��R
(�^&�T{�*�&�9��H��ɰ�p���+-9#�y�쬰�L�4�� ǎ���2~(ej���G+&-B��&�(M4Z ޠt^���r�[����ɭ(�^�w���P��5w���JSn��s6`��%7r����Aۃtn��W{���� X����,�{��I���Z��rkt/��ED��wR+�B��'�<����('ׯ�S��Yh&����7,`.�K����V'$n&š[+E��4E3ij�a(0]�����mj�ק~IVU�Zf�?�V�h@GV��.�nfa [(��d������F��L���2�oޱ[(÷��#B6��3Y9v�99u�Wµ�b���סZ�Z�:pސ�+�W�Щe���ؽ��,���7J��U25�a��E�M�^�0�,�wK��MƎ��J�[IՀt���Pܧ[�7j��-^�^k���i��P�ۍī��֋�.�u����#\��cu\I$���%��ɬx�*r^����m�w؃J��^5u���-jS�I(�R�jF��u��[{b�',��V=���55Г�C)Vm�Y�E�Qވ4S���4Ab�cRPZr�wYX�����M4��oA���u���f��E�~��-ZĻ�p�n����(�)��'ʣ�,��y���$�R�kK�5D���j׋op���]䂜�V�Q1���;E0x�$���09WX��[B\X/LH��p�:�{Wk �� �,��U�4��C+%��7��|�i�n�i��v6���W ���9N�8��,RD^i���Z&���Q�h��eX��Ծ7z���B���������� ,�Φ.�a�K�#p��N�Ȭ���j}��H��B��dR
�CR2�]��ͥ%�͜��<w�^9h=�[�Ҁ�RwT�ӱ���u7N�s��\�T������wD|Y�	H����8�n����rNc^�b�Nں.�s�@z����Շ�z�"��.�]>�D�f�5��lDsR��f������j�\J�SA[�2�Q�b�;kjd�8�8���!=[��[�}����l��$�p�7����⮬�/Q������w /��|��55:��\OC�RO�#DP3��?o��(��=E��#h�Rݧ�+.���dd�)����7Y��KyY�����ʦ��t�\���:҈g��v�A��]S�����e�Q?^�<���,�M�т*�[�A�m��z��P��3g ل����|Ѣ3"������XĎ/o��W�ѽHJys��b����N���qEֆot*J������YԈ\�����1���n�#��Y}Daʻ��[Dg@ �4YJW�夠���/�䒓5Ŧ�5��)m�6th�e�F����:���-��bǶ�k-']ti3Awܚ��7i�V��˒\�1��{b�(l���.WR�ᲅ
�Z�fBI�wXt|��׸T�e�H��4�'daUt�+#���.��;�����{E����u$��E�;���m�f�� ��h�t�o�k���&V.�&i����T]�$�)�Ρw[r��b����[�q���A8���vp8���_-Á�H'V����4dZX*S��'3l�Ыu�2��F�_�ܚھO��K��,5���w��T(1�z[��D-�|��G�`=p�<G��SPV���}Ϻ��qo\[�a㵶i���хjpSh��eerR�)��)�D�y�;�g	I�i��vc΁p�iv�`�p��e�OJ�̘;+\�#���T9>m@����R�鼀
A���mu�s/1�d�)IN[�ײiU}��>; ���.�K��բ���^CzX��RI����Zེ�����VO���Vn.�R�����L'rJ�J��e�=����j��v^��P:����y5��bK��"O��ȭ���%}^���d�6mP�a1f�	d(]�+**��Z�n�S!�S��+ђ:.V.
]wq|0�]<�/�Q�U��Wխ�ܚ�:�����#��"�J�����f���8*��������b�$r5k��4 .F��;�]ک�VfS���˨b؞m΋t��8)ݢ6A�;��"����Υ�r��&s*��]W$Z��N�:=�At�vw�h��.�34m*��2�r�[�uH�@��,{ъ�A�N�A0̷e,�a[��uj����}݇&��g`\�H�ʶ�oT\����3h�	'�]%�X8��c��be��3V0��"�����	\8>i�{r�7�?���l�:���z���o��`
�!7R�H�1�ޞW�9���:~+��Sj�T�n`��)4}�<J��q��ҭ�fY�n��mV��r�R��
RQ-7%��Lu$�2��~C֭բ��j�F)��t�!�W=d�|eIʓ#���/`H�����4dh#N{���o�d�Uc�菤��K!!�ޭ�_^41I �"I�A˕������v�z�����-�EZ���7-��2��U�����m�p����d�Kɷ�ѭ$?�U7)�~�^�c��W:�VK>l���F�^M��[�kC�ft�J�d ۾��h�e�����ۯ5[����<+ԝ�V]��˳�q
��@�5�@;e�{����c�m.�je�<�j�M-xm8���.f��
�5��!�p�=a`s܂�N�M�L�c�[dM|C)���ה/g�-�G��0:�	1�θ��C��{��x�-�e9�:�9�-�ץ<�.�E��c��S�������,�*��,e��1�aꛯ����;xRG���PO�V�U��3:A�<1a�_[gS���oz1�>" -*ݔ�p�u�l<��fެU�u����`�V����Tt���Fb��wS�\��3O��p,��gn�:v�i�LJփ�A,�c&M8J�ch]�T����¢��1m��g]W��9�R+��k%T����W��#Ry�>�|y ��|YW�KǼ�^.0-늶�7�D�@!}{8s�ֺ�v���%�|�T��Iw`u���֜���I2|;!`瘇�n���\T��n�/5�U�%�IaJ �
�؟e�v������j�ƭ������v㻪����Z��_u�N�w�Ob�Cy;JgJՑ�.���
ށT�IX�Ǘc��9XjZ�D���K������U����]C5�9An��TD�,�P�r]B��g��v�b/��2�0vK�0�h���iF�p5J:����R�5�t���:�)��n-4��rj�YV8<�FeD]��K�LfJt�/&�ЇV����p%��k�(��̨n@r/����ٮ9q�"%�T�gnoC�`��5�`k�����KGE�@����j��*�Q�eS�t�9-�1�@6�UtE�caZ�\���f�N�w��k���4�"��U���N���B�4�3�ƺs��34�w���*�X��fb`ʻz�K�9�a�Ŋt�=�R�j0P�����3k�]¹���ݔ�-g��Ui[r�heX�цV�v��܅ȯ9�4޳��G�`�B�e�1ֻ�B5s����ff�̭!����mM%���ߍf������Z���[䷷�S�MW<�T�0�m.�ʛ�YFP��r��u������ڹьkk4;+[�w͎&�tMB�|VӻX�wd�S�ND�£'��Iz����Tj��D��F�?�%
{�Ȭ575#{yڨY�PЖ�"�������_iq�{3EZ����}��vP
���!Vz�m�7��|0؏���4On�;P�y����;q1f���:Q�p�;����AV��Y9ث��@���nu�;yd�v�wXU��*��w�@��zwe��]���a��]	�p@q8%o��kA�L���j	�%�2�G����58<�jvm�/�TF��\���Ke�qp��N�	��*N��1q�����E١b��DJ
�:���!ĥ�L�u2�K��l];���c8�v�dZO�{��u�)*����P��TP;wW����"���*��T�q57C4.��8#��4Wc����`I+�,��U���&�HJ��\픭�A���n�ݮf��9Cu]pf��6Be���[�Mǔj,8+�p�.�Q^���[+R�ۧ��)�(ъ�Ʃj��n����A��5�oy�tu��^[y��P��#*�\<6�ވK\o���t0����ok��ͥ�Tr֗-����u3yx�i]U����"�Vn����]��#:gB��x���������u]���z��y�ɷtT�	Ȓ�C2�h�yb��X�q���@�Q�Z��5ݍ울4%u�CVzu�����gX�ť��gq�j��.�SP���n�f�O[��w#��;p���bт�ɶ����&y_c��i�A�����&&�i��ĩ �鼀\H.9��������N�6j:Ki0��� y����@ح�NY���x�d�^C] Z�b�w�ǝ�rʇ��3A�E�P�ۛ��|n��ۡ`޺+����E�o��sN��u�ڭ�Fk���nbIl�}��Ҫ��{%�ʺMcu�B6��X��6�}&b��(�����A�������P��F�we�t��{���)�W|��L�T�Ú��D
�L����*�h���)��gK�\�7ɫr5RiVV�B)J�ژ^�����=#"9=�Lq��1��옣(=�r�g]o|b)�5Vۓ�m�*9m�ˠ"����=bG����`΃xt&�vQ�q�f�J
�o�XD����c{����϶7��F�r�=����}}�]Bi���G��̫ۦzT�ב9�ܮc�Xa&^J�(�=BD ɘ���3*���r�/��(���D	�Ow]�j���rF�[x(�е�{6_d�+j����WZ%��u�7�S@���} -^�`&,'F9f1�:���S_f䲸w�2\6<���Tzt���WX�\�W9�u�n��a�G�r9t�α����j�N���(]Y���b̔���t	�Y�[�+��5���`v��:d��cmmm<��-]�{���ėwKf28M�����>�a��~���.�nqç+���w)�2I+;+�M�oZ+n:<�*�[aw!�a̵��f��r�N��⼬��[����1Z�(�ܫ��Ru�q��ut�!���.�6���T� �u����'j�v���z삍�r�m��V_מ���e�\[��ZN�2���,9|�w+���cYf�4�p��S;
���%�\�
��ݖZ� ���ϳ��kY"��	OZ��{;��S<��Spm#ʀ��Qz�1��
��m����G2eޣ+�Y��VG/�` wlr�@i����dn)󶺲���-R��
�]�l4��$���o��S!\���/�o4�AgP�6�]�@NQ�d3C�����؝��V����è�،<x��<�f���3 U�癈��>$�M�y�)�`���.^�7.�G\'f�uъ�J�"خ����W�:�*d,��וβ��ѩ�:�5�-w4����H��a|�A|gq˫ɳ5K�u��	��|7��ͬ|�0�w�M�y{Y�M�S�)�9���Ѷ��1wX��wi�N�/��b�Z?	׎�3ڪ�Dqd���,A���l��ݲ��;//D��hE�s�]P�T3��=�fX#��Rmv��gn�ŏ�kk`��в�5���*��h��-�55p����U��o��{��9)f,u���Z���D5 ����C�$�i�  Wb�o�#<
���nV�����m^������[��;+�"\1V���I���f���Ԝ��7)i凸���+Y�ˢZ{�?�O1�Jtr�^�^�
%���Mmv�`�h��I/������Mt��S5��.7m�3�4�oz�2:�:v��\�ʶ,pE���P�(�lv��B#�r=yy�N��{s���{�����&�Z���®��]�[c���[Y�[��Qg�����3.Hq�#6�'~��N���1A�2�r�G)]�>��[�ؔ�-��*��y�S
����3v�j)W��͊:X���͗[����GR�0.���)<}���	���ԕe�.^�p6$c�௴U�lݧ֝ՐLo
'ntnu�&���]}@�E��F+Z/�"�>��C��6ف�ob�z�H�i����Jz.��6ņ$���+>�z�E��L[��p��`sr��C4��
LQ p�b�!ˋ�#;��oi��.�A)�`�!�!�4���Q�k�z�*�I��f]�7i^���gb�kL�?;Ԏ��jA51޸
{|2��\��c=��3�mۡ�_b��soW�2wq�R7y"]jԸ��A�ʸ��Д<���؛��OxA11<�,5��:�,}�V�ֻ�F͙����L
��16�,�j�[[���QP�;ӌ�q�������2�z�8+5�κ��+�:�1<����P�N��!Zb��@����jrͽ����$c�=���wZ���	�m�vC��&��r����+�x�YLvÑ��y=j��)���P�n�VJ�į���Ov��:�\����7���&26��k���wQ�}�ȼ�Mʇ����ic&�Ky�0�R������c�݃�Ƣ�ǯ�˄Gz:ظ;�n=��t�K�v��\���IkqV�	Ԃ�X��&���e�2����w<D,�6�<�R�0S*�tgr�4,,j۹�A{]&�J�d�h��2�j��A��-i���:j�KVz�ks��n��(���Hk5Z�;c�Pw����&�v�R�l��P��sB��F�'C\׻e�K�/��)��A)�]�f��u�Y|h	`T�AY7�sZh��7����V��m��mt<h곐�� �޹��[cY�����N��j��yO�����H��w�PâZ�{ZM
�O����t��
���;�׵i@�zm�
�����8��s��̷z����ܷ�79Q���jӾ[��U���v@�n!l#n)嘰m���'N�q\6�S��������*�-W[��K+r���bʲ�)�~�-YWM�������[�+G|
�4��1�;S.�H��m�4��2BP��}�r��m��ޘ ot�<�]���m�"[��T���ع�U�&�8f.ȥr��VƦ~^ߖl��atNTx2&	��K2f�uY�4��ܪ`��B]ʤ��Hn�#O2���;֖�ô��J���L�ǳZ@���E�[�h�3kB�3&����r��l��k���z�<��;�1Xwr������zq�i-�,�ZjK��"0ִZ�M�ݼ�#a����͇�nV.�oh��pܺdn�vN��`�	 zoIlB(q��P����w�`�5F�wQ�Է��T�;���a������H,��oq֑���2e��W&-,ƻ�%�oi`f ���S�U���][j����`�gZ(�]/�;hé̹dkPV�ד+h;h�>c)	ر��%;�e�+i��7�(��3�N
V:�e[[�]VR�3-��TD�&� @�ou慸�{V���iknd�����Y"� <]4�V��V��]���e39J޺9x��ދ;,��'�&��g+N��0��6u<�ZԔ6�7o�g���1����^R�PKDm��d�<2d�</&ʓn���*�C�NJ�sa���lM�L��J(hd�p�*�כ�F�#��� ]t�:g-Ժ����u���:� ��uoZ�'h�(�q�Rt�(��'�����������ڄ��$���>as�_ugu��aL.�8u2<pg�I5�,�r�L��J�r�\6����(�{B�'����Onk�3��7���.d�k���K&Ƙy6Au{SW��z�`pE�K.����(���]n��=2��A�z��������@<W�Qr�cV�'n��+r�
ح/F��D��9���-�� kdke�Ӥ5֝�2V�D��dvp�+)� Í�z9hx��A�:ƬC��#�V�+9�
�Ӕ��o-��z�ĸ�Z�P�+�L5��!�2mb��k�\��!m �-5ܭ�̷v�i�	_L��l�Z��v6G��Q�Ooe��zM������nd�ѧ��UF�}��Ƌ�j��괇�Mݶ�n�n����6��-P(gG�.��,"���V����׹A,��p�7�㻺����ح<Zs	�����:�`9M&w��j�X˓S�:hn읭���[Ǆ�ett��H�J�i���eb����Η�.L���}J����Sɪ�YwUp}vgE�O˵Nm+���}g��8ӡ�Z�ێ��|�.�&��Z��6P(�h��u꫁ف�<�N�j�Ojo)\)䍬��t5�	�x��<ﲙL�9v71jx�� �wP
򶓖L�|�L��^�L��S�j�@[kM������l����#�4��M�q��)Ci���S-�!�C�`���Z�:�+u�+�n��0E�E���K6O$�E�,aUTR�~/��/|�	�X���A�y��g׼��c��u�\�1L���k�����>*�A1���y�N����q�����66*X����ŋ���]Gu�Xy,�gR�p�#MnJqPZ�'A�č,;w���Bܘ����;��d*Mn\͍D6����o���Qhk�OYY�Q��ވ	G�T�Yk}����#c�^VQ��x��NU���±_#��`���������.+J#�l#�"���O4�Ǡ��T�Q�s�+D5�MT��F����B���[F�p�4*�uLih{�D�M
7�H�0�v!+VRƅ�3U
�����k\�tL4�b���it8���Ӳ��N�n��Ox�e�	����J�n̚
�mb�Ҩ��Ǽ�6:%Vai:�7VͶ�����b�&�F�|���V�N�3k�S:��n��}J�U�ļ�T^F�٣�ۻ��tmVP������y��#���$������w���!��@��RV�v�N�V�Ѫ�7����Z�UY��ֱ��<%r2�sn[5�Ab�U�]c�[��� f�ۺ�׶hK����gV<�U���(G�4�k�����HF���[��MܥS+/�ve>�Pm�蘚A����z�40�5,��Ɗ���W�7���C�$��ޜ_�/{�*;�.�dx���'t��4�:�v.�{���cZ�.tㆋRZ�Weu���7G�s�iC��6�ݡ\��3J��H��gh]'Mp虓y�w���F���s�o-��@ְe5%n}}�S�h��s5c6Q�ɮ��V(�ց�"�ŋ�nj�#bC2i]*���wF{w
��,$-v,,}���]`���:�%���x�Ha�g	�Vu���I����[�����q#�\х�&��Ea�y��cs��YwI�����ҧm��M���]5F�F�Ml�.�8浲�\�*WBާzD�^��@u]v���`��Hk$�Ni�6O	��-�����F&5��.ս�biԅ5q�	,��u*�=}�=��g��]�,���S��,��� ��._A���Յ3�Si����{¶��Lb����,nc��gU���ۀ
�� q�sk[��aˡ ��8Od��/0ʈ�9n=�:�%����+otE��&2K������i�w�ga�-��+;��SJ�B�5qz��׬VZoD݈+��%�K��S�U��sZװ�m˥;���)Ę���]�)��U�S;/����u,Y���@̩7�����Ұm�hU������"u�:}\��hgqSn΂������][�����0:JN������6�×�k�3F���#�H�}.m��9{զp#l=���.X{Q�q�&� ��.Zݛw��}������1D2N�VL
u�l<���؁ɖԕ�H���H����Z�[�K-��J�CS�`e�r`�o%�yz���3Kw�Z��d����j֛�ʚ%�]z���v]�څ�o1�0�;PX��`j�ۺ�-�}6�r9qa��ΘGѭ��f����{/H��_
*�7R��jj�#î7J�*��9�Y�61�[��ג���l���cG0XaUi0�T�K�r�'*v�.�[��)wKhӋ"w��t�_�jQX��{N�K9$N�g��a���=��Hk�q���.=d0�:qн���[��K����,�%6cƛ�����Ί['	�V�ʂ�u&oF�3u).{���[�X���d^L�K7G]2H��{/.����i��Y\MeE}ա<�8�d�ղ�hG���M.ub�
咸8�
�ە����9��i�abu�3n�:�M*��1f���7n��J��F	����*�ޜtϝ"�QU.�]�I�|ox�V�6������l��6ԧ���:e����x��˲L�ٝ�
�PZ�.����h���2�M���m�S6�^�iP����iv����]5.�5�n��Hp̬<g\'�M���F��6�V;r��K}��m�T��u��B<s0�'ȍP��s;����-t��KNMڜ ����Ɖ��w�+�	��^��tg���F��'2)I`TW׆�ΦP�Y��i.;�7�;��X٣n���EN�[�>���WūC����{r��<���ܝ-ŏy�����V���y��/ xܺ�L�tc3����L�o�د��[K���Wl,�2ȷZ�rZH��,�4!�X��ݝb�0��vЬ��|��!1�'����PJcl%[QǸ:lNgV0��32��VԂ������-b�cw�w]X��LWD��W��ZH��&q�y���,ڐA}�� ,�F�J'A�W���$��Fjp�4�,��j1�I
N��8��l�ֵ,���2�B�Y�h+[V�(�k=y4ǝ7}�-�V���A�>㥚�)$a�t��F�dl�Et�-��Vc�C9��J.�b=�J�����zU��/���F�ˡc�:pv𩫺�Se�X5�yx�]=o���n����`	��`�:w-�b�;��=J��˪�;Q��n��9�u:[�Z.�R-:_m��X9���bu�޻1f
ŵ+kD��KMe8�͐.�v����5�ia	��wy�]C��	<��"��+&�V�Z�ߜ˖�(�����lÏ�V�K � J�wV�7�+�T3A}BDp5�r�	�,P5�i:��h���1XC,Qn>�]�t;yϖ� �A�'�F��Gp���M�sSM<fAUm�~�AO`�a��CS[d�� �k%�\i��)_og${��E���U�N�4�o<��14�`B��L���[<�v�>�(n#���e�%1�����z�[��܋7@�dN���`��W܎��`�`�V�܇p`oKz�ݥ(d"���mZ�f�I�;�����MpI73�akz��0�*��1��_!+��G�s�p��~���`ۂ�S��Q��pr����!���N2��Ӕ[nѥO�{�ƇhٹعC�bUF����,�b�̂�cK��Cz��TF���TL5\Pc����5>�׺a���k���m#y�j���u�Wr8��Ŏ�r]��¶(���mn�)�(TG���S�yf�ܵ[L),���_��B2��k�d���3�R����u�t�Z�^ uuM��+��nE;��or��v	�0�i�(�Dl�K�얯վ�q�Y�yNvGcgUCumI���^��L1|sv�h ^Q�`@������s6�C�b��߳��Gp�5}ہ=��'s��KW�ÀN��������Ԩ���	�1��+' �qe�8%�U^�v� ��3%�m�_�:Z���Dr�f��}�%;�t�36hKjU�����7t�|z���tܧ��g��}b6d����n.lN��W�K��D��VT=c��2�<��n*.���K�x���po&��/`�tKJ�,G8�v�2YI�����=Vd�=��S��.�%\e�s.���]nfL��T�� ���x�u��w
SZ2I���[WJ�wK�Վ����%��� f����:%sK� �0�wR��;�8_F��RB�ntK���
;�N��,�U��[ͷ����yRX2��j�ޜ��;�=�u�qE�N�WR[Oov�.V��$���������R���*3[�ĵ����`E�;k)2��0��(�]B�!��R�NG�wM�v�?�Vf�t��S�IKrﷻj���.Va�e�Y�r&�b�wq��,V�
I	�z%�h��zR���M���؜�j�;�`��V��y{�σ�}�<oE�"�uX��&3V��8%k1��`n��T\����k[X�s�:4͚�w��Z�-��o^�t;5��	�<x��zuFxlR +h�罄��:�.��k�A��j$*�b�zL@��@{�޸���g^�4���h'}�YŶ�c
T������};-g��)��Hq�n�V���g;�m��9RbYg���BM �g�uM�'H/�%���!dT��si�ν͔���wM�wAp3�n�2�z+�ex��4�Z+��-�,A�n�N�V&1�%��dDC�`i�U��]$��#J�n�L��e� ۧ�����A���o#SE�9B�eq:�9-���(wma��
N�`I��'c�V��{ۍ#31Z`�؎���e��/GT�9��*XE�LP̡��r�E+St��׼�v�tP�i���^͡{�q��`�t}e\��.�|٣ӣ;���.�4���R�B+��I\��H�Ч��L�U���P����<���i5+��@�N$E���q���VO*��{^c���{�żߒ�n�r���X�v���y,>:Űf�(\��OINz���d��*��i��ۼ7�J;�Zwb3O��6��.��U���8^���w�/��
�k��	muЧaCݵ׺��5�E{X�:Ո��Y�1���(��ؐ�<r��*�(Q����L��MZ�9a��]�1bb���J�촙�.�IL��(��*Iu)�5�r�J�`i��D]p��2K �Z��yN&,���ŵ��轆v���	k�j`���fl��e��prO�-f��ŪNV
����Lfuf���pY6V����М�A�z*���
�t����3i�V��a]���Av�b�IZ^rOh���� {B}sxj�%,}Vz���75�T9/f�<��]m�IA�.����o<P��q}y{P�*�pꬔv�3��xcl�2�پqu]>�2�p��c�k��ً�����;F�ā�㡒��q�Q��X���Eί7%-%�d����:xÎ��`MVT`E���Fi����'t@d-Fإ[ք֟�I���������e�lu1��0�p�
@v��x__Z���[&v���շ��GZ�[�CmB�O"�Y9r����Dؽ,����7YoW���Ԍ��/E|~���A�4D$t��\r�������{���â�L�>FUJSr�P���0y�)��ފ���5;;mC��`�����ˀcvb�Oq{+ wnt^ޞ���Ǘ����T�Òn�i73]�[z/&�6�n��@iY��C��J\�Y�3`H�ީiQ��	�m�Mh�Grp<r,��uZ!e��#�{ӯXv}�#a��_�Ux�*#{�6y�l=@�+j ke׵�
ުf�%��L]o0�3oh��0h�]�� �S�3��+L�Ճ�c.��3�WdP�)v���Z�55/^b'�������JZ%�����od)q\���	�ԲՀ���2��ǒ���0Ĕ��t�� ܛ�C��v�8�;!;�]qg7�
C1�\�dF���[�t}o]��$�}}�g�[�7.���nqe>uq�Nn���G�z�ΐ�;5q�Ͼ*]ZG�
9�z񹏪,����C�@��=��`o���Uk�(Ԇ�4�y��A91t	�u���+2�6�&�A�-X��Q��c���Y�����<$�[R�U��3wj�	�2u3;�f|1�Ha�}�J�1�l�Z��d@ӻ�a�Նh� �ó:����-����(m�x�A��f�>yS��KI̔����nď�4Ho^ ���
.:���.i��[�8֋�I�)�%����5�}w��W]6��g!�/H�.^_G\�WV;vz�ݣ�,聎���]&6v�*WU9�aˈP;Lӻ�2�Mu�9���7ה���gRx��j�GezT6��5����Ϸ2p9ڜ�t�[���l���:o^��OW} �I��Y6F�w�ܒB��URI��F�U�����=����Ww)�j�P�A�����[]h�3Oԁ��Ra��sH�W�nvB��WL�W3[:�;1X�a���;�W����:�b, M48̈]Jn%v-C��wZ���Gi�V�S�J��O[jl�Y�q�%Eb
����;ͥ�@�v`kéi)2=��cguK�Һ,��5vZa���:E0�$�Ii���tr��`��l��,�c,mԢr����e�[-�;� ��Z5�6��B��ջG�d���uB�d���TZ��(Gf��`��&���Tŝ�ܭ:�8�GZ\�=�{�fa�u�
ī�C#���:�-��X��nT�Y#��m0��Җ��׽���|����IM���ٓ����mЯ�8��s^DVZ�ܚ�l�J��:�y�F�k-��[���l��\��f���Xf>��D�5�"EE#�c�����e0cM4i׼;��=	ٙ�ػ Sr���pL�ܕ��w�	x��ѵaT�KaJ�2{���{�֠BZ���@Վ�����
�1X�yl��۾cԠ���Mn2�WSÝsg'+������9A�|�V抜���rc5�
�y�*�8�/�"sZ"ڢ��"����܍�/I�b�oJ]��p���`Ô�+y�^�:�$���ͩQ�C��_WC ��.ї�;i�g,{$������Ól2��`x*M����or[9�Y5l)��	ѣ�a8��n(&ZrT��rT�y]è��M��
ޛ�aB��6T�il\�УW��S�%���g��vi�����/�tT�Tٚ��
Sz^^��m�xu�Ԛ����/rç�)��9��t#F��tgA2ȭG�V[��>��ƻ�h��`t���Vge�(v�6,��V��m��چ�������������s�*�X{�7�]�@���5n$J�/���!ͮ��/xV*�u���B]Z�:�ke"T��Z�۲��
g#���%�X�Pe�K�X�ݻd���[6(T�F�#��ѷ���2tL!$r5�r�]�ɘ�k�ćs�����Y��O�c�h�l�pmѝM�2�A�z�jr�',Y������7�[�d&jWQ��&��N�嬞�(-�:5Y��-���A��@�@�(�5m�)KV��(ѩY`ƕ����d�-��,K+V�A��kakj
0Uc����T�U�*���U-�e�J�"
��V֕�Qh�4BЫ��+h��D�cE�+PR�K��*�T��(��FYB�U*���nZ�`�L�%J[J�-��Qt��(Q����--j�ƈ�m���T�q�0cmZڦ7��
T�[mR��h�ҔTU%iZ�j�e�4����7X�Z6(6�T�����ԫY�*""bPV��,�&%aj��Hk)�[-Q�������h����A-���ED[J5����\���˃Y���m����V�5�h��ETq����)�CN*���5j*"�®�G"�2�MԵB���t��-���rV�k�-���]R�b�i+��5)Q�D˗W2�EjDV�ZVZհ`ĭiT��,�Ķ�k#F���ܶ+�V�����W>m#���[���o�a�&+5��)�utAxvs�.Y�8��᥋��h�[pkT�� Z�Ovd>Y_��_d�x���m��g}u��W� ,o'��Ib�G�rI$�����S��|� fmrJ3�]kS.��%>�y]WC�@�mN{Vv�2��/�a���#���A/���Ya0MC�_�{t�hK�k� �z� �����$���1P�y?sѠ�E|e�xvV��VW�3�M�).����jx��--��	���{�Y��z�kb}��͜�!���=�W�/[	Եiky�D�􎶽��@��/�hWD�{x�rN�;�Գ�̫�H"��\��MQ���P!���^�P�6�R�DV�.��4�	�������"�V�]b�E�7g�Ɍ.�X>��ᮟ%R���<����̲2����T<<8J�`Nؐ���v�YU��~��73��g�r#��km�۹��-�=������O��!�D��x���mB��y�v[M��g�f[5=���(�\
��^���>��4��3�w(}��������s>��+*n�Ҵ;�v&\k��{rqU�\�Z��n�;]c-�F�J��4��Z�W������;TV�b�;�>̆�7�:�*=%sm�{8�2����g)�Zo�R��o�I��nq��1�����m5] �]A�Ƒ��*kZ�"��]���LlEδ�"�n����;���	��	M>�[�EU�k�z��c÷4�%@G�S;O�����a�S��k��i�ī�=w��t��j9u�_<��F}ί4�_Zx%���k�U�Ԕf]�K��uB{W{�S4�3z[�fk�r[�{�R�ЈD6 ��
+�<)-�^��FLw~3���I_�఩�y@�T�]����i�������B~b��KY2+�T���kZ��*��1Rnd��ʠ��/�rR�~}X���?E�D��ڿxn2 ��\�:�})�jr��5�V�ȣ�}o�ω�#!�6��0e'~�YME^�}"�#!�"��.�	+�= j���U�?6��(X�(�F���@����l���fa��+D�=����dg;�Թ.#q���Ny��]E������wDr�Lj"=Tv��w���j�T]9/4����ӊ�=��.m�%�WDCD�@As�%��K�����]G���Ί�E	({�q,�p� ����ȝeL�K�PQ�`���)��N�i���;�,P�'dI�/�w����v�n�P�u�]�֋�� ��dI�Iw]�}��h)��m2��诌̵:N������d��g.֌���XJq�:�*���"��N;\V��Ӡ`|å�t�s{F��N�3,��Y��@M5
�Uk��K���gU�8~g��]��p�/���ڀ9)�[�p��#�3I���<��;���z�R��ޫA�w���K� ^�X�}�J���.�$�;zM�v|s֖�V��6����O�t��V\;L�BVs@M�ѱ����P/j ��A��(����[�=���e7zm�pn�9$J^�U�X�=K��ߏ�;B�^s\�Ӎ�u���/�a&.�9�Cz+�+k�J�C������t�J�LU���e�!K�zw�x�SS���#~�<�i�n����V��ӈ��,�`A�Y.P^ۀ�����n-ҍ��'iu\�SW�Ў�^����44�Q|쿩fq���S�h{=zih�bU���h��R��ۃ��K�YS~,ʉv{�����#��%���a�Л�=���Q�u����e�����}^fe�Xʭ��rp�0d�be���	��Y�8e6���B��^���<F�ˬ����.�]���yT����G���.�K�P��+<^1F��8��fO�WV�
�;]mU��������\@�]뺥a�� ���«��1M�#�:#ϯ֩�՝۶���|�F�BW���%_h��ϔ{�x���z�ޜ�3e�����)zz��tSߧ��0����4������K�����f�X���q{����.S�j�x���zZ�ej�߬��N��a�uf��+�_��r��x��"-t���!Q��t�LW@�+}�]�1h�%�fw4%�f�_h��I�U��K�pE�ux;��3"{���ǇmJY����2[s�^�w�8&Ԣ�z��A}[.�yZ��9쬓P�^m�"�2k�oJ���B��SȞwU�p	:��ь ����<o=��V-{$�7�~'@x:WU�/���rQ?Z�6�m��SϨJ9v��9�HGn9��2�=����+�1��b��'���>�z���]�G��?qI.�]۽f}=������Π�V�^tO���Np�^��d��-���W�E:�}�x���$X�ȯ^�Sx!�EtleZj���4>�IN�W��kc��H��o-s_����d]�*�����T{�0���nj�z�Y���cD�m5(;���>���n���Y�8���6e{=ڶ���l�а��n;��U��U�ug���\�6�e
Uhef� ��{v&C��Eڒ΢� ��lE�f�L��܉ӵ˘�U����8�/e6*{����<���,w����9�L�^�>���:u��VS�5�o7���A��Ղ�9���Z�RUH���Cp!K�uy9՟r��6-8xd��&���Ъg�d`_-�����oi�{qR�fĞ��*����}S�9H=_�`?V���i� �����r�B����9>�v�<��d�h�=y��ݝO�R��n�nv�)�<���^��{`h�D����g3�|\�ĕ�)�Ϙu���+��>�w3SS��}PV��4�k��;����<��X#�n�k=hh�=��z=q�ǳ�:������[c�%���s�	yGxg�f���3[�����<�}S>�u�c�&2;�B�M�.{;W<�;��w�ӎ��@�+��k�1u^�����MW�����7kx{��T�:4U��9S����\�=�rа�xo8n[�/�e,�1�҄�utd(M�C#�F�����V�;�7Վ�V�xEu����'�ef\�v:���[�t��`������uгofb����9������ɝ���[h�dh�Jy1�r��73{���>�PU;��/�I�=U���W�i�H��}S�N�{d���^�я1<63r{k�{��OU>Uk�K),���oy$�N@����������~����nQ�pk~����S�+Q� o,��S}�]s�:��� ��X�[%e�a[qI�s��8=�/{89~^Te����o����v/B�_A��Rf�H�oϋ*�S%vɾL����k�ͼB?OZ��>��_b�;~�����-ř�x'ڡ�N{��>�;�Na��M1	��f/
���Z���`M���+w:h�:�h-�cbio�	���?{�9�]����������籌�}/�OG{��7���"3*�� ���t燱j
��BqI��xO��w��>3��Ƴˢ���_H� R5��]�
�pЖ�hj�8�)Q�����KY&�q���;"�5DU�ף5�yXj�7�+k#����hg'�ޭ��F.��g9��v��o)��?vf��=φ���#�V�^>|y۝أf���K��eo+kak���T��W=����nWuL'i��b�-]���ߞ=
��d��ӻx����Y-o`M
vς���(��}���k�Wu�ձZ�s��-s�ԡ��f��Jw�r�o���54��%[U+A�/O+z��oS�7��;s��K�,��}%�W��ɉ;�g�u(�M	�uڦ�o����ګ44�h��D���]��1	`�<���X��.��`9����1��i
]�l���	��ڡ��:�ԹD'x(�T`��=���=��-�kwٓ�7b�V��|�;���<�B9�"Ou�,��-l���(�0�G<��u�V7�'����vţ �����]Ժ�El�mwN��a%鯹b��d��υ�-|3s�Vc����M�y)�9.va��zf{�H��������b�A�D�7]�4f�;>Q�ޭ�����%�l�,�K�*�9K����{#=��l��[ ŷؚ�=��Fd3CCkۑwR����)��%� ���f;����Nʼ�{m�!{�ȝ���2q�4�����&{���39}v���WR��u�C�!׆�n)���;�فc��ެ���D?R���x���^?^�D?Ez�w��铎��2ơ��j��wfys��Nl��X�@-�a�3����=L����{ �/F�U�?`��=�x�fIv<��*r���������'zǊg�|��Ml�}ڷ7���<����|��ר���Wf.yo^�G�L���P��]��׏ou߹{�=��R"��'���A/��Uv9m�WFWb��Ils;=�sR�	3���q��O� �U�{~#v��	4��g� +�5�=�27��K���E��$���c�`�r�[���{�g��������{��Gl;o�dz�گT���~w**=�s.���8��Ay�>c���ã�U|��j'�g� �S�w����8۲���iD�>�w��������2ov�\�e��M��I��zj�X7n���bp�Y���t7xW��Fy9
s���#DԬ"nK��K��+Y�V^�]�WgB#�v�u���	����:�7;V����_\j�d�VC�}� v��y�����-��{�b�Д�.�\7�i衭�)��6���v���� �gx]��W����-Ğ���޼�h^��;9�6��^�(x�u�ҽ3��w�X~��9Πρ[Ʊ{*��V�_���s���>}[U�����?v��<�X��܇�������^"'+�>�~�tu���������<�5˳��^Ϡ2���c�loT��Ǹ"�y/!��,v���\zl�c�6/O{�
���0�4�;�����b���{H؁�ώ9^A���5r3�=!�Q?{qw���i�>⢩��S���q�3jX}龅�jy)��qο�#��oq����y�ʸt.[]S��0Z��V���r����&�y(�ʒ.7|���M����{g�_5"��T�S���O}J��{��|g��x�z�����=��<�,��j:(͂��g���/|�u_tƷ����c)Y ���7З:LʆŦ��ѦR0�yL�r����Q�oo	��เ��������.�K��`?a|ҙz��LTw�m����ө�]�Obo*�Nv.r����X%�9��K�Tv�v[#�7pE����7}�7˶�֞�.��<�R>�'�rw��|�:��Łg���洤��G�C'�Z9|��.�_�<��"C;��.|M[�'Vs<b��s�T�琱�:J��T�>αSQ����u��\��Y𶑆a&G�Rک�S�Y{F�]`�V<ۄxg3|�䗀�yѻ�"��'Y�G3_1�y*�U��S~���F0�������-W��/s��Z;U�v�G��L9������5��n?	�"{@?v@W�d��L��{���"�w�>��o�%4����`�)|�����:�l�F�f�K�uF0k��7{����sɤ/f��}��-7�Sܾ��y0��mɦ�x�x�\�7uA���|E�){zX���<F�O�%^��q;_iF�݄�s��oA}���o�8��5}Η���v]'Z�>�qv@tk\m�.-Ыg&]ȟb�{Hge�4]�
u�8��fۼ9��D�q�ڥ��ֈ�=V�Z ��b��ϭ�Nao*�1fZ'I��G�!N�Q{
�ͳ�SХ*�f�{�[N�*�{�[ݕ��z���s�[�r��4+�)U���ѨEoO�]�&�7ז�3���'`"Q���ε\��%�1��ӊ���@֥�f����ܛuj�PR�b9,��]	MT�+zq��7�m��Rsgy�N�f���{�����Z��W\��unM奥�\�6%z�s J��*�;vgv�mI.��P�� t퍽�vH�=�[P{y�fH�U6W/�9�q�6�u1��rI
��NEt`G
Fcp�{��LP�n�c��"�0�GW��n3^KK)��v;%]>Ě��|3Ĳ��aeeu���9�H:|+e13�X޴�Ky�z�b�fky�1|2(�u��	w!$�vH=Ww�@�l�WMpY�[¯�з!�kX��N�Z)a��h2�f���R�g�Q&HEF���|l���V�u��M�&��3ag���ε�7B>��Ǫ2��CkW�v��:�K�(-�L�F�K����U�Lo�iMm�Y�Sz@-������h��u��!--T�m%�����͜ã��j�\X�u|��ͼޘE����Us%��K5t���\��i���L�n%�2�����	Nl�cᔃ���UԒ��}u�9�����MS�%ǎ22TsN�yz(�K9%�8U�M�����#���D0��ѷZ!�nXǚ��ټ`Y�7\u��Ф��ܪ[i3;j;��,�mC����5.�qa6�a��Y�kp�y�Y����4��z�����]��!NKHp�̻(O��'vV���̒�$��66U2�'w �ΉEo�&���A{��<(��ї)�'d+8�*=��*�4���_^ө����8u��.�X0u$/5;�%;�w3/���)Gu����~�ٷ{)M`��3���;��8�Z"D��d��y�B�5Dn�Y0!�d�D����}�r�)v�����J�Ĕ�/E�6�&��p["���i'��y@���%�9�|��6�ie��vt��R1}�] ήR��Z�z|�V�"֥����+*��6�.���E�4���6`G������C1� C�����"X�]u�4��=&�bt`Uq�u_�^�7���%�e���m85yV�K6)��e��qH2x�s^]ik�B�=���:���Y�gN<w�m7-D�%��&�C�|����4(�n�_X�����(S�eGq��LW1�e�w����qg��ӑӹn>X)�|) ��Ӊ���`ԩR���$�S3dt`{���������Xw#ԭI�w:a�n���|L��v;��֭w$:�AQ�P�Bq�e1e0:��i�i�gK&�-�e�ܣ�F�h���Ռ�\��	E�����J���L�j��r�֭-K���p�����**V�3*T�֣j�ej��ڋh�Y��[�1�j�m���-eP[)F"1�-ɉ�Y[)mLj�W.���AJ�JT�6�KR�
Ѣ��Q�kkF����uu��Y����Ym��墔��%���X-E���ڒ�0�R��-I���s0�	h���J%�P���PEF֣MfcZ[m�iJ�.eS�m��\���F�KA��P\����a��t�0ƈ��12����Q��C)�"�J[l�m[jX�Q��fj��l�+�j�5�Uj��ѵj��mDm[Z��2�[kU*��EW5�MV-�k[�`����F(�5���-V؉Mf1pm��Q�QdV�̦Ep[QjZ�©iYZ�����uj�61���"������f��73-�Y��+9�t��j�Q��ACv�|�9%�ٍ驲�y�5A(<�֪�ʲ
��-U	b�N]z�u��^�)5l�2Ѹ��L
�֕��{�4B�߸,�Yͻ~��69(��ϼg>3,n�5�9+*Q~���['d���߆0=���S샯��Ⱦz9L�����6&���)��K��տ�����]�,E�9/� %�S|qޝ�[ Z������C9���%��F� �������o�:#}��u���f���Q�R3���\�3���vd^�7OX�u�ϹA�L{V*uح���)�Z��>�BNV2���/b�2N������9 �Ӑd?0�_���G�,w۱���\���lD���l`��NV�.dʡɋ��aN��T����@)��r��E�;����M���G����P���c�u�IU�1s��h%yJ���t�4�b��Hv�"�C��_{t(�M�*�0��@�6�.̱2����5<��i޵>�6�����g�Y�5��r��۔�`D����^m��Y� �
�5��ͱp��!����H]ln��{���'+nh{�n�5.�E�D��\W2b3P�wgq\�Q�n�C��V������Pwҗ
ڎ]-�1���K�v��]�����	�w��LCϒz~�[�d	����jg�*�뻿��:"�o�-��*�iů���9�B�]�:۷wf�Φ��7����>��U#^ɽ�ǻ��;�;��2��&�3���j|Q�ȸ��ŝ9�T=�p>���G�_����<P�#��-��;q��n�.�w�掲.W��`]���{"������+��|�巧=����;=ۣ�Jȗ���/��2jls�ޞg��X�^)"Ľ�kt�9�v'Σ��꿄yJ�;R����dzt��3/�µ��*tm�)Osț�x�38����ζ�ý�s��QsW��&�i�N�����\��Z�_F��v\?O���~��D�s���{��ry�6����K��$}0��c��N��.u�aI]�t���)��g�zŊ}��y7"F��(�-ҝ�x҂M����ꝺa��p��9�_b[�M������Z�Eά�jˣ-q�E��:ݬ|ٙ�mj�Њ�w�?&��-o�Do����F�_wn�rv
��:�Ãu&�Πp�A=��d��Y��pz-�m��-v�������ہ�:}'/��*�s���7�ә)�P>������nԛ:0�~}:��಼�­�cϘ��mX���:s4�W@���54/�.&B���N���w�պJ�GŨZ���k$bYSc ߮ߔ�I�%����m�`��Qx"ھj���f��\�ݩ��Vޫ�%���%-m��§�{h�Ia�z��\���jMh$�\�NW�;x�y�X�7at{��n�v���WѶ��v�,o����bG;
�#(ZM[�&J� ; �.WG�����.�}ܱI�~�X��O�։ko*���^s[�4_����X�-r����ٜ�s��xהCX`R��D;�S�v.kޢ�uj6�;���$A�{�䩱1��ƥ��Ӟ�����E�3�nw�w�� ~��.W�[��̒k-o���c�듕�u�C�����f
�Z�jy�݅����}�^�a���f���n�sW^�*���m&��t���<u*׋C��kve��`;�43_;w��=K�$��D��y�OfP�}JԷ�-K�m���\\{}sw^]lV�D�0�'{��3�����r@k��y�f���a�O�Y� �:E�1+%,��Y���2qM�nxw{Sl�/���Ǚ����l��y��
U�d|y��4��0��o�򷱓�Cs��p�7[NlJ�ם��坘�m�^��s�	��4-��ˣ��=�aҁ���$���He�5~��HMaP�w���ء�^�?��&ה��&����'Xu���C�zɴ�����O�u��<d��{��}������L�۝��$g�V���}�2|�gf��=IXh�0ud�a�X���'u���
�2kT�d�n�y��2Lg�LC�`)�'�����c�"�=�iW���٫� �3�K�}^�I�hi��X��N��&5�C����.���7���$�ٙԕ�&��8�Vf�d�a�Cg(,���}}��1}�gW�=E,����PZd�v{�>a*J���u=/p���,�@�&Z�Hu���9�����>�a���������2o]ϫ����:��v�2�~���R��S�}�|���p��l�gRq����_���E'S��⤕�N�2{hO�,����-� VJ��_�u����Uh��}�ꂅL�S�;k��[��Ϫc��,8�~a���M��&�,���8�&Ͻ�<d�N����H��h�n�1���C䞵���0��H~�g�B���?8�w��Y��Lv�0ϓ�+&��/~��+��s�2��v�>�~���}k@� ��#�Xw�P��r��\�2_,t�/1Q�u�+�L΃n�o[#��&�侠OgSy�=Z`�shy1.5�_��[�n���`ɼ�Q��U�SY�3kh�nw���L`t�'Y�&�q���8ɩ��N2Ol�����~_P���g�0�8��O��'����C��Lf��}R��r����2��[��@�߽gOX$�;��'�S�aY6��O���l�1	������䟲��d���u���n�	�N09i��_`����_�|E-s�^c�����W�C��!���C��p����L?s������E&��!���2~gP�5d<CL��慒z�d퓈��:�I��]��UV��㣪��[?M����=���:��?e��I<C���>g�4����I=f0�߿hXx�|�����<Hje��i��Xne��'Rh�0Y'�7���~s0�����5�|���I�d�{9d�'m��,+�6�OC��0:��rx�	ԟ�3 z�Y1����1��7��2O�g5�d��$7�q&�?"��;�7�����sFw����o�6����I��\ԝ�I����6�!��`Vm�~�B������2xÌ��Y�&3��s	=B��(������~G�����^�+2��m������N�g�?2~E�@�̞�$��y�&ߘN3��|���|��8���?C�d:�Mw������~��~V����M�k��j�'���ٱ����;��(�OP�v�'��i�O9l��d�kP�`o=�m�I����!��'Y���$�&�܇�_���U����柟N2~�:mt ���ԜC�&"��hN�Y3�pQd�CA�N[	�N x��ݲq��M߲�o�&��C�j�m�2����{���J*������?�w�|�������$���P�'����!ԛd�Y�Y2bw�.�N���`{i&e��1��sVN0=I��	�J��7y(f	�p[�T^�W�Zx�ͳY����@��28�L����V�g����)$q�|�0��n���Gy�uj��,c�(v��iu�*�W£��꒑s:�3@_1�h��|Z黅�*3P�0$���MjI�g�6k4�q�''g������`������,浯|��q��>C��C�|ɴ�翵�I�Vq������CL��!��!Ԟ2b,��;����9d�a���|a8�,XT�M��yr���뼿�[�����~��rN2~I���'u���<I�:�~X1���>βO���5��Y']��>d���
���-���u��sY.�'Y;�w�o�m�h�)~w�^�$�C�[C����D?3ě��!�$�joܓl:�nyO�:�hu����ACL�G~�D�'SS��A�Y&�}��-��;�
��&5��߾ӿ5�w��=�@�
ßy��zɿ�����XM3�'�����!���m�d�aY:Τ��rO�m������):�<�����﷗>�����G�f���{��y�����?s�~a�����VO�8���ԟ��&�q?j�~z����N2O��d�C�M�_Ri����^d��u�����w�~��y˭k^{��]r�����7I1�y=~d<���m4�ü��P���u� k,���M��c!�d�l�$����d�E$y���ڽ<ϧ7��,������6k?� k�
�����}8��M��Bq���!��O~;��<~B~9��=C�i�{���I�߰Y6��C���f!<C:s>������W5���褚d���=E$����N��^a=a���̐����OS�'�;�I��'���nI�?j��'����l���3~���u��ͷ�{����8��=gMRI�M�$�&�I֤�>�,�d�5�=�>@�^��ݐ��{C��'R{>��zɌ79�jI�b�?w0�鿷����]�=���س�I�:}� z���I�O��fR��&�������O�<�:����=��0�u;����gs�q��I��>��g[����e{�}�.k��;&D�R-=���ʬv5и@�+%>Ź���S#��P��O$�K���`u�w=�>y��R	<�J������=��+�X���2���\�۵z�I=Y�tE8�������;aW`v$���oSe���_ P6Uf�i����+�P�(_�<ω�
�Ϲ��2N'�E��P�-�I�'��fP>a����I>@��'��q�<��'��{����%���������7�����$��^���aԝ�N��&!����O��5�pQI8��b��P�l�'���E�$�o��	���Ci�	�~��y��=�����y��7�~��Шt���=d�3�߬6�ONy�`~f�?�I�d�q����IXh�(�N3\�I�XL2��O��v��Xm���\�R���<羷����q���0>��+�'�u!�xɤ�Vu�u�N��l�s���6��@����&+5�`N!Y5���q&��Y=�������s�߿k��2��}������}�7ӌ�$��LI�!�#�	���Y���C��C�z�l�W�'�*zsY��I���l����Ms!Ԟ2b)�s$:�Xg|ߩ�}�}w��ǲ9&��ﶇ߿�O��_�J�ɩ�'X���ߘN��!�����Ca�̀��M�^�O�����u���̇�<E!���<�����޾~�_�[��{��I�&Z��C'5��$�&��Xm>a;������5a�$���&�|���?!�M��?O��
i!���3�%IS<�{<�����~u�Y�w_���]���O^��C�5�����2�k��@�jg3Ƥ�d���}Bq6e	�~d�}��q�c6�i�a?'�c'P��s���3�W���<�~�xo5�s�9�>I�N+��wD�'Y�hq�5������
ɴ�t�ý�ąCG/�'Y59E���OƨO�x�_�`q$�޾B� ��~Q�9����~��>�����U['d����:��}�Bx��o��svI��2yl��y��x����+%I�A�u�0�����6ÍlJ��/�ڊ��L;��J�9ۮ�A�ߊ��dÛ�+#,N�7�a�Vn���
vvv��"����i�&w~��(�3t�ݩl=4��ۈ�A)������kG27(ty��]�C��B͐2;J�w7��uu��1���ff�����$��םw��y�s���x��;�'�l���N��l��ԜE�P��Ԝd�9a? u>���u��z���0����q��OΘw�O'�Y�w����ӑu��2��~����_՗U_��C�~d�=C�Ր�5��|�|�s��N"�j~�����k̇�d��s!? u;�>x�x��`q'��A���~`�T_�����r�޺�����[̓��Qd�?$<2��4��3���i�|�$�'���E��ٯ2N2r�I��m�}�������;ݖ��o]�u�o�9�5��'���w��d:βi^�O�d���C�'��(�q��e��i��,*Cԝd�|�a>dѾd��I��'9l/�s��N����߃��y��o}
��M>��hO�%�=g�<a�N���|Ɉl����1�d�'�ѐ>E	�N2z��,7���8ɭ�Z�|��x{��3�>���ߓlvm���p���W�W�����0;9����O���a=�0�~aĞfI�2c8����B|¡�X���h�,�"��g�>I֤�dkj5S�E~���I=�(|��?}�PL�CoRN'�Փԛz���:�xϙϨm�0���:�2~f�?w�'P�&!���`N��k��U�q^o���<�ݭ}R�ñ=ɫ�?���uwU��~@����h@�&���'��!��	��5a�O�������u�xϓ���A�RN��`x� {7̓�m�(U|�u�bU���������>T>4���59E��I+�>�E'X��op��{C�<I�a����m>՜a>a��P��'>����~�_���k�d�=���U�>��?T}���3�'���pud�a�)=k	ܰ<aS�O�I��6�`O����&������4������5�A�ja��C�˾��x/m$�lm����uM�in���,d>DV�|D����a5���^Ac�1L_%'v�ZqD֎���;���;R�uaV�]����#;�Y�P�D=l{7����ɢ"{f�ⷢ�n��!��W;�.��+���?����[q6�{=���I�
���Y��	��_���'��?NRu'��3��P+��VI���$��dRW��ՇJ�5�$��^���;��_�_��9�����'�ֿ4���L�'{`x��>M�u��*h;܇�u����,'y�P?2e���$:�Xk��a:��Կ��LϪ��+���^YO�#��C��=y߽��l��)4��N�O�4��|���d4��.��):���C��Vw�>d�hO��@�-�`W���z���>�Ni�e~��<�6eU�|���f�'�z�����'����Bx͡��E���d�2u'Qy�I�N���C��Lf��>`z�Cs�������S5���t�����n�M��u�V?w8�&05�'�xɶ���O�&���8�<a���:Ρ<}I��E�?P6��:���0'�O{a�Y&?E����w�3�;n��¯V�~�����������R~t��������Y4�l
��<d�8�B~L`j��'�>�d�L&��u���nk�'�d����a�?~�|o܄���p��^0�0�a����z��Y�v�'�N����$7�=a�O���Y�&���z�}�q��=^�Å�L���f�I%��#�'��k�� 8��Oƻ�`u��d��I��܇�8�L?w��I�1�uE��OS�X�����c&�a���N�����c��q���y]�?{�~��Y&�w�y�;l���'Rv��aY:ɴ�w�C�����I�=g��������1�o�d�&�5�d��$5�������_�i���o2��|���Ĝd�2��O�h�3I'6grO��|�����$9�
��M=N�HV﯌��l>d�3 �>d�q��O��.��+�h{����b���5�����Y����Z]}o��M���y�-眞��L�6�lY�8Ԧ;	k�Ͷ��y���W�:$��_�yݷ�J��|8e�g*i�9��D�̝rĦQ�|�%"&�ֈ�S�3��:���hu󤱞�m�����K������M!��4d	�[:��OȰ�e�d��֤�2^�i���=��O�~N�?r�����l���S�d����]Q��_�����B�g���g�.��6��Lg�KI>B����(�N��,�E��Zq��N�"��N0<���'��oRN'�VO���Ru��u�}��>b����?�����Yޚ�{��0�y�C�CH�rN��LE;���g��E�qNQd��L�qğ5%�N0:�I����7��u��;�-��)����R���-%�<쇬�'����	�|Ν��x�9�ᤇ�m�|�u&�1l�jC����h��u&�Qd��L2�����7�Ҿ�>T�!+Z��U	X�����߾}�΄��t�:ɦ!�����d�l�y�I��k�x�u�/rd�R�2I�&"��su%I�k%Ւq�Ȥ��	�G���{����w�r�缿����XT�'ud���M��I�2M3Ԙ�X{,�2u5���I���7��,����O`k�����2�h�0�P*y����y�r��˽>{�}��߷�XO̝�@��I�� z��x�f���$�k~�a�C��u��:��ﰂ��8���N���"��߮���]|������<���S�s���������TRcP���+��<�O�<�����XM3�'���0�!��rM��&���m���O',�!�U~�������u��b�L�c��E����z;I1���2}l�P��m�;�@�
�>�~q	�$��4É�j�~gY5��N2O��d�C�M�}I�N*��9�x[�w�/����v��ğ�8�N}�O8���n�b�|���!���ԇ�?&��,
��m�;�'�1Yd��m3�Ր�5���$���\���fk{q���=�KɆTο����U����N� Ι�Xe��������yWE�@-z!ǚ�SA+�ԓ�E�Ec�u���n���"�V�呫�خ�H-xI���Wck�2N�bef���u��`�j�m��bK�/�Hm"5����P[A�Y+K���JZ�{S��c������.R�I]�Ñ�]���븯��}�ۗ{{W[ ְ=�@�����!�]�L��N�\���:����3�a��w]��[L�B��#n����f�k�oʹǫ%�ŜʴսR�y��=�go�2��v𱙺�K�9�f汆�a��ƺ(�&y!�N����k\1������Y%��:{'k8��1�Ҍ�KA���!Տ���W�&[���-N�EDv��؜�
6�itF�����>b�:�*b��I�N�`���ź�<��Z|��Z�f'a/0���H��4;R����e�ǰü{8��ܻܮ�Dl/A����l]o	ϱt�O�tި�)]���@�l����ؠò�Ņv H�7�Qu�#̆�����ˊ�A���O�7T��ƴ���?K�J�`��Q��m�X�a���#9�O4l���.��,����|��R��:6;-�h,S,��U� �f���N�$�-�䬨z�T��<9�B����9�.���}�.��9�=Vȉʒ8���g�W���O1dײY3Kс]�̏��ǹ<��"��E�/\5m��ݢ�,�5>��s�DӮ�coٯ�Y��r� ��wWyb�����6�%b��E,���6�U�B���8�
�\k�û��P��
�pĪl��7�3j�C31M4ӷ���|��P�d
C�g^����w�
�{Mi�%3�D2�+�*;���z���k$�cٿu?����X�L	��v����(\�λ.X1L�C���6�h֥x�^C�%S_v�ڴ����\F�×�.�c�+t"{�)�ؙڢ�g�ÚUu�Z�����i(��=	|�CH�.-D�|)uu�a�qJpO�;��+ʹ�a�����V�G�etUq�mN�I�"�������ֳL�,=���:��L�g��ҹ:@f�1���awjoyP���Op�:��۶$�[.v��4�2����U���P�Q���"8�%`��xs%J�+E���F��z̵I� ��s4a��C%�e���$�Y+Jlx-��+eɅ}���N`4�4���U��KβL/��#/.-�!���{���d,V��ļ�2��ƪo`��$��h����T��ĐLP�WD�Ś����Gl�( GGUfٌ�����rȾ�-*[W�2�����t��{���$��M���#���.���V/Q�'�*�aÂd�h�F�틅�'�`}�Ҥ�f�3p���f��\mSʷ�� ��P�E

)R��Z��6�*Pd�h��J�cjV�2b�����5�[ej�,r橬�`�k,Ll��m��մ�m��Kh��eF����D�3T�-ҵe�kR���Em���B��PcU-mV�D�[JVQ�%Z�+mU�[V�j[UZ��J�R�
�Kj
�R�.4�`���c�q���Z���m�J�m��+T-m��)��ģYkZ�(�Qj�KB�m���Pj�*EJQ�Vڕ�KjU��kF%�K2�lU�e�m�F���*Զ�P�Q�-q�R�ѵ��UmZ�����-��[lT���TiV�L�Z-��ҶU-)B�Y*6��E�J0�*���Vэh��j��m�m�Qm�[mm�V�R���PQX�4�`ѱA
��*-J%j��[�َ
�փ[-m��T��j�YR��+*�E�lj�DR�R��U�b�UZ((5H
��
�(к����=�M��kOp0��0���doz�V��jX�RwXq,�:������,�&�[0��|^肽ib��  V���o|��=�$�)'�_Rz��Y6���N2r�M�u=�r݄��}��'��Oӽ�G����CôXx�?:��ɶ��e|�hu�痕޻ܣ����~��o�?'���
I�&��'QI5��������z�Ĝj~�2C���=N0�0���q'��'��y�'��6sy?$�%��Ös~���h�î���Ͼ�~����i��q�2m����!�M2k}�d������RO��a�-��y���<z�7ߵ!�S�P���79�y�s>�����]k�O�~�P����~7�����,�9.�����ɍ=�T�L�"ֱ~�-��Ls��߫�A�����
������Ծ��vE]�w��1:�H.���t�	��˛�#�4����ζ�ý�������&�(ѻ��d���w���v<�����h�fڗ+>����v)p��R�'w�g1�=?U�o��ä�-�􋈝���t��{5���ٴzJ+��l"W��n]�K�}<��G�� y�4vI�-G�O*��=�zvȝT������
��K�ߪ�ӹP�;%��}��fNzA�w�u�+.�PoLu���q^Ӯ\��o�m�cWc{(�|Vn��s1T�d�ϹѺ�m�`b]㔙��P��wz�]�"��,-��®������Bۙ��37�n��5#F�e^��-��ˬzW1A��U}�}R!�������������j�ުB�E�`�Y���ϼ��%{��dȑ'ޡ�ì�믃�
�p�$��_�]W�U���*��7�q��)ꋊ)��"���Ĝ���g���Om�,3�Q���~5�fL`��_������Z7�7}��0{y�����!�}�ڍ���R| ʸ�.f^�<�k`կb�����;�Dn[�.W����.�ϻ�g3��#O#:36ywv��w��<�Ʊbs�-���83��¶⏞��w�Y;i�s;bO\��Cw�/h��V;���n�>��G!�/j[�9dY=���w{��n��2�����ҫ(�N�Ԝ&�E8��v;[���;J�vq�ӑ���C�now&�Ϥ�X�L6o��%�>��v�{�Q�5zdOD���2f�8f��;N�� q��<<4�b�Y2yv(Խ�%[y3t�vzCc�h��f��K��<�	�[Nh�L0v� m�n�6:g0�֫�h�nj��s��y�)�(�v{k�]���ķO��MŜ�nL��������G�t�׊�|��6�V��{��W�}�� ��&r���3*�`�흹Og�',�N5rK3�������� O6=e|c����(sU���wٱ���j9n� ���xߥ(�>���O��j�VN��=����Y�b�6��J7��x}��麺|������f7Y �`��叉���ˋ:Lb��^�K�7����y��K��W�9��/�M	�+�R�f_q���b[�}qҳ��W^�&I�1�9�#NA�J�|��z���l���vX�ٶ׋��I[o�eᅟ�c��=�L�F*O*�#�u�z]�}<�R�B��j���m�2|F��Lv똷�T0�X��T����3�����Dϧ��9Y]����:ܙԟ
�Eyiw����'.�jr�{'v;'��[m��t�:j�ɕ�͜�"߯E��M+�����uU�����g��=�W�\�OQ��gܩ1�!�;U�o׷V����t��i�{f������Rfˇ$�j�n��u=i��is�������4��ɂ�i{-�V<�@eO�p��.�-�x���f�bh��ͧ�KVY{HMW�f/�������w(�rI������m�e��`~��n�8�ŕ'i{+F�$�O2��U >���C��5=����쑷ySf�f����ҩ�WJz3��g/f������.c�ތ?����s���񺦩��S}ỷ�Ij1"칲n`�����l����;�xwo'����Ke�t��7�Z��O#\��z��]��ؾ�W�b�|������}�6OG�I�䯏�/�.��u�_O��Ԩ>�lN�:�{�c/�d)��*���Տ�^�~N<��w#K� ����Z	~�8G�����D�ߴ��K�$}y�3��uɈ�a��$�uS��ޱ��/�PJVR�6�;������ī���3�	�0G6��;�}Ɏ��¶z(�J?vl�f�9M)�}nu��)`0z���Q	ި�!d:�\�{��;J���!�z���맏2�o���G^@��Ys����{:������1�Rt�����ω�룖lJ~��ie��$6����'Q)t'D�D�iMe����bՕ���h.��\
;�&�h��0vN�]Jʓ�}T ���gv�_�*N�[��mo��diQM����#[�?*��|LK��+�Z"H�~1u^�y��ʲ&��d��0�{oOR�.�x��JN9hv�e�'����K���5w��KCI�]Ұ=�=��y�ֽ��8-׼"��͐&�������,����a*��8�������71Od�@sy�X�23�w���wb�A�<2૩��1���h=7vz�gҳ�/�땠f��C8�������7��e(j�'.�w��!~�k�'�ԅ��\���=�٦8~6N[tj�kí_t�i{��&�C]��,�/��O�Ko�Ĥ+�A{}�a�V��f�{�c;�r�A�b!�L�[2�m�6��{ط��n���o4�;/s�R���t7=����3�7N���@�s86�XL����w���ǸuJZz!g(�X2ǄG�bux�{�q��VXS�-ث�wa�Y\ݖ�(ގ��'͕w�6�Ǜ�,	����Ȯ��V�4�J+S�������{�\r�����R���Rۖ��n
�:^G��Y����
��pI������Z3�&.^���������S�:݁���fJ�����?䄖�9���V��I�6_���F���Gs޾��[N�U�pʎ���d��W5 ���;}�WnB���H��]E���)�܎�{Uo���%��R�l>�!�Ή���6��oμ���15�ޚttޥNO��n�Ϋ��:<x+���; �}p���57Ν�Ϙ��+_t��T��1�_����U����ެ'y`� a��-�zu�t��>����L���F:K���Tߘ���gQ�#_�M���̙���u��������f̜�K�a��Gc�j�'�=�ԛ~�yr�>Y�Ľ�cla��{��~�.�➼z#�S�C��)=@��y����h��9�<�__vߔ-r�o7K�ED��҉E��<�ë�-T���STy���Π�����M��4�|��F�ʵ�COJ�*�W�V�.��2����jz��i3�����;�mc�lM�t.� ���v��X�+�v+۶�5d�#u� (�f�B����6	[Ygr�W�o�zD��(��|�����v?������2"f�w��9��'0k(�z�/���3��{�]�y�����ޠe�}9ܴ����2?F��N�dB��-��?酏Jk���m�h'�"��87�`���ɒ>�l�c�鼒�𒆇S0U�e���5������ވ���r����͇��s���%���׬�}Pk���N�͜���&���<��Ϧ��oc'����{���Z���7=��'��k(?p�w���vlL���]
�S�+T�[�mq�챂H.�>wU+A��pT�������nm�t����]�o&�ʶ�+w�t��N�,)+�per+PS.�==�A?T�0��vߒ���N��۹6���ި�T�!S�ӱmu.cD��#w����W�����{�����ꮝR	ޥ�.8�}�fof��=�Ŗ�������:�=�v���� �-@��i��t6�8R��k�0��M�U*M �;�*!f��Dv�����^WFq��I*��Y]I�Csx���
�Iˁ�1�0P0�'�]�9�3a|�����%��}�׆j��ӃC�����^��#���ʝ����+Ɗ�HJ#*V���`��}_W�}� x���N�)��v;��(�k��n���$`��F:WZ���s�n�+�'k{�ut����-Ħ���j�=�A�10lf���ș��I�э^���RU>Uk�K��zQ2!�ŭr�ʫ�l�D˻ͅ$�8��}�U��/�{�+ݖ���e���~����A���.�V�R)w�ͼ�sҖE�ϐ�k�wwbc�xb��<3s}<yQPB�o���ϧ��w�r�� O�
�A���m���qWj�t��	�rCZ}�"�v��څ��:�R^l[�3�_���MLrY}���242�X�t��p~�i�� o�w��߫�lL���SD�N�؝yD8F�~q�����09���V�4�����/����:�^:+�����r�a���!�mq��{�<`��ш0���b�R�9}3պ|�7F���.��ѱ��5���w�#X�^�GA���jM|$W5��c]g(�/�8�uw��>g��.�{E��F^�Ĺ�:��㺔m�'�lUo�C�%��{�Cb�����.�%�&V�~�x��$+$y�[6���<c�����N�t�Н����:���~1��{b��O�gO�C����} �]h�}w"F'$��;q*��Yqc�r�|�ze�S�j���v�҂��wt��ߴ��ޮ�h=x�F���C�������m_���v��ݢ0�i<��4��NŵԽ�s��6�5�ew�0G1�[�Gm!%{
�[$����G���!��M�~��dYY���o�tTVT�Ϻ"�l�y�	�8�G�h�Xg��y��ZZ� �ڶ�=5�:{z�ʚ�ǱG����{Fl͉�%����-k���~�B|����4yz���1l��\�پr��{xv��g�m�5�S[�����/�Su�:=���z�ɥz1}{s��O$�'�|�{�c{�D�ec�wLh�fF�&�{���F��0�x�'���z�L�hi���tGN����Zs��],u��mM�m]r�[g{1{�yo�������2�\vXt�dQ狻�}�]ŽFʲ�֜������Gm��U����U�o���s�� > �?�۝�M?�v=��y�^�Z��ÎW�umzlߋ�f�{����=\R�ޛ��f2���7,v�C]�l _!pvJ���@�x{:��q��J�t{%�ٜ��d�C�M���S<,�� ��>���<�Y���{y�����*>2f�h�]��������Z������7K�����b��O�~����v^��=�&�ǩ0$�g�����n�x.|Gfx�����T�� =�T�na��?I��_s�v��ѐ�y՘��,Jl� �ͬ��Fj��KG����^���Q�]�6n���e{�B�p2,huWx)����mF8�ͫ�K�՛i-oc��2���nx�nh%���6<t?�zL׏��ǖVۑ���|�E���H�/��(�G��U���&�JA�Bg��|��i��K�3t��|YpD�V��8�
%�����hF��e�(�W�m��Ą(�si���ۜ\ux2G�n�}�>q�vq&!F��Y�6��ѻ�(IS(�:��|�y�f��o�J�J��X;�:L�	��P��n��s���6������E_d6h췱|𫦮3�Enb��&��{1&�;AI]!ʣ�sy�bMs�۽�`ao���v�R��[{
sf˿�Uu����O㲅9��h���u�	�/����"�}����X^�c��;��o�N�n�إ&��mM��y k$�g�����eӭ���f��2�\�NGl�����me�F�'h �3N���;HLD�K�A�;@�#\��p��[���S^�[��ƙ��&h
њcYr�����N�N"RT��U�,�����_\ͩ����X��Y�qE����Vr1=�q
�w-�`�WD�Z��1뽺�L8p��Ǳ������κ�����{���}�ȍl��
����:b��y��͑�7V�s���&�jWP�[s%,��I���CK�7�G_S�x��+��0Ep���[���eY�}�C4��u�hL��y���(�6�&V�tu�����z�JP@oRv\�N����C6��I�V��@�*��ޮWuWe�}�ŉ���bov�wQ�]��[P���v�%Jk"+w,�p�2��0� !p��pֆ��ƻ�ԟE5+dR��M%�a��%��y�EAjMѲ	C�듾}ǰ� �7G\������άj�6��ߒ�j9
��n�]$�G�������:���c��y����)�g�K���!>���!�Z��P�I�Lp�����O�x&Tal;L�S��mL����ŗ'{0��c�ŵ
�մMaV�ށ�pۂݍë4�F�0��q�@�&5�C`�N���24��=�*��n՝���"���[u�9n��{�OLc(s�4q��K� �5r���Q�q�9"F�]׎���0���yY��������^���.�غ��b�qe�f�0\�H�g��QF��'6��;EŒ����㫾,�8C��+ucS�ߘ�U�F��.cb��r��r,�R�����P�ϫ4����R�����i��w����@�!*�n�����-�t�{2��9m�nݍ���K��c�X�j�¤a�Vf��eF,Q�b�E���5>&�\Z�ػ!l�{�Mܧ��^ٞS辱\W�Ȼv���B��я:,[�����$�_v��t�/j֡֬'0]�QJT2�־�c���.� U	M3[�3��a��f��$�=�*
��wr�1�S�n,���ZT s6�ii5*�݃B�u�ٹ���TÇ�o�o�1 �]�{�xo�,1Ǻ��nӴ(��բ,R�j5ET)cV�j���`�c(�j����Vլ���[C֤�
4QKZ�Q���V��Y����J�[
,m��66���J%F)mJ[Qm�P[J�hŢ-�YZ�-i[m-�TXє�(�l����[Dm���KD�-�5R�X����[]\r�j�j�4�m��D��5,m�����*6[��dTQTb�-X�R�J���
6���VVU)h�U(����.Z�-�ʩF��jѴhRҵ(Ƶ+MZ�-5��`�&%EX�X-F#\�b���Kh�)2�AU����b,-��1�]S1�U��D����QT`�X+u�&%�D�R�՘ʱ���J�kam�������J�aJ�m*�ŔE(�h����klU�"��TZ�,��R�[�N�KR���#+E�Q��T�U5(�mV��CMrڭm���U�@�&)
a�����V/��ˣ�fv��_]n�I�˺h�N�h��J �,0\����Z��U�V�R�8.T|�s:-k8��y�*�����]_����奫g�����R���z3�n�p<v�=CKY����f�ތ�wq[>I�j�=�A�M�ٓ�Q��C�������J�w7y��[�w��Q��ã̯umbK�k���m�|� `��-��Μ�{ۛ��?.�e�XK3�'��{�������T����'v�g����>���5t�:��o"˼cp��"St��}����ۈ��zD������g��cۂ�8X:��`�wa=����]^`��v��ԓ���3�UTm�QS���<o�T��9�ws9�^��m!��Z�:�&k�N�2�#�T/_g���̓]b�A=��K��_#ps�5�yT~\��]�}�!�t����P��N�VP�0�K\��6;��i}zG��&�ɓ��۴Aro��]�z�Q��	�z�T�At+%#��۴H|V;r�[�1b�`��%}}b �&>㽜���W$�Gd��X�=�ׄ�mjxZo�'��ʺ���1L��"��5�۔�������y�W�oC��hL/w^�tੌ�!�=�y��vC�(rl� �r>�Ͼ������.���:���V��o�R+�*���	c�����O��zҼK��q��vh���.�B�tL�28))w� � ���i��O%�|����(<T��lڸ���rb������HCE�T�?$�����͞�'ޛ������GR��8a$�Zk5��w�_Q�7�A�b�z����8�!�U��RN����jo��]̛�?H�5 .���x�v�ĂOJ15���10X�'T5}J�������qdy�yN%s���EW��KC!,��B7���/<�ºgOȉ�ݗ�S�=���=���,_�l�]-ǿfᒔ�v\^+s��{M/_�z���rJ�'wO`����m_AhO���V=O�̆�ە�1�^�D=��0'+>��t����W�?]�q���P�dЖx��V(�!CԚ�{xh�)��:���B
����lS��'��x��u�[Wvs��W�� t����E䙵;��k��3VT���jvCٹ}��:�+���|>|�`צzv��~�����'/6�d�噒eq�5��=v�s����������]{D*��S���ʽ1�z�7�^�pE�Z�|<��noe�������;�_B0/�_����FS���Pf�2�/3��c�~���O���&�RM3+��O�ӭ�2ַ!b���_�Մ�O�	'Ջ��]<���R5�͙%`>x�U�{�Ю�i�/PE����o>����kOg��ȅ.;�=���29[�L�b���5�rè/�h���Kd'�z�������=A9X���VW�˦È��ʗ�=Õ�L6�`c��c�w*su4dG��s���o� �'���f�|zn���7A�Z\����ŻF$�k��ٻ��Һ�ŏM�~��dY\���~��Dg,���S?�q��^;U{����wPw7L��6�Ֆ���6o�z-\_���}c@.���>-:p�;�n�.��K�R����nRn�m��|��� �[�ޡ�sP�JVh=�.}�q�V.bښwsl���ܥ>�_Ν%>�|6�S�*5u5����6�u���[�ه���u�I�%�;�k�x�ve,3�}�ײ��0cFc�2[I�v��/�t{K���gG��}��u'������s�W:�d�sð_�=W����+���_t�7�of�?�뀙=7�Ӛ1+��=�˅�.b��l��h���ތ{q倸,g^Ю�d"Z��y��=&ل,�b"�Y�|;�n��ϊX�Y�"��<U�h�VoͿ����uv��~D���ut��<�6�o�ϱ��]qI��d���o��
|������!���<�3�N�Y�i���w��:���,;h]O��.kk��w/6�������N����/9Z}ȼ�g�N��R)�����}p@�
��<�^xo<[�H��:5<����j�>��t�g&�3K�37Md	�\�:���}��
���{��u^�%fh4bs|�̖V��s�������8�rw�O�Bl�݀�^�<q��E�A�xS���wYe����wf*E���J:�{��ʹ�A�C��5^S:�*Ǉz,��}�����*�?-nn���f�y��0�|9M��tv���^:�����Ѷ)L]XW{w;g��z|9w2-h w/E�K�R�T��*��k#ݙ�M��!%f9����|"�J9���d���6<��d�]������Л������(��*�	�S�z�Mͬ���"�����(P�%M�?<�Z�/O��P����+(��.�ns[ �~�B��.E�Tv|l(Ő�Ň�u�N���n���}�.�E驗u�(*U�䖇nb��jT�`	�g���D���B��m�0 ���=}���ܥ����g����T�������E��W2�X����9���ˇ���5o��H�nTha����8��`�ڻ�d0��P���z�h|uZ6��h��q�����|�Z�x
�+4uש1��OO��/���`ڏ�#-Y���,�̑��B������k��-�:޼��:�m�L�4.uoN_Z���G�#V.{�>�q�|iT3tv�SEȄ��+�|�hV���}l��jɏf����8۠v�4�%u��;��AI�v����ԫK[VĘ#��u�>U�1�t��`�Zx*U�M��h�`֩N�*8��z�.����V^�ڀ�������|C��L�lk�'%@�ܬ~o����T��O*go^]:�AR�x͢��Q�CPE�����j_
�R�]p�9�V���-H6��󏻇:��6�,ίQP�%|���Vi�l-����U�4���� ��4�� �A����V���%a�+��W� �,,'w����g�A;j��}T�E����\��7ޓ"�������X���G�C��9D�+:��*-��Z�:���A]�>�=�iI�V���mN�+��HU`B�@o�D(U�>�Q<&`����>V�M��
E#�Ζ냯}i ��FR��i934y8�]aP�a��&��B�H�<'7��lƽ/�)��u��ה��-�D�D��Ђf!Q���Y�k�%շ�5�]3q��;p�	J48M��`^�y]�䬫ڗ^�!X:�G܀��*�*/v�M��K��+h�=�w��r���ҽ#����]�4T`t:K���n%��vJ�@
�X��!$��u;vG<}�u�5l��#O��}�x��'o<�[R<�Sw��8=@�B�t��[��v�k�`��rS��@L�g p�9�yqo�d{�Q��m'`1Yp%��y�w[�Ka���*��3�n/'t[�#�l+k���P����T[g����ᱟGlq8� W��Wu�u������ur���;Q��]�7щ��ޛ�"9�eK�"�bxleM�}�:4`��G~�A�«k<c��wi���o��'s+';�U�T��R���,�U������\|�rw��˩��NZ��~��`���c�����W�d�Ax�{ס�Z2��]��g��W�xb2ǟ7���D�<'����f���/��H�0O�b��u-
��%��pBUM��2D�˛�A3{ӽ:���k��xT��危��:B�Y�
β����%�������z{���bIwT$��s0�����+~���-�����ѥG����V��R�v\>�S�9c����&�Mv�xWy��&���TEL��H���L��(@�:) K��NV�Vc��d��#�$�tu��0��v���E�X�_F�,�Z����F�߫g�ª�x��'���w�{]o"�;�(_�.���<&Y�;�%�t,�H�p������7�
TPf�2>�FIj������<a�	[.U�Y��&h�G��tHr�Ei�Q� �|�a}��޹�Ċ�_`��w���\'LUگj�Q�:s%G��fṿ��qo��V����x�s�uc׎ì��e{���� ۞ݭ	��!ae~�Y((���_-�z��ಗ���"*���)��Q�&lc>��w�kg����Q��*����:��)E�?�:�`aA������A��'l$���Ɩc�$���U�\ηV
7w�wg��EcU{��K���1_<B�>�{�z�VR��nЋ�u�U-Ё|g/���"�xH���z({�����6��{m�Z�;�������^���
�����Q�����A�~���.p�l��<����g�d�vso�~���E+j���u��{��Һ�x#2��t�Xg��l�:j�ON�u���v���`�I����7��2�h�/�y��h|�׆o_�g>	X�|=Vj?�)�Z8)������FB�m�S�|���ϱۨ]�<3�K��z��9��`ޗ�1Q��z�����G��YuO����r�o�#�q�G���<�Aj�å\Z>��xߤ�Պ e4!�Rx����0��kL�oylPÒ�x�+�+�*�u��c�.�O�v��kSԭ�'UZz8<�s�+��h���A=51�>���<E��GT�3x=�0Ӝ�д�p�%k����nU[~�]�4���2���kl�ܳ�w���u�]$���z�?�U_}�չ���׻�p���*M�b���T���q�q0_��,(��Vժы���ml��;n�+EոvQ����"i��٫��=@��cI��R�^�x��gV�1`�h�9* ���C�5���v�iH�F�t3ݶ����7�DϽ>��*�]z8]����b��*N�$��F�3�n��Y�c�yjn{�5�Ƕ�P߼+�R|jy��j���n�eC�u�5V���v2�{ynR���M���g]kKY��7X+�r�B�X�9Cnd�#���ᮦ?x�:�~��W.�����m�\w�j2�khS��j�ii
����1*�]�jw������n΂��+��_f����2:��#Z0H��T�]��^��hz_��,��|㱷BP�k;:��&���nq��`�󽡒0E�<������UwN���Į���~�k�IFT��А[f�*��K_v��mJ�}�D#�4�<��c�	���.�%]l��^�C-Ԭ@�B�̡>;&xL�3\�N���Jnb���?9��e��i�J��'X�j�R�Z����!���:w>]�	�o_L �N���wb�T@9�\�i��u�'^=����Ҡ��:�	�����]�;=l ���|>�"Of>������y��W�+%u�Fx�l:��C��u/5�,���f�i�)�If��G�J�h���V��T��J�1
�b~2��\>���Ы'�<��yދj�+[y�yS��u/L[Q|`�tNw���~���-�!�FU��v�Z�Xf�dG����B��]�b��� ʨ�Op߃�/�����7�[�ܘ��Zz��5�-��nv���<8J�uut��Z���v�ܟ+�K��n��P� {흨�;�z��Sٞ��w�Ѫ\<2��dI�Kˉf�1�hj>�Dui��������k�8Wc�2���,��k�E��b��m�Y�tBd�@d��i�J���=�E��a�Իo�J\�3��Pw��}LWq�{�P���6��P O����ei������}*OS]
J]���ݮ��5+�;+^�X.���p���p�d�B�u(��"�����{��7l���~�J��{���]s�kƜ�h���u�(��'~�ϝ�r�b��Z��2>�Л�hx���Zn�˫�ԛZ&^f!!�T�7`���m�em*r�w5���5��wJǸK�9.E>�w�VҾ�W%�3"Uƀ��6��k�}��z�P���D5S�"��V0�U�ڻ��ݎ��xi�q�K	6�avN��M�w�-iq��rF�$�V�uy��}y�A�b�c�Q���[�t�0��D���>�ܜ�0>�p�Z0͠��qZh%&^�]n��E�7����M4g��T[���+��D<�w&��\���))�/R��J�=u�%
���`���;	���ڱ�
���H�ĵb����X���gW5�u���s��nlv���Ecؑ�^���nk��&Mo��mE|��-�Fm�5X�(�����u�ޙ��9��َv�s��"�'�w�U�5.PKDwsl�ƒ}x�m׺��YM�)|-��-��{�6�0��{��.4�K�e����aV]q�Ć��$��<շV�_��i꺙����GHֈ���+c�\���Ij�[3��d0�w͞�<lwU�����
��>�UtB�ǚ*� ����Yj��P�uۘ��o0Yy]L����*ȏ 2ʏ�D�B�����^rDV��MвTX)X��z?c��3���i-LH��c�^�qW{����ຩ�?��+%�WW�Z�O7���{��h3��OaAT}v0]�K���5ٚ �C]{�n��ee�B7jm�y����0�^C,j�ϔ\mfk�F8a�2Ҽ�:�����_ش�t`�۫���7���SAgjw2�;�]�#6I���az,g�f�HD���*PEkf�Y��W��r�m�iB�Et�]��k�5kI���1S�R_x�f�_P筎��[m����}b��ٺTKx1wV{xu���݂�X���[z�hA�����>�|�	���↊���xL�,.Bn��Cr�r`��[v8_^vt�����^�+!bq��_&�7ǲG!x$-!+Y$3Kd�K4I��ʐ�q^�0yWR_]܏\��{=���,,�շUn��q���f���4���Sz4�������A=Վ��[έ��JPG)�F�Z6�ɢVn�
:�U��4���_K�h�sdn�2�M毁���;�l��s�;����� �2�$i�r�ٽ�)Ff܅��V��Z�aC�]��_uM 8�y�b�Gy{�N��|�8����׼�Wt��]�v���I�f�Q�Ԁ����q��`�";O�L��ki;�	��qx���nY����"ht�-Vz��i'�Z�!{O84��˵����O#=]ve���I�ZJ�u�w��o:��Td���� ��ǡ���!y+S�{mR(��e�϶%@Þ�Y
:=^s!"�de벻8���@f`
n;\�j���k�4�s���hCv���MY��Y�g<v�d�� �ޘ���{&q˷ϵ��~���4-b�����YYU�ab�T���m�Z�q2�(6֖T��Z&8�e
ԩZ*��jP�ܕĵ��������h��X�ٍ,(ֵ��J�QTcm���Ҩ�ֈ5�A���X���b��J���)J���j���,Z� ���-�E��bV&Yj,�*Tm�˖[JE�T��UUb�*�db(*�R���V�-�Im*���Z�ڍ�ZEjY�����1�Em�-��ŅK�,T�TAEX*��J*�KkRZ5�Z
�2�(�U�Ub�Ym���KF*H�Z#im++YR�*���*1`����)k@�QkR�E
��U1�5�%�*�,Z�E��A��2ت���(�TU�V�Ȋ��((6�E-�,+�b����EEV)m�J	i(�JUР�����AQUUKIJ��`�Q�RUX���mQkQQ��\���m�"�J�c��0YU�P �Q�}G9pL���(RAZ'6��S��q���+�Fe����ɽi�H+��Q����^gݣ��R(W�Ʌq������	w��/m��1U�je���m��V�7���&}�G�.K�
���4B{y����(����������/'A*Γcaz��� ���r:ʘ%רPT M�>����7����l3h�`��|J�ul*tV��w��l1G�Ve$>��s�$6�Uћ��\s��C���?�_���4P���֗�E�3a���eUx�0y�WnqA)~�h��os�O� ��ᱟC�I_Gu���ȃm���ߢ�G`�����J�����t�*��H.ʛ��G��H��mک��k�7�yh�b��eOh?����{�%U�'rvQ]O=����8���t�  �� ���^���/�Ku�;ض��.���Y�Q/>�B�r��$��l^%��KC�^�c��m`�v��)�L����o+oh?jNyg:�=�g�0~L���9^��k!�e����ϰ*k�!uU�n�vt�%���x���,��V֣��M)clf������*����_e��V��<u�+,v�^P-'�(���e�ƣ����Q�ŋ�kD���8b��S��}�+H ��*��Xdr^��R�����1=�ʛ�"�Ʌ��t��&���I��F'�:���0�z�2���;s���G�tr�09{�r"�n�ܑ���;�Y��}UU���@/�l��>�M�~��]r��6`�>�|
��3G(T�:�Pt+�~N�D��`���e�A�V��M���(������I=T�`��P�J=B�'�
^��)�좦ͬ���SDJ��xF-n��K��E�`�,�3o4L�u�>�Z��Д}��=o�_���ʽ�pV}��\�Cr�>H�jC������&��R��{�{��u��^K_t�T���e^���r�.�m{�~!e/q��r<��.�����`�̼�����\���xn��EX[�I�B_�T���f�p�4�����[�n���$���Y�Aô:P���3�k %�SB�L��]a��u���?.*_�5��7��B�1�^4����[K�BFr�9Q�a�Tw���V�X:RPX)3���*��z�����-N�Y�O�*9�/��2��e�Ȝp�������t<G�`�sKI20cO� �OVⷴ���CL2�^Ag�ٴ M������f���gF..6X�p���g"��֏�v`�aӉ파?{�,�k̏]ޅ�~�ճi����T�c��C��.i��hiQ���35#����~o��(?_�.����		�[Cd�hOC��Q��JȦ��3�Gn��+���iR[���;y�nw����� �0M�%J�߇@E�
l��b�K�6�N1G��2�ߎ	UX�Q	C��lð���4M�J�t����r��W�S5��_����4o�S�(*�)\J�\!��႖nzq��k�c7�o�z28��^�<Δ=ACO�m��2�Ь��Pp����y� O_�Y��ʵ=�!�Mo��yϱ1\^-�����I�_�U��H2�U��+�:)�Ym���6/>>>��mX� 5��@��c'���}s�T�}����H�,g�[�v�Ȩ.5�2��0�6�]�R$W�.�Q����l��6��`�)��w.��jW�v�.�
rx��=w5�1�u����4X���@���3Ht���ڲ��Q�ܘi��6�BqR��k���\&��+���T��t2C0.���������ƴJ�e��*����=[X�g�D�(!��~C���K��^>SQ�^=��X���(�|r�Z���A����:ąS��R.X��*qS�"8y*��Ex
��Ie�.������s-�{[����f�LΫ�NrÌv�gP���w�>�+�l������F�ھ�Vs���.-̒����
�w�jr����m�C���7:���bڎ8�
���,��`R�np��ύb�������s`�*�^�{�|  ZS3�[�guf&k�:���m�IsU�|�A�h1	�g9��6Y�)J��SvU���������hi>�+��O�v�|E���J�*�#Z2��e[��w���)�Α��$��]
�9}|,z�bc>�%�6�J=�]]b�h#�ޤZǍx��&wz�eW}�	4����`h>�O>���@�����m��h���Zє�y+=<�^�)����M����/���sDyus�^孵/M�	25|
��3�ws���c=IY��6l���u|��K���S����$�f�E�r:X,m�uEa��8��*jm�5�Ү��C��6��c~;�S�-h�`�tNw��n�ҽΗ��ã/�xx
�f�����6T7�Rc��YR��2�r��
���a������a�R��K7����l?=s8]%;�:IG�,�ʗz_d���`W/��8�"����<�%!\*��VT��`�M髅X�tT�N\�=YW|	t�c�hvN����x�/�D�*��*q���<�B�Sj�T�k�����x��3B��|=�\<����g@��@�TL=��>�3)m>�SM+ǯt�QG���JV��CX�{X�5�jK[�2�)�� ��a��y����l��,�0)�e]�V�$w�[�*������ﾤ3O���������n����w������ N��^+nW�LS3U���~KK�F]���#���-��w5���>�Hm���o'�"?m
,���s���u��;:F$��Ē�%/n��=��&�|$[�@��¤�.����A�: |�iYث�u�}M�����Y�LcZ�(f���2��qf��r9�8�]e(�" L�\��;)i��+��Ai3�B�S���u����,i1��\�C`�[�ҷ��XT��Z��Gw�D��^(�;�E*��Qb�|U����`p�p�W�:ʌy3�CG˚���W�]Bq��
���*��P:L�ӕH�9�<��:����v�k������u�� R��p���7&W�zzs�^���B��H'�[4����aY�=��W��t!+���h�1�x_�߰�㨾�~�'`9Nyh�32���������W�ׄ[�c*o-��ѣGd*�+m=<��?>���{rޠ�r�TF���׶�&Y[�8��<Ƭ�V�kr6�1ëd�U���۬>*���Q���6�$ɾ��Z�6��ש���g�T��d�\p5�a��X���r�D���-��dn�����,M�M&���ڷ(t��]�����Se.�����������c��Ŏ�~�Ж��e߳n�W�����1^�;�7����\9S��y���B�pI��Ƈ��7<�S~'��b�]�� >:�;bg�:z�<��s�q���m�U�T��O^��\!`���_U�G!�Ժ�U�����%��&�y���a�a<^=��_�w���}˻߄���~�s,�!A�F�Z~��d��.'��Y��ݲ��}P���C1p<�m��s��j[N��6�FPc���5��\po���%���o�E�ǹ;�v�r�S�����{=�E1��B�7�:2��E��@�cЏ��)�oz��*p��v�%X]���[�][�9�~Dz;�f��7ҡP�A��<ޭ��7��1:�&�G�\���ª��]�:r�z�M�D�WO�^��U	��w�=;7S�+�����t���Ų._�i���~�x״��싁͛μ��X��t�J��v�_��2������wMT����|��)K�j�5SM�|�S��V�9݇�GϺ�;�;�������j.�R,��Yd\Z���, V.b��@�r[�Λ��T�e�#[��ީ[��Un=�g�LDE���H��tN��`��	��X�_Z]������d���\�����F,�@h�U�X�j�ꡑ�Kc$��>5�?�W_
��%ϥ��
�< X�U��"/���_fz�	���4!��Y�m��M!G��a�oL �N�g/��𲢨*�w�b�W���'l��?(�t�ݐ����5컨4՞0?�X�7�w5T谟t�Ӱ�4�9��x;�0u'�H�_��\[3���,7r���շ���NC���:�i����� �n���@�zzӽ�YO�Q+<Tļ _{�h��(����@�ڕTݪ��cp�VKH9�˽I��d�|�*����ߨN<;��x��Rh�8)�
�W��z%[]A�.'Y��C9_���\�ɱ�5I�щ+cۻC$����{n�z�@D�W�~�J�#����Z1�y5C�1V=9탙��]�A��p��0d�ɌC/E`ލ�G��R����C�aj��僵]�Vt�z��;7w��C��Pʱ:�����==W���u}.�M�o<b��A֬��Ȏz󚾋 ����~/��u:���u���Z/��t��8��GM^��+���=R�
2��B�,^��<x��e�:\]�߇�+-}�-[/�h��i�%N���DC[�X�L@a9���^3t9}���l���?.�\��*)NL��¯��(z�p�T������T��#�� �6wv��+.��>nk�c�����||���}�g���TLg�G�Y���[c�cmX��n�J���e<\p�t)^{��$��|z�DuXĸ�ϐ��Ty`�a�� ���j��%���L/<]����4`�#�ZJ\��n��5���^@�qA>���!��^��װK�N2<hx^V���"ze��5�Vm�9�N."Y�2����!qJ(AP�ʥ���:��mݼRc���Y��L��wa�w����ES��,X��4�%ߨhp�YI�ݛ,ORy9}���67��[�� ,h��W��KP�wXF�=s(����z�`೓=�s_s���M���H!�:'�E
b�z�PXY����Z�z�5F@zeP�#Z������P�%�K��9>�{G�����i���V�xC�_���h��ѷ����*
�{��<��;@����r����[��$��xcD�iP��ƫ���5������W����XT%'��	ձ<75T2����X/~�1
��7L�1�X�7Zzi>���:t6�u���Be��^�ۤe=���Ə�)�i���X�`��EՇ{�n�̱\�d���ںLI�����s"�;�T�~�&h�Zu����t�}KI����Qy�8(����]jb��K���򇹝v-���wO����%+�[~���hS��IХV}�zXf��!��ю9�+۹�g�c��f��<�:���	���!�rr�:�<��W�,t����Wx��5��q1[� a�U6*�T�g����{�����^�aU��[R��Տr�a�(��s��]k�yƌ�1�%n&%���{��ɬ����x�B�9V�Q��\�Kϫn�pOE�3z�խ�jK��;�D���g��ҡ��tq�X,�'Y�^Z�_��K&'p8V���g����p���k{��th@:VM��yM4��*�	/2惠�ϕ4~�h��f��~/u�esܜ����q�;^��!���4lN�V�߂����ʕ{2�:���סT���F�^��ѧO��q��B������a�&a��9iy^�0�a�4�v��{{��<��H]W�Wp,��A�t�c,z�z\)SɕĻ8)�N��^$�XY�s�[�a�K�>'<n��&M�t�N�(��k!bW��/�Ř;��`�[�ZͿO-���@+�=h�1T����+E��#}֞D��ݓG|ˑ�'��9/�5��,Q�_���l���G�ڷ�g\]�>��]p� �9�X�����|�:
-�~���¦�E��G,�k��vx5@�x��h��>YԳ�:N(mea�B����;Ip��3���0�<(�Ռ�\?-�=h]�k�Id��*�������xQ����7]2�;�*�Y�W������Ľ7����;�]�����p�qk�'��6$<4���q�`��#�w�p�|y)��,0￝���?�\�����*�Rt1z�����4L�h�d�[���т2AG�}Ҵ86[���;c����_�������CL7�1G7:����6Z�[7�k�k���7�J���q�"O�qs����o��qK	�`C>�u-����L ]^^���.� ��4nӶ[��!q��m�i��װ��4=��hi�����u�˭�:��^m�	��L|�|�X��w��� �C�顓���o�YσfYU2��Ϛ�^S����d���L��%%�_y�N�Nīz�����-�>0l�x����)�o�&��m�B�"�
z������CUɤ�C�n�ڗ:�V�F���7���	��ɮ˫=
���Br�S��:� ��Z�7�\�A_]ge\UF�P�g��4M�����Hj�'4����F���O\��%�5^����u��ى����O ����u}���"lU0�&�BV���9࢜��Mʱ�Y���M;���tn[W�Um_hÊ��V
!��t�s�bqˇh��������x�v+ʴ��}Q��H[Zڳ��v��5��������� iry�rc`�^��V���2��*���%��퍪�ຑ��b׶��r�e�+����;���0��;��FV���V"Nus�ȫnZ�t%9[��v�:�-U��U���T�&�O���wp��-0*^,"tF���7�ۃE���i,'
Yv���ʲ��Y};d�EAΌ.��ƺ�\�X8�ɻX����ڥ�1�rvkꅝ\�i����(�;���fv�jڣ�1ҝ�GbB���c�2Jp�aR��xNϳ�l��Me�pa������o]e�[\��vG -��
��7��'u���֍[ҪwiC��]��. 鵲-��IM�-V��5)�tZ
���o���Z�[�c�����gv���l(l�9z��k���V|r�7��n��#������nN��[7F-b�m�7f���������&�N:�w4ي���s└к�Rei��F{ԎNw�b:H�އ�m�7�*s�xxӹp۷l���0�ŀ�Z�jMV�+�gu�gk_8yP宙W�mk�Sܵ.�o������B�����qnѫ�V���uk�#u�S�:L�NY��ۈ�4�噵z+^TS�v���:2�����{5��?�BY��y��u̻�*_SA)1����rk�׫[1�w"avQڶ�A�V�9����r�Te��,`��>G���,z`��l^��A������[Z��k?ru�uov�̤qz�f_����-J�|��a�����o��Q�*����aŚ��f� Y#y�v�]Q x=�ع��#t���d7�]���|��_��۹N��tJ�;1vvc�&)[��Qo\�"��Y�5(�'^j���z�U=)C]�ѿs�6����A�����kg)nF/��2��dR뢎)��`���Z%��cA���w;i�w�5�;X�^��Χ�R	�50j����_�P5��W�><k[�q�W��:���eR�
����a���u7�� �g_K�KD�ʃ$36����vq܅MǤ�3汦��l�-�*=u����r��uU�G�Yn�}c�.��ķ�qi�_U��,��h��:���ݤ|4�2 ���9)��}��+�1����1I�C��u�jb���������[�r�B�Gdy���>�b��ʌ��5{��3�N]'Y��'a�:�XETFo�+�(�L�D+�1�8�&��M��TU̬W��=�R�ɺ�ٱJcyV^�V9��c�]��k�Ś���k�&�%���*bs/8S\�X��ɓ���d����$���z%u�c�~u�Y6��!ν�LӒ'��l,��t���R1��5(��EUU��R�B�b[TcĈŅB�()AX����mPQD���*T�Z�j�`���b[`��Ȫ��EQH���ƊZ�E[J�B�A�(��*"��U
�F�����h��[Ub""��V���" ���"�R���E�m����(�b[J""��QDRұ�1**"(�ATb ��*��T�E`�+l���Qj��*��(��R*��U�(��T��D�"��m���-L�)m���Q���AAb
�*�Q�X�X�1"�J��F*�VUV�#ZT���`��U-X���U�ej��TH�eEDU�R�X�"
2ڊ)
F1m**[C�b&U��,X��DQcX�J#Db5��m��UEU��������#��TA�0X�jQEF*���Z�Eh�+
!ADX�R��m�Z�Z�)m�QF5�B����z��i©�վ�͸���x�8��VcǍ�,��$Nz�z�M�˓:<�F���޾9�Z�<������n/{gzey��Q��|M1�����\����t�עv1HB��_���D�h,T�5g��3`ee�wH�{�
����\�q�P4E��q�Q��!�:r����^�C�����6DZs���+o�l�u�(���>�ҏa�l�K�aUC���F��{w�MJy׋V9C�S�����SWQ��J��*���W�_ͺcx��m��6��u��$��7��4\v��R��xz���
��4-T��>��;i�bt�`�OVs��p�s�2}R���/G�MŮat �#�%����PS>��բҴ��L�~ۿ h��P[�>�S��v�%/{9[�,���4��ғ�}
�o��hZ��$��%ݓ��]]J�c����sAͮ;��Ra���ԣ�yp�^wX"�k*ǀ4�Kc������Y���/F�G�l�>��=�
Ͳ�'jQ݇�8��<v�UNn�r����V�d��G�eo�rz��k]�\0�}�����P�|(4P�햰uX+B5>Pi���N&J1c�*{F*4y���eht��E�Wh:y�Mj)��xv�heYƕ�v�s5��pהqS�d�W�:����͍V��{��<Vs�fNr�邳�U:!r˥ץ[1`
���"K��	����톻]�x� d���5x�˝z���+��R�A�N������MOǅ�|�)�(X�^��ӯ�7^�u�y�E��p���q�]�I��/;������TN�!�^��bze��Jj�$�ur�Zru��խ���'�e�*ꓫ� 5��*��c�����?T w��բ���;S�1�;3�FI`�F�z�����Z<�$+CG��}9v���B�P��!�����{���+ٳ�v�G��Uq*��tz��z!�l@���}e)_a��ö�m�x�.��z��;�+{YJ��X��]�o'�M|��.�2p��3���u�ۉ?k�^�e�$�9�fY��{:�m�.��(],��Cg�#�ڱ�l ��g4��eG8/? ����W�Lf�iΗ�8�x��2�й/��~2)V��t&��bl�xf���[��_c\��3��¯F����/�[j� U�w�z��54��%�A��eU)���%^�ĺ��ߦ���lo�L��!��'����{�Z�>}aM�.�"�Em����z�I5�KVR�e���KPW�eu7-)���U��KZ�s��֚ǳ/8U�M{J����\�X3!��B������[%�F�JH�u��v�`���T�eF�농�Cm��Rj]�Z�c��۠�ろ����hw��m��f�t�9N��:\:��3�oT�O�U�����9�^�@�fU�;��R�<��������U��WQB��G�.	{��c�z=Vge�e�t�%�þ��q��$����Z���YD�m#K�\��^���������-�4Ɔ0o���H�o2CG���Q���MeW��{���,ez+=���0|�tOe7	�^ε�x���7��W>/��+J�N����?���#�^���j��e�{�e-?KA�EۗA�F�˫ ��Nx3K+�%(RfPKژf��8��pOo;�v^}�OFS���� �=��O�͏qT7\�[:�e_�Ck<xP�����tt0�& Uo^1�a�]|߳Fp�(�q^�+[ݕ�1�*��ӂ�1jb�%����-�
ܫ]���G��}�4��)���Z�է0��������>��Ò��=BP�5���(����ha|r�B�j����r�'==��Ͱja�3+��X�Bo�	C����Ô�9���GҴ��Ql/۳�˹�3G��r+т���[���XuSy?�!Vg����T��hQ�����ٽ6���kޮݽ�|����tv��K�VS�<��4xR��	�h��y�J��F�u�����JK��?ˆ90�����c
�FJ�������b`����Ĵ̊��vqRVqP����������8�plj�捻�Zh��X��>�h�Һ���U!ǫ���1CA^���yB���c	+n^&�����@ѫ�"�vnHP�+���:Bf���y^��U�4����{����6��r��������V"�(2���z�9�*d���#��Y:r	vZQb��9��%lh麆%���:8�'�Y�5��+�u�܀P�{\=[Ա��I-��)m�\|�T���$+��W��(2��	�u(�WO3�sgҩ$&������t��eT�huewLgƝ	P��
_N�
�+躛�;o���\ɾ�-o�w��o=�Y+��n��ϾgB��-�ᱟC�IU��k�ȃt߰�����k��;y"���o�N�������Px���|x?��o_x�߳W��ǂ��4*��ּ�M�$�1i�GL���s/�93+�J:��u9Z��hKf��@�vf�w1��fB�x�����t��+Nǎϕ7��U:��<�A����J��bƭea��1@v:�]�)�w�:Wgb��{Y�q�cB��o9���hR���뢶�wIzeZ��_nq�I]�M�����t����W���~�ғ3N;Uy�׋��BU�-�eS��v�V�m9���+�iv?�>���Pz�����j���^>XR�ܐ�h����1�8���c��,o���qg�h���Q�'��9{�,}Q�tsV�DϺ]`�/��{�OC|:���1G� ������_�����m� ����RBw��6_�ʜ.6؆rz`u-�fz��d�v��F�|�W���KZi��߃�P��U��ZL������b���<��R�.t�`泗��Wr�T�����bT��e� �z�0�ge?+�냡�94�/{h��З7>�Z�z�c�K7�J�B�_��x������� 6��ۉ���6ѣY����o�j�"s$e2+��#�dI�J0_�Ar�P�;W�D��'Ǫ���,����Y�֋�����k�}Ghe'pQ���SB�<���XK��p�n��T^�z��k�����Jj�9�ō�JP��11�< ��[�J�A*��Yy]z ~��2��$����nad:�¡^����e��YsÜWVf*U��d��'H�A  T�)��7�xn�ߧ��N��m�DwA���q���րs� ��.+:W{��R���b{��yd�7]��ʜ��se���h�u$�'dZxC���5#(?��K{�`/�3ͱ��Rx�0vZ���]7c/�ho0'ֳ����:��}����$�>z�ovV��9��U�{L�*,.�D�=�>�c�x:[%"�q�;Oy��#��򆝴�&��y�#t5*��E��4�u��3��7wmv�e.܂��P����	�k���\v+IQe%����myK�ޚL�-�^Ј��m:!P�e�nǅ��C��f��2�%���a���r� =ݼ��+ݓ٧��g���
ٰ��4P��ڮ.�{[
��[�qg6鼡;��')o(!�)�����cW�OCՊ v��(�;0J@d�	5�<��K�z�6���𠎨+)�t�B��O_�o��%v��evkЧ�)Z�\٩�MhpН��·ۡ������:*�J�����/4�T�[�����N��O}k-���}�\� ̯	aAVym1���x�Fm! 	�^�7��gq�{��s=����Z�a�uܠy�J�r�0R ŕ��l@���YC��}�q̾zSz�s�;��\��z:��(΍j��!�){2Y��!.���*�]^�E��0n�.@�(��e�7�nex�2�w�}�����S�ׄ�:��745����k�e�|Ԓ"I������U���7��@����)���%�+��ں(�ZȞ��ȏu\M��$����w3n�#;{
<i.lQO{R����j�%��\εo��]�g�+f<�@��J�$�/w�eַ�}~���t�ޡ��f�~�F^�q�'B���+��u��:!6��v��^�VI)�1C{�μ�����`��* !+mTvk� d=Xeՙ�(J����r-^>gs�]�g�b��+��×��ez��9�
��\s��N(z��������2��L�kywGn���,���%�림U�.p�+�a�F� I�����Zڗ7�w���s$�`�*���~
�b��kp���aj�=�ᑴ�|����~:�%3� ��n�*3�z��q�B����h��IT����<��S(O&-�\����/y��f��k���К��|�����n����w�h�h>C��\�-�wg��+~��t}Bą{m	C*��1	c�'����$վ)�{�b��",���w���5�i��+ʫ�)C(*^���%��z�S���J�=�AB�ðN�v��WI�)`ѕn׌���씫���W/�n�t0�R��V���z�g�B&(w]^c/�]:���������)�cP��T*���9�Dn9;|�.Ӿ�M�찯�ރh<�7�w\������������ >��tDW��%;��u�V�U���U�oU��wo,�����/Mn��8ῖ��-�� ���{�P�<��`n#\�E��#s����?w�~�ͥs���~�fH0�{=A�0�G�duۼ�4fz��%�3��R�����_+����!L!4g�ND]3�p?3s���d���T���5k&u�d������ze�S�,x땻<u�����J3���W]��>��r�{�V�c'�K����Oެ�>�O}P䭽ȣ�}o��w�K�<�XL�7��r��ej�RX�R�n�{�Z���g�l�,: T�=����^!�˔�۹~���:30�4��xg(����Y�q���R�^�Q2� 0�@�Е���W�4g��r�L�L��9���uK	\��w'hg�l��8g��&�!UD��Za:���r'ޣ���X��Ԗ-��襳gp����w`�n�ET%�PU��
��VJ��]���	�l1G�Y��>C�}��b;�����J�k�ᆘĆ�Е *0U��Gd��B�����</ӺD�����܅-��y]ٌ��H�t����C��鯩�/f��#X�@pT�Ѻ;�]X��4������Jyj��pɸW)�¶�/F�۬��Ŷ�����u�
�x����N�w��k�zRY;�*򍐦�G}ݯ�N��ﺺ�o����y+�Cu�}ޞ�u��R�g(+.8X���Uv�z���d�pU�"+�v{���fW���[�z��iW}�g�;O�|�˺���jN���2��u����ɼ��ȷ> $Zg����/Ի�5K��{s�΢@P��܃f�R��r�h9m��:M�Iϯ2{d��xJ���v��k���i�x�s��M'��Lg���W�� ����^�L��N(ڛ�"|���Jk'������Nh{-�G�ώ�1�uOS������5�c�KD]Xv�r�\w�7���[\���¶�}���P�lA�">r�չL3�
�*��I�5a�J:-u�x!�5ڞ���};DO'��Le���A����Ƚ3��^���w-����O��e)���-Wg��}��N�T��b�M��\\-�˂�z���m�@�ȍ�)ء��m]�Q<�x�aT�T��۝G��y�y�5ȣ��=�x��q���ڧ�Y�վ*?�P�g��G���z��XXꡬ�z5�5g�p���K�����%����G���k��j��y٠�=�R�������(xE{vxo��y�dj��,U���^nt��kiǹ��"E�k�s�7)H�Q7Eem4 ��F�ƀ+\ӼZҶ-,�>�z��Q�����cg|����(��_s�e�w�m���2�ϙ��/�T�U'ˇ�i7K��>~Z%
�n�Z̙��촗7�R=�"�5��53D����..�EXQuB=	�^�����F1�N��`�$��ګ$dJ:F��W���\
���3C>�,� p�<�U你��ˌ��׻$u�l����(q_�䰯�e�������XgK�=R�ЀN�'ы�p�<S�g4+���o����:L���U�{�YCY��*���]\�V�H����@��\۹6�ެgIz���@Պ���O1i�ӹYL˪�+�}5e�Ux�����LkM�����m]p�\�V�kIcFh$d}J����@��Gv�4�.$}bʋ�k��+̛���*������eo������[Z�>5�>ЭYAC�Ph��WgK$$"M�'�D=�:y�)T��)0BR�(!���'#�;�GC��m�E�|.
;c؂Hx_�W�Nס�״�Z�2��[t��8g�풆���1��C�6��m3z'��f��]��2�j{;�0��j�m<y�K�G@�e���Υt�5�$6���C����Y�:���!yCFQxk�s��T�t�Uȣ��a�����빊�Q��]��r��ݶ�c2�[��\v�T���]��R�U����6��d����Z�N���a�x���t�Gn��l�4
��vF=�Ec�9��Ĉ�U����{ae�����6�+�s�3A�&�� !-�\dI�v\��0x��XPF��Χ��͔��j�����}�F�&�}4s���%�n�a�|���B�.+��z�8n[��D��2������
��8���k���S�v�֎c�4���f������1��[�C^�[����V�`2+N��fXy��B���oq@��e�6�/~=nu�͔v w�������|�� MQ����vv���M�^l�I�H��ø��ͬ��Ic
m�1�]�i���������y��6e4.
&���nV�g9��a�V�������
�oC����$B�Y4�r�o�+�G�ӝW�.\l<��`���b��6��8ܬͅV�V�$!)�\�՗���ɡH�i�b��P�qBc�%eZʺ��c���:l��PV@Mm���;�K��[������(a}����{�}y�$z��s �A�;�7ŀ�W/{�i�6�
�	�z�c�r1 ��W
��N��X�� x����ίjM2�qc��F�GFJB�d��īUҎ��^����W�9Vn����6C΀�X���+�,Yo+nU�0�s]+6qLl��%O��_^}-^��)T���U�[ƻT%���R|�8���X�i
Q�����slSb���;�ϩ�Ɩ	xn�{��\��B��H�|�-oE˞rn��ҽ=o<+=�Drm�2�����z��y��r�3w}�RIK/[b.���b����,J�=��+[�#��]E���h}��Z� h�
!|�e �]�]��9��с5F*-Z�β�ɤ��TU���M����v�[G/bW@A`%VRGt�A��.�v�#�ޅ�U��mL�.��Z0�W�&�F�� @-�T��3I�Z������/;��TL<�!��]�I٩�[�T}i�ՙW��5�殶�m8n���G/���[(�Փ���r�k-�ˣ�z��=5�16�K���wh;r���B]�L;�`�/�g��1u�,m<�"���m�cI�����[�}�%&��H��F��E2y�ι�o �qX��q EH9�K�[:��n��?Ck0�ճ1f��"Iqf3SA�}ӘQ7>ꚺ�'�4'r�15(R��7iVxϫ�z��j���a�iO�tjz�_`2�vh�1����fE��t]Ԉ�����!�Zz��kP�v_Kt5}(\�۸'.L�,�x��d}�tEw�R��Y�͕���2�dE���Սz��<���a�|)i����Wz�-$C���5�>���
��Z",TH*�Ŭ(*0QDb�EQIZ1Q����,T���ڬX1��"#UQX���[kE��Q���E��

�1�U���EI�Tb�PPDDX�X5�XQk*�Uh�DQ�DD�2)��.SNh��Z�	iU�QZbD�"�*�*�*�Qq�EL�਱QUAUU�*(�(��Q(���P��J�eE��DWUcQq�E�����V6�Ar�U)TS�b��Dq���Qb��أ%KX�����6*���b�X ��5�(�,[K�AW)U�]YQ��
��"�
 ���,kU���[QR�Y�Db���#"�"�R(ŨT]5�*�X""�X���D�QTDEPQDua�*��ժ�E���t�"�2��R0TA�(V��DT+V5(�UU���(��1Te�G�_  �D�X��:�����V��Z]Z��᳨�eKO��x'f��L��p㗚vFTV�T��W�+E�A�����z��*�gU���!�nm�lWK��z������⨻j�����oOy������'tg�����8r�<d�)�[� GZ��t����}�qI��.k�ʑAj�!��4���Ϫ�Yv+��
�(ק'�b#��[�Y�t=��k:xt\����^C	��qUį:�ĥGh8<n�\<%r\CGjd��T��mn�lVw0m*��{�{��ɨ1rP��n����NQwGN�ӿJ�Z��<���r�F9���Xn����w�C��b���WZ�˥�Ж%g�!+��$��-ٲ���=�os��I|���4���s;p��^;%��18�]bi�3�xC�M�MȎ)E����z�fݎ �_����φ�ez��: ��it�M0z�Kh58Z�-�Ӟ��'��T�4�H��!��]�2�e/bc�S:�7$��m/�ܢ����iGo�{-�3��C�=~K^����M�>_(ee�\�%ɘf�ݏ�w�̃FZ��Š�*��
�**���r;>(��#B:=Z+̉�!�l}^�����[q��\C~����u4����׸�����8<��r�~BZ�'�@�>[{�/={#�T�p˷��pY1�->�&�h���m�K�*rМ
t������GP'Y�����
�U�)�$ʻ���BP���;�6%@��{�G�v�v����K8/��ta��qJH�b��U����W��t�.��:ڇ��ms|{l��S������}�j�t~導~�Z`��v��_bN�*�P_/ja�}K��s#auc�[��<�Z+_X�+����<���=+\Ug*֫���k*Ǹ*�Ю����8a��A�[�=Z3y·��?~d��W�����)d�6��S��I�c+�w�Y*�,�w�`������������k��1mϴ��6<�>&iV)ChD9�b��Q]1䶥X�]��h�{ܻS4��Ҟ[&P�Ğ0�ND\:;�78�>�wl��"P�Ah��υg-($�c��a�J�t{m�{������3ԭ������,M�xpvY����?�=�6oZ��؅��%ܚ��>t*��s�^��lm��0z��4��=e}5�=��"�u.���p�P-���,^�Pоt@����fT��;7$;X}� �Aҙ�lh�,5Y�弪�U�ӽx��<|�ъ�hޞA���D�B�7&��D�O�UL���-7��'�doNl
��kzj�;��^�mD8=���w$����k��܊��+k�,:*+����\Q6̬ߺk׷գԳ@����&7IK��_��N��zl��]��gE��\0�X������P���8�C��3�N>}��Wݞ��L��JKxe�ҡ�P�)�u�J(UJAi��"������0)Y�5{C���Jl����U9 ��!`��a�L(���eY�?}�),��Y��:�DRx�W���=7�q�T��V9�uZ���"w�k�| ���傣��z2�]�cW^�7��;x��3d;GVa�e�oPy�BῙ���Є�怛-�caᤪ�]`��h�rt���1y�%�ݢ���n)gv��$J�K�e���B��a�2�j�M�����z|0Xc�$_��u���x�-e��Ք�1�U�YS�M{"�BV�̈́�՟{���qx6����9��l����;�����Υ4�i1~�
d���%��I�9� %��i!�2�|`y֧wJ�UCY������g���1���r�b��ܯA��n�yE��쭸!+�W��lGsr	�i�eL�����^�ev�/՝ki��$�(�}T}�z�=W*ܵ�hCk%-�;3Vtɢ�>�m"w��L������׎�y�vqdk�3"J�����t����s�D�P�G�AU���m;&S˘�Rv'o��L��٢�P�L;��sQpz"��T��y�f��.�~ ]��Ytʶv���e�LeB�aW���-�Sy1=|�=/�Y�f�=�����'*�{��3��@�g
�`�P�������X��~�'�\j���՜k�y��j�{��=�c��͈P�}(�.� 3��i�j�c��3���3�|3e��A��x��^�S�̪�r��.6�}l/�&�^�r��H#���j0E�����g3��>KF����N�H�^!ݙ>�PW���q���F糅�3��K�)6�X#�r�]��w������2�*T��_(.�����)6�->@��s�~8_����pU�4�s�`\`�u�(J���l0x ���ܚ��J{0�8=�M��b��uB��́�ґU�Ր�o��9�a�n
�[� ����d�ր�VH�MҜ�%���
�Z#C��kJJzm�~+Ʋ����S��¶�"$�D�zN���%q�.��ABa�ν{�Y�2����7��E�U�:�L_�l9y��}��:�>��kT�`_���9''�f2��pJ���pt�4�M7b:�7v, ��Epk�l��nVo8�5��8Mc���j��lA�`��8U��_&2���گ���t�<��%��#*i��]ELk/�㛵H�nIv]=�{��Fsͳ�ǅ�g�	+�����۱����K׻��dGZ�4���:�b�3��� ��:�5���rz�qѸ��X��Բ��ΊL�	�J`�J͛��+8ɍ1�W(/m�	���xR���#Sŉ]/��T�L;��q��Hf�Y*Pl�N~��Ը�pʳȠ�V�jP�z�Z Rd�*��^]Ƌ�q;���:��=�:�@ʉ�N���`�#���Cj�u��	�2�����J1(:�Bsx�ug��R^�9w��J�}��\�����{�.|N�gĊо]��J5騞K��ލMwt�V��y��Y�G
���0�@��c�^uɌ���.�C�؁V4���`��pg3��O=�I��ʕ�o���������t�����R�l>�	�O�����:�5�9��ݕ��u�vȭ��JY���򽗿5S�0��BL<Rvº;1^����8V�g������p4{/�t).�:Κ�Fi[���K4�	
C>���t@q��Z/)R#����Ġ�>2�]hB �fNݥ�>���w[�]a�u'fJӜ�j�(�姷Dy_�`��S3�w["�>��7ꏸw8)��
Ծ�:��ʌ%�(�S|���Q9G��-*�/n�2ɝqP�ծ�mGۃO����h[ub��h5گOZF��5�1?�b��i�����a�÷�[w�ΝҗY���e)�M"�X�z�����O���������[��-�>Aw��=w�.�}��DB�<)}%e�O/�v_����΍d6�����n5��?P�^��ѿDi@j�Al`�:��w�|�GM���E�~�|�q��(-��9�ZC���A���o�Oא��Е�J�`N�bB��v�Y�G�u_�; ��h�sJ;��6u`�3�0b�{�$V�u�|)�=ᴝ��b�&!��:&}��ܚ��FSz��c�}v1�:ط�ku4ڞם�X6��}Tsx�zo��n��c4V˂�;���V�W�=s������hji5�zMX�<i�|6�Ί����g���~ૂ����p�k���/h��ғ�/�h�ݒ|8H���L=4�y��:Ag��R�e-L]JKG����x�]Qo'�qhٯ!x-c�XVL��Y�z%�P��^��1��>�(:����{��BU�Z8J��KN％v8(�ɋS< �y�g�R3�=�2l�o�;��F�Ws�f���ee�[��D�a���N(�:�36:+8�C���/u�+�in�#���Kɸ�ʶE!������7��?"��]}���zm��H����f\����V���;����jwK2�Zt7;i-�f��V�O�,u�љ5u�B+���|@��CLTMR�	=G�'v?PsӔݗ�}@�bg%U��e��z-���(�O����Y�\o�^LkY���e�m��0V㏙_:��CNxO2��c*��<���e>ɕ�Z'���a���]i�V�n������.�(�c���5WSfOx�7�N����O�n̻ۇCᚽ�����q0�}�7�iET``t4�[�#��5e��k3�"���-��ҡuw���6���L�������Fg���jA(��䶍Z�~�L���LtW��a�4�E����xi�Rf����2��0�	)W���&��Vi���TL����x�`�i��H1p���V���h���A���O/,�f����ŔfM���{G��a�*ИK���z��#!�=�%es@E�<6 ��|��+
��52V�f���O2
��U�Q�ۆ��K����%�K�-><A�&��{��0�^�4ȠwyviO���$��dӇ����]��Zz���y��f��=��������~�@ow �{K*�%�aҡ���sO5nsc��I�NY���^j�r��rYH��ϰ7N��E̕�ܭ
Fha�[G�5u�j�
s�g1MY�&�=o�n��o�:��p��+�(�����:��+k��F��*��N�[���f�V�6"�)�u�p��,��yoS�\9z�/�W����ӡMKA�>Lg�АjW�ej�'���~��Wi��^�����.t�o�:�My]g�s�?&R9g8��c!,��U�����1/ ��S0����	_=��'�tN���eE����+��Y�2<�kɌ p�����Or�\�9�ݧV%
�������J<,�e�����4���i����oSB�9\V���V�}މ F�Ḑ�5�>U(1Z9��ۤ�i,0��.�G�EO<�V&g;�]Gkq�{���{��|.p�u�A�C�x��'�G��.T��ۏ���<���͠��Or;�48k���k���Q���~��\�x���z�� �[ݭ��`�7�E��H��f"9!�-T[�s$��v�I�J5(�n��N-����^lu������`t+�����{J
�"�]��	�>���(����s���(����wn�Poa�kd�C������LFv�q�5�E�.�.D�s �\�;	͕Me�����Y�3�wNY7���������S7�K[`�\�k�b���;�nqT�j���f=�6��u�t���z$�t�Q�%���P�'k��E�7/ixbHx��}�0$�@AN���z�C��~��I+��J#ji3�=C��QU�P����i����'S񩖩񕻗�Ɵx�쮫��Ҭ7����X�r�O|���lKA}�]^�k*l��f(T��f	Dvy[�X�^�DS���Y��������n��X�L����y;"���x�W��Lh�˃ �f�nUǶ�%�%��*�@�ڋ�~�5�ό ��Z���������/�?%�CVl�v���w%x���t#�y�D�n��Px�sx�cN*�Tݺ�C�������pA�	��V[i�Z{�b%�ϐ�\>�z���?-�U���\'>�����g�(�1����������!���ݕ��&%�24kp�ƕ���Ȫ�j�(p�,����b�][�+9��y��'Jb���$[/�̭�1��*��,e_Z��¯���\��%|�[�Y*۔������wd�0p>�Tĩw�o*��b����Օw�,���O ,�����+2�9���5���I�� �0G�׵��W���n�w
�0��pl���Y��5�:7�B���w��3\FQ�6N/@[��v�S�ݷ���DKJ��N����|ࡼ���5H�ݫ�bخ�����>���L��}����Z�Vլ�9�܀Vg���w���ʡ̨r��^qU��φܯ�F,�>�+�����8Ż-w�����8_��C�ʼ,l��@�ѭW�X�Ĥ=�.��>�ؿ
�������a�7:,�����EO��0K�W�Pk3��^�Sي��s�WZ�pj�����+����
w��q�A�A�v0c����3Ԑ�+�α(��<���%u�RY��vY����>��p��z"�;EJ���_�r�Vڇ+Hw�2��8(��M�*F�$w�2�xCĺF��.�,e
C�'I�X#~^��|�Z��ya?��,�� �W���ұ=�v@��&W�5�2A~U��nUu)�[�ʾQAb�sˏ�Y�f/{������*4�r�Xu#�EH�Aʎύ���MGG�����l�x��	�������g���v_����g�G��y�u�e@������9�G�VQΝ7��sj�u<nty��3�3N3cErL�W�%������.�ۥSáj�N#k�>���uN8���~��(��,N�ͧ�Q��}KU�v�J���V��/o�������WZ6Xk����J�uN �it����C)���|J�LE�CW����喃��Fͪ��+����C�c�h��x�A����p����\�Ѡ�|����,ma�!�N�&L���72�SDz+"���$K�-ߊ;AU�ֹ�]DN
���T�e�p+8�
�Q;��w�Ls��[�X���Öa�w��ܣMP7�1���d�Cl��Y�(Q���rj�x�^8q�f�v²�0����fӢ�@��{�&�;/e'p�Jp��X>v3ҝ{a��	�%���p�v��q�a���������w$�/Ć�k:ܮ�v��$mn �}،&�a+f���7�]X���1�a�Ϛ�`�p��s<��'!����C�ˉ��这��w"1h��̖kZdl5�y�N_!�w�7扅M�P�U߯jP2ϋ�F��f��(jIIw	�4���;m"�^�T�x-ܥ���k}�Rr#Ɋ�����m�|z8���]os�ǗNNww�oL��ɳF+T�M�yz��-Q�d�P����ʉq>3��T�,�=�hՓ�� B[۾u���<*�S��M�W���!ɛcw7ff9ZN���f��8Ӡ�_0�m̔��dK��V:�g|�z���Yp�����`A��e�e�w+��#<:����n�����b��
��,]6�@2ݭ�u��r�'���D�['�����hq���n���O!A�&�sTT8mQU"��ڂMdsY�$�4;�,for�c,3)�<�rH�<Z#���{����\�*롳�XI�vm�+�/+Y��A�ZL{YI̭�j�y��$���S�e}���r{	��Hv��� E�Uĺ
���U��;Zt��U؛"DU�:��x��𓝵��;M���c��V�EN�@���f[�����Id��K���0a�s{�((�Y�}�n�_�m\h���pk�E�	ՂmKB;9�mK�I��ׇh�ds1e\A�A��N��\��\֋��ѕ��$��0$l�Iq���+cp�5��O>��ͥ����iŨc�%��u3sd0gРP�G�z,~d�����J˜��ko�^4lM�Z0l<e�)�k�@rܜS�u���r@�"Du�E�e<Hщb��d��ky�jL�}�@�[���WLo �y[֫�ʸBՓwO_�@�8��������]%��ܼ�/hl���K0Q�� 	���!3:�[�z�ۄ�(/Y�\a�l�͔6E�8_WR�j�vC�St�8!A�v��l0L}R�w��//]FP7Ns+34Qt�h�� 9+�M)�!���*��2��uVfX�-�j�cjV* 
  �}B.o& �j���U
"�[S)3$��Qm*��k*�(����EQ�iDb�X�������4Պ"#cY� �Z*�e%Tb1UDF1L�
-��U1ժ[F1����Ԡ�ڊ�T���`���U�V�PV*��F X��k
�b�(�WQX���cEL�EQD#\�j���JR��+*���a���UDEEb��*�`���E���)����� �5�`��UQE"&R�AuJ-h��Ȫ���R���
��j��-�R�F2"�YC,�X���n�+���U�Q�D���*�+��X�Z�j1V
*
�J�r�Q�1H��2��$`����$��M���բ1EEb1E�+X�QDJ�Z+���h�V(�Tdb")QF11���E�����F��\�V*"jߟ�
2�qڜ�pm�ѦX�hm������L·:�'l�Z4Y�3ZO�ŉϭ��C��u����<C��N"vy��wY_���]�a_�d:o��r���LP�pW��ނ��A����'��ΘKNwr�C��N�u�]���K﹈pE����M`o��u��ZGzǞ��"�H����ڽ�Mp�w�뇓�K�k�e�n��s�%[}K`^��]0N�V}�j��IO#�zM��l�ռ E/�������Iy��C!���־ǆ�|]X]�q(f��R��!�R��I�~��v^[�K�۬=�:r"�������q(M��I㼊�����7���n�\�{ϻ�b�����!3���+႔�)��ӈ�����fK�j�g���V`�ީG�&׶s�½@��_��<���N�s[�>Z����䠮�e=�tR&������|Q�J�h]C��§D���K(u��T��}�<9̞]�H�q�a����/mh�^4���ϱł��D �4S&|����̓�U߅����p��a&F�[�{}�2(��P�Њ�>��Q��u��UJ�G4�x]%kp����=Yce��a�Y�ľ�A�:��B�H�W�0E��e��e�bXZ�;5�[�{�h^`F́�Ǣ��S4�O�Geu�G7t���;���Wڣ�X��L����BZi�쳽���������C��6��śΈ��v�5ӳf�t����/p�}ר�N}���U�1�`���*��������y�v.��rU�C��F���!��UwU��9�"���D%��F/,WZ̖�4::w�� ^�Λ�A����-N^g[��и]Z=�&��Wͩ����o�A�߸0΢N�� �^'���a���2z�*ѭg�b��m����A[�I����2����fò/��ݍ�\:Wrxld�[��3�F��8_�~�6q�Ϛ��O?�J�v�Gu{"�Xw�y&Ҳ��f��Pg�W�h&U/��Vj��I�����R�f�w�u��n��'����MF�#^�ӧ6<c=]�
_{UU��K��w�o1��t�糥j3�n�W���AB�B��w������߲\%��pBW�Z�	�>�;�M���Tf�M;֎�w��X�
|�#h�Be�G/�����UX�d��x�M�&}s��t1檗2�/e���|R�}�=8�;ZC�������s6�U�mq.��-OVJ�]�{t����	w��s�{�ZS����ܭzwA��N��VO8�`;^P�/�p�ߞ��HP�r��&-�C���2��Jա�M�P�+��Ԙ��^��:����h�e��,��z=�\��˴���ȩo+���= J��]��+��=�m���O�����LN�p�ux�@A(J.� ����L+��O��v�D��c�-	�%����
�[϶���Kxm�
�}p/�&�^�p[��+բT�����r;����mjeJ��
��� i�^��w��ʂ�u�{9��6���]�R٫�Ǻ^A(�\�p>fm��{r+išT0/Qϓ�(�Ur�5nѯovc���Ѿ�Vz�J�'�]e����j���4�r�F���SJP�%��E=��Bg�5}k1�|���lUn�S��M-8���+��|C�(w#ٛ�4:o�>���R�0��߹�J�/�Nb&��I�7���;U����7M�ws�x��-�� ݬ٘�}�b�������F�yQ�A������_F/��*vE���N�{�{�W��y1���1��ݪ?kj�>Ҙ�������T��Y�I�jų+���D!R���Ǭ���w����	S�ўW( �up�]U^�:��=�1ڶ��W!���t��U3��j2Ǽ��טD<q-j�ެ�(��(�OnQR_����(X�(��}���6������p�><t�:�\��Fη�k��rmv��3�n�rvX�3�;��Ƕ�=Ѳ��dr�;%44us[���Sy]kW�[&��;�;D�)r��`�]k����e��AU{m�N-��!��Q��s���}z���,9��Sd��_�"�.4��J�ʳȪ�m��Z풨o=LN�J�ۼ$���v��>�>��Yɕp<�t7�}g�]#�����xc�n<9~�R�g��{�`�Ϯ3��UUK��{�1s�X�t]�}w�*˱\�|�͵R{{�1��j�'�b#���}
�';�}R�
38��W�rc*������>u�^�����,��W�h��d`~����V(�1S���q�����I���L�(�ْ�`�#�K�R�,����X<L��� �������l9���=OD�]FtK�je��l��R�@*��˼�و*���Dr�zL>Z%x�g�Q�^�#�M�ҼܳK0X����=�V�l{�ׅ@c�ՁL�W �u��Qb�J�m�+/��0�=Z@�\G�F�b{��w��]7\�^2�k������gS�
iX�Ŏ&�����mpPx�A�mz�&�D"��Z���<q%gH6'n���tpvKuݳ���y��dn���Pר��2<�-->t��d��Z]�Md���V���P���e�u����K����ڛb��[��t�I�Tz\᜺�Nu��汒8[��<�E�t^Qd���]	�z��/Eo��h����_רdb�,�p�E��WQۮ�U��z�9h�M���ףy��ظ!�X��P�Sh#(t V�#�EH�(�'���#J���77v���m?d��;�i�!�7^���o�j��|txA++�'�0Q���Ҩ��WGVգmX�3<yzr(X�/u��-1���7�0$����yLQ;�Խ�Z&�hޫo��䕧���X8M�[�"��6��;H�8 ��IФ=���0�)��ӳj���˵k;����xs:$qxW�s
ޫ��Q��F_Z��9�J��R�({oz���d�5ic0�F�d�we)�A�[�=�ϪlU�W�pM�SZ�����7V�{o4ֺ{���z���a��7�ŉa�?d׽/�cw�zBPXA�BNu�W�F�3����+�A.'��r�=����
~3~��|7�{
� �Bz���]���ݾ�%�;Ew:�Rǒ�L�K&'s~8�P/�9	�ۗ�y���5yJ��"?�QrF��;�Y�Oc.
�j~5&_�rT�y��&@�oH�9��x�����|�VD�V�Q�ܭv��8v� �{p�L�k��E.ӳ.�p(���ۓ]����;�՘vڲ���8�3;q�8a������괫}LOl������:���Zo�Z�U����9���S�q�`ϓ�i��j*�x��G�đtN�}�f���:F̘j�@�u� +�U�����l��7��ؘ�9 �9�}��|�ϼ���s�ND�^��U�&J�=T�T��5�������^�I��8�y_��~j!�9�罂���AE�k�%+G�=�;��JX�����{��s�v.�>�T�=3>�@(p8X2�*�%ר*���G|O33�&M��u�����7�������KE�C�x� �~3si���:��%��/{L��'��m�����C�UC�dҩ�����lf��a���գ�e:U��U�Y�#^�q2vs��B�'�����
�B�Y�i�xcHu=�pV���ճ�g["$^�d���|����f��>�th�$�mu�U~����BYR�}�����ˬEy����݂
?f�Ǔ��9�-������.��_h�*�k	���-
�Xu{����:b��B��j�Kp���R��a� �nM �8�(w�̬����u�ŧ%�����qJl���?˵�zpU�~�!��O�v
u��M��ۮ�`����i\�]ԏB���}[a��h����_YIvV�ݾ�yde�'��-�ph��e,>~�0� �E���>�Q��GKg����e���=�9}L�{#�|�ۤ���e'h/����a/�L��xO(��j�8o�Y|h^�Eh�y7y���8��9�T��|*Y�l>��|1�K��^�P��O_�3W��7�gĴO9�S��ك�q2��Ư� �Ң�W)j�*�`f�b�V}��	�ٻ�O�a�o��yDT���{�q1q�`�ձ
*�z��������5�c�=Z��p���+G�%�\6|s�Ƿ�0s�U�Ϧ��\[�׺�w�Ճ��W˔�V�A�ެ&��"���ob}��&,[iEӖ!�a ����� Y�{���=<����LFla�S�*p�rаϩ��%\�B�Y�ο-�mM�h����b���Ù�]��-��;�U\�U�W���YeR���bܦ2�ҙʯQ�.�8Ҕ%��zU��
yf^y�uޱ�'< W-�X��Gp?�_aB0��K�ۀ�U�a~��`Yd=;\�݄����E�{y��)������6ebe-��&s��{��vN
��Ќz\*����Ҹ����jQ<��7P�Ʋf�C�
F1$�#B�}.�\<�n�v6�je����vdIh�L��{r*�����6;����բ���\�� �i�\��k��K���F�}wfL���>���i���pxT�q��zͬ�"
\���+i�)(-������x�+{:����Wf�;�k�5*�)�FVV�BZ�"�|L`���aX�jH4=+q[�C7�ç�X�����幔k��W�\��:�y������L�����v�_>�D�}��9��I��ܚ�*�=�-=�~^W({L��n� ���E������ӯ�yZ�"��>�^��R��K�dg�_�������)���n���������xU��r���m�WK�u��Mb���a�eOHz�	�V�B;`��D��_��1C�R���*����iW��2�����TR�є��J��^	���Η���P<�$џ_Z�8W�N�� �5�����f}��V;E+K��Z�b&|01���o�|��ﻗǈ3��]��J�Cx�Dm@�.y�
�*̪�y`��>���6v��0��z�M��\� tS~1�(,�V�0sg���v��YC���ͧu�g�ڲ�}�{�!�)��w~v��H������=Y��g�Qk`�~9�}��Z�}3����Φ�ݬPj�ru�/��
��+M�f�8���&�׎[J�/^�w�u�w��Iɬ��v�(�5�}�hG(�9J�G��>�|�}�r�U���w����σ�u৔��;����HH��"b3��n�nӚ�-r��+��)�-�W��\N|]����'MA�+Wk�;<:�J�bv��x�;�pm���]oɦ
�V**v4��W��Yc���KGa��4]w���쬋���S��9^��Vr)���*�OX*��,!Hx5WzLJ� �4d&rMM]XN�u��ba�=u�9�Eݐ$t�`�m���e}l@E���)�I���k�k	�8orV��Hi8�e@���v��_?���C=$Z�_xQ��gEo��x�y���bS=a���N�j����p�ԪT�@M�b��]�Ԭ�u���Z�$�~�<6���,���4vϴ�>�tVc��5qT�h;��ۧQ�BwV���^�"���Z�$m�V�٪ʌ���m
��!���+�v�W�zBK�C���f���B�pc�s�=s���ڮ�MպW����GK���ͥz����=fI����� �,en^z��m���edZ�5�����oѡ���Ǵ��kT�״I��ȏgX�YI���r�R���\�RuY]B��ǽM��9���mu�C b�agl5�u!3��Ь
�e<��h�!E*���FЍ�"}�9 �#.Q�u����Q��:�-�v��C٠�W�G����c*�pH�g��j�x=�睃C�>�r���D�pW	.y�a�v����AИ ��Y�P�9a�ٰ�G۵�{hz����I���^m���q^�b��7��ឃ8O['��D�ed�5�Z�{�娞�C�iE0Oa�2���ű�3,��y���S�!H�zqxJ~���u ��0�T��
����R��j��.'��iB�VK͛ ���J瞲� �>�-�Fע8J VPc�E�ʘ��u����qf/o0�,�0{�j*�kƲI��S���ˀ�00:K
 kv1Ku�h���.nt;�.���(�/M�m�>D��ЈT'��~7]���P9��{���dޑ�	k�gu
0�.�Qj!�՟0r����2P��D�*`w^���2���YÇ০t�ܵ�����A-���=�|=����-X�!ý�h:�怋��6�����#�م��������7��<%0���cL�g��Qo �D�)ۧ%�w�#F�o-�w���$2��f5j}1�/Zz(�N��ͤ��E�]B���1������3��R<�,wR��t��E�7�=�D��Z�?1�XKt�U��+����:���ۥ t{�/&��E[�A�!:�ފst�F�+z�V�>�O/���g]�S�u��mE���8�3�H]]pb%�|vcTO&�{�7���*�ԛY��7yp��ܦ�Z�M�8"]$$g/�\y��l�f�oNಁ�Wt�Ryǯhc��Ǭ++t�LW=y�f�.�j�uv~��}5uB}C��n����W��A���l�:��pR�f*�=�Ԙ��s���� ^��͗1D�V�h�Q��8��}(��>%)ȑ1P�^jԶ��'�R��T�=�f-�&�lۚplos��d�T��&MwJ���(L�(�ܻ̻�]��Ƃ[m�v��!;[�3���]&�),Õ���TFㆆaj	�2|m ���Ő+��d��:�jC�V��-�Hfv�LN����6Ú����AYʞN-ԃT�/a������)^6�u�L�UW��·.��IFM��v�}(Lٕ��>�(���W,����B8+2EL���@�A\�.#�h�4���+~@K]�fo.�9�I�eL��. ��6���1��ְ�5���������*gd�Fw&�uW7F�D�d�W����Ak�v�ǐ�����*��ȭ����h��t&�*�[Z�X�轙b`"�bm���F�$��H���gSƛNƣ�Z�ׅ��3YraB�h��+ZÜ{�[V(:Fb�<�m�A
��s⮖����=�הks���jJ
&�$����~T�hp���Tov�zBfI�U�nJ���C�]��ׄQԹ؎f�}�"� ���v,-��'weV
��6:����]7����qP�S�:�fwP�h��-c�D���h	u����1q`q�`�Ma��J�'f�d�����e���}ɢ���r�d��5���K'T�����b��]��aR.�.�e],`��P�Ap��b�Aˆk;�+��6.W��ҝ����E���85	�躅m��u�_h>R%��)�zf@�L7:����9Ϟ���Nb�8qF7n�!���p!b��To:�3ݡI8:)�,�5Iܜ�ս��}+B��酊��5�.^�-�gʔ�L�V$yA(U�I[-c�/���PoQ����?��@-��K_IpUӬl���r!zH���R�p�WڷZe%�n����g�inaW6v.�p6o��AJj[pt�\F*�T��ס�&����b����N���|�5�Bӳ;X'4��wYzV�?�o/�=�
"��F#+U���*�cU�f%eX��F
���)�����iU"����ESW0,��(�E��DQ.�(�2��,UQ(�S*F(:K2�Q���*
ţT�H`�Em.2ն(�R�""��Q��k
�T[k��Z�R��E`�*����F"�FbTDr��բ������EEEf�Dբ��J����҂�c5q0Qq.Z���m331��Q+*+l���
��Um�)Z�kVZժ�[��fZ��EX�cQU-H�2�2�Uq�X��`�����&Z��e311QAQAE�W,�U��[]	q�T���*9aP���EDH�Kl�J�bň�lUF*���b�U�������"�bŨTj6�ue��AE��1UX�TPE`�*"��V1�����)n8����-U�ʭTPj���+C��'l�{��G����@·T�l����5�W���tw�ևSۻ�I����@��f�=��u�O0�x�m��o;�6 +�pQ��D�`U�ʯ�v^_Xt;���!ʺ�n�
S����ݑȍ�e�x���x��]wP'�d�p�m�����7a��D����ݭ\�tC�d!,k�jbm���v��P����S�sM׎Or ���h5k!�p ����/To��p�َ��T����«a��{���s���.o��t_�׹fjPByO>����x5�薄1��.P^ۀ~���퉕s��Dei]S^WY��A��ɹP���bRL�-������gz�u:��9x�8�<OGu�b��ʷ����	�����]U�՘�lCή��r2�CpK_��F¥��,l9Nw�?WOMȧ���_�N0l����f�+�(1ɤ:�*.�("k�U�+k�b nP�������9��A6}��/Fw�
�-��c.�o�<N�	�*V| ��)UW�;Q����s�^s6V��%�9���X�[�'L��Ǣ>0JI)DX��5g.�;�F�Ȭ34�Ut�ci�.��u���
Ԩ[\5����&�6�v�`��`z�9�Vp1�J��[Y�t/o�.�0a��֫,��\���'(����"=����xw
{j���&&�~��O����!��6�<Mf#��U�b��FL��(�<�R׎����h�M�0X�f�wDζ?U�H*&��b��I�K^T��X���u���N���u������������|�Hp_=
�}tj�2�g��>��x�<��(�)�s��v%�%�]b�	r�*�Z�Ϻ�I�.�
�/���:���8g���j��I���9&��y�߳߷������C� �۹VC5�E��]���_a��F��a}۔��c��e�Fk�V�K&�/��Ȃ�u��_�̨�
�w�b��z:%����.���<n֧�_��6=�� I�}��9��dt���|J� Z5u��&�׎��/�0wc��l��MY�ݫ�	��?	�Z~�>�YB�F�]C�����֛���V&e�K=mp���=�]JY�fש.��+t�ۂVR�� ����Ω�3T�V���S^�����rw��{k�t�C=��l����E}��a)��]��ʗ�Ŵ{�Ou���)���w��a�*r~,zt[f*8�AxҽJ�#����Z��<�&P��Ckޗ��2�hШ�����K4N�)Xf��[��5��=����<����g�<lb��x���\�R��tLr��4� 8oc���edȅ[|¾�-¬��߭�.+T���F�#�MoB�ҟ�yR�`�R��:)����3���=�f ��{�5y\��+�^��R�2y�+~�����u�#R�!p[����p�~Q�'�P�۽��!�.�h.���;Ol��~��*���!�dJ
3��'m����"]%��7��y�ޞ�t!��g��VD�"����[^Oڲ�}�{���GY��ʋF�[�Ȝ�GhJ2�2C0-��(S'��/�y�
�E,~����ݥ�缳�F�}��*������QW!`��v�&R\�?����ɧ�a6W67j�ܺ�N{s|$�C}�i�͌����u��`�ub�����z{2��{�
~y�j�L����&w�I��Z3� U�6��;SL�Ķ����@W�"�X�{w����SeiE{q/I@��l�A�;L��Ҧ�LrR����R𲭈��T}��w��hd�v�_f�C47���m*{=r�}j�@)G+��W�'f����D��~�	�v�o�+2��D��Tem
�ץuo+֌s�w�K<��P��w���]�[���o.P�sD(?kyxD��֤[Yʟ��D��ƾXB�۝#r�	GEgN���;��jN��N��ʹ�-S���j��r�k�\��n�y�h欬&���~��%�t�oX��*�J^�S�{J�6©PwU��p�/���v�xV���7��7�{�w�;鉻^Ȓ�k��>�>���9T���]�c�O��4�7�H位�8y��xo)���^�5�zYF���VCcl�+�bN��Un���,��t"}1�u/��	������ٺ^WR�o��<"�����8U��w�p{1��?��A�t+�޹b�n.K|�G�56]Z�H,��ԦC׍�>��Zg���W�+,�6���.ז�*�q��BWy9���-Ҹ�	C�����iH_f�z�jwʖ�k�R����dI��l���c^�xg�".���_x`{��v�,9�N7���,c `@=��*]AQ/O�e����r�2QaPBe(�1��u]���U�z>�m����KVfW�W�k�ST~�~.�x�Mo���|5{[cU����#Rsr��5>媼�&z��"��.����
*t@��c�
��&_6�9�"�f:������%g������`���5��0zH����̊d�(�{5�驫Yt�N���(̀������!�/K�t��!r���݋R[��/z��Fc�R^m�s���\���C��`���V,w�Z{���©�2��ΰ���s)_����,%�:"�a\�~	�*�)��ʤz�@a:�7L����d4xb�w���sǴF�5ᨣ/��>E��W<�L��6�U	�J<�x,ʺ���yH��nw����#w^���w�m�Q�^��w 9��.�QҨ�K����W�a��E�_�(���bDb�7̒����bZ/������<�ޫA�s@@`�9z��9�����g>|�P�=| �N�7d�*e;�av^���p��{���.��YU�y#�ΰ��������O�O�p�(t�=J�,�_��J�Z��>-���J�
���=����}�f�t2���z�;��'��T�[��C�Fɱ��y�ܽ�X���J�b�U륻!�e�~�8����]Hi��7�1D��r���Rٽ����uqP��h��#C^�e�-��d�����:��w�t���X�PU~� ���l�o��D�{���^z�;�=���s�CH���$m��.����*�p��O}5��r�+����������<���l:!�z��hv�^>;�LR�Y�7��������҅�:�<F��ȴK���wo:9�}�$�q=X],rq�W׽P���b��^��ho�/_m�(W66+��7[b�b�q^Mo{r���6���F��v��.aO�]�*�G&�0�,:��s�f�	)�u���o	:��I=���z"��o�Y�1�f��W�g(*���>��xpr��x$6Λz����nt������\��0k����f�(�rj�P�E�e+��R�r��j��y;z���:e9�m� ܀��c�O{�������0��r2�*�!B	C�z�� jBV\��tw=��wG���F	�ɑ�.ɢ�,sB2��BL,��]�}
`�����aE�]�������(4��0ϗ��c>�Ar}�p�}�SbT�����$�IX�~����{�'�}�ʱ��((��>��m{�C��`��yK�]53B��}WS�9�`�X�	G�n>����eW(к��`Hk�a2��6/�ҿ��%:�*�h��>9~��ɮJx0�uσ�C!����еS>��O.��2�qR����{�4�JI���_I[u~2�ha��iЃh�^')��2�xQ�Q��2���(/����-˥�V����z�	�Kv�/{9\9��dm|'81{��ABa�;ӗO]ݒE�d�~��l�P�Hm��4��݄��;�r�Gj�Pw�d3&S�a�6�T<����f���]>��u:��cY/���w�M"�S��J���:������8�d̰a��'0kV��|Ռ�k��R����]ע�w5^�[�My��>GH��%u����v�n��0me�b'i��g�i�(��v*�U�7�S��5�nr���]�nt7���k]�\0�gS��pS�Z/�Z3��	�%^��):����\��^����$ݹY�jxxeTִ[Ux�/u�UY�UPt+T�C����*�v�J�]�dʠ�c�D�w�����4}:.�)@��gF_Z�8T����|,5vS�<||�;��B���L�豓*����	[>��ˬ�*_���AV�������ՆϷ���ԫ���������.��k��O<R��(\@x��g���tM���5��N�q�R��F^�8-�cI�����ƕJu�Ѭ�>�~ �⵸��Zs�m�y&m-5�-KI��Ku{B˶9�]�w+��*}��}/CP�4S����Z�%����V���i`藞�<+�YK�]ENƃE��!��K�gY�P'�s!�0�̝�� ������HAΥ����s�E��LK����:]��D?`�&{ԑ�_��oM��܂��&bPgE~�1n+�qM�N�J��/���	��X��v�B�Ν0c[y�r��SVf��X�;t���m��-ka���K��oZ���{v���P���u��`��V*'cA��^�Hp�ڮU�7��Nn�N����פ��i������ �~���p�Y��7͖xALX��������������}�E��Fu;P�"�kqQ%T��"𭛛Ydc�W[�i���)�r�hwk����x%J(V��}r�՛��[��#:.Q},
��t��h6�^��ӷ��&�5�x,�g�őa�:6���J��Bq��yO��8,A+��9�m�}y���זM���Q�7c�G��d�u�X�Eg��	����_ٍW�ؐ�m��k�ȮA�=䏻��o|5���#r���ѕ�V��}ѓ|?��(b9P�V����3��j�Z}���8��x.|�P���2�^��ނ��B�y�R���Ǻ��@�k�*��kU��\�]�_g`����x��T�B��ːƜ0�)�b��:;�eM���f�Z��:)8�~�q�>��̘kB�3��A���Ue�`LF��|D���ǜa3J�~�����*Z�Y�+�^[�Nͮ��'�ը�y[^���6�"�<�O��'�ꦅ��tme�M��mDg')ދ���
e�OLBE��L�x/��G �6��&xJ���\vt�T�7	�d(���7�U�k6���ѭ���p�M�F��?s|}C(@��A�Z&Іg��
�a�ݽ�i�~��ND\��y�c�Y�y_�goǥ�n�����5EQR� <2����Z:�yN>��AYl�W��~� b.;7�XU:�3�V^W�V�T��hQ.��߳�c�[3���gn�I$��-{v��K�zÖ�"ܲ62Ǒ�|2K�u�.�b�t@���[|��Be��=����憢��6邚�%�W����:B���r%�����ur�" Lk�>>{��Xo�/x=�r�&I�D)@�������_��s�OU�
���e��~S�o��Vy�v�w��A����3�KA|u�0w��/;�
��`��T �g�t@�-���Ҹ�P��FX*�Kd���Pe:9�g�|=�)(��3���;�c�	���(1�$Ž�j��V
PD��Q���Ed��< W�+�e�9U�KN��<���;D�I���nt9��2�Є���l�������P'���V��{k!릯�_��b�,��*�}���랼�0.�u��'|m-���r�_UX4X�?��4��ܥ/�
1IƭO�s
�L���*�Zv��+8��tx���vYpvH�6�k��"6݊�5;e��Ւ������ۅ>Sz1�:��n�=���Ya�W��b�oМq�H���HJ�'B#���t�U�<6$淋�h�B3uf��������5:9�w�[����Q)�][�`��Q7:������
Ϝ��6\�f`��0F���������~ɝJi=F�Lg���p�x������IG,����r��Ư�מU��*8��{����_^��9�Z��߱�%��m�	SZ���g��r��<�Y��B������	�{�ٖT�j��^2U��Ò��l�rn��aX�7��[3꛷+�[sOS��ޣ�J7��J��%[F�ǕeT+GG�(��X�Os/N������ ���}�;iJ��x���ge���2�;,P�P�Ͳ�)'(�.튮UW]m���V{|#}�pt5���Y��Ub9L�m�*5��i�ł�S�go\���PW��9Bؤ�`�&	�py*��4׮�N�W��NK�t��0��N��^b�%ό(�7r�[9��3�i�\/��Y���d\�Q���3��Ny�d�Ů#�<	��b�JIL�r^}��"�\T�핖[�]{+��i�:�^��GR^�5"dގ�:�;5�4��,v�#]�#�	�YTG$vv��.ỸB;*!̈)2�Oz1a@��DM�����O�vD衢}WV��v�p���n�զ �i��JqH��(���9[��� �sd��nbY�s�M��E�7lL3l�r�dԦ�4����=zg9X������QX����{i�Rl�o��#`�p�z�ҩ^D��p�l')�؀<�]��$��֬2VS� �[Y�N���:W�d�hI�����N�V7t�v���v���N��LP�%�};�Q��=����V_#cc�5F�pH���%�3C;��}�k��WJ<Χ�k�CG:Q/�o��*&���}�N����N�sX{�t�Y���R�2��m��1�O��{�߆r���$���e�K���tb��6�%c�Y�u��U��@���7������:�oS�,��5���9��+�M.��#�n��ד��m��`���9���R&t�i���.�<7[^$f��S6���D���
�-��Wr9&i��.�Z�cs-�[�l�Hx&�%�U;�K2dK�f��5��Pr�����K�[P12�t���������U��D���UMs)e��3�p�v�;[�Ԃ$��ֱc��0 ��{�q���+�F��4�����I�;��sT8x<��1P���mPaD�y�Xw�P�R]Eةn3CL��8rI%�w��c6����6&~���:HtZ���>�Nc��I˃�U�Q$�ފ��9�j�7wu	��=]��s�QQ݄o����u�Mcgd�	j㩮mݣ;{�|���^\���	�;7I|�v��x�ԑrW}h��_!e�;�I����gubsrΉK�2����i�/�q���Y��3)���U�L�#��ك+�뮙� _DZi�k3�S¨�5x�lpY)f��S�Pϯ,)a^��s�\z؃��`0��J��6s�k�[���ݢMG�=��Z�����J)2\j.���ȡ�*c��xY̱h@��L�Ls�S�,<�b�%���I�Z�%Wio85��v��5�n@r��:�1�T�y���E�~��� e+3Ej�;7$�G�V�-�v�^h���!&D�}ց�W���b�CW�,1!���r��s��Ef�X�����V��{���ݷo.4"�m�`��^�"%f�>�v��i.���1��djhmof�� ��fnub�A����)�K�U_(��[2ކX$�i���ya�H�w��U���qvm�X��T��j�(�K8^�s�wIe#��uE�1b�wK,񎎷�&�������[u��{)֪".O��^�g'd�*q�8[ǭԢ��l,E-���g��^W3�;�����DEF1G�(�8�DX��*�l��*#J���Db�S0�UUZ���UQ�45Md�A��QV�Lf0X����&��TV"�kZQDM7
"�"ʉD�*(���R�u�1�E�QTE*T5s*����ƈ�,`����Y���J��1%�E��1[jfa��ZԩS,VۉkW)T�F��e�EQ�UX�E�1�FщQb*W2��Z�MY,U+m��X����"�**ʹ�ƵB�TbV5-X֥Au�kEfDm���B�T[d�5�ST��(���+���EUMe2ڵ�TT�W*�V��R #QQ��h�b���ZZ�aH����VP`�iq�ckb"�iTH�[j-�J���q����m-�Jg�$
4h�U��,v���ob�m����S��pΣȇ܉��`�X
�ތ�9S��6q��]]�
��\��2@�g�g1V�F�[�}�����h�SȬQ�����F���Wİ�j>.����c��#�YGE�(��RǱ�a��L�%C��7�`�j.�b]+����k@��	��]�}f��lߛ�;�$2-#��z|;UY�Z�UK�B:�}�*L�)����zb��H�W�7����7���'�X#x�){����6��C�fО�a}�V�ס,Mk
�ɗ6�yI�@O�y�s@9�۸�k��)v�'�����	�ʹ�i+�6��?#�$�o63�*Y�Hӹ����3|���o��E�]r���T��o6�^CN��Z��ȕ��Y�H>�.�;%{No�X�J+,���]�Cr��}����B{����1'G�����<�����G�ߋ��'��u�OCՊ v�AX�nqUY�iЭ�Y039Y�������u��O�w(NP�E]�V��4gy`Oҟ��lx��S�/ƒ<�l�:�����=���^8r��2US�lz��s�T�}��b�b�/{0����Z�I���}�t�%�:�y�O'���{Θ��8�Ӗk�yfa��AQΧ�����������A�=2���un�\��!�7!�wM��j��:pץ4Cbk�{���5�SK��Pku�u}�f�E��w�!��GS}���Α��h	ŵw:���F�;����f��W���Z��`��G�нKh��׷�-u�I\|8��DR�г-�r���i0E�U���=�T��^��x��=��XJ��!y�(j"WK����%��H��>.�̡mA��=��>�z�7'�v�2wI���uᾨxz��2�`�%�C6|�X�a!2���j�W.�a���'�;�Z��6k��O��<��z%�r�����Z.���"�#���zz��%��z��YK���;��)V!��
;"�-ښ`��LGhc��e'���6ec��D���m��+.MH�͟���9�"�{N��q��i7L���
��V^:���`!A��zwu��'�2�eWQB�5�|�5����ۆ\ߟ��P[�C��ei�<�;��/�{R�d�9[k��M��f)�0wQ��d����y��~:< ��WN��z�K27x��
*�[�Ԫ�ǘ���{lDq�3���5^�bC��gz������T4m�&��A�)N��}�;����.ܖ�>í�=�y�C��w�!�d���R8ɵ���.����/�yٹP�����ۿgkCM�55n�7���wJU����J�e�=�I�٠ �_����{��^�j�-�i`�AfL�����͞�
��^�eU�:&Uu�w&��с�=�v8�{~(ڢ3x�zo��׬���xy�����F���W�.
߁�P�.y�x��+�v�t;l����#C������Ԏ:϶`�Ǣ�	}��pU�Ю�p�k��� Ϣ�{�0�ө�l..�������,����)�.L]D�x:���/ +r�p*4k�'�����V�N�����:f�7�.7�LRj���j�i,����|_dI�%��u���=�Ǟ�Λ�m{Ļ�f���$�#�i<pv﹫�*��J�%�,_
�	�X�-P*�i0aLΣ��,�t��B�ְ��q�*m��̰�����fg�V��4~�K�@@�O�;i�W�`�m�w�;�\�_�Ň�Zf���7���Zo@RX���u�(pU]D
�	=�Q���ٝ�Ļ 	~ٕ/�ag֫A`��r���B�9�z�V2�7���b���c�I��>�R����tCF��Q����4�㖓Qv�͡BtP�rŉ�]J��C2�I��m��b
n�u������&�l"�d���۫VS�iʗsT+r�`%Jk!�{�����`u�ں��zY�l��e&�kn[��=�^V�M�L�J�X:�q�h��0�ýP2��7ykVf�=J��E&�LgΎi��"�n���p!�^�r����kٻ�"aW�������^�sV����W]z��de�ل�A(1��3*�,Q�Z�� P��M����=+}s_T�Xڞ�E�B*�Q��Gd��Z<��tv�����k�;^�5�W��G]G�| �\>�����h�'����&tU{Yo\A���wf螤w��{߷{�i��?$6��]��~�e{�u�lO���x��ѣf������< ϖ�LS����K�U�r~:�R�K���|,Xx�[YS�RU�T-&��N|���s�œx����*nRhʥkD�X}G��}x� j�q�m���d3�U�\#@'r܇SNzz��K�0�����G)���jH�3����3��|OY��)U�`��b��\�[ٱڱu�mʅ�S����V���k�4t�DpU��}��lߦ��^��"�{��8K�������m��;6����3le9�\�K��F��}G�GѼ�L�@���h|���kn`�h��g�N�
���ݾ����F�׎ZK��R�oݭ�eݪ%����Օqu�ʉ
��ݰ�?$�����|uՌ�,3v�������h\��\o��.�(k��hӨ�S�Q�T
����$=媷-<���r4\��<�*��~�D8�,��P��7��h{�ھ�n�5���6���u��s,:#"�O����c|��ܰ_2�^5x�N��#gN޹�0�J���*tx��z��0�:�?�3��R2.L|;�KU��2�re骠w:v�4�tl�x��x$��ܟ\�'�r�[9��0b��>T)[�/�0bc��">%�݊?z�vQkm�q�x
��X]F�
������u�U)|-f�cB�n��=rc;+��Ē�p`�|}CEϞ�+�r�_	|.���]�A}EW��1WJKN,��弭.Z�5;�/�d���K�]eǮa}.���NF/�ʨ�
�G�@ב���elǶ�������ϴ���
���K��V���RȮ�`�@@U�V�s�{zw5fo^")�������p���Vⷩo[�T���h��,��P�y��FP�繳ب���{7;�E���g��D[�D!R�k�Nԣ�RN1G��v*�T�M��!��y�{�(]��`���$�b�����{ٖ�{�v##����c��/�2Űh�]��)C���Wَ̉�5�LP��Ĥkx2�Z��;76���MY���/^�[*�=Q�����WO�E{v��|����[xNu��SS�����▍�ݼ�c�{��i��Z�<�V����߅���\2���Gz�p�L>���gk���g�[��d[ꜟ���h�^��t���5�ׄ�eQE��{V�/z��F�W	�;'E>��)����\��>Q:�쇨m/F�7�G��P>�$8��o48-գ�݌N�$xT����:��'�7+;��]��֪�2A�����8�[�H�h��r�'�d��	W���U]��.�pUo��ފ��j{S�H/�f�Ci۬����½��/���<�B�Jҫ�^u��=B˽��؁e�����1��n3���w���;%	���OA]��+��qdui0�}��E/�YP����;�Vu�f��x%����[�1ힸ{6�J"tK�hL�X.P�;�먝���ޮ'>.�a�oT[�`Vs7�O��\���i�}C4�Qh���,Blz��9z.�ɦ
�V)�aدn<ו�*N�p�>�{ںq�<��̠�
U��L�{"�:�M0	w�>U'�ڧU]���(�
e{����Ba�-�n���-�ɶ"���/���D��j;�Ls�n]��{�\�{+�-��P�B���kkb�?B.��"Z8��x�����ˑ�ޙˁ�s��z�#���¦�Y������!�5ż�*���uc�x�R�>&M<��"��f��V�+���|)�N����>�����b��VK�GJ�|#[@1�'�ܒ�ɸ����ͫj�p��E��5�۪~~9��eچy��2�Xfh%t�uz����r�e�v��8l��őt���{�f�D�Í�+��y�z3��SS�����!���L�X�N�&�=[��RE`���Ǵ�z�������RUG�2den�A��~��b�Vz�smCеx��6��o�m��5�s�8lm�^_d�=[�ޞ}�,p��hJ��PT���}I�ϝ���h��@�g�Ώ0}\���'q��#��y��e;5 ɇo��D���P�_y�Jf�qLb��4z�5���|ɗõ1�5G1��r��d��ޥ0ũ��Ih𞣣>�@V����eq�9P��bO������ޣ��$I�ͷC�02�A}hxkB3��K�2c�k�*u��a�:����Mc��s��p��/���6ϩݲT4�Iu}@�6��X�a�Yr��Sv�U�r��Ȱm�NӁ�$�yy��%!�3,V���m��)9MWb�0��-Ձ�ǄnvN����V5)��vc
e>��͌��<������
��W`�ӱ�4�ح풣K{+Ou�*�sI�⾩�F���'S�$�qٺ��7������!�������];���Q�������f0o����]�>۶�n�<�}a3�l�r��!���)
�
�J)�ЩQ���;,��b�7���mWί���}\�tB���~6���hz��f���_y0��m�d]���#w���0}G�#a�%.TF�5ጺ���Izm��-&��}m	b��;��!�a�>����\���=���O�P� ��f]�"�=g(z=Cl���v|�ײ��wa'���[{W�����AX=Q�%4�)��3.�{N}H�G�JN�1�[�o��^��ef'<��Ax��t@A�* WF/,Q�릜����,�]�c:'�A�yG�j@�>��B������ʺ��[�c!ᤧ U�y��o��Ŋ��fg�U�m��o}��->7�nXƐ�[�I��|=�pN��ᱟM�}P��7S�
�7B��m��ıb|�]�df�+�}Y�3+�i��7�1G7:��n������^���
U���*/�Lu�,�iv���Q �������Ͷ�ՠ���=3Vu�C�[�{���nV��aWf������}����1�����q��O�N)Bn��Z4e^���v�{[z|W������kn���V_Qܗ��b�A�O[M��.w"�ꞛ.j�x�.����F��g�KB-���� =���6ڗ{wю䱻��^�s�8�?_LS��X�:����	���Su-�\%ݫ��οl�ٌY2�y��Q1����2�fYU2��ƩW��N�PUga���1o/]�`�ޚ�����'���UM��pL���]���o�T94�Q�4)��.��)ՅKs[�u�'°u��]�qq,f��3������\�|��ˮR��7(�ʶ��K�ɨe�fP��XlPCޣt� %Q:<Σ\/M��R=�WC�MvKF�V�����̱)���c}�Ww�9K��}���Q�����*Ǿ=l/��ϕ�gz����M�z�W����Qs��]��H_�^�d;�$�%��]�^X�~z��+����P���ލ�S����\�kYV���T�B��^AF�r�>tn����X_.�
R�^iӛ{n��\~���y�5�|ȅq�Q�.�8Ҕ&P��heC�
��]���������$"�2�	׵U��+E�F�# �u�T��._ݮ;��E�nv$ݗ�
T�(�4u����|X���X;8U>[W�]J�7\ڭ�ef�cԥJ�2k��S�yN������,�Il7�W�9=�8�\��sg�m�'q�$�2Sy�����;�g��Wif�L �J��*1~TUN��V�yFɸqoM���4�]N/S�]E��<��ϻ�p��5B�R"�$�޹Y���}&�n��n����F�ua���+��7K��4�)|{J��*{��6��j��2a�$�ծ��{'�,V�K˭??.�P[e�v��z��q�;�*TG?{�f�Ga%;\��x�pt���1�;g��j��i�a�u_�5�,W�ڑp���u��(���s�l��:SyBWu�����K®���M�á���̵^�\}`��D��x�ôY�1�CUoot>��HP��+Թ�?V��D�uqh���4gK�n�R���e�}5�j�"�ϟv�2��v�G,�_6��Q���JS�eu�%B[)<���JܵI������Z���=t]�/�VU��Y��4���{\�@`]/+k�xh��Ei+
]�3ɳ�/�X�c	������P�v��^�^�˧�݆��߻H@�섐�$�����$�rB���$�䄐�$�$�	'���$�䄐�$��	!I��B��D$�	'��$ I8BH@�RB��BH@�xB����$����$�$�	'��$ I?�B��B���PVI��~�� ���` �������ן;�$T�����(HT�H���J(I"�U
�RBEQ��UT" � *�HJ� �����**QU*JR����HJU*UUH�uY��@�UA*	I"�@�R�)V�R(��RJ!i�T��D��LIUH!z�lH
�)R��$D
H�R�F�U 
�U@IT�QPPED�M�Q)! J�%A(��S��
TR���  n��Z�r�:t.���8֪�Q����4�R�sM���v��H������Su��Ɣ]��gmeWs���Gta]�v�k�v�(JI5ӡRJH   W=
����Z�iCsZ�u��vnuU���TN�8[��*�u�]̮�"����&��U�����]].ݭC�s������vB��UUӌPS�IH�JJ%x   #u���B�<�
  ��(]�^��P �(hP���p�P�B�
(YոP� � z���(P�@l�=��P�@@/{E�]C4��ڥѪ�@���VM��P�%$�)J���#�  ��ǡ���k����Wj�PqC�4٩�M�ns�[M�Sc����v����V�ַwuS���ơN��Tݶ�jugv\�gmZ��(n.��V��`��2�ET$P��/   Z.�UZ�.]�N����m͠���*�SW]�l������K�[CZ�%uk���w�
�q�wjr�r��wS�\6�N�v�jlt�M�]�M�s�QR��$��H�D�   ۓ�ws�r۷]ݻt-�Z�]�uMҮUgNn�;�i[�Y.:��U���]��m�Gq�gu�Xj�5ʗS��ֺ"�:;���l�6�79U��mSn*�"*���+�  -^��]iہ��V�ӻ�n+5�W]����uC��F����u۹q�rM�Sl�
�rn�un[9�qͪ��õ�]8֚��wckJ*���D��@%TQK�  �:��ݹCUmƍDƀU��hE�;�wP
��N�W8� (v:���9��u-t흡�Z�P"�()"IIT��  f���J�u�T����lPqI��R���v����ֻ݊�� 6U��X�8(]����A9D��D�RU!�  �<P�j�ֆ�uب��]v�U`�� +��P�Eiά;kfF���(:9�ՠ ��q�@�k�=�*�� hh"��Ĕ���F a�`L4d�)� ��@  S�����a0M�H���E��w�~�>�} ��>�h����^2�.�1��ӑ�#g�UoOQ$g��x{��{��s��~RBB��@�HH�HH@��HH@�`$�	#		��O������0�?�z�pu5R*G�wt�kv�)xr-.)�7��p<)F�Z��MR^�J�Q� r���״DZZe� �mZ����5$�Rdn��FL&�8�Wj�Ÿ%Ia
RT��7d35���p���1�ø5� J���E�H*yv�jB=)]���Xze���f�$�4(�4��b�ej�:�(����9��,PU�bu�j���i�d�13f̥���-��nm�(��d���"��v~o*�e#u{2�kZ����R��76��0;Q0%bb�9����(n�pQmF�u����k�4�[x� ʭ�X3����H�e$ۻT��tK�yrܖ75�
4ޔ��e73���ѱ+,�ܽѦ!jR8$��mh$Ք�0ڊ�-ӗrf����-�-�YX�(�DS��rܺZ�hӹN�I(����TT !�B�3O��q�����̫w�=�e�/^�c!��d��ӫV#�-���9@�6R�ad&E�Lp��;9�FFsm�4��EJ��9d5
5̫w[��*��<T�kɮf���$��.hs$�@ek�Ii8CKM����A��Va�/^J�ֳyK,X��i�JX��2���:�l&�cTdU㣍=��(�m�����r��СF�Y�t倔�D�,���#v>�?�֓�	N�n�J�����ݼ�"U�~q;wYmj@A�wW�Ss3Kc@XLҎ���5U�.<՟�9�Eϛ�gX BC����h4�	����paV�wY�K�����`�M�T����$wF0E��jQ�w�+U�O"ݤN��7�I�4���*��M�ۅ�������u��HX-���� �5-ǫ����o�"I��Nh���DXJ�S��j��V)���pY9bj9��B�vR��I;gd�a͕v����"ɉَ��)�N;��v�āc��t<�]�y6��2��T�Ś+B�Y ��v�X���e�L�[.��vn�Ķ��@��*V^�Z�MLi*H�v
�]@�0���N��D�],�+> ԥ�4����z��KxLY2&V���1����E]��6�B��F��*�M���{����[�KJR�v�C�N�"���JAA�O��`��)]��fd��$n��W��Lă�+aM\�+7n�����Pl����
��	�
M�x�m�h\4���<��]�"'j�@���ׇ.����؈�0'�lQKks�E�50�m[1c/l"��ɸ�;�P
�nSU�nL�>XKU�2-�����hU�g�⵳dd$� �ȶ�:���B��0�v)d��934,)!�X�J��57k��6����V�$u�@
�X�5�\�Ѣ�%��@p�P��hr�z��YCM*���u�k^�.X雅_WCEc��Q(�e^�b�_��2F�Ku���N}��ѳ�k�6��a-�w���#R�2q��%n	Q,7�F�t~2��6�=�nYDeG�b�͉�%d�����Nkm=Q���V�S���Z�2���e/���]�eˣ���H�feֆ�*e�V���MF���ވ6�*���������e�#�(�H��Tx�Yߖӥ�f,���q��C�v����H`3A��t0��ĝ�c
N�K�X��7��ܴ�K0a��B�J���f�Yn��p#(���(m�sum�z��Z�nϤ���I�ݕ.#*k�����j��s⚛�����h��E��{����ct����6ݑ��!I���ǃ��k4l��bƺ\�3���W�4[�Enkn^�&�9MK��R c-<{�ct=D����U���SZ ��z��z�����곴M�C���i����v��j��A�݇
�P"��-z*�׈�.��p"v�]����ȕ꼖��Z�8*-%=�Y��&�Vٲ�-[!�,�߅�e`�-[L��0Z�(�!)����z]�Яth���ͦlK���D�8�7������7����[r��
� �f��V�g�B�f�]7/)�7�ʙ.�4���M�Z��8�����F�ySX%С(f�8�*�Kd
���*f�L֝\F��ܫ2jQ��^�m���!:f-�[sF���흐}c& �RNH�I�9s��S�sV4Yn��U���a�"�7m�ʢ�j��ò��ki���ʻ5�ldQ��݈Pn16+ic�V^���Gji��x��]�y�vL��J��$���2݃�[[���k2-8��n�Ihڐ�R�$B���2C[���S f��n,Y27���wN��q��k��(R�5�vwr����/��O�j`��Y��#�A@�:i�m[jR�J�ݺ����:4Yi��'p2
��-!a	(-�����P!l]^���)��0K8����7�h�]��s4c%�a
%�����,U�ZQ��.G��ݤk/)͖
��;�:nh�V���yR�T2\�Y�Ա��?bj�2�Ejl\�+DW2�	�T�A;ǋlY�`f6��,���D��ފZ�4^<��E*Ab���6	2�3SD?_��n���0��Nĸ�5�`�i����u���Y,������3�D[�r0�XU�3-T�U��VhD��Z!�$ȝ�MB%��n^U�r،�l�lj:���XԆ��b�Pz�/����V��]J��l�h�i�Y$�¶;���1weXA�a�AU�csVǑ;//Y�y��!Ė�bh��*����W���^,�[���RU$�@$�Ҵ�j����U>�B�!g`����P2�l(
��[uf��e/�]�[���qڕ�&`���{MAl�ʻ� �������W���Ĉk�f`�V�-60ŕ0۫lл�	R��f[.�[�=��A���xVHE����#[U�5w=&	h9����k�x7[9�c���H�HJ�'V��U,1F��y����b���Lb��f�'/tom�F�f'Bs�N,�l�F"���(uY�2��Դ��d�AxL�����Q��-7�A�B%e�U���gd�0Mf�*t7q^9QR-GFtP�-��VBr3)` YC(�%��L��Ԉ��f�m� U{���6��ي��w�6@`��ղ�ȱ��P�I�٘V�P�iY�E,ky��b=�oP;�� �Ǉko^\�Y%�GB�ZSkF����Tw���G&�Y�^85�t�VԹ�^�S�P՝�5�E�#S4�j��ZB��=G>�,�3�퇖�y.�W��ɔ�]��k%�M��N�b��v�%[wu*���R#Z�l�tkLt�պ�1X�66��AA)	���x��R�$�L0%Q�u��m52��Sv�+e*�n�Gv� K^�	�����R�W��t	Vh�z(h#3jQg0n��P2�eM#��2�R6��s/s2��F��-�.�� ي����l�� ��E�fu���q]mB�p�fAAb��I%�;��ޫ��ƥ�(���Ǖ&����\�uؚ�Ae�;ͭe]g�\�؁t�t��nVe7����̰`۶��qJi��x��B�rW/+(;�4+�(C�x�#�d�v�^m�.!f
���H�Աl`�65����b�͋v������P�mn�
�	sM�B�Z�2b��0m��N����2�N�H��KU7D�!��M�F�$�Źkf��xI2���!�������y�
��a��d��^h�GvqS�dÂV^���*�liư�f�ɴ S�pܧ�CZ�EG)b����hdڻ6)e<6@ƚ�3���/n�M6�\efUܦ*�$�@�x��I� ꄊE�[W%*B+�z�Z�H�ʘ�1�lY6��e ��t�1��*��C�(��
Fd�S&�����n��VB�k@X̛��0!��(�)���Q�q�-�V���]k�L�Yh��km�p�����v -����q�0�D/��[�{��[e����汖��Q�l�NY�ł�9lCR��T�K.(.�̄J�%n��lS�[[�c�kTզ��i\��+�ڳ��ʘ�&hۍ��<���¦qy���ctsV��n�LyͰ2"�]%OI���E�QK��-ut6�Ci���A�yX,-3w�\L��e�Z�R�(���cR�p���J�s/S�tT�}s�Y��Y�#�I��z�x/l`���Ja�D(b�-����o
P*�fL��V8�fkNaX�E��5r銘3`�z�i*���iJ�Yh=���p)+t��.�1eŃ��EL�B�1�k�J_ۅ:.�˧b,�jG���.�&� ���2�[���3(���Oi�-��O
������R2%�2KfˁL��n�Z\�5e+V�܍F��-<��{�\*���x�������+w{���<�"����\a�d*Y͕v$!^�I�����х"��2^�7��
�Sl�y�[��h��U�թ>0����h^d�́4��KA�1.��J��g�H���d�z�%*��W�U��i���t�*�i���+v��kl �-�XR�Z7Z��-�P�ʺ��R"�F�o6v�OV]З�ܧ�c������M��e��Z4���&S�%�Sz��r�f�cŉ���ջãD6�V��Т��	Ш�%�)�jy�����
z!�jS0낖i͏"���!��bӤyXN�Cٗq�{Gd.�y�dk����iڐ��	�ĬF�e;TwS;/NԻ
S�����L�Р�4*`˘�[�4`a��� �Gd��,�j�i�"ɲ�\�md8���zr� ��m��&����V�܊��B^2˻�-��,�Y��nU��QT��7!Zf��Q�4���l'd��>�`4�(����(�j��u���O���Iy,�#�6dO�u�jguݻ3#�z�h�͔��-j�M�BH�
������!�jC�ab�7 ����!0n�h�b�Լ�2Kze �C��(��Kn�]j5aq�B�n�6��Ak8��ER�2��l���FAn�l��a���1�l��o@p�g::��&��m �R�6�K	��leK���5T�*�Ф���#��4�3�H�G*��Չ�t��WI���f�kl:����e![�r. ��YZ��VZ��7OU��yj�&ӫ�
%��)�0�3[J��Em'���ɮR�H���[�ɳ^���h���yB�\�t�rα �7%)f��c�(�r�<��i<ͦ��Wڥ�1$��o��A��#��^�CB��#16��X�^m�34�6�'��<��A��6�%+��*3��;�*Xn$v9n�<̫-"�^+���� ��Zr�A��2�E-��]	��'y�;�C��gVt+I��j��Xu:�SI�э^�Kwr��	�73w#��T4��f�mn�J�x�-��G4�E0�N�ԵC�4��F�=y�v��W�l1{���ժ�9�[�+i3sn��%�/"@,�b���/%f؆dّ�+]ؘ��ܴ�M�����ƆR�5�>�1g*��bt�|���*��녲�c�e^�6�a�ɓA��;4n3<�jhH��G!���ŝ��,m�P�Ys�Dȱ]X%�u`�%��"��{I;�����CM�d�#y�	��9�x����̉3�T��!%+ɔm�[vŰ�!A��,��A]�D��rVS�2V&PLc%�,k�y�f<�A�V��W5¡�.� Vo�5�I'�6I[ct����TRl�0��8I�^m:J��WuIaֹ[zKnm�5��Z�4jg�½U���U�c,�4��DF�*��f+Dt\�1W,Z*1 (��\�5�q���I36J��*�֭�T��i���2I>�nP�h��]FrɊ�\�Jh�k�(��h�Q-0�;�V�D�HQ�Z�b�uuA㧪�nX��IWw7/�Mx��V��W��ef�-��i]���d�P����ڡzf#5d��S-ۃ+i�M!z�8��Ax�X���P�jz���`+Q�`�TN�)WYB��/tࡶZv^��N���Y�Y�]�X�����˖N
)ø���+1���w���k(���8��q`�������W�E�F9b��v��7��6i!��W*V�ve�����56
:�[30f^u�[�ek��ll�fԹN²���d�m�v�T�����'-��)f��d�2ˋu=wM�0U���G*RU�%,��r���&*ۣ��55���T�`ve����g5�FKʽpƄhC(���0V	�)�km�Z���Dk��4&��-�i��:�h�i)���$!��B��P^P��K��P��RH�X�P�R՚U�
l���x�`�a��n#��9����!N�녣t!��Z,��Tu`�a9�4�Q�T��U�H�� �EdAe�n9B�̫5�E�tA+
h�2В��fּ��Ց�#E�i���̶�2�L�Si�2U�:�-V��@��F�of��y�lk"��nl��m�4ڻ��mФ��Z�/NlF9��K�P!�E@h5m��h�<��D��2�l� ;�ɧE�b�z����^<���p�h�x�bR�k��NH�ڗS�E]��Q��D2)�ƭ��VH{�!)�����^�k����Y�J��VFIs^ݼp[��wl��d�4��Wqmn)���b�t(ؓ�ƌ�6ؚ�Fih2P�!=�GSs]�?!P���d���m˒1D����N �2�k(\t0g�r���hb9*�J�Q�]5D /b��S,7-�h�u��fY�H0E�#'�m�oQ1��u#�؉�rN�o��1�)um�2�:k.E�m����2N�ۛ��
o�ڮt�C1Vu��S��mK��s^�Bq���uZ75o]��g���JVU�I�b��V��\&Bp�Tg9�|��[֧p�:��}$�;���qfVX�Wv{M���٭�-M���'7l .gY���l5y{:--��ڊ�A���6M���9�<*�{yN�	�Ңº�v���ʰċ��W1_�M*̝˨���}1%��6�6��gh4
{�#�l�:l./�����Ba�A#���f��.y�ٕ���k��_����^&�:w'_]a��-:!J�67r�$�D<�݌��^@���%X������}+�P[�{�Kͼ=�3�\���Γu��f^^��J�Te#��;
�]u����ڱPIL��gw+�|\7�c`���s{�Z�Ն��BN����сV���,}�eF~�C.p�D����5�X����|�M���t���z7��}YG"���~+
�{R�:J���k�ǩVMwϦdL�[�Hӑ��9�#�1	;����N%;������,��(9ԪtO@���,���]�n2+�x�'K��4x*���}��;�D'��!aWl�Me�Yq3�5S�r%d������+���(�c��R)O��b��G�u���޹�	�����\%	5g��\�I9��t�l},�[/��������vF@�8��Ӹ):aNavkwe�7�I��l�kƕg;��z���#}ܨ��im>�W��ѕ�Oi�B^�[C!U;pty��֥p�
�5���O)HvPuc��xǡ'w��k����8!<��S���h�a�s�r��F�e���dT���/��n�V�p��F�n�Ǧ��[��p�ٸE�p+ݑ-6d5,Z�G��r'��8��y���.[�2�2�+�����
��#gu]m����$HiM�.�"=G���ͫWT{eT�i�V^͙�K��aCg�5�I/o���̊��cNCg�f[�jFc��M(oBy�,fe���m��[Tn8z)v5�u��gY��^5A�l�5�g��esFL�� WB�e�a��{
���9���h�]ب�a�|9��l��gK ;���fY�nm�l��1c���JR��p�2�P����.����cǙ�@�ٙ��W�2N�;6R���.-=�ME���u���N�`jgY�g0�������V��o�j���9�u�u��\���&oH-.�3��̦49�f�T���6_g�v�)�|�-��ԋv��Oj�1���E��0!6��ĺ-C�R��$�\#*8���9�[��:����]ۂ�g3u����U�V�;zʏ�2���9����j(�P�ȂRP�Zn��]8�D�ˡ�L�3O1e�j�S+���f�j��0q�ۤ�S�J�L������'��5%oq���DnS����`v�KW#c��<��C������tX�f�\�)�+g���z�l��"�˱_K_MJun��[�.�������;*ޓ��!؜Ìp�r��c�D=E����K���8���S��7h�
�3��c����gӻA�͂�^8��ީJ�oٚd�,�ݸ��ͤ��#�\��t��'��FP�6q1vCޒ8��ʻ*Z��*�vVr�3��z�S�O��]��޴���h�����f���	N�V���u8"�	B���2������7����襺)��u{�%��kbW/�����=����$�HT����2�<·�hN�Y��إKN����6���vU�$0���ƖK�Ǔ����x*�Tq�H|�]n5z7�6Y���6s|��N�6�k��'jfV�C-�w�\�'ۏly��8�*b���?c+���u����vy�1֜_���q�g��=��d5r��ȭ���O w�y�nu<��s�˝[����b��L�6Q�˪Iq�2�WR�E�*�7XWe�[�,`��k���*�ڵ�����X�!ڇ����x���ZX�<��㮏�j�t']���ć�=���iM��՗��X��9��c��\&��f`D�0�쮚�=b��M��FwrE�<�3�c��)]��`Yj��LW|Qug�W+/r<�#FR2�l��;oX{���(��[T[;t����kwٔ�|]e.�#"w��HrJ���mc�&��R��y�i�n�$��K+���ʖ�<�צv"�|�u	N�c�oM#W�6-��w�CV�*XM>�}�ubglY|=J��S�#`M���)N�M�ۛ�$�p�N���"C_QրiWGȎ�}���Y[��%J��ɾ��T�}�i<Eߣ��/j��#���cTh��4��3I�����*��[���o�n*h���9����ʴ�7^*g&6&oM�ڵ���D����%#L�Y`?�+[������^�}]e���hU�U�0����F��V&z�c%����铛�t{6]�S*c}\�T��F��a��r�gjˀ����k���	�`�����1�k{F*{�V��}�1���H7Z5"�gݮ��v�Wl�KF�T�3\�%�J�3"��듑GG����Vevq}���7&Z]/����Z7�o.�]X�Sl�t~�.Xgj�f�J^���5 Z������WS�J]��V�"�A����T�z٩�릪r��$�V^>�����j�M��]�֤�v�-�W�u+;VJL�������$Ƨ�텙�a�tI�H���3z��z��y@k�1�K;&jG�mAf�Ё�x�*�R�J%��I�bV��Dbl�pH���b�$:Q�d�g1�
�[�2�;A��U����`-�5k��@9�c���3y�Z��J�G�R�]�����m�C9eY� bZ�7��sW�=>*����]c��֝�$��R�'ך��Rr�t�rW�T9k�܁X�Pڠeo9nJ��o;Q���ؙ��A�s\d��7���n�d��  AW��ej�p��(�-X��pp
��ڊ��;.��Ԑ�+6��]G:vr6.� ����F�T�B���ZA�_2���+95Nv�'k���a����ݩZ�n�6j��ʾ�wi�B����.�qg�40��k��'ݕ��΂p���Ӎ:��Uʖ��.֞#��O� q
��j��fv�������'X��Dɮ�vi�5.��7E���P�B�Q���h�N�����@7��e�<;7f��[�ozq*V���.�2��K#W�}f��L�������9�fJ��;N�褸9-�y�����r�	ڽ�����Ƣ��ԙ��S��׶zU�]ז۾A��d�#�R>cU���ʟm+�2��<�\������}L���KB0�5Mܼ�+G�OV���elf]�[Bsd��A�ݰ54���a0�����6�n�s�k�Ji�3�oE�j�Ū��t�P�����c;����\�9��I����as[��H40OY��B�":L��	���2���Ռ��7$j\�g6�	8�q@����-��gJ;�]�E�ZW	֩W��Wt�n��9��:A56�9:��y(�޳�.��b	���K*`��q={�XF�G%2���,�[hQL����4E��M�,l;F�;+���;͹��Fq�����9� N�,�/_�w������Q���) p���#m����$.�[��9*Lj�uh��kLe���K�:f�#�������:��8<[&Ɨǻ�C�!.yx�������g� X�.��#�����VI}[C�s&��ݜ��ҩ��8wx3v�^f�)y���g�9�}ݥ7�k�	B�3P�rP,sx|^ev���C�N�9�K����4We+�	��-B��ӗ؁���rȯD0�H��b��tw)�M���t�>���Ő.�7xŕHa�:��i��U.|�{/hhz3#�$�J�@���]�s%V�7������9��m�Q�-�$n��]�-UHv���Y9t���z_tճ�����s�$Iʤ�U�}��ru�f�qmdX�Y>�'s�`FvA-ٷv(��7'r*��-�T��mAW�L9a�CAF�+w��r��k�Ypq-�Xv��C����s�m����մ�YQ�P]oe�����ǁ��:��Ű��o�u\���T��q��_5y���V�w�еÍt{�v�v�-���,6^ƀ�Mlj2���(����M��%�}�.�
y48-��\#����cx�A%a��u�֟��%�����
�F��DZE袪X�ν�p��F�@͋4VN��>���u$<���,{��2��Agz#+�O1^��L�@�ՎiTz@}#t���uEJ]ޠ�u>=°v�N̢w/�`j;.>3�4�ս|�9w��t�8���dJ���Bi{���빣��EQѫG~]�oR��L7�C�i_/�4�&��=;�R�4��n0�p�v��Mf�݋�Ps�2�V+WC�&��@�Hy*Y�u1c���%�<�(s"�7�c+�ϳ����K(�p����{s�)-�3���L�afviU�Xn���BA�V�_<Q�/���g
�2��(k�L�҈�w)�8����U��°�v⫉�9����p[�ȕ�E���P�Z���ѧHkL�"S��o^��F�[AY����Y\р�����ENͺh�� ���N�����a!�V�ܚ�v�ofX�* �0�=#7؆n�qB�����v�L�vE8O-W�{a�-ES,�mQ%LV���^Y���(?7	�,tCV�1��j,�p�e]��q��c���a�$7�{�o7+6���&_�Z� >�5|%�H��ɻ�Al����jL�v:�G&嚨�>v�R��s�1W|��.�aY�N
�K��]�B�c��n�å��y���R�ʶh����kiN[`��{�
�f�vٻ�,���#y0�a��c�Ԯ̔lj=��O)8~:I���\y����u`�oO;�Saa�}{�EEe![������8��v�n�w�d��'820�jH�i�����.����y�5���[������j=���<�S�](��	��e�Cε ���"v���O:�.��h��@��a�wL�S-Aٴ���A<R=}�a�B�us�*�Ǣ�H&�6�G�n]�.֠���T����У��Z�c�
�U��l��:7�^���v��G�,�Z��Ӭ��U2Äl�X�M����ˮ#(S��:�U�Ď��#}E�}iުiح��.jٹ�T�6�kj��yV��J�/����f' F�Z��[�ն�qB���Х��`w�!�!�Зv��+^��bͱ�ܫ���Y��)�ȶ��"-ǝ������2�V�GuH�����]^R/ת��|��v����V�5��zo�T�p�?�*�'9����M����юV���c(��"��;Tqu7��S�-$�ԒxRf��eʖ�Ά�°HP���]�
�7��'Y�~�2�R���,�����fV�Spt�P�G�r��}��Z�'¯y�r��>32t|V.��]/����Ddޚ�'k��:î��z��"�ʇ2�q�;�`\6���U�Rf;gH{xu�ֻ�k��[�dMֆ�v;�/{/]������
��>��*Vt��X��z!�1>��MV���T%�pN[���Vjt� �+��y��Ps�+{�f��S֙޷L�)e�Ұ�Z��b�a{�@�N��4z��܂v	���G�N�zv�I,�%@'[e�gt��dD�� 3oe�Λ\Cd����YG��3�r$ո�3|����C��k����U�cn��[{Z~u4��U�E.�u�%�.Ӵm�t&�t��fKcdޠ�r�A�!�t���#�@�,ܚ��N�V�d�vjwH�����@���pa���9�.皎s�,�;|�O8���u����:�p"��;N�i���b+;�hsfaU.�9<�}x�(�u{�t�r�:���*t��,{Gߧm,�H�4v��	�;F��&"�����=����p���*W�����H�)���ͳi�R���s��ϻu�s0.}2�b�׬����&iZJ,Y}XR�sd�ފ�Ўݒ����V�w�J�����Wk\�,��k�9���x3+D���)ٗm��pd����:^3�Ү�t�cW�+�u�U���vGl{%��l����D����u�y�f�&�oPۋ�'f�ݧK���}׀�*��2�rCt&d}C��tk�6%]���-��68�j����n��Q�}|�m�/10�7�K���ls{�^<�k.\�t���:��',tB��HՔޅ\`���6���*�t+��u�yݘ���-���u�X螨V�wOY.]AϞQVMue�7h�oS�b9iֹcm���Z"͠�n-�*V��}}�:�J�혡�29���' M۵���w�)>B�z��ڡ����󲁸k�X]%��3�tƴus���+�%�R=/rSJ�5�O�FJʃ�
�Obߺ�cg���DoBg"���w�>ƹ
u	��)�e�b�ֶ��*hk}��>g��f^-�ŕy�Z���z�r��%Τd���9�%M��{:��Z;m�5|WKV���7��;�I�E��i�7��(�ʷ[�c(�!��ݧ��ev��<F�[Eӝd�C����wK�U�&�eK���e��[؝w���w �V��!�默m�k_c��S6G���v���^�JK�3*�mղU�V-Q9{�p��B���g-���it�����uZ#+(��XKe�ʨf����������~����� @$$?�������~fx[Q}��E�x��Yn/�-+Zr��2�V�J�:�{/ohp�56r�{��5�4\�yp劋u��vz5��{V�*J��ʛ�$�c�+Һﺕ6��#S�8�`Py>��*��=�"�YݣwW;v�	��@ְs���)[a�KaĒ�N7�|���m�Z1鷕�z����͝=t%K��C��,S��w�����v�u
�R���Q]�������p�.�k��B�Z�*��|a���ٵ���i��y�M/�����Ŷ �-���`]����:�I�<h�c��1VI�YsVVT�Sf�k,�K�(Ţm�Zҙ�ź���g�Yep=��i֋�@�Ƴ.$#�SZ�Ցգj����|kS�T�Mt9[�!��Y�u�bmC�@yXA�:ܭ�ֲrWa\r��B!j����U��Y�t
j�ZDR��l�	�Un������Dք.���F��Q-(*����X!wa.��֭���:���˔]��+�ȕb�i��պH�.6E��fn(�9϶�l�d��_S�F��.qh+p-�7���S�P�gd�L<N;N������������EY��
�p��Z5��
��%�NɄ�{G���B�T�ާ"DY�#�V���7k�}*��J�%�;}��f;���2خ-==���w1
݉!a���<Vv.eы 'Yq�8;�'V��kUuZ�h� ��Ҭ
 ��L�Y�w�aea�y-:f�j��;n��]F�k��K;�/g�76��d�v*И��U�EjV��ng0$��o��:��ƀ�8���������ԛ.����(�%�M�έ��Y:MG�hmF�]̧Hul�C�n.�_^V��K;R�����[V��[�U�}%�`��]��H�#�z�Q��a#m�5	ier۴C$���e��R)e���k��u�Jėd��9�Eo;�'plvA��DyK�@�kH�T.s�K����)��f�qa=��9dd�:���C)����7CS�,�B7,H��:=dY�"��a�C�ܺ�]�L�3M�ѵ����.��b��"V��PX����K9��S�8�����gm�\KkNJ��-Kk�٤�Sz��iU��ܙǩM���I�w{w��K�X�(,k��Y��%�
��=-��ú#�R�K&7�&��dX\-�=ǕӟY�`Q�n)L�Y���+���tw�Q�n��YA�37/E�nvJ���E7�M�]��I�-�Κ�C,�юF�S����"�p�O�^Q�\E�,a��{�kX$T3t���A̮�&�C��j�hV�s(﨑R��j�KŅ!��j��>nw2#OXե�H�=b�Mm�{Qu��!hJ����cp-��]��}:��rι��u6���ͦ��2��:�����6�qȚ4��%�.�B�.��+39O�9��&�R���+n�ஓaV��:�҈�^vL�-s�s�miB
��1�Pv ��E�
�Zr7P�%�f,�����i�B,g	m�8���@����)QE�}���k?&��4�vWf*��S���sѪ�"��\�#�.���	d;�&�h�Ү&��U�-��ZZrpd>7M�Y(u�R��r�6�d�P�\C��EB�U�V��eg�Sx���=a�B��S{��s��g`��ހtOJjͣܦ�P=4]��Yt��S'u�C��8��\�kS�5S�� �6Κ]]���	���mh}˯XD,#N*!��p" ��%�����.���9Q��}gO\5�{ȅ�ќ�^(�}�bw;w�����W�6�)U�3i��YE���λ�Ys�m[/��_nwK�EK�}��b.�6�;�	u�������JӇ��s#C�:XR����Kz����9���R�MwS�{�����}�`�ɛk�۩V.��v����7�>7�q@қ��z��V�k�5]kW����	���+ ��c�r���n+];󯶹esCa%r��+��!�ACJ�٥B�Fl��.6�����@^�I����v�-V�Ϯ�dME��۾����������w���d	&7a�nt�b0������5�İm#�QGda�7���wL3�F#X�b�@���ñ	6
ܰ����ۃ6� �������,�\q]��H+�b�̤����Xv�Ω#<4gV�s;��VK��f��n'AqZ7-Qie��Ѯ�GgV�}v"o[{
���uj�R��a�P�Z��2�Fl`<�����S��H�u�a�"�b�i)�㣆��3-wf4�WL�W�ef��<Z���Ut���wZ(�#Tq���v��z��̒��h���I���V�]��e0�[�D���gyݒ�-�j�<��@3iJ���(f�〫���+��nM��H!���-�]9����5�����ů�Iȯ��W#���s!��������sQ;]�T��jr�|�;
�K�s�.��]V��Z��T��y��Aa�x+/��������q[��^J�^NT@�m5͕�̢4\��*r<�yY��-;���F�>�'����U�Ŗ.dY6̾�D�b�$`j�U���I)�B�'v�L���OJ"�wl�^��Èq7 �r�9{xYb�wc�k��a��x�g�vuǯ����R�,�l����WH�u���S6Z[��X��n�8�Ɇ�k6r�]kj.n��-:6�n5��Tx'7�`L��F��g�(��Y�t|��V���og�Q�T��+�*��j���^���G*��b��3WX�]7��P�j9o���ژ]�p����ZU�|�m����+G�>����v�FYa��{ab������erЩܥɾ�i�K7]�ل��y���&о[\:�c�˶��4脸Ʒ`ڀ��$�")�v2�-v���y�y��V�,Y��-N�v�ӭ�ݮ��y�v�82�ʓ���!���n���㮐�7�ݩ�W���V���'�m!D�8B"k.㕽����y�D��M�oszS�$��Y�g*x��S����WVU��f��։���+yb���:Y�;y!��q�y/;�_':�S �Y���4��0.�Ɨ<�����j[���b�؈��Cu�'B#c��b�,�N��!�cO皏wp��(�)o���l=	��QQ嚛̻r��K��x`�!�L��F��rgB3MS�����y���r���gf��(��i�>��q�K�G�z���PYb%l�p6���
ˊ���'!�öK��c�P�ح5z{o5T/3�ό� ��%�k�{,�ثXD�Tyz@�-�'M����^]qjL���ip�nV![�V�B.�\���^2E6���Ko�&5u3��;���f�f����.�N���pP�B�=��cNp��/](�ˁ9�$���p�]l����emv��;n]f�CT�:r�QW6y�;S�^�6-�Y������S��ov�2�M���h+)�hn���.a��k8Z\���Y��tǳ�K� fW�6�<��ɨ���-uɠM������n�/v�J�m��pe�������.��h4v�	��r��9�B�C�Ǖ���������u��ls:��C��V�]R��.��ݷY�=Pˋ�#+T��:R��f>��̤�m+�s#�YU����Q�-��+�Cq��D.�����i�B��ι}z�\y�[���� ����6vd}ֵ]���F�ѱ��Egs�Ҁ���*��/���7Y�A�!ĞW$��G^��*� ��ed���]7�]��{V�a�6�.h��6DUY���1w����儥Y�nfv>����WЅ�'Zq�ZvJ����F욹,�B�t�:�u�#9;k�N���[�K��C�V�)^�]x��c<���q��-ʁ-zk�R|:��u���t��;�Ƨ�Il���-`)vue_�f��,�ӛZa8��o)KqJo��Kfµ͹�UQ�s:m�ܚ����7�.�pu�X���A֌˲�'"�;VS�*���X�9ϝv�-q���U���I�f�T+:�;]ǅ�R��sf� ��ab
�X����3�a�7�՚ǤB���i�N����A��e�y���W�I�tus�ٷ���� ����&I-,��ͻ--��g��aݛ�t���'�&ά��{���FaS�I��X�]c�Ps�]v���VvI�O)b�X��((cݵ�����N)6#���3@\V�&�6��
�E�D�_�����D�DL�U::sLo3��ɵR�g=g�ц��ـi�����9��2,���c"�eH���M9�K���6�vؾ�|��De>�G��T"r�w�����7�NK���3���=/\ҍ#�ա����!�v��hO���m�s5ƀ���V㺺Δ��� \��zU��ɨ���)u�LS2����(���&2:�.��@��~��Md�A���-�]���ʹ��携�|���U��b�Y�d¨�KN����:B(6�U)H)��+��z�:��J��	����H�wl�����&��ή�����h �T�5)f`�R�npB��5p35�us���2��F��5g�t,��z͹A̋�ձ�Nܵ�Tޕgv��v��f�];�T��Aݝ,t���޷]��hr�[��w�g55��O6���]q�[Gc�zӈ�t)y&8a3)E��B@*[�S�!�T�����@�̙x+��'s�X����D���Z�U��"���B۫�z��U������\L�zS�o7{iě�c'u�c		��;s�����a�V�\����q�U�!!��oV�Y��W;�*>	����.ӚԘ.�A�<ֶ:��7���D�g*�
���3[2GW���ky/&fS7Ɩ�\��:�$��g1^�L�l�M�����U%X�xtQ)�q�9����Σƙ2ޅC�u
Ѧ5*+���°�ݚش��˗Y���`�X��:>�����i:�;�];a�.��]�S���kJi��d�K>�|2�r�<�]-�eb�O4�ԕ�R��=Xk#_����J�J��c��2�G$+&�fW6��=5��ϖ[�R�rgg:�\{շ��?���Ы�F�3E8ax�N^ܒ,��p{�{1�{����T���8EG��pI�@L���SJ����R�`tK�e--����A���v5��&�tE�>lf���B��G!�W*m�e�7"�Y/��/�m��웺��7N�Ɉ��R�	�f���1�
=��#��/HF�]BtPh�D��
�o��=D��T���e^��][�{u#�%����˪gZ���u�7Ǽ��=�_]L��n�)j�y�6dXuLq�s�Ū��Y �j��1�e�@L.�7�l��W]F��b�}V܋{V�����ɽ�Ӵ��"����q�;;�dB��ve^	S��c�c���^F����/���u0�:*�rm��N	{M���_M�W��v��)�^�U�u��E+�śQ�J��91N��9�	����.�J�P����7�����F�TF�:@�m(�X�����1Ln��h<����zW��Wav(.ͥW}2u�X���#QAWHa��e�*����8E�}h�Y�'F�+5�@s$�6u�Fb]�2�ɽ��88���E�>h32�ͳ�S�|y�9��5Հ�-���w�<0BP�;_)����b����׍��Q�.S��V���7{��Kmi�n[�.��͓���-�vQʾG;����%��Y�<�|��-�w��|#��E�2��Uso̙D�\f�%#nѿ�/�+��7r��0�Jo؝r:�ټ�<Z��	
��$d}
�N<�nB�%�p�H�m�I����;XmuNޮ꧚��$F�u�6��N#&gG����S�9X6�J�v,:�YNk��
/�7z�U&W]jr��՘>��R�=qûXh1]��ǒ����앦��F��eUK�e'��&��s-rܰm�2o ��q��n�c�D4��#J6��{�r�gs�ji������ȇ˹�v@ݬA_W]�E
�A�UU�
�o;C�O{�*���=ӴᲬ�[+�9���8��R�-�տ��4��) x2�A�7�)9Ի.�i2�;L	�����P����A����3��*b�"w��|�Z�X��pu��j�?m�򧺪U��(��G����6�̨�Hi�;��8-묏4�B�e�%�O�Q��-�3�>Ǚ���Hsr�A�.:6�Z|qQ�@��ݹS�f֊�7�D�GX�8�b@���"�mHy��	�wb�a�B���Zٗ��,�VJ�5'����É`':��>}n��sJ�=�U���WIJ�SWV�p�+��YR�<Փ!��Kƹ]�l�=e��έ/���:�N���s����-
�o"�״´+/���h��.�*ʚ�6�}.��c,�q#�VZ��j�D؊��D��	�C�Ơ/7�	x��s����:�ݫy;�R,%��oZ���E��>.�6��+�z�[gqC��Q�dn��i=j�ud��}&�x*��&�
�׬Ӥ��˻��B�$X�����������=-��M�\]��n�V�7(j*Vu�/���a����w�^���;C7�fР�geEh3�.�%V��u%��-*��a�Uuo�R�u��&���3�;�&ˊ�ʻD�]��w(ns�H�X+����zy����g@h�X�=L��I�J��6��C�Gk�SzԱ�'�ۮ5��O*��j�����/V�0q�(wVƮ�U�����\k@��Y��nR7� ۳Jg�4��&���5��+��'({��7&�����%�;��x{��{���M,��g�ʎ��+r���ۢ&0+�yW-JGh>3���mm�y��Z��<����pa�_s�'y���;�Ә�4Q����*U�x�-v�e 2��&`�%����R���=o-��wG�E��G:�z��V.
���9Aۄ�L�sq����,o�>���J�N\���n�v+�Q���@�3jB*vYg�%\6��*Ռ22����s9�z������u���낵Yp:�s��ŶI�v�t��8|�q�W��iŋJ�y�v�J	owtp'�ɽ)g��fĬ4OwsCMVf�n��^=	��xŢmۼ+����b��,̝�^<�g)0��w��T�(����\�|�Y]��Ѷ��Haĺ�Fu��p�i�r��V�*f⇉Ω2K)��a��/{�0��{�{*"�+u��\���
7�R�k���lZ� ��̸ƚo�N��O/��٩�Y�)^rɔy���U�ź���%��鮾�/�%LM�hɭr����SB�U�f���7.��o
j���v�$���X����,�2fvp���ā
���y�u��D��g�n��k"4>�X��ܖ�qD	t��_K�����8R	2e��z3�yKZ=���e�,�k�����۬��v�Bذ�ɴa���W����s�P#�OMqc;v ��Hut�:PJ�#�R��N���a�gZ�F��V�Xk5��w_(��̣[h`����>vI��h`���dh���F�0>%N��>|68^����p]���&�:��~�s�w��y���"��
��ֲ��-E�QjT�-mJ����Z4�TF,hҪ,���Ң[Z�ت+�B����+P��-�-���aR�Q*-�-�J�*�T��(�m��"����+k,��*�[mKH�Ū����e֔ID���l�Р��b�Ej�����k*�J�YQj* �,��mAJ�*�-TR,�E��j�TV��Fւ������*[jV-V�KjF1b��-��ZʁRV
���BƊ�ʕX����- �ʖҢ��E�T+("�"ʕ�(�������QTkE��Z�+QAh�e��Ъ��l��-�Z��E��h��
�����mA�)mR�ҕ�+X[H�*�TXT���YU���Z��
KJ�+K-A��(�X�QUB�������ثQb�F[me����)(�"	Ix�_��gz�f�-�a_w69��u�Wc�rُn���f�l\b=[�"���o��8�p�ZW*�bk�/��ESz�r�C�M��N�ĝ�s��kA��I�ufSٙcr�yr�S4%�6�K���Fܩ1ۊӕ.��k�2�$[;�gN��5Xݯ6�od,X#>��\��c�=�35�i���Tҿ�j�-r>��4����z��P�x�[�-��[�ƽt�&��x��Hc�4�D�Α׻e�MP���%kE�-U�'�o^%���:�xe��]��~E��1CI�.��f�Kc�F��k7[���D��~D �!P1��g&�x��R*h�V�r��W�Ҟ[j��E߃��d#{LN�ϖV�5.��w1r�����@�hWUϋu�5O:ldg9�`��`uj"W\�βr�֢�.�K�cһ�݋�*k�W<�S�sY��\T�ʺi+|�c�zzc\.�KU�J���Tl�a��Ȼ�v��2x8�.q�i��`�@�؝���7�(�9��D�g��k/0׭1�EE�
�2���&�lk�]k�c|<���^�v�������������\M-ṈgTr��}A�A�5�X
�M{iF���V��ɒ��4^&^�Ӆ�i�YϷ�u����%ἲ����ڇ����B�{F!���j�ч[�<����M�<.�X��McHY{9f!�B��Y�k.���|nk_o
�v�^h��@R����ԫr�w+�n�ؾ��-GKxæ�ۙ����4��F�D���H[ɽ���J�0{Mt3U�
�1�#k����ۻ��n�ޝ�br�8�)=��:}��.V�������M^s�)��5���E�g0ѹZ���|�
[���A!���ˣ�|}N1��M]���l4��n:g�ޫx�g'�����4�>Ɔw7nJ�
8rݡ�KMs*��!:ȼy���T3;V�6��%��Ӿ�~s��)՚r�A��y�"Np�cQ��Pn�/u;����t}Ox�z0<~\eJ�m=WL�b�T{�Zњ��/%���kx���@�W�u]��T33����q���wed�Tk��h�=5qFۮ�V+i"��u��k�<���ؙ��)��;W4g��U]e���g1:rے��䊕�Tʉ�1��&�i��K��ù}'.��h�{v�-�������Y���n�����Q��;�<���.7ixןmL��t3�'٪w���
�B�YSrCU,M��ܲ��H69c�3�q���Qm�lj�x�mtf�ft�����evԡWf��t�Lj:��J��"�ȉ�Z��_�]�Aa�xWL-��|�{��KS�%� o[FG�ڇө��8�����8b��b���K�ի\�
�Nv�8v�S�̇۔���jƻ�wn�/N�{~)	M����d�}�D��f�z��˧�/j�����o������˭�[�^�А�&��y�'U� ŽF2V���Z�i\t<����
Ӆ��O���o	��s���A0yAZ.#FR{b����R.�Mj�]���q�W�r��0����z�&���㳎�E��j���JJ4�0:�"ys��AM��2V�Sh�"�.�P�W�Q+��e��_����Z3����1�jc��Mܰ�d0-���q}*<�ʐ7S�]���7���k)ӹ�!/�2ȱ�K�9�V\���9]�O�o��7n�X(f�Ũ�����Ku�}�8.>�ӎB�Y$��)V�};]�>ܾmXisR.�����K�]>�tȰY�N��C���ë���J���u쪄LIx[��l�)�n��i�w��S&Jf.��a�n��5e{��U"kf�,���a�[ݩN(�y4Ǆl�9�2vZ�6 ^�U��9\Xb���=�j�ݞ$�t�Mk�[5��Zuʯp�����c�"1sL�5�^ز"�}B�SR!q�>YͥQ��nL����Vz��)������'���L9G��*J��Z�22FMZf4�i��]���՗}�������Z��A8T�y8�WPn�H�rǸ��b�#%3��l�l���γ��[��o�$��Ő�lf�ej�n9Ɂ��'��R���L(n$�#�md�t�2}YY{��k]��L�7O%g����pP;t�Q�εөa�(�[w�B/Á��`��a����ر:�0� ��P���qf`S�`ϲQM��Qɛ/ϻ��Y[O��ʄ﹭�4SA��My��,\���/�0��Ɂ�����#�y1��U޵v�Q�f�S�\��V=�0i+־�Q������{�u��$6i����"-����b�HR�a��������/7��Hoϛ0q�3��M[���b�<�y.�yl�᷊��sY�t��溳��WI���k���p�cO1���^�;-�{�1��gE,9��#'��#f9�	S�p<+���/�� ��qc=p���z��]H}hV_�s
9�lt	a~,xR�j�6�ш��-�ļo�,�^��P���4�/Ҩ�b���u�^�ʠ��	�] ׅ����X�ݼ�ު[@����TEz�1'٦�(B�蠺)���Pp��1�K<7�Po���N#�}�ʟ�}�;�~�(k��4�;�Un�TZekR��a}�9�!��i�x�B�A��/U���Ta �a�w���Q�,�����NȲ�ظɎRyi�)c( �@B`fvj
PT��*�_)�81h�ʮf�L0�:կ�YJ�ϙz|'ɪ:]g*o<끋�7O���)f�:�����~�F��%kv�m#ʼ�4��eO��]^����"�����n��[�׋ZQ��~���"�ml�Nv} 7s��V$�J�G���@"�fcF3]�-�A��[�o��R��_��q��W�>��M�A��S�Z���D6�.ĚLc=wh���s"��48v5Rb�¥��Fr���I���r�g�ZB�b��E��
�7�0.����@�x���Q9+��L�wj�\����.���KI��Ԋ���5���<�<��H'�����]��o��u�y��}��)X�XR���R|;���:�t�r6>Zj���,Z�e�����ކ-�Ljf�1�qZ�>�:[˳�S't��,�I��׃MX�]*�u��\�ߊ�Gy� <�u�yV�Fp�Lk�˃��M��ĕ������
sp,AF,�`���PnО�YnJ^�Bt�Q�]C��"�L�^��s�(/��Ld��ur�,4l{�^N�q��;�N�է)�iG/�1�t�k�MX}r]���(Z@%d��a��Vݾ({����+3Y�o���6p8u�C�qp�ق��G�pڹ*��j�W��Fg_�{���ބ[�#����Ǉ�����!�삳�k���[��l�w���ߚ:=���13�4M���N�S��K�S���V|	`�lWե�C��9���G��f���ްc�����035wv��5[�����%����:_��uk��Ҩ����V}ʄ)w5o�.�]����<56ON�Lb�(��T��� �רwb��/��(�P�=rOy�xg�/���Z�wp��n�7ɹ|놎in����/E���tC���2�Y���Yۙ��EKX�**�P�q�X-<���y��qb����lZp$�؝(��T�7�O�r�뒱�D'c-J�@��3$�q�L�S*��ޣͅ$KFGúh�����>�/�Ogؚ;S����+�T��(X����jU����ip!)�����on��'��W��o��uKN�����4-��^�)�������c9}G�oo���fF�@��*Ǫ�s/M`�V��;}��9q�bV����q�7I����mr}פ���|���vRZڴ;��
}1'��yTH�_W��yaf̀�:�ݖ�Ⰵ�ц!Uu���w΢�\n)]�"z���J(���J��@x�gՔ
�Ϗ���n:h��Bη ��!IT�m"6�}�;�V:b����<�&��F��t�<x)������K��f�Q`A�^�l]��\F�`t2��des�ƭ(4C���ш����a���@��qG��LO 9�..��(����_��ם�p�>�8�|/�^��+jmcD��=G�Jx��[��]���`pJY��u���g0������`��wAPua�u�Ϣ��w:1л��ަѮČ`���(͊��#d��z|��#a�5z$6�v��1���aҰ+0ғ�
&�+���c\�]ǌ���l�ĊݚBB��)����ܙ�#�J2�d�#7,>���TOq��q�=�HL����7Ƹ��3nK�:�z�
:n�zw+���b�n�#��nt|ٌ��_�(�蒅��8�]��V�ڛ{��:d�=j9�H��1��P�$�P��0y�����y�h�2�=�ydK���võ՞8H ªЯ���}1Iԟ�
���R����ה�֩�y���������c��>p���:��yî*6,� �l�p,�:\�(��ɺ*s/l����Q-�B�O)��q�{�E6S�u8OB<Qΰ����p�v�:�JTұ�.�.��+f�]JI�ʡ+e!�-�f:�Y�҃7N���FurB\̌�5]�\��5ٞ��V�@�tSU<#��{"��T�j��Q��@nf�q�3���2��z�Wd���R:1V׼W���q�'e��6"�3�}z�C�˅���,�=n,3�G�(g;�a
�K�A�xq��,U�Ȧ�B���sx=��GV�A=0��%)�}�-���*�	�3�Q����s9F�XD�FЊ�x��,�Dzz�uuO_h��o���Tqx��'e8�f�q`�~�S�O��(;��H�8���t�mZ���v����`�8��������;���@,ѝ��DcH�!�C�*jqR���tifG3���΋����
e��(WJ�lwuF�����6.�.�Î$z�G9�]���nT�N���{E��cV�{�r[��޻����p��v�s����7�W�o��H9tr��q�D��q`�E�	�Y�(U��q�3V�;גݫ!�9:v1W����ײ�D�W#o��u�N������f)CT��(���:���8y���������j��Yyc$��s��C"$n����hf׊�i�Ӣa�����V�0����u��'��`��2l�m@�
�2�\�88�N�F"��6$&}q�e�y�v���n.Z��Q#��M{�Y:%F��Um*�_�,xOJ���K8#C��;�^�KV&�!�l{�}��<�/T�&ʎ�#N�dfDg*�(gz��ٮ�&꜍i�s����ow#9�|ue��jk^U��t�B���70�\-��,!�����Sh����{��^��!���r��<�qM�	��a��1�@hYʯ5:hYQSLj'4Xձ�.sk3zj�iq.N��uV�	>�nP��!#X�ܟ6ϕÆ^��HĴ�{�e_TђTm�8����J�$o>��D�隕luPf.�TZekR����p9�!����ˤ�,_��7����$J�:�t���^=�Q��o�`�tp}j���7����։�;�Y̜����-ARe����]3�n�f��9�'OL�S;{q@�:�R�a�r>Y�/��UBO�G�����.��j�ѧ�,E��Z��Yb��f%U���t0~��B�� tvG����0�o���q[�n ��b��OI���M�4k�'��WR�[��wi�ϴRZx?�T:��
m�uO�;C��g���39d�����g��О<�e#jԢ�̩�1��ߒ���e������P6֖H=�Q�7�UaQ>�+>^,J�/��z}kܪ)i�2F�m
����N,D����5_1$�&� h^��y۞����b�Mg���la+0���-�����^n	�j(�v��2���{�p᏷�{�b�P��N+��8�<u��g�@Uu�r���4c*,�U.E��s���#�u�n��P���]��8�6"皯LE�b,��'�:��!�'f�U��hb�\w\t12!�ȃ>�ZP�&�Bz
���B#����J��]�m֋�.��]t���<�X�b3[�)��B��B��ύ�q�u�=�|�V�(I�����,��v��rv\���k�j���>=��m^!-H���7պ���� ��!l��S�뎽���p�:423*Ԧ;��ki��g�\2�P�׵�oaV�h𕼪�p��2osK�r�I�Y�wSs��>p+pl*t۝$5��I{f����RlO)�r����1s6�h�:j"�u/AB9��5�h�ZBE:���T�C��wM��4:d}٧8��r�H2�Md��_=�)�-�S����
�}����l4�q���mK��c$��j;]¬���A�.�9ceC�`��dMf��,�r'k]Gr��c�P�;방	�2����v��}��9ż���{�2p.α{ε�@l"�;����ɖ�XlN��A٠Ǵ�5@�٫���Wbv��S������jf��2���$ut2��R�d�Ҹ�L9e��r̊n� �d�K���3֨�+�+p���[�CП'��¥�Rޙ���b�JؚI�;W�2�|��h��*����T�WF�Tn_^7�.e<�H���lhҦ0nt��i����N�V4�q8�_EvK�R��ÐG]J�Sb<��P���J�s�[MP�W�P��N�Y�ش��z��XP衽�Fyd����wu�EY�x �WL�^n|r��Y3�-F+[q�z��w�������[2�x0���s�5E��v�&��sC�{�s$w�5j�fm�/jl�ΤKOfg�f���^�*�P���FUo�w���3�-���$��g�U��]m��w,Q�bl<[��'�/ytum!� �:�9v�w��O���*���I����-Ȫ���nYu�����b�pɀ�c%�'5e1q݁�-��]V��ĠGd��[�*�%f�0��t}���Z���(��m^D�����RȉMiZ�$6
O3-���O��U��ͧW���]�<��'��.lX�:�Xo5��"�c�|&�
2�=�*���0D:Q����V��ɱu2��x9��rǥ]��Ͱ+��1��a<	
����(E�*/��ʺ�6*h6i )T��o�2�}����XS)��(�����>��r�P������sp�5�:P�fj�Y�RU�Ƅ�Nv���dC�F�H݋BY��N����&v���dK�i�$	 <��,��o)#m<p�9��JM�1�F��$.͛��'ү	Ѕ7;(����TΚR�gA���[��U�����v�HL-�t�F.oV��W��9a�tmTE��"Z��Z��	*�F�J��Xk�[�����B�����d�M�.��ˣo��x���B��!�&���xe
j�HҭW��<�p�p4рT�
J9la%�S.���*"UBX��i�4�2�,�k�Vѱ�#��N�`�$�yu�jȊ�k��K m�2׊��Ec:�����-4�aY�F��F�*J֢6��d�����J�[e�UjĪ�ыcj�"�ʩm�YXV-eaPZ��� �V(T�RV�-��D��X�kb V�"V�ֲQJ�X����1b�
�D�B�R��aZ%�(�
��Z��6�[[XTm(ZX,�R)�AER�hԨ�6�(�"*(�h��*4��Ԕ�(�Z���jRڵE�J�*��Q����"�k
��$��(�2*5(ȣl����+�4���B��
E�kJ�Z�eV�F���iF�YZZ6ԊV��YYPkb�ؔD�Ѷ�ڶı�*1Qe�QUk*�e-��2ҵ�U���EYR��kJRR�Z�KJ(�
�(�AU��Eh[k"�TJ�m�j�[mh�VT*V-������*�Z�ѥZʪֲ-e�m�Q��kT�R[jQkem�)iXVQDQ��������,D~ ���Q?���M߻x��g^�a�kTm�M9��o*W �C���5�.L�m40l����Sk�m��\%�	�13��T�G^[����%�h�����ON�4���r-ֈ�A<Ks���)11w���r��)>�gv{P�Hjp�W>��.6�]2ok�"�',�VVT���<O-�v�V!��O-��Vvf7HN͹�|6���
���91��>�-N��_>�~��6�r���lm{G1���ݔ��W=3�r���d�&w�:�3�I����4���-IB^/���>8Уo���uϧ��V-���p�ƥ�Ϻx�~���"���RV�`���A�Ɩl vK�^�J��؏0����Ǖ����Fv}x�]@�lÌ�[���ꍾV��#�\��p1S�ߦ�҅��ugO
�A���Ia�ǯ5Q��47�D'wf�A�OC��X��{��R�t�Y7�Ź�B}}|�Hi��<��|�:9Z&�hb���rA魇AB�^����^�Z#�ي�>�p�X�uIn�&& %\�A���L�+�TN&m/Ys�z$�fGtr!�x)�.�x�Մ
慨�Չ���+<�I�UdO ��u�}A���2V�2NJ�1�M]�I�r�U����fi���olb���)/e9,s�ͪ�]]���:�f���e[볼�N�\����7������b��/rF�*�51Ĕ���ly�K���W3�rJ*�H�:v��!��b�5:�c=3B�tǎ���lG9�'�/w�#I_�z&���`��v|Y�66����O��ݖ��U1*�H�|��n�ί/��{cm�y��:a�]�y��S�v��dU��O�Xo����a�����y��M�R�G�M��w\�i���%C�ʥs��}����i�:.:|��_��މ����L"��i��x9��p�]\A��·#�x�Xf.����Of죢���sbV�U������Z��d�ynW+��Cxw�d@���rX:P��f�y�{+�O��:�ΰ]+��kĠ�~���a;���ߨ8�9�3�b��+VX�Zb|��K�b����iÅT־�,�5���q����ÁS�rU[��HAy�}1~`S팔om�f�pu]e�S	
�gz�#$��Q�Q�U0���ʡ+e��R�Ù��fJ�x]L��������kJ��buK�S:n��Gƽ��sҁ��:]ct��<!��یY�*c6:��$M��5�|3��p��ռ����gS	e�޾ί:ʵ`�Z�`[>�˨/˅���f�P"Gs�4�!,n��ϧ�__WLYT�����w�����Zn�wl��Ұ&vly�l�v�Td��h�\v����;����m�
W bmf����r�g>��y����>#�*q>�T�|~�� �nU�!x���{��r��zS�e�Ն�t-���q�iƺ
�v,�
 ⾱ZG���ɢYu7����vZk���_�j[��(��� ��.�G	�q'��+Y�%X�՗}�݋�+�H�I�@#�^WQC�f�/y�'KK�-P+�7TQ�rǸ��*��Ĝ(v�8�y���eIĽUgh3b/%���M�"�c�y<��xé���=y��uq�=�{T��-���W[]U��`�B,=�%Yw���q@�"�w��CX���j�X�*�R5]ifR�@��2o�`NL�/�pY��)��X͆�@.��']=��m�+kQ��$on�;M\L6���E��c2.��P�]й�@�I��7/����'�Ќ�/��-����inh�wY�o����i������Z�$`�ꫭ�ݔ��Nu���!օ=Q�H/��{�Ȗ�SyVo��OUX�g�Y
���P��{�K0C)�:��*aH�tL�w[�eHܺ���V�X�h�<�<�q����^�n��ͮk�&�*i߇Gד��c37M����t��T���u鏛�Kv��Ժ�W���V7���2)�SxΔ(*�`�.�+��l�*W-<�6��(-�ܡ&S���U�[���W�����+�7ANF���S�<���SA�w�z�;1�Ux�?g�GyL+J���ؓ��V�	��qX�$�������u�a��j�P@�J�iIB��(�_�O�J�kU	\H�����C�S,>�J[��V�f.���ﳫ>MUԺ���ouh��0!]��sc�Mm()��{��:z�߸�b���������
I�uJP�ZtsubF��d��5��ʄ���	BuEj��+DrX㰽�g[䠪���A�ւ�;�i�ok��bھ�H����AbO�nW2ņ�
�=�/����Ҽ�{�Aٞ�cI��%\"�n�`ߝ�������2�(�L�/��B��J�ޜ�����tE��Cki�6�M�-ƚ���	ł���{&�������)��Y+�K4fW�����$2�nI�]�&��߹E[D؇J'��R���O �}N��ļ�=7ӈ����4��\Rjǽj�萶{�)��C��,隺�u��p��O%�/>y�)L����
@{���OY��4]*��ux�����FM�,ڮ�i@<�M��-�o/����-�u��V������x,��7���0��v<Ӳ�c��]�GF����u���ui2T�ʑ�R$7Sp��k��O*Y�s�BRGR�<F�D���0���;����J�sM�`�<�F�/����QV�x&�>����c
cbi�ӣf>ֺVU���R��fk�U����@��]f�׹�.���{� q��N���'�@冬��-�aac�>V�t������`����z�O��}[�Xj�$C�J�k������/��Dk�Չ��E	����9�ێ#E�ǉ؆��sEиmE��ux�n��ڎ�Q�#��ǹ�a�+E�`ߌ��Jz���$?�q�p!9�R�����Z�9n�z�+8&��0eJ[Q���a���\�A �M�C������X�Kmf��ko��ݗ�4�Vd�N������0���[�q�S��R�t�Mu�am
���i��R�*����_v?о�_^:���}8v�s�2���ճƹ1��]��������|ǨQ��U�l+�f	�P��Z)ͷ\!�9��4N��dq:�5�9�PCӅ�ջ:�yl���n��
���]ɋw�kd�#�εɧ�R'�ʆ��RY���|��!�+��e��12ڻSg�	���V�J���t�h��8vf<���8s�䢉�]��^^yY�(��n�oU���l3�m�"�^������Ԍs������gm](�Bo�X��O�U
��𼖝B��<0Z�a�g�76ocq�KJkuyҏs+ȾT$/_H>p(ǭ�݆՛�n�C�S�o�x����������W���bT�ЯT{'�a��^�Q���NW�;�'n�$�4X.6i��ݱ�Q��d�Q��$��Բ���"&rp���[��a� ��n�{5��ZS?Y�@����B�"�`>j-��!�c�K���>�+�S]��E�����u��F��f�*�/(�Rg�T�,z��ᛆ�/f����4���
�f9X��ŭ��U�H͗n���mh�u콤1C���A������,Ol^�܋56���ܬ�gԝ�i�L<��
����6m[^<%Vj��⇥7x	ڐO5��ֻ�R�өaG�	.쌈-!O�	?���!�8��g����0�Jɘړ�kj���V&���#��`k+GCx_�$�w�T"z�Ju8t�@�4�9�^y`դ��o�S���n�������JF钁�Wy1���(-�T�j�U��ϟm��G�Քz��)I6����Nv۶啻]�vhL΀m֛}6��en�'����e���B;��Ui�7��F�#�α]���B�R�{��X����!M)o��0��V/�`�h�,���+��|e��+��7����ۈ,��`W9
s��>:x�*����9�N�t9�c�T�B���w*x7�5�|�6��2]��CsA�'=���TlLA`��Q��gOv(�	ȫGOA|;��iIT��q��zk��L oR,�ɏl
r&B�L���.Lx}-*i�^�I�y�橓���Լ�{�_U�A�܆8�>�+��1�mE���1&;+��s��>��4_{��guP��Z��ȃ�棏ֹ|v�A���*�u&�c1�[G�լMp�l��7� �7C�if&_V�����?T�0�C}�5��c��5�f��T���{7#gh�sj3�0\�{T2�_��Gk�	sq%��Ϸ.�f;��
[�_r����E���2z�*�
�^�^��(�qmё��q8E�I^�)�wWE����m^�Z�1�@�J��{$�ӆ��dl=A���*3��e��fQ����Y)��a:s��v��5HLdS�l\'&�+X_9�7]��3O���Lju���dI�p��>(����	��%��T�� ̽�B�%��EF���:���{��2���{ׄT�܃DF�1���A�s�3u���7K�Úmꮫ��� ��r�"�7�9I/��Dv�%�Cj����>ӇG�_xMA�X00'&��!�aNH��9ݘ����3�MV�.O��TC��0�.�"ڳ�j��d��U���:��к���*�����~J�e�G,iGQ�cG@�6�����ϻ(Py�Y*�8���N#N�*Ȁ�0L9�s@�mVr�<�Og��]c-C1�l�Q�I�L���KR>ʳa��]"k+��6��% �WO�^�ƥG^�����ǒ��1�e�wU��-2L�m��"��N�"0w�Gj�<wi{��Z��㊀>��Ø/	I��2�*�9P_Z��P�tXzm�׹%|�sM�d�v���+�ٓ	�#w�'E��P��$;�\>}�K����N X���=w�e&qg������������銍��/�5y
�=�.D�ܾTa�8���I����6�:3���c��mL3ƀμ���(�/p8�4�
�`�-3�z a��ǯn���x�����K�A�է���g��+[W�h.4���H)��:����6�a3�"�Θ.��*vh-�������ݩ��tgaM���Հ�-��H�NLl��v�݇�в���vf�[C��Vc�yd�ML[ j�p�A��������I�J�d�頻��sjgg���Nm*��p���>��_�`F@W�"��f��	e𴌷1��-��;��#H`��"�[B�L7Ch�2F��hw��9R��/Y�K۽����렝%��*jzP�H�����Q�a��=���x<1n��z����m���)H�f���xC"l�]\�wMB����B4MH�Y�@PP�.�{�2.��Ove�L�^�H)��=p�T6z�<�ؒ�ߊ�<�dx��J�:���9�F�=F�}�Ym{�x2�À�s)�ݑ_@��>�+��4b��E�'��{�h�w�UlU�S�t�`B�&(Wu,U�p,����]P�NB�֋�* ���b��J�)�8gz���>�%��ⅳ���5�+�=Al��.LE�>0�;�l\-�hS�H���,���u��I��@`9)Ƀ�jE�(AɄ!u2�kf�T���b���֤���jKx��Q�Wb
�J�mT�.;R25��c�˗�q>@Y��dܼ�LUv�xq�R�v�cyZ���݊X��}:��'�����O*�E7�X��k�����4W��p��<2j��X�wp�役u��^�rE���6�*F�`��g�M��ҿU}�Wж�Rl�֮ʌS�t��v�	eFt+:$� ���	���y��d96�Sͬ*��������.U�r�^c���-OlI��WhH�n}�$k���֫�c��^�]D�lw���T���Rqת"�r��J��1���s>����U�c���<D}�N��^`��[��R?@��y4�w*[�O>������C�;S����ZH�W��l��T�1q����ҕ�q�cRD�:j�����Zl���8;��:��N9*����ʜ�t #s^F!�Ƃ�r/�zBzי����k
+��]���H6�-|��]ܧ6�}IKt%����NB�K#��E�-�e�AC�.=���I����(q�Q����3|�J�L�{>FZ�:�2��uYX!컋�����r�(j��V\��U��!`�Y�f�q8�(�:���JX�����;٪D���ma���P��8l�����
U���>{�R�Ϣ�C^�$��n�̄��`�Ʃ�M|E���j�I����i[iɢ�R��h��8s3�[�� �Az~�ے�j�|��w47Q���t�v*S��o���e��xG�^��C��1\N�F��5��]]a�a�9��^�U�И��]�tN�mCR��i ;��h�A�Y�
..���^[�yX0��m�b���*K4��P�e��x�|Nq��
immi��ܩO ��\6j�w��-�i�.�scr-5����ڑ���#nG]R���}j�͠�/*�z3��{�&���ȩûu��M���R�켢�;�гI���m���p���MU�PDRF��6��I���ATw[)_V殒�ũuɎ��LWt�2Q�n���7"�׋"�ҟm܃�ߥwU�	��PY�ۊ�"��@�(6bй�7��G�0
QY�`*˄U�ڮ�c15*Zj�����,P�z���B5͋�W�_�fM=ee�n���/k��7��\�0�cSEYy,u���j�{^�۷�i_Tl���\Ԏ�Nu�Me����Z�h�������¬���بL�uԪզUhu���k-�����c9���}��[ٹO3�E�r���Ι8Rs�\w��KnnKb�W+���j��m�����<t9�k]�2�uɑ�/�\	��Q��z�9�w`���.��[�N[��iw�B��O��X��f<]�8�f�ŵ��Z�����-��N�v#C2�w	��J���WL�w>�EonF���I��1����
PdEj�pљG9RPr�R�#!�YCo�Ee�6C�9mV���sF���ugM|ܟÝ���.���=5�K��e���|��ū+�ksV��XA�*���Q[ֺ�;.��b-2��yl��*d �[]݊jI�t�@��(&ΔI�V̊�V�V9Q!P^��Yc��j$���˺H3��v�;��p�'H�[�=b�W!��S�.�͠r�muh�^`����l�����Δ{f\j��֑H��B��}�e��qGV�:8>Ru�4�2�1�����&�|�}�fN1�<:�^�Z��H�y��cE��6�N5�@�7����+"D�佨f�}vAt^Է�,%d����}�Ϲ���ֲn�%�X����-d���"����QO0��Zm�Uӡ٧��²XٌfjWt�D115Ɩ�5�饼D�(��*�^����R��]��f�
�\*�ee6�:�h�a�RRU������5�*�]YrLx�`}�gWZh~ζ���6��)�+Y���3i=Y�qε�z��6�)ù�m�|&N7[�� 4Z�"�K���m���Tݥ�u�wY���EL\�{�<����3���Woo�ò�\��g&��	��c`��)�/�g����L�y[B���<����ģ\�&�Q�u���
�0����`'�JWm]];z��Jx7+�f�*Q��\�� #vBϖ�:n��Ɉ*|�u��U��̄K:�ƺB���i�D��,�ik���i[b빫 �>��s	��
�5��f�Ȼ��f�s�O8�;�e/�iJ���+
������-�J�e�Tm����ʋD�*�QJ��)KIieR���+���`���Z�֊ib6��[[h�ZĩU6֤�mZZ��T��F�������`��eE�mB�m�ڍ�B��5�KJ�5m�iJ5��Qeej�ű+-Z#
ZkX�P���R)X��%Ki��E�kH��`-��´Q��KAJ5KR�UP���DU�j���#[(�V��Tm"�X��Z0��)khVUe�T��Z���m��JT�J������j��U�ij��
EFUV�V�Ph�V�hZQZث��mB���F�m�J��-��TF�j�K֪5�Xڬj���-X�j)Z��m�֭lVV,j�Tm�Z���)Z�R�U��(�Jʣb,��*Yk*(#Q�V)P�EDmh��JƂ(QTcF��V�Z�����V�2����K-�kZ�Ķ)U����E�S^;������o�<�Wk���͘i7��y�2n�f��7���I��g>�+�+K����͒�u��I�9�oJa[��)ϫꪯ��Ɩ`~�2�	��3������P'7�)܍�r���������n��<=���X������dE�	�`��$��Ү$Ϣ���*p�\&���}���ד��L?wtFX� D�ok���!�%ny���>wf2:�J\�?��p������׭\ƍ�W�-�H�c�8���M3��g�:~�M�(���;�;���S��d?3o�
ý�!��O�� }aY�%q��K���^'��i�R��AՐ�|<DEG����R�չ��u����gY^���i���y�g�c'������g�xw��֤�βmE���5��*O_g�ɴ?0�>�;�d8¡�?9��%g̔}-�?)�����~�Y��{�Q&��+�I�-Cԕ��@�8��xϙ��g���������*����3�O�:�C��Z�
��Y>����o���z�g��8s~���W��~��4�g~}i$~���=B!T�߷��0�<OO�%d��q��� QVN%f�,��HW�l3�~`V�S_Y:�t�_%�4z���:�Y�J���;�����=��=�~W�%_Wl�7��π�1b"����Bʓ��:�a�y'7��P*VM�fM?0���������bxky%tβQ�d�
,������
M��)�Y��
�Ͻ��N�o�I;�~�?��������z�U���{G�//yh� ����P��R��w��<��L��vλH,�
o��gTR
o(z���8�!�Lv���g��6��T��0��S�w������u��i��L
���!P�J�N���z�����N�D4βVo�{�s(��<��V-C�7��O�Z�wY��Ă�|���i����٪��+^3T���&��~w΅ tؖ�P&�*fe�����ݦ[X�0t������/�V9}�^)\��k{&��Nfݧ�w㽽�m�W;z�sȃJ��Ǎ+�1k�x�m�1,�'��)N��Yj��0,�3Y��8�����sF[QH4LU,B��Mw�G��oi��٘��W��>�����V�g�c9�&2zs��)>B��O'4a>B��Ӯ� ��V��]�dӌ���`�*�K���IP�2m1��Xb�����]���s;3B!t��E�"#��1���C��`z�=����OLV|C���:��O�1=�p�EĬ7w���Xud�e���%}C�<�|��d�=Ǔ�����ϕu����JO�� ����� ���j�O<q��������'{t��Led����tx�A`m�Xu1�����݇�����Ag�>�u���%E���x���.�1�>߱K]_H�P���""�}����1>g��wP�Ʋy�2)^2b���W�f�Y�Cĕ��=��6°�u^:�HVi���l;�)��Y1'�#�;�Nj�r��|��Ϲ�<�/�8��6�{�Z�OɴĂ�ϰ���aQC��(%a���1 �I�yn�^0�%M�YY��1����Rz�g�x�I�*N��P1��Vy���Z3��k���߷��O��VO�3l����U��6�RT+�~���n��y�<a��M&�$��p4�Y3(|�|�2��MC��m �B�Vv�0<jR���y�����<��~����o�?~��|}�P8�8�Xc���
�b��CL��0��Y�K�w���%@Qgy̓��
O�y��zɧ�y�sG�?0��M���3�Jx��@F ��$yw1�ƶ5���*/��qY���'�Ǣ�P�=�A�Awa�,4�V�H,���1�z�Qd�s�I�+:ϐ�Yۢ�C��'�6��<;܆��̘��~օ��+����~ChbJ��_=�}���z����ۛ��<a��C����]�+8��SL�
����X��Z���1��Xq����>g�0/���0�*)�w��:���{��������G� p�H�G	�s_L�#�f�~_K����i��Փ��E%B������O��1?	���a��v��:�+'\g��I�a��M$��=�z����|������I�<G�{�T��#޴�E/�ԡfMP�>XU��N�j�{3BR"���nf�} �Z�˜����٘V:m.1^jWdꜻ]Y��[a��em�
�9�Ø��+����6�v��:t�t�
ߔ�҃.�q�g;n���h|��t�<����4��s�}_W���)3.��۝����O��PG�G�6v��VT��0�N���1+?'���ɴ���m�����{�&<bÎ0߿d4��Y�k�63�� �N>��c������+v����;�N�r3�����O��I���aS�N��H,����2Oɴ��{�E��d�,�������g�m�H)��ʂ�3�J�l*N�Y�qߖm �a����y���*��[{_p+��;�F���A�����	�y�q'�9@��NROX��چ>���ÖM�z����|ř�`z��	�/�,�3�g��<��5���?~�}�%g�6����XA@��<g!���g���<E�aP<�ߝ2|�ϻd��
O�����Rm'�<��}@�3��a���%d㏇u�Y6�U�~��<wY���~��~�߾�����xɴ��5��aY8�t�Y�N�ڳ�i �j{O]$�hbC�sZ��>����>t�Ԭ�}����A@��h�~@!���W+DY�Ee*/<��շ��s��1�,1�z�0�%g��Z3��E��Y9���5`��������&�x§P��8�� ��[�̞&$�߾�zé����Lx>�0�Z+�#��*j���AUc��C��֧�,��J��ɈT��O���CR|�bz�0����׌�͖Ȱ��I���i&!P��>�`c�+��:î��+?7����?u��h�y�c�~�1�=�S�}�߲i ���s3I<B�`T������θ���d4Ͱ��O;��6�P172���1 �M����Ax°���d����"�R~B�������X;�Z{q$�ߢ�P��ｳ�}~@�}30+���n}�w~�L� �̇�T����6�ߙ4��'��&�m��'��\ͤm��O,?3I���뤜�d��s�����V�!j��q��C�P� �pb#�}u�����w����I�٤��z�����x�^�I]��t�01��߾ԛ�J�}���L`l;��O����z�u�i��T�o]���ZP�D]@1~�o�,[�=�0���)/�G�i�uV`�S+ �%df�â�6�*�T)'�vB[�׽��xi�K�핤��ϸ\C����k'�����mU�x��t7�-,⎔�eQ�e���.�+��Ir&P�:K��n������ﾆ���9�ߵ����o�����Y/��� �0�1��v<�g�c� y�0Y�+:¦��5�
N�Y������Aq��]��
���"##�"= F�=�u�|���;J����}���8�
�C�RbO�~N���z�����Î{HT���ɦx§mi1 ��)��u
������è-I�q��h4é�5����= DE]����`	��OJ�:|�oă����=f �aY���~vɌ���y����Oɰ��x�Rz�w��<z��x?�c���M�Y�L���.���8�H)��dE��{�8{�����%?��Ab\�_����zgI���^Y;��h��2xw|�r~j)<;�jOZ���c�c��|NZi���%e<OXmE��&�u�z��`m �b��A��==BCw�0����EL���0���]r����;��Y�O��ϻ�I<B�Y9��ް+T��3��?'�7�����+&ýɤ���&��_��7i���C~q����B H���~S�?O�bp����;��7��AI��z�!���q�!��8�~3�;H)�ď.�Xu�~;�����!P��{�m�,a�~��z�<t��9�m�d��5i�iB= z'`T��~*��	�ꜼY�S��'�Wi;�4è-g�:���m���8�"�Xk�8�a��1��>$�1�
�;�q6��Vwӗ�ܞ (����3�J��y;��O�D��@뉂#3�}�]m^|qsW�0��˔:y�����J��"��%Hh�&!^�|��<<�i��_��}�q� ��N响E!��5��&�C�Y3�����4���Xҟ��㮇|5c����C�"Ǣ�D^���x�a�+�x�:���)�f}�ơ��Ƴ�%�J����̝�
E&!S��:0+���Xu���
y}ϙ1���J����o7~_h�_4�P��B= 1�">���
Az���y�����S:�?Y1��YY�l�0�)'gs3�:�$<�i=gb�\H)��l���Xue_�
��*|~.>����s:��*�M��cm����u�ìB�U�z�̰46);��+WQ�@moR����܌ݺ��ңN^нa��7&��}Hd�0u�
����1�}�,����v����>�O��Ǆ�B�"��^o�༂m`eb'p\��R\8�z=K�f�����p�'�C�}~a�:î~�{�d�����7�w{ ��{��i1
���m�Ak8�~fu�Af0�g����"�Y}�Sz�I�v���*nj⻞������q����~e{�=�d�����f�*O]��&�|�z��ӽ�u�a�q=�kRz�:�Xy3�4��T����4�lӈN�����ϥ����@�[�p7����r��ĭZz7vM�J���z����
�
���8���jM�ө�u?0��>��(%a���T4�_����D��:�-�5�d�:���4�����S�~ߟk��oܿ��'�T��-:�!Xi6n�'�Nv�!���O+���J�Y*Az��q
�\d��5�'Y�1��|��L�+6s;�TR
N���m`hך�^]����/��ÿ}�������=a�L�mH)�����M�(����Ri����~z���ݞ0�a�?Xz�4�̕�0��������ʓ���u�X�|" �x6
�NB'J�}�|��������ݞ��1�f~°�ʊAu>�$��LCHb;�&�Rc1��������k;��S�(z���J��O�N�^=a�vm��+���1��3�%L�M򿏾�{�~|�{������&�VN%a߿d4�hW�'�{�?��0��w'���Ag�~�R{�&��M��0+P�4�;�6�_P*��0:����6���q=a�7�b(Jè{�����Z���>���$��H/�)�4��������u���O�ɴu���z ��?{��r|��Xwv�$�����
ϙ+���]�ֈi �J	z��	��p6�:��]-�W6��?w�8�&٤1�f�ͤ~T���?0�){��Cǌ<C=e�'��>C��<`zԂ���Y<@Qa��CO�
����ɴ?$�]0<�|>�="(z��?-؟�ɯ��}'{��+6�Y��b}iW0�>bԜB���Z�g�|ϝ�c6~��u���T%a��1�9�4����;��0�5���M>��dt�����{Y��`e��|N����e�n0��sǇ�ZtDiݲ6`|w�i�XR���W1卑Bݱ����Jw`����<���n���+>K�	6osz�N<�ո�ea�fު�u�>�x�Ðdy�r��������]0F�;�g��y2r��z���)*���,���x%�PHa�k�˴Nr��Q�y��ݰn4���!I����{���ĵ��𵓫k?`�`
�2T���4��+����a���O�%d��q�Y@QVO��l�&!^���>J���1�<���u8� �K�h����u������S�r釵u�ڔ��'~���0DGB���?!�5��&���b��J����d��!�k��J���1?�m�:¢�'��Ch
,���wT��Hh2~q��Y�|?g����f�D�����]����\p�p���"=�9��u��d�N_�T��]w�B��H/�y�a7�L��w����Af����gTR
k(~CL�8�!��1��bu�M�HJ��}�<�� u���?|�rP��#ޑ @�O�����m��C�J�O���=a�
�Xx�y�1�d���������IX�'ɾ�x��8��ú�|ξ$b��cQI�5�t�bw<+R{)$\Bb$z��؏@������xi�
��P�?3'Y1�a�f�I��2s
O��:�t��4�>aXy������!��O��@QVN%�oZ!��
��{�3���߫����|׼����o�����Xc؆v���%ed�Y?5�큌Z��)���A$��a��1��Ϯi�Y���ӝ�i����n}a�1���T
��}���ﳟ����4TV��.?z ��� {�*��T|�-��R
LLLO<q����,18���3��Led��i�iR^{�zé���[5a��4�{��t�Y�2��o/�:�y���~�{�����or��
�g�17��4�1��xw;�m��Y)��& )��B���
�HT6î<C��i�aP��u�!Y�J�!�>������ɨz�~�u�If�����eiH�jQ?{�G�x	�q��C�<~C���OSi��a������-"��V���2i �I�yn�^0�%M���Vs�La�و��
���I�'P�_w�~�טj��}��>���
Ο��>v����y���<@QVM��H)*��`|�{�*��{d�m�N���&e��\ʐX�52�P�A�V�cEx�����l�[YSәLŏ��{n*ko1�M����y�"�5]��]NNA�5�S���+w^����)S�Z�ojz�3�ҋ�5 IQ�6��s�b���t��jӻ*v�7���� Z��·��hߑ�G�C>��EIS7g�4��c��z��f�M�6�u���sS�J��͝�5'�)'�y��z�L�l��4x��
�d��;`c>d��ֵ�$t�����	�̮;ʾ�.bDz �H���x�������S��{-4���}ef3�*,��}�I:�gY�֐]0��y߹��X����O��1gkBÌ+��o�s���ї�\�U�z�E���(X�������*'��x��B��&��m�NZAq�Rq�P�o;�W�a����O����i�a��eE=����`���4�]�}��ms>M��,����H���" c�#�5���zG�Ϧ3�ϲE%B���s�Ci>B���1����?0��Chq�VN��7̓H
�M��i ������a��
�C_��x�Cg��6�����ز������!�=�S�}�ٱ G�D\w���M~����&+_��y��h����{�M�(�m6\�~a_|�3L�����߲`m��!�43��E���n��o����׻�����}�t��紂Ό��d���xZ�l*u��G�u�Ag̕�{���E ��s���b,�>�M?�,=O���g�m�H)��yPY�z¢�Ru
�3��������Z��y�]����=���R��y�~g�1�����18��s�1a_�>�p�N!P�J��;���*���+�ԅg���ށg�3(�79q �����Q",!���eٟ�����lg���g���]�/䟙�4��0��ϘT��
�SG�~z��������{�;d���v��7�(��
�w�I��!R~/;��P1�������q�G���-�u�;�w�x|��UN�R��Q����Lz����l1������@��'r�����)�G���Nv�$<9�k�
�4��'��2O��u+6�w�`�� �V��K��"�\�����ϯ>�{�l6ºa�r��b��'CkGx��Y�x��%@q��Y;���V
��<q��{I�0��6j�z��Y�Oq�����-*��>��P�"?t��Fv �>퍻�	,;Z����7ej����Vyw��A�7�%N�q仗��x��΁�5����o��^�um�B��Ȓ0K���Rd��̨k�Y}�2�b����b�s$����%f����Ӆu�3��;��q�נ����!Y��v����_���G�0���ۼ[@��X��s����d���ć��j|���%E��rM$�Vq-�CR|��M'��`i��=xɌ�[a_�5��6��x�c�^�1���3�T��">��r��|�����atǢG�)��m�O��ӽɤ���9��$�
��S�w'�����y�����>������b�YXÓS0�u�
��g0SW�����.����ǒ3���} v��Q)�PV>*D�8�����FQf'Va֭Te��k*ƍ�ǵ�(<��̤m�ȃ!�J_E��zT�J2��O�#׫���7�eƓ"���"�7GC�fEtg���T�qA�w�>�Q^3����y�aJ�Ǆ�����Q�*ͰWj����E����J��X=����Ϊ�4��3Y�d'�{�v��Ѓ!�J1���$F��E�5Bc&��"!�^b�m3��W�2�j\s�Jm�򛘻�2�G��ʝ�f�zp�1Q��e��;V�5�G���A�z�������㺡���|���,_�.F5�#a���c�}���IKʋ�+n�W{�t�~��
�i�Kt�zU�������6�S�p.7��*���}%�S�C�� CAKZ��H)��v�t��d޿C�x�sp��͚���=L�7��d����B�M|��TC}]:�>�S�N1+Vo5͙�{p\F�d]ݪ=��d�e��,�N����f^�ŷ�����Z�N��Ա������}A��Or�"��tI��>�i���z���U�a��h��L�j�9��rm��VJ����=ϻ�B#�	�����*!�eA˷�+1�޵�miJ���&���:�έ!ƾ3���fBa�cR;�I�$q�F5AȊ�5B���tPSSaƻ@���
�R��F��{L�ڲ�Y���{�5�U�|�B�}u�jݫ���*5���չ���9�(���f*B�Ȁ�i�Q�YV���nh�FPy��I=i]!s�lh�u���m�/��ܠ�׀��ت�X#��F�ve�_m���j�)�P�S�9�d�k���V�%�����cD��=�w�w�4��UoW>��3ᓳ41���U:�P"�H=�Q����p3�L�*�E+�b\1}c�y+m�S���eƺ��鴤�cTy_����:�	�w�c�Ⱥ�}C��D8[����3��Nw���P�$[Gn�>�����{�^�L:��D�b��OkR��xn_1����zn����R����V��ָz�r��[Ⱦw5aY�+�^^M����c��̞�<yN��\pΕ�����1�9���NvV+��t�����u�b�����7X���i3��庆Z6V��$c���TWsqy��`�Q�W���{ѩnc8ZƔ�ك�F����;�!7�~�uB��Ɍb���ЮD��eqY}t����ł��.c�f���%e���|�3b��k�h����᠂��+�O��T�Sғ'��A,q�s����[Vs;+�g˫��M%7��Ե�͈�v���S9����׌��u�����>�v%����2��.T:x��)�9dI�����n[�i��+�ݚ.����]���=j�#5���τ�!����*�����	���E�X�W�l�c���&�Ub���s��fuI}�9:�҂�.�T��K|e#�/L���\R�o�.<m�;Z�#7k!G=K��<-��Rr�O��B#t74�rr�ˤ�H���ʜO���o"����ul�<�7q���˟��(p�M�ѦXmS��:���	�a��us��������Vз}.��(Q�Ʃ������{�hS�af!��m�Q��#È����-ufn2���{s��FU.���>�
ufmL7#(�Ҳ��x�����dxNˤ���[���	˝d��1C�R�m�:�Sv�N�H)���h�^�x�=]�!�D����pft�6=���R�s��)��)��\WF%���-T˻�}�r�D�?�J�JkP�d�>���"��W׼G|�i����\fQj��.���YF��S{��b7ler�m����b�:�d��+�K�cN��d4-k����j�j/+���Ըf�N7P����MO@M5*�a���ΆZ{N�K�{�L�Ԣ�E4y��a���m��׍�꙼�j�ӥ|�*	6�9����)��Ҿ;mc�4"���s)d��u78�(
ʐV67���N�Р٭;��"ӭ���ck��U���c��5�ǯx��y�N��Y�VQZ�;|f@��嚳�ޙV�#����>4�'[GNX���s;�t!+��ݓyj�[�����y�܅p��❭qL����+ms;τ̱��%Jpj�a
�����\�<��V]H�em�kUmf�!Y;s��.Iw|��kc_	���{�)a�Ex�+���*�s�Q�Z�'|��.	@˝��9���^,���ީd�.��W.,{A��Z����W5�oA�M�$U����v��M��q�W�Q��5�J$��b>��M�4
��s��5ԩQY7�Ň,��T/��W�F�Ùt�kA��1��u������7XX��r���zx-
͔�3՘(�e�h(-����䙘�_V=a7��X4�.
^J,�{�G�xgÄGM��Zj+�(tWe��QgR��Lbç3CqG[R]p�ֺ&9�f�{�������q^��EKD����k��|(	H�c5xڲ�(�i�*T.�-'�z���R�fkcV@V�ہ�.l��9䱕3��������oC���b�.��=�]�Q"�i�p���"�j�f�%�����Kx��D�+�;�hLF-���R�^PܴG����x�N�Y��8�W�#��hUy�_�.�o#u���(�_|iit���Z� X�ō�G�,dh�a�B�_P�@,,{%�Si��]���W-���m�`�qXb��F��7�6+�۬��P����rT�vg޺=�4�1�E#�}u�����z��u�d��rK��έl�E�ˬ�2�.�r<��1��l�Ѽ�:uz%�[7�����.R��"��;7�C�fM%��tJy��!�0UX��lF�����9wIn�J�-����ŷi��
kE���oDc�4�D(77tAê�֯d�D��1��e^]ZG8�,�rZ[mZjm����O)��iŋa9�8��+�2R��V`�O��]���C;ZT-�9���+��V�F1Y���óh��7���`���t:�T�1hq2G+��]ⱘ�C?0I�y�� �Cye�K�«r�f�U��B���2cu,�	suI4|z�~���F�UUJ�$Ѷ+�X��mE��
�X�iTV��F
T�ح�Z5X"ڲ�l��X��V�EcZ���,j�Z��#mTQR��JX��jZR�,mdQdYQV��*�Ԩ�(�j#h�P����E`�,��V��YmT��R�K

���aET
�EjE����J�զ4V)1*!�*�hX��mE��KmA,�J�
�+1�Ղ�TL���*���mVV�Vֵ֢�J%�QZ�#mV)Xc�9ab[��(�*�R�,QT���R���TL�����+PjURT�1IiTQ�+�cdR�P���UU��
��YH�,TU��aX�-�����[j��X��9KX[ciQX�ը�Z����X��kDF�E�5��V��-��P�����n�z?oY��>��|�o�1ؔ�Ǌ�:�Hծs �0����v�]�e��cb	�V	�UV`#��CA8� ��Ҋ���������sS�)Ԭ���]�B����G�L]�5�	����EϭC,��Ts�KNTtP�#jXXt^��W�4
hꄶ�sDW�ƄXo�	��<�E�k���*�����/g?r�4V���3#m::f.��~�jiب<EB	�3,}�/Bz���k[�~U�4+D97����+�����G���+'D�E+.��ռ;�J�����Xr�w�1�󞊹~1}g/��X>WĆ7��`�im�op�I��	�����V��W��)fq��q��
 �Uc�58
u��aɦ ��`�L�k}O{oy�:v��j* 'Nsr��q��t�Gՙ�B���ѰEc'Ԕ�D���a���]*�4�mCP����ԋ;�Z�����KyH/N�;^�@��x6��p.#ǟ*�9h.�{�Vyu�]�w%�CYt�z�}׽���}���j��Ϫ�9��rK�F��?��^�S=C�׭�R���%��Ĩ�q#�]V:u�7���}���p���<#-��BGDiW��KB�h� ��8n�B�Ǔqz�J�V��bf�	뽪�ܪ�:��yRp�����U��m<�Vv��ab�W�U�8
��{�½�.��^{^�z�^t}V�	t���}�mւZP�̵���`T�5�n�S܊Uf�0m�|4N}1��kZ��K2�;�wW"�y�=�{ه�z+,�0.����NH̝L1�@e@�8h�ٌ)�Y��@�;p��ۊ�Vb�=T������S4����O�θ>�z�7��)�!�ڡ�Nur���,�jZT�d\��b8pbtNܫ�5�˺`��y�<�zev����Ӝ+�G]	���U�5�ly�y+�e�D�u#�����VE�H�+M1w�$��C��9mb��q�HY�K-ʙ�l�� �B�Po҅���i�0�TH�t�r��R]ǅ�V9�%�n8�C��̈́�Jj�蔺����O�^R�ᛃn=<��k~�=H��l�����m��w|��F}��H�Y�纰��aOP��'�*�F�j�'㧚��I����|��nƇC�~W��Jll��R5��"��I�O>͡�(�v�6����W>�l�)q�h����ńp,�t��AR�U���3S��ɷ���A�н����{�Hh��$��::���qI����W�Tx��î<�M�v(��Ew�7�s�]�T�3�nbϊ],4��IfM�DFV9m˖Kղg,��6��n�㞣��7�y�ٍtv�4�YݬYS��3��Q�5E\�}ά**��;��n�U���P�NL0�ٶe�^����}U�}�wۓ��wD������9~:�X�vE�����y:6��M��jF:���Į�ys�qne<o��m����F��n`���8eØ�eJ�.�^���m+�%z�m�S�d�ʕ�v�H��F\';�w"�	uFڳ�0|�p��s���syuP o8�J��w<�܎v��^W�
�6�ĩjz%Y��>`�J��YjxP�5��KLu����FVqO�VIZ����N0��"Z���ZyJSna�-g��苽ȇP�=��)�kr��{QҙC����JCj}c�LPjU����;��hE�$���]5�1�ڎOJb5�Eƌ���}SЕ��	;�dq�^ƺ�
N��(^4��-�x���׷T�[�*ݖ0_�ֆm;���=�h�	>���h�
��(���J崗���);Dz�C1q��ܨ�keq�����ؔ]� ��NB�@,�����o7s�FM�)��7�h�2�8L��TJ�ء���3|��L瓏�ĕ��c�pu*p�ت�J��>�݋Q9��slzD=�rF]kl��K4���/���rۜ�,%֯o�.��$-�LZ��^����X�t'����<S�G1)1d}�|+v��+%�Z�39��i,��"��q�̨�NU-�lK�g>s w����7�u�YN����^��bgBō���I�:�ܔ8^����z=�{��̺[�����"��"c#��mW���6���I�n��<�E��p�Hcw]�}�������W�c�t��Tf'�⫫�*�j��p=t�˹˔��.��NwSz�ԡ��Q�7�{T�L��t�|�;���v��N��|(����n`�嗚�a)�T�EH��6�]-�u��(İU[�����+�T�?3kaVxA��<v�=�S�>6=��?�*P\{�)�i�ݱ`�\A�)(�jF��X?N:(�-��H�'���¬9�kf���J��ϙx�Mu���m�P1�㒢�Ǡ��b8׽��;�����!nl5纣�W�؞Ov���m�9H�Ί/e:-d�K�lD���ej�H��XE�d��� ��>��f��Z��7��r�&���6v�p��L�ivZ���ݤG~|#��CҚ��4��<8Qw��赆6�fԻݥ���!p=*�;���j������2���V��ʤp^���f����E�A^鸤n��Q�If����@���^��0��Q�5�|���ڋ�\�R���8��/0n�v�i��N=�!�ھ��@�&Sq�#�����z"=�Mq��%�iE���l������C�p�½�͛uSq
Y��<v&��,1�Ż)E��-���~�d@K�{;c��Ӧ;�;)��{ڻV��n�9�|l�
��<7���ʼ��N�>���:Eq�\u8��x`yZS�#��B1��%���b�3N�++m4>�Z#��Q���
ue٘�#+0P��`7�t�܉�s��I�z+��N,ծ�E5��.	�vxGG��0���AWC�?g��:튭�;;�]Zxڦ������	kؔ��Nh�#�Qy�gL���;3������7��"�=V�
��P��7����'%
�TGL%���V��p�a�~�H��n�g_\�QN�*(jp��}48���F"��;�"��&鎉�ť��∋Z��-���7}�)�T;�Ⴧe�����MɁ��Tb��1~n�y����YRY�kVl���u��|�%Z��O�օp2��1
���8P�)���=���N�eY[���{OfK�8�1��;�8�ܥ���c��0��cw���S	U �^�F�Фכ"�4���R-Men�9mfŕ�	Ǯ>��A1�Y��$�&R�C��喵�� ḙ��ѣ�f[|�3�,ؚ�X�񥣔�tq��Ϗ{�  �Ǎ��50�jԒ�pr~�R�jEw)<:����Z��僧ڱ�fP^>CJ�ã��������UƍȆΎFW�P?�h;81��x�5E��P�g_$Gvof[�֭(�"É�]d���6��N8�!�#!h}s�F��kP�o�q�-�5��$c����c\L!�\2%vZS����F87�ǄnC�ЁU\'C�.b��I�ª�S�\t`�!�]]P��Gr� R�@�c�x2�<%�1�tsubD��y��YŰ���5�wL�����u{��9C`�WM�;��:��_�S|P�!��7c �v3_&-����s��3��S�N��9"�{�jū���;��r�*�����+{M9t˞:N����{~)��0 *
�r�>B k��!m��2(���6�rk,;�1����n�m�m����!�wqJa��gD�춉�h��pA�I��L_(2�)#�j�N\͈��3��������� �,�ƗP�l�~NĦ�tJ]A���1���*�����C�8�M�T�Ы��ѲK��/�����綇���[�C2軦�T���ׄ�s�ۄn��ྫྷ/�U��Ѻ�QT��c�����T'N��،�K.�81��ś�ѝ���lB��s�t2�٠���f��,��9w._sE�����x{2T����nF �Jf��e
�3n-$�#�Α�qe�O*�S�T�#E�F�oW��Z�K����a�6f�<ʰƌS�ڤ�M��&&F>�('����zd�(Rw�%ձRg����I��=��%��c�j�XS�V����@`��@�����u8�w�1ա=�9
F��F쀊z�9%=Y^��VhNEl���3jy���G\�n	de�yZ�4`%<"�]�W�pNb�je�J;4O�AN���j6J��7��x�VN;M!�4Dh�ڲ���3a߲����U���yzg<�8D��n}��nC�x�u����M��3.�9]� �@�z�9��4p;��7�SѲ3��8�iX�X�=���b�rqS��o��B��q �4�^p-*���n�A�r�^c�3̾� �˓S�i�FCr��"�]��2(X�*YQNsxT_Sp�c�c=-"�#���oc]W�o_��^��;SAxp� �O$x�Ș�ԫ�#�{Ҥ��¥��cx�f�Z��Q�ʽ���u��aV�`�v7p�'���]�u�@,�������]�K�W5�v���/$��c��۴R�O�,�DM:�Ρ����ռHTl�X�S�\kv�#���hI�K�]ҴSް�=�s/��]rh�%���1��fd��R2�?�ވ�z�جm>�z�nJ��jd9Փ��|�b�Ꞅ��!�	�p+�?g�����{�sL�Ω��(�B�sz��Ξ.ֆn� c^���4A��C��h)9���֚�S��̮z�Q^�z}�0��1:��O5��M3erq���rA��.Y]o{����W�J������N1�=@�mP���!7�=R����s�1NA��b�׀Y1)XZ���4�)j]ݽ[��=CQ������"�*��:[1�('=	�1�o�A�m��}��kG4������j�G\^*Zc���#�Ռ��jU�='?���F�tm����%l0zכ��m���s�Kg�+�`�*�2;�UC�nZ�6�@S,��.�dN�R�o�ey0*���X<�HX���y��4��A�CI^�����+%FޝΙ����)47������Nt\�!7
�e��{����!ڔ�p5#B���!D�v<Q���TnoLr���j��	8�Db}j;U�,Gf��}m��V�CXw�Y<�/c�e�n�]f�S`�W�\�c�m�ta��}+�#qv컳п�Z��:�m&e*9N�/���k�Ӊ���ˈ�z��IgP�<�*`�)VX��� \�����Ą}[E�wR7��Ne���ouH�Z��:�Mm�R�UU}U􍉹��_ws0k�a�ԏ�(��E�0��^f:i)��*_o����m�R�cO;�Ò�3*^�v�OF���<����=�+VXH��XEϢ8d��`L�g����7�9Q��L[<.�}��]�V�V�{���/�1���7���~)�2�<�j��҇��V&�;4��$]f�l�Jw�oZ(C����ޡ�k�����`}Z�y#�֪�b�k&{p���H��t�a��/��i�-�m74���1@t�Ri=�iM��ݏTb�ze���ꢈ�����ʇ-:a�wZvU7��T=ʝ���I�s�m�
e�ן��a��v��-
 ���V��Y��r��a
܊�q�{|&:�Pb���6��}Q�������J<-q@�qޙ����8~(O,�t��ct9Ε�+\�Ť\!N'rOMʬ��p܊(�kۀ�q���\hHM�V"r.,��t%DȦ(����S�}�sW��Q=�a�j�2���4qB��8sDPcA7���Y�h)m6�^�l�m/3�Ӂ��Yj�2ܽ
�L�G��ޮ��HV�K���q�Y�R闹����LٝiA}��s�AU�����P������%ypm^��ZV��A��#�2ވ�,2j	.5jE���hV�*�"g����DG+���RE��؃�lZ+&����+��3R��
�4"s�ju�W7���:^����bk�&hB_��Ӵ�h�C�~h�y�(˽ݺ7�1y1A���؃U�l�q��sqxw���ȅ|ze-���>Yx|E����m�C�im��1J2�k{��Rsˎ	�S�ѰZ�7ƒ6y]���exS��z�����v3��;��;[�һ��ʷL����X��X�Z7hEc"LxS�k�O �:�v^{ګٙnvkYw���8SJO�j��q�s����eW�P?'�e,���cǅS�ӭ�1����/����@������z��i����2��bR�ԎK�@)����zH��)��t���t��=����v�t����p�|xS^�|k+��+��hr����<����y��rT�K�XC[���c�PA�	c�ƶn8�[Nm�-j��4�А��48�]�؜R|d�B�N�^�~�a���_�=��m-W����uZ`e��k(�����w*X3 �k����(�O5dT�Z��"y�t��-��iWu�5%_9�+nL不��OIj�[X_*�ۣJ��W\���h�۷��؃2����*��E���}ʻvp��u��� A�/��ʅ!���Y�U�Ӕ�Fhkݱ��k�YK�*q�����J .�w������֕eݗ�L
�E�s���8�����sV�n{�__.ɏ	)����r�-T׶�sG]��A���N$�Ri��Pt#�]m>�W��7<�-U�)��1u�n�Uv���7s��%E;`���PwH/#w
y6���Ё���o��M�՚t��f>
��w�
�;t�]á�K�縻(��������{Y���q�3`此p{�Xߞ�=Y���Z��D�(�v��gd81i��aTB�A���Q��k���`tz�4.���U�^A��h���b5�s	�\��µg*���%v�R<�F֓v�|fI�p�za\�Cw��k�L*��/��qZ�
�b�'|���=�������fL�}�7jl�i.]�)���d��^�p��}�t"h���t�*ʂ��˭�w��=t-�w���N�ʮ|q�Iܖ�sA�Ƀ�R�+j����T�D+�ΟnrZ�ׯ�TZ����#�`���rY:�qe�$��}��.�mM���n�&4i�[X��喱�`��N�p�*۔�rg��v0��v�t�kD�J���T<6بU�B�i��iz���GU[�3��[L�;�},0�p�q�݃����UkC�Hu�銣�,�bq�9֞�+�m���̨l.#5�����v�56��SחA�lW���ιN����O�
^�chѤ6�mcĵ1�dWV�֍rf��v��*�'��Rt��}g� Z�Ct��{�1�Lۦn�Y�7�)�5.ʺ��hD"���BR��ǁht��Lk����ڴ�uĩM����aO�篰��5�~�l@vӽ��v�Ip+A�r����Wm1����&	]0�]#�/�0Xn�;]6\>;���>0�+O#S[�0��~	'�sGw��F���B�8%A𨂫˰)8��	@�B��
G��÷�f�v�R?<)��aks�+�<ɳ������K�c�2�olQ��ޙ(춵�ZU��Qת��sN�
Vn�&R��q1j��-=��Y�f��l	Ұ	5�{Bł�L|��E�f����dr��"�m�zJ�G\�Kwҕ5�K�B��/1��
�|Г��2[��TiP�+Ef���q��4DU��x�2�:�U<Yf��f4���(�P��. r��T��$ʴ��x
�_T  |iQ�E���`�V��m�TQm��F��jQ�TI�c����V
�[m�a���KiE*F�)PU��PX�DD-�AU)V��ŭkQ`VR��
��m�k*ơJԷ�����[�H��KFL��V��cj#VE*V-�
,����)��E[Q�Pb���UQJ�A�Q��YX
X#-��[m��PR�iQK"��U\mq*�ȪF%Q��TRڋZ[������*�����e�#D�UUR��[e�-��B��e��Ŷ���lj�m-�D��Fb�hEW3Y����F0�DV[b[QA֨Q�X,bE�㈪�b�������Ш�*��P���AV*1UQ��ԕQAq�"1q�iYYm%D����"%�+P���aUYkeb�U*��Q�X( I>� Qo%d�bt�p>����:��y����n죷z]��52m-���_K��os�:��^���X��>��l�Z4^"��_}_|�sW;���%�%�3[C� h��b4xx��0p9@�=)�3�W����a�-h���SMc�3,E)��GO�zgf\�`@Tg�*���������v�k���Z�ԗGv�@�B��0��%�}tէӀ��x��Ы���r����oEy��.]Hz���-�k����;
�̀�iu�q6Y���MP�k���k;^$͝i^c�S����I����a���m;Y�$g��r���9f���ٮ�@K'B�U��+K��a,�t�8�&.��(<+��jy̗�xC�b Yۥ��8�i��u��8����_*�rP����I��=��%���jՉ>�3e՚�	�o�����-읅��q7
�v|��6UW���Fض}
˷�g�E*Z�|���&$����u����0�M"�%9�ɋ|���̘�7�'��Q��5>��N���iݍ�˱��-zz��}Cy!�7��4]�Ыe^�_�����s"IRt!�<$�-�{FM�&�[���l����.PJ���``���fEy�Ӷ�u�ڗ�T��8�e����i�i���K$'EE�����f��]+��o:�-��7�()-wZ��2^ve[d��U�O�SO!ve�s�2�i]@>��۩]*��]���着;�i��n�>�YL�����v�dk�������n���%W܈U��F��PwtU�n�o9*�U�	�tʛ2�3^p*-#u��_��#�)�V��y����{�J�����rF9���!u\���Ē�%��-W�Z:���c�`\ٮ�|[N�q<ng���7oK��������V�|"?A��!�=>��w�J���uU�ݪ�ku���!�E5:�p�O�xȷӰ�W�=4�1�#�����2 ���W��޺�sO���z���թT_�t��j�C)�!��r�]�D������iX�n;[�v���LHCȸ�ǐ�Xd,�j��y��G�����qZ:٭���=pz�+Ll��|�LK��!���+P��]�ɳ�kӋ�e{T2��Ι�W*)2�m�}i��w��},�l�H�I�,�����u�_��Gxؚ��v�Ѩ�/�r?s��k=\�+�^)ߊ�jiĞÐ�Lƽ��G��p+��W��j�?�o��uH��d���ݞ�I�h D�oc��ⷘԺ�/��
���e�)��6�a�G]6��S�������SW,Ǟ{n�p�F�=�@�0�h�:���=X:`R�\�VD��igJ���i�Y���@u����3�*�-͐[/]`���w�uL[mok���(��Ec;������,� �UU}UE���z�y�Rg�O@�,y�}G�5W�^7D�X=_k����Gx��gA��mԲK�5�n��kbPOʴD���U��`�7t�V}�y7Q*���t
Ó�}�׳�ߴD
n���Rl���������]�:/���$�+��!��A�m��f��qIF��g�\=��/����G!��Dd;U1O;�H4�o�Yb;]y���M+@���8�+��첵��J[Y��1��
D誨������n<���by=nh�����\VUl�Tڄy4�9f�$��ݪ�[����Z��GLϊ�.b8��m+��:b1���}U��Q�[kBحM�x���C�Q�Y�
�0�x�Ѝ.���bKl�T�nպ��K���%!/�yT_��lF@`����#i�q�;���� ��T�*��GK�v��%w˗n؂�k�j��C�q�]C͋nf�-#L�|g�@74�rr�lh���j�<���6��}�8}�2�a�"���K��/[�a��֝�A��kVb����e�������Uח5Ŭ�W��;�9��M��T�FZ��
S2]+�#�x�G~��ՏB�o�	��T,2��1ׂub�˸rɅ˻��<Bp�{�蓠�S�
��F��G"ȑ
1_X"���Y���1,����Jz'n���;cynl��r�'c#Ì	\��B���yJdq�N��e��e
�81��j�0���Df�A-��T�Lw)j�q`���"k!�)fD���BBo��"puH�n;qS5*r6t����i-U\�/^ϝ�M�!��p�VF΂��-�Kh4���Xo����0��`� :��z�^��8�Q��rP��eAt�X�B6r�s�x����K�]Z�ׅ�Z�4�H�,���=�ꃛ]%���o9@���H�*�e��o�[�|�'��1�ޮ��K��DF��X���,��z��*�%���C�K-�>{	n8=�Ԋ�k��	`���l� n_��B����\��0��vZ�D���R��/���e �K�DJ�۷�9ToK��{��ѳ����ծ�<X�)�ٰs�~i��uh�>���"��-P�A�P×��§�	U-NmaȞ��'E�7G_UFj���)ϩ�,wR�F]�t�-T�ĐKP�t���g �fP�K���!�ýS U�r��,M�[�u���O�ڗnN�h�&�$D�	��h]���j�%|R��v����$>}����u�i�1�E��:���b��W�W՛��6���E���2X�U�P���d��7���ۤLnyY��]5r4�3�4�n�rs�"hVML=on�J��-_(=sx�\OY]+|?U���R�C�բ1�%1-D�{�[itr�9���:Q�\�vD��*Z#DY!0{��N���T*q�5��]pA����`m�8�Cpch��\� �WAB�'�2\�pf+d�^���Yǁb=���i,�����w4��@��9˴b�zȇj���bAa�lwU�>?'3]_�1J�^Y���9�<#�Y�`������"�d�[鎔z�Dh�̭�Υ�E�%�Y[L��Hg�%'�<��:��DH�<п:�54%��V�X(�o��&Dl��PHy���]u�5Xٻ�|�	�;N�7I��V����E�q��ig�)��R�� �Z��|���e��|1��1F�jH��E{B�t#�;Ya#<��y�>�qe�A�u�XBJKa�V�Y�������b�D\�T�#��8b�Bm��C��� �l;N@�u��L�N�1
�Q�Vٛ��^qe���1`ќ)�\�r�t�\Xŕ>�2�����oHņhR�p���{wv�Ɩ�]/f�AC&[�Z
�H��}��!
� �r���SY�=�Y��tmF_!Ǫ�K����q[�I޻U��h�䯊#�b��ʴ��,>Г��İ@�c�jR�bN�6~�v��Sכu�6�@����T��4�)ys�
C��F�rWAg+39Y��k���ԥ�z���uo	�+�״+��O��>Y�Xur σ��ck�O�����9T�Z^/WR���\�ul�x��
��i᷒�p�W@[�.�B�̫���/L�"N:�k��I�/���������3_� ���Uԥ.�]B'��Ǝq��2-F5�:̗\ډ���y߻�fp�}P��0����^��I�E���G�^���N�d�Wg��H����;�X�ˉ�G�%��2����%Ź�S�%R�oZU'�v�{I뵒�&48��(<����+�k����UMD��@���p�Jۢ:G��Q6�^i��%�~�T};�L���r�g<W��B�v��V�P�=	P9RGy)�XGDő�m�ެ*_a�r��-�[�3=+�A�{:,_�ֆm;�5��f�8 ����1C�4��Ծ2Bk�Q��b��^U)F0��Ĝ52����I�B�Y1�@�]��/�c��2���"����/��P=��:��)2w��y>x�����PW�\�T�rva��8S�΂�ND�2�y
�V⇤���y�1�ujV��ޏ@��|��;�mX�S}?x����Q1�tN�sp�)�l�B��-\#aЌ,T�SVGq=�f��:�����j��ydx�V��Qht���1\��p�-�S.��덵KGU*�F�'�^��
�N<ON����jGF����I�M��HU�0f�<CG@7{X2�d
�ˋgH�iR�J\gX1�J��iQJ�j�h���h�ױ^�G�$�3�K߭i����pQ�;Lz���`�,��=��U��P�0}�J�l�|�k-�s�q��|�l���-�'�	�iq�T2U�������B��VKx����^��ʖ�W&<�z��o��/c{�W/0�J-i��d᧐���6=�H��.�޽(��#A�؂ ��qj�i���.����H*�3����!�蝕s�`���������!�5�n�`Ò�]9-5%��X���	]f�~4�7�H��iw��������ZWq�=EK���,���>���]���]��t���+���^����"�X�OP�x��
,���"'P�6/FeX/sǝ\����OK����NJ��L�q��r�a�:y�O6-�׽Hb�{<�=;\=�:�(]�EfA�&����)�VX��������qt���V��qu�tF��n�e"6��;k�-��9b�.��K�$��{��Vؽi�TU�8��D��7S\C,��:�;����9�w�*�=����V��Sw%ּ��z"p����EF�A��dYfu:9�6�r�6��D*�� �V�����}�}�3�s��
G�w���W�.�0�P<�m�[X`����wy�n�'$٘uJ����Z�P��&����S�m>�Y���W�g���0��᷈�r�S��]�p�ݸ������3 ��B�v(����GSţ� ����V��W>�v,��������b8���-V*^mzg�t-p/�s�Q��5h�u�U��5��pU]�q�ƎV�}�FUw��^'�Z��X+�����Ϸ�`ݮ0���sG]$���&���t ZtS���P��[bϻ��~H4ԭ�Kk��"�ƅ«���V"�e<�ޑ8`�7OegPY��~2�i� �3#n;��5+ޙ�CB'<����T4F���gy��]Րy��b���������,P>�rZ���&dH/�l������ǹ`ֱ��,ɐ�y$��\f1�)��F�b��`��X�N�U�gr��`���grlJw�Ǆ�:�Tf-��yơy֋��sP�ȸ��%N�ɍ�ڙ�Yǉ�Y*�;|0rPx��F�+r�I(Ut�d�NQ��DG��-�p�d{"����P"��}��%
�00�p�������·U���1-gy�v�[ƍ+~ջd_�p�I���Z��Ѵ,S�J��F�>��\��b7�E='bz޴jíqˀ��p��ׯ�X��^�ڪ�E�saE�Z5��ۊ��YJ���j�q�˼ʾ�t�E!�ß�BReQR�c���ي�=C7r�	R�Y�UZÉh����>1l]臩�_9瀎��IC����+����8�چt���7Ҏc��y�j�����7��Xo�7���˓Ts�&��eƗJC�X��)�0��ߞ|��Ϩ������t�wu��-+*��EhTE�`�W�D����1�VL1����3V��㏝�u�Wկ#��1�=|��!�������)_><2�����RU��:or(��{�L�꾰S�pLu!z�'{�S�*��ꞝ!��Lg���b�n`D���Φ�M��K��[�(��>Ӫo����],k:|��;2�<x��z�P� mq�A@�٦��ά���#hf
F��������)n�k=�E�{թubʻ��q�L��d���)��`fFi��ܧ*數���� yg)ᢲ�^t�ob�����=5ܺUs�u,R��e&K���J��ai��WY���I�mq7����q^YGA�1�ZA�Ĕ�F��z"��L���JHV���#���m�	۟�[�ȇt��/���q@�'���
������nqH��*��y�Z�9J]4(BR�{��@��Nx\�89	!��!Φ�0�K�Tn�/�m����;��ǎ�d߫J�k��P�r�yߦ@�qFE�x��D�#���|�}���;��%X��p��.$�vE
����<�"z�se�d�jS�2�V����9�i �]�����H��m	4i�袱0�w[>�cA=ƕ"�[�y��Pu<m����Ɣ��<�+��8yq7�ys�
_@'+M*7ʎ�˩�ҕ=]ϣ*�X���ip��)��ϛ��A�5K�f3CS��;�0��On�����S���vM��r/؏1�`*���tC7MLZ�p{[կ���l��5;��T�n�5s�֖��z0��2�5���e�e�vv{���*滮��o$ox��S���Ε���0�N��������'5;@#^�#ӑ�˞Ұ�ݑ9 ���0Նl����LK�2����s#B����6���Qk��mY�u"7X`�!���l�wa���r\x��/L�S�éYv4s�]�өh���e����v�q��X���$�'�6n��= �h����?�O���'�0E�{\�яNT������qPi���h$bϫ�"�Z���<^�qg]��dEρ�Fun4Ln���K�2�%cɜ��F���Fq��P}׍a^M	��VI�b��L=���p��mb(�2¹,|UA4.��P�_m�*� �]otX�F���6�8:��M�4]������-W.g<�縮T��L�ZGZc���J�Z�E.�t�ey���v��u�$;3+��43��<��]���Yز�����]���<����r��|�m�":�7��P)���L<z�Ȭ޺�	>�US[�6�V���J
��BGB��I�V�e�B+�b�w�U�4�i��u��Q H��U1�@��cU%��g���tU0�k�s�I ѲQ*�t�)�.8?/E���)��ؾ�<�a³RΧw�C�Y��`��\�Zq�p�V
�Ku��WbU���[/Le��!|!غ]���5��@��f�]l5}�*ﳻ�
��v��h�5&n1�d���Ɇ�� ��9��k�:"T#��*��sN�����u�Ը�#3���d��	!N�m����%����F7i3�8R�n�k/�ճe��ם[N��DS��c�;0�����w�3�>�4����+~Ӯ*d�RHWH�ݓB��XU��xp�ݏ_(�YN�����פHV�D]ֆ|;�wǕVM�TB����ҫrs�D�zZ,'Ѧ�������k��=ۮq&���V(��̰�k���I]8{�k���FA�]f��K���P�`BrW�i��e;^ڡb�3�R��x�3BZ�ݩ�ٹ��{���9�d�Ox���.��jV����r�'v��k^�RK��9��C�+�-wg�ܘsbz����Bs���m�\xe���Zݞ}}�����Ui��)A��Ҟ	y�ؐa[ؚ����KO<{�R�o)WJŹ��؋�i�a7-�u�w�׌jQ�Cp�H��nMiv���Ow��/N�"����,FB�xg=�:�/;��^�Av��.��)����5p���@�5�/Q=3���k�KӀ8a}ͷwtAx�+�'����U�N#]a�����+Z�eoj*vG�]�me:��}���tpR�����	�K=��LBl��ʂ����)j�� ��pJ�O�[�:B��P�
N�B��u�����4��ms�0|���0�kB��mrU�]�}�]N1��!�[�6gd��۴]��WM�E�
��>i*ƔHbྑ,���&���ŃoR��q��h��*|��C��<�rl9w��q�H��_m+��(�Q$J�4#y]�K��[�Dӿ�R}���sl�����إ��IlyIзJ�Z�کĽ=��|)�v�����j:
qB_7��R�VK<�h��@�do(9q�qes8ݤb��m�F�X5��Tm���ʖ �kb��Ԃ�VҍJ(���h��V6֥E+-F?RQ�4�QbZ`��!S*ѭ-�j+K���)J�*�Q��Eb�DTQ�k(�,X���[cJ���D+U�QQ��0QV�%j5��iUH��+kb��
�*,��(������+c��E�3�QX�(�����*"
[%����"���"�5%�c���R�UZ��ʸ�QQA��T�ekk3-�� ��X"�)��*V3QTr�A�V�m(����mƪ�+��1(+��,X�es1�(���J ��e�\j�1*��(2*�L����Q�mT�&[iDX���������4V��s(�*���J1EĢ�ְUb�",-��JZV�J�r(�U�Q��j��"��.Z�X����!q�$r���3,�4E�ƀ�Db��2)UZ*�e
��T��Ԡ�Aī��(#�F
�fV#�d�_#��/(A|L��}ʺr���

L�Ų����M��ܰ�!�[+����[J�gY�:f�#K��:`��)�U�AiKm��;���[)YW�hT���j��Ŷ���ȣK8��"O��<��۫%�sv�od�h�\��RK`������)�o��SJ���5�i������{���^1Ƚw�p�۹��<��L!��A�g��b�����ʠ��!��| �Tiq�^�{ �R�)�Of9����;��mnҙ¹�-kq�:n:��Yk��J�k�9w��2�ݎwuJ�޽7�0�,B�И!M�b��ڨ1�t`�u���w��lk�-"��P��S��{����"WLK�ȬSpg؏����CA��NRT��#��1��-7!���YҕҨ�6�E��)9�,��PKC�\b��>����õQ�zޑ�vM�+3ݔ��P�G��s��p�_���t���HY��(ζ��{�)�EB)�ь�bKc+�a�L�m�2�8�j҃D:�;�䔷z�C13�O���Y��$������m�^�]��8�!���g���E/�8x|��K�+�M�k@JO�׊�h7�w�׬��Y]�	O��Y��w�B.��+a"�&�B��VHy7Q*�}�yA�C�������K���poI<�Bi.��;	Jn�+I��#����� ��{��B�j��r��G�-����<�����pXz�[����x�������[���R�M�/2,�n)gfǐ�h�v�,�#���N��Ⱥo����_"��W�N���.��92��#~3'�[0�6��U,Fg�>�;�3f�ׇ{
Ǽ�.���mZ��u`��A
g�	��3Iу�
�^g���f.�Upy|���嗺�����	^<l��s/��bv�o��b��YUw�Y��PV�o�7ju�*�کO^=���~|P�5IR�qM�0�0��,����Z��N�"?�K���,�ΐ�u걛;z�� ��(�><YPC}��tȲ��tΑ���=\oΞR�\���Q�՞B�o����jtO��(o���k�n�90�PYt�W9a�.TA�݄T��|�">������z.�o�����k�[R��?�R�g̼>�!���U�[�qѡzz�g3#����.�ox��������,�5��5AN�Xo�:�$p�tqw���7|hY:��[����"���C���q�gʝ�\0��*�������Dqml����#�EU��X�֍F
2�y���[�/p޹��Y��@������@K�e�s�t͎�6O7j�Ƹ�U����u��Ӛ���sǷ�]zh�+��=�9���')�)�������S�3��C�,ʗ�f0\�wcY�,rI(�>o���ٻӻDn��]!���_��F�q8�R�n�H�{�"P���@b�C
�3��]sz���7��D�z�ȹi�3J�q�l@��M�^/�RQKhNh�(��9�sv�;����1�)�ɇR��Bj,�v�a�b�呷��Qu	��1p��Ћř{J�OU+��M�II��*�@��Ŋ���v<��^҃��x��uK{̂��[Qס<��6�n����Ѯ}YSC�z�j^���t.��	���*���A��95dnx���Z"��M]*���Ch�����O�1>�[�\�;j�^KF�lT&���Bg�^!���{�FI��=y�mEAv=��j@w�V[Vp�{ʄ�!���v�y��
�W �e���Ý��&���y#܎�i��7�x�fW�HÔ��Z��J�b�=�f��EB�SY��,|�w�����E��p]DW���n"Z�L�MVzz�M��}v�ƚ릎x$"�Nr�w�ܧu�C������'Muɭ�J�U����>�}����G���=���2�߯@ïL�������������<��
0�÷�#.�ߗ��+)W��)זts���I��e;4��Pr����Pt��ss��SGsh�3_Ĺ'V�����*u�xO���B�ga|���כ3�f\�j�PPp&u�֌���ؒ2���ZڦEhTE�L�0{)�#}�\�s�*j������٬˭��u_-#0 ���� tv|�8V���V�|'�)_��ႎ�O9�i'֍�L����<���;��U�u�.��x�}qj���T�ե	0'.U��5�n���,�o2��'�ֲQ��Qge��x�--O.�"�c8ǝmy��i4 �	](�8��AI����&�W�RK}p�4D�d����54��i8�Q�v#� �fY4�����&�R� ��Γ��5e����lvyMXb�e��5��r��]��@���^ob}��)GT%�r���B"�q�y�0�z�K�ΒW#��+�q���=����7�J�k+��4}�P���X.�G)|U��u�6+��C�(s?N��v��)�d~��&Xݡ���R0�v��
���QX���;E싡���
K�"l�ӵ9O�>�<y�ma����A���*p�B�<��!�q�Q�+����qj�sO�P������s�d�O��yƸ��>^�v_݈XU��U0 �"(��y�;Tb�q#p�j#8^�%�lM��V��oA�E��;��K���� Z4�R{5䮗DZ�9�-υҬ���C�n1d�#��G���vu�L���g+s:�.&T�nOL����y��Jsf�mڽٌ�5yPE���K)�'2d<y�g_&믒�򁚬��v�r)�V�H�C���mn��%���=�rF��Nr��s�u�%��iّ�q�
1׋��Uo�E.�5靡�H�C�������e�f/�V8̔)@�z���GLc�~u8���:V&F��g'MB�\��0`Wt����a�1MZ��5{����/~��	�i�ۼ������Rw�H3�r-8�8�P��0\�_95���yԍ��kJ�^�\����0�JE�9�cEj��u8\*1�r25h�4�y�B�+Vr���v����vK�#O�+��H��6����t9l�oz�W�d�bL��ۘV�� �NNQ9�[�܎�s �\!�����#'�PX[�{l��ߓ� }�rm����s&�ݚ�H�u;�4PZҘ*>�E�6>\�gހ�r� ,�k����4YGl��U�Q�׽�W^�����ģ��P+i�|eQ��_W�S#ƹ�©�::� 
|�GeC�<�=8����m%W��D�@%9b�L��b��+f�%}�2�t�1�l����lmd7m�`����u�QE]8�`ѩ&@�t��DӖ�Mk��gF���e7��9&~߳��(M��5���U�r�s�]F�O>(�T-�W��|3e��,\��	�"U�bF��b�ӢՄ{�PC��a�Ǿ5��v���U��!\���s�#({�e2J2C�v<uHz]�9��&��Z�gj�f�������Cl� c�}94����P
�s�sY
C譈f�R|��c�N:ML`�S�͗�R�윩Alќ�Ƕt`bʀ�/t�P��[DHP�������I����:�}��`�gdd4���E�]�Y��MY�⫢K������܈�Ѷ��)��H���X�KU��
��F�V;�,�Q�sX�VxR�|���vm�۞�dϓ�����#�V�y�;�å2DY���Ϣ�Gb]�� �^����8�_��9wV����sݱ�x��*�y]�G<��,�����V��e�L�	)t�Vw��ֈ5���7�0��oIR�rۓ�[,���k��$dvd9(^�L����ˈDd�j#��*Bj.�p)��dX,ΧG:F׃r�.j(�j��v��PW�o���:P;q5{���v���^�gp=Z�jt�=��^+3(��}(�vWp�`�sX�2���jb�uON�c}�V��/
�]�x֘"�f��������X�K���9]�ոzZ�� �z�����F0ʙd��}�:wE���#�Ψ���ا<j������;e�{P�ʷ6�"�;Vs�%��V
�8�m�\B,ËSHx��Z��/��(3�~�\p`^�	��pVcMaY#t#.9qb�th��D@LK@lY
1_]H����P�<`w��թ���;�K�|�ׅ�]A�]��2lgЇFB��$�����8�R�M9�c_V�������֩;�N+$ub�ֶ�Wj��F5g��u7TQY���� �+,^ì�g"�b,l��6�a�&^��ȸ�.AM�ej��6G8�"��`�D�[!I�� ֍푧8�K���;b�s��%Yo ��w� �&Ff�OC�#��tQ�yDޛ�|�5F�vcz�����!^���ޟ��
� �≨:j��\<PrxC2� �
��:���"�Un�F%{��jW��B��}��RUк<:�[���F�/Vx�b:�f�] ���$`~o��[Zh��v���;Z�W�Ѳ�	�5h�}�WU�d�ŀe>��1�Ճ.P>��S��]^�{�tm�m"�yE��46�JԪ���0:�K��=Z���S=���ipnI��j=�8٣��9g[ސ!�-�,��VP�\�ڻ٠e���BVn��BL�5�w�<^��4d����o�w"�o�D���\2%�w�V[B�k�T)w�E� 3me*{c�nL��/��j�E�z�M�X/ձ��	�Bؖ��KTnS��wY�T�%U�)J����F+��Ƀܕ��7Ӣ��
l�+�
��g�����E4ۏN�c�K��fa.��S���*a��L#2����b��3��9MlzU����o����T}$}�k[Y�i��W�_-�ѡ��xF�8H0��ŞslA��V��%���{���F������e{f�8�W�ҸR���=�E�c�Ɓ���݂q�A���U,�|eShx��������*�9�Q��`��<�<�il�qR����G�)�3v8�+)vʎ!�p)�͛��I%��7i��L��^�NV��<�+b���7�xK��B���F!MwEVf������Ti�6�Ϥ-��eI-��
�DH��m��SR�ٯ�G�g�V'i�.�ž��� �6���jW(2���o�a+�I���8;Ն-�C�����W\*������in�E�|�d�zQ\!n2�@����[0n(kE���w��C��oc�X��<�γ[�yn����up}1�`���J4�׏:��9�Z{%nit4�ֽ1:@�y�֫8��zv�]��N|�h��'.��-(N��r�䗏��G^Q���y��ɺ[Am�\�Wf�.��0��u�Y�һ��z�ڷ�\J]MG��1�7#����݈
K,���.n'C�{RU��J/u��`�"��R>�wE�i9��ƨ+_x��Q��V�� ��;U�V;���8[�}��z��J[t2y��=�e���N�T���Pw{"�Da��}9����;g�gg/ԡD���*�32p���Y��r}�AS�r�����*=>`ϕ%H��֙�Ig;D1E�1ך\�DS����W����ZUL.O��1��'yݽ����!?c�ht8.���)�_���4���[�ޖl<��p���bc�U��ѩ#ڈ��;��9��e�Ѕ���(�iT�*�#M'P��nfh=y�[z޲��Ej�wo�{�R��(�q�bi{J��� B�\�y���&�]�5d5y;UJ�S��I��>ǐ�r�C!�,vDMSF<��!��peCD̾�� H��$�sZ���oo�h�LoG�]�sW�T�f����\{E�����q&h�.Ful�l'tny �U���-u�˾mj�LW{5�Y��U���PZəAP1���[���j�6���Z�vdn��.�`���\�s�ʴ���F��$�wBj�))�Mޚ\I��v-S�h{AsA���]�3�!	e^�s���O/��]t�=��q7t�zɞ���Ǹ�\��agІ5���d�M�7�M��'~B���WF����WU�\��:��8ٍ���\ҏp��cAP9�
1^�>y�S��2Ŵ�s��(�t&lYآ�+2�v%V��*}ND�q|�|g̏�h���]Ԇx�W�]wؒ��7%��r�c�,\����bV
bGw�3|t�#%9;і�=m*2���)#@��!�mv�P�$�������q�J��xꗲ�T��*�)kOM�V��r���٘r��B��r �>P.'�I�n�ŏ^C�7�8��뜉�=�nѬW"��\�_w�oIw������Bq��|Z�l^c>���a\\�O.&�=ӣ��v�-V��e�p{�����9h��@��\Ϭ#;��ݬv�s���^BmQO�T��Z�ڕo9UbC�����d�jmF��+*�R�%	<��qڦo�5�>�<���2��m�Ù�PA��Q')���=��8�vQ�t:kQ�J�-�Kg���"���ְ4�Yv۳���՛3���|2�ȯ�k)&B�CȲ�J�a*V��b=��P]�#mdͧ�8�^��s(m�q�C)���1Wl��[��H��m♉��;�wb��r���=���A�/wae[����O��>�ժ�Ȼ��Ol͋�!�u�u$-e�9�� ���j_*|4�V��n6���
�;-J��&���C����*Zۡ�'�"e���G5�o�m`���A�_#k��O�\j�nr�kh��kcT�{��u>�.�.wf��m��4��6�r����QZr��R����(���N�Ck }B�6/�[d��u��&]4�&�q����U�� ���r��净�R	�\��2HJ!*��A��,Ɇ�x ��Qؤ�w�:���XI]h��e6#y6q�]ʲ(���$�h=5�L���5ف���xL����j���%�ޱ������'e�ڒ3�;��˅��3�'�*#�/��ޤ'�ம{�mŽsz"E�Y�e��)A��_8;U:<��;�t��Ww{����8�*ruĸ����X#\ڔ^d�\���y��aM`����ǽԪ���z���NM�HsK��O-�r�uq�w�1���V�ZE����R�Ю��+��ڙ�:�y��h3�`B�eV�n���9;̗ljzzK��`��z�o���ݫ(�#�i�������B\윗��e��E�'A�g�A�:D�Щv�jp���ɶ�2pdr��������$[�9ް��\����b��u��c�G���tm,���i�k��csx՛��s��q�ʖkQܕ�Л;fgX����7��yS+)jw��wW�RA+͇qY�l<b�>P�e!)5*z�؁o�0R�ӓ�+ӺQ5֨�a,z�$0� ���v���+M���	hO�8�{Y;yd�F��jU�W�A8sn�v���h� pPX0�.�z�ݷo5��4��ޖ��ao2�m�	A�f���:;��j� �A��#S�}۔����ie�Ðգз:���q����DӋT�?��"�ȳ>u T�o]����PP� r#-�un����Ԝْ�82��QƐZ�r>�j�]�2q��R�rt�C4Kߎj��n�.��lW#V�j%;]��sr�.�����	���v���kx-��&�˴1Q��*��K.��OM�`,��wt�װn��f�Vr�\�L�z�4j=��0qn�k^S,M��@:��b�\R�Wn%�M���
8��A�b�^G1�2�F����B\�5��[&Գ�j��	6ico�� �.�;��D�R�
Ȫ�Ɗ(��E�墋X�*�q,DB��b�#1����e�V��2���j�,���V�EJ�#��*����#�bȶ�5mVDUUDV
�*�F��1X,cDb-j��F(�X�j��6�YE�L˖�V֊&P+1��Uq,R.9�R(��"�PX*�,�`��E��,���E"1Km�������\lQ�*V�m�X��1Uj�+m��d�H�TQU ���J��D`�G)Ab�J�������QE�b�Q�+2��H�Q��*���V*��QU�6Ոe*�1�V,DUF%l�EEPT���R���J�IP�V2҉iVҬX���lb*�eZ[E����-�Z�Ɗ+��1���+m����B�}n.��%�+���"z���<첳��@�=�9r��9X��NL��RX�����,��f�U�꥙	�l�Ž��)j+������t/:
���yW�W�'ǂk����n`�U`WB/��C��i������"�����/���IMˢ��fǝ�|���q�#�S��8)���J��ե�]1��vٍ'bK ��`W9
@ΖD�1�yX[�m[L�p��,�*��J;�W\bA�`)_��'7{�M�n��P��MUx/\�!�*BnSu[(C�`���Q���(rȽ���n���kKJ��K�4	��Akz�L�#�c���C�q0�=Y�EF�U�����[����ռF7r}��i8���1C�q�+�����4������"�+�aͲ˺�\���z�Oۖ��M.:th��D��X5�����,�+�z�SP�lD��2%׼�}����C�\����t�,����A��F��(��`�n��әo��]�on��B�ٝ�Cl�VC��l��b�Mm��t�7�J楪	ń���(�,�y�א�j*�l`YMv��wr�2*eP>��'�4S��qQ������CA,�5��l�PR��rmb+]C��0z�ՁO���g���-:R�UB�r��t����
W�P]��3�u�L��9�9��C-�;��jΧλ"�M�&��Ĭ�S��_Y3��v�N>i:��70"��e�32�;��g�X���"JJW��ݷK۪
t+4���<n�'��V#��ۦ#n;h��N�lܼi75K���=���,�ٯ_�D>�$�O`U�
��(T�p{��|��ov�S*?U�O���k/t7�E��Dﷷ#�&����Z4�~�Vj�\��#����KX�m���Ҏ$l���Q!����YT5��s���y->�lTi_~�{V8Q�$-��C�]�a���hF@p�b9����t��5����"�a��Ԕ�$�q�y;{�m��G0Q��<89�{���-2-���ŷ��PÛ�w�&�7��ɦ"��4����O�E`������= W,*�C�ƒ��ŎT�n=#8����$fB����p�s�w^	��ˤO��vگ�2�dô��5!�k����?�v�F�bUp����#��^+�>���ΐ�0��Ŏm�>����0���-M�r����JU���)�K���_mC�'l36�� [�T6ۚ(��4�266x�`��R��.�%�V�0�i��3w�U���2ѡ�v��W5���))mk�B�F�ig).�Gϲ<^3���+5[�t2�ږ�^8#p�\����Z��b��Z�|m�O!2�c��"�b�[OVԃ�1�\6���Lj��Rj�+��ۗɫ�rq�����۰&�9���]��it�� �J�о�Aq��4��⶝l�v\.厳�l����������u���v-��[,����A�f$�d�֑�pz�|-����M9H��1�+�3���mudQw�I�f\6���M	}~�b�g`��6���:��VB(�&�ٵ)�2�P|���䛏\sZ4��������v[���b�;z�'c��ܨ�@,���f��4���t���UuL�Yb�������g�G�"�-�Q��-Kf�t�zA����N�0��J=�@�|e_l>� ���5�NQ�q�͸�, ����S%q�)�"��-'@�M�	�*Nϋ���k9�&1���uy�ڑ�Ê�т�]wV#�gEoH`׻�B��Na�Ԗ� �b��e\(0������jF��+yZX�WY�l�R�v�y,�cf�m�ݘ4��U5�l�ڹu�F���B�v)�Q����x�^�:D�C���m:gs�����f��Ҟ�t�v�}.u������i7�}�����Km�&��Hd���^�D��ϩmm�(��v�;�2���p&(�nRR��X'��U�F�Q뾵͚���[T��ח���`k��}�tF��ӗ�����0���F��;ʕ�Zf��	��+����7^4��'a�s\t{��Y,F���):�����LMj0
��H�hq��Dv2����t�Į�-O4���,/
KLn+:$7<$^8��&4ߏ����S�
�w�`t�gֱr��%�<��Y�(U�:!�V�2����i�B��,uc�}ٶ����VgC�6_l��]�-Ƙ*O�ׅFb�S�m�0W�s>>�h��������7.�.gܪN�v��G����sC��1�N�r�����B����p�������S)*���/:䎴��#�#�I��ƫ�!�P��C3���N8�SεO+�z���Y���o��8 �ҏp��cAQȶ�g�\ �g,3��5u�=.�"��ݧ����h��˻��l!`�$c��bQt-��Và�W�x�n/�J-1@`A=4��޵K{��]��Gu��ʿ9��a��F��q.�>lؕ������1N��@��Yo����ooJ��
����&�ƞ�C�f�g5ք���ǎ�p�M��(��q^��o��� �u�}�fweƥ�p�)�Ňjf�EF�cEr�7��8,e�8݌�}:
�#_����M�������ڶɾ���+�>}]�B㫞��b���ZB�K�+EbNcJ��8��i��J��'�9�GZ�~N�,�Ϝ����[Ι�Ϲ%ӕJ�,w*fth�~��[>��QN��wR�aK��onqI��!*�1{���;i"�p~LC�Yh{��)1��i��P�wAU7�卍.�y���d�@wN}��c�T����u�k��i����M���BӤ��3�2a�4l{���֐�kE�kR,yzM`����"���[b����}��1�8,]e
C��c5�K���]g<�)��oowR9��m�#�e�;lرi�h5u�k�4p��J�S?]ѥ�]ށ�Z��r�i[�Ѻ�ep�l��Gr��'S��ug���~���S������È��={2����Nk�qHW��PT'�1��u���}�r�Z�)�|�5��=B�Ɯ��4
����<��IT����P�C%\A��+��C��A	>��Ak��+����)똖�R���9�kJ�!ю.G��P�Jc���/K�ׅr?e�(]���@�fz���A�BU�n��5��RZEXCF�kzO��/j�fO��3��L�>昫�'8����8�t�'���w�5{���2k�a����U�P�so\�{�~��Q�[Z��3u�ѓ�Jf�J�8!��|2Y�&�s��gܒw�ۚg`r�98AR��o�<V�[,�,��'sʛ�MY�k�/�\�Xci��7�Kz!R�]�u�g>�ۂG�Nݓ$\s�ڹ�W.�9[���nE��ݟu�b$���lk���,�⾮ઠ8QF��G\�#C�MͥQ²���/o���b��DD+��Bl�����mE����ߔ|Q��d}< �$�������x�BN�|����uEb�u���M�eվ�9bz߂�|&.֚"�g.��`�׳J�q��<�l��v��1c;v���(	�lJQ���Ƨ�X\w��C��`�v1c��tҁ�f �pn�@뾫u��M%�Q���WTiIcҠN�08�y���g�.h�OV�xk�=�����������Wo"�{w#�&�Sqii�QjB�dY*�l�אųy�#�����}�(^A��3�p8tF-]�-���--�2�l����WC���'_4A��j�m��{YiƦ�-w$���R��X4GW�t�pKNX�yVlp3U=�eB�y(��R{.�U:���a\d1%���B�L����-2/�ĵE��=C{�v2Y�Zg�kr�(@ˉQW��S\�Ո��%h2����"�yX�l-L�3�5��PKu��u6�nqIvo��W�;���6��9In���5b��Nf�e��ƶ�^��Ƴ��3����bދ^b#�P�9M��M�Q�r�WR��a�bjּSe7����9�Ui�:��l�gO�xϟ*�9`/��q3A7Y
m�r+"�����<�Yo8[��\w�� �7Ҏ]�>�N%�U3�X�z�p��>�����]��73r��|�龝p?U��s�B��<#q�b�0�(Mny�Pz*��p�a���qw^n�#9�JBÎ��/&�'l0C-��8$1�@=\P��uk�*�����5,HG���<,z��l����dB�B���^C��nx�p�]zH����"lU�vye�]};^�;�Q�u�Loy\3������dij�V�3[O���+kG��}�7�)d�j�X���$7AE+V��v}�k^'ז��O�,��ڋ��=���z�鲟ofm��״����Alŵ&ez�IH�&�sZp-sgZ����Q�=�;P�l�a=�Pե����Љ���bb�;��
b[Ә�N^�yM��iE��3c-;!SF��>��8�^Nf�;bJ��,�(��i>2��8�`�&ҪQr��1U��5b�I�e��w>��|p�9�&�n���f8Vk��$)�A�v����[���s1ł.�U=�s�CWu����q��������3J��M�'Cv5uKDҽ\��ON�.=��������"��8c����6vm�Wo&;B�  `�k9S2:˾��BZe%�%w�>kU���Y�;�bV#����<�VNA�}p��ȧ�b�j�&]�GԼG-�hSg&0��Ɠ�┎���,�;�/&��sg=�p,� ��>��=��/.|�;uٙSB���ε�wG�Tq��ܤ����A��*����?P�7Xh�1��ܳ}��E��⌾xU��L`p���B��S�Ϭ�k��x�Q�~�rau��z�9.�.I�	���hoQ���`�~��ߍh���:��7}�n]u?��$Ox�։|��v��Uy�f͂}:�X{�������'D����p$m���(�]Ⱦ�O��@��i���U�r���/R�2�-OlIS�T�
9���yE�ޗ��k:�``.8�4�RqW���8�c���� �s>8�]+]�����bA�����׹����>���R?A�� �˨(;�
�}:GZ�R�kH�.(>��c�ǂ���m�r�k+:L�ƺ�	Wt:�KXG�1�"�d��ʠ�: �{e�~�HQU�eu�w��TH��X�mx�I��p�z.�tκ0o\aq�n��aL�6uN�����'�����Kld�;���wc哰D{�1�C�8J�t闼�k��u�Pf,�1��c���3�{�G�O��h ����?.ϖUx>,۰�g2Թ[V��I�vW5��[.;��=�6�b�1�(�pA���ʲx���S(�;r�ycѺ�-��^��-^�� ǒ�U��fj�/9�5�eE&_���n%.�-/6P�:J��-ӽ��7�<���U�����HbŘ�z�"��d�NБ�I�oQ���q8Մ���ǎ�6�/T��+���ׁ(
����`X�`���������*z��/��P�B�^s=7R�T�X5C]��ӑ�k%Ě��@���7�Jj�x�qˬX%�
7x�+���h\)�V�V8Յ+�V֣=Vqa��Tī�贃��������XX{��a�(H���6
&�4��U�'�%��m��"�ݑ��)
u��h�<�އ�]fS4�y��x`I�v�g9�շgU��]�5��vX�͖|��ٱb�4�����$Ъ�(3�&u�{zfU>+������5f�2���p%)4���w������}�����u��0��u���I8K�X�5����y��u�;lq��"7���V���۽n�1�7�=�`�r�����9>]Sr����r�ok�����Ձ���j�n�nkW�t�����嗮�ru�ۨ&H=\��ַ�k���\�d�3�jX�gZs�9ݼt|`�L��hA�/y��e�#�)�9*�ʹ̄.!��1ʹ�˝����/9l7�֖�mR��2;qIB�P�Vj!
���A	�e7P˦<�d��c�0�&/+���*�z���\�P�7d=L��Mr@���3�! &��
���<�;5�xI���{e)�ٛ�U$�/Ч�p��O��t^�Ǒf\B�C�bJ�2vZ4DZ�p��y\���ݹE��y��o��B�z���C<5a�6���zZ�X5�����f�n������6�n�w)��R��.6M�kt1]K1����{�j^� qTB�����8����ܧ;���L�EJ<�����9��(u,�P��m�d�Mbq��w�sE�Foon�����H�=��S�,l��VT#�����^��yŶ l��o�(�ɞ��=Y��˩!�h�|�J[A�5G���Xo�ME���/��ʆFn���g�ƙ�W*0�omlҀ�t���5����>Ғ�
�`q�&�5XW���W;X�hRk���YH�gr7t�q��Ln�co+8��n����.�ŰK��cux+bZM��Çx��������f�@�J�pX��}��g����K0���t�M���]�\�X��y훕��9���'EN�k"+�秅��Gk���0�X��s��M����Fa�!OwR=\�����,�C�gkʬ;2�u�Թc�x���wS��@�ZQ�!�r0]����]I�gB�8H���m�ܧ0p{�n����vu��g�^ts�D�:�;e�ʿ��hQ*���[��T��svY|�j�ԭ�۽J�Q��Sdc�.낯��ujNt,�έ%m��JN��Kye=Oj�G1�����`�h�2'uuo_*��:�ڛΡF'f�[ۙ�g5������:[����qT��Σݳ;F�yY��,>���5�td3 l�gitWBs�Z{I�����S�v�Þ�2��r����aBpF*L��<�M��J�/�
�r;�N�}Nwj��:�MI�*&�Ge��d��9��%��vsOg^t�&�n9Eū�"*V֥�������<�;���R
f����[d��h��Wɓ�H>��u�^پ��t8R@�lɛD� ����P���.}N�,�"�F�v����������+����� ��{�]��\�M�B�ۇS�R���%���(��o����.�L�48�3���*H����o���!��&�ӡ�j�
�S3:����̴���۲�ޢX�b��`��KD�MN��b�l�h����:\���c�(����+���Vun9�i;t���҉ݠV���fP�tAs2]݁O���8]5�!W���d�~#:��l̮p(v�V��),9;:��7�5i��VC��Y0��C`q����Q}�0�mp��䁜ckZzR������m�ʚ�H�wi����%b�Ӵ�R��r��v��V~�R�4�p:��D�k� ���� b��[����]���V��1�Kj��:]��<�-� �n��n7Ϯ��Dt���ꔰ��ܝob5���-�p�ψ�h��c-մ�k������>9��m�"�b�Q�3-�q<R�.Q����6���+%��-q�>�y���.Byˉ���Ĭ��޵�rY.�u<�a+U�ZTIgSI=�u!9�0k�&_�rLT/���]쇕��1&��(]vrY6�%���^R]�j�Y�x��e�d�dH;�)_.���c@%"L�M�.�ڵ`d���me��-��-�p��prk*n_԰;�<<�٠*�
q�R���f��M�����\�s����yK;(�' `��m��f��h#X�o*���դ+�|��f���놊@J׵���@S���*��%)��(�+���Φ@�ks1��W3ܸk�C\9u�y��:�҅��bj�s�Ε�^�j>'o8�e�	���WiS��^�gtm���D�Z�K���Z
�{�l�zg~����Ⱥy��&/���U��//&ĄX���Ӓ�۶Ҽ����N���D���UDc�W*�$2�+Zl����
�,b�[r���b�l���R�����J��ʉ�� �iQR�J+Q`�Kh�*�VT�*+ڲ��W��Z���J�ՠҬE+EZR��%LUm�Z�mFQ��Eڢ�E�)��PmZR�ET����R#l��*[`�)��1����Qj�Uh�2 ��bU,��m��ZQ�q̡V��"�
�*�EQbh�� �֢�J��e+l��2�ڌb���R�m�*���ҴUF+��Kk�e�2�Q�� �Z+,���1��Q�QAq�AaD�EG-1Q���im�j¥���ZZ)QDDF�Tb�Y�TUJ�(Ub���bV+F�m�-�E��V�QjV�Y���kUL�R6�U@Uy��|�޾��+w�ٵz�	N�s��P���*�)9ɋGLB7g��!\�A�`�m��:��x�9g$���zz�ڝ7�<
s��z����"�]W�����2sϪr&)����(��*ّdt��ك37#(.�����*=i�ɸV�ku���-��3}�mu\:����7jĥ-�oke�o*�"�U=�>�fq����dH兂���KT��7uP`YP�@{hh���T�׽��ɳ���oʡ���#�;=A?,G�HbZd[q-Qm����ȃ�bY�U��:5${j�U�j\y0Q�X�"�����x�S�q��Z,3�&��z���W%����-*�0�S�VcfKh���r|O���頠-��a�����)_R��n�S�ҍ���Ӷ_K����p9�!q��u�sΣ��U�qg��dV�d"��.	�ˍ�11eӾ�y��w;ʍC��:�3�˞<_��1=��k�1(2�
[��뻾���3r�_f)�����|���|�-.�<���P�+Ӡ����~s�L���#�'�A��{��uNIxl��i:
{�UC8��瘻�{�VgM~S�Ϧ'V}�f��6䬆�2���m��f9dLI�}���Z]���s:�7��TZ�m�t�0)G���׼>���)����V_�Ù�S�]|{rP.A���\;o���9Ⱥ�GG"���1�3]�A:a ��5p0D��XU/�,��{�ց]��ͦ�R�\{����R��v�
Dxmq�mudQs���7�3��~�k�	9;�s�z;-]ak��DHn;!&���j|�A����zҾ�v϶gE/����En���3��r�:k���8�,�v%5_�S��,�ݺ��V;����5��[�N�p_-k����X��3'8��G�t����DO<`�>�y�MB�"���;N��FY�j��+�R��\\(�L�t�\��5�V�Q����{����ϳ`�s�E���V��P��ӆ�X�>��5����.��fN�	eeM?Fm���;� .���aO-o�,��8[Ep�s���ꏯ�1�Gu6�r�C����t�o90y���4�]�R��td��3MF�Zz%���x&�1�&S��F����͸��.��G�����Q����}L�sb�yX+��P�8��`j)��.��w
���G4��-u�39!U�9��\�������}j�����@2d�E���u|�-=�J�;˝�Im+V^�z
sn�_�B���)��[;��lO�n���2ms���֍��+i�ٛ�KEF�:�>��&����G�q�<g,¦�Z�4ﶳ�1u�9������Ɲ�S����|�%~��n2�I��X��\8��aZ��/�6��[1J�y��E�I���u|���H��m߯��#�Z���p��S���TҸ�'�uPW#�{Nᴘ�̹�2_R�jR���S��cъ��PԹ���B6��kW�'�'Q1ګͫ�Y�p���<�i3�j�'�����n�~Te(.u���q-$��ìL�]�Y9�5bKn�(��k7����k���Ϳux��1v�BH�Ը���4R�Elu�܁�m��v���%�}�+�9����K"x|�)�Խ�����FZɻ���Re2N�߃���=��%�._��{}��B�T3&�ۮy��v�o�S���Q^�Lf�
K�"�Ý����a)۪x�N�v%�
ꁋ�1G-_�*�Ӛ�P�T�*2v�r�+�D$F���d�]�L���ൃ�X��Y�\HEu(�Ԧ.l=�~K��v������ ��/5%^,ܣ�lG��z�,�@�`r�����۞��O�nԢ$n��YnBP9��A��/	�� �
�/t�A�Y��S�Q��N�Q��j��Iy_�d��V5؝�|rq\�n�)mԄ땵U[��WӇV$��^ll�I������e:��u������QtVg��d�����ܺ���q���ˋ}���[Os����/|�9�Wo�=:mx�����'֕�f�P�޹���J.ָ]<ӆ�l�:Y���9��T�LԭN�U	�.�������HdkH�u.P��m�vn�Φ�/e6k]�����9�����sč���P�"���7�x��i��WF�׎�y"��~�|�|��&p�q�H��_�ҹ�ц&셊�cZ��u�VC�ڗGg5��I�)�Ʃn���6 j�6'�#�)e�̑�xn㛛ݬW9�'ݼ�jT����1�o\F/*���ΰ'e�Z�΋e�u�T���1��[CS+��-_:u���`N����"�܆���ZP��K�{C�gI���ZeY|���58���]MRq��Z^�cl�G]���^	�-��ð�x��OrQ����1�yGc�zlv�st	DE֦0ҩ�z���
��:�٭�h�zJ���F��Tn�ʣCTb"�W-��Jў�>({�o����O�t�M�۹JY�A4xj�ʀ��Wcy���~�NȤ��8�z.��,Z=i�����o�{VR+��Sq/Vɧ���Q�ܯ{ht��j����<Ue�W}镆u��%R�̝���2n���R��c
�t�ܥ�C=(�|�_x��pW��K��N6�,���\g_C��q>���-yMU�cV5����"�j�=����r���}B��k�ʫla��p��,����Kh��ͣp�N�mUT,ъ���r�:�o8���N;���FK���댖]�d��6Z��d�I�Z����l�Mf!+�dQ�<�_C�=UґMkt�.�!;M�����K����壏��
�z�^�����*��V{��5!�,�{�h��U*OK�J�Z��Ǌi�int#�%�5��fL��ì
�gq�7!��Cp�V�N�Z�i�g=��;�G�ջ����e�[W۝Ztm��L�ڙj^t�2�5ub:S�ݗ��l���G��q�nc+.�
.��bs��*u3,�+�˾��̶���ks1��R!-��;�t$f�,��LXzd�\�}��o�*,���А�1��������x=:�u��9=��,W2Y�T��j����V���X�ŷ�n3�O�p�ĽؾW�Ud%B8b��:�E�&�#-��'���Y�>U��q1@ԇc��Տv��nz/�T�ܹu��/N�$��d���K܌x�|B�퉃6m%׶u�H��y���`��C[��^�k;���U���dl����k���S�=�4 QT��!C��[���%�����.�ʜW���	jC�i˴�Q�I3���c��U�2���^(s�UY��9�Ӥ���ݏ�nv�jy�o�BqN��\���;!��*����t���ʑ������Ӭ\�0�![j�<�Q�w���չ.5=�,OP0�*���Z�pES�����s'����L�j-Ձz��<�v��S��(�rX�u}}:�b�4φ1y�*���5�Oj�&ӆ�G�xWK��}�}�*L��x����y�opkA6���Y>��8�W�&s{YR��C�l��)�2��W�wř��w!��y�nwI�Na�$�w"�b��w%Ǵ�Ѻz�k�	�>�b9���U�^c���j��=/M.ɕ���-���ɢ�D���;���Taz�U�̓�D�ݖ��I�ݑ���t�n��9�l�)�|�LvU�y�i��v�Қĕw5�m�#x�ڋ�m]�S[����۷<ui���{u�����}����.\mz�(Hg�4`i�Y�$�[}���[��uU��)��(O8ޘ��Ɣ%��"�����	�Wϯfz��+���Lr����5����8�O5����q����~�ݸ������V�Zs^|�F��۝Xо�b� Ö�Bj����=^�Gg++�Ԏ�m�]jj�T�O���c�)As�F���o�B���&�����X�;��˹���]O�t�)�bS; �+�ڗDXQbݑQNhv��݈�5^��7ܻ��9���s�;��z�LԞ<O���+�M��n$�(Z�����6�� ,�Nl�W�������j�����1:ڨK�^�bPE9�z�M׿�8X�`�g!��Ь���e>X��Jw��!�\�h����N)�96֑���[��j��[���"U�����ܝ�f�Q���;�29K��5��˵8���)�C+��k/����ȸ�K�յ%�u},��u�T�X^�ɯan��R���g89��/6�{�:�+啔cx仁�b]�WTX}X��Y~�6���2�M��Csm�01:��}N�y�N�X}G�'����gՍ���T�ꨚ,��ɼ�"���+1�� V�j@��!��/�1���yh3>�Ǔ=J�f�bG���vCu��r��Xaqo�5�b�˹Mw:7�9�d������ ��c����gU�j�y�g>�_M���\M�]�+��G(֋5�sT��=.7Xܿt�1lc��|��iih�\�"�WM�R	�˷��It�n8�V�\%�wx��|b�r��Ӹd�z��P�wX2:�g�<�
�v�`ҡX�"�˚����s��W��[�n��
��s���ׇ�;ay�b�<��Wq[�G{���A?an�w�*�S���*�Yƺ�NYKj2&�^�EQ��9�^=v@4����ze�X���w+c�Uz��"�u>'��]Z�]�⽭����|��㒫�ݩw��E���/u��xN(��͓|�%K��e���hwtcC9��.`�r��*&�h��F38�bKp���H���;��7��ʣؼ��6Y��w�^(+Y�1��nޚ8��V�jec��ڶ�����t�5��Tc
�w)�RWݘ������@�鹸�H9Ք57u��Th���Om�c^�#�_b��n�`ţ�V���uivUן�R;��W�����C��axB�l%�4�c;���|:�,��g���|��*{�cc�E-�էwJ.���?C��LaN��%���|&�1�Lɉ�T1�X.�bY��8�gu[��W���a�L��E(���zP*�zϋ2V»޸
Nn�M┎�-٩���-�1��I��Y��-���j��gPOLldoT����ͧ��k����Ν5��������6���a�I�n�ѹgY�+�k���#W)�#Uo;F�K��3ݺ��O-�+gS�|�6�w-\���ˣ&�4]�ᦹc��x���ϑ�;Iڗ���\�R���\��,-J����R�5F�_,IW)�����N+1�;�U��p���Օ]��GQ�MR�Яg4{)<w�F#�D�;��4���m��Sko��L�A�c�cW=�һ噩lT��ݺ[��l�=�6|�:r����oT�� p�Oj��o�7�O�@e��=j�=����x�h���/7�Ҵ�-�^ؑ���I�X߾��F�r2�t��7�5����˩��ڇ��:���]��",�qή�ZD��#-��'c��|��y��	ԗ����ҫ�q�W}癝�S/����U�o�Z�l�3w���4�fXSVJ�I]��؆T�:yҲhks딗�����^��8���
&�ֹеS��z0;�h@*Vz!�z����_m�g^�*2u�]�m.��{�����'A�ߺ��z����}�|��d�ꔴ�@�U��L�E��;��XFo����i���֩�k]J�^[�G.�[�E#��x��LP)�8G��͢r�y�Z0Vl���wh���-\e��}����a�6UvZ���<orsb���(���
��.A�oל��`��3r*&��5�QG�����ưQs��ԑ�����g
0�M��8�d�,Պ��V[+d�<y��r�C��V]zu����o8�������vrw�	��g9I`[e��S{��f5��B������0�pQ��ic�v;b��s����}Tȝ�in����N�'d��K�@kONkT�>�#��[o�Z쒂Rs�� ��������cα�u��^�63$�*5]%՝��HM{Q]:��q�5 ���`9)LS�-��*gL{�x�ҷ��:��rU���\oT0���t����鬷����ox%u�%��[�w"��Ed%�6e�f�u�u�������ݼl) �5��xGRdb�4�z-�+�:�o��*;Yx�i|�Pݩcb��Ft�=������e��Qt1��+�����a���
_q�sgo]�ܪI^�&�����9��Z�ˤ��	��.Zj���-Z��������\y�W(�΢]:x�l7� �3�ۚWjCu�6�L� ��.��$�/ncW��'�4Bʘ�Mh��\{�5x�%2��v��+>-���P�P��܋����S�>bVwY�J�{�]��{�H�jn�C:�m���9jT!5�3���{��?i�ɻԛ^R���)9��r^w1������.$�x��mS�8�Lf���G���`]9�3Fɵ�)�ͦt�]��9��蒅�r�m��/+!�2
��A+�N�n��lm�U|m�r�����}I��7G%��8+6���٩d9`��h�t��o����?
ͷ��3��Y��ej��u����2V�A���˄&�EGyx�^P2b�s8-�3*3���N�źdY���vAS�a�CRqZ+u]���O�Ѹx�%փ���̨S�%D��]��-���l�3L���;:I�"��9�<#����гi�5���T��T�V�������b�P!F����G�v�X�Iz�!ً��ֶv}���� �t������1�!V�����+}81sV>`n��+����\����* 
aKt�v�:�֭PZO�ldRID���p�IP���9+2WK�5����h�@��:{fV��h��N��n��h� ���T�8�#Y��.\D�0�U�f�<O�'����Z���{0=��v��JS
*��\�|*�CS)��E<(V��*�"��:��Jl��wr��6�:0�[f��In�j��kqʰ[9#(��ƪ��i�f_7�Q�}�1n�5~�ջ��檋mjQ�,k*"��̶
��ڔaZ-�Yb��-���,r�2ڕ�
�Bڢ"��PaUl����E
�q�*P�`����Q-�hʍmjŴYTjZ���F�����Yjڍ0rcj����Z�ڊ������%�6*ePiAC+j��-�Q�1�bZX-QiaX��mD��JŨ�*��QF�J�h�T��B�cU(�R�Ÿ��\�V��
�%J��V�֫T�U����X��U[cmm*�mj����R�-qL���J�R�iW���*,E,��Z���UB��Z�hڵ�,E��fR�APR�j�+V��h�Ʃ���h�k�Z���c�1�U(5(��F-s0ŕ�iZ[m��8aTJ�����6��J��\0���s���~�x��7�{y[�SUʼo�����K��i�ip���'2&��M*����3Zr�j6���#�i���۽ن&�k�B�Z����`�Ҩח풝��˫w�C�BX���S���_&�!f��Q>�N���)ҡ|�(j���v�����4��xb�W$[\V;ğ���M�ږ��k���}G\Fc���F%1�s��&y�e��n���]ʦ��rZv���\	�#�������5i��M���69��oF�2�^t�sb���|��q:6�k�;����N+5�;��Q.�,�8^��ևk�k���}]E��=�٦�y1/ŷC���Ƿ�n�~����A�/,�W� �Oah���������}�K�+�4$�9|���fS�:��#����j!��T^�jH�u'�U��m��Z��vṗ��j��u����T�}l���%=C�-����(g>�:y�Żw��01�9�g.}�����\n:Ȫ���)_�p�\�%m<�i=��+�e�9$��9^��s.����J�J�xp��uZk6NWM�|Ap1�n�*Xհ�[�G���E.��<.vЀ�+y��}+���f	ў�݁����m��|Km�Cm�s7E7O6u���ܲv��a*ܶ�ؚ���ټx ^�Qzu4�j�s�;}�g��O9l�_��������)�N���s[7a���tޅ��}:<��E��x5�����'Z���u+Ԋ��p7�����(�/sx���˅z��>F7�y�
��PƱ�mԝ��9}������i#���D��5>�����]J}��m���Xᗶ��L[�؋ns���{!@�sw\�NueM�}[@C�u��h��#6.zc\v7��0�b�x�Ru��ɵ����IMH��.L��A_j��{�\S�,��솜� q��/�9j�!һ�E��悳i!V��z�\�OCՃBu�a���È�p:���o�'}s�xWh+�um�F��c҉�k��gS���(�>��@+2K�8� ��K�:�r]t��8�·#�OxCKv�^M<�<a���E�4C�܅ѱ�]�ݧiڄ�p�5דզ�p�j�4��d-Y���d��dg�F��24�e��ǵX��c�e�P�_�;⬹0Wn$��b�8:ۼ�vS�lR!�}5=�:޹��Β%O�l�=���n����LuJ���r�*ͤ����ݳ��/�Sۨ�:�2���XW�5�m���Mw:7�����,�˩�]�q%D*{Y��15��r���R�Ԟ��n�9B*��i��?wcw������[�2��z�*�D��cl�u.N&I��y�Z��������M��Y��f���b�҅Q}L�@MVFSt��w<�$�os
���Sz���9�=:/��i��M(p��8k��㖙�{�R�\fw�:_�UDL��]p�N�Oq�hg6C脩����j;O�ꎺ���27V5d��g_.�{��[���˻���Ӂ��-���m�]7����͇rЍ*gmq.��UN�|購5�ȗ]��]Ĵ5�R���M�~Uef7U���OH9=�57\^�LlO5�S�����A��s�m��WQgp���_�7�a��.b^�O �d����;OO]v�'���l�I�aJ��W!go,���2�X�꛽��
�vBd��)U�)�'B�+7k��(w$����ޤ�Ow�e����U:��|'I=X:Jl!r]*�w��*��Xu�2j�>ȷ�<�Z^ni,3�����w,��n�ǜԽ�g^�ܬT�u)wm��aHimTfhe-=V�����b�[cV��Ÿu	ջ�8�����sQ[���2� Z1C����7k9)�<���ݷң��N�����2ׅuxg-c��bm��k{xC~����������d��vE(��q�"u���s֎n>�gjW�"�:nQSr��k3*Kq�5T�ͬ!��';�+�X�H�5��JY;*�N+>�)�j��k\y�^�[��f�����v��{-�6�ښ/4O;�����g��V@F5[��%�f�e�Ը�ib�w~t�j��p�~.1����Xd-���,�竔,���Ro=Sn�6��ՙm��Nx�G=R砪�SJ�P�w�τc�mq�Lncg�r#���7�k�SЫ�  F���LA�J��+��T��ᴺ�g5���i;���1���Ns�,�����+a�0�R
<�˩��ﲯ�А@�+�������}R(�:�3���������.:x�gv1,B�o3�k�g��;n�t�]�):���v�j�s;�������Ϣr-�Χ�ר����Z�x{����' w ���W��N�x�b�D.���O `m��n���U����R�Д�:�@���B�Ԥ�qo����oF~��zP��&4j;���=�����:K��t�V���2��=����Q�8��5Y����p�7V�:�{�w!O*�k#�5G:o�G��t�]B'K�g�_Ot4Nػ�.���}��{*�V�f��;�8��vMg������5MY����E�X��UbF�,�f:�[9�1[�q<��z�������t��MP�rޠV��Gt��-<�P�t� �3�]��oC�G��=:;ϼ�w�U�O��-���p�ү��.2��[�7s��y7�GvE�X�$��8����e�CV*K_��<�<���y�u݉n`��>4Y� �Y���QWA����f�Wb�gX��H#��޽��#�/LͽO2o���is�lQ���,�íc�36�7����ݓ���j��Q�1S7�r��]�#�F*��f�n���H��%��H�ÊRWKO�_nn^!f���f'T�QY7uԯM`ӓ�w�lI��������qo�5�a�wn�kf�5��Z�t�_C�ԱjD^j�|W8��Z��=h����#�+�Aغ��Ժ��J�rj�>Q���W��
j:����ޤ��C���N���7��:����`��Ie:���jV�4�E��4kd���r������W\X5oJ�Z��ɍ�M�\L��6��&,;ֺ�o=/z��N��Ʈ{� �nO Fţ:ԍ�B��2�QŚ�tW9�=�t,�z���^�w�(Ȇ��YN�p6rUY�x�C��n6�����ڒO��ƚ���6�ީ�x�sZ�+����wB�����7^]�E��j;q��Zj�\�f���ET�ʻ}�Ҍ�[�K�+#��J��@�v.�E�{�S,����ى��sFᨼ�q��>��ƃ��Ӟ{�5Iz�*�_V;��Hꡂn�]�l�9�K����h]�n�
��T�܉Ȇ_7�Y�����%�#s����t�]� '-��/v麍*ف���zW;ij���M�S���0�=x��.R�N�9��sZ�Х'�����èq�,���5�f�j�U�[�Ջ�V��ֳ���>�Jmfd8i�/�(�G%�#]���2�{��}��B�E���j[	u��+�o2��&�1��P]�P]�W�����Vbw�z��wיL�f��aT�x4�n^M<"zxڝ9�K2��������z7���w���.���qo�Yf-����s��,����r0FE���%�)m<_=�>S���)�r��z�t�}��>t�m�뻾��r�Բ�.�e.~Uۻ��s�v�0���BC5�ɣ��]n��G:9#Sǒ�b�8�M���g6Lu$'_N��<}�T_S��9]�sf������[g��Ყ;W�o�y�rUp�q4�D�_����+������T]����ym�����θnܕM�3�wf[Hgl���Z�I;�r�7eU*<B�P$��h�7X���S�r��9\�/�!�m.;LF�;���X�v�.�W��S�o*[N�W:�K��r�of>O�!�b���uk2/��n��r�_}�e�<�9����9v�frw�#��<[<���m�I6���WV�������v�:���gu6wkR��7�f�������-*���4g6Ѫ�UO=:���w���j��lԹ���;�_F��(�մ�^�J�~D � b�>�ŕ�<���D��NT�I ��R~���wK���槰RgFr�|�{���T���r��-��T����`�����Ůq΋�\�v�q�52����}kk����o۳ݽr�s��Q{^���w�W��7�T[���JN��r�oBu#ayu�CjjK���w����s|C��4��v���S1��qm�|�Ak�5��3��bYqY��9��
L_ڱ���z����z�Ł�[�N-^Mv'O�V�Ñ8�r��VK�>����5���K;��Z�]�)�n_J[��҇�'�)� ���b��L{,r����T�Ъ�:�\2�����Nޛ9�ji�L�Y(��������=�5I��	�=�)[�ef�j֕�W33�ik�w�W:G�t����κ���pI�9و��h��w�M>�@��i����nuuuu�z�Z_VCz+f�
�kn6ˬ����H+y�uL�r(�+9bT�1���ZN���܆���	,f�b�9;��m�䦱�ǚ��q��B䣥7�ҭ�ݻ����W�����Mf�4�q��V��}���mZ�i���@޴�G��b�>m���ԧzC���܉Y�P�>��̇�w�u��	)��>��a|�i;���y�.&��dn�����v��&!��w*���S�f��/Q6�Y�Lh���ZV�[�'�����Z�ګ׊�"���)gK����	�cE܏�Lk���5[��^u�����uo���{��D�v76��t����|�+������}t}Z��PQ���e�01˯���ԖŦ��9/+�MR���Tb�1�yZ�J�
�,�Cd+.KS�cɓ�gy��K��c��VFi8ٌ���S���t��}	�1'9M	�wn��
,x%zQˏ�G[��	<�6e�ȡ8>��]Te��w�}ry�+����]�ԓ�}BȗYաQEU�m����WW6`�o
s3h���2Tŵf:���S�޹f�������Y:z�����{2d��<ɡ�gR�����\{�����U�
��@|��&���n�(�ؽ��FDZ��,��?.��z�4��������⾩����N��k���Ei�f��y����Z���k��B���Q����>��z$WnU��rVp���tq��eF�Y���q�]�a��_^M�'����w`9��yn�,�]��c�g`��k��qm�F������f�7y�oxM���DcҌ�rjOrV�g��i�k�W�h֔t���p�1wb���܎���64�IuOK��7.:x�x�%ë�����E.F,�~T��v�1q�zE���;o��FN�|��aOW�=� �EӯZB���+#���M^�W*�Ջ'mkӱώ>C�z<1
�(1�����i_�t30Aׅ��}nK�iB�{����5�|7�ؘθ�V�-����>��)'����ä�<{7bbHN��j�C���P!2�n���_�{�K�oδq��*]��rAY-ъ���f!�s>k/��pYD��t�=��T�V�UӫeҦr��s �rX|4��v�qGDs:�c�b,��:v�q�79G�K��y�*����LQ��**T��L�_�r�Jښ���S�+Z���d��U�[T�%��;o��Hm#J�3�AݠR�XzI��ܶ#�o��/LW���k��뵸�|����L�\���:n�9eFx[I*`1�v�tf�ރ��3,�ȿ����л ��V�e��[����1�N� �z�жK��k�V����ut�Q���4.��v������F���j���kh�ΰ�1gS{����u���v8*;��)F�c��u��6��x��T"�!�O���,���(�ht�<�t��Bx��Wm� `����g`Ʊ�Q{�5}pnm$������ht�n�	w�ȂW:��v�k��L�o�V��Oi#��/��>�R�Fg`���fZ0n�"/��ݕ}z[&���1��v�dӹN3�������j�?L��h��9RW�M��g�z�&������tJ�b�+xV�u���j�U�TK���H`��Tx�V整JJ��x���":T,�y ���9����E�w�e4��z�����#�"vb��� =e��\���t�4J}o�,5Y7oqt{S�@�}u}���L�]�_l��;u����t�(qs�R:7�]��R���Œ�i�:�yݱ(N�,���٣,	��S�2 +���k���c�vm�K"9f	���+����a�o^qu���xkKԑW�<W����me�S.y̦LВͳ�,�f7|ܝ�(/${�-�/�X���/y�vD���[`��Tc����Ht7'Y��J>V�V�N}7c�&儷Mn�Ǳ�;��ƞ���m��wQk�[���oF"��ZYb�.��n�☤�4hu#���i:IĒL�kK��M�S�<���F� �%��y��K6�S�m�G9���$k�p��b�R0�;��	�	����p�B�`��U�1��e�8��J"i���ʯS͖��m�n�Q�y/���᎕:�ܧj���n``ލ��V��mT�]k��.x��w������]bҋ)��m�,�v8i�D1�l.\xw�w���I\��7[I����Z耬kŌ��EB�U&��B�A[�3����s1�5}&��(Yd&ȧt%��5��>�����mF`��v;)�q�+�r5�-uyE1X;���R�F%V�l��t�t����6n�1u���}tz��u)��h��j0ܦҀ�n�3���T�۴x�X�wpY!��!�n�E��.[����Y+j�j*�BҪ�ʣX5h�ZV,JԵ�JQ���)e��FЪ+Z6�4m���Z�J�q��(�Z�iJ�+�`ʔ[UZ���2�iKX։UU
��,�T�EV�-��-��Pj[h�m*9J�G*�-+aZ�FUeV�1Ċ��%k��ZR�h)X�VV����P1-�J%KmjV�T*ULʹj�%Eb���lE*�6��ԩhT-��[Dh��,m�+���el�kb�2��U��EB����b��m�Z[
���TjU*)-�b£Uj���e-)l*��DeUKiATUTX,DҊ�����U-V�Z�JJR�5
1�l��*��Z-�eK-�T�Ѷڍ���jѨ(H"	D J!VWH����5�s��ie���d`#)�=Wagr��5g31�{%�c(T�WN�ew$�a1�b���|���,���k���9�j㕺c,�[1)Z���J��O���(�Ξ0n�$Z�r��q�T<g�Pձ�������R�o�9����B]o4 f��8=ӻ~^��b`\.�%��C�c��<5^_�[˄���]0�V��|���	Ned#�s!��$ƺ�Vb1Q���FZ���o6�(v�`�[�[M��{C�#�#y�*ƹ�V��}u����$��skrn̮}�*��Yr�7��{;�ӠvN0V����)w�L����[W�Z��>w��w1M����,f�/v�ͬ��7����j`,s�L�w'����+rݘ�ݺr�Zw �1ʺ���w�j�l54�=0��4,�R��9/�H*Ci�o�ch+1���֬
�qo���1m�I��#8��3ᕢY�	^m[��T^*��I�����������=<����Mz�$v�4����'�t�ɗ�����c�ۣ����r��{DغquA�6	b_f���ط�f)�������\:�$�w"��;61��ȩġD��G��Ƃ���Y�p ��O�M�,�=�KR�����x�I��<�ޮ�����
e}㭇����Kz�p��g�&a�_H&�Q�X�z�-�҇O^��<�kk���u��u.�׹M�0��������/�h��֧<�oe�a�J���DR���[���{|s�U�T�Ԭ�J�.�Wn�ᤚ��^�n܇Ŝ
�U�a���ڔ�C��f6�Z�WtN"c_%��ם�Q��
���8��`��/J��)��f!Kpb���]�.]�/�ޒo�����b4�jw�hZ��{�/��TA�@��U�qY2�RrsK*��跗۫o��$�'q���[j��SE�@w6��ۮ1T�f#P�<9=NDiK,ӿW]�g36+��/��e�,j;~��hf��6����dק:�ge�a^��}#@uW�Lp��rG8�n)1���U�|M����=�#�q��Y]�*��G/�:��Y8V��O��z'��Hɲ�w��b:�j�	��x �{F4 -CP�2jƢF�p�7����7�^���"�F����E^j��;O$������Ū��e�C��]�rT����XP"��먷/FƪjC��-ѽ�v^�Ɵk�ߌS���]YC�x9�s75нӳV);f��1?k���Qn����Q�$v�z�/h����v�)KM�����,ߩM��5��3����5v�܇
��^�us͵J�4�=[�{o&�V'K��ؼG=XS�偘���ɋ�Y�;���\L$����}�����GR�أ{4��a^����R�U�d��I��y�������*{���K�w�w��20}1vu��{�@8���+�ϜS�@�q��\g4`u&�S�ۻ���r]�p�nTodT���L���iC��R>���~��Z��{��It魙���r����n^֌w�����Kp�>j��F!e�xM�]2����f������V8��U�vJ��>�Cb��4�ƺ�Q1�fd7
��qM�j͊���.�ia[�:OV_v+�n7���+*���d�&7eZ��VZ��kF�t�7Avh`u��:ɺ�֌�)]vb�����n�;!�����7X�����l�ޮ�]1�����Y�����u��ۏ�b�[�;7�ղ�&���_��Ox��?*t\pX�r �%�<��+����Jb�^��զ if;��e�SL����uc��mL��5U@�Ut�����S�2�qQ��F*�-c��� 7��T�@��bP�#W��v�E��=|f��t���^�N��ֲk��J91�eL`ۤ �\NݎR��^�N����\�&��n/�E<�Qѿ]eS�<�wb��x=�V��H}6��q�*4<��W�>��䪕�ZL5�*o�;�,�軺�O,Ѫ����ȐU����1k���i���<�Im��)nw��{%a���f�-�釷�Fh�>s���:���D�ݦ���F����k�u��,�ŷ����:Y���6��P��5�Y��q%Du=�Ȼi1<��p�kH���!�e�w�ǲ!��Gt�yI���P
�y����yo�W"��Z�r&̈�Ɲ�	�u�TKj�Yv�NB�a���(wu���#]5^��R\�[VZ��iyе��n�5խv.ĥJ/C�'[��ք��%wS_oô-���3R�wWC�
2۽q=���t�/���z��f`��u|�i
�����#����Ho��dV�Ϛ�ɾ�>��_{0o:��ؾ3J�e!u�:�CL$�-_[��\�v�%6�޶���@��#Ա��'ˊ������imN_j��&�]��i�[�O!��on&3���qÐ=����+���縵�)ͧK]��U굴����뢟-z-���^����8z3�yY:�v��ËhT(�F�8]N��OR�{���~���
�����Al<r���M���Pe�F!P3����F]�9�o�+;F�B�^^_rt��ő��䝎09*��#a�Fb�TZy�k'X����/a������[������ׂM���8ÖU�k���U��<|mo�6�fױ{��<�����O&�ՔR9.�8�w�5���3Ր	N�G��j��=�������ȇ$,3�^�z���\�]6l���$���fb��@�����:�b�\��ՂuKy�����1��E�}��m݌QZ�:]]�y�{{j�[��Ru5"!R�����q�ʻ�Ϩ���]��[�#:\���
�㇌E�[��*\⣓�a�m{״m�֦�;{Ңx�58�v}9�kˌK��
z/���֒��[���������_"�ߓ�{*�ryE���D�\�1�ž�L�Z��0E�<X�[���o#J��]��ד�w�Q���^�L��EAz�%��%i�d]�uٷ��+/���YYk�V���ߚ���ڥ��q�#.o
������O����z�)[�8��j��}��9;�[�����d��fc;�5O�ǳ���k��1Qm��M@g�j���r�x�OB��u�m��<�;]h���W5pk��&3,��ͤ�Ov5s����ݐ9���⻞}��*�t"�ַ��zq|��;��;�1�lX�v-Y�ӳv�=�sj�Z
Cli�l�b�qY.�ui����w�����W#T1J�*��k���2:pѡ���K�8��ᓀ{��ç����qn>��{$JvS��8�2��e�{�}2�j��A�	ċ�I̦�us�l�9���hKWI�yuT��\����Ν2�n�nD��^I4Ri�ɬv<�\���3�k�:�N]'wGx�݉w�ʌ���+�1T;����[�y9{w��Gu��W�r�\6���z�G͐��1'UW��"�t�ӑkp��s�B+��+.�������e�/cQ����/ZǪs����zj\�����'~����^ߺJ�ɍ0�e�K�뇈�pd=~W�7��n�^�*z��WUS�-�d�q��o2B짂��j�*�'���	{W���}k{f'�V;Ys�v�܇-hm��[ʹU� ��O6�z�s���o+ݠ��P���X��}��_%�����)`6���Kd�J����˹F�e�Vv]���(�ݞ*wLxf�.j���7���p�x���l:u[W~T�w!�^�ZͲik��o4W��y�7�2@���������-6�G�����M߽2d��V�E�**��P#����lsk��*I�v����1r�[��S��l
=zVv�p�^F`��e�hۄ�-�Z9q��x���v���m�c7ctU��:Z�6��h9��*����+W�5l��]a�{�M٫�c�A�b��2�%�9N�hJޖ+GJ�z_E�*-4`q\�w��_�u���k2G9��M�gd�o%w��U�p��+�Pv/�S��WW���\�]�or`+N�e�1>������_�9��*x(ޞ�}�je��kj�v�=r/f$�pn1sܖ�g8��J��;��;��{بBa�~���F*��\ѝ�I`�p���7=(�|Z��}��-ힳ��z0;�c�(#1S���j�nf9B���)[B�S��c
����v7���]KN���n<,)�ч.ȱ�v�Vf����#-��u��i�GM:L�N6h^2&>�Z�¡ǥ��S�}""o���]j<-��+�
�����Xb�gj�ֶ�����u\���f]�u@�5V����.#1�-�͊�l�WEU��KZ�ͱOwb�� �>�j�^�Fz���Fo�^�6#�}��(YW��Y��w�ѵ/�*.�*����B+�Q����V�QW
�:�+�ox�afY�KjY������pò+8���3zT��{���SRr�׼��mڳ@ؼ�(NMq[R�`m4���5�[-j�2Ҷ���t�J錮��l��^��ԷN3n�}���8�iX}�[緒�����lWԱ�A{������3�~̦r^��f��e���f���3�y	�q�h�Y�5��6w[�P�YȬ.�F;4��oE��v7w�h��U������e�ʩVR��4�bl�Σ�v0�&'���:��j��5�N]�F�Cӱկw"[=p�6���P��Ť254�mobH=3Q�d��z�]���=KRW-�܆uIU�m��6/�҄�%�.��5o8�V�� 㷑��'~��cK�D3�L$P�=�lW�C���_�m��:jt�Q��m��.U���jA��;7cxo
�Ҽ��<����a���\���U����Ո�O�׹/���IE��%8M#�qs�N�#mUF_\3�b���׎zc<�iؼX��U�n�.8��|:�:��,�C���e,Q�k��d�h����
��qa��윪[�	-�D�u�~t��jơ +�9�����nS���]\��q4�H�I�U��S:��ܫ�o��7k�T��)�c؟f<������e`[�gxu�trU�\v�j�c�!��]��|�2}v���W��ĳ�o"�����	mM'���U���#��.X��W֩vZ�eR�e[�ާ��j�m�;�)R�U�˵��Im:���/&�;�i�P8�Ǔ�	�ti�3[X�@WZ��q���\��q-�~F��5��N�S���9���ǔ�[���Ԝ�̩�Nj0�t_8�d-۬��&�<ç]�Wm�ĕr��3��>�vkˌ�^�p���j�*��P��E�u�xn�nRx�&��,O1����f��qYZ���ŷ���{"oZ��;��'��[;������w�b�M\�7�	x�N�d��|sD���7�Eы���+f�b���Kg����.�k�}^���
����/o/_,���El(�B��9�\�U�w.�*K����|����;��BB��d��	'��BB��$��	%�$��HH@�nHH@�����$��BB���BB�����	'��$ I?�	!I�!!Id��	'����$��IO���$��IO�H@�p$�	'��$��	O�����)����o�]���0(���1&�&^���I��ն�f[V+e�Ym�i�R����h�d��l���MY��KVf���&��M�5���T�b�FkVխS#V�SK6j�љPĭ���+ZB��e�d_pp�0�jX����i$�m�$�����2ѳ5i�;k���v�FY�%l*��ٳMc۝T��ӫk������k0�m5)�����d���m�ի*�V[!���F�ͦ��v��Tm�j�X��mA��cm��ji�[2����Vf���ԙ�Y�ܶ��R��Z՞   6��� ���{��{WZ�c�r]�ZNn�n�S:��g]����zuyQ��v�v��*��XݠηU��BwJ����;�v�s�u�[t�x��e^�N�  [|  w'��ֻ�V��w{�mvtsw���=k�Kvݳ��mv�֐��u��OY��ڻ�N�I6=*��=k�׫n��r���*�������m��gj�����ګm�n��m�kmZ�m������S�  ρ�����[�n�t�f�,�wi��u̬�s��]�m�[n{\�m�^�֮�w�y��n�n=�z]�wS�Y�7��
= hP��Wp�
 � P��{OxP�B�
 �=��kof�-V� hd�J�   ���(P�@�=��(P�B���w�w}�
B�=���C�Сޞ��*�.힗{��r�M��K�6�uw^��������u�u���.f��ĺ�-]��n��h��ͩ�� �G�  ����ת⊣�O{�WkG�j[�� :�u�+Os���XZ=�Nz	�w���*������Exz�V��p�m������m6��V�fefO�  ��%U}V"�)Df�������5֪��o5��
�{�zz�{���v�1ly��֔�U��=z5ε'���i���P ��>   ���T*���S�N��Q�{��U *ꚫ��J6��ށ�,�]Pm��=5�j�k��vUz�G�Yǫ,;�ř�ͺ��ٵfc_   ����P���◷d�w���V�vGm+�Owr��]e5[�v�2j̵�*��wX��ʻ�p���[ǝT+��nW�f�T�NpTu�e�q�yUH�0ՠ���J��  ;�>;m��\ׯ/m{�j鬸lݶ���gu'���m�n���;f�n����ZuJ�t���Sڹ���^ݯt�Nج��]޶ۛ��-æݺ4t������i�nS�ѐ�
$|  no����wn�kں����Ikg/6ἶ�5S{�Ǘ-];�ѹ�m۬�n��͍%rkouOs�e�N�kk�^<�5t��{�[ҽ�.�mw�ʏ*���]� 56�ʒ� 2 S�0��� h�LSUH�d  O��$@@T�Bf��� h �I6U)OSb2x�����~�����s���O=�n�i�]=��Yn��+!!����E���I�֫Fꨒ$��N}��IO �BC� IO���$��IF ����Xh����������đj��!�V����2�B7���(�:��û�hT/f�ա�� �+�ۓ��md��^�+!	v+��fLݠ��N�"�����P�R�ŨwbѲ�nJ�[�T���n�0FQ�R2�3C���d�5vvŭr�����x��^�y�x-�������G�.h�ƦÓ��/^�*;x�jn�� ���I�F�c�7	�O�>F�b�j=ah�PhU��F�k���Xs#A˦Y4�)��U�'S���2�j\�LT7���}�����_�ۛX�S��S:�j3 �ش܅�Jm]�bBj�n��U�(B���j�VDkZXQ,��h����Ly�Z�+s6�ڿ�[a��EE�<M���uf�8��#b��J�.��������r�y�rcN�m���j����uKD;Ywۯ~�h��\%O'N@�����a�٭zp�s\���J�����;W��b�S��(R�r�_ͬ��e�kVI[X�sU�ơ��D-��w)9@��m���Wp�A�Z�*n
W�)����}�ꙒQ�4�
��̦a�CB�p��u�B�=QlV)5����٠��0[Jۘ���Җҿ �7!�B�>��J��\�nG��8����+�js'�è6Fe+b4�=т{���lL8��¤�KU��ԫ�Y��E��A��G`N|�4��[6�<�L�.�� �!��d����C��b�Gr�۔��g�lT�Z��d��5z�!FR92�9��{Ӭr1+1P�U�f�Qaón�ѵw���o\�D^+ٰb�6+U�&:��M�B��n�*����w)���~���E m,a�w��3}�b8$�-�U���Q��#�>�u�ڸ(��%�F��Rd�l�)��rk��l�!�^�2�Y��e�;4!FE|�{�⹹�5�}�n�n��[�
	��u�-I�5}�fMr[ܬ��J%h��
qY`ԏJK7*�4�)�X���f��HccC���l�{je藡%����[O�l���8ܘF��Ec"&�Ȏx�n ɱ�H�Dj���ޔ�ѷ����3���H9����ҵ�ſ]h;�J0�Q&`L7���d��EnVݼN���s�4.f9WYZ�v�ֺ�X�CK��g�n�L˦��xQ&G�h&����M�z�����ՙr�$����%�î�*�ެ�E ��(^I�����P?8��-Y�"	m�L�� ��"��Ugv^7��㢊���)����娯�� [V�"��ݥ��C�n��T�<Ԫ'SɈ���)�z��[Yr��5�"���Bk9M�N��5��L����0,�0(K�.3��O%�x�w�(Y ј�A�vL��En8p�1DQ��M ]���F�=k�j�p#�KD�y�O)G&Oێ��`��M�'�e�V[e�Vv��-��*�sv���ݙe�ː�)x�m	a.�i,����F��)MF �m0.Ր�i�e���-�k4kh����ۺZ���:{~�s{mLe͐�HpʅՁ|�h��n��2�I��<�-TA������a;Ʌ�*;�h0�'��r���HT�E�D3�z ���鹾y8�5��r��U6�ܙ�#2͹���}�l���D�q�D��Ğdh(�7l1t@b�U�>!�y 1]���Ơ���n��w��٬m^ӳ6��5%��=�l��3NÅ����D�[փ��<4��d�j}7Ҧ^˰�ǃ�U����PmC	j8)�e�z*�4�b��ɴ�/i�t�S&� ܥ�Y�І��KS�U�-eP�MS������nOMU�����wI�"�� ڇR͂�d'lfV�Zm˖�7�0 ֢j��l@ܨ!�����*��8"x!�y�kr ܙ��5�ه ��x�􀽲@���kx��Ǎ#Q|�PZ�[6��Ǒ�Q��@V�ƚ��L�kGV���5��Ȧ3��D�����؁Cp\&ODn�w6�`;�M=ip"ڊ)w��ExJ�@�:N�8Ɲ�
zN�+b �'�KPnͺ�Ն�R�3r%�znW5�L��H{j��.��i�*X[[���ȥ�˚��E��2���7+X�+�Rb�:�7W��{��f�IJ{�|3-�,��Y�����dڌ'8Pǣ��4Ԑ�@J��b������cy��y��\����l�/��@VPf��L���_bO#���z�DPɷ���L-V킙�m��뀻0(6 I��fS�6�Õ:�ڕє�cgVO��d"�ɲ\���VЙ`��|p��É8����A�r�T�~�4�k�C%�&T���\q$	:��8�	�4�:Y�%����������E��2�ؖ ���d����*�
�X����w� ي�F�ﲕ�V�J�.�d�K�ĈLg���co�j���F��}@(��t'���In�V�0:��(�z�c�n���腏E�c\��J�F�]n�&�jBѺh���IQ;�}Q�S�Q&�u��:�W71V���⽘��E��-�1��VQB	�i�tɭ�P�itt;�iGv��olE^�Zq��T��r�!DD�Sw5Q�ܢ<k<^K��7ڍ�L!�b��+�N=2T��cF�V��T�HinP�O��H&��x1�aJ��\���8�ջ���1�d��d�L۞���`��y��.8=*󍡱��}�e�ne� �M��*��l��9���b«"u"'0T��I�B��W� �yefv+����a�ߞ1�q�f6kU`v9�m��kK�7V�>����vT�^e+��۫�U%���Wr˒��YZ^i[��wb�j�n���f�1rn�ú_4��"��(4��pJf�g2Z���<Ҧ[�FJa�����J�Y1���'�[@dW�_Z�<����A!�(�ʖ��k�9�x ~���0�63��/aUڀ`ȩ���)M�½t��n��7{G���!v3Bֱ	�)��	�KTh�򈪣sK�5=e�9j�o/L�#��:���I¯�JO�6�r����b(
���z%X�X�3���؎ލ��4����P��L�orc*Ғ�+��%D�lr�̑�N��2�л��6@�R�-��H��n�)��r�/�&�V�^1n�4B�v�	X��Y.Q�-�YF��P�����n1��@�Iy��i�l���;R|u�7��A�J-"�������^"��( ��k`wtQZ1eӨ~�[�Z]r�-Q�[��)��d�V�9u��j�/,P��,ޢ��[�5�H-�F52����.A$2�r�ʔ!��a'^���<���=��<�Q�����cfn�6=�Z#N��t4Ӕ7Z�J��M;�.��ұK	N�m|&�5�e�L����!2�e
N����-5�ȯN7bh���o3���6	��0��E1φmz��N�U�f����������0e6Ag �K$�;�v��eD�)���N�����dD�T0=�W������
KX��̬I%I`��p1��9"V�[�P����*-Y2Cr�M)!o
WA�«KҦ���&�{��]Q4�D:[�(96nK� ~�ց��k�reK]hbT���؟�DY	xT�n]#�Bgl�Q�g3VM�t2�LGyUӇ�)��u[M4��5��K��!�Z5�ͤ� �Z�dn�c6-:7�^Qdp3�7��k��u���ͨ
����V�!�p\W6��2�ݪq�6Ž�l��͛-�݉hj˭g(���m�w,���g>�oA�0�q�߂2�LҨ6�6�Ve��<j_�����r�=�^;�`k4�BfnR[7��ԵřWN��62�ϋ �Br�dm��a��/c���^[��u�R���oZC�:4�u&f�0JE�z��f�5�I;Y��am�f��,��Z��$057n�1f\�E~b`�sN�Kk�su���ܷl�u��Y�)x����0Mh,���S4��h\�H����O���ō�J�n�*��1Gt�7*X-���SQ-���>�ͬX��ܣ���̴���]a�*֙oP
;BQkL�4FS�ݒe�V�V*�f�Zi�y&���o��ǒݐ_+�c�TK
E�Xm�ǓEC�]��.�A'f؍��<�[����;��I�{2� 
W�֣=�������Е�Y&���*��ar�# �X�H�/�$�r�fȩ|A8���!�suY�"P(���=�t;	��wwQ�_���O�@c��7)5�ؓ�a�O<SCkkU0�����ͼ�������I�H�,�� e���7hI��S#P�wmF7V /
� �p��Cji�E�gf��eE���$^�;O`��w��K*3�oc�I��k�����`�8��w\�>S�v����"�;]kJ�vѯ��Q��w-K����֮rđ䚜Ê���2ު��n�MJӛ4�>vfܭ�t6*��5n����i��ֵ��D�\�$�%Y_+k,2|���&KұH%���[z��ԩ���GCq�(�t��R��9E�K, �����[5�i���i��*�Fލq:z�e��H�C�X1�v��ew$�K��<}�iyp�g�ey��AP���-��u����(v���32�5�rə�I��Z4��]ǈm֗t���T�Rgwl����b��C�aŕ% �EL�>z�V^h`!4�rT+nk�7@ɄY��QPlDp#�e@1�����x7��yd��۳�`�;���:̢�˴csi�2m�b�;���h8�o7T#�WZ̸4< :4�,�1
��|5��Xb{L+
�e���[���
���m���,�Z�!���Ɛp�b��F�+aVn����9he$��:���D���-�ѲBOc��Cod#,���DT#+#
�٣4�7^�Y�@T��^)ز2�V{mǓ-s7)���`�p�!�E cz��[������.j��ۻ�L��Pp�&����1���aɁ	(l�d�5�'bp��%m]��wr�	#�n�k6�^��k��j�
T�(�Gj"1�ۏ6P�-ōQ h�Ͷ5��ۺPD�zkp� \Ty{u�F���!��,r�,I3â\�k*�l`Upl@�/q"���9%>��f�$�YM����E��^�W&̻<wd�^����!�C���.H����К �:n�еa#��	+N��Ԇ��**%n�b��r�V��eDo�Z�U���X+\�rj�i:5�;�]��^�����g4�*�6
�TT1dXTd�skeI6ͧ�-��{W�;�JH=��Źv��3�Z��ELfT��6��P�[���K-�����+tp����A爵��	�r��لo����f�&��&:�y�1-����X�n�2�a�&�J���K ���;n��:)�]j#[�!�Q5ѹ(=�n��q�kh��e�J�F&�P�����j�$�c���a�U��T"SW�`�{��IP����^�'
�<r� It�@�+fZ�pS�5�v�Z4s�t��S4����=KEh��4���5�Φ��.>o�㶈�ž=�2���P �@���+�UGujDO}��� �Ǳ�n)ShiaeeЁ�Z���e0r�ܹ�E#��+(�X���<;N)6Ƨ��D�VsssY:D��˨�cv�ZL2k� !Ǹi�2�[қ��p,TF�x�|��a��FԷs7ڴ*Rܵہ:.�1t,i�si��$pdޑX�)��wshbz�,&���<��tnŊov�}є����CF2��I�0f��Y����Uu��l�e@t�[eayDL��Wb�eD$/�V�0$7	#V��{C,3
hC�l�T�76��ܷ��rMR����vT�f0\�	���\)â���R�ۭo��5&�-��%��A3iR�gZ�6e�9�(V��2M�3�x���!���6(�*`�C�ΰ�r���[�\�4�ԭ.h�6�HPcO+÷G��c��8o�r��m���e��Y��n�Щ��n��Y�/0��ߜ-��4A~��T��^��4�lސ�̥UkIce^)J�Z�7幃�z� w$f�H��P4�e������u�X�%+�@n*�*��_��35��p)���Z�O��ɸLS��Sw�*4Q��8�1X�$�f�{Jۙ�{i.u���t�`���(��B7+�����m��0,�����Qe���v���bbV�tE������+S�� �1#�nY5	I?n��p���(���!��&�V��JAD�l�F��P�QcH^���Ҽ�FE��Ƈ��c93@�b��J�V��[(�ڑO�Z��[ ך�7f�ہINX�un&L�
@��b2%�{V�{�b8ݮ�*�1��ɂ�S���k��6*(�:��
�m�H6]�Un�=ֱQB���:l|��71��L��lp�dMt��A^�6�T1��;�Q���6B�9���]�Yj��	F,6[�6�J�f�;�`�[�Ǵ�ELU��%��)�̼�۬��-�d�ʷ"Ҷ�ϞSxe�a���^���$�n�Լ�y�@T�A����1��m��k+f��*����D�P�۴.����#�̻ I"����k*2�e��bց�e\-�G�n�[�k��^C��5�ʚ�i9�[ d9&j.�x��P�m�H9��Ou�x$�d���YϺgK˺���$_Ks����>�SCG�f��c1�G�5-�b�mde#�2U��ꖹ:Y��*K�K�z�/�����9�Ԁ�ܫ�6A�p����t.��w� ���ð1O�Bu����9�ÙUnE(�V����.K*�Q�qix�nY}�v����;K'��c�	���L�����J��z��4�X�z�7]k����	X7s�M����n���HM�W�����E�+hL-��M�9Pͷ��&���"�%��5���W�M@�,!ǳ�"/o��B��g�XϬ��G���OoK�Nۋ|�;�uA��7(qx>un�å�-[͹�N�V��J�TL�ΰ$��yoR3,*V0�9(��ң�X�ۑ�W&vG-����|[�ƃh�ڽ������t�E���P�޾��vm�v��N��Gܵ�銡~���{�0B�����0��&Q�/c�|�`^�j����R��V7 �����j�z���-e3R�kX�[�;�����Yk�p��d�k9:R��c������jc�Th�,j�EGF������oj�;-ey:��	�M�3*>6�Tƀ8*M�]1Ւ]H�'Z�ŗ[Ԝ���P}��������5�wDlA:�imuC����J
ӗGQ�:HM+3�rV:{����tVbJ�Ӗ���xF.�'bw��c�����: $�5�Z�Kص�K��de��M��2V�-,�ЗK(u��=����J�.��Ӯd�}׽������!�ĕӵC���ɔt��> �������1
���Q̦���6K���qZ����{V���99X���\a��屚���y��hwuR����Q��R��xU���]�8LVwi�����Z}�FvA�Qm��t��8 �+�Y_w��->��y�؎A�[;ž�Jݽc�^�M��M�.��^���k�J��Bo(��U���������������N���K��W܂:������_IϺv�(S�*�gj鵭�]�SR�����p��w�A:{R����]
�Ss��^��C{D�����Pإ�;n��ҧk�Ѵ������$�;���=�:�\B�������љKw�:�W�l#�<B�Q�˺9��u�������`�7KZ;P�9��ʵv+H���,�MW�0ԫ����Ԥki�G�*�6���&]��-��NÖ�Ꮒ/��C	��n�=����M��-C�Mos��b
%[f�6��s�!����Tk�38��;�N4�o�}��[`��`��yTXb[.ݎ��R��<"Qbٺ �D�vU�{+PV�]����{"�L@�	X Fd�V�%��#Nu�u9���wwǇ���������f-�Zt��֡���|�`�Z7h�(���N�t������@�����ۍv��o1��l�uz����'����5��=�����=��'�Z���iߧVh�i�s�doW3��@�!ݎ�bh����]ۈ��v�7@��ٟG9��6i@'5�݃@�
��hko�i��o ��_���o1gۛ~7)b���-n�P�`�&x��C�x��>�ݣ�̢>1��k���'
��i�#vWIedU���j��c�s.�.���'�(���2���Ƶ����W����m)M�v	 [(ڠV����r��v�"�Sr.�;�qe�=w �`�^?"�u��4A�KG%�宷H�J'��voU�RQ���WV ���l�����8�iglZTb���6���fujYz[�s��s�V���*�b��'��\0��b�Υ��i����0��m2���%kw�E�,na��*�dʺ��x�����R�9��Ԥ��WU�\L�Cu]�f��ă#�7��`�����`���X65ς���ܙ��ơ[ܘ����v�ū+����t����%t{A�Н�@��R�����j�ebL�߷ȷV#�8��������W=�JK���LrQK�+��8�����P��&Ɔ鄁�}d�iHq�,SE;����}E�*4ٸ���]<��Y���}}�=�Æ��5���/�r���ͺGV�W��x�'`�w�p�8��]������w�uRԤ�x�༼�)FvZ�g7����BK/,��t��R�w��W�ٮ8�'q2�����s���-�hӭ��B@�g�@]�q���6Xٚ�x>ϻ��'���F��m^��M2��:J�E��t����p���^!)<*�
���]N淪۰�3��}|.�j����~�fZ�'�FڭG2��ۯP�n\wKR��P�x��x��V�Z��o.�Q>���m�m�W�G-�];9�v�!E1�(�YG	�[���{Ǫ��zM�s��AQ��zP��k����5XHC�H j����0v�e�y>��8oj��a_U�}���ɒ7=4{@�E�;9c������r�N���r�.I+4
���q-���]�{*t���S=����җYj�ũ㏷�t;XR]e��)=ﶵ��eݗ��0��̔�+KQ���)]��xV��P�@{}��lO��Y�'�5cr����j�(�y\7�΋���ZDD�)m����p�zi�g{�p�$�d�;Ҭ��oi�]�ަ=sw�F�6<���.�@�+0-tE+3it�à����q��RC�N8����7�=p���v�����Ű/J�.����F]�T�ѱ���T.Ƀ{��gm5��F��-���zrX�2��9%��Vop�u�twFs�M�0{k�?�0
��s�v�`��ށ�0�xc�;;�c��pE1���#�i���X��g����<���e��{eS�k��[�-h�5r���9ԮmL��a�FmA5`�emXk��r�@JԎ��<�m5��rU̷�^nD�9��o@�nÜ�91�t�L�J�ս~v'��z`����y�3���-yQŞ콚�]�>��7;�B\|�5ڮ`�M�7�^��q�õ��z�p,ٴY���sF^�:j\e�F&�)��L���:�@�v`���]ۈY�A&�T��n�g����؝�f_d�n{�gQf��a!L�׭]�}�'׆�]�w��*��F��8��	�
ing�Eelg����Z�����J�J�CYݽP�p���Bc/{)�1O��v3�2m��m�����Z����μ��P��C���fMt�C�Ε�B9��J�)b��7�T� ��:JKUI4>��h�熑�ؕD%d�f�q�2���n��Q�R;��o_hxָ	/Eն+v�����kg��<�ܖ�ȁ�5��Z�)�S�׮�X5�-�46B���޻��?9��P�B�K�C,joY���b��������AR�5뛆�5N���ڵ ]�r�^rN�1��y21��=�`-
���B�x�|�t��T��*3[��4��MM�T���ܢ��b��΀6���vC˹Н�jN4���a��5O1������0�gyb��ޗ2��r��8��Z����e�G���F7��\eIW���7Z��h$u],�u!luj˿���|��1�\b*�1�5V�-%��:�v�-9�;�oB�Ox��u�&��V�"=��p��G��l���[���\pܧ|ym����[�8.I˺��XjZ*+�g;�EB���av���+8�.�ַ�	�J���[
�vͥ�+����������a�c���py�F��9z�j���75U�6LR6 'P�_�}��Aח�æUYН�<��V�T�QJ�X��W4kN��,*qh�;��%]Ic�,�v��W���6�J,��142S{������� ר�d��޾%rESon���uxޅ���`{��@����ɽ��8�øb��\ �|���-������L���;U�����yv��.��i�}a��LZ��W�(��ۈ(z�4����oc'���Z�Y�5�@�h�j͞}�l�	���ɀ�M̭2���~gn���PĞqj��އ�-+۬����sgP�K��k�S�U�؄T���9Ai��εZ/0�˦7(��*ͷ����	z+��{���ۄ &�17%��nY[��+ ��>����]@��CLi	�{�ͫ�W�J��_uq�yWK��ʦlقX�O��Nb�'�Ԕ�P؆���WF��:'�|����u�]��#��u]}R�j&�P��*�����\q%_!+������^,�i�N��p��Bn͏N�&v,W�yn������>" ��k��<���'P�͚u9�;����޲s(��_Mu�u������p�C�����,tFQ�CӸ?+NN�5��eθ�jW�T�!�u�j�9������s���n�IE&�d����č�2�=cOz��B���R��;�]��9��q����wz��H/Nu�h��\��^�彨�;������lSƹ]w�K��闹�&lGYtv����A�)u�:�2���d�ij�e^A- �-o�{�?�/A�������<<ъ��똯)˓n(.��^-p�(
�ё�O�ƛ]W1��t�au���q�;/�R�����w�)D�fW�U��4߫��տ<T*?5k<��H㏶<A���j	)}dC=�X���չ�x���we7v� �so�a�ypIR�w!�Si�2�W�M�n-{���a	N`e~Fٚ�ű�U��s�0a�����3�֫wF)u���U�:;���bѦM��t��9x�����!c�ԛ�֜R�_prCղk�Y���3 �]ťU�4�Qq�=/�[mF%f+�R���
^���dP#q���*hY��]�b�����t���"nc"wa�(c��y�]�C~�퉧T�oqa3}8�Ū���B��|� '�7��.	�:l� ٵ[�^s��c�3V؀䖽�&v�9�mE]�pJ���B������d�h�.U��h��$��	~A��od��܆���|k]ˈ^�s�`��$՘;:s��o�o�{2��q��{��!t7�"odx+_�J�y�n�%!�vB�����I��v"��}���W���/KPr��z�l))S;D����f#��'k������\�RE�r�n�;zU���'�Ӳy���{U��
fN{G@U.�>]]����_1�`���-����GC��p�|����e'F�R�F���K�
���Hĺ(�t5�R_E��3i���B\����X5r�싏K��ԥ@���i���y�zx�y�}�8yۧ�5;U�ڞ�Vi��Wi�fpN<����\�S�#���w:�ӫo,�θij]�ۉk!͈��!�ңIn��~1�ڝd3�q⳯y�8���}��i�%��z�ۣSJ�m��f�hS#T3(S�w5�Z�V�E��bbU���5m#�-�ku�$�gA���`���0��I��	;�o��}��f�X�L�O[N4���s�qS�ӛ�p�,+}{F� jc�&�:XS�,@��ҬQ���!WY]W|���Z���;��I3�6�K��}�J��[[K0�G�%�`S�NC1E6zio�}�t�,񱧷CWܡyS���fo��G�����B���
�����M����b��r�ܻ�9��u�)��ˀ��^��a)�Lm�&�m欭���PIP�,��D�8�E��ٮ;|�vr��΋�+V�8�"tr�n��:�x]�fQ�i^ٮ:H�|i۵um(w�sr訫`V����[*L,�b�]:ѳ��\85!��2��b��c����ܭ��vz_!!!BƖn���s1�V�d�p���c�;�a��]��S�7Q>P]�2�7��z�?F���hȝ���]|�w,�D�g\[<�)���v=�_G�ض���j'E��/O^d��3�K �� ��Yzo6p&��]c��*���BoT2]� �����N��l4>���,0U��u�'.�h���{��Q��Ѝٍ�ۛ��(�]�.���p����P�f�fFyuK�rV�/�LėV=w:�h����i,�.�w3��m�]���[����G�zn^7;�Kw6�#"�]���V�����=Mk�K75`ܘ8՜&�-�Ӟ�h(��x\X�wL�Z��܏s�R�Ew,:.ih���+S�u)q�NKБ4��Ԧv^n�o�b^[kg(q����{8�٩MQ����>.
$�P>p�*>��q�Z$����g(�[�\�Q�:��Q�V\1�Ǥ9��yrɯ;ϰ�������*�9wҷ�jcRF�r�&�j�ݿ���:���ψ���km�V�𳠆�3\��T�I�wώ�uȶbv����\���3����#�n_l�e�q4�*�"PbYפnk-n�uz�a���4��f!�uŞ�����Sy�ۚ1K���F7km�r��ws��Ҋ=�Չ˙�Z�߆)m�,��Px�ϭ��э�#���o=��x[Nj�ep��ᦀ�(N'��rٝ)K��w��90�6�Ц��u7pJ�CG��1��7l[O/���<6A����8�9/�w_��l��oTܦ ק��Yع4�:���Pi[�]n��`5mklA�4�W��o��o��غe�)ݻK�H�=�JͻG����B�ڹ9�LY�zpنq����L)�sG�:�t��%��b{M��ؗK����B�iH�l���㭠��� �]����
]ӳF��f�;�$���uت�nn�,��R�HfC,�l(a:5��pͿ��*M�|�q�M�\��c���$؝N��z��V�(ݻ��{����~�����B!!� IOZߗ��6#��e�裧�a�	eU��;����	��y]&t[�[�OLV�3b���tAӲ�&����t�Wi���g��[��ZR=*��wt������p��r�T���r\�&dg�d��N�:�}E�h�=Åt��j�
��~�� ��F�꽸V�7*MM�kc���E*�V|5?U��5��#wU3�aFb �J=�v���Ź��`J}�[qJ�W�k��j^
&��"@�[CvD��R��绵�W��Mk�y�
NG��ȗ���k����Ŗ2u ����H�F����la4z�8����&��}�w��	�贈t�odSk=ò^�r� ��Jz����h�Xxdk/.������5�8�JZa�n���ְf�b=�V<?rٰ9th�T����2��)I���5�w{n�%��Qț�C�)s�#�/)
ӗ#�8�ƻ ��f{�N�.+U���>��ȝJ!㬡s��ήTM�v����f�8E���S+*Nm�z�wwvo�-p�BB��2NΙI��#���<a1���W�/+S����}�a���� ܼwR�\�юB8�?u^x���.Y�E�^���Ǘ,呲��pf��D�[������O�e<R�+GN��74��$,�󟓷/b��c������1���oL��d�� �)�c���bY�9�^=-+C ��.f��>}�l�bN��l�=Y{/��׺�Ny7�8�AQ7�@�i�南a�b�x��qƺ�9�Ô7��'@�׊msA�Y�<<���T���+���K��VN����ӟ:��9���i���Q���G+�-F
N\�-x=R���&yr�i�Z ��L�옷��n:1�(�1�2�P2��f�i�MA���Co�h�AO����ӎ�[���w[��k��S͐�˳_�a��7�6���+7�ve�@um��m�MTD�N���Íb�ױe�r��
�H�%�+'��Y�����JYU�莻��3Wv���M�ƃ���аy7u\��nU8LE�gb`e�x���g��y2��k�Ts����G`����p��aZ0��h��ˎ_qK
�i�ڇu�MGB�<4�����|�ױ�KF\ǵ���Q�ݼZk�D*��{n*�O�j��YhŴǓ��f��W/5����턱�TR9RY|:�Zv���(�����=m�nҔD����P|�Ξ�dF�hC��v������iY�tE2Ӟ�
:Vف�9���ݒ�D�	�j������8I"���q��r�4��ָ=ߚ֕��
;V��i[�;�s�4��������L9�fkTky����-�.�H�=�@rꆁ�y�+��i=�8�VwrZ*&Z�ޭz�����ΖS�j�]����y�/S×1@��(`�UЛӡRN��;i��j����▪�P�d��mgA��ܩ4�N��gr=c@5�nin�\�u �c�="f��`,���Ym�.��.��̓yaR�/;��:��.��V�X[JV�ם` ��\g)0��U��oh�k��<�!:�٢L:_v6�_q��ȷ�½�v�q�	���j�����*9����z���U��P=�j���V��k�]�s�&<��ۨ��p��.2��p+(���dz��Nz����p�U���]����a��I5]u�zTS��^Qp[���NS0ϡ�v�me%G$���bX��^T�!�\�x)��:�o�����Vh<È�i����8�]9'�a�r�2y�N�ЗKsiĸ���;�(�h#]֙���i�v������7�nq�V�Z�$U��"��`���9��lBQ�nR�Y�U��%�6��ά'{�=%0��-�g\4r�٩s�(����Q��*�y���^'y^g/9u��d~�-q��qOf,�ҪIgn���Da��LP�lk�fJ�R��W�ޒ3�s@U�ɦM����ʭ%��7K���9�� �Z��JMOE.9�mK���lS�qh��.D޶Ϫ�*����cdd�z�d�mi�@��$؞��v��U�Qc-��C�A�H�/���<ڻYI0�o�S��ɮۮ�']K7��Rb��[G2�B����)��&���3.�H��G魷ά�P]K�]l��e�}W�V�r��:iQx,�׳�/�VB�N�S^H/�:�S��Ҵ�8��)��m9_�i�dJP�F��9�yԽ#����Q�"�w�n>#N�SBC����|����p䤇2V����U�ꏓ��Sِ���K��g{�7w٫�]`-B��$}��Y#/bvw�H�Qr
�Dts���ݛ������I��.�mk�8�Æ���
ɼ�n��{�fw���g\��<RR%�IJ�c�1.w����͸��MQ��7����%Vu��x�֯���%�ޛ��|���Z<9*D��3��煏�أC+j��sg<�Ͱ��4F#�hn������=�>�ckx��H̆_n�(,;��Rh���
��˲��ż8��uk�l�Y;�����a�uc��x�2u���W�b�Y`ܮd�і�H�pw�;2K�l^Q��K(y�k�"\��+n����75	},��B�b�e�������Ss2aroY@J:�gVoKb|w��(�y��јc&��/^�l>�����;���<%����axK�fQnl� ������|�����dݱ���rf$�R-���+X�\���M����_j9r�2����v�@Ħp��K�]�;5zc�͒{��c֗Q�RA�K�� .���݇���	k�q ��5���)�Egۑ#�[�xC�{}=�{=��1S�l�G�	Ι�Z7H���r��Q��GW�I�en:�U%�c�yWct�A5 ���e������]s���dj��6������L���`Ҟ��o�Z�Q�"�v�gZ�"s+pc�D�^��K�>Xv`{�&M>�M]^��)pA��6�R�3/����s���%O�zD����Q���#�-:Mu�S�B����L]cJ�7�	�Z�t7�,�[�������Ȭ�kn�+�cS&������&�e���pN��m�n��ܸ��Փی@|a��~ջ脳ʞYD��L�o�z�F짲�S��I�F(*dg$��f믆��v�f�Q��:dc�F���&Og�nsy���ӽY�0+��k���-ÑgO`�� �|�9��5?z!��Y����gn�[���
��7�O[�{5��U.�� �nk@��N��s�(�f�S�oUN5l�1�v�E�y{!��IoXc����a6�m��}EU����	�3a�_ ��7yA <�ʥ�Q[20�`�Eh��ٕ��ϭ��8_^˪c�};�]�R�+�)���S��/�s&ЊLҬN�z�m��ڇp:4~�k�A�Zn��B3��٫�[\��LAIp�2���)�m˗yrs{�[�E������������
Z�]�n�u�G;n'��9F�S.�%e>q�2X���V�b���C�nYun�J�m�*δ*���"ݤRN�doč��m��J�&nl��<pB5e,�1/90�q����X����S;��|�� 3N��{�����K�
Uֻ�X����0A�B
�c7��g#h��='��T���u�5��E v���V)�T�s)��Wi�#%��Ԟ��O�gy@	��!��(��N,OZ;l�jڃ��Ƽ�8������/��n_O`R���p��[����k�][�U�CfV���S
��Lܮ��(��N�i���
hX�b���!��t	�ʋ�SfxpMh���g���;6�֓�+`���rJ�Vhүv7�ɈC]*�� *7�*=ޞ�:�$�:��=V���,��ݥ�C��cS'fՅ��"i�nf" V�Lc��K�y��J��N�99���[s���scW@�c���{��7��݄s)��Q��:�e��r���li}B�ܔ�|n��/e� �A,����*�;�r@��|�Z��r���to�ռ>�v�nX���Zg��G��)�z$�e-��^�^�%7�RG���V�bi�>H��\[gD��q���i�o�)�N^r˜�<��:�c��Q�:�+�(4����.E�@�Rf�v�v�����;�[�9Ï���9�y'.�Ի�U����2%�RD��؀�1���:|��}U�yP_���E�r���ߑ�+�ǚ���UOp颯{�7Z)�sV\��H
sC@����2�<�����q�c=�������"��$�ϥ�pv^9mf �蘮�H���wv2`��n��(sP���6�>z�5��0����Բ�+<�����-;=�B�6��u9[�Q�!��J�]���ƎR�+rHnxw�^�)ؘ�����s�C8'qJN=�P�q�ԝ>���lU�ޗl���!�o0��2�u�3�U��'�L�6��'�3UN
��-	�.!w: u /��4T&�����u��f��n�4Ù�$���SYs:�0;v{q�2o׽`�a�|���ض6:�V���!����l�d����l��s�K��v�p�Һ�=�� ���C�:���ܮ�Aiٵ�:�ɥ��:�2�L���T��TqY��h�I�wW! 땛�y7��vC��et7/%����GV���w\;Ip����W֌[\�x��֩@�`b���v����sX`u�ծ�Kc]��ב�:�ܳ���S=Ul�TZg���i�؆U�i����ˣ��:Z=��v�T�ie�p$$&���0r-�otƻ��Ƥ�K�}�-��'q)�_N\��z�^I��VU���K���^�7
�Lz5t�� ����μ���ҭ�ؖ������:�=m��vi;1�v�k�IgR��6:���	�=z��%Ȱ%�t���ޘ�m��o�:~�ﯕYX�xX��,�z�dg��*�'��/w9;�}��:Q�5��>�+k��ɣ��C��i'՚ ��N��a�^c�fՠ��jR/j�^�s���gt� wx�g����B��*�P�,���f�u�+c %���U�'zʋEh"�ٍ�ƝJn�/�{����o�b��3Go
5yGb����P�*�Dt��������u�]C�S�҇:Eb7�emF�FF�`�t�x��g`��s�Nf�l̑�d��wj���Z���T�缏}<���
vD�m:��[&V�`��z�S��y"ē��Ii �s�j�!OG��b����}�}[Vf:��Z�aoCzu8Q[�0�/oB�u[#Iͭ��e�b��1�j�EBo^��5�u�5i�9��]hqY�b�.����,�M
5�sվ�t!ݕ��D+H�W���nZ�*q��_�������6L:ʦ}>�FN�.ٙ��|�z��M]]{<�Uƽ ҆Y�Z�`AN�Ŭ{�u[:��F�.�h���9�A;݊ۀD����Ҹ���Bc�zw�|�gV�� �N�Uf�U[h���i��W���,��1�x�Z�t�6&.��n�U�mu�q��=�U�.u���
��]�5���Ȥ��S�Uy�8�a��l`=��ӔV�4;�ڞny`~zc��;�rB�;#z�AL@�!n��:��Q�读��8�� ���$��
��n��<3ęeח�{�������zlw�/<�g�r�S���M�iM>���΂��'/���ҽ�خ�na��R���N`�=i$�g�/�Ps竦�Z�[�B\��{y�4iʽ�����5N�hZ�vEk������
"]���ᴺ�]`G3a�k1�ߘ��9ק���4�3Bi���
癨��^;�w��uO4�1ѵ9�)��onq��*^��¡S��	s(���T������)�y}�2�$�M]�;$��y�vZB�$8>�ٻ.��>�@ok��x>��g@��'f��J�Rv�Veh$a�{��+������Ӌ��S�}�KX�P�q�z�yN�~[���#�O#L*�$z��x1X�]�7ے�M��}�cw��(K�+�� ��c5�Z3�!�+t�����x��~��qBx@��!�ȗ����2+�qL�7���˘���f���G�9>���]�sz%���2���Di1o�is.�1���p� ���0Ɂ�'f����v؃Rq}ۤ����:��7�C�զ��E��6�Z/7��ݴ����b'���#�F�f���*�G�yV
��f�x��>�� L��G.���f�.M��5�⭚�C�'7mj�jR�S\	Qr�V�r�����ż1�7Ud���ݠک����4�k�Ɠ.��\p�w�Rv$�Df���;D;{K�[G
�X��sE�����a'���A��ބ��쒨��cz�\�)���Ew���8׮���S�gr�b��3�vД)�P6ŭ�K.v\�y"�*�I Q�n�$��Į�5�R��R�Jk��ԗ5p(�6̾L6�9a�B�Ȱ p���+�M���ɲϬ����M�bY�/��{�j�K��J'v���X�ov	��fU����$����nC+XsY&����gi s�-u\Uia�.TSBnJ��+zZ�)�fl�1��*g�[7B���������x�xkt��W��!��sGH}L7j�v?�q��x^_v�Y�{#WW�q��^�gt�s�7�X�+)7k�e\�mhCn��*�z3뻮�U�Dj�KR,��R�ގ�� {��� J+2U���H�H�_RY1�=���D
6�Kd�j�
�ㇱ���#o]i�z4�[:텅e�����4;Y#$-�6�.o|-(�\;_�V{3n'.x�_z�pi��d��f�ezղLIx�y@��i�$�gk�����3K�������u5 ܩ�ʻ9ۭd[W6�8ud�a��r�e�5�v�'qzp�H�nƫΏE�ĨN��^s�J��j� j�3��s�'+V.����{��.Ba鞀0A�h}u��n -�6�L��e���ӽ+A8�w��WK��Z�vz�w8�������� /No=�#&ؔΠ�
��t��;]�bz\�2\%A��ÓG�]�ze�.R$�@��{h�HZ��%;l��D�.I�s����>ư��􆢚=�d� p�;��;��P{Wyb�(QC��(�!�z��9ܺ���Kz��^PszM����C��wkf+�\	�m%o��u�k��Y���%���8��"�@�u�͡��i���ʟm3)h;Qj<�S����"5����h�^�t�V·7�F�l_'AnybB|tqc;�����N��c���7�i��q��j���c���cZ���%x�w�'�5
&�. �����L�=;p�q��NV����ַJ'�ں|�vN8f���\�6�k ��@ʺu�eoTl1�9v2SW.�zM4h��ͻp5�G��H�S"���F�R�#�P@�ɓ ���Ch�/y�Gy'Ċ=�qu-����A�{Ǉ��b�!�)���{F���r�Vi�w�I{[�(�<9�7;i�Ŝ񓑤�}��r�?y�Q��
1�aU�W5C"[��PX��UE�LIbAkD+Y�E��U��\j"�EE�QR�ciU[j�mX�%UV(9J��X�J"�(�P��UD�PSMc�UkX*��"��cr�4ʪ3V�G5qV�:�����TAER"5*�����(�W-�)-�s��QT5h[H1Eb��5YhWNaKJ�+-*ʊ*�*��Z�"�D̡�J�Q�.%����TEJ������Ń����+�����L�����V9j定�AY�4�����TmME��ʸت�YZ9KPiE-�E�V5(5����T)mEc-m��i]9�L�E�j2ت+*ت��墈�����mDEU����崥�TEZ�E��Ыm��-(��U[j��q�5Mat�f%QFҢ��J���e���
�ڌ�f����϶�s�>������f���\��r��i�nv5�B���r��I�.�>����ͺp�ۗs�}ե�cD���xɗ'P*)Kr���}.�>s�{�]v��xϕ�f��
˱�e�}���#sdO�]㲜�gq�T{�q���o�\)\���F?9�d���l���C�
�F͊��k���i@����8�.H-�by�6�(ŞU��s�wŕ�����8l6v�b�]b�:C�yuB�ЉiY��T�t�B�=,�
��:L��yCb�u���Q���:vM�MCת#u�����7S��3sx�ڻ!�S��L��ҿ!	������«��p�Sj�:������}:�dO,k��[�C�D_EX�
6���"����%\P��^��y��}�֯TA׬ٴJ�L�S*"�
DD����$8z-�T&@S���2-����WB��fqjO8�+n���oeO���=��O̖�����S����<*b��T싈u����ϟ�B�֒��,����r<����������?%�Ŷ7�����*8�<��b��ڲ!q~JT
�s���y+�d�X���xt&{W�bW�ť֌��>G��:�v6�E���K�㋟=7�)�2S�V���F�:V/����w�P�g����gV�C���+L+�2?$�0$����^�Hrxp9O����Ӌ����%k@���(r��� �֟qo��A]!��~�eP*�_���yi��]$�**�L6�;���D@ˬo�c�D-#�a��zOg#������Z�x���F!�ԓϟ�3�7
/fm���~��҅�۫��U�*��7s��9����e}��GL���_����^"�Å�k�Dp6����.�&7/}_v���e������t�v�j6��Y�+�nym(�b��"�mTkM��ԃ�G3\��×g�"����W�����	Mb��4�
'fƘ��f��v����m��$���r����j��'�(}�_I��z[zx6�tGjAo�p�l>��jyn��61��
$��p���``�<��җ�XF�3ѕ��q=���黤I3�Y<�o�Z��</(�%���f���x��dtW��5����ٿr��F;�ί����6�n<�;�$�`D_1e���4s��"�������8�������iأ|Ұ�㧖�I�{j*��H����=3e�7N�\�,���x�H��k�g4%�HfQO9�G2� t�݈R4�)H���*�[|i���L��3s/f魜cJ�j�7p���o��Xm�k�����ع�<��U.��[K���K���՘S��7\�԰���.�7R��~�\S�\���Y��n��h����Y�'j��3�P�&!#����4K"v����
���d:������{�o�q���^2�-�+�<lc���T
z�ܐ���;
�+��	�w�V�g��cl0J��b�|�����K�N�J�KvJԗa�uR@�绲�^=�_1k�iK��QuI�߯�7`�x��=�G|
���F{Ϟƛ:�.V�N��3��1�� ^&5ӷ��g�ѱ½���@�]Q�`C�B��-j$�f�4��A��.���(�8����9����>vE|�+ֹX�W�Q��FC^�e��^�M�;Ο+<`#Ƥ��s�P�6��MV���-`�fz������.VD���Y���=�����;[��ytVE�\�Mi/��ɅwC��!�t�%�������Ea��F��Z����k�P���M�a�S8jFO���E<�>�m�w��3;"���Q6�w�G�����m��:й�A#ӳ���j������A��F�����Gmr�Z6�{�ۖ;Z4��+�VLo��nP�rGhA�Ѽ�v�
�[O��H�Q|��5
*s`����*�C�r��ӫ|�w�t�}G�������j�m�����2�=i0��@��%M������l^gvZ�s��ܹr��^y�9��	��k]�bѮ2��U� u�����������֖��ֻ�4����+�D�<��9�o��z~G��L�TQ�ׅ�qٞک��7�jی���H��-l�E�RW�=;)�'i�W`c�0�Zi���N\nM#�S2�f�>������d��S/�;9|s~�"�!9��ᦼ[<H0���V'h1�c/V��Ӟ�*}���# (�r3ڥq��Өl�"[��$`�����uf�XX�&*����ݽ� �b���0��(v�W��q�uX=;��,�o��W�ƖAChn1����Җw�<���C1�ghDD8|p��P��;/I	t���
���Ex�V�;�k����)����B��CGν�x����#A�/�׭j���~԰4�&����Qo]�U]��5#f$Μ�ǅ���`v�]>�9�YO�Z=➽:�U�;��Pr禑C�ȑ�{}2yx�f*q�4c4y�"tׇ֍r��x��VZ��L�1�YU�'����G�W�K�n�ΏC$T�i39�2N��W�;��X�S��v��b���ǎ(��V>uI�XJ��g���i%*7n�}t_N!4�`��s�k�B���\�U��n%.�7��SwI�	v\4̭t�37:������c�B�X�w$���aD;�8�'k���Jl`��&�$�[NNH6L�ǘ�:�Z����+3��b7{�()٦\.���+����v��.���Z�>V�v��+G�D�g`L�X2����#�Yv��� t���ly��y�����*��^ߐށAzF�� ^,/�xF�ψ�nVP�_��'����n��]=[;P�����d^���JLnh�ua���<oFk<]����nI�wk����6:'�����j}�|:?��]�+|������3�O�OTFW�nk�.�o���غ��T
���	�eGk��#,6�����Sq�^��Y
�o$�?l��5����3=�])_S�v5_��S;f,�%C/���(�A��_n����u���E�J}��yy���I�b����{�?�����"��h3�nVt��ח0�xك^�c��"V�Q�	9�@�!�r�m��;zV�<9����#^�P{7RE�2d���V��5n���w����N�Es<��ԧQ��=ZVWj�d]r}XZ�wtkaJpZR��++���>��[��pOy�U�u^3d��/*��U�EoǦ���8jӏVTԫ"�o|�M�b���M����뎆ŵ!YԦ^^3�f�2�$�\ld�5h䘻?�c�H<�������\����~�}�ߒ�X>Uq�F�5�P�Ɉ�٘�*ۯL��rV+�=W�7��77ː�6_���*vX*n-7ZKb�Tt4��ܢBno_��`�ep���r	.iP3�Fh�2���wT����ɡ%�4'U��Z�γI�-ʬ�q�̔h3꡶2����&(k�.9Z�!�
�t�a���u�P�y���N{G���5e��/ʩ�7�'0��)+�U�4'ɜo��7�]���(8�)L��gᗛ��#?��_���t�_��c�y���������dp�wu����r���������7j�ה?:�f�$�0h_�ME�:ϑ�V��-6Fh�<Q5�;^�4��E����皻��∲��,U��*K-`��*�y�0�]��m�Vv���Vr�W����&6�����W@�5�ODd_�:r�˭�r{������)���`��u�.K=�[x�s�[��}|����y�3�+je��nX�$��Ck��jf{��w����|��m��{���|:J2c��WRk����5jY�{kc(0'�,2�O�Q�'�`��ݠ��p��f���e<yL��M�+�޽�C�=������E1'b����8Z��H��S��U�k0�:sP'L��	��C|-1��f����!"���i�!6�*�n
�w�%�W5��f�e�sUz|�t6���UԼ�u��~�DC�1}0'�}�3R�$,��ә��.7���1���^��Њ�'���@�.&����~�ٴ������v���@���� [�d�N��4�u���pD��(���MR{���w�����F���
+Uz�ӘF蝭�$&{��t(�sj��4�xY`�*����;�O�2��og����	P%�����t�=;*�d�|[��j�=�C����y`痄�]��A�f���$?���l��L启d89l�:T�}pD�=��=淫@��v*��^�W���v� �E՞犺�*��s����^�n�7ݥY�=������4��Z�J��+�X^�b��4,�xo�u���J��,�Τ_[Ո�-�\�s�T7��q��U�;�p�hڱ�ؙn�3p̲�3���O�����q��������IM��|��ň�}�����;*dn����8�5��vZ���<v���B�b������\�͋�5W���&#C��8���<k�Xnv*"�ʎ�����	��1�"��T�3�jgw1Kg#I� =�A�mR"�U:��ad1;'�E�s� u	�/��N���C���4�����\kq^�P�~�����G�����7�n�}d�E��Cd��"�b˅�ޡ��ϭ]4�n�4F}5핎���=��j�ٕ�o�r���睒�J'MS��ߕ�㧻͵辴
�8�HvRyn�6a�v�$����t-����|��3ef�u �}S�]u��W��<��$ �A-4sƺ�j�^�#q{��|���4"25�E2�Mm������z�3ׯ��]J�M;�R��Ru��-yY�x�ڳC4mq�>q�l=N������ԢA��Q(����ӗyԫn֡X���>֤\����q��ӫd�7N�3d��0�sIg��:��c1��Py��2�v�!B�(\��b��u.0�=;�=,�C6��EW�Y�祎Czp͏C�f��eO�Ïn�x�؁���|��)r��ro;�m���R��-:�w�4��Β-!tfY��L<�*Wy}DZ�'�3�MLL�����R��|���9�:����y�9��Q]!����;��=[Wr3=�c�:u�����Xߪtc��mp��ݰXQ ��+�3iԚ`�pL��\����n��7yl��ΐ�0Uk5������vQ�@I.�"��v^����;��=' �{	�����7�ވ�eg��{���(FP���x�����F�Orx^!��8�}G�vX5�N��6�ٶ]����s�޻ՁG�a�NI2�q�h�?v��v}�v$/���kA�v�n��f�Ǭc��')��8��,���� �{�}�LbQh"I��u���E�C��l��9mמ2#��R�Ǉ]����aD7�8�9�ː�@. ����y�	�a�;��$��&�T}�VI�Gp����3YA�\bꩁIr��&3U�[O�4'��umrΎ:��Rb����	����S��eڳ��{.���N{g��f�%od]s�t|����{}a��Q�{^l�����6��T�nW�(h%�W�q��&v��K�2"��^dds��d]���df_�������x*3Y㎧���i�~�i31M���j|B:����!��g�~����,2��y+�Ec�I${F?S݀ռ.��D��o�eZ����rnl�g,@Xyx�e���>hv���bs�睼au*Q�39W��v:�91n�i�oV�B֬�ܣ��C�j�l�.2+���q�la�ʵ��t��X�3^ �u7mG5we�Y��T̴E�O#���*���p��9N]��[zA���S�.��3E/d��������VsIO��m��W�= ��ؼF�-H�pפh�{E����rl6�/jxpz�X|'��W��ģl�n�6)�e�;n���^�G��ew��,F.~��`�f�������:1���6��'en���ꄘB���[ٱ%<��p��crFԺ$U�zX>Ur�"9.k>�3����������_l��Ǉ��њ�L�ҽ՝��;{p���P*v_���M�9A׻�r�X0P_ v�/��s�՚��6���[dY>��Ε����JJ]�='�Dbwb..ue���0�f��I��+%{��恟=�/U��h		�Y��}�FWM'K��NbN�׬/G��f��D�6���=�����Sט���!�]i5�E�Tx��[r�!k�:
��O3�v�ܮ�F��X��ѫ�,�'�ob�o����l���}�Of�P�N~����o�Jy��!ݼ*�v+�Zbє�����8�S�v���>Fٽ������ͮ������s�>�ń�v�WD
=��6`$�ī2�z���?s�'�K�뎐���קi�z�3����u��7z0�5�ڹrLw,���i(�.�5<1@����O�)Q��t�[]�]Բ��c��рg5�588$����&t��떳F.��ɔq�y3��O>��޴5��[��ԝ��Z�,cSpt���IA'e_i�w�
)J͎��H#9͈n�>9J�w���7s�4��!��݊�7l+�����S�^c�1�{ P��L�jANf�+�`]���6�y$0���wQ%�$������6��l]H��V�Ϸs�.��={`X��.{i��ޢcP�gS�<���Cּ}��2EzzF�H&�r�)Di�ʾv[�G���%�M�T��y��!2�����ћy��8����Y\�9\�	ґ^���*Q�/X���u�XX��5�>k4-�J��I'or�������ؓ�=�v���)���IP�'�� -��V�p)�^�=�`��=31��X�C�Թ�	Y;k�b:Ͳ1��:��K�nvs4w/�S��4b8����*�,=phS#�! Vf���^��f�(�Gˣyz4��}�-��r�kS�ΣV^��� jGH�49D,9K�A���`¡��Kv�<|���-=Hs�c��׼�"����"�u�����2�vh�W�H$�+Ke�m�ʮL�1�XD��h��Z���T��:��pm՚&�L��v*�:��i�F+����)�=T�+ra�Q�{sTڕ���4P��B̊����ȨDhS�ۊ��E� ��'\-@I˙��X�G�rn`�Z�ކ��[U�$�D�1�S�'�*Ѭi�;��4�
��5�޽�>�g�ٵF�ؐ:��p)����Fn3L %�cCQ���~!ݙ�v7���0�kH�N����%�����k2�.�x��#-U��˸�³�<F{Μn4��&R�Z��:f�CN�q,��mI!!��;��p��k��f���
/���ӨLg �-8�� ��5G��"��:2,�6;�Mcm�,��S�l�4#�T؃��5�1j��`F�خu�Һ	j�O���N�5��ԗ��  Z�k�)t�ڹy�;�S5@�d�Ub�r:�X
2VVis,�����Z��G4 J}\T�٠p�uYaKaT�+k5R� 0��	�AB�Uj�cQp�%L�5c)V�\W>J�Z��B��Ph�V
"�P�j���j�hڈ�U�6�F��,kTE�Q�ҭ��jDZ�ƈ%F�-"eV�D�VQUD���n�b�mU��h6�3-R�FZ)[V�*P�jʫ���UU-�)iD���Mr�Z�[h����V�Z�Z[b�J��r�b�MeEQ0j�KJ��iA��[j�E���T��U[-��5����!�Jԭ����PmmV1-՚Mj�J��%�Z�+V�imRԔi[B��ktآ� ��Q��֌���-�A��dT*V��U�[R�Qs0ŕ�E`�KJ�sS*�+L�cU�kAT�\�731J�R�ĸZն�d�%V�F�R�-(�4-�fZ�R�6���QJ�J6�fcJ+h����Ū��,��TmlmZ�ZR��\r�TVe�B  $�8xޝG����q�%��`�6l��S]�Uzxr����%2��(;�����ம`�A�uiS��%N��:�U��o�z_;:S��G����u�~�|��_���'��t1`�3�:mA�P��o�+wz��Y-����C+����ڨk����*��8yk@�v�R�x5�dv�U~�V#�w�o�s`�k��3U-%�XZe�}���i����"���Jk�?'O���]-s[�s��+�L���n�(�?D6���7�bz���	2������WbO�k*k�
Cɛ�`K2���0�5M��w�j�~�?�_T���[O8Y�-��;X�����!�ol=��]��i��[@4�!�i�4"^��^��h�#�x�uMd٘z���ga�r�mU_*��Cj�*�PK�Yi��iOk�L�s�k<���׉#T�����6|��0�f�.6%]t���i��QWz�` oy�~�7'T�����z�ؗ�sJ�.Ц;X�g����R��-8FQ�T'^ؙ�"u;��4v��t�o��� W��hi�W�!�V��-����7��n������5�U�=R�Z�M.��;2��=�F��K�bfkds�Ɓ�bsd��[:a����l=�I��s
��L��Aƴ��c�"s��,^���T]P�ά�y��jlv�Y��u �����9L��wBx�5X�����Cmٷ��4�ϥ�7�%��R1�+:��+��;O�KH�D���_q��{��N�G
U��{� msK�+���|.������Nc�\H�1Y�18.���|��~�|3�Xl3l�5�s���[>�LY/�J�
]FXV�>��^��Z.��<UЉ��{W��`Y9��\p�oH��j�an��uL��"�/�nTF�Xn�T5C3�R�a{�.o$�e�����Y��3h�G��Y��L���̇�N���#rl�l�5��z|���C+��5��ˠ�ö�auSۜ�O���i�;:��쒽��V��uz�](c��#V]����'�s��ٷs�	C�f�v%S�>��WN�ś[6�<�&�5q����=���ekDp��UZU(Q��rVP�Ǽ��S<�igte�y/a���=�������}kⴎ#R���W�At��3)应�؋�ű]�ˢN`c�\X��	h����d�Ў�D�B�{d�!Y1���;�q���b�=)�Rz��<�W� ���J�˱�NX8s��1���qn7����t�5��1�m>�.K��.I��_VZ�W�S��JHsMH�<�r᫱�eur4�2����B!#b��V��p������>rwz�h���_u��j=;���׵�6G��BĦ&+W���]O.�c�N�Y}���63�s��܌�^46n<ĕ�E�*�u\P�N76|�t�n\
��Y�ਫ਼4ԢA��n��j�7lt��k��gUz���'�{��B��q��Eq豈K���19w^�;.g6�u�i�#�y�7V>�,>�O#~S(@�������QPc��괎<a�[#Ӽ!���-/3�G�L�{{�3%�7�V���՞�M]::� 3e����J�2z=պB���|B��Tn�ueq!�<CѩEz�zW:���(FP���!��0�h��&Q0�=�eu]s��:{zGP׷h��j$�.X��Q�a���W��)���*7�IM��W��!��o*uLc�r;���=1�ާf�r�"�ر�X��V1�R�=�X�����lf_n����5������.䈬�#|9:�6����,E��7٩�U��6#�s� ��>�y�~��wj�LP��<)���<�({[d{��k���S�7�s�����NK��n�=�yv(Ԛ/dn6�[�a��S]]�%0a�����������@���]Ǚ�\���:,k��{f�zp4ߝ��S���q��a*���&����{��w�)leA�ݏ�j�Í�PW�fsTʾh��&�FK�����F��^�����e���GPV]��
�˽�V=�Z{�/O���+���}����.|�W�aؕ�CNO���b������
4��r{���s"��1��ZKV�CD6\DH�ѿ5#b�ٶEXo�ف�n7-���=Ԣ�mV�m�{��J���ރx01�&V�!t��ѱ\>��Z#&C�v{��s��U:w�a:<L,Xu
��}��V��������a0�CF�N�*;^Pؠ�#/�(�ٖ��߬�6wd���:��%���D���3�EҔ��&|Ձ��>�%3���Z+K���,��j���Ġ��a�i�Y�(t�IP����C+��J�b�cM|�1�^#(�	�C/�vbo�{i��{��Ხ(s^�`b�T}D�@�
�l�!�r�nn�z�o+�v7ֹU�w+�s��#�1�1�C��z�Y��F 7�?2Z�^-��{$���y"%��1��w]{��	�C�#�KrKʮ;(�<�598٣�zU�X�/1�J�=�"6Sܵ��u��8��|_\Q�#�P��q߳�o�T9r��*�p ΈT�W~���GvZ���ۺH_j�̌�ͣ�&#�J�ķy�۞i%;����zkޑ{���g/sNwL��3b;�����͒f���;�
�$z��>�9݁��8	��
���R����;1)����0E�i�<E����*m^uKjle)L�� V9q��E�,�C�,zl������b�c��}N�R_��w��;������(i���貌g���oS&��|���O�&�<����i�$�M�q�g-^xE�1�8�*ɚ��2F{��z6sZ�.ʩ�|���[�&<~qƽC�,�����p�g�
S��Z�ݔ}�;A��{�$�7��[�IjC��q�ڨk�"d&$�yP��^4#�e�|cᕣp�0��z�~���㝡�T`lu���6����tG����ы�lY�j^�-;�C/_�d�RS�K~v���~Ú�*9._e۶��e�]���=߭��g`b�{;Gj��5�Y:XF@zo�s�v��6G������{L��{#��|u�ufU[��QY|�>չ�*�^9'u^��Qt<z�{B�^�v�\)ļ7��{漲�il�kg���WkFl�2�Ν'.ԕj�+:j�nQ��;(��':�6�y�a��E���9��+�.UۛS�9�����a����R�S�=�n��d�R]�}�Q��C�O%�Oi3���gN�.�_S����v��՚��I8u�:����d{��5��Mk�cj�Lb��z��_����OU�T��.$��~s����ݷ�e�ZfEz��������`���r��:��P��p>$�������ʿ��zyܞN��p�L�)�+�md4n��
�$se;��Un݇�r`o���H�K����K8o*�����$���`hC�^.;U���lM[����dd���1+A�Η�j>Uue��qc0�I%�0�I��#A*���DyC�t�bUt6p��'�B^젫,n#}��ےr~�;KeW��LUT�������d��v�}�,�]X�H�P�x�gj��y~�du��ү�� ���v,�$�@��-�oh���j��@��՞�J#C����=0��=4�+�u:��Q�:Q3O;$���mK�P�>:��^�x��ڌ+�xc��$�s��ҚY[]�i�濰��.;_o�X�*�`#:����+e�:��i�����)��E�fT�;
,�Cd6]c��T��.�t�ȝMrO��G3�������o� ����-�4��x�C] ������=Tw���Jn`��=O����X$tU*�����ޥ7�g�9���A�B>�ݼjC�7��yN���.X{=f���c�,�GC��_b���
��:�Hg�l1r8�܋��K��n�z|�讍Xve��;>��/�1��O���=�U�ˇ���^.泊��i3c'�Q�F�:�uX��a�<�^Y�P��v�x Q����Ot;��9� v�܌�??k�,�|�a��j��Ŝx�X���W����u��>j���W63��%�bS�2d���tG��׌�ٌ��HX���G�k��sX�=O9z���>;O
>�s��F������#q]������{f��jk!���'���#�&�w�=����\�X���ߵVEAS�������rΗ�O"\m���^&{��]ߘ�M#1�'����ȵ��z1;J/�>�{�Y� ��)U�q�3��Y��jO	I;��V?_�Q5;^b�|�����/2]���6*1��W���;���{�hz�ג��1�+6�&8|���Ad�:H�w.�KJ�Oj�t��m-�j��i��jaz���ֽDՑ�y^�|�y�S�<8�T��(�����P��H.��}�^ڌ�N�}��<�*�V�vfk�{[p5�o��/Mq�/�i�P���W���v:�؝��']py�&b�$0ٓ����ul�.���
r�m��ԪK��M�Wcx��M-��i�����}���Ϡ �q�nd{{[;bS�5���R��8>�N�AS�_v���؈�]��J{��e:
��q9�N������CY�T�\�8xrخ>��׼������������~9]t�����v/
��KI���UF��O�n������=rB��N�]�)��8����֔�ƈ�i�	xoS�8
�#Y�\`��TD���p;�����v�fW-�V^:�&R��V���#�c�p��7dE�C��SQ��c�-suY/o�ESzޯ�'�VӚ�h��-gԻ�J�V
v�{Kg��[B��FfQNN�dݜ���z�q����1��\���s���8�V��Ao�=�S�O�;)�ށ��yK.f�\%��;�<���Uzv���LRy�a���\Ʉ0�x�VFĭ<f{�e^z�{P�_�t��p5T6�dW=�0+��vLO����o�Nu��9�)u��1�����Z��.9Y�_���:"��br?���Ŧ}ذ� ����Al������wmދ�����덱���i���x�[9��&Tv��6(#\Fr�����nL���u>���OϞD1O��3��>�گӈJg >/N��Q}{$@v��f���W�J�wf��+�����p�wy�=��g��nC�<�ɋ�wk�O�A��{ݏȱo�W�۾|-�d������Q?w�&�Fީ��d(��QF�J�OP�d(�,�w՗C���)4gU��3_-�o >�=�p�Q��Ul��ӑJ0�ܷ���E�o�����t��+���|v�6��X�Ψt�sv��a�8h����jR����C�@w%�A�����&39�������3\8��"�l���ؠ�H|k��i=�����44�P�3�����0�w�xݟI��f�Ga�4t�G!Dq�ge����o,HU�ذ���y�w��Q͡1ơ3C�HT�'�N@�^���(t�]�Ǧ������I�/C�ON��6P�~�H�Y�i�eY�u��n�|���y�1��>����QBs"\&��l由U[k��,nuAf?���VI�r�*ۭ�����a��"�HrhaXL�Y��H��i��������B��U,�K��oD����5�hG�O�7���xJ�X({��A#F��Ω8�r��)�3��S��4��·�PזD�NJ�	�%�@F����F���N���pB�+���#������F�uN�f:�жɋ�:�n�Ǭu�?]�T����9Y���:!���YWMl�=��;.m�vwE��wۉ
��8]��^�jx���;da� ��ծ�&�ηo�B�[аm<>RR�+𢡊/('�J�*�+��u��[c�����u�tˏ{]�H�9�ȸ7s���A�X���O�Dޗ�8k�dt3�Qq�q��g�}�y|�%�}��õh{�vl�f7�}c����Hw;��1�tn����C�z�
<l%�댝��d1�{#�Q�X|��+�͢�ew��eF�S[%GP�8!Ç0�Ԍ��Upu��ʵϙ�zN�"�lț���c7e�To��)�ң@���^x���U ��,�l-�{��\U��o�l��`����t����n���(}7E-�#�$����nƪ���^���vn!���+�BFY�	��,k���ev{���^u�&s�5i�r�I�so}O�D2}j;O�I"v��qث0J��кd=;~n�Т�9��^��I� �ɚ9^OA�){q>F���\����=1��GN�V%WCeg(�8p�2�����}W7���ɾ��`x��
��2;͒'�4y�>K�����*BP=���@�
�TB>�����ur���'@t��:�Ίwgit����ZfqutQu5l8���]��m^|U�]&`'[��!�w'��}nm�Ǽi
�	�qZ�uّm/\]�LTg-U�5�~3����{�F(լ�o��X�-��ɛ&oF��q��zm���f�ٝ�zJB��P=���j�Tz�7��ө&.ӷS���o�ջ����J��|�%ҩ���͠�[�5RW�e ��Nm݈߇wL����^�o,ܤ�հ��j�0,��K���t��W�t�5�}/f�=�r�n���F����T���g_Woe
��%��v�4��s,;�4*�9A�'Hr�[ő�m��tZ�JH=�h��sV�y��En�Ӭ��]�mC�o5b�G��t1 T�T;�iܺ����E����:_j�s��Yu%�4{V��I��G�yam��'Gn\p���r�.��wn��]Cb�y�0���vv�dk�7;��x�Q'�1b�eKa�y��Z^��hƥ�GTu��P{,YV4W,?'��W:�Ӕ�Ȭm�{�Rny.�hA����g��}�!s�q	�u\�4����8ב};�hgY���^�ԗ׃y7�J$J9Z&�Z���q�`����yIe(�23�ذ�#����ѹ�OM��ܝͣ���ʝ���{���qz���L5�z��9�~��8]j���8Y��wd�ӌ*���u���sU
�r�n���μ6nG}=;9t�b�:�g6�X�(6��Qo׷YU��8r}l:˷}���\T^ �W�)Ѧѩ}BVȕ�(�AMJ�槹C2�4Bj�m�S�� ��i��ϹY�:�WϻU��^�����XY�.%&��\G��@ ���4)�$�il\�����v�k��Wڻ�<(>;�nu�`�m�z8��~^C5��WA��2b&d����Cp� Z�w���MY��h%3��]�s}�=�~�qR[cx>YQy�nq:(�S��Z5>�3S.�WLqv�.�� �Ҟ��[���#JY�Ԕe��C/n�����O��$v5UٻW����L
7{��U�͈�q�UXYi����Z\Z���S7h�C�`'4�'Ru�KQ��Mq�~ܬ�x2�U��PEѱ[�g"#O�!�}���t�T�"�{�Gj/��������iʦ�O�f�@�ږ6�AX�vs5^[�^��"Mu�[���u �N���R�N@Xl��`�c��t�a���]�ˏBN)�]�ְ�S:,�@J5����57�L�bB�[r�g�r�}���v�WI�(�|�m����-���&'x3W �4AQ���80�гqC�LjSͥT=���2u� �"�NJ�|e��I��g~�w�L��m},�J,�em�=˧�z3�Wk�0N��^���J����1�ƈPѡR���Ru�X�j�Cx7�X�1n�����C��yܼ��E9v�]�z���L`��f�:�aǈPH�}���jU�~�հ�����k�_4n`�Y@��ڹt��j�9�`��Y9z�E��<�IR1Fp-�q��S':s)N�p�]L��sN��+���x=O�k.R�=���M���b���Vj��fzC��mV�[d�*Գ�����J�rb,�ilU�*�(���騪�R������ĵ�ж�-�e�Jֵ��k�Q)u���B�Z�-Q���Z�����Z�U�\K�QZ��!��\���USEŨ�UiKq�m�J�q�TT�Ap�-m*4�f�Qj���L�*R�Zh��-J�.Lm�[kj�+R҃
�B��\V)D,-�i(�jEPe�Klj��SL�+SIX���:��ҋ[J)�)��e�Ŋ9k-J6�)c(��KKQ-t�4��4�JԱ[F�c�Jĵ��.�*#h�KK�B�Z�hֲ���6��������h���GH`�&8�eJ����2�[jĪ"���0���(�U��QKD��Z1ZZTR�����QTE�U�b*8���sU�֣'J|����C�+�͋�#/����Q���tt�quG���ܕL����	!4�b�m��巩B����>�{���L�z����q�,�=εo�zK*)uKd���[g]���f�f�Ә�}��v�^1֨z��[�Q���7>]XI��K�6�6��a���#mLJ��=�����O��r*�1�#��϶�;�UQi���'Uq�Y˷^wQ��gȎr治&y�hM��Bvs�Uul.�.0����P������mT�x,�-���x��J�!�=��r� �i!gN��f1�#�)�Y�=��_Ý�����{�˽�+蜿.G�������߇��a��@f戤.�r�Y����:W��=. ��
���=h�f�����s���^b���-����<��u��<��葢�?�[����<5"��mR�nO>� �g{����g����s%���9����W��6����Ôz~4X��S��\R���_��k�+���ݢ1�Anj̣�ྚ���3A9�F��zl*����ـ�I��w2��!�3���ɻ%��uC@�ڧ����uC�>q�l�����е������;�a-;��뵻��}F���7fӢ�^�ȷ�M2y��;��:�(/��/@�
���o6;���U�y����[Ң]��ΏC����ͻ���,r�[ձ��]\��]XܡR���L��N���ؤ����%[�2�hV��[U+�?xx��r裫Y�ke���}D�Ն�{�5��vGpP�a�K=î!��,/v��_E;�-�e�q���wϹ_Ѹ��KV��67�K1�UXGq]:�V���X�b�ge�8�1XX��V{]Dm���H�B����o (�P^�KJr��P�Q2y��W�{�������/K�����nm�,r���Ef�R�m�t�"0��@o��hmw0�_u�Pc���d��ޜa��hq�bWϲ��qa�OI2�|ډ{���ٹx�[�A��mt�ce��������&�K�W����~�D���|�(��>�4I�2L`L��Ĭy}������.u���U��
.6��f�t���빁^E�+�:�����Sv/s���Bs<���g`���iB	�Q���Q���C�Mv+����0���m�筮5�}:��Oڨ�w�ߚ����F�s(+�Vr'aL��(�Cr�7[�K�'Z�ꍈ}5�G'�z��v�v|�I���)j��^?*VF�ﴣ�*Vw�%�>�����8��tXo��V:��Z����Wj��������/<�p��&n{�V����cM�x��cL`�K��Hw'��u[�F[�3���9V���Z�rO1���'�R�;�����#�w+-�y����	3�	�pb =�������+{s`�����sk�4�Y���ڡ�5��i�6E���9x�;W�N9Փ�5+u��ݯ-�+��)	���	�vF?����P�&	.ܳ�z��ʪs�;���5�ٙ����z�J%�cH`�v��g��ػ���)ZԹ*�pa�W5ޱ
򾂻��CK��q<'NxMD`I,��u�3���|~�]Y�
��d��e_=��R�)uS�kM��e>6�o
��P�Kj��p<�Ţ�yǼ�ccO�{��÷�M�0�W�t_��	6+����Z|>��W�U\P�׆���r��:}�:^�	.�f�Fe!���z
��Jޗܳc<�����@������9:,�(�Q�Wl��pl�&_Fs����"�l���!o����Ot��PǑ�{c��q��z�^�3�<����(}j���C�:����t��S5���(��Q`��g�s���˝�fs��:�y��KԱ: :��Hƭ!�<�w�_g8}~�V�����=�����W�E�Ҽć�^f�c&؊��"�ut{��"|�I�s�| ��4"��KA�:�ұ� l�Wh�P��4b裮İW}S�I�;K�R��z�=�q��bŖ��Q��C�`.85q�Y9M�r�з#���ٽ�l�]ɼ�{���������qv�X���Mz�� �}b.UYr�K��Gj����S��b�XX�v�nxFyf]m�{�"���,��0<'Ǘ�����E��F��Q�P
ØEJC����tD��A o��)�u����2��x�Lt_mT�`/��=k�X���:�Gt����Z<�z�7'rF���k�)�VھO�tZ�"R��?<#�Q	c|�q�n��*!9(�{ug�%���-|�f�Ugj��z�0=}������d}����qب�t���-,�u+wbK�s�\>���o㪼*�eE���X~s���Q&V�������{�t�����4�����[�EŹ�u�{!PZ�<t�	M��7��")_ݨJg5�n��[�]�v|պ|u��o ]�bmy-7�-�	�`<�/hz����Up삩Jl8�>C/���\إVĆ�.tY�~�>
��d��<TI�\�W3���g.��i���⣗�=u��s��X�7���èa���[����ë��ID-&�3ْ{�AU�B�l��ly��VaS��z����)�ж��Ck�j���Y&�f�\��c^�9���
�z�N�َv�s��8�y��6��~�٥������
�S9�3Eu�n�Z�ذE��T��_���T7{ �^q����^����{��y���S�޽����� �Ң+�=�v����s�+���sM�\�� U���<�e�䚲��'���#�#�O�B���D���b�Q��ܕco�a@|{�n���_F�
>}��)~��<3b�A�]�&yV_ã�б��8����,����.Ֆ|����+y�;�z)�f�q`��K��]9f
Ļ5:��Ǜ$9�m
������#^�C$�����o5��af���Z�֡��KP���[%jw~��X�	_Y�O�gW=.g!WQ�\d���ډ�S"����3qua&�6:M������J�\�o;�y��ߣbuNG�R�Ưg�$*�:�җ��^�\,��c	3�t���Փ�,�/�/�ȴX;!�N��u�׵$��M�o���U+^D9<f6M-T��7v��3n�65�(Y��K3��VT#��xkr��ω՗�ͷf�ۆ]�n���⻘0�o�n�s�y��k'�W���g1t�vkn��0��o�/���F߳���U����լ��M��;�B����p3�����^v7~m[5�q��%�o&:ʎewҹF����s�@.I]ѧ{_w���ǂ/s�Y�	�܎�%�&��r�+�T6��{Ajcs:�l{��|�;�9#�o��a霟ݬN�9��̄J41T������r��l`�v�'l��Ik�;{VNm�+꯫�q��=�=�J^o�wos���5)�w����u��=��Y8ry���#Epv��*�yWٮ���JY6�ن��,�O�ɐ�o��t��3����!_q̾���9�&SW��L��]9�1�G2
�,�.S��1#2C��2�a���U������b�Q�]]���]W�E�U�u��݆PZ>c��`��)��<��ᗋ�����N�$xI�����=a���u��6�U}ބ�"q����K��׹���(��D�BW�h�M��/sp�7�j���[>B������b����W���I�܉���b1��ճ�~ǈ�v�S�dڷʲ�s=
5LOG,���&8|��^&�ө�1k ��] �@��p�J����̀Z�԰�dT�^��m����D]0���+4)3��2��r"T��C�@�9�a0��_������m�v�g�9�X�LBs��^D���9$�f�����=BS��|.�)��G6���	�[A��;{*�.'�bޗJw�K���7@{��)>!�$eﮟJCjd�R�Q�e�B[����ޡ��	���z=�3�XABd��>q��Y%���. %9%:�}:paO�s�UW��xOV��!K[wW�">v�W��p(��:ws�K��3>�X<�k��U�"Ƒl�}~�8�z��.��2�=�>~u���k����S��*"9k�X\���E,A�1�8�S�퍜�h����mT���
N߃uQ��VI����l�p,�b���XX^&�k�����g\=\��� ��w�îND�	��<���wq����l:�
�l�x�e��:�E�R�Uŭc@�*Ud����c�CW_�7���x��<�U�ݟ��Z-�y�.C$��&����w����偻oFk8���_)��gJ���x�#�G@��W�x=ѻz��;}7���u>��x{��b��=��Y뙎�����^����*9�z�i����/���*�f��m���*�{(T&>Ir����vh%�_�e#�}π�`k�7h`�a8�t2�P9��XyN:�[W�@ȨP%�D���|[��I��{ȧ�k2���#n�Gr*�X�#�Ed�
�|%�>�W|a�xk��@w(��$���%�����0z�M����/�[և�{��Z�v�Ef̈�0��$	vr�Qח �xw6\N�<����B��;����s�n��7�6G#�7*^>u�8�
�.�0N��ə�tp�E����^����	q��{�.A،� �g+�f��؃4#����=ڡ�N�9�s�X�1�ύ��ߎC�h�:/�*��������q:�Ǳe�P+zV=��������M��~v�Y�9a�I��1���;������1�MR�'���o�i�<x	�	�O�c�$��	׈�݆3N�b��1���ggg�h�H��K�ɼ��Ry�8�����Zb��=f?{`bN!^��|�~`T������X�f��%���
�Y�)��S�y���f�| �Q�:{�>�Ă�'��v���`Ws���rc+:�!��LLH/P��d��!�-�~a����r'P+�?��Ĩx���k�0=�yvpN���|������~��ǽ�0+�?d�E���!�s��<g�J�����i�5�����I����m%aY��AgזiJ�r�'Y�<M����E�ER~#�yA��,U�=����?{f��a��Y����l���Ws����h͜�N���{l<3�AH���w6�Y������O5d�1�=<�i:�2��4���,7=���=q ����3������6�'���a^�x��?��R�N&k�v°:�}����i�La�����M�VWL���I�*
E������&yAH��I�X8��7�� } �q�_n�rnr�s�:��T������~�}ۦI��rO�o�A�%}B��Y=��g/,����Ax�m=��m�4�^����8�@��ٷl��g�3���;��� �Τ��LL���a+�\g3��W����ʇOu���:��3�=d����0����Ĝ��?���g�H)(u>q7����%J�>�����7�d�Xz�M$ʪ�� �`��m���׷�:��}���=$m:kYPP�*���ݞ?$�bO���!_Xz�3Y�4�`q�6k�&�̘��O0���ψ�a�1*}�~��1"�SG�2~|x���5���ϰ��3��vl�U&�~�>��!Z����:^�Yt���a�F�;�)ʜ�1b���\��s�����7G�x��E꺱Ԣ*��#��s�!���s`H9�v`�y�����u��2J ��ɗ}���Q�0d��:�ZAiSo�����3Zu�qM��� L�d�����������N3o�
�����hi�s������1;�>2x���5�!������h.�V��M�l��&3чS#�1�
<�}~��ӰH����UV�C���B��ӟ����'ڠ�_y��l�O�g���p�@�*|���8�R~g�~��1+������-d��w��1��\�l��6�_����H/���o���{�|}Ӛ���% �Ь=C`~k8ϓ���%H.�~04�N��1��!��eN���+P���O̘��W��'䙗�C�Өi�e�O�o=p@�G�����G�V.ttނx1_uW�}u��{��wڐY�%N����Ă�<����v��<߹4���(q/���u�Af�8`q�ACԬ<�솚������;��������Xk>�6��2bN߾���'3�y�u���La�+�L�fm'�+
���Xu��eCsvi�����8���}`T�N&'��:�?���:�'�9��4ʒ�O���ߨxT��Ǿ�ۑt��Ǹ��a�f�޳?vz�����i�
���L���x��8��Y^3��M��T�30��'ڠ����Y�N����b����?;t��8�,^�|������0�oy��������������AH�d��N���i����7<�<O�O'{��C�bA���. ����aL��3�~��J��u��!X)�6�>0+�>a�����C�����~߻�y���{��{����8�=d��f��C�/׌Khm
�̙��}��6��b���;�� �L����� �^ c��SL7�k����0�Ӊ]Ϝ��" �=��cܷ7��fgo�ߞI_Ri��xP�Ax��ި��Xk��sP�'������:½t�L���+
�����`()��a�|t����������Y�G� ��5�u?[�Q+����&�]0+:n����ӌ7�rg�+�'�SI�'�����$��ϲLAv¤�,�Jʞ�I�y�@�+%ew;�M�ĕ
���4��1��PY������-�y�|ÿ����t��vH�ٻ*M�؜j�z�hFt �s�}�o\Y����&�Fum������k$qK"���}v��7r�`j�Z��.�9è*o
�Z1���[��/�M�Q>�tە�včҺ�8�`�4��J�z/C4��w�{�� 	���(��u��<��L~�g���S{��~v�`V�CO>Lv����AH��W���q�S���4�^!���kt�z�@����4�j
q
���06�~��{�Pw�l�YT~�O\#���?{� 	�Rw��Z�`����k6�^��|3�M$P:��a�x�Y=7x�C�K���봝B��&eӿ߰��X��5ۤ�Ρ��4�I���.��/k����vV�������P�����|�go2J�PSG;����@�a�bcACĮ��@Z��b�OP�Ax��hi�jE����x�ݟ�1<����a_�'�Rm'�*~��w�������~��l'|�Z�z��OC�l�C�m3�����4�`T�!�Y<e|`^w�0�I���gud�bJ�=/�z��^2lߘm��PĂ���C�m� G���绳�n�b�4���d{Օ6�;ChJ�S^��~gbJ�OMP���'����L`q����纞3�J���?wz?2i��O/0=Cd���C��!���#o�H"<��:��ÉM�ft��jȏ�錁I���N<f$�
��eAO���i���:�g���:��*sxM<B�S�;��4$���ý�YR,�O��l�¾�����x����ˁ��o(᛹P�ߖ���������B��G3>`T�:�'~��Y�y�
bO�] nyLt��X|�M>Ϭt����1C�Xq�LI������T:�AC���OY�5g����xD8�d�ɑ[�\ػ�ߌ/��z`�O=�M$�*c�N�5�@�+0�u�i=B�̡����,��dP��x��c&!�>L�O�8;�+ܪՓ����~�
���Dű�ڠ�U�eŦ����os>�3i*���ɴ�<H/X{�a�m�<CO{���b��
�q������h��lֲi�8�Vx�H����S��1"��Y�o(u����}z��빷�<��O}�|���S��O\0/y�����>C������)�<�Z�Y�>�5�&��2�O�3�wXM=@Z���`V�.�3���R��+�+:��_/����Ӥ�f���|�*�l�.��u&ۻ�F��k�(H��=�U��go
�5DU"���o�pçц+�C�2بQ�(~ǜ�b����7�ۨ�	����cJ}t8�.J��p��Sѡ^q߮��y�7�of2�H�x٦Q�q�v��>"`Η�<�{�.5� �
�a;!�I{\���[�(7��CW�;4f�A��$1)vV�e���cZ`�>�Mv�3lh�Nj�0����'w[~�41��Ϝ���Uŭ+���K����c�K��f��S������a<�U4>��O�aڀ�p�W�xo��yԔ�n8";���#M��Q�,�=���L��^�К����_x�[Sf���.9�va�'"z�J����r�'2�~���	�F�����C�;�2/�DV	�w��uc`Iz�zKH:�'ފcňvI��w�����
/<#�4�2�޶;p)�u�:#���hWۅq=k:��L�CFL���|WH����Sz���-'�{l���N��g���pm�R��J�2��p�;Ή���uMu�����|@�틒�;�qF��f:�vh�l��3���%r���D�������C���˳��F� �.���z��j�����Y�[��Ԥ(�͜&�@yw:x��s�;��;w�������(�\Eu���f�͇��þ���+�j���I,c��:��=��ݝ[�'>�QL�1��9Ӣ����]u7b���2� �����WeڧhP{6n��aB��al�&3�D2�A]�+ �r,�j���.�R

]F��vݐj!���O���cK�15Y��H���Fha����ص��Z�tewt\R�j��p���mmTq�)��.�ؔzpE��!��6�����Nf��D�3veX]hiX�)B�ٛ*z��uJ�#��qXit��&Ț�ԉ5dDSL��&v�1���� �KVTV�$n�����V��
�� Zt�IQM��XN ��
ڀ�0�Bv7��$��ExEF����!k�p)��u���{�r��L{*\��ۺ���el�p��m�c���p<!�#S��Op��Ѐ��zࠬN?���h�N�����b�B�*ʹ���m�pՇjà
71-�$)FI�d�5�/�|��њ,���a
_X[�K��c�A5�~��Ѕ(��01�d�����J��R�Ϯ�VC
�4꡴1�t�����sֵ�elh�9&�dn�kͤeY,Z�R�V]��k�p�3����u]Fy��IĳD-��N��� ��*��\}�1����2eA���t4�D�f��Xh#<�{-�s�r������{[�6T� ��U�O)Vܖ,9lf�0�Qr����7�]�A��S���j���Z*,UU��Ԫ ��[Gۓ!Q��Z,�X���7�ŋ1��A�����A���+k�`���TZ���[�pŋR��D�-ŵ�QD�V5(*�)F��r�kU1�U��R,XұQkQT�R��U�*"�q���V��Z"1QF*�b��"��8���8�Kh�`ւ��+EQ[DQUZ�UE��Ҩ��jA�ڱ�����b��*+[����Պj�X���E��D�EDQ����i,�V

µjQ���DD\f�!�Q`�#D�Q�J�DX�V1EVb�TP�\Ub�R�ԴP���ų0)q�X��Q�W�Z"��UKJ�\k����W+��P�X�j*
̵3(�+R�E��F6˪U�L�+mD�mDB�iR��/�����ϋ8�qE����[��[�1^�wX*���]t�Ig.��Tv���-<���ќ��j�IF�4v5�l�5����C�L���)�>��mU�~��G��:�����"���θI_�����S�%�x�?w!�J�g��kz+�AH���N�Ă���$�T�x�'����n0+�8�}M��*��s��}߮\�����Xz��!��P�1&��4�^$�i����^?k�!�:ԊK܇�$��L~C��h+=d�{���i
�3�x��.�̆��:��M��!}X���Vv�v[��LxǼ`�x��^�OY�L
��ϐ��q%0���5'�蘐Yĕ_g��LM����ɶx�$�����LAq�Xk%eO����O4�~t�=)���Y���=������)��'O��6
E�Ƴ��O3L����O�`~k�����N!^��|>,AH�&��kR8�O�`o�O&���I��1�k�vf:���ɻƔ�n�?��`��B�+Y4s�����<f��
��Ax�`����1 �Cɿ����Y6j�t�RW�m�<� �i����O�4��Vz�a�\`T=5׿��U�4�t�UZK�M1����0<"=�%J�o��:grM;`W��Oi����R����?wyL�3�e��ԛ�rT=OP��[�<a�ε"��qĞ!Sɽ�_|��^L�Y�Yˏ� �c� �34����8��9�Cl6��;��E�ӏ�w�f�*�߼�m�L���y��]Y8���L��I�,1�5ힺH,�M�X��=LH/���~�O���}��w����&%a��1RW�OɈ.'Y��d���ɷ�1�SϹ��6�gRcy�;�P�"��>a�<�"��.��N$���%g��B�Ձ�_�<��6��;{�����?+8������|��g/N���A�Q)�_d��*Ag�k�g��������O#���jg����Z��fC�g�����ͦ��
�ß���:�$o�d���R,3}��]�<!�+������h�R]��:�i8�g��&�0*
i
0?v����J������L
�������Ak��m�a�����~C�1=�{�����;]�Sö�M�+�e!�3�e���:���-DX7�������=� �`R]`L,�hd��LlѾ1���f�4�m��k�u�;�)��&���8�tC�<���!�;�τx�ûD�~�1Z�ڽ�.	����aޑEf���x{ܮ�R
{^U~��Gi����d�=ɧ��3�I��'�T�~d�R��o�COψ���<��i�~����H�Y>q�xg쒳L�&�O�}�u���F�}#��k�)_٪��� d�{��?t纁�~eCs�������{�Օ�Ɍ{q�&&0ǈb}��}d�br�k'��&���L@�VJ���$�|yf��E�:��#�$`�{_U����t@���~��>I��z�W�O����''}�6��W�Noǌ
����=� /Z�^'3�&<M!���i���>��i�sY�C��`T��}�|��=y]y�;W� ��Q�cϬ�i �!S�T�!�����8�׌�~a�bI_S���r�P��uMn�:�O����w�
�=�R#����C�J�q���׿WW)����@��1�}3�C�~OY��	���a�8�Ag��ox�R����<C��1��w!����ʇ��0+Rz�;M<d����a��t��7�1�9����N�^�����ԏ�1�c��AH���{��L��g���d��퇲�ĜC�d�y�����,��7����Ag\�mRu>Ld�g{��̜La�P�� �2z��Y��E���Gf��~͵Q���0c�7Lf3�I1��i���gg���(i"��7��O2��I�Vq�?$������ĩ�'�=�d$��'ɏ�
�����Y+ư>�u��A��~q�-��3"�ԣ�����2_,��M'O��i�ȥC~w��Ă�'��v�ZE�]��@�g��ϰ�4�^��,���~C�H),8�RW��d��`��xܕUd�o8��x	��j�g7���3�4�b���!���'���R��I���u�N��_5�h(q+��&�8���ɴJ�tk8Τ����w�?f����lt};��Fo�R�����P�G�}�|b�Rz����i㌘�Ī�W�H�y̝Cl+
��^P��a�x�������OP�y�'����m'P�Y<ϲi�PX]'�}���{䝖މ�#�{F��邊�^h���e��v���Q��(ˬ�uj�N�JZ�Ԫ rk�fo�z��Si0c�'-�n������?}SY�zwgn#r��zZ�T�N��2h�������s�Kcjed�-g��̢72A���zE��=� ��RŽg���M3�$q%T�O'����1�:w5b�^2u3_`c��Ƴg߰6ͳORcY��%ejɰ�p�'�T������&yAH��ؘ���dz�a��u���g�*zӧU�m�~@�T񓷙��
��+ῲOɷ��꒾�WƲ{=��K�&:v{|H/���4���^��������8�@�8��g�z�y;p%H.'����ús^pn��{�~�{��~�T6�$���8�0Ǭ�o�a�5�Wf{���@�T<����������'� z8��b���M�1�d�S�x� �'�9��a�u4�o��>��{s<�s��Yn�=�W� � 8���x�Y�����Ԩ��������~C>��}a���4�`q�6k�&�̘��|�L:�y~`W��CL+
��l�I�):��O�j��o#>�5�����-�c#c��Ｎn P�>�|�v�����I�9�=g���Af�����~LHr�x��N'�����>�z����g�m �d����������i����{�o��}����ۨ�m?
�����Xv!��B�S���u����^n��L�O�3ד��6��T����51������2bc������E���Xl���1��\�c�i �`g~���޾���j�����1 �'O)1�
q
��1�N2��q>�M�i*Au���)�:�3���x�Xc�*zw�0:����5�7���L@�+�3�=M<`T7�p�f2f^$ߏ��|�n��_d�;��ʯ�� ���@�5 �l�?����?�Ă�<7a��'L�����(���P��$pC���a��5'Y�~O��y����Ǻ��$Xk=��{�࣡}��]�(��Q����&{��x�:��W��6s3i8�aXW�i�"�ya�.�1��H|�ɝ�q=�v���8�2�nì���P]���I�q�OݳRUI�z����jC�p��ߖ�-����xL��	�^�o�m �a�\�6~OP]0���aXVq�Lv\�?&2VW�޹��J�I����'Y>���K����o��@�T�<�������I��������HU��M��b�u�R� ��y����=�9׽U�i�;3�&���u� _!"�g:�6un��Uh��=�v:zN�)%�����{�֘LQ3��\�p�8�����{�1{	m����th�oW����<QX��}۳��jgm� �'���`�(hZ�t���b��'�owu�4��C�����P��$kg>�ۼz3ml*ݻ묽�{����v6q�bq�?E�'�����A~B��SF��i���a�����z�]2y���u�1 ��Pq
Ϗu�]0>k8��CH*�Lx�`�P��^!��>3~�i��9Oy�~߫���=��,���(i���b��w6��/oX��`x�g�L��;�M$(~7����Af�3��I8��Ak�]�6�0�i4��¸��s�4��q ��7���/��^|�ި�� �c�	>�ǩ?3�=Ă�����,�%`u�������ǌ���9��1�XWn�1&ЩY;˧��R
w9��^�1<�2B��Ϭ��f��<�_��!y���T�q��(�e��W_�|�?Y>C��'x�jk̐>g��|ɦk�5�|���8ɦC�����?g����Y�"��߼�����n�����N���޲i��YԞ��3�J��T������ٻ�u���x~�I�
�7�B��K�=��ڛH/��d5�M=f y/0�PA��o�����
Yzd��_2��j��@��·�x��*T�>��V
|���u�H/P��>� i�Pٯ�M>���ɧ��~I{ |}v��W�2�������=�k�H�����u��U�e��n�\g�T�i��A���[`m���P�=��%v��4w�x�a�q�;�f!����̀�'��4g�z������:�XjOP������I�����U�V�m������������OP�Xw�4��
C_��Xz��O{�m�hu�}a�~��x�`T�O3���d�+��6ԟ���wy&��*��~��Ă�{��l�HD/���"Oǫ"T*���u3��!��`(��C�X|钲������|�����~׏��LIP���A|N�{��L5�!�S�l���m>?wz?2i��O/0=eq�W��Ci���}r�o|D�R{n�=k5ms�0<~d��M=M$���&�C����+��8��01����0�:��*sxM<B�S�;�|�x�_�~C��|`V�O�~�ԛq>d������쟻X��j��t�f�wi����A���y'3������dսx�
���Sɣ9�ras_Z�_^MK ��C��	5;��������Ύ-�/��<�y�R�h%�|��5�Q#4�P�ܰTX�!�:u���	��ݓ�ٶIdm�&�����П=��*0U��p�݆���G�xO�C�������ő4o��$}ԎWX�dw5�N��ꌲ�ޗ�x�l7,�b��`t�a$������V+��#[/�,�pa��KEF�^�C]8�_���QD_��{�%>
��D���I��9�}�{/w��2��ǈ��;���=:���#l�(�y�d���H߶f#���1���^捻��ox��;j�Uf1#��J�p/������myc�8f,��`�[�W�^��:Z���"��S�}N7 ���	״�r[�E2�t�w�q�,+��V�����cڭDD��|5��n$1�{�Y��/(�Ո
�Y�Ӕjv��PO=����׼�T3�?<�4I�閭/!��u��)�m�
��=j�f<1z8�o/jsF[�z���rCڟ<�S��!������Щ�p嬥ء6:l�H�r��Xw�w�<E�κ3�g�<��G���K�I��\D5�U��2�����"�@lбy�|�
�ާM[���of��) ΍rP/����v�C݃Xl�M��ʠ��܏m`�-�z��9�|o{��.W��Q�ި�;�&�������tG��E�wN�l*�\��[B�b�#���l��Ƭ؜K�Zݡ��,'LY�y�8k���Yq��U��U_=����o��K�n��q
�k��\�W�<R5��������Ȁ��EQG��*��kg�2ji���^�����"�"#�ڙb�%ZX)��g���^�(�dΔ2���a�`*ܸ<��ZK_>[�~H���m�ҷ�,�~K��V�	O���HV�P׸�&��wXl��t�����6fwO1��F���Ƹ��'B8��D�mT��(x�w���p����3ƺ>ح��>��Z��p��=��8�NN4�)�3�0�WC�r���j0.38;^^�����ң���4�Ni�֕C�D=�:��7��wώ?�V��/����ѩJ��y�gf��{W-��yh���w���Z���1�ю���t��c<���8h\����R��&_:��N�k�Z~1P�$���X]�^�����u��5X��Rz����m�V�_�h*YΆV���r�ZX����n���f�� �V=Ϋ�wF�-­4ř9��Fs�m��b
-�NDw���`�ޤ��)`��E��+S���tC�cfg^�=A�(� ��.��k�ݭ����k�q�ף2ԭ��� دROz�p�X�?D�D�rzMy�1� �i�>�S��=�����V����V�s��\]�;���S���gW>�ۓ,;��"ii'�Ta�Aq�����f�n�Z��a��$��}.3���s���<\�鋔��}�(�Q~�A��Z�[��훯=�j�u��zJZƕ:���I{�\s5�P�Ô��Q0����.�9��2�VUM��	�kuu��Z��@~�s�[C������?�Q�C}T⿺3h7u���yZ�q��QU4�k[�k�b����C�
Vj�:<U��W���]p[C;�ly�Ě�B�v["��C��$���#C7o�v����]5��s'��=y�.�hK�_ǧ]��6O��3����<ۧf5�Z~���^��+)�_y*��ԡ�Z��lNIp�q�4�&��6�!{���Ʒ�����g�H��M�2�n�0��^6+��r>�泀�K'{3�==��v���mL�s�v���Y]e�Q���	�;¸1α�IR9��_����08 �Z����������	zNB&m���6����+�X��$H�\]T�Z�;vV� �f�V0	W�V�
�8s��f}wɮ�5�H-P[�@!I�h�#ZՎ��pTZ�}�
B��w�H���a&l�n�j������ ��]L�=}�
Gq�i��=�����hbE}MbR�7�|B�-���Ϗ���4&������V��
�%�(G�xʫ(W��e��cb�̿7a��ᑢfv�2��f�1K�uc�b��i#�����UFEDP=ū��\e���st�锢���+�o2�Q~�M���|7YŲ�	�>}�d2OrҼ��̛Hl�,�;f>;y��:�f&G3��,ޓ�R�D$����|�]a��\м�1Ɔ0��X�_½�5����uq��qn������R�Y3>7=��Ǎgl�x/�6�ے�u%�v+���T�7�D{�7=�M��%t�`%#�0HxC��=�j���*%0|c����B]r�;�ܬ�c��O;���w� e�r�g��:-,0��b�lu�
=ѓ=�.�$�ǔteEwf����t�v�Ҥ_�W��!A�Vb��/ar�}`�Vty��:�g���]A3ˢ\���v*��9�ϻ�/"E��К�/1瘮��-�^J�U�xF#�Q���|��F�E}V�:&�ا*U��\��V |�Kn�Ô+�V1��5ځb���A̸�zP�m��O^�T0dp��e��4�ӒKN��9蝇Q���>ӌ�{�;:���TQ��NV,d_R������t�<���ϼ������PwW5���l��]T�8045tQ��@�®	mq�[�4�l���#S����it��z��ǵ�(f�){���і���vId�Xp�b��~��������xU�c�ź�S�e�uΣ�K,sR8GF=�ح���=@0����b�'�g�c��<�1b��f����a�x��ۯr���xن�wK&���%���IxG�Y����G�j�ޤd�ݬ*�����u���:���52�!Ec��=��))[[���0^D�9蹤T �l�{=��/h�'c�_ɻ䖏����Rv�o(:Y�m%�L~��璉ú�Ә��"��XY�(�a�d���G�o�HğsR^��K���L�������cY������P�Ǵ�{�|�����R�v�� ^dև��5��3~��WWY�{"g԰�U�	�*�������]Dg\�(�f-	��o�E��A=�E�8��O��w�3���A���
����q�G`�u��<3���G3Stљ�7	����}�����KZ�:��-<"S��{���tr<�A��m����S'19�p�K���4��^�
&voe!���T���G�M�'b [�V77��.�]�i�݃a����"�5T��+����Uӟ{�x{;���'Vxݮ}�??��=�_�]Z-���N���Or[�tE���NB�����_��;g��هI5�t�*�F�mv}�>YmO��s珼t]U���@W-�v;DƳ�VT�o�W�G2sI�<��ρ�,�G���$Χ)i��VV@�*\m�;��Q|�h0�֪v�"٬(�M�k��(䚨,\A;����
���Ø�w�CA���y��s� 쵄Mׅ<����P�ݵL���k�Ҩ��Ƭ��_�di�{�eo��~@��o��m/
�VѸ�40�A��#��qc�V��Uzu�ݹ�₽�kY�������Y�����b�������υuc�u�n. W���%X5f1��T1('G���������Eo�#/+ɑa��|'���p5��#Q���X"|ϴ"c��ck�S��["�q��ۦ�>���/r����}��Oj崻m��U�5t4��V�i+�1UWɍ��u��3ڗae��2
;�+�t#���(�U8��3p�䗴�_Uz��᭲��;r�Wo��Дt��n1�lL�V>n��.��N�u7�����kj��z�Vg@���=�����}�O|���)�L�o�oii-��^O��b*�%˓�Z�H��0F��3bv�cm��-�=1br�[H��Vآi���cw8�=�عI�?m��t�Q�W�:�-��3y�
�n�Q�&�'9Y�������:c����O�D�E�Y[��v��l)�9�},c�Q�ܶ��Р[=�i�]���_L��;u���>��a�c� w������1��8M��!/e��zZ�y6vѭY
CmK_Z�s�.0��JN���a4WKzh��zj�]W�/���2v_{[�^���>:�%Qd��[�p�}H�5��.y�\E�7-�Kl����w�H)��tֹ%-s:��v��3`�5.�M,���g�(�{�	�#��g-�/��^�Ŕ/���(��4�F���/�[cy�}I(�.w5Pi�K.�΀�\^����⬘�ǽ�s�!U�
��ssR�t�9���ɥ�njӰ��esd�����Y>ܚh�7����N���c�gG�eu���^����wi<�9ʯ�r9�v� )��Kt��U"��uNם�J�D�0�����2�++���u�
�?Y����h�w�-g��z���r����v�`�eek�*�Glr���e<,M���p���-`�5�n����L)\(�C��	�ʬ-�7����H��p�koH��qZ��0I�&�=on��X�V'�&\&:��%���!�e	b�)^��
8,_KSMśX�5�e@�Ad��!9�	��$�+-�wf���Ew]A�u"2�2���&լ\�A���iwL�0�4໣7LJ;�շvB&�nS�,%-բ:�2@��mX���/�%��ėKp܀����Y�n�lˤ�mi���*�J����d{q-;��RףP[��$qI
�g��Ň"~�N�0٭4A���36\�t��C]�X�rTEe�Q�V ,�.'ML2���뀴���i�E0h�-��4n(�eZP���]?�>U�wz�K��D��3d��vn�k[�*w!#&��i��ňh
����˫������#�0ԇۨ�<Z�#{��l�ܙ�^���K���H!Y�x3��\����*ֲu��>:*L��i�KU���)��=�[�q�T�>gX{�θe���V�s¶�v�[P�@)�����~�������C�PGT�l�UU*T�X6�e--lDXUJ6�m�*�j�"9B���S��.�qX�1X"*E�iU�F*�l-)Ec�b)��TT-�UQ`�%�UEQF���qRڬQh�(�+(���b��,ZȴUVF,�U�ekT�J����)r�UU�[Pb�ƶ1�DYZ�ŌPc��.�*�S(T�F��ŭ�P�FUb��Y�U�iKJ�����mQDjFEUQ��\d�(�X��5���r�Z� ���Eƨ�\nZ�P�0J�D��E���-L��Q�+4جF*[,T��T�AV ��TF
���m�QUEqm������dTEQT�� ���PR����D�4EQ��F �b�
��UY�[vy��7���`~�w�c��)g�s�j�H��̔�^���ɧ<{��ʉs�@�ǎ�=����g�
�X���6�O�{����k�b�;`]sR�Q��/?��b��<���vy��
k��7
�[1	v @Bk����'��G��7�.��ݺ]�T9�d
�n.��m�>�c�Ecñ#˸C�:[B�>��������k�iz�=[�쾵#m/TZ��[����a�CD�}7]f>��P���nZ�h�ނ��ۚ�WOD[5�.���)K^j�d%Gl���]{�9wcP~�n�u��:���~�.����;%F�̇�(�[���F��Vo��O�M0��ޅ�eh�{eX�6�2��F�"7Q�rSo���[�r�"ָ�4�'9M��j��=�γ b�GlM6�qs�LՈ�wQ;���{97��y<ՅY>����V�u\m.��m*�������W�Q�^��wH�ߔB�;��oٍ.�
]���<��<]�D��:�s3�,7(��7�we����x��G�P��Y�.Z0�b�c�44��s���1ü������xJ������Q&�FΦ���o m�/e XL�'��.k�v���׸�o�U�R`ӜU�s
/��wMd�V%(�=��x{��Z�Ըjη�f��|9�*���c�Fb�6�]d��-�t�Vom5��ww�+CW����;�m��V��mx^�.q��}7w$��IĊO�����8�y<�Ym���!_B�s�B'轎�2�ӵx�w�AW���(�B��[��sv�=���t�C쉼��t�₯3���N=!S}c�ba����`i"���4��;{Jk���8C���</7�z�o���m9@It�W�g9�A-�wU9��]��g)jKV��O1�Iߑ�v��PTt��'�X)t�v��Cb7�+D�E����O�US�7ޱ�cT�΀mtx(����lB�ʰ�Ay�W����*����Ց.��ԣBߚ�;h:.:�[��[Z{V�CxJ�Y������J�T,oD+��	��SvhzT�h4E�㷏l���d���;F��{Տ^���yN���3��N3�B���!g(2��S���2>Twb#Z�]p풯��#pTo��s���h�<�͆Wp����u�Y����	�'*��S�8�	�6]�sZ�T�������N��k5�앥n��]i�R";��R�I9�h*�����5C�	0>����zJ��jV\6b��ꯪ������ |���w"yfX�YC�p��
�0��áe��������5�!�k����cU8��_d�Ŏ��s}P�sʤ�|���ڴ�W7�o/zvll�^r��x�L;��F�Ɍ�=�����L,������(��ŵV��8o/FK�YA7�E�vP_W�uקs
Ǜ� �8��ma�iVa��=��O����uS@3ީslɤ�hs"3	����{��u̺ʣ�T	-�F�80�{�s��7SƸ��{��x;$��뻚�z,�<'�:��Վ�:�Nz��c���B�ұ��Wdד�}�K��.�1f��^x�ՏM�8�Q�^�A+�gڵ��JX���_Aq��q>%�7/!�N��W%}ƻ
��`~����G��w�	�^�#d'4�Ƭ�f?u�����r���Ii�a/h�7�Z�pZ�fP����;�eUe:ݭ�}1��z��V���[&�Եn���	{IM�W�n�d 5;k�Vf���H�t��1B�Y�}���l��s}s���t-����Mr�8�*mC*Z�s���nE�m;�z�2%ݾB;9��Vf������n��t�aR���s���z�Y�;�+0PڨZ]BwWM�}�����U�2Ȫ;�^���:흤z�d兵�����!mY��k�1=���kw�w��ú��c.���"�����9Fi�+^X�فVk�@����ޝ�4&��8�
��#����Դ�J�q.q�Н�"Wdׄ�{v�{�L:<����вs3��,+���{`��P���@��U�䧒*T�H�"�Y��7����ܵ٦:��%P	0��|�jF5���㛇ohM䭉�{����)�Mn������l�Al��	ֵgDu��F�P4ݬ�.ue�݄���.��Xœi�@������:�._��荦�jM�
�Ǝ�� ܖ3Gd[k�/�Y<,�*~�����輲��.+���X���V��os�J�kS���U�|���*�&��:f�;��ۥ�B�m�����nŰ_XW�E&�7\.��<#�#ʌ��Я�U�}Gϯ�s��~'�~�s)/ea�o�j�^ڧ�"}W��wO�,N������jg3m��+l��JrË���\�M�����6%h]�}��-{ms��li�|½��m�xz�z���]��:�����W�歓�e�Š�0���lk[v�>S������!P*Ұf��#]�Zg#�p��k�m`�L_S��w6j��}8�n:�뾭o%�ݡ���=ڛ��R��Io9�W���Op�\�����]׈=�c�Kq֡��6�U��X�I��:�P���������PS���*	�V!��kZ��1S5t�S�����fRv�kּ�#���3����Izn7�z��7c�b��qfg��~]���'�[S�p�C^j��s9
]��C������,N�g<�J숕ٚ�z��H�W}N:|��E���]L�>[gv%p�Wp����	J(tZ��p�c.nX�-��O������Ĳ\J��R������I	䚾��ww:�9ӷ_R��Y*'����:��<�!<�oz�-��Ϻ�{�]��(�h�fc�Üzj�[��,����K��X꼈�4+�.�*��6$N�W��ZC�R�u�7b6w"V������8:�T9��L<�A݊r�E��no�2Ok�l��pb�5�Y���j��LJ�E�E-֍��^�q�W&Ob1�v]N:�m:s2�/�W#���-~�w/�Gės�qBUq��F���p�z���a����F�q�S�M�K%���X���v�ڒu��14���g3�;���(g|���r���#5.����@�oU�3�z#��խ�y[g�e]�_���ݲ���x�ٶ�9�C'������}[3��w��W��d����/�dB�x�k'8ڞ������~���d�ƴt��:��"�s{��㧛����;Z+`�fe���*���f�4K�,�@�Lo;��SE�~�"���&�v;{Y	�S�.;��{!ױ.��~(͈�����V��.Ê���rX�/u���h_<gMۗ)���y��6u�Q]��T�3��0��(��v�ӮP��E�Xѱ�*W��q�gWMjroC���z�_-�3.^ǃ�LO�y�Q�]*�0�G�uq��̩O�(��ޔ�ظ��Aq�������^���;!N�zn:�B<�
���$�5����ۻ�.a��6��UO>���5�ݿc!�n��5�^J���{DE��2���3[,������2����}�9��W�)��
��r�^n��W��O�{*���=n&Z��48[�^����=�x�����%��!:�L(���k�cN��U ˲�ً3ۗ^��+�p�r�W
�7���[
y�h�{�{�r�j��a���:�N2_d�c��\�T*畫\;�7��ܧ�3-s0Fl]9��I/xFүNfW���o���:)��R�O z<S�w�����q�w4�pu����9��C$���Ai{r$9y\n��Z� 	a�d���\!��nT�qX�#n��O�1(��#NL��|��-jk])�sV�3��miyI���yA�F���鷍^0m�^�,}�Q�D��y�Ń��1z	]7����X���]�eB����f���x��K�2�T�e�����6/3�����j���»t4�U�~��:IZuf�b<����t�X�	*zc|C'���ٖ�,�xu_^�H�1�O�y���:���
�Jǳ���evk��ىĢ�"�Z"~��~��~p������C�Ꜭ���X�D�����t�Q����ܵ%��g��䯸�ؕ��6��}�r�+�:ڭ��g,Mj���q��WA���ۀ;{I���Vݨ��t�Pj#xh�ʸ�8���Kb�uv�9mm�a=�v��:k��7
�P�"��v�/79.gU�4B��F���d0�u]��y#P]��=��2Ct���aX($b{g;�j����}�W��-�;�AO��)��n̺Ev����E/��8��RX��*G*}i����/�'1U���w5̬�,��o>��
h��L�爢�lG)4ȕ�/��(`W�|��j)%�?c*t������:57�!Ah�ܰ���ێ����K���n���˾�t��X$A5�J�(�\i��ŀ�]׸�Ks���`��vt%ﬧ�5���6�tt��+�q�3%��vrӭ\ɽ�n6�I[�{�ꑫx��^�]%w-�´��A2+�)]U(�F6�����tD�z�:/���/}	��U�n�5L����D��o�ur�Ⱥ֮
��9����4�O�aO�d�I��T�&��~����٘�F�Q"a��ζ��Zն��<�'�m��8��S�8�-�;~nvq����R�u��d��\j��o�&�y��9�����7���{���צ{�}�^��w:�Z����*�*���f��Z��Auá���ٶ�9;��j�Z�#.z�M=��	�n߃����@M�+�T�1^@h��%_C�ݜ*f�}���p;ݠ���ׇ�f���[ǽ��g�Ly��s�u����jƕ8���i��y��C{Ab�T
���J��&����m)ϗ}ѝ�'�]���>jtZ	�M�:x��/j��z�Y���Ӷ[�y(�npm�s	�U����b���~ƶ.�U�ԃ�����@Sg9%�d�����}�;�
I�?�n��5mإ:����'X��ިMn\��S{�y�6�K�t�G��Y%�5�<&=�s��z��^[��qy�;��:E�nsz/pGjI۽}�o���M5����ͳ�sOq�ĕs��[���drq���3���ynp�a��M?.�XT�DZB��h�#�q7ƻ�ҍ��Y�:4/:/M �=є�'Z�T,�Q�Ř��k���A�|\�a��3H������.u�L��e-I�B^�2i�%�z�R,�T
�>��&�T��xd�%<�9ϻuQ�K+8���SvjT�(�l"V�yƲ[*�/V��̓R��ξy��屰�����%��Ē��չ|�V={p�2�:��Z��N{�hx�U�L)�k5Av�%dWX��	l�+���=[�$}�1���k��X��'U*{d��-�-�z��m��G��-��/��PtG]}-W�F���U������8���K7'����|ԭ�Nm��T�mT���#2��S��T&ޫ��L<}�^.�q䛧�+z7��@�R�����ɡ����1\#9�S;l>+2Ľ��j�0�3�5n��t���%b'�MGqS�"�]�����a�&��R�-w[���غk�'�Mk�r*����r�vX�u�m�}ZVf%n�-YvM�q��u��D|!�3�A�D��V��żl�z��F�}�(U���6;ND�^
��nPtA��f���י�{x绸t"���T����zV�l�k��ڈ{]S��X���%J�[E�YrZ��� ��<|gOiA�Q|\)TX�ъ�]�TB�Eff���G�N�%Z��,���%��Y���e(���@�I ���oCҲM�8ۮ��[� ��5��-Z�t��a��^u~4�O����j�iZ12�Z��R�=�ܭ��������l���H+ufX����z�4� ��wb:�ZC+��)@M=� �]e��iG]��)Sr«H[��h=�vS�[�CQ|EN�iV�1����B�j�Y|���p=��/�	Ϊ�{8��^ThE��$m�+R�}�9m�΀M�:��O��s�e2GLkn�A��-d>C�^n�tht����v��2��@KM7K��Pv�}i��[ݲ4�����Dՙ�wo\F.s�l�Sq�9�V��n$,G򫚩��uFYͼ��Ų.��K�{d�HOe��#2qn�Ɔ
TX3U8��S�jji��}�b��ߚo��)�=�7�HM6���-��"Q�3��f�)r��ُ�ϖ�W�h�}y`�:s�@��ӫ�I��3w3x�]��X��Gf�vSȪob��ٖx�ܤ9)ay�y)�����ua^�����چ��[�a4n��w���56si�������w}k�Fxp�'��o^բ��
���(�i��$,#����njH��qZ+j@���mr/�T��cWn7[r�|ۧ}��T-ޫzΞ�de6�6�+d�8���9�����ll�T���2.)gBcT��髉+���t�"��a��z���h��w�f��������@m�Si.:ǉh��3|��E�,O׋��T_��:Iq��2�2��=�s�=�V�<�+9l�̩>䫖��A���]�v��}Kw�X~ƅL��[2�.lj<fhJ��κ&��]��{�X0G������,�Ϲ�x��+��i~#M�ь�"��ۛ�.��n잩mQ�݌�-�Rx�|���(�G{���,�е��wv�S+ �,U����=�Ē���Yx{4Y�������ʐ�%y�so��dG�s��X�m�������ɛ�6�wH�;�m�7������u�ގХx=]WAy�ˇX�e�����t�Y���i�뾥wӞ�Y'S�f:��f�Q�nԢf����s��=�e&�:xf�1��ގ���C�u�����f�k�1��ݱ�T(�r�ܙ�q�7�z�,�3��r�+C+��<�.�I���QQx\���>[d�i�j]1HK�麴�;Aۨ�/�ކ�[���w�D��\�Eh��VVd�N^�|D(���ڄ�����z����𗹶|c���C� �%U~���U��`�Lj2V�h��T1E���bfb�2V�(+j-U�PV"�E�-m��Z��Q��9e�6(�iV-IPQ*UQ�R�et�EkE��R��Y+�����%Dt�H��b
""�Eb��"�U�*��ZQb*
�A�+b�������TX�UPAX�EUQVETUDUb&$*"�#X�����ƪ�DUb����U�QD(,EUUX����**Db*����ČT�T""���TUb���*(���*
�E��U*֎P�b�(�*�,DU���b*�*�FX��V*��� �F* �*1Tb�EE��*f\X�"1��U�ȱX2*�-��U��UE�*���V" ��1"��**

1A�Q,�����,UP�EQ`�UX��Rc+0j*" �Q���2�ݱ�:�M���u���Q�'{���흚{#҃�Z�=�����˲��v��2.�6h���/9�d[u�u�.s�&̃�ѪI\���x�]ڮ�Π�r���twkן�:����vh��"���]��tvY�ت���n���o#���Z^ޡ�+�{�����s��I�ǜ�6��gs�*:��/A��W��5��9j��-��F����˼���w�U�aF����Z�=T$�S'�ߧm ���w�x���6���ɤ���H�+�^�w|z�PO(+D�Ur��������M�^kHf�>�D�0�ݵ��_����IB(2������{��	a��Z�>��x��v��N�����C��w�٫^J���{Ctv3y�l½��L�[�i/M�o��}��BX�+j��S�^}��}Xv�b)��pE�8��U��j�Ү�D��[��:��"����b��Z�h��N�V�f�#��o.�hO�GJ��y�2�,'y�
���O-�p���_T싥��|.e�sr�sF>ߟ�a��C;%
��Λ�>�K�q��HA�� ��/WqR�5�|��_��� %$�Y���E�R�j����M�#L`p�^[�3������c1w�~����Um�6k+>���>�	�;2^��@NfP2�ͫ��*r��Uĕ|�kqs��֦��4��NSVb_DvW��׭�1��e3(^Mz�^�y��:y����[��%R\����ҋ��#n���LNtB�i���j�hխ�Ç5k���'�hGj��.s��ɠ�F}�/j���P�=1������9HZ{D)�1R�����������+&����T"+�_.��[o�{>�nۜʃ��ž���T7%��
3�6șdX���o�}�5�B���^!�䯸�%B]Dƴ5h��K��To'�B\b"�ъ��	�m��+��}���3מ~�y�\o��w���KM�m)��`���;^wk�u���6�����7	���AqH)&Ύ����ݽb���n�ޥ�%ޡ���A���2[��q�V�r��L�,AJ��A�<Rw�V�H	�^܆�o�ɴ���>��y�1����6��f�����y��Xr<sp]�Q�K��u��J<o4ers㺺�	�9�eN�|+�Z:��\���MN/q71��|��TC�7hCա��B���ٞ0;x��	��[*n�9�P0���օ�Z�k�wU��2�\��e�ws�x~�1W�-S"n���y��}�a��"->���B��n�ci�轶<O����u��E�s���RZ��3Ƅ�:�i=C�L>��nW�:�k�^C��E�^i�?#xa]׏=��_�����sS*Yx%A��v�]s�fz��p	��;mV3w�iq٦�\���r+a0���	ċ�VȎ}�����e֊{�e�`q�)������}>ޙC7#��=�]y&5ߡM�m�W}6�6(>{�e��
���eJ��אg��u�}t�� ܥ
lŤi�*5�U֤�3�+�M>؇u�3M�S97�OL�@�l�/�Q��}*��my���ƒ9��#)�sl_����X�9X�:��-�d����$�m�K�^�����&�{>yѵ��7Y�˽78�5��>Z1U�7���@s+�	�R�7/��]�L~��W�>�cYY��Fy�AΙѰ��&��fݰ���,�����`���Lgj�(E�ۧ���m����-�Ԇ�n�w���H�Y�Wǡ���,ޛ�y��oG�lX��]/�'~�s�q�Z}�"�w�mg
�I���h7}�5���̄���G0��g��U������(�p�pT����ہ��M�>�U�j#��p�v��.{�ugV0f�ĵ�(�+�֬� �з�����(v����"��Gd�E�9Du�ᚬ�P��U�(*:.Dr��Tvh��b���=ޝ�˶w`îp2�uM.�t�ayA)e���<�G��c]��~۹	�Q��r�y6���[Jy�6�Z�U�r�f9���(e���?I8Y��w��L��s�/"z���HcNY¥k�3ގS�sI���_V7��!��w�2/Uȶ�wdm�+iX����x���L8��恎3��s�Kq�)E���qNf����Ϲm+lbCn���f|���b����\b�BR�ۭ��劗/?u��y������&�6*��1��B���q��E�"G�1�߲3[\���ܪL�7\�F�n3�^+�PN�w�_=�7c�����wб��]��œO����T<
�T>�pͽ+҃�/S����/VGK3x�XV�3��n��7`:�����s!k����Z��ÆqR�߇���q&�6�2��]�9�*d��#iק3
�;� ϳ�T��%�w��0D�����ҡ��ڵ��??�xB���_KU���f+Ò��3���9z�8#�7�Yb�&�U^kޮ�6�\~zN��a���1����L&��G-�:��{)��:[-vۓA�FP�y��Y0�|{��N%���_o%�=A���N���,�~��+�c������B�|x��*Sk������ΰ�D���N�G]Z	Vʑ����!�剝���r]�'�nɍyKB�U�UI֦9o�������V1EkD����Wx������5�cVB��D*�B�~d �nzq�ޙO9J�NS;=�U�t�c�v��u�q�Ks�!P����E�(t�N!
o�V�����~Wʲ���C���Jt��my.�	k�t���*d���(�wa�~�DP��5�y�R�`���-
��O7)�&i��e�b�9��ohu�Bʰ�!v��s4�]��cg���};/o��Ib����|��Np��=��1���9H;��@m�6u]f�jΫ<V1JT �_�W���^iD����E51~����k3���vę��d�띑�2�A�b���7v�DwW������0'#�UI:�{!�.�)���'m��[X���u��r��a�G:��2enU��0+�����V����*���>�o0k���q�E���Q��F���&ܠ��n:�;%�fQ������c̋��_����K(@j45L�ڗ���T'3
{8=�{XE�'[�r�bٴ��,�}�f�yM��x��zn�sW;�5���.�5E!W�Ɣyv1��d`�e��J�-��|�⬫��F�bQ����H���j~W{�� [��d�'�@�BJ��K�{�4���m�sL���:��g_�o�B:�y���ߺb�c�z�uSꡈc�3�z�{�c�D[�zI�z異9۔�iH]�W�����ο�M��� ��,=��j�Wj�z��1�́ٽO�k}�w�j��9Vn�ؼ���p�q�� �>�i���Nw�����+��ӂ�r�o#�7���݊QyD�]k� ���N��1@k�\f������ �Owm�u,���1�F�k�ƹ�
ޟ��3��QV��i�����V�my�[~ׇ_�v;�+���t��:�t+�<vt�4V7���1�'v�}��pS]��>����҃�v^�vT�@�jվ3sx�۠�r�+�����kP������7A��x^�Vx�wMǙ���ʹ��=�`��%���`bv�麒g��;n�z ��aB~�MB��h�E�V:�P��	�pls�!��<�X�'.���i���n}=�о�*�9F��O��.ʼ��V�Ҽ���*���բ�3�A��}	1z7f�%J!���r�6b̅��c٥}��$8!��ˉ���ƺ�����+�m�.���<�b�<S=n���uȜ�yuG�u��}P�r�a杰�N��n��׭�K�����ؓ��WH/�c�ѓ�>z��e�TxL=�i5䖈��u^u9�*����7]n�Y�].�u��
[D�v�$�V�Q��F����`���,ЬΔ�)CU���{+1����n�p��C7g7��8�G����9̇0EyL6������iU��<:�ؓ|i:�:7�p�t3ܶ�����3��Ag/�h����Gۑ-�<��ϑLgG�R�ݽ����a�%�ək�7/:�i�OS�F�?]��q}ip><�b�]�U��}��v�,������w���<����o�򵾗mm{ ��VP���b���:y�*5>�g�����bGJ�o��v�{!�F�o#v��ϣ98�w� ��J�J�I�|�u��3�R�3����c/�M䯻�����H�`���<6]a���ste����R���*F.o'���������ӱZf3�&!3�����w���VSV5\�a���ey�]�HQ�
6���z���ő��i�TQ
����lD$,>R(�cz1�M��c�I�5�{$Ms�z���t�aX($��7�iɮk���VD�k2��e%�M�USϹr�L-l]�K��3h׭�,��N���R�w�P=�[�8B���:�-�M�EQ��;��Q���fq�k�`��7��]:�7�b�T�K��>|nr!�7)�B��ND����&��fv�͙W0a����2�u%W[�%w-��bMپg�C7�+�M��+��ts�W|yb�;Kցӛ�x�����7��=�K�;)+�J�;�m������1S!W)ėr�����"��]6D�/��m>�Vb�6so���tV���^1�)�4%J0�@g���Wi'ӆ���4��3`�P>��{r�7=����B�bz-�O�K!m�j{[���^��Z{�w�_1I{�j�ݐ�ۓC�������Z&�V2";{:#>�e�rpU�z^�׍ݽ�8��X|4J�˙O'�ѫ$t�h����۝&�@(��ȩ��΋MM7=@�E�y��:�����הz�Li=����en1�6�~`�{���Ś��#����롵���	q)S���'�q���q�b:!�}.=3��y����$�9���3�u$�٤���-jkX�9�_b:P�^�={�{��^�]�m�/2��L`�C�ǣ��;��T.��V*�����/��ұ���߽�<�~��֯([|S��Vp~�=��ȣ�g'��Q�^�*Ҥj����oo���V�fP�ȃ�ўD��j����`Enpj����6�&O��t�{+m8pB<!�ה��ޛ��Ն�f*2��:r�,f�>�¹x��z�~}��i��4�]߲<���.���q�w�0����}ͪ�c3ק�T��Q�y�+9�k}��Fz�VB��D*
P�r��fҥ�繞�}1�)h�.���+/�n;��33��h-�1�a��+���
�<�(:��;�;#��v�n1�Vr����S�m��nf�)�w��կ%DL&�<�ܱp��7����5��b���.�'uP)�_�΅�\�Fa<Ǒ`H�m��M�8ݮ��S�yC[�P0����	�n�<�u��9��1T�$�@p9?r�SFW�do�삷�u{�
����4�`�#G���Vg�ݙx�Z��k�d�U��@e�%� fh�Ͻ���E�K���k�J�<��^x���Z���f�^�)e����7R�l��'�c�x{�a�7�ۭw�ug�V2�;�S��.�L�59ME�}�N_{���3̌��2�,P':�F��:�z�ʾVulDó�I�+�O:�fV99]S���!��-��m����s�fY��6����n.Ip�{f������m�[��]Ӥ]�Px��q<��%��t����6m�k�l���*ǝn�x�yB���&:��\��&c�۩�^�PѺ��nD�ͨ�.2��J���;�
a�q;��]z������}Q�w[$=&d���:oG_E�Χ���YU�h:�����wñ
5`w�|G�{�5��"�s�y���Cߕɚ�uI����tr�?z��רY���n礗��N�E]����j��$��.�Q[��f�[�<�Ǔ�=Z��Ei�ze�Yͮ�.���2���Q�M�C��,�y���sR��;հ^���lX�l���ǘ�;�e����u;�7��+f�J�e��4f>
��p�]��>�j��,���	�s;�Y�ب��V��
Q�f�U����u����k��rc�GYi�=�$VX��`��Ċ�͓�B���i�.5�H+Vi��o1�E�����Z����.�@и-��Q��77k�[/�+<��
y˙h��Q;�d�0�:���ݑ�y����̇q1��lwQ�]�C���&]�!�ޛ{�;uw��4L}�*��K�9"r)��S�݋zv^�2/v��c�1�9���Eѣ�2=�[٤G%t���(S�ux^�;�@�r�L�Y�q�K�6��q�k�Ǉ��J3�!�'�M�g�}��0f�Wn�d�sD��5��olo-�}�v��y�<P�cɪ����>�4`�S�������`��]YܸI�p^��Ld�T[F�&ep�ci����я"P�&�1���7��|&#���F¦�bf�QDL`_-8!n� A��7����������E�7b���� `Wd@�0C��t /X[5��� ���x\,�H�B:时h@0]��sp�_�l�� m`�T�et��w(�1��ڡu�'[�/(ٯh����j�T���Ɋ�w���,,�݊FC�@��r/7JN�혵�T�sY��&�m4ף&��	Zqm�F+�����1˥3r'G��0��;����l"��gW�hY`U���#�����(�\��
z!�D�[�LI�ۼ0��F�F�m�ӳN +���-�Kh����&m�UL�`�R5C��WRØ4eJ�e1Q�a�Mu ,L��Ьp�9A�]����pm��!a��pgbӶ�e�3�!D����3E�ܴ��8�ֶ{���b1�X#Eb"�b*�2�Qb*1TQ��*�*��QUF��DDPPD(���E�PX�ADX0�b"�1X�ȃ"��P��(�"�ƪ���DE��QX(��Pb�b*1EQF�&5�
�E"1VDQ�Ŋ����*�#��R"DEUEPUb��*"��*(��,PU���"+eX,QQ���**(ֱQdT�*�X��1Tb$TT�X��*�+���Z��,b��UETb�A`���QT��YA�**"����(,���"#E���
��TEE*�Z,Y,����V1`��DQTR"�����b��"�b�X�QV(��(V��b�Kj�����l,dU�TUE�QQA��X�E��1���
,PX�1�X�mj
"� *�((*2#R�F"ŋb�fZ�)TX ��UH�H?	�$��@��F�U+os;��=��
��Y��6[:�'����u�A�����n.`Q�N�i�j0U�� �{�X팩����}��?[�3��m�<k�4Н�=�$J��5d��n��%o<�9��էSju#6{^Wz���U�:��k�Y9C��@�����y��������g����Fϫ�V٪�Y���.�s�>��5�6��s���]�Aa*���%��wϞ=�3�$߻����.+=w�^s�#�zrqX���T�.���'�4��SV����׻��-ׇ��	#v#�D��;�Vְ�6��9Q5ϐ��5s¤b]��n;z�½�~��w}�3=�U�4;P;�s��g?�(	\���j����ݰ�8��v@��L�Y cy�G��m��� ܒС=�X�����An���^���W��B����+�f(���ªc��տ%A��Z#�i
�����;��}ы����ʃ$��CX��Ȗ�y*BT�"��]���s7��;5�Y��z+Kf
�մ���u�=��GÅv{rQeo���L���F��+^a�����W�e�;w�s�I�W���鳛ӒNn#�!��uԱ��ju���]ٟN0\��v=ǭr��&t-����;���u�L��|<<�K����n�~���u�2E7f�*Q�j�ʆ�Y����(H4���.Xnm�c'�{V����VهCn�y��/��b-��q�i������Ǽ3xi.s��ݵ�
���<�c�	n(9�R�d�t!��5u��v^J-������ �vͻ{��i-&�T���J��V�r�e��ݶJ���6�I,��_+��7}����]x����sd�a��i%��������w�e̪��p�v Ub�0k�޷bOQRXo�ݜ�m^O�_?X��:�T�}��1��hT~���y�jR]�Pi�U���M�=�O�U��f�*�w��d6�v��.c9<G��6���d��(�b�ے��	)=�W�I�m����!%��[����I	I����߶��+K�zzF.o3����oh)��U����.�/�%��"����~>^k�����
���6�����77���2Z�4,r��f0�����r�>!��>�b��y�K��u����JS��_+���0y:x�)gV��Muwc����Ak*�}צ\g[n�<Fܥn=��],`ϺF\�'���[9+�>��ݫP���d�;�w
KL�����T0�z�p�	��2Q��:�\=iv�՛���ɬv8�*���PT���0���6��@�̪3f]����H�����kY���§��͠��DjB��S|��7�wݣ1+�4+W��g9���ұ�0��l�J�6�[�T0�T�1B��[�c�cøW�Ld�U[�J��M�P��k�]
�n�F5�C�=�c����5�Iwz�s�1�p�e�[��S���[J��׾+iN;����U��%����f+�!��!�[fD�ɬOhhW|��eT&�
''��N)��o�U���y�tȣ�uF�Ɍ8�eb�45gG�O˶��e�??n�� }�R��z��.��K��u:�̩X�ŐqΞή'km�/&����7�U*�˯�� }��_+&��G[/��t's;鱈���?z�iLy�B'{�sY��������f�����2MzO�z^9Ea�:�ܱ�]u�%X�����Z����`Xf�f{�V��*�+����ƣ�]8��5.!��Q��:LG�kE�N;0�<�8�5m^�D</���4(;�X����{�}�F{q�uk���'��K}��yt��{&[�T�`�r�f�+ju�q$��,w�J�H/c���VNb�jt�#y�%J�]뭗�.]�a��!3QQzb˅����,�Z�T���m�߶�
+���ư���w��"^���c�9w������7�@�Nu)�tƬ�Z���ܞt�5��Ջ��v�:x�k��Z���P��^��X�ʽe��)��Z޽�Ui=�z;:�>}ʞr���p�<Q
��@��wE����˝o����b6���[�Av^ �[x����=�gZ3�P�5].c�1�Цw�[v��30W�u��Zꗍm�}�V�7)�m��o��A���,ڛ��c�o,Y��l.s���;��}�΅c���!�-o@qx�(ﰳ�sG�k8m�u�nvDX�]v��@�n��Ǘb/�pO�Qy+3F士	�*�9.��g,�^��78��{40(/��b=k�oY
���o�IN�-o�pz��b���o4ү����C�3�Y�\x���<�i��1b�iL��e��3�A����Ggi��59q�BoMzzc��P�9�ѹ[�/�w��U?�J@p�o*z�Ǿ��Ӧ�x��U2#��)�nY}�e˄�9#���NU�8E��a�->��x±��P	0��mh��CX�MԾ)�J�Ֆ1is囩�X+�}�_*�GϹ��j����#m�C0��W1�y�J�cȒ��_y�c����l*]C������yd��%�6�B�3�2I�oZ��Q������f*�z��r�1=45QoV���\�%nv��r�����+ӏɵ�S��׹[~����8���l�ǌF�9��̮�6+7��Et����}�^�_Kۍm]��ON�����7��sP�ݤ�O@+_�;>~�[�p���>o�Xׇ�,�Jʃ�6:��t_+ݥ�iĆ]s[6W.�}h7wɾ�v������!�0�S9���֣M��V{��n�sC�7x�Kc�������1�x�csoU�܋���m��Ϊ��{�z��xJ����Ym(��j��2#|���ψq3B�k�A�����=�:�u��w����Z�ŕ�d@�wR��O�5ynG�6��ݯ�z�:r����{��:g����%�B{�=����؂y~���t:����N��+��!��ݦ*����<�����]���\fl�g]D��]�����cה��p�y.���ZBek�-��;�j�*�C��o#7/9D���گ��M&��C���J��"��]�����OB����1tvk��ZNн��6�N��Q��ά����,m���������^􋮫�x�ծ�[H*l�v%�f�����[�1a���z=>�� ��?cBe<���U���:W��LOH��D�vn�5��G15:��v��c�]Cә�%=����:an�ܘ|��OOgA
F��wC�9�M΋��oE�tONyθ���ә�%c����>��e�5V���R�Ǭf�ڿ%�{*�莺s"3�kk'+�>��\�̪L@�S-�wPQ�N�cc�ru�Wb���kM����G\�.z���b��=� #��9��:[��F�}#��t�d�����Gg�wN���.�ӎ��M�:���a�8 v)��K�ֵ܁2��	�0#��7o��P3��vq�}���Yݗ���F����R���כ������\Wk�Q
Q�9�"��\�94�B-n�׼�k���S�kq�7ϊ�e�"4{,�.��9�E��ݯ,�=r3;q�U�.E�jRy6���f�^�R}�I�{��[�2�ODx�A�@���Tu1�h��g�sw����oHc"b��������Y�ב��1
��gdu���Y\�U� �:�Z_<���<���|���ٱy�<Gw��n:�j!"��v䔅	/���~�(�2�؃�9�w}v1��ieD�����wo��F}���c5�>�m��F��3vf�<� ���Ro�Z�;��_*��C�KX�J1��)g��r��r�v�31s.��D�䆗�}���c�o:�c'�ݚ��f���tUM<�2��x��}�(��W^��X�ՠ��p��_�x�X��"&�w6�b0H��#춛�6����̃ƞE>�W�ö�Z��<���I,"uXQ�<�V�h'Vg=�X�^+����N����!�bw�(6�5��j�+��:�R#�> ���n�J�q8��^��3��,{*�r�X�V��Ia�����7%/o�QѡoY���W�::<tK�yoy�ǫqw.(v�O�I���x��[��W1������įL�{��{|��֪����e�avC��̉[�X��Юo�:��YD�m�$z+]=�����g)�7X9bu��g��#i�JwJ�=Xm=�����ռNb}���}~*m���o�ə��6�	�ʕ�s��Tu�P�J�i󙭽Z�-oHڮ���]<���O�>Qf��G] �7^*�	�I2�R�B��V:s�5��1�ݎ��~]/i�n�>��cJ����>��D�cG}�e���)��4��k�VNV!�PΔ'y㰕+iC������(������y��3,���-���Cr]^�#�sٹr�6�C����,��RG���M�%|�W�-9W��U��a*Q�M1�km��}ˬ����F�Ź���4���sD=�X���N�K{U8*��K��=MnN�U��9&�ݷok��/^Bx�<9�����f���c����Ƈ^���5�^�~�׮�i���k�������T��c��1b�u��{�N����K�E�Fe�b�����4���7��3ux��])���\��� �m���4݁�=�g��s2r��-Yǲ���`�}��-uz^:�ҽ)�ݢ��7
ng�ɨ9on7��6 ��aIc�ܫ�x*A�k��Es�]3���zC�R��н�NZ�d�= ���N�/{��Ǫt|�_i_�y��\.�����]ϢTo5�_B�OE�52��o��tv̉[�p�X�b��g����B%<��ќ�����la�q
Y��n�.�:}�Ҽ��ׁ��L\���ЮGL9�f�&YV%6�O���5iٕ��Ov}�7�.���:����y��ElSI��59��Wº#OF�Op�������LLn�����c�2!���U��n������zy���<�<⳴��	˾1��m�
�������J�둸�D�{��ŷ�v��$!����C1㜗y��3=ax��ŶT�o�����/%�T���V8�3�Ǧ��Yybx
Ӌ�`� ��q�@���o�����;�W������Xλ�[��Ρ�ۦ�a�P��N���Ȍ��dt;kb]�N���u��_Ϗ��<�_'������Cm?e�K�a�۾��/%rn�)sw}�#�O��5M��X�q��_M=��K#vÛȣ���vB���'4��o2D���.�`���J��#��oR�E�;Af��^�fL�oZ��Қ��������M��v�����e���kuf䭗� $/��UEC6���;ݹ�_Wz�����-�c&t:Ŝ�;x�r{�c�j�Ņ^;s�R���]YOiݓ+sF_r�V��I�T�]�-��7|n�%��x�6a!K]5��Z`�w�î��m3&ݾuY���a1گɧH��L�\������ӅS3��-�%�w0obT'u��I;�/c�6�vjT�(N��雔����F��B�A�����\��X5녲��w�v'ͻ4�f��We77�G���n>�2;i8�3'�'�hf��̜(�7���9���܄T��yt�[�nw �QD�\;�bi��o�����T�Φn��ƅ��)�=���C����m)�vu����J�wB�'��5����S8���I�O<���gdL��3&=�?+;D��5�V�γwC�<8_#3����v3C�Q�k9���]&|�e��q��"�����f%��}w�z{oe��(��3�^<�m`��n�o=��c�)U�ejev��I�^�n�B*�����11PwY��)².�o�p_یi�u5Є����qf�W9��eL�u׌iGJ��59w
T2p��ֶr�&zͧ���M��0���]���<�ʍ(r��=�V�T4C6-���Jp�'���[IVм�ٜ�G��`mK�$�y�WQi���п�u�O�N=�u=�a�������5-ޤ �'nop�P���V3���vs����ZNGn�a�Y:5 J��;��k���vtU��殀�����4$ɽ!��b*�*��oP(j��`���Mc�A�|M�h�R�����F����Ox�G$������
h��"ͼ��t��xd�YI��CR��C�����iv8)|9ύv������es����w��jJEr���2*����4�꾩�!�К�Nެ����@n]��`��9�&���\��>��^Z�2l��k"�].�yʻ��������L�h����4:�^��E�E���g�N�&�cUwF���g;a����0.�P��b�#aR��yJ�gT�w�!Vl[�4�u8��{�ף����|@}6��*�Y���9c����p�b��}V�_�#t�@vrWQ���ˑ,N���0*0z7�������i���7�$��Փ�VtbW�F�*"#q
Ên���[b7KB�))}K������TL�^�5�ں���?#v�|�	������sfݻ�U�I��q�t���(��l�Ã�uO��bn[]̒�m�o��#��is���Յ&����W��pV�WB;���+&���%u��܀�8�
׎'x8�X�j8���ŗ�s�E�HCa��Ҹ��WV'�=.#B�5���g��''��\Ysg�
�u>���.����RoC���<W�ҡRRnjEc��%q��Ⱌ^j�C�#3�+N����>�|�*���� ���t�=�t��XR~t����L@۫Țҵ>W�r��n>�ݥ��
���[�z`-u�F��V��ɭ�κ�����s	h8�q���hwFszޑi�;~�.���h�[��,V5�(jT�7A�o���Qx���zAZ�+�#�8���|r�&vnP�9Re��R]Y��uAL��H{+wV`2�u�]n�+"q�u9��P�x4�Y��4�iF�� 8�Y�k{8kBS��t���s[��Ѝ��q@�Z�SC��xini*H� �Q��M���|�@�d���������ɔ}Vx��5G��w�������k�����N�C��	������-�P@g]g�x�{�;y�O�y�s��`�Ab�"��Q��dg�E��,U��AQDQb�UDTEH�"1��"�Kh�1b2�
��J�V�ѱeeV

�F"ţDX#�La���q�`�Ub�1G-Tr����%���amƊ�����Ab�E�b#(���Q`���A�T�QA�IQA�UX�E�����R(�b�[�C��DU�"�h���Ȫ+X������ ����X���V�TTAX�+�*�YDJ�+���(*�#`�EAb�U�R���PX�
(#2�DdF
#�ERH�b)Q���Db((�V""�
1X(��11����`�
����j���"�Q�1FE�X"e�0DX���`���Q�����S-UQEKE��F(�AATQb*�V`�DUQUA�?c���N9pfM\�彮�Kiιo$���H�J�����Ka6��!�2�� ���ιԟ6��a��W�-@)i�}�E��K��/���b�ϥvMc{CB��L)Ε�jbzGj��ӹ��z�|&^!K�h��<̧�γ�<ךiv��=PL+��OvZїO��3_�M׹ņ���r�h��fdʷڮ�b��[3�o.#��Q������;C�T��휴�ץ�;���%�|zjŏ &p��k��ջ��R�s	��F�%au��o�w&�y@s��s1��g��LK+��Mh��`5�#�-�C��۴�um����Y��6�`l������k{jio��������|�R�����ooZ/�wo���2%�� �[�͊yZ�#��;!�
s*:����~�V#o0;O�z�UIB�f*k���LIOa�r�vl�����[��#�5�@���TV*'=ѝ�o�gF�\��x���%�#P��|�X}�u�.���m�*J
�����|�b��;(W3S��e;��.-Z^_N��cx���c���ۂ�G���r_5�u3o[}µd]���w��tv�0bK���7�b䩷<�p�Ĵӵow<ֳ����4�I���t�s :@�"[�\u��A(��T��e�x���m���l�]Ƶu�'��~�1��y��y�5��v�V��2��hɶ{aEZ䧆Gj��n����C��ז��.O����1�)5���R�QV����t��-��N'E��������ڗ�N����Cy��c"��y-2uwn]���aI}�n�ʶb̭v]���U��B����K}�9��sؚR�[#��tV{�����a�=`C���b��� �(�'��SW��d�-��1�~n�*�ǟ�U-c�eP�G��^��&у��^�.^t��yN��g�D���G�i"�10ל+�y��o1����a>[{&�8�N�����/ھ�B���]l��V�k����B�`'�|�l��Du��h���0Mv�Pe(��]E��ţĭ5C/ν+q��]�y���y��>X�<}��!Nd�6ׯ�Y&�AC�"*�U�ͨF�*!�V��.0>�h�[���n�_b��8�=���ǌ���3���sqe�j�w,��j��ߟR	a�|@e<���~9@��%�9�"�� ��;ɒ"�Q�۵հ_o@��bl�W:�0"�;,0E�9�����u��GGvtz�}[����[���4�+���N���w<H��,�q���4E!zk�8ݚ��L;���21�kx���F�V*�{jxt>�wj��)����p�#.)�x:ͤ;a�{(A�
2#�B�:�,@V�oA�?�+�RW|q7CsK�����=��zˁ��������W�(�9A
KGΑ�����op�u7�Oݞ�cV�k���CL��d�Byk���2��'��z���N��[7�p�<��tv<���/������>q�Z\D�X�������ïk��V�ۃ[�Ӌ<=�33�AȞo(���ة�560�@��u�t�Q��X�Ǵ�ǵy�{�O$���4ͩ�c;ґ�P��f",�=G@%@u�(.;h*n�3g��u�<��#���מA�{v������z�39�=�WX���^3U�V�@`!?p�;}�˫�����1���Oҗ���.��┬���s1K�'b��L�v׏��A9�ް������2s�Q�cމ|��F�OE�/��%u8��`v�[Bx�(]�rK�Vn���%D��RH��Iً���~�J����m�D�����f,��g�Ō���*gwY�MO{��[/Mb'��A�%�:5R�Bt���{|�z��$������1�p-��WH��5��UJ�h��M}��=�$���%��qR����֧K�����4�1��/������<�p�x�, F}��}M٫���/d=�X}r���>�k=T�ئ�h�g��OrDTۻa�!9��s���)A5qp�jL���>W(�,���T�7�v�v3mu�
��۷�/�?Ԑ���b�9���B]���ƮA��o(4�Y�x%UV��9]&f2��PW���`�N��;�W;�
�1�ݵ�[�w��׶$6���<u̘�#gc�Ê����=��m�!��Ag͉��5�h3��������Kjs�B�y�.����mU{v,A������a�-lr��:*�X�����#���v#UPQ��n�t����8�'�Py�}�6��^�#�C��8�KWba�V�4U}d>*�ؘH�jt�Q��dr5�`9]��o_JI�z�!o$�kW�F˲N�Eż�cl�W�b��CÜ��U�b���%�֭��L��]������3����e�QS��X��f�{�U�'�S��^����@=���l�G���P{�<����i�Օ��zٹ����J��K��Y�WW�����`���.��ӥ�7|a<5$P����J�nv���Iɤ��m��9� �Rw�`J=y�g_i��)>k����Ȗ�I�U��5��ܨF��O�:U��(CX<�o:�'�Ւ^v�c6U#�J�[��ӑdG͞UF���'��~�K<lyǴ*j��ʹ��b�`]������ł�P��
Ī��Iޢ_	�i����<N7Qʮ�X���	�ߍ���JgP�-��(l�"�����\���|��d�A�0�%�uU�ҽ*�>�DŤ�f�xe���e��Cإ�Fq�Vʝ�Ϟ���ڝ�����ݼ�z��Ao�y*�hÍ�Gn�S��x����l��3eC�	VUZ��c���Ҭ}��
�<���� ?u�������k�(<1"b��ؓ�7A�vVx���5}z�*<hl�qX3��%�y�yF��q��ƍ;
7Վ�TT9���g3b����L(cN�l���%șɈk�Uyd^�ҁ�Z�^5G@{l��E��;���°++�{�Z� �Ȱ�>ޠt&e�c��=�+~�b�v�ЋV�뚢�������ҥ_rHVV[ޤ(n�p�gp���T��x�7��>z����e�X�.v�����_p/Y��ڛuq4�l�d��Ms���#���D�\�$��/�)��Kη��W'_�_}�ۊj��7��x�Z���P��Wx�;���Ӛ�`���J�ٗ�>���R��sbƂWp�$��Agn�s�����iwpdz:wke#����z����,�{@��e�6>�e��?L�vq��>���I�*���e@�	u9����	u�xئ���p�p|�# �����MՈ�<|����-��4i��J�Z{��A�XW6*�i�!�-:��Z7����A�뙺2?q	���`w	��v}��;<k�����M�I���s���IoJ$x��2���מ\م���-n?G�7�p�4��1{�=�&���:��^��$�B���eHvE�|l��2�:�w���1�5Oݯ������'I� j7�shZk^Rʊ�_x��c˗��sW�|� 2kv�'Ć�@Q�ݗ�
��W)X^uC�}y��.��(�q]��*;3(�x8:慁��8�O{��X�:|C�`B�|��N�eOE#Qlݭ��n�j�{7nAck
g���5P)��b�|��ĉ;]�(Wz�41t;cD��Q4^�1cǂ�Tw�U^�fDMn|������l�bѪ�<VC�"3�2��2.[ч���Z��y{,J�Tn!Y������Y0X="�f�L�n�on̾�> H��e5B�u����m�^������|\����~#cmy�:�Y�Q�7�7U0�D���\���B�;0������:�*�5�֡�T:�l��dd�*{��+�tԳb>��l
�|�>���l|D@�S�aͪ���S�^�u���,#`��/E��nˆL��>�!����uT�y��dc+.��I���},��=���v���CP:�c�#����9�~57��o�3�z�@��e��%�q��K�zt.�OM˖��Cj��/� ����ꍑ|��ƌ󄞫�m�ْ��=GX��
-e�놽�ˊ{^]��%y�����:�5��@�7Y��ۓ��
�9>;"2Fc�����:Y�׉��O%�C�	϶�X��*�h��/óG��h��m�����Y��Ή9��m�yMẓ��f'�GG����d-<2�v��`s�F{��<��.�Q�� =�n��%������%"�M��
�n�8�7�������g$�Z]ēM�A���(��aiGyrA>O_�)c�J����w�q�	�C�t�Q���ǀ��ݬ/e���f�\���a�O|��
��L�S�\��U;�c�U�ؐ��"GIg7X�;c��n�'ʪ�gǢG3�
eP���<:�^���H��\v�#�����{�m�tC�Û3�ݞ��Vzn�y�8f�ޕ�S��*\T���Aov���[|��im�=C����fQ�>����K̖��[K�&`c�@~#��fYBj�ۋ=V�Ȟ	��]�^���K�҉�[���ą_g;�d�j,N�Ī���}�$0OZY��:�'��"������#L��ė�h_K��7�\~`Nf.ط�L��M���$����Ά�d����
9�#>�q�/�Ak肵��/��&�](�@v��]���E=��qw��X�����1x��Uྷ�H�����}�9g�<4x0�]�&�wcs
\�Mt��ʶ��F[�d5�Tk��3/��bP�U��bY�n͸�QR�!K5�ϻ�X4��w	Nj��D�㘙�P���OC�W�����H*��{�����R�S��)��e�3��s�hH#v����y��⯱q!麏���nv������>��Z�j8�����ם���^��,9��km㿁
�T,ߔ\���vG�`�i�ԃy�/�M��tDH�Y���tW���*��l��%�cuW�۾��C��LggH��촶�n�O^u��=�� ��g(v[�h�Rq�J��}�m�bԡFq>]�t�'�<O��%N�ާ��}y%��r��"9,�ޜ-o+���*v��dr���Cþ|o<�B��6V}=)MټųH͉.�Yu��3�c�<~UAF7>�.S�X9�7-�3��ŕ����sו4��M����dYr����m�t�"w<,� ���d]�Kc����}����m��ڇA�@����$���K�4�<w��%��fϕ�.�J=�ԃ�2��<x�~��*f��@�+�>�W\E����#+�:�K�l�έ������슸[��'o\�k���������xq�W:��6@�\#|L���ޠ����l:N��J��:�R�����J��Y��V���dd��g$��[������U8@�.�17���ƨ��\�d����pwd-�A�e��=���8�Y��sE��{÷��#~�-VN��gQ�]�1��P^��z���q^ظE�1�燍�vg6��_�]W��f�N�o��J�y�}�~t4�'�P�FX��i�;V@g8}�߆�K�oT�f���\6�x,����K��G,Gxݹ�z�+��@�)�Ѹ<%�4�4�#�ݩ���5�ki��Ok ���փ+�5p����'���[�ßTM�-�Y�iQ�ggO�Q���{RT�x�Pk%�N������䋍�È��b��Hc�	�˯3��N�8^�nd�an�=A,Wm8�]Z}[�{�5Q�s���7�e�{���?pp ��Z��y�q�R�*�_p�1�[m�s�
��k��8
�R�4�CD�mq�\P�Y>��?p�����7tlj�p�m��E�'��	4��Q#:�n�7½�>��ňp>.!7��b(o������C���鵌{WQǰ�r�����}Y�(D�yP�0��%5b������=��Q;��ľ��x�3u�S��YM��*�\Hg���X~�ɓ���IưӸ�w��J}���5ϖ��H�*��jtߙ#~��6�b��#K�ϝ��@�On����^-��%��:X��}7��^����,`�W�����C�Қ��ʅW��w�F��i���L�k��=�z�C����^�(���������=Q��Vw���n�eu-9�06�Ay#��L3��U���Hq�7E� ��g6P.N�&�N>�x� |�Qc
��̵c+!q�;G'I�1Q4����|x�?���L��Gk7�F;K���. XC�LX���	��ӵ�T�w�wH��;��(d�d ��o� Oq�R޵N��<���1m�W�������;�nJ���CI�� ��C%��u�w(5�\�n���K%��4���nˊ��Ŕmf�ޣ5�y׺�&��&wå-y�f2kE�ƚ�֒�r�q�e.9�;5�7%�7ӤM׾q:���į�s�D�uWy�i)j����ݵ��l;��s쥇���F,��N�ͺ�ԝB䫣�&�l�;����ӈ�z5���K�IR�Lų��e�����N��,���p:�c��y�J��r�d���l��J���m�����:�JG��G�p�F�T�L��Ǳ�r�6��`��!�R�v��V�7W}İ�#q"��#�W7&u1�E����Sv8�]! +�n;�����ƺ��8��mIC�2G��{HIyVu�r�g7v�$�⃱a�ݸH�QMk�i-GAe��g�b%7�3ɴ�w���Q�{, ��<�91^�v$��<뾾�Oz�p��*>:�`κH�<�}� �bc�;�ǻ����ڱ�89�xް�6�7ok�9vN!<Oim���Pb-ذ���ԋuTHV�6s�5t��]�`�#��xx�����4�1F���w'�8�m���5O �(�`W�L�����OHq��L�{7J#�}�n��$.��C��;'���Rn�w�y�Mi�]q..��GV%�d=˸�m�Q����v«:v�~�>�DX\G�dݵ)�,A�ĩc^���tn�-4w@�c���c����wF8�����`CచP�!�ڦ�hݚ�ӚV���u`�`���[k����L�I�ھ��z�e�Di�Z$��S;S	? �Md8"�Vȶ"R
�The����8��t��a� ����CB� ����[zN��k�Ѳ�������O�/`�����ӟ)�ݎ0A��o)ۂ�q��DQ� p$����Ph���6M+|�]�3#s>����������M,�\(�a�ɹ�~�j�+U�*ţB�n:k�ш��י~x`ТW)8n="�8C9@T&� jJ��p��[
-Q��똥:�i��f��X�  ��D���ڬ�u��񉍘��W�f��ؖ����2'{HVU?��l�	JP�C�R�i�#e�OC��J������eR:&�%+�9�V0IR��Z�h���>��,�Q�\⻥�s6G/��у�Z�q7�hi��� aa��rʺ}�mu�M�%�w�S !2�qc	�8�(z.�!D�T���÷��5�2�z��6�n�:�3�����K��n�u`�i+��Y(� !��4A,�u�uu盾{�r��"(( �1U*"(�cAQE��j�Eb�DF
�EdX��"(��`��UUF*""�V"�2�"
�F��Pb�b�*h�֢ ��##lQV��1��A#b����B��*
ܵUb�VZ%��R�Eb�V"�J�,UPPQF"�(�DQ�E�j�F
*��d�TQQEq��U]Z*"�V2i*.��#`�E��QEƠ*#�*��X�Eb��j"i��C,�� �c��V*��QT��(�i������TrՈ��[`�T��QEEUTDTX�"�b"(�1EQQc�*�R,�*�����F&2��cTY"�1EFA�Dj�"ɈULl,�c ��Z�Ҋ�EX�Q�cEPX"12��)UU�"�fR�}�~_|�_�c��������I�t�=��+��,'q1����M�!)�:
�ꤕML&�mG��tXy뼫{ZFU��;�l"7k���{����C]"�(�w�����+	���
9���'�e⭈{�0M�SNH�ߤ(��'�X���B����������/�-�_S�Ռ��s�&���n8�a:i��6�[�c`����
ޠ��!H��?z�����5.zi3��4�/g�����D��vJ��?P�[&�}G�`�O�<rȷ֬A�ٳ:��r��s%�i�;�jC����	:�}���D�9�9�mýWθ�����tݜľ�8h��偾W��ؾ�B�=��v��5,�}>_,ϣs',��52�~ε7�ػ� 3�����QF0�N�aYs�[ciC&hl�oi�x6g���t��lXN�D�]x�Wkr��~ͺ(��$��A�d�PW��N�
˜��J��qC郱�Z\CK$b��.�\��fnMb;�M)�5զ�M�L�}k�Jh���C��s�7���/��<&�Cc�ˏy�v�5=�R���*�g/��Z@pgۿ-ih��8E,�zrU޽9^� {�n���ҹi�4!��b�qcT/k2����~�u��p�@�v�k& �Vs��:^�/�.�*B���ޑp��$`��]�Aϒљ��z���Qo�qK�-��ǡs���wTO-��}bU����O>�I�kh�ki�P0F���y�ueI�\���@XL(�1'oN����ݿs���~}�t��`zU(8`xz[Ӹ�߽m)�ݧ5��ku����j��x52��4�o��dvy�<�x��]f��7}��0��%�{,��$A���� Ӫ�%�꒸��Fa'**4b
�76|�t�r��^�u��V��};��+�iz�Z 5��A����+叹�S�f��3�*r��Of{�$���k�۴�;[����Cߕ8��r�1���9<&�]{R��{j��h�~R�V�3s[�����:Tj7���
�w��<~�D�pFk��;ڋ�>3P�
�wb��Jɾ��d� w>���ۄY��V�_���|%�Y��5:��+{�3��l{2�klf�{��-˃=�X-�g��\}���0!�Bĭ����xq"�$���d��&_���G��Bo�/p���SU��oq�W�X�$s�Tv�w8�<ݺ���'�K�1����9wsXhnG���F�xSƫ���|�/f_,<|<�"��0��3���uk�b���ؙ��Xں�����8��$��k�O"������X{���R�{<|D������w6&�mog_�ln�����E#e]�':C�����#NrY�{�X�RZ��}��,���9���w��(R�Yڵl��As�Ί���X�O�{Ŝ��e��,UZo\+�4�A=�54�����5�QX\�묃7�Q���z��h���];��݃�7f]z69�XUT�Ĭ��Ľ9i����(u�<�W����2��:�]I�V����a��;4�Eo*�q��Nߛio�[�v��7͑lb�U�
�n���ޛ�J7ރ�O���7��<I�J5���覦����b�Ie�̝�^#��L���f{���d�+8�Q�@�Y�΄h
�(ǀ:��ܨjgV��#A���z5�;�_;�m�����o�=�-G��[g`W���i0�����)��5�!ݩ�.�b��#,j��(��S��2�i,�>]�i���}��ޖ<E��o�wr�$mi�q����8����<E͆�o��y��M1Ě^���W/{	�J�ř�WD8�ꊝ�����%io�~��p}�q�G�ʈq�"1��N�V�]v��uw��3B�H��Y\���u�w��#�b���ǟ$=��� p�mD�$x�({(�q�	���k�ue͡�"�jI�ߧ_,��5~�B�� .���5w�4@�{N��S�>��	����xV�w/n��Svu���B�Y�mBx�oh8�)S�J}��K)7 ���b�Jr�VnWGdL�6J�5�uj�i��~���x�ɝ���~�:�?%7tb�8�j��1�y\j�c�Y.���-��м|{�s)��l{�.�3{����x�a����#y-�LPE�yf&��ͽ�	Ռ�3&uD6o���Gl�eN���i�h*2�]�
6iSp��<�S��.r�ˮK^���s7�1��bo�恈���L�Q�X��1&j�3�9��4�z
�^)�3�݀��i���v7��ܵ���j��Cd���+����:�η]>v��?�w�3>�|3���aXR����t���]�	0�_zM�a���^�S���ȧ�1}��|�[s��u�&e�%��1�N1>H��ck���%{я��B�~�r��65��cZ�� cbt����W��5�
��.=�z�ˈJ�t!�L�<��=��աg[n����0�zf,��� o�$��tn�	N�÷3����6s��a۔��ȫ��h�ƥL��Ɑ�ה��V=��Y9����%���̘�q����v��G@��OW����%=���h���P6�ڛ�k����
����Wf��>x��igV���.��81�W�+�^�@��Sk�T�J�{z��V�ɰ���z�[�9����6V���C>��^C�n6��� ��K�r�g/-Ky$����Hm���>aZ��t,�`�����t- �:=�)�@52���'h��8ꉤ��P�g���XEj��t\gU|T`�mK*,��U��	��1��۱�Տ"(x�N,�u/����=�v1Q5�P���;|n,�t�ut_�n�.�f�h��:��D;l҈�s fQ�ȵ~��\g���^���.��+�h%J,W��k��(��]n�A��=Zm�L� 9N�k��X���P�p��֞��_��'�+ΜC��֍��X�
��\�)�gH�>c�[O[�cT)q'�_�C��f�*�o�ݾ���b�T7�>J�Kd`9*��\�4��{����<�ЯR��P��&s1_.1�i�$,#H�{�|�FL�)P��
]r�+P����m�^�+-nk'��dA	����0��ݰ��!a�EE$�#^꣆�F�.ss�	���ٞ��܏O�_1�:�ŏU<�x'�s�J���Y�U�:�[��?�+�ߛ���r[�����G��xo��ٕf0vB�D�<Ǹt:q���5i���q^���3R$�ו��^ꓽ�-#5}�������1�\Ti�ӤN����ƹǮu���퓩���7%}��JK���]�;]L��r�w@�k�V�W2�7/9no-C
�0b�����y�W���[�y�=�~�bg�o9�Mʞ����W��,�7��+kI5:�2�]eB:�	C��z=�G�N��4�^�㧽,6�#�<�����ꤊ��ث��&2(w����(��\�ou�<酂� �OW,�F]��� ���m�����c��l[ͬ�^�d�����W��uח%g�\g!I��Ϭz��ԖeM��u��
5c���d�����:��"��0V�XA��𚬖�a�7kҒ�����m��e��Q�<c/��dv>ǂ8�t��w�eV-l]�o#ڈ��H��θ����������I����{R�,d���V�\�T`}z�s�j��Ψ�4�<G(�c�A�S'�=F��܎}O������_�:�؜��<*냇쓗�d��Uf��n}�1/fBq�ﯾ}���(�KV�-��q���q�G�Om���GT{2/ZҺ������G/�3��6N��	*����Z�12}^~���^��9i�k��6�,G�.]��>Yu��݄��尗X�\���z�rMＳ Ϳ�q/��e!��/��PRW;���gR�'{��ޓQ�R��ml2�Ζ2j��<I���qg��a��7�3߻W�e��� �2�_Dd��φi�tk����!�m�,�^+nK�7�Ͼ��dH"�Z$��F�M(]���q��,Ne2���8ތqб7�UȞ�Ȃ��*I�O�ѯn�&e(�i^��g��A5[�1���Hz���r���0|�Q#��:y��3�r]TΦv�:�z9ӳ����K�C�P��
�}��F�p�F�EZ��ʾX
���͑W;�x`0�zn��+���{��w��;�}��	�Q���/+�㘙�P�����ڰ�����T����1w���ѶF	�#^��G�bw�3�ZoBdlF���=!I쥸�i�Yz����cN�OD`�b+yֳ�Uzv��za��r��l�tZ|��8倻׳;��M��z�^;���\#���w��=B�}\Ij+�Ic�Nw�T�R"zc�$˚�#Ѹ/����;z�7���:���`�c�ـ���&J��O��ˍJ�ͼ�{���H�����{kZf6J��S~���:E|-	�����ȬHV`�;��WP���'��
�^	�<���i���Yx��yo����S��><����-�F�
뫸OE|����WNCB�]u�4y�����ϩ)A��#�/�5���<���6�pA���.��2>*�mmp�>�tz�vK��]��ڝ\�;���	��m���̌��![t!��Q�S���J�� O��=�d�����7P���V�T��15Z��>}�{NFz��[�êVG'5�}D�-�W^I�"�lQ+�i�꼈OW-�����S��H�����>���qC_k�7���e5"�ff����>�p�M�P2��U�(.#`"�f��=�Eƈt���Y#y���nzu<��dQ>6@�90b�J�W#�흀���EHl�����݈�8�A���#yEJ��ճ��nfT&*�W:�H���@�L�ֳP��.9���㇌��(Y�z;���7Ϟ[&Xv*:DI=�-����Y+�v��q�t�\sV��F���d��B��amu��.|�ߥM�R�h���Hi>��ő��z���[s�=��N����cVgÖ��ii�ݫ5�"&?�itIΘ�꫕S����5����Vs&�[­j҈��!㶓C��f��|�rfU�.��B���t��=��V��.e��FkYX�����`q�tEg���c�GO��[��,�����z��R�ap+��U��.����X�7�BcRaŵ�3��7�:P�Ѽ��y˩�Kd6�*�?mwF����\�Z�d�ۑ*ˏ� ��k��.���������3�/Ur�����Q�,xz�VA����J�yІ���t�d*a���F�������Nq���� u����N/Օ[��twH΁�*"��>9~~�(RՈ�<�*N�ry%�n���jX�VG����])�U��c�ORQi�S�CO�F��,1Q�0.6����Ws1��o������5�N�B�~�4��bSËX�g��M���_��1�L�lR���{����gW��l)�;�	��hC�зR/}\��3�y��
�wiR����s:�*��
�}Rg��Aܸ�UW�FAkf�b8J�AoR�U�t�ʹw۝�:�� IwJ��S�(V~�}δO��A㻵J����\!�I�|"��-龼�{�����ʸ��{�&V�n4+g jr�Z� j3�:��C���6�V.���əv@�q��N��c@Wƻ�Z3��{����)α.�U|os3�
����{%}q��\�'�CX����X�R�&+�!�=����j47V�]֗j�MI���)yxA]Lf�9(��[<�R=���*X�-�ev#Ð;}�`��j�d�n�c�� �wWoj�&����S���F���u�o,k{�Ќ�;tVq�b�2ޓ�;@���{��A[B��P��tp+��˟w��>���Pr�n,	Y�oF�J��UF�Z�r�.dV�O[V��:�}�k��;�Ƅ�	�4杽;*B��ymZ9�҉���%Ν��uR�Z�[Ճf��0N��v��~���P��[�oo��aưP��z�b��҅��Q3O6l�#h��/��{s6���J�@|��~xf(s���Q��g�wc�uӊ�?G�ŏ�/�}Q�5<��	��Ք��j�Π�Y195�B�e���^��z��P�}�Ձ���mm��s;�e���%��4D��Y5��PҨݺ�N߅tmؖo� g�2��+�����̞��wo�߉�����s�U9w����G֑��FO��S�/Usq�5�zg{���hG�������\�m����.E�����^y]�[.q�q{&	rұ��{w噀��/yg��@l���L��!]�\g
x�Q�]<=\��Q��4��x��g�E�l [�O�۔_����mt� �{�:D/�j�H�*�3y�g��"���#�;��
l������4���DENu�@���p�.��l��}���ю3�R[�xC�U^���Bz{�X�7m�H��%�EO���iҥU̔��Bi[u٤�)�+�7�%I�Վ�׫��vM��U��u%Y+)�1}�ҔTkL=� �����2p�g�b�d1R�	z�:�X*"��Dwv�
CӔ�sYO���tJ8��YT�S�m�#F9K*mM�b��Է�����q��,&�㝕��H2a�E��PeMV�)K��M_Nm��Tzs/t�Ӧ�gnf�L�ꛙ�oܝ.�������B_4޽�LRt�cL�lmo!P�WX3f|;Fy��R
^�W+{&�o� ڎ�����8�l8�QR���Ty�.�A&����Ȼf�n�Vv�|����N���>���OR�DY�-8	� mGww�4��X�י7$��v0����6S�b}�$G��.@+��ۦ���9�T����)��<�M?��*46�;���I��-d����Ŗ�g���3R�w�g�؎�z9yn�w�����o��N1�Cs��YRs��JI��Y�����9�֨P�EI�EE�L١�;��ZZ�Q=���7I�\�V�#�b=W[Z�<�:�eMHM�n� �+V�pX��#3Z�:��(�Ş=���0W
�(Gn�]X�h\�X�l�y��;-�<��w#�x����Y]�!�<���k6)KEdQ�D�M���(��{��l��&�;٦t�5�;����;��?-��fr��kp�[�YM��DgwE
�Ξ>����E;"Zdm6�S[ƴ���5KFv�dx���hc��KՍ$�ڪ;�����0*�+v݀՘o!��`�a�B�N��A�M�:���Z2�L,I���c�jx7te�Pɿ�ђi�f�5Zf�i�NX"�BslAj���]Ƕ\T���a4�;�(Z (��Y622捓�wt�A�2]�(�1^Q�JK�&a�)����	��">nHq��ҍ�q}AÛJ�!Xr7��mT������$(B�/�Z���	�p��rS��M%f�*TӲmPi���0l`�R,�1�B���$}l�e�g��v��PjD0SrKc�����4�0�4��Vjsd�ݨ�b��H�YԺE�K��{îѸ��j&B���J�)/{�t@8D<2b��co"k6�A��/��Wt����vه��f��ɓ�k>�o�+�r�wɹ�FAa
�8K'���5�+����OtZz���Oń���V�f�	tݻz�V6�=ѿc����w4s
sիp�%�ô5�=��	#����@�*��PD�Q������T�EFV�
�r�E���#��`��ATq�
��(*0QV2jʨ(#+X���6(�X"���V(��S*�CIEcTelE����TPTU(e���&61F�X��"���*��*((DDb��("*� Z�(��X�E���UDEF"��cM5QV
1EE@GMB*1jf
�1PPV1TU���")�I�Lb�� ��"����媊�(*�(��A`���5lQ��E��TQm+E��&���PF(��������AdEAT*(1E��ER"��(��QEPETU�*�%k*"i��TV���WX�KT�EU�e��D,�����J��(vm��p�ֹވּ��u/�&�G���D�f{������Wr�����Rs-^�R��6��_+#�晖��_
�c��L��W~���"�V�����$��#�< #��';�AJ��[j�!�j}P���������Q�Q �=1�;Q`�c<}�MY
5	�|�f�m�J��&ծuQ1�wR�9�\{H��p��n��X)'A�K
�崰�^��2iX������1s�(oX���O"᳢�AT-�9�>}��i��H��#}�r�7�ޓſC���	'�O���(�5�!�m����~��M\���Q�������s8�i�9�h�6e��	ީ�];�q��B��y�n��Wd +|́�t���y�y{1��#�R��)*��^;>��-���n>��<g��}�@S��srz��鋺��ae�䍰}��F$��J-���E
C�WK;<�٥��f��~�F�
g\!�� {�-=�D�W���f���ab�$�x{�.�kH'uT�5Z^"P^9���.uY�8��Ʃw;xelFl�*2�,�y��61�t�lOpElI̠�^���n�`���$,���v�j��4�)�N��&��K��ϝ�P+~h.�n\�b��]��Z7[	b�5��Tn_v���ژ<�6�ד˕���jg�nڝ��٣�}�A�ժ��wg:�{�κ��{VӨex�I�|<�8���퀾���k4�`�4}X�������j��V�s���9Ѡi�;��w~������������J+�Mn۰D%P��c�N�>�k�T��]}��w`�Jy�"Vj�Z`>�x�3��O�7��j��P�7��QW���UAF:�n��ɪX��[��H��<+%f�Zg�zr(_��
�ׂ4�Ǯ%u/H�A��:�zXúS��>�*�=�)�a����n�3@<�IF�Nr�����\[���)������5���}���׏��)���v����XUv�t
�|ڢ�QS�qP0n������f�uy�yI������jb=ëH������NK�y��дG�2]�尖��Ǻ���(dn��xmu�[���q�~#aP�.�����V�#:��D��2������ʽ�z��V�MO�@��CʽE�}���6v���
��A�e��=y��R.�<��5py<6/j���`���	�'ʊ�����s�b�^�]pgk������UmG=y�׉�QE�{��:�f���t���~����{�Hz�0�����dBi��4��Ȳy�M�*�|rE���T��w�A�Ng�������1�,��G38���{��U
]MŶEE;0��(��=Q9�Ȩ�򛑩䪾*�ЦHFz�d�l�;�J��Y�5��a���ӧ��i��xw�����}���l�ewFi�u���(�%�~��"ii'�E�BxS���ڰ�0����;�9N��5/��A���%ގR�~Q�<���ɯ��aNwgPG�VP�1�P��º�R����ܶ}B���E�L���|_oo�.����^k	���:��H���yG$su�ۨ��o��xE�HZlF��f�&W�X�n6�ϸ���h}�^���X奀﮻;&%[��j��h�>��{�W#b��C;~���C�d8����1g�`�ձ;=ZI�f�t�b����4���Ɩeqx���K�<�Ȩg�_{���F���{#�<w��+~�<#Ƥx���Jk ��E�.���T3�:t��}g��e�*vh���[��n!L�^���y]��lJY�;�	O�Z{B?6G�X��Y�(xܪ��܄���.c�`Nb�n}���Y-��N����-=�����g�=��w�<�7�U��u9��}ь/��)��i@�㝁���@�g}�y�E�p
���W�p٬�+���)F��>�;E�MOn��+*�������G��b�[�[�����j3��ѣx��oj��jN�Q�ќ��,2c��*&^��7MrK @j�a,7:�q�-�5�P���4�Y�f-�v/%a��rT��I��Y0�3��j���ꊸ�D�R*#EO"�z��$z6�u�B�#�mHU�Z�ޭF%�}D�
��d�]C�,�E���@�H���$��UA\3��v�5���1R�����ca{�q5��t2kl����}k� �%O>|�4,	>bzz�ՍU."b�y�y>q�Q��>�j����OE#P��n�`T�a�uTlz+�\l������:��}�6i>m	��ź����!��U��ҏ��P�\���*&�y���w��9���!u���ǁ΋E՟����w�(Y�36t�Zn�b�ch53b���S����0o���.��ᵅ���<��狳�Y�簚�&nx@е9yCcvv��H�?^U֏ݍ���[PϿ~�HQ���E���U�����rb��S�UK������)�Ϡ�jV��&sdtuT��~� ���75���O�(u�T#�S�X��og��L�N-���p�N�öq���3�0�ĉݶz�^RH��j��3X��t'�u-e����M�hs�0�1WI������j(J飏VM}e_q�x�ŭ�+��;f R�VJk^w)Y�z@�y� ��h܋[t��W%���<�{8�{u�8��3^����(pN�h���)�c"���n��3�,y��ްyf�X��C��Ш�b/��7r��7��O1��Ӷ��5�ǁ�K����V6k���l��<���kǚ �~���ZG�������B�<.ˁ��Wcv����ڱ�����ʐ{�geI���Q��L�©1= =C�;ϱ3;�}���i�_�D5Z���1���zsi%Y�if��w�,�\`<�> l�s��Ih������wo��l^W]�4+3���)?OH�������]"��X�5e.W�� �����h.�%�܏�:w~�w�k:��ΐ��5���EFs��l��IP�cS�ؿ�v�|���2ziBaW�[)tp�z��G��SR��o�w�\a�V���T�g:<~��3�[�d��04�B���"��oglFkhDD(\s�2��Bt:�HW�]n<�x����r�&pO	����W���7�y�Dx���f)b�Er�Tr�k���n�
8!�[v� T� ���)�6'�&�:�|�D�9ۜ{Dѝ��n=�s6���\����L�^�Am��~�i�}_9�@�[o.-V���眿8YX0q�7�6��t�$��%�˘UtF�v���N�l9˷�^z���<��#�&p�;w
��*�'V��Y�(�+�e�Pp�6ŵer]��nYneF����"���l�G�U~}��m/�!] �,�Js��v-YڽCx�C>}��븝xS�s��v+k����+n�)�H�s�Z]_���g��D=�(�	ҋ��)7΂�(�*��|D8nԛGX6=�{�Zo��ò�7^�ei/��_(s�o�P�<�O���9^��� t@E`���.��\�ٹx���nb���؆��� ���5��7�ə3�a�5���;ԧ�ٝ������Y��,?�X+e>{��=��u�
�. ?�v��]Zwm��.�+�� �{�iu��-�^�[#2����(�|'��Q����r< Ñ��E�/�;�^�����<�U�*7���r�m�˞6�t��v�U�M,��H�Y�5�=��}���V�Z7����8�`��8o�i�p��:WE�|'W��a�RP1T��OFq�)@�%�H�x�~�4��g��\6�z�3q`C����q��W|E�B�Rq���|:'����"�1���k�������L&��KO�7p[�{1"�ڴU�:;��+����m�Gz|�		��u]}�<W�c����@���-�c�q�s�5^4J�{�)C�w��=��0��2$��V���_b���)�c�r�	Ҙf��Ę����]�.[`jb�:���y{$��g���o�t����Ǯ�dD�>��;k�"#�Fç#�U��urz�����WM���5H�=*?]�g!3��E����ʮj�'�@o%�M�=S�aH����v��*�e��׷�����14�Y��'��F����0���Ь�U�?��Z����f��/��6=1ty'G�7���xׄηdOq�߁�P�u��a��=��ܱ3�ud�]��A�y�(�i��4��Ov�Ζ����Iv�У�yX��R�g;����#�z��Y$3$�R�݊Y���V��i
��F�aQ���Q^�%E]҉��{-�%��T�R�Q*��u�L���Fv�.^l�M���sqF��V�Wa�Е����[��2���u:�񞾻�]�<�{��$�}2cF��ń3G\g���Pb��	�t9\Q��޽/:�EMEizw��.���M�$�EÝ��n��9+U�ח�(otGL^G�r�A?���7�S�M���x�O4�GY��B�ܻ�P}�3�N;��^�K�Kqs�{F����W`ե�1�e0�e��)r��S(5nH�j?w<�هB���:�67��:�w�}����U{Ҥm3�0A�r���s�֒\���1W��y7�sP6-�;a�@�l�;�|�Nd(���°cY���Oo";0�\MD���v��"�U$_�q�[���)�%!E��V�7[�^c|Nft*�.{�XgL܊����f�!�=��Zȧ�Yzg�:v�ZOE���-��F��۳����cC�-�t��ۍ:������V�!ᱎy��w.6������B��+�z2��0��x����Q��YKz�jo;(�;�P���4�s1{N�@���h0�xć5�'E�ٚе28�yJ!����N�������r�/E�P;�ʱ !���H.�A�#8���;>�(#W��ܬ���4Kl�+�8�M�˽U��<�-N�������&F��u��E�5�����+�>c�cO/;km�Q��7��e�w��dm�������y��K�+1-���*K����V��szn�N*ጧ�7�gf��+�j#M=�HJ��Ү���D,l�_,�7>LY,IP����|�H���1W+��^8�bdV.ն׶�'��76!�B��W����1��ty���B�^VZ�s*�u,'�	yS�J���>9[��U�����9�� �{��Ʀ���V�w6Y���]xM��ޣ���'w{�s 3��́�5,)���5����Ptz� ��]Y�^Ou��*�Gs]��<r����ٻvi���n�[=�B�*��H���	O1��>Y���X�P��[�WzX[�+f����uV��9��������q�8ʛ6ƀ�����^&Ua��]���<�c��V)�`�~ɍӃω�ۖ/.h�U�A��+	�oH�Wr�D�����H��Ɔ���]>v�+�$�z7�(�y��6�b7�z�E1�7��q���+Zف���/�@f"E4N2��H�I}���j^5ҧ�����4<��z�B�-�Nz:Ķ�T.7�GR]�)�*���w������w�=u/mJ������(�3
/W;zj�T���;!�����z�a]�yG���2JHA΂Z>t��D�'
��:��~��f��q�)k\�p��A+�WA鰪���7]��*���Du�N�Ih��>��;��O��]､*��SpUѹດ	�ti�Z�#�4}D��Q-c�K�v�1$�:��"7��9t�rv9� |18z�Ix枯4�u7I�wޘ����Q슈ӜB&oX�"�1�Z�t�Bu�fl��G�Åf�!���Jk��'q��"h5#bMW�K���2q�Y�9t��*'*�J#�W��t��U�����o.� ���������:����H��
Ӹ@���s#D����� o^n�v��.Xӳ(.�,�3S�v�z��Au�l
wok�Y�X"\>���������N��	f�zY<nWcn� �{�H�u� `� p�bBg�m�
���	��D�V���yg=���P���9=,� �͵R��܂ex`��k�[v�鵐(�mZD���.�ө�<�������Y�Mzd��U����LK=����tG��I��]�B��N�fN��`Sꨲ���5s�Y&����&!>�9�p;��!}v6%��ZѦ�#�I����Q3�#_���� �0$�'f���m�r��7�%yX0�5a�G��wo���/�p��A�J]�VS�	�:��ٖ@���;=W:��ĭ7�M-Jh��*�׼���d@�e:$n��l�Zz ���<�>��-��~��g��}Qɞ�׻�K�D��z��6彾��g���]Z��F
�{t+hr�U���Wo�\�B���IO� IO�$ I(B��@�$���B��@�$����$��	!I�@IO�H@�p$�	'@�$�	!I�H@�`$�	'�H@�`$�	'�H@��$�	'��$ I=�$ I?�b��L���\dcn� � ���{λ �����<��AT
� :h(�*�T
 J�(7ە$u��ET�D��CP�kU@
EO6!(�$��UT�T	DPU
������J�9���5M%"�X����cMh��)\ \@'`5 �dY�ʬ�km�j���I*�D�� 1 �ɣk ���
Z	�5m�*j%-	��]hV���  ��  	 �J��УCU*��� 5Υ�r$�34�gN��eJ6��Wc
���5 ,
����7�q����U�,�R���M� Vm@�6F��UD���N��	R� Y�3���T�ͳm��V[dK(�H��f�vf&)���*�Jhf�i��%)@p&Glf�kDJif5&�����56�*0I"��L��6��	�*�kj��Y[Q�f�5ޢ�  S��T� 4     ��
R��bb`�dd0C#L@1�&0a0�` 2i�b)� �J'��0�4�L !�"�A124�O*~�i��i�ɚ�I����J	�&�d��i��dkկg\�uۮo��u�[a�]��@R�RNh*
�O�*5DED���!AR���������C��`Xt@1DB� ��H "��� U!�+ ��@u�ݶt��X�����f

�J�jKK?-R�g�L=s���IE/˷"��κ��_�0�V��a���m��L��%0MˣvV���X��[.��x/4���;z�6̰v�V#�-��wj*��l��m�IU�t~�nbݳ�Š�m
u>Zˣ2�ȩHJJ�X�,�EE7�W2��+ej��u��݋,�Ԭ����#�� �	�upՋYI�
�Ͷ���k7*�%�k�+�iO8mg��(�N�H�8��c��~{-HE�4�̊�b9�A��[(�C����w>$m)YW���p�u|E{s�!�X1��[���YF�51�nge]�����n�b��=�����]�P]�:B�gY��	֫E>6] ��IH�OT�W��-^��HF�c۸�ؕ���{A��J���t�4��*�n��;{���5��pL�@䩬M.�7Jb�֎�Y����#��%��پz�:�T��v�SM��n'�U��v4S;Y2�?�̨h��Y��R��Ӧ�IE��k�qe,j��j��!�g(=	��P��F�n��Q�g�kMҥw�,Q���\ύ��y���-%�#-X�m��+75��̽�

�i�oz���ü8F���m�@J	�co��hGf�Ɩ�$$̛w���1^	��c��Z!8]7��jΌ���$���>7y���am�4�MF���;̚U=T�O$�u���d�jwX���Km`�N�5t,�xu^����oi+`�e��4d�;��6�i�H}�_׏9SoU0�������MuywS=���]Bwn�l�^Ro(�+"��>؅t�
,��gU���5�Ž�.l]�U�G�Wh�h�U�g;�e:=z�ɰR5w�Цh�8*��&@�F�6��L�;dK��nl�����,*�`X�omm�t�݌4��q��;ɹ+c.�j��K]M-�A�a��Y2˛��luzJT���Ũ8h^=uܴ�3��řZ�C3v6)���&��,[�Ƕ�7c.��e?�ѩS��)�[*m����ݧ��[��l��7`#\\b�XtY��ݭ����ĻV(n����)Y�TbCx���^���2���2���{���V3VPm�Q�Y��1[��TJ��w8.����9��|eiHJ��%�����u�L:��)��2����X�śIm陂|X�t�^V,����u�B��[D�^�|�$3A%��3[�y��졕�n3V-;L����m�P�:u�gL[�`�(s5�G�N�M�,	���h��tM�<$�*{Q�8��0]Hw2��&���h)-�Xh�$�]�z��{��,�gq�B��j�}t��R�V�^'��]� oXV��v&R.��1�y�-�� ������wl����xZ�Q���6�`PЭ��6�i �h'�i���N��):��^�,>�yx4	�n���K��`��#����+/[޻!���V�k�����%�E�GVi��,d�ZA0Q�w������zpVjp�w)~����4Eb�x*ҭ�f�Ze<5��@��J�p�ڥ{K�Y�bm�e��Di<X��h^���u\�R�����k8]n-ԣ
R{rVYY�Q�Ɗ�x[Yor�j�8h6F}3u��B8�4^�e�',�k�cnLL��oX[�m��Y�t�Ȱ"P�/�M-V�f���1T9�B,�mA�c*奏q����Lfl��l0��3LZvx)�|�7�a4sU������;�� :\� ��w�v�,e�\<�p��@�(Y������p����fZtūn��&���MyiWt��B�ZL2��W�0��K���L�ZS����MdXR��јlj�
sv��)
�^�n2���{�����B�L���i�!�,�Z�����hj���n�3,�D+�h�w	%޺[�k�p�4��a|�<@���$�d��[Ǝ�w)��r���ޒ�B�܆^�g��c~�"��L�mLA[r�(b�J����`]@�v^�cfe��I�m�U�	�Z`�1}�\��Y��x�{D�oX�;$�ƒ�rR0;ȅ�ɢ\�ک[��[W6�K2*Z\�[q֠2��7[i5�zNEX�i�Hq��v�x�w��n�ձtֵ��*����/��l3z5���cr���D֌[��A�$�[���	0ۺ]���]��.�����״��J7[�g��'�/㮰��5oQ����W�k5��ȔB�u-���I]D��!�t^+yVu�mZ9l�נSc3bnI������C�Rʹ#�ֽ{�e-�l-ն$ʑ�`�3PEڊ�7]��B�̢��oj©*Œ�w;��Y��l���a�d�hm�i���V��6:�j"Tъ��V�Й�d�� %���^�M�u�
�Պ��ҥt�~�@Ⲍ���T�T�J����fݱ�%�����PJ��.���ĭ[�Fbtv�[�4H�|�{�2N����Y���ض��{QVl�.��w{n`a\гvIy���]k!�w�Hc40ZEe�4��7Q�ؖ2M�u��Ἡ[R�k6��4::��Ku�]��ڢ�2�3Nٲ��`�5P��ұ����`���ʫV�m+:n�r2���ߞ}�G��]�����#�O�~S����O�����[���ݹC2>Yg�J�<v��H���`}�:�*f���i��c��RG�&LWR�آ��[+>�S��gl�'�#]��˘�t�wH��S�wY��O�%>0�3�{rI��rl�ӭ>���c��①��n���t
i�Nv+�čŁ;�]�g ��Sᕰ��������ɻƲB�C��KL#&u�V��).��6��\���oQ���7�݀8��գ�� )������)ymñ9��Sd\9戥|�;�L�Ɠ<���_X�+t�M��H�~�n��(�r{�.�Ok.a�swnv��`�9�N^v���uxv�4�w��كu���WD��%�/b����Q{Tۖ{-ӫMoii��]p?���
��v��1t�o3^�.�� �u�-��夅�8K4s�m�.�Ķ�J�ֹ�Z�w
7ɈV�ac8&J��d��N�ɧ->�%�+���}�#,_P I�g͕w�>�S����lz�`�E�h�	�7��w��G=z�Y��4%�t]ݱ
U�*��P�`�%�,�Q��]N��RH,᷹Hȩ����6�V^���p̺�<�`���i=�e>��_�o��2���<�о�7�/s�}�U2dX�d��.��+j�_��{bc��ۥ2p�w����6�m�ξg�����h��2sۜKS}�C_G<ouWMߕH�
4�7���r|���K���i�#�����t[�C�r��˴3��� OC����ƚZv�Y�	�[+VF��o���������-�@�xrM�{����Ο�탔�yH�p\!������;G7�Ĭ�;��O��QE�uV���C2M9ĺ�`�4�,<��T�Y��8-M�|U�3�l���U�:�j��d� �/�%�8�e�n�Ұܝ�Ʀ$2;��;�X7S{fQ�
�Βpjל���K�Xȡ�!�m*c(C�9�#|�\v�ѻ�+-��{GiWЫ(�����	�c����`�};;���R;wD�D�Ȭ=ؚ#&Hr�]68�!�ŗ�1޶&���q����Sh>}�^�����:p�6�;`aK.�Y�p��B�ű!v����{s�g�-��l�oc�ou�*������Yz��w���Q��V�C՛�u@�����,�B�^Vw=��ii�U��7��4��ԛ��eY��2����nݥs5k"c��h�ut�:9�����v(���͒��5@����ɺ�l[�x����I���?qO �mVL�(�e��LJEN�H��wN"���$�B�I]�E��sgoe�=� X*d{B�W����M�,��{��K�ge�>⎥�6����kR.�X�0�g٪�)g8Uu��������gfIi�����D�����uc�]�TkA�ǯi�#����� ��4vg�{w��u��C����Z3@�|�fv�T���kc㥑� `�l�9[��E���m�NĒ��/��;�Y��ծ��,!%����(��7�)���y����\it�'7q�}�䬊�����5	qk.b(��z�ӆ�%�]��tvsj]-��Y�ԓ�.�/�c:<��p���yd<㣐|�r�t�Ct���wYf�a�Fs}rX.�WJ����ń@!N�-maqC(c�T����z��Wo)�}�G&�\�-�Ȧ�l_N{�jS���ɤ��v��Z�u\'㪐�;4@^�6��Y[Qnu�A7(]꣩�;P�m�
�{I����O2V�ղ",�[�ܟd���9|��yg6��|:�KPvs�崫L��TTlf��VN|�k����Ip�뻊`�wq���ʓ�	��
���_k���@Ԡ��S7Kvc@<���9l�s��X �l�{}�{������ �;���M�ejS���z��l��÷+���|���v���u���;\yk`Ū��n
���h���mč_1^�M��+�Foh�ݘ:�7Nn��eʹ�s77	�4�V������+�r�3(F��t��y�ᑜ|�Rr����Χ��M��v�Q��z�#w���Gp�o{��:�a�yy�x���kx��H�P�̑�$��ܒ96 �r3��HJ7"�rG�%$��RXS��gP2Ԋ����2L�܎�qz�n\���t�q���s����4Ĺ��o�NnĊ�sf�^���7��m��Q��!'�c�[��8���)�'wQi�i���ԡ4Fpn��n�<q�x���G}M������Ʈ�0�w��$�z�m_�BR�:�"�R���f&�5���]*]r�8n���-�V��JqX��@�R��v���p���	�uԽ��9��Ok�d�l���XM�|jV��4 4�������z�v�R�NȤ�b��!�fG�4^v��򖫨�@&+Olo�ysa�z�r����mֳ�i���p����:��ɬ��.l�֧
���V���m�v:��a�.h��r��]�X�}�����o���� �`=�/��XS��lӻ%!��Ӄ6�����l��0a7Wh:���q���jof^�> �tp}$s�ܗ�1��|ᶽ��c� �)�ڸ2�u��Y]Nྭ����~��_��q�эt�c?@QAS^��E���*�ݍC�p;�PPT�:�i�c��]v�u�w[O��^o����lB�q�GMk�]ɸ�)�$�6�5��H�X\]��y�;E��VW"�WQ+{֍wN�i�mH�A�R�D;�s���z���V�r*��䤜��T�vUNysb���T�B9v���5���\�]L �e0I�Z�N��k��ݮµɯ;(.����}+u_�v�ۡ�TA�ѐ1\�P��a�+
�h:J�Q3��p���Rr�)��Ҟ�#�Y{o.�[���$p�+�jQŢ䎚���O>��FҶ��>'hsE�е�(u?������ -�bb$�q�SϺ�v'Fn�s+��
����b���|t����W��B��%��X:��I����yu2�%��Xof��e5B���Y��ӷw2�mf��n�/r�Ĝ���m�C�O�:ћՋ�#ثB�֎��Z�J9�1녹Ş.id�n�wL�o��|,���̍m��;;������vx����'D�l��ɪko)����\)�]n�C�{��/�5�9]�#3����7��Yֶ1N�ovM����2��=ݔ��6y��6���n)�㻂�u7%���wV�Mv:�2����J�A���߷4�Z��vW!n��]H8Ҿ��,�x����.�E����E�u�p:���Ֆ@�$͖���.4�ח�kd�*�s�:��^�{�{�5��q�LR��Y:�2�$A���r��]���� 6Ck%�ї1�<�O���oN՜Т�vՌE^PV���(ɝ%M�X"�$b%�HW:�0��и�&I%֜T�Ӽ��Ʌm�w!��㣊�;1����Q�m��k�q���%�W�xtyҺ\���JikeZz݃�.;p��@JdF/���H��z����9%�����B�o$��'�sA�"<kGP}�$U:vB,����U����T7)�����ܗ�1Rڭtj�����a������㹷96ںMU���vS�W�n�Z |.��d�Z�-�R/�j��|&K�A`�17�u��%%��t	�e�.��2��J��i�%7\�RF�]`/���"gX����GEG�ŐVe^�"I�Q�d]c��gY$Л݁ˬյg{���Yx��[Yu���Q�e1�ؙ��u-,d�tb7�V���m�.� h�r���Z��[m��R�ێS_:��ܖŗ{<��&���*48+���h޶L��<�ۢ�9��7E]�q�ӹ[���a�"Dn��}O��z�� �ܤ�[�� �YR�#��2B��6�Y�U���go�(�_p���q�R��
���0�5�69�j:�˾Ðb���um�]��l5|r�°�@�n����1��7��}jub�3f'B�g0��&����*�)�9�c�ĭ��U�;��%`�TP�֦	'u�<�d,�Lͤ��T�������j�6��x0�4��,��a;t-�u(p���6�jﵮZ�ZB����f�M��O0���yP�7�*vj9�[;�8����^�F>5(ʽR�[�kf��|��z&�*�1�U�JB��;�P�98�8o�pʒXӃ�;q�!τE�Y�5�ޭ:2������ڤ1���2b1�V,���o8v��-�C���p .�+���ހ�aa{0c���z�ud��W�0B¶��wK.�c%��z�:�n}�n����[�Z�T�p:��v��Ɓ��h�^�h�� Uh釃�at6�Q�u*&;�#)�f��e.�Vi	�ѫJ8,Sf��#sy��k�1�)]t"+�kp�����4�#!yƆ�Ps�e9�f����n�e��h���5���U��!e��v�^Ϭ�y�Cy$�}�;�!�!�V�6��8�fwWu<��Cg5���<�ugە���]uX��� `�b�Ǖn�<�`�Q�˳�:w�EuCW��;"��8:�ި�"-1 x���8Ǝ4���}���fO�Z�wR�Yn]�4UsUy@cfk<f��%�a�AZP�j�����ә��TllMD8��]&��Jcct���/9a�sG�hj����d�6C��˖�֥I���+m&ݐ�Y`�R�:���=�iT���F��յ�	����[<i��#���ہu�@��'Z�"���9`�l��`%`���i��C�n�Z�HGo���V��޴�ݻ�vBo�0maW�1�Kf67�1�>J�����W���a�y�wA5F]��F�T�M��T꺅 x�����Z��E�B5�x�e``�k���{g�fW-�쳁:pB��b!�A�&�]`��-�w��:�c7S^��������iv^�էX�i��];:��߮�)�N����k�Q�I�={J��nLE�S�d��t�fgJ�ѧA�G�%幆��Vr�Z�]�G��(ی����rbA�-�e�؉fD���+%H���@᧳��Q��+�H%B�A'(�rP���e�q[�vk(�]���T=����i���hB�VJۓ!�\����.Jt��-q�
V�`冘�uc��n��d����DI1:�u��7�؍'^n(6��^��Cw�o:���܄�\e��sa��sUp�'� �$��_���2A�a�茈�s�w����s9߼�{�šD�nݨV���L^��Tf���ֱ���L{j�);E��*j+0� �V4)�c莊N��}l+��ZwmY̬��%ܾϰX�k��.�n��i}{��bjbU!��![Yr��	�N�`�5t�īa�E�������q}�i��,T�^�5���d	In�x'Cx�.�`�b�tha����Z���ű�=�Eh��'.ۋ�p��6Jc٣;��%$����1u�^.;�f���X]>�ͬD��-�o5���Vuѱ�*�B���J���̢֕�ԫ��e�up1�FƶK�ȳWm���LB�*�K1�e�9��
+t�c��miP���X�R�QX��h���l�T��lr�JkU���m��f-�کDlQ2�ZQ�Lpq�(����6����s}��{鶊Ɩ��bd���!��#�TN�ߴ?w�|d&�b7��b�X��Uݵ4t=�yR�*=�=��Ii�N����xߋY]^�����ޕ1Y���OOTy�������,a�����x�<��f�%��m�.�'-\�fq�!ѭ�۸�ܫ�X�j+����&U��	*���,.�^�n��C���W?�xtV�_��:".�薮�a��e�״@�ݙ�#�7̜QF2#�9F?�^^��S�/��R��.�NЇ/1XM���'�Ѻ�5�6����B��4M�0���aj�f٬y`�&�_]\�Mb���O6]N%W^��BBd�>޶�`ѦI�ӗM��ţ��$��Z��g�����{�h�w4:�[��\=Vݽ&E��/^�[i�ہM_n�Sղ�Y*U�.�����X�L9�k ݻ�5���6B�z*�"�^�ò�S=o9��˙2^�x�-Ԑ��-t23�(�n�.[�;i��to�xYsv�ޡOz������Q൑���9��qsO}����0�����5}�Q���'���&j��`��{���w�ɆDX.�)VO<3�9=iJv����QiE$�+7��E�	����S}מ�O�a$2��h�Η�z ��.h;c:m�V^�)���Y���.�ۮ�x�'hUj��B���]%b����J`ś�)�ș2IǏI�E�F�E��s�u	�����h���T�N��.�_��^�#�����P`4_-1uz�Ѯ~@[�/��x�F��p�%ﰁj�uw<|"����8K�X�U��e 7쀮�_J��3Xԩ2��j��m�Z���.���u�I1��A5�3��Ӹ���������p�GsHjqӶ�E2���<&ɻX��KJ�Ax���-̋ymԮs$ek�B�#=�K��r�~�tZ̩L�U5�{G��^�'Ug�ks��=���L�l%\�.:f�/.S?EP��/��Z���U�ci�T�<r9�a�c&�.���'K��.)gZ�a�w76rg�ب��]�ۉ���x�g���U�@�),������ ��?WY��/%�5[�y�Dh-p�2v��<a�CQ�P�U#[1�jћ���'ˉ�:�9�NeE1��mIA#���;����*��4x�\�U*�C[@�I���Z���}����yzi���𭺦�d'�S�K�]ln꾋��&�����2w����e��-w������o�����r`�	��{4.�:���
U�C/�<�츆��Y��۴nL��w����<E�ٸ72tě��9[���exc�l�0�$r@J�wmjOS�(�NK��6��ws��e8Ƴ�Y�5�$�r�5/4�ƙuz�lE���˷��*�@�:<+G�޾Q�ؾn�:s�yb���|M�S�6����%�[q��^;]��jx��oگ��u]r��8�`�J��2`�L��/8�1�n)�o��4���uwV��S��wf=V߱+�n�DU��jNޮv�=^�t�GCu�/��\ NU�t��L���y&eV��<��>1�j_�����1)��{d1N7U�Y����b����dw��M�i1 �dŅ,����_^��+��t�9���it��כt�o�ݤD��BoGXVd��Ez��h�m����z**'9k�����K�P^Zq�9�K��3�߮J֚|<����O
^T��y\=���y{xP�j)���;�\�%�[�]6f��Hu"4�;|Uݭ�F��MT�A���9�(�ԋ�q�I珰�B哻/G��������
��do�Լ~��6!vtC��
�K<��K�d�˴��<T���l"z���+pg�
?~"�l�b���r� �vn!?l����Ǚek0Y�f�~�D%Y�;:���o��IkA��Gn��b�}��lJRi�=�줹�'sb�t�����K�x�ZowR3��N�����H\�A��ܷ�ΣP0�Nn�%�H����#��/��S�F/$�ya�&Y���s��Vm�����^�P=P{��t��OOR��R��)���B��Ɵ#ü�!��'{����W��@�
Afg�ä��%L����s��g��+�>+#�U��C�X	�-y�1}�n�Z��e�V�E�����>�{��o���vW|����z��/�of��n(�ڂ�W��gqĔ���[k���t�f�kU9n�������oKԾg��W_e��ȫ�*9Z��d�/oUr���1`��.����C�F�pY.Z��fQS%����E乚��Y�&����ZB�Y�׻f	
:)�K1�����l���j���vya��!w�m�,�X8F���yA�h]۫��]:#v�M������X�/�}��<����g~b��K�Sg�MŲ���)n��j0�L�����թl�R��ٔ�u嘕�1��>�?}�NF��tT����Fm�/�>9��K6��@��n��.a8ӽ��R��˽��>5GB���;B/�|�4.j��Ѕݾy�JA�
���xT��z��ڡ���������#�-zera� �%*�d�t���oG��n�G�T�cI�ҭ����2�ӛ7;j.<h_sڅ_Y=��$���.�j��e���#�z8����Rp�R���m�2�mZ��ޱ/��;V�%g&�c i�v��oa1�t����;�75؊��aU���V,:h�l��(\J�2�3��2�e̘�J�cKQJ�Rܲ�Ԫ��R�j*�+#h�SX��e�"%�(V�[�j�(��m�ژ���+iFQ�ŶȌ��U%)G)Z��E*���[l��J�T�H�,����.aq��11���qңUm��X2Ҡ��,MC�޹��
Uߧ��ۚFD(��Aͩ ��ʭ��`�Ŷ�w�n�CW�ԭ��M���;��;"��E����Ǿ?,룈�q���>�(|G�_cL��~b�����4c�T��̬�����h���O��K8s�U�(�uu���jf��x�ǯ����
��.�`{ls턬�G���'؃���G��se�ߧ�O%�m�.�������	��:��K�ׂ���cեR�9dG����bV�z�n�3�wX���S���jg%~|��{��@h�(�O+����w��*�)�fj[��c�4��]]�[�ާ�+�'���/b�Iݒ���3��TG4�F)�]��֏v���֓E�O�:g���e���x�r��De��|+�TIz��V.��b���J�Y���h*юW!��WB�Guvx�k���348ԹwE�gS���s~̯x��3@)(�y�a=�d25�&�/�oJ��������<9â���}xπ�uռx�']t�rc�t����]�^��m��������\T�4G2���I���3���\.��K��ȶ�����t��wX�z�5�A�<Hm�d��C�b�#�N�j!�_2Z�IQ��B�TkP�	�!�X��5�G[�}���t�:λ��( i�{[3]���꼾�X�~��e�9� �.7%�Ӊ���r��ñ��L���uB�}o�)��g��9.X*u<�y�s�Lu�P kt��=��|M���1&R�:C�N͍�n�ݐ���jW�I��8���Vw��q��f�t�'�mf'i`��\�<�N��E�QbzU��7��4z_��M�M����Y,����,v�Mt��s�p��g���o&TIͭ����6�U��3=o�Q��Q$%r��B;�ځ�r�i8[��v;��{�qZ��/���G�(�a��"Hg�igwӗy^�w�v�$U����zص���3����<�*�Ɋ���:p��k�n�S�8��pfT6��X�������3��?}4N�D��M�7�v�r�~���)I�E?.������c�c�y��^y��~�U��9g��$�i�W����Q�t3�h���
�]/Z�ze߬��PQ�Y��R�H������[��oP�ռ����2j��x�L��~|�gڳ�0\uHxu*�T�H�7�0u_I��ND�nr̭�/d��SB+�,���Z�X�@�)�@=��K��S;�Fp��<*�>&�j�x�ל]HJla�ٺ4�8�nUQJ����u�u-n_c7�����8'3��S��Uc�cf�H1�w:6���t/j�(Z�ʇ��ұ����Hԋ�5sG1+�0�j~Lfx�����E���T>u���Y{�I7įL��-�4ז'�i��K��D�UW�Q�y�; ����(l�|0\'�X��,�Nߪ�x��S�E��C�}��>Z���F_+�±�}��6�ĚW	+��M�E�<��V�]ݫ=7�K���VR��t;���N�
<���*8��b�Z����6�Z�E��&�3v�2��M9pF[��V��6��ǈ`s��P�{���F�*Vz��}�We�J6���8ˏ�}E3�	��8(�n9�2��J9����飶��[�0n�oN3��+���V����_P��]����ߦ�"Q"C��KA�w�<Es{x2Aݛ���Ҵhz*8��f�l1v�>ęt���U�H�[�y����x�e�J���}�^�m�����}��n	I���"��s��[�*;&)o99M�yJ�獽������w����}�����r]x���*�	������J�Q�%f��-�x���HC#�p�]�����)���n�s�g���v�����o���u���v�¨����mOE��1c���}+;��gQ����;8VW8��wqKT�^��f���0F�Z��˲&�R[l���%��P9�{i�*��F���W(�f�-�_I$g;d�%�+�~2C�~��+"�P����Y�圭�.��[�^�6d�^t�?ɣ�Z�hy{�^����'m�9��N9��U��v2.���w��)�I�ٌ�ն[������#9F�z�Le�ѵяn}W�U
Bq����j�9�k�]3�<юؠ��ŕ�>y�TI���|������M��i�nhI,�6�_��cz���������m�V��Ÿi� ��6n���h�̍C�M���靨�E]s`�Qt]b�\Cty-�mwp+��k
�Х�Wte_=�Y�8u�K�V�Z�Xx^�����l�L^�v��/�ڵ�ڲt��L���s�S�w�!Xhd��U{,b������MT[/ ��Y��0�l�wd
���uhC*��Z���'0M4:'"I�YZ�F�J��ʷ��L�P��dX]4ˆ1��yC�(o�H�cr��\	�45�`���|�J��C��_��~���k�����hW�;ll+n�b���B�NYw�1s�N�W�|�;q)$��#�����+Q�F���A8�*��L�4��Uˌ�(��Xef:T�����n��h��G�9���4�1Q�M����e.��b�-�<�#��
�ѽR��֩�}(mIDLv�j7;.P���ٗ!�
+m及���L��6�#R��J��'"Ifk��Ҷ@"�L���̫冺��E��t�8	]���]���"6e(��_����!�c*�Z��V�ce�ز��S
ZT*Z��ʊT1�m[F�c�-[h�,X(�U��)h�V����h�F���X(TR�b�օQ.P�Q1�j�j�mK�E&5�TbŅE"�؎aW�6�ʬ�P�T�@U�V�,D�ȪEUZ�j�9�
JȱdPiZ�,*-j"[Kl*T*��-�b0Z���)ڢŨ,�%V"��e&1H��
��̮E
Z[,Z�R���ң��sW�z��k�͝=_��2��U9��.3�&���,��hw<�;�����=D.7x|�?���HI��FĤ"�5��3G;���P�ҁ��/(�o�߽�F�$�$(y��{��8��ܬ�G���7Yb�`2⥾˭�NŇ/ہ�U��䮠f�Wֶ<��4�o�&E�̎��4����}��JayҦ������]�6�"�
?�/R;��nn���Nz%�+�5��D2���e�������'>=��g��>wN�����hx�i!i��� �T��8vx=��hxgQ��}ڛ��k�+�:r�~m�R�v����c����$[]�V�O�س�%�;�s�"��VZ\�9ƻ{��m�a�i�ןy�Oq��潥f�lg������s=�]�\���W:�U�1L���]�i�j/5S)�ȃ�k�Fgc�>=����w�8�/LsoeK��$E=��kY1�d���_!37��A8oV"�z��\s$���OR��C}%V��Ugb������F�+�[��C�Ć�� ���e�ז��@o�L]�z[]�י��y���K�\EP\C�5(o�s�ûbut�TЀ믖�;j����]�1r��;j�.ٍ�s��ܻ#�cQ]k]�;Ã�b\С�}�G��Ӥ4����sЙ�;M�ywV�@7;�9��ʍ�d9�̐]3WK|�n�U���[Q��1��˚��Gk�uF��T�=D��嘞i�;e�Q��t�-ϳ�@��Ҝ���Os�H2���>�J^�g�כt�@X���o�������{y��w��t�U��z�S K�^�=���r��"2���DQ�S�>�`gc�����ͦ��x�i3�ǽ;���������M�-I
����fe�$�)�5��g�@2V-�+���m
�~��e�B�q�.����&���Tm%���K�{2 0 n�y�YPo-��w�D��<��M�v����z�)�;���6Cͷ tuC�-4�s�YSV�b���v�+�kQ=����y:�/�7���͟=ܮ`�B�MO*~m�Ew�f��:���[կ�6�:x"z����p��>��������)����i����r�
FtĤ����y{�z?�{_�~5��-���I!�T+�,��7������橇�Ě�w�/?Y�WH(�a�K�%�Yq:2/%�B��^~��6:�Ys�.��lF$^��g�c^��8,����W�'�(�q8�mm�Ym{��>6��d I�b+Ժ��8�&�iG���}�r�,5��%t�,ݩ�nR;�Ǐj)^k�%
�%0�Ӂ��:!pM�҅�%�?}�Q���n������y����We�%v���3�לU3K�C"�������>���p���4^� ����q�X��-9�:���G�uF��y�%-��_;�|#ue�wx_����k�P���9>����L^e����S�2t��O\ǹT����:���oޫ��Z��]��tA��h��4�,ߕ�vA����3ibi�7�z�CWa���V��(J2;�9ڧMTq���%�s�}U��}��~��������s�
�C�n�*�C}����~������o�o	�I�݇{��^D����tC=�	���Ώ= ��)Y����+���Ļ�<��̨����`��"���/ы�7U�r9n��|�&1X�����L�X���mS��F��vA�7V�1�M���� ���@Jϱ���^�>���h���r�!�窢�����ڎc�5'��M�/�����ʊ�GK�>qC���r����p��1�����7�wr�OJ}���6�t��K|���3�4��JmKjm�|�`��]n�n�k̓B��`�4�^'h��n\�y��9k�{Aַ0���z̹�����oN�\��J��h��1��k�zC��6e_�t��X�[��@k�3��G�©���y��n�A�N��p2�qS���_��O��UUV����;��'�V��h`��9�SLVX��3&3q툛���P���o�b.�v��.ޝA��|s�l�<s.ƽ����o�̊�` �u��һ����q(3�t�wq���w�zב~t���Nz����mm�W�"�$��DV(r����u��I�\��'hX,� /��:c�Kk���M >h~/������\��3�w9y�u	B��p� [�z��26\'~��M�Ԯ�+f��	Ȏ��PVm�5�+Ǜ뜑ެ�=�/�Y���*����.�vV�QG���I]��9�F������D�^�e�K@47b��=����"��e�֩�E�Ӻ=�W���Z���i%r��5j��k]h�껝]HmN
Xߴ�{Z��#��X],Q�F�&Ώ��/��
_pi�J���6��Ji�CU�0�a�\���1��7Kyb��#��ӱ���N��	�M���>9�tf�Ż��J���a�9wS�f�V�L��{7�<:S�3K#u9ȫ��9ǹjL6,jܽ�dW;b�(Nv��ofR�J�������[!�?��{/�C6�aU�ݡ^�ZV<��Ԭ��o;�]K-��.�M먴�"K�2�S���X)��t�6��l�E��Æ�qӐӈ�Uίm.��LP��ꖒ�")I�#�r������M�VJ�]����U��
Z��I�N���q��aռ�=y���jRE�_��� *]%�T1��R�R���Z�r�1�EX�J�J����A��[V�˔Z�+�%(�(e�Ld��L�\Ȋ�[[U�2�j�R��2���������UT����2�\���(V�1�lj��[�W��@��Y-�J¸�\*�F�iX�+(�*�1JU����fXcRR�leJ�����-����*���җ�ڭH9B��Y33 ��wYU��4~��7�~�����LT!��l25�'����9z���z#�ÖL�В�p��|�`�V�v9z���ҷȎ ���W+v���%4��0/
�q����{�"1W��'%��W�|��Է�w
g����9��t�M6;� ̫�5��.�~'+�`�_�L�B:K���6�[0��I����W�:aj�F䥷����gs�԰.��윺E�f;�e#+�
����K�Ү5�3p�Ë��*'�#s�UW�}]�p�@���Q_�_�$�Ũ�}3���7@��;}b��>�`t��C;c$�]���=..{&!�oLE�H6���R��s��6{n���%Y<�y����'͛=sM�� �Z��Y��j�2��l�+.��(U_:7��u�4�N��a�r�ӑ�����d�T�v��_,Y-��唤��Ӣ֦�`��v��6�o"��Suc����+�9n<X��E�#�U_}����X��jË_V�
�7�.w���M�WB����'N-Ѻ,��]P�Q��Ϣ{�xΐ��*�Q�Ľ�@tm�J�m�x��w����V�o[QR�H�_>ך��ޭ�p��ۥ�5�|=bG%]5Ƹ>���.s�;�p�n��.Z���tw�J�S�y�3�׌^�~�9s��o���eQ�2��戉���f�k蘤�f�ͦg#�M?�LO&�*990���B�g�yzO���}_}�1���翎>��;�����K���j"3V������ϖ/w�����l:��/�h^q�s����oD��ïZ
�^����9Ӿ�y� ={H�b�}�U=�Ԯݨ��,�����s���7w�g9ݎx+�.��l��]�J&t7�U��r����^!v�W8 ��s}�����e�C��lt��i�:1-�V�]J3���\��8��Qq'�� Y�w��=B�I
�n���a�	�O�x�XO'�m0�ěd�@�uμ��������+�8�q��I�'PIٻ'�r��`z�N�N�%I�6����߽����Y&0�$�@>d��C[�����$�Cl'���q��O/��:�ܛd��Hb'�HtȤ��6ɶHk�2`2q ��Hxæ�����~o��CϬ�3vC���&���
�0�{@��Ԝs�I�{��Fn��w�I�Bs�$)�i&u|I��aI�v��,%`|�Q��L�wּ��o�u���T4�6��!�<I�����a�iL���'z����I�'�K�&��!�l&Ӷ@Sz����6�>BtȲM�c���3޹�C��a��6��O�!���x�Vl�i6�2m �H�����]=�hd=Ha]�Oc;B���2�:�� xB^���xxi��}� ��Y�7M������&'���N��k)����(M)�c��q�ͨ�!q��9�� Hfu�}��<@R�����$�
�:H"@�����l�{����<�HT!�q�Hr�������d���$�C�;d�}ߞ��.vs�C�I���OY�XM�q5�Hz�l<a:<���a���d���>�>����O���X0�d� �E�P��x�<Aa����t�$�;��~����IX�'�S���H^��q@�I�����8���$�{��<�3]n�!R�2M0�'�Y!����q �`|��z�<g�o�;�9� �0��	;dVt��t�_\d��ju̒�x�ć{y��׎�4��!�Y��m$@P'I>`iq$��Rt�
}��9�.����c$�9�'&r�|��m�r�1l�0��;d
�$�l��)=�뮵��ll���m��<�!��z������@�l��Hk�!��I�!'��^����G��l]�6��i�x�b��D�5$��V��A��g+/x'+V�I�TvR�s�y���k�{�Hx�~2q�Ĝtr��r@����I���I� i��t�{�~��L�$�'�I6�h�2\�;Ha���Y!r��$8���q=����V�}��0Hz��q'�������qf}d�2�;a�Ra=3������+8���,8�3�>d���6��t�N!XD��Y ���=��g�C�I4��[�'�=g�!�8Ȳ�d:B`��I;d��������g�}��HC�d=Bq��N�>I�ya�ya��i��$!;a�	�;I6��:��y���0D 0xz��������.��7on���<�\�4\���=���F�}s�r���,ʂc�h�R�X��p�m�W	��k޲��&�l�K�*[wp�ۡw9��f_�ڰQ<1=.[������W��U-���M_��u�h7V?w�ܬ�es�cz�O�m�Tv��t�ćj�G�q� �����Яg�D'��VN>&v�:U}�v�5u��N��K���zΩ��7�.�\��ٹ~�����j�8)L��36�.�U�mV����|.wW�.���_9�R��ە^h��TYQ�:��b����L��V�N�wy�n��?X�{3���(uN�,sT�����Ҍ�9������^���]�ﶧ�=ج�����-��P��ܼyb�E�}�J�e���M��'������p�=���)&��Iz��p����+(���m�m+�G�C{4�^���-G=�m�2D܆gs���{�<l���|�'�����҉cI���yR�k7B,��<}���Fc�-TT	Ʃq�+_eZtf*,ôts2��YǅTѨ�3���ﾪ���"{��z?=L�qn�|��Xj1���$V�����0���p��	}@�����x�} ܑR�]���&z���ط*`�봙��J�6����Ո�D�+=b�*�U��7����hAخ�I����Uk�Ϻ{��+��~��r�kA�3�����յb��h�q �}�����߱e̳ ��'���a\�Po�F��9�����s��a 	��;ɇ�4n^�t�s'l40�6�Dl��q�H��tt����i�+xgn�fS��dG�E �N$��BK�GN�+�p�u��F���%)�f���6�Z���}����\( #��[N��K9�I�\]����Vu�#r�e*=eF�
��eNIwp|~���L\���h�rf��L
ä �2��J�G���_X�����М�u�O�,�pW�jm��kXT��x[�:�����Sj�=e��o&0.iA*c}w�j�Y�'���CU����21����-�c��v�f��]�{�e��u�z� ۢ>*a��:\�2�R��N@%��gr�rt��hu�䘵��Ⱦ�.�R�+
���K��f1;�6J.��{�n\;y6���WW]Q:x��
#yo"�[��Ŕ5c�ԫԏ	��Q���Re����֥Y��2F^���PL�)M�c��ۃ�����q)����r�re��[����]�B{K,�[�}�*u�f�==��D
l|z��TG�|(||��fF���FE�����)B�V�Z���kP��(�j)YV�*̶9f[r��aYYm"2cp�5��\��(`��2+.eB����%q0���(�+ZV��\2��+U�a�R9ldV*�-�&$*."��33eɖ䢉R�����R�%-ZW+h��s&Aq��ҲcU0\���aTr�$XVB�eLeq�9aRS�9l��E'��J[��38�2l�r�qaq,O�%����H�[��>�i���)��4�U��q;�f�mkB�;�'G���dH���w���j�FU��FZ�����b�� рٰ�\yꃴ�#��I�tr�Fѝ��u�h`�=z��X�*��[@�6�$g�-��
�g�MA�-ׅ4g`��6p�Y|>:l��%�\��ўm�I��=�sFsxa��uLM�g��^������3\MV�X3Ơ���Ц*#�\1oq� ������~ZD��i|.�
�X��S�+�%��rÙ*�?o�����fN����I7�� ���9��ɵ1d9�⓿�UP�k_1����E*8p���	�;�"�s����ő1<Hf�r���x�'Qhib��OY6ytzJ��"��J/P�`�c��V97��p��P,���b�Lp|k�+�hŵd��ٯq`��-e ,�}MI���s�v�3����Y���-2}�V|����yS�Sc^�T�����,�Rp����q/���'������:��U~?m�p���<��xca� ����\;*����9�hbB�R��l�i�fLcjLE�36��f��޳V�$&�&�����̠P婰�' S`y��]���q�f9ꪯ����NU/�Y-]%Q���C�"�f���6F��ńY�£sфCX�{[,�C�A�B�h�(:l݇S�K�f�,Kb����#�]*l�H�01��$�\;'�d�fO�D2�.,ڇ��{t�b"]����bA4C"<95�I��VBg�h�>�k �(;6m@7�U� L��q��UX*��j������d|ap�_��;5�~u펝
G�qot!g��%���Y1YY�K�k�b#�V�q�<�?,w�4��yd�l���v�;�AWr]M2ޖۨď.Z`��裟���fm�#�DE?T���*~�էǣ~��
�gd�!�ҡQ��z�4Y���u�i����3�h�C��+VBhY<Y���EE��D�E�G3h1�]!H�D�ԪF�F�uh�d�A
qE�>��BϨ�\Y�V\�1�����Iմ�f%yr��0��hV��vN��L�o/I�g�v}̵��Mm5u��f�����*E|>𰥪ڋ��o���W� !V�����$��u�H���ŝ(��6}����3!�f�y�k޹�7��}ޢ�i�er�*�i.���][;yvhS�-�.�8DpJ2#}�)�ș�9�����v���)!@�|���é	�g!<��g��׿XU�f�A.�;��w!��~5�xpj��e�r�Y�@U���F�#˲	���M�=O��~�x����Ҕ��F�ִ煩�}f���e�^&'l���wl�3��m�tu��V���':FL�}mQ���{v���ooxV,;�@Ԭ�!5�ik��s�k<�0��4��tI�Bό�y�E���]X�G��/$t���4���I�r�.�^�P1L�F�aB�5a4���_�
��]}�{�%�]\�[�|��xϡ�V�'���E��¸�Ӯs$in��B�2��}�}�Á�����8d�(��^�i�Gؕ������,T{��^�R��b�A��5��=�:�4r�"j�y`ǫ�\����fouz�E�FZ㐆GD��HL**�{.5�5HP�b����<x�ZA>�����������5yy>dV���#p�2���{VY0Y�U/��0Gi��l�'��
� �:D5�>h�E'�4UWK�����3dg /<�PCK�
���d.#OLů+\t��adi�� �?�U���.���t�ZV}�KSai5�N��4��Q�T�-��p��Z�U�0���"�ԌC��ԟϾ����~�������R���n*��Oi��Y�lCo&����o�y�;��wN��F���+��$�DY��$�Ӏ��ȫC!��;����?e�����7AV�p٢z�K��Cf`Q�e�f�m�>�D�!�^f�V����hYBfȳ��_,���Q:���Yr��ĺ�����T�/�g��н�Ⱥ��˘&lTk��>�X�xA���B��M��m�����i$#.7}J���U��핧�r�!�v�|�AN.�YH�����QT���N�c�\��N1��ow���Ֆ�?0�� ��CO�AW���4g�cn�a��C$�:u����aamr��س����5�-�:j�p��-_lu�	����}���Ƽ8V]��f�Z�ƴ0������4 �����!_*x�>[���2�Z��U��6
4E@�O��>�U���j�6l��VF�Pc�d+"�
���o�jW�B�X�Pyxh�0׈�Vd��j��^]ڂl�ņ ���
��
�����.�
��t��&¦~>6*�IU�pO�8A�΀]�!rț�����y�t��t�.�����&4��f�������1)?}U�(�l�r�a3'ѝ� ���<��Q$a;�oφU��8S�Y��!�.#C�&�W/H=��M?<u�V��: A�c�iFϸFI���i>s�x�!����M���c�Tv����`EDH��oP�E�:^v�w5 dDز7��̍�ǌ]��k{	Ub��
�a��9�⽌<�r�W�sf�F���daG�R��8�����Y�l�8��i&Z�,��e&�\e^������t�L�l�YWh�����Z3����v�w�j!]�'f���J��E�̛���:T��H��-�r-��mȹ���U��|2��Ϩ�k����TF�B }@\�9�u�V �r��,���{����"ס-Y\���^�B,�g�z}da�HY�u��.m�6��
!c�2D��y��T@�Yq�U��6x>p	�nN"���Κ�Gؔf*��tƌ����3'$F��؉d�T�L]�A6t�#��@H���5{��:d��܉|�Iuׁz�}��A��Yk�krC-��P�p<��b�-j����>�������;6�+�y򓖬���E�7��GG��t�7�|eȡ<B�X]Q���۵k�7tS2$wo��r$n:9Xx<�R���Mw�>o/K��!ã�gQ�{g*�lawX,թ�"��4R�3)�uv���8�ڱb��K�C��e9ƺb�e���z'�7/;��$f����㵱�b�̕��P�v��@��xj����Ӕ��e&�v�,�;ui��#	����CW�*�<��\�`� ��{IT����;���U��S�yZ;���E+����d��6�U��kL�5v�טa1�iCWv�����U3n��Eծ#�mv[f��2�Ze5�����V�.��O-�/��uVs1�ႛ!.�`�]+=;��J�t�ImvoXY��z���= ����\T�k뉼�Vf�-!��1�R���h�� WP��E���&|3���=\���.z�-�������̑�d��X�=�G*Y����Iڀ��svu��U4sDu��N҃�ڝgl8�
t�=c��4�Y"OnTr \0�����t�Ђ���KMٮ�'�M�p.�yY�U�`)���{LG�^�����ݢ[+ �-���aW[L��W�B��cR��jf6&\��&.V�F�LJ�ұT����q�T2�.Y�2�m�I��m
�Ve�-1q@�bLfe�X8Z���.%s(�B�U�kR�[R+mq�]��M.b(�u�2ҫe2�*�L�]S.a�� �²���u+����u�SM�t°P��\�+JPP�t�s��þ��t�
'ҁ4�ۖ����jI���:���Ǫ��Ǐ��1әv�G��Mw�w�����ob�7W{�3�,1@3Zڙ�hx`�f�
��w���
2�hB�Q��jΝ(j�g�kN������A�Xj7sг�)	�$��gr���Lc��Y�����ha��צ}�"y�=�O��8Qf���h�(kϞM)�a�q��W��
H3���"��rY����gKh-�#W����f����
5�l�:����̧m2�{N�]=�{M�v<�s�f���wu�6�Ӣ���L�94�LT�աM����(s�ie��'_^��V��}�xfFӑ$?�� Yh��6k��
ɺ&I��E/p�.�PfȤ��|��늫��s�F��b���M1HA&�԰^4���?5f�RHu�[���T����d��y�N{M����8={Nag�Xkt=.��2e��|�8I��r�L`L�6��#�P�pw�s�8�E�j���@^&zv	�^-+�'0q��@:Px�7�H�B�c3]
6�Ќj�#�dRf�+�'`T�����-�>���$��$Imz��G�S��.iC:A$i���iV�+�Bs5�MX��|��F�%j��L��D�Ν�V>*�V�(������L����u�eb�0,�y{\��!Y/���U���l�VE�t��xh鰦*UƮ�n�)��j *
P��Nj�!�¬|Ů@�,|�Vc��Bl*g��¡b�-#&����jh�Zd��g!Ǫ�p�L���8��cE<5�~�HAa��U��ue�C�s�$}�didq�J0Fh"D$����M1�x����-*�p�Mb� ]����(�!�ӄ�;1���΄�Bm��,�h�|GMs"�|�������೵�z�����t��s�;=y��i����)�
��v�O�E���I���l�Y�}��(� �������	!=�g]i4m�Y�3�F�zL���T�W�(x�ق�^�!���+ց"�=�0���҃װk��ʊ�@P*�۰����ʙ�OW	�V��h᤹h���Ծ��#W��
��N-|��mR�5�&��K����>�D�E���ha�H)���ۙ�����"���p�p�ɨ(������X�6F<���#�:-Q���3���-2�664�## u��Z$A{td��C=���lDp�Y�B0�t��{�+��7.��[NVAVdM�ӣ
mC���v#$��}_g2���yr�]~�ʕ
�Ӄ'�SB��ϻ��sP~����D)'J"]��C�8,�\�q��dJA���G��Vx�\��S��Y���YцH���|�@��75�f�z��ha��G��X@T� tr�Tl�f��(Q`�}�D�j���!X k,Dz�^2(�63P64���b �HIs�ו��E���4�g�YӃj0�hi�����-�;�U٧���*�T���ث��b�s1��ϸ���4x�4
!�X'j�� �畖Ti���LX7N�8�`�?{���r4襩>���R�V8b1ڍ�r�eA���U}G���_C�o�bO�f��b���Fv�(^��ڼ�	��m�"H�g�7`]�5�͙"��g�x���>�[Ԝ_f	!��QhBl���4n�a�t�˖wO�u�h-Af�B�͛^�;N������4����Dq���ƙ�[=��a����F��WZ~(�n�
0A؀�F�㓹W`����d��IW�ԭՃ���4)��{�܀V
���:Yx�>�U���((0�NP��¢)��T��(h�kV�+k��ɷ2����1ڷO5Lu�9ΜE7���g��*���(K<һ1��]Gۗ�q�۽�����cf2����Q�c9E�g�k?\�{v�o����Δ}�a��8�.�	�U8�D��;g���\h�}PA����*�֗)yWu7V����*�FP�����[��şol	Շ�x��YG�
�SOs�3���� ���`�v��3fk CB�L9N��m6�`�ўB�Q����]t�F��'�w��g���+O������*{�� �tn@�d�0|�4E���Fw9V�H�C�װ�
Xk����0؂��r���ۂ�8s3�j/�����Z}�9Se/lIy����%]��.�0l����/BF�X�I�����ﴘ|>w�����SO��G
�t ���~6�祐�S�CW��6!ℵ��x���ffN:�0|�RĪ�p��x��h�G�=2�6E��8� �H�������Ʋ��	�i�uzR�F��+c��u��'CT`b'Lj	�Q� ��2z*�puC=�AY�g�5�l�B��f����\e���XF`�� �(��]p:/��tׂ+��)q��ج�جUd��q�����hF�'pL�N��}dm� ^קw�b
�'��~]r��޿S �����5��D\� G�oH/v�5�:�Q��?}U��s������ϻp"�0l��=V�p�CS[�#�H�
�v�b�v"�����u��U�ia�q�_f<U���/��\�ݎ!�&
"������[���=�
BC�;�V�OK5��X1�QgK�!����e�&)xYd(,�'��C=�j2�=&�a�&�z�� �x�m�.���룖Y�^Yq�y��t�� \j�7�lu�o�+���V�Z��BL�8D�E!n���g��F����������!�N�"3����q!`��\�3��#Ar:�F��}N�}Ko��ӽI��5�\�n�옧Z���� 2+[�	��օ|�Z����Pq��r�7���G$.�2YMa�^V���Xl44�s.�͟g C*xSeTJ�bv*�k���@��Ŋ�W.?Jw�E�\5�WQH��v����%�h3�I��^�1�m��{���{H��4��r�n��ˠ�g;���:^�aY��:���Yr�Z�&��d�(�HdY�8�,��,Z�F�3�dD�D3 �0�%���-�h��N�0o��ن���Tx�WT���^�d]uޫT2n���9BҬ��&��wB�wY'�K�J�)��mv՝�����˽y/d͜��6ţh�&�zD ���++�ì61��WW��x�fv����d�S^Wh��$32���G��XM�������H�[��ɨ�}.�����ږ�:��p]ә���N���2���	[������K��lr�kR�Ŕ� �,A&��!�lE�u:�c6��h����]��
�� ͑��@o�eR���Ǯ2�=�H�9�ۖn�b���Y.��6��AWp3�Zy.i�+�	؎TeSy�Fc�7�D!�� �k#�^�(<����!�r�K�(�ۻ�Ualb��Ώ\�o'G��5V��́����#���-�Q���>2oh,���4]�U��Gm��:cP6�]�&jv��AW�&G˟,��i���㓴`����7��y��{chp�Í��Qw4G��U��;7g\��է"�۬�p&���T+ܔC;+tU�A9!����d�S%��mɘbu���\�(�JK0Cu�u���gi�ެE�w*Zȶ�;lӭ'��uJ���C��Ĭ(划�f8���uh��Ӭ�q�aKV-[
[E-�V5��j�`"ʊ5*�,��(�ڭJŚ�+,ED1.��0ƪ(*���4�J�-"�-m�Ena+ej(*�nV��aK�@�i�b��5�j�|�ˣ`��Ų�Xk�g3D��/����x�峜?.��:�����0l��Ha��*�c`�H�ܰ�g۩$�[���Q���n���}��"��C��#Ada�X��t*�u���Y���J�0�z6^>�9�zq��6��H��J�}X�.[��=��O5w��z�`2	ӄ�E�F:�`U�u-���Ӵz�b�`툅Ƒ�"�d]su�����/�~�"�q�4h������ign,U=�W^8�a�/>�_�BE��k)��T�xb�X*�A��
��٧!^���=����7�����f[���b���5��'�<�v̽E�RE��.3���Ͼ�����~�Lg���o ��*Y�q��D`�6�A>����xgE�"A��E��J̟<�y��,�
��\l�Xd��l��/R�c=���z��Rp�97c���+4C��5�<ũ�Yf8�̝���㤛E�����3Ӳ�;�Ѣ��*��M�Vx�S�'��p�~�]B�$$XZD5�Ì;���u3w�P�����b�$i�������W�kL����h��Y���J�2G3�r�49��NkQ:`j	�"H�=;Ji�6��o���Nu�A�\c�le�7�e<�ֿ�)��y��&-�5�1Mf%	�O�}_}����綩����פ��|~5�����i�AP5"Uv|>��Y�@n���6Ԍ �l��m� ���"����!� Z\C���E=�:0�j|�0�f����ݛ�.���z=���zA�u�O��);(Y�4b
ԑ�\Q�$�,����LMї[c�q�R'P�@����>�,�F�wHv��Dae�2�0��dE�q7!���>ܖ�S��0x���"m"m
H�|���.kY��%��(�Mhc��{k�����;L��h��|���ݵ]yqWo#����Tg��Ƹ8�W���]�#+_LJ�������l�_t
ńA�^�^p�R�O�%M�7U�z��h�ZD%�7UB^�2t�޺yڭp��*ѣD8�b�T}��.�ug����0��t���Y��^�OG�e�H%:`4+PR:�A�5����vubFO��4�v�gH�Vr\F�Z���h��}��iRz���Y���0,,`����"K>�}���:g]��=Ϯ�1�uqAP����Ƒ�����)�[P�8>�j�J� b����c;u,'euu��TBQW#��	+�����X��od���_Dud'2�b���w�����m�τÐU�#O��a�f�-�L��s�V��	!Z
��JY��*׸��5�FDnG�" �/
!�5'���a�9����bř��1�����=F
�k�p�5��V���+Q���CY��D���Hy!��n�6�Y��]��ݮ���
0֏��aa����`�q�/^���Gi8��*���'�����9�7�v��]mW�>0hD@})���*��|�]� v�r:b�ɪ�k�
V�85�8*�oڎ���\������oP.V��7M:Ye�q��S�z�sL����������9�>�`d&t�9������)������sQ��,�V|�"�b��81�Ooyv��
B
�S�t���Z��F����.�(��+��pٳD&�P�C�ZS�օ>�1!꫆�b� W�*�
u5V
��3E�d�'�PE�m�	�=�r�����G ��gm
j���{c�r�م��0U�/�
���Պ�OqR�����(ٕ�{{R��)	�	��#>��M�<+5p����>�[ƪ +G��B�C�E>,��gDfm�����Vj',�*�ÌG�o*���.Ԙ�>�/Rn������1'����������qC�<*���R�%JQ�\<��p��f: aƆ�>I�,�c��ޞ�F�ޮ)z�Y��� ����{�����j��#xl�G����s��Y^F8�?v��b��]�����g�D��p��q�]U��F�WY��0�2$�=;Hua�`\E�O��s��qݸJ�{܉�u��=n��{:LO|���EA{)�^g�Su���u�y�S�N�Β�n��vIJ6dL�	G׻�.����$u�g���:y���t��dQ�[���OG�GPn�P�HuT���=�ʙ<s:zY7#�uoۥ����S��iߋ|�p�����=O�*��tEiܥ~���e��2h/�Kך$�[w�Z,ya�-�r����^�Suxh��m���=�n�9Fge��9ؖ:{ñZ�Yч+�VƦ�})�EݵQƗk��,s-��^����wF5\�]u�;3]j9ڋ>�k��Zrgn���1F�0&�s}��n�fTǆ�t,�Bz�<}�������׶c^M��Q6D���'��;�MĶO$OU�`��CR�)we�i�G�,� ^�XcQ����w�e�S˨ǹ-;ݡ=�d�Q���c�CRw.�bؿVi�Qt�����C�:X�]�[1�R�惛RAgy2�6���DI��Oy�bq٭�&4Y��$����̄�M_Q7�Ř����zgL��z��J�킹�7����au��n�ިC�����ב���B��H;�v�{}u=��$��?#�V��f�#��s�ۚ���Y��Y:w�!w�j��]9��ޞ�b�n�x����'��r�o;��oE"[�hq)�g^�UcD!b=���*e,L(��o⑬�(��m >���Hf��[n����PMTmQ;�;�dѷϤ��a�1×Ċc�^.;���mb�����%������K��q;�"��vKZ���9�r�[L�ם�/(�v���spɷ�+c*۴.��B�,HTR�g�Y&�.{y��E|�+e7��MT-A�f��Q-Q:���˔��=^>�T�b������f�qM�r���Gݺ����ښ��O;H���t�S��n���3�˻g)�ݹ+�t�v�׹|�Q&�/�+��f�7�=<��K{�����Cla����3v����5t��WS���\f�Ճ{&�WX��*��4���6;�2[�_]:�	��t�w��^�O��u���8�P�D����M���e�Kwd��o��u�[�blr�>��[���'o������A�Ge� �g
��z9i�Y�r�,��Di���خkT�Sj���N�G�"�r�ع���"�A�Tf�6��¹�ջ�^��f��BE�<�:�$�������_�2<H�-JT��1U"ũ�IM��\�c�1Z��q�a�
1�p�Ie,�B���r�,�K�j�m��SU����c*b����)Jl��V&Z�	b5QG
Ue������-Ylr�Q�*��Ub%�m��f9s3/�����b�Lٳ�p������\2�e�qǄ����^(>G|�w]? o-u�z�b{J�Rf�[�^�.��3�6�\E�۔�Ss���A ��_���}ҚR6f,u��Ӷw/]RJ�;�U�/�;[�ۢя���q�n�������%���|�kE�O]47�%ſ:��
9�Fv�T[�Ѹ�����^�{��Vݓc�s���Q��>��Y���1��J�tҶ���'��F�B��= ��㞯r޾z����v�[��5���o4��j�_{n��6�zA���{��<۫�t��ޅ��SZ֙]�o-�o}���=$�|�jv��C.�	��[��S��|eE��u�=���f��̻��aG��8fޅ���ךu���"�;9��̧f�J7o#&�J���y�#�e�4��W�����_J��rX�:�j�((�3����D^�ޞu�����|������f�y^YI�i3�qjT�:n���:j�^V��wn�G���,Tq��FKS4��go���	RƕZ�a�0+��3Fn���.�4x���K0Z�:�ճ�|��*ǣ0:O=��5R�re��Z�.[<���Izz���0R���]����\4����mDE!���������w{�cx��N[�'q���z�?#�~(P����p%֖�ۡ�y��<b��u�QMg��-��H�g�� Ƚ~6���Q��#���(m�<��Ÿ�,�(g�v�>�4��Hz��ޫv��Ԗ��Tm��7�h���S3��Y�*|��!���]�͢�M�c���:�b�&��w��2Rz��ͼ��e��J*�E��S�)���J�NL)u$,�Wܚ�<a�����ۺ3�^O4V2��֦�R�څ��'�y�10D�s�όO=��˨�B�.����g�Ϛ�}�&���'�3����w�m��rw��������>c�T����w�յ��J��։ �7��t��(�Wl����);��%@U�����^��[Yj���.bK�Mۮ7�A@gv��®��J�sU�#R,f�I���S伩�$���W��k��	��.W�G�o5h{\�����}���'���9B�aʗ/v7,���3z�����s�"OS�ǲݶg��u�W�8wMm�w��(�&�:��묭ð�N�������C/e�lI�BR���*���(Օ5h�z�*�=��Nɭ�����1C�~�ڏ��aN�������F��\H�f�z<���ɝp�� �ڤ�Iu_OA��k�"�77�5��j�Ⱥ��a��߭���m���j��k(f8�o<u����,Μ�ݾ�&�Ǎ���>��z6����FC�n^s\v�x�ֆ�!\g��.�uؓލi6�t���Baؒ؍����4��;�a������Y7)_�w�)J2�n~��9%��O7��.�R��DB�z�f�s�*�<�lA�S�����ʎɊC��9�Sx�~�� �T¼C��w1��|�^��v�`my���o���#e�p7��A^���������S>�
\�؁�ZF�ļ"��&�K��G;�k���C���iy@[;����v�]�wK��8�v:^���7U�� �oz�%���ʅh�}jY�&��/s��<igb���J���PQ<0�.[�����n�eփ�3˯k�屙ü�T_[3TThQ]�C���lχ:ЎN��wJpe�q�tmRzb�������v��}���[�B��e���4W=�gNZ*���^��j���[�Z�_'^{�k�w�fXa�]����(��M���Ԋ}r��3=��e�*p�uu��Nga��ͻ�{g�fj](�:�K)c���iv����K�iU�ٚ�\�(ξ�ޥ�j��`dHuN��ۻx�cfz� �^Zَy���֥���9�PbCH�����|��������������e��<��5{�Qf�P�v��P˙�Z�p�k�b���FK�J���kÔou��B^����|�6zq�D9��rܷ�S�:�=�k����
��'6}:ج��X� ht;*om�>l*벜��w�5��ӯ4:��	,���Wm�5�q��!�;��@H�]D�&Ŧ�V]9��F��$R���C��az˰{7��'R�%e��TH4,�6�L�����о���Ӓ֡�V�wn7�s��_�\6��V�"�f4Uo`koT��F���>]��;�r�u��]�G)�J��O������c���+XE����-ı�n��1+t���e\<;��ؕ��d�0�\�+�@K���u�Gv�ogF� 2�g,7�W�k\HӇ�NX��+��V��U��ܸ�  Sy<k.�W��!S���6w��1\1ǎZ�i.�Y�u8s\�k��7���w���+h*n-��X8�Ԩ��5m��T�I��J̖�b�&��-_IG�L��F�ޏ+8Qorq��Y��gKX�4o-��r���d��D��B�'v>!�Z�l�As�r[��7���.�l��\#��sX"8=��Y�C.�ڨ��55�j�u5�/7�9�7��*(�dY�U��̤.U�LT�1�s-��$���*�m�� ڴ��F�"
WW2���V�r�)J�mpG-�
9���.8�Fb[�[s)���a��S-�ێf8	h)���)��f����b��-b�9�QLf%	�N��6
,�ofP|^%u����O�T�C�'D=�5~����L|U��Wo(�Ű�C��dv���4u���)v�1
�ɷ������zk�}ֆAݽ����S=��VV�<�.̮Ƌ�'��-��y���"��k�=�$�}u��ʓP��Ί�Թ��N��Yɂ���컜s�;��l�剡��$��GL�g\�W�ԉ-}q(V�c��d��5�-�s����;g���7���}c"q�\�Y}�2z,�26���AN���+�ٙ�Ȑ��޼��30��{/objq^�0(��nX����ã�x�:��>��t�.�x�#�6��	ҋ�I�WU���ޛ�Q:n�2-�#�FDW9� �/��8�ɨ�z�����F�#G+��x*�MnIM�ĸR=��!9�
�sy� 8�Ve�wY$זTY�Fp�,�5��meD'�y/��S�+��p����\���{�%ge��+*5��4��QI�I�+�:�׵��ֻQ����O�W���������8�/�%�y��u(��z���J����_����D6K]i%�����1-�x�Z�qg��[f3���Y[u�@H[�6ː)�,�`͸��e8Ƴ���M���������ӮA����=��'�0�Ã~�w�3�h��o�������_.L�S@�H��ɡ��2�W3]���]xvF+tnҞ��1�5��qY����5��X����V`���Aݎ�E^�J��p�Wx�����"�S)RA���	�u����5��S����LC��2���MJ_<��s��L<�u992���I��K�;w��-�"o�`�ı�t��.�E�4��y��vlQ�s-ݏ74�h���R��zj�Ȯ����ivVN��V3�I6��2hY��ॕ����t[Ou��F.\�A�*7��ͬ�W�Fl�A��fiY��(�8���&�''��V�w�u5��ȳ��FE䆿GՎ�-�=��Ί"#�.�U�KXv�r���׫L���NrR	C�@���EJdL��M;~�;�򉺁kh�W,Ŭ������O��h��e#u��h�x;����^מ�5�6懒�y�r3 ��o�Wח���}��M�p]�;j//\+�|�.;2d;ʿTM���?���Ia^�Q�1lE7��V�Q�^��Ç��#�q�J�⡢����s-�<��n��)c��k풖�V��0�j�ك�d��X�MTQ���%�Jpo/ԎR�-��p�����9r���A^|��V���i���W�K�X��;�em�V�z\㲦&n7�
�BSۧ�ý�\;''�/ZPOd����S�K5Y|wOl�j�%]Om_��W[ug�x���{�Qqbqm�X{�,*���^ƽ��sٙyǕ�ѳ�.��2b���X43$r�
B�m�&h��Ft7�j���)a6����'�
����(x{^X���D	z�YY���h�U���]��W�t�4s�ҩ����f��f�j�b��J�d����/]���Os�yu7U޺�/6g���ڠ&剮x{6��N���I��T�v�6u!V)�&��W��V1�M{bܦ3�^���M�)e������v0���k�H}��w:o7W�)k$9ӞN2���N1���[�J�V:�#����6|~0`��*��ػMl�r��$��IS�-��ӝAQ��ȩ{�!�P��<,�vF5�A=�Q��)�5���!�˚�����*S�m(�S�5w{s�ƛخ���S˼]X^�a��N�;��ؖ�b��΀���}{}������/��Z6��]�v��������j]� *��x���*I�Km]��C��Ȼ��❙���3��;��
��6TM���3"�jח��Z7��;�|5t§��-��gpֆZ���U��n���
"y�쭅k�<���Uc��v0�Yf3���a_DF${]�����磉���<K����v�n�־�60�Jx�u�y6�����ΰ���Lחi�d|'g�)e�Va�>�r��F�+T�cI�mŵ�o:�Q\��a�Cq%W us`�K3iE�Y��>KL��ݏJ���Ղ�BΫ&][Z\�%�Y��AJnm�I�,\�b�N95e0!�Uk��N�7[��A��ڞ�sb�9�Vj[��1��.�Rmc����~���'R�qu���6u��K'|��&�7Rs�VD��jci��iƧu.K2�G�rӒ������˶i�~F	B#�om7���/C̾��<6�Z���]�OC�ok�R��`��=.A7a\,����C�ڊ��arQ��we�'����lUd��׽@ՓF�L�y������Lrb�Q�;���(��Hu}�V{h�nP �5rD�z�T�ly[�1Z'Z�h�.��U-��f��i<�FKm�ٙ�r&Ns*��2�w�kR��V��͜4��=��L�e@)�2�ΡJ�0�5Z՘j�\�3T�$#6N�&P���dFp�s��(�w�|R��Q�p��v���M�`�Ó����Cb�}���7О�n�n#i"����34۬�5?T��>��̵�Y[l�Ģ�\�T�ʵ+��ڦ&[�1\cJ�G�����@�-�JfV���
�kD�Ը�*8��(Q��J*ԭ*�h-�ڣlm̸�����V"�imF6��pD���ZъT+U���(6�De)j�T11�E����W�G�\��� ��I��r���9�����>����үi�=����ӪVc��n�_U��6}p�{-Am��6�*��_��^�Z��G����yG�#9=W��o�m��Xs=~�WT�Luݛ��XX�/�!�v�]���mո�-����ނ,�93)s�x.b���f(�˂Od�+)���
��3�ٳ]S��d\�5�m��8G-��GW����r┱:�2�)�8Gq��/-7j,�#t413�c��%��-G4$���ύ(Zy�ٕ ��M���Vy�%I⣔��˳Q�߼oc�|(#���E�j�z�ls�cTh�A�/_��n�˟6�;�2�O>J
��&<��!���74�r_g,~s�Tk�.���s�cH�\n��7![�'p"���ܬ��ΐ�,��[Sb���ͨ�L���by6��Y͉�2���G'(N�]�]���-D�����#W�U���;ݻ���]�T�����;g�����9����2w���%tV�r�;Z{!ݣ(�坒��g�}S+N�y��ww�,k��g�~[��Vxb[��s4eR*Sz��!եD���Mu���!�{c/0k"�7�]ޣUG.�MK�*N�����1��fb����X�;8nn�N���Ŏ2���=�Lz���q�l؀K�g�q��g&�uP�B� q�����0�u�Y:�;�FS���]�N=݌���'.��ˢ�kP�济�IeܘsƮ�m�Ù��w �f�� j;� ������??C��G��׻��k��d���!}:�Y<�Y=XBP���{7WX��i��*�H�VK��#3w�F��H��?/M�w'�ӻ�nͨ�!��)/9Ii!߷7��L�f\���^M��;��֩��.S&�$�ޫۺ�����z�w�m�ŋ�{M2���0H�Z|��,�j��2w�s4v���嚹���h��"�m�º�T���`��y��|�}��d�ڞfF��͖�;����~������#�Ѭ�tL�j��<�gMҔWn*k{������Yy^���������%9\GaM�v��b�����)���:)�p�r������k7@���f޻��Q�.׀��i��޼�\Y���;��g�J�Au�<˾���C�{v�ȗ���[�a�U���u<���g�Պ��f�%��Sen*u~��F�w�0Z�1%9���o��r��kv�o8�����x�[��d��/�u�w�cM��'�V��� B(m�U��1��]Op -D�F��n2�F�5��Y���[�+�� ��|ߪ?-�����f��!��6]���X{���u=[����CӜ��c�^�R��C[��-r��0�wuP����{�V>ڝ�;�q�9j�S��)�k���j��K��9_����Z���j��쀯ٹĝ�]신��6�W+�%�
܅�o�� ��0{ ���yڃ�I��`�.��T(<�x7���DuABX�Q�>���f3�Mޚ��6K�N]Խ��Ι��]���xP��\��k�q[�c�����isƕx�#a���]o��ЇK���׶�ǳ��Ƭi��-�"��Yuy��H��,ɔ���ᐼ>܏�q���ob:��!J������_�Y�D��[lX�eb�u6H�G�ׄ��ngO?RҨ��]����*�L���ކ^m�����d�WJYR�$jE�ęJ9�9���;F3��W��������iw����XNB�3΢�咵:�V�I�m�99�e	���bX̧�|q�/�!(}�$�~��xm���B�;��p��[�r��Wy'�>13�5�v�u������,����ddӎ�+-�x���>d�h����s	Q��^8�-���
^�ݮY}W@��ܺ|8�vs0�$钳m�1,O���s�L����9�q��twWF���.c��Z�$U���Z���Fkj�5�W⒲o�7�WDy�[UE�D�m������O]ڻv���7��Y�ՊYuO���k^��v���A��̘�k���I��7��s�y���Ѕ��R�x�Ei�S��ggX�2r�ؽ�-�D����?�� �?J�������HC~��@$	��2� ������D\��Z2҄�|��Mv�����G]��=�����5�0X��|�`$2�&P&tK�5�t�fVtH{�p� ;����Lc_�v�v�������N/��൷T��V\*7�m���y�rh�ϗa������Ӡ�[�߄O����1ʽ|� @^�>Ap������	+C������pn�{��>�$�eL?����Yߛ�B$�@PT���˷|18�iw�AKu� .x�]��#a�G̛R�ε	��m�Y�ٰ����K���v?�� PT���W
N����(�Eȋ�TE*	����Jl��Y�9zؼ6L�Ҧ��AS&�����cm�ҹ=r5I�G��\R���nb[I���t�g�Y>��N�����&\@PT�&]E`y&wp���5}�\VOq��M Kz>|g�2�ÁdضC��u`�$;K���m泘���ya�ìb��Ȳa�g
ޒh�x��\�,�H

����у��'8�Wm��D�P�q0,)�e�.3�����q��0:��!3�/AT�č��Wi�.|�)�D�,��OI�;C͝X�	yQLZf��v��H����#S�P�=O�!��4l2�h6���;�����,|N� (FÂ������)��kJ|v�^���(*u��k6F�X��$��0H� PT��[��>���a�A�r�Й�N�hf�4�K�n(�xs�@��H�<����ywi�-w 1!������0�{���[>�; (*q�n,��nH�d�r`A��X��CC����}ӷ�Qd<R��ip$"(*L�O!��ty=<�m�\5"(*p�Ԑr�7������-};��Җ.L�"�|IW���ӱ����H�
�� 