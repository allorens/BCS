BZh91AY&SYح]8��_�`q���#� ����b,            X                                 
��� �ت�8 J�o             h(                     oz�^��*�!"��B��BE AQJ�D����UIE��EBH�D��R�UP��UJEF甀 �QI
H
�$H�V��T��(�b�:��tR�H�lO����NmB�b�]�H)�tq�[��    �Ð� �(�5_�M5J�w�|��=5���/>T��һev�׎�>Z |�������C�]�%+:���@v��=� z� S�   ��G�  >�����Q
���%T�x >�s����{���'��`�^��=�8=��/0kס�{ �/{<�N��w�R��A�Ϋց{�@   ;�ʤ  ��`	�=��
/@nÞ` u�=���� 8��)�=�� �`yz=�<����  ��� c�JTJ��(��QT���X���8�y�=^c����z��K����p<�y�yz{� �P�p�^@=��   >�� �=�t	�:_p�<��}�{�>�y:�z����P8 ���{�����oX �   ��@4���*�����.�J
� Z��݀� �� �pP� ;�r ��:���8�w ���X ��@�8   ��!������q N 2 \�T�@�3`]��t��@���΁!� �   <�$  >��HR�$�� (��� �݀9�Y�R���: d� t1 �B*p �� `)@ x�H  0{� |�� �	 6�$�`:�  �r	. ��@��#���         i�L)R)���00h��10��D�����@h@hh@��U"d����    ��T���4&!� �IE�(    4 
P�M���Bm�2h��?/���o�_�톹2	?A<��9�@�<�n�s|��E�����QAO�������������G�����?�O�>���o����E��2��� Q_ɃГ�}I�*����?����S�^Aq�r�Aq�GA�E
��%A�@\dQ�U�A`Q� \dE�$�\eA�!L`��Dq� �U\e�TdA�@\`�\eLb`q��Le1��S\gI��Le1��dq�1��`&\eq��G\eae1�a`daq��W\eq�1�e1�1��G\``eq��1��\eeq��@� �q�q��Geq��`q��I��G\aq��\aq��d&\`q��`q��J���Ce�1��G`q��GI�dq��Ge1��Le1��q�`q��SLd1��Sdq��S&G`q��dq��e� �aq��\aq��e1��	��`q��GLe1��G�fSe1��SLe1��SLa2�Le1��GLe1��L`q�d1��`q��SLeq�1���`q��Saq��i��\eq��Gdq��Z��q�1�1�1�� �\`�aq��W\eq��Wf\aq�� �G\d``aq�1�	��dq��G`q��fSaq��dq��G�eq��\aq��i��eq��`q��Y�`q��`q��Ldq��q��Le1��Le1��Sa*,e1��Se1��e1��Bd��L`q��`q��SLi��SL`q�1��Le1��e1��d1��Sd*#\e1��`q��Se�I��Ldq��Gdq��&``q��G`q��&SLdq��Gaq��	�`eeq��\`q�ƙLdq��`q��W2�	��G\`q��\a&1��`q��Le�1���e1��Sdq��Bg`q��L`q��G&Le1��SLa1��SLe1�(���eq�� �G&dq��aq���Ldq��eq��Lf`q��L`q��SLa�$�e1��Ge1���La1��a1��CLq�&S\dq��SLa1�d�Se1��Le1��S�Rdq��dq��a1���1��dq��eq�1�1�1�1��Wq��\aq��W\eq���GJ�\`aq��W\aq��1��\`aq���`�Ldq�1�1��W\eq�	��W\aq�1�1��aq��G\`dq��I��@�W\eq��� � � �@�\d`q�``ee`fdq�1�e1�1�1�� ��Q�$�A\�`1� �C(�Wq�Wq��$�q�Qr�`ɿ�@��Zf�p4&����E��G���2�
��K���h�G�$���>�x�v�c:���N>N�s�]��l�3J�=���F��ͺ��C D�Sf'���򈪇Y(; WB@4�(W8��7yM��Ep��j�n�Ԉ9b���Y0�g5�Q��d�.'ع�SX7�#����jJ'ܱQR�╗uIe)�6�����\M��-C�5L��L��P��<�9��n��k��& ���5�t���d��澪���ql�ذ�Ղ�'�tDSSJ,2���ֻ\�8��Z\w8nIخk�����W��2�r�q�8-�J"�֦�ls����7�]]�vEV��ӜK°�Ӕɽ^���X��b�Ȉ��M���\���z��y '*��;B�%N}2����8�LK��X�{�r�[1uDWl�;�e��nJ����P���k���r�;�+$/����E���{���խ<[9���t�{fNBs�ۇ���y�g�@�Z6�u3�yS����y[�U�v��P��{�"4���0���h�]ϒ�t���*��7j��Z�A��b6ۛ:�3�a���x�Ad�M�]��w
I�>�ygC��y�ƭ㻷��V(��@�K9�闔4P�o^ ���;����8��`�m�C�{z�ʷ+�T��q�:��܂�o��߯.�>�&3�=C;&��b�`\X��z�LjG��_5aQ�7��ӌ�v�i�G?�s��$��Y6*S�2�otFhFmWI�0IQ:{z��ɋ8Ž�8�SN�Ɉ�&��Q�+�܇��y��>�4�kx�śdW4�M���5[:�ۤ���6�V�7��U��+�)�t��7Y�=q��a��V�h��K��R��	`�g<[ض-&72�v�̗77y=� �ն���������i�����k=�]�� �V�C��|�6>)��~��[�˧t�9F�'�7�p!� Q�za=�!��v���]�ZuPdwQ�M�̢m�Y`ߦvd��F�9�CLp��c���7���:.����-�{�v�u���0a9�O�i��p3t]�op��j��"6)-]� ��:���֞s���>���6	��qK����X�rm)]�M�fX�.�9;"Эy���eɝV�T��y:P���-�w�LB[`���qɼ�bU
�l���S.T.p�N���뽤��:�%��sz��j�ۅ��jڰo�c���x�/|��nu'w�ֵ�q�B�5^�`���U�۴�:RWK/��Gda�9�;��$MwyLC���[v�n�#�wO_���Ix�����Vf��;p��x^4�ǌ=�L����[1Cù*[���6�q���S�\��w8u�ݗ�yd��3�hLU�m��7�׳�{�e�Zώ����3w�1.z1X�;����������O��%l�Iq�-R1&gM�SҸ��N�U��k�p4F�v��-7z���H7靵���Ĳw^H#��aή�4�.�:���Ǟ�3�-͇�oC�gH��5�1��i��n%����YC%.gF��+``Ц-��S"�rYb6.�.��t���`��ݬ�[������4��k�]��۷LYؙ3"ޛ�u=v��6���J7�ʔ��2�-ä.��v.+���b��GL��������SvKA�V���.=ۆ�����ҙ&n �;��4<nI�h��Ű�os���ަ�������.�s�0�\M3u<�8�`���is^���� ��X�JR{s�O6AP��f��V�kԀ+#�&�Ԝ,�n��j�(�|���tafB..�t��3K�7�ޓ����j(ɼdk�Q>�:�h1⽴���d�k9�Sy76o�h�M�z�ÔR��wec�:b�Gd!3˖t;�KEc������GF�S���;B��tr���5�<�ӐG�GN<���w�^ǝ�,��e�9ې���Y����I��E�=wؠ��4d��O�T�eˊx��rtW���%dX�!�'O�l[P�.vmpq�p�$�J��5k�����B�0f�f�Zy�����b˓#2�#I�ܰ���,(��y��@]��ih� &l�sCa8�<gp�͋�;p�7;����d���ά[z��If�چ���HS�2ԇ\νۂ��뻼�sX㸴`I��E��v��f�֗ ��z�"�3�
d�
�v'�w6��B%Ǘ��;��M�o<B#�R��n
0��qv�nw !�z��ݴ�9�M�LZ�f�>}�o.���@��sut���ӄ�+���tpV9fԆi�a��٠�僫r���XI#���Kv����Ѹt��r�K���ۑsv��Rt��u蓎�[�n\�.���m%{.O����Ӛ2$�B��jNT�]Å������ ��K�{q� �.�������n��ϵ��.�s�~3�W85�R�>�&B.v���OJ]�Qk���Du���	&�9I�<�v�c��)6�<4N�PQR:�l�y<hr؞r�7:+���	p�$GL�����7hj=�Ӽ��w��,w��>���4{����/}�pZ9�loSx�զbNo.�ݻ>S���.��5v^��wU��b�%�i�T�YV\u#����mv���� 4u�P%VF��5�/�`Ug%u�݁i�B+3ynh����!:ȶ�sw�ް+���M����'�5������!�GpVߞ�Er0IR�#ӳ�ݚ	�;Nt&
��W4�ֶmf3���|Ԍk��$�q�0�tke0:��щ����4j�x���gg}��=Ug^W�/wz::�I�fᦡ�>�$�R�]Yz�#MU��S���Ë��}�Ȏ[�8�Fsx�B��:D��c8hm�Z�w`�t���뷖':��������xQ�J��-�<�Q׎S;�K�r�]r����#����k���F�Z^2Xy#ߔ����
ELޠ*My�m�Z��6oMXk�;�;-qn��t�e��M�J�{R1��٫s7	(�>����V����1�х!�o��#&�* Ӆ7�o`cr.gr-�t�"}�:w)��s�l*Aș��P1�w:V�ma�\�ON�\ha��8�L[��;�opwyv�r�]�l��s��� ���{�w��1u�q�d�;��d=�����@���mOGA�KAo6�X���;��ܢT#���Аa$�R��4�pg��Uh��˖�$Xݫ�Ѯ�5���R�$
�,���wq)܇�i6\�!A����g7T��<�Vr���c,���D�Pl�LNrq�B.�3���N�l�e��MZ6�˛��Ncy�n�h7y!�ϹwhQ\�³S
��#����'.e�3���f�5���i��f�.�i|�]���{X�]�n�$o{g�F滅&�v���C/l��/Ww,Cq빩MfM��f�����L�S�L�5mֺ��pRDl��p��9�ȬJ�WE����Bܧ4D�����,�:_q���[���TNF�'<R�ֲC�F��3�<fG3M]�܃�!���@v�#{H�C�y=���6��j���n�e��+d;�>R�K8�%�;��tV��2`��DG6먁{�3@J>���±)�i�B�K�{�[��o!"�u�nj���%�#O�cK��1�硗�8tCd��e��wL9���	�C��`|>�q�voVY�4��H��Md�n5�RVNL�e�D���k�M���&n�/Y�o8;kaMҦ����h�=J�2��ݜ{s^,*f��C�2�}�pzp�iKh}�;�Ų�y���e���"ܽ���l�wg
���*ߨ�l�ͪfm�vcٜ7C�s��z�$p)O��ˆ�w�Zr�+ѶHv�9�/y��Q���_t5����u�˱��)�ӧv�9v��zյ�2��k@'`���iᚖ��C�Du8�2C1u!��T!��'4���+u��m���H� �7�^��钊�}oA�㽃$�XÎZi��#}ӱI��+93���y.�\t��Eʹ��i:���]e�Ԯ$]���'�kK�ෳ�]���P���q�;n�=qÚ0hT�Wt�4-x��%h2��͗�Pല-����mtsv.��x�k����Z ��`׻6ܡ�0}�$�B�N:~��裹)�Ѧ�\���S�%�aMN��7W��
j��]��Ago��9�+�ҳqI���5P:�-k�^�qťaX5���wr`�����I��F�"��=����C�Iu�˩,��iO�\{�#C�n���8�\g9��R��<���Z�#�-oc�Ӹ���We��Rw"謕̹�8�Xi�3��6yP��޼�9:�� ����Q��p����ia�ޏ]����6e�o0N<a���ɻ���Ө׶;�������vrG����E5��r��m�fˤ�׽���e��qM�7�Vx���� z�	��!ۖ�s/gT9��Ǫ�
�����]�{��(�Wݧw�����q��ؕO��=Ӯ�ǀA�Sk��e��v�Ψ��t��W���;����rr1�;��ӳ�����i���ʴ���c�_v��P h�>"d����WԱ��N;|^�OCF�y��͋Vnl�ڹ�Z�c��D2�wp/E�]�LaӸ��&h��٨{`�t$�vtZ;~;��d�û�u��U��C͹�`��Jy���i��
�Xԭۑ �8���Bǳ"��k��2�\�r5u��#�ڷZ�E�:e,m���d���aY&(VǛ��T��������ӝ�TV�V���C0��5oq��0����o�y9�w�s\a�;�"1u`�{�WN�Z	_b�Oh� os�M8�M��޷n�z����G�_t{�Z��hx���gv􉑔��F���ɹ+7;~I��~
e�c�휟�v��k���zv�a�m��p^�a�Jthr�{iع�s����PY^��A�:�·�L��[��\�̟�3�f��zX�nT�Շ{�;�Kr�1i�&����؊�˙a�廽�ٝ/ �o3ub�f��%����{ k��P��2�՚�"�=��D�����2�=s]aJ�G�4t�n0��C:��.��v�d��P�ƹ:��qɧ*:s���B�G92����0�����rg���i���Od�lx�㚏q��mu���ЍX�ǝ��N��/j��w�kw`�T�Z$y����Z��y��G�B81���wNk�c�H)��dwBk�9)���x��P1�{ܜ�HW��<ׅ<�xY���"��զv�Ov��������Ú��x!^��a�4�3q�]�v%�זQݍv��v�N�]�9>�.��ٻm����VqH�7��ï�[؍e�YeȟIn��kvV�w��Y���:��:���nI�*�@z�a8�=ope\�L�TPO�oN�&��p����)Ή>�R@�G:�02x�`u|���3����Wt�dC���G<�#����D���v빻=g"U�2:nS�tٖl�rtfMM�؆'M���u�D�]�J�J�Nf��]�U�^�2�V�ι���7���.8�;�LOB��@�E��B���*�k��|�T7@��s�y��yv):wL���͝ɸ�<��t�(�p%K�N�i	�Aڠ�s�]��9!!�b��c�e��I�ƙ��$�Tro�>�qېe��E���e��6�oM,�h:��Ŏ&\vXt	���Lǖ0�3c���w{z9:n�="]��K�;���>IRٚ^I��Y(�N���M'��J�n6�d��̹�=�ωD�i8��ޚM�V�'1>ޘR�<d�ԩ$��%'�<|KdIL�@�<OPx��'��?[�K~�a/r�|��������pc�SOwzJ�dZOk��Oe`��N I$�|V�о�x> ʁ�0�����x?{��M3h��G~g����V
��,�Q(��� �A�z������@ <�7ne�J�||����M%�7I�i$���.�Id5�%�"0Bl3߇6���(�J1��t�c+��,`$`�T7H&`'��pwc�v!�!-�tx��x�f��L���4�9I�'fi-KQ��Y �)$�MF3��K14�I&V_�v�:��t����tK' �4�n�O\k��)��K��2������>;$��hLb�y�Ρ��gݯ`o��S%�n�t�ASN�A3�|��5�[}ʚ�н'I$���������=���60
w�3*�'��퍰V�/{C�{�}d����8�I$�(���>*�����S�^�F%�y4$�<N��/I�8��4�+�I<JI���V	�=�!D��Ƥ�Z{Jq�g0���i�%���X�$�l��M'���;�L�x���2ߏ���L�O��=N��$�aD�|J��^��>��<;��q�����t�$��+B�au�ߓ�NI��GJ��|_��C'�DRI���Q����7*��ˬ�%2H��<	n ��,�^���:�m�q7������L%
�GIZOI��q�x c�ӫ��]|�{,������ǉ�,�K0��5�w79$J%�� �	�`�z  GX�
����f��Z�'R��Q�أ�%Г���%O=7a�v��C�5xW�ZqҤ���x��^Q�FDJ��wK�]^T(�Jk��#�o�����~`�����~Ӑ��3��P@)h (�
�(���&@���B!H �"%���J+@�d����*�  ��H�A��B��B�䠋H-(�R�d����*Ѐ�4 ��@�P
9-"�"R
��R�ЉJ)J��P
R�@�
 P ��*J҈4
� !��J!CJ�B%(d
"�(P-
-(�P�@��!���@� #@
P �J��4"-�*H" )B%(����*��� *% #@�@���?g�^��C~p�i:P z�;� C� C��<g�2�#�e>�-�]��}�;���=�0��N�ڋ0�Ґ��i���A�6%�{��`qy|`�2��(us'>b>K���$�>{��y �Z{�`|�9���u%'Ss�ò�P�u{�/qěus�̞C�x�5���^�y/����s�w�{	�xwܟ'�8��N$��;�� |�<���C�?���w�����q�@;�~������8�����F=������b�W�~�~����6���gX�u!���@w�{���\)���s��̎w���G�,� ��������U������������ @D7����`|��~c��2��_���Ih�F|^bi�O5�0���q��J�(��Ec�W!��~{����Cn��R���k�X��j8዇d+A�f5�d$�}._U����M�e�|��wa�q'����M`;�j$�gpϾ���OL\�N��Ʒ�]]���*ۚ��r[֙my�}
�]�.�gV���>��&e�0�;n��!Q&��\�r�P�x�%���+��ۻ��œ~�}�yU���z21�����N���������óV��gMr��֪Ͻ�w@:n��~�<4��D�>�7R����������:C,m�{�8�u*"��>��b���R��Md�O�L�S�/��'�0Gs���pE���P��>�d��k�3��k���z���q�^}�F��ĺ������y����<�"z�g�zP�>8.�CEўP/ݕ�����;�*�n5��ж���ˍ��B:�A��{�a�PT�y�n�zl9��+u��HY����?������]�_�J)}yxsn�'R[ ��Y�����+�\�\T�o�r��ϳޞ2t����Fm*w)l�<�{����w�״�f��r�X�q��k>�Q�+}�~V�η�OΉ.��R��y���QOS��3q���=��3��G�e ����f�3���;��{������ï/Ƿ�����]u�]u�]u�]u�]u��]u�]u��Y�]u�]u��\u�]u�^�u�חu�]u��]xu�]u�^�uׇ]u�]u��]xu�]u�]|u�u�]u��]u��]u��]u�^�u�^u�]u��]q�]u�]|tu�]u�]u�G]u�]yu�]tzu�]u�]u��]u�]u��Y�]u�]{u�^u�^u�]u��Y�]u�]u���]u�]u��\u�]u��]uק]u�]u�]u���]u�]u��]q�u�]u��]xu�]uק]uח]u�]u�]u���]u�]{u�^u�q�]tu�/�RfJ=���׽�s3�-x�z=���;�3S}�p汜Y��֞�40"��>b���$q�`W���3�:����)b�9���,��p��|�),��I���=#mh��������ន��n	����S��>�����7U)�;M�V=����w����A��$����;�`���ݜ%:B�2x�#��i혩�Ѵ�rY7�LO;tg�-���N�MK�Çҙ�ڼ}�w�]U���o����o����f�/d�]�E��N!��4x���tj��U�t���v��МĠ�ki���\^	-��v��p���; Ow4g��*�&k��ʭ�ƇG�e��]�/u���\��\��Q}-)b+�&��� L�ؽ	���}5ޮ>�t{���||�է:��^{SFB���q����W`�}]�ٰ��xr������lz=����j�o���eVn�^��9fD
g�m����ۮw�x�q�G���hG��!�ϲ!���d��n���L��<�XB�ݔ�I�����s�z�a's/,/=#���A{��>�;�+3��o���=4��b~��s�lD���.���R
2U�z�Y�y��:��g�v����^)���Rv�O���nww�}�����S���n杞^-}�y��4�m�=��E�����t�G���������.�뮺�뮺�뮺�N��.�뮼�뮺�뮸뮺뮾:�:뮺뮾��:뮺뮾��:뮺뮾��:뮺뮾��:뮺뮾��:뮺뮾��κ뮽�믮���뮺믮���뮽:뮼�뮺�Ӯ��ˮ�뮽:뮼�뮺�Ӯ��ˮ��î�뮽��:뮺믎��뮺믎��.�뮽���.���뮺��뮺뮺�뮺뮽���뮼�뮺�뮺�뮺�n�κ뮺믮��뮺�ۮ��뮺�뮺�o���8�n�ܮ�f�-�A=��������'e#��4`r��}�ي�L�D��G�ЎW�${��w��=��n�spjr��ë�(w��K \��Y���������31n�������w��	�=�� =�ݥ��m��1Sp��g���k�3�$!�׫o������CǞn�+�ϗ��Hm��׆��z�c���Zw�����b��ѳ�ۈg`Z<��l�ټ��C��܈,� ���F�w��וyQ�x�'����^0��/<5�jK=�;�ۯ^,�w��spf���C3n��u�[�Ƿ�	��={��]�OW{�8�.�q�r�Bl��5޻�n&��O��$Bpb�ͻ������gQ�W�靠M�N�]wa���Q�s~5yq/!�5��1�)knf�7��
����;�����O{������;�}��k%`ǣ�̃��}��Ξ^��|�/+Q����Ɉ��f�w?�*��Nx�Lg�]�J��ў?g��������Zrߺ{� ܲq�������NZ-<�.���+���O>�a[���<�Bޗ^����=�����Y����K��_;���	?m�1��o�=H����k�x��c�aEhB�I��u}�{n�k@�ʡ��L�<>���|�L�>���������#=�Z���U��秏^
��ًJ�O�dS�{�;��G�������A�v�;�#���a^�+�p͝�.��>�������fe��J'�N J�l��w����1䇄��3�e��q�_ox�k�{����n��_��`�z;Gv���)l���3��WG�ོ���=���81�^�c���/9��1�gn�O��{}y�0dz��$�7�أc��[��p�z��Foٕ�D�����XT�}tjW���gGy�黬e9����F}��.,�z�{�b��쥺z2w��:�o��Gc�Q��D銽�w��J8˥������^O��:������e�����Qs��Io��{��y�6Z��*�j�a�X�y^�,��P�^a	��U7-C=�z�/�dзK1��VY�鋆.�3�=�ď_l�����³��`��֐۳��������)�k�'E�u�8�ou#U:�]�rvg_<�b}��Tk�~ў�]x�"/%�.�&xht�+��I�^#��y�TD��$�����4�zhc��[]|w��y���}�Vgz��]���0��1o���\��Ve��9'2��of���SRo�L�ŧA�쯶������e�>9�a>���ڶ��"��$�i�$|�L�fvy��XM��_z,�N{����"�����s�|;���g�������-馷�g���&SN'����Oy����T`��g���77��}|��S�
[�=�ܴ��0���y���,�}�M���M]���<��`ޓ�2t���x�������q�B���}1f>�����%���:�M;x�^>��5_�'��ՙ���_f�j���;4��Zb�lW�X+���C�8��-I�;����2���~�#�k9�[ow�]�  L�x{v�y <p���cv��~���[�=0ພO�m�/�6��l�b�|;�+����R�-Y�vJ$ ��D�K�6DK$�9��,xy{/�m̻J���w��煫e>��y�e���[�{q�_p-ܜ3����v��}uwPU+c�z�İ�<;�w�椗�=����]����ʹ�;���K�|Ǵ}�l��;rB\ Q���{�سC[�t^�z�<�w���^^1?Z��OM�e�;Q��۠�xU;>}�aX��Y
C�t���,�O{�j/�X�������x/v���z��Pv���ҳh�n�NtOUnr��M��7<a��x��U�����U���;��|�M׽�fn���WL0b�Os�e�6w���yť��f=;<<�o@]��'oO<X ���Y�;�Sݪ��}�t��[��7��Y��۾>՞1Eȭ<����s��|�=_I|9�0k.����5�L�^�h����>��M�;���>��o�r˥�o����5t�.�㜮�QT���;��Y}�oM��4���ڞz���@��E�/��+a��3�����v��+'��LT�@��,��`�#�G�
�=��鴑k��K�w�J϶�|R\�Vd��nK-��v�\�ϩ���q��*ę�W�y�	�x���Q�sH�ể؝���O����x[��W�A��<��� U�O5�O��T�j���:9{췆9(�I"X=Z�ohq��y(���}��\���CW�~�=��o��w���9��o.����6���n(����=�����VΣٮ��'q��;����~��>��3`��)��\7�8I����_,�t�s��:{4ǩ���I'�˽��o���x���eE
,��տx�<��'z���C�R�ZR���ޅ��p�]pz��}�8[$y���c^+Uʳ^u�:��@w��{�i��F����3µ�NO�Y^���d�X�9K��������6d�3Ϗ�܎弆\��?n��禬3���0y��X+>���.�m>�{��c6����Zh�7��Wa��j�c#��o�;D�|�Tv����<�)v�Xޙ�w�ru~��Ϗ�mz7�=��>٤�����-M�s8�z��=��;�0�b)-��o0���/dZw}��}��}G�������o,��BP�R��c�S}�'{tN�>ͧ�z��~gsig�:Y�j!�����w�v�vdo~���F>O�e��#;Vď`����98\��&7���-/���>B��6k�k��̚tz⦛�{����C���Zf��R�b�b��3�/f��,߻|\
4�@C=���x;���g����k��}uB�����xg{�%�c��� 	��"!��}��!�hx��V=���;xGs�V���������`�D�u��4v{,���aKA�zH�_���$C0������9�{�fOs�ù��������׬蟗���7(�������S���gn�0����4f�VlZ�����%��U������\���������O�hm缨'�}�̌��J����?�w�ii�P�٣|R�^>�=��F����}ޓ��Ѿ�y{�����Tq����>���rO���w��y��ݡĂKۏL�"rŊ)�*z�E3ػD�~�f����n� N2D�%��#�KXϳ��8����/7\�Ui!Ϟ��t��E��=�u�=����s��t��þ�y׶v�V=���d�Ϥ���pܒ�^��<�O����>���޻��I�۹�IU�6/e�}�Cv�9�`܏�xe�������oÎOnkWL�&����;}�<{��ӣ�Z�w��ܐ�-z�"g��n,��|
i�=*K׊�޳�#5ɾ����lCWg�^�{>���/����� f�t����z�);��O��.\�y#:�z۝��ǽwM��
5i�Z� �Ѳych���t�{ZWZ܋^Z���F^0�m�^�z3M��o�[y��ȀPdH��tőװ�'�V�L�?>�Z������rԕ��ܾ��'�w���W���q���=���tn
,���$k�)·�������͡,̓��Q�z�{#{)�w��
�==8��|;ޛ��[��Q��6+2�ޭn���gz�s:U����R���m�ZD�g�+��C�s<a��5��H����-��}�b�_mݹ�Bz��V7�~�L�]�OZ�|�y�oW\�%n�Q�}�v�ٮ��/�F��&C1�\=}���٘jK2o�Ay݁k[�mïAD����v>�ñ���}�Ǧ[7	�|�O��K���{p�v��3��E��#h��h��Kݷ˲�=zKG��f�Ox+MǾ��_���n��BGx��.>^���I�]T�,܄�/����d���\�ݔ�T`x1�F���[�J^N>�,5ۣ��v�s~�q����N�ec��v�0Ob�~���o;����s��#�7��a��H��7�.v���Q�F$m9���=Q�}�A~ݹ�z�TˍG�|�Fy}74S҅x=����3_�zf�}��yo�k��y�v�<��_���C~�o5����0�{����b����Q����s��}��&���n���|�A|K�I����u�#�T�d;��%~eY짼����"io��ǅ� ���o]kF�1�y�5�m�vS�Ƭ�/,��<���r�u���sM�&j2�9O{=��✯g��V>�H��N"L�.��e�������|7�`�����=�F�W��B3�G7C��پ�VXq���Fv_�����ޛ��E+�������6釷j��������3�Ս�p�v����,?z�P;/,��l�����S���nT)��we><S�u։wELsS�^��o��k��g�y!���p���/��̯��.^>�����<�.y�zۑ�����MCb�}R��|�\����#E�l�#��xt�n2�$�VQJ�j9���#�^Nw���q�kp9H}��&՞��W�<*�^�1RVU���og�&�Ϟﷇ��iE4��w���}�k�*�{s���ϩ!#���=m� 5i%p~��ź�
y�mp�ez1���]�9�C#��1�tZ��q�����}��S����oo�Q�3�v�軰f=�PSG
9�yV��e+S�4S��7E�
\�ط�:����<�����3;����.��S�T��MG0;�y9�um����x�|�ƹ}�JI=|=��䦍���������4+�|x����W�F[��ó>-z��|ϋ��"������|;*�j�������	�W�'�dt�>�h���J<�I�+��}uy^�{Ł�돽����y��0���vuy���ǻ������}�6_Nz�өjv��;�6���un�О���;s��U�c�����w{Y�Z��Q��#ۦIc�xw��7��Uٗ�7A��y�W��ٓBϐ�|���Aí���/`z_]m	}�ANm��Ɏz��{V���q�}�a�����w��]�� ��$���i���6� ��Y����޾��-~���ͽ�u6z������<��������¢��֏������������_����������fu��qq��tZ%)��Y�]��z���������MG���~h��lNӣu���Kc;����ƤBm���� 3�S����z�/���`�0�9�!fv�P+s��a�m�x��ev��\�z��ลJ.e����ф�	H3�44HT3c��J�]x������-�-&���WS聝���r4r�����o1m���mKB�l��k���ɸ��<�>�Ώ�x�,3Te�6�`�Ks �s�͔����ur͍�k�tu�{$j�L8-�v!L�[T,����1��$(Ǚ�n����u��͞"�L�LCe�mi�s��9��0aU�&b�Y���G��M.Ŧ��u�XnnaM3L=�m�9R�b6�5��m�ڢ���ض�:;	�ږ�&�Uk+(mH�]-�q�V^�-�͡�TQLf5�.H!m��%�"*ۊ&��0�b�Rg��-���.�FѰv&���7Z��)u�,"�!�b3#"fع��2��Z����Kβ1�Em�ND���5\��Q5���gV��R�/,01� ��݊�@BT��� &N]VEXCP��%�X�F�k�8�f4�2iB���T@�Z��v$"A�mCYv�0�ƚV[G�ږ�4��b��RTFh���m�Z�7%,+e�ֺ��&n2��jU� ����fC��k]�qu�����Si�3C9yH)�8Vh;h Ri�bp�S�`��в�-��9f�%�;]�"5ʅ�Ж�m^M)��b\@D)������,�\��Mr�h+	�a��t�GCX4��/4+t(`V�K������ެy���Ka����H��L���d��"�����e�ʑc��
���n`[L�`�@0m�΄eèEp�-8�����pX�(̐�����Ա� bgK�-۝6kE�*�"�f��j��JS6�u�A!�n��X���mc-��1�\7+@��X�if�+�6m�*2��\��46��5V֓Ph�f#���vcD���K1�,
��8�9k1�q��ֲ��%��R�4��V�g��;2B��[�-���̷YnUm-��v���sI�ƶ��N-��c����SL�-��C]49R�WJ�!��ZkksKԪ�Q�o\�lқYG�)5E8���lq
hE\]m���]B� �/Yq����@�Vd�D!��:a�H�t-ekĭ��#w.ue�5��Vb6����4�#���lŏ
�����8]Z�H2��#kB��,`.�q�
5���]s���̣5tui���̺˳�4�%S&��3х�L@.�L$ccsbR�t���sD,`�.��a�նv���V�f^	��˨6W��6(M��b��m�x�ɶ�;i)5qST�h�6c������i\�
Eu��d[65@q��KZ��1bv���3�D(�jmI�sH��m)C9�¥�c��QD�2����`h�	j�&t�-k�m��b�`��MhۄCU��9Ub��. Fa�9^���*�j�[Mz���h�K2�c�3��%6�`��iu�vh)�R0��jA&��3X�ո��1�KBT3Ax�yF��ЙNk�q��113yI�� �ٰt5W]��Qj�,@t-��0�b i[�V�ҥU˘�К���[ �1]<�&h&q�i�n�h�]�i
��e����[	�4n�j�S5��l�CY�4����:5ae�b��tiB�3Qڄ�5�AYxKs$c�JsKB6Y]c2�F�b \��J$��i��;:� �4Z�a����S���5E�飙�.wh�����Eܘ�h�i($E�f�Z%��jc�@���{h�YI@�%Z0�1����x��J4�ԥbmyvf!pi�h�`�M��kV�+�:X�,ؐ���.F�\M-��4l�d���dqu`�X��ķ&Q�Keы	l,z���ͫ�ˡ��,�K�rj�֕m��ѕRT�avl�
9#L��.3�K6�\���X�)nHMX��ͥ�i��f�EM�Δx�b#��5jr��k͢w��39K-�ZʲZ�%�4��`����J�KMm�e�بL^m�Z[ufv��kG�S6j�ܺ���%̮��k�Vbܑ�eK����aF�4��M�@�[+��ƶ���a(Jh厰R�ű�d�0ı����#Ijm0!v�1n"W3$qNS��\�QM���kYFJÃ�lY�
M6 �DjL�3a�6��r&��f'A��g�0��[T�R�t�n�ׅ̦�s,�uU��j.*�2h��6��Rv�[�vv�A]u��0��b9���X���IAs�b3	R�v0�ѰѸ�&&��Ẓ�4Z�����.�Q���33�:B���S7 �pf[7���\<tָ�@�Ϊ��%�p�)reҵ�rX�$5�R5L��Ƣ$��-t2�8��Q��2�����iC��-�\�X�$�� ��.��X��LkE,���Ƃ�Ze�h�sW� �oa ���Hg[h^Z�[UqƱ�)^���.1GZ��u�[����*�he�l#,��с�aM5���գ��P�`����jJ+q�][�EXh8�`G`�iIs4T��嶯$�]Pe�.��^��R�H��0!��pԆX�$Ҋ����YP�zŌtve�C�X�8��NH���,x
�$1�f�n��]��SU��ĭ��j��@�C 9���rñ��e�΄�ᝍ&����7J��6�������D����g��0����ff.��LL\PA�0YZ2ʶY,[u�a��QC�+1�Ih�R���.��:�0,Ļ-v���5ZB���D������
��5�6�Bi\M��.���5��֝���K��iQ�h�Xi�NÖі!��X$t�Vj4����q�IL�k����6���v�X�aj]�6�2���Y�,�6����u6t�öf��U�2S��;���@i��\�V�����H����e�j�ٗ2�v/i���+�D(A�l\5�E���Z���v���A2Vm�5��h��"l�g�r/*f��K�V�ԁR���a����x����0Mr ��f�Jg0�搪�kb��f���L�T�[�H]6U�1`���M��]*D���u�G��un��9�uF&pm5��KKs�Y��)U-�Zz�EZ�j��̅s��fؕ�rA�"�J�m���-�SBݘY�6�!T�HimD�-�Uv�`���ἷGl���9ƺ[l2�1×M�%�heB�"�e�Q��n��WZ2V���ALH3t�j�3Q�5�[`И�l�&]rJQ��J8���GM[eFf!��fT��8l[��16�LM�,%ҏ1����J5ͨ]j���S)a��k%�`1��l�`�,�ni��#�p�jm6���[Z�!�r��2��qr�0Mw+`񦴬��)pSp�ctYICYJ�e�[nq��`�X��TڹKp�qb!�3[�4`.f�59H[6�l�C@3
���	])�ũw$W�/	��IL�H*.�p��0���MBi[2R�@@���ɳQ��I�1-ҚfKan��陪6��в�a���-`��.�#n��)�	Z�ͳ)H�6r�a������W���K��.M ݔv9���1��ų^�n����&��`�(�;7h�[6���
�4ͽ���.��l*:�����B���n���r�̰+%��a*X[s��t�du�%t�6j2�e��fW&����(�KI���AH�<J�f�[fu��)��y�NYrEP�����ݚP�(�m�cl�]Mp\Aa�L�5Em�q\؎�Gq��-ХZ�BX��b�V"��MM.
r��L��MG.�X�ku�������F���:�	��v%�e�b���fb��fB䱵�mpev�Tĸ�M���u�͖�HY��h����͸��0R��s
L��`��J��M��/6��+4n�ЋF���w5�n�.��*[�v������B]�V�L�Ji�.�VS�L]T��V�G1��9���p��abJ�F�j��C`�n���D���j�)5�%L!�FL��%�c�Mh�E�v&m�	�L�6.�iZ��L�MisZit�A,V��f\Ǖ�L�6.K�m���0�1nq^"k-Y�ˌ�< ��W3l�a��U �k6�l%Ơ3,*�J[nt!2e�#fve֕S32��'6&����)�QH��V
����]HF7�j�x���� b���ږe�Ɓ0��k�9���F����B�L!u
Lسm)����ˈ���U��e[f�*�C�����j�,�塭�u�ֽ��9-&mb�[�a�l]�bX��f&�vZm����[%Ѩ�"������ˆ��l�1ЌGm�[��:�ebŅw,I�Y��M�ڮm��.ԛ
�i�SZ*S5�ڍՅԦ����p��amVZEl�j�a@G(��9�ֱu��(e��]ᚲ��l����t�+k�YX�f�i��͙@S6˪�#:ܠ��֬\o�������r͊��t�RP��ˮi@Z��_|�kP��4P�ݴ1����jÊ���k;���C��o)����%::K�R�Ҋ����h�و������Yh�:څs[oUٍ�j�랔�̢��T�!�u�ʵ-:�,))fdCGH�.�є��Ȓ֍��Mm��K�Fyee�t���������N��Ò���>y�;]��q��X���zw�z���(ݥ�nM�a�L��uA�ືb�6���[�+D��\+e�,�3�ߛY�:f9�X�$��5M7.�U��=[I��Af����fn�j[��T%�L�����X�1ʵ������|1���}W��Eˈ�\݋��:���T�>�TK�^[F�S�mckӤL�X�53�R�lI��x `-�Alˊ[nڪ���`s��d��\���C
(b�rs����L+Ou��G�}-�V��L�S������{u����������]u�]u�]}u�u�]yy����+�����#1����IÖ��E�dU�p�+��33�����_^����������G]u�]u�_]g]u�^S��~�p��l�.A:md�>�zZa��*�Y�"8E��;���uݻ�܂��J�)K*)30��E��OD�"�����+š�L�G>I�˒e��j��%�(H��R���(�ry���dQF�r�Y!�08���
��QW>�"�t��H�*�͒}��#�EhU�AATr�*(��p�Nq)�MPDZ�;J
LI)4������DDQZ��h��ҫ�f�hW(��U,ƄǟΔޡUn��������QVn������s/�'=Ӗ��RE��qw!/�7s��z;�+��3-�Q�t��q��5���I1�T��Y��/z_Hf��_>W�ߎ���RR��͚�GX�,��:�[7�u�����[LF�d��Ӫ15ct�K�ŨaW]B�r�2�x���X�-�WK�+1Q%!�ۈ��25΂�,4ѭ�FWF�m��	�mЙ�i��h�C��iY�"ݮ��5�t��UΪ��]�i���)r�]cu�L�[<s�F�غ�f�c`M�t�ض%\֐��f��rhԖ:��K��9��Ti�[L$]�ʺl�T��t��pYI�#�%#�������.�oj)Y���-(V�oݍUj6���XIvaEӧn�)J�Վ��i�%��j�!5�]�ոB@
*J��rىe+\�c����V�+s���I���y�V�btF�����7D#�.�=�!���b�ɱ*̻�i�j�[j,e�8%CT)b���tt/8���ֶ�阑��t��t�D�a�j]5�l6��k��踶�R��.���W�`P!p�M3Ycr���]+������Q����L�pi�쁝�[����X�c�%T�(����fk�v5%�Jh�fR:"&�]cfa�*���a�a�)h����M4l+gp��4�F5����ac�CLr]H�*]Z88�Ң��\hTw4I[vK� ]��++=e�X]"钬h��"be�n�ZPZVK�+6�Yu�c�j��	Mtm�Ɨh�C�Y��ZY��E��a�WYGL��V8]�l�nb�.�0)Bɮ��ֲ�C!6K

�6:��+0�!6�f:
kt�xJU6�Ҥ IE��M4��dlefЮ��Mv��� kʱQx�cfbT,[s�4��І�<�h&ʙ3�|����WM^p�fv�L���Z䙢%�>ye�d[,ռ]���vZ�\��$ٙ�it��cB;PIl����]+Ķ����o4�޼�7�5�������F�4���Cj��tT0]2<ؤmUk.��;�7GGSE������I��8�'N��x�k���K	wF�Px��V<
�<��B��u����\�r�7/$ȳ��2��e��e,jڶB��4V�#@�j�����Y[Z��PIW�m���{�1�����"s���)"5+��,�2ե��$@��ʃ^Z����6�i.�yH��%�P[(�,�el؊�
�6	����
�
��ZR}�B���L�d��!�	d����ca�VB�)���m�L���<(˘5���[���~��t�� @��w[�I&f�G���5vB�Ƣ��
�P�q��g�_Ί2\�w��L2��nPK��q*��D�^�KM1>��>�F�� ��)�+<�$U�V��M�	SY2A)�g�D�I9���Ѫ���4j$
e7~���$C��Bt���LD�dX �75�݈w���y��Ng�����I ��]�O����o�g��^�'�,�j�\KsJ��c0icm\UR�@���_'�;��6�|j���}��ngY"_"�@$����N�K������'��_L�}�dS��@,@&)??˰��*�o0�����qv!��¾���{��yB	����]����}���C%�?b.�{����6ϩ�Y+R	�������b��{עQ$�v���� ��x6���[��;���+��M���p4^e� M�<�7��@5��Yzw<5���}��h H�^�+Ð�C�%!Vתo���I��� �u��q���Q���{��ǀ}l�0c��;4�6e��� �
���3�xpز �F&I4�ΑD�z�1��g�fT<Ʌ��n����x.�;@��e���%��.� :���6c6Bi�Hm�:�߻K�a
m����5��"�y �A�vF��;�t��ȰK݈avJv��0���L�j��v���"2E82D�x$d��,Rw�F�Z�M��c��kZ�b@%��\ͷ�xبI����O�~��l�I�Ct�	<�?79f:�w�-~;����֒޻V������6�nr�4��޼�����l!����+�-AN�<	b�vZg,��0�/4�<�%m��,�}����!��H�H��LH$�}�(�/]T[�Lwi��,D>��A�<"D�[ I��������h��VQ$�K� �����>��B��sM����
6�
I'��D4qeX���n��ػ��&]ζf0sYr�=�l�|�U�AL%�?�恠��nD�I݇�'P�߽6�
s3���~H#Yh9Z�Ē�ed���zA���N�Q"K�>�E�U��wDҜq����|�v�׮�X�V��<O��q`�$����g�4*�n� �C"m��� �yěU{����!;۰�B�ِX���I��x8p一��O����/d{}e���q�A:�ٍ4�L���U��8��.P���UnR�M}���t"�ˎ��Ǟ�j׾�3i������X�	LC*�V��4�ۉ�f�̄bŎ�S4� I��nA.L:�C���{y2	d/]��4#�6Q$ݒZ��Zh���e���׶/!D��#}�F���uI�(RfSF��m���
՚i��8�f�WQ�Վ��ǵ+�ߖ����t�EL�$����$�xb1//y��"�(�	��̂[`ؓ�`DD�o�	 �����S���$k\\�I#�۰"@#$�ST@��%�˒`���TD4�S��Ȗ�׀A&�'���L�f(���%��ׂ���N<H1�'!5Q/�^�E�n&oޛڒCZ�,�,�;f�	b�s�I���n�Cl>�/[�p��q��<c$ı}͐&e+ǳu1�%i$�%[� H*se�*d䒴P��Y���\�Ǆ>�N���/v�g�廒�wz.��#�Ӧoy{P���2/������^"|���3�r��B�\c�4t����z�	C�H[��[�V��b�PvwT<�,tS�RR[�A�n��L��+^�v-ڤ4�`C�lID5��kRb飬&�xۨ��
*�z�|�ԙ��pf%���
M�Kc��q��2��!��m��.�B˦�����"S`��&�4f��%�B�Ku�h�!�sh�r�D�fGL�[6A�J\�2������m/#�U��.�X+s�3+rl�����PB�m*�Q����&�s+��<$�r��s9.�7��z��{���`ui7��~j�H���Fq!>��:̃�DL�""����e���\]��ce�@���vI�nS�n�o�^Ƨ$ �K��X�%2�����s\P|$�8�˪�D�-��̊4Fc��n)��� ﻃ\� ���ZR���Sv6.���wNz��,E�^	$�͙5�;'ħ�Q\��S~��\�����0 |w������Z}D��2��`�S�9��VhE���]�L�<��c��^ڿx;�%pu�[�ě|�iy��?��>~c�7�wk�x�&�(�إ@�*�e�u�ʎv�X�t-��"f��6JC��}�8q�_�2d�Y�z�`/�~�.#F�_��#��A����X��nȰ�{߰A��2�^禵0?����!�ǩsB�մ�>�:��e��D�2=�S�r}��"����X���t� �C\W��J�E�Q�U�������ANo���TӺ�a�1�;Kh��Q9�lN"/ޠ��b��Sy���l"ă;��>fT���� �$�� �զ/�$`A�x�TV����e~yi>�l��$���E��A͇�|Y79�W"��q]�В��D��BtJ��qg� �l���2�M{s[%>�ƪ$�'�a�2Hn�<ꗅ�N{���SǄ"���eƗF�l���-��3�Ҁ�6��.u|��q�[��wz	Vp�'1\ X�dw^�畍���_.�33la���|0�	|ڼ&p�"ZUƼ�Izܷ���xkɍ+� H%��=��@�׀ĝ����z��fo�)w� -cC��j`.X�n�H"o���jӹv�S���o���"����%��C|���+^�佀<:H��{D�7��H��}��)��ĵ���r4��|/�|��0#���w��\�y	=�ϵk�\�<�Ti�K&Z�uL ���&[x�����־@��#<��}��k�0f?�F\('�lL��X���6����@z��Ti��%��8�X�ݑ&�3���u��Ӻ�ASf�4�ƈ7D-�ۈB˦�͊Qyp�v�74���ﯞ�\��W�(�(�[��~�O����+sfA�^//�>'�.-�I?��n��8�2I[�/ߜ�ힼ!�^��2gp7%�[�- �A�S�)���"�9H�!�
A�ǀ	���,H{n��^�a��&3 EX�ݙ2=���$:�!�w@~f~��؟捭s�@I��������9HmK׮=��13[fn3�s�b�R�}���X*,�VJ�&N����B�ջ�#l��9s�c�b�3�1b�X�w��	�\�����e�l�$oU�� �����&7<ek}.5������;���O�Ly'���u�}��٦��cb$�3y��C$I)�ԷLk<+����g�j;O�Ru�h;_9��+�����3	����!(�72D�/��n�Md!"I�0����b��y$��T]��08�wı2���N���%"22,C#թ��b��0\BI��愲���$��D��J��N�S���I�n������� �ȵ�������kӗ�fЖ��A��X�`�2G7]z�^���A|��$����������� f���_*Gs٠����N]dK���ܖ`su��x�Q�;��Ml�za���׭?{Ʒ�7���v�|d��B��������Ŗ1�!��Ǌ��G���?�]�}w�8��}��d�m\�+�UF�,���73[Xa4��1�N���f�)
�RZj�6�\��VKF�sc�!s�:b-f,��KtM�ᶨˊ�KW0����1�p:�qG�M4b&q���� ���-�Y�A�6iW7]3�u�0F�^�"�K���u�p��2���ە��ֆ��*5%��s]s�X�%�,�T�u�~�|��y@M
�Ύ��p%�M�Ȁ��	n��2��
��4Wy�o�d-S��E7Ű��:oy�D�H��� ��p����ǪMX7��)����$dR�0'1x��Eo�,]�Nk�����>�l@�6�
�I-���ךd��[f�/G��h	'��y<�Z�>_����O��� B��IzLE�g����=���׃�:�&[�@.�~��h� #��u�$�-�y$�b�}�6i^�<&��ц$�^r�r\C# }x8��y>j�/쪒�b���`v��@�|����vn�vu:�=�s�]�(G]3Y�a�$����h�Ƣ����|>�}�����!�<��@�d/1��|ہ�'�e�Ƹ�&� ��ǂex�c_���I$P>��$"Y`ӎ�8<�L�_�+�װ���h�<���1�5�K�6�e�u���ݾ�D[̫P*��/":#��,X���t"H$��� y�T*MEG��}!L���<A�����"�2I��-�5ꨩ>`I&�]����Zc}E�`'	Dhƭ|ȵsĂ7|�<�&$=�ȟ�b��ݠ=_�� �s�j��xAM%>�/zA��s���޼l���$}xc��%�.dEc�qV!��������=;յC;l̰�s�%�%E�3i4�딶2�+m�������ߴ�[Y�x�AO�I%g�$�µ �N�:6dA�ֲ}��� ��˘H���h��C"^�<}�w ��?�%��o2|�~�￉v������*����y�7>s��(��|��I�?�`��X-�������Pַ���GB�{noTY<�n=���c'�x����uY��{��J�n������>y0�^���}�v�c��wt��^�w��P�:�̳Ź3�=qJ��y��)]k=[�t���"q��ޗ<���{����n{�����I*#=�d�1��,"�:/e�u�v�o��7+�"I۬ʯ��n5�,���>�)���s7��i��tP�ɽe�|�zh��a^;��dg0�/���{y���ˌҨ+��S��(c0r~[׶�t}\���(����]�9�s@F���|75a�^>�U7]�b�I�wuq���މz��A]�T�ދq�tt{ϼ��뻐LUڧ��ޒT1�jg�Uv�co�ts��VQ����h{��b��k,�����^���SGn��~>38{��Kɺ�!H��&RL��:n.~�z�N�Y=�֎z���e#T����z%ƲS�?W�U�M3��{�ל�;v���Ÿ�{ۇa�_r���&��{�Wv��f�.��9�9�.-Z�TZ��ѕ��gM�;����[��.O���=��'�������z(��ysr��N��#m�.C�����d{=�猫�Fj�(�ՒL<��ܔy�ˤ�����O���~^8^x��任�C����bf��= Ll�RL (~���X� �g�Fo�-��h�z�OKyI��K>͛���G��)b���EDe�Dyk�%�횑��LK����]���RP_�a$��p53�T�擎�l��uޞ�6�yU�v��A�[VF*R^���b{�8��x�;
�q��9���{��3��_^��|q�������~�]u�u�]u�_]u�^{3�@A^�mC#[fE�x4�)�ܸ!YD�J�n�q��c �$0ڧ��y���KJ�NŦWK5#ݻ����Ǘ׷�_____���������]u���]u��lva��YM�@s9������	j"�6ܰM�2�+]�:�f���ިSZU�&qL�oX��s�v����j�R�ă�n��t*��9�� ��S�H̢K��P�'��N��Z��싑�m$��ѽ�J����a� ��D9��sY$��H�t�*�}�sȜ\9*X��xpvT9	S��x��B�%��B��=A��u��H�y��d`pt֥����E� ��q©�D�{��GƏ#�z�򢫆i�W%��uܢ�r&^&!��&�z�IQQy��� ���8%�$:��V���T��!��%r�Gw�܊/"Ά��r�A�*�䅏�p��IfUl�P.F�XuRʸt���QV>\�ք���Q�����,'�Ur�f�}v9��+��Qi"Q����C~��ѭkk���{g;�3&,�9ڣ����w�o�a~�'�����r(��r� �aDx�����<�a7�5�� E�"���Y�C# 鸇�3��w��z	2���@Y�e�������r�z40�f��,,�lM��CٓH�0���go�q������؂�c��H`�i����� Y�,�C�����c�}�t����OC����fD �: ��!�a�/��}>N|S��-Z7��\�e�mm��5����Z�)XE�źj`�Mz�H����Ϭr�A��G���C#�}��d�\�%�������s��8$���������0-i��zg����К�@aT���bd??����������鋧�2B�"�t�A��51 "���1��E�	��FǽX�o)�nd��C��9Rd9?Lv�f�,�n �@D �"�eǥ︋ I� �E³�܃�B�!�������^v*؊0��?���LL!�!�������`�F�m8����Ɛ�;HC��������|p�b��h��:D9�R�`H�t�d+6N_e.�fY��P�w8!'m	&+�������LC;$7�0�`���~�j=�c�t=�'49��廡R<?A����/�.k�u��K��/|�g�'�uc���MǜkQh *�a�FA����2d��όc)JW�yϼ�K�D�vq��y>S9qU��t���BH��o��$DY�]��Y��Y�U��8o#  ?u����J�� ���3�Ϝ�u
���_3������|�`��V�vi�ݭ4#[9���l�7c
!eY�t�����>��WI�d�X>��dY�$�A��^��a4����'�����c�}Ӻ�3.y�ͥ��ب�Y�� H��y,$Ȱ@FZ�8xx�RxN�Ø�e�"g�Q Qf@fK�OP������\y�ǳĆFHa	���%�IE�D���0i,��`Mu�S�����2#K �[�y���}�&/����؁:$'i;�����0��	`�2�"�xus�[��o�����>bq�.�׼u/Pf��,�9;�27�,?�I�����,����د
��]�|m!��;����~"�2bH�`
A>wK�)� � �p�t�Dw��39�tq�x�@�CL��f��np{r䨇0��G�}( �̈� @E�c�4�r�a�Ѷ9��$=#!8��a:��:lHgHE�C�L��� 3����0$WE���q]A�j���蕛��X}�1�� O`���ā}Ow���>Bߑx�u�G�E�vp�Y7������9�jyJ*0z�?���ť�dɿ������XhSWj�l�i�d���	h��3j�´v�ٴ!�aa
˛����� �i3WL��0�ְіʃ4\H3^ml]��5ev](g\�)�s�����Li�K�͔q��bWhpJ�dV��)�4K-�Y�V5%ҹ�!����]��8�=R�fmi0k`��gR; ��E�ј�5��B�$l�l;Z���e�ؚ��(6).�y9�_{�-�B�V��1�<�i�eRj˕���3�vJE� �E�\R�]�s�ȼ<C�C#� OwZB�Bɉ;�����;}B?Zۜ�����X"1���.�ą��|��s�~s̽d����!�ds�d (�!��9���0�p�ļ��a�Q`�~�ȳ	I�f+����"1^�����w�;����#��K2 "̈˭�/'0s���d�<ʝ<'S��__o�L�sv�Q>��&G=}w�w'p��]�ѐ�Y�1mb�P��8!�s��+ö_mO;�>-�Af�Y����'o��
W�I�:�듡�;d20=�qV��8�T�")��ˈ�-�i�W�~N����=%���m�����{��{��1�$��<����!�`�dҘ9�Di^���zSXaD��Dgn�a$0�^�ud!���_|�����=�9)јd���9�[d�;���K� �lXB��K6�~��!�G���x��'	��$��� ��!�`��.^�x6���� ��m4��mc6P.�5(F�t���t2	s�n�vy�m��B�5�ٹ>�[�?XSߝy�vI�&d�A�l���rC�NI�g7~~~�y̛��a�߮���l�,��TO@aT�1(��_N@��Y�"�ٶ��P��TD/P,�d �� �ZH;��t���B���MiЄ�A�y��z.~I︭���Q�z���oyL���M�Yg��禱��Q1U�S��M��&L�4����o���LN$ӣ��ߟ/�T��(���զ�um�A�����a����F�P '	<EL���I'��	6��RC{<�����[$�S��z�wva�wt���JX�5j�����ꁴLGt������X�$[)�$D��^�x�PI��C5��
�3����o����U���N%�/2]�fY�Ҏ��
�qy�ʋ�G���I�Rޗ�DDPwI{m�U2p��Ʃ<�#����s^[q� A.TD�E�Ne+*�1��6eꖐ�Ò9�e��?/���\d7�t)���'�2�I$7��d�Tћ\k�)�jY�u�ӌ�M���9�K�Ҹ�W���?��J!t`���A�;є��/{r^�g�լӴ� �8	�I���]�;��wvS<d�/:�oz���&�G{!ZHM�!��<;���I��RA${��eZ�8I��7m�l���ΣU���鏼�&�j��zk��W�^�����j羯)�3g�����Q�P"���K��Bn���&M��co�%XI$�[�y�RE���T��W��*'��<K�/h��o���K��=�M)�O�ئ�)�г{���b&u�5�h.NԼ��ݻ۫PǅO	�F]�2��I��Y��{!�nLw�-����w�{���K��uSә!��S$���`���֟9�]Jbb����lm��u����5���ۊ��\Śk�/D���pI�)�2��KяR,�����I)�::�%S�^pu`��l��us�P�($�&�-])4X�o�@I��yt)�gI�P��c�<�'�j'b�JA"K �r�d�K�t)(���f�|��S�if�V�	Y����.RxJI$��T��`�䀯��eK<��r6�7�y��I/FNC*�)%���OL�i����9Q��|KߟV�=��nM��y��IO�=r=I&�/ҥ�I�ϗ�����{x{xH��k�X<�Y��zI�A�b�ٹ�ɳA[y.,����z
��<C1���ރy+nۗ*�A#�'A+��q��643�gggfa��~HͿ�I�·�y/�@NxR�޲ڦe�H����*��K��Z��,wb471�e���j�P��Q��.�L�)osȐ�pM��d��m��fb���L�����]Hĥ�ki���4�P(�Y�lG�~'��2Ͽ?Ox�v���~s�GH%ܦ$:I �eݯ$�~G��*��T 
d�s��	!^U����K*T�F��A!�z�A���M���PΉgo�q/) �=�)#c�1w���	 �kT�ٗ�9 �}���H��޽N�qR��57і3rp�Iu�ʑ��$��᥊vz���r�;�P�E�{=�<���U�>3/�H򜚄I'�^%�A w��g$�%yо	&���L$���<�E�l�n��H���H�:�_�d���a����y�!"P���d�;d�zD��w��Q�
[��sϐ]�f]�:�ԥ�W�V,���U�;��	�d���|^%7�<Q�x�/Zt/U�{�O��@;'��\�D�n-,�᝝�  ��>���^-�λi�Fh�g#`f��Z�18C\gqM1̴v7-��c��3�c�1�qO��	�Y[�F/�:s)����jc)3�]���.Q��K\1ؖ���z��՚�*5Ļ��v��#cٳ�w3j�`ؙ��c3k�
ʐv�M��鱃 `�mvѣ���m,(] ���fК�d��sM�"(JG1Ce��p�;���{߿<h�#KY�
���]�Rv))0��p�s�͛tqh�=w��eY�]�`�Zi��<Di�v�~�l��_9�R	$���q�G��ڃ+������(��p��d/�w�,��j�}ث/���t�>~�)��+�`�Igs��ftd����$���%�=B�w�����X)�)Ĳ�M���R�A*�̧�S"��(OP-�x4��t+J*�x$�]ܪ�g�6��x3à�]�.�S�W��ﭰ6�	$�]���L����	"ȡ��+3�_��W���wu�o0���'<Z�,"pB�[ʏ���is]�k ��sa��H*�yBI���q��"�Cu�T�+o�]멨���?=��<�V�c4Y�da0�E��Y�Z5�v��
O3�	�ϛ�?vL��߳��K~���m�6�= �dR�ҥ+�ċ��q��}���f�� T��	���@/x�5�O.�ƇvI�L?fp������`&��a�8{J��K52����7޽����|�C<0�jݓ��ۛ�����)G������p2G�|Z��������3�K�� �#���d�M�?ҥ�As=nB���͞yx4&|{��1
/
Eݥ���� �,蔓ُ��O�SG(x��.kh����A�"��Y���;��"�C)[$��1��{�4Q��yM2I%��*RA$�okם;�s=Gc7��W1t��*�2���
g�A!�x~J�C�I=��%Yح-
 v�ͳ��9�M�3���]o��$�3�绞ZV5��Y��	;�W�9z���xЋ�:���"\�"��B�ZL�ɺ�V�A
Bq4'F!�\�N���Y���J	_.-�L�$w��BT�G���j�p2.lo*��+-�T�d�gR��Q�W�跙E�&��e��c����m�t�Hv��&BI.��4�A ��܋�n�xW��2���P��=%QJp��4���$�!Wl�I �2K���U��}�?g��?�6��	˴���x� �:.��s��{�Y����ީ���G�?�����ٮ��Q�e�߽�S:~Ƴ��~�>�ק�N���EN�3�3��@gp���V��_}/}<U������%����n�_[�7a/R�FRL�2�c�I�]��N۾z���̀ZNՑ�T��b�$�"�C,j%/-�N��OS�������#k1��i�'��R�;�	^�̢I�~�B�λ����u�����߳��\�)t�"�6�F���Gm���fsU4&�&�`SbƧ�0���~������u��BF�� <�+[�/ʩ)�W0 E��K��*Y$�K��,%!z�V��w��T�n�ꧤ����O��P�c^]�$@8��M�ISmMr���pT����(��.@0+��Ar�!Rʵ-�y����+���I1*�
^O����`g�t/$�D�c� JH�ŕ5$:r����'����#nVp��Xod�/�e$���)�@$C9�R:n��M�u2�`�
���p���/�Fzw\_=���m���oS����ܘ6�vޡml_�fD$̢�a���
��VD%���-L� g��ᙘ0vg�"f��JB,��x<C�%�C��	sd���d���ĺ�����+-=���,��y�z&�$�Fڒh$�z$��7�vL�:��S�P���D't]u��m�� bՔh�]p�A��a�V]v;{���g:)�8N9��~J#a�Y$�&Ka�( ��	 ���'���̅��b�$��"QA$-��T)z����S<:
�-�������L�e���W�7�2{��H���A���I �n� �I2]�~���\cԵ��e�R�rX���!R=���l=�W��,����ٝs���N�i$�.��T)��e%Ԃ؀��P�=䟭�Yu
�-�ì��"j^{��
a��٣@$�s;��F��K�E���u��no-V��7��)<������i��u���z ���u�w�������/H �ǲג%̈��%�w��N8f oz�q��袵���c����{��N��ǋ����xq��l� xQ�A�VF�c�4��L	��ND%��3�[p�����K�4�H��� �d>=��پ�y��緰{uɐ�/�����;����ww�L��e��=/bX`,�)���zgE�`回��ɀz��6?m{�EI-����݋=)�����x�M��}�5�iSӆ$��S3�-8=���ۃ�Wj3;����̬�ᅾנ	˳���F��͊[��}N�|���n���Y��N�p1���d��;��F?{oM7|Y�D��A����3^=��L�@���;ko����8M6�^�k�G�V�"��{qȅ|���c%��=�n?1�Gl)FIc�Ůz�S����x�~���y����7g�����H���X<6y�g��h�ocx[9�0?v%�_-�ө�g�S�y�R�����O����[��轨z�g�y��[P����>�'��д�Gn�	�@�����@ߵ}=/_p�Ā��݅�r�9�ù%���ny�����b����t1HnyzM�=�E�<
�:���cĦq.K=�����¹漷Zc����1�D��x�� מ�C6�=����<O���׮nYKc��㢬�A��x~���Y��Ca��%�J}�9e��r+�{�����x:4���P���{�ӤB��S$�)Z�"��)N�DB`�'Ė;X�[((ȅ���H$Y�8�0�S��=�!k���קˤǞ8�|�/�?y��-��}�����������K��J"��Ef�'PQi�2TCE�����)Z�o�<�N����lkkd��������lmmd�����������XL��E�B*
9i�9%�V(�$\�S�s��_��ʝE�
u*���g��7�w�}߽�x}}}}~?�u�u�����~>�����������p�L�G+�"�,�ei"�R#	*5(�G�W�f}� ��w3 Y���\�"*��C��HlT*"+�d��*�$���w&���#��;Љ �1�Vd�s�� �B�.I��UA���:d��j&t*���E�+�]��$$�AU����Ȫ�(��ʦ;( ��pفd�IQ�3��J(�2���*s39R�M2d�v���p�w$��z"IW8d���$U	�!�*�YeEE�*�XMd*�AD֢�y�k$¨(������(jFaȄ����;�A^l�%��!2, �!A8kv��Y��l����Ǟ�.��3f��Q
��Q�5�)����d�f�f����sSV�V�c4x ��ԍe+�����M�(hYuƔH��tփ��ڳh���6�`΂���K�[ɒaK5i
SV*$��Ԇ����+��ы��g�,e��aK�,m��T4J����Ǫ@�L�����^��ֆ�f�̳ ��1MbjB�5����ᶜ0j�j�ll�SG�%3���cv��iD�%��UJd�:RA�2��u1��q#(6�	f[t�:X$��э��ٰi�]�b&��%��l��`���&ͻ1�Y��e� GWu�2b�������hj�P�fDJ�n˂%Tƍf�	m.V�̖ƼSbE����͢T&�s�F�tz[G����e��]y�4꺔:�+�J�X�Rc-��eց��Z�]]*\�[.�I^��1P�f��l֮ٛ9b��WB�hAM��,�\�������k5̳d�����h�,\�K�s�8��!�*Ԣ����r�g�hh��Fbf�.��kX
CM .Й"p�XB�F]L��;�t.���bVR���]c��6&+�� ����U�.�V�t��蹙F\5������R��3p86�@%��&�.��ڢ���xJ1���2�Z�p�;�LK��-MQ�]Ih�ZUY��:��-�7��ҷ"Y��.��-��S-�Q�F��Q�� ���,�@`�5wd�Jh��̬r�7G���&��ذ����ʷLP6phE�F:�l���#`����W p���#,УJg�YH�����ث+��iSc76cc5�P�iZ��^m�h�l �b�KJ��:�p�ڌ���6���f����IR](�-�����`��"��Q��؛R<���6��Zصn�.��`hF��y�����X�z�f�:��J��Bhe�lĺ��KD�%�k��b9\lJ˙tIR�,ؠgxy�Kh�ԫfn��T��U�2�;KP��)��hV���I���;t�/n;v���H��������ԫ��6�5��q��2f�"�X��[c�nG0a�쌹���e�J)u�D�m�k���V+h�ڤ�k5LV]�=�t�a�Mڙ�]q���X�\ �	�7�ư
����uمu�s���*.F��4e�\c��k��T�k�
ZV�:��bUԖ�M��ۯZ\ #dl�X�v���<�+.q���s��}��bӸ�W+�l͕�q���"R�
$��Mr\�z����������?|�����/��zA"wq�BI�&7ȢTs�י%[Z�<�~a��)��1j����(����1�wp��C*�K\���]=s���t�hc*^}礒d��ȓ)$��ݯR�>�z}4�t*�3��z6"	L��/{ˢ^I��%���)$�[�<}yN��m�Ԭ��@!��!"PK�_�Uf���"��� :�hF��}�..�:��ȩ��k�,�-�L"��^Gy�BH$����� �Y=)���$5��S�/�z�qAr��x{� �-���H%�Q����z��'M�6��sz��RH$�i�z�$$4�u+I�w/ϼW���<�Bl�x�s�6B�h��B�M!
�u&Q.f�������uf���o�}<ߒӀ�����%'U2Y�Ux���f��R���t�׃&4�7��<
G��O�OG�������{?l�`����K��/�pz�����ܾ�<�u��j�&f�~�ΪՋf����O��Ã�y^w��=���C��g�¨c�<<3�s;4W�G��H��q�BG�IC��^d����O]�KCe�°�HK/�?OR��p���]z ?gߝǻm�
$�_o�
�����V� �eNs�xi(��ɍ�&����0�Ja�)ioy�Zy�R/3kn��H2F��-)�@'k/ئ�I��]}r�?�]���I�����Vx�Z.��"�r�x�g���}��uu��9�!��p�02���hwT��BI#����/y PE��D՝�����l�EU�I�$�.�%�@NL:%F�]�Ay�֓kYv��U�چ]<��0�K���զ� �t��h��gl�ǙPt�ɸ�T�E�o,�A ��zEs�g��!)�y�.�e��&���j���a�QG�t#a+����x5��_Җ���K�g�RD���zgH$�kؽ%�=0-���d���oxxr^=Q)�7�6���gI-��.�D�k$�1tz�cdl?��<<F{L@���kX�hY���zɜ;<�����M;�8>{����W���]w�ۓ:̏�@�ygǄǆxxQE���Q� �^���D�d�2m����7��@��p�!�*N��������I?�J��&Ih��D�H�c��D6k�[�cd�fs	t�FQ�wAUP`��>d�.Pa�z���O�)P��k��y$���(�H��Zҳd�i�6:��������oFmtzƈX�kUZ��V]eb*R`v���aS0vaז��탣���tUVm��gLx�k/�v���L���2�39g'w��i���uw�8hR)"�ϰ�$�';��;�
���N<�CY�u�;�ޘ8=d�|f��r��$�,�)@�{��	E���YOPK���}��W��ZSL����G�#�����^�x4�d����|x���̒ngw�}�L��-�y�H�z����xJ\��T�E��q׾S��ԉ�ǨB)[:Y�@$�ǧ��T��|��y��H�v1J�V�n'�Y�\=�ӕ7���A5�����+?��S�Ƴ���Z�KW=��p��y��3ú�緾u�ڪ}��ǁTǆxx�9 �$�.�s;�?u��Ä�8��	zu��]�A/�єʬe��Nv��f�$�,�r�
%2^�x)��I����%�ћ�6Mn��Cz������t�Q ��#*���X����h�����ہH�M	�M���v�xD�Q��BR) �ȅ��$�d�F��5��.�^	=�lƤ���"SK���}o
L�puyww�9=qj��|*����f�9���I.gv���p(
I$z:3{Ȫgz�2o�Pj�؋]�Ev9A�ćt��y�%oʃ��Y=d�nz4{��Ҭ��DPI$�"��&Y ~��Krw�v����&��qg�����1ß�|F�À$�G:�Ky�8II��-@J;�1D:Uꗸ�iE�%���п������U3��<Ė@���!I�umǬ75�$�L�ȷwT��	1��Á�ˠ΁3IX��K�,g&`�t�j�r��+z�ZR��S��r�=��׽��o�2�����s��E7��^�R�r"���z`Ib>  �o�~� ��T��:ȹ�9��2�E��[�5�����(8�D�7X`VU���;vD�\�&屻���tj8�[�BF�*�]�f��,F�w5��;)m70�c�/�P�<�9S-iX�	�XV���6�cD�m�RP��%�]w^Y�k6`��*�&onLK/n�P��ۜR�mJ�n!iїM�X$:˴ �8��X�5�]�&YAYv�iͲ��p��s���ߗ��_{�)86kk`��gl.��̶m-�3�h���g����� .��툱��w$?���� �2��Α.��DJO�o�eי�iOc̢�/~� I��y��
!�v����TȔ�޺oyN�&�k�$��$�	>��I%�=�1A�IC<�|ٖ��~����
��Ӹx.�z	���ڱ�HvLL�A*Nt�����n��Ef<��$� ��:@�jwL�7�$%�^��q/�1"Zg�p�1�GV"����ؘ%��o���   orbBD���������H�Tq�I;ܓ� ���Θ�ғ$�G��q�;�=ySV�N�/�V�Ѫ	 �ٳN�	$����+��)�
��7��6���>�/]d��5 �\Ri�]f�i�����aukT	PV{���K΃���!B&!B���S3J�(�2�&R	 �$�<�^վfnx��4
f��5"�I����w(;�!�u��h��2�^���"�K��Up�0�.I�3A�_�}��/s�=��asv8���;ou[�o��7o{�#�<����M|F~>�s|��}�p<�%Ϸ7��]�5��,�T�Y3ڐ�W*��{~Ƴ�p����c�wi���?�yg��@ǆxx0|ny����i�If�JI$��w��D
	b��Wώ�t3�^ȓ����0��PC�c]��ꙔJ	�y��w{g��n��c��>���854=���I��&�h8r@���S���Ok�Ᵹ�������7���n 	����3�u�u�S;�@(�����Ǹxd���4Z�Bw�ۯ�Vw��)�b�q���~[�&BO}J�նt�z���>�{�E�[�L�M�L��4)��{��u�������vpXld���92�m��������nvX���-�O+�*��������]��E̖�JH����Hs;����D�*�y��͗���bB �3��k̤'9�V""b)�n�*���D�ˮٵK6f����ʌ�g]_k�ӻ�����4�K��\����y�6��T�1���ւ�ĩ�u�I���t |�;;8	���[U��V��S���������`���y���ޘ�&$.wt�r�wÈةZG�}��*6�+׈\E��ϞU�Ʌ���μ
<3��#E�fo4g�0@8�	wk̢�/�G�U������2�5~��%oZ��4�,$����=J%2H?�p��^�w�\�@�(f/(��ٯJ$�c�JR�`���(���~'��n�$�Ć=�)?����[�L$���%2H$US�*�HgtD��Y�����(EU�޽�4�2�IlT٣\�w:�20�Mp����Pxg�B��[T1î$;�h��o2�%��4�%��w�bBH_ue�����)VKȕ��:J#ӆ�$6č��"	�!Cĉ�t�ȝgvuq�
t�w�!Xl%U�	I�I!��Y�$�=�1!$��s�)�y�%#4oYzD�(^�$�1���̑#;"ZRel�]쩍9ƞ�k{=/4�)�m/�1�|��/3	#��hK�B/�M'��[Z�䄹���A*銠�gr^�����%���g'����s3�$�BK�(7V�a�^�ΊyM����{��В�FxJ;��ǳ���Ҕ���ϧמsx-9z�VN	��DD�㖲=������,�����/�9}���ξ^�s�����m��Ϟ�ѿz���~>��+��k��nQ�UA$���.L��%��עzs%W�SF�
��wޗj�e��nk�4�9���Mm�3Y��qSe��z�H����	w)��u�L[Ʃ-�$��Ĉ&I������x%ݫ3O���9-f����I��!�$�+�8ud�t��׃w
_Ӟ8);��y>���,Xg�$5v��H$���h��E{�t�MA��B,l6%���$+zx��I����z� |��렄����f=�m=��I;$��eɐ�;��K�i�2A��P��$z:��}�#Z��RJ��� (��wt���L��޺�'�F��Ha$<��ɐz�x��.Ru�RO��I���UMgx�qC3��k1tC����%���L���ꊤw3�e�{�!�>�a񫨬�����rOS`Ѫ�|`ť�e�!3��=��]�|�s���xa��4t^��ӽ��]s�՛��]g1}��Ol�� c�/<����~��<.�``��P�kv��R�]4�:R�3Va���hR��E1q��F�;:<���F�tD���j%ˈ�4E�����c
�1qZ���Y����4f5�	��Z��z�
�]��"fk`�X�YF�b3Vf9�j:�\����l8i�\X�W�M��bj+�Lj�is�[	5Ih,�!��q��5�^�n��4����va�w��߇��}�ՠ\�`ԥ�%��[k4+Z1���F�6���i1�]��	��g��6����jߩ���B<��Gr^XJI$��TsW�]�^�#:0�U�&1� � ��z�7:_?!��Z�W	����������:y�1�Tbh�w>	$�_�9;̰\�;�I��$d��7n�k��χ����$���8u��t��x{̖ż�L�I#{�SI�It�Ǎt�Oa�^9$���l�Z�2wI(��� < mT�-#���?��N�������ܾ$�Ho��J%C;�]7�T���.ڻ��}�q�n������	k)g�[�R[��89|��M�a2�9��
�y
|3ҽ�ٯ2�H���BI�I�=��3QH�������}����A3�ԈJ<�grX1<d��
���C1v�Ͱ5n�B��uci�? ���  �~|:��8�.�Q�	�U�Գ<�L��IE$��w)5޻!p�%è�R.˗�si_���b�/�իC�;��zA�q�z�x�-e�58g���ۘ6�m����$M����7�#ot�x��U������^u^�Z�q�H�����-������k�7��|sW�a���ªIG���^Y"f�.���6`������0$���T|A��C��wd�{`�zԘ�I����$t�C�9���np����<,�q�**��|�m��jI,��UD$O��>5;����A��ae�t�,���5$��P����O�L��˙	$�v��P/T�6F�i�#ت�IK?� b��	&F�r��������7q��E4�U5��2Q5�X�˵I����)0Êd.i��.rvv�8���!"^)�{0�w�?z�5kCt�.9�"H�{_���Gz��q��i0�DڪD�ֳ��I�>t��A;�*T~�ƕI?�������U�'�l<4��&�����d�	K�V<A��zN��9�����-��6͠����&I2G���Z^^�v��?%>��3�/�l�3Qr���{��`P��L��|�x�^:�/�н���Jؽ%���z�{�L�<�r|�Z��DE!z�N
u���������>	#���[���6y�{�^��-wE������l�ꯒ׸6�t��ݏ6��K��7Q�U;؟s�]]C���~�����E;I��� ॱ���N���G���=��z)9����޼&#/���god���=��6�Y7N���ؽ��2���u{ٺ�Ч�j���Y�z�G����A�;s�޺���9Y���O��z�P_vn�U���o�>� ��W8���WAՁ��x��Ŕ�:N���һ5�
��w�د�{�2�HێaJVG�>�m�1c�N{��}V�s���}���fϷ���9�ۺ}����.��Ԓ�dp�/���Y'#n���&�=���-��=�4���`ﳷ/���(��p��o/xՄ�
�|���X0�9�`	��h�L��B�_pR��R�a-s�=��c5o��kj�Y0G�$7q��!��Ƿ��t�/���ҝ�ټO��Ξ��pֹu$c�ף%E��c�r��%s�s�u�۝�TOl�z�Z����f�ں_",��{���CO�[,�=�5��\󻰬���㺷҈��S㯾�����Ӭٗ��l��fL�ܰ0���޹��/����YP��ܧ\��A����BX>1�id��˥��z��+��|�o^{����K -�DG"(}��¹Ep�G*����Ud$TQ��3��^�_{|}x}}}}~?�u�u�]u����~?�Ǉ�謰�!"�d���8�F**�&��9�)����S/2?��78���7�~������/�����Ӯ��î�뮽��:�ǧ��b)��+���3!E�R�3�k]�,���b��QZ$Tz��J�Dr�.l�(�CRΪ$�$�/`���m0̪�9E&�%t�e��d�AEUE
lYDh�)%�E�ꁒ�U�ȩ��9rudD�I´N$$�˜�z�L=�W((��A˕PU˒H�v�U)���:UE���.ˍS6QEqj	\�}�iW��|����,�)9\�;B�diQ�((�����d�`t���HAW*�D�q-ݴy,r���y�U�'H�j���2���t�e0����IĎ{��L·	"�N�:!yB�PSN�+Ue]�k8\I*/�-�~��;��c[��q�c{}�w�>��EC�l����w��y��u���p��ÚzK;"�E;��:^k(J��'Ƕ&I2I�o<�I$�#�r�%�CĹ�:y�2a������H:�C�P��'�)}�����Ie?U ���[Fh��`ȿ�,���O}OI �yo"QI.Q���� ���n��w2TBwxa�4v���c6�+6��Z��H	4��i�AOMcK��;��w�0�Bx�9��:dZ�J́-Ȅ�>���+�op��wŧP��HZ76ZHq���T�/
P!>��T��M�c�<[�P%��G<I �q���i����Y���x����ܔ�w�UL]������ɒH>x̯#�p ��� "7�A��%�k��~I��/
Xys�h�;���\�h�� $�oyy����:5�����Q��^6U�x�(��V"�V�/g���Ln{<��?p��8�^��S'����%��ᅎݾ����=/�8�s-.�\�a�K�p��3�gg� ����zd�>�Z{xE8ww1�v��\M��G�Ή={KQ�k�H�̖	>{�i��s73fr�@>x�b[K5VZ�лiaf[�.�,�ͮZ��Yb���P		�@�cN�A���ml	�d#g:Y���kx�@y�|���2��t�O�%�%�E�	km�Ø�!<Uw��I`N�$a�޼��i �]����	���2	lb\��Ú���{5=D2	�
X��,#��ɢ���'��QL!�AU����$��`I;��$[ϻ�\
xE�n���Cyv��5��ީ�ēY�2I$��x�;#�m�<	�5����U�I��/
��ӳ<� ��'��k�X��O6>�=M]��,	bol�Q/���%_�~�5 ������`Kww`�),yU�}Ǧ~��G��wd��݂v�,v��qj���q�����㻚��G��!���]�1��b/۬�� <<8��I�����(&��ƭ���Kk�m�Sk
��$N��M�X�Rk��hd,����]�lP)F�jB��[,fсshgE�mS\�%�M�ٴ[e����1ً��1��X_F�W)�j��V�P�óP ��TB��؏cZ�0�m^�(��e-؀l����YC&U)�nf�Jčm`�֚�l�jUu[L�$�&).6��jG(���g���t�_�#�`����ԥ�j��Qԛ$C.��r�:�u(�_������x���-9Q0X��ؙL �Ov��;�}D���q�{�$v�Ȑ�Y�/�:1�(���27����5㝮֢��f�L� ���8�M5�6�_¿yg��H�}�ЅXM6�4��>�ճ4��L�\�J�{��!fc��-��{rd��v��$8���P�����wgq^R� �Q7���v�7	$��d�кQ�z��Kw��m��ىB.A<"�Qx�,<H�ȉ	L����mVы�%��T,I�B�m��q��k���
֧�,���lR(<M�WZ�A�(+r˲$-j:"�0�`�K4'��,ċ��^"r�l� y"I`q��H&��~�2��
������,	c�ZD����N�<AB��x���4�8S��V�R��z)�B�
HQ��`{G'�<n�Om�f�vu]��3N_������}����oD�\s���\'��g��s�ߞ�~��	?N���Ï �<9�|���DO?{�F&o��%�<�[��Z���>�O���X�tb4�\y���v0@ �X���خ�A �_@�2����X��y�c!<<Ar��G��� g��Ř�%�b^���$�	�q��H�͚����|L���MC^�O�b�'1`x��D�!�;"[̕󚾸�Uް�K��HL�-�-8���3'�ug�f�oni��l���10!I��ກ�̑�T��k�U����l�qY�7���@>���~��أM|�tH2{'"�,��,N�!vm���l���z�. ${�e��Y�'� �D* ���wL���Ok�a�]�A5q���7w�I;��E.��W�+�e�E�ӸQG�v"�Ia��'�+�l�gLDG�cx�)����s<S߄@�!�繧�d���I�kE�.�?<��w�K�ڧ��\]�5�!�f9��ǁxxq�QiU7�]}�NaC~��[S"2M��3 ������F �k���I��kN�<��u2E��l��2 ���H��Kx���=���FB�x��Cā`w\̐�Mv�ϢpR� ����Y5SQ�� ��Ϙ�,#�f|�&l�T���G�v�3�k
��"B|n+�3P���f�V�QjZ3���\�i��@����	�IS�$�\�� ����Mı,K��w@�d���=�L9Lzwf����$�]�2	{�#H�(�x%vܰz�H���#+�c ��얒��2��U��xC'�{���VJ|AD"!7���"M���֚ jo�>�w�	�vL�$H1��$��}֡N�i�+�[��qn��g"<�r�C�H$��sGs��$OtĐ=r�mJE�
�S�R��� ���wG=^ޙ:uw'�%�|h�UI�Ō�y\=@���\��G�|{k��^����8Tp `��@3�02��>�xq�Fxxq�TiD(3��7��<�
���b�ш4(�.D�$�C��mzr���`���˲Z���0�'zc��1g3��L ��ZK�X�iW+����&�J�afU�3�����
z��
""�{�Y�d���N;j8�=�1�Wޏeg��� �6�ĉ��ğ�ЂNb���h��\TzV�2":-�4�{�2d��G �5����xoFd�od�܌"�$���`z��\�;# H%�֬V=Xwƨr��A~�HΎ��*܂�0DB��x]9�S�d�V�v�3�9�F�̉#�z�����NC�7���E�z�9t��Q���D�L�Gvl�.�J�o���΁,	����N�����V�ወY���G����8Z���ܽr�0��l��غ{޷���������!�C��W<6i*�y����[�2yy�����~8�O<*��	�;�~�y�Z��'k��ƙNZ�HPm��DA,Yf�]]�dc��Yr]f�u���u[�pP#[b�3�f�,�[���+��t��8m��Ҥs�ƈ�6I���\*�]-e"D&��VB�*[Z���3\Te�T��f4,��A%qU�&�Ch[�ia� ��59��ŴRn+q�i�jUf�R�]B$	Y{R7���׹��Miq*2�\en�A�6��%�ګ�\�)�j�h�%R���b�ш=B�|w����'�q$�,Kcn�����=6c����,���1�Α,	>���
��	��Ʒ�[�&d�eS�<��mPO����	 작.ȱ[��$w��YO^�t�=Q�b�>�/PБNa��+c`H%��� �M�l����Y�#��a'�7 I$ٽ�TH�ܠ����w�Q�+}������8����T���{�&A����]>"w�]T��%�6CLzE|!D"!H��'dK����F����%a ̿P�}"I;7��J�ظ�:WP'��>MxA�Fl&Kn�˴]�+��  ,�b�4�Y�,1�\�S~w�X�H�lL��w�~�${�$$G�R���/\s���艆�wۓ$�p�܂�ш4��r.�^��p�K�ߪ��5��.��׶��'6�dez�j�k�х��^H��ϛo@��g��]�=�����u\wM�u�]�ڧۯ<
�<�+K`Af`�����4 �7��y��Y��r ��n4���^�Q�<<O-��L��Ājw��� �̠����O�$Ƴ\�N_l� $��i����	$�@�^/�Q���kt�]��h�2œ̂����
�@$��U����|�~��Zr.d���x:H�x%�13$A�]D��uR(j�@O�E�j$t�$�Gt�*�����)��GG}e�	e;B�]��.ܤeɜQ�E	j`M�f�cRxz}Ξ,I��(�D�D(�.8�A0�{%�� ����bc�n��/��zy�X�=}�O�i8t�\��TzrbIV��3F�ף�l�L4��� �t���K�ÑOP�b]l�>�h��$��h[y�˙��މ`C�v��sc��»�1��k�$��Qho{^����1735�K�x凎���4�ӑ��s�]y�2л>��XH�d�g0�sۏ3�ÏҪĈ|���2ɔ�� K��G1-n9J���`�j��s/��.x�%���@ �[��D1�����-�����VS}<.�ӈI(J��Z�,�� ����1s��]�"}2,n.�K�K�zgYn��n���>}�ǿ�f��bWS#�v�ˋU�mp)��`��`X�*2��V���^������	G��<vL�1@Tz�I$��� A��n��b�d}��\U.N4�D""
�����XQ�}��W��AbF�䉆�>��-,��,�'�T��G��߮�������;�d{��mD��Iv콚� �y*���oo���&ղ$@��������1��]rU�~Ήʃ=�:	;�����[yjD�%]���l�щ;���O��B�F��;8\������e�#�����p�NoA������{m}��_��8����.
��Q�9z-<~~š��������4*D�R�@���K&M��:D�qƪX�üc[�\L�$�V}"|�L�5��;�o.dI����c�b�o;�n�92p��G]P���4rT�u�]Is�.YC�֔M����΍m�C�s������w�~:�0i#x�dă$����I$�����`>��;X*�b@%�{:d['סx����#�vvu�Lo&������]0, 	 ~̙$c=�lCH�޽�#�s��D�jM+N4�D"���ِJ� �	��	�)���Ky`B��UT���,�	j�� �v�v��f���9qdx��~�חy��c^��X$Tz$�X���용����$Z���^�5�&��,:}`�P����l��̵�tH6�wn:�����-,��tKHl}�t#����n��h�����^l���G#ZW��B��-w*��S����ss�^�E�ӽV��&E3���k�9w�+�7�v���K�����\�(��������9��1\�6���-^o�g*��C��9{�w��Ρr8�a`Q�w#�/y�d�w�7&�;H��Q�`��`�<��~�Z��7���vsz��K�����z>Ī�˳r(b���0�O<IC�'�f�e����!��<����9x>��Ԃ�ç��|#&��T����z�v��u��;`��v�o�����;$��:�]��ٸ�G�.ӎL3�~��U�:5�qư������:-�R�7�:=|�zf=@��p�Lm^��h�km�o6��=��{�����l9B^#J�g%SǼ�x�˒����>g������6t?߮8�IR�MG���}7{�7�QV3S^�~���-^�������P��|���#����7,����x����[�l]_��Xܥ�������o|�"�g/�K�Ž����ot_��_�{��7|��F9k����o����K�d����a/�..,������ ����4���5�47�r�1/L�!�8��e�,y�ɞ��|F���S�n�-I�[ϳ�"�/O;ű$�{z�cX3���n��g�*�o��������'�A޺��^���My�x{�Url��)s�EE]dN)�3VN1�k��OP���=*�s���8K��&�7�y���|����{�2:R�RK .˵K�G9'~�.xO���*�S(�
�h�9y|{~��o���/�����Ӯ��î�뮽��:�ǧ�����32Q~�#w=h�r#�=CAV$Y!�	�mO����w������������yu�]u��]uק]g]u�讲��33&�����(�+,|�*���D�T���TUr(#�����i\���I) UVT��t�J�E�sc�!]�8!Qq�Xd��DA��J��r���\=J
��D�I�9�z#"9��*(&�*bI�Tt�e�yb�ڥD|�Fl)�OU��r	���>��\�tz5�!�>J�=̪���/Z�\.9$Faʢ�SlO���AT�8I_;]\�s�[��=ds�y8E�9UAfʎU_�Pd�L��rNˤ$ʪO����]��r�yRt�J%��j@�B(��G$ ��؜H�Ju u�����/ȉ���0�pM1�����7�I�U|&1��d���5.4t�k�|��MG]l�1h��j a��"D�GB��ˀ���`K���ܱ���o4�ҷ@���Mi��t͍mj���`"1�ׁ��&����3)�ۑZM��/3�S	68�W����X�nYBڶ,re�nHk��K4���#��d��X�ܭ���3)5���1Ύ���2冱��yS6�#T���3GJ0���m"�R��863�J�&��!�6�m��Z�0�-0p�+�W1��ى��S���e�b��-rJ�:�[r4er�ř�,שk0�"]ft���kH5�w-E���K��Q�lG;Aư&h����R�Q������1���5B�X�6Y�Z�w6��-��nM6t��T%�-Bb�Vl�+��B���%L�YQm��ph��ȸ� ���
)V4b�1��i�a��4�e.ta̎m8�L@��du�sRkm���@ �ͭ���0�h�-­�.�y�d�ɐ�yYl�Q�&��k/:c���y㭚��aDmR�
�"��#�-�����:���Ʃ�օ��mѻlj���	���R�b���\�]6��)Wk6��ؚՃ�i��Mm*R6�:Z����f`���K,%�Gk11yf����\�2hGp!v�%)�w^�֬�u�4�0�Wl4x� �rf
��H�H6�E�K�xK�.B*#cQ��M8c��[+M�gQf#w5������
��RKc[�3^��K�����l]
F�f�����VQ�a�ڙJ��U٥.Iy�:�XC��G�1�&H��^Ycq��66�.�&3&QCv�[�^e�g\b� �m2��7m���\�r4�[�X�3tʨ���%�%ݶf�U%ݚ �U�]ۄb�LT�1��D`�IUkaX�h5ń4K5�ZO�7�<\]iU���`��0^�г^�S����Ҽ�`�qj*b��S��R���;�u ��<�|�T�6ݩ��n�Q�{��7�~n���v��ˀD���D��������S腉YJ124�u�^:؄C�*�"	zR�s��i�fQ#]S�,���M��c��K7Q5%Ѧ+V�i���Լ�*��L	�C]6{mH��[iS�m�B�A5"�!k��h�ዡ46�M�)n(���Z��T�Y���9�J�5m�3(+�`-qEv�uٍ��.�<�hU��6�m�R�[6�)��80-�Y`��-X���u'���<\oY�7V#�`ڸM�4�0(�nU�����!��@ث�:;��ъ�Ԉ0[�&���P�$Ƕ�H$�~����u�y�z�]�m����	1��.=g^�Ar�с\S�@��F⛴y�w�כ� C$@$�{)��H|�,H3�+Q���aQ�)�	FEax�e^�A�0ή3���{�9�(��2�H��".��;�/��d�<wE��H(8A@��\���-��H�K۽9۽���46@ ;u� Wi7z��N��29��?�$�$�fĚqW[|�h�l�I���
��m܉bn�τ+����Sg���C�A��OqJB�H��su�eYj�e8�%���x�E�7	�?�`:_��Þj��j���	��t
#w:$j9=�3i`���X����ҥ��x* �Wu̴z<�v�ɥ״��Uz��y��x�=������;	%�0s��vӝ��r��j�̗���;;#/=|Ɂx�'v$�aJx��,���<	<<8�č!J�4J�AH�Qq��_:��ϯ�����ߦX�}������YQ�7���r�сT]��X�$A�މ�@d�}���a����,��0�ٻ� ���B�rJw�Q�(����Z���bM�zzh�|��A���7� �}=���<�$��{!����X�x�D"�(؁d?^3�����7 �v}PX�޼�bX����g�!$P:����H񮗶�x�U���i]�I�(Cl�RSf��F���"�pG8Ԑ��N�<�\�t�ˈ������[{6%� �4ouR�l�����YOX��=u�f��37��-dRta�
c�u��5��l���`$@��CH/�ɡ��
u���{��x�nPP��tb(�kϷS$�Q}�%�˲������� ��~�۝o�.i�۷�q�@����t��BK��.�T���~XE#�D�j����ۖ���˱�FFyzA�=� �|m�
�D��0$3���	��ǅR��)X!@�2a����n�zd�@%��̐&<M��<J�	-���*{�sP�`.m�H*��I �S=�PK Wo@���Z�,��wlH)�4!�%;�(���Q I WfD���p�ix�I0UT�v���x�ϛY<�AwL����q��<t��>pk|���y�hVZA+���.l�Hhk��\����*ͣ��%�x�ǳ����Yb�8�g�d��${�d[���B�y�:�Z��r�X� �e�#��^��×��DY��bK��^ʈ����a�I|홦H��@��Fhܝ�=IQ�u/C�
����e���Y;��	$��D�(̵Nw�%��g�P/	%�wl� �~�F�B���ã!Mut�TP��h�ɰ�U�H�I!��I��pf���kφZ�����/2�K6C)�/*�������gl��J�����g5�=�`|��TG�%@�N���x<�G/1��=9��c8���3�ÏUBPAT�D�R�%�}���5���c҈.�;�E��$�{@��'ݏ�j�Z�	�bA*�$K&T��7�X�Gcޝ�3q*8�'.&�.:	.\����ͳː�Ֆ̤
"�2�/)��h�p�~��y={�O�֢8����M��i���}̉`I,H�� �����=%�"A ޹��_�;���"[ވ��!n!�H����o�H���JH%�o�Iv[�i��ȳ��yٞ���w.\DG�>��{�$��Mw���.�ٯ�ݍl��i��Ē;�d	kd�z
�B!;�h�F߭�Mi�>G�hO�=I$����,@ �w]��G��N��j�o72&���� p��Bs�@��\/�2Ks$�.6D��G5{��N�X��{$K	o_l�>eO�p��ftث��טuBMue���⭳��%�Ng�צP���;l�	|���:w�'��>�ǰ�>x��ۺ���^��O�d���*p~ |Cߛ���7n���L�((�t	�	�O���罄��.��L�����I+��m���hw[�@1�u��ۜ�6�11�2���lcV[f��l4z���a��l-����B�������6�a(Eg�[������䙭�m\�k�ZR�yme%C f�����5�	���b9��F��6)��m�V�)˛#vye�[�A�h�0D6Д[R���<&i�H�]sufFW+g������s��G����g�!��-���%`̷X´t�-MIiT���� :
��{�|�޴�
�#q���n��R������tI$�ƞ��je77���3�l�vc&�H$�w�fI��E@���0j�O�2A�{���D��� ����"A GvȭK���3t!��K��x�"�݋ C$E��ș"Y  �\����$�%���,� �&+vfM`�=�A�˗���G^{��޽$|ȐA >uĒu��;�=J)Oz��d���y��Iч4(�E�c�� �{w�*=��^��%��y��<<s{�T�/:-Ĭ)	#����=
�u&+�4���i�3�t�@r1���]��~�佾�����2 ��u�� �-�GL�����{XFg�>%��^�"Z<meB�0�;�@�D�K��o��r��k��0P�7�H�h.��r/�<Ey� u�Y��z[���Bo=~�O]�����u��30h���,Þ8�w�����ݔv�nUp���2�}{��L�|��tQ���a,H��|�N;Ϥ�m��kL���.��L��54I �t��l�LH/�]�gZ/ѸǙD���H"�&�ޑ$�]%����
�/��Q�J/��I~�� ���,�;��[�䅘}e�5�.D��o�(;�r� �;qQ A{6$��K�{B� ^�r�*� �y"Iy�M�����lt~w�ݝ�xG��oZxB飀-��B�X1X���m�BڎҮu�fn�	��J�~~p��t��.d�M�lKIm��X��5Y{�X��dH'"�D���e�'*��g�X>؟x��R#1꺄���s ��w;�����������"|��˦�#M��<A0�9�E�$��${}Ł ��4{��W�p>/B����e^9z��ȣ�}�澾�7w�rS�_�{W:m֭�_e�^��;;�������/~ϱ��x8^�����>�)���-'��h�A ]��4>��N�t�$��U���/,$�ڙ����1�g�ɼ� �R^{w.�HxxSKg�Iu䴑d�v)�T��묁 �/�$4���3��k#��O�������8��#cZMr�����t��4[�)*U�,Y�ֺ�uƺ�u;�/�}��Z�m~�~w�I,S��#Đ�t�S��s��ۭ���X$쾑3�B��I�ÚM�\��A�59�TC��*�wG5"	c��q�"�t0�o�ޗY@��%�����(* B�Q�,A1��!���&�b����p�#��%��"Sݰ�혈�&'0$>t^����^�d���H$d����)����<�L����VA�no�^yof�P��,U��3?�V�G}������M���߈Y�+Yo�}sFrS���W��y���W� �6�8����������Fs���xR��@�#�?v4�I罁ٱ�e�r	o6Wm
$�v��Kk�@�>��Z�����߿/ߛ���M�s-�P�!�Q�&�7-yLK���e&��Ҟ|���j�c�~���~���u�I�I��N�b�����Fh�_V�%�1��2�`~{r���."P=u0�xLCG�$z��D�Z*�D����%�"xO^^GTιCŚ��8ģ|����f����1�7�r�@$��D�A �,7~��J�q����ڛ\��̉�(����j݀n�"��U]Q�M,i�]�2G+�F5 I#�*�b�;�}y��ď��&	����9��D;�
����#bH&��$ѐ�W9�Y��� �X���!���&�������?g�����,p��E�҉**�70��� a�~���/��P�+<{�S�}S>Վ�i [��|͍�q)�ÇT3Co���q�&�J��[�������h�1l����6̹%���t��Án��Y�mZ���G��G��iT�i+/kf�������նa�&�T�	@(v�e�Yp�B,-X��ե��8�`��R��r�3R�t�;lg+K����� te���LSB�e7Xg���$։+2�������WXShP��5�Y��`��!k��ܡ����Ύ���3��'gsF�q�ۋ�����V5l�36�հ�{�<�Ӹ�@�������+�p$�ٽ�c/�z��A �t\	��"��x$<<*�7�ĉ���_����O��A ��ȒI�ޙ�)>\d���{$�OXK!ˇp��D ׎��d{��A�(��',d�RP���u��<�b����@�R��*����M�=q��b6�!���I�{fI$�{3{cʦ�M�d�ۃ�(�P^ B��7�8��Έ�ʙ�G����������	�}�# D�t������������>����׿����i�"�tGcX%9₰�6��2ۃU������_3�S�Ϫ�n#���68�N��Io1D�@���z�f@��&�/gH�%���D�#G���q�],$��KO{�B�(���5�ӈs�����q	�y��=�4��.6[�.n��R��wݚ�۫���G%Fz��x�ț�/z�K�����8��x�ߺW_\ᇇ���ih�
���y����������4]}��$��p�"Չ�uL>�Β��x$:�3E�u@�K�fK�i�X^a_����$�}}�$�"�{`SQj�)m��������_�/Dǵ(�}~5n����$�z$H�{�H'_�Dǽ�}y�ۗ�͖��M@�<��d�� ��P E6\z-�6��&����jt]�#=�u&4Ɯ�i�޶�X���Z�tg��<��������t�̦��ip�n��GE�l��v�fmjTλT��]�ٻ���:�S]���n��Ę��H$s�K	�|�����lMv�5�c��N�̘�ӑ�L(N`U S�D�1ܩ�e�%�� ;F�U-Ͻ"A �S\-Gu����LU�j�@�w ��� ���q���9�J�ˠ��1u ��tk�ߝB<q��n_�7'�R{�}������ �%�t�����ý�en{�V��@��_�Q%�J.�ﶵU��=��Ç����ڳzXv-�����y��K�h8}ܺ�> 4.��ܾ���V?{�c&r���a�w��##83E���u��A����A���؃�9�%�w�+j��i���}���G�#���7�,Y����yU�n�����&�����8s����R9�7x���j�<S��8��{w�nxd��㛕%ױEԭ��^�GB�>]���Oxg���1�gb'PÕc���q�����T�˔�z��>��{~J�=�Ӊ�hs���9O}��6�%�{����/���1�rc;sG�[�L�����6F�7H�<Js�R+��\��
��X�W���m<�l� �$3㏞/>+8-�Dw�ʝC����;�{oM�^>��Y��<=r���T�!m�#`{؅�Gz�]8�o�����|�!w�gjoƆ�d�ܔ�:<�<~zU����y g;��T����n�h����ꭣw�T'F��E����7���L��%��gF�gg���|¥8gg�b����}'Z엮���>ň�'F,((�Z^x� �s5{���|�j��A�&h��ݲ�k���VMz\����Rl� ��$3q��6R��αP�����ӝ�D��a RG�~��薏���O��p���o���s�gJ�� 8`�b�9�U�<rP�s ��x}��X���w�V�nX�h��~�����������S���U�P!��D�zeL� ͽ@Lj^�x��z��pt���*�Bg�e�Q��U]���8��NT䲋�i&&b�(�ʩ��{{uׇǷ���ק������]uח]u�^�u�u����)����0 �RQ�X�a�{���0�N����Ǉ������׷�����]uח]u�^�u�u�㦨h"H��Ýؕ���r��UC}��ǝ�W�TY����"�N��%WrT\�y	\��'����U�u��FC�YC����v8����ˁG�J�7<��t��IPG�p�_�|��T�J���r(�w'*>�:���z�X����.	7��wDaҲ+�\����(Lդ���/[�۝9Epu;�U˕q:�9�ABu�=B�2�ԧ�p�����.n���ϥ�\����p��'�����*&��Ê<H��}�Is��ޞ���~�D� *��軈gQj�{�(�V��b������ I<�=��U��I#��G�Ο�dѿ���A,lZ?��0� �gD�0f[�v�$<�A-��Ȑ	�wH�5t#��<ke��B��E��s����[!
�Y\�̔���p�a����b@�X�R͂RE@��p����
eq;�#�䋿tL�V޽����^�G�g®������0չ���7�,V���}w��Aă
�XH$��ޙ$��e'��O~���rr"�!	�50p��[\�I�ޗ�$�{�ڴ�McE��$s��	$ow<�R�q'؊Ӹ�A]c��*�z�h>��ı=׳,H$��1�_��͏B1L�=�ݲ�섻��W��/=��wx=2q�~���o�ŋa�e��������&rPyB ���o2�2f���,��H���w~�Vs��!�Dox���_�ɘ�h��j��H&��e�$_{�r�(���7l�x��z]��k��2,�X
�P��;W���Xɋ��Ҹ#�wv��H>�:�	@�]�An�peY��j�#�΀$�@/�r5l�U+�=��*ZA#�2d��*v	E"�ȡ�G����W����n�1��	�m�y�C��wt�� ��{r�J&���U���iZ�E��j`��l�I�`o��� 3�Rk���| �$k]��Ē���	�G��"U��P�\C��4�ߺ7De-�Xe�w�(�_�d�$�[�1����S������M�6����t� A�A>��2D�z�M��{�!�7{f4���#�ޝ�i��25�J;s�~��M�V1��K�m^��.�{=������i��8]�����u�w�������˗���;A�a��o��y�Ϳ��b֌��=���n�:��5���6B��G�����uFkF-3�;E�.�H��+i(�W��&,fƗ�� �c�HW\Yb���ƹ�7LLF	1�lqpl��n&�Ֆ��V��&�,�ƌ0�J�,ur�`\mh[.�uf3̚V�A�vm�H�5�9ѭ�1P3S�v�iM3fÉj�!*����Ea0ǖZ�Z�Z�(�
���mCk��3�ȅyc�����޽<����f�am�h˚�D&�ũ�$ʐt�]sv�X������`��w��ɕ�d7�fK	g���;�FFqP޿TL��Ad��-�9�x�A,l	�w����o���Y������� ���1,H��$�~�ZHR��t�;j-9d��"%����d�B�t4�s�_��пz0i ����(���	p1T:/B��nz��x
���"HGdNvL4�A �mѹ@Wwd�W���Zlc�ᤖ�OD(x.!���)�bK�D�vD��j��<�'�J@�w��H�@'�d�$��/Vj�^��z��hz\,b��0�CL1�@���f�;XZm��NmQ0�����;�y,_�P��P.��>�:��@�@[yA��$߆^ViOP����샭�� ��+zw��R6��xȝu�{��7s�]qq^O��f���;���k��1�U����� {�s�\��1�)�synZ���'���^��?�}� �ÅY��߮��h+7�z�)��v�2H9�G'�T�\\_tm���(!�sdV<ƒHL��S	��;^����C��k��u��%�펗jDU^����.!υ��7���7�=2�1��v�I$�"�y2K�u�K������:���
��^(�fAU�� �K�d��e�?��m�v��}wR$����X��w�hV��e�8�i��������m�
�l��2�-k\2��!��qe����tE`O�B�����.��,H,/{ I--l��t�+�j�{��Szg�Ko2 .ޙܫF�t� A��bze���!UoNo�MDƒI�W�,��b��X�4���{#OO�%)�K��C�hQG��z@�z��,�[^Ȳ8�$X�s��:2d��c;�>��G�Y��o�ַ��޾�]z���~�<���~s;�a�B��'�E!�3ٚ3�v�G���n����v�	�\# A2��O��<	'�:AiD��D��+n@B'1��o>����<'��
� �c�J�n$�I��QJ��@!Wt���~꫐L�L�$E��Ц�([>�4L��4|�s��ˁ4 ��T	� g���X�C�\�l��nMt;�u������:�'���qS.zΆ,��-��mחU�ѕu�-�Ï_~��snt�
���6dAf̂K�oP�zG�$��� �b��1��^"v94Ht;�ZacX�L��FY� &���˩S��Yy����$.�'�t���RQ��ѭ������@�E�QO�2�q �A����1/G�� y��c'��H$�^%�� ���LuLmgw�n"���e�K&H����@�ޟ��s��t���Z�]�Փ�`�>��m�y㓦��T���^����J����qZ��,�i9xn��7|3d��x�>�~8'ܼ<8�Q�=(�;ފ�>뇀C�.bP>Ȩ�I ��>�8�_�I��N�vuP$���$k$	��F5y���x0���g�g�7��t�m\�%HD�lMn��
�l�5��dɭ�̦���|����7�y�sW��$���M2����]]�G���L�eג$=�p�s	��P�Uɺ+��$k'��DyH�9|��<�P�.^驩K?EȐm�8"Yp���{ǹ��zn!C�p��
�s����@c}� �O�|�k+�̐/�njEv��"}dw�>໻�0bI�'�E�u��@��8$xؒI[�6i�.�����/#��p �u>c@
�7P!�	��RΩ�H$�fGoA͓�!�J��	�D� {ݑ,Y��Zy�Ә/����x�|�FQ����G�x�}�}��P�W��ф;��A�䜁��s�=+)X��_%Ś;���=�AoC��&�~ͭl���9,Y ��j�H��>������1l)]�Ѽ*;j�i13�f[,tuU�ĥ��v���,�%,�з��X][(�e���֕��[z���VZr�9�R�&lE��1�����p��EM��zf]p��jt�PK-�R��U���t�[jR�M*���8�����c�͘%�J�k������cʛE�Ĳ�$�e�ɝqz���mK6�C%oυ~>���I��]�����(���q��KQ�m��3�5�}�r	�Wt:���\�7"�|L{/�H�K�tɜ�g/'L�=�ȐG�gb�L���P���{���V�{�˪���0��ȒvJ�2d�K�t4�޹76�@�okc{�J�0� (�T1�f@$���$�A�s|���8dg��I;w� [$	;�f=#Ց
��H�<����q^Vy�x;�v�5	�K���$�zX<:�O��X=�&�M'�\wx0�P)����eċd����c0���,tLy�s��{)��C�\�6�4��~����ǿ?%@��ҳ,6`�rY�JT6�+j��M5��ˡ
�A�vgIhO���WiZ0x�1Ē�d��)��u5<Y�~����� C��D�i��:���\��}�P�,���g�^�"�J�x���U��g� ��k��r��!����I��7��<D�Efnfڳ~{%֬�D�R�E�������e@H�O�>��$������*a:ﯜ��PG\����D��G>�̣W��ɣ4k�	�AA�P%A+X�*f@ �U�D�X�|����1�%z_)����L���<��6U9��D(z���4����<����d�ܴ�U_@栍2@toH*NE�1��]�r�fn��(x.�!��Y%2vvD���k׷U 	Y �gii���HvAn�L����U:2�����h~{���ۆ�d+`��K��b)3���\�7WJ豍[���d6S���a���a��w���}�2bJ�ȒI';zdכ:n�zfjJ~��3S�-�"C�l��GD��x5\�R�7�W^��^��I0ϗ�sy���2��v���9b'�T��>]` �'Q��c�O�Ad}��$� �h3�̮�3N}b��r�"=K�4��h�Wo�\�;��?x�{�p�Ip�yfX"�A|�Q�Lo��}K�t���������\yw�@O..8������mK|fIb$�o���cF�ӠPtT
}�����;�	c1����;"=�S$�����
�*6���6{��-�R�0� (���?V�i�Wuj�������%�6�`Y$�vL�9��}���ߟ���S�;��OK����v��e����6).u�j�U� B���nru;�ߟrgT�t��{�X��ȒX�_����h�*���Z�<W�N�@�̙(l�\D���Nq����-%��^+p��%�pg��Ā]��r��C�l���}�ͺZ��鷔��ѐ<	ab�x�A���Z�bؒK���`���)���0�>T����/�2}�m=���p�D��Sfz*7�lC��%�$�_D�1��M9�������4!ow(w��V�'G���f�����F��G�ī�|�pz$����^���R�1Y��7X�4v�-�ak6��d��x1d�����r��묔�F΍�n�A�P=@�k��1��d"G6�E8��w��7Q0$��!��"X�o~z�w���;s2�Kt�l�W5јc��v�j!��j�;i��l��u�(y���Y���?~�V�H=�ĐD7t�ox��w���<�XAm�̹�H$�èj0�è��'�TWOD�Ls����ʚ�)��m��	$���2��H;��O�?���?o1�����AsT�Nl� �=s�@�	�0�;�N�r|�A�o6$��hP�;
�@���U;D�~@�1ۓ$�:@�މ�9��1^��>�n�%�	�ukg&$�I�fĞy�\�-���*l�� ��Ȓbw����"]�}Л_'��R�&��NY��{h�!S���v{�\>ԕy#{9.��(>O��,jE���{���;O�ou��۝�/w7��)/9������({r��=;�v{����0�sOw,<+�s�{���� �>�o�����g������kG&Ӯ$�<��~?_b�<5�}�İ[����{;�XW��4e��o)�nnӗ�8߯mJ��_Σ�d���{\��š���ny�ܼ�d��q{5�亟`�d65B��ڳ���m����Ӓy_'"��O`�u���v��]��5a$7�zb�=�{tf�=���Z7����׬����7�:���g;��in���8 ��!Y��7���ӛ�9��� <���p�*y'&��{��7�{��ˮwSv]���6��N���x�Zꕹ�Ć���9�}M�;|^�C�i�{���O�4.���X�ẝ�=�>���wzO��{}�Ń��)�|����fv���^��o�.���h�Ӹ�1z��<`,���d�;w�}��y��S�b�sý=��.��{nZz3H���k����,�|�/N}1x'��zA�</���OK/r��ra<����L{V��m]�w*�������b�v%�6c�ra>d��8۾�	�j���{���ӵo��co��+����}���R,�>ׇ ɚq%T�;��P=g�e���ݨayV���v>_yxe�6��x���>�:R5<�\���d!���p O�cr�9\uo>x^�QM�T�/O��돯������o���î�뮽:뮼��:��1��M|I\�@U�o=���d��'��zz~>?{|}}}}}{}~?u�]u��]u��]u�נ��ȋ�Ҹ^�s��>�H��8�w��&���0��I�Ԫ"�ּ��1[=w"�a!^w�̞�SI��@Rq�e��s�:�TUp*�г<�L���!�,��
�D�-�8S)�>��O�9AU�U��B��,��l��b ���]�	,J�.b�e�y�4��$Y܄�ݼ��7�bE^oO@�6��c�h��:v��G�ϫ�|yV�fQ'm'�V���ݤ\K�U�N�L��֕�9=rk�-�(_e���,�33E��;a��*�.��:����6SJb��,�� k�]m�"!v��iu.a�Ȼ8���\��ؔ�8����P�E�CZ�7%�Z�.��.2�M��9�C��]^�74�V���n�$ִ`�VaYm!6q3ؚ��lڃI���O�[�P�G" faHE�2�F6#[���)��x��,�,p��eZK	�Z�٩�
5���%�4&��-�	E�aq �n�Ĭ��.X��3��,������g!�6�i��f��Xb���aX0�RM�]v�3<�q���rp�b��R&�e��m�6�)5�Σ�tֹ!�*Yet�"hjx���Ɖe�4	�!��l�)p�"��SBP��)j��P�(��(�ҽ�CL�ńҷv��V�j	��V���3$��+:L$[�4�,F�V���f���X�J��* RƣR��M�a7�����q�t3^\
d�%U��]¤��i�!�EnSi�JPCL%�Zi�x��Xm��a�t�@��kh��H�K��+��;����-�\�4	��u�,2��
jV ��`�v����6U )��D���XJ�0I��\L�0���-�6�je],(�i�6�B��`%.��`�]Sl�n`j�qҐa��	0��Il��4m�؄���*i���ю�l�[�0m��6�e��rJ�j��Z�ܑ����LU�[�p���Q�BӘ�˭02�C:�5��M0��	�C�͈f룼� �y�B�vIE���&���KU%�RU�v�*�u�zͳ�:�Lmq�U*�ixQظ�-d�Wi�L0�%.�t�RW��b+�,�3B���Վ�n3˪XMx���$"�+�6�v]�営%Er����f5�k0�A�ˡ�;c6la�,E�u�Uˢ��1h2G�s�]���Z�7.TYj۳0Qŉ ��C�:*%�6v��A�"���h:�!KW]�)b¼��4H[4���\K]5�F�Y��&��d��?����q�"�#����\8�9V�lgcG��tnp��6�˵�9��]��M�u�Cd��-M-J�
�gLeC�m#�q�΍�l�o'V�&50�X͗H�0%�JE)*�K��%r��L��Yn0h �K�:7����;2��V�j�isP�gl��҅h$�"�t�&fԄc��0Dv���!��L�0��-t(.��Ũŵ�ԕ�P6ඥ�
�B1ߟ��շ���p`sm9�*70ֻ$4R�\��3���(�`DC�U@����B��t
������̍d��I�ggZ�%1��lx����-{"K[62W�s
 (�
�OE��B^ݏ���H"s��G�y�bZ;��U
d�M/��f��W��8�èx.���@��X ��ȐA	�$PW�A���/\��H$x�	9��$�M�K :%�(��P/]��w9��@�"�1A�K���I �c��y�݃Y ��8(]�xu!&�Ωu�n?
��c�ln�"�᥁9ٓ$�L��d�Knт3g'�[Pb<��^;���� i4�S�ں�44��C��av+s�����*$_�к]T����?<d�g�`H�H$c;�T5���G�yz����I��L������H�c�F�f��o�F���N�����N��aG�uӧ�d�x��7�m�{�IW�c)C�_<�����9l旸�S���y���6섡�3���2fk%��@!�*d��2d�&dcג(�����ݳ32�r/U��@Q
P���H��2I DE�FJ���Uԫ��gLH��L�$���5g!�<����)����z�V�	���e���b$����d�HwWH<=N�ٚ����_L�tzidD��\�/�2��dI������="Ug��;$�ﲨ��I6:D���V�Ro��R�t��q��.��a���(\kEh�kJ�cE0�z��~c���AHD	�*8%��ͩ �A9�:D��N[���)x���h�s��H�u��)ܹ�>�zr`H>SՋݑ뎉oro�<Ar�A#::D�H+f��˸ب��=>��K	�b�Ӹ(:*�z�<���D��dA�{O�C��T n�F���Nd����eJ#0�8��yF��M�~>ŝ�����Vv��<�qi�y��Cھ��.*c�tJ�Z� &L�**�c�1�g����^/U��@Q
�{��2�U$%_s��b�de]=����ӂ<�j�$#�v&�t�C�x%������Iۑ ͗��م1iDV�N今�� �{b�I�L�ΙsDyp��:����G���(�����V^f\�0��Kip�^mh�h\	����|��o��j�ս�����A:���j%���t����d�i�XFه�M6�c$�9"Io�0��HD
�mL�
�4�y� �nE]4�M�.�$H�Ι#͂J˯o%��e�@-�����w.bQ������v�΁)�ϸ�A
eb�l���t̉Ɇ�tQ-84ZzwE@��z��Kۑ�͢A�z�Hc�ܜc@����Ι�h>~���w��i�]by���f1�o,:s���v�\^~�y�/��z���٘=�=j� �׈�s���z�����}4g�|[̙�&L1����;��xJ '���El�6�\�ԛ6po�(��\�G<�D�E����C	=�3bs2���!?}O���<�8J�we��L\�t�X��`�W�ɘ���\Udx����뫐�s?������ %��dI$	��`�2'\V��ٌ���{=��e��"(m><r]�<'(S~�Mk�]��F���TX �u���m��70�A��Lh��Q�uu�A/C�dCü$�@�T�ޙbA �e̒O[�>4�'Lu��޾��d���&w����Dj���y
�-�}��!�,"'�y��iΩ�$y����}���h��̛e^?����P<��F�}2X�~�T_���mWY��%��l�,u���O�MML�ޑ �_��g��r��34��3p+�nw]x��'|�qZૼ�\4������5}�O'=�")��y���,��hy
ع�[̃&L�����t��L��1�+r隘q˱�\�����G$9�l�q�[v�bQ�f��и��`7B���p�<˵�P�X����+��Z��MrB�����,�GEs��Z�5�K�!u��a-öH@�F�V&ɢ%�[lXb�V<Wh����4�DX��VSM3�\X��kb�fc0,�M�cI�[ib��̲���ZWCc*�y�j�(3����O~��!�jV5m���B��aI��K.����&�x[D�zz�Ӱ$�~���@O
�y�fN11����Ol���m����Ev:��b�$��%�z<g!�<���B��������n^v�!��2 �F>��B�r��/֧5�n����w%�C�rEw%�dH%��u�O�x�
]јI,^��%��ޑ'<:��C��r�@A4�h��?��Ǩ�#�6ԉ�湞�@�F�z@����p��@�ODU����ww�
]�e�ă��:$��Y�<{�� \�L�H�ۑ%����c8*��|����ݿ�s]e@3,!+��F�c3kvz틀�9X���3���}@{��i~=��Zi��Xz���c�@�O�7n�H�oƤ{�9�8���L��H�tȘK�+�xJ '�	
瞁lU����Z�~��o)�x#���i����Or����n㧾��l;�?�L�XcR��x�C��T�ȃ�1o2�2��Ă��Q Ĭ�Ƙ�d��gƭT��odNř�u�0�*���A7ݑ2�&/���^M�^�0	n{�2I���4�[�d@w%��#�/]%���[d�� ��ْA<۝��H�w�{B�[[�4;$��R	k������q*�ͩ�X���L�fߌ�/^ �|�֚z�M2�t�t�
o=׽��g�
W�h��ex!��Fl�L.���8.v�r���k��ɽ��ww���S,�� P�1$��9o�u�p|�b�Wy"B�`�V��Pw*�;/2��T�@Zљ��<^v�͑��C�0��ɓ��D��i1�'wrD��P3��ʘ�qx'��xxR+úm�A$�e�2A ��8Y�.;N�������^��=īM�Vs��
/�hu�U�|J�/u��W��,k;�kU�������I�U7��@ɐĽK�=��,I%��A��	�L����p����V��:���F@�K�@+�%�.��Y��=ǈ��#@rYUzD��5O�!���A��=>̖#�{%��.��M�/EzD�_��K���]�s�o�/�I���ϝ��>[f�k���n�ƺ���Q,&v0��1���׿�]����5j�L���8}���$H�}�$�����̘얓�S�'r"]��/Q�U0� 
ڏk�ϏT�N�H-s�2�"��7�#5C;�D�)z(w���,&��b�ʁB�\zG5"G���WR�N�/	*(����ɐ@$c�rX��̧)�(�^�WDt�w+~�@�@�T�nd��SR-��5t�ޕ�]�w�J��zw7��s��b��f��1'�׻���g�'����)����*~G��m]�}=�v��Rn5c�	}M��&L��K�d����C�<�����kQky���Qf}����z�e�A�Y��H�}��I#wzd3#j_΄�[��� [��d&	m� �3if��c��`�ف�j�MXcF��������41��;�S�2L�d��K�H��w�
}������<bP� ���B|3lX]�C�B�t��}Ǳy��:E_�F��@ �}�LFu�H$^�ͣ��9X%�6��iB}�v��%�� B�(��e�j@c'Y�,[�^�^�+���2!ߺ� ���d�Ƣ�REr�Pv>�$B~3��>�'uv�s݀D�	}�!�)l���Z�2<i�t�x;�$��� (z鑬��Bsj�;��K�n	m����LXSq��$�l��ʵ�=?��RT�S��@��Lݏ��[�r9_<�����t��b9��1�zp��W�e@��`��TT,�����2ם�j��Z���͗E�b�Rj,�a�i�]4�D�4�6"��av�,�H�K�qq`� ����Z�n���ؔH��.�&kv)�Ff�Y[��Ҍ������e!�6ш�b�w����I�bq][d�QN�Y�ͤ��"�b\�M�]X�͙���jUPtݵ"��[���05۱�C�la H{�=���J�(׆(�3���l�B��Vڬ	�`ҘՈ�q�9;���G����	qx3��$�n@�H�v̱v�j�J��ªh��a)�$���4-�V�� ��*�
{fK�Dyeu�G��5{�$�K�l�,������e^;bXx@]9��D��%��QۑD���}k��*�����@"��D�A}퉟i;pa:N�@�T\TS�xA�=9������v�%� �_D�A#�FN׎�rw��$��u	8-c�!ʁ�^ǲKc _z$i�z�k�X	��v�_�%�Y0��2����=��?g^�'�35��MkF��ȷ6�f!6��f���à�Sf�˼�+���q\"��zɒ@)��6�Ƥ��":D� f��f��Rʩ�I_�bEF��w��K��5EWtH$��H8夜ZS���g��{�)Wo\���G����z��7|���C�m{���������c�+����O��0mS�t<�ZL�S�@�I1�g�zd >�9��c���AO<"`�<C���G����
j;�$�kkI�b��wW��� ���>b�;�%�"�u�aCÄ�RΩ�[���nK@��D���	$���7�i�]=���8�-�i ���sr�T@�#�\Te"y�Kw�ACևvC�Wc'�(������#Gt̀nC�s�����'�_��.���,f��Ĳ�훮�����[���y�	��N1"��P8��}���M��iX�!�zd�r�w����Դ�<�d�H�L��s<�:xE�A����L���ziv/9�-�:,I �m�sR:���6Ί5{#���O�j�ወ�5N����vC	C6����z^�"+D?m��C�*��	��ŷ|.�^�����r���.���i�x���{QL��k��l��C&�7�w�[�|�����{9�ry���k�!;'{}��n疾������|@�q�T;�.E�^S�1��G�p�=�Zޱ��絅;<�'�x���}G%��7�j��Ӿ/��(�v��{������ؐ��|�8���sႦ���\�!�m��k�	��=��؃��o�#���n$�ᗀ��%vU���=�.8�w-��$�У�V�uy�#
$���s�������N���2NΏ��gO��|�d��U滩k��&Y�������þ��jU�'l��+��G�iƀ�;N�G�=�Cܟ�,�ʕ�W�%��,l4��@=�R�f��I�Z�'��t���dv�� ���:�wڵ������g-�߼���t��y�0vn�0a�z{6C�i����Kݷ�R�G^7��}�u��S�t��{	e=����%��&�:��m�ǩ��N�=S��gs�/BԒZ�񺏣/�_@���צ���w�o��
h�9jɏ���x�z����
vĥ��ѯ��{����{�_�~Ǜ5b3�j]���2A��<�>�|'�m������z=�(ǫ�{!9fk]l���A��^Oy�9hh\��u���w5�/M���NO9o�
'��L��ĵ��=K�q̇a<E����_1��D�4����F33g�y��:�%&(�؛�v��}[�}ȅXX�1�ƌ�������돯���������u�]uק]uח]uׇ^�8�IQ�i��Y��a2�z�������jE7$���w���_______��u�]u׷]u��]uח��2�Ɉ39�
�:E�j���S�\>����r����t�<g��Qr�r��� ���y�r��˼�NDʺM%Y���C[$�D["Ib��."�"��{b�RAr�*uYv]0�;�\�E"8�8vSpԻr�SYaʢ�V$���\�ª����E�*�]ۙ:bO��G%*��e~tnW�r(�Xs�ӡRo`��TC�e�F�N]�N�W���qO�y��BWO��H%������2d�_�0'�,Kd�ȐH����ԑ�P����(
*s��o<MK�@�,�fƵ"	f� K������g���kvdzD�8^Ղ/�@.ٙ%� ��ɛ�����v���k�	���C��Z�z.1�6���v��)֙6�k�Ȗ�`�BUL����6�^3\8����9c�.���=��1��;�}]Q 42g�2�͉tn�%��p�=�=Y�Lh^����g�REr�P��x��d���k���%�n�d�$b:��|����r��I�E��W���O�	:�$U��i/��I =�Փ�����G1$���Bd�d��x���xu"���=��[��`H0�� �b��/�� �G@������G�뜋���zU!4c��4ߖN ��d��*M�j��K������/z�wp�Ӫտ�
>���o{�4�!��q�qD;-,�&L�
��a�%8���8�����$:#"J��F67����%��d�M̜:#�KOY����㣣��vYe�t�aA���L� �Kmj�G6SJ��m0�n�������~���dѮB�dG���5I��<�����'��d��t�H��D�fK	�uf���sP9�52(!��v��?�ӱ��Y�|���,$��eѧv(�ރW��	X���@���;zH�p��Ax��]�7���w��mv4�	m}�N�e��:uk���쎶U�U�$Tg�K�ȷ�$v�C��q���{}X�;Wz�Cl���xu#�V�c	9�ȓ�~}=y��a���ܑ$�-۽2Wp�`���JΑB}�U�3*���X���k��.��_�B7ʥ���E���>aՇ�w�W��Q�^K����	�K�$�w�;W�&�6m��W�fz�}g^��>�=M�sukL�8��t�,bЖ�!��(�`��0���j@k@Wa�]�5�5t�� �5��D�̰�V��K�B�%�h�U.]V���J�1�l�̱.�&�;]B�pq.�h�,!E�ٱZ��01c�#��GX5oC��Z�\�X�n��l���s�4��3e��SA%X,��Xf�C,�b�h
��i��k�M����jK��z�C�bˍ��7�T9��Hd�����A��4YMr�Ͼy�	K	�~�N��us������Hv]Ȧ�H+w�s{Ux�"*���CH��,hgz���E	=�I�;�d��OOG�%�A�y���Au�D�$}q��)e�����'m�:�=Gn�$�e�3�� K�ݺ�;�6)�(��|ɋ�Jc'wLI�:�$J�@�G�
S���0D6��P��$�d�M�ͫ x�1�����4`��>���ݐSù�.����[- ��cb3��Ի��bS����T� ���UD?l�hɗ��\z��Ǿ#�o6x^��d"��IuP�0���.v�ͷF�\Ue}{��<�w��p������^D�Xso Jd�!��i������ݫ�1�=���KI�݁"��Uj0^!�LT�ĝ���ѽ$y<A3/�b<�b��ՙ�9^����}P��n��y�;�n�*vŊ2�X��LM��>~��>we1�4877�L�r��Ē�����}��vN����)��Ɨ�^%�滗�L�Aٱf�������__�@�����	bntKX��ڄ�->�v�'A������/�u߳����;dn�d�H�HsM�U|���GI����ML�ޣ�[�D��T
}��I6���ެ��A;�S �
{�B����c�L
�_����ž), ��,�Gj\n@w �	va�I���WZmX;��Q���[�X���.=�$�K�jh�I�ޑ$�Gq�~�M�F�z��@H,	{̉f
��D;��8O	@���Y �?Us���wsр�� ����bo���-��W�7��;��͜�:�2	�X�|7C��O���K��	�d��/qk!��yOʔ�����
�����ؔ���E7ޗ��F�o������.*5C�፸���Bq�}hݯZ6 $�MU+����285���6C��$��뙖!toH�H�װK@r�蠅S�ԝ������LɶH�n��A��5�3f�Uk�?�j`S%ꬨ3�!>��Bt�<��8��C;��%����7e7u�w���� |��H�;�L��Ƨ�]S�y�Z��Yth�B�
	�[�[ ͮ�l0]7j�p�j���D����[��(:*��$�}ؒK��s���eT�^Vu��b�>~��W޸Ji�M�+�&�����\�]`�֠�=�$�H�oL�
�E�]��q.8�(xP��-I߶$����wtx��º_ǟͦ+h�m�#1`F�L�-݃�φ�"`�oVd���~�`Y[,C�lKB@�i��of�A �c�<��&�`%"y�N;�F�����nh���w��cţ��no��[���{#���>���͙������fP����y."kEؔ �u�[�H4@Ͻp��kˀ�7���ߝo=�l�ܢ�J��/��!E��N,(pgld2d8l4���&���㾈���d�s���<�` ddy�h�v�ULu찔���{ڡ���]�ɥ��@fD��:�dM����]�h���D�e�!k���8#p~8��8�)�����r|�7d��@'4�g�̂o��ِ���i��	��}ѳ$�t-�D�m��0
 �X��:;�Dn�lYr����}�w�s�������������ù�/
|���%���I$o�xwR@<H+ty �ݝ KH/ݱQ�%C��S`��=�k�q9k3Y��KC8E���IbG?t��o�ۘ���MإOf�"�m��AdǗ�W��Qlqy�����M@St�Cxp���
��y�U=v��U���o��7�Oک>�8���2ʹ"�%�x��>	Y�E�����9���y�t>4�!OO�ͬ�9�~/շ(�2i���፷gJ����)��-�51vk�e�m�L��a�Rㅕ�nn\A�Q �!t�\&�e���"Lg5�ۮ���@Ȓ�1n��	q�"�kqcB�ts��[��R,�s�:�kHfZ��C�k����\��.��-�1�V��kl��vV:F��¼6���a�9�l�ং�]���Ms��sD��}��|{{�Y��rl�ڙ��v2UЕT���ҋeH%a��S>3�z	DK� ��'A��E�`��d�?�Dy����ozA�1w.�q]:L� ���M��Y$�xݧ�*%�c���M�O�[;�H� ^��E
tS4�(mr^q��;sg�����,�D�T�v�UM(�t;P�N�c��;�'��0�K�:�d�{�H'b��O� �A�j��ٿ5e�{�	9�R$H%�wH�	 �ݽ=ްL�A�^���]�ɩ㔡�@w)��Q�͆	7ݐ�S���6":�L�-�ND	%Vt��n�Y����~����XU4e��Mmu5�U1�(��]3t�f]N���?����c��H!f\	b�(n��f�Ww���T�`Is��xf��0��I�d��PX��oTvO?=�Ǫ�����������_>=sN����@��y�����5�3���r�&�j��d�w��vmL�^&��%��h!Ɔ�L�&L��t�Ie����7-�Ad�������kI�f���.� ďy���H$�=��L@#̑��G�37}u����iN��nt�$��}2ċ��mb���P�>~��ғ�v�-�(�O�A� �黎!oZ󸴬�N���6�뮤JD!��S�N�D��7��4~��i�<4������c�W��n� K	[�#Z�5���؝/���ҬD#���[�-.��X��4ƺV3q�9;�E+㒡�@.�-M�_�%� �o/bH,Ww@�7F���wݒ$ċ��bEa���S�t�d�ْi�Jo��Q�H$�A8� �K�ws��h��� �L`�ZǷ���<:H��ذH$��� �����3GUǘ{[O����o��{�K},G¥�.C7w��~jzr�:�9}2��?/;�g3��>��������dɚn�s�K62 �$���L��zK��.^!<9�({�#E��P��nlNz$�Aw$^�
���sǽr��=��-�R<�G��0�9E@��Vʸ�AY����:��8 �z�$
�@>|�`$%gt�L��ج7�z��9n���9q��v�c2�(�j�0s��nҖ#���Sg��!
�)�ʈ1-�6���H o��B�:�	��h����˷��n����U́ ���2�wⴼM�qӀ]_������T׼�D�E7GuP%�Wt��[ď#:��|�Hz=N�	���������C62���$�����c槷�b�O�2	,�zZ@��� ú�5K�g�����W�����	�{r(w�#�jTg��}�C�"��kO��J��c��G��|��gG���{��1�y�w�#�v�|+x�����gq���U�cǽ���ۻ���5y�YL�q&�&I�O[�.b �9��!�;bOQܪcy�}cWh'���I
�dy���X�R�����O8e"QsI(�A�9D�7`���tmن1��C9wa��Uf����)?G�����y=uy�����	$&�^��7�2J��o2{�H����H�������DB��z�H�N!��=�� �����ڀ`� �{"X�vI�fyE�dÉc5g��%QTf5�B',��i=�9��>��OkK�Y�c��$O��d�]aP{�C�x��T�w�M��.=c�יD	7��$�G?rzͬ�\���^$�k@��q�&ǯ�J�F�,�� Cz/&H|��|1ov	�:��l�I��8š�!�Ƨ��3T�s��{��'��}��������9�=g^h���3Ga ���Mf�������Y�'���bKC]���(Ȗ���t��_<�W�z�^Ա� 2��{��n0�[�q�+|�s���θ�{���j������Nn^P캎(X����D�8���X���ֽܗ����0>Fy���8G��}:
��-+��/ʽ�Ԁ���騡�����O��C�3���xh�wX<e�ޢ{�y��z ��6{[�K�Of���M2�����y��3ۻ�Y�>[�d�z�i��m�����f���<䨃���^����w��7ݺ��;��*��i��M��{�'x�@�k�u/*�l���H�'��}���p��/e~�MB�Y�vN�%֫�j YG�p��qa�}�,m�9�ƹ�=�{��v�8����|=G�����|m귫}�zn�ԋ��+�2�RR�.]������S�Z�G)��
I[��yM��N>��U�z����ϟ��{��=5��x��׶��n��*����gw�i{�;�)������`�}K�N�����@y�����$�L޿e�㓁�sA�^h��;���.�ޘ!Gg%� �������)�G��:p���g{���w��K~;���<h���E����!����7�wn�����!#���-�ڶY��o��݃�5���8�؜�_4l�.�&G駹����A���\���h�dURq$��w�R2�j��	9城�o�>�>������O��:뮺�n��î��!�w�2�맜���U>�t�,+*�oW,i�*ŞŮb{r����||}}}}}}~>��]u�]u��\u�]u�駜̳�{��ģ1 ]�$k&hT�\�B�O{��<��>���4֢�L�r%QR֒�RZ�4̂��9}vڸ\��X�9p���9�!��B�����8r(�"��+�r��B�r�.k�¢.y������ox�^d/� Q(UQ��((�(�ډY��XJ����$��r�,ɥg�NȞEʼ�H¹W"�3��fr�$b2���Ȑ�E��J�%p洹Ad�$�����d���+��<u$�'l�'Iy�)�*����;��(z�Dh������(��ZӬ�J���N�ԫ�M�wi�*;TI;��$�"��A�߮=���;4!F)�����M�,ӠЫ�jK}y�7yD��+�����Ӛ�`�X1phhK[X%�1��`�7m��]���e[�)�@�c�.`��mmj�fK+�,���E	h֘u6��&β�Cj�m(�@��S6�r9��t��-�	�Ə+���YA4HV9���1Ypj`�fq5��`S.���2�c�/0.��,��)�s�����[�-pVYB��;J�1���h�^1���H����֘�&i6��e�A��a70니�v�f3V�Mq��h�D�0�%�5	���M6�h��
Y��u�Y]t)0�5�u�C���m���X.������B½u�ˇ[-�ַJJ9��Lkt�]PF��L�n���ggh�\[̢�T�4tcU�R��$�·7^�xl�9eq��`Զ�l���ݠ�ᣊ��D�͂���tں�64h��Kv����&��)�Ü�#E����aF-����r�Y�)j)rݣ`�f�KX+	t��vWB&u�"�RgYb�a �{i���LԲ�]5�l�mb�Ëfm��0�ĺk�2vHݍ�6�RQ��4l�I���N	tH`��&nx-3	ln��Q���XP��h`����]R���Mra�c�B��]�l͵�/q[n3P{,yq/V4����&�7�[@�YZ�$]��1wΗT��.��X��ʐeu�^J������E��.B��X�#6jJ,�\6&���.m"���-/*B݊��j��V��*���홬�ŮS��e8upgF�΃\7��vԤM�%m�����V3nV:!v*`KDf�R�V�X5e�0�EE��ak]w+�,E�:��DJi���]s4@J�<�&Aq�Q*�h�9Q�r%fv`�ƶ��Ɔ0Y�� �-�n*ƭ��c1��3��p�3�i� `:���	OW1ϓr�n�	c����ή�:����Ԯ5��2��۪�)%���<|��&Ւݑ��c�b�?g~w�g^���ѻ;JK���n4�j!x�6T���5�+�6�X[Bae�imʮ��c�)2fU�)(˩�ecYl��&V87��g��ԗ,��E�45rٵW-���p,�����c�:�5�t�(�V[��42��tͦ�hRSi��c\���P�x ����Fn�Unk+T.N����2�#�m���vLF\"Ʈ��kc4�z���2��(7k!Xj�����d��6"���5�"k�_^B��`���0��>O�k�~1L{cbI%� 6;�A�A�\&�uV*��f��"�b��&Phgv��V�"
��M��lJwE�;q\�a4� �^z�~�i#����H���n��vHs��JDBJ �.=�"���]�d	 Yy��m�,(:C�\L�(gNɗDl������@x�Pu
*��~�[2�)C��X�7�Z�����T��:v8¯^�m/:��i^̸�	>9%�<xr�
́����U��y���gH[��KltI�>�;�|��=��彩�e����FrW<��3Z�46�q6��"�SK\�	��Yz��{�@7���s^� U1`X�f�Jm=d��BP�в�u��j\KT���xE�DbG��엩C=��;�^f:~����e�I���N�E���������?��]����Տo����l=��[�ܼ����t�����2cYQd�|��'̗F�$[�N�OK���=�F��E?�"Pt�
�h��ı��X�@'�����eV�&��{��i��['b�H�c��|�)C��ID�s�F!�	ǻ%��4�L�vH�d��@vAgwEFI%�f_�:k5�=��j����<A(:�()�ӄggD��Q��^Z�q��3q���?�D���H"���6'����wʅ"��%�5A��F��p��a�mi�Зa���%�#���Jwx��{��FD��ȒA�3��UP+qt�zVvQ���je茑2���V*�$��}��ٞd��w��eR���Kg�hP$���P�uX�mG���$�����D#a5���H����$��=��$�X�o�n��㾀u]�M�W��v��R�X��7Ğ�J��o��ͥ�:���m��.a�jNI,�����gb�5Pgb����ȐK��2V���(:J�[�^��%x\whnؐn��Q���ݙ-�ۯWd��D��X��G1�s�v�P�"Q$xl�L� �f���&��zh {��$�K5v��	<���iu�#ǃ�2>;䧞�5s%F���1q��Z\�ܙc���	v��;�9��P �B����<� srbAb:�Ge��/ۻv4�@#}�"X�o��	}R��]��:���Y3��%��ϝ�lW��}�#s��<���O�2�D��v����'ö�*�$�P[-'��C��[8�v��v��т� Z�ft�%�2�{����ݼ"��Ø�c�s��4i���I��dI��@An���c��x�F��O�����>U�#�H1���Sc����y�ίt�>�?�ˮ�H�%������N_^�,l�st�j�<8����bǁ����J��V�%I@��y��-���s�c���h��骪"�2����:Rˈ�=S�UT`v���ˊSi6G�&GW2�����\�ivƃ���/ߟ���l~����|�\wL�ދ� �Kڿ�c��c�`,m�%��!2cܳ����x� �?VȠr�������J�y��	a�twL�H$�LǹE5eW��{4N���$���uX�e�"H%�w�"�#2�����0nX[�h�%��6Zh�ٳ��s�Ȩc�3��3+A�"�V߉=�2$��V�y	��N�1`;t&�d���sxx�a�H�=��/�cX�~�SܫOf�$n���KFǺ�$FoL�gP�1�S�U�o{����8'ozX�@q�jj���{�%�c��������c�&��n�,%eC�� �����LV�HF�}�9�g/;�׭e���1Aۍ fP\J%��I�a�h�A��vטcU��A!u ����iV�Q�e���j2�E��YM��Dj�]]K�rˌ;��3é��	b�Q�c8���5fy��xkjd5i�G�ƶ��9� �i��.٪��m��f�gJm���{:���	��yZ�.� �l��A���U:�t&�c�&��ğ,�6�.��PB�¡4��V�a��	V�s�5�]��r�BD��WtJ������̂q��1�$���2_�P%jʓ>��-����H���yBq�(�R=��&A �{So _�:��u�s��J�����F����ΐ�U����lc���@w�s��F�>�����ϐӇ��}�.B�耛,�'��C�ٰ�:r]�	%;�J*�~�W����Oz%�c�w�$���{�*-{���<��P$��/�	Ct��-�DOL�A |��1�{�'{r�P$��� �u�e�.8��bMP~oA���t������mb���iy�!XMr]!�uͮ������m\���q��:j$�{v$�Kk�̃��"��jLHՏ�	b[��6��o�����z��ܛ�;����(��y;Q��fϹ�N��R��n�NZ�63�_	�]�=�xn�=Cԥ`�qB��!�tfS��UXg�����P�����1co�I ���2I���(_wd�w���Qm���v�P�b%M���`�[��(�&7ڻ���I��%�_��5�i�Jr�᪁S�������`�o;�Hv+#�dKVGu�:ǟn8WYN樂���%=^�y��$���5�����V���Hl�2��#�"�d��;^Bs�j����@B�D�rl�]m���n4ˈ�URĖ��,�t��,�����x1DM��0�##��zD�ƞ�d%�wKuϫ�v�{�ķe�
jd26!�O�{r�<@N�*��DĒu��]���e��)1 C�M���7���H������g��WPA9J
 �Ǧh���pGo����ߖj�w��	ʺ��O#��N�wڍ|H�ӻ6��p�����sϽz�NћMm��܌Q���`��T]/_���"�!�&�}��d�u�@�_��I/�b����\D:�U�gM�����\���Ĳ��H%�s��OKϏ5�UJz<n�(rS�@��D��w�܁���(�:�^�H}��0�['2[����}��}�.�̇'e)x6���[6�H�pms����եb&�]t6���u:Q��w���a(2��9SN�$:��$�I����>6���-�s�d�t\�P�j�
���#'�#@$&\#�A��w{���(k�����"A�S��*�כ�]�ی��3���*��"���bI̖�tH$d�����*� ��H�I�Α!�[ ���z��� ��};륚İ5>�ı:�r�Sĝ���&f븐z�T��b'*�ʞ�����ws���y�@.l�r+�<E�G�U����*"V��(@���Ǟ!�<�X�-l��O�#�hzv\�ws��P+��,I�v�P�k�}�9�S��:�y�=��"R$���	�~}�|���;�}�)���ٚj����&�\�nܩ�4)��a�����U�CJ'~y����ڔ�C�In1>G���EOGlIǺ�l֎���dI �w H��Op�xs	EP)�bO��w�����=�<�]"A'�����l\���������	��c��~�~k�
���#4��b�@'=;2%�Mݯ�~�C0�) ���޾ɜA��Ռ�Y��X��"G�WC�t�ꮺ^��v{��$@�̙$tq{�Α����J�zd�uȩ�����a܏F���lK�!EQb[{fdy�G��ZA���&��fY��R�9���w��5
/���3�)�]�2��L��I}��;..L>�ww�u����U��=�{V����g����y�w�'�y>��Tcfs���i�jU��[�M*�b�e�K�[�Z,�6nQ��XKIZG"gnR��s���0�cj��Z@l��G3;�慣5�k����1�+e��lG�]��s����s��\[k�#n�0�bxL��!P����l��X��d�_��U�	zWA���WL˂&����!��A��q�͍���d��cB[������uq�JL�&@�6�h�,ک]b�,��Ŭ,��4�hQa��>���;�@."H�.dI6��g6�O2D�~�2Ɩ�3��e�u�L�,a��ۙ����ܔ��G7�Ԩ��ͳ��+obA#� P}�Y"��*A,T�{Ӑ�{�f�����(�ØJ'O�"H$�e�8,r+�я����KP���Hz~�$���7���9H��2jF�䕝`o��1���1,�H ��H=ۑ!�̽nQ׹5~>�$���i"=�W+	�
wbx^c`�GD��:�zb}�q�=uD�B��RH9��5�C�ű�si�G#1n�EϠ�bڦ4���׵�j� ���NasʻEt��{��YpW>ڀ � �,�A&@ͽ�#tn�3����e���!+3wxp\D:���/�I�gN?r�3�����h������S����� ���]Ӆ���C�稃��w3=@��
�m���6qg�]���	E�C:�c�"YSt����zgY ��w�����/㒶x9�x�b�gK�$/�"I�:���^���l��R5 N���%�=~O�xs	BE㶣u<C��x1��z�'#���Gg�N��b�
߱	6�܁PМ�j�t̰$��y3��ǁ�b�|���ȐAc�D�:������IO�5)����H� b��5#�D�y�0Bl5ujL�-��ë	q����;�(��w;�A �&����z�z�]�٥��Ҥ�÷fd2�[ ���S{��H�?�wp��W;q��\�$��y�LI�`H3��<q_9�FfC8}�!N���q�mg�� �+��$Aѡ�z�c�CŨ�o����Q�ɯ{'o�p��S��|�lZ�*�������>�"�k\��:QG$�s���$9ۛ����E��.����;���Cw�*��݈tk�����N����\8/{� ���A��`ܾ<��E���q�B���=/�A9
�s�.�h�7����!�~z�>���=Re�h��P^��U�}M �/f���q�X���9ᛝ����|ICl�;�pp�-���R���5�w@��>�-u��	]��,��\N��0v�����m��z>�S�յ�5���^����i�R4�{Fd��!۩���_;�.�ko�OgCz�v��E����`��u���zZ�����[���_vO/^������^s���eg�j�h��:B�9��s����xs�}*���ϧ��$�`Y���V[�_���l,>���e�<�5���<w�d-u<�|��ܞ���}�}�_����ѡ=�R@>�y�!"�75�c~ć뗐�Y$/Y6��w���x2�^_q>�G�+�i��
>�6E��̶P׹b��}���a��yz^�*װ]�}��9���V�Kb�����w{�x�l�ģ�hyJ\�;ӷJ��_l�J�2Â�D1�R^��v���,s#ޘ�+�������r��}� �۲z�����.q]�	}P��9����^h��Ì_�}E����ш�V�%�鐐� cO��f�;��z�иH$
�����Q!�I/ӕ��+5uݕ���^�i#4�)+ �,7`�*t��Co��������o�������㣮�뮺�㮸뮿�����QL�H��p��$���VUQ�:�<�:�M5VY��fYdp�����||}}}}}}~?u�]u�_u�]u�^^����b�&ӈPW4H�%EhQ_��}�/K2����#8r
���ZV����!�O]ЬbYaR�����B�b�8j����4�wwID��J.|����Ȓ�8��ʤ�y�v��/:Z��Ш���ZKR�MJYϨ�w%��VJR"�$/G|�DUz'��}*4��]$I��	��]'GI���f�C�[,��WV�D�)V��""q�r�u�����K3��Ȕ�2tNp;�G(S�&W�Т����֚
�M<���=����*�EO�x�\�k%E���5B��\��L��R��u��UB�!g�.Nb�E��9���hb����-��0�̉,^�fO�G[�N '0�LTs�`=���O��D�A#�����q�V�u)̲Kg��A"=�^�����e�BI'�$,���{Q�`����Ly�X�LL��N>��vu���s�^>v���m�ja�[�s�E��#tƅ�0雬ѮB5�qN�����>tJne�@����Td,�GoPX�<��dX}9�����y�AvL��fe�����	ܘa�P��%�]m眛ȓ';.��2�v�$���$�5�8�$��h'���(1�����(�@�{#�$�~~�E��*sGU�g���$���1����A!���;���C���뒯����0�!�I)�.0ղN�ީN,Ftk��T���j�����������bL���o/\x�f󞶄6�A�ْ�����[��^(i��{��1bǌ2d�3B>�r�@Na��.��(�o��Otg=��O����$�u��=�� �ݝ��;�a#g�Ѝ���iMPB`ʢAe�%롙v��¶ր�9�jA��u�΃�9�����H�	ᔑ��a��[`� �OCky�4��m7����8(�:9�� ߄�Bs����(�<�|�,���2@ ꭊ�=�{=�s5�.6�0��=p�y��� �uE��n4ce�p�>||2e���{��$z�O� �B��=�f=��	b�o҉$���jj	��M<��Dn�֏�d�{P���q�k�D�2L��{����-y�Y+��{;�A��ٛk&��{/���ϑ�܌����4o�{٪d�|�v~�<�����:���P�?���8x�5 ��{�i�Χ�w���3�J}-Bf�ۅ�l\�
�ׅN&��M���L6�P^K�%ζ3[4ʗ[�95)Pܕ�6%��Ÿ��1��7M�Df�xP�J`C.���u�`64�dYI��Ռ�\m�[c�:fp�n�9�H���q%ط�y$5�)7.M��a�ɵyN:���q.R�B���s��5�sq���j�J�M�ˉ���?����3Z�f��T�2]ex�
Q�+SMYc[��AHR���S�	�;�c|�m�Q$��H�I�fG2�a�|4@>̨�/�fX��up΂xs	9jv��iF��Jo6$�K�;V�\�Mg:%��$���+q�*���J]:�l��x�*C��jYK
�ɒ	cѦ</�j���$�׉$���d�����xI���9���v�y�.@r�zX�%�^� A�칢A#v#�E򕛾Н�b�fA!ꏂw�L�`S�G�>�X�o��B�%�s�Q�tQkƀ�wp�
칐��؎2zgi�+����ⷼ%�Yh�UV%���!i�릶����ڴ�!q[3R��
ׅ6`�XQI�R3�m��h�i���%�b��%�4�BY 3�8�w��[����l�zZA��̐* �C��r�⩁ק�C��v�s��藑�O���`��'<�44��4:M����~�ޒ��Z�K�׼g���3k{Y8��OW9DY��H'���kb˫� �d��K�7�T5�d�pMv�q���|�aEK��W.��N�BOT]��A��$���֘��U��6�����& �ӓ �d��#��hGGJP�h��`�Q|�_?��Z���Γ�$��;-,k{��[�������%w2�4�&�%���N1T
ܘĞ�ؐz(�/_C�{c�3m�6��$���i���SP�~��E��7`i��ԙJ��e��e�.�R]4��3al4�rL����=RS�t�9����$�A쎉bK��J�;��1��k�z8�6Yy�@'2.D�&}�eQ
��P�C��Z}'�ı�O\�so0$��"I$gwL�A�M�v��q�����i8�/��q�P���tH$�z�%�`I{�q�N{I�6j.�\W�)���=M�=�Z5k���R�����*ҷ��5I�_�b�g��2�<�x�ٽ��gki�}$��2b�{�$ȸFwtJd�:]=��'P!'�.��q��"o��1���K!�/*��K��B���U@�� %����M��	���1�*��t�$;$ɗE�N��G�x���ع0�Ww�$� :�����O�p�H���:p/9t�A��"�x\J%s�V�3.��ť�d���&��g�-��\��D$��s�1Ow	���H�m��F�ʭ��8Y�#C^]РL$2��I
��T�P)��P><��c�Ί�<��	d��{�(�y� I]�'�jd]w���{H�%���R*����ȱ ��O5"N��vVz����PH%��&A$�~Ȗ���S�E҇���"u��{d���.��S@H&��d��{�?�(:����W7.+ۂ)��O�sl(ܼy�-k�M�z�4.�^�d�R�$�ڼ���[D�r���l�r�%��p����X��GD�ɑ^R�9�.�BN�h��M+R/:��"���
�	bX��e��$�Vi�/����κ����]5���r��tX�̪�6��,�s�1� K�,���O���2����b@+o%��A,��D�3���D��"�>hd�./���[�.6"p`9��莉$��~�*u�[e�\���4ɒ$,�>d�1K��]��Oژ�zO#/e��0*�8�܆ԛȄ�c�dU��$y��9<��H/��<ł��A��$����/��DB����XQ
���b���� �!L� I�]ٕ��o�ءj����d�x�r�B.�<U=�H$�_D��{��2=�����e̒	[�"e�C{�e��/;�O<u90�{�����'�e"��M� ���ɂ;7c�=44Fvy���.^w hw��Щ�f�m�b~��s���c��m�nW�]"ii���E��K��#.o6Ϋ
J��0	5��H�D3n&Rr0��j,�^Z�Kr�K�	s���h���ִX�Τm"��e�ƌYq*ۈL<l5�Ŷ��͐�ͷ[���Ԓ����w:��c�H��51�F��&2�� 46�[��� ���s��f��K��XP�k���|}q<���*9�\it�聛u�Qڷ�����W[J�Q�%9��iw#�]@��a�(��,Se�bk:%��{��JO��׈���,HW�"I�ą);pQ�O�d��kz^�D��s�xǗ��Ks{�F2L������{�7�䗲gLG�ёQ��1	ܘ	T�z$�/�b@$]c&}k� ��,��@���MI�i��R�
c�u��jQ���F�U��Je��4�K�u������@*k�I!��o�x��*"R�{�7�����)�#^�D�K��2A+��Z��dz�u{j+�jt�Y<;�Bi��k�f�el� �����Yqh�4�0�o������"NID@�5�Kd�.6$�N3�?4���{�yn���$��ɐ	f4'lb�$��'^e��mT����;4��Pv9���m�Go��ݔnr>��ջN����|����}���ٶ�޷��߯v7w2�)N�o�-���,Z�́��nd	%���@����7J\�t�"�E�bv�i
:�v/�,=�虙�
��栎�􂓛�K������$���*�{݅.�^�0�y�L�z�[�z�2
/���t�:�z7����:��I��$�zdO�U�)sE1�ǥ��$�vĀf_�~<�xxI$�D&A�66��xɗ$��"����"A=S=}��9�����j��"Fљ)������@ƬtM%̺n���j�G��&" ��N;���ȦH��-$�B�t�8��=%�Ʃ{�&�*2d	%�+�&y�<�tS�QQ:OD8���P1S$��zf*)�Y"FF��K���[y�GdC�bA͸�"-��bDю	�X��	=�lI�~�&��b
s�׽��|{�X!\�D/z�#�y���L����M�[ˆ�׋��L�Y�fE���:[�b����򶽛��T�iH<�ŋKLtO �k�#�1w�,Mo���^	F�s�JΌ]�~�tj��vv�X�Unȶ��#x��Df�]�Lև�� 9�r�7��.�;�
h }����T nc�{�z�4xs$��GKK��thS���K�N����:��|(�@v�t������Sb.Z��-��<���Pō�mݘs��O� �D9�Í�zd� �݁d���1���!G�u�;���$�_L��d��Fx�/!H�>�L�A~�5��Ż~��#�2/��$k��I��<�4��\���F:)��(��aI�'Θ�@'��:$Lg]?�^=��_F�/��Ē3�	&�pN0�]@�����P|~	ev�mwlI �	l�ɒ	]����c���ĩ�Wp�����Hx(�/,��9�3�Zix��g}�_���[�N���d�뺣^���[�g��,X�d�]�9�ΤS�x%i��=6ԁb�s-*����H��,I�̉ �J��֩���m�ӿO���X\��R���f�v��,�1���2�T�Lk�s�am��?5K���K��%�g�@$��C��2������%�;�-,H��fX��	k�"��0$kx+鸐v"�#����Q��ćk��X�+��A>��y׃�Ŀh�K�5`0^"<B�[��{�D�A�Dm�:0������Iln��H$�d��pa�*#�e�сD���6����H`_/�@ %�oH���Z��{p�$'�3$�ό�O���$�=��2X�+�  �FU���n�VEQ&Y(�\�������'����1ڊ�����"?��7����*�(�(���	p:���U0a!�@!	Qa�Qa�Qa�Qa�Ea��0BTXe�XaE�TXaE�TXeE�TXd�%E�TXaE�XaE�XeE�XeE�XBa�!��VXea��Xea	Xe!�!��VXaa��VXBVX`a���Xea��V��Xe!��Xaa����VXe!��Xea��@�%a��Xaa��Xea��%a��@�VX`a��Xe3���y�1Xaa��BXea��XBXea��VXa`a��V��aa��VXaa�!��!a��Xea��VXea��%a��Xaaa��Xaa	Xd`a��VXaa��VXXdea�!��VXea����Xea�!��Vaa��!fP@C�A� eD aD eD e d dD `D eP eD:�x`` dA!��P��D�Ha!�eQ a a!�^!0hd8�qHQH`�R�AHe!�D���XaQ!���!���Ha `!�dT!����P��P�!�����P���A� eP9�qTTTTDTTy��P dP eP `d�`	Q0Q`aE��VPXQs qQa�Qa�Qa�VEa�Qa�W�]���אa�~_��
� (��
�2?C>7���{�� ?@�?���Ԥ���h�?�F�������N8��������w����"�(��?�/�����DQ�RE����`��0���K�����H4UW��� ��E���,���x����О�~��?P���0��# 	  P�B � � L ���(�)"�
�(HBBH2����+"!*H�H*� �*ȈH��(JJ$��H@ �B�H ��BB �*!
BH��� �$������"!@(P� !H ��(���`����8?j�(#H �@ B�����? ��������(>���A�?y��}��@�(��p?_�������?�ps���G���c��9?'�g�
���~�?�~����=�Q_�E�O�C�!����?����E���x� *+�@c��z`�+�ӱ�?��z�~=�'��''��vpA��*�+~'�a���?D?��� �(�����`��xo���i�;�?p0? �����~�QEt�?y�S���
����:�9=�OP�)1~~����`z���O�����>��BO?.�TQ^���O�1� ~^A����~�M���
(��,}r��"����o�O�P�?4���d�Mg��P,f�A@��̟\��o��                           (    (    �  �R� >��
HH+F�@�   h  � �� h
�� M  �     �                                        �L S 4@�+4*� �@�3� ́@d$b�g ������@�<   ���1��� �4HU�23JFB��a�3�B�<�� �ХCt��\��\���Х�C�
�.@ (�   �        �T*�e�q��s4�9���aB�:ʸƂ���� �U
�c4�hR��4��P��(T�j�wR� � :(d� �@Q{��<   0^y�z9�rQe� s��K��v+NA�[92*UY����� �H�=�5���ԡ��қ��hR0Q% ��  �       <�������.Z�Dm���B�jTT�� �v�+��a
���73Gk6.n��� ��f�tª�w�(��x  :�1J�1�릃 �t�d����#V���F���[p .�U�s9ى.7]�73s*�qt�R��UP ��  �        <��N�4-��Nm�73s	��ݩ�3��v�];Xi�7]��hq���f�p .�j�\�u���]�`@D� @���m�J�����c��GYqj�4�q���۝�IVcs�uU%p �+�[��Mcs���Nv���ΐ
�$�^   �        � ̀�d�ҁ��BE�R�  ,� ۡ@���P*� �*�
�T �� :�����H�iT t8�0��4P͊�M =� `Gv ��C�r�RFlx��4�MC ����4Ԥ��hL�$ƈi�h  "{TJR   j��&T�A�F�i �)J��F ĪJj�H�2k��$Y �c�E�IO`L���IMHB!!�B�� IO��$ I�=���;P_��C��L�ڻ��m�&�p�X$��,N�&�sĚ͕�;�1!��8���P��\�i�1���x�t����`F73��`W��� �w&��NHFo�\Q��=��L�]��L9��E@m�a�����x����48R�ɕ��W�Z����y���s��F!O2мR2Z�Q��K�R˘Դ�&wӏ>��o�Ƿ}ьT掊w18�f��ì&�W{D�b���ʁ���Ť����,�f�$��WgL�0�)����JgQ���e��9�I�Ӳ��L<@�]�x��A��*�].��@i��͑���xVq�H7��ҷd[ڛA���V\�P���s4��ዱ�[r�ζv��wqb9E�7)(Έ9��_{[�qIKT�ge�"�N��I�X�����ݩ��`�ĆX�z+�+ߛ���0��:�-�nwL�����X-9�*�����ol˸fK�5�'8�Ya�Ԅ3^[�zg;���,����hۧ[��K���3:��gn�4e�k.���D�Dʻ ��t��d���xw7s�u��a���;sx[^�L�+��g��P*�;�cݧ$E�-��x����m�0A; �����X��ޒ������x��9N�h���۷��Sz��X�0�խD�%f�g�����U�H��QK�^����o��ි&�i�8�+K���9�_M��#�g@�Lf�0&P�gnpػT�u��np�M�"+��P�A�:^����j/� v�����܄^ȴ1��:�|�Y�a��r����0�@�8����ۋT�h����t/���8�Ɇl�
׊�ۦ����2��.Ӗr�4��iz�v�Ա�έ��؊�uՒ�ݗ#˽��{���[�C�BF9Q��"3C�z]-����� ��u��s�ylKM�X=�0��pby"�մ�޳��%��Ȭ��k&����AȊ)�Ճ9�]�fL��g:���J:NC��@���o-��lTdYZ�nM�޺����X�0������Y�f���~ n�7f��fQ��)��t�"i�J�k�e��K�n��m�7�=�5A�Z�Q��;8��.olԖU�Xt5�,�~X..�Ir�5��9�-4�4��!�gE�gt]�G��ob���7W2Q�Ҩ��iM?�X��L�n1�Nw*]7��y��pss���5�,�Y���!�/n�x�܈�W�ٮ� _��Z3TrpQ��mN��]��L�v���:�4\\(Nh��q��qܪa�l9M�+�����k���8�Vr;��� �=͋h�x���V��2V����^ִ��B��3�T6����9�K��pt9y��7��W{&pevwcE.��
��sC)��xnvӜi��J|od�d�$Fs8�d������<�	[���G��w��!.�+��f��+m����Y^�lh3@�\�L��|�K�� �k�}��mh�N� 囡t^Ә"hS��]x����w^��$�O���"Y�7���M0]x��P�]ȕ �F�i��B�o�3r��s*�}2,-��:5+������H������ǖ����w����ɽK�%go`�5���gn�������Ͱ�Y)^C�F�Fk���n��<��ں�'!\�u�:�Ҝt���g-h���n����)s�ŝ�&˰568��9�tjv�>�
3w��=o<tN�0�{��^6I�&]�Y�UνJE<yy�;{��)��^��:�n<��l��rxv�Ʒ�B��.cepd�#�bn��4�t�ON���Y��UY�B�N]�.!΀9^��$�B%5��e�`�_.Pt�Os]z�!%Sf,{!\�1�.]0�����z���i���2��='+jݱ�&u�ۗ�P�*sr��u�4���ی�8��q���O�\��En<c'�T��5�^��
�"�UBM�8��������ػ-:�Z�������w;�*�G��iu�Y�E���(� �u6N�	uon1��u�zn+�@��l�-�$^z5懰Sģ1���V+�`û؇*0F���jͅf��`{K�s�H�Ɉ�vO^�Q�Y������u�CoY
s=��V��6�g��kgi�i����9q�����PJ�5"ӫz��Smn��Ձv� ����۱9<Ҩ��ö������ �t�l���^�E<c���tW�M�i�՜��,�P=M�ˣ��8���V���x7/h�kwn��&��T�R���C��^X7]�%���s����.$k�|3xwB�t�K��s����L�����Zv���^�n5Pf�%�bSk;O>��N{�Q�N�䝣��Ţww#��wn+ݿ 3X������Z�nov��O[��Y�8�Y[����c�$Uˎ��A�c��dEU��wt��<+���`��s�`3^�b�{�0��xC�{N�ɳ�QEM8ˈn��lH�fFPR�_7{��i#n�u��&�M��S�)a�״Ừ�Ba��]�4��X(�SaI��ӯx�+�n+D%qUl�y�k\O ���+:�q�)��A��<N>G��ff�ݧ9��u��s��X�Wwvߦ�M��[�.���8�[;X�<�o(l��wO�:��솛�����z�;"��I-�!�'(��oF�f�2��6^-�C���D��T�G���;q�F<�'l��ͼ)�x�� Ύ�61���o<F�՛�|���y���ᕫ�21F�X0ۉ�]�"�2����w��7~��FN�6����wU�Xܫ���s&K�ǳ)���{q�r���pü�J�b�#,���˦���U�D�ٽ�%��eņ�N�'f�E=���-y���|�y§'��j��G���I��^'��Z����Gڂ�k�DĞv�n��[:퐬Z�!'2E���������ނ��8��}��ٴf���9-�$��������"H�Ш'ZD�#�JyM]�%�K�к��m<���8s�������1��j�ᯜ6��X���,Q�v��uA�
�٫I�;!:4$��8��n��S�,[�����A�ӎM��kzP�T���;��]���%���)r�f��9ͣ[��GR/]��.�fm����h�'uܙ��p(s���w��N,���W�ݗys
���(��K�m� |y��7�Eܟ�K��G��Ƴ���wJ�7j�f͘Ʉ��r��F� �����b�hs4n [�X܊�\F��1����$vp�ݹ��(y�]P���A7i�����Ο"^e�f�Zu˽�.��%٠۸���G�TN���Fx9��"��U�o-o���4l��z��х�q��jۑ�!4�zBH�̈t�����Vf�żäv)z^g�-��<�#�T^Ճ�w�cY(���K���Q��wb�or��`|'���k˫~#9��`�8�j#ٱ����o'3����6��[���k���d�4h˂!�U�����ڶf�o��caM^��e$��f�M����[��L�����s��@N�oo�ƺ��չ��9�R�M _
�y�N��/�^�2o��a��m�Wq ��	�&�q������3�6]7�(E-����ˊǥ�d��!?h�7T{����㛮��ēӟq�M�4n�ѐ�Sr��p��P��.��l�".�pc{7��t�3�J��%���ddwv!�����\�r�9��y)��`�;U�r�����o�G&��8��0�A���q����r�ى��?N�[�u8j�$�yF����7�T��i#ږ�"/Vh	�J�;=̜��r�Z�
T��4�ޜ@]�V��6�.���V�V,�62{PpO�٦a��'zD�^5i���ѡS��A�>�J�0j���+ݽ��nYv��6V��*e��8,.Pfw\#��G�A����^���Gv��	G��tk��M1vͽ3~{��������6G�J���ћȎ�[Em��/�^{���R�[��mŕ��b��G�"(�S#�z$2��$�L<ڥ�{]4`p���w�C���BY�E�>ٝ��L�{iC�I�G����b���,�t��Ð�<��M�t;�v�qtΟ�׻4���y��:*�vv�/�2�7零-�/n�f��'Q���k�>��%O[o��L3��8p՝��2�z�p�@3��7\x�*o	ۻp����S�iPS��Wi�;rh�> ܘ3Cg�S۳�1�'Z��"d�B������.;�Q�Mc�O�8yr��^��8bwz.���XK
�3b�gKO� t��mz�j��b��Txp��I��wk�l���s��X�t�U��u���E˹U�_�b{�܎.�H��������Ǵ���/p?%�g�u���9�� [�6�n�f��Q�qz���ڻ�f�����'�^;��+T��X�;9�*�>ȵ\{2vr�v�������'f���u�sn�7��n#��!4�5ש��+.�G����3�����Nx�*��5�;n����0C�[��I�mߑrA��������%�om��"0,Wr`�9N݊���Z����i���<;I� O����6u�[��u�e����;v�Ub��3���M����NӚ6,�Xz4�.�xs�=��x&�m���	V���j�V�x���x�9*z����{�#˔4�MIs�g�21wn!������t���n�^L�0+� *�0j��;v��nn�ڹ���,̓�k	�ao X���8M3\�L(f�?�kg�ޕua�e�w����8~,ΏF�����z�y��Q���ӵHvFb�!X15�fww$ ���U���%�9���<�rC��pf��[�5�>�=5q�.]�۴����ʧ`�3�f觐�l�s��t���'u�g���l:�G0���)jg-ޘ�wk$!�b�TP�3yʳ����7V�?<�|n��|c9۴j��p+�jвp����1K�Ȩ�v�^���G\�_�H=����Os��t���m�Gp�Ӓ䳢��-�f�a�.�D�ϐǇs�&�oo]7k&�B�jP���qr���ǜy@ ��#�v�LO��כ�#z�-f�8�V��퇶�X�����p��e��w������M\@��Jpʵqq��²���5��rBm�7[��� �R%�ދ�W9��jó��'���i[ɝeGP
v��BW Mf�ø԰�γm
\�PS�-c6�ݮv�&{;��yC������:՛�E�gp�9��{�M�� �]�@.���S��й;hu�h.�Ǟ��
׼1��$�m}��9�z��7�u�&.��R#9�R��]٤GӦ�:X��u;��G5�p,웻�A�2��KREE:oV��Z�2�=�ӡs�Mw
���̰��]�7R��۫Z������4�!�����a����\w���Z�;N��WĪ�rdx�u�Vv����	Γ$�������R�����ޔ6�,hNy�����8oU��v��<8ņX�g��9�8)��V��í�� �����N}B�F���I<sL��N�����{�lG^ӜT��>|*㧸�Y�u�yx
X5��7��	S�cv�ʹ�E8t,U���
���E���*��N�pMـg ��|�*���f�y���L����Ji���n9NM��1��p.(�6ۃ�ݻ��+�
}'=8��x�vp�7��
�bɕ����@�������.Ew�>ewP�t�x�h#xE�]��\�t�1�V�zr/�׬t��h!��$NÌj/�U��dG9�n��fwS̖f�0��fs*�ݸg|��u�b<23�Z}�'�\=�.6�L�
]��r#���
.�5��W7d@�R��.;9U��}|�>��CL��w�;�oV��|�vo�CU&�9�o�_,���Gr1�.ݲ��u9V�!����je}�n'���^�n9
Bӛ��
q�]؟1��C��f�O]��(��sWVrQ[4��	MFfJH��ɥ�M\{d�����4>B������G�ڻp�oݣsvp=��m\�d��%�x����Y�,;��b-�P����9n=�����мE�glL�f���Y�v�7''�Z�,A�f(��nM��B���N��(����5�wx�E�v���&J�,�gn��,�(ܩ�+�F�KsF�co����R=��8�;7S�09�n�[[�k�v�^��u,���k�r��, �n��K�ݽ����l���nJ�xe�1��>��4<&�����@;Yŏ
L��HEҍ��/tCe��kL��]VY�9e�!s�os�ޫ6n<2�������c�s��#ڲ�R�e�rM��{��YS=���l��m��|pv�/�ń��*+�K��n�;0h74��(���(�h���eB������8Ej�[.Ԟͮt<�Q�5����q���6{R�o*z�-��M�w�MFVw�*��6��)ԥ�n�I���ܽø���f��������N�n����ݧur�eo�~�H@=H
Hd�`B,)� B�$��HT����@�R�IHE����R@P�
��	�� E�XHAd���	 ��������)$"�)�E` ����$BB,R@+ @���$�!�(@YE�I Y$
B(HT���+�J�
�$
�$�$"�"�H�BAI
���$*V"�E "�*���J�I	P�T$�H���@!X T�, ��(�d ��BH�F�		Y�(@@P�P�a  %d �� �!X@���
� I
�$�J�� ,!$�� �B�����g�[��i泛�����r��R3����o�����[��L@����tYk�ÜM����wn���чxxe�;��c�#����l�#7�p�mt7�:�_n�=lrY�FV��Hm��6DūPwF��q,���j�!wA�XŮ�2h^\�h[2��oOu*u�������ǝ�ٜsr�y���͵u����75t}��h(��A옼T�s^*�@���`����D�T
0�I���|�ӽ�S�x��L�N���g���t܌�7�:��Hč���}��\�vs]�1��d:FsUMm走"S.���3���������hq:m�{mNb"0T��z�a��7g*7.�^��$ZdXwz$�5�������]CT��*yݽZ+V���p=y�؞"0Ż���Yn�}-J�G���r� �3üG�7���̇��/o���Obe�(�N�5E-�uG<Q�/w�_6PӾ.��8{�lRgw.��zex���۽ø�y���p�/˻�{/a�\�sKi�䞳;Np�K��-�殾$��v릟d��}�zh���3p�Ś�xk�����zJߗ��h�D�}eo�j����em#W;^���I�>��}6>ީ��K��L8#�|/����;t�h͋WeI�9�O�c��;ý���<�qnsW���<�ސ{�{��$�|�0�]n����|������Y񸇮�c��������?l=K�Հ�͘r;��zw���%�_]�qո9n{y#��+�eͼ��5�f]'!�{]�n�Zڧ{�8�����gٛB*�Aےb��1�ǩ��mR�{N��'<Fqn9��O$ъoxYT�){��3a�o+ݚ���!+~������<��㾡�ѫ�/1U��/����%]� �:�hy��{$~�I�=���-E��q1"庖>��Cҡs^t��%�º��=�<B�C�� ��㸕�g{&&3��ww=�ZZu7����\1;�h�_�������R�elE�P>X�>xM~��#;�f�Oz�������Mk�o=v��t�Sg{�l�Tֵ�٩�BX8ɬ�6�J��P|�X$�S�܋�*9�>K���ܡ�=�ȕ�	�7��L�!���R���S<�~�~W���������
����b�w8u���.,��:���}� n�Ʃ�5�x�[�~�Rb�����1c�'M_s�8s�S���5���^���_3��b���P܏��evs>!��]t��.��6���B߇���;����6��c����>��`Q��T����v�H^r^����������7�}�Y݋�$����N�C�]��Io�U�ߺ�݌�T��{��W��9��i���8�<�x����=+J����P}�����g4��q��PĮ�}r�E����o��u�ǳiƒs�����l�^|w ��Z�`���v����gg�?��jB�`�U�J��������+�yy��vq.�<p�/�pZLl5���6���֨��b��P<x1U��!�齃�j��b>@%e��8�P��(��%]��-Nf��:�Sy$������ܐ*��<f����DBx����-:�wC]}���y�39q��jfnz�� 5/}y_&��Ʒ<��<$�."h�|����>��Րj�{��0ӆ>~�;,�{<�����	���'kH�}�`M�pT}m�}��*8w�:����
����h�{�|{ sei��;��c���'�����ڗm3{"w���'�y:��;e�Vk� ����6�¶�f5�/*/�|���p%�&OxW�����:���vܧ�o��u�G��-=���e�(n��1�ci�u�̯\6nL2�A��ir*�m�2Fᓣdrd�٪�y�y�^�eD{O�gT$�����т�-�e7O[a0-ͽ���,`;���s&;V[~ wy`�����{���9Jཷ��k��"�������VկK�Anm��B�ddPJL�a��BASO���Ή��;�o�<4'����� GN�Ѿ׮���}�0R�C����pދ}����,�2��H��U=������&��1���o�����_e<(�3�����}���{:?.\Sֽ���d�*wg�n���t�4��)��Ys���`dT�9�8Ȕ���a{���ջ��Ce��m��SՂ*��(kUU�珳����ys�G@>>ǄA��,Ʈm�^���P!�<��.�ӄ�u	oz3�c�ۚ�x/w� ��mx�"R"��BO��j5����m�mS�9�3���-;{ݷJm��"o�aߵ�����u���/t��]�d9b�2tA��gm�2q�N��u�v��ȵ��Lp.8�����b�=��o�)��{JxE�߃{��_���� �7M	���
������@^p�z���k�����M������>��֣�P��Q�M�1��u3V���i��oG}E�ʈ��oi�F����W�2K�y�^+s<��SE�N�b�nm�	K맴'x�Hhlt�T{�.��x�Z�� �Oy�Bw�[���)ƓU��핤�kpf�31[���H*�v�0��I��N�<��wO�o5D����b9���qH�G}w9x�m�s���t�����	�u7N��r@(3����e�a g��y���3����NA�7���f�*�/Ȅ<�Fj���1�ǇY3W��{�Ǫ��U���FF�\[����V�Ư^�[�N�N"�#W�ư�����b#����擅i9��4:xW����=zv��V&���y�ZW;�nsa�
�׻����=�>{B%6D�y|p;�T/��������Ǐ������������KϽ'z�~�x����%�n�Hx\Ђ�G-2�ui'5�x�Ά���AzX��$GL��E�v���=3�f��S�E����j��'<^��>��#��o��_���P5yd�א�{zװʄ\��kV�n��J|
���j�1��C��|h�Xů���<�����{��<�:�V8흽xl�Q��9�ҧ�0{=ݛ�Rt�}�r����od[w�{��7�Ë�����~���D�a�<�����c�CĆ�� ]�X���Nͤ/5���>T�惖-ᛢ�m��q��2������݇P�����,�����1a'O���Q�y�_K�輰s�C�x�^�or� �~������5xm\G�;�����1���pz'�d��=y��Oq���e�/MY��^D�/b�zu[*��N�iKB�<�{���,�m<������7ʾ�Ã��^�����N],IH1P+C�(O���ww��� �3j��!�%��}ع�{e�=�e~�ClB�TY���]��p�g�� {`�v�e��ћ�����vS���M����0�Ͻ��u��]�+��ow87s���z�[z�� �:��<�ޥ�Ow��9��*�gR"�����ò��q{}�L\����	Z�z�߽d�����.pg_cNu��Cl��^�D!��Fi�u.t��{��ٯ�t�C�X�/ӱA�
9��3\�����G;�����g�����oj�7�����m>���wl|
�P6�C�O-�	>;�"-���|�����c�nйZ�{c���I�/tfw�<����og�lk�5��}����)�������=�h[�n�[�꽮p�0�c=�<y�b��F���g���^˭ߢ�
�Q�(����� ��zg�	�Z0"���{�J;���G���+�F�m�������7C+�q� �,W����q����U�x����/�y�}�gtv��)%�|��S ޸�&>��V���7W�%�L���5-�òJ콫{��8���M;�}���ۇ���k���7ަ�wqI�6����ݞ�����>7y$N�����1	V��,Y�+ݍuz;���y|W����M[�,�ڴ��a᫓�㙹=&�2�%`�A�����A�&ي�O' ��6�Q}�f�9Κo���n��Q�7O�&��g�ѽY�5L���ja�7�����r#���hY�1kȧJ�����v-FU��Ѱw2\<ףm���S�c�;�t^�l�~��j��:*�C)a�)�	b��}�ޣ�I��ｂO�
��b�C�=�}�g�����K��̼�6��v�.�mJ��av�V7�U�ym�^�<8-y�����8�98#4��8&r�=Y�޹�go�7������~<�I�n����U��r�,P�ƳSxaBhѣ�����y6�=ꮿ>T��>����'n�yDy��������_l��>��/�����/0���Ur�6o{)h��[� ��=�J�q1.x���wV��W+���֎�]��Q�(��C�N�nq*�ٺNM� 
Z�W��9� 
�@񦅸��\����!]�k�t..�M�y�>o�SbL�٩4-T\͍ڽW�7*��.�<{��V v6�ԋ8[k5��J�g�Ͻ����v{q ��]����q�q^�/"��4�Ӵ����%���[�6�����X��܋$N�r���'v����7i��.>�{��w5���u��|&�"�� <$�1���,z�܇{�r>~���owˣ�o=����Α�<[�M7X����,�wW#�1���u���W���.�<���������]S3����w��S���L��n�϶D��n �m+������LD��߼u5L�>���;&��R��E���M�����}�N�<u �5���b~�� {�眒��)Q��c}��̑�ho!ּ��7H����5�I�p{k��w�:�x���˴,࣫�s��$N�H	�=�Eʹ��
K�׿\�}_��7��>�m�yMnI�G���������.�������	}��"��P�:�m�;�
�_��HY�n��we�f�
$a�Z�Ҫ6{ޛ�=���~�������̎�~��v<��9 ��}�S.]��^}���/A�f��6��f���C@>a}�0�.�����7q`=Jв���yo����K�O����NvU���G���%�H��ú�t�9�o,P3��<�y�����t�>,m�=� <j��^W�m���k==��_���O�{�J�{� d{8W����˞o����ĄZ��Z�����V��zcc�W����ODY�}��6�G�Q�y�
�K4��LR�:�])n����rD'��Z�^o�{Ǳ/���^�s�S�����$)fόnJE�؆/܈H}�a�aS>�ūO|����d�{S���t{s�!������7��%���]O{ːj��u�{fz]{��?p渞k�Gs�_1�gCo�P�j��yj�i�{X�u���ۘA�n�Uv��ۂ��NG���O2<h����\/����Fwxy߼D���t�=pg����<�nEE>���P3e��q Or:�ӅK��A}}H���̾�|B��(�;�|�"���ǯ}<#����R�x;���W۳6�==��ڏ9�ۧd󥊁þ#�qZ�Lޖf��z-w֣�g4���أ�OHּ��� 1���3��)ޫ=�݂ƹꌈYHt�MC��zs|U����������v7_�]���7�=����qɽ�<�xu�rFr9��un��w���X�uCD��GƁ=���{�(6g>o��׶��X=����f��1�t>��/u��K�xk�,Xq�D�"���3nvٜtQ�f��t�x���W�K�ߨ*����<{䫍eõ<Lxv�y�A�{�pɏǅR����a�^Q�� ��x�r�-�+
DP/V�6,����u���1z�}3/�P��ږKfz
�o~�G(px������J���|ν}�Yݤ������4�=�;n��.����x�i^e����ӈ�}�@�]#l���|xS�ab<x�(��ʈ��&��t��j�:5�E����<�����\�K���g�e�MVgggY��-�S��tK������,}�Lj�^;݌���u9�6���uY�Gu�z]Ou��G�k��R!��i�g��^Z�M�Xŷf��֝мp��AQ�S�ݑǄ���{Ǽt���r�ӽ���B�U���D��)�`3i�I&{�[�7���Iv<ow[�F]���t3ݭ��{;�y��q�<��ϽS*վ�[�1ϼ<>^����r5��S��P�b|ϝ��u=3��K�~t3��f��3���{���`� ��G�8+���/zr���Q�B[<�'��Qߴ��sZl�=�dzDӺ-J���w�z.��<��V��s���{�>����٥�D�t=6���f���#�[���Z.ʑokv�L^�i�m��8,׳|�l;��n�rY��)�q�̯U���h���;�F�mη���N�t�6��kE�Ӎo�Z=�xg`��@ﯼ��>�a2Kj"���u5i���;�p4z���gy�Zwa��o�inoa�j=�;'Y�����u#W�}����҅����A/7٫�vn2�8�����آP���c�ق�V=�xa,x����(��sP��Y�ռ�\�^X0�9�og��m�t��=�h�c�:��"s���s�/�h�|���7=�-7d���*�����\^1M�g�!1����l ���\'�^���_^��jk~�J���^y�~|j�x���K���Ϡ��{�7~�)>eg�au�]������4�h�y(��p���"]˚
��0��o.�jS�u�X�������}��tU��L�6E�*r�"�cjw�{н�Q���m[����/^ A2ebv,n��9	W�w�%��s��͘%J%���&�h��ff$*sx31e�Q����{��{ޟ{�6����lS�Yu�WW/K�n+u���:!k4������:���]f�$��M����z��ܹt�u�[���W\I���j����5���L��&vy��M�t���1����q��Z�v�o v�K�1s;�ѡݼ-�vݗ�#I�9��9��k��8O ��kV{7]kX3��Oj�;�����x��肎�m��^y�o I���5\'�����/71J%�����u����ۛ�^NK6v8:y�9t.�n�pu���t��mNy�v��n���ݑ���>g�lpkq;���s붑�<r�3vz�k1umn\�8&�gWiݵ�:���q���q��n�;&v���@�㶍۷�6'vy�M�4e:��s�#t�n{S�{EùۮS�'�\^�2��/w�y�Ў:�[��x�m�s7=�c��'y;r��y�mt�9���,�Z5����n9֔�6�\	d�x�4�6=��ֱ���u۷8<�˼��U�˼ի�&�cl=ŷ8�z�[��x�jp�Qp��.�um�=\ٽ�݉�u�:J�`�c\*i��Fs���6�^q��d�h8�۸��7�i��{`�p�b��Sb^w����(6[�)���Y���t�1�d�@wA�N����a{��0�-۹�0�<�E��N{{mh7�h��'�J/��h�"R:;=��Z뵝=tV]s�����]�iy�n�aЁ+v�X�G�g��]��o1�솬�����1ǄБp��Zyz�7F�p�A��Ѫe�R�Lr�3mn'+�I�l5!�n��M��v,ح�s��GEuWXm�h�sb�l��n���۴n;8�q+<o�;Wg�l�ό���8��q��ہy���c;���k�9r��r�um��3��`+iR�7%[n���qӕ�l��#���J[O�][pnݗ���&�E�0Lہ�{F9�,����ܨ����Y�7X�4���ݴʛ���ݸ�
�7)�A�ni��&z��q�{F;=d�AەU�u��n�gi�]�=�ta�瞯>��ݬOnՋc���۵�9 z(v;p���9�%�A�u{�:{m�2���ڞ��76�؝�ō��:x����nz��4 �:xm�<�:P���n���{e9(҆8E.�`|jw�䦨:Wd�nܔ�l��kmNE���l��ɷIx�k����o��Q��
�q��l�Ȏ�n�z��z1�r�Nԝt=���;q�̚���rn`��G��[��Їk��Z��r�.�m��x�ۺ1�ݗ�3Ii�azsƍ�te�c�ku�n!y풺���mzݵ.�+n��t#�GuC)���1V�n}>��o5� 	n:ۛg�]��Nahݺ\(�vdx�=��� �dۊy���W`6l+�mWHqg<(-�s��\�lGpG�PԘ.�wbn�q������X����m��u�w�<{��DY�v�{lB��싻Y�g۶9��g�a]�c��i���-���gt����m���<�s�9.��y�۬�l�*�\�r��v��� k5un��)6�#�6�8.��=j��T#H�Q�v���ֱ�ti�H��I�I�g=�����7��x�H�h�pv����v�ں��:�.�͝&;q�۞"z��s�wn2.�������[�y.�Qc��'�;`��b�mj��MG5��8��$��� q�s�+��R��z޶66Ǟ�����>�n��]oA�{&	�w+�ֲYݧ���k������mW8�z���n��a���}Nμ�v8y=l�2M<Z�soOny8-0�put�:ӌ��)��n�QT��[/���MX��ۣ���r;kv/C��qn����pq7a�źplb�u�<0;�{)�ۍ��]���n���PrkGZk�;��l�ȚӣcZ�]\㓍��Ӛz��N����*������;mY�l],n{{Mc
@ۀ,���غ�����<��n/J�vwm�]�m�;��K�9�u�G<୚y�i�v�{mw<�˻r��mq���k@�c4Y�.䚸�79�y^止S:{p^�7���5��yƻ8�����m�3�NT{g��{.�Z{F���&������C�z��-�����H�t�&��c��nm5�+��p��y,��;.G���p���uԛ�X���i|��j`��tt�Z�8����I��3�
����ʣ�OwO��=>�[���Nΰ���T������rP.�unnv���)	1n{
q��]�R��kl��*�)��t����e@�ׁEe�$Mv9���t=ŷ(��w�$y��v�����=9m���.;\\��x/:4pvޞ8���r��^�u�f3�{r��C��M�r�۟J�ӥiŕ�l@:]�vyۮ3d2��ݮK��X��V���G��)�뮞#��7��q�xm�1�c��[�T՘��;p��b�m�: w���vza��Ds���+�����@aJv��lkN��l����f��#m��7Bn�q�ˈ@�۝˭즲E��[^6��� �z�%ܹ����c�yU�G�N���7&x{[ qvk�^��/7v�O�l��^,��p���s���j���y�C�����B���;k��.�9�_ի��MpM�.]�F��Q��ۍ�]۳�%�}�x,������ݱ�z�]����V���,�ͳ�ݮ�ۇus���r';܋�ظx厇���͇�r�"�q����YS�^7N�nm��ں}�6]sq�Vф���nn7=mг2p�8��]�v�]G�a��vR�y:{���{r⮱\p�c ����Gf���E��\mBr�Ta�9�v��ޚ�[qӮ��ݻjvyŝz�n�9��O7�s��u�N(𼝔��ꍷ&���z�x�8�G�欆�<!���Q���7
�c6��z�q��)۫p�gK������fwqɞ�V��'3�#r����ٹq�r%��rp��>��)���^�kc��y#q�nM��:ݓ�Sň�����q������e�ϲ���lD������v��u�^�&�^�ݺ�|�1k\<V�iPs׎��q���r0yw:�8���x�G�xޜO0��u�3�sŹ����]s�yހ�;6xU�\�"�����v$鲸s�c�헴M�=�Mu����`�L�Q�T7���m�����۞��pɧv�/
@rv:�]�˕�n3<�S�X�sk�M�p����x�v���7j��:ڌ���q[���{r��;q�A��4�7cA\��7`�k�F��6��,q7g���Z#�c�8/nt��'�X8�ѡM��{e��m�^j�c�����3�r��y��cu1�%�g��{b<�8`yM	غ��Y�n�\�C�<����Q��;�۵��x���I��+c.7;U��kv��n��c������Q�<[�.�=�����G`�r�n7���U���5����9��YJ*VWnv����θ��M�殶�c�,�ܮNjݼ�G7�%�r�ź��{\�8ck��F���7d�ҀU�s8�7W)\n6�6��(9�R�b����V�ەG{a��������7���ƻ;q��͘���u�]�.^�N�;X��zp�M����$�hηcv:d	y�]�2������e��*��5��<�����[�����n��������>���n@�k��aI�n�ݵٹLlk]�m�.��]�sڎ����w��gu��t��6���Ģb��nƝ�g[5C��F�س,`�蹗�;v��s<��z87n�[��t�6�n��B]R�h�D<nh����T
��n[>�D�ꍐ�V�_m��d�q۳���>�n�׎HzN۞S˱����Y��U�[���t��یj�8[�b��W��q��{b�nX�Yvw��z�t8����ֺ�VI���k`؎ز��k;�����j�,���v;��a�x�AQ<6�ۇ�&�%d�\Qcse��	m-�xM=�Ԥ�v��v�n�OC[^jv���dwbۜ��۷��#��u����d[�������b�#��Y'��mk#'cn{[�r��7�`m��]Iuͩ��X��-��p������"��.]�a�Iמ��V�z����렱�ڽ�=�;�#{Ͷ�۶���A�۳�7Z��<n�6���ar�דZ.-@�M�<�q�M� &�sǜ[��۱��n��v-�<�ڸ��Nc�"]�`�g��^�5����<�kkg�-��qx��f�m�u���㳳�o�.n9�A��w�<ۃ���݉v�r���[`�@���)�<�k����[�8�9�cv�xq���m[@�1�5��`s����lX:+�d�E�r��.QMq�f������<tj�{]�ܼ���m�"^�3��u��Ƀ��̒�����ǒ�ܧ�n8�8����s�!����jy���/�vŊ�Svn.�G����Zwh[��k����Hph�v��Ѹ���q��G��s��g��y��8n֎r=����q*�j��fm��L�yx��8]q[&j�6.�X��K�[GF:u��N���+{��g�v�D�����#�(oSu[d�v��t	��꭛f��q]ָ3�a�sf��m���������-����zO-���<�N#��p�pS.tOb�omۗtn�����)7:̻�<g����g� m�y����=��V���|gPh��#����t�#ry�:2uG�7fꁪ��̃���}��OK9PA�C�j�'�Z��7O"��.Ϯ' q�����5ێ�g����]���8�ų�y�ձ!4���]hy���l�]�u[Þ�}V$���r�}��5ik
�֪ѭ����Um�F�5\�\ĭJ���2��.bTµ��lZ��L����ѢU��J(��Kh�Z-�T�[֍R�UcD�b4��Ekm�KZ���,�E�R���ڊ[Q���fGF-[�����KJ�[U*�*�,�R��\ml1���PD*"R�V�b�E+bթilib�Z�mZ֭m�V��bYjƕj�[eV� �mh��m�m��-m�Z�ұE�P�+am��"�FŲ�,KimF(��څ�Bңklj"*"�m�Q���KQ-J��mZ�mKJ�F��ZT�V�����Ѩ�R�YUm�Kl�m,�ũl���jZ��TV�2��A�SR�5V�b�l��R����im[j�-��Um)�+��JV�)j�31���[-(�-�Զ�����U(�1�f[m�V�KA-RڡQE��$m��QT��ĭ��"��
����J�[�)m`�E�0�%J)UkVҨ5���V�J�TV�jfQq)�I&m�?���aE+f�քңR�t�A����]��yn_��+N�Z+t��p�'�l���龶�>��yc���/lqp�=��D�;q�z5��9:�b��x�腈YpV;vӸ.���^7ܽ����<����9��n�<�ζ�ݷ6\��m�sn�m���|]�s��pGN3 n[e��i��q�Q�^e�d��P� 8+����&�g�6�鳹��l�,��7=�`�K mX��	���.��3���ru��۫B�ѵA�ۃn󵕶�7uiW���e��8����6����-�󻍸x���r]�=��X�Uv�u���<���m�Ѵ��8����Q��]�z �v	�<����lc��t]��eQ�b�uD.�.�q�6� C�۱�+N�����	���k��qvΐ��'%����j6x7\㧶y�[z�x�@�l�n}v�4px�۹9^]���w��d����E��y���֞,�����6���ˮ׋��p���� ����a����{u%��mr�c�҅&�ƛv���uU��㝭�Ύ��'f�N㸸ε⤻x���1v;��� �Ol��s��q��w+B�������oJ
����<���u��=6Cv���.�)^#�����v�,�ݫ��ۡM�ms�Q�Gm��ۣ��kn�m��ܝ�].�D����G��9���N�bs�8惬ٱo7����>s�?Z�';�����[N2�yz��(�my©���uu��kg�\M�k��խ��]��n3�:8r��.���'�������ƹ�M�'�Ka�%Fq�^�wHu�c`��W��q�^ܼ�(�u�瘌d2lV�χ]I������یn�X����u��^����mH�r����N<����m���Ǜk�Pn�T+Wv��x\*��m*�v��5.O]ls��WY�M���&<����@.�cO����w��m�N�n^�p����|���;n��+��;82�q�gs�og��'<�;cvM�\p�{v�s��g�u.Y��\*�L\kjܕn)l�q.dj��mn-p�E�(�s���.��	��l���۟��N���=�eM�#�9�w;����r�;p���/&��es�;���#��a2��9��og�|�s��<�N��|I�$LDO�2���S$�w\	.'~�~}�wCDUSl�Uf��i��kx���~�<��?���Fj�� ��;�`�{�H��J��wc�#(�hD/(�(D-�_6� �s�	$��u��=�	%V��}��H��)�0R*&%@H�3<��ތZם��D�y\�A�̒^�W�S��[�[g��Uk�%R6B̡2�5��"�}���'Ռ��gg��H;�� ���l�Ѵ����*fM�b�z�whI�ۅ��1έى��=��mŷ'3���P��3�I�G��l�NQ$�����`m��`�I�N|���'��,cX�� �w� eS��'���o����8S��o�z1Wf9�]Y�Ws�;�����=W�dY{n.��p��I�y��B��>�{h3����U��$D��:�A=�̓�O����D����Q�v�{\c�S�0TB15�$�u��ƫH��Mv���z4w\O������r���B�2��SLN]si�eQ���Ă��@'�E;��*��l
�<j�VV�n�pf0i����7g�@��Ѓ9��y�'1ȟ�Df��A
�y�f��z��;#��DL�>BD���i�؆��k�*����q��8{\+�ͳ������	�BgD�H$�=���%U�SlX����a�j 4�= ����*�#Q3"I�9κ���w+�丟כL�b����Śk�ϯP5�V��L�z`B"i�{w�̒���~$�3�Dh\˧�nD�28��X�qUqD�{X)�۶"L�3!��Ў	s+v�OgT:�ȵ�Q^�{3!�y]��v��X��#��`�D�+q�����U�6��0�=2&`��b(�ȸݵg�e��=�6�$����'���ӳ1$�Ă�oS��Y�%�eA���9u͟g8�Su�e�=K��&+7���q Ý}���s�S���9c��O%�k�y{u��,��$hwf���+%�����w?�������po�jv�	�1]�L�A=�D��a�QLSO:��ă���}�&���3(L���|I�p0�gT�R����d��� ��י7�Bݥ�dZ��l�PD�D@�&<���<A��H'��=�X��u}�''/w�q�u�	��>Βh\ mc����x�'o<�w=�	�D�
�ޣnf��f�G\tf>[.��H�_n���?%'^����������m�W�69�X��͈��]E�б]c��=�	
j�mGT�l4D%��p ��]���R�Y��oS� ��bA�}��/7�Tw���/���G\&iVr�n�[V���"���+t뫟h�>�\��;����;fڅ)}�{X�cؐI ��l ��:�(��y�����'��J�&IRbTL$�x��[g�Ƙ5�q}գĀI��$|U��0I��UZ���������C�I0�ȥfP�l��	+^s`�b��n6nZz�{xa�'�HW������SI%���ߥ��i�F���l,��b@ �HYw���H�{�}Ƥv���׹4	�EY�$��� �l�a�|b�u2��Y�e�H��*-��HŽ��}Y2#�-W��l��ۯz�󾪛p�J::/Q��l[ۑ�W�]�Q���E79Qi��n�J:?����� ���20�P�CC!Df���6�]�����=�5���=G����Q�,�%Ky�m��{gY�%���,����}v�lR�ܔ���/G.Nۯ;����{m��ٝj3l=ѺŹ^�˼�hm�;͵�{d�ns�.�@Hb	���j������mM��A�g��mp�����-�§��Y�v�W]��'F�c=Dն0��^�gRtt�m�5lƊE�!ں�ű�g[V\[]q��76��?~K>���DB1n�&��o��H'�o��P�&��}���|��ٯA0��	�]�$	�&eBRؗ�̀I��
���js�.���$�[�b��2A�H��~�U��VL`<��h�7�u�|H1Y�L	��+"q�geE���C�b�k`�DU�6/�$¿"�	�Be�Uu�M+�7�A��� �LWg6';�wH�����N[�fNg67f-@U$��[�����5YKuN���祝{��$����9��-x��&$*$R �vޖ�g�5��ދpq�CV�h|�v7!c��ῇ�3D�'x�]�U�Pd�Nw]
3�s�ܙYS�X
��a����LzfCA$BZ=���>
�~�:�^���y��Ԇ�o �uE�Jg7U"�����5���_�eR������~�j�sr��xpS�¸Q
�v5��> ���l|s��xAjv�������{�cEf����&eBR�T�0�7��>$]��xi�%<��EWv�H#;���E�2�*T�(Q��y=�s�"@1��L�I��z��ީ��Y�8sI��n7�}Y�+
��P"d����s@�D��oֱ�(�H�ݭ�H7�� �׼�y5�ʪ�̮4�LI�	}�lƍ˸�n��gjwQB�c�{<��WZ�s�v-d��w�����_~~�ɀ���G�I �ל�1�����W6�$�{�h�.8��&bH��z�V��E�8�f��z9�[�A �[B�>�y͒j�����WSxr��DL�fL��H����O�I��)�]�H�+��׫U�<����ܐ-mB5�js*3"�x]�H���\����ƖvhO�p0n�l�Q1��5�+����ӹw�A�Gakl�֌澵q��	#r�}Fu�S3b�|RHē2�)�2*���8�s�^t`���5�&q���H���0%E�8��OF\��\�2
���0P�fsn���i���1���U�$T�P�D�ޠ��uo6o�R[��Q�Lɕ&D8��t��Ռ�<�����gO��ǣM���	��%�? Q�$L�-��H3��a�kky���]StoEm�zw'�O�����\+0J�2L����6��)�dfN[� �g��0EuoS'�/h�p�B6ә��ѵ*e����l�YY��A1��т���	ל� o�߶�un6�M�"B[�ӿ0����֌�{ �T�u0A���$�����8�U�1�bv�ݙ�׳����-�G|�˺���-�qv{�F�\���vI���jh�,�|����y%�pU«0����8���0�EgRHă3���ẀA7ճ@��:��7w� 8�����~$���u4��R��K�F�n���A�vӴv��Ö�sI�\ۮ��qn�i�UϳL~~~�s��pX5g��ݰρ��L�O�ͮ�@���Ѻ�*�K�� �E]n�L����/`D�-��sDc�R���Vc>�*{��Iͮ��Ƶ
�`�.ہ(Xl�eU��n�F��Q0L���cd�H;��(swWSc6�^v�>���ǈ'6�h䰰�J�Bz&���0�q�)�Iou��$�ok�W�3�z�0Lm�����a2|���:/��,bh�I*����@2�k��q�ö]q[N���D}:�����WU�߳�4wv�^˼}z:ZMO�j�_f�Ǯ�-�W���4�g�X���%�y��lZ�ڜO�>�V���]��]�w�X�4	���[�۶צ�>��v8-�ckbl�ls]n��=��\��u��<K�v]Utn�ۙ���u�t�K��Fq�苵�5�<q�An�A���ٓ��Z�q۳��mul5]T��؋���.�����xh\i����i���]�Q���,e��^��y�M����s���v���W=�F��p퓴���>��`{�]	�v��x�U�*p���z]��D'Z�;�1睵�v���J��:��%D%>]�w�)$fI��J_�Sxߏ��f�H�ν�`��[Sr8�l�֐|skf�g�E�2�(L�(P39��*䝪ܞ�u��`N�u
"u�S�''�g��������jJ��FL�2�+���םL��5�Jr-U�l��t��L��l�m³��dDJ&}^����TХ,\k��MA �;�d��ޮ};*��39y��̚'����"g��[��̂*s:���B�.���<�7}�(�|%�����~>�M�7;�~�=���?�� MRmҶ���{j�0\������v��qХ{�?~?�fT��ADp8�&� ����'āS��Uӌ-�Dnt�D��l��X8��3$��-���`���":��.����J�^ �n&.�9��/���D�c�x��{����,���pe,�_��0�d9;�w�ŋY��qe�U�hMTk��3Ur���I3�v�>$T��d��1�L!��/Cyn�����Ș0�2P�3�l3�A���`�ӎ0�f���$��LA5;�߉�ԕ�%��&e�W]ˮ1�3������jw9�I>9��k�N���%�<l���&�)�>�y�� ���h�̘�����UXQ>��l0O�{u�@#5�)O6�"g�vX�$���g���j�Iɂ��.���u�%.�x:�u�_H�����(DǤ/D�x�[�'���u2A ����x:�m��i�����lI�����P��*B�ADW�ol��U��w���<��	���'w�}@��!sg]�&tc:JI�bT���V	 �m���ꍾ˺��J�i�EUsp%� ��ܙY�I�x �P�V�^��7��(s��Y���g?�m��Q��G��Ӎ�MY�t�۹��x�]����x�� ��M��!R��vh2���F7R�f��t0j��vtz��w/�g����0I���{7���W��Pgw^������a��Ǐ`�
�msFu� hNU����^�<���:�<�rE�� ��
�ks���<g9��,yqҪ;�]�Q{�n?{���ǹ�q�rz/h���Ga�p�;�_y+`K�Խ��d�b�#��i\u���ۥcZ��J7N����P�^Kr��S���F��p�3��=����J�g����ņ��q���T���_o��0b`V�u�zvU��}�_��x���49W�M����w���b����o�V�����ͼ}����?f�������b�&9���<���rQ>�4ϋ[��پ�(I2.]���ba=�I�����[�]��X�=)Y/��~�/� h�Ȇ Okּ���e^�1�~;�F�s��(�'f�m�}⚋�O!�n�~����:8�WV:+}��;��w�Ix?5o"p�~w8�･�n��}�%=���o����oy�ؽ�˂����&ڱ�8OL��f�W�Y;�{\�f�SnD�yAr^vjC*�ҙ����x�t�	��'��}Y^ף�N��7�����%I�fq�ئ�^լ��'۔��TrF�$���8�ZЏp�R��V6��L�ĝ���HQ��˽��,��:Q�M��y� ��-~�,�Q*V��[Ee��²����-��jҊصKlj�U�*�VPZ�%[
U[�Z(�-�UQ����ERy��Ekb�2��QE+EL�L��%d����D��ڬ�h�X���*TP[e-+R�J�m�PmkEAT�l�
V��R�ҬA��Z�U-%H�-P*[eE(ʅk��+Zʖ��n"�+iZ��ړLkmm�h�"�jTP���FDT4YJ��R��h��QF�KB�-*�F�T��� �!U��T��0f%��m1.[S������+ik-,�XŭkP�kU����-j��-T*ZT�m��P��EZ�E�����D����D�R5R�Uh[F�mVX֣J0F�i[l�����ʶ�P��Rѕ����c+���J��h��P�#k
��6����#)F5--*����j�DkZ�
�Vش�(���Dƪ1+*�(#TV����FUiZ�V�{��z�S}���N�\׋=�2	�" $�Dg9�0NS\#1O\��b�2�'ċ޺�Z��
V�t��x,���l��I�H�X�0ܟ)�@��nn���Z�q17��}�}��:������úV|��1&[a��±�E?���Ab63\=�T�cj��2u���ۏϿ��M���#k�;{�� ���	�}�09��$��p��l2;:�VCCD��W�[7���d�끹W�sgU	�����>9�r(�'_s`���8J�!i����`��9%dLHQ(�_l����L�ˊ�2��	$ι�A3���'Q�QIL��̷�u�]<��v¹���h�A3oy�MM�5��wB�Zy��E��7?T#}�E�s�kM?^��vY#"�O�6L��*�9��ll&�is�������_9q�����3^%��F�`:�=!����K'��Fg6ߙ �S����%X!�s-kz�W�� Ky��	���)��dٹ�������8�:�lCQ��8��M�Ӎ��e�wm�c���<<�#��g���?_�=��u���?>�h�y��A7���hn��ӷ�c� �'�cd��W	#1"����l�rc2&r�i�wN��I2��d�H����'�Bm�
�Ƞ�dl�l�|:�!A^�b��H���d��*�p��FuI�$'^sd��l��צ��U4��7�k�����M�z�q�	�^k~$��1����w}`N^�d�tc:J)L����o�.��A �m��i	7���E�f�q�|LVo0�#7�k�j�If�z�Jr�_���8'��Ud,��������d�"��2��M��+�&.x�ǌ���%��
�{v�8ڧ�t����x�C��^�z�ST���
��(�ۏW�m�=�5U�tS��av��]r�pz �u�lt�ME��*Bga͹�ۧ�wb���h���7mZ�㣣�������z;q����lh� ��7��/>����6��j �����8tά]u�a�8�� p#��WQ˓��w-<�C�N�}:��k̆N��N�ݮ$Lbz��mm['K�Z
���tv�6��̹{u�:u�:g\tawDչv`R�E^m�y�#�	�b"Jx����|b�v���t+���k"m)�m�6g� $��O�jN.!x�$I�l��W�WoWU��q��"+w��Fk�	4M��d~U~���G�8V��R O�f�` �Q/���jEn��V�ט9��P�aa�a�
�K`���Q�a!�.c�n����F�����b��[c7��}KM�&g+� �s����2&$(�Ey�^$�-���E��۬������2|s��	�{�3mw��M������k�F�Rek�8z�F9���L���1�YN�m���}��z?{����j�cL��۬a�@7�f�>$�8��!]I3WՍ_��y�<O�ul���EɁ2L@"$IB�fs����T����8d��jɹ�g��즾[p�µ��+���*�p��~���ǝMݨdٞ��n�Z|��	q��UzopL�N[��f<��W2���E�+�߻��R
r VQ7�}�p�:2VVJ�3wU>�[�נ�v�a�h��fL( �$I�~a��{�{���!RX�a�{��:βVT
��x����y�~ֵ���V�(��}����R�����,�o�VBB"�Q!	� ��eG^^��NOG�>�}�|���������P�%H,.�w�9��°�
���}��:�||�����Z<2|��Y_����N%@��_-Ή��Cfk�P:%a��;�ã�jB���y��������zqEn�, �}�U�	8�R��M������bo�,�|%\��s:k�]:af�[:zv۶�N�;:��o+��]F���Wj˂J ����������~X�n��{���{{��y��#
��%�7���γ����P)����:�Ԭy����������3ݰ8y���p- ��ίl�Uh�|I2�b_��/�z's�G�>��#�d9�eT�&'z�~d�
����}�u�c
�RT����I�
�YY9����֌�^>��o�����T�|?c��9�]n��Xo~}�a��AHP�}߽�Ă��[��5(���b�Uw����#�F�k��8r{������a���`���ݺ�4=�k��1�萳�z���ˣ��k;��O�
���ߝ��ì�%e*��l�V�z��
0"D���g�ς1�eP"�w7��z���ԞD*J!Xk��ݝgY(ʁR�P׽��H,�H/�����}��cغ��x!�����׃7�i��_�S.sC�ц��w���g�
�YY+��{8�P��[��}y_��:����}�9��
�RT���ݝI�+%���2�{Ϸ�
�p����w���P�Hn��.�۶��OC)�����)�C�|q����_����3�c���Aa￹�����F�-�k����$�!Z0+O=���
�
�֊������g�<gD��wp�:�YY*�;u#����L1!D ��I�`�#ד� τ�H�i�?aʽQs^�s��ϣ:�c*J�u�~��P:%H,
5��k���R)|���o{�ߡ��k���с[7��ߋm�ևMˮ@�tf���ΧD
��YY+����Ͻx�G�D|��鞌�?�w�����aRX���}��:!Y++%_7��
��߼;���))e�@��V���xXygC�����jB���s�!RFo�{�8�R��5����u��o��Dd�c�����K儴�*��gy�����-���~��{w��7C�Z]����D��͹���J�e�迹����� ��zϾ���^wP�<,:w��|����p�u�C�:¹ߵ�a��$�B�׽��gA�d����͟}����T�����bV�`Q���_n���\��ۇ�+����w�So*�W���Ԕ!���|W[F��x�Fv��#u�pQ���`��S� �o�χ�!�=��4a���I��y�Χbe++%}�og*IP�J�럽��Y�P�֫rw}�G��O՝B��P�������߷�8��x�ֽ4c�4Z���tJ���}�q��jC��Y��u�5�w��$%!RC�}�9N T�ʚ��~�:��J�P�����k@����7�y���]f��K���q�~����80�%�V�~�gY�J2�g<�-�Oxz�>�w��dJ��X�����- �a�{�ۇR�~<?|[m5��
_��,�ߨYRY����`��2VQ���{��d�T�
$�,׽��C�:°�*J������?a���߳����w?Y8����>�{��=�Ø�e�֓[��_y��=�
#�y �����[�d��������m�0+O7��r�*X�Xk�����td�
����l�IXmד��g����^WP��p�ҟ\��m��pU/1���W��w#]���*knl��D��aC��Kx!Q>���;�&l:B�K$RI�[ڡ�;�3�@��{�o�j����ųF�S=[���IƆ�I�{�S��j�Xz�;��������
퍫�m��Ѵ������qv[������A���]q�Fo=�$+bz�q�ݷgv�8��mێ�@vu�Fd�g��⇎vH�A�!�-F�;�;6.��f}��s�3k�6Ů(��Ü�������e��������dJ藞:�������v���r:3n9��RCɕ.1��s�q<���N5��'��n��7������j�:��0������R
N!Xk����gY+*�S��߸u�X|���0���$^�����)l5����u�������fsC�h�@S�O���6u: VX�Y�yw�w�����=o�����T(�����>�:ñ�aXT�=��gRtB�#�}����ٮ�1�?��N��W�$�_5�a��N�q�%a����a����hw����)
�Z��~��}g���}�<�����5�~�p�:2VX�P���~��:������ZebB�AC�<	쿪���������I�Ib������3��*���l�bV�������
�fG�Z'��G��<^�ۯ6|��+J�htܺ��k9��8��d����Ͻ��FJ�y�|Ͻ��y�I�6���߿y�u �� }�;��$�����{��'�{��p�Ͽ�����?��{lsӄ�OY^ٻE��ش�R�O��LװX�T��Ɠ�����Wg&Ԛ�Ry�wa��jA@���ݜ�H[HV�+�=�{��*}�߼k�Ͻ��=f���w�ì��R
C�{߶u ��9����\q��j�:�C�:�#�U ��Dy�^�Y���ώ���|�V}G��q�vmFMb�(<�sV|�v�v�'*�����a�9u��L�[X�aM)��T�w������û��722�X��w�g�`Q����{�����t��ٍ�~����u�׆��"��)�AD9&&D�r��~��6u:�YY++%}�og#%B�J�IX~�����{�}���q ��T�Oy�}�ԝ�VKY,e|�orpJ�O8�ֽ4c�4[(K@G�2��������U;�����{�����
BҐ�����r�� ���<��ì����v\�!!�iq�������Ȁ����Τ��3z�M��Zp�3p�#
�����paR
J!Xk���gA�d����j.~�� !5�Ő���cX�}��op9i��a�y���̓�Ͼ�\���`�*�*��$l�:�z����<�6�7Vѕz��.�v`o�}���mK�[�_@����l�Ag̕���������P�%B��.��rH,=.����k�[�1'�3���ΤN�����s�w�8���xw5�s֓\	Xo�{�a׬
Ox1W|� EWe���Dx�~��)8�YS\�Ϸ��%e*Y8�u�[�>��|@�G��A�՚�\m5�:�Y�u�A�s���Ì*AID+s��l�βQ��@�uޛ���&^F��s-K*����ni�&�8v�ֶ���f��D�-�

�C�9y=�ܾ�Ԍ���������ru��DUo��{�f]_�d�#�k�}����ZAH6�<��:��Z{�W�4��.kF�9N$���y��}�f�V�(�����^U}�B�����}����(0�(�o����?w��49�ka�OFVJ2���orpJ�O���_ƌu��uMp�H����~�a׬���<ߝ�g;HS�4���ǣ���󜀧*T
�9�~�:βVQ��bo����u%as�|�߽;�3ܯ�<�1����]����m�a���I�8p�k��J�;P~}��=�umu��\s>��|0�����aRT*J!Xg;�:βVT
�}]1dd#�3���m��}U@䴃e!hXg>��ïX�?�kj\����rS�7���ΧbH,�=y��|��m����(x��RV9߼�:ì+
0�o����:!_y#�wwD^�ڭs(�=�9��^���/�|9��9��\��^o��?=`Q�
����9Ф-�!Z�F7��>'[�vy�����G�>�3��}�u��� �}�{��$8}���2�i�i��C�;����;��JjI��*�|��6u�d�*�_w�}���V��_9���k��	Ϟ%ES��~ǎ�m���2�7�4���n����7R&q�3�}��3|�=����z9�1���Ͻ�Wyr��֖���}��IW��w�0�@����-,=��ۇ^�
�?j�ƙ��n�]/ )�'���͝N��*A}����N�[�O��h������C�+���ۇ
AI؞�����������}��P3��|���9�������m��W-bi�D��n6e�kf�k3=9vv��[��L�7��|5Ξ����|�V�y��X�P<ߝ�g;HZR��yϾ� )���{���Ç-��3�w�����u����
������Aa�{����umn�Uq��$�{/�4G�ﴶ�x_+����γ����@����xu�V�+_9���ZA���7xu���V�V}��8��E<qĊD(�e\�rP5�y��$y++%s�w���
	*%a��M�k\u���\�����à°�aRT�~w�H,���������Ĩ~��8h��:�0M@�#�Z�(��]Ade�$�~����B�0+|�s�<	��"^o��gҸ�NTnJ���:2T*~�<��:������g�2�SZ�\5y��
�=���T�
��@G�_o�,Y��m=�N��}�x�;����D�
��Ͻ��)�!ia�~��é@9������1�<��cg�E�#��TF���d���hdn�c6)=��Q���J1(-�Y�� �'��kU$C�����7�Է|��|wS��VS�k�	�Y�~�y�;�Ǖ,��9�;���;۞3\�n����y�f��XU���[q��ػ���q�>��#���P���ID�:��ɾ���t���+����w����|���W�]�����mҨA���^H�n���3u�s>rH��wS������`z,Ӣv��>���.��Zz�����	��'�V'o�X�	�����}T��y������[�zo�l�t����������.�����$<��ϯ����{�苹�^Ȥ��z��&�7���M�TӞTn���E���e{��F{u����N��8s������ұw��y�ț�x��[W����V��t����|�:�Z���T���� }�۞�YP����/Ҿ]�fM�&o\�vׇ����!˄)�GnM�d��N�vT�z�ɹ7`u�8Ɗ������7p�[���B�ۂg���1�?n��dJ]���VEn��yֽ�Xs�8��Lx�١�ײV�ު��0�zh@V9��J1]�$�m�n�6v�;3���{[�y�{����������q���Y�@��54�vƉ�ǖ��ЇM��(-{y:/i��=dS��E��U`Ļ����c=�?p>��a��ձ�#��K�}A����;�f���z��U�=z���4!� 0�TYj�j��J��U���YA��.Zeks3*��,¢����EijQ*�Z��a`�6�R��U���Ucj�kR��b�[h���ZU[,�+KJ���Ԫ������#kZXZ��ZQbZ�E[s(cF��iZ��m-�Kr��!ThصT��U�T.U�h�e�R��*V+lZ�sZ-�+PYi[ZU*�*
�V�Y\k0�U�P����Pbԕ�l`�ʅh��a\��h��Ҳ�EFV؊4�f#l�mԶ�k+V�e0ȴclQB�ҵ�cQB�Ո�*)m
[m��5Q��%KZT�c
�\��"Qm*(�T����k��Z��J�QjZ"�֌U���S-*R����Im�U��ae���m�i[j�m�kV�m�Z�-��ib[(1Uj�2 入.R�
9m`��T�l��R������±[me��5Q����*TF1(�-�����A�eb��iU+F�ib�+Qb*�5*�F�҉m�������\J��YL��/���uD`85�\�=E�!�[:��h�p��tY�vhu�+8:����F��j�p��8�u�힯m��cgͲ���4\��#h��c��`"3v��]x�#�FA�p���o'�[z�p�rcon����[������:y}�;����l��wg+�r9\vN�����\��6s��e献"9ͪ��뫁����k�yl����OF�&:fR�m6�۬��=�\-M�ez���G�]\t/����oK��q��g+��4<\	7]�4 ��(A=��n���C���Y�c�O^d��p�wk[s�F�v�të:�q=����N����q�7\�t�<����0f%���:�v��MKnܶ�'d�tѶk C�WuX�H�X�]���Ɛ�S�����{GfF�k�y���H�<�p(�0=�z��u��s� �ծm��:p*�vo;�p+K���έ����@DY����U���m�l�]�j�e��t>�ݷY�Z�sκ�9}�(n��N����Y|�a.����JtFU��oPq�sϋZ�ܱNݧ&L<����j�E��Ꜥ<�-��\c]	µ�OW�g������ 㖖�=G�wkv��;�x�af�ؠ���Ź� l��lC�S����=n����������;���x��]3E�Vx�4��cf�>q���Tq�����$s���v��`����q�nq���:�8��q�^������W��=�N}�;a�����ܤz]�b���κ���6('�1�ltG=s��u$@u���fŷ�ݹź�<�ڻ+����k��K�>�9vI��u�y�/�S<ͻsN�Vu+2�vy�O6�hڗ��\�wnx���Mh�!n�9^�qx���"�7X�M���)q����&��;K[�`��x�=rs�x�˱�u�C�=�'
���n�9C�=���[±��m��@�^��B����h��q�{��w��?O��!ǎ�h�S���i9s�vJSye�"��m1��pW�l�n'����p�7>)�I��v�d��
]<�;=<n��u�8� Sqs�ѝ�7X��z�˲7r[�S��;7c��ϱ�؃�Ŏ�=�]eĤ��x��e�����xm���q�uK��[�m�R[������	���U�]����]<����̕��h�z�z�z���7q����Sٷa���y�{k�'�5������ܜ���Y��@S�y�y��؁YY++%~�og#%B�*%au��}�u�F�ng�N���ێGxQ�U�hY�>�� �o�w�8��q��u��4k �b��!�ߨ6G�#�"�|���{q�^�� /����<�|+��� )��@�5��}�q �?n��훹﮸�n��x�:�rT����\s90�0�߿}��T�
��Xk��ݝ��A@�P��Z�~3~��_ٿOP=J��`X������i ��?y��Ǭ
��|��m��4:J&��,�ϨY������>�J�_9����J�P�J����!�|�/�>����G�ᖪFl�ed�����orpJ�o��w4in�0�%a�9��É �}���3C{��Mh��������!�
��Ț�}�p�:2VVJ�A�>���,�#��7��m�$�	�v�N�c�m�\�q�s9�;�'i�l���ܖ:诏�4�B"PS&D��8�||��T>*AID+s�=�ѝd�ʁD����,�,��̗��gPɨ��"����H4�-�����ïc�아B\DDĈ	�C{�϶��`����reVF�����ϩ:ЦW;�׳���N�oz����+��zhx�z�<�X-�1gYJ�Si�@^�rh��ˀ���oj��{�o�|M�Z��:���	!>��s�op?�J�V_w��C��A�IS����I؅d���w��ۯ>�.�<�����* �o��&Ɉ2h2 ���noW�$�B�?o�}��)
�Z0+��]s4��s7���
x T��YS^w߷��%e�%B�}���Ρ�%`C�l9*QALJ&C���|�Ϫ���}�����;��8�W��|6�>��:�YP(%@��}��@蕀^(�
;]�W��x����nB�V�E!m��s�w��
��>|����huu��@���~���@��2W���{8�����/4{���Ϸ�܇Xu�aXT�O7߽�ԝ����x�����~!&�F.�(k�2��m�]F�`�N�) `":wX�����f��uH�P���5��L���4in�0���Xo~���q�ѩ���vs�!m!J>��7�	��ƨ}���X �y�9Ϸ��������ݝC�+����7T�5Mi�/!��+����`�"<��-���+W��̡�u �X��w�{èJ��`X����������ܿ�g�Mv�k�Ox�Pܔ0�\DB��a�NO{��6u:�YY+,d������%Bĕ �@6��}�٬�������2�����O�߽�*�Uç�7 ��}����9D}���#�r~==S��V�^eެ�kx{��3�����
 y�}��:�d���e|��ځ� �/��f�L#&� !�ߨ�G��t�Z�&x���<H�?�g;HZR��[>��n
Ag"g���ì@9��W��!��,޷��'�י��*[��=����A���{�#�n]�)�;�|H�D
}�9��u+�`V�}�u���(!���m���̓�Q����s *�`m5Q�]���D�N���v���a��9۩�D�)�/���D�*bc�d|G�s��:�@��� ���8��(��D���<��!��+���{�<]��$�;�}�gRu
�FVJ���=��r^�}�i�Kp�s@���7￷>�#�wg�ەz��������0+���P6�S�eL���nH,��P���y���w߶q����ߟ[���5Lј�C�;W;�t#$�%�V���l�βVT���˟nMG�.q�M?�/�����k��P6�x���<��ۇ^�
�rP�Aq"e/�#�^�в/�9uw�~�,�2VVJ�=�GN!RT(����~�p�Aa��w϶p���n�~���؇�S���RӁ\5!�Sw�w0U�l�J���vNmnR|��}��Y��?���U���ͩFZ���歔&sj�w�aN������d�ed���|����T�o|k��#�hZi���X~��>�u��H	 c��A�x!q������������9H)ȁYS>���ì��Y_y W׿P���|;�+�Ϋ��?�OOooX�n��t2O��i㋧�)�\�9�sp���n|���\Ll#��[���+���oa��ID*J�a�����:ʁD�o����tJ��z.���c�����ZAH6�?{�����'gW��A"A�11^���K����D
�Y���߻>�׼�i�<��|�P�*IXS=��܇XtaXV%M��>�Ԃ�Y3��>��f}���/;��p�識ƚ4�70�	Xs~��p��R
����ii
���6�eAs�I�� H�$x�/�Ì���(���l�V��{�]9��:2�p��
�{������^��������u ��!Xo�����u���T���{���Ѭ
�Ϲ����|~��߈:)K=��w��
��C!���L� H`�g��BȰ@�����}��d�w߾����3��C�%a�;��H,:0�(���}��:!R%e|��op�������3�U�#wE�&�
&�:�7�b��ҹn���}�+�ǝ�;�=��8һ�qZ��T��u�ƺ���0�n�����~�$!%�υޫti%�֮۬�qu�Fڠ� [m7h�Ym)���\ {==��u�`�� �K�hZ�q\b͓	��D�׆��F�s�=�6����wDn����N�a�r�̷m�M�n)��N��춺�u�i۪Dql�z�f጑��=��3����z1�m=i�����-�68��
�Bv��m�Cm<wY�MӮ�mx��+�%�h��yo1�\�a�ۻ�q黫��=�ݭ�a+$�vzɀՐ����|�zh�ִ-1�=H,=���v�XjA@�����v���+X�}Ϲ�
q ".~�A3s־: ��#~o��Ϭ���*!�;�:�bJ�~g4��Y��.ra��}��7��¤�T�G����U�p�T���G� D���{èJ�����>��r����~f\J��_F�xY�֯�"�I���Y�N��<��Τv���������J�T����oos�i�g/��%����I�*Ad�+���{��P�7�Zh�s9�l� d#����%���:�ܶO����Ah��{���!Z0+O���r��>DFv}^|��}&n�/��;��}�Q�>� �yA�,�#��������Y����:à¹����#
��R���2v���n���%@�=���:��+ư,k��{�¡�R	/���̓�_n/��鞈�~��H�`І��F����k�h"4k������i��U)؉���|�����m�ܧ�O>��͝N�VVJ�2W�}��q��RT($�,����C�:°��5e�wqy���,�o��wt,�Yy&J2��Ϸ�8��>�+��+�hZc������>�v=`Xԇ�w��ܦ����=�W���n�����w��J�a�}�K���龒�]����ͥ��}���{K��cЭ��R�]��̪~f��I����9�H[HV�~����N T��~�ۇђ��ȁ���k��ߞm iG�c}L�V��U���i �~���0�*%B����6tgY(ʁbT�w���>ן�>��_����Vk��^}���i��a���ۇ�
���_����bA�10��~#���d%b�v6���4��YY+����J��+
g{眇R��*k���Τ�����u&��,Ͻ��yx��گ H�ݿfSF��:u���"Vߞ��8��Dx �~�������ӻ`i���o���9�*P@�����w�u��D5�~�gP蒰�>��l��}|��������":��/7W�{b��i@]�tuu�3���u��]�\g�����|N���rc�x�[�k��bJ�Ib�}����gY+*A@����p�R�0��_ߗ�-�y�����=�ہ̤�l3����׬
�:Oؘ�˙�C�@S�����"� #����>��n�a罧/z�g��J�IXS=�ra�aXV%�����:�Y:2�w�|-a���O��Y@����(�3$� ��R����>�u��!B�5��{�����(�p}ڶyUy+��*�27�m�YW���H^^�g`�:A������{O�]��D��">�������lT,+0T���.q/2��o�%�_~��S��R(&~���H,�%B����}��v$�=�<���5�ĢT��	>��ϧhPw0nX}�}R
J!Xs^}�Ό�%e@�T�;��:�X��|���p.�������^���HV����q��{�o����s4]]f��:�����8� VVJ���#���}� lE��km��������IXf�������{��;�����W�}��'9睷���9+����	y�,`$�	��H�ʔ�+sv{W�p���U�;���zř1������:�kY���Aa�7��H)�^��vq ��*Al�_o�@�� T��}�ퟌ��0��{�q�%H(Q{�=��;V���̦��Y����8ã
�;?P#���n���#�/s�É�T����@�V��|���p*A�R����ϓ��.��f��ӕ��O�E�$\ �Qd)~�w���gR:�YY+��{82T,IP�IX~�N�y�׿o�<a�°�*K[��vu �u����kﷹ8�������Uu�)Lxu�V}�P};�k�'�?G�	 /���!hR�
���>� )ȁR��C���,�+ꀬO���tJ�Ĩ}Q����.��L����,n���r[|�'�w}��<�F���=]\�w�����>=�u����BI?��gY*C_{��gP�IXS����e�5������0����7��¤�T��9߼�ѝ}���U��j���� `�@.�� :	R��_}��䴃JB�a{��~>����$�_A1P�;X��Qj�[��8wB����J�<�B��`���S��A$�Z/����l�s����d��y��pd�Q%B�<�������g�
n���'����pM����:��
�YY(��מ�p@\��B0�R�3	�#��
���6|(���}���pj��␶R��k�w�
q�@������xY���"<	�Foї�u�]H,9���r�sfir۸q���u�oa�%�(!Xk���gY�J" ^!�{�q�ȏ�YF��d�V�`X��}����H[a�y�ۇ^�+}��;�#̹��]r�w�~�gS�����g���%ed�9����� �RV���u�XV*���l�O�}}�|�z��q������orr%@�����t�\֫WH,?s���`z5!m[���9�B�����q������8�R*k�fׅ�YH���g��B,�=RnյL��͊]<�M!n��Ɲ��A�!YN@��#h�^�yz��-Q����M�� ��0.[��G,
ieW��w������}{�\�t�}%�����틙���{+�Zh�g��q�7��H�׮|��2�ۓ��;kq=���6��?_F�����:wj�k�r`��vMv뭂�:�\�5Ǳ��7�H4�NwGdr�l���琬ct��p�);Ob��3�!��u��n۪쥔&w$m�q음�����$:v�vI�Nܾ����ݞ��\�%sD��]� 7c����C���1��mr$s�W=��m��$]�
W��c����֐�R3��{5�|H+od�H���$%��m�>{*h�V�S�>������$��p;�����.mC��K��E]�g�����#OK��B�"��-B0�J����7���L�f� �ԝ��ي����{A*���I N�kd�ҫ�ƛ�|��FT��{v�5߄��k�&�6��Ξ���7G6����$�n��`�B� ���!H��|� ��=4f/j��v��L	g6H&r��d���f]�e�	�.u�2I-�U�[>k��@^4=Fqz�{t鞌��ci�>�e�㘈�0���Q0s�m�k��7]��':z��}\ϖcyB�H���ڬM���2Y@-��ּ�	��q���ߘ)3�Č�PZ��X��^�/yˮųH����[ǝ�t--�AUyx�ۆweGP;�$����L�w���z��Y�uKU�������W�����Hϧ��3�5��Z�^1�z��"D�
aK~U��2M���$��ُ`I��ܩ�`�n�$t�j,r�!H�*fĉ�o�l�tj��a ���`�I _NТ@'ʷ9��LZ�8� H3��/u*8��bd�a��D���7�*�b3���z(�'���	��� �Unsg*+"�/�����ڸ!@�2`�L��];�9sZ�F+�9����b���}��]��q���A'b"�R;v�'���OH�Unsc��=9�OJ(f��Sl�I�������P����0[ ۽�Ɋ[D��s�N��H;�R(H����H;�`!�s�w��]$Ld���y4	�ה�5����#e(�&�U9����o;�At? =�?J�t�Sӛ�tb�B���L�Њf4�Q�"iSs�x�d�H�P:9���ޙ��j2��_�'��.1,����� h��ڟ��:�8�薏������	o�ڬބx�Z�5��޶�ԑ�E�;8x�}r��3�]n:�O,��=� n?y���N%pd
�x�b��zg��qM��=ނ�5|c�6��u������f�J|�S}5J'yI�B9��4ԩ���ffG�F)�����v�=�ܫ�����>Hl����ڸN2;����v� _S��Ӂs��J���O��ǵ���~��{��Y�GnA�w
�B�lr薎�t2�>�SZ�լ{o0WN��Q3��Y��ew���M�0y9���+���
�־ݘ�ٸ=�����ux1��������ݯz��5Z�v�zv��{�d��蹧�^&F��l>
P�iY��{��Lv�x>�)��=�h�/L��%���q�JV�xm�	���*{��r��:9�l�/�����R�+��ޅ���mC4�'une�Ҭ;��x�e,�_�F�����m�����"��oxi��%f'^k�m�]y�q[wdDFȁ �U\R���3��ڰ��Y�?��*�������������3�=��U���3i�J�ԯy�������K6D+�y_�q���������ߐ�w����3m��t}S�����{�ƣoe�9j����;��sW�|�����Uya�|�/ˬ`�:�hĵR�
�u�V�Z�T[JTB�XQ��)Qml�ZQ[j�����P�V�Z�"�*W)TFU�(֣�m��cqșj����\�Q�b����bV�1%JʅT���Vы��G3rժʘʢ,�9E
�X��F�*���bV��ڵ��kTQ�5�Ue��2QZŢ(�[Ls*��V��Vb\��m��V��DR�kmQ�V-J���QP��1��V���2�����aa�ȵ�h���VխKB��j��U�ib�2��AUZ���*��TkT)q��[J�[�-ŵ��TҲ��J������U���kS�,L�H�j�̢��J�Kl�-l��aQH�1m�B��P��2�Im�[�ȣj�Uf\�ijQi)���R��j�(�YJ�ڕL�f1Vܵ\�nZ�J��VZZ�V�Z���
V���m�Ĺ��bKi�r�Q-�\p`����BC~��y��#;�h�LV�͛�=�(�)�4�gc����d��%]�|[���I1Yx��Wk{(5sB���	ۓD��F�@ĉ��`���ݲ	z�i���1�$ufРH$En�`��]��s��s�y����J�j`��4�����@jμ�O3���.ss��g�3pm�:����w�����৙M0� ��ט  ��ۨ��]�y�r�>�{�1 ;�0� ��"�R�
�޶$]DKqT�7W��_gd��)){��6AQ��� ؿ��b��oVW� 6�p��$����;s>� ./�݇� �F�̷�r�ѿ$J�v��I$��k��ڛ#���E�����;��W�te"j��Z%��Vk�$��㦅��u�ӌ����M��*q�[;U����u���&�m�\xfl�p���y%�������'�Df�`u�E��ׯ�x{��g䐭����C��Q���&�IRT�#���X >��l��r��d�9�:��/W;�H��rK�H,޹m#-��ڗ��R�,$�y���'E�ю�n�d�+I�yc���7e��y-t�KC�{?@O�b~3��︟����V =����q�z�#%�W�������6���^}0J��Q@��]�M0����&K��W]�<��H�5�R�$���0�IE���Ow�����ALA-D(!K,f��C��l>���q�t�s���@"�����=���j'*$�&`�a2·{�>���\p\n��L�:�`��W ���en�ר۩���!� ���m+�{6��
jjI�r�s�� -������ ���n�~H����$I���ߒuNNN.B(�,��~�ڴr�`�#���G�^��e��gr�g6���:��pr[�z0���d��6I
�.I�� {��}}~w׾���;�=v��2mˮ{up֡��I�m���3Ǉ�ƀθu��q���K�4!�L�Y�β(��2 ���la��=���n;]VM6u=�����c���j�'t�]��l�kD9��<2�2v�:zeS��vl7Iu�av%왧X�n���f�=�sǆ�۬
�{=v��&[�Ǵv��ն�	��n�.�h����W"�in��A��=^�{[]��-��݊�X�'�gV�r�~������ 2��������j� �nU�C
{����2g�ݷ9ꤎ��7d |���l0����X�$��ll��~���Ğ[�;��z��=^�� ۹n)��y�Q-U^a�tsX��N�V�A��*�J��Q@�Sܫ��AO7�,�@�,9�}{<Mќ���$�7�sD�~���;ЦSɒUR)�23|�:�2����a8�Ζ^	��m�6�
Mg:�SU�8{�j�zp$��l��ʓ!��"I��"G���p*/�mXeB��v��w�ۇ�}�K���Pd�캼t:m;��_�~,�����&}9�k[���ջz�Ԝ�su�C�[�q��cI�A���0�K��EP:��D[�ט \���u}�fé��k�}}M� [���/o������TT���� {�"3wB�P�0w ��g~.��;�/�W�f��N��V�=W�;�����yї�`�\:_<�ovM:�j�y�y��z�L? <=��ם��h�U<���$Ĭ��J W�Lc�ݟ����ճJeU@T��MCh{���""*��*�ӹ�Qy���8�� >��vf$ �3��t� �12	�Ug�����l�wF�x�޶�fm�DC=�owoo(��V~PL$��^�$��bʤK���|� 7{*�e�I�̐�}��|����kv@�쫈8���{?>��y�qvݷ�͹M�w=W�oktv�6[��3B*�DTviѢ�%4D�I�������E���" ���4�����7ُv� EE�6��s�&�eT���&"�纚LJz��u�W7� �t� #����Du�M
{�e�M�3� 	
�%�Ԙt{9�`�D{��`��!��
Ɉ�3�wUb&}��c�#}#�ؘ��:�K�3ZX�=�g����>C�#�*��1���.��+dk��%ɾ�ݓ���x{���o��F�wT��If������g��,O	i�����m��~�l��� 23:݀��q���َg.?����#��6i3�Q��	��	�%=w,4JJ��;��hs6�KߝD5�	��m � ���fB.G�.�1EQ
����E"k�*a�#�._7];o[\&���e�.8hh�3<����~���p�R'c�F�{ͫ �ʸh���٘:��������tV��� @#���	!�
͡!A1��	����߭MV�\lu7o���)-޹��D�{�w��6����;+�a����jfb�MULLC����M0� ��׋ �"����}U}�����M� ����7��� �!B�S�Q��sح�<�;w��@|{=���	�s����t�-�*3��Ǝ������j܊ݭ�z�+�<��;�L���Nnh�����F���ȿL�F.���Zʄ>����Aoג�K����ҩ�o���{1` ���۲���ɳ:���%��L�K��۲l _���b���u�9xx+�USR{*s7s�.8��0n���փn	����F�6���>�"tp��ރT̂R+>J[�m��]�ט ����t�Mvz����Gs�gy�a	}�o���H�D��M�H��� չ�,����wX���� ���V@����x�2�ՂVd�互�hHPLD� ��n�k�i�J�gT��*/rFf��{�<�(}}� �tm�&i9趲�X���A �����'>�n�C_�?<X ��須>=�y�VKE������w���J`��[����P��9�����*�gf`⽭�	(��7+	��[�}:���)��{ۤ7�izե~��-�F�l�ث�����Z3Wg|���h�]��!�%�!P�����\�k�4��x�g_�HBw��Fh����Y��Y��S�-�|qr���5����lXݺyQ}l���rڨj:}���w��w�M��F��ܙ�e^Lh���Wlz�ƶ��k�؝q\�˶�v}mϋm�;ٖ{��m-8��c�mՠ�Ş}�݄�|N�f2�v�6��Y_f�g�fVP�؁����Y��Í��n��٥�q��i����.6�=��RK�W4U���K�r��F�4�[=r�뇦�e�xc��u<��tI���L~��q��{\����{��8π�ݶ� @{����Q��.o&��ߒ�q[���-��0�`�U�Al)������ZΚ:+ާ���+u�@ �p�ڢ ��caۓGZ�:.���InPrJ�D�fFw��� �x|� ��8]����vL��wn>H�.+v�!�<��s���+6���J2XV���#�v	Ii���^I{�+\�P����M�FsW6���A1�'^7In_���SR���"�����_ �u���?\n�E%�UX夂H-ʎnH ��ّ�����5}�$��#�'��{C83ϐ�Uݻ]��#���C��Ū
غ�U��	I40�ڟ��>�s�I6r9�$���͒iM����-��
�n� ����Cʯ#�B��*�����޼�m)�;"��0�erq���<vla,*>��j�
B����.�ժ��?p�9Y���V��}촯��\�m���Ed��jˌ�N��y9R�{���K��C��>�us %��o �\��ΐ����h��ؤ�Ŏ5b
�_�ny��� ���>�@Ȣ/�o}�W�{w]�	 ��O7�� ��vfz�Jg�UR&�#3��0R��n�$���H$��m݄�
��s��W���y�f-�������$MPR���c�nf *+�mY�h=��8g��"ov���	��{�ɰ��;͊UW5�U�g����+�J��9��Ʊ�W>j��S�8��Vq�ؚ�<Hׂ(�=��Ъ�H���#g�{gl�<�v- A$%N�a�M���6f)�{zy� ������[���" �kЦ&a�6��RI<�1.�Ta�ތ����m�6��;��"��o'lM�OC� �U�Ґ�E)��SP���b� 3�M��	Pks�g�A7O��ԕ�t&���Ȁ�����f��OF�Z�jrbN�΢7�S7��8:��2�ͫ�Κ�:�jޜd� �o��'R����|B��ͦ	�[�
bB�W�aV�P���;�؈��x��  "�y�@|�����b����<��f`n����(!E��m�I���CiC��0�\HIe�u�$ߐ��tI,,��lBvr.��Tuݘ�BB$�<�OSv���'x��Ӻ6�{Om:�8G�uؽ>�e��?x0
����~�$�N7k$�C+��i��5���y挻۾�?oޒC������P�^�9�ٸZmT7����y��EWk�I~Y]؄IS�Z	�����{FT� 
&������Y��=~�iȀ	�{gީݞ&gu��U�ߚ)#��ԍ�`\�! ȃ&$ր���v�]k�聟�-��i�����4�/��*=E�}.l�E�Nß��^�Z�}�L�ݭ�_���8�6p�l@�Ȟ��:�7�p2�Mf�xJY�GD�*��j��9�{C��ߒA��E��pDJdO�)��ӏ������,8���0.���	��u1��>$���@�[T�@��������A[]s��Q���&3i�<2�;E�=�gn�}"<bA!f#c���2�����E������$J�ݷv\27rT�&_��@���#�Nw	E4�`#�}���A�rj�@ԝ���ල�q�[Zƀ�	}ۙ� }tp#��Y�2c��硥�)�dDI��p��9�_�^` �9u�۞�KۺSA;N�	 ���o� _v�buz��(��&��[w��x]�"�Wv�F��ܟ �){���
���b!ӌF�3]N��� �JU5���c��_[c�]�������H3rz�����U�Ͳ�.�{��Ó��դ"���s0��dk2*Wb�v�I�N���k\U'����y��4ۢ���NZ�6��L$H��f�&'���N�8����{�v�������>��r�R(�^~��`�-�ׯL�L��M3l��R��Q�m�xz�5����(�����X���[��g�>��4Ew����hL}�P	� ���t
g�2���4i4a�L�\�ۛ-#��bMe�\���H��až�\��ZGA��}콥y�ݾ.�1��q�]m�ɹ�]gw���/������lFҭʫ�U L�\V�D5.5�ߨ�u#�2BB�C��9ͭ
�vK�d�9м_�E�[�uҌ��j����e���j>�J��r9��TӵZk-N�үZ����+���{+�e�蚊Z�9�6�Y&�.�o����y�{ST,���{�4��N�������#���]˝�q����7��w{-��۞@_t���\G��>�������3u���ǵC��g@�����`-y�/���b�5x�� oק���1�.����UZ�f�gw\m��EZ�
��߳j�e[��	�ܕY��Z11��]��9</����3�z���J�Y}��T��U����S�9K�<��oe���V�pK.�׋�>ŋX:i�z��ٻ�\�@�b���x�5���bL~᜽�=w}Ӯ�9Bށ�|G�y��lR�*#^�Һ�a:��j��3[ ���v��G �bΛ<f�w(	��[ٻ3�����#6��O�"t�`�|L*ZX�h\i\���`��Qij++fe+c���T�Ī�["Ŵ���V�KE����B���V����TET���Uj�Drي��kmS,1��h�Y���
����J��m���	P�kZ"�+��h�*T(�*VUU�U�֕*��U2ʬ�R1�ѕ��U�me�,QeTR*���	iU�KYKk���U-+kik�cj¡kb�h�+	U
Ũ�[j�Z"�F�-ll@�`��X�Z�EeԶ����6EAZ²Ҍ(�J�TUU[j��J�EDAE��D����*Ucl�E���J����()m�"��m��eE��#R��ұe`���E����U+mZ�5�ʕ����[U� �-j��Q�F��i,ʋb��Qj%���cJ�QF"����TYZԢ�,�J�-�D[B���U+e5�=�#t��0��i���sK;>y�	{u��v�;]�\gq]GI[�7=ά/i�{d9ɵ�x��d�[n�J혭M۫cgqŮ[��jg�V/gmg^�=%�[d��ûG/,xn�Wbx�'��wf|��m���q�&�c[��Q]�/X9O+�m7OE�m�����\iȺ��9�sN��ؒ��ruVӔ�Hu��ʮ��<F�z:`wj��gX�[�lsδ�Kbys��v�s�v��\.-ӥ(��{}v7Y�7XM�RL�Zu�K����4#�W�.r� v[n������4+ln.�s؂瑭x�<[��+g��&W�m���m�TV������zb����^Ǘ���s�g���C��_C�ݔɷ(O�yM���W$�;y��7)��8��n)����;֦r�gnI���&k��K��Us�콖��ǀ�z�=�E���Oj�olO���:�.<�����W#�ٮ]g�������g���b��k!q�J��bK���O/���,v�8�a�u˓�3n8Ӱ��vѸ{��v�l�����a�ۡ�^ܽ��È��	�{v�Gh9`�{+�ql���5�v%�W�Q�Y݋]�T[Ǟg���o}o����F:�V1�d�A�"	[[x���>;u��x���.�[�kl3�q�@x�k�t��θ�y9�F!\1[z�s�p�;��&"�q����'��n�t��9<�`�4�E��΍��O&���$�볖��GH��1禹��2PFD�Ǔ[��{Kε�SCH�Ĺ��=���i����8z��fxɳ��\a�"��^���ݸN��B���aE�y�PNmet0�Gc���g�;mF9ɖ����9=�p�ۗ.z�׷}]���nQWj���c��1Q��.���:C�^�$,B%nÝ��J�pc[�q� �hv�r������Z��8�}d��-�U7x�M�;�d���R�/%��,��V�B�=���:2\s�C���n:����,8nN�p�5u��@���76�ir�1ьV�bj��]��B\]���v��}'����\�d��J��[�Ե@pՉm7�Aɻve���ƶy�Wn�F�j����<Y�q�j�I�3X��6�i�q���uՋ��컷�փ��{G��j�Sgrll���t��4�'fʏ���;d�X�ٱ��ïX�a�λdݱ��B��%��u^7��X�m�u����I&s��[oOn{s]�ѷ%���^��s#��<y8�h�7vͭ���w���!*dO�+%-ſ8$�{�ٿ$J3�Ή��a�Q��L:�B($���f �A%���%Jj��,y��^[ŘT'^��s�rA���̈�'��h�%n�P�f�wW�B��	&��U).#/s���]{m� *]���w�_ ��� �����N�"����x@���Z������{*=~���� ��������̤�W\PJ�l��s��2A����Bz��i���ry�;��c�F���w���"�[��DDy���j흛u���$��_B�4�"�D�-bm����v��z��[���y"�^��������tR��EC����0 ���L y�s�䯭pxI���L�ܻ���"�]�6�l_����J~
c���;�ൿ��{y�oՏ��N���w�Y�t�誽�[7״��@�E��]�T?��J,`l��ʒt��\:Q�G-�6�M�9[����x��?����;� G�������{��ڧ��e_$��" (
dD�E���H �w4� tA�x��y�{��7q��w6��b̉���"�<'D=;��)V������j$O�m��>�=�_�|R��2��*rc(RI��ߦ��i��M��@~���#PK�ןa�P�<d��|	�;����f�Q�����F���o\#8�����1�E$Zi �7nNzC<ۭq�h֣��lW��B;s��[q����ߟ��Yl`M4�ŷ��$�,7�#$�T��ٙ�T��ӘNT/Nu��>@$s��	������������  �l�2̆�
�u�TIi,}<�-$=�4�R,`3��PW^���/1����O���@��M�71�/;�`| u�]OF�̊��o_ǔ�>��D�ÐAs��4X�ƍD��.�\.4i��U���X�Xܕ�k)g����=���1�mRs{0�	�������_���rA�
^���@.�L'-�Q(�SN!gfX�K+7#�k�� ��応�"���f ��km�Iv�w�d�O�9܎d5��w�l�Hʞ�DGHOj�Q�Qd�9��4�/�����ﭦng���F��'����S�q�%��>��ֽ��f�磜���uu������=�����χn��\m�1�Ns��%���Ā6�Q��w�^=k��F{�ͩ ^wf`���IJ� ���6��el�z5w
:z��2�;�9�>K��3 n��$�3<��H�ȝ�!/lNzAdD��_{3 "]��4q��p��n:� @){ۙ� ���L)r�X"�D�!"�	Kq�"�F5Yu� �o7^`|�(ھw����ă�RH��*t�FQ19w!�ʈsU�UgdER�[9�2a�90�>�6����Ŵ����K_-��:���x ��B���ݤ�`��" (
dD���ט�D�n~�iΙ���~�[��g� �|�XY}ѹO!�ܫ��v��a��\<b�v��>Ҷ��+.�v�Gn�]An'�y0����h�d"	�"eR�NG>�f` �5��D�����Y�.����\Ѝ���� �|�5�*��
���DE��[�����J����b��y�I"W�Mk��H��u"_���TU�,3lL�:���n��A QJ�&��[HO6�%%����$�Ʒ(�n�Q� H�/]�i� �Ξ�!�[��)�S(�ECf���+$��d>�{�� O7��`� [�Zƀ@뷛�z|��Y5y4�"6�j�8m,��3aV盓�:�טKyU2"��)��D�$��G7���ͻ����;z��q��jƴ]å�}����*v?�ߝ�c�o��޾>�9�i�Go+wG{6{���B�r�S�{�����;	��d�C}� �p�D�@��I�M��SS�A���ַ����v���	��s����R�Sq�Q���{v�n�9.g^x4�:D@���t���4�Z����ٳ�)���77<��e���U�S\/%��Y8���mɃt�Ut��sωR��c�s�^:z֭Ӊ�1:��5;rnۍ����s��V��L���@cQ�K:ء4$�v�\�����N5�cqd�x��v��<&ڽ��Yv9)��H+=�l�)L�*���X�Ͳ A���9 @']��ςm�n����xN�I wU�f"~��D�)�ǀ�_n��@�0�dMr���aӷ�%;���Ȁ=�=c� ���b@�mf�3Ɉz�C�H]0T��2	.[�ÂW����Ť&|ݭ=���yN� �~�dCN�hy;u�b�&��[Bz�po2�Dk��� �����"!o[�n���#j�w�/+ތlBC"x���T�d̦ӭ���	 ��O�t`�.�ec,�U[�>��� 	���� B޶�ewgm�炕'�0fį(�Ϗ�%!{u�1�l]v�%�ǝ;mS��;pۅ��[����߇� e&�=�*��ND O��� F��m4j}ny������3�[I�=���
3��2IH��s���8{�� �Y��#��D�=�/:7-�u*��n�38�2�v�����8�R-��3�6�'^Ъ̫@M+�rE�.�S����έ���� '�y��A[�� z��Sk�^syݓ�Fxb̐A4LR��#7;s0 �m0� W��B����<��� �3�3 �o[w�[0R�d\4�z2�;�F��z,M<�H���wh�@��tK�FO�y�Ԓr��|��NJ)�2LLLCa��I$���\k#d�q� ��32#^�n�"����W�XU�y�O��V�J[2��"  ��>�!��<ܼ]h��u�#�I=���$���&>���v���b
��*�9!����m�I�����Dx���Q�(�~��ހ ����*\�g��)�*�@��U�期�ǚ)ɠESΪ�>��v�I$�F�I!��hA��b3ot��|+
`��eH�e�6��H$N�G6�p�=��˵���U���K�ɖ�ٲ;��j���I��f��u�죹����۱y�c���w�W\�R������)�F�H=}��N��<�����:�}��	/߭�d3��r/O&A�(�;ٻ�T��:���)�̶� ��mk�՞��ۥ�:��,�������H�L�K�wz/\$�Y7�٪�ps討��u�t�2ۢXI.��lB($�o=�Ŀ��~����QL���� ⎛�{�F|��mrn�e�%3���ŷUn~�����`��$���2���@%�#�pI+�7�wiL�8��ᱛ
͐�z��)d��b'��� b��h��}?H.&z�L�Cjj�D����h�zkz�%hU�li���˞с�%1�̂��	M8�L���v�I
î��nuc�π�y� A՞���>��ЏbiE�pC���d���G��V�v4��2���  �]�����}ݱuntMio*6��q3�Z��ںʝ!���������7Y���T(2i�4\{iQ��	��ȼc��1|��?$G�s��}����h ����vf  �kv�g���۝��=���Sc�՝٘��.�n�NL=�����9����Ɗ!Qm��.\k��u��E�'`�c`��v	�X��������SJ����4�� �gk�" ]��K�#2��Ȳ]q�Or-��$�VwfbՕ��&hR�������m4M(;"���WW����W�o���D��u7D��
�����6+6%�����OA$@�"L)�l){�l�I$3��`�l����(��;���egnf ���ҹz�RA1UR��nw��M�B�p���c��  ^�wl1���ۗ+�F�u� '���Ke�pC��f�����sqyY�N��4�جI^f]�6�/u�� @�:ܟf�G�����N�.��O%M,���@}����g巽nz��v>�2�ꊛԮ�7$�*&��$骐d�U�e:'oqSy!�n�ma�j6Q.k�=�.�My��1"P �$|�ڷ��p����l�����ixv�xꋫy�0�x�j��$8b{pv����ֈ�{V��g��-�\�������N�d�"��T�,�ӔC�)hO-z;����Ů镧�z�;E�6�pt�[k��n���j��v
�mq�h�	ܗma6黲'<�wCC���ض�2K��Ϯ��l��b�n�Ɲn�sY�l�ugGk���j`�"���w%��a�{g��M�`^\F�כr�jg����Bh �����{s0 @�o-��;c
3M�Y�3;��f ��������LQ�9a�я�K��3�)N��{�H��G���Ij��Z%�����r&3s�V^�Kye�D4)EIR�s�ߘ �N� K�M:��eDNߟ� ��i�gd�n�Q�T)U0�$���)�{=�(7*�n�v'�z��O7m�  7r��"՞��93�S�5+��l��h�(�PT�E���sV{^,3�S�(��];�{��>;�u� .���DgT�&����>v�=P:�v���#���v�ym�sc��s���v�>�1 ������T�
l����m��$ޞiȀ����b	����啓�A�m�P	 ��5�fP�451���{s	QI�]��J;��D7qP�L�y(�(c�0��V�{{�G�6�
�@3�\���;ۥna���I:�Ę��Ŗ���S:.�	�Ʋ�u�� 	c2���i �����~���bA�`E��wof�|���b�OH4}Xv���Dz��� Dfdo���^x������@#3�[�H>�=����TР)�1L ���lS���U$MU�7� :�w3D޶�-��Iۋ@'��7�A� �I135�k{.�h��]��zc�NF�z˿ >�cH	]7�w~Iy$��7'8N��G��(V��ܦ9qն��`��hף�71�s��`ƀ����0�3&_ذ�����z��mg���@�st��jz�S�³\�1�ZKf�n�$�/���*"LI���x�"@7z->�gU��D�l�uݤJZg��_��ټ�5\������O��4by!�S0�;羴���Xg�1H���q����6���sUZ{^{5\�\X`YL~�]�-���C#��2~���7w�w�Ե1����/g���[���x<v�wn�����i�[��ȱ3I����3ƥ�$B~464�^�/ksL�j�Wu����fN�ݺp%���ZY֏iPU��.��Ҩ��qw�˼�j�� T��\ӷs`�����9��Yvrs?����]���ū\����}�Y�Er�ξU���_S�]������F�sE]��_]��ɯ�ՋL^�瞚׆m \<�ۇ뾋������荙���ݞ�{��T�'A��k��u���gC��g��m�VJ������x�[�ڽ��3G�~��OD�3����&uѢ����(mI٣�.�"AXt�"U�Hۃw���;͙y����ɷ����F�.���*��䲝%)ٹ��w���z���0���={�as�2�]�C���I�����{�̹E��7�[o��5q�^7�ڲ�b�ս[{� �F�o���ؼ<��([<���Oo�E4��wt�uqZ�zN�T�n��ÞEp�����>��{���\w\�����;�yNPzg>f��}�\�8_y��3�w��fɫPqx\���ࡔ����Gۡl��6�)/e=�_{W۶9��(� �p\à���1�%�I�V��6^W�x�P)��m���O]�_W�ӜWs�u.�y��,��#��HK�N��:œ���g�!U�C�B�D2ߋ�����pË�S�����G�|W����V6�%�V*��T`��j�FZҩZȵ���+mE�1EQV��V�AE-�Jֲ(�(�Em*�U[h�2Ҋ1X��%j�J���ն���TB�kTJ�*TYR��1B�kTkDTQ�kR�
�U"���m��FءQU������Ҋ��XQ���Z1Q"�TmJ1Q�6��QbEE`�*5���[KYEATQ�mD���Q+R������EQk,U�@T�kV'R�0�X
�Tf5�.aUUpj,2�DAm��YK��1j��1�q����$YE���b����nZ���&-J*�Z��J�*�cY\LH�[1����B��,DSUR*.Z[A�-��-��c>�^~׽�  ?V~��@| ��6��b�N�5_C��>�E�w�d� /=��`�sv��ft낉5�s������ �E��TХ6��K,��n3n�o���Ki�]�@ �ۍ��>���#�a���k��J�7�<�vti��͜s�Q7	����cUNn:uC�%(JO��	0&�bf_-yywh�Dv�Q~	/����D����7�u4���٘�
}���]f)Dʀ�� ��
�<�r�jcf�����y��'ێ� �y�$�O=%M��$�|	���&f��Z���!���� e���a5�s^�<��Ob9 ���m&@�w7A��	�%4f�s7�n����3��?f�>n� r}�_�$9�빣�s ��,�3�2�(��ӭ�ä��'d�I����;���YSB(8�"�/R�i��t��=��R�Q*l���+S�lFO�O�'٭�����&j��M�?y�v����ݫ�1SW4y���Dù�DYݙ�Y
�ӻ�Ͽ�#�v�ʋ��;us�{I��Sv�N.5Oo]��,�;;���n8t~�o� ���<��6� ��ۗ� �;������ߩ=�o�M�L�����N�Q��	�q��r|}��� g+�G?~��~L ��'u�C:��� =;
7���դDUV4�F��B)�d"�
��u �������ݦn?fLSҏ^\DCGa�ڢ ����g���M�CĠ�?N��zr�i�1����@ ���� �c����w&Ӫ���qh#�v����L�HUR@��~׸ |��m2"���*�j��`uM��DC�_��� ��m3s;�Փ������p���:V��ʳʛpb)8�b�RCo^؁��sRѧ��9�ΝnfmD�SBH��#������6 Q��1�1�;4��<2���$H\ݭ�;2���KTF{v�d�x��=];8�:���n�n'�4rI���kU�Վr�R� �q����y�뱺�	ۯ:�uf�5��x����Ϣ�����[{]5M��OVx�p�sv$L��LҮ��P�qkv�y�1�b�ۮ��(z�WV��^�խ�yNN5�b�P��í�y؋��<���U�m��n..��z6��{[�vg#���{O�ʥ�]w#���S�'���\�-�C��|R��I0��W��|}fFp�%��Ł� F�c��o����4�繾?r��A$�)���;�z���8�iJ
(p�:��0�:�E��x�Q�9�@�����e���z��[�;=���
��bI�$���N��Ł� ���L A|�c���Sq�u� ��nf$�$-�n�\��J�EUH��U��̺��X��D�q�� ���� �t���{^���wf`
3V@ȕD�UDJ�pе�L����CN��g�2���;2#> ]Z�d ΞnHxWD�w��_������џb�xތ��W=c���=m��m&:�Q�z����Vݭ������R��������ŀ�����DDήcH+ۋN9Uz�t�}�v��Dl�,b|Um$S(��s�}��ȉ>�G�~���{/�7R�Z������6c���9�0��LC�T�1}�+zc7��ݲs6bT����#p�;���#���=�}S,X����}�v��F7�餂Ic�9� s+*��t�������E�P�S5*PQC����<�#���9.���E�]�̍��I�Gso�W�>�h�����$��`�33-���}X�K���π@���L ��sD�:�:��b��#�6�K!��"Q�[����K���Բk�&����m 7�<ܐ/;���|��쑷�9�L�q��6�$�'���mv/�#o/==��NlLn�Zi��/ߟ����%PMUD
�b��q��ozy�/;�1D)^�,\c.=|��DA���CQ�	�$�U$Q01��b
�/L�������%���0����q'	�VPBO��(ۓ��H�T���#{�5ȀH%��ϰ ��#�sꎜ�d<z"�i;��5v�&o��wM��qJ���|3E�5yd��,���Wv�a�{`���'n�>�/Q@>V���}�z�sr~	$��}��bA$!��w`$�n�(!1R�6��l�9gn�o�Ied[�$�!���� z:�����\�h;��ԇGaL
Q�&L̶�f]�D���Y����kf�wp�c )}��ω$�?t�7���P�F�FLI�Š\ ۷@F޹��mp��a�mv�]������#���}T)��~���g�
T�G�78�NO�A��b�Iy%���'-�1\F1��m�{:[jHK���(�M̢U�T@�\4�����A+V���3:]� ��w2#��ڲ"'%�׊����m��9	�@h�0��~��q%���LI$H1/�����u^:ŀ/{s"3���vҰ���'�S2P�'��K{�D����Me�=��RXv�K	 ������A�̜��zV�Oe�Ǹ;�i��}��,
�I�z�nK}����s$�|��ݵM������4*g&7b�2Ol�@�1�3�%�Ywwa%��42HBTL"J�)�����/$��fG0��z��p�w]�nlW$��7� �Ѹ���G���ԫ�1��u]���)\���D�0&I,Kf�6��h��-�Zvb� �N�v�9�6��|���>qk-e�?�oAā����	8�OX�"�5�]>���tn;�iR�Q�zd�
T�Ch*���Bލ���+��{u��� ��DD{�z�HW�gj���MM�3�#972�b�j� U.̻��"=�ڹd��'}2�Oo3�����H�������$Q� @J`�1	���3�f\?���[�� ��s%����.��]q"v��
�slR��F��B��'Ƥ���	"a�k�X��-n!~`x�� ���jH �۹��A�+V@�w.�Vv��i�N6���l�/=�
��w��j�m�F�Z6�ר��}�W�wpP-�����gm����V�RE�"B �@���/k��Մk��i���V7g]Qء����-n��9��wGca%	����{I��ڮƴ�ƶ�0��l:n,pE��9��AR�,d����z���XNgC�J�G�t��&$B8pu�������w6�P��:�ms;�kvu�f"Q�7iͭ�y��v��Lg����9c��S��vㇺ\V��\��u���Wj��+l"�vьs�5�:R�p� vC��t�b	x��Ѽ]�0����$!*f	I��Tn��D��fG0� @K���AM��OݤI�⼦j����߅"�^W��~9��Ĩ�FL�T�u�7xȦ��oc������� K����y���/����ݤ�&��JQ1"B�䦜k�R	}�y� \QH�߮
�ۗZ .̎oЊ	!�n���w"	3e@�n#a�.-��]m�6���ܤ�P�z�	 ��7�276�(I��mZ;	9�ؿI���٢rK<@2̘���� {���3suI�^g�˺l�i ���f�^���=��8�}�����e`�KI�4�A8��/���ûY��3�g:1%���e`�K?����*� �ѵ���Zr|���` /u����-��{L	7w)��/��"=�*HBf�I�Z�Ok~h�Y.�ydtk����[p�\^�s[��K)l�}���9u�����jp�W�5�+�����RsIe���	��Y��^L J_n�`D�v6���T��72��f��ug
I�Q��S3\�]�ݤ^Hl��XJ�*�j�h�gI$!��ݤJ�C'���q2w	Q�iR�CaV��m��)������ �7�>��"V��� #��W.i�{z��'|��Mn]�Cp���D��)	TXCs1��A-��2�I�αXO̽���]Z�d {;���^^O]�˺�w��=���[�v�MY��:Mx��k��d�>�x��C���ěT__}��~*�&��7Y��֒I!�N��$�Y}��6�F{t�h�����'/�I	��V�R��*|\���l���Gq�]���Voo>�  ]������a�'r{}U)͛��Oe�$)3 �eW:^:-$YY�E�M���J�Uy�wb���8��j�%�T��:�+���_Uw�mz�|��Z�}�U�ϥ󟧸���g� :��UP�9eM�$��fÁ=uP�o���w� ���� ���S`-���MD�3%
��l���S���;�eLR@|=�m2 �2���� K����jxP��lϒH^޶�&X�IDUETA�l A/�^a��\�f;�u��?�F_u8�i/���a����X��{ ��A��ęea1�G��-u��I̒l�9�'x��6��u�v����7����*�(FG!=��� :���	 �R�2#��i��l��O}Ͷ@F���O�?�NI ����=/�wr'gj��X��VA"W�V�2ǂDþ��"n����W۹q齝a�c�j���(���L7ݵp�	y�n1 ��1���z�@��l ���nf��A�
eD	�2���Z�y$jYnPY�M�%��y� !Ov:��SN�7s��	�v��y>+7%�
��T��4,�;�r�1]lE���(������y۷��<�D��c6��TP�S`n򶉨�&d�QUM�V��������g^U�1��DNy�ǐ����g� >�cl�����q����i�[n\{k����&��th}:CVq�{�{�{\`7j����߻���"*��|�SL %�u������D�EO]�V:qs~Yy��Ey({��6{�̕"�S% �qe�0A=V�:n�}�v�\� �J_�s1 ��[�XJ�F�g,�W�p�b�8��
Tԩ���~1�w3 
{r�` zDGV8���V��l��Izg]�i/!��ixƇ왉�Hʕ>._���N�(̙ //�� �J'��>ewK��=��F�Հ�,%s���K�z-K��&U}QC
{5� |�u?��8���W�K�ʞwfb �;�m�y$�����z�Z��cȣ���w�A�Ci%{�ɗ���~UȻ��<&�ײN���fb>�c>��r��=,Z�n�E��xh���7�ot��wn�fD��-�n٧ެ}�����^g;FW��/;,�@�������2����w}し�����W�5M:d|�:���-#U~^��H13�K5����%�<�%��̐�[�ֺ6�ٴ�(N�aV��ok�^Z�Dޛ��������.)�9k"�ˋ"�-���Us^'3V��6�`7� ߢE"��:��C齰{�{*���.D���3.rm6F�S�ЩE�U��{�7^�ؾ�o����ݏ!͗��m,wr��Sͪڂ2��2�6��۹�oQ�f�����3�I�7|���k �#��n d֍�j���ȭ�e� h�j-��3�\�,���W|O$��榡�V��M�yR�n��.�Xj�f�V�������hs�^��r���O���F��>��z(��'>:OZT����$yP��Ϲ؋�	������z{�+�&m�����|��`��Oa�`��z,�U��ol|�s�Ύ���l��||R�kD�4N�3�f������)�㷼�� <��-��A���_arF��;�r��w���S���M>b�8�Ռ���cVu����N�|���;#:���o?�b����@:��<����<R���W�O��UۦR��$��qx j��Oq܋އ�PS�o�:m�nC$�U�5���S����p���3*kD��	Vu��̳.�&��!�u�]7�_)�n��������8h�6�c�o�{f�bw��՗�u>qy�뿛�{���춙T*�q̫-�Z1[J̵E�,`���2�C-V�j���p�c��8��f��pʕ�-eKj�
�6իJ�(���Q�f(���6X��6��A-s(ֈ[b,��2"�j*&4q����²䲈��1Yj�A����%k��̶VTQKl1-�PX�lX(.4c�����k�Er�Klph����r�Ueh�j�F@a���J���)P��F�%h������"��q���Yc"�T��E�f[R���S̦&e(�1�PX��Q��r��ڢ8��@DUQ�P���%QX+EQU̲�ʵe�0b�30�r��Ƃ�TZ��X��,dL�1�0��UE�d-A���n��<v0Ʒ���2��ɱ<m�ף�6�ۮ���f�+�Ku��m��e;��t�q����l��.���rv�@ލ�[��ֽ0Ɲ��7� 5�PWj�ZIŶ��ܞ$� MZ������g�£�nw\Ӹ`;o;cg��s�mk�;�[g�k:�5�*�)z�ў�Ƌ�y�W�ے��S�Cm�竱nv�b.oVX˷k�c�����A㱱뤞�q�nvp4,�'kz��ޝQ�]9�sf�p�u���ԷsPa���03#ی��5[q�9�pE�]��k{-ۋuɹ�T^xlx�I�;�� �W0^��s�6���C��ՌH�e��tS�v�2��D�y���$ɫ��Q�ۻ8�i�1�xg�r^9�fv�'<��b�v�/��[�%siEء��q��0�][��;]���I�qP�IA�T���Y,Fpv+��(�l;�v�%��b(7V��I`�oG������/Zs�݆ϝ�u�=�q=�F�ݗ��!a��Xն+�v�J�y�W��g��v��/�/�mɯ�?[v_��Q�u�1{O�}�c�V�5��#��iʦ1͞=�LC�!93պ8q.8��7[nS�m۫�����]�M�����T3��nU9ɘ�[�=�����8���{6은�B�Ƌv���om�8�ӹѓ��}�}K�:��;�m����{v�������ٹ��N��,�gv'iӬ��u�����5N-�<�'!�n��K������4r�:�O�]�-�6��y���;/:&8�*���/]���ծ���[���=�q�r�d���.2�[)*��۰s[v㪮-�� ��-�3�� �۶����j��sWEvCR��nEo⹫���V�[j����sT�(3���L;mt�f�ӻA�t�&]�t��=��t��'S塮�����㕭��VT�󭶙ۗv
 w=k�,)�:�=���K�$�L"vHT���8�;����8�l:���.�.�6�;%���ڍ�\��˭y�77�����P���۞����6�lq�鲗h�ǞÙ�t���9�Ӟ�Y���n4t��v��fZ�p9!�c��� K���*y8��-�Ի	�u��=t�CB�U������7�ݞ�sɧ)�{(.��v�ѐ�{X�k�n9�81�<u�oOβh��<	ۆ��-�-��ٍ��8��\��n��)Ijځy��\fݸ���Nh�Pה��8=��c4��hN�a�B�A_O~�ߑ5D̔**���y�ϰ >컆/_u�a\��n�������wa"W���m����	�UME��S`�~emv�,�@En��#��M��p�䖉��y����p!%B�HJe�}�� 5�U�_E�Y����op 
Ͷ�$�,}�߂CC6�!B�$ʹ���s��̭ڽ�{U�hw��0�k��/}ٜ߬��W�;� �������USRET��\��}ӯ�"@������e���5�
-�;i <�u�$D	K�vf ��ńߧ�ߟ܍v�<����u�
⧄���]b��}����s���qã���y���u�Z
^k�iG��lh ��fDU��$��ˬ]z�7�I���v7� �uϑ9{6aL&RE�jO�������).�_uM�ڨ���)uF�}.�,m2��3
͓j�З���W;�i��WF���k����4qa�SdB��]�/q��T�ٸ�<����_|�  ���� K���@�pZ��]�\c��N%���`�0��~�D%KH; ��/a>T&���p�M��e� ���u���	y���}�%H�QS"��w���;/|��Wn����4��){ۙ� �Z����z�?|l�$���3�8�E��L#��3�����}M����T��H�M�"��nf �_[g8�u�����;���8(�ѫ.m����x5ɑj݌�I�M����B�NL���~�{��*�5f����gZN@���������=ؕ��}9��F6!��;޻&��R���"b�����)~��W7���3�a�	$�<�$�N�o��L��I՜�=�뻟O��ټ��j&��(�*������\���6��d~�5������I��d��|Z��;{��o�����~,�[�s��^r�~{
ٚ9\n��Dm�8�q���I��a5D�9� ���3 B�|��;�1�A�q�m�!/b��g�z�?�Vg�}�@W�;a}<�t8��~	+����G�Ҹ��L@�p�ny��k���zr罽�Ȯ��%��dF|߹��G����}�پ�K�]Q$Q���X�/ M�����W]c��,z�b��R��7tQ��ۃ�n����7��"�R��M�9�nb� @����$���a��վۗ��������"�7���	�߫m�������}���1ڗq�$�H��D��WGS�*(̭��5u]����B�HP��d�og7� ���y��A��Vi��|^w� !M �#���Ԇv�h�SD�ԕU.'m��+Ի�u<����^ֱ�D�w7�3.���$��ECS�3�9�7L^h:���»Ũ��᷹��T3iN]��4Q���&(p���+���u�X��
��J��0�w�+�sl�)=)UUE��s�4�/{^,=���Q���/o��6�y� @)~��ς��O����o����ή�DD����k� 鵓{q]�=Ӂ.�����L�B�=]�����|�۵̢�c�������>��nD�@)~�$�������q7;�>�o��[]��!��6�0��==���q�������UW��  �}Z�����$�N.�S��Y�{E�~m��$��!��N��� ���g�ܮ�Z�h���6l��� �g[�H
_��ɿm��)�2�
��#����n` oO�� �����@
u�y�z���[1�<�w��)L�1UR��[��y٘  S�m��J���y۝�`%��lh��K���������f��@�S��r�$���D�\���W�!u��eV������9 �{��}�]д�Fw��=�Ys�"�����7}��g��_���k1�7c��h����z񞘼�^KX����)�o��؞X�=⭎y�=1paL�k�\X3������\��l���l���':��prk =vK����I�]u�WQ�ٻ�w�[��L��v���m$��'���k<l�&4��p��&ӝ�W�}$9��a�ma��\v���x�Z�T�q�ǰs��0Z=�)�5��P/c,V�u�ű�\���l��뫀ݮ�]��5�u֠�ш��� ҩ�#pr�8 `�@S32s���[�0��w�I%�k�i�$�ؑU�̈i/{s0��L(TD�Ȩpŝ�w �W�x�9�ǻ�*}�D���b )�Ͳ *-/Ø�������'�s��x���1O+y�l�a!�M�Ik�l�t���Nn8� ��vf@�;����L6�$�)����^��_@�x g��ϰ��O���Ϻ�ۇC�LQ�1Q��Ā�r��4�����B��� <����>jͺ����7���q�� <����S��Ϣ����@R�RD҄J�J�
r�m	s�U���p�\���^,���������Jd����5R�}o`|����Hc�_�r{{63,�������� �������F��L**��H*�SLlk�ۖK��
��h�W��5�U��#v%������M
���^p^F�"n��H��shSB��uyR�����^�y_��;'�'�@���퀀G�u6|������wS��]�`�0������y�"���� �̼�S[{�7��� ���j�<���ы�Ҫ�59~W��xr�����7{N��I%���� '3�2�>}մmLo���ͫ���j�j�3J���v�L �u�;�?Y9'�Km��O~��$^t��D���Y4��́ӆ �QҼm���/D�*��Q����!���Ïk�ȇ�gr���k�=�c
�m�g��&i??u4ȃ��wfb�)�"���4��'��8��� �	�l�m7�5��b�K�X�N4^[Xg:��T�As�ۆ�@)��������h}���z&�f�v#�E��ƀ��c >	�v��|����X6p�Y�Brt�nх}Z��d���ć��΂�H�Ž�����Q���oN���b�mk��S���*!��^�ȸ���\� ���C@}9�٘���TLE�g��7�Ȉ�Ѥϒ魫��@)���π�o�j"}��&���1bɘ&�L���r�����H"&7�n��9X��s�@N^[�s7�1 �&7�mX{ו/����߿\WB��4�Dq��f.�ۂ�6�:��8�b���h��,���X�������E��q�b=��w� 	��x�>��tPW�T�"��6 >��ndF%��k*U��UE���V�A��u����O�� Z���0Q��v@��T>9����ol{�I��}��-��a� 
k{.���۔�$�+�6�'D��@>�����EF���]����@���؀'���]�C���0-�8�@3�����Q����L�M{��z�Ĝ���Γ���[{�ެpg�o�$p����s[[T��- ��uS�6ve�m>9
k���p$�A���e�H�2��"PJf"�>2;�o� A���m^>��}i ��o�1| ���iY }��DD�_�;��oʭ=n�b��N�]��C�����h8{
!�շ����~��˖�y�?�#��n8�Toz�V ��n�)�oa�mgӛ���|*;|ڰJ'w�^4�a6����BI֍�֞=���Հ� ���M <�����]@g�a����W9��$����!L��TUQC�������U���@����ێ��$�2{r��Z��-����cM�l��6d�/}����Հ���c� tcwQ�_m�i@�3{3trv�8l;�Շ�qV��D(�������SOe��H���wh�� �:��@x����׽V������_���C߲�
a�ݑv��L=u;^�N�%���P��.'D禃S�n�h^���*���s�^0ȕB)O���cDOa�I�N�xѹ�ͳ�݇�,v�ԁg�e��Л�xv��͟:�<j�N&:�s����k*�n�nHOl��+�&�K���Z�Nt�y9.7Dy��g����`]v;n4�kgOY1s�͓��u�9�w����뽧�b^=����]��È:��r�Ȼ7Wg��ٻ(s��x흆�[F�9*�t �A�����Wrƞ�9��J`8DҲ�kAkv.�{8ۢ.��L�$FwK�!(%3U����n��s�� �����@�ḪkBa�e�
L�l
E$m�����b�M���
z���v���{=��'�x�� K��n }9�٘� ��ə�=�X�n�8�^p�#��$LI�Q3"�#�ޫ����y����x�ƍ���	/$�<�d�X���I��#^0^0�,Ʌ	��j;�߸]����up�D�ݙ�����G���\hoΛ@}�w�DUPUJ�E=��� �&;}n����W[���\����lh�����@ 1��Շ���+��A��X��DbX�����,6ٸ ��w��f�W/lFGk��r�������}���1
��UG�)�Ɯ� �}�� 
�9$�P�s>bp�#�%��m�7`�CD��Tʡ�FGg�������r�Ɯ��mR�v���T�=�w���Wt(y��[Y5ZA�/{I�͛�ԣ\�K"C7�]��!Z�
�3q�WfԺq5��o���
}���1����^����<�(�2��A`ŋ&bf�%E(�4gf�f Loz݀T��wFOD��e��'su� '
�d�B��+Ƙl��8b���x3J�w�� =����&��D0����A�W�H�8oY��/e7�vKݖC�E*�������D��n� y�y����^X]���� 1��j� ����9�w��.+p��0�[/nz}I\e�&w8�y�����<�Q"(B�_��_�&AE�e���������Lv��V  <�����cON-�k~��JI$�=���~__�x�l6��N@L�#={��` ���/�%Y�͈E��-1}7#+r2-��I�@A���3 ��v��I���r jK1LA5'l�V1�s��knpFѻa�m�%Q3y�}�w"ֶ0˫�4钙�H��{����L,[�ѡ����Y�jԼ}.eAg����z|��ݺǣ@�i<��^*/�+���p����gbCCs���[S��2��(}�H���{�s�lv{i���y	�����[��@�سvx��K�'pX=���6w�����9
����B���`��׸�\�zy��{�m�V��7���!t$��(�o�&6�m�z��9v�η5� Z��N����ݍ�!��;WP7y�>��/q�nv����]�՘�SQ`��r\���L�h��4M/eeΚ��f�D�g��>Z��'�w/i���3���H�j�ݤ���d<s����tA�SCvh��J���vo����q������owm$�=��G����W;��s@�l�S�Z�����z(Z��{��g�O׺1d���PᛧHȠ�����#^�{���,T�Ǿ�\��&v%
��(�K����|�7	�Ϗ9�ZW)y6�?r*�W�=��a���D�����qn���O��o�!��|d��ɴ����H�S!�޽��G ~����0��*��>}�cՁ�l���Z(��V��� ה`B�d��up�/��'����H/&�n�;x�ȹ�t3�"f@B.�\���`�$N	�jP,7�T:���@�Z7(\6����}5��57=�z*�Źc�w����2����ϗ޾?U��n�[�ZV�aj�W����Z�e����c�k\��AK���QL�na�m�DL�0Vҕ�r�1b�kF0ER�[m��V���(�-Ve-h�F�q(�m�i���-J�QY�P9q�eV�c�i�,���U�*e�3+[l�Z�PDUqĘ�-s3(�.aJ[1�5JՖ��V��U��QҲ�ն6���-*�Z)Tb�QF�&\��Um��+r�̣hT�3*)���q-KP��ƋĨ+i`��kZ�Q-�m��Ȭ\�fe�U+
���yM��۔��m�n������cn��{'���Kl�e-Ei���*̵�
�%rՋD˙p��b����9E�Vв�����Q�5�%��&7)cTR��-j�5�����T\�UTZ�Rܹ�U�`���U�V#�(��գ�����EJ�X�D2�U+A��̪�
.P�Z+1��ƫ�*\�%kUSJ!Vܡb̵�[V-eq̰̱h�k3+�qʵ%q0����8\ŷ+��?S�0{����U�ߡi�,\A��*�f�
��n��k ����	 ��n���լ ӏ�2��!�_�p���úl�p/oԼ��h3�)�9�:ӓ�N?s�$�gЮ�H�c{*Ia$��9�B(%��&��1UY��?���?9_۵�r��n:�b���a��Im��dޏIw/	]�ã���῭d��TC�a����Ӷ4�@)�ݙ�b�����Ay��D��[���H�U����-�H�\����٣w}�NPI���{�� �c@|���I$����웓6��;1���$G�D��[@�ο�� �|�^, g!��춪����E率R@�N>��$�aia"$�0& Je�=x�I̪�����s��D?\����'_�3 @~({��R.�I܀��Ub:���z��q�BMl����3G��o��	�w�m�^�4@s3�ӃG\�Ȅ3�8��s*o�[3ת��w�6�9*4q߀7.y�&FL�1U�����ŀ�	��[Vz7x���k*���c@7�٘� �����w��NeKqUߟ�����'w����+ok��4����i�W=l�l�������>{��P�:8��A���Ȁ	��<�@|�t�����*���3
�!n�:�_�QY���n��u!T������L>��9����ȁ��w�Ѐ@}7���@|1��� 5<w:w�)��j�k������H���w���I9��v��R���
����mt�ʨ���$�^���l���I���_�"}"&fK&�i���/�cb1��cϰ�	��� �����q$�-�4/����&��,gE=?+" gWuD�)�襉e��f��$�Q�ܐ|�;����S��u�w�vdI��˿�w�Ƿٽ�s��:�;=o���ռA��g	x#�,5�<7�o��!i��{ynѹ2n�9rCH��	
v�n:�;
���u�hͳ۪wG:xn;y\i�;a��Ω쵸� ��Fx�k��<'����#�S���y�n5�S��܊/,y���#q��K�i�ma3��vQ<�t��m�����\�ť��lK�@����Dpw�M�xۓ���̞���Ξw���6R�w<�v���=�^��k8#��N�.�4dyjƗ��M��#�ջUy�}%u�8֪��k�dі�q[�Ŷ�ݻ;�`��f	��R�T�r9�n8�>	!� z��@�-������y�ȌH{gJB'_�)ET�D��r����nF��C�}|Nf��_��@ B::��Ae.��(�m9�X e�Wq���Y����EHU"�jh�pp��@A�=���@|B�S��U}W� ��|�;��^���R����l�d��߯{v?2,��� j
����|\�\�^of^�:S�~u]{.	�)�\ؔ��Dz�$�􈙙-�)i�r��&g;���7y��b�h>]�k��gu�" ��٘�����w�|�\٧�h|�֞+eLPs����k��z���݈ۖl�m~����m��&�U�y��DDm��:>�����>��s����a�=]OԊH�-�bR1b�RLTJ�����vfA�O&{ͫ6y	�c�����ݼܪ���<�w��n�ו��3�~���1�)�z*ej[cB�"oME�R��5P�SͬW��x�QP�]�]�X �^��r� %/7�1 �V�FuT\3��P�m�~��/i6�L����fFH ��� DK/�����<U[�� �w7D���f�����53110�Pz����%׬�E�S�V���@ ���� ����V}�Y�P �͵A�|�PTʪ�TL�'_c���d����e�񴄃��p�&v�a"L��KC��F9����~r���Des>�g��=sv1ڡy����e��b�q.{.�U�����}���^��߿�
cƝ ����g�Qݎ�&�ݻZ�M�f�#l�9�`)~����xZmc:&��� .���<�7�_�t �wf`DGv7dDE�\^�'8��|�x�b�R)��*��Ǿ�q� ���v�C����v.�9�s�F�BM�Γ1�fL��íl�]�a�z��zYG���z�L=��yDw���X��r����(��7L�6���q�H���n�%'�ܗ��Z�i&p�0���O�d�����)�q(��x�@���!�>Jqw8��bo �fkŒn'{n�$=��ȴ�-��i������&i8H��S|NEĀ��vfb�>*;q��� N.�ǥv
lΊ���tȘ��@P'���-�x�n׫����z���\ru��ۉ:��>�o�9�-ɴ����[����}�4�� }^��,UG����)�{�^>�� 
Nm�) �j#��$H����N��� ����d�{�~�� ����$gu9D�&ɝYע����儗����0
S0%2l�]I�$L��~r���'�����l����7�� EG�D?�+�u���,Y*E50�U#���M�}T����r�D�J��S�^VO�� ��g8���q�k+�9p���]���wj)T��i�B��c*�z�N�xx'#��g�X������^�̓��ق��u�)����v5�y��lG���"y�������&�9h3N�������{�YpN�/J2�R+y�@|\w7�N=��Sni�8'd�����P$�duk7C��F$���gù$��7`���ӟ&Ւ�������4�L4�m���u��'�I.��P�"���&�#jll�%t�-=��X	����Xw�gIc�6�0-��^ nB����k��R%%:�j�%E��� .�t��y���ڐ�&[����B�� �32Y5*��r���Q���` �8��;*���ΰ 
ӵ�-%跽vM���K	��Q3"S,�}��*�wY*�� U����λ��H���������	&o���4�b�Q150�U#��vf���]D�l��P�ɷι経 �}�v�+�Ov91���zК�.��޼�'=��>�v�<(�	���T��p}�
�����'6����(��oPc;5F�U��0tGFT�'eM��Q���!��i.���6�Wk<�kn�pa�i�2�֎�m�z�+��s�z	�O����^xcw.<n�f	���]��]��	g�N�Q=Y�5�un�S�nݵ�u��l�n�ѣ�[����֜as'@q�㫜Ӷ9�z�g�=���3Z�0l�`x0r���^n۶�m�=��'ɶ�������+5ف�r���k;V�q雭����5�p��{rv��s$�;���%�������J%|��X�	��� ��r�=N�NLΜo�$	�������*h��L��oa��z!	~��y��v�=�y�7 �nf�Y�s�Y���_�"Wc��i,&�FL._׻�"�z����> ;�X]{=*����4 ���ς":���A}�r,J�0c��bO���{e�`��I��ŀ\������Έ-��W��3e�����6���
�2%2«]��D��z9�č�N]fdLJU���I$��]��D�9�Ԉ�v.c.���񾪡�݆�k�7���&�_o\�s=,痰�!��IFP��7܆�`��Lµ��3=��#>�}mP �dG����+�|�wwĒE����H^졠�*����oO�h9%��nc�.+b�E��������y��N9�ѵE^Ћ�q�]��E��;��/^�nݏ7��N�s�P�r��*'�~���׻J�\o���` ��w�X |W�y�y"�Qb�������'�u՘�&"&d��*���3[�_ ���擑A�}Om�������z��� 
�O7�+د�����m$v{��wz}�&5 ��[��� �ms���f{��Qg�q$^�ڃ7�J	��3&�$��7$��Vg;����x6N�U	-��pI/�s�[�IE^u�<�]�Qj����%�7��l�Ā��p�Sv2L��a�����8�E֍�v����;���N�5u^3/������"	��f`RK6*�r���Ȼ�� �읷!�DA?B���Cy��H.���c�)ؙ���<�Y��D4�Sy�����"4NBFC����?�����)�gP��>nO�A8�[�� �{/0~�A��K��ZmN�[��C�ͬ8$@M����0�[w�q
N4�4b��ƒ1Ņ.v��6�*�^�+M�轷9������� ��fbw/"jh����*eL��.�z�8���	�uٻ��J��?��"�Ϸ3> u��߼l�L׿M�XD����3�q�[I0���b�@|��n����,�N�e�@ �}���D�;�c��kg����ӻ"e�܄F/I�:�{�s��Sٺ�WN�2��� ϡ#$��aj�"&fNR��t O��ń@��uOy�
k��U�ZD��mQ �ݙ�b�"��5J�����n�v��uGӜ�{S� ��̈���ڢ"�^���2f�ޠKL,������c3��/֐H���O�Q(%u	f��	'�sλ$���u���ng������PNW��o�����7א�J�s��D����"��^ǲ��� ���.�42n/٫�~_3T]��y�x�no��y8�5��q.�Yt�u�I����~��Mϻ/���v1���vww�ۗ�51J�&�5ES��;~R	 �qg0�T�1��q�I5n��&�WF4K	��NV�Vlד8��H
}��^��gN���<]����vsJ��ݹk��+����[G��3�,L�-���\��q$��m��ڐ +�u�@L�p�)�=�u�~n#@:��j�ȱbE}
��UCh'��IO"OZ��՛��$�����>+�sj������^7;�~G/+=D��PMR�p�.3��� i�ܠ�	^lʊ��L�����w�Agn�^�P��b��(�&a��|�%�,�DUڠE�$�w['��o9ط*��5�(@6b�9^XFD�3&PU���������<.�/�!3��T���}�[��o9�C��]C��f��$".f�'4�Q����a쩫CU��F�Ɍ�F���gaY!0l`��c�usQ� �;JJ�/\/�s${W�]��4缵��#���D����.��OB�x��X9��_E|6��<%�M���w��bbv�D�Э�ov�.Ā��3�FOg�qn�}<;�b�P�{<.�i��P���i�h�W{
2�� ��Fƺ��I<|S��r��;�Z	{̎��wq��F�����,Ъ�(�XUS �Q�����7�Q*/5�N^�_���h�\m�������I�l��{�G2�Â�q�=�v&��,�b��qb���/�7'���I��+<�S9�|d8�{��_����=��<�+ج�i �]h��mD���ᭊ�eTN���	"˚���{3b0-�[1�5��C���y�n�C��u�9D~�^�VÓ�ǹ.}�'��FT8�\;|_������ʚ��4{�mkW7���  v	�//>��RU�e���3��l})߇<��{���$@Hg^����q�q�D>��{�^��efmsQ���,�ͻ��]��ԇ�w���,[�c�zn���8�[@��[����Qyf2� ��[��U�w�o�,Fo��8`5��wQ���捍�a{\�1J6��� L,Bk&��
;|�;t݃ ����vh�l�Re�䇧Pܹ&���/��=U��[�ח@���AݟnYdl�����tcI��/h���rf��ܕ����R}�3E�[�:�V����ب^��N����[���T��e�W2�*ԴB�*W-D�pY�9m2��c�AUJ�1��3.*Z�E�3-J��Q�+��E�
ZQV"�U��V[S�EB�e���DE�L�QV嘆Y[�b����q�Q2���maX��nYL�5�8�\�iV�T���HŬmX���3#��̹K��̵*(��R��P�Jʔ��&\J�)��9J,T��ʔ����Ա1���X�QDU-�ƶ[A�2�U�fX��-i-R�\ʠ�bZ���U���i�pb&[��nLLrDbȣ��\Je(�P���(**%�ڌ--b��̨�fZ��Z�X(�Pf\e�2�TU���ˆ	ET������)E.A��ALs(�-b�F(�mc\�K.[F�R�J��fb0LKXԢ�iZ�X�)m����~=��x�p�{R<c���w8+$�N����t�F�=.���%�ٮ�rs@x��O�r]�4��&7%�uՓst�vc�ṛGM����r�U�㭮qq��;s�P�;ʖ�&)�ہk��8����:�E�:y��8M��zx�����v��uǪ,���X��y�J����`
��H��y���W	�㹳�+g�k��M�Vr�n��ލ�����Fxmһ��:��65��u֖�G>�n[��c��^���bG9���x�7;�P)�ٞ�Y���;vص&1�6����]�6�ѧ�;�ZD�����.�ݸ� sS���II8Ǧ묝�:yDx���&S���E�βP$���b��{g�΋v�kq��׺�ϛA�� ���[Iʂ����-����m�ݮ7&^��,uc5\N�ۜ���܍u�i��a��v䷵�[�:I:���Od�;�vLB��۵�[�.�s���d �{�mu���=��S��6�η�kǰ �M�]n����k(�y-t��AW]fBz����cd6� ��f�	�Wb�\�&�Ƨ��'`����Dlxy��O'.C ,s�s�t\v��F��27C����F�;U���'F�n�6:��O[����B�qY��pwHg�WS�-{����DR���y�,S�ݔ[s�qu���y�Yӌ�[3������s9׈wJm�v�h��(�'b�	�l���KG�;v��g��nl�4�A��ۦ���F�����S[m�>k����y��{%�t��Nnݳ�ɼ�ga�Q"{U���^q���b�݃:���$�w.ϰ5���g��b�c��b�����\�"�g�n}���q�OE�w; ��غ[uˀ�3�[�m�Ϛz���Z�v&h=sx: �_5��eK=����v�s؜s�l������uh\���G4�E2s�� ���>�Mt�4y�`x�0k��t&�u��]Z]�=��f����8�.���7m�� Jz��hN(ӹ�����[р0����Nh��m���!�v.���W��N�.��tn1y��6�q�k��C�Ռ��l=�����k-�\��.�r��[=��۵ս�5�{t1u��\\E�v�;��s�:�z�yN<mf�͎]MIۗ>{nûu������\��Y��h��gv�n\9��r�:c���v.;2b��P9W��/�aDZ�NȖDbmv��'m�t�bXQo�p ϯ_�x	�M����ͭ �o:���.Bs?I,�&6�[$l�2��!3����<"�u��aɞ��$�coy�O�>V�v��B�y�F#!�zDO��3$Lem_�cΠ�$`��9���)`�{<A�����[�oā�0R�Q�����lѾ�gOb�峆&7��\VsgĒ��[�$�3�o)�ȲM���*������jhXpI���0�=w��G˯M���7W�Ɠ�}͓�V�kd�8�]	-����f	P0!]Ŧ'S1�����y��<^�X�Esq�b봢)cA����,�Bi�m7𾞳�0��i��A#����֔ª����T�eX ���ǎ�10d��0TL��<a�H��vr�fy֣`����k:�]�m�.L�ݻ�(<����Etzh�f�j�(UD��o:�K���Me������������2	 �-���$��S�s0d\[����7d�pk�3�,O-��S��d��~�` �l2`�@͸��|�I+oy�A����2C��"fd�=]LTs�xH73�L�ODm�D��sC������o��?�05��b`D��V�(A���a�_���DʪvHȼ�� �,���{�:q�oQ�uUq�+)\��}�v��[�Ϧo]���mֲ$�̱�]j�m��۳�����`�S&B0�Ǹ� ����$�s�͚}��m��`���@$p��N�ʤ(���S0�ҍ��6�(3�oK�ۙu��A#"6�I;����7�G\�4-�޶|?X�&���)�3G�<�ăs�͐Iw���zq`��
�3�]ĳ��e
�!��ݻ�4VyI"���޾�ӎ��Y�z���ް��㚉��J9�j�3�	;n�H����;�D�&HEL�Cb�>�t��RgnN�b�^�	 ���l�|�kκ�A�B��z���"|����4b��S��dI;ϣj{�IѸ���\�sħ}���B1����4�{<A��:i�qsK�b�7&�s�]ѻl�����6���|��^vl�7���[�2��f��g�'}����&н���V�}]��K�'1AU�E��y�|	��������	�77��;�l��P�?Y� ����h����LA	���)�S��dOIʊ�:�B����# 6{��I	�k`�˚10d���(����*ĥ�Ug}��|wy���7�I<c�,�ם �*�����V���s�y�~��ON}E�v=-θ����^�[�7�YS�,���;;��[U�:=U�n=�]����]�T�'�L�E8�|߉ �1�S-8���v�4m�[��9�A'���Ϣ6]�G��ؑMbh�YI"�\<c�`�5�p.6���)� ��?��[������`�(Ȉ�R~1Z�AO>�	��+ƍi�pf�9���6s�W1�&�����"n�,ᾬ��O�
�5�I'�uP�N_������h��nV2|-4,8��)�L�J�׸��1�@I�F+3b�U�uE_	�[}���_�q���޸�I%���S<��F�"�h$���d��}�2��A���k�S�����oI&ޏBx���xM:M;�$��}Y��ؽ��N��Vb����H�f:�	���S3���c'����1{Y�&v�2�-p�pU�!PK�U���b�Н�̲��y�>ݾ��q&�m�=&/r�i���b��{���~|����q���C"��ȇy�����q���*���U�vx.;Qم�x�������qs�=sh��q���"��3�k��ێ�.�h_sͲ��vͳ��&{t��K���ݷ<݆�u��c����������;��kx��s�[g�2��u=O��8y�n����[O�ۜq�	����`lMe�kn���n#F�u�z����U����X\�p9�����뮪���ۗ��#:���l�/$����CI���>���e�X�ĶZ���� "�mW��!��6�R��oy�IcP����T�QR"eA
z��z�{�$[�	���֒	�Q�+Ē�sdeUM�iݸ�6�1FD( Ę�,I���l�s~��,k��'z��� ��9ԂK��a�Me
d�*�<�ƃ��W;���IV�� ���a�U�m1k�z�F��$�]B��X$��" �l��^7��%e�v�f6M�N� �OM�6H]���B%�n,�'~�>I$�0� �6�o�4�m=�gG�)�Z=1�9�k��������1u�����x����~��|�k*xl#ת��K���d��gb�q�@��S*b���a �=�6C��6' �#�d\y���n��g���]~����y�i��r����������tw�����;����wO�`���9��%]�����\��ݙ��٨>����T�QR"eA��|����i��N��el����!�����W}���05��b`D��h�d���S{
�|H5�\�$���g�c��<)o=�K�B����L���ạ!L�eBT����2�I�����˙u�}o���������GFاU^���s��T�s�=X��.ر��\�dwG� �;��׮6��T��r�	��iT��|�!]�S$�yG\P5S5�b�L�}\� }��'�g��l������BH9����$T��A.���$�P��q�ښ���� ���0ؖ����B�z��Cg�
6�8���B��
��t�R��K��'�t-���S	��vU��I��Z���2-�3�����t�gY%vf� �к�i��D�@��LɃ`�s�YU&�i7	���ݴ�A���T	$9��ԅ�ܚǯ&���֒7�Q�A�*&K~5k�P$��shʾ���m�I�u���k%
��H��{�v���ϫ�y.cR]��6����q�u�lX�[/nNQ�$�B�&aO_!��T��H2a&��p �в�	$�=�٪0G6�&����������nB�%(�1%6믙WL�[ĉ����H�q^$.w��{aWj��|��ճFbP��* m��Ჭ���A�`o�z�e\눺�|A�uԂ	=�߉b�q� �Oi����~�}��| 𿮰ӹ͂I]����4�̲cx�a�)��&��9sHK��n�t�к�G���*{H�V%��[���R>痷�	,��6��^�wbln���Rp�lĥi�s8A�X��ـ�Dy$�L�F���2O���x>�%&�
''�[ ���[�.U�{��^d����k��e綨��mX���V�o&�v����A�x~R�e+�ASX�|�w� :o���'ī��̾��s����ΠF�]@�Hs�͂q4,C�(���J�>�� �KkT:{��t�k~$|��[ �mKL�e��:���Y*��i0�`�[����  �_�> !��)�s�$�=��]���v�(�J10�LL�u<B{����<��'����I!k�l�tuޔ���A�qCG���v�;R��!�J"`LC~�����E�]Ti��]J��WZ 
����+�k~$H��*���W��c���\�X4�b�d#���6��}�'���qr��i�M��bg.*�!=�c����C�/G��U%��s}����p����������2�6���)��e�^Ncƭv���s�v��Ρ���<��t�Ɍ���q���D��Fvcf�ޞ����]��%�g��	n��R�C�hݐ��u��9{���Py�z[�t9��ܽ;�9�m��Z�qǊ���h�[sk���s�)waö���[��l�ܜ�{:�		��{mh�c��pu�+��j��!�z���:���e�s�\uX�Չ6K۞���7	K�@��A21l ܵg�K�IO~���O�ǻL�H=s^5}��Z�5�`Fg6�*��`��050�D��l��ʢaّ�r7c����$�oy�I����(<�9�zLK��O�Z!ɐ�O�J���??1�RI Ӿ�j���fe���J��L	<��?/a���a��8��ޟ����EKF�IQ9�� �	�2(H���o���'L��~�]�CL�i��N��5�$�L>ΫήCUr�S�<J��l	��$��ΏfP�9�2Bۗw�ݮ�^�v-эqluy�wnxۢ��q�U�D���L���T�^n��%B!U��ݶA-�I ���E#�9������vGHȁP�=	DH�Q�O>a��Zp������X�0�#>,��Z����H���B���n�{��"�)��`�p�f�Q��KM��O(J�X��{�9L�A��(���o��nU¯T�2NLOM�M(W��J5���ԐH+o����/�+���Z�< �+ڀ|HW�͌q��1�?���/O�1:���*�kC�	�Nנ�
��H$\>��,l�[�{Sj��0H312"`�%����>*�u0v��I�a9ќ�ē�͂
���772���l���כ9D�qO"sD���=�lnַ7rp��pL����L�[h��8}ۘ� �m2I
�s`��_-Pj*��e�ԫ�F�u3�g8�1D	���y|�$Ƞx��ɋ�Q�!5y�@ �{���*�sd�U�C�V����uM?A���!DL�I����X�i�I�U�m�����ݭ���0û�����&o�
���B�x�C2�5
�ʍ
6(]�k�֯5PKy�L�����^����G,��fy��Nl
{�
��p�|���{;��ݢ.���P i��������1cANw��}��t�a��{_`���S�#�+S7�\H�_B�q��{6
<�R~�ןE���^�5HZhq�;=�F1q�j��A�`�Ui�[[Xv2ĭ�54�q���+^�Q��?K��i~�v]� ��#�v��ΒrNR'����{�	�x���80���}�x�
��j�b_:���la��؈=����6d���'{�*{{��������;�zy�-����9�xl�M^A9Ɲ�ˏ8$w���V��$�u����d3�E�����}]���~�q	կ-m��Բ3v�&�x��(8��^�y���)/�r^���[H=Mm�f����i�5w7DKj7!�6��ʷ�EҚ����3ہ�I���5l��G�'�2�^��?���{�'�OM��%)U���XFiO�������}p��[�J)���,�v�UgOk�������;��r���ɫ����$>N��;�n�j��J��Xu��U�t���J�d��<�]�!+}�賻�+��G�X��0��o%��D�$�s��M��w��y��|�������x�n��nN���{��L�x��Gp�?�ā����f{u�׿��<�-�1ҽ=�js8ݒN<v񻣐���zH��*���#-����� #ĐI$���"��EX�(��WL��[j��-\�(���*�A�U\�[J!Rܵ�S���\AZ�QB�""1kb�(*�D��-�f%mh�Š�Fe�L��*��0���UKEhѵD��̦��R�n\�Z�iJ�U
�T�m�F�Ѣ�V��Qm�Җ��E�ZT��\��m��efTKQ�cJ��X��Q���ĭj�2ܶ����m��mm��TeUZ5B�S.2�nZaZU� �6�7�`6�Gy�Z�-�eV�JT���S�y�����ەόa����yyMǷ q������lZ���7*��j6�U�[Z�&�e(��ɕ�<w/�&y�v6���.7�3��2����j�-Gѩe����F[���b-�����Rĩmj��)lLʘ��"��Kh�KD��F����Z˙��	m32٘W±h����6R�jf�R��w�ؤ�.�[$��6v�,�B�f%�f���a��;�թ:�%gf�@$�����ˮg,\#Y��f���d`'����1Z!��b'�$�� �W,����ti�X�([�� �HX�[$
��QQ`�GT:�����J��2N�fNք+<�B;O"meL^�ڂ�uqm���wV����H312"a$'8��l��U��`���P1@���a��|�$��_�f���)�R-�Z��w��[C1�u�x��� ��5�	�\��,�I�Wkn���wā�gx��1D0�<|�>$�֨\��
��N�X�a�X���??��CѴ2 8J���(�DGWU��0DE^/m�2	#�2���՚��ҩ̚������'o���spo��,yS�\�o�;)��k�����u��z�>���Ϋ��z=�yo��zsj�_�k�T��"-�H��S��P��B%�j���m�0캩ġ�2����B�1}��9�\�׭)����!��c�<`&۹u����ڮ8��ۊ,��]j�mۆ�c}��;�������n=�϶] O����ٞ�S��=�����?#����6�i�M����)����3r�NS���O�7mQ "���@>���EJݞ����z6Sl��l���ob ?_�  �Յ�a�y'Uw2I�X��z1}�L�C��$`I��cJL͗�ONkpz�r���5B��G^s`����o��h��f��I�c&h�D��3Ϙgĕ���Q���3m;������D�#3u�V����uX�5w
�Vȹ�6��<Al"T�׭P�˜�����ˮ&ͫ�в?j��>��c-�7�a7^�F���e�A��gP߇,�����t�:Ρ�p�>_Ug�6Sz��K��� 
�N�2��X��8vݓ�-Ք@�(y����q=N��p�� pp�K�F�Vy)h�|^}w-[v,�4�Z�Ϩ�S�n��
�����[gtq�z���ǜq��r�^5�gS��;���TR0��B31L�t��Z�Z�6��L��6�F��H���9�>��t�On���d��玗n��>9籬���4��#	�y�+�xw[q�;vO<�JSP�&3t��{��1(L���Y�Āco��J��C�h=m؛���0�:x���'t D;�a�6lC ��
!#@<}��V�gV*\���	";;�����'ǸY���ĻFb��t2D�L��I	����dJ��LI��F����:UF3�#w��I*��k%�*cm2�����{�Q�r[@���dV=��>";�ͫ�|�a@�F�v0��3�RD���"�n�u�	E�]'�TH�yecw����v���z_'0�#v���Mb!��&�,3�����j(�7f�#�C:tb����_V������۳�"H�����d�W�6� �H��ܩى7���Sy=5^�.y͂F_�y�f%	�;���	Բt�8kIZn�����=u�*b�UX�t��ر�1�I�&�c�Tv��7;�@p2=���ݓ��α����鞽���	";��{������]u`�ٱL�3(DAF��z�$��4O��y�]TsxI*�y�H'�wC�G/a�� 6��I�&�~�E�T^~&�gl�аs�:�>>W��x_wS�ӯNqX]�fOҽ�lbM�Z߃�#+ȂA����d�Sur	g��|O���E��i��Yp�Zj �#`J�][]uE֟Gf7�1��xn�v;!v�҃��ZD��+���Ib&L	K�st8Vl:D�L^�6c1ol-Rh��Ym�A[�h�d�d!D�]A��k,�UΈ�}}X	k�W��^�6H9=}�7U(�����&/��1(L�m�M O�&6���-o��O�]�װ���T����ez�ݧ{K���9�q���13�\БW���}NÝ���
{�,߸4jv"D]��VY�S|	�%g9�@�����nц�q$ܛY ���j�Ӿ {b���>����*���a�sZ`��:�#���f`)������6I*�:�X��˰O���A�9�>U}͏�#:R0��]tƝ�J#��0>3�Z��RæP��d��Ol�R&in�ٸӛ�__?{Ű�l0�i��"�@�)o�ɘ��7�Ӱ��O���>����9�$��0`)��;|߉���F�IN�C53���D�v��E�6I�퉉K�?)��>��<��8R���F�sϛ$���}�"r�(�
����z8�;���ME�6O��)1~EA3�����j���}M�gf�~ Tv�`�A[�FL]r��})�+Y��oXȞ�rP�f��l�8�Y<Z�f-�V	��d����[B8ą.^��s�uB�L�&"�+�q����sz��q�(���a���/��`=�hxۙJ�Gf#��=͒J��l�o9��t?j~�̽�����r/8�}m��b�=no-�Ȼ��q��<X�㭍���K_�����m3b
Bw���~$��I[�Ex`���UR�@��ȫ���!Vv�~�Ka��h��-h{���x>o�q_�p�@*�6�$��揠����x�o:��gx��&0�e�`ڜ'Ę�n��OgtN��aV�>'�w9�F��a�	&F����:�7.J�;!�V:t�$������D^�7d�ۊՠ�e�[��h0�fe	��orh�6��*�n"ݬ��r��`�V�L_w6u�<VЋ2yX���-�����y��w%%��m�/QP��u�`��Mԣc$��۫ ֱ]�j��}�Y���c�=5L���uo����~~m�f��a|�Y��hv��Ȇu��N���p;k�aa��q���ҧ	t#Ƶ�g���O&�
N�3��u���F��W�ΞZp<qj'���y�������Ƚ�:�tkzL��S�6�7��r��kChx�]>�x�Mv{n^U+���8��}}g���Yz��=�P����^��7��.�ޑnɶ6n�]��U�(�<�������˻2�R5��q�5v���K �b�x�nG,��l[�/����l�u������0� �8�@$E�s`�B9GJ19B�j.:]g�"�����G!X@̡1!-���c�w�=:�U.j���Y�p$�b����+3��kr֜��'\uLJ3)B���1G^@�LW_S$�َ��|l�Nh�H9�$�	���2Lg�""f��+k-�KaH.L�C'� O� ���a�����ɭpv����#O��&0�1`��h����HU���y]�+U�\�n�	����$������l��I.~�bL��`�X��v^v�%���.&�ڤ�:x�b�z5[�f��d���H@��&s����O��{�� �W�ټ�R����QB�5�/\O� ��u0O��K�JfT��(Ӭ�l��4���7+~��Kzf�l����E�w���^���]�Ԩ�2��%M;�|	����D�������ӗ57�/v��W��1�H���A!s�l���'�s�:a!�#��!*H��������`�V<�~$|_t���9a�	����y�1�S�̈�S2�(w]r��}lxݶ	 +y͐A��Ev���Ѿ`�z��Q��DL�Ø��0��Q'���c(ɬT	湰H$�5��1��F�z9���9��T�#����	�R�z-�v�.���WZ�ݚ��Wn��N�X�b���7�峸a@�DFS�0J׻L�|O��}\.{FA��]!��6I![�a��B̡2�5�A=�A컘�Q�Fc3C$���I �I���VutL۽݅�#M����g�'�g�?]O�0 δ�FA�QJ�����0���ΤZwC�!�w{s�&�uN���'/Kw50�I�ݝ"m4^T\FE�^���p64�%<K�KuAZ�GB�� ��=FɈTT*��T�k�L���9KTV�uٵ H��Ì��:�;�]���Y�SS*�TI3q�&�B���m�WWD�u��${�$@0���b3B;6ȥ�����EJF|}1�0qtoM�)��s�hҪPt�N�7S��W�x���?~`;pЄ0�T��~$�s���{��knf��w��7�� 멁��cL׌�>~d�j�9Jk�V�S�> �6�H �}�߉3�U����v����B̡2�5�H$ƾ���"�����������v�H �C�� ��m����O��ؿ"�f~�Rm��3P'Ăco����9ؾ=�N)7�i���W�bftĘ���y�����!|����&�^)�����U�M��zo{�4�no�I��P�Ѭ�p���O�mD��F�Y&T�0!4���S��:��<U���%�{`�5�$�L[�l�B��l�DL�,�sX�(Xt�����9G��ۙ'��k!���a���Q�[�����g���-cd���ڿ`����]�O�at%}ЬQ0�=>�1n��FQ��(�HB3�N[����q�M����O�9�0ʫަO�A.";6��o�
�0�I��Q3
G����2	*������U�G���o�$C����*�y��������3(L�u�j�SBj�)�e*���I�*���I=�\�gw~[�pi��`^�&&[G"L")��7�A'����x̬���2iE�~������$�	'� �$���IO��IJ��$�p$�	'�@�$��H@��B���$�	'���$���$ I?���$�	!I@�$��IO��$ I?���$�XB���IO��$ I?���$�B���(+$�k<Q��hG0
 ��d��Dg|v�          
P @        �     P     �� s�Q��
�*T$��J���l��R�T��}�A"vĠUi�M�(����R**RP���B��"��U=�                                        @        �B�1���]yt{��ty�<�N��  ��zà����1����� ��� .�W!���hw�"��*�   ���h�70��<  z2;��CW�Q͔�)����v�;�p���cN]]����6P�<�P�Q+�]|           � ހ�6���5š�59Ru�3��p 8 �sw|n
�� �¸�����ɧCi\ � �PYat�B�ޕ*�2QL�p   @x�):�}�q(�` 3B�@s`�YB�^`4�eJ�{��7����Bz� �(��(0j��I�o3J��;���@�[Llf�H\  �        z��8����=�:�_YJ0j���x���� �Cu�9.�����о�^`�/\  � 緣�PAAJ�� C��g��� w@sw���y����y��T9, t@ �����1�gE��ĩ � �        ���|��^�{����3�j8� `F�����e<Z	Q�C��x �{�y��6�H�k!C�  >����>T�`�x  vg]���� r���ۀ� �7��/3��y��{;��Z�j���[�  >         |u�9j�N!��O!����x  	k��+š�����5�����@�����+5ź��P�f�K�   ���>�[0��:m�x �	{��=���.�uU媡=�.���rU�oV���-J�)9�R�j�� �CAIJ� )�4�)T� � �i��T�� '�UA���i�0A�~�L*� i@����<ԟ�����'�����xh��U�0!�g<*RW��I	L�;���$$ I5		�$$ I?�HH@�Đ��$d� �����>�������y���]��3�q�y�9�f��тM���6eUEr�4/<!�e�@����+r�A]*j; ���%�Y�7�Ŷ�'��f�.zE%RV~c7���^#�Q��L"��s��R��8ݜ/eѶ��2'.#�`��G����|p�_N��'HS���|���ñ���gN�ٓel����jN��F{5�J��]+o34��y�ʲv��j���+t�T����@*���Rg�s/U�K;`�_�������v��-;=o�%�lH�<dm�q��Т�ls��E�ASJ��ݴ��vB�?1^@� �G/5����=��&��֬��oF�[��Щ���oIJADj�hl���(��y��v����ɻ_E��S�c�g��󕛁��d�̌ryM�^)�#��-:!t�cV�F(^ev��a��ܜ�i�!�\4�Uo}�m�M+�{�6n��W�i�6:h�)k2�?3����&�&�M���d�Z�-�u5����%�'�wh@��mM[.���+G�X-�;�[�ןA{�Lch�;�<L�;Z�8[m��e��0oۛ�ec�pj���ƾ7Lޘ���lTF9p��MɪO��`�9��Cb[��4s����b�
p�T�H�k6�5Rv[�u6X��z4��;�"���<�Ѻ�L;�7����1=����m�VrU�B=��wF�-���rE�=T�[��`�"o�n�XI�q0׳��1a���ޙ/u�̜Jq���I��V��W����*2��JNӰ�+���Crv��D�U�8���9Y����f����<���q�3�A�:� ";��C�����~��;�����W�Gg"7�ݨWӬ�Y��9-�t0k�rQ�ݤ׹	&����Ц��޻B6���<����i�k�.q`o	�7xm�V�i(-Մ��Yb���wU��˜r٨M�<q��)�4��ޔ\�w�/����穝��۹�6ȇrH=ɴ;z���@L/ 3���\}zB����m\YJ��ᴛ��Ƙ/-���7��_=����tWvn۪j����}�~x��T�,�$TpS�^T}oðw<C�db��VQ#(�'r�����RÝ���I?%�^v��Ct�Q\¸���xiY�f�¶��6��}h���N�t��z%�	{pH��93��7��Z�s�gn���Ҳ��0���A������s�C[�i*b�L̵܋���X�na�H׷+�I�ǳ"Yya��@�wPb��%��������D�v g�q��OM�j��"��,e�w������9��'M#�㢫���H���r[��Ϸs�p}�gI;�@�(.��ĺ�a�;�t�lY�����*#/��m���m�Q���wc�g �{:3�n��G�n�zћ�Y�%Z��6.n��/��:jWe�Q�����ˈ���K'V�7f�p��rvcl]����ۃy���eC�Ѹ@'zms���|T��z��%�0�w{��kA4Ѥ!섰s���'"�Ȏ�5�=�tn�[8os�}��tY)��+�(����ù�ŝ#:�V�Xq�w���3n�;!4NځX_n�ru�;5
#9�;��tӀҭ��(��bރ�vt;'1�Q�A%�w.H5fӬ��Z;r^<��b�3ook1�3����h]��E�,-e([C�;��/+����r�ъ�D6��H�nl.�!op�Ѩ�v�xNNO�;���4T�#X��mE��!���m<�snq��r0a���x]y��Xr��;�*�c/�V[�N��=��
A�!p�;{3��ŧFŭ��b�u(&]K�F-�l��i"� ��QI�W|N��g<��C9�iѺN��{t���{�[r�[F���搧��Tb}�
��Sf�2}��[�piם�S;�O�+�vΠF��}��mR��Ǘ x�Lަ+VQK��p=whwq�fL��y`��-wp���W���`��Y;N{;���un�X6�����`L��{������3��gv򷜩
��8�̓��Lq�JN%�7[LNY�d֤;������D:~� �"�}Q��יՠhغ^��-gR���2��{�~�S�40P"�V<��.F�������L�j �G/�nL�K�K�;^Sv��{3W�\�i����J���wBޢ(�N x&�$AM^��k�M���ٵ���D� N=���:�h�s���P��uG9m�q
��;kWt5LSK鼄l�(N�ْ��mv��.Uf�g��[��a�92b��Y�ak��
"47o6�1������ʪ�za�������v#a܆�%�T@����1��q����4�§%'p�u�f�����"ܭ�%°��2hO�62u�/t������C�n�sNwb�l�c��%�ݨ�jr���'q�Fi<�����Gx�y+��x�Q�L�Iou�T<���wcp�Nj�dp\�j͔�a��M|e��wD��� PT�Be2뛩��W��k!@~lVN��(�M��-6]r7�E�pl�5��9¤�#��u+&��.m����p��ϩc9ְ��g�����]d���ө��@hʄ��-�¸j��̹��I
�7���N��tU؅�$�s�ô6����.8`a3Y]!q�X5���\��ܨ|�9ڃq�q�6�v���0��!��FQ�V�Y�ᶰ;�)q���6ڈ�<�s�Ğգ7*3V�5�J�l��C1�w�w�雅�:I'aT��5�&�.1�4utiFNnK�6����j\@���2q�q^�N�� �KDH۫�$v����R����kX9�x�䮫Gk�1�������q�Q�o�/�p<g�����7s�����������[�Q�L����k��Eϱc����!��s�s���i��-l�tnH��e� �]��h9V�|���
�v��;!ο"��v2���)��Ġa�p��t�������'S�l��KL�y��i����D��qݚج\�Z��l����ϪŻ{�!����=�����O)s������vj��r��㓵I7
0o�, gU�e���%��hld���l����4�������[Op�W>�5I����Ă��5lޥ�੘6�hQ���U�Eg��Qϙ���V=���=�v�;��.nZr��f�Q��z��l��-gm��ٻ0rr!-qi�k�r8{n|w=����ӛ��y���a1x��RMt[�F��N�Lٚ�K�s���h�v�Q����:/f��v�C�jͯ�D��1����w�c��)��z�lM�{.�xݧO��+���x*өN��gm�q�p�v�]���4��5JLh93u2z:֭:6dU����n�6풃�5��1y��4;2��{˚�Ã�Bӡ @<�%�v�Թ�stȦ��M��3p�.zw����_tz#�F�!���&f��\n�˒��a�b��k�����S�.l�;�t��,�k�R�Axi�^MޜvR;֞�2�Α�'�r�����7 �h�.��6�obC'E>��7َ������x��o"�-�\jP��v��߯mn�Тo-�{�`O{^*���v�W���̗g�6(V'�eދ:i�;�1�Fe�Nڭ#P�7��`·6[1��b��;P;7wp�pd�qfٕ�>w��S)i��F�r�&���@8���1kcbV����Ѐsgv�;3[�_W/&^�= ��콩���o����v�[�Pؤ���B�n�˜��G��&2^�3S�1�n=��}A�j��cWgb�դ�jYp����q���à����1`���:ީ�N}�]T�	��xnm7q��vu�h�u��ˏ�8��d�`r;��/,ɱ��8f�>�ssnǥ$4Y��@��ДZ�ooM@a�lI{�߮���ѫ�`�u���ܲ�c��	�Os��յS�U�[u��t�Sph��ZU4���نҰ�����n]�2�|& �L^ɷ�p��ɚN��u�-B�ݏ0C{C����BKV]FRܐ�8 O�����l�ӹ=��U(6�F�kx-�8a�iv%��u��se:�q曦���٢��2��Û&�_Z�ވ��ݕme�Z���3��U�i�X�gkNս�@�>�l��,w�Iy��=Ü��2i]5,��^Ɲ�z��n�T];I���H��f���v�D$��W�)�;�9��h�f3$�T����j��[Y�@F�y�4;�H;~��)��'��t��^�2��;`��U�8և\95��r����;���rNO�Z�:�61;��\l���a�i
5��F���1�ǼY�9��fL���{kj�txr�V/c��`���r�]Ѓ����q��}#u]��a�U��GŢ�S9���o�iWԺł�h�A{����~t�{6x�Aty����u��tD�P���G�f�n��RAZՇ�С���msy߆p7����Y���jZ-�����؅���ݐ�Ϋ�cF�w�S�3V)7i'7��$�n�Z��%�=�dh���(�p{�Lc���P]r��1k�:S����3��)�m���o���}�Nqq��B�8
Ȧw>p��d��z�܏DI��u]x�	^��&�7��fK-��\���X�:r���3�)��'Z=f�gSb@�&��^�؃A ���y����worG�y�a���Z���q�9oIrc͈v��Ȫ�������ِ��+���v��5:��f��\ ��Q�^�@�s�wy	c�r��LsA�Q�7�,�\�;����-A8�fܺ7�=�n��WJf�Z�2�'h�]�\�A��4m�N�8w�<B�F^D�`�8I��M��;�-eXْ�OjsD~Ԥ�0��{��s�L�i{.J��;��h���&˫����r�<�1+�'�s7�M�ӌwvς]R��wv3��w���e:G;���w^:��;�]�E��'���u E��sU�v��74^��᳍��%��(3��A�Q&X}���XqN�a��A��y���V]��ӥ�l�U�m��uk�ovHt�_X�����Y��~��/k7X�I�q��ǆ��o]
s3"��6��.�^!��C�Vpd���{^>�ӛz69�l[Ŭh6[���`���p;����p��)���;�r�^v�e#��ח;�i�.	Ƌ٥]ʭr�y��Y^N�����e��,��ۺ+,�DR}f�E�|�_�n�)x�19gR�c��KF��:AV�F��s31�}��5T�sN������.$p�m� u��]ܡ�;�s�@����њ^Į��1�r�թs��D��6�ObR�ʷ ռ��b�hZz�qb�n�x���g#f�x�;^�r 
�Kf��7�K֜X�5p}F�x�A��b 5i�_��0a�jrX�m�,t����$�Fv�&�N��m�݃:-�!ι���{�^PmYmKF�����\���vV���� ii��ga���}.�7���S�U	cn4e����W��	��m��[��'���m�ii��N�{�e�W�q@F!�F̺ٛX�NF�"۠�ĬL�k�C6txaN���ڟN�u�1g7��f��O�	ӋK��dзN����� P�	v�6�onv�Z��x�6��X��R��J���<\D��hZ5�VK���gH=�"��������6��;\�x޶<��wV��5�n�GN��ͧ91'C��;�e[om��i[�q��`W��-�vM;l���y�l���ݻ�ӼҸ��`.}ٲ�����W<!�,����\�yx,T���V����
4�L��R4J�E=[>�)�B�^R��b�d���c�]ˣ��d��Ã���7�+pq��bd�� <h�i���H�U�-w���E+x/K�kgڲV�V�k�L)鼦#�b�7�B�gri��qʀ�pr�4Ӹ �nӠ���:9�}�5�5[C��h�y;x�T7��\�.�SI=��j9a9ۯVͭ[e� Rw	����H;�0Deۣ�Ȏ7�:+��e�']�n�6���QB��;�� �&l�U����`X����h����;T���02_�C����[��ݡ	��Wkp92��)XV�tS�k�����l��ɋp��0��{;#H��t�\�r94S���5��.nu;{�n�7F!ܰ�{9���~H���/:������� ��UՋt�5>3lE�:q���Y��: �[��i�eVb%98n��w$��t�1 �7&�2�Sz�o#��F���K��*'�d{�&�0���$`��uK+�d̯ze�#�X��QZ��ӆ-�?�40'@�C�t>�v	V�#�pLۥQs�|[A���PNs ��֍FWK;[���-:�)un.0<�Aۥ��wt��EB"��XӚ�F�Ÿc��0�Ű�mn��/n�U�gs�o��LѓV�w�?\}���'Nj�F5�xd8����#�s��09���9�ԅٸ7��X\#vt	�ۗ5l�{�5�8�un5����2���@��$$�	�I%B�VJ²@�Id�@��$RB@X�@��$	HI$RBd,	� 
I"�$Y$HJ�I
�"�
� T$RAH��B,��HVH���Y@+ 	Y!*@�BH�B@Y���
�a$a$R@�P�I Y$	 )d$�Y$ ,! ,�X	"� T�	Y @�!`H
 BT�@XHE$�"�@
�*� "�"�$*�T	$��IP��H! � XB�*@(�,�!(E ���!!
�@RXY �Aa A`+ �$�I!!� =��z��~�/⊀濟ȣ/�&�eZ(��݌>v��Cr��3<�6��+�%U+�G�����ɚ�%K���\�f��T�udg�Mc��< ^ f�'?y>x��O���c�P��@�;��}���|[ɥ�u*�D5�S��\�i�no�ԣWM4��Q�N�'�<�k�۞�]�Nn�#M�ܙ1��Hf��Qt�����l;�6�]�W�1�����$�y�6#ro_�~�Q�e҃�ñ��	�>�&�[�|E�:��&I��޵b'z��e��S�/κ�_2�B�Ѽ�g;�+*��2uwb�WhY8U�Ե�̵�ڳI��4�����^�ͽ�eY]�ܽ�N6N��[$�w��5���j��|.-GR��=�ySXq%���K��N����;��Yj�a�T��v�L*�ܝ���E���^Ⱥ��h�km�@ў]�u{�J��;Ab�LYDv`���.+���a�koS8���.v�nH��L+V{���2lnT���k��7���QOa����0�C����;�=������=wmQ]
��5t�Y碱�ׁ�p�8��N��Liӆ�Ѳ`����Niaf��2M]֨	�"�6[�=\ ^���4�*�B��%gZL�K�<X�8<��9)�XD�e��/��l��B���&,��NҷVi���]uo�_+��έ�:b#C�&��N����+���5"�H��9vk�Y#�3{Eo��9a��;xm��\;�}��t���b�K�gz>���7p �	+�͏7w{�,FaG4��۹\�H�c��F��xz,�߾Bf�I�K���L��E/�SUB���x�2��,�t�xޭ��9��&�y��0N�#���Pm&�}�&q�ٻ��΍��"�qk����ޒ�;	\4�7[a��j��YRm	���U�w~Jǧ��! ��˪#ږ��nn����KW3�lV臸�L�f�{hn�:%}5�1	�\}�=�^]Mf���^.�*��ou0���v��p� ��{;�xZv��H����g��A�Y�맸?j�Q�'N��\��/������j���$�2��(T�ᄮj��K�y��-Cfλyh�<�L5�r��C��{}O+�L��w3}b~�^{����<�HN=����H��R�A�j�v2T��2�,���'|)X��@qr�-p=~��= ��ζ..\�ͧV���Hve���;��5�(��tc�X�܂�C�z�ڙڅ����0��ݔ�M]O�n7֯
����Q85�Ĳ:6�5M�Df��^�T�з���/O��<�ÅA���}��Y=��f��x o�*����U̒ͅz�iⳛ��ӛ�P֍Y��u'H�X�"ҥ�rfl����2=:3����ut��t?�nuA���3��K�fd_-vl���1e��׶��9j��b*���B!�7�}	�j�'�̀V�X���|��y�C�S��cK��˂+���̻�q�oaV �z�Wc�=�WBn� ���ыR	P�iy���2�m�G]�C�z�2�`�]~O�UM�IĐJ�u��: �WO���A�×�*�܈�����pI�T�_o{heA�L�*�Q����)C4�6r��̦*�,��_U�rڔ�Q����n�Fޟo15�ʆ�-��d��*�EU8��̈́�F�̹0���׾��gQݷ����v����95xt��|��d/v.��6�G)�ni�C�X��sʟ��;_j@��0p�0{��ᦀ],��g��{�:xъ	w}��ɣ�z�G��闭pG�;��B2�mr5h#z5l���%���>F�x��B��u鷙VB^���-����:��{&OH7s��׷Ǳ�����&�|���S�>*8s�Y���2�j�<��+F��Цq��X#b�mQ~� �bI�n!��0lV��aL�Oz�qp՗7�=o"Er��B�b�(v{�{�p�~[9���/+}�K.�Q�s7�u�p�鹘�3X`i`��3��ad�ۢ��{Ś��JE]��/D8�mO:�弨���1���*Y{O�l7}�=}g�x�,�6*�YZ8F�	#:}aA{�R���mN�۫�Kʡ��H{
����L,W���V��[OG����
Vvo�j���\�'yj�n�^���<h�����]Y�}(mÏ�3�:�27U�DH����*�����x�#�L�~��ʎ@����th�;aȡ�SQ�/+�I��C3��W~v�<gwo��_N�xs��l�U��a�PN�8"*�=41�ٽ�����(x��g��A>�e�n�z����]k-�t{n��H쵇�e>ʘ�]�8�����\lҲ�w�/�qTt�^�o>���7ԝ��:_��x6��D���UE.x��	�0����b�;�:z�&{���у��D$��r�T�t�TW��"�c{hlx9IvP��Vئ���hFKVqPF�x�i�%��:0vvk~����NE%B�j�U+ב3 ���G^��=r�{�/gz��*��f/������,n9O��+��ƪY�W�Έ����@�zM�8X��D�˙�4wx���:�-C�쌳��d��3�D�֜Y�y�+��$��uR�Ã+���:=�VI4�&���Exy{�H��t���3n.�ƥ�V�3�ٔ,3�ܕڄ�S�p����{υ�8I�
٫(�@x�Y:��T�/qR,�����nxz���Ŕ�ղL�x@��kT؈}p=��[��$��c�o�wƴ��<�ۥo��U!7o��A�A�%�Z�R�MB���U��f{;���ە�g�K�2��q��ug>�(�l�4S�>mU���7b�6c��0'��n���ߋˇ�7�-�&� c
�Gj���ӜmbP*��ß+[��8]Ŗ}I2�߅��`0�=���;8�-���:�G�)q���hl(=��.�ƽ��w)�$��0�ɖo3�m�c�S��|�b����Ӷ�l(xOr�2.�k��<�Hĩ�q0^��:Eb��ug�,y�nN4.�Tk5�9ԋ4Ѯ���z�gt�n	�,��`��sOs��m�#��u�3B��Ig}�f�[m�~�]Z+x-�u@{|{�l� Z�z��Ų�Cw�}�<q���� 
J�j��ο1Fj=�(��$��I�A2@ �ٴ�קiy��d�lv؆��w�>��������1�\D���T�]�­G�4��Ԫ*�
�Qv�u�"=˪��/{p�8�����|Iy��&$[὞�;Oq��J�&-����o0�&eO:�7�vU�I��*�f� ��W�	}��z'�k�������;|��y7��\��X!�DSd�1i=�Yt)�ĽWZz�.]3�dm�L�;�Z�ע��;f3��ʭ��;��mH��uA���+=[Z-��}��:�9�E����	b~8+N�]܅��Gn�٭�"X3�y�gW]�*�%.��v�,I�[xb�u�)������ܪǌNf��1�fI3`��-饄L�-��b�����kgz�n�*.�����F��8Qn��]R��R�Q9t7!,]K4��Ԓ[��s�C�i��-�2
Ȗ��*SfNշU{X�
�{h�4q��/$*�!�%�y
Q�d��ֳ��q�O���Y�X\�`>槵��r����eʸY�����V���y.S(W_�o��Q��u}ʼWn�$�wM}��z���i���F��yvo�;�kvH�X9.�]�3�9=��dm����s��&HZ�B�Tg�u���#��+�Ug �G��Q��w���`���=�3j�b��P�����N��Z��٥��eeMM���H��E^ܙ^I5�9a$_I��_r�����T2"�ክ�	H3[�g�Ov�7v=�&Y=Q���Gk��Kٯ�X���[�u2��̈́lnx�Ȭ�Z�ǝ}�/����m'�*E����3R�^��Uir����q�E�5���n��:�������DX��Z�g��F�eCs�K���`�6���I�a�ݘ��{;e ����Sy]��W�uQ�K��r�=��r�=�Lń�U��,pN
F��ݽ�}<�Y=}:-�cEvv]�����[1������1�3��K_�ċث��3��ћPrY�ѠO.��>���S3_l�-q"��%q�z�
l@����(c�J���p�5�C��s:���uC�p��w�O�1E����P�4��]�v)x_r4�%��h��w��"��ԉ9��-Q��!B�x7V��ð`[���e�/u���j��E���Q�����xy����bSU�����q�nDw�X�î5��oq{VI�R�e-Ǻ�x��������� �绺}�rc��O�[ڭ���݁N��(�+��+\W=�n�'I�����[ �h��nxg��ǈ�:�'� g�p����{�����dav�#��S����jЂn3�+���I�j^�U84q��C�]�ף|*����9I⏽��g{�Z���築<ۇ;*���u�3��J��ݑ/o�r��3�G��ɛ��g4lD�o�U�bjJIN�6�ǳ}�K�e֤����n%�;�AɈ*PS�y�QU��4*md�ՙZ�j� �/�t:�+�����p�Mkǋ" ̖um^]��]��Ό�#UcUAi��>��{����!W6sޡUTWd`�<�3��tȖ��K{��`�.��V.쾁�)݇�`���b���F���=��<I�5�R�K#F,�<���L����v���XĐ��,��G&-�(Q�2�*�\�a�#�X}�Y�U��3�����x��	>����zw�˩FX����gG&�q�]�	Ѓ�Fɳ�a��Ή�̥j֭��Ӹ ��x�A]���XJEY5Uj.�'C��I��M��'�G��< ��L���qd|��3yם2TU �6�Ml�u��ޥw�؎0)���;�f8.��$wF�\���`T{2���]AvW�����XU�_4�����Q��wl�O{� k��_�»��CO�������k�wE���w���X�6��1����J��sY"8q�h䝚<�/�8���mq������G;Y���^���g��)�����sE��;�����3�}�6���U��狧�����m����G}U�Yc�'��2#����G���4�N�Egv�f���ֶ�����{7�W��`~���/n (V9G0V�˨�_dw[bưg�U"ήİQNm;V��t<�D�!��>k�;L�����u��v=m��!����R�Y���^2u��h�B��m��Q�V��9᷐֘9u���Q����/R�-���Y*m�0���Fv�=JÎ8.�y���0cΚ9U��E&�����hFZ�\γ�=<������(4h�L���0�m�Irtn���.=�CC���v:1�Y���$uUx����t��ς7O�����vL���T�Q�1l�^�5�N��0��"Ag-7�����^7:baeo5d*Z+A�.��ý�%P�[F��9����嚎���nk��{�J<��\H+6c���G�����妻,u	��� �z���!�0T�+�E3I�&�������l��E�wTK���_w!�7c܆���D/ c7�ҧc^��N�8%/=��45�ޜ��CMތ�J�Z����w����M�A����^�4��i�K�u���/D:�jo����l^����D39���!���=�ը���r���璙���YQ�9iD�q�}�?#Iٱ�ğL��P�������>��lX�I�`��f�u��FL=�	Z.jk7*�'�yxׯ����<��N,=%7!�F]Ƞ���)�[��M������:��n�͂��_.]�vS�N�<�v�9}0�k#�Q
p�Y0��Eݳdͦ��v,u�`5�ٮKY\�:�cTe����F>T�	���UX��ӷ�p+Z&I�YMDAuٕL�s��UG����bo�s$��Gg�{�բ�o��\<6��7o�1�j����E~g#�W�����/E����G�wl���⡴[����QfsO)���=���`g,hvP\ndΖ<���K��^��%�xy\�*�ǝ3�̏�O��i{բvJ����s����=�b�MYXz��o��t:s�\�4Qz�»~l1[y�y��T�w��R�${&ԧCVb���Asrƶ���}���aF���nY �,��~.,���gp'�ּ�V!Q���wnU���kw�x�M��ո6��MP�<�ei�"�;��!P��>ś �AF�]�A�:Md�ض-oH�fa|�Ԙ�&��Xέ�Aзq#!ܒ�s.r�Žo��/\���6��Q�#i�=<m-Q�'���9ʳ��1a������6�^u-a�`����>����S�ǔ�.����V4��Ε�b����jn�./�X4:�$vn�T�R��|�bGr�$��y��+��R=���%u����C�g3�u�㲲��
+���<fw	m$^w]:,N~�69�5��L͈��Cnn����`�{R�����V�ur�Ϊ;Oe�=�Џ��R��<��F�=�/=0@�OG��U� �A�o����S��{��pٛ}H��~7�7݋��,x�����8�0<Idq:��r�XD������(,Td�bY:�=W��Vy��^X���D��&��FfQ�w��/dt3f���Gٯw�W�xb��^Q�{cUUD,�qc�Oa�Բ�/8��TYr1H��ۑw]�nw*��oy�⠸������r�;k�}9��߿�$$ I?I4�[���G83���v`��qS�K�j.��[���u�
����=�m��.ݍ��u!��Nlg�"N����sh���,v�8��M�z:zz%z���se�ʻ,�Cx1����]g�qv�۬XY�8Ϭ��ǨZG��g� /Aɹuw)������ۆ�Ӎ�<��=��s�a��ti-�m�9Gm��xV���ݢ��Rl{^�gr�e��]�sړ��L���8x�ln��,�m����l�3��vtx.z�@�"bўԜ���ۮ:A��Wd]���km�l��wn��viNnI����ƹ{<z����OPb_l��t�e��7��َdۍ��c���۷)z�����=�\0`1nxv��h��]��ל�s�덷;c��^�&:� �:nܷAݝs���#^�{=�*.c�B;����c�=�m�p���p���pۮ´��wm�Վ�r]��ǎs��^S�9�o3������`�5ѓ��ǲ����xY��l�V1�n2��.�;�$��d.U�u�ӗ��+4��BN�wXev������onf��{�;F���r�]\�0k��ݑ�m�v��e�h��v����h̾Mb��.r�sڔ�ڷ&ta��G;p������>.B{k�hW[��c�,/$�u���X�Ht���l2��8`��([Iu�9לn�sȇ\��ٗ�����b�yy�sWgj"������T���!��׃T�Nkk��s�^w	�n-�ہ�n^읰Y�f��lݷۣ��۸���������5p���ݷ1�uf�y�g����[oV���ڦ/GC��<-p��
v�/�(G�ct���W��'�{5��[��m��7�Իl��^m���k�"�}���S5��8��<2��mu=����p��{N�C�nݴ^�gu�\�W'�&t����X�<Ǆ����4��fy7n����-��Y�Ms����
TU�km���nW�^U�F�j瓏)��۷���uΉz��'��N[��:^�½�3â��:��Ϸ;�:�J	'����n�n6����0��5�س<=)s۔;<�\�H��ۍ�X;'aCu��ɸ�$���ノ�\l��4��D�k���2��t�*�5͚�vcp��x�mO)��/3����|�*�m��=���vi�sp�k+nB:���y|�uk����n�rd�`^��::����:{�^a��s�8�,�M��9�c�9l�8��	�s�k�Åqb;�;]�s�Ki��4s�O<{<��v���1���ֵ��&�68:C��G�����Iك�ۖ��]��g��j��n�N6<:��ޗq�G�I�kmnm�R�B�5����x;.�w'U�zإ��5��L[�|]�l���`vsmm�@U2��obs���WS`��[=��3��D`^��O\���{ps��[.Ǭ�ר�ζ��=ήٛ�l���O;��:5����b���]�F�M۞��I��P�\�ѥ�����N9���N�xz�MX�w�+��C�W\N}�\�� w�9���ނ��D'�Fɮ�C�.�6��G��s��� ��+���F
�ce1��n^
��^7��lg�3G1�H�5�����u۲�<K��v��COobMۨp��Ʒ��t�%�S�W6h6��Ƿ�Yَٔ3�m�v��"���Oc��<��d���	n���۫]��nK���]�v�Mu��^���b��˶������<�6.�9���P=ӥ4Wc��\���C;���ҧ'��s�*ټV��]c���i'��#�^�v�"�n4`�ucv�}c�On<�I7n�>���Le�/Xx�0��*��i{z�=<ʓ�]�]���p��뭍���Ĉ-���v�n�wy6���;"�r�j)�h�q�m�:���ӻ[�a�f3�=�۱	�h97m�X���Q:ǃ�p�aۂݣ��h�B^�^��nQ�ל6�lg�L�W<cn���60�8 ����>��rg�����v�q;t�oU�������,�c۬	�(u�;`�r��K3�&���:qp�h0�M��Nt
n1Z�v�\K�НE��a�}�䝙ې�p�kk/h��x��{l80���mɰBb�m�'Q�c׶%��1˼j�������Xkp�g\b��5��$����sX���!�T어D�&�!�m��;[8ȯ��<��"�;Wmv;9�D�[nC[`�/G(q��y7O�Z�Dp�w\q�е��>��F�a�t�3s�9�a���]��6��k^�U�ë��.�d��A��^�����6�]�n���֎�uU�p����d����od�b闕�����b8s�;s]�чl�ؒ�k�c�}<sͱ��5	���tv2u�a�[lwk�Y��q�M��{d���Wfq�z�H:�v:W�t�m�q�ծ��b�Ƈ5ۍ���CE�s�\:Am��i�P��0��'�^�n*{I�wq`.�E�[�� ŻY�X뱻/g7�����s=�{5�:9�MS���ݖ��*��J��R��d����mq�n�D[�����2�S���<�U���;qg�g�k�L⵻��ǥ���)͊{'���u�)��k��y��X�{.K�˞9�s�ܘ;]���yym�c[�{BIvm�{Qp&cm��Ћ=���XƸ���<=[�a���n����m�r�4�;�:K��b��޼�74Y3�kn��+nמ�B�]��������튜v�� �b;&U�7[��'��D�˶�ݖ��n�í`)�
�4î��շ3�dC�m��b��\����רW�>�㓳�v�$,L�݆7MG�Ʒ�i�Mg��s�̓il.�8�g ��c�lk�q��8)�A�+Œ�L�7e6�\!Y��=&.A�[�v����!�c��j+8��G[m�l��i#&�G�;*s��mѮ��Z6�5���-ڞێ��%�+J��nM.|�����ԓ� ��댝6�G]�*���n��չ�+խm�\�5\�S� O��lt�v���NM������$�q�`�܏k.k�u\�7<��iP���������B�(��l"C1���p"�<�1���̶�:m�u��նM�OWj67��vCq��s�5�\#JWG�e���lɸM�^�[nӺ� v,��k�ew�GC������O[����ك]J\�یF�;�ȶU7nOA���ηʄs�ykqP��;��W�V��Ե����$XI���؄�J7�dls�]���ڌ���T;o]���ũ"�d��;,S�{Uj�>s�tI��͂K���ݼHk"�k�6��tJ�����SX1�q�gX�ju�ٔ�qڸ �1٢*�j�Bj��8��v����ݶ@�QуD!�u�mK�����c�ș�Kp�;{��r{<n����ŭle�r{����\q�vS�� �&�\�����S��ٷk �{y.3��(���$�8&P&����"t����1�諶ݢ�������ks�g��)ͱ�Mڇ�޷O�y8�7��E�vv�n��ηʧ<,ka9i{nx���26�s�e���G�i&M�<�6��j駭vԺ�M�m�\��\�e��rrq�]��I�ڻ2Rp���fA:�t��޳����I��r鮥�rS�fɣvjne�-�6�����+�����N��\d�{FE'm̅sn�Q�r8�N{yx�\��.b͢��ٹ]'i�NQz�隱q!�:��:��1x�������1�ulvC�Ȱx���ǐ��qٖ�=�;/9㐮�,77�\u۬�Т��\c%M��l��;r`�6�lt�<Dr�q��oOlC�m�v6D�;l�N�ٹ�d�I�m�q��ܭ%��i{v{��XN�	�uϜ�[�/!'B�����ۥ��'�{WOmM�2�q��e{=�!��nm®�Í%���W'���v[\���\����;��;\u�3��]���k��;�첲�zD�^!m���M�>C�ju��ټ�iy�d�\v����/s���O����x��;vp�]�N�mۂEe�W��a�m٬���Uz���Wlvf���>�k΂:�kL�R6z��9�Ϟ���ɴk���[u��$���{���w��K�[Y(�����1ۅ+y�Bt�]�K;���{q��Ϲ���[��:�̋��[�dk\j��J��Z��[���@��cz#���a�ͮ��Wb$}$v��p^�Ͳ�X��z�[kV�f7&i��0v��E�Dy��D�ٺG��8|�����E=/��s�n�,m��2B8�����o
�"��h���v���ݶ��[��+�n�l�;[�x���/6��9���'I�ka����b���m%[������9�v���V-�c)��[�-���z��a\��m�����nB���=����.��qf�e.K�nq]�n��<Y��ź8܀a��<��k��x�M�ۭ��S��P�������`�B�g:�9��s��J���۩c�5��W"9�\�O�M۵z˻���ݚtfD�;��؃�7Rm�����:9��;n��v5�^K�����6G���`�t\d�k�W�����w[1k���k��l��=ѧ�a#�v� �9Ѱ0G��+�q���I��юl��Dy6�{vH�ۍ6�Eɚ�0�[�܂Wndx�u�q��H���� �����Y�o,�Hۋ� ��D��«JrcT{ص�7i ._F�ts��e���`f97�c]=6�l�k��`E����[�snx9%�j��v+��\��]ALm�v�:�m9�su�[�8G����s1�8��Ak쾺�(�OA��w:���h��������-=tk��wVwk�M�^�Є�{n.K���X�����W�lwc{l�[b*%��q���Q��#+Kk�Qf*%Qcm�[��j5E�Z�-�+QEV��h���ūEmX����ˋ��iU��V�[F+Zڕ�����\�R#�`�kU�Um��eJ��0ۆ)���J��imX���F�j��֊�m��Pm��E�(U[eF��a`�kE[B��J�(�
�aZZ�YkB�Qm��b�"5��%(��a[Z�J
�e�Z�֔�F���h�F�E[�0�i�\R�Z�m�-kek*�F�Т��l�(ԩR�R���[mm�*6�ZԶ��aW-h�*�h�F�F�j�a�(��m*��Ee8[U�5J�81J�%T�[akm�[F�b��Z���EmTkb �VV�%����jRڊԨ�lҔ�"YZ%-���-F4Bƣj��*�ZZ+�Z[-�X�-hV�J�l���B�ж�R����[Z�@��mJ�UYL5�j�,�mFУK,D�bƉQ+X�iZ�EV�m�l���X�[�A�b��`�E����QE�R�L%YJ��������EA1.�$��[)��g'\g���k�]v7m��uv�o��ln�n�,c`�x�ݷ6xesrAN����uS�y�v��}n��L��kvU��G6��<C�gn+tn1̧f8i�밓�9���v5����m<�6��&4�nd��4<��ܾ�lbC8�����[{b#��Gg۸����|�y�4�-۵��v�c��\�t���ݡ�W�jx�;�-�����n޴�6�M �rkɂmkq�sr���R �gR������(��z��s���n[���\�N��vE��`g���.żK��Lƞ������q�0rgp[[{k���GGNN�M�n�������r�v#���������vܼvǵ���4�08�&����q�Q���uQc�p��yv)Q�n���mlV�� �*�N����=�lqݏh㲚�7\�t������"ed�c��rv������k4wj/i�bܸq�״�'ڴ�ݯn�읡'���wV����5�bt��۝՗�����q��񺝬�8ݺ����v��A���dɅ���r�Q�w��p�s.^�sq�t�'"O�:yD&8۱!�'�g���ۆއmQ�ڞ�{;Мg�^�d嗗㓮Q��Gv/7n�Ѷ�Hv�`��l<$m�h�ks�F�8v��mg��&�	Ӄq��ql���[��� WQI�^�G�yq�}>]��;�Mn�f�g���Ʃ��m��v:N���9��-�\�ȣ���UI�3��2�VS��'��ė\^�Clm�#N�x�y�����ۋ���-ћl�{v�h������^s���rmا�-F�;u���:u��۶����[�;�0x���ң��h� �ݲd�1�۴8�x�.ۇ�j�<]�\`�϶��t㋭�Pq�u��^g�})�U�!g�;��sp��{A6x��8�ٝ���pl�PMk�jF�8s�Ʋ��Z����T�.��W{���t� ��<��1�=�&�N�(nN8㰛������=�s�;d������|eS����8q�;nT��r{r<��N�nq�vLl��8rgÇ��p;p�*n����<�rv=��W�m�(����x28��r�e����G>y�v���T�m��+��<���gg��Nv�ɼ�C=���6\�"��C���?���=;��'�v�>$={1q$�D���N.�v���U~ϋ��n��ٯ��2�n�*E)�&����9����=uj��׻5@��ίW������Ѭ�-��%�m���nL�@SD�T��wR�6 [�ުAJ�~�3qNZ�Ț�]]X ���|�$�ίPNe�D9�&�PEM|Ou��샭��#~�q�u� ��uz��_vm��9=�ii��4n���fA�0�L�=�꒠@ ��ڿ����ۮ�̫� ��t�|���W� �ͻ��V���]1�F��A��L�S&w/Y���vp�V���#�ݭ��>�υ�f �_�;��dB��8Q96ꗩ��]�ު�7}ٵVj�]�=qJ;PL�M*
�7ޠ��pB'P�T���-�V�S��Rg4E�'p7L��X.$-�3�9�{�/nx�Zq�|n�K��X�%�O'��dȜuA�\
7�.1s�H*�>|���	ѝ�jW�N��]��gW�/�6��V�][�Ut���2�n�nE)�!d��%@�ݫ�� �k�;'[��Lր}���@ ��ݻ��iɉڙ�0Ȑ	}�:��Mn��I#�]0�H���ݻ��I%��5v�F�����Vw�/̪�9��2�D�J�dT8�뭰_��<��!�J7)��O�[��	�ݫ��|}���&��2>�n�GQ��$���s�c��t{��ۨ�t�rY�3n"$g��p>���L�d5��>�����$��٦�d��W�̶鄋�۷j�s��s"�	Ĺ*f׭z����c+7=|����;���ګ }�T1�Q�l�GLnѳ��o5T���870ʯ��^�� m���� |�S��{j�2�c&ʒ,_W=S/*ʉ�RcN�wЃBB� �+��9.�;5f#��/
k����й8Gb������o��C{��WclA��4�>"��Sm�Q)ȥ:��y]^�V҅V�Fs�w[y�ӹuv  �׻5_v�;�/�6��7$��V� ��۵dӃS�2��*$
~H��%�.=�LR��+K٠�oU�o �{�������ۥfgT�.�Iy��忷�V-x��7TOc<]x�T��giH�"��7n<r��ޜ� svƫ��;b9L�Q$���v];���nר ���H:�:�77~��w�[T� os�iPew�N��3!QIk��D��������s[���I#��>n�@+3:��gh�w(�<�5պ��~P�Y��N%��6�� �w����n��**�<��ΰm����t���i��9P�8�0�f�mW�"y�]Ѐy>� Y��Q@$�K�s�oKP�z3U�U:�n��!N��pӲ�Ud�W`�zehzoʁq�a���gF{9�qγ����K������'�S��� ��}%$+F8��U�� n+6|���M��(H-�(:��RA"w;5ص�����|jw�U��gz(�ͻVZ��g���z�B�ۅD��!4����b�O ۷i�@d�`1u�<)h썷������2��dJU�Wmz����}#m���w�ojzj����r3j+�>S��Q.TI��EC���cj�{���ufm�+��| 63�(��рz%L��/��^f��!,1l9�E/���T�7���X n9l�NײUI���=�sm�:3j) �F�f�7�BDqQHH��)�HƷ+c@D�~��6}�ٷv 7;g{���Ǯg�@]q�Q@eH��T8A�L2����݀�m}���.�N��.NQ5
n�BH$w{5شIInv�k���:`v:�����Z�B'�����&)�^k9�f�p�GQ}^^)S躚��!�ίC�X�
ce>�~���*�Z9ֺ����;��9��$n�޷>Q�˹݃�{V�+/��W"�n���ٽY�
cL�S�X�Ol7�@��n���%�����w����#���n'Y�����=�g�&���}�����c�cz�+p��ymW��Z���nc���$�;��K�㶳�[����u��Ӈ��ƭ����E���E�tlkuv�FW���v��X�:a:�wC�ZR�;���X;M���\k	�����t��ӣJ	��lcE��Zg4���$R�~#Jڇ_ �s�j� �s�j�(�T�e�{s+e����/{6��	�N�K%��D�M��v�P�'Ef����^� �^�m��  ���Pς!^Tx�Ȱ��Q.!˂T�E��uM����z��H�s��M�]{���>�3�j���{}�Tֹ@�)�S�$*(�u�
�r�bN���ʵ` �욯�@^FuG���/#��gi [ٗjͯ"-��rz+�q�U�l�;�$��dlհ�
�������z������v�zy��GA?/���}ƬrN�x{l�uv�P[��ڭ��Wk�R�iN~��{�{�~�L�j&�u����>��^�Ā����v��w�vF^m�m"v�&��d�!2��U�#
�5�lT��ߦ*'Xs^�h:G)?q����E��U��h�&�[�7��̥C+�D̾��NI�;�7|'�:z�X�B�H�욠�;�@7{�����no)ښ���D��a�)U|k��G�q��JC�]�>�Z�{螏g� @_l��^FuE9�G�K��B�0T8aN�e�����;���I$s�����w�� nvmУj��o��t�m�]�s�ɥA����D4L��:꾐 ;w6����}x�NN��sT�@n�mCt��f��f�F�a��O����t��e�MK�Ж�|�d�=v�m!]�ع�<�1[���N>�?8���[5q.L��/�4/��/L�W�6 >��ۻ�WU[�;Vuؾ�
c�a�PI���w��/�<H�I#���l�m�ܛ���8���gz�{��Wh�����j���v�@*�>P�jS���uRR ���j�v�I-��~œ��޿c�-��w�cR� �����Zt��Y�'�R�$��r�y�����8B+�i%��\�#�_MOsc̲���
w�Ύ���Ψn� ܾ۵`�<V8rL9�D�Toa�3}�u�ȷ��� �/��{}�v�՝�N2���NyA$����X��QJ&�PH�8�����v i���;�y�U2���vTP |w_m݌@#c;a�����+to�T��`IS�Tλ������-��c;)���ai�����.��8o�����Ģ&	����uR6m��6� �;c��,+]\�&���E ��wa��2y�D��
%�QA�iMੳ���{f�#�V{�՛�v��vE}C���S�E{��F�s0+�� ��)����شJ-Y�Jh��鏠�����o�u��v0��uQW	��P��9jS���+����{.�F��W޼��U�|�23r/�%{�&e�eA�hR�}Yj��Jzx�E"��o�̈�]��mP��op0 ����E�M�=�;}}��+
��x0	�x0������D�*(��K�s�U�JhH�rΨ9��Nmo]��!.��l�N�u�oP��Ψ��w�Gl��@�����~�����;c�8�g�tuq�ᖳ�zmk�p��=���
��?(�"bJ���f�~���܍ʊ>@ ���u}�r��[f���cm�F�J�g�px�CD��������T�^m:UD�*�w���r{
n�^�ފ����Ⱥ��[{��oֺp��D� !eT?%��E �3�R d�".W�3ך���o  F��n���P��r��!�
aϰ��m��<J��duTS`^�ފ�{Y�WRt��u�@!E���w�7JPŁ��������{j��~�3�ӑ����3W�د�:��@|mgm�Vv.W횝r���p��b6q�W"T/X="ds}�������kz?3�E]f��ɝL�b+�T�Š��YL+�׈�+}�Q����~$��$qv,g�B��e��9�g�/vӭ�p�<�Y,����n�Ɩ�p��1�+v�jȶA��՞f첇]�t㊝�;p����W.t6��N��y�_=���w��ݒ��{3�`ܜ�m����h�p�;t�'>�6.DKrk�c��<fq1]�u�kC�ȝd���u5=]�Y��1b3��ӈ���ϱ�۳����qY�S�x��ti�F6����ò�������f�M��G$��0v�tj���~���js�g|oe%4 ����:ŵ��v�SPbÕ��5����4ICv/���_S������ ׯ⯿X�&=�վ�����=�����QHK^v݋E$x���]�Q��Q��.s��D4L�*(�u�Aջ�j��=�Q����2=� �c:��@�����E��A
~�(�%E$'����IwU8������;/v�� ��l�=�O�<8����ѕ褀ʑ���p7
a�R6n��� {��S��m�����WQ�ʎ�$��v��ڱ� ��;��^�������@�'D ���g0n:[��R5غs�͵s.fT�2������f!ĵ)��V{��@|��W` �횤�<[�#�zZ�5�_�  ̾۵`��X��D��0��T���O�<eS������긳��aZ�zX��h�1�G<�	�DԻ^��Ў87�'nE�e0���]��Q������c'�R�{���Q(;�������횡��Dc�w���Gk��~�<���Z@) �W�~�B@�7k�| c���Ǒ]_�b@��ڿ�m���5F��D�(����g���^�n�չ6��	�f�� 3;f����QѝpW��P^�>+�ww�K�zPP�O�!e8~H������Χ�A싑����ɶ�����f]�D�ٻ/�B�3��T���bwX���A�[W#vϩ�7��-�<烪�j�e�O�兮խ�?���\��.����~�����{����@$�w��2���ΫA�k����h��Y���^�4�X&e��Z�����)�X\��]�_eb���٪@�{���n�/s35��`z��&T˘r�EToe|���q��t/�S��db�W�RNk{��[M��>%���)�o��6��ΐ&���A"�u��'Q��d�z��`����K46@��4ZYm�l�B<�ѳ#��s���Kl�G����$}Q⒘�'�.＂�����+{ג]%7hJ���}�uo/Kˏ4�)�Z�&Ay�Ol���4��MCwj˳�SY]�4\�^wj6�3e�<�-��Z��#~[�nN�m�a��:����2*���C0حB�Y�qGmb���x3|��1A*�Ў�T��Ò�6�8+�������&R^�`��i��=�v͊����2���oB�S�B�p�<�a�_�I{�Ծ��/�aw`�~5=�� W�Cq&��>��o�{�X;���n�ᘯo"����h1�L�|�=wa)1<��g��s�ӓ
sVrڒ���s��SlҜ��޽ۗ��8����dt*�	U�b�ͼW���L��e��X�k]p��Mk��_��W&e*�*n�J����=g�1�R�n������<"��nF���rR�33���|nXE��e���<T5rɭj�ӵ�O$�"�4G��-!���J���yi4�1�ܥ�2.�W_R���k�z��@�E��޾�S�9��a^��
n���Ȭ�HR�FcW�u���%�Y�g��K�����-�w���-v���:��[U�M����4��6�b�I�!���I5o��!M[��7�x��U������<��	UZ��ɍĮ�T���I��'x�������Ւ�j4^�V�S(��VE)�R� ��V�U�(%�F��چ�ba�[F��"
T� �%��YYl�X[R�ҖX�Z�+QZ�%E-���d��-��k,Dm,DU��m�����+B��*
�V�QdX-�+V�Q��8d��&(�(��і%�F���[
�*6Q�*�h-UQ�kIl�ˆ`��`�X��X��JQ��Q�*(��R��-��"(�m-�1T@��1����T��j6��Q����)i,bֵ�h+mk(�0�pĭE��-J-��E��EY�bƍ��"�����-J��+�V*a���-�i*�p�%���p�h
Q�[Q����cl��[VڱlZʶª��V`�X��-�"*[P*�����X�����R�
�)F�T�X�c%dJZ[S	X�J2��`��Uڪ��F�R�DP���Ѷ�X�IV0E�"��b$��Qm�[k+`֣���F�+T���UJ�-�#mJ�����Dm��p��[YZT�kP��Բ1ABҩ�z����[e��ؤ�`��Q@}9��&"fd�%8aN�m�7�fJݪ�1��<'Vc�P }y���n_m��/o�p���*ߒ�cٱJ�t��z	|�e�Ժ۔JK��b�m��7x��Sy@���Y�w�2#)�o�ܩ��~T��(��rC �8R�1�9ݜV��hǆ�v�j��-��mjP+�����#ץ
%ɱ� �mM ���H���ۻ	�;`��|sTGm�h����]H��T8qL9�:�[wcq�7o,d;��;����@���ڵc��nj)��_�O���ӉQ.�N��/�|�u��N����Y�7��gw�b� 7�:����k;n��ES����Y
TH���֚�p�~�q}�J@ >��ۻ� nvN����.0��	���"��Y�*����7-'vgzy\���4T׎2�7^Y9vZ�y��	Va��/C�Y��rlV�ȃ�J��a%7�JTLDI�ɖ�QD����` =������]3��"y  ��{� �̯7@�_d�λ�#��M����Jn���-ԳU'rvnv�qN���&���<6�#���=�X�����|&G2G2̎Gx۪R �V��;@|7;&��~��/qNߜׯ�����]�w`���A
~�(�%Cl���7��o���Z�L�d� 2����H���d�4RU4/o��m��T����Á��˚�oշN���^�~�
z+%�'�=QH ���M���5@��^"�NeĸR�:f�޽U�lc�8���{.�� ��U� ^�uE�1��`8:�d�~�u��c�z;�f\�D�H�_�줽G�q�O҂���s�T���]�H���/�����F�h,�T�uv
R�Mք�����J��,���ۀ��t*���j�����a��vf[mY�ePzG-��I��|6��`o��'�A;�k��9D�`��0����@��9��y6.#,j�m��s�k�;ѳ�W���(�� r��d�]S�v�b[���
b����脹�ϣh�=r)���z��n�<u�e�&1���=(ζ�۷m�'��t�nmκ���%,���͹'��Y����N��������{�we�n�Q��!�DT\�띗�}ywi��dl�2%4���۬�{C�1���y���:v����
v�;cC��pWϟ��dt���q�����$ =��� >����.<�\ڵ�fW�wcWl����|�*e���;*k�u���)�g{*�X| <���t�gTP 	�=۪��F���D9$��q�T�B /L�R� (n���5�^�fj�e��P���ڊ@mH��p4��&�#f�n�����F5�>n�9��� >[��Q@ ��]<�Õ3�px$���4_�����ˉq��*��r�H/�A{}�N��&9�)0�����j�6^�mE {}�vg���?508M�bY*w*N�����q��v֬�f�Ş��������>��2-�*�y]��M��v� ^�m�wʢ�[�jN�M*e�v�R/3đ0C$	��QD����"�N�>��#/����;�'V�srZ[���4׼)n�!�w��ߖ,6_�0QQ�*D[X�=3J=E�)�~�9W:�=]�l��ݨ� ���ۻ�eu�7y��YY��G4J�%w��@ ݽڻAT(�+#�5@��� ���$W���о�:���F���������| {�W�C�n�;j� �A��,�i�5�o"h�I	qZ��6��n��D�I�6n���o���nU��� f����ڿ�`2�g��C�&���;�klt�Khlp�%�R��:Ɏk5{��*e.;NS�=:�E$8����߻�ڑ�K>�Er6Mʥ!�{��v6��5A��v���a���|^��Ӳ�Bᩅ2LĠ�U����,&{0¯Ԥl7;n�� _l�/�MXG"j�f�t���t�D��r9��QD����` =���z��q!(��3b���XQ�U��!϶r,J�`�x���hY�sƱ���p0ZB��Fg\B�[NS��\"z�b���tgd����Y�ٻt���E��Pmo��>j%J����/�v���Q
�NQ���իl���b�����lm�=�V$A�I�u��QzP���(�3�A�T��÷��wYO���+v ^�ۻ� F��Ǜ�܎ڊA=�?>0�z/Bdc��ܹⴸ|�Se-�bM�ݣ�Y�[E������#�$�1�(LMw�M����PK���0@nGmC~<��ZUU�݌@$lvlW�U�9��ԎaI��#d�RVs�eg,��g�\��wh�P���>܎ڊ@�5n��8�Z��u����lU�p�"bT*�ӯ�M6��)$��v���Ɋ�T�L�n�`$��76(�X��v�a(�%@��FQ� ����Us���ŷ�o���Қ �;j)ay���T���C�;�k<���I�f%ll�g�j�4����h�㇯dNa����/��k��;\��w��Lef��7Ƈ6�MY����?������L)|�J�%��_UH$N�n�l����pg!K����$�bΨi �
�;m�����s�-�j��О�7l����L2�_f�=v�a�v�Uc�a����r��3ۋ�`!�(�3{*����gze�vݶyJU�K!V)�lw8�Iyњ��%�(�`��2f%��Z����e[�	T9iUnKI ����W�|�;j���&Ɍ��Mǝ*Y��r����DS�+����v�� m���×�=� ��6����;n�>*�.%˘�T*��i�Ѿ�N���3�� o��RR6 ��ڦ� �݌��QU�mw+���LeTP
n���"#�)�7{+U�����R�ͽ�o���;ލ������݊�z�x�r�}��P����pl�ʓA��*b�E�#�ܥR.���������v� ��9�|��pYֹ��J��X��χ�&�BL���	�U��qgs��cn���&ⓞg��C���T��^�."�n��n�.�7H���i����.�x{[��Z�gw��v�`�e���WA���^�pU��/8jZ���΃�������ul�rt8�9t0�n�16p����/c�w=�lby�w3��42�؈�z�y��֎z�v=,�.��t�[Uڄ��)!��B�ƚݙk�cv���MٜE�y�3tѸh��pk�.��Q�߃���L�Ri�	ò�H ��W`��;�7����ŗ�3�w�� ggm݄^��#�J���R�{j(A��j�◯�v�� �ۛ�vI#���i7K=�9=��d����.X���HPź���y�Iz7iE-+��{�` y��Wc �ޝҕ��nT�c�H�W��}U$�S� ��T� ;gt����_Tdl�W��7����*�
d��T/Pot�"� oީ+1��zD������uC ܋��x�m����CG�Z����Q�1%J0f�:ɳtsc�23���Mkkp����7��ߟ�?�%t9R�Q���v��36u��r+�(".c]�X��컱�������gx=0�q�S.e�8��H.�.!���N��jY�?=��0�f�+/�f(��lM��rc�pv����p܋�W��A��E��O��-�z���4�"�  �y�ix$�Hn}ZYtܩ�E {6�:��X�5>�.�9XE���lD�n!�%E�Ӵ�B�*;ä�	܆Uy߷�xD��Ϫ� y;�}CnTw��+�T��I,�Uk㹸��Z��e�Iy+��|������=���z���i�mѽ;�*�]��T�2���:n:������R���1�W.� L�H 7�z� ���g>��z���teZv�	NLO�A	�W���nY��u��x�����͈x�#Ї�\��w���)s0L@��a��4���J�ngmU��3��CV����wEP�3*z�@)ڝRB&"�T�TQ;��v����8�l@��G��s�W� ���M�d��9�N1�g�;�s�Dzˏ��s,��Ole�;sv��I%䨐S���vt՗7�s:�7J>�FXQ�*����"sH���Wع_i;�/z�-ٔ��#6��3�j^mj�/f2�D�v��q�Z+�Tt���u���I{~��`$��}�`Z"����"T7䒡�"wf�,�N��{�y]����ݻ��@����QL.ۜ���nG�-Á���M�ɿI�$���.~Wv��'����jsg�� ���ۿ�g��lҢp� ����.�DI*Q
A�9 ��'<�I`6�������)q\U����~��ˣ�)H�;�F{� }��v	 /{e�%s����(H�l���:�Iy'���iX��>�r9" UHoe*d�3�3��~�ꋭ($�nn�	 ���ɲ	;�=j�{�pV��5�G)!G*S=7{+U� �7k�P K�u�x�V���ۻ��٥@�w��B�q�S.e��=эV��@�I�$����P	�٦H̬֯Y���/����޸����[�]&"֫��oFƯfL�iۉΎ���g���¾۩��G�����[�c]�!1�q�w�����{Z�& ���bkX�J-̏������N����@ ��vk��s#�6{�zu�ׇf5�)��)�e6�#�z��F���z^�Z�N�e�/g��խb?�� �@đ1]�[ۻH$�;۳O� �OQA>��}�M[�omSm�A��>t�]x��	JP"�٨ꤠ&����<u���g3s:�	�ɦ�̞�� "ze�N2�.��zՇǖ݀��.G$D
��ez��A��ޯ�lA��{#;��N�f���3�� ��_P��OQH	��9!)D�F59���:!�ݼ�V�-#<��d�^���I$�Yy�|*k'��{z�O�2�f���"=
e��\�,��OteW�{�W��4���M�?0�$���'�m�H��۵e��QQm��{�b�f"��͝�T�u�H)��FE��:hdv���\m����f숁��NI��q�d<�ʵ�5������nf��<��D�S�G�p��U:3�1�$q�k�����ӲHj��g�gJ.�)<v�;���6�K�{g�ǆW�}��c����x�b�
�[O+�t�s�=�A�F��=��/����M�Q�M�=����$u}0@:�M�~'�:��l��r��	�b��e�Y���̽�����q�2�}���}cG�����o5+��
��N��ue��/{xp0�=���:�O���ujK��Ƚ���'%�9=��!�)�3VkB�JW�K�/Xg���v�iZY0W!;Vy���M^e'�Tv�}���a��CL�����\�����;��4p�Q^�>���z�������>�����:K���$+�m��F��*��k��&D�6o�p�=�o5h(�]󮱗�E[T�Q�ܝ*�ː�=��0�ԝv6�6P<�������K.؞��o�gsg&"��g	b�wqy#�i�����Jz�<Ft�Z���F�?a5K�	�j^,$:=R˗k�e� 8��ʅ3�r�dU�)4 ;�&��nk�i�8��@k/*��j�Ǵ�v��)��L��V��<��'M�3���H�ɣ&/�j�j]�rl)q��J���o�t�{/��ĴZ1J/`�b�,�E�����
��=��w��M�֎5XXN(����g��a�c"
"*���iU��ZU��K[mEEEE��Dh����UL[���Q��qK�+*��؅F��aU�*6��V
��E��6�A�6�h*8j
��)�Xa*,k
VQ1kŔ�0L#Ak��E����Z��(�H�(8�
��E0�*�� [b�Q�����֩Tam�AEb#b�*[UA��aDY�Z*"-Ÿ)[E�Fئ����j�D��P�QR⩋(X��b)YKeE��+m���T����lD*J�D��1�V"[UFA)[U(ڶ,�QiVآA
�F
�T�ia�T�TB�UQ�X�+hUJ�cF�%j�F(�Ɣ��e���Z�%�Pm�lUm��%B�E��m(��Pm��b�Qc1h��
(Ҕqj",Ŭ��E+�T�5(�-,��-j�k-(#iF�H���AeT�X��kYmUUX�*V�Pm
2ڡR��KJ��DZՊ2���ʶ����R,����*��Բ1"��b��J�)lm��%�eE-��E��,Z�QA���"��l0�QU��)�-��TV��"ZJ�H��X5h���1�����PXs��ū��nx�Żh�6�m��9��CQs��g��7 dNh��qZ#k��<sѤ4��{X�Z{���pz�V'��w[.z��jݺA�_2v���v|���^7Z]�=@�GOCԣ��aӒv�cI���nݎq��s���n��rZ����O���ŹLcv�B;ϙ_a�贕#^�Ȫ]=us����nw���2�����닉�zN��wV��Nq�s�	�ϵ:��vwmtA�;O=������\ױs;�i83�	Ӌw`7N����rq
�=�=�R8p\v�9�1�{f�c1���:�;vH`Nr����-���r]�E�w1�i��}����^i�v��d{D�Xʎ�9�1��:b񷮽��/8m����3H�^K]���Z��{�
��/'�c�t��d��>��1������F���^zݯ
̦+\<�7�6��nz�����^�gŒ��Д89��9�q۞��u]�mlO`q�:d���U����ӑ'����c�ym�vC����ܧn�zSwY�KQB���ݷ'E�˸2t:�&�@�]U��R<�3��E�E۷:��]=/Bk�j�k'��'��p)v��ۮ�8�z��ݽ�N��뎱��!ƍx�^.i����ېɎ�Kt]b���iRb�z�;A�`�t�p'�+t�s��Lp�m�Z@�p�v:v�k�c3�'k�<�vS����;=�M��e�-l]��۹5n9yUs��6�#d #ę=� 8�y.�we�n����W=cvK���m��f�v9���<�m�ͬ�˱Q���tnz;Y�Ɏ�i.9����/�����Z�9�s������:���C����u��vZѬ���u՜n���}C�HK�jX�wI۵���\vLS���W.��i���j<`�=�]���5ɸ�\뛷k�e��m<E�=��8��V�)b&b�*9s�aim�S��nc����}<���]�J���ď��8ǣfg��B�]��O@]��{�����u}7=b����kZ�q1�rfn5˞tps�GG�d3g�ё7�����_V�����n���JH�:ݞ��]�5<�^ rQ<]8��ݗu�C\�e��:.���w)�.�kRl��#������N���k����k{�7
��:�{^�G6�9�WU�l���^�j�7K��.�l]�qy�8�c�-��k��
s��).�ά�q԰��&7�V�ڜ�c���lν�Z�^��J|�����l'*�ne�=�P vdw� 2���Q���s�U����76$��'��>�����p��Z���6j�����Lu��K���>���잢���wc_+Uq5�rL�͝��u�.P$)@�y�����Wa�F�{�}s�� _d��<�����`'�J��
����m�V�>��OFxt��wf�݃g���>�6!nҽ�ͣ�%v��	���
�P$)T`S��l�I$ww]9n������z����6|^�mڱ� �ݟ=ɋ��J�Տ�&>%�Lʒ&c���L�m��78��z_SsΞ8X������.��Z(��
yn7�D��su�iw�f��~��gڰ�͋�@ ���j�Տ�Hɑ��2j	*gf�,��J���l�[�_�8���&u�����ro�0�.��P�P�k��9D#q}3���7v��4g�E��>;Wz������y�����=칥�_xJ^I$���l� ����2	?���:O˽�k�I8��r��K�$MW�MV���>@|{v����=Ӯ�B�=|�����7nұ����TR.�\I�)@�3�_���)kб�/�f�<$���s�� >3�f���;�=�������
�u{���<=���T�/RG����$�,�r����ux�^�띷�n�O���gTRA]���d�o�ϟ?��O�[Zr��]p�{n9�k�Ϯ6z9�sv1���=����qQ������G�"��qȜ�ۿ����>�@-�Ψ��������+@Y;�w�h��Y��E���2��\�*)�eW��u�L�gk��X��ܚ��-�Ψ� GVyz:~���M�;Q�ǘ7*�
a�6ɜ�� �7�W� |�Y�-L�O��[N�8f~�V3w�s�׎�PI=�8����9��!�U	c!��%�0n�7����m������xߠ�0U;�=-����{�~�{��A/�ܚ$���Ϝ0��&�Ϣ&��ak���B��hM�
)�RFv��,@}y��P	�����l��;I��ӊ���F�� � �F�c�	���TE�z=Gn_�:�j�H327� �fvݫ�^�k�J�S�C��5����ݎ��"M�c.��j諦�&Ş��xo��p�����W yە���7�7ï�fgm݃�7�jz��+RVHU�ϛn��z�H�վpB*)Æ�w��Z'�/f���wS^Iy$;2v�@ ���v6��68��w�~��[�4�
%��L�RQD�FU@$���i$��l=�hUEP��S��=���3;nՄo�)z�8P�E�{{޽꺘U���� ���R�@ /3���I���ݞd���ש:1-)�����m�R�JS����!���.\,}�n�A�����w��Hw�{b/�U{��6#� ��i�$>��j�������7HrD�$~���J��G~�t���|77��G,��S��Avf�شW�Ion��4�4�o��/���>�}�Ͼ��&�^Jk��k�f��[iL���m�N�P9�KR"f"o^.8��%(�W5T��{��N� 4���73^*�w�(����$�=o�6&=BH5b$" Tޝ׳@(�s[3w7�����د3������m�ң�6�	��xo������A������v�4�ښ �7��8��co��� �v��ӷb����H�\|�˕'��u�qKdĤ�����ly$6;v, Y�=C����V�N^B9��j�F}�`�(N)�P�L�4y���O��>Q��S����Uh݊��fd�L%{W�b���{r��i�L�&�M�op��y2"�l��wH�i���F��L�֌�i��
��-ގ���[�T?I&�}�w���Z�V����Q�>����������PS���ix�Dk�8W��F[/��h.=�s�:�r%J��EM.�{7��
ݗg�py�тȮR�uv�>g�ܜ����ɰ�+��=�Ch�OX7&���hlpx�'�g6�wO�-�c=W	��Nݮ]��'�����W6�m��N�ƛ<��g�5�ڼ�v�=f�W'ex�{]�n�<j6��k�jͧ�(��x&���v�p\>yE��uu���0���RR����h+ی-�����?�N`�'ߑ��۵`�	��fd��2�ߵ]����^�+aѻ�J�J� ��%"�FMGU}}w���g,�3}^�ʺ�� F��7I���7A��3b.T���D�V�*��`6�J�B"TweM  ���T�f�=�:#sӵU 27v)*fOQ_��<8P� Cn*+�w�o���r����t����'h��H��ݺ*#}����,b�@�<qʏ��r����lBI����j����ԫ�	/Dv�l ���@�۷+#fm�=��J�2��%�`;�q` G�������ָ9�w*6�r�;��Yӏ�~���l�ɞ���L�{��t����ݻ��z�_��e��5ܵL:�~h���vm2�q`��at�ZQ��&�$ w�buY��)y�5`�Dە�|:�}��
���B�Z�DK��݊�H&�oYF�P�pe�|�(��]�f*���3����6b> y����Z�H$����t�@�3����Y�{��K���D�B*��]5_ ��J� �c��W1�w�� >37�� ���j�[���ʙ��@�_���w��vM^G �*}H���% �;v��u�v�=�d���dB�"d!������oLݩ�q�q�S��I+�� 3���� O�;b�l��ƶY��!"HJf	�y���vì�$�t���z�7V��N�5u�}�ۮ8S*>je̳c�';&��ݫ�����T�wFƩnQѼ�}��H �ݻ�Q�gG�Cp8S��A>�S@D�)����2{=>π@/��;7n����T1�������h�%?c�9�0IT��������;c��*�s^�a���g��w��b�s�BlN��eqX4t{.y������&��CMս��E3O� 4D�䘀}72�{~  ]���$ؑ�s��� lg�T�iՌo�%KD"�ٮ��,��v�D� �VU;�Fn�P -��S��H����݀��ͻJ�۱��ʙ��z�6�<�K{6h���D�uZN�d$���]�@ tflUA��>m���3�z|�{����?>��,��Ɛ6n4��n��[�le�A�v<��ͷ����o�y�jö~��|�����Lͥ4 ۙަݭn�|Wlɷm��I^]�4�K��ȏ2L����ɪ��g�ّ�.��Ӿ���  ������S�>�؏]�w&6l��]�n�#}��F �
�QH ���M6�t���+�=s�}��n�FgEP����:�+!?s���.%�������z���7Guǩ ������Gw;^�Q���SCMeU��)(p�5�����׎���`�b�����=��3����bVl�M�Ν���rV��o�a���ٟ}��)�� ���T�?X�ډQ" &z+��$�I^���ګ��"+v��/`��s���Ks6�i/$��v��ӓjn�f�ۘ�R��	N ��9i�8�U�Jq75�u��ق�����Mû8z �W������8�*fFD5��q���Hٳ�@ ��ۻH2}�\��o�yS�ި�C�6h����"12
C����f�i�}��A;�f�}4 ���:� ���X�۟j��HF�zwS�?{��G��A�z�+�ꪾ���ڵ`���E�\���{�b�y����|����ۻ���6	�!9U�	�An&̥0F-��7�>� 6m��݀���9�qӹ$<=���٢�A�Xe�RbLK;SZ� �W�hfU2-�{��u_�x�I,������/A���GN���&�E�z���F�6�}8:v��\��&�Q�JüE�$�,��ߒK�:�$l3����r-�Q�����f�ndY��~�����{��߿��]̞�x��Uqt��tk[��T�X�0��6r��Mv�;j,�������v� �1���u���s�(W��c/c���l�X�L��՜\Rvg���q��dK�x��w �q�#����õ��%�[�=s8�������^v�q�s�j�7hŻv.�}��xv�u�ǫ���;�=��6o0t���9�wf4ȶ��b�qb�K�M�teꛋ�s͎w(-�u��lY�e�`�kItܯR����v�h�2c4�?�ɴ�pú�}���%g1d�+%O߾����~f$�0�>� t���$�ȳ��}3�ӿ�����͉�~��f�f�J��S߻�����0�x{��U�d�s[�:m'#�a=�}�C,�%ed�{?n�_�'������2ɇ0ɇ0Ʉ������2~OÆL2�VT�;�u���a����{�~����<��a���7�>]����9-���&�����~?3��3�{�tq�g��3���lo��i��0}zA������O߬�%�f0�L'�߻�e�N2a w�r�ȟ31);>��~0|+�hY>�vT�zO�B���/z������e$�0��3	�w��2ͧf A�@#�k�}̬��Y�_��/~�:�јf*{�s���?30wI���p\M�fRq�0�Ʒ�L�%ed�Řa��?h�2ɇ��}��sO�o�0Ʉ������O���& ��)����2��a��L3=���}X>}Z�q��?�w�a]�D(�.cK�u&۔���n�n,����D��s;�JVv�e�RbL}�G̏�������?D+%Xz����4�YP(%@�����8��Xy�z���iKN{�w@p� Ґ�C�~��C.�>�����\91�\�h�����D>G�G�~_�C* pOe���ƣA�H��q���?��H���y!;ܖ���c�ɣ76��2��;�zY�0m��YS�p�-��ܫ�x{�����Ls[���B�%ac
��~�2�c
��P;������N2�~�0𛏶�b��EF_P�,��=f�&&s��aذ7÷�~�2�ܴ�����ѾR��Z
�1���~��8�<sC���@�p@�P+*w���e�d�Q%@���}�l80�,߹��(�
bRA~|,���ﺀ�b�7��w��i&��d�+���C)`������$#R
{�����w��g3{�g�> �1����v0*^yߝ�ɘ��q�vpI���tq ��%e*}����$��7�c���q������~���Xm�IA
���~�q �q�����}���9���������~���#?��F�Y쬛b��ڢ]��Ug�m��jk;��^��(������������>桔��!K@��������0*_~��l$�9���U״1}>� 	�qZ��H�$ACb���h�
�G_.e���\na�>���8��VOw��n{�>��:������3L�P(�����gk�!m=�｠8���<N�ѿot`��1�)����
��7-Lf�&��q'��>��� VQ���T��｣�8�IXP�#�G�W�`�Q�ֲz�}]�ec�����u���ۃ*�ͨt�ʎ�[K�2k��)L�t..Z�.ųݰ��A>�]V�̨���Y�q�A|����k�rUr�F/jV̇��j>�+��ɓ��zI2��x���g�/���[^T�!a>�m�ĳj\ɵڲ�f�����F��L�2z})�^�*��L�}��h��]f)㻝UF����Ɉ��v-꽂v9�Y�'?mҰ�ւ�l��u��8��d�!a٘!�]Yy3�S��fT��T�� ��ɹ2��F��]j4%�=��}��v5}O��V1�g!os8�"e���P[�T"�S�٭£��0_��&�[Y��oĪ�Ju���.�͸�[��NI�[&=�nn�gn�kN�z�l"pz:���$���}݌�D�{�gP���ڧ�� ��t�+s��"�몹��@]���T�Q=S��I[і���fe0���=�}_����.Ln\*�=�]�M|���r��ۤ	�x1왧ڹ'b몇b��hwrZ	F�j����i�����Y�%O-�)��B�;k%��!�ńEjo)x�H\��{B����`w�şZ��	�!8m+��mdK�����xdqc�U��Xmm:�*��AW�t���ƙѲ_�n�莣nkI͞��w�08
R�X��4�X��*�S�-�#�������s�S<��O}�j5�ws�.�Z��N�d��6Ӊ*ӄj'�=�Κxr�wIӥ߯��F��<:��	��{�{��=��{��m���;~�h*ޤ�0����u���h"�PcmX��-j(�j�F����X���1F(���-�J+F�KETEZ�T�DE��mZ�
�L�V.)UV҈��b�b��D�*U�m����QF��h�
*��eJ*� ֠�	�S
1AD��)m-��b�U����ZTEF��UQ4QQbEETX���X�b��ˊ����֥����UT
a(��1b4b6�%*TmD**���4� �bZTQm( ���+,e���j�" ��*(",Q��m
��kUC	b�1V�"�1Z����,���"����e��R��*�(�iEQ`���UF�Im�UEQ)J�@V+j،PTX�"+���DF-j�A���)�EU0���Eڪa�a����[QUb�**�`�"��Pb*�-UcS�R�(%��AU�Z�DF*"��0�Dcm��U�,b�[Z�*�
�+U1AF �T��TEV�F�1����G���8h�n.X2( �V2�0�QjW�	 s9�tH)'�O~���2peH)=���h���,�D�&e%h<	���;�Mg��|��HrZA@ι��7�B��Z��}��{`q8 T������2��w�s�?��J��$�T>���h�0�,7��_�k���m�1�q�T�}���J�H,=o�63L��������=�ل
����m��� �w��9H6���?o�C.�O~��������{��I�N�ӧr��n�+�
�<^]����9��VA��=���1���?w���������|$ϻ�tq8�R+%O�w���'�J°�)�~�ۆXm�Iwc�ŵy�[�yw���Y�G}OhY��+%S����ND��S���[p8.&�08�����$)iw~�_�������;߀���H/Fl`T��}���@�P+,Oc���2���� dȻǘ��h��C�<,>��]�s.L[����4�l*{{ߴC�(�d��=o�i �T�����8��^{����
ԅ�����R�+P�?o�C.�/�~a(RLJ
C YG�o�do=�eO�����3��d��~�������°�����2�R
M�}ߴq���}_}olu������⨻��[�)�Ţ�f1��@�P�al��j3Ba/Lyܽ#hd��}��w� 7޳|]�lR�)��2�ڼ���nL�~ x}8����eO��ߴND�5��o*�L��[q]�Aa��}�뤅���on���q��{[������q� �O���`q8 T�eOc�;�e�*AB�����8Ñ�a}��=����2�߭��D�%@��a�e��iĩ��}s�5��\��e�#n�ǒ:6�Tb��߿�|���`8���>�
���{A�$����������2VT
�����6��X�FFL��#�BC�w� dxx"�c/��πD,��.P��A�S� A GW}A��O�y���Ҙ�g����}��q
$��=����aRQ
������$N��ϻ��w�;�!��P�,��F}�)A�L!�`pk\���I!e�{�w�7�B��[N���<�y������~O�*X�Ybw��C,�%B��Q���h�Aa����˙rb�8�w0�
�o[���sn�����q&+%X}u��7�JʐP;���H,�Dx$�g}� QؾS0tE����w)
�c��e��?p�n��8�\9nM����sFӠ�YFJ�S3�� 2���|�n���X>�UϾ�2�q�ID*J'~�~��N2�J�����' �@���_����3��|�닕���٪�~��7f�&�L��Cv\�AM�+rL!>�B5%�{e���؉���O��z��f	7����{��q����Qs�pm@�1�����G�/�"Cs���Xg���77:���'�q��m�����c")d(��+.LD��<m���c��ů�U�f�\�Ѵm�iű�ۙ�OU����P�e��X�M�N�֬��&�$�M[q.���-�״�fN�:]c=1�'�Y�Tc�E��m�F��>3�ۗW��=-Mي���=���n.����]ig`HRut������]�t����o�.nL����H,?^k���!m �w����HV�*AJ{�����q�gL�'Ӏ>D8�u�'��Ȁ��
!�}ߴq�V~�W�k���m�1�q�T�}��C�(�d���?g�]{�,5u�h�4�YP*T��w�H,5 ��߽�99H4�)]S�$g�����g�"��r��Us�g�`a6$����8�Y�J�2T����q'�J°�=�����S�����硖aRT*J��{�d�+%ed�ʞ�~�����N��%��)�J��_�('��ȥ�@^�9ִr�<ZB�������)
сZ�����h�"J VT�?}�C,�����g<���e$�T5�{�8Ì+�e�˙rb�8�w��
����"Ib ����u�}�^��O�^��wgjAHP�����9H4)
÷���2�S�.?z��}W�C�ٸ�Gu�Y�v2u mAs���Sr۳xq��6A��OĶ�&b'֯�(PL&�d�I[_�{>��ND
�*AO����ĜB�+
°��ﻸe��'����y���ۿ�繟Rd�����N2�VVJʟ{�{D�'7_m�\S.nL���X�a�߹�e!�H$=ǟ9�3������wtT�U��wwK<�Jޚg�����������ok�2'��Y:�a���\��#P;�lt�5^S��=	 ���׾ѿ�B��Z
�������p@�P+���a�m��RT���7yu�9���x�<|�Ä��m�1�q �=ﻠ��%ea���6ͲQ��T����yއ<�������R������)����a�������9ʮf&%* A���Yx85ْq4Fp;�!Y�߿jHlH'~��D4�({/s��uV(�D� �J����O��ȏ��hzȲ Y8��F
Ra`�g��Xcz�a���!e�{�w�7�HWXu�.�;�R
o��{�8�
���ﻘi�*T(�{�h�A>����NԌ@S�DǌD"'�vy���F����V�z�d���k�m��[�����m�rb�8�~�X|§s��A�$��������4ɶT
%@�{�l��`\m�1�g͝�����k����A���=���v��}��~0c8�[�8v�=��sG82V_��{�}�q�"���~��'�+
°���0�AI�
����w�d�ʐY*_���d>���,�8͢a	38�q�а7��~�Cc��HYh�{���R���9����>����?)B~�>�]�B�RA׵� �˟�e82��I�Ƨ�70��4Bm�9:?i�97�?���8�ޏ�<����q5���Z��8�����{�x���H�@T���;��wP�6�R
}��H,9�{��8p�8ʹ�70�aQ=�u��A}�i�#��OoP�&�P,J�y߻��08`V��y!ۿu ���}_\���s���<D��xI��GS�&d�fbfQ`&�g���N VVJ�S�w��ȓ�����Ȩ�=��������ׄ��Rn!RX'��}���ed����=���zȲ {�m�޴��u��0
�V� k���X�w�v��.�\�� ���`�ɶ�L3��6L!L?�_�~L(&����AH(������
�����Ȱ>�������"�g�=�k�C,�d�X��P����0�
���.e���[�e��>����Ad�ٓ�3����Z?�%eH(s�w�8��XjB����� dxC��G�c镹�����'������0@�Q��
��6>�A�u����?{�{GqV0#��O�ĩQ=�_Ffw���>�$*J������N2����~���
�C�v8,��"���7��W������p��s)�H[@޷���*Al`T��w��H)�
����u�f�W�j��݅b
��̨ϤN���j��z��A����4^�*'
P};��ڔqy�y�Zt��(u��4a翠@��J��D=�~���8+�r�3�	s��Jcp�0���{Aȇ%��=w�7�N�;��s���T���m�ư(ԅ�����9H4�+P�?}�C.�0+\T�t�Km�\�&�d��"	b04�MS��V��Z�F�^�ZA�.�W\7����?�����k�O����}���
��R
}���9q
���
�ﻸe��
���wx��5��0���}������2�������;�����6��p���Xb�~�m�B��/�6�/� �:�E������*Q���?}�C,�%B�%C�����q����h�����y��L�.n[�e��
������+%�+߾���H(%@ּk�<n�Yq�o9��6��k�!Ii����R�+D/}�CN���Ő���d��V�]�����U����~3��a���T��ߴ��VaX?�}�CL60�(�IDn}�P��j�y�oq�{���$x�3����8�@���k��nssqWb��X>﹨i!�HR�;����!_�c쎠m�����@m8 T��YR����4̓%B��T;���G�`ݪ�?$��`��+����݀����L�^��2���Mfˢ'uf�fɏ(k����,��k�� ��-������3f�ï�G��^[�vp��kv��@%�#cF�C�r��#��g��ܻ��.]����[�.n^�����zĘ㚵�Z,Z�ѣ�����vݷ���6|�#�қ\н�嫇����P����p]�(�pX�u�p��1iP��`�rQv���n�;��'��]��t���wu�d3��̰JOS>��`&4��ptGlric�.�Y���+��"/:�)ڮ��n��n4��)yZ�\n�''���c��L�~�;��s����8���L��{@m'+%X>����ͲXʁbT
��~�Ă�}�
����S���!�O� X�<
x#�~����>�mrNP��I������=�}�i�+9�q��~�d�g���8�����w0�¤�
������2r2�M���v�Oo�}�6��;�[������`|5�����i!K@�~�m �ߏ�DTJv��ߚثϾ iP+,K��{�i�d�T�
�{�h�+��y��&G7-�2�paS����_��|:մ�{��$�VJ����wFٶJ2�?~�}��5�Z�S��ߴ����k� ������l
��}Ɵ����s���6��=���t@�������~��9q�߶���{�e�F�����4�q�IP�����l�eH,�eOw�~�9�E���_Uot�0b�A	0Jn-�'t�g���=j�x挋��ݤH��ص}w����si�q�g��`|5��}�CI�B���w�h�
B��R
{�����q����Z����+?%ǵ�CIĕ
!��w�8Ã
����eŘ�r�S�q�L����H,���g�>q���b2$�-ݷG/g������-Q٤��x���Tf�m���cΥUQe��T��b�ҡ;O��s��z�H?��:���q�d��*=��~���+R
{߻��8r�l���w�B��n��xQg�"|�'(DdW9�3��M�3���N VQ���߻��B�*A`�s��N|s�{0�¤����h�'Y(��A�=���D�N S���b�a �L,��@m�:c�|\J�s���HP�s\�F�)
сR
S��l'
�YR���3����o5�)�?!�
!�?w��0�aXY�����L���2�l*}�s�q%���߾ѱ�d�Y�y�2g�\ۯӈ�}�}�H,HR�����i�!Z����jH)���'���FUEk���� �Pf��"'A솭���ZE��.�����sv���_����7�9r��no�m>w���ND
�2VX�S����8$�$�+
���߾�4�l*O~����מ�'bc_w�8�Y9Y(ʟ}��D�N Y����r�6�8�»���w�������{�0kv�8ew 7��2<	D�{��`q9*Q�����چ�	�<���⸁��� ^� ��г��a}��1f+������aS>���'V�~�A@�T��Mm.*!K\>���&⩓�v��a�X�>S_E v��U��\=x��'����f���mB���Pt��[:'Ʋ���kM]��3����[;�>�G� 
HR���w�Ô�JB�!~���i<	1�	�
d�bb&	`!��Mw�P�&��ϭ���p ��O��ȉ����ĕ�aXS���ۆXm�Ib%����8�~�{�L$N���s�蜉m$%��oD�a��0�[_&�A^ä�-!K@����o�HW������?8(g�����p*Q���~��C,��P�*�{�h�@��ύ�;5̑%8�B�3*�Lĥ�����9���`}<��ה�!���4�/PG������^�8�s����T�}�h8!ĕ
�YXz�����L��Ĩ�｣l3!؟�p"��i�ُhv�4�+P�?~�P˱�R�睵�c.Zb����N	=���G�H,�b�D��ُ���'+z��y|=�߾�2�q�IA
������q����YY;�o�1�x|�s�_M����D�8�M����嫗��ذ65�׻�A�t�R���{F���Z�D}}k�&rZ�?���$X 
��?~���m��RT(�����q�V~���1f+������aS>���������p�#��z��>v}^2ɰe@�P/���l��`Q�Hwn�@�j��#�.pM���t<souo
���ףp9�_�~�'�/�6`��;d�ڶ�]�Q;y?߃O̟���5N
cҮ��k�_� �����~����e�0*-��Br��(����X`�O���,� ���>�{��8�������d�
°��5��aRQ
���w��Ă��VJʞ�{���8��9է��}�_��׉c��m�;�n:�#��]'b�kvf�`�d#v�ԠW������[�N�w�q��>$)i
Z���ѾR �`T��{���p@��~������{<��w���a��~�P�AC�IP�}���a��~����L��s��a�§�߹���T+'��8��w����߹�N���{�e�̨%@���߶q�Ƥ���{���R�+��Lx��Iq�^�K��Hh��ly.T¸\��� w��z6�++%e����Ϩ_���G����}��{�ϳ�=������AI�
����}���ed���2����h�h�3�7-\��mȺ������}�ݻ����&�{��HR�7�}��!Z0+d`T������q�@��;�}�C,�0?�w�������)g�ߴq ����0���[j�p�
�׻���q �VV��tm�d����G8=����P.7�������=���@s��i
��wP�AO{y���~��k�o��xv�7�mZΤ����2�`�`�9�K5.�;��e4��F��yx.W���|���Cȉ}�_X}��Zo��.��K��=�b�R�~ΚLz\�xѾ}�ϒf��rZ�R�-�H��GP���!Ow(��+&���tϻ���Wsp��ޞ�uM��>�I�U��M����4#\�:�K�=u��M���^�bl䐋�1�tG���B�r۩��דeK�Q�vV����Y;O	��D�aE&�n]m!��x܌��heeL�D�ab㻭�V-�[��vT�v�;�os����֯dQ�\߸�>\��l=�6�&���D��g�`yb��o�(�͵����A��a��~��X�Bq*���3�ooq:���hh-��G�M�s#pE�w�}Z���/�bI^9xNu��oWwD;�ϥ<��5R�d�2��N%�997�|k۷N��L}��Or����Q�ï��>�ӣ��Rښ��1^-���ݱ�<�Td���ʍ�)���������pA�;Ư@��vQ��4 T�l�\�.�;j΍��w��+��C��>*y־�r�Of�P�mM��3 ��q�����i�O3IE�5k����r��Sԉ�py��"q������Xb������C�l�2��{.�8�/&+mw��#,����t�I0�h�����[��ײ����]��ą���V��귤�ss��Rs��]ZE��4�.�$�Ժ�y�cG	aԏ�Æ�#�w�f�c8�WmQ`��ÆU��DKE�V#TU��#G�*R�b�,A`��UQc�l�b"�T�D�*UX�QX�����-PV0p��#+*��b1�����S "�#mdb�X�K���2	R��QF"��`�ee�b��*��mX[i�\R��#�AŠ��#DV��VmF���Va*�*��e�-J¦TQE�H��(����QU(������m��(��	*�SJ*�QE�
��
+i`�3,*�lUb2�j�E��((��E�kAXU)*�D-ieJV�`��(�K
��AUe���Q���Z�TE�(��ETbJ�PE��*­iQb�m(���V-TQ`�V�X�ckp��eb�[UU�J�ێ�߯�?+�\�nט�I�J�k�Qt�Ÿ�'m�����v�2s���̀�ۓ�|�g��˶Dz;\�j�q�c�ɺ�1I�q����>^ȴ=��熐�-��Ƈ��-���#ٴ��9n���ҝ���s�5sK۫V�s�Ǝ��2�6;+�O8��[܇BOV��v7Is�įe����n����٧ñcq�F�۪�$t���9]v�9���������l�3���n	A���Ǵ���6�q�v���G��w�'ѻ_[�Muv9���͹��y��Ƭ㛅١�ԻN�n�ݱ�Eۧ�GIv�u�(u3��4vW��� d{�mi��e��V�vWs�'i�n7:.��c �6���<����۟;���b��^��&i�Mہ�l��x���5�]���Z����t���u���7}>���S�.պz8�W3t��أ���6��@��ayө��|�;w=��3��V�x�OE���y���g8�Ř�cx��݂��s�����+�[S	M��]q��Ǳq�ayö9z뛶8�����ҹ��9��<��:�^s�9D�n�֜ub�Ń�n�ts�����;�6�ļ<��73S�ʌ/n3ʹv��{=�p��=�mu��9}�Ͼ�7IúS�s�:��\ksڮې�V��'�
���
��';�a]���ny��(�{\x8`�Ac�]�{��ۘ��y[��͙���=j��k�ͣM�ޚ�{��͎�۸������$z�k�cZ�e�;{#.�q�t���7/�Y\p�[��s����g�oq{#g�C-���g���n[��zʏ�n6����i�ˣ�F�n\Ӆ��c�[P�����h�����p�]��ݹ�ۭ�j�z�e��Sex��8�/\��BKG��>�:�`d]��'cO=�vݧ�{r�3�:��pT��M�q�Ǎ��Nc	[vÅ��^헷[(��P�n�Jr�������Ag;���(����p7.j��ow����o���9n觬ݓ���ر�6�J�����yx����օ����K��M���W2vY�Ӑ�m�]��ze7a��,�b�l��v<�p�;�y���`Y0�n�J硍��m�ȹխ��lK��#�j5�]f�8��n�7W�<Wc�)����[s�s�*NT�q�KC�k��:�^M���kv^��7WF�J����O��g5�gj������燵n��`C�6����2r^�i1��������.r�qs�� a?�I�{�h�p+(�Yc%N�����'
°�b���'��G�np}:݁dח�}<��FVJ2�����@�G�~�1�ܘ���H,-ƻ��t���~\���ߜw���1߾�����������N,@�;y�u�c�"#ȁKM_��ɟ�$Gӳu�[��g�?0�
���ba�3�p�AOc^ރ��X�d��=}�C) `�@���6+r�k�|����i������� �B�{���v0CB��Xd�S��I�I[V��?���8gZy�}����d������sGq
$�����w$��i���h�'������k�u �`eL�_sD�q��u�)�.3�r.Ł��w��lv������F�)
�����@��S��O�*Q�����P�6�
��P�}ߴq�V��}�~��qg��2\M����{7Sm=l�2�\�8E�k�[�kѻb���������Հ�>��*g�w�8����V�w�7�J2�Q*{��Ѷ ��1O�!���w�G�y!��� /և�A|f�xQ�7+�`)��8]��ؓ>��h�AgJ�k�MϾ�N࿟��DnX3��&��X�'!�z�E@{U"Uvرt)�eĥ\zs�e,.����C�.�����h��?� ߊThM���9k�[�!!?��k���?�T�����a��IP�,N���h�'T�ɼ~����o�)���z'�8�F�=�LD��BQ`�dx��WP
B�����h�Ax0+X7�}�L�@���d;�f����i "<	��l*%B�w���8Ì+
s��˘�qL��2�l*}����=��k���ÿ�$��d��������M��*����`q�!m=��� w�������"+�	#��[�5q*D�PLJ�� ���2;� �`�R
~�{���x�1�������&�pV�׵��
��RQ>�~��$����=���������b������B�I0���pD@�L�H$�n�K�n%uֶj.ٹ� Wo�����ڎzJH_�������C) �w����HV�+X)���l$s�~ް��\g���4̧����c%Bĕ
����>|�Cy�%`��JI�r0��{�h8!Ė!Y.����|:_n,Yc|υ)��3�#��!f�m ��Ow��@p� �HW���h��� Q��xI� �C>��9��Ip����M�3����$q����>�}�q ��°�����-������w���2DM����Zl�mFF�S��B�9�!�=��XBи�2m�Lٰ*�qY���8Q9xEF��H�w/gw��X�5�Bs���e��
��T�O����H,�Y+*{��������eL��BQ`�g�qG���+��3���;ޤ2ZB���_���+X�������*eOc�ݯ	>�Yy�}�k�����+��" ��Ã
���.ba�3�p��=���!ĔB���O����;��uIP.u��gk�!e�}�{@s��i
�=��wP˶NE�L�ݴ��!��"��(���!z�0�����鰻�v�C��Y��U�!pv/b��$�w���~1u��q��|��繣��
��Yc%O����ĜB�+
°��ﻸe ������O��z
M����h�'Y(2������q��w�)�9��.c����z���������t�7�51< w��>C�|+��"��݁���R�VT�?}�C,�%B�D	�G~��5�}N~g7(a���>�~ż&.n[U���aS>���pC�,B�X2�������2Q��P3��}��ɟ\�����H)
Z}�������=��wP˱�Q���0�

�(�"7��{��Q�aF}��n��$�ȢA�}����ث������� &K��a�EUVl
5:�`��2'gj̣����@Ԃ���9��W���=��k������x��ç���{�|H9=z��A�vʙEH�P"`�F'jA:��D�Tetk8�tL��'K������ߛ�%���������~�s��v�@�Z+��k��u�[�s#�u����k�v��o��;|���s���p9��|	<o���	�Ǜ���N&�FG�e�lG'����\ʑ0���<߳{du�>�,�u���H��"� ��7� �.�hD�_Vg.��D�
H��eO�s���S$��Ǥ�v��ܛo̏6���꧛w ��!J��&)�cw8q\�n�3;L�9UI>o7� �w1��L���ߝ
����أ�<bf�"!2�U���l�H=����Z�EVf⩇�	Jy�x�w�LI�����Y;fj�vE�0���;��~[o�l]�S҅��:���$�<F�K3���`��,��Ĵk��L���&�T:n�Z�38:j�7��=���~0��z�Շn!3l�VCn��=�#��nŞf���ݦ�v���`ݵc��ǫ������2L��9�����5���ώ]�v�5�l7Z77*���W���9��3
g�:]�q��X2�	�n
�<S.{>[+�.ȕ��c����v�l��Fu�{6��ͳ���^1��f"�.�c�O�������9ݾ�3���I��<;���Qq]�e��$�<:�.s�B>�<v���
޳�Ż3�F�ݤ�������F.Q0���I���i�N�>�F\7���B�'w� �6�?0�A�H��Xߙ��n��9��ӕ���}�>$��y�|I����2Ⱦ�f*5�nD���ј�XP:�[����'���0�v,n�1�n:�P&�e
 ����
z
sBI��E��{�C�bVO�zj���}���?��#�����.�D<���#:͢�bLJ�I��c�9�A>:o2����hF<���$MO6� ��`0I��+��	������c���E��n�:VN8Z:�������&��B&K�Uҗ������N�5�c������Nv^�2H:]�Q��&N�X�m�Ff_V��W1&B��L­�C}�����֋���}9k�ع闻q>Uuvc%,lZ��J���=�SP�t2��x�u	}�<8O7�Ȩ4$?`�r,"m���rv�|>'��|�$�w�P���Sjw=%�'Y2	��(Ս�H:]�IY؈f^�cq�q ��~`��N�
�髙P�������o����{X�4��L=�lI�}4H'��yˇj�Eҏ(dl���9b%�RBf&Lx�#�����z�<�C����Lpؚ|�$���k�c����T�ۥ�34�)�0?@��%St˶˛�@h��T�6݋�n�^{hǐ"I�>?#��0&&!a�vs9�H#]�� �1�s�M�d�[̣�{rp��`?u����L#0Q�d�%W�f�a�ݟ��ܪOS�]Տ� G?/�1�s��9��]��QO���Y1&B� Lʧ�mE�;i�@=ޓ����y=GC�kK�3�����Y���h�ws�[�9�x�\�$�ׁv�.�����V�[��3|Y\̣�/�xI�c���QO]��hX���}����~=��&Td@�������}�v�g:�D���$�u�s`�H9��{sc��>�G����Gp�t	k�y�&�i�ge}L���a2a󇗐�߹�kd�ss��J�)��4M�뭳���
�g�I�mŶ��jݡ�=�O��ˡ[�v�ZD��d��幰С�2ϛZ�s�7��� ��e3O�OF�����v�$��w0�,�,$l�om0IQ��v�fGE�a�w$�u�m2I9����skk�忍�_�g�<w�����"�#9����l�YVk���	'���� �ss�����&D�� L�`��M���WU�f���{���{���u;蕚`q����`.����:����GZ=��wrl�L�ۆ�R��k2�n�&lCd��]���iOH�Y��j������ �����?:$m��2��L�m�u�<pT���Q�����l�A����'�U_G�{��Y�ݻ�L7�jIm#�ٱ��F�n@��#1#ڙ��ת问�s۰���߻�ɕJP����EklA>=��LN�}ܣ���D��6��~$�gk���RBR�'č9=��s�;u�eGc�ē���oă��E��U�;}�O���X"!�0H0ߎ����:^���W����d0�[�.���M����Ex�����f
"� ����^TXk�$��l-;�O���v��5�g�ؓ��gg���Ϣ LJlcj��Iܾ����Vɂ�3�������w�@��{͜��=y�E��&��#Al���/19׽����>���N[���L�^r����e���x�:y���LKZnpO��}�~���? ��z���)n�nx��W=��v�nx�ǷOY�Z��m�C�s����A�l�[t<�N;b��&z�7�ֵ齹�sН�U{�:��?^��u����<��@u���yջc�Y-����x��ۑݱ�\݀#��`���m\uv^]�y3�[i����3���Q�2:��;m�=�ۃ%v��7<���ۋ��8�ؖ��5�ůl�m�e��E�kz5xy�2XZz��r�ګ;n�pG1���{Z����d�A������v҄(3 ��+k[d��}RA ��{͒`���~0�_k�����^���JP��ob��V�7�V���כ�W��I>��
'2��$�]���3'fb����	�%$!	(�|Mx���H��Φ	�jf�_@Uf`�`�m;�Ne�6	��,��o�ks�+l��A�w�@��y�� ���tE�M%�O�udQ7u�*!��I�U�|�$������fD[�S#2rz+�wy��A>9��څi�������
�T�6�ĝ<v,n6|utG5������`�m�FR6�ݩ��}w����`��bV�(�UI$�_m0H$�f�s`���º-�������[��hb`�(B�0
���� �N��0#)L1{n�==Qe����؀�`MH짍Iټ�艻���;��I;��<}�}�ܓc��α��$�3omf�{k� i���A9׼��ͼ��|J9Z�nJk�D��kٔ�eHR�#f�m��N��??Ms����t��p'����oĂAͼ�b)R2B��'��N>]ײ�(���^�2A ��ỳI:��C쩃�pU���#3w�cy�E�"���I�������w�%��S*�����I��$�N�(�9j˘Er��L3���ݒ�	ծόWWU��&�ӷ�a�מvױi��u�D���q���Kr��7+���:�X`�@��j�VC���)m޸��MooD�_A�r��Ir�tbX7u]
�����$�E��l�F�}	�g뭙�Uzb�̽ �3����
�(ʫ�>#K��$��_=����LL�������<]/��P9ᯪ�f<1nU��#�kt��tH�}��"�pqq����<q���Zd����_��xd�EW���q��l��^.M7z�x�ȪfB��ݤ���${)|����[J�Z�_F��MV��o%iY�W���^�bǉ>��no�8u�
/v.���jw6����f��^���'�Ç|x��{)�{�w�1$g�]y��v�D��s���ˡ<=��bwXcn���6i5x6&������1�ijU��ۄЅՏ�d!�5�F�Q�<�ܱy��pa15��)O�B��jE�q��/v+Mr��zI���|�@M�l�T��°΁�|kޛ�0�&��4�./]� ٛ�q�tr�d��{w��@�n�t:8�_N����T*�1whq͒��:�]=�Y�oz3���/AT�f��@�j�)�e�Ь�{,��.��Ef�k��;�����ˋ��i��r�����&�xzOL��'�a�djg���ޓ�wW/Ofh�aWw*�O!�r5���R\>kq�^�@7��o�Qe�`�%BȽ�&�����2�X��oʌU׸�.�fpea��$~jv�|:���J���>k����~�!=��%{}ڨ����yn���L�iC|o���F��/m�k��ew�T�c�<�<�C�ʖ5|x"����/��U8��*<�I��)�����Y���877h���y�]uٞl�Av�TX��1�QDQE,DjR"��QKj,DDUQ��B�ʖ*�
�*����KeAb�İE��(
+�*�[JV��`��X�*���`�ja+m�J����Z���j+[0µ��0�cTb��DD�����UK��qj%j+E-�T-+�\2Q��1Y��,�!V�+�YP�-���J��[)Z(�E�J1��mQA��
�`�FVVE�AE	dcR1siR����*9�S�ƴPUT�TF.Z�1Ū��QQPETXf�	���{»7,|	����K��P�Na�u�M�-��mn)��k�;G��m�d�.�}ow�gq4��-��M�;`3��TJ��'��:q�I$w�@����L1�@�n�`�w�@�����p��r���9yh���S&b����乧]v���u�wa9d��2ѻa����(*b&&,l��IK��$�q��`�Ýݛ��35�	#��z�MDD��I�UFV�`�Fb;�E��̓"��� ˾��q��d�������g�2�lD�"H��1)�B���5��I�S��.e�*뺲�$�}4	8�z��dv�		B�P錪Ǵ:��$]�U	������|f5Bd@ގ"����bv��dcw-�M��F� �k��v;2�#\#����T�&2rۏ��(|O���4MqW31!Q�7��$�]���hEFd[bIb�h��{�� ��_?4(���v҂���	L�g^�ɟW�D�M�;]IC��9�T�f�E�Wo͞��3e1[��Y�����|���EW���x4^t9.�It��sD7}�7�h��(��XV�S0�e��ms���O����$����+cʚ��GM|����A�K�$	W�g>l/���I)yP�b��jީ�|O�ou����LZ1D�"H��1)�����g�p�D��/��$t�0I>$}�� ��1=�神Vk��9�a�ʰI�"�VL������ �<�!BdN������u��8�F?S��[���L.W��&��}I�8�}(�oq�%ϻ�<��=i���,�*���B:��&V�v��u����w���7~cq�6]8�m���G���B�3��C=˺�����}?U�����m����l��0�n�i&��`��5v����cc�E�xz5�.rZ��Y4&c�& ��{g�T��=z�b�=�*�����	Y��]��e�)��ú�'XͰ��[,mmH���v�\c$�Lsv��8g����/Wn
������d��ۂ�m�⋆�!ՙ2�7G�s��3px'�7uۭ�r;�=��/��Н�{kI~|����S>Bb
30�{b��I ������
O�M9\����o � 9o�1{"5�0R�(��n>�^P�5np����c����$�y���A��h晬ʉ�w;*�}���^�%LJc'_P�F��(�|s�˝8=pXs�Z4��a����׉}CjTA�K�$	W�u�6+g$Mr���v��~'٢I���]��#j�4�$��l��ъ$�DD	�M��*�w/��8�Jd�_V�~$t]6�$[y"�>̽��9��F�"��
&AA

T8�$���t-���n���s����]��e�>�����B�b�(E�W2	#���e�6�Tf���nq��ޏ1�o��3������YY��!_6�d���M�Q�wڴ7ڨU���\N�&��p`�RV_}��<�z1��!��L���º�.v�4
O;\��#��*:��E�|�$�����$3/�a�ua۳�:��'1<ڃs�����@�)B�|M3W����P`�GdF�Gb�Y]=ۀ	9o�W�e�S'qU�5�a6ʯ���Lx�����~"�nhOe�S �㷽�LGUMHb�<�Ms�mJ�2az�E*7_6$���n����y���)N9��y���&ϣ�_*�$�O�-xO���:�ZN�(���<v��[�l\[K�x#�{id��9D�"H��1+;�(ʪ�_my�6����/L�c0U�
���O�;��ߋ#�1&� Ē�ǪkX�"3�z��X�ڡD�Ge��	$��k��[�|3IU�\�t�O��LGRq�fa����$�w���B�7���1S�'��9��+VS�ҵ�n���t2��ί7˯\����m��I�x�U7&����������'yXgR�����z����۟� ���l	o~�yA�s(%(R���F��Y���ѱdo��2I ��m3���DEF<I"c;��o�U� Ʉ�*����T�m5��[���n�	�x�~$������t���S��z�,���ɑ� ���v(ݵ�eht֛�ΠNqd;�{N�%֪�DK�Ң�^�"Ie��A{��$���B��{����וb�m�H#�;Xz:tj�(D�bU0B����cu���p�s��/�['�m���)ÎuS"۞�V���R��QH� v���O��}THט흗|��^v�?��(S3��L�FR�f����O��2^>$�U�t��d���g�޴:��-(R����g*��F�˺t�dq��jp�\o8$�gd�y�$�2v�xwN�7rc/��-62&1���3��Q+�<��_?��:�2�P2�B�>&��W���oo>���ocI���a�A�{5�A#.����`���'�hi��D	6�d�J)T�۞�&�4T%�����7n��=�W\�������� ��S ���/;$�����D9w��=�{+��� ��6$������b�^�"J�u�`�q��Vwmo2	'�-��$���2A�}�љ��E���u�+��5��Z�c]�p�v�$��\P�EB}Uu��u�H��}�hw$B��B�0U z*���"{�n؂H�ܡD�soy�	#7;{���)Nv3��|D�\�5�u���D�P ��cb�� ��a֯-�1\��>*��|H��� ���m�xb'.DV��&�(�,��h�獣�<[ٜ'p\�m{�O�����Ǩ^}=�52*~ml���7�����8ﶻ�׽e�TW��Ҋ"��Fd�f$��A�����k����ʙm�v�.mv�p�����5ۮ��'nܚ�獦%v�st����&!9H盈� M��1����j:(��E��
l5��\m��&�/cX�'#ΛG����]��9B,Gn��z|NwX5�/j<�X��&N����h|�4���H��zݹ��<�i,�j��*O^D�l��2��&�(�m�Û3m/nx{x�x��i�{��N�x:3�p�ܻ���s݋����W�&��ӛ^�I���d�I����e�)�A���kĂF���O��(�2T� ��ov0�[un�us[4(�s/:��>9��A�/W���Zy��D�D���S��R��%��ݮ�I��}��� ���P�9r�3���$��u�	;�[>�գTIB$�%Jl��Q	Yx��d��}L�����H���&�H��L??N��47��!IP!B�*�zg0IW�QWA����jh5��I�7�z���W�@�a��J�������;�C�۷=mK67=�n����dYn��(9�t�t͂;{_}����u1ۑ�TWeN�� �oz�������U���D��@׶&.��I���yBLÐ}%A���h����shӆ5�{��}{�f���$[t'��MA�Z#c����Xܘ1�Z����wwggon�O��])���5���ɚّ1f�`V�N��'67_}jg���״�$m_�@�]�C<��M��v���,Yh �$��AM�޾��ڼ���.6+��s5��I����ھ�9��*�^��If�U��#:h����筲 ��y5�K��h�%lH�+�Gx���l��Ѫ$�B��?����_m?�^sV2+F�$]k��$���.ﹿ{�ҫ{{�f~�a��57$9��C�n�<��#�����3���U�W�S��~|�-���]8����������|O���fN!��k��@1�
�m�n{ ��{4��DLJ
�-�{�o0��M�@�����Nl��w�D�Hw}͒MJ��c���\��:�ʇ �
���9�D�{y�$��do9����WE�,��f�H�;��p��fIP��W��n�{L�#�{J�k�9�w�N��y[�F�9����횚S�5���n���w�^'Ʈ��I��)�t!Ȅ�)��ǽp�LF��m�AӕD�w{�?of�Q$fc0�	$o��;��I�azdBI*���2A����:�I{�U�
�)�M��{��I'7�Xīw]�����ߔ�X�=Ls���;0Ls[q�n5����ȶ����3A���ϝ�lsn�V��Oz���L�I9���`�N�,�2}^۽��!��\��Q`��6�&�U���V!L�x�E�g6O�7� �-χVb�,�r�33Q� �ao#�l	7���d�<ɒ颔vk��,�@����#7�khDDT��T�>&�9�+�9[�q�� ��ΦI$�nmRm��}"՝�U6��G�������_���������4�>�Io��]|�t�#(^�f.�N�=2��¼F�qp'E���ok��ܢl�QTA$�`���0O��y@W,�7֚��{�����d���F*(M�QPG��7�mX��CQ��5�Ό�v`ݒ�mu���Wk=�� ȑ�y���)r}$���7��M������$��}"F����g]^YUU5\A�����uh�P�!D	�T�B��NWC�q�K��)��O�@ ���|�H;w�@��cw���.r�օ�rD������N�d�6黎���1/�luL͉Ŷ��$�������j-?Hi#sBZ����v����٢�v0�$��A!��1�%,̄v�]�@$���킦"��>&�#����{y�%�L@u�=�8:��$���|Hw}̀o����#-h���0Z�^�^�,eg�s�r�*��,�J2v,6!>T��o�����W]�� &Qܙl��/�G'f������*�.�~)[ �ޛ{}���L�3	��:��yq���|��)n������f��z1���q�׳%�ܼ9G�N*R��Ul�)@V*���L�t�e�����o��ʪ&�Q���Q$��=p'к�-����$��{kg;�uՀ�Lr�I���i�*e���*��v�_bh��)�]Ou�C�K�E9��q��5N�eV�Y���9m�7������^�^Cr��$��;�z\Pw/x�mXwg2��[��p�`Ǯ�9U:�t���7���w��$K��,_i�P�:6���g�;�B�X�W$�;1#:��� �<����.X;+ed��zLK÷h���Uիs���'&��Wb/�����TGk�R�3��z2a���XY��.r�\C�p��s�)���"��hVn�z��:|��1&M�j��a���:�f�"8���sƟI�q;�����{��#�v�$�=����7�!�o{t�+޾����z#�&�D��g�_��//WW�}j�NR������' 6U �>�X��Z�]W�=�8/3��E��}^��b���1ҵ��OGZ�b»���+�q�k��t�8yE콡5�塇브sۜb� ڵ@k�ӑ�����2	�>X��<�Y���������nh�f <T���KdH>0�3�ǂ��nwn�&���f��<�BD��c,z�D��+��.m����
,QC�lQETQ�DELZ����	�0�a���dEb"�(1TE"��
(,`�AV"��T�6��2	�U��S�TkTV1Q��mD���`��X�ł� ���J�*�iD"�"1U�,6,E"�"*�b�آ��2 �S˜(�����"�Eb���EH�EG)EA�ň�C	UXV��Q��(�UUL��m�p�`��bDb�V�E��AY�EV1�PEb1��QA���m�;o'�=�oϭ���ʾ���S[�����gm�7;۩{"&���r(� ��W�����ɑ"gt�&�d��0^c�+�w��f65���$j-H=�C��Ä-�X��ێ�m�q��f���v�2lZMq�n�1��:�/l����^�\۞���j�n]�ػ1�Em��i��g�{v�O.���[���w�*�ņccNǳ�&�m�X��sۉ�C�#�76ݔ��7	�Ԝ����:z3�C�Yg����pg� &k��ٍN��r��$����i왮U݅I_��o���N������e�絻�s{��n~��ŷv�:�tjϞ���lv9���q��%��۵�d국�KNxt��.�l\���g���N�W�B�$����6���\�yu�����/9248�K���m��{����K�u^Ӯ�e�+�G�nn|���+��yj�f�7�lY��\v1Q�k&���k�7���9�}6���vؚ�r�qu����[��J��3��������'n3�[Y����;4����8�����*�Uɸme#[��eԼf3���:ٌK<A����;�6�.�Cq�g>�H踧�c�$��9�!y���&Q����Fx��E����F���/�b�Ka�3e���Q�w1�v�I��9�l�����d�;e��� tc��L񕱷=qt���<Pk�cѶ���v�b�qg���g����niԻr��Cn^{�C���q�q���{3�G!��un���E���=���X޵�!����O��}�n��[[�t�ot�l�<.��v}�l�<�X��=M�7X�.������ݒ�ŷg��cV^�m�e:uV�-v��8�8ڇAǣ&.�F^s͏9�N���d��۬���S�uںi�b�Ů]��u�=ǵ�mNn�9���Ʊl9P�|r�m�<��`���r�V��{���L��72�s��=�U���Y��3�1"j�uF���F�:�:��+���'����ӻ�;K�y����^d㊷=����tf�GG���g���q�h.��!�7c@C�btz[pb�z.t�k�x�ػy,���c�Zѻp4g���+�n}�cϺ�f��]�����p�u-�=���Ȅ�n}�<�4mՃ�C]cO!�7n�����Mv�j�f��>�;u:x��n����㶎��rO\7)�ks���82��^1q^�������{���2WG��I��&+���o����]ۏ����_6A$m�U|	ﹳ��t����[�5&�;[��׉��0L��+Ҥ"�[�Հ�w]n��sU��O�|H'�.�E��oě��N��j�w��f�ë8(��
`L�l�;UD��}� �\r5�O��0�٠Aﺩ�YΔ��n�X���uS�γ���*��ć��� ������]lbgc8���^���3�"�ВCI ���;T0oo���gf�ڡW6�T�M	w��������qmneM����,ѣ5"�iX��i����j�6I�]n��������ɫ���oߏ�ۍŚ��2�hQ �}}���5�k2�973�X!�Kv�u2w6m"TD�En��|ê�,���)�@���&5�T��WudT�9�����/��5iA�T�m��+-��1&��9[U��;|��M�dzno�Iy}��A'^������*�K�r�\��]C��	2��"
J��m��O=�l�U�z�Q#i�r4�}�2A׽����T�@�	�T�
v��͙�{�q"�r��{�A����v{�����f�u�Ƅ�1 �1d��W�Im��U�u���9�F�����B�wF��m��-F:ه]�=]i�*a��1&�K��ն�'ݵ�݇vs�ݳ�/RZ�cJtg����ޭ؉�2e#0D�>��ֶ	^��d�}#��#��n��z�>"����TA�*f��t�u	��ʫ��]wt�>$�^<��ӄ�؃�R�TdWf����K%Ch�q�}_SM�F�������̾,Th�O�٬�b;���j&�9̭ysk��\�t���3�T��V3��`䝪Bk��t4��0fS;;���w׭�	m��ghh��"P��AITf�����F� �n+r� �z�� I8�y����+`�Ob]����}�B)�n%���^�3����������^$+�m�	�}48�|�f��Z7Qv`��*��ʬ�A������JF��MC����t��t\��9������?��*bA�b�\ʝo���:�W�{wS�[��Dk�֡L_e���@�Έ�|��!hĵ�r�̀��z�b2��0|	;o��$��7�$3�ɮ�}Z:��O����/DfV�H��Sq� ������.�H��ʾ��ܷb�	d�m_8��K�����;c�Q �N>�oĒv���|˹���[2�,����S��t�g�|�ʘ�s3WܾZ��szVc���Ly(4�����7��)ON����.��܂x�3� qp��g�J$ɘ�O�B3z���׻�ϣ��{�߉=v�P$s���$��T�	_������d���{��u���^���+�4��f���(%�s0�Uyȉ���`�L)ʪ$��3�2I����Z����� �����}Լ�.�0LJp8�2����c&p^�ҫH��T|O���� ��cٙ�F��:k�2�fbL�f��ى��<H7��� �X���Ϧku�x��;��H;��LU�
��)	���^#r��*q�\R�$��n��������Hn�H�9dm���n�����b�	d�m�޿kmm�K��{Cu �]Uh��wX`�{3���۾�1f���̎���B��dҝG�}��)�@��yh`*�g����6��q�����X�k���=�g��af a!hԉ(���V�Hi8�kذ<h4���msx��q�����.�r��0�7�0w*Am����9m��2�i1�nMݱ.����_JQ�cuv�<W�h��iݗ\Q��P�5��/��9����6���v���m��[��w6�IK���vz��k^�lhv�-՟5���]u��3��2ޜ�a�Ѱ7cmO%9nn��q�,�>N�.��I.&k6�p@n����jws��������:�0��O5�H=��L�N���5US�����U�����l���D��1fd)ښ3z]��}5�yt8��ܦ'n�h�/D�T9���X>kI�
bD$��T�V0�#n��FUR���5��;$����F���$S�鉁2Q�"f�OQ�U�$��>$��׈#�;7WP��%�,�Aλ��d§�J"ff#��#����-�m0fR{[+������7�H���w����m����c�e������1м.N�����I�3�LT��S=�WN}�����ÿ�YH�Ba]������Qw�ߌ��;臑�$� z����H9w�@�/�����Q�LQ���$�E�I(����|��}.�s�i��� �_i�b����)�o�0Ҋ��v-��pj�l����L�%�h��R����
���P�.�f�o*���Nn��Wnmu�g�.Q�ȉ�A�0�(��H ���g�ݩ��3gkpp'���E�w��-a=BaLH���09L��Y�k��I�uG�s�����죸k6�pވYȌ$�[�^��ɉ�2Q�2f浰	��쭚�rH.+��$o;Xd���c}���s�ɷE��0��Kj\�BpԆ#v:9�i��Kk�m���8Vu�ز�g�-_?v�?~wn7L��x��#����H6���#ĂF�v6s(Q�;�gV���(x�����,�0����U|�w�ԜW^w���eD��y��׽͒	�����2���P4+�gj.j�V�ܞ'r+	��0�3$BK7�$���0G{'5t,6���"�ylL�w��xG�,Kv�])����5�QUI�S2A�z����BQ�a�����)��<2�>��I��q$���6	n�e=��D��1&�S&��P$���0Ingc`�pzO���:��?��޾l��^CB���"(�Ue?۾�@֝�7oF�H�v�$�ws��$���~���}��0��m���ճ�	�*ݵ�sY�����n�v�����7���������͍:3�浲A ��	#n�h�wP�Ν���̀������[ #Kt`ܞ�G�y9�
�9{5t��ge	;w ��嗣/�Lcnٴ-����o^��Iw�@�U�&3^����$s���$��E�V�1a)D��Y��{�B����bG�T���`�U�����yT^��+���T��������~���E E�~{s4}��H�\Ok�س6D^Ι����Y[��y�Wy��m(���{;�sΞ��%D�@���cf�	gS����ko`\j�2ri�d�|r女 �w6H�8އQ���X�!��ήg1�l�P v�r��3ֻ�n�K��86y�`)�D�J���b`��DH����ôH۾�GĂ�wS��QV	��)��˖y����~\u�l���ZZ�湰H���5�iG��}Z	��ɢ|Ho;��$x�'og��ͽ��*h�J"ff �k�vVТ	 ���d���U9�d�t]�H$��� H%��{��V2 r�T6?S7��Y>��t��'g�#���7z��ޚ���=54H�XI10DB��o�ݽ�s<+�5��	&�w6I ���k{�t�Ɛ���-�1�0h��H�|Uas3OgV��ni)��+1��&7#�pJ=�Y+\����~�{�`�k��줝���ў��*v6�t�1¦]s9��<6�9��H�ct������]�m�]S�l=u>u�{����\�x�hS����u]NΈ8�3uvz�˪yn��k�2��.�gH:特��^v�-t�ϰ�ڼ:�\���q��;�zv�tv{#�lM���mg�S�k�:C�h���8�����Ӗ�vC����,�帬��ױ�+!8�݅,��۝wb���kS�T�;v�V8���������;|cfxA��� �F�^�
R�i��G���$�7[%�'������"(ʰ��+FN�N<j#�TˠA!��l	;�z�>7��Q�qZp�錛$V�+��3�1(D7�sͿ	��[$���v"��w9�A#^�0�#w�XdP�
Y�DL�A�r{c��,)��bkٗ7\>'�7�i���}:����c�{pOu|�	`�t�5f�C`�|�dm�UNj&#2��Y�� ����`��}4U�#9��������OB�3��^�Q���Fg'���اQ`�um����q�3�S�%�%��j 譮�D{v��$�}4umH��V�*�����m���TJ ��-��j�
ٱ;�E�k�hr��vH#�	6��颜�ӏ�g��{אm�m�=HA�]G������ّr1��Jr�nbn��#��[$��}"�̬}7�Pp�ԕ�`Ƹ�� �LT�1^=��	#n�h�z���܈��fj������H��2uX�>S2�'�U	]*�Px�=u͟	��{4I6�y�
[�����Q�3-L�����|�T$�"fb&���H6�:������l[d�/��$�w�^'��sߞm�f�߸l�`GZ�aX�c惂v�l\b{<\�Wsü2���Loe�+���|;QQɉJ9��we24�ʒ	�6ﹲ�Cx��
��A��N�(��T0T���U��� ��[[�oZ��|2.��`�{�<+�_�o~䛡�`'*�]
$4�]dHg����| (a���Sl�N��A���4��P�Ol�j��4��ҵqv���eR����c�A֡��Z�o�&D�w�kN_$��aHGvy���jw^���\<���gl�y�� ��jE<���n�}{���
�b��!h�M�k�)r���G����f}�;:���{��C�Z���ۣT�a��/�ֺ�]@�>\͐o*�課�P�^�XA�BT�,.��ފ�{�}��nlO���՗�L>^���5�tD��zq�p�ʒ�l���(�X�Gj����ͳJ�U�)ټO
�dŚXLQ��b��Z'�f�G0�{TMFf�S)!�˷����){��I��x]�������G�K/�}�~���K�������xEĔXH�啯s����8��`�"u��R�����(֔+�U<s]�^ΙV�
\M�[;�h����(���_)���8��yoRwCBhԬ�l�ՅmRJ�+����(�r�aʡ�ak3�r�
פ��E��û9�Ѽ�]��\L"�����&Q�$�=��(����X
<^��{n�R��l�����K�����w�QKP�������J�^�/b����#@��X���fi;�pnƀ������7�6�8řwd��\]A.��ѱ���=��R��,^�8�G�^�;�o�Vd�&z/O]�p(�N�{�E~�����؀@b�������ؗ���y'n���U1{�����=���_���҂*��b���"~mJ�TX�"��*(��DF����EXa��0U�"��X�J������QF*�U��H��Q1k0�U��X�UF$TU�m
 ��TAV�VSZ*"�J���iUAZ�%�*�PciH���"�Yp��"��X�#V�b�UZ+U"�*�*"����Cc!hV�Uqj*8�07�a��[��EU�cQkQ����m
5�Ub�a�.-e�b*���EEDQb��R��Ae��Ҹ�Q���1DUV"����֪�#���Uc�a0�(������Dc�V*�f-�AUa�qkKb��0.[h�+�DdQ0�ƭ�Y�Z�D�Y޼#�wj����Tc}�I��q2�����DKr#*g�I<kj��A����>9��p��L�Ʒ��Hjw��l�9pbϯ3,lq6�B�w�6�:*](����H���D�F��6	'�7�Xu=�$������Ko�@y��f۶v��S]N�i��Z��拌�4�H���."e>Z��ɦ5$����jA��I9���Ӭ)�G#�����`��͠�QɉJ-���lWu�ͮF3��bI$���a�s{u����ZEe�(��/Ď��)D�%H1!��k� ��ݠ��mڝ1{��>���� �s{u�Έ��%D�@���Fv��f��$��t�����l�N�}v���5Y�/2�5�w.�	|"�u��oJ��dr�ם" x�'W��W�2z�w���sְ��C�F*�1�u.��W��8|�Js��^������QՀn�Rb�WMk�>$.�(Ƶ��d7� ��0�ۺ��F�}ny��oK��G��2�yޛ���]��#�k�c��Q�흇�,#�L
Qr�	�o�t
g�fErح�����`3�@:]�}{���a��w�u��T �"L�@&����"]���d�ud�A���jw�@�&$1�'����bn6m�;��D*$AH7�����(I'ǲ�9����H$���y�N�gF�J%zT���F�[���u��H,S+A%_sl�N�yI"���U0d�+2�ơsϼI[��Bע"J�>1&h(��zA9��L���⽸�����A��Q>$]��gFh]�j�-��[1�N�6P��'�N���N��'|A铗����L^<\�ط�T��tm���k��+{�A�N�1}���wF���A>	��a���W\�f��ɫg�Ho`K�4p�s�%��ۭ�]�SsnMi(�r&��r��oC�Y]X��5ݔ�hs�vm���]�qŪNs��c��[�<�Ɗy���{�h-����Q�[��F�1�&˜&ն�e`L��&� 81=�Ʌ
ջ���۹���v�#�io�����y�kc�M%��{U����f-m��؝CK�q֮[W�6��@�зm�����w�T�& �ʏ�VUk`���P�A˾�/x�@�fX��@����ĎN�(�6L���Ϧ&`Boa�6$Lᵱ�J<�o�>'ڝ�P'���{����sBj�Q�+u�VC!0�fTh��ڒI�����x]C/��.x5q͒p��N]�0���!pb Q"
A����a�=WCN�BI ���l�H9��b���|��{o���yQD�t���*BR	�Kw�a>$�f�z���Ό��Q@�!\��H�k���'7>�\p�X���XMc(U���ąֲ\�u�y���<��tu�����,��~�r�
|b ��Q���5�u2Af�c~*��z�n���V��+���w��!�'��V,�j;��]^0���Fw�n�U���M�,o��k^e�ޚ�~��Z���vVޛ��F�*�!]��. �>�*��5�(x�YŹ�G��Dű�����V	> �}��$�ss��w��3�����P�U���Fg��m�s\�$��l�g��Q���z���� ����ر	�(�32�4���H�΋\�'�|V�u0I>'{/[$�N�.2�S�vD��4-��m�B��@&bB)
`��� �w��/b�8��׹����e2I=ٚ��}Z�����{�kI"5BD��L�	N��F�#ڋ8�ܗ;�����۞y%�n0����>K}$���F�]*M��6�6�zU�Z��X���ƣv׷/��H�3X��z�DJP��"�o�ڡ$�(�������� �3�9�O�;��G{y����*��1�?w�V�X7B�w�+�[`�.��$�h����:����/���k>%xY����s�z���8{�V1[�o£��n�gm�h�z�8���"��9{�����&,�c�q �ݙ�0A:��P$d�G��2ffBOUOTi�
�,i
�$�Tnc`�F'}�A9���Z��ޭ2	*&��X�)�d��$�㕵'�^�m2�*���ݚ&m`&-��H���E	��ߍ�\�0��o{�$�B(����Lv��.��u��ԝV�Ses��NG���>��}��$>� �����e�d|t�ʓ�̽���V��J��,Ru�$�w�D��S�*QR	P�7z�$�zLnIv�n��pd�F'{�Ne�6	 �V�KEusx�	��)B�B�3%�gf�N��Pd��;l�7-&����oN�y	$f^�e�&����A��
�֟DV�T��J�vn�$9�+���?:����Uk�ZO0���\<ou�� �f��F�|�?�D��m�I��[[sE؍�UK��I�zz\���sEe�9��v�)%����겣B��F�H��N��jQ�� L�L�J�=��A ��lF��ngf���eeTP��ΦHf�mUՋ�P��I��L�0ŕwI�`�4�:�.��V�Ŗ.\�듷O5��̩��v�AFA���+k�A �Π�$��m3j����b���{�B���|o{:�ܫH81	���A�[׬���J'�����E��A>}٭�9��� �޷RE]��U�1��r��DJ��EO���F��d�s�u�A>=�f8thvn�@�]�sd�N^���;l�J:W�wBC����A��C��p���u�y�.�qU�],Z,�� �c�d���f&$H1bTW���a����7}����]�x�$��ݯ�F����ЦR`�z:��8ށ����7��-����;b�W+���w��κo!�������c�\w�z|�_J�T�kɥ�cB���St�g'�o�p�Ө,@b�rG�1�1�:ə$x����2v��>^7Ŏ��l	�u���
�Ʋaz��L��۳B/���=G#[�:r\'�ah.��d�[���m�	��\S�ڳ���0ێ���t�b[�r�Sc��'��^1����G=
�l��q�����s����;;�Nƭu�Պ�LsY���[75�Cti�n�=�7���F��86s�b:�SN�޸v����\unͥ��	�C�S}���I�A�ȿmRm5ם��H'ڪ�(��m�ؘSsδ	7y�M����AFA���ӕ�$@��j",��EW]a$�^�kd���@�'-wcq�VaD@&fHH��׾d���(I���Cs�W}5�$�v�~'ت�(��ژ����EH%B���v���aOrɿe�$��ôA6��(�@���}Awq��|IȬ�#z�D�
}
 Ć	��H��������	���}����A<��(N_g0r���ZOU-�1*D���1<&;uYv=�ֶ:|���[kt�<�=����6��f��1Tmcg�i��O���s~2��Fmb��ro�M�����;��A(+H��7�U�޽�� n*�.*����y��dh�b���30�23f6����Z�p��dlv�ܺ��f�C�ӱqpP{
�j���$�ȢA#/s�`��9W�����>��+d��bfB�̭�>$�ͦt{do9� ���h�@���7%��(���	Xwg���ˣ/2&rEy�h�H�����w;h�<�2f������]�T�DǥJ*|�-�u��nn��-&i�(K"�zh�Hۜ�$�~�j8}݃;t�F��	/�C#��vw(&�Q�m��n*�g�ZwE��ӷcV���|���{��)�(�R7�U΅fgP`/w�� E�^��z�;��|N_eP$R�vA��5d�f.O�d[�J��)�B���I%����p]ݚV����d���H�10Ro�|�$K��I�N���i>"q�L�̈���0��Y���YҾGdJJ}T8����DV	_�N����:��l�i�cF��C2ܬ=wĎ�k�:�� n��H���D�a[$��24Fer�����AU��?�]��d�q���������|�/`vѵi(�$��	�lu�dt�ʛ*v�V^�P�H�[͂I/wu�$b��EJ�gU|�{J@dI2|I!
e4���F�;�����0N�Mշ&���-������,�V�BJ;�m��|^v�0I#>�+��Uߦ�����$����{�\L)S�aH���[�� X�LgL_\�h�Iy���b��DWYU˴�����Z�(ᘙ�D�LD�	t���p���� �o'5x	$����T�(L5D�@2��aT�&����ߥ�~g����O�S�vg:�:]t��8ڍ���e9{�E�೅���������Қ9�'�^-���i�=�����p*l�r<�G �#kC�2[͵?
�o���pd�R�bfBq����f�N�ц�:��Uuc`�}��ENngyy�޼�i�5p��"�0L� ��3g����^!j�v9#�v]�e���c>��� W������1��#;�:{4�ss:�-j������F��s7X`�F&�+ċ�ڙ���)H)A���l���sȨ���I�'�}I9ٜ�$Ȟ���WT{j�n�dd�
T��R�Fq��������׼xtݫ��IP�G����v���_�̙��������gؽίm�/7M�,���b���@ ^�L��յ�'K��#� ��O'� B�L0*�;޾�w� �ez���s��uRu�	Q�6߾/{6�6�J��_��{}�k�*v��GUDh�)t�(.)�rŴ9oP�ݍf`�����"M>+6+0;/&�wFo����eG�RI�s2
+�Ὦ��gv��V)������bP�ܨ�0Wn����V��׏Y��?>���wڸ�fC{�����Q���9�_s�2�nq���۠���6[�*�d����8��k&�uR)��ж�_�R�o�`v,"w[m]WY�-��쳤]Powf������ �H�"@y:�!��n���7���+"yi��R�Q7��nwfcs,Z��{a(Гy�e��ݡ�%'{�M'G�t��rA�n���XF��k�4A0I5�Da���&U�v��	v�P�;5GV��$ڨ�j�l��34M��+#	@��j��UN,�X�EP[���c������nyd��srP+���
�BD���ͩ��o�Bwy{�=[��]:������<����8��r-�@A$�ɍ���R˽�q���wg]<���f���T*n�@��l�ʱN����gY���^��E��Bͬ쫹���>х��Pp0H%�9|4��y�J;�/8�o����C����xm{���rdw(t�k$^(^�eF�͑��}����ƾ]Q㾣�\%�	�;��۞=��:�Ɲk���(���+�����8����ݝ�4�[<�
`>���(�V������41���U��|�{3dZ��D��ĭ�P�6:3�*ߞ{wٶ��C ��u��[ۋ"y�y�N�fKڨ����|A$�<H$���T���LZ
�[h��+keLR�a��JQe\5�q�#���QVj��LR�m����Z"�ll��������E�L6�űE���iT�A�hҩ�U��-T��*��**�kPX"���0ŕ�,X+m@b��TE��QZZ�X"�*�
0�D��D�*�J�UH�UT�)ic+�\1F(�p�U�j�c���*�n,+qL"��� ��"������UX)Z3�%��Em�Q��ԍj��B��QT+%�U0�iZ���qh�\b�DJ�Q���)R�j���C�-�
2�m����Z�)J�ڌ��*"�RL����ѣ�1�e�j��,jQ��+��YZ�Ҩ�дiEQA.1LJ*��qew���ɁN:��J��-6��rs��.�[9�ݍm�q��ny���wsț�ݳ��(qO]�K�]��9V��q�;QF�r���g��v�i�
�j�h:�h�s����.cs�H⃫r�m�v�U��*��0�y����^��1���%���܉��u�{v�Y|�˅��9���gڼ�5�˅M�����Wnwnq�$�t�����f+��W�n8`�b�S�����f�=8z3��i��!����Ni�=+�ڂ��|���	<N�����������4��h�y�e)�T��$��9[��c���bk*�E�GE؋:��6L�;�s�wj�]z�ܳq��f�v��Ɂ�9��<��C���҉�����Зu��+���v�iuѲ��=�<�5b9œe,.��q�S�,�yn����p�a�Ѻ��8n<DY{A�nn9�pIʮ� q�t�q��1'5�Ob�v}�*Q.;\=v��|F�8{]�xŴ��yYM�7�+Y�%��r�q����;N=��ۖ��t܏iۛ�4nv��*G��r�:��<p!����G�u�Y�v�ۍq�Ů���۸"y�	�s���Ż%�5����7v��]s�m� �w�r�j�n5�s�n���>��iM�����W�"�ӧO�'�!,/>-mԪ����yd��}�f�&��<shع�k.�r��M�Eu�A�n�-�A�7�%km��=�\�^)#:�v���lk�-�� \78������m�m�k��;ڰ]e���;��������,�m�7���vV��kt�p�}��[��������z���../����]i>�䝍n�}�,���܀W�-�ug�P��pGū�+i�"[�67m{�w;9�m���=��MײM�7\�ٸ��ӻ=�z��fZ�����k�(�n9�F��x1�v{n����n;�f��e�;���uq���h0�ۛ[�j�\[l��qn�=�W+���udg�#V&�g����+l��\K�ۗn�G	�Փr3��힚��qƹ��wM������:��+rc 7�$t[E�;<�V�VT����g�|e��ݲ�{d�ѮI�P�.y6:�ն����������n���'=Ri�����B��q���7�;a��
h�=��z�8�}t�9��MN����[�T�stB�D۵�p�h��<�dd۝�.ڵdF���b�Cn͂���<@)�Oy��%3(O߾5Ǵ�@|��V� ��T��S�oc���y ����ۻ0�J�2 nfXH���9���J���c�'�0m"��)�-�λ� �/{f�b���zyn~�{�ل����Ծ	Vu�{��R�@|�v�^�σ��Y�S梢���lF�g]�c�l��=�LA��d8jcZ^�N�鋌�� Fg]Z�� >/�f� �Cʭ_���'Bͽ��iZ�H�Q3 �D�LTR3�@1�ǔ��M�w�G� ��˻� _n�P�0��=�9M���}V�T7�����O����7\��m�퇑��[�d�-Ү�θx֒�-1=��,�`W>���� �����C>QA'B��� �au��e��l�T��;��l�3(N�b�P��K��k��	�z���L�j��u�W��	���Yft�A&��n��y#�6��M����T�V��"��#ng<�:*��'��i�L��=��^n�P-��{�o��Z��2�^�}Q����{��$�Sd@�̴�y�������6��9��t���u���7{�5�Ȯ#�+�o�b&~s,%0�+��]י?w8�� ��ʯP�H�#� 2�����Tf��ӣ�$��e���w�*��3� �p�g��@|��W�����N���	�sT�ei� ���O�ʭg��?�?���ۂ�k��ڥ��wc�.8�����zY/T],c�r���b�~~w��f��K�3�>n�A̮=#m�fom݅���}M^�A;�4�`�"��$�N}� rɆQ�՗v=͝�sɏU�nf�~�Ā�+H�@�fom߭to��<�C;j��
�`�`�T���Bu_��{� �����0������h�:}3�|����-^�;*E�6�}w�]�n5�Qt}N�<���r*իE�����+�oK��H �+o�3{n�2$v�d@�̴�m��g�6.㳶/��]�A �Y��v�v�s:n���{�܋���3���<��f�s)���(i�W>�h���l��;U��2	Ё8��| �g]��os:iQ���ڛe"��{���Q�,�S1LC�-8r�;��.��rp�r���bݨ�n�kd��E��Y�ϛ��+�9��QVG!De����ͪv�@#s:j��w�ꕊ�q �.�:�+/Ec\DĈQĞ�HN���<�%��屵,��R6|ff�� �3��$=÷�|gI�($���o�aN%�T��˻V  {���>�A��>�ݸ��n� ������>uP�;T�l�3(N���K��O���؃���v6 �ٛ5@|�|F<]t.#Q�F�g�%b5U*����t5�rg��t�Cu�yƞ>u���:�F����'nE��ƅ2�+����zZ���"����Lo�W��jâ�j����e�So��~� ���C����눚���=ݹU` s:k��E��|z���]���?���Ȗݷ�9�)�Z����xÊ��7ck�-���<��������:���v�s��]cb��K���|G�x��������	�/��j�|�7/f�>�q��c�#���!���32$��o�kt�W+��T��e� �Tz4'����,�y��f&��ĕ'.������A~�����'c�7�+���H���X	iW�yӏ(]q,Q�
R��B�o����6$�/�o� ef��8�-z6�{�� �u4�*'t�m��&e	�|s�i� ��}�j�Q��gy�t���^��H�zG� >V�.�j:�lӜ�-���kl����"�m!��Ks_)��oCw�J�ѻ�3���ˎ�;��;ɷ�Oe�MT����C4��}�4-D p��u��Uc<���f���طug8�������w:<N�ݰ���۷b�{8�A�5mԦv�n�K��g�[v��a�fY��9��S� �t���KW4�{�n�u�ˬ����[��A�����r l�5�v������g�.�ț���x��X�ǝ����}wЩ�6���a�pr���1n8[]r�]�Ar�m�������C�{`ukUA�my"�+�hd��u�#��qs썷���?��[���� y���H �^�o=��Z{ڦ���ޱ`���wzk��zG�U��=e�3)�RG�����Aۙ^���e��7N�>��> ��������&i�����pNv�%A��T�$uC���7�y�vq��}�n˾�� �/�m�#+��Ղ܏80K>��J�@�n��uِz_E7h<ʣ�F���]�� nWI�G��LV�ǟ ���<�iǔ.��8��˪ۻm�WWޥO�g*���Ҷ�ZG�Y�v����tҢ��;�*��3�&�"�p�g�gk��Xn6�ʻT`��B\\�Ȱ��4QN�����Q2��5Ǵ�7�ݮBI?O���&�b�~bo�Z: �N�� .�6�+��nDCdȁ��H��:k�U�w*sZ�=��	3Lj�Mo����������pO��Yiŋw_q�)P�wT0����*UZC��*��q0sO<���nll�ä6+�޻� ���t�DLK�،��M����&�jI�xs��[����/i/P��2�4�.Vϣ��>U��v1 or�j��t8 ��Q���֦����=��q��Y{�E�� #k:j��_�j����z����]W]�`�=4&d�}$���z߅2RZU�(l�+]�7��8i���K U�ݻ�՛5CoY|Cj+�s?���@k=��Χ>���y���s�vӴ�����!�d�����߿;��`M� }k��WX �gR� ��=�;���7<��ջ��b�% ���a��&�*"fP�Q�=Ǥ;�b'�ݘV��Ӫ��ߕ��ef�R���y T�x Ⱦ��a�!v��2 U {[Խ@ �^�@ ��^�����-�{L���#��':������w�mM��mV��c��S�t�3H\�Ôrj���b���s����yjwj$�e'��r��y.�٢ZZU��Iy֜�Fd�*Q�aCL[��u��Ϣ&s���Z���/P�"��| ���[2B��z�S_P-��pA����GP�o���7/:�Y�s�;��cۮ��/~ۓT�A��#��^^�ڲ�r��ksS�S�;f�^��p��S��(��=�ְb���:�QƃX^�KQ$�d8Й�Y�D�d6˚�� e�������5��N�^ڴo�[�4�`E��)ϖʆ���
������A]��ܫ饉̱�޿P E���E��]���[�l)ޏf]vvd��T>�T6�&I,N�2x� ���V6��|P�	��� 
Ⱦ#�$//���YSqH�� ����<��(�r��h�h�x��-���>@طoz�� y��9nB�ڋ3ڪw�ƾ�ΙS�sU���{���*���.Tf_�
s�ۀc�ª���l�ߞ����.&6ۭ��d�t�Ix��SIu�aO�9R���o]j�@�͟M�6f������	�{�� "��n�b���̽[���0��F��Z�Ҿ8Vk^�m��/Kqv܍ܶ�h�!�]�qu+c������A�1�c��K���fgU�|�����
�^���.��(��������^��aI��Qz���g�v���^��_�"Ǽ ٛ��w�y��۝��ݜ�^zI�*��d�Lp5��H���Ӵ =���z�A-����t��X��Si/$v�5�l�Κ����ɇ0��B��2N^����[�3��Xoo6}@��F�ѕ�ro"7s�����]����ے.Gآ[ޤkz}@��Ӿ_�6*������ $y�J� �_�}��#z#�XEJ���H��"Sʙ�.�+��!o�R��ٺ���윳��x�z�u�=t����sYD��S}1�����@�n!�w�D�+۱��N�9��\͋�9�{��vn�alu@w����׳B�*�L�� �!�ڷ����}�0�;��`kan{a9tZ>���ɺ���F�����v�l5��$��6�뉮"c���A|2��Ӎ����������؜�ɵ�,Aص�!���WZb�-���������K��m�z���xzfЖ옼��W�˥��a�v�=	zxw�]-O��z#p&�[s�������3״�JpE��o^��cb��^� �_�����\��}w�M�^lҠ���8��p�$uf���&��"�IΛ������5H����	*hO>��f\B�F�7.� �8;!Dˆ}$��8�]/Pw�� �zB6$��7���w @^lҡ�}e�����ˡBc��
FU>�sW��}������ |ޏ ����	f�%�ވq oO��'��^� 3&a	����� onի7&����YX��_O�g�^z<��^wl�����=V�p��a��X�0dNu.4��s�/VT�$����>�ݳ]�v٬���m��πd���նN��vp}�q{�?~�'����-^�PI:�H��$P�
���Ţr�	w
c�e9�Fl�躎p_t�'���q�#E�x�뿦����%v���=����� �W7xp���©κ7�V���23�����G����n����B��w��=���8^$��GQD=�yH os;j����|���Ƿ�ڀ@+/=@ ^wmڰ~�G�F�1�����#}Ы<�S<p�=>���;�j�� m�K�+��].�!�o�1�U>W
8R2�.�ܻ��D����bh��:'b�x� $��{��vm_�3�m�MQ������o��h��̺�'t<K�� ��H�#�������S�(������������n�Nfa	��1�}� �;�jՂ�m�K&��g��[���YQI���:�ZX��	��F�>o	~���p��UP``��:o&�)$J���]�I��ΕT�.�yP�ㅿ�b���]���7Q_��V {y���@ �����)dQ�.0YW��79�b�u�7m!����P^;&pK޺��-����|=���^{^��;�;�6�>������d��S��Z�ht�Q��`�MN.�ܧ���oD�}ƺ����Mg�(9o���������V��zT�Ŝ���n=���B����Fvs�g�˹�Z��f8�k�44�������-��{��׺6BP�jZ|��ÈCĖ-����l��|fT�L�0�d��@O�﷡��qQ�Q��1�tM6�Z�duF�#`זٷ�V�W���=�E��>�G0<Iv�sy��2aRgb|xdXK�3ze��,{��7d�ۓ���o���5�!�٬.�x!1=0�t��l�¡�h�A,��l"��;���{�v�s;�r�Z�gVNN�G/�?yQ�#<����g9'L9�k�0�y��2�U�t>�$7ݖBT�����y�}�(�K4�8A�([��{r\{�?OBE�t5n4���r"�GC�0b5��Kp ^�[�IChс|�� �.*�i¬*!U�h�a����9�K8=6�sĎ���G�U���,oo�kLK
z�z&,��#؀��+�CyE�M���b���cl��`�֩m@���Y�Nm���u�a8��ƹ� �{�������SU��S�w���xmbL�G/vo����e7֢ȋY�*�7(\����n���E�����\��G�fo[�	w�c3Np��k���{�i�;���DS��$(^�-�v�]Љ���������%Q�*8q�1�m�J�����jVZYl�Ս-Qm��EFJ+UV��[B��б�1���`���ʅJ�ڔJ�TX�0b�V��c���-hֶԢQ�j5b*2�*Z��Z���Z*Q��V�*&J���b&)�%JZ�Ŵe�2��i�01�ˌ`U�B�E,�[�c	��[p��4�cV��&-��*%�m��qDV6��,��KkJ*�%���,��֣[qjE�J(��Dcm�֢�H�Z*��F[B��5��E��k
�Y����akA�®Z�Kkm��%e)\ch��`��jԪ�е�����U�-R�q� �ک[m���AYme�ږ6���֢6�e�Q�PJ�E��Z4A����DiV�km�V����#V�Z�.\Zֶ�j�[KTj�k�Tc-�Ֆ��ҭ�0a��Q�lqF�(��mUKJ[KD��*�����m��Q,Z#Z�*(-K[kK��Ueikm�KF�-�F��ZU `&��U�6�$Vfuڱ� �ΚM!X7�A�JT
"Qpǔu\�Em�"� wvmS��l� �X_z!���C Qs� �ۻ�̏7�TL��䨠q��� $���.I^�Tunǧ �nz�����6j�ذ��y�;�j�>����0Ȇ�D�nβMƻ�ƻ#��:b�ݎz�0�u`z�������
�N��Fϯn�l@���A��c��C̪�Q���� �u����t�^V�Kp�o��*�K���` y�T���c� �+�����,�]w]��y�["&`��P>��� �]��C����=ۅ���j�y�_P�����ynE#|dH�LC��{��t�ݼQf��xېy�T�B ��� y�щl��4wo@|�:w���m�;��Ւ��kk�0�� �#{M$R1�:��b�V]M�r����DSY��~%�C�� :���=˹�8^$�����R!�{�H >�ΫVK}�Mi�@"��i��K�G�_�y��vO?-�]<�W��X��2'2Ȑ���<����ѹsL�y��%�۪)z�ׅ�f�lWͽ'L�� �$ʸ�m\�,%��jP��Ϊn�V{ތp��hg�;6���/}@|�T�\(N8R2����Ӵ}}��XwC�^ר�4��x >/7:��O_G)�o��.=S�
�ŦRi�a��!:�s���@ ��ڵa�71�3|c�+����������Ϋ�SY�l  ����H����1vC�y >=��� >
�ͪn�����2u�m@ �9k�$���C�?9R�7Q_]�v��l��)�%lÀ{�߁�vu_�0 �Κ:2vjGgMJ�`�ȊJ�e���������ޘ����eb��u���-.�b�����ru�y��M5�&v�.a�(BN��!6�h=��nE�mt��\I˞L���m){]�Qm읷9m�e	Ku���+��u�Vv|�/E���v��8���/`�l�n�#&̛���k��`�=gvj�kf��G��Ɓ���Yշ���v*�p���mV�m�(��Ȝ(�9HR���tܺ��W���Y�7$���r��3F��9��{=5t%���YM<%�-���f�XnNY�R�9طkZ�[TO���@�ە�}~o��Å��2C���l�Ϊm���Ty.�߽��U�ޏ >|f�m�Z��"d�$��*�BF6��@ٙ��Ti�R����sj�`ngK�E �/n�3�}Q�I`sZb	0�i�H���ڰ� {����K[���Y��q�M_���7snՌ�3���-2�M$�'T�~�UN��p����W` fl�  ����ޘ����me^�ش���*-%	(������<�����KM����:k�vWm�z�	{�{w` �36j�|ކ6KHh���-���`�O F F��n���-qr�&���H `��v���n1��o������S�*Sq��컰��l��/��]�Y>U�\)>ۻJ�|������C���
�
�D=�{�%Xa>�4����"�Պ���T�Ά��Ɛc��ŷ�mn�ը@�H�D���q��i�������]lD�#��}�a����m�M�C�ޏ$��n��-���1���Vm���*"~j[�rTW��}s���}>�H�*���<���U��gM}C>@,/�,U=J!��)U������#�b�f���6ay褒G3�]W�Q��nw�H%[�iP"iZe6�%DLK�5���#`n��j��w��T��[�[=��D�W��(,����i�")�vx}s��j��ǌ<�9�!N|��SV�1Sn���+��N����d?À&fI�W�+:�@5�Ͼ�����v8���q��z �u�P�0��x&��L8S�*Sj*�ϮŤ���c�.�b@�S���|�v�f1 �_��w��������ɯ���4�q��&B��{^��|��W`�^��1�dB��T�U(���ڗ�D�۹��h��0�IQ}B�^~�ix1�y�О_�A@P���f�1|B�u��������LMs�Uk�k<��/vk�� ��lm�c���LI�ᄌN�n�2��@���� vvݷh���^n�
�68�Q���̓C���I��
FU>��� ��gR�c�ݵwKv��v���^6�H$��{�� ngM*a=]�z;ʷdƣ΢I:wc	�m�.������(�ݲ�-�JġЗOg� �\a�2L�Z��m�0$�N�[����!!�{uݢPH�gM?$vU�����58����>@����X%8�v8	�"D��H��1M�*�#0wL� ��ݻ����5C>	�?tG�ُ����Bx��|dD�
�,[ϮҰ@|s6��  z9�y�4dy[Ⱥ����v�� �Κ_P%~��C<�`PD�TP�k�\��̻��|7A3W�v �73�� ��Jɚ���f�s�@�љ��p�r�Vit�E(�7U�2�����cI����!�=b����3;V�����x�����m��*<����S��<��y�v	fB��DD��7䨤���ר@|��s1���r~�����73�ͷK�G�b��6�ڸ͇���'.%WE���]Ս8�j9�;�r���̅�j�����ۇn�=�O�n���}����H���$�d���U[�#�-�˻V0��IP/E+N)��H�A�uH���?�Dн�Vmo�  33���ly}�� �Go���޽�SSȇc��"TJ�����W��[{>^��Z������U�^�� s6j����݉Q~r�SL�M���yyE⽕�����Ѐ@$���� �����fz�=�v:;j*�=��Py���̲��}6� ���;d�]�z�H��zi"P����Sd��#zEI׾���Zir؈%�	5AɃ5�q���d\��I��{�P݌{�0���Ui��+/,uq ���P�b�ן�nުEU�1��
1"��G�9�˃�������q�}�q�g=�k����y.�b\x��i��/;���Y�n7krm��h�}�*c+��S�sIv��Ǘi����,z�\g�"H�v��Vݺ��(�$ ˮ�ml�k�y��$=�&�e�D�����۰��cFշ\��X��x�Z����$:#��e��;��vs';.ֹꫩ,oe�c�Y�q�X�CkH�z�]�f�-�� };�����y�ȉM�n%ɑ� �r��4 mm��xř��v���b��C��迨`�6�H1\{�Cn��)�z��^�� �=}��+oT� +��z���������:��������[';^L�D�d�T����n�;�ꌗFꧪfc,$��7�ΚD���w�HK����1d���ij�㻶�-�Z@���}@�^n�ݠ�����|��y7E=@'yu^����c�aϥ�AP���7�Z$�Y���Y�7U�}�ٍ��IϷk� ���7��Gl��2"�v�DFD��"�`J�^�Çt��G\ݰ��"����d����ۋ�k���!GJq1
	�f�E�{� ;wv�X �[�H*{ٯc0~�]z�@"��n��y��DKi�q.J�A�Ж�dI��Yˀch��þ��������r����@�'����*o�K�#*{���+ޢ�Ds��M���vD��yk8S���'n�9�,�ؔ��$����7{v��H��n����\�'�N��/X��*0" L��z�� KΤ��lU��E�y�|ޠ�ݻ�X�6/:+�<R��n�2S�'�Y����;+��� t^lU 3;ޯb�NmO����
�O�8�W@�i[�!���'���LF�uQ8C����j�"ԕ�o]�`$l^tW�3�fuy�G����EQ���7��֪�;�GF��4q�g����;�]6��	�붮A4��`?W�V�q�~����`��/6��> ��^��\c�m���Zf��$�b��V�(G�8��̲���^t�Uq鮊��5��ۡu��O��8A%�y��~I��D�%���ML4����]qDƘ����rTW����@fw��۳��vu���=L'Gg.s�:�Q
eGD���5������wT'��v������{
.k�o�a������p�u�sq���x���^<�۵� �2/6)P��ίP_��&�7B�eR#�{u3�]�iUlrugdy$k�r�H�wsk���#7�o�i~��.1�G�}�>�R��n�2�)�g�U@��[����˩��SQa$*/n	$��uSH��{v�Z�5"�F�
�D̅��s�c�t�D����G��kD��It�=�ۦ�&T�g�󡾗a�JY� �o�h �w�P ���ۻA�-��Wٗ��/s�FF�E/�b'y�^��lG�˟��P�EM]�v�V,��}��<��h���� �Fon���	h��XDsq�^�΅T�`�fYQB�몠�v�X| N�mIYp�oEw�A$�k�XI,�ݻ�����|�1&UC	��E���=��n�}�ꡳ�������m�%�E<MY̙*���X$C�w���a�&N��
#�q�P/�_�L��z ��5��s!۽�}&��ɍ�r��'W4�]�m����5=n�Z
�Q	�M�Ц�t��<@�ίS�u�sNӄ�Rԑ��tKI-�ͻ�Im�O��v��i�;Z�L�D)��Fdc����sg�a������6̼��]~e�L�ۇ-̱J~h��y�	gfիy�T^T��{���K���ܯP ��ݻ��r�LB��D�Tv��@fy��8)�~v�Ow�ʀ��ۻ��Κ���m]d|�sj'j]_e�oU�>��"(r�����X|��>m�������{~ ��n��s�j�+y�'�N�̲���EC΅9�3�YE�|A���ݚ����"��\��o�<�9�tz6��iUFQ$g��q��wFk~N��	�� V�g0ﺀ���,In��9�V����h5[-9��:-�HH@�����$�i$$ I?��$�	!I���$��$$ I?���$����$��HH@�Y!!I�䐐�$��!!I�!!I@�$��BB��$��	'��$��$$ I?�HH@��!!I�@�$�H@���d�Mfu���?If�A@��̟\���0       =          �                  � XD$� �B� �("(P� � RUJ=�)*�B�)V̨�P��)
�� *E6b���J ;�                                    �        @�R��vƚ�j��p��r�1z�ڨW��4�)ٜ��9�l7��^�3W[�T�[�w[[-�5Jvj8�T��   �+�ڕ]J�wZ�� ]C�]g&�Ӷ3V���C��z7 r�F�uW�귻����y�:�=���h(�)�   x        � ����s5N��u�ҕ���S�� u幽=��mU��N�u� �W�@^�B�����T*��+�  }�^�@��jtt� 'C�5��t���Q�sk����� <zf���<�PG��T�Ð�(Q*(
�  �        @21z�uum+�5��s�oX� y�� �`�������Kf��z� 舦�
 t�x  �Ҁn`x�P�(^��<�R��RD��  �|���M�
:z� �
�;� �@җV�`;:7���{� 
=��h^�a�g�Q�m3���t��JF(��  �         !�U{�� ]�J��*�4��� ��Y�WN�t����9���:�8@���I*�S�  8�z]6�� �� �.��
�-tm�nw@�6 �� �L��
� gkiɠ�mr�hQ�5��  �         }�e�U�Z�*��Q�[��U9� .�n�ڛZ�[�3en�iatΪ�7 wZV���Ӣ�YU�(P |   ���ܴj���ֵ�� wZswZ�B�ճU��N٪9ڇZkp Lu�m�p������ӝ�P������O@d�* �T�&JUM ` Ob�S
j�  T���
J�3P ��S�)JM�   D��S� '�߿��� _�o�]���)�������«*��H@�����$ IX@$$ B��@�$��	!I�B!#�������lz�:��R��j��BE
͕�E|4���������U�o'{Gi�6NL�i�硭��2�k��3���K�=i]�$)��d�|2�J���L��^�0�ɛ�v����p˻��둼����2��9��ۻQ�s"�)��KG'��Ǖ��M�j�p�����% �J �)O �߮�_ݨ���ѽ�M�C�f�����LJH�ى+��pDs��;D����ݺ�wnN�M]���H�qG���kD�Cs�H�)�ݮ�H�D�Y��}�~�j`����/���k|9G5lY������C4�ӛٹ��;[+WV�j�{�5Ȭ��h�>���.�%�}�{�vs	�C�\k�Ʀ�B�p'��F�GI�+��ʹ�7���63�D����:�ѫ4p��@4����7p��kA�D	��&ܬ#Ķ����X?\�ۗZ�mwm�5>��1�&�w�Ҹ��SԜzk�f�������
�����z ��8QGd�@�� Tu�,��-M��qrtɷ8BC]�WT6vt�sUG����7�Ӎ�A�;b�h���qU���TF� q�X��n	�Iı=%܏�Z{"��z���¬Žd�ް.�נd���F��W�:0�x�n��!�{�ogpk=����5Uѹ]�pu9��gH��N�K?��$I�U���}n2yr��?)ǲj3nnĚ[�9e�Σ��2w��u+k��.L�1��8��*�{ӥT��R�p���nӔ[�&<��yF�]H"�i�[ڝ�	X@��1��nX�Z,K���o��ۺK2�s+�;�2����6��طr684x%��4¥���3����j�q|u�=;�f�C�jû�p�2��hF�n.{�i��l�qח,Ǭnُ�v���0�F^ܺ:=�V]���qh٘2к��9B�s�1��7bW������'���q\��)y��i�^vuy��^�P�b�r�B�:m��ٺ/d	�E�ŭ<��g
˪ �8�zBෛZ3���ם���㷺we�vV���Dq6qՋ0"�ҖɱE��H�"���ᓨ���%�ӂW�R�A��s87��Z�X��ޫNE�j���8
�!�Iu'�#��E��v&��8�7��rL�p鿹=����iO��Tx�C:�8sRf�U����nn$���Ȥ�:0w�!��+#�Eݲk��nh9��Y���NZ�tZ���u�ٲ�z�8�@�AΙ[jN	cΕr}Ò� �i�ړ�q�Wn���\s�)���]|�<4v��� �׍�3L�of���i��{���\OH�<�Φ��Eױc��B��=ɝ�,QwFs�"��i�N�,��#����#��e�՛k�;�9L/�=��P��f��i{�v�.�Zw�wzMo2wi�a�1/�q��NI��f�,�D�q)�T�z���Q��o�������w&���7/S��\��`=[�qpJW�[��b�H.�g�'��s���ٜ7�ZyM�?����j+�+Et�) �jy_E�s���GR|����n��U�陭���������p�� ��U.��j�Ej�2��ʅY�Ӷ
�P)W����]$��\�E~}�Cr����f-V��E�V����@�)��;¾�Ml̓I|�5
���ᮔx��9).C���v8��Y������w:���K����Gvˎ��Tj��)b5$
D�������R;t*�	rn�����pf���l'k�rN�<�õ��!c̋�\���_hq���	��jB��|���&K���#��7������H@��M��N�we]5\�v���,�m�v��sC��Ws�LR�n,f�;�p�)Ÿ��C'�e����jՊ�n\O�TGqB�9<�qa�C�(�;�٭Pg+:\�{9�,�^hr�j�˱����ʂ n#:�/R�0�c�$���ͥ�
6s��ι�1��OfP����@ c��")׺6X��nu#.ˤQ����&�6����i�ZYʘ|i �.(C^Ǥ-���n��_7&�\��v]]Z��S���n�����u�x�a��gB�ą穨�����vd��0�����᜜am�/J���\����ǹ
R�8���<aK�;�Os\\�4a�yv<hƫs�C7;��;4��|�0�Ӕ,���1����{
3��-Zͣ��z=�q#UwK˨�z3f��f)2�(��f�{g�o�o�%���X���7���d㫎o5�l�8�w�-m85�M`�T}3B"M�����vӈ�v��bc4��v�V�W2��l��i7[�ἐ�K��0�*�sCMA;k�)�6&�~�3C�
�+G�@�ۍ���ᔮ����4H/{̫0,E���܅�yE�lov޸(�7p�vA&ob,:��b����·����;ԤA��3w��:h��@�O�x:��@K���qM�-zy>�����S�6�b��x� M���+�~��~��3y��t켙|ʻ[5�9Ӝ��d��i�&by-[�U#ץ�%��2-��݉oR5�e���&�����w7��h �'F�X������d������Cqw.hq�O?�	�����(rvO��Jt��YS#gH���ˇ4?�8V��GH����QXN΃��TX3��n��� &��y3;is�T���oc�A{�q�/mhx��%��o���kL�eӐ�J����x{�Ы{�?Ɉ���*7-��1��d"vhT���B.���ek`!r�"@C��wvobkq��6�ܫ�Г�7��0&�������$շ#i���^O�:��=��n��૷77r���3������W	%z�p͛M=�9:Ȗs���bue��p��ܜ9�y��^�헎%թ������|���9]q	Z��v-9p���"��;&�Ki�On;���-��흛����x��mN��;.�x��t�
��4�-0�T];�H�� �Ğ��S`eS��^���ƴ�>�����9tū�@�r�V�vt:���byCS�H�0n-�of�:;�N�����*���י��{�x4����U� \E�(��k����\wn�v@�y�	Xk V�qhL����y�EUօ�Y�:�nr����:94Y��5`��[�K�9���� ]h�gi:�/��K����*�N��{p��ohH���M9	�oJ�]�p�\2X���3�L�R(3�qt���l�t���u�v��<lК�ƍO�����"[���*w��r	�v�w0��%)d,[L�jI�-+�Ӣ�\�����)�`�&��G�%js��>6G��ޗ�v��C�͘D�GN���V�� nJiE���.G4��WmΘ#$oR��ן$�����t���v�:�qK[O#H�N�Ț�v�?��jpk��6��懻�"�Ӭ�� �e���?�2���9q�Wǣk�{��{yRW#��5�NA�k��Nǥ蚖C��52&�h%��I�ƀrJ.�Wq׺�9�O#Woᒙ�Xq�����53t�'XxU�@%!�xr���;_��O yid:u�z
�7�\�� ��^���ԹCr���۠v�8�ӻܧ���Ml�}|�u^[�'W^�]��I�L[��`oA�~���K�f�ɻx��}��`-�퍼�P������U���Ip�
�}�f�.��$�啱p
��l�V���a�զ#q	I�p��h��@{����J�S��_#8�G�5��=#hܿA��6�.�s�g. �9zKv��R;eJ!�w$�W;B+,�����D|�#��cx?9j�}����:�k�%���B{���
�>l�{)蕸����t��m��H�7���C���-����p�k�0$�KV%(���F��楔�%A ���/�f��s�����u^�B�Z��k�NN��ugw��x)��	W��ê.�y7����mˋ+��םv�V�Pt=�s�Thʹov��ۓ��aE���v���O�NW�(��������,���2��=��s��Ȭ\5����0����N�I��r��Cc��vR��j�-�	�3H�_�"��g�P�t草x%ϻy˽������NV�컕�h����X�׃,=�Ʉ��W֘(q�0�V�˽��m���ƫc\v�u6��I	���gc�8A��5����՜m�p���Թө�n˺�v�t����������D�d�?�=�kkΛ7	��č�_U׈{_)��S"�ۙ��B���ڰG�c�h�]�K{(z�,�r���+�[����
�Iߩ:��w`��p�ޚ1;�ssw]��q�ы��7��L��V� �:�ņ�v�9t�e�S/J�r�k�wY�Vo6��I7 �#�w�ɤ;d<��s��c��k��X�TsK,�����/�O�͛�ol�,�n���J�6hת�_0FpuwN�u�g�X��x�����7-�8��j{��B�&t۬\�S�r<7q�.1��w�t[��D���`�z<,�ZL�gc ��ݽ�J����Q�����RNK�8��2�9��ѿ��b�Ȏ�[��^��{�r�L�s��p�Z�ɯJ��7�kK:I�4k����\����ɩ#���zJ�z%�
�������X�/)O�Mb�0~��L8 ����3�lkkE���a��vt�Ž���o�@{vk�:8����<:7�R2u}���^���ttz���{�=+�y��l*u��L.�P����;������t���b��q�vt5�=��+ �;p�pv��r\z^*<�]6�h��鑺�diAoDy~�gj8;�������{f�B��
]�nF�G��3�I�ٯ{k�˧tTp���]�f<^��~
d�m$&��j��f�P0���9nC����q�8ݛ�2�#����@֝�eG�~Xr���*;��F���	OY�e+�D��b�q˝���\3�i�\F'�3�H���N��}F���:��.@�h;�Q�#_�XgB���?v������������{t�/܏8���WL���7rG�s�ن��ܫKS*�kxV�n�H<����[Le�/j�����Ռ3��Y�m-�n��
-�H�𨾪r��QY������8to�Β�wp���M⮩{��t�N8���q��t�5G��oe��*��#^H��f�|S:�9M[`:�ysVt���ݐO��(c�<xY{@�I����3���^X'��zn
�͎�[[:K<f��k�∰=��E��ۚ����K8f*� �V	�j=�1L�(�B�Ȣ��,Y6f��[�;'l�!
ɩ�nT��d�N6�sOvɈp.�5-{���de�W����䭻�\N�tv��
����jz$�7�μ���|�	_a�;�d��{�+�3��:�{��h�7`ɰ����'p��ڻ����p���	����}���jvp(���@���s�3x{1�����J(L%�2��z�K�kp(.q#����m���dO�v��Ý�]�y[�;����u�y�~aFF A�]<�[ݱ�ѱ�Df�G���:�����V�[hT�Z�y��!*�d��y�aHY�a�`�;��[8�>S�u��ЪJ��o.	R�cp���P1�P�)	%bn2�֠P:�r,Z]�R���f�V�.9f����#3{(=�Ҹ�f�߻.�ه� ����Oe�q7R�j�f����ˤ)B�E��Ӊ�Ysy���rm/�O=]�W��A�Ty����q�!��p�"ABg^��1�d7�c��uú�p����;9����k��p'A<X�����#�/l�y�ۋ�L,>bi�G^;2��\�vu�\���V�=�N4��äIRL�M�n��'	���n`�6�5�;wPv�.��AYߧ{�\.
0�p�$x/��Θ��D���9ps����N������udt�t�}�r�i���Ւ!7\���Yb��-c;j�̲w��7ez�Ŗ��pnh��&��f-]Gc�ݰv��l�����+<�t����:^;��y�1�<�l��0my#< �!�ǋ�u�%ץ��齜�Ǉ�R�"S(�:��'ymxkt�w�=���n+���e`�4وE״��\�@|��=���Owl���8��Y����y3�vٛ�*�,bxTu���7�F��v��A�e/52ՕH2�v���5;m��>C�����N�]��?>�>;n���΀v��r˹�l��Fܐ�\ɝi��S������w;�m�1a[�wV���3V��q�[�>���F����u�PX��۸�<=��e�8�=dy�#gk�W�Mth��Mֳ_�Sςڀ<5�٥���!ju�.��v��_l�*n�_#���S4�]؇w=0��+�\DHq+l�\���z�Y +n�v����j�u6ك����4~PTkض�m��A�]J��������oO�Q���w2�'g_�Y����hk\��'o�&������P�څ#�YNK��ۯ�E�k�xK�T�7��kWW�к�$шE4�Vwu���vwtutuu�Wqwwu�uWYu��Q]qWU�]VuWE��WtUu]Vwu��U�u�WqWQwEU�]Wgu�uݗ�TWuW\w]�q���wq�u��\Ww\UQwu�Uw]�uuu�u��twQ�YuwUi]Gwqw]��u�Q]�]�wu]��tuwY��u�G]�wwwWu������QWTw]wu�eWugu���u�q���quQ���TwU�W]�]��]ݝ�]��YUݝwe]VwwwY�uVu�ugUVu]w]qU�eu���E]�u�$SI$�4�L*i	SHU��]Wq�t]�eU	�D@$$ $�	/wϿ�~�͚؛���#2����ڬ�pd���c�Q^���&�e�q�/�F�k��R8h|��h��D/�����AS��;�|l��P�8�<k]�/R�uw?���s�{��nE��-���'^��<Orv)B�ע��D*��,����|6��ȑ��]��#Sv����ʹcX<�9�9�0�^)�q��U�4�mD�2(�ͩw���*�sk$m.=7RΤ�θ3���HF��K�HsnL��xv�Gu�ZÃ��]\��U�ײgN�N`A�}oygE�(�sP�]���8�]C�:Ӌ)���n�m��L;�k:��á)ҽ�!�Dm�:��Z�0�l�d����(�ѹjJ����5��E#V�`�!��䞺���1Ӭb�uq�}��_�$�{|�F����,�vy>�6B��L��N��I7ףF%JF��峌���&Ω��OM9Z��a��hb����$�y�ү\��wf*���ᜯj�7#�-�3���3.������λ��7�nǬ,�~���ӞeKʱG1价GNI����<��;M�¼��T�β�ӗ(c�s�D�Dz�[�*� [6ի��I�Y��2lb���1C�F�e5nw�W_xh�3��XK���o����=�P����VR����?��!Ǵ�4�"mE�b}��͌4f� ��7J�g�E�엊�Xv Y���{__A��D��S�d*z���$=^0 J�k���Kc���g��q�1b}~nI�HiSYj�4X��sgWn��<�O0m�^�^21bk2� �o+
�ӛ<�����!��vΧ���}ۙ�+��F�|��Rz�M�3ܕ�~N�f���,�C��MJ�b�fv�kU�k;��TS7��/a�w9���݄���n���#�=5z.����VώT,����:�����-���������w�Ѿ�ppa>ڤ<]��H�K��C ���Gr��)v��MU�ooY���G�^�fݱ>~�+�JMf�'؞��;䠻�x�J���z�)��{�{�>:�s�t�ԏl��BHu^=�M�{ M7M���povq(zN�G�������0=�������`�G��f�*���}���u&�\��G����|�\B%�v���f�dv7^�E�<�gי��6��&N�!{������Q��*�o�[篽���qޗ��������|tv�����s}���%�1iG�T񹗵l����{	�x�uwU���ϟ�&���6Ê=B���9P�4.ǲ#��et�w�_����(e��25�pcr{m�:�k���C'H���r궜���jF�*�p�q$h���.�  v#�a=���W�����z9Z{�j��EG���(_��~���7����2RW��@����=�uw7u�'�gǽ7���ū�Z�������`V������|�D���}�؝��$�����j��z����nw������ Ê�>��x<n���1L��r�1mFUŦe��9�4��'�[Hx{8��]��t/c�?y�5�S�I���=��@˂KyQ��<A���H�i8hE%���j���oB챧��]��o�Y��Bp�����<���-¸�LL �4����Y�u6*.$�DC�&�K�n&�=N���k��E�U4�Um0��pK���.���Ȝe�72�Ҵ���Š;�����'7}s���z{4��b|�0�Zc9yS�G�B�m��������"��e9���p&hr�[Qt<��ٯ{4ȱb[��#�^��t�t}O��G�~8�oq�4�7r+�T����y;����i��:-�,<x�j>/�;�8�2��lv� C{%2u������m)`mZ��3�/k�`���ޚ��޲}�������\:�)f��t|L�.�7 �V�?;��~+�s��]�����8u(5d����YЙ����}j����`�:�;-�3&'S�I���e�%t.:��l� �ʬ���a�<k/D�x[�M�bNV^�̥s)��851���[�{F��W�S[ ��M���n1�0���پ��F3o3�?,��5f��I����:�p�Լ�mz�0�3�x뜟�J|ڌ���i�2�kұ���y�d�
�}�8k'z��<0fќ�o��w*��=�nooyG���c������<�uS�fgx�iZ���/&��:ixX�K<w�����R�z�`�Y0��g���ȱ�ux<��w	�>4�?�xF����(��
MWd�������ʏ��)�GO/.�3���zP�׼�����R�Td�*��p\����o�����-p�����|ۆ?/.i��+\��϶^�������*Т��ɚ�
�*񹲨����hV5�{P�[��4�W�c����W����o��g;_�S�6-ݺ&�m�Y�rN���3��=tB"����J"���6h�Tw:a;��		R�AjB��8q�t��6��v����~�N��^7تZ?���/�i��'�dBu#��O ��=c,�F��{��E�ӇK�sOyNLJ9�Ύng��P�N,�̫�<607(=�8}���GR'�:pl�	We��9��:�[��}`%W�Ěfx0���?��M͎=�i6F	ۺ��u{ {�	�z�un<���������U�ѕh83|E�����A��:�๡������LN��EM�d��+D	��D���in����J\����Θ��f��cB��y�R(�5L0��4��{��J���)8T��)�`�3�1!�7�U��KN�vD�j|T�ʻ��L��l��|W�'�ٸ����*Y��[5��*/�"^������[
X�ܴ6	������qk&�X��G���XZ�L���B4�{��" ���b�lc1�s�
I`)��7���#�"L��n�֌�x5��xķ�P_�v��Tʩ�BdBZA�-@uR���26v5����7'M�<�k��d~�_j�{�xe�,����Ĉl�N�P�֞g�>��8."��y��-{:���UmC�h{5�� %��ϮF�-3��L˲��US��0</�w�A�&�����r�;���>���4�V��v��Z�~����o�p��O�o�ju`An/we^n?�[؃���챮|�����y�W&�K��g3��KqR��N���^���VR����O����N?�Y%�j�>�`��UNͰ��;�D&����J_�q���eQ���J��C�h������rA�⯶�e�����TC<�qM����lS�۰,�iƖR�����k��z�f.@�v;7bt!FM'N�u?=�w��i�/�yJG�q%���R�Sn(Jb�d��#})S{TތZ��œ<r��P��O��v)���CZqM���b[=��0�w
�]O ��.�r�^ƝE��N��)�`T�R�8�LV<�A��m-�y��A��H7�vi���I�x���\;��sN-�)���^O����DÝ���L��׵���5��,�|_��{ޭ�Qo7��!:�&d3!��pj�q+���i��w'<�NX߼{;�=O�d���:<9�.�ÀdA�Ӹ��o$]3H�m�l9ˈ�2��YM;�ol�=��f^�N��ɢ- �)�r��<5h�Ǯ|H����с�����f� wN>�P(f����Ǹl�А�{��5J���N�Ŕ���XXP��+e��Y���5U�Pw���y��j'���j�7���+��{�x����j�x�E.I�.�c�Q�""^Y�E��u_�����������Y�7��{&��m� �}.��'wM;�=�4�c��S8��YQ��m�c�6����X���$I�Ow.2<��oh#����� �7�a�e�,]��d�]~�FL�w7�����3{��@)C�f��N�J����ÌG�����儣l���^>/�0f�ݨU.�vj2�G�	�,�j�2vw�N�:��)��-"��o6��JJ"qJeه"�X����T��ٝ���Ԫ�Ѷm26&�əIkU�*޾�Vk��Z�xjӜÚ�Q̣=��;��p2T�y&$�-�j�-5,B:t3����P�Fc�c�����'F��>�+��_����xً�q�	u)�]�]�9��%�2�J�l���,��x�=�ڈӚ�~`\���S.���VwdUa�,{.�٭e�;w(ZPs��+�Y�Xq!F��\��'�wr�u��Z.]��5�>�*#۫/-���Վ�64+�;�Rt�*E96��N=By5��b��z��C�J�u�S+rr#r��jgwD�nBBg]I�*qiCf❹w��s��zj�.W3YgI�0m͹4w �,�g���5��8�{^3��I��-��s���������-�9Od-�ҦD��oY�k\����)�ګH+�ۀ`��rm���̿v-On�=�w��n��r�7Kr2`�틶�b6������x9��pnb$��wT�v˽� [ԏp��\�^����|�jD�2o{5�������w��B^��2r�d�n#eг��Ƚ�i;G��>/w�X���ag`}ݩ�"�{���9������1���9���=L6���,̊�x�Q�����Yk�Hg��iG�L�Y;(����N昘���8}���6��ww�D�Qe�;���Qˀ>��p��2������]x�2+3CA#Y��xިn�ݙ���	��bM����s�7�d�ܯ��g8x-�4���.���Y�t���������{=�}�N�8{��xB�P;J�F���nc,=�KP$ZU�nkJ形�o]:���~�\�l�N,�y�����:�:m����a��<j��2pW�G��x��ע��`܃@�X.ٳ|�_�`�N�3���ӥ�yj�A{l����aL�\�ۯ)�ݸx6s9V (G!�I��ie����/-��8����Nrk��A�Ew?֎MyQ�eT���<������gN$����F�G6��L���~�:�O����n2�)�ܐ�E��_t��7Q��G�.�����0���R���R5���i��f����綐�^ �"�b���3V�F�f�xh�x�7�/FmXv��^��̠�R�B�p�S��7�!M��odmӡ-U�	V^ �s�ˍͫ�..���	z)5H���Db�Vƙ����2��0���2�Еz����&./:XGF����������i����p��q�`R�w'4)�[�<�����ۚ8/`��p�Sg�(Mj�8"0����O%`s9�r��>ns�˨y��zi�ь�02:gU��k���wy��08�==��h�;�Sv���C⹥�ʑ�����HZ��I�Çr �SeM�njim���	����.+MP�y5���r�yO�?gmO'z�����( ܦI�x�=�=�_���9i�w�w$������W��>5OHt�,�
غ7S���N�(��W�zm+jG��?n�x��p&h��gzj`��,�v�S9q�)��{Ϊ�q��;��B�i�A�	mi�%p$v4"����^�1(������V�G��wVM�I�����e�����4��?:��U�v�{I��є��m��g���*ڦ5Dj?-��{��z&V�9�v6���h�_@8�{�{<�s�-�Ȋ�[Ŭ8��<���)��d�G���]���^G��O#{J���v��.�<�{F���ͧ�uq�) �e4��j1C�g7�첮�{,n(��u�4`3q�e�ܫ����i���Ī�&<5s���M�Ӈdi��7�қ��M׋�����-�:��ihG�����r����V�3o�N��¯Jg[۾K)Ļ�E@fܳ)�en�l̬�Ҫ�x�+z��0�jN��d���he����G{[�g��g������ �B�|d��uG��^���^r���܄��$���ĺ���
6�^޽��8s�i���n�]n7t��·~t*�t痣|<�H�>U������肯�!-�i��b'��9�0����p�z��1L|�u���cx�G�\]K�ЮF�5����n�-�U�Y6�fu��w�5��)������w���o�I��0y�Ëo����$��˞���}Q��=�h��c.��o�$"{��{�QDG�k��>����z "�U�����g���s��>w�d����2"��e�&T�l���d'k7U��{�%��^=�9���n[�U�Ц��+���%{�|�_���,�g\�ؙ;���;��?w������yu{-O�h���|�����Ulz��%����=:�q��q/*�<�lBH�vSw�g��K�a�ݧ �\0�2{ ��;���\3y��>�����ސ���D$��h�2�t0�L槲rw%ݶ��A�sR��Q�u��Cq��aڂ��Sj�ۼ�������0����8�kWC��7x�/�-���&xv�5�8w�g���:w/U	v��T����D��1�2��It�8ul�9�pY�t�'e��Cf�lMڎ'��n��8OxrV+�r3�V�ҳ��c��=H�;��J�A,Ǯ��7,����� fP��Wgh���&����ڊ�8�+��K�y�`ut�]v����e�;��٭H��e'3����|=�EܵY�^��գߣ!+�,j���<��w<��[ݾ���9*Xy,[��]���L��B�Zd��a��ԭ�p5�^������t����B�]�_���|�S�^\��X�"�׫�W�����}u��Ѻ��N;�5�$�	/��Y�~~qWb�zk`m��F���;��9�6K�g\�9����n�clrV|����{v�s%O[�b�h���tbUEN:���5�:U�;�;7.��vr:譞�����e�tu�ru�\d�%�����'k�;x�*��m�O^tZ�t�$<=������a�n8uzJn;;�L�u5�n�ě�;��h���]	�v�P�d���nF��XGnH�K'&�۞$��t`=+��4�	�O].��W��6�m�8���/U\۠�n�]��7.�>/tr]���������=�֮C���;s ��iǋ'���oF�B��s��[�blkp���clF����p� s�t�;$��y��t�pu����Nݱp�ˍ[�&4�ހ�S-۷/����.p;�|q�<]�	�R�͞x�6т�{6��-���5F�{u�m�ܜc��Qq���4��uu�-�g�n� {��0)ƝfWW%c���Gm�x��U��J�Ew���[�ю�=uN�H�+��:��wla�r��=���u�kq��#s\���<� �ۨѹ�v�on�p[�^n<�H���{v7\ͻ;[�����a�W7<��":R^���n]��޹��`��"�v-�'guY�[�C�x��qZ� �܈%7A�<�-Ξ�pr=�<�C��\�۝ۈ;���`Ǘ�\-qڶ��G!�{g��N���M@��[���ݎv]�b3�,f�.��;u���^gٺ̽A�z;l�Vw�로�xˢ��]n �5kb���v7��`F�甙�:]��<;���ɍ���^�JTX�bh��%��[����6�u���G=��%ݓ��,o;��#�ێ�o]�nA��l7^��q˺#�<kFz�tt�N����[��JgŞŔ�m�TbH�Y��k�-t���`b֮�ka�7n0�{�n��,��8���9�H���v�8��ue��x�*SF۞64slq�%��Kc��۱���n4H.	�����vw
�����6��+><6���Pۥ�X�N�̚�Vn6��s�Mӷu��m�!F�L�KM��]����Αsm��z�η9�.PIa��1r������ST��a��8ⴙs벻�N�lR-'nx6|�h��]j��vŝ���ԝfz���;��'c]o8Ռ�K�u\PM�N�f�d)��=���q��v���z�by93t��u+�cgI�6��u9��q��(觲Y �=�:�v��km.<����h�m5����-s{W�.��p�z���t�<�Kv9���^yx�۶�-Y�kn=;tk���\N۳��!�mՎ޵e��Z;�!����Y�m��ɍ7#�N{\9���lm7-�%� X�صG� ���G�h؞h�ŷ<m�͵ŷ=��ֻ7��v�Cgcvd�'s���&�yһ���ĝ��$gBM�6��a'QR[�݋ڻ2�.��G	n�/m�nt���S��W 5Ϲc��`{<gu�+|����zA�V��w�[��l������c�l�L��4��d�����H^N:.�Q九[b����Ȼ��8��7c�GF��ik�[��=6{�]0�5�[kv���]uc�����N�bӄ�k({���_i��rs�n��%c�3���nM�ps�'dΞ7C�1t�=���ț�/C�M�l��$76�[jM�ŷ.-�n.���-�=�x%F6��Ψ]ӵ�댧&=�۷Lv���ۭ<���"ڷ)Ʈϔ�����Lv�g�ۮ7j�.ч�|�n��zY-����^u��i�cK�]��X�v]�;K���a���v��۝C��s�X�������m�`N<9���ΣP��9ƽ�9Yug���s)�8y�v�G7��Pv�۰����S��@k�f��;8��֤DX$t:�����|� ���\�p�&�/k6v�v�&;�qd��K��[Bpj��.�b����(�G^�qr����7\���;8���mv�9��Y׶D�;x�Nz�L]�۷e�ɭgՊ�;=;���nz=]n�<o��.v�ht����`���g��6��y�n�C��{n6ʯS����0�C��9؍I�⛃v�WV�5�����D����������s�����������ܓ��]��:�Rӕ�m��̋sn�9yc�v]�^��B�mmS��jt�����rO��Y�elME�d�S�Kg%��<��7/n�z��t���5������=�7{c:�˛��0۰h�K�^�˰M�������:����k���K�dN�x�Ob�v�v��V��]2��lT�����nSh��֧lr�xT}�9�DĻqt!D7`'d�k�\��m��6�7 ��էۮ����m�=�tm�닩�������6�2 �u,�ʳ֎����ێ�s��n!��m��xֺٰ��d"��^�(���w`c���ۇ�A��=pc'N�NƭӬ,�uclsb��8
#�A���scp n��<��K�m#ʰ��&67l��׉�n��V5�۩�̓�=�ʫ��u�Dݎ�m��1�7���0!�Q�	܈X�@����Ю�Ɯl{��v;e.)��Dn�`�<ֲ�uΦ�G�;�6;[zU�y�u�q��f��f���n\�3�ݭ���g#�ۚ 㝻m6���;cS�=�]n9L�>x�O/���qӻ���\z{;�eK�������қ���-@�����Ѽd�Ok�y!�!���l��X9{� �;�ܜvt���yΡ;��A*�p�0�Ϟ��R;m�M��[�Ý��C[�z��э��LcA�8���1��2���,kR�k[�
Wny�/`l�{�Lڳ�ִ1���Rd�]cC�V���v���t�����t�gX^���{&�ͧ�=v�oiS�s�9;;�;\X���׌�r�����;X�X�C�z�����]m\v��c���3t-��{w2�m�q����l��/]õ�n�N���֠�]��[(�w]n�����9���v.��/3��������ԛq���s��s�mzu�.CwB�[(��Y|�Y�ݮ�^�9m����Oq�6��	Ŕ���9�bp���J�N�u'�q����ϔ�*�k)�T���˦��
[phN�Ǝc�\��rU��� �n����Q/g�u�\�0�=�ǩ(��P��ٶ��:�%����M=��WBuZ:�v�z/X^�Աq�,�y����Oa�7.8aG<�X�ˍk,������΅�5�;��q��OZ+�J{o�컩7Pq���@�^Sp,y��d��Smv2Qγ�;a�m��l-�fh۞�����oP�r��h�ӎ���v]ǃP�\�K�v�#��G��`C�L�s�mk��6�;$�1�I;��xX헮�n9�a �Kv�vKy�<qh��R��v��sy�Okٹ��E�Ϛμ	��;d���r�nɭ��5Q\0jV���ꇭ��qs6An2v�3��Z\Y�C</j�M��-��\W5n��c1������<#[�p���8q�v�M�.^���,ܙ���cd�q�s鐶J'n7&�]���]���Z�q�{�Ahy��jK���<\t�p6�-��\l]�����g�+���=S�p7`N���^ܹhz�l�.'����R;t��'����U+���56;V�[V�r�6yH8x[�6'�v35un1�t���v�u���k��vmp�͞���^��>��n�;�]tsq�7<��P9:�D�\W駵��m�ų]pq�=s��rgS�l��wZ��8^�9�q��kE�ǊN�tI�v����;�[��+�k�8�z�.dT�cv���ax*�Ȩ����Q�y��=�8�ocp�w=�L�V��۞����/7��=O=��dγn��l��t.���)����C�a��I�R��"��z��Z�8�F�c:ۍ�Ʌ�M	�<Xq��wj��oV��ŉ�.��X}��`5� mq�����:��ƭ�ɤE����z5��q����,�KJ�.H֮v�$�׷���7c\�^7j�m��5���5vS�p+����Mn�\�G]m��3����p�J�����W�v��ٵ���rY�ٌ�]h[����vMd�'t	��n�v�І�v�a����^]�Sq�:�9����{s\�lp�C���n�]W=��mݽٻKn�r���N,�d=��pn;�ss��Az�:���q�	�6]��ݙ���ݺ�ci-7c��]�.�+��'b��<�;$��3�iݪX�T�x^��͸ϝes�ܷWm�p1�&�e�q�Yd%�{�n��b�i���Wcmԃݹ�du��싹�������l�V��d�G�Zsu�q�u>�ܛ�8�.9���v���q���Q��h�k�rd�������m��Wv�1�=��LӃ�GV��1���}�	��5��<[�3@l�^����쭮i7`K��q�z�������=U.55�Ӏ�	�'P�=2Ӹ�*	��9n)�y&�6M��湎q>^�ˬpSqMة�i�윽��������h�qMm��Q����c�����8�e4l�u\u]����Z�[uk��J�n`kڋV@�qM������nzYCl��k���Q����x��r[v��o`껲<v����D���py|d�ewm�d"w7^ۃj��M���lun�=�y�2�V8JJn6�8�y��Ԝ�nm��[-i�\u8Y�ZC7X�soc�Y�8�����C�c��� y�[p��N�����bv-K�S��N�<���)�!�n!Yu�껌t�G�[{@	[�1�V��e���b��]%��vn�����P���.�quq��xb�c��B�سӒ�͵�y��g����b��+���o|>{�߷y�
#�!ΎC�t�Bt $�nZt9Kn�lpQ�t�)'s�8q�1Pۦk,���#���i����	!��I�ø
B�.F�v��t� \�%�����Q���AbV����8s2C���$w8���t���l���2� �Kk6�,��VZ\��H8�8'HD@\Jp֖n��r�ga� �A Q5�A��!N!�s��p9Cm8I�v�`�	#�ڴ�	�H��p�8I�t�"�(B�D�8��	qӸ�Q9��� "�t��e���9N[VH��2k�W����_>/�v���9�wI���IC�|@���x���m��٭��JX�\�<�m�q%�����mn�&�\n�z�m�r��#��]i��Z�!�K���V.ػ�e��k�\��s��7�iۘ3�\a��v� ��mۜ��%�Y���=hg%�Q��;Jc�]���V��5�`��s��#u�n�q���"ỷ7�>��5nu=c�˧�79l\�6B��p�#ϱgf��M�K�@m��;ko�v�.����ś�=hrz7<��G烰��f�p�ݦN��\�+�F��O=��m�ݱ��ҷ�m�k�:���|�$��wns�����k��&n��tbxޣk<$���=�M=d�冋��B:�.���&��kz�֊y�hÛD;&�P����SY���N�k���|�:y{��WD��"ƞ9��<fԇ�r�1۴t{��V��gF�,�L�tlG,�����ƶ��Iܸ�k�r�<�E;�֣�Z�vym��^K�����'��Rs�m��������J&#��x��k���^��vJ���˺EJ����=��]�f]�7��e:Ź8�A �3��;�%ùںۗ�koTdrg�k�޺)M\�������p�����D��ro`���M��s�1Wt����{�b_cM5`��n�	�wXx�x���v���N�\Mܲ���.G�msq�r�<��g���Z;�TJT���.v��{C��LV]�n�oi�Cny=pn�;�7[onʊ�;���<k9���>Y8w�lr�[��{sɒu�;�\E�lmLs�:;����Wi;\�����#���|�kN.��Lu�<&�h��7:�˭��Œ�l;�:G���6z��]�`ڸĹJ=��8欙�7Zݓ�F���[M�/A������۰9-^V�헌����^S��=�J����9���^��CV�n)�q���^��n��"uf�{���C��܆�v�����y��{�&ݓ*/oe���1˸y9�yG��6��v�la�V���=���q�{Ɂ8�w�;�웳�q�.¼�rm¸<�y��&L����N<;�6���6y^ݔ��9�s���.Gn�.���oc)�C�O��s�*��ύ���y�2`��e���n�<���㼱��{�jy��z����o�����r8�lU�C���7���Zd�n���v�j�f���ϕ�:g���05I�ADf׽VH&�o]��Oe^a������y�|zU*63�r�w��d䅲�mRBǥ�y�M��.ud��w����ȹI�1\�Ē��"�!�:�H��xA���UFd�㰄�%3�	4s�oĀH'w�''�����<u�M�ֵ4���Em��%Q��{B� ��<���Ȼ�������8���H$�^���������a��n�sGSX��[d�Q;+��;Z��k��3�U��-��ѩ�iOL��u��}??QT3yn���Fj�$��dO�{`�U��ڹ�����~��`���Ɂ��I�7D���fj�fy<|x�di"9�Fqժ�4C�X�1�3]/jj^�P�\=h�̍6�
��Xg[:uW]���J>�`l�͸��򺁋�$ͬC"l���A$����=�G\>����(�$�
�E���g�=;� �H��MNpչ}���N���|&��s��]}3t-��j,�9��o&�C��w7� �[S���+a ��
���Z	W��s*n�Sܞ-H�I!�����g�Q��aa9FnHٙ�#�k��	
{;gzoƣ#&���r7�5
D����J��"��X�ۻv1j��9�q�����R6��P���V�%�k����FKǃ	gzl�峹������=7�4�ݜ�f$�y��d 9~��^`�lm�ZZ�QS� O��Y��}s;-��d�o���;���ֲ��4n$��S�� �m�` 5�_U��W����'�כ�o��|b��Q�^����J>հ��C׺p�zzb碚�ۥ����+*U55Y�mi�#gq`���H��cPD��j��3���xn���� �5ݞ�	�>؝S`�H/zxh�"W4N���O��Y�����B�k���CK���M��y�K���c���"��;;�=��l�H/~�лUփ�Ǽ�oո�����U�-���7�x���c^�8�ҧeMuJآ#����~�����UTfI|
in`>:g\� �{z���ǣt]��ٗ~�����ۡ{@IB�	Hk�������y���D�u��Fw��A����#؃�wu0�v��w�?s3��V��V=f�M&��O\	7�LM��;w��H�Sd���Oh{ݻ:���U	t�ߺ�]�V@ٳj6���m͂$n�	پx�����et��1�ӹ�����a���7�Eeݟg�G'�g�s�Z���c�z�坔}�,f��s�rEߞ,N1�?n���S�o߀��xp��$�5BQ����A�w��*����df�V�M��;9t4��}y�L��CP=:��GLL`�Yy��s�� ��c��ͬY���O*6�p������>����k�JS�o2i6���;;��2o��u��K��
�X˜ذO�o�����;��vZUm�F�w���,�3� ������A����Iɾ��A�k��d2;�˶;�ݴuY[-f�3�v���|�a$�#0E�����'z'�k�p	#&��yfa����ɪ�����.:�u]�|^�؂H$)�ـ�O��(q�y0��-8�� �������vuI]�����{|xJ,Y܅w$���7�H%N�fA1���`��_x���3�̏L*�*��:ªq�j�����]㔓Q-�n�j�)��Y��dݥ�����elL��o�>�d;4#W
� �#�e�:@�ݟmy����ǥ�b��j�ֈ����vs�˗V�9qm\�8������u��6���� F�]��:ж�v�F�lE��3��r�Ym8]θ�S�s�����}��=oi�Q[)���ݷ9븝BDro`s[�3��V^8�m���k������g۞j3��m.ܑ������7[:�뷩��Y��wj�=WLq��ܻ���۷Q*� ���������q�Ɍf5���$P�h���N�GN���8�����U\.;[|S�W �>�s �I �7QG�[7 ���{ss� ��b��$�<�X5#�)v���x�O雷����UTfI�-.��O�X�e�>^����=&�������o�I�K�Wѻh것F,����Nvz��4� �Vf{$�J,�Cޞif0���C'k�s	^�!V��3O\��o潾Ohw]��S7pm@�T���Y��J��6 ���6�>y�yT��6*�b�x�A�W<9::��v��^8�OhqZEb$U�T�lR������zuI]��	|��wƛO�o�M�I/z�ߍ��wgbdD�W<��ޛ��`J��(&a���ir�u3����n����N�u���w�t����A�N'�30��C�.��������f�H�n�����%ŷ>�ۍ�g'"����2����I>q;�d�|oOg�D�f���n]����	mrҩ%��6�l�O�.�pH�x'��D�@x)����ͮ�~�M���Ohj�]�R���mu$�x�KX�Impl�\(DG�$x�{zx��=�p}ϗ,�'���}Ѿ�-p��Nڊ�S-f����!4��`�m�Qnai�R>�C���$�ޗ~��X��8�L�l�#�"�� k�7<���w!�0k��n՞y�/=Ͷ��������#��;i���/�m�|�pA$�V<�9k|L���}6I>8������꒻ev�����]��{���]�+y�"Q���'ĂG7L���X�:'7y�ݣ��g�	l`���0����$��,�@,�oE��A��5Ƞg�x;�;���ا6���d�-i����t�5/}��Y�_x(�6��uX�g�^��~ǡƷ۵�I�{�M��}��#���s��uw9B[]��B������t�@�ɡ�(Q�sf� �w�$�ѵ�ccSFI�6�"A�R���-KQ5U4*�ԓ��ږ��Iӵ�e97��%c�*�a�j�fL��W��-Uw.�ݵb�x�N�M���j|��||��|��_.��&�l�Ny:In��������k<��fhM�n{  |*�X�U�Q׼T@}&�Àz��>�[�HHP+��}�7馵���I��ֈ> �Vvg�,���U@�E������pC�J���K���{4���V ��)n�G���=�I>J�`�7餛�:�w�Q�Un�Y����~��7b�a�W���K=��	�oĀH/zZ�}Ʊ��+8D����"�S��٪�|#jF��-BN\��Ql�I���T<�<�@"q{���'�!���Pf*�gn#=N�m��g��o��O˹�Ierڤ��_.��5�O���?d�!�C�4!@W�� �3�W������w_O�/��پ�/cb�gѹ�-���.U�J�1֔
�PThLO�>>�q���o�QԒA-`�%���
*��� ���͘޹;%C��G�m_fI�4��dZ:���[-f�Ns�4�����oq��y�}�ē�JE�GoK�K�xz��M�5Ͷ��o�����r̅�6I'9OX�	>rP��i�|Ҷ�}7{>���wC\��:���It��'v-u��d�e�J.�l'�W$�կ1�h�Z�T5��o����Df����`^�� g�^��E����$Dn�߉����x��y���*�I��%����i!Q��;<���T�L��t{"2+N>�l�̍�x���L�j��9��<8Guvn,8�Ӛ��Dz�m�^���Ɓ"'u'9��^}�s����]��x؈ݶIx��G�ql��N�n@�=�v��sPz{���0�7'nYへw�N1cn�@`nӝ;n�;\�:;���ONW�f�9�6�WG��r�X��:�׬�{:M�6�p3W<O�Z�#����I�|�U�[�ɬ�y�r�4�g���q�.u��p8����c\L�qoYw��X�&�::/)��ݷ7�;��>9��>�;�Z!�S��b�gW=�HZKj�¯�'�4�m�}���$ծ��vͦ򤌵0���>�šu�~�GRI��L^�&3���q�W9�I�'w���	]Z�	0dK}������\�>�-n�ȥ�-c�9{c�? '������O�(���OhM7�=w��������Wk�൝D�D����=�A ��׃W����ݑ�Ѻ��鼦�(����I���]�����1����n���Wd���lI�[ـ������'��{M��Z��WXD�	-�а��`�>$����4Y2����/�?�}ͯ�����0Ʒ'��	kU�!�}V
'�V6T!��h�9��I�u�0���j&(��H�3,���-�n5�GL-I�ؗQ�Hb�k#X�ѽ���܋f�4.�^�o^�6οZ�E5��Y8�w�? {��RK`� ��V��S��*	��y:��|Ouof;]6	�j���Y�J�z{Ikz9�)m��c*y��Ko	N�M�	�Me��q}�r�ţ�������������er9`�LYUӋY�:�C+I �\� ��s~ �}/z��ugs'j�fA��0���{;�M��f`Վ�I]VG��3�I���S�.f���X�[���f|Hq���I�z�첄\�ڨd�>�Tj��n�\�x�xA� x���"�I�8�C���O�T''�{�|tN��c��[����~{��o��>�����''P�uW����$���m��Z�(�(��w����Fo�渊3�jsliGk��>#u��f�Kx�޷��Ă��MISS"d�P��;s`J�t,s�����LD	��ޛ�9��瞥�k�)�/aٚOsu�j����j�B��5�U�Ӻ^}�=�}���1�/ۋ7�m�i�=�����N1M�=*�C+q�F<�vzI(8���:M:���/jgw��E��O����z��W!���:-Un���a��e�f�n�D����U{7�	M��;wy��������Z��=�N����^��;FL ��V��C����k|wL��קW;-��q<=�����fͻrm�5�ܻx[0����S���__<���׸e��we?��͕4&O*:������*�W�U���Eړ޹�?�ε��L�ȽZh#5�@�Y��P�0b.�_���6�ԁ�x����l^�v&�jF0�&��.�����1�G7(�jh×����a�9��9�Q�gw_��ü�/;�g�����G�&�yY$;Y=��&6`ﻉ�gM��xPs�&b�z�/�H��M�>d�`�vH���"|z���ӫwo����~~�H}$D�1�$��cW�y#��.3: 5�j�s}ݪ���^:ޤ�x�rN[�E.u��!f����ڗ�[�;��.�:.2�A�|�8�`��|o�Rle}�s�l9=�w�~�u��'&���o#�N|�O��g�8����il[�L�U��K]�;ߎ�g�+�C��������������T�3״�ma�.Y����5�o��3�9g���M@��=wP���9�N�v���ld��j�`䯼�B="����wsM<�6^��%k���@�0�9	�숹E�8(��H���,I.H�줬�V�b%�u�,���I6܋�M���vc�-�"Hcmah�N��Nv�#l#��ۢ�RH�mr��Ee�vY�tm�4�H��.ɚt��p�ċ46��$(��QvFS��v�	�����!ΑN�Պ\E�vv��-�
me�Prgf�ͷXBu��Gf����w$Fݨ�)qͲ��G$���M�[YNs��@6��!¢�"�f�V�B:q@��8�6�nQD�eq��5��֐f�ݤ\M�ݔ،+(6�������D8�N�N��Qӓ4r&�۰�,�	�M�q9̛t��I�f��e�A���`�S��L���^�g[;Y��������C��QKRH�X&}������U»k���w�~$I��Y �����OA��c���8�`�p4Tљ���,r�X�~����Y��kp��]6I�����=��l�x�uy�v�~����eӖ�ܗx���8*�,���`�[G]DQ��V�3��F�����>���E�Aƺ��I
{^
�2X��#[9]��m�����}ɺ`�R�[ahTrk�I܋�ouS�$�ز���|A�e��M����n7!`��7� Z��]4ߦ��Ɠi���76��3di>9������KQ65K`��ե�oS[�s�ի�ޓF�*�>�GN�fq��u�&��A��>5��k���^NH<��x�8ƭ����#�p���.��,F�T�8��v�U���G50Ay����c�����V��� �o�a	"�Gt�hԳ=�t�t�Q�k�I��3c�0~������QC���?��{>6i:p�}D�����%t�y��۷b��X��p]��@��&��g{��u���-g��2�&�`�x0�b(�S�qQC�]i �S�>�&�ĊH,��&C��`���.��l܉��@�O��X0���d�~�U�,�3=ڰ�,؝R�[ah�����O�"�'vg��C�g�1c[������co�o�I��Y���u�P��>O�`e��#Mf_�s�H3 �t������JvD���ss	B�MI���,tml��.t �7k��x�:yna ��uM�|H/yՔ����q��1�{��R�w�X{��m��c����1]����C1z�o�%ʟ�jd�s9ݖk��l�;\_�� cpw�����.��z����>EK͸h�m�qr���`�;tP���]���c��y�(v���ny�(���X�)�����mքm�kgcw\}qu�a�X��QK�8�#��+3���<m�m�n5����:N�������}g����ں�v0�t������ۅ�Vn�,�q���O*��f�8w�<����_7�e�˔�yy��;V�b��A��^C����ntc������^�u�w��~M�쥐������5�5Ȱ	��/`�Su|)3k�mof6���4�ۊ��n��k4���]xi�Q@�'�A�7��z'T�$��u`�k�:)��w�K]����T�U2oE�7���]W�A ���9�=�ޒtΩ�	$��VH�ڍ�h�5h)-)0������3��&��<;�6$���X'�g�؎��W���F�M7�,�X���tf'�g��m����}� ��#�T:sd�w[�Y��z����'$��5ƽ ��e�"%I���۞��%:��uw:ղ� ��YT��)����i�QDɡ�#j��� �ՒF�k�T��LJ��$�SĀIo���$����DϺ���_�-G�ە�_>�}۫�t��<�CY��f��͇���#���������UÙf�s���+pF���� K-��ą�}~�vs��>m9�l߳�ө�������-�֐A�]��đ�����`����� �qt��<F���$u,�&�����f�l��]�e�0+7�G� ��s	���OD�ޓ����{�~$������6�]!c��Z����,m��oTٽU��ؐD�e3d�{�	/zoǔ�E.ݭ\��@�D��T*��]v��s��Ks�v�u�ɋ�Ll,�X�H4���
�n���1FQ�C�%\|yR��8��n8X��ⴝ};b��=�0�I�H��Dɠ�\�)��ڮ���;m]�t㊞��ћ�`��WOV��S9��W{�M��!%.�������k� ����}Zcrrھ~�`���=�ݘ�ͬ��L�>�dt������Vӆ*�a���d��3[rcj)�3��Ω1hR�,�V���V��J��y���<������MJ��%ONs�n
��]��O�f��A����Ϟ��wg>9���>o�滑KZ,�J�[$/�׃ ��~�K������dw�$���6	�'���2�n�&�[����g%�e�E��<��9�c��Ѵqm�iv}��0$&�u���a��P��*���;;���$�z��H$�q�B����9��p�쟀�C�n9엁�((,����'�	n�$筮B쾬�$�o�ݽ=b=6�+0bc{kB���􉚂dL��W6	�].� �(b�����h9kxI��k�ݽ,ߨ'�H�555G0�J���ב;��Fӑ`����1�~����/^��_��[���+��}:-aV��B=�~;G�����ۋ�O�Z�X�p{�l�}���H)�6=�����?o���6%�7_<�����������C&��U&�g��r�{>ט3l��tT	7����"��=b'{^f@�^Q�o�ExaVwfn#9�v5�vN�-ճ��9T�X��ۇ�1�8����;���d��g��f�o|��	y���������d�r�~��1
�IQ-%�I;��x�?��@��f�㖧��}L߉�#y���?��Z�߬�rz��7P8PX�#�yA$Գ0�E�Zc"{k.�� �R��	 o5���%�5�5ș4/�U̇�UJFne��>'���݈ ��ڼ$�{ӑa���{2��ٻ������Q'u!'�軤(w��~���z8UX�@���d�����ޛ�zn�f�Tp��$>���V�K,��8�bw~�7)9�]��J��'72��B�v,3>ml�55�z��X�C�u�61M#��_+�YDŴ��M�e�;�x���[i��uRc���on;����Ԫ���mq����L���g<eM��o�-r�wh���V(�p�ەNv�Om�ܒB��@��.2�_����h��1wl��y�n�����qϡ�=�������nL:i6���K�e�6�v�e�qU���q���;����������]vx�9�=i���qֹ��=�F��ۃ�8�7`Λ�� 8	���}A7Jo���߻��6�
��I�`�Wn` �ћ�`�#Lun]��[�<8 ��Y3 ��|`ԁQ�Y�l���_��}�ƾZ��=��y�C7�6H ���r�o���z�hV�ʤ��U'��}�7����5�KZ�Lc��>)Wm���7��1�	K���">OO�����H?N�k�${{��W�����(�w����ɚ�dH�;��	�ίŦk˛:� +]ل�f��O�=��i�X�ZWKu��gѲ�)HꖉHfȼܭ;u�c[zV0L�Tn�:F�kK��SR�(j�
ћY�0�t޹�I>=��/Ǹ?��VK�S��� �w�`q���"h�S34�]�d�f��*����)�����^��X|=q;���ÄF�n����'1�Dc�夵��|��&�����K��G�͐�/g_s? $Ϸ�_�����V�s�ҷ��=z�Q�g�|�_�eo�MH��Č�NP�|y.����S����A��|>$t^��I ��cgj4E5SBKKeRs���^����<w��m���u��;+;�痆�M8��G/%�q��19A�f'랺m6��3��>��u�v����[6 ��V|vVvO��׃K�tf�|a �HI"�ĺG���ۭ���/�|��"E�Ւ%u�P�%V(Ej+�ߗ}��I5%:!4{+�r��Ǿ�-��'�ٞ7sf�qV�Cn�	llm��$qw]6���m
�e�\^�����ܓ~ʃ�wnp�Nwu� �O�V�a$)����s[ݸ��5�}"z��ԭ�$���y�� ������ݠ��1���lW�#T��Ss����s��o��UAh��xf��۽�-�f{���Ljm}����B��7<1����i��3<���\rj@�зV$6A;��^��Dp�����'5mY$�uV��I��uƌ�fk�9�|�'�t�gi��ieVZZ��v�0��GjT3W�콘��K1�y^� ���Ɉ��O$������n�'*�b��h�˷���+��l]^Ӽ䕪9\��5�����V�5��o=l��j��C����9]�ˮ8�k�����k��"k�3Q1$M{��h>��Ѯ$�-d���	$�Y��۽W�L�|D�b��U�M����֢�	�=k�0e����	�񂾂���:A]j����J��'�K[�Ϲ�~=�a�۸�����Ń<N��_�>;�Չ]�Щ�t��1��h�ٕ��+C���Q{����qM�膩�+h[/����<�����wݩ�%���f�;�}ܷ�%!���	$�h��}���6}�v��jT�Z�B��a�_U�	 �˨4�3�jnr��\	��� $����.�/I�Ɏ<���_�%J�U$�Z��Q; ���8�cz�.9!'0q:8���r/�~�~}��=B�5S\iv<Ivj�$�S�`�`�;
vx�s0��kx�ٽVJ�A��*��3�uY'#/k�®]מ$����$���d��|z����h��^�L�A3�^n���|^�_�Ps��w���'��|{7�� ��B����vR�K^/��s]��*��OxJ�MR�d�O�>�d�F��ɸݝ&���i�;�]7�ȝ�GF�%��O�x����6[*�����̝� �ZN�A#V�f��&{:ov�ۗ'Ǽ���=�fi��n���y/Fs����Gk���#t�Y&���_ꟺ�������j]��WH�Ã���;f�ں	�i
b������]��=�s��ԅso�gޚzTRV�Q����J�,�V�.=cu�U��6b)#��2E'���u%�Fu-��*��(��t�aF�ʤ�j!�E�fӀ��D�؊�m��gV�:C�4�;�
�x83�<W�E�i�}�O����~M�������y�~�Y2�ʊ�p6P�%]�SuUs+��Bg��]�ς�,����o���^���n�������A�{n���g;������,p��kkܶ���h����;�ɦ����ї�{W�3�ܢ}ؽ_�l�BpM��{{V�q�=wG־�Q��2�ݙ�ޞ�Q��'LE��n��&I��jj�Ҹv;��m����q�H��
-3{�ٹ��q�{��f�nN�([꬇��l�j/`��Zr//vad;�"���ˁ76�<�qP��^&�7�4 ���A�����/l�ߤ��i����I����.ųǡ�}���ýJ�0�S��x{���{��.y��1�{s�x�\�>Z��û}�j����L�0���u�=c�&�����J8�g������S��O#�w{f��fѻv ^�UmK����;Q���;�{��l�6�8|��K�{VY.E��]��{ؠ��l�J�+�ɞ	�>̿'�_w�\P�_}��M�II9�������ݹ��I	%$v�p.RI	��8�9Y� ��
������e�,Й`η���ԓkP�6Ȏq��m�m�]�e8:.���9�a6;8$����NPr9H (
�裳��6��Z%9`R	�$ G-��u���:L�#��	��9ԒDڷ ';;q�#��g
AQ�T@���I9�;5�֭	��'m�9[hfr$"B�+n�%rs�-b HI�:B:D2�����)9)K�����n���ܜ	(��:qR,�B����@!.�ܞڂ���!
8Ok �.)ŵd���YۛX�%$#�Z�<��>ߓ�7��s�	�t�g<�����Y�Gh��8�۵=���]B��KC�I'����vѓ��v�{+y�X��G�x���s.�{Og�=xG�WoA8�H[��-�96����l=m�<H�������lb荀7q]���\���P��	���m�ϓ�l+�Sk�O�������z�ܚ�ln�y�_;�>�9�P;�a{6e8���GJ=P���l'�Y�g�/Olw\���W���2k<0e�m�ӝ�c=>����g:'���q�g�<�I�ۤ{wc6x���A���s�ץ6��]s!v[�뮹�㎷	w��#w:�n�����7�Mu�m����n.�\ցpv*��5���C+�[{3�Õ7�r-6s��Ÿ6�Oi7=L����Wo7Z�ю^�Tm����Q��A	�q>m���\���^4"��qE�6�{�eݝu�eW��]�N�⃷g�Ii�����yWm��=o8�n�&��c�8.�z��cK���E�=�z�;z����7G����mÕ#���W{:�n�f�okkv�ܷ*�[�Cֈ�V8��Ӣ��c��/g�q��N�ܻy�un+nV�n۝=���n�wU[�u�{��v�e�Q��yڹ�kuj��:���n��sэnڝ�r�zN�� ��۞,�O��a�(����c�@k�BPi�>.7p��]Zu�u]��k�;q͖����p�.��>�񛃔�	tv8�.Z
8NDz��ۮ�P�=����W=�����]���;v<tm�k��s�ݎâ�cF�mɺ7Ż���!N��u֛&��V�{\���kz�n���wk<�4eu�j��r-���n6���И%9A㎳Ӈ�V�R��^��lm��K͌�۴;]�.�;n.��t��{=�3�v��㵱����p{C/=v��#���u���N��#�dD�l��n����\��N�;�Ѵ�R/DI[1��۱wHuGn\�Pl�p���Sv]p\��Y#��h�=�����x�Ʋd��bA���X5���<�5ct�؄\����S�L�
�k�cmQ/PL緬n��{Sּ���c�n�+z�'�+�A�pٌq�;���0V��l�n7dۮn����vC���T���v�Ơ�7&ݶ�*l��0�vm��v�RB;'�㋻Q�x��:����e�vH��؃��f�s�`��^��Gc��q�p��z�;�糘��N�՛�n\�݊Ӳ��(�u��;Gn^-��h�?w����d���+��I����ֺ�I j���l*uSx#&�P�(�a|�� W>�'gj'����SUSB�X���B�n��>!6�X��o�`.r��6�^��a��
"b�D
�`��g��X$���#4h�b�+A �����	ŷـ���1^���g�E��w\*1T�S�O�v��I$�{o0|	�*��snÍ�@3<����Ǥ$��'R���� e�rx>�d��X��5]B� ����ʯ��i\=ߗ�v	:2�Tm�y@47\���q�䝹T�.D6�r���H�پu?u�#�%�xŔ,-�c �r�;i��Q���{�M���������9�BY*�SY�/�^����ym�d���
ʑ���nWfG}�|iyV$K�n�Q�ʴ^�	�N�����Ҧ��N�e��lg����N��q8�F4Kq������7˫�I�{}��	�>Ud����y���\�J�喷�"zv�pH���4jj(G+v�U�	ɳt6^i��λ��N��c��VHLn�1S"P0Fa�Υ�Ss�P�_D:��0��ObT,A]�T�l��7�D���ՙk���q$��^2+��V��A{ά;^:[�BsP���3	�!F%6	��޺O���{8����^6x�QO����x!J��A�ۅ�������`[�Y-�������U���5E�S���ӍM�I�+��_�9c���9Q[c6���Jlu?i�#�%���=��[����yz0O�1)�I><���M�d]�\*�:g{�'�#���e����Kw�_7� K��A����`��z�9n��y�2El���1�SWX$N*ݨ�.��"�Ʊ�6�'P�����乺�[&��N���\��N��	�mO�x{�êk9����{�M�׻��I6�M�mE)
��j)��>�A��@�v >��  C\���4 ���a��e�"�b�&`��D\�$
۽��M����K�X �}��`����s��J�����8��y�BhLl��R�u��qϵ]vT�%ۮ�ksWkaceR&��k�\��P��w�4Odm�� ����I>��}�r�C�ի���S�/�w޺n���2UHV����0�+Tddob����� G��3�I���܃}� �GŒp�ARM�|����r�� ��)l�O.��$�y���
�}�	����K�yy��s����14	.�U��|M=��	�������W[��D�VE�QCN���q��[��D��u���u挿���&��/l6ׇ(��f*�q'[�Ƿx��Q��pT��#�y ��{�݅?O�SMIZAj)��} �0g��Y<��:X{I�\E��[}�I'����j�_��dw��lmG�Z�Tu5UM��B+�;m��J�:��z3��8Փ�P��sk~�8Y�M�O���A$�k0�I�mY���C1r�.���s��bm?W�������VוUh#cM�1^��Ĵ�6���}Ko�	�z�hY�1թ:'��;�}X�O՚�-#u!&��A�~�� �<ANWn,,�Mg[�q��D��舸"&������|��קon^�>�5�H;�6><�yث�.M_�w6��3%P5SUB�`�ٶ�x����F���M�W�]s�HQkf�O����؂/�fk��nB�6iI�Ug��-�S�k�T�W�p��5�.2&Ғq��:
�G'"2A3j���j5,F9H�֣��s&�W��P�>}��Hv�Z��&��Y{<=Pm#l���{f�F<�V���eKb��ɠ^�:��s�l�{��evr�h|i�L=,��#��[�:���`�p�W= �ϛ.��J𙻎^����3'Z{r�nN�cg#��W�y�C0�:�^������^(J�!-��Y�ss�n-<����U�%��@�ob陣l1�6��6�����d^ۜ�ַ7[��a��]r��ӗ>˛�֌V�mktn����&͐��m�8�\��
���i=���ƛO�\��͂Io�����ͩ�6lBw���O�-�.yo|"+�c���|?��&����/e�o�I�!Ž�~#�OX�|lc���&	=GM1&��L�<U��}.�|�!�e��LoLslx�o�u�i6�{��$;$�X9-y�7���Z��UY�)l�|O��wS6	d|����_���
������k�Yua ��@��ld���U�~�����ɧ��͂I�\��㖯�<Y�uW��3��ShU��I~)U�Sv��.��K����l��ѵl���1��L�_b����
��Y��lA><���$��Y}����[��eU�%��������2Vi�ʔL����Igf
��:i��N%�kB�����:U�o�'\]l%TH�qz ���|�(��}�>�<��9F���two�Ŧ^�O$�!^��O`��_$Y^�����-ɑ��M�G1���LёRLny���a�lUܭ����I>�b<}�/�<H}�k��
R��[��;��-=��m�i���$��/�	��R�"	/�����Y��j�^9�T$��'���1��9M���$�31٠���"�+k:�|:3���Q]��TއU{
 �6$=��<m`�]��q�ώ;!��.ݍsŃ��i�^�"�M�w�΍�2�����ٚ�mg�{X�$��7�8�V���znQ	j����\$&7l�� �g�g���1G>��mU>���s1�;�Ag9M�@5��M���޵����7\N�Z�K�{�v{	'�%7�I�p*4�a��*�w_Z����U���rӏV��}o���j�(`f�S˪��=��R��>�5���-��8n���5s������g�O�*ǃ���lct�h�D��b/<z�y	�֚�3Q�A�y���	1)�H��ΐ�C��c 3i��'h�+�&�@"h�p���I'K��٣��r�A�{�0��J@o��lE#b�(���\�Di�D�b����nF7�[��<ǷWoL���V��>#Y����$��a�������I#�W���Gf��=Τ�3Ă�56O��&n�� Ԉ�&�m�������^L'���;FK�Jl�I���Y���Xc�
����Y\I�,�� �f��&�~�'��o~֬f���]w���H�lI��Z��ۛTD"���٤�/=�\j�'���L�6A�N�~��D&�8o�A���-RMF+��c&�����Z�2 %�����-�f��$�z�ֵ��n��Iݻx�ߒ�g�f�>�,���1J呕�f$��~�M��˜ŝ���9��/�1�$���������vt�����u�������EQ<��=շ=����������H��c��p�QR�S�����<�Ě5 ��~�"��аF*α*γ�{�U���	$��`+���B"D������n�etx�̟ KK���N*��'Ǖ��]����w��8���b�@��jI����>$W��	&4ފ���'O�s�1Vu�	��1&0MMU
��Y�#9�9̦��'��F�:�'U��q�٠a�wJ � ��VZ\�w"�Q»4�o;�cm?<�%���c�G1���9Nœ�Z�y��\O�qOe0������Er���g`��������-�`��T,(Y��#}V}����������5̩��o��f�k�I!f�T��u*�4�2p�gg�[�v1^7����v��^�^ڄ���^��5��j@�tcn��۳�6]����Jї�	�lu�M�c��{su��7��Oy��h ���-�:���D������SF��O=H��O7n���\:��Um�X;7����k�9�:�vؗ���M�1F��8���Gr�7�C��;�޷+�̖�	[��4��kv�ù7:{��b�ۥ�5�9sv͝m�w~�{��	\�B9��7�զ�����L8�����b�l�������=n�d�[���~Ǵu_�EFܭ�x�ji&�֥U��9�P^$��� x�)�@0����f�(�/�}��C�Hn�p-C�yV� ��H�⻬g(��{��oXDOVa �S~$s�lA�1"*������^T�����@���� �E�6A:�Qw���*{t�bZ���!I��{X �}���M������0
/��$o>���vȞ?[�?��7qv��/*�0N]\o���:Qŗ��b�oK��w�]����:8^f2u(��<�M���&�@o����j<���!���1�w�$�{Ov�o��]�� �X�{�y�F��z\m��ǭUdz���^E�G��Y��o���K3;���Ml�Ә�Y�9����Ǜ�k����Y���<�f;雒v�a��׼�:�m�>d�u!	%�����7M�UQ�?rM ���1(02>������f����{G���Tm��gǡ��� ��=� ]�vL��.s{�d� ���T`߻=��e��z�12�y��z���'R������3�	$�zk��b@/{��b 6k~�{�׾�'���z�Is���UK�^�N�@ ٭�f��S����n�,��4�����db���3 ���z�t�������ښċ����.�njz���(�ݞmG1��D�c�QY���#:���d�znF߾�Ӹ���sy���o}2�!��Q���Ok o\{�D�(�]���צ`OjN�TWL�}���&���oӺ3�of��X /o��L���k�x�Vn�qoM��]�K�ޛő�:o91` .-�K��۹��r)wFu!��3o_�?��+����t^ 
�^��y�{�[e���ꛋ�w�h��c�/O.Χ��i���P�6���l�.�'a���_{ԃH�D�-���9
s���{�4�^��b�
xp�>��nBGHst^��t��ҠH�2�jSڣ��=&�N��m~+�[������cV}�a�`��Q]5����iF��W�k͉��c�<���x����4_.#���"���ײ ���S+�ݻ���}.��j(�Df��7�yY����<��\J�1�sO&l��f)�e�ca-���8��x���7;$J�0,������8F�7�N���a^{��ڸ��(mrlǽ�D.`3d���]n��_�>qԷ���kջ`T��I�3Ui˦�:�.�n��:�	����w�{��F��$p�+D��U�.N���f�L4���:��mŷD�\����g�����*#l�j�m�NiW�y�4FQ��ǹa�D����9il�"u�ܼ�4l���>��b'B6��C��h��"O�.Q	��y� ݇<cO޶i�99r�gyo��1���r�F�;�/dAG��(�z�ؽed'�(1�n��#'��w�I�ُ[�w�'��@@ѱ.%�r��cC���/�z�{=QkSr*=�dSp�؉��@VY�b՛�4��^Լ����s�fq��S� l%�8�ѡ���ו=+s�ٽ�����pG�y~�d�5R�'.٥f�f7A
�2�I�`��YL�����D���9#�՛���2�����cс����JIN�%9/���Μ���m�h���JqGD��2���� B)"6��H�{h�嘖�q%��C���v%�N��Oj�t<�t�����	H��Jt�fv��t�6��)Ċ;�ܔ-BN6�^�gI�8�p��Ν=�s��%	҅b���5���t%mhD$�t�)܎s��V�I��H!$�IKl�+m"G(���I#�Έ �	K�s�P��ٹm�;�]���9�A<�P��8��X�݉%.P���&�lm�1�~$�ϯy'��~����1���>��W��7+��5g<��Ǧ��C}{S�3� Sgk�H�~�pt��: ���� ,����G$B-pǇfss���G)�P��}q8�͸�<�9�q�` |z��x��]���'4�w	�:��)�v�t�7n��s�y=+��޺K
(��\���3Y�"u��E�G�{�\�� ټ���l��{�k��iӫ��{	����@}ɼ����k� m[m�����{�_P�*�i��ܞ���@ 77��� ~riQ�'�2�v���;�����|�N����K5ߍNk�0l'�{��$�K@|ʔz���#�����lK�yɍ����&�έ馹+�Kaf ������_-����,o>ޜȏDG�G)�I�Bo����Ubn����6�hX&���h���Cj��UM	#;�G+3�
���;��e+ƶ�\�6v���� ��~Ӿ����=��ߋDU�1�jiPB ����2.q����/�-��s[���@���Tg���6u�҅�5�Ӂ�$dmZ�n"�I%HC���8��y��n��X��)os�rN�8F"U?|rg�4�{�k�6 >��cς��|�膑���ɍ���=ɥC�1ʒ��!'�|�'	ܺ���/��������@|���א� ��z�>���z-����������m�rGfb2zviA���z� 6^��>{ڞo����6ގw޹�n�����K3>59�N��$�qk���d� �o��<@����]~%��K�{z>���@�V��\�))B#3���\����rf7z���]��w�'o ���L0��k�d�g��}�w$�B*��<⟤��3Co�Z
6�3���N����v\����{�A\|�?87���-:�R>r�4@W�x/�|�I}�}�32i�ڑF2ߝ��N.<��)��v�k�2�<��נ���y'�:j����4n6뱼��,{@����v6V�<L�*��L�R��Ρq�לc�y���ײ��'nh�v%ݛ&�Ux���u'�::�ܥp�W@���;6t�l�TÐ��*�Xڍ��3Ŭ���c��oK����˄�]���p�3,�p�:��9��sq��.x4+�y��s�d���N��1��++p*`J�:Ͻ��/�[T�����SP7��n` lܹ�g3}�l�����596&	0!%՘ ֽ��č�
J���ɘs� ��m�׵�,� ��=�m��-�מ`	��}�s��)���A��H�c*�F"ף����|� 毞%���P�	��Zd�O�W=?~$�:���	���@z� ��-��H��FON�j�v���n��bH�9��H��{g���W�x�|˗^{K~��ʉK3sZ�ŀ��P��SR���w8�Szޱ��ط��<o���҇Tֳľ���͟eR+�:ە���#ك��h�]"��e�@PE���P��k��i��-
E;����x�ٗ�0 ����'�=�zb�����A�I�G� ���ttjجpeǉ�2A��m]�����"�Ҧ#����*�\��]�	����,��ƄRE\�������f}���~�`2'�\���6n����<$�"����n�����wǽ�gǧ�ɥ<��s�:o�������IЉ��J�������`�{=94�!�b�8WM�D�Xyl����NM(y���Ydb���u�${�=)�?)�q ��KCm�'.�ޔD���sN�)�,�]2J�7�DB��,��c��;3�ӳP A�{�29SO9�u���)����DB�*lA��s���Çw|iL�wDv啧���N72�0��c=�Еٍ�$��N�:]���]>p����Q4[Y)g|�^k�O7ӓ�z@�y�k|ړo�R��k����ɯ��-֜�GIB�Mg�������,Z�ë}��{��v��>���h�;��� m��b��gs����ͮ��mV8���;52_ �z���&w�����л�q8�Ԝ���r��Ac�p��p�wڮ�$�F_B,1_<q� �f���Ͻ�s���/��Ғ��_Oxk�e�����[����OӓPg����0_|Y�D�	(ˏ>;��oKs�ӏS� �agf� �|ﮛm��x_N�?��j�I>پ��>1
�de0����,�� ަx�;���y�`�wI��|go �z;�N�����������獭���V)���֋����6��-n|�-��햺���%r��lA��/Ie#��;3�NOM} ����}����g�`C�2.d�$[�m����ϐ>s��Ġ-�o�m�H�l�,��ϰ�{;����ץ�"��=� Y�_a� ��0 Okw�;��\����j�@�G	B�L���ŐMg&, s&�]yn��KrÀ|�r{1A��Y�>�����جqǈ���sZ�����T�jwA 泓1a������L����f$o��x�m1y����DY�٧�V���v�ٙ��6%��&\�ZQmdCc%��o&eF�Jn�����S�x{����m�F���3���,�"qKq�ǧ7vB&�����cQ������%��������ɯ�}��֘�ߎ��b��;@;��v�2Y����n��4�h=$.]m�
���W|�]e����������gf` ���48;�W���{��rw�jU�$��Sk�"R���55c�1����]]��o���,��r $f��1 ;=95��w9�yw{�39�5Ԡ|����U�eT [^gŗ��� 㓓P �^S�����|&g&b �ONA��Ϋ��"$-͐������C���'���2 �=�4 {���/��߬�wZ������3>>�mq
��V���~s'b Dc��쥽=N��LK�tyB�D\�=3 $r�ң>��f*s�8�~�ﷳrs�/gH�qD4w����{%O��Wr0?i#�q�9��{f���f��يW9�ز7�E��:�l�o��)�U�sZ��x�|��jC콇��q)�y�W��З�����<�����]�����>jݹs��Kb��l�6��ˬ	d�7A۞��\����䮰>�Ll@#�N�Ի��=�`j�'l;(�b�m�4�n��ۨ��<n��j7M�a|��<ڪ�t����=���;�ϭ��R������;v�Mgd���n�]��H�C��=N�v�vγz�n.ca���v�(�Gi�۞Ş#9�&�cnK�x;d��P�����~����I,e��F��f}�g���&� ��ݝ�F���}����yu�1o��MP^����B�a�������\ww���ğ���I� �wٟQ���M�=uzo|����؀�v��,�(���!��*6 �wS�׸?�twG9�6��ң��}������[�+B�����׍s^޲d�� ri*��jg�|�ys���-f�G��M%C�Wj
7%��L���Sܙ�0�o||�'-�}d� wg}�@p�b�	5�m���:x44 A;����x�ѝ�7ξm��6<u������r�W hs����u��P^��!���y�{	$���Or}�����2_k�A$H�w2���'���U���6i�P���z�i�ٸ{�2|�$���%�J��/�=S���?��՘������:c+) ��p��(���Z���5��H���\��
����ӽ���-���b@$������8�̎h�7;;��<���F�ho^5�e�g�X6����g������9�7���g�m����%�x�Yt�f=��^׻ܚ4r7�l��Q �]��Y� #��rs��������?��q�ys�G7EiI	0�O��m����}��]�ǰ>�5��k�:k ��M�({~��O]�T���U��!+v�2��6�݇8[y��䒸۬sIyNq[=O�(�����RW,S��n����o�8�0��I�o�_�g�op���쏩��Ĩπ�[��1�<:�m�iL�פ �۲@�}Ӵ��DH �L� ��NMA�&k���vpn��c��s�k��i�7�Gu1?5�̄�$
~���O�|��þ??��	g�+=���={K:�w�٢L�	�r�M�w��@��՜���sȶG��Qj�/������I'�=�� r����ɥ��WYe#e0����S�n>p�߯��͚x����������T�1�b#�%N5� l͖E Y������ =�N��s�;�g�}^���T�y�0 {��Pb �{=�gc2����O5Z	cp�=��=gpke�w�:B셵�y�+6��,r�r�_z����*�am{s����6���6 ���3�k�_��|(}!Ɨq�	$�ޜ����E��M7��,�P�	I){�3�/u��lf�'	$���.S@�;��f(1��;�u٧u|q��ݼꂥ*,va�ܙu���vd�Dz!!EF�7z勒K�jU_�z �{=�_|����,���;5���P�	MB뙢I8���@�&�� ���g�:��t�<�H����y�n���U�|��OW�v�;��^�7�$�>����2�9�#��"�X-L���E׆����_�2v�\���)RY�|�'�b���N{�5c��מg�=�z���=����M`w�3���.��,]���7V䎎�Gv	gE�8��F�2�{iz�G�����,�(��yvr���y�����L��b֌�l�1�zn�@|s��́�-�q�~�X�8Nzq` ݩ��g%�^������m�|���6-�g�7��<�,��k��N���Uځ���-W1��hm��\����_g4KV/s�����|{ܝ�P`��Lo����t�v�Ufɖ�NGw����I���o^�Ő�泳1  wӖ_��x��������iH8R�$����ng�  {�����S���3�FM���	7\��I�c�Ҫ���.+�p�ವ��	[�ʁ�k�{�ɞX]ж[���SUJO���ޏ��o���'���~�dHŸ�dA8�=pNn��;E�l���w�Τ�+֟�3ȼE.Eh�vL;���d�t�n��\v ��}��ƍ=�ky�9�Y��~�aX����>6�/
�|���Kډ�r)Uܘd�;5	�u���ӵ��ٕz#�P�E��Ó��-�ӳ�!fvzt'�5�ʕ)��zI���)����S㋬괗�T6f������e�p��W��I�h�b�K:!���&O�"�E��eͅ7��m:Vv���M�'[Q)�ٗ��3�2epm!	Y.m@�����7
.E�&H����zHf	�4��
�uhw�Z�ݛ1o���f�b0��f�{��w�x`m�x��My<�������,�j���{P�'gd��WcH�F{4-'m���e]�������ٸ�T�Ny)���y�ln{�կ�q��0h� �	�Po��@�����F$���5�{���{
;D�OU��ת���d���tBk��m�Z�ޜ5���v��#���+�y{�ˉju���Is�S�@�h����%�V���F���;x=B����5�s9�eՉy��]0�yGv���q�a���u��oƔ�.GeM7Ж�rr�<�l�"���Y�M_�4={���ͳ���i��Wv'2i3�
${�eE{C���;m<�b��4k'1�EЍ�(aY�NT�}�Koh�GNO�=��<��w��������I$��$TI9�!��/�{ܔ��q9. I�.N��I�ݸ:��9�gRw���PB[��[d�����"B�c��RH�$"�(���nB�t\�I�e�'$�$C�$��4��qy�S�s��eO5�r6��QN*r� NA8���4�8!LjĠ��AD��=�GǸ$��(���:��8�#������:y�9��fHq%���吣��r�"8A#�2	!fyw�Y�֩f�s�H9%8s���3�f鷽�Aǝi%.Roz�D���{cM�&�V���9-�H�2:��H�fݧ�H%�9�R6��kBwl}~|�q�d�����Cd��w^�����B�t����wF��b{.��n�Q���'hYwf�ě�DO��6�`�67��lu����C��S�_�e\8�;���Z�^����l��|��tl/����h�S�Z�^u�qEA�sѳ8�"F63�ůf���s�'��u����8��ёv�g������sֳ���	�h#��r��n�����W8�[)���.͏c-��	�t<�Wn� �B���5�k����4�u��.�^y:�ͣ���}�[
Ɖ��w��:�띘�u=��c�6�b�q�NKҼ���h�oXw���Y{6���W��7N�D�{�jǭݙ�`p�n}�]l�74� ^L����g(�
��D�צ��v,v:�n�&�yxxy��uy.�6��ٽ�췣����ͯ�>_>���g�8�սlY�����[��5���<�'�#�vs�rc�z����ft�gOh�n|�J�����wn�݀��=��pb�P\���6�l	;k�i��g)$\f�23���=�v;[���m�K0��.�y{����R�á�9�ŷ>V,�F{5hNn�Xv��P� ��p�o3q�e�n�dQ�;���kc��A����Ʀ��c���>Iع킵�#�b��ҝ�Z����Kv��BCJi��j�kڽh'�:� ��S�e�su�����m�6�ݸs��v�x��B����-n�K��b܋��P�ٺS�*%Ë�n�M�f2Y}��� h.��-㍭��˹NGk�u���k���:�r�9&�]�n�94�qV[n]à��]��ϳ��0磶CN컆w�Gj띂ŝ�c���uF]����g���q!⍞9���a�fxEm�<��Q�HtE��3%�Ю���s�Z��� �d�t�Ć���I��;t���K�m[�1sڃ���]	��9�����n�K���ϫ�M�@�7Okp��p���wNT��5u���ݛ��,<���lN��}��o|����d��gm�]V�\�諝B�s��y;up�rǓ��NE��c��)bv�qq�]{l�d��C����_��[y�gG�q������gq�����Uv1<';m��Eh��7j2����qrNX�h=w1ȸ7��J[���h�n{<�dȇ<<>�
=�\n+l�>Ic�&�뇶�c��t��@�[<$�u�n̭�3��N�9��C��l�s[v��w;mmv������<E�n�jb�10���?��YH�\��7���7�Y٘  �^SI4�����}����95�����\2[lQ��޽;y�=t�s^�w��{�@ =5��� �r��A�X�~gqD�؟{g�+�Nsˏ�����Wdy����>�@|�yc�����}�ۗ��f>� rk=3�t�.����v�r�hV���=}3}z�w���{Z׶��<s������,��|�v{ ���-�٪��Y;̙� �����v��L��3��c�� ��=�5_�vfmٝ�� ;˯�ρ～�}����;~���HEmi�I!u��k/  $:*��oaz��Ihݨ�s�3�DRһIx����ni���w�TlA�v{F ���-Ա�ư�^���>AÜ����U�YE\�F��'�&�Ŀ��}F|��p��Q��β�zvn܂��+9}9(iՉY�;sx/Y�Ko����]�{�V{X^�����f��k��s3��_x����X ����S~�����?fL_,w�l!F�m��rU��$��:8S3��ݺ���߽;�>���n{���g74�P��MQ����k!�,W�W��p��������N̙��o���MP@�����٭�ilmo�y��5�_Pλ��B�X�b	�L̀Mo�0絵�M����;�4�@#;���1 ٛ�� ���Ս�i�~}"'LTW�編ݡ��ϧ����jY�����Q8+���Ns��:���;UL<n�T9����6f�5��T���;�H{&������}����-eu�|vw\��|�Ӟ{=�ˊ��-�T����0 �_�BI=�x��I�RtBn�ʻ�D�ǌ���(��bks�1 3~���p�y��L��3��~7��Ű�=�Q�t�MKlV�ͣ,��9�ur϶�/\���I���~�nT+~��r{�
iq��x�ݙ`Dϧ�&@nf�L��W�)mtp���!���
����{��	$��M8H;e�� �{�^�{�^;׾e}�f�9��bŮ¶��»#�,����x;��b#�wK�c���O{���I';e����Cܑڭ�<�����2����þR��On6riŔ���i��u��9�2L�v���C6�����Q^�f漲6 ����>��&�g�n.�뜨�5=���ٛ��|}Ǿ�'kN�S=ɪ��;�a{[�����g�@ 93}�� �ܑ����K�l��,����b�����&`{�^"I8O��8�M��ϝ�w�$�n�阀��&�}2�GUqX���F�aw=v�U�rr�l6�d��P������ة�Q�2�Q��׹�LZf�F(��
}�}v��!5��U�9sfaͦ�T�̝��nx���F]��Mɢ�Tм�3�<ȳ�����|�u�3�%���G����;il֎p��;���?���?���)���=�����F�}�_���*��Da�*f��l��S\MF��Q�u��}�	 f=Ρw/d#I�L�#D/]߷�у�#Da�����b�
b����j?s��F5��_F�����Ә:F��mDV���3�0\6��t���F�T�
+C��?������-9Zz��1u�/W�^�ǌQ��a	B����B�P���G�w�h�
f&�g;5�]�Z�j:ߥ|�=�f^�cX�a�F���9�4�l��{��#�j��j�F�4`��~˰ǌ#R�1}�徾>s���{]�Ǎcq���!�k�٦-3c#j8��>�F0�B�*(�Aϻ>��W��+�w~�u[{I��J>�9��Zӱ��m�����{�L����A��5�#���f5�#��0��#F�W�������݌1��SF8�1BQ�N��1l��NF(y�]�l�F(��~��KYh��m|4���n����}}���ԗ�L�
b�(Q����1i�n�F*aN}�w{F0�c�2#���=q�4�o�kO��l��WXq�j0� ��js�i��-�h��}�4�OF�5	��a0q�y���bx�1IA��4}�g�<�(����5oY���y��c����3�>��b�6���1F���6�%
0��Q��#��z�b��]�~�/{��/����]�î�y����ήu+�>��`Z��r3��f����.i��wL^CG�uNl��
���2���9������/0����y��D	�">�3�$l0�{$�m��$�T��*�h���m�ٰ���=E�.�RY�<�:��\7	ţn��Z{HeǶ��}cpg�ή=�$�ay�[����x��hm��v���yynSQ�`�;��5�;ݰ�XO��ts���Kv���`�q�M%mӽYݙ��8賵p��sј��t3H�n��͎i-Xzn� ��9�zw�9�.u�W;Gi��nĎ����ܣ����2\��;QU߾:���SM���F������6��F��a�Q�~�vcX�0��#0��}���h�F�}�����*��g:ÌT˓�Y�-0�*|j1G���h�c4��|s#��Zr��&�b�bdh�絍`�5�Q����^>�\oW\2��,�
���Fƈ�8w��Fc�20�#Q�o=�a�`�a�Q�a���w���W.^�����L>l#D^�+��S��U�n�cF!�����m�b�A����s[x��(��b����1�g��|����{��Ch<:h):}�u�A�H����e��c��Hgr��b-mءhg�F�5�N]	#��h���G
��$��� �S
z�vtkF��a��h����0�*aM��	G�=�4����%9��*v�b�5��]���Q�7/V��Zu�QZٌT�L����k�(�q�0��F}'�f�B�	]S��mb�8��$Ȭ��xc
f#�0�#G��kl6�L)�j0� ��j{�i�L)���U�}��?F�#N$UQ$lB��Uq���Y�>�՗������+@d�I�-��UҎ��R��a<���z�aLXJ�%h�w[a�*x�b�)��k^��1i��Y�x9��Ϙ��9�˴m�	B�*P�����m���p���p�Z�E48��F�Lܞ�g��F�Q�j�v��M3��dfg���붫�B��$�=faW]D�[Zck�q�]9�QV�Hȩ��Mҷ��f���	8$B�(�\M��-1O,~x~{H��v~kFdaA��h�����4c�#Dq�b��ڟ�f��A��j1G�����KT�w�h��db��ه2=��zz�e1c1��]��mc�(�q�0���;�5��l$�F�h�#���i��se��#�)�aFF�j2}��v���5�F���=�4�l���z�r��U:C
lfA���!�F�����������4W��]�k�����;'9f��Ͳ1F��Q�8��}v�a7�����v}|�
��G�/��i��|4�����kN��ь4�a�Lݚf��5�#Q��>��]�5�#�W��?�U�Y�pl:ì�#Ek|˶h�8�1S
b�(槹f����1S�Q�85���4�I���_uϬ�IN���{���T� 2ڏ��5�j���"rz�k=�I�B�}g�5���=[����ˍ|5�&F��7˶�x���(������
�HP��Da��Ѷ�F�|���Y^�:a�A�=�]�Ʊ��5�#��N��0�-�h���^��M:5	��a��>��w�#�`	#�
+�%{�Np�F/���b�5�##d;�w�4Ŧm�Q�8��?s��F0�B�*��8����J�fwx]����>Ҏ.],<ܥejT��-���kz��f�[��#QF���وkF��b��}�U��]6s~h�)�������x$��&_L;T ����1��bI�n�@��tn-������I�3;���<�E����4=j��_{��u��#Da��~���4ŵt���Q������F3#d�g�2=��5Z�e1c1��j�붟��w��~�/�S0�P�>��f�P���(�8�#�}�oh��F��a*���a��߻{��]��yq�5��L��4�c-�h��v|Nֵ
���V�l1�G��]�'�#0�)(#E_��o�(��;�����U����l���;�w�4Ŧldb�)���<�;v�a��F(Q���5���x4F���~�'zM�5��g�X�Uj�,�ڜR��8�r���64d���ltץ� �v���|���;eg�<�3���i�al#Q5F��a{��1�aA��aF�sW�ޘc0���w����J�S���u�����i�wA���b�5~�nь���2ߗ�lth֜�l�*f24{��\k�(��2�Q�-3�s�k��l$(Q�q�0��{�h�
b��aF�^��m��#Pj0�=���{S��S9��٦e���|xjh�4�!5/l#F8�<���0�RPF(J���=q�k��F(��Q��o'�j߹��1i�db�D�j?��nь0%
0�*aP�}w���&��9�^�q��Q�"jL
�
 i@�6��D,}-��p-����a���<�r�Ʊ�aF�F�^���h���0�QJ;��Y�,�=z���ݪ~��
��Q�hnW(��S��P��ȳ"��|��2|��5�17�H�us��s�fr�r�̵���ΝU�m�eP�4��\�_��<�O��b�)�9��6�F(�Y�vM�h��T��m���w|�q��Q�1FP�?I�Y���$q����:��K��@�G�Hg3��aLT��4sZ��a��5F��a���ܳLZaM�o9\٥�_��ڽ���X�FXT�r�Ie�Z� ����kZ4��l�i8�uѧ]n������Բ�E�����G�G�o�h�
b�PF)(#Go_r���1GQ�221FC���l�����5��q�����Nm�mX�����1�JaQP����ݸ�o#J8�z�yQ;Z�N���m�Z�iF{S7f���5����VsW;�����L-߯.Ϛ��L�#�F�����a�8�4GF(���,��S=��|�y�״��ŷw|�GY�F(ɛ���i�P��b�`24{��\a�*k�����ڡ[�L)��0�Y����������o��
b��#���ݸ�ƣ�j0� ��j{�i��[���0��94�HMM�ю0��{�tr�֪W�Z�����1d���\�ǍcaLT���	�w�-�L�#j1F���{�h����:���L*(�B�_>��4F×X�2ϩZ,b��-���jn~������F�Q�j&���=vcX�0���t��ǫd 2$�'�|��� cF'F���%Ӝ�طt��S85���ь�db�}~�l�J"w�p��dʆ�ۊ�f��v���oma���a����bad�R��B�����`�T;��V[�]1�H7͸s�~#�q�n��nv�^�ۇ�8;.�r\�i�Σ� c\sΪ�v���� ѹ/]�l��5Ɯ�ݝnC�JEw�9��}�'+�ꎱ�rmÞ���r�l�	�;�\䵸j���׳�S��n96S�;��wV=u�g��v�2��i�퉄������v灩R7/���ɞyI�kp��Vq$��0;G=[�h���y�h��bJ�ZƳ���/C^U����A�2�H���|M�j==T�6/������ۍc�(�b�"�(���,�Э�b��h�#�w��ь)�0�#/�����;�C|֙����b��F�;;�-��[�;�g�5Z�uF��Zݰƌq�y�e�`<a�%b��o�9��>:׽�{�5�_�?�X�S2�Q���9�ش͌�Q��b�G��ь0�(��{��^��&���w'���q�>��Y�y�D�j�;+3嶕k���YlZaM|5F*aO�s�h�
a�� I�
���x��|������#Dq�b�(�Nr�b�]b��aO�w�h�
b�o^�,r=jD�V0�A�I��x�O���QO�.5��aLT���Y{(V�1S
q�0�>�nѶ�L)��0�F}���c[Z=W��wY�/�m��F�����l62�F��=���&��joi�G��a�F*aLP�����\xc|&�\�I�zN+b�:��$߷�ح��Pq�5~�{v�aLT°�F���޸�o�Q���7�}�~ZPX�����G\y���.�8�-�ENό�oRv�J���(��������Z�:z��4Ì��Y�Yl���A��5���vcX�0��#0��_���cF'F�s*�_I��s��a�*eV���b�7A�ƣq5w��F0�*fo�E8�Z��0��ֹ�6�L)��O{����M�U}�k���������Il(K�t��g�oƽF���[�&��Y�[�nr����h\:v�{�6u{�,�"8��;�_Y��p=�	�фq�0�>�nѶ�F��a�>���1�j0�F�Æ��|~Rj~�8����Y�H�C�*h�i��Zݰ�*aO~��Ѷ��PF(�h���\x5�Q�1S ���<W׺��T����l���S5|��v�aLT²�HR/���c4��S~N�H���Q��4�]I���ݖ����������Q�j5G��.�kF*aL ��4_5�n0�0��q�b�Q+���b����g��|b����S����6������br;a)Y�m}ZC�~��5XҦ��a%
2��r�b�/����>���m�{���l-��G��{F0�`�0���0�Fsw�n0Ʊ��5�����r�a��a+��y���r倢]UB���FJ��臎�����="���vZ�I��ſ��KG"�{l4�����r�0x�1BPF)(#G��ݸ�b�)��F(�'�͖�l����9^5�=�ѭ�}�m��mǗ�]�a(Q�Ja%#���]0ƾC߮��e�;A��y�-���jV{�[6�l#Q��5�4m��_�7��TÏ���ρ�aA��aF�o����`��L)�)D�{�[�A��1S��ns[�}������|��Q���}�h��kUScb�`�ѻ��t�<b�G�
b�U{����[a!B�#��m#~�t���~�=U���z)��+��p.�� ���Y���[���o�o�x\�۬�<8&�wq3eb��m��j�#2q"��3��[t�`L�N�BӐ���f�0v9�ؽ:۱��[NP��+�k6�۰M�c��u�M�f���Ι���꺴�e��S��{;�K�������#aP�j�W'e���=��VZlfEMT͐�ʝ����;�-�S2���yiSM#y����r��~���m�@�"2Zc����ɠ^y^���2d]9�o�j�ĥ�M
xT^DX���O�T<sp;�m�x���ю7mT^�DQf0HL]6"�.\�����g	N8��=ݯ�Xj��l�9n6/ZP��0������m`�8�v�����Q�
f�՗MN�C ^���1��\��h������Op��A`�ûN�3��^#^�r
�ٶ��L�Ɲ��n<3�z>�7̝	�sˬ�y�s������k��k~����h����
t4+����^:�޳;nDmY�	�5����k�pt�.P�fﯧ�_l 4�nCI��!�Y�iR���A%{S���:Fj�h�Ɇ�uB�tdU��4RY���ܽɊe�N��.r�MdJ�Ȯ�R^��c�@�J�=t�������7����<5�����uxL�&��b��x�@2�/]�k��&g�^�z,��!�Т�h�02%ml*�&5в�.a۪��kh�@z�7M\L�̭f�@a��㚛��춽��؈U�f_8;᧫���o.�%��6$�Dp��r:|��јG\8q�i�DD�$R�q 6�AN��:ԤkK�`��j�i��9��$�Jmؑ�Hm��p���E8��$�Nm۳N���)��I�h�v3J!���Hqn��J\I9��J:�`�H$�m[�XD۵�u��K4	�S��5�m��cY�����m���E������\Ysiki'm���rC�e��'@��&�q��vq7X�%̌���3��p�̋9m�쥫tֲ�.1�r�tڰ�gZ��-$���k��Y�U�d�:e����\��J/l�7f��秂�8;�i����H٬[n[d�Nm�!p۲��n�'%���tIg3q$Q61��޵�aL��20�#Q�����k�#Pj0�Tʯ{�[�l#DGyt��OSN��[�ю0�;�s�T޵�����{���|���RPF�����Ʊ�85�##ev{�[��F(�������1��y[��Y>�+(Q�������x�#�����v�����J����Ҷ|0���SQ��>�0kF�_�s�~�58��4�tda!��~�0ƌN0�8�1BQ99�-�e�F*q��j?��]���Q���_�ϥ����tX�	�mpe�����y,9;��	8���9�{֊6���E>�>�m�u�SU�^8Ŧ��n��a�*k�1F�(��w�^�V�Jah�#�s��ь)�#��}߽��=�ӡL<����t���5�F�dd��,�[�=�kM�kC�ԛ�h�q�}�޻0�RPF/xַ��\�Ϻ4}�^��(�Q�221FE=�se�i�db�G�
s޻F�a(Q�EB�'��'�k���/���X���F�s��c<�����ʴ��FL��Ŧ�ƣ�MF�}۳��aF�F��oy��I=�aƏ�F*aLRQ==�-�wA����S����6��'ٍ�	��
֞��i����{��t�W�[Ç;eo��q��q�0��]�嗺���F��G߻�m�3�a��5�}�]0ƪ����w,����9۩�k�S�{{T���B�*�N�bd#��,x�(�vMd�&@�v@t=����I~M�<���󬙷���f?/0���aA���7e��֚Q��y���]��'.i���C߽�������RPF���˦c�[g��φ�G?aDQG����X,��m21F�q�5y��v�a��S0�H�o�L1�4F�������t����`A�ۉ�r��Zu6h�+�r�c/�z��t�F�W�#��s��o�n�`�����|�L��2}>ݖ̓a�F��a>�n�kFda��4}�}�6ю0��,�Mn��a�*ez{,�-��#0�*q������dk��޿~��El%�x��դ?��s�q�j8�o���ٮ�rI۾�W>ݖŦ�L)��G��nѶ�F�0�#Q�n����F��Sn=��ŷ���==�-�[�Qr,��-n[[#�f�U�������F*aLQJ���޽<Mcq��S2M]W��]�vk>��}-�L����1F�q��z��%
0�B�#G����ة�<��q�EZ�SԪ��@�4$����Y|��K��\�F��a��?�~�15�#�F�da;>�^�m��SF8�1@�OOr�b�����ܫ��}�S
b��j<�~�F3��2�7�&�qG4kU�LX�dh޹��5��aLT�Jezw�^�����(ԟL�=a�*aN���{F0�`0�#0���k���5�F�5Fdd���Y<E�$�Z��i:���|��7i׫OV�m�9�F��������C!�Q�4´%n1p9��;�(K}�����;5̽o���Sz[� �Qnܖ�����9�]�����Ѻ���ܛ�28�j��f��Z�k�wZ���5�up��u)�zznRq��67T��{�v�]q���nDSc����]��L�N�v������kF�W��ns�zjwgonM�;0ڵ�9o��-֒RA�Yu��{"A��an݈'p׋��=-;�V�u��L�.�<[��m�N&��ܡ;'`e�x�;�bOU����}e�&5
�N3�ÇV���Z���k�íaw�v���*aLXJ���r��5�Q�1S##ev{�[����5�~�vw�w�_vŦ������1�)B�**a%#��;za�#����MkZ�=h�Zь-��^�v[>al#Q��5�|��>�}�[a�=]�Mc��#20�{_}��4`��a�(���Ŧ�L)��0�wM����wh�y5�57��tl���`�m��[j4ww�\k�Q��aLT��{�^�
�IB�#0�5�}�9r�OJ�����taFA�a>�_z���F�5F���ܲ�m��4D�6�m�[[��3m*�[q���������>���{�l6Ł(#��ٮ}q�ة��b�)���͖Ŧ�Mlq�5���ь7:ﾯ=�u�o�q�z�F�޳.0���Gux�R*֝�h��L1�0��;�-�L-�b���#����6wr���aLT;�}�m���#0�(J'�ܲض��1S�F(�Q���1�1S=ϳ9u/ݧ�����;F���*�6ö@�mm�g���q�3����f��s�V�	��}��M�dz���l]aM���Ƽ<b�G�
b�Wgye�[�L)��S��}��S1�a����Nn�'u�zt<íy����cX�a��aFFN�r�a�[�k�����+Q�Z�n�cF0�;�F�S)A���1}K��U�75V��`�M��3��i�N�֍º#K;$�S�z����u��wѿo�/85-�~�wI�'����B^�Q<��Յe��ٌ~%�2��k��Q�221FB}��e�i�db�G�Q��{�h�JaP�F��{�r��F����b���a�Z֥Z�kC�m�ة��e�����F��L)����6`��1S
h�Z�>�����޻�F4y��8�1ID��,�-���T�Q�8�|�v�f21Fk=�V�MԭT���ٶ-3;��.5\�o�ݣ����(����[���Ŧ�ah�#���w�c
f#�#�g�_޸���z���]��W���mlj0� �����l#D���aSF�֣�z��0�F8�?o�]�F(Jǧ� I�J��'O��I�6>����궩���F(��YlZf�F(����}۴c
b��(�B�����0ǉ�0�{���~t���e�dt�T�����
�bӥ�����޶w��=��3�y�c�����R*֝�h�#L1�L#&Nz�f�[�L)��S���ى�aFF�da'�_��a��Ѿϧ+��eu���jf��ˠ�T��b�)����6�L�Q�f7͓E9R�i٦-�3����'�Q�8Ǥ����T���$&Ǡ�3J�lYe
0��p=�;��S1�a�j3��\a�T���0u0SآAz�>�ϬQ�����)��IU���h�G��]�l)��SJ�߾�]<k�
b�FF) ��3��`��9S���jܟ�����'J�}��|<��O��mY�t�_k�'�;/�L�1����P�Ǹ����Fwv�����?M+}o�!�����Q�1SPq��z��	B�)��T>\�3�����ik����k������	#ꕖ(��;rs��U�ES�q�5Ѩ�5�#���h�
a�#�20�}����1���SR��{�i�7*��f�\�9�F*}�q���e�1�21FMg;+oT�J�J����b�
h����a�*aLTÄ�F}'�f�B���W�=[ѱcb�����6��0��#�w���Q�j5F23���a�[������wr�}<��CeGT��ܠ�=8N����g�9���Ի�]A�3gu`E��9���Qm$�;���U��8ҏ����X<a���J���_n�caLT�21FE�k�٦-0�*j{��㧺{Y���b�bq�3.ь)��VP�J?��s^��ƾC��w��R4Z�[���0�c�׵�4͌4�5Q�j�ǟr�p���u���r��kFdaFF��}��cF8�1S
b�����f��
b���s~�a�}K��%w��`$zH��{�1H��N�1m��3��]5��Q8�E(Q���,����S�Da�7�
���u�ݚ�w���0�##�5��.�cX�a�Q�a���J���J?���ߢ-a YsM�L)���]���߷�{���|�0��A�(#G����Ʊ�0�*dL�Q���,�f��Q�(9�]�a=�_of��4���Cǵw�!m�ʖ�9z��|1��Q+��������\���k���A��2\��wǆ2�k�bz��w0m��{�=$���L1�Da/�����G֣����a�*g�j��>L4�5�#Q��>�уX�w=�W5&]l�1�̌#D�>�n�cF'F���	G5�r�1l�b��p�����f3�7�~'�M_��v�R׊*�{v�&;M��7'��6�SO����<r\��5����@d(�-o��_V�5˙�x�S0��F};�Y��-0��F��0��h��L#�^~��Vm�N��|a����0�X�a�F����Y�L��=7ǈ��9J9fm�_�iƔ~�~�,icK	A��4�f>�߽z�Cm�/�O�k�����9;�Y�(͌�Q�1S
|罤m�e
0�B� +���U�M{��Mn�m>����FV�T�Z�[F��0�o��F!��9������`P�h7>�S���z����y��q�h�0�T�N�i�f�#0�*pj>s��1��(ɿ��0��
f�=�b�ѻ�����߾ܞ���{{t��+j��a�F\�n�m-0��F*aN�;h��L#�L)�3��~�a�?���֋���U;���íi��0�#3\׬���iG�旻Zk˚im���aw٠�x���1S
h�k�\x�1G��E��g��s�1c
b�vk\�LQ���Q�(�q��{H�b��(�JG�z�b����Q���;��Eh��|R�,|��nv�����UI�^�W����G��tC���k]\�ꏳ׾�<�>vA{L8}�j_w����"��؆�t�m�#;7d66��ƍ�n�k��ExۓϘ^�4�a r�i�����ۈ5�l�#�s��{Z����zi�oFh�F�:��q��Dh�Rں��8ru��'��ͽ�"n��u��6��˷�,�]�\vR���M�֏<g�,��Ǻ�8��B����ٜ���on@���gm�qŹ��Y��m��n�C��шy��S۶:k^�����Y1���Qv�>���+r7b p���y�j�'j�'�a�~a�}�٦li�jF��a��n�kFdaA��h�����cF8�4I[梚�j�kW�r�[�ԿY�-�b��L)��k_,ki��ѩ���@d(䶣1[0dh�o|���Q�(�_?�_;c�:�u��-2I�ٮ*��(Q�q�0�s����aL��dF����0�X�a��0�g=�>o�]�U��g�*��ZiG����,�A]Խ��F8�;�v�b���RPF���޸�b�5�
b�{&�����J�3��d�g1i���5b�D�Ͻ�c%
0��Q��H����[{I��J8�f�xT��-�ϕh�`�35=�4�ٯ{�o��aֺ��#Q��>g�vcX�0�#�L)�}�����L)�a���ܳL{2��lMt�h�-�g>H� �A֣��˴c
b�a��>�1�B��Of������5��(��R��;�5��l'����뜭��|h�#����6��3F�3��\a�cQ�j5F����,����/]v~��d�~���\�t�aB���U[��x^[V��ֺ�cm�����#��k[<o�������X�����_!�5�i/�m(�%b��4v}�/L6�O�Q�db���b�
b����:�Cx���}߮ь)��V"�F�Ͼ����pߍs��h���u�=�m��3ڟn�3ca��5��>����C��;��W�pc��=�U;$��{����ҟ�0h������
x�L�n�_S~�P|�x�j��_�}*W��)��˳ɬa��0��#D��oL1�a#�#�{SܳL[��N&�u��$ޯLͿ����R����\־\k�F��Moߡ�B��j��b�0dh^�ǌQ�8�IB��Or�l(V�1S
ph�#�^�s����^w����o�G�S:#�#�g�Ͻza�`�a��0�Q�Y��U��i��z,��,����$�i��ϝ�鼘X(���E���������SE��/O�(�Q�2�Q����LZaLT���(������H�<������� B�� LG�/{U����(��<�dh�al*�l6�Lܝ�b�
k���5Q�w��1�ak��=�}�|Fa�F�k���4`��F(J9��Y�-�A��5��G�=�c3��vK��m6K����b�XB4�9��{WP�[�]��x�fV8F����ɖ�_&���7�h�ʃf�?b��L�������aLT���;�5�B���S=2��fxi� �Y�+8�)��#X����^�cXF��aFF�g��Z������iw���X�B\�ю0�}߮��#R�1v�}޾���R���rul rOrM l7�߮`072W��k/�� �Q�8[��+,OZďCz���y��X6���q�ձ6�����Q��e���D�=4,�thؙ91qUy��ײ�TK�A#B��Hb7�J�;�Tv�kc��t��K҇���a.���g�I@|r���w�3�ߣ��$��SB����e��ܕ�����DD(�s�@������ >��rgK�pzS��tzԏ\4�b,��R�Y���V&p�gݳ!�yKqH5'�!'��_��$�$N���	&���BU�Z����}m=�	���ۥ,K��v�{i������lh�)O��-V?o��`�P;b/<���P@��\X6�������\�	��ɆD�I8g��	u���6�u�=Y���=�f�I����z&�  ����� @-���7��{�K��;�������W9X݊��9f7g�y����s�, >9���ޢ͓�0��S�DG�#�3�VIͺ���%߇b�bz� �Y�k���n�5���M�A �毸f$ 7�ܽ�I��w�e�LO^�cĬ��\��f��_�_ݳ���<"���R�e��t ]RE��K���9ی���j�ޯ�O���l�Z4��{���_�j:p�%VGj��#ݻ�@���]*n͝���U�KO�ă�����ٮ  ��9�}��f�L���k(
 V�Eok���v���e�����Uj�
�5��Z��Y���VGTE*%0�o�9�#m�S�3����RNM�zq�{�)����&xDu�F��k�aD�@�Ysa��۫ϛM�2Ύ�XɈ���;��2"D'��M݊�Ͼ�W�~j�v�*�������\�3W�3�~;˪6|����>��h�����k]�B@��]S܋��N�F�Y�^�C��;��H{|�3S�1,���� ����L��(�����s6���	?�SgjE����:oWJ���sݝœ��-��i��8�o��3�ǹ<Dē=��M3��OM��6�0�����P�ü��=C�GI�^���4���E:���s��{8uG'�fn<�.n0c�X�x}8""���sQu��ұ+7��u^��Vۉ��	DHH8Z 2�歵5Ԩ
d�cL�c~0$d��u�.U�a�Z��PC`hÄ#R�.z�e�]3�l�'����O��u3�'��O�u! G{�WA^���s��=&�p82]�|s�H���SЇ�i2u��p١�p��Q�}����o�7 �88�>J�=��پ�Y�݃'o{�Sht\��c�tq�у�ۏ:�K�f���$�g��%%������Ǻo�G^���t��9�{��c�v�Ga;&K�)�Ԭ���wx��8X�>��\S|��㞫&q���O7�k��X�;�/��D�7w]�f��ݏF�g�R�N�y�4��r�3����4i�݋�����b90.��y-;6S[ع�M�X�uP����G�4�t�{�����[�mY��>7��=\[�P�.)k֠����٦�$*>��d2C��{*���y���>��jNM�TV��7�x�I"��"��7;�Ӆ524��1<�}q�#�V��Q���p3&���B�ܯ
�aк��=* ?x�@�$#f��z�������Ÿ�՛��oZG�2O	f�mѝ��r�'4v�'�h��Tj@�ݞ�g�Z��C�jV����P��طY����a��$Lz����k3
�>�t=p���^���Z���w�OZ_��m��!8vlάMÊ�ˍ�Y�%)�I��������,țY!9ݘB�Ͷ؆ՙח������F�[6ksa����c�,̤��ma�gb��s,qg%��&ݸز��Yۮ�v�`�f6��mX������V�d۳�';lٶ� +�J󳤈�
��ٴ����#�����6݁l�v[n��\"����f۸�H�f�,��i�m�l3i�3[�[[���Ƕ�/ms�I'F%e�ɔ�U�[^�{�s�e���y�w����,��gR]��fӜ6,��6��$�|φ#;�uA���Z�a��=WK���F�Cې� \�����n�]`�$���Jj��m�F6y6��6�;��J�xy��x*�m��FZ݁�{W�W�{7nܘ�Ӵ<��l�֜���/PI՘"�<sւs���T�o��|��pl�u]��F�8�`�>w?'��6*�8Y�l���y��Y��x�Rz6�e�H�P��m��xϮ�nY����1΍�ػu��6��KW=��#�p��=�׷�z���1�<8 mO��޸1؋����h�p�ocvv.�]ۖ�%��^���8v�vϘN��'s�c)|��6���5Ƚn'��ٸ��0��"}���9Q�r�Ѵ�.�vGѨ����9S�rl��Yی�]����i�(q���q@�{�=*Ai��7nS�q��/:4�����;&��8痝�� ���'���I�V{m=�<�<��s�����AM�ٴu��<=%m��r���=V�`ү�ܝ���stt�Cs���zN-�l�nx�l����+:t�͔���)mx{n�GN������m.��4�]m�#��U�͞���'����"� (�Q7n�i�u����MwSq�Mvu�,��ۜlm��ڑ���*�ڽ�vĜq�����]�����b{�zR��º�n�����v�[m��v�hzۦ�k�ʼ�*���.�u\�\�fv��gu�6v�O3ԛ���A�Ŵ�I�!��px�����R4j��ې3��kxA-ׅkt<M���Kl�����W��|j1���\��K���v�t<��@�g�2��ز����c�3�C&��T;���=F��L���j��(ۮ,n��\��v������N���+��k�q{]����6yB�u�X��`�m�6�p6U0����:�u�aP{:�:\n�]aX�����Q����{1g�g���i��SI�Z�tS�.�3�qɴず{W&Mgt���i�EPs�v4����x�yp��a:�uZ#v��=G��q����<nG�p�W]7G<���!�z�=���N��]��a�=�:Ç��a�X�qyz�
[4��tP�bq�m��u�3��v0�U���5%���v��sb��n-�w9z�{j��p���->ֻORvۜ�nB�hz���R���mc�{v�h�Oaj�[�c۷l�kurC�ڱۣ7*���8�n5vu×�U��B.;:ݛ=���'%;��lm�U��ح�'in����A��#+����=w�` >�����3���Mr�^�uJ�ř��t����ꇍ>���QJU%xb{'3�M�yS��*�V��,q =�r�I$���&�p�	ع�?M�5�g6�J8�n�\�{�= �9��� ��l����N�Ӹ 8w�J��g�f��VGLՀa���Cr��=WGw���s���8s�J� o���n���dۍ�����N��"~�{��ب�*�f���7�:k|��K�bR}잜;�o����Mk$�'�OfLcf��2#��OC��S(֬`���l<������n7h�u���[F��u^o)��MF�i�w���NV�b�b{�xe�T w��fa �}� b�7�:�Esh�.�� Fo�ِ5�rh�h���"��}��g�I>��}�v�c�y�襯����sŶ8j��z��1~YS��Ax=��	����W�f��}��u[� j�^saC��vw��<ơ�4�]5����^����1�q{۫�ﷳ��r����`�*�R�+��{��d>��}��
o�緳Z�����g�ώwӹ�g�-��g����Q:�k.��Jg����T�o��d�ɼ����x�/��G�ߺ�� ������R���t�19�����&�^�2wY��ٛ���a��禰 �{�T�d=��sN9�?�����;��)Ŗ�&�u�v��xY�"c;���� ^{8���ߟ��Q�U,�Ws��@ ��ŀ�g��"�fa��Ǹkb)��0I�����>W�=�2�;�bG��M%A\g�����液��٘�@��� ���9��]zk�JW��z�4HTA�������=ɫ�r_1�r]�Ŧ�^:�Y(���7�8?��B{��:X�Ŏ��xh�oK��>����qv1�&��������|���7���/鮳��N�{��a�{�T���,�E*��	��x��w�E���k$??k�p�=�4��称/6�[#�׮�n������f��nϝN�ZˏA��b$�L���7��M��ڒLv9�� v���z{�k��1G�ŝmOM�l�qF=yS[q�І��K�P�s�mN���+�i�#��G�+Z(�t��FMs����&�$��o=���(O�Y�o&�'�!L56=Q:R�T(U,�A��{� ޷�G�\�z��-�u��  ]�ܓH7��f(1����_ge����^�m�2��P�<��e��}�s �A������w��kh~riQ���v{2���M�D�T"���r�d=�7�;��{�t.H���o�m����2��7�]W/UUZUW�#Xv�:��k�����;�����H�9�M���0}������C'���/G��;��nY�8������KçRG
+7P�a+﷤��i��`�;��u��j�zM$�#~����3�\{o���\�����cJ�D�Å���h�㊷��:�t�b.Q����T �lA���Q�|T�e��=#���w}�̀���!?p]��sq���k�A�I���&h%�����1�N�c�y�� ɼ'{�̎^�kR<@|�N�Ā���l��o�׽~�M��tzm؎�22��σ٩��  t��1`����D���S��Mل�I����A$ݷ阀�Too��E(�i�2ǫ�cZ�{��2r6�u��� /M��Cܐ[��]|�g��>�}�ǯ�ą��5����{rj��o~O޼��+{w� �{��@�{�T[��R?oif�����|�[;�6c5!)�0F���3�jĬ�:SɆo[��bc���D2C�=�WI�~^7�����5�g��y�Yѱi��q�/^�����8Ǟ^n��ou�V��ݜ���6�3��ܝ��)���`:�:ۓ��&ن���v��j潰�`s�۷b���¾
V�l�u�n���v�ɗ���w�S$����%U�v���1��c��c���-�VR�L���>'��� /(�v\�9x�:�%/l�p��:�x�A';cS��fŕ��	��V�1�n4k�<����']�n�WA`��[����]�c�����+m
���s�������0��{�6����X�wH�����σ��ɬA�k�Q�|T�d���!��PAy�w2w|f����@ع7�L���H�lw��c�d}���([����1�N�f|d׻3���H������H��Zy����f�A1c��P�\�+��G*,�wSȑo��]�k\5o� ���i� �=�4�|g==�@w����ܜ�ǰ;=�LĀZ������)D�X��oSIQ�y��Y#��O{�����m���1�@S�I&�WOf1�{n��M�߮����=�i���t��<m��"��a��vᱷ\=�q��M�H���G�ąC��z�7/73倐��&�� s�������O:v�n{ݘ�|;ri}At�ᄒ��ҳuf�����1X��}(W2��G��>����?��"j�g�kޤ�M�;��h��${��ur�����_r��}sw���W�d$�C�{�k�l9�Of(01�o8}����Ѿzw \��R��T�e����w�_P���b� >	}�w������g7:�P>�#zH��z{2��딬C�:�"�2s=5��f����o]< ~&My�����pL$v߶1�����߀5jG�{9A9*dr��p5�՞Ȉ��C��9ᐝ^Y]���N�Rs�i �Gy��ā��7�Lρ��qk���]س�4��[(��ګ��<wς��V��C�P��O�
�7b p���ߧ�]E(�u��ޤz@$�{s >v߶ `��'gC�ӏ���� �=�v�
�܏__�J7.k����a���ۓr�OD^�z��������no~�� {��<���\��p�(.�}0�X�p�J���˘  �o�2�I�_�9����=���PQ��woV��3����x���ni���^���-�����7=:��Y�w|.�g^���"Ӟ��\�� �{s����X���#'�i��Ys>2�r��ftoO����q` ���3��=ɾ���Qt1�x{��t.�� >�t3^h���H����X�O����rh����&����$�q�0���Lπ �=ɪk~�k�NwU�����qƁ��p���{q����]d^��v�<GeNB��:����.{�-nE*,�vww��@ ������$o6�}L�s��]��}�1no;3_(���ƤAE����������u��w~����f�V�9�iQ��W��{�l�t�I{�����Qq��^��� �{�T H<�Л��׷��� �7����v�Ҡ�i�!a[r�b���^G�f��%�� :o���q�ٖ�I���%�X"��O��5��r؞���ܺ�N�Örv`cp�oc4jjnn�)k��,�݉ԕ�uv;�Wx����s���JC�(X��S��f ���5Q-e�vk�6$����u[���Mg��t�}ɘ���4��|�u�8�зU�k�������`�=v�٭��[�x�9ޝ�2u{R�z�� ��$�0�pg��[qWAط�d��4� �iP��{�ǟ�7��絓��Ng&b@ �Ü����[�h'-ndM���E�����O(K�x��I�[�� ܞ�� ���x�s+=y���b��7����|�87m�����5C���n`|��J����˺��w;�� �	��4�����1��&��ģ��5����yx��ѕ .��  ���c���ٞo~�-}�Iz}u�~,zЖ� ՚�!������@$�~�	�L���~jy��5I9۪��8gw����&����g�y����7����[�Y��M�`]����+�4��M�/n6w�l;u5��<\���c!2��k���-������̟F���܍5�Q���6ٶ��|N8;.������wm��v:�u�8�ȃ���m�K�.ݶ���]�Ƀ��B����Epr2nC��ukq��ڸ�v�M��hu�{q�T�S�@�n:���A:��i���c>��I��3����tWni��D��l[�$��{<�`7<��r��/nȔuuQ�"5Ě� v�@=c�^����֋����+Eh�T�M؝n=�::z<��]5zնۆ6�<;�5���'uq�WN��;��H�dL�����y4�$ g��` [��&bf���]�o�Cۑ�|�ﮱ���q��t)���nf��}E�w�{��f�x g�� �oݮ~$�������pz�&I�"��A2�H�E���k� :o��� ��;���Ǭ.��6|s����|7�M`N�퓑;h�_�k>=�hQp�7[��A�s� �|��  ;re�y�{^�{|o����;�QF�GbewW����K rIg��X��2,�΀b!��gD��&��{�T��][���2J1D	Ҡ�@�ów=�Š��㬇�
w^����w�˲;![r�b��z�.� >��&}�A��$��34�oVr�����׵˘��/M��1�viP%i�2�]b=۪op�}�Z��F��{��} ŋ� n{>)�o�f�5����'y���Ekҟ�)�;T���pt>�;�WEY�S���{zE� �O�}�& �4A'��V}���_o����Z��늧t)b2sۘ�> ~;˥F��o���qo{���� K�|��@ x�.��7�%RE*,��5�z����q�={'�^���N{sM���ܳH��}�ҽ;=�E�ol��3ۘ�)��;S��4��8O�i�'0�Ow�S!o�9�}_���y�>d���� ��XހF��\o7�v��mU��G"������X�'[�ѓ���9�m�Mj?���B�����v��=�ȣE��9]��93^����w�J������ ��|Ǭ���7o�` Bx�'��4��GHV�U�d��ˉ`��c�C�m��͒�i� };�4����� �3Ny��Xk���g�*��'-e�;ۥ@ ���>� 6 �P��<�O�Tr��)����m�7�����z����uڹ��J#{���y��w�ؓ�o���p����3�f��E�=,�Nn8yL�GY�>�=��ϴ�o��d�x�<�x3x{O�8j��
��墇cn��]�Cª���N�W
�H���[SU+rǘ��ʷ�<G	���6��,��\d����S^�\�_�n��u�u��r�Z���w;7m[��q���T��1��J��ɒR�SW�&*r���q� )T��U�CZ��:�;��Q'Q�"M��͋Z{��l�����w�{�cg�wA�d����w�p�]�_"�nBx`��ɲr����dJ��xVm\�N�խ�*����C�y���u�v,Ѝ{�RDc��g�lOٽ��w�Z.�9�o�_'�ո�;���͎�a¿U^Lz^�x�߹��{���ܗcEz���g��`�UCr�EK&%�P�J����X�Obܿj�g���m���i�|�wf�U9�X�o׉���7o.��������1��C���&/ǵ�����,�� v����)�75�M�&h��yF��g�Rϴ�Og��t�&x�����y�S�;����3u�$�n���8���I��N
���B5q/=�=�ГZs���5-��bv����4���^������i�%�ϻ	���'�v�j��>�<�)�T�P�yM㙤`)��;�lTl�\��օ��[4��:��w�|^��<j����̙����kR( B��;������o4��:�̎��Z�fնYe��kY��e�e�k��:#f�ٶ�-�-sn,�f��h�[c����2�̶��;M�Ma4��&Y�X�V�kb�Gnv�aL��Zi���M�N@۵������0:�B$J�m�L�ܶ5�ۭ�.ӱ����6�����gfv6,;,�C��˶jn��f��5�����"4�����XiiƲ�����6ٙ���[lmZ�Zd�(�gh���m�-��ٺ�m�V��2�1#���i�Y�Fc�ù.�gs7l�e�4�ml�Fh�&�nkZQg���مGvR�ɷYۇe��[��gi��F]�7bT���9�h&�Y�s[���� #��C`�C���w��� ��]Q� �ﾹ��醗U8��H����v�W���Nl~=�&�DDG4�DDF�%6�ܭ���;A�����o}�a*�)Qfg����0:s������^�����u roVk����|n{���S�9:�����]n�Q7cn�����9��t�x������0���;m�}ͮ�����!~��A�z�� s����>s����̜�7g�^L�4{�J� ��또_=�����J����Ł�)������6�{��?E������I��vɄ������Ƈ�qw�`c�j7kAU"���ˋ�g�ɋ  ��Dk1���K�M���I�fD�	n{���-{;1P%M9k.`a�پ����-ӄC>@�n��@��绶BI |~����P����Ή�qyi�� �r��D�m�070��0�(a��5z`�j���)@�3Lb/L�{=jz�9�j��[�dѫQ�6���\��t�K�u8��H�>2w��� �w�?{O��Y�1��r�� g9ɘ�@ߏrǧ��������8�{���u���g�j�;��)��*�O.��a�"c������z���H�E��k��ϰ<s�������7���<ٿsw1 ]��&`O!rr�I,��WWxޮ���:����W�^�}��| :{����r�Q�4yse�\�v���9ox��[�F�PWJ�LG�k�>���X� #[�&��c����s��������:���WT����jg��{���{)�o}��v��3��x ��,�@ o~����{Z~@Y�zf��zb�Z��-�s��@ ���L��yj�oϘ������K�L��r��1 u��L$g��?{U?A&�7;E����6��Z��^��S�z�P(����C���.�:)�����ޚ�OJ=���0��LZ�V�9bK$��wa� ��0*lR�������1;�QO[q:�wC΍�鴆�wg۞x�a2K�u67X$r��n6��^���Ԯ�6q$���lEN��@�n�f0t�<�p��)�Z���$-^G1W��[N= �4�k��t�y�d�5�!\j�n�b:�N���n8�1�c�J�v�#d��d,���5nC�;�=q�c����G�=��{X��v�5=7]��ţn�˵�2slƩ�
�=��'V�ci J�F��s�a޺��V��]z7���@ };˪6����ǁ��ٍ%j��;�9��&<"6����t��"�f��\��G��i7��0�3πGgyf� ߽s�.M�nz��M���"=:$9Tj�LԘDb�i�Z$�O��&!$�z�}H�z�'��Sm�p�&�������^擣E���;������>�2�B	'��t ����p0�oݬ��M?<�f��֌{&��u%b:����06{����DT���@ �޹���ɘ�J�{A�gY�孋1���d��v��F�l�{l`Iv4[�.���q�Q��q�k|��-P"�й=5��A��� ����|$��˅��4�ĀG9�\�3zf�
�V�bFOw�>�H6����������f�}ve{����K5�C�����{�h����i;0���')`W9�o3���i�<6�39�}Z�ne�z9oh ��co-�o�1 U�-�Y����M��U�E���׮`| t��4��x��ξ9^���u�9�7�]`06{|�πS�q�+lR�(�ˁ�z���Avy��9�o����> ��wɘA=��8��=��Wՙ��TZ�e�܏Ưf� �ܺ���>������Ko��I�|}{X B~;��:�`��o�ײ.�{&���6^b�>��u�˼I��Mƴ�%�MыYL�)g:��2���T���/}˘6���!$�ē�ߖ�&w�{y�[ߟN��y]���s����u٥F["�P��#!u]Dz"T�]+8�ʻ�j� ���{ɬ@ >����g������h�y��r�}Y�=I�]B��`��2w������]*6|�7���Z~�V����Ō�٨`eS��r�RT6��m����k8$kd�W������5��}*�9�';�����~@o�|3 �rǯN����U�E���׬ɷs9�����0 ���r���z�x�Lw�dNkN��s�g�%:� qX"�:5r��ңg��{�>���go}�%�Bz�� ��<$f��&���.R���h���`Ϣ@"]�ٸ��[��,NL؃=)2�v3��G��m�����PUE��w<o.�b�H�����@8L��0tǵCި�S�)���6s�T赭�����T�&|��ŀ�{�ܜ�h���f�i����,�6#7�\ϐ05M�kPY����s�x�\úV2����� ý���	w�\�@ܝ��W����� 8s�J�@|��}sf��'-U
+F�����j8��u�{�� �"���  �yۧ� >~��ڼ]sg����N=޸Y�<�4�N��h.��^�,�U<Vz��x��'�K��2���{o�h٘�+]owB4F�;�P������5�J����X�*�R����z� ӛ�Ł^�����8ǥ��� }�;u����3&���zxC���}kQGj���I#����:�j;n�Ѭ�����:ô�M���+"`8sk�����n�^���z�� >���x����o�08#��䇵�s�w��M���0��n`{K�Ҡ"��-��ϑٚ�Ń{�Y���q�@�����6}�w�ǀ�s�X���o��wǣ��ԍm���k��c�Z�A�w�O ��&}�����u�wKӯa�۬�� y���|��s���@-+��+-�K(\zvg�7����*�^�w\�ϐ��\K ��rf �{�Pϣ���x��k����\�Q�UT��Պ,ό��L��rFGj�{�����=�x��y�3� ���5G�`��w�3S�Z)8�	����&�^��\�Nhn��	6���?j�l��ݝ�}狼3}���v̙���o`�����݃;��v���i�x�=n��9c�*z�ີ��➰'�ڭ���1՞�N;vf��d���]'l����8�^(��ǩD��iq�p<����]�Zڎ�NtC�����������VnI���Z�t<���nn5k=���\r��y7X�۫Fq�6}	��ٸ�K��
�kz��[�x����˱綼q��n��M����p �#n���m���W���S�7[�L~q�}���,�J�9����s��;��3���$�k�j�ow�o�w�3^������y���TqX	���q��4� 3F����e]���_`؀��rf a�MQ�7�M��x�Sg}n�������"V�m��ϏN�&%����&����d&��}��� s=ɘ��=ɥA>�-v�mr�eă��-�^뀞� S��ϖ���$oI�{�]Y��m�g#�l�ɬ��b+-�K(\�d<��#��}VZ͍�j���虾&=�Y阀 �9ɪ1 g=��g�|;��z���ɾE�ě�EkPaB��nwa����	�n�����jۑ^p}}}���]�V�o�5�LX �s�IP����>^�C9����<���ws0 ü�����U�e����\X߼�
���n��wH�Ek�gۚ�MCu���nT������Q��lܕ#�^�<�S�ͻK�yk�A�+ٺ����j{�~@|rM|@#7�\�`j�ay��u��O{^��΁|�Q�:5H:5��3&���s�MwW�����g35��� p�&��H����k�Ԥ`�p���L;7܏�sK]��yo���� ����I$��������~=ɢpU���%
�"ˈ9�r�X ���pd)W�=�Ա�M9u"" G.����s������9݆��S�ԍ5�z��ӹ�����>�h�C�{lk��t��ъӾ��FR�El���gg.���}s ��s���A�|�o�˓ྒ�b �}˘5[�Q
|H�փ�ɥ�A�6r������ ｬx l�95�w��d�&����ďs}����%t$�A�k�O�s����}��\i�*s9����n:	Z�Y����%t	ճ�3�M􉘧��<��Y���Z���5O�]P׹�?*n �>�aٻ���Q��g}ۘml�94�G������͓�k'��N?w�X�}���T$���ҝ�O<u�|D^o����>j����e��]5{4�7�\�Xךi�2�p�Y�0�HjR��s�Uþn��uD�N��"`L#n�ł��lm8%1m���yŮ��n�ƞ#��Xx��LL�1Fjj"Fw��K=��p�_��>�}H߁�wB���y�?wo>x3���g8i�o��8�[lwO���&2�<*�{��[����O9J,�N>�p	��H���$�&;��TL	�DM��y�H;�*�� �JY�-̎z�%��	'�:9XA�n�$�M3F�&D���sM���GleŒH%t������w.��d���!^������D��;��d�ˢ6��.�vFF��rF��ʇ}%�	J��^L���a�U�%,�n�=�e�o{�������[�7G�k������j�G���n�m�s�����;��#=�u��|p�W@����<�Ozd�#�g�!g�FG,��ԙN�W�$e�n�<cj��cmۙ����s�j��}>uЃ����ޥ�m����m��|�<y���J�Llf�H���� �p�'�?)��4�+ܓ/�̀��hV;��@�H:y���|� ������w���9���v�棁K����^;��A���HQ0�p��Ժ��,�N��E�7_<�	��lC�&�"&�f{:^�em����Խ��ר�I֛����J�-u�����_�_u�H�RWM'}}����p]���H���qTI�E�K�o0���[������P4򛥙1G�wKql�BnͲd�)�n���a���e���ݝԆ�g����v x���J�W�\�?e�
R����,��ݙe���cE0�� �ل5���A���'\˹u	f�7��Jض���n��Ʈ3k�Ɏ&��y�fn����̈́@�����O�{ѭ�T3�/{�3u��� ���~�T�@qٺm��JT[���&�5��~�	�� ��
�f��d�Vb��&�XN2&୻Y;�S�q~��ZS��`�B;rz�4$��w���S܌ʈ�Q&�a�����UeA�s��dX9I����;�bT��QC�9Bs�"S�574\�=f����DJ�I!iw�)������S���Lb�!�p�T֛��9�l���/q�Fw�{�N�����	=�ޖ�
ڬ�I���Zq�����7Wi��e:��cVW}��T��`�1\0�`y�۠���v�r�[Ԫv=L!_y!�F�.����|�ԊjZ�p�|4mTn���l��Ä�x��z�R�v���(޵ FwwlN؛y�iJ-�$8z�O0�v'���r�<�ٲ�a�nz������v��(E�N����R��n$�g�O�Aˍix�V?�Hw�o����H��;(��x{�5!F͞�_{k�4�FqJ�;�}Udb~�2���[����v�n���f��p�}^K�Jؿ<i����^�����E�s�A8J������w)oVt[*Y��������>�V�ö�6٭4�#��J���ҙ�jl�,-m�l�DedNr5������F��j�VpR6�����2Y�8�ͬ���9,�Ŗ[n��%��l�Xٚie�óF٫m��s;3��Zɤ[2[[6l��� ��n;m�F�嶍c-��&u�mmN�Ցf6�v��ElܛX�쵶�22̲:-�D�űE�ضЊmh�$�v�N:�ku��n��dòGl�(J:�m�nD�X&�Y��5��-��[��vZH[g8@���u�(�'5�m��p�ca���s��D���v۲�"[f튈���Ѷ�d�gm�Y2�t�ڙgXgsl�;s�kq�wa�����3I�d�ڊ3��2�4�kl]�#3l;�Ҕm�:Um��_ƞ�CRjkT��.�:��tCnm���m������K�h��w�x�i�]�m����q��Jq�n�����9m]V{:���g-ֵ�NU܇':ֹz����shݤ��on�6���q�vg���uoVs�cu���,���&���;rw2�r�k=m
F۲.<\��h[v�˼�u�{v��A9*c��g�nN��2;:�p�+n���8B�mƉ��CΌmNr��L�6�RF�Q�k�n�38��jY�g�-��䛓��Gmc�|f��m�]�yƯ3oc\�����ڄy�u�F�Uۛ���NanظO8�gڢ���Yw���v
����K�7n�٨Q�Y�Y�i�,mݵ{4˹��厊�:�x�����m]Y�u]n8�7 k:���x
�vHܝ�ٔ�ڨ��mu�Y���uK���lH�<�׵\�{j�l�S�Ӱ������`���\�b�z�|�Q�v����wr^�G	�����Uܛ��\�-�:��s��u�c%�t������oh�2����Ak�{O[n\P�T���"iKvr���YKm�޼��<��bxwp��ֶq�l�s�nXGd3��Żh�Gl�z��u�g+�]qg���]�{]�� �&-��4^�6w6W�bN{M�O��ѴVX�1��X��M��W�̜M������I�\[L;�>0�I#n]� �!�uH��g�9
���]{@G,��5��sĴ�$��A�g�R4��9�ۗ�(����ѽ��s�U7l3��i���/i����V�Q�'vZ�|�p�9�br��h���L=�6,-r�ݔ��c�t��@���v������<'��qr���V_�].ٹ綅�Ͳ�f�}�I�#��.�9f�w%�ɂ�dמe�N��N���r��9��{G�cZ�h�W]'&��<�� �1��Q��۞�g]�jsOkv��̛
�n�cM�/�j9��[�\7NU3���y������_D�gqE�G���q�o<�m�x�I�s)n]t��\�l��L�rg�
���t<��K�V��H\P"��<u�x=�ڎ��\�m���Mnқ,����l�x�z썞�e-�Q�H��&�&���r3�l�gp�DqtIu'qЧZLs۳��c�fz�V�lv��U��]l��6��sr����ɝc��q��8�n�m�λ �6M��W��q��@��b:[�����&�rW>,RGTM4ϳ��"����m�H)6��F���w3C��td���o0���B������z-8���;���آO�{��g�ޔ��;�TqA]վ�9=�K��#�[��d�WYb|�K �ބ��>$�9tzOne���9wyg{��6�ߧ8k����K��ȫ+�.�<���,�`㗜�$��X$㎠��w�<œ����x.�S�V�*���ݚM���J��2ᮄ�ǘ�`b�y��O��(�H9�4�{Nz,��.��i��9��m)k�5��C��\���0�O"U���t�8K<9�7�����K,��k�'��������pZM��w�Q�P�kR.�L��5�ل����(�aAH�D�1"���7�4I\ө�g20Fs��6f����p��=Y���EC	;T,���mʐŕ*ہ'�$*'�����<O�=]�E)��^q坙����>A$�T��I9�>��=厶M>�vfo�����B�X�UQ.4�V�׈'���lʎZ�Ė�o�����wһ��L���k"�|�rQk���M�I��B� ���1fu�gd�$�p�͂f�:�Ɋ5�S1QV�4 �\���E`X�ou�y�śW6}��� ���f����;��x֗��_��K,l��F�r��ùt���V-�<�[Ga�#j��n�{ߗ��T�1ʧt�y<	$�B� �w+��NM
�<1�x�w�4�o�9~}�䥖EU���F�s�%��`�22]����|A[,����>0tv^mAz�]��v:jl��`�>r�;�����m>s��%�&߮Ψԋ����ʵ��ګl�3t0�Qu��)�Kjn��R��pCD��I(9(6�F���VdOFe�y}u=�'������A�
� �3;�0�Sf�VI
�v���{g��|w#&��>DNEЂ	���`�{T��z���O!����<?0���k"�����'Oj���n���&�#\�|���'Ǐj� ����-���b@��^��h)��tq��]��m�vo3����p�s��3|��ew�+!J�7�6�z�;��$���6���Yu����Vwm��k��T���f�����}Ő��ӕ��	1��I��"���B]B�)8������"��K4�绬L�+� ��x_�<�Х3���Ϸ�M��h��f�2jH��������X2�n��	;� �i��C�7���g$#{5G���$��^l����'V6�J��3-ZN�`����;r�dFh�-�l>��qh�0������
i�:!'���v��k�ouy��b�@�а�$�'�N�I'�u�m�%.'�w^o��M&���_�g�k*���J�kٶä�ϫy��y݂V�t<�L��	�N�<:�9I�����ZQ��E�>���,{}�&���x�3EśE[q�Lv����'Ů�&���vhc+�8X�u=���Q�R��y��f<$�;Sd�K��Apo��5+hvįf������"b��ф�f,;��M�׸r�4�OzY�Dv�:1]{\�lu��4Z��SdU[]�Y�g�����r��x���H�Ol�D�m��-M�T�������6��~f��mI�L��7P�o��w�,c1x�Q��}'�ǌ��d���P'�ܷ=�e�է��:��tш�a�R�z�'��ߠw*�>A%�f�l���+U�0�Dr����㴜��A�sg��o�y��6�1�H�+���%���U#��p`']v��v�L�%3m�vKͻph۷$']�_��5y�99��;����/���qO=��Hqa�ۆ�n�$vܱQ�W���<��^V��p�ļɑ���v�N�{U58W���{vչ�������}��c��89:ܠ��;��[s�67������ͥ����v��I����g��Q�/�������>^ۡw&���Lv;n\��M͈窚;S���g�+n�F�|]^��%uUPl���	�':	_s��h�-w�YC��ZMo�)8��%�-dZ�V�,!s�j,��x�I#vQ��o_r�T��߬�rw��euIPf�X2[�$_7�	 �Gf�n��:	��u	�.��ĉ�5&*�"�VYW�Y/�ƻ�I�=�d�A#w�s	���q��r	#����պ�I�V��z83�gk�e��m��
� w"�]��.7���=�Čz����Z�R�kT��)�[Zv��V$p��n�l;K�3AX�\@8{�Y�=���#����s6��%�0�Iq������3#��"o�[Mo����;��bM�򫊎GQ+���?k U~�m���L��&%Z���p�]ޗ�i�r�ʨSӘ#V��ښ���v�z�Ϣ��2�����"D.�VtdM�$�����$��7�va ���"�sq�|�Xsnc�
V#����K-N;Y.L�s�M��ܚoჼg�3�,�� �߻^�/VV�!K��|���������Y�J�ݘI�cyM�Gϣ<����ө�S}�g;��jwY��8Ueaj��'�d�H<�T�r�f�'Ԛ��A#f�ɦ�m'��f�5�� }8�Ŕ�u�Xw]b�v�W^-��-ֈxw+;����<�W%��eV�g�}�f,m�׾rkĀI-OƁם=x%�Y� �o)��M�Јź����r���V�	͹�۞gZ���Q� k��M�:LlM�p�\U��-oK��f�m���Dk�m�}t���l���U�$���"�f3$98�7���&nam\0Q�9b��o8}�o&�s��8E�q��.z����\���p[�H�]`!=�y��oۚm7��;��<=��ju�bFg���%LZ[��f����l	��ƈ׹�:��q�_8��jm�/o++T�Yu��=G�o^�����km�0d>ɰI%�DQ׻׀���wF�m�[��#����n�{s�V��rk��P��]rT��굵	"�=�w��p����w��d^I���7�{�oو�t�,Hn�9�joĂK�T�2��MP14j�jl����9��1N'��8	�V�$��ل����TQ��}{_k������hXA(�3\��6� ��g��w'o%��\]�\� �Q4�[�oٌ�T\UYk���[�^���=�E�Ǐd0I��PA$�Y�0Y���4�: ]�6U���¥ҎShL����]�}��"�2�f��[�J^.A�-�C����)2��{/35� �~�	�ϵJ���LDb�<i�V�ܐz���?
/�s�斉{�3�tL ̲_�0����+j�.�u��S2A�j�P���`���f��:ָ�}D�n6��T��T�1��U����V R�0��|��;~o�w��ؼoښw5 �}_��?Y�y�� ��a�+�!,Rd=�׃�����ԏ���~�ܳ$�o\�$�=b��ȫ��3�e$��CRԞ|���������|�0��\{�	�[k0|H�޹�L{��صf�F)0?�{Q�w��$�FI �rx0x깲Itr�G��Sn��&��{y���*��v��U-o_/�lI{^��73�^��A`����I=�l>)�TO�Z>��i�HT�Wx>r������۸��R�N+PK�I���v������d�����]V���t5ݓ/Q�* 8ޮl�����(.��:Wdv�x4kf��t.�!۵�2�^��\ 㝻��mоGqê��<��cM֋��&��(N��a�i���<��ص۱��맛�yc���e�ImNL�!ti�m-�n�``!�n^�[9\v,��v� q���x&8��㮍U�nu�"]�<�xנ��y<W;my��'t�A�6�\����]���H	=��Q��qk��6��:�=��OEiň,Gr����d`���_�tq�4*�+Fe��I�Փd�j�! �M��e�O��Cs=�4rI��$�}��&�A)�;��<7��~��ޘ��{$iX�
�f{!v͂|HzE�jFn��e9��$od�'�'��&�!SBN���������W���1���^`�yG8�Y�1A���9i��e�"�;&�f�Ϳ"VF�Q����r&����Ύ�d$rT95�����Z�$^�v$	�Y�3C�.���0�p�I0$T]m��u��rJ'<�T��Z)��X�nfS���vz+�~\^QI �w	{4������M���n������[��ʗ�[h{�'bm�t(���(Ш�y�׸�<VGs��DM�o(EM�ܜ���u.�):�,�L�y����:;���������gN4�.$u�7܀հ���Kr�ظ,6�`aŒ8��'��r�R�&OO{Y��lD��bD��*�I?h������=�ϱ��M� �tũ@��܂	Y�3<	����1jMH�5B�=��g"78�_1 �.O��#1�fz7�v����r-�G������rK,	]���uşy�d�;kb^'�k	�L�E�I!�� ��M�SM�N�urE�ގ�2G�T�����l��[����jӲ�&�)�,�GUM4Ϲ�3���S"�����5ؐAx��	��ȱϡ�r����[j)ߤBξ�s�Qq[Km��Z޼]n-|��Z�eq�r$nm��|O�7�l�Tvgg�s�}٭��!iZ�T�X���x�&�ӽs`�|u���Y�7,���F�oȬ�̩������ϧ`[�͝篙�] nL�y9�g���y ����n��j��z�����]k��0�͇��e�"b&o7rjO^��&}�ĿKQ>��w7�.�}�x�h�r1�Bq�Þ��÷�^�4�圴�U˙[b����d��s�8_6���#:ݪ{��K�h�����22�Vr7�v������\��h�����>��]������j�.����B�P����W.����.��Apv��$��[jm�Gn4T���������s-
r����1�q"ǣ���v���yӓh�����X��3�w����A�2�fU�ʽ�c�!�/�f��Z�Y{L��{�}����Wyب����H�83J�?\�.�b�Y<�]ړ���y�:*b�����>�¥���.��5Ǳ!�^t�����U� tc�R�-z\5n����0O���%�)�#�`�s�81.g8��Z�Z7�=���fT���8hֲ`Wk^����ٳsfH6O$<Ӑ�[����E�þʥ;���j�@N����}̚����������'*����Kw��Ǽ{�0�Em��}ʯ�"��SA�z=�)>�݄�<Wo���[��=X��+�@�+Me�)�;�_sz�K����<������Id�֬ȁ2kf40��Kd��[�{w��틺�b��caUY*n�6!ߵޫV�;G-Ō��6�*�0�vS� ���Jj�<7�Oz�xg=��VA�x96�����W',��k5>�I�Clm��6�4��[����lIIp�d�Z�ձ�+;E��e�u9HVؙ�(;49mY��tYm�8
JG.ɱ�iݘ���S5�C1�l�@��2�]�i���7!Y����+,2�-k�m���lm�9�h���m�m�[jGI8�\[v��Sj�՝�m�噘����≑f��H �pve��R��6섄���9�l�NV�J-88�J "���8��J�AV̝Q'Y��N9[c���m�E	r�e9�i�t�nУ�(�8���;;"qr��ȧD(\mh�3��(	D��:��"r8���rB��8��f��I���Y,r��'9AI ��K1�(r���r'ﯷ�ϛ�w9�f6������jd��vPIT�w��gY�\s	�����> w��/���95��}A�ZV����x�ʬH9к���U
}��-�Z�f/UՂA	�;f\�~=���_���<�.�G7T1n+nQ�덽gl�6�K��a:�H�*'Q��ߟ���Jꢪ��y����ڮ����Js�,ܹƅ��}���`>���p4x�+wp������o�7��Oϯݟ��A�׬��w ���}`�<��\���S�\�v��d����k[����vyߤ��հ�ӑY��k��d�B��E�]��@�q�&�I�TE
�9�.�nD�lpG$Y�sd�H$f�tX$�|�w��b��A�M�.������&EЙuQ��fڌ�΁���Օ�)}�����<sV{��;�	w6Aҳ��i��RGp�}H�}Q��i_MN(�K ��J���-���w��tRP�n���5�OE�`��;�A,������g�o����IjC,Z�j�]k���9Ck����bcp��R�X	Z����X
QR����M��Μ���{�xide&X*�*\�I>=��,(�;F�(�AiI<~������c��h ���H��0�_-�Qf�Js}������)J5t���"o��g����-v���1�+�<I��ǀe���=��$REj�R��;3��o.���'��~$=ՙ����'36s�i9kSY�NG\�V�U���Ń�:w�FZgS����ułI����A=�6Fu��:���r�j�w��$^�����[��=ٷ�q�`���s��"Lĭ�I�V���qDd���w��'�T���хss�?^�ۏw�~ִ��^�8��S��qI�����{S��m�s��b�C��������{ �t���k��w;.v/𺏄�����-p#̫n�W+���qY�b�	\�o-ۧa��m�\Y��d�b��P��C��qֶ�6^N�h0�
=��v8�]\Es�s�:k\�\���&n�<]��l�s8��\�N��^�;�r[����v��Q���l���Ɔ�];mX��'&o��&�Ϣ`�{<�),U/����I#��� ���d����y�r��7���L��e�AҊ8	�}t/��Vp�Xӭ��D����`$�{Qi�^d����l�Ox߽�1�8@�(Q����)[���U͐O<W��^_)�@�3k` �޹�O��J5*D�LX:�:�f/����<O����$����~���o�"�@o3�0�'m-��Uk��E��y����Q��ɷ"L�Er]��IQ��,���~��ϒn����o��N�e�
�BKkM�^��;��<�[,��qwIfk��\�3ê�'�����wK���52_x������7�I'ݳ��.��\9��%�}����XwY�nK BJ���oIF��gW9�
k3�\Z�tǯ������_�ß<q�1�0,r!7��,p��y�6�NWs���U1�o1H'-p&�z����N#w�M��*��J���$(�s~ ��9��GK#�D+�߀ʾb�#t���BL���������·mT�a��۝O $���M�����Q�3�!��;j���NX���U���I���X$��O��v��hT�fl1�f�>�\
�2h�fq�bA�c��͒K��w�F�M�H;��ă�B�Ǚ���x�y��u�&}냊8��$S�]�O0|�b�X���M�k�R���+j�F�ޮy9im,�*��]�ZM��p�um��;�n�95=�C��l�R��O�ڞktj"�����&��k;81���	�>�q`�WV<�I,d�늫�כ߷g^�GE��-r��|{zJ}�X�a'�%e\`m0ff�����&��s�ӥ��*���5���������WM���Y��w���w�T{��Хq8�>���]��0�[-DGX��V�w�ĂAN;�A�+�g���:"�kN�k�>g�}��2𾆻�ڢ|���Yٞ$F�KøF��A!�5�_rL䈒H�V��t����m�x�)�m�����[D�NtX$y��aƯ������2�gk�c�Ù�֮����O	��6��݋���\N�ӖK�l��n�����>���4o��6�ˏ�\mt�4��j��w��-X�A>��s16���i9im,�*�K��E��`u�]�T�csd�A8�a�z��%N�P�9-��q��m�M=�BL��R!n��Z� (�=y�`�N�F{=���c|��f&�k�������"�d	B������20Q�lm��ՙ��� �O�oK���q�D��R2"��ml����Wxc�������rpa���<R�\n��"{xMu["�_[�{e/s�Ԁ��ކe���۽����{_;�K�gDDĘ� ���2��$Oj��	(����u��߉��0����$�����q�:3����%m��z��a��n�\����D���q؛tNr�I�"~����DI$n�H��}�������L���n�����Ђ췘�\ɮS��|��N*����|j6o��s��V����0H�Q`�Kޗb9�z��UI_w��l���U4"$Ps
�|H$������7������A>��I{�͊k'��	`Ii�&?��\����`��i`I����><��ͭ�Q4F����^4�$ѵ�R�K.��hm�����a�����fm�+b� �J]� �t�e�g`>fKP�&*fC'�o*�ּ[3�g���}��V����K�+b:���j�}k*��rm΄1zq╹���.r��І	�&�+�WU���!���;�"TwC�U���㭘n�n��v��D�� t�:v:�=)�xM���h�����H��Y���0xd#;M�����p�u����������ȽmlNs�g�����Ë�+�&M��7:���'��{]&�Mqq�k;;k2��!��x�{�ǀ$���v�]���yC�\gnݱ�:�n��sѯv�9��&��nq,�9�g� ��%ؙШ�nT�"��Ԑ�?~��FZӶ���龚M7��{Hm�׻{�Xd�h1׹�`��w	$�s� �&qL����j�����M��[>�2�����f'a|	:��	�<��a%�zd͎���x�
����H�n �������{��H"�Eev��=�{��IԻ��k���gϽÕ9iU��"�^��e�,�ڠﶲ ��z���|k�k��˻:��|��?{&�������
Hn� ���`(��x>�7��7ገ�Ϋ6	${�v� G�����y�c�W�^�i�b�mXۂl{v���q�qv�^�Q97c9�����ǵa�]����~�KAT*�To�^m<�������zi�R�������_�:�;.Έ��5�T�.C��ǀӈ�����p=߆n>=�n���A_x��%��P���4�G�㾯ݵ�bKޟ���>r���n���L�fu�r��z�x��
f�3j�c�S} ��v�Hq��d�|���跚3[��9nE!$n�(�eSy�$q�S`����2`��F �� ���_ۏ�S�#	� ��ꢈJ�D�5IT{�v߰�nl	/z[��S[����DK՘H琴�l��U$����M&��zwDS.���5���&��� �Hq[�d���t,[�'Z��8���ت�n����(��r���<ε��qt?�ߚ ����V��{}����&���:36����5�l�Oo:⌌�J�j��y�����7�}�5$T�TT��SVevU�A�P��,=C2���A#b�͒H=���kv�M�1/+�,w���.���lrH)/��S1a��Zm��d�I����5�g$�ק�}[��6l������#�7��|Ŧ�����qr��*�����׈�=ƣ-4�$.�D�{
o8�C��6';�t�K&�AHI��;.���}��C�q����4������Ő}�Md��*-�.'��_ێ1Oq�H�X7�=�A{i��uV<j�S�Ƴ��=s`G���}�M^ {�;T,VE�v9�g�f���}rvθ�2��W>�KW[�C��i:�y�ȥev{:s�ʭ�9%�n��~�u`�I;��`(��5�b�U�n)�H'�6�X��xA���UFd��ڱg���o`���Y�	�͹^�Iu��$�oSY��4eEi�}q�&u��#�h��m��9e���]6�y��ki�ˇ����ΖI'u`�	��5�H���$�D�ҙ��zd�3ҽy5��H$gV�H��I�7�={Y%�c����tV޺ᕙ6��������(N�kܼ�5Ǆ��]7���«V�y�N$�tQ!�X��8�5ӻK�5�3�i��s�O'fA�N�*��Ma �3�l��Ӂ
����&��� �_H����eS1Āmc�[ �;=(�\ɷsӌ�v;XJ1��N��u��Lm��χyMM1�z4�Y�Ս��{Z�a8���zUo:�)U��k���gɿ�{�p���m�Ic����~1�5��YS:��*_B�un�����H�8��|Tu9��WR&��BԊĒ�I�z�Y��m�_�0��y�L���ʾ	�<�{=�q<��ڒ��ĵ$t�! ��s����ݸl+���y���|H�S`�O��tS|�ɹ�;��V�ٙ�n�xH_��זo��Gj�N�֤�������%��g9��$�	/�@�$��$ I���%@$�	/�H@���$�	/�$ IpB�� �$����%��$�	/�H@��� �$�	!K B��$ IpB��$ I`B��$ I0B� �$���d�Mg���� z�f�A@��̟\��|,�G��E h h � � 
B- V���TH�
T
 ��ڴ�@� PhUP��)��G}@����CEAB��A�JV�U 4��)T�@  ���E
"@Q R�m�B�(P$
�                     = 
    
                  ��y*��PQ&f�jh���ķs����8�jE�9�!)�]���킜�D�� �U�suT�n�[@���
KO   ���b����V5� �J���m��7-J�Nf�'Z]5J�� p��t�ٰf;f���y��D�ͩR��
T���  �      �
�*U��]�G�8�su+��ז�Pzn ����=j�g��wJ��޷C���� �ѧ#/OGxûB� )��   ��|�v-�;��Aָ ����i�sj9�l�LZrt�{� �Ь��OgB����s��d
�u��@PP�_   x       z x�N�t_X�rUsuA^����q˼ Lۨ��rt����� 9p !���Tu��@ $�(�  >���HG;tY�`ܹ�`[�@d.�;�է �`X�&��5z`��`4)z��X  {G�@4)|  �         �(�9�w�( x��m �` =�t^` 㸠��G6+�e S��t��@^���G����� �;�Jh������EEj�  }|�=� t��9� \�� x�@9�T���J�u��nwu��� �TY�@�å�ۜ�;e�R�� (QE/�  <       ��%�Nm'cU.���)��j�5rª'n ��]5�j��-I��W.�T�K��* :��s7kj�.wT��@x   '*���j�i͝iQkp .�Փ����;f�S���m���vԦ� 	ʤYj%����j��H���"W���CE)( ��b%*Pd�����UJ3R��  ���R�4  )���Q�0C&�!I�
�� 4�&�S�w�O��h��|ӎ���C����>G%}-��B��>��?�$ IX�		�	!K�$ IB�HB!#����{����|���G_�o?_�c[��!w�o%�T.��hQ#%'.��yV��h�W/F��ٶ�e�M40�1��fI�3h����m�X�.�"�#��{���-�6KWM�����x�+z5V��ov�M�[�¦v�8�&֫�h�N�놭MܹLw�i�7���8&n21RŶ���a�M;y��-�.f�]"��MZf�D���Юd	e�2�8wn,�ul��Ci��A��u�CK�.e�ұC�6�,ѭ���B����RF�C�lhѕFmGY�E�q;eHF���f��5��&�!����RB�"��u�
ݻ����	c	�
S(��)��+v�X�;����FK��D��l��
�C����d���tR�18\�s�0)6�! f]��~X�G��ُ)U%�-ЎP�nP64C�jĬ�A�WX�6��!bk�&ۙ�s8�o��J慇
�P���N[���އ���<�ۙ*fk�,^X�ň�����]`KC(�W3-�����j+.�Ub���с�[V���U%���N'��a��F0f�l*4-��j�Kѭ�X��j�rf��y�tՂ����q��D�Ɏ�E��`f�FQ�B�'(b7�t���[�B�%�o>e������q�:Ӂ-�2��͵��7�Y�����YN��G, 7V��N�4+�P���=�Hh(�`��i�B���M�ܭ����ْJ��.m��*�Gkڰ������`	X�ӎ�)U��V,�{l[�lP�jZ�M��-�Wz֪�58�נX���"��n�̣���M�f�#q��kҼɊ�+�J�tT�Rn�-&rY����	���`A��d���҆n��2�<j쩼V��昩����!��"��s.��sE^�ԝ-uef�Jm�Z��2��,6޷G#�'u5��b�	�Ɋ�H��9�*L���ظ��nn�ݼ���Ȓa����q<�wy�WH�U�o3%�&e�t��au����v��: òP�o��U�X��*nҘ3)�R�
��
3qija�0$QW`qQG�6Ƈl��^,�N�y��iȈ�&�M���Y�>S;
�g�5{%������7@Y`�Ib�Ai�,a�:��xr�I�c]��朕�l�ڐb+(��Զ)-�������梷5N+	�Z�Fn`�����(Ff^�Ե�[�X�&:ݏv;�j��K�V���N^�^�g^�o*���y	�]�E*���TJT4mKWaL����mj���e�� ӺY��,Z�kem��$�vv1�ߖh�*�b��NaNnZ��
�QfӺʰ�4�4vv��[O��A��������ܣLGe��[h�L�+���+`"�k�"x�2�e0��ʻ�8m�Q��`׹i��Ŭ�S�nGf��e[7D|���[,��4�9����eѷ�J�\& ��^�����0ӷ!ٜL@.�Cy�$�ݾ;C���f<-�wt��yOC�6T�F7��9#W�OE��c�cw,��D�Y̳���,��]lZ,-2��~Y5+�6���.�wtJ��,�̔u6��Z�if}�V�
Sј~M2��"�#�wv�cNÙٽq��Mݱ�s5V5�5SnF�qCot�<6%Kf6�^A@S�-݆o1 -�D��[���Ӛ��ۺx�ʚ嚂�n�ř��$�5��Pg,�v&�^����ǵgQ�F�b�lRV��h3�J+C����̄ib�˱K�7���j8u9a'��k����ԟT��.�Wyv�ӳSw
�٭J���k5/ԭ�P�&�n��^fm+z�*6/�]D��r�;6�%�L�b�&i���#%,��1(���::�!n��(2�3Cb�e��'/v	�5A��6C�pr�$7�����
jn	�R�<���� *Vf*��]G{y8^%F��1�sn�B��K7l�h�h\j�i�m�O��2�eRԋҪR�^5F��W�v�!hn��%��G/Xy��F�^^,ѹgr�x����Bl�W�B�"��5V�;��n�i��ؠI*m��-�̩P,��Z��;H�M��ͽ�+Em]��~�����b�5��Yѡ�l�WJ��Ln���(��
�7W)��9r\�����T�H�S��n����W��k0�/BB��$�D�m�z�ScN�!ٕ�֜C�$�m₅K�f̴�0%��K~�]�y
eSڍ�*x�d�b2dR�R�X��s$:�'���)M���{uy�����۬�]ãU�]��ۋt˵V�v�� ����iY���e�� �X����x	�-@���+qU��EBpbI1*�z�&�8�n6����5Yx�ݭ4ӷs.Py5��U�Xt��":����Y�ҡ��ͱ�J�A*�B���Dcʰ]�B��ջ�'�w�KH��/v�HՔ��9(�]źeJo)���f���L��&&d��]E�%����՘%����*"�աޣu��Z�$ ����㶅���m�mNL�T��/�J/+/ǜB�%��F�쭔��VW�{N�:��Q5z�l�{�� Z�
�t*�E�?[����,Y�t��^����݌�%�d��� ��HL^IjۂG���,Y�JBfL�Ę��WyC.j.
^wYJ}���Z!
eҋ*�+$ �-���HƆL�d+(��o!�#2*�7��p��1әN���-	D�Z�cf�4*e��V��%��^f��(;�ӡw��x��Kګv*_�љ,j߁4�eT֮hswRX��q�32��4�ZtלK�)�K"���%�e͘R�ŋ�8�^'��Pfҕ9���r�!��.J���d8H���!Xl�bJ`�l�DQ��ԉ��ݵ2Zj�
&�J]Ü�$�n��d����ֹ*��x�o2�ݬ֥�ٺ�bV��33,� 6]D�ݻ�ib�h�Ū���r�3V+G'��DͣV�sIͧfe��M�W)��?��ص�Y��l=)x����Zw��@Xs2��5�X7.RF<Ǒ;Y�fh��ȅ��M�$ʴ����VL�v2ȈZ�\0���Z`�w�4^nYVb��M�۳zҫV����t�V�]�(p�o�YJ!�����Mm{9��u�&���D�Źi��7�F����j�eNI�0�Y�)�RB�DYXB�-�f��]#�)�����č��yx$(�e�����; N��I�@b�G7L�M0�͑���w`�y(�W��%	b�n+�7N�q�v[U95��fS��V�X��u�!0P�uSr��b��A�����!\!N^C'!5��of�,��ts�%�P1��k0�5��wwx]�s��ZߋJ��ڬuli1�Y��Yڗj3�im��;�p7qV�ݜV�\Xۺ�eĂ&i� ܨ�za�d��olEU.��su�m�YX�V��V�cw޽�@��qYX��	��u���r�B4)��1+
��/�J�,� b�S��r���)B٬�
f�uHM�]�W:��Q�� ��V�����S�.��t^� �-��6wsm��g�f� �w��2ys��b�����X�
�(�%���--���Q�p{B�*������C�U͸j'1K�Q�%0�u�q���֔�dQ�S��A��-�2ݘDeǛ(Խ�`^Y�W��@�t������Z�P�6���l��7W�]�S�Q6�"+!�K��g�aB�IX�(������%���4Y�ӂ��x�rb��*t3b�r�<ۭe�v�|���jS�ʸ��A�)���	yxX���^���6�l2Tq|��.��C��(�$T��O0�X���[KuO~֒�U�,K�u�WBK���"�Q�&�Ȕͤ�t�`/n�]갲�]K4Li��k/��:��6�+��F6�V�K�7!z�iٴ2��x2P�o>���\��{{�n̻�ըi�[��c9��Psv��f5��]��ʚr�"�Yi�~46���x)h�4h�[��m
�p@�m`��%�ݠ\�GL���'&n��S�a3x��`nY���Ī�ͨ����*R�މxv�c�6I��R�[u��4�?��L-�1�Y�Z�J57�2�t�h��N��X��o�xo Ů��77iORXj�\���A[W{�^T�k^<��r�0��%��i;����Zfa^���7�.���³O�����ֵ*�]Յ��q
��`.;�F&�qb!ǀnX���n����9�e�T�d�F�8F\�((a����8��mLY�t�"��7��Bhn�;s&��ԕ؋M���p�(�f�T/"O,��J+iQ��m�c ����[��-�6RwW�2Q��ŏ�/P8���Z�Evᗀ��<*JTvk�e�Z���S����Z6o'��v��cWW7j�{-C�R��\uv�H�S��N��L�p\��*,���7�Yh2�ToYrɠ[�����x�vr�
��x�lg1*�z֡f
B����`���fU���!W�������� j��N��8d��oX�R��6�r�U)� 'Y5˹��)%��j��5��f�H�4�M��N��W�#hjD����l�X���[W@fǌ�tݳDb"fe�Rl�w4U�W��6�\�uF
~-2���Nj��3I<��0mb��L<��GJx"h
nǯ�V\���b�fЫ��09�3!Ǘx0�JoX�Pl`���a���C������Z�

��(-�6�yB�T����ܫ���dA���m� �����̾vE�.ljf�X�i�yp���y8�����w(��L�4�JxC�`�˲���#C�ͨ	����KX6�ж$N�+.�z�y���;���ӄ�8-�MP���%L0[a�c�#�F�%U��X����[rU����U�*/UA&�{���JM���m����-�p��L%I4��q6�̼�4*��&u���.�]cv�����X��f��FI�A�*�]��~�-yT�D�8DG1�Ն��an�ZC&���m���3q>)�b��=��jo�543t!��1����*�3f���ZBЫ,Z{k7����p�ӍӬ�yw-�̬��Ue<�FE�9
T�Q0�
)i�i�s%]�U��j�Nn�d{�H��I���#${���z�\�Ϧ�6^�ww�i���� $�&�ی5nm���O"g˻v-�!�)Ŕ�jm���u�^I�ʮ�`�/7��(�]��r�쬳Z��)�9J���2e[����+���6�����I{�wa�ѡ-��$r���sr��av ߅k�4b�������B�t�5-�`��9��X�R�a�pA�I�����R���檠�lf��ѭMq\9E�-���"h+͛V֕%5�����#�m
.���NB��3kU����w�T��:e��9i<sVbͺ�¨mIF�T1իB������7bu�7���w�2�Z�ش�ϝ6j,8�y�r�k6�n��q���d�t3]�x�jt��Z-Sa�jb� j-�cN�-iŗ�)Yr�EBѦ�ٴ���2��� ū-�kw,��0`��m�i�zd�҂�k�UP�cMR�nl����)b5Y�n��Q�(���w����7EL���[�n�d�rӥ��`�2��kn֬�C�Z�M�T��ԧ�siۺ��u޳��fս�TBͪ�T�p|Q����� 躖��R�X�����+��@ڸ��˰�"��H,���`��͔�;�'w��/ 9z�Sn��	��<�V̉�Xˆ���3�z�u��=?$��a�0�h��KK��b�7�<���fڳ�(7P�ϡ�e�e�V0މ�Fn�H!9�mU]���"�I��twm�Qnջ���Y-8��)�ctnCR �Q/̆����I��xpE`�SPh�qS�ldQ�Y��fO�5L�R2�rhF/$Qȋ4��o��b��˕�e�u�W0��L�2�õ�{*Z�֝b��\�!Cb����
�J����90��V��٩�*\�6��w&��kv�e���ԅ^��:1�Ұ^���
������<bC��1Mȋ�`[� �.���&����w327&R�n �mD/4Yf�#AD���ۢ`b8��d�]��!
��LV$��be:̑+�r�҈9-�FRC"�Hf�N��E�ޔ�����6#ZKӫ\��.�?�ʹz��V�-)�-�slˑ�D�36�S*��̬�:̨���r ���f��TmѨnͳx��s��t�)����������Ƥ��śa];�WvO�2V�j�7�2iS,��f����Թ8qp�^�FX�6dy��<����ї���w�1��2�'w�Ȧ'7KI�����j�*Rrj؃)��mz���8�3(�!n�e�����0�7R���e<���T.���\�N�΅����`��f2AѶNM�-%��L��;,�H'x$Yh�+̽����� ��bK*�����B��p�j�ag �l��ͬ�J��oڷkr��F��$Óq��d��0Jh�@Q�*c��Y�	80�X�H��N��4V<I�4r����.X�L�8̢%`�T��Ke�v���*f8�&ݒ��aR�A�:$ˇ9i���r��)�[I�ٗz��z���,�ڣ�h�+�����幫'8�C �.VH�--�,IB�Mڬ�b��K��̫��L	�.<�
h��`��d(�lJ��m��Z�p�sr�@Vݍ�^틦�Z��`'7����{�@D�q
{;{2Y�f�%p�ލ�4U��ٯ�5�[���}��$#�HB?�Q�wtwE]]�guu����� # IFH#@�I F��ꬮ���.�����㻻��������㫮;���⫺㫢��;����˻�.��ʻ��讨�����+��������ꎪ�.��ꨮ`��	 #J1F$��%���u��Օwwg]��U\]�wY�Ugu]]Etu�wuwu�]U�]�Vw\U�]�t]�w�wtu��U�]UE���U]m$$�BlIF�`$�����:��.����# ؒi���#H@�wU�u��]�WVwQ��BJ1� l�B		����=�W�v?_�O�W�3����Z�rj�`n-��oj��k�n��wއ]..������Vc�^�Z��M��v�t��Jj9A����eq/��
�Ҙ����7�v��ڙ��s;��ܯ�ä���@sa�hI������u��e�e*�#<��%r�7V��]fu��gY�u����L�ji��2H�˽�b�ݲ[��	�3i��߯��k*&.bh9a@���kVȍ����������ּ6�����̾�(��^�3���[����Sh��έ;�|hܝ0�Q�.ڂT�O\�Gny*�E¸fS�����,2Q���F���7�*C&T �gwoV�2�&H"�����R�pG-EvJ�gkOe�T��-���o�QoJ�`@؈ir���JD��h����'v�qP��1����t���ae�%)��d�
�H����e���P��݃t�U�W@�%u������.��{r�9�����+zh�^��I��2��@���,���&S�w�C�w�wV�az�\�.�x8�٣�K�.܂�x��\�]ڂ��׎�ɟg��`�0p�kF���B�������/�ai��
��/��V��3���yhE �ͺ��t���#�q�/��+qwԔ����JT�ºk�ӎ�w�?u7���,�5t��z�T���YjfT!L�e��4�k~�ɠ��rHaGL,���:�_g-M;A���Ėu��f�8����V��r\Lsv�/��+рP�}�I�I�W��^f�g�M�k�q��WǪ��kWje
͞aMa�Qy�3;��#([|ޫ�o��=7��y��;ͻ�d౏5��X�l{�^񀊹�VA>���`I��K����Z$���@xo�[^��-Pa]N��qҐ�a�%���f�-��k���ѩ)ddtS��<C�zJwS]���R��|�q�H}![ꑬ�{8��y_L�uvM,�F�U�[ovWs����/�<��ؗ;a�:���d�䝏0KR��������Lf���ˈ�U�DZ�{;2��}�ls�U���&��/�!L�2�����l���02dv�wan���b%
ۡ��$�[y!l(׫���ذ&k�U�V���ә�KPB�L���h�y״P�C�R��K�ȱ���-K,3i;\-I)�f��m
���Vr@[�}V�۔��P�8`��]��7���T�wzl�8V\��
̛$$�����
�m���ѣ�pf���ק]�2�j;�u�5��@�b�9#�x�/���R� =��oor���^N�ӼX��1ݝ�<M�+\U�ź��F��f���ܱܢ��eGWםzKi�ten�t��8�D%���u����2�k���.��s
�zT�L$5h��C^��� ��\7�X�].���ǻJ1򫎶l73�M]�O�������2�w�c��9ZD���n"v.v4[��D1hkąEj���Գ9�,�w\���{�d����4���-]=twϳi��B5\�'�Ž�q4Щ)��8��/�Fѹb����:Ҷή��RzkA��;oL�a�4�������q�ӷ[���̚�����V�]S�Ƞ�̥�um�����n�L�כ�H�����v�qܮD匭;�lpζv������f*���2�(EZ����O{E�\����t���@-h.HV���'u�6\��ȹ�%���N���ʌ��1�%�9Ҵ���m@�,�ȭ�[�[�����^Xb!�ƮV>��0f�Au�>���t�#7�}N30�iN��NJ	���]���چ�5R��ML�`�I���yj�E����n^7��փΔ�i,0�:��)���6��i�.t�.��$�n����^��_)��f�OE��7M%p�MJHޗݚ���E.�H��V�MN8��D=��n�]��:�N�x�-�7Jތ��,��1��Ȗ�UŽ�\"��|hw)�7�ޑ��N�C\Ź�Ӛ�W��՛�-��3W����C!9�b˦�2Q��/�jյO�n��,��f2��̇u�KZ%="�,��ҁ���֙iP뷽g�P͎�2�z$�Z���C��hp��o[���)��U˲������7a����Z��*�i�&�6�����yc���l�����u$����L확kA3K��Q��r�<�&u��:fA�ٕx�G]�m��Q����&%Qz�qV���N�Z4@z���%5��,9�S.Ef\d�a)���}%�=��K	UZ���k�;Em�3�Bs�� F�	S.��h%���=�T�7U1�s7h�9�V>9���S,�P�y������eЭ�N���N��T��.�s�7��o3kM&���Gu�������1��Ų��H�!�ȡ��ފ���"���r���E ��y! ��kgoV�ε��]3����]޻���0��wֳ -�`��[���]wݘ���Z_,��oBe��&�r�);��n3j�5c$YZT툫�P�b0�F-�p+i����nm��H��^��rq�VV,NѸjbƆFPYv����-wer��s�l��(��н�WN��ȕj��^9�����b��GXʖru��n�%رtIK�]�+_.��ڊ���'�W�D�sK\�	\�Wq��b^U�e��*�"~��j��G�J�v=v��d�6U6�Ij��;8�2q$���{�Ҥ�3��T���T�E4�q]�]�'{�����1
�0����(�B���:mN�e�&����
܈z�ƛɻ۔�e\�wA���\c?d�����n9�����4Y�%C��T#��hT����*wT7�uifgE�3��9v�����
*�>w�[�`è�FY�fփG/6��W�WXM;W{	��r��+��6ز�(HP�a��ծv�r�[������%�i�y�3"ޥ����=�����I�H�"�M�gop4%���rs��mrݙ�Æ��i��J���>6p��ѱ;0��� �j��ًb�@��9`��;T��T��lU�tГ���7��FҺ|��Lu�C
��N�*���1(˴���3�k���G���u27���6ʮ9�p��

cw�U��V�UA�Cu�m���Dm�����kn�*|�{F�.�J�V^a��GG���+��!O�V"�owV����.Uݛ���mr��\�G��ZGL�Nq���8�3:mn�a�������\Q��Δ�*wB����A�f�X��V,��f.5�{�zVn�?�q�2e�vkF��:� ��K�H�F�����z��C=��f��Y>�s3um��j�EO�m��p�9ȱ�l�7;e��4�U%���,���M���W�L�f��k��[*,jV><���T��x۾�$Vav��Ɏw)]���P���3o��f�
�ѝg]j��CC��e�Huc.�Uj��ٻu���ݚ���r-x�n�!e�H#��ܫ<r����e����.p�gd��w��S���ڮ���/-�r�����wcx�T�ccÚl��\a���j�u��QL��v���Q}�x��hjeL:H�e��́����S�@��w�nz#u�U�
5g�jG&�����Ǧ����4���#��yUfu5��S;6�!�X%1w�JZ��l�0VT��R[Jؚhg�k$�L����({ �u�wj�ڔ�-5;��/wrF�l� �����s�]�; �P�!%�rF���o>y�홷r�:��h$WQ%�{�N�U}MK{�My܀$�u��vn���.Tu5�cY�
z�D��nQזC��y}�1]��i:�Z{3��}��h���;�ȕݵ�@�q�>q��B�J�e-tmE�HÒR�j���a��M�ĕ��ݛ�w��5�+Fa�Sk^���5�ð:J 5X����^�Ж�ȫ�ꍵ�;p�"�j�Yi�u%��	��8o9�k89lw.�fj8��]u��&d�:u��|�������v�E����B*`���M�,�4!Y�k�BL9��:�N[��]����]�aת��W �V�`VΙ��':벷����ޢn��o�z��z�⾰q�����n�f�����kD��O���9�<b��ז�܉��1.¨�53��a��}O\�A�"{��:J�$y����e�m3���c�ć�u����p��9�;R	j�g=���5�tV��֑듴c���LLTj���j�}��B�hJ���{�u�*��}� kK�j�L<\w8j��7f����YR l�/���u8��5׍���/*�ؓf�D-lڽ����B�Vy�Ga�*��Zȝ�oP�4�C�)�Ľ�V\��%s������Z�$��zB�j�_\+V��y�<1]�;lfܵ.ν�̡GU���vG�Pb�V=�k��8��+5c��f�:�ݝ��I���:��g:��q�oNm�.���̽^0�e]�#KOuΘ��A--t�|p3#�7��P�y���Gh�Z���o�x��<��~�q�}���\��i��T�n��G)XI�S7�hzFe�� �):�\�H���-�s*b9�b�ɂQ!n�˷X�������������[��{�2a�����1��R��lYp*1%YUC�3	��l�E�C)�Bb]��D�
��p�k-q��:�h��q�d��|����jf�2#y��^̱,��.�k�4v�P���9ғS�����uL�M��!���w(�RQ7�`Y�C�0�`�r���'(�ln��"�o$)������M��a�S�f��a���K�Ln�2���*^+Ƹ�
n+��l���Ĩ���177�vZ��+
μ�q�D7s���Ju�� ֭��\��y{�v��S���Ǝ�C���Sr����r�YD�{��1S2��COQ�"h��֤����� j�<��Q�۩��t��P���V[�1�̸�X�,�/7R�>��OQ�}��Wnt۽|6��%,�x�5V{3pͺ��̒���\{��.�����ї#�a��r�L�	��D4��7U�Q�����Ni��M�4%Df
6��&ِD��m�y�m;D�ľGi�U��jRu�ۢ_a��\	��m�,��L0]�T��Ͳɸ5�W3y�mr�̵V�ӹ����Q:��8�&T��eݨ2���2oj0ǫ[ꃷ0ɝ�91����0hF,Ӄq�W#-�K�FV��}A��:�kAZ���8��d��HD���b�9���k�neM.�i�7����b[��6m6�eMc��u�ћE�Ӌ�7��ZN�ٖ+Xý�2����Q�Jh���r��]ݒm�{�)������M��nn����̂-�-M%B�W6�'��ZnjU�ڭQ�i�S�����nG�^�j_]��q�6n��
���YԦٝ+s�\n����I4��;X1M��5�C��!�	N�j�i٥H���E�
�e�+��hwpT��ޒ��9lӸ�p�[�`��R�.�ب�v�A��,�r��g;5^�^)(VE<z����礥IG�"��Yx�ʳ�N���47
�C�C��"���N㢟r1kPBٖ�^������}.�;ݮM����"�:�o+6����Vm9KE� ���̻S�^Ж��ֺ���j�i{u'l!a<8P5׍��G���w���b�N�Hp����P���[�/oi2t`튋p�jJP@�L 9]N�0jVؠ{q��m��l(���m�����նѷ[��uf��|${j���O]9<x���i��ѷ����ڵ)T�-��R������s�'�b�tR{��`�]j��]��l]�}[wF�5X41p��c� �{�*��������� 65{ս�N�3��x^��&qu���<�--&�U�*OR��'��=�{b}[��ȗ��J�z�荜Z�����p�9�����W�諲���oP�¯*��
h��ɱψ;}��2�r��m�.H�v��,��u�t�d:(�F�y`�(�d-��C�si����5y�0�p�;w�����A�E��y���l�p+.�s��Y�Y׊h���N�-�3j���o�O��'m�E��z*�[�F��V/gF&�xq�W�>}r�)mu�CN�u�)�Ƴ��f�s�H�ȸ[5�Hq�ק1Ӝ�3S��kD�p';U"���B�k�����P�1�:u[=HQ���2s�M�mc����Dv6�_[�'b(`�x�Z�A�^4^f��u��\�I�"�m�����v'u���-SQ��4�I�q�sgb��,��+��6�ovօeO��Х^
*�6�O��e�K�����[]2��Y�h�`�zڄ�b��)1���!\-��p��8�Iqo#w��j��%Y�v��^�/�\�x�"���|����ٽ�Y�{:�=��];O���멖� +�,��+F� s�풋��w�.71�S!�GXh�I�����ٻ��n[�53a�"�<�/T�.�6XWM���r�Y��ya����җo���;ʦ�l���W��L�u�Y�����&V�Ƭt�kC������hᷫg��åӴA<;�w�@�:{�k亄�wyY4�Bp�Z�U��;����TF�jIjcʮpM#����7uE�ىe�+wmK���V�����I�]/#�@�8���T�+���9�J;9�1;�k�����b��:eW$#7S1N۩9v,��5F�*Ϋ[�Q4�؝Y�D���'y�@�]ݚ͆��pn�i�E��y��]����=
�ne;�����1%< ݶ&*���{�ּ�]M}ǲ��h�yw�	�q�Uݢ��0�^[��6�%��x�=�z�����2�Δa�o\ms9��4{-���N@�U1�1mX%��ݝ�J��i�Z�"�3t�A�j��lF�l�&�
u�f9Ә���>Ͼo��ҹ\���i����%�K�����2rݸ�*긆Km��Z��o;Q�(�/(��j�zez�7Q&�9�wg��Q;�4c�\���9��#�v��ϱ�-���5�L�,�Pm�i7'=q����B�JK�$4�rs�{h�7`{47Ocm�1݁�Vغ� ynN�z�8��gz�h]sk��j��u��v�,wI��6}���ѝ��<	<R:��=g=u��ٱ6��/fw�[��hf��o2�-���:T��cFȎi�k:^_fz-]:N��r�� Nδ9Q���GH�ns�Ş�e"ڷs7�[׷-�;x�[y���|��IO=Z{����1�w��5�I���(�v��_uuX�Gm,��D�nZ@�q��d�w��sv�k��e8&zI�Q<s�n�/I�f2���)��k�K6��N���EGa�=�d��y����y8����|=��Chm�R��q�.�ܙv�l� Ss;��g�ȝ��\�����y6���/5�uӰa8x�a�Fw5��@ݍ�\rPtI��h�=�kHF�Ŭ�\�Vsu��^�a���)c�l/Y՝燮�n��l�Aϖ�=������h�.=.�gn�'\vn�5�N\{a۴��Y������lo`����[nL,x�7#���lZ���h,��D::����z뎚^ɬ�c�ldI�Rٸ���7u]=a1[L�4���=@.�s��	�x8#��e[(ۀ�p3��{�hۍ��f�7��7��.�F��U����: �V���.'(����\f����.*�N۲ت�����C�s������E n�x����/]ϯ k��`�ݛۤ#u҅�N���E�;{��۝y74c�bm��Z���fӮ��tbNG�D1��z�zn�OU�%����$D�nu�v�m�J�ouN[�v-Dmq�b�m��1�7��/6J��2�V��J9��U��sɞ�gMk,�\u���;uJ�g�χv��[�ö�n�m�pݱ�m�s秎A<O���{.[����nhҽT��.��Q�!\�Q��ce�Z�m�{yX�����l�6(���-6i�xugY{������Kiw�<�����*���5,��۝y�nC3�7'	ݣ�[m؎;�s�[�Y �\u��l����lfm^yn���K��	�ܸ��[�k�,hE��ڗ��	�]-�ę�]!� .xC�"���c�[[�1]睷l��+��]�mc��u�{��;��]p�q�i�8�q2nѦ�6�W�Ɂ�;JR�\�n^�Eqv獻E�/FN�d��<nŦ�8�ܷӢ������n�(�Vσ�r�;b���Ur�7=�v����EWg�N�k��Dm��n�4<����}����8�:ޗv='U'lN-]�Z���U����8u�<c\8�ez����Nv�l�c{m��vx��GC:k��9�ru�A�:m�E�����U���v;c���O���9�S����O7<�Z�9�W'-�o!��]y�S��YK���ٶֶN4�8�@�WҐ;��q��nR0C!r�m��ø/[cITg����wU����#�i7�=�g��ć��65�Cʻo���]���Oo&g[p�z�z�Zg��g 6�g˸w���n����]��v�
9�#�*ڹ��%��WX���c�`��] �Kqv��f����W��;�2�N�ml���ln6�E�;��ROZ�˺�j㴴�������]y�xy��D�p��ҽO:�����`���`�O�g9��m�u�q;������I��@���k�kc۶���v�]<s�QB�T㓶�'j1�ƶ���hv���f��RCa5�k��w%=�\G:��4W@�/^�۫� $�l��.�\�vob���/���O9]mN�]�9� �.X��s�a��\o`��TYe�c�:����vɯ/���s��v��%''�ۙ��S(;n�^f��Z��s�a%�zȝYvĻK {nyM�ksZ$��rq���s=�d�W>���q�ѳ�'h��7-#8��m�Ê��.��7J=T��\g�4K��;s�l'�{[ZǍ���b�s�g��bHΣ�[dY���ݴ{=n��׈�
�b��g\<��@��`�Qi�.Pє㣶��8S\�ݸ^����<z�oe1ӷn�^�lo��N�m�=��w���	�=�&�Nz��Pk�W/n,
N�9�Wn^�����{����CGc��1�=���Y�͋;�4�:�)ͮelc����ˇ���62�;XN�3��9�r�1����U��˻m��ٞ-۱�r%�x�-,��fK�E�lql���<Y۝�snBݻgvb��A@�rGe��N���v�rB�KUۏ6�z�9�f7 �Mp��S�N�M.)�c']������.�]�
1m�#��Ce%@�ɋv�ݎۖ�c{]�==���ѐ�x^0�vVAǗ\��lo3�Y޶7��>�k��EW����{��
�z*��6��f:��#V9ѝ�펎�k�X�/v�[p��@&�n۶=�ș��X�<&\��WV;,����Ȼ���W7n�sh!ug�R�v�G����ݑδ.��m����B�/[M�]tv;h����0�:w������۳��n��=[!�wz;`����nʹ��EW[��jjϝ����ϭ�v�A�t�'.$�:�͗mͩ���6�mL���l�*�<[F9�۷m�dj���D6�u�7��(���g��D�q�k/�
6-	�3�O\�q٨,`����'�Z�O3۰t���k�Ӑ�� �PۀƐP,��$��<�\���2�+ʡ>�:���D�;�jv8�|m��m��@nn�;�\[$��n͝Ɖ���L]�89窹9R���v�FF�t`ڃ���m�R�$������v���]��㌺dh�;nw��<���{9��.�u�oC��:z�]������ݭh���n�v�.��Ypl>Z��Β����+	5�MIS�
����P���A"���6��F�x��cc�S�9�s۩��lX�3���T��*)e�N����l���n��A��;)���`Fn�C�RB�����{�q��g��޽�Ǯ'���닳�Vg]J:.X��*4�٣���m���^��>��S���x�]�y�->��oa��x�Gu/2=��ݨT�j�:��z�p���Qz9�رٺ+�v�Ӛ�d�ϳ�ckn��r;��}�أ��n�����4��V;;vU2�R\Xm7jrg�O�ݕ��-u�����糺�nε�=�ָ��k�qNi���������]f���Ӯ�����m֖�ۺ�:�y��[�nm�c8M����b��v�&�]Q��eތVq�l��юp�d�+��9�wV��QλzӍ�[�\6�ݙ�n�.ݷcQ�q��=yx�T���^�<��:坛'fyn�Z�E�]<�<	��Ms =ȜZ"��{yB�lm��9�8u�������������C�c�S�b��a#�#sN�c>l�:���x�����s���h��sss<�6��2�A����ܹ�G�]Pw;�.8�k�:f�g��n�y���G��<n��j�N.j0N�)Dd �EQ4)c RGI���G�1f�n{]�8O<�e�W��{n�l�%�������Q�+e��c]���v�N2�k���]��[4E!�����1ĝ7��ogtݯjݰ6��^���ݻ<헲<�<mk�7V�m�E���d�R��]>��琸ӆ�=�3���nP�ٳ\H���Wv�(xT��qƃ�cv� ^z:+�\coI.�ݚ���6�[�;F���٣e�n$���qs:7b������(�}\;��2[أcs���M��cG&zLn��vܦ�]���/�G������;ֺ�z��uW*NQ�=�wn@@�g�眏cf�m'X�v:'k����i7��l�N�]-�J4Cӂ��O=n��ȒuHpc����^S��naۗr�9�\k��Q����ku���j=X�ԇogpsڭo3��E���tcT9|s������C�g�fPn�F=���68��K��:�.]uV��Vf���mvj��oN����<C�l��ӓ�| �u�'N{�r�7��k��]Zі���Ij�q�t7=]n�x�`�X�=����z,7!�^����[������9�k��Mθj���z�V��j�{\�q�v�yӧ��&�����Pq��˭�̡��O�3��nۜY���Q��L�b�6ۧ��cXR{��.�r���}�
�.�rv��]�I�i�ۙ�ܜ�z�W>��"�d��m�{m�rm)Knfz1�a6�cxż/Q�k%X�
<��D����)q�:�4�;u�]����F� �p����Z����f��jGw:��yn;Vw��E�[b��6�h�U�uX0��a�i:G���x^э���v��i�on�۶�,����M�<�e۝��r�!�ݹ�y=��X}�oonэ���"����v����Wh;n�l�lY�m�d-�\kVx���蓍�6��z$<n�qp���B�Sf�'7M���]��&fb�a���j�b�ا��I0h�/�����[�얹ŏbر�c�w;�7H�����뭺x��${mrY��w]����xK�N}�IH�G\���w���]�\�J<0��鞄t�\����W�8"0֨�w���ƍ�L��I�����z����	:5sy��na�\�{-��l5<OWu�5�!��b��ظlu�m�:u[��7.<�7���(��<��l���GW]�Ey����Ҽ7�n�TևΔ��"�\=@"�1X��p��\�P�zK���}U���"H.�F�iif+,r@6����ͷ(p�oz����:���l�h�H�����vV���l�;j�9m[-�$���y{����dv-��"S�ȗ���[X:[nڳ�d �2�Ye��i���]�݉:{w��ti����$Hش�HqE'8�fl�{�	Ξہ�'(qf֭6��m��"v�A��p����d^����V�n;n��-lֆۧ,��q�ۭe�)�!4[n5�qD���pm�'F�!�۲tnY1gH�r��)�ם�Z�dBQ��ٹ��R�JvkkK,�N�8���P6�����%;n�������Zm���rBm�ڬ3H��I�m�D�3$Y��89G%:mdm�@��l\�Q�l�t�mm7mnnm�GN��Փ�h9����9ծI�;#����cm�|�{����]6���&wg�r� 琞���v����Kv��m�h��M�*V�9�x�oa.ݐ�qʯY�0�#�s�(��pQ��ݜyv�lg%�`�W��v���*n�m�#�����c[wk\v#����:V�m���غ��-��0�,�H������ճ���X]N��D����U�������w�|�����o[fvӺwr�;����g ����/c�\b�c�Ϯv���vƷd�G�K�{^�]�\,Y�q�^<�8�m��lE���'F���Vۭuڶ닪H|�ͣtۚ�v�c�l�0�ې�K�8r�u�2�m�m�i$i�D����5�d�D�C������<�l�u��¶vz8�g���qd.��s������ϔnƝmq�	jϗ��I��ֹ�XZ��lOf�p^���G�}`ܿ&�M�;C�#��ٻnL��;k/&Vw41��pc��b<l�]7Ii��O��Wl5b9튭x{tr�5�L�/6鮻5�ʛ/�-�=�r�Z�p�[�y�s���m��?3��彜�8�8�g-n����ղ��,���u�t8�z�ۓd7>E�c��g�;�#�S;��n-���ܩ煔� �F��3����.�A�lp�����6�t:�W���#�އ���غ7F�#�س�\�>���bz�8]�=�=:�[Z۷k�k���7���c/;;�8N7s�s2���j��6�:�8J�O́��5��5^�n��.�{.�X���͸��1x�`Cչ����r���;u�z歰v��i����ӎ��o�۵f��m�5��$ �m�x�fC�v��<#"󙸧�\t�m�%˩H��LnC��|)�]��tl�m�]ghۃ�U7n�vN��u�۶���xځ{��2NS�B��շ��u�;*q��rnn�u�n�ɘ�s�s����C���<W�]�x���;c{���>#@e�����÷+��;dwl{`7l��������>ʜ�ݷ/=�0v�<�yg�ޒ�����g�qʻgq���ϗ��2��w��סy�3����׼�f6�g�����H�����{�KK�L��ힶׯq�4�=��ɞ�r��r�ܦ�3�P'�)�c��`A8�4���9{e�q�+�Mʩ�64҄��Ch�:z#Qʇ��an���OĒQ�UV� {����͵��R���J�$�U���Ϩ�&V�
��|y�[�Z �w��U���糋`��;5� >�}츀%�m=��m);=�T&� �࿍�IF�k�f� �׽�����w]�t��.z9�'�FwZ�t�y� 5vjLcV�j)��f�����w�ٯ9|��t�����5�e� ���w���Q&��>�M�t�f��7�V6X��t� _�����ۉ+o}-�@:W��I?��$=��GkGo�}��7�ҋ胳x�^���s�Q�F�B۱�C+{N�R�@����w��j'KB+� ��׌�&��]���I�=� =��ڧ��w�uɟ,�w�q �����r�����a��ݒD�Wv�9�_fM%lC��ĸ�PqF�-���=�t��A��
q��k܃�}6W>���4��[����ث�����|�Ƚ�I�{�?�5D����I$�=}M�����{�����a"#Ǉ���Šr{͈I�%�'����:ܢI'�sN�4I�ܞ�����࿍��&�O�Y~���>W����[�����&�=�{3h '��+��.��_W3O�����_Y&1��T�ϑ��w{P��4M�v�Y�4��ѝ�'��i�����*������<lj��r�R��S��M��"ob��^#�\x���1�����-�i뱜Q
������!eP�Us���ً ��}�ml> >R{ܙ���wսs�>�t<�4�M��J���EBЪ� ������|���ū�k� �^���� �{ܸ�`]��u�M�'V"#��"P��xě7ۻ%BI ^��f�$����o��(𖽃k�Da��ʷe�����t$���z(�`S��Sݵ+�<{��J'���C��M
���V��u��s�� �����ۋ{Q�LUFRȲã^���zj��m��>$�'tl*�&�ݍ�D�$�5w�}�`��ݮ�d/�4|���Bk���Q��h4�"�튲`D[�~�\<��d ��j'6HI�I7��@ �]�kM�S��ocqA��-�N�[`�UWkUn����I������"B�]�����"�U�Z���O�щD�$_��d���7��VM��=#��B ��̟�t#�6Ne]��X٧���$��������.�π{�}�����Y���)���6�S�� 1EK+*��'��L�I�[�� 'q�S�Ӝz�s���s�| ^{�>X3���X����h��+�$ٸ}���C'���� �y�Z� �����������˖w��4�L�;WjQ�ˀ�,�}ض�J�R2�k^�g#�PI����F����4�Z�yA�G.I4���,�I�.����WԖ�l���&�{�����Ta��ck]�kk n��!.�T��f%��L[� Vv�L��Dzo<��1�o[܂C&��!A�>D�m�d�B�n�ޱ7oGl�[��U!�(�iR��^\�k�"Z	�^@�;˦��W�����N��>&�ZNI�{��T��v�����b��cU�ڥF�#3��b|M��H�DE�$
��$�?j����"&��2!�}���Z�rL�v�'�]b7�f, Os����/ϖty�h�I�f��d�M����BT�����}�rs�����o(���t��$����	 �+��8�b����� �}��$��NX}*�(3<���$�D��׌��F0[N�`�6
��ְ������`���hW�G�^&L�	��"�ظ�,�s7�Z1!w-t�'"��'�]v���k�
��X��ή���`���څX��^.iha}ĳ.͛� Sf��&��
�uh�y���]�q�]��9-ͱ��jy6��瘺6ر��{nYz@N�}O�Z7Ug�Zv}HăU㩗"v��2�mu��H�z;=���ظ�V��uۈE�.nnOe6�p���һ{]���6�Q���"�<�%�=�1�Gyט�c�c�r�,�� Þ��
��y�c��py�۷m��������b���zIݻk�ۤ,�ˤ����X+T��= 8gj�]����0���m�B�f��|}��P�I&���l�Vj���8�\~K�6$N���=�U���8���y�A���d�ݜ%z��G�$Q$�W�{d�I$��{m��$����=˚��˽I0URWT��5��w������. ��-���Z� M����� O{�09�#r8�RO������{����$�ɱ�@$�~��$� ��J��uO�%�`B����7΄ r��*��|=�Mb�wrl�2�����C��?_s�(�U�m�d&�{�?���:���Ar�{V	]����ϭ��m���x_Glh.<O���sv$V�	T�{���C�T���9���ߐh绗 ��ڭ�4���g���������Ƨ=٘�Q�P�&�vK��7�"~$9^���_����K����@�����o��,�p�}ux��}(��~��,��X�uy�/wveR�";����;�L����w1�lz�G{٬�7�e� ���kۛ�9��o.W�NZ	�ѯw�
��k4�d�U�>��5����� =�f`���츀Y��H���-�fQl���{�D�*��$��V2I�����'�O�.��gn��@���t��K���7�8'���W�w˩�D�彮B�E�~��ȓU-���Mhf��?� �b�l�
����J�<���N�M۷���u��:��;{q����|(�(;-�����!$�]�|H0r�t*��p��@W���ɯ�4I�'{d�K�U�X�T�[����vg�1 �����N��c҄�$�/���A5P�ܷ\��8�c$�kV�'D�$����۝p˾OkS07��+�MX�c�.�{�K ���oa����7��-�ԱA�����{X,�e7�5�n��1���̢OE��`O��D�Y��_N���W��m�͎�ٿ^�:���{� tI9;��Z��@2�@5O��Tr������|I&�, :&����$�W�m�֗<N�����ˀj�RLhAl��7�O��>��$�}�����n�g�Y�gdx�$s��B 4U��n� �k˽�B��~MqѨ��C�U%qV;771��V���wb@���X�F�5������w8wWL�����fh A���7�����3	��߇���oBp���ɼI&f�F��M���)b�U�A���+�����|�{>(E�h�}���% G��@:%�W����8f�<�O���`ϳ(������d�� w}i�I��yYzz���[�n�{ ���}6�>�Qzb�AƝ�y�׼�u_s	��p���;!���@S�r� �I�W���D�a�y�4\��w7^���ʌ	�,F��6S�R���=[XKU�����_w��rdmwh�GY�zv�_>�Y{6o'��vc�	����!>���8���y��0�{��>;�'�,,�ݍ�	�s�O��6ID��4U��� P������Br/_���_8��]Qy�5ڱ��6w�E[m�n�6���ݮz�NI�d����d�hE��Tg���{�{ ��w>� �}��f�[�:��9с	%_�[d����,�ee��X��X8���֡߻���&��J�z� ?��y���J��V׽�v���}��-��t�`�,T*��Os�p@]�u� :��{�V��{�@�g7٦�͗�ˈ�;��֡�2���3�luk6����#x�Q$�{� tH��s�?�2s[����vb�]ҋ��4�`cïy��>߽��w=��	{�O7���`6a^��MM�{��&���R���AwV	Ɔ����^�^^퀐\��R���*�zHNQy;H�6�R��jV�ɴݥ��0&�K��b��b����Π��+�Y�p$z�7��ۗg�i�d7b_sDR�7h�"Ǝ[�z�{]��I��vݹ��8t>z����=������-�ɶ޽�p%�R�b�/��\-{<��grV��X8�\;�r.�Wc�z��!����;m'9-q[;���ku��u�V�Яk��K� �u�M���9;svp{����n����V�d�[�ms�$��U�7Śg�����g]"�Y�z�j��)ì2�����c����>k�0�w� �^�h�I&�{�$$�ۓ���]�m��ǯwW]�&4
��j��Y�w{�|ߍ���9㹾���]�\���w{��O����='�k����^\�Gj�}U�1���Z׽�`	TI�@�ynl��}�D��?C�w. >��w1��{$l���;�i��:�q xk�"I$��� %B�헭����<_� (Y���"<62��Z5+����{��ok`��)�w.\��sf/{s� ��f\ r����LB�훸o�q�J��S3�!"H�;�1�yC���Wb��*���¯]ȽQ�T�����~w��mAƝ�~G��y^|�A��w6��N{�2|�����a�猐	�����^�ҹD��"y�H0�w.�����������Y31�͏�1���kjVP�{8ڀ����vG*"��o.�M��g�;%��g̮�o�V��B����<��O��ԽH�I37�@%0��m���ܖ���>����oڼԓe��Tf#Y��x� p��ӢI-V
]�X��խ��8����������f}��9[㣂�R
����1�����j�Ȃ?�����fb �k���]�]�F���{�o{�M�����YYGs����$�<rh��J� ���l���'��=�|I$�r�����+�x��7������8�M�������
��.S;q}�S�&5��w2ܶ�S�4�����ޯE�.���͌B@þ�L�TL�Xɭ�u�u"�z5��`�1T=ٱqC��D�b�X$���h���o�{T��y����g{٘���r���nڇӆ֨��O�d-'$�� II)Z�3�ˀǯ{Y���>��w	y��2��{0�f�V{dybe���Y�w��n���KN�R�]�(_X��ބf-�Er�����i��͌cWǬoMz/y��׷|b�Z�:�Τ�Y���X���������ܸUÍ�"Wu0�%��0s�+$I�kE4�J�͛g%]����")V�..���2��Nf��Q�Y��*f�v��R!���S52n�2�}F[�PB����hHH�,acuQ*��3C5�����-T/^��jZ5�z��B ��ʻ�MHq���i�VV"��@�M�j�od"[����w4͜�4�;���8!���y�G�Pb1����SO0��:6*�H.2�*���:x��YAcVY�7�W/E.2ȼ&/v���oSOv�F��gcj2u�X���hݎ����p�R�owۖ�Է{�dT�"u����}����/h��9��9]���;:���J��󯯅������Mr�.aN�u�a\�+@O2��N��4�ۺ4�1y��Ӂ�oHJZmc$F�*�
Zj'�V8N��_��g��[��<�D�κ�+��2�����Y��"U��8�gmw�vE���`�$���Ȥ&�B���i����XYi���"��nЧ�2��"]K:�p�c&�Rr��٩���J�6��*�E7s^ũ�E��^�A�#3kV��h���)�x�5XN��`��n_!���ٚ��|�=h��:�iNV�N|鏜��w$S[Xf�.���8�s2��J�Hd��Z�LG�,�Y8��wX4@94F�V�%��0bL�9�\�Ӹ�f��,�I.�6��[SZ�8$�i��ø��m���K[I�����mm��H�l7.�d�6V�l��"��)Yٵ�ܤ�lr9����j��m�.�vn�b�ˇ�N$RS��Tpۻ�kf�!Y��;0m���Gf��\qq �G-��6�H�gi.�֥fۖ�v�۱܉QE�e��蜝����t�H�r9�ݵ���0�S;N	%L�3�Q�P��%̈$�r@(֑��	m��6�ڜr)˶њG ��ٜs9�K�fs����d����m�C�Ȅ8q��9fHJmd)#���FnrRS�s�ֳ��b���I��ݐ͵�E$��()!�3�����=�Y�vbX0�{��j�4���������g��-�� ��\> ��w5� �^��/�g8��F��LXuo�|tpV�H���g=�Ńg�������r\�Ǐ=�x�h�C��i�h��]�g6C���g�m� �0���H�r'>�z�oTh�F��AOlp�j]v��E��������)e
���o����w�ŀI�MO/t��iL�g�_�Ԁ�͸$��}uq�{�^Ey"��6lG;͒N��Q�f��1>i�I?^�@2MQ��t�5D��^��#�����t33w�`/kΩ�}Gv01�����I�f{��B~$��V��|����,�@���k6#w����W�U�uX
��n� ������W\Ⱥ�^��z j�H �5���BI$���%U�˕Ҭpm���b�<�9���
cy���Z������j��'/&ݮ���J�I6��6iN�D�S�_Dq�HAt���;�i�SWd1�`뒈��5��c�D��sN|��W]�F�	����B{V ��Fd�l�I&��̤i�m��翿ߋ�zҜ��b�b+���xg�����M1����=W5(�Th��U\��>�8+]$UL�o��X��sk` ��nb]���Ȼ׃��P��$�$��t�P��Nuv4���n�$��3�`�i��bsO7iI�S&�$�{��I�I9�r�pI��'pt���5�έ��tgqS�t����{��7��H��Ŭ H=�-t���ݷ\�6$v���� �{ݺ~�qM)�i���໼��r���߰�o������u���dE+�v�|'�DxB���8���*��lˀ���� .k����.O[�����e�d���Q&��wb�$E�4��u(S��5�PQ���<��Ь/����1X!I��{�Ո�OI�{�r�Q(\e&oMo��=]�4R��9]�
V4�&�m]�Ʈ�e��vr��ݜk�9w96����NW�n�����	�ݦ��d9v��4�;2�;Y1�cώۯ<�Wg�2�0�Ws#�k�t.N�-�:ѐ����ݎ�A��Z@��l���z�X�Fa]��t��{e�ù��:����90�.qt9y�Ԧ��%�=���\ۏ`��:���<�����sk�ޕ�ml�ʹ��y�%�ѕ|u%�]Bjj�ͱ]�u��.���vh�й���Zv�h�F��﻽��	$g��d�I=��"�Ừ�~��lb��mo�G
8*�r+V�Q�=��H�m(&L�����@'=���I��Bg����D���S�f��o[�%��=���7iGJ��@���>L�h���N�4I'§��i�8��-{�;�m >��}�l���٬@'ѝ�O�A�f��q�u8�w}f�h����3D�����@:$L��������$��d��ʷW�b�X$��tq�d�h���9��7L��`Wk���MF���I$�f{�%C��O*ƫaK|O�a&u�gґL(n��͸�n�n�G�:�;F�ڭ:��'�jD*�U��,�ꪸ8+`���7�Z�� ._{Y��3=�|Om��i�mc��݈D���"��Xl
��4.�e>�I	�lMj�L�3��zF���T`�6fS��De@Y�]�ը.�>�Vn���R{�z;_>ќ䄲�1�wL�E�z�vb�2�S�p'7ԙ$�I=� �AŽ�� ��US�qJ��q���\����Y�{3 �����4H�3Ԃ�d�$�53|��I$�^鿶Jw��ݥ+w}�m��x��핆�v���+b��d� ��  ��WM���I��]\D3���*�a�"�ٮ=�H{���� �~)��$д��$�L�����<6���5���-F��N��W�A!Qc�;Y݋�ɍit�9lv�xi��e�ᝪm~�>��yO��N�߾����@ �5��� �4g���q�����W+8�ג@j���a��W1U\��'��9��&��+�^[�,=S�(���TI�^�! ���cd{pV	8֡ݹ�f�'�:�ڶ�8�Û߻����$�������*�5��[r%mV�L�U"֪vSP�����m(��u�k�ޞ�S�Ъjd�Q|�Q{ӫsg���=k�\{�oZ�'�I����c7����[���
ݮETo�N{���{��2%�h�^��Ѐ~�Mӱ��4I=�_d���MQ�w����}�<�r47iGJ���o��$������f�����:��է�M?.���> 3��İg�|�}��~�����;���|�G-�#*����������14𠾈�k�#�_��69z����}￟��u�n��������$=����4&{�?�M8����5��7ތI��ӱ����3��4�`c�wy����g���W'�k+����MJ��7D�hL��tI���8.�A�;�>#���ڨO���U��K"y[w[�5� \��� ���}��Rܮ���B@zv:d$Ow��`� �YV�'���������k��������ϖ��������'�7;��1��]��r�j!:Ƕ��	��
�O�B�+�r�`V��3E�S):�#Ԧ��{2f,*��o\1>�3xoP�2�5"`�_/���o�>�^ۿ����"�"�6i�~h2I7��lJ����ئ��	'=ݍ�~$�f�L�I�3��C;D*Iڷ�Yo����X;[c���T����vܛ��n��L�P%)~��$)	%��ߟ; ���V�{��﵀ �{�fŻ�vID��*`����?<�̃D����� ���;j�AX��f���>�U�Q��L�I����y�D�I��齌A�k]*h�{[�|���*�4�q��k5����w6���ywջ��P���~$�^�@ ���w�yf����	�,��m�{�l�ʌoޜh�)�iI$�^�%h��~�]�Zc>{�qB:��;��ѿ:%����B�Et�(�}���q�y�Y�P�]VН��I�Gyw9P�D���{�nV-����wX�ρ�f�{�H���c7�3�Th������T���$�툩a�]{E϶Df���W1Y
]�:�_j�#=�ϧ��z���_�w�x{F��t�On��;K�p@�ۃ��[�[X�.�G��v�7f���y@�;i��mӔ+c)&���^]8Kv�ۛ�A4��y����X�)d���s� <gQn��j�Vu����JZùk�8e2VvǷ^��8�4cW6��H�	�ݺ�j����oV����[v*�[}���Mܕ�]��mPa���k,$bGn��"�Q��&��<]�\MvE|�6��;�?y�����Ȫ����fhl��]�T&�$����m�I��c�C&k�ߙ^� d�5wI	U՝�� fX���ctOMu�N�7�u���R Mo�t��D���{�� k+�����\׷�����j�Uh"�c�{]�7�h�w�p@|܇*���z!��n?�$�;��HA�Iw��A�;�%��lP�.��	#C��$�I<���&�?j����$�D}溉]e#U�h��Fn�e�b���3 �Jdn�G�^0Z��&G�G .�J��c��r�4I����@:$Џ��'ܽ���+�p����T�v	��։�ͷ���l�ȍ6q=�{6m���*��i��,O�ަy�)����3���w�i 9�b� -��Q0���>����hn�k�2��DD)�1a���&㰮Z���,�}����,�|?���vr�͹��"��,��nɼ7�ً��E��iPYt�}���K�E·h7���2ϋ���39�WRN�C9i�s"U<Jv۽���xb\�o��b���3 ��X�r�i봻�Zb��V���$�vr�����]c4HϹ6@?DIw�ۺ!Hf�|H���� ��$t���U���&�U���d'+��q�(�4�s�h�I��2I&��{�^�;�u'E�F���<i
���b����M�{��G���J$Ծ�����i�$���t��*����J�����% �j��Zn՗��܍v�ͥx�����4�,�ſ.Ϋ�v�D�<=��$@����`f���`S�����QG��ӷ�v�d������4f:����B�S��1*��U�z���˷��#��h�Fg��}$�X��w����,��¸��0���ꙉ9�f, ׽�ml�uxe�cW���n��ߙF���)�'��ΖSUkmݛݮ�N/)%���UZ����?=�ˎ��,���O�����U���s��
I$+޺Ā ����kf.��Ȅݲ:��|>q��`����� S�j2I5D��wna8""�l������D�޵�>s�����EPǟ#�����)�w�f^iZX��}��x���T �I���u���h��uh��d��pk�m��7j�! 촷��+\w9�5BhTu]s��ꊀ�u��?|/o7�� A��w1���{�0;�e�8ik���8�W�N�L�D���9	�$p����fa��!?sL�.�Y+�ey�^dD�7��D�I�{�� �1Wujs�yw|�Y�q �\L�YVZӈ�W���&�����'6;�~��,���4I�3}с	=���t�팲��`Jw��u���T�wQY>���W9��I$�s{��$�Q{�]Uwڻ���y���!&؇��^f�j�EVab̝e.וbL�o8�4^c�Ͱ�p��$��r'b�j�VF�'[�?x{����O�:��fE��-�	Jd�$o鮓$�\����~��|�8��[�;��h �ݸ�g�=��h�p�n�_hʱ������4
����1n3�5\Z݋Eɶ��N��vQ
��~����aZ�T8�y����@��qk E�4�+�œ*�K��Q�F ��{�0:ixx��(�n�����b�AX�W����\ߪI�M�v7�&�?�� q��=|��߼���N�J�,�c�E�،���;۬�䃢I&���/n�pM�|I$�����c޽�� {����O����u�w=N��(._ >^fk >k��e3=����1���� �����]�zI��Wm*��Y�{3��_w�޸��Z����"s�L���hD�3=�_G��vjȵ`���֞I�W�÷�ԫWY3����KK����7ٙe��tԟe�P�C��a��\+����2��@��2G���陚s�`�𥻎W^�6���Nw�t�#��� �[i�y��h�8��.6�k���w\7���%&�9+��������VχF5�kޮ{���-�|t��r����w�O�_ۡ�EQW�`|T�8e!(���GX���T�ڶ�C��6\�t��S)�PfW����e짮E�M8(���{-�i�V"E��3V%�2��'4�UpT��� ��ea�G(u��]�Ua
P�g�����ǽ�M`�,J�+]F�/n�ɆN��]�t��v��t6���wP�vi�k)��3F�]+Z�Ƌ��4����R��6���lR �m,�!x����
ذ�n�!M9�lhZ
㭵%֧m�t�c��m��A�6&�4�9�)Q�g>�u}��^$`� �RYt�)-9{������z�y��::6�]�諮�(h���x�l��;����T`΃9���R�謚f*+Qj^�ǚ���-A�#b���.�1G�j�s�B�Z;X���.����y�z�#l&�ۇ�������(�5��D7�ؾɆ�]y+�Sx�_���k���j4�v];V+D�y�$hP��Tcq�6�J��h�>3T�'-�q;Ce�&��L�և[[�e��8J�k�4U
�wA���m��\E��q�uY�Z��F�WڶnN�ݨ�v�ɽ��'E�+�dvI 	>������c�m6���;lvVV�m9�Y;�+Jh����.�����������vq���ᶒvml��:RRP8촳A'RZem�v�$�����։���2L�����M93%i����Ӷ��m�.!-�[h�9m�%gM���M�����nVZ��m�X䴶�Vwa�����ڲ�����fYl�iImiEf�I2�DX[�i�$BrP��I����������d[n��ݵ�pZQa��v�Rp!�2n���S���ĂQ�#���@㎂�R���	�,,�6�3m��lI���gn9�gF�+lq+Z�N���+��J۷S�͹���ܥ�l��q#��6������n�(t�ɧe7/:��f��4�n��v��mm���N�������G$A�=���i�wv�=�t����/mXY�Ǝ��j�u�\'n�q������eՎm�=����u�W,�^u�M�\p\s��m���w#��ֱ�7v�c��R�sq�Uw=!���E�G�]����s�QxlV�i�1�M�pa�3���[���=��m�sfu���J�´f�,
�B��$ϓ��h�v�����pX��֫qm�9R���T���v�F�Ra��k��^N1��0�t��[$xxi��}7X���!n�9����ݻEn3E�4���w\lGt�m¯.x�.�;Iq�.�<Q;`�-��/(q��c��`ŵ'l8�l]l�q�iM�8����k;Zx��:-�^2���beݵ�v���vw�<�G/>L��='��k�����nڊG<��O���a+7rI�/1\�Χ��l�l&�n��!��u�����E�����ۭ���=�[�=��_��Y����1��;\,q�ܓf�pvƝ]�!v��^.���ۚ��W����sŗ�FwNیrm!V]�2q�E��s˔.�l�v�!s�k������q�ۮ.�1ڠz����kjŠ�zFU3�v͓�c��ݜp=v�u�c[n�ؤ+ݏ[F]�ˎ͖ٸغ�wkLv2N=���1��YM"-э&�$򫰹��=��l��NHvg&d���6�7�X��Z���;�m��=b<�랇��wnQm9Ț�)��[s�����j��ol�6�M���=7jᵒ6�3�"�P�u�wm�����{�3������[n����v�z,�M�qۍԘ�Xx��f��ظ����k�m�%�l��nC�����]���k=qW<a��udOuی��[�,��r+����3mo�.�묎髝�q��Ho8�7mSЦ�5a;XVqB��b��;V��*\*�m7�f�����%:�O���$��Cu�Z	%�����gn3�Z�u��7�9[���c�س��kr�;��ł�ь)�����/k>�q��ġ�W�E��l����Ѳn!��ۮ�yL�_m�Ni՘�eM�ځT�Y��@�vֺ{U
;�
�Y�Ol��Ќ�mR�K*e*A0P�����xܺ��bzol��˱��HtQ�:�a܌�6�wH��mr<I��6��:+��G�f��;���۶Liթ)w]�u��;��~��웶B�[�m���� >@�{�f��=���k�<�l	k� V��'���?[SjWA�C�����y�U�l����C��0	$no�I&g��V� �9�n�ɣ����]��b����ོ�b����s{�'5W=n������쎉 ��y�D��?}�oka�tY��X�ib2`=g=�����3�@��M)��̒I&���$$�h���5��H��5A�I��ѧ�$�Jb�֘��Y��{�`���;�X������Q&�,m�I�$L��>�@��`���{m�X��yRψ��r$W[s�-z;�����b�M5���+�r����Ξ�tv�AJ�x[�}�����uʄ�I��'D����=�,�z��|��}�f����鍨���N�0��i0/'{K����8��Fo�J�*�
�%��PPiV��©ds讧"5�zˍ�R���`�9�ھ�u+�
2Yhf̍ˌ��*�,�&{��Bt�n꟤��w�wy�H�R}���.#�u.������z[��D�3��ڵPePǉ�o��� m�sص��Iu8�/z)A$��	���0!&���=s9��1J�*�O5��sy�^�W����o7� ��=3�]��T�Gg]�$�m�� 0��c�A+�2`h�{.
{��`�g�;���(	N�����6|Y��Ń s��koO�r��b�kY �����v��� �D�.��f1X�c�\a�.�9{(��h^��O�V)�mi�׾;����� ���q����sMǤW�k���-�d|�&���lbw;3ot쓃����*��[�=��f��U�ԙ��6� ����π=��X� �ֳk�]�s���w�Q7h�Enc|=��p$���N� �L���b����4��<"�/ {,�[�.{o&c�#�����l���H�ץ��n��G�����i�k�kbS��a|����꧛������zf����k.����j�ʠ�*zl�kռޣ��0����$�B���$}��.�S�Gj6 �<�PVt�|�pMi�gu�� ;{���9�vr��؀�׹3����M� ��fg�2�Ҿ����}�.	�P�dIBص�y_^ڳ�7yu�b�q<Au���"�����������#s��F�a��+�6���b�����nI�<���v>�1]F_����5D�7�f�n�=�Чŗ�#�=��Бɩ�/I>ٵ�� �_��d�$��o��?VlՇ,	[��Z��z�vVB��-���� ���{
/�\��D���v�TI7�u� c�,nlY"IE	B3w��K�^ ���\^�Mh�[��$��D�������r�8�)�t����.��n��N�*5�6^wNm �xPҽz�b�A �����c�������E�Zw�HO�đ�swV '���mo�UT�k���lm�s<��B��A�5x�&H�7�H@��L�o�|N�_ӹ3nh���h�T��G��#�3NB�5� ���ٷl,���%Ͻ:�CtN����{y�` �מ�ml$�����@^l�(`<��n���2M ���o{[���8�u������d����p+Z����ֶ�5D���ލ�OČ>~��k�[��kێ���l�Ov�F�e���������
|��4I&m�׏�%>$�&����ꅀ����ķ�'D�ڈU3�s�p��1 '%Q =[�T&�4I9����_��3GO ���g�=$�}$��[<Xta�en��=��4I���ܛ+|�_o��%���e~^}$���?~}�I��@Vu�o� �\��պ���&�M�^5�a�k�u�ӮR�TM�XfV���5�p\�{o3>b�ggrr�r���l���n�����I|�اߣ�Vϛ ����R��;�����cn�Ӻ�ئ�6t{n��Ip�B�7;�7��vn���3sۭ��x��̭]F�8�;�EE��dܯ�t��j���c���'`7axwgl=g����e�ۧ���N�7;y�s�n��B��;]v����<Y{m�]	�����sF\v�m�Wd���q�]b�y�F+��m��7a�$tvݳKVv�z��u���\�e�ظ{M<g��[{I�XGٙ�nX��n߿O�A������#��s{[m�g�k�@|��?��ޮ��9��k�}��� �{;s�>�LR���'SǈY��1a4O'Y���]�#���isڄ�I&����o�tH'7�ʖ�{\��\��mX�D��FF޵��X mz��ϰ	�i��.�΍s���߁��3�0`מ�`l���h�����Fzo�k�P�OĎ�x� ��$��l�K۳ۖ�]�82I-y�d�&��h�[Q
�`��{1`�N{}ͨp�s�s�V%*�h���� �\����3����nn��}yH4bT �'m�����L�&l�q�ݦ
�a�ms��t�k�v���:�ޞmD�t�q��s�� ��ɲ~$�'������Z��٫X��V@'��٬@��?[[��A���f7�J&�%p�Wsp:�;ĳ$����nl�H�{i�˭�y�r�ۓ�f�g�49m����U݌2��Q�{�����ӽ2������рE�S�� B>�ߪ�W$���ۦ�Ik��1�>&)��/��/Y�;ُ�M]�]]CtN�����i���y�� X�������V�|���@�r� ~�l��yf�6�u�+��ɀ�7���=�egy�~&��O�OĒM�{d���E.�4;�aO����n�n��樜H�`Q�ρ��~���	�I!{�O��n�yvs�>^o5�=��{[`k������cWo�t�����
QGK���;u�S���l�s�`;�bۅ�6�\�]Um}�����h�[Q
����3 �s��o`�E{�0q�������dI�H����P�[а(�0�tm�$o������]kهp��r�D�I��kr�4I%{�6A���+Ɇlwk*���{���KkJ�Ra��g���> ގ�?j��.vIMVs���z��c{�N��ћ�YٚeF����9Cp�-lC^���T��&F�'���J���˾L���x@��s����I$�ﹽ�m��wwO�s�b����95(��9經�����?Q37u� ƹ��� 9����v/g7�����w���5a�m>������{Zf�$�w�t����f�Ww|I�=�  |�ws��\��q��I������Խk[���EvںOG"2��D�ٱǠ�k����Y,O[�KZ��IDǭ�|�(@4H^��3�$�㾏=$�*iy�����| k��ϰ���q�K-��U�k��n�$�s.ߐ��ɣ�����{Y��J�3�I���]Z�6�I���u�(�u�~ȁ�� _�$�Zp��D�}��U���9̫W!$$��y��k�g�ou~$���=���?{~����P�!�f{�R����k:n�	K�4H{#��h���ti�D�F{ݯ6��k��V�޻+����
5|�ԩ�,�\T�=����A�W�7'�6��c��pK��m�V�����2*�i���ff�n1EW�����?��?\XsJ~s��ǂ���%�����ml}��ګ��e�F���� \�wZĀ@��7��o&p��������ƛ��*�M�+U���Nn�a�z��V����҃���pÚs����������"9=�<�w5�����`���vGD��}�żI��{��#!#q�*�7c4U�MLO|S7�t�5? �1_�۽�$�c�r���[�1@t��X&� �K$D�I	�B�no]��e�$�N+�ΫXA���]��O����/�`���y0o/���u����'����ʲA��2�LT�Ll��������I�AD)���-s����Sat]�.����d�q�ǵgћ�B�s�@��U�ă��i�yRQ����[�hQ�Nт�0�u9z��m�
{~Ư�<n��3��g+Bʛ�)Ge(��b#f�C�������]߈��zo��%�c���H�27�PBH86��V�����ep��u�;��n� A��	�]1��������a�=v=)�� J�۬������n������og=���<k�M<E��ݘ^x��ƃ��t��n�6mg�o>0p�vŽ���/fN��d����nt��ϴݓf�<��顧k�]�u�Vzɭ�v�Q@^Ӻ�����[�==7\�mۚ���ݚe9ڸG[QTUy��9�/��D����1�{� 
�k�+�E�?x�i	jU�|!�ʱ�V�IH�% ��vEֺ�9���XN�!6��례�@�{��s�(��Z�C���;1�̞��BFL��:�z�w���W���2��z&�I�ۗ`�J�j�H��.$?D��0�ߗf������&s�$�
�j�A�s��:VLHI^�P�$ח�����/�d��&�*<�_zs�N�Ɯ�KF�w���$�Sv��	�s��1Ǘ>�	�'y�("O��z��2�+��n���i�/h��-��=0Oq�)7��ϿZ�҂�31�T�|=dB}hQ#y�]�y^��r�	؛Ǉ-]߬J�@�Bt�	B"���s.� �M�����u�.��7o���8�g�;��v8%��`��՟��ܱq��>u��.m6�lVD��r�=�m�ؽ��-�� Hy��z�3���(��}��Y}�!����^��+c$�Q��JA�R��D����RO^_m� ���	^�3ى6�Z��ȥz���[�����pO��"�Т	�w�d�A������*k��#I�-P'^Aq,�	$�D�ano]�A&쬩�ܸN gM����,TU'��  }�ڏ�����>��g�R:n)OW;\�8�����ŕ�)&^n:�渿{���}�ں �!��;:���	;�*��ɷۺp��A�V�H����}��)I���H�3v�\�Y6����}��{��n
$�E����$��ܻ�0��[�3M�.'�?J�2�~*kӹ��m�w���e�s���6j�ҽ�#/P7��C�Sa�ɤT Z��坓��9º�Ȓ���O�rMd"���%����%����h��'�m�V���S����X������}ʖ�:v�xf�W8檊����~�SHшnm��P�.�
f�<voS��hJX�W76�5Vq짛�,�V��XR�5���5���J�� N�K.P9)�k|dS�mb@l�N�,�ݒ搁LƼ�L,h-�x2od�鼋��[���^������d����`k6f��|/2�p��d9��-�S�k+��"���*��cB�;��ޜ���EʰU���1TVV�6��jj��W�e�x�����"��� /��KIgQ�/8u@��epW}��9A�A	`D���x����ަ����[
�I��"CV�o+Ε�̃;`Z�h��E3��kke�Të�)������s<�&�{���qN�}�}o��zo��K��z�����C1�av:�x�ۥ-uX���Hh9	�I˽��A�K��$�wE�����.Q�"���͜N���*1�%��{G���Y;q����ז�oCkv�.
�5�P����Z�V�i�ưn�J�z8�U��׈�ݴ���dRݘ���ש'J���Qh-"���r
�':6�I�N f�b�Y����,�4�n(��Eq/b�F����]s�����.�G2�ƹ}����f�~�J
�/C42����r�HW"�emc�Fu��ۙ����^ָz�7�/�=���oT�OVbJr�
����ĂhNB_b�쬌�7"��	��I�.8\♥H�8D�
Vh����i�'-�-��r�p��G��)�N)9����	�rbQ3�B@�kp�Yb�Mӱ�8�H�V�����Gs�,t���-$�ԑB�B↵iE;��r�r�ӛv��RK-˄�D'eȊm�72�8������q8����9�Z�����%9�d����	ΉR�٬�3N㝵�X�f�N���P�t8�h��[HEmƃkD�Qm�8E��(�@pD�&5��3(�N��2�.�G Nm�V�`8:mֹ����6��B�n䳲���$;L��R3�)	�u9$.����m,�6�'f���e�6ƛ~I �����6�w���ld�w.����(%R	H5d]k��*�ӄ�W�VH"1�U�I\�\t��j��;��ϛ~��+�!�J4����14����3��;�W~��޼��6�� Q���{^/��q�u��}5�*C�V�Ns�gtO競J�z�u�S�=k����v.�jt�4�'�ƠD)R��/����o��	+����@q��˰�݂I�}�.�v� ����@+��y�����o#Q��(�}_���V-�x��x׳y��|�Ij�J�W#��}wń���B�$�\��o�m1���n�z��+T������B� E[�x�}�\D�[V	 �g]��$��}g|�����
�v3��S}Ó���TW��'�}�nzw���%�k_]g>�o5T�H)�j�8�J\E��{{E�G.�ݚ��Ϧ���y6�u�]�?��%	JBA)���:A>/�b��z�P�Y�%�Yv	� ��B�����{��2	�O��) �u��,7k	�G�z� v�7��$v{g�r�������0��H�u���D�I���Xۙ)x��yb��F�|*��*��w	J�T!v�7��'���%�Y��vA .�@���}v	��B[9�
�x�&�?!B�$�ʳC>���
������H��'Y��b��嶅��}v	�f�R$�AD"b���r��s�25��r�z�������Ίn���,�tDԹ
jA�"b!�Z�2�	1�rş(�6�P�ww=��ɿ��wy�UG���+J^�RP��E������X�fY��2o4��]��D�<�/.TQx:֕�1f��8�&������b�����͗Ϲ7�-�ݷ&8�ۊv헉�<;hn�;`�/p5랹�X8�u��\v�=���9���#��Mr�Eā��d㋹8[��y�����wny�rF-m(i���v]x���ىC�����xv���h8�#���2'�Лm���{�{=�O&���`z�s��ώ�F;l	��kk%[��zKK����dٜ[�G7�8zZ%���=���sGb����t��]�=�`~����($�)	H7��B�u@��}VIG=˳��dNm��j��I�w_]��k�W �E(�׳��>Od~O�[V%��1�� �ۡ��N�n����CG3c'TH�P��.��o]�D>ܰ,��mlU�E�|��$��}vi���wx���� �T�M{��������@P[9�@U �tt�y�1S�l��e����ZP$�ADFb�O,vA�����1�cj��hqu� � ފ�/��|(=>�3�Dq\������8��^mն��ۢE�\]\Vv�;�b��P�+��mv�8�O!@+�����}�ݒ>1ϲ���<�\lZ:��[�˲@$}�V9{����% ݑuڪ�AQ^��S��|s0���A�Rm>�%�cbԻ�{y�朝��g�_pG3�C��E�i�-�b�����\���z�w�۫�?��� ʵ�C�I�?�˰O�3�4(�o)J��sQ8꯷�ߋ^� �qѣO^�sX���4��pb���H$�>�D�5@�|pdˉ
 ��؞�ף:���H�f�m��
 ^K�(z.g��øɛ�3W�׉�����>Ʊvg8j�*�F���;6��AvG��.��I�\����]wd�瑁�nn��3F��P�:^�\�bLi����$zZ�ջ+j�(J�{k�V��h�����sCU�D����i�k'���8� *}�ϱ6�}���ɾȺM!@-eMir�˰O�1�Sg���g��P�{�u� �OqULΨ0�Ϲ^	A%!HJA��
�h
���}�/����Ӈ�O�J���O���}Zz����&.�޿*L��&U�G�����M*�\ԕv`rI��5.{5_8���J��w��{���ܳ�`-W*����^7��V�28�ѧ�gy��k��b|E���;�n�$繊�1�Qe��{���TNa��.dʘH�e���7Ę}�`[��<i�jܪe�A=�]vH$�=˾��6k��.����ݷ���\�vF���ݎ�k��v�.vڸ��7d� H�|Yί!��T�k������έ���c�����M
��ا`�֪�<��;4s	@FR0`�&��宝.�S�x��ӂ���@�����sܱ`�eAa��Uё*yg��jC��(�l��Ofk6�=����sxPw�m�9���c��#�G�J	)
BR߈W�D�Q�2��J�$|�`|(�� Uf��Ld<�=)�-�9�E�Ζ���I'���C]�n٫ߎų�n��70VT{s�7�kD�W�i
�ڪ�WѮ�X_����Zo���&�J�KH�F�׳�3k��P��Mh+�L�Yl�-���	;w,X$rv��d�=��vZ��ɡ�zA2%������q㔺�2�����q�{5���.��Sl��vdʘAe
�'sz��A�ەd�9;Tm
}=����U��I���[n��l�s*��ڜT�&���l5���G��A'�۹v�;U�J�v�����f�ǚ9��#)0
�n��-uLP*g4��>����������9�o>��Oיt�J�M!@-0��s,�)u�*`����e� �'j��#��Yn*gp&Kz��őȣ�%��!)셸�!��U�'�rS(In]��@=�j�I#y�]���2�A5��0���RuvT�v�*��*�v�-�
�7	�Sj��u�"e����vu��Q}���z�����	 2�V��_2=|k_���M\n�<��ˑٛ��cXX��g�GY�C۶M���v)�yV�<��:z:�P�f�WEw\a�{N��:�3	-���G$c6����Ft��ӷn,n�� Zۄw�˵���$���ü�zNїj���6Û� )��v:BѮ���`�;�v��ݞ�0M�y�F�%�)D[����k���͹��M���Cj�����s�V��]=�&)��v�h+����g�����}d�D�H����ӽwg���uu�$w<��:�ld��˝��7B��j�>��L��*aI�.:��A>8��U�ܡ{ض�FuZ�}���	(��8�#7Vg���:��@�$�MT+�ez�=��V	'���Zz�#ve��|O�uj�'y�X���PID�8���BG\�Q��A\�ݷ�`H9�\����G�6��'aB�BD r�/yH� >��L2֖,�t���Ux�ٷ�d�|c�����*$�;�~�&���t��7��^���o=l�:��:g9�ˡ�E��R�����-r��؞���ڨ�_U�I�z��*3(�,���o��wX�KeUjX�$"��z��t��B��]c޲��ɫMӖN�)$D����5�\�g4A�s8l)M��-m�;�ww����1���k�3��%ʵx[�8�ӵ}��!l��~)��{�ڱ�۞�7e��w�D%�+-�:�J�)L�Q[�[�A�]��;0����w� $�ͫ%��s�Ř��� ��sM{\�!��0�'�����N�Ă@0�:�H$�N���ѕ]-��;�o��QEJ�`&�O,��Fm]Qce�F"4�q�}�$=�t�1�΅�O:�+���^�|��޼�n��YQ;c�H+���3���z9�W��u��G���b�*����u
�hۄ�Y�~�c_:	<��[�f�Aq��U�߁ ���wȣ�%#*�̺	�+:j@6a�:X>>�U�P3��j���ȫ��-m�Otk�p��IS��QQ�^k���^沭'L�Y�k�����g��EaV]f_7N�X�1UgL�:���^��S�����з׫���?b~���V�����Vt
Ś�[��k� ���y6���ڴ��ժ��Ɣ�S%"	�*��o]�Wf�{o,��_s�A$��Dns���[-��|�{���ط��6A+���>�l��0�B����Ҧ�7�<� >����ais�W�կ��3�>��?�?:Z�2bθ��;�]f�/.�;�S�'�	���9�)1h���EJ�TL?�]N�|G:j�� 
���bX���u�B7(%���
��<�\zj�a'0�P��R7@�s��A���� �NmZ�Og>��}�:	���,���@���@�"/ڭ�D|��ĒxSމ��"�5)Z� sj�x�Og>��D�0����k�Z�7ʪ�n �&r�A#���$���2���ǃm9�Ng:��~�|�5gu�hH�����ߦy�]ݓ1��T���5�m:����U�,@`��u���WJYͥ�� =��4+eI*eB�L�O�o�~�!����o(�.�D���@�s5����w��NC���s|��x[>�;�RY�tP�v@w��Ía��P8]v�5��n����~�����N}9̾m?{��4�=�����]�F�K����5D����]�o���f�A#���-l	�6���R.�F��c@ �k����=u�w3=�F���}�V���i
�h�*k^�fX�H1�]�$��w[��j�<�x��}vA1�]��J��%)�@�".���Z'���&�-b�zwz���ۮ��O�uZ�5`�i�B�2�����d �Y�,]���"��k��O&�X����[�`�#7]��#�Z�u]��'
�~���s`���U��y҉�V��IpZRT]�x�fe *e^����&�(�1u5��U�@���8��\�b�r;�yja�	�]d	F�*��"�:�E�7�̀��5k�Pޕ��H*�Ȳ�m�㩙L�l�dfk��fc{�F�")[�o�u�3g�7�d��7���Gw�P��Ԅ>��w^�:�]�sAE�@n�5,Rlv�_`��1�n3���y�,v�:�esy%�J& bnHwv�q�ҕv֣�6(VCZ�Ӕ�fӡ��ё�Cp�c���}[�P�7�'J����:�o�b�bmf�D.�t{;��!�kJڣx�ޡ��:8�k�史����ѝ}�Q�(Յ��ga8A"Q8��2�Q�>�n,��.[f�K��K��w%rJ��fч��:B���{��PRe@r�i�9����6�ki�L�+r"4e��l]:�ՙٰ�[1��n�9x+_Gp����Q��W��4�ʱZ��yS�w�S�7�k�G�5	*܃��ٝے�k�5�+TSҠ�mC]�-s�ݓE��WGF�`2��E������_5l��ɞi=��W�ݞq�<��s,M9�!�Qr	A�ܒ,j�n��I$hibN�
�q��{Y��&r\%u��b���OL��g,%c]��]�wm�͒g�_F�٣���+ߤ����KS�(�ٞc�g-<J�,S<�'Mh�-/�Ջ�C�Y��p�0�^���R�#2V{oz�p�҆�����Ѽ����Ĳ�ڹnA6I��NN��^�> �	$��!-��pHNY���Rr(2�r� tP:r�RK��-k"JN&ٝ�BH�8f�)$�q���JI[nNA���
GBۭH9�$���I�6�㐃��s�K;��:;k�% #�G8mj#�DR�.;3��t���ؓ�9ÔN.̈"�6�!9�as�q3��s�����'f�C�N�8�\pt
	Έ���dp�:9�6�k�8��,m���@B+#!8� �Q�	�H��$��9$�G�M�r��$D�rpP�8wkr��p0��Y��̓�8��?�Yusq�a��n�Ϋ���Ll�����v���8D�u��98���dl�sx�X�U�΢o;y�g����lu��W�m[�6]�iM���[vN�=�Ko<�ڶ�m�Ϸp�n^�L��0�[y5W�n�7qպ���5��v�}�44v��Eq��ۣk�\���÷�ܰv�f���7	�t'&]�ɸ��k%k(˲�gc>7ZH��s����]�덞��9�H�������2vǒL����v��6+vOn���6Oq���5����lQ$�6G��V|۾�|r�����6;�Xn�!�/Iu3��׋���p�aM�6:�<��|��fg]!أ$�"O�8�M�\��;�,�v]λy1Y�^��<W`�X9z;Ɲ�g��2�+ۧ�]�P^_]u�k\m5]Kq�a�6�F�2d0��k/]l�"�틧����[u�a�G\�-׶������lZ��v�t�9��s�qs��cka��ړrvڹ��*���nM��qn�w��� ;��O*)�S��Vx�١n's���.ےsϠ�.az��|t�������ps�S�7Ci��9�C��m���c�hjՎ�ۇ�OqȆ�7kl;�m=ӻ�[`3��Ƭt�Kn����=��=w]��g��Zح��;UG�\��%#�7��;P�OG�b�N.mz�ی]��T$�v\�<�Z�=�|lۆ�C�g�ۜr�,����4��`1h�nc��=�4�U����\i�y������g�Y����nN1��OP[s���;P�歜����;p�������v��p�㞷);9K��
nƺ�S�d7Z�.��Jn.pV�O��5�q������2�������Ok�nn�Zέ��r��u�h5+��yϝ�	����ؾk�+���D����lv�%�Y<��T�v�z�x�uH�Z���E^ܦ�)�sy��oP��;�����8����CƬ��Eͺ��D����:v�a���.�P]��5b�&�H�T3���/�=-�jR�UM0�����\�\mpN9��붣cr��7m��s�if�����,rn҄P���[��ۜǘ�U=:vu�3��(룙�r�KK�l�a��<N�79�����WPLm��z;s�&v-r�b��kasq�|tq����Kn��۠$�u���Iò;j@�0>M׆��ⲕ�zU�uͥ�]p�y�F�.m����k�r����k�a#��8gf�Dwz�s��5��v.JI��g�]w��}�0�S*%�	�}b�I���Y4�<Cn�]�3��n�����G�ڛ��A$8	����-�
O;WÛ�J���j| �}��� �����>����W�k[�w��zw@I$����b����ugٵt+ݵ��qҥ[$���t=�b��"��Ne(R�r���Ӭ^�ݝ�@K���X������ǧzv_��ڼ ���R�f�3.��*D]��@�����8�wumTG���vI ��T#s���Vַ76z7�r	��:T:Q�Z��������g�Î{\7�D,q�!A�BЙ�~GEP�$eA�|,��	�}w�h�,�48L�����s�@
�x���Q� aJHǥ���
��ӻ�d<�eT[�b��[�r\��8K�i�
���-S�T;����zlA�1�)&�V\3>y���C���-��l��Ǫ�� 5|�;��6�ϹSs�۱�Ĕ���DָWA���� UB��UH=�{W�H#4`���t�L�`�v�����d����$�R`@Rn������13R �<�
 �Gf�X���kr;�7����FC�3B�R�"��f]��A�z�Ԅ���u� ���$��� ���Œs�b�m�w����{���TrWJ:��I-uGk���^4�}Vޭ�����dr�\��R�y��ޔ����D_��.��_U�H1�]�*b�-�s���v (
��|�2�QF���7`aP^}������=��V���
�Ϫ�$��ؿn�I�6�e�;w��;��t���zP����I ��u`�do�{0��,�g�z�,�㺾2�2������V��U1t�#��v2�a)�����\޽ɋ��Dcsa��5�Y:	�y\�a��B�χ�<�M|	'��������l��D�^#��[�'��;,�K�ʲA>��߬�v��^#�ɕվ&���$�!�v.�W�HŷUuQ5���⣴��o����a���0y��&��g���8�:�ӲZ����T�mW%��l�\�i]k=q�\i�ja��1����A��s�˰	'�9�ݒ|I�v������:q�(
���c�X��T�J�~"�Z�lN���ZB���\ ��� P�k�������l�o�(E@+�33A@�^������*�p�$5�[��L7�B� �;T��q� aJHǥ
�]�twt"�(�c�zI���|O��j�$�}��J�}5t�aFKڌ��S�lJ�C,;��S�2Ҧ��)�D�h�l{�V���y��E�l�=�ַk�atD�n	�J���n�ߤ���W�z�=j�{w���5�]a1
��_!�7��LN���R�LM�T�$��hP'���vo{���Wc���V�3)BA$#(Ȕ&�n����4۔y^�oqrz7nm�vո�P[�������M���-u;�>�������N���+���n�2�~3��퍡���J�E�yv	|��]¥��)��|H9�C���:`�<gW�
�6�t��`&q0�(�E�\��I��]�,����#/N��� �yJ���&""�Bw�$��F�׳�҇9���^/�gSl��R�1�W{v��w�w����V�`$ܵD�`�@��%���v>$�ر4k 5}�H95j� �޻$��ݻ��[qI}}e�'Ĝ���}%��8F����U�R�z�,�c�T�ET7v�*�w�1JhKY���"��L�^9R6H�qЭ�5�}����2,D-j��C9���-��Z�@���q;�m�'`x�m��{t�8�;����%�십��� ��wl�q���W�i��[lJ���/��s	��y�z�㭛Z6��{rK[�h3�Ɏ{�ź�k\��)���1��sc�1�7gvN���u��gv�sAn�y,m�����$(��]�9�i�˂��{Q��񚛵n����q��-g����'PkPlo<��tX���܃ú=7f��@=cj���vA�(��?~��
�*4��5�f���m>�\�6�j;�n��UNꞠ��Y�	���]�[��|�)P��
M���b�8����\��B����D�Gs��'Ę�ݡg��h���%\�* ��H�"�L�"��̻�>���	s���Vu���Āsi�D����Ei�
a@P%H����"F�vA�OU�B�>1϶�B甽��g���﹬M��Z�/Đ�5ݛV|��z��ʃ"���z��|^���	$�om� ��ڠJv�wdV܋�_ny�lvy��ۢ޶.�3�����\�/i�ޫ��:nvD�-���\���aPYedj�w����x���vH>+��$Ff����z�&-n�{��ޅz$E҂J�3�+�y/j��j8Я,��ݬ�������7�:˶:n�o9<���e:�O_���W�qY��n�1ݴA��1�3�����>���}�j���	��vH$���� ښ(�6%w]�~���>R��BD&��s�d�B�x� f�F��ey:B��>P (g{��$��ڠH��H�"�I�$P}w�gqM��'��<�0A���\���پ����C�F��f>Ƶ�mP�v)���P���t>/؍��@�7C���Q>�]�d�r����`b@�=#�˞�	[�������v��w;��8:6�c{�����/D��G{��B\��_.�r�({]�)ӣ���)n�K^�3��,��}Vb�߽�۱Y���r���
Yʉ� ^�ۿ�����e���5,0D"��쮵���]ɁT(��GO2�
�{."����$NDE�����6��<ڽ��%,�=�7�<���J�-;,I��;xv��;��*V�f��Y�<��wF}��zn���I �ܫ�_��5�{g�R���!I�3����V@2IO��}����I'��(x�'(�&mRrDR2��(�fI��/,Y'��ؼ�y�.�}�.��V�H�]�d�zy������	��wW�mc/��T�F�D��uz.��;W:`C����2�
7��R�ky'AUab�������wU�H=<��ѱ�M�	�=���$�.�8B�0�2`�"(��������.E�2�� �F���$��}b�9S5�
����:��"��ϐ�������`���RnjV@��VA���vH��Ϯ�b���&��X@�^e�r�j��`�O�I�<��Ă|
����A#h�Y�4G�V�����k��������٨�x�qB�3�7���#$����iΫ�gus9\��Ybkі��!�u1�⋛�G�x{~&�����]����)I�fIRlFM�ŒA
s��n�P"7ng�ݜO�]�$��=�`�Ă�jI��פ��L�部-h�R��D��z�k��q=Y���u!�G%"eNU}��=\��fI�3.ϣy��r�@����!�j�Y����U3��!�M��s���ݩ̾!�k.���D>}v ��Ux�\8�]$;�*1���B�(I��""+Ɵk�Y�&�j&pӋ;K���'�9���+���f�!�%&|�Ugu%lNt�y�D���vŒA �Z�������"|I��릢x0B�
	+��k	/��X8�z���¨�!7�vI �MQ$���cI�+�mY+��l����"�:�$���զ0�N��j6w:V��gf���iL�=7�͇z��c19&kn��q�+TE��U}����"d8 �=����p�F��f�m��a8R�/�����n��#@���2�2�W��*i�������B�A�=�\��&낓��뭪������xm�\��;;�z�qp�D����lO\V�f���vǞ�׆��bP�v��v��9�*q�qk&�[t��n{V�8����ے�׶����?;���t8�	�fM���$|>]��Ui�j��Js�ݚ��zʻu��c�N5ǃ8�	I��c�J
SJ��d���!gUW��v݃#���Y��-7`X>$��U�x���""IF&Ife�&^�ޚȃ����X>$��U�|M���������Z�)眦>��O�h`����շB�[�D�w�V	$��"�s��8���o�$
�J�>�}}�d�1
(ȓ2h�W��ӕ��qɣ�P
���R �}�~ ���y�����!�wb
؊���R�ϐ��ޱd�o���ִ�_�5l�m�*$���~";�lY��^�)����շ�mC�,-�`1�5�2�����g��8̸2N�%�&�<_??���	�S�!A%{_
�ݫ��ݫQ��M#����mv݂}{�;�J
�N`u.�6��ߏ��*2��^ˆD7�Χ�5��B��Σ��.�=L^>�b��5������>�}	;y�R�С�ɲȬ=:�r��H�b!��U}DKt�� ����d�v��Gw]_��q�½3G
�b��+�)w��� �ݫ� �U"^v�f��|��b{v	�$�ݿ_
PzpD�Q
D�����r�y�&�vF�$�X$�c;v�WV�.T%n^gUƝ�NJ��V	�CP��D�DO�"����A$.�^�Z�e��� @���t>>���|�<�+��Iw�M}��D��T�UGZ��f��m���-w\���al�1���r��P������NYe�y�w��~$��ز�V�bR�'�W@|��*%�&S�!A%P#;2���ʶ��3۪K�)JW[�|O��}�`�
��+���{]��(Skb}�9V<���zW-�
�Ź=�%���j�^�!@	�E!�%�p�m�W��C^�#�q�������Nx9>34iJ媼%WJ�����V̝z8�.p�!���Q�ѨdFao\�!%We�!�fr���Yy!����Nd+�W,6���S��)����T�h��C����:���X�)ŋ,�n�\.�6���u�a�
�Y��������{�d��c��ExN�"�*��[v]��&��\�@�躰[��_a��o_A��~�twk���Zz�U����%_tZ3&w'j}�b�n��p���*��놡8�� nZ�>��: f��@mr�$�sd������2D�t�/>�)��Ib�S���m��j�ʹiE�*�]vNn'q˳��t��۔q۬�*�\�>���}��`A�{k���jΚͥ󖶀�6rخ�!�Q��erӾ���q���C��
�B1(�.�l���f�|�y����Vq��V�pI���e�\�Z�ԖёPѨv1r��[s�qn�"rT��QE�����U�2om]%Ʒy!km�1H�P�X����-�����'JVu�8k7�&&5�i�>�����l��KMR���e��q��wS�!3J���9o���.�L��m��RctvC�-^͌@ݓC	(+)d���S9g&��Dk�#ut��_Y/5_#�-<F�F���7y���t��]f\�	��5*A��o�S5z�dۺ���L�r]�;,]M���s��V��y_p�{���,!R���[Lַg;(���v�g�Q(���Tm�=��wϞ�T����:��Ɣ�Π���Ĉ��;GXG;n�*9kNK1H6��M�f\t��iۣ�Il��u$�@��Ƶ�k"-��w9DH�P��n�qGK+	-tqHgG(�&ڜN:(�kk3�Τ�vb8H&-�>�,��y��̵�$�98��e��۶��cm�!�Q���`����7/{׮�ӄ/m8�5�{�y�����8�;���,ͻޭ�n�&݇6��[[��c[�z��q��	 �'mie�痺w����n�ol�a#��oMID1���k.���n��_V�:D�bH�⤒)�f^��c7�Z���!�y~�	$�\���ޮ��nf/m�x� �Ǘ��(8�"QS"j�y������p�Kr3��!ݷ�~ �S�^����"���+k�Ó ؈.	�%�0�u�v�.7/��;0᱘ݩs���:��'|���*H����]����m����}�u`�..rFrs ���	�K5Q=xÄL�R�ϐ�����ʸQ�-���dII�A�G�츃BڷT���*�@��Z�!H&B�*�B����j�CB:lCg�ݖI ��P�}�w~'pdv�e(%)��E�is���[��]�FʪH?z{��@����߅ߤt1�4�65��=7� o�r�a`롎��_�;����p+���Dk�3��M�&�����疐�Վ�f�Lo8d��
&��!��G�r�$��>*I"�m�]��A�����x0������b�wu݀I>3��b�h�Om�*��g��0��k��\�[:l!��9��#WW��V%7�gFU�;�����~OөƢ��ϳ3�ɴ��uՂ	3��v��LՐ����6��}��K����ݐo�QA{ӛO���"�;�b�'���~'�{{hX1�g��F�@����8Dʅ*L�����2�mX$��	��؊c{mX$���v}=��,����B�L� �@Y}}y��rs�A ��ud��:�n�I&Vr���dJZ�d�)�Hoݒ�䌥 ʂ(����d���\�aNt{+a�o*�$�v��>"Vr�yY��l�ʅ$�/�r�q�m�s+,-�E��;���s���7��Sɺ��V$�������ju,���[�&���*�:T˯W,�(k����s}B�}���B�F�R�"�3oC��wb��r�n3�j���Y�Qk�8m\6��.2��r���q�M�v��n��U��qn[�\-�ʗ[�q������8뇄��O��68;�m��^k���l�s�z�Ɋ�Ou�[l�s*�q���Z5�l��mGnx��t\�!t^7F�����B�/���c^B=�|��WNưNyg]�p��Zo.���[g6�]�An����%���sF�U>r��W/��z;EX)󱶻�k+�I���|	"Vrf�W	W�(��P*wU݂|H3���duN$H�Tț���B�\�b���g��C<I"{y݂IVr
1"N��1͆�:I��3&'�"���v,�A����&��Kl��S9� ;����YʉXC�L��#>Bl�y�t�g>-��A��TO��gv\���ܱ�}Ɯρ&z�߅��E10 � �
A
�R�ʐ {��t ���)z�T�_f4ܽ��m6��{y�'���L��L\s'�v��c/>���u�ɷu���c��ڷ
J�	%SY�{�r�9F�Ny��sXI��x�we�[��ԡ�'Q��˰|I��W��ے�(�	�RI�w�d�Г��fuh��^�v%Æ���ȟq�[j��on�mG�atSͲ!���j�7�?M{�d;�7�f�L3��L�
��x��/[� �*��n*:{ѿ�*ﲪ����p�y[|�EӀ�%2&��uGĖ���A&��V�c^�z7R���+uQnwe� ��$�D)�3�F���O�1�+��uD�|;{�� ��润(ER!�^�s+�uh5�)JS!wWݷ`���[\׹B��o�h;׋��{�1����g�)�徛��=�,�,*l"f���Fċ�p��n먡�J�6+�6��< ��^��>R�R]�*���{�v�ē�g��n�WZMb�Д�a$���ݒ)�ڦR�d�(Qa��1d*�ŕ��@��d���ڿ|O���_�n��5
U�>X5��Q��P�yw�|O��k�dn�%�Jr�&�E�0IWa߯��(�i�¯�wY�-]�q3~�c�Y��!�(�ے���z�ͬW���(��d�]�U�����l�/p���	3��ő�P=#��(��7`���z9+޽�7:|��WA %�;�g]���PW�qy ��]v	�"�3>P���`X>#:�\�]�c\T`$s�˿H3���`�s���V<�WFLV�K7�] �p�"�It��709v�Gl�θ��:����`�z��mj��m�q�(�*Q!\*����e�t,��v����U��@�e�W Au�d�S|�
d@T�x�ƥ8��g�{+|	'��=u~$�v����X����E<0;��P��,5=��$�whP*�� G޳;8H3����|IλT	؝���@� ��n���0�vh�7�I��n��+Ď��}]���^o�vgiI�f�i~�!#}��ܔ�x��}\�%Lٺ�[�s��Y�v�#ZwLm�a΋ѓ��t�VrZ�"���������|�pQJ褻 ��k���i7Gg�ݓ�`�4�n�������;َ�&����$ �o�{���3pl	[��Gn����m���܁�̧`������MxaBO��<���X���TI���ڿ��L]�z&����`��v���;�ofR�J`�.�_w]�6���+�k�L�1@|Z� :v�X� ��O0�%9B�t]1�dD�� *"��	�;��VA+zx�]g���_�mm�P��ۿ[����N;�����_p�|���|���I��P$�����ה���WV9��n����K�o��0W�8ʫ��� �g�]T�l�k�$��ۏ�o� ����O���d�9�s6Ɇe��I�������= ��e�sC���^�O1��8��M�&�(Lٸ�p�=��mǬi
|/g,��� �m�fz$�mvgpKW\��	ؗr�m%d��=;śMḾ_m�է����Q^0����Z�lm�HV�[�=�#�3Ҙ״#G��mCہ{Oh��=u���q��-q�tq׊gJUq��݉M�+��8ݎΰ���>.1'Z��;/�fx�=`�'[�/v�p9��uD��\dy�����T��q�<v�u���=K�\Nyf�L^wcL�d��`�8����K1�4��[O^�w�:��,�vF��! �L�x����Ao�j�4�U��̈́��l�뇝	��*�����&76��Y'�M
{^�1��������<(�q�m_�>$��v����Ĵ���dʐbb�����w]��H2�v��AO��.;UEGm��F�ݱ~$�>�^YtdǑ�"B���+;"��N��H;u�V	�D��ݐA�֘v�3�����|s�����ȁ���d�%1V]u;�	#S����MuLwcK�vO�2��Ń�N.�^5�8�s��ޜ[�!ϡ	/��U��AD�t�\��u�wi��۷<E
F8��a!`ʜ��{ÿXV@�D(>��.�$g_mY$b�T{f)f��E�Bܭ�H3��`_"�GF	�! Q������#x��6��2�e��5����!4	��h�N��t2��6&�./F�fʶšA�Ź�z��,\c�5�X��z���w��ŗ�[\	������@8��	�׶k�5Z�(/� 2��hQC9�j� �U��Mԙ�/4U����1��b�$��D�Qw2����� �-�~�7U�` �_	�^L >�� *�{|Э�<w$ِo ����9
��"���*�hQ�>=�����zV9�m��J�߈'*�P$�s�m,�����O�-�(}_�U�}#5\"ak��Z8x�em��ۋ0v:�s��9�;߁�����/2?���W�H�^�	��}bV�8��o����M�k�t�N��Ք���^��]�}��+3Z���L�U]Ō#h��)\�Z)�lV�1A�߷�1��Q�m)}��罪�MVo8�����\# tM�`ɐ�(���<	�/�tv�II �=�QyG�8�Augﾋ9w����i��^�S��Z[V��t����Cd�5�|���FCB-�x�c�k��wj�jTw�����)J�ڽ������| �> � �|:�2�MZiF1Fa��~�14F������ ��M}Z4�i�2����6����w2J�
b��4��hw�����j0##.����6��Ͻ���m�����A��o����'�CF�����堇V �`�y�v�b����=�Q�0�t�W�k�lV�i�4E>�n�M���g=�Q�CicQ��>��h{@]�E�|�&�AHQ)H^S[��Wck�\F됝���r�m���/]�n��vx����|���'_{Ai�؉ �{�/ ���G����X�`FW�����y�8��ɗ��)�l,b�o��э�7�����C寴�э��_(1�1���w��N����R)����6���bA�1$>����C�}�}���W��Zח^s��A� ߑ�IF}�B�l���fn�f0#PiF�J3�s��,ah�����N����SG�#a�{�[�X5Pj3�{��c1�=M�=��OA Q���x�{q�[Wu��Y$xt�D��_h� ���GA��y`c1�57w�E5'ۻ�=��K�t�9Z-I���I�*E�sz���M4bf�e<��d7^�9W��%*;�zP3K2�� aFu�@�p��K3�i��(��o���0h�kO�d��i���F�-4FW�ܠ���aQ���w�E4��~ΟO��z����{��ٍ'�b>�}� �"80���"���2N\�#�}z��r��SR����]PWZ^m���<,Yһ�7\�J�પ���Β��V�!��%�y1^sݣ���DҍA��=�Q�X�6�4F�w~�SE������V�}6l#g��v�bK�(�f��r��.^�+���|��e4�hw{��؆�}�}&rm���>�wt_ ��h#�f���!�4=���LCalQ�~��V�k�]�p>�v��G��3�l���8ji�i�1�#7��P`��҉���w�,j�Q�����{��k���=y��W�q��Ƃ'��5�{�d�N]��N�Ȼ����ϣ��}5�������ew�}:t����Ɣj(�g3�`ŌCh��4I��Z)��#����Q�)�����$�^��4�5Q5]�@[9C��[z>����f44>�|���؆��7�QyG�zo=������i�h#3��P������e"��ҌCaw{��ƌh�%���w>��٩��c�w�C�!㋪��J�۔gmv.Ν)��;��d�j���:��4区Ϊ���#����uLɢR����lɌ��G-ˬi�1ơ�a������-S�wr�
;nv4(iq�E� aT�*���L��SU��w�.�)��Fa3C�6/e(���]�/�L�Yz�%k5(��M�ݺ�^:��x⥱���f�7M]�΄*C�'h�p$�4ߝ��ʐ�ns���Q��X�U!���u�4�)�NN�ݙC5h1��ظ��,��o�rZ5��ѳ�S��F�`�Ѵ������#7�B<�y�x�]�E��qn�I1�:М{��ֽ��>�p�Q��X��uk�7��F
�ձ�����=Vf��5��rx:�F��:�(�: S���#K$HS�w���_V����37�phS��f������j��tc['"�;�V}.��53�K��/.]�{�����nv5Ye�p��}{pgM7�G՘���e�
��yl:��w��sjˀ�T8�U��!�V��hs�*�qp͍E�)��SՓU��j�)KKN��Ҩ�f�P����N�B 5���ow��I�c��l�au�lH��UŃ����g|��:��ZW$����+�;ʋeu=��m�A����3�x,�<h%�"T�ꄸ�D���	*9�N��}��jp��ԩ\�\��,�����l�z�T���w�}f����5�E[5��ٯT�D��Κ{���ȃ��'G�N��#��ֶ�F:��y�K���tS�	)m�@���#�H8�Q'���;��ǖE.m֏;(Iq#��q��+s�Nv�;[Hy�IJ8��,���NF�DJmb��e�	���y�N+�\	��{u�y�BRb;i��׹�F�e�� ���	гNO+<���G�n�7mm���C��IטK��[��Xf�o{;۰�{��l�Cnʞ�Q��釃֒k�;v�9�����Bh��2���VVݜ4lvYٜ�ob��)�z�hr�Hy��qǗ��8�{v��{�6��[Ld&�d��:�2��/j̸�D��{e�d[ڞ���V,���^��,�m&x�q�eR���Ac�jD�G\q{[��5e�wn���7�,���=�痛����g��L��\��т4��Ҽ{�85ںy7.��XP��EY7"��ۭ�>�^�S��׺���f��s՜�sG\�붸�u��ݥ��:n�F��ƣ��ꍈ���/��)�l��Q�vs���e��]��us��γT.�������m��.5�T��^ݺ�9��`x�g�r�W)��He��;Q��;�=N���Ⱥ4/Y�iy�ǮB�wm�g8ø������ge���\�l�	,�D�=��y뷶���c�nю ��m��Z�84�:�rq����;�GӗMӶ�cu�-[loo9�r�
�޻��p��@m�$�`�M���_h
��<���rݭ�O9㫱�k]t�l{�8�r��t����{]m��;n�!��F3�l�i糡-��Xz*�;��d��{\q�ư���s�X��豂��g��X|4�f^$2>	��������2s��NM�]�S�60莰�v��v82vKi�}pk��(���ӝנ��� Rݓ����;N�6�c(h��7nwN�!�74��f��c���fv��烹��[�/���5�:dG�6@}�����E��<��nN��K�Z��U}lrF:�qI�W�m���mV�-���m�7f��nn9��/f.h�<��n�皶�bӺ^\�Ӹ����T�vq8�]����;ZK�7�q�7����sj����y�n���������v���_6�x�̙� ��zz�Q�ܷ��]�	��-exׇ����g��xsn-�6�2;.���I]7gd焹xx���ۼ���[��XNI(�+6��m��qdݼ��^��w'z�ɮ;r�q���{t|�S|����]=��D�m)Ľ��;��O=��O���ܶkk��xe7 d��av�;��p�݆����.ժ�Jw.�plc��J���l]p+���;�,�:Xp�rؓ��ѹ޳�-�s�v�ݭ��I\i�qt��iؚ�az��4����.�����X�)�2�@��v����xu�֣�٣�r�l��nsq��������<�u�͹V9�wE�����p��4(Me���j��a����Ǟv�k��xGgp�:�;�\���a�[�\\��u��7hF������&�Vŗ�(m�2�NY�p�$��)ť��z�"y�d�X��Y�.^�qmv�����:\u�6���vl�*u2@�!hN/u�a�^��&~����/����cL#J5��E�[JQ����Y�Ch2{��m�rOolF�e{�d؆�	���|����ѿ�]�,nEm:�%���y�z�f�iF����]��}:�g�ٺ8Ō � �$��-�m�#L���Q�,Q��-o\���ܧ��ui����-�1�9~�����}�B�h,hw~��؆�I �w��yG�h#2���ns3���f����@�60#���H��iFb� ��߽F4bh�͛Sӳ�@RB�~|0�A>��o϶b쩻�:��҉������M+j0##o��lƃ�b$�����3�����o��Dq�����h#"���k�>����L�-^���c0�4�ٯs���o;u��,h�N�ݴSجa�g9���b�X5�{��bf05�陼�|�g�Ug���ˍ#tk�>���ϕ��pN�;[��q�'K�ۭ���n��~O���c���'��_�h}��H�"�A@7���^A�n4����ٌ�=����yu��z��ƶ2_���jƔa�0���Q��!G�w����2Ѧ!�ﯶ�G�{/�ٝ8�����a��y7l|l9�*�5����\�puoL�l��FR��Gf#tU�.�-�"A&�=0#��ە7�4ʥgB�_+hu��E4�5d`C;���h0h#�DR���� ��{�"����#,�ͯ
6|���1��#����_;�-�lCb&����Ō#h�Dh�_{��9��W_2����)��Db�#f����ibj4��(�f���o����}�B�bC��(.����oR<�!����v��"1Ƃ2�}��`F@`F����R)���W7/���8���+=�э4F�gM����>_i�1�#7��P`��ҍF���Q`մ��w��^����{�t�������`�A��s���AA�a9^�E;h#2�Ma����/�?8�q֨�X:����{���V+G.�t>K��7"�51_������k��x�1o�̣�5J5�f���b�b��4I��Z)��| �O؛�S����s�=�M�t0�؆��Q5�w��b�	�y�lq�||}5�1��q�����b��~�?�'z���Mw=E�#���d5�{�3d`F����R)�l,b�/�{k\s�ޏz�Ofz��`�(���2���e#M4FW��Pcb��iA���^�E1�lJq�����-3s}n�VcS9�����Q��]�d���j���Bx!ҁ�+��n��
�<�Nי�(�_s�1���	s���9��}���姏䆅��]�lp��X�LW����x�o;�W^A��M��kcJ5Q���F1c����^�E4X��a�=���cKޱ��KX���iA��r����o�n����}�2SAiƇw�R)�lE� �w��yF�\�x�j7���6s^���6m0#Q��ܤSV4�1F0���Q�Ch��0{�%i�rMB���)ml�q�]����	8�ǋ��p�by6��J��Sx���~�~���u��'�̯r����C�s(����#�߽E��A�g}5����{�s��1B����A�n0���"���;����ϣ��MB�l����2�f0#Q4�U���h���S���M��U�����6�Nz��LCb��b�gw�z�icQ��K��ޭv��mWk�{^Ze{}��f0"ݎ��9�Mj�h1Ƈ��(-;b H"H9�z��"1�l���59��z���]�l�0##4>��MXҌ �@a�߽F4cDh��\�D�4Ϡ�F�-4FW���w}��������P���H���Fd`w��h��h#�Cf�����k��^�ۻW#��X�AP"����8PY�P�1Y��@��ml7��^Yv�Z���_թs�a��t�g3rcT̉���a\9{{��!��!���Ԋv����{e���`4U�-��g~�Ƽ�#Q��iFk��h��5w�S�=߯����Ch➮e��-�1A�b��｣����҃Q��=�&cw���������zi��
�p �S�]�Ŝ��������ΐ�6+�S�ב�Q��������}�2)���C��)�Y �����xAƂ1�k��lb8}w��ɗ�U�:�&K��H���A�0��o~�э��kڝ����}�hƌh��׹A�1�0�*̝������6���u�[V҃Q��߽f4�A��{��lC�"?����}#��'k�H�!��k�6�s�H�7��`6;�t[60#Q��J3^�{F!�������=���=�n�����h���F(�7�э,j1�l׹�б�������ǯ����kVcA�Ƈ�o���>s��S��b= � �s(�"84��FE��ݰ1�0##59^�E55��;���^�%�C`}����64F�Q����vޙ�h���=������6���Q`մ�����;5z�ϿO������w���`�A�"Hk��h�!�GNW��N���͗�����#�uoH:Kܓ�f,�ս�6~T/�w\���w]����8�(��]�(vo|U����MgQS�s�(~��wWjx0n�X��7�'m*	UQ�qUeV�r�í.��rnq��yt���u�p�n�����@��
�-�+q=r��� �I�*A���h�B�������G�:��裻��([���ٹ;z�h�B��;m6.7A�<�vƇ���P�k�g�n���+Nynk���<b�n�k���w���c��būY�bXy�/;�76襉�\��Ý�Ӡ�kg���m[���\qƃ�뷪����TX�r���v�]�ｖ�D�����,�w�c10#PiF�J3]�F1c� �+�H���ŕ^�k9*���}�������6k��hX�`E��4���M|��h��q����툄�2t��u��c�:۽���F!��ȵ�w�3bPd�{)�61FM�{��G��x{yC�'�/C�Lt��0O��v�hƈ�e{���҃Q����Zj؆���k���w��t��V�48�G�H}�{�ADh|�e"��d;����ω#���e��hb�yF3�~,��O�5�� �^iF�Q���bb�!������h�����o��Z�}��sٯp}��K�F!�[��B�cz�^��NQ�U$ŷ�[c�?w��X�5� D	 �7�QlC~%���h)���������c20#C�{)մ�1F�g{�1�m�'׭���v������s߫ǵ�8h�q��c0޷5��q.vq��v[�F4�EuX��uxl��q�&�|�G����w�a�PaP�u��V҃Q�#f{޳��M;�k3��5���~�	f�t9F&��{z�i�O䆍��nZ9�g�,fY���c1��J5��u�7�В2	��7���T����(N���+\��̻᭺2�L��Ȧܵ���ǐs"E42f�l{"��'�zș����m�4=�r�M�����E��j4��i{�G{�e}�U�����y�� 뜓H��		�$P��X�C��(-�$$������#��G��wy����[����{�l�����d�_)զ�a(�0��F4bh��^�Ӈ����6V���5�T��ӽ�~·���4�Q���n���j1��s�cA��q�l���h��9��ڢ�PDhu��"�������'Òho�2�l_��m��J5�����@�Јv"�+��y��N�=h��M�0�Pf�}��ƣJ5Pj3�wݡc1��쭏;X;�y�o?r-�'�8�GGHImK�<U��mVN����U�9�``i�����Ǉ���멭x�A���PX툒�@9���� ��7�3�sݠ-������|�����5J�e"��iF!���{�cF4F�:V6�=3�2���h���}���1F����2�g-�u|���[�d`N���1�m8�I{���8A��o������ڪ���"=�=�KNi��S���bb�{����(�iFk��h�,ah��44��Ә��6��c�P�f*�v��e^�� �V�r�Nh����Y-l��w��2�{E��ƕ¯-���Ϲ��Ze�&f��h�Db��f��Q�,�CiF�5�{�,f0!��#y_���#Qb��,c�f~�H�x��Ϸ����b9 � ���/"84���׹���L�0#Pg��|�kX��Ws_G
{{K���{���64F��kڝ��-C��v�hƈ�����iA����������u6��ǯ���|X��d`C��=f1�lFH}�w�� ����s>E�$5���l6Y_���G=�$�Yj�A�)뭰S��.m�͐(��D�UPT
��￟:�d������g�l�����f�M(�6}�w���(�#D_{�H��h�Y�}�vו����`f��Qm/Q�m(�g��{B��`E��6q:�URI�o��˛�X�5�!��n�7ϟ��7���-�6!���Ｑ�0i��o�(i��;�o�w��׻GZ8�#F�m��	�}R4�m��o�0�(0�(��z��(�@@5d��L�7�H˿x�A�Ƃ8�BC�w��-�yF&����,k�ڛ_�7j�nP>*�K�,�{�c5����Y�S�w�m�4�PiFs�ߨ��A�4D�'ݿR-�ƈ�6(�{�F4����7߲���m˝|���/�&�ӱ�b�F�87O-���x�KR�?t(�4#�`���̽Ψ8"�#�{�R�YAq3�k~[iy�҃Q�ow�&c��i����O�5�h������2�i�؉ �{�^A�k��j���*�h1�h#'��r��c1���j�Q�b� �=�eэ�U]���_z���?�;������<훬�An�xs���!�oQ�;iO��}lf�/�u��ƨ���]/��3��r��1F�m�ߨ��iF����{,�!��͌���w�������$=����#�[{^G�"�܅2��L�
�, H�����f0#Q�ɕ��_;�f���n�q�[��-�X�Dh�}��,h�Q0�Pg��e��j4��>��u��z���o��j�������>z�ֵf1���Ԋb9 �H9�e�Mb<w_;}�=݁l�d`F��j�Q�b� �����hƈ����ܶBi�A��4Zh��w|���W��T��6b��Q����E�������y�؆�`��{�� ��۾����y���k�H������[��SOS�"��+���1�0#Q��(��=��{��oC����Mh�_fR)��Db�#�ﲋbK�J&�3��(X3���k[�՝+���E-&���1h�k(�W���g,�MI�vB��<�j�Y�U��F�Q���-�َ�5}hNY�\��9�\��8WM�����F�d����(7J�ێr��4@�3�݋͑dx9P-�k]!�q6]�<P��5y�N\�ڌ�uk�cv�n/M�Fx��'G����hl��<�uQv8���;;X�׋�z���sk]hx���n�<�qp��b�獣�[��p�l�.zy��N"���Ga����qn��Ѹ��7ښ��v�Kl����-�(q�#���u��9��ݞ�緵p�]��u�=;:z�Nm��/h�I�:n����������Zf��y8�����	I �{�E�Mph#"�sܰ1����ⷜ��{������<��M]z�MXҌ#a�=�cF4F��ف�vH}���1�#;��(0a�PaTQ�h�j�wkM��ƭ�l����h1�!�C=�r�� ��7��w���e���}���Oɠ�F��!H0fH*H�"���!�iF�iFg��Q�0�� 4F�������u����Ѷ��F(����1��Q��(�f{���	��nL90��
L�X��0��/P[�u�km�5��jA�^_h� ��A��=�ٌ����_)�iw���n�{ޞJ�m�0�;�s�c�18V��L��i��#+��(1�1F���_(�5m-{d��l�}�1�U�g�ƃh �	�}�؇�Dpa>��NƂ3Zu�o���ϲ\��[
	�����U0��}a��h�z����z�9��R
��t��U7�����°�|xg�.���1���4�PiFgy�Q�ŌCbDS�_-�6.}�5������rp1����F4��҉�҈j3=�r��1�7\替�����zZ,��Ӎ���[�"H!�}�oL��r��	�KY���w�l���C���p.��FA�@�����ѰT����6f�f3a�n����ɘ��g�hŗ����W]w�J�7����ph#&{�偌�������MXҌ!��S�/�e�+@uN�i��| �E�����>�����6w>��b��4��hn�E�m(5��}�����ys��{�4q���D���3 �a>��N����{�F��I1$$X �~#��c��}Z��ޥ�����o�m�mtiF}}�h�,a�D#D�v�h��#a�9�{(Ɩ���5�w���iF�;��t,�����#��k��-�����|���툒�@;��(�!�w����]�JݕW�q���W����L�>���M[J0��D��粌im?��W�3��f��׿{��!]�Z6�p������#����W@�-����Ν����d�!4Ϡ�#M����ر�iA���W�-5m(�b{��Y����=��s�9���Z�o��a!���� � ��a;W�E;�ߟgeP���X��[M}���ic0`F�J53��=�5Ux�ٯ{���0�b��4=���LCb��b���=�cK�(��'�������WX�C��C���{�#��&������h-4>�{��lD$$��wE�Mq���{��<�__��ֵ߱4�D65L�CD��oA͹d�����(��r���۠L:h���̜-="�U� �@�fi:QW�e��"�A�r�,B\��0^f�N$��2��}��e�s�g��7�fތ��s^]A�ݍ��!�ea6�#����J�:!{�ӽ7����4�TѝKaU�Zk���l�l�Y�]��Z��:b��a��E;E�������fo�t�k���,�FV�l�����)���gV�h���ns,z�S�@%F�5�Ƈ�+3��2D�Ŭc�ŗ�Ա,�jY�ˣ�u�|D����t�C�oe��y�VM�Rg4��Jɋf��޸v^�����69Զv�v��,�]ۗ�+�T�o���u�!t�������UB�b�Z���`�b�n�n.J���y<;AR�rXܠf���Y�b�������b���S��w�n�c;��2j���k����j'^=���Q������i{6@�s~���m�sup�]w(� ���`^��FX��ngW+��'�^876���osݥq�Ŵn&���u�7��04,e�d�N�,�,@�,�P��8�55HR�e�5����!
�*4�����z8���*�����<��	Ar���y�[܍���3/r���qh�;�*�p]&թֵ͗�F9`�u26��N^8������6�L��[��q�oR\:&pC� ��B�V��$5a���ANQs��g]2������ҖQ����F�l���[B�$gD#|����N)��,�8��#M���ö^�Ig���޽6�Q���{[�.w�����đ��8N�)$9�X-�����0��^�o-�6�V��u���Y�C6X9�hX��E��'�αy����{�{VՌ����f������{bR�jx&�9mv�Y�u����{޻��	��,��g3v�����'Y-<�-��q����m���y�[�HN��ý�=���6ݢ�KtkN�3Y��{���=��v�iM�ݯ='{6��٨�Y�a�l�{Oug7m#C����[l�sy�k��[[I�i�d�<��g���`�m;ۜ�m�og'c������3m������@�̼���B8�Z�z�׷�����dC59~�E5cJ1�a��ۣ1�4A�����(�(��a�����o9�w]�B1[ҍF����Zj�Q��6[�}�1�lCb2B���y�wܯ��x��u�D>A��j딊v�F�x�QX�H� �$�ƾﵾim��j(�iFW��Q�XÐ��^~+�شуDh���墚-�1A�b��y�э,�(5Pj2����}�{~zǤsk+N)T�V(��jq��U��9 �G-���]�峺� ����M��vև���SZ�1��پP[�!�H9�v�bƂ8�FJ�{���߭;{���֭�9ˤSVҌ#as���6�֞��	�!?��F��Ͻ��c�W��k=��w�ʙ�{|;��|��_��&��l���o���bq���	
�{���#�o����<�t=����6o\ߦ�5�M}$O���`�y�z�f�iF!���r�b�!�����_5�rp����ƈ�6(3��{F4���6���s��`�`Cu�i�Z%(�(����h��&{Nt���"�$پ���Cp�]�y`c10#"`F�&�yH��:y�~Gn��Xk
�c�7�/�����7��W���P6��Mii���[���>�P��K`��s/�fuwX�7��뮷|�i
B�0�޲= �_w�1�#F{m����kG���э��{���0�(F��^QcV�{y����{�X�6���1����]��@[؆�a7��E;Mg����9������z>��^����x��E��N{9�M�;�c�ړ�4�Z��:n$�f��:�)&"'�&�G�y�X�a0�ҌCe{�����m�4@��e��,h�Z��xwڭ�1pen�tc�X�b+}�(X�=~r��5����>�Գq��7�E1��N��f�w;���5���^Dph#�d+��lf���DɿfR)�iF1F��N������T[F�#DZ��!>d!��h���}�����Ҁ�h{�e"�V�`FF}��7�e����ׯ��Lh:4�"�w�d�L&��H�cA�o�[��Z&��'�@[1�3���U�����)Q�=o&��TҍF�g�w|�,a(�#C�)�6+a�3��hƗ�o�*��LV��j4�P����{@�d��HEJzE
>�hw�n�ݱA@9�w�^D~��޽�֍�A�cAW�v32�;��E5m(�&(�3�x�)���7#g`�&����X�&�Wm�6+E���z�h��j��7X�H���hJ�@�ڙV���*�"ۙ������
�����AJ�Ȝ�{uȖ����tm�3��KAV�B��!����Z�zQ��+t�S�Q��5���-�������m�K�ty6 �-��]yˊލۃk�7tl���[@���m�q�[r�:H�箍Ȫh�\��q�:��C�����sm�.��Z�|1��vk �i�e�k������V���ܥB·P�}U��ۊ�^��n�N��]��H�v禟E��Y�t�Oo#�\������[l.�Ocj�#sK����w��䷲^��=ߧ{��}��~�1�#JF���Qm[JF��ݳh+*�>��z$��ڐ�{7@a�C�Dpa;}�|������^'�+}H,I6�����ь�j&�k�:�߾z��-2��z��1F!�Bz���h������F4�j4�Q������pڶf���}ֶ�B_��͌��])!�o�Ƈ�����C`o��h�PDph#٥����'���u�h|��"���b;�v�hƈ���n�O�nA��4[De{������:}x�Ŷ�Q�곔�i[Q�l	�s��8�E!^�{@w��әS��lC�"80���"��ˬ�&�4Mh־�'�`c��΃5�j(��=�11cS��eq���#Dh�W9��i����զ�{���'&�����'�[+�R15UMb�糕�ьr�d`:z�\�mK8xz��OB*P+�Y��F�7VH�]��eu�f=���]�/[w~)�#dƅ>�X	U��7��{��qj�u{T.j�0��vi�L� �-���Oo����գ��Źop��D�e�-����4cm���Ŷ���OA7���H5����kjUx���h��yHRLDO�Lz�~q�> /v�b� ӮHU��>X�e��!x�������������bd�AF��
�:��wM~���\���|��'�����{�)���tꁯ0������⻵ՂHδ��������Z���u�'6�j;sGo����� Ói#���*V՜1q���8�X����x6��AЊRZBк�p�"��`|�ש�{́@۾o�By��2���J�]�vA5��98�׉EJzB�Α$�U۴iD���H>�����lK��ݶ4^�Ǭ���'�B�1c�O&P��y@
;�Q�0b�V���K<�P��6#�L*ݢ4e��D�{0��ɤR�Ok��y3��~�A?�p5��⪙,��y���i��zn"��� O�6����r�ݛ�$�o�6~U��5ƽ���P�ny0(
�Q$�{��O,�}8"���N7�W��h�9U�f5�ݭ&���5�3�Uq��C7�	�r�$E>�b.Geֹӑ>��	tj!T�ֆ+k�j�@�u��^]X���n;�ұJ�3��~B(&(舎=�~�	#:� �|)�;�X)�=|,H5��g�>{%L��L"�������AuZ����r�_A�w�P[��ώ�na�M�؀��X,���3^%(��
�\ׂ>!�7V	 ��2v�Nf�X�4��O��Q �{����fxNʄ	�H�~;��SJ����<H"�J� �o��~"��������qPȒ�h���G?]�b����ZS��.=��:�Ř�mrux�<��ׂ]���F.�we+��Y{����ښ������������>,vv��	�wlYۑ�t�l�
����D�=�?���/o�}
�RvEeuvA��2=#��Õ����mN熚�<�nҰ�x�g�l�zr.�D�TrI�&���^s�ޯĂ+_mY�:!��S�klf�=�(R�lo�>��D��0Т�g�rg��5<�=,SoȂ�˰&��ݦ�䫞/��o�Wu鯓g��l�7
O�t��I���A%��
�y=�P$�w�.�"��o�Fe��5�QR�^���u5	N>ʾ9�M�wU��I�gv݂<�iFҜ�\!��Yw�V�舞���0�,m�e2A���q�k���w������x��~TFgښ���L���!W;��d �k,�1l�t�Y��%ҝ3�ù���p���VC����˕w�|$v�r(�WFW/1��׎aÞ{u�=s���{ƴq�7qE٣t�QTա�7������z����X�R8���;���|�j�x�f�=����c{�=�H�i�hw6� �	m�L��c��6�n<Ҧ�Q�]����n�$�q���czք܊W'n��!�g��ĕ�g���k��{Xǔݷm�N[��&[r<�	�=��5i�S�fz�hx�Mnju�툱sډ�"i���M���^�|o��Ȉ�T�vӼ�$k}b�$��J{oR�S��݀H�\�زOFJ�H���I3>k]�J������QMH��b.��Ċ�}vO� �R�3<y7_5��|}����m���&AQ4i4���$�$I9xC�D�����~$k}~�@$jQ>\�qI��!LǊu��{w8�&��nj��A'�H@�)�e�N�H�u�/L�^�e幓4P��!QX� ��U��}����~ʾ� �C�!O{.�(��![��rޞV��P��z#��H��U���A�e|��¼קW	G>n9����:�=e"jYD�~O��d���DM=���t���|c�����ԍ�D��0B���������-α�+�]r`�4�X�V���G[�+�������Z9V�����z��4c�Vj�;��WIY��G��Y�Z5c�(K�޲	��(	�ޏ�ȍ�W�O�A�S|eӣwCPffnȮā�}�`	�!����Oc�|[R� S�˲A���!@10"��{���C�c�ˉ#{����X�[�b�:�$�v�AK$홲�Ȑ��
����A��n�!0�8���d�ʔ	�>���H+����7��]�R���5kQ:�p�5k�x�N[�k�鞮��͵����]��k������/<��mjD��yV ������}��y�~3�B6��	s��P�۽�ⵚ��T-��`D��_U�	on݂��5f�J�8>nh�JA��~U��l (g��}k.��ט����n�C�2�3���-�ؚ���b������z�̀�.��3���s����7K�;g�_=�Y۽�pՋ};�o3����S��ŀ��,D��"��iz w�]�����	���(�����$�&�����u��|��'�{��7����嘘� ����5����$s�U�g@�۫E�bH�"��u�d�#�� .�g+7������0G%���W��q�H�w��2��;h��mcu��u߹'�ܑ����#Y�w{[�A���+� �殐/w9{=A�C�^��`BC=�m��mط�2V��\j���A�C/��.� ��f�I?;��n�?~� 9xb�ٱ'wy�|��}�R���L��Ok|� �˭�^�������t���y�	 d�3 >|�j� �{���$i���1�*{'޺)�l�O�Nu��$���]o9�{-�d�ػ4��UW�Aw����z��5���Y��.rWk�m�.]T���g5���'�ؔ�@/m���b�n����)��;Bb�������rf��ň�;]�0�לK�M~%��9P�6��ʼK����D����I$�kX��TH}��*��'��4�B����C�vC�h#�ēê�=,�Kd������`Nb��[�d\���� >���Z >��o��N���l��^[:��� �]�H�wRLbr+�u��w���S6�Q[G�Z�$�D��~$���F�Nj�+fߓ�d�I�b��Vd�Ϣ��Z�u^��}�w6�|���;��~�|�5BkX��E�o���{�}�t��e����o�>�opր
��H��O��{|��B>�j�co���]�|�N ��ǟ$w�vJ�� #�α��)/k8��Mư�j7ك�D��~��yZ!���\��q.n�\��	I�x�$��(k��֧�	��W�Fή�l@��Z폑wyw/S�58�i�t�,��V�)V{����Tv�<X�an�&�`�Z�_2��)_w)�1�ؤ*`#~m>}z�ߞ�v�O����`��N|L���YS5�j7��Eky�)�܈�7�����,���{���f�0�b����6�htd}���� t�ڐ0S�5P��<:�1�����:��6�8�G����n�w*�{��v�j�L;x��h�- .��,�Wqv*��4�w@Vm^fVڻ���\��A����9�c�Ά����c������U%�a7�f򊉡|�pw�+7{oOt�zD�)�+;��w�ئ�ד�ݨ�N�Е�fV��� �3t&5�&�h1�*��r	]nÄBWyH����o*52suu#e+�O���R�X�Ѯ�*������$�;�jq<��^G3�1A��h�;Fm�&��lkk+IV�AnhX�Է�jqE���ST���M�ȭ�WBذ�LGݐ-�C�.����М��8��74h��c�X����Z:t����T�e��I���[2huT��$;�%7���cg..Dsrי+-m1��A�Ox�R��(��To&�WV��2��bQ��n����*���tX�b��<�l�w���9[t��	[�2ceI��7yx�0!b �vB�cIY¤�j�'A�4 ���2����Ms�|��.�%V�;�nE�����:I�$�<jFOQ����jٳ�{V�<�e��if�i�6��ml�q����v��oF�lb�f;v��{yfP�d��{�����K�s������x��56��{d۴;�B�m��+kփk,#6;c��+y�;c����n�9��v�ls�n�,���Im��-n�ٳ��=6�[��3;�7��7mm�vmc�on�mb{[m'���m-�	&ٱX�8M8׵�y�b��akm	�y��ô�����^Xӣ6m;���7kl��R�w��9&ݭ��%���'0�hk;#���8����o4�ͷ�����i��g9#��bn������tem8��oK6�k7.sl�������:<���^M�rYm��Y���3���aŧo0���oki�m�n=�øx�<����m6&��C^]�M��uڹw.���xw[ �9�۬Y�[���C�9@���٤W��i6k3!�@k	x{.ۭG`;u�N�Y��l\m��n�sώZ6�^�;�i���n&�7:X<�gK'OIǡ�]˻w@��DB���kv�xm�tݒ1��f�e�<�G+����v�\o#l�ͷ\��vSu苫����� �Əh�ͷ��8llpoD�KY��:M��q5��q���E��=�3w\��i#���+x�]m��8{;pl^|ݰ�y4�n�'s��)�ܻN�ZS�JƇ�q�=k����{q�5<e���}f;g'���L�:�9�xP㝡���@���kY���F����#Wk@g����냮y�(��#�v���|=�\̺�;n�m������ �:����=�V:`G`\���T�gI�OW:�tVPQ�f��nXωV�[�����tF�W�y���ڷ��mc�QSn^�6E8'u�����`�枎�뮜x�nGN5fѭ%��mó�C�y��U���<o)�����v�������3��]�v�`!�|'n���Y����֭�]�Ab�.M�u���B��a��ßnNВ7&خ��\�-�ktn�rν/�J��U�0]��Qs�U��`�z;p��;\tKF7c��oc&֎�\q�<�+��^{�&ݰ���3q���<Ѫ�U���=��2�<8n96�qz��1�W5���5�9ݶ�ka0-ū-�+�cv�[v�%� �	n��@O4	.W�4O��=�s���պ�<H�U;Je8ꮽN���nc<%����O���S(��]7 �MF:�����'a�c��ݸv�H��=	E�����G�Xݢ�y����G����G,�B�ݷ/n��a� �q\n�=��	*��sm�:�ѠC ���ܦ껯
)�좖��<s�ݭ6�-���B.vg�N�����xֻ��h6w#����Rܷ/I�c��n�d�M\K��5Л�y�ݓH�{lv��Ʈ�����+�L`�n�%��6���g����g�����x�@�-h���D��4WY֣>�.�֢��]�[��m��xag��n}�f�����$\��Gc�!���[�q^_m�z�v�:�t�8Rn8�A��xx�S
l�m��/;q�� �q[��7m;�ɬ#�mm�����wf��v�nܖ�1A���U]�'sv1:.r���w8��3@Uw���"�ENI������h��j�*��luoo��5�;����z�5t 	�y��l��K�6k
v�^�`p����@����I�%��6�M~޶�$���P��d5���	�ԓ�)�3g�������+� $��˾�|{�+������gn�� �~޷�&�M� b�L�B�wm�m	����r#n�}	$�U����h��/$��[�ӀR^���Ǜ�}�t��e��X�����h�D׵rl��LT
��F�~�?I	 �{�� ��y�M2e�w�P �q�FmӶ��F�n\�Nf����]l�ͲsF����m�o~=�h�@�u���=���	$���2I$o��d�-�{�x��SH�;��lb@�{��y��"�(�&6�u����<�~����n{�I����y�]E�[��Vn[���Qv&&{<%����Lx�]ˤ�4��y��b���V�)�͸R脣����#��;��gv��;3 '�{3M�����r�Y�/�*���:�D֦ ќ���-�٬X ߼�Wm���I��&�4U�}o�A$���L����&1����1�w����{�=9�tб� �N�h��w�N�$�o��l����i���LX�y#���ـ_�X�^�4 ٳ�T7����B�̌:$ҿ/[I��4�$�o�������,��v��#vAX+�%�:��d���xN3v�eX��NұJ�*�o�O���5l+e�p�7��`/s��<�"����#)�^������ W��'���N RQǈ�w�o{ �xwCgQڔ8�s��h����$�h���*8U��	=�h:�x���aÄ���5��tɪ$�L]�lJ$�+f�m�����;e��R�lL�/�i.�K��X�Q!s��'Ò�Է�F"���Y��$WY�����O���dy� �;/@��K�I�MQ����ت���4�dZ��Fs������ٻ^ˋi:$�ScM��]�ܢ@4U�z�{լ��s�Y5�D�o��"�vZJ	�c��=�[ �s�(;����߇��i�$�b��!�E_���9��>Ԕ��Vo`ڳ�v1N��w4�uu�v��sn�zI5����)kP��A����o�el�+����,o��;�[ >S����#��mC���9>=�:$�L^ޒ�%͡�pfX)�L+�w�_��DE��R�P�خԺ�$�yv�p�TH���j�97^qCZ���y ��Z')h���s��  �4��I��P�y��y�� �����{ k�����Y��Pfn��5�����3��S=㤒^덈I�B��L��$o�ڼ�?~^��ѕ��e��b�T��1��I�����R��~�G����۰�,���E\�9*��S(>s�V�K;��q�ۣ��/Q$���*C4�:�"�k&|��9�Z� [�����׮�>8�ϰ���'ĀI[���A@'�k٦���3�WR�`X����oo;�l���f�g�ef��=>9��ͥ�6�-b���t,��A8�x�{��=��={��I ��?4�g�Oa��n��@ .���'f��v@�����7���l����q���&��$�$����$���?4��}kԨ��`��:�4�uv]Wlm[
�s���KX {��g��$�x��[u��� J��@?�5O��f���N R�1c���9���`��>�S
����f�?G���� 7{�n�&�� A�f\X�],�H����ǈ^���x����ٵ��/d�o@|g���g��@ 5�������r���A{I���Xӹoy����0�bis�E�I���S"DFYF�u�5v���d�8���^�̶��Ӟ�\�G���C��s���Е�yM�ծ�;v{.0�j6��aQz�8�^qr�u��{[ۍ�Ņ�nɷ,�m����\�:Ѯ�`ێ9���<��k���l�ǳ�����6�:f�mm����A�-�h�l.6�z|�mŒ=��`tv�p�;)&�S��f���Rn�ݴ[���q��\�l���m��87\�uy�v۪�!�o!��Ltq���l8����np�utx��]vyz:8f�{(�X��tv����w�G��F�l��ks�����-aD�&����I$���n�9et���o�v��{׫؞���`zԑ`Y%��h]���*�-�k�W/w��}�t��#��N�?L��I$�x[�9>s;ۘ�����`�J�LzBn�/w���TI'ٻ�UBh��ig�l�ٚ����I�I&go����x�b��ݤ��fﳏ���4N}��w��`|�׼������܅�^�guw]J�D��(ӢMP�{�Q���|o��7����z�t/[�{���MOF�h�F���!�5�r�M-�����m�O�Ϋe,;NϷ@�@�����`���&+,�Q8�@��]yp��$��HHm�^�o3  ��=�� ?J��%J\�ɥ�l"<�4�D�N���8����N���kS��=��XD���Qz�c�&n't�X�q�1��3����j�|R�.�Ԭ��I�n�ja�!��O:��p����@�g��o'�KҪ�\�u��!�I&�{zHI$�+��l�L5�*y�,_x{OF]�Z�kzԓ�)$�8�Fb39��� �Zg�M�����]/ܟĒE��}��|�^�.`%�p����}���{��AK�O�i�I��󐚢MkTM� ����f�����o;���|�=��v��$��0}��� /ky:ex���=}zOy��&�$���/�O���X����ut=	�ҍ�Y9�z�OL{\��&�ut��#����n�����;<7^�g:�)]l[~9��7�`$9����$j��d�{�;�vt�6Q�=�lm���n,�W�0rT�$1���q�@�IWa/Uܻ��P�$�K��0[��O�M�����u�:/{�MS���:2
���3}Ŭ���k@�{�y��;0�%צ���)Ҫ��/[�$�)���2G+��D�OR����i�R6���Tӧ����r�q��К���:d�����c._{Zo��I>x�����f|������m�^���x�s����5����@&�wѽ+�Id���D�w�m�]�8a�쭟Us��٘  ��;�P���k����&��zۢMS;�tI�N����z~�<��w�c�D�����M�&�V��v6�{S��'R���y|�@�{󟢮��*d��̸|��_������3 ��x�=���	5�M7��{�i�O���E@��bǆ�����gy;r��)�=������� ���+�A�{qf�*7Gorg��ϰ��r���)Imw5����$���s�I hdE���-g�N� >|��k���=���f���HlV]
v�%��U�ůjD(�D�Q�ɲ�ML��!&�%_���غhE��t�'��IW;uhm61��&�D�8�w��,��i[M)�8c�yiv�ź����C��
SjB�z?e(���w�z~�s5�k�R	�TrVDDc�����$����c�d����˳�Pk�i� 	��r�h�E_����gzs����G����~�ʣAUU��J8�t[�s��\8m��%5���z{K�囍b��~~�����X�F����MI�n� ��}m��R�U���L��#ٻ�UB]���Uآ��L��:{��p@a��xo=|�V��Y���������@#S��ŃG{}Þ����Y���^@?wݰ���ŏ=���� ��zi�A����zxn�؀�M�����E_�����^.P��-,�ǉ��➫��ʷ2[Ԁ�=�{���6ص9�L� |�y���ҬtI�ݻ�*��g�#V&�00�{� w�֞���n}�U�)�uo���5�!޷L�+s�I�=�۰�WG8}����r�1��#٤Tu�4w�ܑ���igZ��zo� �侚���w��;�8��0�X<s5;z�߅���O��ny<��2x��qWkc�Ξ$��s&:�]u��qx%�ŰE{N��!�f8��Y�.ű�6��mi��K�h*��ܼV�Q���|��SOZ;i��K`y�w.��5��Dժ��e��Q�zy:�f�A�<V�g��'9÷O���k-�d��/<"����O��+�e{Y�C�ӊ1�8�{'�v����X���Բ!�\��I��f�ͽ�vۆ�ua;j�TȢV�Z���H&��䬈���S��`	D����0��缓'vS�=v�
5��T ������Q�L��AQ��D�����ؿ@��j��К$�&����Ě��L�D�p\��f7s��]γ;!"D��@�3���s� ם�,o���6L�xS^��v���Ń ���٬���h�#�lX߹����I�.�����2I$�]�~$љ��}�P��٠{z{~���I����×vPtk��I&r�9P�B���&h�.{��I'��i�I&r�IU��b݂��BFׅ��MH�&�vV�����v]��gv�"I���7���ӳ���}M�1�t*_Q!NX�?Q4�:d�D�fNm�{��y�ӻhˎ[dH��4��R	�TrVDDf#]�=�{@��^�����i<d�"���G$R�s�0�3L^1p�Ǯ�ӕ{QJy�흐�%���4�����:�чv��z�L�V���s� ��٬@ �\�� �#7���&n�hJ�7C6H����Us���0�k��{�ŏX�l������ ⷞ2I"r�9�(���U���S&�Oo��Vf�]�V'��MI$�r�I(��&��{��$J�,�ӄ����D��jaDJ�t.��>{�$&�$���X�8��.�z-�#� i�tx�$�I=�z0'�I��ݳ~��;�Qɩ�
o����kb1��q�5OK��pa� ggv�8�f�.��9Wl��C�<���Z o}�<�T&� �������i��-�5�Y��|�=�{��Mn�&�q�co&/��$��7Z��2yr Oyo������vb���g9���o�ڭ�K ��d��"#N�7�������|NVo��5��KRrz�g��Լ�S�cGP�%zzo^*��I���״�M ��B�3�.�j.^�����N�,8���m�r���QZ�k�͐9ތ�ot�;pe�r`� ��U�u�*wќo6��;w�8��e��o�t,01%%�/na$J��F]3�O7�zu��]I`�b�\��u`�^0���,�"��4L�J!R[.ĸ4ov���37h�R�9V:k��<�
3��]����luI�;hF�u�L��J�{��I�O^F���F��S�/ s,�4��O��{�]�e��ACy]�|�HK��ye6BO��ٜSu��h�]���j	�@cVƍ����FEn�DD�;�Fγ���佔��B�ii��ì�����ݸV��M��1�ж��&!J�n��0�n��4�-�CE��bZ��Z^�g6�V��,G6��eޤ�V!��팂�k�0%0�5�%ʆ��l�R4]��uU�M��Ք7�˩@�΢�(C�P۾/��r���ܶ-9v��h;���ۉ�!����3���\M�x�:�U�{��4]��۠bxN��%��;3����>��:t��p�J�lE8n�;��}ZΝ�z]a��.�(���&�nQ�ˊ�d�`�s�a�ԡfXm��P�g�n�N}{�'}+l�v(z��a8��NXs���]�!�w���g7��m��V�"���c���OM��ok%:�GpJ�ɱ敎�vf)jl��^�7(̛ѪT�q���᲌�����njl�t�k�-���c��)�����G�jske�u�fdĀ��T�ɴVQ���{I,X��W��CXխ�o{���e�b۲v��V�ڋ;m�6�C�4b�E��xD����l��m�\�.�-�������ý�^��^�����7����y��m�H�I��4�:!��̴��{{z-�Qf#��0�����8�;�i{h�n��:��
ɫ"6��՜�%{��ͻf��םy�Y��ca-�2ɶ���{i9�iu�$[޻�5�m�6lvK޷�Bm�Lħ���{1g7bmZ8�I m�mŌ�٧f�m��v�s�����c1m��ŵ��!�۝mbca�l��-�1�3��f�Z�IȜ{`�{h��9��׶�^�D��g^vsF�f��sbs-%���i�����n�I�,�0���Z�Y�HtN۬S-yڼ�|&�L��c+�k��H ����c 2{ݚ}��ވ5eL���!���pv��V�O�~r�4I��=��D������#j�$�_>�!Gy�\��l��������wTu�]Y1�{ط-e[�$��~9}�h<t׽�G"Ξξ�6ެE��: �;��휖�<�5t�y���w�Ξ����R�����(D%
��Gf��2	%C�g�I'���2hVe�CΞ8g-���K=���^ҝ�WJ䴒7��oCq�����Q�$�Ɲ���R�f�$�\W��h���Zx-b�[����Me,M����L�0��k A���X�	'k�
��2G(��w[�A!�]�\@kw$��Ie���w��v2�wD��3�Q&��>��3D��5⻞2I$���x7�cs8��a���sJ��\��4�X���5)�����%>�!�Ө��oaeX�t�v��:�a�e]���;�R޾��H�ڲ�����oO� d�ri��8�q�%��Us�mH�yʆ���T{6����&�?x���I$ё���}'�]mf���;��d	:���������n�Ƭpt��v���&�V�W��#=b�6��6^x8zk�~$�O��N�$�$ԏ�$&��z�y,��.���2Q&��~�p�"� Ȳz�2߲"#��C�/�t;�f��w�2MQ'�#�I_B	(ǋ�}�ֹ5����;���i$xk����b��*�4H��7^�v��S�.uQ&�#�y��$�F)ތJ^Z�[u�\���a��>�h޲dռl +Vy �j)ޒ|I�O�/��Ѹw]���n'��f� ����X;	,������� ��q+��=(�:�� ���y�H�.���clE��c�v�W���6Q~��d(�z^틕���%Ў�a�L��X��V�ٷR�����G����?,X�Ȃ��u7��z���Ϙ򂄈+�Zڌr���/���3�.m��۴�<ث�����
.�<���XL��e�om����&�m8;Z�.͝�A��+:����u��̥�y���+������΄��n��dܜ�&Z�s.��]�i�nyJq]�Vb�:4��[cs�ǎc�0���=����zv�]�lc��n���;vpv_��F8�+SrV�!���1���2���lX=c�����r��L[�m�7]~������YW�\kY����]󹽀 %g�ٍ�v��a�w��۫ ��X�,�uΒ���l���$=�M7���]9������]����=��X0��n�WOowUD�s�J�D��ƈ��s{�s`Ӟ�\> ���g���W�o�'D�Iܝ�T G/��Ł�)�etVK	 ck٬׵���br�Ϭ��L]#bQ$�;�i�$�6���`/��-��Dz1o<̊�V��	D�2��J�q}��d�2����1���n٫�Z���&�u쐓D�w�hI���i�6�K�@]�j�ް%��,����i:��[)R�ƹ�Ps�q�+�8ݳ3f����Qu���Dk��w����7���+�@ ���� 󏺼\�yzú;'I!��u�Mn��`U��Y$���,罙��y���q$��qL�|�ڕ�u�K1�l�i֣��'��h�m�n���BU㬳e,��5o+wkx�X|(��5��;�d���.�V�v�BI4I�^�[�j��d���)����"�W������xQ#j�ce��Oo��^�;��@�^�"�'��}D�h��u�d����Ub wvD�J$L�7����\�߼���KΫ$��y��&�?���������aK���̟���]��H����`| n����������g'�<�vo^�� �	�^�i��緎���\���͵��7-�H��.�]�<7T�D7sd���=q��Z���k�zo���-M��r����1+�6�y4OĚ�ME��'��=�κOx�k�����\�\Ho5&XX���O��T /n/�����gZ�c4H�[�I4b���P�D��7n�ὼ��S���&&fT�ϐVh���@�k��o��.�SҮb{Z�nC�.�P��ꊭY�/ő�ȍ�����9�u���.ef�+�w��Ud_�5�G%�6K�蔢��ut��4^`��� {�o�2@&.�IP�wǺ���eQ1|=�gy#�߷�93 h?D�4I��?j��HI$�U��~���}p[�g�@�|�\H��m#R��X��a�}�vHMIG}ξ�Y���3E�˟ �s�ˀ ��s���5=�����'<hWQ���}U�����Ć7b:Mu��;W�s\=`��c���m�m~�>�W�QP����f�� 7{����  ҿ{���c��,�h�j�N�{��d�̴�7SjJ6�q�����hٜN[[�f��k�Mfot�BH���$��:{ �rwj�sW�t�X�`Yb"4���6ۧ��%p"ͼ��C=��|I$���~$#�u��2àL��ʙ��
��Rvo)�%�� =��f=�>@j{���ٯ{/{��/A������9�a����ժ�hK�6���W.��35��\;+D9�F>�jd�Gw.���"K;=������O����0.�۫��4w�|���d��DH���)s��̸|8-�����Kfwx�׾�I�'�IW�րd��{� }��;��\�o�n��7WA��\�ư3��x�Hع�n,��Py���d%W�߻a��ڑm��w�ol> 4s��p@ 6k���$�8'�c��ޢo�������vb�^�~�+�,�nŖǄQ�D
fV��>��>�I$�T�{���$�0/yc$���Ql̈́�}�� N��EI"A"eA&�5��W���{X���]lױf�:s����I!��$�
�� �D��f�@��Df��ݒ��-z������l�p��g�O��[�2O�r�AwZT��O��+uQ!�N���@Y��˻�Us���f� ����$��%�gf: C��J$�'J�<�'/s�
�!ug	<Z˙��#��j���MP��W��F�:�բ�uY#��+�~��Θ���vo-ص=h	y|X/����~��t�ױ�=��I7]�;�Em�Lc�n7;�kc�×n.��pQ�A�<�v��ˉ�YOT�{����98�a�N6�X��'�۳�Wl=v�`Fᝂvֺ��q���K{Hs���umƞwK��v{+��\蹑�V^V�i-]lU͓��=n32:�,���l�lBGy��}������2�k��	�Ӹ�<vG�vN9��G�$�i��c�wìq�|5��5f�n�+v��lQ��<�v3t=<wdEe�����}�ݗ��WW�<��g�I>y`d�9{���nnOn�n*�&�nS Zs�x�'���8ԨvVԋO������w͐a��w~Į ؼ^�.��u��{{.V9^�~V�[��^�v�a�������y�` �����W��^u�������tI�9{�����M�(���a��Sy�x�qkH ]绬Kg��w{� d�=!6Nk{;���"��BQ&�&�tI^J͆h�r�(�譝�T �g�α�~n[����Ũ�I4I�9{��$�~�L�d��=�;[tq�������]�ޞDf�k�Y7�<��I+Y�,�k߽��~�9V�'�]{�;�Ĵ ���6� 2{}m�HI�Yt�lI��I&�r�L{��ީD�KTR� ���k>�򔸍p������s��o�{�`koG���ξ�O����'�G��V9�{���J|�D`�}B�.kN�����K<j�"I|���I'����2	;Q?C���,opS���,U���U�0<�G�B��w�h 3Ʋ/x�|����$��[���Hg��C�G��4r�e>G�v��>'��{  Y=��ϐ�{�JƸ�};�P�}����wM��pj|ܔm�?�e�<g�$�0/y4j��Oq���l��Q&��u�A'B��2Uqs�x��������ƥT;]Q��]��˨99:+Z68&�N���G�#�XZ����~EN�Q�5��w��@ޏw�X���猓������Q�k�*I�vf�8޸ۄ�Y$���c罘� ���v�kE��"����	��TJ=�i� 5�eo��̎�k���~[���(�6�j���=�b� y��7�_��ʁ����OZ�5�Ơ��ս��Y��1i<Αe��ұ[U��`���u�#93:������6']�]�~h��|�W���:cZ����j{��� �{.|{=;�T5(2,؎x�g�|E��"=qo��`��Ě$L���ޑ슘R�=�`.�>I��P��|p�7�&�$���ؕ���,7+��o�A�X�@}�]�\@ ����ǻ�z�Z��՗ق��*O��JFL��4�F��le�	:ə@�=X���5�aӳ���b!Ĝ�m�^3��p���k>� >&g{����j�<�B�>�s�wy�2�ɋ�^�\���j��*vZ���}�O=�y�t���[*)X�$�+��$�h��t��KM:o^e�N�:��s'~��x޸ۄ$���b1���� ם�o` {�������8���r��#zﻼz{�Pdm��E���>����`�cc�yx~$���'H��/wH$�~�Y���^������rv�b/��f�[�S�WFVtуn��;�Տy��Q���0K�Gsrpm�������/)s����w��=;�T;/̏M����6 w��T�-�ڄؚ��D����~�}���@��f%�c�p�Nq������C�n��u��i9�\�}ٻ��r"��^n���ӊ�����OV�
�?#�{���L]�rH_���4g�R�򀩞̸��y��l=���q$� �%��x�;�/G��Ã<�"h�I�˷�|I���{���4L
�X%���]�޸�׳P��+-���y��� �G�ܸ| ���{҂�o���l9�s��� ���vb�[��!B�eco��ywb��/�Io�\��I�����?Q:��	أD���E�����o��;�Q5���H<|��4I'�w,[�'��>a�^K�cxI	Z��Tp$�'9Zo�B��@�$���$ I���%$�	/�H@���B��@�$��	!K��I_�H@���B���$��$ ID	!J�	!K��$��	!K��$�Є��%��I_�	!K$�	/�1AY&SY�'�l��_�rYc��=�ݐ?���a�`   @      � �    @        4� �
�  IEPR�@��T�@Q@����%@((  ���
E o�J
QJ�
$JTUJH���� �(*J�DJ( D*@@"0 � �IH�� s�J��r�ٗ �{�Oe�:�5��$^=#��Q�7-R��	�Ǆ^�T�=������ N^֮̓� �T��R]��LN�:{b�Eoc�\:��q�zi;�����:<�UG  R�� ��*��@ ���n�
��:��y���ǓPt���S��*Y�{5.cP�}����QB�� z�@�� ����s\�B���}=�A�΂��+�@� �@�v@w`9�5(
*�O  ��!@�)R*A< dz �҅]�Af4/n��)Wl��S��l�ZD[ۂ#���r�U4ǔ � w��T}g{�*�x��T�G��^�t*n���5H�tMҪ�ǯ*w��ɫ�+���U(�'� �I((D$*��D����+�������D���Vl������fUɺw����{�⽠  |  n���zn�Iu�E����a'F�n��� q(�owW}�צ�O������^�{ h�:u>����*������E
�(�` �=$�������QC��a�O�Q���͠=�B��;��Z�T��}�>W{w�����u'���w�G��w���wE�IAG� ���rȎo��o[g�UyerչΑ�˪��x�����K��
�w�aOgs'��   0��h
RTh�F@� �  O�Ĕ�Tр0     D�2�Pҩ�PdѦM!�M  Od��*� F   LF �T�Q���U @     $�I��Q44#j��*f�hM3MO�����?o￿��X��^���;����� $����ꄒHI��%	4 B@?9	 �C!?�I$���#��������?�gi"����$��	P��# I!�I`�A�(O $���?M��γ��?�����.�	$$���ε/��u?���O��;4)DQ��F�_����SqqJj�]��̅8�4VZ��p����.ƚl��˙^p)`�N�����J�d����0d��g�M�T�c���ǯ�>�ޘ����h��=�fZRӸM�P�܎����׮��r�aY2l�]��M��g���]����4�R�j�����ylQ��oCȮ>�ozƱ�{�Z�;������5\ <�)ݰ��H�Q�������f�t�a-S*�\����mLW�`u���'ˊ4��y�������f�pȅ���m�Ub�$�6��a֖t��K��ȁ����wJvk�^�3G�-�`+ś��Ꮓ�i���A�	�l9�����%Ud?wo���.��ݸ����ۣ*Ǜ��d�ja4r��t��헕�D�n�XAG1�Q��wū@
?��	ǐ������X�یw,Z�<ے�ž���g9��+����k��Q�q�N�7F���(�<�wg\�k���C��vt�$�����j�ݽ�:�$�v��[�D�z�1�n�	���+�q=��[��h9֡țz`��m'��+5�5�61�;2�7�sw��m�1L����l�d�r*3.����nEB�)��5���!�)瓍�-̈́�-��Ne�=
���N�X��;��-f�8�.��`͑rJgV�[֎�iTXH���t�pF#����>\�0��;��ʛ`�A���[q[�n�Բ"�t§F���"��S�`�f%�̼�r��c�G\(��ԑf�JFl���n�PWMk���.\�fšWS�)���N=U׀A�Q�V��������t�ȹɁ��-L���+��Ib���$�DJo��M��΅v<
�G6v�#�2ܩ���iQ��;,�ݝ�L��.��8�����q�܂��M�7�q+5mz	4=ّ�����v�v�ݹ/m$�7�]Fi����ʢ��w>���;!�6.&����O�����:�X�dM���ₘ;��Z����*W�z��Y�.����	u#,���4�bB�of��_Kzp»v�崃��;u]/�u4BR�eK��jsוԟ���Sq���G�V嘆j���|��egs����yY�oźA����wo.0��W]��;,�s�Һ(�q��F/|+W-|:�V�*{��¦�|�Ŵ��pcB>��k��ލ�'���!�tT��d�-[��w���[ӱ	��c�W��/��L��쑥��7�����~@>���B�n����wo\�Q{�tU����s���"��7 ��r
zd�h��s
�x��ѓ:!Lwb��}ږ$��(�Dj�Wf��}T��vc����b)��w�J��+�����;HxI�p���s~��D������O��z�=1���b��1��;�b�Z�ܕ�զ��No������J�{�oS�d�������`2��l�4�ƕ��ְ�˹گ<�*E�TCDӤ!��f�A��:�}.���Mt�­���z�F���vt������`�� �%k���^0,�7�Z���+�S���U�6��j�H�����k\�L�L�$זY�wLS;��3�졾��9򺷏|.	l#��1F�s}���ʓ5��B�3g_ ����&��#�j�d�r��!��֓���G&wi��0GE�z��d�S�\�m$I�������p�\�nYǄgN��h�0S�0�pr�7Wb,7Q�	0E�ޣt�8;��w{�r�wp��y/��Ջ��v�����cӜ+������B|���.Ha�N�n���-����/��C(,LށV1��(��Ȱ�v�}7�Ԥ/Z�Á�֑��b����n/�7%�+[5`���7/�,�d���:�����в��yv�E3��,�b��S_Zԋ{�B=hc4�5�9^}���=G�i4���WF;in��Zc�u�m��Ȗ�(ihj�x�)��:��m%��P�̗v-�:��a���dxu�Jf�4���!Ni��ӝҎ�K�P�u�z�\�8NЀ5��+d�v�[��u�K[�A���u$�-�/�K����P�w�wD����J�p)݅�R��+O�n*�h�TL:
���4ɏ:\O�:�wu9DV̛U�}r��wFni͂��р���v]�%7�K9n��5Z��44R:��'�t�F/�^�ٛ:
��p����ۃ�y�t94��������d�v�F�;��ۇmI!�$�VW�k��b�nQ�wJ��9['\���I+�	ƨ�)���I0����P����5�x��gɆD�3 ��rH;�v]�� �R�c���5^�*�İc��:o<|�5d�x���;+C E9��!�k�XV,�8r9��|��u��&��CSu.��*v��`�t��<��Q�j[�m�pӃTz���V�v������±3�����h^G�I	�d�D�bSws4�1�ΑrYfs� ����Y���ۖ>�Y�P�f��7&i
0�� Hd�)׼�q���\��4�]c}�p��	ϖ�P�,���ʻ �.�ݓ��2'����8K��7�Ԃ:(c��׶r��޳7m/�t�n��C��6�&CQ�j:�K�
�+���r���+H�q��O9�{����Ϋ�\�_>��(�B��#9d���Û�D���<ۃ6X���yK������39ݡ�Yw�4z���Ӝ����;�8�8��\q�,����ڞ�ǈ���E3oY1t,܄t׼9�ɽ�����Փ��]�n�N�h���3��OPx�wr�D�uS\��)��J#v��^�DYP�5�%��%���k׼�B�b��s���L;�4;�鹦D:AJ��d�u����q
 (��]��e�H��ϳ;8�<���H����t^8�H7t����ѵ�H��j�=�0w�e�y=![z.B���<F��\�`
v�﹖x��:���n����{6 7�B�*�����R���y������l���z tѬ���݇�3��nv^�rY��n:�VA~U��z�!�N��aF7��4���sE���n����ђiU�k��y�ƣ�LqD87�M�rm��c4�چv�%c�7��vVd�$�����CnF�37�tv]X�Y�C)����%�ݯ����(طu�2��eyMe=�c�iS�9`ǩ#�:��2j��%��l��@���;�����7��
���\�a� ��H�ܢ��-�ƺ��3�M�i%�q�Ac��'��eA��=N
��=��U*���v\��]pd�k֐�b��$L�pdQ�8PӼ%���> �'t�8�lj����/`t%;Vܻ���֫t�\�^��f��E������'{�֖���l��ǩN�w;Xc{&������N[�{�p�]ۃs�is��v^a��a4sO7��*4oa� I����bE�SyyK��,4l?NӐ/���f��޷Z�\����p�q�	��M�*�n����C"�IH+{z���&����h#{z˜9=,la8#��s]���[&/�����.�A�qJe�U�:4fB�'rnV`�g�Xp�2!D>睷j]�wSK��c�	�����w��������#���iˆ�ݨk��i�ǉ�B�lx]G�� I=�lO���`��⸌���Dm�z��✱�+7���8g4�[�^-[�Át��#��8ޏsqc�]E�����m��m�`B���AL���v�B:�ۡ�
-9:^�6��i����uhG{y*l��U�8�+ݠ�a�Ea��aq�'����@�h����'	��>�T�u"#+@eI,���Ċc�eꋸ�����\d:��L�u�]�g^�,��*wq'8��a -a!L��L�
�Ь���&1:��u<@�qŔu�p�L��F�JjX2
�W8aś*㲂���Y;=٩Xs�ݰqίw������sGsS7\+T�󮞗���;Nl�Æ�X��\�b��|�9�ܽq;ȫ��U�����E�x'Y����p
�gP�9�v9]oi���)����s]�%���w`��2m��幵EI �ï���қ�8�U��bG�H;8��e��k�'C޸��p��N`؍�N�ܽm�L�uk��6���\#�;;P�Z�lz.ٜ��`�sj��^����}�$9���:u���_	�p|jk�׺q׌�<9�:A�#�oH.'mW{6Y�Bmѵ�ͣ�颵�bmi;��k��×��h畖F����uZo3��ìӸ/f��l��LNVP��x����r�ޮ�ۖ�9�L��Qz�XT�=��������2��v.���ۚ�e�&�s�:�Wm#hB���<p��2f�z=<R��-���;�Q���%q�E�q�s�5�lP��
�A{; V���ҙ���b�^�|1	 �R���N�������U�c<��9Pv 6�a�������Ӹ3RI�΋X�7u��b��������G�G4!���2��ϫ�x�G�1ͪ��R�,�,W,�����8� -�<ZW��:�x<=��8�M��F�q�&G-��9)��b%7�'��M��N
L�p��1/T��}���i��ǡrk�%f�F�F��)�.&H`�b��˺�t�`��ǋf��n�g��3����Μ�Aw��SO�:s.B��{NEX�g`-��RF+��|�o�n]Z�����${�Q�F�Ʉn�j�֭�G[�����@�����\��Wt`)�����S	������=�)���z�����.[:�F6��^��G=����d���s����w3����Xǀ��V�ʯ�ӛ���I>�Ya9�f�cΔj�o[f�yƈ��]ӳy�#�
`�v\�^�Yy/v�S��3aF��C�r�M+_!������^=�mӃ��dv[�8nEټto]kYEk|VJ�9ɍ�5�����䲘gf��%�ݫ5<�\�h��N�Cw�ɫ!�^=��F�w��h%�HX�MEZ���G�Tܓ<{/=M�c�k��_�ί�xD�ܣc^���y�wU��V�
�+�0C3Q
"����}�?�?h����SbD���w��>��~8vt~F���$P�)� PHC��	Y	 ,� � �B(�!"�B�$"�"��P� ����Y!*$��YH�B�HE�H,��P�a$"�,���BE	$�P	%HH�I�E	��@�$`$ �`E	"��!R@P��@+ *H � ,��a!��RH�	++"� )"�H�$	 �"� 
I� �HB�$%B�$�� + , ������'���៻��]p�$�BH>�=�{��C��@��x@zd	$�������~{5������8o[����|w�㈡�{|)��B�Y�e,\�}�����\��R&������XvU�0��P�F4��KO�u�3�-��u�{_���z)���9�A�����򐭤M�;��A�@6�h�6��-nsч�q���%���vP�c���ӫ!��q]վw�қ3sпn��Z�W_^��6���T�	�1�	�5�[!]�1�;Ԓކe�5��X���#N*�vbu�޹kh��^ozog�-�^����>����_��D���pCqq4i�;��#4&کk�]�o9��>�n�<��Ӷ�������g����!��H��/�Ԙ�r,S�5��̮�J��%���o��*��R��`Y��O��PDJ缑�0=��Z��ؼ���������}s�؞{�����hNO�Jh�����wf�;�����'(�wz�m�
�����$t��pK/y�5Wŝ�
��ė�т�G��*�P���eYJ{�LȬ�'������������.L,�❦�#U�1'�����R�V�^���8�_���7����V��9��m�q�;�f-9�������f{�K����rO�2{��\׾v��/{4��x�H�g�^�ݽ���_sD^�<��B�� ���>~�,����r3�x�^Ea�|7g����
fu�v�rk�/O�f�m�
ǀn'�csgwUpϴ��Y���SjA�1�.&�Ot�~�.J���y�]���m}��>d�.�T7�Q�y�'��Ȋ��s�{���{"��3S�٭Hמ孚�,8��^7��F���8?.���Z7��b�nΣOoY= �}����:Fi��[�ã��Q=&�Q�W<y����M	�{���j<Ylּ�.��)�cF֜����Z���e�E���j/�������}�w�����u`��Z��Y����/��_�0Oj��~�)���{�n���̹�{Jn�&.�<_�{K���_o���Mp��L��]%��{�Ś�B/Kobd�Qn���\��:�N�o�蟼���WϺ�9�e31��^hu�:�{�w]�n�U��@��#Y���<{���/S~�|�y��Z	w����� ]#���	��=�[a�}z����x�K�o�wM�<�v��f�*4�Ǟ9�Ux�⾚����GS�@�u���f62�eU��3՛���z��~Ǩlj��^H�����������2x��f�'tõZ�y��=�`^� ץU}��M}�8ڰ��fǶ�2��[r�k�"��.1�&�����L$s��潿j���j�)[��A;�4Eh��AM�om�8Ũ�t�9:;ủmȗg{�C��7HJ&Q�x#��.ry�?a���y���M�`�B&2�oVFmc��5���Qgx����g���ٝ�ٽ���x��������-��M��;�EMG�Ȃx������0����*����~��>q.���o�q^v6=�w�'c��A'ʳ�:_l��@�ݫپ\[�x-o�ޓk�ilOM�5�wKhF�B���5�&�����B+�~o�cP�\`�}DŻ����s�����ݨ%Q�:/�7(���W��	���{���8=�h98�Mc|9gPf��;ދw4�.q��}�PT�,s��O��>Ǹ���}�`��}�{Xȝ�v�Tf&p�X�Q����kj�ڊcC'�o!���|�4lY;���{���Ϻs���δ��;.�x�:�J��_1�/x��b���n��DfL�E�=���Q���(��on���Ō���r�4�m�:�=	��U+��լ��+��O�fT��!��5�I����e���Gf��>��c�)u��xZ)�{�z�6N�3q�'t����U��6+,�T�5' :̬wA��qtn涞��o�ۤ�6j������ֽ@q[��p�k����a��(9�(xޯ�������Yk�`!��i�.�6={3�s������y��k� ���.^��3܇E���ܶc#�����g�rR7�����r9ޘA��p~��c���pq��g��g���><�ۯfx=qU�����lQ�8}4��tރy��9�֯>�����@k�8�W�Dq �~[�袖���a��0����U��!������W��kڴ�U@���Y�o�Z�Gs�z�	�N
̀�,d:���7��\؝��MƇ��"m�*k�F�3��L;c=.�j��m�$5�dQh��ͽ��[����Um+%�ٝKn�=vk�}�٥���K�9���b	1@_��`>���R�^w�s�vK/��a�� &�����H��H$�rF�C���.)�#>��U��Tkً%D�=%^�R��ŎE]��bY����^Ζ_
gq^�}Z}y3sWS��Ȇ��Ln�U�f��TΚ�ɨ��:s��r?[Y��w^g���y�%��=n
s�/������K�lSsi?w׬��}��=� ֏ye|p��}�2ܱ7!��dԤE�9In�U?O�XF,eb�P���{l}b<�r�`�{5���x�� ��2�\�51�E��b=�{�� 9S�N�@�݁��Ih�L���=N��v���V]������}���.�{�����X��'�����6�|+Rjٳ�qCy2��z���^i�7�l6���m�366�����~�3���L}4�D��5�;��;��DU���#>�o�ޙ�yS��O�������w�}�T{���3p���\�`��3��Bm�-���;xB�#��9s�ʡ>��V��xzᏁ>�`���nnn�*�?��ݗ�]�Ĺ>�&y�я�n�����/Ǿ���Uh��nu�^4.۱��l����ζ��2(�Q+qe�\�;��A���5����}4NE����e�7��{�S�{���9s�WoT'��0�R��?V0�ꃥX��n�\՟V���,����nX�����|r�sϮr��ggj����ɗ�O���Sf�n����K'����bŹ\Xd¦�.�0'�746���wV��@ѨǇK�ǚ����5*�E�L�1��y,j����/(�gM^�J�����z�o;��x���/��-�#7뽳��fy��n��R��8�3r�x+۸�˄��n��#���S8>�<�X�oX��V��oH��~��_]�3�He���E�,ՊQ�.�3�f���]6��.�=Qm�[��;dEm�'i9nu'��ti��� ��=g�.�ל����	�)8�V\�#6٤2F6�	R�l��S>Ք-��'��8eq.��yM��O� �瘀\��ݗ�=�~��Xi��p�d����j�"|���yJ�/p�Pɷ���۱hXqM�,����h)�Q�s��9p�B�/m�t��>�yv�D}���.�d={؞�]=�7�j�=����b��Ə"�x��<;x�����!������yet�g������w�"W��N�:�i#6��f�m�;��~�1S�vz�^��2�L�1t�<�ɰ�y���,�i��־��6�}d��;rH�.h�Ðɻ |A~�ֹ�=��@:�/fp�ս�#ɠ]�r��j{��G��I���n^��N�TέU1
w7tl�1X�_W:�M�j�5����'��7�f�c�"=��/A���������ݼ��<6����Ua�m��sJ����/iY�wM|U"��@�pl�����{���{sƗ�w��(3�1���'f����a+)�r!�cӔ�D!V�.Q�4�[��E�A;g>>�۞������p�1]��{�9�cYt���J�~�&��}�p�����0w�Yݛ:*�;d��$�z��{�蟀{�n{*���4-݆]�U�'zH�$U��wO=�Oy�j;�ol�%�ӥu�Uӯ,�{�^��9mP��⡜X��;�Zw�~ͣ7�T���2;�\|�����3��+v�i���w�8�\А�P�TC��)����N�	D/U�<��fx�C��O��*�Y;6�/�����qK�l�F�
�U���'=��Hy���)���N��^ĔL"�
�|��YW��'�������]�g{u����1��"X�����=�wwbQ��i�×�#����";۝���}�wu"��� z���:0v�)n[��An����^��i~@k�7X�'�;Z�{��� %���BC��z�iDgl���y��A��Y�x��z��-��Ǹ�T��E��ȏ]�4|�ǝOCO{n�Ŝ�����b������x�}gy.�t��{H�L�&�#�<�[:����Jչ|xo?�	�ZA� �RRG1E�B&5�q��n�һ)�G�3-����SP���T��l=;v��y7��I�����I�#�=��]�_g��Q,~�=�ٺ��f�;Q��Z�Enk;�{b��#�j��^�����������bъ�gal�6Si�qN�r�V��Ň��f#�T��j��S��z ��љ������P�5J�x�{=�>���Œ��р�7g,���t6�8.���n��uw�Q�o���3�����M�g�x�]�^]H*����=����x����=y=s�G�E{+�H�Y�6x�J���s����{�7�S�����>���z<�>�m���̀��� 6!�D��B���nC�c��u�;��wP҆�K(�Ă�fe����yK�ݓ~&�g�f�����?E������3S�}��y
D�z��U���A6�{��Q5/_x�9��g/��5��KA�S{s�y��e��U�b'��_K� .��J��̶s�㫳� Rs��/raܭ,S����� [7{�j����sꞡ[5l�aܬS���˶��
�XgVim+X�X�����/n"%��hy��Nn���K��z��2�.k��!J�"��}��dJx6��}/`�篒�f(���f�S�@��;��pe�'n�JFT�F9y��f���5�oSz�v��Est�5A��_�Ns���N^�<�Ӄ"�~N��)�9�=�{{�V��&��q��E�B���$����ѢkM�\���0�=�oBs֓5q�������jݶ�|�>��<����+�x}w���3����힣4)����_Ob��`�re��L��|����,��XY7���!��w�Z�t���VK}�q>�7}��d��{�D�b�2���zw{jɧg=�ot��t�.ˁ�yJ�G/�z��o��Hмg?"��"4��ʵ	,��>�~�_n���)�d��or�9����x�z��2�j���1�w�o���:�q�w�|F?]M��:V�b��x"-5?~xx{��+"���v�"����,�3�ׇٶ��\���`tе�ܰ$�=u%��]lj�����k����x�=v��Mz8�7d�v��v�s����+�茛T&�\CF��lZa΃�1)0}{e�H;ChcjNf�2���],-��Wal�(�fcj���G@j���ZU�ː7&�n�NG]^U3 X���jT��8h��bς��4!��7Gd�=�g\�:��=������E��9��ݶ�n©�	�\͸3��Od3Z|E֣�mI�=6��lrwY6�O&�6�}�����+t3f��nb+gL�e�G7U���Hp�[k���݊��GWO'Pn'���3��:��ta�p����V�,[)��-;��1��K�����m���4T�2�i�4����=� ���٧��º�ch�f;q]�æ���\������#.ά���@Wc�q��ݴ�>���j�qxVn��7�o-�\���;�8��:rqӮm6P�J�֛������D2�'lX=rp"�\�1����;$��"�o����;�hWiYw.ٌA`��!�m潱��m��c�d��0X�Ku^Z�&GY��b�%;O�^I�M�n.����ic)a`�ڂ)t6��m=nr����A�[��'y��9z.��=��k����F�=Թݵ���4���k�$�r��L�"��T�I��Ejr��T4�]�s8Ӯ:�X.�[]0�;�u�{c�c\rz�x���zvՎNz��o��]�����k��N'�<d�-tn%�%S����öȅ %֎6fwj����а�%�������ָwGgcP��քxz�`s&��c�'N���Ƙ�6�5�y$��ذ�6�j7����VذY�֖���3 
Aʚ�q��v}�+դ;/74m��!�!ώ.���kݹי�{n�e�<��W,�N�6��Ee+<�M�c*	��ĭu�29Ȣ��+�J,�$M��K�6cn3HB[��[2B�x+�a.m&���uX[#oj���#TS/Oo%LcBi���5��p �)�-۫9<��8�<];C4n�9L�R�G*�a�:4�n�=�9K���>��.���XC1�5����vU(��]���	���ca�M)���.���,<gPq���eu$�uj�]��A,�JA#i���mqZڥ�6�W�`���1q�)��b�g�-]�Q��<�\�e�t��Z�;0�i�Ś�r2�B�; n*��"��b%��kc��س�ӕ�㦺C	��q�Z�!iBF�Y��LL���HA��])lҹ��<e�c�f�v��,(V�5��7h�9q�D% ��.h'Vy���O&�n��,4^ɸ�:�枮1�c�{$���Yx����o�V��Ʊx��k���kc�/^�L�W���/:��K��x�0�b�Q�8����ZQ㲀����4Â
��rĖe�7h�lM���d΄��^K�y���(�s�����)����׆����S�I�iHbݤ��ҕ�.�F�ˊ�LR*gZF�.��Fj�,cKa2-�a��]5�8Me,��vw=�7�q�+tf\<����b�n�#k	��bh�ȡ)�5�t!�2<vո[x;h3g�U�qs^..����s�^-��_6#�����O9��g���n{9�x�m��wY�Z8��<��v�/d�I����b�x��2�f�M]a(7�g�x�0�`��z���C�<g�i�җ]����g����q�xe{��c�8;O��us�p��q��$�.\�R��2���F�^#�ؒ/t� `Zzx����\���]�јƯ]���y�t�e"�t�j���5�|�ǞT�,a��\�z��<��#ۛy7� L�67w Y���x��i�f�ϧv��\�;�f	BvŎ&���]�jh�����&�.�[�%��\]̅ʸ�U�pݸ{fL:X���A73����1Q�̡�i��$GV�X�=��9��;��c���ۓ�g�(m��ոˮ\�&=��#��`.��+4�m�8G���u��	���<u�|���T[��{)�
z5tu�����*���v���m\���1[t��ź;V�:�ݧJ��)�k�i�yz��3�3C�<��@��Kstf�ʼsM��vj��v�|��#��m:j.�u.R1� Ia��r\56�fc0�K�����s�ta�-0m�\�0���(̡q�G\�ю�ֺ�Uñ���uJj�7�]�Fy��67+�B�r�l�ƕ%�:�V����a,Z�&!���[�#��)n���G��캘��8j(^ݯ<xj��7�ghѝ�����o��s�����oW<�Vn޳���6x�(Ru�� ]���<��y���k�|v1����i�gt��֙r�bn�E`���t�]<:6����c!�jwJ��#���:y5h�kj����e�M.�6������ஈ̖;@���5e0�VXP��g��y�2��tj�=��u�i�3��4l��m&fs�`�n�q�}^���Xwc�mp^�-P��6%�j97�i9p��!��u��ۏoU���,���p;��Z�a�;Z�On����%n�Zƺ��j{���t�L�c�ƃ�#x��t�`���A*Z%���9fI�����]{;8���ց�ݶ�7	��+���ۮ��6J�*��i�����v��X1O\��g#�&X��Ar�
�n�uN+���M"�F�s�'�WgU��7=k,b,�//!a�f��0[awOn�&���q��É�����8�u�PvF!K�T{W2c�v�&���ۓ\ha2�#`�\��v{I�����62:�'I��ź�����R�:�GaM���m�,H��J��eѴ��N���x��)u.��a����IcK6�T
��x�լM���Q�s�3���]�<��Zm
Ev����a	���β��ԗ���ӕ�A�!�:�e�9����:|���>ŋ0��z����WA�Y�e�qy�nD�C�a�G6�YY�ŗ6�B����XkL!me-�Y�]�f�����R�e�1��2EA\Z����m���k�Mv�:2�<pvwe���s��cy�h.�x8��R��JM�EƋ�[f.e���Ҩ9����:%<i'FGi;kv�����I�MJ��:��ʹ��2�8Yh�.�,#tu[��\Wl�X%�\n��8IL[W��r���Z����]��g�S���7Y��T�74[��;��Vy��ӛpY.���.���zg�q��9IzƧQ���AsO�ma���u�s��ӽ����4ۗ�v�2��^X��J�]h�R#u�ٱ�:�����2�`��0l=���l��{拎�y�r<�zv������<�-�Ս���4�&f��K
��\�6!�F�6ۚ�1�����k��K[���u��]�fܦ�;P�כ�Z���5Y�N�Y��Y:���XV�E=��\�����k�z<��w�*�b�;r���<v���ݮC���T(�\�z�<��'k����&���m���"�;V�k�Y�<>s�I׷F�'κ�p���@��g�D(��Q��� ˨i/1[1�e{ w7��t�,�1�-�voH�!˗.��vy�B�T�4ܦ�,8˥k"�%��k��2���<-�C�+�pc[)�)Km�u�S����������iM��u�:�p��(�Bt-<�
/ϰ�_`�ww�?��U���EUUA��+,Q�TDb"�(�PQB����X��Eb�#�@�
*,X",�TEX��D#1"*�U"�Ub** ���*�(�*�`�X��QR1��X�P�*�ȋAEX����U`����j��X(�UY�����AEb�,AX��lAPX��0���+QF�UD,�"(,EX�J(# �Q�UF �D`���DdE��Qb�b(� ,R(�V"�	
@Y(�� N������ֱ˪�f]aMlfl-.A�f64#f.!��}�ݐ8�Q�H\nV1��=��D��\\�6F'�[K�fѶ:�ɧV ��pX)�������D�6��E�)°�s4����
A�q���s�8��0cy ���uM��D5�{hۮ��gC�Lq-s�-��Ͷ��w3ռF�ͬr
�w�X(0��˖S���h{x�����(�(K��Q�M�K`�G'.�`4�q�\�Z��%��74l���N:.�E���MvL34b:�R��Z,	Hpcn�5�]�t��ֽQ��m��o�3�@%����t�\��J��Bu�Ͳ°%���X9�q��n����������8݌6s�p�M��lX�6l�l��Y��iL1���6��یA�v��Es���[BuRެ4:��4�g�rM�M�=Iy�]EθiR�̚���)�)؁�6ך��������C������o���v-WAқ:��n�9�&4ͳ$��-����5q�63F	[]*�H����&��/�lgE�,��퉡k�3K�G;I�mV�2�ݠ@m�eE���q+K��cK4�:N�;t��4&�p�v.��C�Β3��Sҭ����붇��}4j6 �&fs� ���q�A�ۆד�p&������ �v�P�W;���mA�b�`�ќH�E�[.3�5��a���2�u�"��0K��4.V�ř�v�s��mY$�/8x��3ky9'�5#�EX@��`��eB�EX��e�Qxr�[[	J�o�E�e�R�ȼ�XF#[h'/B�Z�X^�B%�my[kBǃce�e�*1�Tia���-$���1������i���� + �Ym�EKV�ե����%�?���r��Ai��
s�׌?Q�O�Nod�3�#��rR���tI㶃�5�py8sGK�R�[[�e��H8솄ݵH�!J2�=�^�y�V�$�`�4��g�ݓ� ��[mLj�}� �� 7�iP�/�3	��C��D�f�ɱAD��~#�jd=��kzfj)E����Z�}�A�Ɇ�P+6���Kxʺ�N�0GP���H+z\�U4*�k\I8N D! ����u�V�u|n$����&��
!��xGCj i�_A �^�Wt� �I�ju�	��}ju?L�t����i��
t5u���2gH�ki����aw�Mc�8�Oy��� 켙0�ڙ�a�f�5�k��S?P���&�3����W�"i�K����㟀/��Q��TS��� Gh8���˚F��T|�ڪ�&m�Y�ލG��� �kzdK��A(*j"�9��kG1��e*o�� ��c��";�f�A��6��7s$ǩ3u���#c�A7}2$˪.6g�Rn�� JI�"�%��.p�؟n΢���5溹�&�;80��7��$�t�N��$:H�ߨwu�d��̂|�M��a�."q�W7�Tr/(�Gf�RP������uTU�Wm��!�;�~�Q�A�v��j[�w�V&��é�ٶ��O�H�c��J�>.�{���TnnwI�a����Α�4Ό^�3n�;��A�f̉$])�ii����Ğ�������RU; H'N�~ ����x'!����r	��@P�P��(���_L���OR�6 ]:x	&�Jd�3��\;VV�Y2a.!������k�u��K�v��Ai�)����ִ�q��~�xz���:�u�zOf�WT�.:�DfX,��؛�[=>�
/b�e-�nZ�:��@��ѕ	{���]Ш�n=�ѹ�<�R屴���n8>��z�eM�[��H�ҙ ������UĦۙ���s���'7�%
��'����	�ʘ��d��O*�{�;o�u^F�&�S��0n!sE�'k`�;Y]ۜ�3��\��'鸾En_*�+{���zlc���˚H��tf�U�L�D�0�;�Z�^�c�qe}��	J)|�E
�u��u䋍v�K��\T]�lƮ��7��4D@0�P��(�"��� �oeO��Y&+����$wnȔk�B�ل�OC�&�Sq(+B;��$�z��@�n�A�[�8��A&�|�i��U�vdo��I'�;5A�煂�v�ݷT��b�.\6K�]�P��ڍ���x �}�� u���f�%H�=5�7���Aڬr&�Vn"
uEwd�&�Ix�r��<�zw/���P|��i�{�*}\�k�3ۓ9{MǅL)�kf����3=�[�y�g�rm�0kk�G�軳�� �μos���:��ы]�tf/ �WuI���;q�ݶ1v������]6.̄�l�TԀg1ܜݳ s��Se,O���D�؎�y�l=�3���tv١7�BȡMl��)�1�b"hL��mM4ml$�BZC��oa���欏H��k��3Q��U��#��v�Sf���<�ݷb6�]=I�qa֖\�	a�wϾx��Kn�s�׺��H^ͺ�顠���YX{��R���'��RD��������s;ލ{5������^血n�{pwv�P�;-B�I1�-�$�),A$W�{�Vg���7���/��w��]��7q�!�󪒡z(hB7o��\+��R0g�FeL�/$��8l�BGtY`�E���mPt�mH���2I5q%����&yu�]3U8'|b-�;s��:����݅�Dґ�F,��Y���Gw�~[���Y}$��$2���&0I�u/�:�Ht��%h$�8q%v̉ �M���k�A��B��kc�M9���/!u��.�y#���We�����m�pY/`l�Q����������Iz�'��l!j6l`��
!DE$��$�|�խͩ|��k"K�|wo��[j ��I��wSup���ZY
�d��H'��S���":,��k!&��b��OL�/��鱴�s�GDq��ĝ�n��0�zjA��r�L˂[I��v53���T�Ҍ8e(����9�p�&G
ز�$�n�|wm�QK"�o���84��t�b�$Cn��� }���[GLcT/ H=��v����~���>����z\HG �\�#�N��n�}��9X�8�eO._�B��S�C.^/���Uȫ�hG�x{�s����h��=���/j{�&h��gw�H'�)�H	�ЭB�P�N�DF����o��v����{�O�x^+N;0X97s(�Z�-��rr���K�B�m�s���F箨>�rB��^�����C-j\v-���7L�]	)4��نm̩]����p��%����,�T {��a౽L��b�D���H��7\7!1R�NY�K�$ˤO6�3z� �M�އ}0�7vJ��/5W!�
sH��B^E ��78��+��>����M9$�� �r��U_Fv�N��i�� ��$?�|�)�up����vt�v�sPy}�m���ؾ��]�WÜ/t\������Ã��\�=��<�Z�|H��F����t��d�Oe�}]T�w� �{j�#z(h �ΥP�[A�v+j�p�dDĒ�m0��^NVhL]�+tƲ���i�EB-��r�-��bToI$�%�B�:�{}Y4���vmRn���r�"ߢ14v'���}5J�< ��'���$�mh��Y��.A.��M��Fj�`��vD�AJ]�mȠk����q����
s���5�E�!����V�􎾩+4N8�al 	�LT�@O �\��R�#�n�{�qt႗:1��*BκQ�[!{����r�<�[�|=�{� �s7v_�)w����'����BB��.��MuDؼ���Gd"LD�f0�a;a��gWZ;v��U8�I0�[�x�[�~n��\z�6��6���9��^�Q�Ϩ�"°e��[��2m��,��H�YtJ���9&�"B��Ѧl٘���!�4��[��S�-Jܱ�I��맮�rݴk����.���i�cN�٢Ix ��Ӭ!�I�QS��2���IR�}�K}*���|&����/g]P�&'�J���Q��[e$�D[�c0��7S��)��(V>��U!vu�E���
/�/K;3q����C9>� �ީ��Qb�r�D^�����$���6��Ld��e��db��8/x{ո C�T|��D��F������%��j"i@N�ݵB�,[>�?����C�ڤ ����t���y15,�	%�(l���*�1,�Vm��[r� ��r�-���"|�9sȌʪA۷J���lb�zwg�iv�{2fA3��&L$�%�X:�&V�Q<�a�'���
�ӛ��_WSD�0w���]#)+f.�5�ֳ���#LaxgMY��	�{�Q�$��ĀN�Q��y �J��'в�B$�ID�n�H>=ʈ`��ww�bkJ}+�f�U ;�������R����&��ָ��;�N�Q`�7������ጭ�/"����!M�&F*ޛ>fft�k�=��k3fH�TX ��}2����-Ć�H���KX�Kp� �]u�n�n�g�ي�ce��%�r9��'�VvO��MZ��_uR8ݙY>&���Ay64	GN@���˚#_R�ޞ�����@ ܛ�u�WԄmF�D�W�o~
�jb!��v�gF���*��>���+�����|$f�n4T&��#j��9V�=p�9�q�:o��۞�����/2��+����O�G�w�~�#���xN�x{^!��\x�=�����>��0:�֨)@�²o��SZ��U{��@��h���@0�ͧ����N�8�@����|&��+�y��0�}_g�%��p�������r�����>ɺz[o��;�ؒ�6rLe�k�����xvo,9�h�#9e��}5)^�}�+���C�Ƀ�j�%a�<q��{�q�3�SV�����AGt8�S|�����/;�'n�p��5�ܸ��������e��=�>AWݧ�V$|�'%����la�g��؄�=H;7/�pF�n��I겦��1YH�ݺ����[�(�nT�8�������+Z`��Ŋ��t��pi+�B����5�|P�9�'?7�?5;�|��?��o���ZT��d�|&���.�z�/�������|�{Ҷ6't§)���>6���0��Z�2�G�ܪNΜ����ɩ�=���y�{r%L^�y3&u�_�£"�fi�r/ZfF��\��n�2F�{��K�F�@@$](�Wd�������b�E��v��%Y����р�Aa�@D#Y'�*���dQAbȢ�ER�)%�V((,R,A��aYĨ�F��q�����X��*J�`Vb�PYDH��E*\���U����"�-@�1��U��73
*�ZDAQ��Qb�RȥkEm���a���+�KT
�0X��Ej�R*cLBb`ɉ
[U��ԫ+AkY�UAťnd�1UA�e1YUł�X������PF"#2�� Y2�b�E�V�X(�f[p�*ޡ��_~"'|�!����H�5���Q o!:�y�qNltY	�A�9}�#�;>ǳ�GVM]��Ɓ~˼��o�-b���P���*�!�*s,S ��!{�P.���w�rU.$�'
 �-���U[��g�O[�p��[�iʇ/�q��dL�^�Q� ���_;;�ǹ�]�w��u�W�f:<�l�	��������`��+8	 �oO����Geư�����~W�'�.k�'�t�۶�|3�%�"���j�������Ƃ��P��t!F.<\wE�X�s^1'��� ���!��;��P����#;������c��jb/ ����h�s�j��_��qت1����;^VV�M2���
���; �"DD�����H>?�0`%U���^��ܓ�ݴĂuI;4"���Ϩ)�"d50K����2�v7B�n�k��$�n�NCD�k�v�RT F{���t�&���B��K$N�WV�OfL�"2N�*4'�Rd\��s����T��U tu���~�Q��{j�P9l�P���ڠ>,˄�6/�y������N���� 	��eĂ��WmR��p|ov��ye& ��#:\��=��":vD�Y�x��V+$w�g�35����]�̐}˩?I��M�΄ѢB��y�ᒻOu��Aj%˛����58�*�'$�����~c�0�o.�OL���<����{��y53-�r˪����v�Q�r��v�[��mɘd�l����۴s��<���+�t����ب6m��rX�h�����e��Iĝ��-v�v�K��]+Y��Hlƣ�0�ni�3i2�5-pZK"W�q"d�<\A�Ӯ�K5Ӛ���f��:���5�j��]��m��v��y�Lb�u�6��~z0�6��}��B�� ���rtoeG�v^�|Ѵ����
 �T{�̓����+."��^�F���$�v1&���N�~��,�M�d�OTb^w�� �8��Z�od�����wdɼr8"Რ'T�e�`��$ŦH#�������US�Nϲt��F�y���s_�Ԩv�%]=�NS��id�{7g�&��A�YKo5�M�7)W�u4��u:��q�J���CG��E�u��xy�Z�\�g�������UH��(�evB�e�D��*��
��j'�9���d�����q��j�6.�#bm�89􈟩����m|�v�cK�yJ��Α��0∬���j���I�}3�I����Fȵ��g���5���KL�W��T��oUW���xg: F���W�UDݚ�7-L�wC��T�o�{�Ҡ[�N��/	��a7�9}3\�`E�i@.F��H�VE�͒�+uE=:ff|I;�2$}�l��߯oQ�ꭧ̈�Ҳ����c5�Դy�,8���e;I(}Z�z4_�8��}>�ɑ$H�,��.��˷9�.dk�\��:HF�LI,"�a���g.����'�����A�60^��c�E�U[\� ��lY�TY>$��Q�ۓ��Ά���FU�V	ua��2]eܞʆ�����'�l��x�g���zO){��n7�Uu� �ުT�M��m��a���ʚ��ckT���@܊/���Z�]	�{�#|m��1�l@�
PБ�|�vl�/�$l��O�oj�>��>��]�-�x��<�O-���[�S(���V�����hǙp�B:��� �n�Q�"�,h�ڣ#�z�Ue*�\Qd�B��A~��.��&�6�tU� ��l`�㻶�#���?_������p@�(hwjfth��ޥ@�73j->����6&����*#�8��6�����i���������z�g�ߝ�~\dt��0j8�]���К��������Qu��j���n�ӳ��[� �3:�����O���%���=>���u3ܼ�1΂�:0��g�}.M�H����JK���L&�X v�:����l��-p�u#�����M���|z�KeٮH��rQ�YS��bØ��g^9���p�P�+z��{�"��"���A}NA>5�čH����Hg��4��S��ki��W��\] �ݥ_�uH�q��ZP���gL�Q&� t���v��.鳦!g��@����l�R�>C�]3�G�>;���7�'�Vo�� �sv���M��7Et����X�k)tU�F�å��eXU#p��Z�#��{�����T�9Ю0P>+��^�0� ���j�+��XE��؞�����ӹ��8�Q����>5�-�q�ܵ!ޜ��6Cv!�ջO>�玽�kd6ݧ��B�&v���#����D�]x�K5�4����j�/<`����4<U���DŲ�t
�:�IB�jǇ�n@�u����\^(�=��k�Z6�t5���@�ⁱe���eܳ��&���va�s*Wo߻�Д2Bb�Dk� ��\�$��Y��[�E�ENfzA�#/nd�'	p�J;�K"�N�b'TӠH$vȗ���`���Q�ju�IuCfi��޷ �V��I���љ�=����$�E�!�q$�C����1�����W����
�t���bh>ڢ�v�����3:&���y�5`d<%������>�V��V�ћ>�}|���	ٶ��֌���4�+lSCLj��jla(�o~}���O"����>ս�G3��*�L�=�$�����ܫB2�ą��C:�_]�/r��"v��U���������h�������(��#*Бv5�4�\�ˎ���~�,|g��d�����m�C#/��:O{K�GƼ^������/.�&�2����8��X�Q����v��u�NGn�|nb��5ɖd�-�t�0�z|����f��꘺�� ���{����U�q`��/�~ѣ��e�bR�!L�E���zZ닌tѝ�Ư��D�8�{�"4�A��bA#o�F�ݾ�w_���t���PH�äs{Td84��I�roo:vv�yl�q�.��߯aLK9���:�do{��;+H��[i�*N:5Α�%	#��JA�y���R�@⟖�/g�_�zQ=�yǗ�k,{�p��B°�/u������T����.�oF�V�XQ��Ov��#���'�Q�蘜��u��I��#z�F��{��"�,Y��D�#'�T��mP|�Y����"�Ad�)F6\&`�P޺J������pkt-�� �8m��o���%��4�X�{3$I#yQX�OeU�f��gH��ʤ
���' ��gF��7����(���"I��Q�GE�6vtd]�*�z�����* �M�Hp���������#r�A�d(�ą��A�1L��$�O�]&I�ܴ�8��(+�����K�h���F��z{(֔#7W(�����<��^]��gVѽ�}4 ��A�}º�d�<"�dq�B� �vȚ�����7^隹O,�ϧw��f�v��_O|��:¬`���Y�.�t��8�%�cj@��0���i�!�����G�2� ��R�Y%ez3��'��`�$,A�I~��NuUPJ�EfL�S���\0{��"B���&fOv��H�pK�� ���1´꼣�w�� ����P6`%�LtFd���c�J,��3{j�=����=|F:���L�yeZ0YQ	����{�3���Fd�5�	;��>��ro�痐;��!�5�������kr�.�h��C�\>��7�)��&�,TNɓ�����{�l�p�l\kG@�oڃkbI/0����m�j��<:�d�b���w6����W7݈�S�љ䦧��.h寊����q���LI����j#Ю��1�淎��˷���=}�8���2-�_&��.h��_�yܽ��샋�x�eѕ�ym�g�z���wܽ6��J�hvK��oG���g{pnAq�
!�t��~{��ye�����ȷ��=�e��V�)|�Z���`͝�9��]
�X����;���<*�VwW���-��H���m&z^��;��E�͛��#��z@w��ף>8}}�܇�q9X���U"�� gE����G��ً
s��*k�1���<�f,{y-�T��W����:i59q��h[�ve����D����k���;�M�#�c��A���-]m��]:�[��^�X���՗2Ij�޸U{�5�����	{^T19f�=��
��Z=��޷����O�Zx�.72���е$A���ĳ��K}'�?��wO,vl�{���|��c	�,B�f���
6�.�]r�dt�i�AjE�)V�a(ʭĢ�T3�T0k�e�X*�B��T��"�Z5��@�9EƸ��P�˘b�aX�$X(��C��µ�X-E%��T1
�b�"�Ɋ���m�2R�-"����25�PP�+0b�9DVLf �T��-X4�Z��Ee`V�ڨ�
�̒�1*LLL`"E\a[Z"Ţ
)���dD�T�dDY�X(���P+(��Z[(T�Ƹ�2�	����rʩ
$�+��-TP��R��k`�UY����*�Q1�����B�2�Y���j�K߷x��5�����tv�sD/Wl��8d��50�%�ۖY�q� �ZD��u���pr�;�ձڷ���%&���ĉtn�unQ�7i@����vg��a]<���p\8m��͍��hMC�[�n��`� �q�D\[X�jb;6�]
�m)7�h����˵�q�2�`�k
78��5�T��/)��{c��@nv�n��lV��tIte)���6C�\��X��K燶M4���Y���fd�l�,�C�v�X��1���&̈́�ke�nMc6��:�j}�K��v	t�fG�-�5%+XU i��ˬ��Q>����Mӹ��p��ێ�\<��k)_L��.��z��^ƻQ�ղ,Ǎ��jwY�6����+GL�l�[V���msp���[Q�!�.+%ɒ�)���m��\<��cr�]s�m�F8Ϟ��Bon��<�]�&!��r�Y�-l�#94��u�ۓ!Q����'��킗�ڳ��q��k�(m����1� vq=m������K[��x�8��n'������W�a-�k�3��ma�Ş�؍����M��>�wH�1/֝�^S���6G]�����	��j|�A��Y��Tn[Z�Ԗ���]�"5��FN.�8�v���=k�`CB�3c��D�����]���[�\�]�,oL�[q���6̺Os*s�*�i��Y�In�^�d�6i����b�׋Lti�xnRnǫ�m�e�:0��K��1٥Q��Ni
RnڊD�tn���Ix�ܮ�dcK�����R�x�֓ϰ/<+������s�8��k����6�(=:�������Kc�.4� W���6gp��潵u"�[�9|One�t[�"ʎ��&���쫅˵��u�k�)���ն�KbӪsk5��C�4ne׮��h�C+L��(N�a���p�2?�p� �޹�!�}��D<?v����>3�ם"o-_��\LH;Ւ|WS9�QT��� U]�� ��9��S7���ښ��!�(C�a�������r��m�\���Fvk	}�'�]�$U�8%�>��.��A���P��Tu����nq���$�w9]� ��i���D�}�P��Vl�kQ�t���2}>>��ҳϺ}����2��)�0[��kv�6�΍E��M�I�"o;���J"���zA ��L�I�\��y���_Rw�j�	�1LԒ�(g���nz��؍��z׵����݈��ȸ�[�l��A�����;�q�k��o�qN��l壴��K!���{�X�� ���$�Tۀ���oneGD��{#>�P9M�Ȏ�Be��@��oC��N�#7�}>=���BĞP����7�����^	@��U�>�C� �=���3g+D�DoL���$�9J#'�/=ԨF�֫aR�ή��:�+�Ԫ�%뽺�8���
�;�2�j�;q��qu2K`�]�9c����6����W5.#��P��r������u���٪x>7�X-{��8��j���Y�$�k�$�w?f3��:9���9Ks���Gs��7�_��0}��UuB�u`v�f��Z�^�w:��<u������������{�ձ��\LT���}���_~@����ﾟI��~<�,��vy�ջX�x�FF@d�H��O]�߄�tsX�1����#a���P`����a�>�q� ���$�6�I����TgB�T�M�yӴ��`�܁�=�,I8�u�_o���o��!|�D쿃�E�T =��vW�f��7)���T+�g��qK����*KΧ��:�U��$Hڼ��$��}"O�U���` +����,�R[��~���uP�i���^�ӳ�#�o��۾rJ�6"\(	�hH���8u�`A�[�T wgU |w\�ɞq�t,*ؐ��W�Z�(���3��f~�W�㏧�l�A���*�$��
]��j������G�[���!o��mQ��b�	��ݑ���!^\�
m�M,�[�T�:� ��_�;w�a-F�����a����@��c��9v� �V�Q����W�&}�}��B;siP w\�7>�]kB2�� �f�J��F������B�k�l�7.�:d����$���F��ý���{��f52�CR�W�^R��,�[qt3��D�@뾑$wTy���(�bl�w��n�"����H2�\��M�C�Mn���
Q��8���n��VI��B.BOl�d���7A���$��I ���A��j���}C��=܇�;�ؽUbw/.WȎ=޽��m�csq�F�+Ff�8p�DR�9�"��Fei����݁uh�=�*1S�!�cF�4��4�Z�jV����<��a��$��G.x�^����U�8��d����m���gfB\l�B�i
�; ��3[����q��t��5����8��Lu�\ڍ�7n i��4���.��ā�E��Z���3�..�gZ��xZ�#�G�V�)
�`�w5�����1�'���#	��齥@!fd�HG���r��7���d_H��p؊�c�HL9�_U*}��rهpz^j�A}p���oO�ܷS���pD�<�����S��Y3��"� �x���3���ۺ4wj$k��M4�i�h&!���ok.kQ0�'�z�>ٝY�.�DW���a�Uw�C�P��s�I9�������kd���_c��7Oh
(�P�p� UKs��h�6SaK�[@\jG|���dL�'��wӥ�7��G��}ٝJ���*���.r~h��rQ��B �b���$76#�Ŏ���*뎺UtJ�������%��j��Q�Mڊ�x��Ɲzg�FX[c8�� ��  "r��77�|I=w��$�z��O^��lě��Z(8ÚH�U:�5�|}^��ղ�������g���� ����"����������]ٵH�sέ���M|�U哤��j\M��|}�h�$�l���}"��D��P�=�{�m�]�u��w�v�4�.����[�S'
��af�2�v����(s1-_"g���s�u�HU��ʃ�=�-Vl�	������6�'�	�a����ﲏwRt�̂O�k&��u�h�{ʢ������ع2�h�v���M�L�I}U�K�vO��������5;��$�RWz�f^Ɲ�tm$!l�@�.wtd�{�<�o�2�*�Z9(f²�������9^�#_�T#����ܢ|��L9������2Ă;j�����UQv��:����*bP����;- �ԫ�7��o~�UR>ι�wo�v�b����+"D"O�&�MA�k���H�]f���J%��=��U�gK��\� }�Ϊ3GuI��}>�U}rÝn	ġ��j�Ϫ�ȇ���2I�Sת� �\� �����]��9���b��i�8^�p,��mW�m+gW������M�Ϊ���!A� �Q[�]
K�ٱ]ZI�	 �n��H9�L(#��Zh�lT�5Ƥ��M����z��v��Gf��C#�Ʃ��2F0������ %}6�{�I�O��/]�0s��X�u�<L���eH��u�r[����9r�N�TωS%3)��5��@Z�pQ����4d��gE�/L]i�%	s�,�}��ի.1w��8�]y"A ��Q�^m�T ���$��t�	�ş��aҤ'v��%��wefdY�Pd$���ު��IoTL�$|VRX��,/t���-RQ��@uK5D [��\������q�$J]��T�I-ꉟ$�R��\C�&��r\%[����0&w�f�$�T9I �=�\5��N
�J;*���7��*8(�]�(�MZa���e�PM�U�I/.ډ��H�����/!S�im {z�߻G�Ь�]�^�`[�Q�����}Q����<�{S�Ev���Ns����wR[��r r˅]Ѫ<s���y�X�a�:�ŮtІ%��pV]���
�퉠L�sz�gv�p�g�zz�u��.E"�d�����16m�+m�@�i.%�\��,D5�4�Lk���7���n��7��z�ˡ�q���k���\3�u\��Z����XNE�mR���X�F�GmXj2gm����ͯ�\$M�����T�K�ʆI$�(��f�E虫���Ԋ�H�Q2�s�Dl$�-U(�5��ݳ-U��֮�D�r�).���7I��{��gU$.�D�30��~�z- _=4�:ɺ�{y���$�J�e"R]��sHC��*uA.s�ܹ�]r���G��$�Zd��l�tv��IKD��hpS.!Or֒I,�ɜ���ֺ*OD���V�&RI$��h��]��%��}��[;���:`��e����F�Le��[]E�9��%hg,�&1��چ{�n�i$�]��T��s�vQ��t�$�M�3# ��a�B�I>ꪤ�;�6t�����E1*��R֕2�V]��j��;��������g;5����6wC��BSv-@,?��� Aٸ�ҒD�-��H��MR(%Y�x�
�DBlBM��m6�^K����D��ιɎ��t$�W��RGz�j��: ��&��&�&�8N�	$�Ja�I�̙�%{��K�v�q���/�ics�Be6T0螇��I'��d.��^R�C�P {� �GR�	R��ee�ufBE�&-(���I6���V�š���dL�0��￯�k�/�o����;���W�[Jd%x�j+�$v�pv�)�� ���13nwc
t�	�ԲQ16��"̵�H��ْI��ԦR$�;9q΅a���&4j���Kg���Ib�R%/$�P��SG�>���*��*#�����X*g���[�u��y����Q+n�{x��o���r�<�lN�F� �ܡ�R�c��$���y�m�����S*0����+n�� ��3c��%EP��M��7{٨�Y����ٺ���"o�/{Q�<�E�,����
�BM)xd	�/0���P͆6�^�bQ$Ztu:�6k�D��}����~/�{���R=��������>��U���}��p��wi���[+ NL��U55�C���No�Z��7};u7��^�W�5��`M�� �d�OP'B�k\�����Vn�A�Sty���	��|:	���g_,j�������q��<�B	��=�[{��=�;����=]�C��<
Au9��[�w1��h��*��.t�T�(�f�8]����wP8wݽ��2P�,�������"�Vkg�bq�D^CB=��oء����F�.iܶpVss3��M�C	�|�g�8��y���ss��Y���\6ٮ�=	>�2�xe&�/C����T��q�3�/��ˮ�<JaC�lMl��`�uz����}7��I�%����B��[eLT�UX[j"�5�UL�̳�D�l�+���EQE��+RV����bC�*�"��(�[ikbʫ���m�������1+ŁF���
�K�aU*b@P���%T*")k�ʋ
�+!q�̲��X)FE��bVT�(��1�j֥�J��6��@�L)q.8�Z5�PRV�V+S̠�%dY�d��U1�d*��T�R�(�T�(j,�b��-f!�1��
T��V`�m��2��Q��	$��wx��m���o�ܶ����xI>�~�!���#L#z~}e�>3�$�7�U �J��rI$�Y�Y�U7� ��~�OF�g$3JåHum�d$�Gy6��^EV��$�ʢI���8�K�0�dc�r�R�$�	���n.�Ő�F�#�d������}��cjm7~���U��ԤJI$��6���y��J7T��Q��$��e<Ix5Tl8)���Q'ycH�;����T�r��I��R�	�]Ɇ�1�S|�:��Ѹ$���Ҋ4�:��A"Mڂ�&#8q;N��e�r�L�	$��Őh)�B��t�eB��y3�D�J�P���+��6�)w_Tհm��{Z����{���U= �2�'T�޵o��ڗ�::��ˇ>B֧I�H1sdn��;Yb"��{������J��S!$��QP�E���i��&����ەR�1)r�NR%%��E$�m�P��ҫ; ��㏤t3�y�[�\ɤ���R4��E��)����g�fa��x����O|�����Ow������&RA"oS.niA��l:����K�VToVa���y$5j	%���R)*ޡl����;�~_�4�_��}�9ݓ$��8�4���.RA"n�h��WuP��bKJm(�OuF�����%�JH�PIa+��Iy#�p�+뙈W~�-�m)�������:	l�URI�fC4S��a%b��>M��3]�B�I/-쉐�gf�����4�T���T�q��VeE<�dP9=r,x�p{.94�>��{ק����W�������ݰIh�m� �8���[%����N�-:Δup7;v�t=zG5c,3v�a�\e�@f!���#,ʛ8�e���.�kb^��"���Qְ�,��<W�tGbieK����<]t���n�N��7�쾳r��X�=j��5�jjn:�OE�'0Wd+,=�����XH�s��l��ڵ5p����{��E��&��Sw�4^I-�%A��k/�q���~h���veU%��%Q�&��&�&�Fud�T�f��H�+;j���[�!$#N������ۅ��4�7:� �e6RO'�U �H�dL�RV�Y�q-`}��$�I-�ʡH�w����8�$�p�Q���L�m����Ol$N^eU$�K��"e$Io*U�������d�*��i@M$�T`��H$n�j������S𹜪��IvdL��).��T'2�j�xdk��U�/���vR;�f��\2�1���m��[��	�&��U$�G3"eJ�]ɓ�p
�Z���� 
o�M�/��
CJI���M��J@t�_�9�Wͭ�K��ϯ�K6�gtG��am�,�^ŷmM�v�d��2�Ky���������������[�D�H�]�ZF/��v
�܌�̓��J��@ME�"�/$I�M�H%�i�a�]3TA$��$�I%ܛK[�Bi��EW����/d�uef�$�G50�)$jl$�H�y��Zڀϥ�Tz�d��r�l�ƐI%��3�N�a���Jʇi$�J�?4RIN�T�\	�/�#�DD0��Y5<Hr��V<��XS9��4w^{|�\h�a���\I��ڂKIOoUW����S�ⷥ�
#�m\L��&�Ac�2	�q!:d��ʢu��UQޘ�I$9�	i/)��E��]�b�$���	4Z�bI{]�U/$�S��.�L���(�_vV+gf����%^d�_3{��b���3ekԅ���ӡ�ޘ�������؟�A"{���S�}Rju�C�y�	��JGz�-v�A"M���+�,�ڪ	w�����i"k���؄6Sa�$�r�R$��ȑ+�:rj��	%�,$��uP�I-�ٽ��A�(�!K�4�� ���3��M29�.cF�s��;МF	f��In�P�^H���&BU5y�NQ/�a$_~�/�n��n�'ߪl��{ ���Ph�WݵTI ��&BD��]��ʶ�tl���@��Ϧg$�d2L�&��=q4�;�D��ٯR+�!�ئRJ���8��-Uy&ӌ�+�H�y�TJI\v)�$�A-�ֶ�����ػ�1�����T˼xntܵ��{:Q��Ni�hvb��#>���׳�����=�=�(?$�o�Rju����a�A���~6;��o\2Pꚪ��K#1L��'�?5�/ ���W�m����$9���
˂Aұ�SmۙR�{��t(.)��{=UD�˱O�$��Aw&��@"E�ت��]RM���RK.�g�1ro�w&�K���Y��wV*�^H�\9I$�]�	~IA�7iU�%֊Å���w\3)n�ZUw�����[�H�m��H�w�2� �d��'N�Oz�� �����A=ĒEqhI�s	8z{��	t��	8g��G�`HjD�X	I$���c4dGnNX��$��v$�I%��E$v��M�}ު3J�8��;�g�|��kvF�/8-���X���ř����`(��:�Z�ڵ��v�������'s\�غ��3F�̳&��֭j{n��3Ş�=n���{<s�y^��1ָ����=�1���P��vH�s��y�sv��EF$�5Ť�<�C�v�t��aaa�>{�]����ٸC�n�NQ1\J��f���r<�ͼI��5]�Og����f�n�z	���v�Od�v�:k����C�1�Q��ع�t���Q�߼�?R~a��_��s�i�^���ȼ���~	�ē)$����P[m&ê	t�P�I;|�.b�쫼Y˥I�P�H$z���Q��T�	36"�	�pӓIw&��D��W��A$�t)��R"媟$�I��h��+�����bL8M�n(���*�*��T$I�O�$�Hv�UI-��.�Cqs�^K�6��A:�mDN]�uW�RI%�-O��\k��4�0Zo�$�Wt�$�GZ��K��j\�ï� �	� ���ـp�&�t��z�2m��X5�)��{��*ܡ��=��~}�I"P��S!$��0��ۜ�i�AuoUR��+��4�j&�p�L�c�p�Kx��jU�+�j(k�wEԛs�;W'7���AE�ٲ�2�ux�я�(̖���=���.��8���T�Z�M����7Y��a�{��:m�i �+�v��^K���L��y5�{6g��՘�4���
m�:����z�$��֤JA$��Ήٮ��H�^mU"O.��$��PY昇:4]�A9��d�0�j�K�/��2�I%��$���tO�8vt��Nm��իV�PC�֦RI$j�\k�qء�IOv��D���2I$���S����0N��S��P��81�y�b:AG.`cl翞x���\�6�b�fI��,�̤�H�($�Ts�k�쪤PI��3䒾3��	�M����i%׃D[�Eᬻ��%��2I$���V�T��Σ��%Z�*<�	��N�d$�=ɴJ	k�z`D�F��t��9�v��<x�M{s���4Fݍd�r��i$>�q�9��YD.q
j�__�YD�)��;Y���|<����t��K��S!$IwɆ�`UBm7	CI�|�$���ܞx^JӴ̤J�M�$Af�V]�/78IJd����!�NN��S�IgvP��bp�5�!�Ԧ|�+�*��D��}Rf���TAIDG6!!	��p�c�����^�.���`;����*l��}�o����F�0�H��}TO(5�.���g���L4�# �2��2c�L�vc�N�a����R% �IV�Iy$weW��Fnzɝ�]I���* �0�j�(i���	u�W��K��'v�,���D��^H�vM
HW:+��8a5Iôo{f��C�=($I�L2I$��w�@ ���nd8v�0%|���,dXg��Dޏ��s�����c��:&�龤�P��0������g0�faA�{��?�&�6�6:��-�PêK�UU�_/�L��뼳�z\���PKI=�UH���J�I��	ZN���Bb���`�$��ЯI/D֦�4��&�\�hg|����p�6ӳ�]ɴ�If�L�D���2y�2VGd�QɴIK2�����LBp�!�[jD�䄅0;�	RwT���+���TA%3�p(0����"��2��:	>����X�T�H$�N#�e!��:I���uU"�Z�S��ƩAp[I���Wn�wf$^i5T��h�	O]P�I�%2d$�[˺����j�J2j�RUΊԠh[�J���[ G��	��.M�I9��TMx$�6T�D���V4�Gl�gs�f�fo���J��}ǯ���u`҇�c�`9C�L��B�u��j�6��iK�����0��̧m巭�x��+�vgGS+8Gi�>}�����4/\������~�f���P�x%���2�D��a�n�fҫ��v��{�(M���g�n^��9��$97� F�M��O�6/����I�_^=�<�\,aX}ܞ�y��ݼG��]7�V�������=W���D�Ĺ�wcN��6 L��[;���b�>��~j����%�7�y�ct}��4n���ۼlI@0�;��/[��H�š�ݺ'��$����X��\�	�LM-lh��n. ��r�kҦ+�7iuw=8�)���YWM+��4mPyZ�N�+#�NI��"b��y��-x����o�ȗL9}c��m��sp{c
5ө����5�h�pU�v�->��{�}�]�p���������Г`�	��v'v(|Q�&��.�ZY|߬4(��wMc\3�POޖְ呥��"�˹p���Q#L]f����B�c�akY��n-Ҳ��2�� #�+����e�3��y�޺(�s��K��Gf���J��m�d�0��0�b��J!X�	1A��*)*J��J�����[J��RԵ-�Ŋ�`��h��Ȗ�f[�f*)1��!11�kh��.6-J�
e��j()\dU���Z
A���I3,*J�b��1d ��
�e�X,�F�L��Z�LL`�q��r�X
�d���+Rcm�"��1�,�$ư�LaZ���
��Z��\��*�"�XK�2����,*`b�
��
�.[	R�E+�����Km`cAc�~���k�fiO�]����\��W�}���70;έ�|[;�X� ��e��%&9�JʐN�m:�vwqGK�����9�)�l��O\���n��b ���Y�P�5"��.������\=�t�u:KԵtδ�h�6X�i;����7��I�5��������ݢ�p`��=[��7R��&�[�\@�n�.5m8%�����	+q	��d5��EIh�bo1�s��N�y,7d�F�%��q���kU<�7<o=b��77��9 .�;;��Fw^�\�\�sFz۷\��c%{az�N��6�(v�<u�G�{h_US�Ʒp���ISb�-����ԑ�H���^�@|�P��{{FݷV����`L��Բ�	�YR�Ź�L�������W]<;�]qu�=F�=t!�5��k!��wn-�8k�,WS �l�������z���vcmz��'����WLq)�Hy�1j�h��2r�� ���x累=4;Z:��n'��15��Z�[&líC(J&�/*�4�
%�d�M���wW@r&CYm���� q�������[�x�J�<�]4����맴���W��L�JG��6Ԏ! V���^^rW)�܄�o�sr�İ�s+��&Jf&��a%(#q��el��K��}q���o\ٝ�n;[��4Ġ���C�kqs'�5WV��ΉF�rcm��v�֧j�A%�j��]���n{V��f�e1�%0�=u���z�@+�F�L&��lB&��Z]X+?�rNrq�κ.
[�:A�8������7b`��r��5�0�W�9�P�WU����v��i��zm���gp����x�f���J�;�y榧�&=�{n0�C�к�����8�.b���/H���ۆ6�FSƺ2�����کv^-�i����׶Ӷn1�dn� 1�973Y���j[�@��Sq�:�+6�����:�0��%o��Q(%��3) �]ɓXut��5�3$��Ų��2�lCm9$�,h�w��y���ݜ�ݪA$�����I.��E%�6^�F([3�'ck�F`��!�]j})$�7i���^K�D�=q&*mKۜI%��2I��P^dd��Z��A'��Jx���ވ'BT�T�%$v�0�IywvS��#h����oq��F�g�T�
 �-���ג'o���gllO'D�	$�U�	%��ʓ]5�e��R�K��f3.=f#�s��]$�#8nҀU�c��o����z+�?_��=S�D��j�K	!��UI�f*']�N�I �rm/sb�2�Fu^K�UU�iM���ظF'v��F6�F%���QpǾ{K����F�ͅnnL�ʸ�{3m[w��  |�WҐH����I$�w�U�E%�H��CyЎE,'fDP�6�6ӣA,��%���I��f�p���'ZI%�K����e`JL(n8�Atu���<��	��r��I/vf�PH�])�؎%X�l+���U����p0�Bt�'��*�	$�d�oc�!$�|�I$n�&��tIr��QW95�zQ<f!�5Э�vS@�XX�&�D��R�Z7W�1ۿ{=�An����	6�D���&i%��rfBJ7�<ʊУt����][�&�s��(��J�%F�H�jw�����'�L����H%�\�$����������-��p�Ma�79T�H%�d	I$���h��|D5iWǓ3G�Y�MC��2�q^Jy�z��ֹ�u���HDM��0v�]ب�xxnR�~I��RMy.�$�	L���M�m�$���l�Օ�L��ޝ���H�&e$�'ߏ��@ ���J��K��V�'ǹّ)$�F�0��(��i%��TI5����'0�=���,���{�)(�{�m�q��W��X�X���Z6)u��j�Mh��6�4�E��N��D�D����I.��J�_Qک7yRI4;\��B�T�
 ��j��T�JDl��T�k*��Vs�$ϒIo(%�n�	�E�&r�#ɿC0�$�� �[����N�.&�v��͋�*⡸�pKMts�vb�V@$�RC_\23���}�q}rk���gF.O
�6!�f"7�+r	Q�i*.i�k��v7�t��y3�h�s��ͺ!�{���])�[��&�Ce�;�z���M�f77cGK  =����{����NTߦ�x;�q��,ږ8���e�Amؼp9v�Cf.�h�}��OvG3�R~'Ĝ�a�Ood�.qa괻P`�n����'��!5�c�1��GZ�;HiY���䌸k�����TN�Mb����ˊH��`���	�^R6�LZ�H��$Oc�Hݒ&s�ſC0�T(�9��e�=�w`����Nvl� �˚져NS�D��a�!�T5ц���>Ay���KG(�����6��t��������>�R���ܱ�49"�w��x\��Esbz�ً���-��qc/�d��}| �[~~����u�=<@n����-JWk���顩8lQ�Nz��`�왬�<�V�P��s��`6�^����=�=��|�otW��c�̔�)��5f�m��NY���,���hK�Kod�.��1];]+qX��Y8�z���R��Ѷ0�ۮ��i�o�^	�-�
�i 8��Y�a�mrL�%cL�S&���>�'��vWk���~i�>F�uPG8O��d�{u#o���� ۰SP��P�_.���k쎘�Yju��w3$H'ܹ�`&]Gu�Ud��Ȧ^'�U i��U2�4���� ��L�F�ځ���P:��E�Yt�L��H;n�	$��3��Sh��i�R��T�l]�K!��
-0 �ti��3`�s�>#��h#����[��<���1!*�HprvL��v���#v���\�{|;aCN0���3�(>4�	�A�͓ٱWu9z�
��dc��V�A73-��ݬF-�Y�����Ὧ)<�%���w�i��R�&�����3��	��B�N�葡fϦcbC������s�O8a�$w~~`���������*b";*�J@vcL@yǍ�Ю]�e��Ƹh$����V@<����hط�H��іb��`�l}�S4��qj:�t�U�a���)��5~<�`��}"i��̜�-v&I��$���B�_>�ཋ��,x�L�-�՘pX�%�ݬu�$3ھ���s����������/y��F�s�!��p��c*��$�sdd@���h����A�R�oUq�}��`�:�l�6������.�&�e�ݤF�`��]|q���+<��Q<1�j��Ae�e���GF��u)(�;�'��.Q�"UU(����{������Fg�4�gꠜ�DT�˒%¥��|OB�{���`�΃�yt�B�R����������E�� �8c�_��V�GoB�������r	��ލz�����Hѹ2�dB�mYmt����5�,ԢE7������؎dz�'� ��;�:��͑����7��I�J�~�[UBZ~$ߧ��E�Ý�� �gL�yt�\e�2++�m�!�
r�m:2_�PP����Q�q�����@xꆃ��9o���c�wT���d>7��H�� #��#�L�#8Kb^q�p����e�%��IS7�P���WЕ�ظ����2����c~ X�y�"|�~LDC���:��$�ٍ8���Y7�j�\u�a�����r���|���|�tr<�&.k�����l�n#[���jxݒm4��ѧ�?�A��9�IP�p�7��n�an�x�;:�|I4�SP�:BL6�Ry���8��s;}$�yl��I�� �Ҏ������ �M�����e�U
-2@$[͒Mq���,-}�I�-�� ���� �D&��c�:��%⡝�����h-�uTtFc�Lw���Zϛ���V��4���vҪ�fZ�O�]����4 [~�v�hx���\Θ�۫��
��-M�B"v�j�Q��}Saɭwr/4Hzkgn�:��H��[[x�����O���-sc��6�]3.j�^WmA�ң�RE�9�d���lD�q��"[!����DLm��]���9�nq�����Z��6��R�|T8�O���6����sk��l΅w\��4��f)����5�I��a����g�����ou�=qÔK�m���r���MhF����u�l7���l�����W�"�
9K�Ă:�GV�	���)�i��ҙ�VC2�E�H�-U�3$¼��ԭ`�gUA ��#��D]�o��)}���L����Ȋ�v��O�"/�bٹ�qFg?���H+x�'��n.�'V�+ak�	���̙�r�BL�
��{�yiWo�l�~S0�m:9��@�u�*��R�SA��T�����۞��;��zͤQt4�:ҖgO��AꉜsjSPd�t43�������e�q��7�j�tu�!ژ	0w6'�w� ���*TD1
��?n6N��c�o��63W)�8�,tJ�#1t��o_n^�tu����m��z:6n�U����'gB���N?<>N��g���R����:Ω嵅�LUvi�6!L�.��i���Kf�*�d�_H�=I�hcDC��ݾ�����E,E^uRg\?�#���͚��%�`�
�$Oi��S�e�T�'a����̕�J�-�T�:�� ��4���:Tq���2T(r��t�⣍����!j��6�&%7��Sa���|[|�z�A���������"[�#�n|ܓ�<چڊ�V�?UUs���Uo	>$7H��9o ����TeP%��T��aD24�+�$��l0AQ�L��#��B?�6	�?P���PB�\
0Ds�n�
��|�&��_-'��hlJUq�S�*Ɗ�H��ոF3y+���ҽ5\ONʆ���l�wr8�t~��<�k���uyVge�Q3z�thɴnR줷�
\E�{��=��F�}�*�@^�r\Aݢ�E�.p{����f_][=_-���[",�_dj=���q�����Ќ��.ozw&�gn��1����v���j�+��nvIޣ��X��}��mw��ogn��8'=������9z�o}��ǧ��>{t���9�`Sڷ�_ɝ�������a^�ys��'�	���;]o֏a�����矰`|֐�v�m]��c��%�.Vk\��WH��ѵ~o�7����"�6h��Թ�,�
�ݶo�v�����|ϻƫ���4u�G5��.I}�<��5���=�K�F-���_wt��۝��l�[�|�����{̞r��ϰє�=�>�cO�i�/wW�Bz�x�x�)>�K�V���'{Kk�=�N^��>��ڴ��l�y{�l����)� ��0f��{É� Z�����.Q1���+
�r¡���ī
��T��2�H72�1��W2��(�1�Qd3,�LE��,�P1%nP2ѹ��)
�Z@�m����Ld�r�)W.c%b�m�%Pq���`��R���$s�� ���!�d��1&5C �D3*V([C���dRfY*�()�s(b[k!X��(ȮR媋%@�aZ�**���D��m�Ԓ�V���(��آ��j
��.��X�
�
����+2�UXb)�P��$�[Z�Vam+R�h֫*-qSAo��@{����?��D>�E�<�?Z�+zV\�i�5�@]�X �oM�S�-e�J�� ��5�6�R6�!�ΥD�Sڵ=�b>/|�.�uP����]~j��$�r���d�P�k�ƽ��v��*�S0���G'��kzjd�A���'+�S��(s}aޏ;vz"KS��v�7�BEG'[>�;���_6��:�0vq䮅�����6�U����mP���3yɳQ����@z��A!��T��hq�U�[E��հ�&s��$��F�X�[�"y��©�Ȏ[r�N��݁O�rv�Qz�Of��d�Ώ������E6/�(A΀�D��D���? H-��mj��L�*���T|�pγ}°�Sl����p�iu&��f߬,���͇C����n��9��˻ Z�iRf�:3m׳�'�j�bt�2O�U���3*�F�ތ	�~��rg8�Q�<�mJ+�K��>k�E4���uP��|4��]�W�:p9� �T'��$��^`��
S����x��ɐI:��m�<3ͨl��Dw=�]��I�Tŝp�=�b�f�c+{&K}Ȧ�C���>��nI����n��������L�o+}4��@�3c�O���'���6�U&�o�W���b_*~ŏk<&xw��HB�{O,]���b�f5Ce/6��Fvm�n��Ͳ�6��������v��=oMҜ���]�vl�=%�Eڡc
k t�Э-,�։kE)�Ip@�[f��Cc��adC�'	��mt������Z��E1Ig ���jkm<�m�ۙ��J�Z6њi��뗋����Y4r���_A������m��K��Z�	������.�����ǿ"7���>4ˆ���p��o��M���41�FC	��虴9]�q�5=�BN�h ���@���<��n�3��jjb�]��ж����Nm�H�ˆ�7���� �T'��ٙ�D�����[L���l����/kz�H��$J�A��37�����h7��ޚe����i�Ew?0I[�>-l=S���U׍v�uN�5^rq�����݊x��&o������ɖ����s-�I�=[�M�ۨ���9
�H$�c��ĵB~b �U�V�ȟ+�)QEj2�S��M��R�n:W����]��Gy�>z��Qe�G{�9=��ҕ�D�J���(x���	���䑥\h!~��Џ_�ԩ��,��n���D0�mHa���}>��L,����ڞ�y�wt�����of:#ɖ�"�hS�'i�� ��x�O��T5<�+���H�?=n��D�GK�<uC�O�g4>���:d�	�Ҙ0|����v�A���l4*���!�d�hlV�3,�C.�]a�7ϯ�~~������ �vȐA#�JfZ���b�w��fu�A3��]��J1��~/9זk�����)�L�� ���툿8��ۣ�:��]j\�?1Z�+z_��W�	�;�9�b�䜩f�*�fFE��ٱ�V���N�*e���ڒ�L�WqN��c���y#�@��� ��?T0-kG�S-C��m�����|�M.���w=�ඞͶ1{�A>��>s�1�������U誷L��u_A��	�7�ӽ�^Z�]1!="$���N��s���ě��hSmۙR�y��'� �*��C�����`�H���D��݋/t�ݳ �;)���Ѓj!�@���Q9q~/9��Mq����*���39��o=$'�L�Tw�Xۓ���6S�Mý촀}R�{��6�:fe�Aڎ����H���X$:�I=��q3c��Lq�am��!��I{��xo��hNK�^���w>���z�!%J�{������2A�l�0�mO������D�vs�m�\*�Y�� ��a�{o��ۓ�����*z�	P	c��gmt��ź�Ѓ�n�Řv3h�n����᪆ᔢ=<���ogU����j��-��Ƙ���D(�Ne:=/�Q��/��-T�@W�Z ^�u*�ɭ���P1�4� ˈb"��B��>>��\Uv�@,�m~�H%�LAPKNe�'��Nc�XH=7���'ĝꍳ�[@��j��=32؇ �Gs�H��*ri�ܢo�|�^��|}�r��kyS�`��l��ټ��D�ݗi�[����y�9��l��`0lj�S��Y���{��B��:��(m���Y�xaۭ�nֽ hغ8��q�{��nϧ��=v+uӏQn�OfH��zOj�uL�:�1�@�v�v�Ok�� 6q�Zlß��=XX#���SZ����-�W�G��ӭ�*=:��9�GQ[=���i긕5V��wA��	�u&p�D�+���-���[a��9�BPMia�m����"a�i��y� ��x�GuCz��j�B���BݛT�u�(m3Tb2���eF\^�6	#7z} �T0IpK��k�C�q�$�m����{_P�\��E�o��}���b��T��&�qDU�	ڧ�Z�$��Rnܿ����o*��7��C�h�"q{:�Y �[�Xo�B�g��#z�.��^*|�.�5�K&�:5(�MM`h��풭4�����9YB���y,��~#;�h�˽��]3S �;j ��BM6�Ͷ:�O\�9��e�J�W��)n����î���GK�k�l{���.�#\���2�5�fg���q�|G�P�I�?��pn��}�O��)n\L����}�!j��u�?.@���h�͘�蠓I��9����	"g%4�U��#���?�m���WP�o�2����[�0Nok=�30,��O�7�߈]�;yLۜ��I8���<"�@�X�m2�f��֣�s��d�;�������J`�ܖ�_���x�Vu���@{�سۑ�3.@r��_!�����9�W\]�0I;[�>$���U�^M�Π*��B%�p�W�6��ΪBר�d��:�h���ʓ&��S�T[�w�����mS���z�;�pog��}�v-�xpW�]�O�_-ݩ����ߪ����$nYV����5�s�����l�͑$��TdB��%͑�,�)��)���*��_�����A�����:@ �T0v�-�[�Vh�l��ա����E���&�(ڋ�#	�Z.n�_�qD_�oC�>9������:�Nz�+P|����K��JZ��?w\� ��u����>�}�_ �-�x�&r���;�_����r�v���e��~��e(�œ�}2}�Q��u0��M��;wj}��H�����Ոv�,����q
;\t�z�zm�[:��̅��ie�fT�鉆�<��(��"n�&qCQ��_��[���+�Ç�+�����"t��4��_��_V�\0����O�mQ��EB�51V�Ķ����Rb��f]��aY�~���	�����}2	ô�`v�f�Xk�Қ�B��d���2CrmpL��EW��l��5��o*Z��$b�^g{������1ݻ���G@�R�L�U�G��%��Y��b$r�L	;��-tDC�q0;^�s���C`�/!�|Ws`wzW{Y&\�=hg��<� a��hlM��s]%�U_�Qބ��*��Z�t##�����	�*"�s��'� �`9R���˄1ۉ���6���5�0��B��0�݌I�Eŏ%��l�|2�P�z����?G*��ȭӾ���Wy�=��N�}��;�}������qw��B^Z�y�.����qG6Jp���n�W0���{�Sb��K�Ƕ��sR���:��{X�`NW��z��8z���N�D|}������v������p��ͺM^rs���J&��@��m�Q�]��������/��y>�d��u�s��ǆ�^�x�Yk��gwH�r,*o��.���mQ�Ѱ�[����QM�:	�0�P;��[HL�ZnE��&Nb4NWh��2}|��:���5�'�z�Ǔыi��t���A��"��D�fT�CX,�i�e/Se�sb�)&^�[���n�D�U۳��ZwFǺ�����p	���CX����1���yլE����X�zl{�k�U;����.�G���lf!Uؤ��Ν/Rw$�f����d��K�c�^�x���<���D��w5�"0b�̜�wu�Jol�u��X6��Ci*�yr+[�383Эz�<F1�j�6���5�u�{�ͱ+��#�fPX��*ALJ��.$�\�1
���
f8�J��"Ȳ�U����V�QH��T"�eB������R�Ɉ�D�j�d(��*B�U-����DU�dP��)�V!D++Q`��#l�U�
�0�J�+�X�KJƔmY*�e�%AIi`�e`�E�-�Eb[VR�ą�5��")m%jV���-1%[jV�1\s)Qk��,��+m1IQ@X�j���J֪,�q��r̭P-�S6�YKd-����m���
*�fb�[b2�Tj
��Aa�����Q�,�H��T�-l�++V,�7�Zn]c�ӡǗ��ݧ7 j|�v |8+qr�4a�B��Zp䤥&�nb�E�,��g�<�R� ��O�εj���	�#��v,ca��ݙ�E��G\mFG&ط\�V��k��]��Dp݋D�K�q��#g�bx|�b:� <�z^�Mv��ŋı���K�:�pk�H�;��vG�m��^'�;�z��Å�΁�pV��z�5ї�pB{N�N���ۧ��^����`͙�Π�e�rJl�bf�X<�lD�Cq\U\���n�+&z���@������m���n�4y�et%�	x�"q.�d13�.`�2ԣt�x��`1��îv�-�>@.�mY���h0��Fg{���	J�yfaq���0X�[I�s����P��v�x�M&�6��z7;a�Ѹy���{P�d�\6I͑]=q�c��*���Y�f�~�7ß�qz�%�������F��ـ2�q�����7��{�cb��m�b�j�H,��7�e��n4���>�=g8�n�njZ)�q�Ϟ��bl�<�r�ѣ�[),���n�W��6@"�Z�)U�2魥�D�@��RK�A���ki(,�=�ogK=��s����{p����'=��^̥�q�9��mwS^=\I� �R9���;Q��<s��y�vs�.@����!K4�C[
b��qX��5�%�v��t$�pC�i[�5�l�6�6�n�㢋Cgu�u&"�٧V����nc/F��Ϛ���۲��=�^4��20�Z��ԣ�[3T�1ՇY轝�u�\���ּ�C<뵁-W!*h&��g>z��8��-�N7Gki���h�l��T�D\��qlG��7k*ЩahF�L3Ͱ�5�vƝ���"�ƒ�8SJ6:{uz�4t�ϧZ۴�k[�[��f���CUn�K�����3�ܭ�̍&s�	�S�bn"U�1	R:؆)s����6�5��G�[����LB6��dU�_vҨ~��
����1�H��6�6#�I-5Y��/�s�|�_ߺ�{h�����ޯ�h&���Ne���GsL���:��J��<F� x��_uQ/ φ���q�\����/ݎ��=,0|g�\�4�&������=�`�m�06��(�lq#����Bp�|��/u՛n�e�sT�:�B}�vaV_��r�� ���v��x;u��"<m�PI���f���C���cd&#��'.�d�	�ԙ�7�}�{O`x�$�Y�"g4�\�m�L�+�Ů��qoxO�/�w,n�d�V�@$��9�}��MZ�~�"���~�^lfgg�^��-U�\� ���@��)dG�~���Ϧ�z�3,��kfzĐF���I'vF�MZ��5������2A�.�rmpL��EQ]���L���$�w9]I�O����77/��=�A/ ϊ��e�����m�Ou����3$]I�|wy�{3�hL-��g���(aw@�˅⥛
`��f�Ԛh0��x*6����S�0ˇ��{�����nM�t�>$r�LZu)0�mI��a��!V.�7i�w�j� �2=p���F]��q���Hư�6���� �oy�H���g7�(�X��%��'�@i���D�>+��I�[ڥe���8Y�r��t�m�-�낶mdGgW< �]I���a���8	��#��ª[��+$q�B�6���/x#�p�	���!�&����b"��߳{Y70�q�g��y0H$��G����H�U�Y8�*�uڟ�7���J�������H]��ݶ�i����K�)�֮���À>7q����L�R�'^��UFT3��lY���L���w�5h���b�f4G����!u�U �3� k�z��m)!0ZmI�� ��|��9v����@����6��L�JF9��̢�-�۱�ۺQ�N�$m�̐yu!ٲbER�5::!���E�����7�=�G�zl҇��U�=����%�3uB)�S���"\�Ɲ��-:9��G�p�쬿��>�H7M�A�fd�'�Rf�)\5e-:0�D�~C�iZ�i���5��kW=/:heӫ�<��}}����g8��b��Wԏ�:��\Vw'�˰�� ��9&.R�%!�ؑ˭�;%�і�f��|A�ԃy1�H�WT�n�r���#��֘e� 'W��rs�	]�گ�/G\4�`��s�#V6�����d���p��7�gӱ���d��ʤ{QNĶ�%�3��;�r�fz�j�Q�^
ꪠ�%������,���	�ᙋ5�9o�H�7�W�nӫu�=�A�n7vv.���5��&M�>⽮�X��{�y��r߈ŤSGј'p�-��HZ�q��m#`$�����f��Ճ)Yet�C6A�,[��nκ�q�VS���G=1·kNq�8���O8�y��q�q�v9��k�Fm�f��n�9�ӕ��<vj�SE�:z���Q�ݪ�Up�`�g��ny^�]��p��=��,s�=��FT���o�{=�7:�:o���P���� w������=Ԩ̖	�Fh8Rۉ�Gv���:��y�ɷl
��� ��~`�Wݢ[���w91���&1�v��'���t�{Źt�� �n�r���#�G�PNg��{M^��%O�@"'9��ޛlA�����31)S��4srЯ���рET�w6	3��>(uU��s�6�^B(	J�L��x&*Ę��LSk�.�]��m���
y�9��ھ1�7�0U��?�b�pY�.�K���s���� �wL��XkF�mTX�}���j"�%멭̬ND���hՄ��-�n�C�c�fe�$��9s�V�f�E�c̭�8�+�$���|RT��)ǐ�w��In��%��T
�n��P"=[�gA�ҟ����r�/�0ɈlO�u��P}���:�~��r'z�������{t�@�h��s����]�	�ձ�ȋ�	��6H&�6D�w�/T�a��Y�BQ0������ �G��g���O�Ġ�������<������ٴ����TU_����莶����!��Es�p���1�l���\���O��ov�Yn��bة��-:D��R��`,^v�GBf�zg��I��p�#P�y �e��%]��ا����;�0��)�����L�d��v��$9�"@$�\2܃|�s5h�����l��mP>3�X$.q�(� Sݵ_����"�	��޹� vck���VFb��uP!u��Ѝ��˼�o�F���>�Ke�bX] B-��sGFRc�nn������`�܌~��fK>�6F��ǲl2UvmP��Я|��	��mĞm��}��C�P �tJ������_l���ژ$�#c#;��d������πGZ�{�gѬT��99�L�)�?Q6P����+{�="޸mgh�\�m�~�o�9oOnwTH��%������~z�X�y��PH^��K^� ��7��Bna��;Ҵ���*;/��'a�#���OwO�صD�v1!��a&�`�f1C1k��5��1�I@I�������)m�0z�A��:���^[��+������P2Il��}.N�F�c}���V��VC�;�21]�!;���L�%*�P-�9DQ&��d�뺩�u:� ���
��=�!sR� �S���[g��H9۬H$r�V���R6B��� ��P�	o;$=i���5���N�,��Os�F����3��m��������;!kw���;�x��0�6i���c���A���3���е��bk�3��Srj��a6۴u����!����7iy����ܮ��u�1��Ԗ�5,@[2���v��8u0��Ԓ[�6�W�n��8n���n�GF����n`ynEh���YԜ��d�{M9mn�6z��h�n�Y�g#6��Ep�Ք1��M&-
Mk��=YʽEm���8P�`�.ZA�N"���2H=��$yu��PeN��XS����r	wV�-��z��M�9��'UGl� ������	��j��2[��μ�(�K lwh�UW� �2_�.'Զ|���w�T���)���*Y�6�ߓO�3"}J��)W���Kgt*Ȼ�b�M�:�F�	FhB�L^���Ԫ�Ǯm�8r�� �sI���DS�v}䅓*4۷/Wʖ�C�ٮ6��ݣ�`��{����<�����wV��my���0e��]������-����q"l���9����.vg�#�����a�ǝQ�V+�_M�iMW܏�{���=���;gm<���ۚ�yo��I6��dot#V�<�̺&j�B[AD6$b�L�:��K4�E�7\��,p&����l���
��-����DV�G�o]�Id�1���{9�2OR<G�B�Ԍ�(8	���o�;|�#B����=�� =��B;�� ��=uWK	���T����P�8�\�#'b�;]u%��;�<�R�trJ;�bg���{��K���*�6�J~ �]l21JSj<�`�u�#	�l�U-���y ����u*B8.'��>�T��_8��e��;���u*!$�����{EUM��JZ�5
��hfK6�h�t��᭎�-�Lcg4�T���H�r��:�����	詈�x⟴A��oQ�[�3J�Чw�̭.��w"��)�mYq�3�C�s^f��Xd��ox��OhB�y`�0��|s��8�����ym��?M���6�g�����{��{���u��'�c�k�ؓ�װK���[}�x2�1�������|�>�����j�5�k�j���z����/vC�m��_M�+`�R��:�='�o�?|��{gh˜�|�$;���o�y644� |����=���y<��G��F��{�Rސ�#Ny^@�X@g-�_?u���=���,λʝ�߂�!*̓f@'�\D��i:�#_>�﻽�y�m�x����i2�ΥgCYy�4G��wB�ygF���Z�ü�_N=��|�����F��,?_s��g�iR�ʚ���DQ�d�U\���{/p�tIޅO�x�\!*Dw7�'W�ڢ�d��};v>���Xɸ���=�ql�"���d�5�0�`��xX�ߋ;aˠFG}�ϳ��7�Y�o?�cB��f3z]x)�uv��o����? AdX�ŉV�b*��a�*��J�P"���X(�IX9q\F�)�5���Rb&2�EB�LeAjUDk
�X)X�%(UjJ�R,���UB�V�B��+�Rڤ��eDAE1�-ejEUEHVڈ
`�E�Z�0�X)(�J�aF6��Uk@U�֫h1#[Y*�+Qd��YX#�Q"�FDIU
 V�R,�m��%J��,�E�E��E�Ԡ�Y
(�(�`��b��[b�,Dm�ZXT��*��STV((bk
�A�����ƍkF,��Z��l�^fqEy�40~�9$MM�@�J1��Z�4iu�� ���t�����^:��+o�f�������[5@�vH�Y�L�{��Vv6���Ҡ���:*�q��t>��=]Ok�c)�V��c��(�2����U�������&��P�'/fH �WJ�]���lO��&I{�G���H�V
��w׬���#�(i��'g	�����M7B�a�\�D�r����M=�ӵr�o�}������*Q�N!�H=�B��b�Y�j,�y�̐I���'Ğ�ǯ#�u��;��4	��>��}�D9�.�)��0�Eߍ��#\�\+���т|O��$L���F!���m3��:5�śP���;��O��:f�)d��
q���k�Ѝ��&=@&a�({w��[;ǣqω6nW�$f�`��ȕ;��~꽑$��0�I���(D�c�Pb�*���ն�l�Є$^ԥ����yWEup<�!A�K����h�=ҙz�mN����\�>��=�&��t\�P�����y���Ws���B�����s���W˙�Do4�wwR���z��yՀCrЂ�G�����=o5�S�ZODL��v!_�!1�������wkY�5`�4c��,Stv��I͛W�bFѻ�P$�wKDMq�8	�خ"�v�8�A��n#v�!Ykf4����7Z�MѱKrm鵶�]����8܈�t���Þں8�}�r�D��`�upi�9e����rj��=pbR��s��Ȯ0�����uu��x\F��h]�T�8��k�������W>5��G.j�W���(7+ƪ봺*���*���a�ɇ+���h#o}�)��2"��ۅ �	$��s{��Jh.��uǻ���N��0> v��Wt�$T�r�Z�Mm��B &ېz�&��I(ݡ}�� 2��������~5.B�19�4v�ݞ���4�	��$�=J������2I�L2���M�!D0�;�@u�C\�q����n����+w�u��J�IP������>�y�R���DDT�p�P��F۞}7!�p�.0��W4`o�F(�i�8��4�B����VVJ2��9捌��X%`r�bA`u=�C��}^��ί��S�ߚ��X�<皇I7�����M�̀��'3�k:d�yߗ~}��5c����\X���W�U#[�o&wr���/���כ��.���؜L��(�z�G�'��7���M��agsΡ���X�ޱ �xʁ���Ѯ�ъ���_p��+��D!�ʳ䰬>�=�:H)���bA|�
�>ï��ff�5�����@����	�s�ChlIP�J�a�szĂ��AL2�@M��=���������O�x��VJ�þy�C��@�+��o�`t5 �-��������M��� ���:O�*S��=���-vl�� �<T�sF��*�w�v�X���=G������s��B�J�g��2t��FT���ߚ��g�e��l_)VW)����]���q����$�h���?~���f�t���?Q�}�4���/��=0*AJ T�����
�|����=����,�<������
$�Vg��0�0�/]o�/ڷW.k.��NЩ��4I���w���j$���s}c��
ԅ���s@t�]�
��F���~E�!T�B�Rq@/;�3��YY*%N}�7�@Dy|�����������r�^mC���[��������3u}��[�rh���sR
m���[tZ�}���]�/\�I'��;Ϸ�d镒��Q*}���6&�~���GZ֝���kk��9�w���G^|�R�`e�ZĂ���;��$m���}�|�6�����wW��>hx��Xy�ޱ�C
�}K��L��Z�:I�*{�[�m�J�Þ{����0ߝܷ��|��O3��� �:�ߟ}�6M�Fjs�5��g���g}oe��R�H�ԛL��C@eb�Ck�.��#���g|/��_�O��#�l�pd�T�<��HlIXV�����6�b%�;�}^ۮ�l�'3��:���eH)�y�����:��f��E�I�
>9�x��	Ϸ������=�=�
�R�T���7*AeNs�5���
���z�ϻ˶~��]|��i�G�f��n!�P�O�;�T����6�FT���s�C�������g�xs�{�ۣ�o�`v5�Z��������Fh����Ci�j�uLHE�!ͤ�Y�ߧ��>��75�ֻ�Ă�ĕ9��Ѹ�i�aXs߼�:I�*Ad��sz�Mw�Ϲ���\ɥ󮽠qlJ�bf��YزR^���ǻ=�^�!��}H�W/oo�Mo�V�7��|�%��@��m%G�_��qiu�i�l��9�u�- %�������}�Tت�o�x_ [�7�@m �s����$�T���}N��|:���d��q�B��L0/���Ƹㄐ{D]M�L��-*kKQ�{��O� �����AO���AH,>���pf�
J��3��5��M�z��{�Hu-9���6n�Z�����m6 T���J�F�����;5��XΆJ��P���>�gd�k��Ѵ�B�+
0�>�<�:H)6�d�s9�c'Q���@��(ʏֻ�H�~���Y�P����ֵ�s4oL�����ݤ-�-�>_S�'�"��D/"pέ�K}����YY+���C���ĕ}��Xæ������k2������J�կ����R�|�|��w���}b��D�o�k��i���vGKǻ�����|>���I����[֛u� ��'3�5��d�
$�ϼ�FěC�=����w�<a�
���{�6�q
��+%O�ε��2�WȏG_|ǨG�}��}����j��6���:�^ӵy�wO�S�y���s=�v{����R�z%$�����lz�[>��v�R���i6b�kr6jJD�.��P�N/p]�����5�n�u��F�nF�j��/�n�,e,�tz�\t\ ֌S���6�����J�5�e�A�i���v�-v����,�B�Z�bi%��M,p�ǐG�]��;je���7T�M8� |f�mm��Md\uʼ�������p0[i�Cn�3IA6i��<	�[�Ã��-!e�<�oX�H)P*_{�����f]ou���s޵��IP�*�3��0�`����5K���]CI6!S�oz��J2�^}�o�9����4w���bV;Ϸ�0:�`X5 �����t��]��W�J�ϭ�i����G��S�;`e�5��d��� ���6$�IXX°޾�w巜���װ� ��B�Q;�oX��+%R
s�sG�+>Jz���ۈS-S>J�>_�kH����z��ZA`e��c���`T���9΀�AH,�}�|�6�g}���<"�X��cV�~|�u�̹���i/\�A�H,�����63h!��>=Z6�h��A�Q���%_ �=����X�s���m6�Xw/}�϶��~bu�F�h����+�5��ZƵ[g�־���j۬�
r2^��ZgC%H(T�9����I�($��<皇I6!Ro箾���u�^�L�����N��4M��~���K�	�����a�s��iH2L�{��s7du��!0��T���P�c�"9��z�A��%�+.�3��埑�+X ��>���+(�X}�|�:Cq%B�*�����9zΘv°��'.�s1�kp�M�S﷽��%eH,9�j m*�^o��^�z�~���k�HRӜ����Fh�9�bM��ytkZ�zi�&��t�w�=��y�I�<*$��{捤�IXX°�s�u��%B�>��L����O���� � B#�c�E �(J��HD1,�65���z�I�B��u�H.��{�/�o��@�ANï��@m6 VVJ�'����ĕ
��u�$�<��:`f,����Զi]+5��8��R�m�T��~��4�5����C�B�o�h�&�X{�|ѱ�@�P*V9�i �'�s���{�	޺ހ�aC�ߚ��>W5�2!-|���~�_|���UuLsޝ�q<�y��&Щ*AaO=�ޡ���Y6'��:d镒��u��L��r���'��O����PM�jh�ay�4v�R�:�=Fh��#�N���V������b������me㽌.��J�5w2%^	��UA_�mM���ȥ���XwRR���pS�e�%a����t�P�J�^s�i�L+
^�O��r��ᤛ�Ϻރ��}����ٞ$M2���:@ؕ �{ִ���S�����/���RP�<�P�P B�e��0ᤍ ,����x���VQ��D�<��hؓh{�&�Q�a~��I�*K��/�u�2t��c*J���0:�����u���~;�s�53��;�0�F0R]� �ff�kX%w�>���զf�i ��>�A��AH,ߺօ���_��RJ���޽^��u}�>f��~��m�*IP�/��Zb��ʫ7�r�̹��X�@��~ixKl�ed���:��>�>�:@�T
��K��u�CR
B�s�s@t�H�(.g���jG6�V-BJδ����[u� ��/��ZgL��d�X���撡+�/�|�M������+���H)8�d�~�i �tʐS�>扴�~���ZW/[`w�;�45?�%��[�$x<	�o7��X �<�4I �`�o�j@���ho�l�3uSm#b��MN8ݰ�z���I�4�[��zF�i�23��<|���#�&[yX�z�O��Vּ֘t0�-���n�r��ᤛ���oA�6�YY++պ�$�7d���+@�#�
&e�:k�H)����6n�Z��C�ϟ�^ C���>�!D\L������׷��%��u���ҹ�06����<M6�_d����Z�ZH,钡RT�}�i6��*Aa~�u��%�|�r�l;d�K�w�2t��FT
�9����5��6���S#���K���﷓]�o>֒
AN�
�w���h�d�9�|�:CbJ�P�י�7�Kg��G�zf�K�ӈ�p�����T����J��A���w�C��P*V���k�7ϼ�:����F�-�~}���n�[�y�5��u9	Dm$�@�>���l�T|!ν�ϭ�u�ACI*w�h�M��ay���I�*J�d�y���On�M�z��YP*T��D�m�wߞpn�ц�]��X_���C����m�>�u��^��@�U} 
M�
�+*}�~�Ci*%B���l�I�G��
�؋���ř���ӎ�U�!���gVb{�s�Ν�˩�⃧��z��ˮ�2�S����(M��=�7��sbG�~ɺ�b�^��qZ��jn�<�
�I~��+���8;�j�*P�jYY������M%��q��}'�1fIF�����k�L��emb���Y]0n��ge��<+������빳�=��n0/g��������?uN��/dx����;���{���H�5{|"������^;s���hyQ��\3��d��L���UT�D�7��O؉�u9+m\ԓW�8���L���Vթ��H�Ϊb��V-��O��jY�Y�͡�Q��y�,8����w���R��k$v��=��!c��Gϳ��
x⒅��_�ӚwtA+�^^�Al���8��X����UM�,�*S��=�;�m׀���ۡN���,��H�aÞ槽C�2������T���m�2mI���V�7';��6oX��[�a#�,~+��{�V���(k�ݑF k�Z�.�C�:���N�gMoz���w�?-#���!���+�d-d�lm����pf훙�1��HT�K�!�KJ[(��-,dZ���l��[mQ����-����%h�Ak*TDmP��)�Vʪ���1U1*,.4X����\���)X��UEX�c"Ĉ��(�X��Tq��EDR"DX�KJ�Ԩ,U"�bQ�D@QT\��(�0����b%�,EDW-F%kF�U�++��R�T���Ʋ�X��TTkR�X��X�YUQQ`�UU�����E!Z�Ҡ�PU
����P�V1D�QdTQ��Q�[h(�V�+��1�;�����f]6�ը'��N��Ӯli�tl��X5p�
�g���1��y�hV��T��]�ܸ��z�uN��sE�I��9�z5xāb��s�K8�Ђ�8��8���lZ��#�\c�Ǆd����p�������Y�-.ؓv��ؤ�ݧ�kmm�vB�1[iR]�[��{v��A�}�AB����n�=x�ȸq�)��l�����n-狣�&�]�ڍ$'�m�N��3��ֶlym
���!ݭ��6��4�`r�h�V�ʊ	qs�c#���7H�ń5� 7��mq���I7Ov�4����J�1�k3`EA/,L	A:ٓDMf���v�����69���sA�ܸu���pe�.fI�1�x���șF*ԔH1.�4�僸�Jg4�1v���Xk�r6
"ֈ[D����t�,kL1�\��d7X������$z�!p���7t.9z�� �'P��^݃q#�{��s'X��n�=뀝7u�MӶ�I�I�՟]���B�w�%)Ļv;[�x8���ֻ�m���֚]�f�+����V�Ü�� ��i������|�OlV�G;rpѹ���.�R�m�9��.�k�O	;4u���N�!vaY;$t�u���)�ǝ��S��0�C�C����6b�I�D�+yI��r����9u\��\�܂�����I�Z�f���5�G5v�3qsq�F-j�u�Һs.P5�M\�Ƀr��X�N��۝�bj�Lu��\[&	e%�ĺ�C+-0Gi��Nw��a��qO[t�a��BX�4X阶�ͱ.���.J2ʚ5 �Ѻ�
�d�;�-#e�j�XW����8�p<c�9���b�ڣ@m���	I狴+im��]�M
� ��f�Z�w=��u��z��V�+�������v�	���E�Y���^Ѷ�s]ˀq	D8bo;�=Š�@p�<��:����2����ѱ�H(J����g�IG�?�馌�u$x$�� ����Xs���t��.���:3Zmvl3�i�� ��gZ��gi�{ί��ֹ���%aF����C���b�����N�Y+*}o}��!L�Ǭ�>?��(m��Cρ����7�۴����~�z����R�T��\���|gZ��x�R*{�~�CbJ�P����L:aX/L�|\&�DBj�,�Y��
�ٲ
�Y:ea��6�P*V�;֘X�i���������vzA}���jM�T�7�e���j�Y���}��i�2VVJ�IS��jо�-�����}��>�w��}b%��/9޴��eH(%O��4M��z5S�-�ϨkF�����pk��tF��'/%4�������K��̧��I���=纇I!��~w�=0*AK*S�y΀�n Vn���4un���;�:Cԕ
$�X�����0�,����s.ַ$�B�5��L�Y��uU����Nd9�[�N�L�4�+*ݐE3���M��+g�l#=��3�٫��T��S}Y����޳��ƌ�J�D��w�$CR
>�>`
�<	@�gz~���u,V �����7�G�2��Zr���2\׺�:++%B����sF�m �!�{r�w���k�\/�/�	A�F��P:J���6&�_y�wZ�:�ƭ��/����&��ף����ȏ�/�֞�k��|�@t�Y�Jʟs�5��^��gz���*ay��>T|��:��9�fIe|�_ Q_���Cl�����=�<Ѱf�:�~��z��BV�=֘F�����h���
؇���Ci>4{o^e�޻���v����-nxi-@I궚�10Ū:��LEw��v�1ᚭ�p���z�82T��IS߽�@t�ĕ ��9�Ci6!Rg}�u;�4�y���N�����*Vg�z�E �7>eAh��Y�Q����Dx$���99}�c|�ۃ'�V�
�S�y��7+(�X}�|�:CbJ�IP���y���ߝy�a�°w�}��̸kZ�I�!S﷽�6�YRy�63h*JħN���{w3��-��Y[
�l��5�{a���{l3�ܜs��"V�꨼��۔(J�Y�إ3M�a��\��H)�s@t�]�+b��V/�*�~$r6L��x�问O��湉�_grx̌�T���i6�XQ�a�;�P�&Щ*��ε����_<׾g��`ʐS��扱6���l�ִf������X}�7�۴�������ZǦ_]���ջ��������H,�%a�;���*$�Q�3�kt°�]L������7M�r����<��=�����f�m6����}���&2���O
^��A�6�Y++y�4m�H(+��k5�������v��ӯ���ٺAl`V�{���6��<���s��n�����s�c:++%C�<��]����i3��G�6�IXV�����H)6!Y('3�k='Ȁ>�ڻ�?poB"f��w���_<ϋ���Y�}�;�9�4v���)l/�k�k�*=�u���<i�e+(����� �9yֱ �{��]8���H)�r�7��������"<	�����P�iP*V<�z�5�cRF��0GL�}3IM]�_+x
"�Ѡ$������^��������V��뫜�31�٬�������~>@w��(� B�8|`�nA��a�3^k:d�T�<��h�M���j�����aX\׿u�� �X��k:eH(J�w�4L��/����g�^�E��1qt�[Y^�\�c���v�h6u��S�a��?3�>(�G}L
��J���=��X�R
t�S����@>�ձ������R���J��%�
0�s�bAaֺ��˫��5�p�<		�� I��#�R��^���[�>9捌��T���k5 �	!��� U!�J����B]���9�v��
��]߫���V�6�d�}� ����RT����bM�RT��/�x>�s���z��T�
���ֱ��VJ2�T��|扸�`o�|ϋ��ÈSDx��_�6r�S�\@zȆ�!K`uw�� �FH)��@tE G�����ׯcg]fR��I��*0�}� ����>�n��ֳp�AO���m���X�þw��Hl���c�G� >����$��S���@nn�Z0+D9��+�(��׵��u%���V�Vd������&x������p�0���-���Yq�|T]IKb��Rϋ�à����/!. �	Mjpq�+�v�$�zb��u���鎸�v�K�x׮�ǥ�U;�v�+�o��>9�J�O0�]��a�V�1;eX[,3���:�^�ϞY�qZ��ۥ��`Ŏ�����7/.��I�t��D�HiVmu��˓@�![��.��e^C�}��\Y�O��N�vt��틡�7n�k^����e��s��.g���+(�P�*y��h�I���Xs���t�hT��Y�|�f��z���T��R
u��h�����6n�f��� �����
C�s}�P5��U�Z0*T
��9΀�Af�%Ns�zدy�S�bW�F�a��p�qE?�� ��9� ���T�v�O��$wvH�oV1jU�X��p/�,�4����׭Р_^����2��YT��7<L�B�����A��!s�$�Gu��B�#�*��l"�̓r�D�q��;㞡g=Le%�ƴCZ�`��^���I����Ձ�~�t�*��_jno'�[��.�u	}#G	��A���>�N��)��M�Eg��|����p�[�x���Ǻ&�%.���4�xn*1W�=����]cܾ��N\�N�3䰊�٤����*�Z�r����4G���wC!d�sw�q˞Z��}T!wK����9�-��;�d+Y�]T$�,h�	 ��/L���Y5���R�bZ�*�ӃH ��<���[�*��l��{�kꝝ+Պ=^&��a�<�7Sюz�azt��M��k{Mk�R�v�T۩��,t�|�����Ž���$���o�@���cf��S	��:_���ۼ.�}��je�v�L�F�t��؜�,`�!4��*",����T|t�n��빯>��X#u9�'!߫X{X"��TsMﲛEN��T�ᵼ�ej���@����;�U��Q�_p�������>�UT7�&��O���`����]�i�6�����n�Y#�2��h�J�Gy�k=آK�~� �g�M���$�����ѵW�|H)��1���ԙ���m��"�Wc��Lm�16�秅[�n�G
زϺ�f|F�ɐ��^�]GMc���4-��[��(�i��.��T��g%�v!3��7{���Ǉ�O�c��J���X��!2!72�'�y�j�ٽ�`�tk|�mR��{T>�C� �J̐��|�{���&���'�y2�vEcW�_t�d�з;JMZ!SE��n��6rl��,�}e�[C.k1D��:���%�t.���]zIQ72|��JL�d
�w$�ܙ^��'����:������cH��=*�V�B�Y(��A��D�K4�z���R;CFfT���������+z�H'���H$��)���c�O�}\�dQJ�P$2�p'��e�B��*��4�c�$��Gk���z~!\S��9cU���l]�B���R۞� ��&���`:z3}�W[��=�I {��^�S�&D&�p�}�J��)~��Ζ4��ݎ��Α���$:�'H�[& ���&���=y	��7�H�w"|M�2�����2���
/�h�u�L�t��tz��ҥ�岯1��Y��4�3د/%��˦	���cҡqQ]���R�I��Ya-��"�އ�J��sO8Sm��{;p��l[�����X�J�ŏ<ナ��hN;:��Rє�8�zz,9�qqn�]&zx�fų��q�Tvn{�쓊��Kl�YHJ��S�Bn��[�2G����<\m͛Y:��ϭ��e�=tY��n7M��u�/h�{8^��za�,C��H�uT��&��w9�0�����SlI#�C���m�)�v������:���7J�{��>F���H�Ux깡�V��ƨ�`Ɯʥ�80u�U�W�}����|�, #}��V�r �s1v���#
��˚�2���+��*��]����UE��!?!2!73_/�@9�[��S�L�GdP���Pz{j�7��|�?o�"��Lj���EX��1M����c@��{�(�7���{q�>Ƶ�#��E�"���I��	���@��{g�m9�1�Tf��u��J[���{�sQ�1�r{f��qr��7�f�X���+�L�_w5�q{����Tܗˉ+��h����M�S��v:�}q�2	�1�|*��'�_v�r�xMCX�,'}�sM��t�[�@��wT -��*A�t��;�k������T����A04�b�^���ѫ��Ӄ0_�r�H��b|	�����&���[�{kBw���5�5Z��&��<�l�"���˦�n����Ȅ��"-�=;�@ މ,�csn��K��׀���x�J3%����~�튟]gԏ�'z�>A�|'�t^�K�����]2%�sF�UP��(���]�8�~���U����D1l)���Cyo[�nл�!�L����Ӧ`9�+�����D�
{���#�^�����rhs�j�3e�Q�4[���v�_���1�=�Oq~n��r{O�!K��}�@ٽ)��a�#w�L5�D�Z#	�����7h�ڽc.3,���Z�Trj�e�ؤ1��m�N���S3e�s�x�����W�gx_2T��'=gy�דs��;����ya���N�˽���s�gv����\�=Ƈ��8���b�G�g�n>�$F�¯k���U�!?��]}�g�{�a�zJ:�-��Y�U�����8��!YÅ����M�".k7l���V��J�/c��[�j-��v���˞�:�`�je3=<>��}�Iι� ��	A�b���9��^�ջ#/�aNf�i��~��s�Y=-�:�ީ��%��_D�������U��Gy�'�坞s�w3����P흷F�Y�H;�wq�D�1�;%Ȟ�=[��w{����B���5�y�Uk7qJ{��dU$1C�3z�ړ�ö�d����G��e���z)1ѭ�s|eE]�K�{t�=׬M(;����oq��8�ӻ�yܵ�!�0��t�U�=�X����b� �+UEE`V�)Q�QX��EQQTX1��Ĩ�¤Fұ����Vf4b"��
�H�T�P@D3.*(�h�Ee���*�DU�V+P*���Q�-h�b�H�Y[TcmEDAX���EX��"�"�b��[J�UQUb#"���#*�"(�EAQUF*�V*,���b���*�&4QQ���1DE���X��Eb���*ZJ�Q��"�*)QDb��U �����""���F1VEQcTU�b���˞o^pEG��~�Ŀj���
a�V�����-����ېI�RCww,�2�Z�:�:�-�򈦆5U-����__7�����c.���lI`Nwt��|�J���V$U� �b"J�B� ��������t�r�c�i��%E�p(�h���U�O�ԗ�A>'��_�3��P�C�B|�Ȅ�̕�fI�[��Q�Q]"H��_�����RR�������>��#I"%�d��� ]���J�.�z���{x�"�(7��U�葑,C��;*�L*�f��7��<0���=9����{�朗.��t
�ِ��jd�߼���P3;˖o1z�O����c�:��
�E�����:�aW�]��p[`�m9$z�dv�koc_Y��S3c@/^���}T��E�{����n���p�!y;���G�ֺA�<9�����j�Q���wt��^�Ϊ�g;7R�0������̝%(p��S@��I"�+r��RpH7ٯ�|��2&�,�FX�|�M̮���T�!r䬪���7����y�]�U@��H�H�h�.�gG����⯲��|#W�"I�:V	p��'����u�@`�DO��s$;�f��i�������I�bI�E���78�'5���n��-䱧���l���5�����x��zj���'"X��RG����|֨ �j�F5$���)M��!�LHb¡K+�\Ԗ�ƦԮ5�#UX$��'𳮧Uta#5s	��T�ƺD�	�Iʮ�1�����3).҄ �����Q��]��z�7$:��r��ڳډ�C��تJp*be�H��O)��#u=�u�i 5ef��1�y��%�N�ȗc\� ���<�׷qa�O�^�[M��I���ˤM�����FWU {=2Aʈ}�������KV�	��B{��g���ul�K+D�I����>$wEH9�ɜ7x�;��wĈ�1f.��ڡȼ�$��<�3�w��n���lhW������[��]3�:lB�믕�2lh]�Z�D̊Q�Z��#�"%�d����g��k{ۓڦ9�P�b�+}�[<j�;�:��(���P�d���.Nn�{Q�{p8��CA��'�%4L���7΅ދ�WwL�heIӛc;n�ӷ_�<˂����.;����謀�7�x�R�QT�z:�F�v�=���w�F�+����b�a�5�,9�Ӈh���8���yR>��cH>���|��s��ՕB�L�
a��I�=�g���O������{ѻ[B3��|��_QKw8"%���Tv;/�k#lX� �kK$�r���_v7���l`��������}T�}��z�cv;t֫,����u���-��aW�(ج��sS:���\F���mB�c`t"����:`��=X>��r"���#�f��l�+��364 u�]E�>q)�feGNe-N�f��OWDP� �nO���r$���4:M\K�T:�a�9Wd?y�=��@�œ�]�ת4���E��=��53ݸ��]�˜�q��)J�/>}��e��`�u,��E�3�.j�Z��[�8$voR����>��aL0�	4;��t�5z�2��=uT|;:�t�Y�U���W�_&�&�U��$�d,�|����q76� ��׀|?~4gYMQ̬�vn�I"�m�ڰ4%����Sd���\��Jk��|��e��l��s<sڪB3�t�wN"}@��z�g���R:aDKD�V�gF���L;�C�ֹ���Ăw��!P�w)_v[66���&fp�x����FG�'��g����@�:�;�ج ���7�z�49N�{��I$ի/ĂNm���d�Y�����k���oDeU�n�ۥJLî���,���%=��ꏑ��� ����ϰ�0�E8;b� ���30ĩ��B�����,�;��K�j�_&/�:&�b\n*���R�k����d��AF���J5���o��C9~�㱹25j�$��|�\_<3p�.������~����3H��t���U���	$��m��+���t>�#��U�΍3�ΐ�f�*v:"��a>7j�$�|�*��>��33I�3�E������>aY�T �[�&��v�d5��)I��!þXa��ت+gdI �w:�jGF�,�{U�'S#�͑ �EwT�S}R;���[~B_,G͏7����->K�>.1zv�'�.���}��&ě���w�ߔf�\�}���Zs.4�]�UZ9�e�X�F�/cI�S]üF�!��.n׷l6�LY%�w�'�ݮ��i�q��^�s͎�Ƶ��	��N��۴�B�	㍣��y:n��i��Yb�x�;Yٍq�H1���L�;<��]96�=t��g���YZ�y�n�l\i��A�۾|mͭ��W
`ч�Z��v�X�JgmA�w�|<����4�������j�+�H�I�;Ǧ�L�Yg�{�g1V�	�E]y$�-yeX����vz�/�o�=Nf=�ܔ���v�5L9�zz��?mң�G߷��!<��F_����t	��#�
�Us�v�ò���;YT�t�:Gz���[2:��9�1<O�:{�!�*��i|���������w��E��fd��kv6������`N�CGKH��2��|����MT�/�zd�w:��yYe�ST�]Zt�_S�mұ&�N�E�I�yq���P�5��D�s�6�:]��d�)�m�"�PT�5s�p���wZor��H?v%�\:����
g6o��n���w��"wios&��E���U�Æ��#�^zA�Y+����1�g����mH�w��f��R�@��r�<��*>w���0b޾�c��k:	s�Ļ�!�Pj�#�/o�өTjz$mv� ��X$�ogUV굜��V*F���#�m�����VY;u���M׮�lb�J�w�n�������[{��0;��ڧ���y� W��A/�1@a��ؠy�H�컫��=MF\��E�A=�� ����ͫ�5{!d���/�Ğ��	��ɝWS��*�s�褢]�e�q0��waį�g���OD#�$Z�������z�Es�1�fٗ~�Tt|{o�g1W�m�*$j�5Tl����@e�.���W�8��s]��SVC0��A~��r�rIv�}G�����=�fΌ��������ﮓ�<�ǯ�j�;h8�k-nX���s��j@�z�ix�Su׃�!
1RXGo/�|EoS���}_ߢ� ��͘}CAZF���yT|l#'1��t`�_wU!�u@Fcj�sˋ�D�\���ڭ#�����t	_'��<�X��E^�)Ʒ�ɋ�b0��r��#u�H��l� �ީ�F�Wa��S&\�M4��]��ˁXȺ�U'�x���-cȼ($��vwO��u~u�ޡ��Btf&����E��m�����]�,����bJzw˷�� ��e�T���Ȝ�#5�4J1���J<_�D���5N"l)�0͖fb	�9i�;�G���p�T[|�H|���:f�1�WvU ��t��0�En� ��*�5�@�S��d�E�L��#WZ�{�jw2���H�yQ3��D��s �=k̾�q�}�&&�+�S�G��d��D��mR;�����!���i�>���:��Ӥ�|�]L�F�L0����L�:�^��2A�Θ�$8��8��������?h?��~�S�ҵUU �BI	!�?���	$$��l�zHI!$8	����/x3
�;�Ο��n�5ўxS�ɦ�c;�0`�HIа>���%��,�A��_h����$��٦������:�:�N�'!��<����î�f��A��_��e�]?�o�����4�O�l�~�	$$��r}������������$�C����CI!$?��氋&��?�:?���?��ԟ�&	�?���~����~��)�����BHy��+����*:&w��~��LCfJu������$��������r!����_�����G���:o�����BH>i���׺����d����HI�*�y�)���0.g��Ga�gD�>�h����C�&����$���?Q���"L����Y�d�?؇��O��=I?��N��?���)����I���I�~�e$$����	�O��������@�iї����g��P�'������~s���$��������$��_�������0��C�C������P���9�	��y��PO�܈��$����$$�����"D��_���hY?f�O�_�A�����)	��@��� Hnl��Tc�0P�����I2ud��@?a�fà5�����R���r���&�O�`��f����`�u$$����?O�����$���a���#�O�����S�߄?��������C���L!?���\�?�����?>4�8�( ���3����<�����$�����_�B/�����D!$����#A����?ԟ�{���🄟�L�Gru��I�'�"Le������Ǿ!���P���_����7<�?#��_�uI!$?3��5���~��?������;�?C�!�ߔ�_����Y�jIC�a������BH�$�ߟ�?�������Q���ߌ��BH~�?a����sa��u&î�ad�I�yg��tO�E$��'�e ����Z����)�(Y h