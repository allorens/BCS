BZh91AY&SY�HW�<_�`q���"� ����bH7�               �T��*yĂ�R�[5�Q)
 UJ	UBP�
D)V���$����*66Հ%%A%	Ta�l���B���*��F�$R���*T�ѭI�vt4QM`����� J�IKf�)B���/�UHU%:�*�P|�%5��Z;f��\� u@D�R��� j�nځ�N �HJT� �H��Kl��PR�P`�6�(�ׯ/P
�R�zm�P��{۶|{�rs��vͩ�׸my�wl�k�uە����s�.�K��wj.���p�Gnܚv���h���'�ҕM����w�u�k��^�A��4�Uj+Y)���Ҥ�P;�󭬐:ν�z��QL�"���)_CA��y�-
�
y^㦯5kN����𤊒��u
Sv�uF�ڭU����ʛ�t��(Upv4E�I�hkm���K�*T�(x��t��i^��z v�U3ǼD�%���x�{۪�\�ٽ�|�
;j����MB#�#���}U)R�����5	^�m��ޅ�W�G��W��PqT���mT��7ϥ%J��|�
��/;I
�m�u��>��|�[}x}}R�E�-��z(��Q_i�|���`�>�痪����y���(��/}}�U�)l5��ww��k#�*Wm�)kP5aa����|�R�J ����@L�Ϯ���������7���yw�P�j��ky=։U�wg�ת�m<g}�Ί��+�S�{� U��|��W�}9�y�T�n���B��s�v�'Ϥ��� ݾ��=���{'�z���ں�}<Z1���=�������z�p 9`�����;�yX]����9P�%Q^Ҍ�ڃFCO���)@�� Q�I���t��ݍ����G �a� :Ƿ  w�o`�^� ��p�;�]��2�5J�E�G|�)J)@���}�������4;��p�E�`t �m :k�8 f�w@=�nѠ�e¨��U
�J�#(@Jla�Wϕ)%(y�� 9w  滃�@m;�A�Ms� 8�ۀ nk`u��0��v��q�Gr�u�k���d'^����m��JR� ��Z>�4��;`�vY� �\;�4>�����GG@�À8P�l��;�P x          jz Ҕ�F� i�`L&)�IJ����      jy2
JUi�р� LF&�jxBi)*��C0�ɐ�JD�UOH 2h    D��zRHLD�2OHm� 1O������������G���'?���k��5ڈ�To�!E�K�절*�\��"(*�TEO�PPU�_�4	�_���KT��� ��U$�O��" ������ ^~���������08�����`[`[b[ػm��酰-�lK`[`X��%�-�l-���1����`[alm���m��酱�6��[al�-�������[cl�cl4���alal�F6���al-�l-�2�[�[�cl-���e����q������[�[��cl-�`[cl�-���:e��6�lclm���q����clm����0�6��m�l-���6Ì����alm���l-���alm�����lcalm�l-���6�e��6��񅱶6�L�6��cl-���6�����������S)����clm���6��m���alm��-����2�[�[cl-���:m��lv���alall$%�-������cl-���-����[alal�-���Ķ6��[f�[al6���cl-����������[`[4�alm��[clm���[#�l�m���6����i���[�-����l-���alm���6��[al�clt��[cl-���F���clm����4��[a�6��[`[8�E1�6��[alm���6���0�6���a�[cl-��-�����ۦ�ala�6���a��m���alm����6հ-�������[�֘[��Ìm�����S-���6ǌ-���e��6�lm������m��-������aM��cl8���`[���1������m1��-���6������-�`��#� FlA��-���`�F؋lQ��"[m��b�أl�"�m�� �-���� [�lQ����[b��F�+lU�"�m�6�M0��m�;b��F�#lE��-��#m���Kb��Fأl�(�m��hR�l�m���[`�VأlA�-��#l� � m���؉l�;`� �"��ةl�� m�6�c��m�6�K`�lP� �m�6�`<b��J`�FةlU�*[ m���b�1-���b-�S���m��e�F�#l�m�6�b��)l-������#lA� �m�6�`0-�6�Kb���
� m�6�b-�R��lT� �m���b��B؁l�؉l�*�6�K`%��+lE�#lB1R�lA� �m�6�Kb%�؉�-��)lD� m�6�`lA�
[ m��l�
� m���K`���lA� � m�Ō� �m���b�F�+l�� �-���LU� �m�6�Kb-�Bر���[`��؃lQ� �-���1m�6�`�)l� � m�6�0Kb%0Fةl�(� m���b�R�)�6�`�Sl�"�m�6�`���l�
�m���b��F؋lA�;b%�أ�*[m�6�b�Fإ�X�`-��lQ��-�6�[`���ؠS`��lA� ����
�t�`-�V؋lA�� -�� ��l�
�m��Vح0B؋l -����D-����*�`�l-���[�A�
�m����l�(�i��b�l -��b-�؃lLP� �b.�%��%��e��:alm���Ì�1��-���6��[alalm�lm��clm���8���cl�clt��%�-�lv�cl0�6������F����6�����ݴ��`[clco-�1�6������1����clclm���m6��alm�l-�lm��0�6��6Ķ��d`[�`[al-��l-���6Ķ�0�6�����`[c��Kcl�-���ͱ�6�L-�lm�l6���1�6����q���[�[alalm�M��cl0-��-���m%�t���-��-�cli������-��2����c�6���1��-���`[al8�cLm�lKcl-�[�[`[���-�LK`[clm�al
alm��-�lm��0�����[���i-���[���[m�0-�lalm�������clm��-���6��l#����MĶ��Ìcl`�lcl4���`m���6���i�4�������������lm���m6��:clclm��lc��-��-�l�`S�����m��6Ķ�-�l�a~ �0?�����D�/0�O�M�j���5n��(�iZ�+��6�+�� ��wI�G^��Yܺ�qz��7&��[	H&��Y�T�\(��Q#Eۇ7�<l�f]��+#i�ܤdy���|`z\�VJ�R���Mh�e[�d9���[�'J�]yv�'m�t��̎�{����A�I�$��pe��.7�����sh��G*[�w�iqn3SV�%��״�q�-�CR��Dfٓ/Bj�=
�s,t1���VMy��XYQT�6]-P����f ���XL�0h�b��N�]�LG5�D�dFP�ܴ�T���G5ǩ%gs�յØ�@�
�\Ԛ7mmڱ{-�iא8��2�H p��[7"ܤsNG �W��M�:7: ��b)Nd�inr�,.n���
7ró/h1�QڄͤqM���
(�[ër�h!�)u�Jr�'vI#SGm
�m��Za�b�_f+�iS)��x6�rfn;y�m���*���(��^2�n�ڻ���BqF5�vHV��[�+EP�CS
ejא-�t��	ӷmJ��ubP75f*i8v��	�%4I���5��%phy�C�J�tӻT3Ee16=cpX�D�#��{F��6@ݷ%b�@���j��n�0����q��c	f�R�]&�'f��1L�xj��`ٕa)��-l�Q�Uرb�U�2cv�\�g%�	}Pؤ�]�A��u�����*������H�9NoS��ּ��ن�V�ߞ��*�n+Q2a)`�r!�n)�=�nm�a�E*y��<���b+�^P9.�Cφ:�y:\q͎�ܔ��pe������kB�/KC�1
LnkxļTHd��j:ͭy67�ޕ��""ՂX�)4��{,��]����+d˳�MY�R&�J��/�L[��(S��v�lԏ����ъ�2�n5Oe�K�WV*85�p\��0d�m�Tb&�f�vNP/
��4N=�)e��'[FMy(��fI\Amðث�.�(�%UՕ3��b�m�qԻ���YL^�%&I�mov1`fꪽ����b3u�<`��*v���ViX2�"��Ck��R��ʎ��Ǻ2=���b��v�[Rε�4�l�V�W��Xͩa��#z���Bڱ&GIc{��Y�J�Q�x��F�"W�n�S���Y��%�����KԢǻ�����@Cm,��,;[ig�����0�#�إa\85k�^&ױ�73o�ER�%�9%�nia�/`��t���n�#�ۻ3M�E�1��
m�=��Zr�e�p%�a�����深���T��raѢ�6M�wxaN�fYlÊ�o�X����W�mY
�{���qGy�]K9�n&��T��(�v���2%��Vu�7��S+��@���u&"�Vn�kF9��X��w��̖�m]1QV+3/a#��Ӹ�AUb��Z:�uDt�MV�m<�%mf�a @Syl�a(��e���ٕ���J�Ж��;o��	����R�n�u�䨘1�A��ʨ ��&�֣r9rkǘ�<�(��4��X��m,���e��֜b��ˠ^� ̸!hRIUo/s�M�<��Y��)-��F�CA�Yi^�"P:Nl	�hԱ��j䠶�zTn����׌�����(��U)!#���܁0��� iE��e��A+r�"��Q,�W�j��%DZ�w@9�.fꥴ�l�r�7��\t�;H�sA;��͉�r�%d� Lcqi;	R�(���(@�,Q= �Q�U�J���F;ګ�21�Ό����B�#�"��Iy+i:ŗ��W���0�z�&S�'�����R��e�^<��0'Y��MY&kX�%��u�ml�hmO��V-m���f���d�'�K!���s3I�HsY4pKq� ?Zӹ��d��Ѭ��À���q������V�0��V0k]�����:L�U%�>�owu�[����,U�wZ�*0���$��sr�Ђnѽ�����!0���;���eT�md�̻7u��IR,����p��fm=�h�g	��6-���q������!ס!��1*�m��V&�X)n�i<����-�sD��SI��a4��J@ ����n�+>�Y��rLv���T�YR(M��o+��y���Kxr̺�z��BԴ)���X��i:����p�N���%<�]ܷ��V���^9wt��-7#��b�6eJ��2(n�W�]�z�����z���Jw��;vE�.kQ������'v
�4�}ou��ի�����5�X�m��Xβ�!����r����7��
D[B͈��r���?hʀ��Y�`�^d�VqU�7&�\Peo$�ڲ� 6ޜ��1�%��*n�n�ǘ�oED��ݥbcys�v
�t�,���yXt&ނ��KV�ա4ȉ�{�@�S�1,9���o,K!YaO���*�f��a��r�Ĭ��3њ�ɖ Ь#�`�w��Ƭ+��\�۟d0aۘ&��t�H�h�WH���`m=��b�ƪaf;;Jă6�C[k)�b\�w#P]
!�����W��fkЄ��n�	��T�;P��سi �Udڪj�~j�p߶�$�9��'���FR�wi$�!5��̪�Okҵ�5 �D�����RB��Uw1fee�{~u�^���̽����,`�4(#�����x���@- �C4�u3cӡ��,C,X7�V[/5�r$�8�d�ef�A0�2;K��\s~D�l���ټ!;Q�#�+c�@˖$�>#��9��M��1yòb����6c��0nX�����aW�հ�p;{�tP�w��JKj�c5�Ũ��Tˆ���֎x
��h�5�*����&�����+w�Tj��>[[��u�P9�]Ś&ݘj�۸��n�ف�0�[/eh�RV��Q���������%Ս�L�o6���H�]7�1a�W�t�N�+ť��G7Ɋ���ɛ����g��^�d�=�d]�2�u��)R��Sp(��rPv7.�K%��dJ���ތ�D:B�C$YfM�&0��krF����W�v��;"2j�n\��YcNv��sʕ��
�n���ƗYv�d�%*c�uc5ԺB�;aÐ�B�1wwP�3b�i-k,X�Df��lm�/B ^�5&��BB
����3BV�4�҉ڹ;vi�a9��c�����)+�-@˼�"����<x�]���"�Zdz15�2s,���j��
��,��f���A
�NV�Q){$V�9HT$�&�5 B�,���S/ņn����fQ�]7�ˡ+-vZRhn;�ha�3h����ݭ1Z�ܚA�y�9!���p���E�<�
�q�G1G4i֍A��t�䘽�4�R��m��eg��9mH�̻Y<�`�y��ceZ#´��R=���X��{{�G�e�wN��Ő�A\Yo+q��jve$�S��&�j����p+2V,ǡ;:j��8�y,`z1��NF�U�,n6؏j����rM%�FYZ�Cz���[������Xκ6�H%%h�Ǹ���
��i���f�b���G[m�)a��	+�5+�� ��a(�e�v��vU��]m
���'�^"4L���#Eŭ�	\A�װf�t ��a��y��V�\�P�Os-гͱ�����l��ˎ�;m-�" n<�PU廕�����)���ۊup1W1��sm�I�Ǘڢ��q�F�*h����i�"h��V��c�7&�ȯ-�������*n�I[�¼�l�ܳ�lQ=J�)��Ii:�i;�C�)��e;n�P��%"�vn�w�44Aw�Bjaq!�3�Y������%��]�Y""!��	s/�U=WwT������87��2Tݪ���hХlᲖ�U2��%�	���:�id��������;QL��b��Mų/E��6ĺ?"y����-&�D��anǰ����ܖ�[m��2Vc�E+�3��<��!��f)D�j��z��zf
f<�ڟY�7N�m+���Y��I����f
b$�n��n�i��������P�v�Ր�)*zwT�fm�YW��ҭ�w�oj$�%�K$�fǘ�k\�m�Ԙ����ݑ-��b`��rմ�r������0�a��.�[�N�%���}xr�Pm^�sUn���U�%J(���Abf���F��w��6��^:n1uuH:�T!�Ъ�{t�-֤��:�xS!`ː<��)�y�c�o�ڻ�dQ��s���-�W��lH�H�A(�v�LaP�Q.]�CH�u���ˬDȭnms^5X���d�%�L�6�Ux����� �`�5V�F(ZN"��A0��'��p���;vŗ�ܺyK3E3����B��o(I�&^c6l6���Y�"+���b!��F�1 F�vE����B典N���RnP��.K
I�n��lٷ���1���n�)�7J�iXoP�q�n=�6�d�Yq�a,�ӹ��a�pj���-�N�I�E�M
)��:YTCJ���f�*�Q���+�[�����wF����[ͦ���d&�̊��1U����`�D�[P�8��;N�Ӻ�9��!��$�[0��`&�n�7%Ǻ�ov��������z�f�B�޵��w�K/H�-��F�b)iۺZ�bw�4���<9%��q�0U���X�#0���W�b�V#�oI1i�J6��F�R��{V�f1i<6ÁX�2)y�=�l	"�n���R�b/h݄�Ye�;P�8�a��ʘ��g5��8kh���د4{YjPƶ��A��M%M�ou�m�o^ٵ{��2��x�=�*@l�� ^��T��.���֥�Ѝ��^����,��c�-ñ�e���+)�����O �N<���T;�h�� ��0]d"��ĳүL���K�彎�la�:�KI�xv^�C6��ƣZb�`:��Q�1�V�敱��%��u-�Z.-����ԏo̓�����Hm�G4�����;�)�T�F�=��2���Fj�)�T�%䪱�^�ܛ��^��Am+���*�� ��,��e�1���d�)Z���M^;�3ˠ]��w˺S�YWz�Ԕ$(5'�k�&�&��.ZVf}�܊^�wSoUm�l�9�6�j�N��
ں�1�R#�f�Ɍ�t#Bz`��˺'JJ�g̎E�%Yt1S�h��X)	�k>��н��tLZ��V�
و��c�]V���G��x���혘+v�EDe,�
��h�6�K�yxgo��$]�&�^�T�9;+)���˅�b7o�K1Xe�jmGr��8BUS�w�eT�OjH;�V����ƣ&a4#�W["GL�1�X,^sӋ���n\7���ŧдgj���W��XR�.�޶N�׹����r^�fSOe]���+�V�<�rM:R�I�4֚��M��Wt�$��oR��u�w�&�����@s9]�f�6�VO������2/�ޣ�j�Q&͍71ՄއՏE�����[DPګG�o5u�{V��WGi\�DV���B��pK�Gp6\�)25��m���<��Eou�X7�&���R7}�Z��)V;��3��^�{,�~����I��K(m�-^\�ۼݜM�@0T���z8J�!i�K��!�K�����uUՖ�0��	��<��)+:�s6��*E]qf@]�]u3��1�I���fOg�,�o�����R\��n�d��Q�e>g��κ��!:��Pc;�X�v8�Н���y�a!�U�];3@�H�M�f�-h�����u��w��˶��Ѻ6Cp����s"��H>�n�u�Y�ҙ�����'aY����Vv�r�q��}lwr�]������������ޠ��L�I)���zt]�feөeuh~�r��o���e�2��wمm�м�y��zX��@�{�۩.�8w{�w;�B6H�AG0]ǔW�Q� ��w\��%r�Ձ�+8�q����f�ȭa�+�w�!iST����i]�����@��y���BkT���n����!	T��[V�U�jᘆM�Y&I�j�,�y�����	Oj��t(n���Tk�&%N�G�~m�÷\��]0�W�w���&��l޼l��ĵ�����O(x�k�Bp���P�a[r�Wɰ�]�jge��,�v&���V�K�K�Q&�Z�ܡ���SvDM�m-/��ps��%��g"��M�J�7i�*!FGHȖD���!f�R������0�1>�Qkb�ʾ�F��Pe�n�,�ES%�>L�Ա]�H�BIT���p��w�Cb��s*��Go��}�0�����vv�a0Y�jJi �[��X�	I$�I[�q�*K��Np�J7��d�����x�2����j����f���z�����7t=�?K6m/�ju�Oj�&X~֦��r��,Y�ڧrC�L�8�����Sz��;�n����tl_I��={I�[nj�ٸ���ƅ�au͗�ϟD�,��l>!��ٱ��@L-X����ac�����lEr
�)K�����g�o�t�Ĕo�����:z��w۰�4Ʊl�mc#-�.Y�n�M؃���t0� Q�o�-2(��_:7�٢μ��4��`�5%�Ə�ŧ������3zmwt�ӆ����]��+f�u�-��t��]���郞.&�n�"����D�-�&-+t:͇N	�P�0Z�{B���;�-����/b��]Յ��k�lt�ZQ�z�K�)Ɗ:25Sn��;N[_\=��}s�	���EQ0₈��f��]�xa=��#t�56R���%ݐŲ�iR"f���-7��-eM8Ŏ=�'C2a�4����ձ��X��y�9�f�4bfS�l\��P�U t�LU�I��śN�(��^����^_�^r#$gH)�Ev)L͛�.�����Z�r�L�A��Q�`�bb'fZ�f�1��P��R2���ߠ���#�}���µ�A*��c��S^�حټ��7�
ڻD��+��Y/�Tt��1��\j�gu�&U�[���AՉ$��/�����O���U�o`�����K��>����V�YSE�B�.d�[������)!���ӧ����݋U՗/;���Ó�G����~68ml���iv�|��)�+�\g����Y�R�"E�rQ�st_r]�}Kf�:=��2�[�c���G7�y,<���q�;Fd���ĵѧ�nheݖ��	�Λю����v���a��1s�'c���j���s���e)�|���}˥N(!�E	[�[?�{�54vQ��YC�%���N]�y&��x�h܅��ڐ����|����(+I�[��_u���F	����,[�)�.t���`�cS[%��n��b>���=��	Vi�ˮa����Bk��]�1R���/�u��e�;曾���3[�&ng%�	n&"�m��Xz3rF'�k^f	��N��hNv�����`_�xA��Ƿ0�D�:0e��r���N�����ncU�Fƨ�}�]l�NGJp� ��2<T����L����h�u�,]��z�vFJ�6�:�3 ƺ��y�w��D�1 �A;��{:./Dݚ�Ϯ�n!��r�U�z�\urG����Z��Y���2b}+6��bg0�1un����]5���w��|�6�i� 7@J3��wI��2K/켪�Eu㰦4(M��EC�P݆�<(_)�]����+i9ro*�e\�eL1OI@�}�-�|c��b�/�}����P�u���6����o��yV�f,g3N�	\���w,�Nq]ǒ|'u������[F�	�N2�0I}ۗi0ͻ��J�$Ŵ�Qv>�������ٷ]Lc]��&@L���6mc����Rھ7(�s/���tp�!�`�,d��1�N�Ek�/�]�6�����F���iE��׊���[����w[a˙m������Я���]�L�`���\i�|�p�F��ꂲt�򇴌��U�:��JI�����b�h���i��[m�յ94Ŭ�-Sx�Y�57+A�kٹ$t��f�����m��GC����g/�w�~�Wj�Z�xfFjSZ��N���;4��s̕!��gKb4�Kޝ�Gu��l���cB\��\^EǻO^]:7)����U-���Ex�n=Ý�#��q�pݰkOTwu1h-x�H�O�U]G�4${R�!�c;9�݌��+�.��(:��7�c���H��	��ս��}��ُ�O����,Xq�D�Ca�*�G�f��V�t(wv��q�3ZtI _NA*o6�n\)�L�c�)�{ǩ-�\#|��o%,R֔ᣎM��!H8��6Vk8�Ʈ�r�Ó*���Q�1��:�L���N�+׎��B��ٮ1��D��.�W8��cj{��S;��������x������17�uO�$��檤�=�Xڶ�5���܆%����*�*ۼ��˦D�H���*�&��yʴ��׵[�Q�ʛ�T�n�.T��u�=~j��$¬R��y8S�Z�����R�*��F`A8�!��d11���g4��`'�I����u�)����u9�n�e�����`������uq���u�A����T�8Օ�=|$&�f��5w��d��p5xU���f�;R3�M����+"sc�&��nU���QѸ��Hi�V��6U��s�e�Sج=��������wn:t
�N��ju����y:9���`���E����v)�}�}���R���hD�j��~��A��n�l�v[�n^T��,�_X��X;2��CCy��L��v�����ů���.��[�ĥI��2�N]%.�|:Y�o^Ut�%�QM�{�4��O�OY��]f�
l=���v8-�ў�WT+L�
�p��a�ZԼɘ�
� �؞@E��Y��qi���j�_>��}{C�gp7�Ωi�n��5�"8��Bq�k�P;w� �Q�F闝��VL̒W%�c$�G���z�̬�:���)`���V�7ٔ����x��މ��g� ���Sv�q�y۵���o��u�#CL�$�ۙ�I���!U��_j�:{�j��h��Qyemr��]]/SW{>2�G�͚�o�Zx��,*��h>p�6,Mf��,��U�q�]�]6ӯZ*eТ�)����Q��8����Op�F���z�sLN�Fc%�vcݾ���n�w�u3[e�����D�B]MGs"T��SI꺳�W;�-곣��lV�y{ԪgN�77(�럠�QC��=dMn��Z��NƯ#ә��eE�E�w��ʻ+Dv��j.V9ZДo;j)7��i[S�8�
�rI�ɂ�����+5�ע��1❮ބ���;K�D�X�c�@�u�+�^\a��U��wt[Q�2��3�ٓ��an��7��u޶����'U[ʶ�F��^�7��c]�[c8AN¥5t�lS��0�Qd�7�
)�����89��*���Wj�U�u6d�0u�����y*ʮ��W਻�<v��L6U"��1�%�vp�z�v�kd�b��,gF��k�^[����3�bjNW�:8�g5�ˮ�=��:�H<(V����<>���oKU�v�I��IPg��טK[j���6�Ɩ�S탮���v�o?<��pf<�Z
�fb�0_t.��@'D�4
����;}OK��\������+�]�8�ţ(i)T �QX�xu��]�Z�6�m	�]Ynƪ�0%�@��L3e�.W�A�4'}���ԗV�w\�dغv�\-ݳ��&��Y�$��>��:���
�S�:T�E���Ǥ�a]�<s���Vo_��7L����OV+�(�⡽sq�o`��aU���V��4u;�ޥ[i{�]���徖���P�-"q�2�w8M�@�M���l���v����#��>(}�ݑ�u1l�U�i�o2�g�m]Ň~GY�A���G^8�c�`�)*�\'l=�{[��j�����%��T8="m��.U6���Θx�Q���ȱo`',e�7t�8���f;�C��-���:Q��	t,R����U��3���QTt���̏�;x���s��u�v�)=�4��cj���I�&�
6.-B�E��|�8h���R�i����|���IA]�E�)<Lk�:�v*e8j�C��M�{3Ol�o�](H�Z��t�P9��5Y�y�Ї{�]����4&��'K�O2�q�ΦR@�k�������<�bl׍�vv1Z����GbEaI�)�{ae�tv��e�V�j��tv�b\zp5�A���C��N
�;��ƨ�:�f�OK�N��=S�ة������λkw7:��C�[�闲e�_Mz;�Z���6�wo�o�!:ͷ�H�J��9я�u �,<]�0��yp��}�*��[:�MҌ�e&�8el�W[xt�*��I#�����agn�nJzOa��rVݓ/�x�S���N9�d��N�ML��^�ױ���[�cGV��c�ҫemګ��=N�!�{�1ְ���\'c��6�4s�{�
:�s�1>]�Yv��6�{����י�t�+[%[�i�Mg��&�Ū2&��˺k��TZ��u�P������G���7NS���>={��:�A���Ŧ��J �Ҕ$�U"�}O-p���}�R���/=%Tp6����I�aT����~�ZF	t��K�|�߾Å���]�����tzب.�pwp��2�vV��|�h�6嶯*�S�s{f�w0x9��U��{2�֟�8�b��U�m\�;O=�GJ\�-5غ�MխJ���upY���O;+��ry2��]ܹ�-ѹ�u���-K*���.T�l���sQ/��2jfĘ�g�+#xvM0����X�IG�Jٕǥ\���f�Z�b�1�,��N�{��:P�]+��K��ʕ%r���#��Umm�WA�C:��׭���^3eu����^����,W�qeX�U�v��4�廖;�g��ۡX('��b�g�-shg:����@����J���U�s�v�%h�7X�Ir����H���ݐ⇕����:��}��<ÕXO��O���q.�J���Xuy��i��ρ��^S���9vY�u���ӹ&�5�Ǘ�*%�N2cSFS{u����Aͱ��V�	h��J۪��^L��VuUT�̸9	Y�/jј7zn�V��Z���NS�E�kS|�C^�2��d%mݚ���OlD�W���s8ˏE����Gי�eHY��G��Ut���x��[�:ݩLXل=��ʵ�V!�n����m��Rp��ܚa�s�}�J���,��FrF�UŉC9]���L�O@��oP�R��Z1�9-t�����v�Y&N�i�Ǫ��W��p}t�nk6��Ќ�������K�y[��[B��D����Xy8�F5b�;�5vGY��J��[���1%qw��\�R�%�YB=(�3�,"��ro�P��t�QչS\���o�bZ�+����!����	���<q�hO�2�>�����} �(s61���Y����ΝMN@��u㴝��G�զ���ūD'I��[�)��u6Q%U�6����6H85��j���%��gNN��Ggk�y�V�gf65Ǐ�
cM����DdR�欜v�h�TVeS:
�8p�bƬk2�u�΃�;�ס+���.9��PwU��i\w�����ͨ�f�c����6�JH�p�^�+�K�W1��$�t:w����rG��[6$�[X��b;W�[z��Z�YeN8�f� ]��L�ꝰml.����׿t�w�q���4^AP՞�M`V�Fp�W�sZ9Kh�! *�^���ڕP��*6�Q��֢5C;�)���C=}K6M�*
Wj�s�΢ܴ���V�SB4���,gu�IDE��D��R۹w-;�^R�XOW4{�I�MOa�wLtǇWvw�ː��U�=V@��L�ڲ�yY�n����R:g׶'�f��l���f��W7N��-�}�۰�-ܛ���F��۴������]�������޼��񨨠��1�9��" �^m#�A�o7�>��\�~w�<�ܰܺP�x��YL��4�rNW&0�9�;ǟ!9e�^�������л���]:��t�N�du��s3wX*���x;3w�_NRn����9�>= ۗ7�*����d��9����xj�V�ދx2��;���h����}�	��_oRA�9쬼�7a�.�z�A��Ϟ��Ƿ�E�@�IciΧj�T�<$7�uafR�>0KH���кY������M�>I5�H����Pa	$PX��Jp� `ĒQ�l�����Y�]_n��2�/R�d�ۥH�!a�ѐ>8�4(�����#J���Z�2(Cm�-8�0�"xx���y���uJ}��K�M�C����;�܋���1��=O$��m*4�C%V��A��U�0c�X� I�I6�NB2���HB�`���-�r���+[9�vU��Tr^VDnHm8���)�N@�`��C%�����HV��+v�QOB�,B���Q��$��T�7��Y�0�[�o��s�����SHYm7�D�`�LMR"��I�E�ܱwl���-�c����LQt�R�Ŗ��Ն)u'(�J��:dRH�!ۓ5=��Iz��l��و�},�O�,��]��DU:�l�$��
Qd1S�2�(BT�5x
�2���T"9�ȳV,�Srf�bs<�0�D(h]��X"v�6�� ��a4B#�AdG��eK�e��B<Ca�I�>a�E9Kbݨv���_�B�sC0Q�<�Z ����n���2lDa�D�8����
��1!�F�{J]X+�[S�p�.����cZ=�V��J�m��)��bN<����Eea<|jJc9wVȢ��m��!U]�፣v�T	-� c	�6a���;Hބ{�N=멈���h(!i��rf��	����u&�ҹ�[M�GQ4��E�hP���p��.�EoP� ��k���e�6�!�-� o�� ��Ż�t�!N�5��+���J(�ܐ2�q41�SR���	�*���p�osY=�r��+��@�&�M�N�S�'PlL��	����	�3�{�Fn}#��w���Ŏc��z�I��[J�$i��<e�Dc�Z;`�ׯ5�$n@!i�ɀ�0�a����ADD^+�^p�����a��1z���$�4[����h�KkjH��V�$PQY)�D��IFD�b�z�C�%��M@I�!I�B*GA�5Q�/��%���(�L�M#�CgUU6i Xz�U77�ޝh��T�_����`
�)�������X���"
*w�����:g����)S;�2:��&j�����إ�>aR��w� bg�Y}��ô�Zvo%p���Z�TdU��pQ\��7����6Yb���җڌFŚ�ͱ������s�-Ҏ���}�/�Et�;�ʲ敘je�x�����������Ʀ<����]. ,�L
��O:����/];�]0Y�[嶱_^u,���NmpK]a���5�0��5>���s�54�Bd⺄2uZ��6ku��O`�.p�K��e�{%+�����5��H�r�-�r�����&.�K��.�q��W5B��'>"���y%O��"ˎ�e�����8��D\��(��&��p��o+i�6���Ֆ����V^r/��������6�[Ш�y�9Kb-
��6z�P�D��B(�
@ɲ�9����`��ʃ�8�+	�Y<r���Tk�u;�4;��X�u�Q[P7�pi��y��J���l[��"y��!���4oѲ�LV{����X���������ت�FQ�x��GY�\d�����og9v@��mLV��	�[��I��T�gO	ET5Gd������s�6	�⊯��4���g������������:q�q��q�8�8㏮8�8�8��8�q��m�q�q�8�8��q�n8�M4�8��8�8㍸㎜q�q�8�q���8��qӎ8�6�q�q�q�8�8��qǌqƜq�q��q�}m��������m�t�{�^�w�ݓ��"���O�vXW�a��c��H�@���{�ܤ�Rnk�Ε�.����� �U���Y�ˋ�#��W9w}s�B]m�δ�"��5�{�Q�(`�hlu7]�e��ASv�*Iו�)�a��2z���I���[:I�k����V;c~U�U]۹F'�lT��8ž���Kՙ�線�Q�oU�f�o:�y�=���G`�V�M�Gn��3�dk�K�.�ώ&+]�EU�#H��-v�N�J�&�������57)u�D��v^Ǔ,LOiX�����ʝ�:;�����I��':��EV.���bxo*~ڏ��
/�A�)�^'�J�ͺ�״�[��V��^Wcu܄�{�����a�ʓ�Q-�^*�]��廣cL��2Ξ!�{�#�b���9�UZ)
��R�Ao&i���iv���e�V�98&��:;�ѲH�2���b�٣3d��ٗu��Iu�5P*��;���.mt���Ϊ�(�o��ZѲ���PA�5S���B�.�r���o�D�}�X�{�j���^�����`��;8-�e;ʷYa��s�C׵Y��t�yST�IV%�ʘ���d�^�y��ޞ>>�;}x����qǎ8��q�8�8�n8�q�q��q�q�pq�q�q��8㎜q�q�ӎ8�M8�8��q�q�}q�8�8�n8�q�q�qӎ8�<q�v�4�8�>8�8�8�n8�q�N8�8ێ1�q�[|}____\q��i�q�o{�6�ݴ`h+Ӭ2e,Pe�@�[[u��"�kN�]�v�� �E�n��9Ox�3��{�z������#w��_Wk���Ә�\�<���M�{�C,�]�p�ntJ|*�P�cjw�-P����s���
է��1X�c=��P�����F�"ZX��ZdY�xh9c��� R�Bu�*:�L�N$�t+�<�6H2l�r�r	wM��gl~�M]z�������#:��Z�X���=ҙ�������=3B^e��zv;��A��D�4����1y�WmHn��5b�Va�W|�:�hG���2��;��!�V�.��&��Ҹ�G:�r�=�k(Aa��a ���[r��}�>��H#H�2l)���ΑU���owf�f`��M��������]��<=�F�b�6T�yc�v��@�a��.�{H��(a���BK5K:��u{�Z�j�J�8oW�NO�*``^�6E��,��I-�|ɝ�5�Q!�_WRҍ[,K�% �Cӛl��,���X��ݾYᠡ�b�AV1dYwV���6H0���wVIv�p�< E<��Q^�3MC��>:ե���S �{�sNR&����{�\ww/;�i�݉�Y|�}�v�%w��w��5IMډX�x���ҽڀ��F��i�E�2�e{�Z*�5�p88��yb����_<�b޵jrf 2&���uJ�� ������E��G����Hۺ�˨Ѫ78ԕz3y���C����wCMٟ}T�������oQ�Z���SY�j�*��ܫ�v�2��LF�ߔ�'���u~�<t��۷nݼx��_\q�q�8�8��qǎ8㎜q�q�c�8�8�냎8�8�88�8�8��qƝ�t�8�ノ8�8�88�8�8��q�q�q�q�q�qӎ8�q�m�1�q�|qƜq�v�8��q�q����G�����\c��1�q�o+��Hm!��������jۦ�D�WcV�ə���.܄J=���,��ޫwC�ʰ��6#Z*�w\j���.;�@x J��b�i!k ��÷k�-Ǐ���ʕB��/�&��3ձ�*�]���`���m�Y�Zh�	h��zuw��y�ݕ�&���nW�����Tz�Э��kU6�tV%�7�i�茼�a�"kV���V�n&�i`�AT(]���5mۗ�݇5��Ybė��`�3s�J��n��iΫ�O3�:��8�uC�2{;�Ψ6��U�lAj�U�]�^f��P2q�Do��,����t+ó޻��N��a���c���{v����#Sx	Ha]�].����u�u.�qq��=��h�z;56�̔��c�FnI��J��f��;��^���]\̼1<7��D7s.�ҷ�}�O�h��gg�<Li��V[�rmk�9u˞,���0F�<2.pc�`�S���r���!*�%+{�/=GrZR�Q
pc2`��̨���ZU��e�
ޥ�N�Eʳ�UX�9�ot�D���V�iP;&�j<�]�Q�C �!��ʳt.�Z�p��ضUgc\�땵���l��n�=9�o��֘���Nݻv����q�q�q�q�qӎ8��q�x�8��q�q�q�q�q�8�8㏮8�:q�q��qƜq�q��q�q�pq�q�q�q�q��i�q�n8�<pq�8�8㏮8�8��qێ8�q�����___\q�\q�qǎ��&wIΞ��m�LcR+A�ՒfU��7�xR�jg�0lSv�������a6]��y��!Z���Z(����[�Pn��Wm�k ��\*��/�"� �\���J*i��p�2�Q�ɷ��E�D4*�1���E�;y�s�n��ō�T�ts���F�[@s\��U
=������:��;P�z���N����*m�CWN��@�y�1)baY}���6tZ�@ȠyJ��p��<�e@�c�V��!+�wZ�C.a�]����g�̒��m�̇'��+dYc/��B�u8�K�.ڲV)��.��.�3�!�{ݧK�E.�R�	���4����l9��X��Y��:õ����
{�u�H�h`ܮ>��z$4�t��d�-v���Ҟ�U�th��̭�þ[Ԋ�g&xU�Nr�f�qw�0��m��z��.�n�ӶT;Di��r����;_־�����=�7ǽ )��̫�1\����z�cW�E�/ 2�eZ����R�zm����;W^��J����2�<d1
��G�c����!�2}�7U��fl�$�����:�W�sٝ�]۵#_O����}�o�v��q��q�\c�8�8��4�8�6�:q�qێ8�q�8�8�n8�N8�8�ノ1�;q�q�8�q�m�i�q�|q�8�8�>�8�8�N8�8��<q�v��8�8㏎8�8㏎8ӎ8��q���������q��q�8�>턄b�HT��
���hn�Ϯ�cT��ђ�ӌ�{XU���ʔB�	��p�6��ޜ�f��|� �����T}K%�X�b���zH��z�.�_`/�����s�n-�ޑVYc�ׯ�[���`���/,���ˀuR�08��>��Yy���u���s��*V!���Z^021�� ]�z�k�����d����:�3nĝp���A�D*]9�,��#6���z���h��ƆV��W���ȧ-���*��t�ñ��e���w��Ds/2��*t��Q"�V�3�È�gK�\�٩�AV-�Z�.�f�\¸���n�:a�f���A�����ɷ����v�$�eyfL����E��]�E��)Kh
k�`Y|�:�.`A�;v�pTx���}�-�$x�Uo�p5��yJHK>�W��נ��&F>���d����B�Ъ���ʼN�u�ƶE�(�kP:��O�6<�ӛ�	Æ�J�����vLΗ�������MJ�A�l]�KP�o:h���&����a�H����B�����C�V�n�.�H4.���>�Q�ם������OOOm㏎4�8�>88�8�8��4�8��4�8�6�:q�qǎ8��q�v�8��q��q�q�8�8��q�n8㎜q�q�q�N8�8ێ8ӎ8�8���8�8��㎜8�q�m��8�8�q�qǎ>��}}}}}x��/���{����w��/hH��u�աT��j�����CUv��Q�Tq#`���Ң�e��5�*�V��IZ��j�;	)-A,���_cYzl�9h^h��}ۘ�Z�%���MwF1g%DVl�I��[�r�W�2���<k2�V,[Vo3$}������q�^��Wa��PM�i]+�T$G.B��nvRRc^�]�Z Qw����ՑU�[���� �{Bv�6�V����j�k��}Ȼ}9.��p	n�����9[�浢���ە�fǐ[n9��FeT��$�agZ�:�ڃPw��Sג�os�܃��豂�]f�tj��ɏF��qz�M�9v�7�{���7U۠W9��CtY���*�쩜�G��W,謜��7��.�wy@�V9m�#�7練�!b�ī�|���*r��cMq���n-4]KM�*��So&�{y4\B��v�u���y�7��$ ��w��[�f,8ei�����	S�q�3K n��^��VAp�i���F�Mu���*�T�R�r��ŀ�v9W�=^�n���n���x"=��@���8_�j\��V���*Y6�46|��X�BШf���Y8:6:�t�/�]ܣr����5ݜn����cS�O>����X8Ұ�4���2�lS�n�����T�6�6mF��W(��V^��y�ѫm��_)к��zGr��A�j�^V@��a�0���;;y�TD!|�
%q�l�����PP�Y'^�Slx.�f�W'���u�Wı_VMt�լ�s��U�z�|��iE-V������*�]"��̐>��������S�(�q�ݹ8Ӷ���
pJ��5��Ǽ����4Pj��V�lAO�H�I��ηK�h֫�r�op<b�S��V≵ҩS7�`�>]���T��Ц:4P��.[�"�'�*��b�� �ź�� M<�>�b��/6�`O���P�T}Gݺsc�|P�-��hs�re��a���.���҅�X��uE:1����VX�CH_U}��_5���h^'�v�u4��fG�6���'w`�t�Crn�Щ��u�r
��w�uL�I_m=5�V3yj�ۘ�U��Ŝ���quZ˦�e_\���5׻��bA:ʽ�em�Գg�vrgs�N�r�m�ڨ��$j��M�ԐF�0�E�DZ9��/��0U[;5@x 0�E5ћ��"�m�q��1��}�o�Y;M����ѕ��h�fpX2���Q<���]����];��v�N�n�ź��0��]f�u�l�����!��ֲ����v��+��vY��p���O�yC��\�=�͵��᧳MoX]j�0��@~A��z�iU8���"���J���\-��٨����7��Fڽ2�����3���yW9b�Z�Xc^�pk�s��2�*]���b��ݏ�e\��D�S�/7�7�{�c塞WX±s1Ӑ%D:)*�{K"��}�r�r�1DEW!�F�wj�^U͹�{2?���<�4Z��Z��c��-�c�GE>�p!X��t�]q�Ԫg��K9�0[k(#�V��]ﬣ�U�J�6��R������tĭ�ӥ��k�%Z����f�6�ִ/doGO<I%\'`b��cf��V����}�ZmY������1̓\�̢,�vȤ����b�:(�MD�"��J�O�ce��M�Ǫ��b����76�vg[�q�uapͼwϰK]f�O7(rƥLB��OZ�b����S�:8�\`�@���Bk�%[6-��6�4�/�v�Lu���N��TP�F��ʱ������4 .�b���<i��c�l�6�p��}iV����9�C�������km���S*k���6+:�о�3��,љWM�|ؤoI��@�<髋�R���x�9P�n5�ۦ9{!�'h\j�\���;+b��}¤�'X������h��Ԍy`��Tb������8�����Kxt��м�8�I
kk-���m�w.^J�:�Հ�j�eՖY���L��\\��\�YZ �G]e�g*��XսX?p�4"��
T���]�p��]8Qg�_%YVBx���'R�J<�Ա'YI�/�e��c��(��W)���į�n�N�C��\����+��0��� ;��oX���:�Ֆ��nfP���	r�ΰkZ1�,Eˬ�5�V+I�.����
E����y��8J��=5Ts�\�(�AТ�v#�C�n���T�o_������_đ����������޿�?��I�O�\��_)��M�"��v?����lD�,�x>W=��"��N��
��֖N�
�#�Vq�
+R1Y���Y!��R��$���������j�������y�j��TU�
�M\.�p��WR���C�k� v�7jz-V]Ed�V�uzܳl���EK�bs.:Yk2����C�fv4D�N�;��M|櫾��{��!K׶�s�}�pc�j���,�580c��gF������3��[��m1R�b��'	!Z��nޖ�U��ղf�j6����.���I�`XU�,���E�+�(�Z4�Gs�|�;���z�Z��4Y�m��\ȇoE�yTor���k��N�a2i�fU�O��Jt0�aTFk��h��V�R��,�����//C�N1�sm%��J�نs$b�3e�q�5_PPб��G�2�����mM�ڵ��(L2����u�͋K��Y-���+r�k�"�N���Sn&�s�km./pR=x�^N�kucǗ1���O�$6hT���s�l]��s����W�CVZՆ]�J��'�i���c;0P>Tꝕ�ôov횩��n��릪+/''��P�g����5@u5�.����Z�iv��f��(�-�p���A�*$S�E23*�mJ!8@����A��A�6��UB�SA��U.[����f�
�p,�!�@b},H*q�(0m���$J��������lAf��-P4����-���fԪ��e�#	"0BM��Q�E�ꣳ@Ըi=t�%��G9@�\�9�g\�_ᙨ���wV���������D
��A-D��#1�׎���m�v�۷���w��[���UG��uYq!"��˅^3#���Ar��	��)E���M�@�_ CTP�!!#o]<i��Ǐ�v���~�u��?aW�EU��	]������l<�\J��8��@�918�2�
�ceӶ@�nyɃ��\�Nv��M�դ3����D}��A@˞��!�çl(�
��RHT10���z=�7��o[����nޏ�^��>�A=R���P�ws����'�ГcJ�X��-u���m���d����y�o���=��������'$��<\I�+��t�o��;v����������;ƫ��C�ۓ��y�|��T��w/�	���䓥,��_iy�u��t�-h�Oo5�v�ǯ�;v��������{fP�OEǯ/����W�pNS��(r~�����aQޘ��������ǎݻz�Ǯ=i�8�BI������9¦�ˑ>};���
y�\��YQ\������$^y���_T�UUWȄP�2��qRXUA	�˕�D���G�ȩ�ǝ�U�D�#��E�%����/�r$E;z�r#�PEv�����W���i���*	�	m���m1k�v�(�^>ՖU��7_u�%M_���Z�����r/�k�g�v�	��U%ʤ�#�ʄ�$3M�
�E0�.�i�{ᾦSt���ؼ���n���,&iR�B�!�7ڶ���9�F��'�8��`@"�7��U�u���={�����7�g�B�w�������BL=Q��5��<��3�蠲s=���59��k��y�*)4�x�Y�h�3o��^�2^N�O��M����j� .��,��Y�򑹼��������w�I��˶~l�9޺�/pߚ�~����k���yA�E*�1D����Hfʀ��׻4�����s��\���-cl��)a(K7n3s`m�V3f��fd����tlF/N�9����!�+w]3;N�KA�A�
��lI���%f���6��
�;���st��z�З���ƃ�)�����<GW >6���<�4���ק]�^@���Fe�k�����[�6��ũ9/�!�8;��Dfϝ�(f̃@%|�V��ϯ���f�NU��1�7��ЎBW�����q�N���@����X:�G���fl4�L��<��9[�;�J���@jx�)gp����|F*� gl:	�-�p�3{SgQ��P;��@���7�Y�<����C�jڻ͹:LF��ZL��>VϦ���<ۛ�/��:h�'�r5PJ��A��ƻր��A65,h!V�RN��ҋ�;H�Ԫ�j��MJ+]S�q�*���X�����>|2�RP���k�g��~�����\�|%zf�͚��VU�sJ=�Lm�n�j�ݜ~���v�1��A���uZ���	kP�g���T��g�%�K񿫸�����m�v��/�N���.�X���y��zj�G�.\g�z��5���i�`f������fkE�V��U:[Qs�q�֔ʈ�EHrF�:`+��>X����;�
���2��Y|Q9bRET�颲<obO�Ĩ�+wHU> ��r��J����>��o���j��ݱ�]��9�2�v��c��CJ0�)������b�M���/�>~ఝ��%=זq�ǖ��Y��(
�>WJ��q��u*2��9���o���%��^�q�͍ɶ�PՊ��6�5n�K���8�	c���s����UL�5���o��k�}��5�P(TP}��;w�tUKR�$l]��d�g*�Fˆ�X��@�j�89��l�����<�q8�ڼ^��j�ۨj�\��i�y�Hb;>�����x�G�f�����W��2�@U�o���ìm�:?��Tו�v�g�o�>WşP����۩��3��>��fᨒ�γC�i���o}�;�H��6�I�@�<7{�dd���v�L@xX�7�(I�����n�lC<��,�����*�ӝ�L����ep��s��}�����yRj���!S�Mc)CY0_w��>�<��e�k���ܺ�)eJ�*,��������C��41
,���	d�J(�E���(@�A�N�����d^s�o'�x/�|����5�Kt8�?����ݪ�������eL��n}��^�ώ-�@kJ<�3;�H����V�:�
�5�u�LO6�=n�{=p{z�-{�:��&V�7|7=��ך�^
���,��ާW:�Z�n4Y�2e��N�sqX4��3�c�bZ|�j�����j���T��4l���ms;qVn�΁@x	�N��]���ym����7m�޻�k��*E�m�F^l�+�ey)�Z0my�wi�����d>RˈnI\�>u��yNG(^/��Ry��i�I	&{W���j���P_wk|��O%�[�oP~����̋����]�������.�۷�3�N�9�a�LИ�U��g�zZ���x�i_v�[��Vs'ƫ�A(�������<�z5��зs"0\�
n�@�eV� �9:Ż�"�$����7�g���z^�1�uw[ϳ:�s;��<fǷ0�r��=�_y]{�H�?t��ge��s�f�s���P�Cwl+��,���J��ZX��g��2_����||_ݑ�4��f>��V�ϧI�] ��s�%h��jT�YV�d8�R�K�{z��'����T�^�-��޳ܮ�v�o�_R��b������������SxҬ��)e�3sE��-���d���=2�ZP���@��o4�m��ݦW"�o�Em�ti�a�ˏ�N�ar�H�$��3���}�HF���rSާ�{������`Q���l[�q�wW1W!����ʦ��msNx���d���eP��G�E�ņ�B�\���U������ �&I�r��h$�R@�C�Io����5����1�ʅ-�O>���g'q�	�wb��=�w{��h{6��ΌG�k/�Ѓ|E�d
�ྫ��ܮO���j����K��@�yQs�����xL�������mm��̜�miQ��AR5�X�7��7��0��Xۇ�G,��6��ǯޔGS:����:��S���o���P�6���v���] �e��u�����=������tmr���ĝ��@��>,��k��d�{�ٛ�.�,)�ˬ^��p��1�Ay��N)�"�{�w�n���g$>&\����
z@%L�&�g��3�)��>�A2��:�f�k��k#I¢����,󾕀�	l&K4P8�j���P5M<UP��$��6f=�s�ϥ�jVekկ���we@UY ݫsi\$�6����F;x�{yΑ�:��V��v����{d�0J�;��ᾯl~���av�_e��S�s�hC�����	���r�}b�8$X�T��ٱT�A^34v�F�������:0���w]ݒ�h�F�ְK{ҳE��>>���{�.:R��7�bQ��g76B�X��t��N��e� ������Լؽ�W���/`�;���Ϳ��ώ���s�e�w���&aQ&5���-Z/-�j7����W�Ν���d�R����Awx��Dq;��Br2ƍW~��'�1��D[��D�SX�75�ڕ��ePޢ�O�e�zء�\x���l��T't۪���6�E�}}������s�����x��n�T�V,~���_�큏��;������T�u�֧lt�IRBO�"�_��	�\�p�],߈��� if��D��Y��گ����*Y����ryC��r�T�
�WpQ��~�7n�w�A8�F�Y�E���9��6�9�ű3-O��mV��V��O
�Y�
�`U噰9#\��N�� g�wȠ�|��V���j3���N��U��s�Z���x���T;w�P�)���,�;4�?r� �SH-R_�i�/��wnF��r>d޴BuOF�Wb��Ǹp�΄X�&1�5��P��j� ����@�Jd���&e%E�%��䆭�50:�=!�i�,�K��U��{ �
�z�KfX>`��
q�Y���{�]䮖7o��Uc��Z�c]�չz�����VmF���&ph�Eܬ����E�J��X��xiKU�άi"�[���EUnm�q���E^*��m|ML�����im����$Q�K�F�|�F��8�Ԯ��-wWZ�T�ط���𲎤�Ad�>`�`���UE�v#[}��z0h,�Đ�ˣO��2fDK�ͺA^7^�5`�o�mO��X}>X�-�;��y��������W`��3b	=r�����]Q��x\t�kJ�Z��9hW;'úW�ޗ_V�TNw����l��cw^�6fB�av�m���ol�fy��`
� &��-z�zjP�z���{�C;��h^���`G>�8�U�W)b���ucUJ*s�����C�Sp��+����v��}Q�O<H¦��{�Z��x;��U�O09����n�tQճN�������|ti�+g��lJt�X��m�`K�����Ow4�n�w
[�]���)ܢM&��:�����65ƴ>�6.�N֜�kT�sP,6אk�u�1_^�I01P�6}/=7  =y�g������lY��o7nl[��H�iZM.��uIw�5��Uw��Tm��]%�������zH'G��v���:�yW{X�F6}��nK�͹��[1|�;Z�An��AaVn뀯��h�j7։��ޞz�/���r�>N��� x��K�M��[��L��3:�J"bCNN:��ө��q�+|�=K7u��Jwoo4}�t*�~1�v$~k^��׾i�#�ަ��>Y������F3�P >)W��7���N�3/ۋ3���T(�i�X��o(������ٝ(��Ð��"��#��`�!�l+��z
�t0A�Y?m�6Hu%մ��&��N�<���g��qa*�/��
a��ٺC�(��ly�:=�!g0:E��V�� �ܓ��MD�乫�ʽ{d���N�$���fF�0I�.Q���"gs�'�h	w�����gRj3r�G1nX+M��0M�Nqj�V��(\����*Ү�2�J� ���8P&[F-�w�v)�Z��Q �o�vu��p�[i(�A$��I�v� I����%q������C+=b��~��/k�:��]��{�.�|��z�� e�їy��Dx;��tg�O�ũ��i@��݇���Ȇ���5z\�٫����˫3�*uY���^�Ꞣ'B}/LF�˾(���mf��"���Sz`��i�5��I��v�!�!��k?+�+�|v����L����Nk$U�L���s��7��Tz2�y�]�x�����G���]y_�[/��1������e��~��/�U�8��8�3��Y�}�Z��8���E�2�fjr��H$���q~��c:|�`K�C�쇻�yk)�\�˻��(^�𞬳5·��o�M�:�W\��B�{W�'���m�5�ر��ݨe���2^�������j��4��=�$�t.� �ݡ����m��}�Z�dyW��{��p����%��K%��<��@�+���Xmk]�w|�������~�}�B?�8MV}�%�{�_��D˅QCD��w�~?T�3w��@��:fRv:�`v�ZK�&͈��q����{%5[��p���c|M���|���;{&��P�CL���$�u��M΋��7_�@I��f�۪�C��ک��an�C�|���)�_|�����o�������k�绲��v?s��מ̭^��ߪ��U�B�(e��y�g.���gm%K�w+�}�2�i���R�d��|��Tܱ^V��A�a�Kq�����O>�O�_�}�@'ǳ���1�2��Yo���/
$�}�������>��⬪.u�z����v�%�mb�˸J��)b�d�w��{ʅx}H�:�L���4�,������:�W�G�ey+VϨ�5,R�q�N��(T�i�^���k ���F滐���>����S�^̂���N������Զ>c��ӉwRs�y������*������=��m������ZQ��
�[�����3]��߄��8����v���V�6�˃H�7j�"F{ˢc)�É�b��Ɯ�c�M��ʚ}�y���mB�m�v��i���[�ӹy��p:��r7�u;���ޗ��W"�zt���Ӓ��g�R�_r�̮iD�Y�����6)�,����|4+fK;F]4�'�"öL���8��j�Ԏ�),��̓+w�\_r�=�)��Q��-�@⽛}�nJI�z�O����Wm��uWY3GQ�^�8/}1�됬�h�u�������}���0{}�Qk�a��H��*�0`�\�������S��;��ڨi�m�k�Po.\�+�[���B�_����S˧N�ԧ��N�#��{�g[��0J�ّ�B��/�u]� ��YheQH��OV�f��� ���y��b�A���Ev�^ Q�U�d��˅̠`�8��}�mr�̽\T�F`�b�z�F��_�c+o�x��U%we_����5�Ť�w��MB����ǛY����;�="�3�eѷ��Pj�fR`�y{�e�Bl���}�cz�0�7ttrȻz^��׷�x��k���Ze�=�z&.�*�t�J�)�����ӧq���N�4�v�:;�yzn5P����܏2?-����3�WKQ{R�)̽��B�T��ʂ5 ���*��vQ��sx���-H��$���ybA���c�w�O�B�!ȅ廵ˑ�I'�w(`���'Ub�4��()�î�w�(�[%�"�����2�+l�"I��a�W�'7F�\sΪ����v	�"��������+���&��uv
��m���Y�o�[��/l��h�o|�X�ŝ������E��R�]�;�B*�i�λ�.�>'dh>F�E9(l�e�A�ɋDø��1�_[��6����佫t��A1v%ٳ+�֫�.���I�֜8�Y�u�Xxn9K�J�Q1Tڸ���D�c8�Ӭ���}��jd�C���n��^�gѕG�8!�{�	�ѫ�f��5�Ʈ-X����!Kn�i��%��E8�ϯ�Ou������x^h�^f^[��9�PG��^x����Bp��qԏ�m��hlL"�q�Z������ZegPJ-ygh����UA����:�ܙ�a�	�ts��u�P[����9�:T̘gY�h�;k��%��ΩX��V'.8z�Xw��61�	���m�ګ{N��ͻ���)覯�,hI��Ω�p�`�z��F�[Ir%��H�X9K&^��X�:�ەsy��U9���򻬲-���R���g��wua\��GMn�E�`1��:��X��t�Z����F[(n��MPlP�\^K�U�fۗ�U����\��r���:�-�M���=��>�}���F��F��fdU2�PF�׉�Qet�<��W�k*(9O]�v�㏯;v����ZcN9"��ߓ�f&I˽ؐEr�QC�r#軛J���Naw��z��O|x�۷oG��^�i��H� �\")�	Ph/�
eMI=�I	UI��=t��ǯ<v��z����>�I#!�;*$�%!R�WJ
��d�Ȣ���#��(񹄭V�����<x鷯<v�����Lz�6�(�k"'�]��������㨄��#���^��x���O^�x�۷���֘��eR���I5A�qT(�:UC4i)�������m�x��oG�=i���*��;y�<BW.QQȨ�Uɔ����.�w<����R�T��倲*���}}�EQ}0��')�	«���չݓ'����x������z��Tq9��IU�Φ'��s���Va����Ћ2mu�QW]�C�{³iOF�:�\f���;�洐All�����Wi�2�W绳��Κc�@A'�����䇗�ƨi��r�j�<*�9�|��=۞���Y�;�w��4�n�	�GxÐ-S8�y��f�F)u�O��<9	��C�s�?[��^5��c
+B?ui��U\��#>C| �Y�W���l��7����8����m����rr�y�f0���>l����G���U#��K���o��B	}ﮖ +�D�b|�� CA�\����O���Fr�brY��`�:b,X��*������+�,`/�xi�@��۝ߢ"W}0���.�8y~����X� S�;���U�%�z�k�t:
pp�<�{Y[� yS��guτ��S��� ��`���k Q�2���g��
�]+i`{�T9�x�q���8`[�E���)���C7�7t�0K�݀>1V�@��o���KI֓lri]�����vϚ���mפ�����Ȟ{�B�=̊>R+`V{�_PF�\���[�|L��Ň{�<H��,�����$�K����Gs���O�4�}����_�O�_mw��S�}���<7�
�9g��ng���0l; |8����i�JP��>>��v6�PE���Pm���v�y��+D��K�tڇ�ڕ��W7���p��U�+�n�U��*�n���ո�ȩ_�C�dQ���XA���#��[����=��G���+�J�L��N{��{M��#~��ך�'�{*d�ݢÛ\���{�oZ�絭OeV������մՖ��K���P�P�Y>�3 sN�n Ku����.��'d	ƺ{�:<#Z+���M��9D+ʱ�8;���t�!q���(r��.,�	>��{�r�����>�\�2��c6fv��9�/�fs��@�G\	>�n?t�Y�mn=03`�5z��4�ы��y��l$�����P��7\qw� #�0xC}��m:�C�H�,��+mķ��wpX�]b:@� v��8� �OcU?*qM�z1<_� '�yL�=�����q��̜}�F���0!���q�����]z7x5Hp(׹?��1���z�Z�F�Z���!8@��21B��6Pftе���幾
��i�.Cx V�g�#���3gK?�y��/�#�;��g��ʿ�/�uk����~�G�G+p0���@�	��	'�`3Xx�}v��0�x@{v��ifNKxa�]/��|�N��n𵮈b��#���w�w����W-�����0��b]Ǭ.��WR��-�^�
�wM�	���i 
�z>`���KƷ=^Ϫ�+� f}���=�@e.�����FN4+�l�*��Zy'X@�3��(
�2P):44Z�h� �NHM��Va�'����c�F�J�{���]�m�F,���M�Q0Aκ���W�9�S��ĺ�Nj�+ڽ�
}��NocY3TT������0�f������̳J�)�ܰ���:z��SC!I���E
��E'%�0�.�g&�h�L��wn�z�]@�96����lv��0_�}�o�Y�8U�	Z���a���� a��E�� �������0��ĞhӴ�nx,9�@��c�ޖ`,���@\�����F7d0VI����:<��'�i��l:�����0h9R`;ˮ��[v������x 3�τ6r�8��^Xf�����n�Gt>gE@��xlG�۬��3Z����&�_�2<*si;��`g)pe$l���4��H.f����w��8-��|_��dk����������;�@~z��y�,(�Y�8���ʯ������	�g.܅�ƈ��$��i�����t���S��qϚk+p�6tk�3;��z��F�S�,�vz��* <�'��s�����q��@9ѩ�&��\��ٞo5@DhL�ԕ�zj�`T;���1$�	���dϒG�
w�`U (�x���9���$�f�OG��{�Ks8[���滻���]�3.z�7
 p~|<@D�X�]���a�^p��g��q$q���n��h铱�NE�ܐ�zp`0�0S� @)G�����/���QD�����oh�D����x�=����ˉOX�Dț̦�r�N�Ne8��.��5c���.���lb�է�gK��޺o����nI+c �:��΍�@�3eX�<L��Gy��l�]���"/(��֋õ����\O�Olm{<����^�ׇ�RT��1�1�5Ƒ9�y���;5���$�������{P�I��d��IH�[��<�����i�7���Zm�KD_=�=i���p1��22ž]$����n���}����� ����rq��:Q|q�_:�f���Q=�Q@���4�Zm�I�ޒ��������V[�k7�h͹Ȉ��J�%]�p���|}&���fc&σ�3P����<����Ϯ��S٭�CN�ŝ��ُM�,���K5�QoSKi��'��ܽ�I�mNM����7/�*�'|���Wu��q�ϟƩ������.�*��j����؀�@D���`�@���4��s��v�*C����z~v�����;of@Gs��)4�p$���>�����z��z�Y�#؟�|"��8٫C�@1i�Wm�-��$Sxw�:>�8�}��DWK�'1(Oh�;8"����G������(W=Æs�+N���ZU}�-�]�G���\=����<s�����0�g��s�������s�1 �`�π	��Y������{��X�cd	p9�D=S��$��c���z1 �#�>>]����j�]�7\?oթ���c��÷w�;���u�V9D��0�f�+&�+�����{f�U�[ԣ���.Ù��$:��bv��ʮ����8�����wIٽ\��ܮZ����w�o߫��������s����]��nn���$�C�\�|9��_��'���@���	��X��d���r��"�����g58�C97��:�^ck����� h'W��#�{�_[�\��� �.����qk��^�����W��ki~J,���N�E��3�{��i��a�_�3^�F\�E��*:[��:�ήJf� 'f�H�k����Mω�4�|�q1�k7�@ڜk��	%b �-<����k�ߵ}C���S�	��x�@��t�y^t�3��L5@\ט�
26}�`���+"�%�֍/�>����݅��O���8>t"�s�{�c��o͎7C�W0="n�Ra��0�NwT�pa�;�����>0]�
?�'
���>~ &���[��@�O��>�G�F��9��׺����� ��ǖ��P%h��Ų����{�>�ᆽK�~@\��>q?F}<�۹$�����<K�kn�$�(�I-�N����#�1�������|��� ,����~�Q;c��� �&qO.|���K���$��|/����Q��5}�o���9�n?�_�O��K��g�^:��.���<}kG��^&\�3Er5�,��(,�d|B0𨸧�6[������ƌ5n�{y�M)�s2�oWU����e)T0*��Nnŗ��ӎMU�7���ˣ��G��|��1Ơ�1����/���:@��>X���S�y�!��Zϔ��R�	(�Gs�# {�@sW~p*��{�y�ڶ5x�fV��f^�<(��Ǫ^���OdE����\�#�Iz|+��3da�Ɣ��u�����|�J�L&�I5�n�|¢�c��H>����^a���b@��K��X��0��F�t`���	Z��-�]���wм���Ǉ|�7ǵ��/B�,O9Ϊ|,��>^4k��G/N�#еf���۫�=��2�s�1��i�ڟcU�]��fcdI3>q��s���/��nH��1��m��w�kxI�=�kbn���ܹ�C������
������Ip�%�����D�q�klڰr(E��vm���k�}4��o���Y8��ΐ/Q���/A9(����z���X�f��~vࠐ�M��u���y���u�/qĘ��b�E�OE�n�W.�M��+�H#��*�#8�����������ސ��q���l8�a�\�筆�ag^�jO7=�p�_o�3�,���P�Q�?"��}�d�A�%�s�P����cD��km�������Vw�~zA��n-��]�YSe��-�dUK:!��'.���QV'ne=T�#��B�j*`��*5HLR����M�S��o9ʼ<�����K��W�.Wgi��q_?7K���r�.��oEfh���04�	�J�uk����$�v�,�)h��cX��f�T:e)��5���!�d{��\��|��e��*8ե�T�y�ߛO�L�i�񇳘���D�q������2q��"l-��xcD��M�y�����b��%�Y�?�j}ѭw�n��FrA��2c�v�=n
/ 0��SǊ���x��Y/́q�i����������{~��ބ<^�=�#��Kb���OF�C�O�0�-<<4�QDH�y01�x����l��Y�9���W\o#$P��P;o573�\[�Zn��8|���.��S��[�9L���Xq�u>[*��ܠ�/M8�ܲ&�d9����/F�9�&D�=1n��v�Һ�,骫��������^6��-eH��"�Ϙ穄��q��_��b�!>h�I����s����'��-�
�x�W�����<��l����}7=v5뫌�.�Jˁ|p��p�#�υ�d^�ܦ�ɾN�����=��+�a��ڛT�sv���uw����a=S��Fw��1�Lo"s���2}ϵA�qGk����x
�S�{"�Ȝ!��+���!�cɲ��5f�W8u1A�_Tr���v��;UA�SK�{��0� ��;m��\M�7K�*�i�1*=�44>�Z$���wU����hL�a-&�O���.3����,郑�|�EFy��ܱ:A�F@֓�f9�;�h��2�l��d���<H�m腨,A�OK=��z���0�N��K��i*ꮍM�n��6c
���/����Q�����!��3�� `�����Z�~T"�|�ei�Ǟ�
�מ���M��yO�����A�7�t��n��7�2�0���0�Vs�=7T�ǯ��}֝�-��v�څ�\ �i��	���6���{���(��=n�j5�4��>�~c�ǟ'���~�2j������<C�������!2����'�ǂp�3:���Z�%�x��0D������E�[��	>7І��y+�>�e|��ԥ�A��͘~��n�Q6�ė,��W���|>\¥'[���\a���A��w�8^��KܧΪ���9��c] [ė9�M�/yB4��U��V�}��y�-�U�9<>��ֻ��C��o��i�w���҄�a'��P� ߔ��C�x�=��}裍V��nWBN��[���X��sd�^O�~�w��^����D��USɤa�H�ӣ�q��nҵI,^�/#7[�=�!�"k�ub�7k6� �{��=	Nƪ�Du�������hl���t�Ѯ0L��ι0��,J��T�s3vhީĢp�9�����y^rh�f��p��p��rPb�����t�O����6G?W�;�9{>��7gda\���Ư�S�u�ffh�	�i��]�}H"��h3L'��2ք�F�wS���sg%(�pӌ"�uH��oj���ʺN��s`q�.�o�{�>:5>��O\�hsk�XwB�ocU��0;�U�mgpX�?}�*�篑���K�~�P?M>�!��C�{Y�C���Mq�AA�N�"0��o��ۊwb!���A�x4:���?�%�k�8H8_ߓ�Z����T@/�9����bkoɔ�Dd��%�'3t'�����ӧv���R�c�wP�`Dk>/�}_Z�4�~00��2�$�2���w�[���jgFޞ�+f�x�fQ�5����z���)0�m/��̄�Ȗ����~S�r��x�5|/�(8�o�,��Q��vs+o�����{��OGr.�=6�f+��ߪ�ծG��/\t|�g�`zŜ4�{�؇�[M�Ui|�l���fv7v:�G�Yݖ� ��u��thCG��l�͏s��〄w�t���F�'o����+U3��U�+[�V��Z6�Y�mu�k{��.WR޷�Ev��	=�]	g�!;��L�t`�\�[ԕ�s��j��9-�v�����$}F� ��|��^� @���^�V�uWaU���An�MG��D���p�5�J	w�~L��������.}����o?x�ĭ����#wGw���PnLH����s�rɤ��0�x�S�:yO;��*k�%@��ᣲ�L���h�!k��cC����i�����J�}ȟ����}�G�������[�Hٵ��((���/�5T���p�n._<� �#�R	\�Y��@ ��p/}��.�j���Ik�X�T��oo'ŶL
qe���\S#�H׬��l�3�)0@:����H��7at�Ό� $�Ͼ%�@�Y�o��2���5��&U�Jv�-�v�P��(�;�+����r���=-T�b��.���z&yƚ�Q�J�ކ�t �d�M~��uV���cʸr��*�8ъ�A�w]p��
$��t�P_���{|粐��e�{��z��v�f��g���ǯT_�i/��&�0����y0���	��L��vʈ���8&�`4��P��O�D9���\�=����nAlpp����������g~��h���F�vQ��������>�)�m�!eUv�'�3���[Z;��P�C&8��)�c�nM������zhn�%�vv�M�+6sB���:�٭]�8;�m�4���7Ý*�y�P܇}{�u�.ٵ�`�鹻[u��Z�7��v�,u��j�]�v��^�	��@>Ck�ef]eLUc�`6U�B�0���.�Z�8��i�7u�cѵ�g.M��5�V�pnh���L܉R����P�Ut�rB�Tv�vne��L㓩��*�vV���f���]l�Ȉ��r��S�=��:�qZ���+�6�+:�Wt���}�����]PȺ;�Qޛ��M�ÃL�Y�� ��S�q5�h��|�$f�����$�@� ���]mm�j���6��d���˛Ca����8m)�re�>,ly����5PfYvUc�]��;iZЄ0v��q�𫬥�u���p�z��Q�&�=c$GVg��P.��%��Y�3;����`J��Ùo���������&�T,�����1�e�4�Iѭ�Ms��$�9T��D�����u\��+;�;2�J�E��7C��W��EsSrb�s�/����>q_|j�$q�,��cl�BƎ��<��J��Tov�w\듭*��%-��T���P쥙�<jHHfM����\
@$�V�t]�6#h�Ne't�G��3�X��GTf�&�[��T�W*EwA<痪�f���O[��2u��2��4D(B���"�4�Ц{�}{SN2�EV�m����F^j���M��
�m�+�$}b��a��D�bA	V%�Ī�˧�A��gk���g���y_;nZ�Hu��ki����KTt%a�IYa��K����x0d�):�V�%:N3ֽ�*���{�i���X*���NܽKr��1�왌gK�$��R=psdS�u�RYe�}�m��>i���}�ԅ3����?dzޫ���7~]�ѕmθ�x�㽤q(,X&谯0":P9���a���9����d�ul���tf��V����%{��=XXm���]���]xn��%��t��TP�S�u&3Gl}yf��&��,M�`p���,�x{��İiS�d���q��6~]�o餃]g1k�TX%v\x��7�P;7���FT̛���w��k5s��"�O��G�vk�bz뭎��x77#��ڕa������o;,��r�,^����065-i�=1��7ls���9����~���z�)2����3�$돡�P�jqK��!v����X��\�
�4���7X�iY����15���6�MU�������L{�F-,��hI]�[���B��0f��m:�B8��	���pA�XPVd��\�U�ZRъ�>Q�lvq�]�5ܾ�W����Q���N:G�Q�"\����D�I���R	DKFj��]��H��b\�
��1RVA��� �K!7.��)Rh�)�p��e;*$�3b��(�,��L2�BҠh��v�F����b�Q7Fx�삩5�8e!Bpt("Ҧ��k��{�)�)��T�ЪH�
�#2�I��	�(��[�+Tk���PdCP!#��'�;�nK�E��߸��'���E��D��_���7o7������x�ۃ�������B)U����$Gs3���\��S���A�%F���6���O[|m��;z=z���{���V�5z(��$�QuC��Ğ%Ar�g(HH2>=cn��t���m����ǯ�k|����9�m$��E@QQ�DP��'�D��-��HȒ;����:t�ݽ|m��x�z��M>zH'���>��ID���\��2߇�]����!�X�����o����oG�^��� ����#�"	����iD�Ô����I�%CoX�ӷ���_m��=z�Y������C��(*���}s�A˔Bd�DT�(�!��</�H(/!;�XAq$����wB�QDs�9L�AD�O�|��[�W�4}�s�z&	��(T���OLzu��	umtM�'8�tΞ�)��9����g�A6V�Hd��"h�1�!����
e�c޹���K�OH4�˗cb�<�AZ"[�}��IT��]H#u5�'���"�2��:NZ4��8m"�!��h�5P۫��"�&�9[�k|�2 �?��rە^>�Ժ�� "T��= �#�	���sf5KiqX��f�A���"w�ި�<��g����ߦ*1{A'jw�W/��ՙ�Ea�jk2!��^�Ʈh}�"	�)qm��bm�ߔ)�k>Y%ry[3�ݔ���ML_ż*ڤ]↹L��'p<#�ކ�e6�J=}#7�ڲik���^�m�s|���8Gs�&���_��J�P8��A���y����&��]x&�[ё=��Tp�x8���)�˼�+d�'�����f�ēa8~k"���w��Ed?<g_p��ހG��s�u�qk$�7��c�G�Wj'�~�r���o�&�D>^^�m�ݭR��Ѿ+�Yqv�Z����`���#��n�اf��)�'f�X�0�5�H�ߴ������n��(E�RZO���M��C.}v���7�4�5���E��� ���n(�>w3y��k���s�.�cm>}�h�(7
Ρ��2���+���7|T_-x����$ <�ٽ����r��u�8��v�i�2��8��B���P�5�05^\��X�΀`�|��}N�}��ok]�}��7�5b���B�2T5�o`�.qPX��kr��8��k�D].�Ø�a~L����x�<��z��mwC_1�$�+����p@�C�oפ9c�r�W'"�B�s^ݞ�;oA��%ý�A�t��^��B�� 0 ��BT�BDnU֧]<�n4��ضiU�ܟs�f@���"�k<4@���<(�{�cs�5a�nz���y$�N��0���&�h<�$�힏*a�ە�ɨ!3��e����,�Rw���Κ�Ӻ��x+!�<?��i��~"���sZ�"��9��QN9�����K�o:�V�ܘl%��w�E������Ƀ ?����I�Gdo��P�`s����x1�ͱ�Zi8a�o�9Iq�p.!snn��9L�D���#�����#<��Ze��\�L����~��n���u���y��~�w�z���9���Y�C�����%�����$F��!��_�H��r(~���9|�E�X�ڙm�9b&�L*�lƏ��;�!�%�5y�S��:���LX���'S��Ff�O�Ȑ(�#����B��厝�y���XN7�s��Κ�Q��B��/F
'X����y�Q� ��")���x'����3�~#�7�WE�D��XoW�}l4ҾW���r��[M�v����v�}�M��v��Ȕ�	�A��^�v�Ҥ�o��Ɩ?���>�/��3��Z {/�w��֨%�vM��f�<ܳǣ��:�F[�e��Xwr��GN�����N3"y�Y���F�z�U�LY�sM�y�7��̙�c�*�9�➉o����`Yl&l�q����k^'n�n�ؾ��j�vf�ʘ}�an40����*xh�G1b㣽��^|��I.k<e܆5���&�<=�ܸ�i0h����`'�±����a�GV�^����KC�n�.|1ٍ��,�K,�Y���&�i�S]�Udt�$O�8�J�64gm��GgNWfZ�H���
����1��aJ
 NW!0�h�Y��i�)W��T�O�-sZZ1;wk������(�m�fB1�7vw���l��C�1=��LL�4�0#hW3uf�Ǐ�z�IC�!��}}���P��-��q���4�@@˥�]�z����H�=-���lu�6D�u���F6yٔ�7?n�Od��� �ù��1M~�Ӈ�s�c�ƍhL/��Gw�[uz�L��*A��˘�]c
C�>��k/��D���.i�s0�z�]�L�#SJi��&׷Ӯ�ǳ 0���ݷ�ڕ;ox	fT��N���0!H�p%�k͎��ч���Ru����[CdC�#iVk���&2ˠ5A:�~W�H?����|8�8 W>a.$��v��R*�b�򼱿n-<!�2��ԣ��zO��g����G����_/bQ�ch$����I}�x����)�����v���cv}�_j���FS�D�+�V��;t�VQNg��"�
��JY`��Ѻ�-�[��7(�J��%t���撰d����ٜX�n�޼�<�vk75	}`�A6��8�d*h]��qX�m?�2�x�	!A�����Q	_��|����鯘���'����t�gy�vCzbO��RÒ kg�ˌ}.0�c�p��)�!�4\�~@ykD2�y4�Jd���N-��)|hz5g|O���uQ:l	$�f|�ޠ�����;T;�jc��Cs�I�1k�}�����&��cx����}�|=b�X�ʹh/l�W(�����q�S�,S��e�' {iݲ�o����j�����C�|�:C���es=L]���]q��K���ͨ !� ���h�r0>UΨ��k��˕�R��>9������<�^Vv�?މ��O�Gw�>��zJ�TM�'��Uʫ#w)ya'��K�W:�M�3G޽�yiN���	�+�W�?L�Z ��=-�)��d�5�I`Z��ވ��;m�T���wkS;�Z�ZLK����O15����+��Gh����D�����x���)wfU�s���'��0�-��:g���=};<<'}�{+�b�ɤ��`�f��tW%��O3�*D)��nAG�;���B���nq�K'pm%�xw;�}��	ߝ����H ��V�"�����:�·�tl�\t��S�j.WIB�_d����! �vZͻ�M���d������7�+E�l�MT�磦�a�l<i��`S;Kг릿z�IE���S���'��R�^y͈��T�Sb�lK|�9�.�����m����J�F�Z��b���v�ԑ��ʂ�De1#mj�S�
��|4� �!h�#�f�����[�Hl@��ă��TC *!C�?<��
����wnڗ�È1���=h0k�}XD��{3�q�2I/�#9���/"�)|&X�я櫜��NE>�_bƄ=�y�x����m����q,�'!T�hV��A�b��u���5�~1�8����cNfs\,�Ά��;�L�I@�(|oc�����ˢC��67�nT���Q��2"1�|�s�;�;ꯄhP�;�[_:|�Cu�@��YH�	1鮉����K?+����V^`��;[��6����R]�j�q=�q��ѿg��7KB��[�'�@[�8�ޗ��GB�-҈3iG�m�\�%K�c�6�|���� ~,LsK��<χL�=�4���w� ��̼r��l�2+\b��R��
ێ��֧���������ʏ��Pᚈ!{Q9�
(�}K�7����.#9��V?a$�F5�g~�-�p.7׏xA���"��$<N���5�}ɮ��y�9�T/Y+��ym/6=ȟ&=���Y��9-\郂Z���v�nʬ#w���s���l�σ]c��]E-�c�>���[�Ǽ�U�z���� ��H�&�nJ�'~ ;�����uQ��A���ŀ�E��!(��1.�/v����4��k�k~�5WwO}���{& �ղtC����f>�İ�A�����}Z����r��p^���+���놫�s�&���I�$��#�Ʈ�>d��5�7�%��N4n�.�a�g85p�D����v��k��`�A��%D
+	DD��v)�
� ����'޺�mG��ja���3��[�7�@�O�>(��ฟ:P����4�����{a��S=|V\��m��,�������-��~H F�@�����ң����@��u	��n� ט"ٺ��f^}��8�p��{��w�pS��_%���l{�dkg�
7��_y����5դ������9X$�l&�|���ď|U�_i�5�o��lS���fpx��.�Z����~�ib<xiN��F��m)՝v.oT\4��Y�1��"�=`H�l�\�z�N��aeM]}x $�{<�f'��=��m������=��<�!�/e��OL�#ZC�J��tw�Ok����[y��w�J��`��ݤ�>�K�����Y�ݺ�UDd:9���{s�4�w0��g/̋��ڟc�ܸH���<�����ˍ��c��-����+_So�4�a��w��D��ce�����_��oL'�j~GR}��C9�g],a�ip���^�|��S�v��<m��<�j�s�����Ovf��+q���9t?0`�5��,@��"HYO�\�:�+�J^]�c���D���b��4{}n��ELKhn��2$�L.����2�o!ޫկA��hDb�ض_gH�}���A�(�T�h��*�T�b�u��"�q8M�Z�t��l�˩��"k��*�eu���)N�;���jPB7pu1r�L�s��8x$�H�$�3�К3�ɒL$(h
�2
2(}��o�ߕω�N���O�oF��%#!�����~vr�C�i�4K���?��(f�3��[�{^�݋��1���j<���5'� B!���k�2f�N(6F�Q|,��\7(���I��)ջ
��xI����V7�����I� ��Ї��m���P�K]3\U�+f�@��g��⡓5Genh�S�xU��s rlL���X�iP�����.9��!���P���/_�_��z\l	�J����߅i��E?����1�F&z-}�A������Y �Gc������6��}\�eDJ���ە@�4��O�
gU�h��߹���UHu�(��ו� ���'�T��l}��6��u��T���7p�Ì���͌�'�q8ΪJ�6O-Zߥ%�A���*�U���:kw{F� ��Jhx<6u��zY9�o.��3�M�$������@%D9�|T8�����^���_;�3l6q���L��ߢ�=%���sdHw�.�M]=�MQy�w������YL�ӤG��2�.ׁ�C�>=β:�����}=���,�vE�����PC$1h�gåm!�c�յbQ!��oMܫ�wvxE����Wf\��%��s߆9e�g��bɎ֍��)r���,�����r�-�Ut�>�'�v�k5=��^m;v�fwMb_�ȓ�u������*P�(41Q���R�-E(�C�E��{�{�����Ka�dD����fǣ���p�:�8��4ў��Cn'd�ͅ7v5��Y�3{5;�zm��f����'_=�����$�z�4`{�Y+�-=�Lt��orh0&$1��	�h1�l�RwV�Ah ���(A`�9��W�˽�&��h|����}��&��=§1CH?�pp����B���M�R36�S�;���5Ĝ�~/,�Ӈ:�]8c�UA�t��Zx�c�[����n�nY�q6e�9�`0��40o��4 �k��8_��̚^�zI��@�h�b݋=���p��UmC|H�6��5E������S���)c�'˾�w��[�l����&IӺjߚΤ�e�FhL8�O{�ir�>v���14�a����g��ìB�5�G�hBu��ëg33�epM��}v����Ag�᜶�i�a˞m��z�O�{ځ|�mL�Eֳ8\�����{�c�>�� ��9ن:�z����-�$��4q9�U�E�:�o��ˣ�v������ؽü[����q���1�5���Ƕ�\��I�{\԰���o����b+���o�6���f�����3
��i_c/9�9{ϓ'���J�Qxt�C���:�VzI���r2���TR�Q}m�'g_���\��wI�ŒE��Ɍ�L��Y0�����FG{��Z�ˁ=�T�E�[�5�Pkl8t�8�)P��R1*�,���[�Z�����#�b�740EL�c1��Lgld�1& O���	BL���Ɲ��s$�0a��"d/U�?7�q��%?�sș������w=��&ox	w�fo7z�j�v�cYM��ow'�������j/���p$�6�C�``#���'+�d��-Eg�����������1X�^i�鐉�0�-�|]!׉�)k]���&K:z���r��%53uNn����cs�k�[�����:�z��H�]�d8�8���l�M<����p}V9��� B�N��+�������?��˿�;��z7��fQ2-ƕRץ�.W����:�D$��͖�g3t�O��ΰ�����4p :�����Z�۽se�q�Y�o�l�t�g1��(�pl��0�L{���'�i�S�@�b�%�	�M�s���^����ս�ڻ�6(����' �l��T�ǌ�N>��/�,i9~���ٷ5\���[c{n&ljA�Anue�v���8�p��[��	l W'�-�C������bQh{-S��Ia��f.��q��<%���+�/�v|�����1��q8Ys
I�.Z՞g�z8Ӻ����������@+�nX�/6��v\º�cqIZ|;��qwݑ�+�����>��A�����U��K�ty�}��&vL�e��ˌZ���A��D�j[SI4�WwU׽ԞsOBDofK{m�R��T�P��hb# $�`(R	x�[���}D7�~���zsLԷH!�e�H�Ϡ�/�m[��Vp�Ǎ�wn�����]�94z<��KGK���hM5�Ǝi@�X_>5��#9��`��y��OY��h9u]w���HW���Θ�ȗ|���W>װ,��Dt����B
I1���0�I��~"W�N-��0QC�]���n+Z}a�ޙv;����'+�>:���=9��5�����\Ҫ���M&�Wc���i�4@A����Sa"Z���T��	a,���t�PY	���k�T5S@v��\��p|g>r9Fz���u�=���u3~l�_R������)�3�6��\!�vTLp@�OZ�5���	ljb���4�J�p�3Sh�A��v
ϗ'~d*��|�3�`�CMյ-�YE�YP֢ i1�kn#���w3�l4�ﮜ��� T�38-V}Y�%�*py�8l�V˼�������M���0oe��s�vz�穑 G;�r7����u���(�!�{� �m�������t�,w x�!���`f)Mc_����sA��z���"��qg30,���`=��f���6�'j��I��_����[���q]�G��9�j_]bF;ޅ˖A�$�%iTQ��oL�b����y���aM���z�sr��+; ���o�X���plU\:�6h��M���z���Tj�[���GC���%'BE�;�#��ͽ嬰���^��y*�vp�Q)���rM!f��Ğ��3�w��JQ�oB��x82�$�Dx��xiu��d�����������*�
�
��/y��PEX�j>���G��fo�溼+ �����4>�kC]V���/1C��:Km�\gf�;-�t��r��&�]�l�ȧke�j�s
�X7������E�K��e�7,w`r���GV4��W%T�_J2��y�zJ��
��k�.ٽx�+���_r�k��z�]���q��P��ɽuo��.�gQ�t��Rq������ۭ��s���%{��c����
��t+����Pj��@�ī�IӔ܂S˭t�)����n�����"æ\չw��oll��]�d����.��g!q.�~��=�|���+�i����l0�
r�lv�V���t��',�}ڝ�x9P�YkXفE���f��v�o%��cE�ޖ�]�C�'.��-�z��� Y{�AF۱PM��xl{�����E�t7�Y��]�6�U����:.i�d*��\~�(��7;:���6��~���Ǖd��0ca݂@H��:�	��)�R��h�C����Da�7�B��ٖ�<#���\n������`���Uq��9�6�;u��c�<i�9���ٺ� ��)����Χb�-<!�����ձ�����
]�<A��ԸI����C�cZ�tx�F�y��ww2u({��{0q��̙�(Y�O�:"ɴͺ�]����)��:���Ͳw.�Mq�i�Θm�cʈ+n�;�LfS�)�ȱY[wGn``Ԣr�ӈ��8�V��2G�^Ν*�#HY�eM9Fˑm0���+��>���2q�44b7ĸmEJ���+,�7N��t�hѥ�z���F��խ���dg�p�9��v����K������R�z�4�3��w8"�N,��Zq�>�m⹘C�#�fA*c�y����"��=v���®�YG�
�&c ��[�鶸��D#�o��%T��X��<g-p0�Zh�/7;��ݍ�]ufHb��'��O�'f�\��������o�ޥ�� ������!v���U���Q�QL�8ث�=����4�@ҕ�u��cSZ��F�z2���o��b���
�s�V�)tr�֎�j�Bq��$VIx��[,�z��yY(��ѩ��K�p�LHu#<��f�]Ų��Q���7o7�||m��x��׭4��d�Gؕ	�w"E�9܋	%K���Gx�����;�r.�&|z�n��m����m��G�^����!p����e�g�����H~�#�$����/J���"�O^�ۧo�<|m��=�c֜=�!'��k��$���z�5
*�X��&��]! z���v��׏�������=m����E�9z=��x���9r���dL�)�W
����g{v���<|m��}zǭ8�dOξ��p���4k�H)0�|�T$�x���v���Ǐ���o�}߳���~Bդ]&�O�>#�8�H��H���.8Q�H"��Y?��M+�~�9_6 �{HzI��.s���瓇�d��%���T����w�����%��t�r��;�V�n����աĭ�*n�����/}k�;�]e�.�`8�X�C��G���ɻn�ɓ0��}v�F��쒢�[��tu,X��f��� Yo��BA���J�P�* 1V��U��"�[��O�~,>h5���\�M�0�����"NMR�{S���7����(̍�}��l�ò"f���xg�0���e\�eZ�[��HS�[r�i癊�����\�Q�;�;3?��x���Pv�A"���Ϟ�|�A ��y��N��e��]�t��d
l��aQ�<��&������C�1�=����6{ e5.j��8ڂ;���-ۑ�i* L����<����A��w�B��O%#/�:�ȉ,��N@c�_�B�CB�ݓ�:��y�;Qg>��/;�"HxD�fZߵ��qoE�]�S�J�w�sE��'����9	��nuh�pw��$��'���Mp���j9��0��p;�6�٧Sf�?�}����r�I��M���,�7�<4w�$џsK�Br|�q�ql1kڰ�b��#}r,�jkrp��Y���y{���`lK��QΛy�!Q{�#�����\Sq������]:��X/��1���>�*�Di��z�p�|4e�d������>�:�\��7�D,-�n�=��Z�9�۽�{�+�r�DV��XRRv�Fr����E��S�f� ����:�U�PB��Ny�2¯3�tP�ė�h��J4�kRg>�UTB�{�U��/	�px�s�p� �q���4gci0FC�"b2`$6��!���u���{�o�#��f���Lo�&����&��*N�60��=�2����Y�uG� H�����3:��$�[ã�H�x D����%|���L��v��f�X�]�D~�&
�����Qϰ}�}k0�M6r�I�����|����\e�1�wHx�z[��z��h�k���u͑����Ǻ��l1ͻ=�71�����x���˸DI���h���z2�D`�G2BS��&Ug.�Z'7����g����5Aw��V^Wӑhc'1��Q���������k���uX�����	<��O����ߧ���P�p��k�S�0v�.E�<�9/�%O>�'�g'��Du��.�;hylx?ȯq�>�EqN3=��<��}��ψs��x�y�y��Y��\+2��r3�-}�ºc�L4k7ҡ�'
��/�Q5�x����t)}��վ6D�ʋ܊|�5�	��8G��o}+~�_�����p���n(�M�����7����r�/8�H�g(�m���d�q��j�IzC��ms�^�I�=>��\ܾ�?\���;�X��[��e4ݼB���5\�����k��lܫ�j+�/�(�85	�w�J�b뉑c�[cWM���t�i�J�ݲ�����t����X�i�{����8��g﵍�jY�>
S��Ts�w$#���21W*�Υ�biS*�&Fj�1H������m��*n�b�T�)D
3��� 	�2bC66���rP��=������f�!p�L�"`��ŧ��%Z'���p�����+��]**��2��Ȱ��q��Є��Wn�������>0u��b&�&M�F��v�:@r4�1�� {S��X��!������S��y��\b6�s�Gla)�=T5I���Jp�+��n|B�����68��';+6?{<x��'ƤJn�\v��
��,�m��Zap��W[���~3�n�c,I>H	h���9�Q1C'���P�/m��0(b ĜN;Yzg��ʕ�ﹺͪ���tD��U2.����-��f��#�A�r�p"�0�d�e�]�\4>ڙ��~������KA��xP�W�O)�G+|�`< �]���Ur�O�ޠ8�Uz5��'׏gbFF��&�:u�|�ʈ>|�0��:<f����23���߳�w]	l��(�/�o�.9�����o8ވȯ=k��>{�����LNu�cp�����tp��Ԣ��o��s]֩�<�`f�at ��WO
]� UU���_>W"�h�ul%�x�<4"�ݣG:�M���D� ̤#�ʬ�p�X�+��bI]׻
��'�$���L�����^y�kc��<����鰘�캋�r��h�|�fs��G^]�1��Cn��f��D��V��CO�P5��j11�3���� ��Z����v���9ߟ/�!�|��Dr�1����W�}v�svXM�.YBC��gv���էs�cs[<�p��FC9�v�k_�����Zr_����F�m��
�M���-105�-H�պ��3�G�'ů� � ����ԬZ�y�ߞ��!��i�H<n�j켈t�Nm{	1�%��+��y���m5�Y�(Z{L-8�eqBJ���';x#�#��I���ꇍ�����w�x~h0n�7��7��v�m�.�ˉl�'�z�+1r�>$�mݑ8�����x���n8{46s'Z����A�U����x����O�7��o�����s��Cd�D{<�g�\p�+�v��3��%�J���&0(�����m���Y�o�p�m5z���"K���;�=�.���'�y��eٓQ��ΐ^M]ޞ^)�m�9�q�έ�i��0����"ǎ��U���K�wl���sY4s�7wE;���R�ٍ����|���f�G�!|�c�P'�,��w�����;L�\d��<%�O߱�|�9��Bۮ�&S �oV[��*#�V�I��?5o��_w��J�M��MqI�}�'N�s��8�UR����Ɛ���/꺻��5'o�r�Z�H"���9� ~�16��@�1�:C$T(b+ T	d 3�kx7Z�4_�ASf��=<}٬*5�m�� ���V¶/5T�� ��,6u��w�����x��d)n�����H��s�$��b�|���ǝ�0Ȝ���k�]�u�T'~�����RmMV��/����O�g��'~�b�� �	���Z!��U��;=t�*|�q(;q��8�d���b`8��kCR����d\����x�O.t�W6�F�ݘ�;�\�)$�EuR@�xm/��q|C	X6g<޳�*2w?5K��Gi��/ǧ�ѳ��v7�1ص!�*�w�电��0`�M(qc@}�	a�3g�<��\]c�a;=EȈ����M�a]�T��'�������𔱮b*�k͟�`>�KmK�' k��}B��xn�)kV�1̭�u�˞�\��Z�?���G_\Y:�C+�������O�*��Ҟ�{'�:#��sٟ{�+����D3�~X�0�� ���%zFeav������9��`&֢��L1��=��� �����5��W�k1�Ks�X�N�sL��͓ �L ��w��W�r~}�ɮ��_f>��w��j�1kI�0�Re<�y�����چ�^P됅b����'U�W�kBԾ��.����eiS�h���kF��M�:��;V'�{}C#�8F�'��������&��@�+CAjP�P�R(P�R��� �ʙ�=���p:�k�A���>XF�J&���giD6�l>����6��g�ڣ��n�N����nME����{��ϱ�,�����^��bE�p3�˝��0pL�k�|w6�~��/��V}33ݻ�:p��%2�a�!���������ƚ���E��{�~*��w��Hk�]|g�"_��Q�L�K>������G��u��m�#��m�͉Vw9��|t��̙rQ﮶�K[�م}���s��Ϛ}�P�ᩳ4�[.��-.�O��%�"�N�����؟&7������*�ÒX��l�8ld9:kڝ)z>K��MtÀ�x�v9̩�MYg
Z^-U)|Q�L���i�����^>�:������g�Z��}|��q�Ú:V&���o'^��V���=.Çs���ء�� �
!r��8~O�^X3��I���l��"����r貥(�k3v�x��(��+ц[�gƃ�.0������z������ir����ɧZ<f��#�/��}r�3�y��WO�����1�N�0�����g�{�Яؙ��iގ<��C�TbTM$J����U�*���GMy����f<��Bɽ���]i�yR@%t��4��	�OѤ�5§yZL�bU�C�a�B��&5�ܾ<�e��6)Q)Y�������z�����&]�Y�4�h�Um	��R�4j�F�����4}�C�b��)CQ

��!�-TB� �� s�Ue������|5D��SHc������3����F�Ui�b ��7l.�]��>Lp��E��{��5]z����xt@@� Ĭ�4B�5����,l��
�xn�|��������ܹ��Í�p�t�O��5��s��t�Ij^���8}BfN�I��PQ&)o<<Eh�*����)���ė܆D���y
��@��U򏯙�/���Ax��`�̀�3��k��yjx7�f�%��NF{@��5ޡ;�V�<�"{4��q�,�בL�u�.�1�(<��u����d<��@yX����6<�1�Tax`���Mr+�79wA5�_`��
������C��!��!H��ޫ��Ic9��~ Op�d��9�k����f�@�'w�ew��w��\�X/���k[��MZ��mM�+�K�k�Rj�Ҝ�I��;=��yL�L�xRD���;���)���DK�[��Eo?�cqg	�ɉ�[AP�(�>��f��ޚ�
pvM��|��^j�Ϙ�LB���C�������N�u�F����ʤ	+�����+F��eْƲSd�j��_�Ks!�O�S}'֗V������a�x9��/���R�ɵqm�/˭T�)�3�:���g��1��S�`��=�'8�m�Mҫw+`�Dݮ�7LJ߾��e�����{&yu+��/��j��PP��V �@�E�j 
��,�Ȣes������K�\�Ͼ�i��sΩ�0W�Z[�H*�ݞ�FȺ�x;�s��)�]�͓Z=��uzMj=v����È�I��K���}湭�j����A��n����d}�w��G� �����d��xSvҁ/�+�O�y��[o���nƀ���umfv�f�l��'��F���BQ�L�h���k��q�ځjK�XNAz#s	�\�t�n=^Vo;�u�g�BK���Pm�.仲#�X�{����Ϡ����>��.�>~pY�7m���A�C��B�c���� �Y�ó� ׵���Q�'�3�@�~<s���Rw,˲�����W=����4rgo�P5L�1�~�p|��pJ���q-<��,���\�_��z4� Ѯng�,0ލ�̾۸pC�?wE��sM��M{d0��!�g3/�=>���;�ۇ�1��S���hg]�+����K��S�i=I��q���8K>���E�/�5iٱ�s�����'�Yf�jY�&_<����uW���=0f�+��%?�ߟt����V-ĸ�au՛7�T�eo�s�Yzw.�{RI!K�s>�W��s][L~��LW��������K�SLq���U���E��t���XP��w*��Ȇs32+R�я���v��l�B�C�`�
T(`�&v��g &v e0�!I2��y���9y��䄬�[�ɜĠ�N<Tl�^!����ԙbi�C%M�4�:-�-5����o�����H��cX{���%R�9��I�퐚��ik����Ґ<��RD9�k���RŰǀ^�A�B�Zb�|�D/͠��I�a�n� �����Qގ�Mi�{�m�j�q�`�u�1^k������K-r_�����߹�@��@d�|��ڂ}��<�=ډ��덷A��,���~}5�b��x��ɥ���7��A�Sa�>����^ϧq��� ���\h��HvG7�s������v�ok)vHnù�(Լ�d[���@���#�ē=��D��r��\�^t��k��{�UfN�n}l����OG
��H$,3�aQy��m����i�&�]�x
>�����=2/Uٳ�k�T�
W�a�ȇ�s���E�2!ٰ:xק2Gtq����3R�z��N{e�d��O/\����0M"/��]D��c�>|���_k�ɧ������vM0��n�CkT��5E���ܥ����G��e����(����oa�Il��I;c�(�l�� ���p^=����k��>y���74sV{M�&����6���7sz�Zߺ�՞��z�9��^���J"/�b���T@(`�"0cQQL[�U�ro��~?&Ӳq섚M�m!�y���6A����r۾!ٞ��G���ӎWV��<i~>�z�d$-�g�>�Kډ�S�E���|���w�R���Q�ϯ��Ϸm�h�-�� gfz_����縲	��S�{�4�yUy)u4�4���?��G��?Ox�N����380��9ڍm<m���[�0�u	|�0�S��������<N�����~(&4ǥĿ?sg�\��#��Y��tY&��5��x�]�Y/�{����/����a0P�Y�^���5�0�~��T���	�0]��Z<���Ū�nZ���ݱ�T��{�g�������=�b�L���{�@�T������Y�=�َ����4�q$�r!�xpCk�}H-���9��S �K���\74�2�S�4�>or�3޵�����&/� ����y���2�rq餙�$(ق��~�"���|���s�������N8���'�*	{�ҕyE�.���
��ݏ������A�-=*T�Q��ݶ�FS����| )T΅�3.��y�����9%�kK6b��ܓw��X5�*j��
��s*Epܚ�>%k��^\7�j��]���ѷ��9��{&p��C����1eK��x��1�[���1�P����jfc��#���U�i9�V���^jI
����4�Yis�w�UW�8\"�Zxp�m���e!�����2�.���B�M�F���V�YN�{��#�V$Y1nn[B��<���{ъkw��:Wrnn��KV�Ul������6i�43�e���o)������)پ]�ON�֓��޹���iVݽ0]���6h��%���P+ح�W�F��I#*����&]`���Gn����֝�`�C��ul�R����>T]�3g�vи_NU�U�Њ��[�y7�D�6��xA!>8�u;9� ���n��t�9WB69"yY+)U�-�O�jA�E��x�xl��60t�XUǺ�M�L�a(�}�4�:�����;.��9'L^�-�Uu�ٮ�nc��c��6b���k����[�m3�m�P,dQ���<�0���6�H���L����ؤ��.�"�n�(���Hh4�J@n8l�d��/q�q�@�I�AS@�6U�Im��ti*E�r�+(Z��4�[N� �HR�Blf�25T1zGa3'��e1b4�*�Dq)�A�����CUJ�(׬�V��F�vg9z��<�A�Z�����`E��+2�b;{1�#͸3�;�-�0��M����2�/{;��w���ݽ��sb����D�ƙ����ͱ-���khѵ:���ESy��u��ո@���W��4��uu���������j��-b����\ �VuILK�G���W�:��t��EBIǭ�D;ɕ���T��6q��Ò�`�T��[�m?e����e`�}�y*g:�_1��:�IV�b|�Y��t����0���TݧL9�q�Λ�[�IǤ��c��c{<����l�
�л����/�[2�W�J��F�j��P)��k�M#bj��+���2Q��5��]��s����T1�yc��m�-Jn���ܷn%�ۭZ�[�'4�	JO&p&�2@�3]�m�b4��54�p6���>I�P��z���Tm��,S\�kb�=ɬ����DC��U����ɢ��;��W�.y��9Hh��-Âmҫ��.罽K�+��ب�� �rkP��M�g�*|�L��{����u�\-�s�N�uN�\<q�ʬ��dN�Ǣ-����HW`��t��P1�0(.�=�.�(G�P�'<�yIF�	P²�,�L4�uu�\f$e7�B��6�8S4"FJ<�"��>�MW-�K,&���v�Y�w'(ݳH0��E,��!�'�i��L�����Xt�bF<4� �~/rക�e��@��I�J�A,�Z�P�xdI�����B�LEuBɥi��r�^oB��p��C��ߖ�˄OF�xZ`��EcUP*T$q�c�N�z���m���o�ߵ������*9�� ��v�9~��.L�4�	=c�n�=z���m�����=i��D$ߐ^��§"��+�)��yх��dS
����gv�x�>6�m��c֜=���*���):d�ȩ$4*��m��v��׏>6�oG�X�������4E����ӤYJ���Ahr�TV�~c�N޽z�����m�����{!CD5RH���ҿRK��e�+A�=s	Þ{�Z�y5�Z��<v��ׯ<|m�ޏ^��w���@�~���H�r�~��)+-)��5�?�wo+K��d�A]�*�ל#�QUq"�D����9q2��I�|�y77G<24��K�����T��W�h��t/.vS�����^;�O��x�P��p���1�'<�BF���G�Oq(ח3�w��4�N\�'�NJ~n���j;���F�9eӕ�f)�x�hn�G��fS9��@(Z�I�U�2�L���l)�����"Pd��q��F[	��'Ȍ> rs��><G�1 �C��
Ț%E�S$�'�礿g9�{��ݚ�dA�� �ĳ�%D��k��c�W�6�1���ʀ ��=����=Pֱ=�6�{��組3�u$w'�a M;r�X��Y��H|X)��	v��:{�ױ�L���~Ȍ��e��FP��=CC%VSӒAkẦ1��<�	�&�?���������מ�tue��Os&a/=��
��ibHr��������ɯ���nQ^4��x�<6ߛL�97���¤����߶Uu�r�>�5�!�=�r>J�;J���\�\���>b�"��q�{4w]��]_2ʛ}�ϓ֔�����y���^ȓ�h��f�ry�ӷ��f \���g �g�%�M�Z�B_m��Q��� ��'�= '*�8�������z݋0��^�������a8��Ăܘ�:�� �l@0���@�/��p����_5���X�B��!bf52�$������k d��m2�����Ҳk<��@^i�N�<�D;a� D�֞����0'�-!�K_�=�{��ڢ^�a�km�>�s{/]١��<�����*Ѹ��_��gL�o�[8d�X���W�C�m��٣��t���z����MN����{T��B��L�9J"���}�{0�W��R����q��������������D�A3�ќ�iS�<Q�qH��ɚ.�)P��o5-d�R�٬A.�Υ�����t]'f������� ̂41Sq� b���$�� �"������>jj���r>��Y���y�<\r�I���W9U�J��P*�Q����Lne�[ʤF����ݪ�$
�c4��/���/>`�ku�,i���mӃ�3��Z����ᇞe�ϭ��7��=��y�v�L��[
�|f�j	��r�d�sx�K�{���]���˸(�@P����fY��w|cZ�9��/���uF�o�|'��-�����B�E��
:ПN1��:�8{��협���7Mإ�M�v�zm��ǻ}�՘���ќ�h��q��F��A��u�EM�=/h�Qk�>�jZ����0�Q���#��z��6��x�JEt�M�@ި��=k���DM�G����c�Aۻr�\�s���e%g��y�Z9��%C�Ҹ!T
1�/���%:YW����l5�6C�qx̆1��|`d?cm{_����䮴h5.�[ ��ܳ�;_)~���'3 `)ϳ�r��2/��_7�i�Z}����ik�2�Q��֜0�r��ɩ"�%��t
ˣ7�1"��aʦrg� G�H�/ӧR��y�fT�6��ξ�l$���[�`:��_tu#O�LY|�`ێ�����ʪ�4c��>�1)���g/yM�zu��q��o�O<�|/w��UZ�P>�`�ȋC`�B���|��m�V�s�����'�k����,j�"k�>f�nփ���Eq
���G��՞j����v���k�O遻b��0� c��$�,0L�{�ƻSy��z,��d��-s=�ȸ����&o��$��Tz3S�7��'��ߙ��0Y�C[g@`� ��B���h��Ս��Y`5�#
��D-}��.3dF$ޖ�O��e��4.��%S���v]P�w"�>P֪K�>����(j��aG��au��R�h�ޫ8�XYS7f1(�n�{��L.�QX���h4w`�r�	�X�T�p��H��$�!o#�D�\���8	Dw����c��_ܻw�a��l��~4~��5�2Ә*&e,}�=`�ok�k��5�X�WZ{Q��9�������E�3�{B������}̀ߩ��
���[�<y�5�@y�9
�c�K���̜��R޷S6��B�X�׊释�4�6Ϲ����$ewFc
���s�5�fޏ���J��7{�#'��������Pt��ܚ�PG��PqC-�^N����J0Uqm��b������:�6mr5����ԫ���Y��wT�G��ѕ�ԻQ-�ȵm�݈6�\�X�^���j^h-��MD�>Q�40 �P�X1VG�
 �����|�ϕ��󒧝����~�f�B�,LȘoi��^���	�[�|�;.�}�ѝ����
�K0♄�z4��@�q�����i�|M<�x=��5G��ۆm$:0)��Ȱ~ڋ	��Hi�)�_�|������s�ȗ��CD3�����Y��������hM[�Eྶ���W��f}4���ؗ	����$l�
LH�����4z{c|kݖ�\m'�`����(v�X�c_H����^�ɂ#�=(�5�z�k h$�bn9�0��C�����{�Gy��a��L2�����[Q���2��8f�	����A�"�Z2c)�B��/v���ފ����%��}�"�j�\�[ �=�(͚�C� �	��-�	��ׇPd��UW<�݌BD���ƅ��g9'*e��WȐ�Ck+m���z�Sd'Xݽ�>S�wm��X�W��!b8���
��@�zg
G���g�
�_@v]�N3��y�DZ���7��tI�w&}m%�����~p���B����	����e���^?7>������f��M�*U[[���W���V_k��w֩7���'K�)\�v��{�sb���kj��c�7��pHQP�k�B0В��I��F�����um:�(rJX��l�vr$�}����#�����688R
����cpP�����
���B2j&J.����Џ��BW�� T�(���
( ys���~���������@AL�p�~�P�*���H�=���[���WcX�g�q�폘�)�[ϖVY'�zY�.�9͈����(_�����4C}�k�A3��	�z�׷���� O61Σ,rZ�S��ee'kɂ���#�))�vq�����x���SH�p!(�K�N��1��[U�������^��!���( ѯ]��W��O��N�/�m<���4���vφ
�Ӓ�|�ws�k�.^���k�y>%`o �ډƋ�z"x�%���d i��]U*���>��B��#��zq��hN�	;���5�-����ي8����4���r�!�&�96��ݔ���L?W ߐNECˑ����]^(0��q՚7�4)�ڸ�D�C�vsݰ�N�hM;�;�?0��t*l4#\1}���9�e"����څP�W_گ/J.Pk X�՟�ʽ�>�>���M��̸����������4����y�`b��� ����l�t���|`%�;\��������9�����ŮɂVf</�:ȕ"��v�/j����i��=�A�G��^�.�ڔ�	˝��.�vas{J�����X�}#��A�Li�q�/�f3�Beh#�n��)]�EH-�������Z{��(�M���4;��y�R�`;>�	PZ� TZ��D��/tR���ϟ/��������|�]7"}��T'�I���oz|*+��L��Ia��m�u̿9� E�5�`B�t�I>6��a��i���#���p� ZæD�s��O���C�g��s>u�L���丿4Ȇ7~� �t�@G�:�k:<v_�n���$\�o;�0�)+����������'`ʉ��W��T�s5�������!;�c�7���*��`�c'4"y�uϮi\�5ey����Y[Π�y����~J��C��`q�}���0&�u݃9��t� ���(���R���5`�~5KK�4�&�s;��s=�D�b#�2J?C~��>L-���]v���#���~��7�P���(w�X��x�!���e��K^d{ʚ�-�]�H��D��,\�(�+�S%T�֬e1�����F�v�c�vĐ�
�����Gp�*���3{��@ꠔ0p�XJ�	=���dn��}�~�Qp��)҄s��n�0���^n���B��n�㞋��v�7mh�M4�|�\�T~��+:�n匨���a�%]0R�3�z�~T?oJ"x�s���t}���=�|2�`�\by�`���+(����������}�N�A���v���z�G�^�|�鈷=�7�8gp<]/%fm�z͍���y�I���CFa�PR4XP\�`�**+�˿o�+�0���o����=��;2+i@��� �w��v�����˭�4�E���!�x����o��2����i�u�MS�|�=IP�j�mm@�Pׯ�h�]��t����� D�'�y�Vd0:�;v6�����wR�fg]�Y���E�5|>�ns��?�餧�% �Of��o9�6W?�q�[!��z:�߬P���ɮme�����Q!DI	�m4u"g�3>Lsm3x��Ə,&������5�cφV�oc-��7t:Y�6(=r#�dy4���7c+\�z��]�tK(u���Ƣ�W־��)ک���ר��[�����rϘ���T�|��E�eⴉgP�c�3�T��>h�:��hk���!�2��3x�'�'�P��gVG���M�{-�MfA����3�Cp8�ɹ���Hdz�4-;[{=����/����'FVq�)4���۹W���><5�����/}�s�9�t�i��X����/-���G?�5&���t�r��8�"���j*���Mwq޷K2���pw�6�5\��F��t5X!�j`"H$�m�c\vd���}b�#&lν�jqU��ګ���aV�R�A_Lz���u��i`���w8�7Y��*k���^��I�}+�1��#Q(b�ѝ�ѝ�d>&1�w�����U:	Z�~�oD�t�x���+��������U�гB��_)��~Gw&Y}5�z��ibZ!����N[�MiZԹ�#�^��\��v*^����#���|0�q�nw�Gt�9l-�9c�Y��������i��Td,�}d�;���������3��N;_�"��T�ܬuM���6sE��d&�&�Vڙf�'r����+}�	7�W�n\��������9U�qJ��>B���v��?�����w^1�B�M�9��Tֺ�A�TF�tg�����z_��0�5��W��+�W��A�\3�>⫏��sA��|zj�l��n��y#Y��w��,fm�oHֱ+0��KA��q}8����!�;ې������&_R��4�3kVķ#i�
�*����t+a=���׀�>*K�qduy���42l�K�]���U�(M���^q>UфH���,0�� rb��	��ô��ʮx��7��յKd ]��[̼��mp���Gx��a)�4{Z�Vt�r�E��v9�uݏ^̊¼^n�EƆ%��5�۵Wr�7}9svS�g���7Z�Cn�,��єν�s}-f$�uʦ�ۏ� ��מ6U}4q��[���ډ���������Ua��U,q4r-o:�[(������E\����������P��ǃr��7oS�����<aC���(�Z,p�8y��9Ɂ�c����|�mBn�L2�P >�s8�?�`H��QBcɧ��]�c��`����1�舙�|��N�ږ�:�Cy�N$�v�a̛�)����o����w�by-���y�#��u���7�u.A��Ƿ�@齀��}��xy��VyH�+"Z����@�3	5��7��A�}9�ڇ�����{����_��w	�
����������sf1����0��e4����h��>�"g�i�������+��J�ـr��~$�(���Mї����å�_f�Z�~�Օ�;�ϊ5�u���]�kB�]H+޹D9�R9�*g^ߧ5�i>�uy���G%�я���s�v��������!���h��v��C�!ur�<���f\5Y�2�/�3iÐ��|�-ܗ��{X�E(]x�Ծ���x�sv��$$��n�wm$��=�E12A���3�8���G�7����ެO;��g�:����e2.W.��$.zv�-|�� S�;�-�����^�;��{v"u��j��ʗ�B���ⰸg�;$ƭ���ݼ�/q�us����sOF�QCP�,�)���]o����8�Ѥ���L��k3��ti�y��hCƧ]_,Wg���҄�̿w�WпC����A�����40y���23��sܯ�57󽯠9�6�>X��۴�Oug��`ދ9=�ы]�a�8��OݻY���1$���!f�c�����6�-wB��P�0�7\N��x��e�؅�"9%��#�����{n*%F�V��z���{�@�i��!W��֊�S'=���Vގ}�h6Gp������Kd� �d�v��͚�lo=N23_��+���龌X+F��7��x[\.�`C�&\S����WŞ_3q�qw�p,�%�a�z�k+|&x?��Q�h�{�#ù�l�ż`���&p����8���"E���ڗ�.L�LO$�&|t����� ��;y�ܧ�^m�t��s����mg�/�ϐ�|�Q��/�Zʃ[�,���{�Y��2�Y��L�F���'���/��M9�^.y˹�H���f�D�v:�C�cȶ9�*�{���#Gk��亮٬�r�^�zy�_J��G�/����/ ɷ�0��6�rI������P���2k�h�j�"߱n����6[�/sO>�n�����
���ebq&8u��|2�J�s��ٌB�_%��nE};��+q��OQӭëuK�)�>�D׬;x�̳�]��j�΋ys�>0��]��bn+A=�jm�c�M��D���&���$��㡑W�[�[��8dGv�v��/���k�9���1��}���*{.a$V�e���]�$(�O��ݬw�I�;����'Z���h�NNx�&a�7��$3��n��9
�d�4]�]N�w;G>w��=or��Z�o��"U�b����a	i6�Մ���	{Y�v2q|��d�C.���[s+�%�TA���z�Y�2�&q�$�s�̻p�T��8:e��.�(&�.6�2+ �y�5ǚʎ��.��D�J����ٮ�9FԬ�-�{�i�ԀSs��v�fj5�a��<<�69����J�9v:ffoU�ӊ�>�-r�N]֭Pk�:E'��¹�U�vU�۝=���Ps��J�w,U��;�a^z�$���Ɵ*I�*Q=���npf�K���z_JځR�=��흤R�'(B"b��`��|��s�B2��>������f��V��C4�o����֪"7�oEGkW�i��1�y
���:�y]�c�OT%U�r���&B�T�kb��h�ǵ�����C5%&�j� �<}V�<\�,�LB�oI��!���4Ϯ��������&�ؖ,c��:`��O���H�q�E,���p�B���"E���)�d�7�y��TI������3.96�#u�^��)�iRje��q��4��r���D���O�̮��s�l�5W{|S�5�9��n�R�����)�ƷPΚ%:;O^���rڭW�,���7$�Aj�9/X��:�;��ŏa��#� �o���*Ƒ��w0_N�T7k��}����wnޖ+�N�Wuuj�9�Dfr�����ؓ,g�uwi�I��c+q�I��T�;U+�����:/�w���r.A��s�
�˲������]�+*����%G�$��v%���C������eDӍ���ʰԄs�7�R������n�����v�:�y^B�jQ������Kxj����%���"���v����U�Χ�K�(F}TN���r�os���Y��*��ۯ���؍G.r�� �]y�g@5q5ktQN�
)\���t
�Q����2�5�_}^Aj-	�j��uk;]X��4�"�;=�s��V=k�]��u����.�������|"���ΚVܮ��*���:��b�*��{�plG{�%��㜩��:��j$�����*$H�#�y�*ȫ!D�Z�8�c�N�m��Ǐ����o�����������SH��&/��5():��ϧ�`�߫�n��$��D����:v�<|m�ޏ^��\�!�Q��T�]m�1"!��)͒E(��(H�FZ���+/�AC���׏Xӷo��x���m��8��z�8A �;�K��I,�]���JYcKS?�)�5aF��T�O�t���o�<x��o���g;�������r/$Q:p��w3����t��,T����0��+��������oۏ<|m���X���*��
�RBUe��F)4�*��8DQr��z�.���Dbf����S�v���޼x���m��\�T���>'(��H�:V�(�Pй(&��g-�Ӧ\�8����u�y忽�����';�f{�(p�J6�I��!,Yt�9y�H�\�.�z#�J�18R�����o��">���+6��iE��_-�:ES��$�2,�Y!!<��'<��>�'.I/<�]�⩬k�]��(ꊈ�ǒb�9F�d↋6�ѓ�7kbi�� �'�W��|	��?�)�Q�|v��vT H�>����|Ϭ�	��3�ƀ�����9	��p��ϙ�8OBD�-#��3՚�_/d����TGI��=��"����~X��:�o�e<��!yk�uǄ[I�\���)��K�U�S#�}�p4�˺�vW"F@�N&C�J���������
�"��!lq�PA��7ٝ���_����_��V2/��W@�BQT�Þ��v=����y4u�CG�/�~RZ�_e�o.$��E�ܠ��_BB���%|�ü4�sU�O+Q3�}8Gx�ދ��k`�.|�q�Kڔ��a���#�LǠ3Q�_IK�.#��ӆ�q�A.7�}-ה��1�r0?��|��kv
��*�9E�b�O�h8W��4��N�#}�P��y�W5�����,�:닭��;pº�p�ܣ�.:�)1K/P�o��Ƿ\�	�/R��Z��E���U�a�գ�J�g�O:B�b���u��Z\VJ�c|�K30Ѯܚ崟w6�tX�/�JU��|'��ߌ�Y�|���P��zi�����r��bs�<Ⱥ�����+|�a,��?9J��D�ڪt��V'���`��2QՖ�U�La����3HzV�@� Dx���aM��j>��ѝ�}C�����ַ�����4�^L��қ=�-f�Ls��kP�/t��'�� ¢P��C�P� ¢#����;������эfQ�#��9�DBL.93 Q�Q��.�1��Q���������Q�7��9Ks�g��D��ֶ��x}+�^���:D�)h�Bmf�| \:����`;mm�~Z��6�-�g�A�`@�1�-lPoOF�g5W�q�ېN�nK��ښ-���s���OLI,�.@e}�$�?j��ԝpً���g�4�C}6���/I�F��=�g���v��u�ݵb�to<�d���<�%���m�����	�w6�i�I�L�Z�4)���c{�G��l,Z������kJwe����x���Ln��8��������v��&�ɛ�v!�P�F29p������gc�C�y��Z��)��=1�U�]�(�;Sx�/��Ty�G��I�n-���S)	\��wud4��s���������!#���'�%��w͞=��&-���3Гe����F��3V�+\�i�����'���y��5�HB��_���h,�����˞+����A�E^��;�.epW���I:���Gί>��0��������M�ݮ9�
��s���qaڊ��̚�[�wvMD�T��j("�-,��6�ޝ!93*v�)��#Osa��֚/Z�AY&G%]���+�F�}�	_A�f_#�<	qꂉ��m6���%��m1�j$�)F��F�����8x>#	��2j#W;���������խ�Ke2�}9kig����}{Pw�w���n��`E�q��f|����>�Ȍ�B�z���4�F9m�4���n����:�K?@c�dS�"��`3@��";#U����ݺ�E�k��J�Ås�G�l��l� r,�I��c��޷�G'7h3��EZ�ì�9��7UQ�z��m�׹��ٌ*uD��m�*�ֱ:�'���ˇQS����`�
�בD�O_֪F��g�&�A}ў�6><�y���:��B-tٖ�p4���z���4sS�.�/����.t���Qnk4��ń�m!k1	�2��Z�1Dv�����R"=x������,"��)|�{��\���4wߩ�Y�ײ]��=����(��D��n>���kL�&=!�v���~a/+��N��@�+�R�A�L�fk��]�f.�7�0�|�u��^Î�>�f��:�d�Z�K�p�{wy���R'\���uƸ�Ϫ�/���5܍f��n��8,�>�v0�K�v�R�д3�WA�����]O��#�t����N[x���75�;-�����^k}�M�"��A���:��/�c�E\�U�weM���b4�uv�qIb��*7��o�����k�
�>��}vMCC5��x�G�����3���?w�
a�L�$��P��"�6<�D�˼�.g���ٗ�xB����s����H�1��`�C\L_H���ʃ�([�j;�ĽtN�H��Ǹ�޻�Ϛ��$���2;�p�{ֺ����|%u�ESg)l�Y�y;u*TϺ��<W~a�1</c�=o�������
����KY��:���l]��z'pj=ݝ؆ճ��O�(���^;1�Dm��>^���1�˅N�a���ؿq���~�91	��nǶ�n�g}���\�]�B����'L�#.��]��Gw<�Pof�ٱ[��q�7_ݽ��q���ܖِ �11&\�S�Q��>}=�r7��r� '������)v���j�rS>����q��=��k�X6�7u�>����"�ob/����v�.s�je2o����1.�/�:E���z��!Q��©���k��z�iA�a$���6�E7yV+�Ӑѓ�!P��; v���<7X���]N��)�D3e���D+q��-�coH>�eK�o��RJ�jĥIG^b�j�L[��Y��n���^ڷ�9��w�/p�k��d+4!KT���7���~|��7}Y��Z�)z=�e@��S���r�p�A���Ѝ�ލ��ceH��Ϗ�Sû+���Q{��-^����5�ՌGh=n��M�����lQJj�n]t+a�(�@,�p�7���7�r�֟C�'}�r�pu�/$�i����zE?����=�O�����Y,��L'�HuL8JC؂�6�w��O����9UM��!d{�����
\Ʃ�Aֈ���w#�j摩>��2�س�`�1��<�;q#��5�\�q�3{v�[�^C��ms27��x{��	���/ٴۂB��oyO��aRX��5��N��S!u3��$n��7f>�w�j�{o��������W#��2kg�S􄪜%�sY�f���c���=r��,y�`��Wwl{-t~��%��w!�V���[���� )���Ox�|�=�N�J���sS���w�(:�~���X��[�a�<#H���xQHG�V�2�!׵�FI�*��^ia�0�pHLΛ@T�'U�Ì`�A[.��1\u���e繿5S�\�����} �U�Pa�4�3I/��-ν|�3�>�Qs@M�1'ȷ��c��3+�o>?f�:�A9�{�S1u�ru��j����PhL5�M���n.��:u�N`�}��g��$^c�����C3��A.N0��5�.V��9̨���h��$�8�G�]?D�Y����b�.�]���u#v�+L;�z�X4�w�Xn�4ES�k�v�;��e��}���������*6����N�|��d&����G(��Ѻpkafb'ٲ�W��v��ֵ�ny����j}��y�����X!g��0^��/c�+�Q�	�E�w�ezt/NUL����w7~y��N��e�[�����u�R�s&�;����:/kloKΓ/���n�9S�Y$�*a���d�<�9I�ZCn�D�v2.D��f��W8Q��sb�}f�w�O�b�XǠ`�������zӺ3@�}N�n.�����v����I��&b��`MhI�GC�ʼ���ub��Pd��]��&��Ö-Pý��1&�:@�#m��⫭���Ʀ-�R�3�X��*�bmѽ�ކ^�M�����-Ə���'I��
2JTy �FI$�q�|=�	 G	!2���7�ؗ뿾7ߨ"�L(�L�$D	���&d��׵��vS�=y_:��l�u�!+.#��tjy}qk�'���$.����q��ȶ�C�<�*g�Uw��7wo�j��'��<��1�������T��{[$]MT����[F��*���aOw��^A�|�M^z��ݴ0ܪ��л�旋�I'�ݼadgz�j���7f��Q�]OAp}B���R~泑4O�sX0lRVn�-͍Gt�.������>gۯV���!��ʾ�ݚ��ژm�J(O;{��G-� �]�7}!��(T�NRG|�f'Xpy�X�#e��s�i�>�^h͓��2��g�f��N�A��p�kzu��2Ӹ��L�x���T��_6Ӿ&`:=/[����*;e�8>�'2�û=�͸��.������WDzn%��j�ۨN�B�լO����Op]$��c��XY�^�ub��Saf�R���;���5|Y�ĽN��m/Z�.�� ~�Է��3h�3~�r^n�֎�=/��Öo
��YBS
����6�Ut���Չ�:�8��S�I�|<@#��G�,}����wp����)������lO���Wu\���"���>��'�LOU֠�D]�<��v:�r�	���l���P�A%���E�/č���l�9���bĴ�й�S�U��{i�=T�J@	5�h�z��۵�ۻ�z���mØ
�bo�x_L��c�M����o!�����D��pv�`���������t3��TyEsz�,6ӊ�����u�Z�CC��2�g�qU��T�7��}���:��,���C^6�z���H>�X�K�t��N�^���gї�j��ڏC%Q�ޚ�����xWvM�Ԙ�yS���;
9Ut�t�(��-�$�Q%p���ɛz( ����Ϯ3���Y�����W�5i�nj��6B̼5��^dڥ�h��ݎ/{b�{:��f}w��=SvB�֜y<զ�A��%�.�Թ�qpV�X���K�<P�ܳ�:+%8n�Y�:�H������2*{�7:��&���ig�x���;Y�}�U���ʫ�FάV�� �"���l̹+�m֡��sh]_UIL������#���(j�L�|������Ϧ[���?����s����W�ˋ��c{x�ټ��J���tb7�
As��%T���z�w�N�e�����m/i��/1����K�2��_5Ő��şy�v���^�����=L�]u��-�ib��Nd�#4S��6c��q��J#f�y�XĤ��OE�=�����$�@b��W�{���ݛ3z���V�=�G�������ċ�Bw��k،�oNj|�)	S�Y��8�f�r��]<��kU3ץl6x�������y㔦�F��������2�:�􉮙}T����E��
�a^x���4�t�S&�Z,3��n����Q6ѕ5��:���$�Xg8g�u�ռ�1"f�YC9�u�:�wA�(nz�⠱7B�_��<���>��3��w��)3;ú�B�\��ܭ�s+�8�ȵ��{-�O=Rw�A2�_^v@9'�u��������7wQ���ԝY��qRҩ�;i���!�X�����$c�:WR���S��.m��]3�l���"i��NS��� ��<H�#��o���+��o���om%��0 ��	�|�aN��&h̸:������v�J�Rn���~�ܸ셒)'��T�T�Ƴ�����f�m$�kV��t���|��}UE�m�R�@����߈^��O���V��&���5���^�}�������#eK���úb�㪯;��<��K�ݹ�z��ΪYV�=���m"v%U��-�@��L��8�s��ym���|aS3�����V��T-̅��)�θ���>X��vs�=+��!�'6�R�H�3�ٹѰ�6�;[P�r��N�^d��f��߽|��~�}}}����Ogo�/�s̙��x ��u{��s��3M��
Fgw+�N�08�����{�x�N�8՞�S�=+zS{��J:����e-��9}�ə�wO��y��,�	1ϕ����k���@́�v��S��6�����Q�v�����pi��F�� YD2���Wr��-+��u��k2�[�Z[xj�0�\��w
s��H_'x-d�����Zם�*Y+�.~GZ/��rgh��u�M��'�����5,"kk6d*�#ת)f�ͧ�)��e�0ݭC�d�wv�Y;�s8��k�Lu�ܮ{��?C���%7/b��հ���I�*���U��3�>���Z����Q"�U�v����]�k[�m�oN���v7���T��V�y����qǳ��﯑x*S�&��'u�T!�u��b�]�U3�3�v���k&=
�{�쎩�2>흂�V�(�^�7G)�	�i����ɫ(G+�^��9{��ӢEd
�Mj&�m�)�9�gW3����s�}w�6�� k�Y��f+�&1�.vi�#����\�ۜ�ANuy3�M�۵�I�s�q�9z�ۙx�[�X"&m����B�F�d��,��"+7{PkC�]�sn�e$d]D�YlY[O��^he]`)$+TU.��i쵵����W ��:�u�Z��Y-����q)��6���6�L5}6��wwD
��U(VWc�ˌ$�r�nHM�*���z�0]���ff
��}ڕӌ���R�D���^=�L�GRu	�ه4Mh#���/��ӱ�>M6k��	4ɸ؈�.�J�T�'��W_pG}�a��j�l6+�l2E.���#�/RJ���9T'W�����!1�n�.�u�vݘ���g�����2^H�o���]�ё��Efc	�";���A�G����;Wq(Tؤά��Uv��;��,�ge�3�e�� }2$3{>:�C��E�S^�׆�	X��wsB��Vu��˄�vc�(���^�z�2��6#�N觷r�x�e�0v�H�ys-��U{8�O���]�ʬ3\�ޫ�p�&Sw�6�E�r���6X�7�ynZΌQ�E�L��r�#�#Ӎ��/s�C�a�Kc{��j����.�^!J�$3�}�\�s��Θy�����s�+��61�]sח۫3� �����$
j`ܓ�n��`*�׼�NZ!ڜjm`�ëD�7e�9gq]�kn�%D5�8)�oa�j)���q�su�hC��	Q�	d�ָ�}>��	�@�Cճ�[+WK�}s��0j��L����U��u0e��e6���x�� ��qx:��)fR.�=��i+�3�M���Q�m�\8���z�+��ւ�I^��Z�^Qꎓ��t�$��:����@�d;Wh�X����X�b���'kN�}{R�Г�9��(�Ρ�������5FblT���`��y.Q��A����L�J�A,��K��>�m0��W	BI3M���K��faf���6Yj:��[H�&*xJYr0��E�#�n��B�n"�N�<d6H�NJ�>*��s���d�[��(� ��9 ��dD��"F�*Do�f�+�6���g	F4$��C�㾧R�]21+8��@����h(�BG���7o7���x�����z=z�>�ȑ�I*$*�Eq:�!�Bxp��S��uqBZ&e���}��y�߷��zx���m��c=I�ey*:���C��X]Ǯ�x��aܞ3��d$֨_+6��۷����o[�>6����1��d�J)*�Uc��!|c�iJI�E�w����`��>$�)(*�s�~��N�|v�۶�=z8��t��a�4*5��z{�d��U��>2�Sב�TPEhiG-1# J�Lz4���ݻv��o�G�X���܋$����ؔr��n��R �"᯽�B�Q�cѧN�m۷nݶ�����}U~�|��0*�����R��AF~]�Ȏp�=��/���RI�[�YUV��uJ�ۓ�G9W/�wVD\,Ȩ�ʤ��D>D,��7�#�x�ç
��J$�ӎwוDP�U�_T�����2�B�Y���^�Aόn����*Q>�sȳ�r>R��HL!4�$"4�Y�qkՂ�:�,oe
�}�,ΚwfV�\۠vWY��0M^ō-�V�����Ԡ��h����l��
t�^Uol�!X��S��T���o��� Dp\�y�MN�g������l8b�Bs��*`��-�w���Y�{�P�q]s7�g��ݑ4m	f�_h����A�f_���02Mٹ�!'��P��<j/���/��F`�[����C��Kd��:��>A�vK��\uCGT���w���n�I��&���v�=��]�+�t欫��r30؅�E��9I=��^k���FOGg��hgګ��7˵ÐO�r�ר'�9����@�@�Pk��<?\&��c��ԡ*U��cA�VY�3-fw�%��~�fw�K�-xT��D������ɪ��i��v�H�{#��sft�DKcU2�{���\g�<��K�Χzr9��AO�rOf�����Qm6f�n��AF]n�s����SO�� ^�X�w:-��1ݖ�[d4���S	� �b�.���06{�Vgg0`Uv��G�/ �u |�X �f����X�R�k\Q<��S�jeU�DRw2�q��w�lm�N*�����Ԩ%�2�u�Z0@ss2	��e����f�9��Z˳���x�T�꒩Ƶ�)����]�@�3�����0����#��=�a��7v���=ϹD�碯�lwi�س����Ǚ��%6�V�d�.:�oZfpZo��_UL$�[��})v+�R5:Y��7����i���Jk@hL`�o�}�y��D�eM;�dwG��7/��[�j�켤�*�t��O�ٝ��ͨ;�w*����q��UNVv�4����{+9�^[�->�P5w�1�B�'~��X�5��|��ij�h���C6�un���=���6P��]?Fެ��ZC?Ƥ}�Z��P9��4'�w��:��]���g\�����ţ��u� �����n�3g#z��,�Q�x���-;�O�9�C��8d�Syj�5���vg6�\��J�{�����~�G��{��q��<*ߺtS'� ���ϭ&����&Y� ��F��昘��Ԯ>��G
1�.v�TXW]��U�=����ܵc��ns�)=�toɝ{�ph���)MY���>଒èxą�Q���p�Vvc�c�wt�٩���fo:�ZGu���\R���X������6t� ADy >b�ku'�nΑ��{��휛cX^�
P�����qBM�5�ɐl�<^��i��]�]-x�M���,�`�Ր��IRݐ9�P�?���7E���Wv�r�e79���ε�TW���_I��+d=�2�
q�/�ݛ;�]�{O_b�~�9�Q�Wo�{׷�`�[�&�)0CM�w`�ѯ7Ɲ�@�(B��@�����A�o`	gs0$�w�&2�rsb%�qu 4`˜5�5���D�a"~���/7�U�ծ9�ٌٓb�y���������x�c����f��Y�{���z��m���}��o5L!y� Mf�=nہ�'=bE��:}ʽ�驢θ�1ՙ.jR�+�?~Q�����}���G�K�B���]vsR}��'w�Ϲ>���c�a����o����}3˚���6���n��{_&�-�G�e�ޭO��S��#,C/��%w	� SՍӲ�]��2%�n�o���<
���Ob��C�I�zFup2(�{o�w���1�Q�#I�IG��u������d)U��_����N�Lւ�!�9No}���un<��l-���GeQ���������G����=����f?]��(i�SqbȒ �z��d5PGT��oh˩���ƨ{�䵶�a�N�/�k"7�}Mb�/��b���]�q�o��~;B	��j��Ñ�c:w`X�AǴ�X�u{l���J�{�:�D�g�k�Q��JgSd�� zf6�F���a�C\{�9�*������_���pȀӾ��5q�	�޷�k0?/���O}�7\fH�9\]�J��Dn�%�F��5.~Y��H�U}��9-�4�y8Ɖ�#'����#��S@�7a���2kP=�{�!����g������[Q˳mMN@�T_p���f[% �w{���v�vݤ�}@G;@���q{�/�nC�_?oaQ��N6v�_g�rk�V����H�Lfu������C4��̹�]ۙ���w�`� ����;�]t\\�_���-F�L׵P��gq���r���EAj�ﶝ�M�}�>����*WT����&�Q2����"Z��$�
3榑T��4k�9�ۛ�{���彝�Q����[E�D��H�5:��j[��W{��T�`�n�;�t�s�F�@�DDW	M�$0B%���$(�r�89� p��h�.nS��y�왆�p���"���.��ё� m�l�������i ��H��^˶�WU�^7){�Rބ%s��)��� �v�'7 ^����^؀�Z�]�ݭ��$^`�,V�#��	��zkz�����]S�j�ڒ��\������@:�W�8����^6��A�a��a���U�vW�grS2*�4���?7�Ϝ(�Z�-�G��q~]Y�s~VG]?uA2��ۻ�{��^܀2 ��t@�5�����T��ս9ج�ܞ�y��NXwv��w�&:Qb[�B�킣#��	�|�W5�`�3ٓ���}�+�Չ��O�����![�����)��n_���d��5�{�M��kZdk#�9I^/ ��U6=�z
�k/��>�o�CZ�����󥣀�.f@s]�@g����"�x�	��������+]^�{�+�M��9���.���]ۂ��?v�#wO+��S0�>ܗ��s\A�x`�n(,�P���޾Y�f�[�"�]�2��K�6���$�U����s�̫�C�كps��vy�����A����n����*b~��U^�rݕ@����4o��^XU(z��5��,D=rĝ)k˅��Q��9uUtK���)���Q��]h<L�׉`m�U��1�	 *�J<����n���V�	z1�����=�"XِX���b���޹!;�>�Z"���w{T��.̿O������RQ;6mS^+��k���툀�כ������lu����}iN3�
�����r��:����:�?4y�fߛ�Y�y���Uwdm��S���l�߬��Y+����� �)6�x��P�0Wb��:�)��#:�<=�wg�쪢��G�^r��{��D�|]P/c�'y���{��\�᭮j�����(L3'����6���Pm-b������R���pCf
�����֥G]�l�$��V+��\v��8qs,l7��8�|���"�V*�nYE���������}��𬼂�,�3�z�C�0]1A������%]�76���/>�|C�lkcט^	˔5�4&�,���-��� -�t�м��(u�V��]ɯv'D���Đ$p��G
 �7����LM����?
�U׊aCCe��w�KA�4�h�Gv���w|�z:�_�n������oL發��H6zt���]�M�,�+�]�b�����:+�9���a�5�
�j�n����x������L��c�d�g�z���ݵ1W�y�k9CT27Aڃ1Ȩ��c���bK1��[Ĉ��kvoܴwn�9��z����O.s[�'Fⶆ�k�і_6=]����U{v��TzTd�&�]�����ݶg�.�!ӕ�3���F�)��72-�W�]���)˼Oz-�p�[*�3 yq��Q�o�Oh�y�%�zn�_`]��Vlլɪ����6sv(����n�;�f�zG4n�;[�����+�h��X�v��w��k>�����fsdsg�U	+O<vTC`u��U���l��3��� �>g1+5Z�6C� ��4��٩��{��<��&�L��`QDK7��3r�ӼAѲ�;Gtg*k���9%�OknCtB8^U���Dp��`��27�}U��w�ߓP*�ꐟC7@�hj
\��Y�.�����37�Qb��芟b86���^w]�hCk��wT�1�]<���:�"m,�/-O>���n�|�6c�;�o?%�ߔ-m��TN���:��G|�`ZZ�"�%��M) Fg��]��[�o��8Du�d��s,��@�$�^n��ݭ��R�G`^�·�!VԮ��ٔHΛ+�u��3\4�fE:�������B��I�v��vz�k�5)���ğ���f��f�}�{�p6
�n>���H���#Xg!�Cn�j�)g��bE�����6
��;��L��P&v�Te�=���ֳPw񔶴z_K.o��:����Z�k���k�����1��F]�V����gCI��f��vb��ȁ7%���[��&�;*]��=�;_r���s�t̗��q�۸>~���P;���ɏNL�s��tN���1P>��x��8���zV}ZA?C4��<Dh�ܻ���&�Ճ�Q�B[��D2��N�y�����k]<�����!}T���bbѾ��8olD,N|p��z��ǚ�7�#W�}|c�r T(C�MDP��(�b4�U0�aC��'�~� p�G� ��1l�=���sc�a�G�������I���jݥr:�&_CQ�總�Y��T���۴�n�m��#����7�u�u�f�[n����:���m��c7+StdԾ����@��(�W'�o�#����"q��rt%؆�2������Y����ndw+�����s^@��M>l�r��TH�K����{6�Gv��cbWN2�w���)���T�í����3u狀;[Ϋ�]"o2�D`�ә��/���&"<�)q�\+j܈xvg����bݶ^����jbR}P����|�%q1^u��k��6ȇ�O�`E�&aӑ8�WX���Tn�>���C����ar&�Ҕ��e���%��ԧ [���ߺ��f��CG�N��z@�\|岹��#2�u�8�����z#Px��g��[lGn��gc�D�˝���K�V�԰���UeBꢽ�uzl�"?N��hѷ��>�Psm�O6��Ql��4�]t9���:�lѲ��ub�4��@�4hr���R��ڵ�}]Vs�S�n��%��m O���na�#��y���wDtA��4��՗\��s������Ӗ^E$;a��U�E��t�n���y⺦���	�̳� [��i�4f�H��kP���:��4�7o�	
�e�3��+axGz=�J�r2�GKE�w�����p[�z�/�e�3.udxZ�	����{�E�]v�\����]9�꺠![�J�)�Qj�����:W���B�q����h��,��n0�Z������At���A�޸RD�sL�H���D�Do�����GJT��$���m�}˳"�(	��F���U\%Q�s%��딌��MFխ��U] n����ͭ";=�G����r�L�|(�~�CtjF����n��Q۾�nQ���`oke�DG9���n{DWA�8r�3{�Vq�]�4Y\P�ͿMw{��ȾUC�R��������/���#�߮�Fq麙�R���&�G���|�W4��� )vȘ�w$컷�z.��Awgte��f�\��������E�٭�끡V�;�8t���	ǯ{�Y�H�F`�s�.�P��D������b�qլ�Y"��������\2�/Mpʹ+�e��e��P�˽Ǝv7;d�e��wT���ެR���RN�<���n���ӵ�`{*��Gl9�r*�e����9������:��[�(kv|�I�Tt3��U�n!�k/�d4�[�u�r��۽���|5�!�Xl��j��z��pql=�x5���u�f�A
b&��2㷵�&�f�ʻ�m�ۤV����d��ʖ7�U:��V��2۷h}R�D����w.ۣ��D"���ps�qG�k����k�����wzo�#�T�!�+Z�v������ōjA$ױu̾Y�>���;Fp����+o� Fj�CQii˥tjD���K�kv��Y���ސ�ȶ�Ic-V��.�&��Ԇ%n�Wl����?��A�^���-ȃU�mǛt�C����1��7�e�ۊ���kz����[.��xv��Pqz��X:��ъ�±a :�:M#�ͷ*�O�ݽ��4m8Z+o)����vɍ�SC��	�<sn���X�g]N"�t��[�{�UWJ����ˑ��r�?^�M���)��nw0\���?��~�!C���}�����K�w��%U�uf ����5�ܡF9٪1�.��ku�\%�p���\�U�;}B�v��d��h���U��ל�Z�rp���!^Z�,һЙ�U;Ro��ʽ2
s�}�-ڼ�P��B��0�N��hjl��&[�un�"�+���w�m��u������V��g)���r�Vh:��h��X�9j�T�-��v;��y��|×�xy�%E�����yk{�k�����te�-|S�`���{P\{S��j"�ǙS�N�+v�>�7ρ�7��&mnP�J�
sG�������[����֚���wF%Ɲ��v�]�ܤ�=��1p����+e]�ۘN�sW=9}9+�V�}P�[���3{Y��j�u}¹�2ć�b�w�q>T^�ݻuo���vSf^�o-C�ʌLڼ�։���hT�-uj5�pL	�fc�'���쵁R�b�֜ܠș�],�0���db���nP�SU!���^��{v]l�F����{:��4�N�[�Oy_��V|���D����yt�gV���s���k�9�gwwEh#�:8`���l�CT��.�C�).m���6!Z�4#�f�$ �9�1���,�Ą����������r"��$_T�ȫ�$���:t�ݻv��o���������F��H�8�d�R,~����Dr��;�F�~x�j-**W�)�
~��������v��o_G�X��d�eFI	T#���եUj��D���\�����O��.��c��N�z�۷n�|z=z�<���?A�wS�T�㣢TQ�"���U�	$�Q=�/�s���&=t��nݻv�����1������E#�ҲK�˖��P�˨��,�>���2J�ߍn�o��y��m�m�����>z��$$	$�XI)VGHW\*�䨪�"�o^xuiUE7�h����kv���nݻv���q��bG$��J�ۇ������o���G�w��ʪ����D�h���=BHV}���Q^H���;-n�Q
$�H�hE~v�$��.UX}t���!dw���H�鳑G)�%���G%B��K
 �\�
�l*���U!��s���50׷��tR�J�(��xs�)_t������7���w{�a@l��$��.��k���f�=��{�w�׾�х�hi�L#��<�pC�oiT�6?�V��k�c��@/�Ϊ@�����ٶ����K�N^�vv�z[�7��!��/�C�i����i�*��Q3�(6�Y�c3��c� ��=G��%��[s�,�1V�dnk�껽Vu��_L���}�z}��n�Lc5��_()^��H7�8�̛��t��z� ĢI'	R6�Uϼ!�2�nޑ/�*��Aš�bi$�a`�����;9�7
4�W�~����N���s�O"�L�A�S�(��%��72#efK�ލ�f�u�/>N��g���ս~}���}����5�p2�'.�'h�VO��A�ίϚ���'CK�z�lYU���*sF�{�^�T��
B����e�*�����ΤOM�ݽY8Ҕ�8���n}�~|S���O����2W̖j�/���1��tz����Ro�t�j�{t�[��fF������,��s��GWg=���i��=���x��ǝo2(�ɲeT=$쉵 v�Cz�D)ʿkc*㪽���ח�D빚������h�+Y�2�����נs�M)�F����=�$kygu����ʟ��\W�>e����Gg�����%uo^;S��ݜ�Ռ*}0��sMw�8:)��q���{_c��u�<��F�"�<+#d�N�f#'E��g �3�c֡Md�o?zF�gL:��"7y�wcռn˵��~k��s7�zO{-w�u@eٓ�n�V<�v`پl�L�}y�P�V<ҦyZF:aq��˦Ei�F�]��2޽�Q�7\��f�u@�,̤356��b��0�;b/z��d�Ƭt�>��ז��lB���-]�[������m^���}m��[���N��I)�r��y'F���gp]�uJ*��.4�=z�-#=��潅4�5�J����E	���S@�v����I�8HV�ѫ�<�
�%�KO��8X"�}���Y̑���|Ӭ����dȓ�_��w�Ά�y]�K����� Q	\n�R\.��'^�=2[%L�+&�7{����E�C�h�w����f'�f�D�:��#�YM8zC�4�Mb�8�	����D�iܳ���W4�D��u��V�}i���*s�q��������
+���\E�[ՒN�p��XD2�6c�0���1��A-�a�)���
��ap"�K��G��<H�7d���{.p�G;�# Q0�Q	��e�$����կ�h���Z��զ7��i���Tב9��S�w����v��o ���)ܚ��S^�g\�%���t�&������E���퇌衳l3�����(�������ZƆ��Y�٤�t[�4A��x��j�3�m%UW�=	h����n;mE.0�iAu��<Hg����^�-�{"JV;Cy�}�V%=/�Sg�"��0n�D�e��c�T���	ѹ��C\��Dh�A����j�uә�[�G�z+�n��G��V6èfѶ~�l�%���b���3Ϣw�ބ��
�yG�/t�w;��2rȼz�W+(9��pn����	Qi����Vf��X ��q4�	�������m�f���ɽ��0������/Z��'�3O�=Z�����Bu/N�mfv�*{\����ؽ
Xl�z�TvY�y��S ��Ư�\�����uu��\��FU��Q�J�\u8��I�6�$���v"���v�ɈyM/+�r2.Wk��;��m�׵}�r#N��&D<����fPΒ�8���4�߫k���Y�Z��������_��e�o��K��k��1\����n�ٷ��"�_}�KClD���zluBR�[1ܚZf�xE�����u�l��XQ�M�{��Od��Cof+��7_��Ek�܂XY��`[��^�r��;F�\v�k�i��gpɡ�7�fa׻�M�c��T�p��&��wi���0xOF@{�2�u>� !�Y���l�5��p��a횭�ל�q�ކ���z��n��)���~s��z����'�ְ�)��^��{CN�4���x�9�e���a�������Df�2��x�m�|�ē�4�eS�3v�[�H�-ߴ
� s�2�O��(۬)��>��c�'�n���^OTĩn��fni�b�_v{�_{jz�!��X�1n��{�ڳ�r�Z��W+��zi�K�'�|�ed�2�}�]�w�ɛa��⸢��Ri�yX�r��¦���cuy*G�y�dKr�\x!�_ty��>�Ds���=Qg�RNw:uĄ��;U�V�SRx��L��-�>f�:��X�e��j�٩�خ�kݑ��o�m˸����G]n��^Ji��Hn,˾F���Z����&��f��Y��ڭ�|9+�͓��;3�}�0�i���Q�dn�z=<�ҭ��=�n��'��b�ؕ��L5ץ�ڝW��k���f;���w�wK�(�|��J��՗���aa��0pX���{����)�t,�C�p��	��讗Y���rp����J�U{�s��H.+�^Z�#sݹ�U+�g���n��	�!�	�U@k]w��>�q���~�m+��4�^�y��^���Z��frY���e�X����+\v��Y�Ev53�q�W��ݞ�?��p��:�Ts���w^qm�7ʅ�	z�ff�s�����;��� �6A�
�Z=;ձ�P�m���#�w��vD�X��E^[���5;���$�{�nYdt�v�֎Z�����-	��AG���^G����+ܮ�Y�SL�q��oW4u��g;]���R�b|2���2)��x#�&)�	B�P�$'�Zb�6[�i�����/��g@q�m�]_
���A�.���Ѿ���է�L�T��猓̝膘��w}�w�+%v��}2���澉�"�(���wM�^���g���fh��rn苜�y���9p7���ֽ������+ʶ����쇶�}��t��c��f `ֿ�%Q�ǟ��-ݗ��t�BS��+�;=���U��ԃ�Z��$tY����l��oG@�5��o{u�V��i�@Yj��X�wu�s�J����J���s��v'��Aߔ��������N�a��ߘ�	Dc�5�͎^d�3��m��anJe܅��RS�؂ fw�.��3>(L��'G�C,O�����ߐ:�[�}�&�dwK�����+ԛ-!�E�PK?-���1�9�����o�=Q��Ƭ��`5�uL�<u�d���5�ީ垓/�w�
�<���Wiw�Up ��Ԓ�:y�Er�vBj$8OR�ti��!�<HQ���hz�^׀�Um��:�;V�t��]1��u3�c�'tSwF�N�<Ft�oX�[�QWzq�$p#\R8ʑ�A���%%"dA-����)��Cn�!�<n�`�K��*��lTuӪ~��r���fLlȣV$������%��&�z���!�`��|�a��$�QW����r9�͒���m'����h��F�Ƿ,;p�c�2֡�tP��VOY���B��x���S/7��d���my��>�7���U״�����Tb��N[�v���.�����K\���J|CPZ��lpm��|�ɰ��/Ct�D͸Y~��?B'S�i�T�5�G�h���j�=�m7��Q}@�D��v���,N�x����k�ً�K"x�Y7{�I��%Ơ�N�@4v��c�g��y܈��%���ԫ'��\���'8�a��3҉�>��԰MW�rN�ĻR��qI�)�ӧZ�z쫓8f�e��,�[��ڈW)�]#z���-؊{�ncN��ZT���5����_���$����_��wXP�Ӈ�Wc�bR�G]ٹH�������V5�a���;|X�w��ipQ�Y� G����g̣����)���WS�{[k���6��b���wJ�v6�+e�9�gj��-\S��)��m*�H>$x�mB���P�̞�F��fW%̾W/r@��ϫX6���EIGmW���RGp��H�"�/`��[�mt�ٝ�i�6�'Na���-���LVZth����T����q+�}��c3z�9:��X�C3"N\�#֖�oY-�乼sV�{#��_?����̍��,����v���c�/��91`W�?`/{sO����]/Z^.Z�Gb�]�wk�cꝍ� Uz،Fs��ON��t�����6BJ!Dd=�֒��\�$!�7���E{ߝ�0�M�Gn;��j�@}a��#٤�$^��S]b���F�����<ۏ 882��� ١��hl���:����E�;S�t��>���r�<�@U��>7u%��J�]�P7$��_�S���KO��M\�����ݽ�֚@OQe��t���gi-
��]F�k���)!��칪Z&q�'��kR��y6�*���{{缏��*|aYf 6C�b�#�ތڴ�Z���z�7�Y}��M�Z��i��1�\ Q.���q;{w�� ��_0���7�Nen�Ga�3��*g���<޺$z��ƹ{�6������i�L{rmάg1ۡ�X;1��kS��Amw�U�{�P
�������m"_��k��0��lO��T�	<��*��|��R���鋚�N�k���lY��_|��G��b���>��Cc_�oiv��P���5�-SE=�n>�wv�bfb�7�#l�%�,�S}�̚
�uo� ���Ļ�%jUp�.��3����Ѿ%7����J|�z4ϻ�!^ǲ;�q�c���dP�iz��+lClsa�{���kG݁Cv��;ɽ ��ޛ�uN'�����F��\+5��@|��Ņb.1���Õ	�m_40��^��؎���ϫs76g��k��^z���]ŉ���}��=З��,W�9�[� �k���ΏK�ݼ�5]��<�����I�"lٺZe�f��]bYHIX�#��#+�^��Ij�\�n:��{^���&>8��s�) (��1����zWw*7x�wl���v`���L"Z'o��TZ����/*>���F���N���� $p
C&½I��]W�7��^�:���g!"�^O^|m��������]�[�-}�Ku�`i�ڷ}0�yf���ds��D{
�٤ܨpǝ��4����.�
�`��G
E�#{�&>״߽�@�{T��Wt��c���1}���TU`n��"�#�З�L�N����Th-��7�S6j�m�����դG�C��AQ�X�ݖQ��3�%�z����j͎��.�M�u�v2��m�Ƿ�������V�f��*	ii��}�.��z��͜�y����*�r�����jS�X�uE�[��Y�2�U��AĂh��m�-��@���I�oMl�mzO�W����q=[��������W?%Ei�?L����b��E`g�嗞���[ܲѸ�jX���ݻӘZ��d�d4��pe�K�����J�߿>�Q.��;ļVQ㼞L�q�AP���;�p]�ˬD�2�����UokU�̬�}��L�V�d*i,��;mB�oScس{�,goof��]vl͒��k�=�F��i��U�w�l�䐊���R��a���*x�Odt�KxV�bJӫ_��4�Ȣ�T(�[�ԮyӋ��z�U��wvf�shO��t/ڳ��]0-δ����~J�r��M�u�}vN􋊂�1���S��������K�V�L�b��Z�p��p��+��3U��OT|M��e��N��fd�k&8{�nܗ�Qɯve����IJ�ZjҊ'WF�p�3Ei�����n���Mf��R�z��n�ͮT�fGUz��o-�Tmpj�8:�B����f�8�����L��:�;[����n��v�MS�[�f��W��n�\ʻ��v��������9=�W.�����KbKD��y���:�gV�)r��j����K��	5<��I*�4�4,�^w�F�ͻ��m�jc��f��R=\ �3Y���cc�w���uד�̾��&tBޗRYN��Sb���h���A�%����.�_��H���ʧT)ؖ�N��KP��5XrV�1m�a�tqJ>�Y��ў-��M	Q6�	!��P*�9-���*�wy���Q�&�'w�ގ��YqJ���ӧ	(������Ҏ��Öj �n��$1�A�Y$���G�����B�c1R(� ��d`�k��C�4d?
*�E�Ϋ��m���&�ܵ���[b�{�}�R�6VE��[Ӏ��j�0A�h�`�^�LT̬�+m����aI�5-�o���ѹ*�B���Vd����Y��ZD��n�tY�Ԋ,*L4'^�Ƴ�$\�op=�V���z���yk*u�e�R�ۙ�iګ��,b�j˛�����pY\a�����`���_Q���޽���o3ZUC��!P��uC�J�t�j:�fM��2W?v��\�-Y��ta�ސ跬p�Ĵ�X7���՘��X���,s{��5��&	�G0�>[J+e��Vwa�r�<e�wk�Y	��S	���S���j�1[��kͧقZ��u%�ď5�m�RWu��qMT��q$3�-�{�]��:Ü �-�f�l�Y��ʙ�U��w%l�~N�C��}v��]ڣ\8h��on)Ǯ=2T�x��T������F��*%�����Q����:��K3]�7�3���׬��K��-X��}wd��	E�y�oZj��`�/�yꔮP3��V��B�ʕ��軦,û7x�9P��mg'*���t��b_�-�N�d�Li���
��1�M���9#��mCua�ZLUdBX��qv	%D�0�BF2J%�&���mR��9�C-��BH�i��	q9!AtDaPA:Q��FȎ��z5��A��IZ-��@R�&a�$�T\7#�4ҿX7f�	.�"F�2D*1�L��W�<���Bg>$3 ��8k����p�A���+��B����ɭ�U%K���/��;}m۷nݾ�?��a����R����G�"�_�y'+�I>Wj�J����t�ݻv���ǣ׬f�}��z���<��'a�j�tD�keB��zy^\��@�T�@��ӧm�v�۷o_���g;��{����|����T��yܫ]��Y��֗��J|�ԢFC�T�6;t��nݻv�����1�qIG�.V�\֙Q(=������M���������fA����h;�GX�v��m�v�۷�ǣ׬c���t~���-�XS�U�U\�L*��$⅛+"}��۶�=v�۷o��G�X��)!��QQ*��ط6���	�(���k����FRd��\�"�dJ'��D:�*����lQ���{��|���3G;�~�$z�Q��
�rr��PbaEr���<qx��(��(���D�I�	(�9E�v��Q�}�(�|��8��ɌB�F$D��Ut��1���td���A��mw_��;RW+`J�W�"��ZqEv�G�H��6Dzz5;_ﱤVբ�l�E�g��,���i�ۀ��7�� �s��v�[��,w����څ�~����qc��eK�f�#_E?��'�=�W����bK��>���h��*:گ{؛zm�j���`K�;F��͈�2��2D�4ѹ����yJ��yzg���4�=�,���y�����"���ֵm���8�l^!�Dj��kzqD_E�3m��j�Ҁ�ܽ����5��M�q�p��'�uD����<��]��X�s�%����+Z��3na� N��,S�����`�'	$��1U���Nl6�Rܷ��ec�h��[��̀����*<k�[@l�[�����j,OT�k�`:#U>�2�4�Y�f\�ꍋv�r
����X��s�>,"/��%�	��-3{Vnߥ����=�72GD�؉��m��os]�<L�����)��]n��SNS(�@7QĐʼ�g�y��/�<�v��Bs�����^*�]icz��f��2�7+�n���U��9u���P�z�O��5Qg�w-�L���^�Ҧ�.�	�W"{5��jw��R�8T������Í������ s�$`����H���f9�_R��'/����c����� ا�B�k��ÝŚ�����͐K��μ@���VAh5��7y�4�J;4�Fe��P�T�.��wQ���oO��8n#|�V�}��5Z�;U׭���9�rw�]"�������s �@��놛,��f*�v��C}�̄bY>r@kuϖ-�9a�+"DS�l��4	�0x�����J*���{Ƅ��%ϒ�n��ܖ�-��:v�q�9t*��Y�n�Kdv%�ƶf`�<�g;=${����[�ܧ3c!tm�t�*�]K]��)�#�`�4<�e��oes�#�ݵ�H8��3��ɤ��	��O6����M�˷"�E����d�ɷ:�Ts�6�a�WP�*E�݋���w������l����F���M~�دww��_�+p"b�ewJ}�[�"�i$��|�b�Ma�D��p�+���t�9�,�w�q�;�2F����rĊ����oV��6j���
���(κfɏ0���J���>�u��c��iͦU�ͅ
���%�V(}�o�=�m�-���3t����!
��}�L�����B���5h��N6�l���)^���s�9��R/,��pYܭ�YK9Q��mO�}%e�QJ���G���� [�e��I�e�B-���i�a��9�!��WU����*f��yy��g�ǡ�������z����Wv�mT"�o=F���DP9�-s���.C��O��2`D��f �{ʃ����la�íNK��,)�YOc��(�M�C��2��Vb҉�፝��w����7�V?��V�=��2���
g$U��::�J;��ɾ͚�j����u::��nmS�}>�q��3��11V2��;þ��3�xm+o��o`�w��{�sq>����y��.�{W���MN�t��C:�n:�{�%x{��${\�����C},������z<���-�يD0�k��U�K<sA�v��6gu�,]�UƟW�UQ؆^�x*���os��{s���@���_U<H�<���)R�gv�s�m�����3ν��o��3s�s�Ӹ2�pp���}��[j�xj��2̎�ņ���k�����^��uKQk.�hm�7�}w���� d6`vB��ꛛ�w�]o��<�uv3ĸK������_4LEe^>�6��b��Z�e���*nی�Q��1򛡢sc������|ך�択�� �N�O�[�F\�7��my��荓"�t]<��v�5�Px#�,G{�C>yt��)s�̇���Y���V�(�#�t���
�9���gu{u}(�٪��e����+�2���l�޾ၲ����@g�-�9����w��c����b��h�6�!�x4mI�,�d��4�E��pռI��ѨӯN�KU��B�T����N&z�L�&%������||��빹/y]+�{��t<c͏��X9�ð��+y���T�k�"�fe��tsAe��d��n[��HWg�$)�֔��=#.wWi�բ)�wgo	'�P�Yf�h��:�%�odF���.N�]׷�%W�C6�Y�7$���6�L+ �xF`�����xjR��JN���z��֠Sd"���˃=�ʿqq��l_�@wF�w��������B�;�����n�n&`�oӈ�d�F�hu����){�~����tݳ̵�C��;��M^wr��D����H}2����Z)��z�����j��'�s���x�M˸3]��^��0���\�6�kZ%�Qf�[2j���ݻ�wr=���.���YAԳ�΃Sπ��:m��Q1�Uۑ�P��:+����7�@9b�u!w��c��.df&�i1v]]D�nl�p���Q��ZvH$��f�.ͻ��ɕ��cu��tNlS\�Ŝ ?z=�� ע]ok���}�����ٵ���J���Zf�D7U�A*ψw#՜Q��X�>r��p֞�z���j �Z����^��ߦ�>dlh�?��[���8aհ%*�r��l*����̓���H���J����{���m9��D�vޅH���Į8�Q�|.��Z� �����E4����7mH$�^���C�k�û�f����s���2W"����w�[CO`��x��p*��G�� ����.x����rs�M�O�z�����Y��e��ݘB�ޅ�ڝ�<jwU�����7ok�me���c~�}�Ѧ�5>��m��}d��M캞�0%uz;C)���\��ϺF��;��]��[[����g��S��L�@Mn-�3V�h�v�]����E���UZ��w�A�7'�V��q6��4؝K9&�#i5]��t�L�\���q.Kg�f\�9�lL���r�Z�S�K�J�;:�-��I�g!��K	̌�7�uT�]L�M�;�٢�}~��75��;)�xY�ų�� %�vwT���=U�+�W`�>�uwi�꣣��H��<Of2[����$;׻�y{��ua.t�\��>ǰ���pB�h�l����|��E!�68�]X���[��wv���l�}�V���*�,��|��SC.���7�sW
'�(L�.�s�T��Zؕ����]�wZn�����M�|U�50G�Mi �NLn�DZ���N�]ܭ}�wVI޾̄Go�L���#�(7��/k��`�u<���m��n��V�I��zj�Mű�`��޺n��BH����/y��#UU~^v����d��N�']��;��h�S=�1�55*������pA����.��^|	�k��6�K���ۈ�Ȫ����Cd�f,�e�����ZO�T��y>SGA�k+8r��F6��5��b`�0|���c�|�3��C��-��u8�����2~�WGN��%kw�7���u
ڞǹ�T3\f��W=�����Kߤ�6���lg��y�;f<���� �n�ȥ�'σDZk�l��,S㽗{�yy�
�������r�9���"�
���8�XR$t�Ⱥ�{pk��b��{�Q{qCH�5����z4�Kt;�f���PE�%�c���`��k�r�[>W%�� �#�����v����9s4�9����3crv$�2A���$�癬w7`qKs
STt��zn�2�伄,�	���7�t�|�rȐ���˚ݿq�#db1��u��Ju���e6�ߺ�q"
#�f��_dv���gAG��x<#�30kˬ�6� ��gY�đ����L秼�[t��pfn�0�P4�2�5Bd��	�|�u��N-��+9\�)�Ҏ����L�3^kX�9��������k����J8���9�����M��W������s�����7�M��98�lL����U��B��z����h��8
��N�M�;��]Ra][Y�z۫v��y��իk��ovd�O�����G�Oc��yu�'�Gd·4U5�ޏJ���p5M@�,�V"�H3�M�ZV��v��3�gk[<�9:\�~��=�s�;�z�|�r��p ueP�[}5А�D�i�/F����,ԋY�}�V}��<,���o}/����wܳk>�xF���:�v;�Έ��M�n����ow�dO�5��a�5}7]w�Aqǅ��������s{���Ͱkt|��"g;�H���*XW�U@��5������K\Msq�n���$b��#k!��;���&�$]c9q:�+H�.���G�_��w��;��|��N�ni>a�i"E+���j��염2�M�Y�bVd�
��b�#,(�=�`v U:���M��,��2��=\�e&C0n��w!C�!L9 $2v�6��a sNݲ�~���^ٔ����->{>��iC��g+p'���x�r�Z�W:���ĩ����M�����͆Q�޿>I�>A}��yI�4_5������Vk���a�v��pV�G���ݓ;��Տ�w:�_j�RDZ{������j���4�}*��ـ�����vMvjgoj�٘�1K���%
=l�����7���3��Ƈ����'!�yw��B���[=�"���v�s�F����5��VuS��ա�3�Hj�䥟�%]�7��k�>�QD �6�:�jL��_eMf�}�m�-W�s����z�2ݼb<�W9�q�F�G'��4�D����d��'�"[�3����� ���|��Kk%�#�v�\W�XܶN���XX��*�e�+���έ��hawݗ5q��X@��/W4V���fr�h6�d]�A�{kv�CcY��w�>�(��㏻���H��Ǝ^>��*�;<����.fr�3��J�s`ۼ�m�
=�gi�,ju(n=�ƭ��<^ڸ���O'����r9�������ڬ�m�+1b�˷0(JdoZZ���"<:�wr� )��b1��A��5��G&֣�3�;n%ٳC�ױ�7��N����S�{������Ŵ��k��:�F+�]pm�������ϤE��ur����Z�y�Q�;��o>���ޮ�
\�x/Xǜ)�sעn S[�vb΄��9<���Z�މ�l�yv�T3�B!�?w���<����j����*��x�QB��}�v{V�\{1��6gs���|��eC_�]����k�dM�J?5���d�$�q��QZ��3v)j�9�t�@������E��>��.����B��.,��	K�h�a��}�^Y�Tst�f�2��r�>�>����y:�'��WG.��c��ol�����*�T�5�y-�˞0���;^�&�C���B@QY�K��y'��n�̕}�;�4_Z�l�B9�D�r�P9_L髋���h�M��SA���7��L6,渹g+��!���վuL��䆃Q��]�[�}yI]�AA�l� S�����7�����lZi��;���6MSoxi�ѴA7�S���W�ݰ��:�W�f����E�
�)yWZ����Tu�:>�l���ݾ�����t�;r�p�{޺�#q�����z�7:ă�O6���ה��oLҬ���P{.{F�/y$�!�;���*g_&��˝˙�Ǚ-tTt�'T������*�9�%���	�V�-�ŭ�w�fӃ-G�]BVڲ�J�B��^�oOt��ʇe�p=�3�H�86���h;ɹ�pq�X[[�C�gn3]���m�\YK�����ᩞNXe��	��Iv;΄�(�E�8���Kd���gT�)���\Κ�(�d�4o�xh�+�w=��vA
����5�ԍ�(��YS�]����B��L��VJ"��̦kv�2c�
���0��!�<��k�,>�3Pb@�����u�dC�!_�����Sӽ����¼�>@Yt=�17��Fq��N��:*���\��/�Sy�:�fFP$��}�^x֎[鎻���]�WB(1)ۊLw6�*�_{��T-ͨ�V�.���[ML��sC�����(r#+o�N�b�e�[�*���CB;q�sT� Y]J_T�y�$��'a{L]��>μv/��u�7F֋�`��x+������-NU�9��^^���"���Ѵ�������'v���W��&��VW��u�d[���[�1�*�PW�	ͩ���vc�xi���)�m�����]�^�y���>Z���V�y((8��y}$U̘h-t&^�ʷ�n�Ѯ��t���2�Œ��7&s�ĥ&�M�J������:ŋ ��v�ĳyd�oZޔZ雳yIΗU��{և�X�d[���$�kiO�.�/,�f���=2��ݍ����d)
��Fc�z6���1n:g�����u�&oǧ.�]-�
K2�G�֥ݵ�i� ���x)����	��3���&��ț�B��T�#��{������FMǸͤ�+p�HA]�aG�%����;��@�R��
&��ʧw�\���$D�F�h�&S\@��HtC�\��:QT�%�*�ILk�:c�ox�۷o���1�~�~}%>�S�.�1N����~�Q��O'&���x��o:Wr%5:�:v�ݻv���Lz=s!�,1?S�>��ό���9YТ*#�EPA�AY	�($�=z鎞6��nݽ{�k[�o�Z��/�r~t9Q7�ӹ�����m�Q�z�B����ݾ�<v�۷Ǭ}i�o�������e*�fQ�@�kN$Y�8��"J�T�^�cǏ;v��׬}m�߷Ϣ"���XeHrL+P�YUo�re�U~��0���Z�/��"���~ݝ�ox�۷o^�����̒G$�E$�� �����IE���
��_��Ay/)2���5(Ϯ��*�!�D$�c���e]$#��E	�i���aW+�JM��U9,YDV�'�8�IfҸDD*��w�r��Q�ʪ�UAL����k�\eQU�(;��>B�,����B����:zu�/j姁��o�mҭg�\CF<�����6;��hMU8-�Yv�o z��k��lC�����p	��;+��h��}Pzt�%1��;�+�Y�_}A:��5��Y/=�ω�j��odN�D��#z�O�L���-wVo{./��_��>�}�*�M��4";�������Nն�:F�<M�]ٹY��G�4ާ����v�a���?���F.�t�[����oB�\�r_�8�P�Ij�IUBK�/�8n��{s[�Q��\�uv�\iLb��S����޶�����1�p�!�1��ݻ�oW/T�I�0���j�n��c�[ܷ��.sr�i/V_�o(�F�/4H�yt��>V-ފ��M���#�_FzRt�Ʃ���&�c�v�u�'e���y�&Y�x;X�Zt�����Oq���*��b� �"�S���k����p��DQf̮��dP��NhnF-b��J��jWwggq�Hɭ��uY�Ղ�ؗ'vg+5ֵJ�q��:ޜʺlޖ�8�f�{L�W9S��������s6$����yew	;����mʠ��=�>��^�+0GX������]��4�� <��>0UJ�iJ>�ɮ��+��d�)��FoM��'Ҷlw]l��ȑԶ�wqT8�}%��V�y��5a��+��e�T�О�9������z83�m�����,C��,�҃Y��g7��ʷ��s�X�7"�7�j�WW�������kD��u�N�g�$T�5��$����W�yW����5�c�C�]���{��S>jT�9G��n�{����Źv��%{�S��f�<՛~���m���S�ޝ~]3��r�މ�P���U��w@bG�|u]����0~[r\�[`�ʋ�X�q��j����t�][���f�,f{S��~M7�9wem摭�3|<9�cj��s�[^J�y���q��z)ؑD�x�['X;I���wf�3�e�y[�������.���߇%��8}�������}�Z��{��]�,���U�.�=Y��fS�o;W�י�{+$�L�ɝ�W-����8��m�w��,�Ne����(Q")"�/]B�3���O~�H�����]S�\�B��Ⱥ�-���˃
`k[�d�E��`=��7/�5K8�ڞ�9��(��脘 ��f����AфHaDylB*�1*fC-�ʒ"�#B|0� H�P�gIIK7t�M�,�Y�{^���+��@�})v�t�tu2$`�C.�qg�c��T��&�M�S����t;�ջ��d	 ��O�K�b�bz�5�{1���6�h�<�+�r��a��[/�����������KQ�'U��ˈ���I��cWŽb��4��:�Vخ�74ވ�v���B5�y�����p��zI�#���ř{��A����_7�㲲_�j��'j�ݦ��V�Z���1�hFM�����<�5\�;�E�O��T����3B\k{h���Nǰ^����rddWKl[�rd5�Ud?"#������N+��/�Y��`�z��û��kw�n���+�2QD����X7\�ƿ�K�����F�_�S���L��C�G{�������.���()(��=�vY�R=Ց(���b]�j����W�(A��?^�Xč���ʕǻ��GS���O�J�l;�t���S�po|2��?c^	�������ǰ��d+�bo`������fLz	�	�=(�xu��a�V;lM�̲�׸�wk=ý�I| �#��z̞I$�:4��GVL��u���4w�����LHm�G�ou��rylY�����2���ΪxT?��.pk�-�� ��'���k&wq�a_w0����|�3�N2�}#g'�ʽZ��|�R���2���:�7��ܒA������yN8s��u��
��&m{n7^E�'g�Ⱦx��]��B����~`zt���*�htn����V�t�cq���ow>P�ؿߵꟿz��~���'<P�v���_OG��q�ٙzv�!@���5���N�DWiv��\�^"�5�b��o�[���$������|�aճ��oB�醈���qj�j�p�+ҷ<�Z�Ƿ��ܬ��l�߆������ǅ"NF���m�{���Z�����Rx�'�����u��6�wF屛5V6�uk5Ys!$�0>���.�Y��vsp��̬B���Ab��.u�JTV�X>���D{��Dz�O��Do�Lu�ι 9r����v�M�<�m�p'�\�ڔ﷦N�b��#�M��(����i{x��3��vy��Y#7��4r��y=�����0ZG`�C�F�r�d�n1UD�)x�7NԲ<�37�G?����П{��(�33�m�3i���P�d��5)�>��g��Ӿ8Ε�^��o��D��r_/��s�A�E83%�3gm᭞�nיmH��\ʒ�[��h�3��%�ڑ��͗�J ��S�w8��>Vck�&�	)���ʕ|�ym֩����X�qKg��v��4�F��@��]2�U6ݻs%��U����E΋��?wd�Q��r�t��v.*��b4S��X���"�ǈ�f!�!�H�$jǽ Wg0oY�vn�p����:+u<K��n\����� `�C�5��j�O��;��r�����q�<����\�T�ێ�n ���b+�|g`7ڹH�zu�����U��"b��ͻ]oqա����f�8�t�uo�s5.��f�)��>FĬxEBf�D�W��5�ދ%s%�ȕ���O�0*�nACM�*E[U�]��'5i�"�6�v-�nUox��aD��@� ���6qJ7��ZR}Z��U;}�����P�/P�^��y�2��\f���N��B~{�Μ7ez�!��F�T	��cꝍ��غ�Gg�����4���ֺ��E����6���~v(��P�ǚM>7�y^�uHܮ�Lq���!V���Q\���x���T�L�F��R7Րb���>�g�/U�w��o�|����_�z�~ݮS���S;�*˗��^:�E�/�i����ݓ���KX��{�A���hm�ۺu�[��2�g���^�>��*�t+��avʽb�����7��x`H*c�K?;�b�nܗ{��{z
��v�u�z9>T��f(Y%�����$�j�y��[Lj�Ѻ�f�p�'�o0D�.^�kw@�G�=�S3J��ZݮŨ" ��[�&��}Z�s�����(�b˛��:�O��މP�j��
��v�j&&^j���å�Sܔpy,k�`.OVU B���~�X�	�Tu֌�beq�e�E���kELBmR��*�y��A( ��3�N�DwK�BtRu�v�!�P��)�T��HH*�ϵ=�;�G�he�ٛ�c�'��q��8YC�	���Bd�$M�Q�m����? �ؼݽ�~ޚZ�Q@�f�9G��Ş�s���	~���o�.:Ѯ�sԱ��/�b�wyr����Z$H�g�<��<���9~ۆ1�W�G��N$��_�ٙ�.B���%\�[չ9Y���f{	Tݥ�S�ݾl���G��)hZ}}|���/�юf����<s��j{\��Gyp3ܷ�&�ը��|��Wս��ל���W�ݨ�erj*����0�ٷ)ߝ��es�c+z�t��.^:UV�Xx��Y;��Dv��]A����W)���?{�TCRJ��E_V�x�Z^:4�?�_{1���7ɚ�a�R��W[��(���Nk6����;}��Β����|G4e,�|�\[��l�x��U͇�%��.N����S����﮽�BP00n���*S�cj/��:�&m��ݾ W�vr�Z�T������ɵ��u���캷���{h�dw����+�e 7��?)�V�ps��n���Z2l�TZ�{�
Rp蘅���h"u�0����õ����J!�����>�0@d����G�ǑW[�J�=�3/ ��Ӝ�	���w29�[��l�j�aS�Bf�x=j1��,M���~xyY5�:9�U�z��D�����S��o��'��.����1/��oOt���.�	h�\��V=`5~�����nyz+��I�����.v\��h�qm��"��Ԋ=����]9
<�WN�qb	�fr	�Ez����
�!8oe�6k��z��暵+�Y����z�����4
ޝ!�-���Ϯ�}ћ�ȂO#�yܟ}���n����Ѿ����S����n��{"y@�v�in>f�?p��`]���
�W��azX����3�Wj����N+�]{z���5C���[���y8�y�'���ͻ�y�7X�f�Z2*iU⶧�o�1�]�E����X�������כ�E�9�\۱�r��qlA<�c})�f#x7��mv��G&��a��}`��uj��Z�V1��!��	�$��xI٘}`���IY�O^;��v���˒d�8G�Ek�GQ�:�v97��Kq|��˯9�/oķ�,<�� FF�n-E��b�Gxf�A�����1αV������Du�T�CeCS�փ�ՙ��m�&�[i����A���JT��g��B�t��@�s���%����o�=�kf'T�'��@��ZEC��w�9Ugu���'���]b�l����Ad��;'7�ξ�>�,����wW@C`��	�lw�K4����\3���̢I ��K��#W<79�l����o�A���׆��V�u骑T���u����P��~[���!l�ݦ���u�z�lt��^�LX���؋|�ʺ$�L���;�&ݐoݗ�rX��1.�u鉰aQ狉���o����'Ɖ��ߛy*V�wUL�q��w0���$�s�eDI��_"��̌nGa�Z�����yV%�Y�;�w��
�޻��*��a���i�fA����q:A�8r����9ͽc�8��&j<��FM�S����ƣ2�v\	i���=�R�D����ɣ^e'��n]Y��M��^�������mb���=�Ԝ{K�
}bv��ݞ@��y�oxc����JdA��Q�"H#�������~������W:�"3ag�uZ��ۏ�Q����"}[�â����3{������VO��$|�68ऒ��>c�Y��;S;�n�5ww(� O�5�z^�k2���Os�D�vOqA���]�P��V�������8��K͂[��.[��m��vڝ�z$KU����Wu���z���,'fb_Dn�Y������k�v���k�/V�웪��f8�w�G'7R�؆6�����9�D��5H`�D�����8�$�gT����C0:�=��kᡗ���c��=o�����ī��.kA�O=6*���v�W�q;�z=��V������טv�?bj]b�����6oGo��M�dC��B�����i�X=�S�ݚ�=��~�����%�R?�� �_�T?�����(��R��A�DKZ���^�-�� 2 �RT��`!EF��Q`�Aj�`�`�@`2D`�`0 B*@� D !AD)���*P! ! !T !5��C`(��"���ETFCt���!�!*���i�*�!P ! P !P !  DTAn%U BEUQ �@��@��A��D`! XEF�� !o@!�A��T`!@F��`!DF�A
`!@��@`!H+!!EGZ�hA�� !ARQ��@`!@FQ��@j�B�HE�� !DFT�� `!A�n���@����
*��"�	 B��/������=�O���?׿����������y?�t�d���{���7� "
�����?j���}`� ����?�>��S�E��@�?z�@D�������A����?G����{�+������I_�B��E$Q$P�ET$QdX@D	X��D�E�E�@RAEFEFDE�aXE�Q�a�Yb@X@V Yaaa`�@!�X$`@Xa`1E�E��E�aa X� !dQ�#a Y`�@!`�X�`EdE��001(AY`@Yb@X�c`�X�X�F �V,�@X�X���A�@X�DX�V,��X�F`�"0�DX$Q�`�
�F0$�`F#`�X��XE�@X0V,E�E�`�@X�FV$�bE� � "@X�@X$E��F�F0 ��A� ��VA��E�Q�E�V��@Yb�d�EYaad��� �@XDEX�dAaEAA�Q Q@ 	ET�DD��
 TQQ�_�(�?���?R��(� "(H �2
���ϰ�����}�@���`������AWA�P~_�����Չ�;O�� �����6}�Ђ ���!������ADAW�@D������
 �����*"
����%���y����!_���:9��6 �*ϲ��G� �*��H�w��?�~�C���D�O�?�x4��*����D_�\���H����%������~?ۀ��:��<�� �*�."y��% ~��>� h?����3��A�����Z����>��/����1AY&SY������ـ`P��3'� bB��7�%"*�)�ʶʅ%[aI"6Ŷ
RUI!Q%��P�3aMR���(����
$AIUZ�(�Q��(�l�3j���V�UBB)6P*�R��*��U�ZbE R��UJ�**S��Q�F��«�����ZkU$�LRP(�t�EE�F�JW�$�B��)�J6Ȫ��@���EEET���-)��1T�BUu�%-�$%�*)P^  a}ڦ�,}k�����V�6l���lim-(�me����-)
�F�V�f�d��TS[Ҷ��,�֙j��UZ��i(ڒ�:`*���(�5�H<  =�z6�
(��r��=>�P�B�
K�9����5�J���6�5}7l��C� -�*�m�T6�([*�e���j�0Cj��jT5-����mt��	���/��R�H�  �����ԭ�D��IaUQRҁ�����:PB��U�4Q(]8S��l�j�-�`�Q��$(���P�DJ�>  ���*l$¨�Um�+mQ0�M�kV��VQ&��j�mT�ګHUBբ�"V��)"�e,�(�m�"�ڊUR��������  ��Q�Mm�T%��R*�ƛIB*�����j����(���� �X�Y���mjTCU���J��%EH��";eR�R�   g��(U�f��ҡ��m���p@:0 4�e 4�04 �F 4 �j�  ���kT 0ԢUUO��TrPi��   -� [��@ 1� 5Y�@3S   ���4 f���FB���CBʖ Y � 1	(HQ)T��     tl�@ 
�U�Z 4������  ,L��Q��j�a�P �0��ڕ#��QV�iH�D�G�  � ( ��� 5�` �!@ �j���� �54�� ҄��[  �0 �)Xɀ e+�_f��*�%A(*T�  >hhe0 �Sj  fT�h �F � � �0( �XP�(*5�  ��@ h�O R�@  E=�	))SC@ CM4R���HO��* �Oj4T� 	2�eT� �jy��5���j��_9~��tm���$���urdT�;=�tBޞUġ���>�z#��z=��ϛ��������?�`���1�1��]�lcl���c�����ת���e/l4	�Yx�C��v�y�3F��0�b�n�U	N���R��Ү��G�?�F*��Tڌ�dG�3Z�n�
,7��+q���� �eBmhÎ��6�I@��Xe��Sv���gm�tDT����d���r|D���H.�ә�XC�^\h`a�1�ƪ�`�4��8���K)	Y�&�*I`��Z̺b�=�k@���NQ��kX�%�32"����F���j�skٴ1d�o[')I
�c�T����6��Z�n}v�!��Cƈ'wm��֬�p<Ԏ�-hʉNm����Z#T��B�:��I�wc41%+l)�6����W�`J�he�Ai[�L��N^�D+��;�ӡ���y�p��[JPK���v��������3oMJ�\I����ZU�����ol�A�wC[7"�jd�J`kC��EY������bp�5V=��r��2[� �`i1(�ؽ,Ri���[o~n7�X�f�Ks4�Ov�[�I��X�(�Ul�2އ0�],�Q�x��b��L�$*0�0���1�������lMܷ�fDԭ�Y8��p	,��ãjD۫9@vo�h�P��7"�"�n�j�Vbˤ�y�q6$���A�Nb����v�JHJcդ#��UmJy�������WY��A2�X@<X$A{���WX���Zn�S6�f���DĪ�n�䘨ɓX4�QV`���H#��v1��-VA�-�CPi�r�Hi�Z�SQ̭�+^�R� �.[f^ʀ+�n #�zNl�6�Shk�;�mkHU�R5�w���ѕ�M��Xb�J���k\l�G���4n��IhA��a�� �����U�f�o'4@��YKFV�S��@����ui'p�&n� �����KE];�ۙ�cA�ښ/�b��O0�C*(�U7\�Bl�Uw�4iÄT�n�R�u���^�m�s3�>���xmGX�7:�-G^�tSz��"*4�Fh'q�Ud��juq[�R�Z���SPh�jհ��Z�-�:m<-eL;� -��\��N��UnXaV���.KGJn��7b�ي\u5֬��b���7��%�u�y�ZՒ���{�8�SA%���M���޻�gUj4/i!N��Q�r���N���`�ݔ����n��7c�r1[�`,R��l��1*r�	�̬�ISx�(�e(���v��u� ��؏6�����2��(NX�֫t��Κ�h�*[��6e�F�V!X�^=b�3ȜW�Rly�s`*�֣;ZJ��9- �ƍ�[N���Զ����k4�ю�����R����<���а0�ym��Dv���ɸ�x ��l�&�)�u]��~L�:΢�.6�|�2�.���[�q�H�`�ӳC*Nc�$���4�D�m��f$�;Y��MҴ�J�yVb�r��YH3-˫s3%���ʰ�\�V�b,��q��C& 35��M��\�� �Z��eԇ�X�z�[=��jH�j�`�����i�� �?;YKD����)�ڑm��x��-w�oj
��쫵h2�Ř\�{�[��F4�ݒ��5�j�ʳ+EʘLc���ض�\�nh�!E�Sk[�r������z�@fV�Ьl᥺B���jhw�m�T�jl*�6e&�YI�6qF3
DȬ� �gb��r�lf��Ҩ6i�q����G^VvQא�s"���R5y����N�n����m#����[�qǬL�R���N�R4�Ka�CC :WB𩂫S�
�Ϋ'u<���u9��MF�0�snک��ea:iL2[K^����N)�^�$��&5!kVEV�J�^�s���n�8_j����fZ��ѻ��[)drY�xF��^ ���!�>��T�Y��u`*�)��X��X6^#����9�6	Kn���͚Bf* �ɒS���1m��0��dR�v�a�	;b���g
�.76-j�V�7wgH�o��eú�t,VTB��N���D.𛲆ŗARPᩗHk�z�^�yA<�@3KM*ς�#b��4�d�4����]-.ӛ�{x-b�)ӡGRa� Fm¯nm�E�n��N�$��cvEw�i������/y����������s x����ɫ�X�Y���.�H�D`�;�C�.���"1�̛���*�̒H^q�e�C��#fa�ٙ��ǖ��ɥc�m����`I ����V�/j�j�o^��P����&#"�7EfS���ַ`7�N�� �6@|~��c����O�;�1�DY[M	�u2�ʼ�ͧz������$�WOv�ROpY��R��<��(���%m�듒u����Z�5���Ȍ�k�ح	@��^6=��u��h0~͆�вAGE��@��33{A-������rPN��E�9�VK�Ua�2U��gUԩ��b�NG�R�lm�)َ}�0�ُ,��B�,��T[M�� �i����"�*��[t��kU�Z%�6[N�T;ٖ�V�j�|]�62�(d֓���mTa�ڵ�M7��n�X�)�����y���6͢�i	i�A�B�7�Q.�ԩ��G�&�W�-@"*5[1<7���f�z�
�e3��I;f�;A����J��v"T.��`,ě�͸-�et���a��o��l2�㚩��ה��C+J�)�:WX��~���`n�AM]��&�����Y��4�t^��D��<�m�!z�-�����U5ouxa�ҧ�bJ��Zj�ő^�j0�V�e�/^ޜj�XeB����°+�&�s&eI�E�9�,���;�p F
&Õq�q\EB�#{�vaК�5̗��;-͠��e�FPՉS���Rd�-M�عr]�@!�.+��̆l���Ool��7�XN�@%z.��a밮��U!Q�e�-ũҼ�LYGkY���k,�x�䀁y��t^�PH��^6�%h�~ҕ�^�ܔ�!�'V��d.���;.V�jMub�*V˫lc�6Ӳ4�4�&05o��>�n�K"Fcoqb�?^ۉ�wI튵G��e��ٳ���zY
.ƍ�d$�D�ebj�K�8k%�4���m-��P �����"N4�M�@�����+v$�]c�q�HM	j�e����#�[�J��.٢v�y�,�#YPa��d�>�R%yh�X�.r״�N�����-� �ߖ�{J� T�w�Zs"l�q��v�+�ܷ���*+��oAr�&���x�jI�y6��x�ej-RÛ(�;�4�7�*��p̹��{v��r�J�&�#�&B�jB�w���WJŪX��h��ۇu:?<��˺��m�r�ݫ�KR�Yld:I�5�z����U��f��,c-�dAj�EBRC.���&�M5��y��v�Z.@�\M3w�J���]h�4eYҊ���M�ꎜ5�ڻn ӈD�dc/t�߱K����w�����c,'w��b��"h�-&�Z�6�K��M����fu\�r�n:��$7Y�s)�D+R�Լɖ�9E�Oh#'}~w����PT��*
4j�Yr�#yiM]�ыZO��N-8M�s��{6��)|)�Z`��,@h����'�2P����ۥ�i-ll�d�5+X� ��A���;L�f�p<�4�m�IJ9��h�M麔�34p�
�J�]Jl���eыmfD,��+��:���5����j���hn�y����>H�-j5!Hia8uh�h��rY7Zڵ��1���Օ*���1i�&��*�V���z�%?#e먲58ҕ��%��j��p� rm�V�M,{�\sCZ=L�o�̡d^���6C\a[�YO(�ٴ�^�Al�n'@nh�M)���`�lW�M�lM1�C�e��r�K5�!������f����xk�#����*F+^a\N��h={�-]] "�m�C��a5�Ҽ�=��&�9�YIGB�`P�ݓ���QC!KJ^L�U0l{����`�H5 D�įj�K���8��F��&T�Ď���j��m�k1
�2ab�^��ŭ�6%�%b�0��E�X��L��T��J�E��a��v҇:�<
�U��n5�Ԯ���:[ِ:�L�a��lGR�
�$ܤ]����Z+e���v%��X���>N���$6L�Ҧ�V���WyyD����R�^Yk�ۼ;��e�Z4��le��@�A�Ǜ��J��:��Ѥ�gd�7�!���r̽��Ք��Ҋ�
�rm�̑@!�Ȫ�dfOA�.���ݨ��X� t�"MSn��u��q�޵G� �7�ޯ���6daӵ���b	f�)i�UNԿ��;��T��,�x�����t�����6���Ą��w-/��h�Xrͷ/t�GEǭ˻nL����NL��;�*4��q�hKY��U�UZ�[�0��6[�z 5���Cn&�J^��*��Xf9��<�+R��b�����|EJnXgD��@���#a�{%ۗtU����a���іr��X�P��km�r�5G�(F�n#-�����;jF�e8X�$tQ#&"�c%�.���l�%Rwܻ4�vСS�Jԑ^݃u�nk�]�W��j���N�*9Cjq���%.�e EJ�mʼ-�em��dE-�Ga(�wMT�V�[�	�il��B6,�[� �wufP�!��Pʹt���V�b�/�P3(=�e���R�nfZ�U9�˴˹.d
��ȒSj���8�Rf�h���t��p����R��U�-��!rjБ:�b/I#]��,ڍ�K�Z↵E&�WF���3����)	.�V:ӕ�A@d����v�� �T����u��އ�5YN۫TY*T��[V
�U�Yym]����jB���CV�U��FV���dQ]h����.ɖ�5�(d��/2�X�]��:�,Wؖ~���&�.� �)VQߥ�ɑ]�U72 �IX�A�p��W���M�����ŏm�����X[AL�ޢNSl]�3hm&cCb.�H4:�oXT�ShS5،��^��� �p�y�"(:i;!
�3l۽�j��+Af�T�C����6��ӦU4�C���0e�u�a�v[�QS0�RJ��	(	� I-���,5�SY��n^
й-fmX�;��ܨp't++O4 R*,۩e^<��B��tDm%�@���dSыM
m�I֘(8f���_��l7�����j�Uɶ[�����5j�٣6}z�mCx��6ڌ%@:p�س`0b�� ��8$cǹ)3���vAF�s�^$��Xs	Uu�j`V��Z����e��&֥�U��B�iC-��Mon�[w1�9��a� ׆��Ց�Wr�i5��%�Q�_5GC�!Զ��"��I��Vk��� ո~ NIwVJ�i�/vY0غ�n����v���io.�oD�������`��t�E�VC�Q;���T���86�H�4&Ue�@�f��[Z�SIX�U�eՃ��i�"j����1�[{s~8�B��5��S�ܐ��r���M�̴qX�wCƗ�K�Te-��1Y�,T�tDi
�N��h��n֓rҙ{��Ǵ���!�l��X���7Aԫ�so\T���5�2�+���T��m�h|�y���]��ӊUl��¾��Ҍ���b�l�/]�	@Z>	��r�$�4�D��gt\҆ա�.3��44]��y��Y�e�w盋i�����,��fR��+J�3W��l���g&�n�H��qb�h���h��V��Q�0W:'�S��g�%ݲ�i#��WVa��U��yt�����T�i2�I�6��;"v�R�'�2�g/v��Ta�3ki^d����\Kw��V^��U=V�v0��a^�/i�R�]�vó��0,��C�l��ǴCY�:b�VR�Ő��В�`�kc{���2_ن�ܸ�6�`_5����j.�	�Ƣ�4��ʲӥ.Puf���W��d�ǽ��[��7�/�S �n�RlÆ��>o(k4��H����N��g(��yZ��f&�J	xI׬,W�VD`M=�/$j=�7&�U�;���{��*���¡a�l���5�jEn�٨L_L�Q��b"�ɶ��^*e͑5�����%"*�Xd�\���G�2��4��n\�����^�VS�u�UL�Eڷn<��Q2���[�[݄�l�vB���)����IQ8�lw��p�C���V�r����u^�f�US�e��ԣ�. �U�In��L"�;z�)�:�WV���QHRǎ�����^9d���
����wz�ñ��1^tݶS9��Qhm�`��o6�˸�TXr�6�1��)�#��O��-�&��ZD�6�Z9��	"�Yh�3S�]룫uh,8��M�ZK"�b�WR�R3����*]�1e^�X�o��SF��������D�.�0�PTOA�#%�j (Gނ��(kypJ���̹m����]�u6m^�-E�4[�]=��8�n�֡���PI^Z
Hn���嶞���N�n4�ۘ���+H�mV��Հ;�켱[�R�4
*��r��(\)��٦��0���b��T�6��<f��r	vج����[zhEwjȵ����l���g%��T��2m�KJ�0aW6�8�Z�kʍǸ�w=�7p�fT�>�bx���3��j䔡eX�n�.�w5��LF�c����v���Wl�R*z�Gm��OOn��t��0�2u3{�LfI �˘�S�;%֖F�`�^�/v��I̩�6M�&q:mm��0%�٭X�دRM��Zȕ>ɶ��Z�
Ȣ�NĊe`�kg)�3�k��;L�-LG��-TKW1�w/���X:s�0��omf<#�+���s��cY5��l�ϭ� R�sVs2">�Fu>�{�P@ţo��v]b�0D���#�+|��Hum�iglEI5<�m�v-jT�>9�3B|���u�9<t�] ieuZ������qX��xr��ݣ�V�ߓ;6�����`�G5zHNˆ�Qy+^�W��k5E�Y��dO�:N݆���Z�TF�nXX��)VԔ#�G^�H
X�-����44��ĞJ�p�4ӕ�VHDZ �_b�Kz�Nٚ�=�!V)�eEg�>�W�i���ՓUvq_n�V��+��'��e��ww�������C3:���N�<{˻��h5��k�f��h����6�^.[�z>sn�Me_lT6�P;V]��-�e�ugn�5cf9�@�8b��V�Ѝ�T��.�ys���[b�L��۽η�I/�ڡ"Ne�\h6f
M	΍��C�(R���αSv�01���{�[�l�t��͋cOx�eW&�*��1�N!���'���j��b�,��U�w@P�E�̀t���#��stȡ��+�=��@v�V�3Px�)��c�n�ou
j���[��(CM��' B������ͼp�5���l�Ⱥ��\��0n����V����x�0����N��\�O6�wr7OQk^��ˑg_���\�ki,�W;�[Jõ9�9l7u��!7*�і�Q����P�]�]=&�pnԥ sVp�G������gH��@�3Vk��yQ h��uB�\����L岻�KQӀ X�T.��ap4�Ci�ޖnƯ��s9W����Y�.ѕ��u1��(]�y�_ʹ����]$�K���@�Y8:�>����;��:�,��l��e��쬽����t�Nvn9y*RS�� ��٢l!�2�.��[����](���}�xq*h=�z�@��mm
��7����6��D������@NP�|�u���)2�������Kp1�ΠӃ�:ԅ�A�nE���9��;�V%Yz�[\j	
v�vK�5N �I�Dn� ��NJt�N�k��`���u�ƓՖ�ìQ�T�ֶ�60.[�u��<Ճ3H���\�I��C�!K�kÙ���)�Z���v֪N��[[��A� �n.N�]�i2�Am�vn�jAC�镆p�������wKqҵ1,HCB�$�gSȪ�є�f�Aw���WW�E��}f�a9�uS-1SnB���M�w����x<�JN�%]��ot�WI�Ԇ�.d�)R�Ӽa���wt2�s�`br��HbO-�������2��[/y�+@9�>��eZ%�3��Jv�^�[
Y~�@���)c�,�m�w�;�ú����2�B`��!�Vi���uV�k�.�z�#�%�j\Ӻ;ql=Q���n(�1�gX�Wʾ�����GW�k����9��r|wu�OS-�*���ASo�������g5g&R5��	
���Gzi��b��{�VFێ�칕��[;��^�ʍ<'{��չ�c�k�C�r9v�|���sI��F�@�Q�Ղ��gv]�p�ĭ��K�_b�)��@ f͝:�kK/-0C�t�0*��y�<�N���gX��u�Ya�t�����aj�`_e9D��?�ZZJ�s���2f��\��s�S�X���L�{����r����:�e*k���^8�r��ؠFg�Q	�_ʴT%F�}����]`�H�S@��;,��$��#.^E϶�r���ŽZD�':KͦD�"*G���1��ecX�
�}x:�eL�z�_׭5AWRu�+z�]��;������O�=;���"�a�T��Y�А�5�����i�}�2Pp��Ս����quku�[κ[Wl�qp�ϯg*u4j����pfdT�\����Qק2�s��[��`�y�NR�ք�˓D�!��P��.��e����F�m��e�h)���� f>k��$=Y�ޤ6���[������E���E:#�d��b����m�&i�w@X��-�n��:����e�q��0=|�Y�޾��HW	���e��1��{S=yڈ������*S��S�X:����n+R�����X��\�ھ��x^�s�]��e��vġ�IoHgl���I6�u*�� �dαP�QOV�X{R�KXפֿ(��Th�a;$�����J�S�!J\��K�f^-]o�$�7խ.7g/d��#U�&re+��� ���g>�)��2�����%�r�Sąˎu���X�@a˥����z�과�-ߊ����s����w�����q��C����}�����#I*u��<��R�wyn�얪CƺQזz���Q��=��xX�U���7S�b���}���x�	m�A
 e�9��\�FlC��v�<a��[̫p<y\&�q�X1�fk*Ro-���Y�aY|�<haq���}`k`mj�G�N4��ǔ�8r�XU�K���h���U��n����=N���B���!Yl��0�������ڒ�%�����-b�����C;���/��p�ǖ'T���Q�ʹ�u�P^H�^�W�u�K�h}fS�r�&�RvEe���#>Pn����[*�Ԇ��<�+]"1:�����v"m[R�j�:����iS�|��+v��ʈC)@t��&s�t\��p�ɩ�P��98^��%M5�y�hob�xa|J̏\����.$q=ݾhn��/�.��9J�	�'R��yCnŭ�neD�3���[��w4mWv�7����N6�ӏݪ��f��p�u��֡$Swh�\�m�����.�}�Bmow|-l�K��\t��[���~.P���ڞ�ɸ��&��E�x���86�[[�L�#����mc3\#�ʚ(]�u�x�>�޴�}�u��KӜo!��`��J�c�:��V*.��݌wGe��lX=�è�W7x�p$;O G��1k��{�{�s�0�8�ۣ�)����*�r�0#��fM��L��^i���'�Xw7�I��)�ߘ���e[��]G8�F���:����K|��oG�-�z�5��p�Y�f9Ǌj�l����lh�� ��!�*�mѭ:��=
ͣ�L/p�72�cy�� G-m�㾟)C�l�A\��;YN��V��e����sm����!2���	JpZ�u�w�gM����u�� d�ʬh'�9kn��$-=�����Ժ�lt���u�����T޴Y��\��OX�=�{��p���Yb�V%5�cɊb�[-��	A�n�Z�d� h�U����/;cQ������Ɉ&Rv[5Nds���c_�J�@]e*���ʘ�,��H�u��i�n�s�y���:����A��Et��:�9t�pYljn�p�I�F��RL�nwȧy�����xտQtÃ����l]�˿�e��)��>���"*M��X�ٚ� #��[x�r��6@Z��2��LK����!�.%���:ޔy��+��]b����%7��+��m+�ʲ�O������1h:���ۓ���1��R����z��
�ҵ�jE�o8�5�.��mѣ����������,U�������E�TY(u']�x���h鵫*0)��K+z[�l.}Ƌ�^�S������{��f��{Ԕ��wK��2�T���$ �u���JsoT"l�j貒=g�Wr[�Z˾�n�#tc��ľ�|;kl��ݢ�s�}r=G�Q��}�]#t��u�ec�S��2���me@��5��X���{v��ض� =�u��"S:�sN��s�����%]�AP���5o�R�ֈ��O\m��4n*��w
ݲzY7�����o%ܗoSٝ����YLS�v�m���T����<ݗ�g*�i�M.�#9����<7ޚ�{U��v�:�����O*̵�`w!�DK]b?��<6�j��T��,��1��N�-�� �ќ��ͳ[�h-|��yPA��*���v��Ψ;�:g-��1�A�bGw2^�q��\��z��+����N5��e�J9���֮���-o8��O���tNK弤 q���&%�m��)̫z��
7���^�^}�J�=�2ܝ9𻭒�B����JCH�
�w�ӵ�]�_*w��G��9�R�eJ�y�`A�[@��2*����;C�u�Sk���n����s|WM�m��Ѷͫ��Z�N!LɖY�5{YAIq���$��Q:�;V@1Ǹ�<Ŧ0f��Η�8j]dھ'zb�wF�
���T{ B���⛄]qVY
�N��K7,\ֽ�4/n&;GQ��Xv��ժ� �5ȷ�򺘬��*m�R����-�뗥qu3ݶI|{�\]�1���������'%Y�'�-��s�j���Y�$R�Ө酣Mv����:��_V�|�^�t��+���չ8Wq�5}�.[9�;v>g�����L�pN
ˀ�e����;4�x^�ͫ9l,%�Sp���jd�QO�*�DK�zry\�:DJ�Ǧ�]a.ȓ&�e=v�����f��>�1i��_k�4�5�Emw��L>^�s'�hآƩ;)h໏ܫzIgX�;;���댷3��7b������.C'_p(�ӥ��AK��5X^.�����9f s.�u� ̎R9u�i�9rZ���7�D,�ń	D;a�+`QZw�B��ۖ�J�KK-q�Dl��b��쾃m��p ��9��]����}�=I].�#�)FM9$����<�G��s4��
�qWSDB^Gk�E���� +)�E��tqe�єu��tpmo�X�ܚx�����p�wgD�hQq������X-N=�h
va��N����D��K�}��B�V2�}��k��VV��J�|׶/m!Ӎ#�A:���M�1P��v��DE�퓩"foX�@�Q=������mTMhKT�AW����1�Ϝ�ڶS��Vj����Y�AԄàՋ�+4�zrA�����Z)Q�Q7)��(e:-��79^�o�h�ʇue�yc;��Z�Zy*����Θհ��	b9�!�9�q���<��(�v�ǔ����8_e��{�`�Y:�7{��r�(��B�5�#�Ӆk��4�I��W؋<�#�ҳ����e�7#[��L�)жC�P�\F�fBsoS�i�*�cU�e˽bI{��y� U�a�i��+Euhm����C�%������ޤ�V�]����>�y� 5n����}����;�+��Q|�΅=����Ѹ�A�7΅����p�1�e
�;kB��2��﷋�yA��`f<������MKQ���x�v�� ۩nQ��h�]&��V��,�%���6œ���%`��T�ύ&���mɖM��%��I�}Ȁ�vVw'��8/�R�V��Uu����E6F!��|c륗��˹��kc{Z��V�I
V�Q�����Н[��Z݊�Ԉ�a�,̤l����6y�z�-�����tcTٺ93z�ƚ�Z�"5�.hm`̛|�K[V�8vh�{u�X��t�{Y��+;(wRc�gӰN��.�J�K%�:�}�.��l�vb@jShQ��wI��Ծ�V�j�KoY�ؑ�UzHc���t�qi�� �ݠ.�W%XZ:�4ܫt�㮷l:�^4+S6"2���O��s7o��j����L$�	K��֦�pp���о��Ym^mc�E%�r`�=BMZ��ٶJg��Tw1�>��ﮑx�/�݄b�ؙ�F�#�g=�4$����R��ۜ��t�^e�j��ZI��{s�o*�f˭�瀠����]*9�r���P�{e	ȃ,�5co-��]sP�S���2��d��|b8���X��Z�`9��CqL��]����}4���O���|���
�.1Kg���:^�Ů�ιO��U�L�6�6.襅l4�B���a��@\nm˳�]§u݈в���PF��}N.�K.�%i���ۦ�����ro3P��T8���FE���C��)d�z�m!{I)8���Y]�>��;vA�B�m�B��hwX�	�t&�Vn�jG�3U�y�y8���爪=��G�_i�ԫ��mlu��Na����^�4�^��T5�)R
����Yu��Z�WIJ}R�77w���41��ᑮrY�� }�.�2�����T)���;��(2>r�eem�&��].�ٗƔ�4TY� �_#*�S������Һ������GҢ�{����$�)oJ �2۾���]w����1�gN�4����W�ı�R�x��m�*p�gA&GKo\�w&*��Ы�9��:��5������+�
��fe�j�R���M�����n��X�9�J��G�;!N y��ֳ4�*�wD��Һ
�x�4c�%��a��.R|�L��f�<�.�4��Of�^-����lu&!�&��+��2�����l�"iNZ�wV�&n����#Ğ��buy�� �	�<��1 �;�圑�euv���Q�cQN�3�vfQK�YV!�,���,��!��W�dW�[�ݷL큛���v�_Cέ���J�+:f�Yo���뱥j(b�v���A;�����YE�t���xm��w�ul�����S���5��kgVh��R�5#�l�(����r�]wz�G��ѥ��[D���_e���NvD/���Z'v1/8Qa��Q� !��T�e$t�b�"8�o�� ���|�'8�Y�Z1lǴ�����q�ƫ���눑�@�I0:���WV�ͬJS��nֶs�8�S��*i�egT��������ͣ�K��G\Ř���Yn�ݺ�;���&����5�5ٱ���dw�"��Y���KR�E̡V��r�fQs��d9�v�t����t��9U�;��Y'ju�(ɕ��D�jg^�;wi��*�oJ����]'cW��:�:��>r�w+�)t�I|&<��|���]���?���wz��������ê?��~=�s�ޠ/�n�9̭ͨ�4s��u�E}� j�8����>�����"�Б�ڍ'��I��2�&oY���z /����p�f�#/��2��um����`����h�ˁ��-P��/���+�U���4戲頰�vC�YJȔ{r֡�喂x�h7�{i��4�[p<���Z�.�ӿ[�7A�Y@N�֪�l��I���t���[Z��Mq�m�==���az9Q��m�T��t��:n����*�醳�>L�o�V��εIsi�sFəm�����+i��rA+9WS̏��|�(�V�u\����(>�9��]&#�̔x�Y][t��TV	������Xͺk�x��b:�Sq�v��gRݐo�j��2�<z%�g���]Е�+�r=�����l�v�c9E�s�����C�,/E��ˡ�.�P�[c�⮫�f��w b��oU�ۑ���x�Ed��Nc�P%	�\h^�C�JV3ށ���Ǖ��\Ȼ�]j��	|�WnC�G��r��u���k�7��D���C��5ր�׌�r [7)�k�z��0bz��`�yl4�v�ب������uh�
��Egsa��8	��ˮt��Liu����&���c+z��t�˂��|���-67{�5Ùݖni��*�YboQ�{��.�^u$7;\pR�`f�oF���%u��ܔ�}�^�q�g&:�AJ�gQî3\I:rk����*�](��1Gk�ejΞ��ZO@@�F�=R�ɢ:�4e]�LmK����P��Z6�p�׉�fM��J*��:V!W��No=P�~¥J9�����\�� BB��W$GNrWa/Q��e�t�h��N�k�y����;�*۠���v��I���)�5�ю/t!+-��znm;�2jg6�_{{�����@��N]J�44pe����<��B�����N���V*�-�|��*$��ܮ�(��g�i��{��{�v��9OvU�:LO>��<ź���wIRN��|��gP�#�Bo7��.2�iZ��N�Rn��-s���������o~�.ʴ�R��B�a�ć-�L!�I���M7]���iU����z&��ƚ[@��wLt��h���V��WL�-�=��q�k��S�{���n���͠��������o7��V�=gP8w�á,��H���Q���Oe�&�̹C���=��|۷l���]����CY�h��i����+vb��A{�9I+�6�_!b�:��X��.����Ӹ%e���:I޼d��*&��E��qlS�coh���$:|��ϡ�
:ݡXqA�"��7,m�ȩ*�,z���Ӻb������+VDɸ����i��F�?=`�}ʠ���rΉ�5��>㪨�
Ψ삯��rb�c7b��k��V���4��.8+hWT���'�0��7�˦o����@�\�p�՜{(�,N!�)Q��k�����wZ�b���MkfL�-���{����J�Ne��u�*KY���;�$޺����S�f6�\m�b;=kV�b3*v�9G��C��is�W����U�Z#���G1��X�m&+Q��5C��C�ʹף9�;r�Sg�:�ifdokz�����%}�#��0��vK�Rr�o%n�f�M�:��vRՒJ)2�k�$u�F��ԃ+uI�7k��
�n�f+C��6��"�����J�QB�kF�TܸR���E�<�Ϲf�Ղ���rr�(�v�
{�M�%����s���=����a�e���̼C����u�	�"��pw�����n��n�yҋS�Pxi�ѓc���}O�ȃ�2g�$�}�:5Y��pVj�Vb)�uhcn˵Ke�l.s)h����u�ZY�*�O���wZ�6W	XlG��!�����t�ÿ�Q�������N��
���G�s��6��5pS�"�^خ�x9%
]ɢ��xf��R�U��È3]�Y]ܤ|t���������㷣Us4��uPTw�G��D�c	 �Lɻڕ��a�֡H� �G�@�Ѻ���j�XY
U[)�M!ٔ�����T.���u;L�gWot��l��ݽ_iQv�TS���2�*�h�>�&��O>{��NL��V�ꑻ��xr�5�b�[f򮓛P��rul��n\OL�
؂o�dV!�6Mj�|�gf��7��1�8�=�,�cb�Be�l@�^S��z.���.�»��UZ�2��ٹ�h����j�U�d��ζ	�)��o^���Pf�'�n��F�4ѱ�0�fi�TFH��NI�,e	+��E���bB+
���'�GM�.��D�[��]�$���I�3]�3\qN���gQ��Y1�F�6ȹ����I�-4-�i�6Xԅ��]R�v\�X��b���i��Z�!S�ӫ$���fYг��w.Kj����q�U��:�n�.qepЯ�=��&i+2*8ᰂ�Ùw�aG��ҧ2j�r{�[Y�M���α�Ws��״��F�e+��'�Qҕ�T���W�Y]�Mc|FT��-��B�:��Ʒ��ڨ�{�=����Nģt�d�s�SR�ZkfJ���:��(�F�r���$�ۦ�&���ye�g�L���w������-�֨��9�߷C�9Ln�XF�r��)�ޤ[�,STW9�]ԭ�����M#�f���n�+7��{Z���{X��͙�˭��h�M���$�m��y��%��9�]���)�;��N�n%j�tg��!�v�w�t��4�8�>�K��kԶԋ焳�C�]�gq���Y���ۣ���]b��[��W.��w ��Mk.1������/�^f!,*�z� �'G�ʖ����)'W��:xz�T��CѽC�0�j�J�Bާ��-Ძu�]u�� ��SwϮ�\u���T7��C����������ea��uڋ�7�&���u��@�Z��dێ;3w�+M��p�Ql����]�,Xc���WGX�r��͉�y�/9J��WW5��8�Uz79��)5u��L�%�7�;����޾��E*���J]Z��g�ËV��!���;y���5�u����1+{���;%�F�
�-��^�g���oR�����oB=��	�`G��ŚŨ,����9�hӘziZ�6�����X,�۫ˊ�	u̬f�\� t?;xL�wI0�b��ݬ�%8 O79uh�]J�#J;��niۨ�u�>?%J��˳c6س��Rmu[�d��ۏ��]��I�F#z{8S�݋�[��htV73M ��$�&�ٜ�n��`���E�bV�cPnS�sM��$���K����Gu,�;����|�f@���[5r���\���M�W�!�l�|�]��4�Ms1��)34�w�V��e�>��3ri8�����d�ږ�c����t"5���͍�L3��X��U�3f5҉y2:`^w$�T�[��%[jNR�Q�|���y��h��c�+���Cà8��2�f�D�:�v�_>���r�����������Z��udԠ^�����;��f_q�\w��{�}4M�����ä�OF�>�c�}���=\g�Oe�U��X���7>�{w�*�t�.�/u������O
����ޠ"􃅆��-9�Ǝ��j�gJ���W���Y���5�"W`��}S����ww������r^4lR�,�W �n�Yyp��'r5��X�Ю(�g�*�S)M<OƝ!�%�o3B�s;7��| Lmv��.�r��r(s^�ٔ�Z���i��/@
L�K6"3F�2�Ɗ����E[::��X��������Д���]����۲L41��%f��u�WoW�9�QC.Y��;3��Yb�8�]���%��<�R� �v�I|�k�}}n���VG{�>Ǻ��vYޢ���i��5�����N�5)'��I%��ea��u�ٮtg-3N�'wL�ܕe�e���N<:+� �z��iI��G
�-�t]e�Qd[P��RR�n-����-��9WM������!�]�n��Xf��Y�$����sN�T-��6B�ܳݏ-d,����x��*�{�U�׵O�s���n�޷n�X�0��>�eЩ.eb��l%��b�c������7������kj��|��Ø�!�)LO��|�8{csg+��Uj��T\V�Wo%�Xb|v�ײ�6��)f�GT�v�ۛYE�]�g%���ڒu"c��LH��^�h�A�P:H�jQ������r�Ԅ����V�i4�ژ��Md���mN�a=t�p������ֽ�h���}��*N�O~ӻۢ��A�n�{ة�%�0fM"�P�JmL�,��J�4\�N�F=
v�Q�.�=ֶ��-V$̨V'�C���'g<r�>���-�d'��v�8�m'w�溂՞����өD��;+3�7�� tbLSPJ��7��0+�B��I1��ӓ��SH�F]�,,�n� ��o���{R[��SXz����f�+E�����:���{-��VR.;[���wBQ ݔ�+2��m��kt�Q��D4�9h�Wǋ��G��5;'w5{��N������A�WŨ^�J���ES&Jƞ"����i+)��t.P�p�L�=ᩲ�M�
����m��t����`����TLvΫj��1����f��WGob.[\�KS86�m�y�P栽�8���s�$�|p+��c��G1�����Z�j¦!�8���zK���[�s(%������;d�V�
篂:ހ[����:!X������д1��eA��`�׺v������(q���p
5+a�s{��^K�]a���Q�7��*J�ζE�;hS��b.<�[�jY3(ҷ��ytλ�F�}]٢�����V�N�x;��q��/����׼؉��'���%�)��9m	�9��ƶ�Q��v�K�}<W.�d#�[��/�ukR�2�)�5��.d�D*B��R6dǛ���Vu^�أ:m<F%e<�r�U��38�;\��Ř���+Cl��%6ib�oQ�+]i��ب��3�X�9`�%���}O�����+�}��b�Vܰ���{Bݝ�Ѹ1V��j)�0JWcsQw�C��2��gߙݓE-�,�:2G#��؍e������i h���ZţKG^#+<�ס�lAH��z�Y-�݁���></ࣈ�57u鰛�'��q�yvV�i���.��i����yof��;eN����N�藃t�T��F6�ײ92�ً���x���
.>}��r�%��<��3e,`jͲs��`X�y��3�oS��4WA>JboL{���VBFF��3GR���f�s�+U(���b��A�7�d���2��;�q�9�|/vJ�X��Û�ӂug[Ǹ�%���Q���Z
w��ހg�D/eE�u�Ő���I���4�^�3�:���N%9��l�M�Ք���gJ��+�m���!H�j�G>ܵ`��r&v��\�2��z�v�dX���֠��Vq��Bɗ�:���D���^���,��-��H�h�}�̾ ��`[c�o�E��[d��3���|�I��|5��ZP���ͽ@�%X)n��|�+��;��ݾ��t�F�5'�r�+t��<��<���o��:�ѱ��^Ͱ03�A�kï%r8��4l�0ɼy���-������T|p'����Y}��}osi[犱Y�ڜJ�m�q"6��M��uLv��Ԭ�'�m���_	�����0�[kO�K ڏ����+��ڨv�Ç�l�B�Y9*
nVH��Jʾ��p��f�W����K���s�f=�X�5���ݹ���|�*��\PP�亙���ɼd�6nW,�2p2�bCX����Cy��Y]�Ygw��~��f�E�תe�����T�H��.^Y�N:	�l�{B���pc�̺���h��B��҆ �@T�gh�-j7IV�Ph�Kiv	֐��5��:��B�\M��m���.��_ۈj;��,|bTv�.+��mx�u3��Owu�Mp,Ƌ�+6�Ćd��zoj	&�v�Ě�ܙi��HG�N��E�$��k&]:���%6�li��5�U[� yR�kv3k
�E��`��{'u<=KnY��[��w�p����g�����_wY��k��uv8��3t�.W2��s�j�n���(K�r�d�eEm�5��r���Ǫ�|���HkJE��_vIN��̛�'GL�.��Ủ����i�5&3W�V�m�J��[ݮ��h��1Eck�u���`�J�*V�S�sA��t�s�y�tP�p�����޹��-��o�W[WH�r��b����tns�΢1O\±Vi}]�	MI� �;r:�P����۷f�����Df7��4���_!�����9o�B
�@�&\���ܨ:(��6���6�'sy�j�k�qWVڦ���CY[��N��He:�Wwl��r���%�j�V�.�lWr+M[Nw"�Gg3n����Q9����`�������;�(7v�L�]
��+zu͋{��d�}Z��B]t:���-k��Ry|tu�tj׹aJ�U�lWAR'�;��wUEK��{����<���@J;$`WR�5�5��z�T���ZU�閝fZ\{P���\�豷����-M�J�Y��7�(<�4���3��ƺH��S�(
R��-}/,B�`��0vc��e��
�Ɂ]�*ɫPxR��h�u�C�r
���:�+B���hKX����YpT}� )���J\@?t3�-�[_l�Ŧ]�V�mz8��o���]U���j��z����LukZ��EJ����+�bֺۧx���ͭzժ�n-�8͟�@ DE�x���,ٺ�3�|�r^ �3yՏ:���=��v�vM�tb|��7p��:[�>���|�Pٔj�n�g;�� ��ܠ:ؠ�4n�K�Ѫ�V4�/�Y�ϖ�odx.���v�/{$i�4�w�UX�����zkdSF�瓱��]b��ۿ�إ�M%+���8���R�m��u)x.ؕ��V"�ڑH
����P��S��4.n�7���e�RX�_p��lTI�ڌ��"�n���yrj*}�z��>2��-VQ�e�+�H�|�.�z����(7�&��x�r�׻�]��;`��,,Ҟ����vN#���T�%�j�� 9o@�L*��]n�an��;w�u�	%����Bh��L�ɵS����'jdnr�9�
����hf�ˀ�z�]�@�]�W͝82QY)n}i��JX)uۗz�7Î�i.�E[Ùѕ}�j��3���s@:cu
�Ԍ���Z�iS�\蝭	�,��:��%u
���9%�	Vj��G�g���v��hȻ+j���P�m���X���:�Ss_E2�b�/^��y��r�3��x���r��rvx�䙹�xڥ�Ȏg`*5Ls�'��Wk�F��\��L����w�����.?���vA�ޓ`��O%݇+��¸�tE�eM�ћR���fJմK�W��8�q��t�D�L��

�QE�2N]0�!PĢ�V�ӂ���k.�p��ʓ�QJ�0�L�"ȹU��!d\�2�Y!3D"��9&Up�6�)-Q&D�N�t�d9	�"��H��*�C���h`�j&Q8��AT��((�tK� ����p�Q����4�e�H��i�\�H��G+�#�D�J#(�i�9t�9r�.W
�p/+�u	�P�Q(��Ji$��Tȹ2�ɚ,�=�"�����E�8��$����\.V��r�B�*H�Qp��gH��RHRKCJ.\eQE�H囝\�r�&�p���(�)Y�IQE�*aWe����l������7���(� ����Kڅe���h�����eZZ�}*�̮Ĭe!/'X�}mi9�G#/���NV�unt�|��Ͼ=d�'q	��Ȳ�����w5HR���.묚.��p��!�}b�
��+�-Tƽ/��9w}�6�vk@:K�~+��ˬ����(��*�x���ӆ��M�vj1�դ�M��e�;L��`S�
���>zǍQ�y����+j�)2�]{���+I���{���*k�1/7���z�����+N�[�UL���ldv#OY�2{���ש�z�m-�y��5�9U�|���ɌR��v*V��z̠�`��/2XB�ۋ�5�6a9M�x��(_�²��/
.�p
�> ?��瀺�tB���Q��͆��*�dL�6-��:f��Ńg���>���qk5�	���*�@o⻗�ם#Y�;����i/L�>�Bt�������U�-5^�v�WT���m��
���41���y����%A�:�_�wҍ�yJ����_Y���u~ף��0@vS��g]ӕia��K,�}�vi�R�612m�3��T!�C[�����d��cT���!qڮv�Q����Њ~�� �-�k�n��6T�`�g$��׼)�HK��e>T�Е���жe�j���u���PP��9�5��7����6�ݑ�sA�.E{�l�S��J�`|�Ac6�Zyq��E�Q�v��gN(��z1k��z�|��sս!������x�g"�W�eu������޳u�'�:���3�ے�2gPc���l �z��Ex2B���K��T��7i�+���/h���&�-���f�u�� S�Gʽj�+���?<j�~�uC�d�<OP��=�`���Ϯ�h0�v�V8uR��3��Z<=��4>3�U��O�<}Y�̝H{�%t��cƥP�δꟓ1��œ}����S�u�*�]S3���Xk�RةA]�$ ��=0Ci:�R��ŴU��J$KX�G	�7r�p����3zVmM`�
-�5;�:�Ӂ���!��t@ v�K�M�DT_G�Sݷ���~VӋ/�|x�Ĵ���aO��{��t�HU -�N@�>ҭpu��B��:���M����e�C�Z�y��|i�a�Z�<jt�S�-�I��
f�`ÁyJ�;%�(�~k=�=�AP�<�}[���,��x���1i��vЃ���!>&t�,�V�DB˚)lp,�����j�ҹ/�����߼�՞Z��ufd�Uګ�=�V>  �|�^�����sׂ�>�ץd�a�g�$e,5�f��U��E�r+�/,�\"˾P�y���])�]�c�p��'�c��sɉ�l,��\�A�-���И��b)R�Z�;��ALEY:/���z�*["+Tw����bL��}ț�/�=��iW{�]ݮ�l�9�&}B�]W�T��b���;e��b�'�^b�xX��ڒͺr��K6V�]��Zf��˅x?dv�+�����7^aX�|@}��,�w��%Sס�ҳ{��w��e,�vӸ�V��+��������j�b-�g�@�/ڈ<<����2q^�;7�F��O1@Vg��������g�?�o�[��Uw�?_�mu���&3�O���j9�!�M:��<�6�	jwd$���$n���*�p�i��>Ӳ�g=[�D//I�@Jz�9�@���Aj��j��-tޞ���oUip�$~u\�E�^{M���j#S�أ�u^��T6�d��b@�O�%�8�Z��X��y)j��O�E�1r:��嵺�����Y��Gkf���"T��*��m��`Xg^HU�.pT�S���Yي,����'w�W�c�-:�`.Q�ق�5J#�P�^�����-ڻC�;҇�A���k���rA[;�y����w��UJ<�uOyUt�t_�@�[K��6���mz��a;�q�q9u�*}�e��&���G����%���}ݝos�Ӿ֓����A�{0ٯj����W��x��rX�̑����#��(P�jɯz�t��aK��o����QiƪA�@�����Z7��ل�H���it�`��M��+�.�]�S�ݻW�G!X!�:t��TA�|��2���|���>�W�}�J��K��}���ky3�k���^�_��~u"�]Y�^N���t<)�}��7�0�O��4�v���L9��&�ܸG���E1�ō�J��~GX�U��mp#&�xk�
�1��f�޲�E0� 6��t#m�ou��N8�2��6Y�$*2���t~)1��M��g�Y���U^ծ�W�� J��^3�(X��[�=F���k}���x���ab�����c1��V��4��S�>�T%V�����d�^ÖjW2˯thWv{�E�T�YFK�u�)�^��(z���m�.˺ٸp�[#@��UX�*�m���b���up�9��t��j
�ʄ+�vK�&��@mַq����H�����u%N;����X��֭._��{5�D�D1��ճ[��H�.%�:O
��ͲG���)h�7y�����h!�Q�VG������[�dVϽ��Wؐ�����f������e��arW���.��6�يT���6pF�n�y&@us.�.\�z��VO�����vN������T�Zck��S�3{��vNNu���>��7��ܝ�ܢ��i�f���������b�w"��ܬt��s�'�Ϋ��6���'Fn��MX�NQ��d7
6�Q��j�x��0)��} ��muEq�='1[MH��/t��^]+�;¶�ӣ0�6nB�Mg��t6C�:2ݟt�ܻ�G�^�G������:#���؂�A{~{��'�v���'�����U��x
稞=���g�_u�����~Օ�}�K���F0O�( ��M]��C]\���l�n3e�5>�ө�>s���:|�t&z�e����e=�+���W�#W��X�y�س`�Ƹܺg�2�aT���ة!��m \y*�?�OD������#=*�2�.�1�F�$dd�g�z��]f�fW�d��>���	mS	��d~�2��Y�Ɩ&3=뷼�p��=�.t�B�����?��4��H�����T��`1?���,M�{�a����{ۣ�z�Q�V��p/�cUʦB�P�ێ�:m_��PlP�����	o3�/vd����p�W��@a��^]b�j|@g��	�M�~ߗ�����zI�5LA�F�f��t�-%�+�t�w`s�WX�sۖ:r��j۴3j�+����
��m7k����syDݚ����k���\ޜ�f}�)���2��i��/�*�P����]���Z:�r���&C���i�Vr����|���Q����?@�kz]�� _��� �Uz�>^�"�P_Re�����t�E(U�f�_���?e{�<y�u]? 1�x�p���=Cxρצ]��2��X�]ڲ�Pe�����F	�ʃ��h�\��m�`�λ�d�(Z�o[����K�v�V�=ظ1�o-f�����]�-4�ַ���F�2��\��X&��ĕ�m�Bvh����wl
Ϸq�4H�`�|�Z�a���CRL�;��*�D*��Zس_@��4t�=j��[�Z�5���a��7L��J�S!�#h�8l����&�oo�3�Vy}�e�=�籍���%ڭ���-���f���r���Pd�ř���kB��3ճ$8kzw�5��2�V�!U9��m���|���Ǫ��޽o+�z�ͻ~�/�1����SQ`�k�A��C��;�"���(ED46��R���ǻ>uF�Jt��a�oT�b����TzӶ 5so� �e�<� �: �/�(�Ư-�N@n�d������ n,_��\�wc�-��9��kVcΓId�Y�#�������9b����񻩻�mը���)O�X���Z�&q�(��`\�o%u֞�RH�*�2+1�II[Ӗ���-�}@n�ʗ3��x\Ů�n�u%M9����7�鷙8�t�ې<,��7^F@�XS뵓�F�2Ac�/"�G�V��N���\��]ɮ��V7gf��|iL�����n`!Al>�2x?�:u]�8��R�WE@\�a<pu���m� R�b�۪nO�U��5�V��^r�S�\<�<V�x^��^�k�������C}�<��F�C������������^Bcl�R�B(�6�q��E�d\<Na��ɝ���=*��s����m�*��kO,=�r����U����uG�Mg�DȰ��j��j$l0�����ZgH�tC�G�ϼ�V[�hf��x4Z0G���u���_�gL���w��̽j����=r�jX>>�w�N��Ws�e���ۧTP9F��S�a��N�����_�ΠA��V����R��^-�|���Y���Ј>��T�Q/�/n�{O���w���ʃ�>:�8��Yb}i�D��\H�3��;J��-[/�C=��!�U�l�vשw['X�|a�u�a��UvJZ*�/O\]��>��V�XׇL�Z��L�������$Rk$vh�y��S5���y�-{��'v|ѩ��W���[<
^�t���J~����y2"���(�:��aA#�i��Ě�u�uR�\F�p`���ض��r�p��٤^Y ��ܜ/�ޤHP����*&����@��C�9�B\�K�sN�`�|�ď,eh^}�r��;B�b|z��?%�q��}xy�U�%-Ww*�IΠ�FdOtm{��\����he��;aU�h7K��;��b�rz�C�VU���y�{�*�P�<��T�\q�<)�K��J��E�T�F��I��Dz��ޜ֪�Tū]���n�vSLVnO�K1�
�S0m
���lm����:�3nB�c:𜀠T*�(����D_3��6�ac��κg�M�a�C�i9xf]�Ǉ�[i�#�p�ʬv99�0����s�E����t���n��+�i?:��c�yf>k���Lo��[O:�0]�j(�j�5y��x��� n�i����c=�)��]u����V(��Wx���%xgz�Gqy(߻{N��~�� 2�j�AV�������G!��ȣ��ռX�y���S���ٽ�[�]�af>����`e!��Fӽ���7U�V< �3�'�y���S�v��uz��+}�ó>�!��x���VeY�z{���2�_O`���'p~�uyx�V{s��R�DS��5YLB�;�
u4�u�:\t]�I�ˢ6&��w����t�}�b��e@-��:��JT��yL�^dl*�Ī�=�z���v��3��3,L�oZ�݇x�"��D���b��}1��}��
��*��[61=����zyi�lvR�<�u{�z�I��̎�+3�����B��_�� +�$8\�8'v|7@�K�b�=������.���z��3ٹ>��h��<�>A�g���_u���7��xo��\*fx߷<0n�7�cney]5�hBY�2(f��Q �W'\�f�_W�J�P���.j�9��w�w�YK=�9]��ǐw^�����N�OOu��8�r��-`v[��z�����Ԕ�2�<��LثF�)�-(l��--������¢�,a���T�F�R�z�>�٤�[Z������o�62W��6.������vU���B�ý��&s�Q©�}!Ǣ��䠏��Z���
7�Պ��m��`���͚�%c�������6�LH{�#�����Ր-��h��.�s����6��:5j��f��V��
&!�u��7zۯ�6�)�1����HӲ���w��@��k���m�1�=S8n@�M�f���-�º+���[�l�>R�LG.G+���u�g�9P�c�yҎy�p���֞Q�c��쮫k�Ty�]'h �A�ׁ�Sk�F�|>5�F��`*���Y�/�-��;��;��~�*.3��yX�2�"��@R� ̐�r�w;�%;�ad5x��}�0ww58�^��I@c3�є&p��m!��b���/|���?0)���l"f}d�`��ҋ�$uØ�ݥ2:�߽�y7���E{����MY�3�o]�X���C��u��2]f��Ke���Wc�\�Ա_�:���S��b� �gݘ����U��f�f�)��TƔ�Q�����!n��ڼ>���UZ�g��	��n�7�y'sΖ���"��<�j�]������>7�קʣ$��(k� g�� k�����ͯoWx�#lg���v�B����ܴ0׷]�3<.Ӫ^}�R��:�p���aL��)+mK�BfIH�-�����)>���`WNF�f�z:�����ި�����ʥj��<>�!^���\n�3��
�|�M��6��ԓ�F�Ԡ��>ب����ִ�F�*sH�6�Nl-�o$Ā��!QOXP��v����җ�{�t珰��9��V������Nڽo��$F��B�1�W��w"�8��P ��o����?�c�eok��r�]ڿ�����o�a�hǲ����=u��[�S�e���:,��W+uY+!;9��f�1��w���z�oA�f�L:ر]�Z�nY�W�jCJ�_�:��
�Y�r���b.]+�\'�*�]�\D�A�݉9���JC���Tv�A,�{��Һέ/w��em}m]�\�����Y�j@�>�5�qq�O8��%�΂���&��}�k�m�<&j*�}��,��&�uu�_5��^�g�4@�l�\��y},}��V���:�+dI��g7�V�ST��y�V����9�$@�����D+Wv���4F`�8_s�y�]��ܠ�lA1W1����lkz5ͭ��ݥwEoQ-Yt1�vŪWe��Y6("����;P��tLf^�����A���_Sv��-ݚ�Ya����}ħ}7�t�Y�1���3%h��u�k��ehw�Q1�
��En'
oX�j��u��E���`0lv��i���ܘnbǄ�ו;ZhR�A��QwyK�����	�(ԅ�.Q	���@����iK�O����Eu��˷��.G>�yf�ᵔ{��[�����±,��x34a(3�Pص��}�3�Jpc{��!��5܍b�&z���[ъ�23f�ý�Ǳ��-U���J�k$��kCkT��ҷ{��g-�z���EHa���є���͡Zu�Kc=+�L�B�Wt��i�b�~�Ws���v�1�w�ZΝ��=�u�ڭ�6��4���'��۹�Q�Tj�Ï�+��4M+t6��Μ�BCdw{�t]Y*�qVp&�����ʴ��;'_y��+ �ݬG�D��ã;P�;&��`n�KC��1eK���+*�+�������l	|�q�fM��{߼�}ʲ����j��ө�{Nŉ�H�e]1�n�s�*�-�yn�.���q�W\���W�1�#��ܽ��dX�w8�HX��j��f,r�7��e��:M��@�3����.�p��I8�)�u�v�b�t��V����݋N�Y��T�zK�=�:�PP[6���6��%Jo��ܝ3��k.�JX2lbo5w�P\�(M�]L�� r�ͱ�0�^��N��3/E��7ۀ�K�۽�9��g��$����4��۽���)�]ˍ����X����3�v���cN���J���<9�del�&(]�� �A���M5�9q R��0�z�̩H�� }qu��܁THr�u-5��ܥk�\7�U�:mJ:(JS9S���]H b"Ú'=}ݣ�4�w7�)���ø�ݑc���|-t�W�y��(��	GQ�0�*�v)Ca춆�r\ƨ�.����9��ٳ�>�U.�f�6;�u�7˳��P����]��\h��'p�.�`]���Vl9�l��q�U��,�\��MPS�ϔ��&qs.�fmp���'nk�r��щ�t��ɑS$1Zo,�si�Q�R�;6ݝ�O^��Iu<u2�����=o��<���4����B}�ջVuj/nĩn���!��V�Fo)�|�脨ERt�F�	�*�UA\�r�#V\�BL鏑
*
/9svª*�ʢ8U(����W*�աʒЂ��
",�T�b
��BL�ɧs��v����Q9��*9Ȍ6���p��TeQL���.�ΐ��d�^N{�xe\-IG;��J�*�.wZL���"%G��Ad@��AȢ��*�
5"��Dy�tH��Ev�.�g8*�&¢�QZ,��-J��
��\��TH�Q�"�U����d�H.��J*�*�E��M9vԊ�+�UAIx@yB��|�K����:�fvY]xG@�s��3���-�by�7v��::2�����4�!��w�����4���S����/�yL*�}�l��?]ɿt� ,����<�q��N��?������$���{C¡��M�O\?%�����U�HRO?<�poH��=��6��(��V�o�k�}�����O�|C�r�}�M�	ޝ�߼��pyw�i�~����}&}O��I7ו��p���}O�����`��pO���y��{Oh�M��;ݾ�����`��` op��=����!]�Vn���������>&Prr�?Ss����7�$��o_�{�$��ҾO_�x�nBq����9����N��������ݗnAC�^�z����]O���uI���������p�t��.š�!��ByA��b<�z��_�$�
��	�97���|��>�~NC���>�����yv�;��~�~��N޷��+�4�w���i����p���=���8`=z��SLmo,n�������=�v�{O���''�o+��z�!�����Oem�~M>���o4yL.����x�m����������w���m�������߀�$��ʢG�z3�f!�n]��Ӱ��[�>G��S��ăG!��>�������]�4��=o~8=����ۓ�F���_�?,ro�O�o?����C�k���ˉ��L.��ےM��MJa�@f��CVA��4�]u]l�~|�z�_����9�������'�I!�5[�]�i�����zL*��={�����_���]��!��S�o�Iτ9�Ԝ~q{��ϔ	7�$�w8��9	N�����|��z�z)54-��� �!��8��w�;H�x�?%�w�^LyW�??z�<��O������?�	���8�]�7������>'�®�{��xM�	7��~���!�������NӤ��߿'|��.��bz�H��p���e��H��4���yM�	🝻�`�w�i��o߿y��nӏ�m�<'�o�+��8�����9�vC�i��|�z��b��>�>��T���)������./m������Q= 3�<�����������P$�������r��x@����ğC���<�{I���~1+�&���~�i�	��|v���O{M|���ܚBw��7��~������X�G$���iLGw�Y���A>y���;5iݩ���:yWJ��oo�ͬЗV�������,��R�I�^2�K���q�C3���雰���}���o�o{
F�-�R��y�}�+$�ja�*���̶���j���)
͡Ԉ�&J՗cB|����c�ꬺ�a��x����L/��?;xI7Ǖ����q��}O)��><�w�?'�	/�}��������߿����]�o�ݼ!���8<�߼x_�$~&�v6z0��R
�P�r�H������@e��l.��}�yM�<��z��{=\����!�v޽�����?���fr"��Ɉو�">vK��Ź3*�̴����<�́�7�l���hM�	'��/�o������y@����{�>7��n@�z�cü!�4�ϫ�}B��g���o��;����˴�����>�<��~>%���P
&#�<�m��{�m����sf����bC�i�_������]��?@��o���O�}�)�M��Og�L/����x���$��v=���s��w�������o(x@����~�jw���Q9��y�G{G����#��}��!�4�O�=��Ǥ�!����ϯ&<����_�=x��}������_��?�q��]��}y_G����0����>�����=!ϔ���x@��~����e�NV���T۰7�A��k��ڝ���P�����O�9�����q ���7~��Iɽ!'���^>�z@�������ǔ�	7��{�<8�O߶}u�܇�>�?ןݷ�yv�S����,��ư��n�(�v�gV[�G��R�q���}v��q��C��?��<�}C�x���ߓ�9��}��I����������>������9'o_|v�﯄܁�/��<l��SN��ͱ�p]IF�ڱ���f��A������M�?y����ޝ���yw�����w��M�	������_�	ߓz<^����a}n���o?������r�o��?��oI�������v_��5��\�nS���d3�f!�~�>v�����8�;)��N=����HH��n�����w�V>��?&���=��RC�C���~B�۷x���g_�xt��� 7��i�K\Luu����J�s1q�I���߽xS
a|o?|������Y޼k���̃6�q�W�CHo0���{:j�NL)�׾ǷyC���ϻ�q ���?#�ԓ{B����18������˪��&�V^�Z"�k�@�Z�<;N�7��C.-���-�����`PJ8��Uú���aFoFTrņzS{B�.�:�a0S��U�&Dr�o�Սy���l�L�x;y7�F��Ns��O�%}�I�|������[}�(xM!�������N�?}��?%щ\y<}���ߐ����.	��>>����������X��M�<';y�8ް�7�3vR;e�e�q�{�x�\�V���`0y�38n�s��j̃��';���M�o�Nӥw�׃���ߐ����|�=&��޷�S�(�8��x��w��������Ϗ ��
�4|��X�,}TEW����..`ˎ�꽸��Fy��z,�3w������8��Ct�K� J·�-e��^Zl��т���.��u������ߪ�V+�jó/�g����rUYg�ʮ<��>�i�� ��9c]�6/-���&L�����.�5�����UM�0��}��^}����y{f"l�ؖ�cp:��,F��Z����
�v�ך�|�CuǡA�J�e_��H�/��U����H>P��!��|�|9�C����WB,m�/��HӅG����-H�2J�Y�:_F侕q�zH�р�Y�c斺ٍJ�ɱM��{��V������J�1{Q����M߀癉T��%��#Ryk�����8�Z�a��}�R��p�R�y:�6Ӹ5AR��˸̏��8����ڣ���;�%�@J3g0���,4�g��P�P���	��MӲ:f}M
m����������<�����vgz�IF�#�b���gJ�?~�/=��%>3_4e:w�Lux��1^d�/1R����3k ͞�e9��8S�B�C`i�5�{4�Q:�Cu}�3����'��d�ue�::*3��yC}�k�X}��d\ؼK��������x��y^�Y�bf���}�k�%�ޓ|��ۤi�9�ؼ�,pn�E����|Z�5v:ŘxJX�>�2�ϑq9�2kvqq�q<��ܔR�b2Ʃ���)���U���c�}�����R�3L��3bb��U��I}+����@ALM����uCdj,�;v�i6�
��l��sw��9�5�0��j]F��<�/|��^@VWá�בV����q�^k��4��rk+���jʄ��x��
`G��X"��)�і͈B%l ��1l,m/q^��!/R��Y�:�{1o[T�]�Y�²��N� ��W��AUu�:{��-��j�asZHǖJ�[ 6�_���厼2��U|�(�\��������31��_�/Oa�D.���}�c�+��7����c���^��� �?���1��<��wy���0f���Rʕ�?i�qb3�{0?�w[8r��:���m��
�<�3��ܵ7u~����v���\�T�C;���>�zI!J�w��r2o*
��,��Q����id���&��D��zM����"��q
Ӓb��(ؓ-Ҝ�MΠ8z۝��>��of�c�.7Vzݮ���Z��E*ڄ��9L������p�&�n|�o��_V�W���7�F	�ʃ�Z�d���� ��˲�P�S�o'�7bQ)^vl�u��԰������;�R�cG����j�8-5.��C�g�~d>>�d�5�>{��
s���݁���gؠ!Tm-OXP�[�n�ƉQ�m�f�-��ˍg57��l��A����d��{��+6:��o����?�c�eok�8�M�ޣIM�1������ �F��د������'[۳��F쥍�ĺ�ꆱ��C^���d1�*��Q�lx­>%�dbX>��B2�^��·�*�<;��E�V��]��{�)�ջ�ݶV�\>��P�S��K���f�44��1Ѥ�[�gm,Ƈ�D�E�mV�"��$
HU=��+���ǽk#��4� �G\�N%0B�n����&��L����M�����Fq�~u=�.��oXu�����Jo��ֽC�z��&:å�h�Q��yz[ëy<��p`����J��0b5���o�L�P��k"�U����<���PAR��ExԮan���|����+pRt�Cn�t�Γ�������:�8l(,�Ӌr������� �n�ؖ��U�[7&9G�eVI`���`�GP��.R��Pr��m�����6���bH������Ns�y�����@o0R�!�[tܟ\��]��j��8�+>U��}z��a���<}��kӦ�XG�<�O$+�������u�0ud��^�t�2}p�v{��p<�j��%���$c���U�?�����/�U�@��y"6����Z>f*��/R�a�r]�i(}�oa��Yf�a��
��P�e>}�D�Q�r�
������
�pt��&Nד;)z������\��ʦri��o:PU���
CӖW��>��t�^��n�]w71��:����]D=��j���U�u�2����HV;����\�=��<�o�ɾɶ+oz������
�|>���N�[��g��*���p�^8;��4����'V��Ǣy<�vj"�L�5�&_�X7�Y=�)�UvJ�������%��2��ZM�&� ���,�i(m�[�C.�h�
*���2�
�)�I�����לE\d��e�V�(���ި繉�����U���o��Y�^�=�Xr�gE1U�h7Nx��}F�D�}6��xd�א�FPNn��vG�fV's�e;]���S�*e�����k�<��b�j���}5�R=a抽�7�)��Z��ɻ�4:��,����[[��g ��/���xr`»n�3ն	3�����+�&���+��K�n�D>����?]�����Uw,~�;�h����^����<�g^�6�,I�����^�)Vx�=�����B�횱]��X=Ǫ�Q��W���8s3`Ǔ�G�����$�X�H	�>�E��wD��3���n�Y
�ׯ*,��_�yd�d՞��m趫�3�/�]�.��0ue�{/�i?K��Y�^Oݽ�a*�rՅ��m"`!��?��X]�G>&�ܼ��x�R)��,o2W_�o��䒞��-V�M�����Z6�>�Uzv!�V;�`  ����O���x�=Sj�6���}<���:���tud.F;�n7�V)<5X|���Wo���D�D�答j���:3JG7���M�������'�Zǂ�U�����yK6���J��+����K�����ƱS�P����l��Vs��`�S����VuҫW��>�b�/���h{&� pC¤徹y7��)�׺�d�=��n*�48Q���s�F��U�8qzR�W�s�Hp��e��W7�`a$l9���O]�5��tf�p\��K�o2$�׏�|�,�/��8h{g|Fvv�ӹJ�+<�|����v<�j����$S��k�ւ�C"�0�+;��$"�Sw:$u�n���v�q�GE�fp��Boq�����$�������v��}�o������2�Qi£͍��-Č�t�0�Q"
ț�P*!� n��4^�lO�Z�cB�����0+_���W'�v�f�
0�^z=EkՏ�7�}-Y�U�����{�m�l��6����46�ҧ짍9Lװ@���2&�F�Z�e��3a������td�K�<�wNK��4f�am¨��e����ތꚂ�9G#!�t���4;�Bp��;n�fY_=�AZ��G�B�����Oc3��|b���w�=\��y��3���5��p�5�f��ʬT�v�<�`�K�%�KU�C]E��ҌUNم��Q��mb_f�G�L�i�*���p�$B��Y�s���S+��^��P�̜o��Q���a�V�b��%�t�6; BU �N� C��d2/�F�03�0��oHĬOq�o��{�X�.SY�V%�c��U�2e�8��t@�[��z?"����l�(P�=�]d��NgW+� \��\Y�X��Y�L�Z����-z��0ױ&T�H�d[T-���@nh�S�oq~}�Fr<��~<P��}�P��Vƽ����%0w=[Cܘ��!��n�ԸҚ�4r���E[�����Zt:�1�ay��(��#:��׊���g����-��1��@5ܨg
�Ռ�R�#��Md����)�j�s���1�^:+s�f]޺]�Q,z2ұc��V<)��X
��]��ׅѵT����P�Ir�>y]J�����.860��H+�{��f����xi�xx]
˾^p�Z��f��Ј�#V�kUcD� �a��O�%)y<���B�|ok��y�+���z��������f�m1�o�81�K�k�+}=��	�ϳ��"��3<.���=n�&�@E:Oq����v�i�6�MF�b,���cf�h1��V�fI�`�z-7����j��fu�d����EY��};�t��ia���xϰ��*���n��A�k�d#�3L{�l�E,���ѕ����l�W���]�=�{g]��_t}�J�zxJ��G�b��.����4ڝaRZa�c��*/R[���z�X��O���f��:�u �[⧩�KCI���nG��R�('�*�mD�6�V>�-T)d0���J$e�L��c&���U���õHV����x$��J�d�0;P����������"�U>H{���maC�;5[أ�b�?]�I�\�A/\�}]0�-���Ծ�ú�>}�N{{�|��гM�GR����ǋ{C��Wwb8Պ�+�����t��q./,��*>ͺ�j����K��5	���kX�k_V��;�-y*�D^;�gT�Q� ��a�5]��)G;Pս�<�Mmd���D�o����yݺؕ{�x�9���}=%��mp���D46�cS��#(Ʃ��v}��zϝ���}:iX3����6�G� j:�Y�@)T���TI���uXEl�)�l M��cp���i�>�*� v�{ ;n����t���DT�n^R��FE �[�#�u�h��u^��zU��p��Vu���H�Q��^(m)`vy���o����\�������@Z�=�i&��jC[mN��^���!4�}ʢq��n%*��8,a'�r���W���k�<�A{���+�y���� �8�74���S��x�y��^�׫_ Zx=J����x���u�*��������eW<yk�gz�y���Y�]^S�֍/����E�Ӧ�̀!��A�c,y"YT5��*�d��|ij��
)BQKg0Or ���^@G���.ZY���Y��5�W{�w��t��X��dg'L���4㥽;`�C��ԃ�^ժ�U�7n�S\J�ϭ/i�$U�/��pW��r�~�����k"�z����5���Yէ��.%������$�1$Ѻ=,�Pڰ4�{ɸ�WU��<��vu��s��)4�ͻ�7�e��V(��x��t����d�y��TX(JoK�ي��5˅�� |���֩����@aoi��b��
�{.+���Jfw8�1e�%u+<3��ʳi�
D80���evM�9�!�i�sU>)n �w�䨚T �{��s���Je���N�pg#�\;F�[M�$jwГ����q�볳p�ȊA ���L��j4��ԯ�4o�ȂEwA&p�P���&`�]�H��Ǭ�!n���n�wAp򡶚Υ3����F�_v��F�n¬�
�2��e}%ӋlH���X�!�Wm�k�;���o2˚�����7\xZA6 ƌn����*\8��D�n�,�x�6�oJ��0��M�ˤ;���Z��l���m��Z��T�B�Ή-�U	Gq+�)�s��z.�DJ�s��H��{F�:�f��\uŀ���/��K%���yZJ��wfi�|���OU���"�%ԑY;D��BPw��펬K��_Z�x�"��u:���b8����/I���SlϹ^�-,��Щ��ү��ۥ���F�:��-W\%=����\n�&Jٔ;�3�vq<~T�-���6�J��غ낹C&����M�Z�uq�,�]N������6�Ǩ�5���T-\i6	�����-�$slpR��Z��p�$,t/*���@�k�r��4�Cq:�֠����;���XCꔦu���c��Y�<Z1������}n�<��&��vҗ�zc�އcYj0hab�ۚ�r��Qm��q�@���[�S��Kdʵ��M�sE<BCR�y\�����zmfW,ŗ3� ��Or��1R潸�|2���Lٙe�*�.�K���rɽ1+	\�m�
���v���{�
�U:wLf�N���4f�Θ$���� �7z�\b:'�U�������ţX;���f���QS��Ԙ�f�V�kN��qa��t�	�!�׃���ö�򬘫y���*�<'2�՝5ol(�F�!π�3�;0G�]�q'����PZ��^�#88D���GSYP�V�e�����Wtx���]n������C�*��Ϭ�:�3�c�D��<v�:ڊ+����e�`�]��ܺ�j���l˳��if��A�[�U�GQi�C��[zB��̗���qU�n�sz�����t�ul�H�*�L�hfAX�� SCi݊P�4'cDS�ɧiaE�/��vZ����Q�1��44M 	K��gy�b�ဩ3��ՙt����[��Wg��5�ig7k�qY�v�>��/���HJ��m���e�	u��)�paR��i�J����U\��_M����Q�wI��w��M+2��3�W�Q^��P�AuA�W����2�yPR�I�IH*"��j_ay��T��`S(�,��UEAW#��ZUpww
��@���\T(+,iJAp)�reҸ��v\�DE�YDf*Ft����˧B*��E�0͔rIVӅP�r�g<��������Q	˄W�ԙr�28QvQqѹ����UrNU�+�.QsE\�K��i��6¼�9pJ����*�˜�Ny�젪(.Ah�B�L�*R4�vPڬ"��wK�"�2�r�Ԩ"��NwP���˔Q �� *�"�k=�u\���V�z��������y"S%h����1��2Ʈ�"����c�x�wF�1L皴WVoq��o�m(��/l�5��\��]�Vܜ>�A�F��:�@�ڍ�UZU��}�c���s�3b���`eμ��C���l斸:(����Z�-]�UvJ��������[��h:6��5-t�ڎ����cխp�Yδ<�C.����>Q0�<�"��$�D�)�Y3�x�}�N���$T��ڲ�"�n.�Y^�}��[	�u��f�f����ˆ�˹������ȉ���A�P�s���O˜O���{گuWw��5Խ��4����I^��ۣ��;�ȱjV��yR�h���@L����%�R���cL���2��v�v:sN��W�)�/�}�0q��}f:���@=G��yR�m�a�Y�N^×@��d
iq��4%,��dɧ7$ִe�!���ޟS���Z�=�|�u��^p��FQu��y}~�)��o}��Y�GW�\�tS��rlz�`
?ox�)�㮑Lg�%v��sG!����Ee����t�����*]�YSd�!��l !��m��D�X���y�?��c�{�߲�x�^�A��{KpY�\��� 8v���F�f�XV*�j�_0L���Y d�+��߅�AS�fz�޸!a����:�v�e����1��q��oe Ȕ舢{���hB��tT���������y	AoqL�����.p�Ξn*��2��.�c�ڵ����pUL^u�eN [i@�N�W473.[S��8�������=xKhՍ�F����J�}�jó/��-%U�}<�n.�&+x�mη��{�T�o�K��O��#,�4E^��v|71S����h{%k�%縔g�^�����V������d���l,��;e3���S��M�d�q+�~@Wu���5ޓw�q$@��ؑ�c�]ԕx�}�|��`��<��qؽ>��_IMӮ
�)�)��oQ3"��wњp���斺ٍK(U���d`m���^@�z��J�[�a�[�b����B���9���CC3򂏏x̊���Vk�,��\)�ܧ����{��W��F��'�d/ڎM�N������.�h��a�[~��8�(�Ӧ��+�b�Wx�����n"/7D��Tc�δ�@V5���]r���{����
��O��Z�gս�W�m˵��{Qq>5N���k�Y��ժX7/�����Z�4i�e}�{�Q����4[ �)�9R!E.(Y�C>\ߵW
x�s?A�1���wz5h��:m3E�3 2�k�6�Z�en�tS{��I]���F��wo#*6kn��/;�(���Ҿ�Is���>�n^�qg�L@���]��&�D���G��}T7I����
_N��=e'a���b-���h��^}QY,i��P��|L�0޻
F���KC�S8�b�,�M��|�]:Y 2ҩh��.���d"��7��1+}8����1��z�62���;1���5�[�l0�-��m�ke;C8Ԧ^n��R���J�[��G�)w�=��ϻ̝�]&N��-���ݨ���1J�q�M!W����=+ќ�-�I◞�v2�x<K �B�,�UV�n�kPL��9u��}�_m����ױ�Z<�'���l���qH��%�ܝ���K���ߧ�h���1�8�ɳU���oj�J�b�^���ƕ��66꽕�O
�?q����=G��tY�9y��x��-�a���tT�ֳ�_5j���TmP�
��K-cc��7t��[t:gX�搻h�NwΗ��͝�3Z���T��a�ʶ*���4�Э4���S/n�o]p���dQ�%����:��E���3K���Ҟ��爱�z�Z������X�,�gʝ7[O���Ҧ�Y���7�6��j�T͈Mb	�hV�3_w�,�Ξή�\�;�UW�W���H�{l1l���[�����z2{�v
��nnaƂ8=�����\y<��q��q�{Վ��ӯ5��mQ�O}��\u��Y�7��Q���қd�)l27f�nǑ֨b���k~&xRٜ�l>�6t�^�5��P�m|/�P�O�f�IkܗOT�M��r����>���%:�Ľz���R�Ƶ*m�ʁ^�}0�Yl�	��[��+C�wvZ~�WS6rC��d�����|��_�6?�R$���0ws1�b�bV�,�+�9҆���i��1Q�6j�SC^��0M��i��{�ݪVD�U��/%,�4��ܶ%�j�E�i�/;I�i�!�c0BSU��5���gdh��tش��M��H�e�ĺ�Ǫ�j�[@��b�ږ���ͱ)d��M���l�T2OJF�kL����=��cUZ!;��k����\��]�a:I�o�v���n�Z�����g��[Wy)�O��;r�F�q�Ά��4���~�&�.�F��۴��6m�c��8�����.�QK���rhz����]i���92�:[��G��Vm'9&y^�F�19�~����鮎��
�ɘ5[��������=���o��1�e��9���{��AG7}�.|���^�o�,K�*��[mBlͤ�%�]��avIU���_9��d�$�W�ʆ��s����u.�<��P�޼��\nG���frj�=��^���������c�lz'�/mN�c������^��v�X49��ho�6!竽�׼�B�y��z���YPÛD9%b����_����с�fò����>d5�s������L��E56�J�j�X�T�i4��R��׸�Z��-�O	N:۰��mہ�[�3���^�qC�S��kz=;1�j>��	�c�b}D庭j"]�y����W)��������l�G�*����[�*��P�'w0�U:����y�$�ۡi�m����g�xJfXF�UxjfeOja?e�z��#҆��fCB��=�����c*Y��,�!y��ޝ��ۍ�y\�6��E�DsF:�Պ�2�eZ�����Q�%j{{9�*�U�:�5��U)&V�S^;,��.<Y|��Z͗d2#�"���m�k�S�V&mM���΢��o��꯫�
La֭z�ku�6��rlWN�^��3�f�̶;*@��Y�⊭
򼇆k�����tZ�5�/{U�P�٢d+rj�/j2��'i��6\��V��[���1ҕ{��kk�蕑�%��^cfn�։|y}�ҼՔ��z���m1P�R���t&4����ս]Z�"R��T�}�1s4ZO-�ޱ�����N�H�FI[[�^�Ȩ|�l{�N/YKk�m�a�OJ��U�I�jT�׬[Z�Jk�Ն����]��m��*�~��x�=���U첶�/s�WI���/o���SE�T�xFޛȽ��Y�4c/^Ĕ��-��+�q�Cm��Κ�j��'Ʉ�6m-�Z�+���sNl,X̞v�׼��gc�g�!X���|a���OP�ۀ{�=PL�|�IOە=:��׋�d�nO���σ:��/4�x=c:�]�/���g	u��ǺQ���Z��a��"���u��Op�t`ވzQj���F�c}�r�o.o���w��CO����p�:�sҸaޒY���
Os%��)ݍ����|f�	Vt��T�81,��æ!;f�9��{@�T���T�?`w�BҞߨ����E1Qs�]�;	��JqP�����<�l�=��􃫱��_VN���{�纜oT���Gc߯�-��{݊��O�~Bo�T��+���-�����~>܆���i7j��Qk"66r)-9M���/vXT�fO���m-�"i�Y2�7(M#H���˖�t��0�i!Ko�P��[�4n��Z�c�Z�KE�YY��I�,��J�*�Eݡ[3>
^�v�|��Lk�m�F�ir���<�}F�nn�WS}w:z��3I����3W�#�Z|M�
d�)b�vݐȡAM־��8x:�����}�ߑa�#�ʦ_>�2k1��V���j.�w��dؔ�7��ng��OK�i󱔼>y�P�9^V+9<�5��<o�Q�$�z�?%}�o�=r��9N���t�@���&1�!f����D5��]Z�re�}Fʿ�]����v�����b�Oy�k#L{���w�����߻�7{r��!�gǻ8)��X�v5>�*ts��[���t�k�:��I؍rH���yǜN��<�w���@�w|����ɝS��[��5{&f���������n�صs!ۛ���N �T�����?{�t!�����q�B��҉��L&J�&�mN׬qB��{,�i�ս�+lװ��vPz_^�hg�_�un	%�j�xi5�Z�AD�k^b;P�u��W���s���l����}S��K��Į����6�]�zqc���8&N�Y������o��X�Nxr����\��U�^<N��ƞ�k�'���o��s���a9�����~�9���2��f��<kI����LKE�՘3�z�����6q3꽖d���R��~�#vh�ﯨ���,����hBSs!t�Nz��	�x�ʞojs���eo������+�~B�4��o��L�ǆ���7v����D���e��O�Yk��ӄ����{}�M����G�� u���/b��=R�q�ҵi�j��ؖ�p0���� ��CY��N(q��py�����c[�:]�;%$C6�9�xN��3
��O�͗-����'�p�M<SG,����3k�SC	yg!��:�	��%+��}�s�v�vD�Gzb����#0젨d�����+S"������y������[��(��0�ܭ6�ji�1Q�6j�����Ǉ�>��ص�kj��)��'��{�z8���lKڪn�����Y�To,̙�z���y	 ��F;�#i�ء9�}e�K��3�R�Kʒ
R��ˬ�lpu���L�B��L�}i�HS�w$�L�ɵ[h�1��!L�{�ë��-�#V/}-O�Q��(�:Ѷ��OF��5���3�-y��nu�M��SԖ-�z����ֺR�ٯmC%�p���^���e���ۤ�>��t_T�_yk�I��[�����IKpZ�;k�þ�^��3o��O�bWu,=�o�/i�N�c��\>U7Nvms���'3��r��ݵ+v�Z�������6����Ĝ�4i�r۹fUՍ�0�N*�_q{J��Sӣ\{��ذ�WO:�W3�E^B��ir6�����
�z����:�6��0Ą�n����"�go%���]C5����W���������A݃Ê&�K�{��c�U��ˈJ�h����N;���P�
έYJ`f�����t���"�Kq�\�z�=��A^�]x�E+~�TIΚ��򪾯������(��fv����O��ގ{�NG�?[�{T}����ޕoz��M�֝w9��J{;���Q3�Ot�;�N7�>f���{}�Zx��?d��#���{��.�pۮ^��-yğ����B�_���`��=k���T3}R�������u��,֗v���v)d�ܪ���wz��e���&+f��}�q+�P�m��*Di�Ե��QlWN�M�fF��Zf�C)�U�)>���eO��V�lt�	S�A��e���\�2�m����n���.̛�
�{�(lU�r��վ�X�g[�g�YSP=�^�n��U)L�n�omy�n�Z����/����_N�)��Ҕƌ94�lgt��̆���mC�̾��~g1�?����?;�����F��"�9�ծ�5㰹�U��m�>XW��;;l,�ež��h$���iw��}PuO�c�{�����j�m�1����j�[�b1�v�JK�U�T8��x�|,₀�6���<�}o�-�Z�-X:��.���u�l�}`�x��xcB�*.jE��Z�U{�7��[�7h�hI˓�8ĸ�&�r��ɼ���Ԝonr��A�9Z�vz�}�fW<�"���]2�ɤe!ƌn�:�ޝ��m,v:�������#؞Θ�[��;�қ���m�����$��9���둌���d�Q�k6�S��{v�i�{b��/N��oP�g_q��q�-H{&tmWd9{�m�cq:����=;u�d�u��(]I�u�ΌP.�8w��I\��Z%e��[4SHQ���F��f����G8b�t#W�Uԣ���r�7� ��z:�D՝�.�v��:�տ�M\%���*�w�`疍sf�y*l�St�ʙ�_\32����w�uX�du�>B�
v�ޡ'Tz:tEbt�Q/�5c/`�<�m��t7oQ2��Y�8������k&й+�C�`�/�C��1�[�}|���Iv1u%s~�]�����]�:�W{OD��܁�y��mL��������SĤ�3k�m^�V9W2�Q��a�Tߓ�e7t���
y��<�0��6�gv�杬uט�F�8:��M�[;;u���u	�wJ�Df,	���5��B�P;Aı�cj�x��$����|����V�]�S���c���d���%/B�2�yļ|[Ǵ�{��'Ww�ά�t����Q��S�cq����/(;�p���EH��We=r=̊J�"m^V�+տbNd>��j��*�����v���\
u˚G&p]Hz��)�ŤZL��ň��4-C��
�/�ė�
��2�vpً�è�;�P�ܯ>k6�O��Z&U���\/&���
��v�	���Lp%HQ�I�듶�S�w�BcSNjs8�T(ly՘����\L��x���j��ŷZ�Z��<
R��N�z)M���U�$LN�km7��VL|c�X��!ܭ\�9�w���Q�ig�f_�4]�Ӂ!Y{�ĩ��6��xs���6�od���m�˹��輸���.,��g�^5,#0;�@���I7ѭ�s��YS��M���ل�
ƸY|)	W O:ȯ��v<�y�&(����v̫����%�g�iV��²����_P�)%w��:��D��d��.���Z�-�Vs@��	T�`���>����נL�㑊Ԕ�)��W�����3��T�6��g�7E����>B�� :��Мg,G�Kq/�ŧV��o�3��x��n���Z�j")A�;A}P�1$�r1����ָ[����]������{��|��i��ؑM$�I9QʪdBK"�oN'
�8\.\�DDd�\.�.ɡ˔u�TPzNET*J�3���PS
ŉ*�BUW#=��̚Z'��#VĒ"�U�U�������dvQfp��(G(��D��C�LU����s��*��]rB ����R,ʜ�EQTP�9DM-H�N9$�zbs\u���-CJ�'�(�˲���"u���.��:L.$W)2ndPG�Ba*�;u��̼���ȧ8\�
N	�T٣��8Wj�d!��=L�DB2r�0�e��e{��L��P�89�@��nUM���8�	�L��g������#OD8����st^ޗu��1=�w��c;6���ލ�=�+i�^G�;��C�[=�5o�0�5�}_}_W�|�]�������>OO��T�	e��;^Z����]K�PX�F�<�jw�2JKY���n��oqY�y�{ܭ�^Į�Գ�Z�<�^��ݎmuY)��c}����ߩ�[��	ӆ�aV�;x�(dJ���dbB�,�k]b�|Bh�fl:i4�J�cw-C�)f�gzvk���~�l>^C�*�]0�;�U5�zƽǍi3���4��_n}G��ܕX�s�d-ׇ��]��k�We7������!��<h�����}ۓ�3���Z�_����~�6���ީ��B�o�W�ɋ~��kI�4��k�/W>[)K$ݻ>P�x�ZV�|�S�i�I�9]wD*s߷]ך�i>��'xit�Ǌ���kb���Д4��Z�&[E�oS���X�j�U��[��d�2Mˎ�[��=�fֺ�/�ޭ~�
�g�]��p�9��Y�&��z�J���ά$��|=[�'�}�iK�%���P�r��|�D�u�/�(�l�]b��C�����s.��ҮLfj���»(v�w0�7\�Q�v�iTV�ʀ��W}4�.�Y"�܃O�P�-q4uݿ�aj��ztR5�������?���}��V�<9�;�+_�cy���UD�������mZw�M�u�9zkw�B��TB�ZU*v�f����vb^���,j�/[I�֩��5�@�:����q��sAd�ͮ��Kn�'<��\��5A%��?�󱋽���~��a�o��]�M,�4�ۺT#������]���,���-q�,L��cW���������^1fO��eiR�JJ�=�A�Dd޽�ؙb�I�JDTn��@T�̓*�Vǚ�S�f�	�_U�%4�V/RC.,�nZ�S�zx���9{D�S�z�'D)�KԻX��}S������$�kO(}n��'��J�A�),��)��^��ͪ!v��j��S����_��^��{��9�*Q���j2�W{�lu�]jF��v��s�<^�c�]6MNR�#��}62�:��^]4n�d�[��d��_[p쫯OJI����ާ�S̍�l��!�fb��N���>�]��<l�����Ӿ����I��I��2�o -Q+(�a�y�s���@,��;�g���ǣܱ�G��Z��4P�$8@��Ʀ,T�woR�.��\�shgW��Y��*�rZ��t2R+�UΥB{uQ}��q���^��A>�I~���f��D�c�.�5͑�{�z��Զ�<$�۴�%��n(�{��6�em{���++B�S/�������^�����n��Qm�q�lK�|Ǥ�V��=�k�ě=�y�jR�7��|iv�|o@D�z����s����y1�)���lVZi�,��U^���|��Z�M.���W����=���<�o+�살J��[�[�s�W;ْ�E�l��~n��ZU@����hmJa-��ny�1��#W+с������(g˗���<}^N742��ݍxف���˻blP���m5���^��Fx�OyJ�~�������T�V�5�Q+ְ��u�Bv�LT2OJ|6b-H%��Ym�^U,}�e'��J���cs-T����٫Z�W�u������!��"�,;���]{u�g��vL�{�~\�I���-]K��>�3�+==N�;=�N?kαfP�K��U_vb��e7[n{/Xpum�-���ic������}�����S6&#���|h� _�Kv�+8���i�kTR��[���s|2�n�%���{�x�EuB�g8�u)Rv��g��諭��]��r�P����[Ba�Q��'Y-�g��OWQ�Lyj}@Y��z���'w�!�-�4To����f��6�%q��T2|�����0�iG�6i��*o�Eu4�LkHyb�6fi��J[nJ���:�8l^�U��
�������s0���MBMsb�����Wn�~�ro*ɳ:��n����o(g�.T�2ӫ,��4ͩV\n�^��V���f�%8��]�|���0��?�rt'�W3�v&=��<'Ǻi�τKi�[U�v�9^��-�O{ôP{c�%�v|+�T
��bߞq&����B�A���ߗ�;�.�����7x.��0����,��g3�,[C�$��I_{��k9�����U5�*S1�P1X�f�����G��g)7�|+�o���f{���܍�a�V���/N�{k|��[�>S�xjӅ6[%L���i����[�\��W�pn�.
qch)]C��7�V�mcyh-�\FU��I�L��5U�����T�U�����~��:T	�lxn�S.>�Wڳ��Ch�� ��GU�F=ΫR�i��6�	����:x�f���{�/�'A�qa쥵�����;�]�Z���t��aeK��v���?������ٻ�l�i5{6An�����#e��w�M�u���J\��xVœ�nldM,�Í��uuO�jjlҠgU���'��^���k0���;�D���-e�o��9W�R��~	/#�:~v2�u
y�lՀ���u�����prb���ѐ�Y�s;�HCͯ{G3A��P-� ��ci�w��W��t��Cޢݗ^�
��>��+6��w�A�һ;���4��O���ouC�mX�2��V5?�5ѝ���{��3m�{�w%��yꆥ�٧֓��&jl�^VoL�@�z�F<���T��{|���.���>C���{n,�e�5榣��7D'Tʲ�҉+6Z���7[u;6�ee&�3Le�T�5��1���vױ.��^�t���Dt����s����a�����o�������C^0vJ������-�Y:S�M�u;�/p�G��(_D1���K���7���)��b�B�e�d���bd2֋�g�y�a�X����o/�8/˰i����c׬�oM�x��q��6h�a�f򩽓Cnػ�f��o��5ץ��
����k3�^�n6nu���Wu��������\���;�����u�\�(a�wg�Wv���� )��z
/���e��Sy)�����ܪ^ͥ���B�-	!�E�b�������I�݊x���ح㽻L�/i����[P��e@��},���{n�TMf�݋[�E�E��jBڙ`�fXl��Z�{��Z\�l��J'=�򫕻r�g��bg
�t��xl橺��e?�{2�GJ���T=[�ޖ�Lv��/��v���Z�,��cKm�aq�%�$�.^���eTz:���ʵiCD��[�f74�ͶR����`����g3|�����;ˮww��:�� ��Y��A�-P�#Ք��eXڍ~6{�-�?#A%�MH{մ0�h���rs�1�NP���1z�P|�}��'�6��^U�z�~-~�{k�Z	�]�ĽG˨��'�ս�|kЬڥt,�_U�ң��iį�(Z�C36�X�#���d5�v�۸r��.&�uK�E9��V��JS{���%�f8S�u���G���p��}e5Y���܏.��R�)Xk6��
t�$�i^7��f�I�Չ�7v,Hb�G���\��Lw�H�;S�
]��[u�^A�����y�ӁM��$��3����tǖ<D/j�]�ǒ}N�xd���>ŝ�n�H����wt���#�y�5I_v��SN����֒�f��Z���*���J�>	Y�c$����ym��h}�ם�T�l�4���Y)k%w3tn�ñ��C��f�>�O3i�e[6�h�a��rJϼ|i��6ѥ����è��3u5��^�C^��j[p��)�#v}E�wë��W*�X~�y�c)<�(a���=�CL�a�nCM��,Ȭ�J�.���afF�F��t^��3��)t�k���r���	�=�y�-s����艾��o�p��a^Q{�ޢ�B�5o�U���
|�+Y��&��J��������;�Uu�Ek>��Ԉ�֦٣3ҋ���w��u��β�N�es��_Om�ffh͚�
�c�ذ�ĥ�6h��XΗ��?����3�2kU��GK}|��iG�����}ί���bsJ�pV�ݤ�Eyyeܤ�?v�Y���.ʋ��ʖp�Q�i�[��ܹ�snWe���Z�uz�nV��%m�8�v��Z�mqT*_u\z� gK�j�U�S7�V�F%���k|{��7�w�ذ����K��}^�TJ�JZ��n�7'�ݻ��
�0��������v������LT$��a�Ԃn2�|[/��r�im�L�j�ƪ����=Z���FCζ���S�l�a�Ǻ"g1E��-��d�e�9����[�K�>o�L�~�Uynz�n�/�J�7�=[��k�Y��>�*v^������~]K���}��d��S�}ԙ�^�4����ʫ���'oy+�ױ+���=�m���:�4%��{�ͫtL;��Vv�>+ӻ
��n<��̤�6���uM�cH��ӘEd��*WOId\S���vvY݆��ś�[:��A�]�g;v����:<O��JPC^��Gg��Gw������E�rs7S'�Z�i>n�dV����6D#��p���4vx3�6��U8��(��R�;^�qP��mc��n����V^1C��M���崜��������ŕ��rbu��F��dg|Y�͔;o��|5����������A��b���3h�sC�.U���]�sSA���cNQ���Q[�믍�'�i=�|����oS�IGr��7 �(���>�n�HJ�k=�^q&�A�tҝ����]{V]u-����F��8ў�����>�a'Ҩ2��Ql۟3��1JfDnU(��6��sb��P���^��1���M�*CF�j��[�֮j�C�ɰ�i�sSۍּ���}~_8�4��mk�ՍLϰ�A�ݭs` ���Ĳ}}�e���E�c���Z��qR�a��l��̞���OW���y�­�p�g�ggiՎ����r^��K��]�6�<!;m�)��Ȍ�5�`�S�w-6<DZz���3�p�3$ݷ,�}b�U�W\3Z�^���P7h�بmV4KnI�ڝq��l<��\^��|�)w���RǍQ�E���m�rm�Z�
��������Eo݌��_JD\�OpQ��
6��ĘLۦ�ԡ���1̈́w��>>�k�[�6��%s�WV�!����v��ȷȊUy�Ұ�G.�5��0b�Qf�.
c��V�024^�A^�?x�B9r�B�VH�lmZ΃^L�D�{�Sۡ�y{m��8�r�ꚲ�<˾�=
��8���
��џf�����Еe���x�Ku]s�{]����κҿ��������8gz� Q���'9�[6kL[/F��K��3�
	����͜lY9X2whb���|B�#ӝ�G����q�*=�{[WsO�����@ÎS|�OWa�dT�vZ&sc�w��5�L1�zM�Z��֍K�cY���[��S���yz�k��䕕s���8�zwrI�R�JO�YFckF�M��-,�jMO�P����A�q�d�S�5��R��ŵ�z_QY�˽����a���͵�̬S0�B}�ۮ�PԢb�mI������R�ܹgJ^�Z�.�-�
�慹*Cƾ���i��:���w�.p�:��
�5�rx�BM_�~~вm��h�TPf$�5��;�r�M�!�-A��u��0{W5o�^�y�W�*�_?	��V�+*L�~T�爻K�}e�K>�"�㌲���ej��U��<����"�V6�T8bg�Y[�*�Ȧ��f+�Cz�+��R�#K*�jcz��¦�L���&��Ԡ������p��k"�)_��]�rQ�o��ΕB�a"�ns�(빢��WQKdgu���)�_#Xh�}ϲ�wM��v֧X�Пu�煰�$QL�ݺ�dfv@EwtL,
EWq.�u�&�3��,�ׯ�
0%�;H�mT�X���m�76��yj�o������yE�T�33n�d�����Q��āь�m��,�5Ԓ����#���ٛ�rն��7[�FPT�a�ٱ�`��|�Xp��ͼo+l����F�ޗ1�vҾ�7!�����[Թ"���\�u�)C\fV=^;����]L䩀�ˍ��{d�o5�n��.�'f`@���YW�"fN'��;J|��i�X�����*�2�G\��\�Rw�ݗ����t��i��{K���b��5q&�i�n粰�����(��[K���̧�IX��-=��P��C�f�M�
c�Kυ�_r��ݪ���HV3}�E?�rD0�Ζ���B�d�eXM��۩���tc|�A��%1�(��ʲ���Υ�p5��U�SU�6k�.�Z��Э��'qd���,.a��C�Y�gws��3]�
�x;n�ln���ze�ǰRnK-U��hh)��W��w`�\Փ��봷}�tj:�r�S���9�V�m�=��ĻeV��UǄWa�s�̬�!;���2�Os�p�pKu�S�y������n�ԡ>1�sK�-ٲ����WL���l�ų�T�p>j�Q�x�'�s���.�h���oy3Ӄ�:K�=pV<k.��9E-R��8Z�,�>�u�����c��+�@�t�4~hөȄI���&���V�*pܙ�)	�A]Ϩ&��dU��d!��a��o�_3&�� K4Y�k��l�����X�c���[nP�Ky(������}�N�����ξ��Z}j������<��v���Į-�woc��h�=��ڵR4W��S]�B�o�1&�9N��&h�w����ŴvXZ�,t��;RDв\[j�w��������j��ҥi�����n�F�nn��&�	�X�Q"ګ�����Q�#o�L�f�l�X�'8����!�.|1��j����eͷs:RF�RT��TF`Km)��5����X�u�
�]%7ql��t�V�>f�(j�e�Z$U��3���S���*W[�I��VSGyp��{�2"�N�n�6�J��a
��1���v�Y�Q H�@_c�i�Ľ7)ϪYe�&nI�y���� 
��n���l�V.%؊���CF�>���:ej�.*��p��k�dF�	n8�@���فTr��'8�T������T�c�T�"Ĳy��H!\أ0����s.卌JK5NF�W��R5���C���k^��Rp[��V_-�r��K3�BO�.F��e�W\Ї��}wlfjN��pm-���ܳՅ�{��a�H��vr�������NF4ѶW5/#�WJ���ܖ+��U��������z���
�$���Iƙ��DHw!�.�f9� ��tp�S*Ez�dH�J��(��%�q �uV�z� RQQWs9w"�0�!.]�\��iEER�(���:�ShMd䓆L�r���2�'2�\܎Tr�L�EҸS13�7i(ҹ�id��಻rJ�P,���Ud]&SEL�PdG4)9effFIDT;�yTET^��:�Z	r�Ȼ9�4��GX��ki��AW�]hfl(�.Y�,� �d��WZNI:���a�S,&�9܍N%Պ�BB@�i�r�IRkY&�Z�p�bP�;�蜪
(�5E�UU2ғ����,�M39AA�R+�H��͒BW*�#�\��D�H �ݲ/�Λ����A�EY��HJ�)w9s��=�z��=k�޾�9���7y�t�_SN��*���C�ّ���_W�U}���{�)�F�~�Ͷ �l����U��*�U[>��/�Vt����Y�o{�ۙ����5����Bg�EF��#j"Ԃ]hʆOj��M���X���>U}�z4��E�S�1�c�t����e�PԶ�Խ6,�G�;�ݨL/�n��:4^&d�f<�/jL�RjW�9Z��	�Vj��.�4��#g�u/v�LY�?!��,�~Σ�rכ�˨�c��/�O	������Rxl�}�zW=�=;�䟡��nOm��Բ��K�I��IY�gn��պ���33;����㳾��t�{>�����iu�o݇t�-M���3\)�����Z�U��l�CCk�&�[{*�.�7T2y��͎�p�>ƾ6��jv{&�gV]�4�(��4��I+���kϞ�Bw��7��;ۆM�=���W�+G�}lyfu�R���	Դ3L�3��Q��Y�[kg̬T'�A�ltOUsA�vYJ�G�x��R��h��.�v�7
�Ț��B���i��P�N*wb;}��s��0y׏=����O�1�[��I!��e;gQ)Tyc��j�+����β��]�"�[�p9�l�����]�I��E��Zsu���F�����e���O��\*v�S��k�$՞�O=*������5Ԟ ���jZV������ט�Q�Њ�-�j-�f��BU2�7*�|��Y�5v��w���E�s{�_����Wi���K�+����[KO��y�܃l��wP�l��������&ź�CP�ke��OA�ۙh���!�����ST��yXFϱjlP��Z�g�Xu���=[C�Vj�BN�&�6=U�N�j��S�F�C����duhS�-�7e�Z�o��A�sU|�A剩WT�Z�z�-n�֭�Tc�;[�Cۏ<��30w��6=���t~)bߗR���3�[^�4�u���k�WqhrU�y��{�bw���p�T5�g<����uS>(�����1x��)�c��W�b�@�ڡ�>OT0�Mzwd�ɘN���W['uϠR�Ű6b� n�Nɭ�f�qw�pY��:�"Eͱ�8��+�j!�0�x-�8�>i�{��
��[��Zu�=5�*�ʬK�%��h�C���ea�3V33h�{��T븁�b�K'��ʘ�]�*�&��]��t��].ً��S{��or�	�H�yֽ��֡�74�l*S�+q*��kc���j�f�p�תͺt['�'��{�w�mQ�Dzx�ϱT���{�^͈�+�y���m�a���qΨU5��z����L�#���t3^��V���i��`�ec<�]�I���t�{)�:���VL�O8֓<7��6��8�Exwγ���L�c��=k��)҄�!>�Qm��V����W�N�[�PO-��b����1�*S����J��i'GdP[N�dM1K&e��5��z<o�}��D9�}��ڿ+{]ɶT�f�}-Yl5�b�kJ�C�J�V��������>��nrF��S���S�Za��6�j��"��l���ّ���W^F����ZM����TZv��lP�(GT�P�X;��3���[5�m!W�޽��]6���W��I���
���P�U�{�gLXn��ݠ�p"�w�������|����v��0c���^��ع�S@�W��o�ee�4�����ћi��	��+vBKS�NUk��2�c���C�"��L:o[Oj�OM�Eդw�n�W�v:�f�u�5��5�A\�QדI�w�������xD��Ȥ����O���{�Lro����}�����]H����v�&`<�p�Sa֕��Z���{�T�l7�'Q�Oj��^ԙ[A�%�%��F�Q/S^�m|g��ї�C+�x�U0ؐh�,�m�~���B��F����imlG�5lZjz�gj�G5j��ۅt.=�B����uibwR6L�D��7'MNʢ�$�ǩ6m�4֘�ni�m�[)V�V�1�5��v�]ȫ��fE�U\�qQ��N4�s�(�;��P��܊d;Q��)�-z>�������|�$�dU�x�&v�<i�r��Av���^t�iV��ל�6��2�ӭ�9c<kI�[�0̯t�'���ܯ2�ʸ܇[�>Օ������n{6��׸�L^�Z��\1_��r�.{J�Ы�2�mt-��y����v]o���<:!]ƪ�+%�-W���2�-RWu���牏�i^lRrN3+�x�UC�~��x���*v�Y�_�a�y<�Y���)��1Ȫ���݊�����s�wm���>�����l���3:i�`{-�����N��)v�gf������m�jx�=;��r��}�C6�ݜm�M��ŝ3�)Lȍ�y�j���Ka�+��
�*��2�^�M���
�tg���N����5~��j���h,�}��>�8���˞��
�~!|�i���ϫ�}��է:�s��(tZ���b�s
����H)�R��6)mt��cJ\�62��ҋ�>�������,�"�47���X�]Z�. �Vs�K��P��	V�e��ToH���r����"Tn+�ݚ1&���u�!F���Ցj�+��&�$v�䶁u/�dU��	����w���,[K�ci�
����տG�CR�)L������b�p+�0�2�^��~[������o�.���WӨb�Ѻ�P���v���S[4]=�,=���V�w��Θ=[+�����R�c�z�\ȡ���:t��މ[�=OR��$ϲ�F��d�C%�5;ml�I��+507�g*׹��÷����Y[O�����^k�ZY���XڷYl��C�guꝋoJ|����*F���5N��ѷ��$��N�	C{<����H��5ۦ��wS��K�}2$�giq#G���[y*�ǥ������{��⟪������޽V0�ͅx4����v�eh;�N�OLv6�%��H#�x���4��!ӏ�{��k�U�]4n�d�[��fI�t�m4F%u`o7r�ޑ)&q��xz�f���Gt?=�k�5��5�߽������Z1ʤ�VOq�kF6Rgר��h��a�v�y�<�yڡg3״ǻ:�Ƚ'���������)�Ě��4��Ԧ�9^O&��wf�c�����f�_2�i�ѯ�%�c�E�n|�)�*��蒾���>���e�����읈��T/�a`��M��>�[<q�!�r�OZy��^ݓV�
����ϧ��㷘�hd��O��b-*gh�E��2͠1��o#Y�h�O n=���~X͗a�K�m�V6Y��'�*��.�jDѱu4�U6���LľL���)�E�P/Z�"60��I��$��*ޛ�5�Ij��m�������*���}]sS)�Ɲ�-
��L�U���m�lD�� b��^fG����9O����������f�;����38mGܞ���J)-��fVd08�nM#�:��D���6ac	ٙU�ȸ�ɍ�����[3i�%��-��]^�j�����AT��2�Py�m9���KR�r�����T���ڬtMC7�x���_��+�|�����I���-]K�O�B�V-��ǑO�}^�B�|����f�T��e�m�,~$���0�;<�↣���A�gԽ++���w�f�q-�|���\9Ա���c�>e�8څJ�H�
T��-~ܩӆ�o��O.���iz�<�j��=Q/M�s�Q���3�3��y�+T35�c)f��S�LM�hwh����u9�Un渠�Ս
N���je;-9�'uK\n�^�Ǘz2�wtK�v{i�����_g��k�u�_W7U���)j�<���S�\}�cn�[��������ӄ�6y�OJYw	�!>[�v���S9�k}ɑ;�`μ	�)�b���S���e3^�n�X͐�(���!�(-�״d��R���v���u��u>eh��t%d��S3ik��^�9��/+��w�h=��U4:m�S���ܺ8Qv�U7R̙����|Q �����A�jOv�Ԡ�1�ú��`���j]�.�^��/���@�1E��r��{��bb�w��fl���Ϻ���˾�UL�z��-eB�wS)f�3�KQZ�a��fk���σ�uE�S���S4���]�{A;e>@զ6BU�{�h̸q������&p�Jo�9�{^��lN^N��T��~���O��뻧5�(��w���
>����n+��\��ߍRLe.V2�'�����<f��
.�ҭZ"5�UCM��6�W��a�7m˽�ɪ�5]p֬3�Ϗ�]�����~���^պ��ֆ��j}1�1jA�I�Хf�b�5�M������^p/R���r�ά��ꏇ�y��U�#<C>�oH׎'g��ݬ�Tu����������KԼ�EU>�S�ó��{H�'mD�^�O��g��5����Բ�k͢�uNaMZc��a�n���Ć��lj�Kt�ޱ��k6��z��� ��z�W_D���;�����B�>��.[�l���pʂ�b�׽G�T2��u�kF8w{D�P�*���ǡP�����>�T1���I�>U�z\'&�n�t]��p�E���]��?ue��sL����5���N]LuN��@�ί����:E�(��*;�I�g��ҳ��?�ꪪ�>Qù�&��������W��?y�v��r*��L������p��-w�6CBP��[胇g3�d�b��ߦƠ7���W����ȩ�ڬ7��ݹK6��-�|k"�
l������z��4ߵBS�wf�n����)ބ4��՞���V#�c5����
w�K��im2i,�4Ǚ'Ҍ�0i;�mYJ��<վY�]N^�&-���&���K���Z�:�+{:��hk8;;|������5u��Wv�O�[K7�Dߡ5ڟ����>3вI;	�Z�F�>��%'���LΝ�6۰�b�k����/:���6sE�g�����Z���G��,)��,��joe�K��2��Se(N�H��J���r��no��=Ysm�~T�i���J|6ے���;£me%�u�ujo�u�T�ŝ��:��U��[��5��Z���j"ԂL����2����߻���fzs������S���Ypu�un��P�o>J��ZVf��һ�c]�hOc7f�+姒t1tJ�UЋFعp���N��X[�8�W�S��s��ڥw���=��Ym��j!�%9\��:�Nȡ��.]�~�ﾯ����r��Y��T��٪z�TkZ�J���?>~�^�xpg�T��=��?Vr���yX�AE�v0v�����%�|��,�B����n��{���w^��A���s���O ��YP�z�,x���Իi�"T3��U�W�=�G޵��r�׻jYl�ܡ�T7a(V6��O����kd́t�r;em啢e�_sҼ�fŚc�v��kuH��>�8�}~
���Ϛ�zZ��<�q�OJ����r��F�wYB��,���yRh�y�!64-kh׼�y߻�R���^=����#������O���{��za5���_�ѡ��kwǖ�\�#r������~ɉ��_�w2nv1fG�mjP��R�EHG�t����r5t^a�۲�bDNx���c�5)�wxwI���O_��GYlzT��}9!�6��S�U,��.�m1���iM�Q�U΃t�L�X�-�u��΋��^\��v���*�6�0*+%�s�\W�����P���� %���z���ƩyGi`V�A�f��c%up�@�==0Iuj^+/����㍷չ��w�q\�F�O�p�܉̚S;[��G(k8n��Yf.Eka�P
g�֑E���˾ٗ�Ջ��\�2M��'��X&�4��4�v$��;�{ [Cn���a։Ս�ŗZ�V���K����l��V�� ��]6��"�5��+���I��Ϝ�Պ��nЬ��H�9Y<�j�><â�RKdm_�v��#���v�ݶ�Iuܔ��6 ��Ƕ�&�����_iu��Q.��4XO��SD��.�%�`�7��Z��q^�����1d���Eeo��y�^c��EWu�i:����kM�Qr8����g-2	�w���7��I�'l\��ŬƲ�V�5��)�g8o:���{IS:;C�"���b�����r�r��f;�׷���VN��s�b��6��[�)�c�ۙ�'�&�=Q
�Ј���:�Ϋ[hj�Q�C��x�J�fW*�GJ�Kd����U�z������M7�mW2�X�C@_>�6B�'']�X[��IT�����3pɻyK�MeE�&#�4,�h!:!�
�,[$lq=leh6��uF�;Ϻo���mtke�7Wyjt�m��
���a���_&�j4��v�U��v�gv\Zws�ת��46��/5=\�V�K9wx���ˑ�:�4_&K���}l�e+�z����q������X�ts���&,sbn9�����v�-�u�m>����+�`z�[y%�éUг�ҫݸ�aR��4�vl�,`��-�]|�>{��Z�0�f'u'��,f�6%����ʓ��A��,=�wl഍�j'|����H�v����o嵩�C*jAG�(�W��e�)��R#{U�>��0���&s��p�1��rR���+	��%r���+޺S[�z�:�B�-�Z�?��^�k{�e�蝅
'w/�ZE7z&
n>=���uڲ��s��)N&�M�]�ט9�w�yyMQ;�#A[�qe`�fJ����&��w�G)Hp�����#�/��n��Q���t���,u�ݽ�\oN/C�GS�O�J��jt	�"�o\�Ӵ��[�#��ޭtZ�9�N�cAp��M��8�qv�4��[X�u��IIX -�:
TL�|��y(6�sr��Wz)�m��1�3m��ִe��e[)����v�T��y+�T��k����Ν���M6�嚅�I!h�vi�f��EQF�}z��-��e���Iou[W�L�F��f�lT!�z�}\@�ŁJ�uԞ�X\�`{m?��=��s�}���.G�;*��i��B�D*�t$���H�*�7�B�i�҅"eUTAp5
$A�K�eV.y�Ju�S���EDZ��E�U�� ȭ(�5P�e�$.Iń�	0�%4����""r�+��FsB��Β\�,�J*Z!EA�7:�]<�ȣ�TQ%D&�Y2��Q�Um��#��Q���
�JE
�v�&d����TVr+[��Ad�w,���%- �P��瓸$UV��Ԣ�$죕TVetVFE�sS� �F�Y!�P�ukH)+��UJ�gs���T\���"*'%����NUbH�����k�rRiD�**�:$�J���Q��Ԫ(��֑�3��r��E�T���B�q�\v�QD\%hV�!C]bD\������ii�IE�YI�Ȫ�B��A��L�e�U�d�Y�fNaDU��N�u"dD�i�P!	qX�Bg�g\�*�*
�������ޟW���?:��qe=��3]Z��w��Aݕ������*�wU�`��yH�r���C۰��%7:�f��n7�������U}ܜ�/��հƟP��M�*C<j�Yi��~Zv���V��ɧ�L��,ی:l�w,� �)�&��M�KTl"��W��c�(�]����.�wLV�D��Rx��lq����Sb+m^590ρ�w=��{�Py�{w]���r�T����#pM����xثh�y��Z�����fo���++�����K�|��3��{�z&���md��F����Ϙ��ŏ�s��a�������V�(*����6'��Җ\�HvL�5��l��/Ozi�����e�v�ʯ-~N��Y.�8�踷=�V�3��/;���ӷ�jw����m�rW�%q�2o
�+���U����4���9��2�4ϝR�6*�Y#-�b�
Ȇ�1�z{�St=�bVϫ�}p�yVW.9�sa��V7k_}�7.���\`ܙ�:�e�*�mEֻA�׆3[�g�=�&���stQo��Ί�3YX'�V�"�WdL �\������a��$���@�s-i�+Y��0��e�}g�M[TiI��l�ޕ�4���[��oR0����G��sp������W�Cf����)M��:��+�����&v�Gw��{�E�vZ����ù���7�O)����Q�F�kk��ܔ�^uro��ݼ�|�Vy1)�7`&�u��rj>R�R���w��!]��rg�o�8�l��\ǹ�y�Y����=O��MX�ev�P��XСT��4���[y���,����-t�6=GC^�ГB��0���w�ik*{��=*Cƾ���r����d��-C��R���tf��;D��UM�Mh'��xե��	���z����#p��̞]_��d�L����{j�����Jڇ*��@��N˯b�"�(�b�nô�c��(g��"a��zh�/k~4���cx;ܣ�̏Skh5�1Z�����K�m�b���U47�F��1ۖ7�f�K5W[�*$�}މ��*n�����sl{��+�v���䊍OF<��=jA���*<��l�#k�y��/^��#�<�gʅ��ҕ�pY���y3��l���D]�����sr�e�����hX��l����z>m	�<��uo%���E�:B�]#Q�W)p)���
)O�^�Q�G�hvx�|n��}��w�/� Tm���ʶ�D��q���u��\�
c�<ɔgj��ҝ�U�V��ћ�W��%�A��c_�G�{R���R���,��Zrꨨ�!����ɞ��?B'�9�d|�񤦯Q��N3^�l�GuV��s�v�	8QL��\�U�}�س��5�J��:�rךB���x}y���뀤Ly���ܮ�gT������J�e���j�ci����ǈ]��Ŏ�ީ�iCJ������o�^>Ƭ׌�d�,V�q��t��3�)٭�gU�rlEﺄ9����3+��Ξ}����wa���W=��x���~�����{�@���Ŋ�ik��;�ڝ&�Yt�oT$�'w(��@�SH�2r�e��L�^��ǋ~�q��'��>�[�C��=�����7�/��'g�f�Q�[bN<�H���m��^���|��ek�W�q�̆S��e���9Ɵ�7Xip:T�s��W<C���#Ң9ȞP8�-nϨ�\�=�b���5F��F=��ݍ�9;����Ed��gyl|ڝٹvUŚ�;��>���(lTN������n�A8�dL)h;C9�*y]u7Y���oz�=��y"��*�l��EC����&@�V��(�k�pŁx#�ZGD�`Hα9-cVmJ�q�FOn�����fl�X��}��4~bz�s>g[����Q�O�`��>��iM��>���RQ���ј��Pu���ޓ�N�Y�ώy��� Oāo����{
��3�z�q袄�6T�5��v�9�����s�O��E_����㡗�����+�=� È�'����ǎ�B�2/vcl��q��|�T]����,3���\!�=�1�5ܢ2߬��q\s�\H��έ��Aǃ6�Zr0�������g�sf�*ou�ǿ	�o��+����&x�m�A��*z��ې-v��x�e�=W+���!��tAfTd8�뜦�z7�(���Vڀ#��Q���Ʌ8������a��0.5��d�\�2��3t�{M T2��14�|�h�Ns�y6������"n�>�M�q�N�ԿZz��m��,�씏==����+�F Usl�;�FJz�d�W��Pz��Oa!^{#��jղ�ף`#�d�Z�K^�!�[a��;
i~j#v�s�m�F�fI�k�0$�G�߆�dHH�0'����;�*tp�z
[%��=�TT�Sֽ��h�\�76��oK��P^�N1�.x��v0�Z2�YQX+obҸ&�`h�S�����U0-ͬʓҵ���9K�F��7n�̃;��Z�K���mwvf���L���f�oJ-H���ǹi��Zە�r��}K��;�����FF��B��L�������}�-l!WT�5O��z��Zk%�)�S�ir�����9Y���sw���{D:�w����|'�hׁx�e��B��Y-}��e;Ѻv�W&K2dR��4yƋVJ����a�h{��R�7=G9U�.FZݟQ��t@��$M�(�yf�Xb�G,mm�q�;2p�@��j�ؼ<Oa:u�D��"Y;�&�r5��s$d3Otءx�U�j�y��]�x�h�z4�0:{20t��ƻK1O�#�)�1�����u�[��G`�vz�B%�vs!�Q��y�L�(sjۗ�ZU��
�~'�m�i�~���� �a��R�WBa�g���T�}�c����rW�v��k��s�]a��k�������0a�8�����C��S[}UI�4CQ@n�&Z6:Aq�uꡖz�9���%?�׿�?	U��h��\��qj)�0uX�@<��lD�ݨp���J�O��%��«{�y��Ĺ�Y@9b�R���}?c�ՙ�/պ��X���5�E����P\�ptVy�2z�������3��:�����{t�WNx���88�:gC� �;ث���m�Е���"(aw}Z`���r9��a칲��<��k����qw�뒐ʊ�g� Es���G���ᝍ��7�)N}��:$y9p���v�p��\0X��:�g ��a=�%ϼ��l��$������
�l�§��۫�M�P�u'J]�wM���{Jd�5�z#"�v[*����Ѵ�P�Ztm�����r:�! �Lpy���*�E��8ZY]��1���)����(r�k��Nn�䉗�aG����h�s��r!s�!��Y?Y���4K���\�f�ꛯg`!h�l�0�{�,qV������t_Q��~ƽ��)�#�Ϩ�V-;SU��"6�E��݇�B\J��ࣽ��O�^�{�L��S֧�Q\w�.ڛ��*û��O=]Q{�/�H�7Ef�|2ҝfǸ:gծj��)�b�c�`J�c���Z�L�xz�̚�c۴q�]���-շ�(�wOKtW��9B}nΑ�|�Tt����?�_F�:IޚI���������j~Ge�#�w�8'ͼ�u�[��=*���GeL,?"�U�ZטŒ����0e�/����SB��i�b�n>aB[c#��sT�
Z�鈫���H�v�d����z�̨���//g�w�`by�p5j��R��-7�>�s/��_��/��'�||�-��&�}&�oן���V���h���f�T��],�z�����R*Փ�6��:~փ��߲V�X�����zB�7^󱪷�O˭�3+�F����I#�E��NV� ;��4��C��h���{\7�S��k��+�c3i��i�y��d��n��|�f�x�N��G� Ͼ�!T�������r�� t��sZU��D�0�ra����j#���Ȳ;%�����jW W;)�#ܦ9��(tO��1踱�j��[�e�r��Α�e�b�����@v�$�7�3�0آ8up���2W�����a����c��h������)x�g>�1��6'�^=q�?�!Kp�f�R�}����\�-�̆�Πb��Cn��'��s��ۚ5�	�m�=��]�Y��~�vׄ@��qӞ����E\��}�(���S9���Oy��g���X��f���!�]�Ҧ�����dc��Q���.�(�S���J���B�;DI��̝�8nz#E�zh����)���8�SF}��.[: ��mc"�wQ}[F3��O+/�ɋ�7u���Nt�S����,X;Q�`+S-N�����S��.���uU�\Dݢ7Z,'�}�Q"+�u:�m%q]�ݍ���dL5�l��
��)�܊�q
�ތ��aU�n�J�y	NB)'�:��J+e�i�(�w3�N���gLK�\5]�4sA��u�Ws
���)p��czc�3޼QM�mfrt��@[�K�r5;Pc�})u�ǚyV�f�����yV,�7�ֳ_��,ξK��7걚��o7�X8Z�����J^k�ڑ0պ���	ղyV���+*�]����=����k��!�٘�f/JVj�4b\�@~6�e%��8���#��y����٪9�����-�Y����ڈa�7]	C�u[Ƙ���Q���N�j�h�#!d�,�N���?�����O��dC!��5�m���ŇZ�r	�p���.9<���ŏ^�x,��T+��׸��e�s!���#+V�@חUH�C]e�����t���U8���	dg�#���#sd�E	�`{MQ����PLE�	��L�uQ���O4s>Dq��9�] ot�*#������~;���b,:4��ɂ�3��y��-|�s��Ct6?F�K1��-��å�T��a��{L{��[,fƱ.��&����&��T�ױ�b��Q-��mx%���e�o>3l<�
倍�+��ݷU¦2"e�.qimB�ӼCmq��-�w�8�/�p���혇DJ~'�;���k�ˈ�rݽ���6�c��ւ"j�G)����\����6|l� {c���q%�;��헎�Y����v���먷3�qBw�C�k�ۢ��d̲�3~T���Ǫ��/�k�#��.T�ˇ�CV�@�ݶ��1!��w��5x��1
�2�Q���+�]���t#cMe�rN*�4�笪(�Ow���K����w١a�9��n9Xw���qKK9������PK&�Ԧ�;Ө�g
TWI���������z�v����^h�f�R�q�n���y�;����
�u�� ����.ZY�S����`ԡ��o�՘�O5�D�aq�=���]o;�R�i�������Th�қ�����GHp�`��~�:�J�Z��o'0��Fk��w�*���d�#��Z�>yLj:�;-y�W����_V����K�ZW� vY���!TuN�P�M�!"��E�c�7	��������,p��)��Vp3I�R��?5�2��[��+ϲ����@���e���Zk%�,O�u�?ų�\��DckK��n�4]��=�n���\�^��'�s�c��m���KS��y�d��.Y_!N�p�>?MDn�VN���JQ�mw�)ncA�:T�\�	�X $vݟQ��t@���@�:E�u�X�=ˡ�|���t�Rq�KWT�"T"tO��fݟ�h�"�+K*9eL-�s���;�gaY�`x(�d`㯐��i���O�)f�0��)�"b`I��y�;7Gc&��-���(w������~���V�'��i�<�y�a���`/צ1���d(��O�e��֟a����Ο��о�%�z�T�Jۊ,	��X%��7!�`1�-�XV�1�Y�o��4�+K�Ձ+j�\L-����z�84�Zx�y��q�b��$R��l�Q�]�f��]�;NVb�����;53P�}J��ڜg[-��]�z:v���}���9�*��wO��G���U�ˤ���W��-c��I��fUy�&�J�x��g�=���ܓO�: =����;���t�N�	<^�s��������x�@�%=T2�]G9����\2��0�ja;��
�Z�M�������T�>�n�������@��FG����ŏ����1���|/�lC�aͱ��-|�z@��|�6�g׺�D-�#��<���a�m|���=߱v�U��
�k'4	P�3Zq|��:�aK���k5�}?b�ܶ���W~C#�/����C��ʋ�I�h�x���<)��$�Zp-c�Վ���S���Gi������ˣ��8I�ުڥ�^�pvF^�=�c��m�f��M��W8��B���V�>Sg��(�z��J�,ff�����@�<ڙ�l�A���i�g�k��������;��5��)�(�U7�]���H�Q�{�r�z�el���]l��r��fH�] ��_@��UL(Χ�.��uUΪ�j�܌؃i*��0o5o3.��>��w3.~�*+��{^���֠&[�@+ѳ���d����!�A�ݺ�����J����+��]z����Dq��kYԠ�@i�:hz�v9�Z&��ᔡ��ֺn6.;��-�}0�+����-0���ǫ$Dv㰣%@Y�R�6+�NV�Q��dK�iJ�ǫ�x�(�+rJN�
z��Q��:�b��=y��Y|��vlꩭ�2\�\�T.�ҧ+���Ǫ$�>��j
y�{�i����a[�{�;>YNu�%ZX��8N�����$|��A�֕�f�wN�M��P"l��a7�[oP��D<�b�����]�;a
���#�����������#ڳ*Q#\��
���Ӥ]�+���w]A��i�g�M�y]'B��z��w�4��ϦͻyW��W�E�Z�O}1��tP[���ka�I�PX�KVr+���å!�u�`����w��}���̼���6!.�[�*)��>wg����JS�8� ���F�`�4�<�q�3��ռցï��c���-zC,���x�'p�>���S2s�V�Î�÷ ��:ԏ�!�;��]��/qB�@���U=��V���u*M�/�U��e�sU���X:�݃����|��ӫĊ���7H�ˈm�>�;uٽM5�����+�7(�\�԰��B�qM˕�����mV�B�����EG�Z;�G0�8��]1��m��	�W'1�Ri�� /e�ǰ\��3(�i=@#)���ӛ���A赖��+�m`���T�mAM������ӕ��N�]���Y�ܭܬ����r�8
F��4ݛ��\���dF��$Nmm�Hj˷��0�Ƕ�e�-%ҕ�v���b��6�����ѻ˹�����U�Q�I�&rՁ%ef��x��=f�:hT�t\����\̖l�7Q;Z��^���v� hu�#�`��5���R: :�^c��]gN��Ge1�%>eWF�I_gY��aE9��(�fQRa���{ˬ����6VYv�e�������1�p��b:���5�%@-��.B�b+��}B7�*K�j^�N=�w�}qp�y}���j6W7�N��6����lw��=RqZ��j34���vt;�5V	���.�)ң��ua��əAhT�VJ�ױcp�LA�tw 搼�{k)�p��a��_���2c�Vܛ���ǖn��r�+:�4��gj�j���̝J��e�NbMe��Ս����CWϖ�u�q��vW_R�ͳYn^f�lv�F5ڭ�t_b�PQw��3��W�Q�s�$ثU�;oSk������ysN]�ѯ�O/8����1�F�� o��ѭ�>�7��Ywx��5[�y���^|����Cf�6V�z%��#ڪ+�׮�By�g&t��Y�z���+L��1�L
��q�7����ǜ�r���\�a�?&�5���L�]=�Ʈ�iV�]��;���c��#[��ܦ���O.���Եm[a�h�]��+�����oj��jIY���h��o
�}tl�u�ݐ���w
P���$�(�U]9F*%QVE	V��TW.D&t��IUr���DEk�"D]$�Ϊ~t��"<��PC��4�8W )L�EGR�N����!���%t6AD��DQEU\�9TQr
��\&uA3�Q\���9W"���"�D�*��P������S�쪊.HNq$�L�-���D9T�
�*��^�B�DDEE��Au�s�p��9Ar"*�)"0�����2�w\Bf���)����9D�ɧKR���IcH�J:(���Ev*\�AE�EEUȈ�ar�\"C�\��p�rE��*�JX�QQ���G+�9�U�t�Eʊ��*�v\�(�SL��Qr��\���Uf]NTQ�@�Y����r�Ñq;H�DDEDʢ����g8z�GB@��TEy,(��=����J,�59Q��H��h��%��N�EY&asR#R�58�QE)�ЕKQ1<�2Ga]F�;9��	�;�jw�*h��(������!�n��츪q����F��� 5/��3�sԗ���f�6:����:=����!a�N,�wOKu39ڞ���)�tl�ݰ3i���B+2�NuS��X�e�hW�tpz<��d`R�������VH�i�T�'���YHȮ(]T�ܳwt�{��wd)Ӆ�oP�>�Mi�b�,������<�N��/���Z����]fl������[bXG�l�O^$�y�gl�4Һz .5X��Q���#Ͷ�:�q�V1�j9� f��n�H�����,�� B��%�`#����o���j���*�a�UM<�m�gT�!�5��9���eY o���@�c�����]�g�u��/�x���ݹ���_[վ}9�Dl��%ߙ��Iò�O;g�3�0آ8u0W G���Eķ����|���e�f��o�xfi��a&:��46�f���\ �-�[\(aW��bFEŭ��_ �D�;}�4�fmf�FM���K+��]�Y�O�[! ��(�-��ۧ=���z4���Ω鿹;J��'y�V�V�����0���~ɵ�:��5���Ӂ}9 ��(�S���S��vz4!�V5������7Q9F�D��\�9�(ʁt6���:�xUR:�3>6�hfu���;�.#N�C���Fᙀ�3������G{FA�?�9HmÜ-l�w�Xmv�Z��� ������l��;ս&�.Xo���R��A���2�B@�g��3�v{���广��l���7���(��}�B��e��<�F����<����ɷNZY�L>��3�K������m�S���ްƚ�;����4:�{�e
�:g�����ŋj:lje��N���Pn��z�t�fi�΁	v)���>�Rw�(�����+�!q�y���t�`nݟ��s�"�����(OMft��jw�=X����(ZO�v�����)����*�h�;:/Kws��'��-�6nn��/z��� O��x�ӤvZ�G#�_F�'�9|�3.���ԌOB�:�����n�n��r髛��זN�eF��RIZ_��ڸ�P������&̥ �ݙx	sN�P�5��8�鹱L��7M	<۸	c�G<�>uU
�2��*�ĭU���;:��<��}�}4{�y��pZ��$D���K7(P�v}G)�����@����cg`��WuQ�;u�.�\�͋��[c&`ς����t9�z\��F9�3��d�][Ǐ\��Ԯ������{m�S��`C(���a�o>{a��K�=�c��/���z�r��Q�ϐ���y�I����=�`��OVȵ'�8k�[��e���c��R����Xi��7�٧u����ͻa���c7\�b[�����毘�������SY{i�݁�z`�aӋ����u�Zw�g0�[��0��c�[#�Ƽ�{\t2�py�=��u��ْC>N)Q�c{#v����ݐ>W�a���]��f���8�x�C�7�f8Kk�DC2��=3ݹ�27����t۫w�G��6}�^��׽��?~�k�
��kɽ�2����tp;�-�<��5Ә�UGUY�
pB5�ꋃ=�"��p�
�2��-�9M�����(�zvEhy��Z�n�%TH�a\�`�򈔣�#]�"{,N	޸q�k�=�h���\N�Ҟ�'l$�B��@MZ�g�aۚ����aq�9���]o;�e/֟�*���N#Mf�H�t��*���]ph��ٵ�����z:�
&��S�i�$+̎!�l �5����W'Kj}Y�z��9��O;:s�d���ne~�t��U
�
'Q�P�M�!#8�Dz�!i�iP�]x4�W��LF�L��&�:z����[�H���@Y>}���� MS�4JN�,أt��SS��KM%��*�m���O}pk�j�>螞��V\$����Q��!U0�S��y�;%�w���<�g�ī7N[u�TG⩸���[��$��=���X�^㓻�r�ғDܚû�x���x�_��٭:DE#wf��i�Μ�2T��_>������c�_Ϫf������w/�ޅ�q��.a�q
��/wn�<L\�|��q�^�,C�mkn�`}�����=ǲ��4��C��9TJ����nk}8]8�*���n��{��s������m�=�a�=��Rq�WLr����u���,�J��([B1N�1O��3$���V��	�=f�;1�v3�ƻK�q�%S]KTJx� -����?E�`�X�KSSt���gљ^��,CMm���j��AЭ��<(:y��ϲ��9���"��Պ�W�n�,�y��Cg�^Y�!�_<Y-��Qnbʳ�,�X���F�4���M��S�T�o�Lp]�#Ǯ �Jz\;�w���[rʚ�9�5�d��.=�e�;��*WG˿b�e�À��߽������tE�B^�X��qX]��^=��Uoqn=��bc�+]M�.]���5�kK�'̳���_DXyf>l��9f������r����׎�ӳM9̚��V�'�g��->�eSz9�_�a.z�vY>�4[z�嘐�z n�Nn����`��8��QJ��8:��L�8����@�j���;
��.�m�����~ց˱l�Z��ՉL��՘� ���9�I�7o/���ݳ��騶C\�-bR��v��=ykE��Nl�i��-C4��:�*��f���s�w9N�\6s�t2�y�v�7�E��p����nl5}+�Y{�{����Gb�)�f�Z�3c���w�lB��j��P����N��k�S����Z�|�E���*F�4���ޛ3�ݗ(!M�>����v�;^~��!Z�h�ujw�k�N� �z�L�egfte�կ�w-T��[�vlVu�Gkݐ$] ��^���T�i�S�p�W��Z�;���i�ې���d�1V٠�홥д��t���FĢ�8
s� �4l���f�Ng.#π��dݭ�Q6��lz����;��6lf�5�B�h�9���n��
�gH�Bl��� oHՕP�Ua���NsB�>�F���������߰��χ_Q_��]M���a=��O{�OXh�_3A��`�S�8����4)���wa����(K3��2Ǟ��
�[v��e�x�6U���]t�J~0�&~ҭ��z�gk�i�t�kĮ7lYI�g�o��ƻq{�f��j�KrUl���͏с:/��nPuK�M�P��#x�C����\�iV{	���݇�~�ξ.����=��=�6�e�z �`� <����l:	w�j�rpwp�oi��O8G*l����vXV�3:*ҨZ�\Pŕ�ЋB�&5��ɣ��Ke+����j��y�[X.�e)}\뺖X澻UgQ9p�_.VvT��Eh�C��������p�%�Y$/�9��oVL�ݧ����0���͛��;���r����魜�E�ܿ[���,�������s�й��3ìv@��(��w�4:8��k��ʞJ�k�oc�m�:w�gy�2�׭�v〾\ �-�}�0�2����^y\�g)�>��y�"�T�f��y����w�&���evW�ó�+<�Z�r~ CgTp���)H]n��M��tH���,7����@-��k���k�����N�? *�[�_D�����Gl�We�=��nQB�ϻ,F	fJ���n������u�t�ZY�`��?�{�<q3֯0ڗ@�d��vl^Y?F{���F�]�	.x�`��E��l�R w��b��4L��/k;Y9������"4���4��Q;-}��o���E<�	�u��y3��n����~��*��`|ڣ�"i��Z�֞�ǐ��!"�|�����S��4�[1-�ϒ�e6��7�4��QN_4l��
��O�^i�;-W9Z�-�y} Z�����4ffz��l։;�2{��!��9>s��즍�'!T�RV��S�[>��(K��}S�P�/|��!g��YнὉK����/F����Wn�FϤ7��.wy�@v��;w�(\�Es9lL� �trݗ{x~E�y]�ڐ*a0Uwn�tA޺��0�hZn@]a�ugoAMp]�7`���2�(�7�+w�]�Ժn���$o��7v��0���ˤ���R�WG<��k.ykw�����E���Y3ܱ�c�~*��Z�P��5��]nE����95A6T��Q	ȞP8�e��oNEGtP�g=͊nMʃsy�Q�bv�n�26��J�ˮ�7�`����r%�`�y�7�w�P��*���w�k�ӡ�6�.�A<*���)���hf9�>t�ܦ9��W���pMU�A��[[����72�&��b���������gO�뎆����;�f���<m��Yٲ��n�j<��n�=��k�DL�X��,��;�'�^��1�[6 �y�[V�9n~��9�S�o� �̵���>�����^a}��\��`�����5��Rhi�����k�j�����dK,���T[��w\Pސ܌���2T��r�����C[NIhy~x�Aw dt ���(\2͐!��"�)��lLP�n�Ҫ��\`�~������ڟ�q�rh���\]sm�s6��v��qi��x����p��'��rtʷ�R �s����9�G�n����0��}kb�	:{i������}{�Zn�]���*��#X���Ss������n���:.���1+2j����z�qɃt�w^�
�p)�X��$Z��E�M1��JF���N��q/�8���v�4��hv;��g.�
���掐.=�F�S��4��Uc�Y-��F��A���d���qF�ۣLZ���==q�����c��l\fx�9�)�:tN���w�f��ެ�	F���q1-��YO+"7m�Qq�G\T��������h�e�:e3쵰��-��Q�PZw%�*y4�G�=bk�/k_y�F�i�];{c�����_b��������j{����	����fxc�C'l��f�uv�z��U��n����5��4��B)�#�V	kv|G)�: \�M<�-Δ<�K֭��̟��V?;�=xVz��M�Ü{	�4�=Vf(K't�D���G#M�\i�nO)�����[��}�/�=�b���F�:3#K�ƻx��$��MuK�S�݆�.;��^>nV����r崳��ʗm�`r��3*���	
�~'��}6y��˪�m���vm<rJ5�i���κ`!����	mg�0�2�ی�d�D�[�
�E�1�@�1�vAl�3���3�7���p7�<@�4U���Ac��JE1���<�^����]a�����E�Z��N�[m�F�J����}*��x�뗃�]>�'�{Һb�F���lȲx��O?=k�y�r�k��R����7+@ �m�ݫ���#�H)�f�_jB��s���ҙ�mZ�w]s-n������[���m�V��Gy�ܞ��C���6V	�u�����O6�Ɖn���>�pe�u27"[9������'ǫ�Gd��g�so<�q�nWD�m��|~m<w���>B�����@���Z�"��u�	�~|{��-Seo2v'�H3���wu��Do`��k{f����(�R�O;{�}��Q�&A���E�λY�L��Ù�ѽ�t���f�|�6�S��[! 5C�zmQ�S=˖����[���[�f��+Fs2ʓ���>���{�v�K0��L	�{�\@�nB��B����p�"氎͜3�a�=Q�n�CE�]ƍ�r���C�Gi���je�ڋ�2���x�)l�	��T�u]�|�Y�@�n]44j;Z�tp�(�����pt����5�f�UL)e�lL�a3-U箽�Ύ��V\w'�,���f������3���L�F�8

�P���vPN8�я���V�Wl*��%,�������v�YLȊ/�=-�2�A�{���=��eq�&�xl��s��s��P�㺓 J}�O��d`D���>�#��U�N��������ye���;��*���eQ�t����ڕ3q�B�E�/�K�J��<}�
W<�@ܝI���;�������w�f�§v�O�h�x���Wuª��%ӕI�+6:]����,s8�6R��ۍ��.�{s:�v6�vE�����{�D2�a�6X�W�s�f]i�b�kc�'c#��Q��r���a�-z��
�Kv��Ќ����-n�oc�1j�U/$Ʃ0vTr_���U(����6�Uh��;�x��qП5�-�ryT����qy�/& 驂��`Dی����d��NQ�+���Pw9�<q����� G��9x�(tK�F�p/��y9ob"���ͷ-�Yw��á��!�6��v���b���� �����ϥ��	�?�7�;r���;�h�g��=Moc��s�/�GKp�p���}�x��:QM4�*l�����_�77wX3�H�5l�-�-�
v�fm?yl��� CgTp#Q�co�fBd�?Y���}_E�?m��/�q�p ϶�?=�^��!�]�Ҧ���SM{�ڥ�\��֫�|3^lU��P��6���yn	�L���tt��;�l�r�&��$�4{��u	�~v���]� ?��QyS-n�S�)�`i�����b�����$4+�/5eKem\³��y;.��{%*j19�]h7����@��բɋ1�=�#���CN7�YWP�Z���.hȺ�VvNyqnT�}\!,���e
0����@�Xt�ei�o�j:���pӜ�׬���)�P��8ݔ��U�6��	3R�Zo��gҮ�����Oĵ���T�����dN��Oq+{�49$����2�����n���w*�Θ�.g������r���ӼT���پ�Na}�F�5���\�{7���H�3XCz�P��I���H*j6;����1�)������>�l��7{b������E�������+ݎ����{����<��4��b߆w.R��؃5-CS+���(^�%�1
uuB�$A��oVڹ����!%>�ݛ�j�t;�ӻ�CE��5ր�j&^vgR�Է��/�^k#��[�R��0V؈�#�[���b�C3����w�RJ6��9Q�gRɒ���ɵ��5V*%ۦ�WH�\h��]E�YBc�SI:w�zf��q�v���.��ʘ�sm(�(����fU����?Z3=�ez���ossn��EA��w�
|�ݝW�۹�u���e�Rl����r��(�=Lg�����je�l�殰V�{&vc";�R�L��&��N#I��/�)�I��.�ѝ#7Mns�w�ǫ�Ef�O�n�	�Qs�v7�.��K�s%�}[li!P�|q�����J![���wZ�]�-��:�f����J<�R[�V-�I+�,� �o����ī:�7�g噮`�5�`M8�l�#�Q��V��1}/f�>�cn�apl<$+L�����ً���u���U����n���׷q:�F)+L*��%-�Y(V�F��E	s紕u�vRtB���+{�~\��/hv# �ŝs{)�ؤtw�!q)�x�W|�;�sJ�n����L�d�z�C����W�֯�tkN���X�+N;KU6�]7.���k�g8�CN����՗�H���vH���j�0ܖiT���W��^!+I��6�zyI�;F���w]xf,]O`,"��h�R�CL��Z�ˮ�)C��f��v]p]��ؕZU�̆]Ð�14a}p�U2�m�gD�뗝�D�4�]=7P�l��0q��{�gc[�KUR�YQV�"'w�+6�/�Ĵހ�ۛ[h�Oe�|�ǝX�4���R��3���T5�c� �3���Ug���Ν�˲ſ�L�(�w�=�����x2��@:�*트=]sWc��w�"�����`	oW�	x�]����E+F2��T�����Z�Cv���������zI<�+E0�<�G��Gv�����=!���ޤU-��X+��nď���9G��߲��+���.���m�KzA7(d�ut�=�ht`Z����`a��a\������+�$�v8�3�����%P��8}D���Y+Cn�f�d���s�tr�B�  h
>�kY�YUY�,�U�l�5K�t+e�R:DI�T�QVi���'���вQ*�҃��R��ӥk��vP'B
���E'TH*sa�W9�N#Փ��i�T˕D�TXt�R�#J�
*�UGJ���)$��Ut���.r�Q5Xs�d��΁PD�J*�QG"��J*/@ź$t�����QP^qɹR��Jʷwj,ev\���Xk�QEʢ��Bt��J�9%��Us���ETU�4��H�E\*Z���EȨ ��P9EQQNIQW.U��*�J#�܈��)�Y�M�i�*&�yG(��9^�I]$�
���QIӄG&Q�@���$�#��"(���,�(�wAQs���y Rl�$(�����\�6BaQWe�W�p�\%�r4Y\(#R��J�r&Rp�6TfQ9��*&L���K*�HYQ�-3(K�iP9\����o>�����%�GgzY]��Qn;�#��DM�@���L�"��پ��WR)ֹ�Vu���b��tm��I�ZК�#�ʬц����d�;}N��鰸J}�2#�{S���]J[+��k��'K�e��tF�ìz�m������N�P��3��S��Տ!)�BDRQ�kS�2��Yzث�A�yi��M�����2��`�w�6O�+�F́�
���/4��5<�Fulh�lO�q�t�h��h�i��7�[��W��]9M��ߨ�el�c�Qú�!Ōu��S�/4��Tf+�4����vk1Ef#��ӦѰ��$�СŲ��T�\$��wV=4s��gΪ�-z�d�u/v���\�y=���g��G3T��KWT�"T"D3?)P�,q��#(O=���Zɸ�&wP�oC;F0�3$'�Ct��#L�+�rW8�0B�J��"_`���9P��-��n����4{Q��қsk�0e0(Tle��,��y��0���T�0���$�v��\�|g�bM��g�ޏ��,��,���c���z㡗���_�7c��g1�f�TE��f�E�W,.�a�";^�&[���]�T�q�q��33��iOP�X�,q?�O���.Y"�ƌ�y��&�P=!��1%&Rb1
�N����q)#� T�W�|��U2R[3RRվ����8���Y%���k	�R��;�V�PSM��e��|���qd�e��h9W=}�Usï9��/-��m#��1�O�l��"��l�{����83_����ٯ&�X,{�?�˩� 6�-;n�-� [;�Αێ�o�-̲�ͽB�GFC����nP����{�@��wy9��5����,�u�ƨx���WmE��˓�[z���n��/^z/4l�泥u��I<jx�M'n����aq�-�X?�ao;�)��YWm��z']�w2i���cu�dd�i;g��q`�GH�ԘM#$������"5l ��cQ�	�����ӭ����\sj��l�_�S�ҟ#���U
�	�;�4J��3��
�q�v�c�tc���]m��3��q���=�AK.��YC����]R�S�3N�-"�77�uY)��&֌�7��1��oo����^ר(���'��tǨׁr�
���b�2^#�Z�K�u�;���w<��.Yq�;�wV{M�p{==<(�=@����#o���kGj2K�5�ty���ziY�<i����l�=��<{	�>�㊖��{���u�Y[�V/x"����K���b����;H��\5������{6V�)��2���vS�S�7~<�x'c��R@ν*"���u��q<-�Pq��s���-��w�G`��6�Xa}4�Ƈ�����AJg�+Ⱥ�7��ɼ�܏k�Fut��s���M$\zw��
c*6Ͱ\u�O�c%ݥ��R�(툺�ʮݭ��޻����7wI$�;�8;r�@�4�^���̦`�Tk�<!��4�.��n��4�س�"�edTG
��P��`!Ga��;^Y�!�_<Y-�U�������<��u�5��r_q��ߴu�+u�=�;��]r�)�p�� �ʠX�fy�J�E�E^�u���L��u���%��!�e3N��0�� ~+��vy���!��r��aw��m/����d��]=QWb��\����N�hXE߬��:[��^�Z㣸�.����oT7d���@�z��پ��js9��ѓ����k{f����(�R�1���N�,�v�5ǆu��
�i����KNa�7�#����0��t9�{Jd����<.�A�Zp-Kd8뜄 v�1����m��K)l���ޚ3֦hbU���>������j��L@�w�2�\�j��p��#���7�F�y�6��Ӓ�߶�|�c�)�g����A�b��	�C�Gi���V��'�_Q��B����TY�GZb;�L���>WY��\�&h:;X^��^�)��q@�KbӸC8;^��Z��ӯM�)`�T�8��e��7����J;	��+��Y�s�x��ĳ�u�9S��96�-�0mc]D
����{�8(%Vpu�$4��(W�2�ꥱު�6D>���;�X��>��j���b+:;>��"P:����=�2��k�v�`���u�[r�LO0�ڄ��q˞�]���;Fl�;��˟��(���PQʵ )1�gcܹ�Q�#���ޅ0.z:h	jz����V��T���>��lo���ߚ�6�0�R*����`����a7����
@�D8��D-4(ҍG�ٷ���a�;���U��7]
)���<�;�t����r.Y�r�2ʽ�a���>��0,K�TЦ2�m�f������9�r�k�u#�m��J��]�P�����Ϛ���ǫ�v��Һz5�W�6n��3�=��XK;&�=��4M��?� ���yWK�����3�_�`*��s;)�)�s��x�Vk��ɽ����\��e��e(~r���m���m��'2y���%j9ޛ4u��)��������0�Ϋy��T���#�Sp�a�Mp���nO���/��.:خ7�FJn���h}g|�π�\ �:[��k��?:�i��mcVE��~��K�䎬�7;�9WYI>�y�0� ۬��Cds*���b���s�޳����6�ᓗt����p��%<p+,�;S9Su�Qvl{�4��v�e�6�Qy�f��׌=��+@��	�uDi���8{�z(���z���%���:k��?5���A|�����n�7�
��ř��1���������Gol��������0�����WSȶ޳f���}�� 3y|���.���c�k|Z,R���{]29��[ ?k�/)GaU�(\��+��)�"ŝz�p.\�46�;.4�4�����J���ㄡW� ;V��^�c��]֧�bs�:�I�@�*�=��]5d�Q�������]T�4�|�-OѼp��tȍ=��yS�2�'e���rx��Xֹ�-YB:fa�_^���2�yt5�����P��3�jwZz�BO���d�(�m��9�%�w��g��[b�&x����I����Xѳ`G��Qj�x�Ӥvi�r3�cGWC[��_nzh����,�.�z���*P!k��tñ�P�d*�'�N����Z��F&���63��`�#������ٺ �����ц�x	=x���G<9�2TuE����u�W��}��>�l6����9���PG殩"=*!9�%���ɚ�8+J���k�=c^J�/��hUm.���it]���ck����*eu���5ʕ+jf��0��0�9Y2���������]!�@%�nΗid�V�"7��`�N�K��XR�F4VŜge��T�I�6�8:�_fs�Y{�[wMC�sPs)t�}]g,kL"�V͊�u�D�1���m�M���)�~p�(!ٺzf���5�$�yfĽ��������?D�Ә��[ĩ�0%����Q��c�k��q���é6c��s��O=w]m
�^���iQĀ�u/q%,��&��uX�j/���������(W��CLbJ^˂�^�Z�ˡ0��5XY,yd�q� ��y��S�X�q�q���Z�B<�7@h�w�UW]{;Vm�z�k��#��\���Ƽ|�ٟ��^o�h��~�k��m��ou������(�ƥ�rn�6���a�#@']��t���E��n��ľ��{fY�d8�ش��*�i��n�F'nӽ��_<�����1�jQ�x*��]����r�Sa�����4h����1����l�4t�P�q8bY����}|���<j�C��#��Y��ܮ[.��[Ͻq�x�oo��6y��씍wNN�"�¸T`M;�3N��a!^dp��al��n�Mݼ��2�ʁ�6жon_z��TJ���rt����FYC�)�:lN���w�e���Ȑ���x�l4���G^)�>m�u���i��3Fj��M���!#��V�KU��u+w���� 8�q����+�;گ{4�H=Y�#ȯ���j{�W���|
cϞ��a຋��^ޑN���P=N[�%$s7��WȎ�� ����خʥ�9!���iEA��`���n�-];)C�N�ᮑݛ�-�)��4p�6�-���!<�C�S쵰��/�O��i��%�nl��u�՗�/ڠ]��B
��G�^_O��=<"� "�˄�[����\W5�i���7UK5�x��UE�z-�_Z����F�YXy�bz!����W��	+i��d�6��5���nRs����@�:Y��i���|���d�#�N��s����W��k^�n^��͎<�v}��rE�Otء^2�l�:��r�;�k���q��6�Q�6�.�؜^��~@w��wE��|��RZe���vW�d�r�i�x
���v�z[U֔��ŭ������pu��{�X
iS�XK��.���p��>�x����w�W���E\��;��tt��9��nN`�o8��x��h��r�"f;,��um��d����ڟ�W�:m���l�����ħX븾��؃�s: �+��F-����(Vh�t��#:��"s�N�;Fs�͎�������K�k(��n�e.����?ۮ���ʹ�̃���?^>[r�k�^
�.7��bt�]sh@Ȯ��hf
hF��U��C��$���뾍�֌�}�W���?1�������E�͙��X�cr��	0�l��/V�w_gs�ײ�[���E�s�A0��K#3a����;���N��S��E�X!T_�m	C�����=Qrk���<=ݵ��\͞����!X������Y�N/��nU0<�3n��[�s欇7]��/�'����Su��2�h�ҙ"�bz���>� 3��h~ɯ�D'[�	��ˣ�9F�?gFaTܢ�KvT�5*��i���XM�������%�����p5m�6��6�L��x��b���y�(�۲�ס��%�(p����:��d#��-�B�Tѽ�l6��Az�m3�I����XQ"7�Qܿ*�8OD�دg\v�� �>O���j��baή�c6�Ȩ�z��[�L(�s�<W�۽�S�e�qZo���e�tp�ة(�����%۫xi��=f�JO��<�� o;�5q���z���wZ�B�|�ն���Zp/��k�+��Ť̩Nm�pOWm��:�<����c۾�~�dK��Z>��X8�a����ݮa�5t����~x����o�tҟ��Ss�R�hG#E�
墦�1"̺�v�{0ܥ˧8�^^�IS��49���`�6����鈉P���P9<���j���%��GO�-k��v����A�>罶�j�n�����Ok-� ��]�A�un��]�K3m�ur��s�3��D�T���Y8��T�{]]��U�,fі�K
�+b}�n���_o$C[sX�&]����]�t
�!ӵN⑻mv�Ǻ�מ��-�yh~�og�?��������� ���3�č�>�7�C��dsH���Y%�2*��D���9˚m�x����L�c����4k������a6NC��� ���%���k�
�Y~��e���{�G���.g<a�Dp���<ⱶ�TYŸ�x���>2%��8�2�G�����|�� �-�u�K�����9j(8�{�>��m�w�:��[���͝@�A�'M_FKu��]�Y���1��wu����j��V3B� &�'��:����~�Vj��_�׶��a�/���虾O�+l��[��7	z%���@Z�Sjy���GaTܢ���n��Y��8r��"ŝz�p.�Y�zuCl{~�Z�KC��Gy����5�;�l�����1�Ѧ�U��֝�!)��r�ԁ<]���vY��@�GM�{T�4�iډ�O���Ήõ>��O�gbvZ�������ke\�86x�εB3�P�zf��:�Q���	jwZ{�Ѐ�(�=<m��r�����Fa�Շb�ua�VPM���.WM�-��[�F_i��ڻ�/n����;vB7��ζ����#�D��-Z���]�!�{�/Utʋ�.$(=sN&���I�;pὨP��v�pֽh�Rh@,hW$�\���;�!��=�L�A�o�	A�R�\j
-���p6ףf��l�T@�j��/E#�긡��5��)98��횡��s#�YOzm%(R�s���`����o��6B�}T�K���LcO^�Z�ʻ�:���*�ا��a�lv�d�b'�K�,������'��p1c�s���T�ej��<��������[�#n�{c'��6s�;,P੺`�����l<'YA&����]E�ӑͽ�t�':s�%�i�:J����,��|J✕��L��_JZ�Q]�{mj��"?-`gŮ��fɀ2&�ۘԟ��0(TmɖC��Y΀y��Q�sJ��]��vê VS�-�3�$��U}3�z��c�kOc�r8\k�(D�s�f�1ͳ<��Ԍ��rF'����`#ͽ È���&k�_�������X�u��֨Ee���5�sr\,;fcD��A�%���Kot��*L[�BOZnz2[���ܲnh(�'g&5Z���R&9���9 vm�']눝�A��Kӛ�u�	��|7M���*���F����ߍtиc�\�^'E����:�K�ҟ]��ΩK���m������^]�3.Y��������a�*�
�Sy
1P�o�d�)�ӎtΤ�(�EG�\������j��	;�C���pѴ3u�ed����kz�Z�a-I7/S)l����ˀ�웘����RJɓiS 	:�ήV�aQjxؕ/�.M�I�%�Y�r^�1u(u�q�����gZ�ݓ�$���Vf;I%��o�t:��H6]�HH)��ҽ��D=�;n)݅�:2c#����UR��b�C�n�H���
�a���kW3�0�W���@h̰�*���C/�]�%X�3�4�J�N�5��V\Ŷb��Mn5�ޠ��B��P�j>��uʅ^W:X���q�NoV0�ܾ�u��x�f��s�����ƻ.��Qor�+J�Q.�3I��H��z�qcv�EKg�VW
x��J�tqU�َ��@�]��2ZH&��Mp��wZ	_f���� �x��"��s���uy�P������w�!��o&|	�*J"Iܕ�=K��BBmR�J�R!�ɪݥ�F�e�V0����U���՛���hN�R�*�E<�\���ס>ݍ�).��3ˎ��R��T��W+y���C�:��|x5);�F�W�("�����л:-'�on&Lr�����rj��]ŕo��GK�y�t��e�������*)���bڂ�A3��%qI)�`�tAV�q�����d�W7�V�O{$�F,�ǲ��ms��,���v-B�Yq�s����і ��׉�a�����RA;�Hg�[Ň����̩�����'��$2S_�ˇW�@���Q�ϑyYm^א�Y�o89Z'ܕ��R�1�6v�AQI��J=)�S:뻪�f���8#��`B4�5{{nL����a]��ڃ��FP�t��wp�)6�`	>��s1�X�C�͉j���T,�,���(wIy��c�ĩ���Hj�a-
Q�R�4�n�b�;'wZZ*�Bi�tM��L�)C��x.�37)v�;T
 f��Ba��K�R)T�z�J`���*��o
�|�e����};sZ��;Mn���ݗ��W�ǏG�ց}�j-F�R�m(�`���$�q���Z�4��
����5�<�M�9q[�<�/1�ɗf�t�� �O��iM!��V���k<{2���P�˺�
c�	�{r6�>���.�R.�K�����39v��w��ʒI5:��C%:��n�o���Xe�̆�{�)]��9.S��:��D\b,�â�\R��Qk�����m5J����ޖ�
<֌�� �qۧ�V�廐&��l�Ki� �X a�v�S���Y�=���ՙ���*��V�תR_E%vd���Nŗ1�F�ǔӑVs�zU��}B��"�Ȫ�)K�ʪ�#���E�.U˅��Wp���!E�"���d�F�q"��BIt�A2�U9�vI#"����H)�y$UeQN{��2nt�T䃙Uӹ܋�E�q:t�\��.U&t�a�("�.��bHd'(�e���Ut�ENa�Ap��2���!��*�	�듑t��@QTD:�Dy!y�4����q.C#�IE2���Ez��T�΅QȊ���\���D�@H"i$��N��T�'r�Ζ�]���S.Q:1�*�Õ��,�T�D�J�N\�����E�wi�nC��*���NGe�
*�L�*4�$:fpL#G I�QY�%2�ӚRe�N]P�MB�� �]B����"i4���HI���ފN��}y�u�[SP7:��3:����D�	���ƀY��n�PW+ӵ,;�1m���d*޻y�/���A�w�f8�ƽk�q6��7Y���<��ϰ�����#uG�L�.�Oge>�e���O����Y��s3��)�zz"�C+����|�h�O�\uϱK�[��T�Zz�K'��m]�.����#I7͝��鞷�R4�踰v���+�Fh�S�iU�w%�8HU�n����="ﲖ��&��?{'dq�][-��t�]��\�)�:teP���w�g���y��U�}�K�ʊ�m�Bt��Y��岨\g�cG
��-���(x��-l#��@�ϳŖ}��ͨ��=�g���K��>�xe����z'��y�*J*�	<{��@�������Y���b��?`���e0�z�w�v�5����t�YXy�b'�J�Q�Rl�ᯄ���M�I�&6�Jǎ��Q��l@��$M�(�y�Xc�w�������i8�T�kM���N�/;�� w�c	�-�4Ŏs$d4�M�eFٻ�l����q�� I�����dE�Q`�L�-qr:J~�'��uSE��Ϭ�O::� 
�r�e���̯0t+{&�l���\Nd¡�i-����"��V3g�x��')�K�kQ�;��r=U�ø�b`B��*�\�o.�����f>�7M�G�%U�2U��Wa�4\��Z#�p��_Ts�]�}
d8&�Z���X&��os�ʵ�;���h�S[Zi*�&aAU�2��ˤNV�M��ԋNVV�u��zI�ݏf� o=3�c�S���������x�d�C4�[�V���ѥX�t��������s>�m�C���`�.p7�����W G)�p�Рq�r�3��ul&��t�O@�H��m��66�{��w�t4��_@�mt��O;C�|�[�b����jx����Y��?��ᶳ&]bǊV�'C�M�Ku(�����_DXv־9ob��NW8�m��������t�r�<,��ַ�g֜_>����\�:�s��!H�������������4�ߘ����A��"���־��j����C��-�9c�j�|~�۽֫���iT�zd�O�b���:ZY]�Xi��~�mZ��>�{��٧Fʚ�n��0�x�l�\��$Col ��c��6���Y�l�A���i��?KX�a-�s˪ݪ�3늚���/�h���w�Sx���s��t֣G	}ء,��M� BX�à
vꈀ�ﱇ;[,f녀^�B{:�S	��疢�.z�vJ[�k+��\zΨ��"������[m�=��������&�l�G��0S�v����F^Iӻ�z��j�t�⮶�K"��cX�=Mա���ӹݠ<n;"�j��ݼaun������jΦ�p�]:�Ӊ�w]/o����m1|G^*r[B M�_b���NR8Z�[X��l�p�-̧�1���TBM].L?7���d�7:�Tl���S@M=i��N��f����Kk[���t6��q"�LY��AN��<�Ӓɰ��vt���@)��ϲ!Q�%>��j~Ge�#��o�e����[v��؟���#��ҩ�K7tq�V�;�v}��g^2�M���
�w�a���nq����v2:� j�WT�㻅0�mq����v�\���kwf��E�F^�}���]���&ѻ�n����ƙ)�'�׎ l���U=0��w�4�R��LLN�ͭW�yƣ�� f�]�sz�a�%Q���3���΀�p:����V�W&S?\��������r��	�,a��98:���[�e����k��he��|=�fu]`��z�S��(��_�Op}��������q�#�f�������ϳ�{ty�:[����a��Xk�:j��Df
�y���L��[�ِ�������f�l5��\�T�k��c�K��4��ܢ� r��Hʣ@���=��*�\Pޚx�9��'�g���"<��__2!ڭ�M�����}3�N�|��@�P7���|����vT��+ZS:��
δz}������_�3lV������=���:8�9�����o�m�L	���4�}���.�9m.�x$\��69�d��?T��/�#@� >��/,�v^�3B��r̝
��X�(aN3jJSZU����QW��0��殛��&��YL5lw�y������=�jtSv� �j��=N_�д��t�k%�\������忋��V��&��;M;���ap��:dCi�O�i�:�e��L�5Zk���j��R4�gI�<������:�I���	�u����%9H�-_����2xI�ɾ�.�h������Zj
-���&S�eF́ʅD
��_�#�k��nV^3N`Z7
��B[7���ǻ1�=-�l��˄�Y���r(^B�F�Q��	77737h�m<�Ǳ�5�	g��2���9Wd�bzT��e��,��\$�n�j��ԸK��8ԷV+��uT(��{��n�9����#�{�ԩ��y�ӑǹ������U��7�r�𓃙����4\q;�b��{�lJ�|!�m�L��2����ۄJʬ�]w���(���q"<� v���9��^M)�0&���
�ʱ�5ؿ'2�?	�ߜQYet��q����n-.Wi�*]�i[�#v3���:8�l,�`7a�
�'N���t�6�MH>�R$�:��*�[����������ݖ�`�pa���[aǀ�S}x���'�y��tj��}���C/��6�~�7���>�.���w��G���#/��][���L�e�SϞ"�*��t��!��� O�Y�I.�u���������������x<��(�3�����m]�t�c������7�68��`!��qܜv�TD�u���ʙ�㰼I�)O�x�K9���t����3Kk��!\s���|i���-�B<r�u�z2[��mȆvp[0���S*�Mpb_�{ͷf�q��d ��O
�y�%�a�>�}�+�(KoP��y��	�]&<�O�\���c��c̳��~x��l��8S�P�����w���U�k�3a�1�RPq���͝p�a��±�t� �U�sK��~U+<�yM(~��b���[��'��zX�\	#�b�g�)��'�O��T�6k��6�,�<�t\X;^��.£i�і�~Ұ����q�v�P�5��q�;
�{�a.ze��L��'Km�wG|�����`B�T`M;�"7�6t��W�9١ms�o(��ϣP��Zn�F�O�(<ޞ�� ��(}*g�k`��˅��	vW��j���h3�vS�2���i�<�n�G�����=�µ�
*��I�������!���T�X�x�a;dc�f��BO��3��o;��m[E1�5�2`�-��f��չ[7��6�I��J�} 9+X�Uc��Y��=��^.�Wa�}HJw\�ukY� ��]���XC�Cy��wN���V�Ns:����~hO�:�����yf�d��%�coF�wXy�4;����V��w1��/'�0՞�7�� b!��X��e�ЪfQ��{���!���8�{	�x:h�@��F���CJ{�����s���$D��s���~FZݟB�h�"�(H�hւ�G�#Pzأ������lO�4��:0�����/�.�	�)g�h��~���%d��'�]ծ�'^ig��x�m7��q͎��oe����<�w]0&Wa�;^]���D�-��爝ؖ�mZ�Y=�K�;�����9,F�t!��������L��l{ Y���;������O(�q{��:�m����u�Q|����1�<�~��Y���+���w����Hܦ���!��7߽O^����1��R��7�Y��X��!�ݐם-ӥ�%�gC�{����w��Z1���~��ܮhN.�.w�X�������?*x�X4���a���k�aO'�`!�l5��9��Y6f��cż��=�{~���D]�lw����^$Z��L��4G�~��~#��1=� }��Sg{���˖3ƻ�C�x�0�[:��	�i�;�V����x�d]ywu���d�49lm��c��p��T���]����u1��ˢ̚���oO��:���V�N���6���v��t*��O�F���7��a��/�'�x_j���og�:P[��SX���5<5U^7@�O��ڔ���>�;jN��v!a%lCU�ej���1�o^"gf�z�n�m;A�Pj����l��yfSg�����#F���FYC�Gb�n݈+Q��`�@\�����9N�7���lQ"7�QܶT��;';`��:C� �Ug���)�d�����2�tۺ42�T�Z��<�p�=eT2T�d�\r�.~�e��l:v󹢩ʭZ�[pN���t@Ój �3ϰ��l���S@M=i������5N�e]���n]�/��,��c�z[��j:
X�v�`�0.["iF����v�\[����Lke\�:��D,:)���TOiS��%�Gea�xuS�οEZ�۳��"��Ϸ�ʅ*ڙ��]��`�<�86���h�!��T�
Z�鈔��L��[����9�5�g�F/�Y��{_�~��5� ;�����/�=e��O����@�S� <yS�(v��\�@��v�o���-9y0t�]�sU��D�1�쳜�� o��b�5�@A�e�p/�2�(����h�;j�]���7J�j��P��[����x��u��83�ۥ%'�3���jS'3�\l괁4�u�����%������Ԋ�Ź�9ʷX=�Ii�ޠygPo�+��ݤ?]�߽�����x�{�_����f��xaI��P���3b;\�� �������m��n�*�Ўn���(������Dd�1c���O�A?	c%=��s������{�##�#�-��v�<�9���ep��|���?�ʺ3�G����k����Si���:���$���߿2���}��V�t�*_��6nJs՝/7vE	[f2�7C�;,�%��38�ً "߷���Mu�A��m�{����~ U�5��䣰��(�pg��`J��L�F�|;��2M��h����~�s�q�9MM��Y������Tj/M�r�U�6��V(��&y�u���o�Xc�r�#��GN�V��'��i�}N��鰸J|��"Oj}�ZnD��յC�.���:��R�O]�䣴��D#,����ٰ#�P����(O��i�ly	4�j������kw���@�m��y���a�Y�=���m��<��@�q����U>�y}��90��D���Aݹ��6<��-�cF#�o�Ȥ�����N�l�I��Xv>Ê�Z�Oϲ�^�}�  4Rk1�+Ύlw5e�u���[�w�����:�1Ӷgs5�(Ŏ��^�j�����ޜg`յ��eN��]@tq6U�����T�ݝN��E�����Xu}g1�J�#ٓh�s�b��iw�^�n˫wo|�_T�����-p�ӏ1iYZ��z<�FaBY��0Χ��v�'���s�R�O'�x���a�`퍹v�c_�U�ތx{�d[(��C.17��^㑓�`�#��WT�UYE��Y���˴Kɇ�r����F�.���T��ٿ��_d7K�F��r��u����Ń7;]�����S0�N�I��;��[�J�si?a�
��v{����/nXz�Or��4㓧<ñ�T�c��u�i��Fv��9����c���:+t��pr�H|m۽e���69���7�vs*��o0x߲�O���4+���³�����t��lL��H�/O�FD:��
���sc?>�����<�s������Ǡ����W2���rʽwfZ�Gr�c���<E��Jƽ���=ݱA{�++6?K>�?<���R���ԕz�,HtU����Q��:¡�`F�C^�გ�{p�tXzP#�j��.�q�o�
�u���o�c�\���C<�iC�[����q� Y�F
em�u.�~z������Q�t�d<�n�2����u��h}Ѝ�����wh��ùI�P]��g8�fX��ލ0p�ީ����&�p�E�����b�o+��j�K`ל����y��;�ESݻ(<��ؖ �]Y'l;,��3x���W�<�/�oؿ~-���.^x�����]�Q�¸T`M;�2�N��fE6��U��D=Ix���h��'��xP��A�?o>6�l�R듥���D"��)���*�Fjv��= 5�{��&����D���dHH�0.�!i�Ut��&tp�z
[+���P��nS��p%�n��hD�ML9�w*@��|Fi����8*d����p̶��c�:8a�:y*v�����|�58�;�5�����Ǧhׁs��L(��|jvK^}YP�y�N�Xy�hmK,1WC����/�5����9��4�6\F}nψ��|SB���:}Oݯ5���2{M�]Ȱ'5	gO'���[�x�2�}�v��NpS�g���W�䋆��B���7l
�ӹ�Q�'G-���#��9�O:8��?0S]R�S�9_Y֙�g��Ms X��r�N���jl��QQ�Ok�k��E+}sӾ9�>#�-n5,+�!�Gi%ݵV��qW3��*��1���Pc��Y/�zʲ�Y�8X���o�8�ͯ;�x��!�OK��3CC�����!��dT��1��k�Z�������Vp�V*B�����+!�ŗ�O
m�eqC�˴��E�iݙIc�w�cS���Vs�c� [�C�ot�ה�nOv�~�\�w^�\1T�"� ��4k�a��J��׮�z���GO ������Ń��`�l���
t��,q���RȮ�
�^�/:�NF�X\gT-�囕�dS9CF�p�.���w�f�OS�T��22;ٗ��.꾚G;�wVҖ��p ���WC/���r�ܠݥ{�^�VIX�����Ե;pֽ7�,X7f�EF�Usw
�Pe+�|5T��a��x���PSu�\����j<0���\�KcgU�e&[�Fl��w�ÙC�1on�8k��+�����E�m^K���T��g�Sz�Lt���ե�.R�j��]��v�4�츢�愲�J���#F��k)]i�s��F
ϛ3�#�����������V�}ɹW˶�[�쎈q��qO�yݑ>ƳE]!Ţ��+���O�.����-�vGܕbA�8b̀/{�n���8>�/V%{�9�7����9�tu����S#U�;�"�c�Ghb��]3%Y�K-�w�%�Z`gH�4{H�N
S%��b��۝��s[.R��K��I����g��k+���J�hoZ�R�GW7@��Zs�pV�f�1�(Pf,�7w����U{��]a�x�"�� Y�B��7�K��J;ϵ�
֨�(%�g������7�[a���+]&�=q�7hu��d��U�N{��{��H���@+.je�+JC��8m�f�}��h�U9�7c�VKwj!e���E��\�}=h	��A��;�,oz+�u���C;�S�h���\���m��v��M֑B�Jg7�W^�]Kx��'����H��#ץ��|��� ��mJLع��d���3j�vdNm֨#��K�O��Ӫ�f&���!�,�"�-[�K��=��(��o.��*m[���ك��Ǡ�,��Q8/��{J��v%�z�1�DZ#�JM���{�4˷��v��S�ce,�L���c��+\��:�N��n��2	O��5����G�=��g�M
Ո�U��O`��T�.��<	�(͚�L���:^ڬ�t<�awfFUnҏ���V�U��Lj�|&���Hj]��sv㡻9U�B�
��9KE
�䣬諬S��&LU�-�W.3�9»,��/;�H�/#Бv^ʷ�Nm�:+֫���0�`�Y	Wr���*$�9p��ƒqn�]h���-�`����lg1���W�ԭ�5H�������}6Nup�E=*��K�L�}�+��X*���%
�B�/���6Gb��-VWp��Ǫ�Iғg��B��@W��k�%;}��+.�����Omc���O���1iΔq��7K�3�+%a����{�X���D�M�[#����<o's�$ɐ�F���ͬ}/�)�Wk��h���]�l�g(��n��ԇ)ݻ���=�RJRcm����㧠5�V�U釅�r��嵱����o9�_<=�j����>�&�
��(�d2�v��TxM'�

H
�B^�� );L�$)8��l)�QBg#����'"�E	6�*�kWq�r���n��"*N2�L�T$��wc�Vs��;
ng�˄\�W((s9�9�e�"��5�\.S*�\�H�(��nJ�Q:ĊN�ykL�e]���"!0�d\BH���I���3"*(��죫lI:v��Q\��� �T�H�ȳl���FI�9$vU�S((�(�J�s�p�͔ˁ�.DEf�9J��EU2�t��NTU�gJ�
�K�U��+Zj$\�$U�J+��KYTQuA%!I9M+8Jй&j���YVa���(`#�S��J��=f�~[\ʥ����mOA�����s�b��O�,T������O.��c�@z��s]�;w}�w�&��(*_�������k���9���K��.;�f��:�@�0غg��魘I��Uî��:m��2�hD��?a�M��:ջ���>�O�(��n�e*st��ңM֐wj���̮"��w\ЖΨ/�c��<.�����F�Ӌ�a@K:=�6e�Ov��l�ͦ�ڷaM�y�]�vu�B���`������V�����hM4
Td��l�D�w@>uÍ�� �6������r��ݷGKJ���u�Q�uv����n��s*"'�v;ޙ�s��[!�,��#V���{_�\��^�F��I�zyln��:lؗ=Մ�S��r�:�@G^�4KQ}�4��x�;���D�m��w-T��Y�'f�tt��_��b��j�E2<�~��C�^O�{U��u)�OZ�}E�\��.�b���������/�-�>Dd��u�S�d��~��q�筐5[D8�u�=i���t�с݌�v:�a�kB�w`VH֍ݒZ�Qnm셆��Y��a�
kvt��� ���ϲ!Q�F�hui�L�����j���8������*!˴��6sx�K)u�t�S�`��MC��O	�.��A8��>< ѽ�ں}+N��]�����U�U�A`� G���#�x�%�ǜ���z����|�t���>�(�w7�R	ɢ���w�;������J5��ͤ�W������K�ÂY�����#���S;��Z-�9�����}�=��\�ݹ7uV��/�s1��n�?�0�h�(��9�8�]t�CJ�e�'�ۡ<������8�t�,�p�J�耑���vTc8?m��2��8'��ܤؖ���8���g��z �>@�����o=�Mm1�*�a�U��3����p7�k��xm�mB^`���d]ۓ�_0�9C�/m���ݷNN����n��xf��F��M����(&�䫼\&5�v�bt�lB�����s?�E[��\U�[�����X�q���1��Z'�$����h�[#n9��s���S!�:���>�s�団%���^-�YړgZ��{�q/�f�Bߛ#@}xDΨ�%��	�O�����-�V�yɓw9D��g-�ٕе4�-�=�Qp˚�6L��}-���� n'�.�Y^��j����;�z���y߳S�i ��'1;�bλ��E�D�\��d��t ��Qy��h����;-��ZX%{X����}]XiG���a�XJR���/3J�ʾU����X��u���g`�T	�g_�wM1X�iZɪ�{��pj��v�i7���W�$)�塔Z�(�Z֫=�`xc�[��=f�YyJw˩�\s���Uƺ�q��f2�]a�uu����}�z8~k K|�,X;Q�`B�T�>�{N���ڟ	k^uP��|p�_%��W{�m�7k�2���+�OW�D#>��l��
��jz҅��5�趉�h�}V3������(�"��w
��StV�ui�(�Sw4t�N��6S� of�F1�f�y����T��~�\z}W4��E��Öˠ���n��t�gH�;��x�ƝQ��7��ys�,sleH'��S�[5�	~|�:�*n�"��(qm�e��g�Kn�����>p{~�p;��5�\��UP�&V��\2�9��<�=x�9T��K���x�S<Y��-I4�n��,��a������\q=�b���׻ )5��ə�#K���/tUѧw�����9\]�6�����%;�l� -2���-�& ȚSn`M.�@�N�о�q��9At����o����v���;wT�,�_����tό>�t�9X:�oc��[�<��}�U����5������J�:qϮ\wsr�F�#ܜv�TD�u��v��K���$������+V!���hWR�y[u�k�hTp�h��.,fPlf�N
�1دL���z��5C>Z
ƙ���v+�[��}�������󆝍A���r��]b����r���r�_��]C*^Y����'�8��\w�S������k�/���fc����D2̞��ˢ��-y��K���]�� ��&w�:���8�&{�v�_�U�ܲ�w�meqǟd �tp�g��܄����w�KkT(���V~�d�7��+����/��ٹh�f*���=x~e|�0�� o����V�RSwMM�;�np؞�1a+�E�'�奟�O��g��J���F��a�V�J�+4� _0��J�����zow]�e3vܝ3�od�i�.,~�*�\$6��1�v���&��Kz=��Nw�?o
^�q�>��"<ڶyo)�\��a�1��im�����)ߣ@�Y.�:x�\-N��cyw�X��0;�w�Y8�f��ZqK���:8V�-����#$��I��d<��k2���*����U� _��Q��t��~�l��6B#�zx-�kw���u�E�+�&��qq��m�`��u���OK�杒׬�e�Ѻf��Ȥ�\œ�7����4o�J������:_���[��8��*�ЪQ���~�yf��d�����o���
9��w)wƑ��5[3�!��z7�uQ��������ȗV��y�=��⮭�w�\]kh,ub>E�'��^��r?N�9��th��u��O�ʹ����P���kF�ĨjUy�M.�mug�߱y/Xg{����t�]ٲ����= �|��Ǫ�(D���E�ͻ>���rE�OtءLeFٽݥ�%R��f�%���{A
M��C1O�R~MuS�4��@:�i�s��즹�,u4X�׽����]Tu�����(�w�´�</m�H�7�6��n�%Oa>}����t���w�r�ckV뒛V��%�e��3Y�=�X���f�6�@ލx��FӀ��p�f��Q6{�7r��>��z���R)��I]�����"��	O{�u�0��x�� �zKI�W��Z�h����y�ˬC�I�g"28e=E5Qg�P��PY=Mٹ���u9ˉ{�WWͳ�{ׄV�3[��y��Y���.z2x]=���k{f���ȮkG2u�=��;q#����n}�v����P��&K^���5��sF��L�Q����I
-\�ՙ}@Evk��=|�_Kd8ۜ� ;5j�������:ZV�Xi���z>1�R���'�Q�e�SZ�����ޜ�^s��j�A�Lu���4W�lF�}`� 1���]vA'�A�KQ��?5\����_P�c��u������;�>ע�/�'z��
Y�I֨�ozfv��Aܴ�{�}[J4�Cݷ�j���m7�,#f2Σ��1����X�3$�:a9!�Ci�E��Z�#��*Y}��a�nNUq�~n���OCP�U4KQ}F��u��7�hO��;t�j�G�a3��Ū�R���|ڲ]X�Oxw�H������fX&��FY��K��%�)lS�q��mj�A��ꭷ��{1G�k�3�讞�ר(�5�I��P�hفf���������Y�|���] ���(1s��^2��*{zsKaYgx�=�=-��N��hH�N��t��wRd*�#{��r�opkM:������VF,������וnGC4��g��o���6X�V�l�ԝ�3v���L�c���У/�ov�
�0��{~Fq�0���S��,C�Gt�	��_�Z�n1�1Y�w7�'�}��]�4�J�z5�W�,���(�S�O����$y]'-�޺N���E攥��}��x���j���(�=�'\[��0J��i��e[z�y�j�9������G)���7NN�X_-Ց�߯�O�]�k�=�������L"�s_{]�;G��lQ:��>�`��~��ʈ��e=���f���:ҡ2��h6Қ�ͫ9dx+~ԝ�lFQ�=���%k;g�h��y,�=�yR�N��gվ~���^�d+�_ܡ�7t�� 4H���^����sp����7wZ.��=�3ݔ��:�%V����9Tf���)���7��̲�A�h��= �3th���\t0�q�θ����uA��Y�֛���n��Q�!=v�������Lu���^�5��ǖ��������=���B��7u�	ޫy�%���w���^���,�e\䲫��3���r8q� }����v���M��S���g�e�gl�b��v�r����ȸW9M��|�e0�e���.[: �u�S;�)�D"��n�{�&�d`�ۃ�����̢,X;Q�`B�T�-N����OѨ�	 ���Us�ľVne�eP;�wq�2���v�f��<v���Sˠ�6l�DM=iBߦ�`#rb�r�r�zݗ���q	(�<˟����tf�[;��
8�+^����l��[�U����q�l�s��)���?#���9���؟��5�p��=M¼v��U��'��^4�[�I�j�C�a;�
`X�n�RIZ_=O�l�f%�:7M289O\�b%Nˇ�he���e������nY�ǲ��#5�� ;���w��g��r�x�ߋ���)\r#���U��n���0T�kl��&7����vEz��&_`�����g띈W:ޏH�.�4�N��'WY�+�P{+ՎoQ+����A��*���mAK�V�{��Ŵ��CV^n훏��^���F�QX��[t[�eΩa������ī�<�7���f�,gs^��}ڹ�m)�9�*#��N8��nϨ�E���6*��׻6Ī0�|!�3��V�&,��k��k��M�~�e�8�$CJ�� �i�y���0E��m����S����>����&��'��G>ƻKq���v0�r�$g�~�.��t�a�"��S��1J�VN��a����蜍���M�������(x�,�t�9�����o�� 29#=�Gp�������Xq���3%�ܢ!\s���ƙ�����^��_�%MI�!o�S�;�p��p=��m�j������r�[=<(��#w%�]w���n�
~ۇ��o��G�{"��mC�n�#l�(�q]q�ݷqe��/�}�0�� L��)C(�Wʣ'��}�F'�zy����tZ �ߞ���V�V�7kk�Lif?���iŧ]o�&Z�vMi�Fx���a�j��N��?.���m�:a��=�ٞ���h�a�£ ح��\��"_-� &� fyA�[�i�lw%�8H�հ��)�\��a����lM|"Ne�
>��mU��Y��T�i|�p��;c�w*�y�>�}x�DE�-OP����g�'׼U�Aι>� C�tyF�i��j��i��CHb��^l��yb��ѝ8Wl�/���k�J���t�p��Wk��i̺�Foa9ib��姧�#�֪�
�(�3*r�]}n4ν�dFh�D��nQ�`KS�q��~��3�O"��-9~�q���z,u7\�n莎�6a�m=�>\�ܛ������ꍎu�5�u=�I�r��Zr��t�b~�}(`�BY� �"�*W$t��w�G2�T�q����Q��S	j�\^i�-y�eC-��55\��敊�l��;rcO2\c�OO
c��T�< ���#r��e�M
�`e-Oݯ��R��>�TR��km��� �j�:��<V�U�⥫�H�J�NtW��~Fm��,���.{����᷒j#y��i��Jac.���;�k��O�#�-��c=��`���4h������Q]x�V6������s%��k�9^
���xm��ly���s�逕a�����6�9��u���x�۽x�YkUE��=g�
��G�y���mx��i���ёl�ӏe\L�T֨�xj<���"f�Nρ��oQrʚ�9�5�d�\2�٘CI<]�"ۧ#.�|6� ���C�S��A�>��a�����z�
i�1��W����9�nʆ�����!z��b���x�C�T{�#��R�7F����3>T{��D.W[�ls�n�v��W�H2F���+'�b{���ɽ*�c��K� u�5+PWcJ�o�vc�{�a��u�:m��2��
(Mq��z�R�<mx_�7���l}7����M�7/�����U~ǰ�ݳBs���]�_>G
5Qc���</e�����7|�RP/�y`�9k�����O�!g=7mC\OeѢ��_,�C�7��H�ՠf�6�sc*�V75A��:9[���jru�B >������S4//�oKJ���3��*&z����Z���W���sv-&]C
=׵0'��h�5[��&��+]�1�z��Pѹ����~l�������a<�=t�5l��SD�}ҟ���t�H���w!��#W�"�i��ٳ8������*r�o� S���X��R�a&u>�tWfʨd�Fkd='Ț�˼��Ω<���������6=Aӗ���� X�*��������q�j�q���fmvOF�͏!)f�;���dv�qf;���)��9B��p�G�5~<���	��̧ �{J�?���Y<�?#�Y�";N�m�ҜQ���6Y�.�2�^��ü����cIK�[k[h�^�0(K�SB��,���蟿���޾?��_�����[����a�����v��1�����1��co������1���clcm�co�lco�6�6���6�6��m�m��6�6�clcm�lco��6�6��`�����1��m�lcm�6�����6�6��co�����)��/>6��\/�9,����������0���J��T�TJ�QR�A	EJU
EI$�	[0�"E)R*J!J�UU �ER���j�QTJ�s��A@��@UPJUT�H*	U؈����K�R�8*�)t5	���E[2��-5T��Ck5MUID)@� �b�%I��  ��  ��  �0�6��aiTlT�2��+j¢LXؖ����j�h
��U���s3j��E*�R��J��(h6�J((	I��  �-A�Pm�%*�U�N  r���@�D�� in� BPi��)�X�A�����	p ��L���&�R�@IhRP��V�R�`� �T �I��)��j�Ff���dIf6eIJ��� �%kFcH[5U@IF��m��ѵm
։Z��@�8 &�k20������х�i�*$��-�J E*��H\ ���I�J�f�J��@!F��j3�2'�J   �44ʔ�j4i�21i���Њ{FR�����@0�M40��4�ɓF�� �0F`��T���h�4���C@ "� @)�1M4FA2z�F�jA&�F�*�&&�	�L �l�q8Ӈ�o��g^�dR-�r���"���iK�Dx���<ª��S�@ �-���>���I�*��p0�d@X&~2�(�#D�*��@��@[�wy�t������һpAD�F��M #\0��&��w(�$�Dg�=T�Z�ؖ�uV����\��ܒh��,
�����ۛmm`0\�ܗ���3m���J�)5c�Mn��B6+r�2���n�z.��l�7bt0�h}h[���8� #7����@�mn�����:�,���6��5d�0��}))� �q�Й�5�6���s^L��A7/a�n�Qص��P3R�*����q�:H;z��ՙRc���ŭkM�����z^'��3�T��<l�]��(�MA%Y���Q�vf�����2L�X(��5yA�-nAj8ħvY�6�����Y�22���]nP��&I�����i�wb��a�q�X�m��۫�BI�*��A��aP�Eѐ��Wr,����lԷp���]h�,U����(�� �RQ��7�Y� ��7r���*��ާ%��z�}�%&T�d�Q̨�PUU���:,U`W/6L��ZMc��OU�ie�,�Ln�e Q���v.�U����&�&帅�)�5S[$�2Uf��U.�t�
z���WMXK7u9x"�荐Dw/SF���vjC��#��4�����ժ�aXҘǏuܺ40á��VVVIiR�Pq�c.]e4F�.��ݗ�!
�5�^�!^��I��@v��$�&��lw�^2++2ι�	��e5f����Z�)bw2��Ӽf+��P!Fq��C%X���Be����H{��ē�țkc{a7�Tz�UMŮ ]^��d��KW9p�WN�i�h̢��k\{z�2�8�$m;�m�� �ِkQn�9��^ͦ�&-���2�B�e��L�@�n��X���lMu�P��f���J�ڹT���H�3K(%u���E�Ѩ��y�p6��q$n�ո��`�*�RVP[��ݥ�`"�� L(/l�2S�2:��޺�X��E���j�Ȳ������8к��&�-D*'J�ׄ=\:7+N�%���=����tW��h1��H�FP���똥-��a-�m��]�ԛf�jb0	�^��(��5��S�����-����q�����f[�ٌ��zwBh^dM�f��u)��)6k$�h˫b�۲Z�Xr��ll��[����_4�|C�D�.�j@/T �!왙`SP
jQ��R�2�ͭ�-�l^���GD�ḴS�RS. �|�N�5ø[j��4I����\]�ܬ�܈�wOp`/]0�JU2�nt&U�Z�+���ث���!րn��;��B���Q�X5� �_!u�x�J�
�kbc�mi0<��	GH����Ma���X�ĆR���Z�)A
����pV��a���F<F���ȶ,�){�L�������\�6
�kY3u��bk[ &3��4A��[30��^��V;����`��6v��c���6Q˨E��՜Pc����-i��#՚�p��yQ%� �̹͒�L��WzP�Q�ZQ8�4V6nXP�d�^��6�����tf��l�YwrY�;�Iͦ���%;�K���	��xP�x(V���9wV�W��md�U�z��ɗ!X�%u �X�^�$e
4�8�@�M�U��K�& �a�X
��d�Z�+6�v̥(+7�
�@�N�!�.�1*�Z1ƍ\�QػR��^`�u��E@Z�,�\5$��Q��k���|5��h�sU<�T(�� �B�F�
V��>rnn�4���Q��c9ǘ6���7w.�L1g�%{���V��eS݇ ;lL�U�'��
��x�a"^�nn���)�i�&�a+e�R�
�ɲ�]��սc"�B��Y�v=��Uy+��N�n��c"�E�
��n=u�)-F%�qK��o�ZB��GZ2�;�x�%(�կar|)YJ��fmh,i��F�Uh���N��.�׏Z�`�;�����ʌ"B	
� �K4�=�!*&��n����v"h_İ^]M���:�OQ�{6N�5�a�1�Tq�)P�7`��{)�2��E���؆��)�
�I��3q�����p��y��C{7Y�f9�Z#^虅fA!:0k�Z�݋Ϧ�WOV�S�R��pI�� �̬Q�7O��u&S�w���&́֊xU�VUK8��6�#�S谚�q���\���+I�>O$+]�كBg5�r�Mj����?PŸ�2��`F��.�Q���ôO�~�w�=�Kȷ��M�aR�6Z"RZ��N���E��J��+FJ� ̛
�*���My` Ω�F���j���i=v(����T*�B�;ͥ:��/ �����cS$�إ�FVV�,Q���µY�<ÃHx�����·`؅�:����t��1�)L�FΫ۫�bd�NmVJ�/*4^���b^Mř��횥�~'L�V�%��L&�I�6�ٙCP0-��;�>��L�j�c��((34�5YOvbЉT�D"�Yt�����i�9n�>Y.�m���>nZ�E�өjY�Y��	G>�wGmKTf,��.�+�KsC��G(����U�aUjLC5�"��]���ѧZʪm�p��W)*��`�l�����n�SX�iǆ*�7�2���Cct�R���N�Sz*]^�⽄Уg(O�dvRx�Z��6T27qm`0��I�(f"f�w�W��.�����*b�`�u�h�e,F���Ԇ�mS���Va�1��PN�+.����l��k�p���-�"��#>�3^�F�)C&�V��K �Ė9a�\gp\��
�0�)e� ����.���xJ�,$u�v�+4�`5��^BF6�+Xr��B�ʶ-#��X�v�X��C]�Q���2����U�)^	.j(L��R䭠΢�������>N�Xi���u
�7z�*q)[��U]�E3V�l�X�Ƭ1��.�j����M�]fm�F�ؑ� �N^;�ЃN��&C�Zǵt��q-��ֶEUT����@��y�#6l��"�nA>�����%�.�\wb�mhxâ]�4]ƶ�e�&<�c�e��(!M�D�Ŏ�Mz0ZeL�Đ˭~b�"�9�R�t&��rٙ��NP��KYF���{q�7.�bM�����,:_!Z��&X�;&���<�u*�n���.5N��2�tT���Xh� �󅂺�e��rDk穲~�Zq[�n�)0��h,9N])qam�d��l���[�X�j���8vc�C�c%�$�#,b b�&�EP��G�w����� ���-��F�(����&�d�!U׶�Ԛ�]4N8o�e�[�ɚ,�b���g ��t�]����t�6�6h��м]ga{�/���@��B2'm�J��㕄�*�Ze��MV�}շS%י�*�������������T�58�K�e+��q|sR�P�7L�h��+��Yg�5X�jS�s;�ه���=������g��)�Wl[�[�ڰo��{9p�Hѽ��Nt |f�9ԫ)�f�O��Fd�DeJP���թ�w 3�P:�;���\%i�m�ުYaG[$��#-���s��`���"�]�zi��[�%�}co1�.��1���W"��.<�/���	�⼮�E���B�"��WK��PD�n�q�x\�J�>�p�z<[$n�Ю�� ����k�ؚ�iC�B�7x!��݄ýpVj�B�H��Q�Z�yE�t8Z���*�c����,��xP�a������z{�^�4*DY�u��x�!vu�z���;{[6g̊ǲ3�ٷy$f����f2\��\6���P*g���t�LF��46���������z��v�xF��N��&i�#F;���i}kI�������r=8��݁"c=#[����s%`�x���]=G8N��{�gǲːa���؛R�·�+���z]鿷֬��7ƍTev���켵ךn�� �A������1p�w�k4%�{d/\X;J�:��H�,74��,�_s刳�8uȻ��L�	KQ�9�UtӺ��$�V���z�;0k��
�*�J�$��:�V�}az�>=z��%�y�18"����=�)��U�oԞ���\��l�sj���m';p�6R��a�җ6}o���Lڼ�r�8�'��Tp�k �������`Ԙ}dPXJ�E�KIΤ��]Y�vl�t�8J;u-�������a�c���O���[�n�ޡ�1jT;x������*�8qJ�V�|��l�ݥu����-���3ռ�sZ���S
!=�{ySN��[�/J��dۍ�ؗp���U�|Y�w	l\����|�v�5�iKٖ��:plI��z�-�Y/�z�T@�ñ�[X�;n�Yè��p����u��m�!'*QV)n��$F�x�˷�q�x��J��]_Ƕ/�����+�H+7w��k�����ϲ�w_,�!f'�����5�Pb�t���걦��3�9s�ɝL����Ma��j'or��� u�#�՜�q��u���;��%���Ne�����i�ͳ��C��;1}��H&h=�O4�=�R�7eF����*��v�4<��o�D9V�o5�i��j
��X�t�b��J�X2G����w:	p��J�����U���w!4"��Uu�ζ��F������� �Z�����7������m��������ة>��m����YT����m�97]}x»[�����H�		���[ݝ��C�U��:���h��FABfB�ptFb�Ah��V�Y�a|��롛7�85'fK��3Na|jJ��f-r���;�6c�n9Z-Q6��R]Y��9\@b� (a�Zu^>˴v^T�&}N�;��a���Z���}&��z~�E�
��w5VԮ�+�A��'q�����c�ٜ,���l�P��y���7t�f�p�R��4�C��yj�7$�qZ�fC�B����Wnd��x�Qa�S���+z�y�%oݎ��:n7��N�*����C�0�p�U���<�`���/`�b�Q�y.�Pn��9��[۱w�o/iwv�mSH���kP����S=V�]*S��I8�ɸ�Y�]0 �]���Į���r���4n�uN�	�GƗn�^暚m𹝺�;]���nD貦j�{g �-��zu���o$+Odg�ۘv�:'�L�ݒ@()�¦���U؆��)	���{����1�=��ۇ��N�V%rry(#X�G@��ZHn�*={l*��v��������2]om�Ch�W�I��Ucgemw91u�k8��dHL���7j��t�������Wi�e���`Q��Op���;dg �T���[y5K�ջ|M�XLvņ�&�":�9����f�I�E�s]����M�Η֪X�x� 
�gV��5a8u�
���eXʵ�UƓ��؝��b>97��!�$��0��-"ip�8�e��0@z�}(���ۜ�?��N[�r[J�Ҫ۴r��ꄌ������u�9s�(;�Hمnq��{�&Lwy��%��I�V&�գ��w2t�N�K5'6湛��ifm{s�|��j��_t�֜<y/�
k�Ǖ�!��%N�+�6^t�j�����=�E#O�������5�4�H�+�pU,��G.f3�����VvC+q���)��'��C�-p�;�p��ŕ�����n.]�Wf�v�ĸA�8b}$��;e��;h�k:6�s�h�Q��]�Cr��-�]�c�YJ�e�HF{v5���`w��]�FWo�e��<��VCu[ܩ��3`�G;C�u�dP۸V�5�w7���D3t�ax8�7��nvT��QK�Zxqd����ݰ��m���@�tUr�%�0Y�Eqw�iAMN�"�֮�v�� »��˻����(�[h�w6���HfE�~�E��㢣BD�S|���_=�:���%5�L��a�G�\@4�����(nU���Δ�1q�u�U! Z�����Ek*J��9g�*Z��`�J�˚���f�I<�E.7.o̼�5��V-���~�J�wu��Iw+���
�C��{��3.1��3;�nsvd�|a�iUٛ�)���3z֪c{��S��I��T��1R}9���`��� �
��v�5û���s"����C������hU�6�f�#���U���|�E�����w�e����F
;��x�@�*ѹ$V��c���}��bE
8&�K��x��a�Udȫ��oJ�c� wZ�˼=�<T��Fnv9�w:㪣u�q���sIkCV�C�;(��f_&7��)�^>=$�7��De��}z�af��!�0�Tn$��{�RS\DO5���}&���ژe��b�9�Vh9n�[[�f\��|V·�u� ]׳��������]���Pڈfᝲ�;�%��s̭��f�f��g;1�P�݇��%ꒈ:o�����bN���fx�Av�=w�m:be�k�CH~�UfI5�삢��D@�L�4D�r^��?�����c�j~�~�%m��s�ٖ�{v�!��b;iV����aqًhZPwֳy���,����;W.�9z"�#s��S�������eL&�����9�y�ȝk[��ͭ��>�(���xt�Y;{F����;��R�<�:�q����1��o�:m��j�qoe�X�]�"Ņ��V�[R�V�f�h�u�r�����^�YkFs����0�S+W�;Nu��P9"5�(��@�``u��u�[i��&:(�Я <��Y�٠eH�>�4��铞�oYyu���#C8�Y܈1�d��Ҭ�!�is�s��s�f��\�)bކ.zAׂ@���n�4��r�o7��c�c�zpԳ)�ڰ�V\����MS��/l�ـ�7�L�	vz�X��sv�d�:8��|���F�X���-��q��;��ֆ�uJ+3l��>�S�v��0+�R4�δ��Uv�4%�RK"��9�@�|w���dXNF�@��C���W�RDr���tQX3�Ѽ��Bj	&_n���9��VI�Μ�Ư+3ޮ}"�\2��O���f�vY����Ï��kr�U�bZ,E��3\jڻ�w��5v��c(��0lW]R�4"op�">�X��{�Vɧ�]��@����&X�;��yQ�ٖ<��K�͙D�]y�ft��Q�F���Z_Lx�nör,s{4�ʺ��H��bFYzg-#C�Ҍۛ�i�IWv�wW�7����uWDb�J���z�c�t.���Ib�)n�r�$O�gsB�B�yغ7݂Z	o �a���1W��U�W6�wKc�G�]�����/7C���Vȭ��;S�52NƧv�cʛ-���;���:��\��-+zN[o"|�{Y�`�6��A��}���<��؞���7pѣl���o^.w=r��<̤�<�Ҋ�ڑ9:g��6�_Y��E�@:6+4�omb���8�GmbE�5|�j:Hu�C8�1=ɔ_Ɲ�\����9����K���7��R����m���!TR6�f\��0�y�[�C,�q��,�=�g;j�Zema�	<�Z]#�Gem>�.��v�
S΋��rΛƟC��I5��Y�s�]t%RnL�Ե���N&:����ˈ?��k�4Q��w��N@TZ��X�	�&�J�٭�FU/���wH*�m�H��5��Ы�Ɉ��͂�x��M�r�eM�O� ��H˖����׸����8���؎��W���2�5I����0�9��o�<}8����ImH�/um�IQ��ђ���r�<�hn��.��i��cE��u�z9�Ҕ�Y���O��Q��{{������ܡ7���3��qZ��h_m�b��3=s��'g=�|��ʬs=8dj�٪��T1�	i0���75et-ryD��b�:M��+\<��������r�� -�M�gj���:����g;��j�B�e���N�#;� �)�����^���l`�IosV�d�[�Yd�e�6��:���c��ڨ���v�Q���q���4鵎��:U���A�#:��
�Bnt/��w���$�]q�
(�8����u0Y��[���!u�Q�;���|w]�+>9O��w��b�лu�	uu��.Hk<�턜���[9v)�7r����z���,��י�@����w���z�b��4��f�1�M�ޢ4^��������#M�7�qN�a�4����4�4v��Ո��ܼ�g�Zӷ7\��u�D^#(�%��L�i*chͫ�ü2ov�]���Cw��b��#�:�t��js���44Q�������N�3W�u���-�vN0q�,�����ecG�:��X̾�]����t���ۦ����S�ăJ*�X�A,��t
�f#����}zm��uk�W�lE��c����UM=��գ^�{G;v�y���8���4�<�ALe�Sf��.���JvWC��k�%�S7n�AV��3��i��b��J�L��H��f���]���Z�[C!]r�`�+C*�m�����5}�y\;��7w�)7���́�4�e��vуx��w��Zf�i�]X��TV��˱bo��k�Ï
��������t�HU���3z]��\fA�E�9\�g��o�R�ѷԊ�O�L��L3]�x�M��v��g�	7M�]����q!�ɫ�G��b��+e�X����䶳tgs���ܢ�k�j��W��ot�
�s���/�%B�J���U��螝�O!1^�j�lp!R۹��:���b�vj�$Zm݃����'E;9Y��ef3��ۗ��d�#��u yD��y��;gU;={�6�V�Շ�G�Q�{��*pٰ.��]?̸gՙ�^Nܝ��rkv1���L�6���ot�W��q��]�����ˮ��5��/>;J��L�6q|V�e_l�Bs����p�B��y�Z#�*�v�^�:�Y�p.�񽽠Y[��2E���.=R'�Kn�$����N@�{�&G B	H]�p��k�q����f���bb��f�L����aX�,⪙*c��ȃ8���d��8�,p]�\3��`��޶r�3f���K��P��I*��mhXu�I]����4A�)�:�ga\%[wR0��99������6Գ/3㯣}�N��=���G�s��쫽���FO���^�8%����˘����҆%��o��8v���}-h7<vl[��)Q��N=Q���S���ynX�Wº9V�v�h���(:���kY�K��^Z s�]^����qˌa�*Y1ퟡU������TuHe����t�5���2[J�%�S�Y��k����^��LGos�ɤ/#��􃴚�\t�D<�ؘԓ ��`��X��'R����T�|��ސT�a�f<cr�%x���S<�W\�!aoC	���@E�EVMp2Y��t�j�ق�^����γ��8�f�)mt|�����c�Ռ7nV�-��v�\�_�2w�l�|��=�\锦c���+���>����������i�c�H3�_c�#R\����,�Y.��pp�����Ҧ�lXc�/�!qm���K�",�U:��K:�z*+����(h굛ʂ�e0b��u�	���r����V���,����9��N���]wx)T3�qt�C+6�Oq_eg^�U����V���z��{�a$uC��]�={	���?p�@$����&H?=�=�~�`w�?U����˝���Iۯ�Ҵ������7B�
����s���*���M��X�7t��IhC1"��y4�;p��J.���`Oe���r�L�Ybdܜ�FVl��,��I'V&3Qe���ڒ>·-��2����x���X�+"�s��`�Ɓ�%Bn�����v��2�v8��K��!������0Ӣ;�l@��Ә�o	K��;����ܸ��{�����GGNP�`ZN�b�:��wJ��P��\1��}D&�0/��X�dCP������#�u��YoU���s3�뷕�L��z�+xJ!Q���d]K�)Z��՗f���Ӻt1-J��hVkj���rb�6y��������[�r�7�ǎ݊�I;�H���k�Γl�����2ƻf����o�/�<�4�����FF7���[lՅ���-��(]4��k*ɉD���t�	l�����j�驪)m�Qբȸ�(��5&�*�r�34�MEX��b�EU�t�=YQV.���H��,��%EF�Xb�����őb3,.\\�Fڠ"Ĩ��Ҍ�ީ�Y`֤Q�*uJ̵4��,��/YE��`��� �V-LB�b���c*�$�<?Oy����������wv�:��Ȍ}�ų`�.�5D�K���_f�{���i�:�ܹ��=7�޲m}tRl I5pY����{-�H�H������3TN7��`6�܋�t ,ɸx�켾�&�zTv��<�n@�h$Y�ki8�Zv;h 6zk:����o��j�$��x��<�dH-H{�׹5�4�p�t�r��Q5��2�fk���a�����:�}�u=˳�+^`�]q���;�N�v�\nE�1���A}ٍ!�4��G�7h��;�4Vt��`�qR��s�h��/m����f��y��W9Wv�&�W0���s&��d[�x�(|dbvT=�].�}�op���6�I�|0i���:����ٱ���]���£��M_2��EҾ���ȸܸaB��E�����Pױ�oMnC�2�;p�ݨs���3���|�����C,�����E@i
}���ڷ���9\�U:�-�+H�������9<���y;�پO�T2�a>S��|6W����|,ӯR�=�K#�쫾Ѹ0��R���l!�y�ˠܣ\��ɧr��3)�؀}�iWc�+P�q-���p{pR�h���F��]����Q�I�F�����4�	��a4bQ�u���V���9V��0'�Rބ�藶��MJ�Ѻ�b-S}�:&+]3��,�5��T���w��iۇ��*�6��<���������Ƌ�Tk!�n������7����y�)]ճ�f�/i��ިDL����當!?R���J��c�;��P�vl��㙎J�Lo�Qz�ٱ馳V|n�5�O^-\pͰEy����gn���3\�8�8f�;K�1.㧡��oK��'5�gn��Y�A��
<�~���>��k�"V�Ѻ��/fc�V�1o�n���|�N�0�S���`��Z���O%ꏞĕs�U8<�y���#��v&�|q_�Xoˢw+�vᾯ&W2\tK��g7��-�QS�dױ7�,���[�+֌��
�	��S{/�9\)�r�}� �x)�W7��q-ܬ��t,P���
�c�@���UۗZ�M�p	�$��q�+"��׆]a�V���0�H���f7�,�Oi�w��ل����r�%���X�Fq?\d��ͅ>p��� "y�ŚakY��|�i��t<z��ǳZ�����D�ŝ�p;ܸ�t��Hq�tI��]^�Q����S��'	28]�k����� �Q��(��@���x�BLX�ܩ�,DV�#P$�������(���+�ZZ޻�c�\\�	8�����z�A���B0宸줮z��Ӛ�\[q!�}���m�G�t.�^�F�k��x&�_v�֒���5Ŧ�o������
@
��3�(6�-����oe`��R�J��CNz���Æ���ZYo|N�����'���O��zd��]x����vk�o:�H-��6��_Y*"�\���^���hRo&A(�x�B�Z��of;;�fB��N�ˬ�r��]�
�w��8�j� s���	�6�q�'�Qnk�띅
3M�~л���Ep��]��9��-�{Jg,c��;_;)r�[Kg��9^vs���4�i�y�ZR�����R3J���y���vX�.W�ۛ�=���wO�ΪnM���3vNP�3���<Ǩ"h��p�f��[��;�x�[p��D�����窴���5��[����ʞ
�
�ɁZ��I�hz^��-���Gn�Z%9�c]�b���4o�\]������A�E���xm��U�̒/�����P+w_)�U��P�#��ķ��QF��N�0�n(��1I��>/s�������ů%9�(�ۛK��7Y�ELj��en幷1-�qi��O,�;���?[Y~z�0I�=��<|Y�kGĠ�f�U����n>{��c_lZ�6)��s���i��g_]� Y���c�4���l��i�fq�YE�5u�\`�,�t���O�@��}[�}���KsD4G���	�6TiN넞�_s�Nm�7$�o�z�Wm~�$Q.W������v�h�0��Vr��Ӱ	���zW��+"��@S6�!�=�-�:i�J�% �6E{'�^�Vs)E�����!y�IX��\{�)�h0�dk�׭T�͹�<z���-�-�{��򞚎����gq�S5j��y���.^����<�%�p�u�7�}\�s��	O||��œ��J����׬+�Ae�<�2�M����k:[J�ۮ���61�������$$��b��B��}���T�Ыi��'-���_ &Y��t��gU˽�/��yiI��j�1�yW9y�d󗭐���u{r>T;���t-cBʮ�Unޕ*4�Wb5��/C�T��A��޹�!Y��rW�P\��� ����.�QGC�JRo������깏��.����������~�qm��\�Q��l6RJ�:v9wEnXo+��W����(��d�]���:�)��mm��M��En7؇S������B�����)�?�x�2��g�[�����"fBjWa�C���|�*x!n�O�ۇ�]��t���3kί���L��`U�y`���V'0�����NL��u��iڶ_l2u�|1�ſf\�,ٳ���A�Wp����t�ܚ���nl��Noq-���w�re�>�lu�����<;�88�%LkY�p�p��6���k�B'Җd�,�����s��bo�~��40��*2K���7٩�-�L�]]�^�Fo����T	f�Sa���ⰲ������8:N��oV�
���.��F��u�.Y��u8��-fl"���CSb:�S �R��݋��k&��J�6�w&�ݝ�D�zkӇ�P���i�*of^]\N����dix~��z��<W�U1[fԲR��T�MT�5+��%`s$&yN]�l �X
�A��L�-�*��&9>��>4R�rJ�c,�nd�U�b���jʱ��Z�kĈb�0#�M�tPb�1XS�5G��*�T�*0~J�4�0EݙT��ud��ς�]�-3�����7U�+�c_G0%Zf|]3��Q�T5a�x���T]Q�SɅ�Ir�r�X��R�PiEn�#�t�Q*�F�e�q�x��S>/��T�uM�4�ǌa�D�S�UB���$����aX�b[�h��2&L�
��[�X�+3�� �[�Z�~��Z�i�Z�T`�Q-�Q���Z��#Z�J�Ŋd���m
�b���UA\e�H(�b
�TVУ��Q�.S�TulU`� ��,��m������V$ĔEU�T1*�,UB���"EE �1Z�(��`��T�lPS,�c!Z���TR۹�g����\�}vk:�]�A��w��P�XI}&�<��Jڸ��RoS$1jﵔ�T�p��e���*�	�A-���Gē�Ҟ��5��]1�&���ѥ����D�v1u���<��W�3�������~�wo ب B��PS�氮��<�z_U{~���e���X��iy��F+W�5Z���ذ��-o���;%�Ou���T>P@�q�R��8���ʻuӨ}'G�;<�V�_yE��S˚kS�cr���ǆT�WW�71�ta��p�O�\2��}�kf��"��b=�*�u�gve}r��mK�p	{�|s+ڗ�졜�V�Z�*�ū�}�^@W@���T���J��o`R��!�����wے�6#��8!�;�x���5��~z���u�p� ���t�.���y�Ͳߩpd=���׹	w���#�+���y�9�%��7]�ώ���ٹhÉq���J���=8z��a�����xo�W���
�)����NN:��|�}o3]k��W���^~$N���j��E�\�k���Wu̩*@�9�L�7�Kp���xOp�J0�NX���\�\-�w\}[S�t����w�s�y��wy��6�;Ձ�M�q �'Bą���L�@S��ջ��%՟f����T�G���z:b=p���0�$=N�z�q�����R\��c���<���޷���І3��|�f�6�=Ad�aā�@8�˼�0:f$=a�C�M�C���������HCԓ��RN�m�<a�"�m���|��i�H_i� q�%�ϻ����ξ�|$�C�HAd�����!�a݆$����$�N��q$P-���߆^�zn��m�zr��$�@Y!�,�@�L'��m��v��N'I�w��6�����=`�2!=I��|�pI�N�ë|��a}͝o�k�o�I�P���Mr��l�=��9gI�@�$�������Ւ��E$>���]Ryw�~:������Ӫjɳ9I�nV���;U�yM���ֈ���Te)L)(Nw6Q�EX3'���<�c{����O�����$��Y� i�MNP�2��L&�I�&n��I:w�w��w�����U�z��q |�t��3��;`��wC�v�4yd;d3��`wLaY�N�:a��&}�y�k�'�$82t���!�'hM!�]Ӧ��0����L��x��	�q��5�u�sߠx�{��;dY!֨C�H�'ēl��VHS�t��[��^����}��r$�����6ȲgvI�L9I<`V O���C��Cה�h￳�m��ί�|�C��	�O�k�a!�6Ȱ���i&��� m�vH)l��bI&���z׽��I�B��'i<@�����xã�8�3VI6���N$;I���1�9���o�k�}���'l�$>�=d;`k�'̇��8¥B�̞!06�THc�}y�o�y�$1��$�;H��)6�;G�2c!�"����@8�ݧ�8�3��z~����ONXx�t�J�ORv�VI4���Y!��,���P8�gԁ�}��}��w�s{�~����.�ę�ۧU��yCGK5�p��=FЏ�yw�+���Q���CA\�+(4z���މA��=�_}_��Bt_���!��%�� _�I�oHC仡����_=9��������Ϥ=I�FIP�$5�<C�_R��yAI<BLI�l�������&��o[���~�:H��@�1��'�hf�"����8��8�v}d���$Ω>@3����oׯ}��1�N��XB��8ɶ���|���M2��$6�g�&!���� �'�u���������i"�=@�ߨC�v�2_Xx�<{Hq w��OLHz��#ֹ���=������t�����O�I�O�!�Ci�}��$�yBq��i6�q�_�w�:��o������x�t��$�%dP��$6�遣�q;zd�d�$s6}��ϯ]����N'��d��6��!�6�i&�@:d��CYa�=a�Hq���Nw���^o��$7�g�'�d�,��8��j��I��:d�$��M 6u���w��!�I��C��$��B�;7d;d�!� vu�I<�0�s�
��-�q�ը��K�z�6m��r�+��x�m�nΣZ�>eK~�V��+�����[��wT�͑[�5�:�04�S��-��1�������rv�!3�I� �$��$;-���o���6�8���"�kVl&y�;�����=��4���Hz�$���O�I��&�$.�>`v����q	R���1�������g���>�F}�@� @�	�!~�t�v��_d!P�|��"��:�4C�0�:�'z�<`t�w>��!�$&0�v�T	�=MRv�=�9�������T��0<�����+�u�>���)�6�����xy�&�#�\�l�"���V��v�ޭ�t�ЍaGN�żx_$U9;�ƍ4��J:�dEaW�C4xF8�3��kB�ɍiU��N�ѫ���Q�oT>�I�m	�gdX_CF���ӕ�2�+j��:��\��a�c�o�4�d�7�W�E}9.�qN�o{�Ü��Gno��ӓ�kKV�i���m��Z�O���t�����i4���M�i8T��j��2��M��+"�<����?Q���gn�c+ގ�ں��Ydh򻛜������,���5=J{�7��W�!����-� �{#�)�S/�y���8�&F�$\�=�>�o��:�Rsk���㷢�ί�!&B���%���>�P����2�Gб�Тf��J��p�`qz�9DFT�ܴ�����e9=Sz�=���t47�Yի��������2v�8'{9��2��<Y���ȫ{�`��=w|�f���Sqy�d#ʮ0!����KF;��-�h�ܵ�w"H��j6�$2sj�tl�+��ךS8X�����tz-~��
T톺�dI������)���v����Ϫ*ѕ�(h�&<�V��̮���8�nLN���l0VYZK��竅>����AF,ʷ$�x�j=��gws&#��f⛳�S<x|�#�'���{&;����iY�^?�_��_�_�*��2��kQ�(/U�K�%޻�rxt�y��-����͛�/pOS}�x.��cd�[���ې���^�\�;�w��ҹWk��W[K7[m�")��g���Q��	������-��k�ģ��.{���1U�76�����K
��^N�ɓZ�R����f�t<ݧ4EN��ۓl�ly�Fn��!���ݹ�g���W�h�a���9�n	jMÂv�1[O�zz䭤1wVH���BWn%�(��y��ZS��S���?���=�Ы���uK`�#��b2���g�4���uy[
���t1m��T,�����8�y��"ӣG�K��6qGت�Q��>^o�eg3�;��j�tt�9.��q���p�����J>��M�W�p�׶�I�p���*	�y�� �J�ق��E���f�੖�D��w�ؽup�\$�j�s��f ~��^�Ċ��ϠL��T%���U�5�`;<ۛ��u����z]NsH)A5z��u-0D[r��t��9w�t��Z<'0��e�[6 �� I��`�QV�v+�1�M�Y�t�[��*��;�;������� �u&\�ΎX�t�w�{!���×��Tۢ���:'�bʼEI���s�m�^�wA��D��Sm�/�$�z�_E�6Z2�^|�-�'k1ꩲnO')��0U��/4��i�iP<���M1��L�$r��.���n�s��<lr�UD���k|� ��^^q�;�K׃/՘/N��of��)Z�t�>���U��쫵k5����T���V�Oo�=�,�Fj���	p��U(�:E7T�ϭ��X��9J�-A1�5$V\#2�X.�U]%L�o �ј�ݘ(C%�^aU���MT�BM-�R�V*��pI^���+);VBTqT*�"�Jd���VEZhRE 須7F�����o]������%�e�Ìi��SM�HѢ�.$��jfQ�bn���7T�`&�XkZ7x��G��T"~֡��-C&dsj��AnJU82Xm$�t��*S�7XA��0�-݋����r嶜WR^��9�U�l�Ia
$�	�YYDГ*���,Fpc"�T �j�~a��;D��Z�V�Se��}g���~:{a� T]J
#Z�m���Z��(��XT�%T�J��Ձ�E����+1�V
�F�i�Z&����£iQmim�X�fc-D�*e��J%*7FT���խ�F�*�ӆ6��
%��,Kj�--*(Vk�-՘�#��ˌ��C
�#U���Q�U`[a�ㆵ�o�~�ʦ�ۮ�W��NcE�+A鉽vb��x����}T�֧�h���ւ���Q�˺��O#{���uk���3�����tA���Bf�v4�G��%ܗzż"�̱�-�Q���=ȧo�Ob�|�g]>��ʁ�^5Vq�Kh�f��a�9�n��Z�^18ťsM�+��唶�[dG+ը���t�<������s/�Qȧ8m۞8������8d1y�pf�����H���|���C(qc��\e�m�zY�&�x� ���3H��2���H�Ig�N����/���W�9vz�]�5~�b��ghwS9��E�GL���UODM9+4����<�}Q�`��'��M�x�1&	6y�.+��-�%te��A.�8�c\�#�L�y�SM�w5eƋ�e��z�3#�i�R�ꮀd��ܣӅ��Z�6�ձ�j<U������}��>����\�ު�7�
~�z�3�E��ުfj}����MBjQ_�gP����3e�F�T��Y��vIr��uhx��|��.���c����p����v�'�j�>VdFg2�,	9Ǐ��D`��y>��v�=;�W��}�jK�ig��^��f)����2��S��{{Qe;`�f��[�F{K��Y�n��⏍�#�=[	��B�JX[C0o�q�q�\Ezýa�|��cK\XI(5�j�⽷=��=���"�.$�������Ib/pE�lz�{=�G�N������-�.<�����?f�����f�$`��������^��>�!�C�)��1�5�tg�>͐�h��Q2����D�� ��QVX�N�@�����m"yb�'-0��>s']�y5W(���'`��ZYa��L�'e:@c�-k��(�L3x���｣�[�ו�u��Of~{��D-8���Bt�?Ev�����E��� ��52ɜix�r�R�<a���Vzb�դi��B�qf�+kx�><Q�g�*�ЏJ�*!`mu�����J�c-��v�a��DPd��9�];�z�eĦ�r=���<�;_�!3>�1�H^Aj��s�e×�*����S�]��Q�P;w�ڼ�vs�P#K#u{��9���͌_޷㶂7���,���?x��U�p�ٗ+�6Fk�OG��-:Fj�X�Cܰ�|�Z�rno�Y�Xx4>hi���u�����O1�^&<�n��������tp�3��]���I�3��un>̝�<�a+��)A̨0`T�1E�Ňm���X�n��ݙφk���jyZH2Y$���%+�"#���z�|=�5<#�jȅ�#�
���n�sIv��=x�ڵ*vf�s>�\v'����/�Ee�!�W��{X�U�q��鐄�Jg����7.zK���V';�]M?i� s9�i��C��t�#�&#6��V�1�'L:p����>8Y�V٨�e轤n:��c�7��g����,�PͧgS�e���e��}�x����܅��x�8NSbޚ4�!\�Ks��4׆�9<�k����b�"�<zX��l�;��8h����[�d=V3��%�fP��A�M�r�'�},��<��9	j�ߦS��5cX��[T�����QS�e��b����E��,G*Ħ�uc�����K]������t��X��̬ݻ��w����ݽ�,��5�xѨ��ˁ��g��Wc���n����i�y�-\�@ӹ���(*_ː|�=�c'�'y�����;v1Q��E�ǦXF���;g��i���G��Ok��k��ld;X��!�.�������M���_dY��N���B�H)�Ο��Β<w���H��NcvR�з!�!��������'�#I��o��������v�D�GhsŠ�|o�9j�cw������Qx��DC�<�f6S�9�:�w��᨞|�+�P
5�?9�r��O5YP1w7��G5�ӹu�U���x�C������*=.c�rq7V܈rf���2����;��s�;�UW�U�[���n�)���-��������c��_!�l��ֲMF���ϱq�_O&t� ���#_z;:��R��up�@��ő���x��C�#�eg�&�	���5�x��vZ� T̿����f�4T�_1Ps�:v/l��,���V_��$x��:�p馎�ԼΔ�R\��Sr�ҵj	�y���- $����i�^�ܬ��{�M�����b�����º�>�R|���_pQ���L�Vr|����{�>�8X+�eZ�wV8�_3޶�b�\��ҹq`�%�t�(r��|��8���(�T���g�ku$��y��$��7št�V��߶�T���Sw�X%���A[�iV���S�P����#�z�I]����J�;��lk��R P�N�I�6�q)U^#i%y����I	��s��_S��Y��̺�^�	�`�:��ۮssn��"��yaChA0�!�,!��c��0�{�H��8�CA���S�aFyc��2��]�GL։\��"p��1��YVt��Q�#ʯe��6����<i��B�c����O��\��Ƿ�y������Ə�U+9hCgu}�ԆMc��>��<�v�p�	�
>>6I��#���*y�;�}:��EWo�V��D{�)lA�	>>:p�}�鷪�Z��ߥ�<pΙ>���v�ȉ���G.��ޛy�@p�<9�C<����,W�Q���tT�y?6S��/�p=f�p�:�R�9�����z��P��dvG�U}_}�^BߣW�����!SG�B��g�����mU��&V�Y�`�7���Z�#Xx�Ѩf��&!�EQ��I?3QQ�h#����L�g��+U�ӟn��+/k�L6���;9A ���n�śj���>�NMl�u%�~�K�i��)QG4+許h�P�+d/�5�}D�gָ�.!|���WA��:d��l�Х�"r~����1�yq:�r��|h�!,W��u�g|��ւ���K#�^����C���k9���/|t��)@'��f�x�X��@c�Z�S�|��P��x|�����o��%�j����~�]k�L�a�<{�v��J�(�I.Sf�&�St��cfn`��r�Z�;��7���\�#ޏ{�l_k�~5�ك��MJ��1�F`���3x!�ԅ�V���0�%C��N)j�Nb��C�HC��Ogvy�+�<r������p��qQ���Տ�	Ƴ�{_�\�7 릩�o<��W��)H�V��Nڍ��G��>��C���u����Ӳf�è�q4�]��g_{�Æ��s����VB#Zd��1�Q�y%w�o���U�j4x�!�t&b�GM������>D`�ܙyDB�7��o�Qh!�;3�/��ZG5���m�ٞ��Օd{�4l���:@&R�-6F��}}왣��Ha�r��v�^"[��{�JN^b��g�j�o*]����	�P�q�P�"4���h^+� H�䷅ɺ�$w-n���ʆS�0�y���eBM�	k-���X�Z}�wd��S ���`��y;�ja�;+s�����{m��B���+ݒ4r�[���5�(�Eߊ�E�[箮f�@���3�4s�^Sꂚ*{�y���U}�M�;��̲�,v'vf����粷�B�i68�d��!��Z.)�j�8�9V5WR,!���1	B�,��w�j�_
ˏ�5*;n���w�����Y1��г�kr��Mp��UC�z�uM<J�}��^u)�)ɤ�5�V1ͤ��X�%�T��"�Ҙ�}���j�#Nև��\��CƂ�U��$�n�2�"˰��<F��	{y�2Y�C�]ea�D}nA�Wh4!���-�x]�>y3#S:WeԳ1��L���Lm��h�T��HeXi�N^�I0r��i��(�i��و�a��30�A��Ԫ�n�
m��m�@�^c5�*�J.�Y9vq��H������o�c_%I��[�$�0�i���t�
G]X�UWL˴n��&�������CP��k'a�`UWm�P��-�v�QOoH��,�P&�����u��C�3�ֵ�-��*�\``���U�[Q���(�Mj��������,PS5epm�acE�e(֮�sY��-J(�ҍ�V"��b��c�K�XdQ+b�HW-��`��(��"--U[j���E+*Z�+()h�UQm-lTmR�֕����%�(�[R�ι�u���E�@v���O�(�vݍ�$�yC��J����� z�no�~��Z���Q�q
����K���Ү����{޹p���+?,C&�Q�Cډ�x��c��ے�U{Ț�T�>$�Za�$x�\B���{"*���`پ����߰ٶ�5���>"����ۈդG��zg���[�.U��g��;�{�/�H��0�f�ӧ�^�G�|A��9�25i�K0����w�ig��r^��rӶ�E��Z���f^4v �7/����#�0�5��v㛞�+�'ۊ�e�ZQ$x��E����h~�X��[;���MC�W]+�+�44�Z@J��l����>tb����I��S�*��
�Ita�Y�<�L�\0r�̮,v��M�W,���F_v��'_4�acop�[@�m�5+g`�e7�;*9 ����������y�Wlδ�uW���f' ��$@�x:i�c��:�iu��2#��V|�8l�FLd����K�޽u������Dȇ|��֭��8�#I4�pY����F����6."�STEe�Y���
��6z���C�Q�����Θv���`����mZ~���{V��a�8�Y|��
(���vG����4�����/�cI�7J��D8E��$�f�gk�t'܈���d˔�dʘMu�fΒ^���ûݙ�4�Q��<����*+;��O�	��]fuf�Â�t�Y
�g�G�i|��0:sa�_��+;z��ő�e�/$�ù]>�ݗL*��.�����=�nw4�>��9��Y�	.�ЏV1u�m��]�7����\CŔ�������"�	�����z#���d-銞�2��6HC�n\��t���y}�}G�7`|o�C5o�CiYun�(y1�m���̈́-Sɑ�7�=vŎ��h[������d�U[=^ݯ��(�#0ࣽ��\�84̧����}�Fq�C�|�t��(���O2��~�%��g٬몭u���k�d���G)C8^���Ҳ3ٙn��VVJ�͍��H�i�*"#����4���OИ���8��%�_1���\j�?���*�O"�8q�]&K�S��Jn��`��=9�'%�ܾ�b�_^��0�9����ͬ��FZ�Ի��j��{����sݕ���kO�E�ZO�1Ǐ�q���5p�̻�$4|�����c'�#A���yW���6G�O(LL��r�	�.*؊5��O�x�Z���d��!����x�Ms���fvw���<6���u�M5i~B�xG��f]��7QJY��v~� ʞ| �1Q�B7|��BȾ��D�|U�6oP�!E���Bj�b�⋈Y�N�K'����O�!x������-u�r�����������c��p�Ȫ2'��ښX~��y��0����<�gm���f�#<��Bڣ�Y�R��c��J;��TA��6�=�ۼkldʚg6n��vf�Y�d!U�K�6.u�U>��;��ּ�#=�l�p5owo}�G�ޅZ�<sj>�W�|�6L���s7���,(�k
�X��:���*!�o���_h"�Ό����|N��ss�ȣ{�ZC����,F1���y���^:l�����$�YGi|���HA�xlӥ����WJ����z���zl���do)�0~�!@���q��׵�����G�,p�\���?,C&�Q�A�D���"��j`Jk� ʜ����:��13.NCz�gQƓ/f�]�Ĝ�	�lg����[�3�@��3Ϊa�S��|!�@��J�W���'/�9���-��C��:��j�?�ç�����p;���]�ȹ�)T�m����d��2������Fn��n��r(xAj_,���e�]�/Q`�E�kʫ�*�����.P�m뱮��)�8,�r�x̤����w� w�ם��Ǽ�q����v�����˄Wh(毹�:�ve'�;��v�D&� 	�O�?e��{y'�V̓��F���s|�f�S������Vaq��hQƴ���x��im��Giy ���W]-���TVv/�1���&�љ�q�l震Ǟ限���<l�P�A��4͑g���P!=��r����uu�0�q�
�1x�%|��_�:Ifh{]�A����-S$(g������w���Y�Q}Vx�� מ��3�iy[�_��U�ڬ49������x��E��(���d�~���:t}�7�M��{z��v2=T6l�6�լ�����玆��8��zC���~��=�8Ż6׈��hda�*��-`�=��>=ȝ<GmA��9�Լ�u�ymx�G5a�
#5���b%��_|�V����{�T@�K��X,��=Nzzc�RIj�up5��D߼�񲎑��?2=��Q�)lt��=�~f5�B�8t�b�^�"0��H��oG�6�ۓvm����c�i�F�����fZ�#�ռ�e���!������^���Z���Lٳf�kOϪ���=��D8�!e#t_���;G"��������s�wf��}o��1���E<�8����3Q���g�����V�-��sj����3��j6U</XMv:P�R�6�/�6�if���)�6����v馊���^>?������ni��B�$�j+?����C�Zk4B���7;����udL�����d�����P�'{�ڼ{S4o���1�y�K5B!�9��I�W�8�����/<<p�ֈ�~��6��qq���Hw���kǩL��T<��螙� ���X�l��Oݙ��ֽ�M��Bs�a��n$���)����d-���=�1�`�/�� �4x���&/<t>ĳ.������~�D��C�q�^8E��o�N�z
�b����;5��m�"�xG�ުX;]T՝�e�����ў���÷�Q`� �|��6e����Տ"�f���n�)�%�>\�s��Ϋ��`�Q[����7�_w,�%���ݎ��Ǻ3Vl��'�&���K�� ���s�����J_��6]�"�L����]]��5x.�s��6s��²8�W��ǥ�]kM�>�-���	�5i�b�(�d�N��q���6�%�1�F�{�{֘j͚#׮��̈́h�+!�20�Z�������'��y<�x�r�3�a3)imQ"�e�ت�<��ʆ�g�� �Z�x��s$>T_��v?�[���h�֘q��;l0h���$p�����F�*����Dx���d���هǋ����a��f߻���u��$8��1Vk��,A�52���2��[S픩���5���>x�NPTy���+=9I�|�ً�IL�"�z�C��e�Ta���8���<!n��� �A�U1e�s�EOJ"��m�_G���Nu�]�&�O�Ww��M�+��:|v�u}qUr�x.��rg�AD�H��S�8��}����!�|���ǲv]��t��H�g>0u=0y����B1ι{|U��xDq�3�0�ј������V�Y}���'��k���"`��V��|#��]F�x�����i��&hᣖ�4M���O����n����_����������-C�����D���M���|��9��]p��^\GDJTs�mpH(��Ao6Z������,�?���1/�+4X�a�Z�2���vT��<0�k�!z���b��t+^]���C9z�/�¢kt�mܞ��[�J�u����|iR٫޼��Iv(�TЪ��[FJ��']CJ���6�fV�қ����j �d�΄- ��(5g�J�+\���˲�68�������̒Ըn�׮�=�A�]�RO���Ԗ���)7��m�!O9B�ej����SWa��nr8ƲA-��]�ʒ��h�w��+뒴��.2��zF�V�ttɑ�r9��Mg0�]��O��A]���2��:oEML=\�<o6)h�_�1Ӱfv�Z�30�K|�P7�x�տ4��e��I��F�2:�h�H��&�)��d�c��C��C�HmJ;X�ř3���Ȝs��3r�/F�ED2�Z�4�֭�b�Pkˠ��[����*	I��?ab^h[��o^��Me�$�h��م�.1LIٱ�\���ww:��S+o����x��#9lfZ����V
�i�s]XЦ�8�9\m�*��5��rC}��
�X��9Z�n����:�v���G��9�E�74V1� ��u��oNw��.g-�隶�]�qq�������{-NP�5ѽ�fR��a`�n���{�V&��6kk�s�.�`�Ղ��N�mJKl�am 1*��Sr� ����3x��u���}�zs	��
�W8޴��ݑ��n3I�j�!�N��,�<d�x7����a�9麳u�d8��F�ؙ�Ӯ3�)��D���d���}ww��P J�T��J ֭q�-�Q���9pʕ�@�Im��+
�*��Ɗ�-�V�5*��*Z��ܸ���إ*��֫Z"��P��Q�b-����W��"[J����h-+*���-QFE����YR���ei-�%�Q����E��e�Kj6��-�̱F�i��-���J���J�Z%(Ҩ�!mF�ֱ)iR����F�V��(25�u߽�=��7n�r�r�l���H��uf����΄���k|>��,���Y��C�����B!B~dA7�v1�q
T����~0�Q,�f�����9��x��b�!DY�}Yp�z��ې�ه��P6��1��p��8hj�:b�:�^z��>zD:��$8b�C���qp�����R��Yw���d�?q��Xƃmx����v�����C؁/��x�xçym1�wu��̥��^-�Z|Y���>c1Fy���2���ЕHf���	/>?X**>!��#����>uݱ�ZY���_5�a&�����O�g��&.?Q�1
`s���"�AgF"_ݛ����3�(����U8���Čؼݑܼ)D^�5"�o�Yl{��js�cC���CӹE҄����g
9Z��"��&~�����W�Ų�W�A����X {�}>2;a�z&T��h�Do��ywD�;lUqީ�l���v��mN��pds��*_�R��>[��w��;�SP�^�j��w����O�E*b�,�^"5��I�ԗ�䗗�F�^1X��Y'��<-����Y�n�Z��nv�PK����ݓ	-��P�9�r�J��z��w�~bX���eOL��(%F��������9�;��-/P'�XZ��XO��|�<*pW��ZR`K��q�}�^�t�j�����Z�ǘü������{{�Y�l����B���GR���7����@ߤ�
��v�'�'{�v&�=��j�ݠ���Ȏ��g�x�`�������}���IV/�������4G�a�Q��E����<�~�̇����y�-�&�� �k������.ܺ�FGZ
��	�xx�v�9���d3�+s�Ǔ����E�o1���Y�y}�,�)���J���],��J8V�:e�����z��(Y��4�3�����<�
pK�����Z�0ܵt{�)���iU�&�9�,��>�0ѯ���d�Z�F;�K<a���j���j�n�>H"0�,�Q�nX���}\�r�;b��M"b%}j�ZQ�0��+wݿpjHFŔU�7<�8����uծ�u�ʿ2�`)�������gYr�%�ۆ��N�����gq�9����.�m��$:qG6^{ԫ�}U�|FF�{�,���t�iIӄ^y�/���i/�O�a����|l��}�ȢH���^,�:i�2
�2xX�H��.�~_YT�%���x��iM+:@���!�A0�������W���u��K���y���0�iT^0Ѳ	'=�V*�Uuz��b��$
��S�7�lBȣ��=^�>Ea�Ø��6�㽯
��j��PWj�-���_+���4��,�޿M4~>Tt�sym���;+z� ���Ix��xٚ�Vsįs3�Xa�<�Z�Fz�mh�'���\qyU�}짫5<�qJ8�*"S�HgQ�8�a�*�z�;t�(tnک�ݮ�K�]t��8��u�\��z=�0�|���y�r��vFI��?_We�c5����z��~?�(�)���dO�ݘ1T�U���;0&��C��r��k�@�d��yV�*��z�*^�ϜVd٨RPQk�8h塄O�(o���oɍ�<Bl��%daZ��a��(�Lus��a>>*�"�Tl�40�]�G�cO�3�<t�G����,�q|�?(��� �_U���Ț��Zv6���B���&�|j���:Q��K�{�}JvT�+ Z7��À�繌4Gb�����9���p��+>�`A���߰���v^]�.WWN7��f�>82��'���VP� �����W�b��o�ԍ�'�=�%!����3�t��t��;T��u��i��|��{�1�SyV!��	|aN�^�>�n7�n����
0RU<��2�G52�QG�k���b�[�Q�8�j����,ãцz_�g�j�ĆxZ��o�7j���.|��:l���_���|G�$&�T}�
��Z��DG+�O�:�o�Nw���
}ۋ�쌗p?[>����Ob�����ZJ��־���&-�ٕޔm!��C�礘Ѕ�0�u�g���k�����?Y���r&2Cʌhd����($���ga�H��(�à$)K�v���4���{8���!3�8 $��
J�$wl�՛ݻ���Z!��Ö�{M}��#-~�&6֐�W�!F��d��b�_2mQ�\_��O޾ckr�����:L�xʑ;>�f�e�Fe�u���:����f?�]��� ��y�0����3\�����F�-�G��
(�����5����*��M���#�_f�x�C��A$��v�}��l>��P^^�2,69�	��ӧ�^�<��֏��8r�.���ϱűN�g� !vz���~�O��lC"$��ǇN����ƈx�g�t�}�(�G�_/�"{���],8-m�3�Gv��S��Ո������ť���id@���}��ū2Nn\_V	���]�3lGz�a]���lZ���>�~3kgm2&��pфk2�үj��8xE��v�6,+��0߀�����Ԧe���#G���Br�C�Ж3'ϫ!0��I��cό�˩G�gǈ~\E�-2�4m�
#��t�p��f�5y$לU)�*۫"��Ӓ1�c���^��j���g���}X�?9����^�ļ뼲J$��c'<.!"x����B��֯��
t�{;����<t�M�:@�L��
���W�^��?����ƾ#�Lk�D��{n{F���!���`,]�r'����E�Y����S[�r�{���`خ���t�=�t�M�bZ੻����0rYRR�<�[�5��ٝ|��Ӻ��ˌѮ[�ɛ߾����:��>��u-۶��mͭ��9��+n�����5W��-0@'�!�h�Lx�J�zf���U>#'�|5�_+-�����_VAWʓ�]�(�M�r������^�j��K}�9�=w�ެ6~�W��Ob�x�g�=kh�D�G՗��c��0�x�D4���j�BȲ[��H�a�ܿ���||^�#�3+m�Nġ|��Xk�/��1砢���Eb��v�gw�z	-�����Pᶾ�_i��F��^���T)n�c�f�L[�<�����G&�/�ʧ�3:u���I%���w��W^!�'xo��!�j�˝�v䏅iɼ��L��\����Ҿ��}�#�*\ܒ�6���#gL�p���:�~E7�{�;��P>#�cV�Hq�C��7;�=�M�WA�q���ܬ��1���Q�S&�,���l�0E8ꌗ1��$���A�=�����p���*�Y�{{�pި.���/���g��	�=�kv�2��������O)�h"���D�>K0yV��ه�k���thT��㬚�0��B|�ݗ�\�OG����%<!�欌��R��>�=G��HY�H��7B�ݞ�,Z��*|��2
�W��n]vn���P$����O0�.��5�ǖ�	�*o���<sľ�"�r����6ܘthE8jQ;ʅ��	u�W4SKf�s�M�-tר��Np���XjŻ�˘b	�cފc�kB7`ɖ��;�������pơ�����E9�͞{����A�O~/�oE�;h�)�ZA����d H�۔�o^*u_Rr���Nw����dQh2�V��U�}��s��.�µ^\�F�I2��S��ŗ �X��:�i�sj��53�u���m�B���j1�L2�ů9��	�3&�I�݄�s9[�i�C�$o���(���]���(�I8ý2m�����B�uy��ۭ���n9�x^ӗT��t��S��j>2-Mb�#N�p����t���"Su����5�W{!ZǓO�_�0v8��6�Z#3���2ڬ��)��
¶��1�J[��˲���f�޺Vg�n�/�®`�-Ǔʻ.J>�o7&�1F�n%H@��z���s��Ĳ��),ټ;�qs��
����6�bGՅ��k��j������y�E��m��ngu�os�:�
N@{l�k5�tVJ��E����:������k��c�&�k%t����-�X�/�F���^m,ľ��0�8��b�Que�t&���f�֤Vwŧ��7T��.'�>{Q�θ� ɜ��sh$K�''E�6��Z:Ji�V�����^MӁ3��P�8:y�D9u�n�m"�]ª�7.��%�����ř%rc�ye�;r�U�%��Z#m�*�*6��n�q
�
��b3-ʌ(��V�DUmhU���Q(�U�Z2bc��b�\����i�%Kj�l�*�����F�b���-�-e)\akk�0j�KFZPb��Qem�c�Q�ڊ4mTt�U�UQ���%�*��.[i*���2�Z�K�SU,�ш"#�Yu�b��QjJ+�]5QE�b֩���I��?z��[^ڌw�oU'FԬ{Ba�PV���R*~_Ԫ���۞���������P��:g�
6Fк�����C�/R�Qr�d�3�vL���G�K�i���꠩��4t��!�b�w+$��E��!��5���	�pK�8hݾ��$!ч�tr������z�}㶾|��T�kM�3J\���[��.U�/��#�և�Z/�KzY�t������EZ��_�ۏ�<й��Yf��/�����3�w���4�.6~X�C=��s�����8N֬�����V~z��@�!��&��⋟�1�1c�]N
��ߘ�V�$]����u1�����{�_ќ��2��wk�>�Z�BWD��wE���μ��������Ñ�� ���^����z5��5�kY�91��|8���&ӳ��k촎�#*]_�a"&!��=hYƸÞ����A�Y�n�hY��� �,�,<e����6��	��ghT��مE�k��^*au4��SΨokV�£0�Fner
�o�n�;7��2n���Y�����<lr�M}����$3��������&�G�Pg�4F3�&�:�ٜ����Ϗ5d3�:C8E�b�i������-s��_�{�x���׌"Ȥ��:rF3�|�/{��!��5-x�ds_x�I9��:5���o�$�i�Y{5?lL>��Λ�;I���+\W�#��Y���wpc�o�dv]�öx���WF���x���d���j�Z/�o:NӜ}Ɇ��0�W��[_G��[��ό���������(l�_;_�����[s�a�㧉3�K#JV����?G�_�k�W����"�n0�̑����z}�J"4�.an8`��l��d��b��G���D������.ڝۣN!������\�� L��e�p�Y�&C��.90�!\����A�$�a�y龋*C<��{��GN=[���e��Ey}���mw@K�t�!I�tC��Y"!(X�˵f��@�Ԫ�&x鸁�!->�cq6x�V��������O�뺃>!}��V�dU�7P�TT�b�D-tt!ځK,`����MTm�8��r5e�m������6r~��m
/�ag�l쮟1X�E�M�Fe�	y�L٣��V�9�Ɛ�%���B͛�ff&M�LӤa����ԥ������b�0��2On�1�Q�!�ǈ�M�DLTY[t�,��w~��H�ha�g�����bhY��w����� �N/}ꝕ��YE�!��{;h~� �h�h�g�!���E{��CA��^kk�A�����{VŤC�X��N���8I���[����W�㪼�����Y��,�{�Y����%���Ԇ�t}\��'�
���$C��_y=XZh�Y����WK<,�.��u�w|L6��sw��贙P�>���8��宬1CZ���Ә�p���G���b\��{�[����0��2��� �<�G	�����7ǈ澲*�ļxC#Z�3S=}u����m�+j�I��v��-8�̶Y�Q+j.(��7׶a���}�B{G<���
�׌~�Z�S�P�/}X�vg����}��ɎB��hz*�ߵ�E����'�KQb��O�ΥmסT0����&'͎���{k\�.\�'w�#x�\*r�C�}��z�T䴹��f�|�v4I4om�����+\ò%z�xۻ\�˴���I�;&���[W{��*��S���+��o�����芪�f[�.����qД�S��gV�ڋ\�u����
�)���N6�g�')�ը��=�t�x;ˡ�/<�!t_��;�2�9맫u��@�I31b��ޜ�g E�f���1K���D��Z7(�Ž�9C"��ׇ�T�0+�5�7���,F��k�l�Ry���Eh1"�����}�M�No��>q�$7������P����5[p��:f�9Əa���y�t��^Ϡn�v��,�Z�N���W1jRmⴒ�'T�����AT��F��uaS�f���+2n�D�!�}�x�ǰ�Ȝ`[�k�+^Zx���ҭ�*����ڏ�Z�T��|^�!���:�@.Vq��rmwJ�Ƕb��Kr0t�V��Q�w��&������o0�����Q䑧��q���;��d]-�m��z�1�s_��r�e6��S��j)�W"��"WW]*��n�kk]�ݙh.�_d���).�k���������!V�c��0�ǆ��Ϧ�T�lt���b�ğ��=)ݜ,�B����&�&ݿX���<��z�\�c�	�e������H�1/2��yE�rn$ ��M��^�W�op����,vr�$�v��}�;^֝�xW�⧽��=5��N^mc����}��Z�8���^�cl��uC���zd7��v�pf�T>��^��\��}
���y	2����9��`R8�6iÚށ�CؤH��5��;(z���8c}Zk r��]�R���yٓ�9�����Z\��/'*�b�59��#|�,0�g���͜y�|D�_k>�	�MؼQ�=��+Q��yN��u���F�H�W��|���S-���h�:��ibO�
J�@��u�gn���8����GDvF�׍W���Y!Y0T���qR{1O���=s;��wa��@�'H���^���hqt�7�:[ه�BF�T��5����)�ݢf�[��F�a�h��l�uE�;����B��{:��5Ay���2��E�e�_oK-���w	qgI�5M3�[�����D�x��fp�U�Ր�+�W��XK�������RGZ��OMZ3y!���W4����sٶ\�m����9��!�S���c*���sxZ�èW�wt=�m.���� �VJz;h��;I�1�*s�i�����B#�>����eG<��E���zNط�-�'��,x�W���>^����֞$�11'�!1�}=��y]��4+xI�����JȣK�rkA���i�2��xa�v�W=�-Ҽ��f
��a:�x��tŜ)S�l>PTֆ޵sJ}H ^r ���`�T�Vպ<:��7�ur���\���g{u�G�o���n��嬡�r�ݥ��r�F��;�Z��)r��l�#9��I�����P]I�rX9�Z۾ͥըskee��c�Z��"��%��W�"8Qxaiu��W]�c�QTl�������:��n%T-�nm�6����LP�ܹ�2]�$TAym����J�$ٽT�\j_7d	|�g58b\�!v��Y�Z䃮� Tn�,�D�Y�K��Zs ��a�-��0��:Cf���.l�b�ӕ}��>�O�h�y�R�]a���D��*�K��d�/%�T#s�ea�-��R�a��m���diA���]ݫw�Z2�� ԥg%���X̬T���-xH:�1�`a�EZ��x���R�0���Iy�V��.�(�#n�B�L�Y�I7���X���a&���i���n���R[3h*�!V����4�;���]���F��?�j
�bx6��ˌERBLy.ͩ�Q�����JƝ<��-!QF�5TFŲ�%�f�!�D����-�s*Z���u-XB2:�"���a��31��k}�w}v��,�QGY[�
.4����Pr��d�V&!Lk�Li���nc��J%�ʊ�f%]fG(����bS�%F+\q��V�ʫE-�F������1b*(�K�\�Q��*c�"ʔUE�.b�*(�Q�W
Q�DF6��*)��+�jU]STְ�ְ�i�lkDA�UQ���E��V�b�[�ueA�\�%i��K�q�5m����,U�Z[PD)��@�2�>�k��_X#��R]J�rN%Z��o���Xo��巚�M/�r�J�*#~e�a��ƅ�c����k=U�ӏ>���rטy	�{��|�2����f�k6��{��@j䥖0M�ξ�t�yKrD,�/xi,G��#��GyD�G	�M�[=�qW�<�kmV#��mv���;�:#����Oۍ ��+4i�V<]��}R�u�L3꣕X-��>�z�_mq�DQѵ$Ѿ}�}���r%cq@��+>$�;�R�:��JM��=Dc�	t�p����[X^�|=Q�ݫ�v�D�J��#�_�%�U�:���l0�l��#S�� £bVħQ������I���O�
��J���lw�Q�Pu]3���c"m��3���KV��m������)�;��ы��|m������͚�][fT5�g���5i��z�Rv��
�]{ET�u_�s�&R���R\
�Ǭ9��{Ӧ�;;����
����y�@����w�h�RٴE��y������V�)�pҍ�B��c��m=���ۖܲ���]8Z5�f�{����u��dk�~��<�g�'��$w�f_Y`�q�����:��u>��\MVdb�ݾ�p��:��X{6
�F�ܳ��M]d=ob��3SX[��
�t�e7F��|��ʖrP��Z���ݼI���6��78���p��A���1ޕ�\iu�!�C�mt@�G��;c{0�]�D[e���:{���V��^ms9���_<���s*�3�eLN�ɲ�+��ã	�w+J�o����.��I�f��K7�����5�au��
;�m`�f8�}Ts'݈�CKG�v�3)�:ڢ[W�(����V�c�ݘ�:�5�����saft��	ր��Q�<���sWi�"�w4�s7���u���'.Vt�k[�;z�mzY�z���Z�%m>���W7¸���XB�ߏ*��]h�ȘzMlj�k��B��ihȨ�i�ZS�<ޖ�Ul,�Q�BuYם�u�ik�td 7e^��+h��m`<�`��+r���X���ٝ6Y:xsfo.�L1h�l�3
:��w�u��q��4�e�?�:��Z�:����2�h1�!�v}ݤX���ԫ�Ԍ�&�;��>���R��~b�VMOu�ҫL�u�T�2*�`z��԰3iwc7���t�P�oZ��<���[��LvnX�va&-�.b�nvo��e��f��D���TZ��.��"�3�d�e̋�ޜ�ŝڀ[S~�yMc&�+w�gt����y���i����gU׹j>;�cC<���aF�X���Թ��5/ �0�:���w�U��޽Q�n�����owa�1�:t���}舖�q�G�{;2�v��1c.�l�o���E�myu�֧a]���w�W�����k��H&n+�گq��4S��M�a�wT�vt	y���p}������T�'0!Ji�!���[T���3s.:��y�z�ƭ!�Jc�<��ef��1yc��M�^�{�5uBFi��Y�1��,�������ޞ�0R'�T�Ռ*�N�v��}j:`Ip9k�-�P'Ԋ����ӽTt���B	���£
1A$��X�����$���KP	_����Ͷ��o�%��EBjr�q����7�+n����=:�쏉��;b~���� <���h�u�=��;�]�7�Tu���n�(kB�a�<�&o�Ⳙ��v�,	��m�[�J�h��J�勇Zf6w*Ы��z�rtEu9��&���|<f*��n�%���y������"yfCnR9�C^���Ձ��{M���Q�%���E�9�� �>c�a���
��b�:fw*�nn<13h��w���Z����N\�G����p;˗��w�8�|�@��<�0�# L��V���f���nWUנ��D]�>Y�WXBU����鰬�;0�;]lM��8�ᱎM�R�>�ȫ���]8��<,�=uȞ�/t	� Nq){�j���l�K׷	
�6���ٶ�~CD3�/0��Z<G����x?6���5���顥�'��m��{�i��2=a�&�xN�/Q2�Au�f��:v!P�-���Ӌ�5��0���p/��ѵQga0��������'xlw�BQ��{� G"����7������vW�z���N�3AYw��y�%���
��`�\��o�п.��ffW���k`�~a�>[^�Q�)i����X�O6%I�>ps�}#9jX�P�@�劻:E���p�劝ԫ���/-]&??7��jT��w(6�r-�f\��VZ�{n�!u�ׂT\�3��Co�>'4�+F���n��w�'�.�t�X�B���*��VYw�*�S�y����o�m�-K@��������._٫$��ꪮ����n����2����W0���J�++ld5�^�ɕ���\�9��ԑf^��4���yt������w�O�=1�*췺�����:hOn�*����k�b�3ǕB+�0��Ezr�g�I�' �Ԅ렦Dk��Ww_�zeN���_��e�cc�F9��9�W��;����6��:��_g���%0�]�3FN�
��q��'U�d#�-�zN�'e ��J�xQ��Y[Z�_aDΏ"qϱ�,�)�|/�fu���r&�p�-e҂�]���Ws��D�����Q�)JB�-%BۭDL�7�6PV��vH��}]�gt=�mX*������[�$�}��b$`�����p�}twoe���?t�+6�����[�]��V윘eI.{�^ڋF�dި�i\7Ь�2���qk�f�ս{�8�I��<�\O�,�NG1�u�sAduL�2Rr����e�����KIp��q�,Y�3����(�]�ܧq\A��q��YV֬�\,��j���9�U��I�ʏ��ˇj�2�f*�r�v"�b�rFp�h,����@��$iAy��� �#r!B�6f^]��FD$�-�är��Ŧ���@��o����G,�����q�H�+�^)x���q�l��B�e �S��/.�;����8���QuS�!������˻�L�.�!�
N�aDv.�y�aW�ݘ2���w$��%����j�r]�X��2r3xM�B;��d�B�ʒ�m*��e����)Q+	I�ZL[�.e���n�x�d�VdIBpT�%H�'q�L̫6,c����7ލ���;�5٢(�t>E1�PF�+�b\Z|�-��Uk�TS*Q��h�EjT--k�����R���@ƍ,i3*���(��Q�T�a�E�*TZ�k4h�i���*9K���s*�he��)j�m*��AU`�fb���WeU�QE�����Z%,V*���Z�f2���ՙR��cicJ�Y)���̺ц�Vbe�Tb�4]:W%im���h�.4Km.�Z�ʈ��uq1[j)]8	)]a�DB�Դ(��-/�_�X��qt�[�]�T5��6����1�wu�2%t����ì��8�
�7������te�,���|� ����m�'�n�3���M�/�q[��~��x�j���L����^�YȾ�OT�~湬Fk���7�}��󃀻�p����.'���V�]�$��>�K+Jɣ�>� S����c�se�PB�z��-t�8�޾�����0ӑev��S�=�<J��rt��^3v.^��\�B��!qhehPs;h�y󘦏VڳkfV������a��jnWS��JQ7B��aW#�I�ߓ��0��sƼ�_~Vd�T�Y�3ڶ^:�.P>���0����^��e��2��V�p:����[����Wtf���Z+7^7�L� �בyLf��nr�"�5$cdrʾ1�4w2��:	۵�ަ�tʳ�����8��^K�7�����Z��/{�jP[|��d�na�z8UfB��0�4�h�/ Ƭ�ۛsu����^��\eٖ���c9\/�T�b���/xL:{�z(������
���\�������h̓�`�����gM�@�Ax,���}�ԡޡ�	����\���ރ+�s�u�+B=���*�����䟃�2v\�`+.<�&Uωd�;%{hל�mN\�D����y�����z��'ma驜9��u����@u��pˊ��O�+�:��_M��}��༝zQT������k�������[�<��r��C�S#T�7&zT���{V$��(�Bw%�7�Έ��u���嫱�P�Z�7t���h��w�ޡ|{�Hz�Dϩ�y�F�V\��GW�G=��/+��lW���Y���>���i	ڳu`�Wk�TqM�=�W��sӓ'��Mk#V/>�K|��Q�4�����3��KE�NU����?c���}��ǜ�1^z~�|gB� ������V�:J�T�tA+c+�:i�4f51�s��z�f&+�	�a�	3�d��wM��\~c�CV7�3'\������^�[���
���*X���me��b�*��睝�9�Fqy.��R��<��.������ԭ湯ԯ���=*K�q%n�®N���=<
kM��C�T������`�l?nPk*Bocv:k\��So�I��� �y���HmҬ�Nk�mP��0^=�B99����y�b�S������is��D+pSo*�𜳄�R&Cz��&��F�6us�A�o �Ws��|w:ò'�h����԰��~&T�s=�h�
[�Q�C��,�\��Lz�_	}�]�|.��G��z�fhyo6��b�"����}���a���l�ME��7ww�0���N�d���S�h�o� /���{�P�����p^�Ͱ��$'.��v[�S����վ�W���a6'����Y�)�^�����q�v6�Nd�������(�V���սqe�܀�<����|+.�YZ�����S4�m��\k��ѓ]��ͫ�ջO3D�릠��B�oӮ����d���kg#^��ǡ��*%;���Y��j��F�T##3�"v�޻�.;;8����^.�%��+��R��Ż[��7n^M�L�.`����<]8vs�Ǎ1�#p��F��u<b��0����3�e��W��a�j�s�J4�q��cѷ�0��[�X��_;�Po�=����6�p�Jw�뷶mԪ����švwB5��H�wz�[�}�p��\�7���|b�"P�Ob��f�Λ�{m_Y*��GN�)�� U{?j�k}WVw�N�5�
�Y±����̬G�	�uB�;�酄fn�Z{N��k����&ɫz1�Ŭm���s2=�J�mԮO;�#k�U��ۜ�ě�*jr�Z�׫p8U ]nS�Q͘�c���i��rMs�Re���k���{I#�^Qʴ�*I^���E@�cJ��=u�:���;|�i>�*������9[�E����<�����eWJI�b��Ϯ�L�hת�_���:�+�����=;t��|���7h�:�K�(�RC�7�m�w��s�Ѓ�{��n��&jt�f���I�;ތ�AGG�׺��f� �fŝ�(<�F]c�*ϵt$v�۽�9���������k+�+�]��]�o� [Cءr�z��TFW�"}�˱������`B9(nE�5C�ޒ4����]h�|��}qiƎ���~{Y� ,��xm�2#zv�dI3�՛e�6v�p{W
Y�hG@Kfo�nQ등M<�J;P0�9s��WT]1�3Og3��ǕP���b1z����0�fg�y�^-y���]M�<������{����\nW�����Y2�ޢd��~��&g ^(�*@L�'&���r�ݒ����Ϧ�8�A�V=����l+�#ouk��\���]�<bʡ���x�n��+|�9�f��'{����en[X����g5�'�<��뇘��B���uܗ�.�������>;��9��krT쒚ݱ��q�j3[E.6�.nI��_ϳ=�z֕�_Cu;N4�����X��>"=s�sDʶ�r�]B�H7Q��Eu�Xr�������/�[��X�F���Q���P˒�S9��x�u�&�����<�؜�b�d��IО�{}�`��:�C���c����pϳ��K���_2PݧZ�P�}ۙ �ΙB����3� ��{�h��\�+�v!t�&	��$i�*��s�;�P��P��}̻�r���uݒ`�	��ZFe�)]���dŊ)\h�����ٳ�ҲzhiA��o-�ѳ)�~�9�(�5ݣ6W<�F��:�1�d)�4Љ�bb}ʒyfF�;��y���;k�0�$X:�|8e���P�R�-�G7 �ń~���ܣ���<U���iynI�+Z�-k���Y��.�����F�	_e�@���r�Lp�3.��)��(��W)X��c���d�2/Wr�;��駄�S����w�R_s��iU���N]'���԰%Wa�Y o�/w[�eXT��Ɯ��)%������V�I�6�!�r��JX�f"򍺼�u#�l���D��#!�JÁ�R�}�����UܦP4��	����l�rf�5p[���Y$TTD��&����D
�,YtX�`�a5�����P��"cˢ�Uy�K
xc5Fф�4sX�n��g�i�yb��8�j���F'��Y�%S$�(�T��yt.fe�;��k%`ΖB$A(�E��[t⨶�E��h�k��Qb(i�Q][�%�f�+JV��1bL�Uq�b�,e�U�k4�VasW-+er�`�*6Պ1�ƈ�j���b��c.��+0h�-��,Pt�P�(�Daur
2*�r�L���V���Ӛ��1DDj]WT�E(�Ī*[,r���,���Z
f�r�U��sN��h��K���j�(���Jՙjܤ�DV*�̪1K�%�H�����ݞ���z�+�������n�/���Y�㇙<�n]��8�����3�R#��tk���@��z�9�\u�\��ccg��Z�a������e7Nl��ik���=��)�Z��nw\>��N��.,�[���w�/���M���Q���[Qp����j(嬍볚��ZCm��ߑ�C������ī�5�vno�g7���OGr�M���Y�3Iz���Wwx䬲Ƃ��x��v���d1ntoX��
�qCi9����qQ��qY������(���j��]���ƛ�n������0���utw����t�J�L���/is�JNYc�ɝ��B˳ �@SX��n|���+�i]y��*d�{���}���f�i�+456�=GK���}z�N���1i���h�j��tsU���ާ �q�J�}�<�rڪv��P�摘Ky���f$P����Ӣx��qپ�:Ҕ��6�sW���c��a12@x$7�����=;Ι����<����r��0�֙�d�vy�Io�+�;���ӄ��RR���T'2�:Q���^9����U��D=t���jC���)U��j�όUއ��h�XNN������n�Yf�Б*�YョG4��}�b��ܠr�jc�'�J�ړ'2�*	�� !���j:���gN]��"cG[�&�����k���_U[�vg;Q|�j�(-��R�m�=� #g�eA�[�b����U��9l���w|*+���E�/�n� +�1X��'�&�)xT�V��z�Wc/,S7�]Ξ֏A��qDvqd\[ˇ�H�=Zu�����}�ע#�V%�c��sg�&[Z\7;��-;J���m+���U�xM�ʧ�uC��-�3є�Ļ��h�0���228��sW2lj��mA;:q&pĭ�;!\v�$��\lM��|Oc{�_B�>\-��%�׆,��!-��~b���Ns�*�۸�Ϲ�Hj_�;zG.�ZƬ��QQ/l��лi���n�������~�	�G{��Q������A�2�����6�@�2��X�ݎ+���&Ҽ����X�l�d(^�@�VM�Gg���iޛ���q���`��RMV.6�v����x�X���F�&N�WX �T���f�$�p�]#���Ho�k�^�ǵ@�RyL�=ai�zE�l�٧C[ڥj���&���O���	����]n��T���zD�jFO^��/�:�m�-��P�>��զ�-��ڭ�]ϮE�̆��.P�p�O��[�1��l���[wO��L��3&�S��my����
��UY��NC�ܒhz3t+pq���~g4Ku��;�z��nu�3��nĭ�O~/���p�]��{6Z3��L�*]G\I��E�\��i�9�]��{Zŉ���խwoHf�Uٯ+��R���6�{�� �����3��L���_#s�~����^� �EZ-�����-O�]S��z��=b�V�b��38�ey�k�k��|��؞���WV0SQ�O}�0����5�P�����ˑ��j�gB�w0ao��2��g2;�!�T�r���{'����t膝:�_H]�j�ɥvPo������k����i�>ZtR�l~��� Ax"���cf2
\h�Q���,��T�t���h���p��0fi��ҟ�\'������W��a����=��2�2!A̡�^��9Z �B4�������*�D�|y��7��=^NB��?�c^%kս�2�]��]�	�"��^�ٚr/07�w����Η��6�|k��nsNE���7�2���2"\�Mm-��c��ebRz҄��Ba8̐q�6�Ylzcx��#qV�z9άW�i�#���[n!�kdJ ���^X�*goq�ؘgݍw����)�w�Tǲ�q��]�+��F�k�j�� ��rY�#9�2�A�w�Vʚ�rXt%�d��u��;GG�B੻��ъ)�zֽ�z2�a�Ò3svz�_r�?Jc�~{��llygo�b�QM��(���Dj�4L#�0��q��޸5�5t7�=���aȪv�_N�5u�Q��;՞� �!�ǧ�U�x׵���S�u��i0���Zk���C)Z�,�ݲv<��Ɣl,k1¹LԹu�6�a����Yx��)z;{y=�µ�����̶&��2����S��N:����Z�>^�u�&iW^�f��,>�vD2vΓV��gr��tZr�f,'f}B�R����ռm=��8Vb���"�6�%������g��	��Z�E�E,+��LPƅ�V�鬩�m+����+��7o���Y���TUݑ�c���k�h$�x&6��^���!݌�Ls��A��fO-���v�{�P��#�kE�K�WiZ� ѝu��x��uJ��u�J����(��\�97��Ҝ~lN���J����NE��-�Mwc�OvF���@_qv�K�t�F`�dtLHo#"1�T����-�#�Cۜ,]k�b�)6��{����|���4T18����ZˎX�� ����gm��R�H������{]R,p��<�C����c��*�\��5��i�㹯T�2�����,[�y�A��4���wf⧫J���S��C��Y��`����x_�%�M����st�<Ҟr�52�@⣘�F (	t�k�%�1��/95�'gK�g��&T�w'��,oTDQ�~}N�q�G2!R��0Ψ7i
��}eA&������K�7��ƌ�-*LE�����D7ӆ�z˾��ټT#oC��3UdB=��K�}}�;8>�a�4s��t���H�m;���X1�޽�$�I���N�^tf�7�u��e����㵥�X�Z\��$��:�&M�mѥO���V_$w.^��&�zڦ#�I���j�hFn�ᝮP*�Y�2�Ȱ�$ ��V�ҝB+J�G�ڳ�V����o.hw*��ƴ�@�ᛍ|��ՕYհ��@��O���h�AZh�b�e�xp�����6ʖ����wP;0b��cO_|�;�m�@�������ܶ��ˊ�IR��G!��傳���u��⾃�\��	Z���Su��e,�-�Pn[���{�	����`���:�f�_[����b�7wՁB�٘ݛ
�S��ee�ӌhC��Z&(�m������r�{�2�5��k��r�^Ⲅ�ܕ6��6���i�Gi�˭V/��`��"�NFf9�%�մWWX�����xm@�����iIr�Ӥv�.��wٛ��/{���?I��$b��鬭��\j��撨��բ���Tm����J��90cV��t�VV�t%$�����T�c42�ʨ�q�KT�%T�ԳIZ�JEr��T�,Ӗ��b��5s��Q-�U\�\պ��XVi*�P,Tr�AR��,F��,��VTMĮ\��0V!EEejbX�PS�+G�I�$tf����]Ů�54�,-���[E��SY�5���ՙh[�AV
�GI.69f���띾:��A����q��n��d+��L��:��$�:�mO�4��vFtm���Y��&�*z����u���·9��U�讶k�!R���8��r y��:��}v.>T�n{���ڋLC1������*1�fć^x��м��F��0���]1�=��^M<`M��z�����}�"9앦�6s���8�u���g�Tj�ON��B���g�+!��D�֙7�/���bL�HuW4Yg�7�MX�n2k������\2�4��.Y�:Y!�ە��Ҕ�n�r邷y]YH�4M>�����Q{�2�#���$l����զ��0/ѝȖv�u?{������8Hos�hϬ�������&�4�*Ѽ����k��t�o+��Vv(�	�ݩ��S�\�b���uyƊԮ�[�����8�kֈ��>��Jyk�����r��x{ڪv�r3�Hhl����'r)��2(�?n�(=�y����G��o�)v�øKU�Of��W;"q��t�̺�8Ľ��T��A^�����6J)��J����fa{N�J��(u�����v���Pz�3-��ĿFwwf�I�F�b	ޔx��gpu}Y�峇����\.^w�鳜]F�	��g��=8��e+�N`�s�͕�Lunv�sL[Ӕ��
��#.�$�ЊH�ٞ��aK�t��U����;���f����y
p+�G^kV��)�X}��;}����[]I�������Z���\�s����Z$R�J�8k��C�c+ҝ��N�����-
����}*�n�U���}:Y����s�Ҋ~�+i�V���������7n�������D�t|��WyWGE�*���6��$j����%��.��K"J*�ùXK8u#D6e�d=�����wv�RWs]w9���u�>���Az�W-�OJ�{:m����|�{W�LL[s�4�ⶼ�3Y���q<f�X��Kj�<��.��Ց=+�-;fxC���{ �@�%EP�:��(g��hu�uo��e�;��ҹ�t�+J΍��r͸I
�'2���d��'�{�uX���M��=x|�z�i=$p�C�z�v�Omf׎T:����#�����R�"�>A=�Eߤ���.jg��ЅT"{�f�^T��X���̮�U���t�
���,㩝�>�X�z#0G�k��@�*����޴*�"H����t��/���$U<�m�����������v
��[j��أH�s�uѩ\#�q�_�Ć���5��U4~�m�|���O�iu�MJs�:&�Լ�����
ZL�7]"��N.�@����z�A��=�:�91�yai��B�3O�s�����X<�O'���I1Ny���x����u\2�lY�q�,��� ��%�󾁖2&4�k�p�ĺ�6wv�ټ�-[tG���R��?(�Ff��u�=��'[�v�X�Q{�����Hor�
	�@�1ޤso���x���*9�ibԧ��A"����b+;'[��~��v�;~؂�3����0�/p�Z�V�qb-��y4<�}���5�qt�,v��t֧�ށ7���k�$޵]O��\iԭR�*E������!f�F��e�,���8;��h�܋�|��eC:��xv$$�o:�5��뷺�����o��.ǏNv5��_tiL�NX[K�[��Z�z_�_��w�sJH���Ǟ��5��V=]�Խy���.��UCɬ��P��q:���<�օ]uc��VS���0�Ѿ�7���lg8�F��O (V��uڈ�'-vuL.>�f,g=��X����v4.�	�EU������G�U2���_"�s�5������q�n{x�ҳ�h����B}v7˭M�F1B�o,o���P�qu�ͨC1Wf۶m�(\x$ƽǱj��'�1��mjȽ%�1A���x\�Ļ0ν�2���T����Kr�~�&�SE��o)6��۱*o;���U��g�h�a��~��r]u�+ z��:�Ʌ�/�vo'A��0=��{|������=6�)[g���3֤�]�-:��[��L�<M��f���:i�)��Cy�Ss��d�Y�k���e|1'ҏ+]���j�__,C`Y�+]�$��A]�v䙸w;��r6���5���̤�f�Zۗ���Nyu�������7��nz��/Hߟ�r����=���+�[[<����}��R'�ӣᴁ�	�z�Q�b�:��_&9����f���b���Onl�Lk=qF[�����H���t3զ������C=����v�cߋa�ƭ��ڙ޲�+����1W���waqj5n�l�1hްF�K�B��ϲ�م36�in=8��o��+�����[뮧�}䞵���2eB��չݘ}Y]�\8=�Ϋ�׵�nַ݁�{@r�i�zs�c7ji1�#�^�RW��B����3x#��K���e����Wd&l���P��8�k�{�����;�A�����FZ<�U�q�x��r���W��X���X2n�Z=��,˒������d�?n#�2"�LLDDDDG�L���$��AD�x$� ���O(".��,3Re��<)���������z����������d'�na��֣�A)�`j��B��uC[k�72����v�PQ}F�#(����_e��&����>SNî�&��#3Vy�o�;���y0�/���+(fY��5�$@_�3��2�^�L}�!T@_�@�@P��$��O��$8�_�p{��ğT���q�K<u�"N^(���@�7l1:Xi�1[�B�6K�� 6�Y#$��j@��֡3�K���:�xu�F1��(�����D@X�ќr����"�""<�TFϦ*Ɋ�D)��Jms�,Ҟ+�ɯ@�T��AD�����Ssm��I��!��.)P��@h%r5�W�fW��}�'���H����&�!��۹�9b��=�������ϭ�����9��. �{g�����""ɹl���1N�jC�_o��p6�Qv<Hc��=F�&8�q�}�&wN�2:�El�h(����b��NrLJ��3�x��	а�˟� En6R" ��4hF�����P[60 ]� �Xk�Ȧy�^����B�iD/y;�BL�X�\h�U@\�w�ߐ�ӂ
 ,W��������G���������@N���Ue����r^�;^zD'�=B�jS�Q�W��IAD�]��n��1	2J�=��#΂�+�`�s�?�$�2ݡ��=y��������f��`Cqh�z�ԠAE�r���m�=;��-~�dC����z�>�9f�k�u�����e�p��Msʥ��H6d��o��:�Í�~%���z���h`HD�X�`ڃ�<_?��Çb���Gy�6�º���7mf.��Bh��,]5�D�|	����s��EܑN$%)�o@