BZh91AY&SYP)����߀`qc���f� ����b� ꂒ���                                      � �}2��}�   �    @     �      J  
            � �7����
�))DT���J�	U%)����*���EU*""E%
��U%R*(��

�H	��Pn���I �J����!���H#�(��X�P�n�@S�����
0-�Pv��;���� 
 ��mh�}.;�n΀}[�B�^��H���� A�6�m WGy� v䀛�B�lx�B������ �  ה� (��Է`*�P�B�*�T�T����(��� ���
���h� tN�Ԫ��@zn�^�{��p����`�7�$Δ)�z� 8( @��J����{�I�.� S��� ��{��` `�f� �T)� �� ;�!N@�=� �  (P��  >�*
R�BP�"*	S��A�0݀7�f��@ wxyH^ �ʞ���< ��rt ��!J<���`4�`9@  o�)  p@|���@	o{%I.@}�㗠��r ݀�� w$8 -� � �`��@   ��� | R��T�D�T ��@� @C� c�I�(�<� �`x��z�T��q��q�J� =1] n�C   (:�=( �����&ℋ�c���]� $ q�G $r� �� � wϒ� RB��D���� �w�qAn�: w)
� ��v"���݀]�H����l  
�_T ���2>� J ��@�r@22 a�� D��2@22 �� 
QQ  � ��h)T��@     �#)IU@��   ��T��*(      6J��T�      ��(�JT�P22h�	��� "D��JJ~�lM)��2&	�C�h��F�>�w�������k���|���v�f�s�0��T�}q���
*����(���
����
�W�������@��v~�?���ˊ������*�I'�TW�*DTz�����%0_���
b�%0`4�)�S�)LR��1Je0H�)���#LF�L�1�L�LF��1`��i�1H�i���L�-0Zb��0�1`��)�S�)LH�)�S�)L��1J`4�
c�1Zb��i���#L���#�+L�-0ZeWe]��mvkvV�ٵ�0i��0b��)����ٵ�k��n�ݛ]��6)�S�L��1�,`4�)�S�L�%1J`4��`4�i�S�LV��1�0Z`4�i���)L�21Jb��)�S�)L,˲۲�e2�ͮ�n�n�i���#LR�F#L��1Zb��i����LF�ٶ�vZ�5�Uٵ٫��ʻ6�5�+vV�5�k�B��1Jb��i���)L7e3k��e��]��-vV�����ٮ�2�e��]��5vZ���٫�WgeL�LB��0`��1i�0#F����� -1 
b"�Q� LZb�F 4� )��LAZ`��� 0
`���P�-1i�LU` �@)��LPZ`�ԄUi�`��V����
-+V�Mj��U]���թ� S  ��%0
`��E� �1#F�*4�Q� �0i��Ri�#LZ`b�S � LQ�"0
` ���*�-U]�\J���m�-Uq+Z�-�]�ծͪ�U��i��SV�����!L� 4�1
`"�U� �LEB���H@U�(F !L
b��i�� )�0�-1Zb��i�����+L�(Si��3k��f��]��6�-vZ�١.�]��5vZ��٫���]��5vU�We3]�vj쫲��]��6�5vU�k�Wf�-v[v[vV���J�]w�S@�z�Q6r���~��#���`��ӎ�B�8{�g�T�:������~�ۗ��pc'.�A�_m�w
qW��Y�.r�ۧ���;��|�1&����Ku�n�خ:� ��!Ğ��n>Fh���uѺql�Y�n⣰�ܴqsO��.W-x&�0wV��ڻS��X��۹{���f�E�]�@�)qRp}��g��Xq����h�tI1�1ݳ��n]3�QN�z�_�@�v��&�,X�;؛�d(�x�Z;^��H��)ڱ�x�Ze\�7[4�ʹb���;2S%�.���8')��ⷲ�Ekz�"\��r�:M�N+H�����Û�>���9I;��n�z��_h\�6��z� �]W �"��dZ7�+'9,�V���W0B7~ݥ)��9����4v�LvU���ܬ{�X�U>��G8xn�<��6�x\��9�x��vLX�cqռ�u�,�L\{{�̝��{&I¾��n�y�/5�J�n�t�&3��(NƆ�9� ՝[��nlz±��������_h�8�Oz�5j��,M�Ld]�� 9�q�9dǜ�͹8�;L��p>d7�6��	!V�iBy�wR.p��L�l�.
g�v�)#9
�:��y駶n�jO[ ��N�����VI�B�ǩS������I���k��ŢC-�)�θ��ؕ�e<,)\�uPV�ے��';H���6
���ץ!��`��a	��w+���nn�EǷ?,~�z�{�c�V!̸�V0��t��	>~-��H//9��S�e�C����\`�i��E��:��t����w����ǵ ΔVr,����;,S_p���@�̬���P�Pt�ۺ\�K���w�n�д����_ӊ�{E�=����\�d=>�|U�v�g�l���	X��� .J����J��5C�����P�p�f��gvQܺ`)A+�g%+�N�ksrj�qu����h|�'l�h��r=L��y>���G�sU�{�����Zq#rܯt��dC=5���#�C��-��!�u�d��g)ɻz�͠+z�l�QP,(��t���..KV��򏩯�z=Z��'�S�ͣK�D � �ݵ(4`��Ќ������o�Q�Z�՝�K��օ}Twa�^z8^���v��X�1rQhb�ѽe�]�s��_'ٲ��;#Z����Jٰ�����\sm�hc_g1�ϯ;E�2�.nj��Q0*�X�k�NoFMѱ�v�沱!���ϧ���BÈv���[P5m|���}B�q0��
���(T�D$���֝�ROHx2az[�c��y�YÄ���(�#���
ݲҭ�jT�viK U�-�2v�x�����p�Gq7���ۅ�1�[ןbS��H��w.�Ζ��k��ÂI�3c/����r[�-wq�pX��p�j׵h�,X�}�Ģ.��s�{���M�ay�,;4=@��*��l[Vp�r���������F��Е7on�5/��a�P���F^�-�AfaE�B�)��s��6���$L�gmܫr����L f�skʹ>�ۇ{v�pb�kk�$){�%Ǉ�L`�r�ZzQ��q&l�s���J�tj������[��5��v���E;rI�%�k�B�ӯ�3+Z>��s촋��Qc�;Ԏ�@#�k������eɋ��q�OA�MvM���Vܛ�0Td��i��޺ma�D��$�)�X�{MWV�m�<2�dsz��呩�>%���{����$���w{�%q
`*�������Dhl׫9��$��gg=w5ٝ)��:��ꋗ7�{��nܸ��@ F���f��f��[5^�8F*˔�#$�6�k�aJ��l�lKv��7����r�p�w/i��S�I�f�5M ��;M��N]���ǩYrd��"��un˼:[�6'ٽ���C7)�vh����$^
3NK�a��1<tT�ɉ�{L=����N���e���sА����]�ށ���n�t�t��{9L���e ����Y�^���8]���.�l�l8�;uO��"�:F�1��3L�Y�W�����������9���y���d������r�Q�וev4�]Њ������M7&���HRZv�3U�s{�RGlp�g,M�7��L��# B�����Wݳ��hH�!D"J�wF�̺r���	qǀ���j)��
9�8�ͭ����n�4�b�C:���)��U�=�Ȏ�0�qN�<�K�p!Tp�A��T�����X��s�Z�.i7�o'3r��Z�#�uF�{�%���eYfl|'6Q��<�j��Av��ٮM�\zgXr�9oAuŽ^��L��Vnnu�pgkۜ�v�����cr�뺀�tN��+�t���X��)�b	��@򡧹;"���zP�ۜb|Wr�f�΅��6���W�X�vJ�S{��(��b`2e,�
���9�8@[��U<�?��I}��W�{sp���'�i�A7�y�-�i a��8*˺v9��5�{mSD�HL�����-܊��aӭf�6F�CD.���C���|�|�=� ���B��'6�o��"�@г���4ko5��c�u�yv��s��z�Y�/wn���]`I��:Z2m4ˡYVj�Of�J��&w��uyF�+]/�zP�Gw�PHNA��!�V�"���̗5�>�=Ǝ�W���Gc3(YHs�v��b��Aݕ��]�(�v>ߧl�?	Q�y��gDѷg.�e	Ӽ��:�%z0���Msה�n����#z���X؉����m87'cw��:t撷 y0��7&���O���ĵ��0W�ɡ�P��ߩ�+z
��drNÎG-pd#�8�^�u՘�=�9�Z�c�.O�԰2[�k٬�R��1�3_M��5��߬��pk���A�6��x9��w/p�{�Y��f�26w�����83��/Y�T���;`;�qm|]ۀɚi��r,t�S�tnS��n�������ГT�%$��,M�-�c�)۫n�n!i��hv#�+kt�jh�رf���-+x�=9��c+��ݝܘ�;�or���#����i L�}s�p��G��<R=/"�a�Qܘ�c=�`�g,\ I�$9���jni�\2n5�+֜Bv�V���a�3G][|��������8g-�n�� ��w#�B�5����C�j^��.ݎ�;R�qh�{��I�Q��$�ڇ3���Ӗ�e�7q�FM����ŧ��q����7{7p�ʰ��x]��Mn��j7�hG{�ܺ�^��跸c=\1���N����� v��È���z��<X�o�h���o�u$г�\�8[O*`�qp�5 �nveH��c���׹Z4>aDq�nR���Zpw}�,uQމq�c��n�D�s�����Ӽu��wC��)�<d�r��a1�כ�r��9j�=�]D��sYn��[Od*dk�����o�k�w'qٽ�C
ٳ*����=y�p��bS9ټP۲���n�ɨ�0�Kw_\#jz=���Is��!�@�ם�mx��2�v����(�c�#�D�T勧9��x���1��m����/76�1�a�^���]�C�wd���_K������95;{d�|WL�E8��P.Lژ��Y��&�@r�g���Y�]z�qd, ^m����m�s��7�G�qɈ�%jwq����B�VB��ů�o;z+�:��v�\]ۋ.���NE�F^�!��R�8��٫5>��R�j�a���;�2���![-B㳙sV���ݓ^n�Ye�Ǻ&���W;���s�g7�c���y,�K�{t\�y��+sj��:[3l<5=����N޳!���/R�C^�~U�1�soZ���۪�6��s�w�0�l��s��6���,���6`�.ï`PfX�(J�N�u];>�'���d�(�F����f��±�zY�L���N�8{rpiz���^j�W&��{i���(�H����w8Lv��HL+�D7{y�M�B�\�,��e����<�8y�@ٽ��\f4����0D\FL��"j�Z�H�Ѱv�o���ga��^�s�Q^e�V�{�`�g.U�@���kc:භ�3W-��+rf¬yt�˺8���!�s&5�O^��h�k sx`�ջ����<����S>ˁn�Uk)eG�\�	��W�����
WY�t�ّ��Ǳ�O	�pKriz㛈��h1�9���qr�qK�#�>;��#ŦrV!J���r��;Q<�d;>7KgF�Ep�u��xw�:�^5����W���A�"�!��6t�Iee�EP�q�<!��f�7�Bx�zӓ7��"=�p��=��qd[`+UmaҧS����؋װ-ĵ�>�B#�"
�P�L���z��죃L�1��}�#��ٽmVk��--W��yQ�"J`;����W�N��v�7�"���q�`@o.��R��ws���`�;��%�׺��u^ov�j=����5VLٽ9-��ǻr'�}�V%��zv��[���c�z	3�H�7�#��Dr����d��#�ټ��8�z�X�{y����n^��b�to1�����=���cX��̪)���Hy���YqWe���wmd���ڮ�b�E�b<ɹ]�Q1I�ii�p��7aA$X��)�zCǿ#�m�wl�ґa�n�8�����a�D���;����e�QX2>P��;���}�I�r�� #�z�.[�פ�� -��h��HbQe�T�kzȏ�쇎�V0��.�p؀;�_��G`;�4ph��=�t��%4������U���;���`�=�p�8]x�]'�#�T�v�;�^��њ��p���"t�B�bx�yW��$H��*�Ӵm�(�>����twY���8݂-�sֻ&����AP϶q���5���x�3���gmvO�8���]͵����[nɴ��G��wZ�������b����p��!�fkz	�-Y�xk�YnTB�Q�y��vܝ���j�l��s�=�jZX΋s^�{�w���[&1�鋆�Ɉ>�e����_�&e�M�N<���ۍ����e�����ݖ�Vvm�q��[Z{&+�{8!��b�g^�CᐖCv��痛�g<�N�V'i�,�v�ݜ�����:��vf�Jݬ��D�1�^��3�Mi��gFSލE�@�Va(��\:6wLb�۝{�{v���7z	Gșu��%�*��cl��+mw�ӤKct���^O;'�]X Gsb{��+wXs7#@UZ��H\�C�Ov�xa�_k�,�5=Aח���r�N�*�Y�K�=������>k���K�����n^|�:�xuU����npz�Zy`(b�\Ah��!�z�-ǹ�Q>�	k�j�P����Ƈ��`rx�j�8Pu���n���6.h�I2����h!����r�*�x�e'�{ۏ�]��n�ѯ�P�h�`@�Lׇ G0+�ebbb��9qz;ta�w^����ڷ��/�������nz��¼Wmҹeu	Ȩս���~�-���){�n��=
�Y	j7�Fp�qś!2�"(w�sC�Z��{b�{�q���N���w�I��=�E�;�Z����4wF:��1\BD�L�Z��9$}�:h�tk�d������"�g���4��dM.�n�����e�i^�|g��g]�t�ұ�[D����d�K��d�v;��,:��3s�9б�:�S�Ǧr��5N���QZ���֩���V��ݺ�1�LK�C�����H�ed+�`��Y���c���3C�`����|�U�cD�4W��o�T�3��,Rȹ�43�[��C��f�㝃��
��oj��#�6�&^���plq�[����@[�3q��ys��{�\��G�"K�G�nw+���B�mƺq7��ln���T�,��x�z���F3���zt30���G2o� z&rT
��;H�,�ou�p�h��v�t�V�6~�yM�S�m��9���%A�f·��.o�װ���@}:7SO�l�E���)�m��O�����������Y%�!���Q��Y����ͥH��5���[�ڋ����v�Gn��;sCR��^��n��u��!ta��CY�p�-�r�%�cL蔐)�k�ZA#j���o:�uA�iy�����C�L��۸�\��v��Oe�	���X�� _��ُ�O��T/��Wo`[_���݄µ
u�݌�|��Q>=�M�t�2{ d���S$n���.�`W���-Vr	T����:�{���8�ۚ����4-�)Yd������-'|ۭ������һ�H�����;:[^�����3B������Ͻ���q�)<2/M��ݜue�t��F������ٕ��P��g ؑ�>�����+ۼ2���ϲu�	�yg�ރӂ��n�B:S�@zg"a�������؇w��w��'T�"�x�Ry����8�&�*��k�����"a2N���xi����W�d��"Sƕ��o���.:oy������-b�#�=����n�ע�;aw٦�}�o赟��~�.��g� ��c�n��.\Я&}U��a���0�u�N�u���&ۺ�'xq<�h���&�|1���d��\���vf�\}I�8;}6L��ې�d�'�|�����*J�G��<x���k���e;�xŧ'�Q��f:^A���VIK5��51��j���Q[������������: �d�Q	 EP�Udŭ���V-���+V��j�֣j�mcmV���V-��j���ƶ�kk[�lm�j�j�+k�lV�ն���[�Ej�ڵ�6����k�h�Z*�Z��ѵ�+Z5cm��X�b��-��[��m�5Tj�F�Q��kcm����kETZ�E�m��U�U��kkb�ŴV��Ucm�m����j�%�clm[Qm�V�֪���j���F���mj��mj��E����j�m��ժ6-jŵ�Z�5cZ�t�$	:v���3�O.����?������6�|ч�<�i����XL�Ƞ1 1ce��^$����<||�_ �S'����z��,��-?pd�̜�=�[�s5��<�K�5 G���g�з�-��qg����E��uĥ�&_*/�P�|�4���6x  =�1r��) @Ky���x�J$s��	�ճ՞��n���x3Q�8~� o�؝׈�}����>�r�hzlRK�o�)w6��tġ���(��|G��Z�I�wo�HO<Pћ�(�_DF�y �x*U�����˾��Y� Q_��W۠AT@���>�g��_�_�| DA�'��/��ߋ�g���Q������y
�񙱗�#=��t$v�UEy.�E����y��
��t�4�`�3}�5���>��^p�v,|��J�������nn�i�ڷ=s��ta@�P��v�H�f��c�5cҩ��d<}�ҽ�J(s*�F� ���s ^�un=y��Ca{!��^��~̤Sh�,�����0��t}�wn�o�����3C��L�=�ֻw�8�{7�#��ᐼ� �{x�}���޷�_�փ(�(�/p2��@�X���4�Z� Z��Z����y��/F��(~m����e���S�y��ny�93O�h�п/w�ɧz�g�/%n�O�<<��oi2�n�@gD�P��V���ti�����.M�}��|ǽ�|o��J��j� N`�/�{ޣG�"|L[���f���T3�ޓ'0��^3�c: �7%e>���ͨ<�S�h������7�1���s8���w�c��h���mŵ�X�C�LKxF�o����f���j2�ū�K��ۀ�x���sYٚ;'r>���իӻ/b�<�4������ ��%O5{�&��B��4�׊�b�ཞ룴l��2��xi>`�u�g���{��������n"4p=���]��Q|0[�פ����Ր/���޹L��o;x^�Ǟ��7&��.i�b���8�{N,�1�ݐ'2ߎ���$c ����{��/Gzd+�ߧ����~�ǎ8��8��i�q�v��8�=�㍸�8��qǧq��q�q���8�8�q�q��qӎ8�n8�8��8ێ8��������8��q�q�{pq�q�q�q�zq�t�4�8�xӎ8�8�c�8�;{�z�y�w&N�Sc�p��[}C�_m��/z�֬�!�X���룎+�f͏��&ʽ�M&�aÈ��ə��7;�8��×~ћwc����5����w����^+�i_)H�ĝ��cV����'�4w,�����M(�S+�w��W�3�a]�^�Ft�6{���;�s}�9����5������Bվ��{ob3��;L�@���5�:����z�_�<�O^�,�K����.ڝ��\ǜ)Ze�F9/7�ޖ���e�C��\�Y�2�Cd��:�{��:;WuG{��b�H׸��4{ӣ`�	pc���Ä�큸o�O�K�f��]���I��5�3i�t"�{�ٸl˽�q�,��/z22���o=�	��<�ɯ圖��G�	�{ZvH���9j=��L�㛣O�g���������v3��>6���+1Ȼ�^ixo�������z;9�O|����1vу�yo�Y�:��nl#f��s�q8No�ӵ9�6g��]޻���3n���j(��uGG���rǛ�N���y{z��;w.�����8U �Z��$�r�_7�o���߷λ��gx�É\������w0��gz{�f�4yr>��4�d� �2���x��̓���\z�
�3�O|Vj �>ɾө仼��1[�DO+�n��>��P����+�aὧ�)��N���09�m�=�q�8�8�1�q�{q�q�m�q��q�q�x�q�q���N8�8��8��i�q�v��8�8���8�=�ooooon8�8�8��q�q�zq�t�4�8�8�8�8��8��i�q�v�8ێ5�f�|�p�}���&2wp�~��C1��f�P	�s¹u>&��\��������JW"/��;�v�v{�kd~�7��x�P��WX3n{��|�.�v �;��t��]~Ǆ�{۰�o\�WZ���_��_���T��;p{�ke�Խ�o{n��-�c�<�a�2�2��h<~9�����o{@A���5a
P�v��=�����|�R���k�],�_�D��:s���JzgL���ڻ�f��:�*)&��G���2���x?8a*M��^On�`���6]x<�+����?N���po��ϝ���G�=c����n�o��j�yɛ|�����iF���۹�w����&E;C^N��[I�u����˖��u7nt����e���UU�p�*�'^�^��*�S�t�_L�����ۯ���>�-���� �޸��y5�D�w]��=m�r%�U����R�o]�}=����/�r�f,�v�E���,wԿ�W���z���0,������K�N��>��}�a�fL��󧒔���/V�2vvO�zc����|I�ǏaإGa^�׍��*��t�����znaK;9<ޞ{�`�����HL�sȽ��^��ؽM�����}:����a�6�A����#�����Wؔ���������|�7z��x|���f�֢8N���{.���䂗�{�i��{���!�1����U�E�&d9�O���~׋���糑~w�q�y�n;a7�Ti���^����� =g=�u1H�;�sѠ2{�E�o6��3R��
�r��ݠ�Z�
��,᝝�|�]�0O_I���صr�yA�w)C=H�{�8�����~ʒ>	�\�>m�M��i5��H>��o?xO����X�{ϼ(G��}�����O.���sĳ$˽��	Z��&�2��P�g����f��w�.�+B���x�!�^B�3}��1^xi}؄����'F��0��s�)�ϝ��F�n��pݱ��)>Θ�2�Đ�PP����{r?���x�#K�~Azu&5���G%=��9꽞;��ެ��n�L6�K܇�E��qL�Ja�(c~q�������q���y�T�컻���7�/_Y �-��*���t�݄��R��'r�w/N]��z�|A���2��В���qݡ��Ĝ3
ͻ�l� �r��NW���۳;�f�g,S�}�z���u;}W�o�nP����֏��W�����(]���⸭�Td.���B_��b��W�w�sw����!Hw��<�����u�!��m�<�>��o�K�\���΃{�c����$#q��|�	)��{ܞ�^O.2��4?v�5#�|O�����1q�g��䞸_z��/n����3Vu����.�r�Es�'��x�r�&^�m;��x��(�u������b�K����
��{]�7�\)�'�,:����@�O1?g�h�'J�y�{�jі���X��Q�}�jr�t�3��v����x����8����<�>��ukE�l7�4�����.��;�'�;r��b�mK9��f�-܋|}�h>�Fz�A�f�����5��\�k=н���{L��T�T>��=��sT��8��w���"=���xe��/<�=��5����ť�Ȳ1�cE�=s��=���9ø]�>��� ��=ۯ���IR����<:�0-De�ww�7�$^���/|=�-/�g*��+~��6Dp�'��ca ��/b��o��ӨҼ<���`:��w� 5
���tN�TZ�����v;�2���06n	�#��}�X��q�6���4���Bz����q�}�˼��{��<cA�Y�e�:xv{pn����G|���&��C�� Z�zv[��io��d�����5��.z������*|4��>�V�����t�򷙸�^���6��`I_�r3Gf�Q���s}���E��e��
����&s�^�#�3�.�.�y����'۪'9ݫ"q��C�S��Û�� �t��=�Њ�ǔ�I*d�y{f,��ـ�o�j��ܽqׁ��=Ӄ�ՂE7o'v�z��3���<�''�+r7�p���g` ���bs�U������mA�0�_��jӒg���������R�� o����RU��'[�E
��A�N1Qu��K����d�!(�\ϖ�6A�=�;���_���O�������u��-�ߺ}s�T�E�(�|���N��M5BL���o{�ޗ��%{�On��Y��z�G�w�h��Î�w���Fb����_nN{s�yÃ�fs����M�7���v�z9�>���˛�=��F_)�K�4��������;�����非＝oޓ;ԧx�CK��	�n�Pʇ��S=�b���^K����f�/G���㝤n�N�qlr���9o�w�~P�*�.�xӲ�-�K;n�=���E�v)�<��<U#P���s����x��E�"�,'� �z��Ui���n��`����jW�����L�ǇS��)7���I��Mcr�V�ͯ�����r^�C�rYÝ��tt�|�
�z>�y�j�N����>><�k�����Խ��}��{����&��Wf��{M��76���Pr�旮��vh�=yk����~̦x��x���<�S�[(�f�]s�=k;˖��W���zg�k�՛�L�"Rj�ɒ��I±IQW�
b���o�핆G3eW��ǐ�pv�"m�^�|k9Sg�/:=q���[���>ݥP�D9�}:��`��Q�I�,��C�S���\|&���Uv/d�����N"���^+�ǋweI�n>�Wc~���Y�>
���ˇ����{;x,��7���1F� u��w����bB����;&�Y;!�tN`�̘~��yѷ�^s��=�D���|0��W=��<z�d��nv��Q���ek��=�:?.�|>�z|���=v��۵>��N�_��6l���ç������kV\�t��og`�i�7�^�r�>�wX���^T�[���-;%L鸸�r�ߋ׌�*�WPd�����<�赮λ����w��Z�� �����xM�mP�E7��_|�|)E��mXͭ�y�³����N�X�Mh3O���ΙX�8ϖq1E��ʗy������gs��$��F1��7��t{�q��#�$�f��M��V<��}1���f��N� �H�<���ԀuH1�5eG(��I���4���1�L]<Ww��`*�}��_�S�>Ʈ�3�3�˞��#�k������gL��{�t�z��Ȓ��h�{�wV,<Q�L_�Y����K��������|�9ۦ�3�w�������l!�X�����@�o]�V��G>}��5����
Q�3W�);6'�k���v�[�啴w�g�+ٛ�P�^�k+O�����r�El�����G�k�0��h��h���D��
�n�T0�on�r���Z��@����/&�Ї��Fݻ7��z%1=Y�&	�w/<=����d��G��''��i�E�&�{"���.y �n�ŉ���3��R}=�`���V,��scN��1�mνhWn��_t�Пxh���[�[ޓ�c��$�\;���6��WX�{�v{����J��P}�r|��(��.n�~�6n�l��ަ3����*o�� �{�nZϳ�}}�Vv�׽���ݴt-E��v`�zGu����p�ח���{���|�*�v�Oo�CZ�X�������ѧ���n��>i{�x��>PG������{�,۸�5�&A��>����~>>�]���~��F3��.�6��(Ly�k�x1s�g�;�B�]���������ܧ��0"ef�x0�÷yn��F]^�NK�$�e4x�P��ư�ܽ�����j���7�H{��`�c�7db��;��>�]���ճ	Z�����bq��k�E��]+�7��Q\��L�z���үS�x"�LY/��SH��{غU|W��%wۋpr�	9�ۏ���r<G4��������?$ ��$�ǧ���iڹn����L>�n�pA��fNW<��4���g��O$�p�4�+)�wv�(�*��,>�rU��;�3=�{�����S;����ɽ���x/m��zq���J�=��[��R>�3�%{�	����(Y3ݢ���{�j�78)G���n\����N���+�<�q��)�&�x�m��ڍ��;�s�1�l��T�(t�T1��K۞�~��6.oo<"><xr�5�R��':��%�na�Z�.���с�W����,���^;@��V�ݳ}y%vC<�wg�,4��q�%�=��������ʯ�zLV��ܘ�o����v�旄�~\���}��Ѿ�_9��C��b#��x�*<���Hz>���k|ig4����S��a+}��}���JeKA����=�߄�����ѝ}��}g��K�	����.����Yp{덉�퉟"��o=��^v�F��l��R;�ώ-��)�3�x'���^��7�L�K=�җ6���Z��O���ɑ��.q��t�������rv,�z<����>�����:��� �Q��>��幯In�huO�3��妕!$g}RZqߗ�q��b&C�y�#���щ�E�O,�x�-���ޏ<��P�n������;(Z�~Z(�0?)�����QGW<<@��Q���S�����Η�{�;�`���/x���}�ӷ��:����Y��Ǜ+<�S�wi��k�|=y��x�& @������5}G��q]R�>��\;��߱�E�F^^_r�2P�/4��u������u�!�;r���[�:͗1Y��y#A��l���=d�e���`d�J!<�˗N���m��wVC9���9��7�������Qc��Ŧf�r���,��n�|��^��,��2/A�q��կ�a��������������_��@�]FU���������tn�&C��t��=Ēݺ����>yj^�r� Y'o���m4_C��N�`���6G�k#�{<W�@�.��}�¶�g��9�=9�+)�Eoo�����˖��w��y��^�w�N?Z��?�7)~6eXt�Y&4+Nk�78?��~7_'4a������]�'�&�Oޛ	��c�ɲ��G*��yИ���X�S�Y"2.�|b��������s�/������R�.���c�s�JԽ���a�!�r;�z�=��t�����M׾
�;���{�������n4=�
rOw�I"Bf��ԫ�pd�.�*"e���\��憭38e�6v�J��>t�;�1��9��W��c�z;�</^)wu���Uu���V��"�+�����7���g�_�'w����O�����/�<�Y�֖�qf��j`%b�\�4/��y���0�pې&5�%�-�(]S>sѾB��g!��d;5R��z��v�ƨ8��d��U�.��M��L\Б�s���P2��
�uub��ٹQ�T�,�m���8
Qc\�ٖ�X��3Ac��y[����(�^`1xn���u�V�gP�Pdŵ��h6yp�ڙ���d���e��L�E,t�m%f���G(�^lL&4���V���厴n�b�Q�3�6�j�*��XZ�Ye��R��]�"���k@l�m�m�V&XΡe��r���o.�	䭬nGk�$&��0�E�/Z����)�\���խv2R�4e1�2��̱D���d�-�����Ł�|��R)v�ӓ�fŤb�6�k�����Yp�*��&�^�T4.2i]�pk��N��Sm���j�j�"�rVZ�S]��Yi�Ԗ݉k�c��]��f�^�A0l�Z�)�+�Q��@��mi�B*�Lh\�&�e#,lMfͶ��� FL����X�ɇFa�І�\k�ȳ6��Nne�b��@�B���#m5��xSZ�d�)ARZ�`Vm��Gj��m�MM`��`L��[���SCp��m�jh�XڶZXCmmK�&e�H�H`������r�{�|�v���R�kz�ܫCu��8�b;����[����5�#�#`�;��ڷm���]TU�m5I�uP�7���Qt�h$��
c�3e�c8��J,�`U��ݮ��\��͍%u�3v����0K�ᔰĦ4!3��#v!!f)fn%��m-����@C^)\�oj�:䄹�qB)J�d頗l�v��`��T,�ͳ�Ս��ô�1� 2[�
�kJ�9�h�΅`�j� Lh��thB�2GՌWi��6�D���5l��:���]���溴��-��و�Sn-����C[� BPلsk�I�j�Zkh8�L4k��Mn��k4^��P�n-���bP��1]�b�P56�����,n�<Fl�5pٳt�F���	{[�A�ɬ�MK�GF��0aF�f/f\Ǝ�Z�4��� �h2���1p�%4����n�i�=�'b���T��s�Kж�Z�W&�ͪq{1�1�Mn�6.� F���ZC���e��lk�1�]+ˤ�{`�M�f6��az�<�1�1rL�=oiB��Yc\�fm�n�aB�Vh4E��fQL�L��ame+�B�p5RSY[�k5%q�hױ�t:�rZ�����6�0��gJ��3�B��M6.v�XR c0��İ+x�u5Cc:1� M�˫�+����Z\�&*���E\w����)3h1�l�YA6 X�+.�ҙ�������k0MFˠ���:�Ҷ�SCk1U�L��f��j�u�UX��T�:�ţi�Y4��t6��rˉ��x����$)�;52B��@�.�:�,4��4ʭ���AU�k�JD���ٓQ G#���9�	c�a�c��mķXWK-���f�ٕ�)�Ќ ����1|,�P�M5��&����їB1�ke�aLiYTĤ��ml�Z5&��S0i�A[�i�k�4v%Fh�2�U���X�N0���l+t�*GXG9cr��a)^���D�4�\��3�쥔�f!D�0�,AZ�.�˱+��ՠ�&/R���]��h�5�Pډ�j��:4P.��ؕ�n1��qt��o +؅�6]�r�2HZ��m��B�[(�CJ���%�[V�,-�;Pvґ��ؘ����	IuĬHg2���5�=�p��&�"�Vt���YEUH���#KW�f��ͪY����X[��E���ֹ�D�g�(����B7`�u&�t5HR1 nf����%�A�gLK��K�[�\śm����B�4��煮��p��rA�h�-X�Ԟ��y�y�X����][ �!��iFm4�Z�qWG9\�e�3�i�:�ȭ4��E��32�uvh̗��ޖ.�ɴ��fpct(Ye���0qQ����d4�Da��5u,�YKh�nr�U@�lͮ�-�nqHA�Vg��������Mm�6V)	������[�F�]�m��r(L���*6�R�m���`��lp�`�r�V�Ŵ�e�nI��3��[(J&&�m����.��Z�`�P�8���Z��ZF�٘��5[L5�x�b3±��H9 ۔��:3r6/h�v�\Yk�0�cK��ffKJZL��8i&�3.34B�4%��� F\P�`�&��gF��\�k.ej��)D�n�6���ƍj�&�����E�7E"M0��is����KM�ȥa���m4�B�#��Zm��f�iD����4 A�	w��#��v�K,��-ųaJJ�FSK4�hY���{L��ZD-6� m�ݬ�Tڭ�#�ɦ4)V��Rm���e��-WX��9P�u��m�JR%�����,1 m�s	�o3��Y��Z�-��L櫪�P�e63�if�]tƠCj�f��`�pl�C����.���ɱ�*Au
2��v�,9h],vЅ�y�W30m(K2�k˳�tV�-l�3f�;�����̬�bDҰbF���l��j��,�Ʃ]Eq��t��gW�B͢���b	V�S�P4�Nm���;fcH���(hس���[\ڱ@�E�<M��2�:���K��Qm)3j	�icb�aYdc0C;��l�����a�܊Z�lҸ�y��rVi���Kqn�.�!Z�nx��YI�Fm^fj����&���]��mL:��&mAڐ[-���h��c�5��L<AE�CcjFf�m�C��i{,u����skqηb,�ԯ#.e�eX<�v�5���G3�;i��âKKt�0aJ�4�/X�*˱��Lh!��y6MKIV�"� ��a�f���!4튉��.�&���rJ�z�v���� �1�X��v�]\�d�7Z�0�Mjj6��̮8����\G��6�*�f�6 65ͯ�>K)4��1���c@�ƫj*֫u��W5ѥ ��6���W:�0�[�A�ڄ�-�Y��BT�
\�hR���ka�kY�Ls��a���`�c5�fH�Yf�H��ؐ���1C0vx�ٚ����i��̢"�I���q��,[�syk�����KMM�6U��Hj��5|/�஢��V��[+�&�;%,�]��Պ9ɜ�����	C�;�
R�#R:�M*J�L��`�D���,WK��jm`���Lǚ���0�
��V�]Y��D�uR�f��3Y��))�f�"6i1q�H�(�Nu�k265�S��R�^�6�]sqr�a�[��l5 ��҄en�{L��Iu���dA)
��:F��m^b�J;�2�MulB�h1��Sڔ��ݐ���J�u�d�����SZ��,�C0�7��rv�٥��&&�Q�ҁ����\��6�]T i�qS��cfjB1���n��M���(�8�G;bm̹\&�[
��:@�T��ntJ&e�At�1imb���8�!(b��YchT.3îH�#j���4�լ�b�5h@������`�ԗ2���f�҅	tЃ5�^�&p�r�7e�6�e͙Nf�6Nܷ�m�h�k����V�%���-Nڲ������axź��Օ.�\���X��L�Itm�@�5�T�����,��]4�'��h<0�Z�]qS[��ƚյ�@��e���:�Ibcdѕ�a�M�9�i�\�6�9��,��iFb1���r��uZj��)��CUۈ�����1�M�%.P+�v&y���-P��Xd3J[(�5�lD��@&��j�@i�ZcBj�C&�3f��W7Lllʲ٥j�Af#j�4�)Ŗ�9p$�L��3CJ�+Kkv�.��6�bV�,`Z6Tڊ"i�z�7.�A�]��8����ML���ZƄv� lCV[�����k���Ss��պ9gRiK��bܓ\�T�����8te�Fe69���Fae{7[�3M��{70��tE-����	M�uJ��(�t��f�uŅM��bL�	�3v�h�Z'x��mMui���e����P�$�K+�)����Wm\����[3��h��;k=�&*���"��4��Fn�j�qwdv \�Uu��M���<��ڑږ�]�1�0@f�Z�d���0��wh� ���t�h(JU��P	��G��W5��h`�3Z"�b����!��x��]	^1��M+q���	�մ	��ycY],,\2�	sXi`��Xp���"���fܤ�6RY�4MLޣ�2�i�Ś �Z���J��ۅm!K37V�Ds4���x�uht�U9b�&t^��7b�u�����s��fp�Us��-��ˆ!�[6��6����U\=��TmK`&Bl����ҵ2s6��T�2�1�]��6Qi5�e��7-��j���V��f�&Ҹ�#�3�h0ٛE�K3�3xB1f�3@j��M�h�%�dڸ���f��<��[��!1*�_.�y��X��]R���A{&x�����l�%�q��qZWv�S��a-����kf�˅ֲ�1IPe��e�T�h״u��af��nFY�X�9�+Cf&�X�A�Mse�5u媕q��]l��ۮAP�mV;!X1+Fjmk�hl��˂�+��h�Vf�B�HC�nR`��L�ܰW[�(ˉ��5�\�\�e���6�d�/�R,]wak)r��*�Q�f�ܙd���Sd����kD�,��ݬ�y�0B�Ŵ�̔n�@
LZ��ΆI,-f��i���v���]��$>��	q*$�V�ΣPdT�Qz�FF�ʷlt����Ǐo��۷nݽ���IQD�AP�*����{�n��ߵ�4T���r%�ddI��������v�۷n��� � n5� �H0ۑ����CW�r0kr�B�����Db>�WP��! �
��P����2��mr75�y�`��k��.�]\�T�k��ދ|p�Q�ݮ��tCRbŮ\��W�ؓ����寔��^h�5sn���5�Hä����e'%:�!%�'^��Z^5Yq�̳�qG]�w�t��׺����c4wn�
�\t�Iwe�w]�u���q5!���I�4��w�{ӱPK,���q�I��.�����1�۰"Y��WX�j�;�
J��m�;$�ιe��n��*5ح��x�EUM�jCsK6M3��[V�������:�KY�I�D�"���՛s�R�n1ka��0�٦��� �0�
�����kM�4T�c3�C%s���[�u���&͜if5e��Κ)*jK3na�,���l�.��Ech��3X`�e8A	t���m1E0\�d���Ԇ�-�T��c�9k4�tm�Uf�0ֶ�WipYtD�t�)�%�$�ʚ�-�鰅[a��`��F`x-v��S����k,��^�;CYC+�P!m38��8��r.Ë��'932��f���Y]u��Ufuι�!X��%vv�]���@�CRX]0�˜jh�n;,\ki��2�����2�!+�enK����o�:�Y�!Yu���8cvX�&�obSc]u�\ƪLF�\@:�R6�!)j+i��@�`Ɋ9&�b(D�Q����)+,�v�冓�	Ll	*�C69p,E�*�ѽ�{\X��
R-sir=@Z�^&��uv��4��-�<2�շn]Dasv�3oGp�ƻnBm����j7��P�d�ٖ�r�cEvvز�K��γbl�`!c��L�rT-���H��7�k+k) ;1�[�R�cP	��k��8�:]j�f�n��|e�%�՗�5����l�R�+���ڵ�c;4� l�� �\ufb��4�3S�m
U�U��c��+�2�Y��Y����;���U�8b����<|�_&FM��l;MC2�A8�.��0K�
b
+zݗ.�5�EjR�t����J窹���t8��ز�e��&-���Mi@��榹��z�lɠZ�͎%k�Au��V�S0�(Vj�Y���\5��+����i�Wij���4�XF(:��e5�Ř��u�ww��זz�z@��Q�e�[R����Ă�!�b6P������R�@��iz-�XØEW�@e$hHV2�[b�iX�8!*0 <V%��m�a_d%���cl�e���/q�{޻'�{��r�Y)+����,"�X�� ��Q���m��Z�i#*,�|��g�����'�l��Mfv��V��VY[��e�9	��s��dv�����n��6՟ZozY�=�u�,�8ȝ���ʰ5[�Rp��ũ�-p�g��'#�/<嬌غÕ�6T��l=X�gI��i�鸸���*�����_[g����0|��!�Z�,Mnh�e����Sz�:LU�T��V�I+8(�C{.�&��K7�Y���r4D[�m��qv50ů��)F��]�ݖ}�m�;&Uı��׼��ӕ����lz���^)<�([j����I�V���4@$C뭬n#�c��"�q��h�dt3�;Λ�?=�>|=-��ۄ�GwL��9x_O�o��i��׌�QY��$�'�Uf5��N��k�XFV�i���6�c�Κd�:)��a���0�FM�4�lM=]4��z:��E���Ҝ��э�??Y{T��\�8����;ie��d�����E�Lo�(nK599L�+�㸆{-�z��p���i���͑Y���e��-s��
���x|m��'��C��{򕟅���,�-[���Z�9x_2є��k���5���[����m��k��J|����"5�k7�.�f懖��wx�� �7�EY!��rI�t��N��Ĺ��SV#2��^�B��W��.�5�����ٹID���|�_��m�N�5�V핛Cr0�)7Z�fh�h��s/fKw�G��`����L+#?N�+*Ni}ܽ|�.�2��M�8��-ډ���շ��$�$��$�ա�%=��.�_�͛l�w;�;�
��Z3��C.�5�H��qT ��~^'������I�������^�Ogp�>a�}=��f�[}���7W��E�Hs�{�w8�xn�|�/�/� ���휍9��Z�[S�O���c�r�*s�V����]�H��"c�N�s՗'5�w��gJ�_�Y0�w+ĩg��z�t�z�>K�ِ�\VR�el��q�(8,i.e6�� )�pa+�m��s=�|~	7�7�do�VM����GCni��7�'����I��?����ե���;]D4q����˂�
�|�2ʍ���� >�ass��y'�Y���M'$��O�%^N�2�����{�p��L��q���}!̐�o�yʌG]#�o:_��wo��-�˻��!�e]�Q�w��Iܝ3t2�+�UeO�nj2��#�
eONt���M�k���fyy�2R4b7lUf�Y��A��M�gXz�6٠mc��&I:J�8j�k#Fb��j�m�[��YQ��l�$|�$�&o�e��?hC{�����T�iZ��0��ڵ��te�ez��U!Z�	���<x �e�Y���}"q�N��E�ͬƊI���Gt�wf, ����$�Q/Z^*��pM��
��ܻ�}qQ�Ww�ao����ڼ��Ԝ�2uY�g���r�����[��^\�KVFX�Rmh��Q䓷�LL$��T�L^3m���t�m�I��*��{�Uy��-Tʌ�+S�=�9*s�M�v�뻀.��l�aV4�V16�b��}��Ww�ah	�I�M��ͼ�.����K�=�g�z�S���Q
>��乼����L�w��ON9�������y³����/,��{ã�M��0��b��7`=�`�oy��z-D�Lsp�Y�Q�6�&2A9Kp�F[�]v�ḓ�xV�6�NH#��9L^���YtAF�t���n[
�[�EM�P�&RRi�÷1�in��a&v]]�m���2��08+ �4L:���u�CX94�k��5Zָ�ΖR%r�mYf��:\�m���u�1]��M`PpM���7�2�Z!�v��CZ0nX\����|?w����˷7f���5Xյcb�L飈M.�ښ<Ev*�e%�}���=���ݰ����w�V�\�Rmh&i��b5���aw��	@�U�dU\�*�����Wj��k��Uy��-T�N��J�[w(Ci���]��cy&$�-ͷ6�!���T�^��̫��0����U3x��U=�r�v��A�,�zu�T��.��!j�˒�&�*ol٣(nz�)f��g�X��&�aTªZ�C�A��S)�cuM�>^�y��-�M���ST�m4g�^�w�r�~Eq'[ƚl<x�u�meaYD��؃���j��1vd��I�|�y�t���?�_�MZ��sf6D^]U�T�0�;
�j�K֫oU0�$�I��I�Ą5�
E�������<d=&�X�� k=�NN�(E(f2/V/��d��J�U�ԩb_a>�����1*�d-i<eA4�G��e?�q����%j̛��&��Q�m5W���Z��{R��a���MT�U>�E1x��s�[+Z�n�,̈�L��]���g�u�ꪵ�żQ2��g���oU0�;y��!�.j�L��g/�vl]�~C4{;N{���}��(d#�Һ�ו��S�׹m�م��W%�M����©��)��͉�`�@"Rְ���9-�X�rѥƠ�#�G0jD..��5h�;�o�[�MU���j�qfdER׶�:Oq�(iV�@)��xUUUS�SfM��PX��6v�r3fE�\�䙭��o/Rt���V����ɳ��3���wlG��c�1Tj.�ƾ����l�fgU�S�utL0�7n�s�%��jA�OYyҥ�b�"=��
��1�d^T�8��Ҿ�*��x��?��3��5�ׂ߽�/���S� ���_�8g�'1""�g3.��v�Y��Y���h�$�^�8�M����~����=���?wyNsԡ����u���;-�J��5��0�oU0L�#:�����{�~��ÑIp:����Z������Wl�Iu��K1��?���z��ɱ�,ɍ����7:��N��{���f�<~��s�������5�kS�v`Q>7�<��/r�2!U�Г^.u��4T'���ˀgUmcU5S�	9o�gEfV%��"�d��Z��OP--�H7h�J��P�I�kPL6�©��-ɍ��WFn��7��2���ւ!+ўl����Gعi�>��]yߙ8ff\�/q�2��rC�P.^tUf,�j�-YS1qE�L�i4m�QR����g|�j�����z�ެ�]S�׸��e�h^��fd«e��0�+��b��f��~�H'b�#�M��s!k�X �ñ���!�+�ft�c��
3~q��O�׌Sz�������ءn�-c���Z^bRI�tC�n�7�S_�Rvr�N��G]὘��L�����U�7F��7������y�[�>Ul1UG��x��gMk�>3m�VQ��Ƌ��ɋ�e�	?�u�Co�L3�o�6��pj���U7�&�726([�嬘>���0�E���1y�M)7�5Sv+F�N�N�:���ݕ{7h�ѽT�o>�T��zh�PxY2	iM��&*Ci��bұ��nr�N0����{�"���o:;[<���c��U>�����-d,�P~�ی�ڠ���+gC�y�f"�;bgm��KP��LzE�|<!n�9����z���ٔR��̃kf�����ڔ�ܸ[-n�6(�nI�Y��ј�V�ـR��6����7"��)µ4n�E.����a�5B�42���s�M�4��y�e��ۙ�%��	k���v�P�� �з-�v�љ�$*��8q+�Q	�j̲�F�LT�	,Cm3-��%D܄ƻU�D�1�� ��Pl �ǿ߂���,[?Wm��g,4��Z:�]ZDԮIkS��g������M�T�2/5^4^�fL]c-�͚�������x�!�����}���|����-fCz��%f�c�+
/-,��y`%7���u�O��M>���������s����?E(�V�%u�ֆř*�ѫ�ka��ژ�`*���ًD�y3�Pqd�E���S�͠�oVfL*�u��]Eݦ}����-2��`�,.=v޻j��r����3o��=��u��=^��L����$���|�=|���޳�v�>_��ʹm�͆�ʳK*rU����e�t�h�u�h�M�OS�o�ST�Ͳ�گen���mъe��D�*��I�T0M�U0�i�̟�^�3�o�4�j���Q�^�c�Ȍg�v��2C@݈k��-X�!�R%��!�X��N�$���"̹G����d+�7�{��.��h�N����V��C�#�>_Z�S�!��9����]N�eK6�X�'b¸̬�����JaT��d��e��븯i��,k1��R���ܙ���;m�����*�U0LR�v,.MYl`u��I��vºq�r��j���o�=ETz�*d㙝#<�=]������٩L�[��HF���c.��F�!��T�UL�]Y*/y��ϻ>~Y�՞�YڽO{:�+�ʼ��b�ST*��K ��U0�U;���Vd9^U3acy�CPܺ���EJF�M�M�y#�%�라���{��ք����g+9S��Q��5B!����X��͑�&�[���1佛�����u!4{�sm�$���=���tΛ�
�4��Jf�ƺ{�G�S����>�}��n�w��ݫ����3�������[��؎,���G�ʘ9&C*7���}�������4�:�Ĝ�έ�VO������{_ur{|�v��kӖ�v-�!��W�G��>������=�z`�q�ꔐ;�_����n�鑒�m��<�U�ײv�/GK��яz�7\�{����v?m;�wc�V%�[�Q�3���+�=xf�ڗ\]�p�l�2�d�C��(Q�0,���s�����ɵ�O������>���؄�چo�]��W�6&�w�K�p��=����ӥ����^o{o�����k�8d�A<`��v���Ġ3S�j�P�X�hώ�G3z���{j<������w��b�}r�}��z�t��OEϷU�����a}���Mk/��{�Ud��ئ��3�x^xv~Ro�4ro(������{��C�۾>�٩��wf�ڈ��>6���g�7� ���>�u,>�>�q_2	Z�4�d��}U�=��$�N[��VCS(�����r�\=���>�{/[�͖��)�+>qا��A���#_6b=A�<���b��c�4�zYUS�p���k}�=oB ň]�m\圖p\��xd�Ë=%��u�v7n��4L�'{��aB-7����H���J��<��b��4 ��ܜ���y��vGwZ?]٦�ouؘ�s���w�\0L�;��9p��>:��$�J��=:x�۷�><x���nݺ�i� K�UJ��N�*�)5Q�����_V�C�P��ZK(l��s�]�.qLt��i����>>;|x��Ǐ<�]�.��+�vl���k��﫴��Bs�WX[�hhw�J��g���W����ǜ�`3yۋ�^O�/o#u��4����f����r�{���<܌)�.K'�z�����Z,:�<�������b�~��۞n�t;뮦��2=��]Wz�.�(*\�ss��[�|���疹����N���Ku.�>/^�[cD���E�߮ޚ!;��/������~+����^��g��^�͹汴l�AWt]Ml%���I@�	��ħON�[e%���:xR"@�\z'���$ֆ8,;kԐ��:�����D�����mSM(P��tg�=��߹̶������A�"���N��	7���\]�.���m����o�����v�qW�*�9�����Y�o�4޼3�s!P���24y��	LcOy�.�v�A�p�&`��Gh V������_N��䢥w�s�� ��	;������H����=Kkt�,XaW�(����%��K���0fhDԆ�m�g��|	�g �����|Rg���6���^SUU�xŷ"���R	���YI�	�Y<�@&�i{h��w�̧F�~�x�x"58������lV�k�Sm5����w�N�6�ݰ&�ヮ�f�{M�= 7����'⊏4�o�x����n7G��A�s��%+|s��<l���7�ܣ½,�z<�ȇ�*Yχ����ն#}薠A������L��YCE��e�5M.o�q0^#���g4��,cՕ
�&Z�}ӈ�{wW��s��fHw�ZX@����l�����fE�y�c<�U�l4��cfs�b�K٫��ŏY�/'}�����h �������,�Qp|�|�B�=�L܍u��
�~���JZ��6�7����o)5"��Z:��7BLh��ǣ��j�q�!��.�	h1a	fu���*Zjǩ�ƺ�����4
�s1L׋�I�rI��K�czw�+%Kh���R�Ƌ���@
�
[޾oO��a8 ���8�0z�޼r6Kg���}�l��A9-T9O�ݗ��T�y��&W8	4_3u��&^y\�w�Yl:兑!��HM���$�paor��1$��bX"�q�n�/-�{�S ���v��I���5�{�t��!�%�̢�{�0�ANM ��=�loN�ed�����L�O5ގ��8>���o�6��Q�W�J7l�Y�ݷ=w5OGe�����y��u��켖�����0>-�����E�o0d�Clu���N�
<V�=���;����qvׂ��p�s?7nms^���s>u{����U����{Q"U������-�7T��!�������J��O侢�W\�c��{�ק^�gN���??�+��l��A4#[%�qQ6-�n3`���-��e��ڤ�46	u��BJ��4	0�0ƓL��[�f��i�gc\���
B:��Ļ@e�6h�[V�$�dJ�à77�%٥������h&K�J]C�B٥ ��v֙�G@�P�b\6�:���.���Fl��Xl�\͎�ܳP�(F[e-55l�aG"۳��G�]�7�߿��/���ոûA���X�6��+me\�+s��"�u�	r�ŜL�`���d�A���?�d|ʭ
��<���bm�������&f^r�������@��r	�f�n@b3{��k���9��&S!�h�Yf�P6:;w��h���9�	���rp�%���/g�d��8ޓ���(�&�x�ͭ]wkzP���:&����d����c�i���l��尛ݗ�G9�ӻ��Ժ+8=�����T���a�L�qU�U�q��Uw�_�&� ̳���~
d��ib%�^`�[�l�H7l�,"�έ�h�ǿx+���C�k"�)N��6Qs�y8rw�	�W���Q{��{���� ,��+]�ae�	m�.��*B�
f	4�[-ja,�y'��;��r�����Rj��W&j���0��1�aw3oM�髩��5İ���*��`W�O��$�	E/�!���쭂�~
���xR��*�,EKN]$���O"�/3���7f=��J���2��։aW�b��&�NE3��a�~4)M4��(��v3���*�*�~5�C<��
��	��9>��C��v<k���������:D���8�"��Rq1��L�"�LǇ`�{]l�b	*���f�z+�O�0T�p|@M$9I�����D��-^�sX>sQ����}��/l���u�R�1����0pE=S�62ֱ����4;���$���>I��oCֳ4��s/+`�8�3�^���ݤ+7'�<M]�m����6�|�8 ��y����x����V[]��)+q6T����	��W&�l
�S-�3V�J3X��z�w�{��p�r�.A	8|�@�����U��8y��q�E&��vCN��\�	�s�v<����|��JM�Y�Xk�L6r��.g�7M�*Y�=an�6��x�s�r��z�
(�um��c��˹4����MNF��.&�e�u�h�b9��x��왳ݻ�MJՉu{	(��#��3���痷���I�=�(;ͯe7ѭ�m�� }U��9'�gf������뼺��uo��ƔZi�DP�n\����s�3J�V�7���f��6�C���%&pB)�E�n뇖gv���>������N����6q��=���\<s����㇙�Cr��L�)=�m��Qe��V���Y$���s{�Qh���:�1�.X	n��4'����eo�8�&���!&BO�u?��l{H8ϷG������A�m/���-��R�Uv��B[�vSs��Q��ާ�_7@��o�I	/D?���	���s�3YxշG�a��T��S���O�?a����$+�����s�W�j{!�ʲzس�sGF7����A�p��P��=�wyaJ]�|6��<�8!-����u�'@����o4�AL����&r)6v��y>ݍt�գ�+C>��}���h�gM�1�\���H ݸ�>�5��U�d�%�"iÂ;��`�t�\��1ș��j�� f�φV��Ѧ�u-)���	�f{�˭�˦�v�����>��/���XkK��|=M�`��dΙ�!�b�؂S&�6��">�i�A.e���&��۳�O�N���?�>IßO�I�~W�g �X���-�w����E.���g �poH> ���Nݞ��$/��~���^�~Ϛo:Z�)�eY]�M7	�:P���3m@ؖ�hD��6� w����w���e����]���vX���z�م�J�/�>pp��Ƽ8��T�.��L�`�6�BL�p���=1*��7��c��7�\���:��\��1������M�T��탂�>w=�=�N�Q��C M�e0�i0p)8s��9�8�͝�v=u��>k�j�A�o|s�����@ �Nk��.�Q�g �]�s��=�f��A�`��5�A�&v�A�e�v�aj�\<���;l��R�j��f��X�<[��9n���pA'+�6�׷U�ݾ2�8��j�y���e���n �T��	�o&pA�I�U�A��P��B�!�zuPf]��J��ӷ��9�u��4ەL��MF���k�v��j{܇Lwd6jBC�d�؇I���f�v�&�'ru���jY
��ߍ*Mq'N��|ߞ�]�rL�60���褢�
�YcW������R�'�����PAN8��5-�V�q�v��U�4,h�"Va�]��Ď����HZ*ut�VQ�uY�hgfTM�9r[e��6fGDn�)-�]����H���0��\��)l*-��:��ݲ�(���sMdH��� ��1�v��.���Xj��YXݳ���9������<����VSb��#[.�ǚ�Kն75�G!4�}��B�L�'�h!�P�9e���[v]��写��#/��ex�Y��ꛛ�-�{�ɽ��{��h�}�d"5�r��f�� oŁ�`�[�����-QK�x���c8>>�>mr�o<�y�[��6k,���\�Y=es�ZÖ�m�<���u�SuN����;�x(���+n�� I��6�`�����S�Y���.����j�9���!'���Ӻ���ya�s�o��=�k���+��o2{��)<!�m��}�nc��'1���'O�ن���D����<e��y��Z&�;��L& H\�q���c�dZ!�Ɩ+�kbY̢�L]e�f�[FhiA�D1��A�Mil먞ߍ��:�tW�K-�{��-����r�M��i�5SK.�n!�!CT=�MSg�t�g�6�C��ϒ`�!�I����)���K�~2�ݷ-6�A8엣
�BP{%I���^��Ͳ�;�^h�|F�н��������+�sȣ�B��LY٪U��zկ�{��o��*�}i
i� �wC����3�?ە�n����������. rq~0n��f]Un{ޠ�d?N�����mӺ�N{U���ʼ��4fSrǣ^����e���O�x�7��ÔQp|I�x���ƶ�Y�f���[y��n����Y��;�xUT�����ޙn���9c5���f"�z�Bɜ� �uno� M�Il�E>����]| ���-����:����x�pG&I�����4�{��m�� .}?u�0a��p�d5��S��T�)`6#�C�P6eHй�\���M�w��~_�ĉ7����Z�/�[��y��1�o�N�*����T�ue�L�C{��ot�nI�8���6���Xg��o8>4ȇT'rst����/�0��8 O�ca�n[��:'��)W`�8^a'���XY�E�4MM�f2��sF<�N������UWF̵OU=fS�Uډ&UT3���T�_??n?T6$�_@�w-�wֺ+\�_+|�j�_2��~4��4�"A��{�9��]{�������Og%����݅���l�{�S|����o�i��Bn>�jx���8ji�s9����-pc���>>L�g=?F���P��	<Qr�q,��N(��$�H!&�m��:���a�&�)��è�U,6�p��SG��g���8 ��X����.bGWf;��3fX�m�ٰ`<�Sc.�I�[if�bh `�5�K<H���0&��Ǜ����2d�����[�GD�r��3�SG�Nn�d�)0k'<�r�0�vYuv�u�4i8�9Z;h`m07�����تL-�`8��&�Uݼ�q�I�b�x1��)�!�Â�'a%8� }��H�wƏ�IÐ���d|i�j�L����#�h�UT��m��x̳��md8)3����a=�)�Ks���{�h�7�{�Ã��z�{�5no�����{̛���r-��M�Q�wji�Q3[����I1@�9���WG��B���L�����h���ϡq̃����^���E[�ք��y��n'��{�ߍ(�M4��st|a�,a�a
M�&x��"��Y}�֬ @�;h�[1�A<5��c���`���_��D�=B2�F<{�=V%���e^�Ck����f��Hn��p���M4tha�$W��._ņ���I���"N��Qy:8]M,�n���2�RhǊn����������ǀ|7m�6D����r�zL����)֏S��e<w@}�y�ꪮXR��5�q��#S�#+�\aT��|��C�l�3Y�2#�4��k��Z۪�:��!�B:r_~Ђxk[��������g$�I������㜸�T �h ���<Eny� ݰq}aK�p�u���w>�g�҆]�9ݝ���@e��)f��RRo�Rp����e���άM�u-��uLUu�Y=��	�*�C<�L9�փ2�$Ҩ!=|�E-�.�t\���&&^J������ א��K�Wn��3��l���r�9���K�}���uy���lP�(X�e��b�	�US촯(��2+�;�b����D�ɮ�{����7nҁ�R��{����C~�����1��~��C��܉���s@��Gp�j���垊˳�|�a�9�w��K#M���^����y9,�����~�����+�E�e�� �����PA�ڧ��N4<������ȉow�ߥ2�,7�]�j�6����Un�.j^s �'FѰ8W�x�[��H�~���yx�l���x���.y ��yذ��C���=���'�&{f�(�9�:�x���a��<���+S|/2�e�{�=�%�kΨ]�����,r�0�4\ei���!��x罧ؽ;[�1`��p���ޞ)s�=N���t�~>��~�9�k����Ipga�^�`g{s��3G��8��]|2�}�Y�{=��b[��]�Wv1!���L����2�|<���tG��E����P=�!��x���s�E�����{�з�����l^�U��ɻ|��Ѳn<������xN�=Vp��ݾ��Dc���^��ϸw����{�*�(��r�g��s��>�r'1ޞs��L�E�S����*�{i���iف���F����5���l��q��{ӼU�� ���]��z#��F\���^�y������c賱{Q��v���3�5:���NJ��yy��@��I�Z:0���������.xwUj�����k��+Iݝ!�����/; ��8q �BA��eih�{u��A��<�>x"аiAi�:�v�z{���{؄��P�0��7���)m�z�F��	d�A`������;�^�zm������o�<x��ǳ��[�y��~���o(痞Q��Dh�
�T	T�_��ޞ��v��<x��Ǐ�"d�Rp�h��T�J�����wo(�y��r��]k�'F��֡kJ,�X%�f$�rLZY)�I%�$��M�{�7�=�;��}W���cN�\.r�y��v�߽x��Ѽ�y�̻E���r(ϓ�w7�ۺ�ƹ�������Q�N�L�o<)�������Ew|�����:k�mw޼�۝(��܋��˞�o{��-�s���n^���d�y��̑�����u�GH�{�{�[�|o��:2�^�
P(���?|���w�<�5h�ـGg�ʼh�du�pKW+P�&BL��-ٗ"���ttW`ұ�ipe$)5 ͝B!z�df4F���R�r�̓�`�]�,Z��5�	� ��KSa��[e�J��sJHG`��X�jm]��iRZH�:X��e�Z�sY�v�4+�#��D� "�3�]�g0�cnm�A�����ŤM@Uce0ƶ�&ea	L��m��<��`��_,m5��Fb�Ho"O<��ұ̤m�u������؆�[��P�t`�ͦ�(- Ή�lZj4�.�s����+[n��e�5ңbs����]�����OmdF&�R�v�SQ�.d��6Ur$�] f�cٷ6Ҙ5�X��5%-�V�%.�#��h�%Բ̘Ęl�h�l4��1�4���\.��k��������*�/1s�Mcɥ0���3�q���GP�a����(�����C���3멜�hҲ䔭"���\���+v!L�0�Kck4!-���m*,��2���cB#�G`��f������l��T���Se�[���06��2ܓL�Y�l������M�4*m�7W6­q.�7R�êg�&�e��LM�K@.��� ˘�n-F��͢98Bj��G�B�A]K�y�7��5��D�Ʀٺ�a�^���J0L-��bn��0�,�SX-��#LBV���S8M@�*�k��Y�2l6�Fh�͚R5��fQ%tF�3f8�q�9��4��.��iF鋞���e#��4��\=`�ۋW.$b��9�n�-��*��J���6�v4v���L;M
gD��</�/�<���νe��P�Xdu�A6X��a��ͥ�#����%x�^�L.�`uu����i��ƨMۚ���óH�]yc�M4&�7k�56��;��sVإ5�jd!��u�*@t6J��3�D�c1ik�����m�o�\D7�,L�,<��x�J�؊��@�SM ��wԝV��X�Y���5U��t^��7T\�5�Q,͎L�f�\��R��6��+�!Q�m��+firسX�iH-��iir�8��[�p�dA�uu����[s5�X�X9f΢ҵ2CB�һA�2��в��lc5�ʆZ��h�m-qth�FR�X9�K�a�ٺW1��32
�`�j���u���Ԙ��3��pi6A+3q|$�ܿ�g�Ie�k����%�qC�/L�Z�e�q%�6Ƃ��=�Wф k��=�-��\HM�7�����46.�kxS�R��Ѵ%4�40��{\c�Wp�9k�t]2�������y�X����x��z�l7�8[��^7]� }���M�)4󰌲���s��OY��9�yEs���*�Nr�-Z�m>l��yK�Q5�&�W60�:�ϩ�'��'�&	3���W��䲞����v�,���_ŀ)3�Tn./G=q�1���{�� �`�1$ZG�wju�K��V�����7��Ci����ɺȬ����f�R�Gy���۶�|1,��mg�4�JM�>i�N�bl`�f �,	�fA�3��6m
Z%֬#5�μ�;[[4(`�X��)\�n#��snX8����h"���^f�z&�d���l�8�UE1c@�����7�[Y��I��g.��v0��K����n��:�3��e>nnx/3��)~[�We	��زh(��w}�;����Z�;�J���*w������+Ư���s���@	M4 {^��
�pA��g�=�篍1�\��\��I�c0ǋ�k��
�w���$���"���]���җqG�1T()˱�f�1�����`�탃I��T�	H>9��T���6ӽ�; �iƐ�����7;�3}=\�R��60�G[8"�
a��f�o#�Áx���v�Gy�f3�A9�ݳE޼[�MK;UQ����z�Lgy���&�+�9E��W�Y�g������1��7=����Қܖ�̷[��viLTy�e�l��ܲ��l7�l#���71�J�1�qf>ݷ Bld�����=��4 ?�ZV�r���� ��m���F��h��"�b��f�no��+VRY[���<l�ƧBH��ɮ��.w���)����E�A�M#�h9�2�9����CI����(]��ا����;ߨ�e�~%^-�'2o*�[��L�Rɳ��Kǝ޻�:��>(�Qi��T	Q��|���y�����~	���"�Â�L�x��@D���نw/�0G٠�����;��"��'���_�b�~V��^,�9�e�O�s>YQo^��j|Đh�©��Ѣ]��p������줲{͍����l$v�tȆx:�R�u�p,KU�_;�A��mֆ�4�14ԁ�"=LfQ���D����9&��&=�� ����-���I��&)#�״��hN-w�m	��[� �
?���,�C�,� �wl��SOr-Bo���66���s*�xWRŘ������E��k!�I�^���l�4�3�D�v���C&
(��X$��܁�h�!�*:k���Y�k'}Y�{9-�=�a�Q�h��.���Zh�F�u:���1��87���8d��̬ښ�(N.w����`*��f����
���U�
|;{�5�'?h�9�D;�駩�`�+˰ض���\C�M4Ⱥ��	��M����ǹ�Xd�< �}�D��E@�>��\'�l7��Q�9	?]��-w�c�O�D��o�[���%�����LK9l�&rvI���Ŷp�و_`����U�-�4��vѤ1�3�Z	V�Ye���J4m.N��x���F3���!k��F���\8���͢����d��x�M�s\%U.͐d� �N��z�2!�i7���FG6�uct�6^��SAJ�nV��P�\�q0pA�s��EC������k��0�����	0pB���ȇ}�h�1dN�?um��V,�ˎV��ĳ����)3��Rg"���b�9��KYF8�f8_�$��r��;GUv+���c<l�*3"!��ê�|3���щ�d,`�4���`���힎���cͭ#^�N�En���X�\��`+�IE$��v��mOV���wF��q��,꘳UM��!cm/ �����w4Z�`l���;�{�Iy�D�����5�� K�Z��4ʩ*B���D���iN����~z�>o�^S�!m�5h�*0[ÕD�Ƒ��r�v\����2��U������ݥ��ْ�2��6`�X�M�Q�he�q	�\���Ma]&�b�qD��bR��Ĕɓ5�2�j���WV6c���&��+��`�J.ט�S��u�� =S3X�nf�ꮣ���Etr�(X�5�0t����R� >l�)|!t�5�U�
��O�y�k(�n�tv�G5���6Xb:f�\ٖ�ۡF^hxb�"F�_8&��"=��,.���!�uk_Owt�N+�ˎV�F4zޙ2��J�`�1`�0`���Dp`������7t��.A�p����'^g��\����p<l������%�\[P�vi��P7l��i3�>o2L�i ����R朕��J��ԭ��b�6���q�������Rp����S�=t`�i�����?��Lef���˺̹�m�>�o�����q�E6T�s�W�q���j��/Ɗ��.�_5]n�Kiڮ�#y����'^Z{�\d���rIl��98q`�y�R����K���\8�Y����P�~)����a�t��ڹ�	I��3 ��Cmn�Ί�����e����^�����̩��Yʭ����60�G�D;wGNd���Ȭg�?��Æ�0�okP�s�cŇ�aL�����T��ˋ�Z6{�����{���n�N�k�= Y4�()yOQK�v�;����'�M�,����������w��P�"���!M4(�9ga{��~�=����f3.�2�U�� �kL#�&��v-�.Zz�0�W��d�p|s?�I��o:N�ŵ-n���ed�R[$�v+|��&Sp �p�$�p
L��D)�]�TN�d�wCU���&HiP�|��̩��[�h�����s{S6�#]��ka�� Q��X��I�QE�`�$��
zi�.ek;I�9�ͤ=��ޝ�n�̻�ʞV�A%���dC�L��Rd!�=�l�u������鉈SJ�X])��<R`�Kc��T�i7���D�Wy�0}��>0l�pAn;+0d�}���'�˜^[K���A���Z��)��M �
L��B7[�ܧ��ϛ\����r��JM�ګz惡x�1�;��g�o��@6l���GM����P��8\��%�̈R]3�� g�4ty6��¢�"�T[�L,�R�d�5�'�RY���xGV=� ��Z��C}=�t��l�y��FG|�u��o�&M�~4�SM  j��1}��Ff]fT���2�"���� �����,�0���yz�g�n�9$���0c�}]X�s|��t�pFH��]��;:�"��Y3��{Y��a3�@)3�_��I����)5�ǌ�v=���r��4!���su0pG&
(��	0�3-N2���a����k�	J�6�fʌ.�
9��p��*�Ѡ�~m��e��KI�S�,�o��;���;���z#/.��y[q�03�ݲ �r���&�*=>p|R`�!Ҭ�u��SbE���ї��g��Obi��T�ӆ��� ��x�|{���3�����҉\�ƫP���Z!y�[S��w��A&�|4/y�5-�̺OsJsH�/�9�oj`��+�8(���	�9	?�LM�pnn���2`�"�y����6E��c�v�>,�˩�m�L�8!�����#�XpC�	�8��U�j3�����S�rh�(�Ɓ�ꃍ���y�>�xB�H���w4�ˮ���;�u��y���� ~4M4�/+�|'2����Y�����T[�E�,�*|�����ݳ[f�6�?�/����;lObi��7� ������I�!2#�����������>�S�)2�X[@��O)��R����+�k��F8�[�f�:�Q���~�<�p �l!�I�������wW)�(f.��!,�Zm�[�Y�/o��`�;�O�p|BS���=F33����Ȅ�����Mz4wo;�ɼ��V�A3,����(>"�؟(ґx�LK`�T����Mw�,![�ٽ�iovt���s��z���g~ڬx��;���Ð���	?����J=��]c\	Í`�._��kϒg��V���2%���q��L|� ����JFW>h����E�}$�r��`�n���Gj��;��o:Zך��X�.���{����pA�C�v���Mf�kdVL��H<�(�~�A�{k6\�OA�?Yoqo�w�V���|�t�ӧ����{ާ~t�>SW�=�t����,J2�]�*���!��J4�*������R�C:��H75е���v�WZ���f��S4#�wR�a`8Hͤ����<'���[-&��J��f���m4�cW+v�`�!�fJ��K��2��5�a����d,�P��f����r�p�r�ʎ˱�يk-In��D�5����aژ�"hf*R4%��⚓gqN�]
�.\���f�.�!�̻A	p�-6Wz�*������M,�Ѓ,,&��hm�bX\c-$6�W\mˋ�6�����6��>�v�pQE�)8p�{qx_���T�Fw����V�7X�s;�[f��;a�.����.��ܭ������K�}����M�
�<A���S��3z:fD�8�1�8�0r97�Feq|z�n�6߶A��G��=�.�tQ�[l9VEq�S���n6��@�Ň�d�\�,n��r���M> ��;y��e.�E���m�Ɔ뷋���@I�]�Ō}3S�����N���3M�#~�!�t��r�5�֞�+u�a2�.��-��s=Gs\ftlL�Xqhc���')��G'QE�)8��O9='��'�>OٷX�BG:�-[1�=�f��e�G
��R��y�����D�a�8\���BW�md8�ze����d�dO,n\FS%m��{�q��[I����L$�R� �M�l��^�T_��1~��hqk���`\b��`��8�w
{��3��=�n�L�^�²��YB��<���u^��t�k޳���S|� ��hV�hJ��;�M˄���\X��a�y��|�Ss�p�pA���BV�F���J����gwY�E�&pc�$�q��/��X�P�}�"VLߥL��eJ�a��l�ܸ������^���y�G)��E͐}z�|l�S��Y�J������W�<����p���#22^hb!L���$��)0rIÐ�S�gnl�g��"�ü*�۳�/=8�;���|�Y���N�0d�r����%b\IK4*E>0[�Y�`\�tx�q�l���[M3��6mc��et�~n�,���I��
L�Uh\n�s̋�l]���A�"Z�0�� ��ÑI��$��I�BL��oN�,��6�T�6	��8�<c�K����<�|�X��1L�i��o�� �3���	�`��
`�$�)8�z�n�GG3{%:I*���K"n��Dad��Ii;���v�V�B�2C�C���l�H仦�@��'��J�)��3Vj�D�,b��p����x�|9���/�>^��yy�Ύr!������@��Cw;����^}�{D���z������/ye���������
6�����;:���p!޾����bX�j��ӯ�]Ä�[��1VGn3�pH��7"�wt��~/.49�xgz�Ϊ��ۼ�zg��L`��/��fy�A�B��H��o��*��^wzժ�[���SN��O/|7���o!���/.�t��������fP����z'�}�{u�%��E�w��΂����<�=�9���������t{�ɻ���O^F�ǹu���@d<aT#�ힹ;�ڶ�=�0����r�G6�{k�v����.\y�����\v>`�z�����7٭uZ�����N�����5�������vq��<&u����ݚ)G؀���n����a��דz�w����>��ٚ���yq�-�=S��ݶ��Ee��L�l=���S�V�R�f9g))}B��j;S�F��0D ���vf�� �)�,;�g?/4�~l ��.o$���=ؙ� '��W�������f+���b�����v�_{���|��W�w����[�tY�K���gk�/�N{8{.�pe'A'�>��~�����h�0���0협�z�5�xЅ��zO�<��<Xm6�D�G�[x�N�v��f�����]�#}\����P<m�6��Ǐ;|x��ǏK���{ۥs#έ���b]�nbwD���}��پ===���<x��Ǐ4�T�$�������t�%��_��̄d'uӜ�r�o���r;~w?K���褜�뾫�~���)�[lc=q�pu��-�!m�l���S-��S�����y��!���w���an"�β؅�[ŇT$�w���77}�p������[m� g��-�՗���p�盁��ȍ���"�.��/^W{�fg�$�Ͻ�|�y�BK��y�\��L\�ܹ�s�D�J����o��r�:!�&}v/:d"i&J�I	%K�.���O���J4�@�� �5����ODC�&��7�	������V/�Z��Zq|$(d���+kd�r��	���3�ա�]��.��w��,8ܛ�c�f����Bg���	8�0I���,K�P꺨�d�_}c�����[Z�8=�$�:�����e ���6p�jx��l�c.��HH�V�t,.��evN���ڻB�	v�%��I�.�%lٌ#�#OK�"�QpA'�V]�j���v���3k�ź���x�4����2!�L��Rg#T+�zdo�}4�A9�7WCgw��H��š�w�S� ��'�(�i��0�6?��w:\�p����|�������D �d�I5�y	>N�n7��S9���p�`�$(da��̳m���?A�|�����,�L���[gz���l�3[4㠴Ƴ,�F��A��V�)�ѥ����Źh�`��|NQ�yv{���t^�{l��.CPu{g��Ԛ�/�g+eu���J�H H���0�|W��1g����֕�w��ЗċO/�Y�6���U|~��=1#*��9����A���l�]�Wb�=q�9��g�$`f�Xk(�Ƙ8�5� ���m���رx�-�,�m�\1f�ur����J��[��R�!&�D?�jkF`]����>O,n��t�a�f���Zϒi>I�N
LW�<�3V�%�(ɏ�Ç�����[�͗¼Ks�p�F�B^����m�hd����e����@ �Yn��%&�}���Rh���O�*��<�
�š�s{i���98pQE�"6Wc �9n�Z�p�aS�4��9�Η�l��?��q��MO#���1x��'�7|b���.�o��D5��9��;l�$� ���!'Ra���w��s���8�����KN�1ˌ�2�����ۀ���I�������w͌�JVZہ���s��y��P3�����K�C�Dś����g�{��M�|�$�zV+Ƚ&���~��G��؉�G_ߢ�ņ��xA��Xt��S´�믊<~4�4� �UD��Ւ�$
�v�Y���H�mD<(ؔ��2���;9�M�p�{n
����{DKsncP-)I�Z�[0�e"J��	�˺��Х��X^��	�5R.�H$�Klk�Z�g絛{`� 0�F^%fA��\�dLh������3ku3L4�#1�#02�rełiq{(��9:�#�a��v��i�������6n6�;hc�3`�������uC30&�00��ղ��?[����ݺ������g��g���ޮ��7B��p�nC�v��UW3��V�;f��AI���L�`�"2O�1YӃAN��"�5<�b=����x�X�A�9��/K�b+�O��3�#D _����	�`�����8"��p�OM�8)���nķjls��f1��su�r� ݰp&�i!���74o"1��o�0����>)3�aU�Oo���8G������g�~�&�[�:|��p��	G�`����v�Ȼ��`�z���ȭr�|E�󻔳ak�x��3�73L�G��
L<�ԉ�/;pK�y������汆1e�1���k��Z�TRc5��tuk���z��B[�G������c����O>'ᙕ����a9{4��� �}�V!���1K�4��	�o_�Ɗ��2�guÚ;�ф���� >^^Z��j���v�\�y�m\�:�M{�����,^�Н� Ɨ�'��f���A��ק�`���0�eY.�M�	 B0�C3�<+���y��	���&p|���
��g>��UإX�1�`N� �z�4�wS-���[Gz+�8#i��t��N0߉�mdciA�Î�I��\��M��7�v񚭸L�YM÷En�l��X�sv�Zߜ9<����z��z�e�xB�I�/��'�"���is���e��������a�#��a����fm�h@$޾mv�&�Ι�&成��, {����ѳ���J�%����� �p�Q����>ux���3�3(�siw5тj�duf�J�g1�1��^��f�Lm�o�}���[,�񍞽2>!2!�v$�*�?�|���m�ǋƈ����YwY��&o8�S����?��T͑Ϊm�p9GK���Gr���WQ��ޗ�� �vr���)۝��z��`�@v��cG��R`�`��M$�n،��9CVp�����WM�6�e�aV@Ӵ�4���qN���ƈ�����f�}��Up�]fT���<�,6�"�I��� ��{�7�o7�����c���WlG%b���l��0pG&�'o8I�J\X�mi�v����gś]�\���
LF�J�A��X󜭸�f�Ȧ�H��
E㰀�8 �LS�������7�{�kC�?�mޗ������b�K�m�Ǎy��=��o?��t�ŧ�"4�!��Z;���U�.źW����-#��G75��v�M�Z�X����^0H7�ݳ�A�go�����XIb�c�:�ߵ���m�0�AN3��)8rp��gT�I�z��X�F㿈;�#5MfUp떬e�Y�ۈ&i������k�dT����ٔ�V0pA�pࢋ�@I���ي�M�L��FR�F�/�/��g��ڜ���ȇ)3��Q���k�h�Ȇ��Y&��]�T,~���ҕ��_/��ŏ&DH�j���1!�(ur�GN�ʄͲ!��;�ŕ���R�Y/3�GRsW:�p�}����9�y�1�z�+}u�+g/ɭ�g��li)���A
�ό;ʸN{e�{���7�BNؤ'�v�}1ްi�?%t���u�N'Ǭ�m��g �M�A���N��� ������X&G���B�)�	wj���"�JA�6��k1��.��7��ߜ��	=����>Iŀ�.ۛ���O#y�ޗ��v�]�����`3%�AI����I���o�e�k����m��w���֎�Ub�e��9���|G)�!&�l�-L;A%��Q>"����ۈ)p�)��h���Yj��3���9\y�Ajn��Ϯ�|}v�B)�����ٗ#rᆂ#9����`���۶���<��̬�K�/�C]q�����p�>���$����#�8g[�sz�Ob�[Y�F,����5V.�_8F��� ��O�Q�I���ƽ:�e����
*Mc��l�B��E͒���ay3f��i�Ř�ʱo��0�u�،�Y���c��ݮ�ݸ�è�p 	7+_�i�� �o�������j\�v��6��sWiX����l.�j[h��Й�D�,�eA����me��Qѱ4��bn�)��HցwV1m���Urڑ)!,*h9�8r����2 h�t�!Xh��u�Ը3�Uǲ�p�8�ZWR�Z��\�ڗs�q�[Kh�L�F�k,p�36��[���6#ƨ�%�2�e�Ț�}o^����sk���ZMs-�+jL�+cS][�S��t�S,��n�|'��v�������"N�)�#9'W��t��Ȋ�V��0��& �Ky�ҜdA��r)3�~af�0&��/G`s�n��Ѡ���|w�@�����5���Nw��8'���N/��s�Z�3��Tw��OG��pAm��"���%&J���`�5o�(����4��������'�(�	0raBj�[�����s��:�9'S��,��ͶK6�(�5����ۼA�g"�khv�k��߃�M\�~ok3�/cd�� �0t���o��]��ˉ�3��< c�p��lZ�To[fFw�ڼx.\�98rw�	��Wn�Ƹ�{���}#Ys��"d�FXG�nΖ��[KiP�K���KU��A�}���^'����~�H{L�x��d�;��>v���Hd,�s����pJK�;��;�H"-��L����p��6������ޘZ�)Q��̕4�&����!�'��O�����fy�����:��L�{Y)l;ÚՃ�0���9�3����p��|����|D���?��2W��G�k1�+��A�gdC��;Vl2�砺��3L����	\�Ȼ`࢏�aQ;y����.R�h�cf�_��l��8!'#�Ʃg_n���C�Y��y����wϙɶ:i����p`NS!���Kʋ~���X$�����[�����%_������{[��y�Md]�5r�৲�1�+U�	�g"�>I��ϋ�dtV��Ф�����^^)+����Y��	�8h��5�c�ݥ*�2S��c&����`W}�n�8�>�_ߌr�.kœ�p�ԃ2��K��;��8���L.���禲e��+��G�n�6�A�I���3��6�D���}�/�[8 ������9Dlu!��pc������ܜ8(��nk;��eC�#q���gK��Rp�$��tGu�<5�E���{F�=��/�*|���s90�e��Jۭg؀xq�����~e��(I�d8*���1�
u�&���=���"����f�y���k68Uv,|8������[#�k�M�T�|�\tuT�4�|A�i�> ��8��e��ӥ�m�@�;��IpC?�_������/|}��0ZW�4b�����X�X(޳�v����Ԇ:���p��� �Û6_��KDR�8a��Y1f�|=ϹR�fd��юy^2A��x��j���4�s/[���4Fk��>q���I��2!�Me�dp��|8����b���R����"�8�ϒg��0>7l�zf9�;5WOw�`ѳ��þ�2��j���~p�8p�C��p��q�Զ�3Ѭ�sR�s��E%&s�D]�n�&����*���1�.s�{)�����(��NN��q�Բ�'�F΂2�8#2�<m��E+���5�x�r땰=�@d���v���a��E7���sQ��t�^U�Q��b�F�&t�zѾ���E��vA��'V�E����w��N����ьjA���N��d!7�Y��QotYM�v\�kpҕ=#��C�W�98j�ĵ��=�]�پO��<p��8&8&D%�������x�?}yU���J䦤�	��B�4nc�4��3��H[���CgWZ���}~z�~�	�>��C�>d��&p�U{���c�z�����H��j����!���X�p��E�')�
(ǡ��2�;1n�Us"v�am�Q:Mvfdu�|9u�y^A�g �i!�M��ǃFZ�g|��>�`%'
(��I�㥙��T}����!e\�Y�پN��g�L8��Ȣ$��1��B�-���=���dǌ���r�&m����U�Ԇ=b��{����`��O9L/:럖ֽ7���s�˂��J��E �N��SA��Sm�5���-�̝�x�n땷�`��3�}�d87l��& ��uEs�oMކ���C"�,�M�SVz��{�P�����9�f'Q �s=����B�T�����Yh�4㍋��ۏ�n��N�W]}|W)㳟ik�3j����<5�L�j�.BN>k�6���	Ĵ�1�C����!�Ӓ{O�_)�j��<¾������.d�&����s�G?-�ď�2���V��u=_;�7{>y����R�����������v��y���;���b��u�`�}�;;�]�p���؝9 ���z��n������q&��{�o~~=��&w������Y�'n���{̭��Ju���^o���ǹ}��nFC��Q74�!����Ϋw���=��Ǽǔ�j����K��Oq��x����x��2v��ܸ$p���^#yxӃm�}�^`��q��%���0�;p�K9���p��|�^��=���[�q͓|��Ѯ��I���j�c�m��=����YOQ9��qij��Ԝ����j~��ͷ;�<�{��v���I��:�u��Q�7G��~����خv]�{r{:.�m�w�N����C˞]�=���ݥ�&�����|փ��L����k>�U�����������i�+����A��`����FOJ���7��������p�<n�91�U���{�Dm��D����ŜB��n�����xذP7G^�a;M6�����\x���q�n���h�0��a�P��G�x�Hήoe��8=����H��==P�t}��Z�}����=7�sa-����l{)Zr%��cc�����|"x��|�%Ԟ���I� ]f!]�o.����y�o�z�K����yi��!����,��7q�"Yf�t|]�Vv^�h�Q�4��ޞݼq�o�o���7��HO㓗��tE�I�s��b���^뻮����t�8��n�<x����t]7�ݽ1!cw5�C����%�����ק'�O�\ܮ˗:���;�/D�`����=���ˇ.��b���#;�X�/��ǜ�7wk��@7:Ns�����~{�4U�e��w�^n�$����#^����=���%�耴�)6�8�t�gu����eۭ�<}��i������+�"���&;�o���y��'Źi��S���wM$4/whЖ\���O7cdI�� ��9��������d65��|p/w);��/��ej��I�������L�	����׺�������{��6o�;��/'6nHYX���@5�y�a�X0�l�\\�0���$��Y�L7Bց���h���.��T͸#���$�鶫��	��`�5�V�!
�������-��	���(���v��Ȱ��m�l���tumf�����m�Z9����ᆶQ�c1����+j�f�-�֫e4��d�Xa)�a�06��1�6[n���5K����jv�+l�K�`�ZՀ�;8I�R���˕��p���\P�cT
b���J�30+���L[����Qe̚e3r� ]u�B�-!a�T
��*ږ��V�ޥv��l�%��1��  S:;j茥&���R1���E�k&e�����V,GlaCk�b�3BU�cRX:�id��l���d�<7��/Y@��r5-��JR`��@�.5�20:��0���`if!e)�sm�*��sVbc��7,MF(ͷ"Cj�-Lf\*8�R]t`R-���!ҡ�K�,f.r��tv��9��mT�Q8���k����H�Hko��)Z\GK��ݝyu�n�k�A6��֪h<�1�مu5c��i��li�!���jMj�9lFVm��[Dljb�-cM��]1LY�v�u�7$tܫ[�)Lk�4W�k�e�--�r�R�[V��Ѡ,�X�q�-M�`�J�)1���]��гTB���R��e�$�Na]����K��X�jM2�R�̲̬ ����<ʹ2Pe�A���kKU�1�Z\3X��lWm�Z𛪘�3e\(Yu��Xٱ�0�pՍ�s�]ˬ�H	Ĩ�Hk���ã%�[�-��ƳH����h:P�cc�6�!�5���L��n��9�#���f�Z�v����9�\��Df�%e�К�뉈�R����6bb4�W������pevh��`1�j�sn�:��,���K�5t�x��in��kp`�'����ax�΋���M(?��jM����B��1R���j�9�	��Y��X��S���	HCF��l1C�LH@3Fg#�nR!�2�\XZ�3#���fɥ(J�-&X��Sb0�*Y��B^U�JF!���q���݇#LZ���P�j�rsl�b��ո��݊q�U�� �ZQ��	�����՚�`�B�Fl�k��5���~�_�ߺ��Q�xf�õ�aa�������pHkq�z܎��Fjn[�8�9N���BN���b/��%�7��8�5��p���1���O��N�����&�|�z��t�F���Dcw4|V�T���>U�$q�/C�0 �0px���FMl�"�U��3�����!92\!�Yd�oz-��p�|ax ssPo�o�ݻ,Ne㢲�[qN��aV��A�S9ʾnBY'4P�P7:�b�R��j�V��Ã�K�
N��sb#�$�񳼝�8���|z���;.2*��#)�Ǐ��$�AL�pRgif��\M�U"����r�v^��91����`A��?�8pQE�I�םo������UZ;F��E��b`Ջ�k�6F©ZSd����I�it�c]�O{�e<h�_8pBN|C[Y6�cv��٘謮�n?n�j��|xoRm!��g ��&�*|���j9��FK�8�gP�R�A���Y��1;=�A��jM]����w�.�s�M��`T�WR������fos��s3���4�B!"Hז|p�pB��U}����4����x�6x��Â)DJ���;sCVyi � ǜ�@�b��B(�&�)2J�e��Cݮ����Le�c�?��058sE$��I��U
G���.l�)8z�<�>L�{�Nۇ3�v^8K+�� ����uE�ؑ���cy��;��M� ��9I��Ṕ�(?�\8�[���Z���M�LÁ�`��5♼�?�ݓs÷q��|�/�>S��c�Ie��Z2�4�)Wj6:��:U�p&��r��!�|o�<��q/�a�n��ݳ�U]���+�&2���������Фp�²1��W?�0�BN���EC:lje��08"�����#�4-���V�WU�3.�@L�r�n9�a��,`;L�lX�^�W��(���]��z{=�}u?�&h�Q'B�����wu>���O/������}���8=�玨ů�����-,��	l�%C��PD�c"#�O���o�$����i�HҾ��L������$����2M��"�۽���V�4���>�֙��g��Z�l؅}!d�g;�	��^�N!�b���p����pG�(��)8�Y�픻y�ϭd<R	�u�p�p�W,n �2�A�!!�f	�����I�ws�Ʋ�N� .m�������ʒ�Kj�î���6��֚A�Ÿ7�X?�#1ÔQpAI��V��s3�ꢻ%�ɹ�]�����zD�r�A�B��D9I��Rgm>�O�&����j�b�=�ѷ��ۡ7c,����s�q����|��͛9Ɔ�xk���3!Q`�N ��?���ȍ�i�,�y�)�i
m�f2*��y^�E��r�מV��U�4d�4$o�c�l�筹��B�x���<�n_A��%�ɻ�	�gа�x��� �7��� ��R0E�Zm*B����p3���vۧ���1�vK��2�\��<c�m�3,p��&�I'�c�Ja$��=���-��[7��B�y�"���$�eC�b�g��]��	�d�_:Fx��8�e>�(�n�uj�1}�a� �y�Ò!��6��,A�d��I��&�3rJ����4c487h�6�~�=|�4p��w)���DuZm'o��i��Xގ8SV���vli>Z��o]�����F�V���D͙�՞⌐w��r�ᖃ*�I�%�ɹ�<Qr90pJ��VD��b�K����ȇ����Gi���
"���	2�R�F�����e���	��g/�#�����9E�0o$�Ȅ�8�9���>Ԍ{'J�Z1Ñz��BdC�7i�`��n���Y\��3,����h������"��`/��!C��9	0Qm3R���`�%8}����LU*�����n'�J.A.���L��y�˻����L�2�y��#���-��LP��}�Iʘ����;��)���[�̲S&�Pp�i�*R>�����Lu\%��G���ߙLѢ7f���E4�@�"ɯ9��*��]��R��++WFc0%.&Ό���l�T���72�.��%��H����n�2mDM0"�`�Ѷ��Y�u�[��뱍[R����R�f-p��gPn5����]����l�����*�yI`
%ҖZCm�l���6$ձ5���\a��Sm�)�\���h\:�im��l[�*�DXir��y�M6[5Ϸ�_?��5�:�l]b���B󥚚
f��`[	nd!aH��骃*o'����[�K�3�4��v�%&p�s;�曘��0��5�<�f�
�t�����0�Jd_���Swwh^#1������3MfGƜ����	�g"�pRh�L�C�:�{���`N���Ϙ$�F�'�n���m��gyP�zU��{�#��>jp��`�>���T\�Jsc�h7T5�}mG׭$���fwʋ=7/�	�3��!u`��fm0�7�� (���^.�<M��͗�	0rS����]]/��n!����}�xӓ=X����o8L�pRg�4��\��B/ �9f���`Y����!��1���J4��`1�zܛVn#���%��Ɂ��/��p�U{�0rzU�͒������p�.�j� �=y<Fb_��Y��6����𴡉v�캞�����3�;��[�b~�=�]sM��fm۶'<͛��CT[m�{g����d��|�`v���11���Ϲ�,[�<�||}�I�7�ԙ���w��;�m�;�0 �0r'QFzg�z��<sZ=}h�#O���G���w�醏&D7t:Vrk�P�z�pN�h�iɞ�n ���D8)3�)3�N���D0��zuP��#ۮ�Θ]�ꬽ�c�R��l��&a��#��S.w��w��C��8 ���&D?�MX��0�vF��gu7׃�cb�E�b��x0&郀A�8(���e�m��.xϿ}[4�e�E�Zk�Mq���#U�X�Ь�a��f�]��C�3GI���x�pE�+ħo?�DD,��}�/2f�����1��o����%�c?� ��y�*�����&:纜\=�+R�}9T��G";����.A�u��!��.�#/="ۈqn����pA�C���~!F��?�R+��Pg�$���]Cx�f���϶�m �j��u~p�� ?����ʘ'��e���y'�]��>�:��u>T,��r���}@w����|:��Lʁ��'C�0&郂���E����|`��׹�L�A�]B��h����������3;�/2'�� ��^���J�dV9�l�p3��3�f�7��=y�'p�\/u{6Nb�z8p�p����йU�8��������[��zBdB��|=gX9$+E �xAr���Q��̥�%m0�T�
%�Z�ٵ]���G��42�����C�:�)���2M��R�j���P7��d�c��\d��Qz�����(��p���?�E�������XDF�x�:D��d왝���Ս���5o�l��e�W���]��ҩ���,�`|b�޻o"��I�ʝ{f���B���]��c>w��?��-��]�k>I���r#sN��GE�:t�����wYwm�0�s���w����E�&������E<Lғr�K�%�4C��[.�����q���9cL�����f���n��R�X�ɬ��ͅ�/4y拪4���j�g��d'�,�����L�5��:��Q���ÜS>��ǈ�Uד�bwx^4>OV7 A3L�"�r�8 ��G�$Sִ��NMw�~$ٕ�
��n����Pkb�BU��E�U�]��I3čΰ$	��`ࢋ�Rq<ks��q����|�kpqa�E,=[7U�9�F���H���3��o�0J��_5IZ}'���	�g|��y��w;*���x0&郐u8Q�s�iX*�����pA���	0��y�"!0���-����e_Ƈ����&i��dC����"��d���>:V���>��Zp���l$]^��
.���7���l�pB����:э�0���E�ݵ�M�9W����Ü��S\c��u\�7iґ��'�����S	\���V9��<-QG:N�_��D��۝�xi��Q �vwo��]��>�=k�g�-��t�<���#o�=�9S�:�(��3sι�I�܅�uuQ�*W��H��#S���ߒ��eG0s��+���ȴf�
`s��`XLJGhF��l���;@a�kJ�&u��)�.]S�H@3(�ZEC8mE�����$ۉ�E.�h��eմ���X���#ڵ�i)��VF\f%�VX�Z�le�1J�ѡ�mwi�!�Ljh��j&���a��܎��gs��f�M\���k�6�ѹ=!��}��h����1k`Tyگ$p��4�	nm08��e��5LD����t�7\?�I���F|c͗ۛF�wx^4>OV����=��/n-�k�h�7l��7�R$�ȋ"g��)�ښ�&_�(�#5��W�������l���;x��%����^%rv$�f���C�y��n�3�}mg�m �
M��6�;<U_��Q&ꄧ;����y�郐u8r�.!'H��/;�P�_���W���4b���vp����x��5�Z� L����Eﹶ�Gt�e7��pB)�oR`'BL��H���{�-p�V�o?G"�}V��~�,�o8n��Raq��������za��¥u��v�Rd��\�F�jV�rC���Z����J���w����/_��^�x��8{H��z]hs:W=��pt\�� ��g� �6�8#q�n�|QP&s>'�yO�:����UR����DW���,���E�V��=��
�w���{|�I]��;މ��Zzb�6�j��M��}�Ʃ��A�	�>��a���8��{4=T��g(��oq�`a ��0��y��z�X�&AI�<y�F|B�b�S�T����X���]�[dw��fK����I��2>I��!�a{�����|B(���y�훭ٯK�g�s���`M�^ws\���n�lx�pA�|C$_,��2J���E=9��j�w��3Ս��j[Ι$��A)o�:����	pIg�e��of$F�60Ё�U՛D�[kJ�1�Fҵ]9[��D�: �0�� 濑FA	0y�sy�)��+l���8�P�8L�eǡ��.�9�M�GԚA��`��\׎"(,��D�t� m�ƀ��~WhsM��t� Ͱr50pQGZ#����7_�`w�^C��%�7n�$���@�i��EH��􇘕>jtA�h �J��z&���.Ls=���D��!���G�>�<�y��&�{���`oؙ�NU�j@ūh6L�S1-٤FP�
~���Ä{�np��/D�^=���{�E���|�� ���r�x�-�ؽ��w���:s�ڜ������@�OwnD��!r�{w��}t�g�����{ڸC�Л�'��=�;��Ľ��K�j����߯�!�T�i�����6�Q'��n��;�e�-ª����ĿrW�{|��9^��	v�$�P|;s��`���ۇ �6R���4������]��b~�����g�b�f{xa-*/3G�F�*��%��٣�ܞ�ɾ*��O�x
�eu�=fX
��2<���κ�W�c[���rK(��|��}�cW���jznyb�d�9�zH
겞�/f���-�!��>�!}3֏gF�����-�s���;<C8vhUX�>^��צ�9�b��}��xn:�i���|"�;&��o1����Tq9�5 �h�@yNy���'��Ҿ
sǞ�$ߊ3|�'^���y������^�Bn5���B��E�s�r�x)Ƿ=�ou;���wo��n #��2C0�p��[ܞ��${~_R�>k���
��3:�;�S���,�IZ�4 ���>U	�l7=��\3%��7�잾�(��n�bҺD��w�]c=O��KU�*G�mĜp���f͗.�><�l��}U�l5���CkUe�x�Gq^dB��d��tp��9P���^ϖ���'���������� �;���D���E��~��&�LE|\ѹ���l�I	$�J��a	�4�ק���Ǐ�<x��� ��@� 0�Y'u߼��Fe)��*D$��I@��M�i���q��n�<x✄� �-���*(�[���5q�a"(�[��н�t�����LI�ͮFM����'���4��r7��rC �u;�ls�Ʈm�{��>q��\�2s�Iύ����h�Q�7;��#W�������M���漯.jJ-���nRZ�c����Q>��4h�l�W�y��Z��nXž�{�Esn\掻����yQbHlb�+�4cm�|k���U�E�C�\���A+���m�H���j
1?N�I��%%b�o��f�Ky�<�Am���5S��p�)�M��&e���)7����H1�pϘ������a�/0j��o;������v�6�땶G{]��n!M��cn�����V�w;y�a��SP ��8)6C��\��ֳV�v�+�5������z-�V�8�p���r
N�?>z����~�lv��f$f	M�����8h�2�&��V��bc[\߾u�zI��Y��<J`a>�Y�t�N�v���m��5�Sεt�β�	�U�����Gֳ@X�Lol��M3��V�j���ΊTg�[�h����rc��$c@܆�WB��c̩��s9ݰr�?�%&�=l�[�0�aO>Q�购�wp��Í[ �mÂg ���	?�V�,�YX�k�3x��D[�� ����W�j+v{xS؛��[۷����k?��q���z�9�i�W��{�έ��c�]�2H�U3�݈tӢ��L���0塱e@Y�v��3�_�]��Z����w��_�쳟-g>J�<��p�������{�t��P����swgT�3֭�;������pA9n� ����'F\G�K<��|����Qٷ=���а��g%1,+f5yvE��p���Ō���~p�0v���x���,���?�e#��5քuݨ�6�\k���<4��_��K?�z���U�1��X0dL�V�h3�c�?uh��%c�W�ͯU�<0�T���Ae���&�s�BNv��m6��<����'�(� �'a6���NkS�n�F���#���8><d��Ð��?�D�|Ag��p���  �"ݳ�JL��R;�3S���v����m�0D8��,�r�(�^0�^`��QE�I����Z�����l���{s��޷n�a���M� ��r2!�Rg �Rl���ֈi���{��{<�l /��n���	��a�k꿷BȎ�j2�G�_�|m r��LK��"7VV�r\�f�3߹ﴖ�F� 1u&F�'�=wn�v��b*4�����>����q#���͡��kF�����p^�ՊP&����M�.s�U���"8e�0�.�,`�b�6��c�W�m����lX-݋im�vh��궅���e2�V�a����'j)0&�JV�����õv����P��v%�3�,Ch30pb�ˍu[�f�H�����S2ʸgd`8���#5�ؠ0nYj�'��|�4��Q�a��U"�^�R�ط[%SFlZ*�k"W|����F�`�qÔd�&���u!X��Lw�9���wL����@\��E'"�~�]�M�9�z0%�m��eW5u�Z��zb��_n�F�:G(��v�nr��e�ws�ue��L�"p�pBLR�Ȏ��w�:��Q����bj{Sq�zdC��?��o"��'�e�13��.XIiÎ�dp�]�[�|��R��d��<Ƌ���Q �D�X�6\?����&&D��n��_)�U_x����G;z^��_��G;�/��`����e�E����?{i?��ܨR�Ä�q0AmYb-]�͹4&���� �V4e�qe���~�ۋG��>�r!8ȉ�c8�Ve�{"jwi�	�`�lk_�>���֐A&�*X
L�gc� �*b^"M>����	�Y����R�鏏��g�H��;���-:�W�g���_!$�B/U4�1��{���C�U�����$�IJc����R,�� B�����?<p��������ɞ��8 ����� ��x���*�<�B�h ����mg���ݲ��O�Ce@zj���VQ��V��c����ڜ8(���/T����ΆF�VͶPo;�`e:�MUy�}mdO^ӭ�.{�S���3,��pf��n�i��� ��E ���)8r�-�A�v�>wg͞�+��.g����d�bp�tX���^�>��[{�x���FU��Y�&��Wkv��0�نm׷����8[T�1ٽf�F6�����ݴz�u�ҝ�;���ry��� A������y��Q��X�pF�-_B�:l@![y���?�U��wv�;�USӭ� ��p�`ɑRn�$�:�l//4&pD�q��r�%F�@I�U7РKa�Ǥ�ߴ�O���`m�WG�} n?`پ�oga�%�߸��9Ox�zs{�\�z9�Lݯk%�M����w�r!1�90���>>>�ح7�r��+̺���y���N�$��@L�pRg\\S���bnp�a6�汜AI�ԏk��뎦�J�1��oe0r.�hnࣅ���&O�U�~����/>`������mFo=����q�ݗo�
����`*[�;���C�v�A7l6�gmP�����kAg�����˹r3gdԡ����b�����s�˂a]X����ǿν�����`�\�q���ޞ����Z����I�S���+\ُk\8#y�"����n�ȯGI��̓�܏�Z��6<�;ѫ����ҭt�q��a��(�[&ˑ��Ɲ�p�+��,�.An�N�2"�D8�� �Wg����>5-�DII�JM�QNׅq���¼|�p�:\�p�Uص�=c���Z���8 �� u�}���� �4�Pv%��D����4�8f9Kt��c[G��[�J۞v�7��N'�3�{t 񇓪��@����?g�jI�C3L���x���Ds��6�y�L� ��$�o�ToUݽ`^4�w���s^��U�����L��N�\����7.�z�vY��IQ��?�f1*iF��32��Rh8��5�IX���j9����f���w��ҧ� �������!���	����̥+ܵ��������9��vܷ�A7l�|��C�v�FNe��N�Ӷ/F���8q��]�uX�y�����p�r10	8n7:�\��>����C�-�	�g���
g!�1�Ʃ�n�f�>�J�j�U�qTr�.w���H �p�\��p#�]��鉽��Ŋ���mG��Dˎ��ȣ^1Ys�&�6�3jz����R�vUMo�sx}V�A��<��R�8I��Q<n��*�T��2��oU�{W�Y���<9n����!���#�����	�[����}���b�k�B¤����1��x��x����CcL2j������{�!�^���g��_���� �w�;�~3�z/�q��/)�Qҫr܌L:�B;m\b���L͉f�� �[�<�+��\���i�2p��bJ��sk���0L�cJ���c�\�������1�5�ɬ�]�#�"������e�0]wvAꠥΚ�6�uPu����f��#��;Z1��6d&�BT�[��aXŅ��[SJ�u�!P�3��|�.}[�4�}����$˴�U�.�1*r�M�	�M36����&b�X�i�����_�7���7l��n���Ž[=�*�\%��	�8���L�r�����4s\9�e��������'�AAK��f^�d7��y�g�E�m�1p���3z���dCx��fH�촺j���w��4���ۇ|�$�q���o#��r�Ռy�ˬ}���%�#-�y��&�D9����=���̶7歫�ɚf��쭞�G.��x0 �0�V8�k:�J>���	:\�v��n��Qko�c	fD![R��T��;��m���N���ow��p�ٲ �]�R���b����<����Ѭ��$q�CV�h�ٶ�e%ClnE���F��p��~`��f���qט3{:�؋̺��mpp}ٮ.ݮ!�0�uOY��[�<uW���/�v�]��^3fdBj�*�
���as�ز"�3&�ʇ��[Ƣ^��>��fdc�Ni�A)���=Q��_������O��o�l�p��mS���|| �$p5��k<�����0�e�\���57x��d��2TcXʷ)��h��L�`�޳d`�z�eݙ����H˘��op*��2!�R�JL��S���Ж�z����a ��s�Ϝ�?�+=���?E�������̗F�gS4��^���р��m!�Ri ������+)�[�o�@;)�����&��V�;�`A�`�N<ȣ �ɫ�<&�?�g`��&�	L�(6�k
k]��MH9��a�ғfd��BSG�U��'���.A���&�(��j��k�#.b�u��R�M�Ŕ�p�G�&���pBL�JLL���e\͈vc8,���8���6��腗t����t��u��@aw
��A�#<ɼ�y���ro8&�Cy;UC7=Ќ?�'ɥ��/����uK��ث|پ'�����'e�����ܫ�y��{��Hi��
���͊�e���x���g� ���	@�GF*~��#����*�8#S&>	8pBN�voW;����1��,���)w����+1�]6-�Nd���{��r�j���"ځ�3��$���IÂ�wջ��]��U��oWp��Z9�������8�� @f7�]���oc�CL�FQ����.����8�ə�i�3Q�#����8����&-u`4���w쿾��Ǜ�����y�{5�GX�VҸo@�5�$K�XU��9u�'5���?��w��Ȭ��������M���?����cse=f�'1��u��7m���	�x���2#�����h�w0ۇ&�p�f�I�nO�|�g$�z{j��,V/;�\V�8�p��I��&pA�H�O��Kr���sv�A�I���u��B�eVҴk7x�U0��{�&b���B%��u8��^D<����m���r�t����^\eT���Z�|�^��~6�!K�3���?=�]��N1�oM���=��֌�[�Prۇ$)a��f:ٖ���^�����6cB���A�)7�oH&p|�^�[���*��l�����������IZb���m�,]\\Ӊ�&���˴#W-ͱ�����^0�� ����Ǟ�������냄%��V�:�H�o$�kV�9�x�x��u�g���M���+N���r�eV�Z�A���#S�&���~ȶ��Ek�!K�o����p�]����5֨�a�P������1���lƄ���L��9I��&g�]��rΰ@��N�0p�j�|Ǽ�P��Ѽ�]6x��`:.�������3b�_z�x0)�>�Pț�
M=�+kDB�"�ϊ��v�5u󪶊�u�����#S�4�9'��yՠ1��q/O!����P$�s�'}t{��!����~a��uN�ýr[i���K
ۛ��[�6�^̾kW������������k^��+�O��[�]�_s=�^p�q�4��Ƀ�Om��Aޯ�S�|9����<k��.��N��O�Ms�5�5ҔG�>k��J��Ν�!8fޜwOlˠ�Ĝ�p��> ��x%�)��*u���d�������9���h�q|��V�\���{}X<�=A��)��˿OM����a�[����'A��%�u~9�gk�\M�vI���O;/��	Fqu��ݐ�x���`�}�Y 쏮?w}����b}����l��Fw���}��Yg�y���I�6O�*�UX��^^B3w
	E��' ��tz�_\Yr�Gsfܵ�`}�&���w�ū��u����{gu�<g��׷�{ף��Ǽm��c��������D���G3�8�A�J�=79W�ޛ���.�H} ���F�x	�!����f�~U��{��Ø���8��3��Z�ś�L����X=E}���=����<�xf萃����U��n�w�-�p>[���s��b�6T��T�A7��������yǷ��ΏO�K;4�H[q��s��#Í���3�+��'���{w\������}���(C,�,K�U �oy) I���}w�ǝq�{wFI������r�����.���q{�IMIx��|�8f#�NÌKZ��t��p��6���2iY�v���� ��$B�cy��>�������=����� k��<D���Z{K�k��y�G�1�o�Gz��>~��pI�K�
�Ѥ�F�F�6��BZ�;���4ۧv��x��׏9ȒN�w�ō�nEbH�f4��㲍��HI$�t��n�qǏ;|x�o���_�F��fQ@��4?�O�ۡ��n�{��V�}m�0�X�AbLb�XM�9���L�TQ5�%�n[���TkwQ�������	b��l=ۚ��m�s� \�6�6$(�QDZ �cmy[����&4\��$�	��(����b��F��7��1�
e��ܠ��ۻI���b�Y�\�EEd���4��W2��%{�#h�DQ����X�ưlE��F�QPY(�弼�����0IlEI��i�h�XИ��l�eb��:�,s�kԉ���e�u]α$k��#.n#�.����6��-p�h�J,�3Z^h����YJ̄�v�qc"�����:Z���2k՘H�.�v�sEl�`K��9�r�YU�l�J3iX&��R�������2��@����h�`�[Rj�ܘ�!��^�bp�xX�TW-`L�e3[����&��]ec�ICP�e֍�M�pi�����L�h�4����q�%�YnUL0��Ybb�g�[Xiv�$�PHR�ZVm�����T�Eģ��kVVm�P�T�����M���XQ)[�1(�l�Ҹ!l$M,1fq����5�z��]	�Z`2�Ŭ��{c[�j�,�g��L�nM.���XST�ژa
�62n���Q�v�kv@�˰؍a�����lb]M��E��\��v�
�L@b��6 �W9�LK�0� ���m6�L�7E�V+�)+�@;0�+Y�c���vBix��m)06K���u�]��`���	��a� h�1�(8��a2��P��+e�� ����х�k��@�e˻,a�%�k�h�HZ��Ц́P.%�ͣ"�X����qX�h�c7IJj�����66��ˊ����j4�Deڢ�	����6���U�Z�!�4Y�ˮL�����de�º�-�ו�j� .%7Mj49�A�,���ZP٠uRT&�2��iHVLl��1[ q1�XP��3^�`қ�Z�k�kE�3E�=e�X���ܡ�s�-�Z��*vH�Z�RSf&�n�����@X�k5�4#R�6�Z�TC"����5Ι�®	u�΀�{m�ǌ�v�
�2��Ԗ��Mu�z�7`��f�j���ƨb�lU�Q��[\:\T1�Mn{mB-����M��-ŊH��͔,�r��;,�t/^�+6���M(͐�Æ�+����31�:��5���`���d�zO?|��!�����h��4)�1��;��e�q�=uĺ55��bvv��*(�͍G,јt 4jC:]45P���`�"�cDm�M���5 ��n@ηSJ���7iD,nm�Ʈod`�]�jc34e��#���f�h���mc֥��hŬ6�P4u���..n�eƖ����`����`�˥�k6�P���n��\7���
��c^-�ҫպ��\�x����i��j�W]r��@�>xO�g��嘇}�p�����0�>��i3q[���h]��j�y�c���6h �T���i���|BM@������NP�b�9�r�{ˋ�U�'��b�?�0rZ���n��.�����ʞ�.8�4��������?�&�L��;�1�WW=5+mUl���p"<e0�6[�0�|�� ��ka�L^��㠃�N�������{tK\N�y�e7JL�]Ǫn]�d�H�lg��d�� g���(�Nci�A�v�S�5ֱ��ӽn��7���$���L8L�ׯ!;y&��Xl5͊�ʞS�djB�p��(CK(�nq�Nj�u5��(�v�]F�Z*�!��f�A��	��80��%&��pw���sڪ�ᤝ��x"���KC��ec ���k	!&�p��R`��B�~#%`�SPVOZi��q���Ʃ{�m��t4�ş`fUB�ڍM �ӿR�O�k�ï�r��F�k}[�æ�u�����{���!YQ��[���5on�k���1�vSw�%&���dK�]�R�-����pA ְr�"��	,�dY��m�12��������YI�;ظ8%&5�����y�Rg|�l�Ě�3u�P¼W��  �	�V�v�$��)���u��e0pX�
���[�]���|������)���P92�
�;���Uݢm�{�Ñ}���I��$�$�%&\��[��~��'����O���vi�LJ��2�nX7kb���uKRرDmdJ��:�}��>|;נI������uy����J3;ظ2��h�&M��$�H�`�#u����r�y�RoeTq���fp=���x�X�w�ٴؐl�^-����y��8 �p���J�Fݒ��t�lg�`�ݰrI��	K���ǔ9�`�L�6W��H7_+����d��_5g]SǤ�,��L�V5�q+Pi^��N��L�-F�����S1�vV4[=���������{��1z4������7�'�����A�I��`Z�H#�Y��s�m�4�����!'���#_:i�*f�y�7�&��rح۸�0E�8�w�<���O���g�	o8&��ږ��,ó�c��Qԋo\؈��mn��� �N���$�/F&�nk��P��t�O���ͽ����!�c섘6jŕ�*���̵�@x`^ �ϸM�pA�`�v0	O��Rq>04vei�}������w�f����zP�|������Rg>I����>)0r23���;�(�3�k��*�S���)�Vg{)0y���9}�e�����8�$��i>�c�������Ϯ�/k![�d�
�Fz�ݥeSb/x���f��Ra �����>'���*p�z�f=/���a�����G;����#Gn�X��q}8�A����2�yZ�d�j���R�^��F��*�b��=�gƨk|����)Q_�YvA�[��}��[��1���q-�L�J���T�{����� n�� ճ������$�JL!��emX��{��F����鞮+3���8 ���A�=���?��\ЉFN@��}���P�ґ�:�J�����77%��J�a`�Jkz��L�R���ya���3��Z�$�|�8��k�m\�JlEp�n#&4�]0����A�k�5�������M�0x��RV�:�?oxψlp�#u���`�v��!��_N7x��y�'�^�֭=�y���[8yM��`��R`��n�
���)�M�������es�&����	8��Dv����U�SV���������o�����J0J���3$��F��*���TF_��P �8	HpAI��
N�,]:�	v�8R�t6�B�3=�M����A �>g$�pRg ��i�[4ɼU���1m��s+S�M��{�I����ӽ�λrb����3K�.��HW�qWWQ��SeRO1��n������zX�AA�x� ����qĝ_'��f���C�!m�j�Qs�����^35�)9�8!���6hXg΀T	pd1K�Fz��@�qnHa�+�j���<+v�s3��[��cd
n6�1�`B5ZQ�����+��bfi���!+��Q�HA�j�tZY@�.�a�B^n�Ǚ�p�T*ba�̂�\`��	MPQ��0%.\��J( ��-�/����}����)��Q�j���, �C0�h�%�A�d���.�Y��>��~]RY��.ot�v[u������j.+3��!�J��,�Â3�m� ��!����*��'�c�QXw}��3�N�;�]��Ou�cݾ	T81��
Li8QwLZ8�A�xu{��h��Yɒ�G�ۦo}��m$R�0H��7|Uz*o��k��i��6l� ݳ���<�E{x�b�2�a����;���M���>ш���d���>�푁O�Lǯ<7�G;��dC��ݴ��r����f��R_d��|\�g�,�~���f˶�K�;�oM0r���(�$��h��5���?��C�Ƙ�/ɫ���.�S..�fY��m�K��8��LCD1.�6HO 0 ����]�ȇ�w9�4ToI�/���.=���o�V�#Y�m��&�*X��0X��v|�λdB�|��e���3n�Qչ�t�^2n�T��!<�Y�;��:��p2��Og�I�y� �.��[�e���`3ʦzL�,����or�j��{���ba��g=�]���0#�vy!x峂9��Q�k�s붬Ƽ͈�zy�<�U�1�7��1�8L�L�\�$�7`2]�
ͬx�8q,-7��'���)���k���[�Jh+�a}��9��SAV���	7`M� ݸr�2/#���a�v���U=�Z.�;�y�񢋃>-X�BoO�"вCUt�仝�����[�k։S8`[����)0�iNK���q�ڛ C��h �:�A���A�L��v��]���1��/����b��%�ن�%0pQ���:���(���/J�:�LX�'[�M�=��t��!5�t�p �)��I���,��T�Xs���)��U�BO�H7�޻q>��j�����@�n��É�G6^�{�n;��]���ߢ�����p��(&�Ty\��^��nn{�57�8�#�����H'Ȱ�p�z�V�ȸZ6\�o��pM&F&)��0	?�T�htª��������eǜܷ���Ͻi�6�;��.���U0�b+���fO��YE�L�{��M���r��{�S�wkx�H���?�F�\���D+{�X�9�m�87l��3��9��>K/����*~���g.�Ҍ���������J)�0+�P�dJ�}�=x|�y>�^���bn�8���'��dlm��js;�y�T[<��^�c�ޜ�2Ϩ?��9I�t+�����􇉫Y�\J0N+��k���P��1�5,�Q���ADW_#�'���Z����5������.X���������;la8	7��?�f�:����}��#-0��ڶ�L�9�E���X>������&�6��0^p��`�8q;]�$>�s�3;�x=x���`�oAŐ�0p��uT�=MT��y �����w?.������nh�w���g\�\Y;�� �uY��){;�j�		(�Y�w��g�'�$��sʽM]ˮX�u��	�Q�wM��m�̙�JL���'̓V��eE��� q3�U���V�	
������U0pA�9I��BNuRT3a�hN�foŢ�ω�fF�͵��5��)��y�K��˰'���7�#=��|���A�p�������*���ս6���u[q�GcwW,d�A���sH ��x��A�&Z�V�<�E��y��@�0r�8q;�VH|�n�hQ��S��4�8 �N��JE���go[����ٛ�4ѽ��&��a&�\]Z3x���w'�����~|~ �L�eo�A�p��
p�#��t1�d���nl����8-Nopjޛel�W�X��3�B��\���+o�Rg���r���i�0e�	������n�me������v���<��Lq8	H$�ˆއ��]����ӆ���;��L��q�/�x���؇��$�D��d��4��E<��#���_��go-�������с q��%��}|��wԾA1��`\r�@*$�^���\R�dA4�0صIf�u��CA3�ڹ.�F�iJ�zԥMa��ͨLKM��`�t���0���	��5r���k�A[3��]���+*�9z������,�\@{ε���u.��*(8t�774�R&]v��V�22��d��ƤR��m�)� ��k�u��Cfߞa��A��:ܫ�+qbCH�
�с5��@G�[M���CC9fč|n>�o?���&p>&o?�qc�V�		����p`��]3����f����Q��8q>`�8>0Qւ�ދ���"y���q���n��e[=�N0}4�A�����3y{������9m�t=l�u���X���6����#���ƌ�������pAFː}���I���M ��=ڍV��d CIk[�
L�z��VΎF������sZ`;W��\i��i����Oyda���;��p��I<��Sk�A�$M���ѷȫk����A�1���Y
L������?>�_������]��k�����i���6Q��%��m`�&�4���/�p�K��F_8�.)8p&�s�w����;�y�+�Q���sǜѯ�WK�"����Bx�ju�z�4~uq���㋈��)եo�y�U�G�Xr���E�q���{}#��M�̜i�)j��e��)ML������W5��J}c&��7���'yY�s��w���P��~փ����pQFgo���6��[��8!s�G��'�`������,��Z��n݋��E[\_N7x���}V�pRo?�L��m ����Vj���[��F8�������6ۻ��K�u�.��["0��.�{zpW��댏g7��3��n�ρI�I��s��fD�'e�wb��[��
c3�cp>T�� ����\����[г�ߺ����ueŁ����8�?$�2M��i��	�Bb�)2�� Kǁ2����|���_1����̐�B�l�wF�t�X�sӍ�*�9n6�ڣy�렇��[;��&�V��g%�&탃5�!6n�m��F�Fs��GY����ȹ|��z�`X��#!-���i�(g�ȟ�@�k?�x��������U�3�ZE�uE{ �
�pe��^�L��*�7���ó���Kw���n�j��= �NI�Q~y���N��ݸF�����co���z��_l>O����Z����S�z���7V��O ��n���(!����\��|�ƭ�f]ѨO ������Q����G�v>���6��w��Of��9�����{����ƿOp�f���{�{����Q7<]#����� �ӽ2U+���{����+.���xp[a��"M�ͼS��v�=����w�e�8|�����HF��FJ_OY�p'/
;���v��Cc����O�ņ�~�^�{���wG�;J#(�=���&��;�%N�1�s�o}/��%�O�1ben�����E���>%���+�n�^�O[��Ta�Ĵ��V,�X�75띩#������<���;�ܙ�OQ��Ӂ��v�~��n��N�{t>�L�����y�x�N/��ǱÁ=���gw�QLG�7����;��_w��s��ڰ�o����O|T�c9#�-ɥ�%ӷ՞t��B˽��p��b�S*8�z:��j��~�A~W�0P���X}C���x�T;0�9$��&g*��Ŕ���,���~����tOlL��b��0���=�A-�Y7�=+��{}����~T�ႬYX����M�=��e==�ȯf�89joЮ��� �I6?{I"c���n:�>�k�}�ۃ8A�/Ca�T�K<#�!��/�>y�z[@�:��<��>�.����4�V�1B��!� 8p��lSxN��]]���>�~�����CF-(�j?��łѯ�r#B,d���m�n�>8��ǎ������H�Ƹ���t�b��nPnU͊���L|i����O�8�Ǐ;|x��~&lj64E}r5b�A���߾�4mb�L0�4�bѣ#I��`��F�*�\�z��Fח;�����;�+��m�(��F��2Dh�,�F����Jm�(ح�E�F-�/�k�Zœ��\Mr��E�6���|Z�#��J6��F�w}],m���]5\��h��mMc��E1��4����FO��Qb��b�1�U�Ϳ}v�b�mE�:�z��;�FBd	4ǌ`��9���n����g���Sj>`�|�'��8�B%�lR��K�"���C�Uۣo�R�7sӍ�#�,���]ي�3��j�֐B)��!&�5be�ÚUv!���a�us`�)�/���(����p��dC���R5T�"��A?=��A�(�m����*M��ηGcj*VnEΖS���l�d<o�3�0���"�2z���nZ��"�fO����Fh����-G�_�6u�LL%����9ʢ*^%�ln�m���j�Syͷ�)�5��蘿�v8��hO�{q��H�I��қ�$����}�a�dm{��i�e�7��4e��8����x(O�AL����<U��忟�׮��"
m��Kebu�X�=������U8մ�㮓��ڠ��`���3hl��h�l�g�f�iG�`'�=���G3�y�����v��.rɓ�z�1�rF{�>> ����-�&	' $��g�V8��]SQ�����޹�K�b�� ����w8�u�S=����~Li{�Kqa*����t4bZ:��v�v�B�v����;��=��䓄�f�M�K���F_(�����&K� �BimX�v���y�BMo���&�3@Ϋ��m�{ۤ�Uc.*�a��6��� �ά���ߛ\m��[��&�IH�׸z�Lkl�s�E�%�w+�tL3��=n�	2I��t��t��[�V��&����p=�"�/�p
��/#��7�<��m��?�y��)���������d{�8V3gx*a�%>J��m��bL�hz:,L��T:�i�LMX�i��u��]N_��#kZ���ݐo�n���Ӽv�E�$��0g`����6-�V���׼ԍ�BhRi ��gI��������4ri�E4�cf�[2�n*��6͛�X͆�J�`�L[�kձl����U�%���P4�K\Tps�U�lmE�艱Y�e�D˯a\��i�(E!v�Ի���
u����X�3B�Vl�\A��`�2�[��-�b5�Fљ+a]��Yn�T�åx),4e0a�1o7���#�a�b�-�<�����j��>7�T����b �vk�bn����Z7kT��+բ��=��	��I�J���{c�.a,{����9�ܫa�\K����)�I�x��c�Fs��������k�!��.�ԍF_PS�Eہ��k��2�>d�u�m�'$���E��u>�lUYQVo��c3�*xbd��.��]?I��Y�+����\�d��x$���z9��ǸK�x	�;75�)�w�i�on�I�L�Jj�+K��nc"fs�@Vޮ"�S+�ԍF_(�	�X�I������0>ih�	�/9�OeVͱ��]���fW�M$v��,/k�B����#BD[pu�L`�]����&�a���|�\n�ڦ}s�rdo$�mՔ�,Ow1�v��p�2 �Z�2��]^���T���=�����;;l�f>�
N�c*�Ws�,�=��=��,Ѧ��de'[��>> 4p���Z���f��E�,{�S��a=iM�4>D��}|�S9�M��f���޻{x�z��FbZ��sM���Q�
�2LI�X❙����a�bv\*̯O�[5,�O���c0�w�)��v8���z����n=w�r�]�B6���{&�]�k��(��P���-�n� ���D�<Z�>0�ׯg�'ߐ���a��5�9�XK�����F�R��3������#��ӌ=�%1�k�ӥM�\�l͵F_(�7����E�"�2��6����Y"��.�L�R`�"��T�^#1�b���9v88�39��TڒUʌ�U���@��I�L�U�ϑ==p�1`�MKr��$��|� )�y��_��6p�=ȑ��<�oWIg�`b�+��ܭ��NwL1X���%�c~9��M���۾>> G�F�n�l몜�P��	����S�	0��6n��iS��"�k$�u�B�'�m�2�F���[��9,��J��8������x]�z=wQ�u��k��s��gnƇ�g6p
�gߪ�ڲ�yi��M���JN��` ���
C��fM�f�Sa�m���!u�����g�=��#'��k$�I-{8�z���j���QWv<�i����˯�&I8I�z�kiC�͵O����azxԭ�zf�c/�pt�|}��oPr��+�'r�EZI��Kj;xK��&��9]�,!���L���)��e�J��s�ԹlS{V�I:�w���ƕF[J���)��;J&��l�/���emZ�%D���d��&e�inc-��Y*7"�����y�Q�6Χ(�50&r����3��xu��|@�����s]�R.	&�ܩ����0+�m��`��o1��8(O�(�I?���#��O��7-�u��4@ͷTbΫ����b������ ��m�]�HI�kr�Ƭ�%���͜:�ݬ����<��F0�	%�W���� �6�M�L2��,�|�����M�S+D���+�a$����5����2��I�I:X�Ļ��q�fX���1��8�p17�m�o]���N&����^�cs�RM�n��,����͜����;�(vؽd��*s=�]\y�z�����N��n���_�Z<{�n����\��,ʙJ@��ǻo$�ܹ�f��J�Qʶ�[ɰnl�O����=6���������O�?)��e|p��C�0�� ���zs'��׃~铰. ;�N0���2z>#4#��K�j�d�q��?7�徬)-Z����Ҡ1��G[��GFUet*��\�@Ke�؄��,��$�������P	T�L�e�ˀ�,ΰ���9�R!��A�Yn����4�2��c�a��̚V�ڶ��:D.J([M�.�M�`�5��i.u�$�����M�e�TA��:�<�d�e`�ttt��A��SVm�����f���ߧ�b��*\i��̌�[r�ɣ�׮��8i,bmp��;��{*����$�>)6��7k��K(���Q�6���e�:���T���y�J|�m>lN���wd���s6��2����A����T�گή������m�[��8�{2�B��P�BP�Q"�A�T�]ɩ��T��&%rI&	'��{/��n�l�xe��+�7���{����P�1nL=F�p~a��Y�m��z=�^f-�Æ�y�68�S��4�kw�0r�gL51�J o��XZL��)%!���ǐt��+�^�ʦ��B��ȕ�֌k ](M������vg�,�+Ӹ'e���0I?���̭~N�B�yX]��5����q��	$��7��e�-m�M<U�"^�1�).2�52�m��v�ܚ��*�+����g��z<x˔���|!�8i���T����9nj)C���T��Vǻ�||@�1�շ�ō��
�Qr�}s��p��'�(}�v}n�S�/{6�)���$�0K���v�;�ԕ�j��ۺ�p#��G�����:L�K�ڌ�T��@F��I.��,���;,hU�����1wd�u�X޻i�y$�K=�l3�������[�j�^���p��(�J��I��������s�?g�����F'l�	�V�H��M.���,2a˦�Kfx��w�/z��~F�m���-wk{С�gH������sF"dCW�Ӗ�$�&�I?�,ZlP�m�p���5�srvXЪ�0�z�%1Y���L)�r�')�X�I�'���f���6bK7'3Q<��3X&��eCD���y���8�R돟<C&�nk�>#|[�����z&�ݼ��7R�n���v�����A�tuh��r�����$�d��5����jr�5xtی��$�U�{���(P�\����0�In,�����o�	'�L�]����.�᥵�\污T%��O�~$n��۵t��[v�}��R�favK�gxhgg��J����d[A�rK��J��K(�:=t#���O���^2I�M��6��k��r��2ﻵ[�xM�cy�I��$�y�����b7�[����L���
�[;�'�aww��,5��X�+��N��I���>c�Ϯ�𵊵��d*u�:��M�?�Q�yk�c�d��y퇶���\�o_'��	���^#�n�����h�wJ�̇r��2�F��p�Z��x���-!�渚�*]�(��ix������4��*�
o�����-�=�e ��||�z	��$�$�]���x�0�a�zn�t��(FT���m��%��B�����F��v$�3̮�L��Gk��,ґ0�GBV�;D�]�iTjGK\8�4��7���xt'Ԕ�ݶ������%S�嗑*��=���y>I�z��}v�T�c�����v��uw�ov'���λu�|��ܺ�\�T˔S�� X]��$�$��z�~���Hr*J�[�P��}�&��뻀.��l8�u1�z��<<wH���JFټ�3���>J�@l��5wR�e���6�_p����� ׮�`�����3G��5#����l��+��Z*PY��B�I$��y��"���}ҵ�N_fѫ	�sާwO������z6��bo��4n�j�e��}-���Gp�Cy��z	 ���K�A}^��v���$�J-���KN1� ��Q���=8�;������Q�$n��*�/n�z��N	;�S4�F�}�3Ey2{ڹ2���x���G)f8%ig��l�i��A0�"ޞռ�3�e]�*}�^�~=�~on����Ïn{q�v�rҮ�Rޒ������wq B����/�[[�܊$��7�e�;}�B���1l4=�w<�.��:}�g�s�g����ᏸ=�>����_cC�hՃ����
ΡM��w���ũ?�;������|��[A5Q]�<�fp����<��]���Gyg�OF�7�����U�ѝ�^�PƮ��W������w�Oʔ�,$���I��C}�p���,��UOi��Q�y��dm���O�ecf8wU8gPj �DT%Ys*F"��W8�x��r����G�sV���C�Ǒ�%Uosq$���Lf��"zM�{��O�<����^]�[��;|�Y�+ջ�)w����f��woP=�^q����3��Wo=�;l��p�w۝�_q�}���w��{�n�e���+r77Wa�beos�`���{f��=�a|yƝ�l�|�]~���U�ߦ�*�X
9�J}<�뛤��M�v�(���}�Ŧvw��^���?_a��w�e���'n�|�#=t3���A� �f�m};��Г(��Y�G����޶��Owk��{���$��`Ɉ���%��l�Y�ۈ�����rOO�<������[�&ȕ%IEcZ*4lD��T�� <���N���8���۷oo�n��u�dE�������~���}}W{���l%:��J-�����x���ӎ;v�۷��o��cAb�N[j��j6��#L���d�"�cX,G���ך���E��m�Y���:�+���U�&��툱4To5sQa5%{�Q�:�W�`��6�`5H���QF��CF���ۓۼ�4��b����Z-���j*�����2Q��&�o�r�X��ncW��q5��͸V+%^k��m~�{�b���P�|m��F�H����k��e�!��|k��4QRI�0T����{��������t�<eg���9e�����#]��b���ۍ�o.�B.Rk.!t�Tڳf�g31���F�z�b�-b�l��S�J�L��I]z��pˈ�$%2,&�Z��]1Ml#�m]s��B��&JX��#�́��%�c7�l��ճ&�gBR؅Ê�f1�o]a�k��	��I�-4��&.�׊ԥ��i�C��.�!ؚm�4�g�9�AX.f�\l�Di��-�s�	l�ݝ�f{(չ�5Q��(]v�m�[z�`܅J\�*��C嘬��[4m���B6�MZۊ:�UQ֢ msM	KN%���Ke�54Q�,nh0̰�SX��Y�[�Zr:0e��(�spJ�Vh��LDl(s[�#M�l0�d�հ�V��21.�"I�)b��	Q�KHPń-u�jSFbb��h	`�t���<�+t&���@܆��Y\u��P������ 2�FG��%��ڸ������b4��3T�����!)r�S,�#�s�J�HJ�.�]��_k�,��C*��jF�j��˰�ՙ�ś�X���aЬc1�(��]�`�څ�z6�l��6[�Ph��C[�W(ً����` j6[�
�(e��15���ceg�/��!���!1y�����c3��[�J�3M�6Z�V�j0�1�ҝv���.�q4�J�=bCv���Sb��Q�:.��UU��7��f,���Q��f����Pu6�J<�v��W�`�,5��B��6��m����m�y��D�ک4lw���læ��f�����ڰpʃ6׳�1L��,u���[�p�3�]��!Z�]��K3�-dɃ@H����e�ͅIR���4î�lneU���4X��Z�R���1J+v���r՘���9�fG;We��� �Ћ�ؕ�J;CHL��J[��	�L�ex��i��G�i^rj����L�<����i��r_��{�޽d������m�g����sauZ�0�qKoV��ݒ�HM�[,&���f��(�k��\L2�.m�pj����a�Qmb�,�L�i��K-�!x�/P�d��`��L�F5�-+\�i�����s�"���+n���B[�Q#k�p��	Z˛�"�h!1�6ms�XXƔf`���=����]]�`��l����f�W~&��O<|�v���#�ۥ�كsr�3KV���S�ƹ#�l&��lM����ΘWc���2~�v_��aQ�9G���X2c�p`�Jd�a�L"8�5���7�eFupwlR�	��$STB,$�&I�N<�����/R�oVyC��b�X)QY�9Bq��S>*S�j�x�s�*jQ��ޏv7����-�]���NQ��L�v�cGC;㗉��>�L0	'	;��q7Z^Y��*mȌ����b��yv�5P���)����\?���o��?�JÆbƐEfb�Φ�&�1��Ҽ%��9a�����Ii��_����q�N'�8š�=��M7Eg,�ب[�UG�rkӍ��I8	0I�c@��t��U�`�p�3�64_C�Ƨb1i1N�I�d^B��	y�ǉ�b '�ph {�������o\:�|�(�}����{r�E4d&������­���ݕ�
M4�������d&�������mꆬ�I(o�b+:�a��A>���	�v"��
��0�No�	(S��3Y۲y{�({���HVc��N�h�9gzb�$O'�Yq����\�|��Λ�$�^�ORƞ��[�W��k_T�i�=�i���]x/P�~��|���){�O~��1�[�R�V�B�<�qYM�W%���mSB���~������蛽�ݾѼ�y��;d]T*�i�͋}/0�Te��{����JRj�̜K9�7'q�P����ոݓ�z'1u)����o��B�n�b冸LH���mη�=���T�&-�b�������Jf�"#'��;�����هw��}�Ѳ\nޘ���Y}��*�`w�ՙv�U��ۈ���0g�x��a�,-���IMY&���j�O�� �I�#qO�/�����q�K,ݙлk�;d*���z����k�9V��=��I:LI\�m{���_И)���2�j�1agVpR��$9$V�������۽H%��%�,���e����&"�<�փ��λY��h���>Z�Iy�e�i�>�'u�=d��oD҂��n�wȫ�	W��]ݏ?4�ugSO2���]��ѹ���d*���?���#��wN���̓$��6Ѯ&)�Jֵ���S�/:s�53R7b�֭���[n<m�Η��
���n�N�Jz�=���{��X������ZiFF<�eR�yVMU��~/�	^/��kvo��]e��1�st,����m�.�S4ѝr���j�b��o�������Ia��ñ��5�qAV��F�&2.�'@�a鮸��x]��/yک9�
z��[}���V1��V3j9��^�-��o4�Q�`�w����0q;D[�	'�Hn]�_l�.{J,^r����P�5T��!���䓤�7�ZZ��Cd�l�n�C�u3�7�k�V�m�J[��P����w:L��Xii���t��#��Kڌ�Ld]VL{C��T��
�BoG���7��뫑�C�Q�`@4�����lۆ��|��iE�Μ�	�x��T�i�[�"�stg����J_�mOq5�낦�[:!��!�U�o�­���'#s�ٯmD.xW�X`�e7H^:*¤6�n{���$H��i�<G�;ڸ4�I���5t�/�m]Ga��`��S	TaQN�;��z㍜�7F�)�ip��x��gnE�>��|>����K����+�p��.�M�E��7���S˼���ػ��U�va1���t��!B3L�u[4SUδ�Hh2��̎�k�c�c�!.�n@*�%m5,4�Q5,�$���"`��X�!��*���%r��9fn�1�-u�M������YX�p�lĩ��u�`�-m�T1��	�nf�T��j�ixY�lU�/�P�o��_�ɕ��GB� ��.��]:IA�\U��-F��lg�ߛ��. �o$�$�`��Y1�Ę���LvNf�6�.�m$�$�$�M)��ƉFv2�(�{�ƶ��ؚ�Wf�8	���Gg��)�d����G���I�`�E������*e�,\��Cn� �w����m����`��َ���52��|rs��;�5suY7�
[�xx���}n8�i��&�]����&�����zZ���6Uj��Myѽ��*S�n��	(��םݞ�C�,��������1u�;V]�i�fQ��6ČY�Xk��6�X�6ih���ޮ��'Y*�t��Cn� �t�lq���}�/���o$�.T�3����C>]�r��ܠYR�h��s��`j ��i&�l���D�Ǚ3��I�;
����jVM�.a��3U4X*�>�b��s���E�|Κ~�)L�d��W'���<�fL��I�N�كxe��_�S���Z���ם�LS�I��I/B���m�h��5�ۉ���4�m}WW�u!�� �w�0M��AT6�r����8I�����C�WhSt�Bow_ò�u��v�aJf�'Ex�+�����<����,)#�g~���}jm�Q���c��7r�yجi�J1�ZjA�^ � X�U���{�awo�]���5���,���:w���M�/�Y�� �s�%�s^����kk�%p����z��*ra�+�82��{n���^�[Ҙyn�	7�Ii�m�=J�ik���/�W=�C�[�Z�m����{
����g��8�5O��SC�u�vr�p�r�Oy�7��>0Lj\�.V��`ED�������zN	Z��7C
S7Y=PޮIJM	'*�Av��M9e�I�̹~���I�+kΝ=�pǂn�5�x�+�C���);J^ޭ����q���j+�eFA����$��8��pN)lz�K���l�����lN�f�j��2��EvJ�
eͩv#����S6b��Ϸ�����{�O�`	'�'7f���
S7Y4��΍W&�p�f�z�IO�i�8~Ƿ�ͨ�8�� ߙ�ۗ��<�=bk��`%Kݡw�'u��M��R��ky$I=^�ۻF]��s/f�	��ΊO�o������l� �q���K����9�I8��9�TݼT)�������F��z-Q��{�����{˖绽i�KwO����\>}{�j�Ǡ�K�~��{Ϭ�Z��㼜��n����;o;v�͖��>>xn��
�)�`�I����l�9��K+#��OX��:w�*_q(��P�oϿ?Os�`]F�)[��ԋ��3
�K����<��������������#%�'�u Boy$�d���W+���7�;#�~��f�mX=r�˗��̽e�O9��.�,��%��l�G��WwM5�
�do�CUs�,;�E�{�9��.ϙ$�$ͺ�s��ɨ`�**�nR�1=�t�	����0
�R;��"�����/gc�2R������ғ���V������¹8x�mwwiF��jd�U�!���M�9��O�#�T���}	0�xz�w�츧z������{�轫����T�L��)��(S��6�M�;T�b]������M�n�)��{��ؘYyi_m�|�'䲉��(�6�߽/^�'z����~�<7�M+eƊ��5�J\�v����-k�;k2@X�:(��	�l�92�*0Yr�6K-�P�t��*�\��n�E��`teՍ2��K���t.Ĉ6�e�<�kW���96�e�6�oVK��9eK����X��!���4m,���\Dؖ\Qe--�؄3�vˠ�(��r@9����Z��&����/��[����a�9�5�s��ML�.��g�(h�y�;3�xfc�b\D�����l�"��0kȾQ�z�Tb���؜��ܾ�F7.n��I������[淵Z[���q��8�]��2�.����J^'����u2�a��>�uIM�m�*ږxb+�Mm��J���}䒑~"�������!��%��b��xb��L׳=�:��b���`�U`�m��}
�m�I��JR^Qӕ����)�M��9[��2�.��{$��,��M �`�z�{s/o��[����KBD�J�l� �,c�, a[j�h�s�ZN/R�����wA�SP�#��[�b�*�{���I���I������	T)��-J�n"�V�{eڍ�{M�'5k�ov� Xu���e�g�#!§Q�b��Ŵ��P�T�VF��x��D<�>��ⱼ�ҫ�vz!(��Ӽ"ǯS�vA��A�����z�{`�p�yx��5�C�����Ɯ���M�m��m�own.ҁ��_��A?s�����m���v���y5(�|�>��;f�k�C�v�ٰk��6׌Nd�B�/$�dv�O����J�g6�J�Sy�;�!?�kΙ�I����֤���~?=��<��]��R;B�装��j�rsn��lMr]�x��Qc-�َ����d���OU�DbG*��ˀ5�~1<2e>�J��wi�z����v���׺#��f�DSO������g��z��M�h�a\��_,�ȹiA[x�7 bJI��,\��6�%�Cf;����^fC�r���OC'bC������<�~��s���=_s��s�p�5y�C;^]��̓}���$�R���-�]�b�0iŁ��&�yX{V?E|#;��=+w7]w �4x])���c��{{�Y�Dw}����fۨMq��O�}�qc#�Gj�{�3��~��q���)�_s��x�I��f��|�K�c~�Ǔ�X\�������*��;����_F7S����B�s[�$�t�U�������#|���U��L���u��U�}�٥du:ٹ�o�Հﻲ�|��Dۼ�B�/{��|�p˄gx�x�nH<z]��G�k5��R\��b�t����E�L�~-��,��D4���ߴ�ؼn�_a-�rj�N���t9}�4�}�Z�=��Qp��j�e���YӉ��`�9�ό�=�V�ɽ���-]�s��+g��(�׈�+=�@ݤ`���=;��Z63��� K�
��<f�ٺ����CN��;#��-���/�t�fٞɛ�4�/R��2Of�7�:�l�A�l�㞛�h%w=�����k�4�on�wQ*�ؓv�A{d֕b�M�:�D�e=�g�ݫ^��u�X�UTN9������ޭ���B����Sþ
�)����?aX��;{9�1!���Em>K��Q��\Ж������+�p�Ozy��c�wnF�%���8pD���/�����{��Es�C����)�m�݌��|x�����ȫ��8,�zO"�Ř�L	v����31d��\�cƟ	N�[x�P�úQ���	�y�*�_¾w~��v��������v���㷇 HH��XH�[aI�5�U�a	��m�=>>=>8�۷n����ߖ�~ڍ��Z4I�lj{�W�&RTDm0my������m��\ђ�������E��5|W�6"�Z�ōsk��\�ѯ��ί�Z�V-r�~���6�1�yW�o$�ny�yh�ݓ��ۜ��v;��3�^^c��Ū4Z+9��ۛBQJKVcY��/.ȱ�E�ߦ�F�����myW(�Ov��Eo���5�\�5&�i��4R|\�[��~�v�Q|s�����l����_%����� �|}ގY�����W���xo�n�)M�U݁s<�S;��q9E���z�ϟ5��]\��u�H�[u%�0÷�6E(�ɏH��LI$�lu]x�;N+p��4�q3�I��4T��N����O�75�a��z��߰5��a��K8S-���;BV0{�,�� �w��^ ,^3��3n;$�I�eOV��(���^gF��ƙ6@��Z���{vG�'&�M�t۱v���w���K����ĎU��]��[�vֽ�XVL�2|�n=#�&t�%.��f�9��n.�kG	֥1o�:+�S��y$�Ƚ�}l�1n������K����޸��ԯ3���<[ϧ^.!����N��a*j�|��� }fM�L+���.��=�.�Ͻ7����~.��f�ar_�/4�MQ������ ڷ�]���?�ݺ�������2O .�m�7+'b�I�M�޻�wwb�΄I�~4z�^�$��h�6�)����G&�8�	H��Rm2�L�(�aK]��!��H1��{�v�&$����4֎�Jb�7�A���4 �O�Էx�j
M�}wp.�oKđ����s�N�\�dgg7d>`��3�t�ο�s��yn<���o{��I8I��sp�7MM��tﴫcf�I�M��G���̒poR���g��1st���b���0V�l�
��/x{i7AJ^�;�Ll�=��أ:jnu���ly%P��o_��G_M�
�я�7ٯ�ׂ��΍��}�I�I;�Z�*�)e�c��[��M����wHb|Tؐ���36#�W�:]���+C�NՁ��]�W�V����훳��~o�~>��¼fܶ,���^�����OR��F�&�e-����9La���`;�1�1P��m���c����_	�sm"vl�M��.�51b���J�2���eYc�[Fë�eyj)�IQ�9������a�Dk!�1[n�݋/0 �iqe1�R�lhs�jC9ҼX�,.Ri�M��ф��H�rm(�of�+��iQ�S=474tV3e�\�i�ѷ��߿�RnƠ�i����[e��X��ͯ�Ie,�\̉()x��@�gޏjp��l
r�����k*M�n���4�o#�.��ʇ�0I�I�O6�b��gn�����qht^�N��o�*�¹:I�4�9��]��� "�&$�"4-��d@�Om�6��J�/�{��q�j�	��%n���f`����"�7��=�xR�zkl���TM�n��c:�VЦ��Ef8��I `��<Dm�4=�>��X̝�WAWo� �j��$f1Ay>� �hO���;`0�X]��4��ۡ3[�l�ڐ�:8�!�_�Ly��e	���y����]r�����aWn�ng{�R�m^�M�m���]П]���h~�1���ֳ��o������ b^;&��-�ů�����x��C�s���]9'-c��w*.�Д�1�� ϻ���m�ެ`6��-�싮TM�n]��jK�RrD\�����C�0	0I<���]�P��g���a�p�ލ�y&�����o�	'�{0����^��\�0�t���X��\�����7���٨��|�7��Es����z��.��g�B�]��j4�BB�z�kU֏_{��y��H��24��2I��M3�K����Ёa�.u�g]����K�a�\������R}~w}�^0I�I=�y�s�MÎ����y�.U;�dO���ҁ��|G�٭S�{�8�K<F	�I�����u��77�����9��vz`T�"��l�#x��U��'	0	n󎑘MB��2!^Շh���8�p�����1g���W�q��=�j��lڼ�{[���~f���7��~8��T�2�Qh��q�rF`f�1�g���Ο�V�.u$K�p�|;1�cwo������MM����怒�/0No�����[�L�1��	�i
�؏�Ro �y�%o#Ls1�L/nU,«�e����(	+��02wU]�=}iu�\�m��v`a�.T�&5�ц�.e��a�0A`Y�c��[�ǟ�&��_C�+/�R&1k{�O��O�����C��֔��y$��v���؅X�w8	��n
��6�9>=�o�S0 W'�K���T��ǈ
Z1b���'>�0�h/�c8:�
������^_F��E���l.��`�":n\>!9��v�$|�[E�=��X�6�.q���N�Rx+��v3��	��=���3͵�|��T�;���4���V���݀<H����.�{ٙo�	�Uq��ӏ,��h�3�
���P�I8�$�έ�6��3�tm�F�q�y���*�	�pd�(O#ˬ�?~{�<�<�?n���F��L�F�Ƌ5c2J.��aB�(C�v�x�]���@����ky$��0�ʹ��L���W�ѽl��C�����N��n7�I7�-�l,��z���$�x���>d�2�ܬ��H��k��E�{S*R#M�S4x�0��]�I$���cAU�M"�����j��?�`�I%C=^X�*%���^�Z���cz��=3�e^_F��� PvQ/�P��>q>I�7�x�O䧓F
�r��]�!�e�^f�bH�<�G��oV��[�Z�~���������H��{���<����(��\{��FwE�]�Y9�۞:4�t�z����-޸k�Z��]�)�=������Gt��%��}�������i<�;3\XT�u���֋vI@U�(��]Yv�%�4�ԍ��81��E.�vl�,FT�YA�J�]�5�3��[�c4�
����i�������F�KZ��s�+���R_9tW��s��,�R�M�T6�k��eI[ġxh���y��s�ZL���2�i. )k�u`BT����*5#V�֎�t�b�&�"������q�?��_H���bGf��͍)��3m�t���e�]-�Ts3��a��K>�=_L�y$�lؽ=����W>[��p�u����R�������}�
a�����cz�g��c2�/�{��8��d{���ݺ��L�I?�$Έi��n绻<#���.�$
�<��Z�	'&	7�n��\��׷q��7v��.ٻ��C�<�nپ���6����������ݰG��'����F�2�U[�����ey}��D'�o$$����/^���}���׹�����a�S��-��
�'7ͥ�G�-�uj��H<M侾E�<���F~~[���Y���u��*���̶�j��nn�z����X$�$��=�c���Y픐wk$���TW3�������u'�rj?�˖��}����=�T�}gytVaɂ��P��M�5�&������x���_�V�W���7u�\Z_.7�*��T'	�"2��|L/�Zd����,�c��I	uɉ�z�+�W�� s�q�J@J_�I�\�_!}�Ȋ��1����9X��aM��s���R�U���珗����w����{5�	�p�R��-����5������k�����E�Ӂ���`#�o�ͳQ����,b|Ct�	|߲���@a�֩5�Bg8*��R4�\s.L&f�6�H%����D��}��N'��w����ɪ���my�[�/|��^�ί8�awn�e(��8X��eX�a�^u�wOE�*]�?��&I>T��vC�Mny�~E�[��I�`�S.�l�sIp_�<̧��Y�y�7P�<�M4�����g�uX<���OYivu�Y<��I��ǈ�6]}q��^�;�>��V�)<w������2���Ϋ�[9S{�?�`�y�����K��ګv�����t�דի��2jk˼����'�9{X�l���e�m7�rS>!&��XGk= C8�h�1.͝�ț)���]��(�J���ᝐ��E���	 �+�������#{F��Lj��-jV$�h�.��jZ�h���>���8��y�v����/9�����;5kX�ES�Vﺵ�&�&����8�l]����p]L?rp0��V�ݥ���e�_@�<k�>�f8��-��T�m|�Н[-o$��7�-;��;T�r�}���2�.�H�+�܈�-�Y��o+��`O�|w�]GV��x��*r0u������{	�#S�{�\YL�`�.��1����,^���9����f{L�-�޳�s�Ç������	'	2LT���-�񛊋���-��i������=��ۨ$�5˳�e���˳�8vx�C��Ue����5�2d�-��C-(�Ͳ�a!as�~�žZ��	7���M{�/��8SZ�	��*��@joO����V֭ƵM��ڔ�0�o8k���*�eM�zS�):QN궥����/\�{�-ޟ]�Žں鲃	�s�z5�1�Wy}�k�u=�@@I?�����K���ȗ�8 ܧ�cy&�ܦ��iZ�8S]u?v��!�pV�����c�bh�N��	0K��L��ۺ�+x���ɤ�g������0��?���G�_��DUEk��_���2 " ��G����ʤ u��H��kfUYY��Z�5R�l��Ym��WYU,��[e����YU,��5�ͬ�[,�e��e��[+-��l�[,��*���e�Ym�V�5���Yk,��5���f�Ym�Z�-��l�Ֆ[e��eT�[,��5��l�j�kee�Ym�V�*���f�Ym�ke�l�[+-��l�U,��5e��f�YU,��5��[,��UK5��l��,��ke��e����*����Yf�Y��me�R��e�VUK5��l���`�E�cZ����J����������E�����
����������#J���
��������
�����
��������
���,��� ���Y��̙���e[ləU`�Ej���c1EX�1QX1QX1X�1AsZ�dͭ�f��U,�+wcq����!���a��"���db�`����
��
�#@�*�fUK+e�T�m� `� v���2ͬ��Ym�UK+e�S>v�T�[{�v�Y��Z���eT�[,��6�f��9�?�]������ 0Y EH��^x�w����������O�?�����t~!������J�*�w���|����*��x~A������E^񀊨� ��~������>��柼>���UEo�����贋^��6������N����?��(��b*(�U�A@$AUA�TYAIE�QbDQaE� �E�E`�X�@V)E�DQ`ܔ�-E��bEE��Q`�TX�"EQbE(�Q`E�0TXE�EQb�XTX�DX�X�QcV,����k%T�Y�[&�+lj�k��Z�_=j���~�~d�eDER@@$A@g�p
�O����@�3����@�y���"�+A����}�y��\��M�>�;�xC���>��U�>�?J}�?�4�
r ���PETW�C� �h}����}��"
�+�
~��Jߥ�3��KP@�����}Σ렰4�QY�!����������I ����O>��/�?1����>�� �O����cH����>��?W�*���ٰ����h�����|3�N��	A���[��;\�ω�9��lU�($�͟zR����������"���:`P|z��+�u�o�s�����)Ξ�1AY&SYn힐�(ـpP��3'� b�>�         >�                            � �                                      ���R��
���
UJ�B �TUT�URR��
*��$U�*A@)J�	)$��TIEQ@| ����$
�J�x��Ч�P���04z�����y::�`����*���(8J����޷
�ـ   �  \7�砠�<C\M P�U\� ����E�(  q4 ���R�u�sj
�)�@��p{0�tJ�g^��޷P     {�  |})J�Q QIR�'�BB͂�3j}��rb��Τ9$��N`h�Ew;�mBO;��T�%I�U)3ڎ�Oz�H    �  ��pt�{��P=�"D{� �sj{Ϊ�J��zj9�r��^z�T��'{u��z��=�seR�m޹�     |   9�$�
�P�����QW��f����*���[��
x��P󒨫 �m�7�7w(��
M X����p
���   �  �����*!�& �� �f�n�*�n�
�X N�� ��v     {�  x� IT�R@�Q@$����@�7`�(��u� t��l � �`�@    ��  ���ȷpt7D�� ����� gڝNv��)΀� v�`��u�!�{��   � ��R�J�PJ$�
��+��� d��E�:{9��p�� ;��@n�8�Y��E��
RY�"���9(��`   � N�%L���>��p}݇�v�-���!�$c�R� ww��p<@����C�w�!�~�&ЩT& C@�?M���   ��5R�hԑ�#�OM*��IQ��i���*S�4��d��$�I=�T��z��N�e���G��rI'��/g�'��n��?�wF���@�f����  BI��mm��窵km�5V�m���D$� HI	�����������k�u�h���*�������tYPC�.�e�Ǧ�R����2�M7b�\�W��Oc�=����CSvᒖ�X�t��V(�0p"�J-�ص!��U��ۼ�� #�q�����T�wN�I������X�դ�E�T2�w������ysd��wop��ZJ4�B��C�6�8*��&��R����ILVJ��&#x�Wd��el�[M\�E�t4Y�b`�"�ӻ�YJ�XDî�QЈ�e%t��X0�ڕ�Q�Ʃ�U}�dҖ4�l׋,b���Z�����U�G6�2dub�Kp�7fY��YgP���hЭ%�X)�rjY_]fTo/n�*�ke�j�U�p�8��"V8�ce����,L�w�]�߉���fff�Yh�mU�s[�4��̽�TӓC�͚W����v�S��x�`�e�F�R�v��m
աa�Ƕ�hoKCL�cY���%ǫF�CF�Ec��ǰB~9*�$�e�7�r��懻w�u���5Kj�/*b5�t�U1�6UL�d�ʼ{zi�"t���9
��[z���/�P+M�ӴbN��D�ѵ�aM;�#v*+v�G*�x���iC*�<I�*e#��RUop�p]u���Ug�@�Y�5UV���A0�������pÓ&��L=�����	VB˩Q+XV)��{Va�[���D)Z���8ov�Ѵ�"^���5�0���ܡx�8�A���on��ov�&Jv鷑�t�h�Ρd�b+�f��B�7b�r�b��<:J��l���l-4�h̽�+F�U)�����$�cq=�ɺR:m2§��'M^�Ƣ��lY���w4�N�.��X��%kU���J�\wL]��,�%�N�ѳx���f;!<�Gm�ov��*�ؘý����I]���.Q)+Y���/qA�����ș��,8����n����^J8�U@������Ȍ���lv��)4�^d�tI��u�mP�/1ѻd��*Ƌ�����@me^��U���pj���m;5T�&��V�w��"<���6(^J��Yf��ћz�T�5bPmn�>�<3[MM���YgE8~CC�*��ks�ȍ�S��fD��sb"�X�CZJ��iZ6֐bt�����J�Q���8F�$#A:@�D�U�V�˕����1�yd��F��\���ʄ�de�*��-*�:���[��m���W������Cn�)U;R�SR�<;���+F�nB�R���Z���*�8�[3E���x�ŕ� ܼ��ɦT%$0�UWzr�stf-:�+��an��jZ;��];�2�iXd����Î�#�՜j���b�(���1���o6�ۤ[�/��kku'�St�V�ªm����Zǟl{yx.į��ܬk,��8��XZlћzP���V4ƕU��2�#��#�(k�w�����9TqiW�]ܗz)b�J�iI!�j,J�튣��+j%&ejJ���T��ZM���ڡ0^��yw�����pǢᚊ_���oC*���Z��L����ݠ�5CݗUJ����^kyI]���"�]����U��5drG�7�M�$�D�vŪ�4iOK���ŤKM�+w)Kjp�
���fP[ڍYV��B�e�̕i*��1麊h?aL)r3��T�Fܗ�Svp�u�*���(՝��)R9 �r"�"���Y�F�PE �Y{U�����QŲ�%W��֘M[�BwV�35�:/*�sY11��1�`�y��i�U�6�[���n��*���� B�g!d`[Ud�Ǔ*o>%��|ϻs����{ߪM�h0D��5#ڒ;U(�LڙJ�sj���Ye*�5K����V�ҥ�!f�T�fiق�,���jC7�0;��ݬD��c#�UQg뱕�#gf�)�����j]���u[L_l�T]�LJ��}$X1��Cfl�l[
�Q�Yb�Q
Y6�w��ܻ�ъĽ��sv�E',d9��F*t*��3�TP�0�sm��ɚ�J�nfm���ɐ^��1�xiְ�^=1�VJf�u���VN$�)�����T{��2��j�M�کef�ĥ���V�n]K5;T/n�-L��f�3\#w�M���e
�n+���b�*�U��׭�3md��+5&�d�Ī#Z�c�qm�+Bb�¹&(�/	�����3siQ��4�$�����6	�z��8�G]��^����P�i�;6��,�E�YE[�Z2�(Ъ�m\��Ҽ�j�F�.�XN���p��P@��X����&��J{��U���H��FL��R�]+��.+'e��f�EE뻐�6]��IU˽�KB�,Ʈ��U�\T|͕�#�wm��c7��G6a
�<SL�O42��$�sUe�Y�Z(2�ɕ�V�ʥz���X���\d���*��b�՘�e�R�h6�kefی��6ؓS���3���yl��˽[��5���%�)(nj�6���	-�̫�5N!x��,�y�#�x��bڪ�s�.�,��:���­wZu����&܏9�V݂��A
H\���٥%��*�A�]��2&]]�F�Ʈ���\R^�.�Vӫ)��{�Y+;N�^]
�*�LL�e��P�n;P��c���ܥw�^Zͺ��:(F�JM�)�x�De�vF���1qmKid��n��*<�0v�%�6Kj5)e}CkD6]�����&Z�X��Ը�O���.��՛���=��e��%a[wa���]
F�mj�qf9�]�UL��;�R�Ͷ���� �-��T��sk2�����4M�`��:�mV��/I �Q�&�ub�`��P+�u��Ŏ�j�çDU���l�2�PUX\Y/	�:�
��K�3�B�b��3T���-O�6�LmG����"�T�(�!�d��E��w���^��3D�֖2m>���㳛&�۹U,�C$��&/DҲ�4�h��I��BH���p^�{J���m9cTW�����T�y�fn��[��%��t��	�5�j-���9�%凉}Z!-%�@�j�&d�w���N���j���P���I�vN�l�F*����tA���hS�y7n�57R���U�9'��a&�nѱ2�6�³4^��"���-�	�p6Q$��aՓK6^�f�T��[�j�?1kn�:�Q�E�Q�ѱд���D9��ؔ�බ������r�7D˯���%렮3I�WZ���-�m�ͼj�
Ǥdj�Dj���-R���Koa��lۙCr�n��F��.��#pf۹ae� �o-��b�#ǻ�h�h��:iS6�BU+MmJ;�eM��uWvmP��V�j�%�#2n+Li�f*���yT�,� �L�{�R��۽�Ud��h�v�	��[�$&���*�*��l��5=st���Jm�Q`�
(;c2^��`�\E���1?���Dѻ��zn��wWSv��Ks�UMM��&�i���V%��J�Ņ&=`������ǸsNY���`������;�^U�U��)��"ɺִ���f�,?��6��G@Z�f���4�F����9�K�N���d�i�d@J�Y6$�hbH�,�oV��1T�Uc˪�R�a4��n]ݰoj�p[UǫJt��'�EД�mXB��Ӻ�2(����:����J]Z�re锞&����w�g3��4��*�Z&<(U�2�1�ʎ[(��2L�����Y�i�R�����Oh��w��'�&-Ỷ���F�y� *m ����4h�Ef�j���7q�[E,x��x©��^�ʗ�7n��gI���yʬv&5�ږ�ӵ�J���T�I��q�U2��;��wwa�լנ�X�3K�D*ӕrM	Uff-�(g�ji�v��)	,���P�2I�I�a���SKwc�s����l�՛���v��ٺ��J����lD���]M�W�p���1��I��h�uN=�XSZu)Gj1����b�;�Y̟f�֓�"�WzN�[�U�oE��Rڣ�C*�Ac�o*Ul�d�kb�����\�x��73T�~�([�Z�2!V����N�nl�[J�2t�S1�a���T��W���(2�V`_`��˚��$[r^�e�%�8㪹����jWX2X��;`�yL�Y�z�>�r���E�m�6�j�j�P��1���g-=��乄���w��p�J�U��,��f�~Z+F�f*xeK��1�Re����CU��`�8ܫ�N|s�H�m��c��O%m���Յ6�*=�r09t%+����VX�jXy��$�(��63Dh��V�^������kڻ�wuzYnnU��u��S��e�I�sj�h��I�B�e�H�u�[�[l���Cnn^��!Q�-S8�B�����o"�43X��M���U��ym+FS�p�f�R��v��lV��A�B\əj�Z�m�#"��t��d��������!�ֱ�EZ4���:�Y	J܋-�gsi�����di]�������2����̬ݩmݧbeQ�`�;sG��5X�H�r��SP(�֭���d�V-�Xl�#�0�Q�33am��ا�`*�ȉ�Pl-=�-�uC	N�8Wΰ��m�j0m�[{U�]FY'B��2�G�U�p�:;��U���Z��Ut�.m��-[bΨ�A���Jg�[��-,	gd-M��f�a��yz�z�����KT�^�.�}sk6�WgP�_��������aj�T�PY�T���hi�j�7�Tx]U�w����[q:��7-=�7hT��De�bu�e1*ie�Y�Q��SQ�305w)��J���5��)�gV(m����gBXB�l�3���p�ܕ����bXA�GQˤ����j��]�������K��te�8o�Yu�j�C���֐�&^R��]R�y,����X�6��CܼkpLa]�h7�ddC69uE�"Y���WM��ӡ짴*hܓkl���Yc4TC^�b���s��nB70ѷ�����<6Ȑ#{��ujdr*#75��ԭyf�ۚ�w�G.E�0L��o&������F�Eq�Պ�L�F�A�Xl���D�`�&⻀���հq�=t��Uz�Y�TK�k���י�������*�M%J�]�C����
������ݬ��yf��r�1�6�eT�������5�݌�����]�d�iLV�#��8I��+^-�,��
�YoUIU�Z,T��锋�k6CY�D�ʠ�U�ջ��M����������JQ�c�k甮��X�ļ�p�4J�Icڴ4��퉽��UUq�aLQ�hk���)��n���@�B�h�R�)�U�E��&h�cUoC��UM^[�r��P�2��Rͱ���Iz��X�Ҏ��w3)���|~R՗�KA֜�-�4��ى7�z�i�YXN�M�4`�j�%�2l�D���4�J�,ё]�ygk*(\.P���OV�tA�J��Y�2����vrT�����͝C7&e�m����&^`��l��f��ţ�R�h��vdmވ�`/q�`��.�=��5�XQG%���ٵ��f�N�f�]3�nVڬ�Ph�k1oN�$9������� ���QFQ���f��U�_ْ-B�2#�n^Vc�����F�#M����D��d�D�m�'fɰ֬үn���M�od��Y�*���1�O��Ũ�.���]�+�BGs.�Pa�{zwbAQUor+Aji��ʡ�mò�͂��o2�V챹t2����c[u� ʢ�&bÛ�&��;�*�]Xs�K

��7�է����ff�+R�D�ncwS�r�I%h�5Y*[ɺ���V��Da��d�ʻ�E��h�*�h+���u�$��6�qGH�a�Ҷ��n��,�K�W�B=��D@��j�N���˺8��x(ϘXX�I��[hA��XZ�c.Y�P�M��P;����l���/дl��C.�ݲ�7V��9s1�6�f�4�I�f�D0�2��cYv��{�I%nݼ��c4�R��Kq@��5�w�P��K�P��)0���Si��1�����p��VR��`�UJcj�݊�ʠ�ʧEVEJd�G5c��\̭��x����R�U74C̳f�m�&ռQYI�8�9��s�2�g7!D��L���8�ެ�ۖ32��\���n��+4�<�mYպn?��	-M`��k�3 y�j�2�卽�!6kr���\���l˨��ݘX�(�S6%�F+W��cJZ��B;[��W�ùz������b����ڢ�f^���u����ݵZ�B.�l�f��쨛@��9E�f̻ÏN0hiy����uGN显��e�S�ܼ��V�GZ�r\mlQ��Ŗ����Yq%y�s�7t�<�v��B�4�d;�dں��L0�[i�n,�l^�MK����tc%]S��R�jrf�ܨ,����a�r^��KJ�Sn�f�֙DZ��ȆQU)�F��ɗTL�ZkK�*��q桐<U��-�qT?W�Z��Q�i�WT٘����1�ڼ���,��o%)�4�ee=��=8eJ�T-uj�.��d9��ի���h���[���Ó0$��͗z�R���b��#ܩhl
z���t�gf������ѧ0M�Ԑ��wJ��+v���b��^�Q�Х�Nh�!KI^R.^�wM���-�z�b�{���O�uCf��+�f2�2���v�#�{j�a�j�tf��b�w�%*����$N�J[�jUb��nźvn�sj�[C/e�cjmi��Y2�?j��:�A�Wk,���ӊ�j4�����Xk�"P���Y���U&h����b��,���׸���t�Fʘ-T[�D&h�MmbY���J�����&L�%�� D�W�*�4��[�"hR3k.�ࣹ�oN��r���5v���][��7���6f8�Ch�	8�2��2,����J�f��\}6�tE�W�U5��D7FeQ���6��k2�Ix�yf�a(������(�-Kx��-��m[up�b��UX4M�4̗������*����8�AU
�Qߺ��ڊգV��Z-[E�j�j����m�Z�����mlUm�j�*�Ŷ+Z6Ѫ�j�ڨ�����E�kmZ�Z��lmkE[bձ��hت�kX�Tlm���Ŷ�mm��b�Tm��mF�UZ+V+X���֣j5j�ڣZ�mF�6�QZ5Z����mѭm�m�T[Z�TmQ���m�֭b�-mQk[FՊ�Z���آֱmFڱ��-������Z��-U����mj**�5Q��Fڣm��ڊ�F�cU����5�Uh�mFص�kZ5�EZƵ�-j��[_��>���G�/?~n'���(ɟT���5'NU��*��u�|�(C�}Cz����t�#%K�Y0,�U���Mu:��')��/Om��&�O�Sp�
��/ ��mJ��Żj����w����Q][Qְ��{��P.Ro\���|Qz�I�eu��'{���}P���7>�yˈeݺjө\6[�r�o�����n�h�;{g.��J�c4�x�n�&fӦ��.�s�/tΏ��N�V�ZtRF�Vdݾ����]��I����Ytt�{�n�$��9��<Ƭ.����x�`#7.�y]�d�Vܨn�^��,΀���B�O77��]�ݐ,�f9SF�e�P:\�ۣ�/#�w�U1�&n����wkk(��0�J��Ҍc���~n���j�9�P��]$��7Y�4:�o,������wAآ�k9i7ϥTY��|�i]�o`�z�NUc����6�C49Ջ9�Uk ���8���f1t%��b�of�VE,n��ٷ��OI�y�j�h�{�ﾦ�,����\�H��j��`J��b�+u��N�}���]۳�a_
�%�r�R�^|�.���N�Wg�V|��%X}�]��g�u��?%B��Fr]�q3tj�Ҭs+ʈN�j��B��B�N����CpJ���S[z�-ܸ6�;++��uۥ�-6��#S�4��TL�V�{��f�7܅����q���Y��N�=}sV�����ۧ�6�Lgχ1�F����|��J��+.���kq+�N7yh��V>v���mg,܅�������o&)���<�Yi��naO�d�U�w�Wo��*�^a�x��=�I��PÏ3�^v��&8+5A�j��ޮs��Vc��-ӭzNX]{Oj���,*�bUi�>��X4��Z�^��f�a��\��d�����Pj
����w{�:L�#j�ƺ��Q�p�jX����z��{���ϙ�Mu�ZZ��7G P��wm�;x�6�RJs��o!�B��r��N�6;E,��Ϊq����g5%���N�{�Q��\S
㚜�_^��.�R�ϊo�$�nh�:1I�Y[\����Z�7�N$�n�1���%w%��_.嶍Jڄn�[ס:��ngŜ���圄ʬ'z̩l�������J�(Zє�x�t��c�~��r��h4�����}�����L7xWf�W+1ut0��Q�����p��i���k���g��v�ɕ���N�Vt+�	��C*����l�&�7y�pV�U<����\1��ڄ]Ҭ�r�d=�]"�2Eo�@���YP�5�6�Q����Tj[�x��-ǕԞ��O�5�[�ͩ�X���goJ�1�n��]f���0LR�e5��|{hiBͬ�[�ƃ��-ӥ�UG\k��b3����U��4UsF������r]��շ6��T��
ב+�+�Y�^.<�]�j&å@�I�,�SVr���n�t�M�[��M�Y�t�닋kl�7i�B�ʔ��I��R�Y��ɔ�R�k/���oqp�aV�ʠ�=7��w%_3�7�q��=��5�ϥ`31]:�s��s�6�WZ���tÛB���'.NrГHΕ�����Ý͝Ip���R�ެ���=���8��:�e���ֹ@jӵ��jkwL<�򂬆W`�7&�Og1^n��(���Q��tu�QJ�<�T�s� vc�jEU`����U��2�ỴЃ%	qm�mS.�u)-%�'��Vc�\�W�.]+�r)Xn����6���&�%*��s�����Q�H���лK�#UՄf6(�\�T��N�]'W틻aR���v�/7kFt��X<+��5|e�e��v%���y��Q��b�W�h��c���U�j�!L��(��ܹ�����7FF�n���acl�8����M���m�Vx(j�h;w�.��Xz�fE�r�jY��̓wf��-�F�+����Ǝ����f�vq�����l��ܵmU���d��f�R�d*��Ґ˜2��=Z�]n�k�f͸��j=Ts��\���ꭘhY�|���Cmo:��,�g)O��Tni��]��Ue��/��C�	��eJ	���\��s+�r�g�j��h���m��o�d�&��Ȃ{��Oi
W1;�5ͩO	;R�#V��_<��AQCpfS���V������;�NZ�胚�Q���v:�ݻݭ�6-R6FX%��{Dڹ��	]WK/�'U�]+k8ޫ�Bʌ�ћ4��ͫQmv�;��\�/��W�]uh��-��e�'���5}]��fZ�.fV]�C]�/'q^�S��-�
�F�����ڜ�6v	�
���í��vnS��6�^WmPGMކ�M�U�dޜ0���(T�CV
�C����h�����X�E���n8͑����Q��r�f��*tz�}-���v���Ҹ�Mi�d7f�t��zd�y20o���#�)�;�b��\�5̨iϛn@�F��{�4�r���F�u��/R����P�����wǐ�Qӛ׽�uq-4w��]����,�uL�����əˬU����t٤��I6�`Ô�g�nn��q���R;nIsOv��}�Ydpͳ{�:eƙ��}��z�qI#��2���	�ut����+1뜮8.LV����/�XmqM���Mk��̃Z;����}}�3\�+���[�`����+��<��Ռ����T�Uޚ�]��8h\��r�8�mK��AuG��Y�&�{�q���������c;�X�{w��X�f�a����^���̢3A�1J�_p+Ъ"�u���w
#�K�Sn&d�ه�o;T"�ʚ;w����ƎVA�z*���U]�����Mk��vmwf)�J�`ۡo;*�٦��fV�:Y��缆Lu�T��l_oi��Ⱦ�ݜw%H�ꝷ4����؎p��ڂXD��rn'�`�~qe�L�������w�4U<5�n�̫|9�̲�u�e��m�erg����۴��ڲnaLw����Wˮ��k�&JBef����#躶��{���mG�RY��˺�����]��9�U�:�y���au��:n�=�;d��wnrZ��l��.�����I�fD7#�;רZpJ��73���n�oZW.��͆WT^%+�B��{����9Cx@yZ���ض�7��UnYU��u�S0�)����q�Mg�^�o/p�`ՙoe�Č��7yQ�ƻ��ٗ
�)�L�W�α��k�]{�]���iӓvE�Y
���֣�al�|�E��%W�=��\w�����]f+��j�S��t��o{[���J\��UT���ҏYMm�׏)��M%Vk��;D�����2�%��0��vc�ǚ6�fQ�ʬݘ����ޝ&���mՎ��7,9[�e�ն�����@�mayGH��B���m�
�ks�u��W��n�V�&���9���1r9���4�@�x;Z�W%s ��7�7���y�{�ؒ��I��K�i�p�	��t��yB��cˮxfVh;��ts�Ǯ��_I9�z.d��s�=Sl�9�v��򺘱ՕY��ԭ��c�h-��ow7� 7�sj򵟷[��I1"u��݇eR��uC2Λ���Nܾ�ª����`��uW[��|�C$x�����"[�/y������Ϊ�Y�����|���dg�`�;��{4z:`�����Zn�pSn�>D]�15|�Ƕ����5��j�Z�v�|pV�NhCl���E�F���B���^�E�4���.�oyk�	*aVvHa���nL���Q6M<���������������໽&�h��{���C�83�UWEn�&V#do��np���IUw_]���ݱr4�P���[��Um#�����f�,��X�b�]����b�M)�q�0.�U5M��|�x�[�sv#yYc��W�LӼz�U�y�����5�qs�n���lw���yl��Fs2��y��}�cKʤ{E^�P��Z�j��e�c9W��GT�Gf��9fJ��tw{8]5��-���n��,��E0�n����^U�n�V��N],�nխ��R�;6�5ʴ'ef���6���$�4;]'�b�Χ�E��X0���B�҅�9�b_]�x����8bǈv>�����1��䛘��30e�����ڥ�;�1��-q[�y���|��R��X����y��pUî����P\���U�.��C���z�fm���mp�|�oh����=ٷju�	T)뵘s�`��3�,W}F,��/�l�srr�S��F���D�t/���Gp�YDJ��r�,�\�5�_aӫ��.�uOx��:�6>*��T���_KˣY[��:�L�yHr�n�4��,��^o3����c���o#V2<�wj�qtyV�8wUBS�NƊ���51��7�op��a��ˬ�!���i��b{�Y|&�^>Ӻ���¯2�WK�M�Z����D�Wx()e�g��P�Ů�v�˖DÔ�r���{B@թ�xq#�;�R2:���\�3��ꢕT�5��2��Vj����V��Q�N<���:��}zhw^���a�Mf���Ϭ�G����X�N˽�pv�nWe�k{�����6�V�ԫn��D`����'��g�Ƭ�������켾�x���@��{�_�%�w2��ku���I\���_n;rƭF�`=SO�F{���[�2HM���}(ɫ>;����;3����h��V�Dӏ�,w׵c�J�jP�lm��o����,�voPt�Y�fj�9u��]ݮ+�U��]��w=o[�5��u'5h�0ܙw7�xUodwy�7���M�.��eu�[gZ�.���\�|1+�M��zsZUl<m�d]+f�/>Yw�,�5MЬ�ح%_a˽����8*��T��٘kS}/H�!$�W��%d��i�m��o��^]��,�Ӓ�V�7b�i�2ۋ,�3+7�t/�8TY}���5A�c+�*�M�wj��;;���M�����c���m����t�C��^�]��e�g.M���Ow+z�P�����v�C����wyN]���X�n�/��]�a:����d���ڵn��,5�\�2�N�p�7V��0���\K�Y�%ow;6�݉Ն�S����aZ�e �&�����.ٵ����Y�0��]�fMͧ���]qK*V�:#����h���ۺz/Op�P�a������n-��{_-�����5�2;���XtvmԮkv��ef��}�V3�vR.�nv�A���F��L��^�;��Y{.��<�r��/JwJ5*��f_j�2�`y��Ux�ܙ^�LR��i��ٛgg<iܫ"��y���"�׮R�u��ۜ8�=�ib5��u��8y(d�E��0��Opod��2��V�^�����$�t3eI]�*E���	"�Dy�T����h�Ht��d���|��c���X�W�.	\��UbZ̛��2Uj��Qc�+��M��T�$���r�o�ne�i�;p�3��R���kZ�~���n�����)V��'s�=՗�rYǺwL&�յ3�թ�Q'n����&�(��,P�:/��D|�-���<t�N�f���|�-��5Z��خ%O�.��1m9���6�Z�P�H%���s@To*��,��hZ��x;m�wR�{n��6�]s�G%�f�j��	�����ڔ��K�o{u�۟^n��Kn�l-�ub�0��s���ַm��h���LXj	y�)��gug��b]F�e���usr�`MP�gq����>��	c�����Qjo
�W�|n��u�z�%vf)����E�c�94�<�zȽ�G�CWp�n]Q��0���"����أ��k٦�h����z$���R闚�r#BಁЫ��ƙ7Tm�,��3Y����:�X�����:����f��N㲎^
������L��;&��ʛ�k�u
]�nS0=�6�.q����FJ�0�QYے�P�N�]��3$�L�r�s�n�N

��m潺V��i1�ne�	����μb`�cOfnV^����7�j%�L�D"2���;6R�+��32J��zwZ�8��Ԭ�U���Y���e͹�!]ǚF5�-5�4���aJ�w}l��s���^d���^W]p�ᷱ}�T�/�۷b���Wu��5'�nU�(�D��l���CѴkX�,�ܝ[�tVwF�bޡ��M��]n��{��b�Z/.h4Y��S���q]�dP����y۱��];�E|�Jc����2��͓[��WWQ;�ݒ"iA���wo7(aٴ�k������Բ���Λ�N���e�H���ʜqb�+��ft�Ln��ܮ��\4/Q7w&.�t\�>��(Ld;�w�8����u�A�����h����k�f=�������kGD9.wp�ʼC���VK&�G��9�k*�4'5�z�L�aG�gv[]z��x��E���#����W:����&��@��ėo_P}f���z��fP�����-�.��|�e�\3P�ζol��U8�TB��j��� b�ֹ���J�j��g�te�`ɥ]f����Ʈ]�Bk���)���u�u���˪��8vq�Clۛ���p#��M�-��j��R��[]Snͼ��[|,�SJ��vm�GŻ6�7	T7��df^��hmuv,r�M�zj�r�([ಫZT�b�����xl-�7��U/~̏`��.Dm�*��j5F��,8X�y�tʯ����A�͙�w���	]�
�&�^M�������6�f�d�;1,�U��A��S�N���޵IM��^�\��{ٛL!Kg��X/7�g����I�9�ņ�H��3�^���E��o����<���o֌�ymҷHc]����N���Pʥ7Zˇ�Wk���m=t�����s.���Gq;%��Z��%ĳ\�M��Q�cfbD�,��:��[+��,�'�Ғr���f�O�����K�h̳{k������lr�l��o�m��u�{�'>R����eL��b�:�v��{�leu���G8۠]�J�G�;��4�a0l����)Ih�uVmDQ��XEY�A�v�����\��� �	%@ �ռ��t���cW5�Ĕ;�Ǆ�U��[�d��Q�Cs�SVp]&�imv*��,�,�.X��Ҍ�\`�^��j�N��=�U2��ѩ�S���G��%�jH����R��xa�m��EZ�V��N)=v6Gl��|�^W���Gm��A��sX�<@�ojK��-�R$\1E-v�qd�Ì=m��vk�ڲ�t��G�Q���eZRFk���W�<��H���Ő�n��H��.���gd-������bVa��]J�ًb6T�i���N��c�;{T�#�.���%pQҒ��j;\+��GM�wn]�{�<���=1��ny�`n-��z��u�M�n`�8�̽4C�1���ё�-�(���dr�u�؏\n�����'Ieܒ�ɣ��k��駪��Y��qO+�d�sn-�c��m��6\������:�A�[[�r3�)�p=7l�j����;#�;��Nk�ʀ��x��L��X^x�x<v�M��^���1��z��7a��nj˷n���v��z�pF��z(��b#V��Zy�ePl�F�w6-��78M��R�sΎ�k����b����d�+���7'F�
z�z.�^qf��d'<k���s"��H�qm�.	.i���I�u�J�i�Ϯ��/PƹR�y� P���"E�0K��Fa��w8�AY�;s��cl��D\����/k�R/'d|f���ݰ�O']W[W��=u�r���y[%��`^�!�2ę��K�[��{�շ[�����0�Ce��������e �N��H��g��l�sg>�<z:ѣ����E������l	��˱رeqs5ʳ$���k�%�0&��ɵ˝,�V�1.�T��ǵ�;��wps��;'U���N�8����2��+�nʜ+�luv�GN{�r��n2ăl6M�f��6:b��20!�"�l���aۑ�pF�]Ut�kI��뗭b�ݙ�m�q��4 �x��q9�\�n����SqVÔ�8�nb�;s�:62�N��@����#�$�����B(M�Ľ�����e+�[�c�b�#���u���}��w��ѹk�$z٪$C5♚����V2���8�c�0���y��8���nM����P�I*2�Z\��Z\�
6�$v��v�ǣ-�:6<����,t�G�2�5E7��u6��Ut �g����kq�Hji�]�a0�,�#�z�X�#�ȓJk	���!����<���۾���[Be��T�b�R�.i��������3ݙ�1\�p6p6�ۧ���%vN�ЦC4	Ϊ\��6M՝�nk&([n�:õ��e4�ۭ��n4[7K��疻h����d���I��r�×Gj7Mi5��rĖ�/G����{#�����^�8E|�ָ=�a�V�l�E��Xd�^�p�^]�e��ⵛ=�v6����\��uf�i��@�9)��"e��1�,u3bC��Ύ�L*�q��-H::�Wc�;������Of����jp9�ۀ�qȨm�v:��벝oS�	�j��>����Y�M����;\�;���u;*S'[��98��s��X������X#��ɺ}��a�V�C��W���u�����ĝz�n�v�VE��q�3���X���L�vҹ�Z�l�ua�� GK�
� �f�0JCEN!���Kn�VQ�D���*��ۂ�H������4��s��1@p�Cvvw��[��Vlf�;=v��Kr��v�Uvi'����c��^��K��`�[v�l�(*�;=�����J��:�E:͍���K�G��3k1��ާ�ܦ0�ǔy��4wjU7v7spu�v��y�^����%�,b�x�	e���ڍq�,>�ӥ�y��vƳz�F�hL�j̥a�Z�������џ�pȷ�ьR �¡)�ٲ���j���飜�&�v�I孳v������t#�$����.5�Lb�i�2Uŕ%���'v��g�x����Y��u�l��8|�V�Odު0�:����c��C/W�� ��69���q`�эn����m��m��J�����B��Rh�8ah�k4\��X;4�8hMtCvk�n�t���9�o,�Yz�VW��]�umQ�8�i�<\��:q�-�nK�Q[m)��Z`cMs,kJ@�0�Ko���s˼�x�Ӄ�x�N�Lf���S �ؗU��6i�	M�mN�y�^�f�nb�E�<v5�k#�Y��ں�ۏmq�u4!4��r=z��Ya]�\]����w2���=wض%���i!�2]��/L*�bT���k�YX�M4
�x�۩ρ���j9�B��3�@+4��飺�f�=v�r-�:��p&�*,e�Vn�Zt&v^�gq-pTs#ǁsa�_[����I��uvbCq��ƣۮz���úq�0�s�ں��{e.��Wj"�8ϱ\b{oyF�x˞���<���ݯ�����LB˹���wZ��^2�]��1�p��<�78���o)W]���I�kg����%�z�\5'�G}n����Y��(�r�;P;M�ᘖ�ݍ�h��2�����{s�r�e��W���[Y.�[��}7����	z1�Ӹ���.�	\`\]�ˮ9��kp�=�v���6S6ա�TH3�d���Z�[k��b��͚���K�]�F^.6���.��퇗jq����ts�sv��}v��=��q�uӓz֊�����K2̾5�7i9z	`��������f���- �F��똺9�7Y���6�5��bfMl��P�k���sF�ؖ��e�x�!-K�[a���e�[v2�[��#y�B��cf�tf�3c��m�6���k���N3��ݒםжew`�ح��+�QCtȼ�z����F�iE�[r':���&�/�]����Zc������E^��uv�Yp�\�HZF�ڍ����G��KԬc
��3P,6q�m�^%�U�,�$f�lAj�c���ݝ]''cq���˷E�ݢ9:�n��؄�;���a�SJ,ˍ����-�&pXL̯GB�̎�Ua/nf�("D�um�#�s�\�Uc�ksV(]3a�zHCY�b-��!�o`�qv��p�״�˞�u��3e̵⅏ike����n:����2&�7[�#T��+����Bƭ���y�#���h;6����غ�`qn �ј�f��ۡF�l�;9�t��\�9/	�i�W��j��`�V��v�k��4��:p���tu!��g��ܺ]�s����3v�v�I���ϡ�	�J�e�cs����{MX�1`1ÃPЖ!�v���wm;sagsօ7;��\ո@.���&�P	�8�,6�[t�*��[�-^h�&�k`hpT]���.&y{m��7P�Y��<n��L��9|</mn�u�}��	�Z�p��Yǭ�y�+�5e�e�`�0w+uB�#���������ۉG���Z[�ʑvܚ�ꆬ����7�6�.���[r��o"��nL]n���t�j��r]s�K�gX��C[ﶓ�>�֞�<hn���Η�fd㍏]mn�A=U�nդ��[�AV<m��nk��E�;s��h�al�a4L�,1��;r��^�<ڴ�m�V�����<��l���Y����m02:xQ�Z��u;��X�m�m͓��%��V	\8۶m�5:g���ɽR��1�����t��p�M����9q=2���s�����),Q���s�z���=f��X�*3lPI�gn:����Ѣ��s��ޟ( 2���v�&��2ʬrE�MtТQ�������ۍ�����T�g�.^���?}���R]�{jI��I�X��֊�`U�L�e�I�٧��̖�Sv4�¤u�eV1-���;Y]hgGf����Ν�q�Zk]ӝSb�#�B nۉ�E�-q�]7F8�=��og��u��n9��};V��#��;d�[[s�d�����К̣���1�=\�l�=�d[��d� �{/����c[f0�YM�]�q�,�c�K�4N���br&����c��\��f;v��4��)Y��Yl����\5��Vl�S/��u��gu����4�S3�s��;�"-8;F$�W�T,f�����p�ccIi #)4�qRj�R.�t9�8��[��M��hm`�\1n5�ԉ���z��3�n�"��V٘K�F��]��yf��m�A��K[�岹��m���y�Nٺ$.2�԰a��.�mX@��f�u�+�4.n�L�.�}��ݻ;���[TGZ���z��Nƽr�W�뗦��Ӵ�v�jݽ�t��c���T]t:���U�t�֮n{v��;��+baIN��X��h�A	����u�t�+�)��up.��l!�]2h\��Z���
d�5vĻ�
�[
�
]�t<�XX��p<��tk��pn�Lˍ=u�m�a.Q#���A����N�=Q�I
����uu���C���X)�Vi�V��+3N�dx�Ev�MGf�9�%!��k��֑ ����I3����5�J{�.���PFO�s��I�8;i������t�������ٳ�%0��De	6�j#[#�	.�`��s��q��=�4}͉x�h-����Ӷ��%W�t�!�6nk���:�ұl�m	�p뇥�7k9������CW��<P^�S���h�q��q§Z���7�� -!�k�ٹ�;VǛu���-n#I܄cp�nֻ����46��V�9M�p��s��6�u�/P����㥧�t�=z^��\�h�AE���G  @f���i�ԓ^��÷m^m'/#÷�����:��=Ul���3��iz��-nt���ՋpB�m�:�[Kj6���t�;R݇R�]n���S���p�ݭ=F�-r�;]UV��W6��6��ۮu�\�>;{U��h�h�%nh��r���ڌ����`�X�ʢ�-����ܫ��k������Ζ�$��H�0QE�J�rɮ�]6��^���5��Z湭ˎpm%���Ƥ۝7*wm�ѡD�1�A�&4�[�64�^��3ݮV"�����sq�U��r��Q@c9Ҙ]��]�s��]��#`����EF�Axt���{��h�"4Rl�}����׶�D%�6(�4���h%���7;���&�y;��N�l3Ym\Ɨf�F�b�13F��]�Rʯ[nrv%�.ձ\����W!6�@f�-�*9��@4ֶ*������m�j��ic��u5<�1�am۵�u������㴸7B�vI5Y-s��ӝ��.�Ƃ	H&h)Pv,4��۶ͭ�S�iZR���͸6�e+���M�s�P� ��+�lV83��8qf9p��y��W����6nU:!Ү���XT�e�#��b��Z�$�����LТJ��]�u��Y`�[9�ay�7N��x�˪evy"㨶(�`�&�lFb��Dn{nM�uy�W�v�)��gPI�+)�f�]mb��#��G�ՃOfP��������G����s�ώ��	oCrz�M��.�u���W')n_,���j�Gw"�d�gn�X��G���D.�f*fP���̖MA�,k &�Zg�B9-r#�ݪ�;��n+��nn��ܔ]2�B'^c��s�hci!�ڶl۟'��շ�c�����q<�;���f��:DR�͸R7b1�mc��E�����2j�U�`��h��k�v�3��n�j�����-��oj��qx����F�j�.B�cj������b᭒������E|lq�i��w�5�tk22s�x����gx�Z��rm�K1D�ib16�Cr�c�f&ZY�Q���0�6�'��6�E�����9���{og���-��EՍ�OI�=d�ڲl�yv�y7.� 2]��5]�,�]��Ӫ�9�:�]�:�q�i"���mO��tn6����&&v���6�`�� ��]��� !�6x�[�)hK]�;E#)�l��9�3�dH],���T���^�x�]b��g�¬U�(K<u�m�s�v�az��,����5�:m ]&�դښ������С�I!f�[ޮIuJ�@%abƋ^-�/Em%���
4%a#m C�=@coo+�-���*u��B6YK
���j���B�[j��E�F�Kjڅ$��IX�KD��Iee���e��`�����)�����Yb!�	m���( ��ʹV�A���!e����������u@[rqm�nj�>T+�GYN��\=d�/I�g4r����*�� �����YV�����r�_P6�U���� �"�hW��_� A�W�7�=������}H��)�y/}5�^�EG���?J�"�z�Oz�E����q��;���e��m	�,J�l;ͧ=~}s��r��j�ׁ���־n��e���m^ᘽ�7�7��"�� ��[تg���ng�p��<(q� �d�W��r��px⯎�u�,��mtXݥ�Z~f��=��\��n�W�W�(x�P_?7X!�)�n�{�g���F[f�Q!�����պ&V�k��=�����tàg�G������c�e�����g�z_����m��K6��H/=3�QE�A� �@�,��	n�???�˰����m�ϕ:TZ,�H,�nD�ܹa�λ��=�u�g��%�Y�ʂ�ţv�Y�ϵ�c�g]٩G����Ck���o��X�V��xW��|A؂!��}�Y"�y|r ���x����e��Z#�k����+��;�����v�]�U�O|�7�T!� A���>�t�CL���_l�<d�WŴv{���ݬ�v����k���_��^�[����s��{ԁ��q7�,dn���l��L�ve.��!�{�I��~�ך�Lg���R ��U���(��:��i`���w�m�Ղm�;t��Ƭ���;�On��Xj�*ʷO+���f�e��Xͻo;�g_��+��W|}��7^a/}��o���kY�2#��.wV#��q6��`�H(���;
�f�����+������j�mxA�~־n��g��8���`��+�.%�t��2-��MM���o�Ӣ(C�+(x�������_A��i�s�jz��lт�.m�XgQ�,u\��}Yt��Vv��o,��$�lyZ_-7[�}X�j?-�k4�fz��H��e����_��=��6�q,�f� � �.RYewp��˾��{W|}�P �@DQ�道�͔E|]B ���!�~n�Ch"u����jeyw����?[���n�
Y����u��n� �YzKU��OF�@ӱH"	5��7Y��6Ӄ���1�ْ�7fr�nüY�[�{��+�����B��HChmx;��ߺ�cY�3�P�w1���S���@B������|A�Q��r���Yl@^R �����k�����_s����A�T!�UӼ9���,]$x�{��e�_���ӛf�Ԇ�7}�*35�vk��4��4~��A���e�n�]2\�_Ix���ﶀF�T ����=����Ք�L�<JD9�h�g�W��Sw2:3,V��sd�cR�:�Ws����N����E"�u׃;��M>4��X�r�7j�Y�l�8\T�Y��n-��vΡ_7A�|�,��!���K;<Gw��ߴ�R\8������{-v�ڻ����X���\2�.;�Z!�����������~~��}���J	Dե��p�:���uf��^V��zw�Z�/%�Ϥ�_�����Y���,���?m�틬⽯|CyW��}xa�[_7X̳�x�AˣRW?R��^�5m|��!�f��y��{R��L�_d��D2���_�����ǽ_/��Q��u�Ye��+sM���r�a��U�[S��~��V%��X���q6����fM�uJ�*@�G���z�ϫ��o��غΫ�?{E%�й�����+�Ht��E䗂{�A}<.�_s�]�[�0#=��H��!��|�[��W�.�ݵ~����#�S�O]Q���
����p<;����dmr�ʍFC���y�)�d�;�_�2׵粳����3����_ϓ��\�E��H�6�n�ڴ렖7h2h죌b���K�����RK
hƽ�m���<�݅�pp���%
���E�C2��Z�O2�7>fw6���i�e�۵�T[�S"i��V[U�����9�c�vS�yx��� �1�:](i�/j(]Ng�Z���^�&�����Ѯ�^��j�;�C[�:����:%ܝ��v¬ƭm������h"\3J�5ƂU(V/8SGS��us��Df�T-��v,�&��_Ї�>|A�	e������U��ʻ�k�tKC������A׈GҐ ��e�[������'.K?h�A|;o}��==���.��������ւ�	amb^�+>�G��u �t���|Ct�v���߰_2��6�qb���i������m��
QtD��2t��ܑ'6���={��f�EL`���X?���g��r\��7H��/B3���>
��Ќ3,��ۯ́��\��/v�={JV[��J}�t���I_i��3�u[�Sꭲ-[��u�-��l�[��lZ�xŶ"]�s,0q{�����ŧ`�m ���@���'��?{��ϼX�z`FxPS�n��^��ag,�댳34hs*�q�9��W�q^�	�ѽ�C��T�s���l��IQ�.�f��?m�\ɏ-Z<U��z�s'Y'.�-�OI�uZ�.�G�Tԍ9��,�Y�={�3����8#�o��z����W�r �����I��n�4���+@�b�?I,sܱ�z��;.���Ê��'��� �,Y�����%��/sڗ�{��q#O�ux�AM��ݺ���b�|X���X�u/U�hcg,H!�B>!�����~���X�%z�=h��]��}�3v'e�~��NA#��4��@�20����x����G��Mh[B���Gnu���a�l�4�QtK3� �Qĥ������w�Y( D1}_$�����?N˾�3��ܯ����4s�*_��}b�r�@�
"Iv	����OQ'��[J��͸����,g/z��u��/Lg��j��ǻ���^N�n*�|����#׍���hs*َ;���8B�+�k��	gJ�OjϘ��ZÖ�������۪R�!�t�9���׏������r����Ma�O�r���ù���Co��<�"�� d��2 �����j��a�ԧ��`���X��������ۓ;N-�� �:W�;�b�����0\�A��҈vВ��m]k�ٍ���}kP�6���{���`����j���h]Gŷ"�T���^�p�v�
Mˡ�e���n�a8͹�zAճ�wiFk�B���?_d8�}Bw�>��@,�����['�D����3�ߪ��s��^���Z~����("!��H�5��l��,�<��K���׻���ۗ"�8�+� x�_�d����3�՛g�Q��k�u�B�+"J�*���fg��.���Q�y�mA3E��>~� �5��!����p��y4��Tw��٦ρs�_� ~��n��@�h�p�7�[��^�vveg�A�e"і_ǫ�B�]��Y٢�n�'��2�����{f]���	UZ*�h9'� Z�9���+ͿUm_��\�O�j���($VA��y�.՝^�ϻ.�J�:{��ٷo�iŻ_x��D��/�%#�0�_g�>���%�+���ޢ�nf�1�h�Bk�\�9�lvavEĨK��X���/ϟ{@��� �0�d��H���~����{T� �=����Ow����G�����X�%|�0���}z{��^vW��en��;�qd
��F]!���D~�/a~���B�S�/����c��Ĉ D1
��%�h��;�kt&8��sn�WiŻ^�����b˔� �
"Iv,-��˪�h ��B��dAc�}�=�ߞyL9b39�_v�NҪG��B8�_:����e���܉�2u��|,`0Y_:Ѩ�×P�^j��~�z� ���+��(������~ͣTA�'��-+�7m�5R���$D��Ң�ۨ{�	T��Vvg2s�z���6�4����^�1�մf���_Ă�aU�j�}uWr��6�l�Nz׍��Lr�F۳�v�c[��1]��֖���gl9z��J�u������r`�s=�)�Ј��u���&�rts�sƌ���U���Wd���+��z{o:��I�j04�lu��K6�ē���A41�DR�	���e�3��W<�cq�3��z�P��<�K�3VT��ߟg�ti�P�[m�%g�w�`�vb�ǀ҄G�����N�3�1y,�|�	��$���|CnD�e�ݻ�y.�Waś^?^{���[y���͂�ߴi�U�Gn&fhй�	�;ygY���Q��O�����Y�7״�m?UX�L�wܬ�JW��������ξ�Y�IIZA��J�A�G3�DH��i���� dމ��	��qX"J�a�>��8�N�eZ����C|~�X����;���%���qn��>:P"�s��g�v9�ѠΤ~��"H��( A��H��v*�Qjốv��i�|�C/c�n) �Ag��{���o^}������h$z��c`�,��6�u,Į���*�ؚ[�Jo7��|>�n4'��|�e�3tG�nYb�b����b��u��F�#�����E��@C2����]�T;c���];5���x�"�[#&i=.���]���Y^ͻ��%SAנ�u�**���cu{w�3h��e�>��<����/j�����|o6D�e�{w��p�Q�>� ��O�l�,%Y����w�:QDv�����!$VA��]�Jע�D��ST��yܩ���X�L#�}�� � �������V��z�7�O7�u/�̲����'"�7�&"]l�� �m��`�tF�,����"�$VP@�gWG�*{�-���݋�bO{�?zmu��6�+��(�5�d�?a��C���]�ieQX�V���:6��Ȏ�㓖hy���=���I��2vwYw���1g��a�m�7x׽��W���Y�L�L�i�|�?��F�e�\e���Q̫�#����j�Y4�e���A �ҷv�#qN*���`9��Aˀ� ��!ړE�V߰�Pb��gʁ/�VA ��/�|d��u��֏�X�(�����Uj5
�,�P�(�C8;��-\��ܵj����s*���0\��"��C�{�(:�Й�n��33��u���P�Bb����jU����򪒳t�s�FU1tv��٪�v�ڮEO���R� 6��.��L��:_	����.���~����s�4b���^g\5�]:D�*��Y(�L=z.�����gZ{gkV]�A�NvPz�j�Tģ����T'3��0vT���7�}Vꩈ��J���:��.�9n�&eЬg[	|�gr�[Z�t�)VH�V;�`����U�&��7�I��q���VxS�����5��#�����Wu�meU\��7�Typ���۠��{h��RNYg��t�A�+��ru����A�ue'[V)���)�|��4f�k#���K+"�P���ۛ��T��3B��r-��K{X��Y_U����5:螒�S����:�;0d�h�\wCP+Z�]�V�����h�Z7	�JE'��g
«]	���ޗmIQ�q�ٯ��7r��3.�������b6�������@�*��[x�Uٽٽ��ۼ�.|�U(��Ð��fX���ȫ`�w�vA�D"����\�db#��gMh�|��3�+:��k��'��.�W�U��[�CѐB�����^�ܗ}�AI�j�j����n��!2�vwQ�.l����Ьz%M�4:ç�<9��U9�U4N�c�j�%��3�Q�eΪ���u�ޕU��d��!.�v�������+���ř�:�[fg^J<,�_� IE�2�C`Ѥ�q����y�\��wusbM�#WK����T����\��wiwt�[�oz��3����t���]�wuͺP��Fܢ�q{�cr����h�t����0�5˧M9wW+��ʹ�st��f.�t�ˆ�]{�lU�r Cw��"<-���Et�8��]���6�!b��ѝܷ0�r8=�xb����wnEr�˛r5ʝu����ܝ���;�y��t��\�v������K�u�ܺQ	Û�ogov�F�v,]"��o9�+���[��snswyOv���\ܢ�Ӆ^\��WwX1I:�kˁ���:hۚ��<眈�w]���\�q��Q�Q'������ݽ�ޛ]|��_�Y ?�ZAH,����p)D��XQ�sP� ��� s�ZM�Y)��p)II�9���AHw����k0��H;�B�A�ޠRAMD
a���L�d���D9�4�_����owo�~��Q'�G���@w��i%D)��ۆ�>��������������<?$�$���h.�)�������0)���B$��p)	) ��s��>H,>aH�-&g*�s����v�Rp��A >̃oul�-����'ᕖ~H)

�7�- ����p) ���s��i�2RAB�9�,��?����+��LeU
��R�n=���y���.��U�.��=etqh�&���Yi���i�j�RAH,9�i��) �Vv�$�H/+�R肐O�3�H�}\w�/׺�8����I }�-< RAeq�}�9���Bt��-�r�R�) ���ᤂ�P3�ZM�RAd���p)Q) ��9a���R
9E���]���3��oߵU�) ���i �07 I~<ߗgvǚ�W��"{�Ȃ�a�$�!L7�\4���H(9�4�Xi ������zǚ� ���\>H)�E��) ��J}˸
AH,5�sP� ��aH��R
Ay˸
��_9�L�r����:(��?�@wƉ!U@w(����RAh�u�
AMÜ��L�2RAB��H,40���a��$��9�s��p:�[��L�����SݳI����]��TAH4T9�\>H/�������o���5��νH�E��
H)���) �HO������}w����ʟ�F���PQV���������Bfa�ݵ�jM�^CL�y�ޜ���|��uM/�O6�o۲�U_�f��)���� L�!Ԃ�P;�ZO��R��@�D��Ü����R@s�ZAH)�*��Ü��LHO��3����x��C��\�� ����*��W��� 8A}?w. h;˄.!3*�&fX�?}��o���2`n�����V
�.v���sX�0��-m�����0�V,��z$���?BB�(d�ި�Rg{�|�X|0�r�I�) �Te9ʁh��_)�88G�G���g��)
������_7��ޢ���$��I4�L;��i�FJH(R�H,40����
M!L9�\4��) �a���;E�����:�Xi �r�kTAH5*�n$�������w���,�=�@���� �,�Jz�ZII�fsP� �r�I]����>��:�Y1��*�i) ���X|��RU�����$���SHÜ��L��I�s�i ���^��WN�y<�r��t]{��D����'|#�H����i ���4�XH/9P4j�)�9ˆ�
A@�(���Yy�=�U7���"�*�������>H,>RyE��B�%2�r�Z���?��W�k]<Wܷ���9����!EP�- ��_ܜ=��������L=�\4ρ��
!��I���\��i ��)�9ˆ�
A@���I#�H�� ��d���g�eB�t���)�}�$����={��~�&��|נ~@��ZAH,��O�P-$��·�j$)���hB�%FS�T@�_/��ϸ��o/��e�Nƥ��U.ыnj���4L�٣���\-��עũWY`�U�c��V���d�Ϟ�݁�N�.1�����;���;��C[kT�h�¶���7k��V�]<�B���q,��n���-�WO=�E�K7n�,�:ks`�v@ok�<��7U��Z�����ݝ��?��}��5�Mj�g��jGFd썵gu�|�lw</Ϛ��M+���]�;h�2"�ZY]���isrog������X�鳪�0j�4fժ����m��}cv���b#Q��L�������b ͋J���#z��	9o=��D�����õ#E�Me8?���Ͼ�� �?�T{E������P) ��0�r�|�I
C��I?	��y�t;�u^��|n1��ZAIY�����롌=Ϯd��H(s,�A`i���v�h� ��s��
A@�(��$P�O+��
Aa��O����uW�aĂì)yE���Y)���p(�$�{�!N�
�G���� 8��R*��QiR�RAk��@���@��.ek���G�{��H(�- ��������@�0�=p�AH(I�Y����i ��\
H)�9ˆ���9���s��#�W�>����'$�|��#��,�d�ջ�HhII�s9�|�X|9�-&����C)�r�R���Ü��I!|�;��_]w��s���ZA�D) �?^j$�0���L���
�9F�o3��{���n_����~�$�r�RAI�
a���L�2�
�o_����??h�o�Q���\��D�Ý��I�`R9E��
H,���W.!���Xs��i ��aH����k�˩���\��'����W�Q _�틍܍��WX��'�9���)
��E�B�]��$ЁL9�\4ϙ) �PC��I��a���}����*bI�	��;�T��]��1%��O!��	�\�]3�b�tI�?_�ZAH,3|�i ��=f�
AH/+��� ��.HW�ݹ����|�=�g�� �#�H�,��9^��r�����~��
H)����>H)ޢ�m
H,��y\�����Ü��I!�P�G����&a��ؘ�;�<���"�o<��0���G(c}+%�w��g(��q�_:ON�=�SX+P�h+�;��������BI%޿�) ��@��.g�%$*!��Q���Fۥ�6�U�C�_}+���>�@q�">����.d�e$
v�$������3���fAH?��
A@�(��$Td�+���II�9ˆ��R9E���R������ޯ�����e{�Y��?p�\�����r����R
�9�ZAH)���RAH,9�\4ͲRAB�r�$�) ��Xj- ���=����^0��\4�R
ឳI�����p4]Rs�$���Ͻ�߫~���٧^��7E��
H,�J}[�����X8��t�����e>����R
n�I�B�%2�W� h�I�3�?$�U�Qi �G/��I4 Ss�1�w�o5?V~��
C>�I��y��w����s��h��Ă��\
H)<Ssw2|2�
{f�CI�r�j肐h�s��|�_��wU�_~�?��߽�Ď�եic�@˒*j�30��l�`"��o8.ڒ���'�I�zD
H,�Js.�(i%$��4�R
9E���^r���7�.5�u�*�Q��|	�S�#�+{�+:���勤��R��5�
AMD
a���L�2RAB��(�Aa��^r�4
Aa�rᤂ�P<f�w���^�
AH.~����
A��������=�����ގsYN��n�O RAeFJz���RAaG9�C䂐P9�-'t��������_��Ad�)��(�߹p�AH(�- �RAh�5�
AH,9�\4�R�`��H������\��zg��|�+���G0I��$whi{*��m�+Ǌ�h�V���b�X�����CG={(w���j�C�2"U@�O�N���HI߹�����g��>�v���Ă�wa�RAIHSsw2|�H(;�4�Xi ���D�R��r��A~��Qi��I�e�=�{ܓ���) ���j$)=E���R�]�P'�<�h�ގ�UYJ8x��?
x�G��@s(���!I׳��������ހ���L9�\4φJH(P�yF�0���.�PaI%D)�9ˆ�>I���I���Ay˸so�������W�n�� ���{�|(��5�����w�;�/%����- �y��n���JH,9�\4�X|9�-&�) �P�9�| ~j�)����D���CIB�ǚ{d�<y��(�BOc��u�a#%�*�Ի�M&��H,/�����R
�E���]{�� ��
a�r�|2RAB�9�4�Xjo5��9��m��>߾G^�$�.�)&���j��w]�p�\4��RA@���$��_r�� �
�9ˇ�~yʴG� o��j;�z#�ԷiR��?�-٫W����fv*�nx�/���-��7�n�#G���G�־�����躮]�s�%��g�|���n�f�x�}��IIZ&J$�cڷ�(t����q	��VA ��޴��`��M���A�W�G��=a�{#��|R��ݛ�u��k{(����Nk5�Vq�(:و�K*)S5��k��ҍ9�Ҷ�s[�dM)0�o�=��	z��7ڱ�}�ʿ�%��۟���P�3%�|g`[r�p��y�y��X-�}`� ��� ��"�k�W��t��R�_�
(�C.��έn��/2=�+i筴)X��.�o�����������?܉�ݽ��]��]r�^�x���P���B;b\�A�� 6��n��9Rsh�xT袀�5��6�w�	��	�����U�{�DIY�v��N�~=:ł� ��D�ŀd���J����^�'����v�3�kE��`��@I�P�IK�+6�J���\q��:�:R?����y�u��4�&�ލ �k`@���6�<�0`<�|A��I.�J�"H�^i����B��uIӜ����&�vW�?zj�GuD����,o	�j-xL�x�!��_��8s~�н��^���-�jm�^��'o��J�܇J;�T�O��#R�3{Y��ɚWf�N6m�8��������?{%Щs��K��W؋�v��nj�unj�7=����Lc�����vn��K�6�92q�GpD��mk	�ur��V��9���'Y*��i���fkf��J[	�n+c��{^��f��z�L��mu�ď��.u�����pHr�J�.ϡ�u��&^Eź틸�.�����d��nMÜ�0i���$��y�u������Ɉ:�W(�@������ZL�Xm��Ylv쐬	��T��B		>����܀y?7x�/Ob[ûOg��vmh�<,\#���(���!�|�����D�IH�$V�L�>����9�o�
�Ckv3n�o<gCI�5>�o��� N���!�%���Dn�u�D���m[Д�"��m��bw.ma��J�ʍ����jA����܉�DQQYOc5!��)�wc�p5�%X3<gp������X?�xA�^�q��ϳ�۪�4D"J�$__� $����g�_���X����=��W��9{��~�$�oŸ�m�͏F���!�I$JJ$�l�;��7&�.���=����v.ɦ�-�v�����8Cq���Ԑ~m=J��o'�j�a+Gex+�/j��Vˑڲ�;���Y��%"'
��W��O|Z����*<�.�˼;'"�����S�
��R��5�m,�9���89��)fX{������ˋ��3�K�5}���5��t~��r���B@�g���H�F�!��K�{buLVQ�[� ���s "�^����jͽP��_k�$$A�|~�XӜG������v�JOr7�	j0r�k�<��$��� �%/��X��B��E`��9�Ϩx�:�r�A��쪹;q{*o������}ھ�0���{�~	���Ϭ_�J@���Ib�2T�����nj�K�qz��x�^G;��=����N�����Ekt�4�x�<��%|���,�ZKT�m ��/I����w[x� X���3�{�n��-H�#�q���"Ef�k�����7y��<�B!�i�逪���sa A!���� ��L�A:
�u��M-��՟~�Az�*"[�Ŵ��g�l甂�Aphia����������:@A�
 �,Y��%ff�}�	�]��Y^�J��Y�W+���!(�B���Zf�0��ʯd�����R��W�X��D���]��޽�J��|��/|���խ��8��+;��?`�6�_��H��$A�!������6/�����,_��{�=���6�����RvTsob�:�X<�����C�@�"d���A"樟v�8E�A�����{ْ��	��o� ��}NA�K����Q������1cZ�0�u�65+��9��#���`��qIv�k�C;%	7����'��!=�X�%|�"J_s�/Ys�U?ە���z={p\�{+�P�'v���A�G������S��gw���_�dH�=�__�̵�i�*���o��俤�w����+�o�541�(�G2�̽�1�*��ُ}Ҫ�fwfK�M��|�3ڬ�ܾ`_I�d�=�k�L�<���h IK��z���)�ۭ����������9�qU�eV�yq=ǗÁ7qLk/4A-�om�fm�x�Eʤ4�n}Y�TjZ<om��[��*��r�bW�Gf�*�N�;?H ��<�7zD;�,fe�.f\�D�K���k������z�{�"�
���i�l"����}���+Dm���z�V�fa�ne��P(M�=&�����um�.x�=k,g]����&����{�bBX�m��|�	�ʈM�f�S:(�g���kx�����|�@����%� �_"�5B�����V��eG�����zw���k������2Dx����sH�� ~�  �}bD�D�2Kߪ�G}^�/|��S�[���^ �7ԁ9,_�JD����m�h�{uT|�/( vr��B��j��gz�Jᄧ�o�@�=���%��+pZa�~ؗ���� �)�Ń%fjS���!u/�z�n�=�k|Mv����A{A�P_"��3=*tY�C� ��k��=gj����_Z��j��ϯ��]5����c���M�f�Ī�1K�ķ�:�����0�"��]8૱ک'���5ʫ�J����)���[�,&�����t"�i,on1�uϲ�v�H��ʭ�*�	b�]�Rg�L��L������4�榅V�t�r���Xkj⾭��ԋ��;�U�F�3nv#Z�f�;�p���$CU����&�s�oVG��)��k3qe�f����t�:�+\P.���'9�r�hn�����4p�p���y�2װ�EI=7�J��W��t����\Cr�,-u��GWR^mY�d��Ɔ�Y�4��M��}��0��~�kw�RG��:;�k]yZ6��E��ֵ_8��G�wp�Cˮ��h@�X�e;��t�.��^-�2���\�G {�;gK�7F�.ܓ��/�kId˅��>�$�.�P�򣒍��h�;����@�)me��q��������[���B�eW2M��8�N�Xq�/���v
��I*�.�ݳ'j�����J5�M�²�77wN�ٷϺ�oS�B-�(����Nt�D�����o�v3�w]N�G\��3�����*���wA6��*���p7�}�&:�W	��;kb�Qq�Y����Z,f���Q6�ks�δI�5��G��eF��׼Q�˧VS��(�������]��/;�&hH�NN<zV�q>ɻ�U�̭��{��9�����ٲ�7�CQ�뚝��,� ���R;��b�Y�s�_q��\�:�9U%T�u��q�΢���j�錦n�n����/sVs�|`΋���Υ�ӧ[;ٜ�g	��U2�*UB�i�R����1�nn�۔�ws�L��\��4DQ�P�$��wjwF��n��uݷ9n9�rs��U�wn.�	δsc�T���ch����w+�ݸ��4�ۖH�Ü$Yr��e�6���9�\��,�-t�s�v
���:���W. .W'\mȈ���\�u�\�r�s]�9��݃%t�,DG't+��"����7w)�6�ws��cE�E��p���b64s+��wv��� ��v�;�L�L����n�ܹ�������h��v���ws�]!4hws2�0h�����(�G1��w\�Σsr+� ;�߬s�pu��z8y�c]c�z9��Z<Y���O���轺���n�Q�]D�ޢl�\�
JE[�u��uK�2�)�g۱R��j����-�ǫ9�Ѻv��f\�Ŷ�y%�E���ts�t�����mq����[��8|��t�b����u�ԙ����]%�%����T�b��,m.�.�%ӯ%J𛛍��5R:3[1X�H�HWYf�)d��h�n����u�0��L���.�	�&99���b��+���M�=Q��8��rs��m;��8�u�E=�q��=\z��L�r7n5��"��ۢ��ϧ폹�����ڱll][ZFm
�sڂ��]iv�vx���6�/n6jB�=��8Ƙ�e�.wb2�r��0	V�q�E��f�jH�V��׃-'Xy,󻡦&��o�F�V�.s��-x7Q����ѹ 47����\�g�q��=��}�ع¦;8{b�:.Ø M숉�nVֈ�oC;���s�x�����f���n�
7��GM�Iq����թz��s�K�����ꎑ��f�*�J�J��+u#��E%�8WEMW�q��^u�m���/=&�g\t���Ls��'a��p�[�:3sfܖcĻ7cj<ǘj�i@�Zlt�Z��^}�;e��ŗ��:►S�����t�H����.�`�E4�YJ���%���Vz�ͫ�΍^HQ{�^vËG6��P�'� ��ʼ`�g�����W].�1m��ܫ��ٝ�wd�t���{{JQ�����k�HJN3��͠e6�����6��\�U�X�ǯ&d�y�s�6'���w=3����e��v6+��p�1kuI�DO�2�؞7O��k��_}�z��w����6���aNN�p!�aD��-=.�{�ۋ�r�-��Ph}�ТXˋ�F��smliy�W\i�q�\��2c���N�lI�c��-��u�gYxt��*�HͱaVl�'isH���7���u�Wc:�6�_�$�f^�4��.��֣cb�h��1���T0p�=������`_WY����%�f���u]�A�l�[2���>�:�ܦ�uU<6ā�[�IL
{ls�וΰe����ls�:�3ٶ��v���\��)�4�&�t�BfK�׋�9^-��SZ�UVI��-n����L����׃�.=B���6S:-5�g\% ! �}I�C׫~�~/�O�\#Gp�v���r�j���tvR��.�=M��rR$�\L���>�RF���|�mȑoZ�Y�pگq[��ί�۰�yA2���X��p� ���߄��n ��md{T�/��/�}��:�ݿCZ(�g��/|��ً���ֺؗ1�:�s���'�}�_7![r$�"�يY�&���Cn���<�W3�7=����{� d��+�$COUeyڿj���~֗�6�H������j�U�UVF�@���`���j~^wa@!� Cng��"	n-�G"��q�"`7�;'je�k>�7�^�~�1��D�� ���-����ڱh���f���:�<��l9M9\a�C�X�Sc�UP�3�G� fB<�$�Hn��̛Ot��U���`�s�^*o-��P�|��G��$V����u�w�Q��5��-�"��l���}������\5��������fp�ei��ߺeV���i|�ܩW:����w�2����� {����x��=�#wp{g�,�U�W� o��"d��G(xU
��7 �t�{������/�	���k����y�׾�o�~����w �"����XJ@���8��y��A�n_�+~ �d���x�����K«��A��=���1������<1P5x�r�+�d�Ȓ����v睫W����_p��p�_ZX�W�^ ����?9/�+@ �(b*�G{�9ۤ�.���un��(L�]nB*���t�mWH�H�$$H��`;���ڲ�~�޳�7�5�[�����D��&�V�F�P?܉ � 3��VN�����A��R?C�}�WZޞ��Q����s��{A|AW�2D�~|\����,�������e��y�E�/"j��t�Nf�R��d*���.@��mo|i�@�ݩb��i�Y�^v�p�7su�Cj��/fv�ne�{����ﺲ`v�����c_m~����|C�JD(�$c̪v̐�Έ���4�ީB�����۾߾�lq~��U� �����\+p"j�#_X���W�6вͯ`;.mEU:���c:Wٺ�%^��%�q4���A5pq�/�mH!�fr���V��
`OĘ�C�f��qژ��b�I�<�	ٵ~��-�}�ϧ*v7~��{jA��.���nD���W�sUX59��E���I��{�'��>@�
"H������r�$�6��H���]r|�W��1>�E����>���;�@�b��|(B��X�������Y҈?6�H-���e�{J��Ȕm����UZ<:Z[C\�A�@ %q"�A !�(K�]�Ӕ�d�-Y- �P��m�כ�+ّ�0�i�J�7��O��u{�Waə�jU}Dӷ-�:nV�2��iv�"�Y��t�����J���Z&���s{���J�k؟ok=�Q��1zڿPz�� }�Zx8)H����`�(/�&J�N�ٺ&v���e�r�S��-^��7�^�~:����G�����o��}�Z9�'���+��	�S��k4��	����br'A6u׎�-���rY�����
��z���H�#��J@�D�����v��b>}Vk(k�K�ۭ�{� ף��^���m�oW��k>�l�ȩښ4�����zswE^�m�i�Jr>�=�� �����\�N��E� T E�H�K�A��H��0�:��J1{�o<�u��r��h��O�����&�X�%}����K���c��l��2R �C��ި�w�o�օe�rP^�������`����4�"��X �"�ܗP��&�D�bǴ���|}�lL�.���s���K�J�AIX����q�T��x�V	�KӃב��X��/k$˭�֯*o-P�_A�˼:��������Ke�u��h�]�lEOj��$f?�|>s�����A�%��$,MH7i��j��M!�2�ob��8���m�M`��)-����4Kz��Q�E��5E5��ZvNn�0q���`�������ɣ�8���{+����͎ tel��ktA�PA��;�2.���XujZ08Ә��;Tݻ5�I�K�ܝF���]�v!�s�e�%��m�ٶ��ҍ;@�~�<��iFb�ێ���+BA>�6�����ȕ��i�a��5e�pg�K��	̀�mI���b0��a���F��P�����n���#��!�"An>��>S���5&+u��+~ ?R�o��:n��15������������j�8W�d:�4D�����+
�	_�K��r�y厷}���>ܽ�{U���}^��F� AK�J�	W�MKǓ~П�q��#���$A�^�){�Ҫ_�ѯ�� A~���"��d!�Sۉ|C�fJ@���IH�$�,�^����f�E D�,ױ�}���#��P.މ�@@�s#��� ��תEV���u��|��e#��{h1vыQ���z��۝Ů���s:$�� ~:��z ��W�Ib����}��V&c�{�-�bn,G�58=U��س�Wȉ+�"��#����̿�S(>�Gav]Y]�r̤Ŝ��]u��s7q�ïO�]+XTõ��sJλU-Zzx�-Qy\�*��7J�y7^q�|���p-ڟ�?g!;+�
�yފ���k���%�U�@� ��F�]����e���R N�Ib�J_$�]��rϷx���ڝ���Z�j��nz�m ��A"�����=z����v)��~�/��X|z��vJ�Wr����^ ��@�<3څA��5�����D6�H%�Kpm�U�1e�^�����l���֡����	~�`�=�"!���!�}˯������u�gS\��rm�iz��Ãh{]�;lMnι
�6,� �smF��|��~>�#���% &w��;}�R����������r"�~�)��:�A ��2Ed ��^��eܘ4g|~�,XE�O�ʲ���ngW�<P �,X2U�����ۘ,���;l}�}*��}r ������=捅��#�͓���q��͝���ݔ�V��˾|.�&n����1[뼯���MQ��� ��UU�ז��}c��{�$n@���nD��"0�en�m=��LnŃ% A0·��[��<��v��������i�͆�6W+�x���"��"�A���麋�9ҭ��R7���X�b*f�b�3����9�% ~���J��S�)���#B�ՓX��V�U�3�k�e����뜙E��b1�����>��2|��m��6��躪[u�8��}�@[��X�bV_V�9D<~�!��D?w۹a�*��:�|~g��z]�G�ՃW��_�h"�� d�K�u�֏ƿYq1˔1���L�.&8�rƽ�K2jln,�z�EL��O��� ���K��~�!��v<Цvn��UAF���pӾ���1y߮�Q��o��ڬ���bKtk�z��v���;�U�!]W�	mUG[�W\���jT��5���T��//���P��5ؕ��4���ѥ�V�<���=)���LB�����?_ �9�"Kp�����[��(��k��?R�/[�~ܯb:����!��� ���+ ��즕�9��F�tRZ� ]q��S�C�,l�\�wf� ��s����o��1�UIm�{��}��&z˃3.�32D�w����tET��3ꬍ#5�cܷ�؛\�!`Υ��$���i��"��Z��j��=�����N�t}O��
��? A~����#��(מ��L���M�R��$�����D�U��������W�u��73�-�'h>�	{AA�A"�D�?H�??*���U���U���u~|�����/����o{�m��f�3��Aԁ�����ݍ�8������F�D6�A-�@A���!O���#��l{}xE�H,��S���N����Ё�T�A���|D��y�{x���{��A���v�g2a���Kؼj������4 MV]4��Л�gP��ė]�9�kR�ܥ�-�y/�:)����woU�;�qR�9�����>��>��R�f���{�{�FG��c2��7l��w39��e4#��&��dCa����]����A����Ϩ]g�v�͢�Mz�b݋7+C�p��ݠ�e�7rm�!l�\�)�uj��N�Cs��Nʻ�U��l����\Xw/:mh�.��q�i���v������Ro&����GA�6����U��@��mЬGS��W�����@.�8��]r.�㵛�����\�3�v��[�ASvy:�eG߈���{vD��7
�u9���;�W������s�h!W�����wW����n����ԟ�$ף}z������u�|�o������Y������@��۟������U�fn~�N� �p2E`�+��[�N�cO�ی��|��x�6�D��e�@�u�~ �h/��������{�6��[;�\|��H���@�%'��oo�<�^������g^�����f��A�G���RA������%Gѱ�j�~�.D�}�������__Y�����7�~r_�V�A��)-j@2�d碪"�Wt�U��F�v�MҎ���`�<{��M䷿Y���."9E�f^�&e�>��w�}�G�*�/�d���|�=W��T��Bwv[;�q���N�#2�M�����>��U�WR�����ݓ���w���A�P\�6JC4RҤ����E�T/�{j�%���]���i�e��T|�'�SQW���S(݌_�����̏�#z���-��}����q;A���	�AL��$W닧�!Z�k���y}%�+�$��;�`�W���o�߻_����oo��$o�\�,�H�% D�ń�1@;����K���Hn����֧D�e����)F�3Y{
�{ừ�y"An��nD�nߝ���m{��^�yo�=�v2������^���H���}��g�y�oѿ��K��n6�&��Cl'���nN�%�u͸z`�؎���v�����C���ͥ�m	���Y��`�<�'�5��y���&��*b@ �������Y_ۙ�A|A�d\���f^��/�����
����謃La��3 "~����V�*��-L����ӥ Cm2R�a�q�G�Cc\�)��c'����Ե&`�z���o����F��`��[*���̐t3[S%w��6�pGH(�����U�V����N2�ꘂ%��ٚUg�࠷�����Y���շ�k�m�W���Nvt�ug0��F�m�7>��js����Z���Wr�U��������z�at�tL��ULYڝɝ��M	���͕ەw�Q%\��Zx饽J^��A9cY����:�%�+oz���rb���=WJ���E꿷;ۘ]o<�ݎpi�R�f����ζq-;��bn�T��)�W�7�}Ɔ_wDe��{��/��2vWw��IUV��ml=խ�z�p�r�-���`�e�K��75WF3���%����k����N�ۣ�k�YSE�ͱd�º��Y�U��卬��*�P�	�������j�DUBn��f�5F障�U�������C.;e�Ui_%x0ՋX������A�64]���+��Њ];#��/{���;��Y��h�{\�^��ٚ�F�,�:���ٻu���]=��wgf�u��"��:�)��v�:4
��h�R����0��YV��;�_ق�\,<#�՝:�x�,d7��,-�pm��ac�ԕs;���`�6^)�m�̬����87�5܁[pt�]�O���2���f��ӏ8z�ǵ[k�Ujϗ�s��>��U�$:�q8��*1��ʾn���(0��v�j�`�wڟu�Y\�pU�ྺX�e�.�vLՉ�ai9MϫyjT/0�5k���/�:�!��}a|���meW�ڜ���@��߯�Eˑ\�4��Ú�t��FR��v�sF$����C�W.��sswuЈɡ5�ur�Dئj%wk���6��:�dú�dI��k4D�f�hĕ�wv��T��e0�s����65���"J��3��	&e$h���)J
� ����!0H�:*��HD)`�h��X�)s�Ra��"W.bis�]�hܺ� �)�\���HI3J� 	�1�vw&n\�"	��)�"ȹ�Q�RۙΝ�e
%	6dN�$���.ƺw;�{t�y�����/h��!"���O+�p���W��={��!�!_I��}3����}:��ίN���c�3��X�<lL̳C�E�eb\s2�v��o�K���m7̃�Q_�u���sG��_6�Ҭ��^A����|u��\7V��\�U�c-�a���"�����j�.�V�Jُ׽����߻����%-���<�{t�y����^����Ї����d�Jd���ɵʷ��Ѐ��/��b�c}������,��u}�7Ԉ#d�`+C�K=~}�]t�s]-j���b���?IA$W��7�D\�5P�#"s|*kC��謃��~@���� �;�@�"_I�V�5�ܵ�^u��;*�����D$���;齛�hŏ8����,���vu�T�W��U�c� �7���z�kGp;yl��,�]���9f1�:�������<����p�]�;�y�M����q��*�u�=�NYf��~ �ڣ��n�v��r�s2�̲ٙW��L�d������,w����gwU�|����� {a�А[��!�U8l$��l�y��f&�&M� �tn��D����:vq(걼N��gM����Z���z�~y�@��Ąۀ�m���j�誧�e9�Yo�Cz���U��k#�~�K�$�`�_"$��s����^.�x*��T���D=)o{��of��1c�'(=���� Π�2E��4h;uuJ���A�����"�K�$��]6���媶��v���X��K:�:����dCA���)$�
�ot�:���z�����h"甐~m*7٦�����Ed���}{��i��;�i|C�`�H�D��X�%ooG��Ū_��#]z7�~~��`ś�NP{�	{A|Au}$ZA��
�m֋�����^hWu��N���X�zc�g�f%;�zZ�d�<S���}��aV3-�בn�\�t������:�9���{i�.�5Ul�X�t4䌊Avt�)�g���<�fѼ�-�S=�FV:�*-�bV�m4F�����Z UGc�+��y�W,�����rg��-�q[�gI�g��0v��GMEQ�m�I���.����#�"Ԛa&հ��;Me�[W6�9N�p+��x�n{U;�/'-��_�|��nՎ���hW����K��\P�5:��O?_�l2�4К�v���Bh��`�a�� ��w���u���	1sz�����?���<�B���_6БyWsٵ��ʲ1��5��g$ț���yT�s�g���$��~A�� l$��9WLƜ���2 0�RAq*3u�T��%z+ ��.>�R�A�A|~oӍd���7w~�y}UA"u"$��+H?%	�Xu��M�a=�W�ٽ�1f���X ��� ���H��"�I��%�v�IF��U�#���D�Ib�}������:�#���7Ԉ�.��->��=)|AwW�M�A����d���^N�8����*�D��/'z���Σlq���/گ���/��/����Ő���М���n����������@�P9ͺS��yte3h����E�Ӧ�R��>����i����_�1���S��{�hś��x�Фm$�n�������D����o�P޿x;'�IIv@p`���m1��x��l����3��e����9l.앬��wf:�	���s��%י�*{����8�8�㛲/f�{6[��8�B���	��|�hOŸ�3���j"���`��7��ѡ�;E��X��e�fY�����ã��gMM�9y:U:��X�=(_�������D��ʱ4�����͟�x���,��[��wh�{�C�@����Q����da��d{� D1P "�A�~��2����:ŷ������r��YJ��|Fz�d�`�K�"J|/�/wǪ�)u�	)��ka��ףB��^"�SQ^���6�s�-���.�ɕ���	d����k�7Y��=���Y��Ё�sJ*F�*�O��� ~�X�%|$���/���gef��2�4X4�H��=��wS���*&��D=�/h A��H����x�o�_�ի��^)��7K��
�D���$�[�S]�:��e�W��zdEyXkjg�7J�&6bQ�3��x#uk0��-jV�ko�����Wu(<׺�0���ik^�)%�b�����SwY��s29P��q��������%"$�`�q�FWd��@@�b�Ch wۡ���QZ+ ���M<=3��#�0�0wP���ۺ��d�$IH�$�,�X;��M�jڠ~"*ۚ��n�T�N$_�� ��|;�g�H����1�/��Z�捥�����˪�2&�����]ɸJZ�$�:���5WWuF�}J��w�}҆��|D�ŋݶ�6q��Y�3
}���cBN{v��V�u��C�Ո��V����E���/���o\	:�O�����t54�c�+h�>���ߍ�_����F�:݋��� �:�Ib�2R$��/"���ѷQ�QR�wW�eLa5���6����O�"D�J�k���s�n�|#y��J�H���y=���s�]����3ԁ��j߹����q]3Z�'R��r��C���ߴH~W�	����յ[�q1s���|0eR�����׽�k�@q�]W���ڵ����|�X�^���F�"s ��q�muz�ü7��=�;���M���{2��t��__�~�|�2K	7VL���y�?���bՇD��]���iuU�C��۶���.e�-�4yJُw��}����C�+$IK�3�xgye���NP�=a���
�Ҩh{AV"D?H�@�d���7��u\������A��7�N�6�����i�>WnD��#b�Uz�;��D'��� �� A �ڰAE��[��a��1{�綠^W����2���?^��(���s3,��U���Yj��Iź@~�;}��%y�p��;�b�DA�2OX&mY���Ezu-p0�)��3P_�H�_Hq~��p�nxh>���ϳ�������<-ʗuv��A#=_&��%i�$���VxU��
���]��n#.rK2�o�q��E�%٢��[�ޒ�+ȕͪ��L�j�էkv�fe��7n�Q}�!���^�X����q��0����i0�E�L�Jӹ����x(<h:��������6�؋I��0�vM6G��*]3ƺfx��(���Ӭ�Q���U�::�`���X���K��4�d�k�T[3H�R��MP���8���[�s�Z^:�q�=�nu���q�2/(�!!s�l��;	���JՍjF:S^Iʭ^�1��6�f�}�:�Ɏ�V�k��V3M.��:�����5�Şk^�iNl��48�
�d��2��9��n�F]�Ave����[7�[����e�v�灓}�2�w�`�������Ň�xK���- ����mȒ� A!���x�w�rƜ��}H�җ��O�^5����(\����AOu�%I�Ϸ�]m ���/��}%?H��D5K|x� ��N2p��.���x�>#=H��,�HARI�����A	yA|r�I�u�p����D�P>������q��bgO�~�_/�w_�V�AIH�$�fJ5�����lB�Lz1��cb)N��	o~�K�A2�_Kk����-լ�l Ϙ%T��`��I���vl��{m�Q�q��ˬÿ�Y2Qg�$�͒����m}{���_܉����Od�R�������|�n�g�3�ŗԈ&Q��~-�@��������n类�*���ʃyp���wc��[J��a͕]=�V]��p{9`n���U]4EHn�Tٺ8�%P��|�YI~�#�=S�w �u�p�����k(b������"!�鞯�m����Q�jя^6��f��W�8���w4���v�s<$���!�~DA�g�١�~�ӏ�̽#&e�M��n�r�v��̉�}�"8�W��$�:��9���dד�����A:P{{f�������uq��i���2��!|�]S`��cK�{Y���X�*����f9С����e���,33S��|7��O����ı�������aGam5۵�,<���n�e��ģ���o�z�!=�
��"An���{����Q:�c�=�A�LQP+�آ�� ��"g�����Y�z*l0D�~��<5�xs7�֣^Nf&k#~ �:Q���+��{���:�A�J �Iv=���BH��� �Iؾ�\����;∮iȯ.Ժs7*X\y���	͋�U�7}���&Խ�Hb����bZ�#���k7����t��r��pT�Ws�*�~cy�i�yc���5���w�סe�ffY�s*��}�w�;탶}�p�.�D���,���Dz��1+C'�=/���fe�Ѹy�ȳ�Ղ� D0�d��D2�.\�f�w\r}�����s�"�wT������� �/�%/�?a��>�-Z=�`(��vA$F�hJUK{f4!^���gi��1�kHivL���z_�C�~X�!��m����GwXp������
b����E����RS���"8��|D�ř)~0 �Qk�ذ�cc�א��8@�p��y�)��T�O�:{���@!�� d��ds��h��o�/��h AתA6������������z�{���\~���N�����Rr���H��"H�>�����f>`x� ��G3Xnw޼c�3��M��j���VS�U��V��ub�F��k�w��g,��12��Φ֛�C��Y��o=�t����`�Ye^T�����Z
��������B]�|Mf��\���i̩bfT�33S]X�;w�Nd@�+Оq^��*aN�d�	��X ͠��P_"�D���ߟ�o>e����w����<u�4���>��O��Y��ӗ]�R���5h�n5����=���k����ʹ$k�	���Q4�R���(�-�c�p��sa!�DI�d��(Ep��f���k���"�A%�oO�����~�`��D�M��i?oۺ��W� ����d�A��*��/X�mQ�+;��VWe�'hL�mA��PFH��$_	 N�����V)�A|~� ۑ:��B{��J�j%L�G���D���ŻC֋�e�ɾ���K�$�,��@�_I��k3ڼ��z��l�����f�Ϯy|���tA|~��RK>��G�]�ۮsOW���N}�0���x����8:���6�rf!o;/:�jS�5C*S⯕.�qqh�Ǌ�����}�E�]��z��XŊG꾼�mnd�cp�L�CU_=J�����n�;�n�E�!_r�2���U��
�Q���vS�rk�p)�������U"�l1*��j�uI��p�hf�<4�<�-��}����r�k8��|�W�]��B8���0�Ǭ����_Zگ��u��.�\����Ќ����`��r��:�i9��-WaU`҉�Ӷ�eJk��17�E�^ڃ���әA�ra��fs�]���U}3:��*�[­=�T�$�6n�㵭�i)�ogNJ���(f�j�c`����vd�h�C���Gw�n�UF����+!$�)-w8=.&�r2{OC����WEZ�٢-����K��]��*��Ro��y[�7�U��v�h�V��Jf�i����כ�{WW(�W���*\��˘��U�����6V��]��܍*�J"U-�%e_[ɚgU��y�3�ۨ��pY�r��]��n\?�ɧD���09�X���mE}��^J��u�K6�I����R諾Yw)��{�+�2���S!�Ug�v������º�GJ]D8�**�/)�9�6���
���*曫M�h���v�x'�F�fjS�e��Nc�c�õ�v���M���b������.���[��XyV���m�ެ�j�-�&?�������l��x6�]�~G`1�:ui�k�./t��Sta���"���mZ��<�F��I�����nw.BA!wtܝpH���ewt4I$d�b!��UБS���;�I4�#��]�I���Y��#4)ݸ S��D��R]�Ȍ�v�vc	˅$��`��1�Ӻ$�0�)1��!��Wwwt)�!����4"J(�F�� AH\��ّ1��;�
�"��j
��L&a#9ЄR3'v�G:#K4\�F4X���!�t��Jh���ݢM��Mwn�ł�\	�+��Dس]�����eΓ77$M�f)�.Era3��D��ܷ.Qg\twWA�)!&@fE��sL�)H��c$$@����I�ܢ�b�/=������0��/L9ͷY�]i`��7[e/]��29��Ӷx{F�L�m�VQwK��n̙
��i���X�3�0�Z�]�{
�vG�����k��y��;��� NX�6���%�n��8%��Bb�Q��0�d��͋�Qܶ2��:nW8�8���M�Pv�`眥��^1�`�lq�v[lCT�.�]e,λ1���0����JʮPw'F��Fxyd73ڹ�zN��iuX5WW��k��e�77
���t]vX��a�z�Փ�����z6����a���֬� [���]:�g|Bg#��H�X70�/N�q�1�}C˝����i�Ja7iؐn��i���LeVnW���R�mA�\3b�/n��8Gia���s�����ɼ\�՚'�����^�'jlJS��L<��;2�' 0mg�9F6^cX�8�6�[n�������&�W]����ݻ���)v��mY�q�uV���ib��6.M�1��T�F��|��,)��r�����u���k]�>��\;���n9^.�j��s�\�zp�0mQ�.Z�N�
u��upYi� ���,s�8�S-���v.^;Kb�4 b2�nu�ݚD�m��]5�1�F��f�H�U�N��f[��:XB��G��X]�S�]��۬+���˛i	�gN�[��ܶ�f�vQGusrIM��� ���5m��X�m�e�Ya,� �+e��F8k�ݛ7X�ӓ��a4��VC0�p馆�R8���n7,v*�g������֍)�+	)bMK&�7@��8ٝ���r�6�ti��jWL"v��Y�CJ�[�)���!�b�J�l��9)���zo��ѡwn]�k%du�G�5,meu\�8f��N��(b;r\���K��*�m�݃rza
x���2�R\R�5%ڲ�C�p�n�g:X�4ŎD��ne��)��m5�:8�$�]e� ڕR�j]0���v�q�z��5�6���׮�k�:��G�y����j�/j�_in�mdzԝr̅�(Mۜ]��lb��x9�`9vn5 ��G���ld��D+[DV �Xݮd�}�'#O�qɏ1�km0�ް�ٛ*��cVW�Ǚ�-�����؛��7��Vn�c�>�A�Lbk������s��r:�5��VvucB{[[��^�gwG'�h�P:eu㷤���F�⎧bc,�cn/e�@շ�Y�t��զs�:�C�p�XV]����b���F	>��������"p��iOsvJ+UC'���H�v�겴h�p����D��>@�"�~� �r�ѩ�
�����m������oI��Q*f�7��>^nD�[�Y4!j��E�dM�;���{�,E̢��e�#�a:��O�a��c�o[��|͍�\��_�_�t����I,Y��!�u��T}���q���6�iOsvT����_����J���e�CO?/�NA�A}$V2 ��ZGNn��/���J��vL�b���{#~ �1������J߈ �+q3�J-R�ݐR����4��ug8A��;j�K\�ح�]h�N|H����J��2E`�"�����m�]��l�g�[�.����߶ւ�ˌ�n㙚49�b)�Sn�Uv���.R��F��Ea����#�j
��Dº����J�O�s�͵�.Z,�hi�]�؛��7.�ӵ�����[�n�|AgB�=	�ը�����^� �@@�s "�Ci�1�*2�C������� A~��2/�����$��W�X�Ƴ����s��Ϊ���+�C��N�d�?%"$�,��\��$�Au���� }��&���>��V6|�P ��I��^͏C�6���vD�% A"J@�"��t�n�l/���^��V��\��A~��?f@_"��?H���W���Ο=�J5u`���nv{F��-��/"�T���b��o�磅v��c�� ��^|��k�A�A|[r:�Q�{�fk"!W��i�/W����1���?J_AR"IX ( C���n�J�C�VA�A|{��=���}}��L�g�_?5d� ~�{�x7;}q����ذ\�A"z�RK�� �$��'���p]ذ��eP���X�{sM��u�s�pM�op�j�d8:z%л���1��*��Bgc��x�k�yXs����G���;A�z��@#�_I�$����⮎��:�v�<�ρ=A���m	�h��=�35�����Ҿ�ݽ�4t�-siHr�K�L�(/�q!���t���>�{�wx���.�ϔ�@��+ ��𒾒 �0r���{[�M�Ww+?]۪��=v�u�b��z.�yރ���r'nc���*��ex�n� ��_�V�@���^{���A�^��+D�R=�W�4�ά�_�E��nk2�fe��̽����ukº��~�/��X��|������5K7#�|At���b�2Wf��.8r��|����l� �A$VAqn�ǝ��g]`���f�;��f��2f�,c�ݽDNe��˸�f�e\N���ޣ8�w_X�� �_ ����k�ܜ�Uz��<��A4����F�-z�}��Y�ef�0>�X�~Ei�O��b����q{}�2��C;µ+�f��79���Va�[�꽩S(��w�+��"�Z����|sھ��͠������:�ùNv�wJ���oX�;�j�Ox]�uU,��^ >�� �:ř+�����}���w�s���4�2�j�!-��Ah�E�Aၦ�n�m�p[�5��%��3߫����~���2A���{v+^����]P9�}�n� ��a�ɝS� ���u/�mȐq� ��b�����x���7ak�cs^�Ԥbk�}�l�W~9�-�4�0�)�H#�R��S�6�?I_)%���l�o��^픛���T�oz���Ԉ2u�J@H��D���ʳ��ݪ���ӗ��h#;�ʭ�5�{��]Pϓ���j�<^�[�G6f�O
c���|�rŃ% A �)�Kd�Y�u�UwB�X!�-�&�no���Q���� "���-IA���̭ܿ깙)�uu��Q����ex��~V�f�����]_����U�]����m�'��ݺ�K*𬵕B���#T�.�Ձr�����߀��뉺ڒ��az�6�Q�ƫO�)�-�Xo�K� 5yF��jlML#�(�CJ�5&��jU�73�۲���փ�ҝf�^�P���b��f,Ir�Y�`K��Yc���;��gm�D�#�B넫Vz�u�4�r�	[���psu���d�;k��o%р�I������e.!1(�8�-jT͓�}}�-����:��Ǳ�Ke�u��v �{� ��ʣ�V��ku�֯�_ф����	��?I_ $�,g<�Wt�����Vm��K��n5����*F{�,����]��,�ʂ�W�~���u��������ML���{�d��z���;7����ذgR ����X�% &h}͵X�����I2��9A����{A|AE�����På>���f�D��N��I,_����y�e��*�8�H��<�2�P3"���yW��34���-�ŋn�Û�P�Y>~��L�ѵك�sA~�$h ~��ŷ"h�N�f��I���5�T�Q#��[! �gJ�I��]��䂊���p+f?_d8�|��|����/���{��R��Q���E�<>u�6�.��:O+ �"�I_Iv��Ň�\��Ljy��_W����`�N�H^K�V�t�Y��ݔ �Ew�>���Oa�/���e��nb[���M�w������z����,s�ނ�o4L�9R��@~�r$���P�q^��:�h#6�z܉�@D���+"�ڽN��'*^{6p�gguS��~_M�$��?H��Ib�2W��C�z;�@ �z�Y�A�%/N�������p����/h�9J��v���z������|�_O͠��M^�j阴{��01�1�����w,��%{�#}K�q%|6A�1�>���c5�SmD�ļ�t�+��Th��˺�ǳ�r�u�ʈ�F$JJdH�)�y�g�m��m����{��*vwy��ͯp�_b���&W�w/��`D�y{!�j��\CӁ�~�{=�*�ܭ����s�Oy;7�%R[oW��@76�m��'D^ҫ�<����lK˥��&���8����fM�5�{���WM+/�����W�[W�31]1�ꩣ�l�]k6�t�m��/�Y��w����Ho�a:�>��	�_^��2�7՘Ϛ��~�6y�Y2߲�ݽ�s�ؾ�D$���I�=��U`߯4p��/oY����i*�ܭ�����	"�M�ot�	�S��l�hFf��e5��b��(X����E�{�#��!*d�H��ǟw��_@��m}��|O��3 �'/'�q蕇}��1J�۽}$@I@J�5�!Y_Tc{�y9_/v���ޕ�<�
{bl�|�����;]osF��I��$_d��p{y�&+��T���~��n��n�ovy�ܛi���5u��F��1��������9y<7�]wS��A9�^��՚�W���e�F�2�y#ہ��,�Sfbjs��J�Իx$�f}��T��V������l�>�#�$��+�"�o��=�++�]�;f�-�yS�#����"�I8�{pU`����R��A1Gi�vZgc�����7M��BSh;�UqA�h}�������+S��y�77+zg�b�%�����!;��T�}#B M�<�N}m�����r�D������k�!'��f�ޑ��{��j�$�H��G���w}����<~�ٙ�q��|����裸e�U�YoO���=�P�I�±I��x���ޙ�]�^v���_9BH�� 䐿yn7�����q90��o�������JIG����ݪKDo�"���Q,���7�2�]�X���C�n� ��a����M�����W��^W�u�oI�s�z
��iD(L)2JQN^���v�<����).�q��]���ۮ��I�u���mj���w;DΧ0@��d�Z�a{1#s�5u��;T�xj`���5���erֺ8h�\�-��{%bc�,�;"ݫe�m�S^ےbX���=���(8�v*K��eY�9�c���������hL'�]46l�h���n�E�Zg��ߟߥ�2�t�����vޗ�M�\Iٰ��1�����5�$���t������?���5�^׼昍��m��\ꊍ��m{�8z�m7 6��cȜ��{:�n��u;��
���{�*C3r��x<�:r�h�m0�/�m}�m�C�����x���^����8��~�_k��(I$�{���eo�5����}%/M�O2߷b�+ٔ$�I��j^��[>�I�I�I=�޷��� �-�+W�{�iR���3�<����M����ߟo�����5��q1R m�p�ltg�����\v�ҷC%��Ƶo������,��ki7�	��B�+	���M �����T�I�}����2;_vn]��m��u�@�kɡeu��l��UU��;����෧ne�k�O_�Q؉r���7;����]���~���{Խ7ϼ~��AK�GI�@IBH��v�w���_or�H����CTH��Ov�^����ѩ?{��UH^�V��|���$�	*H���9u<^
�<���r�I:�I�W�X�&��Fz�q
wYǸ+c��$�	*I$ۇN��+�����s����T�-�1������m|{�c����~�8� �B�C��u�.���!t����X��JD�&(�"�2��M�������ow\DH�z��/@���Hڪ�w��Uj�n���6�g�(^d�$�#o��Ւ_�?{8+�r����Hsr�f��Ȁ}RD$�I�2ꕎs��!���{�ҥg�7���\*k�kQjM;e��ڹ2�;�}����mR��K�������X����D2΍߬��y���{��d�K�YŸ/�8,m-*��؞�󂄍D����*�ԅ��t�G&9*K�&����\[�+�������$\P^CuKk�SQo�ʔ�&��k�[m1,�ѐ�����[�Vu�//o������)
ɐ��s��	Z[�:�U�W�H\��;�ѥo����������;{��������k�˲�E[�k��ܷ:HJ�LZ��Wt�X�TOA����b���7}��f%�S��8<Vi1�t��ݞ޳�;���i���k�u��*��A�"f�qgS��T�h�-NNǴ��U:V���@��z2n<�8��q,�ڴ��=�F��'����[|�zr�o4��N'��j&�$X��T�|�2�K��}��Wf�X�=W����5�û�ч6{g�z!���c{�3:��	t�=U�m�6��x1��e�C�u�h��Ь[��Z��9Ъ��5⿭���Y�:���=نbz���z�̳uC���I=n�g��Q�<�kw��u�z���|�VBp��)+�n^8{�2������-�F�8�_T	����UN>Zɜ����Jw�c��}>�Z��w����)^�U�mR�ga���9m����R�;6�n�b؝z�u[|&�:�;��oU��o����5$��R�t���ں��;�:�%l=�5���v;�=���\��0&K��e�βZP�B�TBk� ���&����n���LD�d��M��r�F��0b��n\�����0b��r�$���F�d�ŗwM�JH#�k�4A��1`(� ��f4RD�D��B�4BI��r�Qi4&��� ������RH`�%]ݍ�˻���!
P���2E[2r��Y��LBId��͹\ HĤ�F�7:J
L9�A%���f��!�p.tN]ݫ��Hs�&�Ɍ%�`�.�p�m%Ed
���%��F1`�Wwb�P�4L�"���RVMwX̤�A��t�$�Eѻ����.��77 ��cT�(�Y��߳��M��R�#���5%}$@I�&R���3a��q�*H�>��~���b�r����]E�d��L�P����@k��h��7�VyR[1M�����^�n촯6���.�'���	*I�2�{x�&W�����v�lQ���)���ţ��Q2��X
�Z3qK�	�ut.��5j���6�~��"Jy������ht������Ό^���2V�ޠ=<��`�!��G7�G���_s�{Ͻ�PX��[�=��A�����Q�e!�Y�պ�Ӽ��I�I7��M�sP�c�]�)o�9��f�'�wd�*H���;OM﮻I�|��v�{ڷ^z��m	'���хז�{y��Ə�\��m��}a��6j��V�\����}NՎT+�b�ݥX���
<<�����Pt����뽙�}�=����RW�D$�A�	�Ͻ�֬��J�٣R���j��z�����$��������]=��?�I�ᴱ�nx8�k����Gl�)�����6��$�% �_���s�/�ty�'���G��Y���0iv�՞�ӗӨ	"D��p��{�'|��5��@w�L��{۷�=��M��}Ҿ�M7Hu1@KT}���n>mɩ���1��&,U����d��[�x����%	"�Ѩ��'`��-�� ;�kj|��=Y�2�T��{�V!�;zt_�d�	�����q�����lJ�3y��ڭ׻{v�2�򖆹���I��uª�I����׻��xa�"�+2��V�r�������7+�2���tf�>�����c+�^yf�i���v�����Ƭ�s�Wr���͌��e���9��x���t.Ԗ}5%���[sf�v�0�"]ezm�A���:��[KRJl�!(����[/Z��Ð�b����	��Q"�L��vF k����7m]Ӻ�Lo`�i�ո����FǶ��L�t�;:8{&q�c��M͸�uг��fY�����:�OV�nƊ��Rm�����ɺ�6v�Ϟ�غ����kU�v��j1A�ms,�F�ܪ�h�+�7E]f�Y��^kC��RW�D9���N�Ӳ^f��=���w_^\�*φ�@7�𒤈	 UN�M����˻��{,�o�W�������_}�I�j�Q�ѴM��P��}_	$�@��)�Q�~7�^��y7ڶ���T�s�?E�J� $�J��7�W�o�_wW�O>���]m�Y�{�y�����lٍ�oOt�I����=�c����=�^��Dʉ��}5�6�poL`rwEW�o���^��\՚8JhQ����:�J����S��L�T�ZPq��&~/��Y=����L�c��ڿG�wT�5�l�$�'�}Lڏ��)+喇���ͨ���{v��ZЫ�uX�-�"�/+������eU^���f�g<�O2�j鴇
P&ɨ��ې�/}���!S�(k����^zw��̵�{�x����$|�̛=X�Z�-L���_I�J�)'�q��깪��װ)������{�}�l�����9#7�R�ַu ���_�����Hk��?D%j�֔[}�܏�Ӥ�$_	$�	~	�-��,+K�u�{+l�Y�d��};�D>����2�5�I�cB%]ګ�d�6�=�ݨ��^ؘu���hЛm���f��f��_?l����cm���sr��B�9�Ϟi��1��)�Emmj�=�{�$�	"�J��zƕt�g��~W����E������t������*9݉	{�`]��u>��$� �\��zR\k��W��ף�9S�r�U9�)塝,&���X�����#׼��h�rԱ�`�b��.k�bыv��Т�������[er�ݑ{�+���B�n����,�`MFc_6Н˭�����ͅw��"��W~�����E𒾒)$�<���_f���·�j���|j�l����/��o�׽\�~�L�m0�\��1�	�ŮA�\t�=��p؂!$aL��&R1""�������|hk�G�Z�j=*1T{ͭ�X&v�o�l@���� ��}%I�E5������B� =�����O�l+���hk��2�*�}�k��m�߳|������J���"�=��t�"��$�����zяV8�1z�f#�1�8��n
ߒ�Xa�����S�%u��͗XE�v�����;��9*���@�3/t��r�/5*�.������}���=��Sٺp�*�V�p�C��n~�������Z���Փ|7�{����{���W�H���V��=�UU�tHRB���-�m�=�����h�X��f�3�&���__~��t����7fV�c�;�05V�~J�iT]y�λ�I� �c����e&���C��#Z�=�+�ݑx<���Iس�������؛��L��%���E+B����n�,zÜ{����{���f��t�FԻ�0U��/�r/��˭Ʊ�kn�!������<R6����z��{��������lS���^_b��ລ�Q�������[�/|WӨ6�luv{"�Ψ�z{4S��wF����T練6�f���gv�@З�]O2��h��/.�-l�vA�u��o\dVb7Uq��C��كt	�vj�ѳ����ڹ�l� F�n�����6�猛I4u�)Z��Ne�h����� a�p��c��V��X���\�`9'��������|�����vϝ���\B�)@ɶ�qt&�m6�m��th1���F4���Jaԥ�fˈ�K����5swS�8�v��饹hKs4�Y�gg]`��ٌ�%�R�������,�Yۮrq��%})]s�v�Gu߭�=U��+i����c@oW��������̾�ew���ؕd��ۿ.r6�m���{��:d�|��=��A�����>w���|>�����of���-�-{�u|�A��h�����­��F�v*ݑy�9��7M�� 莧�ڳ��t�o7{���s��{����{�k=��g�W�ͼn���׈��v'���k��8!���|79}��:����ՠ��]ѻ��N��tY!w@\�=�No<v���;�+��Lf����gr�n��p����X;UnȽMy���#��s ���@6݆��6��晈S5|W��m�U�\wLύ�QwVWN{��C���w�w��uV6�=��R
��0�A8ݩ�%^����ޮyǷ�]�w^�J���H���{k=Ο	�f����ΆlmpfNd��N��ޯ��h6��f��5�"���~�R����pks�ny #���h7_7f����x�읿vj��|=�\+|�6`�9��k~�����S����i|5��m��6GwRh�;���ڹ�N9��N	馂���·۱���7�z����\��7�FQ�Me�]/�-���6�N��� Cq4iZ�B�"�k���m��o��8���֠`���V��{����{`n��v�n��-���o�+�~k�K�^���;��n��]G�Vk��W�sm�Hώz`g�Az��=t�~�>�m���f�Y��F!r�]oH�33eupg��dfW�v���Ih�=�n{�Ʒ��q{��L��vT�@��ʻ�];;f��`�ގǮ��j���7�n���6���V�vN�S�X+�ϬI_+}�u��:���pks�ny
"[�͑���[n<����|��m��^�+�����v�}Pm�N�oJ͒��y_}:�m�ߋמ3}��'�(�W��V�+5eQ*��,�g	ZF)2L m0X�l���1R�J���k���w��Y��vhn�xn{z���A]���&Z�L���_�2 �7M��t��Dᘧ���Ɇ�P�f�nb�ȝN�V��}�t٫�6|�0or������M�{[����K����8��/J͒���N��@6݁Kg{�X�=��������w��S�nz�W{=Β��[�4�e�MP�|b�˻vs��-n3־�R��}�t�iHZgr�[��N���]O�h�v�mz�6v=���漝E՜��G0���;��d]����u���39J��=|0m�I9��ޫ�8;�����n�mҺw�ϲ�Ͼ3Q�]��+5��9���bݴmẓ����w2�l75�V5����\������i���6$�f�^��;ӽ�ۮO�=��>n�n������b��ǭ������g�/}��	��!]����o�˹��ׯ���/�z���A��������Os7\�j�r�{��_GA�6��y�G��xf��!n�gݦ�w\0!��%xnU��~�w1��ؽk���m�����=,՛�sWVY���}�����6�D+���s�3bn����?����@���,�2���I�3����촞�������44p.�eކ-�٦�	N�*���-ϻ�l�Iօ2��V�ʫ������ya��q�K�R)iyX����օJ�\�b��9�I32��.�N����ǑZ �tF��8�ш��sv���p�롶�Fx;.��B)����1���c�;� ���ƗT����֫^Ў���`�ʙڮ�pL�g��yI�ڼ�!csqY�*��j����S"��Q�_[Tv��m�B�e:��z��}Y�kq ��l��Yփ�ݝ}ō9�*�R!>�ø3�3��قйc�����#�\�ѾɌ�"��Uh[=]>�)v�xW�<me���㜎ba�Y���4Gh2����dc���O]����fG��v�j+l�A���
�K�T�S�X����U���k��]z���y]��cՎ�t�vl�]]&��t(,%>�C�����1�W�Y3'ur=ݭ:��n��ǊTm}��)`�޵5���x�e�]�m�Wy�f�)���j��o6f
r;�Zb"�U�\۔qUr=��`�������/7v�=�R�!L�uL���%Zq��7ݕ�����6_-���f��曭���{���!Y��o�Ѿ��ss���kɓVMs�	n�b�;�����	�﷛�s�h�Ug�g����5���}3���Y� s�༧}u3e���y�:�0�n���yϳ���ǽ�d��u�ק���~��jۿ�b��Q�F1�����d�m�!lP�.ŌDQ0 5�R&��E��t�.�@M�LB��i,G9D���'v��A����̀����"!
�A���,XJ1`4ȹr��LEcb�M��)"ţRlF�&�`�0EdѢ(�#DjI�"�`�F�����PF�EF!(-E"D�"�"�&Mc%�64kMcRY��1!�Z$�ŌQ�6#F�dɱF
�F65&�E�2Ent�P��"�c&�ƌ6MD�-��cF������1F�%�5��X��R����X����U���Lzm�V7f�#���9�p<�v�{suۤ籮w����y�{%һrI�e�����]Ό��GP<qn�LW�3(݊��ȘH%����u�-�٠��jm���ƪvrKR
�H��uъ�5�шw���=��m�`[�X���i��������!��0iHlG:�^A����;j���JZ�#�I$�ٗh�[!��@�6�p�ؼ����u�˳�+�秵�]����F���QaŹ�+��)�'m��.��ٺ8�k���:������zBۢ��\؈�W\茊��CMf-��Ge�8�.�j] "@���8�0[��7���v�n�ok�l�����ᮟ/M�b��k[�Y��:��r�jB��l.{y�!9�ֺL��P��Z��0�Z�]f���n�) ks�1-,G������
����[=8e�8��a��iT�Oi�k=��rkN�	��ۖ6���x`�9ӎn�ŵƺ��f�Wi��,4W`�U�i��f 8�n��
eռ9�� 	%1��m����ٖj��r5.f#�kr�D!7�Tn&g�98�&���\M�<��9�V�ś!U�-F��f��]Gp\{/:4�㶛:��`�ܑ�-I��)�K�9�� ���+q�9t������,1��L���0��L�{r�"�2�e͉u-qŕ�;�fdR��E�n7%�ZCh3��um��nlWR�J���m�(f�<�������p�(����iN��A�۲�u�F�%�u�&���4�\s��H�K��T��=���ĭ�lL֣m��D�u�D������m���y�qZ�%���Y�2�h��#��ܾ���ʒa�U�V�vث���:�^2��h:h,L�lg:,���3ݫ���Z{�:ۊ@�W<���ǭ��ې�{c�wtOc���"}�u��43�J����6͗�Gl���c�d�ݸ<IvB�k��p�����y��ꎖ���Zru.�֮�8�eOi��������Gp;t�Ƶ��)��Lh�"������rW F��]�N�k`&��.u�͞:б�}��{u�DT��a���B:6*�YV3_W9��GD���jA��vJ�[	��wc/��r��k/g�'�;��\�W�4n��뙸�,g�y����5��8T��uV�;�n���`����Ŷ[����5&��ay�iS?<�>�_ٰX�겐m��oV������M��N��M��T*����#�G�}�_��M�n�\�oڌ�8=>���<�ٝ��,=��6���}U���J깜z��}�@7SOv���yC�a��r��M�S��V�+�����@7A��k����o�����o�m��W{<9�F������f�1x{��}BH�n������7�8m�{���={���>��鼛��u�m6���s�*��̠=��Og�D A�l��@Nm�m]V)O2x�����	��1�&�!�o\Si��m1.%�ޑ;в𾵣q,��߾ֆ�����}���<9�~���g���Iܸ��i��M�ϛ�h�x^2]�s=2��3i'�M��B�/�r�9�/^.�B�u�9��=z/�<����C^�*z1���]��5�A�)m\�_V�����oxL��{���Vd���6�=���t����g�G6ǲ�����t}v��ug����Y>�;�8y�U��_�ݡ��m�������-8��r2�Sm�����m�������qnY�f^��_l��_7_7A�w�jw�R�w��7fN����}��#m����rb��pU��A]��q��n���絖@�<*{9:�Ǟ�wV��՟$X߫��@gy7@7C���/�5Ucݓ��j�OI��n�tmK��{wv���=�5Z-�NuT�>z>ɏ�����s�[�����/�}�A�m��ʲo�T>G}��̣6�Xi��S�SV�i��r�\����{��p;��BgVm���Vu�[!ʙ�;qo.�'WJQ8 m=�U���M�+!�X�f۶yY����w᷹�<�����o9�n����^����n�6g��w5R�)��{���pW��s��<@w�7M��t�ö���ힳo�./,�g{���$M����l�n-�v.�P�n��	U���ݘE�اty��)�b���ݼ��Nu6A:^KvW��m7_wy�}�^ۈp��𩗫��g���'��:�m��7BD���QW��s�gK��>j�*Su��7k���n�j���3�r�|3�Mh��6�W�5k�3Ԭ����ڜ�]��
=u���_6�����k��^���71}wn�����jZ=>��jw�[��� ��$��0�oMnƷr���h_bQ�<�H�Zk�5O3z��wVl����[f幘�mKo[�`.��:���/W�� �vh6_�?Q��x��_1�5���|ʙT�����u|�@7����ɕ�y"n�(]U�eU�;�m �/nm��;��ԙZۢ\�KFe5���O|_sn�k�g�V�N+S���3ۂ\�c�1	���i�=�]J;�ꤠ��>�_{���b��^ˋ�����s�t�}��c���h:�w�����t���y���q��7\�v�Sm�7_d�+=������z�z#�Ug��[Oي�o{�]}����b�7��_{�xu�tyt��5�]��yl��t��Ƹ����B:��6۳M��|q_����޾O~�]��b�y��x+�0?V�֘��<5O �K߬_[k�+�F���o]��b�nV�JHKAP���"��cvx�bu�Ԅ�#,�gV��+��h�s%����n{q��b�y6pl��md������.{!{Qmʼ���6�W��f��hS����H�Og>޶9�\�>�k&�Kq��QT���[P�Kj(��MS����������Wf(|������m�jZe��.Qqädˬ�c<5[��dK����&�5���_s���	tq�q(��]ok�t�X���Tx���uŖe.�&��{�;ϔq7_7��读�\��*f�<����y�x�}�7_���_(�D����t����kϴs���8�zfU�����o�b{ז��^>�������7A���΂�p��J�Z6�����}1u�P����Q�n�m��z�b��F���ٻ�t s��{)z�S6I����F��{�}z�n�m����מ���Y9JP5�ì���]TL�f���d���7�C�|����U"�)�"@�-�(`�u�5�+�^�Zn��4v��,�����?Wk��~��k��g�=�=�.�x�'ss��x=��>6��<�z�ʹ��u����Y,����P��@�9b���uN��e�+LWca�����HNk/X�˼����S�`�%Ռ���hn����4��NT�پzp�o��{�0UK��ݯ����Uf�������#_7A��/x�p�o^=ޯS�Y]3*�oxz�$ot��"�z��,]���|��p��=�'3�[���o����$��J#�,��H�tth6nUa�6Up����b^�(�{��k�y�����}tz�^}��_�f�ra�M�MY��b��6�]�Gt�;�����AK,л_�����n�mh����.��y���x"��ψ������W�|�6����'����g�2��/�����w���w�1�<���s�u�u^eQ�?I�C��|�@7_���I��ٺ��m�n�d�˃V
% s�_ҩ��7���A�ST���ڲ�R��c^��{����*�|�w)1WPU�^/��.5�y[Ck�ms��Y�b�rx|��Sm|��W˝�U�yӔ>m�'�����<�Xw�=t\�8�w[��%��΃m7_7_�U���P���z�%�Y������|�ߐ90�=�����T
�ٯ)��N�wn��������nZ�WjF��mvl�mU��t2rn�n�m�~S޲�r���nxw!�T�o6��Wso�s����d�`�;^y����ǹ�9u]�t���;(d������ �ٙ��t�_|���C�׻Ao|6.�%�뺛T�s���@F�m�B���;�����Pr���+_{<_CUN����t�ߵ�����]+)�~��O��+g>��"u���iG�]��U�yʛ���v0F��͝�7�c~�[��th7M�A�ݢe{3�5�gb�:O�ۘ�S�Ѿ��6���oc�,]���.���J��I;�jS�|ЛԠX�k�#[�esk�V�]������{]|�A�8y����Ֆ��M���(�3�����=�ڎ�m��|���ƾ>��/�*z�ە������5U���n�P���_��U��P������6��ر\��uu��/ǒ̼�K�Y{��24�7A���3���y�|���O/���7�{�:z��ک��ڔ�x�_��;�~M��m7wSݵ�m]]��N/{�KQ�����_IA��O�Z�^���:Ex<�}׵[T5e	�}��n�>�u
j��(&hi�V�][y��%F�VVҌۡ1��H,�ꓫ;���]YK�b�B��ڎtQ�a).�X˝n��(�MenФ%5�E�Q�[�sX���\�f���sq����뵨�zN�7A�]��ζ=�Yz��]�k�p��0j��yE[�x��<eǶ�=zu=�:����qv^�b����nb��"�v��n:�x���y]����?f�7�C;��\né+\#ۧ��&�G���'��~��]J"�љ�[�j��^�Y��w[�X�͊e�.�-F��k���'�?!�:�m��}˽1Aו�t1^���*����}��u�th�30������s������R��>�ʹ��n{��_G@7��[n=�1��u ��m��|ڥ�����O�D���K>�3[����W͵�t�vn�+��}�i�5 �A����*u��13+�P�{��y������w`�y����cJ�mj=���O����ǹ�6��n�m�Cr6j�^n�t�l�����X랂ط:�N�:녵��d��%�P�YD����n�o�Qo�{חl_|�\���Л�;��.u|�_7A����S�9.��V.���t�-�:��V�Y���N(wn����b3�­���o�ՊY⽻�Dw]�6*�r���Y��7r��y��o���O_���2�V��΀��>��2�n������������G5�ݯqtig�����.�ɹ�������_7ClU��a���ۡ�A�|�Fn-��+�=�^��^T�{���/�^&-�|=��m��`�/ys��K�sz�e��V��u�H���9~{����1lo��J9�i,����ە�is.���Ei��h�V�Uw�E
*�"�}�����~���^���j�7�����J+��x������o��V�Cޯ��|;M�N=^�5���[��^P�m��v�nO]�젥	���Ͳ+�(��b�J�*=���Y-�j��#D�v�j�r=w�㧞�5[9	��5��Wop��7��o��t�+!��o�j�������Emݴ���]i�kX)J��у-t��zm��&j�+n��Gt���y��f˫�}\�).����t���(p�m+����yU���y�Qטz"��F+T�f�Y]4�����v+^p/���]����%}:�Q�Y�������̬W֘�tr$�";D$$��nZ{ �bپ��T�n=��t:�n$ʰ�y�l��I����fւհ��D�,t��'B7�ؒ���E���l�;"������VCK�,͇�8�j�vK��q5�r�[���u_mf�J�B�.�=&��
����5����R��ܔ���;��f]	��ޞ�֬J�$^)0�$�B�]c���BM�ZD7iů\W�r];�Ň�o35q�}Zgk�U�D�Հ�R[�U�v�A�Ǐ/��Vnf�jT�ձ�,�\�詷��'�<Y}��5�m����Y�/����r��a��ܷ�hصx��[�.��3�b쫾�A��;��W�mZ�9}T2��:\���V:'9�_FkfH;Ac�Ukw$U���Y���]2cΘ�ld]���"�zHG�X^�U�מ|�vͪG��Sk!�ۙ�TX�*�UX[Jv�6"wx�l�M�����{�[��y��`ї.��31���oX�:��Xg&�٧7J�k�Ǖ�n���O�kw���v�\�;.q���^�����ep�_�n�^�p�������dP`?�R��ȉX��b��(�$��Yݹ���Q�b��2���#T$�(J$QF��Y�9�4"j5�Ě1���i6���dѣ%cN��!��X��VI*36b�b,lcL�nj�l�Qa��,�cD�h��A���& �b�b���`�"#h�u�#�ԔM��a"Q��b��0EnW,fUsW-"�3�2����h�4�I��Dh�)#@�0�P�(ؑ,h�j1�N�膠��}�s�:�����o�<�d����_�޹Ơ(wD���^�v���]��M�}�ŋ�x��x�|��
�9���m|��h�c��2���	���Wfym�������m��+���r��G�x�ʼh]q�\�R[�XŴ���Z�������ƨ�į�Ą��˴���p�����~����0��3���}�qMenu�����Ch߀�~-� ���x����ez~��`-�i���t.�76�_?G���Af �-�vڧ
�n�kT�C��� ۑ �[A;�q22��n}�7I{�ޟ�Ј܀��������zgwg۷z���_[����-� ]�-��ۘ���
���� �ݸ��el/Ȓ0E����B�0�^�7�	맕�j�P��n�ǔ��`�)�r��|���u?U)��U.���z�Ӕ���NA�^�*������	�7����k�oӐ,{v�v�{��%znf_?G����1|�}���n{�`��ڳd��ʿ�B��)-�	u�oX;����1Q�#	�Iu.m]���:9@�[=����͠����f���r�Q���;ޑ3|��c����#og�����[j~#e�/9o����}~=mM�b[ٺ�S�B�x^��y�_G�$H��F�I�1�Z{�ӫ��"$��dA�<�[~�.���+m��g�;����w�M���3F�"-� ��2�����h�����?^��|�C�z^W���jϽ����BO��ב���:�do\�?c��-� �ڟ�-��q3=�"�Z'���Mn�CYٺ�)��!S</yo���p� ���mF�xY����+�k���-�p�|������������zU�/^5�Gx*�^�"d����[|:��6^X�[Y��.���x���e��w�].}B�$ht�Tr��PtQ�1n�A��z�i�zΪ�{=��A-�JpYGiFٶ��Ypԯb9������:�R�Uȑ�Ga�ۭ6nH��.��K�W�u��7c����"�MC��m�R�vwVd��ԗvݒ%�s6f]�ك;��\q{cHG(ݕ���dT���f�.�c*K09�.�2P�Bi4	�|���>�Q�M�{mn����w:�	�\��U�q����QNh��D����B �������/���\�x�e��fS�8�G�D_���/e��KG�S��;�� ��_7Ÿ��~���6/����O� ��ߋ�V�]��!՚���ס/`/�m�^��F`e�Uxg�J�D��A6���"�Z6ph��M]1�W���˺B�t^�����G�H�[��h Cn~���t*�rz6��s���ւ#sdO�6��{u�����y6�'�q����$w���߃��7�D���~@�%2I�n'���z�V����Ã�εþ�Kw�H�
�����W/���mȟ�͡]��R�H眎�� �jQT&`����>�"�n�cӬa�S�V
�mƠ��a��*;f0��) ��[���[joǱo=���y�M���eʽ���]��{y	 �?6�6�A-�9ح�(���A�2��r�f�Ѷ�o��\v^hQ��{ڱm�Z]9�vF�����T���~��['�8Y�ݻlq�%�xE�������,��3Y-p�D�/����^����&�R}�?\��3 "�{]��6ă�T�Gy A΀��$���htI2}	[����Y~�Z� <�>�o���^�����͠�q�/�m��}�gT�A���/!Am�����7�{��h����@Dzz�}�)�޿d�= 3��H&JD"�$����u�6����h/��s�����f�C�8�A.�}9�"�|����Wi�^%U�$S���SY�3	�ul2
�/O:�0��e�]7s::C�Ǡq����|�x��kw���::�����~sQ�d`2`����<A�W������mH#=4#�����^C u��9Ѐ ����Ƿ#��։�w*�'�� Mtx���o�}�%�DK�;@��H�M�"h"s�h^z����s�;�T�	�	��~���(pY�� gnT#v������Z^<���̣����u[ר�J�"�`5�I�UV�{����w+j��l��韔�s��|A-� ������v�� �ܑ ��6�7x���L����z�=�	p��i�DW�|F�ȟ�`"� A���Am[�8�wK1}#ɬ|�O���G��։�?B���{�����p��+h���i�b��3�tn���m��ۧ�F�^�����8���x텺-<^w����}�,L���s,����'�����6T>�!���7�,��e�eK�f^�2務E�������d��W ��/ !��+��8�'=\�	ӄ=A��PbL/np���~_n�A��2 �����쵻��y��N��*���&�fH��p��o�H�R�ہtA�w��c�t������_n���Mv�Ùʇ�q�A}�${��k�H�jԭ����Q��7��)%�d{A5j��Eڲ���h�ne	���V<N`�~�^�v���]�������m���w����m����$_/���D,+��g4����<.�]V�n�"s�c#���t���������ڡ�������8�05*UH<Rp�f�Λo[k������|�=�ֵun�1K��X��2���Qne\E�jE�<����<�aUD��Q�oM��8�r� A�u��[�PM��2R#���=���4�Y?O�=C;׷ʩ����XT^����) ������\l��?X�:�Ip݀mȟ�p�?6����'k��l�B�O�د�	�2}<2���8����͠�-�"�����v�Z�r�D�Sc�"���D���U�� ~5���!��1Z�;�~7p�6�6�A-������ �o��Ω��6�2����<�>¢��p ����'/�� ��~ѷ�����X:���W��+Η�+�1�㻻�y�T���-D�wam%��l��-#{�6�cl��;��sq긅��v���Q�h��m���*�)VmK�E�e�Jc���.�7F�Sne�	W3D зSb	Z�\�"-̫��a)�R�+��Ɍhy���QwkǤ.y+G�2e@;S��
���֜�Lt����qjz�� ��V�"��ۉXD�0�=m��);l9�`n0`��{�����!{�g2��p� E�:�l����v4�TuKK���u9	������{pݪ�\3��k�����47\�g����6X�BR��S�b����}�"An��n��3�Ƨ'�,�ڬъ�|�܂#{��"E���L�X#����]Q9�~=p�?6ԋ����O?XUQ<�_W@C��$In;.7o�2�DF��z)�dw\� �D��k��(�w��;�2��������*/��A{�$ �-� �ڐCi{�i�5��2~ݏ~m�k�h��l�T��Ŝ'�q�C�[31�m�&�D�F�� 6ׁ6���[��"���O���o��y�ª����?���$H-� ��s�~9
�{}9�?��;��f3U��{D�����Y+��*ۜ�G7d]@�^�	�r� �� �O��m�w}�Y�{�=�"��p#Z�c�z:S�I}�o �=�mx��/�p"�~ѥ���5�����t�G5>^�t�,wާy�2�����}=�狭O�4ej�!�����)^�E�VD��Ɋ����8��!���e��1��GeG���� �������~�r�"�|y �9�� �s�Df@G2>_ڍꆗ������z/+�')�U��ƺ _{2D��"��!��s�}�>��Ƃr��S�p/y���{Eud1�}���^�I���h{T�e8Y�Cцj>G7T��� �s�qQ��cC�}Z��ݳps�V��.xp��;�j�ר mȟ�hNp*ی��|�+]r��itA��!��;�Ӯ��n�u9;r�#"
S)3
7�,��) �A� A��X�|㶽�z���\��0�Z�F%�����@_~�Ap�"�"����F+<� ����E�;yǟ:�3�|lb>�q��RA�1q��_�?mCw1H!�@�w` Cm|�x��ep>�Xv�׷���9b�iMU��㢶�PW���(D����m�f������;�������k���=�N߰G�m�=9�����f�3K\�U��s�C�W�l�33Z��X�T�o���G�����8� ]�|q��O6%Q�{�	���"5�TF�\��I��>� �A�BKp����s��~�K�B�_{�<VG��F��}��� ����@�mV����N�#2�s2b����X�\�rFr6�tpOn��֖^�13�t�?s�[��m9�0͊��hL��p��Hɛ����e�߈��Dfj�[A�-��K�+�9�w�>���B��oyM��YխJ��Tk��k�<C����\g2X���&oz���*�3,�33Z��f{�pLzj�s�|Ѿۨ���냈�7����;��PE�p!����Yt,@�����_e��]��D�\�6��kо!���}:/g�@2��j��~�e�V}i ���m��ط�����e$�H�T���s����}uY���3)�M��Bʺ�}�מ�uc�8Of~#q[�����@m[����2�ݜ�jE��OV�K�EQ�x Mt>y"Kp��0c�E���{7UŒT�[�ՙ�6���jYR�݅ �g�����n�����Q,�tZt���<�X�����S2�;��}���b���k��X��}~�*xfߊ��.=KWo�ٱ@�[jHmŸ=S�;��s.Q+>܏ A�q�^^EѭtJevLp���A5��^ m�E�xVg��@�B ��R-��n���ǲ��u
�b{�*���L�5\�@�tx���Ch/�m��0Z�=X��D|�Dgd������m��5��#��q{� ����z|��}���Fvn����� �mȒ�:����_n��[�.��'D���p��ƽ!x�!�3�m�o�M+�#��1G/M}/qՇ�h`�Om�3����,Y�k����+��駮]t!E��NR�䮍�fm�-Z�WZ��2N�����=��'î�������%�Ajp۠o��ƞ���'w������2�4w��W�z��mW<en�h�f��鏖�W܍�ȑ���]�G��7q*\�*I��U�qZ���r�]�W��:ю�`�6$j<�Nݽ�}�}�]��e|��/p;�a	�����՛G����vN���N��3����f'Uܳ��"ۨ:�WN[U�4��_!.���[f�g^��:�R2��SrHg(V9�a��e�3;`�󶂕���b�i�d��c�ٱ�`�ko�%�73Z�=�|���Ù�k�A7�L��ɵiս���N��P�-vn�HE�#�+7�K�N�|�[�ʏ��6�;M��n$I׳[�T�QۗYf*�ۚ}�/z*�*glj麸X��Y�6d^�KWp�������p�O%����۸�*�-W>T6�݂v�̺eڣv{ZɊ��j=��)��<�P���tgL�z�T�Չ�q�%� �u㣗.��ć2��:�����4gi��Emu�	U'3i��T�ño9���[̪�B�t㻵�Wת�H�H��x�9X�F��9i9�eUevous\G8�*�1n�ܣ�PX�ir��rb�Oc=�p�}�aL.�徥�C{n�Mͭ���>�=3ز���q������7m���_�	!��9{{k�vFD�����Xw���E׹�܉��Q0���'}��g���T��ʢ�/41�m�ĵ]��I$�b����lX1V4h@�h�E2Ƥ�&*2�rLR��c%�4PA�,E�6�6�lh�Q!$��M�U͍�h-F��4�@��Td����1�Y�"0W-�,S5��r#UDL`2j*( ��F�BQ���Dj�QY�4(�����TY�n��FزE���h� �bD�h�5���

1�kM)D�*5ݻI���`�E��AD@<����UUT��vrDdq¬Ke�f�p��NS������g�Om���]��v������ys#�
t%�H���{J�� �̖5�a�6��e�v��a�U���Oe����wfz�l�Ji�l=7�AwN��.sx�*b.b6�Þ�����kr�k��x�Q��%.8;���<��9���v4p%�pS@fi��̪�٬Ҹ$b.��Us���d9�k��3v��-p�v͚�2/�7��;��G6ܪ���T(���;�"�Վ�OC�u�.+���[s���v�[f"^띂��s�qj��e���H�9g���Ž9��WN�q�p�v'�tjl맳��\�^gG-ն2�޺�]>$����wD��V��I��n=��@snX��t���j�&Bhz�n�U	^�ȱ���ܖ	��8�*�gs↸�M۬�H��2L�f�V����"م�,����Im�DL?����]� ���i6���P�l#��WEP���-]�;fz�N܂s�z��s�%���;�9��'5�邥���]�M,k�S�Rqd���y�P3y9
U�.�
=�;�Զ��vx���c�.���fbf�l�P����L�Ў�k�Ѱ��Y�&4wh�����),���U�o1"1��R�p�UE1��˘L	l�Z¼is4�
�s7���`ݤК)�;��B����o�}��bs{M,�;��Mh��)Ur=z����k���v���/LG����i��=3��m��u�BR��뎹�άs�nr�c��q/X�Nv��܎9�ê�Pպ�}F����x��x��Y�v,�����2�Yt!6mь٫�rn �
���0���Sظ�Ec�X�=�m��5�BEl�2��e��:�1�c:�Lm���
�0.��]l����]�۪2!�N�M��=W,�z�/.�[A������tt-�Vf�@Cu62��6��n��0[�@Ԇ�m�r�1�ř�m���1]вř��t���4cŖ��\��l�v�Hc����bm�<qE�b�ɭ�zY��ʝ�\���Ws5K���V}�v�^��P�յ���^8�v��`,pơ��S�,s�ks�p1cT�G���fɫs�nJ��px����e|��e4�z�FZb(�Q�m��uz�iTe�ee.��	J�1Q�\���lCM*:�Bm_�ߧ���0]�]����P���of���Y����}Fw��������o���y��|���/<y��\f����U}N""kC�B�3�3aD�|�N�E㿽�߈2 �I,X&J@��&���*w=#�/V����}?^����}���y]�%��%و/�n+�na�Bǫ���S��?p6����6�+���o����F�2rKX��9�A5�@�x���������u���U��U��Z�{� \�A2E>u��ޭ�^�,DO�=�����"�N��i>��9��=�,M�h4.e\G1��ф�f�yH!�����z]�%+����ܵ �����/�mGV��W�!o����F;�AI)�3 �BL(H5՘Զ]�I�+���a&���B���H������a�v$�� �~m���ѭ�}I���ΑK�����5��y#� ������@��mI������D�P�o�wM�ꋵҨWu�k9���9�\]T7���i��u׆����a��U�}���f�}h`Vde΂�[���A�w)���/���.��X��ṕ�� !��[�q���\����Nl"͠�����~�͏X��
��f��M�1)]�8K�_H�A�/�͵$6�M�ձ���Eޡ?��hm������eCS�r�A�ס��S'm�=[3��u|�P �[j~ ����f��dLB����ʪ��o=Y/��,D/h{�}� �<�?�|!�+�w(32+��|�Dw���Xn]k��щn��L;�b�ܦB�ifX��k-�&�L�����׈"k���7}��1�Yu7��R�pN{��z������#7�.;ʱ��s3�s2��o�u\�(�	�/7x4�@��<�G��N�5Gpܮ	�G�^ �mΛXIz4S�,w�O ��H����C�������rꙉ;�]P�!3NnNU�,�3]�L+ι{����u+;�Yj��:�����Y
�,]��u/�#�����n��C���X}nqP�U�˿S�~�L�F� Mt��$In ���܁#DmG�:�Bw@@�}"~!���p�޷
�=�J���Wڮ�U�Y~��;�����V��H6�I�駣4���4e��w`v+z�;���b���?W�|A� Cm}!�5}��p�韴�ʒLL��R����eP��GX:�3]R�r�� �k��kJ����>�x��RA�r$P� ����}�e?{�0R�`=]隸�DY�$�@��۟�[��,��o��p�D�ȟ��;��<7{m��¥n\p??j��|[��װ�L�kﯭ2A�=�I,H-��w�Y}f�#m7�gE{n#7��p�p��H&��/`"k���p�:��b�ۺ��j��ȶԋ��Og{�O�f�����k�~�܌G@�����2�Vt����Ӫᗸ�ꄥ����]�����r�n6��,��FOC^_w[���V�����?n�wGD��h\ʸ#3,�L�?-_>�ͯ���B�;ō���ǰ;�A�/�[A�"Ŷ��ƪ��dA-��
�\{]v�ƈ9�:��tt��Y�[�x�у�f'65Z�\�/G�b�(�g��5ʱh.o��q}=�NpǸny
�=���~w�v�#��OŴn��"��v�m���=��7Ё����{kӮ�9�aO�&� Cْ$��U��߳+��z ����Oz�H�I.���ӣ�!�N!���Lx{����T�\w��������|�m�!��m^�>�E����ۑ �G�����>7�=��y��k8H&��5�ƽ���]����$n9�~9�"�"-� �_7��ܽS�u���-V��ܽ���^�\2pS����=����/�?6���}x�{���'��jȁ9Q.k2*�qy�s���c3��<��Q*WZv���Э�A��-�*s͆�N^n��o˰b�j���ee�!}��_UX�Jx��z�]��Tm��]]E�T�s��s�kr��ɺ;;���Ε�7a�L=�%x�F�+�d���M;�G	�tF.V�t���S��ŗ��lq��[�P��l���A��������:ֻL@V1��m��[��m@{n��`lf���9��Q���m�M	H��F��`�z��SͱƷ5�vx��j��-nr�w:�}����xw���RQƵv�adf�m��3��>�b���Q�n�(�/��Dv@@���Ŵ��k��ssT��
�ˎ"c|zK�;B�߻ޯ �t#�mI�� � 6�c�:�'l�N���@���Cm�����VJ��7�i�	�B �z�6��l}�;�O��{N�RA���q@��X����k9�!�g�5�pd�0�E�|�����BKq���6󽊸C36���@y羟��������uU��ˎ^y|�6 ����h �}����	-�$�
GO�j3�lG��/U�ېo��ِ���o�j�{ۙ��{>n�x~+CB�x"J"�PWvj���1���A03me�De���ރ�����H�[(I�o����I_/���ڛ�۝X�j���`�3s(N^L��p��'�s!-�D6�H%��s�.vzb<w��r���yT
2E2^��M��b%0�mǻUt%�\]Ů�� �i��Z�Vu�Vz�񪈯\��8����Mר3uÈ�韎���Z7��.�:�b{�A/=2A[A(��~g��U�
6�Y����?6����|Am���$��'>�Nߜ\3�y�`�|6�O�p� ��Cng�����'9ʬ���ז����Ŷ�77��M_mDc��?ހ�"�E�n��>��g����r�p�-��m�yY��ʈ����Iy��uJ^�����/�����~-�����~��K�a�[v��]��sO��M���7\a<hM�Ra��K���?�?�_�$'���1�A����{�z�b�4/���H용-�w3~�ԡ~�A;�} 6�n>��mHoT_;~k�E���;�^�l��*�ڈ�)�{�񮀾 �^H��=}�U%�Z�� �wH%�D�Aۑ?����Q���+}쿊U�>����V^�M����_7���R��UR:�pv��eURb��^���{T4/���pL�y2�+%�ye�j�T��*w.8�y�$7|q���"C+#�!-�P`��/�~�<�c�ȾC���3B�k|'�p�~��r�9��
|*/�YX��Ÿ@�mH ����o���:�y�U� ��#����F�Y\1�</`p5� ���������>�h�n�V��.��wb�@��:;+����űp�����f5����6��|��A��Cn~��m��G{����^���"2�ϪQ�|�],��@��S����^$G=����&8h4��2�s7�M��"�/F��X ��!��S��d���A�K�	�ꟈn-����m�0nt#�pF��ڟq�K��c&x^��[}�D��"mmȐ������Qo���?��w{���E�TK�T�\w��U�;.]�NX��~��\u�4[�#��!M��5/]q(+���ż�{�_���6��W���!*^�����y�^ʬ�	S�Ȳ6�>�"=ܧ����D6А[��5Ǫ���И�������q�瘊��H p�7�!�˿��?v�5\�|dZ/�P����6�X1�ƛ��z��\k,9����P�!j��t�����Q�1��o1I�/�q�-�?�j����Y\1�</y[<�iO��F#���t�5ذ}�D�A$�)v����B��߈�zg��j��G��^�D�N��	y� ��������x��G5ڤ��}�n~n<�2���8/�U6��3"�<</E���R���m�����u�O�2���F�|������;�#�=�c&tk�հ" ������Q��"��K2W�DH6��r}��C=��x;���T����'3�A��q�|[j���ވ���;��P��&9$���U�y%���c��z񸰪�39�g�.�Y��K֐�y\��x,��;�Z�t���CQ@�S"&P0�p����]�dy��
�3�^.	٬��\F�Z�Y��clҚ�Ae��2�2�3k��`�c-�ƭ/��[]u�8�N�8�J]b�@�Qգ;�v��;����;��|�q r�IwnɃp糰���������X��An���{�X�H���f�G7:Z�tR�2I`�d3�NN��vm�P%���}���jKbֺ\��	�4+1�]�\�kq�Kڒ��ݢR�cJMO�|����0�ܑ?�[Cy�u��v�y�Lx^����w�w}�b������p���@)�H�jS���\*>�� �{�@~���l��T^
{�b����Ȑ[�ʳ��j'4Va:3 {�'�d^B!����'��hR*��Pn�"c�a���y*��#�����h"� �^6��\����U����H�{a͠���^]�M�A���A5��S��U�7T����f �p� �ڒh/�p��{it�J�`�R=�s�.�t+Y��&�^H�[���N�~y���1����׭-%��*PZV�R�Vт6��z�ڲԢ�O��59��Q@���jotegz7Mj�%i������U��s^���D�^�ȶ����Ÿ&�x��n�
��:�z�0��r��fnf3/=^>û��`�`��U�6UQF��J�3��O���X����!^�:Y�&�����8~��������ro0�P����N>��_۬�XU���>R����`�")�����h侢v�nWG]ǽ����X�)�{� MlA�-Ȓ�|�h/�m�+d��j�kA7vg��m�_.��WޙyFav\}��5d>(��z�-�}H�������P�=�n�������`߇R�������a��|��O��E��k��&~�TGˆGW)X�R$fT�Q���
�[��c��h�?v�_����'	iy���o������ ���A�Am�翺3�;��R���m^x�)8��W@d��?���D6�H%�@�s���������� �޾]ޞWޙ̨�\�8�^�$@�O{��g�K��Gm_��������g�4�_��[��@A��΍�cuIf�j�-��V^JV�֧r��1ܠH�n���>�]yz$�
rI+�f�˙�0G���goeeIc�`�r���ɖ�:�\xF�w�s��ZEۢ�4*��Y�Nn��^����յt&�:��We�e)�'p��=�l��sǣz[���40M5��se��5m���؛����ttkDr�se�0J�X 72��ˋ3�n���VdS�%'OTA1u��܊���j�s���A��-�z�ηo��E0��*�kl� �Z�4�m^������y�s��3.���WyۗWt�h�z�Hn�	X҂���/BW}[�U{���v�*�=�S�[֝P��Ο�Z��72��v�,V7OM��]b�����ݴn���BO��H��Y7^1�*Y���}x���]*�����zw'�1Jv�ɜ)^l�\�.�CTM�)���Wj�ZD�x.��ңYԷ��S��U�U��r�cQ:��v�pij�����>�J��'3mf{�v�롧����]�r��וe�U����jUK*�Ki�sytL�꾕�ݎ�S���CF�vK�b��tٕ�oG+�kB����ٝr��{M}K�r,�
��u��o��t6��M�����j=��G�}��}J�Yq�ܱ�����~V��{��^��lf۞+1ܿ�̻��J��n"48���L��uc�1�꺂ӝ���U�U��k�]�����UP�:w��Koy��bl٦bwU.���X�]0i�u*:��.�3�G�lD5�|��e��Z���d�`�*1E�4_
鄤�1i
J�QX��Ւ�ŋEF�h6�&#X�MQ�*f�5��J�A�ݸo��"c&B�61�F湶*6��h���J���3E����#F�"KIh�!W+^k��<����r�\�Q�	h����s�4	�1�Q&

��.sEF�v1\�2lb�h4Y/{�yX�������x��F�y�%�5��~��ר߄�Ch [��u6jı�f�_Pv�;��͵5���=�]ފY%)�9}�#G��f�ПU1�kc��CnD�p��!��Fb��+'n�~��W��=<��Nd�� ��� �mn>E��_�WL�z7z�$)&q�u��xհ���(�:��>z�����OFh���2���{�ݑ%�_Ch!��w˪Dwc�1(�o�W�5���滺� ���%d�A ��E=��}ҚϽ�� ��V�w'���RX���|}����H-�a��B���A�П�t|�mCm}?6�o��d�OI�<��)vzZ��9�
���~__� ����EdIC�wvs�l���"�$H6�����ܾ\�#�a�F�m�� G����.���S���K6���1���ie���2h�Ǜ+�*O���=���:�ݧvGW�o�SǬ3��8��.e���jL�G<�?o@@�H��+ ȂJ;~��f����4��#ݙ���k��I`Js�p8lG���"�}��6Dm�؋��&T���:�û�Jx���95�:��&�y��h�pJ�jrA<��"�Cm}!��wZ���Ʌ��і��U^ծ ���B ��Rm Im�_����:��m��PB�/�u��0�F�m�H �B ޠ�m���8��no�Q���0=x���/�p� ������z���=w���U����?� ���%h"J�܉�ǯ��&��^Ez�@��������z��uƱd(\�w�K�S��o��{B=����$7�ۑ �U��{��v]����׌�Ftm�_�E�����p%i���㈈�/h��ѯ��o-d�؉�����!W��n,��=�w>:���lof�YZ���c�Z�Uʯt]K��2��i���[,U�tY�Zr���8��IF����.5���re�;bNx��\W��.��LY�p�9�v��z�-s�Ju%t���BeŃB�u��=�uXnr�]�;���9�==T�����#l��in�jЫ14E��+.�.k5�/{7�s`��\���)������sӅ-t�F���خ���Cs��f8�\�n�]�.`�rE�V�r��5�֓+�|����0��X�����ф�n���@�Zlۙ�����D!mG7ؤ_/���ڬ��O˫w�bp��_!��5�_����?g\�;��!�!�2	n"ndy��^�韏׈Vww����֟b8��q����k��^fm���_W'T�W�9E�32�G2�"�%h��N���M\��^���x"���_�/`"r'�A|[�A�9�>ܿ*\�:�S�oor�]]�A����� `��Ѿ�� A�As ��h Co=}�:d&|g�;]�o]oS��>�q�q��^� �m|�W�[j���5KGQ��rKj%S*+E�����m��k��b}������<<Xv��Ĉ �ё�}ْ$�[A�om��Qk�/B�s��7ʍrF9Wi�9A��G=����E�@�[jA�Cռ�l�k���q~�P|dWK����T��Z��I�&dժ�V�x�m�s4�u�=H�Ee,��{]{��a���d�5�xg�;�ބ �9Mf�r�S������@�}�Ƅ��e0�j��zc������������|��r'������^���~���#���A�RA��� mI�q.=�X0tɸ��7�"@-����{sn;�b�/B��s:A.�'ۏoк�{��o���z�-� �[k�mq�����v%!���Y3������@�}��9�n��&�٫/�}k���s
n^9��uc���.f.����\Z�DȒ���:A�l A�A�_H�����u�O�<}1���M"/V�S���}m}�~m����@��G���we�7%�'��t A�{ٝ���6{r�D):73��p�z�6�on=5�"�R�ߧ�d"	��Hn��Kmb���F�}���`�L��q�J�Mv�=���������n}�z���:l��߮�=�tX���3�1�Wry3j޽I����w`�WF�~~@�}� ��-�����܉�,q�SK�q�z}�?�h*��޺�u��"�28���"����B�o�Y�'/����-�[�Y�!�F�z�U��'F� ��c۳�l�{0����~wK�~A$�$C#曨O�W��ϧ��/� ;Q�܆�]�i���n�$\kI��n޾�`G����P�o��@�<��'��O<��-�����\�f��R�,�_|��gc�����H#�����D[s ��|B�&�>�(U�'�1����u��Ի�71ّ��w���E��� �s9d�nR`� �/`"hIn ��a�.";�Lp���t�^1R4=ΰKt��K��"D���S���]C�y���}yA-�/oV��NWu���ap��>�4E�����r�]Ar��7G}݇�vs��>����1�~��| ��w�sZ���N�������)�I>�1�!z���t|�Ƃۙ���r�!3��ިߨh'����;�%��+�#�'q��[_7A-�w�g�c�j};�"�J3����K���T|gi9�;m�7�p�n��c4r2L)�av� A}?7x6�������=�x�EP�{�!�ɲ�C_��b����g�� p����xz��m�oaM�S����S�]c"�\5�����9b̔����!Ǻ������p9����ü]nn7�Su��z�p^��� ���RCh!5o��M�к5l cr$�B ���íw�Ou���P�8H?�A���g{OK��@��_�����%/� ��A�d���u�x];��g�A��y/���,��J!p��{������~��;w���*<�t�Qf��$M��(�F�h�0�[t����#��<n��K9ҹ$v
9�:�Uy���P~�0tg�e�{�w�����J��G:�����]�����{��Rîݜ��G���^��mՈ�e���!�����f���o�t	,�&�-�W:�E���1���`mf�Mx�g�l�t�:���3�;KpV1w�k!ͷ��c��zc�ݖ�����E��Ն,j�Q24��fR��/lp�c���Y�<S2���eWsW7h�塂�b�v�Lg4E��O>�����kb�g2�obBKӷ�����)�1S�H]���'�?���F�o���]��}�j�Z��g[� ���Z��x��^_?��_�@�m|�|���N�������C��!C�=�c����.M*/s��A�� ޤI�w^y��^��}�
�>�@���j��-�?6���<�Ow�b|�s�k1u���ap��k�/��hH�D�D6�G�i}��[�5{)��D�~m��w=������,�=�p=�I�Ln�q�Q�{c���Rm|�-�@�ۑ?���ʵ�+�8.R{z�E�.�,��T8^�} ����@I6�"D�iHй�7�"��J�7V�}yK)�nN�͕�PB;)�ģ;Kss�++*|؋ �[�$�|�}E������d���"|�.�B�����A�d�����m �_7l=㙫oc=���(��7B����m�����p�2ʩ2�aQU��z�z�鏘��cՐl�u����u�fR��&�!\8�����{P@{=��y�+��F,�=��5$[��-��6X���c�����	 �܉��HD�n�2zW{C߮ז��{�{}|�����8H'�>B�����m[�Dd��uC�1ǽ��r��y{!Am�o�ٞɮ�Y+ȥ�_}���#=��O�3X�}q��
!�2	n�7~��Į�Ȩ{���PB��_w?D���ŐWy�	�k�q�p�%��s���~���6ZF�1�f\(�m�z�gq��ۛ���Y-�4��M�z��K0�rX��,����7�뽃�]:�)z�Q�{�!{bZLg��$�V�#^ȟ���p� �[jH��ļ����v�������}5�VJ�)h��k`"7?[�î�tΜX;�b�}?O�!|AmCnD�ChV���������5�NsصkɈ�zn��~��+��Xʥ3_Y�}����"�_wy�(��am3寮��=�T%ܱu����Oyۏ�w^�*��p'I:Tb�o�4�0b�+�����S�6�n(��RChn�]�J�ǲ�c�iezD���|A}w��|{�vR��Q�oxH ���瑛j�b�@~���~�A [��m��E���y=����v���֞NV�r�\�^�@�k`"��%i��~+s��o�>D�V�7(㋯5;S@n�WA���,<�Nۑ62ks����o����~ۄq ����p=�[���&���X!o�q�y�{g.(gN)��;����_7�n#Zu�1QQ�flȈ��߲M���,�{��x[ސ@1���$e~hK3�9������jA��q��0������I)麹��K.�%�����D���x��"�,n��̍�=)������@t��{z�%�Ã���;�	�b�C��Dʯ�÷[>�5����͗$E���e������O��q�;tg$%<��2]a|re݈�7ڣ�q�vmm|R�l�&i�c����c���&e��m�%��м;���}�F���E�w�c��C�wH�"k�m�~��g���z㇄F�1�(@����lF[�0=�!�I�'�����l;��T�}��������RA�^��� �ڑ�\=���]җ���{�yg�{\��9]�W���Am������" ̮�9��Ԋ��#����w�w���o�Q��q��) �$A+s��~I������	�����ǁ6��sv������]��-�t�SY�Q��{���"���m|�}s��c�{Cv���~�A|o�KmO���������U
8^�Ӑ8�[݁��B��'}Fj�ng�������+�6ih�V���:z��ݚ��{ILF��u�n��@�u,w���! ��a%UY��km�+U�[o�Uj�ۭV�m���V�ߵ�խ���Z���ڭZ��U�[o�j�km���� �	'HI(�@���Z���Z�Z�}mV�m���V�ߵ�խ���j���Z�$� �	'��PVI��f����A���@���y�d���vO� PJT
HU 
��� �AH�( @ )@�*�D� ( 
 (
	�  �(P����
	 )@)E�@IH (�P�B�J�( ��>���(@�I%H���
D�ERR��TU	IU
�BT�U*J�E"�QI
 ���J%
*%QB� x d|�Wv dTn���(��!�A�� �r ��[�s@2��D*�x��<���=� =;���H7w
)�P��q⥳*���W^<����Uͥ倡s4���K��͔墊�U�
 (��(�P@��	EJD�T�|=
�����-U!�Ԅݜ�W:[��qUn��n�9f�*�TQΩfjE9IAEQ@��(͠U��&qHn
d4����TM��J[�ê����������TDPU�� |��D�QU%IR!PD���:I[��Rf��tR��Y�r)�B��n��� 5�QQ`�#"���H 
�� ���pt�%(��4 �j"���n� F�C� nà�b@� 8(PJ=� DB���T�PH���� 2@�`�@]���t����"#B!�@�w ���
ɠ�5  �U�  ��=R��J� �  r�� 뺔Q��@�@݀r R��� =�� %�UJ��J���L@۠���� �u�A�uT ݃���w�p
��� h :�$
� @��d �%Up �8�9nw �� 7EW :�� ͂���A���      jzh4RT�#LDd� M Od�JU(       ��T��JMH 1  �&�M��L���       I꒐�T�      $Hz�Q&#F�i��G�mF�hl�jO����>��|>����*=pu��q�ֹî���{s�'��(�"�
>����!�=����k�C���%�(
< �zp��G���G������6� ��;�A�KH����j �
<�>o�5^j��@���~?W���{D{��y�iD�j����i���7Co�է�����_iƂ��H�|���=:��Ó�W7�W�Y��xR��]��J�uf^�Җ������Y��%�v)�-���B�S:���;��[�2᳋��Ѥ7��vrđ�d�@�6shl�I⢴SD&C���n�����n5���j-��L��b�;.�Y�w���8�D��Z���M��o%\�9��V���l����Q�z�۳��b]f-O#�{E��]�7��ˌ�q6�[�ѿm\�M�cj��:��6�7q�4���`�^�Zc5�2M�1a��,]8��{-�Sp��{����dE�F���D��u���lr9s(X���;�Z��f�)ϥ��R�R�umMI6� Maa�V#`�T�$	Ŧ�]!G71Xw�-��t=CW@Y�N��deͅ6/ۨ4ȹ����)�����jh�f����dLj�[�n������@��6�Y�.ΥzL���d�����9��t0��Sҕ�5�QC1Pvr�ِ� ��V۵u//V�j</sM㩵��@�]��a�#p��,)�F��~�8��&e%sbDK�BX���M5�&2�1n�n.:��s���u?�M��R�q�ff��0o#02���8�h���z#i�D�XBeQ�R"V��C�cP���Qnf
p��o2��hdVm�ڱ"�."�WM]Y�OŚ*fO�g�5#Vm&`+*�H�)(��2��t��4�n���,�h;v�	����7Naϐ)˫٢f�@;Ue�_ѻb�ٵ��ǒScu;gD�g.V]�&hF^�1n����qJ�����i<Y��U��J=b9���U�%��{w�a��e��N%v�`iJT�<��'f��*ڻ���3�>���������R�j�s c*P��˻R���ɨqS
�U2h�#1��TF&0J�.�(SeRa'����CC3.^(Yjˠ~W�Ǚ���l%a�v3k.�k/6�KV����d�3"��˱+\���^Ԏd�
1�h��ɩ�+c�E��	�ܳ�݃9'!�3$��PM��NPܵ�Z]�;��b͘wO,�l8݋ۘ�ؒ�	+҂57eٷ�1<A)0n��e��z�Z���r�<# ��hhb9����%���t�N��ܶt̋�*W��0U�T5��MU�J�S.�-ݫF�e �K������&==l`BJ�U伭1��#r©��P�˴��k����h�&ݰn^4����E�@��˚��*�m������9Z�2]�r��e�,jc��l��%GA�BZ�8��pR��M9̈́���u����VPk]X�+vmK�N�;��V`ʼ#&��n����)J5�ҋK)��۲��c�6��K�B�e5��#��Kʛ#*�f�J����a��֑Tk��y�A�6�vo�[Z2�f��V�7��.*3s(�î�3����ô�H�mR�Oq�@�xͥt��܎������c4SJ�e�Х�-e�!��P'e�K*ٖ,�9j4�RwQ+����N�Í��f�Xl�w0�'S3	��"\S4)�B��L�mC��6�iW����q��w.KUpF��m3��$�L'.��JeЏPY��V��뗧6���9�m�K��ABJ�zܠ�0 F���f���Z�kWw��0�ɻ�<�#V��$����eh�V��*ܷ��lw��,	{sB{,�0æ{4��^%�`�v×���z�XW1=QءG4����V*v-�
}�RLԲŝ��5m�ԅ'�����+�<�.p���� 2:�#7/���Ҫ�
 �YF�3���Ȯ�Ӷ�v�	��&�֡94�V����e�!�lY$Ay�+�14&�wV+�����kV��r�(�

	�j�ז0�I-+U�Xf�Y�bR��B�n0��y��]�D@�W�f�I����J��a���u���
��ݫd�"�Am,�A��J5h¡�n�2��NC�/�b�Ô�ɚ0<*l �B�h�)*­h5�� [jJ ��&U�&;8��RO(ۀ�#)��I���%��5��6�)�	������+N�v��pœn� �kV�r�{�Q������鱗xndW�����@�J<Wa�ٲ򲭙D��3Zqh+�!��@�6��݇73+&�^m��XKF��<��d)�HG��AJH.ۧ�㧈����j���K��d�.��0�]1ނ&�00e��U�(PAL����hm�*��Xa*�+.#�ɯc��y��Ա["ڑ�.�/!QVEDE�,+ �^Z�K�A����Ҳ�VM75��B�����\��I�V�ԩ	g%f�6�Ա�X�г!�D�l]nn��ˤ.��U��e�Q�@A�#�@ҧ{[�
{a�vt^eˎ;i�)�[S&)NX܉n!Z��[q,Z]`���MӒ�w�EK���� �nԖ0f�n�����(��+2��3[Uw/�٨��v��]�n�v�k	(e�|����w�����3T��� �� �*�[Y�.�j�b�rG7�7��r�U:4QQ(�IA�'��V+!�l���܀vkZn��
�EZ@�Z�m�&�%t�X{j0e8�
��n��3ţX̫�2U��2T�w�tKBkۂѬxu;�w[WJ82�@���1U�N�a�[b��Y4!wPN3&H���M���:��B%���ؘn�ʃv��XF��gY&�7��f���z�����Li,Hh틆���pU�2�-�j�wO,��'�W������$͙���E�����q9,d�e���1��Yp�1R���q�Vسr����Z�MC
+ͳ�v�P����ܨb������`'jv^��薀��aL�u^X-`y[�,���$c6=y�ai�okC�D95�jL�6�wz��À�=�����e�qY32}I�.��K�%���ٗ����o3)әT����Yy{&�jE S\�Ә_���L�u��!��pKg���4Q���w.%���м�)����P F0��5"%M2��M��&H��˩���*e�XrY$l��i����Z�7)Ϥd ��U%Y[�&�v��w+&b @�5�wVl貢�`D�ۺ�3	�4J�w����ܭ�sI�2���G$��n����V���I�Vi���f(���l�Y�(�φ�F���J��AE�M�z-jQ�qj��;��saB%�T��T�NL�I���ɠ��ܴ6�(jv���HE����%[2�Ej��&ز�F@�mʶ������YenB�|�%Z��^�0�Hպ�B�=2�+a�j�r22��R��;ck"�����l�-	c �+��XDU���Iht�S7h�E;קƃ�Zk-�I�ĵ�%���z��6 �#��y������lcU���L��]�[1S{��^��f�(�P�x�%�T���,�M,���2iЁz>X��Ĥ��C&X��K� 4�ֵE�Xpl�n�3�ZH$i��YZk,K�I-j��-9MÍe�xfէ@���4��T
�許�Ņ�o���P�Ö�N��5��P^ɏ7�1�ՕxP�0fr�׷+3�9*�-\�N�V衊楮ѵ2C�X�89��x.��j��-��,���H���waj��2������ⲳ@ʍF�(��n������Az�Ee+��/���*�,a�wn-��+���ʶ�wF����ge�@�kUr��ږUhtȤ�f6��6��]LxVD��ʅ
��V�$��M���4�8nՏ���GBd�r�Em�1j���؈�x��ʄ�R�6cMe!NƢ$��Z�QY#%۟s",0�LJ�M\f���x����ӵ(r]�ɩ)�����f(����'0�0�B�B�	�CJ�Pu�E�6.m)\N�eC5
��F�ʡ��嵂Y���}oꎳDՇ+@�ؠ��w+,Q�+YչKm����c���@���ӺV��l��&�*VJ�Cfu+ธ�Tv�
Q%���`�"����l��Ē|"������[I+��0��nF1Sr��M�R7"�d��e�j�.f��X���vo��D��d��{�i��.ԩq-�Մ�Yi�q)N��{���՚��(eX��5�V�t�[^4҂�a����m�I��)��e�ښ65Z,���x[M%c*�#-��l� �)[����e�Ԗ�2p(��ޫ���A�B�'������c��m؊d���z2��U����h9�M��hZ��VC�6�"<��{�e���f�E�El�c7aRE(R��t���X�Ytմ���#��,�ͭ&��S&H�yx����4�W���YR鳢�<����$y���Ikbۣ�\��JԈ�rVLv�Mj�°�li�V��9������Hve�m�̬�N$l��*R�cGIFm�*w3i��H�4R�
�׬"��5��[�l�X�'.j�x��Ŧ�sb�y��|�:l��7KSv� MX$f1��6NF��f^���]c����3T����:�$i"Ő����b��P��n�Ҁ�x�[z�,U�h�QSf��Ej�F�&�6i�W��*Ӕ�K*�Т�Hq�XRؖ�sj��%���q�2�06
qT�M�V1�@�`cp^BJ
*��A,&�s^d�ȷ�����Y5p�� 0Mb��]YD��rqV�k6^]�m0�Q�tQ� oYuf��qa��ɇ"DA�S�eQ%L7w�wb"᭧�r�H�P:RnZ����J�X�A�wWx�C�B�B0Zqf�+fı�c��
� ��ՕY�����[�L�Vº�*�lB�d�컕�5�E�s5�U�R*i�R�f���[�����Ct�yo0lݗ�S�%F��{�c�Z#@�X��F��ov��Zݒ�ĴŊ]�v��r��љ�5�AX�+��]�Җ�Hm���e]�sN���;��fL+��a˨�-[!��,T�vt(�ӈ���B�:�#f�m��nT�e�sr�X��s6ϬDa��;I(8pзW37 H&�%��i��0GJі��l�&��Pnz��ו�T��'�b�� t�X�ks�щ��n�fI��AAtN���(JдZz5^k�u�D����,t��P��A#W��4�]i�7a� �\��]�(����e"e�
PGr��/ZY�q���ᱶV�7�4�G���	5�k ��[%�ŷ�5�١���Z��&�nn�*��oHơʂ����qG��J�5$6�Ūv��N-/�x�tѲB�#r[�pҬ̥r%kpAtp�R�p��^�z����C��#�*�����͡�(Zf�����K4��/�hV��e�e�P�u�T��T�9�Y4\�2�Cb$:�ٟa�-��Yíૻ�6,��R�����^�hnkUw��t\d�jVͼ.43��w��ޡ,�sVf��P���I�ql�9��/E^*��n��O�]�m��Z���(�����Bu� l���ku�Rfҡ���nE�^+�,eV"�&[�-�;Y�
�.�%�3�Q���ͼsK�]䩐�(�;gS��]�,l-���R:#)�o��N�Y����:Ӗ*�����kk+JԮ�dؓ�YY��ʀ��wkvS͚�+e@޵1-T%��L��	�U��j*�LiG�{�l�y[�ޝ�K���4M�ne�CS*[���kw�X1T(�-��ܶ]	�3��yu�;I�Z�-	J�N���n���p���	���i�;�T��8��L%؉�i�us[��I�t�����^��y���a�ZQ��[X.��e��E��!���J��RX���p��ڥ.�*v�J�@� �hj�d��(M!�Y���m�4]�N�Q��3V�0����X��!/wt�F����6���Ʌ�N-��&�f(U�����S+9Y]8���"�!��ɪ)h��,\PJQѨ��(㘶�F�I���z�jߦf�t7�yi��"/RY��B�D$ڬRq��t����˸(�&D��]��o�\�$<�L�d�y�1(�ө`os*����G@�b14��'Z�F�0�g$��۵R�b�E劗U2܌���1��r��{��Ϻ|cP=�����yaGI����w��=U'�Mg=qǻ�ttr{�� =�5�[Ջj�-kcm�(�kcmX�����ڍ�*ѵV+l[[h��X��E��6���֬m�k���FՊ��V�F�Ƶ����F�m���TmTmUF��[Q����[kF��Ū�j�-�Ū�Ŷ�mTUQV�*�E�E��*�-b�QkQ��-j6�VՊ�ڨ�Z�mE�RV�F����h�����ڱ[Tj�-j�cV�[b��5�Z�m���TmX�����+mcm�[kfA$VDA$�D��o����Od�<�g��s���_�Ukix��AQ��_���J����G�?�h���#�������,X�k�8�����s+�'���6VZ(;�G�]��U����9���W��IS�ԭ��؞ÔpP�̲[���'�7U�u�h
��]]e�U�����ە)��^ -��J�,�fI9"20�A�eEƊó��u]bۡ��#��H:+���Z�h���>h)�	�!����E���۔��$p���ѧy�owc)�WAP���C�)��]]�M�,�2�Y�C�]�N*�*С],��U^�0d�%�2����*\BLu��×V� ��1�E�F��]���c�m�,�����)Z���ɻ�ጫ��ݺ@��m��
wF3w�]f��9�Ŋ,0N`_!4i�O^=�\r�YV ��Y0,�5�C.�	�J�56����bf]
7`˾y�5��� ���*����6���5�r�1e�J��w�����R��q���f ��ӓa�{uِ��AA|��@Y���ʰ��5K�t��A4��÷�h��p��*�n%�'PV�G%Ό�1jFV�sbB����T7L���҄����P�X���f�0�b���nJg�b��oWq҄�+c\e�%�m\Bs�3pE��뜙	�R�R�[��<��v���L鎕�َ�i��Gk�Z(���>3���r�hw7��"�
Ά�Z9x)��
�P�2�F�:��|h��P��I��J����nY�*6�F�k�N�4Vľ��f�3���˱O"D4d�ز��Z-�ʝ�sa5uֻ�ӌ�uv1a���D����4��b
#�]:����ªhm�f��b93��T���h��Xo&f|B�Pu��H@j�bѩ��ۘ�.ui�&P{*�+��G��[`
�;�J���8OQ;�X�<�uJ�S���ڼK���r�7��/S$E��x:��F�%�g[N�-v" �Wm�����M�	/[t$*gqҐtτ��r=-��c�A��pǋ�7R�a���d'�{"�F�q�{fᛴ�\1Xϯ��'WZS�7��٦�F�ێ��ݥ�Ɍ�´L���amt�7M����)�� i��sw����	�eԆw4ea�̧sH��N��4��V0m���ú�*��y�U�ʰ�^�2�he�g1{��l��;��B��WL�x��Ὦe*w����F=䀙e��+'l��_c��Iׁ�9f��Kf�nh�S�$Ui�aLy���Rz!	Qj"�,��)E�ɶ�������J�NJ�����
+��a��%r�+t�p#���l�b���7b����jyel�!�ѧ��L<�*�[հӣ�t�轣+�o;+3x�㙲b;F%H*]ԅ�y�*&�.�t�_�h���"��@�Ș�g!e�U5�lY�*PQ1YqET�*V7#%,f��/��Ђ�^�W��C���!��6�\$|ʨ�q;K6�v9e���XlN�ll�Q�0'ƙ��\=���NP��udN�|Ve��I�n���hKW��KѻN�[�bm;S.�7n�W[wR5ѽC2»kUq�Ƅ4��^`�Y�!��e�tn�M"��y��Gw*ेj��켨�����+Sw�o!�ZϠ�wwYC'2�����SU������m��/B�v�D-X˻ޱ���']��~�D;9�RZ.��nN�whl�Rv�p�pʿ��à9��m �W�jޕntkfQ	m��o�)�}L���A8èI �YG�q��Ґ��7i��e�g:��dU��%$�GD��3#.)3�0^]�m���y�L#�ƹ��2d���YYb>�4�j�L�`�9�R=�������*[��Y$����#2�l�ܱ7C���ŉ���Z�Ȭ��*1�T�&Y����Ah�yF��d�y�IY���H�+ �����C`�N5y}�w}έ�G�$�/-_Lh�]`�ՍH�=u)!pu�̻��1���
�6�:	��ؘs-��n@[��o"�G"�3�$-Yr��Z(K�2���kqF�f�w'8D��+t�0_ەם��۩zF�l�1��9+1�������f^��VX�e�X��aM�����M�+*آ&
��W"�,�V��;2�fJ�f�'D�m��ey��L�����-+��HY�N�"s�DiVD�KN����8�.D'L[��>�ݾ�9��̮J#�
W�ر�u�_Z�Nm�xt�b�e�̖�<ʈ.Y��a�=oP�Y/�j�)0�b�l�rd�8ܩ�ȓ���m����Y*�Fa�X�˸�u�p���3��eҀ�K(h��]���JX�<@�$�c�CA���-oB�=�a�Yi��X7f��h��.A�;ӗCf��:��\�-_Y�ign]�-�Z���U"�,p��n��F���y��` ���e	�P�)�msV�x+�g�w�kC�D���P1�-9pW:	�`��d::�@�<2��J�
L��мk"�4$�g�0���RƦm���[�}���L.3���Iǂ^^�u���.Ta�#/F_�b��9����~��d�8�U��q��x^ �Pc���@3Wdݛ0+3F<��xuB ��<!���>6��\��9���&UJ��|����s�AS(l�m�f�v�)�����=2��ɮd����V�ˢ�I���ڱHkk���v�y��N�B�Z%���B��q7H��mK�M��nͶ:�T���RUK�CU�="}��V��q��V�6��X-�ü�mi�����^�%�3��'|;�}��R)����if���Z�v��O���wL��	�M��Vq���#dY�&MY9L�D��0�3&T����U�KO[*�HpV/,E.����awBf�IX�%�5��X>ש
6"n�R�n�<yEA.���՜s��!N�9׸�N�A���W1?���5��)��`W\�u��}H��o�1��)�M��e�eH�l��dR��[8B�(j;�YP�Ϧ-*�]�$��ұ�J���)��w[�cqwL�����&S�l���e�C��k�y'�����c]L�*&Uڋ��IoQ�zc����t�r�.��,��csm&�+�� Swױ�٩�z��֫!f��2')�(�d�Ԓ&eZ�f�\��,&�Q��S�B�`ژ7.�=*�oV�W�9��_󮢩���ֹ�[� �`�Sx��>���m���ϤUu�d��1�9B���]�+�������E�V����#����}4S�&<��^�KH����B�;&od��[N��b��v��7]��t�ۏ'hW�Z�U��!td��8��������z*^�ɜ#7t:���[{M�^b{���r� q��i6qP�f�`��7�D�[(���Ӎ�b���n�9��k��f��v<܁�_evbjE�u�*"���8Sޘ�&�F+��n��r2���k;oI"1ba������2I�s"�D@{�Ժ3v����X�-2��w�*!���9oMQL�"g$
�I�Ktuώ���:�{�kwp)�J�[��9MZ;�1v�����]u��2ne�w"�S�#e@���N
ȓ�,�BEH�8�)P�Q�+�y�l/@�>ΰ�ȕ��K�h������B�Cm�'ڣ�� �D�0��j�l��ϢxPT1���j��S��i���}ۉ�ERs,���lT�@�ݟn�h|h�dm����y5SAm� q���ShBB�Ʉ�@���̠�Z��l�(6tÚ{6��w�Xg��2��u��U��g���zA@�Y�3�3����G��>u��Lxe�2茼`(���eˬc��])U�[p�q��W F�k��hKFt�xa8a�6�M-ͬ�˖���~���`�Ƈd�Cl+��s32�Ѯ�W�nd���u^XI�YO'��u�7��G��q�=�־�5�P��ݺvI�����#�e��:��X��]""��.���D5���ܛ�
�ܿV�r��DV�l I2�~ՙn(k�)s�Ⱦ��Fep]�V4v��(��];���0���z�Ѭ7h���moj�f��V���n��"]�K�xէI۱�Y`�"��,��7u[�!;���-��e��SW�����"���IX�\(ƷLWJ�]*�V�j�̖w�%'����W�t5��f5�͊�2��c	��mZj������&tS��JB�������{@���vt<�b��Qm��	���,KF��g��{W���b��m��9��V���6K��\�V��[ҚC�ػ�ִ�-�S��/�i�%oK��
�ފ\�ʴ]�B�=nطYz����N�4��uvpХ������%ӥٕ%g[�ԁ�b��V;T%ĹV��:S$��YۨhqY�禍��x�(=�@�U��NQ;4K��d�C&
*b:�VlZ0�r=�5�k���/��)�A��1�[�A�<������j��sx����ؿ�umk�S�=�l��n�:�9"�����%[
_K]�i���Ŕ�όoM���fY��5�
:��UL�&u��n��'4EZ����ŗ��XN����y���n���d)E���J`Ǚ�i\�.��4��hm^�U[�8c|�e,��i�c	"�D

l8[R�+,X�0�T$�F�4z�b�`���T%��ܼն��}H�����u�3��lqXf\|�\��uz+;Z����#j�7t����c%(hI�
�SP��fst���lK������IHⳛYNKz�x���b��sEf��,��2�"L�e]�{e8fT HVAk�[����(,�b�=ytoiL��>��D�)Xܭ��XÙ{�цD�GnL��Q5��v�PG�t�M��]�3���AmuN�8�q<�����P6�ӡ0]"�p���e�Y��7+r�;W5sc�8�2�*ݖ�j	iÇx;Zn�y	��]uk��8m]� ��6�` #ݳʌs��.��ﳊ�&���ù]��_pM�eY��kt�R<�d0�W��t͘�kl��	�!�ٷ�i͸ծ����}��2n�M��)�w��r��Xre�a�G���Ul��:]ܻ�U��\���&��UgL�6���N�h����/����y��s6��m��o/�J�gA���fo\������gUڶ�pΦ�<�s�CN*5��J}�h���S�s.���M��k�	�]�]8�����e��<L��Α��+p��q2Md��� *B�|��1�7bف2�E�Z���e�-}#g]ݼ%�J��a�U�B�+o/YH=�kn¹Z�
�(<��N,�}��nM9QfR:�1Wq�"��yˢ���u��Qˇw'n�ֶ��GR�%�K&�TRYV-��
� WY*�3�%��J�T��Q�s��u7���[&��l�Ү	�0�����(��b<e�����!b�/��cD���E���V�m �6-���.�D�f��U�53.��qC'*T�j�ט3T����-}��(6�.�\���&�^�w"`�i;��a�����45�L9,���Q�U:$�e��a��a2��w5�ߒ�۱�c4��me��P��2�m1���6���%عJYJ��R�cY��p�5� mk��A>ڴ��U�����гn�]}8ۉn Nbp*q����x�E݌S'\�.ގ�"7��G��u�0�ͼ�Z�&K0<x����e���(�u���|��M�n�$��A81���\���W
�冹����>�(�M��Y��}`��]�N�D[�uƎ価��C۸��X�4��Pg[�=[�`�$�T��%=�:���2�K� ���Di����5�)ލ��6Uv�X;/���ܝb�t(2Z��EV������Bn�Vb��4�����r�$O�fl����;Y��,�Yz4o+@7������WKv�)Y�t�PC�3���@����u״��3�b�99SbҲ������α�f�T��IтE���$E�ܷ����-�mP���{]+Z�ѻ���{��`[�����6�)"$\�2��I�>PV`�� I���r�ԇC��;PE쌓.T���p��򝛚�ռ���N�Z/�&�"R�q�e��ّ+BF[1�X��ݙ�Q���M\P4���Bg�? x �+'�C�ErM	"�D�;��|����� M??<�Q]r�(��G��Ɛ�an�g�u�wɷ7���bZMPƗ%�� AƕrMN�hmi'b&*� �k���8���XV��PmrMM��&%q��ő�tbm��Vh���K80[�f�X��ֆKe3�f�
������@w�Z���iWb�F�i���l1�M5�a���6��Ej�95%�f`b�Ye;PM�����h]2\3l�N�F�uM6�1�ف��.�	A��v���S&SWf�eWZ@#�/��Vo2��e��a��b�jgXXW����<�C.B'X���j\ݙYcu�F���/1�c���U�P\��v���8m�;VB��t[��.�F�c,�Jvq�����^y 	k����;)��A��	v҄��i�+3A������ڻ�Fh�lve2��֑3Z�JAZ�����nE+ѻ..�"����]<f]�k٩ue�u��U�qt�-h6�5[���f�La2�\T��i�vD��,����6�ESfD�.Mjm��֎l�K)3B4J��9�#6��V�J�mB��V,`;m�]XWH�u��"*:\�SWuk���]a�݁��Z�4b�&�1T��T�ke#n�sҪ�bn�&����`�W$]���Xy]2�\����H9Ys��WLq�@Ŵ�LH�	�hX�6`K2�n.`�f��XIv��u�9�m�f 'k��&5�D�5i�v���6�٭�]�8�� J�cضZ�t�u����W��ڐҦ�n)l��ǲ���6l����(Śi��u�m���#<�;^�1��[L.LTIM�J���ɘ�6�K�M�V�WM4�a��{B,�Q�ŕD���f�0�&�-��mk�L	�.�m�vv#M�
L֒��l�c1*��GY�(�ф+���V�^t����
k[-u�4�Zk��Bh�R]1����a�Ԍh�`�p�g0���.4{;Ul�ڴk��R��#)�3���l�#���6��A���\JJL�w8�T��\�hIjT+��É��2�m3k��hU9jb(iv*���J��+1m,0��aG����&ֻ%�š�mΡE2��z�f�դ��� ��iai�3�1vq.GK ��&���5�T�5���R�i�b���e�G]k5jb��o.!k�,�v-�M�bj�2��2�lд�`�y���ll���uK�E;Y�[g��ܛ%Yf��K$�P�نb�R���̠l��Ɔ�4΋BB0��Ib�jk4dmԙ��4@�QԡI�Xl�����Rn�\f�F4fѥm�u�m�&�c[V^��e-�f�����\ͦZ^�17R�.1L��蚖����i4�FԨ�ZmffX��on,��s�ZV\�n&"U6@հ�]��������,�H���M���lƌf�g���89�e��-�I�2�1m��kr�X��se�l�-M�=����ĖteC0�ij3
�u�V����b���e��x�F�7j���e��KN�rb�L֜r]�֮i���f�Ƌ.F!-�9��MF[*A�,���Jf�aڧXF����\�..1a�J[&�F٤��H+\lb�o/�p�ĺ�65�����]�Kh��5-`GKc�V�.�h]lhs��8�5��SD-"�a�ְ�5�P�1a�l�.�[��G@,f�f���^r��Z楖-�ƙ��Sb�j��X�*�Msb^&�]E��lB�Y���� H�S���bҔ�m˲�l�2��+X�Ȥf�����R�+Į�#5�ɼa��[D1lD36���p���1CM54ɳn��Xe%�+���A�$K�]�rMcLk5@Mn��w��D����,�*͵�`��fmq4��S�����V&e��%�й[[�.�y�f��y\��l��[�6�˘�Yp���C
ٻ[v�f�3[q@]YQF�JK�� N�[%��Q�i�Ҽ�s+�f�V˵J3��+�����	*n���n�ЀP��YD�Lݳb�L�e��[��M��f��W����m{bnm�R�0Ղ�oo1���]4��RM�B��G�k
�Z�Yp�f���
�ᦫ�s��k����`Jh:h�\@r�nŶ�D5��L�YfK�[^�e��`5\��۠�mhcCZ���]hgAΎ)	��%ˠ��e�ZV3L	e2���iG��3�o&[�٪�4b�ԥ1n�.�͖�3\�4dѤ�o�\�+�kh�Բ�B�q��.��@a��f���1���6�/f�(M�V�%��L�f�,�,6m��.[JG��� ��hFŚ8�̮q��
����9�;'�sS�����\V��og;�i�Q7;[*جMv�:�4r��tok�vخ�,˩.�����%tcv4m��D!`�f�LV�Ik��*g�R��n��\�V,�%p�ӍЖb'YEū3-f#����-K�TZmD�,�pl���;j��4�`�L�]*[�ךW]���M)a,%k5ĥ�݊+gn�$K,��!nses�*A`��f��M�f��9��m��{
�҂Yrض[�Bh�P�ְv
��c�#�Gc1Ț�Q�f����n���G3;#�s-Պ뉣��Ԭ`,,� &RZ���`��P�2�[p��L٪76�s��,�XJ]oP���,-�m60-Mi �aP��B�Im�J��c[��KA&�-�1�+s{�s�2RƓL�Y���(�����z�z�K\�H�K�d]"Ep��Rݱ+Q�5��Vִ���3����#"[+���ihUlבb��]��+Q
�e��N��Z�j�,,�s�� ,J"�2��FҶ7�`��$����q�Ř��ݨ��F�.�� �"y��Ř��MA�ṭE�e˩�n�Q��C�#�2�N�T�B�h���%.�jhYlֵkE�!P�$,.h,j�s�VEd���DԄ9c��Q�A���.�e��n����<BX�R3m	��0,�S6QfI��T �N�[�k.0��K7j�ꦐ]0.��T�3:"��[lV��V[I6��%/-G1Ck�V��ڭ�(@�`������a4�c8칩J��:�b�)4M�̬���]5��
~B��˛.U��E�MV2���B%��Y����L[V�H�j�f�[p�h�lY����5���u
�jͶ��O�Bx��<��V)n�N���te�bL+�z�m��.2fT�A�[)V*V6�F�j�X銱Z��;V�1/&�+q�m�e�����g�� ������u#�TFm��7#z�`T�af�,sie\�wΆ���4q��v�\�2��e4p;d��[�Z��MH֑�H��n.�qe�ƭ-��Cq�Y��NkHRïJ�Z]��0��TfԬ��m0aL�[�獞`ܡ]6�1n�:Y[�J��qB�3,3&J` �S-�E.�k��ӱ\�B��.���6�cf3v�����+B�!���e���͢ȤbXٶbK�׫�۝�%]��p̵��Mfb�,��qw$�v-�6�0cu�5��\D �pͳ��F�ͦѰ��v�����Py��]j���u�
�ID�:�H=E�%��X�teBR�⒘
T+2[ee[,�ȃJ�C%kq,k-	�@�Wh²��r�RT�`��E��Lں:�	6�p T1a�Ƴ8\Ҵ��rX;Q�uܘL��k4(�ƻG�6�mCe��JAK�b�YfX�Y�C5��(��l��mɥM�V=�"��!|��"h��\���a���ue�f4�])4{s� �5�%1�����j�n{m�����D�6U�h+��b�g	��R�)3v���ZĻ��f&2����L�v��v�-+DXU��mT�pҐ�e���`[��b�C0�W`�.e��wV]Z0@ٳ:\�61t�̸l4ΤԳqe�<�A�;�XJe���4�9#��R;��v�x1�;V�����^	�Snm͔�#m�VPn���i�+�X�<���ړL�fe�#˘:����,W3��&��!^#�)\h6Ҷ��������vڒX�hX�mq�*-���Xo<f-�3� �-ejV�Eh��M2E�ݠ9�4fic�h�-���K�����]4�B/.��U�m��f4ڤ��d���aK�,sk��Kb���7Ty��Ͷ5fpf8�2vCCG�e�����;vq�F���s��h]�eΪl.u�U-�bK���j�ݖ[R�U�s��0UٕF�UUU�Te®ʪ���������������������	ha�q�]���\m�A�3	+b��i�v�V���4���#�2ۆi�4�RVVZ�ڑ�Kљ�-��g]�nŁO^y��_)�4[1e�&!6 esuWSB�^F���Q���.�͕Յ�U_���X@��K>tU�%~<�74�*�t{ίӛc�h������c��F���[��ypϯ{��+��sU�����){;ۉ�<;��6���/��� ����A}�G�ϋn_�W""�Td�|j��wrǗ�W�sy��Ư7G�[��;xlk}wAS�o��;b��=��\\�ur����>'n�9�t���y���y$�z�:ww�a�>?=��qE�[`��L���nKSB׋a����dB�&�\���U�JB���e�p0�ͣ
���̴�ͭF�%Z�p:�YJ:򑣂mYi���.��"�:8ز�ᚊ��`M��]�vR�TA+lg2��Qa�g*k���o`2����
��6Q�J�V�Թ��vY4�3���ִ�lKc��PJP֦��b+ahRۣm�ka��4��[A��+m��$�l������e)���cn��crdv��n�,u�E$ڷ%-[i�� �[]�Z&NK�V+t�)f�=R�ln����`It��L�p��5WGg[���i�1��\��Ѓ�f�a&-)�Љ��h
�&�q[1U&�L��13i(Re��(V�	�6ڽ[m6JD��b.(/X��f4�]����me����6f`��V'mb0�5K2���p�Y���nvldcu��X��<��i��޷a��� ��=�����]P4GX�n�K6W��1,]�
khs�l�3�H��MK,�C-����75�j �B��j��F:1��ltpQ$%����jPM�(�V�i5t�f,B���5I��QA��0�"�fѣ��f��8X�X�V���5����g�	trGR�����!����Xu�R�6 ƚ�@��Ĭ.MGW��r0��Il`����!coU�h�m���al�,�j��`�X�t��	�F�m](f]��&��YI��,�J��)�7@��GdkP��F�3��a�le��Ņ�G1��o��%e�,,�!*��&Cf�W:2c-ƶ���&��Zi�K3]h3lb�:�%��тe٣Jk����\��Z��]�������e���-�V9�mH+�U�1�@YLUӧwgP�
����-���9��X�*B��*$FXP��ז�x��ba5i-�,oS��e"�l��%�[T�h���V����[j�@�j�d�m�%�Yh�c�"Fշ�����-j-��iA�Ye���5i+��#E�jW��|�_Ԩ���͠���գWF]SH.2��+��)B�Q�J��4����=��Ӱ �9��UZ���Y��0F�
���mlu�<^��6�6�A-ǔ=�W`�GWL���3S\ܼ�.q�r�A�A�fͼį���*�H!���@D܉��p29���!��{�[��ܯJ�8�D6��iy�[�E����"�����A s��mHɼ�3o��-���/ #�˅��Z��=p��"s� ���A Cn���h�A,5'9r�r��p�p�@��[h��D�m��
cf1��!�R�[-I+�V�U̵^���2�����V@Df��[�Cp	��1�Wc�w+ҧ�D�����'-(dcA���^n(�m�#�S�M9�y��>T>U�-�����-�53k~;r�u8;��#X�k+����G>�����|v�WdP��ent�o�N�R2r�������5��7�ۀ�A��"Kq�::�����w2	�M��܉�p�8��ΰ�ަ��y�p[Q���^�h"� A-� ��38},1���rP/�=�����PB{��\�+�^���{ax�d�<�m����	���p�ڟm[���&m�����>���r{�A(p�A^ ��[�/Б�7|Å����S$����cec.UlbW@k��Zj^� �+c��Ur����=]s�D6�|Ch%f�O�r^v\�p��_P؋3�����Ax�B ���v �"-���s�sk��H9�*Ov����w+�3�A�� cA��]��/<�<�9q�y���mp��Y�f7�Z"�]�ݜ�p�[�eN��'���@fÝfuEg$��vn���/#u���W�����˙�;W��;X�F��&�Gk^n=`6�6�תc�N8��A��s�A �ܗ�w&�e�mG_j�D�s;nГ' �l#�Ƥ��/� Cmy��r����=�.g�/[�����H ��,h mϧŴ%���o�K>�{ ����:�f������c-��l@b�fGx�SRFlp��jBu�.���|7o'�HY%��(�A��ȓ�<�
!�3������T�Go/H�Az,ܜ�};�N��p�&�T�s���2c����^��׵��mϛ�X�{�;C�����uW2�(q�A��Cmy�[�Q̓/����T.ן@���ŗ�{<;N�L�;Ʈ�
?]
Z&�4S(�ȶui���<s3ۛY^�T�d���æ��n�|��U��5���(�f�L���t8ӏ!ڂ!�����!���+'��Ju��nU;�%� �j�G8����lĊݨ��e?Y�s�b�kY��B�Ѯh�b�L��⩢3!����2���;Cݑ%���Ƃ$uv�w9����L�W{��ct�����������q���:-��[/����vꕆ�/�nxs;��o��	 �
dl���a� �Nd�[Aۑ>n����qQ���S��\8��R sA��my�t��ȡ��@D5�'������E�vsSs+ҧ��^"�s�vg��@uV���^n=@�Ԑ�[��w���0����7;#�����o Kp �r'ŸD�V�n�p��23s[h�l��H�}ZT����BW|�.��Yu��=v��t�+x!�����o�^�?/��X�䣙v4����(9�11z�ߌ��uC�҈/&0�]�R�0�5�	�qn���S,&�r$V��mI��(�s��08)k���9��w\��xfp��V5Q�d�\�i��45�f5 ^Z(�]\n��뙭�#@���9X�V�6XjG]a����"n$.��(�a�c:���,5�ʱ~}�_�7�IZ[��%���B7jX��kL�`�ՆPP�:T���d Az�!�3���A]�e�w}$�q���',�\�1��/��-� ��� .��p�b�cӗ���I4:�K}}�jezT�{�u���:��x�u܆A����_�p����yl����sn:z2��� � />s���-������3i}���ER��CI�[s.��]���%Î>��׵�V���K�����$6�>-�@��܉-���Q���&GA��Z��T�zT�A��ւ!��!��7
���`�e7M���n�G�Y�bl���L��b :��˙r��، ����-� �mJ����g�C��b7�Ȅ�-�\�`z�D��@m ۹��'Js��e�
�X�M���
T���	�<���	�"#,�f�cT�R�����+��ll�*ʏ&��Mt^]�Ϸ�K��ϳ��A'Z�}�q��ܤ����,�{J:lO�_)�����$����1Y��`���"���kmMLǢe{\ph"s���m[�X�iN�V=�ju` �-��[jB��v�zU����o An ��We����� F��6�H%�@�@6��ڭ��� e�����U�Y95�I�q��RA��n �ڧ�&C��[�c�6LD�&DLK����B��*�R��-U�b-�L����{���ײ'Ÿ�m�"#���E�J�D�H���vb�ݐwt����D��꺇�*��h3��^j��v;������o�� A�r'Ÿ�	�C�Dv������y�@���|�U�c XOi9{]pCY�׆/!�FY=��H�<�Vֱ��ۅ-y��<jV�hn�f��.'�����z�T���XyyR���q�;W����"j�א{{4u�1z2��v���� �l��,[AUW�6�3V�R��3�}��\ء�/$�!�!�L��h"�"-�$כ��dݰf����v���7�[��oy[��;�D�� Am׮XYg���=0La�*}�$D��PB�%�6�B���T���ۭH�r�\�!����/o��ۙ�m��,.�ȼ��$�\w��vAʮ��ҰA��A�@�[jA�/7&s��.`m�����#5��G�Ӽ�T��L�� G8ۧ�"NnU�S�ۄ}�T�h/�6��	hި�ބi;�GZݝ�b7���D��In<�@6��4ĳ��if���s@s��BU+ș�ˬ�}�dp ��RE�q��TȪ��<i��1 �\<MM8�b�=�c�qي���t�~	wM�ӹ����VO�:�� 1�p��J�6�m�z2�E�C�t A����� A�nD��
5f<�ɋ�`�A�DD:6��#71���A{�s��mȟ����A���R�L��)28&P���.�
�m�)�.�ؿR�z�I5p�Ŷ�QW��w�bݝ�cW/��A�H�{c�6�mߤ�"2�MQj �k�A
�9���2���	���	��$��-Ɖ]��܏Q��>#�/v�^ ��O�q��t�����QGs�hSs�Sސ|^Ǘ4!�>���Օ�'b�n/h���9��A-�}�k��Sջj���@Dc[Y����6�iy���Cnd�y�D6�-�!��{T������m�^ff�; ����[�k�H�����!Zݺ��Eh�]u ���kn3��3m�Smጱ.đ�͉E�
�m�U8�;Xn���$u62N��30�2P
-�\MX��t��m�:ZU�� :�`a���Q�9L�B+�jg�2����an̹I�ks�[��ZԬ��qb�� �b\� �Z��
�-���R�	�R��y� �Uًi�c�jl#v����(�٫�2�l���ˮ��f��ks�mHL�T����)��;ܔ؏f��{��9ιvG3 Ь���]��4lÎZX�Ў�!�TI32�X9�@���W��Xl��b�:�z���x��(Nx�;R�V^ǰ�!��m[�%���6�,�&� �j��Zצ��9=[��o	쀈#uȐ[����,��� W ���d��~�6�Tr��WI���˼�qaǸ�� @ւ�n �ڒ^Bi1n$�C�����;� ���6���"'Y�¦�#Ч���"/��U�H/Ot]�!�H�ڂ-��^��@�"1"v�v)��=���9f��b7���ք��!�}��?�{��\K��X�䫚���0u���+�
��) �ɝ�����K/籖Y���k�A�9�}��y���.�=�1��bi*�v���y�^n� �+��}�L�1I�c�������X6\ž�����Yؔhޖ&5�%��g2nz/549�k��r�0�<�Ō:���t"*�V�7W��U�K��/�FT@�(p=��<�@�ۓ�H��̖�6���@�j|Cpn m�	�3SX�;7��5n����d�а[�AmmȑY6��  �Z�ݑ>n=J��_,˾z�;A�}�|F�����gۺ���p�>n&)bU��sC�	=;��ʈ��{c�����B�b�wϡ��y�u���cK�
hM�.p�&�����n{K�):B��M�25�y��n�Ԛ��u���صk���;Cs���ѹAU܉=Ј-�1��An�s�]#9Rp/�7�'�w ��θ��}�N��缧�k��qp^P1�DW�R���']�l!��53*�fQ���)��2�ϙ���^X�W�Y�t��:c\X�2��f�[�K�6}��Y�^���㭑��v��D�Z)Ec#�;'KYAn`,�eҾ༼]�9�z����͉�ql-���z�5)Q�,�B���/Z����"u�3I����2�ǀ܉,'��.���/�'.�L�ۜ�-t֞PG����,�R��ܬ;�*&	F^�����6���;{�\���!��T�۴efɍ�;z�U��nLl��	�o%�s\]���1���wp�if�]cj�1d�6�m�B�[��p��U�Y>}[Ye�^�籅4Y�H��k+0<�[���[�i`"�1��ٗ�dƞnh�	��ˮ�{�R˩��;$��r��"j��"�u��F=-��6�)f`�;�ku蔈�5�`9;�s����$,�:j�AiTA�W{�W/�G�O��ᮠ��,RY��>�,s3��㣕
�3�x�;%ofS��SP)-�il�3��D��U��wkm-����S�%���X��#�ږe�5b�(J�ZI���mLNжF�����w��r��i����V�5ЦzGw�P�0Wn�VT켾:�ir����������xL�/z=�X���-GnQ�ؼA}���f�ٝw��v�%���a�&vD�y�5�뼤�\\C��"�{�1=���{�Yɫ��u%5l�zR����`�2�iH�EN�R��@�-�d@�$�7�5�!��T,��w[\�y8�͸[���6�Ρ;�#{^BJ�A:F��){�͒&X����o�oIj���RS�)zZYS� a�:d��	�6LC���Ĕ��81:}l�����|�7.n�#��L(��5�rK��2�>�}|�����tF�c��
�v������|yF�HE-��E��B�M�R�b���}es��C��
z}�y��|F���vv����Ʈ1Ii5sa6Ԛ��OO��ײ�ƈ�H���D,f�:~��'rEM�q� �A�ݡ>݄;� Cmtڲ���
e�����u��%��N�)h"�/6׺�xo_=}�}OE��E�KrD�8:\2��p)��v����E�)�U��?O>�7�~�=���MYhe���Wz���ʹIi�&.�:��N��F����q�mzm���.��(мA�B���5ױ���ƈ�@�pZ�qu�X��ޜ*�Z� "3�{\z�h"r'ŴA����X&��.�i�9�	�� �5��nŶ����;���1�<�Z�$k�$��CpI���Ѽ7�C��
xO��x#�6Uњ���P$(G�9��j�V�f�.�ref7rf�Z�KT'�/�!M��쫣������A4�9zu1��	�AQ����^�����Neq̽3  8�蜃�P���8�~�5����0\5�#��ᘃ]�Q��	�����)����&֌�m��0�K#�qȏ:�{kVLL�N��H ���9mϧ�6�J��)_s��v-��ns7�Z1���n �ڐCq��G�d��;��"�R5�h��!�@�= ��΁^!�&�*ʜ����Ϲ� |�) ���n m�!b];�w�]}�'e�cհ8��In!��6����	ŊK��9P����ψmjh���p�N����|}p�x��Q"��Ǒ��>!���pm-���ɴ F��ܤ�v%��xw�pD)��t/Frۑ>-�<�(���V+zuo�]dRKg:��W�%��WFhC��xvw_E9⧥F'���闹D��wg%��g����x�	���4�.+6�Ut)4�R�Mvb;b1�%-\����F�:�6����9[p[�,��Z�l&i��
,�]��g�|���\�k��$rKGKGZ�+h!m�Q��01��K�]JV��6R-��`W���15�.��&�%�6�:�������G���X����/P4fK��-#ĺir��v�.쟯��-�~�]�lS`�A��pZ�fTkz�wZ�,=qv���,��Y�q�mI���v�����q�;�ޞ�Q�|N�T��+�$��&-�w���ں�=��VCLOg2�V���y�`6u�� ���){v���f,��g���'dJ�>�s��^����L��!,��09ϪHkRV�ϙ�rN�}��M՘}��������$5R�G�c��6�[�]��q��I�y�]�}S�v	I
z���XQ8�l\f;lL�bѲ�eq1�����ft��C�+�f �y��d�c�[��FS���gd ӷ��m�Lu^�����!�Oʄ��泂h
�8k�X��.��yLg�[��ى,�M�P�x��wZsMܾ1U�-u�4�:(�,��-���i�_���{�{�տ�ߐ��/���?Wbp^��`��� c 6ϋ���Wp�IT�]~�gӕ�'��<v�ɧ|�߾���l
��}ٽ޿���*+ʱoFdy#1�.��\')�S�oCh����*�G�d�� ��9wq�or���ڇu��랩�H4��M�AU';�c�{���,�}��Ь�pV���QN3-�V����v�أ�FÙNjѾI�"�P�������]�}Z�I���򪥳rHdUH�s�����\�c�Z���9NR��+�Hfs����סA&��H$�q5����2y���Ru)�F��Z��P"���o����&G\����+5�n┹�;��\��{��DN�1�RjP'��xx{�_oO����/U<����xf@�$�2���X���m|�9��A�P�c{1�ۍ&�ٽy[΅b�I����ʐ}���%��ڱ��]���̝�zϫ5n��������O{n�'��I�* <�[&�:ƴ֤��.7��b��F�ZB.��g���C���RO&��m�v�] ��	�\.�d�e�y�� h	>�����u<�o���4
��ր|< fǀ��ݣ��mv�i� # ����v���R%�s(�q:�5���\���D큽n����
��@/34�������13(ku����3��£-.��#��s��4���G�����X%�̰4�I2�. ����N��vq�;e�>f!�� P>��^ Oջ����:�W}V�<�ȉ�edD���Y��>�	��	"W��R{[�t�97�R�;#e�m�#�dn�����!�ub��˘����V��TN��Ǯ;��R�Ɵ���3W͢y�B�	"f��fXh"$e#lD̠K"9��39�����;����G�r7�|�<���5�����D�<ݠwH�|<� �m� !��K��0�ȁ�m�(X��a�u�b񰶹aZ�=�Lf*�Ғ鈶�2����a!�؉���M@s)"e ^�8��^y��f���qa���<k�4u��z�zb$9��,���X�e(�DH�32�󾫞���W���z�,��;9x;[����KYu� ����!�P7#���C��h�J���� ι�H]�7#�`�Ds2��!2�9�κ��㳺�c�Af�W�Gv���?x���w� fPDH@��@�����כ��� �aGx	���L�t��yHX@I2�,��s^J�<�l��3[@ָ��$~R6DNg�n�Ȏ�ݢ���ȁ�H6@32��D�e���s^h���^ O]�'{����G Lx|D3��$��H���R�HD�  �Dc��f����1�cV�YM����]��wՆ���˫b��%fKK������	��v�q&��}��$���[���u�*��X�XX��h���nv+�kR�J	���&L҇K�79,[�Z3f��l۫P����:��-�s�eм�%��K�ٹ�5"R�Ҍu�+�d�\Xi���k�G��L	V�����P{3j��ю������в�X�Vh9�c�j�e��
���f�V��� �6[}����Q#�GiQ�Ɓ#�c1���2Й��ai��m�j�����a�D_9�l���,�9�~��� �>ݣ�?>���� ��>]�;�����n��"C2�;�^ fe�i���HD3(��VV��q�}"i���!lA� �F���Vxy���k8��Š�#��7�	dG3,���;�n��;D�.�. u� ��僢"L�:�E�6� WP/��ؘ�̟����G��7#�؉3��&�9���HD̠"fXh���x�f��<�
�����@9���"Be 躌��)v}��Z~�x}� }���s�rk��V�lD���@� ̤�fP6�Hff�4@qǀ�/j��A�ʀ c#���9���Z��dD� �t��N�@�6�O����N�4��7# ��o�����0�8�E�JB51I]�4;V��1�Xx��W�m���w݃��3v�dG �� k�	׸�~�}��{��z�y�\o�;8�:�B���"u�6��]�D� � fe����I����x���~_���p]�nÏj꧙Í��0�Cp?�̬ݫ��g1y{K�h��0��R�f�|�m�]�c�Q%e�m�_��x{�| �x 3iЮx���|K�N�73W��WA�"B�n��D�D�#�@Ww�7��:��Mu�@� 7����q��M�B�$��@�;�7[�s+�N��Z��������w�F�$�v	a��LA̡2��"MhÞ|�4]��k�,DN<��)�6� �{ow����a;�� 5 |��"�@�3Z�3�:�D����=�@32�u ̤m��2�-"9�`N��7�w�"t�/t�ewϗ�o���~lʾ�h]؉ w�DO��<��ǀ�� U�Y@e����O<�yM�l�.r�k����L�3b����e�ƥֵ֤w� 7t�D5��$s}�D2�n&e k�|�y{7����Ox3H�|<+��/��>��p8���"N�����$�@���Aq@32��0�ך�������� #�=x׀������`�w��:��w@�<�-D2�羸�!<ާE`',M�. g��h����@����fX"`����;��
_��m��}���S%昽�CV&D֫�2���?bn�a�S0i�Џ����pu������C2��ʋ���  x}�WԒ��עWA��H;݃��:��,"9��032�4��������nbq@��I��H� ;�!d�3(�u5�;�ٽ͜_}kh�"$ �;��]W�q��8���.�w� [3)��h����G����b4�go1(=���)�h7�{�+g��q��Y�w���w�t�Y癤M0����9��L�֩�c+�"2����0D)�H%
�l�3�e�JZ�i��.����ɝ�������$�z:w޽8����fX"$��H_u}y�p�~��������V���\���݃����D�#��D̴@���!�@�9��3�g�Å?d���� 
����||3` a�s��s���/���k��H�7�#qu�@32��g&u{��"@�T�q���� ��:��2�.#�@\D�̴٭��<�7W����wy�w�sA�+�� �����HrD� � fe��&y�\�y����D��X%�|��t�̤
㎺ם����fV��9��@7��>���'�7�(?g����:fGr�L����.�k��%j�V�<0׸�m��"�D�E�*���DCr"�o���� ;ՈzR/�}�h��#̠m����"j�HM�U7S�NUN��� #n�����j���D�}�6DI���9�`h"$��H�������{���v~0h���%%�Э��ܹ�9�A��H\��Wm�:I|�����q�`舓7be��|@m� $}����}#Zu�� ��6DK�Y{���]!]P9#��H� =�H��̠"fXh�� � w����L�5�7f�@:�vq@{  ��f隿��gW� Z�>����~X:"$;�D�#�@rd�s�.��(3\�@<��"D�y�qff�4@s)`$bfP��
�H��9���W�[_x*׀�<;����%�̴]3)�d ���_�VkB�r[� �����L��-���dD�̴>gxw�x�ի+W� |G���< Ǫ���q���� �C	"y� Y32��G��3,�#�����������<$�� !3y������vu}�7A���~X:����K��P  6׼u�}Y_���י��a]�5;6N^,o�h[	�@������=RV ;6_)�����G-1,�A�Y�E-ɓo,���6�.��	���� 1�$�o�J�����fG��̼6S�J�[��2��S%d��:�nG��p|�����,���VsJU�h�m�͛OF�pb�4ц]�-lF)LS�,�ܔ7��K+l�vv�Q�׎�d����,-[&��y��t��)Y[�;��Ĥ�:�F�3�_wA&���s�c,�h�yD���o[�I�G0Sƨ�[$��p�{4�Cu֕ �!�c��ƍ�������rR�W��c�6�I��7�
9hecVA���z��͹ע��W���U��yb��CA�x@O����!��j���'_:�I��Ie̓{�J�g[��)�m�v��+|U{Z
#����r��K
(N�b��\��׹�]8�:�&�����V�b��Yk�0�u����[�D�'V�	�%��$�Ͷ2�C!n��_a�}��S���ëM��9'"���']���5}Sh\���U�ru�y�����|�SIn�9]x�8�h+�����=|t�O=���F�ꨕ���V��3u����UnYW�-LK%]^�����1�L�4��q�\�+�EU�z�p�%*���Fd)�Q��&�z���ֲ~hK�?��@��>�-�?��G鹜��}f�$��\7�����J2��\/~��ɞ���]v�d�wA�Ԕ�lص�B�� R��hu �)z��^�p,�K�JL˜���Mw]�뻀E�{�L����9̑�}�/]�w2����@l���:�8��bk�����>:�n	�L�}7}\���:9č;�hE�~�&�k�z\�3	7��qM� ۫��>�'����hؙ�&�G9����Q�a,Ҷ��nt��ٱAGuLF0�pe�;�)Ԍ"�z���h��.�\8�d��f]3T�eT[k-.�y���Hk]��j,&�ÔM��qu4j�5�sui�U�ڄ���NctT�[Sce�4�ST-��7
\Gi�Q܆#ux�2F��̶�٢�J�H1�m,@̱l)nKd�jc���661�D�j�
C6l�5�Ԕ%\afA�eܷ)Թ?�i|�W�X��?�-�#�Q�hLv+#�2��ۂ��ֹ��b�16nh9x���WF��ԉ(c�LI�f�I�r]&e�`i4ҏ;f�c�u�1YW+��2Bk�Z�0�u)c��[��ܓ^Y��4�X��຦�P�c1iol�XY�Ya�-��)%n��jmn�����kF�WՄ3,� ˬ#,�k����ɗ]��YA��b��.��C@Ք�W�m���7W��bu��Wb"�k1΄��1a`�m�7$Mp�Y*��K�h�-�A��Vi,vu��K5�#jDm�e`7L������#ft!k��h2�l�uT���y����B9��n^¥\�*Ji��ZM�vbYr��,k)-G<�v���jL��p�Ehg#v��^��M��]�8�c��4+D�9B�08�KȑWh�N�4��9y�u3l4��&��ȻG^�:)J�3�H�@��.ΤwXӫ��P�3�yԹr���R��y�:�P&�M��U�EԵ���n3R��7T���wkH��	S,m6!anC���c[0�T��f�wia��+2��Zʽ��,v�u8�,���כ�Z��R3j���-��c���r�kL�V�vUUUW`�a��璷x��V-0��(k���FS4�.��#7�	�.	^�,݆��jǈb*��gZ�	�MiIt\ZL�V��j�b��Hۋ,�ͷ:[�4����/$Qn)vnŋ�͞�CJM�*F:�;�P�4ƺ�� d9����!\�4��:�
P���&���GF�#Y�����]t��¬F2�a*�F��ё���Ŕ�qY�)C8
�bֲ��(#*Sߟg��h��\B��My�Yl�Q�5ڏX�4r�B�����I?m��D�ￗ��w�~����P�$L� �:����*����/h���D諪�����<���@��|�,D�3(8�����%o����Y���,��Ȟ��5�[��4oږ�l� E@�C��6DO;�D�̤7�N��u���qw���2�ȁ�\�j"F�t��N��̰9"$`fRk�=�g�f���}���������H�yh��3(��h e�N��/�l��9���M@w�B�	��|:�5�/u|��Y{@��a�� �Fȉ���Y�'@�b:��LD�;��".fZ��D��ez�י���Ծ���&�;�^ H���|8p�d�k� ��>>�s�ȉ;�"j�HYs( tЈv����A��BR��&�eAK�wkr��֌,6B0��F�8��_�I���ӡē��#lD�y`���LD��@���n�6���� � }����{����6yb�R/:����|<>2 ���S��>IS�Վ�Fe��	d.ޒf	�YC���m��4Fmk�K'v��DF�A%��C>�����֬F��:��<��+�������l"u� �.Ny��~��޹ٮ������D�}P�o;�K"=u@N��^����i� q��̠m���D�#�T�D����:�y\y�;냱w�h��N/�&��{�d]���X>�j���>�Ĥ޳U��mj��#=~]�zVT̕p�*��|���n���E��9pN�o���p�iG{�=[�'���l�����;��:�F*�W)$�f[eˮ�����$" �D�����a��.��$p�-���c6}]���!'���[��6Wq��h�â���jC�[��D}[���J���Vh�B�`�l6V��F�\pFNZ�����W�ƦE�'�_^�����vE ��Z%� �[��V�{Bv��e���Gd�;u���ܖ�ſ� x{�$����o�'�8ҏ�뭑wc��u��^�/7�� �U6&V�������ǖ}���	�{y���*�M�lS{�*�t*AY�W�C�9���(z��6)1�~��G��ѵ=W� ̪�F���J�\Y�l�δ�$tsR%�*kvÏ��|ǿ��G�FI���o�g	ƒ�&on/;�f�l|���^��K~Ş��^^�-�m�YU5&x�����]ڝ��¯)��LSb���\�
^��8�]�sӨ.�k����m���f\�� ���r;��W|*�K�t{fz�mݓ(��'���ⴡ}p�đ�Mk�3f��x�\d�S���Kx��[r^.��g.3g���Y24H̓/pۥ:j���{� Gߪ���m�[��5��G� Y�w��X��h��79Nx���ڰ)���h�u(�(�l�$9�"���e�4),˫����ӛ��#]-j�������q�f-��ٚ�����_��;����#��N��5m%�Ώm���b�7!�3��=w�<.�x����)�51�先��}�WkyT�l}�+�\/t<��
�X�f�v��s6�[úA��GHy s����]�������P��V!T���}�yA��%w��b��7=�ك���٣/ph�=kc;d�"�p�@�Cq
;Ǖ���w"ڍk�g��p�Ҟe���?����L-����E͹&������HKV&�,�]���e嚖Y��	�#XL2��r�5�c(h�)�̺#G�Xu�3�乥��I�BY���"�`P-$c�]M�4�K)��O�3��%,�¢[V�]t��pd�6Bщ���n��e����T�vճSj�II�������h�ƃ�6����a?;���u���#:�F�XJ@�;[4qtk�2@S �)�R
��T�;�w~��sqh�~�z�$�
=ϲ�O;���Tئ�Sb�h�P����
�����Z�{}Er6�������V��h����Tb�6>��X��.ǘI��z/gp��_@ww"�.�'��A��G#��<��7G͊�e�����1$�=U������#�`�pl}M��ܗ�t+4�#6;��������l7���'��d
� "M
�k,-���.����Vыue�P��s�2\��AM��d���7����T$��fɒ���^�}���o>n5|�ׁ��n�Wo��g�@;'�Aq#eL�W��\7[Y��=������k9���)�%��mҦ[��rہ(O?�� C��F��w�؜_���USFx��p.þ3]8
�'�ww"��N�(v^�r�,c���ŚB�T�lSm�cjJNZ��Nj�=� kz:�S�|�eՒ}_?��c��řc�S��v��Sb���c��ɻ�ɛɾ=U51�[�c��S~�^<���([�^U�U�Ķ�.�6��Ja�clM�ee����}>{���עSb���+"���k4��[���w{�Z>l6>�����VK"��>���N�w�-H��-��L�Iu|1
�p��c���m���ʽ��gV3�23|�/�]�S`�y7grzN�[�:�#�{��ev,�x�������͡0
��_�2:N�_GEMML|.hl|�l^�����}��=��M������o���������gsP�_D+�6>l|�o�ukp�>+s��{˗$I�S�Z)�M�wݕ�0��3��׌ͰK�sCn(��bg!q�\6�.�բ�b�\�ϛ������+4{ύ��+���y�K�N���w
�	�lSq���J����}���H��o���ת��m[���_h!Ϟ���ϛ����{����圈>�����m���<3p���U6{	y�ޜm{X=U'xڡ^3�PO��_���I`���u�z��\����Fj�����oF�=9����T#�kDE�E6�J�d��-ﰩE������< �����G���q��3����T�p^�@A�}��Qe����Ͽ?=�l�/��~�yj�.�3.�&iIul���#,(v̬���!D�30�5�l��w"�=;:��`:�s=�}�Ւ��u���p��c��w�`�s�үA^���x7��V/c��R
�hn��=���X��6>n=i����(g���Z��o)����X�E���G�mg��}��9}U�+�7Ԏ�Ø��Sb�l�� �ϧ�x|	`�T�Y�c0z��U�o*��]<���?c@���Ci�.��ʄ9�p"!Ƴv.���&�fJD�:ƺh٩5;�(p�z�:�}}ڵm�EQ����)ހ0 A��I(�`�f�[IA�V�u�*`�[�����]c�+n�4eZ#�Xˊ�m�]��*b̮�f�GR+�i��f�C[��ѳ]0����X��iE6�Cpf�Gmh7*K]	�m�:�8*��5�[�z��ܨ f�T���b��k�*E
��
�t��%,V֚�v(�X��v�Ņ�4޾_��袯Ҙi�������ڤ�3ͦk2�U��G0�8	�?R��hl|�y3�(yk��[����Â�;{��m����X��")kul0�m���.�.�����CG���������u�r�b�����et�L�y s�]�����߻X<�>������ٲ�r���!���YՐǔ���͊l}v��Ή4�Frc�9��b�]L.{��Zz�|H����x�_y������QP�� �](
&�Mq#yW@a4h�s37Y�`��Sb�#:���un3�;y��0G�N�l7wx��]�fr���Jwb��!A*B��|��vi�f��+���Z�)�--5;�`ċ]�]7t2�v뤦&.�� ��9��𼹏�I]U��G"�=�R���-�~�������b�lSb�����H�����3�WgmsQ}U8R��a������[u�w��B5D��c��+���/뎂��Ԋ�W����͊mF�G������r����nL�=^�T���͚�"�b�@�[k�^�ֆ�^�$9��3IK�V�c%�4�`,\�bߪ���lW͘V-�[����v<8s����\>��b��]�u�*��.�=\��^�0f8=��Cvz�v�*�V�l�q�w����=+�*T�m����*ʼ,D��̴ƚ9����x�P�W��J�J��U�]�v�1*�b�\-L��8Goa1{DK"��F�u��Ÿ;jD�M�r^ܷf���Zwq傎��`�;k���Yǈ�����i�]��V�Cm�/BRR��ث��N�Y��^ݠ��Ǻ��ˣy�X��k~�+��#@t�}>u;����GzʡB��[5wW��F�ܷyt�8��Y�d�.h��W��v���Cՠ}��U輧:%�e�=dg�h+mgν��n�Rle�2���dNC���J�N� ���脾"�J?��Wn��p��7M�+s6��uuc�vu2f�ö`�t�l+�ʆ�M.�e�,-�$��y�����YwXnY�gM8���\ҷ�>2n������ܭ�Q�D�kK�$����f���]���w�V79�6�x%���;���Su��j�[�K����2��6���	v���-�o��7�)�=�Ń��e��r�E)��&�u�M�U���Tœ%��L�Iu�^_^^.��3(��/Ty2�
qp�:(�Y@���:�5����NŪ��;]��[���Z�g5�ܚ�G3��#�|&i��	�=��Ȱ*r�S<�k����۵�e>ԑNѢ7gQ�LU�����&�4˩�_��E�}ר���:���߯/;$|��J�� �"��f_���v$�;����4�U�-�,��YBP�p|8�9D�˝�\�/.s�Q�d�nu�r�w�뻴SΨ2��v��z�z�3�n|n&��ouq��1%�z	m����Xf2�����磝e"ܷ(��n[��uɗt[��u��{�P�h�r�9̔�"7,���KCK7"����hĆ�Q�� �UtW�q`�wV��b��ԕ`�>wMK�c>�V�W���".���'T������m�� ���y�C����B�m{�zmo8�}���me^o��|�6+��6)���]�;�i�C�5ܮ�2������;Lc�c��u@��#""B�fDF�lY�8ڱ�-+�.{P4c�&�A���v�߹ߘ���z�N��Ǯ;Y�I��&bm����[_n���q��ٮ��P�G��U,gi�u�#�}<>�� ;Ѯ��y��Z�B�M���k�f�y�č��dz���=Rh���a��x�h��v���Y���G���Hrת��$Pl9s�nE&Y�2��m]�%�r�-\K�rd������yAvQ�C�e7c3�-o�/�n޸�h+�Y��P.`�����:/~�ߡ�_6>��ͿW�=?��Q�y�6~�	�^\��q�p.���J�L�z����7#)1r�m��E�4nu���e^k�ڰ�[�ٕ���]6*��[\�xA�=//=^��k"�}�r��)��b���R`��B�fj/���1�wZ��k�i�>y簜k�ww"�S��;�[O8�k�ݯ��k����+�o�խW������B;Mr�A}^w�}�8*��"����]͏]������0:|ŀ�zo�ݭǪ�q�U{�����rghm`B{��^,�3Q�����V5�T�:�t��7�s�W����!$�ɉ�a�c#v�͛��~��7���A�J�k��ML1̣�Ba�� f�h�꬙�,˥��iV�1Y��
�x5k^z��r�s��!l�q���+��&�jVZg�)�ۙv�H`����f�⥹v:��vu�I�����L��b[5kkG+���I�J�jv1���V�ivx)d��& Z�.M(�X��v�гFZ�w��O���Ю6��u���N��;�]�va��ZDB �RJ��1���:�z�iT�����{A,�W5wcԴ>6�}M��c��l��pL8u�^�:�����ܘ G+�힜���ъ����V[��4@Nt��/7�1��h��c��cZ�c��uRb�p��L)<�;��\��3�o*�w�$�^S v��66hgǫ�[j�k	�g��+�|���+��7��6h�Z۩��P�*�>�D�����&%-�Mk�"I�,)�:�����M���d��^i�޸�W�a����~^V.g}�cx|�y�kk�4Z�:���oU����X`���">|���n��K��h��&���ߦ�aɁ�عN��e�b?� �_z�~���߯���wG���}�S~�'��Ҷ���ݕM�l|�]���d�����ܥz�+z��U{Cc�l6>��cν���U�!U�Sc3��Vc��y�]���@/y�z�
~�
��͏��M�b�<�
Ǐ^J�{N��&�n�l�[}��d�bԙc�"�"�#en�@��J�[4ѩD�F�*fei`K�^�Ϯ��[&�˶�� G�]�l�5X����c��M
-��A�y�����9�����F�Ü�m��%��O�� ]���͍N���jM�k&��Z��X�|.K+�ʷ���_���|��\��c���+e�iԋ��:�7"�k� g>����8׷��:���6H&t�g����c硱^%R�\}�<�z���9�u'�bo
l}M��l
�
nK�������נ��9���]Ǯ�<�G�C�q�!L���B��%&tT�뢹ubSi]6ʩ�i.�<,vr��������|ف<]��h�Ӷ'���K�G�����M��6���t��C�b�T�ޫ��rs�����s����1{;"wA��M��6>o�����=IWl��)��\#\8qw ]Ǯ�5M�Z<;:�E6+;��램:v���7�%n��ΡӮ۱�"ݕz�N̩E��٪��1ɅUtsU6�M�'���n��=T�&gf�W*�ќ__U}z{ϛ��6߸~Ӎ#���機�I�@�z�W�Sa�Щ,��Uz�P�%�i2�,��M�xe3��I�n5�f�6(�GG*d<��z�.�Bꇚ�f��.�~/�����ϩ��lV�i��Ý�M��\�|3���mö<�<.�]yj�@����͆��2��MwG��&��3ò=��z���4��.\��w�Sc(��Ë}~�U{��!Q�~~�pD�p��|ئ�Mc6���=M�Ν�����޶��vø��z�s�$�z��!��P��9�RV����ܖ,v���B��Q�<�Lɖo��i+zT���R�n.�NGn��uް��Q3뒄�h�����X�f��%+0h� 0�,���n�3.5̤B�+څ���*��5"���ͳ[�]6���LPr\�cR��h鱌r�̬v�)�Z�����k�Z֌s�#�R���@h��]mue��n]���7#v��m!�;QKx	�ei-����i�-X���>��������QG*<Z�B�v��L�*m��@�$�~/3ew���>l|�XN��?6x0�{�3�y*���C�?
l|�y������m���}[�/B��aK�^}�W�k��C�䫐��6>lP����Jw��6iL��3���ew�E(6ޮ1-O~6j����7^����f>7k�|xȘ݅�<� �w"�=M�o�jM�&��s�3��W�ۺ��:)�����z���y|�	6�Z�L���Gkl�j�n�l�L��C�Cضm�no߳�j�sy�b�؞OoT���S]�}�{Fy�;�������@���˅���{��i'Z	�3�bܭ��Bj�(�Nh#&\Y,��F�G�[�Ę���B���{c2�6y������� Wvgk�,|n,�ٮn�p��P&�;��z��E�m�[)��1��s�r�q�N��>��l|�4���ؒ�ǟSb��y7z�{W,����*��ĺ�*�@�lSa��w�ٶGw��!qgm�gq�o��o� k�]��6GGOoӳlG\�.X->PV(�V����(=��.ᬺ�#f����\�;��>186*� ���Y����{�K�������\ � q븻x7e���ڑ
�ev���:s�Ν��F�w@���ٶo�!�1ٟF)�M���W����Ý-�,�w�D�����ΛFAQH�s� �2,�}Z9;t6m�nU�jW�o>c۷F�.�T�_���o+�.�J_3�q�n,��_G��q븻�0�h�\�x+y�y�Ov%��^������{ޓ>m8=��?
l}M��������O ������G���o��`]����KY��b�� �2!DŇkD�F�
ͪa䮨�!��vA7@���ʓ�����Z�����d>7o��lH�'.G?c͛���M�l�����oזw��)���8��:���1T���}t�Zn���͆���ǻ�?Aޙ1����45\���a�ا�M�3�4��ʦŭI�<���|v,�xfǍv�q.�D�F�
�]�*��\�q�;��H�m��n����z�f�G�·6
9�L���n��bn�h%ţ0"s�xz�w�܁���6>o�Y0����X�9���/�u{P8=��7�j��׽d^8+�Ѝ3+]R�.���kfY�i���m�c�3������]6)�X1L3S�U�\�V���׀׶C*�S+��͊��n�9OS�'@7c���iR���Y��q�p.����sZ�4{Ez
��b�v��7�����s��2R�=]��{��a��c��fٹ$W	����v��]��4�d����2�{��z��o+�g��m����~�OûS6�Z9��pR�p��Y�n5����6�=Di�2Uz|���<WMQ����9Jo��Lpڱ.��d�"�Sh񋯷M,ݻ�3!Ω�٠�lVI�[S4���]*�Bj�p<����d�*v���f���2�^i��q���o\@ɧ�"�Ffֲ#ܕ��דs-�� *�őӼ�g]�`�އ�J��}x���je�J�_Ϝ��Sk�����<�|�Xl
;]�ݦ��̓ngӽ��eC��'M��hyN6u�u�����J�ww>�����5���5س��O^���1p��B:�v�/�f�	�髶�&�;g.�8������|5���|;d��cl�x����/i���<��G��[[�*�
��ٷ'۠Ж��
�%ݵl�U��+Tt��g*[��{,+�(e���*b�[3�;2u�PsW���Uz	�SJ*�����[����9V��� y����j��d�.Ll�n�lu�$��n��loj�CVh����j�l�鑮�]��wT�U�<�>ǂ�/n�s{�e-j�:�v�)ݚ��vTD�ͣy4�*��a�Ĕ�m�(�ГW ��XU'e����x��0'ZH��Ț;%}}�v3e..�I�GE�CZtV�)�"�W�ܛtm��J`\-+��W=��#�����#%靬g7033ɣv�J�������0B�`�<��E���U��/Ư4l&�d��d�~�IE��\��cb��+�n_K\���QUر|j܊M�cj5�rܭ�X�ȹm��6�ѫ���E�6����i1�֎h��LV�wG��zJ���,�ʫ�D�~70X�h�wZ�ۡk��������Id��j5��#F�ca	-ͮlZ*��nm�cV1�ǚ�M�$4lcX�yr�[E��ۥQX�Lk;�ͱX���W�T��Yy��],����B�PI$BB�Յ��qW��QuF�8�+b:��A��f�GST�V�	q]kp
A�8v�-n���P*�ln�jh�cb�*���˄�?����(�<�X���ڎ�ʩ2K0����ۋс�Pvv��j �+tc�kWXp���]2���XF�v���t�7��`��WG.���cRm���6�5�m�lG%����j7�Ϊ�P�MD�M,{&	��!l�5l�/�ͨ*j�$�n��%���vƘ���L3 �1.�g.кP���h!y���@T���1�ض^�7l�s4���+iJ�*�m�Ύ�h���"V����Ca��سn�,]��-�"V��nl�;R� Z��lC# 1rK�kb��,u��,%˵�+��](���mt6�i
��l���郎�A�/R�k���a�9��Bs�"��4�PL�e��M���y%&� Xˍ4ч]��ZXA`���-��i�Z]H^ek�pDƍ��Ƃ!K;ji�&��h1��ҖS����[��_8��b!!��5����+B��d)� .&���Ʊ-��@��6%	`6jMM\�Y�0,	u,c�V�剮�)�#���`�ei�֣�qj�wT�67��.�f2�9����j�Q��yk]"F��M�`�n%�&�J��U8z����8�T�5��%�]]�їMī�R�p`�/]C%Ű
�E��4%�a���:lm�������]V��R갖K.��H��Y��9�%d+wi�� qW�%�,��a5s��,j6���.������q��dR��q]q2�6�It[qHn�%HQw	6=v�z�+-�-�3e0Gu�!���!-5��*S��utt���	�ńm�r�#s��̹u��\�����lx�M���i���^,r��ę5e���d�x�"5�Lc �9q1����T�jL	1����d��n��4�EMf2�m���$8�O1�Z���������4#�0s��"ǀWhj�-F]�q�A��R��Ypm	F�BkPB��#�ĥһ4u/ɭ.�j��p�]�H�]vłP���J��hj�T��P3�võ�t6���?S���l.��)h6d�.,%�]A�
�lu�,Y�&�%�2ʙ�z\���{�qKj��3U٣�`�w,{ U������pl6>l#�����T��{vuC�˞���a�Qٙ��Y����ئ�7Cfy��Q�8󱙫�F��m�}]��Cb�m�p�*�u�=�>J�ϪppSa&w�q/N�vy���cD��� ��M���c������� ��\��zY^l`����wr=wuuy��uLSXI3�d�0��d��l,��u$6fs��Z�HD�붖n��<�>������qQ�Źk�a�;�Ĩ�f{dv�Ȼ��1�?}{�S-��`S��1%������$yj*H���y)s�����oUs�3�ԅ�O�n9m�ѵ�Go��e��oՐ�GU��SS�1�0��|<�dvixۺ�xy���U$>�6�6Z�[[����`e{o�������ws�B�u7b_8�G���=wYku��a�.�� e��g����63;�����`���+uA��>���XW�Wl�3����.�ۃ��/�	8`ʋ�T�.�iKq�)�c���/)�Am*�������<�Sb�e�`磰�`"Y���F{�����M��8�g����Ӈ��+Y�{��1�kMG{6���1��Jj b���6�a^&ݟqy��1-��P��Z��R2�x�D������>�Ӧ��*2���vx�}�;Jw[Yz��-��Rb2����&�j&�8>�����6)����"�j��M���]W����̂'���z�\��I��1���;�]ݹ܀���#��0��y���q֚��\z�=w3�����Z��Є����:%)��Z:\6RkrA-�1I�,(��:��������c�Q<�b�:��f��.��7稘y�Tc���͆�6�*y�g����Xr�S�]0s� ��|#�xd>o5�������m�|��F��x�c��'�i�{���v�l6�UJj8��/E�\�]�4��xO^h}E����پ$>0�A��e4jvkr��7�kh�:gT}Raz(�ś��.�su=ƳJK�<�	B5�!�7*� �}�c��Sa�7�l�6�ew2��qg�~�=[�UlSe��^�c�y��Y��hcZ�k�jln3.3���mئfUYg��|�l}[���k�>û��׹9]�e�ؙ@u��z��E� at.WWe�,V�颭x'��k�uo��^���Z)��0Im�6߶�W��M{ފ��B��:zD�O
�Sa�����0y�د�؟���w|�s��+�^N(���r���������t�{fKʋ�h߯����8��'T�k�O�R�M�n}�غ�|�"���Hhy81҈�.��v����;Ae���ʯX�1�w:p뎍�T�PP����V�8Y瞧����IO���C2�A4�BlA�dMa�f�u��ŭΥ�Uҩ�Q@���m�w�x��Ƶn�-eh[�Տ1�cZB��&l���{i��e�(���+b���wbF�#�Q(T��3!q.�d��l��U1�z�tk���<�Ms��.�6�B�m��eァk4v@v5i6��ܥv3s>�����Vf���Q�@̱.̢��cf��uq�JT���xs	�����������R��r�zzD��ݞ5s0k�l6k�^��\_}]����|������q�.�K%*��Cr�
�a�M����o0י_�A2�m���V�-
�M��]��#ouV��)��))���N��=O½\��o�=���S��Tئۣ��k9|/�nM��>G$P�T��Mm��9��}]Wx�K��4h's�����ft��+V\��-��2埿:!O�b��t���N��a���M6q��C���c�L{Γ���V��F�K�s|�9��3�c5.����T|��,�[cV9$#�ҏr��|��iY�iЌP�ʊ�����ݱ���_���	���C��6M������b�6>oݗJ�y!={mX����,2(G���T����Ŝ;}�׽�l]m���ֲ�a��{�-\�Pػ��y���b�^Usϒ� {Y'��˞��~��}Q�5r
�s⭾���;��{T�ĺ�nt%Rc�f�,�i��T����b�բ�e�l N� ��G2<�b
�IO����FD� S�+��ۜú�����x|dA�G2= �@聻��<��(�3s�����ň�lA���D$#t]������/a�@fG�f!��P�n�㕷b���٭��c�a��azr��_��X����t�����43{�����P��i�����{�
���ӓ������ ��G�b�dW� �G�){)��ى{{�,�:�� �1-�w�syb̫�8@���^�vDD�;�x��9�����AF�@}�k�^rd%[W��u�{��W���B3���^ ��̏f@o���}�'���IsX�#+�t]:��Mn�-���mRnP`��AS32�����A�DfG�a���S>˞ބz��z�&���ǲ��/Nd{2�>9�"�^������ݨ�@�/PB�J��ѹ��3*��x�!���^��<�9��n�� A�A��26r:�$����Ցz7*��6 W�/�@�3�2v�������3Jf���]f��(F&;��Џ�7��]]��Ӛ5}]X-_^��]g	2��Kw`����/���`*��ݾ�<���=v-�ܪ.�¢�ܱ���*����X��B���{2�'2 ���d��)�	�b��	���x����\��"h Fdyf!T����*��`|�M>�	��p�C�V�әc��DJiL2�R��Tf{*=�z<��fE@9��h9���1z;*|�]mRpf�D��qD��̄��#�k��
����Ay)��Ů�\�#A9м9� s"n���j^瑱���&� C1d Fd�Uk6�T�,���2�r��<�h"3^9� s#������:����D�����d!29��LV���" �Q{d�2��^@��� �@���fA9�3^qp�/PB��qK���Ʉbc���Fb�@�A��U�2#�
���]d�#��lC�R�n�tX�eL�Z�PVo���-�5�*�f��ΐ�)Lػ8�t�#=����ÿ<���2�b�Qm��h�f�,��1��X��^V�h	��MKa&��	.0�j�,
9�[1��K[c�Q��@)��XGp�%�q�e�ˍ�d�X06&��f
dkGm*�-��mT����0�sa�WR��Mh]���t�Θ,Uet��Ļ-,j�Yxi�E�n��lݙ�nYvZ���~����C_�T�і�M���B:������@�\U0T�333#c��lAZ�dz�����t�gկ�79~K���$��E9�9s��^#1��d#�����[
}9>������)�B.� ޠ�s"������ڀ����D���4�?i+;��w�z^0q�ty{1<s!x�2#1;f�m�ʈ":r�G����s������f��w�>=������Sy�]������Q���A�ѹ�Ywg�g*���;Xtk�]T-rp�2<���W���q�o0�T�0&d(A)�;%�(��nvcml�������e�?�~�&�|���P@����Ay)��1����p�1�>ٌł��Ȏ��޶�/ax�s!���2"w�lo:�Ĳ���$��
���c�σںŀ�u��k��b�_��pr�N���K��@�z�P=�p�v&F52`����s��A�܂�u]X'��f��p^����#3�^��=�^ &�2��ly�9���!ݚ�� ���w+��}K��g���*���d A�b2��x2y��x�p!���b)��Y:�)�
Q �G�tNE�b������w��H�Fb����I�̇��=ӫ{��|A�kAx���#˴j�9FE�&XD�k*2�v����n�b%�R��2���ڏ^��s!Ā#�a�c���5��Z�=����*B�øA�AxۄA�"3��#ݲ�n�N��/�PP�޷�u"
���S���V[򊫇'\".�#�Fb�dP �1�����c܌�I?8pv����NbgnWFbڰ�<1L9�npɜ;z�4+�� 6�+�%W^M]�qj��pD�[hc2�.ṟs���g�����Τ@��.���w(h�#��p��F�`�긅�;a��ۨ]p�;�[v�;�Y�Nv���YN�d2nl��nb�Ň��Fg�Yǫ��c��4�X�"f��k�,gX�|2�G���j�ZU�^�Z���n
#(p�G,ƌ�Y�G�h�}�gI��u��<�t�5W�b�|�ѝۻ�;{�umr��i�MQD��^�\�1�r%L��s�r&�{�on��y[u�Y�Tn��y�p��%�����Cf%��MXؼ�U��_z����K`�Z2�$o&dX�ƽ,;�� ���.������3����x�i�nqG+S7���E+�X�!Yx�/���_&z��� 3�RM^Ǚ��P�|_��Ml���
�4F��6�����SI�����f2Ve�M�6AW�mw[��z_d+��]�6�0/NR.��q�en��@q'���ܫy��-�N��R�V�J��:��B �`��nJ�"�-����0;*	İ�n.;�n:�jś�QP���p�d�&Y�U�1���vS��y�C%W���>S�`�*���$�7�p%nl���W�����Z��r��zK<�b�D�����U�HD�W����'�� r���k��E�75��
 �sTU�X��FM�DE�b��lh����b�2V'��������߻�*62b�X�ck�ms��Usj(�m���m��4h��}-�*��~��Qb���W�Z"��F�DRG��`��m�*��m�>��(ך�k�ڍ��b6M���"�E�آ�6���Z)6�nX��(�jf�j6���[���ѱQ����V�D[�5JSI�5$$	�z�w��a�F{��{U^K���@�5���K�1dz�I�����4�H݀��^ ��/v�;,�᭕B�8�
ȉ1Y���g* ��"3^̄A�"3�%Tt{T	��j��)�Q�	}^�A�@Nd]�z͡; �2H؉��GCG�H�]ή�b�x���j��Y��W/������Fl�Y�!9�W�u3[��ג�;"&h��`���"�/�̄A9��cH�w�"�� z���Af�r燻*6b��q�D���gp��Ǩ$�ܯ A܏,��/�1�b��\���ӗF��Ȉ��|{���s!9���/ e�Zv����/c�و/	������{ћ3^��@�}�F�X����L���<�3����l��-˱Yph�����+5b�*��]���n�[��t�*@����_Rhߗ�|�9���^#2=�R���]r>�^؈_f��^a�1B�z�6
7 ��kӇ?%p�^ڱ��f`N,L�jа�&�1֘6���&�]�vve��2�>����3��b
��OSު���""c��D̙�V��$�A��7��Fb@��ѭ2�i�Q70X8�}�9�w����ͅ^K��B�DfoB��Qj3��y� ���3@�]_� ���
�nx�:^�/{
��p6�z�9��A� Fd����ઌ���z�bޔ*���t�dD(���/��8f��!j<�[��3����2�gg]8c�
�ٻb�g��N¯%�oah"3_\���l�������~Wk+���@ ڛ��L��d��\��S'[왦OX�e_�)�ʱ���6��t�Wf$07]d���o(_X�60��մ�Y4�MChFTM��qp��y�7���Y����[Vf$�n���:9�"�-��ئ�uT���у������^*銃�k1Y�.ˬ`�G!��r�J���6�/na�jW��Sq9�[KK*����m����[лM�����(�n)���r#��&��°�Er������a���a�+Ŏ����.�H�X�ʝFb���*�*+�����?.�'ϛ�o�&�#l��-eP�zی������ Busax���̥��D(��H�5M�v��В;�^=�(���i�UeK�1��� �AȰ�f臭إ�"|uG�P@��"3 /���fh����k��Y};
��ۄ͠3)x�/fEx������南�:�Gv ��5�����=:7eP���{���}��J�ut��H�]��W!��ՎE��HϳEZ,�7���� $ �8o�G2�A޻���k��
	4�|W�5�-#K��kVǃc9	i��ڗRfeUAƁ5�6��̏f@�Nj�]�v{�aW�� :�u�Ax� �d A2�u+�����nkI���R�V��V:�<����}�,����y����$�̅J�Ng6�v�bvI��Ш\�[�z�����p�}������vU�z��^��̉����e�`��^U ���Fd�Ax�1	y�](]���t���Ddw�>;Ё���2#1 �T�w�f�5��՘��[���i��.ҫ�p^y�7[ӷ%B�*���F�^>�A�D����9��ՙu;j8��+��<���b�z7R��{oW�#�ᘼ���;��X���j�b��bR^L��b����ci���QS0��؁�ysA�Y�(��O���5}�"##�=s��p�A�Ds! Fb�j���LD@fr S���nj�wi��]��p�!����{ފ�u����h�x��|d?HX'29�W
)'k��96M:qT�T�;�V;�+Z{rK�����L��׎���2v\Z��<6��L��`��	���Mc�zU>�}����~��?��7�q�́Df@v��:Gtw�;� G4��EMB���{3VDFGOt }�ƺ`��c��&�<��F`���*�Hh��4�����'�S�UI��0��&�"�Ax����3�)�5�1Q�`G�"|��D�2AQ	D�f�DL�	t6�h��`�cn�;;[��w����~�:�}����=)��_iV-pCSO^t>�%�j�wW�ǳ g��Kّ��櫡[X�m �����wN�����Ȉ��=Ј _/fE���U��^":��h�u �W 7W!�j�E�Bu>Ě�U'��%�\>6��6�f%�3G2#�`���yvN/k� ��T��	�hƌ}�lZ���=ջؤ/Pȼ~���ٺ6�#W�"��'�d�9��]נ)ܐ�����r�^Q�8�3��_\����"��{2و+���}clT����j�9��x ��^̊��d=��ۺ-` �8L��	svsL�P41Ie5D,�K)�]5��Er���{T̀�d"�C�����HN��OĊ�m�[&u|�����Sb:���l�(�,�A-�S��O0�Y}�`���E��dg���8�� ��ix���L�qF����<�p�Z��FG;�Ig �p�>-�$6�֮��r�k��{9Q�E��7Am6�o+;*�ǳ+�.5���➋��J�@���܂�@�mI6�-ǣ(Ňc�S뾻��'S��V\��΀��hH-���B*��t�q�I����*��9�::ɢ�\╇3�]�Kf:t�O8R�r���5�[��tyF��?/���{�?��~�?"�nD��-&��+���;F�
@le��B�t�պ$]pu33�Yo-.ؚ`�(:��[����U�e�iv�[va�E��q�H�3�R�b�-��bAfev��k4ubslB�W ��5u��7Ul���X�P�sS[���.(�̱���-��6����&�����[��Թ�[�߿%��J\�F	+�tl�M�g��FP86�"��L��fe�C����Cn}>lU��}����;t`��t�D���eU�mp� �ڟ�y�YZ�n���ԍ���!���yU��8��ۥ�ka4��*3,EӨ���\�܏#o��Ch [���ڹ+g��D�fS��iX)w� ���>-� ��!�"D��7�oK����m7
�{����n&2 {���}��s�t. ��Rm-�	�"Kq���Κޮ�"X�-�&��c'�_=����>�� c@6�|[@��y3s�|�FY������`0�4�!c�̵i��q̣Rh�r�̙���2�I�nڛ���+;#na��b�!�N���9p$��Ȓ� ��!�����Ekz�U��yJ�"��_�����BMΘ;����u�.�fE��0�@���TpT̙\F˅R$��ɨ�1d��9#*����YC�>�^�X���o�̥���FG��Fj��uT��W�]�w@��"mȐ[�>mŝ+���z{���b:���zA5���n�Ŵnv37�8�_JZˏv�KmM�va��㶡��b�	ހ��^B��u6y�A�"s ��/Ch"q�n�Z��_�U��U%��_%��d\{�;�{6��	m�s�E�����lGH�F�bT@�����o#���l{E��1/M�32����w��O}���p�!�کܩ��Tu�����.�6���i�z@��E���m����S�ir��-��]��a��㶚�1b�/w@@�ּ�N@�nՙ4"mF�Ϥ�����	�u�LM�ɇ�犲�n{�V4(�bFg;h�0,�yW5P�9]�!�i����2s��T�w�G�/�u�vuLf<q�q���R#5y���6��t�K��� VZly �uT�T�q*+�u%�zA�F`X��U�����'�6��Q�Ԑ�[�-���O`i��f�sW��}."�.@��o\���ChI��;����UD��L�4�����K(9�2ؒ;A9��k�a���ɽ~���"9�D6�|[AH�+��Y�sp��t�[\8L����U��A _@�d6�%��B��c�0Y��/�AN���$���Iy%�A5���h"yw���f�y߰.A��;���[�/ڶk.���wW&Sc��gX��{�/\�����6�zDډ=[���/�����T�ҫ����1�.8A�k��V��^E^m�$�G2�"�9k����H6Aqu���չ"/��A�y��W6�
�;�Z�����wJۏ��q�A_��ߐ%��6В�GV�����T�*��J���K�.	��8�@�^��8�*��������&�
Ts�u�K��ɵ�ee(�jcR)
@���
eL�q�NW) �/7 ڛ��c:��mE�\���;r��;p>��lY�m-���*�K�f�F�7�D��W�Ӌ��nT{��^�3P@�*ќ�Cu�Aiq�D܉�nׯv���9U6U��	y$�[^Ƃck���[��T��jc![5i��;  l/6ԋ���C���FŨ��<��~�K��,�΀v$�y��ε�&�j���AJ3�/\��a��T{�sS�3` [�A-���ѳ ������b0q�%L��a�V��f�@sf��,Wb��g���j��>5��ˮu���]�hJ�f���a���B��i`X=|�t��|���Β^�;��ڲ]w$� �ݫp��B��-`3����}��t�)
���3wD�0��4��z�p&7wV���l�%�.-��؀<r�h��]yw��cUs��WG�����>��F�r������թ�u�.�Zf��ěŏ��T��ѵk-�O�����Nf��@V�DY�$�ʵ4E	Cf�Uh�H0��9�%^��8�a�c3����p��{��|�X	U���r��l܃���Pk���{������T�W�}}kۗX�y�W�%��ʗL����H3���!��ܐ�!���%gWJ9Qa/y�d�:��ū��J�o�U���VV�De�O��A�+�b�ҝ���y8�P�u�m2�+�hѵ��m]ޟ`�AM�[�^̙xh��6� W��a�8�C"�bcU���%F�
�*��̤Y6�&"�$;5��nf��#T-���3$��[���u�g`�h>��͕�V�":��W����}��;#<1Wu\��Oaw[�>�Q�|��,F��a[���V��a�E"t9�4loF)���c� I:[����z7k٫�/�*�9D_�ocޔT���6Ʈ9�0&�4��套\�� ]C�D�yZ���9�@�h*2�"!Q��1���-�E��]771�wQ�ݹ�kܺks��n�b�c���z��n�+���xZ"�c���=�[���j�unE���y�i+E��ƪ�Qbض6��[��jJw\�U�h���b�b�W5I�\����U�ﭾ����W+r�F��ƍcW-��E�ت1��{��V�;\�2_J�)H־��QU���sk�lm����כ�ADj-�j����I�W+&�O��{����������wS����}��.��@s��D��e��̓J�^8y���&�6G;Q�֋�[��-�u;�"ݻ6��n!.�T)T�a�4�ZK�YeV:[\�5hW�EF��n`Tr6��Q0[1��$���SF� �';<w+]D�k-�f�#���m3,���e´�	.)Z�+@�-�Ft1k�Ŷ���lJB]b5 �0��M*.)u��ͬ�KjS,�2Y�Z�KjA)pli.�6��Ycr��ܚabpn%��� �	VW82���!���6+��L��#IE�X��#�����w��k
ۥ����q�LW^��B0��h�-#�WX�9��L��ѹz֤C�E���Q5t�Y��M��V	Y��G)���ย��R0����6���2X-�K�I�Ů.�Y@�1e��3�bhm�	�&��x���q�e�r�T��z�`�A�B�A�#�S9�4��R��-(h���5D��.^��a(l�)�Y�-�Ύ�҈��Aa K��si�l���t��v�V�MMw��"�쌵���3G��Q�b�k��h���Qr�h���m�[�A���\L����)jm5� aʅi �s���iZ�M6�l��Y��B0��S.]q��f�;C�1�kjA�
,Ͱ�4ˊ]a�l����LM�,��49�b!��m�.�L!�.�P�F؋a+��is`��at��ЩTم�`�Kp�s���.v�"Z�LF���՚6�#K�6�ىM�P��4�MkLN��Ȓ�;,]n�W�f\�XF�*@®�Y�ޫ��ƄP�V*%�������\�3W%��l�A�	��4.�3�,1aVR��²�3l��i��UUUUUVӎY�Kqj�(�"�#�VR��u��6�˿r���˸�����������MeK�CY��������[C`�b�A���Z���G.�@�Pq*:V��f�O�����(�J��L�V�R)Nc���Ƭ-m�[��+�T�[�o����B5��s��8�$����xL39�R�!��v���.HL��� Ħ�`E�4��bD��]�����w�_ߤ'߶ZD����	d����5	�ceR���ªǜ]����~�/_����n ��O'�����{v�%�C@ZdFł�A������ 6Ղ"�NO]�<����z�n����i��綩�/w@@�ք��)P���� ۱>>m	檣!v̙U9����̇'y�H�A�6������S26������[� �:�u��{v�Iz\y�R�q.����s>9���|^5�my���T��X�NZ�v�������i������� -�����f ��1
`)(�j)���ʶy]"�4��1��B8��\��]?/�>}��_ �mϧŴI�����}��&8��9+�NwU-^��k�>m����p�u)�g��G.�e�|D�h���#-��]F~�.�2�ue�<%�x^Ʈ�6�б �qX+��E�{%߳d�MJ�Z��?zZ��7��}'師��!m��+�.�Ml"4���9�׫ۈ#��׭O�!������X�o&��sub2��F�.@���\��������-����t�ǖ4�����hRQr�s�ʝ̇�5 �fmA�س6p37 ^��l An ��H-���"�����-o$�]�!ugi��H&�=�k����6���Ѫ�k�HAY�����@���s,)Du��]��jK#���3A�E|���~�d�v��p�%��^����w;��6)r�U*�w@�'�	:��CnD�[����9SqS�������&f����̙��q1�s9I5[����p��V,!�@���܉ Cpd�~���y��MX/l����*gM����*t�{���:MO;�3iׁ�c�L5�ar�t˭���3Zݹ���o�FN
ͻ�zb����K�H'n��D6�|[A�(�j���(tR��{z<�m_c隫s;t�6"���1�2��5��:�@�܉�p� ��DcgV�ף�� �H��z�����C��>��$h"�"-��>�<~���~V�����m $�Nt�9�!u	���d5�jE2�����ϖb~|cǾ� �=�v���_i���F��v�����-�7%���Ɠ���(�B�ܦ�_L�Q��ݦQ�J=�zА[�AdF�����[@>��q���܉����%hvvm��-��v���� ��ԑ��|[jHmyz��dnY��6�y���A=��e�ȣY�r|�C���EU��<���\� ��

ͣUZ�nA���X'�^�yc{�C�s���^]��݋R�T�.�Vn�ؼJ�Qk%W�V����z{�nڒm[���\M��JB:�N���/*nw�hR����@��BKp�-���U���:<��fO�)�Yu�ځ�mj�rH]L$��F��F�9n}����/o��v���U2"E�v��S{��G7_o�1)�kG���p,� `㻵Y���X�q�7����f�^5��'�.�AۄA�{ �qE@zߣ Y�� m�$7��mL��a��ިۃS\��cc��lEw�>;�^�-Ǔh Cm��u�lDU�(���Df�ψmS&Q��ޗ7�\\{�sR��FS��Ex�G���$7x�CnD���2I������sW��ӓ�	�� �������>��O#3&��qG�ɶz��tn��� �o��.V���������vɽVp��)�"�fGX��n����^�OI�%Բ���z�aih�5�=��!uP����jƔ�m�@bgbs��%jm�2´�LJĬnt�hMA�h�ee��4ZYe�����r���Kun�l��0����(ᒶv�lBg+*���h6l���Y�����R�[l���-�%�Ibi����(j����Ֆ�&�Lb�ie�س��~}!LQ 
�f������b�i��u,d�����(e����:+��F�-��S��9NUF�o�lE@JC���J�` .�D��D6�m�e�@��n�v3��۪�)�k�7P��(���̫���㏯��A�@�p�qؕ ���v ��In��O��uy�yȬO�\�;�g�.�N�y����k���'e�-�� ��8�x�[jFes=9U�f�v����p8��aQڂBW�$�B �9 ۱ ��|��Qk�)�*�E�T�);���L��qq�5�H �A�KmGfڠ�1�L#�lJ(S4�E�k�X�k�[�����`�j��l��>|��_���������Ow'[oY��y%�2��ѓ�nN	�d�E��-�7|�S�\n��VO2�cFR:�虫�O�d=�(�pUP��6���ݢ\��X�K�ǳh�.u�aP\�2����6!=�����>9p�>=�)̮霝��<���w`"/uy�ێ=v�@���M����|[Cmg)�Yx�s�UN81����g3!�Ǹ����^-�>m�!�S����Zs� 魟gE�|�
��5���a�=�~����S\IV�6��
s=>;���x���Rn�n�sQQn�� �ҙ���VVƻ�w�_/n�Dnj��y6�d7�����^ }@����V�a��0�H-tQ�S0q����n�C*���0�����혞���i���nz�r}:�μ�f<A�A {��mH!��	n"mO���vd3Y���:yf��9�w�K��p�-�tqLc���������m�!�� A�m��Jh��a������Y���Ɩ�,ݵg%��=}~�[�'�ŝg�xj\6��eL�����K���Z,�ƚ��t���]��s�6"�|w`"��p��n�m�j���;';T`"�ǳ�>!�!E�^oK��C��^/KY5�]e��L�z��/a	�כ�/7 A��In%�PGtGUY��)���{�����K���1�k��E�ۚ�5Դ&L�!A��"��Ai�q�R8r�,�`�Kq�{B��
�����A��s=���ox[jB�n:��v\_;�b/�C���Ju=1�_H��"��Cnd[�B��O�{�:jđy���"��Uo�RY@�U�ծ��A�m;�sQJ�9S�;R�\Amȟ��2w2,�k�o�l��v������pmz�h"�{���[���V A�A ^���ԅ}��e��j�n��� �ʞ�0y�씼$?e�f'}{E����ʸ��n�0���P�E����~	2�r��_ei���3O}�hZ4n9\\?��|~��}�m̂p�n!��R"~�{Sh�~���B���7�����qq�A�j|Aւ-�m9U��,n.F�"!,%��DA���Mv��1�M��%�"�Xt�"&�2����,������o�h/T�D_<}1�.����"T9��Ӱ,����-� ��RsQ�+�g��A/�w�}=��ɸ�{��A��{v[�$�+b���ͳ�G
��D��|@6�|�LI�[;�8&�;w�<��#� �5�p,��mH!��3QVP�)-���u� ��!S�}m���/�.�|z��c��%
�"wg��n>m�����V`�r����LY�Mk=�ͱ�@���[����-���UPni�"�cΫ<��f�)�|�Vu�u��l��n19��lRJ�1�T>�P�4%ge֕A-�']9����".I�m��M��Z
�l��)+)y��P��w��Mn���Crp�7eĢ�u���h��6K�l��h���C0���+�Ќ-�D��1�э�f2�E�u5��6�B\Q��Y��tj�6
���lvDtt�Kr���#WJ���0$*[�����$k���ԩ�P��-���U\��w2��}����q4��\���[��B��/j��i�k�A!��W�oݹ��	��n�ŴHQ���݇r�d8��Ֆ���s-p �A��[j@!��	n�d�pc��ҫP|j�G���O���V_�] ��^ �Aۻ����U��'^.� }�T��p� ���}��y9v%��lY��m�b�}¨��$��Aې$+��8"!�H ��#�O���HQՓ�[��-8��A/��D�LP���]�t����א �  ۑ ���R�E�\K�N
e "Lp��z�Mz�����4h��ϋhgF��T	j��"* ���
�ɥ&��r�0fd�il�C7i��fr���!�|��-� ����:�wyU�Z6"��pvdq����gO���n!�2�`��A;J�Uu�5��SKze�J�)fJצi+2sq���c/f#ٮ���+v��Tt���$�iU����@��|C�
C����ntkyI��A�j|AZŸ���j09#����k��,� /6�In �Ї3sr6��5f�}Yn���$8�A�4����p���!,��g�,�p/��ڐ�s�S{���kG_/=�����d��:�GYʈz4��#v!�"A-Ǜ�=���V�{��끠9
�cv�:3qԸ��A����ւ�D�Ù�g�߿^GxF�_��,)�;�����l�GQ��1T��32�Ї���W�����z-+��w�ۚ�򄅙t6z�����o �����-��d8��������r��εMS�c�Z,E���� ���-�.��m���E�L�^�!���m�>�W��fp|zJ��*��b^2_���
�Í�x���w��KfM�w�*P�p�L�Ԡ��R1���
��X���ہ6�o��kv����Ow��F���ҹ�n��n�3��Ħrބ�p/G�HR��:C1��,f�߹cP[zN|�=�_:�(;a�vW+a�w3o���h�g�^�"gFM��U1E�m!vma�B��'��`��=]N���.��D�'vP��o�+)A��-b��Ӛ�3`cKg@+��O������%<��ou	��
��a���"�0�=�h�!���˞V�d��s{�,�Șr�e�g+
�����c���q`V���3m�.Vp����}���>LNY��Ό�6�;éMr3���[n���w�b�$d���['�Y��>w�`��|�ܲ�N�3K����M�}.^�c��M�`�Dȷ�n�a;�H��.�+(���uso!I�����KC�14k������IT�9'ٵ���ʘ�p��(h���(�dѽ�n�e�':��^0�K��PQ���������{�槖:� ���8cz����F���H��DO��]�݆q�Vl�4�m��һ^����j�>��&p�F:�i��i�zaZ��uE�����㱛6��y�E��Kc�[� ����"�+�X�ö�:�
�]�*��T	��d�U�l����5ceNfi��wx��igK��t��e������۔��@ώ�� D�'ĔE�k������@��I$Ow1Dc{��M,�r����y~���Rm���7$�#	D�$Ԉ�;���Ηg�t�p��;�@�&�]�MΣI&�"�\2F�tRw\���Db"R"�E&� ��\&�]R[�p����dd�MΚ&庐�	��e �s���.��LO;"&��sp�� T��cE�1�5\�Y6	��Ѽ��ۑ2�sE��ͤ6�\�^W�{��ۼ�K�snN���Ӻ�+���s��3�V����^_�k��^\�_�y�N�ͱ�Z��`�m�\��[~�\��*5r�TV�ymsX��b������IX����cF���(�گ�U戟;\�E��r-��(Ԗ�b��ꯦ�d��A��6�*�_O6�5�E�Qnm�|my�9�o��/>��?����7�ї��"���_)k�7��RCh �h��6θ�9Y"A{@m3�j��ާnj��.�Nt D͍���1����z|s�@���Rn�����eT��zZ�׮�b���kh�k�����"@-�!����Oo�S{����t]l\SB:4�H�k���!6��S�!.�Ut��i�Ǟ��'�4���W���J�\ؽΌ�u9��9o�t�X�A��mO�m�p2�]Oaet�l�B|{����苹�Q�Ֆ��a!�:c@6��֩*�:Xi�/M�RCpn���V�L���p�o�Tmf��cyy����O�p�-����W�:�=%�N�Y�v ���|[@э�gs9Gܲ*�q�]��')w����%�;cY��;��!y����ì��p�����z���x�h�;ڼ���k3,���I�f���N�F@��T;w�`j���Ё��5$7��mȒ��������GE:y S$���q���ﲮ�z=�ۙ��uS`F�������#��k3m�V��CBj����,z�aVX����I�^{� [���ڕ{�h�S��11w����ŕ�{ ^[�7Cp�$�����j�X�E�^n���ז�j�u����A٨"��\cA0��R�H��r$��
�7�9�,Ԁ�y�y�yE�����ʺ��@�1����7�%M��	t��4� 6���u�9O����1r��^Z�Q��Ϊ�wE�A���r-�!����Y� A��q>�m��>�ܧ�Ws׺���x�j�栋p���C�\|7�z�	�f`�w�(�d�qpq�9"�oJ]|Tة���Ntf�V�(�9w)d�x���g�bL��,/[�U"[�u%EMcC#�]q)5�Ju��!.�R�c	�@!h���4�֪M�&��f��UC4U���r����hC��.�M�Q�ىBсH���<�!f��YE�lh �:��;m-ub<��X�3\bf��gv%t@�W8XRh�bs�b�`cC+�-Fm���R�;���$�MW'kv+S79�VR��Ħ�ԋc�er���n~Y�}���� �6��������wu~�]!��tfl�OE]��'��E�^ ���������4Џ����3y��m51@��#5�7	��|n�����|qǐm �^�К�כ�:>�sV��v&��'�����n�Ԑ�	�E黑��#6�I�[AN����=].�o���Ј����a��Cw>�����[jH-�79�C*'��R.����;K���1p@�����	-��:*ڵ:�uK�Y
"nH)�d$"U�4ֶ�T�s��1�luؑb\�r��.%ϝ�h Cn}>n��u�^�E���NFG67%�͜w�6U�KΚ��A �Ԑ�y���C�'��ݑK����5V�ANfHk�E��6���]�
�َ�|�4S�9��Qu��`6���_���k�SF�sn\��+6G�������A���bz��S~0�}�q��m���"&��P@�B>�jHn-� ���Cr�t�p�6��z��\��9�D��|��bEg�W)b�f=cZ��O�h(�y����{q����H.�������F� �椆��p͹p"���kW�+�?e��l1;�)���	Ώ/cA CnD���ʜؼকG�Д$	S ��(KA+SP�.��`�1�k6����ʹ�2�O��9���ߗ�����jno�-�w��5&1w����Y����g\y6�6�	��/���n��vlY�ώ�G��^�u7�bnp ���Ӛ���ڝ��N�.d ^Z�G4�;�mȒ�"hU�rb��&)�f�ݚtB`�����RO�iha�u��9��q�[f]_��+z9��~\P��TƷ�o�k���ҽY�U�M�B�O��q�����h [�Q��!t���ɂrЀ ��V�gfzr�9��I�\��}N���y4��H<�{P^!� H%�^ ��D6��3�&�(�Q�����]��*�o���8�9ڽ>�A�Am����/�/������W ju� �-�h%�ZԉX�d���6.u{j�gl��D7	� ���7�ʓ1|A5���3&����x��O���q�[jH��eM]�ݡ�6 ��J�u]u[ǝ8�cy�y�InH:(C*�Ν"o�^#]� �� 6�!�>�A�v�^�wN�;�ù�{P�A9ڽ��n<�mO�n=��,i��_@�eȐs��	و����H̙�(] ���aێ�|F���������B�}cDy�\�\c�F0 x�lB�jWne���eJ��]��8�b�A�.�?�P��ק�^n(����y�)�Y<2� �㸛[?_Mm��>�i1���@Dz�H-Ǔh`��J*�;��f#�/J3!L�d)�]�B��6i
#��-%�R�WO~�y�>�CߺO}���6�[�lCW|�*�����U�322�_�q�ؠ|�^n�� D�t�n_�k}w���j#Vpm��5�O�� A�@��c�������
p(����7�p�A���"��x�;�w�e����t�/Zp�-��m̊U����H�3���A GoH�7
Zf��Z���U8�) �B�Ӕv��6ƙ�D��A���!�>n3j=�u�R��Ֆ�h�댙�BK��!�����k��1��b4��뻻&8�]T*�=Jv/�_R��-e=���ᘭ�{3��r��B)�T�{6$�Ä�{��\ي'�^��G�<��-63��u���Y����J�0ʖUfQ���f��.-��Eb���Ya�q�A��ƶ8*�u9��e�c�g]`�n�9ޚ�m�5m$!H��i���+���A����%Jff\ʋ��J��Yo2���YZ�P�)��	�n����dJ�� �i�F��4���V��jӬq
�|�߿l�LCpFY�-�fif�6CY[6b�]��=e�V�S3�Q�W/Oj��mM�u��WSz�7c!$�%\�k���������D<k�ő,���e�]	#��|{�BWld>fU�i��'�/NjŸ��⮯��zT�ܐ><�/� ���n%�F��7Nb0��L׌.�Ä́!�n���@���u��1�k��Ax��>m����]j���K.��t�&�y�YP�M�@�B ���6�H%��p(��ɉ�����Ajfs�Gk�W���6=ǻT�sW��W�mUެ��z�����`��)�� �6����X���
�7kRT���2�X{�M�f���In �Н��k�	�� �Bм� O��A�ڲ'ՠ�s&�VDD����t��;�X�)b�}�-FI�p=�}�L�
|Fs|�ڏ-CB�N�y�[���..0�A��?�>9�"	��R..�>�o_F�X1r��ք���GY}=��	�~�wG�h݉�m;���YgFf�7��M(����RFlp��j|Ch!3U�+l-�uO^����$Ј!����q��8��a!�9���j#�A�nl�ٞB%!�$�W��nڒm[�Y�&�v���Ήx�쥃	΀�5ȟ�x��*yq���+��f B�$)+���؂AK�#6+fq	�мd/X�Ζ�e*�'�~0<�t!>��6����*��k1v���eF���=e%zk��9�#�>̅�3�@^"���������@�A
�1��C���Ux����D7x��ڜ�,���<�=��W��e����&����=��N�SMKB7���ծX'A{/�]��z4vv�
����Bmv��.9�)v�'��G��8P�\��8��/� NtA�r$�m ۱#38�Ɏ�A]W�Ƒ59����9�,��+/�ʍ��R��7&�ĺ��m�7�p ��"Kq9C#�u>3bƤs�/gq1�=u����^ ��6�O��f�k��y�}��D$cD�T��H�������a)�";T�ūk���}�e��ּ�z�mM�^�[s9��jI��f��*a�
�Ȑ_B ��6В�/4#�-��!:�Ϗr��ۮ���eF�Oo) �^n:��'2s\�ʭ^�� A{n|�X ��+3G
��^s��rqex�C�������7{Ÿ��p�9HM���Gvڑqw���g6�-I1����~��cu�&y՝#�EK��J�NXeC6�_Ƕ^����1ӽ�\P|�����sy���u{�Osw��ϯ����7�D6��	n�!�l�����{��W8�oqڬ��*68����5�^-Ǘ�m�����~���%6�9Xm��\@[�X@n`�����b��H�D��/:��wdH-� ����=S��}�W�.0��<���==�;zg�6��n�mzGgNGY��G�9ܦ�;vo*w3��LEw�'z �qHv��v�@k��fǓh"kӍ
��KF�ݾ�S����_i��	��> ���D�S�A�	����f}wr$��7:OVVr���R��R�H �����*7�������[�A�m�Kh"���u��{�O�7q��[��e&)@�s:D�p�Cp���d�3y\��&�f��I�y6�K8-ܐm:X�0!W�8�u�V���>ˮ��4Nb�A��ǽ9���(���ʍ׸Q�!|�р�r��0���!�ܸ
�GÖl�	�U��fR�U����r)e���_��m4�]��p}z�^�)�)%	���\Q�z�虚�õ�H�N�f�Ď�;ǉ�����jƲ��k�����z�.9����t�g#�K�|�EL<ĝJ�t�W,��fd�͉�w(��J�;ocw7�$�ے7d.�c�Zɡ�%���Ue����������a�RX�w.�2>ˊ�CS�S3h��w�ͺ�rw>ɔ�^p�^�gbVͥ����f��S�s���X�^m�	�v�����k&]_Q�.uL�q�B��.�gM���wRHp��]��.�d�b�j�Պ�iz��n�F��d?k�6�C��Yb�еJ�WC�XT/�[�"��1E���Hy�]�l�I��ݝj]����
�
�6&�
T�̒�"���ߺ�����^��m�YV2�[Ed�C7��c���ݳ�8~�NkCtq��`�q�;�(e���l^��ױ��2՜�0� ��z;"�,�B��ǃq���Ljh{V��,`kjn�3��mk�g$uN�&f���L�v���[We��:̱c;Kїo?�����qTh3����[��5�6�Q�IlEhشX�&��*9m}+sEcc�lW��j��\����X�j7���*���Q�1jM��P��j�j�v������j �}+������y�ب�&����-�U���_=�~u���\�ţV-��Tgv�mҴ[r�mDQ���}[��Q���+�J7~z����[�܋c�Q�-������U�p�&��^�:	�'n������-�͹ ����vG$��S��b��iF�R�B��Cg@얖�1��C�],]�a0ڰ)�aJ%^8�L�\���5��isMi4]�Wy|�/�T�(f9A���Zj8�D���4�]���X�K�F�ŴU�.�CL�4�ˍr�٣���61�,�K�9o���fj馁"�3k+B�;i��"X,����H S��Ex:˦<[q��R-eڬ�͍U��c1�h�c�\�U�eu6�J̡��1��b���LP6n�!��9K*��a��Ji+*�����c6�X8H�T��`�e��5Gm�`���XcYr&�h/j��5��Cg<���#KLQW%f��F[������aZ�,1b�ڴ�M5�CplE7Q[�ZۦYQK^��X� � 4F�ۑ�]t5ص�T 5�Ne��V,�깘�D�!k��)��:l\DW\�n���Z��+���2jF7B�K,
���h���v��N�q�Lܶ������a�*"�,�ZˢlS)%����pumډ�Qְ��e�b1���.�]l��4�rJ���6�	�)4(vb s�v��*�k��P�ڕԙ�e&���uXWn���]�%�mc�Fl�]*A�ɦ�����̳`1A�2�h�v]�e�e��n�n��1M��H]��5�ʌ�w,+.T�CC������	�B�R�lͷB��7l���(8UsZ-&Þ�%B^��c���R�Gf�R������$nD%K�9�Ե.�e౰���8Ի&�(�kJm+e��1����b��7�nG
���I]le�A�͝�3M�����1GkL��+��T\��ܮʪ��h�M.%�֕e�v��#Y�L㲖�j~��������ĖQ�jm���!Z���Bh�ke�se�k�M�W�`�4F�l�4��0��MK�FЮ�E���T��iplX푖ЌC�rij'mJ&����,�p��m��V7&��gbi�N��,I��%��Wq��k��5�n�κ��
�vn�ۡ؋LR�c2kF"�ƃ�6/��_K�A��&ba�˭�̐JMv%�K5��+����&p�m�~z{߇��πD6�|[A	��/���;�2�c��De͎]��iYu��� [k��@�� D��t��^�>�B+I�ܚ��������ly�mܽ�����ek�OcRAm��yx�Ԣ�x�xF��(WI��OPB�}�F��BAn�n�dYKm�3��A�#�����f]��.�v�Q��{T���x�\B;�T/s� ���/@mȟ�Q�}9FpӚ�ԅ���W�J��c+�H ��!��s�B�af�gG,j'�J@G���Bd��驌X�swX�r���X�YV�U��濧?rC����{��͵"�&�^U���e1�F���bo�/
�n�ϻ��-�w ��"W��ރ��ns�f]˲�n���Ѹ�Ŝ�	f>�;���9m;�<�4n�Z[�a�{�#��ST$:�>�x��O�rM�`?}�{.��2�c��j����[���,�ީ#5	�x�s�����@�R��j��e*ۮ���(] ����ې'�6�-����e���W�`o�l/KmH�ɾוj��Z�1����C2���wc�u ۿ	�q���ee�up��P��כ�ymek��L���\#Z��l84�(�˫#Q�*Ld���W2jk�k�p�R�m-�&�<�W3"���@���D��[AT�\vfǋ�y`���+����מRY���*
"� ��3���Am�!u�Iq�v�����A���7��m�s�S\'� �Ο7��f��]�@���4��������;/���J�ɡUaVn?�z�ܞ�W<���\�ͮ�-t��*���{vg,���f]�	��F�O�q�4w
��{���%�8�eF���{��5�^-��d7#"�U�R���n��C���<�G��Υex�����YM���N|y��p�A-�> ��n)�s�����R�}�՛1{��uRb*x��Dfr[�A�3�e�k;q(&$���ɍ�Զ%��ν�#���8�����J�_'�~Ǽ�w��ۙ�p����3/i�q*688M��h<�����������Q��q0{޷�OiU���v��a7���Y^)t�� A�h�v�K��Nn��ms�M�) ��@� 6�L]eę�m��en(�ܶ�)1K���^ �Ο7-�w#/����`����PDn��m]�Χәu��Ĩp�_}-1�F鮾<�m�ao�]p�s��C83��Tz��H�;�C49v�xF4՞��Mj�s��ܒ7)t�Wz>~�#�� �@�� Cm	-��&���r�T+4Ѫs���c��y�}it�s����'�͡���	����G.HFV
��JGk\�B@�v.Z���f��k����1�g9H�-�� �ڛ�ΛΈ�춶)1K�C�L���/�` �v�H-Ǜ�@�܉���1����_t���U܍u�ӗM�dJ�� ���H#5p���3����>#� Aހmϛ�!��I��_cK-�+���I�΄ 6�����ŸG�{��nz;���A��^�.���ޞ�#�W~�G�'`�d<E�a3�����Aۑ ��� ��B���/M �v��S�ś��FG;ܤ}�� �E���;(��;�1�"��׻�"��\�.==�أV1,�u��KݙVム�;�j��=S��N.����7�ѵ� �e@D��*%���LX9��a�T��{�v+�JcKfI���i�"X:a*$F�a�ֺ�[��!�Ye�))c*�k�n�\��(��Ѻh�1	2�Q�;6R�氰m�6�ՙ\�����I�ֈUe��0��䷛#R�V�kl&]r�%g���Yk�ܷJ0�t��E+K���6����E�Y[m*�,S\%kmc�x[��gfћi��V��|�4�Y�����<{�@��)��o���n�e!Vp�̮Ah�g�״��#;�O�k��KƧ�dv$��Fj<��Q�o��Ⱦ���6�3N&)p^퀈�hIn2��YUQ\��ݹ�A{M��m���кz-����nJL�w�B���wx��uy� [�A-�$6���enE\��@�7�ز�AM��;/z�������h][Z�`27rg��PE�@����[����a�^��U����}W��-r�lA�s���A�hup�'<����_5��.��G�qW n�pE(�J�7���UA&J�JffP5hq��A���7p��ķљ��
!��<#�9f�?ft5$ڂ8�Km{�	nY[<��c�>�6�8�&e��ʺ�(��NҚ�6kC�����-��uTw�+���b��V���>�N3Tj�.f��UH���F���?Z�}��I\�xġ�<�[A۪�x�_vfߤ�}<�/�@<�H ���W�%��N9�
���9w��Sڸl��/� ��@���H-Ǘ�A�C&���ѭ�������m��u5Y��b�(���^��O@%U��X%
v<�=R��8�"�r$��D��;��}�kw:"��x���c�^!��-�R���x�.MK����^&O�A&&h)	u$�Lج�+�n�,��nU����a���x��tǾ�>-�Vkz��-���k_ TGd��iӀ�A�D�q���܉�S���<�Հ+��7�A]nmR}��{c+P� �k��P�ōl��Z�K۰�"|q���Ng-F�\U�Qy�b[ɭR7�!'z��n+��L�|J/����cR8�5��v�]v�&262^й3Q+U-��t���#{]�9���WU��p�-���|[Ax��O��Z��p�%����n�лk���{`	����u~܍�/�^n,���D6ի5��f��Ayc�u�-f��*Qpz��ւ�Dq�f���z��^�Ɵ��3P�3�m`�RY�3��:�A�sv�k1S+�C��z @k�[� �
�O_GD�n�K.��'����U��s�#[Q��mڽ!�n<�m�"��\�C<sa	��vgv�9'���B3��=��y�ͅֆ� ��$����b~�v�꾃�fR�"�1;z�c��o)�� [� mI�������Vk�A�>΋�^*y�#U��!:���C�8�貥t�(��qk:���d�<�Fj돧�>�V��d��<��Z][�}��:�ͮZ�\�n���8ɭmQS���έѝ�s2�ff_�͠�n����\f�Q�f�{����2�T# p=�ݎD��m�>9������9�ٮ�һ��L);9
V�������#������s��!��1=����M8�V�'���e��� ��h#�6כ��pN-��mUf{\i6�
W\8WM��.��1<$q� ۃ2�h��v�� �uǐ9����-��Ŷ��Vo{eKݨo��(��� �nD��"mm��Ő�w �]Ƃ3 "3uy�3��W:��;*&##��REL���y�����Hn���Ȓ�Xk˺����;OS��^��Q�I|fW�#�-��m�����x{T�'G��$f/S)hј{:��YE�9{Fty��i":e��/�9�w�Xu�o-��+E;HF�oc��f�f�+ƈݒk����XkDb/T\�	�ݵ4&��Hb2ʉLo�n�7Y���b3U���8�m�;T�"�f�=�a*�,�]eQ�va��+��W��(m���f���Lu��kJ�Ŕm`鐎l�k�X�Ƞ����X�&�HVӫR�Js�q,n�Vkk�Uj�\4�c���?��m��(�n�tN-�E;G�]n�*�@b۩��M�r�c���s�e�^ �ڴ��fvl�::�C������q�Z�$ղ'�/[@6�A-Ǿ�T�M^����K���]n35���QA;ܤ��q6dov1�H!��t �A�����Ԍ������p�;z���L����D6�|[^n(+��/�rJ�w�E��\���6�9d::�C����e���]�0�Dw �Cng�� ���&s~ʹ!彘�x�O]B���=ܽ����mP����5��g�a0z T�0�$J1D	Jsm���UH� ĒL� |Ys����*����v
X�	h���� a�s=w�7�3� G=�O�mp��mIqu;[�W�)����aJx�K0b��U���c�5zqn��.�ʷ�S5�4��J�c����2�6lhL�,�~�A<�Zu�m�u��::�F���Fs�%��w&L�00�̂u�7s>>m2�.�`ՋA�fVu\�t���e���v��p�ڒHC�J̫�˘A�q�A
u|���Fe��L�n���;�������d��h"�"	m�!��g�<�^����%T�zxr{��U��� ���	�n�Ϊ�}SF�l\Y�ty����3��*�^vB�͌��������VP;�H ��n������+�힛����Q�8�UU�&��"yҲ�P@�� ��Ԃ��p"�w�v���lh5q�p(
wz���P���fP���1�����gu]�vbx�^��>��A6�������ױ�`�~Bb�j�t�J�I�^W¯���^�6��9ˈ�R����`��]9v7)��NY��uR��J�Cc�H���WF����W`����;N����n`oY]�]�oN�s�[��(1S�}���x�	���Etz���g=��!9ub��y��X�ٹ�uػHi�VTh��7"�"Xy4ZѪϙ�7h_ hTtv����lְ<2gY�	/&-�p �;�ʾ�k�rE�|_'�r�Hl��T�q�Q��e#u�,F�gF�kȃgg,bB �.�6l��][5���EwWd��4Z:;��AՌ(E�o��h�wS�'h���H5��9Y\��ӷkNf�z�LDE÷x:���o; ��nJO��j�R.�vr�v\e�08ij���nd6� �������Vv��.g��r�0�{p��k���u,�td�sT$čO=b���7sbh=[�rGܖ�-�[k��"�tf��4!8��[��b�PV"���]�рC�W=<6k,L(G�oۣv�d�E�ְ������R���.��݌svEȐ��F�2�HP)�@�����G\֡��j�*���=b��w�	�c���c&> ��}k �뻯��ڮi�i+�ۗ|)ls�o8=�w����X),����m$�α�}k�zXr��ZI蹵��sQZ��+*̼�(�
���'O�7�(�ڹ�6w[����3�\�+sW(�k����<�o�[�ە�Th���ۦ����6Hhؼ�F�W���k���*����h�Z2U����lZ.�ך����ž3ݶ��T�Pn[�X�d�M�������ƾ9�W-���nn1RQ;��o�rѷ�# ��ώ�h�>��,cc��ŵ�˔N�F����$��Ja#�߯���~}}㮹��Dl{�/������D6�D�W�Ah �k�Auz����u��(�A=ܤ���;S�\���\w�'q�!� � Cmy�CX}Ϯ����f�Xyw���ȅ.��3�=��1�v'�6�����L��a-�2���	��:m�l�fP���Wz}��ڒ|��n<�m�8-��}]sSR#x!\3�&�TE�' A�h/۟	�:k��wj����3�ψ�Ay]_-鵺�u;J1@���h"�e�[�Ъ1�2�e��)"�v��$��������oU,��gEz��S��>�,h Cng��@���{Fl�2{%q��%��V<��<ޫ�b�H���9�OL��&�d4]��+�ټlg[τ��f?���`OoayyÓ��Vv����G*-pR����o�`�`�����q�,�8��Am ۹�p�cAl@=}&�_@�'w�6�^WS��28�{�H#\p�%���<��Ǭn�~��-�`��1�#�����2�ֱ6��H�ۮ�a�Lʙ�ш=x��B@-Ǔh!B�8w��j]O�e	/��e_da��^#3dO�k��6ԑi劘��!	-��T�x��y��R�����;\��Q{�E]�눪�qGc�${c�͠�m���7l�]�W*�k5ݨ�����Rh"�"	m�6�"nF�7�+��p8��BA{��!B��hk�_I�u>S<$�I^�_t��Ϧ|Gj�y [k���/a�WhR�w-o���5��I��"7�Ÿ�D��[@�i�y�l�оd�V䲶�c`���㺦�'9Ru��5�(��NX�U_M:�຺��xM���f�����SL}?�x�ԃf�`q����e\l� Jk�LAF�fi�]3)�`(.ɷqs.i3JuA�+{{j8����h��Y��a�7'S.L$ ;`�E����H[2aHm����u%X�e-ٔmlTљ��Ye�M-����vp�͍i��@�J�4��c����cƻ)�]��9[�mՔ2����ͬ��v�Uź��c!Ε�2�A�R��ZJ��jJ�_'�~��A�D6ץ�������q���D8�,��	��q0�, �A��[jHm���vŒ�!��B 栨Uծep��7.��g��Ё6�6�h=��կVǨ�Rn�D[i�D.Օ;K�]�5�r���"7���{\�-ǐm ۹�q[�m��ra�R����U\f�}m�uy1�'{��"��W�Z�{��Du�Cp-�@�r$ᶨ�X�(�'cvitth��7.��e=����܉�m�^��n��`GDǐ�1aE�
&o{r[KE�5g*��f��b�i�d���H}�E��y�Sm�}--�w,V���[q�u��9��!�ϳb�n m�7�L��R�~fL��`�z��l�nX2�1bWh���r�Kۏ|��,� �^\��t�%ݓ��Qo+����>�4b
ܮl��d��'{���-ñ��A*����^n���D܉-�6�t̃3i�1*qdl1ٶn]O��	�^!��^��@���aE�蕊�A� wc�ڗ���iw7i��"7�%�=[E��a�=��#9mȟ7��۷=p�g�n��az���qX�l���3=�{��4n �[k*��6�e.YǛ״o�VgrU��1�h���H���`�L���YtV1"fR�#u�� '�"Kp� ��)]-�;6�˩�B-�n"c�#u��O���n>m�#A��j"̅��} o5oǮ����j��n �ּ�@��ɻ��
���r'��Ch�ϋhwdt)�Ĳ�����W�z�|�� T���J�b�+�h��9+�t/Ψ��v�j�'d�o;���7�m�4%O7wo�'&aǸ�r���QڐCpLV����Ȑ^��
�M�=��gY�u>��8�Dv�ru��aڼ���/6כ�e�Q�D����x��]���R!�^n>hIn͡Ss����|���>��+�*�:n1#���R�mH�V��ZͲҡ-��r����!�����{ￏn�[�^3۷=7�G����v�r�P ���آ	m�!��p!�[ِdtown�˅�jP������7.��3ސ|{��͠b�����H z�^r�h"�#���'�idc��:mns�b�H��[��!�>-�Aۑ"�!gvJny�e�/�����WS�c���.јq�A�� �t�7Zg���M�+�����n��0�V����(�&�u�
����wP�烣hh�v��i�U�ڦH�u����S���pm�n-�#�	Wa��4R�+t���n\Ϧg�����܉�m�>����G@� Ж�3enD���ٖҵ��XF�f�B	v��ϯ��e��Ԑ�-���Ԇ����v_Yb�H�!ʜ���=s�s�7{"|w��6�!�"A-�#&����pq	��ώ��o0���F��	����-��v�g��r�Gj@�p�[� �mC�}JhD��4�N3z�ә�̡Ǻ<� �s��"� A�p���L<���RA�A��-�ܻ{9k����D8�d ����Q�r6���n8���!�"A�D���g!����b�(m�j�oe$n{��� �pn��it�n-pEl	��1�{p�E�&M".����Y�bb�d�ʆDJђE�9�d"�Y2���Vy���=�|�[��ie��L�� jҝp�\��8�ԍ��x���ư�Ζe��Gb:ͥػ@5��:�l�pp#AͷMa�̢ـ-Z�6����&�Rr�`X�]���ډ̊\���m��X&r�͕B���a����Y��l�K��$.cIil����R�H�������-m�h�3�j=���V�ά�����=jpϴ5�\:��e�j0���j9pU]��{4�eṫ�. C;dIn ��
�1}���u�>��T���Cr�=��^#;�����@-�$v��k�Ķ�7���>y������]�5�D>��D>hIn3Qjz�3�h
�H':�^!�"|@m'H`��&����ut�v�$r{����כ�Qm�7hMŵ	�S��]�Fnϻb�!�
�Q}���;��^���A��&o��`v#gB��ϱ�E�D[k���@�Ƶ!���~c4�{��ߛ���CG���9n<�	��EnUdS��J�*�E �[ա��-�a��m��L5���,�[+L�WicT�ƶZ�܉�m��͊��[Β9=��V��y�Ҭ���� ��RCi�[���7��4������Cj0���x��v��Y5[H*m�,q�"s��2�|��3N��_x��XV�d0�'�icLR�v/F챉��C�l A�T*h�f��w��3(q�>Ƃ �߹��s[�rh)z�(f���G �H�پ�髇*&u^�ڼ���$C�����ϛ�!��6�F3}N�}�#j+ce �܉�������s}{\�Qp��{�[��K�˄}}�|Ciy��܉�n0o9uy�q��b�'j#s�t_;��^��A=мCp�|[^Û]¯9��*",�3��*JJ2Q"@� ����	�j�֥��a61\�������w{�������~Ȯz�CElc�IB��k�tyc@6а[�<��N�Nץ�Ur^m��^�;�[P� �h"�Z�T��fwT����� �^n�-�D�Q}+c��PX�Ŏ���PY�N�ц��f����AilOؤ3��[K�~3���[��0��9�u�jsz�+%zfzA�#�s>n<�Q��3�k�Oz)zE��Ǒm�4�y|:]�[!�@�p���q�8�� ���6��	n ��6��5]u�\�
ܞ��w6��-��|{�zy��q�[h[����:�JRaL�R�T�e	%�� MFlչ���0�3]�+��>v�현���{�D�T�Ƿ���U��̡ݬdػ��� ��@��@������&]���ڟf]���vUC�[!�n ��%�1�DD�mH�� F�p�!��m�O�B�wm�\�dTSg'��u�k�E�A=ܧ�s��q�[j|Ch yh�љ���Ȑ[��Cp($hoޛ�qW+�3�=мDxNp����8oJ�"`��]@ҧ84�hC&r�T7��o��nwP#�5�A*Q����S��&�����<r'���qD������3�0r�۸qٶy\��b7�&��|�H-�7 �*�U��E�ྡ���E�e�FZѴKwR%ʸ������ 왙��k�K�Dn�D6�|�+y�����-�����c��ZZ��@-� ���p�������b��[÷���U������q��m�ŗ''foе{*(��jH-�7 ���l�@�b̽=�W���P:+��R!�BKp�n6�H�����]tƂb����	R���]��:�j ��� ��ʈ��z������!���p|)�#�vXy( $)9c{f�*.�zT��}1���2������ԫs�0���9��+�:v� (ܣ��@Q��^���F#�~IN�����)C��~��:?-/�����1�B��A."��E (�?�( �Dt]"�3�"�����a�II8��=�kҔ���ю�jz�'	�Rץ�>��~����/s�=�ǯ�a��؞���x�D!a����,=���4����)�r�Y�E/{��^��@K,7�p�qӠ��G������� ���b��{�D�zP�Oq"$�KgҞ���}��4���?��?h?����?�->���=C��}?� �������������� ��a���x>�솈'M�G?�=�� ����<7 k�u�����X{}����X:�O���9rݳ�A��z�i��]Y�n~�rC裁P@S����O�Xځ�MI"�|��z�U��'�΍	���?���}������	$Z}�!����q�5�����)�U����{��'�=T�k�?׀��?�>��Q�?�;�~�������� �
<}�@G�lOx~�=�/��������rh(��{�m6>	JPt)��Z��i�����p>���P{1�=B��C��W�~a��` ����E�3�������q��0,�?�
Ϲ>�G^� ���}`���O�?�)�p~�/�)���6�?`�W? �% >��<���(���\$���[d��X���d�Q���K�����x_�g��	��Qh��_9j��A�)����pi��O��r( (��}o�}���ާ� (������  {_���0C�z�C�i��_ �'��}�����ܾ��g�>�@�{O��a�>|�~)�����2��~�D����@���|�o1��FO�Q@����1'� (��<?����	��{Cc�����>�}j���}�^� a���*4F-�M���?�!���= r?%< ~�����?y��o��8���=yo���#��:���Xz���L!�tC����f�O�%=:�s^�8H����|�� (��1_�,? ,��p�������{��ڂ (�K���^@�z)��4<�3��p"uu����r��H����P�o����O��ܑN$���