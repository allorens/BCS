BZh91AY&SY&��_�py����߰����  a{���E  A�   t��
` t'h �  	 
   P
 �   ���1�hJ���ӏ
 ���]�	D(IE
P�� jw�{��]n�u�]�G
�m�:�v�lv�n�%�8�}��+׻�IE�Oz�g����A�}s��q(_x�=�i���V�v4[7�"95[�A�	�
�F���u���T� �H�;k��`7p���=Cl[�*0ӝ��V��[h��gw(�s��I��t�t;�ml� ]e��1b���۶t�Ӯ��]5w����7��{��۳.���!k]E�#����{�=���pzwf�e��w���v���ں0Pp �,0�����wn���ݓ���ѱ�f���w�׸S�=o`5��x8�۫����^��Zu�lt�5�Gs�]uI��wa� � ���n�L�Z�s����ݳ�����w��S�t�
���j��ws��m�xt݀ݨ�������m��/�b��  @���E$�i��h��`P4	� 4 � *�!��J��� �0#  ɦ�jx"$�Jz��4�0M10&��L��J�d�M       &�*JC &�i��0!��4��@�
�A4M4�&Shj���)��z��O
i‪i�*U# #10 M4�`@��}���{���zqT�Y�a��[�bl�\���(w��s�;ۣ���r����BH�+(p�.I�zQ$M!"�`�"v"~�~E�e!$H�sX��������>����6׳C�����%��Ղ~E&p�%FJ9��x��1X���=Z$I&��$N)Do������
d�@'��=2y�����o,vI���U��͙is6�ٽ�ğ�?g&���rf8X�b�L�&J(J H�(I�LQ?1��=��,s��g�ɉ�L,G�ŵ1ӂQ��$� �>AY'�P�H�$�Btk���&?�<hl�i��r�t�D�ω�D�3<������s�tOՓG���f8?`�X��b��(��ُ���G�`#rOȘIׄ�(L��c��L �L%�1�Ǆ�U���<:W���@� ���eG�z�x{R>	Q,��ǆ�0�=�����>艅��r�xY��&10���O�-��:r#���<1�1�-�r��#�G� a��x<Lyʞ�	����t���D�==�H�ُ��>��UT�ss#q'��xY��I"�(��P��O��&��1�a��$GY���H2c�&a$N�ra8#��L8Y�r!��tNx�'���L��!(G���Gc�	���`���,���0�+�0�9ل�gO�	cqd�`�&W�2��HN�\�X�\�(���(I�&0Ef8`�{���'���YBLBI"�L%��YB\3x�G��1�T�P��#
��ω�.a!=�a,�V�|�2>���H��f<7#�%/�)%�1��#��ft��,c&Ň�FY�xN�p{� n!�'�Y=.G�迬&#�)%��IN�t���p��#p�;�1����@�,��H(�	��	e�����ھ1':�k�Nգt�-գ��Ӯ�s	'�<�����;ȄG��0N��pN�L���Y�ع��2��Dt��B'����>&G�v#)����0�3&�ǄI}1������"(A���zb>A��=�&$�b:Y�3���ْΝ�Ѣ�����ӷ39�~k�'�a0i����1�1a��LtG!0��}�za�}�~���=�9鄳��I��=���C`��`�\�Dr<A	.aG#䲄��Dj�,N}���DF�0�'�GМ�D� ���3����������Ŕ#�H�I�5�D�c�$�p��Qd�&RQ0��T�Y�G�"EY+QÝfdG2&K*b�r<%�pO@�'X��
$O7����DQ��I �"Q�����h�L=裠��O�(y	�$O9�'X����~A2'����pJb!:x�Q)b&5�F�a�dO���%	LĢtO9��.#�t�9�$��Jp��F!<"5�pk���Q�
�Ĥ�&w�L���DH�"$�D�bc�)�K�H<KQ(��Ƣ|Q<��|�"Q2�Ė��CY��9��$���D�j%���O5�?!�q��(JyQS�'&DDs�>:%�O�?,O�(J{�%�x��pF0��{2�;x�ysi�'��1Ǔ?aU(Os�(��&rfN�%	�X�8q��w9�'\�D�F	c|*����"�/<ԴP�GȊ �	\��L#w0��3FfY����G=3%�I� Fa\ϾFٛ�?"g"��&�fj��D� ���c�����A!fi�,�g����fy"{2%0���Ly���e�DQ�A�Hfg��L��@��;6�J��U:u�]�کGUg'Q�:u��C�����H���Ώa8'N7�xN�ώ���	�<�g�	��͖y���AӌĤ%��-D��ע~~n%(N[����a�x�k�Dj;��"(��:KQ(�9	%�F3$����j'0}���ǉD�bB����C1(������	��b!8"tˏ3"p��S;	�7�(x�NDI� y	��2"&1�(L\�tN���\bx?I�~I8q����&�����{3)F~�&&��%,L����N�D>�ҹ�$p�tMexe�x{�}�P��dτNN"]GOpy&&	f\H�%���Y�D�Bp�(��K52�@�r	d1�p��%��0�	d��xIn%�_���N�0y�x$�@�|���IDL$�ID�牓�P��T#%QOН��x�v8 �|�^L�I(J�J��BX�rc8&D&	��"Ag�����JO�:$'���=G�&K<�,�$�J8�̈u���$��o���Ù�͌�>-�~�p�����sؗ;�Jн�>A�R;��=���	�&hI��N�&fI0�LO	N)�̕�8��	+3B9�����D%�Jp��=:��N$Gx��0�>y	O���g�bw8R�#JK�&�s��&VX����-��ש�5+{�f4���]Gwf392��$�H�DOy��&��,�jf["����l���ǹ	�'F!����D���JP����CP������=0��"~����O1�lp��D�7���bl������$��"�Jt���G�J�D�y��G>�za^���-�Jx�Dؖ9�>ď��IӴ�� ��/鸔�&؟8q��u�JX���ps�L,o�=�Ȉ�I�>�I�,�,��{�X�OT��B3"�?!�0���D~���"7�1�)����%[3ÓId�p��G����Gv�-:w��lM�x(�D��/"S��~���D�"ȁ<�%(E������������#�'�$���(��2"�<P�YQD`�z��;܈�S(�* ��<p��D�AG�"�a��Ν��rYx�'r6U:=����&�I�r=�p�&	J*�"a<�%��:�ŝb�x�XM$t��Ĝ�9S�u8"ǄO,�G��L$�."�&c��|#貄k�)��a脮�Ñ�Ƚ9��M���Itd(�����
�Ԏ�?J���/���}ҏ̽Eq8�#�����u��5t�z�CfK��|��}���m�r1�]z���Q\a�/���pi�r5�Hȋ����ձJst�cg����¸gWos��/T�9*������奃���̬&�7�۹zw}ۤ�(t��T-���0���O�'��b��`��V:WMlȏ�s�tǠS��Gk(�ׅeh���6����W�.b/���YӺ'a͛�S�� �TzU��ms��Ν��]��;c��z#Ӱ�	�e�2�
�3Q�RXI޹�/1̇c�k�w!çv1�г��erG��;�k�?���l��������W�؎W%�v�DI�|�{�/^Lk��L��B�K���՝'�w�W;~��>x�8�g�����*�_}C;�+��4�pE���^7<��_ٯt(in�[���<��0����Q���yq�lh�4�Ʈz�(�e����w'��ɫ܂�NbLg����ٗ���a�M� 2m������8&S�*�2x÷�BAo��V=�kf�O�>=���;������DM�On4J����p���+@�9��dc��18SП/�ny������u��>��aO�u�cY�&>�=�{��o��]L������A��:Iz�2����t�����t�	�c�+J�1mU���'��/�;h��ɶg��?}�X�F�yq�:ܐ��!��k��s���:�L�C�y�ƌݱ��w=��6�kWp�J3�Zw�4�G�?g]�:c��(F??���Wξ�GE���$/.���Od8�����3W��(��hBwf[m�}70�G�5����܄��*���c=�61sf͈�w��:I���p����szCP����=K¦��t�y�|@ƽ��MUb�2	V�����|ʭ������TF�ю����i��'�3�w��̈�g����~�*����rsj�GI�g��9����d1pa�ս�6�A������ݮ���s�����g��Y2<?��x�΁��1|�z3��~u|��~Z�Gc6�|});��G�v��'׊���p9��}����b�*��=wG�.�ۙ���B�9����,}&��X��[���{�ўYޝ��+=��O�C_r�:^e���sw�o�Y_�^��E���;I%��N`��A]:=���ܧs{���:S��+��Ic��a�j�zo3l�n�u��m>F��ÿ*pB�W�s%�D����ʟ�J����OH��1t�*&�C��.e�Lr=w&=�ow���	"�����P����-��[�C?����;B�Ű�hȜ;�ӄOݝ7M��r´��ȧ��Ҟ��Љ�����#d�C昘P�6M����ӱ����NH��z�6J�a'(�s��eac��=��&Ə�Ip�#���~���F��g&F*�}[O�����z9<�Pyx7s��/)�º���`EC:��:a�=}�I��z޹�_�zV�a���w	�����[����,��=߽������A���ۍpu�M�ǻ���O>6�l=Ɗ�>!K�Ϸj�u�J���yʧO��Ϛ+F�^՟'�b�f��S��O�0�<e��Y���I%�IQ�\�d��ώa\/�d���i�����ꛊ���޶cy����ٹt���>Y>t؁6b�}�N32d�7�M;N5��G�k����qM*��:���=wL�J }���'EǸ�q�V^ۘ$��4X�¯�:�ۄV~Y�9zǾ�?n�ު�U���j���3Be�~=m'�>�t�X�"�o�>wb�c��H�e�>{�������o���^)��T�{	��'Ot,M�$��c�˶�/��f���?J��Z~'���ː�gi���R�!��aK�ߏ�� ��ܞ���z�M���ӻcs��zrEn�N��i�|��|�~~�ݱOx�_hٲӆ��v����o�\y�+��O�����w4,>����a6?��̵���7����1��f��|�3��;n\A=�U����\��v�{]	�|O�=��:��Sf���s>�}��I���.�5�`���+��du�p*|��i��-�*��8}�p����h�%y!�֌�$�u�/�[��ϻ�o����M;}����Kzr�iD��1u�ҿm�<���E-Cصe�����Ǖ'[��[QE�zv�%}�d�Ni�;\�R�Ṹ�ڢ�ɺ�|_o��u�۟t�Ǿ����.=�=��Kp�M8}��C;;��`m�Z�`�|O�9��{�f�zfc�z�3V���W���7��(עC0l�)[�fT^�a1�\:Y��nۂ},Cd{;sk�U�0�O������N�!�	}�������X�O8�itӘBi�����G�Y��d^��I䅈�1>��Y�WXd~0w=)p��"��۔�AԎ�>*\k�����jZyU1Q��I������?9��>���l����'ϲNݽe2}ͪ��7c�Mp��E�fr3C����!Z+??87~�-�<��s=�+4(a΅�L*�65��,=6��"ߦW�$���yL�>���m��4t�L�Ύ��>�7��ͨFV�ߣ��Q�Lqt�I(��2E�Z�l"a�0���c�g�t��g���7����'pJ���K;2˚�gk�=�V{g���_F`8��;LLf;����Ea��a���V{��degLc˷�ۥ��;3	�E�i�31d+t��v7����s�}�!��S2��q��n>�-���$P�]^%�Y��~xd���ܹ�UL��~[6��?}�
��W��&߻:�Ǔ/Ӟ��X{g�����gc���wp����d�:����>���C珯���(%�;_ek\��a? 	酚{p)��=���E=;�w�/aOK�e������h�C�}�5��'�Swg���"�a��wP�d?��:�+Q��O;�~�~�HQ=�=��Y����fwKO�-48)�0k�>B��b����2�<45�mv|�k:�d�;A5�r:wNH��z]o[$�y�g�6��D���a:t�%�p��*ܧ?�2y����n�c�My:�8�*�팽���vc�9u�g=�cgbz��6�N���p��t.��R�kR��2������s���|�_�:g��g�����n��O�j�=y�vF&)U�k��o�'v���� ч�N��� ��^��<��V<V��xp���o��gl�Ӫ6n�M��+���ۓ�U*/ok�m�1��V7�3��~
���oWb��5���JF�[J9[�36&3i�a]��42�q���V�ZF���H�(�.�N�L%K\�jE�X�k]	��#�;��]F�W�D$!!Cj"̄@�p���t��,H���tSNEt�d����n	v�I��1GBI@�)#H�O��D�x��
I�j���D�K�O\d'0AE@�Q��V~!-[)����x�&�j���\�ƒ��р𐤑�e c%bd6S	��}W��=@�\%�I0aa�bp6�G�D=�xx�ax��vpM�\A&	$Pdr�A�!�c�2 ��Θ��V�%�gu�MD�`RA��8-E���I16a��B)#L2�h��D��$����D$�� �k�"�?6{#"*0�j�*DCH�T�8��Dt�u/V�7Kӛ�+�'(�jHϡ�|����G=4�]tF����3�K��@ �����F�Gt5z�H�]څDI"���01� �F����l�r9��䡵�~_�ҧ��&Ñ��A���F�e�^l����Gbl2cyP*��@�瘇NP$Zl6��B� ���
 B S�G�!��>0�1�c1B
��lD!0��Qh=���,�Y��B���J����M�Z�����K�c\�o`�$� k$0�,�b!�Z��;�k�P<KKE�kA�*��p&���$\LBAq�8�$���(�G4���pe���a	�������XRFI�c����Xj�	�BA�~�����D����D<�+���x6A�2� c��O��*�5�~4Zx�Gd�%�:km�+y�-�0�PB�(�!dB'�D6�X�|�E	T� B�T�C��ܷM'ۣqMǂ�K%��@�Y;���2��c��h���^&��s�i����n�a34�B[n �ump�ۮ��q�fB��<`�@��S��ρ�&�֓�g��L���J��~�8�҉���#���G��" #�|�xa'��@��P�Y��xO����nv�qDqa-�(��K�T��L[Mh��&�8�347�@$a	�B,�ģ�)|���U��@%hP�1�\�\�Ҳ�d�����se��q�T�I�C���^-}�v����<Ro�?���_�����i8;�I������ỳm�߿~���ޯVUqU\aU_+J��|�x�Ux��}�{�_+J��ZU^��YUV�Ue򴶼Uz��U�ª���|����">��!%��RI����򭾼EU|�*Ҫ�YUV�UUQUV�UUmeU_x���*�
��0��k*���EU[YUU��U�iU�;Z1		I!�DI;��]����UTŕU�^*�VUU��U\EUUEU}�z}�*�ª�"���*�Ux���h�����k*��^-}��}������n���oUiU|���0���^*�^�Ҫ�YUVՕV�����^�Ҫ�YUV�UV�U^*�XUUŅU\G��{�ｮ�Ja TB, ,��[��$��dH�RN]=i��"R�U��-�g�v�����8�&��'q��w�Z��ۙ�;��7�ol�ٱ0����ĉ�(NxJ8ID �%	%��ı0��L<%�&	�X�<%�g��J,C�P����I �$� D�<'D�K�"C�uh�Ӭ�2�#'N�|��%$��"""bFI"$�BpD�'��a�'D�,L,H,L0L(Lĳ�YQg�	�H�'D��xL>m�M��]FV�ٴ��#�����s����*CT�[���V�V]z��>[�V�?e6�	�î�eٲ�mn����+�)J���$#Bm�Ep4�A6�l��C��[�i��d���S�$]��06����3b&��f�ɕ�Xۥa��������[=1|�[6s^1�F�6a�c�T:�3d[v��-Z�f6��h�ZAcF���e�6��ebo�z�#�j.�H7��U��&CK�YDĠ3�,aaUA��cd��H�Τ!����h��P�$�
@���p��CŘ�R	�!�)�C-�`��Ą%�D�ʢ�J��Fcq��(�D�fM��|���Ѝ4��H�h�@��F6�4�(��R�&퉶[1Ipa��0�`�H6XWif�����v#H�2٠���.�ԟ�;3�k��}��R��g,CI4�I�[/��e�K"';,�Ɠ�`t�P�K)�L�ih�i-�)-��n�ֶ���E�.�r��&ID�]Ik)s�V1�\�s��dEm4�S�G#��
a�,�S������eaR٫��(�]���eٚF�K6.X̔��8�õ2ܚf�؂iwK5�8�%��[2�и�R�hJ8��$B�"6ex`�B�p��Yi�	B��H[ ���0:���*�=7���5����t-��X���6aPˉ"a��J�BA �h�m�+afZ��&�+���z��"�BV�����.�b�҅M2�a#o.S�	���$��%B�����M�{��)7$v+ɶ��k�AvcS�p�]����k���l�%t�^N�����kt�[fN��,6#KآT,F@@�Sh��Ɓ&�-	N�g�g_�=�F�L�`��Quq\#�v��բ�eǝQ�BL�K1B�h��;DjX�r�;���s[(䮺���t�l�!6%�ٝͺ���e��5�%�����e��k�X�-�/z������O
��!��(؂D"O��J(P��1{�h:ؔ ��S<d!�h�1X,�5Nj��g�� ����~�ww~ݍ��������������>7wwwn���ݍ>>wwwv�����߃�>����:i��a��X����%	Ft�<'+����\�F����U�2:��1��k	�G[\#E�d�rg6�3^�[���ާ]�)8ح-�Yrl�ѢE�#f��Y�B�ķ�C%j�Z�mC@(e�Nl��]u�Ď�~gm5��]eq�),���ݯQ��F�6�� ��V0rݳkΫs�(�\l�A��P�1��!��H����ڕ"�m�[m���zC�� *>�rƈD���ř�x�(��eP`a�X���h�:�ծ�U7yxk�ţRPh���(ǖ�Ou0l�i�[��U�+�%"�b`�5%�ea54��c���E�l���aF��a�h�����ю�Z�ɼ@P�h+��(�����d�Yb(��C��(�!���	����(駋4�?&xN��&q�m��Mݳv�l�;��6�XQ�V�R�ld���,4vs
(��s�4ɵ�L2�;�C����e5Uӹ��A4Y��(�l���vt�(����R��A�T�7U�i�,3��}�\9B�FN+a�i��(�gL�P��LClX��-��3����d
E��!�`����0��tD�(��'�b �J�x�4�Z�1S��� �7	ѫY�8^��	�Xhٲ�0��D�/u��3��V�>a�猷]�9�A"4!���L�5C8�	3q��Xw�Mʛ�0j�`6�Xc��1!�ɳ؇I$��i-��'(;�A���j����a⨘��,�����Ο:p١8"P�a�L�w�]���Q�&�*U� vt���*f��8jN�p��@/)?p8ǹb<�FC	QBCF���5WpƘ��!�A��;]�������y�G��;iZ���b�ٚej�_S�8�qݓRJ�hĠ79�ƴfj��S����'���Q��0�D�Ή���tx`���'$�m��+� `���Ƃ6�J
�*¸.&�|�{�M_O]�6��YF(��A8�q��(� ^w�Pý�%4�U�5�='h���Bk��+<k3+v�9����xM�I�,��.���l� �C���R,��P	��ntѳ���X���f@��DU}ql�>��=&�����j P����Z0iS������a l�G��H
G�|˹f,#3�&Z)F��Z��T0nk�j��F���I���e�m�q�]q�N��:Î4㭮�\3vZ���a&���@�
i"��'C�V�n?Uj�>ju.e��a]H��@٘_�UI���.Q:Fڦ��ͮ�ۯ��N����[;�$��j�K�p��1�0c��B@�-,�sU0�B�RٸY��c)�Gԍ"�v]�jI�ޓlD�_�A��8&Y�����%�,��'�6o����b:k���
L��\�e��В!�=�4��f1@Z�ɳF'��F���1J��Us%�N�x�=�tA��|RF�iBa�����)2�@��|�w0���T,��[m��B�F�e�;$��Y�it�Jm��k��#���p$|(����o(���c9�r�+����#(|�O:X�a�&tN�%a���u|�)$A%�
m�  b�u��^��}�N�����j���j�1R�c.��aS����z����b�Mڨѳ�"0Ȗw:�$U����!�a�0�.&OC!������a��MLgZ닗��HK�ثJ�9�{:h76�;<`�����X�,�""&pN�%a���ض�	�J�BL��]�Y��R�v�x�sS3��e�be9$b50D0��@e��*CBr$_�9"��
���"���2s`�R�'���ea�oL=ū�����Qz�kE��zR��F��ГpnOt�W(�����C�̘<f�
<bP��l.ו[��0�&!��]�w&�X���є2�Cq�=껫l��"�&�fg��٥���lV�>��*YS�`�!8da��h`A�%�K����(��<a�"&pN�%a��P��a������r~p�:q��}�bV)t�]� ��8���

7��<�D�Ű*~ʷu�\�W�tpzP��(��<HPo;�s�t]��$��e����}�B��%d�p�J0��t��B�C��E�/$�:��}x�gT����q�S��s�Xi&�:&��JF��PX��:�d�S�P�I�+��<z�o0�^///�/oi��F�4Bi)I)��F�����Yf����t�:JQ8�e�^������O�_�<�&̥����co4Ǟm�>�#��1��e��O<��yk��<��yH���KKO"'�O/�_�y�u//�\���io'����<�G�b���<�'�W�4��??7���~0�h��IM	�I�4I�'
'HD�!8N�����	?�J�I�8�1s�lZ?'��=���������x|p�(��U̧g����0a~av�[�"y"<���N���׻��ϳ���ǽ\?��O{���MBB�|���,�b����P�i6��gsA�tw֧��j���s���y[K�q��,�GMwc���׈lѨ������S}�I�L�$��(�1��Q�5W�ћ�v�{ޭb�<��Uڡ5�79���9U�?�d�'�ϳm�����.=�o;�������_������3��}����wwww�������www�oۻ����̻��4���if�i��&�&i�M(�N�O�#%Q^UX��" d?*(��C�C�8�Z�Oֵ�Q���j�m"�2A&����><�P�DD�JJ!�*�AH}�J>i*��3�Щ7J�*�f�@ �=�f:\9% &ٰ�Y�/�FH\
���haRR�d�v��%+�DB�J���3��,2p��P�@��r�fZ��O���%Q�{�];
ЉЩ$��4�M��b����HM&I�j�z��Iں8�"3WEv��`s�5v:05vX}�0ܒN8p�����X�i�iG8&0����C$�#Uڦ�ʪ��������/K������LD��0�mc�)Ѓr�**.�D)��,Į�	�	���D���� >�l9�Sr���b����%+tT�J$9ϨTk�]UfbL!U�B?R�����R�*Q��7K�U�r��5�.[J������[��ʝL���ᑖM�1BɖBĩ��H��5%�u#5O�Jm�Z�)�!�b��b,�B�*C�h�,��tK�#؆Cb��ZM��d' �pD@�ȈWJ��T�Y��*	��C��q�矜<`�A��4ҍ:pD�Y5<֯���*2�|)L�x�a�c��(��Ek��h�6˭	��N2�BP8x�4+l3��@M��(���L���i� ���hE�&��2�$�֋7�,�����s�t��>�P����8pW{��A=�z��a���iݽa!���pҺZ(*ð��2����2�Bu���#ȈW�(�kJD���a��H	#
*�241E<���e$���Q��I�T(4	�KI���!`"�4PT$X)�0B�d(���FR�T�&�	B@d�t��`Cb"t$�LzPZE�`�2A��%����Q&� �>·E�RJ�4B�Б���д��i�Y;��	�%������pDLs��x������¬�����k�*�'����!Ҋ4ɀ�إ�&*E ���Y��DhA�J�(��KfU%Tc*����R��eƞy矜l�I��4ҍ:pD�X�r"�l��*�"%�C�p����M�C �aR	U"��d���6饶�O���.v}n��FFN��������Q%RѤD�"�;"D���BRI�
�H0�P5��[���B����P��d��eW��4�UB�`18"2JCp���F0PlhR��@�=Y������2����K3�C0ѣ����Na��Mq��X�`|!A�;������T�(�0.��C&"jK� ����=d�@a��������d(0QE'�:Q�1}��2Â"%ʣ싛$�!��K�L�>�kQ��,<ۏ�??8ۮ�[�2��<�.�ۯ>MH�I��f�,GI$� ��@�h��)�^|�⤖�Omh��:n�����˹��#O��ҥR��TIb���E�0!L��`��(D
H�#"��Ʈ����)�D@�����%��'e5eVO])��2$62|%!�K�5��T��dDD�wY�>�B�I��Ӣ��%�8ȔQI<l��O�%�"&#	�;�\5�
�6!q_�*�##e����ș�c%�7CQ&EJ%�0�����Zĕ&B�a��bn̲G҂�gD�)��I�2�,K%SB��DD.FJ#$��RhB���*�P�ȅ�r]5He*����g]e�_����q�[G_�[�0�H<<0x|4d$Z0���'��#T�RK�`�}�UDFC�&�B���UJ�13�. �Ҥ؅�"A�h)#�!bB�. \C�}sBX���Q��l_��5��ⅲ��=;�)UF�MP� T���"OF_-�D&�D2��ĉ>ޮ]�5��TZ�-B��u"զWJ�lVcx�>�,R����Z]V#�9H:�m�Y!��T%CI�-B�zf�!L�dI��-I6fP�`�\�X:�暨0��AP��c�.�m�lh	�0$���,j��J��B"B��d@��%($�6�i�mG)h� B�5�`d%P�1vE=5.�!���H��%V6����~q���I4ҍ:pD�YɏT�2G	�I���2�V±�3�BdBA�?�rP��9�ڝ1"�E,�2�Z	5�B�բ�Q�x�|k\6�Cz��8į\�P�Kf8�Y!A7O�I$���
ls��{�\��d��!���$Aa�[�"H(����9��mG�r���$6�z�ab%�mxp��m!���^��	���I-1
�@���FLM�_�?W��S1�5R��|ut��eR�ԇ�a�'S�YP�abFM|$� `��E�4PnBб�t}�vU�M�4 �}E	r�F�2�H##e 5RDAd��,`�����1Ć���'���8�>6b@��1d2O�)�3TlC����۱.���m> ia��DetZV+�%-%.�
E�ܥ�&���[���c|d�	(�EH�LQ �"�$�ˇarL��Vh�v0��a�����F060
�Q�}V^'��Ϫ������~q��~q��'�I4ҍ:pD�Y�E��Y1"-�#FP��I$2$�^T*�"�(<(<Qvq���]rL����.�F�s%�`�q:!�SY�Z�$Cѿ�����
Z-�86Ş�Kn�
	d�J&
�bf|�a1H��0b�3�]�
��&m�-���첈�'�%����c�Bۅ�c(����$=%Gx>�{���n������ce�X�QEˡ>�ܢ��-�=a�f�G��y|єTBXF���<�.U��Vml>�aU�y��4�񇎈'�I4ҍ:pD�6W[��ƨ�[z���x��'ơE#�(j|`>��'��>2oZQe��b4C�&��d�m�jܮ���H�����LѿB�Ֆs%Gꫫ�DɑDOLv�P�,�B�֋M	]����Ul�j-�-5Gn�l�b��
d�Q�E��e���e��-�C4�
DN�&���)����ɥ�v���4|�0�%\Hu��4�ꭊ��c��]�~����"�hh�j�2����b�ZFG�Z�OmvUVpdHVaGi�[[�F[���q��~4�a�	��M4�N�<&���P&iWX������UTH3��|�p�vfy�`JU|`Ѫ:$�E3�-�;�7��QH�/�b>=��Q��l�u���0�r��I=z�鴱���BȠ�>���-�F*���1u�2����^V«h�J&���2���eZ!���>�]�M�Ȼ��ǙB�C�,������K4�j��1��x�`N:!P�wUZ��\1*�v�3���*��9�zQ�Ъ�1���|i�>|����:���?bu�:��O8�8�M��o��+�y����6���,Zx��<�-~`´#N��O�'L'HH؄�t��"D�K0�4�#L'L'K'K'8�ɴ�KZmט��1�������<��z�Q~'��o1�^c�/�/��<ϑ�.x�_�0�,��Q�&2f�\���=O�Z�av���[�a��<��=�弞z�b<��'�\��&���~m��Ϙ����q���W�����I�5"L4�ӄ�mFLp���V�q���/��6^�\O'����4��N�N�mDi&�$�	�IU1?_�K�Z<����Z�<�������|}�����4�F�����n�7@ȋ��3vu/�{E+	wZT�����" �_N��O^�8�wצ�P�0�S���$S��X���0@�o�f�p�L�DP����a�7r�K���H%�Cs�9F����U�u���eQ֕�nS'�Or���
9��O��æ)��6����I.�b�LHh#����z��tgV����B*�]+Ɉ�r�.��?j�<�����0�Qh��B�I�R���1���#�SY��d�lјg����ąX^�b��ŭ�r�f#nc��yR�1+O�W��* �D�o��c��w�������޸{d0Z�%/*f�ס��R���)M�1��C�=#��;sH}��˹�����"�4֧�i��ך�i*���7{�Ã��u�K�؊�M���-�-�w2��������s,���j�>!W��n([%	!�eN�[�����FX��kLfWlA*�Y~�x��8G�7l�������� ��&�}�$��K�hh7���зj]���Ȋ�IaC"!�#H\.�'e0*��E����\H r&4�������~��7�~�'332���M����������UU������UU�����ߎ'��0���I4ҍ:pD���h_x�x<`����,���a�Et��XK�x���);(�[hi[0��5�tJ���
YV�H�c�P���͋���6�.�óiL�� �l.[H��IA��%s���⛴6���3�
;d2���-�j�^%5#�dͤڦCk�u�f���2�h��w�Q!c�.нDs���I�a$�A���ڑ��WC�Aͻ}�[$b�`@�za�s�/V��{:9���ｮ��uɜ������E?(�⡩y��K��,�ǥR�4d���'LK�d�J1D�.��~]��k�IiոuU�l������253��Zĝ�d��4\��4��s�;$���~�.��A��3�50d3�f_��m�.���FLC�r@���P��tx��jrR|T��g��6U�}���sfK�,��Oƒi�t���<l�Y�]ы���UTC�~�>����4�qx��,�}�4(�69�d���ó�+�(ɰ��|`�u��T�3CaE��Ż��q��JJ�$��Ï������C�u��x�-��A�騆Ci�cfH˔���dݻ�yh�����c������4���]��>�q%�:��I0���܍bun��-�󏟝y��t���y�:pD�Y���QSPW ��� ��QqUr�%��UQx`>�w�J90O�8-vd|n�����3G��q(�����T�)�e��Pī(B�Nqjdg�cIa���^�Dp(L\J)lJ���!�l��KH:�7�;��ee�b.;$�1��O-�6yxE0���wy�)�#�t��-�f�L��1h���$iH���ΨRD��(�y1V�4��x��V_�,�o�??8��a��i��4��'����>5J�6B��Pm_eUQ���N:�oV��՗i�n�k����=�v!�~�xن��.cx�n�[xn��8�6a��P|z.h��ˇa��\�qZ��
�.,a�r%GO��-��-�ծ�l�l֙?1U���T
�A��Er5��M�a��ɧմ����F�k�����o�]8\eKC0̔�G�)�MffX��`0l�b�ð�jl�A{��F����y����m�N��4ӆ�pD�,�����N��&�X�J�6]�����Q�J��,������-�8C5��aU��&�)"R��2p6!�O�K��JQ�2\i�'M������ @�d% @I$�~�*f~KŮ|yE���#�?AO@�.�n�y�EwW�Hג�^Z�|8�r1�~��J� 󇔅�T;*Q�>ҕ����Y��L.ߪ��5�k,�
�}'X�2dC�9+�N-b��&�eH�����kIg�ٞ"Թ��)UrҊfO���0�fgPf���2i{�wim�Y���Xÿ�ΦabE�����b�Q�a52&$����l��f����r����ww{L��sҤ��aלu���m�N��<�/0ˮ���[ڵ�^-���UQB����j�d�%E8Y���B��ǰ{x�<ѮA�T����T�9�XU�&~���֩h�ͭ�VqWK�����v�0Y���et�X�,�n_�_��j��h>��_<����ӌ_�3MQ�1���O������S�[2L�:f1�.!�3dt`Cv>y�t%5Hc�*.ٚ>�ӕ�HY�o��i�Rj���YF�u����m�A4ӆ�pD�]����TD����n(O��U��9��-M	��[j�.�3K�<�L�Y��$.��$�R0����ƾ�>>��`��x���t�સ@-VW�6U�)���~<J^	0��p�>�UUi[3}=���p%Mq�L�1L՘|}Kd�񴭴G���Կ'ŖY��т�Zl�����3K�\}wq�����ŷ��L��JRo���m�y���[iӮ��<��2뭺�P�Gcҵ)�#��x���B��G�0�UQh�,p?P��x�\B��L�����%4j�(>�F)ڲ�4յcS"bQCF,Ce͝��de(��1�'Z��93�!��smb�t��@���\I}7����(;
&�3���w4ؠ����.fL*rjb�>�78fU�*�s���-��խ�ԋ��1��AgO�~4��: ��i�J8"0x|���0� �e���ʌ�D�%�a	�b���-�J��Y	0A!�	X��-�B�J�'8m��a��.7�Ɗ��o�S��Pb�C��ĵ.wĶ�I ���f���ǋ��o���Z����B0D6Ӗ��"2��ף5�{���=�s5���w�����Т�����}��:k��(�Y�ШUN��M^Λ=������1A��(-���g��ɛ+�2J��5��2�	ǫSNg	Fw\��sÏ��Tʯ�E]jo�W&"d�Э��'ڇN`6�����6E�)	��ce&ՠ�����XRx=O+�'��qB�*bd�$%�i���: ��M8iGM<i�(�-�CJ'JUU����2Y�?.��5'A4p��}���1��!��A>��ʆ�|��6	������CP��%�O��SyfN�'D2D�.1'W���Tye�e�M�8�T.�/�6f�wM4uK-��x���{��u��N:P_иw�M7&���q�eݛ�-�s�������hoM<�q�~^ߜc�����u�<�����N'�/��?>���e�I_�^_����昴�yq�X�y�dǉ�c�����u鄔��	��Q��gIM&�$��l�<^�Cg�MS⼳���i�y�'�^�_�̯�b��y������Oby~y~y~l�2�%Oɵ���\z�yu�e#+Ԓ�Dy#����.]�-ů�/�/�o/�\��y<���O��//����<�O3s��o4�����?8����X�;��.�W��q����G^�\��ΰ���8���N�\�{H�ؕ<ٍ&�'H��d�E�V�iE$Ys�-k��:��Z�KyhO"4W�<Q�%Y��=7U�7�0����d�i3���!I�I�K�0g�خ}Ԟ�Q"ɹ��fiy⢏:W�pi��ӷ��Ln������ʞO;<z�^�s���έpj�pgG}.�S)��%
���RK��ٴiI�Z�'�뾋p�>ʶ��^R�k�D���$Y~��9\��NPmn�b��9r!(��wGَ����g������������{�����
���fff鱪������}4��a�i����i��4��'���Ɩ�U�㴕J��'�z��p��0���(�"d5�,���1{�������/Ù2G3$�t&I�Lk�s�,/{����-�c$�JHI&�N(��3��øo�K���;{�	-��,������6K���ܻ���lɣu�+>�>Η���|�Rn��%�~����/h�<���θ�ʹ��Pi��4����4hfb">�Erb���l�UU���\����.p���^�͆8.I�æ�1G�%(�>�նAl~$�p�-�E�!&�p>R�ߓ�c-WX���T�D�l�-���f���Ԉ&b�����E�g�>�N����4�P��v��Uȴ��i+����f�֫:h���f1�0X0�C_2e�N���y��|��ʹ��Q��y�^u���G��<��4�H&@A��j���20B���x��N�#��t�j�J�'�[!� ����UT&ȋ$6j,��%���e�u�.���M7�Yr�*�������+�x}.�8m1f���r��V��wg�J���1�ӛF+�K]�����`ܫ�-.���qS�8Q�e�p>��/$ȟD�0h��]J�vfN�4$��K,G�����͟<tU]Y�r�J-C�B���}���V��`ݰ�K��&G��2��a�Y�n�?>�O^��A$p5�>��D�2b�tQGOj!��%�s�'���>$0Y�e�<�ʹ��Q��y��u�OM͈ʠ���UY��`��G80�G��L������щ��b\�F��m�vd�>�Q��b̤;�tkQ5�꫐��l�p=�d+y_��
�\���O��Yut�U8hV��*�.�f����r`0b˅SÖ���;��f����`�>f��z7��ɣ�Yf&���A�O�i��&�pӇ��4t�i;���QY�k^.��v����*�i��(���6]Æ�E�[TJ[/�eש穊��;�s�-�G��,=c�fa,=_�U�t�2G ��OPf:H���4w���m�>aP���:w��]��yn����@�~�̞�f�ίƞ�ota.�i_~Jd��n��Z!�Zߟ���d�8��W+ϩ��?0�6�4��4�ǎ�"@�i�NtO	��2�6:�H�
-�q�_�I%D�h>�9>�|d���d��ܲ��CR����F��h.��Fʯ]�T��D���Eʙ��*9tw��B�A�I���������{��p�Ը;��:Y��Lb��4'R��Q>�5�7
'������Ͳb����]����]Z�gIfym�L��4��θ��D�4ӆ�4�I�d�DTMd�k$��j��H ��$���-.q��0A���6bǙ�(�4��V+m�l͕�Wـ3(B��#'��h�:I$�@^۠���nь���i�x/���/`s�b�����T����y[�-h^��J�s���n���ᖃ�w�a�"�n�<�o�̻�D>��d^��6!���z��bƑ�nd(5�8�ȟDO��L��������V�W�)g�u���n�uuVf������?A�u�cNW{V�~۩.4L��l����H<p>
4ܟB�g�Zi�N��U�A6'D���L0��D M4�����a�.B���<���H�<0���ڪ�o�Z�{��7�Q��|{iCY��t���`6z3��2sM�7M6�^j��q��!���e�B�\;�;&NC�qh��O>d�ܩ��f'�4`5��_�.Jm1�Ar"cI�I	$S�z4w��e��n��m/�&��v�ǔn�P�1�ŔdC��t�fU-���Q��"~0���$	�ӆ�<tѣ��w�k��b��������V���'L?ბ77'�����RC�E5 `�J�S��30X g�5�I@��29��Pٸj(�1��|\1�`k�#$6�M�i8�#��,��%]}��ת���>%�oI�Nx��C�T�~7��IO��ЈXng��%�)"���t���H����������?���ʹ��Q���/2��͹!�HH�*QA J}�I$�9F������~,���\�2`��MGcKl���AH$�a�Aԛ�p���V�9��)ay�~d���T�g��s&�D��Z��I���F3
�RA;�˦��s8pѴY�2�ͥ���_�E�;�$���iw9M��U��r��m0�Sts7�ŷr���#1uM?:����~��~����byzym�?>g�q�g�/�N��y:��OISi����[g�~ez~[/�����k�~\~_��?4�=r�i�>|�<��ί�u}L��ז�<�N3�W������qm����&�)�k�y����y��y�<�i}O2��b'�/�_�ɗ��c����.|��Ǘ����E�����fJ�Lܗ��4G�<�-~a~b����y<�؞^�_��/�\�v��=r���^���_��1񿭪�~:W��tf?iZi)D�Y��F���`���>)<t�/���|r��el�]S�����e|M<�'�1ǖ�y��>M���EǮT�yaxL%��(G˲��^\��2��q��/Y{�fם��.�
Go�C`Z�A끲���U �@��T�;�����C^v�����T�iih�`Q6��!��Gw�7Q�<��g��J����C����p���؝Ǖ�T	2:Q$PB7
ID��@�L,��!!�����p�FUMJ�4]��q<��_p��l�$���"�X�h�C �r=W=W����&2y�=��W�Y.�>����z��K����B�Ǚw5��|���^{��&���pT^����X�d�u���F"	�\��*J8���.b�;9�K���]��YwT�l&�`[�O7EgJ�ݘ���N���jES�A?2Gr0��"J&A��h�pX�e�V����-]����FW�0v�M��cU�-�S:����\e��ôXM��I�R��j�)q�Km�2W[h�k�0�L�#%�Q�5�F#㠫h���Y���0�cL*�@�W!r$B<)7\��_�f5�k��v��"?�3������������{��������{������]�ffo:i&�i�a�x选&�4��xQ����h�G<��l �jdAp�G1rQ�.	�3��OK�o[�r���,R�CU��Mյm�5�f5 �K" A	�bADZ7��B��VY��#Z F��,�>��"�UD�ƙ���Nqp��7�c�l��b1'�&�푼�(�D�"���L�r�QaqVcv�elX��,q��jW[���H@~�$�A�|1��4�ؼ�w0�	�:��A�$�WHDx��B��q�;|�������[-@{���\�|9ɬi�l�Y֭֭���aގC�'��D;q�p����0\1B��r���i7�ʓHB�y��4��}Ga�>y�ك ���C�E�(2d�jϯ�]�P�l�)���cɽ�?ZZͮF~�1�-j���\`Ɖ����npp�}ɳ%nc�J�gb}T�W,��Y=��iF$�"h�`�:`"@���������$f2�8J�!�p�|��p����()����hɃ#��^�٘#
OC��k�ZZ�M!��zH�yש���0�ڥ�c0��k]j���_HlVE�W���ڥ��D��2798��!Q�:<��Xux�+:��'��LB�%ÚI:v���bV|��������.�0�ͯa��E���0c@�&��ɠ���t�p�<&��	�$�p��L�:f��j;�j�[-�����=ڪ�w}Z���540ܼ-�6Ô�FX!u�խi�fs&�&'��q7�0���vL��b�x0P57�6"n�[-�^�;gM�:�f��~�qclbym�?�b���m�)hf��e��G�f����X��d���ܓ4�s���K�iT�g!��5k����,�"h�~0�<t�D���2h��%��V�)�UDv�b�������{�.���u��iV�l�9�٩އۮ�k���ƪ���Ib'L�����
��Èp�_f+���ɰ�(��9YV`:>�4ͭtz����a�**|�sE'֗yF�F馟���22h,�32L�|�9��Δv�̒��ļS��e�������u��$�~4�p�?Ks���䩥���P�ě0E�a�r5Ñ�Ӣ��\���ⰻ0R�ĞD�<.xI4�d&���1�.�d��NA8:I$�@�{�4^��(�f�5�v�F�(�S�%�;Ƀ7t�^�k.j��k�nj�n�dT�&OB�4d�D��_k炥7o�NBt9 %gƌ�}�o��ԱCB�M��%�W0 � 0}�`H��(Sm2����/�������p�)�>sK^�Qx��4`Ɯ{�n�*ִ=��Mɮ&�,s�M6{J���O��q����i5�����b��պl�?=�`�w	�P\ S��Q��ɞH�.���y����ο8㭴��H(�N'���+xAʞUTp�bQ
����_�,ƋX���>�/�W�w�b������0�nK�aa�V#\�,0`��:G�~�w$�|�7L1V����1�:'����A}��"�|r"[d�!I�@�LK\do�>��L�!����P�^��29
��jfdC���|dG������\aƖ����8�m8u�u�0x飦�Q�آ�-�d�k�	n��\�0�Ҫ�7ۥ8O��o��2~�nZf���ׂ�S^�_a�lӥ7��.$,��@�>K53�]`���]ܝ�ss(���"�=�`������ϋ������%�C2k\*�ğ�	�@���a<��֩��v>,� ��`����ԓ��k)�#����i�����L4�Ku�g��	�$�i��x�`tZjۥ�m3
��nkZ�W�Χ�v���y�V=��������P��B�W��U���)"���x�ދ�Db`�l���:��63 ࢎ�0�X�I�UUZÙ>��a��e��u�$�}^�/7y��[K���$[ioS,��>�z�ٙ��(���f|{!e�,٤�~�����J4ӆ�����=L��A�*\�^5^Jm��<Qq��$t�b���G�#�@x�D0�^My`T��H&��TQ&&\���0@a ڈ�DHRh3M<҉a`^�I$=���vV�Ź��8���p�	a�0�`U��,�]#ɲ���{�y��;Vn�����Y2�����WF�[����$����U�K,���1�5&��a�E&ʱ`�`��f!s�6d�!�V�e�ɾv˻ݣ�'i�NaӴ����h�|���>6`��5㇗�&�Ș�m�Q��Z�g�,�u�锹�t��P(~-� � i�H�Ē���Sf�&���>�կak�jC�&�+Si���+a������u��:�:��2��F%r>��̥��F��D�dYV��UQ"p3:bxK;���m��!�}g����ˣB!�P��g!��w���e���h�l�K%�da�e������j���I�f��3R�-1Ì�w���D"a�3��-��?p&9_-�j���?Uu��<۵�z2�C;�h!�#�1�_Nɚ�ϲ�0��̸����Q�`�$	e��Μ-2���y�y�y֞e���`�aB"`�,��P�ĳ�'��Â��"I��Q$�H�$�"Y�:��:�:�udt��0���A�$�D�$DJ<"'�� ��(N	æ�if�a����"&	E���0�,�0�bt�:&<t��%�:p�Bx��(��D�H
$�������6#�C�mW3ĕ�=]�3��Թ����4��P��(xT<�uk�e�L��άX�̞'�c<GU���]׹ ��]Z��e-�g���) �[*j�&=�}ɾ�A�8Y,�ܫ�nc�>��v�h3;����o��ꏈ��o]�����8BH2A�!�i�o��"�����-]�c7g��o�|����&�o��̽������W2�337wgU\�����ݝUs.�33~�M$��0��LH,����:d�A�"nUSU쪪 �5G �2T�j�<�d7��f��E���|0d,�`唭}���y6-t�c����}#�|F}?0��L$[(��>B�e���t��~0p��ft`侴�6��K>ɀ�eˇ%}k8&AL�-}<&���wuD��!�R1O�z�n�r�-�`�u�i{im�ͭ����q��0 D�4�xN��񝸘�I���C(�R��{��I��t�T7�5U�g�.pLJ%C�5�qp}��>8{���o\%]����1,^����f�}���b���W��3rۥ�O��>e�R�+$ہ�f��G�p��B�<h��&�����B�H�a��1*�a��[Kg��ſe�j�.f�&b���.�����>���2ی�,�Ř~?`�:`"@�Bi�D��AE��_���p&�,Y��DCĜ\DӶ��J�D4��I.0�U"(�Q"Ac��<��i&���F�J&�&�Ae�D1�D�C!�[7�R����i$�A}�}��D�x��r�������i#��a�2�i\��|����kK�Vb��bt�6,�猦�H"�1B��d��fK.O��ֳiMߡ�D5Y5L��+��a�=K�;O�2�k�zI�Ū��(��.��!e�8y�E�0D��W��2�2��f����F�-�r�`vj��ڜ���쉔PK�޳u�j��[���c��$F��̸Q�	��'�L0O,D�����:d�8r(����
��u�UD*Q�,�L3t��C),�0!�6Y+���}UZ�a_8�U5MR6b	���91
,.���]\Ѱ�'��l�|`���h���'��W덢��'?^(�FY���%��ҕAz��T���0a�f��[&�ҡ��&��r�*�Q0`�d�R%~�}1�T�>[�6Î8��KbJN'����و�<�$�L�)ۡ�Z��3,ˍ���%gyn׊��\瑈�ɘ0�m�d����2{�.\%2����i��M���V颂�C2XP%ù��Pv|�oQ�/��8���c����/�g�a�\�̋�r��4ZS_��m�<ˇ��www�竔�.���<�D���e�v0Y��w}�����>�S�����<%�:~(L4L0O,D��ӆ��t���H(�|\Ls�c��!�PTkj�.&���r�T�Y�[o	���Qrњd�������Z)��1e��	�8<��%�������C���%��0i�im������;in�����fwR�k&!�!C�=jr�j����&�b�=�t�>�p="Q�ᙉige3P��\��ي.(��~0�L0O��Ӈ���E@�u�A�m��`��'�� ��=*�x�~�H6 q���K�ⰺ�*��w`+��8~�����T h�с&���T�&9�p4��;�I$�LT����}f�$p}WCF��Z���|�"0�.o�ى�(�aWn{s�y��i�PIH{��4�0CP������~`�O��[&�Z�S4�3{��,�)�ܲ�~�,�쪲�ta�Z4lM�N�&	�g�Cpȇ2y5U����)ÆD�a��ˁ��A�>��Y7�U����	�|�v`�-���]ҕ��RUU���;����~�Jg݅��0N_��k�&��O�2���~~q�[i�	"%	��%�2���DG���&1���IV�Ҫ���2>�CI�:q��}(��X��a�\�â�����G	W������9<%�NghK�F���01��R���E�|�f���E,�逃M���A�+r�h!� ��iIA�n��S4[b�.��7����`��prdU��g8��fZ�O߮Uޘi�Ct�-a��������`�"P�p�y�:p"d��
̨ذ�ĒI��Uт��>���(�LD��0\�b)�5[�U�j��|x'�]^�h�N��p��:��6<�	�C?���He����Z9N[4���nS��[H:sn��몤����R�P�c��.�k�L�J���n��|��񻫺u�A҅��.��CSp�Yӧ�M����%������6v�껬�*ʲ�\qUQ�x����RO30P�>�M�*0��ʚ٪����y�媓t�֮�e�e��z}A8��C�,1'��?��4�'+Ϫc��:\(C��73
L���]`ɢ�Vya�Q�g�B���*g��8\;M�ec˩#��-%#Y�U.��7R4�+y�w'ζ�N�nN6��I�t�0D�����	GI A��$�N� ���MDJ4�D��X�H�	�,�GD�(J DDDN�0D��	D� �@�%�tDD�[GN�t��-Ӭ�a�AHH�	"H���<"'D� ��(N	âi��i��"h��0K:pK�ı,ÂaE��ĳ�JDDl��'���`�gO� K(�H<#�ĝ���5r���9��<te8�ӣ���]u�%#׭JXC�!8�eO0��D��B1*C�=8J"���m�^���ײ�K�C����q.�&��Pxt��:��Yչ&а��DdT+�*!Ot�eq�ge���l�aA�
�/2�&H ���b&�xW0�
��X��焎���z��]�F�(2i2Ck��ܶ�����Ee��҄�ih'�i�tLdjA�Cc�S��Λp����,��}���"=����s<Q�t
vP;n����s73s�3���q��ǲ�Q���rOp�{ V�As&�	�wnw�z�� �����jw�b	���a��.�ڬ"m�J.�N������L��#T��kQv��դ&Bi�i��LuKp�a<�cQD�q�q��%���Bӱn"�!ᥓj��21���S4+-첈L��(4�HM�,�ի�R�a*��3ب�5.��:l[��9�Jh�l�P%��Mf�|�5��a(1�X!G�Zh�&Gh��#��I=9�"���}ڽ�s2����ݭU������ݭU������ݭU�������M<i�4M0�K:&	"%	F�"YWS�QO	�����}��ie]M�F""J�K�����c4n/0�S��mhںf��a}�dc�{�	���uŶӱ�[b߆>5g�Lp�:��8VdH63�k9�K�*��\��@&6q���|ņ^.B٬%nũX,�aq*9%�� �Y!����3@&ζS����l3�t.#f' ���hEX��Y �06ΗR�sIc�Uu%�Q��J���AS��IFY�wIȁ"ZD,g�VQ�@Ģh��)�l��"�D��BF�9"����5DZů���,�L�q��̜>�E��2�l�f���Th��a���(�=�����{mSNLp5G�ΖQ�����-�D�p�\N�m��}�ΧA�T�."�a��^z;>6Y�œ��)���uWwu���wg���:�{
��I��T~�����DYEY��8h�a��&	"aFh�id��<��pP@�E½#��x�I �D�g��c�N�e��-��UM`�6�V�����<?P�\O�3�]���i+,n���]Ԓ{�S
h�.C��1����;CG~���c��	����%���u�9������ߤ��*�\�k�ZiF�sf����~汒˗dk@�1(,ӇN4���4�0���$L(����G�C��|*4^q�fDJ��UD2v9����+�4��h���٣�i��[2����K��bϦa�C��+5mȘ"'�n��ߜwFqa��%���S���Hmh��Q��NT93k�!�R�3�C����DFiVYf�s�q^��g�٘fj�E	�Q��_���qÔ�iȟ6�"V�y����Z|æ	���ib`�Fa�0���6(׮�O$��uA1v�<UX��0�e畊�`Q2#G�,xP�3�X�eCE�"|(���+E�$��g���D��m�����Z��)�Z%����T׿"噥��L	��h��'�rfP�.n����}�6ddd��Qݧ��"j��撚1R��b�Z9K0�5�_�Z?*:F+u�f˓�߭w���p��tD�&X�"Q�p�L4и>��R] ��a �F��E�u	PJ�*!��
d:	2`�"���5%|x0J$�j7X���*3D�L5X+\��~��oYg�ф~CZG�1�I-q`��oHU�h�U�|Y���]���d"����5��r�u��fO���,L�!�f=�����saBz�:3�KG��=�^1��!��V���2EQ=%'�����r��/�&�q��o'�f!�A.x��W� �=���C�P��P�ZI�Ώ�~,+*��dh��j�!���\f-��W�x��m���e�G+R$b�}K�ܘ���e�δ��:�ϝq�Xq�q�|�IR7r��]T�}ڪ�F
�|Ŕvxab&��(/*�B�O���g!�0���C��a�c2�>a�9�xQ��4\�<7��������5x�7��gD0u����(�'؃e���	h�Y�O�F�,H*7A��<�*�}K9kDr�b������go�8�#�u����q���1�W�j�ü03�EIJ�-�|�q�Ϳ4��θ��\u��p�������L�P��F^�V"jQ�e�Q�g��p��v��z�#l-�j��rט��Ô����n�S$F��Ẉ��R)����SE�EC�|\��M�K(��B�07"K(M�ň�S(�hqf�M��^`��!�ؗ*���$ș7�T��̘mk��s�_�����y�Zy���&X�"Q�p�L4�.�F�rn"��@���>�m�D�(�SX��~&hvX�e�~��0Q�!�  ���OJ4Ieq&R�b��
P4;I�v�pD�����!�`r9%�(D-�V�����{�[0tq�P�B%��"�Ǔ]]n��-�FX0�WXZ'H��MUb&DN���!�3��<h��gM4�&X�"Q�p�L4�}�9�hP�]tNb�*Y1`b(C��$����
����q�3a��bhLI"�-��#$M��	�4�	��@��>�I< �l}w^�*��������9XPe�g^ǐ���%���r���G���-��vos�4/A(2e9OR#��m��u���s��v����+���#V�-�Ye�%q�\?[O��+�NDk�a�G0ȉ�L��0d��;e��ШPf�0���l3sDD�T�,�7%""v^����7t����z�]��ɣΓ:�&:�ϟ��ր#�R�%��'�	M}˂�K(D�J�_��ژ������r��|�o6���<醖&�aF0�/�"L*�fj�m�-f�9K=�U��(��B�3m�	�Q���a�b(�z�%Cy2\<bL�^4�U���6&�t�0�N�ٟ�m2���bPfXk�Ϊ��}�&���r��a�9
�`����U�)�q�KLCɏ�x�(��N���P�ħi�u�C/�'�T�Dd�][Z6dݨk��Ӑș��B�)�%�ԁ4���g��0K0L/�:!�:'���8I'��$N"pD𞨄�0L<'�D�&�p�Ɯ,K<'�"A���%�	$�!(�D� D����"%��:t����Ӭ�e�F:"@�@� IDDD�"pN �$�pN	Ӣ&�i�h����tK:P�&	��bY���g��?$"'��tL,��<@�$�'�I	�X�=����zo2��g}�k����������t��s��k�ħM�����3ק�Fh��sFw&����6�0�G:�g
�o��>Lg�t���pw�x�lä/ us��ݶ�&t�}۶�r�|a�:�a�5���0j��wp�I�.�^
adZO{CË!��ɞ�a�I���7>�{}�hP'��D��A4��+��-!�`�^���7}9�6����}'�b�z�+6}�J��^fe������U�̽��ỻ����̷37wwy��f^�f��O4��&���&�aF0�,}� �&b2����¦!˵Ʒ�窩P舆��`�A��2~o8�u��z��x�,N��^D�"W�m����m �e�g;�����H`#��{E\(�diy��d�Ɋ��'&lɩ�-�/��B5FJ$,�+%��1
0&�jT;�A0fwԕ����BhJ��.σ{Nl�ǌ��h�ib`�Fa�4|4Qt���QB��e4��$�*#��<����ES��SK[H������ϗNA��uK�%��V�u��:w�4-�Z6���6�#Bd�}NqY�m<�'���ͫE�Q��i�SE��!�9:�g��֌pKI�5p��`�*b'gao��I�s�iuo0ұV�0��ŝ4M,L(8af�Y܃�$��蠢�ALx�����YB����`�ԗ%���A@�����ͪvaTm�J; Pf��WĒO#՛�Ƶ���%u�����h�����CڋUR��1Sf�z0��Б� �s�(�׏�<'�����2olZ2%���8\�͖�G�#��ob\(����M	�vJ8h��e����`�;;���p2}�&��vIb'J<Y�p��V��51��~ABԉ���#Q>�����OէP�3�1�y��N����6�<~?	��%��aF0�M,���r��,�@�	F�dB���UX��N]V�Z2p�"<"�����hL�8cK=Jɍ�2�25Xy�I�H�|�u�I)}�Vm�Y7	0��j(�dMN&�+�Ÿj�
H�.�҄�b`xw�p.A,Mt����3'J�U7h�Ð�Â`N��l��\f0|I�N��0񦉆�%��aF0�Ǎ����eWv��g#�P�ag��F��=]a����ڥ9�m�rF2^�
2!���7�Bw���>f�JHI2�A��+��p~�;u�_z�-*S�	>�>ih�I0���ȟdу�E
"k���Ȗ ��*1;�j�kw���	�k��.ҭ�C�t�g?%,O	���0�ı���<x��=�E��UX�p�GM��˒��>�g��Bx˅��g���h��O�V�����O�]Ybl��g���ᛏ�����0�?�dO@�c���nҮ�&�J;1c:��0dM¨�r{3�5��
�P�_�~���dL�74���߉(���~,K��,჆�68+n�w��z�͘r����%�L@�x���g+�$[Эh����b�f@�V`�6�1i��Mz�%��j�&�F�Q��d�bzI$����M�����`Z�jD�n.B�k�X7��I��@�zv�2�Cz��Ɣ�{؞N��_�y3PUPY��L 4���;{���¸��bn;Z<\7eqhЙ7�x[��(3�4l�dM�eR�i�z��9H�n��i���U��6QG�,�5���^*�p��22c+�V�(#ӕw��R��X�6���ġ���g�*ǥP�R.��Ӈ<Y����0�ı��6x�,Z�U()m���D�~�t�<��L2�t��V���y��nr��Gйp�)��(��?i0�5R�b�6e�&�D7N��,�����N�����>1���r��3F�x��UQlŌ|')x}*PY�Q�a)�˧#H��=Ky���q�D�����%?>�+�m��ߞm��0�ı��Y��{�D&*�e�&*��UX��P�C��=L6Z�G�]-��/�a�z�f��)��}d�2%����`PFA�	l4�g�!QƝ���0V�eZ/rnJ��6n<�*������
��ɩ�a��o�A*rz|��t�^�d6&D�l޳��]^+�pȘ�>`�s�w�J<if�D�K�J�8p������.֒�����Ҫ�MCT�ٜM7��l�W"H�oj��O܃��^��ĳF�`�EHs��ꮪ��EUxM=������o���3	Z���t�p�A�39��1mjvd6���R�X�	��j����CF0d�E�s�K1%&A>�����IM��#�E��)�^�gM-&0�x�K,�`�&	�	��t� N�B'C��8I'��$N"=�O�N	�
��,N�4�0�<t�4<I�"""`�4E �pI�xO�bt� I �N�a�,�2�:u�GN���D�:&	BQ"@�E��;ȄO	��i��i��'�:H�&	��bYY�Ibt��x�"$��,O	�Έ�Y�:\���I҄$� D�9�;R1��֑zB�Sd���B�u3�F&L�(�4Lf�3y!I��dTUQ$Bn��"A�,4,�W,a���n�˅6��!�B��손G��2nn֡�T8R��`I�'w8�̓�Ck�w�aYG�Ut�`�T���ܤ�ε)(���9,�J����׀�P�7�K
a��p���Z�(n� �S9���K(�Ͱ�Ẽ��Ȃ,󫽂�d2k�-za��k_G����z��;���x�KB]�>��Qú�w��S/w�-;�͕�}v"{�T�0^L"!�U,�3g�lR�Y�9�=�h�Q�d·L@QB ԅ�� ��c�MY:�A���T<��R��k8�/����X�JD� �0Sl%E�	�͌jb�f�V1kG^$&B�1�!\T�&��f����l8�+[n�Z)<>� �+��(��N#��6ZF��p��V�1/77�7i��r������:�ř
��j�z�@�24D0��L�"P��T�`!%UB6J���0�Q �����l��������w~�w��wwy�ww�wwww�ww{w����ջ��m���N�4�<i�a��b%	F0�M,�/�f�hj�-��1�t΀�`,��S[
K-�h���r�-��ؤ��v�L�`RZ޴Yl�2����]�z\]��3F֨*�2�b.�ìn䄶�f�̶����h�x�.Geg�hZޞk�tԩx�aw�Z�4n%��[-V�ԙqW6:��׵-l��sv��0�E`�j`��B���+X��$�xA�x|B���n4!$o��¹���T)���,�P��i�;�R�:s�\�՚�3ʃ�l��>;6^�gKT�K
*���Y�7�6a�RJO�Cݩ�jhM��+��i�sK�6��u"尶0t�Ț���3��ǎ�Bf���i�I�I���c��^�>0(!cI�q	1"\�@��������fgD�C\�cU�w�]�E���,�O�	���L4�,D�,჆�6^w1T5���	�U&A	")�1� A+���i��I��4i��5]�������K�����U��C��1=	3���mr`M	�b4Tu��˅���&|���R�p�I�2p�50T�������)K�!�6YH������.C|z<ˌ2��.�>'��G;kPɠ���M0}�}���{�-r&Oi~�ڣ5��M_OW�7L��l�y��ߟ�u��>u�a�\|�ϙ2�rf��wh��nH�D���G��CFp�dKb�[�2��5ɘ�|�|��h'!&��FY��C��	�6�Na�e��I	#���$4RH�~�`��E	�������[�מ�e�l=�4�"5O��2�V�r��+]�4�Y��LS2xʹlȝ��O��ؓ�+�6�ۏ�<��κ��"P�a�4���{&&&�>(��i��Ub%Cft�읱���3�۰�����Ϲ^|���X����-�Ӌ�"�!E&MC��#T�?nL	�b�}
�`L1��R��2x�bQ̢R�U�,��Ԅ�>���4`D'&N���f����	�6&�O�qu8YX� ���a���K4��c�������H�jʐ!��Hl�c0B�iWSfc
5-Y~�4>)��L�4��f\Թ��ȓ7`���!C�$�xA�(w Ҵ�Xe��		��i��О��O\�v���� ܻ ��U��v���	��l�=�C�]B����+в�%�DWE�諸�8h���ݪ�QpMΝ=��^n�X-y�D�5��C�F�ܘ�3�vn�A,LC����\���<���n���v�إP��97�=��۬�N>e�]/��N=�L�1�Ζp�i�4D��,D�(��i��z�虚�����UR��V"7��v���G��J(jҳ����<2-���ҫ���0o峢sF
���4`D�jR�q#�e�>>��_䑶��'0"tb0��͐l4�A"�N&	x������ɼ�qh��C	ګ�e'�q7O�Z#h�?����D#FYo�����o���>m�ߝm��&�ib%	Ft�M,��f~����KJH���-XlĢ��J�1:r�JU]�/���Ҹ�xtM���:n{�6%I������1�>�Bh�/L*��"v�M�C��E��	B&�e����s�6��1��6wFD艖n��CR��i�j����>�4��|ɔq\�4��$��N	�
D=�?�M�	y�Z%?[��s	�~u��[qǄ�"if�h�%a��4��z(&�-���$�K���V"rM�:��UT`�nc%�����̜��İPC3K�[("�(���\,��%�%Ý1�(���
��-�9�e	�ϡrT.(�<n͕T�Z�j�Ŗ&L�W0�!�2�̉���e�)��7��ʙ�ͣ*~m����$�n�Gi��^���N8���~"if�h�%a��4����Ƣ9��0�E"�xP�������c��<��l�o��K�*�l*�-@]/�bh���f��0�74��.�6���1� l���5���_I< ���{�yu��1���@QO�$�̝�t�?
5L��H���T淛��//S�D��U�g���-+˪�4�Q��l���j�9B}�*�F�r"b}Oъ���G�j�#TӔ�M��,Й�%C��|�i�Qv%k�5�qXqI��&sG���2%��r���/~(�4�<i�&�if�GK8pɳ������J��ܪ�DCAe�QŖ&�8h�8��Jn��8zI�d8#�i��7�aj�b`ؙ�'���yp��"`.�z��`5b�M�����;߾���A+	�V���L�C�duK:!�5ȕ�,���*Y����Tݚk�]TѸb8L����	���L�V�E���N��ߜ|���\u�`�`�YGD��D�'�e8Q%�"H�(DN��Ď�`�B'D�D�0KǄ��X�:Ib~ �y��i���I~HN�"'D��b%�(�Ӯ��GN�dɖQ2A���$��"""x�$J AH(J:@��4�D�D�M4�0��&	���,N	�'<'��"@��:"Z4�>m�m��]De�KGN��#��=�v1�g.>�Gם���p��^�<�˹"8)"OvX�b���7���?x.N���|J���2F���ժz�^3��ѳ�}�|ޙ�_��L`>��D�G�h�dY�w�}Ǒ�v6j{�O�3�l�����\�ni����o{�ww~m�����ww~������ww������www�����4��4񦈛y��:ì8�N:��nI$���+	�yzxѝ�j�X��gJ,MO$�/)��A�1�t�Bf��vVI��N3#|
�da�ɮ�avl����,� :x�P���U�mD�8��ϖ�,����h�>�R�����s'
2&�>�WՏf]��r��5�#���{��i<xӧ�M,��4�P�a��>{*�ĸ�j"��IX���`��2>с�mw�u��fB�	�ЬQGU�Qk&ګ��h����*�=�ndD�3�'��̚��UUN��C�&�̊�G��lɳ��>򢍗0hD�M�̙$�15=��c�v��WrK�Ju�Dq���k|�֟>q�Vh�f�x�(J0æ	��LE�9*q#,��E% �P�4��'������R�T��pWKѐ�r�V�����1Ts0����O8��u5�[�2�����A�I'�E�?u�;��$�S�����N�a��f�ǒ���YF�6�X�μ����p٪�^��8�!�\��_\2pNJ59>�,�,�,�5Ӆ���[ف1#Q�Q^'��քUvpK����_5��q�xM%�]mrp�k�"rJ:&`�7�ST�>�b3
��l�mȗ��WUO��޸�����+fmH��FJY*�ܜ`�X���{�r�$}�r�a��|��|�믞y�D�(��&�V��p�rb{\��|O��)�"޴k\UX���a���Q�2��F9�+x6SY�e��Ey*l���vtON��S�4lM�b��χea�7u��:=7*n_3��( ��tG���N�D ��Srx�/I�h�3Pl`ˆ!f�G3e�0%��o4��&����N���'�K(�a�M0K4D�O6�:Î4㭼Υo,^.�R�%��U���(�s���<}�͞�s��L�E��c�e��18Q���dȗ��O��ڦ�ҭ������0
���vYFä��P�(��T�%}wĕ��au�SV��B}<;�k�T��2dMڪ&a��C���|d�;��!�t�Gn#�a�Y�af�x�(J0æ	��B'�����8��DD���Ub0y��oBɳFD����Y�B�0u�I$G�A�@�@�0�YJ��Ȏq��Y��'����,�I
@�B��dȘ����&�ߘ�0&��zcEz��(N���/���l���U�=L��|�6�O.IW~�Fi����y�Tۨ�;L>wL6��l?b����Q��m��Y�af�x�J�0�xӼ͖��ňAj��H�ؑ5���Bņ�H�0#M�Yj�Hi�%P���k*;��ܗ��ò舉< ��I'��Աk�oͷ��t3 �Dt#�~GDe{�^>'ؼϭ��\�z�au�`}�O��3��]�/V���dØ���Y9+��K)�,f���P�����E7�Ҳ�����.{NZU7V]`�g�%I��Ħ����!P�͛��%n5>͛�y�ʷ\`�}z�$g9[����g!�%��!�c��R~��+)����/�4��Ϟ4�ƚP�a�LƏrI!���G�6�|e��DpA4�I�,8���34mu�kA٘��\��(�C��f�097��1&I�^�;����{2�կ�fx��C�����N'!5���$,�C��&�>���e����p�
�A>89�aP�,�R�6l�x)6 ��:X�x�4��Y��4҄�8t��8�4��J�aO�����Ҩ�Y�PA� Ϗ9��
��2�j�VN:�2��Ѧ��1�K7�E��(̳p���s�}��%d�����I0Lc�A��ph��\C�T;�AT�f�hȋ��fD�<Yߢ+�b`ؔcb��==��\B�a�T�a�pɃ:9OG�x���(�Ή��&�h�Y��<���8�o%Q�R;7B�a��M�1'�1�k�=m�Z?H�K 2�Yq���3P�A'��ܟM�ʯOSvn"j	�΢��;S�7�ك�gIf��,��w'j��v�Y��y��ӫ-]��ww�j��ynS�8�|����4$���'��H�0_�V(*��!"D�������F����J��t}(ɒ��a��$�I�Ɖt��p1p��.^ �"�b�!�4bJB*�	HD%AT�"HB�����Y!J��JR�JT��J)aJR�JRX�JT�����)aJ)aJ�K�BQBR���T%�IaJR�K
X�JXR�,)R��JR�*R�BQ�J!
�B*��JX��J��R�)BUB �P�JB�	HB��� ��UC��BR	U�BR��BUA���T%T��� �B��R�JB ��HB	HB�B�������A`� �DD`�!#F"D`�H�DF"D`"Ȉ$" �DF"#""0�$�F2�2"1FD�Ȉ"H�#dD�ȐAA�##dH$D" ���dDdH ��$FDA"A"0H$ ���$F�F	`��F�2"# �#""2""ȉ�# �"DdFDDH�dH2Ȉ#"�D�"@`�#F"�"$"�`#"#"Ab$F�Ȉ�DF	F#"0DDE"	"1E$#"0A����H1#""$D�D@DFD����F�"Ȉ��"AF"2"DdD`�ȈȈ��A�2"#" ���A�A�"1"�H0������FAFA"2"#"""2"#D�"2"��$#""0DFDD`��"��D���D"R)���"1H0F2"�Ȉ#" �(�0D��FDA�`#"0D�#�Ȉ#F�"0H �A���#A �#"2"D`�#`"$����ȉ���A�	�����FDA�"$FDA���� �#H��"R �H�*%�`"D`���A`�DA"ȉdD�ȌA"ȐH�D��F#"Ă"#"$FDa"2$H������# ������#������"2"#`#"0D�� �0F ����"2"	2"DdF$F�P��F���"I,Q*��#aURT)RE�IU$�I*���I	�BDF$�JH�QTJ�����%��% �IHD�f��-i|�0����� ��B�	HD%T"	H-�"B!)�BR	H}�BR	P����JJ\UZ�JA*��d�@�A�A����EJ\R�%!J�!A	HA�1)BUB��!)BRL)!PA"A"A�%B�ZP�%����BUB!)^0\-��B�B��BR	U�1"�"�"�D*Q�BR	UBR"�`� �D"�"�DA�A��D%!��EBT%�BUB�P�%�BRA��"�K�(�B �"A"�$BT**��JCV,��,��,RU,�Ɉ`�R�B!(�A(�̪i)�J!J�D%!JBT*RP��B"	HD)�"DA��b"	HD%BT"�"BRP��!J�EBQ	JT��QK%*R���*���B	UBQB�!�%!D"����**��	U��!	U�@�"	`�AA�3���!�"��EBR�D%T!	HB���%!
��!�P�!	HB�
�PB��B��PB)�JB�JA�P�T�"�Y)b�J*�)*�)J%TBRJB �	!)
�% �%T*B��B	HBB�!(����!��*TA)BR	U	HB)BR�UB�@��A)�R��B�!�B!*�JB JB�JR�,��K
,��%A	P�D�%AJ��"��T%!	D!	HJ!J!P��(�����)K%,��E	Y�J�`�D �2%)b�JJR�)K�P�DDB1`� �AdA��"�!*�)BB��)�A�� �"	dA��dAdAD �IK%%JX�JY)R�JT��,����*R�JRJT�E*R�%JY)JY�R��R�,)IPJ�!!	P�%!���%T"�	UBR�J�!)��%!)	H%B� �%B*�JB����A"����J�D%!������R��J��K"��%T))�"��%!T�B��A���D3t�!*��J�!*�J�B��B��%B�@��JB��!*�)��b�B1B��BUB J�BR	HJ�BRT"�	P�%!%B!*	P�PJB J��%BJB ��!IHD%!*��
��!)�BT"�(AbD ȃA"A�=Hy��r�4v1�-�5��0�f�7*vJI� Z�H���tb1����ٶ�Sm�\=�7do�}h�}:٘x9�M��l~��h��|pn>�~���4�	�0ܮnZC	.�c���4��a���,��2�3��2t��lm�����������0��w�7��0�$O���'�o���$�l��~�8I=%�H�?9&��K0O�{�w'�s|��:��}�'�0��)?�G號�Rt�G��eh�9+҈�7>�D���?g���UM���I�w�G=�hO��7��c)c�6G���}��gPb`���]͡�u;�펨i���ٔ�Fu��������=]�#9�I$�F0αr�aL�De2��":��2��3���(�edX�S?4_��Z�d4~[�K�u�?�y�:3&�Ǆ3�ױҚ'��1
nb`�ZU$�J��iT���$��$��RHI.No���wa*pF�6�;^D���R�$ݹ�Nrp�F�N��3%0����퐳�������(�"D���L�2��I�j���i�I�w��(��C�t����F6zϣ�yZ���>�S�F��E��r+�9�'�s1���:<����W�<��'8y,�Iw��|�R�'C�������>%'v�bG$��H$�U���"}gj|",���:�iQ�\������29&�N�N�M��(�5��Rr��ij[Z�	�ۉ�4�:��-�BH����P��:�)@�a)�lf�%�a,(�0���DƲ#Hn�byA%��0XOܗ�L�C�Hp��t�$H��ԛ��~��;���g$���"z���"|$��:�2O��Hw���&�:jd9��uEFB8$u��|��v�]�����)&<#(�+	�O���N�"D�Ɉ8�:}h�RO����"n'kC����~����jO1�:Oq��G���i��Vh�m�nH�OV��1K3�\�0�ix��da�S/T3��'��OW�dS#{2t��=-c^�f�4&i��ƭa$J��擒N:��EŎ�꜉�?ل�3:S�I�6'����m66��u-a�Vd�#�zӃ�|��'O�`���%��O`�sF���/�rn���z"�:�8`�g<�lI��]n�	��7o�A�},O$[+�(���P��ޟ�rE8P�&�