BZh91AY&SY�.6���_�@q���"� ����bD��       ��R�l��-�M�e$��[-���@[�m���MV�����UT��
$
��)"�2V�bl�\�������C�[6�
���4lm�MZ�ٌ�U������ZK	IA�fśe2�l�i�lidԅ��k6�ڵf�U-��յ=����϶��6-����n⭔�Jk�wNkf�ȩ2���[2�Km3����6���l�ef5RZ[E*Uj�)F�CF�2R�����j٘�g`qɰ�Kf�l �   �}� ���huB�k��Zt������WN��고�\ĵT����֭�����f��
Q���L��&T�Y+x  ۼP +hm��(3����(��� ����ЧN9� k�Yv��9�(4-������{�JR���x==:R�����(6֫i�ѕ68  �z�
R�N��T�K{ǯM )��p:��� iJU..������u^�@*������J� ]yp (Yǻ�P�kVɦl�i��m�,�� k��B�m���:�i@WwZ��mkz��=��J�oh�*���{��� =��T駻���G��pB������CM����[fm��R�Y�g� ��i�

C��Ӧ�q�t�U:�ƨtI�]�
�r�T�
b��Z���: ��p�������M\,�4�H�f�a[ex  O=
�SR�*��c�,�
��g0 :c�Еm����Ҩ*k	��@eT�t ��)T)���t��)�vʙ��XB�f͡Tm���  ��( i��n�U(.)�t�m��0n�$)��7P��@�F� ���A��)E ��8Pѡ�w hf�e���Vkwn�H��M��   ;ƀ�=�h�(�  ;�� ;8�
�v�� Sw��C��� 
��8��4�Sm2مfd�-��   ��  .N� -Nܠ
�g 
	�`h���@ ���;I� �-�Ms��h ���km�Ef��V��-5f��  9����P�;e�EZ��ࠠ6��� ��v�p �n�:����@��@O�    }   ��2�*�0  M0 j��b���z��	�� �M0�����)*��L� �@ ���J��      "oSS
�zLj!�0&�04�ڔHjaLLji�OP4ځ��H������:6:����t��(\��[d��m�T�qN=�|R귔9	�)�|>��}��
 *��*~� ��БQ_��G�����>��qS�h����j����U��|	S�Ң�+����A��G29�0̎`s���3)���fS2���as)��L�S0��̎d�fS2���̦`s�09���es3!����	�\�f�2���a3)��f0��&e3)�L��S2��̹���&e3)�L�fS2���&c2	�L�f2��̦as&af0��̦e3#��fs!09�̦a3)�L�f0�Y�̦e3	�L�fS2���L&e3�L�f2��̦bd3�L��G0����f0��̆d3!��f0��`̆a3!��f2��̦d3	�s3)���0���&a3!��s	��f2�̆a3!��!���T	�G0 �A�#�s�Q	�@̀&e̊��2��E£�T̪
�eQ�
�� ̨9�0�A�#�A�� �aÛ9�G0 �D�#�Ps(�e0�0(�E£�s �`���0(��3�d̢9�0��@�#�s"eA�""� ̈9�2��2���W0 ��sd3 �`�
����e0�̂&d3"�dĘ��P�(���0
� 2��� ȫ�3*�
�d 3 �aU̢dA3!�Qs9�Y�S0���e3)�\�͙C2`s	�L�!�L�f�L��0���&a3	�L�f30��&a3	��f0��̹��̎ds	�L�f0��̄��29��ds�L��L�f2��̦a3	�L�0�C29�̎ds#���	��`s��1��ui���?���;1�����z��S�vӴ����r�h[�n���m"E�dKsN�[�ɻ���-��D��	H�.�r�����4���{��ۛ4ٸ¬ǫ���O^�ܱ�*�F?��^�f���Ť���h˶�d�F2����P��5,��EZ��,���WyP2�����\ٞnen"���ƥJR�cE��2�V׎ڵ��+Ew���f�F�ʗ1@��f�S������q[�]±�{F8�b��r����A���+|<ŋ
�návsYf�l�bS��l�m7N�GM+�z��d�#\9Hѽn�ᲊ�D��hT�Ӳ���[�1iw�ɯ6�f&��I�(K�`t�YT!���$�;f��M�J��933֘����&�9����2�3���y[������em;�#���!Kvv�̪��xUX�X�!�7Vc�]I�n��@9-UҊ�h�͛�`�٪�V\@/(�wn�V+�%��v:�l�f���U�#��Ȳ���B��:���(7c[X5��̭q谩&�`!��u�L��^�E��tv�m��ʕx�u��7swݽ��l��"�ͻ�� ����@�-"�Z%[=�B�Uˍ��n���;ǡ�k�kջ�
;�����H�;n^ɚ�d���)m��5G��{�]ͺ�kpje[X��Ӊېf
Wۦ��,"Fb�O��?<r#�V!�*9��8�(n]�4��)VL����[ɗ{��77�^��M|����!y۫1=N��t�����FX��1�+HA�j���a鷺�,�Abʓ^��Yh��z͆խ�����P�S�k*e�
7���3�x��5قZ��T)�����M6KY��[�׳_��d�f���e���^���I`f����P!6h��B.7�5�e4i�	O���B�$]�Ǵ�#j���1n�k0fb�9��];C6����A)Vއ�+f���[�2�Q�<���^�6�Պ���&[j�4-�n��2��Y�X"�ܘt�29"Q�P��k����7KR�ڽ7m�6Iy�@X
��Ø��r�c
�J�s�*֤[oU���[=x��6M�a�J��Q w[�Zq+Kd���B��o��7�J4�S�jٰ/,�"�sf�i� (t��q��J�Je�5^���������En)+��H�9{
j��n�"��E��E q�5P�D{j^Z ��tFܵ7^�.�VU�l�	��U6�8�7�M�R��Ք3^ZM�6i�_��/H{Z�4M�٧��SF�^�Ɋ\�Q��`=;��F+������j��j����h�F�]��N��/I/U�L<ˈe:�QH��nP�B�Z���~�ȷnf�Z���Ŷ�Ҡ�e��W&c�bmJ���y��D6�B�S1gr�b_�Ų�,(�if�QXܗ0lM]���n��!��80[�4p�^�wZ�>F㭹�Z]�cou���=�A7���睡�yl-HS�������9�.��@���5�f��,��61�XcYX���F����֊���]�=݂\0ye�K��K����R��X��Ԛ�D5�R#����-צ�	VS����0�Ku�N�fZ8�����z4��q���/h�w67�:�A���A�ӫ�U;x5���5��Nu�ò�Mm=�#H�!UUQA�5��8鋨�dAԮj��sQ�v���t��n��F�^�e %V�����/CE��a��T��%uT2��x��5�ᕍB����H#h�PSN�x�'oq��!���-+�Ɵ��x����w���Gi6̈́V��B���uK2�$�:�P�xd
��e���t�s.n��"�*�ɘF+0<ʷ$�˻�Z��Fh�A�����qޠ��L���!.�ZFJ��3A��v���B�����5[�ڔ��N
�5��/Q'���zQU�)L�+/s@���-�I�	@�A��Pf���Ɠ4JɴUl�-��C@�f��f�J�����!�4��e�Bp�&V7JKt�^���auakf^[�os[A�L-u��e�Q��/�,�]Ve���.�[�RX]��;���0<���vPU��N��6�5�XZ��fi,l����ZK7.��b�R�V�@*:bSS��	u�F�sFҘܻ�0u���!�;�t���@`�qC��V�E)BBF�02v�Y��T�.�G��s3`{��g4�I0�o|�'�haٮ��E��=:nd�W�PɄKr�ʺXh�립���OT-��/N+[�0`�.�MR��\�U7x������o蠽4���9�R�0��"�5j�1�b���R�
��\����X�ݦ��kA��Ĵޗ7hj��QqiQ� ݂^���ǵ8 ڱ��2X�y��fX���4�&6�GgX{[Έh�엵�,���ܒ�;@CbI��dB$��9��R�i�ܖ�� �[Wh�����缕��yy��v�+g�m��h{/۷�[���0-m+Ȱ���ɀ�e��kbm��%�񭣮,;���&�n�FYѦ/sdX��	�)����(�~̙B�6a���u�Q7�˳�c�hhZm�*A�.��Lܙb��Gv�ռ8�%r���Qݙ����k�bZ�01�i����O�\�����1��[w��ddB»:u7���!\��r+�kAN�̽0�F��L�4��l�E���M�q �@��TjQ��A�n��XI�c(V��*f
�]�̦��H�f�n�a�0����Zm����A m ������e�:~Y�{q�7y���fM؊�/,��@�7�T�ݢ�!j��Yh�s��n�	v�+YF��$���z�@i���>�4�u���=�jv������A6��� �ՙ�9sF+w$Ĳ�=H�(EтKYx�`q�v�{i
VV��122�e����!,�f��(��w�(,����[�N+Ic ᦵ��`�6��Y�
텛���Xgt��e�î�캗�bT��e�d�+U���ԍM&ވ�3����ѳc3ܵq�u��FIӷ�jD�)�n47n��L��A��(e%�#O^���b+.+z^��D�
��ٚ�x��$��l+wD������'E���9��;�En��-Ջy�Y�y-���;��3g���%�rm��7Fe	�T��:o%BK�`�d��%�	����z�����ѫ�*����e�"��.�Z�-�m��8e�Ę��&{2��/p8�M�qF�i�2�ɑ�NJ�Qa���3VjئĬ����OY�k�Am�8jn[0l�����R�+r�6��Q10K,<��PaZ���8N���$xp�;/)!�yk�NTvv�0E�ɂ�p vlj����&<4� &�w���J�E�H�<�gk7�3˯u���U��{
[ �o;Q�����Y��ژK��u�`n(��A0c R����1h@��Q�'3,f�`+P1h8�)���aF�r�!#ˣQ'����@�t��^�lS^�����m&%�㶫K�����m���;�����E��U^Q��(���M�a0h^� �iT��`�R輛�ejh])�e�c[t��^ZKX%F�f�8���Co#i��Yû���m��e�
k#��4cm�a"���ǆr���;�U� �
l<��d&dqG���h8f�J�n1�ER���Q�j�5����Y�6C(h%n{d����K�����ig^q�M
Er�v^}Mڿ!�����-n�r�5�\a�{fh3+,�h	�~DJW2Xd�a��R`�WLf!��.��*B��,���fŀ�)d�(��b��*��n9��RM������+v�T�^�H0\��xF4NL�r�jQW�B�:�e�
ɺҶ(ZR��L[6M&��ڡB�y"�ѣ@�aE�e�2�[�����U�1��壂1�,@���V�f�Kv�`Yy�-���3r�Ū(�%��^��6VJYBK���Zqb�����Ѯ���>�'��:����t᫫�
�y��fb�ⓙu{I��%�����Jղ$_^���Z݅��[՝�KI�����ԕ�wI2*��n�h�e-sܔ^�:ʹ�^���v$�ݺuR�g[eSՆ��I��ee��#�o%*0U�*�k����!��(��t.o�u���U;b�͑j,ʽ���łJך���l�j��ʥ�q�n�4��;A�ذIm�nM����8^���u�q况`�X�\*��V5�aY�u��eT�ط2�jSSh@٢¥��(:�E�Zm���26��r��a�Ƿ	q�bS,���a�HM���2*=T4�p�5ͣv�s2M��`Y�zH�Њ�K
9���{�/*^(�7w��tM�,ێ�	�{Yp\ �ˇ,���(���v�o-�$YO���Xj�PA����Ckj�jh�'��a���GP���!���a��H�ݳR�8�Vf�=��sp�*:��-��5� ��kZ�:w	��!�oAx� ����3i���뭳]D9�N���T��Q^�-hR��Z���ڶ*�ܭR����ӧ�w��ۺ-b�f�I5"j��I��s}�D5�4�m��t��	 �m�s-)괫AŎ<Ƿkb�=����8������6�Zr���t�cCX�	�V٦�ɚ�wa�JPųZ%��,f�Ɠ�i����+������_�Ⰺو�7Dy2�Vӡ��Ӷ�n�C�h7�6�n��/ҕ3�0��Cr1�(�`�졌��Ԡ-�2��ݬ8�d��iԉk&�tLQ������ڊP�����̭�l��z%2�i�f
���U�K5Z�hZNc��Vc@Ƚtٺ� ���,�l�f^d^~ùu(�5("a�(�gU�L��4f�t��z�a�]*4��r�
{��m�&:
[B�"։���0����ӌ�'DY�r �&�Ԣ1�a3㶌��K���4�F�k0V�E[�R�m�ю1S]創Z.�c[N4�d�$�v��cX���r�eû�u�ڶ��"Y�M�lb	q�َ��Լ(1���}�z�E�7�H�*�Ռ��gڝ�R�@��㹦QgM"Z�A�O��m�C[��c5mǊ��7(䗬�Xc[3�=��YǬ���t',��H��Ef]!��2n*����9{�.X@�a�U$y�5�B���$�,���f��f��k����+q���kP7eM#uxn�m�OcC�D��D�6�&$7r�֫:C�kv<؉�,��JV�72
�M�g/D�u�`-h�������-�3$KpC�z����PbB��+¶�����Sw3CH���Ê�]9SeZ����=����0�0V�ݽ]���ـ"�!t�]��ѡiюX��!�����1�N+t#vk0X�rD�د^�7�kd*��}���j�ȄŅ�JB�#.�@�؇4�Ok$z�i9�լ{pܖ7�LZ��E8U=Tv	Gl�����{�y��YJ�B���D���yY,bZL2��)�:��3
�Db�*н10X�
lT/�e����̡��(Ô���b�jd�w���n+�H�FM��ՓY���m*���b���ͼӲ��D�ާwnM���ې���V�v�NZ�7i��ku�����g+6�����l�\�m�јH�|u#ֵk��l�mUiVW)B�o֑���{>F�`�6���W���ݜ�[45Yu�nԱ%�c&�{FꫩyE�w#-�Rm�WWC{i��N�bn���*����S���FM����,́J�O&����c�)�
�����t/T���4�����n�)�I`ض��Y��T-���ze�(�����"�t5��-�Z5�zH�C��pd��̵pK	����B. �ʽz�s�K*���ztX�s�;-��wEJ�x�r<:�VH7pH��3,a�x��a�sp����b�PÎ��1�YTm���Em1k,KA��*��KZ3�hv���y���{���2�a�9��t�+��+`�* &h�J��hŎ� !,[�3!�W7�gu�lnmֳ�lR� ��v^f�(:�m�*��\�Ǚ��]]\��B��a�g���s�j�=����L-�%)yq`��48YF�8�Դ&����
��NH��ʬX��M�`��T#n�;����M�o6��ARU�L��%C[`���f�3	Yv �.GPO]����ofk��k�.������@���c4Zٗ�ѫܻz�GBh���b�6�5fIZ\i�/NJ�Aͤ��M�.ߒ�0�w����ȅ+��V���+�!��<*� n2`�I�mn����SN�T����6�d=�Y��c� ���j�*I-���p�Rt#�bqb��ܪ���H,����J�C6�M�x5�ݼM�B]E�J��d;Wtpm��*���_Q��^��_��^�E�b�n&�l��ԀU�͈�{�0 @�������{,%U�1��S%�gQ.��f��3qޒy%�!ٗ�u��lfr��h�ĢY�����[Ht  Cؤ�'c��c�T[Z�p�}���ɩ��NC�K��b2�g��.�ِL����)�����s����Ћ�XÕ\�%j$▲+�7`�&���ѱFm<�����̡p�$���%�~��
>=	<m]r$�m*J_��B��Ҹ��#Bі\2��X����n+�M΃w��Q�*����36����A��P�
�M��ԱZ�� �6�]
�Bt�tk6P"��6R)C�6�����jh��	���TD"�͏��`3��H����jTM^B�l��I^��P5�̡˻P\[/j��Rn��n\�M���M�nՙ�ʽ�ցE+:�\�.gY�7�)���×'-�7z�Tڒ��mg��ت���ct�4��6-���/����q���p�o��f�sissiw�*�'���������I$�I$�I$�Fd�.v�["h[����3�2�m�=z�@`R�����zV���嗦�\DoN�I֌�w�jC"v- ��7�,�-��V�e���uɍ|��\�θ�U�e5�WovǕ�����z��^Q��Rd��Y��a�f�2��#�tT��*�N������yÛ�ǁ˺5��Ӗ�9.�Ý��8kXz��;��̆��xH�
٢ܱ�2;]!¯�Tf�)�2�-KvX[bUI��,��)$�t�_��y�+!B��,��2	�x��/��nY�x��If��d7�v8���8%t�"�
�uq~9|�9�96�w�{6���/0Q}4���f[�8���޽;�����!��qH�jU�c�3j�W���ج+��k��n|u��ѣ�!�-|����q��L{�>�Xĝc~�o�p�0��K��*|�W.� �N��R�UY���57!���ʠ�wR]&ѧ��I���1DЛU�V̻7�sw؜�Յs)���묳X�v��U0y\��M=9חU�U���4$��Yu�dH'3�UR�l�4qVi���&�F�y	
��UYN������E��]��xUly�E��j���c���ʽ���t��|�9�%�ac*�iӐmtq-�3�n�9�b�K��� @�wl^Q�R GٮH�U��X��<�*/�]o�T��I5#���E�m�E$��*����nG�κ�\�J�d*�>��ȳ�
���`�[��%z��� ��H���`U���.L;1_�m�7���L�9W\t��y��Uϵ�����K)���o���&Ww��3�N-�ph�_ j�T3��z�(Z�l����'�:����j���k���A�I��@���&�}���*� !<����`.;;Z�{U^Y�F�o�Fi���k��έ���}�R�@�vWlԂp���B�o@T2λ�]xZcb�0�����a�WK�EJƳG[W���{gY�v�:gB���N���y�{���(
�oGuΖs���V�M�Xi�R�Ia�2�s��X��T�[���0]���8�wm�uo���Ԗe�=Z�uT">��e=n��ţ����b[$�����Ó��l�����, �;M.8u.���3��ޔ�u��5��F�#Z�+st���Ǉ%����U���b�K
�Q�Wk3��WTO)8\��m���8��v��#P;���u��u�0��j_X��C��C�v�9����z,�W:�w��o��{�q���'U�WB���n�:�mB��u�N�І��3���.:N���X.�fbͥS�Z�3�1c�c,�b�jV�=�3���u#���ٮ����x�­}�= �+J�m��y���ԍe	���z�Irpyֺ�ɝ�_q�KD��oyEC0hZ�(�,0��{�\^�U�I�Õ����ҸCX򋤱�T ��I\��u��V����n�`������Z��DOM`�v�q�ރ'9E���$4�k%,t��b�;��Sf�	F*���u��k�m��c�:9Ш�J��ŉYSnc��҈b��
� �ܭKeL��E��p�b���<�%�[q��ٵ}�+X�v��4M�������Q�!mf����ۃ{.�q�p2��:v�V���s5��hY�
�_>m�˭b:����nNͧ��91n�í�
7o"�t�^�b����u�2���m���KU�vvӷ�n�t�Z-t��hs���bݲ���xz�Vi�*'��vY�hݐ��<����.�o��9�E��ٺܠ��V^"�5n��+	dᵮL�\�F�n��ލ�u-���Ksr� ^l��1g�$�7gT�k���k�E�ҷnSns5i�R}�b١��M�#^h�.�� �WX2� 5ԚV;��q��ᾞ��fV�������H�Y�����X��)v҇M嗭�;Պٰ��T��>��=so(�]���>�Ć�X���F+R3�bǬUNiV�%Zs
�+��9�2�S���L�2�y�"$�Pl���w]!7� �`:��C��3�]����ւC����!��9�p�aζF)J�f�-�3��p�Sa�=2��؊f�ɬ:{[�2gIj���qM����-�Z�D���eX�X��,���ȇL���?+d��#/��ݏ��ȧIb��3*�)���@���=+�����R��U�릆��O��JB��������<���V�-a�h̵;Bc->���I�̧�l��ˡ�pp��<���f빩�/�J�p�h�c���L��/�������C�f���b�uC�e�`�i5Y�7���	2����y����n�� n�Gi���`����s���Ɉc`�S�je��<�m'��h���w+"��]��{s9Sy��z��������:9>�
���a��No�m!��ʷ��s��Я`�CX*:j�]h�u����_h��DD�f�5����j
��R� ��sv�Cin�1�r�J��,I-�$�C��*��>*��&��{���6�l�V�ۻ�GoQ�޺ŝ�z\���ZUU�"*��H�VQ��U6�C+m���x0�D�R��
���w�����q�ڂd�k��&b]j�8�U��M� r��I�j��E�}��(����MRj�w��/,�V�;5"㡢�ގ{@�2ܘ�Egm��F�o7�q�oc��r�����e�zo�-X���7b���dF:�,A]7T�e�4�4����쥶;�1A�k܆>�����j5�:䡕�ͫw����9��nF��!�z���Z��rځ��T��LM	n��G+7+R�s~�)Y`�9W7��e�[,���f�t{��us��Gb��`�r�e��`�6b�����@��#8/t�{��6M�u_���:nL}�h�Τ7��k�G�"���S��Ǥ����Φ�ݭygn*Jk^�������.��yٻʂW{�KV�Z��E���sb-W_1�,��)��35R�;r��s9���r�-�q7ץ�j�8pQYhiSc�{SuX��ua���f�{-P[�����h�e:�p���<ʶ$ƚ�;3:�P5�u�Ɏ.�-<k8��V�}�#!r�u�6��l�C�.��ٴ�ԍs��~������D�0!��W�J��k�\[Ӧ����6�n�ݰ��+v�LXh��T���I�v��z�7V��ŷ������M����d�P�9R�9'V�i��Z���-ďJ!�K�L��wv�vۖvL��2v��r��L�I	˩B�+��T=Z��YɺxΛTȄ�COoLSj���jm��t����-�M7���,�R�Q��;�kj��;����(q�-�\�0�u�n�ۚ��A��Z��C_�2��?7�Ҹ�^<t������k}��L�B��&���;�}�̌�b�R��҃1���о���w��k�RAH�t���މGe�	�K�G�z��g}�j��خ�M�bL�ʄ+��Z.����F��!�i��Y�����dCS&����`6�Sr�jh��QU���/�
����5<�	+(�M�UJNx�۴�W�f�P�(E�5�"���yKy�ׂk�kmm�DՐ�n�xZњͺ��k�;І؋�d�(�x:�eߦL�grװ�㗂���Q��pʅfkd.�X)� s�*w�
��h]{�کm�[��ƹ�+]å��n����P�fB�3�e�C3��C>[�98�]�S�{�r�.�J�3r�f�k|��z�Վ�]	��qy�L����ns��o�=a�I���۽���V�ÊgU��6�8�$sM9j��EF��$]�rQ��,-�Bܼ��sz�V��4������R��m#���B5BȺ��
��j|A��&�	�bU�����a&��l��bj,5Kuٺ�� ��h��MVCQ����x��fH�\{�v���������D9C��T����v�}�b��!#j"���4�)��t�W=q�Pw�=�Xy튗w���L�Z�q K�W�=�.��b$�g*c�"�=��Ȥ�mke���95�A]n�ݾRþ�b�/���4��gp��9��A����#�8��9c.�\s�sk���	;��|z	
�Mo1{(�r �ۚ�N6���'9��N|�2�e�rwx=7[����d��v���|��a��Ӳ��b�����]�aZ�MJ����X0��7Ms�I7������a�yKs$�*�ƈ�B��~9g���*)[>�����,t�1^�ȳC�9q���K���&�1��AQ�̦�8��M3z��ɛ�VA�:l��=S���=�s���"ѵ3�9s�A+픎�,GBјz�p�Y�Q��GZ�0��	Y��X���}]�ԱJ�9Q�0�ݪ�}���[h_h켈�~o5�-� ��{�Mu�d2&��A��S`b�w/��gL^�V�b6�L0��>�ם������v�0o_ktk��KÚ�k�s�m�t4㕼%ev�ti��h�R��aۖ�VV�}DI����%e*~��Uc��J*�r��8/�b<���	�/�U���0D�2a�\��r���/F���~��1�z{(e�NdÓ獼w��>ǉc�~��I)��r��Z6�/ �S�u�vS�ډ�ŷ���S�a�_f�L,�7hV2k�FH}�np/2f㛧�+��C��;CnF��`�|\p)�u���v�I��mR�֌6��-+ŕ�zþ���BN�-�Yں6�T��KT�{�^���cz��ڟ&�5�ЦS�V�2��Cr����l�W�k�rN���'T�|
辁X�����]�|�!Jjk��܀�ڵ�:�h�+]1���n��b�e[8��D+Rw�ڤ�k�Y�Z5�D�����`��z3q�%�^:���T���v�Y.���s�f1�e�� ����uO�sw}��'yu��.-J��D)�Z�ַ�ЪK��yX�Kμ۹f�-�T���e�a��\/qY;z~�(I�R�9���)	����)����C�Acs���r����[DV]77��,1:C�@2�����7	y�VV�H�in��}��� ,�Ȫ��jt��0��)����7{�j�;Mm�n�m-pG�1m�ڗ/����W�1ǎ�t�U�ێ7�s%Wl��Ql������l��3�ӣ�1�vlg/r�R�T��w��������r#[��+4�0S�������z��Drm>ْ�1{3\�PBW`�0J
m �����
��	6���1���䒣�{5D�V��,}�b�7C��#]�Vs}��0eR��b�|=3����o47ڐWR����(�-�d,�SV"��98�}���xDq~|��%}��4Ív�v�7��*��D�稼[fN��g�j�Bʡ��ͽ�1�{�T���u��n<ł#�-�X��b�Ct��r|+�3��A�u�+����]j��3�&ۤ8�N�m��I�n�����m\*�= �ug�pw�n�[]�/;W��R���"�=���ȥԻ�ei�����M�����n�f\�;X�N��h���*�P�;N��S)�0e�-L�	6���f�g4�[�ͩ�}�󍀯N;�x�͍���}U\gEճ̖{Rܿ'�R��]m��Vd>���=���kn6��m-ꕵw6:��G�p�4�z{):�0X�����U���M��՘r�/���y��n� �gZzl�Cӡ�^Q���xu̓M�`8�v-EQ�;(�Ժ��ݬ�id'T�{`xN�$����<�K�Sx�YR���jDrǔ��i@���{�(p�̺	��E��f�A��3�ە����wV���
��oIrG����{�$I6l.��Gb���e�ռ��{�V��z��R:"+Rs�׻��X!s$7D����cO�}}�f��j�i��[�b�jj2(4�oٛ���C˲��Q޽���
��S���R
��2�kB��e4�b���ëf>�K���������bSZ��|��5�V9������,���nk�[5��;���v]���^��u�z���w���:��z��j�c��M��]�[�4b:��53d���k]�A �u��v��Q��'T}c7dvd�e�yK�G��a�h�f%.�s�Z�z�z�]�|7���[W�p�j7�����
�'I���5.�qGY�Dm�x���a�`�d��H�.f�n,4Ӕ춻*f��c-���V��Vw���F�V;�O�G�/��#����4�%]R>m��]��ɯ��V0_KW���|�8�H�C��I|Kؑ�GIU�.1<#���Y��Z���hn�ڣ�.�+�3�8Gw���s�9�0J�עÃ�lcQ��2�����}��:]�0n�u��wFj�G7.���J�Xu�p�j��N�Q�=��7��J���;:�t��qȳy%��_:�	C룐uS˗W~����0�vo �Ύ�SMT�x���y��"��z�1�x�y� �ݐ��я�Q�\?���S�/9�r��9}�������o�}�@|��Z���OwR�:ϗ�~@����3��@{���{���!���}�ݾ��w'��t{��Q��	���;C]w�޷R��Cu�/��{��_
�`kG�z�v~�A��7ξ�Q���G�'��(u_�DAw�?���U?x߳��=���g����f�i�ͭ~�χC7���G.�WUwW&���o)�')ᱛ
��8�����)�{]8�@�Y�To�l<7���ڴ,�l��g�t�:0�U�tU�I��˗W�B(�\Y��dn��bw�i��Vu�CkȻʾ��V�����m��5�S��� �W�6��
[�xiT�2z:��Lu��� ���5�<n!�&�O؞��X*�݌�r��ncI�fu,Hu�5���BV�m����J�:q�\��P�}���y���!�[0�'Z��)�r�D<��
DU��̻����]��־����41���شN���� ����sڸ�V*��^U�A���_hq��m�VO�GǊ�T2��-�#�0pL��/tR��G#W��Y�F���%,8�}so����O׭�̼m��̴	C�мa��V�*�]�F�b��@[���Č��!���y�v��l�uco^DW�v�+Lv1Q��֟B���A�Y3�V���:u͡9B��N{�}e�;*(���uf�c���K���Q�rqw��n Ӭ]�R��Nk�n�r���w �]~q�h�	��Y3���9D��>/����Ӯ�ʲ�h{j钵�؃���Ll�$�tz�d녡��dOYLV]2,�	e�G0��K[��{;���^%���T�7v�u�,4��r��p>�t�w��d�ά�,�����������ǎx��ǏO<x����<x��Ǐ�3Ǐ<x�����Ǐ<x����<|x�>�<x���Ǐ<}<x���Ǐ<x�x�}��o����Ǐ=�x��Ƿ�<x�x��Ǐo<x����<x��Ǐ<x�<x����Ǐ�o=<x����Ǐo<x���Ǐ>�<x�<x����ξw��U7r[(�C���wK	X2��6¨�H՘s0l�`:c\�1�5�J嗃9�{\���Fm�oy)�B�@r���K�h�x�9Tݩh)܎l�����u㳙�$ɗ�:�B�B<��f�`v��]��@n`��C�D鑝���`��+Yh��:���;��L! �<{��̋�^V���-��.Q��`\9v�����8l���=y�-���<LݙQ"p��p���{2��.���G�~��6��q3�FƼ����-!u��zn�%����rN�0�<��*)�^����rM[2
 9
})]捱A�J]���m!`lqx��곜�=�pYk��	�w�b]Ƶ�NtN�-x��k��zV�Ħӱ��x�&�e�x_wS�l1�E�I��ZS6�X�Y���xkF�"�a�;��T�rҬ���J�쭃U�]��:��f�GE�6��	C�ν� -*���&�Y3E<��h	�Mfn����¨����++�ϸ�����������T�
��o�m�ܡU^=V0ek냱��x�92�2�4Û��,/;�I�ڒ����W^$7��2��i:ك8d[dt�v\4N�-k��K��Wt���X���yՎ������}��Ы�(+�f�W�ĒS�;{m%e;�#���u��_����v@�Ry�Kxj��Ȑ6%��ƅ:��r�un��:kMJ0ɫ^�Zo.�ğ���í�~=<x����|x�����x����ǏO<g�<x����ǏO<x����Ǐ�<x���Ǐ<}�x�<x��Ǐ��<x��Ǐ<x������Ϸ�����Ǐ��<x��Ǐ<x��Ǐ3Ǐ<{x��Ǐ��9�Ǐ<x�x<x��Ǐ<x�x��Ǐ<x��<x��Ǐ��>������j.ֵ�u}oqF:�tG�;?5sZ��q`k:m=��bUïf�<+�怜!⦕�:yKv+�aQ��`eşj6mfW;VP������OjU�a�m]������R���6/���g3�6U����vR[�v�CV3V�=������8ֺX���g��{f�'C&"��Z����x����m,��b�9����m���kt�Y.E�@����Ӣ!�8W+
��뀂����ovrwC�2ތ�uve���@��mB�=�Nc�l�[K)ʯ��A�A]ut�N^�P�IU\�pv�����iV�X;v	t�ø�Rr��®����C`�Ģ��k����;OngY!���n��=�<}f�@/��7�����s"Uw�ɭR;k7��˸'fU9�Nr͗�,U)l�Zn�9pb��PS1:�f%�U���Dzk����Vu�[�Ύ�gV���欖�mk\�W�x%E)���.Wշf.��ó����M!Y����T�aR�cۖ�����Vh�ӿWX�v;�E>s+�r�󵋗WJc�s�h�*͢�k��d#X��.�R����v��c���vs#6>�[*�5�F��]8y����`��o��$㵷��h��	䓗��N�LUu�CT�4�Ÿ3v�V�@��4C�#R������N�w��v��T���ڽ��0�캊Z���ʹ��p����{�����3ZHc(�]yt��0����,1h4���U����%L�7l��]�g>p_N�o(�;v~��7p}[�j�8�Q�U6	�	���V�4���5�1p�Y+^��cr:���`���5+ki��f\�]k�G:
o�X|]��Z['ªQ�L��q�*8D�i��/4%��+�B�V�����l�a���]э+�Lp��Qq��*w{P=�s�lU �̾����ʁ`�.�ӳ��:���e�OmK�T������P8ň�U5[�wW[Ä#y:ִiB���ڶwܪ��'J�EsN�Z��}�g$�U�0R��O�c�F���y:E"4�O�锝-���yHZ�*���*,��+�`�G��/`�zN:J+]a��l��-�+�g�DTd&k�"�S��2�z��CE�bWO��D��էHW�L����D��Vx�7&�	�i�gA�ëh6*�s��%嬛�w|�Z���&Q��%���ﰸ��휾�C7WF->�в��v̈́��&��2����	;�qp��v��5��H޽]zr�Hh��Ur��Ve9S�v7ׁ1;K�̺�P䳐�Gתr�v��pp�;O�|�r9"���B��I,u��;�|� ��j���R0��oI������֎�,XT��(+��C�0i���Wh|�k���h)7��I�{2�"inL-�&�S��3��>#�Ioan�e0��[o�[}���%2�x�����vݶD&�B-G�LȜ��!٣{�����(R�[�^n��hٹyс�p��N}N��G�7)�H�x���Y�r��ي��Y�,M�	�OԆ%�l��MX���OO�!�ҩQ�aɝ��w8�����⅓g
U��ޤ7�{��l]�n�:J����]�ֶM"V��
�8I	����|��dS�tN��f�#�j!��uV@2�Y�5<�J���L�w�P)��(�mm2�j#�F��q��d4�W,���d����R>�6�N\��˗����g,�F��^�es}�i�����P\�,�]���	�}��ZJ�ĸ�{���C��-w�r��u�}��U}j(�}��69R����v)ט��=�0�y��Iw_@��c����r�ب�k)���	�&�7���^'�%ɼ��I
����������a�s�xHC�צ�eA*�i�od���gi���D0/5��+�u~����ǐ�)vk��&����ד
��漳0���1
ޙC�-��[].��8&�E]�N+^5�`NV7G�_,�%��{��zmf�����RKk�#J��УmcXC��ʬ�,!ļ��S{x�dR�]�E	�/�wK��N�)�q���0�b�jY�|���gLg��O����+In�fn�3�l���3����ӧ�i��űWD7�tU��ց�\�,����X��9���O.4�v��o��e� Ws�[��(�=�{��f��KD��[�����)�u��M��`Ⱪ�Z��L�
���whű�����l�ce�r	-�5���-���(�s#t�xldȳC�����v�*�G��9�W�5v2ۛN�G[əC�<,��-���ۦ��;n��<:VP5	|.�V5�P�֥BF�}��8��گ�p��U�Hq�;�ĳW����P4���v!'�/6�BC�"�]1H�y�j�k��#�[�z�#Z=�R{�Z�!����0`|X���Z/&].�+cFm�g9i嬠LK}!���<1�vSyc&ֻ�]wG/�A}�x<p-{n��r�	��:s�j��)B��b�j����p��)[,�e����mZ9���U��~�|�Qv6�eE`��Z�$!4L[1"�B��sk�U�`�Ƶ�oz�.�^�ʕ����#,+YO*2t�쭕r�m�jKS�B_s�R�N���YZe�cO$;��-ƣ��i��α��m�Z�p��hLQ�nZ��`�vQΝ�.�t���x��)��k;Pa�m��ԑ,�Sͼ�7N75�J��G2��k�eG/�"�Rxi�}AU�uwe6�[ba|rbǹ��bPa� �8���N�guĸ�Ǆ��]\Z���	iPQ�h�0�N�X�Sf�Z:p`��Z����f�|kq����ec�i�Zs�1�;ڻ��oWE��P���7��靳��V�Td������l�񭉝�	��f���ue����l4.Q������{�@q��h�'d2E�+�f�:sc/v^���<�*�.��:6l���Wͺ-�T�������ѧ�F�K�t3��
钇+�pj4�î����}����.��Wni}/:��Ws�����O��p���_+?�óU]�(9�m�'�jY}1A{�ko�b4#uv�1����c�-�Ƅ�T|�D��u�$y;�d���ݲ6l]5�=4D�z������k��eċ ZUz)��J��=l�Q�]��!AA��8:�Y@�؎���܇]�~�I���^�^Y\�*�ge^����=����},�Q��*%v*�P�TE�[�i�����o-�+=��%�4q���ɞ�s	]Y1��\x��=�f�w�	i�x��
Ɋܽ�=[}F�f�x�	m\P?T
a=ʣ%e�ԓU���C�"�Z����!���W�o�kPM�]X^Sp̼���Y�i�jaE�l�S����{S�{�*�6^WP\:|�L��֚2��*_nG;+4���lW����u7��
.�h��h�Zu�!ͽ��W��%+���F��R�I �lut˺k]^�/fE���U��oRa&��Ã�[[��1��9&�tr�/�����e�;���rԳ�(�sGpS��p���F.�-�^.��u�8�]G*��ܽt'�=�J�9�:��F��&����[[��.��N+�ۏ7X�����QX�5{r38���n���:�yc郘�w� 짶Ӊ��
jP�F��IN��8�v\AY���aa��|�V���4�e-yԋ/dH��6s8m�X���}��S���yBi1��s�{)V�
����=r�69ut1,C�<��Q�Q��B7����E�)�]u�{��\*X�9y/l]C�;��N��^�I�CO+�B\��^��`uu�"'�j��h�|��ю�r�ɱZɉ+�q��� e��f�.IW3؅_#�}G	��#ϱA]a�Q}5Ѱu��r�A
�w��|7����І���frݫ\R��CT�Wm��Y���t��L��չGH�6K��_<`�$����VhxGp��ǳ�a:."]b����LP�Uڙ*�MJ�,���:�*S5�'};:�%
��)%بmh&�U�s�T!1 û�����CC��{�®eZ���+�W3Y�:�1,��TB��qg����.����]FNʖ�����!��S�ַ�Z����/W��b��*�eņ\=���bi���Eoਊ4na�=��lw:Nƅ��Rۮ�Ԉf��S)��+k�u8*Bκ%�9}��˲�0W! �n�`��S�`r��Ps��sK�%���B�9�:�"�
-Wہ��7���9q�m���(�#a�(�b붶XFo0��l�v�b�ǹ�����1I��W�m����>˻�`´���W[�wX�uc�V�4�jv�d�u�xv
W�ԣ֊��MØ�I�9[o����0Zr��ݖ/(v��)Fɫ��wf�]*��u�M�܌���R�'�Rʝh-4�x;γ��}Bȭ�OvdMb�Me�t��e�J�/��U���v��
��-��a4s�dk���Ra��'V�lb�y��!g21T��5'����Q��^�JyϽ|�0u��
Re%2��S*Je�7I����l�[�%�n#+���g �I�坮v[�U��snZ�)��L�v���UZ@:_��X�̢�ڋH��H��{�T�MvY�Qw�-㏬(0v�B���k/�����E�ڏ*�=)�<��W9�+��7���J�T�y'ٮ�K�	�BǟVv�,n����LW�h29���(�J��޴쇨쩧��ݤv��7W����jL�s9╭�����xWjJBy�yw�����73�:A	%VS���0�]��<7�j�]:�v�\.K��c�_)JX�3s���w�]�nUK���F˷���w$핫r���*�b3��r[���ř�8��1R�U|2���e�5��R�+:*~�]�p�����Ͷ�jvX�ČiQ}Z&,�N��fԵ�'�V�雼���\�!�,_����{	�)]p`�A����u��s/��;Yc�)���4q<���f	+r�^�e����l~��=i�]�IT�=;����m�y@2"��[�B�5.�:|��0SՎ�6���y��O/2����n����]A��v�Z�1,�TgSN=̭,�P�7k����6`�;�i�M˳b�f�rƓ}�u{v��<8q}�ld�iW�a��ݗ;b=�n�p�+z�2`�fS�̸�F��a:� �-�Tt���Y���w,�I�
N��Z���@E�Ѷ�=XF�9:���S����G �����t_���ܴ����S+�@j[Xe�:O,��-;O/l�Ż#��.jV�5��b�C�(�����!�45׆P�%
��Ԣ�vѩ��-�;��1�q ���uz����
[�-#�����zk�]j�F���?���������/��w����5�T�/������귣�Xl�U4�q�l��)0�����HQ�f$�e0&�m��!P�G�:m�NZ���A�H,�����Qp�d�!. A����U��j�"Ya��.C�0��S��1�͹N�A�����9�G�L��X���IT&�[5�|�"5I��/m��l2*�u��Ҹ��f��<��Ŏ[���s�����N���h�Z�	3&vS�rTj:��y�J9ˀ��2�\a<�}��:T���8V�1t�,C����*�w#�����*�������y��
\���D!��gX��-�r����f��7�S�i�[�*`�Mu�Fo{C�1ތW��\���Df	ۖ��CN�m�&L�u�r�k�:��by:M5�a���6mH���z�o)0��y�Vk{c�e�X48[�.a���@�͎H�BL:�=�8%Fq6k�򭌨K2Qf�9�H^:q�@(E��
:��s8~l�R���48�:
�\��d0iXʳ���v��-a�i7�mN��0�y�[�StKΡ��T����R07�sDvylWA����lv[�^f�w��*����hn;{ǅ���Ԩ��l�n;��7��p�Ʀ�� �nc`���B�w*�q��uƵ=�U��Mz�y=�sQ�h�`�+�X�L���X=�*�dP�����]Oa��X5��2�CE�z^�؜%L��L�:$�&��5(>Uj�9%�up�ɳ�=��zM�#C��/��X����S�X叩h��a!�О��:i}�â~95n}����QM�I#��?��̡	P��:��1BTm$��i�4��"$$�J��$(�L�	�O�E(`���S1p$d�����m���M�?E��r0aO�e	rAZ����#-�$-�B,�"1@��!L6�RF�7�A(?�8lơJ�_��`,0XDD�(cI&4�)8S (� �8�R@Z�LR&JUA��Dg��Bc$�	*���� =d���)��WO}wgZ	<����z��RDL��&�Q���mMm�(*�Z:Ʀ�"(�*��v�=>>�>>�?������|x�q&�(�bH��v(�Tm��h5�m��6��AEiڰPD���v�=<x�������~?��Ǐ�$pƃc1kSA	:�4N��UU@hq4Rh��h4톚	� ����tUѝM�"�֊4��
�g��(��(��ET3EIr�e�F��Z�E30{�[kQz�_sZ����*�"n��Ѣ�������m�CDT�C�uS�wi�����&���:����AI�QDUAݢ�Zj����*��f{a��h��*"�f�c��u)���`�H+`����:��:�1��M�V�':�Q���ulDh�`ԛlXƄ�v��8�(1m��6�F�;�F���j*-�lgVذ:1���A���3;i�-[kK[k&k"��֫:�Fp��|S�z����]���WF�u�e�!uf��&;��� Ks�fhBr36�Z��Y�+���Rn���9�*�U4�w���WZ��a
���8���j��]Z�1Q��l��D�d@�M�������HMN&�(#��IL�I�l��{�ޢ��ަ��D�c�+�l*Q#v��������
E�>�fμeȫ�6f��5����{�����w>�\C����5#\�zI5��ܪ��\�n��̕ף����5��G���4���p�3v�C^8�$�1Ơ������9ͻ�3gn߆�3z�Ɨ<;.^�뉟{ҏ���y�����@�{!l��ť6�1�b�,A�������/ٮVV�U��t����_��8�� �I�g&|;Ξ}L��_�e�3�7��R�q[�pr�G�Ux�>o��g�^���ъ���/���ήv��)ڂ���y`�L�}rL���=�n^��o��(���z�/�W�*���&�3Ǡ���λ�{�<���Ǜ+��s�_=���LR�Y�2��NS)�A�0�����q��T^�l'Hc�t4��{_���~�\R\�<�eUH.�{�"	����)[y��c5�r~����fKR�[س$FXׅ�Ov�ٜr���n�Ps�vc
%�V	�l��+�Z^��=ǡRcҷ�BzK��䵯����Zɷkn9�ܫV�rY�CGٓ"J�i·�{CŢ�`1_1)J+b�Ǖ��]z�N���j�#�ܞu�n.��~�d�b!��ߦ��1�M?W)~��%�;7�S}��׶�zL�5�����=� �~���q��G�[���3*�I?����ݑ�\cW~�Z�kࣰ9w��������*K�uo�;ҍv�Y�䕌�T�y�3�Xy���r^�Vg2�a �<{�M��iW��sػy����|���p~��C��<dFou��"����\ӆu��T^Y�K�F׆��sK�����\��C��g���}��x5d룞�����{�ɣ�=��{���y�bw��޽b}��4�̍wg/o[������x݁�����l���Ns���u�৛��{��w����C��H-P�T�͞'��=>�����m���Iy��)��Lbe�4-yfˉﲻn�>�y{M6�T\�ɕ��0����DܼɃ{����f���<d�ةf]Ѫ�Ư���{"N��"k�d���dG(���ܲ�����|x:��0�P���E{��]��� Y�������'*TQ�u,�j:;�V+}�wh���0l5���`��fɫ��:��4tدI�zS�L�P�W��w�ޝn�{U�%�C��,;��,�Zx����OC�P�=��/�q�K/�).yJ)�z��:�t`N��ݑ�	^�=������?eee-z�W�N��I�����j�
���~�s��?v�S|#�����10�#r_>*�w�[�zc���<�S���t~����?+���^'�Ķu�D�/�2��=/���W|ֹs�Ȁ�)�$ ���̗YF��r��І6�o��{AX��ܸ�K3q��3K��mj<�9Ep�����uC�7����U��J��}K�w�8�fx%�z�l�7DU��x<�8z��8�憐�jw2̀H#����{3SӴzs��A�ȸx�
�����|���ޮ�ߍ�;/����wh=xi�x�y��ܶ��H��w��E:�W��f�=\C��M㞞u�?v��X{k��u�e���sH��,����K���ʘ���%"�}�D9���Þ�qo�8��Q�2d�cj�Va\�ÝQȨ֊T���{M�ٛ�`x���	k!�}�3'L�Ȼ�)����u̞j��>��,�٢�=���Wpj�Q̢�s3��\��Ƴ�������$�0x�r�F�9�k�����-��bMm3'h�K8l�0hG����}�I�s��&Ox��V�}����E-^��`�W��!μ�}=84G�5�ٲI�;�6�O���g��~��͘:�=OM�����?x�6����G�l��G�V���!��̿<�ta�T������=�TPЮ���xI��<�M=�|�����>Wݮ�\z.B"���߽$��_�4F[\0��x�ޟDa`swCOM�e����<���ss4g��nZ���S���A=\��[�˦����aO7 V����^��v��Ǻ��v� 剝����X��^�p���~6 �ps������~������W���=�P^bك���z�1.nm�I�jno�>阭�I����1��%��5��IDֻλ`���r�$+_Q;�+������\����̘6�3�9	o�T~�0�6�k�(�Z/	y���D�"�4�-��s&���S�N�Q����'[ӯ���>.�	3XI��"ϥ�xJ�>����T��LJ��͹�����2��n��=�T�V��LP����#D�:Q����$��j�
�G��4�o�ߓ���D��_�^���k޹W�0�X�<I��ڣ�	��fg���5g��k��dl����H�����=v�:ӛ��'�;9@\���;C��A��=Xy�|������򷖭1M�^�c7�F3_e�����'�lɣ;�]���#����F[9i�J�a�}�+N��#|M��=D��7����۽�nm��m����*/z�X�~���k^����Ǫ={�+<E�v�6��}�2j���8�c��>K��_��f�kez�>Z��~��9^��?_����t����ma�ì��r	^5���k�(�y�N}3�p��J��<���,7��wg���n���]�&V�
�S+"��+��k��V&�N�(*#�V�~�&���K$P0�_t��t(���`R]�f�i�HKړk)��Q�ܵ�/�UcϾ�n���fx9�]�U��>�w���q'7�t�v6S�hb��ϦS<S�py20��(?�q��:}��7����o=�]c
��%'xoM��Z���P$xh����UMt߰��m���=A���I�=�R�F�����0��z�x*[^���������{���y��9=�z��.�^{==ނ:�����v֏`�*Xb�bQzQ]�-��v�U=�-�q��d���o���z��d��1�����	��
=������Ya,qC�ז�Op�p�ws��/>��K7����$8y��0z1������pL���^���xg�5z�~���ſ�y��N��{���la�;ǻ&�{��[^�Z"��򞊯��73;+qOH߸�~Y���?���6#���hFDf�7CI�@��r܍�L�ެ��ph�%�GǷn��u����8C	I��u��j;zJV��:BzGZ�vt���H�@]nQ�\y�s��#$�U�B�=�ʶ7��l���}�A���G�7Gw�ftR�.S�3����̰���e�ך.s�v_կq=qSL����]J�����A�κ��c�i��ޚTeyd|4�Gu{}�K���	0k�6�X�c4�:��`�{�gy{w-R�m6��W#x{���uᮑg� �;�t�k�:����	���r��������ٳ��A�u�Y�����2�ۺ��l��u�팱>=^	�aO'OS��q�|��=BL^���3=��g�3GH鞫�>��(���n;����/J���s|���[�0��g|�k���E�ܪX�Aud	ؠ���9���^�ks��X�B�|&<��+��"�v���f���Yդ+_W�@��9d/Bo'Rt$�|�y�Vk��N{��R^^�����z�{�7F�43��nci���9R���Κ�qtky�oI�{�1�uo6�B�cfMY�f��d�]����%��Ӿ�yy���n	�o��\5BR2iK��;*�]ޟh�{QHq�Vo'���%�;��ڙ�S��|zN���H��]�����:�Z��=��2�5d&iA�����ګ�t�.s��9$]�<�8�H�PWRV/�;ӵ^)����������Ă�ϥ�s �'�X���L���w���9����oMx H��F{�6������99�{��w)�E�e�E�g�x86K�~>ǽ�^��Y��E�j���S�fG��u���<�wwz+�4���c�V[��[@���W�]6�����>�f���G'���~�����U�=���4h��u}���;M3v"{�#:������>�ݝ~+K�0p�1ч*��s5m/HR<+�}^򓔩ݩB���[����+N��49��&��T�D����4pS���e�9>�y�c�e�fb�9��3�����O"��3pd.��{���F��ו����������~�r�k��~��Jc�X�V�9M���|���]����<�2�h�ߌ�ߞ[���].�����L=���S�m;�G�d�ǂǆ/+�-��3���Ǉ��ȭS���vn>�uű��ת��t�[O<Y\^�)*�����+k6�8��}���mGS̀𛶦S�)i�8U���y�c��P+���D!����1H���2<R�'�u{[�m5��~\�pl��D�{=��G���������4Ȩv
��Y��1��oڴ{�\��ss7<�p�6����s���-	I�iR�y/�\�PU��
���~2sڏ�D���{�hO<so{Շ���z7���C�����?zJ�����崕�C܍x��I�K�NN*�n
�k�xz�5C�V���=�g.���51K�W�i�ro(�U�9�����n�Iq~��vXں��>C��No��=���	a����I'd�|Ԃz���C|��W	w������w��������a\�3��U���6@�DO�p��cb���n�w^+T�ÂV95���/،��)�y��7=p�w�OY�|n�q�i�{�gf��s�!�O	���=˫�{͋\O��C�*�ڤ������-�ʖ�㡍^f����gz�ea�(�p}[��o;�N���L�1�p$����R˥[���H�t���o]�Ԣ�[Ji�{\�b77o������j��ƌ{K��Z��Y[���q��Z��$���iG����;.���ݷw�Z{��T�Ģ���3�Oe�S����>���/���y���㯇�>7��{��䴴7��������X�Ƹ:j�5P�Թ�<}<�tEs7����&	�쥏>����$E�:���x.��n��a݊#;}3|�G��N4V�44��c^zζ�l��ir�f����u��}�a�u�� �s�T������87���`Ҟ]_�R\qn��(���n�pKѾ����S.���2�Γ�\Ͻ/~������3��<���}݊?����M}J�J<��"��I��}�7�&���7���L��̝�:��Dol?�i��1�|�����A~�wW��v�}�����r>�W�4"�3馌�)�EK6��~��g�m�Mv\.���W��m����s�l�{�!��R��^�Z���|>�p��X������)D��XM,o���5%w(��wk5a
�Y��d��bFPu�.��f�P�',����ko�`�vLӫ������KN�w�'+��p�-�j�Ს�ҧ\՝�{`��#���l3*�4�h�����x�f�b<ڥX��"�<��X�
KkL��h�g M��r�L?8Z�kh�X�7Ưo�η��~ŒK�Ga�W�h;��m��]�j���c�S�Hd����O��2
1pܩ�E��*�Ϩk/����^�x�EܗĲĤ"�x]	��r���'Z�&����A�^�.�a<��z�nQ��SM�[l�Vˬ؈R%7VΚ�Vd�/Q�Mddޫ�*D��r.�T\�I:��8�݂�J���AQ^�[*�it�DV��g���S����ݰS�;���t^����w65}j&����oj	�]��k���m��z.������҆?�#x�͋3WO�,�h��ѧt$m��/r1�50̍��8�4m�*�AƏ&��r��sf.�꺷�_*��t}mV0�JYIVCO��{���.
����͢�hΉ󹏲�m>7��N����Ah�b��\�
@�
��y������:�	�!Z6��d��u^79���4.��;%ɼF�w�c������ˮ�m��R�&q���{V��+���fvj�ټ�@��:�r`�����4['`7�
�톬�峐�<�kev$��^�a;~P�^3,��W�����ы	p�,㥟~�׻�}X�*�6t|�9�=�mZܷ�cӵ�c�Z��CJ5�L�k5ъ�1P;|Zyuֱ�M=��&�A.���n��Vq=yҘYG�ir�ד7틶g^fq��˒�b�n;����۽4�3�cn�K8�D$C��{Z�[wo��������o���-��km��ʼ����+wc�Q�x�n�c95�*���&
|u� ��Ê��73Y��ET�����B��OgVq�f�89�[՗oi泪�X	lt͜���9��%�r=��	�]�i��.r�
X">ަPķm�k;�񋒂̨�W!S��7�r�<(ss��=A4�����K3vB.�0���T�+���73���24;gt�F�+GNDʔ^��Щ�2��C��ٚ����]�B٘���{��u���iu>�R��������\��qC��nJ���"eFr���Y�ԋ���
_PǞ��[˦A@NvY��Ox���t5��w���V7��w9��j�!9{R�Ǫ��>���n���Uɣ"�Gغ�v&��g������s�з��ji�;�������2�X��oEL�$`�k�ӄ듮u��Lf:�Y}�'����*(A��2�uh��%�o;9�n�\�":癲�p9��wD-n�T��8q�k_r��(�J^o�U��A�m�mX-j�몌�2-�_:��km�Y�b4Q�����k��u81h�'j5��ӟ�������~?�����������[X<��I�F�L�"'E�mf�-��f�8�'U�l�h[F4�S��cRA�==?_�������~?������x����k�����4QTأV�m��u�DfMQV�m��X�TTMYɪ�bB�ER�ة�Ө�a1E�Fz�)hb�U۽�7]`������h��&-.�)��cE!��)���'�=��'Uh�PSACEETEKACE�P�m���h=Zb���$��f;���(��i�"����AMQTQ$]���v"))J���%u�5@˨�����.���ERP{�� ��R�*�(���
Z)�j%�`�d�(oFtQATғs��;��~��u�wߟ~��Gu�~�����-ef��p���rE՚�T�t�F./8�S�ɀ���LY��b�p}_W�>O]�������,Lṫu�?n��6�M����C�"	5%�[�[����g�w��s�>��e�Gq������Z61�;э���c�׻�5�,�4��,:��PFL?����y��&^J��o6�Pͯ|?U����څ?���^ z��_���^�{��)S6�e-�Y�3q��*d���3{�m��G���zجu�*�����67Cg��Q��=_Ua�ב�����}�[>O
8�J�k����3ڇ�G�,��
�/aWo�s��っ��[�|�,.D@D:�E-�W�X�ڱi���Cǌc �o9D�/i)�W�F�]�u�753��S۸ ���]�+�18�l�~��Q9tP��0=��}=����8b%<�S�+i5�����5>Eê���������-3��u���	��R���Ⱦ�8�E��q�&~/��I��y%��\Ú�=_"�.vǄ�;��֜Hz�0ѩ���XB=�9��80�{\�^�v�0���ܢ���2��'�kP{%�����K5��v�@7�,�`�GP<#��> #��[L������=���7fx��� �Vɚ��qu�9���6T9P�.��7X��+���XeԹ�A}�C�H�U������&a)�3�UJLx+')n;J���U�OS�sr�[�T�m�.�m��F�n��j����)CH"��M��MtJfe7���:�g@ݡ|E}����}2%2���E�n��;�K�7��:LK�G� �v��:��6~@w�A�?P����5�����~���K���[�ס�a�¼�z�j�ǌ�����8�a��[�=��9�A^b�L���]^�bS�Ʒ���zs�W1n����(D7n�X~i����AԱ_Ti�ɛ}�b
�����C�w�B]��z�F�ί�pm��aŜu�yX��-�Q{�ݡ��O:�a��e��]�{�����E���Bi�Lus�Cv�kϳ�ׄ���^&Z��y��5U�nA~�w�w*3xii�C�l�D�y7��ul�wA�����|���
j� ��7���	�i�/�n��i�Wq�~�C�q�mû�m�ʇ)i�[%���u��a[v��U�WXݭm�:pJ���M�Γ����pq��0|��f�c�ٳ�#$[/�@RO����25���ԯ�M[M����Gd�����?5��$�Ɗ��z���ʋ�4.3��_[�
(?z6Η[b����y� A�8�x�o��:�����
�e�|���Z|�\_�Qo
j򨶞�u���P��+݇Ed�?MJ��N�%;�5���Rn�o�I��Vu/���K�7�����h��b5�⠘�й���<��u���"�-/`��h���yg�\56饫���lG���'+�ӵB��l�z�SK�h�RsrX�-b��#/0�{	�a<\��kp. ���v.l.-	�T��U���!	��m�1�ꠧi���E��殈L�و���R�V��qo}I�.����e�;ur�{`���{g���Vy�¥�e5�́�׽.ӽJ�,�x	��d��oo��{�z�2�Cǜn:���A\tߐ�ZdA��1�Xo�k�����/��Y_v�/oLyEݳ��a�4�1��l���sp��#k�f�ـ�~||$<0|����>�e��e}����\��v�%!�<�g�
��o
�Y��B��/6�Ƈ-�o��+r�cm�������5,46.�}4�����U{�z���pEv���.����������i�NV���ҟ~��}�|ZkQ��C����-"�cSX�zi�֯�dȸzV�NK�LUG0��'X�΍m�"cLZ�F�xOyk`w�6�����@|Nja��{E�5���P6t�=�i��<D��f�i��f7��z���K��o@���gR�w��ǃƈM~g��~�fI��]�FvP	�_Iat&V��]M9��KwT��_y��9��������B���Q'�����@@��a���?{�g*�g�F��x�0G�u�;3^K�5�n<0Iϝ�٬L<z�]bU�R܊�-�R�G�C�fJ����z�:v�|�� LNf�5Ϸ#ҟ�U�Ɂ�Ëx^���S��à��*���bNX�W��v��j�ˏZJ�����J��o������g�o#-��ivo��r3�kL��bC�*��lD[.x���π�	A�h��
Ll�k�+tr��v[��تt�i�a�i����_9�
��B�5曍���{�Zb��|�}��y��՝��ORn`�����&.���cJ�UKcP�R=��PY�(��u�����l5;<��[pZ�U���C��P��)��6t�#�A��J�j[�
�"Se�R*�X�Rw�eFDR���<�+��ʹ���z�o"��ែ�`$'_*`%>k��B�O5t! &T�I�>�惇��c�5h{��9��o�8�x
��������Z-bN-�N�|��<O>�˥��H#n��'1��({83�Ȏ��İ]�4�F�
��W8���!O����P0ͲCL~�g�6v��ZΧ̮#���d��H�9W�s��E�T�齃�)�b�v�1����`	����;��aG_7\!��Ŕh��sƼ(�N�YU��-E��T X֩.����]��[㎇���W\�#C����ؘ:ni4F�C�u�zK�0ǎ8��E���r����r�||���a|T;j��ӭ�����|g1��^��1x�����n��8��,r���"�l��ŭ�j	�;D7�k�v�O�P(oqT���)I'��y�{;�m�`�6M��H�{��(aCcw���B��$�Tޏ*Rą[�#�V
د������{����u�ql����;�o��Á|��ý�=Aí~��lT'h���A5�(q�k��I��}Q[0����n�C�ʹe/��~>����g�]@AC�0����h�~-V/�h�Vw���zs8���E����-�^�Ǣ�`inX�ʁG�9�x??���pė�K��ݳ�v�m�d1�s|ε�hr�l�l�^�'�1�Iz$@����1�LZ����g�������VE�n�־��+"9��V"�w��@��<7�!�OB!�#����A}����~�T'��c�-,�'prus[:4���R��?/��!�%bk�Vl�,:��W�����b )E4n���d�7��5��{�^כp!�^[}�SH4&�N[�/��{lIK6/����b�����59��B�C�Ϭ1�m�S·B;��h���P�ռ����3�f\'b���"�B�a��nN�܂<q��1�`�,�Ӄ@Zz�+�O�}s	�����/�~���Rc�I�C���)/%��N�-��E�l�	Nհ�!8��%�t�K"��k�X�^��+�V����xާ��t��y� ��Yxt8%͸���L�y����w�����t���om�JP�+�Oe�{���hVȸ��DsyE�p�i�]l����w��=x�e�Q�],KoX޾5#�Cr�'��t�A�9�s�������+uH�*:��J�FV�?���� ������+��p�C�,�ٯ���#��.}�N��4�K���[]x�I��j9��-���`X����6��L�|����al�uL����f
= _Qw��4�˼�-���v�,v�֖~狼�e��QS�z��4]���y�C@����&����"�y���0�v�0���Z~F�4ŷlW��^���\G��1��֐�4�OGy�����(֑G8�{��ۗ�S>�N��>lN��+��m�4�n=����sl=�^��äצ�0k�b`�܀��z��j�^��^z���[|G��s�j͂�-���6�t��L���wf�vD8��!��O��8��j}kV���d���O��Ȫ� f�x]1�e�a�V�5\g�.��N��G��Wީ��}�G�ٟ>~�W�p�0�h5��@PXH�R#h�I�İ��n�b���R8�����X�oӟ�>u����OC�E�����~��a��ݠuAy�o�lY�.�L�azV���3�}Uk�y�Q�<q�!\"��sͼ�τ���0h��8��}q��@}y����j�d_:.��1cϯ�ܣN��Q�k]:0NS���y>�dao|�пi�nr�ܤ�b���:Of宩{oTF�ʡÇ� n��Y8�t�m[�^A�m����A7E�����6�gD'Bћ��9x�w5��u�z��U���>#����`<�]���$GoK�	�^ 4��b\Fo�t��5��z������b%��=���i~���	q�oW*����V��t�0݆�i~m��6߃s$�@!�gY�6m�dgO<����,`��l3�]����x��6i�Ӕ=�z���`^,���5.��=��ז@� �]Z�F:��ʋ�5q��&���Iƫ@\:�%�5H{�8��'\mzw��x0����o-���X�ɒ�"Q
�������î�B"����
8QC�>k\���g��� ���L$�{�0_Jnj��JQ �Js~)P���^s��#���wx��a�<w}N9�����m��z �c�H8ȯ7��W��A�^��#z�&Tn�Z^Y�ԯ��������7���δOOh��:l�y�-��G�>5Ð����/��Yd�kK������ֻz:t�0쁺�^o��"�xsb恶vk��������j��r�jW���[�[�w�<[%���^��0�es�U��^R���i�Jxw�����е�1�Zc��)9Vǁ�{�k聭��KοT�6��c����c7J����O�� ��XV[�������Zެ��q�z拭m/�Gq�)����cs�.�>CV�5��J�(��r�=kF�v�X����e��>���B�mg[��hR��N�Qh(�/3a�[޲ $k���u�i<��Lut�֍��_=|�ι�ʁ���@�r�i@������'��ć��7��6!ۼɓ8�����@�d�BՏ:��:���eA/l�Q�9Fp�XZ�E����NG��F2���`0t y������0̲E�&�֯gB<l2�uB:N�T/owߧ �I߇ѓ]��ܩ[%�?�4<��<.AV��7���`3$�e�L4�lE�����fr;Wd���>#���9W��D@�V;�3=���B�/�k�y�0'C�|����Og��-�-c�����m���z`ox��L�/"��{zB!�0�L4��	ƚ�D�� k`3>\4�~�x5)��-�n�A�!����fH^Ǧ���fƴ��♄S^�/���B�&���.�P�ڤ;��uV�쎑��fҽ�5��8��X�/�=�ʩle���B��eȓ�&��=�tmK��^�V�������?tt�~�U�����~��~h>S��2W;R��WA�/�����2���o�S�k7GHC۵ �ut�X]�Ӛ��U�j���	 ����u�Bo�x���<�י�GZ7}[��/5���#��9��7�j�[�U�xk�<'���Z�� >_hX���|�0�K'�_%��z��;�5eH���%�|ԣxs!��
Ǔ�ݕ^�s�#�
��w�,UM�>���c^ݓ;8��}�H@�q��M�:�S0Q��;"���ѽj�m	�Vk�y�OD�Fv�|3B9�;⻍�k�lq��.SC�/�=?� �s�C@�(>f���y0�q�s���ק:e'XĲ.���m��F�
}���s	�_ZAvl{�=:��s��т�1C���uԺ�,��/�;��QtÔ�.�<S�*�\7X1����7:�g���X+�W³3Hz��h�f�t���-���B�N�ENëQi�����5Iw��l�������mCicw�p���L�Y�>�C�u�zKHb���4����0�-Gs����\��M�la�@���=ZY�E&5/�k>1@n? a��k�LKb��-�d�Ͱ��k$�̠�7*����CĘ�t�'�{��ԓ�9�A��+�0���Q���D��<ȶb�W3��/[<G�r9��cl����O��1� ��1�������w�\%��ۿ�rM���8�^���[D�=m��n�.��"�C�M��lc�\��@���ð��g�]�V_.�_f��K[����ꘐ)�
��1e�^�ұ�A�6q�6�$= H�D�MC�O>h�S��<`��\T���	���j5>�Lo�����j��'ʱ���i73M�,9+��^519_���R�'���fq��`�f��R2	�N�g�o-CX��s���uj� #���5��;�5�����ʳ%L���ʥ�hݢW3�a�}�����w��c���RZ]�k�]��6�Rh#'Mz�T��˙b��ˁ"���:UUh�V�J�ZD�
�)
B���y�����}��|?zմ�+��bU�ZfP�a�a�
1�����ח���֟v�L��z��j�>v�+�;P���܎N0��rC�͛OC�/�"���[@��<�.y��ƫ$"���l�P��Z��ͼ�~��C����<o��-�Km�T�ɨZSI�ϖ
���*�\8M��~���hS��jk5����^nW&��nC��u�L�<�: ���"���+�I���S��*�ナ&~������oR�Hx�pq�6!1�:�@B�����>x�Js���4���m�5��p�������;��j������>b�{Н�#�~�},�H���$oQ��E'+<�$�HM�/�_j�N����C����d��T��[?d>�G��|ǳ�~���4��.�]7C�=ј��[H���Y\�n����>��t�_Qh��0��^h��aG�=05��F��U	�(�H)���Ӭ1w���ܟ�t/1mK ���ct={ϹQ�
<�E�xQ|5��.�i��L&��S5)�/f���=�._������3mZ8�'浦M�])�S#=yװڼ�E��nD%Ҩ!z�~=��u����E���7R*��
�=����ή�H2�*��N�Vj��!��:*R�� �l��c��6U����O��|���䭞��{׈��B`���,E"��+��Xm�ޮ�S �54K��d��&P}�콻�]����&��ʎu-
�jtnۖ9��:N�u�����f���".�I��]���]�n~ħذ��g��d9b���,��,{x�ĳy�ݻ���ֿѹS�l�1�u�q�V�w5K�:[XA�ˮ&+NX�������+�":F6�Ż��BU��8��hv*.l�B1ee��.]j7ÜBh�vb��U�JÌV��*î��IqT,�i���=��b���� n��r��j�����Ep��C�l�Cz!�7zZ�{[�&�EN̠v۲m���D���޼F����yz��uo]��s����cnF���ř�)b��}��=�N�04�Son���<3ꏩl��R7V��w���eF����G�p)[{
3T���M�a0\�8�%!���Ҳ��Z���9��P�d
Ҵ<aA����2>��R:�V�a�f������NB���t��o4�ԭ�EQt�9���pm�Y
���)3U�%\R[��+:צ�&��+���*�wE��*�Ǽ�s��3�o;��f����VP8j����I���lP�o�.��`S4+�܎#�;Fb镂��ϒTr�6��X�k0���ʯ{Ssq���֣P���� �s���*�s ��@�pOf��ך��I^�4��
e�u�x�Z��O#E�x0ȴV���;��ޕ�՗��J7~�ͯ
�4�,e��e9�e��ʰ���i�+n�m_^��B���Nr�_L�l#����kMnWSܻR(5��aG�(T�U�r����͂�id��Y����6M���!�ư�Ȑ�0��>�@��{l3r������ӊ0+qR�)��0�CeЮ�t�<�9���1��ˌ\�R�V�$%�8���(Hõ��6�3l���6�A��5س�S���n1~l���%��-��]Y׮ɤ��;���%�_.B�WV4�ݚ��̶�:��O[�����moopA��eK6��z�l3�"Br�7l���E��Zv�Vs$7n�G]fM�<�3�2 n��)�VLo����Œ
9&̪T�Ԧ��8��������f3�t[cȭ��;I`8�1�]lx��Y-*[:Z�ލ�d�n.cj�a�A�w�au��w��(�	�a%�o�(��i��+�[�@h���S�_�E�1��Ѕ�Q&��Αb�V�,�+g3|e娸>��I�u*UΨ�8n�k|�u�
���3��u
��|�U���'��I���v=�̍���LKG[ty���S�u^2C;Bḙ�>`�*�q��ޏ�v[�{dN����`~9�Vc�g*�D07��2����*��q�{�j�ś���UP�@B)���QT%PPST��M-4��=>?_O�������������<fZ
i�������*���bi�i�����+��x���Ǐ�����������ADB4�CMP�HU445{B4�-1��h
ZR"����)i)h����h����hh��"������
K�ZR`()tH���$���)
��b(��Z���������BLi��DC4�4�DUM4��x��uM@Dwh
�J�Z�:����AD�I1ATvƖ-�Ge� ��A���A���(�o��z��%�Q�F\l��'MH���"b	&�-wn��<r�o���'�WG��mseD��B/HС�צE֑j��w4r�[b>k,R�L<6E	��S�%�f�p�IF&dRC�$��P �!h��2��	�X���j��߿	��������+ܑǪ���%���H�CZH?{��4in*���/z���Xw1�e��G�;ƫ�A�G8OP�n� \��x�(A���/Pzg��_����z]����Ѝ�����E�3L(qh��+�ղ�n��5�;9s��]]c��ăVl�H|12������N����ƲG��k�4&��i�֣Tӽt�Ỿ�hY٩�e�;C�~h���!��h�昘I��[e9͏#��^���-�ũ�cݑ�ք��� N2��٥�Y��r���l���$�<!�n��6�_L��D��Ddwt�^�Z��BZ��IQ�g�ٶT2��*I����	�~��/v�ϫ�+.������i�y��wB	���a�@�5⺵��S�g���̶��Q@���������>��?hsʎ|�sқFL.z�D �^��):��P�t��j۔d.�m�f�ahx�mati���p���3Ĉ��t)�5תv��f�}	����'�)��C�.���W��c�aG�o�n��]��D�v_����A� �~i!�e"�Y�k�вL��5�j���S>��Ъ>f�������+lx��R�ta���c��ҫ�`������WVX5�k��ñ=����;���^��S�)Q�v�ڵ�h�"Cj�|�M�٘7�^pNn�� -B���cp>�w�U�)Lam��W��}��y��p��ٍ����W5�^b���R~UƁ�6^��[�	��|ׇ˨F<9d�^2�m����[���+���%�-�k鄞tr�d]g�x`ϸ��}��Z\Ws��C�Q�ۋ{��:��ek�-~�`�5k�A|BpУ~�I�Y��֣�ȼ����`���nC���QN*�����C��v�5��iz��uSƅ�d�⤰�]T�n�k�/�Ru�!ڗj|
��,p�\0g���|���y�Lr`kl�^���d��ұ���8�Ұ�D��z�i�[����|���$��u���3�k�>^���/g��}��wjd���Aʍ�7��.�z!����#���5T�5.�e轆s>2%�=��dD��G�#���'Z��m)혔���5ܜ��P]��W��/^���8��Ya�-���r���8�4F���k�c`�sC���z`���s%�!y��zB!��@A�/tfhv~�r�>?���O0z��������ڄ/�F�K�n8�Fd�{��^=��ƴ�A!���G=r�"k�7N�G��)�?)���V��n��{�u���i%�1sGհ;����82�GjwY�-���D8E;�%m�?�n�ܣ���6)A�\ ��˩6����n
nХ�q]o_|��!�Z��:���af���oa�������n���|�u��z? ���p��8@A�����-R��v=G�>"뇻���zi�ʩlj��!s��A��B�J�� KETO<)�Ų����8u�,�.:kuB�/;�?~br��sҕ�Աnt!5���>zǚ�6�S_����G�MkGp����W�h��K��\OW�,T������sv���w����}2��>�/�L�	�IT.��x�m�z��Yĳ�Y���X�S=�[zW]5����|b�(�� dޚ��L���"K	NŲ���
}����'�^���2:5�+G��&b�F�%�_C�t�zג���H�,��������\�����At5vM��9�{i�f�\3sO��suz`&�ƅ�I�U*��E�沠��9!���٪�l1U��5�Ӹiܲ�]�j����y�kO��ct<JL�Մ���Q��p+睶k�18{i�Wv���@eׂ祌Oܼicm��=#������i��d��H�9vhDXh}�r������l�I��X*	|���u԰�:-����3Ǭ�?�n>2f��=��
���u��9к3u=��"�n4�6F���~�h���r�=y��@�Ӫ��*��ul/�r�@��û���_�d�WK��8q�2�Ҕ��-������*<H����e��1�LD��f�p��,@�������m����}���?�{�xe�blp�ɚ�dSg�M&7��:�/��q�~c�Ǟ�;q�3?��'-]O��vs.�9R�z��x$mݢ�K�v���ق�Q>���/@ vqy�{�DS���L;�v�D�l��'D_v��[}��#��K�X��ҿwPn��X�D�s��$F�MC]�7�%�f�}-
/��}��,��>vb1�d=�O^����y�5�7:���d�I������6���;����AAy/��ZgK*������ǔ�ٹ�C���Ę��Fο�wS�����_���҃*d����z͛OC��WH�x[Xd^�\/0�o�[])Y9EܞΦ�7����J���%6r�1���ڮ�`y���[�z��U"%�U[�͝[��B 9������74z�e[(�%�{\��_�Mv":���;�h6{�@��E����Ӌ׳��k�$�6И,�����3|���Г蘉Nlj�Lhi5���86���Y����q*�������-�*Y��,��v
��q�&Rr�)��*��bg���W���_�(k(3"�/��D��A��Ά6����������MF��eh:�#��oj�&Ic�J;�m�ԉ{�ם�nvfJ��6\��HeӶ;v�����-f<;���z�c����Y�Ծ������}�/��{���{�8�����xx{�L�`�E��nhe��966�D�\O8@��UZ�5b��|�>̼zm� �z�	�����7��"(��R�}&��Q�	�:�x�=�ܹ��.PP	r5���a> r�>p0����k��ֹ�����q���}�j���ƫ�<�H�0��w8X�;LK�k�;
Y�������ȗ�^\�7.ѦS�^�Ȕ�BT�n��k��%?5�2m��)��^�H��A���W�uT��c5w�9�C(a���vO������7���$����Z��O�l�sH���o�?��j�@}�Uwn���#-~мS�>>3�}l/^�d�>�4#hgRN�Fi�{ËG�fz�6DX��s3D#�w��[,}����C�*jԐ3�5��q������dc�Fv�3��wZ�N��&�S������f֟1��|tE��sͼdK�#4[�?8�?�?5G"��9��I���p�T��l#���Vl�C��;W��d�&3-a�~�ߕbP�*�7������1�i)`jv'�`;O�KZ���ϫ,v�_5Ь8�BZ�Y$5gY�f�?V1e|��Iz-��y�b��ź߲�J�v��6s��5��#�@sOp��nS���PQ��I��f��*gv깮��q�=�~�H6P�1�a� �����x��"�ʒ	�XA8Izma,�	�:��K��]^J�K�˼Բr���l���~E���Z�l/]��?:���|�r�w�DO���p(z�ޝdD�Ѩo���"1�D܄�^m�9��� ��YX�\k=o�O.$𒉗��9o�{_5�:��P���l�X�N2;a���&��\���2׿r�N�-T)�UDe�tvb�ص'DG�	_���[��o��j���_���"�a'i��nЛ�}�	�|��S����Q׮���K��"�TS��ٶ��WE��XQ����Ҷ����8<�[Ng2,wwl�ϸ�/v�Qe��X��E�����A�N͔��� G�ivv!?mJ�ݹ�훜(��u�0%��|i�@��-��|��Xxؾ��Wu=O�'��Ƕ�R�b�M&U��E���@C�b^����Oo&Ves�Z�E璒ƽ�i�O�xw�D��wMG�60.�b��c�����@���/:��fÖ��qvE���e2��+v˷��_[MNB8�l�k�E��V�c ��|}_�$>>4���8���"�r�q�ǥk����&���?>o�»���P���l<	�@`�#�����4���Ƅ�2����zY��w?=��7w#M���^;��ڏ���r�U�*��k]lWu�OV��
�|Z��UizN�h�i#Z�*��c��+ꕈ�3�K�3.��`%�{7��^�l.�����z<r7t)S����\�e�y�����\�/{�}��|.@\�**>�|�;��t�v�����c�(v��ƥ��8�-V
��$�p�	��$O���}���&X;OW+3��rf����f�ίe�<LIza۵�q��:��@�r�6=!M�0���e���]�.A��+�^��}a^Qm��ݦa�e��C�@A��iD[*�D���~�S"	�U�����ʅ@���'��OsQx��3cZ}xބ��U��E\�("k�YV�csS��,�o6�7�տ65M^(U��>����Af9K����U-��@Z�ve�m�s�`U�Ͼ��ޮ��N���	��]�*�Ȃ	mI�lS<!	���i�9�lc%~��nl�g��WZ_v{q�xb�HL�)�N� ��4��X��v@���8���"k����/4��R�^���KWA�X/��JS��B�ѳr������Hql�V���V�:_23��\��0Ǜ���*��L��<^%�u��)�^��]r鿒���S��9ו�r��ݴy���c"!0����n�|$J��.�}]0�U(��4��@cU�4�KA�s����o����T���ÿ�H1�bF���Xb:°T��qf�d�b��U�1�x�5�2{��y���L��P�X�4�_'��v#mT�6��y[��%ѻ���)�+`+�k[�&�vju�񵳘��uq(��z�In�(���sͽ��u�u�\�\ ��D���I(EOZ�{o��[ý4x��lgp�ݞ�	��Ȟц���*z�E��ǹJ{�6c��]�y�:��cjvu�1a������B�鏃�����N�#ư��o!F�T�Ԍ����w���s8n9N�^�.eT���9��8x����:��A}��g>���g6�Q���V�Bkl�nb�mc=�PKܽ��tG�N��B�9��x{��e��|�B�WtR#zs�(vn����6�qʓg�S4�c��q��1Ɇc����y��W?.�*E�+6s��,:a��ߥ۟f�C��,k	E��s�	P��DS�v����ޟjźw'����'hY�E�	A�8�D��{��t����ٵ�!����"���q�qC-l��n��J~���k"Y�p���yC ��=���/V�lf�֐3s��Rô����_%:�I���@k^9�4P�0��^/V;׹��u�,G4��&�FFS�j}<����|v=z�����d+��6��HY8�5x��6)>�ռ*���[E�E��䃓�T�;>ϖ*����悈��:o�.n�6�w�x���mjL�m���I�ay�(�yּ)��N��RW\�)o΁��%�1oPφ[ӛF쒖�L]>f*7J3�B�hlJa'_
�U�7۔�g�m�>o�0�`���:�bq��H����>���=��8���<N�Mq3D��|�n�O���5*;��/����sW�دN�%6X�(2j���j0+��	�ǫz���-����Ɓ�:n�S�M^�U�P��%�O��~��HC�6U��8��%�y�Ji��F�]����l��p�Tv!Ѣ�������j�~D�G�~?U���gB^��N�ሔ�T	c5M�KCTP�;X��1we)nd#�y�ϑp�^���"�)f�M��}�g���O;���ަ���j:�h�u����@1�F�Qa̋�Qѱ��h�a�"m	��m����Q|�Z�4ɨ��Y�B�L���;k���9�=��,��2�K׵��İ�@~o[;��`l0Q��GW�T��+)��ܣ�K��q��t'��e�	�k�R/jF����w=y�3����61��y��?P��P�)b�B����D�작M�wU��ޔ����{�v�W���6�;H��'�W{��}y�Z7��C<��`r�C$�!ع/B]��E�j�Ia��5��=���e2��������3{��y��!݊�΃�x�����a|�����4#k:�plFi��z�����TÌ)�� ���K����
�WX�4^���/:�3��N�[�XLk͂������gR[_j����i�Ɠ��2>�2fri&GiUA�sXf�+]��_��Z��'gg��1���5:~��o�3�p���^�z�Ͽx}�~9�a�]]���\-||h$/� �����(-10���d�v�k�J0 k��8��f����BQٮv�#~�b�1p�N����y��[�����h.9�'@H�WS���f:�+�����.)g��O�זhMoJ�j	N05{���o�i�sͼ���	K���c��u6o3�a�[#�ؚ��+v��v�8��<^Ĥ�kYFy��t�*��/�y�a�i�{�G1�>��n����!s�f<��D܂rg��˜��d�,'�d�bWN3�f�����ef�w��UoMr�`�<9���9�2�����M?�����2��r�N�__�U��Ll�S�ks�P�@Og�U�Q��su;k�;�]��������@��n/��4�ü�iJ�����E��]㟸�L��f�H�hU�oG�Ƙt����-h�v�1�������m�~�f!�,�m�R�p/1W�"��+��_]��H܁!�o�t�h�az{WMf�p���R%�o\�R���}0S��d]^�k��8���<�w�eXy	���&�k��v]ٯڴ��=�l�(���&���q�w;��_�^�阷�]��-�wj�;&�qr�"��܅.�ռ�q
�u����LS�M�'Zz����h���O'wg0K�bo�z'|�����u�����:U�SM*1!�$�5���{�6A�74�^M�ם*�r��Kx����|�3��'��N��ԁ��)�
hu\����ڍ�����`�F_km�Hc���zޞC��\�Uke�G;�0�6��5:m
	�PD��(���F}c�V��%XUR��U�_N7�N��{��:�SY�\��ZYr���f�SK�rm���X�[sy���y�	R��T�����dL��ݾ�6G�
�$C\0t\*�#�b�o�.�Xj貫O�p���
a;�vC}�|�;�ٴ�d˥5�I�-���g.�&Nm��M�*B+2o�G���8���y�-k%0䣳���8%Ж��+r_RS�ᓑƝ�K�:���ffQn4���{ئS*u��5э<xTز��`|�_>�Y-p��M����ٛQ�g7�3��j,�9���}qx���fk�����I.��m������t�yȓ�}�h��A��J[y��#���սN������ݗ��U��A󪇂��C��˶�FRCt�t�j��#��3����ԌѬ�I���xo���3�*y�7^n����J&�4�ym�ҷ�JVE�l]�Ht���P�CMfccjڵ;\�3�f�fG�k�a6�?��C(!��Dv�1]NC�lM�D�ee:jP��������75�roVE*]�v3q��T��.ͷ�|�]�Ҭ�����48ɐ��6G5W����z���&X����t݆e�Yfa��m��]�W��U��ě>Ӵ��	�c,�v�#�M��,�+���WNN���������}o"����@��t'jzXոN��ne`w�ovU�|����(�z�e�4�IR�L5�
��l��Gp{������4ػ�X�Xx`s*إtb4f{�vmJw�{��Ҳ�#���7_�������Zȝ�җ|8���ƊMon�Vz���9�5ֻ뇒�/$ۥ9f�ZA�l����c�p�;f��&�jï�
��M���f�E��p\y׸vhԝ�C��@�.�%����v��Vr�q[�u�8�y���v��=�u�����hk�����n�=}����:��:<뇹�(#-1�^m�NR�c��� p.9���E�ı>���������cY��CO��u���J��;x�3u���CE���ዝ0ps"������<m�����)96����Õ]Gn:�4/��1e�**���4q�t�GJ��U@Y�}�#-n�M(�e��4��b=��w�%+ѷ��{��߯_���>ED�CE	�4^�IT�۹�T�ϧ����������������y4�}�U3AAAIQ4?%�DPGNg<x�x������������x��

��J=A��
�	�
��������|Í�%�Q��2R���(�&("��i�1��i�:�U��z#MUMM��QICQEP�U�h�����!(���MUT�A�Jh�H��"��j-�KSHSZ5QDTD�%U4TTRRTTQ�1�4�ݦ�V��G]����i�d�����Ӡ*����(()Ji1�~�������sD[��_�l����5�ɘ��W�E������\��ߖ*���D
����a�ter���Uz{�x���?����3x ���JUsN�%�2���6�a�`
z��~�2$ٔ�M�\��j����в]�bv���e��w]���)0������t��^5�	�B͹��.�E���c9�Nq�3��Mϳ����ϴ�����C����A��r$>*��C���CM������!�6�nU7pyW�t�toc��,�@�J��S�'�bi�V���!�>�Ѐ��ИfX%��4[�*_Q]�^�{�|��e�Z��k��E����,��Ɂ�[02"tBa�T�Jw��:-,b#�V?�-T3v��� 3l�e	sʇy�ڻͳ�
��sW��X��_Ul�=,���:XE�C�sD=���ݦa�,��@$���Pi�z���-���4Iγ�\+qZ�xiW���J�Uύ+�_���a�{5yh~�����#���ccj|�r��q7;�����B����X~|]��9�O��a}�
!�����.�Ztw��Vq��F��0���v���w"qƏ8z���	׫]���p�k��g�����=���u{PݔaϯW|g�3���n�2u������^�(��<�j.��鑼[{o/��o{�5��Q�i4���V�^ф�=�F��aO"u�I��Ϭ�;�J���`�]BEz4�������7��8b�=��.k�ON_����T�we>k�+��}�|~?�{�f��aY���[~x�	-���&�X�R{U��c0#;�X�oMl�z<��C��*�9
�w�f_��ws�~�B&���Y2Z�A�xNx%)�e`�o9O��/�(�܇e���Fn�MSBN�8gA�K��08s������^�oL��<^%�u�s�1�Q�F�s�2�۲��i�Vs:Qh��J5��-3d�s�@K��>�%U���p0���9T��剗j�Ȫh�]��#�rK�^��\i u0��y��~y����1��ƅ1�P⺊��n��9��9��5غuۮ�Vs�.�Lhj���A<y�N�}�?��_0>OP�y}S���ܟ�tq�{lZ/��7:���h�ը�s6��s�q;/N7 8�#Xt�������2⣩.��k����֦�	V0�]+^�PKܽ�)�U0�����3��o3��ۏ:����ɧ[-�h[n��Zaٲ�EgM�~R��Q��c��q�sI�T�FvZޠ��ʢV �vv�O0�������#�o�Y����01�/��(�\m$n:��m�,��+u_{��z�E���X��V�9���N����'�鱳�|^��L��ޖ+���;^F�ތsio�1b"hc�H^�I�C"Fm���E��:3���V�������%Y�aw���gZdQ�JS{�Q�ڇ��ww�y�_o�Ȇs����Û��N�w�T���1h���U�4�����[�+�d(�x9a h|.�,+����@���3;�������*d����qB?j[u�����l��%�<D���A`���D�[��C[o\���g��?N]�C"��~�̈��$�ǹ�A|/%��R�0j�X\Y�|�,Z��٦�W�^��7ڊ�˿>�����ב�i�qTͶvP�+c&����3�x\7�򧞻WF��T����l~�\����<��!;�ɜa�1�ݼ����MiD��]8��վ[ռ���	��L3�oMP;���k�l�H�"Xc����~�X�UmC�N+ܢY���+U>,��ڌ���j΋�\���g-N����(�I���d�|��?#�Ԗ
�p�Dٓ�])�|"S��60����ޘ@|�a���}��㹙8���ۜ��ȳ釯t0�K�m BRͰ�g���+�.㥚h�Pu;̹7�����ÆoF��C�(�X�"�U̘����}�O���G#��Bm�1���9Ψ�53�D�ڼ����[Qu�]�Y�Jbj�v�HO �֢�:�M0����`0Q���ye���[Dݫ��l��y���<��
�׹�$�U��OK)�Ɩ�.n�gM:��-q�bC��[��.��yh����6��Ư2�ۼ(����V�6�t���C[{!yL��R���Y�ۡ�dɛ��׾��{?(�?� �8A�E=s�|�v+]b�.>��ާ�i����Z�a�^;ؤsL?���3�/އ��ve�:}�3
U���P�(C ��!�>���']W��SW��=׍v3�'�-2m��O��dw��:�����hڜ�x[I{)_c �����@]�ߪ3��UՒ��-X1%�S�Z�9t�l4����ó�V0e�׾g�Ya~���~��B
��rŜ����ȭ4#(gW������ycW��hi���s���+����^V�)��/���?�z��1���d+ki���
�wN\Wg ���H��h�W�2�X��q�DYz�o�D�����|�K��06��,�-۬0���\�^͟FR���+���G��L�M�����o�E;�u��Ӯ��J��h�(��a�-�<MG��[t���b�\�
3��3f�v�c�,�z���ѳ>�V�1/�p�2``o�5���r�񼨬j]'�va�j��͏�X�\�X32}�5�_wb���}>V���l���.Xs�e~�G�z~:2?�P�k��+	M�=��f�lju�hjk�N�]�&��X��	o�6��;Xw�󻦲S�u [�o��ۑ�f�oL��x�ЪOVք�ܧ��>��������-�]+;m�cݖ­�1p���)��ʒr^�[k#�7�����>�>���?��<�QZ�V����G���*����PꋇT.1�C��(2.�0|������:�馛x��eM�퓝]���1�=��No�*��N+��X;�}ހ^�@�H8�+%�M����B�I��1yG(�f��/L�N�L�����E�WO�b:l�;�0���T���f�����}������}�	����e��4�1|�S͎Sl���9�o<�;�����O^����߼���Ax�3���_����
Ŭ�X¨Y��B��/6���DTm���X]̔C�kv�'`���@�5����ѱ��*�j��z���/I��IaH�B���ح�_v���B��#�qi�V�z��t���C��憛�N������{�/�g"�S���=7�����Γ��
�_¨��'Z�=�~��p3@#c:�S��� i� ��9�ͷ�;9�v��Qaͅ)-��@#ӕ�5-�@�/@��s>2%�8��R^-p,(���pӿhZ�<E뫓�pK��n�a�L(������_�l���B���9M��r�g��z9>��f���m��˲5=vh�)���Ƭ�)�x�2k�;��q�W���*FN����x��=�śF*��*�`{G���G����J�{Fz��m��s�7����ڽذ���ю�j��6��0n�\�/0�����s������
- �����޸o���?��,T	�h�_<�y��ME�7��fy^k��	S�|�L2�u��C6��UWd1�u�7!�6��C���МEx��p����p��׶�����H<��#��`<6�nz��K���g�xf�0*���[�\y�k��E?��v�!���=I��C Q٨����d����vWg!��\�(�B��Up�7��M�S^�le?��5�?��Dy]�>
[.�s��6R�̱������)����a�I�*�g�����o"���1l�B��Ω�����[й|S ����{�W���P�BS+�x������MAIT.�l�>���w�Ev�M}��xu�hq��\+��y��|k��	:�&Y�ƼQ���1��k�#j���J��mD���/P�fɈ,=K��7�D����>��.�r�E��]#��G-���v�6-ݧeAGS��0�65y�mi�#��`&����9�)�K��J-恼ye��׽ܲ r,��q�*P]���8�xXl��lD�ߏ�i�zz�G<��f����͝��r�]�l��ֿn�m��T�挛P.��$+B�.qg2_5����ŷ���z�fg>�p�J����Ո�әԌ��fʼ����0=1����g]���־��K{����0�j�-.�h4��nomV��AV�9�:wן�����G9��R=��y���z4��_q����;�\˰�$���"��1^P��%Q����d������^�<n@p��7���G�UE3���,΢�o@[NW�%�W��z�[Mk=��z�B�sO�Գmt[�!�Lv�7�a��dU9�׳^��]ٓ�X�f�-泦�_��&6(�|��}��;0�a>^�����������A�����2��A���59o��~[���������HH;wn�,��}SoX�v��ȧ��ՁY�T=����!����*l��{�K�Cu��m���F�\E��a2�{=Q׽�\�ՑG0�_E�y����L���~0����5g�2��.w�x�P�v-����W���ޖi^9:ëﲇ����K�*����
v���t� ��-��c�9O�Gi�zj}8��m�G0N��l����	���S��Z;��h�4��O�get��'#�D�hB�h}ǐ"�ӕ�U��mEz}�D���(2j���ڮ�a^=�'+[6���U|l�ڳ���џv'߹r@?���%��@D:�En�q\�u�|
��'g25sK�j�"6#7��̈́�Y��o�xs�{�S.V���Z�{k�����Wgj�b^p#{��E
������@�U�WFoJ<�l�|;�5�I-]�#slM��s}���X�`C�g0�[Vvmj�ڶ��+64%�H\�����~P=��
g8E��y���#vR������E=�Ǥ(�9����!0Q|$}�"S��i���e������:��w��r�l�n��4���m�5ȳ�~1�	�c��m���̳.�a�5�j�=ӯ=���s��הE+t�5��lÚ�	�/O���h���r!W�sE'�wء�Fwq���P�)y�6�ʡ��&�~OI��	z�Z|9v�i����!�}��c\�?C�<R���g�?p��B0��U�ޚn�g*ֻe��#X�ג����I�wg�4��D	�j�z8wm'g`�,vn~92']Q�B���x�TZ}b�ɷ��)�Zx\�i\d��3��f0yCu�ݘ�t0d�J�ݛ]�.��zdR�Ia����VU��K^Z!�Gfp���]�β�a��D��0ƀ� ��\|Q�~]�a��za�/����D�w6����{��A��0��;(w�q��\-xו��T��E�PZbac��<�j�mK,����Y\�<���6��;	�]��f->&:I�_�)��D��A�5 ������Q��Z(�.N�o VL8� �S�0��P�1'��V+��:|�b#��߽e�H3C��߹w��Q���^�����6�l�.�rQuZ*7$j����ot��0oՃF�0j�_e�Y�2Ko�&�9y�nT #�:�Z9(~�����~yǇ��� xш�? ��k�-�_!�_�fϠ^Y�5�'���dQ3>�ƴ�<���|�}����_����N�X�:!0�=Ŷ�������j�H8�0���Hj(γ��{Pb���g2��7�e,n^�ϯ sӼX�#(`��	��zaQ7 ���l����]�k��\&�1"�c+�B=zjٙ�l�#o�����3:
�x.3#��������K2���:#G'G>�;�����]�K�y/�:D���
j[s�C�.U�3���
�������B��-�IZcr'�S7bۙxtAd��D�6J��
��q�l'�-�WN7��ck�Ͳ��I{_R;����>k�n
�N�?^�v����M8^b�sȢ�\���g��'f�xa�5�(�UY��%1������4Ai��C���#�o��������E�IO7�m�xX Ďj��m�y@�U9��إ{�"���۳{t��`u�C���@K�~�2$ٔ�O��熯Z�E�]�t�sŉc��"�Di�孨fm;	�i7�Xv~!x�l|{ʢ��}�+�������p��-]y-qr��{�\�ICk��u�6��moZ�t��O&�h�ih��|�N�=&L�T�>�%;8�@���;ꋬ���
�JgA��0�;�J��o;w:z�]�õ�=	3kY���t�N[�k&�博�ս,w	�������~��� f�Է��J;;�c���X��R�`�����ώ=�11�k�q��gH�¦��n���5��13��S��`���Ts	[bu�{�>�3���3�Q̣)p�1�M��9�7���Ѫ�2{ ��4�w�P7�KƯ_f��ƥ��ǠYz}"^!��?)�]sv �>��gL���B�[m͉�mN�vY�@��,(9�_���C�#3��BO�S��W�U����k�����<���`L���ZFN�ޱ7l�&;���^��{�2N�efb�w&V7
=�JW��x��9��`P&|�Yq1�ݤ�&�5�:5��-#�S�B2�S��Sv	�}�뵸
��_���x�~4�/�����:+�,/�B ��y8����s4ۗF]��~���%� �����\�;���su�Є��0L�!�5'��*61wK��B��6j�-��D&���ʂ�B��
�h]�ǹ�����Q���~2Lt�������b�C\O>��O���5�nt!1@�JsiJ`����]��� �&Ye4��v�\��f#���-B��~aG�7z�v	J:����(][�]Z�V1�R��y��r2�$�2�njc�C�졚�Gw�d�k�&�5�>���=�װ��Eq��eS�{c�P�{y���ƽ�	�2��fYoN��w���-�;+�.cҹ���ñˋ4���/w�|Җy��ظJ��d��c�mk�[@�^h�����@m�ܘ]_SkpU�4{�#�����k77�R̫h��	�Oܩ)�����#�������2|�kg;w��2���̌j��ܴ�9M���t��ݓ�O�%�=*,U���7��nN7��{7��ێ@�]���w6�bW �<z+N��䇖c���7�L�vX;�oI�yB�sCr�n��A6����'�k��݆f��Z��:'��Hܩ�rk6��,��k�[UA�R7�U�Uk�f�.gL�.����&����&����U䑎�kT�Ga�њ�7��f vE1���ng`�I;h]5��N�.��$JL�s,�xx�ܒ��I6���[�]:�9��n���t(��9n�W��T�����/l!{Xq�%N�Xj���͗�����r�N�*[C��l�jK�C2��.#�����������)��^�z��`a��gmn����uؙina�۾}o�lo:���:*��B;[��kdP7�S�s"Û�Ya����﵋�����Z�����T���t��pu��\A��l��pcᛳ�DՅTs\��L���$q���\�_kil�ՕQ��R2�Mq8��`���Z,�hr��e��֣���d�W�ο[�dc��aD��[�;^t�}�Q�Sg`�8��V̮�������w"u��UҺ��n�]3�vuohh���D�����Y����ő�U���Z����}̲���^TU����.�1s�`��@r��d���gR��8���.[�������ϊ��k�/j�,X�[}��?66����$n���J��S��
��j,&N�J��én#�2�pɘ��'2��
'zԈ��}�7����uy�DV^��a{���4�uU�ەYD�&��1x;�U�j�=c)#2���ӷ��r�9���2�QFQ=3���l�)��c��T�n�9�/:b�8��z�p��Y*�uV���V�َ���au��Z�λ�6S�x�	#u���(+�sǺ��7%���}D�Ŝ1اu�Vv�,��D뙜���Yrn�q������I<�1pc�h�-^Ri<����t޸�ʃwUե��<�	������r��N�Vm�H/'��1�<�m��F�ں���3s�����m\����P�Ar�Y�Ć�[�c<؝��V�u.��|qQo`�U>�w��%WnƯ|����R*�p]d�(��OV"��$�X"*���JH��������������||||||~����j**a��)
�"�h(�ڪJӡ�;fs����Ǐ�����������r(~�#K��k:k��*(� ���@LEE-5U�3D�؋C���STѤ�S����
4ik�:�Mw4����*gy.��j{����	�@�(*���MT�ErG����1u-4:4Ę��M!�G���Lu�)h
oXu��PbLl����V�:]����"�kM �4h������[�0[[��ѷ]�CCK��N��:��M:T��(����V5��:��UmE%SJn�բ�D��E�QB���&2Y�C���"�sQ�ڶ���$"�}�l�([4u��E8��m� �Hx3�v�5�����9|�[�)��V-(�-8I���&B��3��P�i��f&Q"��_���/�����f�"h��m�hǋ�d�+�RI�P^�'m�hⱪ�k7�����7��^P|�0O>��3�ޙI�g�E��c\0���k�8V��ܥ,�b�u_�ՃU9���}ʢ�=/����0��]0d�8���Y�l�*��Y����]��S��n/���6�;�@AC64�8Bn�0u�	8��X���s�M���Omv"�%4a�֢��X	Ac��7'�����M��8F�Hl�-��ZeUYk���S��Sl5�ye�qT`��Τ�����1ip���B�T�ء#f
P!���j/��������ίN�kd�Ͱ㰱�O�W�ό���9�������?J1eV��2��;�s�h�f�y�gM���I��Q��ޱ�=8�8�5WV!�<M�Ż���u�3�jC"�;)�΂���Cξ�vO�/$;d��Q~���"�6�cvj�Vmݮ/Bh^E���~=A#��q&>�����!J�/`K�:]���^�DVa���|���XC/_A����D�j|_E������
�/~�u�?|��Ziu�<��.�DxѸ�1Ր"�7�\=>#+����T���]WH�FS*y�iþ~�yL�=f��PdQЌ^��& JBf	�VuFUY��mBH��t[��A��QW
����gs�մ�Ǆ�|si٤b�7s����C߼<<"����~��v��<j*ٹ��;��,:��PB���p��[�6����ޡa����3��w���12�w��H�����S��(�	�Ɲ䩛l�ƖN0M@�m����Ui��l����wY�����]�d6]�ƴpt^b���j��W����)��JZ�*�{Uӌ.g���7GѬIL&�[����h�"W���xan���h�d�殈A8�r�d]]�%��D\Ef7-���%�{�h�؈�Xk���)ZLA�2��'����A�7���X��;m�HiES�����n�R�n�ˉb���}B�ߊU�mq�<�"��?���	K6��Z����5ܖ�����9���z�$�/M���n�Pc^��sP&,�y�<��W�B=��m]����[�� �j6O��j/c
�i�~��/c�Zsɠ���.�a'�?D�p�ٹӦY�ZgA��ba�Y�p����;�M�3�k]�2��R5�=%�౜q�o2u1/�'��*.��E��?�0y��Zܨ4|�͇��7P�궻ғ�Z�&ާ���1<ᱮ�-�"bB(e�������u�]��i@%����A��$�4��1g�r�nFvT�@��ֲ���}��r_S깾�{Z���a�\� �����\
��r5*\�������V�<KJ+w#6����.�P�~���޺���wWd@c�3nA/N�ȻA������Зm|�2)i�,:��F�y�!?,l�E�������|_l<y����:�>8֜��#���Ԭꘇ��'�����B
�����#4Ë_�'9��Z<|8�߼x/�n����5h(,�Y��-�2�5��#�V[ژڨn�my�@�<bK��,Ť$�w�C���C`�M{��8�Oj���b$�~~1�M{W�#���c6~w��'s�#�Ώ��r�٣f��雁��$��W�F��V��V��%�N�4l	�!��["�髟WXݭi[	],�Hi�
�
��h�ǋɵ�Q��&�������cW(9RN��d�$s"×�yQX˜���V��G�������s�ڴr���v�gyV_���(V\mz�&��@��Dz���2g�8�B�/YiF���Ѽ�Qn�Au�Rt�H�@UE�5x-�ơ<��p�1�="zi���v;��շW�38�n����ۺ�+��殈,�ߌD�%)�UE8��l'ݑm
�N7���ҝ���1n�V����Iv`;�$���;Kr7'm�k�5t#�+N����ub��S�� �
�)+25c�V6r��sD�U������I�Z�3#��oF�@ml�6�<u��5W`�Z&WK�|�[Z;@��;��E������xxU|r����W@C��6�l� ��ޗiԩ2��c�Ew�:� ���o���0�ۍJ��kE����L!Q�����/���ޤ`��;�l���9�j�z$�5I����{.�@L#�~V��r�e��w��T�:�	y/��F�L*�.xm�wy��m�[+:xGU���yC:S�;P�3��܇�`���M��6�2�On�VP뺑E����F�R��,(Z��3b�k	�=���]
����J����7�?;8���}�WO]��!s�Ebs'p=��zdG0��'Z���`���X�3NW8R��!��8��6��h�mg���z�0͹7�XkPΟ%`������r�Է5�e�Pg%�n�KQ���|�b�:�	���s`L3�e�g��E�_��v?�g���gb���@������`���-�V��x��&�&�#>ZF:v{�7h�x�^s�A!�f8��efxYۨXk��d:=�m����q�{`'x��g�"�1��qU�;����:�|���Hg��]�#P�AX�t�!��J�����Z[�u��, *��$�]�3r��\ü�lS�jb���lwK�L�]S�=T3�d+�,�ۜ�Ӿ#3wM%6G�4~�\�+U���;�/�:wz�d^U��y��iX����3/L��_j����v�*bd�����{c���ܛ�!
^k}�M��.W�)�=�����4_ؓ��Ffu�����=�h��[f���@�W�e
%I��ýs�^�M�[^U�ʼՏ
����e"�}����Os�-�^�BSe�R*
OaWm��ס�V��9>v�M�(��2�2��Y���K�	�xM�x���<�:�ȳ�s�JSԤ���l��5�\j�u y��O؏�{M�L�lS���cP8�q�oW�b	s��Ks	�/%��kc��:;۫[P��,)�+�S���k�@�a�'�	��.Cu��
�K��Fs.�xJ�.�;�u�ڝ|`�ݩ�޻��_�����R���ߒ�C�L�1���uγ��ܙwVz;��8^Gv�I�w��]B�Z~d��:���Rq/>���G�:nm|u[�a)��mZݒ�/LJ|�&K�MȮ*zZ��3a]�X�KӇ�n@<�#q䧴� ��^^l1�	�Z2=ϝ�k��Ķ�N�kdL[k�K_(��/)��]K6�߯1g�axJ_�����&l����9�����7:E��ݦ=�4\�kZ{��Ժ�	|�j#�da_��ББ5U�J�;�0�K��Z��N�bE�Ѵ�n,�;�4LŰcV��(y�|�r����#�7Գ��ͫ�����މȦG[�^T~x(Q�	`��.x��L�Ͷ�ˣ�&6�:�/��q�v�(n�i��Xq���c�_��&���A���0J��O��� ^�3�G��rE���6�$i9|��=Q�{���z����u�~��Gƀ�Nq'�_�������6��/x��{�TR����{��A�����B!��I�b�)�cw��^�S�=0����ws��zE���~խ2�^��߆�n*f��é,��dÇ�y6����}�,�Of3-B{^�V�u���V���ы�S���Jz��:R�m�vPcAd��
;A�b�����)��(ۭCg:�S�!�)�<C�<��EG���0K�ڊ��x�M�9J��)��'�����v�ˮ�95���Y��Q���6��<�Lq�$<�� ��<��A8���ENYh�7١b���[����=%�Du�5{�gO>��x�`bx.͐��/��:91nah,�J��ogWj6���]x�JscT�c@h�>6Gd�mz���#����JZ���H�45uC��SMU]�}�&��s4T�B|�t�Pfu[�g�WΧ��ҽoj�Z���(^]X;�X��[!(FY�����Q�in��4�jQ˕.�Mǳ���w�c�	^��$h�w��g*ot�Z���4����E��}�~^o0sf�T^Q���2�2E�q#GQ����r�t�4*��LYz���u4c
�50L�y3{mj���3W`���[P���"�y�=�R��W��n��Qi���	}��t�ɚM*9�Vk���>
�-#~#��B�g�U7�7_��ny��"�mH�0�?s����gG-Í��8�Ļ�{`����ǁ�02U�=�-Ѭ��c)!roW9�]�TQx�Lц�v�����0�Ud�<:�Fj����A^����_yW莬����|B����z�Z���\OE֢�?
��xO�>��ݕ�z�5�C��1�>K�av�EsS~Ʌ:�z�3A�����mgQN���a\Ze1\�_��j/a�G�G����#��O�J���8b�sÅ�eϖ$ܫ6���a�:8�j&Y��0�/C�m��rm��L�$�庅��`솅�&;�\ŶS�l�����ʑv�Sl�PD�2�e��'�B�7=�or��\↾u�6���ѡo�V�x��X6��c蚹�ݭia ⅘� ��B���f0�I��Ϥ)	��H@W�^�᤮��7 p�!�̗7O]�g[���Q���Wo�g^��+;��nR��:�ƫ).V�Ř�N�6.�FY����RC��f�z�7�	w��Ϩ��!�b�7�;�.�I�7��뤓6�ϼ}@�����^B� �V�����Pǂ&WƤ���"B��\��/8�M`w��hH��r��I����F�2a�j�+����[�Pʋ�5�`�'�����4��^��u~����ŏ�/���8��Lg=tA��ܡ2��P�j��SQۜj�.r^�o��9on��lMW�q]�rem�B��ݕ�Л�z!2Of"S�)PT��N.�6�}�Ӈ�H�g���c�>Q���n�:��Dz9��!�2�],���oB�Ǚ�n(s�kw��Ь�7,�U�Py��WN�QV��DcH�)���/�K*�4�7�%=��S"ꌨ�=������_�[/^S�Tvk���kÇ���e�*_�.z��c"�P�xi0���Y����\Z�w�xde�/iAcK�C		����o������d��ާ1϶�'��U_tp����YyT�8�*K���f�WZ�|��ۛE�E�y��`�+	��-#n	��o�n�=�o�g�|��Z�P�nd�=��^�¨��ĺ�W��h�(j��d+ߕ��5�Uj��EWVI&�n.�}�9!��!��e�\�.3�.��^��&��zK(�u����fd��p��HU�w���SS�6нy��Qf8Ox�[�A�G�(��S��Ƀ�+.�X_X�Р<��X{�/�����
߶�i�ua�u���j�x��p�Ƒ�<ómȬ���g%@�.�ǿ#r����,�(t��l�=Q��m<�T��3`���s��e�\�2O9��v���
�1%���c�9����A]��Gv@�t�n��l��]�.�4F�C�{aB*-�ݿS��rb�3(��Wp��<�XZf:���\�!��4�� ��k�<7W�3�d!\O��'��x��,���)�J__��h�՜4�a�Y���^��PDךE�\&�f2�*�X~!��e�J}�*��_ea�x�k��-�B���BifP5��(�
��C��P�E-���t�X��5F�Y5�l��F<��d�����"�v�E�(&Ux�ZӪ l��x�+ٙ�$�e!��7�������_Y�<8l[H.%�}��C_g��t����%9���	�9
ƭK��ڈ��'?�\�֚+WߩZN,����ʏ�	=�pF��קL�N�u�T��,τ����]y��.��7P(�`���1��׵È�}�-z;r�2�4��K$�z�c�����Um��}��rcn�^!.�ly�~��p-#TY�۲S���J�Wc����g5Bk��,��!3]���F��W�q#��JX7�w29�++^�ђU�;ڈOf(���+�&����/�u֜�l��2�����x���'f���[�>&�矘 UI.��)�.��u�j	��3���Hk���-����g-[-��|u�C�P��T�ċ*z�9E�洠��R]��'���@a��r��ۡ�X���ۺ�}Dv�z+� ;��T�gg�����j�YB�qTa�>��J�r��� O*AW
���M������K�7��B�!��C��~��ŀNЦU�l+yJײ���{���]�щ�[�5N����bض�����~/>�mt�!ٲ�@��V#��r�y>������[���$��i����#ܪ�tzk���?������%���FN��y��9Q��rF�>G�Sl}�����~r���ʔ�5l�?�J��U��H�.Q����#O�X�~����������D$���_E��kt�P�+�#�Op�L��)�k�+�����8�%�ގl�o;�m����J�!�#&H���'��xe�lEn��Y8;C.�4ΨE���P =��u�s�/^��n䥛A�A��'��C���y�Rҋ�/��\]����C�:����Z#f�1�ѥ8���esj��w-T�Ys8�ƶ&Q�b�e��.�F�o�_��D�Xf���&��e�0Q`�&�yGbr��d�R���-��B�V{`"� 1pF'-BGuAэ���Պ�Zt3&26�G6�6�4+2N�iCPJ�3�76�P��<��S}���vY�۹#�Y����9rd�i>x'F)WU�� �d����$d@Ų&��k�y)�h�|����/5Tcy�>G5�.놙�����^9V������0��[ƟA�hfs.h��y�3����ΠR�0��*�)�Qs�KE<��V◕w)�����F\����l4͌��H�K�=�Qܜ��u�0iWnd�z��;IZ�}W��j�缜��ۖc�������=�b�j�jd�SS��>ة���W����V��-9k���f��tri�J�t����^u�����Q\���/:���v�K�Ǯ��uh��1�/s�0����:�Iϖ�3���H�|��έ��g'"�ُ���l]�\�����w4����]�ې
��W*Wܖ�M�5^�r��u��. n.�C�*�Q&\�r�����lm��cH��ur�.0y`�4ǉc��:��f�/i���8U澖��O#�.���a�e�g�b���4�=����7S9d�����+�VN�oK���O�f�RY.���h�i�<u���G�4��n,ʼ^ �B�^\9��QR��]��]�]�^�,{f$R�,�ҽ�����W�I7�Y����yh[�	��l�"��.�oDRT��Q�u��LN�#��IJ�;LqѰ:�Lo&n[#�έAS���+5�ҡ^�غ����5�p�l�+K�#t�ly]+4.Dm�������v]�̒����LS�;U��vӮ�c_]nD\�H�����J�E[;�lީ�vֿ�c3jgkʬf$D;g�mA�\�̾p�F����z5>Է��`�wĤ�<��s�3l�`�諮�)'Q���K�} ��V�!=4�v�%��*��)�]�['r��]x-f����T6�䳠����~�yG�`%��+;36u��e������o��{�1i���T��C�Ы����w�a�A�����sxTV�Uy}�C��nA��;MM�J����zD8�Թ劭��;t
f5���Vik�e�Ǖ�u��6�s��xV����yu�Z�lnsp�H6wו�!W�^%x�)�t���$��׋�[��su"tM+/!�7F��u���vUG�i�{�^h���ޣÂR��TY1V��yq�J���p�5�xZ����k<PWhJB�y��M�Jf���u�v�(^�Gl:�y�v�F�e�`�A��Z�zN�kB��盷��
5�����cA�����7�k`�c{c��:��X�#��poPY��h����������!h���hh}EiJi��4Hfs��o������`��qSN��A�a�Ѥ�l3F�iր�hZj�A���s����Ǐ������������i��i�()(
4Rh�=E�
<:��+�j����4kM]�4=X��e������)Ҵ%[z��i)"��-���HoY�=ADG�EF�3�h�mbu�ruҝ��P��㮺���-�0X�t����@R�kC�']`����^c�[���1Dk�.��'D�����N��Ɗ(���l�:Ƥ�5��*�����4�i�еT�k�uՋX�@D�l����4��S��&��hKc�����z��T�os�R΀��������ZCA@vV�t�i#�v#3��r�ѵu�呛{�q��-��ec���ތ!���([�l��N�U-�n��G�������>��q�Mf����X[�z�;O��h��^@��L��`M�EzW)�� ɮm3)B��yi���e=��n������j���<T�P�|��pǸ<��!U�8W�ԍ]G&��R�~�ѹ=��q���΀IM2RdN��|j�=����x<f�t�o3g=�Ңj팭�1��ݡ	)�z�DI�)��N([ �X�ϵ=� \:�:= ���(��C���#��~f$������^ϒ��T��t�&�h��s�]�����b�湦n+Z��,�+� �a��yЍn�LW����dIz�R�s�,��$)�s��摋�F��ټ�u�{�L�]+a�|��vC�y遯B��U	�(�r�4ak����ۭɛ:�g�� ž�y���N��l��}F���z!�q��:ꧤSuGu[^�tbr��]���=����#���K�ҟ*�{���"
H~y"|��gM�A�����I�s��5�w1+�'Xu1���tzL3���Z�I�D��;��CBp�ƯU}�sn�����K�6P�+�9�w7}a��^C��v#t�nS���T��Nb�k�Q�:j�xQJV񱸺iŮ��97GpP������/�����	]�+/�
S��C��.��+�&
$v\��Zn��r%\�nu�G�pgC?!��o0��c�{�Ҥ3�&ک��ϒ�0ŉ��[��8�4���yu�	�]&�����>i͉�&,(geb�3��7遬�f�}y�a�
bK�x�f��:]�֊�֪�iEnd��j�V;�X�j�K��X�[�}��|�����//�%�<�~��P��鬻ܜE.��q�U�Z~������2E�����%\�=뉶͘$8�Nwgn����Y5cudv�-́˝\L��^M2��xO�KӼX0",BO^��zc湬��W\�UBaQ2����ݛ}��#�S��B	�(ʖ�dy�K��t��!0.}b$�Y
����ZB���Ͷ��]��[Z�c��tA��ܡ2X���K�����\�YL�W!�R���r������o,���&7]�^�B@����=�	�r�	�FAJd���ɦp��D�z��֞��\�4��m�O7�H{h	��!�e V�7���*�,/1V9�QE��ً�Y�nn���܏��֪���dA�����}�懇,�C�~��#���w��bf��γ��Ց1�H0U�s�O��6�U�[����T�B��X�A�24�����ϻk[���(՚�D�]⇯}�F����7�ߵChAA�XͼY3�f�a�(��41��oe�|���I��vv��
�ڵ뛊�:��}��_P�<��6���/y-ꥨY��<�w��_��7��-	��AQc��أ\ܪ/�M�G�X{���"���9�=�؋	ێ�V�Q{J�a�'�q�݇ח1�AH|w�|h{�ʤk�}����[�z;��)�uH�)X���U�]<�o�"|���U�P���w��&�b������1��ZdRn���x�%�Ts	�&�:�����<��O;�k�Z�u��Κ ��`��b<��B�^z���0�ϒ+k�&���Dۢ�,��KsM��S��b'{f���1=k����+}?l����Ƈ�7���3$�3!�&�Qa@���x��u��rjs���v���n�Ylف��B���r�4�oh|/0��<��:�3)k�*�(--[Y��ǮwQhW��# ��I�c��k�<7V@ftxJe��I�덛Or]��8���롑���]�d(Ƶ�[Gdz	��5曌�F�GmOڡLX|A�zN��;�ߺ<���������OU�Kd���Sve^[�6�T�p��6�E�S� �Q�!�b��7�Ͻ�n�J�fFV������[�u�P3G	�5�ѯ���^2L��}�C��OfpT�pbW�tw�;5B-�{�ȝ�}[+D-ȵ���˾�ۚӃ+��Ւ
���]-�U��:�Z�Pt0��9������zck3t�y~,δ@Ɓ�F��t�^�.� 0��79�p#�R�B�ڮ��E��܇���hx�֮�cռ4��эA|b����}���j�	MC�Js�؇X�T`漧�<ks�vs�L5���B�:o����=�ć�����ǂO7�|i��7��*Zx�¸�mv:<��ı/z��lliC��tIq@=��z��x�b�^�!���p�Үh�}�~��w���0�U(��yc�b�_�λp��� ��*�[{�hqU���d�-��0e&�i;���L+��brܜ�>�%ߚ��f�{�C�*��v����Ƕ8t��D��g�������g�;�o�*�=j5�P	P�u�9��P�@m�M���Z��&ƈ,�0=�4~��ճ�)��a[�V�����w�ƂS��13�{��x�U�,ƶ-��\��A���^D;k�vf�{�6��r��V"+Z��X�G�����'�+^�G1�ɾ��`���(p�	�y@֜���+>547�:�:cw+����4ڽ��T����0ڮ�緪��:��b��0T��Kw���d��C8Y��O���v�x)f�A�mJnK�ni5���gt�x�r�y�`ʾ�[�ΘF��sN<3613h5X� �R�S(U38�	����^����^~���iNy���u9������@ۡ�����]a�Ʀ������}Zz����5;�y�B��ڻu�rطd6�M���s��$@$���_E��b*�ល%�vs�ᩓy̲:f�۝�4�B�`��ض���y:3k����f��,;��R2Z^;�O�o�}TOӰKT{oӺ�E��z�3��S�gØj����O����ѭ�f�rn��&���3��xe'�_'{�~=��&�����ج��%a��Xr^b��*f�yQ^��JmxA���������Û.:����Gx��t�=ʭe������P�|��L��Ǹ(�d,`&�s�������{yc%Aq\�Y���+
�
�(�|j�Σ�"����	�5�]�Mc2
�S��&�0+ĉ/����Y'�)�P%��&��ۑ>싇U���S[s5�پ�3|�=c�5������*�A`����_'ҕ1~w-�7H�T�nŗ��׽���<d���M���X@!���^���7�$�_)v�nY'�r�O�4f�.���y@��c��ʏ��L��f����Kw'����e��y�[�ǖbv�e/׷�b%$��eo�wLMX��3��gC}^��P$�{ڻ�2v-4�Dkf�X;(�ǎ9تlC;$�5���2[ށ��V̮�u��.J}�B�@�����G��� VOg3Yw%�7���]��xE�|���!����zSu�f<&�
.���j�:h�5�� ng�W���2�k�,��^��vcǛ���k�ޡ ����Q��ћ=�W>�}���#1��~}���n�t�z�_O�}Ro���H�$<��w��|���
p�ܽ�#D�������h^ߜ�a��������֒�a�#hC���`�48ey�<�%��U��%�Z����.�� ^�C:Rpl]4¹4���b�N[K�`����k�pnm�vng����Fǐ��Zیq���1�^�>4+�bK�0�ͥ��<�S���z��F�&�S&���R¶��k�8�����כ?;������فɕ_����+�j5f(��
�Λ5��ܥ��+��}�����2/bj��{К�5�]{;�zz;���e�b�UΆ�Q�ב,�tgO#���X0"ä�꘹za(V �쾺���]�GQ��e�?5����ĭ�g&:�K���~�	_�����0ת��T�?=��_����
v3�84jy�����N)� �v�b�]���W���\[�z�������ɜ�8���^�sۈ1c�x]{d.��͍#r���t�(3ۙ���nA938C�-�Y,&���'6��3��+߫�<+���`78S%Gõ���|w;hУi?lP�3E�]�3��C&?;��}�*
V|)��,��+9��O*���_~�n�XθBok��1��@����ss�d]�Nl�%S�W�2��ݼE��>�U�F�+Qm����mC���=C)�l�pi��$N�z��[o1I��.e�4����i!��j���!خzw�xa>́ ��u�d����1���ʅ��n�RֽcFչ��7�k�����'4 ���^���H<�0���5�{�?��Zd���?e|�z�>�(���UY��@Z�E�(,kˍC	�4��7�CX!|we�~ƥyN�g�hSW:����:0��~⨰�k����4��Y�W�PXA����<<+�g�q����s��0|acuz`c)��j��@8���r���*��H[bu���'�����kw��xIŎ�>��3���0ǡٕ�O0Mz��A�Mc߂0'._<�é���"#/��nov0�3X�\h�zW0���&��X�fI��3��Qa�8� �OX��V��5u�{�d�y���M���ޣ�r��f�ng*��_ q?���/�B\��y嫊�ZzV����lӅ^��:�k���KK�����*޵�m��L��g�p��Ǥ[�S�2�.\A�2�������������9������n����������+��N��*{qs�|��mǯq�tE1��HƂ�)���Ca}������l�&e8!���k�e���,��h��;��� ��+ĚaC��*&v�W�P!ߐ�;�.��+�hܷY�M�ƾ�X�X�H<���<�\��Sܺex��S::Tt4���̉i����'�A���8�l�U��5U��[g�)����ܷlM��AЛ՟��s��闓V�)���lS9-�k�v�q�Bv����%6_�HL�,T)=������ff�'^.���ޝs�\60���*�4�Q �+��5�m�	M!�>w/y*���髝��r��u�jR��ټz׶t��{w������g�P�����Ts�z�6e�������vg��/Ƚ�QLh�I�>�r���eD�p�3\���k���S/6�o���̮��$H��]�z(�a�aK��@1�\�nY�6��zh��#�U�4��M�
813�#��Lm�����I�YQ��9_���ZPX׵Iw栜K1�w��~�8��?T��}W2��ڙo�͙����E=���rJB
��.�s;2�dL)�%A�˹r��v^�o^<D���U>�X��K��T�����c�ް�H�IoN�U�S����_f�je].]1+3�}���� u��r��狊%�L��s/����͜G�r+GF�o���%C���<5����T��&�G^�e�zp�}�}o�ã��ֿC�b�NЦU�l+��V��d��uO�k�8ǯuW>K�Y:�Y�\��o@A_�s��w�~������ٶS,������M�3w�/o���_/��0�s/͠�c����n���(֜�0x�}�9V��{�Ouc�;3��(�m�}%_��KuY�>��5��4X��`|���/��y�Z���hk:Ä"nu<66�ݠ�9Ռ!�wA!�ĈA&���o�w�~{Fo�m�K�V��u[:�Br�!��=z^���oٵ���f�ޒÒ�#,2�k�pWη�=_b��}�ZgK*�Bin��=ŧ6&���W��#Q�jf8�7]fOct���������ֽ��fu~��w���z�������@�W�B�a���ANz��9��A�^<����{�����൹҃&��$�x��a@�^=[ռ���'v"X[�y����>sޗ�P�~uSYc>z}�A�Z�"rJ���ޱ��-t��v;��}�R�리��w�X��Hf���{����ۣ�q���Ⱦ�p��ݰ�(RC�wi���au[�i"�f�
o�FŬ��!���0k���&�a9
�g�O�_P�����~ƣ�dr
r�WD�P�Ƚ���)2'B�O[�X��t�@=��.:[i�3�x�>���ݯ��6��	���]������ʑLhi5��3{����cة��s`�y��wn��Ӵ����5�0?�	���kf[�;��i'����(�*��2�f�=����r�=G�2-�x�#�����}y"K��]�ܲO^����׉׻mgFL^)��b�uvd-��Ɩ�*�٦����l ���s����wͨ�����Y�8�R�k�tv��&^�$�zJ;��,g^�2-��!�6|��<�7���n?����#n��M�؆�·1@B�ƻg��Y����O�T���.�wf�`ԃ�8�~.g{6QU�/S[2Pބ��]K���
m̖A��u����F}T6gZG��~Ǣ�<��P����/�o�.��*, �[&�tڞ�۟/L�ѝ)86t�
�eq��_��ED�=�yUZ{O�w����>���������k.��p�+�$>=�q�.�	�nb<E��kX~�*Y0;ӱ���_��
F��gb���P�y�P�h��q�5gf���-����N5��f��f�;�w��=BF�ִ^�J�F2bb������Mj;Y.S��Ѯ�T�*rꛬH'��7���3�щb-���Ie�c���kN���gJP����q��V`�&T�58$�ͬ{R5�zz�UN�U��9�4�m��n�,��,x��#�]<��%P�",�ݾ����sw�:��.&N�r��h��x1{���@m^J�+oF�ݲ{q���b����n��{7�h�8)Z����6	v�un������XKQ��[o%�E������c�K�L��B��Y9Jk�ke��:�k	u�+�	�\U�]i���m#a7��:N��ㅞ�p�����m�����Q�9r˕�<��H��$��a��KE�Po.��2V���b��`]S5�qk�=�LFsb���ܾ��T;�#%��Uy�Ń>�m%dՑ9�r��%,x�ae}/S�n_f꫷0�u���b�|[�s���8�_d콹�6M�B��x#�k_�xp�k�Q�CE��vУ�r��Ն�Fˮp���c���B�	Lɐ�l9,�ɲ���$��T�p���.ݹՖ�wM�ou7c�\�N{��Wx.q(H���']�^;mgZ��m��J,o�a���
��-�����{�w9w�+2�gu��4��n�4��k�	ϥkZ%��3N�c^�U��)���;ܺ�:g-�$�K�m�����j<�f����.6ir��S��܇I����1�X�{5�af��"��n�+�A��ȶ�gZW�ty���G|��F�6��b���ιK9�@�(����;�Egs+n�U�&P���XmTC)D��)u4_e΋�5t!�k�qj,`�^�\����C�;VM�JU���c7:[�ɛ�xmOlM�P`�6-�$�˰2Nh��vF*\��wC����)Y��/�k"�TʢEX�%��:� ��=�Ҕ�����K�����1�N=����$^��C�������O�:s2��b�ЏRO.�"�9i{���`N^�֨�g�n;a�����*q�ob����u9Q���Wv/����� ۶�n8f��f�Ҷy�ݶ�aP��1�aE�I"�ۏy�cw(;OXJ����W������K;��aK�]1ِ]kB������X����V�gV���[��R0��j�pk���>���N�UI~��e��r����ދB���ZÐ�֗pn����Z��JPy�R����q���moAYV���&��w�b�[��s�ޕ���V�η���!Je1u���=�A��;��=��\�:p�S����9�ƭ�b-��ǲS�� ���Dѱ��^�� ��P��C@i4P�AEU:R�F�h��uPfsǧ����������||||~�����n�ƜT�4�ӡ�URQM�M.��������z}>�<x����~�>>>?^<��?:܃���Ǯ�wGrkZJM`��J�T�Os���@i�F��QF��lBS�Ak7X4�mN��]u�6�&+e(+F�&��I�MB�I��B������PQF$�kZT��C�X#XwFtS���i8N��P�M[;a��qԴP4�6��J����h-a(Ջ��E�&�5T4�J�;j�Ś���]���
���X�MhM4�1���MU��GLQ��h�l�cF���lf-!�thj�8��ִj���#X�k�4�h1�m�E��AD[`t�A�Puf����;��0�(2cA��B�M�L��8T�\���v\}Y@��h�t��3tV�qnl���ͱs������ʋ%[JX���iO����$�l�LFݝ�>�ɫ��-���A	���?�@4P�	��r!�a���M(	�D�b7�7���/�o�������G_l��vL�%�J�V�ב�|b�_���������0\s<:Op�֜�Ƕ//�N^Z��������coyo;u���É�i/��U�Z~��;�E����6�瓔�#��黫5A$͹���9ս���}75%rCW�2}y4ʽ�-�<�ӼX0 Xt�M���˅d5�fw}��6�v��^�0@D���TV5�S�X: ���Ɗ��z:�H���5��Őc��ZY4���Z"uó�ضM�&?;����(,T)XU\���'��U�n,�PN�2�oïk�<���ä��G	қ���$�M'J����8�Y�����=Fwv+����O�"�;�����] �a�`�[,�oO�
�*��
{2�����_���O�7�����]�:Oq��!���?P�s��	e[���ZxKfv;��O��t���vnR��*l��M����Lx��q�h�����HME�X�!�2��K[��	����mڡ��]����
�-N��P�r��*w��>M ��A�Q�ru}������ųw���L�X�&���f�t]�GK�<W��핗���y+�k���>=�9��.����Æ�ki��=Ҹ.��9��YW5*Kc��VwM�@B��'�E�N=�͈LC��2oog��[;c����C��1;3�FԾ���y��z�	�$p�����'��~�2	d㋱�QaV�y�ں��kO=8z�U1%L���w�kGgQCso��N25��2oM�j���ǥk�*	{knP^���j�V>
�W/�d$�TC<@X�k���Z�g#����y�f���	�9*�t�;�����a�v5��.��.��*[���Zz�3�C8Oށ���C	�����f2q��Ʌ�Q�2o%t�ӛ���[ƾ�v�}耇�:>��Y^S�I���c|Hz�O��~�o	�1��+:v������,s���e�����x�z3=�كS��P�΁�#w�E/tNU2+C�Ю=?[�=[�,�֟^G��� zK$!A^i�ƇGm�����S�9��Gx���S:��C-qqw4^�5����=T>x� �@,�o1*8sέ�ûr��v�������*���@��L�K��~z�c+��a ow��ۀ܄�Fj�D^M��S��g�!���!�M�߱��e��f~�nǼ'�_���qI���ߚ�w��j��en�8�KB�{�K	���.S�o5�ܥm�9v��籙o]���͞���vY�ݒ��������yĩ4!�Ǩ���|�b�3�Ԋ�5u�6�t�����qލK�:���3���m�NZn�<�^�[\?�>����}���cp�-���Ҿ�6��R�&PT��7�Z�Ξi��=!Ŵ'D>C��%7B�fD��-�nk��9�p^K+�7�Ru��K"��)�FS���!J�?�j	�2n�<e3�w=�{{)�,�?�k�tf�H�ҝ�z(�a�aHs�1�b�_��3ǚ����P���h����Y!��zz�v^�
60�w�Ut?'��Ȩ^N�`��B�K��B;ח���U���f�ʀ`���#�kH�P��8��t.��Q��-F���*��/�s,�Da��dh�����_�ǌ��a1��s�A�W3t�������m���@p��1ܽ�]՝ܳ���/b�U2͕�loH���o��(���������}�E��{s	�w^��8S�(�[�q�0mB`�ʁG��~(�8y�A}�®�0]�	׳o�_#�l��]�������]���R���gу�*h&�kþ��;�3m��tXP�P}��5����ʼ��R3�CH�C�$@2	5 ��+ɶ	��'k�M�wr=�P�~-�fZlQ����M[1j=��I�5��j�	��M�t��8��.��tLeǺ;3_7']oR����}�ι<���͊��:�~̂�k��XM뽩����P9r�j�@��m⛹�g�]����?�
�����4��mٺ5?dK<h�\v,��[Ѽ�����No/R`lJ��ԋ�E��wX�9��������,�41	�=ŧ11�����Ԕ�@�N�vR�vr|1�U�]��878��u�5��z�S�x`?��S&��Ua^�i�fU����;]���~t
�>|��k�o!��Km�J��D��Ӭ(�ǫUi�P�J߇�e`p1z�|}e��W�'�cM�c�A�26�OW7;��Ó�.t��eaQ�U�o��L��S۽,���R��vлSw	��^ׂ���;/D�$_I箈L�و��(Ǌ4��u:�|�Up�>ߊN���K��F~�m)���c`z
<�+a#�����r�W��Q�m�dT��N��:��;�0,�f/�_#�~�q<�CЄ�Bc�m�4�ц��o���gF/w�N|�W4�n�Ϳ&��\�9�a摴٢'s�+"�=05��O�3���7�L�s�s\?+��Ξ�B[�ېKŨ	�?���3�/�����\�ɸ�9��K�����訉�ÔDq���e^{+��;�����9V����-;���V���wL�2�@���1���MW���fM��}�¬
�*Q����ϥ@N�����R�vZ2�[�kv��Z�"q\۽���S��<��}C�����~B�-ە~7���GE�H��T���E|$.:ݮ���Ξ/WJ}U22��n�ш����%��^+�_|�}��'���^�['צ��s%����yt���gZK���wm�����Os
�;#S����Bd�?7sЗd�>��׳�'.�aɜm�8�s[ʸ�S�"Uv�']i��g�ج$0���7��|�v�ď�t�z��ϰ�P��$�-�y}΋�*,���1BdЪ?z����j����q����I�� ��o�?�H�/h͟b
�U���dn��+:Iv���dLDy�֔增l�g	��[ql��ת&O��;{b]# �J�=v�x!Z�>�>���%����Pr�x����[!����a�1�r;����1�M��z��K�2(�4WcO�U<9��a��5Syz����	�к��G�/���J��!f��ύ��T��XrG�wkC��s�}��\�B ���u�K��#If��Pm����E\j�n�&8��)�g���!Q��ۢN1N�u�u�qҩt�[aGf]���L���c��g�X����ۻ�Gx����c3�m=.����s$�l���a�d5�d\� ;�nn����]#u�\�:��P�JJ/!��<�WZ?O�
����H�c��,����ͪ|�#�ߧ�#�-�C�_��bs�*�	�����ޓ�>�����:%sAҸ����s9�# :\�lmB�8&�ev�u��b��Z���KT.$k���t��ᄠV���c�4�[���u�;#��#}:E�x�&�d��esҔw�o����ò��8��>��U��_A�X^ǝ-5������T��޵�`�͐�ag��db�|�:��[<��Pk�����oM*�{�c�(q����<q�,�룼4n�H|Έާ���Fט?�)���
�M�*�rD+�ST�43�2z/,gAȽ�om�ةލ�ڬѰ�G�"ϗ��3��꽑s�9��VOg>o�{�g�g�(q�L�g��Ɇ.f8d�ċMy�ѽ��.�(�����t��~��I�K��Z��@E�!Ṫ�Q��7UO�L��Z��T�jݿj�=3?(��Wb���MN��P�^��	c�N�*[���1����S4�ө�1U�[x�ý��t(��{P�Fk8�)=A#������[aE8΅un�I��5��p��R.T9�W�}_ J$}:��X6���z�"6���7��3M��u#<{�M�&���6�-�Ot�Wh����]\3�R*�ɡk"�-%����m�T�H��޲i�vM4�.i�a��)���r��N�i
�ͻ
]��<ԕ~ٍ���rܷ�������ʶ� �,����5�h�S�^e�5j=��[��խ�=��OR*J�٫����E:�����drd��&_��]�r���;��������#X����=�7Q��~�f`n���D^�ؑ����E��R��O ������n'_����Զ1�]Y�{m5����3��;��s׽&����QZ󦎫H�F��縇�Ҝ���5��.�S�(� ;[�uL7��T�wu���tS�ޫӴ�ս��k�6��^6������p��Db��Vw��$:'6�cT���e�ꊇ��P��Wt`�.�A:��=�ㆉ�cN�׽V"{mMev�w��:u�б�v�bE���RR��E��
�;���(�wMa���BN7&�d���S�sw~�%��tSU��%_4
��o7�L�5��=9��~s�ג&�������~���1x�\���>N�$B���Qj�#ʋ�Z\)���� ��?H�%�h���@��Bȼ{�b��p϶C�܈q��� ^�6�2@�|����'_�ޱ�W���f݌�ջ,E	PO�M���f�{}�H�	�=8h��6o̷%�c�ĩ������9�t?$�n^���b~��gp��j��v�o���D�?��l�S��g�Ђ��E㣰neyu����͆bE5T�Qf�*��l�vU�`�ѧ��^(�fʩe�l��7au�ʅ]i4յ�aܼT�۞ͤf�(q�ސ�Y|WgQ�ɹ�2(2
���Rs׌l�m����6#;z�n{]���I)J:0�\�V�v����݊�pa��l}����T�%7����5�<�{A*�Up2��^��}=�U�C��l�d�o�rv�{2�B�����4������S�
�bi��^j�Fc[5s���1e=�Q�}qh��z�y���T7�N���A-���k/��ue�4��������6��:j%0���7j�l[�^�����ꑖoj��z�Aݮ�2_����r�?�T��@ޔ��θ��G�=Onċ�۶9��Nv�x�y����ۀ�]��p��&��}�
L�7}T���i�"r~��d����k[8������Y�r:]�6�4��X�^�N����]�s�:�U�+�ib1Iwj��a��Hf�OĨ}��{,�}�LH����N9Ruɺҗ{�4'�?�d�����K�	���v����΃$0a��i�q��I��{����rުvP��8�6�]��xOe�����>u��H[|w�x���u�Ti޴��G'n��^=���E�G�<Y�u�kn�Y$U���oo[��o{4\1H��:(�/[�v� `�gI�Q���.A�T�l.&�ݖ�7ڐ9����!"0�<Yj��ndǐ��c)�s��{�����i�w|~�鳼��7��i�}��j�f��������c6�t��]��2�|9[B�j��Q~g�#�7e
ᘶ
ǂ�d�����6�˒f�v��c�s�S
��o�$��ϱ�ֹ.���uLY�a*��m O<J\HGݫ��������� ����n[�Y�iU_d,���)Q�U±��t3k�\��1�c�]�؄�hӃ. z�UiW�b���m{�|A���W��!u%o�1�ݹM}�=�Ӆ���i����.��@���B�b��=^D�A��3����n��/{���Cl���MS9˽0B"��V��+���o3�	X�+�i����ō}Y���]�����)�庞̉�$.D�X����.+���e9#��iN:����%q�6N�j�;Cu6��:`b���{%�6�I���]�;uE���]%P�q���.mӳ��="M�h������p��nx��jczq>�~®��~�H���yԨj��A�~�����"����!���ޠ�];�8,����Kw��f��e3��|~������Oi�~�_����s#�	t��W�V�7:udx͸�h9Ur j�;Ԯ�fUz�gR���7Y�n�$���Vldt^��[ɺn�ʪ.�KȎ>�C�7ͭ��Ձ�F�fq�ʁ�H�4&p=Z���Ir:Pܾ�}.�3YR���J=Bh��D�3���T==�=5�5�{.���#��}gsl���\�\����i�j;��ݥҤV���S�=K�X���8,�&Ʀ�g�R�J�L9w�W-�B�q����Y�g(9��Uƴ�@=�<4p1���W��<f0qp�G[S^)��4���ol����{9��`k�}�hԂ.�-V�.mI���!�,SA:9�������q�������SېX�s{6픰b�;!�P7}1�gWX9d��Q��Д�J�����.nH��Stq;�j�u5�,r>Վ�=[ȒR)r��n�o��%�K�]n�آ�l^��r�M�{٦��cB]�k�f��h�D�ӑ�c�8"���Ӌ+I�9'��XW�D�:wvA��;5v��n�`�Xn��x�\�q�S6�zq�4r������d�|]fi{�vʛx�a�Wn@�9] �1��d�C�yVp�̵$�/q12xZ=+`�)�BFT*�&6�O	C y5�$����rd�R&Zy0V�7��ݜ��"�T~��6�����5I����g��z���5j��A	a����P�\�[�<��P0��z5v�#o�B`ɇe�Ⅳt���
���sp���t��m��3��Ǵ9�[�D�>Dמ��am5����q��a�r�+؟�0D}�ш9��LAݤ�w3�9o�<��^;�S�����x�3"=�Ub��}��C5AS�)A�v�e4^�Wݖ�b4`+���DgL���W�Wi��H;�ol�L�h�Uw��ŅL"Ƣ�HqU����CQ��4_W�{xT��|Q�TorBo�n�ܶn9�+$e�K�m���dq%^�R�'yU�0ఠ�v�R[яa�#��&�!u���_,��l���ؗ��!м6�〾�9ݹk	��{��e(��-�4V�L��ž����{7d��d!��j.
�uK]U�v���f�9�Y(%��Bh�ޮ��A_9R������3{.ciӄ�|&��[z���[B��[�G�����]�QȮmv�fܜ��+��r�T�Y���]Q�l!�z��Cr�Rf�Ժe�L��S��������[��\e����:�g�!�s"�q�v�v��u6U�7:6A�	�;�^۱�F1�qٷe��+k��S�7�=�Zk�B�d]�m���(vZp�k�o�d��`ǃ
yH��lVl�,kf	OI"�i;k����z���dq��<^���UȴA���`��z��Cv5�e�C���a������͇�iޝ���v�hBpwQ�1��[��]���r�4ĩ�ȯ{ճ�-z�*��6�X���4`���gI��z-	��S3��Oo�����������������؋A��WF��F�q��>]GRm�mkB_n�3ڤ5CY��l٦s�������������������G��i��:-�6��U6Ԕb4�j���-i�ƍhѣm����ڤ�ŋQ��]�P�`��5�[!tj�j�4�(fӢ
���*���*��IEAZ���TG�Wi��:�5�M4m��,X5�+��X�AC����:�ƴ�4�T�Aw�s�SQT]�LKm������;f62�EPU5A5DF�1���4Z�آ�M�Q��1�l4�X��kӉ��5�����TTQ.�M$Al��b)�Nj�b�ݣ�lm��$b��d��1���E�Q���kX�r�U���S��tIC��Qh�Q�8���j��&+vn�5N���3�i�L1CDDMm�*���k����Q_M���:���׭����KYuN+i�o%�T�R�s��A��l:�s]����MvSFKqP=s&�#�vTA��
���{6��û�Wa��J<��ύ7G��4s8#y�a��Q�屙%�����/�����澛��������b�F�#��C��]�L�x�����.!�N��\ViT8���X	��=����d������e���|��i��y˸u���M�F�K��P5����;�������������<�`��a�T��z�w`^" 	gg�"@=ɶ����q�"z\�ӓZr)�fz^�V,{�/�+"��Q\ux#���P$F
�מF�=��؆��Hͭ��[�T��+q*�Ow.e�^k(�Q�'q�xgu%^�>T�Od����6*��7&��"�)*i�ȃFd�n�z3��pIj��t��	)R���j�i�	�����A�M����`�
ѢiR7�%`�#�;x�T�]-t�OQ�ٚ���:~2:�`�����U,đT�ThA=��Xw�q	iW���Gd��)�ݥ���¹K�c�E^Tc�i�vF↌U�̫���ٲb���\��.�E�n����ӣ	ĺ��.[��뵮t�ӄfU�VH�ʧ9��d4p!��zC
�c`�{=C���`ѶÝ��iX���oP�
�g�qn�W_*E_<���>�5�H�#72�8xEO]UԚ��pp�O�U{kϽ&�i+����-i	�["���[o3*��qV}��yE�m�u �d��P����s%.�O��֨���_�����o���&�aCq�.������u��Bp�����f����딸��L<�P3BSy�ȹ�/[>����#�l��n��ܳxr+xo@�HA�5��5���|݊�S�8��9���Vy�R�Q[��n��;n�v����w����W�s���\��O�,_P�gǸ=��Om��Hcn�ეyP�l����n�dǬ�y"�!A��zb�etk$��D����I�m��ޟ`WG�L� !f�I���{��[�y���[�K!Fj�r�oS����s4q����s9,�:!�T��h�&�O���%�c_�S2ރ0�٧y5��-��3/~��m��&�E��'�^S� ~DB#��ZԧY���<����=zӭF���i�U�@�\��̕b1[0f,[g�P�ީ����ɺ��h�w���������tGb��ǣ��\�`~����n��b	�˥�^��I�^��x2��+*�귂�:@&үu�fґt�a���~D֓ٲ��Q�ʾ�s��)J��Ϳd�OR(^�Ar����G�.%���mN�(���UD����5a��t@��"�k�v *�+���
zg���q2��h�(th��O��u�@��U�E^�/�O��49��x�E�����2ɷk[�N�Lgvv��[9�t�:��HP~
=85M�4oJITU4�5�FT��]�]y��Cl��j��6e�n�B�9dG�s{o;P�_t�-&;k����b�ʗ+O���ͳ��R;��0�-��w�i�g{�P�s��Uɯ�{�8�8�U�3��E#]ڱ�g�k�3SvoDR�Ù��i��rG	���L��NmF���u[�+�邒���i�#���h��5�V׌�P8%q�_n�a�A�k0n&ڵg.���ݢ�g#%>*�Qqg�@�Xw�غ��
��=*p�=s[�S23J�n�5ű�E����,=��-�oɅ4�{U�V���\엮��r2�8�˒����7.t8��-���'U��u[`���ј5��5+^!3%�*I��4�?/7�x����z��YA�xn������@YZs=|�Pc�����K˰gB��Ѹ�ۘ��Wo�t{�W��0:�g���WP�If��B��O��cLM����q���t�R8�M��S��C�(_3���&U�lګU�c�#o���B�\ ��Yj��ntW�WQ9�m�bɗ�K^�uC�~ ��~�����H��rRD�D����n���u�y�_A���}vGvX���kUE\M��d��䶻3Em�GZf#�o\�sp|7�z��{ �>�6��o]���L�b
���[Ü��9#]��v�L\����k���Y�Nc��d�7���-D�O���$ W�jں�U�l=t���ݕ؏Z�<E%&8�=ґ�n�3 �nB܄.������w���}�r{�7��7����?�o��J�<�q�P}�S�U/L�>yrg�\�u�8����ɞ��'[�U�z�ڲ5�����0�u9Z��W��� ��x�^b��ho,u�K��Jk3 �Or���y�gd�C�v�D��<�[M���]�˶#՜냳�ɔ:�T�+X�y�oFbs.���}�x��y�"�o#��c����ڠ��EI�%��Ky?�T.7�tqsn{X��ya����GoD��	΂:�Xm������RLY��䧽es�*F��;λZ�G>P�r�u�,j�h֯qa�˷}�锧�R�]u�yZ�1��48���j�v��hBw� �C	�a�6�a��.�����zڼ���[[lo��&_30�בZs~���;~��=>j[�����Y�2��6�zֺ��fl�l�m���i�M����4I���Y�#o�L-p����a�B�]Q7 e���ʇ2��+�Ӝ޿S�y���M�]�u��NfßP�g�V"��o-�{B���{~��k�~j�`�F.z�Wkw�M�^&���s3I���Z�\m]u��z�s����f�˜�^��T�a��I���WVA�����'������8�
��p-EsD�r�r!@�����<�3�Ԭ�{�n��7�.�R��r
q�a����i5���I�Y4��.j��㘋���v>=�<�Gt
y��:=�+2?,魠��Թ}��RU�1\��L�Զ/v���EJ��&b��uý6K�qD��n��5][U]���������6�������͑��O�+��MA�t�����<��n�-󽷹�WlwGf�w����R��(� ��ײ�պ�l�d�	N�UF���Y34u=]���{�=��B�P��)PSE]��O��@�g}�yW��u��l�A�����VB/��.�Q�8�M�ֹ%�/�<I�-o)����>���u�
�Fl�W�W�Ee<��x�����5���,rksY�F3n��@��>����а��dƭ�^��S@�������5G:u�������<����������~�UFwv��a�)���\篣��H��y�}� ��6�M0n3��o0[٧T�Dԃ��zkK^��>���?u*�+h$MM	O�e��Š��<J�:�薖��]����є����2=.��c��خ�O�e�= �nF����Q�a��cE�98m�o2���Y�e�)�zA���^��)���'j�� C�դ����BZzA�o�n
��M��{�������󭱕r�_^�����$lݣ|Zk'���&��7H׼�u�U1lw��ӻVH��4�@��6�s�����z���#�s�rt`�$��E�J>�-����:`+���>��=A�L��;ѹ��N��;>GRA��'�A��ۇ,�
���ٙ�h��>�$�~9���Wn����F�}[��-��5t|Ю���IXy9{�1֌��δϗ��;��'��g#Eb�x���b���g:  �R5bTH����ެV��C�@�(OZ>&�(�hͥ �P6Y���t2��k�ؕ9��Ր�W5����.c'���>eo�q�Tz��\��v\�Y�3��Lq��#���d��S�B{�"�l�U{��R��OM��ME\��	A}ٳ�o���yB��p]w��"�^�/�H�H�<5��^g�m%��f����^~���s#��d���,�`� ^�_�9���c��P�{�����6�_��l�����l�f<m�����c� ��S:<O��M�c�7Z�7��;�)WF�ګoU�|_-��n`J��;Ps)[��`�N���o�k\/+����&�{�u7�,��ڍ�<���]�g;�ԩ=�r^�d]]�f��,�d0�wm�紅(lp�dS-��S����|Z��\�}q�ݏ�'`��@�u�|�T�7G�[��w�5`�z��U�]��9"�Dx�wGh�S"�בE#�Ռg�kx"��G�_�0���/�w�CϨ���3��?u�o,��5�* U8�3���*�?��a���9B�y�����7qow1�w�\&�i�4����ţsM�U�Y!��|��1�?b4 ,�ծU�Y8�UC���ܚ#7����R8���/�d�A�p\8o?�8q� ��]Q�-��-��p��=�Wݽ�c�G��T�<�tQ���� c� H��)6�m��C��/F�MZ��[���=�t~~[�t�ĽkK�kO�*����j�dഞ�S����Ga#�_ҕ �Vޔ[."/{7p9s�n�����)�[,���X�=��Ş�zй-�;2(�2��9}z	��={��7��b%��]9TK�\6o�(F.�ئs����ˡ�N��(Uޏw��ŷ&[t�5��l��a��+a��K��Mh�2�t��b�U�pujE-o�d|CF��t���W+	5�;6Y]��}s�sV�fڗ-��b�n��w����}���2��3�l�j*%�	�����<�Ѭ����-��U����9ݠ�Noni};]:��^�M<xM3�f�X��?����i����ۻ˙��)����\U��j�J�8�=�ܧX;2�t��]�VWNo��aN�15�q��b�`0n�f��[�k�*���+���vZ�̲̌ŗ1�ڊ�A�o��qj~�f�t���*���IU�W�ǧ6Ȓë*�̳��h[2{��[_B�.��T����P�U+�E*F��vgTF_7Q� �E��o^Ǧ��}�K�9�z�
~'�����M�ս�=l$I�N{k7���gn����=���)���
��v)�4�M��#/���e�vӕ����V���ة�n��a���9�zo�SZ��5��~($s��{;<Q������lѰ�=��ߞ�&5'[��廓�49^X���O��gؤ4V�������^;�>7���m�S��޹PVW�7˝i�*��F�k�-��������U�2�uu3m6a���%9a�w���
�,sQ���(�hS�K�����g�y�ޫ��۳��Y�ah�(�ظ���2	r1�����r����p�#��y,�۴ʄ��^����"���� ���"A%��ꆫ��M����guU�c��$����g!D����ں����4���E��<�6��q�v��ܱwi��t��}v�݈$�3)TM���Y_�T�2wi�s;�{eŽ'�� �]�+�����&��5!T���GvD�;k���t�r4�=�gj��5�P	P��W���;W54歭���C���<��\�����b�:'�h�e��}΂���%*
J�`v����Jiر��QG:7��c�t�O�p��O\�[�w�%`�#C�<S�n5=>jmj5,�[7��t�_\̖�s#�Sz���@�
qh��_�R)76������n��ۺ��^flA	�,�F��ޓVS`'�}g&X����[���'�k�\Qɉw-䚹6��S���r�`�ٌ�ͪk��rBWM��B�9Y���X*3��,A��r��X��$5�&�]k���=��v�C_A%X� �"
��Xx��z�3`��w!��o�WKt�t������H��h�<;'oUqF�����10���寉�Y/sF���x���U�lT��v�-�Ik�K]�IÇ0i� �0���o[vݒ�"�P�-ٳ�؊	7�����i�P�|B�|#���3ܮ�N&�������:z���l�`���&^c�/� iWۙy�KzD#i�e[��*7����1b5N٤D�f��rv�n�N�������s~]H[h,l,Y�5G�-V�%k�B�)����9��FQ���K`�S:șW+�	�f��)�繉���Ƚt^�b��d�9�T�^��-�
�:�[�7)�Z);�V��ɕw	K�y+�vl�����Y�m��^]���ukS�e�[�Bl�7rm����%Q�ک�:�vk�y��1�p0�Q�Uͧd�e+=+_o:#�a���x�ݫB�ur�V�3���;�v�p<�{�tz�Ŗ��L�}B$�T���d�U�����=}5�v�x���k��h�OQ٫d���uC^3(���j74]ۼr�I�SHj�Owuf�=ǗO%�vn�2;��"�ug�o_׍��ˮL��`�K�`�-��$�S~ῷ10qzk]��1�X��_/kk�i��F�Ѧ�$��FU�(<�j�w�~�.�t����[�vw4��W�z��O��Ԙt�J��s�|�9�q&���H�7v\��Bf��M�[z��;�z����"6���7��!�z�42_.͜<���om�4`cH:E����Gf�b�;��Tu�j�Β ��	au�n���@Jж���R��W��CN���fvC\�@����	rwr��F;�9�s�H�~��;@�C8pC;U�E�o\�W>�����F����l^���J�$��m�="ُ�\��|$±�u��o��l2,��6�W=�n��q����e��s������D��Åw��Hyw���`�nn��}#<��`�U��,I�:b8`U{�k��ٗ`����;�ޡ�A������uyҬ��WN�T���ѩ>�l�m
+�L����Yy}ABj���L3KW�s0.�1l����cf��e��V>�|�ZvO-��&Z��x�t�r�٪\���q�{dɲY��R[�v��V�9Y��
bK�rk����Ô�_ː�M3�۩�}xDx����n�=x�yn���t�-�Ÿ����!ջ��E6�ˡq�ʒ��2h�iߣ��)BX�qpެ�u���ZZ��ap�UXF�s���c�(�;�w���:���0v۬Fl,hZzW
���3#�,�2nT�LR߮���羿NλӪ�PLk0SN�IAF�11���h��(�w�j��F6�u���kK総o������~>����~��~�~ъ4�E6�W�u=lm�kkQNڒu�(���ڨ���ѭ����9�P�:cX�h�j�g=�_O��������~??_>��i��֭�}롈.�[E��@Mu�$�ލ�Tbtk0�l�hm���"b��5�G��.�m��PQ6-Dv=lh5M��]���b���5Z,�q1���6���h*b����l�h��ձ�� ֆ�:���f��+RPli�kZ�����z"��� ���6�T�GS�������͊���5Gq�T�b�L[m�:(�*������ƨ�M�X�ֱ��]V��ZsQU4VŰ�l8�DmmA^���Z�&�=1���cUQU��5S�5CE[b*�(�����D�EUTL�����A��k�Ƣ(�+�i�*bւ��H!��Ѡ���tF�Uu�uuю�+Z�"����e�U1AN�V�"�խQD��F�Z�ֱDQ	QIF��1�=�G}b�BYPF�☄8jX�xU����b(�j��iiO��wlR2�#���T=�d�[�6�7Zv�S�M��ƷA�o9T�!��!�'�1�P�a�H����Am����QG�U�����<=���)}�c��u�t�gw��nq3�I���r���Q��,�?f)��l^�d�f^d��]���q�He�g>����O�0n3�7�0ޘ��d�����N��7�T�S�}�W἖�D�°f�h��뎗y�8�]��������`��ۘu�+B��=�,��Vߠ���M�?kS�,8�q�0��E��Ys϶d@WX_0^�ɑ�$u��զY�w3�������K��WN�mf�8wG��X�+�{���ܻ�؅��b��m5=}٠����x����~���t+��O3�����K�r
�gs��_i꽉��Ԗ!(���{�!��D3�z��,.9�m�v��k�5z�1�)���D�>�C��F�:�3iM^�`�
�2֦��~m��F�9�OV�k�7�R[s'�[\��* �]�@���������ޫ�n��H�B�&�{)�Z!��ؑ�d�{י����9��>Nl5z�uɪW]�m���������b?1�Q��p���*�[m�;A�u-B'�\��P������}�q�k+G^'5�u�`�v��*s"n�&�6:����똻�~2�o)�����W>����u��t
��Q�R�����Ys�u��،��5�s�V�5l�Lj�"�G:~��?�{e��Q3�C�w'$7���*����u�^���CT����G�������r�c����{i�O]Dٟ6c�h!t����g"�&�;-��������q�oE�w5j*7�.I�E�l셃���L�:-��B��~�����P��DFl�F��_)�Z�(�b��t�ƀ]�j��&�p�F�[�;��0E�[�J��MG-�S�y)
�zhIS)�4L!}Y���wxb��m�>za~���p��ٹ��O�z�Y���&Z7���8pV��ݕj/�ݒ2F�m��oo����F�dz��D�jf�|6��-}������%�$q���}�h�_��%��G�������x��k�R�c��ُ�&�!e���E�Rx���n��6�Q��О�o����l��=�{n�^苔����9��:C�e�&3a���~.5�\� �ã�3��ur����j�_oe��acKw{��f�1�F��y5-c�����������ovx�\����}jF���gÏ9�&����g�]3��k�wc�~a�8+��|s�^����˽ǂ[�?s�,�C���2��oUY
E��7���� H��C�ᨚ��y�":�/��	Qp��j��y*�6�4��ŧ{Z���	�U=Q6z�b�.Kk��5/1\D�gD��u`�g����Bwq��ED��,�+�g�����"��~�!g���F��Fn��&A�$Ʃ�v�GM7��:�Z�����,SQ9�.�o��7"Wn���5�J˼#),���{5��+/���v��s/��cم���%�B�
�j��H�:��W�&@+����R��r#`��Օm[ܙ�j=�ݣCÞ��pحR��ŠWIU���\o]\���.*��"*zꏭ0����!�.u�Ž��U(���"s��O�pfО��ՙ7mj7Ǥ�	|��}��˯4D�k��
�gv��c+y�Ñ���T�g0ޓ���F��X��S}�0ɵ�N�&�-9�a}�x��p�}η�4�=���A"������V�J>�َ���%f11�[�zh��y�[���fp�v�t3������՜�R�&l���Qe�X�F���Lvwu����*ݕw�u0�`F�⺄_���FǪ��Q��]�og�n8�ݗ^C�W��R�J�UP��n�H�ÞB�jh*�N�(��d�J��W��^V��u��}۝�ɠǆY��m����om�\��s�vT)G������b�\d�/��LG`�xl���u�������Լ,�}T��ktl^[���9&�c]wDd:啺�V�]9���6��(�!f��Bud��ot^$"z]V����E����4�6w����痠6�wG�J<�rk�1�r���ʖ舍z�݇Gv�v��v{\U�9��rU�9��B�#�y!��n�B�]W��O�mؠ�x�W�"q
�iIP��PS�>;W>4�j��Fv�Ve6;#�FdUp�V��RYei�tնz���[ݳ��䄛Ǟŷ�C�^�0��!��B���3��#��6��wV6��6�ҳ,�aM�W{tN��ڧ6'��Z�]���d�L"�N�:s��(dqy�/o�`.���ہ�f>��z�Y��%��-�N7�g�k��y�RQ��H���x	��ߔUG�U�gԪr��:
uB�JEI�;�[[wi�j��}�C_�-Kϻ��
�\FH����w�%���)��n��7w��0��BA��Z��F�3�EV����W�f�$Jvf�t��d�v�1w�;����gݵ�6ߜ���(F��ޒq���]�$�{��ʋc���zS�?{/�:v(l�!�nɉX�4�*1Gn�u��uG��k���I�\����O�0�ioTh�'F�d��r,tb>P7���3;>}����[ISR��\���-�l��,֬��}7j����#�h'�>�ܤ@ܭ2����eɽ9C�l
��6ڳoĒs�q�����ci� �υ�{7�����1�\͍g�-j��������pׂ�y^LϷE)������e� �0b��]u禱�&���n=��|>���Q�7	F��s��\-����-Cx�
e�A*������Bk�3�OK�侮�i���պ춥ӃT���9����iuP1��n�8maf��ôd�.4�UBE7�:�_6���v)b9\������{����roK�z�w�!|xHD���FF�?NC8A�+��%����Ҥr����l�荤u�j��W�WV,B@D�WP�b��B�sf���p�FWwǳ�� ׍ٻ���J�3�!���m(�O����W��B�*�2+���g���V�1F���z,�����-��q�v�y�q�����8��w�9U4�5�a�Q^���j�����T9J&�ݳ�51��wSDvdu����e\�V�}V� ߡA��"��|zZ��6;&��^]G9��=�ó�q�t���(���=�N��q�H@~�C�^�E��n]��m�~��xm�Ғ�uƃl����M���X��y䱝59k���>�.���ZZ+QQ\�r����Gd��n-�zm�g#LK.��jF��:�R";dF��_)����H�]ݫt�ܜ(hS®���o8g��-�J���Us��X�Qǖ����xֻ��2:,�����)�u�����k�P\�B�������b!ouiW$�Q�'y���,����-�o��z�){7f߱#�1/�U��O^�%�5��B�
߿}_W���92�e@�gq	�����\f#;ʧ����sy)�W�Ӆ�D@~1�xl�'s��\��3�3d�p�y�qXi7q�*�\2~������{ otZ���9/h6����๻�4��/���֔���G���M_��|����>���eh����¾+T9��0u���nϬ6ވ�ڳ[t,.1P�G�r���6<���o�]_�cgnjb��A��㫁��T�
�d;zi�������<%$ ���嘯OC���j�zn�����" �P�h�M]U�r�#�_ҕ�*�ɷQ�4g7����A����`�;��?����S�޳�6%����+�̾ ���0i�j��Ǳ���ED��,�� ø-�)���]�1��e�j�遝׭��i�FLI3�l���OL�������8"�]�@�Q�Z���r��2�f�RF��;��.�i�uȤT���ӫ:��1ڻ�u�&Cw�u0Pl��YX�]]�K�y�ɮf;�DMR]_&SZb���U���;�+Q�j���e�#n"�B7��"Kg){Ŗ8/�}_Wի��纹9^�w`�U�κ)X/�m$��
��dn[��*���T��S�Ț47s\:�^�Z��̈́��t��sɒ�������bm��v>�<d��9�� �d��Fح2��mt�Z�q�tC�6�Xn�;����nKq���0�.�r|�L.�\g��*�+��X8����>����z]����<w���)g��s�e�����	Lq4�7�g�vv@����˟N�nul��V��˕{�j���`�-���`Wn[bn��,��ɬ-|:���*;�<�z�i՜{�][Cdu7@�0��meuݰgZn#S�K�4e��>q���Km"C.�]߂�����6t�l�M��1��u]���o��{t~x
��� ���D�d�$u��Ot�7����#7��1����}����E�uF�}ѱyo�� ΖM{U��_����W�Xb0i��
�;{�\�%�ے���=s��ފ���0u��ck8.����Ђx�׷�x㢖�����Mni���)��];"��[����Hn8d(�s��ܒ��w�d3�GZ��v���5��+��h^��������8:�N�o����i�2�R������޾OtV~��t�(��0�}�.@����"*n��{��uOd��=��M�{�m�)�هqC�	5��'�5���7+kj��[d.�z�ۼ�ߎ�d+�W[Uʨ�<6Y
���R���4e�W9������.}��j2#��+�R3Dɯ�[ UTӗ��z}7��;o�[�n��g�F��9M�Au�޾]̂��P$�JJ�[��8&�\�ov�xV��4�o!|%��w�$Y�&\fo��5�<熞�c��fr��]-t�v���m�].�ǫ�~H=�U�/)y�$�����ߡ�`�۽����S�v�Dj�T;�ơ�f!S�q����ݍ[�����@��<zz?i���E���j<Eo�A3�Y���9"�7WW�\�.y'ؠ���W���*��o���o6~�9tL�e<��q��y�R���oOR�t�BO֑Q�yu�8���y���p(N�Y\A�r��B�ɻ�gZ���h�r	�j��[R�uoj�eT6&5�����56� D3��e����3��Ȧm!��1~�����͠y��W�a0Y���Q2��k�o%�%"na`�}���Ӽ�r_��gi�쿐���:ca�j.72���;�nŇ��nF�❞��E�F�j��i��"�������x��bm����/�z�-|qX�0�>KMnޡ�[+yb�r����:�?����w`F��-'��5ksuN\Wg�	r"|H=�$��7cb��d3�
���,���R�#r���ʊS�g���w�4V �|���.r+��<�Vm�`�l!f����l���}��P���u��	�h��9���]D���UQ#gCa�
�X�w2:l���\B�䂐�:ڃy��+9�X�w�Y�c$�\�B��ni�E@�nx_�j�p�u�*v������.����kk��7��F�]xM?e[����� �����MZ����Y!�-<<�e5����뱪�a�6Ι$�x3+���u�h��4K�A�e�kz�iC��9^�G�Uk�<W*��O>O%�e�����ĸxyF�n�r�˙S�p"��Oft�\������L�W���E6m�]�N����Ğ��Q�9������T�����Y�n(�1�	��U���i#M�kǙ�� ��<�����sp� �,H�;i�,�c�7ri,�U�}Uc$ ȷ;n�}n��K9��3��M��}鷳4ƚ��k�U�͒��2�ҭ/�xK��L�j�U6u�Ųr��rFH�b8L��E]>��1���z�u�*¦�(��ޝ�e��8�+ueQ!�o�9�%i��޺��[c�n���[c ��l=��e,�YAs�)9�7��e��-iٗ��H�];O����9�FQZ���if�wa��<$�l���E${[b�%L7ɟ<����ω�{�)eޮ�\�������:��W�)�ۡ�ͷ?p�) �Ly1�ٲ�p�♾�Ǻj˲��eM�c(T�wR7�"�_!x��]{&�ȩ�L�{�n��-k�8-���+��;]���TԥB�w][�F�A�k��GT��-o��6��9k�v���s�<Zč��[�it][ؖ�����M��E˘�|�볝�1\�oKɷ`98և:�rm�^����KVZ��2���:l�dS�&|�f�t��ok�J��0�8.����,�K�[�1Yd�J�nP����>�B_i����>j�g;ݷ��Tst�l�Ȧw����b��=��Ln�Abb��lmuH֬��:��B�Yɦ��:Wt�w*E�ר����GQICT^�kr�P�e���W
�6��,0R8����22� ���l���	�ճȽc�f���i�e1��Z.5�wn}�\�L�P�o��6���Kð��{��Å�X���wI�1����k+�ZY�1M�ji����y35��n=�T�>4\-�u�n�쾱w��ZLvݙy91�c<Gjb���:�BZ���c�Ŝ{f U�(���C��˝�uպo}�=�?pg�1�Ee�H�ǯ*��jM�cE�8�\ݭ8�ѱ���i�Cl1%�U-W7cX���W؆�*n��V�,�u���i�=dގ�1�v�u�.�2L �r�.����U�B.�热u6�[��f�-x����;�w��-`{�"�43�d��k�l�w���B�d�u����>���:c1S,�8���5�&�u{f�E���*���(�r�i����&j��n
���R�JK]E��B�nr��)G��`N0ƽ7��k"e���z^�%v����sn���f+�v��!�x�\�م<�-�]V���U��k���m�2��B�tv K!1"
t$2�b-h���Pb������"b��"�
j�����	z*������������~>������ڢ&��&��d�����آ����V��5T�5M@W%��O׷������~?������|�Ѣ��F)��-f��"J���X5;:�MAA_C����RV�㫣jk�uu�li�F�c������r5E1QQ35�S=gUX�61Q4Q0M�LL�E1UUM4IM,CT�ÛK�6�D��Q4w����3Qw���(")֦)���[��D�[a��mj�ъ���"Ys�j�)�*&�!�`�i�	��v�7�j��ƪ�J��X�T5EI7X1U����R)���
*��������`��������`���E$A	T�Ɋ�J�Fb��ӊ
�J��RQ�@Tֱ�JPQQQTD�Hk5Q=l��
� ��f��r��mV���v�Y-cٲ+�f�ةR�mi.L͎�N�h�g�:Jz�s�z�8?x��O�'w��]�����z�e��o@ɪ�����3�J�^(���]r�����ΐ�v3r�-�^l�F���;�ɽ�ނ�|9�my�㫉��lǍ�w��e���ip���)��Q#k�0lV­M���*\�'�Z��
7x)�4�m���j�j��z�H�L:����#x	��k���)��s��J����u�����v���a�<���{o�2��k�i��d�s���]��N#;�ߣ~D����"�51����x�����0�ۑXi:Ƙ�|�������ۯ7�S}���.��3��2v�lo�o���~�{KF:�y�q�֮ͼa���vH����-�vO���h�������ظ���zr&�k�s����g�5�Zz�[c��gǣ�o6����tQ�j-2�5<K��9ǣ��LE�q=�m�1x����BD@=����,C�D�m��3�]O�r��U�Y:�ZԻ��AwMk���b�MF_�y>���}�+��4E���5wM���4,*�n'�y�uW>b��W<!�;����m����pZz����to`���0t�5M��X�w�q�Î��W���c�ՙl�¯�B�ߧ����Fݣ^�����&�$vm���R�2n�-�t�vX f`�U�Ϋu>,����=T�z&�d=T5NXL
������Sё�㗷��`T����n��\�k+�b	�/�rv��xt�]����]��zt�r�G��&��UGo$t�Ǧ��<j��4~��:_�;m��c;���U�i��H�1gG�IH1�i��JF�m���B�0JU���Y�3�ڸ]���V�k�w��c�H�W�y|�}1����Zw��v��D|�-8��Ad��}�}2��OAHj����M[8���[׎x7Wv���I������V��\만wz�*�	nz)�U�H�z/3;���s�%��c~�y����~8LU�(3C�6�� �6r.+8=M9���/,��{���U�*���n�W���-��3X�Aھ���c�XC,d���P��f�SF�[17�M=CT����}�)�����~��J��h"��Je���-�ZӘ��N�(a������s�T>_�C�j	{���%,f��#��c�ZcM�`_����Pt<8E+��VV:<-��]m�@'��gr�ͮ�>�����2S�H>1�����<��B�j��Ycz�n�]Nx�_T�܍:���J{|�������'�ǣ�X�(8��{�~�׾�	�Y^p�<�jo�h�H�)�UߗFH���Du��%���)~����R�ӑ_�xp���G�(��E��Jظ�D񃠑�<s-��)��m�nv�f��]DV
�|�dX�hЊ{F붹�q�͊���:&wNA~����	����?x��gϯ�^��`=%ޡ=yvq�3�5˨Yk���՝-;}�h��4�Ҟ�xa�t �a{�ק�֭}���VL���ڼ<��@�v��ƛ�R�9���}G�3�]�����A�peè�q'ǿ�֔�zҕAO\����p�+"���z���"����e�>�t�~�l}�s0�/�_.�t��J��/Йּ���S���zE��f��|2���+���J�7�s��MZ�u���b��r;ډ��ˋX�����l�D8V�����п��� ���UΘvbk�:q���b���P痓��G�ڽΪm��"��w�CY�iN�Q�n��,Iu�̮���'���ٸ{)k�̽Z��'k�m�ߒ۷t����y��m����N��g��𜝑Ǌ���k�S�21��l计$?5pLd]�� ��w;Q�y�w��f7R�~�6�g��X���An.-�/
٭�&����kx��-<Vƚ:��dj53����g��6b�W�8���4�ч��np� F�&��mQ\^}K9���I�
_g��3A4�#Gv�4�o2^q��F'�M�=�o%�䉩�K�a�i��j����-ᇧ^�7ٔ��w�r� T?�јu�+�`�ō}S��3��g���]a1��9�����s;R��\L�a�̈
�V'��S�aS��K��-�i��^�n�֦W���F�]>�����t`F²Β��t;�A�u���O��-Co���w�H$���(��<xs����FEq��y�'���k����)˫9QW&�^���i=io�
��WJF�9�n-3s�ʺG���d35�E��"^��-A�,m�ܽ��J8o�)f�v�v�v(:���ܭK��{x'>x�������竲-۫��ڜ�5W"M���͜*uBlΖ����:be�7hW;}(���CB�g�Rm�4QUiSA{NGT���}_w_&<ٵ�4���Ή��Y�
;n�.HOZM#���Ny��lv�iWY��ѽ�ZFSZ��bn,q�&]Ҍ'�c%�䂬�������9�Ol�S"G��KW�M�.i�
P(G\��]�E�ܸ���M�Il��܎��#�x�ޕBSt�����M[<�N_��������⪛Y9�z62N�8n�~&���T���}�t�F��o�Kd��c��'�9�P��5�JJ�:�6;�-�>�������nK�A����CZ�i7xV���R�5�kZ�dă����zy�wn�4����Kl�ah��\sD-���S"�k��M�Oj���=��#Dm��³Z;>[\����W���U�cz�S'ڬA�ۙ�{wu�^�*NN���<�!;���#߿e������>5;�s@vn�J/���(���Nwi��T{������j�,p�"m�Lu���9I}v�K�rj̜�7�uyX�w��d��l*��ZKN��:�C=O�M��	�mI�xf,��	ԟ%���e��#c��gp@�}��{�{�$P��[�����Lue˺�n r�oPn��s�`]YG��U�O��i�uH@�W�K���SP�ݓ�8��Pc�j1q9��qWV�p�{ƅ8g�ꅩP�^~�0�#F�j�%���M��SRo:wZ��3��K����-�Ri�輾�,;�Ċ
H�5��,�?�۲Fh��s�]y^ط3��(�(�{�z&��5�q�t�c�����}�?+�D�5�@��:��E;�A(z��<xSۉP�ڟ��C�n޷s�f��;������U<?x��:
�M�=ۂ��unT���t���/�m��{z18��9�Sl9#&̚�U^;y t���aW�����$�	HdvLn��@�u�K��5䒐c�W��.H��dЌ��k螽���գ�l{�2���!@�Eo@͂���r�<�66��u��7��5��3��+{�n���e��DhhyeV�l\��%.�h�@+�tw֬E��?bϧ=�N\G�:�7drߘI��Uj�K��c���y.D�R>��Na������ԫ�N�0����),&]��}5D�6�
���f������R������D��v��Z��&���F������p������>	 V~�F�i�K
i�+.��2����#fs��yӹG]t�<�v;%�
�
�~�7�x�I���7�d�*�s4�mvr���wa�Z��v6@a��	�������%L�nڣ&ꬵ��ӳ�ײMπ����w�n�W�:Xe�#4,T�[�C���0�/�h8+|�;ȓ:E�^rnF�YC�u+U�dm�7[M�VC��(���w�!���T&��g$B��]ݞݼ.	���o����$��&q���_T�U����	�q��٨Y�v��]�mݹ�z�fD�+���t2�h�0���K����5S�ʰ�R{��=ɻu��;��V����D��Kפ���K���'"���L8��z{g����C ���H�z}���;ʸv�N�^��ۇqC��$G�bV���;��_�Fk74�T������-�m~���2�&NY�y'r|Ƚ��8�ARU�U�ӏj��}��]�;:�X��&Rn�2>���w�2k���ߌ��+������;}��@�e��݆7��a[^o7��giw�¹̜x}�ˌ��KO!�]��]���)4烇���e��wU��ܶ#��������q�B�)"-)T���2�6I��hiy����{�oRd�U옾���z���$.�2�t�t�P�ݛƷ�٪}��d�Du�+[9��j�zi����W�hN~���\�b)&��~�����Q��@�G�;��ǉ�f[)�u���y����� ��M+/��O�x��K�2!$���O�&mn��c��Ru��Z�ِ�;��\�0�:a-�JUI�QZ��4uZDϵ��2O7oU���U�Y�����g4!�����r���,�N�k���Dr�Qk~ڲ�l�]���}`0���;���Rv�y,K�e�m�띩눺�u�waQ�1z�����G�c��Ǵk�7#զ�t�K��\�J��|�ѕ�;�0�^3q-�7��n�o+\�A�{�%J�|c\72�0\��� y�-Z]�[QM�O�`L�SSX�()Y2N=��u�*�����i�\As���Yv ז�u�u�Ǳ��Wc3i�qi����.�������ΛZ~�����^��	�Clg3��!}�"���v����2s��V� �ξ�׋�1�r�����F6L�2M~XC��T�v.�'0�B;vꈎ�#0dz��N�"I�O9�5�ا��g�L����̻|�
�M
��GS���^���sI�	b�E������9��7�z�j�V��W����.�k���==Cs#˒ևI6�)I�ҟ��om�o
��sLEmd�6��=q`�{���ɸ|����S��f�f�i:����ƃ��N>�ǧ,�}���#�`���T:������w�Q5�۲{k��}��R��R��W�-��2�H�p��S��4����Uݚ'v&�z�#,!}�:��z��4
*��Q�N�i���6M��#s�+�\@|�|8���)+�u�g����l�
g�?�V���S�8�<8�	��r.��uF2pd����'F=ކ̛�%	�^7�s���#.s��]�ty�Xs�*���nc�+z7ю�F�R*I�.gn�R��Ć�����H�9�k{vX�[R���YW�Z^��Yy; �ɳ�8{,]��m��[�S�S�"����G��5����9R�a>���j�����ӥ2����[�����-b6��_�k�Ge���q�A=�mѝ{\ Վ��Uj�uXś-��͆����#O�IVk�N&ƞ����s�Eκ;�Ӈz`�eS�����f��]�K=E^���?�����]@1Ք.�:rFX���a�fd��z�|�1X�a�v��f�7+Ne�M��iW&�q�;'9��5x��B.neQ�"��0t,S>p������]D�Zu� �:�
s˿iL����b���tٕ�z��t���j(ft���F�W�����|��Xl�}�W?N�zt}����(Ǟ�qWU�����=���{v�cv\n�Da�Mp:,M����{�gW�����׮��������d�QU��A�'�?�@��"����tl�����v*��X+��C*��*�ʰ�0�C*�*� ʰ�0�C
�2�2,2�0�+C*� �2� C�2�0���C �2� C*�*� �2�2�C°0� C*�"�2�0�C*�*��0�2���C
�2�2 @0�2�0��ʰ�0�� ��� �
b22�0�0�0#����0��^ǰ{D � �� �@ �T �D �  � � � �#� !� !� !� !� !� !� !� !� !� :�zD �T �T �P �A � � �a@	�Q �D �*�10�0�� �C L�*�M00�  u�C�2�� C"�M0����0�4Ȥ��$0!��@�!�HdB@�!�J@��;�zP!�eXeXa �U�U�!��ʰ�0� C*� ʰ�2�2�����(=|�����AD&TE
QU&O��o��?�������O?O�tK{>m�~۷oW��������3&����n��#��Ը�7��`ETW�����?�?�DP��"*���/�?�?����K���P���C�*�������������� 7�=�D�����O;'���_��DXR�@ " � 
T &D �@%$ 	��@"� $� !�  ! a 		@@ �� !d 	@FD �! 	 ��  d@F@ �e  �d V�	U�V !�d�d�	%a%Y$��?�E��O���S���-("�B�߃��u�?���o�
��}������ETW��������O��O���'g�������g�����ETW�~�?ԟ����O�
�+�QQ_�C���?O� Q@W��=��{�!TW� 3���`��k���.�����?`�����*������~��*���<J��������S��x�?������?�
*���x����DUE`��1�=��;
O޿���N�����f�?��A��?	�'���"�+�=�C���S hv�������O�}�/�QQ����}v"(
��?��OO���2�?�1AY&SY2%���Y�pP��3'� bB��>�H"Q!$���JQ"�IPJ� ���(�!*UR���UA
){a*(��U*�%!EH�T��*��ER� �"���6�*�ک%TP�%*��@��(TD��JH���)*)��Q�"D֥JUM"��R� �T(%�`��*� �))B�Q!R���Zʪ(����
R�"
B���UPEP�*����*��TO   1����QS�_n�3DcJ �������Z,
��Y�ke:;��,��M���1�Ͳ��tʻQ��((%����JVhR�T*R�U(T�   cc�����٭5�S��p����{d���U�k'z{�)��f6��m�<�f�����U�-.���Z�.۩*[h�#h�-��0�V֥�k�m�)�A\l�J�-[u�(�(�lBIR��J   ����467��ͳC��j5� Ȧ�&髵
[#)*R�&K4�ջ�CjK
Q݅.B��Z4�5���M����Lj�V�5n��U(� )*�T%"���  ]��jU֑�b��12����[V5V�"��&����-*�b��e jL
�B���A]wmf��(	�%@PQJ�*J
J�U�  �j�����UEl�fiF�{w
�*m���	���pSV[P*�Ѡ-SEdT�j��Q	*R� ��*C� ��i���4�*���J�Ko]:+@
mT5k`SVR�Ӷt�b������-J�%J
T
*T���  ]*#���j���SṾCiY@�ElF �L@ pv �1���Hqa�'`�w l�sT_Y!P�*�T��)/o�  �� h=��@n�����w����Z(
���� �A�  �Vul���F �0� �]B��*!�	*�Q�  68 (ۜ0i��ܕ������ @�A� �� ���C�(GS�vP )�Q�ts�8  ҩB	PJ�QIUB��  3� 4 �� uӥn�p  ])`h
kuV�Ѡ�����mE�Ph ]E�h�f� �kn����S�T�@4@��a%%Jh42 ES�#�1T��h�)� ��(� ��*R��  '�R$̪�  ����>]:B���IΙ��"�{Ɔ-[[S�}Vvɝ��3��{՝v����U�m�kj�mm�Z�km�uj����6�ֶ�Z��[^����������?�F������t��ʷ	1��,D�@t[zi�T�RnIU���&��*��l�-�]'�����+$+!9�F�"�RяqF��,2/l䎤0��ۊ�Z�(�b��HobA|��DPZj�Z�'uT�In���۬Е�k^]��q�a����d�oM���ƑĨ��H�cYKUXMǀ9Zs�r|iK2��Gu��8v�b�X�%,nb�*]�6�������w��G$�ᎉҥk�Jع!On��[�H�u=Fڲ�S`k��ɼ�0�KVUܦ�����V�,u{��ˬ2��\�� ��Z��*��ȍ-L���'`�N�
��د-�xj�u�m�v�M���7)#bMו�����z��\��2��qa��5r�C,:g_�{������65Ea	/ef����]�����{'*݇��LK"�I�oV��\A�:��$qںL���.L�5Z��r�(8��y���,J��`��d�5&P�Od��*��b�WV�dK]a��+l�0�G)̈́��lՑ�[������ς�aY!xt'�|`o2((XP�R�v�F�i+E����1�y ��nE3N45�Օu�b�q՗�UҦ��$� ��NEFTE�ff|�2�e�D��c2�Վ�� h��e(���L�7)�!�x��^[Xf�˺����W{��(k V�փbŋ��{ �u�L<�}��Ua�3#'9;ǳ(]$Q��:�k��9WYXn��t���%G�f2*��9Nm 5�l�һϬ#m�ͅ�+�[hT^55�@:5�ݕx�,n�+r�]c7��N��{vVk����J�Fk�{@D7i�(7�Y�����m+�v�Ȝ� pk-أ*�X�/�6�k����'wp��U���f�*ȡ�n���Z�O)Q	��U�ˉZ�_��=R'�;���N�εVf�L��h,'���,��Z�(m��Te���3Ee�j!e��)fVZ�m�YZ�!en�
���a*��x����T��`��P�׳4�������8j�5H-���b�PnH�+k
�*�w0��v�F��,�meҬW1�'fRX���m'n�ԛxM���Tv1c#��I�f7�[V�6���J�Hd4~M���&ܽV���f�5[$`�U��CHaM��k3Jt�會"Be��:T�͡NS��G�=�v�sHrT�Q�XVT
%]��̄$�֤�Kl-�(��~-M���B����t�I
���D�A7���ؚf��-�κ�UvA��o%������-�B���č�z&�{��xiM���P�fH�4v4a%�A�� [X�ݴm�p����]��̺SSU%xm�1K3>��\
�ɏ002e3N�P��Uf��"� �b2��|���Y*�q��N��P��x��֥a������F�Q�Xv�2�] �w�N$�g��[�e�體�R����	��.����Tb9a]����Ï(�4�˼i�DbWw��ʌ죨8I$-�N<@*�ۘ9��ALR2�I�F���t�3��ʘ�\��:dҏ7uJ�J�/n�a6�i�,At׌�Yu2���d�� �S�7^�a������؋$ӷ�Ȗh�c4��1T��X���3r��*7�փ�m�弊�S����I�V0Y�l��͉� +J�+�X���&VLm���{�i^^P��V��j��+����͗�w1Ū�"�����Nnu,�An��e�íGX��v����R��t�`6-� R�Ӥ�2�PWQ%):k��1�����&YEn�.'R���Ԏ;���
�6�����;�P\�N�kCF���u��/*k)�$b���n^n6��Z�Dk�:8u<e��o��-�6ŷ/[�:B$�zW���vf�y��V1���2�H*V�b�I9�6G'ڝ*�j��ͥ�d�0�[$y�X�=BU�d�
��H)�q5��ݛ�kŚl��N����d�r��p&ۗ�h�L�Pc����X�!�k"�X/^������hIm�$8�n��׷������iYWRlW  �向b��7y��VF5��V�[�-#UTEڧN�1-l��J�������h� c���N�XZb����M�ZѴ�=���i�` 2��90�$�1��:zM)��!�7�S3,-s\6��@����ZkRKMa{��K+�I�]0��寕5�{K r�B�'ka�e�ぬ�V�x�)enH[�
��O�	={J�/�Ob��Um�B�	F��ˣEh�7.��ME$�5���X�n�d�D,m?�����^��x4`{RhR�=��`]J���m�.�w0��cQKj��8�%뽽� y��N ].]���0p:�Y�U+�쐃X�6\���I�����W�E�tmEu���8K�+ef]�ic��;
���[s7,%���"�j�;#r�&�F`v��
��yE�uq2�ֻص������:�QaZ���ˊm��cPG���dۑ^C'�'n�G>���J��d}�/\�d��T�S#u�a^�۷ikE�X#-k���͘��KRlIZ����pVb�SW�.]��$�j�+�k[�YV�:�Mma�q�.nݫ��,�ux�B͚L,p�邱@nL͵��.�9���!"�X8�SW�$��*���C�[�M�֨Z��^+�`���P�F��Jd -�J��3twF�˛�$b���hlKOU��ɑ�`%F֖��6�,�e�1� FÂ2F^�U�cIb+1Z�ݵnQ�3>@���ء�+MW��
�'Y�]�� B�3.P�x�z�1յoM�TL�h`��SʷL��(LI�s�+^E�f@\stq#��َ	>��n��Q�^���Ksf�yh�8Ӹ��Ҥ�̠%٥��Z�S�u�ҭL&�G�\��j�@Pd��њ;�Զ�tp�؜ߖ���#�[m��N]���&f���%-�K%�ɪ%C!��1���7���-*yt"./�le����6�jn��TTķ��+U���̱$�����4H,�4��-I����SC[��x��̰�͚�T*� ��tk"v$4� -	��[�*�)U�S;��Lܓm�xৈ��*��u�5�`�{���R��4�UެG�86�G�j@�,�����15:`��ӗbVĕ����+/�<�#�IaB�Ѯ�0�6c�(M�k�5y.(Ӷ��t�[A�BXĭ����ȭZq����n��'��"��Fkz����2h)l{%�sP,�aa��4^��#XSzѴ�`
	^:�$o,���ؼ�˽����,VdK]�%^��^u��iۓ	�����0*��V��r]�f�̑�&0ͭخ��QV�e,���H+�!B՚�k\�dA��w��In��R��в���f��y &aF��=���L�.ĳ7V2�K&U��PbbT̩��m�ڹ�3KB
sPڥtIq`R��V�N1�1��^S�&Q�
Sq"�2�o�F�"t�s&�QX�i�j�
^�ʩ340�B\�"�W��� ��yW�Ɇ�F�$�E �ʹ�a�B���lMX� #Oaò�4vqiO�\yQ@t��E��/ p�*C��;[B�j��5B��8���om��(Mi7�fB�5Wo#����WG5���������&���
�f1�`��@.�	"q��e[L/�1��'���M3p<3N=�m�!��k��80����P��f�"w�v�R�T3d�acY�b4D �Fݜ@`{����h�B�����d(�aG3 �����6�����@"4�7>�L���'X/�6���Q�aݨ�$b.��w`��QbyJ�R��gY���Q�v��A��k�2Z�ݙ�k*�#�Au��mF��k6Ɔpeh��Z�=��[`�O@ǚ��Xp�Vm���a)RaW���fd�ʄ[8��N���Y�*^5lr�Y�')�sY*�����h�d�[���u�*�bϵ����b�	�2�\""�I�/v�d�ɩ���ᔔhiڰ�5��@eHl Z����:����M�0hd��+�a�y����1�*r;�yj�U�s��\�QS��U��5�*e�C\��m�r�լM���;��E�TZ w.��V�k5@��aV+xjH�4U6�̡�o�-�6�CD�N��M�y�'Su_�wh]-:)`����$M9�Z�pQ��SUA"�*�R�c�&B�� Nc�,�t�,��
�"@��#Q�n;�ٺ�"@�v�n{u���@L �F���+ѹ���W[i���ƀ���v�66����ݽf�Z:�������m�D�b,T#�D&YX����ˆ�բ����w�s@�6��ݒ���=��Z�2�a���35
������p�
w���tL��Y$\�I�{/!�kS17�l�.��۽2e�iH���m��t>9iU�G�=ӁXR�ذln�����:�ZeB��[�*K-���5�0�ǔ[����L4nG��T^,g��l.�s59��`�#/ �C��k�4�gn���ٲ�{n�ڲ����q#�\͌��XƹcZ ��m�@6ܽ��mm���;��nP��x�Ӧ>9I��Z�2�9�vN��Rdoi������F�f�T�R��^���91I��b�r���S�["�]��h6Q��T��KN�^��D#9J�����e��2i �B��Z�pm�H��������յ�N�e6v4��w$�MK!]p�b� UC T�M8>c�I`e�� 1KU�I��S�Y���e��Y�Q�:�ӽ���Y:���Q�iU�XtD�ݗ�D�j�S[O)&�R���� ���zEI�*�f���6�T��`1s&�ݤ^V[HGj�V!5[�j�n�J� �A�u��B��
� ܏.��F%M�J�J��6�͢v�ͬ��-\�]5��J�ÆVeѺp�R�p(e ���*�NVan�hݻ��wE�oo�=Xi�U-n��2ؐ�v3[m�X�~%&Ι���x#�-J���`"�޷�,V�x�X�6l���#+v�T�n�d��v�kbM���[��e�.7S��ZNVd�KMʒ� d3mCC��u\�r��9, /)+�r�5�E�5c%6uS�xJPYZ�TBXC&�r�ud�,ڣ2��,�O컖b&`&�P�h+�wG
읷H�1��(n��<,��r�%Zn��U�#�sC@�u������z�s!T&�W���qK9d̗"
�+p�V�r&�T�td��F2�T:�c��eU�۫V��gM�=ȨQ�"��%b�[:!��S��dc ���,c�>i�lح�bc�hffekxBuj"Y��7F]��B���5��)f�M++Q�l�N���PP�:u5V,aջ́�K\+%۴6�h@Tk$����2Co�ut�觕��ۗy��^�`aa�-�&�z� j:�m]��(���k-[�*"���+N�̑×�n`k���J�PI�22ԝ �#`�t��I�3h����`�ч7n�f�n�P�b�w���z��@��˧/Q���n�{r�q���� ,�.L��N
��A�IzaV�FS(1�/l
m+�b�/vB�w3^+zUҖe��0�7oa�T�R�j�d;W�1dwV6�DTd��A�yy(�n��05�V�B<`LU�c���^����׮,DHx�IZ���\5��RH^>�kj�{��#�"��6X�"f��;�fT�!��ò]{W��\�I�v�fM����U^:-nl����2:�ȭ�1[Ibͅ��� �PIF�!RG[��RB��ʊLXڿ����)�u�*R����<P�?E.���-�mY@;;@d[Ya-R�Ř�䛕��╙�"�j'Yq�m��i�QQ��֋Ub��f�R���^A[�nR18��HY�V8��𧙂�V���5�m�*Ө/��y��ް�l�f�vT�R��/�ȭ5sq
l��c�JL*��e�Ŵ�X�8��6��v4�gD�Vc��fZ!�iU��*l\���0ֽ�U�FGی:�5L5m�	a5�[N�Z ����sl�0��-S�b�;%����̻�&o���۳MǸY�֫�Ub2mf�2�B$�vJ�D���w�mPnS[���80F0��v�N�觏��z$���]mի��ʄ@\�ю���1��]b�J�ݫ�+'��xʍR��`�d�,��j㧢�YY�IQP!Mwz5�2�N݅������jƁOv��)��l����	T�.��"���,֑�wP�;x	fnCH�D��*�����y��7��m����SY��w*Ĳi��Z~n�ߚy��Re�쵈�9uhn=ߦ�i��w��k͊,�Kԥ� �WWzնn�:.�������0x�yl��J��^$�ٖ�^�:3$xx%�i��	�L��l0�`� eH��o �9HL�#+1�2��{m��e�U��ѣZs�n����[��ef"����A�{�@kfhf�]b��^��ԇ�&�,�C27�]	ETYs�si�NL�k��w-�Ż�]��)�[�%�k7V�4v�඲���5F̎�V�H�Ѝ(�;Z+p�u��nc�z�RattZ��cBL�J#BԆ�+�!VF�P���Zò%��WƱb�.��@�G�U'X�3���,�M�2�v���7@EKH�轎qS`��%f�DP]�nS"�".��Q8n���bä|�j+� Ns~�#&cH ,����Q슭mPdI����RuN�;7*U�N��:�X��f�p_n��HDr�m��%�i�gW}aCy�����u����)wp9>�@�����ɽna��5���FB�^�->�p��;�M��K�6͂���N2����8 㙮�N���0;�w z��V�ǵ(Mar��u��1öf��.*vf�N�a����q���	�9^��+[��[��Ry"z]S0��dV
h.��^���d6/_la��ّ�K�Yt�����=�B6غ�J��\sD�A�Ӯ<8�;��9Ш�Z㽃p��Vhɏ������Zf��E�u�qG {')[B]:�N�&�U����|�'+�l;bnF3���h��buet�x#bݲu��Md���B�����|�e��a�\��S��5�ܫn��yt�*�4�{(ou�$��2֧{��49��rU4F*U�|�΁�.�<��L��N��ȷ�aK׵���M�K��-��U4��Bþ��zÏ^c��3�RXEbw�X�HJ��;�Y��\���SUg�*�u�+���/"��\��Zw��5�J֕�uЫ�+�TB�>�C#y9@e;[��s�͵��S*�vf����AR¬Ρ
�&LO%���{�H�Ȕ��r�u�枽�$b�؈�*�}�(��LU-bv��'�'&�-otmc��b����x ��ʛA����ފ�N�"��v�A�!����J�\cv+D��r2�7��
��`��w0�.�gu��	n�,*���k>?Mk���L�p(n	b�lq0v=8�[v�]�Nk��{�9h�l��9�\�3jb8��҆*x��9]��x���=�t��t�.Fe��˺/z��$�;Z�8��;8�H�sK�`VR���B�Nn�ƐUՏ�OS�g+��ۥЊڅ�ލ�����d]3���y�4&b&���YR鯞��+T"׆cg��W)NS�֜�(��xoX��=Ҧ�]�/�B�^�Q�Q�α�gN�8�匤nǵ�쫘��6�u[l���W���V_���x1-譅�D ��]Hj�9����,7�E��}Δ�4u(ή��K���E]f>YĽ�$t�<�5��GEe�[�Kr� �}v�k�X�����JI�4ou۾���fA�p�Ƈ�Nzqk(a\��<��}@�ԫ�8i�I�5[��b���'*��@qۥ�݉���$�v#��@4��Q�vE�9佪�MVG��5,V�\�kH�a����򞮾�,͈K�oi췣�!��5�n�ke��gI�3F.�-4�0�����M��&M����F��3/�(�m�u��Eך�����
���)��E)�x���+e�V
�̘��ߒ2=�^�+����w�Q
�X6�c���<��ХE�˯c�RjV�#�#��F�����4���hk�㾾�fU�q���`�i��ϯ"��u�
c���F��q� �x�:��;7�wtg{��GƱ�[�VRlJ7W{��C/;F(6��T��ޅ9�F�!�`B� s��kjqv�"8�t*�8i*P��_#t����Z���ݛجĠ�mSе��Ҍ��0)�u(nU�/m�\X��$8BA�ݶ��=A�T�����+9%�Z��B���3�N>.���7�Յ7��e�{|o���$	��6�c�ܶݝ��ib{����}f�O��P�B��ݛM�GVt}��V#���֒�ݎF����C��ش�;����o=Xkʹ�2�Ĵ�ըgP˝�EU�	�r��OoSΙ��IwK��bU�pu���-���m���:��%Ge"q���Ό�]&�]���k��J�G���W�VU��56� I�i��^�7��K.��7�b��<[�%�suJ�ct�@@���B��J�7��Υ����q�lQV�6�
�U{>�Z�]ٸ�=*���tٝW,[�L��#\Z�T��H�kp��Q�RB��m��S\*R�xE��n����̵����5���)�bjz�mK��j�8^Q��a�w&��[ݱ�Y��v/�<�;b�4<��-��%n���%�'Nɒ���yZ������r
�9�%1�(%�P5�F���ՀC{Ԣ�gIXU���*R��7Դ�ڗ7����S�˧K
7W�l`4,	�G+���N	���;29�փ���;+���5'7J�9`=�]��E �z݀�Z�>[��ީ�]s��gr�z;X�&��}��珦�&|��')�b��A\�}�a��m���WJ*s>�{�-��w�LC�V3�zՈ`�J�^�����jQX�z��GD9vF�j�B9XҡqVwi�eӓ]���ص%d��W]�<z9	u'v����|m35���tUff�ͻ}Q�i�j�0y�шu��C�Rg���Y[O�!�i8t-�k3��̎�b�f�[}�sI���v_��ǚ`��c��>���:�`�Ce�Գ��J��� DCJ�巗!��׋���q���P��8q�}���$w�Zx�˕;F�T�e��#�%9��b��ï��5rR���c�뫌љ���LlZ#�,d#3��b�m��8H"^�\�=����ǜ��=+X='p@����!�r�X�tS����C2񩪵�}! ����]�ff��J�2��]:;���Z�Jʍ�{)��s!*�	JB,�YG9�ʜRHi��V�� [�ņ�+�r	RN_^�}]r+���RƄx�w���`��d���	�y�|�[|�����>6��{y�!�}�k쬩M6�<z�n�ݹ��N���Hr}��������9C��8�]S�T�P̧7gNE<��f.���ƣ�O��+r�<c��ڒ������%��bΜ�2��`4
�K�z�)��SL�Vnv��|�q�,���(ٝp�ȷ�[��wq�l.��"s7D���˪S�ڏ]5؁\3V᠚([doN�l֡{o6p��c�v�����x`�K2�Z�}ܖ�}�յ�,֮譅��u�K��Mժ�u%�(eTL�J"����p��M�W}3{z��tW]��a���+��zk�lsO�Ol,x/���}��{Z�	�N��/��n���Z8�/���)Q������z�eu�ۏy.H��$��ip�9����P�V��Ia��kݗx�K" ��e>���-��V[*%f����TRɼ�z5w[�=��Q�����8���9�	�h:A
�oT����fk�{�g5��v�T���wc묦�'v_L�.N�c�5�j��-`�Κ��ٮ.�g+��|��ڡ��>��-ް�+��y�MmX�t�4�{͍�����/�q�" Nwy�xk��%@!ly�H��E�C���r�E3bsj���2^T7��89��-�u 5��q஛��yt�.��q7%*�t"�Ķ�e�>|ɛu#!����:�)4!��2�JN浢]�������s��I�5в�(ݮ�>�)�Q�ظ���	fv<)��hL;��q4�r��4b�밊���Y8+1f���A�Q��ˆLf�T�ٵn:U0���õma�[yZK�\+*
�R[#4��kU����]��#C=�ۙ�L	2�z�wm�6R��.3��
5���K�m��X�ʗ'��S�-7�n�ɬ��(ꋙ�T:7��b릁rX�7�jѹ��Rۓ#h2c(��%{�sV���gr�b�N���]���׀�����/�Y�:i��L^�v�o�8KpF��V̲-�ۑN�f%��J�ɥ����5�1���#�KjZ
�V�rV�@f�ⱎ���ř�7Th�Z}�R�l7�uAM�^�I��UK��w�����J�W��;4q)O�7I��i��v:������|Ca>��4�t�S�B{[77@y[��ѩ����j��ʙ
lﮈ���KF���˹Z��e䵸"Tr��g�)-�aim8Ƹ�+�V�+[rF�d�W���c�&h��� .Ŷq��L��5�2�Eq�9Ke�]N��4���.L��#��ɖ�⊘�72����U������2�ٴ�D�f\Unc�)��Ǖ�7��۽�\��&e�3��Օ!7�f�X��Bh�;&��L�i
<��G��P�+q3����;����B�V����f1�v$]srU6�W�{��4��li:$,�N����f��نGθ��YtU"��8��+*Jǿ=wp����l��p)i0]�t��MňZ�ےb!�)�����M��y^tu������Ô����T.oh6	������{��&gL�3�inO�Ng�����mKR
����Ӵ�3joX<'���P� ��(��.D r��c�/�c�
��yD^�[��ٚU��iq��4/B�j�4ZȆn!m�{K�����qƝ��g�������rh��A�k���Wr��0VGE��x��.���	i���Rg$T[A�=��w܆�ҽ�"��x�X�^��Ͳ����� _m&��+�C}m$jU���}@W.Z�a��̐6���478��s���fq���X±ܖ��§���mE�Y���7]�E�!����㻷(����M��}\���v(��OLw��X�8�F�Nͧu���o�uf�}ݼSvл�p�!� [T�9��E)���@������Y�W�$��\}���*�K�ƺ�i�[�-;�s�ΰ�%8�����6���jv�Z�P���	�Nl*>�v&�x V�=���ef��E�L�]j�6�-��n�m�ʥĲ27�w�Xxo�/'���zv�IѐP���X������u���PD��������%��3.���`�J�tK'%vWp(�&u��c2R�s��Fo�6��.���n`�l,�k���1s��J&m�!�
�e��J�̭�����Z�hZl ���E�0Gc�kou�l���S��λ��8�Wr*rK�L�+:�̫���Ogo:.�l�]���wc"$��/c��'�E!y.u�9-+7��
��X��6ղ���83��+2ࣙ�$��Q�Z�*!�[lE�;�U{���t(�r�R<�m�>x8��mg�L�"�{*vMfbǽ���Jר$r�^�E[�J�љ���`/3��R2��d[a)���'u�Yz��v	�w](bբY��/�lu��mDė��������xZsBkn�~�\��+a����4$��[�<;��p�2�hb�+�JE�4�@ i}�Ņ[���e�V"��Ӳ�9ʹvr�KP:ob�U�N�v��څ=�oúv�W�K}�Mi�ңy�{ +��G9k\f�8rfɂf�kg(|dΤhm��AM�/�}���V�1CG1{�K�p&�N�xPu�FUp�/�F�|�6��D8�v �EЂ�K�n�L���@��d�ô���
��U�ac�[뇭��wiܰrcapk���&Q�v� �=G[�3�G�۰�Tw����6��R��xK<��RM��,�h�s�w�ym�X+�E�4S�}ݛAv	<L�{/�=�Vjg�gnb��!Y/Rf�͉�/��jj��ԭ�r'�h�N�ài}|u�*�b�n�r���x���c'�s'AyNށ�-3,7.=�5ا|�8![:Ć����糯�<q���*� .�1��h���|ܢ�n�M�F���FE�T8�͖�p�{�R�^0�q���T�{vM�v�ޛ���dK^�D炬�q���t++e�L�F`E��v�������=R��,�ʎ� WO '�����޷�pww�ʮl�'s����l�]%�.���4'�Jw
ӽJ���x��Ğ�[��A��y{K��n���+����G��;D��h��u���kZv�q�sl����滫FrP�]���u�����y4:�M
�سg-����2�OV�����ڧ\�nX31 ������[Oq�qøtc�y�d��ݢ�Ǡ%u�'|.]f�-�
՚�t,�fw\��C�X�K���$��u�6�P}�b��b|������E�j���a�v��x�d��PCj�L��V�X��ᘖ���'L��n*("��'`�X�d]��`|�t�sZc���V�V����U�J"əӝX<��Ѱ���k*�p���s�v��oiN�&�H����i�eɡ�(V�����,��S�5u���o.�j��T�(�e�C��ޠ,��M�(�	RZv��9B���j�j�.��Jku��u��.]��..�U�Y{�<����ܢtuN��B�v�E����B��T,���v{X��U�
��uP"�i��Y�Iju i���o\*>҆_U���=�f���{��֤(�k��S*�C�Jg�8�-"z�G���p=Iܫ&+��n�\�R��X�'D)Hr5rI�>��53�7��;�^�=Iw.}�ʌ��&��w��4�]�ۛ|������k��k�o��a�&I\;���8���*�m�-�r�iF�tr�ջQ�Ν���xV�`�2����s�f�塞խ�7fC��w�WwA�y�5-7�]][e�����_^M�5;���S��{5fq�'ۂ�� �W�oK�S�"��&��[O�����g^L��W�|n[���� x �^�����R����s,�oz��'�����vV��ِC��$X�*ŔR������[R�<��dj��;�١ZM���%����ݠ�b��{GHo��u����#�21�W���uJƅ�]s���dtۑ��f����}trR��n��;
E9	�F� 33��Zt�o^(�h8��[�%�FQ�TvN��xV�٧׋����v�a6L땷3f)/p�=w1׮�\ͫyb���۲���o�Ӷ譾���fJ넚 *�P��&sX]qຕv-r����̬���S�]�d��U�Mrb�S�������ĸvT]).��W��i^dY3���vZ��;8]��K_Wu�i�=-��/�)�"�_JTP���kq/�<<��x{��������k��(��HO3g�'���o*��j�Z��J���䕡��d�zp���S^l���!`�� �+�d���;���}��rږ��q�i��p8I圠%�w�YAmmjX+��OovFS��g5ѽ�3���٦�����_;�˟uk�V�>���Os�B�򗏔 �4P��qPW�N����\4�a`۲OŽ7EY�Kt��]�)�ýu�a� �_`�B��y*�}��{X)�%җ�Q]��=/6�o*X�.��S/`� �����[ڟe����"5v�_'��w;�U�F�����Ի��U��S.F�/An�׫�����w�6��`Vթ�W,V�
�@Ƿ&�i��m5��9���Jv/_+Rn����4]�dѻ����\��Z0fۿ�g㫈�ۖ6NN�XC���r���T	��7����c���%�k(��UX�ju��Cw�U��'C)�U�Y5/4�QۭF`��P�,�XZ��@�B��]w*�	e�*�]�v�X1�[V:�ԥ����J^`Cw.a2���>]H��Q�Ӳ�+e�ܒ7!�8�_�C�Ve����cp,���+8-l_�j�`�+شuY
�ͩ���5�:0-s�g��{g;��[��Sj���0�Y�d��4(e��Ǻ�9ڝ;��0��W�0�ll٢	���;�����[3_���c�ۊX%>�k��e��4�+Cev&ҝ�v�b�|
[x6�c`k�]]Y�]�0��0�|hZM��鷣�Dt.X���!t�
.t�s]ۍ�ioXհ�w��#h��'���$b�[F�t����-v�CI�b�Y�|.�U�딨@�D��:j�K��Ⱦ"���]z:�R2}�;M�a���]��5oRʝt�"$*q�}��MM.�Y[��{Zؽ��nS#���;�	�#y�T'o���5p��B�nUݻ<)�*�,]�F�%\Tַ'9����}�m���c�������W�p��E�I�C����㠅Wb�eu�[p��J�����)��kl�]������V�����&�kY���q���s�YS�Jg-�����#�ї�⃂��iNY�h�<꧛�����վr��>�#�lލ�rp����.�TԠ�F5Y���d��n=�{
�h-F�.�#��۶O.ͤ�!�f��c��S��Z�oJ�ދ[�.���k����3z��}�4ם˙�D�:�;䉰���2�u�Γ�O�[��.��:��#;J�3�$��uh@+�΁t��ö�3�vnf2+.�F��i�k�]���nWq�1�w��cP���q�84���;*;�R-�:�A�Q-�`ᅞ_7ƬL��C�WoW:s,�ܾ��9�VnM�le���H�X r,��Lc�g�R�⮍��U�p�#�)���\�`�b����W�O�9G��`v�{B���G>QY養�_,����ѣf�#[N�Y},���g9Y�}V�ui���W)�lk��N�A�g��H��a�U{���ܪ���3l�����S::�x��^���v��M��b�^ic*����h?�ٺ9����s�T�B�鼶�.�m�Ќ7tO#!�Ή�q�,���Xהu�[���In�k���mI�is��9��cm ����A����(��VH�ؽ�ͼ9��E��E�O�Ӯ�w��u�v]	Ϯ��0s���dCz��� <U|�K!�Z �n��p�A�\��K�� ��j��0�0\k V�W��W�gwf�
�;I�9*��aꆻ�R����$�N.�2�8-�}P�Ǜ{�iqz�=�����
\��t��I]����W�N/��ef3B>���i�r�¶�N<p�%�����N���{�X�^���f��:ޗ��9��5��&�
�RL��↘����8�$��y���.�
j��ĭJ�<p�	I���u^'Ga��X�4�eD{����XXU��;��]dC�I��P���i�gpÕ`�p��8����OI�Ve�T\����o�L�6���i��`��=ړ���NA��!�9������M��ɕp�p,�B�#���ˬ�6朡`K[�ʹ�NN��Qf���6�ۋw5ܝ%J��5��q�䡤�.�K&�^h����M������2%yG�@�1uj��"
u���0��+��=B�t����X��`ɎJTT���Xݦ+�S�8By���Rt���݀K�"�e�����ns}p��`�TQ���U5/���3��W,5�w���{�:�h������&�m�X�2�v��̮��v�wM��;�le�t�Fh�ώ02l.s�{O\��b{3
ؓ���vW2&� �)Fe%��=���WQM�Q:��:n1,@�nл��]nV�2یb���
�<B�W"6~;]��cR�2Y�rc�U�X�=;BL�8Uh���Q����쒗�)_w��V,Va�,�U�d|㮺M�'�\B���Į���0:�n�g�@�]�����`k#�:���}���rͱ��*�v�]U���8=��	bw6p�b��t,
pݨ,t]]ɖys�V�KS[���NG5H��rD'�X5�j��3A#0�y`��ض���F���$��j�0<���ev3aid.����WU�lN��T���L;֘7�GPC�!����ziɸ�5�[��OgGh�v,,'��t�n�y��ň,��v�U�y8l:R�:�[�m�J��
�F�_c�������z��A�c�-��ξ�ggn$�e�i�]�{��H�۹a�uN�\ݦf 6���3ݹ��T¨�%u4���/5KK�1o0.8�ٺ�����f��RPS���-a|�|6q�w��FѦ�.�&����9� ��X�ƨ����8�2�,�A-���T}�L�O&�%��T�:�7J� L+����Ĕ��ٍ)��5�yP<hX��c̨����k��J�Xq���v��voqZѮd��կ��|�s�;�t�+2����p�=�uiL��)X�&v�V���Օ����WŬ��n�#R$�y��[Z����K�E��Vd�v��8� :�^1`JB��܎w�pG��w�U;�"m.���;�½z��]�y���'n@�U��"�B0|�j^�I�]e��M[� ��dۧ��Ni���lYvc���x)�^|)D-boE9-ܣ����n�L�\��׍RQ�B��x���gRb(.t;s�$񮮆;�7\a��#+4�m7�TA(�iҠ@�ǚ�}��p����)l�ܛ��zr�%�L�\���m��r�m&������jJ!�>E�K�x&�aOyV��{*Y��ܳ��;��n�To&B,�^O�Ԡ|j7|dQ�,�����'M�*��7xn�nf̤*ȁϺ�r���Q�z���N� �4]3�+��뙍Y|3]�Ƴ�A>S�LϴC(q�i��g�Šk�8o@C���S���mM��V�8U#S(|F`A������7z���Í��bu��[jocyY�&~к�u�a�C�Zn�U"��[���E��u��e��Ǎ]�]z�|�Mn�.��4U�V�y�*�u��Ϲ�Z5��QB�6���喉#����w�aG�8Nu�m�lC���ޠ���wc����n����8��/X� 6�t2�*9���5��uyS�HU������ۘ�q�j.X�F@N��C�Ca�=��6[�ޮ)������7eZ�:�w/��z�Z��鮜Ƞ>��K����
��WD���v]��9�Yȁݫ���Bن�0�q�
w,,���vY��y��W��vБ�R(�_/�!�/�N��y]�ܮ�9�:�)�{���6���]wdѮýul�w|�� Z;��^�r����Q��v�Э���Jۗ!i$n�RV:�0�6M�7c\wӲ�]GN�X*�c#�p^�睂��ޮD��D�P��-���T�)�C��ϸ�����l�ϖ�Y�(!Y+gT����<��z�ͺ9����E�|�����^�4譈�M�C�Ӝe�𲦧jK
��:�%_Y;;/e�sT�ÊBcf��DS@������y�惣J��!��L�͢tSU�Q�a��W#����6먐�Ngj�h4�3G�M������mM�z�F��_[�$�������S�s�Q/�TQ�;؎�ENu��ܽs5@3LFM����Z�"��������۾|c�A��퉼�����Lv��e����Mܘ���gkYShR�ݢ/�c�9�8pt��`b��(��tk����5ufuD,�Vl����t+�8�!\[��lᛧB#B����o��i)�{zm*9P��]! �F��Gm ���T��nЩ��vʉve�
��*�Ƀ��k8c����|��)8e +_[Y|�:�v�F/�f
���'J��C��ݵ��w28a��Q�XM=7!mv�}Rb�*��4٬;i�GC4%{gOe�u��w]�ŵW�S���NF�+3n�,�e0��)�xkhV�lR��\�|j�z�բ�-N��-����&m��7m+c��6]�P���խ̖��⯱����;9�)��y�%sZs�����ѷD���,��{ǥ4ܮ
 v�֊���� �9�mu�
��Yعk��9ے�7�7%�(x��v�|�|��5Nآ�m�W�l�'���&ܻ��I�ۃ�q̝ʄ�p��rp��pB��'b���	u���+�{�z��9����ws���:e�c����(�EP���}�������Z$�̠�r��&h��w��V!��b@Wt̠�qtZc���.�mc���ڂ��B�1Y��a�*�����B[3���-���X��P�AL]7,���������Ev�y��N�VCx�������N��i_�Q*�ڡV��J*��r��tW���B���j��&�u��v<3yki�"���(�
�䨝�ll�k�7��Xk����s2;"��+��D'W�q�����'g:�<�,Xs��7��rR���a���2�pԸn�MTq�x�9� %��-�}ͫ��[�������θt��fW5y����m^�Hs�k�^1�`j�gk�77S��*:0��{��Vb$�p86�6�'O]�2�@b
�&agX��8xkcqt�}�yV�Cy��YG9:����T�V��J��Q�qf��ߟ^Tٍ�۠�b�ëw��&C�#W��@K�[p��T8�F��(+������Y|��n8I7e�:+�Vz��E*]�x�]�fk���k��'H/8.�
ğEM.�R�.o�N^���zW���R�U��;3m���v�oo&g>��&���t�UA-wCg>�Y`�Mn��� Z�MU��^�6�C9,�gb������]��w&�ʒ��/m��-O*E��,U�u�痄WetӮ�t�0a�[�1�sU���z�i�9G;��uv�(�7,q�%j�̫Qu�Ү��֑���Ǩ� U��0�A`��̹��¡�RO����۱y��rݦ�mJ��G����m����ͭb�h.��qg"*��tR�f3Fɝ�

)��oa����wmڔ�n�+���J��wX�u�0j��e՞n�7LZM칢h�q�ӹ�̻,�(_%�I�����2n�>K-e:i��G�(yPǴ�F��\��|�n�c��=�{-�D�:RX�]e:�0b"��9���f��4m*Fm�TwO�*���=�_K!�ŕ��aA�X�]7 *�Z="_V]ַ�q��0A�TM��]�ۭ"Z������	�7�K6�M�C�����Jܫ�X�X nڝ&}�.��EZ�X+�Y!��Y�}Yy��������q�v��V�)JY���r�ܹ�tS3��[(�0>�Gi���+y �����m��0��B�P�/�l�+�:H��t�*\üz�X��S���iX���hs<�J�������ܖ'�j��#��M�N��WwB�*ۦ�v�B��ÜH�F��EG.X5�j�J`Swr^5PY�Wwu�W�킡}�r#]}Ir���ʌ�����a� �9!LTM��+�7�9�*�%D�a�2�&��
������.��u��l��������4��2Vwm�.Lr�����[[��RWXr��fVA���I�����S�K�Ce��{��2�U��UҭԜ����h�̮�\�}Ό�k!�`��6�3Vb1�555Υs�w9���c�����j���y&��P��e�ř��k�9R.Y��5&k�J��2@�{yqr�η{�\�e��sl���r�[����S
\�U��ʎ�f��P��/�Zѽ5.��ק���J�h��j���w�!/qB��]d�&�Ϥ`��ئiw��E-�_�Nj��#�E;��Ґ��w'����μ�2��E)pH4��&L����.Eخ�Em�Y�k�s�j֏�Lș�R�ebj�a*���v�ԦU+��Tn6�Ju� ���g�/6��xh����Q�����!]�X�ܳ�NǼP�+�
7oc�����O�����\����t��z��s/��A�N���m���M�D�l��Zx^Q�������S罂vee�Ż; �:�&����%ֺ�{V��T�9�t�+�Ye�,b�W`*��U��[B��Ư�Ơq�!�a'H9(%\�̳K%q�;�i�WS�LKwsO��em�*.�=���d�'��B��]�3@[g���`dQ=�h�x��{U�ô�Pb�銓0v+�P�Ѭܖ�d�����UwS�6r	�5\{�ι(�^1��)�vn��� ��auq9��O�����˷Pq#��]l7s7	z/�C�!�P�6�0J�m�6e�EE�U�ΑQp*"�nr"����{ξ	��e!ٹ�x����X�o-�|�4.5��P�t�o"F\=��S�́}�*Z�Bk%3�N�ۏ��V<}]���^��2���9V���<��T�G�ـ=�����L|�_��}��V�5z
wۼ��5mp6�IӺ�����*]��Y���P����V�xr�����'�������#�]�\�C��T��u���n�Y֥s�^T�������fa�/����ŋ��D�%�S�W|�G�D�a��O � �ma[�uW`��}���f`Q��j��$xq���͹��9]m�c*�.�-�����:���.�
ӻ��#��k���1�!9�8�O�=�`�l��8�Tu�9� b�!Z��PϻC<M���s���[�1<;�Ra���Q[ڌ�U�h�Gn�p{:+]6�R4�]�E��ղ�[cb��¸��d#��@�}�9���k]�w��/Aʶ�u���3�q���F�ep�.��ΕB�t��j�p�兘)ǃo�>�Uv�'�XoF�,��\��6�iJ)W%*����w�Z���]f6.Z���2%+���b���u�.����R:�O'l�Ċ=�F�m�#�[����G8�`م��L˜ZT��됳(̙�݇VARs�{����e	�t��'9)���V���3��.�O4���	fd�9����L64��$�;Fi��#����)�JRa�2������!C&u�Wu��s�:�wk����;�vH.�Ѓs�; C 4i3$ƂH��"E�B$��cnn�F[�\Sf2B0�%b;�n�� �&��� `l�d�l`G8��;�h!��2��3�D���l!�2 �.�[���Id��bL�"iwt�wvr��#iLIwk�F 2X���,�.]$H�JJh�$�s���1�ٍL��Twndh��a�Y Ƀ��PX�X"Ā�dLi2�� ���ad����(P � J�;,^N���;/J�������t�_�qw6���h-�1L�}I>�T���^�]��X9�il�[��{��*�r��nv#�*�Ψ�]�	�|��WZĶ�ӧ9��ݭP�G������s����ٷ��}C�(���������_�����:p|)Z#n���yѫȰ����o.��0<���
����	�ؕ��b��B���Q�\����>:Қ=@0�+�j��=��f�~{j�nd="�b�;5;_��i���6hiD��B��Z��tR�mNA��z�u�#4��x��T�+q,1�;�S�w<�\og+�h��?p����?_��t�]�-8��R��á�8��T_�%��&��F�4�ђ��N��[��H�7�m��fz�G<��Cd�B��|N
���Z]m��K8�C�cd�"���*�l�Wn�U��{��7�1ŉ�^���hd������4eW�H|kHBHܬ,���L�6��ĮK������5nF{"�����-K��Ю�lwʈ�C�
I���CJ�ـm��W�0/:���{bA��-��9�_����k�:.q���6�QB����=6{��ކ�(�:˷v�i�ikbf1�vi:�z�V�Q$Sn�NwxT]�����t��t�k�[���:(Vjsw�?aNV�B��#�V��Rh���0h��{�*�ʷ��gW���|X�U�o�����s��
Ŕ^C{b��|&�,UU>9-.��Ȼ���9��Nχ�{�Z���:ԝ=`d��9��-rQ�#y糈݆Mfl͒�pE�DD'n��u)̎��']%�~�w��p']��z�N���>�[��$�;i����\�G�P���(_0��T��Y��`�_	^�695J�H�l��L^��oҼ��|��c�@-򸚃LO�~|Y�B]���g��fϼ��]_r�"õ)5J���k=�����{�.�Y���t�K�w�:�G��s���Ҹ�9諱F��W*���U9~o�	��2m�Q�C���(��!�%G�T<��>8$󜀶	�8ƴ���{܇���XX��Df��&��B�YG}��=#��rsv�6z��G6T�
�i�b��$n�{f�!�<�5)���Q�{>��x�6a[�JǼ�'�Т�с-e�b����6��O���*C�� �gZ���!�yg`�/\�fc4�'D�uo0�ɭK��dטڶ��\���EV�s�Ҋ�:Iw�ۤG M�j�x��������qv��Z
��|�#!7yS,�]w%(kyw/泳(�S�dΫi���8Qed��!���sn濃�a�Jy���n��N�QOpR���i��Q����3A�.�5�,��u�B���BE�5Z��,�'Et�l��k2��k�����b����D�窟vˣ���eLxE
,�������T����̱x\au�����_fv��b:K[<�����_�a�
(��;{$�$�:��/j��7j��l�K.�Uk��']F�Y2w"HkgʆJ��aL�y
n��TgG�j�L�eD+��-[��v�ڼe�#b�����>4�ʴ�ǯXt�09��mX}�V�닀��3S}x��sL�כt�vI2�3� �\����tL_�K��e4F�p��.���.���Q|�Bj!oђtЏr�"@)V�d�+�tZ{B_���|v���~̱4M:��	��T�%q3LaL�48�B"} 4�`���I����>W�5�����4]v�+Td�G���󝬃c͹�O�݊O�H���ڡ4�㢝!�+OG�(�k�{���v�j)^ZF"<D���tl'#�8�9�d�F�"��EG��o��b��Z�{+�n�����F�
&��P���SÞ��+�'fM�9]�C��I����
���.2�T8nm�H�=�}���IP���zk`I�sK�e�/)6
�FｗAы����>�uv�uӤ{I�4�]E>-�{Y�V㝛���r&VV"@�J�=n�i@iX����j�qv2��<=���r,O�����Pt�^�k�N�.�|�ފ��L��u��?u���J�9'���/|���Lŏ���e�E��ހrǾY�;meH~�l|�8+�@}���l\ed��2�v'P��e�O�?��O�zD�ͼ��Ӳ���cB�Y�m�xώc��;~�)�V*��Jf��q�U:�l�X�9o
�tr�K��wF��9p�{B�V���
�د�j�c ���*��6g�qz��f/ MT1�N����J������ �X{�l��.�	}��wruڃ��M�7��9���]P��.!-4��T�#�z�u�BNA����FZPm
�N�[�*U�83Ǣ�L���P��3/iw��(�ΡN��dg�F��J�L�O�{�o��w���x�� ��>3���S=��U]%wl6�{�rnש��!�@�Owna�2���\���,�u$�>!�
��G�ݗbY�Z}�*xd�
�/�5�N�mFLi	���i��Si���%W� 3S����9U![�W���]u��3����3�խ^�N�/3KJgz�Ik��Lˍn���-�xս*O{�.��z�K�U�7�E��\��ѐ{�g���W��u���h<�(�\w�S�7��2�J.�����F�"���=����ک���_nr�盫��+���+q��� ���WN<�1���u��K�P���8�8ܘVݘ��ѤL8��3�J�&��q!����kP㶨�Ǡ=#���Ѽ%;l��ґ@9��+ͺ����ЦJ4I�����i������:N�/H�Ƚ�Ł[!FX�*���\��(��,���V�	T�J�%�������ܮ�-eft����EzNÓ0����P�jW0���O��*d�f\G>�x��[כ]q��=����bm �I܃1�l�(J��9D8ɬ�
{y���]�N�o�μ�qx���wf�;�U|����?���~�.�ڃ���0ǋ��u)KcF!���[�r�/0]-��.z7��ku���P�m��q~��g/�8e�g�'ʦ��bU�%'���^I�E���o��;��>?̯0,4�s+G;�U�hf��ѿiD��B�u��3�p��I�ьʌu.��%NXΥCq�1�;ʜ����U���1}�R.��oJ�y˧n�.�]�1q6gJ���(��]4u4��ן�vߟׅ04z����׬h~:M��+�Ŭ"��hc�e�}f�U�:s
���=�(�o]�0_�R�ic�/㵁��_Z<��p�TW�rć`ά֌��`4c�
{�WL
�ae@Fe��,a��3h�w��uF� �:W[�֪.mY�p��Dj�9�b�7��9Z����g�$��x�)�K��C�cd�b��Fw��4.1�F��4�f�}��4m�/d��m�2E��$o�����5�5�!��L<9�[�t��Uí��n�F/kQl���{a�.Z����
ɥ\pq��*�]\~�b��F'j�ɂ6�ns3���\c5A�o�s�#`(�:.q�"ࣨ��8��/�n�BS�ٺ�uZ�
�g��UI����=�]�Z'�d��PuA@W%4�=h�O��ڔ�W�s#�3�� ��pqP8buѱ�[G�~/:��l��?�2�J�\Y�-��R��6����¸����ht��y|h%`j�cb�&�FyˤH¨�I*7������i�pN���=���ȑ����1"VӣtW�޿8Ԍ��V�IQL����SҐ�%��P^}�� �>�V��Z�%�w�:�T{��x�%^r���&v����Cl������LP�<ɓm����o�Y&GHG��9*<⡓G��y��� ���f)��gJ��%��>��k֪�~T�騌yaZ�ũ�/��b���F�
�8�Q*r�p�����N�����t��;(
E�c\������D���ܖ@��s[Bt�Yn3�p�q��k*niN�]aV��p��M���B�^�,,	;�Fs�K�]@��ޙ��*ΊK�����W������ܲ
�k!C�GaȞS����w�Q���:}�5:�E�s��� �Kq�dckܢ{~�c�A���PsrCӾ%FA��u����A�A֩�k`Y�/6v��k�V��썲����j�9�����>��QU�Ox�}ws�3���x���C����+=ʑt�|���׾�{,��mh��
�;C�S�F�\�ќ�|2�B}�,@�fU�+�x�R��(�k��e��w��}��%{�p�1S&�:<�%�cǷx�k����n��er�-TI��}�R�eD#�S-������zCj�@~��9e�vW�}s���~��2*g���K�4��+��aҌ��B:ڠ��>J$Dh��Pyv�&T� �=Ug�6�$3�]�V��zS�*\d5r�	��==����x]	�:�fO[2:������(�o`2� �ZM��efB�tb}BKt62�\�̣��`��g+^-U0L���%����7Ż��R�a�Ux:�g*n4�,�k�G��n��>���sWR����ǳMݠ�n�qm_]��5Y�-c�w��i��y����c�#������>8o��W�u\Z��N<\B��w�\�P���}�*pq��G��l
��$�\TF�0��U}ݴ�r.L��u�������`�{�@���Ru��ִ{T�j�_xK��6�@�y*J���'���3��&=�y���$m{�[�i��4�|���6���M��f�ڜRv�ݓY�g�y1e��{+�/~�~B�L���4�T�^i;2l' k�h`���0F����Ѝ&����pﯳ�o��^�V'���X���6O�wy�4w��r�	s�=��S}I�&�c:�`ה�v�d��"wO�K��~���{��0Anׄ�7�O��H�[�xm��{���+�ez�5b��L?�ƅ?��7^�p����e4d��.3�ҙ��
؁����Rv����C���M��8U0s[�h���u,�
��s���eV����V'�q9s��I�[�L��8[�E��<
��,��5�ڿu��qN���ٲxM�I�ۭ�y��{�9��o�九��cگ�+�Y�x�8*H�T���
��.e[��<@�E{6݂Puxz]�/�[�u����g�e�1C�s��p9���T�&0���EsN'�Z��r�՛�春�.��`۬���I:�C`���Hѡ�{�FM��2�+��[�ֹm^s�p��y;{g#�t������<�a�7:sL�Z�r�+����[��Jo�*?QPG_��F��5���P�ua��"��J�-��N��6a�^���>�~@ Q�O[Xd4b?{�:�O�[�L�JUP9in�0>�
2Ҟ�����c׈�/v6�:��_�Iw=Y(�i'�2<��te#�;.ĳb���cjJ=D�O�2{�v�8=��O��O��I��0�u���#�*��
�8j������ƾ��ج.�;K����;Ny�06�mٌ���3�v� =W�2�ε���w_Ma>���T������S���M�H�r2y�Br�ݳQaL�}%,��fs7s�l.ż�c���I�sQb��`q�
���]nCj�,1h��|W]���5�J�I��U\��,a�%�GvP[f�#�ȡ�i]^����k^iK%�]]s���m.'���wVVtEs�"$tC'p3��J��3������p�,��;X��=7Z��TD(�����5~.ϢGK'�A��jz�n���ţ���t2�j/���Ζ�|�
݈%M^�7�5��`Ī�i4�u/���;\�St3��e1]588�U(�QcG�+ad���3����whOzq�|c�t�y'�օrbK���yԋ�Q����)��x�uMa�Rn2�}S�[��PP�r���i�ա.!Y����`��U~y9l4���QM�5
�{w���YD�ܸ���D����y�m���G/��)�x绥3�N��
d="�LW2�s�l�ҠT9�rm�m�˭Q��t����(�1LF�C����ɼΥ[�`p�]�NqԦ�7Uo�L�x4/e-�ވ��j��X�#�U���U�����(�`xK5�M砍O���l󨅕;Y��cfs;��+�����_ѫ)�ʝ4=��C~'u'NҘ��5P�d6L,���.�-��{KZ8�d�~�l�\_g3�C�m�� c~���Uz��ƴ� �[5[b���淨�m��U�3[c.��|�e��5��m�ɣ�&��pq�� �{]u©��Y<� �]�xr��Gz��܈f����+|ps�e���
6��(�Z�]`�� h� 	�q����_��9��>�]T��)��[=9봎�����q�s!@Ro]H*�KO:����ݸx�h���P5�$2wڬqP8buѰ[U�;�Q���1�=��J����
&�n�c:dE��(��mXm��2������8��u*�W҉��t%ӌ��9�����)-|n���ύ"�1�s_T�m9����quҼ���X�����9�{5�S�U����!�*e�t4�#0&wP��.(���͏M���[�6��1p��v@��;�5�:��qptj�� tU������ջ��|B�z�u\5p��\�:I����&�ySCə����4�gX�v��a
�ӓ���H'�[c+uoƓ�G��+�*շB��//Ω�oA�;����՛v�f���,9������'�_�o�ܮb�X��9�;1J�+ck�v�o����f�RSS��p�F�ky�b��B���wa�E����)1Y�Κ{]��-6Fm�����T��n�N����+K��@��jsk@VS��Vuط�F�;�҂O�;�P����&�3��}0ȝ��3x^�bGa��naгx��N���[��?#�.�FnB�jl��d�΍7�R�e3�g^�3��<5�'�Wk�S�����P�=qn�v+ߚd���<��pu�c�Mh���:�JKk�޵��d�M�ʞu�Z$nnVMg|���U	���łVZ5mS��8U��*-���]]Z1]�.ǜ� ���]�C�ZdY��,�9Da0�X�@8��zu{(v�6� � (e��n�z��.R�s+a}{H"&����Ϗe��'���}�b��</�a�y��G<�-eu<�{��]9�kk/� ��܋F��yAp��[���j@�;������1��L��&������f����h��+n'{G-�`�(���1Z�,+�Y���*vr8�#s&�C���8��V�u<����ri��j���,��]�gu�lɶ�~T�h(�f���zVk7���xi]H��Eա��\R��K3�ۼ��Z��Ŋ!<k���[ur���Jݻ��'{�N�%� _,V��e����O�3VKt	P�
�Ihh'����M�+�f�[��upu�*Y�ь�LȐU0��@�6j	S�C�Y��e:�����n��H�}i��5�x�+մ(��KC]H�Zy��7VT���[��(ېf�M�uRW��U�F��A�f��K�I�y���+][�쪉�VG>=S�f�n�1��3z�v")���J��:�t���7�uN��_.�5��l&u9��]�w��}׫�I��WֻuR`}��9a��	n�ࢂFVm�h31�:;:;�Vbʹ�-�wp�-{y��Ù�xȚy_Y�p����Jo7i>]�w&p[�����vS�,��Y��}�2ED*��{��1��C����;h,����'��J�dء�u:T�P�e;��p�5�d�E�f�Ic��v�t�Ң��e98�*V0
����a�6�v������9�%�-�#�ۮ�������E��f\�[�k�P�����a�&�ܒ!�DCI�)2"&Hl����!	�I2��	�d01�Ia%��v�1JL�gwDd��e	H���Dc;�YE(�3)DdDT��M	!���fJh	�ID$�03H��sv@�`�2)F&�	LRd��J���� ɚ��2R� R���L����Y2c$hb��DTd1DD�61.�h����0�#�&bE��B���щ�سa$��i&	�"��Q�1����4"�3EE����33�C� ����J��K����OWQݷO#G��a��뎶ze����Eu��c��{a�	��x����U��{\q��l5���]#���3s�R�����������潾���^�v�Er������v����W����m��h�z���m����^+��[�~��o�������=1� t?��qq��+%ZK4`I��.���t��?
�(��x-�y�-�W?[x��|��ݯm�ۻ��~>�kF��|�<�}x�_ˆ��>ux�^u��םk�������k��׋~^��o���꽷�����A����L��5�Ҳ2~��xE��?W��6���W��m�v����K}W76�����~+�7�=u�o������ǧ��=�xۖ���ߝ5Q�"<+�\�p�� �'�♹;��ɉ�kwǯ�$}�#G�"0DX���S�*<�����( xDDxg�:�ޕ�^�>y����^/�x����o��\�/���w�-�oj�~��v�~v�/�W�zZ|�/K��ͽ*��hi��
#�w�a���}��}g�ϼ��/մ=�����;�߯��������_�ϟ}_�~>+ţ���׭����x����z�����H�@���Ǿ��M�&"gه7����{k)
��Dx}�y��]��->u�������ܫ�{�]}m�x��ܽ�~y_U��������<*� c���u]�x���	���B��Z7�Ͼm�����ޯ��������t��䪣�oϼ��.(}C�}�z�_潯K����7��^/�߾y^��}k�w��_�x���羽�>���Ls2�c���0j�d5ssn��}�騷�r���[}y�ֹ��]�����ve��v��!Z+�01�}���齶�W���~���潍F�4��d�*���Q�	�L�d�zZ7��ǽ�_[⽭��u����]T�L�} L	���0 px�0�#��>	�u+����U�&�+]���H�"!�UX��">��:�������|�zU��_���5�����5�+��m�~׾�[�x�o�w��7���-�x��:�߫�ѿ����<*1�(}̣����Ϟh�iL��lE��}��^j���77���Ͼ���o���|�zo�{o>�����A}m��wޯ�x����߷ߞW��so��^������ۿ/�-��Ox��;i�� � >�ܧݣ MȮ��7�1�M�	�ɾ�,
D�S�g�+3�k���,�RT��+�&'9����^4�r���J�$]7�9/�]�X�]��h��){Y�)^����!�{�nXnf
�x����]���2�XC�6�va��t�i�*�<�gv������c�<>�*����T|���޻�����m��o���|�^��n�~^|�Ƽ_����{W��}k���^��}W��_���������x��D�ǽ0#�{{/#Y?;�9"��W�zk�sz\��l[�ݿʯ��$L{�:<=cn��(�P=�Ԁ*<<`W���[|U{�|�E�o���_Ϳ�܅���4�0A5�H�S��H!��ޛ�^-^��~����[�޷��x��{�ޕ}\�5���6�o0.H��{�ǆ,��.�Q�=���7�nU�w�;;�7�no߿<��{��!��,C�:�z�u�r}|���wh���(��K�Y=0=�1a} d{��������5��[�u_���o;���ln^�{~��x����Ly|}�d{c|\��xDyG�lk�ǔ�<"���y�NV=b&�~�q[�i�z�������6�����6�x�濾u�o�s���ϻ��^��\�^ﾼ׵�:�7���׮����W����wu�<`�Z+�޾|��߭�η�ux��^b>��;�`�V�έ�o��u��@H�������W���|�ޟ�+��wڟ�A�C}8�#DX��1�号���������^��k����z^�x��Z���[���<�ƍ͹o�����[���|��x�r�|	�<�f���`x�d�	�(���t�`L�ti��G��\1�0?��{�\��r����_�o��x��wkү��~/���-�����[��߰&=�7��N����x>�@���v�����*�������szm�}�������X�>�@�tLg/��<{����\׶��Z=����������D Dh�<�~�@���Cq�!�)��饞�=9T�}"�}"��H��W���m��׻���KF�W��y������������6������/�����;>� c�ޱ�(d�� �7�{�����'?}$��"�}�Bj:w���s{�s���?1�x�=10>�sP<"�[�����zm�u{�u�7��^/֏��h����۽y~��^-�]}[�lxl1ᖧ ��G�xh	H� } Ǻ=㑷^�����zRy�g�/�fkG�H����D������"zvN��ች���Jߎgbs��V �n��&���N>}ֲ�3D�:5����.��2;�i
�I�u�n�0�WU��*b�k��4�F�s��M�aa��R��iFK�cG8jC���wr�Ԓ
v�]%W��Nr�����sQo��~z�k�|y����7�ܾ-������|�M�nW���k�{k�\5������������Z��������~�kF�����7����o��ך�F�#����ݖ 6br��r�c��=��{r�޸ 8<"f|&�x����痵}[���������ߊ��������[r��~/So��w�^�����7�v�[�{x��y��Ea�������������D�XG��?Z�okƯ����M���Ƽ}W����Q�D�19 �����q������^~��-��m��_�߾W�~-���������W��=�����ͺ�R �@���&=���>��}_n��R�*~��� 1���"�TDx���5
=�:G���܏�޲}�
@:�z��wu�?7��b�U���-����ۤ�-����	�����@0<"=�:���l �	���Fw+����L0{��~͹������C�b��Q?|,�_��{��zU�s~5���o��-�]dT{��1�"=u�� \�d{GL�齶��o���}~4h�۞���4_Qc�C� ����#�!����n��m�/�^vb]�~Q����c� d����^-�����om�+ƿ/�׃\�[��yش����;�ͽ*����Q�P(��<0��0�<b��[u��A�t���"��>�����|�.r}�r�i٘_�Dd���`��Sbܮ��W��Qo�������u�o�_��/|����k��^>7�;��lE�u�+ŧ�׿}xޞp�zaG��-��#����pW�g-Mη���[s"���DH�� !�믾�c�����������Z�����W���߯z�m�oJ���}����E�}ί��^|�^�鹷wm��^���U�!�Ę�&��� }��i��I�jvڒ�>8b$}��<�\}}��&�������3��
 P�O�z���k�^���kם\���>��o`�1�p�$�������Ȩ�G�d����@ ǽ�(��9��ܬY]zg٨Z��|G�D?��,} }�9o��x�ƸwT[��^ z�Z#�ǔ���d��	���_��|o��|���^�����~��PW���U��Ub�~|�UAG �b����/� ��.(���^�o�?wR���x�J���Ê�V������0�Ih�q���W#�onA�h1'}�b^�˹����G0H��d�1�r\-�8�hP�H��.��g#�9��k��](I�;��f���&�cql���uB,كej7�$����嫦=���?����K���7������^-��׻��^��\���?��o�齶�����7����)���Ͻ��zb#�Dty>����.X����$|�H�0��}��!>�o^�n�[��ݼ�iG�?�Z����{_U�i뷻�W��^�����ݽ/KF����w^����x�X������@�>��{����-W���o����_��-�\}��oK�� ��/g2�|^�����[z\P����L	G������=�O���ۙ0<"=��w^��_^ش�����<��U�y�s|_���-�^�y5�~��^5����o�s�ץ�����Z|�#��z�[����g.�,�=C%F����{�������z`{�����<�����K}W.m������M�/���W��ƍ�꿻z[��x���|_����o=��|������?<*�T�3��Q���{t��S3�1���ju���[ʨ����X!��.9u^A��_w����]�	��2����˥O��wKg��{��H��̭�%����7����-���ǝ�N��Bjx�T-X�6��Ai�nU��ۍ`q���S�wUq�]ҥN�̒���;�IC���g}yS����!+�x7�>/��5�M砌�_����C^ݒ��&�w�ug�7=>�/}�D�ƴʇ��J+��\ςӏ���/�\6���Q]��3ؒ���b�a���Om�p:�.�vJ��.�C$XI�����W��=��R��9�t��.��J�㐋H+٤7ַn��a�r)���6����4	�i�-r��)j�ض����]�k�8p��ӹ4s�t�E�f�������鯺�fc
;W�e��1A,�X3{ncc�!����k+l�e��ŹW�r4�8�?��U|�w��t��k(?��x8�zpi��l���N8�����iq�I��\�������!˯x�~�g�ia���P�t7K	��{M�e��F�ΰ�˜e��b�9�z��pݍ��:mY��p	8�~ϫ��9M׌6z.7���GCRt������r�f���sk��E?��^�#]�b�b�<�s=*buѱ�ڿ\;�Q�aq/Ke�i	[�3ı��Xe��q��V�C��XM%�z���x�J�X1������4�.*&�chV(�IC�L�l��M�lE�v&��#��4ɉ�����7m�WLh2�V��b�T^z�F�[t�����8��P.!L�:iL�A��q��Ξ�;0ߓ3�&�.��۞��/��ӟ_�6�b�O2d��#Z�:���I��Ni���M>�1q�o�G-lFh�P�f�����Fz�y\���r����5ϙ5nP����	-Ŷ�61!����Y��$Va�9�vV9���g=$Xݕ�j2_*}�S��+y�P��-�q�=y+//r���ꔮ�
��2������W����Y���r��&�����Κ��rמ���W�`p����قQ�E�Vy�$���3���e�[Õ�YZ�Wm�\�]o�p�B���=��Z%��X��9�Yz� R�=����(�����G����8��^����a�s'�}�ٮ�5^�w���*�+������i.H�X�:%��퓲��ٶ�O�~�Zw,��/�(��#ܾ,�i.�;���<�yg�U�k5b�1aӠ�,���z*o�藫�L��OB*�~~Tm��R&�p!��3p��,B�K,��2�}n������
(gNI�>��4/B��2�[���}��,g�%�;�Y��0�:�_k����e�ٰ��V
n��TgF�\�˽y��հ�}O]QZ�)-z%VH��i0tbv�׬:Q��"Ԫb6�-��/;�f�B�;�.��1$�*!P;��|��϶GKҟu�B.^<���~�ɺ�;%������`B�,a���y%�� �B$�ZM�y��C�����-�Jyf����uk���aC.���n�8���fJ�*k�D"& ��l&��.U��m��Ե�m�'��~���c�^�N�0��l�9Yǽ�MW��I�$O��+��g�:R�(��W��x����^Vp���u����\F/j�]�=v�����8{�7���Ӊ���vL]xP;-<�Z��>�4����&*���볚�<�	��|k����.�ht��`�oM�Lv�;�G�����tmF��G��kvE�U��]�5��ﾪ�ey�S����������|��w����]NGC�M2_#[�"c����`����&��{EQJ��K�x ǆ���Zlo:�v碤��Iٓ~N@�j�����b/��֑]\�	�=�I����>ڂ삺E�zT�5~9
6��'���v�^d��7�Ϗ�o���� %��U*��h����j�ePY���s�lWJ��<;���4B;a�bլn�b秡��R�x�C3`��S�mȨ��c��@��2�c��;~�+y欷���IQ��t�巛F���g�g��������|W;�y�lj�/K�d@�gr�&epI�ݤ��&����D�J<6d	�XxM&Y;Dj<گo{�oY�*	���5�,��ιV-����6�=�q.�T�V��W.��x�*�N���a��!��A��\+t@���K�9�=��i{K�DV0�G��7���mj��]�����|mӧ	d�gAvT�P"7�(�|%SKt���]͊��i=}��܇ޑ����%�3��X�4�:ݙ�	�.�ئ��Y�GG���4}�J�;��mMB�,�kx�teK�T���+�up���
B�v|%JjՄ.�����ov�M����满k$���z{޾�^�X,�? �
�i�=mD_n�}�$(��!ku燥et,2J4�U|B�2��뀹A��ܗy����:�T&�[>����s�dm��ai{�1�����A�{�5b<p��+��e[�^�b�p�YM��\r�V&�\w�q�q�06��f1��5�)�0)8/uol��Ņ>�ex^?��|tT�5�]_kѶ��Ȉ�)��^mМ8�"�wjE$�v���[�a�,z�8_4Ek�#}�Q�R��/��VWm{�[�[VYٷW'���.D����H���SǕ�ҹ��}(-�ME��i;���;�_��O�|��}��"�}��qgޏi�q��N@�qD�z���՝5���W�f{��@X��vf�jE�+�����[}Utlaq���0��)��.ϢGK'���97
����x�W��o�cի:p}�N�斎�����!�ȘP1������_�p:�YY܅�8m�/f1�O��qx+�q<{�gr�y�L��Xi��V�w`����z�^W�l{�Ӗ8�O&��V�
]�2���u����E]:�7\�N�S*S�-�:8y,"��2[��y5c[�>em��|S���2e���y�d�8|b�|����@��X�wK<fqr�<������;}G/�Ķ:�jØ��{3���{��{7�:����0t��2�q�B�T�W�x�r�u(�q�3Ω�
��R�$��G7������x�+gӌ�T��`��tUp��x[�م��U��M��.ή��ِ���K�}�)`���C�v�o�������.=��;��ݳ]���'0;��GB��e��P�����"a�r���.�;
5�����C%TXI���TW:�}�Hຫ���ar=2����Y���.���8V��l��8앷в%�NG}]w�4�N�}����-�Jii�	�ƣ��M$���a����
6�y�C6ˁ+C����E̱�L/����l�4
n�����8,(��iIҐ\`DӺ^��z�̕lh�>Q(+=B#���5����a!��Ճ������ڠ6H��D�ح峊�������btߢ�Ϩ"!����z�Q/��n�bD;�w�:}� ���[�r�,224u��	�"}����1>�����ܕ8�k�X�Em�N��h�嬋��e]������	�T{F��2������{׶�>�s0��V�_K��Y[��@����r�c���J�&�r��Uu4����)�tč�a�Av̧�7�j�.���g���ƤX��苏�� ���4+^dGi��=�8֌�JC��n��i�GB�qR�U0�eU�x.������0��:X�T��o��n�U��gh���69>�_�U1h�&O�Ds��6�E�k��u�����<~����+�^<�)�k����_m����MW�N��^�>d׭�v� ��jʊ�v�=K"J�/��8l@�E^�AU��0_�9�5*�LLd8�ʟ`�td��*�2R��N\Q�g����6a[� ��ʬ$+�nW���XF�=w}ie�gD��t�������v2��a�|�g9��85�|��hM>&��v����Eb��v.n�N�{���	�"8 �{��~u�N>��a�]��t^t�^������9	�}Yv�������!��������6��cfX�`�Y49Je�ۿ8��)3^�]j��^��-;�W����yMh2������U6s���`R����7�岳����e�
;�Y��m*A���B���T�$#�L�tXۺt���;q��(��.��Ku����G��&M�cE��Aܦ���8��]����ƭT蚋��nmw,^�)��c�c��'�_@.�V�ck���iRǋi�Jo�ݥ��6�@r���]we �n�{��7U(��b�/+���o�TC�KBw�Wkr�c���@��Qp�h>:�9��Ρ]	��Yv��Q����iA<�|��VX��<�.Z����G��su���f��Ә�l�1�9zL��T��ǙKL�r+��T鼔&�ƯNn�iֵK-+�a_��Dͬ��{z�N`=��i�v�is<y�sl����f�YiV��*=���C^��o	c��=����]�%�}�uK	�-]�n�3�Z��ܭ��s؏�U�p5 to���õ��%���$I��r�gCksVeΓ�Q6J�Ai;α��K�W
��e7;�i_GmJ�>Sj�2�kj鋻'�+f�����!�+��}!�-�Fb��:�*ٰD�M�Qp�6�[7���b4�PWW	�.뫜@Ik�ȇZ����z��ڏ.)�y�hywF��]Y}k��{��+�50_@��q[t5�e0�R.�̼κ,�ɣ#�@�] ��=1fU�>���9����kQz�
k|������i�.*�P���ov�u�}u��Y�r�ֳ3Bt����[��J�M�||՝x�Z��dZ��AR��L������	ǲ� ��������b�((u��ܱ��G���B�9P��3.��2zefk�wy�5ϓ՝Q�e��h2���q�"ouk �t��ݜ�������R��ɴ3��F�]Pc�5w�VkJ��4w8(��\�Y��Bgו�.�����\aQ���X�![�:�N�IV�Yt��@&(�f����VNa�C䲢��t�vu�CMm�-L���m�բ"ɭ����RE^}u8ά���mdH"z��*��ȼ�ki�P�ኲU��Dqɻ��pJ*>݉�{g%����B������Zoy2{fڂ�l&U�t����I�t̽�$��pD�k���;���y�m�s�㜡��h���t��/�nv=z�Vq�,U�6C��<q�2��/��cr����M�����4mԻ�6#�0#�uW3o�驭��W�(.��V�mJ���fByKw�Y��n�t��u�j��՝�jmj��s	a��R
]���:�賜c9�d5l5�[*�������Raa�4'9t�3@�Q"�KΥh�(�o(<�ؖa���^�v%]��;��ca�<(�?݈�'�Ǵ��T��
�~�&�r�p�������nwE}��G
����5}�N�y�&�\�#��qw_=��+UU�$�#3�I�t,Ikݟ*�Kj>��2�W�)�
Ψ��&\��V�K�ɻ
j�׌Z�%i:�n�yrU�x���[$�d���ʮbӔr�d�hZ���#�w��YDû���˧v��&4,��2�����K��X�z�v�$v�s���ߴ])�6�(���XMH�Nu��IB6�f����Q�u�X4���9�H�\�,�F�N\�s�bK�`I;��-%;���r�AHY��4�"�5ʸ�fM,&#D"����%)Q�	��4E�'wB�˰�1r��DH�hC��ٍ���v�L��3IB�(1�,b4��.q
���hĖR��!�5Dn]LL�1	(e((�ܡ�P���%F]�6i���Ŕ��4�*D62ĶI"���2j��Ɠ0ɀ�5ݮX���%��%�6"�~���������z�y9�e=d��Jޠ�0��u�Ԅ!}u�P�6���p�AA�F���.|'-sJ6ܧ%�=H�c��}U�W����,^�g��u��.��X���B8I�W ��$:>U�el���tЄ5�]�]�SJ*qlZ��(�펆<�SD`���.:;v�Y���"@)V�`�ea��Ԃ�*��w"����ꍾT%�)����룉����U���#�� q����>��M�<�Yc�3o7�s�=������R�7���G���f���n�"�V@�
d�w�J����o���5�������\
���fz6S7�<H��.�F�r:�M2_#[�V#��M5�7�k�
�Z��늏�)V졮å�^:f���67�L;󞊒N���כ�m�}�u�N�#Ct�2OC'��f�vEJ�%K�VB���(�e]'N܍��jc/��*�!#
f��Mr뺘xDTtJ�bC �3��:���_)�˧�(}Y��Z=U�7�R��x�G��X���k�
vx�`��#1Wyu�h�����{��mq��d��.�<��*p�zKR�4W�;�v���h��s^��V��vx�'�he���[��r!�w���kbbd�#g��Z���/�fZ�nef~��|��Ft~�շ��0��gV��E乘��8�6k^�
7{VW$�c�kn�m$��X����iB��`` n�5:�e����%%.�c�Λ��]\aU}_}��{�m�)�6~�;=
rgL�̞(l��PjL�(�Dj=a�~�s�j]̊#�1��+;I���`Aε����^f�\��mb\O���Y�x�6�����q��Ӯ8�y�����L�5^��9O�� ʋ�3�D��S��;~��?]�ȭ8ڠ�����溱�!yP)H�xS���L�qeJ7dD�&d�R����~���.�'����-q��f��S�1���`�B�����w�Ĭ��,�Ti% g��|B����E�V��U5�?�j��]qמ��fC���J�f��0��ީ�������܀�`O�*â]��2�ya@�@p1K����	S.;��!�il��E�U㧆�ph�y^R:8�;b�*�A����:LG\s�EAL���.���)�dDV��.F@���Nc��?`�Րn�~�'�����H���Hy��J!��������F'A�� �^��/�Wd�Κ�=�}Z�R����	V��i��ȶ{M'Uz�z��~#NC�U{v.�RR|¦]$r�M�8;R��_�E�^j�����F�Z��ZA�X��ub��� �g9b��9h��(̯�۰�=J3/��l��4f��Y,ݬ�jS���t݌t�s����JnH�|gnޞF�`�_.����9)�m�"��z�#�{�x ��r���\d����F��Rj�/2�;�
�]Wy�-<N0P�3��t{T���uqmFm�au�62V��S�q�mUѼ."Sr�4���o���H��&Տ����v���)��p�r�����j��"�6���7O\�lҝ�}���˥ݙi�Y�� �����s��.�ظ��C}ƥ��Ը�9�)��u�S!��̭�v
#f�<�7oWj2�,�G T,Y#+�t9���u9G�"x�r��J"���̺-դ�r� Ϋ1����lb���6ƪ���[ƻ%���2�����2��������3a^h����;T�w��D���������N��o��t^���,�����������S�B�ގ�	�jgn#1�U�d�b�����8\���]��]����XI��G|s�du�T5�;z��s��0.ϸG"�Į����Ӟ���l�%�q�����A�}55���zA�3�xA�52��λϮG^�/�R�CK�����;[�<pJ*Z���K@�7\>f/�y���Y��m)<�l�A!m-�l+�����y\���|.���aͽ
j��3n�#�x��ż�mgm�����7t|���2���x�����Sh�m3LI�ڍo��s�[��n.g�C���㫏lA�7S�? ���{ӭ��G�d�����P���I@H��h�>��T��M׍ [=��H�����fL:̛�䅮�5.=��A@B�Gh{�P@�a!�;�WZxV������y�6{�����R^q֥F�;��n��Po��ƇZE�K�[��iߓ��^�ץ  �'��S�9+���M5j1ˤHp.;��lC�v+A�ʃ�C�w�,C-��mm�]E���󺲕�.�iڽW��H��	Pr[s�Zf�DtXDdD�T��M��2��Ie]�����lE���,����ȫ���67�q����H�b��&Knb5�uQ�nQ���x��g��E �g�,w[n.T�W�ۋ͐�ꫠ�u\F#�H�I#�	�6��N����5�YE�zqPU�ʳ�҅+�+�+�{X[ο2�����\���fw�{�{*;�sU�gє�⣇^T���s4�0�b�=5�Td��6���X�v�l�����PP೐Z��F�1�^��Pʺ���K'vVp� �h�پ0:���@J���Y���7Jn�7qg%w��T}��ѹX��L��%�5���[��ue��iE����3��+�kw����w����tp��^G�����F��w�͆r�����(L��R���U:r]gwp�x =���j�u\3�&>2�+�q7�Y��t' s�]-��9��*�b4���a��;DS73��]J�0vG1J��rF��,B�Yd�)L��w�e��Յ����VD�0u� ���޹���"��I�Q>�%�ѥ�U6s���}��>Q�8�r�A��
L�"��-b|����c����ϾӢ��x�8�P>��]]6�)�-H�5�ۏF��Z,Tj��}H��[q�z�Z�v�j��S��P�d�@��$�9���xos�BVPW��mk:�d�]r��'�FE��!�6rl<�PN2K4#�zA��H)V�(�rtU-��Vxd�Q�}V��7�Ԕ�l?t��s����1��(�
d�z@k����l��vtG���ݠP~s��n����b�^��#��r�n�#���g&�%��c��;y<홷g	P�T�S`�D&z	+NFdl�o�x��˭ѿ'#�8d�%�.�y>&]>���Q3�m��:h̏zv�^:f�^��+7�x�H��^z�X��u����>�j�A�O��y9�3�����Nc`�VA��Hv��0%2wtHum����U�.��\ݵ�9nnmn7R��'�y��4;M[G��,RN�ME�oeZ&t���7�3L>3����ůn��T@�1&9FrЌ!����x{i�����}|gh��ܤv�����$�OUP��:��]��E��\68d{�4���}��t�eTd���@ll��Xj@�5�L�d�FH����k[�j����؞��� 7��;_�nׄ�7�R��Ǌr���k�����7	�y<;����#:[rtR���F2�'�N�6*dd�Ζ́�j����T�4s��=c��΋w ŅV���_���̆�Ҕn�"�0�_��93�jg�(�ِ/���*�L�f���]n�����u��u��r5>.T5���#f�%�[	}��_1�W�pi���2p���3a{�w51'�^1��cNA�@@p;�Qt Ξ��O����{���'�����ь��CB��i�g��t5�1�E.���@V_���W��>.�r�yuv�A�*�9�3(�b���y�����$(ǲag7~zJ��B�E �U�yPPZ��v��n6��FwJ���K6(�>�R��9�F��0����N���#�ڞd���uk�W��(�U���"o����߁�mK�;.ѷMG{���F�Z���+YZM�����d��.�߹JV���p�3EF����;Iӆr�H&(n-	Huѣ�*��Z�S�M)u�����Q,5ze�B��M�㝊Ys��=��3?�꯾�ｎזq��� 	",�UK�[����6��bne�q�C����06��1���P��{�l�Bb�*x�ɘ0$0cK&!ߡ*�P���=�.5�]]S�Ȉ�=�t���DDӕI�\�vvD����͒x�9#Ǒ"��b!R;�LO�*�e�2�X+��E2�PK6_s���օ�2����VY�1h�a��R�M�2��	V�|٦�"��I-�u���Y|��}���&-l[��(�!�O��L��ˈ�Q��	�8�v����yBv\���5c&k�q�p��3���Y���]5F� hP��0��#�U���L���x�m)�U�K�B���V�lΞ⸠��Crr_�;�85:�roB�����%�)s�B�e��cغ���`�D��q��Bn�e����t�o�����zE���eowijJ5|V�;�y��s��X�C}6��F��J������9G��,�Ε�n5�Ģf!B)@��vcw5�Y�-{�?8��ʹ�N3�en0xU�[T2����p8����J����y���ɷq���BO�9}+��pfzo���r�1������b���%R�e�yS#�K�9���������m��W�q2jqx�B�91�m�f�MW(ﺭ��u�v���Γ�&��4���k�U{sb��t�3��@�9�}@ r��w2h\G���4�рK��`�^�-��w������%+ Ϭ���כ�b�oL��{״>6�\��C�cd�"��B�8`K��yoϢܶN0.o'�_U�O�w��˛<Q�����P�9���m*���]=;p��"�q�+o�f�qm<�v����oF�����'=Ih
�v�v*e"8�w��ҷǙ�^�F�M���vx��Iq<^��2����0Qa��+���k�J}}uI��7^4[=����z2�r�B��⬓�h���W���^�(Q(��b7��C@�a ���\*M���i���|��}x2uEÞj�p�eF�u�M��:o�T���D##�\�,O:�=��^����d����������1��~��}ɫQ��]"E�FB%�9�݊@|+*�	.�g<�)?J��l���+�f���o#��^Qڑ���9-��-3N":,"2"|��:i��`��׽���<��_x�G���)�x�9�i����T&-d��ۨ�{��S];S���c#��y]�L ,�S�g<��]qN������:ʙԁ-C�,���M;70�m�&��8��ڃ{;���,�9��ps�&U����d�EV�}K`�����v,�X3�Jj5b������ӂ7���f�d�f��VT殝ŻS7����/�4R�bR���U	+�i����LxA�v���+[n/6B�CU允'v�ƽ�PV@��������@�ӲU�jx�Tc��Dp�`�
�GR�$o�eC�ňLW*���g�c���_�7�����>�����+qp�����B�y�WQ��2��#F[�n����l�yL!�e�R�1�SC4����EoK'v����Q�м�bW�k���G+<Ĺ�l��I��Q��S��9����{��J�{-@�S�'��^^�q�����5Mك�9�uH�\�ѿl���Y49Je��w�e���Lq��s׋vu�M ��pz�"M���Қ^�Sg0�;������e�ٛ���|��K/CqY�f�������H�żD� |+����#�����+56�z,��[{�;�Ԓ��]��Ȅu�A�ZϮ.�GI=DX��HgʻH�y�~��s�W����'k��r�"��)�0>��a�A��۰�2K4#�zA��nD���̟P�q���b�b	�s,)�&J��^Ƀ�Y<���N��V�H�G��3k�*��gu���u{����
s�t��>�������q�ifι�+�n����,{{�vq��5�W,tљ�7�\��`��q�u|��^��� c���ET]�]<O�'����щ�	�Kv:!Ծ9�n�8��y����#������W��&��1."�u�("�}&�C�{���&�6Ps��m�}3��Ξ9��{��.q�B��D��N��hC�z	+NFdl�o�x���]n���t�^>�"�0�z�=Zr=�w{�xTAӀ̎c���&��3�Ҵ��hy�)C��p#ԮQ��7:�}�z�$?'�̛	��+e�k�'�nz�+Һ�Eʗ��1��b�*�9J�+��Gf.6)��~ض��E�f���MH5�L,��#$wX��>y�y{s6�c�M�����	D1	u��Hz�Mˍ��T�_�'P�ߋ��;6܊�N�֡�%y�����]
��:NV:�
x�}T����iU��*�w�̝<.�	�Ԅ.>�uo��=�J�=�}8��ne����\\b���+�x��|kUV�3̔p�o���ʦ�,�F��L݌̬&�ۧ�ޖ�����V��V.��ٸ�t�I�6,�cڮ�.�UuTϹx��%#"�^ZOR�ۦ��w���p��h5g�d�l�y ���sy���)
�2�ĺ�/���:������%�e��Қ�Y׽ʹR��jZw���o���������Dv�w������b����#Si�6�gV+�V];�Lh�]v�$8�}z�f���q�4W>`]��QwJ^;櫥�qv��w.�I��6��
�v����0�x�ż��؇ZBTsm�R��V6�Ď�·_�|�,�qg�����:�.���Lt�[�'�i�j6e�y�҃*�p;Q�@���}���Qj�.�*2S���+I�ld��&�ZF�	�θ*��:���;1�=��iF�l�^���=�6螕�W;5S�9�+�]�t��v3Q0Ǐٱe�vh�O���SU��̅�wo%�jJ4̤�n�[r��2>��\��Y��t�o��ܻ����� oi�[���}����ȭ� �	zg�m��`q�aǣ{vC
�ˌ�W�8�Y��^˧R�qGre�8�6_=Y+R��:��/&��Jl���b��۰�Øw{f�f�ё���5���9ӼoVYa�C;��S�acG+��&]�޶4�.D� �Y�wU�W˟U���÷퐕���g�ȭ��ApO64��Ι�r��^�{�y+|���.��&]�bUalo)^��$~��^].Ʉ�9Xp�]a��Ѻ�7mc��b�hb�z���鏆�n#/�2��U,S�;@�WF����#�며�=�R�{M�o!w�Ys�fX#�Ȓ�Ms,p�N%���Ѵ�,k�H긳��ۖë�G�u��M�O`�1�d�Aق��W�#y�i;����k�d��] �
w�^�޻tD��X�g�{EIJ��=Nu:wtU�p��Z�[[�D�*E��x�����d�-n^'N�����A�TV�ɜ�3)�y��A˻�D@��_+��Isދ9HA`��W�t�S��Ǒ��d�R�͢Md2�����
�WG��Cٸ����;f�m�{��A`V�%'����7C1�g��e���C��А�`s�>V7Y��3�<��� ��W48�����9Nʾ�js��%������y���n�l_�$-�|�
z�7�[ "e�oa����ù,r�{�o"��b��?D��P�J��Y0�X�n�5�@u'fg;�%L�®���h�Lv��؜�
��U֎8#\�W鶺'����Y�$��U~�j���QY ��c�]LY��Jn�1��k�lʘ/qO�:ё��S�k{�롽�Ȭ����n�1H�99r�a�P����W@�Zf�%)�sh*����nlf�Y�pRg7+;RyH��ķ|�s��r��r�۸p�l1�ҹ�.�S�]\��w+�v�q.tb��ۢK���T̺	�`��79+��[��ǃ��F�w�VG.�)U��9ΐ���
�sZYCU��!��hUP�*��P� P�
��#��I"q�KA��1H ī��(*J�	H�2�D(�L��ADm�4���L���H4��$�;��i ���wq�nɄ�b#BL�3n����S�sF3iLI��h�P=�)*�L�a�ssb�X(�BRhđ�Zi(�1L��.[�7)65"$�4b�F����!� i	�k��
H�$ƈ��334���lS �`Б%œD���	+��!��1	�1ll����E,&��I�BEN�^;�9�p�ق��N��asL�65�^�qZ}���V����굵j�h�e���R�>5�n#��c���꯾ b��Iv\������N��S�3Swƶ��8X�
�ep��XxJixS�gP��	�3c&V����X{b�U�"��J���N�&/�[s(�" l���,L맲�ɹ���ռ�H�ĺƣ�Y��D��	�wpin�3X��,=�[�<<�����QQĔz(T���'��'��*���#(Q��ݗbQ�Z}	K��9�F�h��oz�6�'�t�J��W�S>[LA��X ��]���P�T��q�\��}%��l�;Ny�07�bD�G+f�>�=J�������5 Em�m <�w?�3�/�B�CWGd�m�_t��f�maMp���;8t�T��^MМ�wl�ZH�u�Z�b!#�����*�ZW�m7-�Kٴ��=�{�'���}!�E�|�OJ�R�Γ�+�������4v���9�p���U�O�"�H�V�֪a����ҦK�e�s�FDHN���� �,4�.w�Y&��۩����o$���!�M�a��7�یmUѼ."Pn\F����lg�� eE/����4��;5����.1�Mo���C_oy�7��ԥ�J#�ݑ��)\{.�z%���Ժ���q��99c��T��[��ȓ���7b��w]��xCх^5�ά*F�U�JÓq&�K����]��̙�����Y��~�x[ŝ��&�̢g�A�F0�t��:+eqh�	Hح��c���S��&��(r���W���>xWXd�i�J��k´*1p�-}�/�f�&w����k�+�V
)Rrֻ��u1�U��W�w`����"�١�2�B�>���u9Dœx3�DZ�����qI�2�s��v�$�c�oҪ+ӝɋ��k�%���%�U�|+�x:���h��M�s|��no$��!�D�w�b��y��t���:�i���&n5�}��} P6n�������x�"�r�[*'�Qg�p/�[&(b���9p5K��VW�vTƽ�0�2ڪĥ��f�,$�~mz�BH|vQ�1+��qt��8Y~{a�.Z�,�gv�J��/{���'*0E�g'Z�]\~,T4��XO���ps�e�U3�F�ݥV�|�3���iu���2�A�(�J�z�iO�u�&e��r`�p��ٙ{i$cl�t>z�#�Iү�.=�ꂀ��{h���@�a ��n���L����zC(��}z��������N�n_� �V�Ln�<5[��@d�(����f�nKݫ��Ds�+WD�K��2kw��N����*�u�o$�S���!�k��!0��֠7��q�WG�P��p4�o.{y�m<�s�.F������䳖�F������l`�����Tn �w~z�N�2��\hq�(v���ք,�/�x7���Ĭ����o��KUɫQ�]"C�p�m�D0�
�Ad_*��ǔf�Z]�o�R����",��c>ӎf�8�jF�_�T�m�An%�F�"2"��fvCm���9�z�f}�/�tu|����ff��7�����ΐqO2d�i�N��-���.��Q��c'ܪUj�N���y�[g毙��+���5�.�o�ǲ�c�{��:�h��d0��V�;a��7�/L�5w2�WCyJ�hW�W���Fo���Tg�c\Qشf.:���0ju��>��<U�0��1 l�ϻ*�$+��*�̵�V��..�
�%�%�\(9x��E�A��g`�T����j7���rӹd�� �Wo��� &3��B<�ޱ�m;#1}�Xi,�;t����ЋN�d�j�ڮ��'�L�ts��I�������k�3	�r���qV��|o�@h�̱
�K,��)L��^q� ���i� r�#}�Xݽ{}'���96�۱���m�*�S��im{çA�mdKP}�O:p��j���*:�o�gyN*�^�kE֥rp��t�kT4 <�O��Lӎ�h�FY�}{��|�'r�..�lH�Z�k O��Z��������ϝ􁠍G�?J��U��LD�TN�?�X9�GR��/��*��;�$���w:{����]��8$�����	t8:x�8���\�k�+$~|�=��]����f�T�X�k�1T6
�J<��:Q��B;A�a�)�@�
:I�2�v�Us�kDn]S��pc����#���^�%#Ls�}��I�λE���3�^@�"�O�F�a]C��"��[�U���Ė�tqwO��;J�Dm5
&qE;��G�7y��4�p�`#D�������&�AwW����9����;Y"ͩ�OPk���V�հg0?}�ؤ�"xj'���� �L�M��l�oO2�.�E� 縗t�!We�+U>�����oIx����8��*8YJ�ժ�r�+�a���V�gu޴i��]5�Ӆq�sܨ�!4���' kQ"�l�1�(��>���
.�xl�S�N=��^���V��y���X�s<-0� ��<���F'<�1�s�b|۬�)]剱�G]�������Ѱ7T���P���,F�n��d�J�A;�Yh����{���W�@�l�{C�������]�N��I;�U��y�L�c���؅�L(vܫ�Y�kX�f��m�eZ�d�]��GL�4����ﾯ���!&zc)}+��v��y�6�9}x�f�pO�y���4�Τz��W��Ta=��7�����ꕑ���nW4K�i��'��B�9����yA����S`;U��
��*��1�Go��7�;
e7���[��w��P�Q��=�>�T�g9���D�9B%�;[���j����y��1h5�����]�~Oz�^�z/��h�o�����`�Ϙ�����~FZ�0��a����\�?v)�Gb�Lw��oR}���m�+��'_��tʗ��+[��ǰ�����ނ\,�_����w�:�� ����a>��Eԥ��I����[a�-�<�^�v �ށwWR�����~�$'�ݴ��X���-�O�� ��u���*awt��c����Ni]����w�ބ�H��{t��R�s]�du��g�|^���n �u�#�c#͆]����ak�Y��efp�{Z��j"�ڑs.Z�fQ�P�΢���e�)WWI��.Fx��%d�+�#.C6�J��8 �@��!����,�|(c�ue��橼�(�}_U}Y/'_[lW(�K�GZL;�m�n�� �)�L.��'�MzV�k1;�%�ŧ�]OWK����-��� �5p�C�ͨV�!R=�A�Q��]F]��!��N�Q������ğH��}SM'�cZ����(ոj��Ӕ�lnsHE���
�/�ɬŻ�6�k֘F���7ٔUr���s���/�_���<�����}RskuS����xG=�]�b��s��ӷ�/
��v�����V}4Fb�6������ܤ�Dp�e��:���!Ύ�})��~ۛK��i_ZZS����y��l��ӑ�n�ƶ-� ��9�N���}]ڙ��m-!mN��U�|���L�bmV0���]���q<�abo�E�����%�ky�3��S���u��t%���Tޱz����a��-d7��b�}`K�Я�j�%G2�����WZs*�g)=Q��"��_n��{�A[j�,��Y�jܜ�7V�5s����/����-�M�jG��[�^y��o�%��WQt�z���݉���HH>�Wd�]I·z��E#_],��M�������2�TwOd���{޷Թs��WRL�lGI|#��/�m UbT��Ky~�ǭ��a��M�keb�{�y���'�.����(|�IJ���W���y��ƥ'k�Ssi�E�Z���a8�����E/oB�>��OJ|#|���<ј�m�(�k��>���eT������%�mnD���QƧ[Fӣ��Fj����-�~�V�{�^x�PuNh#
{ˉ���M ���y�Sȍ��Mzu,�-P��k�I��h3�+ͽ����3�Қ�S�P����:�D-s�V�׳y׵#��9M�4���d^6�}���Hu�k�yP��nM	O&���<|U33�병u7��J���[�Z5؅9Z�Ď�Vy���k"As��o���^z��uV5=�8�9��Wu[��*~@��̪��~��y�^P��S/��ϗ�
���S
9erU�[�o(�~���<1��?]�7YM�C2�*W���O�N��4��P��U�4�־\���,��\���P+x��2e]9N�ިF�jw.�uE�]G-�n�1%�je��ǒ��N5�\	�u}��:"��{���e�{Z�{��3���M�e��&9��1��YT:��gFeʃʞ\��cy�-�1��o0"^F_���2�;S/b�O��s�����Vo7�wa'fjUo��z60U�rf�`��u�B�(ޖ���u���T��\S��Mqxb{%��h��M޸����W�{K
��9&��˱�QO5��s�p�0^���NytQ����P��������&�=K�Ls_\`={ڹ�p�6лoT����ª�#d�>W�=ޝ�k�v]ِ�np�������^�5����w���E�#�ij�c�ł����2�mC��V���)i�Ry|��Fm�r���C�]����1��j,�Ǥ�/W�>�˻�@��aZ���f
��^z���wX��{��.`��f2C�t�[]�.��&��z�[��٪��/#
�D��!��HN�ώ���~s�S��]p��H�7Wt}2v��ZrЗ����v�guc���]֥���|1���<[��us�0�Vb��i�w6w%ئE8�����#6�r�} �:�����9r�>OM��"Tn��h짏�� N�6���'��OEtۚF�t�M�w}醳�G�}�]vS���qb�{u����KK�;f�50*Q=H�w��vyZ����8%##�����kQ��gZNx&ƻ��vc�n���G���
'�F+ޗ���.b[ɬ��ެv���L"��S#]��4�rr�@�e�8�\Ќ�ru+0�׽����X�L3V�o&��q������$�s��О�T.��Ok]b���ە�{=}u�rj�F���1f�Vm�Е�y)F�ǽPU��7��c
/�;�&V[YC3�n�[�;���[W��};ܜ��s~ZB��KG�5�n�.�nz�(]m��D�^�����DՊ`"���E�)-�]��VQ��whC�a��|��ע]u�|���<>��^�j��6��o�����Π����=ϙ��=I���j�/*r{�����#���f��F1yBs��!Q�^�xse+�ٰ�I��d��\Ze���=|������;2��'T�,�ȥڂ�t��kU��4�Ǖ��R���]��=#nZ��n%V�ʜ]�ڗ.T�q�K�&������vS�͞(�| �P�Ά�*�ĩX��X�Ya���i�����u_t!bo�x�J����ȇ�F�k1ܸu�u�)D�O9��x=��1V9� ��+{8��t��{{@�{w�5�O��*�Db�$�,�x�N⣇i4�6Ӌs)p���C"ءj��Ҟ�b�.s����oi��T�>a֤����2�D-�}���P�y�kGpSN��Ȭ���6���Ր���o&��v��*��8���<��lnߞ�zn(�㊵���"؅�4'VM{5-H�Z�Iðc]��|�+yP��f��/w:UʛW�D$�.A[�J��f�=m���Ѡ��+���9ٷ������rXγ�襁��y���{�1M��N�pz�
?	��)?=���q��-�O���e�Y3s�[����ξ"��[f�\[�3g��-�u��97z�۶�R���ҩ:�c{J
�Z�&�[�N%*؎[��5�Xi۹��&��8ڊ1�S��U*`|V�.�EƎ��������R�mS-�����Η%�4�wQR�3��c��䃛G9hS��Ղ��&�H�*��97���!����Wh��rdf�Ѹ��e��KW��S��SEj�R�e� ZE�V;=P�n@W06�-M��k�2�qʌ�Mǣ:��T�b߰M
����kq���7V�-�*d�y`�Ӗ�\�W/�0�Ss��p��޾p�wY4P�Q[���A*hB�|�wW
��t7'R3�ML�S⺂��l��&�3��郩h`�5
��>����^#��ŗ����*
Γ;�ym&p���S#�aj,�gv�T����*���,�o>�#�1g�֮�T���56�t���)��뿮�\G/3V���Z�<��yZ���5��B�<ȹὓ.�n)���&�Yu9s0��Vb���u��A7BP'7�W̍������8��+�95j>=N������!`�O����98ɒ�-�ܻ ���<(
�ǐ�8g%X��,U��t�o{읯�'^c�������Ȭv����8M˃\,k���T_,���C뚨-A�y�z�kږ��L���#������Jrg2y
�MT��ಫP��e_��f�DL�Vk��y.�H,��x�7��Z*DҹQJmN�t�� ���v�b�����cY׃ ���}+���+�u�{�L�Ώ+���KX36v����*�"�nU��}���t1�pڏ��`�9�m�š�k�_㹕מ���1-��ފ�x��;�Y�@q��u=��Y�Ƨkt���V8N%���0������ju���uR�4kv���Wk�.T:�1#ϖ��������9�`STw�-���4����zo]��Q��%�(��E����>�x2T�3,<X�`R�o�c �t��k1o쾺=�7��fEYbz��e��Z�'F��2^����m̚�ɑ7�-�U���4vk����j=�m^��Ƙ�$��x��e(��Ysq��-nU����^}����u!��a�n,�/I�vd�ޣo��&�:��;��w]Y�a�c����q��Y*ak��0q��k;��}uq0\3�ܻYzљ����<�جrv]s}�:vs���0�S+���৑E{w[�I"����ӥ����y����b����e=�;er*ۢb���ccط$�wZt�ܮ�|k+�4�%VQ�J ��ڎmoP}v[�NYՙЎO3�K۬��ǘ,`A�fa`�/�u��d̦�5�V0�J ҩɆ�Y�hh5xӠo09�bz����f�kJSʾh��ړOmn�07�W����&����f
*��x/FV��P�G]�0��^8�p�8�n5M�bwh^w�����oM&���Q�fd����g��s`������Ke.WM�v�B���h5WwRRT\���cn\6�F,�&(�\�&�1c@wd,dۗ4E����H�$�bB@��4TlwtT͌c#lQ��\�X��L1��4�Ef�s�0(�*�R2�JG9F˅wU�I1�w4`Ѡ��ɱn��(������Y1d6 �"59cr�F4�뤗;�F��1�cs�+���u�Ld�hP�0�S�I`эw[�F�B	���⋮�e�3r��FJ,r��.�����G�d�{�UgY���ХsEl{�l�?cS�j`�6�L��ۘfqiKu���_V;�tw�E܍�n�� =yk'v]���s�N��m�k5�v;���w���v��](�Y�+5�/��u�Z������H�|�L�Mgm�*ͽNj�2�u��(q)78�͛��_���r�O�/�Et��`��ٚۚ�G�,�-��w_=S�����];�S�z\��	^����{����X����W����2o�����d�"
�K�\W��-���j�d��3Τ4=��G��V���ﳤ��S~�>[�
��T���ڝ�0q�D��kf����oo?><�z�^7~��>Cz@(� CK�B���7��V֍����6h�5mj�:����+��=���y�v��z1aP9ֶ�T](��q������7�b��݊x�W�*���x'	�(*�sI��w�R�1��QZ��wb㼚HC��R�m��qF-����1��I�f�D�S��l��A��^���΍#E�u��T�f7�����͜��*ֈL�O	"X�KA�NݔF^aW%5a����dxmv���8_XK��
V>��s/�$6����F�#����s���%>�N�=�E��F�c��x7N�ync����Թ�S��9?Y����75+r�o<\o��~M�=�� �3Z��В�>���V̞�d�Sx=��췷�gyfҜ��x��B���H���t����z��lk�$tbyFȋ[B�| �{r����s-ken��<:b��Ͷ�W�0�hFo�ʡ����V����$Q���'�z�[�(V����ܬw�__�0���SYU�7C:2��M%�C��)-�����F��쌱���>S/b�|�xs���7	q�Gp14��^�6��"�~��-�5�#p�q����5��p��]RoVX�k���˶j
߾��w��������_RίCHuMC�kz��/R�1�����g<�?w�(Cu��	���>趐T"�0����k���v����n+ւ����i�����[�X|����r]���#/�wE�0ݺ��(�Yx��/a�N�.1tOBn�vW�
�r��w�^1N��w���b�d�5*�
X<!���w�S;�t����*��en��δ�u!zI��q�ˎ����+�蕓r��i����W[��/�x �o5��uK=������'T17��V�����+=�nU����ج�7���c�=�o.�(�� Ry|��{h�q9oe�G�%]����n��)��0�yd��1��G>�]؟-�5~>�W��ג�� ��
e:2�ɮ1�� }����.��ұ���6�h�&B��R�}8�$�sw"�oh9�4�.0�#`����y����íy�Eo%�e�2�jKa0�:W���ʵ����Ȩ�y)�e��Nue1��)ndf�{S.�}S^i8��O�f�w���o>�w�TZg��8o|�+ѩt���K,N�������M�m\^�02-A�ǁ�S�ês�Oe�f�-��;mL�'q��Rsߚկ��F&�t��we��{�$o)N�צVElm�'�|�ј�M��FX�N��I�^R� �!TgG	�/r#Gd�iL��>�o:9�~�lN�oP,�fQ%��i[:Y��R�j�s	�1��M�*i��@�I�Ɣ�u�S�V+���(k�$5���]f;PG�[@�kTǖ�����,<x�G�{L]��n�O�Žןb��xZ�g���>{��:��r��dc������U\s��En����ꆼ��z�ݖv+����S�iAx���5������h=��ۼ.o�����:�%�q�fD��{�ާ'u���g���<�,�������O\|r�`�'���#����u{�1�d71���}b_>�9Ժ��·&�S��֪k�K�}]I}Ci�J�4���5��m=��SZ'�aBf�\%���&m���{Dp>��^����t]JQ>ԞX��^F^V:rKY�ː��-%���
W���c���{<�J|w���ȹv��=�<��H��7ֻs��m���PW
G{zA%�p��oVRĻ��*%:�wt������ܻ���Y��<Ƞ�9N��yS��t�����CLZs���ȷ��T�`����2�g7�A���6���*�����G9Y�ڑt���v>5j��RȦS�X�Y��KC�3u�+��/�y�5���j������u;�p����m	]��ta[�U��pe�(���N#�ds%�z�n�z������"����R��v�ga} �k�˵C���/�/�N��O�������f�sթ-s^i8v������Qpo��r�7:#�ן w+��L;�M��x�6�m4z*n��]����Ce�	�!NP�������P��^�Z�ueU�R��h��f]=�V�����i�H#Bڍ��V�5��/f.��-�O-������gFW��/��l�t�}�U���2t�R�0o��&Z�ǯ��[��H+��&$��b�k;Ov�_8�A��H�N�^�\���?{�t����79^�}ׅ	��讖��+9�7�))�H{S����x��3m���:�������KU���rM��*y�Y�}�;t��9'��Kyy�~OdA���܀yȂ�Ľ����s�XZcq�}��iu�w��.�����g*��"�Q�uH�1=�]]�#�hڇ���0�8�+��$TZr�FU��Zq��t�hVojc�g����y��s�r,����c7�gR]L�*�7|��(�1�L���IO��z�N]�)�pwt������vl��5sܡ��;8�KG /���;���9j8!�S�C�f�wB��j�1U��oo��T�W���p��B�wDl�<(GR̎���U$�!nzw]e:)颓��k��{޶.Bt���R;����ɑ�3��M7s����[�&�zo�>�o��;kp'��TT���W����RFo9ձt��>�)�|y����]��o�4�����FIȫ�](D�٭/j�,za�M��A��;�Oe�N{~]ߧOe�����Y�3&�,G���s��u˄�|q�>_co��zҜ���WO@r�? ��e������Xz�h'�lc�s]�Q�ևQ�W}��䊳15�1�V�N����5�+Iզo�c��vs\t���<vz3Aۓ���drELe&%�P��w[[���9}������5��F�4wU�a�f��Nwta=�Ǯu�V:Y_)؏��do�|�u֐A�*�rGl�ˌ��q*��^uj�2q�Y�8��=���42����v�5�"��Kpv�^���.�ű�CD\V�盃Q.4f�� ւ���i:��6���S4]_�yHNs�ol��1�uC����{�
�#��+�:�mj�l\Q� ��ƑFu�X��V8c�l�T=ʋQ��*��!|�CMǎ�ga�����b��gi�I�<�jz�C�}aͬ�g�:�
S��q�Dܞ�����Z�q9=Y�y��i��>ߔA��M���pzQ���榪�ȍ�[2tk[*����|e����h��ThM�v���t����,��4���S��.�U9w�J�7}�5�agי�˶�n2����\ˮv��	���F#vAi������KM�_���ac�7��)���oF�p�T�\����*9��Չ���އo�0r����a0��OK��ze�aO{L}���⺱v��=g;XQ��<�m��)4m'��E ��i�#�.�؇����9���4��m�^F�1@{�N�	�j��	T�Q��ѷ�{	G�`���)Q���OMר:!V���n�Cq"b��|�n��/�,���}%�x{�J����V��6&J�79`�����z�wg	Y�Rp��e�]�Q][`S��PG^�,��J��e����t����W@X�r܃p;Ǳ����a-�IЬ4�t������De�Cy^o�i��c]��S�9F�甅x�ٗ��uYu��sr�i~Y���Պ�u5i�kͱ��Ŵ����o{����}}�Yom<����I�Z����0�잹���!���׍�]يY~�{�Y���W�{X��Jz�-�7Sܔ��j��0!�u�r:���)���uC�hH�s���1������r`|0��'�։�}���ng�O{
^N-!N�P�W�ńe�����msk�6\O�|�+�<��w�vm���ga��8��k�0@�Ƞ�m�����z�=.�Xj��V0�1�� ��\�}js��5'��f��x�u�:��e�؎�� �%��n%J���X��[葊�<rsj}ݻ(eF�2�U��r�#d>F{�EPݣ~}�c�S��#Шb׷��{��`M�"L�rS�b��nNs;�*cq1.�sk��q�S�!�6z����u��%r��^�#C����J?����1�W�=״'Vl�	���3�Ƀt��8=�q{��B���1՝E��3��y& 5�0$�밻��K.����{ӭ�W)��/xم+��P1�����<��նbn�Vx7�0*Y�ԇ��|�z��w�ٵ#��>2!-������/�2�j	�ڣ��9�}�m+�V�Ov(<g)�4��[�h�k��u�`t6�vi^�`fv��W��T1q��W�;چ�v��Mŉ�詹��]��^q�P貵�zV�׳y�Ԏ%�x�C�����O@�u=��h���^���enM<�k9m{y�U0����곯�<\<|♮ǧ:~5}�i����3�<��}�VD��\���ao���OB��ʟ	��닞�:���6Ќ�7�C^�)o�U�y��^݇8����ʉ��o���X�����k5�ucʥVn�ZW==C��g1,Y,��'��d�{�Iyy�H�i�S/b��ڦ�F��D����Y��E\F�K��+5�n<�&<h6�w�v�K44�Eke�J�l[wM�6=k�k���޾3�e����W�c�l�VS&j*�
�Ҡ�Xu���Vr�Qᭀ�\xSu��:��0p�aòup�X��w�Wk�9֞�ss�V�����7q-�_��"�tqi�^u���ܥoe¥��ؽ��9��&z���|6ǜ5���i�,,��5�z����t�RJ�lk�grg�}�(��wo�X}�=7�HC���؍Sܐ�N�Ӭz�1}��л,�����YԻ
�[�P0�P�ݒw2a��bhͺ�F��A������,���+�	lGB�:\���s�tu�Z��q۪�J�ץ-4Rya�k��gU��N[wY7d`��$�+ ���"�>��r����-�X�o�<��񜁙����_.�x��\&�0T�f6C�pQ@��P�������{�J�7��L�U����[��y�iñ��9W�a���}En��L��i_�y�.9"��6�OyF�.T��C�môpHT�GR;^�΄u�+\Ծ�b���w{��[��:z����Iլ���V[��+)H�萬�W���8W�,-��*WI�yS7Z��vOs{��V�%�7%��0��0򶋫�/v��0�Ŧ'�qݨ�;�	N��]w�d�J��t/��@�z�V̌�Ԡ�|8Z�C2�m�C(m�r7����ˇ`Kj�"��]�w���#�h��$+f�*�!f���g��	Y�0�ѩJ>H�c����W.���MӇ��ʍ��JXQt�E��b��՚' �,[W�:�䏈
� �b������Xz�c�	��-̑����C�J�%gu�h�ϕ�0eJBɲE&�(��ô�P�fj��FstP��V��Dm`߷SJ���n����k�,�ݽ�jܩS9�[j2�X�5v���]K���q�DF������N�7����C��JU�
�u�*�ӛ7��1�=�r��L��u�c}��F�k�@��h�LKU�m��0v�읬�Β�mm>��ȫ�ΝyS��ʍ>iv֎��.w@��;C��@T�F����gq��Ǣ��Nr��g��9V���X�.Gf���;�i�3�K��㻐�ۓk'4td��+wV�}Qh�4�p���,�����͵Υ�
ƻ��M���VV�y��Q F���w�uY�H���|ru��"a�RB���o����v�P����,�6�V\���-ggvv"S��%������eվ7��帒�3�2�>&�4	��M|�;�f[�S��� Vt������/���jN��b#0����M��gkM#�ZgY��5�L�5�Stk2���[UԮ�� v2��YzWV�����.t��q��,w���tL����-U�{�����\	_i:�do�e���l#*�ӏ����wX��2�떷r����7�tҚu�k0dk���t�Zb�"�������hBU����e�8Y5�٬�:�0�H��yOy�xj���;�f�.��p��9V�58��dD1ɋc���T�Z;#�f��.��v�|�p�i�W����5%Nv��gv��a��u*��W
6�m�t���`�L�VjÁ��*�	��/�������`uqށ�!g.>}��J�,��(��o y��S{�EwĲ�3[�5���]Js-�jV�x�XJέǽj�%[��R���Y���8����] �����BD�J�Vh�Y-Q�����f�Y/7� +��̇����qk	P5IK�N�X=�B-������׷��@��ɹ�L�9��CR�P�׷w�[��s:i�UG�E�RAo����Mcm^�5i�͘�*Ĕ��ݭ��(�W#�qL�vʘ����z>��ɭv5�[��+]R�/�;�B�6���Lb�v.?�Wc�^�\h������t	��3��vJ����(]���F̀�j�-�t��0q���j�n��-a�cE��?q$W�@�*��)��Kwj�ɓF,H]�2k��1�v�$�v$e�;����,Hh��t�����w]ݮ�6�D�Rd�(�k�l�(��.�Ѻ\�"�����)#Q]ۡ'qr��	��s�1����BI	QDj9�qi(��nh��*$�"��tX�7��'69��k�[��b*�r�����κ��'+�4H�]܅�K�Q\�7`.�\��b�#m��]�.!��9I�r�GN��q\�r�s���\�>��ٵ�-!�����$
Ū�:�$c���]�n��=i�qXoOfL�����s"�1�5���`�vL!Yuݢ��Iɯyl�o,����?W��ci65߂8']���6b�ס��m9�}&a.ki�Ej�����٫uM$�����؍�yT5����F溁��7V;�<��?G'^�̡<��絹X���10�uMe+4iwZ�M���Q�c/Iת0[��Bm�D�����r��S/a����1]]U+���rN�v�����.߻H���히z�Ҋ�;��R���RHx\���ͳ���kYܨ�Ո����p�9����֖�9Ua���^uz<��DG��\t�,��Ob*�6R��pZXĮ�{ϵDz���X}6q��:_�����;��5zg���QB�.�	����G)��wn�;���F�����6U�ry׶�ʔ�w����V���������qRm�Ե�F�L��2�)�Dd��>��^��_]^���)<�����CHϪ����*B�3Հ��]���[���������5��#���/�1mפvM�t�S֨mo8]ՙ��v⾧r�}�5�r≇�8ӈ�K�b]pU���뉮n�d���0�}\��e^��î�㗂��p2�D]A�5��Κ�#�u5pg���m�}�9T$�!.�/�u�S�@��f]�����V������/�N�MyR;��-��'�c��r�V������uv�T��Z�7�c;�@6��uNh/�e��v��N���>�h��{���M��u���+�5p�CqJpJ�z�y󫻭� ���Vu��1|�jh	�C9���]7�5擇a�5�8&��C9��Y2������輧M��^��+s,JY9�3�6U6�E�1[�e�9t��A��c����[ڌ��K̡8��w-ܛ��']�D��1%ލ��]���Ê��N���<���"�P��Bm�	屶7S���mӫlJ�j�\]^�3�`6�5�����}�k�k;֖�~��}��u��d���{N{͈���dc�����Sp^v��f޽��Qju�}��=�<����o�,EI蚮�9���c	�m�.�{ݎL��̚��36)qA�֦����iV
4��G�+��:R��L�{sM�S�q�ڃy�.�c\�Mb��L��	��S)7�,��f�*V�z7ze���F��!u�5P�}2�w�FV���[��`K�����&�tP��s���S��9� �d�BVE�S���_���n�A�R�u�L�~��V4��oT�|ܺ�ڽ��7�k�o�LD�~�eUlF�n`�I}^�@�ĩl7|1����n!7}wY۲���7�Į�󕈸R�l���)>�+e*'EJ�Vjh:�Y��ֶ�7��|���[A�-�񻋅+��
;�Dwnf�K��)f�����ۜL׊}�9�\�/:یs)h���ހ�2FTet>Eg@��y��J7����������ýZ�ds�r��sC����.R�MS�u]��`,q�A�SR�e�J���y4����~f�6�n�N9��c�gs�*�N�(F��e뚕�5��R7�s����"
ܾ.��>I�Ow��{KtJ���-ኁ�m��9����rS��{E�Q�۵�6���Wc ��e-��el9�J%�C����w�rưFL}0��'�|:#��Z���]ɫ5X	�тwzF��������,��<!�3+(Jr�>����_3u�������3��i�W!v]������:97���RK��N�j�{��q��9����lk�B��5ى�1kk����[���ùG=3���y�0��~�<��u�L3^��m�^��-p��_X}���"wtV��Q��>��wy��c�^���5�c{R�5cf%e�S�H_Gj�-�d�b7�	���Z4�VR>���r�)��i����M��$Ϯv��|��s�b���C���`�N:�"�tqi�N�v��=�D5��ս=�����X�=�9,m���9�.z���W����d��p�V"#z%�M���?:Mk��ӡ�D�˥(���v�ǜ��a�m Q��O��L��M��彸�I��P�;a���떟X+9u���b��~�SW/۞��l�od��=���ByѦ����amy����E-����S����6�Tc�<�����~���|
O-�k�>��}���<oFD������lh�h���w"�u�jܚ􉞇�f�����Gj�%,X���Y�kw{<*>ܶ�+�öD�ok��էV]Ҳ�z9��X�jv�u��ϓ���_ʺӳ���̜�T�ϳ3-cJo+�"
��*YR@�p1;Rv@�_/��B{#�]���1>4[�v�p�b��Ha7'&;z��3�uf�'��K v:|Wb�94�q�#N�Vإ�����ˆz)͹��=+�6	O��ne��h���C9v��=�Uhd�a����v���>T�z�ڃνp��+8�S�w�����qk3#we������T���lk��	��1#�h��4�s11�ՍsE9�歎la��������5n���:���m���<�׆�o�&�&����Syp\jt#3�^eO-}�����~�/�ؘf����qym���O8ų�����3����{ְE��U6��y����D��\���BuYכ\��&*�ڻc�GPǛ^Uf�g����D=|�V���Vz��Ǟ)�ߜg��ݗ�W$�Vy�5�s�yͫp��|.��5�+5F�8�:�.Y	*��{41��NRP�h."��Y�lk�έ�r��{^����V�2�f��AA%�b�+�E�͉"���:���Y��,𣏕���Z#��8�4�4%s�{��b���՛�]�Xhӧ�2��$��ҥ�l��:����KD��l" 0��7-�9�3U�|����6���Q�M�-xέ�{r��[�A���겔U�]�����Vu�VáTo`j�������NX5� �/�j��JWxio/k-�-���8{b�Ѱ{-l<]"��b.6C؅%!�)u��.�-4Ryc�kdtfMW&�]GV�>J'����I�t݁
@^ސP"q^������%>&�����z��/<��,�WF��O�[��:j���hWn���`�Jd��[�z����w��w���}ʙ܊�l�s�F���S8���Ԇ�c}�k.3�\�<�*��+ܹ��C��
�8%R28��
ۇy����9I&�V\�+��侹���jEכ��Iÿ2ƻG΋�F��{y��7R�.�������+�^�_��Mf-�x�Խ;��ng�{�e%�١y��{��$R�l�Y��%y�y�s4~{�[~��uu=/\JW�ːT���M��ܽq�f���:c�X"��dJ������-V��!I4Vw_K��P�ܝ;�r�7�{����1�[���_sc�z�ݩ���.�&(��Ja�I��%��T���[�k�ǿU�6����T����+�YCF�S&�-����!΍ej�Ɣ�Ĳ_<7Z��o�b�	��'���"�/n��%ֺt��km�er��^�i�k5�u}�mH�8��_��7���\�5Dʼ�Z�ΖKQ�11>�\�)�R�u�Y�5�Pʳ���M��6�j+���
���Bnr�X]��r�a�}���B�y̧/�x�I�wtG���e��ޢ�F��u�W��{��6���1�2�\\�I�v���Ü�[�y�T$����U�R�-��]���Mm�\��o�ڥ��N��i�����X�l���ʽ%'}tS�wGX��w����u��V��c�[a�,~����A.�5Q�#tKm6x�Iב�ɌƲ�ؔ�׋}���}�m�:�}҄�~�c8���V�Z��7�[�ו�2h�dceer��p��S&�.����Z�փݸ�36��(3}A1�� t`�(��fS샖Z�qJ�a\�O�
K�}*»�T�d[����g�i���{*���U�n1��9��QR�D֘�|��ב���v}�-�1�rV���D�w`bU�q}X�u�Ҹw�p�b�3���]�����*��ۼ��{���+]���M+����Q�b�I�%7ۍ�1�#)�x�-P����	[�Y��ڑ��\�����+�)�.�3�������g[�]���=#��<qR��=��]�2�:"r���4����[�/����6ƻ�(k��Q�赡��OfLF�4�J�ռ��>���������^���V��#ֺ��{�v��;T�s>��4Y��J�/Dg��^��"�2�[l	Ocou�r���/���uCU*�f�MFW#ǐ�o==�I��cw�.���t�X�{Խ�ӵ2�-�]cUf��Y�7=�ӷ]\٥���M\�����p���g�޸:�:�ٱ���ެ�Lz�z�=��;�㲊�w�\�{i�K|G?%���-���%513}cjE2$��+]3*>�fܾ"�FPǼ97���[۶�k�s>�8B���,6L��<��4�F�u�
��)�C2��R���4m?����-6��y�Ӻ*���>���e�p;+�2�|��=�]�]�n�9�.s�Z�~���=M��/�l5��3���F��0uT��\wDq�t� ��G,y2tk];[��Ym��->��AvU�Mm��k�n�E�|��9:��WUB{��i���5�簶�Ol���f�tE%�v_H�{��ՓY�|#vO����-0��k��{Ob�]F(�j�ؾa15�����xX0���վ�]^���}��k�y8Psx���=$��U9�aO�˧��������u\\[@Q���0�/N�}k:K�;�����ۚ��#`��MJ��	�������rf���*//s����o�����T�z�ڃ΄u����>'^�A��v�ֳw��{�C��_7�4�pSc�k��7IΩ��Q��jB/E�`G\�����=��[CUZ����i�}�P��[��%�N�}%��(HI���P��9��*Y����x�9p9(�Cyo�r�n�k;�؊9C��n�3�P���0��V���7��W9�H�
�)���EP�&vKwW���s��L�W������M)�](�F�Y����)v$�h��7�Ζ�~��쪲��Ss�o�9�*�ͬ>s��Wz�!ͺ�V�x���%���"y����v��w�-e��K��w��)�G�hH<�� �k�dw:%m�nG�l�^�����r���	�N�][�g!��}z�m�&�0�r��Sq�^�5^�8g��ZB��P�V��_�\l;+X��cF����XS��p[yޕٷ����;�����I�s)��떷�Tֈ�1�%��g��Q@_�+��l�{}����8������M�s~�6L�<W�ܨ�w^7�ҟs���/W����Ҩ�SY�u��~���v��V\9[�
C�RR���Zt��#"�$&�^4��j�mF���v��i�LE��(I�K�����˳�|��V���(�i؇o��ڶ�)�)��)�o@��� E�����Z�\���GBU�.0ͭG�O��E�U�R�kU��^�@���4����3�)F�7؏J��}LNd:��#SQ���</2<�1؅+��J��uf���;)�1�i���f6�<맵�+<�V̬��ms��7P
�4y1��'��U��)5P�YX�p�H�,	�h;}��sn����>��iq̰��m;�Z+>�_9P�g�t�惮w^���!�3Feqok=��AE��c9Ũ1^���H�%�[�&Y��1�-
?h��{�`5r�'����uY�Hv\3s�|6�P����e��ה���ND�wy\c�dO�.!""
֥[��u��R��j�����}j83^4�`��hG��䮦���T�����*�;kpR��5)�Xbm�w��\e�uǁc��§-����g@��-�X�tF�]=Ē��񅁵/���ץ�a��M&�Q�C��:{B�����kz�Q՘t��ǉ�Pw��x^���z���,L�;
="������:��6X��u�
m^�R�i.�A*�a��63Ū�w`�E���WtZ1�i69Ծ�\�۱2����Qͼ�%'�pճ::��ջI:�jbZ�x-D�iϧ
��Vu$�p�.��;��c�%���Q8o������[�}�� S*�����7S���x��ĺ��e��ޝ�,ދ��n��K�d�8�zuj"����\�]�^�L��7�C���#Չ�-<GZ��3va�"iԈo�ۘ�+��Z���v�*�l������,����wP��m�a].ĒA��٠�{4��w��J�p��DH�zfY�P^F���R��ĭ����)'V3����:��+�}�n���C�W���	k����]w�ڞ.[�'�aʕ�XGk�ˬf�om�CGrho;�܁�K�b�հkt�D�$�k���x���:k��t��I��wu���|�_p�ؘ���y��y�0U��\���g8�ݼA���h�t�¿�k��t�,���"�*w#g�㛷$���Қ[�H9V�.5f�e��d��<]��f�a���1%�m�EYթ6��nI}��-�}�з��ak��z�����2�{��dv�ѤE]�}��\:�0U�)�ޭ�U�1�F�QU�a�uhz*+E�y�����/�Is(���ܳ��l�r��s��*�v�����fl�\�G҄��>�RR
�W_��V)�	�`��L��X|����<�� ùv�3���P�[����=��v���]��Z-���Vy�乪��Ҙ���#�Vm	�coh��u��R�׷Ekõ7���;�+p��P]���+�=E[�Z:.�eJHA����]�r\�]tnj��f��w}Ւ�a�_n���a�q��<��]5ui �5�@c-��;�~ݸ�b����.��QWԯ�Ph1�~8��.Ir��ˑ��K��Ź�s�p�S��Dh��F.���DW-Ȏu�n]9S�;�1���Quݍ�����s��;������nU�2��%$b���\�ѹ\�j*�r��7J��̚�.]���`ܧ8�m���]�;�Z���;�˚�uڈ���v9���Z�e�S����kr�F�'Eѹ��\�98���
�uʹuۦ9E˛Ar�c��˚s�k���scr��������.u�.\���ѺS��uۖ͝H�ʹn���u�b���wv�gqXܺ�û\�;���w����wwaݹ�멚.�7F29���ʻ�wb� �`�o3�P�Ӻ39����"��g�|�3��W�
��)��:)X��<ˬY��6�v��n��ɴ����F���c�����b{W����'� ��Sl�:�4�)�ڌ2`�V;��O�ڿg6�w#s�ts����v�(W�pO�#�Q��y�:���*�g`A�^��+\ץvMg'@jE��;擇~e�t�ÒA��~]˓�������v��u�d���T�7<�=��!��<~W��N�.0��=U9��pO�/����<����UI�{5HW��y�6۬}���[~��졍�m�8�J�޸�o�Fb�M�Fs��C�W5)bU�*&�1�s{��)��(���Ci�eB�7_j��4&��M���վ&W2rm�s���/9	�|��e7%���m�ޯeY��uɼ}����]S�ѱZ˹�צ�A��(O��EL��s���W mm����h��M�����U.z��	^�j��i��ok�D�0<2��{[Y��V-���+;;�8RW޹��w�7�fک(g���*Ѹm�%+f� ��T�;����{�b����d�7�C�u4�a�W$�evF��7vI�������y�)ƅ[�;�r���S��)^3)�B�y��q>[+�hk�}��Yy���vv#ps�<�I}^�@��%I]�t��;G�.C�9�v[���r5�o�Z}~+9
��lF�@�*Rq�5qx*�]�B�kL�lN:5��{~��ak�Y��w�R�� �j:R%�Y���n6�]�J��-��e��5��͡m�S�J�"�fe��b##�E'�_t�V�*�-��v'�Ŵ���V��{�^x�:�9����[�39|��MDc��b��V��qJ�q��&��o��������+2F�re��M�gf]�9=�h�g�
U�jV�������\�	U�#U.R�5҅����X֢�*Q<�D&6��5<�x��R�S�bn����B[����R�s�@6ƻ�9��`�1kC�m��Ӄ#q"݅��7�(��.�io���R��u�a���m �V�5��n��#�My7�]E{U�보 ��^��9C��Av,��Ӫ��{ �m�:����>�{��i�J��N�ӆ�=6z�yN��ӹr���9pSX�X�n��+�R�i^��y6�F���wq*� �c+���R˕3�$ṽ|d=4Z�v�#]:r��yS��Ȗ��l��k-�9}x��k��ǔ �Y�7��'�Oo��,�֖��ϭ/n=����g!#-�aL���\q���b� T�k���������n�|.�辡�梶z⾭�����@��wB��,�T�j����Hj���{����Շ6��d�H55�S,��Ė��]�EX��QA����X�ٶ՝gg"3A�>��.*/^ΜKH��G�璮~3�����bt�KqV�X�z�->�}�v;�h[V�SW!U�E��n9�ї��t6��Ou��a����<�{`�ol�4{�;�Kհ4	�F�C��+eBR�@���ƻFs���O22m�K��fJ�4gD�c�W
@^ސP"���-�zYo�ֳk�*�E�u�I��Vp�&��Px�ӪSH;ˤC�
[�����7� th���v[]n=�PM�~��V��]�ה:���kZm��,H6Nն٨��nS�ZϷ<c����ST<���^A�j� Ś�����\u��us���f�7�p�ǐ7ܚ�d;ͺ�e���xDWeᵽ���.L���3z�w"���^snh#
zWTl�_EE�O~�W�g�K��-�%q��U���C�9�&��mÿ#�U(�GpA�%b5��9�F�k����X�&�s��_y��i8<c]��]R�n�ñVy����U˶l��j�n�ne�o+�V��V�'SB�כb5rJj+��oGnVg-o�]O"I��0ӎ���3�K�3����Z��=�����;�R��X���s���D{��i��zA�-eY�ߪ�U6��VFX�N,m��M�9ݪ��w���a��g:��c͠��닼*����Ez������J�_�;�s��)�[e	�ӿ)��d�]a��}�6���3!R}lm�9��p͠�U�*z���X�P䛋����ʹ�Vv�U4�Vo�CO��~�*m`��J�����	^�넣E��,&�X�϶������)��̲p��cɢS�8ˑ����v�Z�3]Bąm]��jY���G�ƚ�L�����Z���FW�,�>1�\}2��N8m������|ĝ��0�]��cq�[aau���e ��m�����{�<�'%΢�W.GەƚVS�LWL��;h�)Awu:oe�2��ꭈ��j@�ʤ�V�9V)*V4��0�I���t��eq���S��:X�ݶy��\)b:A^|�IK���)ieb���]��yz������v7����9^N���R��>(!'�K���Oc�5'��K�1��'f��f�}��ny�Ͷ��ΩMyS���OrR3���cj��ꉥ��u݆WW�wt&�ޥ���m��T�0���EdiBsz\r|��D��I�s�З�,��r歗��P�X+`���o]�����ŔX�썹/\Е�5���_y����p�u[Nw��Ss�Z�ZB������_���?�a�~�/�t��U�e��q���{:WU����&��Y���f��T_�*Jt�����dDl�v�iÓ���<s��Z_5~sC�G����}~����o<[�ˍi�i�N�ro��	�C{��o6X<k��c�g�����߸N�yL�s�۷��ERw��9�s�]�B�a/J�������alj�(�����K�*��u)�:���z�g�|E�xp�ù���;�Hf�)+�Ҡú��z{e;�ae�'��vtm�˷
5����4p����{|4���U�k��GSg���u�h�>���n7-\?B���=�N+�Z��~�y��Fl��Y�Ŕ'�L��˿;����2�\a��nO�5����@vy���*���Ȋu������]���a����2/+}���Uw�ϋ�8Ne���/��8r>4�ތ4������ʐ=�*H�팢��կV�==�rC��?}N,jڞ7g�R�!��_U#u��K�j��[�/tz�8�u�n��������ܹ����S�q^���m�Βt����=P��h��Ug�ѱ=1}K�e�ﳫ	���t���rY�{p�O�)�c���/�R:	;�(	�>�W'�P�����a�*S��g���_��ޥoO��eizJ9�<녡ϙ} �iAy�z��ps,��8�ڨ��T���5 �T�{�n�Mķ|0{�;\q��;y�����QoG�ӕ����E�@YPd��S�"��}>�P���}-�C�_��܈N�I\�EA  &X�y��6�e�Q4}T�)�2Q�"�:L\�QZ^{�BW��#E�&���x`�4Um��O�;��~��7v��vz��)�Sk)���8�a����&���/��JL�9�.v��/*vԠR����d��qJ��)m_b�;M�{�-��Y��x_B�>��X���p�ݝh�1,�۳'�u=Av�ͦ�s6���60�Jp��K��d$n���O�3n9���3�;J�����f�CxzK�=W�Ss���0�'�dB�@��(�e3gg¢V�
�vNc������u�t��t���Z]wF���2m�@k�UC/e�d�L#�P}(n�wMc\���G�'��:��b��n��j��^�'w�=�S�~r��n��Ɨ�|s����[}Y7/p��M��/�	�Nةxp\W*�wѻH;�ܻ�ǹ��G���V}��v�i�\�^{L�.G�U��h�s�x'0¿�����*��Fu�g��ˬ������,��%���Mv�;3�W&/�<�:�Ow(��,�]t�mᅯ�x *qrĚ���c�~�{Z�/���t�%'�j��j�w<�Ӓv�Y<0�g�v��"�WSkk������zf^@��XW]2o��^Өl���k|��:'�Q']%����~�CÑB�6v?Z���=�O�����ɋ��P�7�Յ�.�7�A���ܶzZ�{�Vq�G��8�5��wV��KOkP��ں����凕���v�ֱV.��,��k��q$w�P\Ӛt��66��l�2����[uպ���s��6����� ��w7�W֞9�� Vl�΅�]o'Q:�"�8�����/:.OC�����	��n�Or��/��p�wO���ᑷu<n��Ĥ���8��Q�m\=�ǨKq�˻9���B�Ps�6,�.�K�2����$Qr�O��Q.���);���h��'�u���٪+�vK<i������H��a@��q6J���
�G_ʄ������h�y'^緽Ǣ��ޥ�q:Ѥ�s#5���*r8�MArDĥZ�
���4�cM[�:�\M��b5q;H���Kg�`7۽��5��IB��q��D�{�.�u��y�����Щ7����S��.5˩��N_ϡ�����؊Ͳb��sӵ��7�������hE�߃���J��r�����'R��tb�N̛�����j2/�.�˽oU.�m[2d��Iu��%x�K���OM{6��UV�I���r��t�X��G���wc����� ���/�yRl�z����1��0�t�/����q�ylv�݂��ɔ}��X�d],���*U�p?�i���й���@��������^�p���m>�r��S��(c���u��P�Y�X��ǩ�,^�ow��ڎjp��մ��k50+[tgu��S���z��dQ��M�Ô�k;���Z�t���8<��>'x6'|�z!:�[2�G�v��e5�al=�arg�̡4����U��go���.�Zf^�S������<���s�>��`���ex�As�7��]/у�~1\��u�>{E�L�J>ɗ�=�\?D*�L�s�s����q�o���L�/�Â��n�,��`�ϵ`=/��gGI�83�N���P�U�n9Re�.[9���5:�c.zy��Ϗ=�~�uuE�g��\c��=S/��j���i�x�@��\19l�Ǵ����x����m�cm�Y�.;������0��=H]L��n�^��b�����Wr��5��Qչ�ߓ��?���s���<�Y�x��D��Ό��/�Y�bv.)#��'������E�8���ŷ!��|��Zo�R2�;��ĪR ޚ�(	��T�S�?C[}���h��8yV5�O�'������=���|��uh�$r#��=�h�;QFO���7��h�kA���{e�up�Jv��9��G"��7��ۇwlМ�~QZPE�͟V�6�̢���Q�A�hJ8ϟå���G�9u�����,���% ������w�qfo�}�>(��T��.���J�9Ȧp1����RL��A���r7�vھb�w���n;�%��o�[7~۬讜Ĥ��'`���Cs�ȇի���4�7}QK�� �c;i�YjZJ^C9p����c���[Xegem���$н�Av��e��i��H��"~��I�L7�w�+�[N��EvMgJ�+���7�t/~W����ٷ�j��嶶���y�3�k���`��A��N�2��`��x�g*�.����8�ݻ�G�d��p�Uѿ7@)�n�_�
hV���Y;@�v���dS��$V,����[��,�Y�/t��R��n^\w�������'Υ	�o}b�����x�:�߀B���o�\��a:u�%K�p��or���*�zc�ӊ�Vk����~��l�3��j4f�?����R:�|_�Ϝ�
�d�w>���u"s�Ԁ�>�c�UI����Q�Cuc5Q�K���ӱٕ�Ր������8�w��U�aq����)�1,M8��'n)N��tV\����y�ZQ��/�mҤ3O�9�p��ʝ7��Op0����)s<r6� �������m�dy����x_�3���?�����J���#v.t����4g��|^�#aйQ������L��'��-wp�9~=�2��C{+�j��J���>%T)�Iڙ@w�n�y0�3��&�s�}�l*�mVt�j�1	]�@��q��]f����ZN����@���sw&����tO{���{����Ms��L�-gYu�V�_]�d�͚���ۼhT�yD�WK��m�ۼ3U0ݺ�j�[�W�d�Ep!n�v�1o	o�Vֱ����c�u:i���t��>ӳ�h��t�~*^xj� }I���fPi��^%���j0���B�$�ź�I�B�x��EVq��L��ObtI�����ӡ]�<0EX+%��tk���횅�s�E��x#�9F�mM�٫�v�0���Cς�^a�򴷍d��gv���\o�9��Ŧ��
�]� y¸h��'YE�/Dp��l�#���mD�R�t��8k�5X��r��q	2��b�P �]�u�u��ێ���s�֙�:N]w���Ω	���"�v�
JH�&��%��rgQ�:��ݸ��lϜ|k��gs즕��:�J���7��v�k�BFz�_$m����� ���-4�k���}vO��yGYxဌ�{��{����u���;-T9]�"�w~K2�ua�k�ݡj�t��;��m���ٷc�tP�m|��ά��
뗒Y�:Z����������V�p˨����f��IwPj4;Fjsy���wy�S�MgAl���+6��不烈w5:�e�Va��S��T��͠)�q]��L�sEn>�0=��C9��Sʚ9�Vr��xo��] �vm��!��\������̈́�Q��'+��V�,�'bƩ��/3��Z�*9X����X&۲��M4U&�7��j��β���h1��5��rI�q�4��\ׇ*wKF�K��ÛU��g��[����)�ąi�m+���8��ot�\�^��pj���6����]�X�	�y�\�a���x-��M��S��j�䋗uOT�����,U,���t�����̃�E�9��Z}�
8��1�´��u#b��-�/m�B�t�q��u8{��^r�m����ꨕ]��΀ڗlT�R�,L�+��ݜ���W9��Y�08�l٨��������K��P�t	YF�g|r�޶�10��MNb8�Ɗb�%��2ږ��ݜӊ��iv�)�����Z�g�5y�i�u5�Gʭ�$�wۻ�xu��,�` ,:� �]�̽'�7-�虸��G3p�,
+�į���ON�� w.�����o����SO4��c�W�`$V�윴]�/����A�ڏ�&_�?�b�H.c�)�n��j`Y1ś<3�V3���Z�]���7����3��ڧ-�z�c�2��ӅN�v�S���y�QV�AM#+	���mnvԝQ��w�Z�v*�a����@�i��Z#�g7+�i�bE�!��G��9���`�3�eWs��LQا�,M���ulʈ&A(i�n��2ӽ�/A{�
A͒�!�p��@�:26
Û���p�j��wd����@}cS����I�W 74��wls��s�����]�wG9�w.E�����M(�]اu�:ۮ���隹�\9��:vnT���ct���ۗ7v\�Diݫ��Lp����F����7wW;�Et��U͍������ܸ�iˮ\��w\��\��Wr�j9s�wn&(4sr�wZ湹�1��1��k�l5˖�tss\�˓������*㺸TE�H�Fw`�ȍʹ��������Ɨ*K�\�s������\ۘ�����]u�uˣ݋��鹷9��s�Lntwj�.Ph�ss.��&��-ȹ��#�r���:��r��3s�;�\��h|h
@a�ѨG%���N�ȭ�A��{q��l����ޒ�h�4h�ɋ\4�,�;��������e�ǔ�a�B�Xz�N:���{�S o8u��?���z��:�ea_=���θ[�.���Gپ�V�$��yc/{�����ft	����<΋��I�E7\&�[�=��9��8w��Lf�9COxO9�c/#TU<b���q��2�R�"��}>��:��D���5�Q��U�����%��9;��}v�)Q�"����;FB���q�K\�3y���\��N��37����WR%���D�Cn���q(�3�����!/k���nj��}�J���-���="�e�Q������p/�� k�5�R�@�t�tS>���,)!Ԁ�+�kkP۱ڐ�R����7�����������2m�@k�UC.6_�MDt�=+VĪn�٪�gnD����<��
r>�T�;Z��^{���{a��]��K���T�ר�Et�MGk���5��}���L�ad��b���W*�w۴��˼{�t�����s�֞w�-�8���}���v=W���_�|o�fc��
n^��XgR z�SV7��*<�*+.������GS�i�����xsp�xZ�}$�i��Y�P�5���MJ2�˶T5n`Fg9�/h=z��oP�GX��ņ�7M��7��K������0Q�ة�Ր|v�WI6�s�P�8k7�o8�+X��SwbC��Ή_����?f�b}S�z��ySjY;��!�~T�ʭ1%�Jx�6�8e���^ 5���.SrT;�����p�s��q�9'h�xx�g`��uc����Td�1}�У�W>�G�zG�2�+��Ȧ^+w��5c{ ��8�j���~��OR���$�j�D�-xn:3�%ooq����&tm�L��t%�'4it������n[=�j�����)}�<w޸ɧJ�Y޺��rg���Q�\�q���>��s�J����\9C��Gs��+v�}���q��m�Y����_#��pq"���}޺�wI{D���	�{)�j����j�ͬ�I{e4���*�p�'n�� zK5��f	)V�q�=�R+V	z��H��ȿ�l�׃%|$��A��|u�����HۇwhU����t�rD�U��j�|;�ٓ)�Պ2�Y}�S�5	��ƣy:H��ϴ�r�`7��ͳY�%
��\}�Ï+h���r>�l���T�G�ѥ"������_�s>d�B5�R�D�]g��0�!�f�������$x\oK�����e���&j�@L�4l����M���o-������i��6��P���M�}�v��������0է�vDU�M�3�bt�̽�Cc{l%�y�[��\��M-��աT�5�ۖ��[*�w,TcUoZ�n�Ⱥ)���9��pfcl��J�f��9�5yԴ�9���1m'fJe�ǻ}{(D���#ڟ{�!������P������m���vW��K�]�Hmƫ�<����GST/�[ewb�V�s'����>~����/W�y�U�a����2����������H�U~I�^���+�:�7�K���Ϝ�S���X���H�O��̘[^��{�9�2=�>�=�_Q�~'iH��-[�US�|�1�Ns����<���\�O����^:a��+,]�.�i�'·�L�qS-���2�{��}&y�L�����5�;�7o�8{�?�tq<U���_��E���?��:�v]iP}>ɔ\aV���Re��M�������A\���5��WxYsFy�O����t�$�9�j���i�{�.�"�ä0å]�|+z��p�W�����8Kը�mK6,�'����T�F�]��O���,]RʫB���me{q.��%��{D-���q/%CQ�Y��UD��x�A��]�U�6�:��MO�~��ԯ�UyJ�מ��)C����F��n���Y�]n��W2��Y�q��|��8�6D7��t��L�ӑ�O.��\~�Xڱ�˯8�Z�� /3xTO"�f����B���[���؁�ˆN��vt&j³)�Y�MHk���Tθ��U��n�Ds����KΙN����)���U��Q3�^b7r�лc��,�����R}q7-�q�=����n<ݑ��ѫ�L�������8�h__����s l�u(6 ���PZ+Z�%�m����m�s9��n�v9_V����=���כ����c����H�y�;�d*G�rax�>߇K
���#/�[z�������Jv���_oֹ쬯���44E+T&���;bf9؝��Vӣ!w��҃Q�\���EN;z�9���:�D�C2���n0�GJ'`���ED����<�Uv��OW�>����c$[��������]���
n��耦�\k��<Y=�ñ'�wt��Pt"ǯ=�gM�8�¸�=�i�v��X]��1:ɸ�;�'|�����>��X<o��1ѻ�������#���\W����ZN�F�or���*�zc�4⹕�F��=~�y�/��4{���;�}kdΟ�Q��X�8�I��k���Τy���O��Z�G	r���=u��V>ʏ�ا2���+���H<O��1V�0j�%Z�K�9���{ռ�������˽{t�ֆ��t�x\�49Vn�6&\��ժ���Sj!�gtB�t���.,����֮*�s�ݰ7{w:*���7>@��9�K��)\bٽ��Ng��+g�N3̭��?�+�����*@}�i�T�j�}!+9��ǲ�|�.R�������&W��\3O���y�S��{��3ƾ3�
�W� %�hn�c�}N.m笥�ٝ���싌r���,=_S�q^�ژ�<I�W�
������슭�o��;���}�tv���������c���|�ᾟST�z%e�^���:	;!�r����z�o:1X/��\Ǥ����u(�SBsR���k����Qۇ�p���2���-7�����ݫ�xv\V� �y�g@��O@���uJg���r����x�q��p�HQ����""\����4b`�UV�FIF��z��AKd�'�O�:P�N�h-�AWzwdlw�Zt3Ϣ�w'�g��ۭ�n;��q��R��@[�	�`�鶴/=j�����%��Szwَ�o��Ƞ�|���n������mր��J%��@2#I�VӢ�H����d!|�r[����7�δf=�%���i�`hO��WH�3��3)��wW;n��h��������6��|���(�X�j4bG�vm*�j	��wZ%
�;�	��`|i��
�@��8��2�J�[�N��{:$���3;V�N�k��|8j��:��2��\0Ԗ��6$a�~��f|9���[74�r��=ܮ�d�p>����>��鸍��UG���2nt�S#�/�&��hm;[�tg�����lt���V-�/�n�Ӫ�P����'���r�ꎅ'���y�g�$��z{��,���}8�R�ฮU��v�w�w��s�ދ�R�.{��RgҎ�Ε9��^��~�i���.͟�V��(��c�}s+��S�%N��@
�g@*j�&:��v�8u]zr��(_U�#��R��ʘ�~'3A���?*�Y��-����k���2N��䝃?�� y5d_�N�rq�F������������:�����k�#�_�9��5y���zzg���*GIpFL��)������K�f�[�3���%��5	�F��t���E�MCX���*e���ڡ*n1:��]0o�:�>����C�/�S$����/=ڰ�	*h�/�� �<�/�S����)�֕X��N�Ѯ��mn�7ɽ��#�Y���ٝ=��g�4���]c0��Q���OQ��D��^�.�R���s��h�����4v^)n�o�,{�x��ΘE_���N���]��ΐ��j89�K�|�k{�ժ���u�����YBY]�8��$<C��Su�s3�͇,�_Qܓ�h��u�[t첀�c*DdIoq	�-$m
C(�m��.�U���ۙ9J(M捃w%_#�����j��:��=q�\N���If���"�u��/��m}�v�z��<�<5�q6_݉�Mħ���/���7Z4���n�ЫS%O ����FO)� e��_P�c���Z�ݦcܝ�}����9��[u�9�f�)�P��{8��X���;���et����ަ*���������q�ˎ]n����%�M�_B5�g�!�T`+q�y���W�\�"���ff;�uxTK�f�Ӟ�W�KM��Ά��Iْ�xhV�ޢ�y�<�{v����h�dWK�x2w"��	~1_J���OM{6��UVi�偐"�2��G��s΃IPS6���
�*A����[	�1�N��t�/��=.Z�zk6�~�t���)��^�W�S��N�3~uaN�y47�T�^J'+�|72�W���T��Oç��6���>��Z'�O3�J�S2�҆����c��؅s�>���bxQ��؋����xl˯g���V��d��T�5p�<�'���{�ڸ��G;�/�S��+#�XC�G��U�[%�F�\���yl����K�ݧ�{6&�tu�gR�r�-�z�VB풎Q��*�U+__^�5��i��Fz�ɯpp�H34�֧3T�N�����a\��gN�;��v� y�qdιj$�U�\]Q���u)���oT��s�Z�'�%c�'��e�P���R���>��ވ­�qʓ,r�͏g�7�=/s���vb~z�x��mO�ĥ`q�S/�ꐊ�d>�t��l�������]���-/����ee}J>Y��Qb^;���ߋ����)��f���];5T�)�u����b�"��2����D�s�=��Cv��蕕�E��B:I�a@��������@��6���c�㪸��]ĳqI���D�o��!�ײB��:�e�wl?|�U
@ӽ���<=�H��ȯvS�4�Vփp��=�a��SڇKw�C6�a8v�<ݑ��ѯk�iP��u�JǇV�ew���x\GA� +�s��3��
��Z����0�u�~'"3�C^�&�Lo�����mc�I�o��"jD~�6��f,J�f�T�h�Ã=^�՟~Ӹ��]��q�/��%�1�^�t��W���J��l�^���ϻΔ�[����D�S�5����r,8z��_ɪd�B7wR�����?�ӥ�y�)����{�C�@��EM�*���Wb�x#EU�**�������On�:�C�Rݷ˛�&_�L7Cb2�e������y�T�?9�>V��'h&�+	�7 'Y��r )Oo��e���ø��V��Қ�kr$%����e�h�����vu���{�)mFaz��mUѿ�� �۶��
he���<Y=��-=�����S�1��<7z4�<	�*Xn+'t�9�wJ�q�yqގN��:�'6�X��3q��莛��Uw��W}K��gg���N��1��u-'N�L��Wʦ����8�edk���C|Ŭ��U�<o3�~�=���6tV���>�~��?P����N�]_��Fu +���CUI���x��{�Yw�NZJ/o%�z��o��{�2�g}��pf�K����T���鄆]�v�S�����_;t�u�.)�g�N�f�|�����qe��fax�څt���^��.���kfN03�����إ7;��ާ|�J��~kjc��$�%|Y�eX?UJ5}�`��s�q�(�a��Y��+�^�.�Dc���=�o���1މY|�ģ�b2�z�F'��U|�2��q3�HݨrJr��z�Q����jV��5�ei��(���:�j�s�w3@x�Hs��ƾp@�FX���ZS��}t��7\&������\@�n�cx���`i�Yo[����S'}��4z�xn��<[��$�J�t��|o��|�k��8j:�*��2���˃��a�]�i�os����^���|�;�a��v��%���A+N5s�Mt1�f�)��H���l6񸵾���I��4���_�wl����k��A����O>�{�҇^'|4Pc'U���sgs�y���h8=�hn}��7��Nwn�(�qT	�bg�mK�^�cl(y���h��_f{�;�.&��r0.]\n���g�ۜ~~wQ
e���!#gd�#t��V�׷ܕ}�+Bg�R5q	u�-��[��#XD+�GM��-���~��tZX��c�.
�
���W�O3�o:V��{p��j��O2d��|P�P��V½�Y��u����c����tm��+���ชŶ��v���W�	'U�:#�ro���Մ��������r�ͼ��8�W�m��Y(ah���'�9I����_n]�b}�ת��{x�5��EשÎj�)Y�k���w�ū�O�O��k�0�z;�Ƽ���Oz�I(�[�����m� �.�=�ރ�j�9\�m��<��V���������^��x	��y{�����8�mS-�K l{��/�I�8�WO�Uý�o��gNIۋ�O�� nk}ճ@�U���q�;���բ����f�A�>���i*�_�t��xυ-o�G�5E���Ia�� ��n�;/�}ip{�u��&�
K�o=����b��9�h44XT��[/f����L���ݩ1T�ݘ0j��\�b�pzGZ+��R
��8[4G�;�Z�t��j�+Z��"{�*kD��jIBIpV�M!�[f�-rO��f�c~57� ����^}j��7��N���=E/*���tO�VHy�Y���3UrPZ�\��e�]7m��ux�1s-���mG��b˵��C+e��9�uJֳi�J�#Ji��f#Sc��1��!ܫ]\V2���C�����)�7�R�[Wy,}
=�Q����k+/��շ�p7x
pm�Vi�b��+��kTDm��ƻV$1�����Q��V\�*l���B�թ��ۓ8��ʢ.���M��tr֨�<��0���D�ͪ|��:�m�r��a��N��Z�30q9�8�� P��Ê�_Y�6�ʳ1�L,]�&ou

EF�5��$�֏��y��|�T]gY}��7�9�jԺ��鐭3s^�<;�:���o��8��/@�m鈢CJ�i��:��;Y�톩��Z1�/9|8���J�� e�QG�Nv�^�`��H�T��	do��8�1J� �n<��}(��8�ٕw�,R&��"�h���l{�Pr�����R�}�{�Ō:{���V��G�B���b��c�z5nY]�+Dg{�������e�����:|�[k��1r��r.�m�;M_V9�ZW��A��j�h���Ǘyʵ�
��sT��K��d�n�v
��q
�w���������+�yD2e���8:x����*��'f]�5BV���qŜ�Y�v
k�u[h��,�y��k��t��'-�ɳ�^U2�_sWώ��Ⱥ7���Yp�C�����Pf+�����s���F8�Q!\/�kj�i���AA�g+Yo�i�a���
�h��\d��f�	������=�4�k"�]�̓{�\@��j�,�W���-�ӵ>l��oB�WY�M(fY��\Z-����Ӕ|k/�Qi��2����n������y�t�;-	yx�j��3����N�0;Kl�Q"�M��׋������T��n�	*\�	ZÇl��5���.E���z��y��+J�\���ƍ0:r���=Gt{�Rz+g�;A���9�w��@r�a�]��M0��Ǡ-{�6ɛ>�Io2P5qG����1���t�GV���X}�������ެ�(fM�F�!��Y�J;'��{��S[2h9�łwf7�� D_Mv;�qPH�.��G�Գ9K�u�2ۮ�9�!�SU��ס;J�}s�,���i�Rh�.�[�gf��%���|�dnV�n=ܜ��u����u�eu(�{L5��x�V�w��؜yl�A�e������Y��}��
���xo�p�KD�}��PP_H���vw]���#.�1���]���v�;��Q�t�������rnWI.Yݷ*9ˑ�#s�rw4��Gu�;��E��nfssgw,9�i(��ƹ����[�.��4�!s�t��Ĝ�r��n;������Ӝ�BF�'uڂ���9r7K�볺��湢J�ȗ\��b.[��u�Q���nȱ�9۠��r�Rsn�9�(�w]\��˕;��s�wF�ۛ�&�ę!r�#\���\�Mt
Q"SbILw;sD�Φcs�7,U˻����J��vs�FB�;��;�#��nnY2\���$����	Δ�Wwk,X�����:z��D�nD��Ŝ��j�8Y�����Xﻭ�bpE{Cn�]�z�"��w܎>�з�-�ݛaVU�k�gwv�����QZ�ϛ�l���p�atɸ�R�{�n�ފ}q���!1��⼺���.���]]S�4+	'\�BgC�����ڡ*n1:��9`��tX|ܶ{��v����Û�׵{�=c\u��4��,�ײA���A|P���wN��-*�7������
�^9��Z�졑��?�Q�	���O����Q�t��e?�H���.�w��_��tDң{.n}=�x���1rА�Z��O)�����:�p�'n����,�" oQ�P$�ZO�=� �B��u4��+����eF�x�\M�-��z�>;��h�^9���Ы�2|�q {��6��C�)��{��X�D�փ`�+�&�ƣo������Ke�����ͳJV�@޴OO�^�S}o	C$��g����]JӃ=��L�.5q˭Ѵ��,����Ѹ�dᘚ�:B�����3��@y6����G�f���R�Y�qN{_�Դ�o:��!��tWw?ޯ�@���4�fH{��_��s�;�f�����AO!�?Y�}��і��}�Hi�U�л�c<���g���+�����lJS鯱v+��b�B�3wG���}��8�ҭ�����\'~�}:�S�W3�d�8�5ٜ�(�+h�@� �=�d��\!
݁�:ԝ��!W��q�:�p�n��3;���pЛuq#ʴ�7�йz<ϕ��tͷ,��Dkʐke��=0��Na����ax��%� -�}ے���9��cF�z��uO����37�V췓Cz�R=d�r��L�q����U����?���=N9�:�d����gKf�rձ�UOI�5LsS�����h�W>��a�5Q*�g�]�<m^��h��eᢧc��Zl��F��,
�5p�
��,��:�zWէ|p��~*@2-�U=�V��c�fK>���=P&tuԺ8/�J���L�:�
����O��G>�,�3��/�m�'c{<��d^���v~%+\e3�Ŋ�|n+UW����)�z�����Kי����vGN�?���K�B�i��*Q����>��R3�r+��w>�q�����t��9�_����^�����-�C�-�c����O�VWJ8��z��!k#��Lª�U�^|����Q���gt�/]ĳqIm��JV���r��=���2=�ݰ�Y+b�A�^2���}�d/X`	�q'@�����uX\}�\Mķ}��ϙ�8ܜ;y�#+_���gD��{��/Ǭ���l�C �ڂ�ixm3�ה6恰�mpW'g+��O35ɀ_l{*$|u��
;_�A��O�����S�����|Y�}Ǖ��4�&�c��_d�z-�3���]m>�w������'͞��%��ͫ]ݽ���F?��i��_��.�@r��L�����b��ޔ�#������ݲ�q;U����߷�T�/�N�v����uI��DĞ}4/�S��qav.��跎��~Ǚ��)O+,��"W���
�D�Rv�%]���V���3�}؞vZl~G� ���O��zǤ[�n�����*d�|̰5���+��rt�v�B�p_�:\bwf���{=����k�����e��q�����ګ�y:Kt���)���� �K'�{Hw�ێ���;�P=��=?x�����[����Ţ�zX����O}��M��t��yt=��vN��^���.���<�
#Ŏ������c.�����n�f�-\?}
����4⹔���&yT\�}����oƜ~w��6����m^%�1��SV�	E��'/9�Y�ކ[��S6�4��y��;�������x��j=���o�]����N�{ �/W�_/���*@}��S��X���s��M? �b�[���9N�=�u�4����\geN����3ƾ3��Ϛ����lM � 9���}���Z��JG[`�چ��ݛQ6��o[wJ��	^������֦�=�\@����ا1��/뮣ާ~��*g.Ee��-)췡cm��"-� �+iZF,K:���7+��v�,�r��UG$��6�CJ\�8/܁ٗ~�/F����i�eք5���p�*F��:I�V�U
�B�������.�F\Q�f�ۗQĪ�tF�O2^On閥�蕗�tX�i����c���ܲO�d�$�L�T;������Gi*�7��oO��rZ|�J;�4��u6�1�'�=CTm�.�J�>���(	����@-)���ϩ��7��|0,g�)��r������ʏ�;E���;y;���х���}�@ޣ 8	l��y��å,jX�ݞ~�N�ߣҐ��u���/�hn'[���q8n۸�FJ<�t�<�h��<���ry>Q�}��N�����1��h�� �ˮ%����m����&�˙�$z��V�v�a�~���f���'����Y��9Y�	ԍFZ]n��6�~�i�5���] Z��5*p�vߥ�龥�3A��l���{X*�[9F�i��ͫ�7S̙7�n��ƉSS6X�z��==�W����v\Jp�;��Â���ݥ�Uz�l$���BM�hc�U����F����'�^N�Z_��/S;�<�nSU9��n^�[M>ONc[�	�k�k�Y'a����1\��G�i�݃����ʾPR�]�.��Y.V��X+�e���nT.R��gRZ�!���'�eJ,��IwK�߱Cs�R���7��E���P�����b�Y4�3㡓�=0��VqR�࿫�i;��Aؽ����3w]/go{ۂ�����Ի��n�9Y���z����>7�Ne�f9�	�0����������]+}�>�S4�8]hY��ǕS��5O���W���E��Le���wl��˄b�0���"k:8��d��.�['�K l{��/�I�9�5t�Uý�=��9'|�.��U�6r�L��ƮW�!�65�L�Ơ�T+�u\v����p,�G�X��6{�O�3X����>�v�r�[��Չ%�c����/d��,::����mP�7�Յ���qtXw�@X��)�5+gw3ú+��~�s�Q����x�;�Aڃ(	�BOOۺt��iU��BѦF�d���z�qף�����C�(��j��
�f�zJ5��z�� w,�K�ì�Z��R�d-�z�gO�V?1 ���a���>���\N���Ie{ �(c[�]k�;B���_����P��b}q7�{�w/�780�Hۈwv�"J���K��¼���2�KK�X����e$�F��d��a�CY�����{��]��Ֆ���Q����^�{�g��5�ݬi*.!uWG��ę
hPn汦8�Ѝ�G�αt���q�~�m�ػuK��+�ቦ3��{x�M� ,���y<i^�0��.5|��}g�[,���mށ}~���k��}W!�q�tR�=�gd���EJӃ4�F.5|�����,��̪{`frs}o\V�z��<��+���]r�d�uxWҧY�,��{�a�s!�7�M����{}���Ǣ��p��2n>N\~�F�"�e��<;af����/���4��YF-�9׻��w]���x-�ۿ��wC��S=ܰ�
�2l�z����1ݝ|L�BM\�s������3����x���R?�����/-�s�|}��f|悜�oj������D��(}=���;�U��`=�|\AިS�|v�V�8�s���UT��CT�59��^<��z��>���\{��!{���ד��ˉ����"�U���O�ʁ^��M&Y2�#��d�2�BP�:p�箒�»/dK���z����w�l�%�o����5�����]bH���`�8��(L��x��8�{��R����\f�X�w��S��{�����(_�2�Ω�[���3�(w�p��U�7ЋK��f��+i�R�ӨN�4+�ݝ����oNd]j�Ro��܁^ưٵ�\��铴�}�d�&T�������ו�X��jȤyv�����A�W��s���H=�%���qe��{��j`��n�w#ܠ�[�e�\c�Hg���z�p}肫8���*Q�:I�3	�3Ԇ�ץ
���6e�]����p�I�][���h��n��J���QCI<�-JU^���'�����r��E�Yv%�o�N���>�!�ײB���F_�ݰ��}E�z<��N�v�y �F�p9S�#�갸�)>���[���.|�il����)�{�6��td_")���.W$�F�i�|=��}���+��.�S��
���U2�77[�K���g��q
g0�����û�h\)��uI�d�I��BQ�}��ںc��٪7��o��ȥ�� ܾ�Ͼs8�LLz+U��;�f9��w�+�[N���e���P���ص�qK=��vil�OZ�\7�t-�L��|�� �ԃ�^'X({K�ݳ�|��Qmv�E��ջ�$����,>�����P����m�Cj�������K�d{5��Y�3~��է��|�P���e����9>t�0�d�/�wJ�q�yq��������&���[���-rӯ�Ƨ��ڵ��jq��5ց�ĕuq�~�0|���sբ�����ϩ�[ҕ����C},^�ש��b�R�mWs5��r�-<p�vƒ�ոj�[����Ô]�h�\��S���Km���g��|&RKsGJ��s[�]]���1��@�W�8���~����_�l�;�e}cԩ�:}��n7-\?B��������P�5�� ��|��u���Wx�����_���g�O��?��#h�������[�<�*S��=~��d]ی�5�S�G�Ռ�F��1q��7��faz��(]ZxS����3
n<���E_���� +�'hu4���-��:=�����M�e��+.j�N����7go7�i�O�G�*�7֨��������)�ܷL>���蕗��]�#v����g�����H�z�6\���?E|onT	F�1+�^�.�d2���7�覩���T�iwlvf��D�`��gA's�C�qS)K��ԣt�X��R����2��}}ޣ\Pݟc��oH��,�	u�o��e��Qϔ7��~<} ���uJg���(q�s�?)��u;�v�Wq�Ãk�9����w.ݣ
,�r:����H�Mֆ=�9���Vq��f\�,VƂ��~�Cq:�&�x�'��qV��k�"��N���pq��$=�]2a��ozf3v��9}�/[9�	"��l�Q"(��2�W#�x�h1ٶ��t����ڲ�@Lm_����BD��7�O��@��P9h�ӝmQ���?b�5��#�+^a)�L�ڥ���n����S�#�K��������^Vx��f��K�Q�sK�C5	^.���9uĿ38-��7�~wJe��鉝����U~���Cи�$9ާF�騏e�3p�5iu�7ۮ�� ��F��<��zf��矷nOz��mL�pfW�Ǣ^�
���Q��Zoy���.�f���2D�"K���b�.��j�:��/�&�a����Cl9�r{�V-�/�T��Ok�e��{3��5o�
��[싗�c{�zK�� ���囏��3�q���=0��VT�8.+�i;�b��s�_M;�+4�yz�Ã��}���o���=��*\͞ңvL�B�e݌�Qa��͉v��,Ү3� =ki����-K�=�hf��k����z�Y9�=�,Ř��:���q^.�B��V���O{ {��:\��u�}��ގ{|DL/!������L��N"���kg���d]C�a�ug�����s�J�#���-_��3��{5n��Ӓ%ǯ^��9'E��v�x8'B�T���T%M�xU S^�k��n,z�Z.�����q�G������0Խ\�қ�pM��Ԝs��#^���D"��i�/e��!t2xTz�.`ɿh}yсja|!t��̥���ՔȢ�C4s�Ȟ�R��g����3�����t�RO��Z&���)W�n^����7��)H�����O��=�Q�� �(��B����{wN��.��K�?D��5�w�z��z%�vƏF�t�z�GnW|Uc0��Q�t��e0q#�B��Tm�"br���vx���g�S�ԟ�H�����YM��p�����;w�=%��z����J���bn/��)�(rp��+���}����K}���S��h�o玤m���
ۆz�y����꽋������h�w:�`-.�8�.7��F�t�_9�il�9��Z��Q�螯پ��_�,{��F�9�P���?�n�)�
����z4�f����u�;7vR�j�n�/�c���I��}��C5�#H��S�ff9�ë¾�:�	g�k3�i�ߌ֗��^���|z�J�m껣	�fM�r�kBcћ/�I����[@��+��=����j��n�w=��MyJ���'wB��37,��+�~�'pzc�������.�$�3��,;������u���ܼ�=�NC2�ά)��{V.:�R=�DW8ə�o3&x�	w��BO�lVA��y�+��x��z�흦�r{���pݥ���"��W&�+����,��`�wd]Z2�8;�s����aR�湡Mד��
��s���Ñncp��f��9J�^���x�o����94t|�Q�a���.t��gh)�ͩ�d�f�5�g5	yC#E!�] ��qw̓z���x��.�K�]k�ŋ\��?p�rc(����i�pʔp�"۾�U��׸n\Oq�lD�^-z,�hct�v%87��5b����=6ie�o��	�G���W��v�ԥ5�մc�ug$�Z�,�q�����>U�8s��-_ U6�1�U6V�-3���Y��C \�rgnP�@x��g�;�4I�c��X��g8��`_'xqtT2Zg0l�J+U�&�#��Cp����wd�H]>8F�W
dP}}�Q�g��
��8�+��)�)4)��+�����0�5���Z%���:c�b-�P�(?�*;�!t�9��!�e�[��:�IՔ�tt: m9�����y!*7��;~�k/&ɝ2%onQ��_LNb�O�m������A��2�Y�+�wt�GPGb�W�^��/g&����*�@��r�gC�F�s��4	h���nj��'N旛0%;�:�Ch�\����\6�� 	�����j�o|������2�׌�-�z6�ƅj#_�϶�j�fU���,�ыRf��+�Ϋu �}���m�;��Ϭ��M۽2�Q�*Ș�^��(l�}�@r��]-���bҾyLl!�ˠ[|����:����;#�ïc�
k^���E8��]�ю:e]-�5h�r��Z7�/\�Ğ�l�95����lK��f���Vy)]O�[�n��yD����Y�9n�;����]0�gD��d�xU�QG�� �s�(7�h���Tv �\��Pytƶ�F�ΉS�ޚ+eX�S�e4��㝐��ʻY2+�@]7([�#]���\�B�|�KA�jA�dp#�JE}h�TF}�4�������+��}��ؓn[1�_1`�T�+hs�muq9���_S�e�	��^teE:N��fҙـTݥVNK�s4r����@9���ɔ��8p#��v�z7nX�8],g2���ì�P�YǨwn��>	�ܕI�i��;M�gN�o��I݈7^�u�a��:U�{z�;�ϭ̐t�33mv���&Y W`��]����k�ŕм����5���FN|�p�x��0R�/q�k��NXf"w.a����A�i�ۭ��c�5➼	���ڼ�,�v�α��ʐ�A��JysH��i����B��")��A�ooo��"�Ԭ���utډpw��E;��ԓ�Ј�����ҥ��cOwl�;Q��P�D�#dv��r�EFbЖvw�R\��p����ǝٖ�sŝ9��fA�ù�6�J���ve��}����k��v@�uB�������4Id�;�$DfRw]�룜H��+����q:n!�.Tu'8  �qw�6���XwrN���&������r��d�؎\
wk�\��wc��\�4���%��HܸR@�Wu�.W@.naݢ�&H���f�˙ݮ��L���$��wHŌ����!spDЦ��̔�Dl	##).���uۢ�A�v�����Θ�B4;�w"F��H�r2���s���$d�I!����G.F�@�be
MH2I;��u�7(�v���A��⸘��cEw7!e��t2
	��DI�$��)s�H�Ĉ�n������#��P�B�L�$eC@hSRh�1,*�UX��]×P�D�3Z�/p%Z2gs�
j.�Fa���<q�Į�,[҈S�⚻x����}/��֤}��v�:N�J�GxØ�����$�'�3�3�J�S2��T�59��m�͢fՉQ�sν��g�Y.�Q�6�J\��^��V�'�<w&TsU�U4�d���~�s���yU}/4������M�Ԯ7��s�ギgDs��.eA:;�R��J���FL�9�����S���."���Ni�]:H쮨�o�ޣޙӿYd�\C��=2�ߤf�l��c`�ױǭd��4��4��:1ä3�7M��<��Vq�]�(��N����\�7>`N��y�6�z}+C���q�t�?E�������薎{ ��A��Y\����(=��z�ћ}��R,�e���v��EL���]ĳqIm�ܥo����|��Zo�R2*��]F6����t8���'���,J`X=�m�X\}�'�r��|\����ڴ���3��L1J�wWI0~k9Qq�V�Z���4�}2��A���x{�eq���}��??;rc�ٓ��ε�+xzZF�W"�s9��Cn�v�ݳB��F����6�#�M	GY�z$/Q���<�۵�OH+��t�\����Qj����L�p�}B���X��2��'�I��o��''EJ�v�8�u��U��4�	A��j�.��yJ��l���R�.�,�i@:��G@r���|�gM<��;���\nVe.��Y���e�2��\�v�W��\?C}l!�r��>�3���j2�1>�.OX�����C���p|�X��ZW���w5FE��N1R�ԮC�]иiS%��`kB��d'�](�7�̋V!_�y*r \��6�����:������r�#2�i���ǛUt|�����`i~���OV8�14ӯn�}��� �K%�>��O�_�N��d�/�wJ�q�yq�����1:�z#ױ���]{��U�����6����/&}{,4},u������1�Դ�>ݔ��嫇kUA�&���ҳ0�Ⱥyf5tN������^ӿ3�g�����,~�8=>j����N��������k��<����;ݷ:�� ��ߒ�����E���_�J�x���亞c�$�f'3l#�\T� �	`o�Z\u4���t��S��������A��7'5J�����*~���`R���9��TX�<�59JP[*�!��Y|.��1�4��꺒�S��O�-�C�g�l�b%���y�?W�s\�Vz�7�uG��w�*�(�ݨ1��M��yc�y@�1y�:� +���p=y�R�����A|4�ڻ4E���E��Z"s���50^Ց�qe�o��$��m�m�W94nt淯;F��۠��\=w�V-�Z�t��]{�d���U�F_<OsL��FP��ܼ�
��N�N�����u2����7]�bZT��緅�]I��YC�i�Zrx�녾.�����J��.OPJxz��3}�� U�r�C/�W;�QrЗ����o�9��8v����wv�/@��j>� o�-�;e��0UR�Ο9��z2�s%8:�w�G��ՠ�!�	��7��q8]S��FJ5�@]<7�{}*���`Y�����a�Mmz��Eg��CX��`���"�IN����h�D��<�J���YS}o:e��F�g����m:7��*�n9�ԍFZ]n�nx�� �{�p�V����4iQr���Qofty=>+kIL����=��ᶪ���;�*FgQ)�_V�[��ޓ%��_�
�e���2k�鯏�����EOa�qX�ؿF�-<����̉f}��v{\틝Q����cq.M��6�,ޗ�|t2{G�\�
����u��j�z�׏���nl�z���q��a�Ux1���*_?~��؟����vl����c�nQU޿k��ق��x�]����0/��m3��{ީ�ӗ=���+f����f����;e� u
�J�fY��7;��9����>�mv�aSNͰ����K*��û���5{��6l.��6�.�v��6-��G��5�6[��(����K�q��S�_Ɲ`9��@
�>�=
�ރ�W9��{^����H��,�Ju��Y�WO!�3��YU��Ua�����F@rTF�:M��wQ������m��{����0+72�����_��1NI�D�ˉ���w��U�h��f\q]2o��^��TMVǂ�U����aq�6���3}�|�q���Iڙ��L�W��H��Q.u����q�������j#]�z����^����'-��5p��<�>��+�MDtW�_�����|%�.�4U�-4f�L���w��M�vƏF�t�y�v�p��V3��Q�GI=_@_F<��uEu��*���������=;�|�u���'^�SG��=~u����?@��n��L��_�{ڷ�z�.Y���H��S=��\o뉸���<_��܆�F��̌��3���������JwT@���i_��gĀRU��+K�	���L�o:�(�����cU
�����3�K�\rw�-Uc4�%��T����0_Ң��/����e3���0��j��
��Aڠ�5=�������g`Z����'|�j��i���M��+�=�j�pI��s�YˬK�T)-��_��<����T�;��eJ}��mV:	��x�92�M�H�Ԩ�檲�mCUk�Z����)��Yd_H��](�T\%<�g�g̗�k �Sh�Qr��R��>��X��v=��U"����.��o�"�YkUH�o�����'fM�.�#Q�[/�I�(���[b_�T����j�o�e�޺��:r���+��o]�!����t�e�sc���k�H5,��j�top�Wq{��ǜ,byw՘n+��}��Ƌ���c���؝f���|�Չ��9G}��϶���.F��D�@>�̘{^���������ҙ��VǢU='�Sԧ��U0���oww�7�4���yW>�덖������V���d��FL��_Oef�+��>I*ܟ������<��������x��o�8/��8J�::K��>4�>��^5�1>7�]֯9�^�i�h��MW"��*Hﾥ��N���kK���+��+O����6��[�8*j�ѥl�>]���A��3A��#���R��N�>�Y�.eJ7��$�Y�%�����jk�����gՂI�sn�^��b��x<�KG=�c��7h=>����'Fa��&7��'�j3Bw Ǫ�ȶ�Pc�)��$�hI��w��}�+=�t��'d�Bp�0߮�a���(	��[D�kf_%G�����Nm3�� s�}�����2�uב��3u򵊚ٷ�#Ƙݍ�����QcM��ieIY�Bԙ��v�?3ĝ�8E��}b��Vye؟��}blKV�����}h��O��8��yu�_�2ƹ�U��>%Ґ�Ԕ�J�W����aq���z[���D��ﱯA�	�B���*>s���O�8�vF[��j��(���&@s*�l�z8��Jr;ʔy`�MKC�K�;o�Rз<A~�H�9��nw��١jd�Q�$.��m2y����51{����v
�5v�u�^��[{�/������%z���+UQ�T��c�ԕu7�C�U#=��iGb��Ö�Q�<�k:X}�\�-���pҦK�3,~F� ��(?i���-�J[�?ӷ���:~�U/㞨�[Y��R9W�p��o=�=�j�����H)`��/z�&^>�z=�ʼc7J�D�����5�OT�����R�<g�az{�V��7/.;���Ű5IO6"�f������C������w�'~gn}��Ϯ6X<G�>b�Le�u-'N�L�U�AX��3G*|Z���6㔙�0���{Tp�^i���3�qŜ���?F"��pOVٙ���<~U��=��	�˻�<w���u�%lS6�����93k�ǡ��8���_�!�5yݵ{,R=L\�u�U$F1�ʺ�)�.�(�h뺫䮹�e���t7m�\�X�fCwP9af�ڝ��r�v"����)�9֩t#`ӓ���}�u���'�	�j�?e���ê`��Q��uq�ε�s8z9����Ż"̸,{XSyx�k:8����9�7R���L
�ܭ/���S��z�p�>���_��S�z��/D��;_��Oq������23 ePw_U#~�u��MPa{�-��7;����;��Y��3�*�Ỵ�I.���*G\\�'MIl��z�]|v��(�*��W��!��홬1y��n�L��n`J+3�Ǻ��.�_���|J���$�}2���
�^����O���c~�ƥ;߿O�u����9p�x��Z}d������_��(�B��A�q�niOm���S����zޡ�/�Fq׋��LM�w�?:ZT>��n<���wv�/}�Q� oa����@��LM_��[b酽�C�{\�����'|4� �����n���O�����\#%or$�Us�$˵�M�8����iQ�������zF���ա�.�����術+n��,�ݚ�n��	�>q/�*f�fGq�;$LK�td->��ێgR3�K�Ѷ�p.H͢�ɖ����^N�,죅��w@eF���#�6
�(�cʝ��&e�Tl7�CG[]�ّদԷ�_�y���N�����6l��OVΚ��r�j��I���s���b��:�*���nY�'j�n�ddg�+:��[�ddXPR���,��3r��Lާ��������k��S�h�2����V�
Ȋ��Q�+�=�s�[�D�����k7�n^�7:��p��5�*��]̜�zh�P�|�Oa�u���H��e�i?Ӓ�_�o�v�E��P��[�ˍ�N�z18�&��@:�z�}^������2�,����,)���T�%�����+�����"�z��'��>�br5ʌs@��^��O����ǂf�7=�����n�=!�ہ;��z��=8�Ԁ��ǕS���>r��ucx�^�	��������|����>'��_T+�Ua��L���i *=�Y��7'!�F����"yǌKl��������-w�Y}���Zy+����3�v�@h�f\x]2wޤ�;��R盾3����7���#ާ������%g,GD�j$��.�KG�K�*���J����q+�("sLy��e�a2�ce��ʂ=�М�zZ�{�Vq�{�^�h�A|PU���j\r���m���uS���iՉ�N���p��=����ڸ{fY(���'��p��r'mU���V�/��1b�>Xיݕ��0��H�5=w��Z�i������//���]��ix�������v�p�.)�sb�r0s�tBR���I���<�;��^�e��j�˫]�lu�M���o	�ᙎ��x�6p"��]��Q.�yu7��)v���;�E��>��u��K�$�xo�e4y���������Y��Z��Y<�O�YG ������)֓pO3���\n1>���o���_�����Ѥ�r.J�|�oTK�������L�~����.��`�� ] Pҭ����ơq��ƣo���#ӊ%fJ���o.+�����M�ӓ�\&�@�u^f��2JRWM��"bS�%i����6�����c�|{wu}��>W�m�|K>�3�K�#X4��;6fc�t�(�4���~�Gu�tW{��M-�����C���1m'fM�'.�B5��d����Z���&�ձ8jhrW�ˣ�<�wW���^�e!��w���wt/�'AL��ܰ�_`���*`�om�8�_�ھɝ�����cf9؜�S��uҴ���4nW���uO����3>sANJ5�����<{��FW���ߪG�K'(dfL-��>7�L�'qL��VǾ�UOI�����s�>ϫ�},����v�/�R�\�O��||�ςU�73̞>ɕ� �?��?).kJ{Gs+(+�Q"P�&��Į��)��]����/���tlK��~{���t��l{���7*�Ҷ[�*��S�K1V^��4$qd�۷�&��A�`�t���t�]C�֪�n��FV+lp�	E���6�΄mQ�7y*�5%1Y_re�#���+W��8�a�L�rp����3���G���umL�9�R{=�=����C�`+�0��_oW"��*H�u�o���Q��ʝ7e��
}����R���/<tI9��W�L�k�av�����ވ�\z
�������ItvS�mE;{�w^��M?�+_�)�����)o֗�B�in�z!薎z# �۴���P�O�z}t�7ς�]1�:X�K�d1ʃ�F\wS�?����ݼ<�js�����}Ѿ�~ip�ݲ��/�H�uL>�|J� �(		T
���;>������\�g+���ѕ-�g���n�"���Ӊ�þn���;�F��(�Ax��J�	�����t�f�z����uԩ��*c�)�F=_��,�x��m�N���١B�(�T�����kcCrg=�Ṿ�~�U�x�h:��9�e���Fr�c�r��>s8�^f���;t&�2��e|v�ȃ9�;����%Y'��Z٭RJ�_����4�����C"? �������Z��mU�m���V������mU�m��V����Um��m�ն��V����j�km��j�����Uk[o�֫Z�}�V������V���mU�m��Z�����ֶ��ګZ���Z���ͪ����j�km���
�2��x�2$v�������>�����>�<(����b	I
)R���k	%��BT%lb��6+"�kJ�i�m��e� �^�mKm�ͭ��
��U0Y�����t��,�Y���i�m�Z��k-Fڵ�kRA*��tz�;޶٬�FٱM����EU��%J��V͘�ͭP�l�5U��TY�a�ٚi�m�ٍ�M��Vǟ9�<M� �xx�`�VwjS;�t�{{vd�x��Z�{���m�Xz����v��oh5%��n�vۨ=�����j���� ���ַ���%l�U=�s^� ��� P �XO@zQ�����  Y{���� 7L(0��G������}E5�lٮ\��WN� �>����^=U4��]����=���:�u�m��S���d���t֛{=�z��{ƧOwn.�͵��nv��MZ�� ��м�']�{�����V�ͽ�4�9Ǜpj��w��ܼ��{oz����Uӽ��j�5�z�W�մ'Q���L���̦�m�8�l�w�;������h�q���嶯W���թ�=n��T;�wh�{��vz�Wn��\���\���^n��]i�q��xv�;�y����w����S�ʽkT���e�I���}}�`�}��[�t�y����j����궮���N�]��t�=�v޻e�*ݻ]��]�Z�׻���ob훮ݨ��N��^[����K> 6����{�s��oov�gM�W��f�7�n6ݲ������
��Ƿu�t���{k�#��M��^�z�&�v��@�[Tݬ�4mͽۚ�ѫ'\UCcw� w���{6�u뼽��{��-B��G����t�v�vǧ�w���֫M�kv�[�g�v��Tu�lжk��P�v5���ם���[*Q� �ﾴ���nv�ww]ۮ��u{̎��g;�u�[p�ݍk{�]:���/;��=�έ�z���[�^�����[fUfۙ�1Yi�{�ݾ�v��T����x��Z���{���3=��RǸ���w]�݀v��I��j�H������     ����RJ�� C@ � �)�)JQP40��b S�2�0d�d4��"��4�)H&�M4`#�CS�2��j� a  !�i�) 
HКd�h���MC�7�h�0�#e'�������G���ӹ�sT~��8+�hRY��+�����zL?S�?�"���"""���c�a��TM�-y�����������h��)4)��)&�w� ���&�@�`J@�PE8���.>��}��#��߿�~��t� �u���q���}&0l~Py�:~���'���M��4~�_������L�~w?Xأ�D*�	*����{I��%��;�b���[�(�h�cinP�(���2TU�3��v�h�Ȫƈ�R#sk7d�3+h��P��ڔ�2��e\�٩x�4��YYi�t����l���,�2`[�����������	��&jw�V#���St����yr�'+l�V�4B�����
�cè	ZmC-�Vd4T���/>d��̈́Hr� )�6g�k7*R�Z���+*E�29�#"�3�!fۦ�9��e�y���,��k�{�i۫5��n��7*�z���[G2�-�n]�6���ݸ�F��i�V��m�R)�1�f������� ��]�~-K�'Ea�HՔ�v���ي��(@޲��<w��L���L:&ڷf^֚\)aX-hXn�h����ŹƞLKv�r�*sJ� ����摵�J�q�l�����7z�z���7��7��/`��$�S6��2ٹW�ba���F$3e�hK�'v��������4���V�I��H�S3C�Zi
��;����$f���U/n�M�����K�Zk6'�������:�؛�dʀ=ۢ�2������4��ĝ1q�چ�༔���-ݦy�9��hH���;a�j�" qT�A�zћ@��*V����%+j\��.��T�Z���Vl��RT����h�$��xb�I,Ӕ� m:9-]7�U)V�".�5� �7�A���s��ʻ6̈��)暎Ik,7��K[�ɲu��,���{-�*�tzK[�.��AmQύk�k76[�5�Q�R�Ԕ!!j�7�9��[Z&�NL�ֺي�^ Jڼ�ҕ*���e�3���0�������&��]&F��]�Jޛ0B:����{zƔ�;b�Ie�r-a'����+N���y�1�!���,���ˁ��l@jZ��&�[J3���oPˣ���� �M�n\�u�mTxK:�V�h�9n�ȼ˨ �$4ȤH��NeZk�3J&-JܥQa9R�Mv�
9Zie�.$�S�����ۘ�֔��9j�I����b5�c^��ޙc-e@$7a-KUh�Z�J��q�˘I�ƻ���?�0�(e�Gwjűx���5h=B�T�V�,;�.� �4�Q%�fG�rj;cIV�s�Qq�c1�3@��`TY���%3N:�ZҬ�N�[n�4ֶ�Ek-������6�N���Ohl�2�E�׍�;�ܗt*��̌�%e,ջN� ^S�e�[5�%,�[z)V��^�f�k0��#�&��X���7A�\M#%X�F���Y¥����+$΢2Ի�A����-�%�#��nA�^���Ì5,2��mB85�V��W��I��0u�#cF�H⼑�k6���*7�T��kw�*Hk�f�����(�x�<�����4�&sQ��*@lỦ�����b��К�p3rU�+[��0 ̱���r�Xn:Ŕ&���0FT�ۣ��2�S�c	�!�� (i�FGAfa��7�*}n�F�Ǔ�Uۭ�̆�@���0����ӗRc6�{��u�)�}�QwJ��ӏ'��co!���;��x�ǲ�Y���1 ��3n��[u�c�8-eZ�ɣS�Fa���OL54� mc�a����y����h����N�-�A#8p�-�3`IY�ʎ% �ȋ�ϖ))o�o��T9G�;��M!r���qF�1���]�"5*e�h����� V�kD�n�E�X�T�ؕ�mJAGq���AnKL�)�Ycc�81�"�ۏB·�va�X�hC����i��`�3Z�)���a�8!ѻH�O�(0d�+4�^�mVҧE6Z4%;h]��XBmԽl���wYh����U�D;jb�um<�YH<��Y8��W���T!���%'��e�&�3kS3.j�D�1V�-�5�B�`��xhU�7[�
:Z�-nP9�B�iJ���T/����.kո��1��)Ò�w[�z�{��J�zbp�M�/jeU쩥�ap(�����m��ѵ{��&���೬�*rM�w�JNa��:�ʶ�-�=����.M����y���m17)i�8�E�Ӹ��V�Lb��V���݂4��M�f^nmbFQ�y���2h�n �I��-�C4�ώ^���{"rXn�ɀe"�"����l���JLk3 �uqB�m�űf[M�;T�ѹ�$��M�R��W42�8�۸�k��JxrY�/7r���gNn�m|��u�oa��8��W��̔��E�z���ʼ�@T���C!j���D8L��;KS�5tj�Z�Q�57��5/u\9J^�iL�^��
vlROP�ǁ��S�t*4�!�&K�S���"�lĵ%�\j�ځ��)��xFX��M���!�MT�0�QKcyH��w.�h2������9u��S��3.�E�ncj�bZnl��cz�r�ۙ#*�:�n:8Zå�Ʒ�.�V����X�R�֖/�ן
�n�XQ�k�1�̽;6��5]��q}��ܽ+E,ٺ�n�팎7N�Be�b� ����;�_�;ؘ��I�-R�P�+.�N��* �Q��M'Al�6���f&6�Q�mԋQV�m��`M��h�30a��4��^/�b�A b�� �j��.	�74I��w�bf,�7d���ͦԭ�p7��R��u���͌��հ˭sxK�����m��썑X��m��5hzз�e�v0�@��n����|u�ʻ76��=O"�31	X�s-(tf����;socI�A��F8ևQ,50��5��PIh=ޤ��������ޒ�L5ġI2��0夶�%D���*n�cP��Y�.�V�-�n�v� "�0CU5�ӭ��Z��� XU�C4���$f�]
�LYZ� ��ff8��wt����Z+45��Z$խ��T�7��	`,�N��V��݌pA6��I
�Af�ɿ:	݌�x�r��rk�� n�4YK3��Ie����qԦo6��Z��9����c�n)Sj��^:e.�6�˘\.5�Ɲڻ���2�b"�k�W��E��pjY���Xu����kM�"
�F� �wa������0;�q�Z#9��Ʉȱ�5'����pd����QÂC���ken�X�2���0!�q\�fMY�VfV�tY
Iu�C	 ���,)�ݩ�#~��j�4���)�X��d����En��;vi"%�2�4�4r�����*�|�<3l�d��k]���@�[Vr�
h�K��д�v�v.W��JN�bt�P�XXP�D�x-��j˗�5��v���9i���SġF�����dH7�[{l�07���0��A2���!t�V#d�Ty������,]:�bP���6N��P�J��\�f���6�֗��9�'�(Z
-������W����'��
��Ԅ��pv�7gi��lShq-��LwR��To>z�i4> �)=�3f�9<x-Y�U��ŕ1+�i��63EC�k�m��T�=�rh��;������p��"S6D��l�Uy���˃U�O\��"�bx���.���y�ϫ�m��q�Y�����;�ꆞ��ݽ0S �ť��(䎦�%<]!HT�N�;���d����nK�2�;Ш���0;�6M*R�V��$&KF���طAd�i:�X�yj
�nX���k�-Af��q�y-�2��S��Hڠ���E��fB�Z^���ص�h��֮$�{���ͮk*����`�(dڃ�O4�&��'t\��D���n^T�Ph���m=7WM�s~d��j5� 6��&b:�gN)H%�	%�}7# JgN�L�I��YBJ�h�VV�����^i66�I3���n��tr�Tf�-��5.D+&�o]l���-�Ѹ��R�tj�],��TnLY�Yוf��u�2�0n�Y�`47%�aT�v�e�7De�+^�*�G��I*�,P�.n�͍ջv3r�7`R���^ek`�	���0l�9G#Uf�śu+.1[���HZ����d��:��VV�D+E��[�o5�R���YN�� X��T�v�n f+YMi �J�.�n�n��KR=֖m%K�E��.��w"wbˆ��V�+wD�'0;�5�VNcO7vd3.�*�[���Yw@��j�6sc*4��1�xz�@u�����N^�!���x�ʔ�)�OE�t)+X�<j�>9�5�u�`�2�1@�4Ф��CE�P9���s�^�ͦ�JWt�˭�Q�,�[�]]S��Ïr�\�@F�廭:�5 xt�V��3Hj�,�ud3����Dų5Г��Bǔ[p-�$]L���T���Uy���.hѫm����I�����+1�+�Z�m2s:eMVmȝ��& �s�S)ń��:
h�����3FlSvI�p�q�x�4���3������z� �lYF3~�Z�so"���L�P$X�ઙR�"� ��*��޳��ռwaL�d̚�$��Z^bG:zPw���$Yq:��t ��u�����<���1іb{�5h�u�VQ1)6��l�ݣQҴ�c28��[]d��oA+���wA���(<�4�<�i���L1�;�s%�y
�r^_l8+2�(�s]���^�Ġ$C#���l�6���yV�{7e�J�X�6�A�ѡ-)Dl� �n�+hJGN`�t�@Jf��xT�\�6�T��z������������¿ld�p~&�E��8r�Ο�����_Q�}�f⾪��?Ϗ��?��                                                                                                                                                         �@  `                         f�Ix;H�Yzr�%�v������Ȱ����[ ��x�O�
��� ����v��H%ܬ����o*oy�Kv\�uSM�9ԝ+����/{hJ�D���n��{� �!��ʴ����u�y�hDrr�F<�ke1*��@��S���s&�p�=^�sZ��z���`�v�	��I���Lar9�y5��rmb��Egr0㢥]��S/:*�K������Q֗v�V��PN��J��4拘�cR�*����|�:R�y8F�$�ͱ��`��7����l�J�ha�������V�����i�ݶ��9+&7�s�;N�dYV�C�}�%�[�N��6�_Af>�U�v:��9)�F-q^ŤXt��~�J��k�聄(�1)W�y}�v���u���'�4�~��b��7�yJͤ��p�R�[�g+c�[�^�_6ݺ���/Fs���Bq�lfX��[Gv�c����
�Nd�2�lԴ�ܝ��-9���J���N��V��t�Ʊv!j��D�
*�{���Ē*�[-�"6����.C��9pTٵ��u9�e�]i}'9��)W��Cw�����7�#, c�'�vq4X���6�k�9+�щ��c�Lק��U��H��t�ʻb�#��3�gZ��馮'hf.��8�E!K���&+�;��a�e�j���Pmj��,��ue�C�U#���Z�;�s��Ҷ`�%��:�f�t,�p�}Gw�q[��ŝj�wfB�Gf�S��`tQV��&���T�^��2���ˮ�4�����x��g�98_�����8g1�.�f�=���3ɠ:DЋ[w�W2nf�S3�lE<�h-��u����+]ʷ������Y�z=�u�:��Y}6�3I*.��p����:;�P�sz��'��2�1l��`���Ml��y\�t���2��m��1�K6@j]��v��y.�rm��Ł���t�`E�I˯��%7�eT{x���r�e���y�V�p�H��s{��-V�m�m ���J�j��h�wt��v+J��J�G۲��q7L]�u�б��S);��#�7ƻn(f+���Sj�K�%۝W�p�٤����9�+C彸�QAv𔻱jw���P��c�}!}ԭ���*I��j<���**�ҦŮ��{|�z�ҥl�BvN����.� n��؄�͵XR;Y>/�b��e�\�[|B�!np�˚3;qa�5d�5He9��� jr��e�lc� ����$���5�s&��c���>D;��l+�q�H@tէt���M����*T�0Z�38(��r��
O��̵Yr���u+��8Y��$rv��%�v���+L�cr���+u7j�N��_w��r0m=
luح��s�ʘy:kU��k�� ���
t�3u`������,��/"ػ&M���Q}��L���r;�D���]r9+���{���KWʭAS0(���ʹ��/�\u�F.c��J�����p*���vT �cy�˻���4��l��� X��׭S�ҾT\68��y��ҙZ��-^�����KsB��P��:�O���'n�d���ZuIc���o��$p:�s�|�n˼a;�����n�
|t�g;���E����nԮ�ZTf9>�t�;�}2NhkLG,�_1-_)�����ecs䄺�z�R⹡�m��Khf�-�X@���X�K��p��Y>��������L��1���v"�}��7��%B�4�{�;8��N��e�&��{ssF�A+�s����CxA�����Lezzb�����O0�+3%��(x�R�䬗@��6��:�-�: ��b���H\��-�\"8�^Y��u;���	q�m���g�ɻ`���f���V�A�쌿;~��@�4bA��^��]�ܕ��KӶ(@e�Gwq�N�����a˵�P���S+5��#5��9�ԡZ�gd׮�R�ה�H�r�'� �c��P��:k_bc�;1�;B��^F�d]q�.?h�{�{9m��P�������%�
jL�I\�&�s-���jjⶺC��y&p�Yϲ�#3�4�������]�\XT�`_,&�޶��I+6�h�#�3�|�&f��t+�m�z�S�,���N��x��ULRQ�no"��Ե�Ϭ�tH��n���N�1�����&yx�ͥ�w��0�r��=$���"Eu�}$�R(E�ᵋ��/4�RP4���}���-n>߮嗝����m��'�!���u���l�滺+%�o�!g83KYƀ�=#�_:j�Y�0�U�l�/���9]@j�{�&�MC&;U�sR�t�"�v��Q�W:�t\Y����Eg0��n��"���ѱV���e�J�@ê�񿖙q�,f�p�{�.N�ji�nfn�iw&0>e�ar�eV����Վ3��w^@�I�J:aܮל�a�(qhG��uM� �W&Ӂ0+�v�wk�Qz����Y���c��P��U�{�4�x����U[�M��;;.�9ۡ�Z~y�;�o~κ��%��a���V+A������3�*;6�(���t����m]�q\�X��/u��@I�f_
�16���^:�*8MC����g
����h�k\�|�V�|/�*Z��n�܆>��9Dn�F�9L�VQ�j�Q��ّ��J'�ө�l��� C-Z�+/�H3DZe4hΦ�����s�g�]��9DK�f��I���^�g=���i�A65�P�Uw��Ӈ�-@L�70RMgrwCi�/�7;�}:��FdPq�F�N�w�{a5
}^):�At`o���c`��[�pf�!��Ux��Z���]E��YH^.�y,j�4Lvg@ōjD	Kz��d���4w�	��\~s�A��dD,ng�0�.�)�胹hs�qP3��;{r�l��t1�{q��+�\�i�X_Q�B�����q"�����VF*�����駜�c���e_!�ݷѪ�־<r�j+{�^3(�����;�cxdne	S�=�&�]�P)�mLN:⇉�S*t��1E�V������7�:�94����g��cs�ކ�=�z���r�;������:5�j߲����%LA;��j�pӬYr0�	�
�p�&,j�K�Wo
&��ħ��k�p(l�^V䖜Pwv�I�]R�j���)��뻜�|6�]�)���d�;{�vRl�2��/�h�+�H��^����@�1�NWӊLǘ0l?>�3:>��J� +�-͂)��nW+-=���e@�H� u%/�����EO�`v{U)qf��ͳ�F�p�/��i_ĕYx�m=߮�f��J�����x�)�:����PR;��tlu����m�j�X�[��f�J�wk�ލS����xS&\�p�'S�&��bقJ{����h�w��Cޫy�U���;]:��3���\%�.jKJ���b*��s�uj�V�L5�1WrwtL�,E�*Mv��r��.�)c �9���%0�8N���q�arr����@ha���=.kE�g_g�[��<Y|V�k8�r��EI�,��-�be�c��j^ujw�l&��\7�(cɅo9�#MH�-�L�[͉��!,��\U����\�{;�8��i���!	{v���?�tk'%D)�.n��g�fU�����3FMk�0��b��M7-�
��9R�t�BS��2%έ�BJ�w.�*��mJ��vγ#`�ף6�(��h �?����u4�KI�/U^�k��S(�d�wdΓ�:{"�E<Z��s2=�۩a!p�V��2�+J1�.�r��n�I��C��L��B���	��%c�����љ����Y�	Z��J���Y �^�^�7Y�Gĸ֋��Z9�>50�q�t����:����ÉX�iv+;EG�
��b�������AT��n�bm��CE
�v]�:d�L0�o�ۼ���}i%�l�N� �m��:���9P��b��<٦�tR�ct��]��O�*��+r�o�?e�E��]3#���Ϭ��ս��_:l@�zH�v��u�wN�����8�)<�-\��X�i����VBI�\�����p�qzTr�7X��eNxR��_���m��M�d���>�
�7��:��;��I�yR��.EI�tgz�X�q{I�/o��:��ۀ`)5���>�L3[��p,����Z�f��܍��Q����'�;d8Кf(�����:�7GOܕ	�/�y��U�q^f]$���7�����QMZfkgttrVs��*Kh�9*pi̸�ԭ��8���m��'��l۫��l��<Q�����	�4����%��ԟ��?=�k���&}��5��vL&�����jUc�<�;�LhW&U�Rr�	tW2�ns��I��&�[����N��1oZ�)X�J0*@Q}:������uQ��3�����r�0s�[���F1�k���s�y�Y��b�5���t�(a،{��#;zty�X]f�
��)p�}�f��5��b�*h���YJnJ����M�m7;6F����E̉�Ǝm[C.�-�,���ICHYg4�j�K���g����R5���vv�v�e!�×�9��O��V��D�ʾ)IE�Қ��$6܏�H�F���(Ǝ�FF�Ե�&ΎI#�;��O�hBï5f]ނ�M�9Q<�F����p��0� K9H�\a�A~�@    n� �            ���_3�����w���ѿ�v�@��)�R8�]�
�|��B����~�vU����E���_�7l�V�����'��Ō	��*����G�y9�s4�bMi���v-T�ٗ��˵i�|	�bfN8�}pVR�
���ս�ϣK7yu0��
���,����59m��e���3Em���X�T��T��� ��MR�-�e]+���=;}3$b:_V&n�ə/���4'0��h����rm+Y6`�*i���;;vn��C���ͣͽ1:q��ңm]l�XMv&aH������E����`c^�:�{Hu�}HGq�ChP�,9�&���EϺ�[�͡��u%*Ԩ��u�b�Xל1S\8u��]�ڱ���\+!���%R;gZ4��M�V<7�{L��&앒݀�#j��J��&䦞�Jͷ-o8[�j�P�����B���̐C�<�e����wi��t���7ie�5�xL6�m�����gXI��Ħ�C�8芌�9�vL؎m){m�صs��y���A�7��t���&63��
ʛ6h��5�U�ɧ�R���m9�����[���A���n�샼�ڥl�3y��6� ����7�u#�c�x�_�@Z����-sR��-�<
�͛-]O�;�	�_�]��X�Ć��49��b�p�-+m��k��E3*�1Υ�=��3�R����\w�LK��+C\9��E;uחv��Ż��uw9���SNy.��:q��e��c�(ڵ����ͨ��Sn�,��[�p����QC}e�u']"�tu�4$��]M$�ʖ����R�H [�{���i�n%�L@�N�,��j�H�ͺ_*�fpˤ��Ǫ93)���%1�3�鮩�]�D����N�(s��bl��g P�^����Vؐ�I&-=Ħ�H��g1��L�̣�#�=:�1V�kK��7�d<R�����4��2_ks1�`Vi`'�I�;���6+-[/�z��	�`�\�i�����v��Fݯ���$C�_R\�=�5Q@���
V&/���=)�6������b\ܡN��F�橊K�v,�<�:T֤�A�WNM�OC\�X�xM�cn�+�c�b��<{E�o\x�{nz�՜o�sV��l��ٸ�Q���x
�br�ͨ�ZǴ�GWP�α�zo��M��X��
�̬Y;����D]ZBd��^S���if�cL��1}t�L#\qT�1wya��g8�k*�*��V�#�����d�e��F�B�f"]��)%H�nK�@u��9���NV�ds���}٠�
0�n�Scl��ԑW%]��:�,�Cz��������[��p�)��KD�2e�Np=����Ld	5�H�2�9���\]��=a��}k�`V������Pn��mȝ��(m�o��n��晲mi|v.@�N�K�d�� �mw����e"n��JI��7x�c8gR���42��4��F0o��h��*�V�4d�s��˽���\;擥t���_X�YZ��3�I�o���>��	�7�m 9V�[�J:�O�%�]@��]+��p�t6��)��դ����7�^*�6f�y��	}Β�˶���V�vM�Wי�\}*!Z���V�N޺с�*����Z)�!��@jbV;��[��f�@��ۥ����ul�t���	{1���:���\�\Z�]u��o�$��T�
v�e�;|�����{:T�N� �v���.��<M��ƴ�ڜ�b���X����J� #�T��*8���[X�����˖ԀV�T���3"��x��ط8�%���.�Qٍ��ni�v�QٽĘÔ�s��Sj�DiG�摔Z7�BU� ��ƕ�wkqUA�[�6�r�3����1;˛r���r\R�B��ca+[Y��� ��_"����Nც�eH�k�-Ss����9���c��)��z鍫%�٤0Si9I�Ы�r��{k�ivk��n�mI �����[{�uȄ�Nl4{����I�%	�d��!u�ai�r#i���W2u��Q��#.Q�p�M�bg�A�(�0�-��eb�ty�p�tQ�̘�+iR����"��[@f�il�)�������W��/Շ�9FwBEP����-�δ๊lͻ2�u���u�n�!�6�8hڀ�� ��s�N��7��r3J�F�0��ަ����݅d��,N����f�$�_f����e	���RO���-º���* ���"��9(*��t��U���k��b�*,]��a�ɒ\��9���d}�z0!���62�>dHj=��,�w�mn��b��ݑՄ8�*��;i-܎��&l�IӘ���R���z���ygffc`��I���Kz]N��h�f�S��]�7X��RH��̑,��tl��� ��[EcG��JZ�t93m���yYt�K�XزЌ����K�KM3�d�Z}�{k�N��&NP��M�VtW>x���-�k�˼�!U�Ïp������]b��j��Z�o�Â\��i��G3�Ń,ʊ�VUI3E�H�}���$�7`��-�[�bDa��×e����w*�ET�`Iw0ݛbcۛo]J�br�Õ����x�kOJ��i�un
�ak�s,���-�Ƕ��m���&��t��dkh�p�8���r�]"�R�"
���FS�f�Xޮ3([!����̻;����yf���m���N�2��6I�ۗ 4B�Xc�ju������c�6��u�a���>.���{����1�Ky�B5XO\����A\��;d�8��EE�j�"ã,kB�v�[o(S�;�"�P!��f�{�����]8뙬�܋E�;Ť5�C���t�Ǐ%�vr+���$+Tsu|��b�9�͋���s�l��o-dh��owt:���mt���6\����W\�'1ꦔ�a�I�"pN3x�����i��$/S�Uyvm�t���h@`�L�m��K�𕣰����Di�H[�z�
�CZ�C�Q,����zJ͢��27�L�nl�}�㋪M.ݬ�N��ٯ^��z�D��#j�M������+���LT��}af�:�����f7��i��++e������e��D�ӫ�9�}}ծq��	�,v���+��˔�<�]�ۍ�d�%7��S���ڕ'U���աبԤ���Lr�qv�̥:3v�o5x�o�S��d$$��0"@^.��t���dP��%Z��m�9y.]5�����e��O%L�t��.�.�\QO����έ�@ra��o�:��^�V��.Q��n]֐�r�:����xV0Y�qo#��Ճ�vE��@��6oI�Qu9�@S{�pe��x�Lܦ�U�U����uNO,
ڌ�I0������є��4*��;tZV@�qV�kU/_�]�	$x�'��y��rP{rC�8][�s{6w,���gC��V�۫�.&�JP�<�9���ˬuz����O�oP�����Dc�/6]�aR�,٤�҃�Q5W��ͥ�QB�7|��y���&�Z�u���U��i]HH>l@�V ������kZ�j�
ز77+&���7eZ����WlǎF�����U�O4g��%��R,�����ᒖJ,���ʦ��3L�ɧ�eM�d�1V
N^$昈���n�d��9H�l��q��O2�l�.,����� K>G�VV�	
�p�z��g6�/O���g~��Jݕun��Q��Na�,e��q��e|v�]e����1-x@��bĲ�)����E��B	A�-U�;T��X�ɴ/BE��r#�.��N4�t�HU�\1][+�v��$#]C�wNE�Z�ڙt @!���(j8�ݜ�V�c�_���Qt���3�r>W������j*I��o�H2����u�1�d-oa⿴��(�.�ҫ޳�z�23i�qc����+hq&�--،��,F,�gS*��G�ȡن�\Um+�6�*x�9w�$�c�h��G	i.�=�M�;❑�+1=�T\b��� rmbL5Nuhy{�&��B������f�o#��+!46ҷCd�V�J�]�ܻd�DNIVXGs������9LΆ�6���N�t���͙f5;��ۂ�f��j��y-��Rwʥ��ԝ�'���3F8+ywW��Hz��ć)��lv��9N����\º���0"d���Wu�z�0K�`��F �H1�;o-�����C�݆io0H�x�'@�z�"�����`�"7{�D���뛡AM�+4�,J���OI�L��;� �e\�k�ޙKb��d�҃]�'Y��e��R��FQ�X�7����jJ
��&�h�͛�Ci�YN�E�΢^�����t�ܙ�Aiչ�]T�uf�j�WI]3�BRJ=*�3�Օ�*��2gh��U�����WN�ڲ�h�of�� b1��lTYa�L[��')i��W1w��ͳ�m��ֽf��� ���\�[4��ܹ1��s�K@����N.\�v&뻴�5�ʺ0�K�3\��X#5�$�w�,Z	��W��&�!2!{)A�i�2��Q�鱇K��:�h{N��J8�����k�j�2����!�o����
.�ͫ�x�g����*Q��5N©��O�]eѧ���͇`�H�6�.���3�:R�X�9/+J	s]�3j�C�ܡ��i�D73�{��]�k�v)1_!�*ZK�����Q��,��3��N��B8�˕'�L��X��=H��m;P=�*3�dK�+A��0ޛ��s���a�a�eZ
����h��	X��ne����ot�C%�˖����\w�|�u����DH"�����B$���Hv�"r|$(ї�o���`               fN���8!R���t�ٽ��S,����@X����M��s�}�2u��r5����w�EWm������ ��J+%♁�]?I���Kvcݳ�k�wB!����F1�s��Ze���%�3�s�Zw/�gs���R��|�gE�Rm��	�2���S¦e�U��)�9O���+�f��՚\&�2�bԖ]��,���BbBX�O�]�mI(�����}� )��|6��gU۩�h;vs,�ᐌV�����ۣ��]��N�%8f����LKl5`�lk�u����}rR<����:ɺ;i����suF#_�r�η�^;)�"��򎉽�*3�;U��,�rQ�}p̙�s�k͵�c'��j,�5xo(���M%C���q7���!�k���!��Y+��le� �	k��b�dqi��e=)�&��ؑi\gF��+hK�r��)0�.{V��
��dW
�#�@� I	#󙟟�Q�{�O#��)x���2��
2�
J�*���2���$���) �2�b@�lC$32�����j{�7�Ȣ�{�2()uaPe�%�S2I��TTQI�`jP�

�ʒ"� ȈJR��5��NNT��3Y��	KA\�DUPQT4D%�r3s,�R��u.�X���JhZZ�h�(ZX9�d�I�.MUM��i�5k1i7��T-.�!(J�$�,���&IMvE2d�CB��@`B��"	��>�MK�s3x��]�M�}��5�������`���oP��إx�sI��aغ������oF�o~������ib������t���X�`�U�s좟V��~�u.зϘ��Cjj���~�ɻ�`rcI�^�xk�$�qy�'G�\e&��|�*;�Q;�_��Fc����"�s������S,��-P�.�Vѭ�'�q�;��ܕ��v�b��\D�@[x�7w��� �{w���v�d���ظ�q�;���/�TM�(�ů\U~^m��N�����Hp9��Ӭ��jI��?{f�)��m���ky\Qcz�7��2Ns�ǎ��廫��'��yT����9�bѹ��u{Z�K����ɗ���Ek"�19��\�7z4��'�C�^�Z�o�������t�N�a�cŋ+�-޺�{]]��V���M�=p{�y0�1P���W�pgo>ւ6��s�2��=JV��K�&m\
��YԸ�i�YG��V�Q�q}I���7DX=y��u�P��)���窝���jÓ,�$7ӻ@+F͔{��O������db:�?v/RRou-���Z�ZBs>:�-�s�'���}�+���LZ޳4��yW�5'L��~^9�X׏��q(�Qv�uDXd�N����V��
��b��彯�(%�t�C�%iѥ��}���0ڿxZ�Q{�g{�9�1� 닾X͉J^������վl��G%C��x��':���u���z)���Uf��� ������V'��ʪ�w�3IM��tǦi(@og�3��S���|���B�	r�����BN�\}2tvjQ�cӁ�A����7�+hއ�Q-�f幘��b�xuƘ�����d��})�٬x�q݁ݦ���������KzsI��²�{���֫��.�F��h'm�'շ��ݷ��Ե�ftq������w���m���c��BJ��7�v��r��V�_c�3W�ʡ�#V�j\k�wg4ю���7����Y���,�9��-.�O�lܻ���{��ƫp�E7�뺍�꺩���������[��6\%�9�흝�X��ePJ.��P���;�R������7���c�"V����lW�k/wN��ʲ���<�IևdhU�yhi����k�|̪p)ڞs��+����^�i�-Wٺ��~��� ��+d�^Z%��c
��`���K�w;����~�lS̔�W`�,Xh�{E�Ցr���`��2�D5�Z�@�M�ۖl��}���@��kWC8���̋6bGj�z�HMW1���r�$.�e霅����성�<��</���Ӿ�S�[�-.'[��D�i�)=���4��X�C�v�D�BK�*��g#aޓ�{�s�;�7���8����ng�,W\�L�K8�#�fħ�ps��m�ˌ�~�r��`�Ƚ��>���;*#ؗ�0MT�ojkb�%����Jػ)���}ބ�����[�����ےR��y���x(*�&��yFj�}�}�{��f���U�}+&�("�_f��
�ɂ����S��U̸Bo�o)��u޻�h���+�w���	��q/����'�]{K�)��&qn���ߴfRR�4y5yb�[��R�3dce,�o����1B`�p㰜�ϑ�6Z6���2`�T����M=�NVYΧ3r�,�]��w���
�wڲ�4����{��3̑��V��M\bi���?c�u�[�x}i8w���h1ҕ���5�e��e��@orNs}�����[�<9ak�X�w��~�>�f�~��ݬ��t�t��r�y�'����E��Ю�i �{}F�:>�yw^{1�\0���-d�$č�z���������{S����|=�]q���œ��d���_<��>P�q[�2��A}�X��ϣa��t��o~�&;���Ƕ��J�xc�foIX=r3�3��%�^���N��GTt8����4��c[%����������F6��TQ?��b���j��KӞA\��oT;�<�~3'a����=;�s��3�ȹ�=ʙ�W?�X/h>v��n�Z���9˩E\QQѫݘ��d��Y}���ۿb��%Jy{_B^����{�z�d��"Fꜛ������fy��Tfo�c��	��旷rt���>�=�w3ذr�k_��*0{ˡ:�e<W��t��<����j`*xJ?{�g��x<�M�/{f.l�z��=��UŸp�vTi���rR��Uыc��J�0���*�?tT�/z�I�z*}�zp���{��&�*X�{%Z���ﲓ�͈��_��g6�1=Z線��vrjD���Ɲ����Ɲzd�|j���'�]t��5���tu7���X�o�w�7�p�&q9��J��Q^�Β����n����xv�i5o���V�f��R{X���fc��W�%i�Av�Ѳ�!����|�9WlDwf�:�ե��,��'��T�^dt(�\�����.ۉ�ӵ�%��{��F��Zة���Z������W��EZ���%hr��2\����u��6�'���n�l��{}դ2.Ox�Y%t;���펷�k��]�g=�p���L�LX�Z$'4��Y��|b[�Kn���������7�uWn�5N�v܊mz�8��W�O>wvv}/��`����vT7���m��o�o�׎�����v��c�|�uy��l�+Uȇިxx��ni����>̟U���q����=���	�`�<�2�CȦ��=w����k%=۽󜺁��m$/V=������U��_��������K��k9�=~��Ro^���IF������t���Yߜ�"ٝM�~F"���w��!�q���4Պb�Vu��<�a�d>����eZ��fbu��U�t��]�1%�Y�YY��8����-��l�wr���f�a}�gۛ�;d&b����/w��g���ww�fѤ�����������و{�^�r�l���]ٔ�y{v��wâ���F�y	Z{�x,�k0J6����ͩ�Z�;x��ٔ����b��[�/��,	[���c= ��s>=��N��7U�	�ъ������'}��q��V�#�uSm�%��.������'3}�An<��"���ɟB��j��u^F��Ӻ7��K7�%�^��>��[�_u�9��;�{ǌ��'���l\��Ag����&�E����;��<A���X�2�.<��z��Nȼ�s��+RC*�c�[�\t��-
���qN����$z����g8p�o���:�����%v�x���Ke�U6M{��{��q�+*Ñ�Ӆ������m�ʪbg��Y%�h>�fѢ�W�OZoq��eFd�nMnӺ�3��N���֎xڿ�Q��*���C��:�����Q�7��m\��q���Yq�������7� oa�h�|:�8.wf�Ԝ�5i��ж)��U�ٺ�����:���IgփC�yx�6ߣ_�<��c|s��K�gj:�c��qR�ݏ,�f9�������歿;Mg�u2A�9{?W|&������y
�|��G�V���T�tl����7�fkXo,~�V��_n��z#�u�O�S����C٫����&�*�)�(#� ��v�i�n�wK�
���l�����0��ݽpܚ����jvGNۨ��ok��9�CmK�]Wh�놙��,T�}�99�͎@���.,���'X�Τ���1����_��w\��64mҞt�R����ϙnKp�-tl��uF�;Q��2�b&�#�����͈ט��{�g���Cd��>u:�?�A8��+�gV�˝e�쫡���O��F޻X%��%舰%t
~o��1�����W�`��M�f����//T��M���N#�<&�T�d����+���9�3ܥ�����xg7�[��R��2��iʌٽ�Q�,G��q�w�NޙRa���V4���?.�UW��}�]B��D�@�o��N;Md�(Q>��rs���4���!�?�~��UN��y|�o�h��Q��� ]]H����� �4�;R�+���r��NX��[�w�pr��v+)�ã5�/4:z�bո�Jƹ#4�tF�%#�#����u�w�ι�6��n�%mmv\ә�HmX�ے�8�!}I���'3����Ʋ�v�X2*7�e3\�ە�weɥ<ν9��|��V��UŀV�vdWXk�oo*7{��Pr���=k����mN��5b�q��U�h΢h�튕g8��.B��-���j���]���ֲ�U�gƖ<�f5\yVn�H.�Q,�o��_Pںztv��4[�PF�ȷ!!3Wr�&�e�!���}�jc��]�C�X��J�g-ʱ�&��A���0�c7F�q�p�qN��c�{ox��Hi�r��+!�,��m���d&vb�!���b�C];�PY�d��B�Du�¬%X�_\�B�9u*=ooL��}'/�q�#�T��e��Pn5Wm�e����3��o'&1,�+���c���m�+�wSD(E΂t�&��gi�!�ދ�o.��b�_�}�|>�߀               �͍��A����mi����e
�e�6�+:�܍ ��v!�%��e]��؝�Fk��!jn�O�E1�����U��8CA	��Mo]MtK��fH�`S�m6�i�W�l/o��j�v�6gsM�/y�̽��#B�,�5�)ښ巩R�wR?0�[/��SWwAu�Z31r�멆��P��֋�47��(^�W(�۫��'�
���M�ɨj��on��ˋq�WXW�5���Ӕ�X��vH�b�7I�@��L�VŐh��g@�k�6�?L�k�Żi����b,gv�Z�+$gFnM��s�]�Tw楺X��_mi�g�&�2��T�oMU���AA��.,��
`K�������}����|��p֕9�N�ťx-&C�雴�Uq���[���D���cv`J��AMܜ5�ל*�J��'7���ε��ܟ8������n��]�D�� h �C��{��U-ĩIE)E�k���"(ZJ(J���(iW�MCk���2ZQ�i)��rF�(J

H�dd-.B�eITd&@����J�fb���4�C@S��B��R	{a�d	T�AHPQ�d�R�4��IT� 9@RR����̆E!H%B{JR���*P�J]fB[����_9�NY�YֈS�f��/�]��8�y\o&���V���ޣ73�%��8�$��D���|�ˌ䯦9+�Oja�)���/�p�m��usG�?|��?�[_��Y��j�s:Y�U.�O�ק3۲��a������b�~��֕eE���d~<M^�ØrN��Mǚ�C�V^��/o�-ޗ�=�d%a��o�����0���{������C"�1Fn���VD�#|�,��x��s��/��Nn{w�}{�d����c����*�rt:_x팕Q�^��aܹ�����~�����ʐt���c�.Ą� Y�~�R䆲S�i��]�Z��:d���Y��+5�ʾ�&U&������ř�u����}[<2�	��Q��ҭ9�a�=Zڀq�j	*���B�u5���e�RY�{�f���F �.*�P퍸�\�/&ws�݇B���R�;x�J/:��Z��&���RZ9�p+������r�ߺ�_��R�2/U��T��qN���Z��.�ڥ��f�	�N��>ԛk.*j���~���ғ���-y�7�뽅��N���t+�����#�_�����9����Z�#�ۃ������*6.-J�����ӯ����~�����Oyor�����n2Ԏ�s\��v���"��?�˫\���%����Ot{|����5{���o�߫�9T���?�k�#�{0.z�j�^�c��G��7��߫����O�<�r'���:�Yz�퍻��T�-���m����<���;�@8����򔵘���>��r�]�����~��q�H9�����S��^󽹕Y��M��,D����P���f���`��7ݱ�������&Ǭ�hƵ	��怫��ҫ�������i���Lv�1�/�싌�t����+ﾯ���{R\�k���f���E��2':�څT�=�5���1�'�nΕ�L�.���]J���>�D�b�Y�Ӻe�e��BN��z�0����R��'yrC�b�\k�q���9=Q����Vd����y߷G�5yS���;�=�0t�0@���]��"��{�S����,��ٝ��z��,6���SQi�fo��S=M\�TU���"���>�=m}��ETs2Ї��������A�o��߫Yy�Χ� ����>��m�=��=�n+@gZ�=��]���y�E<}͚i*������ڸ�ʔl�p)~���N�軆,�mO�^�Dv�/�tw��P+�L�ln�U��Lm�n���rUa�+��r�u/�[�[�0|����"Κ����)ĳ��n<�{�-VHD���ee��[J���\��}���%�,P7ם��ͮra�\�rP��Z�խ�\�]U�s|�ӈس�j�n�Y�S���r�z���sm:�����#�ewۅ{D��X�Y���->�7����q���^����2$T�����c�o��g쮙���}���7�=�m.FB�����v5��/����{��6��^����%5�=��&ϸ���d	���7�9��5���Ǟ�ϝ��Pq)����<�w���y��#!z������y��k��S6�ռ�R{)��r�&{����~���{�=�ߚ��}�Jq!��:Je�]�<Й2�y���|�~�����ii}��a��8��S[`myg��q�6=��s����{�����䧧�!A�p{���;��)�t'��9���2e��}+�w��-�|߭-/2����w�M����Y�k�0��=מu�|z)�m>@�2Ơx��������_# x��<C�>�A�̽�a}�߾48+�*�~�M5��D}�?����<>�:��}:�=�ѶNІ�b�r�[���{>��Q�F@���C�������~����}�r٘�w̃���tW]��{�@� f��xٙ������HغgK���	���tïP}w;��}'�J���Z^;��t���t�-m�#���5os�&@��\��J���}w�������<���P�P�d�q��솳%x��!:���R�K���A�ɿ8P�s�jWy��e�������<�ˏ|�<�l��^e�w�@C͹������]`;ǒ�p�}�<����=��)w8�{���ی�}��9�}ֵ�^�s޹��]���o�{zw+ܞ��2�q#�^h�_%�^6�K�/m�����pu�)�m!����G�J�m���Hs�q�^no���u�>{ϣ�>C��ww'�xysܛ�c�>��͊�s//�i{�������1��B��{��[��~��!�Z���Ճ��T}�D!��ܾ�ħr�&��ġ�X�2;qh�x���9�m#�&�bҜI���q�f��y����y�Cx<�h��+�>�����ҽۺ��^�v��{��09�;��l���w6�8�����y.�u��C��{�7�y�mϻ��}����L���{�%�
M��gcF�>����J�;����s�KܽA�'�=[�H��V�m�6�u�x�ν��6��z����t���2�ix��sX0�S���4�퐽�������8y+���� ���k�yW�zv~��5k�$�H}_`���Ԏq����w����w�.J��ɒ�.ư_%�XjG�y����U/�������ߟ������|�qz��;��qy�茑�1Jy=u�w��� y�o���]u�I��!K�K��s�s?������n6�v�||oo���U�*���G2�:r%n%��X�`v���,�7e���ܘ�����L�xP=#�X�qe�[:���tj��s�.�r�\�!�r�HZ���r���ۮ�o��Џ|�\�޼���h^ ���e5� Q����c�N�69�IA�AN�y�a�X��x;�K��[u�K��瑜���q�^s׋ľK�dr��c��!��������FI��D��N�9��_#$��4&C�;y���O{�M��s�[y�Ͼw�����˘^�}š�CFb{+��o���{#ܜu�o;Jo�I�8=��sK�~�8��}���^�g���%<_���}��ڳ����r�W��G{�
`#�pO$t�a�m#�;�jS���.�y'�����I���P̍���d#��y����w�q/2���;
m��-B����{!�`��ls�w#��	������\]�g�����u�z����3�.�naԽ��;��}��o1%�^��B��<Y h��}���^##�S�����M��}�לs�^wיМ@q)ܽFO�`=C�a��s��=���<��x6�K���B�!�84�s���<->��=���ǯ���~���T�߼j�
�������`�'��<���X��+ܝGr�q#�8��0��_ ��#����p��^~�ն���#f=?G�/�ຐ��^��x6��@��N��2C�0{��|��O%����p�	��T��#����1�����)��!~}}z��z����R���J�=����C�����/VI�Js�r�/�ps�y/�m�B����k'���l�\ieGP�;ն�7J��~�=�f=2��=5����3��vs��mf����3��%���9ߐ�K������.��ȋTO׳�/m��";G���K��[�.�$Q�D}b#�h�q�]w� sq���#��.����z���J�z��2�v3�_cm�0�o��� Py/�М��P�&ons�=o����<s�{z��}�9���Hy#��~i�y{�=�ͱL���`�y��:��{�tb'���:�W��vq��ah;����O�^}�}_�&��k�6�!�/�p{��m#����x���A���\�4��Ò�.@w'���Ǻ9�x�m��׼��}yǢ�.��s��`������ی}����8����6��'���Z�<�s���ްrrGs����v��x�Z�ms�=w����9/����K�nm��/QĜ��Е�&��>A�p%x#$M�:�Pw	��� q.y�}hכ��ߞ��=w�]�ө^����NH�-/��p����S�M�ռ/pq�)����9�x�F;��p�{��w�w�����m�^��q�Pq.��{��9�c��m"m��\��~t��\@lk6����;��O {��q�1U���UUq��3�����j�I��~�����̼��Ϻx��|����4&IԻ�e�;�K��0��q!���J�y����8�`{�}糮���ݮ��z��^��'w�AԞ�a���|���M��O�/���ļ��\k�_eߞ4��w�ąo>ǽ����]���w�~��H��mm���unq�ɯp�6��w9��{��߼C�}���0 9��8и>�xk�W�xTr/��?7�k�@Y�f�4��y��j{r�|�]��4�j]z�O_��~���c�wR��^�+S�������릆���R�GG5��ͱ=��~�Oۛ�L���΄G�@F��}��;�~�C�f���G2���A�r���K���'�wF�:��|�߿4w/��u&��S�5�]�{��ߟy��{�l��v��Z�=��6��1�@��awv�A����'P�/��̏r{'Gxy y&�Xy/�b;�Ou=�w[e�u��~;�o�6�ˉ~:�Kܯ6m��I�d�u��CFgr�A��by������u���b����{�������́o�u���r��s�~��%�Gc�u����߸	����'y��d���<��%#$�5+����A_1�Uf]-���=���m����ﹹ�e<����^��{�z̕�_x�CB�;u��:���Nd�;��}���O'�;ۓ5��6���Ϟs�j;�=3�}�����_. ����G�u!�Q�X�1����Hb���x�@G��K�$s�M����z0�/��Ogx<�=���_w�;�S�w��$;��8��2^c��������A���Z�ٛvs��q�=u�Ƽ\�������t� ���7�#����{d�����Ķ3�.�2rk8'��7����y���s��w�s���z�x}�yC�b�d/7P�=NKˬG�|�m�#�1���&�ħ�ܯ�m��/6����y�\���޳޼�Ө����N�����_6�$��}.FB�Z^��6u�ܼ��ة�o#ԛ��Jo����8ێ��E�;sm��q }�Q�NL���`���G�ӻ��+^�{,��7��M�bnX��&�zVsѱ��4�oA��F��z%vW8�s�����N)�ݺ1(�Ɵ����CyR�E�@�m��8�~��|���>:�8��8jS��|�P{/���!�_6�R�I�|ir �g�-/��k��#P=Jq����mw�y��^�|��|zm{�!�{)��!AǸ=��qK��^��C����2e�lW�{�-�|��KK̆�U��f���߷g{��琢��}�񯾫����!�m��.�yϸ>H�r��~��a�r=�S�R�B���~��7+�%���y���+�W�;\Hzf'r��0�@�7�B˼�uu��A��� q=G��ɿ�C�}�����Vw�{�q�>��ߨj]����s
m�H�B�!�c���'P:�%:��qx��}�~�G�~,�Z~��}��裼�I����v���d�U��Pˊ�E�'7DTb*���Ɲ�؞�^�3>���~ݕ]�Q�5�U+�^���.1��z�3&�7�탅�f��m�C
ܫ~��z�}I�s��e�Uoj;7�U������in�կ+�r���7���~N��)j��W���&��؂������\��Vm�-��{3R�3h]A�E�R��Gjݎ���\n�;?�E����Y��2[��x�l�H���童6����qe��y7�8��֫�'����Ԣ�*�@#H#B@-
4(R-(�%+Jд%%PR�$s��q�s�\��F�����/bw=��k:��%�Ļ��|�匷w�*z.g{f9��֗��E�BM=�;�s���+�Ra��}u���
鲭�_n��'6�Γ�EuD�w���&Ƴ��C��]}���2�e���z��@B�4��X_��I�5���0��t�:Wr�� ��Ucw�pd���5m?v�S��i��յ�C�~�kMu����l�MQ�J��7�t�5�9����76�J��[=�vl��/ڴs^u�p�xΗo{חV��䣓܏;\�^�n�1�ʻ֭&�Y�fefM[��Q�<<6sݒy�G�Ǌ�눝��s[Z�	x�,Z�V:�v�L�;>�Գ�t3;������O���sn�7�����r���ѼR+��b�q���qȸ��y#�� ���,޳���ȬKm«q̼�/z��n;��h���V��09��cq>/��cwP���LBy�j:7ջ-��5B���Ys;s��uň��30`Co*ﺘ\V�-���;�	��ĕ�Y�Oc���r����[���yo������W@�W%X�U�I����}}M8�VC6����$�Ф�*���];kz5��z:G8��yщ݀��b�/o)�K�:WX�^�xئ��"��nX=�DMJ�Z�]%,ێ8�0��:}j������_fwu/�V�ltˣ��
������1��������eX�5��`��ݶAѺ��N�����P�J(�g.��uz��AT� W7�1�@���P��]��YRpy�>8> e8�c���eN�(l^v8���n��]5�ÞTt���q&�K�Jz�m����f��DB�"v����~��:�U#��               ��=ݒ�6�Y��8��K1�]���e*�)I� ����f��n@w���sa��A�_QS8a�:��F5��r���
�Z�SW��>�A �v��x/��s�5����;�8�$p����c������=k�c�Z�]H2��_�A/D��{7��
1Yi�މ�quv�}��ܨ�v��zr�Q�+��Q[�=Q!�A)�7���\;b�I���6<C�M���U`��;��Kc��]v�7��m��U��]N�
r�1=�f�r��-�*<��7@*u����#(������1�$��Y�8n	������l%��ɑ��*x�-#)�m��*�f�xD��C�3_7;/I$�u0��5���7
V��<w��M��R�����u����lv�S�mn���lc��Q�xS��8�m��eǋ����ɘڧ��3^.�o=Ǳ:pu�Y��xP� to.��N���30�/I�̅pG��%�\����������ԅ�m:* (B��)Q������ԥP�B�o�NK�Ҟʹ4�JZ� )hkS@d�!HP�@�HRk&��a1�"*�y�7�P�#BP�͒E)AL�H�9-�Jd��H�%	TH�ILT�#͐RD-DJ�P�QCAqШ���=u�?Ey��\m*/�EM�a�0��N��.�wkS�' x���L�W�q8�=���">�#�s�q!��mP�5�w�UQ��~������~����u�l�Y������j�5?����z��U�{gg ��i�]��^��ΕT��Ϩy#5�����x��-�U�mO�/N֍�X�*!Z����'�������g�QF�efz�p.Wj���E�ҋ��X~�5��TD��ۏ"�٘���4>����^b6��R��;S�L92�Ϝ�Z�RJb{b���=���;����]��{<�}=�ށl�-����,,E���v�e�yK�b�bI9�2v��WO�V�c�g�f��3�h�Ǚޜ��	T��J�Jy��W�%�l=���).�]�	�9µ���s4\�ʰ��]�K�Y�35v�#}��:�W.a��d��=�m��f��k�^+q���;��K�
wT�۽�f$���)V>���L��ϼ����������Xk`n0_�q�ᓴ]W\ڸ�y>��(U�(�T�$��sa�z}ܹ�r���P�n�b�:�������ن�����B��aoC�����=/�at:��N�k5��z�k��������4S_ZopG�a���v�XO�@f�������ETs1{��j���c���aΪ}�*��|��9f�6=ӛ�5����96iz.��of��J�zW;�#�I��]��]�5���]'��s�s�S�c����4����Z�keX�/p��/��e���6mG)+ڎ�Dr���5)���[E��mv�U!p��_�[��g�0o�۷8��-�H��ʂN�s����b�p��d"��3&N��U���6��p ��O^�^��v��"��c/��V�V���!N9Ɋ������M��E@X��6�!�O�W��h�g�ﾪ����7��x�]��=����un�n�*�ڬ�'��vt{ٰL!h�J===p���:��+_ͦ� Î#~��I���@pBy���>�~Έ����f^��Ր���/�¦o��]]T�huu���S5K1-�mz#<W��,'j��I��#�y۫��6��w��6��J7��+��ᓴ[�sfW��k����@�S��c�ʯ��C=��O��+�L;��o*�)�^W��+*�0�ʎ	���VّI���$��|�޿�vd�p\��=o{��8���W5=*�w����V��l�.�Ϣ��J�{Y�G�J�Z���0��^ڜ��'�w����Ǟc	����x6�~
�r�p���?����{�x{&ރ+t��{o!��j�躈��vv%1=g
���������I*����gN��ag���e�ѩ,֏x������"��s�������x�j/x����U�'F�폨�p�q�F�nl�?U�����q��J���Gd����Гs����s���t�<�`�j��u��2��{O�1�3U�\w�I���c�r��Ⱥ�u���4��������آ���B�0������S�^��O/�ӧz��Ҽ�'�=*h.,���{��z�;y�Ū��޺�ؔ�߻�e���8�����ok3��յ���u�+�3�媤�6K�^���\�����첟af��L�%��әb;�9 ��v>a9�]��'I]R{��m:CGٷ��n-��t�4�����&kr�3I}�n)0�Iw�:!��M�t���.�����&�E��m��>��菡���͵s��wYS]��J�y��(�+T�va�'1�zO-{z���\!3�YJ�ݳŹu��j�9m�g�}��ٚ_���s1ƙ�U��?M�ep���غ�k9��n�~�Z负��2���W�>�$}���roo'��+9ܐ�k�����|��QK�>�W��dS{Q��sw�&��ռ���gHS����w�LMOy��9a|HJu'+/�=�����h��h��nξ�0tx���C9�����ͭ��2w��{:�V*�~���CP�9�v��j/7�|p�u��٫h*�}#�{��t��	���=E(޿�G0e��ZfmeMY]w�9�ވl5v�$�:Y"d�X}�3s�Go8�"�PdX��N����x��fJn��W��]�$�/j_���e��Qk�U}U�U7�$ߟ���C�M�{Q��bTu+WMY��_�8�YoϦ��s#��,����u���$����E��i�W��l��W�3U�T̠T��x{U9�q߇�}'�)���t����*����k��z�1j�9��4H��K�k�Kj�vS�j���WOt˙�|PΛ-â3���k���rњ�*2&�Sݓػ'�[W}B@����o�ׯ�$���0���亷���Hvl�ʘ��EY�k[��嘉���)����*ߢL����u��ޡ�f;hB�ǥ��<U��������9W������C��l~�Y4���7sl�`��d���X��!�.hed�M�ԞwC'N-&�:��,��`w�r�l}z�D*i͖*�� �'M�^Q��ފ�n���U�c�ŝ�r9�������&�c���e�j�ٮ�6zW;�"��BP[%�O��=�Ƹ��hTlޣ�r��F} ;�*��7�_�5����=�&%쮵e1��f��y/~�V�VJ�5}ԕr�Gt���Zny���8��A��O3S�r�9C^2��h��E����IX��8��\B�EW ����%b��w1矵��g��>��|��<���B��wʮ3E��S��:Z �Y����Ȳ¦o��V��ȥ�w�R��G������(H�����s���݅��%��3�G�L�I���ExtS��>��9�d�^ �_P*���	�0N���d��>�h0����[�����Ggb��y*fs��y�/׃�ٵ%҅U1�۽]�ru=�q���%���c��Wc�v�}��yK��\�ΑO��W�|�v�7Wsȍ����{u�.�5���כ{8�`�<�ý/�JW��j��Y�bo���Ŝ(4������-�z��70���9���5�OA�K����>���"�Q���[>��R��ȷ+�$���H^��]/9�r\���2)�Ç��֗oHs�g��q�Fm��Sя��L6ol}>�3z8g%B�&f����u>76�wP���xnD�O��Ҵ���a8u�e�,w�VR���WVj��A�v^X��p�����6������{:�hgWs&_ϟ�K'9�ه۳��c[���m{v�
����룩~��X���S�[�|�[G����5�:ҭ��}z�zMp�4���8S��o3��AǛbұ����{�ZX�����I[��������JG�q8���K��}�}Dr��&%������q�va��ICyk�F��vh$�m�5v&nϓ�#�9g*�p��:�Y-��c��/e/`������-P��y8d��Ou�Ev�k��n:0�MW��k�2q�K�g��I�m��~֕k��(D߹zj9QvR7}�����Q�KY����ֽXsk0�et\������������3�;f6<ގͯ����}�v���4�5_	��u����:�֪�oh�.�d����!��sy��9y5���ЎU�ޡ��mB��*]�/�L�W��m}\;�z�j����&%K���:F����T�L�S`��ףw��]�;M�n]*�'鹊R�1V���Y�����R��/�k��y]L�U�;ԙ�7�r�A+�E�#'��~�">��Ә����D��L���	{/���^�M��S����a�9�%�o��k���<�����v[�X�+7\s*/�Y�����pt��J��2�&~j�s�)�߮�#M��t��M�s�w:��On�׋�&D�ב��w��Ԯ�|�X��g'~��� ���Gک�,��6~ߌ��N�.Ir�޾Y��Q� � ��*�=���1<�R��5讳5I��wVN��(偕ə�ta��u�Rd;q����ĘL�����p�]uM,�yQ궻3�e*����=yC.�����`W<�w)���������?~ڹ{W����$��� �wK�]��G;k��*W�Vm��s2l ��{��p���7�bwHఆ��k���C��]4�K5�LR�]} ى��C,��r#4��ڞ�*����-.5I�	Sg;��A�"�3�x�Zx^1�h�q(.��&ei����;lnr]	`n&hJ���Ž��%cï24z:�Ob ��T�:��P��`�z��er��9��Z9���΢7��C��J(��n�L�
iuedT�>�r���[-#y�*҃�{��n22��	�� e��s�
�_n��EÑ�U0&��G4�*��W:k6!���m�(6���v#�y=v:�=s/R[�k�9ww����Z�2!�~QH�Lڊ2iFi�f�d%e_v\�Iv�Q��e�5_�	�ZY�\|zeq�+���0)V2U���!�;�x�O6�t����Sii�xӡ�2;2,�N+)#'��w<+���-us����u-᫊�j_6p\����i}YSq��tw+��Gƅx-Ͼ���)�^�-�=v�睆h�              $�k�$�;s�����G.R}Sv俒L�����Vt���8�pk���iK��s'Pj�&��!!��j�;z9ty;��p�w����K�R�6�N0�!��#��o��6�9H�mNsv:NM���I�!]�݉m��[��N��<6KT��
��-l�\9U��BQ�ZD�����H��':-�r�Z�t4��|N����˽2=4,��3j��zw99ZL��1���f8@!�9�֙�Z���yᬛj�����r�DB�5���"�.�o52>�r��G#������d=�M�B.t�A��eZ��5�J|�8o��;8���#ngE�x����v9�W�GG!���@�����k�R�;��,�hTS*M7�쭁�}�lJ:�e��q#&%;rj�jݭ�Q��
��ܣsa��P}>���e�;�/��T�E�a�:h��t��N��9��ʁ;�"C�7e��c�SpE � �7�����|�"#����0��D�0J�^�LDs�탱R;T���.��A��fP�+f6`dPX`�B�9'����(�j��L�0���0��r�y�k�� r�]BR�&�jʌ���V��2r�G`��B�f%e��X��J@,�������>#�K����p>Ow��3�k��
��2[p�yɵI�mъ�*ö�'�c��g�-�����#�^k��W�����)��G'4�o {��y8z��h�圽��{��?z������^���S֛�۞g��=�Óe����OU��'/�sѭEB)��Uy������`��7�2����꺠t/�!Z;�NZQ۝:Jqi�Xngr�7�o&�$;މ\�G]�3/r�T.��z���'I�hTl��9R���vίx����|�\��	���U��o),���^Ν^*[��ߎύ����f�헾'5e�t�9�w�)u �]�Ɵ���ೳ�,�Ƞ��:��9�o�mM������W�ʯ$����.�/�X;K9"�*�Ki!h�գH���ǀ=�Z��{�))1�.٢����뙀��u�v%�s�q�<9P��g�XQ��B��g ����%G��h瑋;�]�q�����������:��?�G�+ �Ypݾ���љz�׷����[[Q>p�T������E�U^�de�r9��&j��Q�]_{�v��;�c��H�cq�|=P[�e��TS���6}�sp�ն��>Hޥ=$���y�!�M;cJ�W��7��#Y)x��総cӱTyKU�{&Ҵ���S�;��/Za��ꚋ���&���d�w���ǳ˽1&��C��@�/�V!��fP�*���G�轙�)�p�gs�%��3̷��۲�iv�z6��4�߇􏌊nj�)Ǽ�_�ɛ5��Sݕ��\�
���Q�\��Da���u�5\&��.Sh�x�Ԧ{jf�I�M�g���H�a�v���jȹ��V�G�ewd�/,9K��ͽ��=�"5�X��܉I�諭�?s^~��������^��
�-܉��x�=��m�kF��j{����9[�~j��W��"=מ��������^ǧ���pQ�F�MVOi(��K����O<oR���wձ�eh�Hu7~�����������=�~V���[�i0�(��?�Ʒ�,����)�T]�ڟ*~+��43x������#>�u�^�u�x"�Џ_�6.���/u�����it���ی�I5���Py%�
���'�	���'j�����U]��k:�_�����˞|��dBxܧ�X���^P<�߫�b���ٻ����UZR����;��z�c�X��Vi+�k8�J��|�]���Ls���;Ս	Y%�W2�ڈ�ի�3r��!�����(+ϻ&-)>�~��ꮵ%�W��=��g'4[g�޸�ܬ��t�B))׷���6�����[*�5��I�سx��/�p���:ɗ�I�{R�9�9ykyhC�і��������s�{R�֤�ˬM��<�w����b�5�L����%To�=ǟm�)���V�GG��u��p���PoZ�$�;�V�L�]�Zt����%�\��[�_�k�G/i8J|�8Ϳff����\]��%N%qq��5\E#�7�\�'oٸ�ռ�=�$n����t�z����i��<�(�6����GvP�&Z5��䮥B�UC؁8)y,7����N����N%D�]���Q&���.��1���ͪ��.���O[#s���{�:>X�y»W���q.T��x�؈�2[-d�׆H���@�ٲݞq}�@��=5����S�}���y7���X��PS��*��&�@�3;��	�G�0� {�4��	Q���s��)\�����U�
�z�T�3�Z>&
�˃FRMxx��I׹��J�R�#K9m0�t�D^�hw��^�/�������[�3��Yj�:��
�.兘�<GM��P�6E�O���j��-뭞�Ӳ�&�jA
����,�0H(o(�5�B�]h.���֑\=]>L��X�p&P�5���Pq"+��A��<�Թ��G�4�>����O��U�����Mp��N'���\��TX�Nz�ݜ��ő��:�긆t�o���e��q
����f�sg�n��2�8
�J�/�����P�☻�r�ܬ��v��U	�AWή�?rJ��,��'������P���/�9�����ԋ(VR�!lV�� ����x���0�A��ȫJ�+'5��
iv+�y��䍙X��wbW%�s��
wr1hU��s�O��1��C ��fr5�)�T�
<�zl�J7R��#�z���d���U�]��\=eِ����4�કʺ��፰��X��72���F�ABF��b4���E�ڬv�h�^^/M�jk��{�g�ޥK#��a������ۃٶ�hY�X"'Ǣ쇜~��ܾ]�ܻ#�	�:�-�U-kR��D�c:��x���o���6>��R�����D����5����i�=�Y�Q+ٱv)���x��������j������,3a�h���F����=���f��Q�yhT���"�o]�	-72��rx��ݬ��ۭ�G��E�u�����z,�X�D�Ag�0ke3�;)o�U��&�����xe�g��0M�����Eb�~�V�)OnA�5�fl���L�8}�ЮkOnm���ц�k<�J��� ��M���������[\����Go*i�P]S&>�Z��C_�uԯwMv0�x�''k�.�3Z��pM}�)в�jd3W2K���]��7Ӌ��Z6�
n�A^�׶V��(�����SZr�<!�G���dg�{L��js߳�]Lw�g�\zآ#�&$��Ȯـ�r��3������w�:��d��QW�~�R��I�dz�*�f\���Z_z&7����'(]Jdb���[y����bF���̈́���J�|π�tH�=����;A�����7ݮo["$0�Z�ƙ-q��\���$:�R͈#�:fhk��n9��v�h<��Xl  ���Ba��\S�n5�1���f��s�̵�V��zP�CZ���uR"�#��������2�/c}9�Z�j������Sqߝ��F" W�f��Ź9�:Q�����v��/uS#HfeR�b�SE�Wk/�Ȉ*U}�G��-T1i�q��5L����wS��R�sl���6V�g�1�m*�(��(���.�T��X�ڵ�:���7�(�	��FX�3l�ӝ[����ŬB��Wk�����}2FN���W��Y�?G�DKW���g��IU���<�R&�(1�M4���x�}w �>)@kO���� +(ziW�&2?��qyA��˳�
��ݻ@�w��^mx���T$���<��K�
Ы�p�#�/a�����-����S�,��s�,X3�t���xK�+M�eC�`N��\���"v]��Tz�PƬÆ��%x�pxxh�u��a�����/9��$6-0��f�!Ƕ]���}��Ō-�X��P�+NzG�,XC��e��
�PU�ˈBM��z�^ʐ���xb��w���˨mXb�A��@�<X�g�k2���_9�dGs�s�$ƕ?z�W[�0T��:-�������t�uD�E~��y0�Ø�y��#�z�Z}�o��w��Mʁѣ�Q<+�"��O}H˾��t��r��3xVkmu�y׺�wQ�䗼f�/y�<AkQ��Y���o�J�Ex)��Ps冭,�ŕ��զ,�Ż���w�;��m���nȥ������+�Ie��癗K�_\7�g��9�s�Z�'�,�6�D����9[�<��zZ�E�R�<;D�|6���� ���r�a~>�}�5Μ׫���j���P_V�;>C��`�v]R:E�G��&���C��f���c����iK��P�����(�X��i�y��^�)����zH���S��*��i�C1p�K�r,���4�(K�{����LJR��^��HT���}�}e�3O��Fծ��Yt�����Ɵ���-�Ez�C�D�=Ǹ�TΨ���=(��v�f��,L�Z`�-d@�k��K���b��;j������2#k��qxD+҃��^��/ C5�K�ȢDot�2>�^��t\��W��"#l�l�=�F�x�]a��8���B���2�YD�\ј� boY�.�:��\��\��1�`�ᖺ��HF7W[�yVDwR��o&�]w���JwhNd��%wWv�B1u��Ö��b��f��tgjvk9v�O�n~��S�;��͌�^S<�OZg}��RP��k�zh_�Ι��:Cx^�R�b{D��w;���E��X�w��5�Eˀ�?���.�Ѩ>�d|�*�n����ņz،���8�q~��z{+/��P�m�	��çfv�!,�"
�B��ү�k\���uÎS70*x��p&�^��;o8ُ���n�ƇG�[HTit��]�����曮���w�=��o_{{ٲ����BD���w��tz�]�iV�WG��(>!^X�D�1=�����/x�W�+������mmq�&f�3,eql']�_�tZb��9Sb�]c�;��;��qim�q.�����TJ�3�9����l�oо�T:0���V�	��AV ��`�_:*�a�fz/9ƣ/A��dC8��|*XK�P#�:���xi�	c�R�z�v�ے�X!��� ɩhyS}3���J�dr��8�2N�M�E�Œ����8��<�ƶ��2GB_b^F�h�H���d�2�&�g�/RU�T�
�l��R�պW��X��we����B5�0�mhㆸʎB�V�ek�B|�
g
�v�|]���i�yALw��r�Ӧ��o �v�=�<��[v�.MgV��H�m��G����4���b�\�m�B�`��N�C<��n�����>��]�x:l�{FK;f�ً��/�fG�۳���u�R�ge{[��V^I6�;ڏ����y ��?���Y���(�����(V� kzj���Ĩ���(f�r�O���z��\�
��"W�(�6�vbc�^�.�޸b���{�B�knVQ䚈.��{��L2��f�r��K:պ��]#�;j��@�`�ݒV�S��(�i�W���x��K"���{�=�����t�3��TV��_�í̏m��qB6Ҕ�Ć�8�sg�$��y�W���$�c!yB����a�,`�              ;��L�6�
�:NIVɼ�z',ӫW��vk����}xv\�/��m=c��J�vq��g<�)���mԥ�����a�҃yK`\�Ģ���5��p�]��RZ�d⺕l0\3��N�8jgi�慽QÅ3`F'	K[�[?Sn�w���V"��91���r+�t8_3YU1��*V�rR��J��A���9,��PC�d�d4�d�Ɂ㣇]n�m:l��Yx�̭�lp�;8Mۤ�VE��l�H4Or�u�b'XҒˬ�js�� �sl鍶�lܬ|��*���N���P��,@{-�Ti렺m���\PO6jW��*��mJ,�_�E`tZ*红�QhX��B�K�N�\�(��T��ok*��:�=���7�׳�7���f �R�a�Z݅i̩y|�+u�ǘ�=4��$�4�Uha����V���Kev�L�K�Y�vb��r�ܯY]Y�|�cݎ�dՈ�ْ0 9 �Aq_�=?D\�鏢eh�C��2S�4@m�jr\��WR�ё����uJm-�i2���C,%)h�Z�Py*e�Z
�(\����(hA��P��#��R�5K�`�E9�o�i��ʊSQ��&E)���d��.�� �2�2$��lB��"�J�IY���_��<3$��^w۝lI�Z5k���-̖�c��C�~JyINl��_P铼�1SO���˪#.���Zю�JD3�L޺1A���$�ӆ��ǹ��ӭ6&�# 
3����]q��X��!c$�����ٺ�U<��}�O����e�/�� @8ҾU�ҋ�C��Ų�s�E��������+VD�ˌ��Onm��Y���G��
�4t[[�7A���魩渹��.K7�Z7��&�9Z{�Hvj���V�g�l~)�^f�C�A�o�3Wե�T���Cs��ɉ���
����)y���ݷ84��O��0o1/��o]�ا����t�Ų����=�^����D�=0_T$�.-���C{z櫖��i,��u�N�2�W��TMhTM���"a���rÿ��H���o�L����{�:�~~����\k��O�,�4]��uY�&����3���+��d[�Ea�YOҲ�?�o�����[�6����ffd@���WMR�8��1;�����K`���b�w+��\�u�e�;6Gf�.h;�����%����ݻ����~��r\f�Hj�+8�$gF���e�`�[-KgsU�����\e:�F({���{m���fL�9����wH��D�	��R[�{1�i�
��Bf��-�*dV�	�~��,��[D�E�՗��Uf�lb�I��r>���t��e3�x�t6�S6"�"��[�����w��L�2I�Ȏ�AI��B&U����ơ��'Q�*�Đ��B)K��f��,��]u1�xJ�����&]���CxA��)1s����$hz�(tޱP�a�G�ʱ{�������N�zT"���&���Ψq�T�*J��w]]3��}`R�\��{��p��'�{Ve�·`s�y�R���\(u���΍�^?\3�(|t�ڼa�}��Q�����hOyL6MO%\���t�/���c13�_uC5hkb��"�q�:]���ʌtΡ����+N�ǜW0R�>>�0>�ى^g.&Z�(NC8�Dmh�G4bY���o|�:��;�;bѕ��\���+n@(Ě98g��Ev@Zێ��RG/��<m7���a��,����ty`8i��ß�	��)-q��t�L�]�`7��y��[��yV���u"�gV��T���:�-�5z�]C�=���o��ϝ9�',��e����g��R�*�:|�Ыu�|�F��AΙ�L�t<`�qc������ܨ2��T�]|�]ɳ�qV�*\Kܡ��a���2��q�l{W�%��*�!�E�}���y�Ь:H!�ຐ�+qb]�yl4�Ac���a���'�D��4�bY#0� A!4 �|�U΍o�2i�#�29ν��>���������o'ν֍����\�:�/��@rkI��9�S�#���O7y�2��u(v��)�ΕDI4���4�&�-*��G���Ys�y�<�$v!�Ԩ��S/:�;n��l<&�q].�.aP�{A@n�g�����9;e$���*9������+P�v�'M����$|m�< "�b��{���*�n�lҥ�5��3i���	�Ѯ*�u/�7iU�9��w#��|���'�L~�vND?�tK��a��ur	�e2���W��s7۶9�)i��p�2�D	��P�1Gh���7��o]����D�
B��!���ق��S�c<,yx��J@�|��K�{���Z�)��,V�i#Ώ٤C�Ȱ���G�=^/"�]�f�f�{�EA+�P�*yH�Uzm�a�|.���ʧx�c�ê�u��)���Z]�.Ϲ�nv�{V?*��t����FT+'T�!2���G�:`DA�_�����3�u6:P�nu�Or\:����BF����ңrd����Ba0Ī��垾0�s�S6&���YN��"���d��K8x�#e.�i
�.����-��)��i��Lm��I5����zmu#�
�"�K��T^�T;-o������2�U�Z2�S�Z�cV��J�ĥ��Ҏ� ��k��<OvDRYI�c�]��h�;mW.	Ȃ��+���ܙW�%�t���m�7�>�m�����z4��z�;v���(���B'o/)��u��-��^��4�wdZ0���[4`�ۃ�X�ϕ�K
��ڼ����|~��c7�eo넮���?��0ԡN�Be*��'����>��c6{���&��gx��������� (�nʫrp�?4�6��:���O3L�>X��"�z�5L�aQv�=|�O���4�d缞L�i4U�C�ѣ�M�ޡ�U�D�\h՘D8���3�ߦ���7�2��R.����tJ��u~/Ư�ȓ�h�qe�ͫʻ�b8�1��^-(�-V]�̖}���&�W��e�= U`�~)IxBE� W��rx�|�le-��yB�j�+��ɗ�K�q9*{�zvZÅ����Ǎ������58�w����f��I�GE�q���v�=�w��'�U����:����Cy�=����=�5r��V���[OGw1Mۍ�Έf��&j�X�϶P�4P)[n��V;�ǲ�RJ���r���si,��0e�g(5���\���\���ʎ��ׁ��#�/3F:�~W��d�a/�T�U��-}�v%��SP�BϮ\r�^I�U6G)�!�Lz�"<�`a�:<��8� v`����C�n�h���ގ��($4<�DȠ��A,K������Ԡ�Q�|�xVg��Y���v��c}�ή�8im��n�Q� D�a8��+D�k����m�We�ś/���36���} �y��C[��j#\l�_������g|�.�����3$���E1hR��ڄW{m��ɗ�0:�I=K2�{�a�my?[�@p�(�������k�pU�5��9�A����u���|��ۿ��Cy(�P���>c!�d����5��hI���R��-�?oM�7Ά��e��t�Y�+���gl+>=yG�P�ZY���w�Gn�@j�:�@W�{��IWI����>�הR\Y�xyc�J�'�;�hK�f�Glw��Dզ�c���*\��]�̳���1V�
��X��Z�bs2�L��u��Qm\�4!,���>|�7PY��v��睚�����{�}�vn�)+���d�](x/Q��"'YT�,ּ��mr��'�sw���5kUڿ�*��hy��Z�.�H~�X�;������K˸���X�	qɟu�*���E�PȄ��[ʅ����;��V2{��9uH�;ј:���C�^�h_��ȴ�,z�;䩎��i�mCv{=ܓX.1h�a�L�}mA�4�3��x��a��謹��7�_{C��S�榯d�7+�����e�Հ�(��i��e_p�z��Fnپ�U�����	���`��1
B�%�/M�pv�حE�G�G�Q+��L��cCŝ����^��wC�i�>c�׽7��xEϒ"�̧�1���k<<5�#�c��9��Z��˪bGH��7�i���区'p��I���R���Q�eŷ�e����ѻ��X�x^2�r�ܲPܛ��X7��՜�
��Q�K&T�![Y��}���:
ب�����j��b���	ϸ5 ���k{;g�U}�;�E�oe-2òG��(�ą}txR�
��g��/�t@��)
}��q�Gپ�-;P�ݕg�P��h�J�/t���TY�`�֕����O==,8H���^~Z�qp�Ε*�iM	�Z�z�߆�q��N�w�Ic�}�Ŝ��C∬�L�A�huD3|�T��2�j���&��������ފT�^^?�*'WCB�K�� @���3��I�V��FZ�4�04��k"�Ap�����Uq��;[�Y�eI��RG�P�6E���qzʁ��QO]s�R���U~�b���J]ի��̈́�uO����~
�Y}zD:<�[��4A34Vn잠�&`|�8BD��<��r�{֙�s�5O��	���������ɶ�z�
v�N��Pjf[�g܃�7[�[���г���b"�=|�׋|��F��d�3��wVMKǎT��u&�$]JD����jm�T�q�Hj��5f��D��f5��e���+7�9�'P����c��v�����í�;IL�ğs��T|��8�i��>�ג�#2�ٖCD,�ι��K�U�ܜ���.�J�TQ�ƸV/R�8x���(<չ�O��;���z^4���Iu��k�0�bfRDj]�2!�X{��S7�^�����k{^��@Vh���y#�qq#�h�v^
�؅�맫%�{jk��#����ݺ�S(T
κ4�#Շ���K����Iz��c��z�f/T��2/��y��������B��&�Q��Ø��Z��T&~Z�U��hxx`Ђ�����hyb�~���>��$X����^�
&���F�����i�演\�����2a�F�%�]�Z]e�u�qL���D�+��ŗ����#�<��7^�:�^؈󨀦�	��X��ȅ��I&�P�Zƽ}���Ԙ�h8����8b���K��	��j	�J���A��!p|.1��^�l�'�7�r^���w:�>	��\%��c�����NV:�/2�X�z�p��"v+��E�Й��B�N�n�':���	�'��N�Z6z���*zj����~�v�gͦǬH=�B�L�L�C�\�xt�7��#�X��Y�p�.+f���?)��>�tz�����߮6m�7�n��g�:�̟B�=VC5�<�#\p�U��1~�ڥ&7ǃ�*�V0f^/��������e�7�>&'¯媥�����x�J���;��ӭ��'{�E��AO��7�����>/e3|��Ų����oj�t��ѧ��Ƌf���Y5ƂX�Th-�/.X��q#��m���fwH��3�P�ng���\�>���4'	<�E��G�Ȃni)��?%p��~��+x�m�S�b�j��Gz����<�AV�')�o�s��J2X��Bԧ��3T#{�l���,t��|���8/��ߣ_E�~�}�U{�V�����k]�������B�p��%���.�r�O0�j�Y���S�(�h:��r�2:$�.�0jUepJ�b8��б�O
x&���7�B�u1U�����N*��x�]S��X�	��<�V���Gv��3А��Ԥ�@f��۾8�=afB2
U;��Y�6�eo^�s��A��Ed��Y��m6��'9�Y�`"a��͛��i�9<db�c0���ZnT�
�`	.�y`�!��&۫��pD��n>��Ǆ����������� ���B��ۼ��D8�� �n���}:�fD�]����O�wG��WF���C�C2d�[qǒb��J����vy��T�@koɇNv���G�V��ﰁ�~NJ�;�@�^c�4������VE$�f\���^]Ї.�V��ܺ�����X�f�R=��\���!��1�3��W���b�����K��h���T�ݐ:�4���&%+�GDs5b�㜨�h�֔���^�a����P޼-�jT��*?�SL@0               3v}���Y�e�����s_B���)��GƻI7���|L!�>�nq��=���q5n�&��6��jniܩN�scse��ko1c|��Ũ��ipV-�a\Jp�ͤ1�̓�d/�C�\'Bi�5���*+��e����D�z�ؾ���R��zI�Bss�Mn���u`�E�2��Jr��-��n��~�VQ3�O"j.��;��Ծ��S�p_�ܵm�9��� �j��J�P<ac|�է��/��%��Kx��[��p���R���]�N"\yk*=���n���%Y$�j�[b���\GQiaWNA��6y�Q������,b��8��6Kg��Z����)X�U��.'X2�	҃�j�f�O+,ڊ�MT/��f�^q}y;HGW9s�u�VGu3�H|v>�9�w�;��-�)�n�K��W�c'-��o��;��
�QW�b�K�sq����@�*����r�� #�� �C�Թ�C&�(<�D�5	��CA������j5-�Z�Ֆ�(
S3)���2�0��hi
ru�5d�eE�dO��Q�K�I�d1FaQ��MXX�FfPee�V��ؚ��̌���(2k'��QfU9&E6cY��ט��,0�,�
�,����L�����2l�̜̌� ��Ȍ���"b�(�r���p��0 ����,"/���{�:���:c�e��zr[�2co��(v��v�r�E[,�����#�� �f�o����<����R?�z���BփMj�#�Mg�p������ӗY��ɽ�yLs:=�/�#�]% b���B���i�ȓC��r�Tql{��Q�}a�,!��KZG��u���!��.�!���ss�I�Gŭ8}�	Vx�R�H�:���1�imY<ty]����-7�`����E9<>�� �P+*;�2H�yV,nR�;B���O�yES��z9݂�%�+�A��+�!>�qF��f'ΖH�!Ns����{w�ݝ�Y�K7=/�^��r��e�@FoTK�T3�J÷[�ɱ��2(4]F�ۭN�jq��4�W���h������U퉳�φ�����ł�٘�'�ByaX�����0�~�@Zk�Qy�<D���aO}��}��Q���:�U���B���S���O��~��u�!a�y��q@�$U�����G��c$O�!�bY��2��Ī����5L*Ddj�j#7Ǭ�u��5]��i��NأU�FW/�s+&wj��Fw���ZI��fq��߼Vm2(s��m9�,��� ���o�3d#nW/e���b�^V�J�e����k�	�b q'�L,�.'��o;��U����i
�Cr��+P�z����*G>p]{�e���z.h�%�7iI_|R�ŉv���B�iL�Ww��tR���>�=���RH���8@�<uQ�I�\����&��ř�[G��>tgnغ\�8ʳt��}��_B�a�T�:�@vP�~�#o=�rt��0�H��h�����uJ�Y&��!�\��'��_??t��6�f�yP�BZ��TE{�2�uu���vMP�B���s.���ݷ�6���8����� d��o��F��^M�'XaW���5�s���b��"ȁ>�AzTHEw�r=�pwM'3�Ifp��2�^Wt�@�a�ˇ���a���ȡx�t�rYq��x�9i'VtVz�[�Wүk�DY���S�ro8Գ�yR���pS�y)\��4�v��w�\~��Rg4��6:Y5�01Ly�j(@�ߍY�R,�,��]��4��g7��x��+�x��?���g�eQ�^x�O	�߻k��H��J�{$:�+������q{T�b���7�/�ő��6�Ռ��u�c�A�q��qL�X�=�;]�V+U��.���B�eֽcW^<8��y�<��~�3�,�J\T�"ݹ��}��S�3��g��ѯ�։FH(Qf%V��,��!��l�P�6���3j�G��b
�����A�!}�G�[_Fz��e��(�{w�X���i�Pw�Y��O�'�V�i/~�v^U ����g�n�I�[����[mw�1�ΣYQ"V������<���r�~m�E�\FN���23���C��ָ�@�4GT7p��%�v#�E��{(8��_>R=��8��:o	/�me�b�
��6�)��sӍv�{�Q��ܒZ����%Z9y��'���-7So9S8�.U�+FN�˭�XG��cz�:i8���d�oL�[�?(P�.�P�we@�ԏ��,]Z�&������};k��p��t�U�Lʻ�5_��V�-g�+U�2�lK���Yi?/{�c&*��a�AP�k��V�oP���B�.v߉�X�����mLI,i�6�:�؀��P&����Z=~W.͵yY+��Ԓ���ץB�|L=iV�E�x��G�[t��v�}��	�{7�Q��{*����⽴��.�+��Տ.��Y����jU:�Ʒ�6��m���#)3�ڲ�K<�#�'�C�����n}8x*��'Iΰ�%v�G��#��3ddLy�)Y�\o�����˸d�2v����H_Q<!L��p0��ܦ�ؙ���jɣ�o�Moܡ�\fr�WVpj'�a��/�.
�W�1��̫កl�fD��wn�WR�C_����uݖ"�\�Xn�\p���$�M�o&HJn��al�n���:��b2:�~ʻ����ot�z,Ҩmڥ�;U�Q5���Ч�^�����eG���چ
���q����\��3S��I�y>W�ws���5���oX�TwO>8�$ 8d�����K����r�'b�WZ�J���Fy2�+K7��F��i���9Kq�`��vs�,�K� ����B�`N��ڄW{m��r��{��V��8�ϔ�S��W��H�3�4��5��T�$VpU�x�4Ъ4���0�ڤ%��aVi>&U% b�j~�"͈7�>+k�YA��R�oP���gJ1�	��RIMt�N�*Ɂ
���v��y�D��5�"��a*�*P�ؕQ�R�2M-��SZeP�Uvi��93���2��D�T5�Fm�ȉ|���cE�أL�htޓ�zv<R��{l����X,��\Q���f'���.�[T���k��͡R�\���V
�.ylӾw,"_C���YfG=��w����6�,��{%B��V��sq#;�:�w@s��7�OW0���@����"�]@��=τ�}U�O瓗�,�x%��z[9ʋ��2+0���&�D��v�7��`�,�9^"FEڸ������0�p�xp�.?'��hd�0N>�Xƍ/N��MW��qQQp��T׆��o{�����.��gN�cbx���A-���Z-�����V/;�����X��F�u8�m29��6����,����_ˁ�}Ob>̧J.��9;)�mW(U��q.�T ��lZJ/�6�{s�;��$��ϖP�."XH�h
�c���+L�g��o%Cm{T��f54�{�};ס���#��R�r#Af$4���ԻT���}&f�Rfn�?y�k�Ce�Ń��]T�������ȾA�!�*���}N�Ǘ���h���<����a��ݕ흆� a.��t�������~ܢ͍[��xP��٢ݫ�t�EfPݐ����u�m�#-����)�i%�P=�ͱL����p=��Ҷ�X{C�9���ͭxL�g@������9����sp�] �}-���qϬ����~Z�5�
��]}�if����ዦ�{;f����ѣ�*�*�	()T�L�������L��q��N	�"6=���SV࿼~?8��� U��C�^�;@;��w��s��8X!�"Gj2�)�~Zn�n-(@s�jTt�������t��钄�I�p�>�!و	CBe�ѥ=u��K?Jk%��n�΢'p�Cv�+�^�%膕R��=�����8לZ/�;z�U������5Y���z�\_^���?(�o,�������U���g�氍Q�(���"�\]�.ϹE=�=S[�M���f���a:�"�1B�K`��|e�2͎�0۝p���ka�Iy�q��-]}�Ps�։F6+�a(l0�u৵��\�`B��,-���m>��q�H�(7n��֪�eM1O�ޗ{���]���6a�>Ų;�*�A�%-ƟNK��k-��v��/;/7j�KKऔQ�ub'��U��E]�^�wZ�w�>܍���R�I7=��HbS�e�zȺ�ǆpz�Ϫ��(W��SΜ)��w7�8�#Pr)�tk��b �p��[���t�.�����|��6a��f�F���Vd4�
�WV�ȺF�0�<�y$��ۿI9VX�Ev�U�yA���g��^v;;/qC�@���w=��PR�O(P�.�P�we�S:a���@V��6��d�籾xt�l�k">����]gL.��xV:\m
�c6zgG5�Ϗm�f<4���_$�ˬ������j� Z�&pr��IU�}��ъ�KlK���:�
b�h�J�v�)rR鸽{:�$Пg�%8�ޕť����ge,O6���+rn	����?g�:lm������\>S���ryA�U{�5�I}���^��@sJ�C�f=q=7�وtC�c��������Z1D�gݘ�Q��x�n�Z�u>��R,~�D{�suu~o/5͂���l��v�'( �U�ڃl�v�58a-��o�q�Ls�ꮙ�I��B��a(h#�m���Q��^��9�ws�J�8 �*�����w��=6��?\\'�umKX/|�+��6�t۝�2�
�+=1ArJ��d�ߍ,5�x��?gI���n'����Zڇio�E�^[�5v� 6Zb��0uח��B�N��o}�Bp,!�8�N��}�3�� i,p#����w[���J�֤�C9sH���L��cH�![����=U���6�������"�Β�`�^P<��Wx�s������B5�i2�Z�����I�\��ĸ����CS����yB�m����G�B39�\y�ݮ^wk�3��ؑD��xsЪ:�~�tM<]�^�ߵ^�]�q���f,����7��2a)28�Ϙ�lU��	^���d���7�����P���%m\��)]�P%Ӿ����S�Mޒ��������B�w8�F$"i��\7��n��{�.��p�]�5&,���k����ꦬ�ԧ��d�_��=��H�L)�$�]#��N��;�][�e��`��V�yzR�^dx��|%W"�"�U%�MmV����c*97�$��geT5j�i���V:�YL��K�>�Fs*�����a���ɶqan$E\vȫC�5J�d.(�7KN%~����WY�IՈ�.�6=�,xߑ0��/�+���ʋ��2+0ꡖ���Κ~s!d��؇�8p��������D
ү�z�}�#]���7n�<��u�����6s$�ׇ|u��c����z9#��J�dx�����#��O%K�8�Wkk)���TܠL��=&�w�)��q�"Si�\�;Nz�|�{�4�Wd��nz��M�3�"Z2�(_SK9B��̷Cś덇��U $x�W����k���KL�Ob�Z���%�*M����g8^97
޶����1����"=q�s�u�[�+m�u&���w�����ɟ
ĞS�����
�MQ`rtӴb;�Zt�u�(�%�$u��}�˙{�'T��e�txt|��	책�T롵�M;;�����r�]����iΕ����'�c��}�C��@���/~�q�24�2�8�F�*N6�
���.����Yg_p�â59�޾X�&��r��u+L������eB1�m��3q�#���X�ٸ�JG�0�}�B8��1���Xk_�;X(i�2鲚C[�A�ї�B�z��+eF���
S9_��uA��5���%<,78:N����6��-�[�D��k�3ej��oGyP#�dI�cyX�M�W���uɞf���j�N�|z��z3�U�[�y�"��`��(�uFʼ:61����34_�|�ձ�9��1�QcnE2�n>{jw\�x��,�[����{՗��WlqPvb��             I$�A��_&nv���x�g����A��
8��t5�i:3TX<ْ�b�	�D����:��1��/oF'&��*V1��xZ�d��Y(�۬��D����p�`�.9SC����WJ����_^����
.�Z��=zyUXgr��:m�M�K!��]*9��n�Mh�7I��WWF�)����wo_>�:B�����Ӳ�F[q�wL<�l�l�1�΀�E���&�wt��e[�t'
��M�[2N����Ձ��?�k����UL�t�:h|Dy���[;z�6�f�\2��{��mB3�T�t�
�f�<k���d����:n�����Ɵj�yt��Q��`\�1W�-(�ՃR� hZŻPn�V�_;(�oRn��f�2��������i�ۍuӧq0�e�9�z�+9Q����Q�[a��6��~�^1hqF�ᇃ�[�]�Vftf��7���|�&2O[U�噛��:qO4	RGRI����(P |ɡZ	��Uf`��ޜ��9Kde�I�Y9$Gs�-fcFYe�a��dY�E�A%F�A�NYRQacUj֛2����$�Y�F��F�%���"�XeSDT6��;�5���1k(%��0�Y�J�,�Y��1�2*�m�(�efY�����LS�efY�OX`C�¢hʹ��u���eNѣX�4h�#���ֵAQQU:���D((\�6=Xb�*�R�h��E�����S��u����.�B��tx;#�/�_Ϻ�6�̩�z�hg���¼��/7[(��/;l�o9����=jTO��ٻ�.�1����c��s�v�L�a!���@x� 4}�5O>k�cӑ'3��\�?n�ká�]T����:z$#���h�}� �{�Q�Q��5��/��#Zg^U����ĝKuC���]�g������@OU�,x\7H�C����E)���Yd�j��o1#��y�����~������W��xD
_j�$�POF[�f�j��s[m�K�VP�$n�i})�p]q��D�>��<A�������,y��x/Z��<l�$��v�!x�-7N�E�d@�������|7��ݶ{z��BՉ�Fg��=@e��+<�Ѯ�;7/}�]b�0�w
��(��ưE�������ʪ<�݀���g24+�n�^�����Yqҹw�C��F�#��+�Ey�;$�^�|����͔�šP�tSV�c+���|�Dz�t�j΢�k�K�c�6�2�4-s����hv�6繱�l~���W_	����=��^�z�6w�s�_�.�L��G���G���qf�.×g��o�ͫhe��R�]鯥�b��9��H�X�K`��|e��Y��0��p1[~9��_��O��h��d�8���5�Ō�kE/ΥHp�*��a�u�}�X�{�
��ڎc�q��6��[ ���b"���k�V�A���%�{�l���<#>ز���r���F��bT�>���YKK˽t�_9�V3���K닽��&�u�Ƙ�x���U	!֦���m�6UQ���bK�n
�/+�g¬C�F8�*��[����Os�}��y�٭�P �X�R�S(P��Lި}���`:h�d���]��'/J�^�*��I�`���2�=�ifS����S�R�/�x���"H�e�E� EO�4��n�}"�8ᵠ3ϝ͂�gH&���N*KWNn�%�'1�����S\Ma�K9&�Q�,��ץ�>Gl9�)7�vk�������̹��L��ME�dq%��^�-e��Z��}M��{<n�t��߁kq%�tb�J;���_DG��H1�����L���F�*�w�sg�X��!x�%8���\ZX�8n�����y���P��=��ٌ_ABJv�6g���L���B��Jo�θny�f��:J*S皙wk�o�+��(h������X\�0�s��������wW��}G$����Q�8�k<�_
d�~=OM>E�Іn�t=o�F���1]�3�:�wYLߋ�`�_���^<<J�dJ�=KG�'<���ؾ�~X�̩P�WVwQ=k|^�)�w��$�������{�(8��}�y�v�;�ga������`xP��N���Y~�:cb�T��h2�2��3�V�kP�2�b���9Q�Mk�-��R�rݩ'vc"q�Δ�C�ci#��]��tё]�2�n�\O&����D|iI��"�L�z���}��]��(5b�c��3�<�y�jk�I��{���d�&������-���M�\&V�>WJ������!*;����DOW��� ��J�:���<�gu�j�o{m�|V<�e��ۯ�I���#wr�wH��DP#OqC�^�y�5+��İ�Ĝw�SrsuDMU��{��ac�躺N�$�)��������>h�6��]�0X�}H����A��!�J��G�jR�M"�H}};w����_Z�di����
�2E���K���D����oO1����T6k?CM"�i�,o
d6�Ȭ�n1��zl��m	2�!/i{�i���J���e�(W�)�k:*~'�<a=����*�.��a�\.0_�޿�)�᠎Ʃ�ݻ�gS*Q�Q�ǌ�jPzz�>;����GB��W�`T�=�t�g�(!)%|��hU=�w0R���/}��惬��!C6�b�Qr�%n�aѤ�QP�'X휧�=�:`�pT�L)�hT��A��P�Fs�ي���Cv.�����̻��ww����L��L��^�wM�%^�a��0�e��ׇ|]�56s7E��Z1��ul0?}ե���o:�ce?,�49����/
�7^*�:��J�5��D4=]lb1���J�G4�Ӟ����,h3=��׽�GΪ��1uP\�W���GCś�q� �U�$�w�����q>(A���!�.��u�^,�U�cY�׻�������S�-�pP�6��Ԇ}Α�3���y b�X%,߽�����qM�q��ѽ�cp��<���N싥,��%�hAS���x�m�$kG@�L�H^+���u�z��OX��\�ԷN��C��G='��1ġ0��hp�q"����kY����T�W���v�HH�y+,̻�v��B���t%���#�-���(�u�֩p
�u�̉c�S'�9����}v0�HM��2�2
�#������r����Pۃ�A��B�CV8]�V���l-�K�u��#(3��/��#�����
l���L���;e�#�<�����\TJ��Y�� �0ר�õ�{y�x�lQ�}�Y�2KV=�E^�]˧�1&Mw�/1��~�	���u�o�B��p�6�.�X�u�	CBe��m�7�3\~��c����U�R��q.��x����E�6":��ͯ'�o�\���O*�yhW��`�K�~��.�j����gyf����9����o&�0{ƫ�x*�6'�E�W�Q�����5֬�f�J���c��}�}k"1�2�K`�񋇯���Y7��M���:$�~S)W��'}��9jB�3�x��Tb�bVw�)[������^�I-�wμ_&d�C7�E�u��^�|x��Q.�򲣨�^�re���3��&�t&UlYX�"���W]�1  ��`�3�k�l�Soȝ�a�t~�9���9��ߝC��u�7u�sͤ��Vnq[�#�6frO:;a�S��q<��mo7�]�^�1��h�_�d�����t؝�;g�Kz��4���iW�*|��J��j���S���:Uջ�0x��{�O8��%�GyR��tv5�L]Z2A��f��V����ڪz�8��>�!�#9o��BP�i3��Ѳ�iL�j�����u�K����\�K�c��>5�G�S��iu�
�"ʫ��m囯%���v����3r��^��͇���8�;.�Z����y����^s�v���@��<�;�%�7.�Ԍ�H��9�Q������˗9¥m̬Ӭ֢I�B�ҡ���_28�iY!�Ȟ�wt}�w[�K'�W!�
L�cr��,/W����r�iy �Y;o:HȺ^��~uǂ��p����z�C�=�U�wZ|��Vt�	jϷ1W��@��.����+Պ��  ��k3/̺~�Mw�,e_ʚ��f��S��w++��cN�������f��Ô���}�L�3��li��5W�J%�W��aw�72+��d�a:�=]s�$�_��5xط�?�Q7��*K�蠐B�@���X�hY1�L�d�q��2���Mwc�LA�fS�)��;c -1b�:�J {�7�nI����E��̯t�{�5>C9w��@W 4�;q��Z��yα��3��D�4x�w�p�������]�[Jۑ�j�f����$�{TE���E���#3�˱�����Ky<1zbv���a_��H�]�R��$�B��+i�b��q��
�a�W�gN̗�������ù�o� i�!t^��S���D�O�r�������W���˩n��`�݈��T��d3��@ޛ;z�}E%�8u�HxD����X&
�IV�"
X�r����龗pR�Z<�5�&���<|8^���R��`�*�����X�f���Fߝ����W��]��N�)q�'`ڴ�
�[�C���kc�l<{Q;�ˊ�|w���\в��;�4U�μ!�+p�7�iNL��0%��n�j�G?)������&��x�?%�S.���@ծ=��R�7��.��>�G �V,{)b�LZ)�L�#��v��
�z��y�����P	���zwu{���DVKU�zú�\V��x%�^��Z�~'�`�r[p��Z��B��tʆr��M����Eާ�S��׽�F��zgv�\� �(3BK���g���j�{|p�Ç~�����Y��c�wJ�ҹ+���0�/G:�ce?,hsSW�P�̼7k6�Ƿ�IѼ�(��QJ(kThp�S�jdo:�Ӟ���]~���(g����0˂���)���]CeSz��Y��>�=�K�o>�ӕ��铸H����7��B�2�C5R�nW^6q�zo;a���=���3B���|v���;e3�4��u!�<f_��4;�C�@e��rҮg'l5n��;*v%J�cX.B�6Fsw֖��fvZ��)�w�%�$.�s��w�p�	<w�X�T���s�Ի��ifL���}��ͽ�R?(T?��Ǒ�{�����t��"H�N�D��
�\К�dUݱ��VD�����ׂ4�`�ʳ�w���Þ�^�F�io��q�'�����x?]��۠&8p��#W\j]W��O�
Ă�Z�C�8�ƇI$3�4�u\}��3�Ƅ�BP*��uu_�����7%.���@���_Jj���Ʃ�D���7=���,�]�
8k<*E��GmYC��@�Z��?�v^r�t�������y����&�����<C1Gh��Pύ�e��'��X����mw�ޒ{�[�����ńH�u4�t�E�A����}dAnM��>�-����oʏ�=�bW�Ci��9S˃���3/�{|�{$�*�1����ŕ�-Q�<�^:_J���28���6z�c�Z_;������o����n���Y��E�\�l��]��7��>D�g[U|'	l�-�u�z��0;��ǙJ���'�s��x�}�[��S	�sdn�S�}1h�9���k��Wƕ��A%p�U��$�W�M֫�M��̊���|Y
w��u^"�f9#�e#[ݾ.7>�kx�D\8�)@���;~J��rY��V�\�L�q*d�jg��Y��ks�m�����$l4�w^YI�@'ve7�
�a-�.�E�Η�ϜX�l&ڔM��ot�a�q�sNZ�-���M��t�v�@M�ICʜ�l�����҇&*�2�Z?05HB��{���5��8�s<B�
�]�JwxK"(;n4�T ��<,�J.��+}�!u��]wD:�,��I[g��3�|E������t�t�3h�]J����ηW���R�!u�ʉMǔ��Fb��Je鿘hμU,��6�y�xAhJZ�+2���,�Ш[�V��2��;Sv�ށ74�3�R��X�-��;8n#~��}�                �ގKfO\ס�/,����Wu�N�0��������Na�Ɗ�Q����W�U�lO�Wh�<l����̀L37]���כr���>' ��{�eN�Ĭ���!�;���A9s�����-��ws���Xn�"=m�d�3qN\����v��Α�r�ȠF��5f��yAR�mJ�A-Beh���p>j�u���s��1�`󏸫�j�$���v�|2�n@�%z��6�`Q����>v��sa8CY���F��u�W*�zU�e��>��fot���Ņ�M�!�m��5�8b��#�&��L����N�;aTwv�e�&(�
/0��tGH�Y(�їԬ��8P;u	r�VԎ�\O: ˭rpҲ�Fހ19Y�s2լ�v��'ǊUk��%j=9xc2������wxc�(�8f��h��u�Lٮ/z���G�b��o�ݘ���mm� "% yV�yx��;h�; �U��8m�l���]��4�4sc�sJU�,���ֳY�FfQS�f��F��URŕ94IMfePsd�TA����5��E`��U/�dfX15�d�a��	���ىA3LQ[ڌ���\��#SES	����Jb��VFW8d:�$���i�N�H����5�A4HZ�55��"2��r�*��b�EZ�
��ZH�)
 ������ua�"��9�Q�EfPd�IBPSu��E1TM2TP Ǔ݈�%�y��{L����u��WA�P8�<r�6�u�@�ȤX��9C�){��P�Wgy�;J���uf\a�f�Zȋ@�A�^����,�2uv�~�Qjs-�'��A:����/����^Hi�b�|Y�z��VW1q�=:�-�����u�4����2,+�z��ǀ�R��-r;���C���?h�X�/�V���U)�V=oC$�����s2us���AKL�T^���P��=���u���LA�{A����f�{zw&��N�d��A�V�림)���F8�/���9V�}�7�k���GN�AhX�
^ը �uf�mC{(f�s`EUX�λy�cy��h ��ފǅ!��`$p����x*UVC!a� ��Z���cߘb�����Cb�.�x	�!	�{.�9G�3�L��&�����C�S4<W��$�tb�J2���H��H�~��K��U�b�˺x��cd�s��*�ӴR�О�d��:K�.��V�g���z�
��ifSQ�#���'1�_1��u�Vh�s-U�J�]{V�٦�������P�P��<��>�[$��^��/�e?"J�@��mS��%�#��U��<#t����&��@�8�~A�J;j�}���+S?g�2�*�K�$B��qva�6����!r�+
W���/
�X��:��v߶;���l��|G���r�-\���i�v�p��e,dU�3�D�M�U�u����oI�l�k֘�:6�u�T��] Ua�ω�	u�Q��ٽT�=W��t*��������5*s�к�����*?��0��1s��w*7U��$gT󂉫�&.3�H��Ɵ'�Gc��v(
�*�O$��̼K�`N��,u�8��A��}6Ƒ�B��i�ե��N�&�0��ύ$NJEC�T�qϪW5��iBQ�4o[�����FW;Ѻ�� �کVGoY��̎0z�չ����,)�b�ttS{�R��3���*��	b6k��osJ��#��e�d���D�v���ܛ��7/#{#Q���]b��W�r?�\*��V�ͻ�G����M�y?{]���������p]�/���|���&B�48N�����^�sn���p���%Ktí��aR�b>$�s����B�?>���M	h�LƑ��0�<;�8�`�_;������=�nNv��d��T�Ӥx�F��؋P�������W��@�Mq�ηɌ�K�G�Z�֗˳��|�0�u�J�үzU��'��?tVL6�ӷ�V6Ҵ��"*��l��8Њ�A:���&+�|ݖQ�w�b��Q�#)rŪ�\7D�|�=|�Tu�a矻L�i�!|�,�D��~�g�>:lj�Y#�ڜ6MOJ뜱%���ދ˱��4nP�%P�L�T/������pᡋr�OMv+=3���ۡ��iW��U��0����X����49����]R�����e����oD%�(&@^��Ybn��w,�c�km�Ti\��|-���T쾠��<�I���H��1��r���&<N����4oy]�7˻\�S��n(Z�����~~��o�LX�!��T���^\C�A��s�;-\���9��=�v�|��}��f*�[}@_(���fR������&z�~cK0N�6;Mf��s�Z�B�2�C5�K���R����rmf=���ݦY�*{U�4%�&�:z���,�H��^.;��K���>5����IL�=Hѽ�a��X̩�}!V�8l'Q8�w�9���Q�I�3[�L�v_����e#�3�*͎��N�7~��ec����O�Z<�K���:Z���N���m!��'����� ��D��5�X�˫�g|�f�Ÿ�KC�|��_X��<�q+Ύ��1����TV��Gp���ƭ;�����Ȝ�'��������J�_tט��i(�Ñ!֡�Mv^�t@o��)�؍,���n�Nl�%LUP�9h0��龽�^
��$�`&M�7����1@�ߗ@���O�0���L���ސ�n�� چ��E֫�T�V<�R���WU�����{Hd?�e�������"����T"���h�vz���H�����+��
��e!f���ritYI��=~�d�c�wg�F�]�|~�^<��qX�`��X����]�վ��	��u_W���I2+��r��<KL�D#V��Z��y8�t����"�M�������$�^ͫhg<���3B�dVt �U�l����EΡ��9zH�t��Td�S��nw+/��Vڿ�E��=:w�e՛��{ѣia�\��3�l��P�(^�|CW\O� ��,�^�ޝ7X�U5��^�?xFr̆����2`UK�V=oA���'�)�����q��t8ԥ�_�.�ʡ�g�UZ]��jq� �#g�R�%���2G7x�A*���^�/��\e�qw��Z,-0:�龼6����{(s����-�{jH]��z�ZZ=�(m6��gb�d���)�Ef�.��NV��M�O�=����Ee�Ҍ��.��%�U�V�����q�������A�5� ��bH�V�P��먓63j�C5�i>�5��=�;��b:xvEc�|v##�RU4߁�}e���r�oݛ<��������KG�֫��
�
Љ឵�xT�N�ގl� �;ȵ��j��<�9��PIC�e���##�^V�'�k�l�f x��L��X�����^��8�踴��Z�r�JS��[u[��,� p��v���| �P�6;L6����\]Q�q5��{�����^B�K��<�U���N��69d�pO��+Ӝ�;�&�F�OX��㹾��ǼUm��*{
�K��옡��S�5�y۠�1%	N��86S8�B3�ߎ��`5����&&?V���~�y�ghh3W�W��cҧ�ə�\�G�՜�O{Ŷ�
C��3����2Oh���w0;wx���.��ڊ��2��2+�3o:k�i�y�`,�Cz���wB���Ҽ�X�F���ӄ����]-�u2ޮu�R�Ck(�5%��FѺ�z��I�RV��`b@tx@���O<�f���7�^^{{Ϊ�1+KO�8�/�yN$|�rH'�1�����g[���>Y�Sʹ�  ��<A��y�-yA�|+\QT�Ӊ���G���/�F�o���Y@=j�dv��tyz�E%�Q�/z�νR�Q1F���~r�H�_B��;#{�B��u���UL���=]��l�xʂ��x�2���-�1�L�C�ǚ)��r�\~�rٱd��b�Hz��aFwPq;N�b+��qmrJIH�<��tT*�f�#����,%Jj���s,1g�sߖ��`��̩��	4�{	�C��ū��!B�"���˒��lzw>�<d����9�b�)b�*y]!x�υ&j^-�Ui1�'ƀ��0���c����v�{�/��/m��lF�=b�e�N/��o&��,�6�WA���\��� �W2b�)3��V��7�J%p��nh�Q�?��sQ������#�w�����L"��Z��j�иn�����a~&�E~����zߎ�ze��-�_?\3�2��᝶Dg8�*��vd�sS��j\t�~���q��c13�_(g�Ʊ�4*��e_��ҝ��NK�$��t�)^*Ǩ*�q��0�zPȵ��榪;�͂���E�۲cC��xl�
�v�J�W�����Ƞ9�f[{�~�%���mcQ�̺��|S?��6g�lB��W�P��%�2���ٵ�m��WP!�[�G~r�̺� iR0T T~̤j���7�׼�{��"Xa��A�����5XB�k u���v�_V>s��Ä�>N��K�?/j	^8.��lU��R$D;�!u��o�Ӣ�jj��YAB/��l�$U��Ƈ��ʲ��f����]����4���f�� V}]�ޞ��	�J���:��v�Z��Fc�v���Q,	%k�o-����b�w�����5���x�M��Wq|�\��nf�f>�������K�މ�������w냲����֟��D`htww���ɝ��yy`��F�M\����Y����#��^oFω�}i��ڱ�Qx(dB�����]�]W�.����dviޮ�p���	J�0�ϥ��H�4`��DR�C�_��ٯ�d�3�t&�j��@�(/J���A���p�P�"��Ž;��^��'e���7��^�;�RńSb��4�,�%"c|4{��]v��*f	�E��#�vE�U�b�8k���/��p4����ϣ�����G�Zgg<������|�#e鲎����\]��&gi���XnJE\�sj����Ҙ:q�;x�ꑍ��2��z��g�\ڇ�ˇ�YP�4;LFX*㾛�qz�ɍ쨝`�/0���0s������WJ�����
_e����X]�}�a�B�W�:�61@u�Wc��\�rh��b=Bڋsh�Q��ͷ�����m�n�wK�n����~K:�k��u��xBpr0��f�m����hf�s�䏏찋�I�I��,Ŵ�˯�]N*ȇ�]S;��hp����N��*���Y���H����KL�T^�"��LUA5[�N5-M��V�^�x5�}�
�$ljixK�Aq���P�,'\w��	ShU�L��d?j��| �S�ABĪ��j?]D��P�=��ߟ�:d����.<<ЂZ��X��|���Ϭ���? ��V�kV�ԧ�xq-A�_TP�X5\n*,����Pd�dX����C���qI�>�p}�-u�=�Q�C1T�(z��h�%�7.��o�#�_9[t�A(�di���]n!z�Lr�oҸ��5�{�������yA2�zҵ�D�b��P���m��:",�]K.x��+�r�ޥN�4�\{��Q ӽ3�HPRվ��j�+]`E�	K5�:��Ҥ�
Y:����O��
G��#���OE6�5[�|�Z�����QYSj_n����.ν6�)��9Ow���j�Kp�ī4;S۹�C�*�l��$�5��DV��{�B��Iun��gϰtd�/)rL�Ic�.ht��u�ml��g;�4�۷�/�B�v0��|��[x��*>�����W�bH&gkɍ���lM�n���v�;K������X�e���9��=R�e��NR3y�a��-�zF&����.T�����Ys;�hF���PM�BgF��{7Q��]��^�2qZi\:�ݪ6QGp��7D�N��O�Q"�d�B���F�&ՈP�3�v�{m����Ms��d�^���0'����h;& {U{};6��l����92����u��W��T�����c`�5>��\lmt;c5[��]��V�VR��|�Ț�ϙ�pk+�&̮�2���x��dM���.����$"i#���ͺU��T/X{�[pv�!                	7�m�G���곜��a�u�G���%����ܪ;�7|h�]���4 ��b���*��Ԗ�J�cd�b!e!�!U��ih�$��8������|R�{�ɞ�ݢ�xܕ&!捉.=Y6.��v�0Q�w����9��:i.�J陼P=���]��WAb��v�^F-k7���ĕ�:u���&�����1��&�0��':�l�$zU�v�'Ss�z�un�mG�����	Mגn$7tX6��
�_-	�4�pV3� uER=U��h��.�֑d�3�\bҐ��Mj�V������i�I+9c*y�=��]���'ܽ�o��:�+��*n��+�*�m��I�)��e��RG)��q��ݒ�����XF"I���,dpo-��->�h�0N�3]ĥ,�����I��"�UÇK�R��/T�6�����_o"B��4�L��j8^*{��$��b,� Z�z�;"&ou(�@Jq��rF܉�
�C�+�@��ji���������

YD�R;a�4�Q�2�(��"jR�����*$��JH"����,�7����i(j���d��$A@�-D�,��U-	ԙP%1%Z�ʶ�*�hh�
����������{�
)"��J(�I�*i����(j���iJ�"��.Kݒ�!B�D��TQM%4M͑HQCKI�[�ES4�R�PLIT��KHR�U4�̱L�Х4QMS0������s�i��ӈf�u�K��Lzt;�o�������((ˬ��y��ج��؞���5^N�=D��}��}��=}P��0��ip�����SGE�B�<8Q�W^^�tp�{���s�o'�C�W���o��jlS�
�j�]�$�Ap��]���ojـ�r�c�%m;Xpl�q��=����뢂@jY~5~�̴g���oU���W�0l���}�V�ؿJ�A�f1r�WVk=M�^T;$�z�a&�XtN?/��f�o�L56/ah֢�,K�rq<�����K\lYu�`�c��>h3��w�pg�o/�,�缩i����ix�` 4a/�mY�o�����>ē�6��V7\~�$�w���̞�9j�{H�U ��I�5��,4�V���{��O8�}E_����m3Fܾ9�����GbD=�/�ҷϧJQ�2v�`H_��3@���2�a�#��.n����-k��ȗ@��2$�kh7F�ѶI�BC��o��ڧ;�����2�q�*nI�v�NQ�����饤�����#z�;��J�f�M��I!�M���6y��O�د����B�Ň�����L��Q��aů�vD<w�^gL�wGY\�'٨�b�I��.�A��f�#���(��I�Ni����߿$e����>Y�_��j��.Z�T�Z�L�"n�YS2*f��+���R�܈�eV�Y��}f#N��KdW����>�6Z�]��K���h!�Jg�K�Y��������%�-��u:+:�)�u��������Q,��yC��x�~�E�R�m5�ܛ����q����/�7O�)աƤ��3�_(g��������|�}{7yZ`�漢�����C�g�
��T��/��X�?v�'�:ϫeX�6�J�X[@Ԯ7��4{�İm2�T�>Yie�]����k۔%O~��9^5��R���� �b��K�V8�	S@~�Փ�������M%a������c��B��xW�;ł�L����f��
�w��vbCu(�M���S&;����KxIu�V�l��;�5r�A%[D�#7 ������5_�fgObM��{�.�F�7�6t�w��J�ͭ4+S!�D2��X���߫w#���:�i_�\_�z�g"�C^�|�	sp���,��Ε��q�s3�p@h�B��%��<���7���Z_��5�k�rH׫���j'K�ȭA�6eZB�].5�v֙�^��O���ɺ�笷�:w�ĝKuC�*���9Z����9�6��=������~���KT�KZ$��4-%�0y%�%T^�},���������3�Q=6�n�e�(^����]�^��Q�e���{<���|��A*\"�<}�6��GMY�H{�fP�I�\��x�i�2�؆��J�:
���o�A��<G��T"����Oy�wdi�(����Y��/���gW�6F©����S�ġ���ўO<�(���庺{��k�ڼT���Ѝ�J3A^p�c� h���[o{F�p�n����������LN�������%';&r�Fp�v�yh�q?�;Rl�?���g����b�(K�*�p��\Pw�ׯ޼ަ���[���o�Mw5{�+y`���䡱��#�!��6��<j�N<n"���8���a� �۝nmn:��0�3B�E��
�W�L�q\Y�I=
WCՇ�.���x3�,9��P�
��t��e*�'�*�=K{�#�*�{������*w��t�g:���hf�Ȱ���蛨.���=�����Xt�u�`�����VDNV��V�e1ȯ����CL}1��nnq�Ϋ�$O��)iw�켪E}�ߺ�|nR�ˈ�v瓊.5�{��hT�D*���  �|�A�0v�k�a�뎠��c
���M�ޣ��[�;�v^����h8�������"�u^�C`̭y�����PǁT4�<ЂZ��X�H}���xj�0�i,P�k2�P�s)�y�P���-�G>юIB+��n���[}����Ϋ�r�=Ѩ�8��.�"1�W5p�_5�^����ՓԾ��<y�N.�M�����ƻ�k���_�^,�_ƫ�(�-<[���|a'�9��	3��-��Xz�-�U%$�tb�$������f���2z��(�t抮7YC"ȅ��Iq�P�=r��l�މL��;0Y>�#��n�kE�:��<��U��>2��9��7� �T�ޗL����}�]�_�F�k�_,�-}:�\w�. ���5�&�,�����ݏr���!a�������`UE<@�����r��x�{݋H��f����~ږ���f�7p�S� �Xڐ*��C;���k������Z��1p���z�_�O,�fT�Fz�Y�1�{��V1 �x�������ʐ��x�ry]�y�T�J�t'��������%�\M�|����͐<�����M�R���f&��	6،��DĪ��66ȰO]X}]����%�ۇv�H*�|�v�=���5J��&�R�1ep�ػw(	{��\��m��fAj�m��m��r9���j	��/ѥ��D��;�90�gֲ���O�zp�[W���]��Q|,�Z-�q;�~�\ց _���N3��M͝�ʂ��p�*o����v�{v�|dB!L���<`Z��j���;�p�^�}5ô`l��^r�Sh\*���g ������곬O�/U�q�DoNW��)v'5U�5u��s�B=�d����97Z��D�|��a��vq��@�Q�Ƌi=����=�T�:�ݡ�1��z��h��,anV'ƻ����=O���x9d�m��W7��fzV�wyf�s��#���㣓�F7���ָ���.��yhi}f<-k��I�sw�8��Ѯ�{�_��;"e���Z���P���k���bM�
����;�k�W�5΀�k/����hGY�]l��E��WF�s��?q�������/ʲV�~��s�)�@�j_�&��o���OY�d�dǰ�����E"�y*�uH_ts_�NޛR�]���]GE�׫G���$�z�}�x��8��H��!7�퓧bW;�>�ۯ��y���l�K��:OK�*�f��ԭF���=��Ru�}�!+�����7��[)f�)(���i�Ӌ��ә9��o]ǇQ�{�r|m��-��^M�DsK����>�2"��9@����|�^�0.�n�;���Y[;��vz4��~u,Q��h�,���xK�]���8s������q�M������" �	}��+�(.�f��W��3�-"ӗ	b�楎���*��jL�irk�5�y��i�<<1���ݣ���uܭZ�<wQ�;I CInicYK�$p�ڧw�U�\\���v��q�~�i�$��R�5_�]k�%���0�e�޳�^��z�#.V�;S>�d�P���I�F��}��OT��WڽT:2��7ؠ68n3�Is鴬����:��j�7�*��=�u��s5~P������r��J寕�H�eeVaט;��u.:�Sz�_K����_�ufIQ��I�Q���s�@n��?���;u�18e�1��\}j��[Oʄ�_GF��a�\�<���\b&�9�[����2�������)C^�g,��Ñ��no���~�㓣f��o�	nS���o���ϱ*��󸄭���[��u���2Ҹv���-	I�d Z7[s�?JT��P�}�X�W�J�6s�ѱV��K������,�J�_�Ky����]��O�B��͵V���B���$�R����2z����Zǝ7�9U�uw�s�έ�J��	�F�'{�|�G�֋M�F���/N���{M/^'��o8�8�[�d�u�O���,�`;����;(h�}�DJBY�Dh��=!����k�<���<��L0k%���}<�ޓ��-�@G�z�{��<��H������J�&F|5��Z���.�(y^Y���߭��'���;ʽ�.UU�t�v:22../�gR���9ͲusZ��^�7���EZ���*o�}�|�Go	�ҙ ��tǣU�8������x����וf���@eDrsQf7�޵����-��]�Y�����-� ®���^\�n�bS�!aܸ�]���`�lN���-9��B �$3&�ܰ�/�6�<뮜���#ǋg1V�h�l^*;)�;K5>���e�ιԯ��A��n�Z8g�V���z�ίZ�I�سz�Ή����^7���Y2���K�w�J��8�UZ�!>���6����!���%\;A8�-[q{��E+���3\7����}���c�T��9�͝����sGn�Z�Nz��+x��r"]�Zu~�ûnw��zly���K{�T���A������73�����"��U!w��=٪�)i���k��1b�H��8����WIW���O_ؕC�W�+��ȼ�7���d���&N�On�w���|=�ٚ��M�w�ypn[��ǕLꞄ:TuFluv뾬�*���Xu����K X��;���,>6�;���Ԧ�y��{�uj&&e���+�����6;�̨;�����Uc$R�3A���&��/�<�f�E�{��;�/�PF��ǍC��Z�eG+�ԥw�-��Mhs8.�%�,}\E��A�>����!�l@&U����a���{Ud|���@"fI)��E�F���$����ǃj].������c�F�2��}���
��6�78��A���]pG:�]2,W�B����;�fT��9��8�I����|��$nOUݰ+o}�Ә36�V8�:W]��:���75�]�Z(n-���1]�u�I��q82����%�[B!v��%��i��h�u��N%����Ů�+�OU��G;GP��.�g%9�B]��D�{��u�_��4:�[��^�9Tӊ��r���R�u�ʍ�v�ևo{lF�P6X�n�,1rn6��
Zg�'2���t�Գ�Ns���z�g.FQ��A�鋍.�ٳ��]�����(���:z��u]\�WG��                 3c�v�D���2��H{�/Vu�J��<�X�wfn�-v��]8�,}�����wc�q�+��\d2]2�oY�k�:ZۛZx�����#�Pՠ�Œ��
��I��@{�6+\�Io��U��'ea��]�[�s��]����1���T,�+�P�S*ﲳ��OEƀ����Gi����B�m�Z�1%����рi�ʄ:�Ȅo�;��4�qڬVqp�G6�N�O�%�3��N��@gR�/@(V	��i�1�ջ�������V֫&n���a#�n�)�//l��M�E+��N��Dkv  �.�*�Lg.ȶ�{P�2�n��:a���n0Q�tL�ꎛ����u<F���EWor#aTWO�Qbr������>�X6��T�Rѓ\��We,���K���H�.�os[��]Y@RIb�nc闼��Z9������^��U{�kȠ�$w�Yt�����P[�ζ�������{;�oy�# �� �~$ HR��%#E@�7� \c�����r
v��c��)j�Z�A�Z]A�Ԧ@d�T�H��2��P䔍&I�)��U
RP�'H�
ChrfҴ��M)J�S!h���'hPP�)�P>Y'2�$H��aWd�9��@R���B$���� %W��d��eno�l;�u1�;G-�C�6�S"F�CC�ua��vչJ��ģn4��3Ooz?{o(�k��{����	t�K�u+�"�Xg�mZIA��L�����Usj�&PUn�����9�'��u�T/������=���J��j�l�-�WGP�}�_yTE�n3���cc���Yq�N*d��oZG�Z�bn��0��>ۧ���ΌH���$��c��ry����w6��_�Gz�.,s$�i<Zެ��s+�w��]QЄ��yº�ư她ד��Xl���G.�g�{~�Gl�5خS�9�K�0ed^o}�m	���ONB�f���l���ŉ�Վ'yR��t�`��*�T,��%|l��E~�b�'�2oث++�6<�Y� �K�k�)P���fʽW�Eᗙ}���Bfb�F���mtxn]�%�vEܘ�nX��Rq��7[2�V��<�j�9���ʐo�5'�ƚM�W�N�O}ξ�U��s��^vRl���"�v�k�&��W�
 ���S=	�֊�yq={q��qs{���)��oy�Բ��s�F�p
-.^xL\2F�4�{��w=��9�؇WI��Q���hЌ�Jb�t����d�f��W�^4�����	u%�Ng�$�3�K+�S����I���)�ybu�o������l��k���6���˓��N�^1�Zi(��([x�c68M^{W�z��[�:u����Ïk�~�~���M���I6��&s�&�%��r���� �+�j�V3�(�����sdd����>ܞ�9��3�s7R��M��Af�[xj��z>��X���^��1����K��3�kdyr�	nD(�4C�n��ҷ%͉��q��Zq +:l/'K�]JПn!֮䆯fv��tg=�'x���3�~�Ky��s*�=�p�P�j�uy�L����]+�5�s�9��fSy~�{^N�(*��Vsi�d�:��}9�J{=[�'Q��W{xY��v9�o[�e(ct_K���q��J���O�U��;q�UGl�uw�sø��~[�N��ۉJ�y�f��^����k�D�ڿ�����/���Q�/�$�Ýj�OGf�{D�k~�oF��^y�F��K;O����lyhc�r.�+�S.c=z��� ��9�,�W�U3�ؽ�B?�yn�6ז�;�je�7\�x��p�������{�3������9ߛ0�G�Hh�R���M����CWk�+g7T�`�N���T$��. �g���3���
!u��Q�n�f�&�P������3�t�5�0*�G����\j~�=�o!�F�~�muSW/�ҏ����ۯ�L�x�T�*�\����:ql��5ݰ�*��M<��l��։*S�ԧ5:�龯N�~��*u�^,���������u�����e~����E��z�7+<��H��ټ�f����W���������3R�~̫/X���]5fJ����=�W��bY�^�m֓m2����Y���w^V�u9V�y͛l�U��s�e�N-�]�p�'nrV��=���Nw�j/.�^+�Ob8�	�{��o�̉;z+iɤ��xs�|oq�>����bf�_������W���u�z�����L�@I��bũF�[J�'���4��a������w��NZ����eE)iliu�rL��;D��;w��.ᘅ��V	�j%���{�J5r�W���_�ю�UD��s�=��()i���]n�s�!�/�'��k�h���65�=�S]��y?nߧ��,0��q������װn��xb�(=�%hr��ם����+��g��f�*���yy
�<�������j����}�,̓k
IT�ܛ�<k q[%@nw�6����}��'��]�^�B^�t'^���>�v9d�S�ʦb��y�.�x��%�d�=�n�oC\�L�갷�ӥY�O���jە���_���7V�|l��};��MG�$M3-�=�oy�%����=�<��%MeQ�5��s,��;�E�m���^YqHF8ngX��{׋�k\�/S|:5v�Z�	j1''S^��19Zy�<�_t�e��ܧ����S5���M��\�W�����ݵI�Ӷ�렫�t5<e�lrTkBkՏx'SB8ycz��G�ݲWzb�;=��+�YX�ѥ8'�\��N��fN��V^���O7sH���o����]��L��l��\�����"��5���v�O�^�^~�yZ{x^'���Y�o����w��E�r�>�GJ�^����G��g�7��r��dq�]/�{3�dy��2Sy�L�)�8LI��n���ty7z��!e�ê��B��Y�6��z*��XS{S�܀��;'	�{]w2{zc��T��+���}3K�RH4��1[�f��ʒln�</�8�;jlsǲ��n�=�k���FK���yin��7n��	M��� ��o����oxN���)m��pٺ�e�X��S$�k��J���rG�5�l�]�䔡��g�b�������)���B�7�S�frڝ��U+�wѾ�Wo��>쪻^��Va���jh��۱��Z�>���k$U�>�謢*��arn&�=�c���d��@����9�*az��z5��r�N79^�#�Qb흥�B����g�ʃ��@�G����EhE�sYΣ������`�2�R���~��U�{�슜7����4����V��ۚ���K��P:�X��I�>�_���Ni1<��hf��׼�K��χ"��	̣�?(ϥ�T=]��秽�K��_�nw`���!�Tk=2r��.�j��&�[GO:E
�Uаr�ێm\be�|�o���s�(T����!N	�J�'{���Χ;��@v]��C[�[�3:⹢-�L�ܤ�S�qC[�K���	RԜe�2��~�o]Q���b�_LV������Who<{�އ�r���F����Ч�<�B�6���Ss�,'f���S��۬8�קX.��N�;�wˢI��3����w���uu����b�e��WE��������%�WC���+"�����o�X�#93��z��Bsje����;��Dq����ߩ]T]�N�O������μw�T�������!�˛+<g������o�s/
�����W�׹=�Nɞ�����W��E�����Z���)��}��ܑ������fd�[�2h��!�s��]Yݔ�n�
Uy���̷	5gSx��r�K�S�5o3�1�e��h������sv1KZh���Iy���ލ����%�VG�;xԒ
���vf��.l����+�z�0KxH�AW9����ry�7�U��^�/���&c��k��_��$M�Ot��gX>ډ�U����>o$z��pZsg�y!�&��'���;����o����q��#<}�m�F��6���u*�^��������l�:��:��e�ҹޞ��W@����|7��ܞ��{���A���my��;�kl�!_ ����LS�2��u<	���Vx_�{��590�'$�j��a�]D�q�<�'��9��yW�rv�cc�`9v���K�=�X}�b�����׽�L^P�%[�poCgΕ��} }ﳄ�}k.�y�݆��}�-�7,�+^�d+X�ˠ���M���F��r9�����N�V��+�5sm(��$;0qi���� ��༳)�v�CG3�o�^�o#�<�hk`���+�^�:����1�f8pFwE{=�{"y~�sj��n�𼣷�����.�	�=X�̄Bgzv��o�9��U���S=�eT<��ۚg���ݹg+�T��=�?m��+0�����±�M�'���^���b��+���-û�2��"z	c��[d���~0j�7�~��Q���`��޾�1�˼�{�ܓols����ns��\bt��\lޣ������𪮏c�T�6Vv�2�>]��guƯ$�&&2�&:���7�4Ӓ���v�9ʯR˿��5\�}U���Oz>��y��Uk+QC�g�!������?�?<~���ʏ��h������SV��AE?o�&h"���'�d��?�a�h05��:�>����?�}���w���<��QH�Q@��(�a���( ����;ߓN��nbbs�h1��a3����`|3�_,P�7L\���u �"��|�`{�����-�������4��c�<.����A��l`tl'!��\�<�|:0x{������As�.�ψ���D�������W���X^@>�QS�B^PTO�!��Rb��������'�����A�N�bm�?��A���I���p�C��-����"�A�T���t`}�1���SB���?TlBr�8�k�7�O�a��S?�ə���X7�~���� �s�����G����{�� �GGѹ��;��Ѽj��pDl� �lm�-�e^�ڨC�����2��o��ۮM���!���l|��)�^�����8��;�G�m��~��n����o��p����?%7�~��n�������������j�������QS�qg�H}A��p������]���8���S�O���}�������kq�����}��t��k�_������9>��E>�>�X.����?h~��q��7�DG��y����L'1M�B ����H"�����Gan|�cX'�h�?x�|l/_�#�t�S�n���iA�8��AI>�E��C��5�(")�.�.����}a���óͯ��e���\���0�W�Z��;y}͎�^��N�@"������O���� "��_��B��!X>��� >������||ρ?��ԟ��~bh�� �����g�4_3��=��������O�M����&���F �"�a��=���|���f ~���/�A����x]:?�?����������O����'����'<�(���~;b���~Ȁ������������T���?��W����'#��|��[}���A�������m�'?_֖�埧��:#��G������'�&|s��WF�l���ø���}00��)��e����??�N�S쿃�?��{���E>���~i�|	�N���`�2�פ?-ks�>ILA}���O���Gߛ�����)��g|�