BZh91AY&SY��_qׅ߀`qg���#� ?���b@>}@  _YT��QUCf��m�l��%V��6d��(UZ�)SZ#f��QJ֍ikQ5�h�l�֔֔��%j%���m�18[e&M�ԭJ*ҌF���ְi��M+6���UV�eV��IZ�ֱ@�j��fSb��ͤ�2eVj�6k@�dU��Yf�f����N�,d*m��SV�f��*��M���ea����S-�m�Ҫ�Zڶ�j� `�h��S4�6fU�U�����T�S`�l��e�Ƭ^N䵴�KF��  :�ᔡ�V�յ�EKDU�������l���-��V�ūU ���ԭj�A��I*�]�
&ړ�:�(�ڶ֙lj�(�ʦ�  ��(S��7e��@	�\���Cs��t*:0
 �Ρ�@
m;p�
;#  r�  ,��4�*�efbV���kL�  <�(v��0 �m�:  �`m�M맼 :S�ǝ�K� �X�@�u;�����Ӫ��p{�{Z7�Cm��ڪ�m�lkM�  �x !w�����g��:P�C���� X0 �{c�z �x �
\z�����k�UJ U�W�=@�i���iMYjj�i�iUCF� �� AD���� 1�����  �� }�f��@kA�u;��: �ݧ��(okn[:��(s�� ��\��X�m�����ͩ�ճ�  ��(��n�Ε  .��
 +���J����R���N�a�;�9��)n�� S�����M� u���h�[l�I�
���L�   �{��\�΀h� ι�t
)�&�
4��
 �w)Ӡ]\ ;��ӆ� [��4j.EYl�Z�̪Kd�[   1�  ���L ��S���m� wX� ������� �r� \�*� cuVZYl�)&�+$�jUme�   �x �  ,��P;�8 ꋹ��(.�q� �` �X � 4�P4�ֶ�,blf�Z$҃�  �����B�v� w��  � �,    ��� �� ��  ! �T���M��*�	�0b4� &�1��1JRUMh��!��#�"����J0      O�OUU �4 �  R ���CB���ڞ���j=G��zA���)&�$�)�M���#��F�z��yy���n{E�+�υ�\޸�k�f�����1��|�3�i�iW����3*_:����� ���Z�ն�v����~��m����{}����wA��*+�Q��V�����������[o����_���si5�&���*����m��鵺kn�ۥm�m�[WJ�-ҵt�]6ۦ��]+k�Z�m�m�M��Jۦ�鵺[n����t�����ںV��k��j�MV�]5���t�����U�n�Y6��V�kk���Zɶ�m��V�5��骺[n�ۥ��m]+k�V�]+d��m��mt��Mmt�]6�魩*��J�j�[j�-���U�tյ��mVM�����[Z�M��t��WJ��ҵZ�Z�t�ڮ�m�t�Z�mI[m]+m���j�[Z�U�]5kWJ����Z�j�]6�WK[n��dڶ�M��t������J��J��魭]6�]5�KdںU]6����Ut��V�����t�]6����t�WMj�]-��j�]+WJ��j�V����?�^�������V�S�ѡ��j�]���2�]hY6�C�0^Ӊ�y�l`%���I�7�S^k���7Hd��ڱ.��Ԗ��U�z���7[lܷ[&?�?fnݪ!�\	^��)6�]42dY	rL;SA9)�v3(��ٴ�n��o���M�X�/p�.�����$n��8����7HJ�&v0kr����)v���U����n	�G(j��%l��<��M�y(?�fL9�j663&�q]C�7fU�n��r�)��&��2��E�:%#9X����kMId*��B�
��`8Sa��6J��z�[B�Rn "�w0Q��3M%��][464� ���Q���mk�r��%%�D3,KCi�BQڐZ���u{F�@��>J���2$P�2�<�[��Z�n�T�M�MX-�t�Hh�ikl�o:����.lS�������i>A������i���YXXWB�-i�M^٤�f��X�o]h:T�eA(=�DH���8�a��SAe�ȕu�Z�[F�rnc
�7)P��p�kY5ԩ)�����u���E\�L[�֝�N^��n\.�[��u%�L�<�V��)��	{Y�e��$Ԯ���_c��Ɠc�U��%�(�E��X%)��G��XN��(��e\��Lj��(̨`��t��w0��(��&CEmd�CDOZciS7��5�o	v�/C2�6��z��Yn��t�W��u���Syz�귍3m�ǎ���e�Vv���x������;�����0%$R�79�n��T6�dx�`���jB�9Twx)Xe�-l�y:�l52U��ڛ��q�f6cͰF�3Ք�Z�P��h�n�,�gD˕���R��?Y�7,Ce�����[�ǃ����^b�����u��U��ƺ��W�ݚ�
٭���ZM��ɿdW�r�w$�͙��N��2�]GaGYy���H�
�[/�۟M�-�T[����p	�V�_l�@�J�I+n�*�NS�(Q��r��I;�����M��4^bUkaKj*Z�S�r���w���X�J{x�b
���� ��$�F�tژLavwuS�js0��4���h�Pl˴w5&	�m����r����̎Sǻ�6	ƥ#�b��]n9�l�� �Y�QDk�NƇf=�{$�mm��m����k�P0[�J��-6����Zx7F��=E��t<䱰�xH`�H���5��4��աM�Y1�g�O,�Ub�̺pI��R�d��U�i�_GYXEM.�*K��*Amk�#O*V�3$�,a�< m7��ŰP�&��.���$��ɢUԶ�]hW�`i�ݸYW[���H��NM�J�YKl0������ތ�%��#4�jGz�J�� M��+�*�
ʹ��^�hb�s�Ŏ��[FJ,))ܦff۫�Z�gn�ց�ucY�J�dr�9�o15�Y�P��-�N��Wx��j����Q;{,{�lu2Х���v$%�1�˘�[M�W�dUɄ�XjJϮ#k�Rݣ��Z��
�<��"�cǀ�� �鳹����Bt�:`q�T4ųv�![Vu o-V�zu/Mŕ"�gZ�"���ر�]na�jɲb �I*9�m٧zt<�� x�cI!�Tf�1���.)
'aâR�Y����aT0�V��A5{�cx�hXnk8f�i��ܻ�gy ��
�}�Zʻi��Z�ETZ�A��æ!h��;5���Vpd�iaV�Y7*M���%�P�^R/K��d+;*���<vCG���,�v�����B�if�ۇS�?�۳yY�b,���R)�+f<R�L	���a��+�٬*lֱp�dknI,��/u50m5���e�%�uy�֪H��7l�Рu;8��vo�{�C�LʔoTŸ�b��U��cj��VSq�F!D�$lm��.��5T��������X萖����w*���*�Cv�h�
��+6cF�9@�[c�R�'1��eE�hl�r���+��G1�-խ��
C`Vjf�w�J�5f�.����ɺ(��1�����]Z�&� ��i�՝kU���ݳ�B1�aӷ���Rǈ��t�b¨�E��R�(�)T��Xº�F��x��4�IQ�ᅞ��ZGÛ�*-f<��.�(�������c�H����	��J{uͪ�8�Q)�m81=f��P�˔k\#�1@t�2��,�KР��C4D��vCm%�7 ̥)m�9�_%�զ^�Q�4�.�*�tf����U͵f,tou��f]�r�^�Zf� d�"z#���D��6�YH�p�mb5� ���M�H:ul?�[Cr��9�L+h�������A��[��+:��n��h
<�q�k�%4�!ǗK`ø��4���U��n��5�-�R�8έ)\�弗�jl��M�W0/��բ���6�ju j��E�V��U:B�:�Qb��5���Q ��l�R�Y�ivXsj�V�����C���hu/���I數�Pm�R3tS݃N�ֲ� �c�dT1��9��!3��^��N�*��h�e���%]lj5�(����JOj$kJז�U�d�q!Led9�T�)-�Eգ.���:��g�i^�Mne���5R4�{�	*,�y.)(�E�bѤ���I��!7�l�P�X]И�#&�I�Fǂ-+f9�� �;�5+켐�V�({Yq8"d�qR�7��n(�����f�u�� ֦��T#i뼬�o@�p��,����n���LG!��XN��q��[�%]�Vuu�)R���A����Y�����7�u<�e�[Y��'�U�w2no��gb����
z�@��7k-�Rǌ[��2�F��Ӻ���'�fV)Yˢ�=�k*wUa��h��[%��j}�y��tvP˲�14�V��4��9g���j3[N�KB��r^��Q��)3U��<[�؉�/S�͠u �㗗�5���H�r��9 :7��F��nѬZ�Mkb�ܱd�e�yJ��CUa������9mˋ�B�))�����vv)�i��7�%n�]�	^�Ti�R
lŕ6�[�z�Mn}*�	ImI�l�q;&�َ�&�͕�\�P�L�J�2PI�ʻ��VØܶ~Z��M�/p���J:��~ة�ɌԱ+��mh��^ j��oD۬�n��X��ņ�%iK{���,�h��Љ��R�R���˵Km���:�*�3�U����4�ع�uJ��Rc#* b��dy���bw,����ֈ�A��.��:Ȭ�2����<�RjՓ>͊�H���1�H��ʖ���������{��)��kh�Uw��<�Sklʒ��nJ��&��-�rV�"���iQ���t%)��a��7"�5,%C��F�j񻪵x %"`��M��G+6�u���f'Y{w��b�1�*���%�(;�|h�Ƶ�ͺ�{�+/Z}z���{.K8��K��n;
�Sv���1* ���d�P��wg���ع��x	ݖ�f�M֩J���D�p�ړd�F5�t�n�̔�Vf�u��5'&L�5c�2b9r�3e�R��mi�gT�fV�KX�X��XUa�&� Fe���B�<Uw�=Vd�t6��f�A��l�ON[�f�,Z���5��İm�Lh$2nl��be��z�6�
��̭�y[�ڢq��U�-,S�2�hMJ�b
�srQ�Eaz�j�Ǐ.�व����L�b^f�h�N8wR�zML	Z1�SS���+F�4��s3/{�bJ܊�c��KR��� !/1U�'>3H[�3�f�0M�l�����8~�3[E���5M�N#r�Yh�[�Rэ���r,�&n�&�1V
u����$� A���H���xq��-��M��,$�LK/:���{Yl�{�,<��kIa�{�H�+^���쩋��u�SX����.ۼT��f���A2�v<�Kq�����]
VL"Lb]@(i8�[Һ�x����p�HT)��a���(R�p�xu%H�v�#ۢ�(��!Z-eаe17��.�=6"L����RR�!X�*�;��}�+8�Ɖ�е"k10���Y>o����n�c���&���tK���6�ǭ�R�ς�K����Ty�eE)�x��s`�i*�&�5���-ʊj��?�c�t"-��b���|BJ�Eb�E.Y�R����e}����@YX��WLc����E��H��eɭ��༧M^�V� ���Ak�I�0��̋)�Ô��5�EBwN�z-;t�M��٢��g�sL �#;x�87��81�+��V[�1�Y
� �/N�D8E,г(L��=2^Zʉ�{#���ve�b4��&��6��3	�-�Su
3H�6V�č�0ē��0ι��6�c-[�=U��(�u��d�_H�ɶ,�)
��>{I׺4}��V鄖�v�ɰQR�Y�3�i�<WZ�YD,���0˭"��HP��D�DK��f�ג�Z�pb]<�Gk5���˽66�ta����R���1����
bo�)�iX�d�� �p��f�M%�A��m%��C��*����,�T\�opcwY�,�.��$P��r�Ѝ�Jb�)$���4��� ��y�X�7Ud�M�@s7�����o�����q\�3Z�Ҋ�p�3i��7u�����Xά.�BѭLҒ�$1�aa��2XW�ΐ̶1�� #�Xr��;HZ�%�u����\��LK�=�ϯR�����2d
�ؠ��\��m�0��d��G�p�.��i�����=���2I��'�,k��r����JL�͹MH�%Q�6-ذ�|֪���A�&���֖�'oa�X�� H$�N�@,e�H�C>���ƞSsjnfk��2Ra���0�Q�S+#�+.
'6�*��Ej�=�og'z�J�l�x���^�	hw,�ʉn-���2���D*m����ŕØ[�9�\P�vB�i���PJ揶��7C�Y��@�*c�6M�IGa�ʼ[$v��d��R�n����2mЃ ��a,�m
c)��.)y�QL��8�*�o�<5͌���E�����M-�ZCѸN�n�/0��o)�����̰�E�Wf�Xh���*!�}���ה7@�-��������V�)��I��9[W�Q�V������1mC���a�9��-��m���W�j�>�o-1��u�vlQW�j���a�WH�*=Z�t���2��G3a���(SRd@�l�P4q�m��ҡwJ��f;�y�F�~x3TܩJ�ELa����)4S�Y����9��V�!
Q�V
b�.0��on�"�k���7	��c�U��mA�%����35X݉��L�p��os��D�s[V+p���tP��h)�$ᱛ/e;,ZĻ1�U�M`�(�X��.��X��[��XU�Y���3A��e�y�1Y±��5�e����Q��t�T�"�]X�7D����*���j,]ŷ����pSq���Q-��4RR��Ieb�k
�̹2����4
GQ�F�E3ldA���b�
,Bo+�,����hd]�6�BSı���W�;�Z��h�c�v�90h���a�+F���O+@ݶ�G���Y�)\�� V�1����%�©�1
�	(�i��^e�Q�[�,ۭ"�#�E�k,d�؈�1B�[�nK��wЙ����[Z���� �1��0�Ѵ򈽶�{�0�<���y��d�b
 ��3�)�f2��e�Ee�z����k@7�6�$ ��43w�@��̲�Kim&�e�F!,�u�(�u1rN'k���]If��E]�ݏre=�I�x����&)�V)k�RF\C�R;ifm��6bЩ�،��ܗ���ˬ��R��;Dˎk�R���t]����Z�ɴ#*(�g������l�5{�J"BuK�*�ct���67��i����M��#E|�j��^nPC	6�d:��YIiU,�A٦I*� ֪k��&3��Nk���sFf4�z��s�l�����)k�p��F+hd�M�[��0g�*A�q�oo��ELe���V�j�V6I�N N�V�4��1P�+F�z�݂�n]����.R��]��髨KL��BLHf�w^��B�9w/�t���CAM�Q�2�4��;�B����Bףp�e�Zu�IRAL�|���P���F���;�҃ �0	Ov��AX��vHwF�
ͻIm����9�3w2I�˙R�b�S�E���x^� 6�j���;�����F͝��l�����Mm
*�`]k�uʯ3.�\�^�th�w�ެZ�� N���e	�d�'VK���X�Xr�7Pn� o^��"��CJ�Ul�[L�j�[�V֊��PxM�y��,����M�qƯ��Z`�Sӡ�5m*�!i���������ό���j}��,����r��T0�hdP����.���[c�����7.^顅���ś�uӊ��G"���ٸnZn�TT�,,H̒�W�Q�j����q�7p�8V��E�X�;̡����)�캁��#��B���h��wsșԉ*ix݁i����`����HwC�:���p
-��U����8�E�.��̝��O&j2��`ǂm�k(�	�(ݛ�å��Su��9�vWu�V�#��Z�D��,┳j^�U�'q-60���(V�c�W�õ�7D���8&g���n�Y5��ۚBUpU��R����u�kߜy����|����b̉.�[-c8��C6�O�3��tP��&�:�&�=����Z�j���2<8b3a�#Ș�n�\U'
j�,Y���&ha[��@Op���!��{�bZkq�h�W+��?�g��V@��߾�����?��h���@��\(]emaH�\}���Br��JYҦ��t7��0�bbN����;��/"")�QY4+�y֕�j�Ept �rAJ��ع������d��v��pީ���u	p0���"&�\r.�����H�<�Njč�.��z�od�d��;��:Uj�`�Iz��E�hd1A��
�C��Y 3�u�DV^^_o�m��P�eМ���z��}�6mh,�vV�^�f���Ν����Ѹ���>+�db�f�_8$�m��%�S+;�MDV���9��.�t��b.���݁���-��e���Э���<�W[pR�|r�76���&�b8i�]% {���Dޖ̻�|:[�ӆ��s����I��ҭ̊뉌�GT���bu��K��c�ǀE�uʼi�1��W�b�c��.�q�d ��jPTp��;9�Yz��Gt����*�iym\�8a��e䘋��.�X��sY�w箠٥��U�qn����O���l�Iw��5=#��Kk���0a6�t�{�<W�����R��{b��tځ��]��|Bw�3�8�9N&��˒����%��0o�')�ۼ�t����vE&�d_Z��)��Nj|
����X<����Y�!�J[���v��6[�v���p�u�I���*h���pͼ4r� �� k��D�U�9aG�ɕsUB��� ���M�$�Wԥ��wTa���+��`�	R��չwb;l���m�iєH�LwQE+fn�{�Fyk����޹�)`�ش��M�9CY�.yu;�����aG�����V�x��`h��`���le骊��u�t)��3��ٮ�M�1��M�݌�,�+��חS6ڣ�B��j�p�$�`h��F�f�Ŭӄa�3X�+���߳��|�*L��J;��*a��'b�D��D*p�w1ϔH�q�\�d���	�ʺ���Wy�(�YM�Y����:�r}M;̞WH��&CUg���vv��zW6�
ύ����В�^h�u<�C3��@�:}�A�+�-!]��f��h�IR�Whn�;�^�-ڜ�2����m�چ���V
H��1��>&�*�{2���G�Y�q}
���mԆIy���Ѓ� άx�dw'k)�N����c��1*���l�(�5au�w��WàM���i��M��X�ML��aȴp �J��,B�԰����˹y�3�e�j[��o���*�$w�����1����E�rgL68K@�Ey��q�]ө:u��K.�[���S1��O�.5�OW���P;^�Hv^+�,�/��Ӈoy�VZ7NC�I��Go��j��|\r�����_�ѡ��3�j�B�v�Qa��|��MK@���'c���v����@����2j �a�F���ǫu�E�g]��u/X��7����Tor�
;z�%˅d���La;z��s�bo9������L�����7*3�����9�)4ΕY�Վ
�+vM����}���1�h��k�;�{�'�[�1�,j(����}��
��un
qǘo�S�gz6f�����-6rkO+�sd���-�Ś�}wwN��3(�ϥ��N�8��ѼV̤3Nܧo��;k��D�Q�0m�&���X�Z�*TV�n����֨9^;�C��j΃E�]jķ BC-��-:�/7',Ճ#�3P��ݞY���p�j]��f��f�]@��9�ɛb���ȝ#����ݒ�@�o�V�T�-*뻻��v2�u�Gj�꼧Qh]f�,˹�� 9+���A�����G2�֐C̱4�s���.�����͠�؝��ũMb�m�N�++W+F��]4�Sʙ_ y.j�,s���X�}��A
��uA�U�lfѵVp�r���:S|���%��=�O_�0j���_:NW]q���m(�^�c�r�K�C�Dx�r��=O�,oZ�*��G�,�� ���T�ʆ����ع�cs �T|"��L�ys�� ʳ�gsQD+e�U3����ڲ=|2��!���Y]���F7}%\�$7��/^���,vC3m��ZU�*	�F,+w[�DǤρ������k��ƉH8��U�	��9��	81�o��Y�bG);���8$]x���{�8��jyt��k�G/�;�@�;Q��b�_`�t�ԕ`����zzlv��D,a�$�qR��\�+:�X#��H�{;�\�`�ר19���v� ��M�F��}��mb����s��]�UȺz�g�s��T��q	-���f���� �W�U��ޔ(Jڲr	B�9�{7��x�vJ1cfm����G��'�Ъd��_C��1�Q�nmͬ��+���OR�i*�9�p�"�|L�J�ǹ��Ro����4A�2�hs1���\��"a�wRè�۰�6��ƪh�F�߷�;&�M�1 !\�����2�1��g_S[R����ڄlI��Ꭶ�P�#F�_5ם�w�H�_nGL9�Q�6�H"Y�^0�"�̓�ea������Lö�Ђ̆
�SXx�j�ŎJ�'e��[���nT+��l���HNX�vL�v�.��P^�Å��݇3�i�_RY%�Cru��Ŵf�rY�,5 �K�z	K��wc���V��_�Մ��֥5A�׭�m:��_eK�9N�$rD�ެy2�N�C��4���6���=��iؼɐ���D[��\�u�IX�i���<��.H���_��x`.�����O�kb��:�"��<
��������α��p�i�]F�bɼ��=�Kާ8Ȁo�̙��'K9f){�jģo$"g�M�+6�;�:Ρj��f[�7�����t�\��lR�|;�޿�\���ݩ��i�ݛ5�S+�H0T.����[��Ҭ��pM�&u��Lh�-P�vY��؝]��4� �>�=��|�9� ۣk&�k�A��!�8֗��\�5)��W���J�]���{�����+�.Sևq�`�R����#/��C���a,���B"�5���R�����r�R���YQ���:�[S��7n����P\xv3��/c�5>�hZf ���Yf�{N�vQUm���P��;��#5$���*����ޅa�y��k&��h�*��qJ�O'fj�ھ4 �K��Z�Ʌ}�s�]n��j�7��zY��V�&T��ǔf��q ݁�be
b�R+�y���nc��B%��:X�*�W>Y�`�����\�딥��f�;Iވ��f�*�������&ӫ<1�["bX�-e�	��>�-��S:ѵ%�X٭nwAzoil��̨�U��ΐڀ]�Z�oZ�S�"�
��%w3'^X���+Edi�Ԩe���ԏ�e�W������*̇C`Gf�T��f`�6*�����)�e.FVۗЬ�j��)�b����^N�άE2�Tx���X�q�tz4��!���:�,RI��Ӂ�AY�5�okU&r��Pk�dXU� <H)Q�ѝ��-��.���J���aT
��^o[`ҙ�
6�-�p]�gAEG�7760/�4s8�q!�1�֦��.�t�.{���*�f�,���F�O��ʐ�$����k"q3�m���(!�Q��݄Ag�9�3�CbLN�JW��hpv�r��`�݊D z�Z�cfR��/���S9jd9Vk	asv~Ք��Ч�ՌF�>�NKYv<L�f�o$n�vA\t`$	՗c�$����䈙�Y��-� }�{���d.!!yw�]�qQ��h��L�����iGR�8�S��d���V�W�	�;�+Dr� ��YÈ㗜I�9Q��P&��I�v�n��.�v�Mۧ�G�k����Mھ�₍I]��B슋���Ģ���wC{�Dd��X��I��×�d�V�%��ꕩ�ۘ2��4!ݩ{��ܝevE��f��,)T��'+��1��J�2V�c��Xd=T�f����[����V��t_r�]N�5glENюfn��Ύ�n:U8�YJ�7X�5[|�6��v��
wpgf�Ni�D�&�V�K�S��7G�-2�k�mC��%y:�I0(�i.̲U�S�ݵEC�3�ki���� �X�Z�6�,��lv��VN<�B��]Ǔ�����6���ޜ��6��:�c[1✛8%0h��;�v-�^�ۛY�ΈV /x�o�p�,���q*�����c����"�tu;I�*�6��shY����a�%_n��y�.84��`��xt�Z��q����6xeEM�3��h ���n^���^�����2g	|�V;Qa9:��{,������N[ue�He�}4)[*��J��؁�\�(�1ެ����6/U�9
Z�ԍ�w��8����ƖV�g�H����������@��|�%��Pu�ɋ4�g���GVY��ALn�i���Fs3��Kbz�`(P{�l�-����8�pe����ח|4`�f��u�	7��4��]]ҩ0�m��)Cɞ�f�w���u�0�:��98sHv�X�d5�K��,�\�̋sQ,goP�u5�z{S�k���N���U��u�90�a��pĳ��\��z�;�V�"W4QYM4x�a
p�5�e��|�{�حWU��,)vＷ��m��
٫N+����Rb��v}��I1�\�Z����\
t89҇v�{ h�q�ɤ� �oY���;Z�+��5 �cyt�1wS��fΤ*���!s�v�:]bS檱�:^��
F��[h��i(�-Z �Ó�A���W.�5�]5����e�]�Q�]W��)��߹
�셳#�@,� F�"�z�^+�e��K���<��͈M�/8ۀm'ʗ9u0R�y0�r����WD���+s�wq<�$UAwY0���O�����S��V�V�Җ�^��'
�%6K����AF�`Bּ�2NͶ���[����]�O�f���`"���v�$�xYTu�;-�6s>p���걺k�,j��n��E��u��;j�].>8pA��:��T�!��vԋ�ݝ̧�J���c�������r���=��;j�Cӛu!�.��v�؝"�ot]Ң�VQ��	��,�u�hjB����]Ne��a�{������
�4�Suz�ays��SOUK��p���GptDr���KsGj���u�rκ�&]M�ײ��jq��i&N���V�P���R������|�o��t/
s^��m6+�M"p�.T�SbWY�97;��ҥ�'t�shZ��B��N��w嬛/.�}�(jR�*�`J�<R�IwVU�빖��)����9}�
�TR����kF^��_��.�EVz�5�Ua+ǰ�W+zQW�ɯF���A��PК�u8�x�vA�c����.ُEYi��D-^<xn��U��)l\�TLY��G�RU2������Й3B���9i�.��p���ˆE)�V��9nH%;a�#z�]�7h�l�c�1TyB�V�'�@��&Ɗ�4��Vw2[��M\�j�Sz��5�7� 	aQ��e�@�M���+#�&��Ҏ؝�[�7�/wf2��԰��Nq=B�7����
�G��M|!x\Kq7�Y�c����u��k�Dn��c]��ɵ�;a5���.�v�H�(r��,��&��)���EW�F���Q�p�����ous=�PHm��5MC��.�(� u�LK���H�9��$w���!_cT����T��QVaIb�}K�v�،e�������ѵ�SN��Km�r����7�|��3���v=۴�j�k2�{�;�Z�q�l+�x��*%;(�[s0�,��#fн�X�r`{��ټ_X��$�����������Nf�R�ha��d�P�Z��f<�� d�A��[(,M9׼m��;6�t��]}8Ro5��SM��[���W��_l�9�Hn��Qn�[W�%��	���g���0L�a��S��˶La;PD�2M���q�۽U8�U��{z�	�P��������"�1�
���ۻ�Վ9J�mkAn�mB�+Ɯ�K�ʧ �Ρ6��(rU+jg�ڰuTթ�ufl�]��2�y�ѱ��AI{�`�,�y�n��4�D>�N⸋J�ƒ���
�*2�^v �U�M(Xl�)	��V�v[�W2� B�p���EI�K)G�[;�Ч���r\'�l�W����Zp���]�����8��қ�i�攟_�S��hȨ:_.M�ok������j�_,��-!;�Շ����ܻ�)����1|v�	�[9@�w�B�_(]ګ�'(�3iF۶MՕeՎ�f�bv�����a�{��'�9��/S��b�(��Zfp|u��q��.��
��7�v�襪޴�aZ;{���<�9VgS�ƅ����B�4}QA�%}�/[gKVv���&L���7Ș<<�N��]>�pK��҄`s�ky��ffܳpH�JGJ�72��$���,��	Q�k	���)�&����f���o�99�:�h� ��",`p�V̊��;2K�����2�X� >���'E���f�Wk�J0Axw�pª_ @�}�)I_!��b�S����}׋Hhǻ	�l�w��It�Lغ\�]ݖ(�ɽҍt��>�Z3�+o"�[��El2Jˎfj�x�v#��(]���8 [SfV*�����]�?yWj:~�x���^`TG���]������R�c��\�ʆ
=��1$�X�#�1���eP .ͮ���##�8�F�p\��j�I*�J�rM8�%��;+N�Ώ�5[Zb� ��9�~,f �����mb� ��c��У���M@ۉ�>�S������`�i��
H*�t�8�j�M+���a��E�a�
 ����mЩQ/�V�o1����-*�q�M��(KK{�EWSߺh
 �f�iQ|���jx��(���zg�u��볖��{qⷥ��˾t�1;Y��/�Fk[�g�EU���;�'B��]ꭨ�浀�����F6nW���n�;��Å��s:zk�K6?��Ր�KU�UqYD͜0
�X�\	O��8�r�*%un�O�)tz�ZM<��=7d���˄�7CVY��SUa���D�e�ڄg�l�>���xU�h��{����e!u��kK���=��}���s7}Iq�&ވL.�ܒ�m7Oa���{�ӌ/���G[�K�L����2Ĵp1ف�%a�9g�gXg�n��=�~��v���S���hl媕 �c9j�|y�{_eL��q%���}�|ț�yPe5�h�GN�/�e̹3��qm%�r��ءkM�F�P��
(';d��n�,W<{9�	Y���<"��]�>�a0�gYcfK��J��T3͢�j��/z��+��v9e��O]�Srcld�a�MӸ���u��V�םu3@�y�����3�+�f'>6(H���]	������ʬ���ܝ�V5�l�k%�XE u�rc�M������L]t�`A�{
����T��)(�̫f���$1X���k�+�v�7Wɧ�9��w_���h�A[j�V��Q֪��rc���2��ڬ�;T��:�1�d�.���S��ь�Q��9������AE� �0A �A�@ �$H�AE ��A@� �4��t/k*��6��݋�����2��69��́�F��d����ʔ��� �5br�j��)�hQ�7pe��M��̕;a0���9�3���� �r�֖���w��K�<:��F�\��V��~�F�+�ewH��,��U�[�Ox�Q�j��{d8w���)9`D��A�k�2�[q9���#Z�vӂ�d��-V4�+������t�&wd׺��q\�㖕@r���m:ǎQ�%�v�Q9�
y3�l2e�Q_Z���;��Y�e-�`��	�Wa[L�)u���'ST���P�C��P'ؔ�
��yQR7if9K� ���u]�-�Z���ͥX�T�ɮ9a�@R;t�#�񨘝4JW���i�I�;���[`ji`r�b�]��w�b�[Յ�V��j�z5�f�ѩآe`�����n�xbyR-�B����&V\�)����x������U���Cj^:�e�8P�F�X<�B�*͚BsJ�oY�E%��ޣv@�d��UL�FR		Xn�Q�_Y��z��!�O��E㭂��6�����狪У�wP]ѳcfk{ɐ���U��<9V�c��re�ѡҬWBþ����Hݪ�S�J`����6��c=����/����.��-�5�[ńg+-���jiҟ`�#�fIW�Mݠ�ue�l2�Gǧ�X���+�@���,`����� �#� � �E �(P AA��AAp"ן�����K����xζ�<vЮT ;x3(�f��ɸ��@*Z��ۙ�Q�\4��^�t�V��,\�5b�V�F1s����Wgj��T5գ�a!�&$��"�`���i�n�M��[�[C���ʺw�}��6\o�A;�@Ҿ�cKf�C�Qִ�j�g(�M�-]_n�)��]����h�h����B�X�/Sa.��7N�N�u�4d�0Ma']vݨ�挵�m�d�Jʙy�uriԕ-X�&��p�X�ﲴu�Ƒ���Nf@�6��^P���u���եw���i���	�*T���y��S����A�YÇ�:��^kv�������[�x�5*{{�k{�E� ���+f+�+�Y��\;���Yܫ�N�)PcwJ��V���ua{���/�b�AV߮��HF��4��K%�(����]M�"�j/'Z�3��v�r�ˡ�#��7wւ�S�0zIU�TTi���-�����o)�OF�|�{m�G#m��-U��bt���dmq�ulĎ�#�,��(�%���vښ�R����n�kX4ԍ�b�)����Yc"��2�}��,g �E��7�gŌ;[�������:elSgW��B���Ҷ�������v������go�mD�Y��p�t
Zz�p���oqj;2�{o�3ֲ*U�bE��S�W���g/8>�{Mz��#�nFj�wi��3��)ʒ�
B��aC�#��[n�ɴ���4��M���&�vbv���PvflCC��ɝ�@���t+E���u\@\�4�ִ�Q�E})j����)_U����Ҟu��7ǒ�h�O����ѨǗ�J�QN��L�Na�����-�o�U�[a��ά��Ǟ�H�h)e��*V�f�Ts����&]�N,�p#��w��gN�Im!thM��[V�n
��Mgt4l@Kx�ݐ�D���Qh�t�r-��O�L)�Σtİ0��K��+l��#�X�7��}I�#&q�u'�x-f��Z:vcv�([�NR�AL�{�[���b��)	@�zxA���Z�N�F嗢�˖@�{rܹ��
�ݤ�kf<�D��O1t��Bg.:�'�2V��ʗY/�j����9�V���V��E�ڹ���C6Mv?�Os:���_-ܬ5'��g>�Y:�����a�:6@na3j��;{��U�`��ܧ�}�ņ�"ʽO�[��Y�����_�.έ���MyZ��_Q`�<��#�fu�fn���_-)��0)ơ4f\m�5·�h�	�8"m��ی�ٙ� ���w��kT)EfS�g�U�E:G����X�pQ8fDuf*��i�/����h�MIܙW�QqN�w@
�֏a�zoI��{I�Z)=kx f��L⮉3�i�-^�����Q�]o��<tu��^��'"��K�;q�P��[�*;�2�K��E��hr[�;�3�ޠ��=Z�6��*jn��A홽�V�r�Z��ɖ�B�Tn��dO�XV�5:��*n��A�9�sl��Ĥg;P��RV��Ҫqe��L���h�MV�r5��ǆJV�T�:w&R30j�p��%���-�y�;�gu�(�-�K�%z�I��TٛD]L.��]&�-�̱�
�l��^+�b9�q�Hk��h؝��=�yvAԷ^�����zvbӯ�8`S�#�Y;�<���آ��Z��fg�Qt�(�-�+0���[0��:��T:�!����.�t,ˏ�gD�L����\�pT ,�X�O��"�,RC�M��u����7���m���8;�/�3k�ʏ*������<�iJ��{��{7dKGN���sB0��ڬ�z�+���ծ�
E`Ď����� r�.�V�V��c�C� ���U�)�X�ɥr_3���7GL�R�y+V�u�G'`- �f\o[�0�@���^�r+Yn+�X�2����A�1$�-�kv�䬮�Z����d(V0�{�g:0��Zt�˶M�bj2/`t��,�:������6-`�[[���"�ժĺ�$�ALٙ�`C�p'�r���Vj<�&fU�䫤{1s���U�#Z�A2P�7�X��f���kt{&	�k3��iԠ�^�)r��b�&]�Z4b��k���	��UyWE0D*��ye<��4����oV�j�{Ja
��4���@�uuj�앖�\r�EL�aQ����' �..�׎T�h^�fn:�MMK㏊@�I��-g�B_j�˱:��V7c���V�ss��]Ī�`��^J���������]WK7���R�<}S��w��gjP�()S>6��;{�\{�k���*m�68�m%�.�A��t\w��4�B����w�)bWE�i��S��\PAdX0��;j��x#Y�����:4�)�����uՂ^nCd�pMX]��ӊ]C�˖.ed�'%�� `��f�����F����\t��}���L��JH:�1uu}�����&p+�00'�Q��Q=��n����Dʵ�yۧK��%]pϥ�^Dɵ��)PV�\);ӽ��
�
��0ѩK*V���þ��4��3 `�ׯ�6ְ���L^!Z�PN�L�Ùy�@X<��&�J>2��jQ��(�J���\�X�`'���7a��ƺ����X1�[b�J�L�L�v�@�Y��.�V��0Ro1jO 0f�N5dΘ���������moKS&��s��t�6Ugm���+��+����v;�4�I&i��7+���%]�;n�fRmB$�w�n�!��P*�3̌Psݕ�H��~��km�����M��<&c���t	�jLf��q	�~E�OsŦ��Qԕ�n�H����.�)��,����TȌ�B����o&�GO)�
�/$NQ�3Ef\ʗ�ᯨ�j�k;R
F�}i�9�_9R勜sASe��8��X��C7Pj2:�	�]�a���9�-J�̩ãw[Rй���\H%\n���WL��lRܬ�U��ķ`��f���3X�ЕҜYmoR����5Q7�{3�U˧:�GLXG[�RM�B΅W�F���Ùm��pҁ��7�4������R��}0��+/������Bʈvt�L�f<i��7*#�'7���.�TP˰�p��`�4�9X��or�'�SiZ1:È;�CT%�<���q8o8�d����9��T0�)�����6%y�ͥ/`4_��*|{峺�)�Z��i���WK263K�X�;���7��F�� �c7m�r�^L��]�k�.,�q�4v+��՜PxMJj����.�E;f�"5btjs&i��6��Wn����x���9�"�FMcNI]j�S�I����ӝd1Z�á5���;�y���b����]���`T�6�%�����%[�U9�̵��G�lL5j��EH
*�%��fu����k��T�O��L�Ǆ|�U�!)_l+y���^f=f�v4�f[�غ�����|)3n��(鋐۲��[��tqv��W���$Q�tV�B���-������ѳ��gP���sG&��^���W1K��]@^$ �4���	�H�>�Kz�q�ǧ*$�(b���)�MQ���xJ,����(�],+��V�]�o ��I��Y]Õ܏V��Y���@]����|���g4��\���v�﹖�4�ې�����H,�i��ʺ�e$Ԣn��2@u�r�j�{nK(���x�L�}r����dTH��.o.\��w�����}�@�(-��u�u�QO�;���f�5�sW�3
�3vk�[��hd��{ƶj{��C�%=�U�M�������]�RY��YaLS;G��Y4Xg{�k����Ad-��5����ۧƭȇ���gj��L�O!w�g]�p_bH�b�`�%��.<*v�23��.�%�P�౗'c�Y�E��SKlw8��H�X����S��ɬ�gk����KzZ�Y�Yή�.*y��4���'���WSݣ6�A{�}��I]�r��\#�Wc�g'fN�5��:� �9�0pͭ���.�l�ftQA1E2cR��z��ؔti:pewia��Uh嫗Wf��HԤ�t3tA�B��c�0���8���R�2�o)V��@p��j�̕�1}�[阱�㵷�'O����d$W��K��뤵�2�6ԤM���V��]���rW�.��Ђ�s37�`T)��-���n��(�a
����+#�X��Tʱ�
|y�f����z)G��Ǝ;�����jN����3�#Ytt���4��#���v����*���@T��;�*vǬK�2-�{�2U�r��U��@�)s�9KdB(�X�����\	k�;c�חavu��R���������9"<*A�޷�%��R��|Z�������Vg��fd.�n���Ltb��a�I�ճ0�-�iI��-e��$�x�-y�N�|x���6|B��X�tVN�c���F2���6�.n���$ه�VR����C�;����U�i�fw,u�6�tU,'sn�r8喓& &C�S"u��(�qp���!n�ѳ\3w0��."�F媾����G9.(���J UZ��*2 ����*J:�p��*��[U�뷓������u�h���CA��hA�W$}e�h�5�_u�cE'�F�
��ffV������ݥ�X��?3���R�dǂɺU��,cy���wR0�U��z��y �r�\��`|�	I�ǘ�Iq��A;b�J�YCEj"�/���
�Z���ٻ��Ie��%��`|�⫭��5f��ԑ�V���d��Ƙ����u������,M�bBV*P��{��*�]M!r>����X��0*	��
Ԩ��h�|�@TJA�;�U}1S�h��7��y�9P�F%{��2I1#�뻄,vJ.$[��y����I>͠��x�̂��-�HeK�h�v�����Z����)][x�Jh�����bnV�3���S.�lo��N[���Z
pr��F%�o
�f<����5s+�'�5a��|�n9�U�)�����R��)P���ŝ]����s8��vr�Wϙ�{.��7DU�t�<��3U�JP$��-8{�8��8�".f�&�p��\Y�)u�x�P�b����1����c_pQ��d.۔��}]�d�bl9��i�去Wv�Wa��횩h���1�9i�qե��fl��YIh`�%�$k[�3 Mz+T�t:N�7�t�Jݛ�S�J�=v�!#o+�)s�.c1B��:���*�+sn-���qX7Q�Y�*U.n�\ޮ�!	�1hXfaJ�Sr��0m^R�h���ڕv�j˖wWT�E+c*�t�Ŧ�Nz���ww>3��[�*^]��<LgPlKK5�9{�S�n����J�Cbc�&e%]��f ����� �.�.A��s	��_6l0���i]S_M����+d�\Oײ��w37��%*��K�Қ����m*��<F�*�zv��Wj��#��X�v�ú��ʃC���Q�q�I
���5�0b(0�$�2Lf�JeXy*�ٱ�hv"����������Nd��؄�o
��O�xE��-ڲ��X�Z��N)\�ٽqJ��Vn���*�rJvj�V6���dt�ܐY4+$b�֖�s�
�9t孵j�%l�G�ʹ5�N@����pɓ� ���v�+��S+��oW_rN^&��5�m��ȭk̕�2�9]smu/�N5��B�kḨ[
�硑���F�@롭��C��̩u���rZ��O��)�棽m_l2�D=�rr��wT�a����po�{b��4ɴC�^W�V���;Y�C��8�O{R��c*���q7/+'+�.
Y��V�y�;� �@V�1Y�D��/�U��=t�M�2�l��wO2&�r�^<X�+�Sb��RP�'c��@��^'����vP��vQ��խ"-禣쥥���%5{S�)��mN'q�R��L�p�{w�Dģ{��u��)�a\725KjT{)I 3I�_:��Y\���YrM���Y�r���9��w2�$[�-��@���lV�7W�{m�����g���Xҗ��H�C����[�; G9{�!�v�t��>��n���n�7�T�ʰeh6�fodt>*f#�/��Uy��*����� ���uq�����}��u	}-�(|�+�Z��{Ⱦ�l�⠵�wt�i�q��
�,V+��!Y$�M�<Ѣ���!��0���ʊ�j�.�r���ҥ�����y���瞻���|��Ф�$���&@�8Y.��ι̂	���7iۯW��}^�z&�������ݝ8�.�	x���P2I�DĀ���x��]]�׻���{��F��[��BW�ג�RR��:�gt'���뒸듻�wM�.�w\t�.��7\җ91�n��)7�tfW::[�Mp����k�
^7�wGuە�n�A;�ҽ�ㅋr���M2�;�w�˞a˴w(�]d�W.uݹ�$��I��t\�ch���s��r;����$��t���u�-ˈF��9r�C��4D�H�r	x�M\�B%���$&#�JD���yq`�<��wd��Rj�湸$ȄD�<��d��*;e`%|��|���������3�,�eZ��͑׽�J���J��IgLrb;��	#1�{H�b�06K}ܫ�:�Wu[��0�a�l����2��''��*����sL��J����ov��ٳ��@���ʼ�B����U���������F�D��b�m�����*�N^u��v�Q2s���s=�X���+}��h����7~�(^q��zP'�J�IXTVGD�n�̿A��`�$l�m�O/�bhv�CD��g(v�Ԓ�f�W"utf�ε3�!$�uz��M�Z���HeJ����REy�;��ƫ=�)՝���u�f/z�S�o��Rn�z���!�໅r)F��¯����ʊH���	���5[7�g�?y��{.��ZϮ���ʬƞ�oO����~<+���xlf�^.�T��r�����bc��jZ�6q�s0����P�U֋��4�SY���y��I��}�kݴռ��⦲�Ow��*�	����ܯM�R�
\S>�3ޛ^���xݟ�����/�ɥ��{��|�^�5�⚻Jĸ(���W��)\{,���w=<�W�"2�%�*�d�Z\1�6 �7�
u�:�W݈\r]���u<�e�9	뀅_q
C[��d��_,녓Y�W8��.��o+F���Gx'��qrUj�:� �_�׵��=��U*�K
�,.�HיJ�S�G�M�*A�;w3�z`2]�����\ȫ'=����z�U�(RÞ��U�(oU�4B4D¬�w����-G�`��+P�����jǅ\^��h��=R�e����Y+��8�r6;���K�Z����Wٸ����
c�'!�x�]��;������t�n-���´����kt��E��/BF��j�b��Y��� ٞ�m2�ކ^ԥ��U܂�qA^#k�,"�	��wR8��{��u��늚gW�W��~��{�u�G��f߫���4����[�՜g�T]�q{���.�qk������C%#y��ԭ��o����������g���g/�R��f��֒*��� F��V�]NϽY�X���d�^�缟ׄb��3�֒��+~��/wY:n6=�F�H���Cys.�=���"S��
���ܚ1�8y>e]�!��;$f�n.�
�n��vں�F��#�ۚ�
�(k]N�h�Q����FG7/3#̀-�Ƕ�	��!q�`Pi�XS
��`�ts�^�s=P�UdZ�c'����Gb\j.x�8b���j��t�=>����<4��~��y�ϑ�������X�~ �z��]5~���{�:^�My��^�w���o��[�s�{f�&ػ������Μ˦�W�8��ѻ6h�`�$�}"�HWz}{\��`��x�"�V�,_[�>�Ne
^�)���{����(���[(�=�'!�me3V��j����k���P���Uֽ�{�������+��EB�S���8#��;i�N���T�����y��$Y�r����ʒ�*F(�a���[AWmoҧWT9�2	��}uh���cn��P4��k��Q��[N����{�+}��&΢/|�,@�뿫���:����w{ާS�P�n�>�s�J�z��z��Y��o��yk��]^����;���$<\9���,҉���&,��p�+�n�3�ؕ��nL��ZH��g��]�"x־�蝘(N6���ِ+Z�F0΢�������ܯݝ5S;=�v��(\�8�:�r���:�U�X+�v3m+�(_W]��N{�-P}�p�4ǋr�J�h�VҰ�E��ڹ;��,�W���H�w�/�&+��V�ߨx��B�T�Q�(��g��y�?
d��U��2��2y?;�yG�W��5�8Wj��#�H�ϩ�'��rW�Obo1t�|�o�w�|��[��u�ua�z�FJ:��W@'zr����^�x�SuB6eh�ܔu|�S��i^}�X�k�yt�����|�w�O=���-������y�	M�g�e�o��L�Dx`8�~��|=��[yo�bRL�鯔��������z�.ҽ��b�9{wǙ:۔1��Lu���IU�oٞJ���7[H�Д�Uֺ}�z�l��OBQ�ˍxMr���,
��>3˰�s>���`�8 ���)r�Mg�+��ِ}�{�����j^�w��X>H�Rʝ=e�솼��Mʑoa�W>��Z�̊6U�Y��y�d���|r쁼ca+�B�?M�\�Z2h�ʸ��Ѩ<f�z��ê虹b����>-Ѝ�N��MIm>��&e�ǖVd2�I�)*n��{{{��h���Bu4���+a�Nv�����MU\��*7&9���{\j�չyX��u+���~�S�ߛ��t2d��V�[�l�E�9�ud��Qy~.��c��}]w�:��/�-�t�4H��^���J�Ֆ�T�W'������"+�L!k�ݎ��xG�A�C]n���=��ѧo ~���=�yz�5���ި}�B�$U�gVJ��ѓB�N�u��'�Ƕ�:jy�M~pi��?V�٨��'Qz�~�q��]Gi�}�DYjl����i��� �.�>����T�m{ۋ���u����/:��o�c��
r��d�=3�g�&#2`e���4F�RB��"��\9��%�A(��)I�1g�5�m��!��8]t��������{]]�{�${F�APV�b7+4�ȼ&;��M��P���d�xz~�F��J�ga�����~�^�>��cԑ�{|bߟ���kWGw�ٸ�!6��]�*i�=,��U�* QՊ��;u�_<����T�[qs�y���$і\�u˱�­9Dj��-�-��PX^��ƹ��[��A��W[Eb���S�[��#i�{�+���¹R�=%����OƸ��0^'R�I���MMvX�*�i�ba՛��;^�Ii�Pa�Cճ|�����]�e����w��w���h��Z�/c�ܩZ8῏��*����e��[�`�^��V���ti��O n�jw��ה(�j�37�{���g�����§�\_�$ގ���nw��.�} ��C�#ʶ��=ָI
z�ۥ���̪Y�8p�z�O��F��W%u,R�K�#^e*PnU�����4���"ɲ�h�&��k�+����T�T�t������^����Ң�w�u �k���
���l"���3@���uT���N[V�&��]��w�m��Ͻ�׷�������M��_�c )<x�m��+-i��>�/�A�=P*����w��^um�Hq���M����u�=����Y�����x�Zt2�l����mm����w ����O>���&��%#��<�j�+P�Ϋ�6�k#OT�E��T���[ˈ�q��^�5�.ߎP�l��7��
�5412��㸣���Xt��s����>"��n��M��>�X;$Ӯ�۲�q���Z�.�b���/��5��z]^q�ڏ9�<���ޮ��1TL�|����_��~�'�Ԍ�Ѷ����lm	���2��<zt����YY��cɇW]�F���_�2�x��߳o��վD{4X_IH�)hSIg�u�H�Ϩ>f�G�;�+i�2ܷ���ϼC&tj��-���m�Z�8�ޤJ�͢�:���٩:�[������NF�w�*^��c��ὖ��M��^}�W����>�=^C�'����K�W�V�<v�*��}�S���i�-�"�����-��x]G�(�Gծ�n�5~�6��2�3"���n�M�Y+���f�	���8�9��q���,���)���
^�����fŎG�ڽ:�k�)�c`��f�^Z�/k&3U�ʶ��*��}��_�ܶ���70^���71���lx�3�|����ρP��To��+��7�=I}}|��2�\^wۗm^=�VE� ��r���"����;�q�����)mY�Mzp�N�\����i;�"e�<�E���6����q~�X��zv�^�I��tRWu�ڜ���:�h䦋<��;�(�ʑ�ԢT��
�����.+����$=�5�pW��}�:���K��W܈����x���~����Q�D��j��[׽�G��7p��q"�Z��ψ:% �C-�y~��z��}c�=qV[>U���u��~��Ml��{ޤ��I{*P�Y���� �H&A��<�1��t��i����Y�k��c�/ ��W)�V-�����/W��<k�j�}L�`
�y۫�c�N���
������wy(��!�V���-�IFӫ�%^�jg��3�Yzns�M��⎌@l����Cõp��JR8�}�C��M4�o?u�!s��;�Hn�ڔDzA
x��f��Ii�P�C�b�0*'R���g�zR'��\FҮ�z�$��a��>�JΩ�;m+R�A��ᘷۊ�/����ʮ�Ѫ��4�����k6k�ڨt�����VG���&�{]��t� U�,��Ҁ���� ��mb�������`�x��K�zW�z�qӷWS�����S�8�="@��}�-���Χ����ȳ;�;�G�����}���RX�"#-�V��}�2��wR,N�kp؎;[�� �n�).W����Ũ�b���&�G�J`Oll@�dМ�g�hĬ���U�Kjy����GvA8�s����f�/nR��
_\�ޣy/m?5��*��3�:C��4qb������I]��_�ο>t�:�p��k���՟[5zȯN(ב�q����=x��C9ع��K�V��A@n��LZ'�#��6�K>è�6M��}�ڑ�^���w�ya�}������,�Ꙋ�g�=�f��7M��D�=�ԇ�]w��Ϩ��P^B�B��lxB�:< h5_!�w{��Ω���Z|�Y��GS�x��Z��Eg�_VJ�����₭�>6�xe �5њ�q�J3��O�{���Ȫz;)�n0�r��Ǐ���[�C�~�=��+|׽���~�v�{ƽ��kŭ�V�W.��5Ql��0��ۦ��1����5�a��˖�agKz,:Y��B_iGґ��$�̴��v�wS�pQ��純�+'!����b�{U�DY�}�
oe#Ԕ'b�%��)12u���j���­염6yϳ�����أu�����\�b�/&�"G�l+C�V��G�j��A#���zR���q\N�j�����������VlH����4I
��5ֺ���^c��M�F����k�ޛW�E_U�HeJ��{��3*;��}��^�R�h�Ԑ͸�C��;er�R��z�:ɳp="Zmud�Q隣��f+;:�w��VH�U�V�� |��
�8� JO5S�]�z��ŝ���R�/R��3(*��;�E�Rza�7��mפ����*`�U�{d�~��O�Ԃ�`/5|}��,�8��z�'�`(��g���z�͗z�҆Q㐣O�nd���C�	��T6��>�Z�I��5�;P+Z���rz�4���#S���n\�W6�Uөb�W�|1t�k�O���r�xP��[~�!֊*'�`���|,��huD��᧾��| ���b�q��E\��`�.�){��]T|�`�m��"�i�yp�{7�cZ��S!F�Y�Z�%s���r�YZ��1J@�HN��oA��+�H�1����R��Ѳ�n��U�h�1��c����۬�'�R�R�2��.��,��p�I�^��ؒ&b�	�Ni���ۗq7t���BIr]D����-�ը�/�eⱖ�5���lf��im�k�u,!�v̠L��I�ᛥ���N)�b9л W��ڼ���$`�7Q��o�L�����̶K�FY�f5��V��tA�X^&�����K�37n�W$�t�Z����l�%^�,Z���3P�ӣ�`K�wUX�d��[0�,�B���izAI}�Ku��BI�,��/Nm5��Gs�z&��X'[|Q�X;01�]c�`�C��5��: �g��[tT[��N!��ܤb��A��]�D]�.��(�..1�g�j��u�馊�淖)7y��Jzj�U]�oH{in7@p��������[�htR����Y W�E��j�u�Kú�s<*N�H��PTt�0H�Nu.��9���	�����kc���ݳ�ʼ���ٹ�PG��(��	V�p(VT�5 ;╖/��^�ޝ�ۆp3qҴ$�]�D�����SyY��N��˴6�*=�҃�,3�D�N��gKT ��Ջ����gq)J��V��Z�7�M�)c��O�_bC���5v�9�ʰw@ෲ��0�v��U.���l��TyQ�+���նx�P��r��*M|1���q�˿�i�����^K\&�aX1�7���kZ�h[�P�h��4ڕ���y��e���������^�c�X��7�N����f	�v�B��ӳ5rٜ��'��ܩ�v��
VJ���j�>I��-��d-}zV�'Q��'���-�
�L�V������x�(*�9
��
�]�<���.��W�U�,�M��W8����ƻR�^γ:C�+�Κ�V��x��7�,��s��W�r��A���#tY�'=���f�֓��=�:ݤ�̼#�=0�i�&S�,Io�T�tF��6r��#{~V��qΨ8]hF��wk;�-P���-��E�ή�\>�:�ڃ�b�e�e��������I�f󊦇9� ��>tsv�	�3��Vmd�gtf��Lh���)h�8�y2q��ѻ�J�
݌�؀ą�gC��[%Z��`�Ɏ�Y]ƍ��=��	9T�3�Rʮ50u�i�:�#mEd9Qs�R���gn]E�{'�t�j}{W�X���[����w��
]]!�l�ۜ�EqXȍ�!��PX7@��.�g!$��ٛ�4sK�ð��������+6��X~]c��M���ds�->��uo%�;s�hΔ���w�#-(�u�-��kW����r��+�=~��b�v�2�|����5}���*k�C����0��9�Cy{�_p9䚧`�W}�U
��&F&���2	^ۢ�8.u0����^^����{��|�6
�d3o��Ő�\���dЋ����ow�{���R����r�#DP&)79�v��
(N����sK��G5Զ#$aBaL1D���HQ�\؍	0(��p �E$�&4�i��y�&I�2PbŢFlR�P"X!�0a!�HA�Ǿ�1�>�0AD��ҺjH���F��M&��f��k��/]�cr��&4�V(4cF��Q���㆓Ih�KL��p����NG�}{'4_������2��a�)r� �q��g�4��W���D���7��lc��=͸�m�ѳ�qس�@P�W��xN��?���)O�%��ݞ��Z�Ė�-�������UeI�U���1d�]g痘�ղ�1��`u��9�9Ӊu�a��yX����c��2&���͡Qݨ\�^ڈ��E��B�(}ꅂ��W���Y�����n��yt.�!�V�Q��������U��-����%�^��Nl��ldτ��D�6=~���w�������8�:�_dع��`�x;����rf�Ӣ�<?r�2̲�Vp���ʫVRb���6'F���\M�;�h-*	������#�t�HJj�ڼ�M[�"��}g`�,Bb�_ᢝY^ b�w٢N���\�s�ǸXb׭�&��r�i�A��n2Y��VԼ����痪�Gm�گp�=,�c�P����r�B+��S���x���U�S���1*�@���kDfߛ�v_����O@`x!_W��(���"}�{�@\��^�� .��~�a)�lh}J[�����mM���#�,5^@�ؓbz� :1�ԠdX���gNm���
��_��;��b���y�WSqeM�P�֨��J��pZu�kV)!Mnq��ۺGd7����n��2 網
�������8�Gwn5W�2vܗ�oR����sjQ؋�K�6�����N���e�V�:����;,(z���3�-h��q�=�7����3aJH�����s�ASs0g�`
�I31J��pa��,d/��pt<�R��z��C����%�A>ϙ̱�Qb����GE_Q�*����/h���$3=Kv����_���C�p)��Ӡ�a߭V�=�~����&`F��������k̻�Y[{������*9�}j�Og�+]��Z�^@z�Xgu��ゟ�L�P�/����y/b_�+�1Du(�WOҶ��Cd؃'��8���o)�bw0�˥2<}�����H_�tN����~�x}�r��;h���,�l������"+�ELy�[�`�!�s4�4�SzJ��y#��6z5N��xX�V<��lB�O_��������C��/$�?5.;��-!�����4��N}���rf�*���76+��v ~j���f�w��3��޾C=���VlcT����(?P�x9�8��}쭩Y�"%�C{#��!�ѱ]|7q������r5�V)�U�bv_Ji��~��9z<�z-⁑�=���[Rݣv4DG������������:F.ŚG+����Zw::�B����ލ�i�w]X�ά���<���k�!C� ?v����$�Y]^�2��I��*WY�.Z�S'c�T�Oy��K;��HIJe���w����-�/�6����N��2�ּ����Y�tV	����q�.����qX>�2M8nw�Un\mXס�'#w}@x��݌����F̻��kb��G��F�RؑuԄ<�M�!|���G8~�M
�/�y~�;f�Ev��D2�D�rߒ��
W�:�3ޚ�q����躟'>9a8�������q��i�]p~��r�#���5{��*>��b�g��7�U�6$O�����(A3�Y�r�؁�����O�OgwY�!�����7�m��	څ���hW�$�_.��Q��׺v�grݿ2+�ʼ�8r�z�||�N>�r���6�)⁃Y��y�,9��c$N��!��1��U��#G����C��Öv y`���T�ft'IN�9jA��b}쓶�����oۜ�bgnD�_DJ�]	򕝗�e��8�(ρ��'�Ҋw1��Ϫ"x��."�øQ��CT�*±s4T'��5]�t{.!�zM�]�P)�
�{jw��5Y�7d��0�f�N%w1���V��CbT�M̰�Vp�"�~8+TX=�:�Қ�{;<Z��s.��ZX�	��c��;-Ԩs_�%q%^�}X���Kܗ%=ߡ�]w�n���|x�-�p,�x�@m�5R3��ҵ�������[�Fj�֝�.*7��A]�fn��ݽD�9Mz,ݯ��Ϟ�Ȱ�Sf������ޞ��#yD5���l4'��Yj���¶|j�jH�߇��lN�z��f1�t�Z�T)��^﹂F���x��M�bj;�����#�]���ږf�o��a��ʼ�E��D2c�49���<�Y�{5���1�{2�c8�ϔ�?n�S�dO�[t��9�&�3O�Ͻg{x����j��YMx:Ʃ�|���1�X�*���~X1�r؟!��Կ?�`���j9����^� "l_�E�>Ⱥ�F���|��b�p�6��z�э���~��&�Ĩ�0ô�nׯ}8:{�Nv=3B��R؟`�����(![Ϡ���ڽ\���я⪗O��n_��C���>�Wƅļr�h�_:���|+�|m�|'~���g=��Ur7��B5�E�x�T��c�K�j~~k!��g&*Y*3�6h�kj��6I��W+q�/���*~D�G��
�iz�H�.���rcCt�c6�L8"{cٻ\T!��^�u�yL�m����(�FU��5�n_��`\���\�tL���3��"v�@��j_�S���VތĤW�W�,�G�J�޹�DU�V�ԡ�ɛ�#*h���:4��̧���49���]̫��F96�c|kb@�AR�X��_P���30h|���A�c�����%>���)a������0��w�3���,Ǐ���d�������L?��H��P�DQ��3�������ݨ�g�o:$m�������uvW_{�}�
�:�S�/<�F��*��X�\h��R�������7���c��7fw,̩^����$�C�]�Ɏ�Y<U}^���˶��0�� �Bk���WO�Ӈ�e���J��*fk�T�=B ��JN���	�TP]�V|-p���/|j�h1*�nk�23�M������5���G��Hujӝ��t��B���S�Sbq�A�,�������n����_NeEu��z1��ؕ!�q�;�Y�����8Q��yX�n���1�ړG�o鲹���?v_>�<���C�V
��pc�
���������J�}���A���?����0*���ݘ���Y=O"���vQ�S�Å~��%e�����e���6�t����l!^�kq�O�zx H}5dC��㝶o�1���lҜ>�a��ׅ���.�bc}�v��[�o�㱻�܆w��Sx�%RF���ڼ���8ݪ>�A��s�vfn�expc<�T��Ձ�]��Z��W�Vg]ֺe�Wg-o`w�-&x|5�-��v��b��0��v�՝�9��'F����Ǥ�+gZi�����5��{h=�Աn�Ѥ���)\7*��VE��B{+uHh�ɜ��_ꯃKюq?#�"�Y�u��T�}h�	5n[�Uo�{l��zY�ϢO��յ(��f��0m�9�s�"��2b.�;�8;,�^U�~C>'l8}*fܦ��c>� ��"#`Ѽ8�x�����]�������b~�(S��}dA���:;���pnpZ�*���ڌ�^�xq��_0r~�f�a+��	>z�ы�@Ȟ��g����Q�u����m�Ys��#�=%˿E4׬zN|U.=3�x*ɘ�]L��@�f���%g��2�*P�P���x^3�Ms
5�o=�%iʏ5K&����Qޭ����I�"�BiK��Q��\����לT�f_eA�/��][�p5��J5���a�
{D�`੃`�����3�<��1���l>�B}
����������Q��܅�9W���Xgu�3�$l��
��F�F��ϻ���F�"�b_�bb�t��]?J߯�t6M�H]�-��0�L|��/���g�Ru�/�̇�+L�齚Y�.e�6L{���嫯B��&���jȏ�؁�W��sެ��ڸ�%��̛�VU��ۚ\�fKE���'��v�Z�-���EZ ��nX���p52�fs�W�7%��pT�RW���;���\㍪�f�u�$�����Lq�������:�2u7Q��wS=�\��3�/���7���+$G���v��H�ж��~�#
W1{=���,��d���S~����f��r�Ӈ��P#��>�2���![�?C��"$b�1
�b95}��{ �������C�<)��ܚ)�U)��k=��a�1���w�	c��aa�A�.��H�|9�8��}�ܳ�h���'�#c��X{�)�Ɗ�=Dea��7���fpI�?N�]c��[@[�# g���Lh��A_���x�;�OZ;�X
t�>_���-�{z���pH�T�Ъ������{ED�{��tTt��y�_�=N�FO� }[�~��XB�*['�~�qA� �<p�V�\��ܯ��Mj��&�b�3��m+�1ɨ�`�l1WR��n�
{຀�~���]�/b=^./���Y�c^Z���!�| �a�MFC7�ng�&|��R������W��f�1��R���#�Բ�X���ؠf|���Ք��	څ�v!N�Q *�_"��_�����]~�W[>�><�1�P0T��W�f�ժ�t�Ҟ(�هz1�@��pOF��43]it�?�~h�|���W��,,F����x�J�s+%�+�L�\cv�(	�;�PZa����� �^Û���A����*��FW�_.(>�4�c��b���^�!��cZ��dۧ0�Cw,�����45�`����3���ۋ�����q�ިg7s(@��%GX�&X8xX1���[�~�J��gS��cE�jE8�n0D��O��������tL`t=�/�@�+���#�W�.!���\��9�9�(�����{ތ�6c���c��Q?e��db��N��aX��!P�)��5]�w����J��r0oY�"�fq�3s|�r�,�p:�0UL/O|�����##"T��M���*�|�¦��r�W=�@�<�Ծ��}���?}[��if^14z�BHN�e���¾�xj�ju��T.lzTM\ǘ��vە\uuFCh�3��ޝ����-�� /S
p�a���FϮ\x����<�o2�)�>���kU9��*�H~�{5Ḳ�:�;�ɀy�f|��orŖ�#"|�N;dk��uh���	e��e��Rs�YLW��_�Ӌ�f;�a�z�:X��U���J�R����7%���IܳK�,T0u��p/Ɨ��
鱚s� �х��f��|#��=�!�p}�sW��'n�I���͞��M9��� ?N�R߄T�����\��#3�;��=\��u�W�=(�d�q:
^7ܑ�r�Ʉ����(3�/y_��ޓ��faZ����;����t7�Z������gգٕ)qBd�2�I�k� q݅�j�j�vuM�OO:BU�ڲJ�j٘ӵ�-��M��r9���:�ʜѝ�Q���C�G<P�І�ϯ���r�MCrٚ�m�p�զFN�Ӝ�=�{��*U����]_���G��w+�P/��ep���K��:�Վ\��Y<�LR�Q�L���F1�{������=���}6b1DS��6,]�1.�R,����U�Lo�҄�*������o����zD����|��)
�9}x���e��vԞ+��w��1��2o��.����25K
vD��)
0���"^�z��s~A���X)J�f��K��b.2٤�ntcv���*��X�> Ж$��*c�Ņ�e��Q'�Bj.���xrt�K铲�w�ڂ��ch�,���
�1�|�n!`U�&�T&�SR�dx��Ű���$`�<��\�K�Wu���kE5�!8��g�V}`.��>:*aY��ǖcï� =�Y�הwA��6'�E�W��:/��-y,���S��lN6(0�s
xl���]0�Ǜ&���d��L���º.-R�˭��E�ޝ^��<�"�z���Q�ǘ����dz���tfg���T������u�@,+�j-��)��f��+w�k�4}��#*���t�kƴ�FJլ�f_(���I!�����?�]G��ѽ�w�W	�S!--��)�.����SQ��(>�W�vp�b�i�R��IIgQ=v9��u�KE~����4BG���k��Y?V�eU����pa��/�d?���gMVǃ-�A�r|��F�f�˫�`t�o��bK�N{�\�ޜ٦h\��Hد�KS������S����O�]�v���v�I�����B�;AV�8�j�΋f�5�Nl��)͟L���®��QU.)��soۧ�es��a�����	4Ñ���nt6�#�[X�v��}�K��ٞ�G��8�{�2�����'E�����LH��T��,1g֌��V��/@f�CϛX�c~��1��z]�u7��Y��53��>~��PU�-W���dC�+�����d����U�S��#{�(QU!���Y~Q�G�@Q�t���z�V����P���D�S���Z�8����Lx�]յ�>�����4�5��rʚ�y�nz�ɍ�"����g~9�y����g]��]2uY��~�c���zN U8��; U�1@�D��@�f�K�W��1�mg�Oi�ӴǮ|�e����z>�#mʏ5K&�;��Yw���I��6� #�-�T%����**���W�q��T�Mf��{�O�ȑ� �yȭ%N�/��@���5a���
_����)�^{�5(59�����Oӈ�����+T"�8rݐ�إ�׀��ӫ.�T;�}�Rn�{vH���$���.�GU��Y fV-J���������$:^II-eӼk&�y �6�'ڭ�,vg�s����t�/�-�o�Eo������-��'-���U�R�4��U�UbX����B���l�IF�V�#�W��+i@T���'�u�� �s:����D�͡�0g�JZ��H�9�4�I"��&ڷǖu-���h"NU���ܒ�5kc]�!B	եgm7������d�qbeHSKq ����+
�VκT85�xh��/	o+v�Rサ78[Fl�wxDb�<�`�ܙ�3|����R�d:R�mJ���U:[��)g�VL�$i��sk�a��_vDV«j���e��))����2���B]�8��WQ_V���8�ktz�T�\��+pI��e@*�4�f�:�v�_*9ɠnm�����.�ԯX��O��b���� va��CϷy]#��@歇�昚S�gw�|�{j�f�5�;�	�|v�]#C���*�S3~�qG�/M��^�i��wOc�`��]�vz1���J�V�
��W����.|�%�r�i�����b33F�!@=hLB������rIp���Hi{B�3:�bLR��h�H�B�U�2SGF��d[Y=z�y�Z���Oe5e1�������mQ[YY�������3v�u,�M]D*TX��`7�y޺}n��n��۩��l����J��t^ts��,6�I�\��懀��&�V��)]-X+���1��h];!�{�9�f�`�o-������6F�/K;�Y���XA;���Tj9�8���c\��^�{�FST(]�JoݙR	MhԸ��fN�C�]�K���h�q���j�e:.}��:T{]*�$<�;��<�N�����3�wU���=A2�wVw����V��r�!{:'�\��t���-�E۸�V�;�p�8����<ۃ�P\���*�G2��L��Xg+���ݘ�Wm0��ܮժ�M.;��
]��rǑ�|�]��Z��Do���YcS�u�q\.AA[c6�PB�l1I�{�M�o�c�\���I�Eq(�__S�E�b:y.�Su1��eg�K��7ylϯ#�WܴT��a�II\V+!4b����]�+4qܾ�]��l5�����Җ<S9�7���\w���v��{�d����p�y;&ٍ�wo#���L��+�=Х3��iպ��/;��2m�6=�-�x��i������t	۶Zb�t�]pZ�[X�9ۓf��ʄ���]wH[��8L�L���;Χ	���ޠ_'�o�`�7G���D��4�0*�P<�8Oￊ�
>��˵3,�0#W9_��4��~o�����qd�Z���DV!�cD��ܴe����{��xQQ%�����Ԛ3�W(���&DR�`/������FJJ�nh�Dk�+�zv�QX"ޛ��Ō\��"���u���t�|5�"5��7Hъ���bO;��cˮ��F�/O"�M�J񻮊+s��Th��r�Ȉ[��oR%�s$�z�����įa�끼rK�t�P��t�L���Z�.����^�\���ۚ6B5��o�D�w\��]ݯ&�$�au���\��z���.h�%nrTE%.cu���ε��^,]���x��/J�.Tkr�`�T�<���*����+�ͺ߆�b��k���q"$滩����b�m���JͰL����l`Aז�@N����n�J�U}[Ԍs�}��wP�K��ʅ<yX��aMt>��}}Jo�|��O�
�>��K݌�ω�#�ٽ�<(z�Uu,#�e=G�px�qv7!8UpN,2�ڏS�6���j�ա�w�� ɇ��dW��`P"LLx)Q5/ew��:߉�Wxۋ-޹�V��l�ں�y�f��1Ԧ*�94�ݪW�}\]�鮙+�Q�mZ�^r���;+�����'v��uy��R�M�d�7�c�CZ�鏶z5�Q�٥�u������@.���:���F`�TNoV�}$W�_��5Y�ϼ�1!zX�	�!5}�{�a�lK�rgB���˛����r<�ںïK�=;]���ef�|�0����s�?P�x�ΉRvv<=��*���޷wm����q�o��uc��OO�����_=���!��!���(F=�@�~�o�\c߰fә)�cԓ���Y�p�KGʹy�r�5�z����~�
�ܺ�*V��n�ډ�2*z��<Ĥn�7�,V�<7����ږĉ�B�B;UT]gs�ڽn]����b��-��V+oy5w�㐞��f@v��2�u���Wi�kW��F�R�m�I*|�	;��#��jW��8L��˷���cN���u��=n��E{�,+��\����n	���җa��MV�+�h_wyt|�1e�8o~��6+�>�!��9�47��r�V��ꜙ��@��A�+�b�'>9a15����qy�o8�︍��q���E�����{K�*<�P���F$��g�Hfo�z��U�9��j��wq�t"�X�Η�f�ſ.����?}�m��	څ�vTjf"��}=��ЩK����ǂ��	�SB�C3Fl�_vnZZ�S�f�;�y�-�������B^�r�*�$Q v;�ߐ���*�Ѓ �.X���ώX1Ǖ�eվ�T}%:Jv	*3l�ɉ����z{��{jԸ����V�@�+�:Le	󕃲�`�� �.o Y����S����v�u״}YD�	<�Ϙj�0�yp���p)��+3@�Bk��T�v��츆��ʞ����B��EG-��4��z�8ujcW0�q+��\+aa��*o��i�B�yN���ݗW0ý�מ'���9��O����Z��|M���t�-\Ņ¶�ɨ^����&�74�C��^�{�l{E��xWzE��{�fV��o�4�s��P�,)?'�cK>�;^��mU~�~ē���˞��������0!�u>�".]Ժ��(��YR,)��H��MF�7�Z����
LVt�*؏���wH`��r��\)�j��Yt2�"��7[�M���^����ޭOq-k�c	U/8��o�6�De���ۗ|ޑ�K��PsIV���������Q�(+�ʞɸ������ݼR�۶cV�e��A��䅱�ۃ}Nj�v��s�t��(�~���`^�eI鸝S�G�J�T�3���}�3�,[�|E�7];U����|;��k�/���qp���E�,~��<*��U��g_�B�1�ie�����t�c�����z8�ҕ���q��x7k׾���M>���40H}7R؟w�y�ĸʜ���os�q�9���Z"�X~y�5M�!M\7/�����|$hU�DnU9��=a�������ߨ�Q	�tt�YHB��b��u'�n\��fS�d<�90T����1G�z��>���b*\�1ZDz,S`�ۃ��H������\�nT,K32��+�<����'�T�{"�M}�Bz��_?�GD�=���◫/`(\�cvnO�n:�ӑV�tfhN�iN[�	�?P�NȚ=BE+�\�>��W��j2�"�Ș�u�ןs��l��BزY��6�%>�IN��7j0��[U�bI��Tة��'��W;�2����V�vf *�%�������ܕ��qT�]�)� �2�>+)���ꘘ쑀�m���7�����''Ƣ�����۔�ع&�t�ٔ�0��8]r������=�*�9�Pg}�Z&٢w2�oa�IG]���l��w��t���ﾁ��{���2��"���ĭx���4�{AW���*���q�0��B"A
���:Ɇ{���8�j�^<T�Q�R�ʅ'u�����:���'>*(.�Ug�
�Q�詄o�uB�����-�,X�@�'���w�k�z[&�z��a�lKbC��~��*�!����6�Ԟ>\D�?1�YR�5�!N.-R���nz�oN�m��	��N}~�*&����\���7����~�^���h�)��qvPzX7G���?YҊ��9�@�*�1e��`�99no���=D�'�G�Y߫`(�]�ef��Y^�겍`YGߋǏ�"3��,͑1����F���o+>��㴫b`֯�o�3�kޜ9��]O0������Է�K����y�B�O�>���v<�殰D�َ�L9�up��ͫ�z-�q�*��џ;����!}O@���s���S�K�pY+��]4�Z����V��ʪܽf�C��8�]�����ﮣ(z��Ո���p�յ+ ��EQ)����!��W�:�M�jX
��s��]��=��6حͥ9�anb���J�r�3�WFc6�C|�e��1�Y�����ab���5S�m�y�AS�@Ӻ�����,]j%//��A���+U�[[˜*�ie�����s�^m�
9�Bm��#u���-K�n��]q�2y����}��;�W�i-�hص���f|D2�D�x���&t���}=���(H����_Ypx��)ߗ;������b3,r(�9���V���v�eM����hؓb,E�Ϡ:1u(t�5��~��5�W�?4*��#X���5�]��S��3�9���Ss1��D���4�L���a>����[	��L{Oq�8��^�})���B��g�unTy�Y6����˸�`�٘��t_	t�*I�����ut.&0:��0�1���ʃ=�X5�έ�8�C��Q���ό`S�'�w�뇅��n��O���ۈj�E� A?VQ�W�^���џ��<w~�X(�˱�	«�ӊ���/�$'lJ}<�=��1��ʌ3�dP3Q4;Yex��k�v޺��_t����s��#N��2\�>�Ʈ����70�)S$B�;rA�٥�b�h1"��mʺnY��Y�-� ?�����#0�����Oz�RL�?�8�DVm���a����ltc���]B�tB��+(x�x1�e��߷�M�=��y�go���E)lH?/S���#�W��^�ϽCb\�3�;��8ܐy+���IF"�����x
}6�\6��gү���M#b.�@෧4�^d�=��(D �����TP;˔E�@:�*�����o�Y�ًAڀf��g-IsJ�D�2).�����p�Z�w����h�����8w�L���������@#���@��Tq>�
q�����&��r����Y���aɍ��8�B��͜�T}>�x���p?ތ��y	�7ۼE��}Z��W���V��h��c4�C���<$��:�r��`�\$J�UU�a9*"�x\�*U�<����Q��~����A�x�\�ܨ���bg����K�R[���p%�g�8������l��>��xo��a
�X�lH���zj!3`��41a�)N�և���0�<�j$8M�61�tX���eL{f�X#�(0�z&r{�}~�+^�+}E���(l��>^YQg�m�iW�ԿB�c���o�ɉ3�"}^�B�n�e��_���~?pc�f8G�/�U�V��pb���f/[3q�j�nm:P�������$��|��7�Viff�ܰE
Q�T��9���+VnJizFqO	�lô1�x������3z1v~�.tO�#$K����@��N|r��Ϗ,�V�A�&ٝ�[�����l{cS�:�S�[(�ac>
tL�T I�C&0
�+��w�(!6��>����O�����D�ٚ+�2�ڋu9G�\�U�,����*��X�.*�[u���*LI�`d���Pr��d8��/���W��[��vֵO$��|����aT�:����GJ�&*U����C!��*����:�'ٖ�\����|>#�����)�1�&�_�J��~	���<�Q����V�\�	��W�U�%�B<:^\uӎ'+�x�3\�+g�\B��ؠbUjc>*�JUS�l,��ؕ7�M��
��lY&���_i�
�,Tڕ����	ȁ^�ըMA!'��1W1.�����%�Q�ǯn��KD<���E���gpu�n׌�oú�NwSbj1z�R��c�K>�64>�LB#���zX�y��ՍY��J�`���R�>�Y�~,��f5oݙq��������؇�q���v�(^-t���vz���a2' �{@T�#�q`�z���|1\F��޷����uy���y<������a��wS�������`���߾�͚��ؘ�:�,9��>��إ�r\���J��yw!��8D��� �p�M[��8��nׯ}9�Ozi�}�����r�kVǞ^zw��^�V'$9�pB��>Y��vܿ|�����C��1P��|j��5����٭"�~�Jm�fQ�,x>�0z�6�W@jM����4���ϫ��ymK��k!��90h��O����gM��_l�5��H^����vJ(���R�N�!�hC
2�]ѥ��f]s�:�S��d�c�T�(We�F�d�H�7���PT�@ڛ6���K]���u��\Dɣ��v����rm#��C@{�t�{�^=���G���� �]��g|؋u��ȏMH��a�G���h�a��no�ԋ#S�S�j�rc�9�������yS"/��z�T��"�M�=��r��"�}}x����
0.]�k}U�f�M�3���{n�ĉ%��Ԍ�׸	������S�&�P�Ę~�k��H��z��.޴r'o�����.J�
��y���	}$'IN����F?m�D_�R�#4&�QS�ĺ�Q�c��򊛆=u�u*�E[�@sG'�����*��.ۈJpD�R"6�ÇK��zG��U�!-��3���&����GX>�����!=��U�X\+!AW�Z3��eզƤq?�|k��F ��ת�¿V[�S�����V!{װK��lKbC5^�˱�{����$1�N���?]bQ��L^��0�X���x�>W�ב�
3�O<��
�s�Uu}q�5\C��lƌȜ��,���X鸚�Fu���G�,��q��݋����`�('���������y�̣�W[���F|�����8=9�O��5�����-Mn�o�g�B��2�f�Lu��o����w���}��)~����ÃO�	^U��]���m�p�to�\�{�����q���)gR"�5+����+�)U�'Ǘ�(2�	Y9D�mh�����N��P�O4�L�ę����9�q�����v\�~b�d��UU*�@�>���}�Y�I�Wp��!��8�yh��Y,[��U������3�p�����~=�!����J�I���
�싰�����;1�i�#up��ͫ�{mc�ڣ��%���?Geر_w���l����ؓ�JxW��q��8$չn}�/C62���:[hR��A�mz�1����v��k��z0
n��!g��az�4�z{�>�;�y����i5���9�&t�v0�˰�1�*���z�V����	B�v�"�{�����'���
��>u�?�Ҏ�Nq�j��S`�W�7QF��+��L:��nf:�n�⍸����V��Gr^Ed��\1�t��:�R�N����<�&`�D�����ٔ��Mت�^a��f#��+���pXV�Ѻ��F��V]�S��� 2����f����v+��|^�^�JA����P(!<��0e��T�����C�p)���Q�����1׏hvh~"x���xe��op>7G�}�*a�`G��@1N]OG���9��`��.��-U���F+�C�5{��U��;����6�f��6�����9�Mc!��{M�ߣ�j_-�A��A@�mח�x�g�sF��A�(j/�\70/�d7/�^y�����R��:������*���>�c��7w�-�9�uU�tF����__�տi[d�mW��__7�ߞ��/����y��~�0`���"�3Q5LW��WOҫ�t6���2R�41W,������=����Lű���`N�8�])�ki_��B�g�钽F�[V�}��n��7��U��<���`xg����2~Ȋϸ�S�����'ޓs�M�׳���7�B��b��-��L�&�zè�~��ᙷ��vVz3Λ1z���1�j��{����6%�h/�5ٓ�-��jU.f_��X"�́�]Ӱ�;{�Y���aɍ��8�B��l�D�k\)kݑ�"����p��gR�����坆��~4��V��o�9�B�o3�M1ӥ�9}^n3�o+��ʽ��}l�S�]�� �ݏ3�U�S��}_:W��]71�Qp>��8��\3_��߽��c�T�zSmeƺ19�o`X>��xo���'Ѣ��"�n:4ݿ1oތ������0Bn�?|�,p�������p�����>��r0P�
a��c�N�ʸ��Mw��}���й��X����TX>�nsJ�����b�#W`�w�F$����D��2K���ab��7��ufh�d���G'+�E�J��2�È`}�m��7�%���Z�+�N���ũ"+	�Ǐ�����^�kU�2p깳�Y��5wQ�w�0��R���kWɓ8�L���K�*�v�lpšf�rg
���򖄞��ۇE�@C�+��Ȟ��	�Ev�Q)�ז����D�v�M<S<�k�*��oEa�x}<��rim�Sщy�P�+YK��%@���PN��sh=�r�.��χ���!gqy�5+<vl�b��(�u�B�=�h���w-Q�ep:wFM��*�K��mj#��C�iP=H�[�'=66>.H4�����˦��UϺ���,�ډS�W�u�Tt�;N�QPΓ@�B�q��X���@���+��\��.�ڑ�Ed�h��U)�ڼK�YF.�2�2�L�+4��7=�v▚�5Yޤ鰰-�qY�1K���tNb�L�Ш#�2��/��Ξx����՜�ڋXR��am,���<蠷��3{R���n�䶵�pB^��xʍf)��ѵc�������r�t���ʂ��1������j7��,Ln�e���9���+6Ve>�͓A�r1��V�>C�#cB�Ϳ����V`�[z���;&)G8,ɑ8�;���S�76��`�-�|*0�[�MV�ˬe�W��][��S����(;��\��/h��ʖZ�:[w�hJ(`��X�Zj.��y�kxX��<��	��6�2��Q$_���V�6�/�\;�;
��mJV����uפ�����le.b����[���1���743�i^��$[S��(�V����oRg.}7t,ү��mb� 3�HKv)_A�n�Xu��=HVk���q�mi�GVR�ꭼ�xR��I�8/��������j���6�/&f��e;�����okP��w���9�n�R왗W�>w��^H�b���eT�(󓦇ԩ��&�Gb{�+�<\��E]PJJ�j{��q.Փ_L�����M˼�,��>����dC&w�]�Y�ĸ��͋9qBo������..:�,��kHfJc^q̢wT���m;�����vsd�S�:���Ŷ.D��}�T5�pr�%�����ƯO@�D��%+�u�(Mͥ�t�Մi���ŻD,F.����C��s�-�n�+<)J�����jf�u���B,x�"�����v:4�*���Q�/��,z��"x�mi��f]ɰ�������>օ��AU�U��f*���k�Lb��R��&RZ2�k.�������ҕ�ɨcv�c;�n=�g�85wg�b�^t�pcb1f�N�;��1LT��׍1暛���l�SFomq���JgּA���!���`���}�Z�n��g
Y���!g:�*�䀆��voY�98r+�p�i#�|���� ��S��*LK:Mbe[�r��p.�n�C��*������՝�y7��y-�],��;A|9E��zj��5����������y��;��o<�WM�r����Uͼᴽ�^�w���W5t�/K�zz�ܺ�H�˥�����k�\�=/]�5�)r�1sW1��<��u�
�3��E��׎QWǯ^z_�󷧋��SŹ^��/J�5���'r��,�y71W5�\��f��h7�RF9N�r�x�K����ux��:+��J��u�w^J�Ti�r�l^wc�u��9_r���^<G�x�4!n���ͼn��k��E�.lZ
��%��]4�b���d�wQI���Ws�zn��s"�s�ί	l���9\�>���y_����u��-a��Fտٹ�
&��k���AN��2K��[�eH��v�oa���Y���G�}U���ZM����������������7���_�$Cs�+�=��p-m>��9IM�FvT	��bχn
׊ث�����阇{S�a}�T4f̾7��U��
x�k4a�y{Ut��~��#������&:2D�`1=�	�1t8X�;,�:��
C=-^X��I�wU�(�ό��%;�MH�tY�&W�T I�D�:�X�>r���P��89�£�]� �P>w�����97�+���|p'�
1���*Ջ���T&�S��m���V�M�����N0;.#��7l.�(�Ujc>*�N��-p��*M�S��L�\:]/-������*�]��"{e������o�׉ȁ�N�4MD�!`�s�ұ��מN��c~Gs��ޫT֚N�R�Ɯy��9"�6/9{N��PB�0�=���ҷ�j�V��o� ��C���[R�h7�48R�^�E����/2�b@ve��A������k�Ml��/D[kpbJ�H�8�����?��
�/즿�S�'���[��x;&�9���m��n�5�!|x�k4����*)�Ω�w���W�G?���1;��D��OF������2��<X0g�c֥��^J�SUv{&��&�U����o"|0>�6����\򏭊ͬ�;=�K�V�u��5:�����+[^S���k��jB�A  }��o���3Z�=�-����8y����j��7@F�Ӟ�٨�ؘ�­�r-	�٧��⁨8��n���)��|�/*1�	,[��M[��'j�v��V�_0���~�������__�ҜbM�<e���}�.�p���	�n_�SW���k!������
c���z��S�yӛ�f{UzX�,*���T�3&�\E�x�s6}X��ߋ�j_��C�z{�;)XY��{�_�hze�'�Y*2dGMH��:��I��͇nZ�H������st3Xr�� i�NCt����Ar.D���O��pc�`���׊^����ES۞����/�{�k��s��w�p���ς��4z��b����J�9٨
1ȅ��O�T�z/��َ6�y�3䍳:��ntcv���|�`JT AD���&;���m7������.s�Aw�z�p�9�������Uٌv�B�Z"a�L�믯���������C��&��7Sn|g~�rs��}MI )��	¢��������T:U�ly�C;�+�.�r��j�#�3{�D�蓻'J߮M"�V�݅˰�Q���Y$¥�[q�}�}]���SK4V��/8E�!"7�:��Bm
���;������]F�w�i��1ʺ�?<��� @zVld2�����Ir����x]�_�m����Km[o���Ϟ�>��>L��f:?�*aXW3A
�X�>WB>�w�v�{���B����N5M�t�2)�:����Z��B��1<��z��ӵg�Z�G��LQ�����:�Տxќ��@G(�涠���Q;��OM�d���	����ڙc}z��B�֖
�\�x�dx���М���=N�Z�Խ�dg��}-���Ӹ�+��x��gɮ�9�s�ӛ4��ɟԋ���_������ӵ���Ŝ��ݕ�Y,[�ߊ�!�}�^9�f�>�DW�9��4���!z��hOF5dݾ�c��&�?z.�bt��0	4Ñ���s�6�!�V�&���CUa�v$,�3��l��6K��$�@�A�
�E�! �ќ�W�s�U�gs���2<������Z�.~��r�R����>��#�t��;;,�y���`/[�\��nd���l�=����w�O��S����ǂ�0o�W���W���
�b�����;fЅ���!�w�u�"�ϣ=/�n�-���.��~�a)�S`�xlϑ�&�W�+�����3O�0v���$)P
+����`:W	&Q�%�@;��1�3�dO@s�{k�3�%�eXó�f<���b��x�L|�"������g{^�Z�M�{S&�:�,�����gE[w;[xS�y:�sM��u�v��j�lU��̩�hO>�|��������V����&�ַ�������%��]��V��9W�px���y[SY����eǦr*ɘ3�0<N1O����g2|x�xJ��:��c������e����z7Q��G���k���#�*Z��|s#��ڝVx�5��F<�#�L
KSu1��*õ{	X5�έ�8��OL���o�by�WR�#Ċ��%��n��6{D�}����fO	15����F����G�x��bR�"D�**���Q�@��,3�'X��6\`S�dAu���������[h��Z�8K�twO��:X��E_E��w�c���E:S"��Z��٥�b�i��mZ���
׻��ze�������~�~���M��u��iL'[Af�2=��f�igXɝ�̝od��h��^5��ьk�º����ٛ<Ưc�lH��bc~�#W���1U޹�Y��Py�3��~(S�cg&h�����]wN�~���ef�2Ň]�Ü�.�b�q(�S�Nir�Η蜟l�?hۚ��B"~a��J\w��1��N��BMS�/��֮�L5;���/w�7XK����26f���RH�J�n�q����eD���0�N8��:eCE�`�h�Z�+�)�mP���1GS0��,�{��L��un�R	��7O8�S�"禛�Y׊psjHwpw]ݙ��a%�ׇ`a?�U}_~���� |> }�u���ka�gӅu�?�⁐������mKͯDՊQ�J�7]6�N��B��=Rs�>�|�y���1
T{��Un^��kט��ߨ���}[��}V�D�bD��hӍOw2�o�s�n�k��qE�����8���ߌ��8�X�7�b=�P4p��ȥ���j}
������:�:y]�H�g]�0}���{�B�b�b7�o��s_�(���z����^Dܿ�I���A�R�9�9X�o�=����f�fn5e76S��6� �Ν�[Έ�JB�P�@Y��f�?��*���S��yc*��7~)�]��W���:0�q�:�Q���b�aN�����Ȟ�,!=�OA�8F��r���7���6z|��B�FB�U�,�)�߭�R�F`�H*'�+�c���B|�'7�=�m��fw35�Z��p>n�_97�):��N�6hk�
tD�V.f�!P��H@�+�끋;�}}��*��j�!h��6�bBF�*�LS��+���r�46%M{�nN4����ȷ���/gw�o`�c �;sr���K��γ�R=t���m�Y�<É*����ڜ��ίV�o/U+f}�J�2���u�WaS����#��囙����g�k��Lt�]��Nٓ����0o3��y8������	�O�*[��c�iZf���b���j�:���@*/Ս��A6���P�"���mϠ`���5�ND
��P��M���N�e���P�I�v��4���o_�10Am^�C��@���J�uQ�Ox����>��;��5�0����8�k��6��f�^1�{��ck�.0�mJ3q:<)@�܋�{5K�f5of\lW�J��ϧ�u\��J��tD7�i;="}Ր"-�U��v��K�D��5�b4����W�����F�����\8ϥ!n=��|���>��n�o�9�͚��ؘ��U�o:j�����9m�/q��V'H�ӟQ'��`�Ÿ{�-:P/���nׯ}9�ޚs�M��u(�=�v��Ƴ3b�f5	�"���R �_�&�~M\7/�k!����0g�ylB��MS��_!�/.DnU,����GX�p�)�K��5��{fܨ�ڗ�cQG�=J���g�F�1Ϣ�Znc���� ��S�+b�u�R�`�aBϗnZ�H�T���*������|㤾�a�ޗt�3J��E�+�Q�)}ʨQ���R��럏��x;ߟ����-Y�53r�-lw�ߙ��r��U�p����\V��\�ç��:H�>�h�Y��]v���J�����*m7:�c���zFC���*Y���a��^���Y �����$�+!��I�t�[�-p6�	�;����}|^�}}yނ~���Mm�k[m��7�&&���fG�>���W(k�eހ�3����❑4z��Q��"���9�סϣT=�Ƽ\�;/ �1��t��9#l�r��ȕ�ڌ�qN@��bm8������w���1`K��6*c�Ł먎����Y�~w��8�s����Uٌ�v�B���f:��s��������D�\��GP�B�����vT9=�";�>����М����kjb/���*>�{)|���1������!@ϸO���ީ߯��-��B���u������,�}��?�T�� �RʋS�g������\M1J.,=J,e��sFs�{�eX��^N�W������>h�Eb���<	�]��7��s����_M��ç������k,TE��~<�/��O1y_N7~�[��^�!-��a�����Nl��c&|�4i��!S��/zߣ�z<x1�B9K_��"���egıN<U1
�y�4�uט����@V�y ��&�/����C��𫀼*�b|4��'��t�a�������7�O�h%�9Q=���Ȋu&������+��m���j��V&�^�뱀Dso�ǔ5�'#���o���|�L��c�&�f]�u˩p�����@Mx\8�Wlr�ͨ��qaBeа��{���c˓�9�g���\N��a��ïisdN����>>�~}~�U~��RV��z�����y���W�a��Ԗ��+����Wμ�6$��N�(!�Z3�jܷ0�h����Ι�����6�ӭ;k�q��|�1g/�*���׼�ٱ�O����9?GǴ��7�8�O.��,�>�*�r���ǟ>� � �yLz~��
��W�(S��&S�U�(��mu�_�y,ΧB5��{�urʂ4mù~�rZ�C���*l��R4'���]�ѕ�E��ے|xjP��#�]*�Ft��A�y���mMg��t:�N��}?N�ϕd�g���-(������No2�&}�~��%e�e��,d,
�z7~Fە����z1�т+��o��.�������dLc���ml�G��A��3�ԯ�ʃ=����][�p)��Ӓ�hb(b������c�'R�O|g�e��|j���jH�&&�LE�(�*z<�eC���Q��p=�.[z̾ROz0�-\��5p�8���c�6\`�N��@�D��Dy_��Z��}Y�Re�!��������p�3\�F���
o��^���N�w~�K�W<x[7��T��B���ݓ�?b��L2��z�;�I�.)�_#9�.��iU��8T������N�Fײ�왡f��_	8
f�]�5P�q۶]��".�֢u�����>G����)C��ye��-8�>Z;��Y��X�yZ�ָ0�����n�Ɉ�ʿ��;��V��}� }��  � �����@���K蚓ӿ�Y~��^�P��dE`�iLg�ߡ�-T��z5���G������roTia��cC��u,�jݍ�ϪKN�.��/z�z�bbc~�#W��ϒ��e\xk#ٸ����@t���W�_�c�^�u�n�������Vla4Ó��r��\���^���Y��������>��pc1�?0�m�R�FV)��}2�L�Ǖ�6�<\o���؏2#�[��/|�T��O ��x'Eh�}k_:_��?�`E�s���{���m~><�����nd�P�ꪷ-�c04�S��J���S�G�,1^�����/\���w�{��v�X��mp��� �>UP��p��h8OL��8+�7�pL�f������L<��twx� �<+b�x:���F��^wQ��m�h*���Ty��ˈf�425�2��1/�m�lO���>� 3;R���YX�o�=��c����7�m���2[�ɥo(����}G_�I���(�v#�ѣ�]
>2»nKгpjߕZ���aG�\�<��6�ds��dV�Y��J7W�*�unT�qGj�T��G�b�<�]/���MtY쏳yK�h9Q�}X̓]2��4h��V�*n� �[�!QH15��`��Qh-ᰜN��
�6*Dhotԡ��<�X������{�ǯ���}��{�����m�&�h��֥m�pg�}{�-�@��=gdMt� !=��1�PT��c���	��={�;��'�����I�gS��c~�MHgQ�e �@� ��"�u����<����=cם���^�o�^\A��� �.o���t�'sS���`k�"R�S8Td�����ֵ�����=V<��+�T�v�߽�\��A��{����at�J�ap���V�&�eɡݏrw����k���s<��+�n���u����@��P��6��b%��HR�!I��^�E�9������Z��Ɠ�R�Ɯy��9"�63��H���.8l΄8�앵R�U���Ϭ!�,�,m{%�u�,����D7#@��٪_nٍDX�$6����Q>��B����2�;��1>~��<FD��q��{u�+VD�.=��Ҍ\ԉ��3Ԝk��y���)L>�0��e��,S��+�=�to�8=9�Qc'bcg��߼�O��,�C�ܽ��ïP�	신��9�g��zK�5}/Bv�8���tW�},| !w9��<�M��GH�R����ڶe_��2vVa�q<��n���>�U�;/5oI����H��U���'-���#F�л�2�Q�\~E�����|��}�wt�K�`n�\ �`��5b@p�g��V�Y�W�00��n<%D!XA�2-լe�9G"�;M�9E-�
���'CO:���b�7�Z"�]u
��X:���y�[�\3q�l��p=���MyͰ�;Z3o�pWZt�i��̊fu��5���d��J�VU�u˅��2�'z	֑�؏h��˭Z��ÔzF�H@[���6��j53J���(@{k_$�R���}�ZN�����.@Q�w�D��A�f�wy�H���Wz�)�[(��؍�;q��K9�6�i�Ju�C��>i]��n��� �F�4���hn��u�,u�"ҐZ���)N��}O%�ɝw�Vkj��<��{���Р�8�븶��2<Y���7��ϕ#�}�$�{;��8�U��,��pחy&�v�;|K�V��n�on_ÐԜ.�
o�T�����	MB��$�N3t��ܺ(�h�٨�˸���*�� �V@MA1vWU�'k����)p
"�)5\�ͩDL���}R��K��SU����Qr�㱊�mV^��ݓ�t�L�k�5(���f��)�U�Pu\�gz-w$$v�}���郖.�r���ἇ�&FVҹEj9Q��pAR�D �\�Pf�sn�E�.G�{�(�p�fp�ˬ��\��0r=�`���1�
��gXrb��p�%��:q�!,�s{�^%�9ٱ\|q�*�]�s�n��X��N�4Z������WF���~PP���rC+iT��X�]��+T`Iǋ�
F]r��j���2�*#c��2�l5�:��cn���n`�wV���5T�t�l��FY9|���+Ε�[!��ڱJM���ޡz�p#�%xNwK��t�F
y
S�m�,�3��Cq%�o5�;oB�VrJY��9D��Y�5�����v[�$��wG/*'�hֆ Ĺ\�P��1�8'5t��b�%�Ċ���6C��Q�ԑ��a��
�H�+$Sf�"�*��K@����@�Y�w�{6�efA)ip�SS%����م�r��Y�g#)�����u�?X��id�\dG�b/��l�-�I���q�F=.-w1r��s�I�=qPt��ɰxN��25�Yy�`}]1�;�H�4�X��Ǌ�R��"��.�.��5]�XLP�w���ze�Z�B�O������U��n�����t��w)�K"�k�nf���˨LuƔ��P�$�f�a��?su�ko.R(j%��N�Tsz�yBL�%��7� û\��F5�Jk}� ˵N��e����.]a��l��2�Z�f�2Rx�m�ʎw7�\N�e]�������3]+�p��)mH��br����=Yk���zI��4ЦmPA�Mz�w�z�׫�JMW�r�p���(�4����9�M&��믻�����ĢMF�!�N�A��rኔ�鳽�{����65�r.c����J4[�4�i5��w��A�^3��u�����&ܹPX��\׍��c�O%��B��sEx�[��-�6�����E�^6�j�wnW7rܵ�܋b�*/K�E�^wF5&�킷wF.��F(���瓻����%���t���v�r���F�r�mG6�m�) ��Qbɍ˧;6KE��s-޼�Y�U�U���d�j�x��=t�CGx���	|�۷B��ۊ�Cq�T��W%�,�fbcY4�cy≮쳫o��m3�%��_?^�:s����+ZJ�k|}�������֜�;5��O�l@^����E�A�E,�g�M�r�������=뚪�lZ���8b}.�?��L��ۥ�\"b����T�38r���tM�t������.ak��ʟw���:��Y���!R�Q#�C�[��Q�V��[jǡb���t��~��[���%uH��a��8��r`���Rc�r$��+��qQ�Q�}K�o:n�=�]9��g���z��u��{F.]�w�+�].��	��<g쉠z��Ř��>��{����~��oǇ��H��X��Ә�a�w�6�NR��_cv��S��V(�MA��)잢�Íyz�G.~�#�$D�`В$�ژr����Gzpw��-
�8[�sG'�|U�}8Wf!d��c��C�sml�$bcAckDL;B!�"o�56M��N��P��u����jN����&�fc7K)x1�F��zwOAb����:ݥ�H�rd�Q�)m5�Smީ�}^�o�`�s�R��
W(����dYj��!)	"n��<6~�:�*O��u�Qq1�Qe��sp�<�{��Em�fB��M[�"�]����]���N��s�%�(����tUu��C�݄�fb�����w-�<�B�[�xVU؁�b�1�#��nH�5gc���+��7r4��
%}s#�8֝�ce��$.[udqT/k���r��f���r�������]W�WW���x=���$���g���p�<�"���p|��1�ڙ��s�7�Qc��k�b�>F��T��u;>��>��.�/��f�g��[�n�0so"��!����5�'=׮s�Nl�qk���!ǧG�-K�����$���9�b���O��Ct;+>%�q�[�Z�rm��	j`m�W�O�v*��\�����X`����xU�>�"�6'OPBu�Bi�"w�����\ө�]���z3����8]��pp����X��_��D��\)�b�����y5�r=댋���k�=�ê�/Y���V� �>�'յ/��PU�Sw�;,�dt����9�A��<H�
 cN�H��cs�U�S���0%^S�O��
�+`S�G��'$�����1��������7r��ׄ%�ȳ/���-z������Jx��y��lIK�=v,$�x�{Ώf�<@�6�:���WI�������y[SX5؁��p'D�V�=3�5��'!��ɮ�����n��i�7��b�"`~���WY�0䬳��,d%J�1nLj4rn�pA��"��xY�7ꪩ*�>��[d�����_��	}�pi�7���X{�n��}�d�7��
B�^ׅ���y��E!��«+���>�ƹ��.�¡�X��ʳ���;Wmb�nXa��`b=��lr��g7�Vn��Ɍ9�%Ӵ��_�}U_ʺ��G�}� I���A.ؽ���}wzrf ��!�0)�*lT�NgT��ni�4�?#�!͗�f��U]r�,�l��۬1�Om���b��jH�&'�4O�c�݃w����I�����?A��^�eH*\�N,3�ؼP���)�2LO	11��EujQ/�����,��ߏ�����]��8 ͮ�����1�;�qJg�`DW��S{5��\ɟu6�˺g��.��F2��X��?*�U�U!�>K��y�8}�z����Ldz1�W��+���ѕ�b)�M'��ɚ���v�@���j{3o�:<k=��6$g���(Ϩ7�b!����[�mgS]���6�Fu=�{��y��ӕ3���xW9�:�v�������M0�c�nIs9;g���p�[��r�T.|SLN�]=�ʗ� �CtM)q�����}'ј$�ڧ��ŵ��Ŏ�Ǧ\�B;өV9~jŵo�v�<VԽ�D�X�WΕ�i{�Z��ٗ~��n�w���Tf�7Ņ�Pc$ӆ�@UV��m`ס�'#t
7�.�μ�1_�+��?5+}M�M�]�Ԩʕ��.���>��5Y3�ZSnJ����z�0Vu�
��'=�����L�S���B*�Y*PP\ח�i�����7haږ�,7}�[� �Gj�r�\ʋ�
Xfj�̱vJ�9�r����K१��-2/;��SB �U1�<��Wx`N?T����HA�7�H>���v�0�P����~�����)�]��pa���;�7(����B�B�R�"�XAN�./<��}���U�Զ!P0\;-��3Y��}��	C�L�MY�uF$́"}Ćf�JL�X�+�����f�fn<��f���1�#��d�}n|�e@��b�}:$O���6*�����/Vn]l�5;�Tt�mJ�2|��zF���Y��<��pOA��;� B�r��AS�_y\G���W"�'O�|�F��x59��GS�a:K�ا-H!�c�V� ��#�Z��y87�'���ޔ�ˈ=�x�asvro:W�w1�	�C�±�"W-�z����p��Q����%��̱��X�Q�ST�V�츆e�&���ؠbUjc
��ӟ%w1,XN;8i��m�ۊ�^�b`3�2*��s4��v8W��M��{~��NDzup���億��������a��b�?�����+a`�f��P����+T��zے3+zv7ƟN��-����n���6��tB���*u�EL-;*��'Z�Ռ(�f�zh�t�t����լf�8��΄���\�K���Z���im�7��i�9���޾r�c�x�'�\��ʝco:��sZk&��y�;�"�F�î�8����lڝ�>*��V>����X�mo��ɪ����>~�}����_�����?���?>��~��4�迶�����K�Ʋ&��(�[�c��f�yn��3tΜ[�>�3����FC��a��!��XO�9����-W@1N:ɤ���w���}��%z������/E�\��x�?,�^����v/&����X�x���3ԍ?B���/��C�غ	�V}�,||��)�*jܽn���k�
��T}�ṡ��;�光�?�l7)_�G*�ux�C^ڳ����)^
j�B��jS<���ǲ �ˢ޵��#�wn���=,*���T�38R�tX����u5'|�j�Y�Mn���'۔B�OGSu�_��p��]����Ȏ��l:��I��Y��t\wB�~�=����~����ͩ�[�S�Uk�ʄ�6�L`r.D��G_܅3ġ�M?~��Y�wq���-߯,Ӡ���\�<#��'�s�k�eއ�	��g�S�&�=BE�x�Q�fA�NO����u�_P�>s�}y�㘣a�^���o�K�����t���29l�=_������У���e��	��)*:¾�$�D�byB��RU�(��֦+s(n��'环�f���$�+!BR�H�pD���y��(};{+�A0v��� �e-��&w�(m��n��=SoCg�p�cj�|�������~���>��>5�y3^�A�ww�X�<	BZ���q��Q��񽇿+x�8�s�*�����A��][�#8o��'n��쨄�5�&��DI
���Հ��8���&�j�ş�"�??@H5wsK��u]3_ޱ,?E�
���\+!F�������P+��"����ޖ�K�p��9y��|<w��fw��y��)KbHlPa�u
xl�c�����\M|�zTEtٍ��n���ǂ>���ye_<��Nz�p�	��z���]��7��z��ɨ�����V�=���C��%~b�Y[~	�Y��������ȃ���p1���k�'�g����W�x�%����_���:�L�6(h��ǯ���[΀ގ�ϬŸ⩈.u��5L-|�V�uJWK�����b�hϾ���xM@~A�'OXCyጓL9�8n�˼}^�	��a��K3ym�q�*� >9�����X��@�A�
��*�&�Jr��RDP�m�F��=�7<��)�>2ª�/C62|���Y��ږO�J� ,5�07B�;Pe��wM��(n"^|����f��YT�~�:�m��I�{�����Yw
�{�V������8ݥ�to��[j�M��8�C�A��.]H 9ݎ�Vʹ������zu-��Wr�J�=�fY�0<����PX�%Dd�<�-�H�:�ç׽?� 1 }��|>�[��<[��:���\@kԪG�ǍπUX�?A�� }��	W��Ӄ��� @��A�(:�9ӽL��оs½�6D�nq��U�^��
�r_��Js��p5y�=����X"�w���6��slM�`{��=�KE�5p��ͼ������ښ�f�����A��Rwy{[�0�R�.k���s0|I���P��h"�ur�?�I3u0䬳��Yc!*a�x5~r��߭Ӯ��m���N1lq�&":`�q����i�n�Q�^��2�����eA��y`ז胂��1�z�w��"�P��Q����Xc��?X8*`���LM!N_�=R�ѳ�wlV���f�k�*wڬQa�7!k�y��ņS�Q��.1N��bbxI��(��؉��ޞ������Y�Ad؃$.���޹�N�_�ҙ��7�K�m�]\=ۨ���cfh@��*�f�c�Q������4��	ߡ����uu�^�_�BJW�3s��"q�U�e{U2|�@�u����fm��G�g��6:�_��~��_�u������\y�&�r�Zh�(�t�����e"�,T!��7��]����J�u]�;r��ݏ�۪"[s\�|�zV�=
�f5sQ�Y�ҝ��d�Y��9*n={��C+6��՘��kj�֬�Z�3��+,���3�-\h	�
��YҸ�7��g�؏��}~���C�S�H����u�f����^���Á�����"�����)��Z}5D9��9т�*>�FemJ͡,:z*Ը�sja�W���b�`�Z����e����)��ϥR�:�r�Ջj�(�hΊ�����ҥ>�is��,7�y���c+�O|�*��O��p����ߕU�{�k�19�o`Z]~�~��t�0^��u9�{���k1��
ؘ�$mu��B,+���<p�Hp�lc�ʰ��B���&�{U�y��Hɗ�/�l���
!^�,99��)����^wQ�e�8Ud5.�3+���q�E	�P����������w9�ĸ,H�E1!��� ��5�V�����~]�,R��ׂb_�*>���g���G%�p�;|���P�5�P/��b(T�o���.�N��k�룊�t�ϫ3ǐ��0�«}#Sv�!�هv�8��&vD�hOA�:3�2c$y��G�ϕxK�>�	���׿:���6��N���rԂ�fe�JDo�ǽ�U���k���|ukW٥�eLάR��k����\Cd������>���S��V�0�;ڳP[E5ǁ���&�����m
T�e��v�q��4,^�r=��K'h_i8_.kQ�m����.���w3Ĕ�� �R��y��3G2�;��W����꺿��ɮ�x/6f��#�c����<��e�|��87a'&�x�c|�\(fF���]7�����h����Ս�Zi���Q�G¥����d`{�׼����)�1�\��}�W�&<�]�X%��_��1�V�Ρ�&��Tΰ�]�^D��p�{��s�2�۽��k��W��z�b_:E��*1�^�>��:۠2�j�Q�5�5�Ꟊ�n�=j�U-Y�IV]_���~"w�z_��5�^����Y�X��K��j^�VR�)U���f�j��8y�G��̙��/�t��j5u�FG��a��!���1o��2'8�����*WMĸ�n�Z���sY��M/h~��*��8�Cz/���)��*Ç�?,�~x{y*�J핞��Be����~�(g�VW���Z�Rs�"ϝ���X�B��'[���#��{&Z��~U{K�!�+�<��\w
�eY�]
���z�O�A8}�|��������X��,�x�y�_���B�f;$�u�p6��̣tdF�S�}�z+�+������8r���.���T9j��[����g|v��� �g<�~�e	�56�]�g�� �]Z����'�!��/��N�_<�� cu��W��idG9޸����"#�wZ���uY7��$����� Z��Mv���lΔ{�Õhɰ�w!N�V��}_�
������s��$�z��O��X��o��/�d?3s��d��Ӳ'"�a�G��N;��"�P���]���Φ*5����u��g����r`��B�mT���\��z����;�r���0L���8k�Ã�P��(î��������3�I�����o,$?P�ʅ;"i26x�U�/x{����bC)@�����Uu\s�sl=�΁�4m�NR��_cv�U蝳�y�9p$�Y���&1�s������4�7�Lt��LGz}�x����p�9��ǅ����9��z���k�}�n!b�0���!P��MM�S}>S��Ou���v�5^���ƽ��Ŗ�S��}hN`*���n0���b�>R&�j��˔n�<�s}��T|�'��ܰC����?T�j��8�ņ�P�՟���e`L^��1��Z��b��ݢ1���	^��JN�j��R6���Ȋ��p|��1��S"wՎLVMFL��|�n7z�ʿv�0�%������f�߶W�/�3�7{9��W[���!�o�L��Ϸz��T���2�A<���ǩ�1�Sv���.�չ}QZ��0)��a3�!7p�q�uf@�G�a��Z(��9��<f�Dɋ�lY���8L8R��c���	���ki��Q�r��v�ԙ�J|�sm�oh���N�;74�;b�*�-e���T̖8dPT��3p}��4\�!��j�f�f�&�YK3��gb��K�C���j`5%4,)憬o>Y�y�3($N��<�J��[�����qYY��}�Dp��f^�u2�0Vo<k
��k]�/c*ԁ�ֺ�ʻ��B�^fd��9Tۣ(���Ò�y�%��7�ꗵ5��Yl�.����(ݓ;C��N�s��V�G�W\2Bs���G3)-7Y5�ˏ5Ku-sM�]v��ӍU���j�f`+{�oR���^�]��%tZ����y.X�'�;۹����#���1�u0���B�K�:�c��uט�՚�H�Jp��c8{1���@���F�Z�f{����f�k�,w�����������`�?)V��X�S'Z���`��@H�j�Fm��츢X_�Z�=x�륗V���;�X������k\���%U�R��wZ�͐����Fm� ʙl�᧦#�0�fQs.Z��;��Wy�z)z�`�l�'mu�x6��p=��ݼ�d*�I���&DmE	��q���]�2��R�3�������PS�k�h�ܻ���f�E��9��ʶ~�ō{�^ч����S�=��.��N�7J���Lu\�V�8�#��w.���+F�Z�;�F�D�2r�ڛ�P��љj]hş\� �g��
�/8`x�n�K�9פs܍�r���(bӽ]B/���Y��9*5	��3�L���Li%fWTz����X3��n4�/�wY��=6�`��60Ùm�1��+�R���F�p�ΙFNAZ����]����<ݮ����s.�^�%),=Gn�p�grv�u��m�:Ws�����9��G����S	�Ojn�}L��&��CƂ;j`��`��vs�;��O#��4T��:��>c%�UjMc]&�B�����&Z�j����xQ�Q��+�ne���K�V�@)�w�Z��D�tMYł2�V뷮�΃ζ�������
�s��'	9���R`�N�=�N̋��;�7��+Y���e��Raf�J�Tb�*D��/��
ۭ��ίav�
T�c�.��Kp�\[�擲�uݡ�d���LK��Z���Ce)J�l�T�Y��7�$�C�9a㩇J�
��m.�䲸��@����q�R�z�և>���K��Jxۖ�X(i a�bhW��ǘh5�6��#�6��z���$c�7�^D�8��k����4�ZR,�'z��l*���a�\�9��2,&	R,�+!��k�fu�p𥖯�z�U�i�
KoV�.�\��a��a���f8��|��s..r�u#����7���ߏ���������ܭ�lmr)J@H�^.T�ѷ,d�z�/����^Ѯ�h
5��b1Esk���)��yy{�ޯw�k�V4a�E(�]�#`��V-�mrK����bo}��4m%��p��(6��Ț��!DF�6�wW5�t���W5�J��6�9�X��V�l̔[ƹ��lW5�"TZ,m%�cWMs�x�W��#]6���r帗7#s;�sr7���ƍcE�]�i8QIk�wh�QZ捱�B&(6���dwn�ۼ��G�j1�Q���nQwh��刷wu�p��z�����Ē���:ٮ�[V��M1�ڀ#\��I�Xd[�i�{֯��)�W�r�ͮ�P�����n�Ԥ%w.��_W�}� }��<�{��vg��l�ưl���G��<�}~���w�]��X�n;@*؇C��Z����r^Զg���U��7g�e���8J�yV?����lN}��!��#R"�]O�sC�^W5�j�9ζ�!�6d��x�Ĺ���N�/%~ fPk¼d�%�����x��r�`*��%U�n|U�z͌����64Q���>��xk頪#cw�P�?z�j;^���-��X�Y�����n�Y8��UX�?�<}��J��'���nG�.���|�7���N�#��0xW�<+���^�9ߗ|����ж��~��*l�o�2Lƭ������^P�p*}!TF/���fM�\<1�<���t:O�g,�����}�'������l0i0v�@�3]�4�L�L9*���N��
����s�jk!�Zԝ�* ��a�˵�{����q�ճ1c�J`RT�Lt�9�ʃ=�%�f6ǲ�-���"p��u[�TOC��F�ö�(����Dr��F���}G���%�{��@��ҁ�k�͚J��q�^��S$������6kl����b�*��t,ұ+��Gz6�{���ŷ+~��vl(2�pk�3:�oa<U�=�|�v���hYww)��ƫk)���3�����%oQo�>�hsoU>��^2��o�z|?�G�#���XX�:󨻟�ʎ��K��\��Bqa���s�V|?	D��@�A��� ���g2����X]|�VŁW^�����CD؃%w�8�޹�	�Ë��S!p�SI��~�M{�r�ֳ���_�V钶�!��_�t��9~��^&���jȊ�IL�C����n�g�1�.���z�G��~2��+ҫ]BVW�M��X)5nǿ�KC��F:lH�~:Rˏ^��m�C麗]D\1�քg�+�O��}�����Шzǅ76:�v�g`m�@fp_�y�Ow�y
�k���u`Ʌ�%�(?P�|47Y�*N�Ǩ{/jW�Dy�CoEZ�T�Y:�=�~z��t�\�L�~8a�
�#8$��:�r��5��o�����ڗ�^��SQQ���g�G��m�vE���ş[��N�
�ܽ�6�kwi��(���A�G�??nF������*g����޿G�a
�X�hH�!��7�Y����M	��nN��f����蚋d=3L'F�NL�f�_Pa��L 䟁�)��./<����ۜ���[�b��$���Tc����ZW*<ܖUeaV� f��|�V�[�J�RmL�����(��lk�zuДá��Ң��$J�o)��ӯT�lCB�XƮ�M�/�8� �l]���}ӛ�/o�`�X��H�8d����}r����Wb �;\�S	ƚy����@�����7�o>�1&nD�(1!��� �Ϭ�9Z�pb��r�7H��y�J�z��ǝ�7�m���BA�ʁ9����>�'��\�
�,��k�з����#mޯq��?\�����UZ�S�f�;߱�1"#lOG�쉠:D���x��@��G�v�~�+ǃ�t:� ��V1��[�)6��t��o��5#�r���=PĎ��Z���<4��e����/�=J,
ܬ�v\A��� ���'W�-;�ß��D�V߷t͸��s10��.�X����.���N�.!�z	��aw�@ϒ�S�{�N5l��\�*:sOBNb�⪘}¶��²�����+T�M�����%�Ȁ��Lk�r��v3=�ϢȲ�Ls��N7A��Z���l35�P�:�D�B�1Z�_�~�7.�=E;ׅ�ᕇ	J"�p�9��C�ƗN�LMF�aN'�cK>��\�59R������J���}�3�������3^�+�#�t3lƾ�����>�<��x�-O�3yا����Ҏ�����d@��k��ٌ�r�E>� g��>���{�U��j+X�@M����u��j��žz�������J��>�cH�*n]�ԷEz������TO7)���ͧ�ϭ����X�3$���T�\|��$P��B�Ș=Oc��*�~�N��N�LO�4VG��]tz�R��w���e��,S�*��ߖP�r���q7�e9.����O�
@G��yXuƭ����7�u�B�Ÿ{�SV�xI��])��{}4�ʞw�'��׾3�;�xʫ8J�F���z�e��xϻ,�gݞ"(�O�|�g���j�~�Y mc��kL��wn����
�=uN3�)^]^UU,gŭ��ޞ#v���SkՊ\�/�A���n`�J�CJ4`^� 0;�O����g0�TF>t�q���6���0�pbлL���y��8�A҅��U&1ȹG�O~�O����'�e����VmP����h������W�b���'��5�2�~{��#_X�9�'/E�B���I��!��&�"C`+��D���ב�~9�6���@ƍ�:��n]w�>��{�Q0��9���yZ��_]Dl	F��	bJ���:\_��;ӝ�{U�p��tEp�"Y����er�,����}8����qh��j�D��
��
jn����Y='���S�N��f�&�$��A��邅L��Z�ל2cK7�\R<Ί��]˧Z�Q �2���u���M��N�>9Z�� T��I��K2����$w�7���FM��Yy�VL��+j!�3�_l��X�o){=3���Ԁ������'��b ����_�~�'����>��VB�EL+5s4��p�R��V�B�`��k
�=��%�W����K�=��T؜	���?�՟�jQ�}��� �ڼ1W�\��H��!����7+!9�f��W��b���Ȋ��@M�8�L���׮d�V,�ԑU�NW��Њu�P�M���+�qd:q���J������'��� ��b|�~���o���L���׽�P��(;�G�8��Ve~�ϨZ/h��}���_�F�΀��V}a-�y�ܶ}�]�R�B�@�z"��j�m_�`f����^��%T����m&*�|�z����{�4a~��=�]{�.���\7:j��kn����g�v%�F�谨y�)�����5U��;��u�9\�?�E�/��1�5n_��*�r��ld<���66���}>��f~�L���0}w������I�����\G+�!w��`/[�N<n|���~��x��yNy�P�>��ץWV3>�����m�`W��1*:���ެ�R�\���q�pZ�v����qy)�����TG�\�kƙ�ܴem,�z�]�r�ܖ]�E�u�DvWWSˑ�7uh`ޟ=��xg�tϷ7S�ğ������A�{ !�?�t��������k�&��-��#��jrΡ��9�M�ˬ
Z����p�s����_�/�������`��y�bM���F,T���a�7�pO��bV���+��q��&�Ñ� �H���78�d53�D��:��	�0䬳��Yc!}}m�y��W���z��nY�ѾT��g�/B������4�@��l�>�·�O��T�KS�C���t%܈�ݬ�ڑ^qs�K��][�TOC�����j��~Δ���P;G��ڷ��~�+�Zȿ�����*J�s�*���D���-ʼ��8���`rFˌ
t@��y�ѱ:I����y��=N���.�b��4���X�'ޞ4S��s˖�H�OnK��湯y]V��y���e��{4�P��H��cj��p���d�M�_{�<�#7�6���Ds�:\{�W�aM�y!�n�/g�T���~c&hx%Mש`�M[��Ÿ�}�������Ed矕��b�DH5\!�{LG��'2���j����	W\�R��ַM��w��z��u�}��_��<�o!�H91�u1����6s�p*>�FemJ��a��beRk��+'.�ks���O��`SgDv�a��}"y���1z�q��HYX�s�ٍ����q,���1���sV3�³Y]±]���ɫx+%�:9���t�A�N�rF�q��mR���W�m+�H�+�
[x�)��"�O���:���z�;���v5�.3"�7�l�>��
�#EM��+�1��L�c���ܧ�c߭⁑����G�)��wJ�CN���~����0}ﶝ�h�.c�z�>�8I��7*f��͌O瘜�ڍ����a�ǜu�2��lR��>�D�6��"��y���B�Tx�x��M	�R��Zf�R��̙����:������7�pL�f�_P��E�Z)'~̰���\<^yQ2������nV���(�:���k#���*f|�X���1$���M�	��X�<{jlyݙ�����Eo��y��0�fn3�[m��N�)Z�ʁ虛���A[��\}���3Ӎ�����I>7�*,�zo�7��V���H�)⁚͘w��Xw�`3�'�@��k����0��	y^��.�!�lpj�xt���v}�k߀uo��6����S��[��g��}+���Y�=�^�!����4O�tb�O�����(&��z��9<;�D=+=B��5	�?K"7����gDJ��\�
D��N}5]�w�q�&�	w�@_eaB�&�y{��j�8e���	�0t���+<�;2KNL]��������޹���@�����VӍ��6�>��2��r<)��}�A�l{����w-�����ܜ�vSr��ɟ�#o��ca�{�^X�+�@l��v��պ�<01�����;��|0����"��A��>J�b�
�FFD���72\'�xT۟@���5�4^d�j�v��;����MA�)�Bj�-p����f�gP����E�+T�[�G����G�߭�,��ǽ,��;�K�>�ؚ�^������Ϣ������K�'7j߈���C����=��4O)���=y]�{2�ш��^T�<ۃ��Ȝ�{Mk��e�5ؓ���͵�>�)q�ǵ>������
�������}��\Ϥ�n<U|��c��6e.�zFp�w�J�2���³�/�u�a�ÁHN�����9�g��L�)���(.�^T�;ʝ���Y��ӌ'j�����]��xf�¼g�g	N�{�Gޣ신��>�g��(M�v�n+�����־*�zK
j�~k!��X�T��5�^:4e:����^�'�ma��m��]��Ѝ}�b�����V9p4�ԿA���g& �d��ӢX��sbviS�퍧��>�f���!C�����j��-�v:������\���(S��#�x�4w�⦎�R\��o�"'�U����iռܠV\�(�	�M7b^+7��9�K��:�w_l�����}���w>
�ԅ<�H��VB�̭���=���X���wE�6>�Ӟ�$%4���q�ܜҡ�{������3;پ�~<��N+f��:�Bo�
�h@��D�=���B���{�I�ϵ��e���2���b*�}�׉ȘC}/흑>�A`/��~�/���ב�Nb����t��l��t
ڧ6���cx�:�S�/:�X[��k`I�bI��T�GK���Gzs�oa��n��gU��-MY�zFd���s��W���*�� �n!b�0��B"A
��Å?X��𫬏�p}����3��mzғ�)��	�TP]��ϯ�²0�j�X����X��{ǁ����
�Cjӝ��%��B�ݞ��p5M���K*p��z�*O?P��fy^~���������K��_���l:,������1c��"+�@Ym�C{��̉�P��x_��}lY�g{VG�UYvP���t�0��yx8���%�fs�7{ͼ�+��f���ʮ��~�����T�<��F���|?}Ho��c&| lf�jlW�ao:{�Y�0�:�̩���Q�=^�$>�?��!М��y׆3}�zp�٥;��a����W�]�Ĳ#0@zB���ueg��N��p|\C�UÏ1�шY�z:]d9�L����Y����䰻��GIy�s��e)z����������OS�����ɵkW[�#t�P�t�8mbY��
t��N�$fFr��M� K��ݮ�2L%�ޥ9|*em���E=f+��w��%+Q�U �aupٿ{+���~��v�a�8�>.%}N�*��邮}Ty�dή�.�W1���@z�8Z3�M[���U[����xX�cEY��VԴ}�*b�N�ͯ\=J����Cx?����Eם�,9hC��/[�۶�Lے�P��}�&����\�U��/Ud�nv/"�Vܹ��}p+`Pa
���N;>�� �={�B�u6\s�*��~��좖n��ٕ:BU�E�%�jl,�+�hؓbz��X�@ȱ]WΜ��:y፼�qi���x:;�r�2�M7�:N|�9�L���c�D��:��	������Y��9)J���Y�V����	�aF���LjV����l����n�$�(?Q�W�=�)[�H�P����:�2�*����][�p5��to�:-V���O�
�7�$J1�d;����~�|;ϔ�}خ�*z<�aOw��Eu�!'*�N(>Nl*��L.̏Z^So6���֔F�!����
11H:qut�+E�����f�x�����U0c��_���~��b��[5���ھA�xM�jYͼ�]c5ً�̱�u��C���Ԃ.�v�� mm���P=�i���I�רd3�/�s�X'W-���3'NkV����${���Sy �l���J��m3�P��G)ݞ�+v�1(3U��Lg\�[b)���J8@���B�]����5>���F��hM�N�(0�&�Tn�G�/�]�T=eNʵ"�2�4��mı���Hށ�Ԩ��+Vz���.Ҿ�u���Yֵ�QR��GOL��t��`A���n�W(�Oּ�k����׮�*�I2�[ݳ7t�w�Pu!1_%3PFRц�֪�"��0`�;�̲3GFӝ��1Eo@�'���y�VE�B��F��N���7v���/*�f7z4�#N�s��9"={@+�ھ?H��u���i��hl�l�����[��|�昭�;$Or��kZm�Ɉ��UfNa9CBɕ�_8͘;�i�u��V�����Z`9��i�%k��剢�e'�UC��F�?J��8��̽/��[���%˖C�|�<9�����NT�P�����3�s%k��m�.L{�|����Z�6�oQ:����ź�K��M��4{��-�X۴��H���'� h���>	��|�TO�w�Hڼ�(��V�f�ZK%p�LR�����]�jX��*ʁ�z��͓F����%�GD�u�D��]Qe��\���!��|�����]�W���8j>ɱ|v�u_K�vcfu�S�P:g:�Pp���nͼ|�9��vG݂�	��`B��Vn�Ӟ��.��h�2&s�\xBGz�
���k1T\ւ,l<�'G\Y�Iqn��n��ő"�n�	B�ڳ`Q�*.P�3.����#S�`��N��;2qS�V��Lwj���xv)6$��0�����.����noaڊX�Sζ��a�� ��Y�f!l�uʝ�L�����b�W����7���M�����]�ˉ�ݬhc�p��>���]Xm�Fa��#q��x.�n�T��k�v�VT�9"����u'k6��ʟ��Cݺ��5]�N�䜄B�.�sf��4�s�n*���Z�Cͯ�3���1�����r/��K��`Z1]	Z�9�]�}��r�U��왚3e��+��^��L�wJ���i��zV��ptX��S  �;Ί�Ǡ�h�dK�A׼fU��gN^[�U���e�5���Q�mN�P=ѿq�
Va���ЭOlNl�ǡ�ݲ���4�RD����i>y�.��kst��2�����ca�ľ��N��Ϳ��;c�Ґ.�f��owo(���!TW�_U�����q��繚E��<q��V�gT�G>���y�eC\�cb���T܆`͖,G[&d�|�dM��CӮ	��ҙ�/��%ңSyf�:�+ڱ���Jz,��qQޫ
�ԨH(Qx7ki>Rn�r�"�68�^��}w)�S���Y�>��z����=y痫ϟ���\�TG(�qݮͺE`1䥃����/���,]wQrH+����1G69��vr�-˻��"�r+9s/w����{��kE^wiδ��Rk����\��6���\�;��͹Q�����W�փy�i۹�utŻ��ԑ\��ݻ�����TZ�wk�úwQ��k�X�M��s�q��]:FY�A����\�������*�wv���sp�ҹ˕�r���r��9���[�wu��×-��2ss���˕�sD�p�[���]ݻ����U�ܣ����;QW��$Z]ѸW-��+�ד\�+��X���(�'��kr��;����;����wW�y�]ݻ��r��ܣ��wv����6�nG-�r�����wWO�ϝ����ה�0,��ɗWY��d��D�����,�*k��f���pAEˍ�.��&,$�wY�D��vD��2:������.Xb�Fsّ�':���ҕ��+�i[V�}�쮏�����̵qB��y���D�ڦj5hU\Cۘc���%s6z5� f�iu��T,�]����nn��_L���_i�y	�y�:DH��LB��،��O��}�����Шzǅ7>��J�z���;>¹NY{���Z;+60�aɍ]L9��B�o�<O�=��+5PdĪ�����<̻���캞��Oƺ}A���+��������=���(����m⁑�3��x^)��Ux��9��;��'��j�S�����0.O�~��qX>�0I�΅Un^������:�d�yg�>�}�k��5<�ا�b��~���躖ċ�!��qE��u۷�/n�3%26skw�x^a0�E�sc:p����)�l�=A�'ѠT�䛠����:}��w:3��Q�`|��_�sG���R�!}@Ǚ������fĉ��$3>8 �2���w��x��7�����מ�94}�E��l��j�noS�>k��[��� �g�87��K�??0L��+r�pw�+qe��q�Fr�TT,�F��(�7�F.Aó���V�_d����.'FV��������� F��6��<���痌���n��o���ľ4��i��H���NQ���{�t-l�;�b=�X}�?�����2���x?B�g�-�9J��.�U���
x�f�f���E:��tN6h����SEu�z�67�s��b;��@�
/��<,��`���'�&ٝ�:Jv7�tԇ�����{��C��Wx������}9$!_DKF/��+e�>�Pg˛��97�<�y����7ӵ���R��?e���lj�"W+3ABhp���v��e�7/I��V���$ɜO�H��d���:�1���]8��ŀ�V��hlL3�{(��`?��J��v=�\����9��=��Dzu��a!8��Xi]E�¬l���P��"'��\�{MVʱ���'��`���~��F}�eoNǌ�O�-��k���X$D���Ǎ�Թ�yLQ�s��{;Y�S�� ��H�_�����0�.=���*b?nZ�dM��5��3|z�����ˬ�&n%��<.�_޺f3��}��\�%�q�8vK�z�������c�7�����|�?�w,�갸l';)��"П`����!�b�a(}Y�v��t���e�w(���^��^��/��We�E[A��t��ơ]�<8�K�wXo9h�/Vt�¸ye>V�]�s�T���G}Ľ�-�.d�$3Bӛ�d��3���J�W����a_^>���[���������> V(����a���9Dץ�ä�gW^�pt����zg�ć�^؞�A3��r�����=�${v��o>���r���n_��Y>mp�&p��ۧ9�OE�1���7�f!�Ճy�-�P.�V���ً�{M���4�ԿGVC��r`�ʖJ���'�/+0߽/����,x>�0z�I��6%�b�|�H���U�L7<�iT�4�������-�����|�r�y(����H�p+�P'���
�8/���`(ϗ/`��'��5�2�k;آ����|�d�H�,;"OH���0�5�}'E��sӘ�a뷝'ƥ�B�z�����n����y�4��Όtb���v[M�b��A@��x�[��9v���m����z�<����j<��8[�9=�_IUF8.ۈX�0��B �"l}�N|��go�\n��W��O��9���I��B#��3�'�"P*(.�Ug�
�Q�P�jgS�"�b��K�٧���v�b{d]_�T��{��%����S�Sbq8�ņ�TXS�g����(����Tw���¶ճ��o������F�q�t�K)*`s����U6��1؁B���2i��.���R5kq�r���\b��]G��1���q�`t�r�j�SB�-]�"����2�f��X��|�3��}�i�iy(]�n_�߄�@ ���7^n#%�J�}�`��/�5p~�b�g�ʴv�y�l����c��l��{0�޹��D�̚>���ivPu��tx!��|�p�۹��z�c�w��&z~s��l0�����E���@Q�$���Ϣ�i�3�64CS>����y��#>��g���z{y�R[�<��5���}��bkUni�l�4�u{�͚���>�a���U�~79"�o�]���F����Les��a��3�4Ñ�W��ڼ����2t���`������w���hX��W�Ouա��������E�,�ќM[���U[����m�q�h��x�|�P�؅��z����)�~�����B"�6.���ϻ,�y�q����d���L۔��lc�	؍��+x�����~�Y��8����0�}BP��]`w��)���,/S�r�H����Oۘ��vs�1��t��*lf�Z6$؁^��s���\i�L{��t��k4��ػ�X�����;�<�a�Jk��tL���<\�Wƽ�c��$��Ò��X�0Z�}墻3��*^F��1���u5�gP��Ze�ʓ�nf�:�i�z�i�V��� w��ptO�����p鑠�I�u�J9�a�&�>����2�ǋG!�vˣn�٬�+�h�,���!�폤7�����:�od<3b��֪�~�~�!4����G�ݗ�6���n�mʍj��ۯ�>YvJ�VH��(�G�3�5Xs+�^�nb=w�ǃ��Lt��eB����unQ=����#W�̬1�Oh��ウ�xO�v�Kq�uߑ51b}_^�*\x�vT9��X(�.��/*�ߓ��u�	s�����1��Ș� ɇ��dP��M(��J.���WP�m N3k�pV��c�P.�%�����#W�A�?��V�+�+���5�%z� �6�MKr��[�D������BH�'>�E�d�9�9��!��W1l�k� ���α�5���lO�h���jd!C��k2uz&s���y�/{���f��&$g���(ϛC���m_�p{���$F�~�@�T��M�q�㛿���^����^��Ӱ�X-}�Y��L90�Xr��\?���tNG����T�e��׼�a����zo1O���5X궓�Y[�cE��q��L�b�snS�X1���@�W�������y{�o�Pٕ�����X��� &Pk�"U^�8_����I�Ϊ�r҉B]��٢��;��G�q��B�B�o'j}M�OU͆���t��o���=h;���6�G�����3^��U�:��{ssz5�^ы4��o`��ͽU<͙J�&#��Q[$ޮ7Љ��-_�uمt�6�5K�ږ$���\��I%EOR���o`X>��y�G�,!^�-�:�y�����,���4��H{�ޛa��9�恆�͌r�Vo�pN
��@���(0�z,T���9a4��X̅��=�z�^�#6ظ�yQ��4��j_��@Ǚ������W���_�+�	�V��z�^�Nyon���=ƱЋ٭����pb]n��ٚ��V�si҄���b(���γ\�ͩ͡I���!�� c�[
�P�5�^���^
�zF��@��Э�y�-�����3=�2�q��ƺo��~�/�'�L+��1t8Y��; �X5���'�&ٝN����:[f!c�jȽ�jC�N�Q�Ή�`*��+�:�]	󕝗�<q@0��L�B�C��>�n��(��ό����	����#CT�
tD�
���!P��NL����Cr��a�+޺�/��7��A�Ң9�X�74�;�at��]�X\+a`46&�O�73A�B��¼�'3~n�]ݠ��޼/T���@�e+����X��l$%9GkK*��W�P�Dx|$�L�z�
�3<�B#�H�7uJ�r��+;�)�_Ú��M�j��?�3�ֽPˠ;�mn��2����#���|NۅR�Ϋ�"U�l)9|Q�J����`G�w%]V�Oo74wX(9�4Z-�ɪ{y�B�
_A�,�؋��/?��`��ߩ1��xO�G��bs�+zv7ƟOt�&��S
p'�`ig�ck�.��}To6�%�s9S�k"k�+�V�nG�޼S�^WF�eǡ�A��*b|�-�W-Zw.�L���dKn��52+FJ�U�^2��.���Mw��u���8�z6�da�N&�+c�����Cb�/�a�X}�w�o�8�6j/�l�_���O���z�����Thؼ�6b�22.�1�|�e��-��*&��v�8�i�ݮ���v�9�ٚ�/�׷:ݵ����o��? �S��ayg��7m�Q5�7-�5��6���&���;�Ns���[��Q����rǽ޽����NGh{�]yW���Ҽ|)�Yh���Y=�:�0�5W�n�d^{ޤT�y�"��"LP�j#�b�������B�u#1y��8��n�,���ɽ�lG�T�`t����B{���%GD�=���)z-^�Q���n���s9Y���3�\�iљ�8#��9ln1g>~��8쉯H!�0�5�}'o�#����a�����U�o�.̬�$�,;&�TAM��Zi����=4Ќݪݡ��W��8�a6k����°Wk��K�`B~U��߼jVq��w��K'S�n�a�G�t�a#������a��l��C��չG�:�Y�κ�l�Xh^����r;�����Ύ�6l��?svL�)NZ���`^ˈ��l؁a
*o��p{^Wb��zxW�zIcj��+gyVAn�8Z�������pvcm�,U�&���NtJ��ux��={�}ex�CۗSnW�E��';�Du�[Rt5��8
���ϗ	�Q㢦�|]Tp���us�flF�<�_�n�N�}^�o�`�}������qA���e<�����ΩWs=���%�����ʕ�z��%�F!�Qc.��+zu#c�{��"�����w�����ߕ��+{�tޖfz��|�MW��\]�i`��\�^>Q��}���qN�(���;�� {c3?{.=ք��#�欈x����`���9�͚y�2f�$lh��}���~-O=��g��^{�]�g���V}`4��⩈p���:�~���� �͚S�>���t=Xk�n��T��{=�|�è��iƮ�FW��&�r3������:j�a�>�Fؗ>��تr��ۓ��>�Clu[��`tdHy�X@�#<$չn|U�lиg����fFp�_��*���.�F����M�7M֭}��S�|/MUr.l���a�u�*P-7�@���j�V�ۜ�!��i��r�]�8�A�,�S�A��c,X���[��jb����of0���_5���A��$4u��-[X�le4�»����`C+�T��q�X���mdF�Ԗk�j"�̏�����ȇ�_D���E��<n}������=�P�x]9��5<�[�^(�ī�pO���+`0����8�^L�n>�����e�eb� &���X5���5r����S�E��$lI��W�+��*P2/�]W�:��7F�z��Ź/8����������v��v:N'D�9��*jf0ע`S@��Rݩ2\ݿt���ƠyD͖�2�包�Z�F�6ܨ�T�m}����qέ�����"���❠u�\L`U��n�:Y�8V��eG?p(�;�F�`�y��c%<{�g�8!�#���}B5/����ƕ=k�Rm�	�&�����ʜ	��r�Q�+8a��!�5���5�O��ȷ��i{L�Ū�p{�)de�pn�GuDL`���mE|�b�d�Lh�Ս1-�Y��`���Q��[�8w����7��I-���}�}���'B���Z��N�� ^)ܬ��52��2+S�n<�I��M���T)
�3fM#)2�],���@}�?e+s�<h�ʔ㮀��hƔU�}������g�N��ů	]3+�c�f���(^B͋�h��ys�Z�1�ccOB���׻�5��9��Y]�əʾ��;�y�<k���X�V�,6v,o��ײ��!>p��r���)z�n�U�ܣ�.��<hu`���0��u�X\���������wS>΍D����C����<КA���n؊�,>��_����]���Q�҆�����DQ$!�/���]��A�t�Њlg;��M�u�n�������]V�G
��=o�%��U�=R��h=!te�_��6�]��9������Wy{=���m�e��F���J��u��C����߶����Fn�GL�vۼ��$y��ٱ_@��GN�]׾љ���凃���%WG����̟�,n�&M��������2��3�Jʬ�q�����ޡ-�����+�Xf}ŗ��u���}���{���yv3ۛ~�96��H#�}�}!�u������5���U�=�LId��k��֊��i�p<��IJ(SJY��jǈd ͼ��$r`�� ^G$��e�M�v�8�I����C�8��D��g샥Cz����ئI+�a�Ǖ3�+�Ŋ�R���q_q[Ҧѩ��\�7`�Q{/y}��~����LX�}��8m���Ҫ��%���f�˳�R������%�r�:�=ܲ�z�9�0oi��y��'��"�oy�
�<�CڇO
�)4�YtVc����a"�mMЄ�䢩�n�u�헴e�1��o��ꕯ]S�7��uZ�3�)��+�M��nf�CCn�t|5'A�X�v��*���>|��P��
b��Ϟ�;kl�ה��V��o�6(�,r��'."���pд����{�4r#t�p���U#%���s��F;jęv�(�;t��b�C���ȷi�uygh���1��Y7�L���%D,S�Z�*�Qe��4�Nw���uq#��V��!��2�qP�!nK�B�X'0��a���ֶ-�*�Mw^�\�kM�%�^�wN����f�4���� ae��AH�0��S7k(nIշ�F�,��q��#�IMH�������.Ws�o��)/!+1CY���N)q	��Ƴ��X��>�W�=�{�����e:�w������OM�9cA,9��c��w�#+\������u}�ك�����OR2
Z��y(��J���B�l��*�ʕ��CL,��e�}��]�գ5ō�y7��ؓr��ӷP���n��~�f�_{�m_X�n�%i:-�2fHT��l��g�Ŏt^�x�*WR�p�j���n�{�a�l��f�)�c�|���eY�-�f�k�B�l�ԏdY\j}��\�p}�
{S2�C�p.��^n�{��uI��%>
bV�<�e �!�Z�uˤ�핱�n�nt2����P����
�� |!٪�X�p�T��G��t��*UV�:��o���>�u�Ʈ-���]���8Ʒ��\2+Bg4�`�S�25����ۧ8D�կ@���jq�Tj�>���]��	��:W9�_b�ۚ��)'�r�Ƿ���֚w􃯦�y�o3��2<Q�ۮ��k�e���E	�5k�]��m�9E���'`���5��o2`�#��C!|q�}
�Łvg]j���jY�|­����܎�t�F�d�yh��e��dmo�D��l͹��Q�h3��;J�AnvƊ<Z�NF�̂e铤� uwk�S�.hAmN��3LV��ν� q.�Y�no\m�"(�U(5�Lu;u��R'���K��fw}hV��ܫFn��]�Pk."��WL뛂<ٲ鰘�_u2DׅXz���������+�wJ��li�Fҭ���c֋����
/
��HoR#�5��ӑ���]a�K%�}�@y �^�[g~X�JѴgS��F����ŤԷ|�l,��n�>��&���z[����%�b���D� UD��pO�ݩ+��R�w%\��EF�rŮbNYy{�7���mr�so�^I]�M�p҇+�˙ݷ"���ܢ�W9x��y�nk����w����4�guu��c������m�nm\���-�rn�A�5�.���E��ۛ�wQ�X�+�"+;��r��+�ׇ<�!4Z+��F�;�'Q�X�k���b�d���]y��ĀX�c��cT�acX����x��	�r��Wwh��Nv�n���s���]Ӹ��Q�\n��v�r鋚�����9�b�4��܉�9̖�n�
<��	�W0'wW;�%�仐�M�s&,DWȤ�;�2E�-��i(��wW9WH ag��^1�r�F���ƹ��h���t9�9�m���C˷-�;[���x��Jy�"2��b����o^fb��xw���qM�oX�Y9�4�61�3�t���7>�Z��Rͭ�:�%�볤��3=��@T��lg(C��_��5#���
����c�5���o$E���%�x7D�!������&OԄ+\�E�dz�-�łH�j�]�B�~T6�y_g�=ϐ������>���*��(<�W��0��G�UgD�=�w�yߴ�	���/�h$��	�JW�m�iM��Y(xeGz}1��&Lϝzm)xD�6�����&��FF���؛Z��V�h�Q�����`U1��Q�i�&+���7�\O���7���Mm�n��o�0������}�ݳ���[=W�@/wE���m��=���ɢ4s�ez���M�i�rW��	�ϓ�Y����7�o%X͉-��C�"�
�A�g��/+'�c/E�k����6�BA�i�	�;O0Of��_�lP/��ȝ�C����w��zw���慱�X;+���m��������t�nKi�q�~�i�C�E�Wy���a����Br��c�9E�gJ�`�5p�٠�Ȳ�
�{B�m|FV�MKK-�d�ʲY$�PfV��	�������6��ۏH��w���U�Aw�[�q��:�<�"o����f9���l���19�G�]�����41��׎ ���k�)�/`�ᯣ�x�5�S[��e��""�iC���d��c���Ŭ[k�݅���|=�g���T���_u�FM��E���i��>�8�>�!��W�����+��_f�&��w���+�Y�ak�ϖ��z}ʄ��ԵߘJ���'�s.gk�]�E�����$Y��YYo�P�[�@?@ Ā�K�k��t;�9{�W��~��yZ�MS��]����
�������L�~;���j��i\���b�mb��%����#�I�
��U�pě<��:w��$�׋��P���.�c�&���+���D{S�i�i�c���9�k�S�3�ʕ��c��Y*Ǫ�TǗ�����}��Pgfs���R�,�E��3%Gz�H�1Z�ͷ�r��'A�7@]n�r��ޯJ�t 9��w�D]�Z�L�;��8ec�v�{�_�$>���-|:ɽme��hg@9T�7V�ƪI�挗�t�c/�їJ&�:f��Q��@s�k�)��Sy��J�v����ǚܘg�A�$|72(�jj�6��L����Sf�v� վ2��I�]�=��}�������5�~�v6�]����-�n7g?V��"����|c��-g���a�û�qh�u�>����`f�!r�q�9��Y�u�w��W�f!���["����#�O��չe_|'�{')l_�>9�'�]Ww&W������lH����"�y����lGShĤB��U�����{���Ψ��1>��>޸ܓc��A�lt��HN��XJ޺��k�����b��{�7�d67����U���O��yz�]p��_J���g�ki�{����Vd_�^�J��^'���3�u���Z0j�@f���瑮��~G��s+���5u�ז�����8�:)�Ϥ�UO��q��62�rM�F���S�H#҄��t�6�X�*�ك�g ��ϭ:yc�dKj�z]鼟^�jg�C�p+�۰lX�,jS$)���D��E�"�����=,�	���pm\�<��&+y&�a��'hE�+�[��V��SR��m^L/d���u;Z4 �u�X�9$Q���+��:T.[��q=�]~]��ݱL�~��ߍA��Y�Pޣa�2%G!ݦ�[1us�P�[Z����,�c\J�w��I7JK�>����}�q11������O�5R�˨>�*z�^h��M���]�ެR{f�����pGTO5���0�31�Ə�咽�����$����^z�o_W��زk!*Ⱦ0]�R���V k%X��?T�n�D�g^x�μ��m�b';/qx���6	!@��!�ǆ>׆�U����3#q�����V��	�^f��5�x��W�a/0��쇾�k�v+�J+��3�^�R�j5fн���ݶ��������P+��y�g�y������^�
���dT�շ���P{�V�U��^d�����DVz2���l��/-���5�}٬�w�(#N��-��G���Y��6b���� �3��s\���:ߏ�]��XC���6��s�va�=��飼�������
S�\K3���ͻ�pOi������b}0�{!����S��d7�ԫtP�U�����#�<��=f�a�EB�.S�Ď���-�׏W�9u�oWs�b�7���{�|����[�v7�"]�4�#�R�h;a����蠙o��a驳�����
����;{b�熲�s̭�Y�
D�lj�Oy6�"�z�����-r��n�r�V�g��r�p�tt�{r�;gx����+w�;7�����rCwF���+�to3�|f�ō�|�6��l��z�!�g���{��̀�#~�P���o^+�Y����CY.�8�禷d����h^ߛ`�	��@c�@�BCj�Z=�x���=>���T��S>�d���F��&#�A��8�~g�T~�
$1Ƥy�����N6���ks���Lt������97���3�<�b�
�D��|��v�^1^yA��͞�=�w�=�w����U�eB�S���ʾ�sgy���;�at.��A�����{�� �����JB�ɶ-�4�c��\�˝�u�ҫ��\ܔ1Ď_R�������}}͉��j
��1*ed�u�u���m8c;M�ߍƄ�Cu���m_��Nk�ټ�=��?���i����8�)���8���,
U�Z�@q	���˲M�t� *3ˀ�]$)ʉ-cv�ۖ��A������S�!RQ:�U��7�fNk97�07�g)0���x�MΉSV9�dZ<orSG�,^8T/{'�rY}t�p=9���'`c�X�{�=7��z.B9d������V��=����l�|��,vܞ᳄���߸�;{���d���[���b���6�Vlham?Z�c����R�_�KQ��Fy��^F��f�H��v����������ظ��f���h�*�zI���=�n)v�)m��[hGZ��x$骿�J�h�Zu]�9�)������#a6| ��?/9����m7�sy�<.���	��'���1�zfl��#�}c�C����唹yͭ}^J �x������]\cځ�_��6�Rx�tE��uOϠ�<+�<��$<c�P�
��5�jo�{q$j�.�XwZ��-� �	`��g�dLI0��QSz&�.�O�kP��8/6���iee��rǽ����> �J�Mf���P�^"�_j<=�����m���;�*h���.���"��	X�LÛ�_#��+��K'�Ҡ�M\�#�a�t�ԧ\��}���3!��g1-�8�ܦ6,�n�o��(k�R�=O�Q�/���9�����A{��f@�n�W%��'-j�L�5��󋛶�*H5��gj�q��6L���|�p��<΢�N����z�S�r�z$�1/V�^��=�4s�&�¡u����^]�nW��Ί�E�*D�|3��At8yD�[]�oA ���:��e�؟^��V�`��f:�BX������w�aU5\�o����.̈y=bz���x��O	_.�?1`�+7M�ߺ�A�7W[��u{q�]���"�ϼ�5�&=���ku�4/{����?�������,^��d�C׻��z����
<Z��]"��0����^��z�v�j[�������]���ɻ�P�\)�
Lzp�'\s	�.�mS����'d�B�$�]�Pٚ�1�͊p|i��Ӂ�B��4ڜo�b��],�s�͡��U��W���f����7�:��!��HNל��]_K��d�W�ch��M�Z#�X��%�����mJ�u�P��)RVI�����|����֔�2�v�[ӗp�q�C���S�c k�9 ���:�t�ok��ɦ#�ă��K����-����wJ���u&l	�gL�����뽘;{Q�r�7�gr��U��R��iS%:]7L%�ݰ��R��pcz��f�ϴ���g���[7�[䣻������#�]�b�dd߽-�㷽ү����5�)���^Y�}a���Y��:��g�yT	���f�7P��N�e���k�hH�뮾Y�J����ϵ�E)���u���j�,7	��I���jbn@�/�:Z\�j̓��,jS%O>�Q8mx�tx�&&ɽyT��B���ް�`�@���R�]��pT��4}�T�NU���E�yU�YED����f�t��������T�Օ���N�bݾ��;����o��l����ɠ���BeAp�f�oި��U\4���ԩlLN�;ش�{+H��>��M�$W�a��^Ń�d�FS�[;�zM��M2=�1h�����=5��ɰ�����[gb���/Є��ji%[ꚺ��ɜ��B�O��q ��ho��Y}���]e��>���v�3��\H�%I�������XJ"��<[�j����������ȎroЗ�h����m]�E賁�#a�C]ͽi��Y׷��](��RRd�VsWo�֬�)�˳i�q�t6&�M;��+����hs(��o6����\�;1Q8d�ow�z`��Dο�������!��"�͈,=�V���ɿY�f;m|
�*����w��ؐ��1���=o�YS����֫���gk��SM���5EY��`�e�ޯ�!�����IS�f��׷U�1��k�b�(3c��G��f)�e��F����z�<���S��ަ|4'�}`�ϝ��<v۾V�PY���u�gg�q�\�hϷ:������+��P;C==L�yg�y�����ςv	�@7fr��uU�&���w0���>T�T�/�W���GٜYy���dY����Q�CP�Q7H^�i�h8����*�Ƥ6���V��2���Z����]�0�'���Ȣq����,����q��y��O�#K���P!x�Q����q�k>�No��z��]`�Ձh�J�~!G�)��`�SP�$�_��h1+����c��Ђ��"*�䡓{f�+;8.�݋��On|�ׁCk*�#��=�9�}�$��]#!�ڽ:nmT�<�VŃ�f���KU���qv�F�R���ܫ������v��=BV�p-k ��5e��Mu��O&�"������	Z�*�*��g�Jp��E�z/�g;��pe����B���M	��>��5��}�BID$���0"$����[��^=�u�(���yed����!��[���a������ߪ%(��k,�|79Z)Ɜ����c�Y(�g��@n����+�X����`8��!̢�9ۜ�_ d��\r�g��ݏ���W����J������<g�f��r���
��B���j���_����,-뮸/���q������1�/�>g�ό���$[��O2H;�=�{��Ǿ܎�ά��œ��oB����z�Q��B�J�m��[k��V�Og�݌�q�lU�r�����(ܓ~��қ8q�
}��4;m'��>�Q��w�g�}=��xBEDOz��dٱ:�d�ǨI����ym��y��}^qN=7���y��^�^�bb�ē�y�����b�A-' P�r��L5'S��a�O�#��ν�E*Xo�0�MT�Ȝnc�U���)�$p.�Ffwu�ViܳZ���N�톰z�Ap�$���F���.}eޞ��.��2�V��dk���̶���|1��خQ��Qn�ʻ�1�H?�u͖%19�D��]ڳ��yƝ�c[�\�PZp14�������X��s����1�)���;�J�V�(ROP\�Xqn��!�1����*�<ۭ��T/6KƸ��K��*M��+�Ȉ���)vݹ���Nƚ���8�X�h��.�Z��Jý���k
H��ʎWk����jt�N�T{��I�a��:-���
8uQA�W	C�ٓ3�cy�Yߙ̮�i.��|7Ao@���N?N�<r�����	�!8&�X(��pwq'u7i'i�o�X�8�u3�m`ko;�ʺ��`0��Y�	I�ܘ�nM ���ι,J�]YM��ek�ku�L�2�ʷcY30�c�gDԧ��@�f��g[:�,�}��ȥqBN�9ƹFh�f	�P�Ԥ�Ր���|�w`�[e��c��jQ��dƆ�vm�B�F���;U'�\�v�%�Ŏ� lf,�;���;˺]ډ	����b�"�-�xFFV�DwL�]
���e�	�{Ɯѧ�nd�x�1L��"�Oe�v:�8�a��e֨�o�K��Wo	G�\S���J�a2�j:9;A^ofc�);�lp�㐴����^�;Sc��{��n��Vלz���ysei�5#S�|�
�e3M����JU�m��=�cD^�{��gV�sh�����{��`�/���F�7:P���`��&#۲II�N[����*M������(��N�',��}���+)g'�l2V|;�w[�!۽�Qv.\�8S,Qxq�>�c3u��]ir��J����vĉ��Z�^Ʌ<'[�8��U��o��f�.�$��f��2Y֒��C�G3v<X�c�i;�:�2�{�CNM� �ݐ��:Fj5��N�C�݇U��'�Ie��tl�(��/e@9��$�w�6;|�z���fI8Y��|]�2���چ�FR:��S��q�Û���	Fn��&WZ�B��`�t�ˆ���n�̥/��O!�v�	gii3�V�Rmc��;ٌؕ�5�ƣݡP�Z��[���I�9Imk8u�gY�
����l{HPj�p�zÎ�[ �X�vV<����V^�u���ꮕ�oq�{3e���V!s[���x�3W��d,lBটM����I���'��;�w���{�1,�_�=�i�]R��Ҋ�<S��z�@�CS�C�֘99��z:�Z��MusR�Y�C��3����w5-����a��Na�ɸcq�j���� XU㫘�t��Ğvo_d���a`�����̨���0��UJ�$Q��$��Ĥh���_AW�B�.b���#wq~;�6#�D/;�w�&ww.��~/�������n멷7q۰s�s���D��35��h��M��{rǥ�^�w���{��;�v$wWb�$w��WwR%�逗����n]#G'\�\��Ʒ-�e�W4��ˎ��LYr������.R%Fa$�����q�9��E����+�9��t�j�ך�%0h���$�21��k����R��k�����a�w��guЕݫ�W:d��y��:���:�%	Ӈ:��r���:B��\��y��W�I�(���®v��:x��<� \�we�"ɢ��nsN���H�p9�t��&&��u�	#R2L��v.�7us�9��:��;����	��v��v[��]wp��8�NsK��1�k���k�{e�~�2��O]�s�������wX}k8WZ�p�ܐE����$��k+�dR.��-r�ř�ﾑ7Vc�2��$�W�9��&����W"�GW�4Ѐ�An��y��l����hGg��oٟ6�_���+�����z��U��瑣����>����=b�;Z�^\��_,V�`T��/�ɥ�O�X���$�G�}S�.��+����y;����_|���!WW��?���{^\s��\��c^;��q�y��m�-ď�A��բ���Z'�i`�6�P�qwb,;C��t�C�I�#�U�5%�ˀ�z��|ނA��:��d-�3AJ�;q�|>a#8����VI�T0��^K[ߍ�b=Q5�+2S�T�{x���]�7��M`o�_��+ᛎ��U�ƃ6�j"�o��ۜE�z#9�gܣ H���/���5�96;�V�[�]�~y.���ښ9��FF�ƻХ{C���I���m]u����0�k�a��ϑ��k�WgM.��x6]_g���J(v[�h��z�i�4n��*=ܜl5w9��Bݼ��E�"��;K��<��ƨ\�.���-qj���[��ܽ7K욇Vԣ5u
F�f�ݵ�]�r��.� 6nWS�޽[}T�V��4�f���8q�1�:��$p[Z)�d[b��'_X�a<.��ڷ��������g7�0�E� ��կ�۷�e�lH����CpE4�HЂ�~��蓗ձ��P{��v�w����>��m�#�O�,l6:x�t��Nߦl��P��'b{|�Wl�V|��V�Z���K���zz����>���+�w��R����'�b���|f����c/S��w.�V���G�\Xvr���J��O;������>�Y��:��g�yTq�����6�^���9��`�PW�u�4�pT��ɳ�k'+-<��LGy���7?j��dL`�d^�D�G~�
�j�6�w�5)����\�^��2���{L��!���=���:~�A��K<��*}�!_ky���K�}�3����Fd�^�m�p̈́�X|1���p6U~�P���0�ɠڲ��ճ��s�������>ወ,j%�׻.kׄT�F� ���l9ar�X(:���>=����۹�%������µҦ�M`gu�%1Գ����7�d�64#!b;.0Dv��w�����溏"s���	Y&Τ"N9%�ܘ6��[��D�[���	{L�#dX��ˆ+��J��
f�V*��a����'��w>7���Ͻ�M�R�,F(}�l�3�}�:��y7��P�C�5���-g�����a`�+�b�l�f���c�/�d]�;8�&���ʰ���n����a~�����<���zi#��s�C�uI���w�_�;��ג�P��)m��!��"�ϓeHg�iEqb�)K�U�_��o�������K͉�ΐۊo꜊ܜM	3{�ǽ��{�)+2�z��m�!YY�K��.�D��׫)�?�����|�|�_�ܽsA��P#�����e����D��6#rRu���įN_�B�ev�#��Xѕ��#c���o�m��X���9��0q�N����q1����o�s����C��%��F�UtN�hjfo�8����,�.��c:z,�GOuZ�3��hU�8�݈�Ћ����r(�q���B����ax�=6�R���s$q�[y9M� �.uy�;I�|���ż��W�{��p�u0�c��M�3��2*4t5%G��=��0빔X�Ȓ$�&���p�j6eQ���eШ�e�yu����(�x�1);q��p�x��Q͞۴`�y��"���pu��#�P��	��G��UR��o-�J���~�"OX��Y�����3˰�q�h�pX!Q�"`1ŏ3��+fG�����^T�Ǖ�%��si����q�]`^X�
�UI�ᄛ�֤^J�]Ƭzu5�X>���w��+�,�^J`�W�E�}�_mK��]x��y)����U|Ƹ��z��i �ڄ��������#ެ�^V]z�SvT�~�z�U�8�T�ɫ�zۙ;;��n��r�����Ǧ/��At`��"�./}c�vć��ʞ_b̟�������
Z�[W���E{�Ը�wɇ�i=#�������%�����UN��6.ҵ����t��ȿ]�=��kV�������^J��c�W�y��^3���JJ�"[����Q�Y��+�(�(i~���7�T�s75����l}�����n�@ǽsi���9R��(>���*EW�(�J�s���6�w`ٴ"��S�+|�	np2��u���2;'o��2Z�Å�]㤋r����<3uׇ8�hO�|���Aa�4��x�<���}1Ҧ��h�
�SU쭭�S��>݉��hz�R�!�Ҭm��M6��Vj���E��+��Qk�O���Fܭ�M6����V����k㶓����D:����9��oُ�W����M��u| d�ǨI�9��۞���(/$�S��,�XnP�����ŋ���*|5r+���OϲH�}c�ol�-����ksՕ�׍`\�1&���ܫ��_�|���!��Fz;��{G���"/�� W�l	��+G��ʗ��8�YX-����r`��KMM��=յ�Q��G�}�Ƥ$�z�{�mpT��=~ϸ��Q��7�-��������d�L`�?	�IhMv�����l�_�7�Vę������N���p�TO��,��@�0�p�&���|ޒ{x�������G���v_T�x:H�v�Xr�=�5�L�TL�)�]�uM�^�u�"�M>�+�G-���vq����hܻ�����{�J���J���20$}��a�o�]Mk LQ7�u}���9��� ڝ��>���Q}x�����K4���_������V`��aS�Z�f�C�Z��G�
Nb)DN�������j}��o��Lp�k�d�������JR�c�}��F�T[�-�[�5�ͱ�|¿��x����}��o%�A�.����W2�ȁ+�꭬љ����o=u֋�a�t�.��`#Q�"�}����yy>�������hO�yƿ��e�s��p�:���]�m�U��]�n���6(/�ۊz�x@�����2���zs-���0B^>�A�y5�)<m�q����"���{bb+5@����ȭ��,����JXJ�{�2�ϣ�Z\�%�b=��o��=��ԟ�E�mW��|{�܊�6��Q:���l�e�>����z�X&�&2��� �������f�_}cN�	����� �����p��>���G�*�[� ��U��ғ8s$���\P�a�[�N�mg%NY��&�Ј=͵p�v�a�8�q�v�&�'���bh�
*ÏY�T�L���)^ѡ{� rV�m���]'k:�%:����\�#�Bj�W`n��LqN�u5����i%�Tk�;��Kd�V���6������V�]|�X��K�ɳ��WMO�z��%{R=h^��� O��=�q�!�`����<
� ŗ<��ה�lwU�q����)��]��$��;�3_	>k>��~�/(��{P=Өb(��h��t��;:��O��q��o,nz��l�)��7s��`�i{M�h�`�	(��a��|=*�zz"�חq��]F�z<A8�;jk���Z�G��$��|�9�_kFb��v�\�w�_��Tܛ6W�c��ִ]� �^�6����ޱ{5[P7�0�ook��$����+��F�B������fsX]a��$��=��@�_�#:�¾ŊH�IG#��r��X{�Q����[�4�8�ԗ��oy����Y��"=��)-4�_<���7�_^D��|��՜�z�9�M�AU��M1���*���a�/��WjN<�8k����5� �5���?Z��FK��	C�ܳ6ج̴�xL��wR�	���d+uS��܆�������r6�d���"(�V�:BQu������;7o����t�ݿn��3���=}-��i��*����ܖO��5��ז�3�~��A��x��ᜄ�C�hHb���iw�[oL�l��g��]R�Y����v9��6w�g��/9��7���C��e��q���c3�"=3i������O�n�W��Y>n���ғ��K�Qg����#;�JW�_/%�]���G���By�Ϣ���x�S�x*�:R�Vq��/�{ؗ"���}�����v������Fm���&hl�ox���ε��p:{a}��q�ՆpY
�D
�AQ~�p�[�Vv��}��<6P�ޮ���sesi����^���,\�Bcg����n�6{n��3��D���q/{G�7~���V���^��s�{u�E
�$�+u{���ڱ��Ap� j�4�g�|֒{ڦ�)
���o$@�U}��
wDѨ(���k6�[����Ǣ��)����۞�g����aY��ė���W�N��d����(�]fԴM�`
��[���5rY�hi��;5�+wX[jŅ��ӆVK���]%�a�kp��'�wb��[���l��7�e��|�U���{�����K�(tܻLK
��Sm�^{�޾G���:d��b��(�V
�-�}o��M�����{ؼz�|߷㱳	]��Ǭ���%շȶw�&���&}7��m��c,��ʡ��P.�+]:�}���X�[N��x��Ty������gm�m��d�V�\YW��P�Ƚўv�ߡX�W;x=�-1cO ��Aa��Nq�x��{��%�_������_fA����c�"����}�T�'z����S8j��L^�n����R�pp�F��eKO��|����ꠇ#��ի��]\�m:���-�n��u�t؅BO�1?!�}̑���n��۲����ݼ8L���q�<H�\d�S���@�B��}�����=��}��E/��ya�g���f�b󔻻����쉸S�2���Ln��I�j,�N��AAP�R�5l�+æ��͝�J?LΗ,y���h3:���B��b��I�5�j.���{���=^�P]�X�2�"/s���ￚ������w6l_�̢��A6��
w}]);�v�'���:<N^��h��]��@�<��D��v�o���P���e�M۰h�ϑl�M,����T��S�K��]�of��e��6�������U�5c�w��q�T���B�.�צ�����lA1��DN����#��H�~��'�X�C���)��(�Ck;=/�h��]3_���]eQ���،1?0O�Z&���l�#�C��)���ub[3�=������6L�>�ud�L1�bߟ��"3�<VQ�R���݅����ǿ>��'܂�����n>�����:���Dz��]5��7W�59���>�[ɱ���Z�&�>����k$3y;�+T�����"�r�}���۶�[��SȰ��L;�K����e�o+[vI�5�*&�q�X��7� a�`���-�s���~�C}_�eJ���-�L즲�'���&;m|WY�)�۷�=�c6$PR��	���� Mϣ����&o��n���=�U�@����)� �}Y�z�zƝ=yYs2�]3b/��Y���"jn�%Z���"21���Y��ne�E\2��FY�Z".�� �;��"�0���e��q�{F��v��sNSZ:�tO)�T�ՍN�h	1om{TD��p�u}�+��֖�j����Ya_]7��[/#���cU�Y|d�R�77���2�,B�#x�[�\%���.����+j�\�ћp���1�]���n��
K�Ӻz~=\��CG�vP�vh��:�fPY���L������ۣ: U6����S)���+;��w�����żΒN4�!V1S��B�qR-8ro!�x�Z��]p�ڻY�`�Mp�|-�K�7���cg7����o:n�l"7q��3��k1�9������YK3(�:i�At{(�ʮ|���tz��}��Q�Wo��ž��:�zM��B�R���g6^sk�R)�U�Ȧ�\d���Q�AӋ�N�VRI�|��� �5��3^kp-Í��+�M��9�$[�/�-)L�y�j��;-^�EM]��b��K���M<�(���!W�2�J�c�tkc���
�P�<�4\-��c_��3I����P�Tl�JM�aLβ;::�&�b�bԄ^�>����u��ҙ/$0_r읙��<�֘��Jɮ�Q7k+��ۦ#�㲰R�}�P�>s�ͮR��#���z�rj��.���Xa/��kaL	Yqe�3'7گN��9��76AyF:�#=Iv��M�r+#6�K�x�TU(hcqV��ke.��n|���i
oXj;�N�����H�"$[�V��iT�4��´JMl���5`�oD�oz���9�R�����\�z;͊�ކ��% ��#Wwg�3��7`���t�yG�F�Z؇��L�+`�Μ�̼F��:ZDgFXoPMHL� ���ݔD�Y{(KuQ;K�s��Z��ɂ"r��k`�Ǻ���jMLBƏ�>�M;6l�J�9��:C�=2Ët�|VL�7����t^��*v1�J*���r�Cd�WQ��V>����҈HorX�0��.E
)�u�Y릝��6���v^��ۻt3�ݏ�r�A�B�R. mUվ�����y��2�T����9��s�Mu\�kQ�3tA&���6���lJf���u����i���m�������M3pP���������	}�y*�膍��󺸛՘�y��H�Iu��Ϻ�u�в����*w���[���m(fAΫ���%w��U��*�rP�����6!ıg^�i�)���bgx�cjܩZv��<�6V�m0���JI���h�p�8�ݽ� �V9!�#�v*����q�.�U�,����r���[�8VKɝ,��ҩ�9;[沰MY��W�q��-��ܮ�9^m�ĚY��=��Y2�GE��ВKF%�&Gr �.�[�:���V��q� Y]��� ��庄R4˺�ٛz��w;ɛ���}_���{�♻�&��!9җ��<�cnw\�5���B#s���v��^�w�����;��;��wv9�F��	����B�ws��y�����a���b2��8��%ˍ1˧wwv�@wrln���#%�v��r�wx���u�,!��-��\�N�������ۭÄ��u��@���x���Zs�Δ�wtwn�鉹�K�9Dd��\�I2�%��wW\뛙6b'+���Q�;��!�Ls;���'��^:���s�ww"I&^7/:.	����\H��0���,��2�w�:26c�����d�N��9p�t��"r�\��:\e��s��/���\�F��ԏ<���#����w�/Ȋ��gT��dY�8f77��Q�/M^BAi���2���V���c~ݛgpx#tB��&�JCfeG{2�o��x�n{;�%���/��� ��(�w�E6���2w:��e���ś�� �ҍ6�edu�	s8�ޚ�\���V6�׺����X6A>�q��m������=q���=j���^����u��p�y��h�d���u�j��������am�&J��9��&Q3�l�����j 1�Dy�hK*믞X�*^�M��h��(�]�;�`��n���X���!�e�>��X׌�5QXjf���2Q���0�%�һ��s>����4��}k�>h�簝���؄w7�jf�'7/��8���8f�N��~8!�5�xD�`�R�	�z7�u�	B$���E�$�>��*�Q_6F�p��`
����Ǯ�q!��b��M5}Y�h�U���	�R	�ˢ""k����z����ֈ)��P7ȸ������f�N���;l�[�9�;2�e�����n)��m1|������a�Tݻ��u��+ؽNxdvn۠�9�ö��cf���kD���WE8��/��招��R�*m\�S��/N�s��i�!Ē�bu�+��5(~4h����]n��]�7����0�����F�xy��u�J�z�,^�{��e��07[[�]�4�]e��M����D��Y�>�_@�'�ԏak����n�{�%��%f�F�V��xw޺雭��:x���lSN� �mXZmg���.�_��h^D���#ΤK�h*�N�tk����^��h�"�Wj��t�ޅ4��RU�w��]+��W�ˬw쳼�y����u��HB�����-�b�6Uc�J�W�ǳ��'p��7K���xy�=���@�T��m������ �gu�%��@����s�|*�0���=E��u�ax�\�������F:O�.�,�"mq�l��>�d��<��Rj:�t��Ư>3�š5���{0�^d��}���� w�XC�
��1u���'�����j��]���z�����VR�:j�UX��1j���M�Zf�U��6eo�	XE�u<}�C���o�Fˏ6Mɔ��8=�#�V��
�N�X',5�L��]7î��`A�C��S�][�Dw)�yՋ�efĻLC��N��]�}��>�o���yާ���y󧶏>(�h[j�8��������W��ڣ����8���3a�yԎ{ ��/6�>;m׸�x-G�W�x�Sg���b2�b#����b��pz�w�v���*�����хKkxnp5�H!~��ο=�f�X\5D�[Y�H5���o�~�(Іh��� �1s�
S����N�aN1�WLl>���4�A��l��!؛�{�/!;��<�	:�XBD�4W�Y�VM �T��ʂ�3���iθ�Ϻ_Ox�K���e�U׳�4�~��oq|,&}�~y+�=N<)�-�e�����2��D�BG�u;�q���G�{�ŷ�Z����ֻ�N���j|�w}>�1�pLK~ؐC��^��la��>d�s���{��*�]��1�a�Tա>�녷�4��hz⛰v��U�~��{�~�xЀ�7ݵ���s`�7ɉ++�����3xP�hc8MA��-�
� 0���ҿ�z�?ke�|w\q���đEf���ѳ�4cnϲs���S7{z���3զ�~���M�skC����;�s��Ns,�Ԕw���$���m�;&�9��9Y}ފ�c�l���"�`�����w�!�%���C^�w��:� �M�sч�����V|��=�n߻��6!GT��bD�PE�9{d�vͼ5�;�N�����4��_,]!���<�Oz<�i�j��u�6�\����xiBxz�����O?_��~S�.�_�|�{�/1���qk�u3p���H|�W_<7n�Xl�ieS:�{v���NzbFe�g��L`���~�CT�5`u����Ϟ*}@����Q��k,r'R�՟���~�g�W��uq�O�5SڬW���yGg+#L�+pK�k%q�,�+�oP��UEp�lF���'�����rȸ�.�s�6��G�5��Tv�ސ�{~�ܰS�\�1ap۰:�O�1��
��P��ށ�x#�}��N���j��[�]?�Bo�qK�j(�wՒ����8'Ul���
�@2���Y]���rߵޯ[�h���/���3��\��3UAw1Ր��U�lF�EwT肍��Ⱦp��K��e�JL�*��b�1Q˔�qyL�.�̺��<e�K�=��yg&�{�ҟ:]V�g<iZ]S�4�ɧ�y�Obˉ��%t��j[��n�m��9����X<Z�k�;눺��٪���Ϳ��r���\N�߄���O�^�����N��盵יS�D߳}*�i[3�Kk��m�!�������0�:��뽈��*�1(���%=������չf�n�=��� 9C,E4�۵�UVm!|Ͻ�{�,2��%,��%�$��i�'h�ܧ�r���e�-f��t}��qۚ
s�^��|��6��,��:Օ̥��{�{o���1{��eq��ԇ�����X��},��ۼ���:�=c(�
��-{=�"�ί��_�3_J�W[&���W�Ҁ�۬��)D�ؗmU�&�v�u���f�L	퍠Ǻ�C3,�������,T��	;���l�v��[v��%�ʰZu���; {�{�!�k~6}>���yHB�䗰zzco�U��c��VR�Xサ������$}��SE�QN�BD�M��t�D�s��$�yӍY�7B��q���+࠳�JQ��o�-l\��`x�$�o�qM�7�ꈩ��b��Ѻչ��s�U���%�3�J�9M�8d����<�Ǻ�
H��lA��wЃ"T��>D���9�ʼ��hx�K��*=L���?[ ��f^Y]���s��ǔ���>CV��>ZH4���F����V���j����],�Ü�u�6�u<PcU	���՘5�_/{P� JB�	��y�aue��4���o��V˱�D�:��wZ�w��yz��l&}�cX�Z��g���uR� <��H��+����n�����39��^?{E/m�w�v�;�W�sO{��k]�	��G+*�_��%��7�B�D�*;:���\c+��7ܞ
�7��[V���|�>]�����EY��0��B�o<״[mh�2����}})��M7�&݅EfN�xo�/$�:״��zQ��Cu���Zc�zE���m�O��Aw�v]j�g+�*�S�/�W$��᫱��IZ3]�h�Y/��g�ׯ;De5kݎ�/x�X/�l�N�MK/�p����r���a:�(��G!XS�*.7dF�2����V�}6�.�"gz��u�V&!k������MntTh]c�,.ނ&"#�H�u�d����C�.~f~�@��y�|v��M��D���eu�J4��1}	�#���0-���d�-/]����L�����&}�>z�#7�L���.�@>�}� ?Pϋ붮��,�L�{�u���}��|v�	E��uO����ۡ�W^�<����VRi?n~�=�`�G�[r������q�3��Y�Qcz�͹3��ʃ�0�/L�G���ʽ�{�Iu��F�-T�z7�I�������Q#���i�Xn����e`J�d�����cW����2��|�U����?p��bm��|֒	�^�tL�jǾ����'�hxa&Wo���ҚT8e�����Tƪ�������sN���2��{�D���W_rb~��ej�%���Ʋk�0�9Ǒ"�~͝���Ap(m��-:^T;ާiz��W��s**�Y<f+xi\�E^u&��N�S%D��J�Ufn#��X|�W�K��:-a�TW;���5L �i�w<�����Dְ��Hv�j6��>|�t�Aز�K�P)�����1�*,�3����hw����s�gV�M���/�Ϣ��cڹ@ѱ��y�9��z��9��X�<7�.��ϛ�N��?g�jۣ�q�Y�k���<�0N�D�C&kV^U9�#P~���:]x|��2��1�t߅F�={^�r���̞�뇢�&�~����M��a
�*7ѧ�>�G;��ޫ@����%W��H�g�F��ʖ�ga��lRF�H�������܋�el�]��v���!Gl����#������r=ƴe�+������5���c�.z�L�<�=~�Kfo0o�J���t�����t���ׄ�^�	5W��l%�-s1>��j�q�u����}����VƎ��p��x۳GV"����s0k�+�#3a.�/q}^��=�M�;��s,`*��u����<Kچ�L�Z�������δA�O,ڱO٧���5fוu�y�]]E�6�c�ۼ���y�(��	���o~t���+�$��:��=�����+�]���؞�����I��z GT[D �:��N�GG��� ξxF�,��SUɽ5>8o%$��3T[�v���y���P6#�����mz���NtF�t�����g��6��F�\1��'�v�v�+����F��ߏ�����+�wku�6/���3|1�VI���*���zWzx���eU���oMZ{؄��%,o���P��}���M��D�z�u_W����Y-�6�G�}S��Q��ko�`��k�b"A�{Lz&}wf���/�r�b��"��G��"'��-��箺�,>A���t���Uh5|��*����#�m\�;ႋ���b���n�b��j��{ڒU��B#���6��n����i�lH��(bs�=S�`�(��q��S���x ��6sk>3IbO6�A�;��@�����2��s�G�_	���v����4�ރ,���es8���U�D�Q[Ё(y��D�%�Yd[x����/+W���/�c}��x������[�	��b�jc�WԵe�ސ��IY�e@B۴a d�8LC ��:�m�F�c���Z*,;��WjJ��r&%u)��9�{�Y��o �Q��/��eG���E��!��j��_Y�W�:�kn�e���ދ��=�};�vW�/\��`�S��﵀�4%W]lἳ���a}=�G���MI�ndg�2�}L�?���Ϧ�������?eh��ҵ\�{/�kK��[��4��l��.Gr�i�yc�; H�Ї��C�		����2��W���Ȭ�W��,8Jf��}��rR<`�b	���ؗ�+#k�c�V���-sUbw�6������	�)�~��!��>b���7n�z�.�윂,lH��Ĝ��i� �W�yO
��`b[8�s�3����x��؆d�sB���v����k{�}�jd�&���K�z��
o|TŊ�L!ϵ�~�4/��5\Y���s$��g����q�[���rÖ���H�+	j��7���-�b��~���2U�1��hwu���L�BnEe�PSV������_��յ�l��w��t��W��R��R&֪RժSU�D�j���$��T��j�KZ�ɵ|w�z�[VL��^M���5j�-z[m�R��M��Oj�mԭ��[m��UJmm���*KVSm��km���l���)���j����l���)��e6��Km��:�����e-��Mm�S[m�ڪ���e*�����[m���mݹ=uv�m���e-��M��Sm��[m���l���)m��[m��^U��)���[m���l�m�Sm��[m����J֥6�u]��նR��SkU��^���fֶ�J�PD!��̰yo𿷍�c_��yV�>.fw�ۓ>�Y���s}}9i�A�}��������h�����v@:#S�0�����{QAQ_>~W���k2"k���_;�_����?��o�����浵�l��I��IkU)m����J�کR�T�+j���U-fڪmT��e��m���l�km�UTj�ښښ��Դ�j��4����m�[Z���d��?����}��mj�mm��������7����֯v�w�_�g�eEz�3%�kRuY���� ���Vڶ���~�O�y���kmm�ڶ��������w��嶭������yj���}Yn߿�k����ż˷�f�Fￊ�~��s~7��[ն����W�������m
�Ѹr�۞ښs=[�wõ�����m]m�mm�������{���ޱ_�g�$m�`����R�"v0�¡����e}o�Mo㼷�����|_��W��߻[V��z�o7�{��ն�����g_fC�?��e5�	ү�;�� ?�s2}p$q����`( �A�h� D�0Z���@V�`  �*)Mh+j��j��A�
 ʅ5�I�������l�j)j�0��"J���fm�X�)��&Zmkj֨���A[m���wf��e���2̌��Zl�Z��Kk+&�A���m�ff�����͆QVkZ��5�M�l��sl�L���k6�%[bU��Kil�fKiJ��1�-ZUU�X�VZ�iL�%SE�F5�5�Ij�T�u��k-���  ��}�����]��]�{��{^����t=����鳭���n�iJ7�O]�Q�����n��v��v���Mv��v�u�l;:���;޽۽�=���GuR۪[�7OTl6U�T�m��T��   �0��hz>�C�Cy�p��_c#CCB�Co>����4/��ݎ�hy��p�(P�B�w��.��k�ܶ{mO{��-����ޛ��^��weoE7�wu��݁ޮ5'e���w{��ݻCGi�l��I�L�Zڶ��ٕCU�   ���������Onk���vc��ws�o;�z��nwX�5m�嫕׷qճ\�-�����i]<����� +�ݼ{�������=R����U�x�7�9�]�������SU�]v�m����-�   ���ջ�m��ۮ����ܞ˺�v��]��v�X=e���rU����۶��c׽��{��sv����ζ�i{^�������Z�@P��pWM	�Z�km��,��v�\�,S,��   ��V���敪��,Aʹh;��v���=;�k�V�؞��
�͹@���N�t[U@�����P���Ul�����+IbS�>   �Yoae3�Q-;8�P�n�Qv�p�[��nƌp�� hv%�U֍�h�
��ueփ�bn���k2��Z�����m�3�  �{�I��j��T���Z��U�n�������-s�8�Ԙh3emڸ:���q@���@�/Z�mEU����Fթ����  �� �z���J����竀 �4�  ۪�� �� 
y{n(*�ܸ  ���z�TZmV���Qd6m4m�|  �y�� ӆ������=� 7<y�Pz o{m�������� h=��@ <�  �� ��;�  �{ܓZ�%�L���ک�-2b�  	��@ �� ��=g^8 �`)�@Vw��ր]K  �:�
 ={ך� (�� ��i�  �)��J�� E=�LR�� �a "�ѓ)J�ѐ@S�����   jy�*����4 �*DM�T �1?���������n������N}�Ir���*\�!�E��ҲW��P�������z�e���1�cm�m�m����c`���������c6���6>���y����?���[f��6P�U�I{u������ ݷs3C� ���ͫ����� {mu_� :#�J�;5и��B��V,+��Գ( ��E�:�
�:=�
=���8nq���F��s�E��ұ��QD�U�כR�ӷj���rb;������1ł�13fȌ�#gj;�1��C(*�a�Z��fՒ��?�ͱ�e=��i3OQqђ��yVEk�PaJb�uz/-%7�y1�ʒ�' �c�%Dg�1�A�f�j�̄�YuK`�eJ�@�\X�Hԅ��o�,�pY��]�[+d����S0t�Z�n�(�Y*���/M�iC���$���5���b:<�L�gN�ŷln�m`Af�ٮ�GF-6e��Fl1��|f�^ؚ�a�d�&��B�h��c@�sk�6�m�bnku,��t�
`��Z��;�L�(�
�mLkgp9� ��0��dŬ8��;�s-��#x$S+C��]�ل����١Rq^ʹd�l�E�%�2t�����a��YP��,+w%6A��)VR����V��\����޲hi�WfRE�ԩ�R�dҤ��JXǁ*�Kn����z�{��e�1��wKY����Y����ӬYy�����&���� V7*�Ţƽ�ug���G�;)-��k�h�[HIaK��!�0��D���.�ه3wZ����k��巪���G&]��Ӣf΄���m+'T�m��x�\ȮK�Y����ơ�m��.�by&`n�2�zl�%��S����ɹ�K�~&�_��R�hjy���]�t�4�V85e�:�-��|n����t��/_#��"�:��,��v�P%fUֲ����SO.�����V��ѹAn���f��*�}u��b�Z�n��c���8��[�������U�,|�{PL$���Jjܘ�� �Z�˔�Y��:L��4�S�,��rݝ ۻ�A�,����պ���KGZ�@��DԺ۷C,u���],��-h��P=��V�+н	q�����Z���:)�r��Xy��h8wMm���HLۊ���pf%k3wd�O(㱃]�ɕ�w�t����	\�]�f�W;z�jw�� V-W�zs�w�Ye����;V�u�#s7L/wN�vie��B�qc2�3�O�-J���;�VPNIM�-��mA3Q;&={�t2�pY�K�˕����yzM�5��,�����.�r�n�R�'m�(�4��f���m[wi�x�K�D�"�߷-��(yZ7iy��՗an�a:l^�X���+P�F
ۀ9%Z��ߝ�ͭ�Z+S�h v�n2��]ô
5�X�^A#V��	I[i���L,M&7/Q�p�.`{�M�Vٴ���caJ����YI����&sE(F���e�5t���mE3 r�ԋ��۽�:�&nh���K����]��\�{���h�����`�^���K�;�Ri����;���չ�Z)n|,��y��+vc*��Y��*�L�Yn��ȠC��Lgb��f�X�觃]�÷V�B&���c/Cm��I�v���vk�J���&+Hi�^�7�
�m�)3P�Ӂ˭J�2��8��	xpe�ͽ��6�� 5��p�U冚Jf�݇d 	%͎�mk䬪���u���V�V��V+��n���l�l�X����b��H�{,����ŁЊ�EmJ����zlm��΍ߓK#��Է9��d���Ѣ����e���
��|�r]W�����qZ����ԡ5ކ�0��&i9p/�j���� U�7���/V���/S��J�ZT��ٵuegF��\�n����>�n�������0�D���<5ڶ�6٦�)��W^����L�����"���μ�i5Eփ݃�jk㛋YQH�NXtl�m�w�����w���[�1d��m�Wk&d�h��Y0.�坭��t����� ���86��a���J`���Lf��/ ]��/)�f6�X�mX�wy��^��FsՀ���Dlh�E}�T6*i�(A�k��-��,H[[t3㵅�;{��kt�*� �E�7v���b��-�h�w둲�t�s@��V��n]6��D`+m�����bugN�h[�Wg*�����%ڬ�+;���J��QXm�Y׽��7hj�FFP�<+��4Wv��صܴN��Οr��ϓ�U�N�پ�D�*c܇oF*`����yz�z����U��V"΋H����Z[f�wJ����[��஻R���)����⺈oAv�B�LcT-U��T�-o32�5(�
�ca[��·N@Fh9d9jr2�6�@�]�ends4`��րF��c0��n����$��(��ϫsko%mcx�Ӯ9x����Y�p�	N�dP
�d�	�VH)��{Ia��Ӭg2�����eU�X8�0�>KC�v����u�'Tk����!6<F1!;�f�vf빡`�Y����IY�eb:$ei��2��Q�&ۭ��5�YB�:�O��ÔY�2'�����VN�1���`f�3 	��^�P�Z�f �d�
���tV�ɶ�w����v�z�1��J�����+��A�զ�����wafK{�����Qm%[� y���,ӡC��xp�ܨ]���vr�!JR�Z�w.�Y�;v�fe��_m,�S����^h�r���R�y5�iVF��#�'�ͤ�u�b���(��#r,���Ld��p���	)t��tmS���{\���2m�RU`���x7U+1;�vi�N��
��s{I@�A]m�[n��I��{K�5��	'�%�ĩ��R�$͋��yAj��dىҡ��v�˭V ˫L�B�;����R�^�fI@���]،���$��
k�q��$����{�o*:Vݑ�&^ڷ�f�1�Q[�CX�Z��F�ٷ�𔊱���m�1��Ŧ����_B�܇SLMn�N�yxm_au���f&�d��e.7�ڏʠ-��wF]-��o����#��"�Z�+K�˭DԷ�t�.�jn
Y,�=��" �(��R6�j�j!�ҽ�G*ʉءE��h��N��2����ݵ�f�Y�n�n\ۙ��@Vӯ\�b�!��x��b��F4"YhVlL��v+r��D����Z��h���׎�M�����X��L��̡r��H��Rl����N��<��jJSMf��ܡVh��h�Öƚ��Z��������Ѵ/7�x�AJL�V2kU{�]^�
��Շ��j�Y�C�v�"��Wq�F6LoP�[N��
bn�z(��S��qe�I�̉m�"�Ő䣐ǆ�m 
�\?Z��`[� ;4���q+8+jc�BV��.���7M[u�Qnde$3K�ku�L��+����Q���b�f����(���#R��pn�À^�u(�U�Ӎ�&�m��!���{��2R9x0��J��"��x�]�r����:�[�@�WXr��i�J6��ۧ���B�S� :�w�G ���V^lȣX+D#6=�e�@��ej�ծ�8�Xwe�shjf���r�k�
v� ^uve ��ƒׄ�X�u)�۱�Q'������ȬI+���m���&{
Jw5��U���<ZeFk�MU�)�j,e����4�A8.ˌ]��75�)]�,��\oph��ɢo�굖	�:μ���rn��Ҥ�oS�A*M�m^���.��X�8�`	��b�oue:��We?���@6�6(�9X��k�7�TOU<$<I�76�Zݭ��
*XIR�Ě�z�F�2�Nn�����Z�R�Q闋l�b��� �B���A��{���n�ݥ2P�t�4+t�[ZE:-V+ys��Uu.!"�P�J�#]Y�*R`�2�V���-�����5��*k����-�
��l3���XIC�V�k���[l����:Hx�@���xe�5�v� (v#w��L�gX�o�+���i�HY+9i}|m���PU}���)�X-�L���XusU�+{z���d��r���ʻ7-���ԑ*V��Oo/��I�s�r�m�6�VSk�逍��=K���	�F����@����A�h���^S�b:Db[	Of�`f�r^E^�$P��wX4I�w)�kI�.�:-ǯe�-�j�*Z��fЦȤ�㦶�øqP���:��˓)i����nY��4юf
���	���uo�mm�c˙����D
�'��W���7���]�AR���I!Wa�i<ђ=:Hջ�=�Zh�v�i�^�=۰����-�ؐN�ÔІ7**31X���ˢ��hBֱ�C9�(!�/�oq�6!fݍ�q��Z��5�����R�0&�z)J�Rû#r$�	"*j�%DjI�a�`^�m���� 
�J�Wg���T)�4iǉ�Ód�+�d|F1On"5R4,mE4��*�t��P��/�K��mc�t�c$��Wb:�ט�Y�3P���Ygp�9��4��v*��Y9w�n�v�h�,o^�����x�ӡa����(ո�Ժĕc����"F����ʋ�X���ȥ�M�8���q�D�ne��ڜ"-F��o:���H�l�������!4�RX�o���w�o��hUf��mT�d]�۲�f��U�Om�X.��p,�z-&G׺���6�5�Y�o^#�9�,Q�u|�Z�����{j�:�yL B\���G��������w<:���Ҭ�P��z�Y����0���^*0�6��3(P����+�坔 ��	�f��k>��dQ�91h�*����/F�щ�Wo.�S{��n�9C1��a^ص��a��O������Q\��i�Y)�o2�-�u�HXa�IW'.]XRFkQ��o6���i�F��imw&�:O�]��+���:hf�yɸn��ӻ��Ɨ���dYH����x����Mj��B���Ņ ��am��7ko��S.�
�w[¹2�k�|���e1L5����n��)	��KV�n���{Y*2�#�c 'l�\�-\)LD��(R���Iǭ�`E���)Qhg�v^�l��/q�IY�{��%�Xt�j�9�I����X�b�qh��;�iP�@+��ojT�7F�kX�͊7J�n��Fk`BV�t3j$0���â�V��j�����=%!6m�ti.�m�ܹkU��)-�U��U�JL����+D��3���-�z]��)|U:�2мH�V�����Zv>�K7(�L�t�֮H�̼�я*���e�:q���&��k��5(��T+.�h;&�i��@Р �.�K�i��0#�����ҰCv,ӇM�H��
[�E�u��"�nQ�WydSnM�0�fE����@Z�O0�*)��h6.LKk)֨ɂ�::�X��G�&i��{�^�PT�8Y��!0Jm�j2�fÉv]����˾dB�I�ύ�e#L�G�Sm��*^������e'G2�:1�X;��Iwg5��۫Ժ�t�-kJMw�aq��0��жKs�ɭG�˓`�!X
�ɴ�j�*��w,��DZ�3N��l"�4m,Q;��yJ��W&�N�%Yt�-[�� O+JD�Qb����8��cz����b���/bĨ$��� T�i�GH�n��أ�1�&6�ݥ���u����c�z��ʼ�Mg��T%ͼ`ƶ�0��m�Y�r�߮ ���ZST���YoC�j15�ԩ-��&��X��T<A�U�݊�ad`ҏ3��b�e�u�R��?I
�VTlm<.ĦQ�"Yk�m�<�cV�
�Ц��E��A��Wmee��),�}���wLpy���� qaݛE[(���(�P(��5=�7��pemҎlk�Ifmn�
�:x�.I!��՜�����U�g 	W݂�]il]寍;U5,���,T�6��,U�g#�)���X�J�C\�ࢍ[|�˚/m��$�aW�If�yE+>�q�jem1�6-,7��-�i���{g��',]z�K)�+�&��*X>)�;��|��N�.��%��h��+���ݧ����y��+4RL�hr�G���� lU�Vf�v��)f�2}l1�)�?���J��,U��*��.4{�.�0uڮ���j�O�!�mf汉���Ύ���l2e��R��B�/7cҦ�U�0����i%J�:�u�)(�ze��i���&����p7ȶ�i��R�q�禈���m��@�W��R��X��ོ�v��RQѫj'WlS;x/fi8�ukf�Y��,�m�F]Jr)c��j��t�-��Ź+�F�PBPdb7��c�62V�j�l�y��!�le�X��yvn9 ���1A�ʨD�Snŕ�@=����rL��<�x,v��u��Kᄓ�-*�w-b���qPQ��sv�̊�Ct��9�Z���ܡX�L4�+^YQ]<��#{�%ڄ=�L=��aj�J�|�[�m���۫��<�75ikYX�I�̆�L�[!WuV�;���]]*�
rR�Bͼ������r�K����l���٢��J�.`�6��k�
�J�I̺�t&Æ�0e�IF� ܣ��K�|�S�F�ViB-HU�AY
����Gv���>0�� �jdt3��E�e��:�Ԧ�7f�n-%�1f+���ںj�$Ϡ��k�o*�%r/��TĶ�k�y���a?uu��$�%aXw�lN�-�����Fe������5fT�&E33Ճt��(�#T�Az��Us^ڼ1%�V�b�IY���
�v<��(\�I;�CZ/3-���O5"q���]�wx�!x�U��+%�V�K����B�%�[�M#.d���-��w&��t�j�R��j9q�FU��u��I�we#h�7���Y}yN��]�r�ZJ^��\x/0�b��,4B'&@������WA�Ţk;�	V�$_^� ,g2��\���I+4��]Q�ˇ`��kim��a���ڐUuzg
�`ȓ�L�vV���VB�����&�8-Cx��f����9�w)9:J+�-(�l$05� Z����g����]�9�eBI�ݷ �qk�M�6Jq^.2rqT\��Vq��H�Ե�k5���<�ؙ�CIˌn�Me�x^�Ա;W׆тid	�W��#[O8�Z��*�͗#�7���+Fͳ�+ŝ���tV�ݙ��C9 �7�
P�Eˡ�ش�b�M9�5U�j��T�'�fG؂oԤ�|A{wLdC��Ƌ�,�ǭ���
���)Z�	��(�QVT�bi
V���4z�D^G�B�h2SSeں�@�U�	��4�ɮ䕿b{�0grwZ�4�g]Z��/m��1����
�7�r�]|�'�b��Vx���EX�ֲ1����8Y��7;��suB�kqB���U�H��&'�)L�l�i�m\������VƗ����ۂ=7��"i-C��m�КI�O��%0`��G��4/os!1W+�Ւ�4O=� I[՘�Z�(-��|��{M�7$�z5�h)���2�=ﴙ��{�"LȨ��ˎ	�s������C���Θ�Z5l������ނ��]snUn!�h�qXR�*c@���LF/��Y�� ͻ�A�	�h�r@4�E���>x�TDZ+�L��I�(V��?+�Z�@آ��k�kd�Y�e:�K��*��^c�E�5�[N�"�K��S8�����\��Ҏ���F�oqծ�l�G�瞤�f��\�en6J�6�eלӏ4q�0S��Cb�B����{A�Ѥ"̤��� ����u3�&Z��ӾكZ]��dbޚ�T��,��P��+�m� '%��ʝ��J�����{rޚ�}�ItTooRu���:��k��J��VK���fm5A,�IP���g(��5Z�Y8�sM�{0@`Z [J_[+�6�'(N��(�(�¢{k,82t�)W�Vv�ʺ�N�d
�f�*2/��r��=�gQ��u�����7Zr��E�I�W:^�Cy���d֟}�I��S,����;$)�vm�}Y"�/t*P��������a�K�®0 �R���-nr�8U�t��Y�up#��re�,p���(�Ӷ��Zvj�?�.�%��N���w�;]��W�	5�x�e�!t�`��>���Sw#d�&:�m^�r������&�T+3�Wl'���en�V�;.�m�N�fn�
�r�.J�����ܘ۲㔭�ź��eVGjj�sj��NT6�S��ά�@A�;��)ͻ��l�;
'2��X�o�u�|֎j��j`������r&ޅ��xZ�W啡��y�n����y�:�o�S�;LK7RԷ�J2�������VX�N��,�!IF���W2�Al�o$�$'���K��l0�;�X/�Q.m���IӪV��H�
�/7-���1��00�%lux�
q��N��N1��J�a��R���H�>'�N!*��-|�b����j�����V�8��9��x+F���V�6�r�L���M�T�w���\Э7]�m�qknz�^M��6��]p�u��	!WZ{�rf�R�I��ʻ�0Z�r�6�{�`����S�jNk9�ú��dѤ��e����qR��Fs��T�=��sw��v�\YM�˫f�Ir�^Q���b��8�S�r|񮸔ng��*�j��e�-�K/8�'���ǉ91=�oj��j�t�"mY۸� �����1�<�֍�Um�Ԉ�̭�f>E�[���sDC섖�{}�ތ}�R����Ϭ��m�� �� ���u&���R6S(.9�jl��o[�{Ҳ�$|�h�L�k�(�[I�N+�H`]d1`G��R��w��t���S-cT�r��J�n�:	!��Ӊn�)�:w+��ۡWo&dDoe��]I0k�D��j-�R+C/��ʵ�+�$ˈ'�;)�Hju���h�;ׇ���tx/��V��Wo�3
�ZK`=ӫ��m֨\�'r&�[�0jg�`����ۊZDPH5�t�ؙwŘNGXF�i<�i�շ:Fp�b�Dڛţ���%�=���q\ϕ��n����n�ـ�5w�w �E̖T��g(Fh֕%[.�G/O̡���1�����R�D��ͬݽԊ�l�]ُ���D�\z̃�5���h��E���="�,�A��7\���ƹ�P�VX��^\8�=Ω+F��h�0����uj�8��=g�{T�l����C��ٔ�ٙ��-�H���O&�`a	�wKY�{2���w�d�W��'�H-��(�^թ�kg:�X�ڼ��6;H�;y uw�P�����m�.]g8g\')Vaq �3�;��{X�S�k�6�om�.��DG hk���u� e��s9@@T$��6;���Oz��� ��4=��\��ndn�M��p�Y%c��
P򝝭�}�*F��z��om6�n�*�|�=�`�ZT�0浥oR�Djtl52��y��]^!��j��n�t�;k;�� ���� jh��ҫ��tczA�C����8"���_Z���ԒO;Z�7Pk��0C��:"�p+�ð������:�;�����#c�ܫ�RD4>���^���	jthöڳzR�Ö6�S��x��6�q`��rN7�c�IJۤ�!�M���rn�>s3:��۩��J�i�RFK�~�V,��܃��gi�y�Sk�Q����N��7;P�om낄�%#R��mn;��^R�ڝM_gS},-%� rjѕ�5F®����=�H,rI�������c�/�q��mk�cn\��Z��Y55@]����{�̘��U�]��#��P��-<7:�/��j'`�J�n�-���J��9�����4��Ŵz�m��)�]��8��Vw1R�|��>�(:KZ�d�*d���X�����՘�曌gbq�=�{
����Z���+��gY�ހY���㋣W���O1J+5y��{�j��\��m�q�e�=��V�����a�\4�EN�e�NEa�;K	��V����!��	0�Xp_fev���B��v�hb�,E��j.��Զ�\Oj��*��~6����o[�1%��e[�2�9���]����v�/;¯7��D��Kw�^:�S�,}r�j�ᐧN��wq2����[�ٛ�3m�k�M����Dk:��_]�
�����b�V��J��.�29M^��\��m,ڜ�,2�������ʲ˙s�$n$��S+(}�'GR&n;3X,��ʷKonY��f]�YB���I�D%���}|���wɭ�m��� ۧ�p�X�Ǳ�Sv�c�AƦ�t.i�.�S�6#����]�^��[oN`�R��'�r�[G)b���V6�#��h��D��Lf�jWqM{n��8�޵���܁�u�U}��R�K�M���hN�4��k�����=�{~��[����p�[��r\~�r�A�-e�4��֢��dn��˛:�T�_F�L���@�Zɜ���ĝ�bU�P%�ohN�]�kg�lvI��Vt����k�z���7��f��C:�$�����n�m䗖�c����yW��*me�I�V#s����&��˒ы ������A��� 7E����ڵ|�K��ɏ"o'ml �֮"����m��qӕ�W�^ܮ�V��sm�.���� ڢF��K�4���A~laT���&U�ygf���e/l�*��Dڐ�/A�]�Õ��^`vԮa����x�c^kF=j�V�b��YS8Z��'3X�]jQ;�x�$r�K�#52�T��fa<��z=�0m����F�,n����H�'5�<qq�R�H�7�X�9�����&�X��sEK���W@I�Q�8s�%��ʒ&�L�k8z�.��W��*�X�$�u�-��em%��T�Mp:%��u�T�[&�+�!C]���Ԩ�QR�q����}�}o��]z�%iH詭M�v8����v�{ӝ�`�����9n���8>@�j1X�T��/���~��ׄ�*�.ZQ�.��ݭ�}�\��P���]�yš1*�J�,�9!�śq곦]o��`�m�\�n1W���kw ���d���,���%7`�>[Z���Ҭ
�Pɟa�o�K�󌷗���;��nH�G�⅍<8�M��[�,:e�� `�  �rq��e��Z��VOuk�4$Y�0�d�#�E�O;��pjV��0ma��Z���Tˇc�YZ1i�T)�![������V#EnU�ڠ"�wU��`r�k �B�-m�ה�G�N����^f�Q����x�]s��Y��/�J��ۂ#�.���!����v��Kj�ת����u�7��Ж�%��/@8!�؅��T_`�:��|#{��pw����@w���Cv�'�a�[�9A��ccNlp"+U�W25WP�}��KΈ���;+i�A�W�,�:�we�%tT-i�C5ǔ�@Lk����o�g��EU�A@��<��lUw�]W�m,�]y2H�U�_�Ŝ�˽��n�ԧj�iE�X�]a�d�)���k]]Υ�
UW�
�N7�Lvn'6Q�Q��2]%�E�D^�J�"�]+�Y�����\�K뭡�ilBv��P��������WҎr��Ҭ��p�rIȭܫ� T�Y�u\VK4�J��ѻj��z��u�K��i%gf���ƀ� �k�\\��h�H�N�'_�8k�u��<b-�sf��h�'&�`UJ�c���sn�ȱ�啲v*�gwXV��P�\����q#�P�m�U�zU#��钶����i��c+20������Z�۞��a�+�c�T���u����3�<����6m��}��[h�R3�K��<��f^��3�� yg�W:J������̕9V=8-Yů:X�bhI/��L�.�?{6N�L[wg�طjsz'��ց�I��9�QqX�Á(D�f]��S*��l	}��t�^��2��vR[Z���[���/9>�|����6����GuLM�#�Ӻ�RR�T��{�N���kF�-�ju�I�uݔsPՀ��5����yJS� ��9�?s�����m8�y��BF�IFiޣ�Z�݂u�� f �j����o�Q�ʟID��[N���J:�O�nZ�.�mi�%�X��],��N�oj૾|���Skr��,��k��H�B�ջ�Ң�Q*�Me��.�o�׃��T���ffA���я�-e��KYsu�B��n�T��կ��?K�P�Ń��{7�\�d��I�����.)G9W,�����ߗ^�82��j�Z0ٕ/��6���zKT�)��j#`Y�B.��R�r&�|cxU݌L�^�dڽiR��]��wMr�����I���ͬ�U��buZKf,���˲+{�XvN9�*�Ø݄�m�gb�ܛ;�Ŋ�+L�<Ay���1ǫLZ�m�]�)�ׇv�\MfKR�|hN7�m���*�+(t�cJ���w.��k����2�����w#~vIg��k)s��s��OF G��nо��h�;:FV.��Y�`j����a��JC.Y�Qv-�ΖS�qQ>�Փ���,�71c8�M�kM9:�]Hμ��ou��Z]���Yȧ��˚�	�����*����C����-;�]St�%��"���
��|��6kw�wQ[1���U���s�a�˨������{�;*�n!�J`�b[K�;5��a����lKW��p��7l�,ܾB�,Җv�Vcs��]�ۑN��ƀ���� ��2����]����˝�qu+Sr�f�����m�չ�.���#(�M�X�cV\@�]n�%K�F�`�ֱ�J�PP}M�ŵ�z<ɚH౫�w؍kXRɯGY�\4r&�(��un�0A&I=����!Ҙ���e:%ݑuYx�m��(�3��\��`�;I�g+��رٔ�e]/.�f�tiVb��-=�w�Z�XM�p7��vn�#�KP�S-#D˩�}��Jp�l�ܭTT-�Vk��u��V���;��]@����K�,��ܛm1}/V�F]aܑ�΂����F�c.8K�M�u��#�J�H+r��aݖ�v8)��@wz&��a�tp:;p�6�6Ѭ3esՁaxQ���Zq������j��q	���'�<���y�qQU6��b$K�nZ��.t���e:�ݮ�:�=7��h�s�ҕp���iC�"�v6�M�)��D}LY��jW-����&f�Z��@Y�^���Ph��� Vr���`���ѻQ���s:�54��:f�����1��0^�K�TG&��H$S�L����jɎ,��Ɩ3w@އr��݋SB�)� pQ��/�;34���s�����c�FkS�������c3Q��\���V:x �����.Q�t��B���tcR�	a��_c2��#w-M�32Z�k(��:�9T��g4}�hd�L�]�YR��Ws�X��h0_^ڷov�L�
�y.�qWu
a�Oe	d+˽ć@�ԅ�{qô�;`���s����P�Q'�W�s���7��z���ݎ*�VN�@�.t�K�S#a��K˘C�C�V3L�BNk2+��0��jn��{/)3�IwM���E�;��o�\�F�1J̑�,J�$2δ���8��Ú�U�ODK�u���]�Q"�q������8Eԣ<����B,���:�W�Ճ����QJӴ���T����\������L$�Y�<�c�׮��j�����MĶLR�vr�X��)�ڐ����MraJQJ՚��b̲f�Έ�����ӑbổ֓�gF�Ir:���Ak;�Iw��C$�9;���|����߿��6���,c`��Ͼ>|���s�+�'���K�m\�kd\�w�*������lX��q<��sir��� nv�L�w[����Ql�u����Ħ�l��f���f�6sK��2l�Z�&����X֮ #�=�VWڦ��!KG;fj����1�R�ٛ	L��x�.qօ���\��@�%rT�rƂ���l�z�Oskle
<��mv�3WC)��X�0;��z���J;C>� ob8��'ua}qv����]��a[�� �[&��Tbݢ/f�⒣����mJ+0ST��֘ �؝i�j�M�VI2Ν�3n�7(i��sm�E���Ԧ�!Ś��ݙ��{-�8�F���?Z�h����w�+(Ƞsz��qۿ< ͖u*�nD��!]�9])�nL��BN]�B���F��Kޠs��KX��>}@�Z���ˬ�|�$w�c�*�Z6.aZ��vYX�#�H�i����� cǔq���B��K�c@�;��KZxL��NV
<o�����H��irW.�7��sf��r!OJ��q9m������{Wj�MU�ܗ[{9>�4ros1��B��aW�5.�$&�6��`�2J�㕆��n-��(��-Zl��̫a��L���9rV=���PF�9�9�kݥj��Tᬥ�
�{$8���@3��G*|������jӰ�Q�"쑒�s3R�Z3QdV�j�&�V޲���f�5y�q&f�ڝE�W϶�T���������o���Rr�qJ��ͼ�n���$��cc �ًC�]ԂX���'d��5V�͡ҟ��j�Q�	/�:�l�PU�G��-Nͻ T���Bs;��J���Lf��fU U�Ki�3d�Щ��Ղg7��u�6|�r�R��@�y��2v n�ǈ�q�.�Z��f��r,"��5��7	����wH�̸@Ic�TT�(\������ȴ݃zx*��ww�G���)0�9�6�wL�-f,���m�U�8ѹ�eN$�s�kr�ٙڍ�7�y8S�tN]���k���yM��sjVDގ�Z�X�ї���1ة�����n�=��57A�s1V��4��$�3�t��8���4u�N�U%��B<��5��'x7�B�68�{K�ʼCE�&�o��T�t6���kzd]�|͡���4��:�ə��G������ݸ����F�K�ͫ�yCj�PV�u�O���f��fZ�p��5w�`�g����Je���-��r��DX�]ժ�a�WF�}�u�ъ��-��\��
Wq���I)څaܲ�^C�8h�E9�P��m�լȴͱ��ƩY���3Z��2��^4)\\����X
��Rú=�۴���ʆ��Z�J*v6XlVt���$�X������/*�E�k3�u���-�q��e�ɕt�������Á 7�jn�Z��r�u�3��V���0B�V����P�tfB���Q%��WMEZ��,M�Ӽٙޘ;2�EY#�u��C)XE[>H�_w��j�AH�GbO����3Ќ �ZH1�ƫT��ǹ��7DګU�Bm���O�T�nuY��1��7b��0�q/M9���4�:0�X5]�w��R�g;�٨� ��۳(�W��>G��M���nDCCJ޻×�=X��q@�Tw/,JP�۸y���褄ʶ�Sq�|�Ѵ4=�B��*3��Fiq9]f�l���m%�3�,e�p]��h��S���%�����U���,Ʃ4�eL:�Ma�pf�Ah������nw)j��rh�ˮ­����=9"QJ1�s�ƥ�+^��b�/�r�x���S���?1�B69h"��m��YN����͂�[�ycU�3I;jTG*�"�����Z�dm7�,���Ԩ����;��[9��:��
5�����\�o/�K:IL��7JV�N��t;vM��6�Er=b�+Yf��t�Ss�U3a��ozR�pV]�0X-YQvS��`cxsv�����:0GBPF���6��H���C�Q��:�����e�ШK�u����|���҂�WZ������z]c������Y%L��:f�
�Ww�6�� ��峤��U�>�\��$L�&�FL�z�#�-���T�L�b�3D�1�
��-�ǻ,r9�j�MP)��8/J��-�v�M�譫����ٱHP�@%i�4x]�Wg:�JSi��� �Z:�b�ؓ��;��ֺ������I,F���sǋ&L�]30��y6-[�(�NgyR8.�Y`�f=Ȧa��,�����f��*��t��g3$�-k\g�T��v���j��޻ܦ�c|o���a��ȥ�QU̬;XT�R�8��X�gy+]Szm���߻h��ԭF��ćUо�����fR(����ˡ�h�M㥮�p�&�	[���q1D͘�;ywB��QP.��w�h�s�+.���쨍�դ��Κ
��c��P�/9�E�Hd�Cu5CJo+&���Y%;=Mr�ܢcӅ�5��ܗN�R�^n�R�K��G۹X]�&h�k����-���h*quD��ڱ�1W:�-m^ٜ��Х�E���'wk��Q�\GQN�\��zij�7�'���������BK��%�p�آ7օ8�K7*EqIcV:[��]-Yܻ��ۑ-X^ˆ�MB��-�W�IݹI�n�!mѳ��oƎk6�sӦl]G�Ҩ)V�҂s�1��z7�t��~�3^v,�^-���\o�"�q��4��،�Y�Zw���懲c���X��ɖ��j�L�]��K��j� ��.Z'6���e��|嵘V��pM9���U�q�ݕ��Po�h�f�z���
.�u�zaHҥZ�Xܤ2d��^�t�@�{'p⨕[g2Y�D�.:+�	|�.e��N�ƶ�nJ��!�������5�����Г����v���B�1��t�0v�-j�إO�%�Y��C�Ֆz(���Z,Y�%w4f�{So(V5�R�an��a��ͬ�h�-��4ӵ�VY28��>�T���V�xf0�n�ȫz�4�	�Ū���^=��C��`ge����<�yJJHrwj�WPjN31V�����+�"e���-��;�m��9Ds7@A#�"d��t^;Zxo�Pw{7O<˶��k��YC4�R�7��}*d�V�`[�;k`3w�6���k�VهOD��8���y��ۚ�7v5����v�=�
�0F�T�oع��GN�4���s�t[��3��ۂ����bΥ�a��d��*�w��_B����]r^�w!5�t��kN�<ծ�V�-�5Q�d�̾]�%�RE�� ��d�֑��\�+����nzE��=�O���I+>��P��5kwJ[cA�	�7c�E"6"��X7�̣�#V�#����lM���"�anb_�wI�>�Bt6[��l�ك.��s!涭���HۧB�c�9ݮ�
Qf��w��X�2�̹>|e��1����k���)�,J#*����r`7-$!�)�Fe�v���G�X�m(v���6lx�]��lj/`j�v%��+0���n�=�!���8�HTڴEVS8��f���諹R�����N�g6��J��A�u��7^!�h0$�Y�!ֲZ��%)'У�X�=#�Dj ��sS��⾕m__ �6�:�tu�Nj�YR���r�ڽ�jN��^�D��'mo�u����+�/U��VuW-.���cq*�"�:ڥ �m-t,^@]
�	/����.W�c)�Ӎ�2���Ź�u)��n��]�΁�3CT�d|�u�W����ں8�bYB��^��v��c�F�$�[��lu1��2��{�<��*k&� ��Q�Q5������m>V.���رbU��W��iCS��5U�شʀ��u����}�D�8S�j��M�t��H��/ji��X�|�8EQZv��r[ODۗ��m�H�_B��n�Zx�`�f�H\���²��U�*����۝3D/D�J�33Q�1�f��I�^�I{w��)Ӣr���L�p��宀�/��.��4���m�:�oU*2DU�j�j�[[S�i\���Ǖ�5q24�09�
�&ĺg
�\z��ccdC{�I:���㣲������@�fs_v����D�����H��;��c�u1Mi+i��3R�]&�a��tp�M�M�h�B���ֲiI��REYu�1w21�/nf��wKĭ�$��s�d�0[�`F*p̓�W`�Sh�̺�X�F/d�aR�:�;o����74�h�����NekslQZ�TCn�fr�K�;bM��St�\�[Wot��Ճ0i�z&���U�J�a2T�+ ���[�u��ZZ��75f��Nbͮ�+ ��=��ʜ���%��S��mՁ���u�P�ڏ���Qw��+�>Q���{Q��Y�"<zIwiG��"��L�V�j��!�hi�M#[�	fRydC�.��&D�_FT0V��˛�95��(�Ӻ���G�>W)hI�W��!;]@�v.��	}a��eKZ��l�x
��@i*ߛA��W�t�����f;á�y���ܒw%R�gr1W>�]�}X�֞eV}x	�n�-砛��P�AhT0h�7�Yc ���Nc6.㚮�o�ҝ�4��X�a�:�	O�G܂��hЮ���+�ݹ�>C�Ĳ�ơzD�S�iA��WAl�3s��Ԟvފ�R�G
�U�Zo�n�kw��8��I��ޕ۷�m���̎"C�Ycr�C�伫��p�/�r��ݱ��x�W2�	���N8�k��5���ۺo3.�hrF��a����/n�E q굏���Tc��ް�eS�o]�T56s��J�o��Egb���N�b�u`�r��,���4V��AVա� "��Ke�5+r�k��)�X�I���s4>؞޵�{%�q0�Y8�9X��Q� �\���U[9/+n����*�4��S{�}�$�B\а��
F����\KN�|��W�r$�bs��t2�;[.b5��I�b���Z��]�7˲�Ҷ�ܿ�����(V��(G��a��C�u��^(T�Y����
�iS؆k���i>�6��F:4���P�K��B{�/��OPӺҕ�s&..�ޥ���%�Ĭ�El�q_`o9�����0��@�"˼�M�U�d�(�c�Y�/�+J�.���2�L�0�.{����èJ���i�te�e��1���XGf<Ӥ�c��
n�e#��[��T���N�#���q�&�ޢ��l�nE�����Ǆ���e�鶀ٶy"ڌF�C�+�A��h�WV�T]V�=0V7u�V���$����PΑ.4\5���l�ѻx�̅�\Ǐ�fvO�7�Q��Nc/U��Rұ�i�fֹS4�]���o��P�<t3%�n��I!t��<E���c�o�ծXѮ�z�J���i�v;� B<<�=�-����ia����<\e�(��9�讲��LU�4���T���\��)I�����.�&]hՉ���U����8(]���}i�6YV�v���dՐܖ�w��z9�v��f��Ia��j@�H[����`2�fs@Ү0��_]�[��{q�QT�bw��ܘ�˳CI�o���-_i@�����k�oo	��e���m�m�8�����]X�ҟg]N{�4wc��ʅ��V��ťƚ���v:�1cAE��[�wכj�Azq6�3a_iyx�BT�˺��uyf�ʹ[ޠ�W2�µj�9#��ZI}�>YE�z�6k �Vm@$��p�6+��J�I��	n��O;���0�w�5���KJ�����,�%e;�u��iÈl�5�f�I
J8��2o${^c�{ir�z�lK,6����hα�zM^[�I��l�
�]��+��1���Fh���=�hLGv�'"I�8�-VWW �oM�A6�ŻI��3/o�x��������]+i�a��+Q�Br��6���,E��j�+e%�fX��{�c�r�F��a,�98���p��n˷,�[L�P���C����\8Y��sw���0�^=j�c뽗҄��5&��Y���ٷV������r�Dݔ�P��;�R��e���;��0ŁZ�+s������A��wI�.�k>Ԏ���q�1�!�V��Ἒ{�b_�4�B��0����=�n���������
�;�����$�����Z�X�h�b�f�zU\���}��e�[v���Vk.����JN�B�S�:K���i���p�X+kp9kS�6�K��ͩ�fn�y@��1Q�V[�%���m-���)T�(+b�ʛ�:�k؞�Q[�3Yw�.N]�ɸvn�]�Zԍʽ�7�Vޱ+v1�a��*�f]�)Y�
}}�4� ir7jظa���޽)��i�x+uw��vʵ1�v��E[|,J�#ʰ��n3��!t��fP��q�r�\̈́�쳒������+�B-��ϥFH�p�]<��s�j�U��fp�g2"41򸻶����Vz,n���X���p	l��!���h�]�	��6��z�EN�]�:�uv��=ώs`3+��0���F�dBm���.(���]�6{�h�&�cEV��\#-�K-Щ���a��K�R��A`���0�C�5w�o!�ӳ�²f_\�'M�����dwru��<]��_]4b6k�n�{����E���g[;���בoU���Rt䳫;Yn����uZc��d;�U��b:�L��V��V3o���f�S����S�{��o)�x��tk\��������)�	�T��b�vh5WO�k��Qh�Ǡ���K7^��zDp�1ֻ�jr?��������a�|����x"*�o��<كZ���;Og��c,1��`�[�Q���Sg'{�8�Y�4����90L�89N�*�}A��q�KMv�ZգiF���Y� �顷�4�b��Jm�������m��#�:�`�41�e@��6'�m{�� ��M��.���nXo(ŐtM�r�WT��
�����\н���YM+����}��'bu���	u�J���g�����#����a8;d��͓��؜��;1����LN^�Z�5�nT}��C x JWN�Z����W�)�dws���P����M^ń�+��Х��ö{�Ȓ�;:ij*][��/ckK`X��I���C�:� 3 q��׎]*R���Ž�)\|^2�<�˭�uڷK���I�ײv\ֈ|�V�j�4b�|$��`;K�1*�Ζea+-rg@�[��F'G��K��V^q�JjtS�C����B7��9�G��W@��%�[�6��z�Rf�M�NG�;'w�R����O���O
���0�2^U��x�0��_��Lx�on���ys�Qk�mQx�V��;8��u��:G��K̅)�F�m�����Z����m��VEN:�+{lnu`k6m��М�	Or����*��Φ͍�q�U4*m���9�f���B%���&$�v�8�^]�1�V7�2�RJ�U��@R�#����NDl�9@�L��y�9(���N$�N$Q܉�#�TQC�iG#�"���Ur�9Pr0Ȉ�"��"��ʊ9ʨ�r�L���Q��+D��E�"��eQDE�TA9�p�2�ʮEDw+�
�(<BQȨ�(�Z	�\�W�ePQ�)fE˳�r����J�#�<t�E�r���)f�ghd���-H-G+��(�"*���(�QE(�t�*ԸE+X�u�D��pyi�(.E^���Er��ÔfF�p���T�Y�fYZ�"��p�%ʈ�����DuB�̢���#X��ӥ�J�fEvP	�@EB�}�}�{y.Sw�EsH�^��c�F�X`�b`_W�W�q��|9'��˽�F-�ZQ�݊�&'��Сq�w���].��7�.��X���;*�b!h�k6�4k���^�f�g��k�	����cH֓�8;�2R񍆖�+υ���q�l*g$�]t��~���+PY�Ѿ�$.�qÛ�qz�m����l==�eѮ������U��v�D�u74���UeK]����5��+�z���~5���Cj
6߱4����,%4D	w�u�}��*���ւ�.�3y�l9t��wZ�'W=݇��'�U�Y�`�zS;kNx{�s��늗0��y��7�n�T�N˙���S�ϥ�64����g�+�w�;x�¼��;ԟ]�<;1+�bMҏQ�%�
�����s)o�^d����'-�'���5Q(�-�cIs�VJ ٶ7>�{���V�'K��/��j��]EH����1��	{��\��vƢ��
Y�!�x�C^���kDtPp$�%�W�T��u�?E�<.BZ�k$���1�ھ]�$)�N26�a����=x����ǯ�l]T����]�ϭS�p����X���%M��N�5�b�6�sV�ur�\:�ӱ�!��T��`�WL��UY��W�ZV��� ���VZĹK��X�k��:�[�N_%7D7Ӏ�1S�8&�Κ�PS����c,w3�)i��Ǵ���Y��Kޭf��E<�H��>q������-�9<W<H'G,^c��΃G�������^Jt�/���]x۪E�tBf.;2g~��}���l'd������:*�������-ș*�5f�|r��������N�Lٗ�d��@M�N5�ֹ�ۼ�|�^���/��U����zOJ�6���`7^� g��Re{��x�Hc����s{�6o�5���W7ȧ�w�1|;V�X�:��H�&���l$(o\奣��i��76���Bn�K׹�2L5�)���m�?JK���oh���7��M�/��<܅���F���F{R<�U���7����Z���h���Ϧ��9�c�J׫2��x��N^D���
�v5ja3_֛�~9�Q|�vK���w��o����INpQ�U�^��ب�®�)����p��9��N���\��j8�mR}!��L��Is�@��R'r����ݲ�as��Q�E.�=�^ *���C:�{č�`V@��s3�=��s��ت�5�%k�퓘s�*:���U���zs�j R��P7�Rga�e8l��,C.p㶺CԷ���j�9�!�n���=�\7O:��7J�=������W�1U�+hsfO�7�N��v�s�M0���Kv4�9�9�·�vz���ti�W�Vv
���+]K��n���q�.�
�	�zG�Ϲ�`h�0�;�����y�
�Z8.�iQ0z��ٶߚ��+y��R�/{�%�K(��ŭ��o����N�>��﫫�Db��Z�K�GHS"fq�\���8�z/���2���_��t�,�����<s�s�jwC�C���^��W���A7@�T;S�9fW�J�1Jf'Q����CC!v\S�oL��*s��^�B69����924�f]�9B���Ǧ�ң�.~��)����$��P���f�;���#��ݪ��Z��ɸ'`����ʻ[Q�	�G��8R���Əs�t��ȊLtc>��X�!O��5�9�=TY����ʮsd�qD(��%��)��Q4��0TG����w5�n��YJ.�vo���c�3r :�O�� �>I�U�z�G���}����.b�2.�R���\B��y?"�K`�P�I<2��x�&k��,��=�� Є��,�a�f�en\�`�JZɒ��X�r>Kѫ���H���WՖN=k���^3�H{�G+�ܟ(�}����D������2j;�Π��&Dø����ө���n�e��ԇ34��Ĺ�bTY*�����ڷk+RUn��:5�~>�"���i_-��5
�󌟥����=c�w�����Y��6�l���ݎbՋ	�ኤ��O̯<ÕR�
�϶[���v��v�1s�b�Ti�J*f�͹<�JJT���4��!X!7�bx������/+�j���i"Ϯ�{��d�m�eWmՊF���!��\V�89�Q��8i�YT,V7�KS�<A{S��&�.p6X%4F"Q������feû,07��;>Mg�>5�.&ٲ���K�:	}+|$�B-��}�����z���7%V��+#�C�����l3��j��]Ʀ�+P6۩u�e������PӖ/=���N�\t]����r�؞w��8;�g:s:l��e�CXŞ�������A�c�U���8�����~X.��˛��>��ϗ�+�ǽ�q䨇�r�x�&lM�ao����;F�5>��N|�{�2k�R�v��^�ؽ)��[����tr����n�",�޷$�U��r���-q =�x#ʼ)��ݩ���W�b�+QU(�m#�n0�r�ލ���I�tVӻwo,>Z�#�7@�J��ڨh屼*���"U���zz?Vp��l�fEk!U�*~�+9��\S9Jj�%�=��\�'����A��Qh��<.TU6a8%C�]�R��.���@Obk�Q]����ا�WJc�rx&&cN7�g���HJ�uK̅K�� �o�۵O�e���;S��c�3��/Y�$'m����:��M��wlTڪ	V@k���,��b�JoC��g��~���C쫗��9��
r���G�؀�������AUL�yVֈY-�=�Y�Etl�D�g�-�O�tyWk�Һ����5�.r%���V�{�K�2X�'��b�57�s��V}�� L8c@�Rxg����H�p�ʇ=Y���yn[5v��Tk���w�4����
Y����v�^Zoo�}x��:���Xm����9 hqU*e���V%m���S�0p��y���(m����ObYf�W�6�J���`s�j%��˵L�.��7���c �,�C���asY�G�8t (�S��.|g�M���QdiM�z�)����v�}�4�rZ��ֶ���׮����{M��N����$��Z��z�JH#uv��2���A��g����̹��s5^*w��ӎ�ڲ���=}������8C����w�(�$��ʌP�����Vm�bD	��f����~g#�4f!��I�=tˋ+,��j���i:r�󻥌�vM��1��T�mɉ�4v�QW\%-�9��+l�N�:<�Kh9�]�B�d�u��^!�&7c����� �CҜ��sv�̃�G���3�wj�����ͻ�����F����E�"񏈩Y�^�'����GpVZX �+)��˫^$�h�
�}��=A�n�<Qc����[��S%Q۬�Cg�'k�lFC�n{b��5uN����u���¼:ʽ�9�}|\Ζ�� ps�.j�x�-]������mi)i�*��:<a%3ϝ��OI�<	�e��!]#�|�]���.`��A\�!���9���B��W� �dc�u�z������ru��c!#Y���������pA������y�瓮���8I�
���E,���к�*��z�4�|Q;�bB�oN��Pe�.9g,�=6SX�~�g/���j�a���S�,�@n���f��נ���d#OJ������X�jFL��7�(xꊵ�Y�ʮ���zԇ�߀/�����S���U;�C���x6�߇h�^�Z5Ruc4�b�=��Hv���W7i0,bn�K�{�6D`}q��\)��מ�m�^�\	+!��Z���qg![T�P�p�&�Z�Y���P��a�Q�U�-v�\��0P��mxǲ����\��N�m��@9Z���\�fu��ŔZ.��h̾�\���]�gT�{.����mM��E�����[�s.:d�Z�h�5�� ����uG����l�c��囐�y�C#�C�>���w�6�D1���,E��1{n/;Q��|�n��R���8���J^���
�v6v��ڹ����z#Al��Q��p�,��p7hr�kg
�ܧ37���!Ls���#���eA���*=��V=�ǧg�F�&�x�ʜY�?�x�E�K�O`U��g��	�n�P��tL)��9�J�뭊��_i��ֻ��8��pWV���ٓ��[L��l�v�k���]�ݭ5�QJ�rg�TXe��瓣1ݑ��}�YCf��i��p��'������w�f�*���
WP�ẘ�����̰�>]�_WW���Zp��EX"��0F{,d���c�(p�=��ߎLƸ�4����?ds�jwb�C�5�Ί�>�:�׾Y�O;����}�)�a�N��
���N}��.)�xf��J����Ѝ�S��O���%�Z{�0%H��������� &��Q�N���S��o�;�KzRU�/k�kQ|:+U�3\/��U����\�E�>�6^.6��u�>&ڭ��X�v�ie��BI#�wW����T��4U�f���dc��;�Ab�:u��_(��5�v-�}�,�Z;���B����<�`o��i�:���'�
k�k'mzg�8!7�Ty.+�<�"����D��21䪰]&"��Eޡ=��\������[0��od`�ɗB��	o*
a�IW�����m�a�������	|�H=H#�6�N��9��U��B�UU6�O
P]�C�c�t�$����Ө驼+�a4�d"�Kϝ�$�
�Ds�y3QO Z�w�ndd��v�i@\!�D�m��ӽn��uu��W�<˜A̺����I�0�v���j,^�:��eV�����E��cD3�]��|��T�½6?1��߅i����Kmt�-t�^{]X:_�4��[�,��ʣ���2CQs�Bȣ���+�e�`�kj���<�9r6�` t�%_"CYq[����8C��6^
���F�x�?qق.���==��%"���a�@p���8�UQa���P��5�5X�҅�ޅj�D3m�������e��q;��?��`s�-\�[����P�.
�Ñ���E�ʰ��#D�D�3"E��P`d��ъ60Z�����Y�SZ�鹝��"m�S8���<�D������]���dě�{O�MsX�
:*O���֨%{b��f�G�V��R�d���β	�e"n�2���n3���r��&#+M>]�i33"ޫ�L���
��S9����*�]�6��T5�B\E�������O��Lt��6��̲����)�K<눜�^�cP�U��}�7�Q�֔~R����+���7�;�Έ�\7gjM���Jxocg�8��f�?W3�@��l�cX�Iʏ{S&FT����B9W�v/T:%U=�Ĺ�Yo�=��0�jP��vi��=�}�&:��#�U�[¤�j)lU���ų#�g=����^EdU9$g�T9<5:�����N�O��Au(�c��G���L�M�+،�Dj���	0��"��F̝��3�!��lŦ��C�b��U��f;)���v�ɞe�)��.��IUɷP�R��d}�r�@m`cb � ��oջ�آ~�fjp�5��$�j�=Z��0�{�)��#���=-��z�沥�K7_\4����oE��F�m��}����c`=�����DR�����;A��RH�z��j]l~�돯r�Y�u�.]���J6Ϩd A�CΪ-7^�����폧Cm�>-��
8'�E)�hl�Cb�`;Ph����n���L�u�B�5k2�+Up�e8�H�&��=d�q���)��	j��x`r�MV�Gr�����9��/��y��\�j&(LY���m�x��B�9K!�2��jW�GX**Kq�=�Y5>E����G+��V�ϓy�l"�eڭ���;����Y�Ú�r[�N�f�:ǇQ�sD��PoLg�{}����s�ݖWqJ-�6��`�� �=��f���er�[㆚蹧.������\z���ka���\9�C��;�'M����3 &EQ�tdOsJ.k7Wd��W��ĵ�+O�ٷ~�V��yE����3��?z�ܸp�p�ԕ�*���>��9��<O��+����_�E��������fbLY���a�z���z�w:��
�J-}���p�#<Y\���.�QR��ҝD�w� �u"�W���#d���8|�nF���d;V網�K�&�C������u�oY�חϒ�c�I�ҿ>�m������G�b��7ޮ�ג��x�+T�D�;w���q�`���w\ˉu�+>b�b�cm��K`�O����i��n�L+�9�3�޶�������&Z�lH�\��ԅ��N̙��DKΥ==��_�_)�K:՟[
��9�;�ӝ�q���S=�m����.j��ǔ2�೺1a,|���%�T�)*0�9��0�u�r�%�!~b��l �W�ynӛv����N��Ro#	ŷB�M׺�Db��tF�N�*���'a[�W&z�|��Kf3�HdwR�EKs`�Hr�h�/�D'���W��|�&��]@ż��.���#�9�C ���x�I^v��<,�]I<�p���6�]��(�m��a'�#�!���R�8WX�am;j˽U�|�W\h�/�k�4�C�k���4t����������-���Yj�78^�1�}����� Š�3-���"�]Xޥ2¡�B2���k]*������ʷ!6�ĬA�sp�h��%׭��Î�]�%�i�|�-���3n�<%���9�b��%�o���\�$��y�����{��3!�r��Z��p�����s�m�%͖;>��䢻����9�nh{�H�X�Hإ�QWs�Y���5ڣKfB��U��X��9Dt�&��.R͂�v�0�cY�� 6e���3�;Z�u�����)un�vp��OR�GR�)��UJ�����ÕJ�F�o�hͫb�����m3Fh]�V��T��62P'	�+)�7α��1+hf��蘓n%�R��J8�����+��,A���D��V��Jc���CA�ǻ&\���ZE�j���zR��"dZ�/n#���u��h��F�Z�n�Y�����҅���(�i�ow7�Ϳ�f����H���Y�d����(oHE8
�Ix��=of�K��c��"w�I��\��3;$���P�l�x�7@��Vķ:i��qΙ�t&n�NGOR*�'\�"��;*d�ّjSqk\z�+S��w��a�LWc���k<�,�0��We��(bHW5�r*T���Va����!�A�@�,����1H8^wH��� �ɉ�u�h�����>y��@_v���j�.�#H[���f�+wr�sE#:.�d���vE��B�esK���yg ��6͝�G���_�꥔�kG���W3r+)sP�i��kkR�[�S)c �cK�
Ջ��&^�v��w\���+�GÁ������܏wt�}����w1ł��""�&�a�pTߌL��3N���́PZR�Y�m�����:��t9r��^��F�bֵ��C%NX�c��ͺҒ9FTd��@Kز��JO�4����6��pᒬC�\z�Ɨ�0��׬���޺�7�����}�ld[4�c�ܒ!�.��t����69u��)a�Tu�_5L�d&���������T����<)8��kIʹ��WN�Z�ku�:|H�]�1��|[M,��r��J���eʙcD͘xTC[���e��K%�����v�ˊ�f�2k�Q���M�m�w�h�hh.��f�I�*�yN�>I[e��l�u(��:�b���Ly�mܟ
� � ��h��t���B,P�r*9W8GN��9h%J��W\̓%NE\�*�I�.EL�*F �&QQr#�D��N]9r��ED�+X���\������T�V�Y�Tv���d�EÚӑQ9$�(��5(n$��EDgdZ�q�DR�QTEDQU��F�Rq+�T�W��`TEVIyB&W��$�J%�\�9c�eWJ�uI6vh���h�ʪ��.G*��G*���

(�EEr����KR�8\��T�,�)$&#���AVT\-jaEL�)BJ���V��"�Ds���bED]C�R��J�\�#0�Q�T���WA˜��$W3�F$L�:g�%N�s��DBd�(ix���UI��hD�#Ǐ��e+TE9f��2�֕ ��f��:��Dl��:�5+y�A�{)�G� ิoVnӡ�!�h8�K�
��"ŎX3z���()����P���+�������u��X���&N��E	<C���r�N�����v�q0�n�������C��7J���c}��v���o��|�w�䓿�{��?㴃���ǿ߾s�9��ػ����k�`�b��!H_~���7�'�ۉ��|��N��V�����0����7��޸RW�� �'�9�����;OSv�M���ӼOq?!۾�<��®�4����u��%��~�E�No�Y�՗T���B�=���:v㷾��S�~v�oS}��i�Bt�S����!$v��n��C���@��������'��vr?8�\��x���S]�}������b��˼��G������^!U�U`����`�ߐ��;�=���i�\~��:�t�����#z��n�{ͽN�N$�������M�	۳���-��M�u��0�q��t��ۈ$8�wߞ<.�"�a�TJ���T�'�?|&>��-���o�������ߟ��B�����S}x����:�S�aw�>�y�G��a~����QC��?�����w�bwO�z�O�n�����y�۝F����~��dq�Lr��n�>��30'��@������:W}v�<Nκ8~v���]�����;;q8�|���t��'�o��#�v�~�����S���6�7�r���{��ڸ�����=��O��]��v�ߓ�z��O��~���I���{��8����Ü�
��j����8�|��wô��;q���x����[����o�;_����n7�I��m�ϱ�C��>v~��>l[b�/z���7?tŨ�����p����v�}O��O�c뎕�����>'ht����:w�q�C����aw�}w=w�t�U�w����BM�p:�7�q8����Rq?@�a�0����	���>��j,=��g�>�	�������M���\�a�z���|?{��۴�	�~���;��q���C���;����q7���ޡ}�u`��&����:w�v�]��?|��|q��:"��g,�dt�!۱���8;�f~�f&b?'�8�s���щ޿sލ��n'���7N��=�������©��>��������=��w�i����Nݺx��ߜ7�t�ۉ�I�M�	��x�@�6�Wd�{�6��El�x�p�p�c�  3f�IEa�t����]��?�z���f3�W�
}���5��g7Zc� 䨋YYW�)�^Y54��у��SЯ'(y�KaG~���/72��ѓFY�S9 ��v5��S�������m�B��K��{����{N�����M�9wg�=�n�
o>o�ރ�z�r��缝'�8�&��~y�0t�S�O�8z���r�ۏ�8���s�	2�?;q%�D>����I���_�����G�e2��<����=&����|�q����|�����ζ� ��<M�7g�r�Ͻ�O�@g��4��=�ʝO������=���zwn��
z�&�BC����C���>�[�q8�\����פ�!'��� ����㏞s���]���G�~v�:K���u�������?��@�����G�v�#>Sq����&��r�TO�*c�?���Ǩ������:w��aw��A�:q��8��ES�]>8*1'\�|M�����5�w�m��o���s�G�>g�T3���@�<��b���_OE�f}��\E��Q'�}�|/YC>��>����xv���ۉϛ��4��O\t�y�Ӿ�][q�:@�?G;I�g/Tz�&9���;w���j�.~s
~�����m����^�H��xu����]��q����v�P��xn�x�������I���۟y�@}N����|��۴�P�'{�|�I��~���n<��8�Gn� x���B�>G�Dy�S�)�yy���9;�Ӊ�8���&����&����sN�]�>s�A��aw���~�|w��8>y�:M�	7�I���F�'S���>��O���7OI�@k��*D���*�=*�3r�ϰ6u�_}��v�_P�V�;w�i�����N��~�9�x�����w���m�o��7�����1;����';��a|�?8�;qǤ8���xn�P�O_���@�>½�e���&�^�Y�T�S�7���OC��-����&!ޭ�Ѿ!����߽���+���}���;O]��;����0��	�v��|;L)�B|��m�w�bw��mV�='I�ec�f�V�ϯSb�r�O�Tt=T���M�'�\w�i0�8��:wN� �����q����_S���󏘺����L)��\=M����8����1אI�������=I�����}o��L}���:�TO�����3z���A�5oa�}���/rE��xRI�9�g�(��Y�m����ީNnk
��x�1+JXk��5jި�>���v#9��w��k8V]0��ݓ�a���:�}̭��M�K�;G���Ic�a�)�7�}�U�}�����y�o��{���?���8�wN�G��;qӉ\v}���N'�㰮|�N����|�!���x��o���]�v����_+� �*���U��y���2i���lo�8���u��Rq�]u�8��ɽzM�y�t�W�o��|���0�}O���v��o��8;qӻq��:M�-����9���wǈvr=C�����՞�fd)�1P+��<�l���S�9��8����8�8㏨q>���t��(u�~���\m����w���}v�s��N��?�����U?'��c�����t>��n+��]���I��؎_�Ic�S��uP���y���B~�S��p)��ή��nӟc���z��m��t�����z�&���κ˽v���s�߽�����}=��;w��'�}9�7��aw�'��>!�1�Iv�J��z�MLmǆi�ۥ�O�cOt��$��x��X��N��9տ����'�����8uo�'oy���A۾;H?w�=��Ӵ�|�S��Ǯ%w�=�c�Lzb�!O�s1�f_>�RxQ"�@���"��u�^���W�~E��PR�{��]ۺw�q���+�	7�����oP�\���۴w����v���z�����a_-��:>&���y`q���g�}�|��*��]
^No۟c�ȏ�	����Ͼ��@Mm���v�7����uc�:��N��Տ�N8���n�[����8���]&vQNz���ガw����>5�}�V+������EEM��-��;~�{�g#�'���EL}31�oﱈ��8���:��n+��|>�ô	$���������n!?]��;N����Bzv�s���~�t�V޿���;��D	�8��>��Ȓ=U�����oe�YD�q�o��������~����}~3�q>�~�ѼO���'κ��I��q�<�һ��������L�����z��w�|���v�ۉ�N�#�t�r���aC�;~y�������_��?^'ygsq[��>��"=��?>����t��~N8�į���~N!�7��!��=�|C�=N&��o�;�x��}9� �\}Bq����#}O���v����>�g��E&���~�������IP�ӡ1���a޺�E��v��;��?�nݧ�S�"j�2�Uϻ:��\�w7:Z��j�&Nǚ	��R�oZ��qW����c��^f�7N��_=�dz[��]�bf`fذ+r+T].�&�v�
}*�K&53U>�}�_��\|M��ޜ�ht�W��?���B@�u����t�ݧ�����v�ӿ��s��7�^�|翺�W��ݟ����ޡy���y�o�8�S�*���x�O�R�O�"��q�wv{��s�~�f>�WeO���;zpU��ۧ}x���vV�:L.��
:��L/}s���n����u�~v⻧|?�p;@�$�����u��;I�B~^��nӥp3�~����p������V��F�C����-�/�n��ڭ�>�*awn�}�^���ҡ��c���w��F'x��9��=M�;L.�8~q�!��}?�s+�M?�:O���a�	3(ߺ_���x/^������?|�"N���ζ��v�o��z:v���=�I�BI�������;w�i^�8\.��~�I�N'~C��+�M�'O���bw����p�����*~���T~=n�=�>R��}��?)���;�z�?��:1Ҹ�Bw�y�!�a�7�����|O��n }<��Gn'z��ǧ��q0������nГv�s��IӾ���@�!��I�/��'�bb�JU3PG��{�O��3���}W���:���ߐ��>o~w��7�8�������t�\z�q���x�i�]��uС�!���tc�>���=�c��0���{�c!�T��P��b*F�ח}F���޸\�TQ�����_NFP>$��]�㾻I�w:�~;v�W�K��8�����>o��7n�ڭ�?��׉�0��k��oܻ�i_z��o�A�}O�=�;������s�N�GU�}J�ҭ=���zt��'����>��:C�w�m���O�{9��0��E�~v��=���]��o�n!�9��\?}��������U�������/C���z8�:P^�����9׿.[���^Q�0����ad�%�z���;u��4���{2k ��u��=�0q���+)��˫\I��Fx����Z�`��;j��w|n��:���YX8wE9uҟ\�k�c�H����J�f�-X�ZQ��α�g��C�[�W���4�-!�Z�:t��+�u �����-�4r�(L� k�ˠ�诞������S���j��W۳2����ǷV4+CӰ������a��S�C��x|�nF���d;V��I1# ���']%�W����#��.��}��`�E��3_l\���c#`������.�]��!,���v���K�frXf�r�
��M��u�1M������+�$8��>�s�ɫ���UpOѾR�2��� ����o��R�&㪋U��f/S�&v)��d��S��b�.�|ԅ_j�������l/��hq��@�ai4�����A��6�Sh_[�����ŉ�S��Z]:r���V>����jꇅ�%��X>t�p�:��B�y�d[���=˕�u��oqyr�iߺ\i"��t.vA�|<� �u��\�"�\MP�f/�3WlLU�T�ii���6�\�:�C4���+���0e�>JU>�'z���P���n�+���w���Z��3�MÉs�����G[8�����\r��I;�+��}�e�[n��U2�Z:Xjb��r{S�C��@r�Z�.���*�qY3z���.z
�v6!jad��!ZZ�Z�Д)1[@|��%����������,nu}\Ya�V�kL�i�v"���{�T����y�����7jq�B�ذ:7kfƬ��hl:�^s�3Y�G�K��JWWipu�i�����V�K����ڐd�_I��	�����s'��R6u1�n�>�v�ҳ��(����]t��i��U4e���mz�j�+����j���s�9��7c<��(�f�C�g�|w,�,�k��vnp��$�owo��j`�֒���32�wymN�*���V�ꖴ;ՈӦx�'��Z�/j~�d�R`�A!����<���j������s�'!ј�ȇpf�:���Db�T�{��fz��)�3�
u���yvn�۪��N�Y�ۑ.e��������"��.�+�yK�7�N��>�� �W ��x?��o�]��|���;s���;S��P�9U@��W!Ϋ��j)@[�
�>���4C ��hI�&��Uvۥ�����x`�ýv�/ ��NE
Y��+�e�F����ː��&��ö2L��T
;��1󱪲ҬW�W�8����B�:�=w^��?C��y�	��ʀ���'�P�]W��|$�aO.����TE���t��3R���qBc��d_�;HK0�k�l�qD�qD(�؄��0ڝ�S������floϘ��݈X�PEN��f��F��r�V��ygǪ�]*��{�nM��1��v7.�X]1���X�i�ĶY���ǨJ�?njKBz��`IH>�ˋtI��i����1\棢",K<&6�ق��={I�i�d{�yQ	�f�Tw*�ũs������>W�}�s�'� 1VY�/Vn��]۱N�#�n�x-P��)< ��]�y����$�PlDk���5{:i�\��%��/��P.�t��b�X>�OK�Z��K��^�Q���Rx��I	y~�J�&�Mw�.u�ҀԽUz� ����:���|�*�oX�qD��Z����=S5G����6vn�6ՋԠ�U{|ǋ���XX��k:��ҫ �;ʂ̐�D�s]f:�S����{.�i]�z�p��݇��T:��N�hdCYq[u��΂5#!�h�vzW+��8��Vo�J�cE�`!��#6�UW0�ss�rs~N�6��Eu�����%�8�z�}�w)!�|��t��[�:���GW�g
�1q�TXr�c�";�Om�&Ƭ;1�L�k�R�ʑ�7#���3��x[i�a��Z�=����O��_W��k�v�l�W�R�o�(��s�,��́Wj��K_#����d��̈́�G뗊�W�N�p�[�Xz�c�=N��z�J�^a�jV���y3z+�CEn5*-�ڴEK�	t=,���/��Zg���#q9G�5�.�ZfM��j	}J^�]��O1�$�:�d'{���Q��^o+E�+`ej��`Ye�%�Sѭ_$9b��:[��*��e�0 �z5���O>|,;��-ZZI���ɬ�m4�JǷ8��e£\2+C��}a�z�gg���ё����Lu�4xi�NX�%y����!R��Ra�-6�힄B\wQhq�\�	"����-CH�.\Qn��Y�vyq�`M�tlMWt��[ɑ��ocN'��
��ծ�w=�g:��	nݑ�RDՏrD�=Z��+-}+I��L\�u�������
8�L��1��.y
�ConS+s�}��91W	�_W�W4���a*���t��#l�4�c���Z��ǬD����f�qJNUu��w� �3��}Ey�F��YP^*]r&�b��VS��L�ZR�[&C�U+�U>|]�ͫ��L�)ә���M�/�Pi�o�.6�J�+C�ԍ��li�X�:��Sa��UGM�v���)��"�eڭ���[˹�j�)�)QҔ��h]�Mg,=���%��F9�r� �!0��,�C�	ݖWq\���$	�Ol�-��W��m�p>T��eԯqW�b�@�q.}�')[�\u�ʺ����{Ҏ#p��C�mp#Z�=]V=��u�l������J;�%�C%=�T�f��u�c��J�Q���qN+ڴY����V��w/�ZZ��vM���<��
���w��O���a��!�]�+���]&����P�����w���^�5���M���7(�A��ǊO}Q�.Cg��x��cZo��ʮ�^��x������}s�<P_1在f�y9���b��]� ]^;�@Ê���@=ύ��7垽��ͻ��{I�&6з1jmw\R�?l�l�J����T��pxik�m��\I���g����*?:*�y�O���7$��x5W#�EH�z�d#.��>r�>א،v���ê٫
�bXz�yg=�y���$���.%���C�Squ@b�[5�[�~.��F��O\c9
s�-��V!�����fh������`�+�$>[U�;n��gg �x��.�� ��Λ������	����|0�D	�!|�v�ڔ�-�tT���s�/=�2i�$���`���R�}� �z��-l�KabB�Ӳ���;���\�������\�C�'�n]�A=��u���4ZR9œkEL)��@���T�݉�Q��Ƕ�]H�(
��0����8t����;eС�b���x��'����e�R�L�1Ȫ
�T>��#-CV�I��ë�Q���%�J�D��|��|+p��;/�I}J9��gn��6�S��-$�#5��ItE>곫x�Yj���j'mU ���^�巌�x�o/�Vz�3���g�\:	�2�nfzs�6%ȫ�.'��[{��j+����Zz��������c��F$�>�m]M�������/^�M� ��3ѕ��L��{��H�P�p9����W�e�g�l��/��,܄��"�p��k�� Л�8n�]�[�W�C�tV���*��Y��7��^@ڦf�(���GY��N~�B�j�q�t|qnn){��b�d_c�,�sFL�z�-ai]�z�!Qf�{�_XE�v12,R�#�;{���5���F�K�E!�V�7e�\�Nb�^���8�Wm@v�8��E����X6���w&����q535Y{R�C`(u����t����gVЊ��تZ!��Jbm�c�.j��s�㹕�;e���D4'�L��
�ǟy�o��%쮷G��WڈXI�e�͵�r	n�. S�uN�	�u1z�����#>e��0�*<�����μ����=.���49�E١#��/�|+��n[�Ϧc\n��S	������{%�US��ū�A�W�
�~QoF�JJ���94:k���[,9!`!�@��-�B&�l�'��mP��:�nQژ���!8j���֫S���ֺ ��@;ң�21L��B�4�`�_^+ϵ��d�*���I𢴅���i@xlf�
���
�������y�{��t�1�s���kc+�8G(��N��9�yVg ����[k*֘�����lk���\-r����|�]R�x���h�,�4���Q���of�!Yќ��yʃ�6��His����g6hڳj�m#Q 扲9�S����ΜY���uI��w�`���%��P>%�bm������� =�ϖ�)�K;jŏc�e�6��f�wq����|n5z�K���K��;E�]m�C']�Oh;:k5��m=�~���jQѠu`�{+{	��EjU��-r��i�s��\�11k$+y������p�S��G6��+e�@� �6Q!S�mgV`���(T�S�4e�q�縶�>9�3��Z �v�^2��NH�	�Y��EA�y�k�"��΢��eM���eXJ�0�ދS~,�����{��Bյ����B�����u+\�����1�G[������a:{��PUˮ)�x���p[���猩N8{l	pm���Ji=`f�&K���V�d���˛*��u^��Z��)����y�F��m,yr=���������M%R��L��`Y׊Z�ܜgZlSR�V�wS������;M�۳��6𛢦2���V_�ܦ�F�6��k�ƫ͖6��f\�����"��$��t���#H�/a�oo3�Jƻ1vGC�X{6���!ݲC�%Kƿ��,�ҝ����]�u:rTV+m�w:8��i��1����;�L<˧GB\')ŝi��G���� �!X�ǭ�Y��z�9_bEI6Y��r�Q&Gw������j@��(�[��3Gb��I{��qU�a�w��X�66����n�e�͙�,g+��,%E�W5�t�x�+)��
����Λ��-�}y���y8*��4��P���]�IL���	TN;��!��m^;&���&7�ݴm��ӈ�[V�hK�����\I����6�{y�Q�� N#�dfg2�r���P"�h�n�3fOg��*��3軲��j!��"U��f��7׬�n���x+M>�ƘS�)��{��c�N���5\ȭWn�{O3��xT�#�M�k�V%�\;�]|h&\�p
��֣ j�����`�����c�,�%�ǝ!dr�4+w4mج�NF.�Q𗕭tZ��c�;�[�Fչ0�	]��É�ǽ:�ud*���b�F�N[$W�Zx�Ӥ�l�fT7VA��%5�Q��"��J�t]4�,�ËN`�}Y K"X.�gR/HP��jM��փ7��5i�	|+�!gKH��i_gb�����¹�3K۶kBTP?r�����+YeRI9p^�r��W��W<�ԣ�
�t�(E�fL���"9�sL-9�
rҭZe�JYZ�$�eG�����.YөH!�ST�Ε�gC**�YNq�<HEU�S.fb�]�!aE
�,N*�CI��H���8�[Y9�/(h�Na�*񤰐�<�'�r�2�FU�ÔdFyȨ�S�%q�ĆHar�P�i$�r�T�QG0�O8\T�"q9Ès*��(�Tb��FT�\G��9]:A�n\:x���!��9ƔU�BK���b�x�xJJ+����"D��s�J�Y��E�r�q!x��b!�I�5,�R�3$�B-4����"��RÖ��WYD��!2L&�Ef��(�g ��t%Y��e���	$Ȉ�f$�)j�u8DU������5L�N��.�,Q�(����f���Pk����*l�Ҕ1Pu ���t��ޔNWn�]/�rJ�q���ﰞ�f�fdԝ_RQ����^>}�g�}�UMmx��y!*���z�QW���b��ę�W �����*@g���y;˲��'KU'�m�謹R��#��C�#E�W
<s��z"� �s�o�D�찀��p�f��vQo\V���K�;�Ed;yp-����&�<�~o�u�P²��ܬm9��7.�Q�[6��ZAR�]Ј�SoT�u���tY����ʯs�&j����
[hO}��Uī��Hیz���|���{�aZT�O�
N=v�
Xu���fg���±���y�C�v��H`���R����^J����B�ab^:3t"�$�PZȌ���HWm9���u��ԧ$�v�y3J�K���C����u��֌���^}��;~������Rz��2䗏1��6�j^������sH��T1WK��O�)��Ӕ���<�w'<ڥ�=}�*�w�0T���3�	ݹ�Υ����$r`�"m4�J���fHs)��W^s�I1��'ʗ]g�'�H�����bw�A�������&�9#ێ:�����c<�V��/�������T�DR+1�S��Wm�UGG4r�FH�ë"oxV����݁�!�K��e��1�|��KSIn���A����v��W��WF��J��0�Ι�z�7��J�(���U�s�9M;���>����ٽ��������E^�p�����XY�3�
����CzY�ύg	ڻ�.0�4���u&+o��A�U^g�{w�t����U<�¡�_�Qa�ߞ[`ʝXg"�I����e�Hc�l�!6��R��w����𧯘��7��f�?����u"��y�Kr�U���^��~�U�N�c\n�Z���*���^�q�:���<��֨��$���{.����;�8�s��eiO>|2*�ŀA�lݩ�fz#b*�rJ�w�?�v8V���y�P��Wؽ>M�Z�G���'m_j#=��΁d��@D�w^��2��pg�\�Q���y��x���Y�}T�(C���S1��7�wZ$�z;���I�ɤ�"a����X�����I�1�B�\j6d�'���Ԑ��f4MK*+�[κ���t�[y�9��*m�� ]|�����f�M��:�9N#�(�)�z��aQ�D�e%����Tҥ�$+}8�q4����F6�:GG��zY]Uxtգm�4�]W���hb��2�����OkD����wXn�����5Z�b�:<b�W5������IBե�ut�(�zz����ۛ\�s�J��}�( J\v��Rp:1̺� ���)'nv�ɇL۩���j?���qp�hA�DD}��ڊ,���Rg�����5l�.��{�����1pB�;M�c��<�7�gCؼ��r=�yo^�)T�d�^[�ڼ��N�2�ӧ'Xw4GJ��Kd�@uh�N�w�@��k����kAh��O����!�����bo 9��}�Hu�Z\�!^�R�Z1x�������@S<�m�����V:n���4��س�UP�9����̊7��ZQõq��^$@:p�*���$.P���.�f� �rU�r\��5��]��0\d��)��؉]��M��o;eG���c�o(���%�+OCf��ͫ��u��h� �2o�y�9!����������(w��a�2/.cz�K�^�Ia�
�=%�Pc ��'��swm���o��x_)�)��~<�)[�T�he�k�(m`~��d���F�|'>��X(�� KcR��Hv�o���p؇F�룪����^LS��9���OÜm�_�Jf�y\,������Ķ.k���~��Vk���LF��ߥ�+�V�t�[��Y|�w$v��*��D��yNW�K�ik걆�}�W���U��ZX&�AZ�{<��rX�a�r��[LR������j��G5�m̔:i���~��w�x�0KoN�v��ˑ�V�:0K��j�mǼ3�8ӌE���eq����>�˵��h>5�F�܎
&d��LԚ,VG
H}�.��7�n��3��{[�//�*s�tR)O2�m�C_�W
�<_҈:>d$k���ԧ�%;���v��<�������w�k�_�� f��8dM1�șJ�ѱ��2��o��Cl�9܌�N.�u�s����m��t7h�s���s�&]:C#��6�,�Q=���j��A��r� �$R��ܢA��K>s|и��+�B�vd=�nfzs�2eU*�i��:잃�v�<	�+t��u�魛�%���M"{��JИ&�d��������,��ת���P���^<�Ţ���=�4�u���<��K�q�r����k�@�R;f����h��v�# ��^ش�џG��jЅ���TwiΤ/<�J��NN��e�w-N��seVm��0㊵0��|�nhɑ�s�M,½�� �@�3�xh9O�a�	܏x\۞LӚ �ou�)�b���cUs�;��<��ʧ����hzo��Sz�1�H-�	t[��,��&b|[��-K䬹e�\��),���2J�}y�K3m\�L��q+O)���nm�����`�eX˓�Ɏ��:]���mE�_���/�E6�J���5b�$�#r�4��N�"`X폐;(ҫ�j��j�sԭ�����}�|�v�zL�=ke+�@��ؚ�35��^��ʆ��u���-Y�6:{:��T��kL��RB����N��i�f��UH�����C�7\;�(=M��U7w�g)�=0�E�U�$�'G0��]n]���8��/S��GnD���6tdU���-5[u��al����Q�XB��"����\5(ߎ�Ƹ�4��<}o^�/z���ݫ�2ק��,���� ̑���vc\���, v)�����U	��qN��v�&͖q,�r�r�h3�ὶ�o:��ɑ��V�:�5>>���a78����uUFC�ՙ˶��#'P�d_�u�qE��&���j���ԯ�&��Y��qz�df�ݬ�7�6�)�i��$/��6�H}�Bc��D_�S���u�����F5{3q
�`\���Q��l�	�E���af� J-�"}�V�P�V-J:�8�bua�DX�ivu34��ʞ-�羭��,U��x��U�]�?�*�A��4�ԋ��WO2=�F�=����͵k���U-�����\��������x�,^�\-c/t�Έ%�i]�mg,����7ćH�;f]�t��yB�rظ�x���u)���J����&�(�%GFz�7u8��{y�O�,�d��n�=0ȹ��ܚ���r��Vj���� ��{��7�k1�F��d��`*��(�8��1}�Y�����-��7�W�n��}iQ
.�zF�)n}�:]�u��<����u��g[�����p����Q�v�j�]Ԃ�}.'8��T5f�\�/�q�NDN�S����U���<���kƐ[�hS�����If�;�<��ս��Nmo�>����:cd�l(�ÎvD�uY	�����?nt��@�����v}Ui���.*R7�8W�DhX�ƳQ</�AeV�}v�]�s�v|�ό��e�v_L{[n��<=���PѹNv���N�OW-V��+>�P�.
�Ñ��Q�ɉ����Z�d��0p�/�w5p��p�\+ѕ��P+O
D�VV�r���y+E��Ŕo�e�#}��闝
��|�6�<�,�
�"��C0D�p��n�����q�*�r`X]��u�+QJG�u�d�r�쯹�C��w2�!�{�(XtJZ��SI9Q�It����g^o0��糀̸9g��s"�Ϭ>XJލ.����s+�k6'��w�Ûae�Z�N���w�7UҚ�9({��R�g�sZ��e�O�,ámn�`BhZ;����3�VV�f�����sM��ݜ��l�m�n ��RV%z���Q2&]n�-�1�m�S^+�H�զ��nQl�8�И�V��� x-y\�5��"L�z"��Q�0�G�ד�m��+*��3���L�^7�tu�l-�v�jާ�䣷�o!^�HJ�DC���B]���M&�j6d����� �_ڧ��_I�/eŸi]x��8����ߦ`����s�&��f�r+�<�9k�����_j}����n��|Y�ʭ윗���UW����G�\�.']�z�)��#�ȿ��CJ��6���,�yk��r	u.��ʕ9,�}m+`=�t�K��$'P&*@tH��^T\*��
�C��牺ޒ�)*�dod9��^㝆�匝be��t�x=[y0�}$0�pB�6�b�9-3�wف�Y/<$l��C����0���F����j�{�p��x7Ҵ��x����	}6j������6|/>��V��9?�ܔ=u;���8��՛���ݸ�b�Dg{&ڐТ�ai
����&n�@!��z���s[[�1@��q�<�Z�Z+�cY�w��2<��֖��@f2���x?��9E��������к�9ΉU�,�y(��ǘ\��g�p>�Vv�<�Cn�.:�jD�]�D���҅'���b�F�o���RF�on֌�t�.I=�*�r;����J���v�h�r�K�'O�y+- �p��Z�i��2����$B�\�zy��\�¨�P{.�'�ј�+m�ʌ�w��=�1��3��>����~Hq^�˷$@=�>7v��YΧ�4�.�������5��z�Pg��؉/2~������s�s�+/���]N�e"N�Ж�n�é��6{�d����?5�ύEHB�Գ!i����Z��;V����=8�˧�l��IuY�l�&@�L�ҍ�Ö����6*k����u,27��z�[FT*A������#,ad����`L��S7�I��W�Ck�"/�wG�ma�������2��uV��u<Dm9�o�P���2�o�̅�5�Hz��-�tP}���%�7G�,ͳ~�o���_��k����_u���^d��Q-ɌHG�zvV��e�\�Z��w��P�*���6��p'g�k�n�9�@sU�7ELK�*���KJ��̐��t���/�]��yM�z�|����d%p�_ɻ2Ļs3ӟ!�4��
��̨��%�p���oT%�(����̋3jKk%P��=U��+���A��%*��w�K�5�(%�؁n�[�e+��ͷ���;yL<�ŌU�b��� U�:\��ʄ�o�=�׀�p�]��W��ܮƀ�I���w���|5���RR�A2�V"7���  ��ΗkU�[�f��2�,�(r'U��\:D��ksS���������9�5+|�=����VIU�ZbxV�M?n������J5:ODoWR>i�f�}}׭�f(�B���1�
�'j-a�'?�)\���
��`S��/ǠE �y�X�3|S�{W\U�������eژ[�7�sFL�똵^��̠��]��&GbE�S�y9 p�]ln4ڻ ��	����k�rP�9��N��U�p������,@�P��R)]�T���eg�:�ÜM��C����/jueC`1��b~���ⲁ�Z����Ib�+�ѥ]��p8�y�2TCBy�ʙa�ʢ�<�>rqј�N&0�t�$�8ʃ�l���� VP�@+��뺌�⺘�N�Y�nF2��M�U�̿^�U��z$%Z,?R0��
�3�4Q��� 뢸@�WZܷ�1�7*.j���sn�sEZ��$#�x�~q���s(iMd3�
�"*`���W �<���w�MD5T{�����;\
p��,�sRs��^�B69���qҭHr�:5	���P�*79s��kGr8)n=��}���!d7dN�YOr9b�%0�\C8燲�SS�>سy�L��R��MV��l�6��2�r���e=s��։��^�.Ț�L]aGMج�ۗ56q��pV�c��h�9kN�ޅ���[ y�;��ܔ������	�������3�;<��gS7a��3��#�!;2A��1��	�G�m�P����g{�����)�S�S��M�!�}Bc���\�!���66 =���^�óZ-����}��쭘6�c ]v*烺׹V���OH0)o��>�<)�zǕ>�DV����˵�6��;�� U��CNQJ���x.U���-�F�Ȅ~�~����G�r4���1��:�(U� gPsD��P�M-������v�i_-��6MXy��[��;I^TdT��Ϻ[ww%2�:sSpM��u������],-���������9I,rz�,�0��s�WNx��1��ܱga�d��T�<���Ѐ޵�8��|b$�O�}j��^9��7�u1���1�Gvs�"_:�N�hd5���s��i�#N�Vc��\t���T2�	K�H]]D�V+
cy&�*�����3��>'�B�;ڽ��k��9쩲�����R�~��YW��y�_1�CO�uiU�G������V5� �>BkO��Uֹ�1� ��}�q��%VqЫ$ʒ �6 � �^k����k��/��pj5�+��V�ηJ�����e�7堥�b>ձ���Vn���H30:W|�G��.� Pe:�!��}D����)*�r!/���_N���f�������z�.�-�՝�����8�m��Y���iM����kc}�d5�ޥ�X5�Q�ft.+���㜪�O��u2)���ut��yY����l�E��R7Ӎĸ�jzZ�j�iE����۾ ^���R�ږ�ˠ�#(i��$\mu�Ω�k(���Cq�:�����fbO3	&�a!����ma�z�U���&k&�tveX�u��M�oKUe*��Y2[�6��w�$	��4pj"Ep[zV�r�܃�k\��&�͚�YE\'n��2��K��ћϤ-Z���׵�OP��'C��Ar sy��6��2VU���s��+6���ȳ�Y��k_KYx2Vun�J�����Y���&�BH����V�5��<Оv�����w%`;!�M>����P_9C3�:����¡2��KIk����Ύ�@hp�^P�%q��Ebk^�\�<�����rݦI�i��G����������^�3r]�+qw��g7b�::F���b\;n����KE�)�+n����X@IJ	h�Y���7��=9�9�*PQ۩��	���5�1�\70���ܧ;\鈾8g#&�[C�����һ���	��:� I:�L���u&_t�C4�a����6Q�sH��q���l��U�1yJ�0��=t��)�%�YٶQP>�-�L(o(/�P�Dj�d2 lѹ�)vZ�g�������S�$9�R֔�u��Y���୺��_$z�g:aW�l%ӏZ=5�����=g���(e��A����h��w��cif-g�j$7��^%gB�C$u�8��Ū�h?5�H�**Q�� y公$w9�S�����ɉ�;������g�V%9m��v���N�L!am^D=�Vd}��;!��쬂���<��	�>̬V�Eu+=�)vb��F�Q�����/$$Pz��h]�o"唥]�o]�j�2���,��rf��';�ɫ�u�3-�5��L����A�p*����_#]�䲫�)+-լ�2Z-!�G���I�3�{�B|����s{�vV���7Ǥ*��v+/W�ovkM�n���QW5�7Z;je4e�ε���AAC
����7AK�W�c�/;U�dVrp�#D��[��e��ռ�v&��/d|*!v�=Ү��ω��[���&#�b6��:U�p���/I��ʱ�JXo ��.�W\f����XV,i�f�.9OFq{c�O8s�kh�+8굖wp:0��ǣ�z\�dZ�ب�HZ�V�������?]��$�.\*�B��в�L�b�*D�f��E)RV)�hHY"�BD�J`�J�V�X�`fD��)4�$��g0�P�J�NGΔUQF(Qd!Z�eQ!�!U���bJQ
N!De`��Bj�H�����%@�Ӥ�$%iXjEb���P����e$T]34��A*���fFQ�rYW)�LRT��T1!V(��"LH�(�2(���
��R���\�#�LJ���$ْVL�靦�UE��#*�RVUbf�9��I�B*���I3H�C����Vap�
QB�fW9�E�����4�9&���9I�gH������E�at�RTd�V�*��B�NfUE��XU�iҒ�:a��	TN�����BU��Er+�"@�M&��+�1L|f�{-��,��ΐ%I�,n��9�������[�0.�m����渖�|��ٳ2����	'�?���ﾪ�����sR܋C�:���s�i�p�\+ѕ��+B����Z�AQ՘t�:�P�=-#ݑH�==_LڅJa�M��,�;�°��q�7f��U���U�<�fW:�����&.:j�UY#�3۷Q|ǼU߳�7}����بD����}���o~ܫ���`+�m�돖�p��Q̊c>��})S��R�vk���5�خ�Qk);�}3/mkd���@�N��U�Z+���v6��H���k�����Y%']�;�q j�Df�z$�(�c^d*]���һǄ)� �6d�Rx؊[�U��1Fˊ�=���&s�/�>:�>���7��U���s�$If�M��:�B��{��˃�x<�'�)�M�#����_U�K��)��<-Ø'SK0��1����t;�{mlTNs����9ʹ�פ��U�Y�eK�f��ĺs%�_�"� :�T��)w���Kei�U����!Nэ�1p��s���:����}�v;z��]n����F���u���$�<e�>�=�̓ݔ:e&����v�i�T^��ـk��;޲���*`L(�f�Y�R��u��r��T-ycBԅLN��!P�y������d�eAzLᣓ���vEgq��v�9�u��Q���}�4�o.n�$��2.�J���c���A��J��v�\�,uG��ʵ��/�򜜓����{�zT33׮����H}8a�i��<�N,�T=KF�-G:6Yt�QƖ�b�x���T#k&�O�U)�&��3�q}Y������l��=�4�}2|q����Ƙ�u��1��N�Iߣ�k=ii�@]�\;�^��x��&���3�n�}9�K���̙s��8ݖ*Ht��ht�r���b��0ϯ.c��=��Nl.��pV���%���dŸ�St��j9���C`M��{n`�;�>�U�~}����"Sqڅ��>�>��ޅZ�����z�)�ndk��ط�9[��!�չ�(8asU4a<*{�'��5+UzK� /f;��ʋ�uL9�]P����_%��.��EH�$]��o"�����o�CR�6�S��0d�;�+6�O&s��{���jY����g.��ĵ(�*^�w�w��4����?�ʸW0���QGT}���@YY����>��/�{1��5���}:a�i��k�t�iV��R��<��^��˂U����^����jU�q��
<���B��T{Q���T�,�:+R���m�Y;��ȹ�+ v�f=×#I.=��W�
�n�\�J� ���9X������ﾥI��/V)�r�R�}>�mdC��:~N�[�M1�!�`���-&��[�.�?p�f>��a��\�3�
O9��c�@����2�!˜��[2�\V�StN�4E_9m�G�\�К��62S@��Y�h\rU��ݙb]���Ss-Y�Ь�u������W�W��Cf/��`a	㌘&�����QRV�`X6+إ�؎b)^��v�SRT��r، Q�`���u�~�s~GZ[��|����d�yS�Nfն�16�٪ݲ!�~��۪��tu�g4�_U��*���̯ ���/d̘�_&�9����"��끶2L�'l�"�����y7%�U,-+�Q��I٥�����s�O�Z��j�s2{]Ü�)�b�;>�2��]�e�&��,qh'
܋׽���ivEXo�[Q�¨�s2q�ʓb���}E��r�op��q0��lF=�ו���� �b�ad��2���#�̬��U�������Zz �_�s[9衝���oܦ�M\��rF�G���8d� �{6�OI��n.����kui�}�
Ѷ5��o�+�5/S��i؄���]77mR�qu�[YH��OE׎��]ôjy�Gw5�7+3�RA���;�HNY��SI{�z�kޟ��ﾯ��3������w~�u�U�p]�I� ���Y�v�ڪ��N�].����T�q]�K
���R̻���r���~�+t���9O�Y\¸:�n[�ip�Wu�Ӵ��_\`|�5|�"�)�N9�#�;S��p��g`V1��M��0A���P[};�h��޾���D��k�d�yg����52�:<4.8�X�E}�n�������n64�����S.D��/�7����v��[l����>�Q3��M2{���!���ᄙ��i
�p�S=? �􎐈z���h���v���a����}�:(gv�&x��}>շ��\ɁN�'����R@�|����Y��򡈁AG��V�
���K�׸U�ںb��W��y����$�hiTR���.U���l����^R�^���y#Ǻp�����v(n�9�&<2:�254�b�Y]H'�(��:7�
3�{����7�I�
u����<%���A�6>Y��/�Ct��޻��yq?t>�g��
��G4�|��\�K�F��2C|�P��_�`n��Z�/e��뫭;vl�K(E���BÙ��]��ά�r�1�Wy(���ue)S��&�:(8Z=[ʘ}jK&����r��:+�����\+3�"Ȋ���Tg��>��<=��ь�V��)_h�yFa��8�'o)�UN`��ܱe�\�`Ny�+�VD(3]j��U���tD���i�;���'��8�h�j������jw�Cˊ�|-+��[h�W���5Q�.������I�ޜ-O�!<";8�v!]������c/��+�}�+}b�ԛ?67�U׈�z���K�:	}��:2��=�(����#Ү祡��w(��<��^�+����5�sz��TU�2;qC5>*12 �
�d|h������w�=�:�ά��o%���f�:S��wF_/�f����	�ϑ�Qc*a�U�r}���l�Ĥ�V�S��;�k2al|Cw�+}J�3<�����n�Z%дa���V� k�rQ�9��� �W��
�ie�7qL+�ҕ<]K��ep�QG���U_�v9�/�Y��|�@�v}�Iމ�&KC��A�����V%�T䑁T9<!��q�F�[��'�V����ܟ�T�!�K̄���@����j�]���؉�U��^��U��u,�wЉ��YLoϒJ#��;�ۈf� ���(oVR1xJ}���G���u�n�W@�Ez�pR0���u50��B���;l�l�,#O9�=��J��ډ�{ƻ,��*��1U�5{g��D]=�U�t��n���Yrb������J[LO꯾����$g���k�q$W�f��,�}��L�!�&�ǜ�����|�����o�	�J��[���Qv��g��}�!��T��6 �O_��k�4�.'XJ����iK̲��i�B��$�]3ˬ\��㍊�T��y�T��f����l��̗�d���1 ^w�D�S���1p��?��"���'���Z��Ժ������Ӡ��.m:s<����NZ�Xb5;�oxL�S�_�j���vg�|[�D��0TAO0�E�˵N܃dF(���K.�K�(���m���ؖ]Q�u.Ȗ�U��X#�W��`0��O���.��tW
���E��v��@���"��&�����F�
�n����uÛ�EPc��Kw=���f&�h�=w�JuK��ͯ]nt
{6�XP����v���yW^bY3Q8Oe�F��U��!��s&r"v\�axX�ߖ'�N;���w䁨q^���QL�<u�b�6z���ȧ����@�0z������M����&����s#�ve�lV_����c�D9a�q�u�Jq��3��@SU6Cn���`�n5j1�t����}v	�dp�k"�Wk�����J��d�B�X������d�4�љ���������X��;��V�Nv˧�7)K\>��qm�ȎotQ��m�N�OH����*��_UW���{�^��{mk�?Q�&�� (s�0:���\jY���o�����א؃�+�0��-L=�>�.�6��O|�J��RX�&����R��@<���/�!�n������vL'��y�)f+��p��r}]��%-:*�ՠ�������d.��3�qm��sm�������c�)�o]�S��ѵ��?*�\�4x� I�25�H���,�yѭ�խ�u��zGLbU���:�Ր�[��J�}�*1���-l��� ���̧;B�c��ݴMy_�J�u@��`5#��8u�Z�K��C&ubȬe��KmI���kf�n"8�^)W�fOJ���[�q~�j㒨tɻ2Ļs3�#!C��}+w2�:nJ�g;�=X�"��ZO��D��1|�.��ȁrX�����>�m\T�Zm��+��v��M�-�u��݀Xq�nd��e�CVI_E\btqp�����sOںo�m_�T��t~�Τ�E�$�F���|�a��΁�}w5β���h�"��g*3W��^@�� �A똒����Ǝ�1zf�{���k<+�MҖq!ݚ,1ڌ�S����d��B��@�k7�gR����s��f�A���:9i�Q��e2��Td*x�Ώt�hF�� �3�x�"ay5KI^kr���a8�U�hV<���q�M�b8���MnAr��F��{����:�
���6wq��u9X:�K���A�jao��î6�XOcXtq9�E}�q^���)gy�f�lx�6-5�M���A��| u��^�1�Ru�B���lv���<����8��gz�JH#��C)������_P�L�5fh�/jv!eC`c�����xpt���J�[�mO,��h���i�;��g�hŴ�>'A�������� 0�����1SKzQ��ޭ�\��ҁ�_z��G�m;�+�}�
�ߨs����=��K�ߡ{D_��XQ�淑���r@��n�	ۿ��!�Er�"�+�T�pzܷ�`��S��θ��Z�ÅW�56����܍p��M>�m\Mɢ�MѴ��<�%����r�el�<r!��t�����֎��fv�%q7+s�j�k	��]���ޛ���:Ljd\:m����}=�z}�^�H��E=�ĥ���{4��v�p�J����݄8�#z
idK�moZL���a辴M�"� ����Ѽ�`�{SS�i�~�� �mE���C2�}yv�Q`%,z�8�햃��R�͟X��!��e�'3]����}a��ˑ��&&z�,R�e�aW%&ȹP���U�W�R�Pgw����Yjc�(9�Sr&gE�7�t��N#����kR���Ο}�l_�ب�%�J���5f���!;��
3�����ę�+����¸��ʭ�q��^D�r��" +⧢K�{s��G�z������z���i�2o�����r-��!d�ؚ*z�quļ��4c�Q}z^��r�h�Y���#yr5k�wW\:�M���_j�5�༚d\�y)��nd"�
{��Y�/����T�|�ã��u��q:o=�-yoE�d'��.a���>���;�V3��v��w�e��S-&�eM��-fkV⑊�߭{��>��+�j��Y{�MI�Qe�yM᙮���Ie����k�����9:�ǃn��զj��Q�����j��Ʊ{�Iݕ��4ʹ[���}��v,5�v��,�Y�aL&�!N�:�;���KS��dŊ�ƪ.477�܄�8�ȁ}G��@ovvxjn�V���r�m1�)���j��kQ��vIͼ��ˮֽ�,�fR
�ӕ������g��Ǧ��څ�U���Ѷ�]�KrKj9xt�4�F}r}
��]��9QZ�Nݩv�X�,�+�f�|����&<ͦ��H�#�� ��VK����UUW����O9;�o����3v�ED�����S+X�.y��'fDt��<N�j�,�ޛj��QI..:�K�3��$���"5���3�zc�����a8\Q���"�&����k��JNzRF_���7&F;s���D�e,ż��o\cs��
BU����K�"8&�P�f�;��Vz���9F���i9����l�nv��
e���z@,��K�E��5;���s���낋Y-�y�\5�Bd�Z���"G�衙��Oe�u�O��,���-�4�n�N^Kq�^�bm;��EVZb�d6�2ѩ�!���Wûw#m.��]p�׍����&�X��l9��x��K;��	��e�-������%��D����c���1n�r�j�܊��:��X}�2׎et ����t���-�w������ZU{�]���(wv�d`�q�
�oZ����id���Wc$���*�J��.�(�V��t���LF����{ײ�P�spp�m��mw�R�:07�s~(��r茤�jeuX�RH't��{.q ���t�
�� ڝ۬4>;'fY
���K�j$N�XF�)��A3mӕ��R�TfvtM�/�\���g�N�j�ϬTF;���͎*C��T#��jM�L��;t�r���蘍�b�Tsd������v��iA�f�&3k �|�Wd��#��L���G�wP�Q��i[��W�r�9D&n��l;@woW_ ����JK��I�Q8(�3�<��
��Kj��7&����"9�n�x�ڃk����W�M-�)��yC�Ufu�F#�@��q��VӋ1�s�����i��l�& � �=�����
c�����q4��N�2��|/:�E�TD��:�t.��7��V+fEL�����^�L��"�Rą>Q��;sK�r�/V$E�3�B`�oFU�w�ɹ�o6��*nl�a�Q ��ص�_Y�U�jjq����fE�����+���.�5�L �Fh�;M �;�������8�*�MD�Wu��ӦN�Z�f�g�54͢�vm��]����9�c�ʹJJ(���n�f��*�d=����Y��[V���ޙ��.�����b7Km�sZ��c��q��z���pk���+8+���]�W_����t��J�䳄3�g�ʨ������pE�o�I���G=;�K����UݜX��84Fc@݁���D����NL!+�]ܳz��4���<n��%-ɽio'��9�r��NنKvY��u.�R��b�*�S	úz+�4�@��6�S��+����2�s�Kl�� Z�;Ao\R�ah���)u�S���]�,�wK���,i�;�Dgk��X�%jO(�${:�v�1���F^L;*I�
7��ǒ����uݻ�dۧJ�,.L+�G�X�QF��4v�x�u��Or��k@��^�S�v+��uwl	YO��ob���;�G%Z�@��k�!d8uk�v�m�]*Y�zi�l5�8��W�v�@`@��/�$��E�z�ͷ���7���}etH�w��r ��VY�X�a>�)u�a�@�����Ed��f+&��:�z�@�֩oq��W{Pgw�F�RξH�ls.�nA���0��9��MĨK9b�&q�b�ʱ4�%J���6䠵��fmK*d�f�
���ס� x�H�9k�X &���7׸�Z-�t+歛Xw �2�1BV>"�n������C*S��#,���ۣ��)g�bՂ� ��+T��H�;J|��W�Nm*�y"U��>�W�.����!�\ۀ]�")f�b��Wb� ��E�z�r��6n���,;`�R��9��4��B�7)`�G��Ӯ�s��t��ϝ�>~!ʋP�g,�����E֔��*�5�]#��dEBh�4Ij�lH�
��",��jaVV��J­�H�l�T��3�!g5d���)�I�E,�]"MR�TS9��#-dEU��kjKH��jRID��e�PZ)�H��e&G""�P��i!tE�%e"�̉Yfd�Y
�4��9X\袒���\T�%(-Z��N��,��R1P���*�D�jĔ�Vt�*9J)e,�Ee���L�U9��fe�Ģ1i�#�Y&��#X�)0�2��CP8�Q�4�M	
��Ri!i���%u8FI�I��2e��Ȩ��u"6Ri�Z%�"�Yu1"�U��f��$%D��
sIj�,S��L-��)!J4.�"HJ�!�"iR���$�L�+��W)JI-��*�*%�VP�O���:�G���00�����;�C����[7�Cic�mD\:�K���͔:K�TU떆V��$/�}��}�Fl�M枸�����?O<	���~ ��W�z���^�e\TvHC�c��J��S\b�x��9�:{Z����9io�j�jߏ�'�%���f>�n��늌,����9����ܪ�YE���^�����Is�U�z��2%>�U�G[��'�����"�l<l��E)3�����0Q}|�[�x�L�|��q�N���5+]-�8l���rg�E�e�w���z׫��h_��E��YW֓��n���I�Q��&r��M"B;w���K��ӌ��i\Mɯ����,dpI*�p+;U��]��W*�Ew1-��֎�8޸��o�t��ʣ�2���a����T[Dc���v?��7�2�J"^r���������ʽٞ�ͮsͰ�F8�"&���uDu�4�%�/%��4Ϗ+���>�y�Ηa:q\�[��#Y����g6�51w3�f���o�1͵:T�����w�9�ޛ�җ(X7��,t�]f�T5Ct�7�9+&�i�+�FFY5%�y�,��m˺�%,M�\�l�ja�+c���y��+(�P� ���">��Yk����6ǵK��OL�u���%=dk���M�p��(B����[��H�����OTHN��@]�q�_V��z��ꌓy��y*\��6j�S��SVێj�c�	�r�Y�o�o�ZF���ѻ'��v�l9���i+ʌ�v�v|۾�\��|�x�R��K�U���J{-�hY6���9����lu���;�W�:���S��s-/=��e?uKIr{دJۺ������XU�v�p+dM�<�����T���~��5#�*�f�nX35�ɤ�H6g2U�eٽ�ȚNTk�/�5�Kw��"�+P�z*�-�7��hZ�[�e�v����*$q���u}jȞp���y�u}��}�[]��Ď;=�⽳����/��zד�|{� �7�8w�j)�%%��J\���q�Xbl���>�}G��3���e�1P�5&��j8fT�k��`*��!���>�V���V�y�f��]�
�C�G��+�yD�I�U� �c�˚z�4���dԨƭچb�Κ�zXk^@�v�}(��1Kr���z���ݧ
[XA�1��y�z7�8k��bf.�R�Y.m�L���ﾈ�7�Ք�F�[�9��[��ޟ��[��u��}�j�nM2@���8թ�Uf�-`�_�,)<��7ÂOKƹs�����IL�E��:��/"�^W#H���j@�k���P��?��n��O����\�a�)S;��|�Opڝ�c�ԙ���	:��~J��i�I{�4�S]u���>��s�뭽�۲���lT!(�J:e>���F'�e�k�h$�֞�}�Nm!do�r���e÷,��
�OTH.���s����cB����!���:mh��%L��L3�����m��7����������M[��b�jx���5��	�݊v�]h�$�R�
�Лpr�V	پ{Q���|U�fmĦcup��i��8���yU3��ã��e[׺�m�º���]���Dw>�m��Ӆ\N�X�D���<���e�*��Uj�
���wT0zc��.�ok<5��k����2G���-�&���.��ҸiŤ�o=V���7�䁿U���lŘ��j&ͱq�N�H�9i���i����U��T���+�ȕ1��5mdˇ�u��"C@���rؘ���j'��h��n׾�������y���7ڬm�ͨ��2��we�D�U��ܚ>��N�j�xk���OOB��ݰ�����w��>g2��c=j����~z� k�5�Ş�ҧEA��F�z���s���VyMh�;%��vGVe�>Қ��\Kf�ݘk>�v�[����M�����Z�h��w�هB�
�͞s���%w�����T�`W�+V��!��p��]i��o��n�L�����H\j�D��3+`(,���Ib��{�w:[ӽ�p��J�yfx�'�	W]<zZߦIYl����U��ߐ����VO1�K3#v�)�7��P��yv�{��4��r:��������wx��\,�u������ޭ3>���j��!���<�M�8tFFzz�%I�j�#w��b܃�4��֑����5���%�/%��5RQOlDU@� �b'�Ǥ�o�*�,�w�dw5v�]�_&�/zpƛ)��<���s�F�wW�$? ��%U�tY�C pK���1��v���.m��:�Y��h�������N�E�W\�su�J.�n��� Lτ��͑�Uy�/��}���٤�.�K�ʮ2���)�sA�j�N^Kq�!c��=��m/ ����;���{�����@�@}��^��yu�"����-p��-cl���qj�{��Z���Bˤ�NT�,�]����H�-��?t]�W���t$6�{v����e�aQȇ�:�UWB�)~ϬǵiM|�=��j���/N�oϛ7�n��g�lff\΍}��{)��}�B�u��4���<Gy���Z���:����^B���C�]�ڑ�Eg��v���1�t�8ViU���,�ý�ɧ	d늌,����.�՜���t)iy�yv^��"$I��c=���`�H�q���	d���[�xنqڳ{;*o)��6�����|�ݙ��ĕ�#���J�����=��+#��ysԳ+��#5폲�4T�PP>�U�ZOXp3M��U�i*�5�l��`;�6O�����JNmњ�U��y�Yz��{gp3�̮��7L(�#����*k�Fe
Z!w��qֆ+i�Ln�ú���v�it��8R����>��[JXS���2�J
C�a �LH�!��S�H*Y�KS����[Ž��q�A֧1��v�[o����' �̨��X�v檠��̤p��iF����� ����kG~�q�q��ۤ��T~$�	�w�Rt��wTΫ��/T�:�9�m,���bnv�t�<�t �����v3E�2���U�>u\u��aW��)���/%➂��6]պSb���_>���#)D>�R<�zes�H�S��|u�O*x$b�2�=����1[�6��2�嬫�l�]�u�a��:�G_pj��m�b�������ƣt�9���y��#�	���Ӌ�^+�=�e�՞#r�ؔ��w��{IS���j�BN�8t_����b�K18���;6~֍%�j����n;f{#y���ǐU3������0�&f3&�sa���q���+*�����~����N7y�|ƦZƯ��M��������o�rt���MR����B��3����Z�8�l*�*`YJ�c�`��c�1f�J״KCvz��\�>ɝ��t�L�`}���U�S_)��ʘ�+eYju��u�@xv�P��]���{sm�׉���l�&�m�}_}�W����R��}�2�ݸ�r��f��"i9Y:�,e�4f��=����t���\�g�VQDvK��XMg�9l�JN���ঘ����Iv=�W"���.�x��v{�����{`˨:�{چ�������r;i?�77���.����`7�z��D�Bʘ���f��l����ms�����M�Ds��5���4� [W�ܔ���p�v�⅝��U������ϗXw�7������Q�7�1�ڱĦd�w����F��T��r��.��8�a:��'%k=LL�8)iɶ���Nt�� P\u"���'^���A�F�0jj��8�.h��s؋ؗ�7	���⫈������uM֡����șw��qt����H�����6eÿ_�4>� ʧ-g���&C�g2�CY�&�f��ʸ�[�����B��}`[�;QN���t����k�NQ�w|�(l��Y�sp��C2�:@iw��z�Ƞ�����
���q;vJ����ͮXٶ0�]�Ȣ�V��Օ�I��i��r8�f�w��蛻	�o�F�}_}_I�{T������}eu�&�ٺ�I96�B�s�5��x��\wb+ήiW'����졧w6������7�>I�\-p��c�	Ⱥ�Z��$����������WF��E�/Tv�<��g!s�F��Jithkq�n(���(��gj'����P��'�UW-~KeY8J���=��Wm��!�)cV6���|��;�T�U����h�HUn9����鲶sY�V"����%��oDg�oR>#�����ڶ���W+F�z�?��rȝf�CrQnW���g���jY��U�Ij=}���EKԊ� �W��,�v�[�����9���_|�(P*���|��gA�L�D��ti��
�V�a�}��L�f�CE�j�!�W�qJ��鹹U�2h/�Q�i,�u�E7��$��	�
0�*��ȾQ����7	�����p�/س�^�a��KS'K�7�ЅQ5N��gs,��#嘯>��.�k�t�^"�QSnv)ٳQe[�}��!�͛3�7Z��}{�:��Ii�x����g=��Erc	�c�)��9����G�}�4�՝�QZp��c3��&����>���$��>��Y�n�n�<��j=�r��ry���{��!P\��yC�r+��yP4jmv��5��E����z�8K>����ݛM��C�2����I}z�J�F��,�ٍ,�P��;%���7q��:��D�e�R�!�H@i=�5����-<��jj'u�;�;�_�l�d�4�l�\$���n9������<O�uf��lM=�{"^P]���_V�ҋב��t�d�m�g���ڼ�����<P\����{K|�[�'�=K�ff��iu��i��ʞ��Q���:8�[��b�K3���zO��Kt�ͩ�|��"�<�8\��Yx����:-3CLnmAڥ/���l��������d�Vy��
V���r ��Y�Qnqޮ�N�?"���Uo�F��/f?z��2n���J�Nw)�<��]����	�ڏsV�cM��QޝNoU�B�k7��i#uy�=/!u14/fK���N��WLt4�\Ø��2�� fZ4XZdXn����u��>�1Պks�s�\�+�w�G(�Z��J�UU%3�6�&{go�:�����i�Y�*0��+-�;o�!Y���y9n����V'	V�]ϞZ�nʈ�˩�oZ��'���'[��E�Q4�gU:U��O�T�%�����@�����O�[���~�q-�dzU�l���J؟�FI����UFL�{�l�45=��x����WRM7�v�;��ML�Қ#��]�ou�:���]�ҹ�5��������g�<%��Y[8C���>}|�d�6w
֎��7���I\ܬĻ�3��N�D�Ⱦ�\�\�3������Y/9r{�~��@��#6�g����{4�	��;�%�du��~C��7�idKf[S���M�f���wkuweXΗ�y��.��	\�Ѥv�sڽ� 6������'�h�-�<�8��^}��
�T�HN���/��N6���u����5�Ev����}׫��;(�YP��)��*�dt��D�RI|)*�J�.�D�&�k��)^�j�)�=�*Զ�6�����-<���,m�/o#!���T잆�JO��t���*�j'��׫{�+�
���[f��T��4n�a�x�_pk5<6��2��m�Q��+��&Ӭ�H�Y[�g���Y�.�:��=���V-hs��7��=j	*#zX���-����|ή�Wfd��6򡆣ғ40X�V�Gh�cu�,V��ڙ;����d��%*{�����c�9�i�ƅk��󻝁�8���bf�tT1f3�.W!���.�s97{GJJ֖������9�^���vI����W�RŤ0���ٝ!%�de�W)]�վ�
�=�0�q�vPq��T�w���u��].L����ɴKW@�����NL���|S���X�t�r�.�q��ы��)���aR��P!�:��u�%��C������G��e3چ�����NB�in�a���r�4�����XU��-�l;]`�����U{�]N�I�Uy�5���wC�i�oA����Ud%.� ��G/l�ȯ{��纳��t�>���P�7�v�[��&-�&�9��a\(|ƕ���p�Cʗ�׵�.��LN�5��)�X��9z�DWpAF%�h�����X��P�ޒ�VoBlP��`�TK,��o�J�-hG�[x�X�(��f� 6�1!��ǭ������-�P୥G
�7Ɠ��j֊��v�"�8�<�]�\NHyt�գv�s:U1`��[��gB�v4�]�%��`�v�r���K+���XU���]���QU�,bU�!Y>�ԘY+�#�ZD���y')�ޖ��:4\\9Ns-�	��=;z���䢬��*X8�^�L��t�BǓ#�%�c1��`�D�U�{Q�
m��B�C�j땺���}u�^6#�*�l��|�^V�Dj:C����E��{I�[���X$��R��*#q+[i��[{8w7��W.Z�I=n�[ia�!T��7Vei�c���:j��g}�QU�.�x]+�%����;�oQ��XV;K)��"�f����*f�۶ɕ���r�����ڒev��Yee]����S4�A �G��&a�����(�]8��r���^Y�M#���;���'�m�Dч�'[��[��Y��#G�H��)���ツT��S�wb׌H�ǂ'�J+_;u�����Om;{���,Rh�u�Wv(1��M��v�rK4S�]]�/Tclj͙Y��'�\���E�^��&�t
*����j�	I����Еťx�񭾇�5a�G9*r]ʉ��!!������������j�-&wL�#6,^Y[@���1	OjR�V�ĺ�����>�	�6+�+���R}�BD<��;b�6~Y�kܱ����ήБuZU�f�gv�����!�8ҷvbB�-Z2�$��9FeV(�5eE��RjGM���s#J�s3eHQ�4��Y�J�23(,��)��J֢$��5��Y	%@E�EGd�ĢQ*Q9UF��i���ʬ�+Q1g@�4�gB��$-�#T#f
bjRU��W"5�h֑T��!Є�Ur�����ʹ��Qj������p��r�UgL"ꕩdV*�Y�h�J(R#Q"�%A+�5@�s�XU��b�D��C�����,[@�]XV�QGI�\&a�1�.RGI�38�g*�ؒEu�J�ڋL�VA����`�Q��N\��8DkB�D�Qq$���e�D�XT��sR���UPPHe���9�4*���"&EAETZ�R�a��7χ}�������R������[p_Y��qjAy�G 	Zsr�)�q��*xB�x����=IzJ�e�ו�ul����}��t��;�:[UF�4��ee���M&�\KĂ��%�䆡��6ۭ�ē�1�:8��\CʭX3T����-�CfU��ȝx{sKN�=�6��F�w��>*��̵�͎�jm�:���=;����q�N췳��V>��pꌷɪ��oɖ�"��PH�����d������:�ih�*��ŝ�y=p�q��t�9e��ys��&�W�u�����^�l���;v_�j�9��վ�ղ�3��Eg���rD���6UƤ�|��s���6�-L��˕��1Z��G�~���5�3��.cW%����{�˽��USl���4'[�.�4y"�O��.�S�9�\+W\���s��#\.�M>��f�Kk��F�ܔ�G�ۍS=@��$�.8$�XwM���q�GW+]XL�M�u�fu���KJf��+.�R�L0���3���k�e�}��Ζ7e3F��2�qޭ[w�U@IV�*lsq��D9ۻ��VF�Mr���\c�!�4a����kRLޡ��t�Z�O ޕ�Z�����E�'�n�M`�U�9z#��n%��
{>��5��
J]7[�|��ȸt�ߘ�ѓ���W?.�E,ť��J������]��L�X+�#�u@�^3;�Ef���~k����w'�/9�y���n�S(�M%q= &i�6��[75|R�o,1ˍ�K:Iq������6e�r�dH
�*z$���.b���<=���_�>��[\K�L;�7I'!��,�t%,*���k.�{=Q4�H����9@���m������7�!'uk\:M��w#�g�ko�K��U�8��5Ɍ}��lS�4�����ǐU3\L��|c���Y'�q�ԆR��d-�̪^ ���_��������=�d�GUe�Ư����s[�j� �2��~ͣ�2�����_�C��+*�(.�Ȓ����ͪ�)�;�Q���|�Wd&�7��<\�o�bu*���-W����N�+��)]Y��m����g6B��n-;WO.������xx�����M��d���oR+z�U���Q���\m�Շq��7t��#f�ʼ0v�ˏ4��u�C�T#���3sTg2̥���ko&Lţ�N�ʝ�U�Er��-���fz:ո
�|�76Qn�{}�f��м���Q���|N��[Ԓ�S������]:��	g���F�����&��e��!�q�SK���k�(�b`�w��Z��|=2Ú�x�$IJ�����ÓΔ
��n�k�(�%�q]���ܚ.d��|ʌ�Ib�7®�M�մP���a,�R��Yi醻\-�ӊ!RW7&���>���G��.�u�eY��<�Er���������N3Lcs��
�BU���Wh��<�u�����.H���Q'ig��ߥ�ͦ�m�J1��w=�}��q�J���Uf�}�7z��(�W����v���ȱ�b@�t�Љ#�!��]HF����>uyh�għq�m��I9t��.�I\5k��IY&;��v&�.z%vK��r>�/�#yu��^��{+ GNf��O���N�sg[�~�}Fz���n?S��)k-a���C�z.[n_�+��ISx�aķ�7Ս���I��k7۳m&�����^#I�Ķ;��`�`�|�£�7�i.��eW'Y�3�_����f=ν�I,{�pbSȔ�]�T�L���sϖ]s�4\���]g�o�+c�ޭy��2zb��fu%���r2���\Bn�|�ã�>���+Ѫ]N#q��旅>���С���\��S���QfSױ	�i�b74���wZ�P�	r��`����I�-��V^��9�<��hܨw��Bwݝ��3ѱ�Z�� �B�J.c}�}�<r�q��"iCY��,�U����EF5Z�v���ɿγ��X�;�_�����G.�UoZ��y�ȝnQQq6Y�׃-v��r'5-��ޤdg�k�#V4F.p�P�k^]r��BDǵy�/3sX�W���.q����n��C�� _=��x��\��f����sp�&2�@�Bָ9`�Rv/�}���Lc+�ZQV����9�O��3l�R/c�ߡ��Z���)v2����7���Ih�Muմ��2�m���Lj]�m�.��n$�w�as2p���uE�v��K7Ҕ��g1����Τ�b��ˉ[�7`Ss�z��	���0YN�k�.�<�K�ه`��͕��2�j�+6��S@G��]eҒ�.lWik%J�����ۦܲCGT��w�t��]7���q��L�m%/9v�}��9t,�|�S��p�m�����2��0�OH�\u���:1ʜ���Uʍ����b�÷��*��L��{jĔ���7��5M�V�U���ǂz\ROz&�F��)�e�n5�,��S�!;�9+��/-^Ee�;/9�7�={IS<z���TV�5i��.�����D��Suu7����j;8����D�[ϭŉ;���}C��V-ƞ���˞g���͸�����Q��h�o&����[��z��LoeTٙ�}���������d��
��4�w ��e���O<��}�1f�QD�Y�!e�^��X�e�\����5��4�����gry�\�H|�R{��[�Y�j��[̢;v_�暰��f
��z�<"�b�]S,0�xi�1N�K�:�v�;��:��"Ѣҡ���f�Gr�k%ke�=wh�+Vc�w4����C�5:�7cu�i�H�E)til3H�m]<��a�B)����*S�9���TGh6��e�շӎ�gL��w�������[���g!��Ϟ�3�m)�߁l����n�nJ�zY�zv�����w��k�����9�>�|z����R�Y�Nz���,�L�`D�7t�g�0+�j��97�����4������j�.�H\j�EO6f]|�%������7��OM?w�խQ�`�$��q��J���*_j���U�eE�)t������52GV�*饇|4�%����1nʫ�(�O�c��*�5�I\�6���T�-�k�;Y���Q���<<:ᶖK�o~�{�p�ؿ���Q��l�T(��꺊����}�8��{��#YeI�-D������_T��������^�;��y_�Wh�d���t�rCn9��!��jn�}o���9$K�r�;��@gw6�����ծ������ٻ/SNl��÷{H�YV�Dc�-Avd�u�
KF`%�Q�Ӧ��0ZSU��ѝI��6�47Z�8K��7)ު��Aʣ��I�p�{]pR��Hޱ��K;��֤�5{�J���ځuL
'�[IUܖ+&V��jx�t;A~Ƥ�ڼ���e���E�˔w0���1�������-պ�9��Zw��Y��i��p�,�z����g�(G8���+-%#�����ܝLg�"�x�|�A��}E�U�4a�7��l�v� sot���[�n�E���PPi��!�{6�����ݸ*'ڠ_�od�ʶskAH6s��k��+"u�A�\ [�X����9��is����k��2�;���K�9�پɧ	F�&477Qnq�}�
�v|��p�oH �G-��*�I��wt���%���F�����&�Bn�"�<�wU�jV�����C�
���T�AWti��0+V�d��AM�<�oO/F��,��}\������j{7&��5�P%��ZIu�TJqq������l���Rh8�[��}�_���	tM�?3�@��Ҏ)V��F�zsQ�t��Z�_�l�l�+��z��^\W�}',z{����!��H���&ťX;�7�*�R����Fk�R�f�Z̃�}K�rVJ4���3�u���ғò�o8�;n�
�b���1�yx���%�$f�[n�e.���ݩ�JC��
�n�,7^U������rD:$%�y7���8ޢN@M(w�(��6����0S�h��_61(<Mxʷ4Tt���Vm�7q�����Kf\;R�m�J�2�M_"��K�Y2��{*�Cw�_β����h;��t
���&Yq.��9;֯tn\۝�� }=���Y�������ݯ�(����y�ާ��9#��i��O�Zn9���x��~��f-���o�|����Ԧ�4u&��+�mz�\v�,��Y\��=��G��K�U����[Q,����>���qR��ԯk��T����ka����5�I�v�	Y���Lqݕz�}��e�M;������UE�u����bm��v�,�\%��qـ�9�T��mwD҆�'\VX�e��ӫkMjQ/v��G�@���kǏhJ�_��C{u��Z����|zw���nlE:Y֮�fe���z�F�^3�k)�A�$1� )��x�|V����l|-A���h���ut��\��4$vI�e �J]��ͻ��櫷���&�����.���+z9%�`,�)R�)���y�����v�$��� ߊr.��y���ȍYT���p~�p�]:\x��J�ot�%��p���|܍p��kl��k�}7&���
lt!��UJ��x�Z/��n����7b��g8k�\.�et�]7$U�jZ�U�&��-mQH���p���]Z�Sd_���c\��o_���K��4Ao;/W#�:��n"nM?���)��-b�婓���^r�q.1q�M�:��U�|ھ���aS�1����[� ,ձ�K���r���� |J��j.h��sܥ�SmdT+B�A�D�6Պ��i�k�x��ް|�+rb�q��l�0�2�[�y *@TAS��t�,��]pˁ� �|뫕>�
�m�����xں���Zn9�ˮx&��7�f,؎j�����l��ݘ��v����[�J7�'Z�®q�s�m<~�����ڃ��V"1Wꍝ�`nltn��C��P�|�VQ��8w8U���5(#D�	Z�%���R�^��5���q<�7qM���X؛��k6�˹+L��[�ce\0�n��f���GD�,v'���c�.�%Ŋ_L<�k�E\ʲ�ե4g�t�������P|��#<��9ś�G�o������7�Jv��~�Jm>���Q�˨V��:�ۼ�e}�W��RnC����r��C��5�j7��!�Q/�J홑��6T���X�s8��;-�;���r �Vv�R��,T�����<Ty�o���/G�_/}�Y��q��(�����;=�v�v���%����h���9GZ�C���
�S����nBm�v�`�����S�	����^��h�v�M}@�E�uѧ�s�V���}�ŮO�Q�@.�R��� �@��n]D2k�D����|���l�͜;��^ҫl�m���$�va�Ӣ�G��̓onc��(O��?p~�}6���Ե���v��'(8���^������XCP�P~J�\�	t����J�<�A�9+0�Z&��ʮ��{n:�V%AWE�գ�V=MWT�2˷��:�^�nJ��t�:�+��bN��f�f���������_-�n��RA.)�kL�G�TL���0��1����żR�%�fj�dr\�+����!��wYՋ���g�^�P�X�*P�Fqۮy%�K*�P�!*&I�u"��s�y������Zk1vH���g�M�k��}���Z.��<��S{b}������4^<3T� K}��e����tIHrr���k4m�p	���罠��Su|ˡ,�4��m!�,�s�kX' ���\Y�pV��nn2�P���KY}y��e+1-�H��v����n�b�y&��f����B�]A�Vz�:� ���)&��E��o �qf��[�m-����]aƝ�d����ٌ�b����䥳�Å̽��ۙ����[�+#<�w�xl+6<��^�s��"��n�vڥ�L��ڑM��[�o7��7:��2��XL���m�D�+���Ҵ��_d���ˣĴsGYh\��f����2n��Hr�֕�m�Z�a���s�؍`��jGZ��f��ۘCh}��,��XF�
�X{�=߭嵅ک������.�T��C����*��m�p性�t+��[i��<4�(n�EOo,��QB�j�XOCݨ���=U�,�ʌo�S��\���M	q`רE��er��Ӳ����$z�e�&�G*��F��U]N�\�l�����'jܼ�bB���Jm��� ewX2%���(u��Z�x/Ryѵ�(�]�3Ήy��%��q�� ��*U��H������(��F���
��2;��e�pW8�͑���4�L۷���d�7�+��P9�[y����ʕx��L��Sp���B����yѳ�G�Ӫ��؊X��9 ���r�l��9[5���˿�Wf#��}y݊�`����!��ї�I�V��g^�M���G++_�qW�s>U^�H����kV�tJfoܪ�V�ɿ�w'sz�8򩙬�U'�bp�f�DHTY�sVIѦ�;�85e>�z:��B��Ʒ;)��j_/�إ&ƙZ<��=/�⹲غj�����xV���[բP��Ŭ��eB��+E�:�n	�2��m#(�K�H���={[դ���6F�&H�%��f�n�	��Y��p�{W��Z�Uh�.��16`L[)�^���FQ���N��G�iV�Ջ7���i��3�B­S{�኱M�#dHf7�d
 osyN�z�i� �R���0҉ꗍ��陴��k6j��b�j�*(�j�F�}���4�u��h�\�#[��6�W]�iV$��Ug0m�dF��b�2���d���a	(.W%
y.�]�O��'��
���WE�ޗ0݄9�����Z�1>&��^q���\��ڱ�B����ð�k�`yo}���P�
�ZJ�G0��#S!#	3""�f�A��t�HDWe��PTG5t�iF�+�PDȮ��R�iXQDjIU� �"�9!�#H�	P�"�!$�(.R+H(�U�%e�\,0���5�2@�UQUJ���� �
�L��"�E8�C!D\����PԻ*�˜���I�BB
�L�"*L�L�R
T#��ȉP*�NUV(�PE
�\��#�Q�f	$N'1)V�r�"��V��#[ ��)D䪴;"F�QʹQs�5*VұJ���Y�m ���+8G(�L�*�D�"3+�\��Ȩ�)R�2�G0����E]R吆dJ�vTr	,DK5*��i�����J��-�Ad�˗L�:eY%�"9\�rN��\̺�BAD|S���,F�1Y94�k1�2յ&��:�zu�ctg��s�d��RU�5�J%����+s�vkf��Jf5���'(�ތ�G�du�M(w��̒�Cv�!(��JR���݇^��qz�8�uK�^Uô������W	�/>��^|�*@Vc(�wO.��E#SQ;�"w(w:�Gk�]|�m��I9��;1��M�'�[��(}�f��	=���=q/*:�-��+�lza�ێ6�Ʊ�ͺzS��.gќ\2�5*���b�^R��+�t�y�>6�;_7ze^�q�bĽeYE�vT�c�M#��ã��[��b�7�*<�g2�Ѓ�e%�C��G�ܺ�R�.k��0��1�&Z�j�߳O����v]٣��NK�v�M>�,�S<7dN"i�1�:0������q9Տ�eƻ���q}�	:�TL���Q!;�:��M8k"u����Qnr�ج�rƌb�x���^�1���/��}C�*��l�Z���޳+�(��D�Gl,�i�Y�E�]&�v�K�/7��.�]�gs8�ѳ���m)��t�a�7U+�����{��n�lюF�VT��nW	�EFt�3b�������V��ڗ���}N٧�c�?�dK9�F��g{թ�Żi��s�J���v���VSD=���τ�}aͥ��ƙ"L�=���]J�X<T�71���UFL�ޞ�F��Yl���ʡ(_���l�Y��VkyjԈ��1��+�����.���#���IEI/�<�+Dv���݁���X�A��Kp�'!��ȊL���+��z���:��ಜ{8�nu��M���p�ݝ�G�q��rig��ؗ�6�����	-�c�^��NH��g�x��H�j��/������E��[2޼�Z³(��O��/c�]�U3Ad��Aw=�:��G�>%;�h2D8Ga�
���Hھ|Y��]t�yK�n9�,��d/�U@���G�2��jj��at8y����d9G�(�c2�z{Խ79x�����2ɦ������m�Ԥ^O�~]�s��^�c5�B߫�1B�K�^�Kk�� �$�����X�C*a�'I�iV,1�`l����4�򐦶�'ݪtjZ�y�u'�1�����:��i���`�s��y����vLL��}�^�Nq��.��+�q%��٬�֣/{z[�;10���։,��X��!�O��F�h|��
���?��b��A�g��_gYx������y�[ǻ:�D�
Y���}�O�I�}9�7�Ee�D�s���e�-ν���M	S�a�l�+�S3!\As�*�YW��"iCY�0���Q��|C�N'�v�盚��b�vȍ{ZF�Go�/�hCV�����[*M^�Ͷ�uM��:���m.�K\�9��[퇉�v_`��=�n-L���H*���皡ݩ�(�[{=J��������{���m��v�Mq��J�흫�F�E<�/�%<x�9}��,�����_$�#�z#ި����ɶ8��RЪ�~q��qoM�ߗP0"Ib�$�u�ϩ�.o���������02��rgz#=l����R?�O��F��{��IYޒ�6�ɉD�ؾ��(�-v�y�uץ�Ǻo�a�BQ��J�z@/���}�!����w~��6�^ܺ�y�� Y�eSW�b��^�{�Mv<�fp��Ts7Zh��7(�r���VO%F�#�E�D��7�{�s�͆����h�]�S��h.�H��]%m�{f���r���r��]�7^`N:f�A�#�CD�J}��PݡI�B\ޑ�ӒF�NTx_���Z�jk�܀p��-�_���j���"o9*py+�\$]&̵�k�Y ,�ꐜq�y�%�f'سz��$�V�R��/�VA/�x�5N�5&�|��ؕ.��Ҏ�&Ɲ�y$b��\�߭��K|���yl{�wعë�z�F��ޚ7Ff�vo%�eo;�e罃��N3s�� S��6��F�w�� �d�I�u���n�o�C�eF��Gm#���iKKC�%>���+�	�W����Oq�'�a�Ce�����άx2ʝ�*"YF��U���#&59ے�N&�Gr�s��`²��;��Z'>9��6��в�O*Y���;u���R��s1�u��va���[���}���v<5��p`��B;�y�t���8�$.��]N���dpno5�	�s�i����HUua��>.e�����I��]�#��^���'���wZ��C��X����K��9�J�z��u�P���Ir���"�c�r>��Y���)�1�Z��nLR��Y�!F�O�k˛t�o���V��nd�l;��Z�' '5V�&5Ȯ�ܽ�M��3�6�&	�x����Y����F�����M�p���{+�6$��[��_pQ1��%�ҹ�5�s&���28$�u�S|�m�NPΔ�謴��Gc�oc3��*J���_��Uȭ[�:E�mc+i8��Y�.3��0����/�nv�!HJ?%��z�n:���z�x���j��	�c������Y/9���6�طl)�f6ka��әs���H�Цs��g��kYqV�2�%㗟,�;e�#��Zԕ���6�z�ԄnNK�[��Q+Oܘw�����t�8�dr�����kY^�m�>�g�^�Z�U�����{��(�=3eě/��4wG�X���/Q����m�lf�Z�����<)�����ër�����{c��^��Y���r��9��b�N���'uKQ�7ޖ��t�`���L�l�.o>�kl:����\=�,cn���@,�ǩC��d{�e�ۤ��	���r�^��R��+�@�L�R�ɝ�� O4�t�uT�#��<��ī5mv��7z��T)����n�w���Bf-����p��.A������0�8\���x��1��i��ͯ���.w|D����E��s�Z�K���Ț�''Tae��E��z�5�Nq��m����p�y"�\����C5i���쉥d�q�����;o������.�4������uFv�r���Q`�*[*CV���z�g��Ǝ$>}��:ʽ먮Ǽ��e���LZ��	Ԃ�:��ώ`Hr��2��9@U��qW��).h/s\7��Zi�|/��7$���@�R4�n�۽޸ٷ³�.�Q�n-g�����I�v�Zq��$W�����+'���u�c�I���_b�l"�_�Ȱ�9+�N7���H.��5x�%Z��i#�Sߙ�"]7�5�q�\I�	��/9���7V1�7������z��u�1LJ7��W=#�Y�6������Qjc�ǞM�Aw�յ釷���q{�#5�n��M�ض�]�.�)#V�-����:��s�KNf��<��Ј睻t�vf�Ay�$H�)�s�Z������m�ھk�p4/(��§Cm��S���h9=Ҟk}�e�J�.<�NO���sy;{���2�/��s�As���G����k��髧����D�燮����Kq�>Y�5OT��/*���t�FhV�bU�j�����J�{_<W	���I��~Y|�N&���&�ܣV�X׸thNY{�Z�<^��o��.p��>���<�V,W�̛����欣3n%gF��X� �3�����^|�����͎KEƌ����d=�A��2�nwl�Ee�M;�yEn2��1��!è�7�ks�s���g�,I%[4�J��U�7�x�J{��R��ꇒ7���\�$�l<������F���+
#��_�Ї*K}u[��E���u�y�����N�7�}�<L����݋S=PV�i�$�@����Xz��Ƿ�aA��p��o��񸛓fK�E�t���w�+U]��"�.��N�tf�]J��Q�2r�o��R�rD[��f��돗Rn� �nq�(!݈�	�C~�ۼJ�Ï��GX�rͥg��P��A-K>�}9�M�g\T�rgh�z�L5��'T��x�&eopW[���A���!����N�u�oae����>�p�f�]���.�����!�8�nz���P$�/�K_<�l���ұ��vl���v�*Й��3��¤�&�Q�����o�kv�q�������ζa\�jz[\3�}�������a��%W����꿣�٣���&�A-8�UÞwm���/"^)j�U�e�l�ʍ����oT;y����A�HT����S��E�l�R�kW
�O%C���Q1�P��u�izV.��VƝ��,����֋ן6��jsW��y/!�:���o��Z�^��[e�U���ً��������ē�0�ís��9��ņg_��=嶡);��\b1��=�]L���~H����&�^��I�����Μ�x��~ �)im촥����`[<�3|�/;]�����^b-C�ɰ-0�Pn�Ӣ���nN��{��q^Roc�N�ey�i��x\�qx-�	��^�l����%!j�q�2U�|L��c;��>W�L����%�����6eԧ&���^`���+`����Y���y5>F�FM"�a��Y�|��e�j��;:���v��e]t_,2k�YD4sg�l�.'\VXȅe��z�"D�AΨ������z�I�Y�����U/z�C���;7W��,�j�7%�C��;=��Zjf���+^cX
�(�"�̖9W�9�]:�P'EG���[��]��2viުY�Om�z訥�8�z���S=P�U��F����j��7�.����+	(��ꨮǦ[i�@�����Ca �q9+�5M���dW�d7�wp(��j�����I�E{�'������g��*���q#��&gʯ�e�v]�^�'w��:,w���N�,��z�:�GC�#7��=��b�T�-@��r|��^�{}�u�����"�ײ3��G4.'�lD���|7@������g�J�h(#�f=�,���#E�>*hA^�6&��B�>X�y
s��ʓ���X���,վ��W�,ϵ<�V�����$8��(���j���M���\��U�)�Q�U�Ϥ��{���K��p%7�;��m�w������]�J$�K�{[hU� �*����8��V"$�d�7��Jh�������
SFunE����1��l�w�k�[��Ք?V?�"�!��G��M-t���n;DZT���\��Y�*����绚��W.U�7^
�oQ�/}��_A�]H��0��20{nU�;����6祸�ꋔ�5bw^v������S﹫��������4i`���R80=�6Y;�E_��:��<�k��>�=�<��7�����{7=;	���}s>�[�sۗ'�(f�9'B�z}�"�m#ZN�3��������u��F��{G�
�PP�K��y�EvG�{����h�������͎�E��0Gz"��d�?W�f�a�)s���dq2-��|o�+���`���J��G���z�;��������v��t�No�(�8sׄl@�s>{=~�Y����&�����i��u����t������G�������P�H4�`�߬dw2�ğfL;v�;�$�㫊[��d�1>���������>�U�f��C# t���p��Z��o�:{����K��R8p�Q9ِ�>�hQީ��lw�e�����Eѕ�RN|�N$B�_��q�^�f �"J�~W눦*5s����a�6�'V��-;��5��VG�U��k��R2%�MI�-�c�&��Cr��yn:Zw�ݑ���}.i锶����]v�,Ʌ]u;��+m��j3Y�u,�w����G�!G]�ج,z�ZSWrL ��ú]bN7�a.�3{eoR�9�Hm<�KM���cZ��)v.���"�\�See���n��4R�l��w����������{C �R=�$���O 	����syV��aP�s�d��1!.�XK�Q��k���=;~��c�B�O�����ƛY|�����yWBHǺ���&�jN�S��q/iP�z[{�f�/�z��ֲc:��Nu��u�C&Қ��c��v��1��SSkU_�s��1�D�SѥV��e����(�D�����3�|\|�/��ML���X)����#1�X	�������e^�|�L
��
��
��Ϥ�f��ݘ�,�V��wd[]ר��4���yY�ե�pD�1e��৷\`W�~���z�Y7�
}�t)AK31��q-����̾��ܠ+bm+�\9���l༪���������g<tj��0��#b�fF�^�GCr̶gRJ_R�V7z$�e���f�Dt�j�Y��x`L�Ò�E˷-;���iWC�]c�����/��t!a]�-N�R�3��bMWw�,X
��A���[�V�սG�̻��nƳ�vh���gCm�O�lY����������0��.�e���;'z��ϕJâ ��D�Kd�2JC����h�*�
����g#����[���L�k7�bk"#m1��1��̺���Y��]%"RS�i��B�YY���s��fQ�n�k�|-i&f�7WfU��A�oaWB�v���U�S@
o��\'����`�R��ց�7W&9��L����z���FVn�u�ډ���d�|�r��Ԏ[��� ���z��HsUr�a�#�k�S8��dF�����A|�7���s�ͪx̬!��'f��	�X�ݽ�F�=��!F�ͫ�W,]ؗ*��#�z�VΌL��Th�n�$x�c�
�W�i�EV�@%ř4�d9%�շ�$XWT�u��K�m�0n�NL����J̋U��v�t����ѩc8�R�����v�w�{ܡ��o���.%D�`I�����m9]][r�L@n�	�)�Ni+�����np�3a#�O��{qܳۃʺ�f0K��[�3�W�5]n}��/%�o����M!�&�"�YJ�Z���˻�mҬ��5�\���i3L��srY�z��"mf�!J�E+X��LP�X�t��L/�B��;���ξ��謁c)^�xeE�c��Ru2��MEWx-9u��˱Iv5}*�"�=�#���U�ml۸�A)K�
u �%�x�y���c3����&�8�	��wK� �/��U�ԝ&�n䢁D���*�ݬ�$:�ӝLM
J�"�#�J4""L"
N$G*�\L�:fQ�N�Ȋ���U�Rt(��f�EQ($D�J2(��Aet��hAÜ��"�*�"�(��E2�"�"
�iQI&TQQ�DF�AVE%�hd�ȨP18W*9ª�9RF�$�h�('"Q*�Vfr�(�T� ��"��U���EDQs�Z!DEʊ�G$Ái���"���E�T��qVET�k9ʸs�W5�'�%ª9QQ�.DUG"(��I���G$��
�(���QTG"( �UșD嬋8�
QA�(���Ut�3�B�Y�x�E^0�MbUPEAQfUjQ�D٭���)1ȓ ���*�8��,iE�`E]R#�a9�9Qp��*r��Nj)�Y�4�C�ʈ��A(���~��'GT�KEh��ʵd�j�&�c�5���4�T]�7���6��e]e�lSW#8,����5�yb^wB�3�)0;oKE���B��,�B��˯���E��B�O�#c�R���,���y�H�.�=0�n@��5'���霩f;k�x���������o֦���HF�{�Ds�O�o��;I�V����)��VY����!S��	��t$Kf��u�5�FS*ԙ���{Ny�z�\;��>�����Xz@�jy�C�\U�Y7P�D�*��XŔ���/���,�3���F��4^j{�p{Em�'�8���å�4��U�`�EJ��v�♿X���G��n�@��$���G�9!j}�Wa�^����̟k���~̩
�nS# z�ulɑ�ɢ!��3և�>�hzW���L������݅�s>��޹��{�7�ڡj�!ڧ�ߪ.j�O�:��{g}>��g��A�~W��W�Ϗf�4�vD/��_�-��r(�����D�*}�..��yJU����R<��zV}=]>Ϫ�|:v;@4��4�����ll'�^��S>;���c�k4�j(��sG��똵Z�,�P;�1�����X���v��9���L�Ǒ���B���;+�]e_s�A��d�}f�fV��D�{���y�8R�m��,(�]�:�=Fb(e�sx�Fu�Apg,
��T�;���6�<\z�xj;���4��p,��;Ys��J��[-ط}�<oF.[,$�e�;�|gBKCS���]���v?S:��U��m���w����/�%b�C�~�^5��g͕�7���b�´�K2���g7yeO��������x��yFO�khv}�����Q�~�|�⽛����=��{=^v<��Ic~ِ�{��3�t�<}����,�����(���ю�*����δ��t����������˵us�Lsur��z��{�>��z��=�#�Ea	�oXS����~�*����BB�Nf%��Ӗ��y�]xdE�דY�������7�R��j0� F#웟QЅ^�r�0�(����|��O�|���ߪ� �6雮�W�fj}�{�:Q��aͿg��y�E����p^��x������:�\��e|���J��?�g����%�l��/7���wD�{$w+s/+��맀���'�=~ȫuA��-��hME/Y��~���K�~���3Z��,-���!pq?cc~��Z��=��g��ͺ�*�U:�NG©�]��욁��[�uou1>������m�cR�x1Q͛��?W�=��lC���V�Vn�8�jŨn�����\xd;�fzL,|�*��R�r)'�6]%|��F+xgZ����NU�E8U!���e�qť�G2M��Tqnފ��1I���:�Vm���ܘ�wI��$Ø0,
)lv�5������bS�>Zu,�i쫛��t��_���J�cSK�_�"�䭑�׻#��̱���2��'�t�c���9��GI��P��q@�=$!���9��pΜv�/xߤ�5���[���r��׺�s�:�yev��F�VE�_��ã���5�����U�;���ڐw�8�ӚǆQ��������]Ng�}�+������~Us\\ITA��e(�+2GP���U��������p���ŀǡ�s7�Y��w~>��o�Y��l��hjF���^�dV��cW�{���^��y�����蓫�=Cb��`g�+��pJW�^��"�ݓ��g��Oo��q�#�UӷT����yu�S�J�K��H�Nׇ���׼�\wh���݁�޿sN�CZ��qvyW�{���!�hH6+��E�]��w4럪�=~�9��=n{��wW5u��{���}�vuצUp���5ŏĘ��^ҏ��-ۊn�\ܘ��N<0t����*��e�>����\�8��|F�z���� �C�!+�a��U�l����\mK;9�r�.պ $vdFs�vtk����ּC�Rx�bܚ�nႍ��v�� 6��[�:W���M7'���&�M�u�^а^�ff���X�ޒ�fκ#"fйD�<�dxr]��0�/���nfV���t��Q�E`{ڰ�ZP����'��E{���~aw��3�do���v��D����*��G"_%�Ń�l�F��9B���࡜��+=~Ć�]����fF��'|)�p�0��k/y��*Oy�R1�{^��%jFM=�1E��>O�؉�����2��3|���O\cq��u{�〻�=�*}�U�g�.�,�bCB�V;D�)ϲ;�*N&��#��xw��Y��>�5[�oq����7�;��4�bMT/dM-t���}��{�V��~ʟJ�������ڪ�����WW�}�q�*�ޯL�;���캑j����d`��]5}�c����^�כS;J��ͯRʌ�I�����{޼����3�ϟ��4k>�L=�4��:�pz;���B'p�9i�턼9�4<����
��y~�'w�5�\ϭW�TWn\����S�¶r�=���]_)�凷�;�����^琚���O� �,�o���G�s�/�y�]�~��(���}c�D����W8���/<t��B���;"�ӷ��yW{��E��U<����t�~��=����qxi6-yb��_��Ql�II��(ޜI�h�R���D��FY�O˽w3=����	���r��Y1f^��;�q�.95�9�kF�r:X/������j9
(Ղ��JoLe^X:݂�P�O)�F�-MÎ�2�3�'Y��U�V�������ו\��qȢ��Y���L�����"�j��c�{O�⯺�i�����Z�F��qiۮY*��F��˿Xώ;�n�����5��^����qK�c�A�	ȍq^��~�O�ǳ�H�3��� ���,R�va��{��M�ou��>�׳�ݎ��w"�Ϟ{2����n��WC�I߫,�ȉA�
��N5��^�>�|	>ٟO��s�e�=:�]xe��"�w�z����ީ`�o�	�ul8������9#=̟J\qo���e�
g>���0�l9f�Qo֦���HF���C���@�1X/;{{|��p7�vEM���2��X��١8iߘ�(�eZ�*)�����8�}Cy�׫;����<w���=^���(0�麆�&�Q�j�B�hx���)Z�U����>K�n��T���%�G�hlD��Xu�ɗN⒦��T��n.��Xq�˛}@�ОpGx�y�õ�	||��r#�W�1�~���zf{�!����eH�^&�K��"K[vo�3�����6R��Z�v{ԞuYt�.�vRT�&	��i�ڗR<�x5%ꌞ˰��S�3z�{Kҭ����lJ���"&wϛ�奷���� g*/�	3�vU�'J�57��)Lp��0(D��*оK�tX�b���E�XJ�NI�4�r�[+OW��)���X�
8׈/�q��<��S.����2|��z��OG�a�7��.C�	=zVD�l�9h�&���?��z���#��/���n=Y)1�6���+��|��u}�mE�/�s�q��9z�7���X� xӟ8ӋcӮ�ݱ�=��v.ڼ��Z;I��ymw
��ނ�&�u��혵CW%�P�����ŁK���{]36)KO�����5c}������e��^I#~��f��u�Kw�T=<�,��4IU^)�w�Sdr��>��33���T�����O��x���{fo�5�:��	xEw���^���,W����(o��g��̱���$�������K���p��,��tep�>�K�b�Y�8^���=Y.��×n�3�錎n�^��p��T�>�����<��S��a-k<z�\G�F�܎� إ3Q#�9ώ[{���׆_�y5����>�S��4��z=���8�<O������X�<����>W�3R�T�t�g,϶/��5<q���S(@�z���b���[�6ü^a�����շ8f���AFc5:�*T��FM�mr�9��9K�PV�Ćѭt����0sgl��s[��b���Q�xK:�|ݙ�{�b���ms�ó��PQE����H�v�bɬ�f�\�1=��(謿9�r����x����w>��ɒy�$ Gt�U��ٸ��?)�Ll�r����Eh���S�W��Ώm�?Y�}������"�֡2ؒ�)��&;�§�k�-�\��4ݏA�l#��hTq�?cc`{֤xh�ۑ�w�7�b�U:�L�{P�]���$�y�MEq�7�,� ga*~�Bয�|�^@xl@�z{��f�wn��f)��މ�wg�UT���s���.s��~"�+dd5�g��,FD&���f�*�l��� �}��y����D�U��c�(C���״E��Ξ�^�o�q�͗#���׉���yמe��U����u��sG={77�n����ʆ`wG�gpV��d����'Ђ������z#=s��9��_���>��/�ɮ�3������d���R܎��׾.�Eϛ�ïτ����ϣ��=;�Us���;����gմ79:���ԩ�^Y���iw�Ǉ��n�t�����oW�zv��`d<�0_��*��>J}�޾1^���1;&�Gk�����O�-���{8e����5+v5�QnQ�Yϭ�d��s�C94�����Bm�c��g[e_�f����1��9	��7���#��:��<��QL�V6m*���5F�b+dBSD3R��|���12:$�w���q:L�����kc�����;G����xzv#�^�9[���G>��+̾j���'�W�F���тe
}��!ɺ�X�匎~���=~�>��VU�k+�I�����)��}��b=��|"�cP��@k���#K��+�/V�t�.h_���y�+��[��]��;�^���\�/����*&�pC �T(�W�]����U��4��k�G2)�~9��{���y���ddo���w���%}�N����B��5�/o�ZG�w�g�d�}�Mo��;ƣޯY#��x"��g�bw��+ݞ� ���7�zw;���5�{�C(zP��]#xR���D1E�B~��O��a��t�}��ߚ��+�w�ol�9W���uc7���R��d�C�������hg��c��N��kT�n}�Yl`��/}묠�����f�J��f�����30�����������r��<�T�Y̹�~w�2=������~˩
�&=��3}���zW����j�O8"�O�zh�'�(
)'AP�7���t8���S�u�+���4����	Ԙ�c���'N3,�mb"�]d;h���ޘh�C1����X��U7l��M �RΡ��q���[�ef!F�#^k��J�TZ��P��AZo}l;���t���q�~���z�}y��zd�YW<�F�i�둲Ȩ�v��{G{;�\��g��|m��{)!�;�����+��6����lx����͑�eά7�hu�U�wǼ���#�:�9��t�����B�d�?�ز=���zy����Փ9]�1��g�z��=���̏�q�"?	ѷ�R�q?����w�:f�~ ��3��#ҝ�g����@������=!������F<������ʉ!I�U�E���L��1踱�nF�ޜƷطM\�d����㑿{/��)�>{QY�u�00<s�E�7�����z��)�zVnM�Q�9ze/I9���	��^�����z�O��VY��Gn��� p�9�*���?�,;X�ye_X;���z���;�|=���C#!�ߤ�Ee�Y# ^�����9�1���q�˭(���)���ps�����g.�+ި�o=�W�|�}�Y�~��p�q��p��^�7�H�_�L�Hs9��.8RAN�#�|6߭Mg��b���؈W>�q��I?��8<�;�P�j���*��A߭��5���	e���d�F��-h���,���l
�6�'X��}ي��5��IN�\%&��͹FK�eJ1��N4�uړ�����{eS���:��8�	� ��̗5x�tu�E!��}$iy�ݱ�
&e.�"[4'`�y�B�J>�&e��}m{�&}�u��2����|;^)���޸=���[Y"�@��^�c �4<J�p��{�3�)��]��A�i9Sӑ���t{ր�ϫe�鹝V�(���
��GP���k��0,��M^^��d7cݔ�7��C���..7�ۿH��O��2}��f�ؑPi�`����'�W����X��h��l�r����6��da~�l{�2�}���c��d�b�K���S�[����;e�C�-�UC�Q(N|��+����;L�־矸���وC>���n1i��U�q��sW�ܣ��勄=��g�v'kedU����X� w�6�������O�56U	#�o5�[�WK�︫L>�+ɣ�׳���ع,�P�f!**~�a��[Ͼ���]f	�w�����
�~���j]S�#�C���?^I#`���m����l�����=�c�#���;Țf�z����%�W�dƯ/mN���P�e�ᐼ��yFs�PӔ���}�+~ǌ�ݡ��^���	2�۸��å��B=��[�Q��S�ߛ^�ň�p&�3���^���V��)��"S�F ���o������Ty�6�϶>׺��1P����I�o��̡��7+`�%5�M7՛����a�'!B��{v�0���ֻM��� `�#%<��_$h��M�oe^J͛�({/0B�^J�m�S�)/��N�13&j���yY� �ZsX�n�\e�b���ɻ�]𖶸����(�S�J��O�9�«���w-WKhe��jk·�l��B�jՋN�WrٔR��7������i�dWB�jY���c��Ͷˡ��f��o.�|��h��앳�9��T�ޒ���]�Jhlv���AM�Z�����.��/�+���-�����㚶kR�nLyd�C]^p�E��Bu �y��G3�f;l�&���{0�0*&�VՎ,�"�u�8�6�í���A����֌}�sy'w������$��t�B�Xw��]usa�I;3���[��V�E'uֵb֥�.�UK��+�С.=��_f���i��}l��K�v���'k�����2�]Ry�s�.�7U'c�
�η�����f�m3u��ָ뺔��J�EBnWcxoڀ1&���:x3�_�G�Z;ws��V��)E̔
�إ�2�xLI�t�Kk�}�Rl�$�g:�W�X{@
Ry�K"�؝�O'x�:Eu[->4��x���t�իo�g7�PE�]�)�N'x�����&A�4�w�6'|BjJ؍E������׹�k��w˸�v��#c�5
��7\�HX<�P�4��"��Rc.�ӛ���X��)�z�5/s�6�;g�B�a��7��8�1�W�f-.GB�~�����v�����~�w��	����<W�ڕ�U׌ۉ��S�8�k�Kee��F�P]]�$��ݣ\Wۧz�Ԧ-9.�xK�J��pɆ^
�pΔ���7����m��++��2a��Ӥ�Z ��Wb���+S��moTx������򅺔o�P!��nv+� 0t�ӵ:��r��OsS�O��ƭv�}x�����x\�72V˓���ff�#WG�+%Ij�xm�qf�V����A�J�7��֑9m=�E�|$�3T�xv�9(�5��u��l�ԥE��} �.�5a�9:�or�[�z�v��N�ǹl�x��Q��gd�۾s�Nf�t���U^�}��E�]�[�t�V�T9���czlY�r��wyyYE���`�����'OCv&e�F� �(h�G�o����Lf���`tK;Aa"���n<M8�d$p(>��[w�p�X�1����v�Dnu�0&�39�����q��RR�hsj,B�v���9���ݥ��m�V8����	/��w�*&�۩o�"vW|��r
�F��ݜMa:�ك����#���G�;�����v�Q�!�t ��
���\�8�*ʈԉ�V�*�S��2�W+�"T.G9Ȃ(�T�'j!�rТ�*�q�a2�"��(�
��S*"�څ�$�V���2i�K�� ��"9N#Y3�Uj,�����	r�����!D�(��#�:K �EDj&\��p��MȋLNAs�r�W&�)\��Er��"�1�D\*4B#�dQQd�
��YE�'r�QTUU� ��"(�9r���"IeQ�"58fTEʢ�Q��&u�r*�"�9U� �����dDr(��ʮW-iE�#�TDDUEDh���Q�"�\"��ET� ��es�EI�%r�T���PA��( >N��PoNL�U[��vY�WG��U�-�(�WF]Ġ�C�q�mJ	EC�"xl�%_R�8��,=l�W$�d_���_�L��	�h�z%��뇑=���/�nC�[ő��9�2����n�5�Gz��Y�����>iA�%_�ko�U����1ނ=~��T�=��{�+�i���9�K��\�t��߅w�QX�r��H}��*s5<������,˦2;ɼ+��3t�ތ5�[`J�m��ǖwUE{�ڪP�yd3"؆br�L�Hs9!/UNA�m�7Q�:%x>~�S�m�/y��\���^t���A�����p�\,�����
��|��3��v���¼y��.0��0wЅ�C��q>�>o�~�$��N���
�T�HH�-Dٕ��)O����<'վ���]$=���C9�pq?cc`z���~�r3�;ٛ��1A��jc�I����� .}��<�%~��Ym:�?�!prY�����W��;g�&���Xp���W���W�$~:|���K������.Ws�׮=�{�2�n޿GV��u�'v�T�z�v��,z7�ė���>�@d �7����¶��U�3~Ԟ��1�i!ulkǘ�H����h��m.�1pߩ:�s�Uە6���` N��������)[;��]�Oۙ�1J�ߙY�ۏ=}Aj��9�g��76\��s6g��
N��Y7/!�Daܮ�W1����j�,�&pR��'b�AJ�]��T�[�v��Գ���Iub�J�F���u�~�4s׳s|��o��Ug+΂B���R�p��L�K h��<��~��������N��ߐg�>Ǎ��`�^ʩ�����D/s�^�"��V{k���xk����^ p�i��o�zv!�ߏ����ly��dv_M��m��rշ��*�3�)d����O����`!�i�ޯ<��^}���pNzfb�"��my3	VM�# Sq�AȪ����Y/� ө���/���1;^���6z+�W�y��{:`{H�Ga�'}z�\F���s3�!O��!������c>�~��s��=������^�+��>����^�/�q�PQ8��r�5P�KJ���ڙs��-�����Yu����:R��^��{�Ν�E{ö#�s,�[�pU�
���E���B�XK~��'Ö�峞S��e"������o=�W���\�#|�N�v���0�zab^q��K�39U�)�z̃#�3pP�~Y���$4:�G?WI���O/_��"�4�=��
{}���sR�(Cʿ{՛�]y8��"�O�F�c�$��6�y�7\�V����*����:-�84Q52¨����	\��u^�yY6��FT��	���n���e�6٫	�*�r�e���+s��b&��w���e�rO�e܎X)���j��(3��,!�Z���aW�/�`���#h>���8ث��ۛ��qRqi�
7�^��<��Y�R�W@���"M��"��+>��>ϻ�*Nwy��(��n�C�ŝə��dǷ���>�~�ȕJ�L�9�5P��GD\S7��xW�{{R�û����-��C=�t��2ٻ��6��g�^�>ב�Q�u"�0�H�E�=��W����b��;tK]�^hye{��������U�O�s>���=2F,���R,��Q�
:g[�'s�e�u����?}��wY^C�t|Ux�=���W��3���~;qG>��ϙ�7�$lY{ _��#xR�X6B���OWO�*�=8���!�3ز<�W�z_�a^��q��9��ڊF*�Q�~���hϐ�uN\����w�:v��B�s:��=:���6��\���j����dz;/�>�BO�
ڮ�ۈ��	�r��%���Án�|�=�Υ�y�ݹ��K2���}��b�9潞���xt��{Q�uZ7�\��J� (�D�����FMN]Y~�?y1�a��}U�F�<@��OW�y|�fR�،�q�<R��E�[��g�ג5~��)Ց}۾T"�O�ݜ�O�;ǎ�g�x�:�Qۥd�x��ǡa)C�ĥ�Ԗt�}���oj5��KKp	ڣ�����13�m)�f%�Fb9�ʏ޵����۷�>̘}>���<�������>��Ee���Gn��0�(���U1���Z��|�z�Ͻ�jǖTsy��_�oz����{!���������$�1�_�^g�oU�V���r ��#Q�촃�n�½���{���O�#{�,C q�yo��vl��^�H�Վ��O�,?���#��	�+�9���^��
L#�|6-���E{ئ5�g2ț9WR&Yֻ}ŗ�;����x��}끾�b���P&R���H��	ߍW��#d�9LO�������~�$�Q݁����Q/=;�����?Wp������Mox��&5 �Ѳ�n�J=q�y�5^��V{���ao��W�9SӅ{��`{ր�ϫe��2�\Q�R�9ʌ�qb����ܣ}����^���{)�oR���A����ۿH��O��2|�&{�v$G�a�5��=���<���)X>�U���ٺ&�sn�cada~�o��,d>�K��޹����-L��~Y;K��,��Aj��J2��D��V�g`�Y��5��7!��#���۬?y=ɜY5{��$!F�V�Y�:j��Ŝ�����x��ߥ��"`��3��qs�$6�����;���O�G{�յ��b[VEp�;EW;��#�l�Jn���Vn�Ԍ�`v���\T�I��\є��w��Hu����̒I��%�F�A�����bmq5!ԆW磿R{A��:��#��`z�v��D�l���xt�,v�<iϪ}��w^
�d*^X��a�d�U�������g�sF7"���LR�b�(�b+/�7�y��ˋ�=���Wd���)���,��;�g�l?Yal?^I#Nћ���M�܈F�\L�9��Ȫ���-�w/Ѿ�����t��bz�3:���.����\>��'~��f�Mm>ݞm���*R�^BZ�U�@����=�س,a��KbO������xx��܇��L��l����G��.?"�?��_��𻈓_����=m�j����7[ߝ��=~���q�a@En����^!�;!��EjfJi��Y�Q��+�׶�g�~Y�Lc�y7������˼��k(�Gn���r�ns��K����lC3��&|�9�����>5M���ތW�`��Q�pqޢs�R=�^Ʉ���>������ڸY���&'���ʺM�����3~Db��*����(ds�ȟyZ������fH������p'���L�~#�[{t��5�5��Tg����L��!�j��;]vƱ���.�b�i��tj�&N����]5*��ɹ�F��p1���#ԮP��WJ�B�_mf����(e�B��JBuĮ��瀗��/T�:�eܺ.�;+-A��i��f�����z��t#��4W�\9�Q������3��nFG���W�<����c<[��v{�W��M�*��MS��o[@ΥO�>�!pq5����^@xu�(�U/]��7yٻ��Oŏ�&r�?D��<bҕ~�X��]�s���,�l���q�sn=5�Kv����IM����{x�3ޯD�k��#�(�A�n>��g"k�#���$�{>�*]�5Z�ٸ��)^Tg�O��fɝ���s���>�����ϕ���s۩�S��������1����6�x6:�x�a���+=&p�nzu;� Ϫ|,��&�<>>۩���}5@�����(�*�>��-T?U�y�t�7�i�a�Y��w~>��~�^u���\Wgݹ�wK<G�{ה{	�x�.�*�m9;*��ǫ��^�b���5Jけo�t��|���3���u	s�����*�Z��}
����]+�h�Nv���+>9~�g`[���uzV}������_�f���a��H�qW�u�d{��cز	�z�\iۮ���)�܊!�A˿X6�Xq�k{;K�V����R�x�z�$��cΠM�H�S��wT�ّ.�wK�WѢ�T��F�Q-������!ȋԽf�{.��S]ύ$n8�"JauG&"�oQ:��	`�����i��Fpٽh�Yۓm�GH����B}2�V m��bi�<���@M��p7�����{_��}���Eah�����~����N,�c9�Hg�W���y�ɇ�{�ӽ�xv�z�Y�~�>#b+(���\%�&۰�'�~���m�n�[��~��^����s"�2/�9�M�l/T��؎�̲3|�O:�/��=�
����_%�Eo��S2�]4�H23y%�~Y���$6��Ds�O�6��4���zyp���"�Q2�_W�Hn��"����b��sV�m?cb4S�#gվ�/u�z��^߻G�<?{ vz�¦��� ]CphN�^Ur����#��Q���ɘ1�u��iq;�s�9�̶֥l1����\lMC�u3p��nj�{>�: 3^���KT��R�qY豻<o�4z�ź�ԥx��O�>��e�n��O��'���٨~˩��o�,���zyO��E]�sieq���Խ���<6>����9#!�vz}�WaC�\ϯ��${a���mԇ@w_��eף7�z�,��|�|:�^XH؃��<�C�;o.^�#���}j�>�ۊ-rq^��3/&�h[�o�"+]�\��z���O�Ե%E�WY�Ӡ��1�G��-�{eZ	سi�N{r�[cj��2�K�˶�~r�ğ���$Jg�VC�w��c6�S�$�Dn���x
�Ki��(+�1�'7�
���z�2>o"��s��U����X�r��K5{��Ֆ�qö�ǽ��zd<u�_��{k���^�p�=��"�~��q~b�d!����W���WKʻ�:-_�;Q�2���������>��t���FϾ�/��e�a��I�zDo���D ��υCۚ�U�YPX|�5{|�sɕ/L��ff�}�^;��6#�~�;-I#^ћ�;u�00<��G���Ӫ��:��)'�g��̱�{���I�d���	��\�����f)����7���ӵ����v������ ����(�9V�=[w4�}��C؂=~����x׭S��Z�X�j�8zB�W��D� �z���R��*���ǧa���ȿz�h�~���|U�(wE4:5y�|�
'�C�����+y#$!jϕ�s0��"�Y��~���E��a�q�ي��:�D�(��K�:��>��s��{ vG�؇�L�X����j��w��U8�J��мuE��N�q�J����9��{NzOC��F���z�qWPad���&���y�>�"yh"z��;�������G����[F]k�bdӫ'�Q�3"ᖑ��V�u�;/xx�ڴ�\�(҄�]&���Y��ތjd��J|-�b<�o=�[�+`�r��K���xu@p崕7��5gq�gdKUt�d�bI�璛wݬ���.�^v?D��=�p^G5�&S�.�hl��Xc&y�ȫT��nц~����О�SF�>2��|=Bk��n�B���a9�#�bද����H�ϯ�2}��dG�����>�#��yĲNw��z:���RC���齺^`�T����֮�3�}K�X�Z�|��ΕsƊ���#"{�'��ɶ=�A�U��'>��l��9h�;�k=7�o�d��Ϟ�]��z7ތWyw۽�6�}hF�V���h�z�����,��k'���]��N�v�-i��y�;�+�����wfl�����g�|�9׳sp��Z3����7�>»�^������G�_�@��#�!����v�g�a���w�ּ�\�h���۩�T��%@�1��_s���K�c�<���Ț�'��]��O){�6=��[��)eq�tT�~��x��^_�ge�v���KB����X���"9���t��kˆ�~�G�k�g�j�֩E(�-�/"�t_�ȓ\?Q0{>����_����Y�W�_��Tcƴ^�vC�3�RtX�U�\��J�VL�xkol*�=O�xlT�=\��Xݫ�9��.�c$U�r��or����^���e\���w�$T��)����m�_^j����ga�h%�U�V��[ch�2�!�w�7�䍮�L�&�˴�C�7�ݣ[�Q:���M���i��n�ܔV�v�5�Њ��Q�ǁ_5�f��Cݺb��8[B�H��rw˲(���R�I�>�[���\�q��x������< W��DHK�R7��]�rǛ�Mz0����D#����3S�M�:w��0� ����Z�������Bb|��i��9D����Y����z�g��@�k��!��Ȭ�_��߃���~�$�z��G���y�N������i��A׾�2����5^vda��9��4.}	�=ZG�'�["��l�}*��lX�'���������#�<*��@&0]~c�5O֦�[@��B��w��9�k=`wq�>�}W;_��J�r��@���^�ӫuU7��!zd����\��E�BVȮ M�K���uW{t�=�9�^��s,F??`��D������^�@_�0��G���¶��>vW%��1~������ڽC�҂��כ�o�|��\���s�|��>��~�MY5<�A���v���r߽�ew\tb<�p�}��$3����f�S��Ϯ|-o�l�ڹ>ʡ{_~��4�Ar֛���oβv��_^�� �ಝu1���Uʆ�K��Zңb���mK��.���Y-L�WK���\D��%�����OQ�1���Q���pkҬ���.6�X�º��n�3�9b%F�+Γ�R՗ɬ$��7���R�% }G]�p����v�cܛ8Z��p�F���J��V��[���@�;���f*b��U�3[�0ՠ��ZAoy��t/�cxJ�)A����gIV�Ii.��uf-�����J�D9�9Y߷1�-t��}��D4�TMü)��qs3�O�M��x-�5i�������)A��W�#j��.�ݫVZ�)o�%f�z� :o	V@�:��b�ct��	9Sӝ�W-�kl<�2i-Ш��2�n�,oY�Ԗmir�~gt����+R9�UZ�E��0��	�+|*�������*�g�s-�v�����N�eMd�IF��۪�B��+j��rه��{êfr�����ԯ�H�e�"�B�{��J(�wiP�˺2F�eX5����8E�e��d�����蛹N��:mD���'6��p6�X�ށ�)H�ut���%�K/h�<�b���W-� /���vV���)f��q����U������b��鯶�u�=%N,Xsk`��r��]�F#usQ,V���05��:*�k��M��x������0T�k6�mMY����±I$���-a�A���t1J$����µ0�|���v��K`�~C׮���qb �]^0_�IjE�����u���}��w��T(��W�W��5݄��[oß@�ptMk�#��:]o'�nr{�+�WQ�M8��cO�]�H6�����y�������<;��}�����v-������td\'T��Nsyt����M�}M��/�j���X�=aѼ{��a�an�;|����-QW-	�];��l)wz����d�6Tt}�p4%Z���;,���,���c3������Co�Jg����o���"�WrGR�ҳ:���w�mF�d�f����i��n�=K|�h�b�R	���o%b��s[t�u\v"�{��6����]���%ֱ�`�E[Ԣ��wи�%XΨ��r�lvԸ�Ef��k1nm�5�\�|�%+�9Kn?j=5Кke�ʋVZ/ti���k.NL�X��[R�����D2���֎v���#���z%<���2�'��#h���A�B�B
fX�(����1��Sմ��b�!idYo3D��Vd,�;����6�VP�d#�e�*��l��Xskv�A��勬��@�� �!9jݼ�%��O׎.�D�9ґf��	o����痗��pi����C[+SK& ٘��q�-�qB��ӡ����e�-��y=���I����a�����#����R��ڎӳF;����p':{07�2��(   U
C�T("��UG&E��+�.QQIĂ��r�K�QTEUr�ȣ�Dp�ET\���Q����o��9G"�EE���EE7���Q��"5��Q2�EQ*9QDW(��\��e2��8�r��FVEs�D��DDEʮ��ˑATS*�Q����������AAETG$���UG9U�"����Ȏ���ʈ�TAG""�FQGer�EAeE�8E�9r�"��-i\��QE��EE�(� ��Ȫ��e�*
�(�*��9U��BW�A���*
�eENA�NA\��E\��r9G!"����ǟ������������,�\&��Ozu�a�y{nv��Mq��A�gn6@P!+9�X��z�b���VwR�۝U{�ƽ�$��
�z�,�E��]�Za~�g��W��J!��y����xz9g�QE�9W����ܽ[��P��}�YIڅ�aꉺ�V��5~Y���Kv�<����%~U��/9[�OH���M�&���{j�qz�ʧ; Zr����w>u��J����&^��%��M\�d��()��~�:�d�;�"�N�pȌ,�S���C���~��75�r�=�}4y�GX��AGu\�G_�Nk�_�����=���E���!� ��*��Pi��-����N�gFyO�]���n�W�=ɇ�{�ӿw����޹�q�����wY�M��,�Y�hiή_�LR6@�
&��3&��D3�����o=�xO�s��̲7ʄ�1�׻�^%g(�f��s�# 7��^��e����l6j�Q��+#��Hl]���l�b�Z���]B}$jx'�[p�1j��+�&��22��繊(dG5jU���_\�5ờ�� {Eo�xּ^=G�ϟ��;#�~7�TІ�$ؚ����!c��v/�6y|s�o@�'��bJ�"箹�Be�����x.�G8�o�=J�N�H[;�����Sڅ]ް}!ަ�X:2�Zv*y�TA9Ip�%m�=]����ZܻW�A��NALq�3�^g��3�]��'.I��vj먏"e��$�*J��9�;�BԔ]*�t�G%�'�W�r�{���V�Ǯ6&����T�75P��GD+͞w��Wf�םF�6jW�5�cݔ���j�� ��O�#�Y�-���3��#f�~˩�*`Y'�vb~](����3�=�qu�����K���q�d5�J�y�Xϟz�}x���#���r)���F\���}x�u�����D�8ul�~�ì2<C���dA�܆���L��}j�G������g�����9l>?�,�����8�:ƭ����7���Dq��{G�\�j�Uݜg�YU�u~���*�0��2(�߯x[��������?�����Yх���盝�ǽ����άE{�sud)�z׳�7�|��~��Ma�ʭ
`wg¡� 扺r���oz�og�̏W2^�_�o�^��R�z�!�/�^Z�F��3zv�``yv��.ɏ��Y۬��r�.�=�J���ݎ9�obO�&�{���{�z=����ڟO*�2`�����V�`�>.*�^�ߠ̦�����O��#�ډ�W_���1���Dz��c�S��{���ƠW�qg�~d�Ď�WyԄl[�P�t..&�޻��w�ܫ��h1���>J%nZ
Q���Sr�fi���'1y�md蛮a1����*X&vM{P�{o�K�y���p��T��Lj�h��p�E��z�u���8�ĺg��"�.�M���z&#IY(?����/�dH��*r  9���+��-��f��דX[�E`k$�váf7��-Y�U��{�K7�!��V0�FHAD��p�3Q*��a�s��kv���j�_�V�(��N��\ע��=;���Ɓ��}�ުb��Ũ)X����١6^�ע���׺��Һ�(����|�Y>�*G����{NzOC����A������n�>0����fjq�`G�����RCǘ�/�ʞ���O��hG�K�d�x�)u�*�~�Em�A�ʊ%�'�N�>���XV<�Y�,��1p[W��{֤z=^���u5�r:c�ă��˔w���L�R�^�W ��U&2���o��rׁ���22�d{b=�cq{&�}���ǝwu{���s%�2l�mP�U*���ǆK�9i�k�}���0���%�V"?�O�wnT�����B6#��~����9�����g�v������w�8{�̮��\VwF������ә��N��	�Z�}������ٹ�^ۭ���"��ߗ���,�P=�(�n
��M��y9�2��:����ey���\X���������5�j��v5q�B�m�B� qbĘ�']Ve4��W�y+��J�;�l]Y�D8�P9�38���(FQ�R��3��˭=�{te4q���9��ܨ��D95b=����/�2;~G��v�g�a���s���w�H�;Fw�U9���]����q<�� zDv@�q셝�F��~�O_�f�w���a�/z����ߗ��^��O]d�ӹ�|�=��p�iT|g�V�v
w������sٖ�����^}=~!:^9�üތyr8�s��������M��#/~O�`�Vd�@^�r��Q�q�1�s���>�0�N�WW�Ig������r���xǑ�*uc[j�]��(�A��66�����A�������\\�����G�u��}�{=&w�������!��x�@����9I�k䓕Mj�#���������j��5UO�UH�߼r⽟E��f�7��+�~aq����R8d;w,4+�:CᙚsI��zbr�)L�|YW�9��s�Ȭ�_�������2@��z������@�x�R��{7�k�uP��lKr��#����G ���66�H����"����ii���Wi_?�ɟ��D���^Sʖ�1֦���2z���B���0�U��~��(������3FP�v�F�SWm2��3z���ޣ�^�P�T1���"1��Ֆ�������JSDf͊����H�����qLqR��d͢�yJ��c,�H������J��}h���&Vt�w۴�/yg[ĵ�#�5]챚9 Ǉ�|���:�US ��P���f���v����)6.����st��<H:hI���,FCo�(g��z$�]���@)`;P�M{DWt�϶1\W��Y���[V���,�������KWy.L7�˜�޹��?W��������H����Ld��=7���x����w�^b=�~��+�yw�g��|{7=)�x�ީbϼsf��
�8ƾ��nnti��pw�]��+��@눑���w\xVߐ0.��!�3سӿ;���WC���ա��}5���;QH�W����n�������P��=B&�O�adp3o�_vVB�����uA��^E_u׺�li�y�H��6���:��]Y�����w��w>tVx81�jn&j�s5���)��G�#<�xzF�/�^,�uޡ�n�f�
s�"�s�^�G����Uryy�+����+�U�Q����k�_��������Z�D.ʤ``��T�}��=}[w����'x�@�{9�W��[���ra��t���xwz�_(��s�6�����"�ȥ�ov(뀯���^�1L��]�)ڬ�׼2)�U0�bޫ��k��T炒g��jޛ�E���яW*zϵ������l���v�n�[�e����P�Q�F��y�0
��d��u'b�",ЈU���"���L�����ܪ�����;��G��p`q���U������_�r+"��p��:;޹�C���C�7`VF�z*��3^y��O������!T��U�A�@n�# �l6j�_[�Ȭ���Hy�=y�Y��q��g��.���z��1N>uRQ2����ё�E?=�1E��(��j���>gQ����G�N?��m���!����~6�U4!��6$J򫜿K��
3"��v���9�>lo��/����ɬ����,��q�5����U�A��3������[���?Y��nRf�a+���T�s���e�6��{g���y4��R1��f�[�=�=q���H���H��;n/�&���S`���dd5��N����|��3�ȇ���l��\���4N_i֢����>�;u"�^\H��:�VA�a#bSC�t^#"f�4�vF�0yW��n�߈����zd�֜��yu=+*��NG��6�����y{��WM�Dq��w��R� �w�|�Oe�o�}�][!�{�k��G�dQϿ^����V��<:�>�������yw�:Y{�����v�)�v�!�ص��4)W)��d��|\�Y�~\�u��:K~�5���z+Թ�UJFd�=k6�k���l�ڮ�2:�Q��^�wCr�[�,�r��nD`V��Y`<���e�M(Fd�C�v�J�N�ԙ�G��@�h���`��p�����~�mL�gylzu��zG��Ë��k��ۮ0;��P��3U��3�켇2��E'^����y�4�g�6�2�W�xT����7�e����RH״f���
�FE8d�mI��&}�%Z���tHu�8�,g�=s-�I�d���	��\�����ڟOwI�콿vǙ�|�{g^UI�Q qC�_�)\<�9W�V��1��d=�=~����''�J�QQ����Ą��3������:eD�aW� @s9>W�6=)������&����^-�ۼ�1�U,27�R����fE��D�����L�\@�3_J��Y��s9��C=�u:�]nu.���U��G����DW��zu>�4:�x�{ vz�y�Q3)O�K�������Qk�/��ʝ	 q5���}jL���x�}��<�~�@��{ pȏ_�*�b�
���ϙ��qtR>�}�JՌ9My���ړ8��9؁�Z���?y���_@~h��4�:m��؂y�W?���P[��>�n��ٴ���a����޵#��
��c������c���,#�گ��wxy[t~v�5���Y���:P�ɛ�,���T	��v[��i�]���\{l��$�6�J��-��ss����f�N`�bJ��&^�E3-f�'o;����5Y�-:TQ��c��6�J����jL7�]�S�꛳@�3�*��[7L�M��ca*dc^�q����s��yUayf�iԚ�5G�c��P2=�\���=̛�=�B�C
�m99>���r�t�Y�}��2��Dꮏ5i+ʌ�����{�dC�E;�7sG#׶.#��Z3�F�j6�_��A��=����{��C���������4�l�u;��؆}k��U�r�ٹ����F}��ݜH�2�c�����'љ���xV� �-Y�ڎ9���|�Ӱ���º�x=�F�v��,@�M��0*;���b����}R������+�+��~����]��_<��P��o���u�k��=�p��k��`�γ����n4���������o�ݎ�S��}S-B����+�#ɕ?D楹�hi����d�'Mm��@U)� e������S�z�4�2&^s�{�9>���H��\�>����y;��@�-� �3��/`�����!�h^��[�DdC�^M�~�I�>�[���\�s�����D�� ��]-���~]�E�u,ۭ��J���.V�S������*[�ߊ~n�G��V�KZ�4t+�6��Q>:���&�v^���/�w���;W@ŵ�Q�&�%�q�˳>�����(�5"��3���]c.Q��Wy aCڕE/�VW9pb�?O��=V.��EJ�(�RKU�dϤ{��s�Mz�ˊ�E��f�>���:���A����#A�۸{��Mk�c¼p�((�GS{�&'�����d�z����s�Ȭ��j�����~��yC΀d�W.���G�]��UlוPT�e�>LSvddA��t1pP�������6M{����7��n��2��rp���6L�����*Sʀ[BC�)����2y
~��\g>�dzc#'��iq=�pz3Ѥ�� <�վ��fk�V�T�k�T/B���G��{�!��}981;�7�={M�~F�z��G��,F6���{���Y3�k�(,ӵ�ʁ�zk�gQ^��{��z�-2mW�[�~���K�߳.q��}u��颫&��UHP�g{�'���#�z]G�MwyV��l,�!��g��A����U�C>��9�D6\y\?M��|V��u�;�|{n�s�W�둲���+/�!t�ö��}��}U��j������j�oGX�=U�yq]�}=մ7 ��b�Ԭ/�P7U����5adp:>͇T�f/ߒ�s�L��#�$�f��+J��s�9V��Hb�z�y�ٛ��Z\���^�6�2b�E�y���襱�9��.#�IW�%��PW���ۉ�[N��\�1�%�x�Ɛ�&Ry%�Ź3e�)bq�H��[�d�\�'�a~W�u��_~���$�p_h��t�/P��T�o�2�_��wz�UG����������k��O��
v�=#}���<Y�B/N�p�����Nuۙ��7���c�o�B�,�63خ|�'ג�8z�"r5ǯ������j|w�XD#�H]DR�ȹT�3z}���������jp�۷K2��x�&��t�z+���g>~�> �M�G�q_/A������zPȇ`y[�ώ[���ExW�n(7~�|�ޙW1��ڣ0V�>+x(�L����Od;�/"F ���*��w�Sa�7�P��qN�w�]�o���8D��Ǿ��G{�<Do��{#�lU�:�(�Aw��TݙE?<�dȫ�(ߒ��\�j7�[�{�؏6�c�x~�@�]�T۪V�n	�ŝk,dK1��7t[�=��n�|q�@��z}��'!5��3�+�Xc���L�&��ͺC�7�C�|9j�wж���X�ܦ�ZUsYR�!���I[���̜W?��l���1��Ɍl��1�cmc6��ll��1�cm��c`���X��������o�c6��l��1�cm�1�cmc6�61�cm�������c6��l��1�cm�������6�M��o�����)���.y���9,�������_���1%� ��K�IQBD�T
*AE$BIH%U%$*EUUT�@$��  �P��@E*�IJAJ��$*��1���%D���%*�(�!)$
�%�%T��B�i!U*�$UT�TH�E��!IQ"��f[�ʥ@��NYR��JZ�J�)"� *�J*��Q*�D�
�UHJ6�I%RBH�*��A@�(R�UJ�y��R�b�  �rB��уV���P��!��M�%J����b�hk 	���-�P(��)�M5iYZ ����d�T$8   lࢁSK4
�V�(�XMu\Wn(���QEݶ�QF�X�EP 
P�����QE^�\tQEP��V:(��(��.�
�EH�R�)��  �q@��]YZ� f,$
�k[ Hjj ���TZ )M��k +`���%k����R���Z2�D���  Y�
{V4 ڎ��
��]���݆����PU;T�4 l]à(�� �
�b-ѧ@ 0ª�%$�*����	�  ����MY.�C�mTij{�e�
�j=p�@R��q�,ʦ�d�uJ������� �Ɂ� Rm���cJD��%B�`�%U�  ���m�`m�Z�6k[ ��4�d%j�@R���$խ�D�h��Yehh6���`���@�1�j��#J��D�"����  6sM��kB(P�F���BҬ�jd�V�m�A�md��h6afڱ���V��5�Ph-� ʂ���Q
 ����  w\��
4Ͷ�*ڒ4�X��T�$-�Z�(��&�@j��YB�V�5Vh[m�R�T��6���b���M��Ti�JBHJI�)�
!� ;�Af
�0�*�Fh`�J�Q��b�lm����I ��P��b��(K*%i�`V�ڴ�Ű�(�J����(��*8  ]��h�U�iZѱL��,RL��4TCCB�����m`mJm�ڀPՅ�F�*�� ��l�*��I@�@P   <�ʒU(       ��a%)Q4�24�4C4�1�	���dɓ#	�i�F& �)� �$���4 i�4h (�S)���OBmBOҟ��H􇩦�)��A&���EOP����F�	�vu��>u�kΝ׽�iϝ'αX�,֙"�q�5l�
W6��[N"��/�t���,��A$<@D^A���S� P�%X>dLEl�x���A�_���������0�'�	��@@��T VHpJ|�� �d
]P�@��Qs
yx{����:L�A�y�yWϔ��DDDDD����$�PB��!PB��B� J��) HT�	*$+$�
��
��HBQ&Y�Qb fU&f f E�@FaTVaP �! �	+ �+ TP��P$!Y$T�� �I�IT��*B@�A��P@&DH�B�QUUQUUQUUUUUV߿g�D���S��w������%�T��#G����H=ў��@�P������$,~�������1u>[K\�yt�����֘�w�r�k��7�**1x��-6��N�,��̫������VQ�R5�� t��n���k*J��m�;�X����4����	B�P�x["o)7*�)y[�ݴ�Q�V�m`ت�a���X�l�M��E��e�&}i-)����d�L�k1��d��x.l��,�!�<2�7z-�`G�	g�G/
u�ՠ7�0�c�A*IV#�:��"D��w��1 h0c����f���NQ�y>�wr8T��H++JH�1<��j��av�T�X�"�7��ZS*�2� Z��utՌ�V@3\�;˲��i8M�)�m˹��R�&L��y��	�.�լ5NZ�ܣI�rYN��$e?�v�*�fnZ;`�d�I���e� (�C�d�.�J�n�ءWX܁�P�h;�P�VG����ӛt�bR�h��J'{g(���߰Lh�V2�T���H]���	ī6YJ�xe^�:���Q:6gbW�Z�F�Q�-�+�*F�:Ч��u�R�	ddIJ�&��a�J�H�o[@h���+T9Sx����Xp�V/e�*����-��ڄЀ�f��,ݺ .�5��݋2�
�(eG���k4e� ,����eֺ�j×c2��W��m
'.+a�6��VT�+���re	V��l"���[b�n�Z�&����f]�'��,/f�V�{Ge๱&ʡ�^���J,�'��r����u&�-+r�v�h�r�J�ˬ�--���ܒ�&��*�z�����e��J#oJX%7�kpY�~C�DT��b��X@�0`��CP�Ȟf
���V�#��UZM`�q�ߴ]6GfI@3A�u���FRz�|F�u+�Ch�	�ģ[��zH�GM�bP���"6�����wMB��ݔ��Ϲ�!���رH��.4����zs^!�3F��5X��Lݪ'b�V��̌m�	6�M3�G�v��ʧ����XEȉ�m�u�:K�-�F'�ʆ�Yyt���3j��[��/`͕��^��GbV�+Ѐ����1fYNĂ����8�wH�����U�jɂ���Įš#tr�^�f(�q�225���`͈���e:�)LG �yN��#N�nY��n9�2��K�/U�����y"�Hl�������v�n��1ѱL�Q���-�:�@�ނ��-\LD�on ���l��J��*����"l�h/�4��:U�M�P���ܺ�rf�kB)V<��k.T T[X4[�U+hb���^$����*h�o#��۩Sh*4����F31`4�,�QA��-�K�o��:���nGJ�2G�u���Rh36�� �ʠh�fZ����@`|�;����[t�k�MiV�M͊+�DܻTh4�I6-U�x�(k&^ˀ��
�&�2� I�U
+1��-J���' +Fm���uq`�r�U����!7i,�XI�X9Wu� �4lS�[r�,4�j�h��;l8�}�4�f��H�!{�K���ˠ��F����+$V�Q},�l|Ԭ�v��kJ��AGY�l�R�Z��5+��3�lQ*e�k��pӵ��Pܧ�̫�҃c��J�ЋTW��E� L�2R�R�c�MA�����bbcMm��֚����:-*��1�H�
m��M%�V�TW��^<E��L�.ܳ*tn�����	�h�j%z!\S�w���fnB-�lj^"�"�j����WBC�E�[�57V��5�ە3A��l5v�h�����������j�BӲ-	��߱�ѡii�J����38�K�m� $v婑�	�gC�h+R��'�?2O�ȅ��)�$u�К��vd��&�2u�g3���Db�n�Mn C��9��,|�%���L����敎�G��bc��Y,���Y1�	�!��"��\4әw��V��t�
ˤ�Y���6���]�.^I@1K*ebВʋ�~n�sO�d���NhU`���Dc�����dTV:�t��]MKD��*�!�b�9 ��6v�T���<�nL�F�����:[��rAR7�kt5m2�u\L�r�YtV]ͧ,� �R��v��3��3]��28��Ř�%Nc*�ɃU��*�Hf��n�#E2�Rr���{�m<SYyK
���ֵx�;JK����GzF��`�3�*&T��E��5Tj]7YY�-�$`v�ye�u�n�D��wiZ{����ad�T�1b�VM Yb�$��Bl:�6"Jp����Zicx�KeZ�J���x��n M���T�S��GM3yt�0f�Z�)&l �V�Em���)�l���w��v�*5�3�t�6M������?�Y)Q;(�K�$q��@i�u�,*X0����ń��1.�$��X��v[X���S
�%E����,N65ݙT�J�ZT��Sձ�(�×KUK��o2�tv2o�%�^��ɋR\wf��ֵ̺���W]�ٮ���8��G������kʔ�Rb��a3�5�[w5ӗ�IQ㡆+"��P1��i˭��h�mr�*���F`�켨k2�@��	�R0,���LM�%i�j�pU���l��7v���J��l`�g^�I�J1��@�[[�7W�Vc1�NY.� Z���Ʌm�,��h�V���B��Ci
�z��5���w��%C�H�U�[ȜY��(�����ZuH2��EB�6$R�E�,��Q��k5�h��6�@�3WYX7ij0f�]��f�\��]e�:�=�b�Ӽ�Z�1����*ܦ�� -x�V)��p��?e6��⠶7Z� R��
�Ø��jԔ�8X�:_�t�`��-�t�;�f�d�[�0R��)�S�X���y)�4�P�.-��7�d5����X���û�2tc6�͖Z*�F�e�CmV��vҙ{,^�M�b�;�iT�5�`f��U�t�ta�c�Zst�Q�I���	<�ff�n�pFqf�
S�-Qmj���hҕ�$p��AIx��.Q3&�p-2���/&�
���5齁T�\ 鹵�51=���9Dcڸ�Tݫe���;�F*���{���@�ٸ�
��6�j
�f)��A+[{u�Y +�(!k+w��Լ��e,��ַ.�c��G&-P'�)�� ���FÔf�ɖ��U��&C�)��SY���i�	�Q]؛��H\������-��$Ͷu��,��Q�73wv��WB	����!Nh�2�QP���Z���b�lZ)ŲAW��%C�{����5o�oHʹ3V���m�p�
N���f�$F�ЩF&�^fTFG��Ŭm �d��QuK:�&f55V�PH���j�бR�F��^YkD>�uo�G�}�2�$
�)+ox+�@���0/A�>p@+�f`���M�Ba�I��dn$�F�~S2�6fS�a���ƥm-u2*gdpK���%�u��tcn��@�+~u�� f�!=���3wǮ�8�Du����-V��V�c]Z�G#	�a\N��Ǜ��m�{o^n�Q�wo
�D 3ItVfT+�d��Q�H��X�T�Q��{�+��Z�>WW.�"nnkxpa����������6�%�a�A7<�f�Tki:ަsK����;����YPISw�T6L V��\rYH�V����¾EK��h M�ދa�/V���ڙ+"��Y�Q��7�w*Up���JWX0T���&Ѩ���D��ŚCmh�ܣ"zE͠�CX���n��4�Q�hSJ��^��J�I� ��*F�S�ё��]^v��+5XA�N�e�⌺S*�72*\�P����ן��`e�u�5ZR&n�u���*tq����`�V���vf�N��YmenJ8��1�h�b�Yj�d\�b(ՌZ�F^�6�kM
�Nm+*e�t���+
E���I��&$x��ԓj���h�'eX�ӧJ��
���Q��\Z�m#zJX�;*�ӨH�'�f�{��\q=�$��U�A�
h���n��ܦΚxl��r95��<��"^ݭ��Q�mM�ADh�J��*�*�g3/6^��	a�Z����4�yb��4ͦm��4���K���4�S9M�َ`Wy r`�o.��r��ZL�&��(�˂�1�ff�kO�iJy�E`�W��{�4fӳ��ԷX�N�6�w��O�TˎĦ���SU���7x��n�I�FL9J�Յ��$��;�k1�&[yLK@�k�t��SU5ս�Tt���`�Z�)P[�
��+lL�YJ]	�j}4�mӷ���,�ө6V�*�1jJj�cIJ,�@hAcI�J5��L*��b������MϞ�٫�[A֡b�jlSxH<lS�[�^PG�ӔK����;n�L����ܒ�C��#B��c�q-�R��*�P�F��K�	!�T���\�{d�.`�V��
�#vV(��ŗm���/6�̩6Nࣘ�P�حA[tU��3�7D�#Im����A��
��w*�rն�^�t���Fl�=ۥF��u&���K�?	��0%諰�XV+1��M$��I+Cf�(�wUM,`�Û�m�`����V5*��k[{��H���B�R��b���f�Kj�IO(V�����yw)�Z֯��������O-mf
a��+5�f�ЍևL3� T��~-LN��z��݊��7.��PT��f�A�1] ���Xӕ��y�p�X��j)oEnP���Ӧ��eU���#:�"kٴ�U*X@EM4���ׅ԰Ke���E,���
�v-'ؘK%�c�P�O�Q��.[��EN�e�Aޏ����1e��wa
�ѕZ�ZM��8� �J�$#to�	hD��f�:f��*D���x(Vs# .�X5�W�q��*��ppV�zy�X�r�u��ތWkK���EP՗XQ��1�sG�+]ՠ�n:����~Y�J�Dc��b�i/��m ,���R�L������� �n�.H��,���1T�Q�+[�%��i��LME�D%���kV7a��J/j��31�T���R���J�WM�z�B�i,L�A��R�`�yZs~,Ӧ7s��ůb�Yv�+T�"�[TN��U�1u��i�F0uմ�c���2LY��B���vh�mAx%*�P5Wf� c��V�Yb����Q��j��Ø�ݐw)]�U��x-ɐ��ƞƥ�"�,�i8uE�=����0����+�!4�-��3@���r�ɶ�ء��V�k�1����+ N���82���b�k-Y�I^
�$ŕ�C�nVͻ����@�R'�a�g@�4�2f"�[i�k]�1�[���VXX�Sr҂���ԮGR�0��r52�jl hT�0n�B��JY���B+J銽;�b �T <L�wV����a�Ce��)��D���r�L�S(㳻L��d�c��w?;��Z�"Ph��:�!�[��׈��a�(�cX	�k]{u�bCE��bZ�@0�)���#z0��Б�v�nܧ��W:�m�.�)�P,<��.3ތ.U̖���Q��j�M֩n˧��YUV�a-b��R�JVU0�Øoiv���P>tҶ�en�
�dv����x����M���)�\b��{b� K�،��H�l��R�	�׿@ėÔnCF��/�*.�*�N��q�Ƴm@�e%�u�@n��'k���hL$ZUL�������^�oh/��t�C*[Ne��;1�0َ̑�jU��b;�X�hܰ1�bX�̢~ �ݽ�j��`��$�������4��!T//w��Y+:�U�ܧB���sA��7c��5�v����YrV�����U�K@!d�a�
�]�T"�����.���aš�őB0���b�� ���d"����d�N�в�k&���fh5NVd�c,��Hd���
��q"�U��	I1E����,GAl �����Gn��m�"��PY�T�d��}�	�"ڎͩ��{o1��K�D�QI��'�Ҭ :�pJ^�g�3.R�75Pَ��-d�Y��l@�)X�l��G�T*m���,K�VnlV�;�o]M��T7�-�3�n]f�Л�\gArl��-3�J9��n@��X��%�%Sj��)0˘n�	�oU^ �t��
���F=Ǧ}���+�pH�V,�U�7h�F��0�(P�Wrc���-*��v:�ʴ*J��ݳxkd5�B)J`��ui+�ۭ��nb��Z�+6�2V��F�Ys(��D��
ND���+/v��Y5]�=j�7�����n��#h�U�+Z��e�J�-43f��E�����
�vIr[�.NL��聳l�%�t����JӬ֯)(W��.�I�`���͸�Vx�C7j0ͭrA��7t�X4�(�
�]bl;��o�dS/E���4��J9�X�u�#��!7Z��hе��5���YPD�& U/V#3~i`���Ak��4������H"� �5q�r�ᚯ)��5;5.ej��H>U��ڤ)X��WG�.*Qm��դ�]�j��!,���VF�<yk$N�L6Vb0R�96�`�:��
�M)j6�(i"_�Р�B�De#T�F��)9���'�kR�XO���2��Wh�6xU�Ip�tuT�F� ��d�S��ib�ur�K0noJҙֳ�LZ��0�s#.�C}]�����织:�!H���]�f�v�����m��5�`l�2�B���{Q�k>\;-��9ۺ�u�N����9wSW��o�y���]�2�\�ۺ��Q͋����y�J�OR��M�}tD'=�+`:<`˘7��A���e^��S���U��:�s�������4���s
�w����*�ﲎ��s��9��X���d�ť��"���s9f��]��x��f%�T����ڝb�,d�zgwB݄���t\����"y��);�f�r�{��|�!(�\{8f]l�-Z�.-[ �U�kJ=�M��|hq.��t.�VaX.tW�c���a.�	��d�X]��sg]oo�W9��)6}"��e]a�ε��f^�|���
�&�U����0��Rޫ5�m�	��b,�S�-�����&d��a�������Y9�6R��Խ�կ���v*��v��-ا�|�g.U�%��%�)mo8�����F�㗡��/�T�D͇�d����x�=] ��f�V3]�2J[\�,�'Iȁ����49h�i�ϺE.�'w݆���r�ߜ$�,�meujԏ3Yi���({���j�hs^��y��WQ�́��*�ժѱQK���N0֋�WK�$�T�ƴtS*�w!����39r:B�I
�}�(J��eY=pϤ�]W�{��V6k7���Gs��\a؛*nc��l�t�TQ��m]併���X�c2�Wt	�xps���
'�)T�V�˸��¶ͻ���7D���U5D��02b��Y�S	fH�ܐu׈ݲ��(��H��u���'|Ɨ��SXs���%��f�٫��K�CM�̬	���L
�~���mv��@ ���s��=��rK�ŷ�alؾ�7��30� �1�	��*:X3s)P�{���x8]�A��D�E��+so��Dk�K���4y�1�R���9���e���h�7�мV��5��7	�ʬW�U�Ԭs�_*��<j�oq2!�J��}�̑�2�r}ז�$��Z������j�WA�0��;u�ҕ`ڼ*^�,�W�|��x���H����]�ɇ],���/3�Z/��h'È�C2�X�57I��[՛]�����d0�VXx��q��=�6�%�c�����G���8�\+�A@m�����_U��Y��*Q�i�4o!��d�k�2�p��uv��¸�"�9����OW�=d}�ʻ��3��*;���V�N:����K���]:}-�אm�t`�ͼQ�L�,�z��I�v[�RC�l��t��2����	ܫ>Ok��Ч�L�)T�сH����$�k�pr����U;�a/loZ���Wp9�#F�`f�X Z��T�WW����J���j�L@�4M�V�*�ͽۗ�M��-��|�ȷhv$����`^�Ge��PKh(��.��n�B��N�Ŝil��b��r��r�R࿘�&<3��0�1�J�u-��'r`�nSp��F���!u���v;�Z$���R��t�)wʱ��'�����6��7N)n���O�u��n��Wm9BG
�ϳ�-=���L�����]L�HԳ%���e�
#���orpJ��.�C {]�0�&pK۾�+u,�2��v#�̭ � f;��v��qOn�8��Ÿ�l&/�D�u6%e��j<�R��2�E�]��9�������Y�G�:H-[��<�����={�	�qj��/Z������na�l�����;����2�Wd(ֈ��4'u�L���1;gm0Q;�ֳ�@�-��Ee���>]7,�S8q�grZ�K�bF�Q��i�5Y�>\�6��d{+�GV#�����]W����(��B�T̗&Ag�B���Y��\�t:��3B�Up����Ot�0��u+���Ւ:G���yb�=H����*��Iu��Mv�����>5�A�9�̊�m�sOEs,�0ɻi��[�C/7����E���nc[�}u�[���B7b�� �w�딁�<],�*�Xn&�*����xh��A���帑t�q�0Γo�=S��E���'{ܕ��t���H�0�H��Jz��n��]s�B�k�4%e<�"�K�4A����i��[�/�����&	��EI��n�Lm��g�~.�E��;"�o�v�2
o��鲷��*X��G^��1�m�Y��w]�5��&��u�K�A����wu�ޥ]����+�1��T��h�n=+�7;����Gp
j:E"w;R��AhK8�7�2���GX˽��5�qq��F�\���'�
���X��r�@S�Ǖ�TC0'ԙS�$�pJ�5%����֤�wl�\��"���-e�'yͤ�s�����0�]r�ĵea)�@��<�1ML�vMu�U�g-n�3�K�g]v�0����'m���˧z�ڱ���F�b�۟tam��ECr�V=Ŋ�����u�)К6��htԴWf�G�Հq@K���d��m��c�5�Єe����Tޘ+����C��3uwĎ7�SM5ʋ}φ��.��}�P���{l�nlÆɩ�'q�,�+Q��	�������,�q��ɝne���}A�,��*�򤠭T#��7�G��j�Ζ8#n�e�g�5����F�VX���(��ӟ-ޗҊ�fo(wvP	��&����m]�(f��o����If��J���K��h��[�����Z�L��n�W�✧gh���^5�ٮ[��5��R�{C�T�`Χ�]q6i��k��j�%�a�uZ�o������.u��\�K�.�@�����tȯ���*t\�Xd�1�\�Uʮf��k�X�zk�A��Ϋ�.�f
�S�_Po�r}|X�I�X�
�݀ۆ�f�]Τv�v����*6�,��rb	��M@R�f]Ƨ)�{�m�⫋���ss���UϬ}&�#{�hν�D��{8��]��×#�=��]W]�u+�ܩ:��A�3���'C�e�+��̒]˨��T�M=8���{�<�6�/�� �w��M�)�����=��B���uX!0��E�O+^�omGqk��O5U��\�/m��tWԲe�#�ʓ�';9nN쨵;�W���M4�ˬJ��4�G�=I}D�͔�vK�vW�)C�;��{�uyr���]u���f`Ԗ���Գe���e+uϝ�R+'..�ve�֐ڲ�7��l���_,�)Qy}H�5+����W#d�� k=��/g 0V�z���AwEtRw��^X	���Nҥ�0�ޔ$ܮJ�q�e��v^T1���9UK����n������t�dܙ�n�]*խ�D�X�z�6]I��V7+Z��3&����({��J�N�F�M8�VܙO��۸!ر��卬U����R��,{���7�������!�鼆�Vrq�u
K
}b�ݘ�e�sLe;�n���-c��20�Č���Ε핂��)nr�\;��w�wGL�,z�;\�;&�\턨��yX���ե���B�'�l��=��lZ����vk_"T&���v_gG���˻�IU�:k#L��HfQP�2�����ܵ��c���+�c�	/�?��E�w��)o\<y
�����aӷ�A<�ޤ�&��]e��U��%u	�ۂe�hj�#��nL@6:!�rT�:K�tO�ά'N�#{m��`_V�����@`4H6���65)[��;6��-S�J��1�a-DfX8c'� ]���ڦwvA��m��p���%D.���tM��v� �L�gM�CB�J6�7���"�Ƨ:i��-��k{���|rV^�� b�֕�Romɡ����q��z��t&�ɔ�t�Q�/�ɾZ>�}Ǝ��V���k��ć�����d�"Z�ﻖʄ���t�j��I��{�m^��hc�����J�q9Y-I���m�9�\0,���)�K9�{��u��f�Ď�'�o!|e�U�������E㡢�L��1s�^�f�q�M3�u��3q�z�N�o&vJWC]��u�*9sYł�ޕko�Q}��Y�˴��K�3��I�Q��쐜���1�eb�O�%� A
].^*�ڙ�zѮ|8�kR7E��/�}%s�f��î�E1���{ɶ��Wr�̒�տ�u"�
6�\�B����Af�e̳�uP����cKt�39�ņ�drX(�ۚ����Jw��*=�N���TgS�u�� ;2�
j���X�Mr[�s�I�,�ܯP,a�.��	1�XB]>�;n�vRZ7�plڑQ˄չ�!�`�ñ6��]�4u �ԍ�[O@�+�P]v�K��a�tk��o9��NV ��^��k���]�Gi���m�V+3������Ww�U��C.����]i��N���3p��է��і��Ҭo��\��Z[��6���ֈ�m�EK]\��82޸h��tL�I����|'8���5����[��;���]cK�}��u�;>B��(�X%:aā�3Qt_Ö�����<�urJbw�i� ̍��V��:�[P���6���y�gC<�^W( T��>���`�1b !2�����a��v��;o:�b}���I�Bd����|�%�����ޘ����Yger+��۽�"��R���wWC�fX|�0�� 5�!���p�[�_!څ7���9�n��b��2X틒|L�9����{�ƊN�ZÒ�������ے�@v)N�����/�]m?�N��9�.ojan�N�h9�Ε�*�(qA�H�(��<�G'K�W4ia�}@T&����� �5���+-$ wG-�q��z��C`�(�GN�w��" -���5=/5%փ��S~�#�Hӽ6���J�>ᷴF����Y��7qt�ƴ����G��u�ū�/gw�5wu���.c��yK�weʁ��& �lk�%�����tt!�v�ա��JR��N	i�"�e�:��O��`[kN����i_����.�]���vɏ��D㥃s�u�\�8�of��o��r¢8KI����Ko.��k���u�YA)A*'��o�X�&��l=(��b�62j/0Ȇ\��]���w�2��_s��Z�9��튪�Y�@�%$�or �j�S�yZ�+�4��5��z.����ټTK�H�^oZ�7�T����ʌQX�����a� BNvf\��\�j��]��t�eh�wHV
=����� -�]�V��7I9uo:��UL�_��t�*7p��{����c����ٹ4��V�6��˚ i/��T֮��B�3]��P=��݊����`I/r��ͥ�Dr����N���L�V�=W>%�����U�D�N�7[��՘�	M��i��Ӭ�d�H�1gI�ZGR��U�E�z��/��e+x����Ϋɵ�oZZgt�+'�u ��H��Dz��Lq8ǋ�U����{�ee[�8��b�9�69w}%�|.u�:r5��Nn���Ƅ4ӎ�'��w����<�Q��낢�8L����{R�]'���wQ���t��\+�;��	C��Ĝ`G�u���� dp��guY�Q>����K/�[��&u`�+��;�����Y�X�;,]N�pX՚m��p����+GC�y\��Z�f�D�	�tCTdf��2�N-��Z�+�,V)a���u|�i��qRl\%B���5�W�l�%Q�X�u[o3OJ��jF��ď���*g-�������*���0�W��_A9�Zī���G@�}�K!�0p���ը����zh��8.�(��1Y��m]����Gn�3��:D�b�n:�SY�̝�XD������"��Y�����{SƴWV��:):];.wi�l]l�gD�q�$K���O�Z�$j��Ն1qkrJ�+
��)��:�U7QfS�FGK�WN\S9�̕�d,�A� �)�uA���l�2IܟR���p0�׸+���R��T6���ŷ�_Pz
���M�܅=(�����/�]�:w6�M� ����A��g��v(�� ���3�u�X1�1%,�� �)Z�$NWR�`����O2�m�@Wrts�1�u��ɽM�K:�=z�Cm������Ȇ��A�9r����ߘh�oX,�}�B�nL���'mm.Ck�ǯ��u'ϪC�����:���}]Fqs	��cWC��=�:�hÎL�e�M�Ή����k2�K��x�@�f�(K����N<C��V���B@�2f'ى=9���!IZ����C��кK�B�ٹ�E��w^r��+]ir0���L�<����cnM�Ո�y�3�^u�>Q�/�s$��s�geL����y��I.I$�\�.Ԗ�и;(�ܖmi��^�X��>�μ
�;��sW��Bp�!�n�Z����`�/R��=�^̛��|[>Fs�M�a�C�$�7s��"``KsBގطQ�=�I�j*�\a�;L��ZV��H�Xk�M�8[��gZ�5�3RŎ�dJ�q�	�E��Ǡ���+���y��p\k��u�ΞNj��)]���7���gۜ�X��)a���%.;8�M�֪�T���,�Îr�֒�YJ@R���]fmt�+�z��3OW(��)���f���y��o�����em\雺����2�L�ݪN�f_ Y��:ю]�����Ki�,���pvY��r*9b�8J���[�(K�U��b���@ᶠ7�:�0�=�tySFH�H�3���q���빨ɽ:zw/ǉ����(*-M�+�m~w�@E]���E�
��p�y��|č���T^'������]�M��k3�����+f�w��`��VЉ�Ǯ�ћ��5Ɯ�ޣ3'0/4Fo(q�Pu(�[+'Kc����q�P���f:x�!�GKl��]�	46�	w�ld�fn(�n�?fv�̾��í�/1^N;�-Hڹ,!1c�Y/�D�8H�W�>���HJ�Q�f���#��+w����
��&�����t����0o9��slW	�>8F�����-R�ݰ��vhLX��}b�������7;G+|�9Ԃ9����z�ݘ�w]N�oF��A�j�Z��6;�'ʒ�9.��8a���)"��_=D�uԕ�t��N��!���Ϯ�s��fI81�X�Y�0#E($����*�9�/E`����T�4�hp[�	yR���pK��f������P������(;�M@F�W����YH���v�ݢ��K��&��ƅ��I�eT5�{�}F�U����Hjj{ٕ��n8�(Q�٥]G~�@���9�;�8�qk;�Z汐vW�v���Eb*�<8.�O02a�7w�A۝��b]ж~+���[l�\�uܤ�V�,=��d�X-Tnu��z�N�����*֭:�6�V�c�h@�k��¢zg\YG�1-�ٴ:,f�#C�VC|{,��IC���ں�B�tT��J���8�{���sdWF<�$���V�)(I-P�$����KJRI,IX���ӹ�r^�eeC�y�`j'�nT��eۯ���kb�C��ih�z��1���&�@a�-%��G�!�Xv�ӝ��h�#��ޒ��>�m�H����h�/�a���'-L,�3��V�.J�g2s�3v�З[�zy)�v:�Hs��2������Qo�1 �6J[a-�h�+f��e�<G0:vT��w.-J�����=��͛�:��Oa_GQ�O�%C�Ve���ޠ�+!�X�d�o{q��j����Kc�3䒻��;�&�v/��p�RJ���8��ӣ�Գ�]��8��<�fF�$^�bɓzr�q����}Z>�ݹ�	���V��X��QY�P�fTw�k��n�а;��� t���J��(��b����պ�̥�f�%�j�1�u���ƚܒ`�k��>����[������A,�f��m.w*���]��i[�x�@)ځU��r-j�4D�Q�Y&*���SlI|eK�ɕ�2k+��j�j�M�*7{Vڕ��J{S�Va����·��gk�5�Pl��q�t*��e���א11,�t�ʌ��m�*t(j�����t�Ɗ�]��;�\ˊ�GNV�̻R<�q���G*Y������S����*̙��M��+HW&�i6:����o��3]{>�G���f�YB�*�
=�5*wwwwN��IbJRJfeBI$��I$� ��_�٤b���m�u���y��ĝMp�3Z��V̧tr��î�z�zӡ����]�W:��@:9dF�
��˥�A�י�\2N/�0TTE^�v'r<]�_H;)�ڔ>�\.�k�72�rf�םY͊�L�����ZG65Fq0����H:��x�ˡ�C4��C�J*B�v�.��Lӱo8���H�/$oFΕ�1�=M�Z��ka����ڻ��N��)��e�-̔�.�wv�]����b��(ݽ�fU��R��;m͓l�垬�b��	�Y����Pɔn�J�N��H-�:@�֐��6���ư����U��2�$F=��F��V�m��v�K�nlU�-�]�Y+��U�xp`�Wt�(%��/�ST4���Y�|RZ��]d�������5�\`�9$��3���5����3���8͎�;�Ru�]��y�:���Px�d���N+3U�'L'�H	�b�J[��].I6��iL�v��փ���Uྋ0u�O��=7]���[u,Ŵ^��(�7*L%��԰va�Q��bBk�(�Wv,���'J�ᲶR���s�P���<̋��C����F�R}G*Ҭ�P�Ja���Zˀ�o�ʺ�k=ψ셪C1H�B"���I`�w\e�hˠ�����A�X��m³�֩�[a�m	}O��I�e�ū���Mk2�������O�M�\��P����"�u4jJ�+w�s�&U�n�&}���	��Y���=��Ն�X�E���A(�'r���_]N�������/F76�aq�]DU�)�[](��*�+��L�\���`�����f�r�%Z�ō�>��m���&�i+Fl���(�{ �2:_�k���ې��'`
�;�GLh�83�L��g��䑗��d�ʐ������/6�_!�oujX��t�(�k>�\�)�#����*E�7�d���(D'+�uo��7��HpS)!Y%��Vk#ڷ��Q��o�޺�6��[�j�4�u���� ��]�ޭ.���OmA�{�it(t�B�t��d�7�μ�,�j�cc[�q��%�g˨r��<����ɂ��=}�Gͮ/t�T��ԑ6>��T�����"�X_�μUi�⽃��nh���GټB��ı$�-�o��g2��������jqf��+ed�}��J5����+�^T��|�+!	+%mliM�-2�^�%X�ܧv=tqh�m����BTڗ�i�`t�,�ܰ���7��n�P˻��(�Ӻ�[��P}��3�����K��:V3s�\I�3���&�.��N�*#&�YV`C��Y��9�U��֧$Ki��m�n�Y�]!E������&r+���s�ʬ�7�
��i/�V:s&���N]n8��Y�K��s�wU�;0)���p\!���*�`n<7g
��)s�3�К��+�w�ǀ��>��C	B�S�I=.GҌ�\aå�{У��]`�\���7��`[���.�!�w�MF�^,'�4�xH�&B7�B��HhgL��x�M�{��
�-�g�k4K\���_u���m�ݘ�45Nz���G�iK�@eon�S���_b0d���;)����\A�k�T��yb�\	t7^�V:�sZ��s��j@�K�Wu�W-�lD]MN��Z�ަ��O]�)�9�W�jx㣙JY����8�M��	�����*�L���{ɭ��2Q�n<��u09̓l�f�E�C��X��Ӷ��2̷7��O�뻝���7MfK���&Ixn�e1�$��Gf��[��n�D��O��c��@�����СKWp�/A!=�[x�
u�f��hVT�/��n���.[kO�mc%*y׈t�z
�ہ�sj��M��^���o<���yR(����$�-��`��AX���,4Á]|��f�>˺���K�P���]��gj��6�v�C:	�+.�vRWv������ݟ1���r
�oV��&�v�-�#�G�Sb�ј�KU�X!�YO�(i�y��֮d��k�tN-��^��n�>4���yET�|�k5�%��G`�M��[��Z)���L�:7�lZ��l�S�
�2�.
��f���ɛ��R�[8�w|�K.^r�&l����R�M�\����yYD�Y�"#EK�=%�^	.=�Ү<�63�@�nU��#v��#*��bs�����p���R��r:n����m���V��u,\�Ѽ��.��盼��o.��l5�'m$#�A.���O^��6%�[W�DIHGz!Z �0ݬ�	�Ү�jee��]�j���:����\p0�Vm˭	�i����AG:��u��{p�H���x�!��.z��Gb���G�Mge
�Ȁ4�W��Z��Z�7�q��=71Z�,��v��Ҕ�F�h멀ݮHU�[h�+J��#B������� |~nt�В�L�_$s�k�ԏ]��	��w(�{���;�"�5���
�A�S�V�+`'%N
�K�)��g:��7(��U��-�t%k���WYFb��'����;\�Y�;\nmJ�il���v�0�Y��n�=��TF�֤HHq�3�_1���jҘuݥ����M�A2�c�O9� ��[+l�o2D�������{[]dPc�M���V�w]P%��x�Y��F���Jhb�}���0tVݴ��zHt)�.�u���r�t�`��*�{x/�8O�X����`p�r��_;]XNuʴ�e�J�M,P�,I���֠s$g:�Ո��e����*����f�j:)\���#[�;/��m�	ܭ�س7u�d:q����ŋԲ�[�i�j�s��=[��4�Քg��qc�S���e4���/��No=��z6
�V�Ҋ� �>�J:�;�wpި�]vԶ��w �/����԰���Ǵ�
��ӯwq`JdR����e�������c�RNO7[��  HbU�A�u3]j�>Z�]M/x�kf��<��P�{B�Z�<EYH��
eQ��D�X8�gR�Y�+��[��\�R�Bm�u����8	f�i���4��lB��y��)Yy�wp�E��j:њ���"�h�������*�:��|���Ś
��p�q�J�Moe�[v��3f�Wiʒ�Z�ܻ�pqX�u��E����V�M���/v�r�p��vW�z�>��OU� q�]Jo<<�f��.�C#�5�#�+2A/��G�]1K��!m.s'/ZOUL�ͪA�J��u���O��}nV0�����T�	����V�&�
6ɺ織�+���q	��9S'`'��;w�k���PǙ:��O\
����ï����y�Xf[���3)����A8�q��bX��3;�*�U�-ƙ�^Z���]�ka=re����D����K���ܕ�;ڽ�|VLܨ��o�z���x�\��@���7�:�9���XC��xt�%�o����V>͹w��%�=@kW\:�!V����f��Y�ez7���̗N,�|��j�	��.�-�b����}r��-�ĨC2V��:��]�i\��_
�Y�O���ܧYn}z��� ����-���.����0k34�4f���p�7b�N@n������Y��c��Z�kz�J�6<{0D�����k-Y(msW����8.�V,�1�P�R�_
|��I[s(m�G]�i�<�8�u�R��"���R��ͬ��Y������3�:�Ɔ۷�&�*�:���R�޽��t�#��{�����s~�*�,��:��v!2`r��zl;���t;e�Ӥ�T�	n�B%�u���`��Su^��fӜNV�J�'j�jO� �[��K�X�h�YV6�X��U8jj��\Z9����5�p����Rݴ[]!�:�V��~�WY�Ƅ�un�n�oUK�dᩫ\n���e�/
;g���x�4e�(�7�\r4�9�LC)խ�_^�^�[����s��7��ǷEq���qap���SX��k�g>-]^�f�A+���Y�	��h��b���!���6�0c��T��nQ0Ꜻ.N�����yf��0�lX��v���+��&u�|&p�Iu�X��$�f滺�Yn)��E��仟F_k{�5y4��'�l�����[e��ٲ��T|eC/Z�.��-ނ��2����ـ\���%�J�JfVXQe����͸�J�C�5���Z���<ܵ�V
�
b�fU���w]r�$UGlfI%�v��A>$�/�6��v�a|�LBie[�V���L�%	��Ft쮠�;P�͹ڞ�P��V4c�>ݏc�gY7Y��.�[�R}�Νj�0��%r����\:�ot�['�\6��*�N��kΐܕ��'��&�os�©q��Lu����3�s_n!��r�R��NS�>ꜳ�:�2�4�r��v���7�������]��K	fKZ�,N�V%Ifq�=�N45,�}p��tB�Ŏ�������L���]�������{T�(}%��u�p�����$�vV�Ov�&��_i�����P"]���,�����ub�6�F��Mvt˾h�X�R�5�յ�.���?���@b��;�|�T��'m��yZ{�v��dg-����i7]m�V]��+�$���]��<m(�уq�5�	��dY}ձ�'V�~tW�f�3jޞ"�4�3-=Q���ۃGU��cS)S#6���0�Œ��Fԝ�%.quZ��W9��m\�8�*4�--\�v��[�@�$��\A�2U��/+k>w[w�	Hg
w���T�2r�:������[[�� Mp��3&4��7e��ԥ��n��=�KM]m򂻺v�gh3j.S�!E,f���D5�-�D��� ^�#��묆�)^�
s�a:���e1.�ng��>+,d燀�`��Zqn.;c醹gT�Lܣ&p��2]��C��2'�g-���l#�`�tñyӪ����7���zy�k�s�M=���o��H�|s�TpKj!֕�\ٰ*˥V�;;޾5k�S���jWq0�j�V����n'9���7����{��U�xu�@n�Ρ���ǒ=I�=��sN���ݝR%��9������ t��n;�f�7�	lCm�i#��F�G�`'��i�/z��M��7�r�9�t��U�K̙,e;}�pǋd9���A��Y�O+H]!ׂ)�s��v!�EK�V�`��U��$M��Z�{I��SB �ۆc��+-t�aR��yW��{�]�pr��B�q%l}����Da� �ݚN�%�r�@���q� ����]��A�����EL���2z�xÖf�'vji��5�2�L�Sn� L:q�t)[��!#��
���Hlt�D-��v/��s��HH I�"��p #�����~?+{뮺.bló��B�����e��L�G�;qb]�Ye)���H��I����<wS����K��䩰�7��3JpR��הD}�w�c�W5�|[�ӓ�O�{&]Ө�v�̝��;�X�V�8�|������+CN�#e
�ո���Ԡ�+�A;��sp�ݒ1}J��Y����玕g�٭-v�r��cڑY�]�M�-�+�O�K)v�-��wYZ-Ө�O(	"�e��0%���Wy�)^�}.P=D5}p�3(�4�N��R��O�Gy]e��/GF����S�����_2Ҽ�^`LX�����%�y(��X�\Tζs�,�%�H��S��e��ec��,>YR�VjZV�[��[k�z�@���y�@E��+�fWWJ���˯_����;��ƫ�eu��!4�e=���;�n_\"��R�w���!c;Rk*��٭�9C(��oCv�a�e!Mh
�q�r]M�.qe�"��t�.�gI\�v��!Oo�b4n��h�'[�Z)(#*bPyGHװ������t�� 'K7�q"�qR�{}ۃ�vcĚgg-ol�z���z8�L`�5���Y��c����M�����v�rL,u)��,�:����܃	]I�v��|��{�5>o�=z]`]4U(��]ݴ�8A�����������ُ�sx�ڻ;���-�K��
�e.]x���B?A�D{"�0!E���ִ������TQ�QE�+FҢ��DK���}�ڱ�t�m�{˔��S2�2��%Ģ�)��Z�TV�[e�s*"�\���~K��kl1�QEb���q�m�8�F"6�r���U�LRcKrܖۘt�=R6��a��±V�,m.eȰ���Jم���UFی�QD1��+Z����V�bʬ�����&Z�ؒ��h6��1b"��Sb--�ŋmV҈ތ1��:�pȨ��˔�l�Y��l�1LAfR�j
���-�[��X����J�b̴V�E�ˆdQ�R��S�%�Ŧd�	�fTb��V�1�KmTQ�(��pq���q��bcT1��\q�֘�Z�m��p������)h�m-J��UKK2�aQh�k�KV9[W[-��,�����*��Q+2���r�ب��P1�\-���E�cV�mAV��� �-TfZ����e`��n�<�d��^�[��L����r٭��Y}7��=�\ǝ�_P�;��,X�v�Uq�\e��9�Yb`c�&شxv�.3�V�>��Ϊ��1t��&!+�|�����٪�x�����&t�Z�c4j �����4G��w��s&�-X�oi#���X\_�WL(s(c0���X�u�d�_w��I���>�7�����׼��*�~��/�)��/܏E*�5���X\� 6
�!j!L�B����
f�-Ha�H��7e�O�)��ŝx��)B.��Ě��ѡp�V���ʾ�(��냩��e�����BF�UdC^x�Z�ׅ�g��'�����hӞڀ�z��_��8WX��
���].��]
�tY��L~�A���(c�,f�˔*�n�{�]e���qP�4/A��!^��O�;��I+i��x0��y����c��ݕ5*p<�@v�\fZ���չ2�=Nm�D8ۮ	�u��BuB5l�(z��&V��:2��(Eq�F<�^֗C�5���}M�Si1�%���&�G�ҹ�A��uL\=t��b�Pۛ�ceB��ٞ�ȭ�b;�v���Qrr�T0�za@�;��gD����AҪ|X�.��a���O=��P�k%�F�h�)X�F�I6�]B��t?K�}���m��篝�3)<�˳3�l�����Z�˖��)yL���\83���;9Ռ�ً�84�C'���s�� ��dv����ِp�$��{`kvm���ewv��j����d���9��cs��y��)FE�G��Ic>���Mu*�<�&��Y�{d1P���sc�mIùO_vy��{�Ы�*�N"�htvJ"��ٹ���D��$!L�)�Ł.#�#X����!��G  RVz�p�^aV>l�tu��[�������Yx,i~~��y�Ӆ�T"�2�g|<-��w��L£P�����p+ǥ[��z&�j���ɴ''z�����c�#E�ucT�X;�50`���M���%
�ʅ
���1�A���t"ow}�g�������/s_Ib�����J���K��f���6���8�>�W�����(?
 A�%Q%��uP����CrQ��7q"��fT��.�!z�^��Y6{�5�'7��J^WT��H�#�ߤ����M~������})�+Ǭ5�Ӆ�rR�+�KݻP/��vc��S�p� EP�r���6�#�uK=U
���㽮|���3�	*�j8��N�@�nq'"8�5�TŬ����G�K�x鄖W�Or5i;ޤ5�*gn]�S�6�#�oSǉ�f�����$�<�rg1�ϭ�A�wDc25㼓+m��F�9�Uh���f���M���b%���_���ht���wF���Kŭ-��a荚�f.����oY�gm�b��j�C����B�`M-� ��yKA�;���Y�4����nֵ�v�猑͑���97�V=�^��T������Jw⥊.�d=Ɍð΍�D4�f�M��h7G�%"�|&�'��uk�P�MtU(8k.6��]ȱK���{�nK�(ve�����!8��b��%W�1��K��/%��*{F����8�j�����y�1P�<�#�sP��g�r�
T��C,Fu��8C2%��d�l.<�����T����G!����M�@��:_�}0��ù�*1(�٘f	�['��A���b�֫�NE��9BNJ�FtVV���c���Ւ^7�4eӻ�U��6�����roN$�:�tӓ,;��N̋����/)����ieoi��A�'��4��ʬ���J�&�ryw��������WQ�P��J����;
���̡�x�a��gכ��ue󗏡�U�9c=���{Uo" T+Gk4��\�.�
dzgq�r҅p�Aa#�:��3���1ԩv:���N��/V�����Ui��4�b ��z�F��R�����;�&�cw�iTJ��x��;�k��M�L{l�8�+U��� /��}�kg�}�-kO.<^,�]t�E�J���Y�WKou�'9)�ޓ��Klg�Y��*b�D;�b��I�<KK�j,WS<f���x���|�ܯ�R�d}<�a����񨾾ݥg�M�SMy\J
��!Y�K�5�@4�8k�&��oj�����(��(ؽ�RMB,0�:�ے# W�xk��q�@{(y�qX�]Υ�?b�s���M9J��
Y��A��{r����^S 68��
�w�G-������ ���^�����L�>��Ql����x���H��Ցpͅ����r'�9��S�6�ohC����tխw ,k��^Y��d�[�4uu3�5���
u�u8�"�е���k{	��إj�T¿^��̌�bᄿ�����l��u�h�Wm����,�a*�'��N�b�q�[w�<�&��7N}1U��pP�k�%a�K��s�3�[�����m=}(��\�jPw
�\<E��1�z����g� �E�s�z�N��t�ifbL�Y������$o�D�M��1����e���T;�:�n��x�nR5J�f�˚29yɼҡZ���o��0�Q�{mVvlΑ9��]�k*���i��X@�qBS8�]3wE5y�Stιcz���Z�s���� 3z��Vt6�����
&���={�포����͢����S�'z�����+YY�5(4lHb��L:�U8+�PDױD��Y�Ɔ:
����p2������o}؜p[�sdXg��Ή�_�=%#����0p�]g��f�A�p�;\������j�Z��iD���E�b@������T¸���Ȃ�ao�8�y�����E;�Î���*�U���@�r&��GĿ�}�R�S�5	�v�QQ��g��w|�h��@�θ��5�lo�Lޜ��vbE��f��
�k(���$"J,*1J�����c��r�OfH���/���W�X]���s��a��Q0�]b���y�ʚ�ĜY�B�s8pu:��F)�0�y�*��z�;�vXW���V�̗k��軆ά��}	h+��`{`Ln��9%���l�Dbμgc��q��$�B�hпE@�̇|�*���u7�B���>�Z1�a��k�G��xK;Vs���='M��~p7K�X�{*%�>�h�d��i�mN\�x�Z�6��ЯmyQt�*�����z2�&q|�5_r����_�@.U��.�rYJup�&����<�X���OF��6�RS(��hwƮ��ٵV>�%2����j���>��S�Ϛ��Q��W��c�te��HD5���)��z���E�ie=��mW0>������+\N���[�(��Y�!-K�f�hS���2qf`hvN�&')�j��/����z�������_���n������;Ն:l�����[�m�y�^���g�z�d�CԌ�L^�t��kk=o�i__<�gv��l�ΩnO.��;G'��	�Pga���HR���w�[��yy
 �	�=Z��#�w��Mf�00%G%T��GLW&1Cc�E�0o��i:3��1%m���9��ZV�J��bƵPM��NHmF��B;�����"��V���{�)5X����R6G5:��xu�Ӓ0˔��V�2Y��aZy��U�W7�z��Wn�dF����Aе��s��H���0��)"�-'�����,�M^�s��w�Q
�`lU)����A�?+& ������+b��Z�V]_XN�79�*�uj��B�l�?:Ո��,w�8�F��Ҏ�ڶ	D�g��z�#y�Dr<	�l��7ؖC�]-�v�/%^��s�Cz��;�I�Qp<�{"ޅg�&I�%K�m�M9�C`���5�^��+뽂�^�$=ӆ���W�,����`s.
}%]f��=w�H��N�;�����W#���S��C����i	��y�R���hu��juM����K[���%�8���=;z���O�)+�R��w0U]{����j��v�79K%v��?o2%k�<ڊo��<�[��{ʙ^)��;˹<x�w�Ӝ�z�+f*�m�oiƬ}�����+��-ϖ���^L\ҝ�{���9i?S]��m�8�mc���V��f[�^x�v7���e���백�������}����u�.�¥���T�G�g�'t��WZ|���Eeʠ�/��9,,JN�Q}	��fX���^gjr�ںN6v��rYp�ι�th9��*�J5䨸�bET��{�2|�����!��7��.��b�ԩ*�Ccy�=����ۺ�5��viWD���i�YF�Ý	�x:�g�+�j�%2�.Y��8I��}�LHюk`k3���>5�X$��Ƞ'}S���:��D�Z���7�ב�4��vt�ˌbrT��+��Z�9�nN�E.|�gb�0j}Q�'.�KS*N�������x��x�7�n�w�;��#^�(E����x���=Y�V�^��3@sj��4y��i�{\J��O�m�J�����Oa�T�q�W.�C�L@M�啽J�O/���������ӭo{��b�N�r{��6��Z�����>���Q��x�Ylw>J˩8\�1���O����Yq��ͷ2� 
C��}5Y��ѯR���}���]s_k�e�V�_����S@�XZ媛n��r�Og���TU����Vk"b9���ʊlvE'�L��cF+� �jNM�.7���P[5?iռ��.�y�+���Sa`�x�9�nj��c�}�x9�KoW��3s�9�J���o�<��pm�R8�q�ԙ�^�Dup�~�U-Sa�����|���Y��ޣOW�[��7w��o���΍��龎2�;���_���ZhĨ��W�*j�F��B��$DЉ��6����d���G.�&���),m]59Ys	�ɿ�.��	YR*\}�cC���A�zڹ����)I�Ɗފ
�q�f�J�A�R	Ե[�%���I�i8��ne����C�^�7�;�5�����Fn�ݟF�,��۞�X&)���Q��]B�f6��u��&�T�C�J����6�y�y��-c�йѿ1�"�����/qn�59;�b�,���m'J]>���ˉ�u���w
W��qW_:Y��9'��C�ދ�6�r�:����y��myR��Fl8�����*�w�\:�3����{�"\t��!X�����z�-�����30� m┃�8v?*}�6FZ�'�N�5��
�i�F�{}-%܃vyQ�Cސɋ=I��C�nTC��*�o��+z��M�\�@,]�:1��f���omE��n�QG�o���Q������[���� �x�����I��O;Ƶao����i��s��v��%"*5���77Z�Nja>��Y�OQ�;h���P���Dۜ���]C���t���ʹ�U������=ztt�!�kGU���rvO�=�T�yk!�s<}��YsOk�h�-G����sn��,sȒ�����w�ox���l��Pw�GR�-L��4��r��8�z�V�焸��$��{jC<��[�y�#�ӱ=��P�O$�$��W7�Mg�
�7���TSc�I={,�G9ɒըjǒ��nMF��]P�#)���<���w��I��gS=UЁЮ���V��͕�6V����{��t�/���F�Sf��	��6���+7w��wA�v>��`�s���Q�-W���w�Hz��K���GF�7Fr���׵�~ծ�8څ���6fNr����ME�\P�Bg�l���w,�~�Ɋ[]:�(��\�m�h<o3�M�їb�lh�O;/D�.�ݪ+������
6��.��������W{����_n�O-N��phn`(YB^�P�&.���$&�jt��k{hgr0VEef.�uW)_>]�g���05PrUA:�Tt�rc668T��7).tJ�B{��-��-���#l`Q>��']�������!�P�������Ƨ�_OX�9��3E��9��'n�!���VP�܍�r�+������wh�vR�\	�78��Vcwq,j�/��+�:͝C{,��ovv�֋l�wQZ�_F�32=�i�4�yN�]��HqV&��w�����i��sR����׹��DE����.k`�ؠ�����{˸�F��a���U� Ոgрp�J��N0�fk��DF<�nes�&�I�jM��P�wp]��q���g5���ɤ�/u��������%G)�+�Yj�k{V%ǁ���Ѯ���:�g<����{��L=Mp��gVqɛ-��4������V��k�u9V���f8�������J�]���j�([n>H����Ȫ��%9�{G�eui�PkB�U�����`qfYn�K`=WDԮ��J��Xo��{C�R1[3�,˭gK�T#�-�ل�<�����`��>�F��5���oT<W4�.\��(���h��LU��y���o\��n���]�q����GX��Bcb�pϒ(�Y��,B+��k�ss#��NP7��#��3��Pໃ�Z��V��W�r÷K����a��%3h�������[v�<	��Ν&J�:�c�ft��V�.�����)���>��w�M��̫T�����!��k��vW��W[��;LK�����1�}����-�����L��KA[t�SW(�v�o$Ya�L�&�%[���q�uֳ�P��U��9ͤ������oRu[5�mo+DtM�k#fWޏ�=�L��i�^g��"�u��\˖b]d�3y���Ž�X=�!C�np��Ϭ�ڡ>Xq�1봓}3�Ew��g{�*�ƛ��wf[ޒi��=S&,8��'�;(W[K���ֿ��"E�3���eTz�u����V.4T0pŷa�ѫ��Y��:���%3�FQzSFK 
�#�4�`�uy���.���N@���:�����ٰ��yB�-V�˨�U��6x��"�_V�ˡ�iw�X�䢎�tr0_a���������-�ܮ��:�ơ��{r����cJ�'�j�R�jl=���{|XN�pCN��"��)f��S�NV���"!Hu�7t6�&������X؏U�u��Sw B�0�M�v��Z���<�>�"�6�>vy��>�[�d���6��J��I����{Nވh�D�[�V��榴�|hj�Y��Wgvn8�+��W�x)[��_�񚻏<*��mqι9><tS|�N=g3�jZ�7B�a�Q��z��]FvX�s�M\��05DJ�죚P��t2�u�Уa�^Ҭ�\��2����2����s�&� �W;N���`]ӻAˢ00�k�o'{�ϳ�Iu�ǋ��nψ�x�%[�$�?>����z��#�K�Ow��kgK�I/��[%����=޹˞Nk:�S��ٳ��ʈ�QN��c��s1[*�b�����VօeȸdU�p̷EG)D[j�nu����<����)iUT�3
�Z�8�m���LŠ��̸�ƹl�1AEʹ|���F"��!ZZU��a�	�)m`���`b�.7(.Z֢bT�Q`�J5�؎\I�Lqf+S.%@�J�\���FԩQQE��2�E,Tf9����"��aQB���c�W,�̮F��!Z��)r�*9`��%�1�ŵ����V�QJ��2؈b[)E�RT�3-eU�*�ZZR�Jт�a�",lĨ��Ѷ��[j*
(�mim���1�%X�EJ��ZъE1.-��F+
6�L��b*T(R�F(�++�e+B�"�e[J��*1+**�k�(
���QaU��̕�6E�(啘��ʖ�aXJ�ڋ��W�*#Z ��"���b��R���ܢ�����#���b�J�,Z�"-©�j
ps5����w������:ۿ`���(�g��@�pV*�I'�ۮ�;Y��)NW1���;�#L���J���R5W��%�')=T��|f���y��ٖ�sˁ��ғT���󡲤o�Pq09���]0o�UGok�\{#K��5/���������g��m��շ�����C"�����nȄ�Y����
%l������ȷx���'n9��]9ʕ�5׸��#c�i/k��!Ύ��׽h!0yp��m��ձ�k_$]_XN��T>�(pn7+��Zf�V���혎�r��	)�����O����w���F�^v�\��9&x���U��u�N��Uv�mK ���^+\�����s_Ma߮\h���.F�j�Gw1ɹ�'J
�c�J�Ub�Fð��#�Җ#�Z��Ra���"7�����M>����<Z/��&2��X��ף�Q�Q����&�؞Ur���ӫΧ�u����>�
��(o�Q%��=�V+�=��'u�GI�ҵv�ܪ/UE����_�u)��}\�jևDe�"�cP��6��WY������h���1��j �]"���Y��j�7}�p��$�\�Dŵ�����a�͆�ܤ���ٝ�8��3�^x�s[F�Ao�P��rMVII��p�(e���;lL2��D�:)�{zy p���*��is�&cv���bzt�/�vck
��.������LWΔ����4����ׯ2{�Mc��x�j�!��˟J1Z%�^��b�OCq��{���2+yFp��p�ӱ�e�o:�׍=��w������cs~��MI���n
��B����ڵ�TB�����Ϗ���������V��|I�. �U���L_CYkB���M�ȿTs�or�8cc���h�\���:�\}9:�S��Th��.��dF�����=·�1+[���9��Pz�T��b6D�G'c���|�%���뽲ںC��6flz��m��C8���ڈW�Eo.�0����v��C>}���\�T���۽��W� �^�9���ne�)�@$8}=�[G�U\m_w�I�c���J����.v]5a��s��Sx�2�}������y��)�ث뀛�8�ҰWjU���x�y]E��8Q�]���̳¶��Fb�P���ܜ.��j^d��+:b�j�D~��<哝��s+��rM嗋9�gLd]z�x۱�o8q�}Q)�16��x�˩d�J`�v���tːǽ;�S�<�I�JL��ƕf����ȟsm\*)���c��go�R`35�ڐ�|��E���].sWyk#{��o2'�\��T7|�������ZYS����k�6���f�uu)E^;Y���5>���q\�M�8g�3�[�^H��~��9~z�>�o�m���uQ�r��^M}^[�H�����'ܻ�J{J{�|�o�oW$�?-��I����j;w�]T>i@���P�k���N�K��m
x��EeϺ���*��˭ޡgO@�Z��ݨXq[%F�T_kcg��s�|����|�.k����⽓6�ju=�z�Vh�pnXHe(3�����ԅ�'�/��-��᛫.;��^r((�/-�/����U���C����㫒�P�=�M빚8��h�nnr�{_���t=�P���H��ߞʧ~�G����&C��r����+o��+.h�Z��+n�Jl��y�wVkQ�����T�ʉ��l��pK�o+�|���HH������Z�����.��K���q�����D���Ѻ�]���{r���L���o��fZb��E�wZr�hr�v���Sb;��@]".��~�}w�nS��T:y�a�U�(��V�Ӯ��˙ۧ���۸��E��e�S�O>Y�x-�Ѓ��J|>ZF�1Qn�kwms��]�^�ެ-�.���;��7[6����s�}�H�gni�.�ZߜQH���D���E���Q�4���\Cn����͚+2�V}sY��^��|
�{@A	/TԪ�Ƶ ��x�NچWó��c�ޭd��63z�Wr�AN�U�mc��0�J�1�_V���w���׎N�yH�W����ݒ�)|/ɇ��}��S�a�W�]-�ʜ����=�O�2ݫiKVw?$�R�ac�o��}�>v<>�$�l�z>�N�8��M���\y	�3Gس:]��G����w���'�>I��y��'^��z�ѿ��	���d�T';�������<d��g�&�5凍���b9d �/��L���՝��O/�޷�N��Xx�q>gv�I>By��z�2m�~k$�2q�{�$�!��2q4�=gf�Ì�J��<� q��i<��F���gH�(�����;��)��MA���4�;��t�wkbҩ��g%��c��jr�w�����}mu���������{[P-�jl�(���6�2G.���t ��K'���־ՂlN�(75]`��8�s�Y��]z�oc	���M!Υ�[3wk�'�}Ϩ7G�6#�=����p"'L�J�zͲt�f�'�Y�5C�8�tk�P�h,����z��8���Bm'�7�N&�'���a�M���_5���5c�}nL�2�~p�;�p��{��{���=d�:�d��l��<jN�m�2��:d�Vm���N��$�
d�&���)6�l����6��>뗎f쿣uU���ϐ3j�p��D`�}��6��y�m���|�m�Y+Y�Y8�hVC��M��S'�q5:�����6�Ĭ޺�]��Bڡm$�E�q�#�#�x��3�ނ����8��q�r� ����M��'Y>�M��&��IRz����lRulP�&�YLd�����w��:o�a�r��jE����"({ޑ�N�G�����y��6��hxs쐨L����>d�'f��8�'l���!6ϙ5�d+$�7�J�ԇal�
ɴ������]/���5w��[|�p=C�N��Y'q:��C��I����m����l���2|�w��M2t���x��;I��s	6�2h���w���]��vҔ��.fg�}" �!�"��Å�q'q�0��$�tk�'�d�f�{��'Y���N�P�>ɶOM��;d퇬j����zín�[�5�ܬ�`u�~�z�p���@���Ω*
��$��J�є�m'��l�����&���xB��q��s{��1~>��X�ywq��g�����������O|�Ϸ��4��w��z���I�7Ւ�a5�m�d�+%I�2}�<:��`a�28���Dg��zB=c�59�D8�>��ߒ�ʳ�[4�c<a���OO���$��9��t��5�!�<d�zæI������I0��
����Y6��':��1=�=�C�VП�|̊���إ{��xMj���$[%]vì�������P��[����u��խ㖯�uG�����{�Ӗs3
������ۋZ��V�y����>��k��f<`�&��y�3Qd����ss�ce��-v����x�E:tA��9ø��3u���*Kv�����v�R��l��y�{�G���!]��O=�2LJï��q��5�d�M��59̅Ci�Y�C�<I�d�<B)5>�$��&��,�3Y�c��a�������zG��Rrwa�'��A��v���$�߲��'�=�8�1+���Y�'N�m!�9�ěd�+��8�ĝy��G����k�9������,�/���N�{Bv���ԙa�$��;a�'�Nӌ�I�j��2m��ԓ�8Û� �LN���>J�s�;d1�h�=	{���J�&��oW=�6�o�TP9��I�&��.�z��je���&�P�	�8��a�a:5���8��<����4���u�'�q�ܧ.�}�����ss��_��~D�~�2v���`x�l���������N�u�D�M�5<��2m52�v�&���l�ĩ֬8�l'F�2$�
�)��D|=�@���L*Q�e�L�϶3�~�&�mO���i$����o�	�=Ì�d��'��<a;z��IY8����t�hh2�xΙ8�2ͤ遢$E�����#ޜG�"a}�oWp���~\�^�C6���v
M��=Lg&������Xq�a8���d��	��3�'�̝����I�Y���q���=J��M�Yd<gL�N�w�}w�h��ε��Wϻ�2OP���)&u�P��iX;���ҳF���t}̜��8û����O<�d�}I�d�dy�\���z8{аU-�Ҟ�ӷ�oG8�Ҳz��p�C�t���SN!�k�p8�d��>�m�iXn�a�N=���rB�q�����m��N���{���LDBG��>�S�f	8��S\��Ͻ�+$�8}�IXv�tZq�I���2q4e1��&�]{��4�c��o9����N2z�����g�{��C�˞���f�\�r;$�	7-R!�(���G3���n��ý@�캟z�ܠ�{��8i;ˬ�Ġ�L����G������c'A��*���W]Dv��+	��/��6wΞ��/e�E?po����r��'DA��5� �0NI�O�g��yy�޺�bй��̣�k��a\����*
=��*M����>I�N&��O�m:5���	�w���*|cч鈱�����\4�LJ��%��>l�'�'>�=~d퓤���$�m���{�y	�4ɩ��,�ho�%ABk�>B�q*FP>a�O�XXM�q:׳�R}�1�21��j�uЗ����H��_rC紞���''����a�N�O��0�&�x���2N&�=I����t��sX
I�:�$�RL7v��|��I��=y
�����ɓ�f�}�����tɉ֬<�O=a�7�+�&�׻ɴ�w�I�I��a�z���<�0+�z���8���sX z=��W��x���R�TW�M<�/&�/=�^�zo�sVO<�8e'��2|���m�޽���'8��7�+�M0���u$�T:��8Ì�l�:d�
C�s!P�OY��!Ğ2}���yOw־�w�y��w�y�2ORs��$��ܑd���)8�i���6�t���N�6���d��������I��t�'�LN���6���=�ߩ�gz�����Ǿ}�T4��T=d=a�'=�0� j}�I{�Nk�$��']Xm�S���6�u����d�y�y��&�w��'�T9���y�z����V������}��
I�����M�Bk���&�=Jó�����u|a�C��wd��zɶT&��:J��I���:I�	ɮ��4��I�o˛��ѳ}fs~|��n.�W���G� |�c�����98��z�7gm����;I�'��<7@���N��x�6ɣ�O��N&�������I���x�����t�s�wY���g�u�V0�j��L���s�`(z��6���&�q����L��w>�N$�+!�)�N2x���TN޾�IY6��O���&�ۧϧ_f��uy;���hU���3v� I3�64�i���W?~F�X��K���;��b0f��)<g�ɏ�b�����J��\s1�
E^��yP�[�l��ti���1����Z|V�gJ�����<] hQ�j�<;����ǽ;��ɱ��/e�nC���L�����֬>b�:���'Y<���6�ĩ�Vl8�龰�i��*v}�N2}��s�q$��G��}�=�|'���;�q[��n�&����e��xJ����VN�|�d<Ld�<�>a>B�Z��
I�z`m��R�삓l�J���!6Ì4o�8��8ù��|�_)=d�:��{���Z���뭍o���i��5�����sij��!հ�+'me���m�2�$��h�È,'�F��m&�X���'9�<�$+'[��sOW�t}�|�r��^�|�xÒ��q�'�;�x��~d��d*�7�J�ԇe��+&�Xu-!�I�hˌ'�6��P��#eO���#����ݳ!�|9O�����'̛{g���������N�;�x�;I�s���O�9�%I=g��$�,&{O���AaԴ��m��_���=y�w8lS�W�`��]���p1:a>g3̇>��<����Hzy�6��	��xq�N�:d딜f�4ä��2��&���&���$�(I�B �{�DA5��賕��}��m���<d�8ad�a�u��m�I��{�m���m��9�I��)�&�O>�x����y�d�M2zä��}��z,G�였=�1���?s���f�������ܒ��9��%d�'Y@�M�}�4ua6��:��8�6��d+�'�����I�l<�a�I�Ǚ:d��>��({�" ���NF��[2��>�뿸�=Iϵ���$��d�*I�]�T�2�u2�l��q��Մ�Cy�O��d��:Cs�r|�bpz�,G��1�\>q�_u�w���'�R��!P�'�,��'񓩽a�$���+	��YO��:�I�IۏS�2m���}I���a�z�"�����۰#+�CJH�FV��}Er�4*qiI��ٽ)�����r9�;Mo?���fe�����؈؞cF����=�����X��$�=|y�ӛV�ml�������2�z�f9y["���=��#,s����:�Wt���hM�]�����ؕ�=�Rq��>�:d�Ӝ�T6��V���O:7�:d�a����$߶E����P�$��5݆�6�$ڢ����q��Gͣs����B<�y�>� |�@��x�z¡��$��ߘq��9C��I�*�Hq'��u�I8�����$߶Ol�Mu��o��9����p_f�no/�#�B����x�u���d��xO{���8���I�C~ӈ,'�s~��M�Bh�<I�OYP�v��2u��I�'�6�5���3��#���1D�D��&�A�0�&ٮ�i'��Y�M�@��d���N ��I;C�{�2q4�=gf�Ì�J�痈d��GVVI��ӿs���Ż�z ���M�{LwI�Rt��k,����IY�I�Vt�q	׵C6�ɾ��=Cl�J���Bm'�����$��y�g[��f���+s])���!�`c��9�={I�k��l��Fk$��`u�'�I�M�S(O�N&��l'�*u�Ad�צ8�ɠ��"�i6ʛ��a��}�b�n&�!6��X�1���X{�$���d��0�r�a<|d��d�2M��d��������a�<�!�tɴ�S'�q1���&����}����뽛�����u�6���<�)8��T���
��}�8���N0�z���'f�p�̚�M��%��Rz��Z2�m�N���d�l�ή�]r�x�Pin}=�!B'O��P��#���M�`h�x�q�����%B|u�=|I�'I;���퓿xd&��&��A��E��x���V���	��f�}w�/�}�'HVOXp�����I�O���r&�&7�d�� 6���y�m�ԓ�|ϝ�v��'a��_�v�O9I6� w�N��u�G�;5�O��`��4�-]����8��v����Q~rq�Y
M�"�����z{]�6�;j��8�χ`��q�w�����K/�L]<N���O���p/V|��v3�#�N�8Y�%�j�������vOQ	աukb��9ޭz}��{���w
�tÓΰ�	�vq
����I�(�|���re�m�;��8��w/0;a;}C�>ɶ{G�֜���z8z -,�݁3Q_��ߺ�<�w��'���}�$�:d��x$����(Ln�VN%d�($�O�Fl����!�&ٮ��+�=��s0ǽ�
�c;J����_X�Ϭ�OXOx?a�&�x�ٽ�8�2zŜBq=�I�:7���a6�aY>J�ٔ�@�'�SS�	����"=������pe]�#IZ�Fv}�
���>�0�Ͱ�)�d�9Ld�'h�2�<Af�d6���2M���y%J�g.�VO��5$��{�=�Ý�����U��D��9�2v���'��{����v�S߳����{Ì8�t��2i&�R��B��OY�C�;I��ēi=՞6}�0�
ߋ���}���%j���<����d���jya�'wf�4��=���4��;=�8�1+���Y&=}̜I���9�ěd�+��������e;,|��*�a�ٕ����x��{�+�I����O�Ya�I��væM�k�<N2v�l<����4ɶ/~�	=C�57�Ad���!A�Z�}����(���D�EOR����<�̒z��"���M����Ěf����q5݆�m����z�d�N$���O��'{u�'�#���Ƚ�n�o|�k)}C������l�J�j��d��'2x����ɶ���2m+	�ĝ3ɖm�x�4Ì6�y���M$����[e[�_lg�l��z��p/9}�P��O�xk�M���q� ���Ì���w�p�'>}I�N޷���q��5�m2�xΙ8��d�0D}�eG��֊�J��We���5nJ�`�l�Y�obIN��h��ʙhSL^9�>��mhp�[���we^�y�x�%]��2Ѩ�a9�u��,{-�Z��-DsO4�b��X��["=Ks!mp�w�D��Yj�INa�1>	XD޽E�6�m�1fjt%��ӕ�L,YYF���T�1^)�H}��W���y��.9��.����Zk��f����s	�sD�W)i���_g^�`��:S}�饮ُ�5�]F`Yy:�İR�0�)Be�ʗ���{�V;�R�$�yy��R�J4Ju��o�dbq/�66˶����@]f�}�Q����Y1�Wu�E��~ծش33z�
Z�e_i3��D�L�iƝ;�\���KR��#G]W%HqB5X���i��� U�ݺ��D�l��T:"�Xis�5�.��MN�&sF�J�w`�2>������r����::@N�c�s��So���͗Lӱ1Z�/���tg\緂��Y`qSm��woN[(V��Dv9{�%g㱷t�1��p�Ytg__v�gJ.�*�<�.D��f�s��iq�oF�{r�/�n�t��ꘂc�\I��fV-�n��z�M��d�Zy��FI#zӕ�U���6w�D|N.8^X�%6YY��c̗v>�&ՇcP�GV��Sgd5;O�j�fW.878I�y�	K�wY��㴜��M5��K����V�oI��
l��l�ڥ\{��<�q�Uej��F� v��|�d�Ӭ��ʈҬB�b�_��_���ͿԿ$���u�\��⡍B���ä.�n��8�G�n����Rw.{�fΡ�z������3%g4���:_~��VD_�|J���iX�K�sZj��=�%p؏o��y�hu��������q7���� ]$�y�G��������՜,�y�;�5�S�0crP5}x��(eC$������>�^�[�}��7@�!�H�y�q�iGM9���4V!�fK�֔t	�Fa<���+��C{D�p_kf�������Ji��� �}m��(�Vujt�u$v��;���-�蝡;���Y�k��m���X�6��-u�i9n�\�c�w-YVZ�,0�5��PU��
��}�Q��h�L������MTɷ���OA��{;�ER�+����<k6�4�y��C"�W��/-r����Z��ꬆ���{�;0�Ѱ�;�{6���}�i+���2��v�MZl�g���Ϩ1����qu���L��\��Oi����.S�}��!�6��5c�0f"]Xr�}C��a�m���5��P��nZ�N��l�����*a��0%����3P�Q�^:����ؒ�ڽ]�h��gOoRs�&����W��L�h��ܘ�*�c�1Q�wt������g��qyܸpG&N���'6�<���Cu�����@�������׃���?䯛;d�˙jZ�cX��H�ʱa���KVێ8Ԫ1In\��\�
�Ե�Hڰn~=�}����l;j�̵��+
2�Re���Y�e��JG*+mYF6����9J���}�:c�X+l��N�X�a:�]Z�:@�B����T�R�zK2�L�bU̵\��oYC-�N`�\E+\C��9B�hQDƕ����D:C"�R�*�*$PU�ʘ���V�AƥLql�+RQ�Q�XB��z�*(�ҡF#��TFҶ���f,�[i��1Z*�ӌ1d��
�QDdPF-�iFڸ�&W���&"����b�˘9+��mZ�k(�,[�cW-�κ��[G�!SR��mX�Q\̓Tb����-j��X*�+�[E*j**դ2׫\��D�Ke��H�(��W)m-�Ė�PUF����Z %)+�Bڈ�E�(��X�E:K�he��fl���=Z1�܎�q��c�k��r.�v�Y-W�[����#
���Re�UC��+�\�|���
;�������sr�nN�1��D@�}Y D1�w�AI�&ҳF���I�4o�8�0�a�~Ì�|I;��N0�?2w:�I�$㩚�+'O�z����g�z�8|���ޥ����z��z�G��m���)&{�2q+S����m+5�0�@�}̜��8�v���N�;�d�|I��d�a6�|��y������\���=����y%a�!���VN�|ʐ�d�*T��6Ϻ���I���l�J��t�2q��$+'迧�q�1�P���}1��y�ŽG���}��{xo;��m�'�RVI���RV���0�8�ëH|�8�+	�N'�{��4�c�>�q�~Yt4ɱ�|0Do�ހ"=ص������ϵ�9�]��x���'I9��<d�I�9��f�9Յd����$�(L���&�Rt['�6���I�M���p>f��7���;�*~:�B�$�^q[�f���˦���Uy\)�7��Lc�un)&y%Z��y&�<�/;:�MYu}a�Z˜�ˇP��^Hpc&@�}-���7<�'Q�����w�UF��9k����	\%P��}�.�J���ms��� X��<�jQ����
W�Y�W��Ey���u�Ut�wZ�]�����c��yetG�u������I��B��y����¬W��r�=f�b��ܵ��Gs��]�	t���j�6���Qn�!qyD��_[$�ɨt��@��!��%�6������Ӛ��9�$�r�veJ�]^>�J��T�g��.�vW�5�o�0Mfά�+��c�ovI�O�Y��==��"��I|�g.��U ���.���/ϭ���:�d=���>��V%�GwA����X69��+0��-�~����Pŋ:ҕ7{�+}2���R��{�n6���^�}���vq]��ǲ��N��(�k����Xu�>�F�/+[��N����Ч����HN�Ȭ���sޓݚ=�wh��7m��
�A��j*�S��)t�>�m��I3|�9� f�)�Z����@ٌ�*�J�R�����HR��}��6�w��ME��s/w����J�}��T������x��'Yq�\����eڅ;�Z�����!�D'��-�����م#f�k �U��M>�[WQ*۝\���(<�]���ĬޕO���]Q��)�\L�%U$\V�X5����/׽N�o!���%�i����̾�T�T!z0I+~�T<U�h���x�"�;����
�J��1Eŉ�U� X�I�M쑜�gS��Q� m/���*�uJ$�_�K����)�*�?��HG�r�:˾��v�q���Jj�k�T���Nef-'����ԧ ��gN����U�D����W�7�������-���w�i���v�

����y�����(A�A	<�jV�^���kI�x�]qOc�m���fcü���VB\�T۱BKw�#���X�Ist�8{ƽ�)��Ro��P|W�䭩�mWvJ�U��{R��G<������%���F
yf��s3+VwwqkSP�(�6
�<�S
��Z��{R�!�{x�l���l���~�����{ς�[�Q����+u�R#w���Z�=��+ʮY�ںي���6��^�u��6��)��&���{��ò<��'(�Kg=E�])�d���Ƣ�6�W'[kZ�ݣ5c��|Tޯd��V���8�����Q}>��k�\m';��ӕ7wR���fb��13j��N"���kf�� �}��9.��1J'a�(��7 �qC��
u$w�o.����,���É{���f���μ��k�������o�
�V�B��Ol�SC����;�b�j��R��Y�q���D�Kr����4�>��qյ�9ۜ�g,�u�K(u��X�{Àg�n�joVE�T�v���ߢ>=�g�m��[�1��Z��}�[�ƳL�3}U�9*��0x�t��'���)9}b�����s|��om�b���p��0(l�#I�δ�<�d����
��m�C�ent��(��Ά��}��F�J]T�[)I�Ü@B�b��5�F�5���ި�|�]oU\�X�b�|u��vXz�$'"�Q09ux�9��*��y��Ȝ�"2��h��dQp���rFn{�k��n�q�ʮۡO�z[����C_(ж6�������1�Z����pv�c���n�.�0�P����E��B�Sbk�ֶڣ{H��3GUjE�MC=mp��U+��T�MF��qի�2��m#�52�rb���꽚ȟsnj���^�
�=���ru�-���o�oc.OU�Nb���ou;��D��c�QM��e<�
Lo�-�],���=��>�^j�� �ydIR��:_^v��]��PnU��c�-6�hߚ��w���0�V�\>�Q�q�үy�	�oW6����#��O���F��/5��t�v��N��]Y�yB�3;:�9km^Jp��g�fom��{�~�=�^/��o�ܔp?�6}����㼴���L��/���8=H[�$nnE��!Z��Y�)Xq݋E�d�c�Ȧ��R#^�)�v�y}O�w8�jh�n������Աn���hW�b�y�6Wf	Tm�x�MI�.�k��I+#���
���\m'J]e�9��[�U�*���(aq!��W}����D�jlQ����ה�v9��6�&���c�+��!���лTJ�,ܺ�<�"TN�b���o��
4���FP����&N^�O�l�Y�ҫ�y\�E6*1Cx�>�7�ld����|�Ԟ�gcs�{�����=�Gg�'ù�<����\us����zm��f1pjs|�T6�2�y�OCj���R ��^��r�V�.uGT7[�i�����8��=leޢ�&�]5T�g�9B�x1'�8��᤟q�l\v�r豋��H��j�\1A�p��ċ60�ݵ��[[�
��.b�qMt��gt�+���8��0o�X�o"��`�էaܱodUu\��S����y���S�8{U��-�(̊��~�""=r�._|'�yA?�x�W���/�s]ͦ�l�vB�*n"�R���j��ŞDh[.%�ޣ�������]5��br*�U�۱�i+z�WtfH�WE������+5�1�Wʅ�%t�P�8�z��;��ӋS�]yŏs��c��%����nONx^�V��掎�~���d��Vε���!R�;��{*�t�*���$7lhյ�m84�gs�$�W�86�nӹ�p�}�׫��o�Գ:z2n��R+�k���ȍ��6�9���&�E���ܛ��߽P�,��Ol���fr��u����Z�\m'P��_6���V����e�"����TW�h)��O�D�5ژ���r��_`��t��9�ܭ��;��MfѠ�#�J^A|)A�Lu�$)bcv��*AVf�o�]@�Z��YX���t����}�����2�~�y��z���4�W&*�h�z��'ݴ��+'f�E�k�nd3��w4�R�b��X���V�;cr�a��cj;V>���#�
R��YNPw�]H�q��:��tk�'.����#���K����au_�<�r�����ǥT��\t�$6ΞDH������4s��Qʟ����[�qC�t6b��H֫��ֺ�n�M;|�{���?b�����e�)u�nT:���
�
7{j���[=�un˃�7N�
o���զ�e�S�O��q}�;m�^ٴ��<�C�B�ץ�^0�֢�'�Ao�uuӽ��$�勌bF�v�i��
1V)�q�dC��#���VlE�*��kԚP]4�7�/v�'�m-=��ܕl\'�� 
C�Z�%��k
�w&9	��$�NO�t/Sg��gV��mr�%u ��\�Vg��^R��[
9�ޔ�JTo)l�����D5�My:QP�X6�yev�l�^/G�Ɯ~��.���ں�y�-F��^\����M��q�'+��OUu�VUh�	���<����wC��3hA7�����Z��Z�V�'����Iɘ�V���"�YА���8-�Y����r�����2u_U�4�m���3yw݄u+��S��ք�u`���G������v�$�z=�D@���-i���3���^�
�;�Z[>��O���=Oy��|�w��b�M<�>l�9�԰o��+EҚ�:�/mc�su��*X��<p�]*4Ԓx�s�ߜ|ڪ�uC�h\�y������]Ss�M��5�
��V�ozc�~s�����U���}%Q�tW	�P�Y���/c4S6�R���`�����Mϑo.1�ۚ�F��W�J��}"���;�w4F+�c�r�Cb��>�����f��W���hi����9u�ؙ2���Ca�n���Ӯ�x�B����â%nt��-p�X1#���<�W7ؔ�yz�c�H��aD�j��)�oQ��e�+O5�Qo��p�������<[��涟��T*b�;���a�s��*�i=�U���qWr�/�ϝ~���q��>3w�)�B5,��0�b��6jz��VZ�g|�� @�aKXr�U��Yy�x��|zC�x�6�I�5uē�H����9rV�m���]u36-�@nuq�@��.���1v����-|R
LEh�֬+�~�p�9��N|�U�v�Lܝݹ6W|dp�V����5x[X�u����~�@���]j�6�@�� w��_+����'Y~��f�7��ˠ68IO�5X�J@2Ǧ����R�mT��;��uW�"�;jÕ��p��R��]�F�
�8�o%�7M�D^89�'^_^��Tf�'�r���l,���3gd�#�)׻�s_��������o{����ou=�G-pg�ڌX��W:�8̿r�e����>[�m�2��8�;٥x�e�S��կW���?>��J���Ǖ��K/�o���C����Ǟ�uX�/s����i��j��ٽq���-hS�[�vv�����
�e�٬�[�sT�q��͠��c�F����ڏ�ͭ�z�nEe�*}|��M�!��s&rr�,r'��pS�v9�E�&��];�6�{�\�mv�o����9<�	������O#�\�?�_CB�`���>�
�71��Fn�������^��¹fޖw7D(�a��^�:BzՌ��t�wmt�s֓�xd��\�+�+��q@��˙a�ɺ5���#��Z{�!ϓ'���lX�r7w��,�"�T��No7�_6ժ���J�jy���뼂�b��s�k����	Z�o�[&�;�*�Phl���@j��F�$*#7��7[6;v�8V�y���s����rS�V���j��2�uJ�:�w��e�ֳ!���e���N[��k��V��K���O�nT�>�Br&JhG*�u}�����ܮ���*y�_Aϻ,;�R��M\۶��t�+��EF�bovf���V�l���"N����)���E��q&������s��p�ڡ�6eY�O�\��{bĖ�J��u(�:�5.w]5~�dF���Z2sN�}�ȥN7�7�Ӵ��ek��}[X�CAU{5�<�[c�@`]�*�-Sl�ewd8��dTr��s�`��q�S��f�d���pn�j�{���ɼ!�7vƦ����s�%��Ū��T�*.�p���u7p����)��:���S�^���Z|��y��2��X��^�G��N}s9k2�t�Y��0��=ϯ�\��u�G�)쩦D7z	W��t��2�7Is��3F��'Q�2,��z!��O������2C�l��Ū� �jO��u��52�7����wMLo8[���l���,[����.u�. ��!���PƐ�����J�Wp�E��]+��Zj��ƹu�]�t�/-�ˀ�&�wP�eJ�՚�}f]@P�G��$�)
ym��2+\R�F�]4���f9Myc�]eQv>Y�U(6�&���Y#�]�ڱ�q�[Sp�*����,�����ɶ�^eI���]�u*f����$)��Vh���R��.��u�����ܕ{}�k1J�͡\:�"Dޜ�B�zfeM�	��	7�4�[��Z9]�eX�:���։B�Xh�m�g4#��h{�6뷳H�5��.
�mϱ�&��њ�*ak��O�
e���S\t�LX�ӝ��S��sd��w�ڦ3�\�V�4,�H�.���u_0�>e��e��ݩ�x�㙳"M�]"�s���,KWT�:d�,����r'�PΣ/k���C��g;T���W��醀lU�YS.��,*�L����� �FNM`+j���ƅRn������8��;1B��S��f��\n�\o����|P)-\�,��諫�0v��:t�$#H����)���K3L#0U�O�V6��x�3��e�� �,ŻƦ��̘�;�u��[�y�D��u��K+l]�wu�8�Ͷ�q\���9it_����E����Iv)X�u1bow>�v{����t�9���XmS���������bu�v����< �ޭt���c��a�K��(&oI�q�"�i.&2�굻z�&)��m��MwC����{L�V�K].���wD>�k��9���ƻ��\�ve,�y���Y	��Ja��;]����y�)��q�u�� ��N��#��a�#�*�]�2����3�v��(���+�;�G̀�sB�f4hV���ʃn&(�t�U������-c�t��j^��GJ����h��H6L��Q���Y{�+����d੾z4�W1'�P��LΌ`̶-ZЕӕ�z�w.!r�.r�r�Y�5��P�9��o��7w���b�R����L֕�('�\0]�։ε��Jv�V��3��k����:���8�u�����=�ΠĎ��ԩ�'{���~�!q����jz5���H�QHO���۝BS�[+E�[� ��у��Pw�(�V�R�	�K��Z����4���>y*բ��`��o�Sl���e�u���;��s��ho�v$�ˬ=�i�����R�|4.wk#��W;8���K�`׃��)s�ȹVG,<��Z�s�u�v�ݐs}��m��vE�+�B�qd�S}i!0��ڭR'}���� `v��
�%�����E����xȰ��F(#�E"#s�{����Q�*�,QDEE핑�%��QQ*��VbP�����DDf%�AE�,�PUX�dQ� �v�6��`,Qb�ږ�JʬgV�Z���¬P�+PAb����iR*ň��X[N�(�[�e���JE��5b$DDU�1�AV*�(*"�QA�DcmH��+�AE*V(��:�A"��gMQP�`�,[e���Pr��
��Q�t�Db��`(*�bUA�Q�EPX�A
�EUTEc�
�J�1Ab�	�Qe(�����"�cZ�r�EQUD1��DU`�*��ŀ��*��QTE�� �����_O��t�F�HM��p<ݲݭ�!����-��i+pꕮt� 5.�^���������py-��ɚ��ί�g��(1"5kgY��f�Ο��ɫ�כ}N/�X�9���зQ'�ryOWt8��j���ֽ���[ܝ���V	�'>��Q����N���nDЧ��P�ڎ�4Z�y��o6�q�2m	ꃊ��4���Q}��IҗOP�jy�}H�)/���}�s��N���Ѡ�J�9.�����&*/�!�oT����x�a�4��T�'��Z-��>�p�u#Cuz]��\v� w@����L��թ=�P����������n(���r5��D���pp}1�?^+����J-N��ޣE$+������j�]���)�����Z�q+dd0�oeoR	����,��̶�z)�ם*I�)�v6�r�p�"[���1�b����I��-�k#�w�H9�{mN�����ڜ���UC7j��gmЪ}r�z`����2�Ԛ�a��ʞ�>�'���j��ouP��B!�W��p�� ;���71`+�x��*Ssc�v��y@�Z�k6�����𫩝f�k�JOw�
g ���6vN.��ԌVr����|l"v٩A;|n ¢�� Ξ���G+5a��!H��]׫�G��G��{� z=��#1��ߪ��������N�.�0ԁ�Hp��j%�ecWV�[�D�Na<��\��wn�ܩsTScn�wZ�k���^���B���Dht}w��H��E����z�R�dJ֦�����䪕�)8튚\S�{i.�byE�M�T]9�]����S�z9u����[\����6���u�~��s�T6^��P]�EҟU�5���Qq���KZ���Ri���X{��J'���;2^����N�{*�^8��5�J.2����i���ڼ1U�8SY+�5Ɋx���g����V�t�련��>�1Y�6{6���)��IR�Y��P��ܫYQ����C�ꋹG*�R���!��ȯ_G!KS�/����ۉ�U�CcOI�Jv30fzVv�L��d���B��Lb�ð�G7��-��z.��󲰮�#�>��]ɑO>#Tڋ�;"��*�Nga�uq���3�����^�}S��oT��㗛�=ᗟ^��dwG9L��ƣٜ��t�N�sXծ��$�O.�ҩ��Uڛ�Jui��w�����y����p"��m`ձ���u��GxEH�P�����yp��������uN�x�B����|J��I���Ӛ�|��:ñZ���6�8/jy9LV����+O5�ι���!9O��\��9���ۺ��S���;���]Pc���Ui=}��o�ʽ绢�ps]��ڝ�-Ӝ���+�>T Ơ����8W7S%��=$�z\�m��w��i��'X������+�U �"���i�y))m�Z�L�����:�ڑi�\����RY*�q(�x���7����|�B��]5:�/�mo7������'��G���A�Q!<�2���{�sO��^��a<�w��Ϫ�-f�S��D�k�ۓ��+t+��1$��1zE���=��z��s�B��L���������6vB߫�_s���������D�.�/v��l�y�|������T�ϓ��!r�?a�\gR��u�0�u��~��7RTu,�M_P�ׅ�^_U���V���#&,_]�Rb��[�R�؄�|��^paʱ���熯v�����]d+z�r��yVΨ�PK���t�id���{Q�Փ:�/{�U������wE�"K��|�����ߺ�(�mc��7�Z1n�ݘ�ª#0J�6�T�uW��y�i��P���5�=��\m'P��sk��r��Pf��3�ٹү U�����)w�n]�k���5yИ�O�K���}�(���}���E�p�#1�gQc׃�tms��_���V�{c��vh������j�uW*��%T����׏J���uѯHT(n�h�S�w�YY����Ů�T�N7u��o�޿�_��\�!����;Ζk&�i1Z�{\� %��le�fF�1+7��>�mO:*D�
$r~�2��|�9��]�S����ॕɫ�MUt;�+�*�V/9 Hɻ����	[C�*��51[�խ�e&������������9`/37pssv��w${.� <'zc�x_�����4=������+;��zo�;욑���}e/?^�K���C�#�\u���0�q��1�5i�lt�2��L]G����L/�'Ѫ������9���s��r������o�^ٗ��wVz���+�a{d�Ϊ2&��^-NI�k[��1��(Z��g���5����t���+���]�mg�g�	���ڋ�;ǧ�/93��y*u�O����u�U��8�=�;}��C*��F����+Vw4�\o�6
�K��7-ԫ�/2WsT*iꮠ�H�3�J�u�}q����O�Cv�\s���]b�+�t��RչSf�ekK	�W#uz��ҷ�L��x|�OW{�k���7�S�z�Rk1���R��,q����U�LSS��Z�^�u�R�.9�
�w��&7��{^\sw��X�M�T�iA��j*�SI�5�/cl�Ȝ�\&m�\��Oy}\��s��(ax_
Pv�x�����I�C��Q�8�J�K�p�y��f�*[Phl����D�׶�r2��M�r��'X�V(O.�1ޗz����l�}]��A^���ڛ~�et6&qT����b��Wk��!7Ʊ2�Cn��7,�Ry���n�&�zV� '�����j�#���G6��rn5&���f��6p��)�vn^IV�ϝwʔ���������yåʼ�V��浽��g6�5l�[���� G�e����v�Ktj$1Ry��
�Na�>�ޮr����|ޯL(N����!q#yW�r��ޥe7��߱-���̶�k{�xˤC�ΔҎ��V��cdA��L\#�z������ݤ][ѩӾeO�$��5��w�RU�j�S�R�A�8LAj�R�}}�u�~��ۺ��B<��I�;&�����_d�M�ź{P�� ��9+E��]x�������Z�7����.���p�lu��,�U+�������v�=͜���ΤI���m�k��͚��M{(����Q�%T�o�Yrx�wZ�|��nw^�S�Od/sҴ��ɾ4��OPŏ��Š��u5�ԁ�uݥ���s��_mCgݫΦrf���+}ʙ{�_7P�ƥ�y[9yMַ�c˹J��v-w����U�=�Ec���>��QyZ�>�rn���Iol�jS쓢�m��Ge��YG���+j.ep%¹�7��/�Z���)��J�N���	Źʶպ���o!�u(���.�-	�mGZWAp��g1��WvV�oE��������y\-�=��5�T+��5k#pJ��Ub]׫�DG�߄z"" �DG����s\�m��/T+_���n;Z�ܬ=6Uz�J�:�V
o#,LUԄt�-�P+o��{������ˍmk��1DU��A�`�G%���	�!�]��W%̕���]�Td_CB�jh�h5n#͹�BF㺚q丫�5�:�-r��FK7.��U�Q�ɍ���ﹾf��g���첤W��ގ��]�F��й���|5*�uT�9!��m�>V�L��A���bԒ��V�k�c��*F��F�Pc�oI�x�YaZy��Ia	�9���z�CW8����ܲ�����>��A�&.�w�7�Yͧ��չ������p2ﬧ����;u�n��\)T#Pb�.���Kn�w<��F��ng'�	�[�Rj˫�	�Zn��u
U ��M��P뛹t����"489{%�f�=�t��~V[br*��m�e�ݶ8��&|T��hX �]�[g�w����Y��Ɲ*iW�\�VdƕД4G$�=�YF:�ww��q�Rt2�ޡX��u3����t�Ƒ}�S��&��'t�h"�* ��u1\![b�����h��u�s�j��-�ur��s�k��� �D{��K�h+���m��*�/\�N����Y�Vk"}͹NTnR<j ������N.�ʏ�9��ݿ�n�P����J���71Wyk{e��dURGc���N��(y'�8�<���=������Ux�;��~�סu���k[���;��Z�8��/�v�lvd�V*�E5Gr��,}�mr�o9\�JG?U�wmt�[X�9���օy�-�{��V`�6�0c��f�&�fyU�<��ut��(�N��ˎmm���r��m��ʭt�)<���;G'�v��j����� 0-��S���:zv2��(���S�i��j��W80n�9n�(��Q�uH�=X�P'��H���+$�����D��Zoanw#3n�u(��ãT�C�aߦ��L�U��j<A��y=
H�b�ɞ*�>�Ҝ�Q��vB�[��d[}K8+��rGW�Q(�.��>�$Bg��1����L��Pښ"l�2NǳG*�xXO��L����?	�rh*�^׆�i�?[ ��؈BPM��_eʔ��l�g7������f�u#��CF���'l��˥�hɷO��YϠ�-�Z���q��Y�D]�bU�Y�3Ämh�1؟ӎ�Na��vO�o\H�r�&��.��*%� Lr��̑<�3D�O��t�l����0è)T¹Jޜ��q�D��*95yG!�N�:���A��ZZ�Y!���� �R`8JNQ,4n&[�a2�^�H4r]����˳!ծR�����G��vX�sK쉇�$��$"jT��⩎���^*#��H�7�O,R�\�����ܖ{��������ڃ�]�)_]ba�=��ҧ���3��za��U<&�^\�ϻQ?N:�<�o�x�pؕ�Y�3TȄ3���ʍ�xj$�yq�كzm>UU*wVin�r�ή-)B.��Ě��p$Pl��ĭ&�XڃBCY��X���uh���mg.Df�n慡ߊp���8�5���z��b1;D�e7Lh��� �;�vF���`/{�;=䠹
�ze\\K�<�map2Έ��Tm��M��G��Y&_O�^�e�0�i�m��͛�~�-蕇	�g��_�σ�����F5��I
��]���0r5�0��N0�t��2�V�WE`�C�Hp����l�M�JU�^�e�YJa�CX��{���U�GWl�B��4|��Y�4�3�m&���<�gr��̸�f"u�d���)q�+u9�cBj�Y�������F,J�!>;�љ[� 5H�u��:�s��o)�R��������W,ߣ�;�;tb�,�aD�7'DPB0�U(�,(4&LPOnܸ���)��n���uu�Y�v���6�������4�>U����.㶥��u>H׸$�_�bXF��S��.b���86���뛯�P����9��������~�ϻ�$Lh��1��D�!��h�(,(2�xŭ�ݑ���O�Y�0�R�ge��bv�(+U!�,c7�০D��HB�xzI��Q���Y�Ww�1���Z6��r�Q�:���c�P<7Q|���K�xb໭Ñ#��Ub�1Z ��Es��YJ��qf C�T`Li�Y5��A(=��).����Ku�f��E�U$�k�j��K���;zlh�N�d<�f���0��ry����C�:��:⮭S#�k���@����n��X]� 9�tc,V�p卯;��
 A�Rx�+K���z����Z��Sj�Pq����'%���q"�9�a`uJ�%��,mC��°H}e������Cs��y[Kk;N`�X��'�$�޵𥽛q�N��YV衜��ݨe���W��ؙ���ͧ�Wk}8�������\ ���q�,Nv_s�£eP��� �e�J������YH��(��y�::\�af�؊�Ԛ��
^Sz�Mid��uخ�3�)���CuQ"��+˭������>w�;�|D<��KT��	S*d���v���U�����3J�얎a U��H۾A<EDY��ڽө�����;G�Ⱦh�& !Z�QXMz�R����w#���>��p���_JJ�t!��g�R��ՠ�z����`j��`��pǽ�Wue=�jf8����[�叹��#v{�<�Wt��,K���Ɯ�b[h�g�(J���
�y�LJN��A� ���ۅf���)4r�c�Vnb��72s�U-;B��II�si��ɌV��9��k��f�����'~�cN��������b����8\��[T2��}@���L	]�pc�B��"�V���Sw�zE3�����;.k��^-�s�U�ot�:��� �7Vvue3����i�/�qv���= �F��5�n��Z7_llG��1��e��t:p�`�� �rdC{���|�Y�����x0+S�(pǠ����X��G9#��s��玲��D�Q8��� nNT�>1�sEk�K������v��GRG�4a�ұa\�0a�0�ͅZ5*.��⋗C��'30���ST�2���;G`�7�8,t{��[4�*�%1إ4�� ��C��鞾����c�<m�۹��yG��Χ�O�[]V���b���p:������]].�ba��6xu�%l]�L$
%��%�W��������)&h�fr;�(���+:�\�=$^�ؾ�������3�����o/����W��3��[]7���[�f�G�'%�iZPך��������հr��X��f��p���G{�ڍl�+�ja�f��vZ���KT��qZ��;�wq�u��uܬ{x[z�k[��)�z(�l�yK	�Z�H]��^�Ԧ��I�h�{WLq�Z�@\_ʳ��{)3C*���8 ��71�K�dmj�fx�AM��!�WI�ڭ�v�L�su�I�,�Ҭ���l7�5�έrTٷ�Aryi������[4���
��]+�S��Ʊ��i8��a��V���[�¯.:�jfS:�}�zV�\jH���-6��5>���Lú:*'�����:��,�t 
c�$k�pU��.�q�^�!��d���:�VX���a^Vh�p^h�'���Zy#R�!#��hU�󳋥vuJ�+��f����	1u�U�(r8.ǇK�w^�ψ�� 6'-�jƳ���Zv+�2���wІ^v�-.j�3oV��b���R�0�3��'3�}aQ�[�A���%

�UOBũZ�&�t���4^*�F�q��x����}�{9���V�X,QՅH�D`e�R(�
�ڢ�)
���b�ɫ���f�jJ��,b,X頊�H��cőV"����UEY����4�Q��uh�2X�"��
��TKh�U�dYX(�X"h�Q`�c��Ƃ�b��QV
(#b*���b 届�k�-T���E�EFՎQaU�2�,��Q�"
1FLe@EQ+V���B�ETe���-Ҫ"V�m���2�J�Kl�h��b�-�1TY�Ze�X+Z
��q��
Z[lU+��m���Tis1r��³*���&[ET���
��R��̈�H�P��#�l��m�U�s
+R��1,F���[Q[���8�c�2�UR���+T8W��������+[�#L����Fu�Ԣ|�µ��k4ƶ����esXf��kf��j`�D����^J�z��t����u�6�V!  ����/��'|P��
���ר������Ӽk�}(D�Bwj�$!��S<���,���sS�TX�e�2�ͽ�6�N�-鎢��:�m'Q�TtO�8�e�i㠣�t��_�Zj#oi��8}9U��N���N[�<2���"�VtK�Yf��`�1��%��p�R F�[�\L��?<`{��`��נ�L�!�\��i�-B�3l�1.lv�iD�����]hW
X��ֵd\=n��65ZC�ބ�JK|jE�X|�{�7%��T�e:����7u;�#�8����p8on#n�w�T���,-�9�}_��U�`̓�Z����Le��֕�y���M_D��DW�EO�=�T��E�£J�uQ��o�i��z9O$w�=��l줰>1%��?09���b���j}0�)�<4�6��� '9��u��#�c!q���Y8K�Ge�A����Me*l�qݕN>�xf�So�*^=�9K�����)���L6l\k�\mؘ�2#@J�g��~0P}�T�ȹSӾ�m���+׸���������.hǗ�G,��$���ovuEDV�ɑV�
�T)K�Y��岸��*�7�H��F���LUr�J��2un�M��Y�f�8*9e	˸�������㜦=V��`���xu��j�Q�nf�����k9�1��"�$@�%��6ֳ�v���'Z��]գ���,42r�Ryܐ�Q�8C�>'�똘�ڛWO����s�9'pѩ� %������R�(�8��ѯ_�yH[��v$	�r@1+��^���<�$�2\��j-#P��04�J����8b��'.��,h�w�~��*��euf�g��CHq� �.��Z��\S�/î���2}��	�XT`�����}��0��kUh��ê������
ꐸܒL�$,6�O�����V��h-�RJ1=��58e&�-��К;�[۰%$F@u����7]6ٳ�mY/*�+�x'K:��7��$�X�������L����k� SyH|X��\�;�e0�ұ1��L�?��K��"l����޵Ӯg)L���\힌(hk����Z�-�	�~���j��5J�z��d`�ND�G�ti�n�V^o8��VMa��]wg�笸ژ�zu:/�]"m�ֲx����B�x�����]�mO.�e8�ZdK��r�s��P�|�W�cu�<��f�l�6�����p��*N�qDggl){��d^�>n_\���u�bv�ʝ�Cس6VeX�U�8�5qs�
S�Ԁ���ס�˵���l�|;h�:�o5�u��ݕ�1���9�έ�@�=O���wx�T�]��\���R�5; ]C%�N9�w��d � C�:��o��z�������W3��,�4����T W����o�׷o*8�ES�N�{t��5�*�)L���V
\]#l��VqR�WAL����;X"�Ę;Y���Dfb�����7�)���:i�
�>�z�U�)��(�>W>9"�b�=뼒�	�-��_{���.��Xs��%#~�rE�û#�AB\
�%Pr22�F ��]Э��\V��M�R��
;�k�"b��ąE�ͷ<)��8S� L���T���y[6p� �����z�ĥoNAs�8�����W�s�%���wg���1�q�Zi3�)lu�0'�s$���1�j�7�T�G%�`P�"�TA��JR��ow�a\���rr*��n }���J�L���Px�RGQ���w�n�؀ڔ��w�5?X��X���r���|xR�J�Z$ԯp[f.Z<�~ƴ�����M�T�g%j'z_wT�PS,+�4�ؕ�b�L�B��	�yK�Z<%�N�/	�q�)��=�K���o�1R�܆�>':����b�𭜦��$��̏�p�*ۧ�4�Ue�i�ݲLН������s�W_�ޙ��j�7L�仛M��X3b(3t�9�b)���w��q}�k3|kt�H�LZ��w�����W�QI���vu�4�`u���x<*`�'��͊
�"�?W��m��;9�ފ��]�ʯM?T��7r�檴��|���\�b{�L:(aަ4�$5z'�-�V�Wr���(�-�^�U\\���ٶ�P���>n*5k�N.g+c�@prnH��Ε�\�&s���V�[1�p���m+�\�r�����㮐uZ��^ ō�z�������-�w�vΌ�tYuVx���M�e��)�/��n�j���[��R3�ڞ�;����ߝfΏo�2<w�g��4ϕi4Rkcy�͊�h�������Vq����^�)u��63�]!֫,�/Ǆ���K���X��o4�<��Ӊ3C�_��&G���!��������*w�\-�!ݑ��۷`G�cj��㭓ˆ�e��+��L�L�⺨A�OR@�-��"Vmuܯ���&y�t�j�$����VT�aWTmQ�>ޒT�3q0Pu��<����.��9#��![�ga0P�Hݭ���'0�yv����Bk����v�/w���8N����8i{o���\���䮛�5l�r���Y[wR๕��wP�է�t�|/���:��sR��k1��t���� n]gI[�di����l��k6��J�T�+^����sk⑪�����s��tx@b �ZL�wz5��a����Fl�*"����Q�>�ĲO�bPu}JK�t�j?�/�}Js�Ǚ��{�K7Xޞ��~�Ɗ��h�yN��\S�
Bx�G|u��kɒ�>MW-�/�ڗ6$|=��<cR�iAwl|��l���3�w�����`x0��u�I6�=k�3�	��S��������,��+���0�:��(l[�6��Pc""^V��5�Ƕ��߳�lM��c�*���@챹Y��4��:���*���z�x��ҷ���˛om_���l�G�L������t�E�;��:c��q�뉸I�D�Қn b��w�jw�g�Ot\�ݫ�UA�m2���<�)1Z=�Q;yV�{4��*��D�;�/���Sbz�����}wu�KT�ci�����rV��u*�"�`P���{�4�1�P+o��PWJ�H;�(7Z�'��:�6ͅ���Bc��o��)R���<��:���R����enʳpk,�m�L�881�T=t�h�U��Dl8\�+�a��Ǳ���kV��;>Lu�:o�R멥�����P~6Mr�ǻ�خ7����{h�q`,�V�q���3��WI]N���WpV��=�7��߆Ը7�A	x�I\�F�.���ܣ�A���Stj��q\�Z���@L���v���h���Vϥ%��\�*OiW�9�q�)W�4����]=9��'+-�ÔB��\�o=�|��a�ͣ��X��� �K Z 6
�Q��aVmd��w@��1Y]���c��W�EG�ؤc����	�T��L�SΨNĪl�z��q@\<��q�[�Q*�$<�V�g��F��k�\o��Lu�`�%@�'QwJ��s_B��*ºm7+�����}�v�:"�jw���,43���,*5�^�T��	�y��X�n�ɦ�-os�:{��e�Tq,U�O�D��LX��Mfh�x���g�LW� |Ϳ�ھ/ӹ֩�Y��Q\t��/����Qz�C�FL.�+����0���7��;��Qo5��{������cՐ"�<KKµB�we�u�2��L Y�O3*B�x��'=t���(}�'9#ga�Lv�����NCh��*���Mc�Ll9_٬��3|�26�Yٵ��Jҝ�K5�W��,K�۵BV�"����.�7]6ٳ�hz^U.s��k��۰��;��'��T�n݁��Sג�j�B��ۊ%7Efw|�um�^���xv!.�{ds�����ܸ����č�R�W��B����l1"�a�{�����q]�S=;P��W�4:ģ�j��9��V����}`�+�-[�Y͵�� � 1
�j����+V���*�W:v�D
�����침w��8am�-K�ή0��=g;���FB�T�0/��G�PCC���HZ��g�o�d���r��0]����oI�?L�j�*�L\b�c#nU�u��n�E��H^o}r
V�e����z�gf�����L��Ms8���M��ڊ��OqqU	��b�Cea�)M�ù{��b�qOe{87���{���Cn���t�Ғ��e.X���}�2������Z�4Pr-�0�9�]7x%=oH��a��5�ԖxF��jNQWgC��P&+�S$h�ʼ����MB��QX�q�DD��뇈�aи�;���L�U����κ<�'�n���v�rR2���KMQH=��C�1���o�a����w$u:�8T%����|./��a��'Vp�q��������D�oNa��#]�Kz�B�����B��+VG�왮�''��Rp����L"�<!������*��]� .<�L�.�J�Á���s8��F���#���A*�lqw=�-<��5��{�����^�U��^�����Xt����U��ۇ%��+���/�[���s��햰ht8˓v���I*��J�:�L�q9��w
��"Q��;������ DG�չ���`�������C��r`O),���9��Wq�VP��y�U���.������S�Iio>�ia�ť*�H�W.���L%RI�RB$�­��:�:��W�TGY-�oN�c���לfY��6�.����Q�
�aTu�&'�	�7�R�~����R�ӄ�oˤ3��额�ޒ�s\�=�¿9�@�6%i�S"��&�vq���ځ]K]զ��)
�R���l�r�"�y�I���H��Pa<X�hH`_.e�{]�-').O	�HQ�~��.⧆i�,U�evOY����8�\�q:D�e(ݧڬ�GRx�ͽ�4]\�Xu�f�X([7E��ݰ����:�����i�|5������f=�|��� &�p��k���5�~�i�V����������'t$uqSEJ�P�N�4����H�z�����+Ю�5Q4�"r �f*�45���\���2��D�m��;������n��\�w7D1I	�f�v�d��;����E�mm0m\};J����9t�,�<w	�e($�#��<�*;u�r� �5͡z褴�h�f+M��\��.r�a�v<���;��y�]��l�eq��C��2��Gwe������{6�(a�y�)"�u9���fsy�ݾ�w������G�v�?�%vh1��"c�A�Q������:�������Q�r!��P8DŠ�?e��;;�3�4n�~�T]�I�b���D�!����Ce�b�
��A��,�;�rkZ����Dhp�N
��s��
�I.�=lQk_p.Wǅ�|Z$w�oZ���hk�#Q2��@��nӮ�u��4o"6�:;��&
���y.����F8�ybӥ�h�CQ��z�U)l�c��"%2`Ti�Y'�f%}*K� �MOK��睩�H����κ��%��9�����]��ظ��`@�@�7'����k���	Ř���ٲ%�WIb����CYݰ���#�f��X�R�h�N�$ֶ�us�<����=W�B}{����w�\HL�8ub���Ö4C��y��6���A��ŏVXD*����E�����,R��q$�r�MBwjS��c�#���#����M~��+��d�y��*ab����	s��U��J�� u��s�ڦ�ڒ�i��>���Sg�s]�����H��k���pE�;������-�`��I]��5ሻ<���n�9t�fm��S�,�(�9դ�̗3���%�X��'�����K}�G�^��j��}��a�Z��-]ֻ������ed<��Y��踟����~���_���x�#�e&+Ge^\ЃWM�ufOpʣ�4�<�n.V���)�
�s�� �o+��;����\F����n�]F�ʵ��[}������$����������
�G�~0}��d[ٌ�Ō�ʐ��p�n�v�#�q�fg�[��Z���X)<���5�{t��UNΌ�E��޺b7"��ƭeDN�d��s�����7�hq;&�� ��LMtL({!oʼ��N�����1�j�Ke���^7u'�ݥt�����ؖ�RKG�?0�W����l�g,��P�mZ=�P6X�gA��_�jᗴ�����uIP¾�l�qxt��Z:|��?x�)�cy}؈Ma.��9Һ�rD�R{|+<�6/��tT:PdF 4��ngYw3��NN���$
�]4d9�]��b3[�Qok���9^�£N�S&L�o5��N=8�u\�˨���*zC���,F��n�.7�*�y@1"�w3���{�u#}7����brz��(8YUJ8rWm��C�>Oi�ͥL���t5w&BR���q#�෵���]�����E����Jn��[�U�g[+.Hh��t0�R�u�d�v���Pkݎ|1i'���c��%���àm��QmdASwa5-�e�`S��y7�p��9w�q�MZ.BՋ�����"��J���E�#�4��#m�M��.�ms(սȕ���֔*Y=Vr�{-�
�k�������Z�ZR���F�u��k9MS#�6:N�P�OI�{cqsM�,n�^S����8Wwdx"U�ҳ{c�ܓ�kI�7#�4�gn|��4]g\�qQg��c��>��ڣ`�T�!+�����A�w]S�Y(=�����% B6�7����;��7`���u(�x/�wr�o_�96�����wjgz�+��;`���M�f�[�����10�Db7�:aQ͹�f��.���zf�)�8kz�G�Fc��7C�a����E�۰����us:^=������mA]וc�^ά�n܎�
j��V���v�b�k2�Ir�� ���7w�o^� ��uo�g7����ZWu���u�,���n�>Ǜ��T�b}��Ss���s�9�7�\�Q�N�X�l��޸�����Kpŷ@L��tV�\;����R�aΘ~6�̝����k��)(���yh�]B�V:5 %�;� z�Ƴ����;3�]8�y��X��b����'^WZ�9�o0�WoH��u��~�#�2&G3��<�n<\��suۚ�ZK���@�SP�s��}�y��!P�w���:��Ԑ������@�u�ʜ�XܧB�osf��_(I�+�+
�r2�Q�dz�Dm�Z��F�
<�(�88�[W��=�^#/.�y�Ճ<�0V2�D�����{�}�x��9����:�H�% �WS���6��,�p�
ޫ�+n��K�� ��ՁwH�"FS�Q��ޛ9��VN���Y�z�U��}+���pt,��r�Ob�� ĩM楦����:R]����W{VYN��o�7U͢��;��c(��j��K������7�C�@�)�j�4�<O7�lx�whan��#%����:��9e�G�vz�޽�0���2�I�*���p7[u��L`���+�e���uχPT%�:9>�t���KC���	�-�*q-
ʾM�˷a�q}�u�dU�j��yG|�9lA�;I�:�g��
 Z�1R�l�9�ED��-���'Z��w�;;�v��ȗW���Q�r���ciV�� �옻��8�`7	TV�Q�H��jU�w�R��i-�/U1qg��՝ի`�^M�^˰�1�ժ�I��j$Y7���۱R�WK��k�G�lMಭSzFX5K��]��r�������������\��Dj�&�_cI���Wl����|b��Q�kn��ǠD << �0`�b��E����"��������"���TQm�f`�����N�J���ְTKj�(�E����S3�D���\��1�,c�Ub�+{����R*�*�����b�kUA�Qf�Ub[��a��+q��J�DX5*-�`�b[G����#�F,YmU�B���D����DT�"+�J5��Eb1r«2����\kA`��*�Pb5�+X*�2�3�c���qF.4QkU�n3&!\@��-PX��0F#
��)��j
9km
��Q`(�e�841	X6�l��\���d�H�[AD��"��
�r�*"�c-ĬE�T���-VcY�88ʈ���Z�ڱR�J̶,�������KKZ9q+q�+d�)P�֋2��J!����S
��"
�G��o�ޗ�k�w��עwPB�LY�A<۾p����/E���$Ρ���_ut�s�!��G�rD��Tz�:��{:w��U.���������7�c}���UZ&߽�)���fatFLhu��Y�ᅐ�a�w��4���c�	���˚�TW�v�cj
6đ)�D�ϴ�­�ajTQ��L �t��yz�X�������ғG"�a�+�*!\�[$+%�=;�<Û�<�#[8vا�
]'YyRK�:�UJd���4���e�@tr%�^_T!���zo:�5�rr�e)�t�oyԃ^\�	�S*� �,]D+��}�p¾�L�t��fᕉ.@f�Ɏ���y?���vOY�1���C���������A�����ꖴ�T�9�e�x*2�u���s�Tdm�k6:)k�M��C���=���̇���y�Wn�H+*���&X�j-����)�6f=
��?Ż� f�u��Ý��@o��޹�٨�aKh�=�,�`=���μ �Apr[�����7�2vAر:��=��a�za�M�g� �ȓ�E�N;�W�3���Y!4du��J�������^����uDg=K[;6��]���nl�أ�2�ռ�nI39WL�/��[��EDHb��}Pf�J\��NT�"�Xk�"�\]�0k��V��Qj�4�mM<��^�u���Y��=��#�z"=��;��G�u�l�G�ؖ��{^��o�#+���_w,Q�:``0��=���8�f�/2�j&�aQ�;\qx"kKsϬ�V�5����q)�rGS�#��3��^e�'����E�[ 2P� U鷛%#�|7=w��R�ٲ��s�b�{:�>9�ՙGe��ؙ�S3���F�@~�%@��4uAͩ�<����Ұ�&���b/ �'��s��[Z��b��N:���d�J���r�ɯL�ѹ��9�����J�"z�N88�{����oq��U�h��nӮ�1ܻ1}�0�Ю���$"J,-u�뚦Ё�}��x(}���i�"�0Ƴ�ܻ�T�㘑�B���tI��C��G�����]�q��yyM��}��cጷsy�G����i/͉ZE�Y�6�1�ox�XU�	�KV+�;4���W�g������w��~��q&��(6T
lJ�n:X٣N�@��7}��hb�Ԇ��tK>��9������1��i=�TM{�+wU�+��+�Yذ*�Hʙ:Vf\�w���t��� �~}��x$���:Χ5�׹�V�&OU�=q�v�b
N��c}�tq�h���':�oj�WS�������[�Z��,��-�vm'VVq��i�C
�f53���NVww.\�G���芻�ږ}_։���Z�`ǋFP��D�:|W�/$��V�c�&y`�/���%\���M��#��z�����V��
����0y�>���������\|�7x�D�jT9���RuB3��'����p��8���Ί�;��/'��n���x�B�Zk:�YA��;��݋�1�b�[�*烿M�R�,�[/������\��Aa�\�鸘�}=H^tJ�>UO���f��Ӄme!�B�z�*��)���GX�~���Lƈ�q1��Y5�C-��
��0).w�:����X�ΜAÜ��B��:��vK"���ٸ��u�B	��`p�^���E��T(_B��f*}��v���.��qP�T:J��ޒW�	��|��Fq�=����^�Z7�ꙵ�n+. o�M^
ȋt�ɸf:�"%2`W��,~�Tø��>�u8}}�Um>U&�VL���#8�K�~�N�CNh`��S��B�T��3�d��u�B�J>}���O�t�թ���H�N�ye�� ��-}w1� |�|[W)�q�0�H&.���8�R�"�Ǻ������_m���M��+5'e���s'd/�^���	d�K/�=�ߑV����Z��� {�8�8����Jt����n��.1���CY��\@R�с�ZE��1�0�x1tT��5����.M�Q%#�3V�T7%֪$w�9�a`uH[bP�$_+�;Ew��U���F�������H���˅����^�7ґ=�*qN
5i�X���/k���@�%p��d�|@���.x+�w�o�c���^���B���{�D�u&[�T���g��
nq'=�魹aQ4^t�i���/�qM��O<�U3��)gU�2:cC�\�q���Qo+��;����_�@l�I�7g�!�O/*���/�����hxkM6�콤g]hw�,P�u]��G�ԇ<lk�����^T��ڜ�w�7�����+��V\u�O)-�cF���Ъ�����r�dv�a���z�%��Ie��ل؝�h+����e�&�LMlL({#�6�ɚ�T��k�	���S���t�R�E�y)1Z+Ω0�VZ>=),����J~`/�� �p>*!�Q���5ps�"6��j�����{ëb�Un�͋eM����T�P��K��<�(i6�"��\����+7�;HTn9��2Ū�Zz�8w��'p⠫�D������xO+�<���� �S«��b��R��K��w����z*�79}��#e�S��~���q���f	�XXPA��W;�!^V(;KjnH���Z�w�e�f;
�F�)-��a�b��t97<dF	'I���=�~�2����$~S��0E��Ԧ񡀷/w,E�kw�y	�+�a�'�ܑ*d��j\f��X�����D���*�_�&7�=u�ZT��yQ��*���MnFyۧ��!�!s�hߴ)�h�_J���G�tlH�  `C����f���+�dƇ�T4�]^Y��+��T�e�;�]kZf�wa��(hU�v$�nJ$TI��>�&�ag*(���b�ۤ[�l����ʼ:�#_�S�ģ+9Wau�p�I>�#��墓[Q06�2���V)��ws��V4��ՇO�%Ҟe�wU�$E��^WU]>�dp�d�ӆ�Y�1�jRKFr䱷2r؋*��&0v�f��H4��P� T7(���sP�;(��0���<��ͿgK��@���:�*��x���۝��B�p$R֬�g�x��W_\w�^��.IM]�Vzי��f۾G�|�]�}��n��̰T'J����z5��׻<�Z�G�Z���)����D���eh]�6��ܺ�3��L[k�D�d��I]�7�֬�\�V��3\���7M�k�
�Q+b�{��r��{��x�z#�q.�W�P�8ҿ䣎��F�3��[F2k�S3�TdF�F�~�\�^Z겐�ͻ��}�Ʈ�j}3pZ��ުU���d��Dx�|���Ip�]O/9z��墜Z��ˮJhP���;o����+�E�<���z/f0H�(q��l6n%N�Qj����l��軋gr`���I[ˣ@�PV��Ä�aPc���f����R�ꑶ}>��x�������I��F��zH���7k��T>FV�zW���3�(��B�"`Ɗ�#���p�vW�EV��AK��\/�o4z���Ǹo��d���~���\���ܞ]dppM��'Dux�Ƣ+U�M����q����P�P�{"�#����^�O�U��~�RW+�A���t����Db����Ss�ބ=���),���V��z0ӓG��p��I[��Ã���|KK���T>���hK�������>s�Gχ#y��]`���a�n]��~�r��<��P�!V�#�k��9M�i�D�Z�H��Lґ����^C���U�B��Ög���y����m�:4��4�'ΓX�a�Jtv�@���{1�����ȯ�)o�]���{˥E��>��}�Uڼf��y
��P͹η��zPܙ{��e&�H̜q���wz�a]ѳt���v�]߽�G���=9������F
?�$��q#�ܻ�x:�Cq�H��*�aW]b|О	���t��^��#9�T�U�b�ޘc8�sy�C��a\�"�bV�=\H�K�t8�Ѯ���ǉro�"߶'0ԞJS1V�o�R�]�y�I�[lH��P (z��]�]�G�sЎm�ᷗYP�k��Y�Mx^Uqpu.��q�j��L}�յ�J^d�t,S��l����r�c:,��bݮ�T��'�Hc9E
�ʦ�ʠ�sƢb�m\�[����ԟw;�}$��c��<���W�-7yL\i�avL�I���!�Lkk�Y�*��(��%�n�$F{���'T#/�4\=n��ŝ
��^���H۬��8)o��-6�P�����y�X�@�:&�n�w
���c��D6�t��5$08s��(d^Y�:��K\J��q?�,��S�P"�z|3����Ї�e�a1x_�N"J�{z�7(�v��=���Q�``:=��t���D�׎�d�b��{$0�� ��tT*���v��:xZW+(3�f���`L����޴��c0�r�CS=�ީ����z1Z�_RZ��`�r��}T�Z[�;�Y*<����g�Z�Z���YrDGvʿ�kv9��e�inVN�q�(�0�+�P�]6K�b̛���[������DDL��9}�}����a��rr��
��Q��L�x<ˠj��\��� }�xǎ��K7���!�wk��ƛ���И��Fi#����3�F��\���^�՞*�'z�2+wLu�q�u�s�3¢�W���'���5�@�0��	�<K�0�T�����כ����A�?E�t�x��r%͎�Jw�sCt[w|+"U����U���f�
N�k���գ�^0���e���RX�Dc��+R�k ����R�ѐ5�2�U·wF�*��{��]�8 �D�nKeU���ݦ�7%�֮$&i�]��ذ�=ǫ�d�]�A�Cll>�^�Z�$L����"�<�:�0�٫��Vo�"Mn�obdkr{8��]g�'��Ӱpf��ׁ�7�+�>��
�]
b'���K�K
�W����K�{I&L�Q�x8IP�TM'Q�)��t��/Mm�
���3M:5ʥ�[�7Wbe�IL�/1��z�kk���ΫdgLhu��Qe�"��TvWƲ���������$�n���{P^cf2h�.Q
���lm,�I]S�0^�y�CA��h��Ņ����D@��V-♷�3��J��8)�Ρ��j�\�.�"�t�v��gu�Z5E�A]|�� �� �bޅ�	rﴍ��}�߷�W�P��I/�ϪO,�4ra�k�xp�,\e�0�#��;R���"��F�ȆpV�9�x�(͘U�V>��\����g���~��QP�MtU(8o��ۤ��gB,5C^��j�w��.b�9�w�u��pu�>Kw2�N&'ձ0�T^��ʟ&s*B�0d�jz��:����ɼ���],��h�(*u����qĖ�/ -��MR��w�:���(��D@ޓ��O��<6�EC�p+�uL�����ps�rZ?mF6߮�	2q���Hz����Ko�d)���ppk�1�.���`J��%�鞥�C�� �#�Xun��9xz�b0f�QV���U�8�7��
yh�\�Bt�c��H�|��.�"�O�Ke�D��*�����/AyQ��T`���ddC�K��ڕ�����sڜ,��,k���� 0#Gmx��3z��茘��5+����0��=j�#��`����kOlg	J���a��X�v$�nJ&�3�%|+As��wr<Z���ܞG���E��Ÿ��eך�~;��>�p�U��4�Tkv�����*�<6rS>K`U�������\MY��M41^�̅�}J`Ȓ��Om��;v��.3�nwm>՚;��Og7�x�9�[�0e�a�wli�B�'����L�������߇��.�|���}Z��ѻn��UF���Ȱ���W(R�$�rB�Y��;^Z�)����Q��31��=Y��g:�i�N�@����ªf{��B��%`�w����M�6��)�SՎ�'�Ucp�4���:�^D
nP���:G1�9;�*f�߽<�������~����E<��hTZ���K���KZ�.���Q:7��*C��0�e��Xv��G��d`��A�\�1Q}�p�F����f�:#jk�=}hS�x�rְ<����~��;�`��p���(�q�ٔ4�e��B���b���]�k>�gen(�D�#��y'�gx���xe����+��KL�<�ʝ�� ��:�v�j��u('�=}(��P��Pw
�\<��-8c��=u�>,V
ZZ6�������~)���F���/�=}J'�"��[&��zy��y�eaў\%�w,T������Z.o�ƥf��B��$�'q[laM�,<o��V�5\7Ը�s�H��U��?�O�ʮ�]E�SyVlz�6�դZR�2��]sD={�%�Ae<�	ػ��7\6*.T�U	c8p�˭�$"�5��[��7���o���7_<�r^�YH3o�1� ��ʼ���_�j�0�ꏍ�����Z�]m?�sټ2�����w=��sip���Ǘ�p=���JT�T�����]�q��}	�\3���B>Q��x�-t�m.��Jyզ$���x+�Y���x�����f��t.��GOj+�@F)�Ҧ�Џ^��8M"��V /t�,8c��Q������e�b��B�T�ځ��5H�
�|�V=Wͅ�N�В2��4m�Pw�Z�s�o�+���sN<�^9���B�dd�{W��6;7,�D��K�;M�ʏ[L�{+T�׼V�A��LY��W_m�wp�[�)p4U����Dq8-�H�Ln`��NqJ�b��Zl�h��nv�JW	/Uؕ�7RyW{{x��5�츯Hp5y*A�X�%Eu���Cv�-�o�{|:;�㔺�e��M��m�5��6-��=�y/_wD	=�ךwz�fT��mX�\��|E�j��6�4GY�K�VX�FZ`9��q'���l���&�C��hWb�f��'����r��o> m��Ok�S�/7�.��1ӻ�
�a�!��en���I�j��θ��+���e&:e5�z��i&����YT�V�f�,�t.�Zfs�j����"^Lu�H���u���x���e=������J��P�ý:=F����&���l�
��x��2�I���aGm3g��v���mun�#��Y ���Gzi���9y���J��6u(
���c��R3{��a�-����LR[&;�;br6o7�r�,*U��Z�*�'�� �3��A�ṋ{�L]aVΰD,���Ƙ���Am/�V��s�ݨ�����R��h_�x޷�A*��5%s��N�V��=%n!�P�����9�Yr��h;dV�^���Q��Э����P��X��|S�Su���U�;��������[a�ޭ�k68$�A��X���p��
]oI�M�m�uk�C���R��;��l���f�-r�tw��L�!J\C�	��
�\*m��bL1f��gie*�J���8���p]���=.��4.��\�u�����st�O�����5VE���RXvQ�ڦd����s��s�;�k$,;�:i���[E;�Y�g��Hl�B�U_u�)��zܧ��۱VX!����np�.R�w]֑y��Y�Yj��h�rc�\
:/3*�eA�z�g6�g�lfmbʑ��Ɠ�\�۲iA����[/9��.�R�{z�oa�T��x]_.ޛ���Q��-�vt������,[�}��q�j�3�0�]�9E�+%.$�����������W*(bk+R��Q*�Cr°+X,�����p�,���B�+2ب�
����
�J���IU1��YSo}��p��b���\jZ��X*���#��P��j"���b
j-E�U1(��+�eH��X(�LqP�LTTH��j�j���X�
a�QJ�dU�$���+P�6���3,�V[k��c
��H�6��UB��B���1�p`VVB�1k
2cdɕb�LV��J��kKAe���@��q�U�R��\�f[��fJșk"ʗUCi�c��br�R[��2�J��q�s3IPq1�k�VbUk1+d�E��q��@���آ�X���X,aPīi��0E����[ejUb�2��j,���LC-*UH�1r�H 	H� @`o��D��+׹���Z�g}�|�B��>?wp-�e��
s1R���X�7:t�nt5zz���Q'�]���yG����Do�˺�������7�H���@�'D*�"7�V���-��+=y�m>͔�%BgSi6�.oyD��Տn�Z��p����+΄�ȖF@0Ĺ��
��T�)S��ʹc�27Fž�wJ�����1^�G�ٺ�^��V�:�dЛ���Ip�YCቍ��o�r��=9<��&P�:�v��K������vbE��f��&G������aUL����*:E&��b�^x����	W�;��+�T��Č�P�*�aW���Ow=�{�n�Qg�C�8̱��za������!��
�9�@l�w���z:�d�mTwt�o8OI]�#��&6�'�פ����TZͼgyJ{΢O-�$W�e@�`i����+es]S|��q���'չOF��Hf���Y��k�鼹B��3��=f/S��v�CQ��
��Dd�cQ�YY�l�}|G[�׭�ݖ7��^��BݙC���B��n�ep�2Z�;�K�5=�tt�:"�ܜTm�v��{:����[yL\i��a�-�����nB���J�5	NFB���7�`}�1v9�����e�ipa�.���޵�������euJA��-��ۙҍ����걧#:���n�NP�ǜ�/��Ok6i�-�n�䬦�v*�s�)��pTjj���n���گQ�{گ�~�G���D,�֟�_N�����"��G"3���uB2��@Žn����*��QeL��ܢ9�}��z���-颐�\R�甴z��:&��H;�N�_9����n���us��S�S�S����"G@:\��vcI�.'a��PEN�*�ŌR�3L�4Ocnj5�n�G/�z[����#C8�����U`���U��Mb�˿=��˙@��ʵ�$���G=-��Z&\;��J��J"ʙ�u�BDN�p6�AG��C51��/���I�]JM� �����B*<¬�Z��`��J�`�թ�'yt&�K�)b�\
�EPc(Ï)�xrG�E��e�B�'a<�U�<K���uT���I�wE?LK�Ӓ����sc�ubsC�n�g�U
;6é����-�o)��6��\���WK�Ìrx�F�P�Awq��t`l֑�:.�v_h�ס�W�`ݩ��'A�I�]_��ݖ�7%�֮$Rsl�A�j4����6��X41���������ֺ�p_�Ηm'7�u4챎������3.����@���L�ڎ��AN�Β��4�&9+6u�!�1t:V���(��R��)���Γ�,/��{H6�G]��ؤ�B�{���~��{�����,ϭS�᝕�X?.���K�d1��0=�f$�rj5��9��徲��_Y�x�D�8�`���S\��nJ;q
X�N�)�d�{�^�B����-��(���g�+w��o�>O�:����&'a:���9�t���mS9��G�T�LQ��X����z������&����,lvu[##�4:\����W��)h8���ه���R?��*����-<�E�K�g�4o��1�d����Ì��ԱCE�jȞ�Wdj&'X'>��Z��|DM!��ce%��^ue�\)<�����<}�p�%�l��F�j�l�3ov>R.�8�{_�eӎ�u�/[�1ҩ,g�� ��ElL(�qdU�Pu���[�{���|mZ��V��EK�7Z+�&n�'��3<Ӡ#p��ȥ�κ1��	�� ��ml�h7����Q0���q���f%����6�W��Zm���w�:�v$�L�ѮaᷲB}�4;�^��=K��
��P�z�ɏs�nk�4K���{��ޟ)ܥӂ���c\����\U��v�r�vFr�m+���V]�TW��,o����y�`#������q�l���Ra�Q}]��֢������]ʆ�\IN�軩odqX�If-G�����u�Y��\�~��<G�Ww*��%n�;�+
��
��Y�r�=9�����*��#Cr��XTL�i_"�)vBoryq!�dɁ�#�_��U�Ls�]G*-*zp���
b�o�5��T#m��wY��_sX�=,E�d�rۿ[�� ���*�U3��O��`�J���́�)܊q#r�Z�K���LV�R��9cE;�b�ؘ"e�(��ϴ�pˋ�m������9�K9k���O�p�J��uQ�����ȸSMB�AQ$�7$,7�s�&;#����jgR���!U�ꓘP�'���IA�6�P-�"2y���B��!�^�W]`���j�^7�����kו�
Ɍ��{Τ\�	�0���@
���<��emיL-~��sz�8���k=�QZ|+h��`T�2<�[�oM�g��s��ʍ��˝�Ե�/U��(���oG_�^).u���T�B:�3������Ǳ���uxk�7?Vj=��@"Y-�Ք��|���el�z&P�m�7֪�	�ц�JT�JqUN�os G��]U����J�v<��Xf�i����D�p궺�2�giX蜍e`S/����v�Ӯ{�>��.���x�1�v��ԋ����m�;]��[�G�� �ú�&�wh�X�����;0tߒ}��Puxkñ���[��ǻޫ*r۩O3.AҪ�~�-�+�1�v�c(Є&�����~��c��5�b��3ǺI����%i�UX�p����]-9��]5��*�gŊ�KJ:]xޒ����kk����q3��P2+�S$^(�ɿ=�O7�<����a�;���	ņ2�zʎ��'��v��*^�L.��j��`�"wآXz��t�3�8o�q���f�hf0A�ݤz�إ�´G�kdh=B���+4����[��Qx�����u���fJǦq]��,�c3r$?u�y8ܠ���� _���E@0���:�mLu�y���9k���q��1��T;
t!�l���.Ku~qwf��PTL�)�ɨ�A�`z��p��3"���K$��&c�A����tƣ��u��+��vbE�;�y8�&B�"|�HD���I��i�җ N�8*�R
�T5}&�p<�˺ad@uHnD9�#D��i"D����3۽�
�&��"»�b}{7��%%\߳d�P[,(fQ�{��ݎ�6ͶTV�����ݫF_5�q3O2�V�è�i5�e+�e����C50W7��>�+;Y�n�'!��(1�����%�)6m��w�+���sꓫ5�D��O~og��&]n�:�S�@�P���T�	Og]���)!��� �:��S���];�n�H���J]-��Y���)B.�y�I[LHlh;�Z�M���+x��%i<x^|XB��k��P��F�^����/�|��&ޑ�}�79y6�=Z[n�/�(���Nа졧��{L\z@Bz�>�2/rmeؽIz�{|·�<�k*��q�Dsq1�q/q���{L���a�]E�Y��ex�:�I��SM�w�{.5��~�ͯ��2�9�l�z�����aT�E_)�Rg2fse�C��_������0�Up���a@��2Tm��;���;6��ț˄dcO%��3I�vZ���ԑ��F�'(�x��51� �æ/:%n'B���1��[�>bvs��O�)U\�qȸnpm�e!�tG���!�cw�D��A�,��!�
A�q[�b�$������!�YB�T�Z=�w+����x�@���IW�,lQ�w�&�rZ�yrs��+��k���Ԥ�A��rn*�'zHQ@�L׽=�d�s��Zk#�$I���ΎM:�gJ�����f�H���·aöVw���3���JV<�B���[��s�/.4F많��졺噮�fV��g��]�L̅XCn}�h���з�k 	J؝;H��E�;�����fN=��h�'=��Eh����bʘVa��{���[�2�I�aѤ@�0������u�&�.}]�
%j�t8������Ԥ��LF�D���lXi͍��
w2�6�/�l�����sG�Wl�0#Lb������W��q�O�Ԫ����ܴN��V�)�����0�jяc� ��pH�9M�ݖ�CrQ��j�C<��L��c�m���ya�������Ö6��-`�&��Ğ�n��Q���'��{*z�gr3+RA4�ēP���R���vԱ���1~��p��HzhE�z7jػ�S�^O���j���i�yOGY�>`<�T��e]���7T:ʳ�kDu���g��һ��O@�E8k�U0�S���X�vuZ#�`k] �� E7��B;�E=s98a�M�J��1n:@�5%ỉu*�q��h���W��j���?
-o���^���L5wmWB�;1��F0eFL�p�f&<O��^u��u<���h~[���Z�(�(R]֭wͳ1�����iC�(�
7/0�\;����r|�)@��U�������a�{���f����aG����0[�ʓ�˻bח׊F�R�tA\6��r=��
8�6��WG�B�KϤ��[�ʔ�$�=�/�F�rs���O���aW#c�"��o]151AP,n!)����,4�b�(]67�;�M�R�$Eo+x��$j:b�9y��/~n�W:L:Yh��K�*�Z=���ОV�f]��7{�. M r��f�7�x���\c�f�'	c:
T��V����M�yj�NL�w�ؒ��F3�{$:����1�ظ���И��,R�'yZO�5܎����x�A�Mf����s_B��Ξ�/)�̈��*-�r42r�9�7���Jo��ǝ��"֑�H`���'4�R�[�h��s��n��Z���%���z0�}^�=����^��`x?�}� 
���ҭ�s<]t�N�M�r���nߠp�Gϓ���S�iB;��6ܻ;�rƇPX�v$��rQ5�g���Z� �}�b�;A{�45�QF�:a*�p��ō�rh�#
�Ut\tD�U�":͒*b���ޑ�Wu���8�6"_�j& *9��oQf,o9�{ЋRuJ�$F@A�ȅuP�%�;դR�:�x�|�k�oS��e?g�R��;�{��룞�4�7J�e�+j��Ѯ�9K�,��f>������w�y�VzO�k.�Q��c�ħ1�@�&�`	G���2�n�=�ZZZݎ��M��(���w�P�@��_l���\l�.G���Qss�OR/v�7��A�8V�Skפj9J������l5�<�>d
���D��-U�ɉ������^��_/���(��m�|+J�zm�p��{����/Y�Nd�U�ߤ|$s�B��`��k�i�[��J�ȗ:��ӛ�Wȶ��}=Ҭ��ÌԮ1;���t��{���R�a�iT���J�d��a.�y0n�"�o{
OveVGc������(B���Bf�;��-�+�1�v�c(Є&,�l6l7\�W,]2L����Cp}@Lz�O"/C TF)AڧW<���<cA��ytY���Ժ�����Yʝ���G��}>���6T�H�Q-�p��>���瑖�xkBw���3D�.I��{�n^jM���ai=�&cT�0F�AQ�X{���V�5w��I������ܕ-��s�ť�tH�uDp'G�7�z�����L��_��)�#Gx����ی
�e�%l^�W�.*�W�@)��"�`@�
����Ԇ�u�$�Dˋ7�*85�������+J��Y`Խ7Z�8uܩt���I{���_k�qQ续�e��X�������I��D�[o6<�I�s��t��i)����O��D�݈�쾓�qK̦�8sr*���.�I��F����[!���r���u;�V�^Y룦�Mu�Y(W�Ɂ>�%�S(4Lm�`��6p9���|��O(Y�a�����~�t���wX-+�r�ćE�wWDO���r��QE#Di/Ҧ0uL����������Gy�w?���e~�bF@�e�Y�V}���5����tI���%
g����&/f����sy�C�@sH�ԧ/^���k�<Ps�����dȄ+l	�P�^��Tt�b��m�;�P��o;�&K���5A�W��g��B�xz������a
XC5��Z���^qpu/�x� '.���z�Z�xÄ�Gk�TMbv��3_�Y1�J�L,�'���{��+g�V���J]���W�\9�ePp/��DTsqQ�]"S��xdC�ѵ����a bL؜F4N^���O/U̐����gE"/.�6Fu�:��e�:h���q���u+�ٌ���9���d��8K��M�eS|�^B��=Y)j�ؿs��1��>�7	����3��v�fE]�ۨ긮Wy��cʷ�"gƞع�:��(9�j]՜��b��k��{p�Z������W�0��#���&c��Eӻ����=K������M�'/:�n����q��m^�U�;�w���{J��ɝ���:��3E4	z��3X�H�6��\5����f��|�N��oF�Y�w�W[d�|��%��!H譫�ܱBT{��l�����Q@vp�`�(��oѾ��h\��*���6��v৷Z|;k�^2��[uݰ�Kn7j��2���Yf֊Ke��<��s;wV�#Z�L�2vm�h7`Ej�Ѓ�G+E���8p�i�7,Cb��4��g��Y��sġ��u�4|�3xFnv�47�5T���)T�T��Ա*��gcRrWe٧gm��������M�ܾ޸. &�j;[�vVr����IJ�J�Ws�F4��iGZ�=aovʽ�r�gV^�ې�+	8 �ub��
}#	��C��)�.'c�ٓ��i�wjh�T��s�R����+��A���u�"U}�i��'E�[�G]�j�Ã��nY���V9��s��{�6U"��y��Ȋb�y�=|9�S�#9�`�j�YB���N��%���em�ؠJw3_fv1f�U�b�I���� ��קJ��:q�_*`)v;i��7\�������b�N*��`�$%m�5�
-i��j���T��V^GK3~�c��]���Ӂ�%\��͘s�k�<V������w��n:yd��::8�C��k���m����̔��@�je��;ǮM��������V��m�ÔFA4E[���qr�]Y��ӳ��w��G��bZt�\�D���z���	f�g0���z���l���QB��w�\f���|�OZ�G��3:��XMo�z��b��8�1BJl,�u`�"�����Юe��M���h���me�:����Q�(�1�+�~ܡH�N��BGi[�\���s(�S����{^���4�F�_+������=FsZR�Lf��eD{w]pt��u4�(^�\��q����)8>�4yBv�N���7;��E�ѽ��V+4��#D��2gne�21�%
Wd�sVp��W�k=)]�f�v��q��:Z�*�C#	�Vo�ɛq>��՝�9ѵT�At΅�7�N،[@��-��9H�5Uݞ���rΦ��Ϋ�!=��L���P䤏@N=4z�NXkFtb�N�s�9��[k{Odebe�gqkM9�Æ��J�&�oJ�$M"U�����ɴs+��5��e�w"�a���wl>��-e���%J�����������_bp2��z��7�w|�9	����c�m���YΈ��K3�5uu���_R3�Ҏƻ�+&���R�{�#��Ҿd��ü�.���+`�	�'� �����C1�2V� b
ɂ�V�s�w�p�`�eE�P-�J��,��VT���Rc+
��L����X@�ڔd�%E%B,���-`V6�Z�@YX��$�!�-E	Y
�E*�2�(�e�2C�0LL�bIQ�k
��UI��%r��q*-�.fb�C-��)Y�k��CcZQ��*-aXX�Ĭ��2bb�LeC2���-�L��%baB�bm�1m�E1� fXV�fcjT
Kj�
���	XVVJe��`��10AI�\a2�Y2�0�b0�ٍ-�*�P-��T���q�¸#i�!�d����+1�.P+r�9m��@V�զn,r�Ĭa�Aۊ
]�c|�ۈ��S%M*��;Hɇ���mغ:�anp-���o ��V�n�wj��*��6���|x��򚳣?�n�a@,䜣ӓ�a��PED�A��ț���^O�0�p�~����
�b:��(����^�$��Ԋ�z�b�8<���'g�};�ԣ�pw����KT��Z&\;�Ш�Q �l�L�51P�mV�^�`]�#"�NS�n !h�9�}$M.�&��ߛ��!�1��TD�I
��@�ޮ�}g��N�:6���ï[wbʘVb�M���ŋ�:�]e!tX�����E���M974��I��]FE�������%ڔ#8�hk���4�ƌ���U�we7y۠�WLխ���)�@�90 A�bY5'��C�"���.1���þ�<MG���=�]��^^���"l@�$kH�,f��@}�'A�<˫��&"�i���F�ͣݒZ8⼡��z�us��Ȑ�fَ����6%���1ףc�WXDUb$h�5�ˀ��<�l���N��-���ޤ.�y�I4��P�ځm�Go�X�N�VM����� ���rڑ�%�����X\#D���y^�����&��O��̲�;X�K����7��4�t����l����ۑ;�B�U�����3x�[��<�}��J�G��!����g�`[�����6�i�oZ%˽g��<tj��.3���&���i�]R��˯���U��)�����^\�i:�����p`(<��9�b�ۥ76z�O-O�I8�c4�A��".&��(o�����.vB�`�o+�N.w�pֿ'2a�����s��� K��Bx��X�e�0�p>R�2r�d��tWH�C~$�q��d�V���+0&:U%���.:�K��б�Ysӗ�1umON�������+������ì���²��Ps��c�YE�� M8��du�fg��i7y�w '� �$3�O�=�N���K2�f��EsL:U���JK�pP���I{���x�۵0?=`*|� �=���E���L8G�o�EC�b��TL�ӎ2�Q���Z�����s�ܙa�s�r�ﾒ3����~�G�}؅c��lk���O�1{��{6y��?|2���
�:ʺ��:��)�Ӑ^S���z��#Bjc�3�\>@ZX�//Wb��w�z�h�y�'ܑ��
�����VT��v�����ym)R�嘼��67����\n�-^�j�`�e�]��K��"׶���m��.�.J�ŗte��&�o��4�Ne!��ٶiI���M�����;J.���e�E�˴��G�ˑ�	�AgKf�&Q�[�nj�മa��}��H_Mf��9��o��zG����yH]���b@�  `F��9��f�Q�	\[�S�ݩ��ڎ�]�,�uxad1Xm�vw"���ıNđ0����	��p�j9���y�}*A��X5�Un�b��p���ɣ�jaiTP�rI�-�{���)$lN[c�c�u��k*ޅ������%Ng�(nH����cm9�Ad�zΞ���y��l��E�ڔ8��Z�J�&*��&2�l߷�H4�6�)�����C��ʌ�sΐ��m�q�t�mCQhB�f;�綊+O�m��B���U����F3���pk-g@Cչ��Y9���EW	Yb߇0����晊����t�튷���I��j3��jc4�ΊZ��%ޘѡa�iT������D�a2 ����=�7-93u�,��Ko(O�V���	�T��Ų�C�Lv���ʃB��d���f\���g<r'�!�\�`�Z�Z�vE�*� ��(;T���"�i�ߌҘ�A��'��u\���%R�%�K��|����w7����з&�����9��M`�b��k����EFd������tUE@�ƽn�Fg�i�u�ad�lofL�� gYS3oP�5��2)��7!��x�ocE>�l���y�.G��b,�}��'H0z�����Ғ��/P_=��$K�^�3�c��7���xt��K^�Md�M],���x��:͏�tl*������X�A%b�a��!�M����lu��b��9�F�󧧜�D;�:���@p �I�j"�ݱY�Wh]02�OmIҦ4��%��\
�>�"}Oz�E��}��ܠ�I6	�,��0��1��r@�$��O���>�fa}�_i�88\iXb�5yGKut�:��\�J����%���衚�����$��E��5g�-��.��K���E��=��i	��}tjo$���n�Sq�Z��@����#I�s�U�S�0xﯤ�f�G��wL,�f�c��5�wk؝��m8�a^,�=0cf��1����G���LSp��G��^"<�e�md�_Uv��M���ǰ��a��L����Q/D�2�[1V�o�Nκ.���-��q
��拼���������4H"+H��;�%�tP�Օ�Զ�y�	�#8�� ���K�i��,.f.z1�&�.�P���Չ�4M��G�F�Xls�x2�����A�'0�cɼ�+��{dd�!��U��s��	6�.or�{��뾁fN�J�K��s�u6�Χ�8o\����D������/K�Nw�x��d&.5:�%s������졧��Y,u`7E��k�ίv�{��kvG=��E�Ί����}s�s"�9��ۅ��6�u�tV�S
�⽴�,�ۙ�=3<�����eMDI��"�1^7:%q�Z#":�s"/#�4[���Y7n�b��yNH�4����CH�l7tET#K�,(4&J��A��;�0&��Qhs���U�]Қ���h���ݚ��D�Y"��1��@���L^tJ�;6u�k���y�@�DPY3��j]Fi|lb��n��^:%�s2D��T� h�����I�w8�M��d���/K�0�zܕ��:,�<E������qF�qKp�K��kҫx���z_:+��0p��+ާ\)טU��Gc�QꮜNFξ���\J��6�c���
�-]�����)�OgCe|��s�B��1�Y�u��NE�[u���ryp/�T`M�O
�҂��A��).�1���K�4��=�P`�Z�Huy�R%i{6������*�)h�cCUe�ɷ�+� ��z�JG8hG�A+\�Z�_f1�V[-�取��_-����=ޅ�]0��ҠB��>���7vd�òT��g;�\Y��?	珺tٔ2@p���8��$� �����zN�(�}���]�G��V�b�
��B����<�\�}.K�rx�F�P� EJOX��Z��`�1�g4�a3ZEÖ6�`R���N*��8�pU3�l߾�T�sx�y��U=��$?'6�,��ġ�nX�wTK�#�Fd��S&��]��*�������5R{��I�'(D�wj�%�)cEC��.:ѳ�}Cc7���-�͞�o@*���(t�e1y}V{�:�Ι6��D�1*���.��ڸ�y�<����y��w��\�! �?���9�C4��í��.�V>�@b��Y��+܋�O+p2��&p�=�����j�]�xmR;fJ^u��/K1�	��~��c��>L�0ۣ����y�5��!����^�Wg�	u�"'ف1�/|��U³�yM����e�9�o����ƸsUNΌ�XZm�#r���+�Gh�
�3�Y,@�#raEj²�]5�����\��@��Q�*�f�S�.:[�7�¯#u��t�t��GǍ��me	޺����$��p��Ǉ�ORZ��%�Φ�V�{��.x��G"��w�v�@�� OÙ�k6�4u���)���Oz��α*ݞ��2tG�f^�34���Z{,)��Y�Hץ˼㫵njK���|gu�t�J�6��3�ʐ3�Ҁ���-��D�a�@S�oT>6+�v�\˓��-s ��G{hi�c��DV�[��=-���<6�Hum�!L�#CY�o/q��P������	�^2#����uO�Ԭ�)����1�v9���Ԛ��W9�b�YK��V�����e�z"1�f�!�������V󎦎�ݞB��8����N9-w?M�P�����F�MfPǎ��yHX�y x:���P���*�9��ߔ~J�kM�<�jyeD!���׹iB1X[.�W:b�;�b�ؒ%�(���I��z�LY��D)#�\6v���X��w�s7�n�`uQ��d�j�ZjĠ�/bM�m�q.i��TIq�$f���vP�����TQ��9}RMy������@���6�bEq��\�O�էjf5�vQ%�����K����Bj��%��.��yԃ^\�	̝��S����]���nel {t. :���D�ƢЅt�g���¶�)�	�dx��v�[/��շ��J؜�#��H��QзB�Uw!��m��Jǻp�|# 	��f�'������y�n\��DS���&�[��q��b��8�\�M����ys���Y{8�}x�5��iR<�����5�P��	�����uwH_LcI����K㫐㵫"�����b&2����s�tL�~��^4��Q�Ό����QN{oV��uʲ�#n�Y��Eyk�M���e;v�֒����c`�<��M�����H�&��v��@�۞�fa3Щ�Ɔ�%ڔ7K�ٌ�Bۮ5�Dmܘt���Q+�J��gFٸ�:DZ�&�%�.1W �(>U5
���p0��b��{�f��Y�������'7GM@�(�D���K�����)�1�Qi�E�CZ�;����b���Uʕ}<7��<���p*��j<�EVzSn
��&�KGs��Yܹ��}D�F`��v���}+J�8��ù#�!���p/Pd�d��+<�#_eFǑ�X�yH\�Ĭ@<A�m��f��l��6�O�tF� ��"7��A[%1uU��Þ=�1�\���L�lu�Ұө��l�޵�Qϟ�l3�\4hg��b�Be�=h	[4p�(g���6�B��Y.��s��Z)�Ӗ��VY����1�T�]M.�U�v�����Wk��&��J��]�[~Ë���ֽ��^⌷`aI����w�f�w`�$Ƃ}0��w���%e�رo7��f�kH�����4��ׂY`�v%O�e�@6M��w��o�<{�wP��)s��jk�d���}N����$2kҧ����U�H���˺a`uHj*��'GFHV�}ǚ�9�6��Ѣ�)�*$��!<MD���|߄�����z+�Hy�Ǝ���<p��^8ߦqA�m{�y�]�לő\-rB�:��z��h��_�i�^��yC'�C�b�1Mo���;���5�{m�B/��P*����chА�qaTl���R�i�݁άt��j�!v�8����<�Q���8���*&��=��7��i���ۭc�s<�I(���k���bym��pg��b�n�{�]e���<"���F�-v�����-l��a��N^-�͐��N�0��*j%�yt�Y�H������4�Df�k�F�eS4�I�����9�}U��ۤt"e�4D���a��l�A��o��ɿm���F���K����ͫ�iT=0��ݕy(m���yh�f���
�.o�0�i��P�\��|�rfspvQC����-[�(�����T�3芭{�W�:��2��T"��ѿ�W3481��`��ڷ{[�ӥ���gBzyGl�.���Ӹ5��G�>���gN'ϯzl�aS�S*,w�<ڍ�5;p����#ef� 7I�:�3���'�e�W�qyOL�Q��,�
_DgI�B,��ഠ�T�Z=�I�D�P-	�"�ݪ�ɚϏ"W���I�:6����WJ�A�OR@���Ϥ���j�x ѻ���B�f�`BlL��U@��������Qe���3�����_+�%L+1���=���*"�+�N瑻1c]��n�;�k�`u�����X٠��=A��â��Ν��"��p�g"^V�N�X�״.���&k���a�����W|+R�D)���'�j$�Q��l_W�~�rx��(���^�u���t��d�I��%\\�:2f��r�Ӻ�$O�%14��Z��*E�ŵ��E�v�����zJ7|�Ċ�sl��ꖜlMط,mC�����DPb�{'1�w<����l�ԺE�K�����{�Y��Q$�',D�T�o���ũcC��9���WŻ��|�4o\c�qj�7��awLX�,W9�ys���'P�T79��BԩAl<Ԟ�oNU����L>l�gՑ��l�ML5�*�)1�S�����:���ys�%�G���7X�xG�SWY�U�]ٮ���JP��)�W�OD5��^�Dl��p�\����-X;�����#�8,�%�ɱ�[у"�mf�yW^�@hgnUn]b� 9���M�j�e^j�S��|;��bf,0���^���;���j��Ku*[u�J��4�wn:R�^��J�NیS)�b�]3��x.3R�w�;׼ҫ�����
6�j&������}��鏠L��u�)Ɔ�`���Qtr[�@hcr�Yx�,v#4�,��bҀ@�M�2��[Őj<�|�W�n�(��P8����5}\�d���hȇ���tY�;T�d�
���j�̬��쏞;�y��o�$�@�s[�mqw+���n�Mz�	�,wP��-����K�g�4��6 �.�%\yչB,���u1�����HF32���j�'88��s����E]�tn�۫��+����'��z<���ɵ;�̆Dv�2^�qm���`g�`j^��^E�F�iĮ �
��d���L�����Q�ʑ	�Rx���D�5�Z��n�d�����
�	9VN3n��4pV|"�Ў�R����32�i�Pp��)]o��Z�����q�vo�
�fh�C�=���p�ˬ�ɍ^��ه���w��t�v�N���jV�r�:�FT��;eН�B�M�|��� ��#IVat��e��w�+]��FKyJ�dV�nV���@�����P5��+��p��a��j��(S�o,���}������ƖSӚJQq���$���M�׷�w$э�w�+|Vh^��
���s(��V��m�ޮ�X,kneܗ�.���V�ǝ��*V��:��-�z�{�ܺ�'yw+�+\{ah97�B�Ӎ'v:v��s��KVEKI��[{�B�'`i�e�YDN��QO�Ͳ3���Fr��ew��3Myf���2exxktV�C��O�O��K&)Q[��ۺa�j����r�D����y�q�ų]�]��}�֠+�=-���d�4���b�J[��6F�\9��[Uy�a�B�z6���Oo�
ҁ7�å��xe�0@6p�u_a�M�Ki��07x5"��x^�+U�X�N��Dv�N��vk��K;�G5^ �]M��:^9V�E��jf�w�5J�Ff;��3�[v`�VlU�R(��0N�d=�}{3p�x��v�2'��
}c����9�i��2*7��|���b�ԻE�W:w)��as��x⴯E�w:\Ogt�鶬�G���|՚��f�����e���&�݊�NM���ϳx�Mu}�j
粯Xױ�D�K6���}w�v��5"K94Z�����,lōd@ukY�C�� �"�.������γ�tM����к�MD�ΐ��[�'KE�=��u9fP:�ͽm��]�{�;6yE_]�_+$S�,�$�%��WLF3���Z��?w�P�n8��*�%�H
A�T���°R��Km7;����ڠ[I1PDPĢE�[IPQJ���
��mb��F���(��X
�(�PQT�b�6�TH[bő`�P�J0
�fY+q�b ��� ��ʒ�X
VTX�

�ŋ$QB�*(.9��AL���(�,�T�b��X�0dXc,�C
���#e�-YR�X�"�QҪ�U	kJ�Ҍ���q-�a��Z�Z��R�
����0[lR)r˖J�"V��*����%B�d,���A�Ƴ+m[eq��HcU2���m����jM%@V�;����;��3�%���;T�S�h.�mD2�gm�O�DJ���at"�+�Ӻ�rrv;6�@Y�ݒI�G�/�s�k�9��w_�󰪠l=y^t�����'=�/~#xfЃl�sݝV��M�}�a�S�4^�X�O
.;Z�.�F��3�kѷ���P��O��aq�
<^�����{�m�P"���q�H;UNΌ�E��޺b6jlXłX�f����.���Ƌq�t�O�kq�d��$Q.�&&�Lt
��Y�>L��;�/:��8�ͺ���&�1�x�ۛ�rc]>��}�%^i�Ɂq�$�z?0=�����s��W��^������RN�M�E)��Ч�ʲ.������K���&�Sd�pa��{$:�o�
ꈦ30k9s��V�*����_V&8 �T'Ywg����Vd\�ON��ef�טn���Uw��CR!�ms4)�V)�rF�*�'Ä( r,��]몚:����i���7��ʞ��Z9̺�ɫ����y)��� � T+GnɱM#��]���%kz:&K��5�cp����W�1Xn5�xz�i��~�?�đ����k&�]��Q����.����;ˢK�Ҳ]��U�����C���X�ړ�R��¹ǗM���wq����j�+̭�+��m�����N ��L��x�=�ͨ팵>��r-Y�V�˜{����\��J���զ��wȌ��#owr�<�:O�(GI��l��7�f�(����˷p�:��pܚ9���<�'i>��Bz
���I>��GY���Rk6�%{��Vk��Pa��R�3W��a/����������tDlg�۪�}�Ib��^��:��\2�R�pʡ�}o�u{G@��j�­w3���@KɍD
�BP����D�Ҷٳ]+VY���W���w�Qh�Z�wv��LcUv�����<;���u8+�Z�.����b&2�ׄ��o]%xd��_����jSw~�,��:b�j�C�����Q����N�7�)�ѢcN�Fd�^�P��nU�QhʽM�����NeMDZ�+�k������U	��N�46Q.ԡ�]��L<�μ|���'�!�5;>J��m`.s|���D�z< ��p����]-;��,	��T���PΜ3���Yg����6Ϣ��]IH���d�P[%=�#.�R���z��3j�u(��e=�~5��}s�F��tL1P#�������T�p�YA.)'�i�V�w0��W54𸓡v�]�u�ͧ��QϺ��ʘ܀�N1���m��cN���2E.w��
��C%��~�$4�egjM.��o��x���{*F)�ۻO�ip[�r���[<���nQ�rMdl2��QWL�����F�H����d�F�w3�KV�5�
�n�Qc ��ǜ�;�9̑�h.x��	�Ū����[�����w{��ĿN��tPA�F�)oTH�+��-�C��#�:����&c�n=ɜ�ڙ'Pѡ���An��S��2^��:���=�+B��]5[�P��e�Y�W�[ rRֻe&�I侩��rt�~|v`��f����Y�G=.����9�ى26Q�ܳ��X�^�k�[��Ȏ%�^�|߆��GJ�b�9���H�K�ae��N��S;8������iʱ��1�TE��u��&�pZK�r��>o�LSp��G�>��p+1��We=�k������l��9> J�x.�!��!\lW?R�.�u��xS�������}������\_��"�7�Ě[m�P*���ckƄ�+��
��N��h������Ӝ��C��^��\綠s���N��oz��}}Lm��)�1W���\��Î&lc�<3NQ�6/6퇾쮲�dG9��Tm�v��z���D#��/h�;m����9Z6%w̨�l�4�УG�c��#<��.t%K�VN��Ύ���~ە�ez�z��f����̚Ae�����z��kɏ������|c�K��,f&v�9#�u&M]vM%ϷsxY�/Rq�Ӊ��}��y�x�ȭ�0�5���+�q�p�|E���#��w���6\}n�;�=/v�%��˝�5VT�q�L��'
�b��^����`Й;��.z����w�Cp2�n��]�Ī�����t��ᅢ<.�~1f��t�����f�V��n����'�`�y.'B�S��)u������RE����D��m7\��7�ef�ȌY�ƈs�1��D�!�y����	h�|�h�ѥ/o�^O��)g���s8C�X�I,=���z���ӏ���R�G  ѽq0�d�(�FNˋ���4�^��:����<��_+�%L+1�n����B�*�W����C�Q[��7�8���Y|aQ�@�>u_L��l,;��>��R^9b1�lnj���=�h���+|���mڣ�&^����}��W6�P��|L�w��T�k�m9,uW8ѽ��R�ۙiڼ�h�Xx����]��
]��٭"ܱ��+�(��Ԕ�R-!^F�ت�I�ױ�-.z����+��͕�mᲰ<���<<;�GW��d!1�^	�f�vR��+M�L�z�c��� ���)
�I�85u㬋�ݜЙ���\���-��j�";6i"�V��h�h���+p{�1�O�l骮iu8�}�6D��v�����Pl��8S�1"�9�adT�����r��;�\,D��$S�/�����جO""𿑱zԧ�����^����})�����nJ;������}�y����9�ߪ,C2�W�6��}{�I�|�S�=k���ӫ+{k��7�#8-��!�b�ĴV�۪B�d�/�L5�U.|�જ��<6b|Gj�5���w���Sz��������r�X����t�Bx�Gp���ōE�ӱ�rA��2p��i���S�:�Я�X���kVE�ݨ�8΍���^`Lt���J^u�v!�|��u�]�>�5��I�WC���}����o�����o]1�����X,^!\漣��+� �+9�5}�a�Ⱦ��*|��T����t�硖#6f8C���R��Q��s�O.!�&��B3<Ӡ&�%�*/����Y��a�;g8�u���P���Ŋ��f��8Kd�$�q��MĪl�q�&{$4��O8�{��4��@�*f9%;ʶ>�w��rps�(�^<��n^gz7���1hf�ஃ�&��}H{��W+��8�[(��1�^���l�]Y|��VU�]v�o;ؓ}kz��+��쨯�%
xy�*8����)�|��&����SZ�b41A�.���"4I<N� s,��qJ���=>{�&a+��1*�OM�Roϕ�og����W��
O;��s�hU��
��ȩV���Yn�T� �Te]��¡Y��q�iȂ�;<UF���x�a��yH]�<�>t$D�*N8��g4T��$�2_�Lr6��]1�]ǥ+�� ��0�9���tr�1B��K��	�+�}uy�ڤO$0�Um�d��+Qb�b�g��ל�+f�n]�p������ȋ�
�h���7�Յx�w
�P�$�NHXn%������|~��b�{�Pa��g����"��}���w���`?%$F@���F�"O�>��yT���*qK��ur��z�s'��/!Q��u7� ��/�0���(\X�Fa�e+�dzo��f��
�u�FԦ�㓔�aq~띳�3��.�E-jȸe_0�]e-[^��w�6��:�,���<���U�;U�Y�W���W�h�=S���Q��&��)퉍4a<|ƴ�3�T�/�4��]����`�Uթ�C�	����|3o�D�z�5̰��b��p<�~mW���{P8BX����\��{�&v.�S�u�z�kU��`�ǹ.���"�'M�s��t�|:Vk�C'b��y��us����{;�Ҥ�ort�G{��p�]N^�l��y��J��n;�܂�D�r����.�xY��[:�^@�X��x��+�倹�	�tKd^*���(;�N�Ymy��Z���WNj�,�S�a�uj�MIg<=�%�9E�<ܨ�S$Z��**�O!5Bژ�QYصP.�V!��Y�W��F{��2���Q�4��U��+Q�&c]�U8*����Ks���/@Oo�y�,v��!�[��X�/�q�pW�s$w�bxD���!�6�#@r�_5��Dl�[�q7��tPA�:�o\H�W/�q��ú#�:����fNmn�q+f��0W���w�a_�;zr��B�i��.�U��:�0��xPb�ۓE�w&w+�����&�9,��A�q0P���P�
	쬉tƣ��u���f�⍃SO"_%����,�4��-�mү:��[Ȏ%����6�TgT*�Y�D�fg4������宩���9��C8Ò�t2�L:��?�2M*�Ik��9�~�\
1��^ջZ�i�w����=�4�[y�'GN�
k쾲��El�:�WaR����W&녵՗���#sE�j؝�|�]u>t��
���YyV�]vG486�v5����p�9��l�}�A֠�.=J>��z-]���X�wy+Q;��ԅe�aXsH�~lJ�!y�2!
��&8��Q%��e�RP'�e���^vu�1��$��hпE@l��c�8/q�+��^zP��|}��Γ��[e�����笣�|%T��(�綠������U��l��t��]z�ubh���X�Wr����61_���o.P�ͪa�vWYp2#���\�V�D����w��u�-�4�'�;8���{L��F���*jT�yR��ΊD\eֆ��lx=YF����c������'q����@��������C8�e�O�(F�l��M�Lճ�*:���Rm�\� ��.L��^���(��}&:���Dx_`O�s[O�U�-h/ڻ�a�f>r{:�@�Q�pgD�F�B�S��B�Q��Օ��8a�,4��h%�[�.�Y��'�.4��p���L*�Ȳk�Y��C>,qS�ah0��pѓZ�L4��9�c6yp�d@�������L�9Ԑ6�^���"�m*<hߢ'�bi��ex-d+1aWYfI�Vh/xj��^�V�f�8lZ}S�&,��3;�pK)��4��X�7��-Y9�)X���v���^T3�1M��=&qN�v�����bè�:5����q���4_fpYj��;���y�*I��y���Wڃ�F�_�na���T���s|��쪅�/�n�ن��t��\����[s���mh��M����*5�|�K��zPW�A�J��1;%Db���Τ�K�+gf�ScFE�wʣ��)�0 F�Y7'�똔:U;��ά�[�I��Ag�`��<V��r��U�W�����Xڇt �BRx�<}~~~;1��{�y�Yo��hU;��CrQ���$Rsl��T��bhl\K�[5�~�e�HdX��I�yY��H�*B��,>fa��5�+7Ҥ�NX������Q����"�tr^�m��~�vYk3.��u�压����:c��{Τ�\�%:]BԴTsF�S|9��J5m��sο	�Z6}*�U�G�K(p�-��¸[��Y�1��zT���q��x�U{��XL6���Y{@46�e;߯!8�h�`c��>n�L���Յ���bF����1�\3�konB�1Ғ�}��Y�6vj����N�x���j�6Q����@)}ү���ܭx� ����S͡��������B�v��o@�wS/Ec�ޓ�5��S��v��k����Yc�1ǰ��0�'��f+[oc����,���]2�)N�sO"��fNS��Yru	Z�7(�{enʳr߇���~�UN΄XT=t�nDT�Jİ�3U����˺���[ðS���,�cIص�a@���p�ɚ�v��8�z��C���"�r�`���o���Q�₱��Y�I`|bKx��`'�� u:@H�e��L<�1�]��sc�ާ���⻢a��#
�&`i�p���頮L�W\�ĕ-�;\L<9���u&,��7���*�$'�����l_����k��`TN���珢+GJz�*t�Ev5T�RZ��+�XF\�q������he���'�$c�0"`p�`�G�I�mD�n����p�oFGS��*,_��=9��; ��\�̡�,7�����<���x$�5T�op��[��	[Z@B�4kx�5��ߥ+����
���tr��!nO� [�,}�ܵ.ܫc�!_#ēµ�oY��4�af�۸XT`��,�ca�͆�D�l�i����XTI7�䅆�%���B`m<�j�899�o��r]�3:�9 I�w�cqʟ�u���4;�[�|���`玘���ƌ��L�h��c��b�s��^����@�TͻXց]���:6C����v:��ӻof���Z1���uk%n����S5P�t�.��X������;GF����<P㣽R+�e����J���*k/i�5wSo��b�f��mVvu<An������Cs���örq��m�x���ЛܹT�ʳ��m���VNk��y�Y|��������Hs��4U���N�l�� ���b�$@��U����吟��4�W.c%��qNKq��kX�C"冲��z·J��L�\G�{�����n��'S��ή�G �P�c���}]c��R���֫�w��z9G�:��)m>���<
AC��X�=��Wr)i}��;En�s�ά͜L�AjS��5��{ҁu�L����E�u���&�$3zdm�*	���rIу:�Z9J'wr��:�Rv ��73a�˦�/ ���3PX��JW[�������!��{����`��ëf����+�%\��-�.]ens��G����7���T�:"�)편��qˆn�w�M�����՚S}F �[�Q'Bv=z⚊��L̸����V�.�y���Z���]â�	���);X6���������[/U'q�Y�c4�>}0rp��oqҴ�q�j����41�lܮk�㹦s��g��+w�Qo�gB��H�˗"�q7N��vb����f�G�M��0��Jf[��=���靇���rp;D1ã�yo:��AL�u&�V����ܱ9�J�mJ�l)�Y�&��j���[:֧M^\��h�ܺQ��W�*s��x�Vs��>-�Z0eZW��8�ݕ�@	�f�F��:Z�Tζ�}}���Z����M�6Ьn�4����X�4�\�PV��9Ԟ���t�����H:y�І��g
��꧒�mLUn�&�b�)qS;k��K6�<IҐ���IK�K���o;�+6�5��.]U����T7S�};�Ě�����\�uڀG� ;9D��I��0���;��Wy�:����e�c�L�R�ո�X�C���S��pjܣ�5nF���I���hJDp,e������ⅇ� U�RZ���y��mXbQ�q�VN�r�Ԉ�/�.��}���.���^���d� ggY���
�d(�Ԡ���V��7MeC&QE������b��[�uL��Gg[�]��[r��.���w8�z2��`ήJ���JTT�Zo $WS��ruPjάrW>Y�Q�r�mDR�n�y��8i�V���0Y��'.��1�qux͓�%*�7ݲ�ewdΗe�X�uXRs�KR,5�Hy@���Y�ۭR�l��Ȟ�%��oU��^�`���T@XƵ1�T��+�´���jV��A�h�������}��v�!R��@�*5�X���TH���%*c1R��,�s��﵊#Qb��(�*�ؠ���H�QZR�׶�B���Ub$Zʈ����c1Y*UTe�+-(((
F5��-�iQ[J
,F)+-���b�R��aX��(�IQj+�QE-��̥��ˍD�T�A,EA���J֌�YV�e�lF��+-Rш��EFڅ�mPQV�ęlDUb(�X�X�UkFF�¥h�-ePUQQX���,Vm��X(���10V,UT`�FV�XQ�Q�V#���l���(¥���b
6��n\(TDk�%���j�*�`{�o�>���y���tbu���!��/M�T�-��u-�$KN�ѝսw�7[�O\�Z�!��<���{�􇤬���g$22g`~�)"2y�����e
�>�וK��qK������{{��꺱R����qp���s�&��D�@���R��w��8a\t�.b����ޭ���=�ф�6�
��G��g��.�B֨�,v�����ʆ.;V�7�V�y\bz�ԞJ���L�ȳ`�S&��9�L�?~�{K�����]���&�>}o���z��tR�08]'J'��(a=�r�E��p6�p��7
��n�'X����V
�ו
I�{^\s��XB�O��ץRV=d���P�[#b1W ���Aº�����fՅ��8t�.n���f���Q"�.����
d���E�t�v�u���M�QX�͞Ծ�x�����sK���M��tL!P#���3خ���X�Uti�P�or2���A�cI�����CQ�ug��j�h�;�:�Q* �a*]H��G�0O,��WĈ��U��q7)�'E>�t(��q"�\���n%�H�dTS�̤ג��xIh��Y��F�����3ԮkG�W: Hq�8h�_ѽ��玙�:)͍��%�#.�4��d#��q��b8��q�4�۬jIONw�=�ӗ�`�c�����X:�XΨ9��-9�r�򅉉��+��=G�qr=�;�e���:^ ���"�T1�Qީ�r��9\��9V��������]@ΙT�y5��2^.����/�K�&�ɨ�A�q0P��3 �O(g�wX9�������.�������.�&'��EH�W.��ȘU
���HD�D�aT���*���&��霅�d".�[ܳ����n��S(c0���0�&WFI�]�i.�-q����k�Q�U�m*7��Q�7����ީ:,.i.���0�"D!���'���#}�z��[����v^g��+ir�x8�(E�o;�5�ѡp�V�,mxА�妀,��^��Ԗ|�������i����)x�;8�.{j��1=���@��f�H�5����W��<�f@��}W-�*?�A}
�3�B�j�����ˁ��xE.qQ��8����.z�"s�H�1��*�޼cv�{�g"T�w�HW��E�ֆ�0���x�w��u)��uP���H�=n����*����(�f�O��aʯx�žF�zd~����s6��t#�z� �ף�y�Ou�o���k���\�f�.c]��+��m	=@T�pRI���)#sv���C���Vb�B*)v�N��{]ut�C{�*K|3T6;���Ԣo;�>�:�d��U�#g��4��WD���'Q��;���2�_@��"^� �S�������t�%�M�-Yؓ�`���C�^���c�J��cK��eFҁy�,#s�P��1D��U`ܬ�
�n��sV`���1����Ѻ(�����"�D���d�!�z�W�|X�*w�Z�0��d�u�MÞ�:ӛ��Ã����DP<73<�WU'� t!l�9�/z=�	R1a�݊�O{������!(�b)И�2t�IÂ���A�*ag���f�5޵�b��m�j��5��j:wo^
W<��Q¢���<�}��Qr�0P{Ԥ���Y�y����fM�*b����R�x��^y�E�9�!#Wp�MI�{7N,Z�s����=ѢL���,\F9<b�*����������9��@C <���R��0����t���)��Ǥ��b�L�y�(��7q!3L��T����r����yr����h`q�$�B�RX�S:P�a�6�>.�Α>�/
]���ڛ1e��t{���'�_ZՁ�&צ�=S;$�H��S'����/m�h���QV2����<�6����vN��?:��V��]9��<�T��=���-��&&�����9�D)u�he�q�=� Oc5���fVB�MM�`,��I'N�!�wy9��E��jс���	�٨
�|81վ~�8;uV���؛�⳺��W�r�FJ5�������<Ƴ��?r�����?�e2��i�xP�C��k�=|�[���/��1���`MB�`��(n���{"�f����udh���ĺ����)I<X��{��M�G]h��K4\B֬�{�����!��4�Uּ#���-����~Z���u���o�J3��+#�誝�0�����ʜ#:�=wf�t�����m��z��z%�	��V��uW�f�TBf�S�c<y��衊��,�1˟Xͮ8sn�PU��0�n�e%�����\���,Q�@�B�,�[�ƒ�{y��N�]a�nnR�������|k�T0�d��֦:U"�r�6Īl�6�wɾv5s��QШ��$uZ}�VC��l^�����q�'Ģ]^�?�����/�n�=�;P�쓽/�V��!�q�i��� u,��C=i��Y�£N䍥T`{�(ճ�DW�FWL�˧U�.��5�>�(�`Z}.�}���feߞԒ���l��$Fv ��j���3���a�V�<��d�,�K��Hs4�5�:p�N�����>�]�Ĝ�Nd��Sq���|sOjw�j�r �G��t�![7�u"N��4�&��%��ONAyQ��UF���ex�a����ߞPs�9]���Euc/R$!) 0��l�E���6�+�8.�,T�Ԫ�����CM�U�~���#���V*���ı^�D�rQ$�'�f޳|j��9�L�V�/zdi��f>x��g�#�JM���zi\J�I2ܐ��K�$�~GmIF����'�\��:�)ӎ�+p0��+�TnH��P�ªf{��(Wh����cGf܌��s�Z���[Jt?��F�s�%|@Pؔ ��⹨w�p¸��.bf�����k9�$�	�YS}KK�=����G�P�	czo�H��Ր���X����`ʨʢX��b�OA�HWl�&�ә��*ًͪ�;nzʌۨ�l7Ebt���Hwf�[S{�|7Ry�|٫�~@ܽK�lL���,lZ�#nxC�ڨL�uQ�T�n��}�l�E8Gi9�Y-�ꘪ��C���X�1r�\��>�|�x �ǳ�9L�1�QR|����J���ҳ�W���Q�B��7�='��:�8��\�+���e�i4:�h��2�΍Yv�ƅc���]L̖�B�̴;��ی�Y;�0oa����!8�ѵS/8a9��y��5���+�5y�;/uwH_A��I��z�GWU�A� 0��U�C�����K�F��^z���啶� �{���+�\":�6Q"�
�[�b*��y�{<7�	�7�5'����_Z{T���c[���o�
������\b�a�>�z�F�/�V�i�j�h۹#����@N��0T��B�@���-�IJRޜL�0We���S��Hj�}��;����t���ier�#�2Q�����-�Nޜ.U��s�{�V���$���^�/o��w��~{+����M	U���ip�還LV�W�VD�cQ�õΓYM����~��XT{<Ee���J��f��Dq-r����z�U3��ky�dk��u�]�(�����}|�:�7<��p�.�a��L\$'���<g9뵢��+x
�Ż���mU�qy7���RU��7�C��9�@�ĭ"�!��D!]`L,ƚ�{o�U�|�y�<��K��
k�\�Tbμgc��q��$���ѡ~���+	��cT�7K>���R�>Yu�c�*��p{73���b�os�R
_x���-{�w�м�z��3:�1�3�M�����<PXwna]-u;��hv8�z_O�0����vu����WC.�k�C��C���F�m���4z�*��|�v���N�s��^۵w���\X�nu���^�K�xNEs�ڀ\.qQ5�ڀrչr�f���<T:�q,a�kс�Lz'�
��T�TW�b3�e=�\�-�z�UOd��J8�풋���n&��B�k��m��<N=�1�JÄ�3��N�+�q�u�I(G��lżQ��N�-�m�7�ٗX����[�z΅92�FM3rxEP�	|6]��i�Ӟ�<Ufܫ>ã�7�H;T���Xay��;��ߦ�*��eD�d#a�w�wSr �Â�8��@��Ԡ\FtJ�c�v�ъ]F��X7++� O=��@��gKTyt���bpu�L�A��.&:�"ɨ�!�^�r/�T�|�7F������|�O%F�g6D���w��@���Ȩ�d���u}f&�U7`�~��~a}�`�r���L��ߛ�"�F�v�̢��ߵ�B�܈�vxٹ!xpL��A�_+�%L+0��;y�����Ry�zmp[��X�xT[�x"��#vS0�� C�:�t�.����Pd�;1j6tQz�%���9KsCVm0��@��L��6�\(�՛���[��Ҙ3��]�pV.d�g�an()��KGX]	ϫ��Ė��M\o.��s}%tn��tN�h&H�i̓]���1l$��u��e8�v��Ό�l��"�x_q���/q����tH��`����yخ��,t��O<�f*$`@���,����BrO-��I�u)�N&%^�NK�O��J��.�B.���c5� �Z��eu�uK�.����@q�&����Ꙅ3׺i˜��w��HL�0�<RӞlM��]Ѥ/�!;�N�~�&XDW
�H�k^.��]f��3]D���%��-�̋'%]�������[�7F�ũcC��3��K��"Ą(]s�*�6�-鎢�e��z,�z�3�u'���%mf�mu_��<ê�߄��l�}��?�*�����EF���\�R��xu���cC�\�	[,���0���W"�f�Oi�����*�rʑ��i���0?a�0���{ѹ�a�G]hw
X���kVCܘ�:΍��&e
��l{.�B��I�v��C��Iv:�xU������<}S% �U;:aax���s]{m<ͭym�$p�\
����c�X�JK�	qz�?OD^���7
���T��L�Y�eޮ�1Vї�������*�Y�N�{h �ȭ.5��Lw�*�:��\�{�����}�Vc�7��v0q�Z�C��㚸f�"��!؛�YH�%� ��r�OvohruoM�U�)�0�+�Ndw�vF��9ʕ���;ۥR�E��3�c�=��Lv�%lL�I<Ӡ&�%�/�	���Q��4_B|�TK�l���P�Y��j����F04�8Kf禂��3�/"��bg�_I���W�T��́;۲�7bc��$>���c�����v&:���$�*��P�F���*&F�Ƶ´{%p���Vd\�ONAyL���@O�moi��A�'��J���t5��.{).��
����b�Y�:�xE���z*���`�M]�v�ڹ�];]�-r{�x�;k�0-���" ��J�tQ�S�f��cp��JW5fD1Xy��ʖk���mou6�������!B�İ�.����#�Є6b���IF�L!�Ͱ�W������s��o+|U?U��VyI��~SMy\J�rIl�
�z\����링xy==��<�h55��Yϑ�û�Ih�°�����5�{���׵R���8��8��/��>s%�E\��,l@\U���s�'aL4@�lJ pb�\�>�6a_�>���	V����x�<��w����ϜY��}�u���gf��&��ѐ���m鲁���匿��ep`�cT�x����IM�1On��^�����䦕l�R��NTs':]Ô�שּׂ[�uwhɧ��R�M����\z�����v7իiE��N�{G�3��_x;��	��"�ͅ��K^NG,�!�	��[�+�ܮ0m���3�kın�6���ͻ�2#nzʍ��g�ptbr�z#��R<�:��Rbzt�N&4h�84:�G��%�dK��yx|�l��y�qq�P���МުC��lor�^Y\�-�E�O1�v/f0H�.��s8��`.�0����N	�OIi�Z�W��
�]C@�R��*up�r����k�{)F|]
�K���y�:�b�/���������dK�E⏩�N{��D��n�N���m�8̞1ppL!ʄ'V�Rهsx��Y�z�U��<8�}R�܇�C�1���[]�#TKF����}�;���	����O.�82��
'�� �G+]��q:���:#]���$*/�s�X�G#14��*
��I?:���EI�Y����L+�����a�+Lg�㵊�%MW>�b�Sz:�Ϸ6m=佩�*��:�39�fmBsqf��3�S?�y�ygqBB�������e
�(�QW %$� V�I�}�*/��$��VS��A��*	hP�D��7"�t=����g�r�]��0�`�2��JY-) �R�$�Zu� ��"�L��*�*�R��	?��$�1${���3 @;t I	=@5�ZP�(��AA�EPU;���"(��ȣAEQEPQ@T�b���<H_����P�I�r�*��dn��H�O�0��"��,B$J� ��ya��G����~k�����P��8�
A-�Ń���T��Q+��7�S2He�Q��d���F����!H�7z���/� W���<wi�sS`,����\u�* +�(D!(�{��h�����?��BG�˽S�z
�����N���a�w�Px�Ğ�T W!ֿ�����a�! � ܱ��h>
b��Q�K&Z'Nc�2Vа���P�'��̟ڦ���,UfnP�����;:Ѐ�q����7H.� ��<�?�䈢�ENV	wa5�
8i+��]�Ԡ�@���I BP@��<d�!풌���2�1b���(h?"���X�>��D�.�F�ر�o�E��RC�
�$*HZАA�(r.(k���GHc�9=��	d&�CI���tǬ?�	��Kl�R�0��4>E�à�`�>H�~G�i8;���&��� �+cֲ:(�!�G���>bxv���(`�I�o�% ��ݡO��$��x�{�A��mq�7<H�Po�l'�:B�J����y����@vMt���1Cc���` =��t�B�}���Aݑ$!�R#�Ѐ
�A@技
�!�?HMX�!N�%��:�P�����AqxX>�8�AL�@�(����R����
3@��E��,�ea�L�ʀ=�hd\S
m!	r��L���ā�eV���*��R�� ɉ(Л�@�GE=�/��J��� ����z(z���gBQ�h* +6�=b��@��/��N�l�S����c�~A�q�N�{��i�P׸J����;��������z�G���t�lxBy!��E��O��s��@��>G�H* +��yX�Y�9 0@A�&Y<��4����������2�������zw�<��'C�CD�}������ ��
Ђ(-�8��q Wޅ�gՠ�aLOb��b��?ȋ���=�,:
��ơ�n
�
��1;�^��C���C!P�/3`�4@y`$�>���:KnN�@��#B��y�$�h��ބ?T$`<݃�u�0����a�h�@=݂m�AN�G��v<_WX

��~��=�rH��a<<$n�	 ��2��Om����)ԑ		D�� ��Ew�p����)�t�3(