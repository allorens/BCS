BZh91AY&SYcu2�w߀`q���&� ����bN^�         �ʃ�`�mZ[�V�bim*�)�S%Q���k[4� &�hj���U$�%ClR�b�)UF�F��
j���H�Z�5X�v�fm��Q�m�R�R�6�TͶY����A4��Z�Vm�V������l�4�V&�V�&�V֡Z�kEfc&��� ^�ǥ=�f�
p�v����q9NY
����RJ��*6�b���������YfYj�M�Q��6�ՙ����c靱j����[l��[Sy1�ٳm��>    n�}��W�C������z5w]�CZ�J�;u�iv��P�ݬij��ۻw��l�V��ـ���
zm�m�b��{�l���نhV��՛kV���   n�o�-iJI]���G�HT������J�����>|�5J��eo��M��[,�x�D�)7���Ӷ핥iq�W���oL�u��B���p}���Ւ�T�|VU�*�ViKf��aXp   �}��W�g�>�����*U��������`e{k�{��͵PϦ���馚ا�ϻ�}d�����m��P>���K�N�]7��_{�ڏf�QVp��UW�o��n����[di4,&٬Z�   1>}J�����_{	y��Ͼt�}�.����ޯ���}3S�_=�vҔ�j|��^�V���w|����2�k5h{+��A;[R�χ�{�J����}|��.ڦf���l�R�b��EiUc�  nw=���^�y��m��Gϊ���������y﯀�}j�����)����n���;�����[M�^�{�S͕�V��|���:Mm�����T��5C�C�i�N���M�Yk3l��f��ʱ7�  ��gpbU�ޯ����=t��r�窒��km����O���Wr���}K�44�w���*���G�_>}�J�j�_j�ﯬUm����o��z�"������P��髾{AL�h���+M6�[k`e|   ����(w}�}����ش��y�>�孷Z�}���� o9�������A���yx ��z�\�� �����ח���ե%U�Z��d�5-��   ��vn1�5�����W;��P�=��@=r��tH������4;�{;�֔�k����q��hw�n��4�W�mD-�ZSRl�B�e�    ��@�{�P:����Р�]Z)����n ���x�
����zֺw�{� +���t ia� (��zm
�2lƲ�4i��   G�:=�5���y�T�t���UL;ݡ�����J.����Tx�j�4u^��ꇭz��:��  @   ��R�Q�  �b` "����F��P�4ɦL��L��IQ�     ���J���      �"`T�G�4���Ѡ i R�S�d)��� ��y'�������i�'�Y�5_k��\���y��ebϝ�3�Ɯ��5ߟ�HBIs�7�aI	'BB���I	'� ���~�������ǒC�p�$���UQ?�I	'�H� 	I���?��wa�?�����'�?��������Xxa�2DH��tIvP<2k�'�M��xH����xI��K'|P42:,�.���X�@����:$.��40C�@ߊ�A�@���,�@���>,��B�<$5��!�����<$3�!�!�C�~,������]��҇��aHxa7���|Y:0.��x�xH#���!�%�@��׋!�	���C��d�����|$3
�B�,��e���P<2oŁ�|RQ�D�d�ɯ��d<0�e!��I�O��:2=,�����׊��`xd|P8$.�C�&�P�&�R���ђ�<2k�'���< >(.��D5��ߊC�A�d�vP< kŁ��)7����pH]�����R��<0ЗŁ��<2k�!ѐߊ�œ��Hxd5���O0�<0��Iѐ�,��C^,'��sŁ��`tdD�(�@��ޗ�(N�e��&�P<0ߋ'��'D�e'��R�xHoŁ���82e��!���9�����< kŐ��o�82x`>,��ؐ׊C�~(O	œ�,�`��xBke	�oŐ�|XlgFC8R��I80&�XHZY			�!!�e ��	!x�$<$	7℄�� >,	�	��xIkŐ!�	!� � ��@��d�<$�5�J@�I����@|P�: H]�����R7�� `���@|Y �	���BkŒtHH�`Hx@ �� ֋'Fh�< ׋!�$},�Iń!с�xB@׋!80 ��$�$!� ���@�� ]�$	�`@��!�H�HB� �(Be	!�C^,�O�&�YO���I|XB$]� O	�HHxBHo�$!�@|Y$�.� C�C0� kŐ!�$�����$�рB�BH�`Hx@�ߋ� �D!|Y!	b��XoŐ!�@|X:0�.�	�HMx�BZY$��� xBH�� ���@�� ׊B�$��Hxd >,&ĀI�`HxBBkŒHp@~)$����td�,�5��C�0�x`>,�e�ၯC�&�Y<0|P:aI�,<2o�'�M��x`�����xa�O7��▔�]��kŇ��Y<2>,�]�O��I�&ߋ'�G�c%�d�ɯ��`x@|Rt@�(k���'��Hx`;,�e��P<$7���|P: xL�``�׋�	��G��%�@�^,�~4O�K���ɮ�O��xd|Y:2]��tf�Y0dߊ�œ��d�^(�Þ,�>,�٪a<$ߊO	7ғ�G��.��������5(>�,^�1�5�8R!NH���ˏr���6�C���V�u,�4�
���R�!�P��O��-����A�srޜr��s��V�V��]�@ݲu�O'�{���tNYG+C��=;-�+e�r�ܹ��t�Zr�!Bfg��a��a�k<脑8����Ӗ��X%���f�����	e'$�3hӁnm��J�+1Z/�{r�')�h�:%i���`���ظ.=&�̠�f��)�@�{y5m�N͉-jK�8��b̈́�%?���ٛ�ZI]X֚����Y9z���� ,V�*Q�ч[-����w%ֆ7�F�1��jݦɱX�dU��/ܫ�/CR7�U�k�i� QZ,�w�y�����䩓;���P�t��pL��Ҭ��5j����K��/tR̚##v8�,�"����'��W�;İ74��r�$�����U�뽫�ǗF�J� ��*͋�R�m��%�	g�/qf���g�����U}Ǒ/�����3x��K�jB�T�sb�w�x��V��7�D�A5��E�xM��i�f�!���a-)�Ae�>Uu��[��n6Ĥ�JX��Ne0d�Zqޗte�n� �`m�*LJ�el#U#�F�z�=��v��ѹ�������hl�1zŒ�(ZءmV�^�,X�3Nk�_2��5+]jded�Y��]PQ�M!�4r�96*9�Am��"[���]k�oD�;�w�!���R7!��*��-�˭$B�,Fh\eft�����i�3r�Ve���(�u�۴Y���c��+R��*ЭźP	cO����M�6��u]����Z���.и���@C���� �sD�%\w�r܋ej�N�]�m�h:�xS4�#�k��@*у6�k��Ր�
�7q�ņ+f�u`m=T�1Ų¬ڼʷ�����"��>�f֪8Fmh�V!n����0aZyj�6��u%�4d7�J���\�̡NM��Y��w�J싸�b�&�;Ln)�V�97�+C�m�v�w�{���\��|����@WkB�6l"jk�i�V�����@Y��VeP��i�a�,j��C�-$�Qw�E�]��,�l�U,L�B+r��h��7T�Yt�zwp�]�)"��v�^5�u�T��\�1��Re�g	��*�'gB
�Q���ޮ|�$���˳j�Nit���ut0P2�mH3dҡ��b���8Z���� �u͊��Ğ��ַ�DTZ�т��дR��o4%Z�s"�2�-��$ �X$N;��QAapT���D�����*�n�,��"Sim-��͘�m&�KQe;�&�Ẑ�;��+���-���3)�.J�hn�ݛ�;ò*{��V
nQot�SZ�PREn���h�J�`�]K� @)wy]=.ޣ�ksX�)�˽�͢��(J�trK��GZ(�4�&��B���n���E7Ya��):_<�X4l�Z-��a9�*F��`Ϙ�+FPOqVٳ��D܏u�0�1n$G�p�[�����\[�c��{X�flY�_��u&vmi7R�`R�V0$%j�i� '5=.S�6�b��w�f�MX��)v��bbr'"��9FfI�6��W�5.��ؖ[V�X�f��R��D֑XJ��q3x^Poe�k {t1�z���d��Q�	��ˬ������ߛ�!�xH�F��r�|>�Χ�45�ԝ�4�\�dݩW1�Ih�U 偻2�f"�%�Z��6c���X�5e���&R �j�[	�b)���������rY�*��c
(�m�֕��i�-��uY![x�֤n�v#�`�.��6��e� ��LAhP�4L����y������׺x:��~ݚM��`����;��m��q�j�VRYu��Oe	�d��Øba���W�aӴF4Rq��Z���o�g[k	֞бK�]F�iF�=zwEGO2�pǆ���$Y���$���Y�I��He��v�������cM*���q�ڶ&Z�:���&Ķ�*
���V�a�!���7��Y��2Z�q��ؽ�D�����"�4e�è9�M�(%�<�eRܫ�+&�L�c,d�(m���U�`��,`�a�m�(�Vֻ�&Dj�R7����$FI!)b��DE��gs3i�.6�e�� C��Z��m5Xn��Hn�{{Z�i{v�e���v7P7�\����Uc#ka�f�u�^�ILeG��]�m1�LJ�L�kFؗZX�{\�Z�鏭�{�!�� ������n��wYW�-	��b��ȶ�y[���X3��·��Yf�!J��>��]�S�]DV ��=n����)�ra#f#�{��U�.�L�MP�Fb�n=v��H�Yj��=/����`PbfܖL��d�ތ0ܢ�Ńb�І��v0I[NV�l�4�4jmĦ�KRX7�u ��D�wʙ+6��
խRQ�	�{�v��4�.ژ�����؋S�w�4V��@M�N	�
jF p����ጊ�ΚÎn�Rj���.�2�P8Zq-����[&�d�3>Д@^�Kd�5���2��$fx�7S�KUu���B���c�J���9��|¶��ݝ��=��H��j��r�^:��K�F@�V.����\�xm���Ne [Tf�r�i4d#wm�.�<�e.7y�֒�i��l��{Թ�r_�m��Z��[�H�6mɃ�̗�����u��_��z4Ld�9�`VTT,�4D(�#X��Q��'�n��b�a�е���n��)��SqA��)������R�������D"#)��h��n������S�xl'>�p���v5�ا�3�NPYCm�*�U��ҏ�Yce�Ԋ�+є�M-�ŵ�Yjސ��������x
��ti�r^��tFf��̳�TƘ@���6��e=�0v&��B�k0î�q�����*��`�����3>&�����$�&�:}��+������*�پ���f��x��+P����VMɩhI�ŷp��Ҹq,ݭVE���-:lm�ut����[�cb�.ͽ��2�Tm����Z�i/TUv�/���xum�-\n���Y7cv�z�ϬL#4�[�Pu�܋>���+�N`n��Д`�:8q�0-��A�w*�3p�Q��w��i�&���-��.�Ѣ����h����4��\� �� �Z�Y�8���%�`���#%B;r�ŬPܬEw*�ܵ��]�!��l��ͳ�)f�t-��c��s�(��29��[Z�0�*�t0�Q˰kwk	��L��yى�����o�[�]  :�l-��zݵWR�4��m,x������̬�b���M2nݸ�]7���u-�F�h�77or���p�.�6hō劷VjH6�����u�7�ͼy��b���0���7��v�{�;�m�nⱄly���1!Ii�Ov�P������-���`lϤ�/U����3n�X��S�xFIz�t�Z��-5F3����~��j�'��s6��R�?{�D�\����ͼ�W�c[vU�Dd�T76������x��R�/b{a#GsON]=�����"�e\���[!SU�k4�g�z��<!�0��bS^h���𱷊Wpy�z��OuZ(�ʅ���^ ��ކ���
xiEF�TamG*�R@fÊ�2h��%�e�lM� �.��֩�4e����X��l�Q�

,��ѽ��`�5�;�7.�^�y
��Pܺ��5XE7OZT�r��akA�[,^"��h�J���+�f\"��/$�B��ڂ�1�(1�%7J����ӤfRJ�S�2̃K�О�ư�'+\�f�B�e?��3d���[8!�Mh��(2j�H��t�)8ͫ�F�b�L�z�V��	�5�fǸE�L&C��*�I©�B�a��5�mE�LXx�� ԦJ�᱀^�FRJ^&�e����(�~ԏЭ�wh7PX�r����E��0hh̨�v��#[��071��d�"A4$vݣdië�2e�j��u!�m�s(S�[�nKxD�[�6I6�F�Ѳ��Fb%2�+�iK`R}r��A,��e��w,Mp�SJ����J�/6Ȣ!��4��
dj�e0�n���A4�m�*[�4P�z��jU�T�5�s[�g��H`�y�s%0�Q�"�%7N[ ��۫u�ǡoۥ�����<t�ǒaͧ{C2Qb,��[p9����Y�Jו,�Al���W�saZ��{�^��P�y�yx�����kfn�N�`��D�[[O,>Y�H�,�0���������Xtlǩ�b:#ʷ���ʗ�)Mõ��q1��2潨0;�(�,-CV�vN��R�3L��+%�����R ĭ���,��Y3U�U��O��*$��i!+5E�'�#u&Mc�=�N��V�h�i7��p<�1n]�hm��_=8��h�J	���[V:N��-b
�
U�q,f�CA�)��Xj��	��Z��X�?!�Xu���u�ͧp�th�U�u�^�5�Db�h줌nXj�B��Bf�9<�S��s%
�c�W��&��GA~T7n+��i�!O	�Owbk�n��,/Q��6Ku*�n��-C�J�&!uy���$�N����oL�3j�Inڗ�cZ˳do�ކ��PH��x��Z����)Sͳ�� ����N�g6�T�7J*�Ջ�AEEXSq�i�����+�u������xnFw[�������ŷ�Vofh ѥH�����p�/1,�mN��u� �l�Ur���8Y�nU̘(�˙��ڐ�5u��UQV�S)TӏA�*^1i� �em�D��4���l�%(��Ӕ��4�f0JUD[ԝ�f�xm����[�ѫc�-�3Rcf��Au��z~őe��>��'��Yz�pn@v�8l�9o.�c�"�`��2sB�R*�	�d�l��cl�n])e?�ܬx�1r�E~�6+h7�5��Y��#�q��� ���X��A$��k8ҭL�B�55�&eH�)�43U��)鳐H\$Za��\�W ���茷s-��/�%�+j]5��2��j����V�	�<�a!����y�0cߑ��f�`4]��ѽ/s,[�.��3q�jʂ�-У�6*���m�cp��T��s2�=����-��P�c�©�ͬKFn��BB��� ��v�J2R�T&ҫL�n�)��E�e�WR���XG^�X��Tñ�[�۔Uen-�a�E��RY�A�[�C�ީ���n���7���
RS:&'�e�Y����%c��W�!��5�Ej�U�Z�/@)�kn�[�����Y�/Yw�0�h3.͛xv����.yhuуU�)�7�sV��`�]�n�tnj�j/�V�0Ez��6nb��!�k0ڧa�J
�Hk�s#�fg�t����V�&��[f�1���R��N9b���O�=����2_vܩ�kum21�Xt���N!�����C�a���g1aj�� ��32.�+Z����eK��spi#4a������j���ϑU���8��n�[�c��E]�%`-;�nΰSe+@fѫ���6�4�xh�Ufh'�)�Q��)GZ0mۢDa ���)(lGN
�R�2.�]�w���M��`��z��lV`yc�6�5��Ðَ�e��X����`����E��<V�Tj[oJM����8D��`n`qV��tA�/\ ]9��Xŀ'B�%�>�l�u�#3Kfv�I��7�9��#[x۫�C�Ǥwg>�@z���M�Ϻ�!g���ի6���F\ߕ�=iK�KskC�@>f��"ۼ��Yk�cf[&afȼw͚֊�lfX�AڌU`�V�D��[7/2�e��@(N�zE���C��),;��Y1˪�BU�t(7S{aPf�P:{t�U����9ukc$��+¡��
��0���y&��Mد�=��#�Ûu���b̩��A�mC�,$�z!z��aͼ���mIv�w5�:6q��q���x�4I��/&��{B�i�f��NB����)�CA �1=��:ɲ�8v�*��ѥ�ʟ��(E�Ƀ>έ[���&e7aĄ�pL܁ɕa$�0v�[;��5��SVŮ�XdyS����_#6�'m#(-5�\HpM�5���^����gUnͬ.�F2�<b�� �׆��n��r��h�K>ȵ���#�Ԥ����-}��ݱw#�G+3Z/-&��Z�v�!K#�6�B��:7�K���������J�e�����ݑ����b ɣ5,N��I�*�ـr��;4��Q!sf'�����'-����[��ʰiJ�$��ͨ�E�9�Yy���2�);����}o�VLZs����)Lt�J͐�W�Cbฟ���ɃF��6j�@�1�)� V�[����ʖ�7���@��iB;U��2�L�I3��!�
�L�!�Dڲ�2�K̗^<N�"��ƺ�mV9�(�lmd��ˠ�Ȯd�Ҍ��gj<��+L\:vh�ț��0��
#m
 �"'�8�-�ACW�U� �1^k�*ޒp��a;@��tW;�h�J�F�Tl�aݎ�3B�u؂�Q�|����KN�ء\ra�-N��v�M
Z���޻X���A.�k��i{{I��GPPh�!ݲ:�k�ڐ��ú��Xx,Z{
�>P�2��":U�zsp0��[k,:��%Ip醼Yf'*1VQ$:�1&����iD�J�3D!�De��0K�J�YJݵ�)�K��,����i�ƧI�
u-2�cZ�*����8�*��%�0>� �h�w�����> Z���h!���-BP�ӂ�{��6�����|c�l��g���_w�8O���G��|������g�֦�q�_���Wo%)�`$3_@�\V0Wm�'p�DƹG�P�я:q��7R	u�9D'�����֥jUʮ����֛Å��P��Ϫ4�p}�۠e̩�D`�ǣv��{�i_U�ȷj�*m��X2�W	��o�򬂢|�"�P��N�sn�bŗ%��Y�d�����:�V�sv��I%�:+a��Ў���X��6K�S�̆�����MIF6��;��L��c�wn��͕k,�U�՞r�h�3�j��p�g;jfX�7+��O�m۰m��V�Q�:�ժ��!v��s���vP�y&`9�H���m�:��g�ʃ2��L䂣��W\Xr^nԋk������w^��h铯�X#f���|%���%�]yi�L�o[��mgVP����Z�ϲ��Ѳ�\���u\{��n7[�8.���LZr��8gv�*Z#�I��[�;{n�D�!Q�kԑ{����I������:!�%I�@L̍b��
�L�8�S���
�Vb�j�/u1�����(1[eDOɇ[+~\�W]Q[#��ݘ2�j<���L�՛�G��3)��K��,����E�;S/u������y:3p�E9Z�"���Vg�FD�Ms�-��X;�=n��PNm�Z��6�vַ��˼���D;wB[��ӵu�j� �k��ܷsp�L� �V�f^B]\ϱ�ҳwr2�6�D�3�{�|�
(�U�ӦC�����ΰ�/�K�H*�	�[�(XB���ܺ�b��M쮠$�0t����kӀO�w�eB�%�7eS�$�ޅ�b6,��Rخ��+R��MU�+�VM�䡬�]�6e�ö9T���ø�=���M��c���n���t*������I�����2d]z>�]�]ޒ-�t�[�}V�M�tZ���鶲*���69Y�f'g)g�z��^��0��D2�z��4h��t��R��Nuu�8�mUվ��"�$E+��5u/�b��������s�+Yۨ7ۖy�nf��2��N,�s�`�m��u�+�O"H�,�qӭ,�,��ʛ��QZ=nEչ�:	-�i�u�v����[8GZŏ���s�1�ΤӘn�kl1)�T���1N��qA�ԓ�H�A�{]�T*-GV5�O*lrŭ'{jh�Ļh���_5x��Ar��f�o+�n�+JG�I�t�� ���`2s��D��8]dMm�zʫs��t��36K(�L=KE�#�$#B<�R�ݮ����U��`�����+���uoo/���M���wd���=w��ӌ�e�PX���퇶������h|`���z���x������W���%�j���.���wN$�6�C}�;�a�<�_bX��V��W��˭���=Pa˫��T��N�t����솦��	ԥJe���]��������X�ů�Iʗ.��:��F��\�ٶՄ��뚐�D�Rfe��/i[#>Gq���)xwޜ���ұ=GY���zZq�#$3��EӊL�ؤ�e�=��4=�;�n��%��%U�ۦhT���	��^tП{�l������\�6�s��X��h�`���}��z�\�o��ʁ��O1�n�F]7��]���sR��X!�� z�� ^J��]J)C��{k(�v!'+��ʼ����$���Ad����j˵wTw$��+)�j�Fn����lۺUo6��TrH�1�/����K�-�7�w���Y g�
��p��̘���fB,_p2���x�i]n����ٶI+�N�:J�cʫ��p�u�}���e���N&oJza��:�cN�$z��B�7��̼�VIP��S��Y.5�J���&���#��U k��>37P��z�Q��/�j��g�#`��8�,JoQM��<J�U��E�n�͵W���(�ɕ��tl�\9n�Z�㋽O;9V�Z���]�Yq>p�삦L�7�L�c+{@��[	��\�r0��KnV��[�X�q�0��Fg=}`��<V�(�ա�!�%P��|�7�Xηl�C[{[�8�]�4K�W+�~u7mM혯�},2��Gtr�m���m����Ɗ�P���y��vR�ѼxK}WE�k�Q��kr��-(�ѹG��J�a�[�Z=�/8j��fSͥ�0�+�[VmQ`��;f��J�E��%�D���y]�7�4,�6�Y�e���Ei�d��t;/nea %N7s��E>첀X�����R�<�-D�`���R��gk�/Z��[T�R�)���%t�nV�`}��XHNo;/]�ѧ�r�����̤u�����Q��ӑ�lv[�������h�J�Z���h+�v�ml��pB�+�^t=9S\�{�L�o��O U~^���`�\�2��,z�h���M~>o�N��J�>콲d%tLP�2�剺�D�gX��Y�%�.᜞'u�zԅT���H�7p����c]۵ر�ԥ�+�.p�:��ن�mdA�o�w�pF�4Q:���Eg�1Y��z�7�BT�ط�ʈ'���Di�c,u=��H��x�998�,��@��4�c��*Z{�.����a�V�"Pk38�u����4"��	�m�k+(>�4�FR�[f�N�f��f4aj�E4v�@�>�oL��J\�j��5��P�]'2�#���o�ձJ���+rB%�`���<��֌�ĥ��J�����T�r�҄^����ua`�qi�,ղ.��Gn�U+�}���f��X�����]��ُ��]�x<�2.2�b���d�dP��II@�*����@�9��㯲	��;Qk��{�h`ۮ����P���>��������B�XkG-zz�eE��܎�\�උ�]�otl,��Y��cr7W������?* ��S�r|��n®j.f�{�1fM�/j�:�`9�Ѝ�ڃ�nw51	�Z1O.�� i�s1# �H�;u�n����'��12��6u=Z1A��:z���O�en�����p7ʯ>7�{��⵺/���f,���w��.pM(D�3�Q؜�OE'b8����h=Q�/ "ʘ�4�擮�?(�����j��j3G�:��N�H))b-��p�}��SQ���D��s���$FU�4uv��.j�6��kNϡ��Hju��s��=Yʔ�>7� ��M���S�m��=�y�v���)���bW�� 2��ՙ�1�ڣ@�zh��7�MTDvJ]X�Ǩ���\�6���P�)��&����*�e�a@/:���G�x�U��
�2��[�RY���oTx́�ɽ�D�;���z��OOD9�M��o&���)�WY���kH��� V.U��%�u���hBG։�̻�� �E��5f�V���H]Z���Ss���ʅڍ�LPJ�M����!2�	���£�yعiJf��v{;��Ʃ��@�*V�w��X���.�sr�r����y�\O$N�[j�t���k��5mǿU]�b;yT����Nwn	�m8�a�.�[�S�͖���{&j�L>
:|�$�C(^�Gr�lL)%�����LQ�ym�WE`Vd�ufkM����3g�g�%��*g��K*h!��Pj�4*�5k3�v���w.���[�bu+Q/���2�}����ʛG3C�U+�C�K8�(��/�v6�u�Ү�]��	�J��w����=6=�u>��)9��,�נ�� ��A쬾M�D���Y�-���+w�a�W�b�{��6�yhE�]�X����-�ʶs��hp���&��Ҷ��S]���)�45���^�<ޥhu�MmX纕�Z��-�'�g1���bܲ���ѫ�0��L�Ҩ{��:�V��3E�m����hP����Y�7K��:e����� ���y�ݲ�6ӎJ3�d����,�,�اD":M����Ϸ_.N�f�ޝ�B������*զ��N��*7L�"ЈmR>�3��⽺;�wu"(��cd�ZkX��=�q*a�{�f�ò4n�9&�sm��cA�W�1Y�y�*c.��+��;wJ%���9�x2_eH(N�ZR��^�ɥ!p��XH��ai��h�b��.����yn��D��U�hv^�qYAu�4��Ŭײ�0KaSޮP��:�D�L�{dEE�2,USi ܻ"n���۱�1��I��a�,32��Uؘ*���F���
�۬o����il���l;˽��+Z�ռ���Xj ,jd�_�ú��Z�d�f�5$zneD�u_8F��Ĭ�W_-b��+�F�X�낛�S7-e��dQ�k�U[��2����H��ٸ��[��V��"Z��BiF=?F(����s*^>��s���y2.���{��ah_4�����0�u�`V��7c�D$=疝Z�3���23��˙����nP�΀�]P�l�Q6pr��K�콒�֦cPԛ1�՗����,��u��675ͮ&�kL�,늎_SO��!���O���\Yޚ���php���ﶸ*�K(�媙�u��ܫ0nF����^$�K�.�F�٪�>ˈ�|�&�BA��Tڂ�ۋXwd��'ٕ�Y����Ԩ3ac2��>*m�i]�[]�:.�IvO��xh����%"�|6���zSx��S:�UQ�Ut�ct�Z����K�h��ݗ�R�m ���h���f�ι��T��F��V�����ۜ3Z��=���/r�uk/ 81�wtڶ�(2�&�!�b�)������L�/i��s*n�&�s٢G/6(LVn<"s����k4X�a�Ʋ� ��)��KP��̮���Y��Dѧ��̓!�Z��C������s
��J� x��r����, �Zm҇�nf�E�m�^����/��ϻ�(:k ܹj�ډ�J�nS����t�;�v��͜���Z��c�W/��_r��|�<�ۚ�5��h�v�n�vjݙG%�|��ξpm�;�L��-D4�B��� ggt�ؕ��0V+`�j��{,;W�����k�GU�ʀ�[��У���k3mTB������}7S�s��Y��1@�3�v\�Z;3JҿB�.&���C��O���'q�7)�\ھ�p�Y���?����
̻�w9C
C�.�9����<�����X{�uri��;�Y/o�;�8��y�W�B#fҖXS�E0�t�����6A�2@�QV���3�rk���"t�7�S���YA��JG����3,�ŕ�ms؋Ohe+�+�?�>�,�q`���7gX2�D�{��#�*�V{�(#߻4���pE=[��2��h��\���fve �Z�nͺ(&L��	DoSꘃ�sl"d��n^9�L�r��L���L�P�7��l���փyØ�d��v�5�OhY#ٻ|{�+;�H�V7��6f�#u����Yo�G��6�b�E�����c[:ѡϠ�ZV^-�whg���[�:��O{0C��^M5I{���+�>b��o��v_ML�6��
q絸�.H%��8ÍRZ`mJ'"N��7tT�Ր�w�a���/����m��6n��ko���:���xW3�,��tZ�#MjR���q�U��+f�>�0��u����/N���w��y�;�S�O+w��XW�������lJ�����t榔��ь�+Ty]�6.��cgm����U���V�8o> W^���V�����R����ܾ�c�v@L��Y��m��a]٤@H5|f�%e�-u,mf�^wgJ �6�l�6�fG�%2$�c\J�>s11C����g�F�Uh�Y\�$:_�uu��K�����t���3f�`짴3S�`�yӃx�R�Ŗ&f����>����dVŧx��8/���b���M���U��tՌ��@�f�T��oP�#�_Fkeՙ���h:��QZ�h7����E�AS�V#/{n,�?P!���ov_C��ɡk�;Cm&ΐ��x�ʝ3hW�yp��]��{h$���KĦ�K�Ko�`m���5�7o�Y�Y6^���[�bֈ�2;u]h��D��M�Xna�e�XK�a������<�ۻ�&ڵ;c�G�t]n(��
���}T)�*:�.�m[����2ݙ��Pj��F�(�>�}&���wZ��t�����]�=��c�
\r���%Z��[X�r����/��_o&�fE0��:pg���,s$�[�eqk�:�S{!&�:Ap�:��ٵ#/_M �ܤX��N�7�!�f���f���3I��Fw*I:�[|�dV�y�6#�n_U�c��:'�7�Wgsky�m��/En��F��tJ]�Pڼ�'qe�j�nu^��Y�s	N�uf�w�h��-u��T�¹�q�j�k�֞����M���E��aX/4�����Ad��(��d1�Q�4ݺd�i�L�B`�jwn�qGx5�?xu�F�5��W���\�8�w�Ҕu��fk2�ET�+ʴ���.J�l�č�'�0��0e�9,�!H#D��2XJ ]Ug���Ő�A%G���L_�BZZ�"�[�ȑ��b=��l��Cl4�9�m_;sG��B
M�a6�J �QWz�
J�9ѓf���%�qmS�G��(*9T t���L��L�U�L[�̎��ҪD&h4���H�M��IQ��Y`đ!�I���K�u���m��"n��*��[Ka�)ˁTH�d�q	TEFS"���m��h"ֱU��ZN�$��6+ıC�/��<�!Yv�$�$�~ME�Z4���i��2	�F2\"�H�B�������C����QE2��T�U���*�}��H4�GYm/G��Q	�jC:&�NL@�_�31'�?a��� �I �s���6H�>B ������@fw����_K�����2�'��P=����}kZۡF+W-f��=�ӯI��s��-ŵ��t�����N��r�̏r�����o.��BW�y�N0��;A�oEM;�;�����S�huv��=53@�Kh���ܬR�Cu`ě)*��m8�����h�S�DkH��nr���R�2��Rʅ���e+��>�Nf>ɂ��Ɗ��F�U���I���Z�y{�e�ӝin�N� �U�@�f��4�n��C�1e`/�rj|�m���f޾jw�~I�".�-6���
g3��� �9��<Κ����eıu���Z57a�uZ+s.�A(�i���ʋ-Z����X��"�k.�.��뵺8�W�q�u�'d&�g���#r)M���d�sf��۲���$U�Աʝ��Q����\=2�r�Z�V��9���v4��a�F]��(k��y���;�Lv3k+T���ߢD�P��ú��<�m�"�N�#۟�%�pQ����/^v�mF��L��5B0\�Pi����w�T�x�5Am��[��jt�]�>�	�ֻd]�4jV�k�)]O!�S	Q��a����^��&GSj��h���_.���
.��!)��0r���*�#�#���\/�m���盡��޼����SV���D���Qp�&�V�ɭ������j��6666664�c��������c�������M����6q���������1��=��ɒ�ę��݉O{:��f56S�N6�&X���f�
�Jd�aǜ��,��O�M��5t�lĕ���R�����n�䡈�8�c�p+���z
�pf[�vq�/5!���k��9,����I�Kf]^�#5�Rzq�v�T4e,����S��M���Jx��)2fP���>�sy��V�]pJgq�!8yn�t��ԙ����U_V:Xxov�q:`,@��X6�()�5r���
�*�z;��5�
�U�̧��R�g^�Q�`�vb���-��c��q|��vJ�Y�K�f�*u�}׭<�2e�j��h(�_ĳ���qj<���HA`u�ui��6�;��E��5����fiU�*�3yG/�;br���KV��l���\���k{oh쾕&�,$�[��K��FU�n�,�1�n�0�Ģ��,�9�W���@��O�N�c�/�k�6�h�U'd�1��z�Z1pɟ��)�8F^ҳi�����x�z���x���ћ�&P�Tg6޹>wŋ8�]����N�큅�Vۻ�6�[;7���lGW�d6�9����3��́Ju��O==���|:�d��6d֝��U�;+�EpL�ۆ
�s��sO	M�z�-
��+���V]����<��	lllllla��c���������C�����4446662��ύ��������1��cccccE.Q>��J��A����[��;T�ne�it�����9t�.�p�ܬ(���4��і���;ǀo`�#ux-���
�k~�ùQ3s:Br� ��&�����z���nFq�Ղ��'�jt��v�:u̝1j�w�;A{�\�Ҹ��y��DiA���������s3�hK?�j���ѣr��N&x\�oJ=��[0E�����ǹ����e�����is��/���Ӏ��W��V<�!*mIB���s�&�����9ɳ1>��E�dZd|���d��'D`�;OA�c�ف=������i�T]�b�V!�qRh�\�;	r�rف^����[t�_�tL��[��ei���څ0ys���;�����p��P��jΛ�&M�!F�+U8�9��u@���ݤ�^�|�I�d���wcv˕����2[���n:�G��oi�º�kݡ�Km���_>r\¡'80�r�en6��:w�`	�%�ξ,��F2��c�V����%�;�f�V8r�9��r���h��2����xD��gՠ+N�:O^�M�F���vb���T�pL�dzK��`�plw!��a�5ŗSx�n�QJA2�6����H��'�̔ ��쏟5�N����숊,��o�������klq��������663�ccc`@�Kcle���pű����cccc`��M������ፍ�� cccc`+sB8Qt6��VX���݌#,��)�X[@r2Y[_UP���)��{�Y�y�Yu���%�x�p���	��_io*ډX��Err!��{��l�c`���T�ʌh��0�m�9�	4�&3֪v��A�;5�v�m)6����sn�]�^՜��`h��{���i�X(p��p�E�k'���I.�r�f��qFm�dY�Ψ��w18�Iy]I.�&�T&�ɺxw*���X���̢]��∽4�9^��Fa�a����	k�V����UTV��v&�T�6�N�[k��X��],%i\%���R>m��� Y*�:���d좺�mK69��͛4=�$�dՂ*$[wX��@��*��
�t���Qy�[��D����M�8+IV�jdZ��PP>B�'E�������P�I���P��aeQY��)�N���i0B�-��Y<SBN�����9��<1��Ћ��Ko:��fKm�]檹��z�m�a����e����f2gF�8j�F5ʩZt���u"����ʔ�>�	��p�kz���ٗa�f�l�0h�`�F��)�k:VXO�^�-��i���l
	�G+�iuX���mw-��%��;`.�m��,�jc��^ͩ�TA==H�{��K;y������llhla������N66460���ƌo7�� ccccc`�8����l�ccccc`�q�������Y�TVL�9�\Ҟ���B8d���߿7p�͕uB�4�[lue�u�m=s���7m��r���Z�`�&���&��[�Ž����(c��ܡR�y�*�P�ל�a|�9��vJ@��k��lj4(�3h��*�o5HpL\������:Ɩ���4�u޻�к���}B�wN'y��}AhF��:$�V�]z�f�\�� Wgg7����Dgq6�^���,�38vgF��
��l�o~�(WQ8�V^W�Z�f��������ub��]�%�,�[J攅�͹�5�V�C+ED����\��}�5ץDh����#׌P�6N��V�L�o&����k4�R^+ζV�<���e��g�꼤��ְ���58�/T����J<�Z��[���n�B�X=Aj��Q)w���0MҸ�\�g$!R�7.ŗA}�HXا�SǸi����4���¹W�ԉ+����|��'kd�;�&�����R�r|�^V1�M6Ѿ&�[�{j����Գ+2\�J�?}t��G�} 4:��
kk^ib�5��t�	�V�n�i��oƻFٗ���T���$������ƍ>+$�Yt֚Geȷ�j�'=/�68ɜgE�Ѥ��D�����eNHS�ޠx���7.�ʹ4Jy[�d�9Jۉh��#f �
(h�F�8p�Æ�8!Ç8p�Á8p��@�8p����Ç8pᣁ8p�tA�+�����sV9}#h��95pާ}��8^�UAq^*@�pL?;K��Ș+��oz�~Sx��Ŏo7Z{G	/rjڢ��Dq]��fM[Sx�
�޺hf�p_%ek�+l�8Ӈf�Ϭi�m���T.	�
����{'6��سnk��8��V�Y�$��NWh{�3s�w|�uV��;8�k�o0�XJ����Q!ݸ���Hct�i���G�z�a)�.��Vd[�3`i��)�s��^��� ��E+��]�=�P�չP|_s���xT��H�V�e|�mݰ��t�
���FD�6��ڞ%�WF(@hX�׼�h�T���^fZd#���$�Y+�Zu�Vr�ka�2�}��R�����o7S�v�7uyr�Z[gR��\�/�ٽteқ��Y��1�����jc��<̮�;�`;���YK�zwY@��Ѩ;L)�N��ћThwU�P:�EV����؎�`���O�����R��ڤ�%k_}n����	�J)��޾�RPv�в^�o�\9�tT��5:�sĂ�T�:X=�S�1������5�2�TG���Sh�N�U���oYԶ)��	��C=O): ^G.��+��\�8��cל/��4�QRM�XSB���[f��F���"�ư��h��D9T{z��<�'-��+��[�N�J�b�p�Ç0p�Ã8p�Å�8!Ä1�8p�Ç0p��8p�Ç8B)�&�׼4Р�vnve֊v�2�4�f�eŲ�wS�]�g-��\+c�zl \�Վ��'��hU�F-Å�Y�.S�	C�Y��c.�ڴ����5��])�&� p+�'4*m���ܖ��4�;f vU��	��U[��W]..Dp�:���P�g#9�7��OP�8W��ưDE�Y��^��[��vnʳV%�Ȉ!q�|��	55����"��]�h6�36���	E�)�uw!�����'x�mȉ�:x/Ѹ�9�{B�xd���*��k��E`L���@�q��w�;·D��'zo��	N��_io�vw<Ox�:VZ=u4�|�F��emMH��.��m)z-������cX�J���
�oBf�P�lM�2�dh�zrr[6��(��{t�s�q
�Wh�B~���)������2��`]3��l��
�d��[fm�>�>������mɴ�&����L<���Tpܼ�fJZ��h��o9�;_.��]����7�%���si[ՙ/��ϊn�w��mC*�th���5�䌵��r�m�W�\��Uk�fȲ3+�6tMj�Qѩ����.���յrY�+����A��3R�J�׎H�i܌u���"���6�����쉪n=A�w�.lٛ�T��*���U�v3;�?��s��8hv�[���ń,X�F� �Ç8p�Ä8p�81� c��Ç8p�À�Ç8p�Ç8p�.�WG[��:陝�]��!Eǰ�� ��X"���Yk��:(^eA��`�N�e�:��F�B�(�\n��8�]��.�e�S$���V��4ʪ�� :�W��tc|�ِ� &�1ue�[�+s���H��6�۠��6&*y��#PR���l[n-]�_-�,�]vyh�f0k��YqA��c�ӮiV�bW6�Zb�V�X�*E�&�ª�{A�YP���ɟe[m
o*Z2�׸�� � 8'h�L����)���]�t;)�I���#�T������v����/38���dyu4Q��Sd�ǔk�r�+�j,�̏�WG;4���6G}�̶���� %�m�1�g�Ԇ��]���y3^�� ��o�ň�3o.a섃�X�����ԏph�������umn�X8SΔs�r���m�#M�		��Ǚ�ػ�s��4����;7��F�3���2�8�T�݄v��rU�,�[ћ�}ikF��F��ގ�	�f���J�
����Y����UN�����l�={˹+㛗B:�H��\�R�̈��2o�{5�!�FU}R�	�5�,AY�3���4��W;�=㐉��P�{BK�T�&]�B��6#��޼�t�\ӬVjf���ƺ���}�����/�Βcy�vJ=�ͩpY���!=�K=�w)<�RI��v�6�h"�,pᣇ8p��8p�8AÇ � �8p�Ç8p�8p�Ç8p�Ç8e�ٶ6��7k���E@3\���+�B�����*�^���9�`��Z�U���0�1-�Ft�Ď�:�8�V�x��I��m�a�U�� =�`�s��\Lum�y����|5qZ�nإ���P0�m�?�"��>��R�ɻ�)r���G����-�'����밮S��Lܗ"��"��@W, s W9s<-�)8�%��D��:��x�]�<����L�f�xl�b�KUږ/5��e	 B�v�>Ҫ��WՒ�'3��_�����P��՜
����d#e΀���{L]|�=F�A�sf�1sڗ%�݉�v������]�.��}nʜ����k*s��q��ڇ{��nP�A�\�����{!��1��IF���Z��tճ�t�}\�n�E$1�̻��Γ����Z��Vu�ϸ7���|n����@�7)l�[6Ѵ �'��6��)G�J��J{�܆�a�8��dOW�Xt	2�J�m�7�aqn^�Nj�����jm�br}_M�i���9�;��0'edB�2
�+3a'~}n�nI�=�,Ü�c&'eE̳���r���9h�-pm(����L0L;�"�%���
�7oc�����+�YjV���:t|-�����fnV�Iw0��q'�uҼN�W�T��Sq��;�h-�C��+D,tý��Qj��ٻ�[���]!�6AmeF>����**���r�o{���g@@��M8����Ħ�����ked�j�_}X�GՀ,G��������Վs�!T����+�V�F��Ft߳��kH���W��˅N���݆9F�vY�E�������W�*�JW�6�������+�t�`��>�p0{����0�5�5���Yъ.�]c�F�P���7�*�p�h��t\�%о6%A�����Y�MJ�q?c�L7	�v�9S	�S�>�k$���{Fɭ�sX�2]�MR9q�Ѹ2�=��4ͫHf��$���V9ҴN&�y�Ż�<�T���1
��5tKT��Ãv
�X����%�¬v;Wl��O]n`m�ތ
��WfZ�H{��d"��椵�n�z6�32�KBB�F�t�n�E�p�[W�q
��٤�K��ݥ�����gaQ��^YU�Sͭ�me��┶~4��QGb����EG��D�ᶸ�����g�Q]շ뼂�(��'Fm(0���D"���d�v֝�(A�}/XiV�ܖ�NK���%J�0o)�w�w+�G��
���uR�3�
���*����l�/��f�`��jղ�Pl»;$��م5i�tɮQ��]�8M��Hf����Ru��q���];a�
USJ{QTNw-�m�-�9�)�W2\�ri�.��|̙���ͭ�����G�u'.��0�T�/�����L1=�.�I���!K��eW����?�`�37�3����~ɟ���3/�����~D\��@�H�OȚ(��Y(�Wԟ�O�ov_��m����㴩�*$&�v^��k[+���,n�����M�Nͼ�i�L�Y��VPEnlY� �K��]����aŻ�	ǗP�^i�͒����i�b�"��%wV���3�ݝ��X[2���@[����;�kC(�:رQW`�H�Md��Ϣ�p��.p�G%���&���P�3j�]�>�n�z�o.�C;�-��V��e1����w�f��ޅWY��fAGtw m�I�Ε:41��T:��ܘ]���g:�QAS�Y|��@F�8�:'/������es�[.b�:�h��F,3G�WhQy���oM�D��x"{:�S�\t�OF�ۋ3mcwgk%IF@�Y�O��m[n�];	�/#�!o���'FVY���6rPb��,+{�#"�eˡ֠��8��fn�Vx��eL�`���f,!�.�[%�r�>��i-Mqu�e�e�������C��E�t'(��]�y��՛R�+��v�h2�b�.4(���}G+�e�}� ��W�(k�ܬ�=m���`�s����.޺�$��@�:.�X�$p�3r��
�z���!�n��mr��dW�V��k��Ѿ��m�vd]�pXh!��H�S.e��'ФRC�r��."qH E��i��!��.�H�[h�/�7)DO �@P�2%h�д�[p2
�D2]���0���8&��R�sMU�Q.�EUbGz0ִ֦
�ĭQE]%eh(�E-k����CVd�������w�eu�[Qq^��L�Ւ��֣�r�Q��34����**+�бk6�Z���2��N��NN%�f*&5�&YF�+)b**,*���)�,R��)��E�������d�����qx��i�TQ���^[�f���WY�P���Q�U5J�.Xڎ�DD]X�ʹfL�����zv���0���2��؎�1��b���2�C,��T�я-c6�M�UQݦ�kuq�m]��p�5SE<x��l8V����̵����s�,E�f\����`��n��F\ͺ+uec5r�"w3r����WP5�V�(�8t��\�lg/UdݗT���\M&�.��+�ʂ2�Fcp��˙*�[m��2�D��.V���f��2����q*���憄1qL4x���f�0I��V�K/u���J�.!���a���R��m+�r�e\$Kj[Ne3.e��l���*2�╢���Zd���[eMe���c�-�f�;9��X�ԣ1�2��^fLb�z�5u��U*��H-��uf��R���dE�yn54]
&6�[n%o.*�:k�uK��L��D��Y"9�`�������S2�q��k��t�f���KX�P��kJj�r�̼0��Kr�b�`���ƦEt�Nj޻��o���W�x����{|�a�:��uc���U�{�p4%"��^t�V�4�r��6��y�ZcJ��	jB�j��8@� 7�Γ�sH���������7����8&W��K��E���O�;`��ڱ����mV����������uW��;�ׂ~&?�}��z�b^],�<��O%K&\�z��k�{�K#�j�*(d�B�ʩlט�r�L��}&��w[�C]��KQ�r�t{_�\��L���{���p��z)�y�w���������߬��
����Ϻ�+���,�**��]qO�Ln�+��ll׽�|b�ъ��u�m~}���C�~c��:��h�LT�g$7^�o���Ĵ�:�������\X9�Kj�z�t� �Z��<K�רe���2`�<�������w���]�t=:�(aT���^�y�FN9^�i{���.��D_�`�}>�o�ײeV��vZ��aI���3S�e1¤9şo@�O���@ͪ�{۸���?JfM�׫��A��c�X�8�Y�Ԣ��|�����IЗu��\�x^�=�e���Xb��i��a���
�^��$�[^�Jn��=黠���&΋��T|w`);�F�y�ce9P㾸�x�lͱ3��Y�O\�)	@!wp�H�n�LZ��A�6�┪�4>�����޾��Q*�.kr�l�1��a�jy�ۂ�����<V'����P�o�+��UvLu�)�Ϩ#6��f�h�ʼ��"�.{��<<�ۦ�p{��:~=@�1��h{�^�lz'��gR�I�������Uo�ۼ�ⵌ�;�-VW{��|&߶e��������{�˘Vǳ�B����E߫_�;�F�Uƚf�{��4Q��y��Q�յ}=C<����mW���W�ʇxc�ލ�ëik�=�u�I���)����	����51�t��1�$Q��`u��{<�/b�㒬M1o���q.��Ly6 ���=���;���wֽ~9�'T�&/}3�uylqg/{�uO%�U���~ӣ���'�g�~����Oҧ��1�*o�*��^���^u\�ǖ����MPt�~/�ik�7y\�:!�!���uYͳ�$9;л,R�t�r���*������^�ʨn'�n�B����z	�#sc�[���s���e�
��gj�W0t��W���ض��Y.�� .�[�p<}���]�Lg�^^�s/�۷���N�y��4�?rs��5�%��n0�z��;��:�m滣�jw�v�J7�����~�1�6J�[�Ǟ<E�sV�2�����Ý��aN{�M�V问t;�	�b�q�R�:�;���]���+f�z�|�\�H/1�<h�|�+�B]=���f�`T*�|�m���1���3_5�
��/ejn=�]1.6���{����;��W݂­�b�(���ݳ�b�!�����;	t[�1'��6w�7ȩP���UnZ�����T~��b�(�i��)I�'�Jj���S���*fͷ�kje���[g���Omf�>~p90*>�
9zo�g�-��{���׾i��3���^
�G=� <���&1k�,��φVE��ΪV�����~t=��}Ru�r�}��$T�{���ۿ|����*�N�Ҹ��O��8/b3g���{l���-ö���h�|;7}�_W�N]�꫚h��':����Q�����v$7�ՠ��v�s&mG'h �H>���WYt�.��Ҙ�	�[�}�JR���N̏:"�5�{�5��e	��3VG]�[�0����ƴi���PU�d�}n\ҘH��p����w��)�6� {�*��6��t���5Wĳ\E��f�ďI�79@i�;�}�f��:I\��S�ꪼ�K�)��{W|7�{�g�<[����|��h�^yw^��|��l�e�k��{^�[~=�+��n���!�	�Ou�sF��H=��~tEP
{U<���e͑X_����h�G=C���v�m6�e���o�z��}�e�%�L�&���=[;�v��l�ݵ�����eMV:�G�O�q�����o��~`������~ͯ9�ꭣ^�%�nzOIy2>��K�āF���:_��^��fp�a�޽�s!+po��JfP�G��g���k�����=��0����5AV�Dѭ�������E���o�^����y� h�K����d��G��9ny��F�s�a�GuWK0.#�s����ʹx���G�!L�W�P����`_Jŕ���"�TrG"W����n���7�%�9^���nڛhu�S_^�s�*S��s����ݺc3�wdG)�|�c�g��j���w��L=g�Gs76�%;(�!��ڒI�S���[�g�?������].���A�Zơ���Ws��4�1և7��ɧQ�˚�n��ro��~t���;ɇ�҄ e�{��Vm^���/RI�IΥ����⬊voӪ��Ss�n׆b�Vi���K��,u7^y��8I[3k�e���;5=�����]�]Vf��@�햞�1��S�+O�^DݵW���`��A�h�"�~	ݣ���{��- C��w�wZ��|:Cڷ+u�a����<���E�����+6J3'�<Y����ן���3��v�[������!cݿ4�>����>*���lXu<ZBW{o޹٧�z+�����j���������W]n�{�rmA�9f��9�i���t}��k��5m���{�N7�'FWEnS״V�"����6�ڟ���1c>��8��Md�o�k��+��^�����̭�O�Ю�.���U[;]�~~x�5��8}�A�Զ��%�SC~��-���Z��_���bAQ��/uh\�\GbS�^o.�Uoы���{L�O�EN�/e�Z
�m�필_m�����|+WS !�H�xi�V�ێ��5K,���;N���w-�M�y#7�3Op�=�x�v��|�������Ow����o3W���e�����wz6����_���ܑ���sfF>�v����������}v4vk	�����=+����9`�w��b���%�[~��~�]�TfB���8s��P/w�<�/K9ר����[�?	���g�y�{~3��Rі�T7޺U��xa������=�5S�a����+2VR_]����Χ:���)
�O}�n5���-J�h��)��U`�2
1�9p�CZ�0חB1�E�M��D=�?V�ހ	�bɽ��~�o8��l^x�c@���Ŀd���B5�4&ߘ�����=������~��{Xǰ�o�s���M/�b����6�ó��ǖHGn�aF}{4n�kFA��Cܚ��O�mJ�~�r�yA���|��Z�ۏ��m:r�w��-��5�X�)L�ճ}�N;�c�#u����S	�#|��F���0V:��ȜŢ�ܥU���&���)(��˗�(��9ZdS-u-��|��ԭPՙ���%��Hu�l�)�mm��r�RM�S#���Md���3�dT;���g}��[�k��y�Y�C�w�:3~Y]�Ew5=^�t����7���Ψ뻮qڠ��ޯ"�)����O3�� z���	=��*��7�C�d?�����Sв#c|<�^Mma�&��>��-z�����g��{�'����'7��O���9+~�������^�; �~�t�P"Aʾ{���z�a�@���{M�����x�m/y�/��à��U���|5�^`(~�r�;�����\�(�ٴӻv�L��;$�w���m,��l�y����M��k�|�xE���=��*�y��z	��Cԁ��=��ʡ� _z/�]_��=k=ȱ���������~�������b�(҈�3Er����E��5>��)�Vz������f�F�Ln�؊��6�b݊�,p�N�*_��u���TZ����ߖu�0(��O<��r��v]��7o����AB�.o�hZR�X��̮�t��e�#�QN���Wq�IP�4��>ꋖ���TV��h�K�#Q �/@4.��[n�L�q�g"�k\���q]�)���1�
%�r�t<Ȅ%|�M6�Z�n���m2���Q�v�r�ϩƶf���U��2�Z�VJ����\�us���C單���T�Ϻ�O�t]�^Ӗ~�oX�~b�,��N`&XɷS��[�-`T����^�.�8K�U;�~G��U�ٯ�qs��y���M�3��t��C}V���f����tײ�o,,�'"���	P�z*7`V���K�J�3�FQʱ�՞��p�G���}y��4�n�^�3���㫾������j�u��-֒�{x��,��=�7O�.5��A�MF\�,�ӕ7�w�?l�da�$
x��^�����U�i�.Y��7�hX�1��=���ˎ�C}�����D7�\<���9��HiW�����^fQ��>K�����٥^�ؓ�p���T�+٤��^q=픸���p^���]1���!3p�{*�p���[�S��#�7xy�Y�����.]�k���_ȱI��)%�IW�������շ[v�W'dM��w{�9�Ǡ\��2�oLk�d��jW9\��mq|�Nb�߮��[�d��jU��0���h�ћXE!�)#"��T(U�����8 e~������5N�}��&ۋ�|��{��f�3�}�|tY���7V�!��E�Ӽ���~7�j2�4*�^E����y�΋�'[�ѻ��>yr�������/�D�z���z���k�M�.��u�����lת���C�f�۾�
2��z3��|"�����[�{8��^��;��^��x��}��Sށ�1�{7�Q������2�o�phN^�����m��K�,y�2��.�G�E٭'8@j͉��o:�x.�����`��w�L�6'�s-��}Uf:��.g�����@Սk�M.��2���$�.bVҒ�Om?hhY���,�Ŭ팓W�u�}P~���k71|���{'����
���z�wמ�*�0�	ŗ}��]+�=�Vo_��%,���n{���~��u=2���g�O]63;��L^o��ֲ�4��6�eւ��K����*L����5�:��p����.�~�+zYuÈap�W��y����j�}T�m��{�.�}����_c�
ȸ�� �Uڐ8(N=�w���;/1Ι�8�OnU�Yd˕�W�蹍*�,Zr��[����(��a��N�G����������L���t��fw6c9��B{��H
���whH��G|�����u,�W��gb�e6�X&������y��2��RO;�8=�}@�^�w�s�s��{=�bt������<���ٯ{����82S��A��{���q�������My{�+,�N��?uA�w�mmOyI7�7��;��- ��ڛ�=NU��z��W��R�ޏ�M������]'K*�Y�7��W�<1�� �5棾	tf�2�F���;�u�9�T�Xcɝȡ��&���TN��"����A�P/v�/O0Ϲ��-g���q�#ܬ�jߥbeK�o�AS�+���쨽�w:�frd��U����?F�-�I�H�^��yoo��kj�ࡣ%��VC0�7�v�;Ј���G�T�S)?������vSR��w����j��5���K��L�,p��(2�{���4�"pU-��7�a���l�z������`Xu��Ϟ.mZ.��C���j4v�UN1��
t�oh���Cg[�6i�3�bU6�dX��+t�ȸ�J�J^P�F	��D�M\��(����'��w2��gue.��������+�8��;����V�53UoFO�8f˘���b��ݙ�0�V��|r��ظ
Uj��ñ{��r
��\v$W�&J��:[sҪ��+(�e�TgL��Z�0�,��#��o��9A%p�m��i�t�vu��ݭ��$���V���wf휷�م�(���_t���In=�M��G=C��kd��Py2:yJ��ͧ�:������=�gV]�a���T��)�/�*3�D5dt�*!��i��U�<<�ꏉ@)��7���t�\�ٛ�bչ6��h6lh ��y-�p@�ڇF��4���E�H*�喺3W��y,�ʮ_3w�����n�2�awk���_;��v1Rp�_=�SC�-�ŗC���1<+6$4���>��8��j�Y��]�3dŷA������d?l���}�dj��G�
�BՍ�:�RS� �r�+�T�|E3;%๽[�����qY�]��[sU�8���5��7A�����t�dX;��g:�`��6Y�QN����`$d��Vu�{����-5ZyE���'t&,"��f�U J��+�f�\��buȊ��zفU?���]��oUN�|IqĤ:��b[���	�ӷt�M�ߺ��yL٨�c����U�$��k1E$}#vEq�މ���C���n�4Hx|�T	��I@�1�d�S�k���j۠!�yKwf^��"?=��$u��+�:Ǩ�3#D>�]�N���~�/�I��byRL����sw7���Z��r�Y��1��$���N�-T[\C�.�=�L�f
u��4u���S��ĥ�Y��w�0`���:V�WZ˻�On�T��-{B\�s����ٮm
�ԩ�θ�]���ǩ�r��������
�]-MK�̩o��n��$i�O����h�)�c��Mٔ�F�PV���v�]���(Z���F��4� �����I�(�.���To���"� ޷��q�4f*�� qAu����w@f\]N��0T�b�v m�#b��CZ6Q�t��E���U�,;\�Gzxܜ{���73L]&<o�cr�9�jO�Ɍ*�ct2�B�:+/�u̴��	�Q����|�>�i�1��rV�8���P��ub]��Ƭ�[e��l���ܔ���6��}���w�[�c�-��<���aR4�8fo�A�FV�
=SL�bnPW}ǰ'���6���ݔ�!�%ʔT�7���T_��7k�~澅=�h�F��ı����qӈ�9j���"3z�f�m��<��ct"�*���
�f�''&����Ӿ�_Zi+Zز�6���k�h�k��Y���dG,mә�6�4��5-t⮭�3:�0�z�������ɫu8s
����7�横�X�eYmQUu�p��1+DN\d�-+���&�q1m(�,�����q���k��*(�E���:n�S`�t�3F��UX(�{��2c�54�6{)T576z;��8R����,�eq���e��f�PPA]0�)\�fSxLW2����kWE6p�Æה���,ٔTUU�)CmݧR�DFj�R�i,t�{�"��⡚eEa��t%b�)��8pt���9kM���T��~�̩E����E(�����SB�-�l��g+(�̢�(��<˓Y��Z�[U���Yg�1r��b��Z(��2���r�E0���Ç��TdDX��LeF���ب�,U�E���Nٵf�J��m3(�����H,�-��hj�k%T`��3M\�kD����B��ÏGg�e��x��`��E��z\]��H��Z��/oAGu�Z٢�L�8ntf*Qp��+C�!��^B��z���ح�/8��G6y*�����y�(�ͣ���k�gcA~6�%x_bz����@K��آ�]�$�����-�^as� �׉i��)���S��#}ϼ&���cz�c�$)$���N�9㺃TS�ږ�l/2��Kf�1#:83ú[�E5�O`�V[���ܮ�bP�:]t�0�ojbj��03�B�<}�q~�B�Y!(�Vf�h/Aԣ!?B��L϶�� �PMM.�x����E
Ǘw�^H/B1�ʕ�˝�`2��)�\Ԃ��2��.5��U���zD��6�r�sn���x-�� ߀ޯi���9�@�9o[]�7#*#����he&,j���6�Ioܷ�<�����\���b��27�uf�#�`j}�{>�"�)U�^t�Ҥ=N���P�\��Bc[�C������TzӒ��^r��|׮�i�gZzC:���Vv`�8f&�
���h}s��/���aD���HP���0 ��X�:�,�9�H�kx2��%������	y3*��]R�0��'E��r��ϋ#�.���Z+��鼽�g��2��HTٺ''�x��������8��YfP�#i��ylW+O6�ü�ħ�BZuCvLA���uU��JT���f�@�$�i�[�r�X�`�t�������!%R�{�8�3M��\�ޑ�2Qr�H��C2)9��4'*��]�3�C :�f�n��M�Ʉ1T��������C�iu�7�	���dzb�&�A��篃�hj��]�ޖ�s�g�	�͇n���t?�x[���P)k�U�QkOG���}��QS���2�0I!�n�%������5����¹h��i�q��h��pG%��\VUzFz�w��	�������C����ѽe8)@�z��~�UZ��c�j�0nh��/v۝�~����̈́��T�Ftq�:�5�b[)���\<m�c�i����.Q����v��zS�!�Yt����i�����b�$r�M$�;��8�y�W.�5(찄љ�"n����5�- ��M���(J�w��E�Z�� #��N�Nr�[7Q�m�od�N��:ĕy�7&nUo��/-R����RMoO��$xoz�N&$_+��&Pl��V���1�VK��~�T�s��
���C�)�
������A�Ej0�Ȓ�#�RQ�����m;��;�<Օ
Y�cث��g[�x�TU�{OL.�=[��zb��+$V��X�SP��IE[ˮ�Fi�sF|��/=0*�Q��C���k+ �1}gMvJ����(1Sð��{{o`�Cq6(�n�"�	G�x�Cmn�#!XD_����ڷf�r����wr����')3�ЎH6��eG�u<��N�mVQ�����~QwN�!�o���-G
/���ܸf7֗kZ)�WO�1 �dA*&�w���m�i�Ra�=�ڇ��D�ף^�Q�ՙ[[�9��,���`�P���5Źw�Yz�����:�3ٔvqF.َ���g����g]�����51~��'~�R;�A:����Sy�j�TE���(+�45�ԲWH9����BA��
����\vb����z�q�O�uڽ�����~`TE1��∿���&o�+��?[ *�����b�Zb�&�S��}� �s{��>Z��I�%R��N��Mף��0�#�݈y��˛{L��SBb�����X�a6��O\��j�R^l��U pї,ڮ`Q�˓��0�W9�B֜EZL,�w�t���t^�N)�9ƛ^�2���c��3	0���W��q�c�Μڎ�iIk�b-�]m�rٱ*���ɤ2���k�dJ�˒A �1Huz���?�w��KFv�cq)1qV��8�΃��!�%Ь��vFm�w� �/k�oJ ��,�
��'��M�~�G���}=�<秷3.�����k��� c���f_D~�Y����A�Ʉ�� �<�`��� H@I�q��D���F�Up^!&�J'hieX�۲j�Nh?�j�E@�;M��)���-R?�(�v�<{�2Zr3�c�c��kW~���a����>g��`�hT�&!gJ|{T03{|�N�1I�� �{y���@Wo6��%�/�k��]_����*(q���L���t�,��k�1��U�lz��I���9�ςU��y-��)�2�u��/�D��� o�|2ߩ,R1�A�K�7��0'�K��X<�������l�_ftN��j\B5���1�doX����(A��i����50��(�;�pڣT[��V�6�c9oo�r[�O���z�-�ex����kD&�0e���X�6r����N��,b��s�xv�QN�b�Ta��$��J}m� n6�@*��^j�X�0�yI���Two�;���z@�Z������n�t� G��|�:�P��&��Q��CU���k�M�֋�i�t�[�#tF���0������s(6o�x�;@v
�5�?c�Oߖe�u1�:'�/��je�u���Ӈ&����̳Ð����pz5W����It���ۼ�-���:zU��8<*�S�`���߽����\�WuW�\��-@�㋴��P�Y��\X4�����~l\ʹ��~k� ��v8d��Tưz�
~���6�EP��9���LY"��[,�p���UrXQ�8H�uT˹
�����6%J�&54�ѩ�=��}�{<��m=γ:pͩ��)|�r<���s��1���Y3�~�ڿ��R�\���榞U�;�������Y5dˎѽ��[ՍH�=�^������!��592��0���G�]�IWꯪ}٫k�N�;�a�P ڇ��_r�"~ F��z�@!ٙ�xټ�ӈ~cR��IS�����i��(l���T���&���c���1��^������������g{�(�/�[��I���E~9[��Jn�������I�V�l�;�6�6��Խ� y�l5�fvK����\Cj�]ˋe���>���~vGA��_z�h48#���d�??�l٧��h�T�_Y85;
��	
z����צCǉ�i���aw(�4����yX(�/dөv�N.���}W�-�=fQ��s�+��z��MF��#m�D�j���[e�F
�S�ã-ǻf�;"EU�."�~g�ڡ+0�����b1����Gjj�]�5�5�3���3��Mlv3�T7���sQ����L���`S6�r������"��,���|�v�C�*p!�a�����j�?�st�#+�i��y�Y�1�W�D5s��1+�Ƴ�O��1X�w���ϲ�\[Rل��F!7P�=��ɫ�`��0 6�+kZ�j�a��<7z�Q��Il}#�U�UiWNӱ�Ɂ>�7shP���.A7��͝�0>6U�e��sc�Y*�
�}�0,.��ei2V�11Μ4$R�ݡ�4���p@e�{�%���
qn���E�Z����O�,;(���;�q���r#_o
{�}�Eb����_����zʇ�Ҷk�7�'q�Ç0���:��Vυ6RSx�`���z͏p��͵ܠWP��L�y�e�,��p;����kL�M���S�/<�A�v�@XY����W@���l�mc3Q�f�]E�5+�>�$�P���aR
�H�]�Q�1HH�}�'|��O*L��
HQ�6����!�`4�.�����}����#q0�SzC}	����bS�0=�gWY��8������{�/�5ۋx�t��z-^�ꑲ!�%�0�p4�w=y�?�H����񊩩'��OF�L���.Y# �hNQ��9��'���=$�ý��sߙ0�s�z[�%�:�|�[¸�O��S�yT�UܫH���+���7���7�^+`�M�}��c2�U@�Sai�}���xZ�2�p��o�Y[��
o�N�`vx�IN741�Z�����z&03�k��J/�Sf�\������$L�&�#��8�� �ӛ���;�����8��O^� ��6�B���ǃd��.�X��y`����u�V�q���ܻ�v�Ȣ0�O������`��%
�_֟b�f,�˕"�\�G�t�hjwʞM[�P��"Ee��#���ظ�fk�ۢ�e�G��y�/zX^��w7�W	�ԡn�MRJM-s7���\<j��*�Si��SGmv�7>-��d�d��hus~V![-���69�34)�A9N��K���ls/ڎ ^*�r�o�15E�����U}TG�<>�`�&�f�V2�gz���O��#�Q�Ed�,�4�t��1�>T�͝�$�,��1�>)^���ȋY1͂j��R��<:LS�e�{b� A�DW(A��Ϸ��~3�h�>��˚���O9L0�?���NO����X�H��acM�X������t�����YB�۞�K��Y��\�i�H/�g���ϫUvF��#s���1Y)�c�r�^uG3�Ʈ�L��b�o&�"��ɪو8aWT�2Gm7R�q��]���c��m�m
�s�P��o��E6�[�a����c3�""�{����i{f�P�t/�(�v���2"��}&@�?v��<�0�7����V�r\h�$M�E�<�3+����}l��$����L�LW���T�����E�{�۳�>�k�^#Eu��jC30f�eգ!��uZ`,���\���YVh�j�C����k֊R}Պ��n��geM�����)���Jp&�|dÉ�j��J3�˓�0�F��$��j뷒�jK�ئ�����u��i�V��h�jn���Tr��Չ���^���K\�W����6�	�H�6[+�7>�Έ�K1�z��|V��1M��w#���xP�t2�4p�4�;�Ή��/WU�u���6���W�a�à�����k��� ��՞�=�$;Mļ��d]�P��E�޾P�Vv�=Q��-tiz�{���l�uجª�g*�s���ab
�	:��DC��������ޮ��N0���E��Y�������%��i^��0���~^�� ��C�!�A����}]�U��04�sT����kU�]}���Ip��ka^&9��>��K��c�oR,my��x�dEj�"[�����y�U��Egiz��Ⱦ�CQ��'����S��vN�G��0]w�"Ħx[#=�X��Z��9&�������E�Y�R֍�2��|�4���Oq�c��A�}@~^�uk���JEșlO�u{­��@��;��=!�_k�y�y�G���S�bu׆s�7��0"����� ��#�����������2��th��Y(��^�����W�Ф0yeg�¾���0O���ςm�s��C]8y�h�w�#��6���U�v�(�]qd࿉�=끣\���
��ůaN6h�x��\��s�	A�f=�ɋ�yz�n�3m�ҳ,]��v�g�!s[�M�f~ o��'�x��Y�oք����ܺ��e��ۼ�u���5c�B�9�U$V��N"�c�`��A4��.n3G�������:g�nY�&���23h�#�ҽy�&9��%�ṩ�����e�o�j�Wy��:�'. X�y���,AbM\R��]N��Ħ��,�
�d\�\��e�7����y�+���ԍ`�DZ\�Ҏ�z~BX���gd;�ϡA�N0�����d�\�m���z.&�m���aUR�PС�v]�y�n�Y7P8}$�㖇�\hC�#c�	sJ�|
�m?6'��o���Ƭ���9��{���B
�#�DD֩�Ck��d��P[�	�d����K���XI��I�o
`{�l3��ٮ��Ɉ��S�u�.u��>a��"б���K�0wt��*e�E�-M،�
��͡sR����r���7�P7	��b��\!�]k�o!���X�d(<���(�M����5��{m��T��uL�i���Am��y��gZ��v: ���Y�@%�Y�~�Q\���(��ыL�k˅�jT��q��6�;�驯H�r����?9���J�4!�+���u�f'l:�X!}�+h��ͯ��A�y�:hs`w��t4W��j��/:�9��h�y��̫��<��pNM����:���!E���[U��� nq8;��8�v�5��1U��@ԟ-�b$f�^�G4-����u2�t}I�ø�$���{�`��x���C^���J��މ�͏w1�C����q�$Nظ<�X��D8蹠a����f\�m�cb4�n���\O2�Z~~DbF0b���;��s�����˒N����UG��?��A&r~*���y��um`�ً�R"��B��tc��d��K�pu�H�o���C�J��cJ����S��v�<힗��ƽ07{X0�=��kxp�D����<�5�.�,����6^�Pž����=��G1����
:3;ON���U�D\.��/}igCj}x�{�2i��=#���r׼�98j�tc�1(ǆJeK��A���'���;P'������]�C���]�I�|\fӬ���	M���
�m��YX�f*̙������9|��aM�t��n�9�O���E�^s�7A�_��NN.�{%��­��x��q}O<��15���^h�'�O�Q�t%��aG�e��2C������d�\ݘc��[Gv��դh.~���=�!ϯ)FP���9�p�J}���K��u�Ų�c*�Z{��vm��-���ZVSө3�c�C���6h6��[ Լ_=K�~(�}�Г]gLe�(F?�nMu=��	�9]n���ßfi�ϝ�m}�b6}��ɄJ{�a^ȥkoҏЃ�~��-�-ʮrhD�h�48A��:��lѤ�VَU�sb]\c�icd��E[�e�Yӭ#����7�ݔ�f�tMw��`���r���}���쭫��a_us�V�*���DnEm���Ϲ��[����}��3.�+Y|p�.���2���&�Rt��ԐK]Ni�%���G��Y���,�؋m:㴪s���A�{gQ��7PySv
��-_�]�n(9��X�'��g\F̭[�cM��1�A�U�u��S� eЫ����ʰ]n1/���I���AO@N�ʵ�D��d��W�?C�-x�{�Y��dłqm���{3W�ȋ;��9��W.�!�!����Z���Mn-��
&�l��o.S�%%r0�h^)�_6�{!�ʳ@� <(� ���p����oC�V�J�F�H�T�+��h�0����(�ZME�C��S��n�C2�=�l���׆�͹r�a�sE��Ԫ�D����e��"��0�[=��F���z�����;��A��w7]�ӽ�i4�r6�wcY�'�����FZ��]� n|M)���ywn��wA�9��јѳ��A2����&�V,�s���ً�
�4�U�]�R�!a�P�Ѿ)�E���E%@ֱ��#�w�����Ϲޤ�*����]z���q�E��N��E��e�խt�r]_1x0���,�rIA�Un�
��R�7��,300���l���Q]�Yi��F���{���_�]<6�~�(�Vk|v(%LD�C4)u�Orat�n�T�wK:q���ϝ\Q�Fo(�Q��3촙ީ|òȟm����D,�o�-̓�W�f��o�op<�&�Ԩ���@�Sz��BӾo#���\�nT��9|�-[ÛE�ѻ���&��y�F����m�IΥ�b��B��38��֚f���bŐdW���!�Q��w��zᮾ�q6:�v����J(�Kך���g�z��t9�ԃE�9��#����u���=��~���,��4�;����\¹�awo��C2�{Z7f�X)��5��������M�2AxV[�εW��� �T�(iY���W	��M�.н�0�j�Ɖ�K EN�S�ӻ�:���|�$+{1�2V2�%�(:�?�߫]�^Z�/N)P�J��{�mͦBƢ�'�`���V�7�eg�fU�<ݾX�{0eM��V���[fXD"�1|��\�1�Tr��*l�1� ivs����[v��Du�i��rv]��q�z:cN��Ⱥ���B�f¯���Q�Rց/l�}�v��nV
ƥ���f)A E���ѵH,���	��w�>6���T����bAڴvQ��i�f8/����-��ۃ.�Pkh�ջ�������Ih�9�U�#B ���ɰ�`qpOl�����6.���A\5�rZ8HM���TD����@�ȗ�(Ѐ�R_�zۙWPէ�A�(Y��i�b�N$�iBÖ��Dӫ!CLSr5,*A٪��H4���3*��n:"Wߘ�O0K�q�Z����k.���D�dEP(��E�j-�d��DUADV(!gggg'	ȉƕZ$PAalR�b�b���Ա"��fF*:ֵ�d=q1UUFY�����Ǒ%V�%��(�Q4Z,Lj"�R"�(ʽ̊)F�Q�\A[gR�-���MN�N�+jJ�[m�b2|s%b1uJ�Eb�*��)T��Z�3T�YgggNG��\B�`r�F"�����r�dX��f��\�mTY"�Ç@Q�3((��Ƃ��&Z�P��Z�Xc(��Mb�Zy���%m�E�*1����Mr��x��+D�)ƺj�Z՛�F�D`���|��AE�����h�!R0UfZ3F<x�N1X9J0U�!��F,UDQ�VrՊ1b����4p�Ò^TH֨�����mtZ���fV(
���#�(���X��Z�хj*e����,ƺB�(�5b�j�+b%~8$�k*"ۼ�[J����5�o��������^��/�͜$F�[����k�g���)��Ѵ�<��2�g+f��/-WT����-|��Fp�Y�f][���c1�A��!'3]�tC�� ��0�=/<��b����"��ʋ�3���ֶO�o��V��M�AF�C�zDvMn�`Ã6��OeAWK��R�%z���@5�c�#C����g@y�]�����GL�Ʃ�2.���b(;āNu"�5���Զ�V�@����r2�S�8�lj�F��f��LD�l\��W�J���=��v���2v�<oQ`�g^�z���5;����k��FA��>e�%r�(J�̜E��;�>�D��Z�'���ڿ���G�ko�d\��y�|#���Um�>EOz[_W?�~q��~�г^�|�\���S�o4'��кa�ce�[{5�#A�Sy���i�����IC_D�s�P��o�]�Fә�x��ĖE�a�~(g4~�k�m,z�#\�<'�B�b�C���R}�r'yM��Q�؛�w�ݛ�%ؔq�5�v�Ѫ�/F��S@\�}��y(��dp�>9��Z�Q�9˳�vz૙V�V�ӘN�����ܘ�d|,Ax��Qv1������	kĺ�a�Z�e����`��ks2���'�:���h#C.��Y��4��a(l4�{��~ҏTXO�2ϲ�{LA��B������9g[e낪P���}�]�P.�������2r�pp_9���q�� ����&�PM�-�0�D�*���D����=�I/���0�1��0D'׷�w�_hs�R%��ȕ��j��Y�5����qԸ��T�Z9,� �G�b�j�L��C.�m��f@R�F���N�'�=�)����}�v#bjذ�J&���ط	-sU'�*��Ӱ��Hl�^ה�,��2���fqt��2��3E���[���`=?�Ru��Vw�n�����+Z��5"��X�_3L�цO8�f�X`
L�G����F��m�mZi�:������1��E��:Z��Dlq���2&�r�/�vF�翜��c���61�M�9���S��3�N{��n��%r���BǁXA'��"�l��z�il��V4Z4큙���0(�0���u�T,�f���#Q�Ӄi�̀������d�c3NFѴ����̣���Y�|��$n��>n�©lC����s`�oW��:���\V��q�x��C/��)@���#O���سa!Ԭ{��ٮ(��-��]v6<~����3&%��\�;̈́DT[�&e$��X��kq���h�����d'��A�Ή/�ٺgvҧ&���Rܻ���?G����]0�Ji���纫��H8o
�����YE��b�<��[���ݩR-^vH�(��2:%t��@�l�E���ʥn&�r�a�'�x]�<a �q�\�
N���̃:���{\~o5��-���c�?#�c��A�;��|�^Z����!��8���+=��W���o��v KH��od�b��}�pM<��K���64sh'B��O�28˯��P��8j��3CH6f��׉�2{s���<�^4iM�t��X!G��~��t`sr7m�Z�ݔ��u�rƼF��Pz�#�Wtχ�����J��)���X'�5�AYo�1��G{[�t��`��	О���Qa@�V��v{`��k�κ��..86�Ʃ�ne�R��`��7Ց28�^��^�:�!�Ѫ�9�A��L-&�Jn���� ��I�c/pn�s+�3����T��7����b��>�DSu{ &�cZ3��.-�*)P�DO,4�φ�NCA���r����+�������*�F#k%;P[�p��LyW'5�)��dK�О���8��u���z����jĐ�,x��T|C�������;c>�4Um}�b`W��^ᵍ��y׵DQQ)G7-��}1\=Ĭ�pNl2q@�ѐ��4H��M�*�Z��n��iz2��M����l���:�P��3tR�Y9%��k�H�46���j&l�{��G��Sb�n�2P3c�os���-kDn���Ԭ��T�H��k�S`�b�g;��,�2`%e��`��S�s��sc�|��-��~D���,  Am��ܞ~����E5w#I�5Ig��W�I�i�� ;0���� Xא��4!\���e�Po�gguX��~����uI�\�Q�{��Tsa���8S}h��7�+3�[2tbus�0ݼ]�edE1*������z1�b8���c�AgM�I�JǺ�V���#3��`����=󂈴���L�a44�9%������ݠ��v�X/6�8��^��0������G2>}/
��X|�J�(�7ɜ�?|���GjECaq2�	e��y��l�XL������Y��J_�i��@j��+�^����(=+T��h��W�;�4��V7&�̽��.�
X#zkۤBI�5G�{�Cʜ_W����-��N�B���R.�A�� ��xYE��B����sR�m�u8�{8r�f%�m�����kUb����pܣ���@��沗��4 �$e�..�:h����x:����s�~!l�lJ*ޜ���SL���ɼ�����H���;+���b�ڄ.�Yc��\p~�K_<�Z^������|b<b|k���6v�+��k�f�T�;�v�)>��7��3�>����ԛӑ,n<�:�
�J����U��u���W:Y�^�\���6�a�C�8� h���u��jb�3]��^u\d�v#W�O����÷h��j �V�BA�S5�o�O��bH�A� D",����UEۘ����uD�!��������6aR�M0�L#x�@}ƅ�&�Iq;%yᖚU-��T)��pQ��=�����!�aE����Bɹ�C/�}L�Ho��/Z(��,��\�r["v�7�KOm'd�U-@��]`O�|˝��NP��e�X�q�֑�/�TO��M�s���˘�+pupsT��T��(�^k�B��݋ǯ_\���,��<�����7�v�Uz*�^�����`��K�t@{��1�EPʋ�a�gN��=G�|E�4���y_q3a����u����%�|T��������c�y�Fȡѽi8:��i�GFQ���wZ���t齭m�&9S�/��?=D.&�(%�S�E��[t�Fs�n�:��E��溞�֚װ����/�������!C��;]4�A���s�������.L�mx�j/��"gӾܼs0?�PtS8v�5�K�s��R�h�>�^J����'-Ş��>�Bڅ��-\G���߬�-�h��#�J#:8�Y�I4��*\��]�d����&&�����̡>]aI����J���;X���\:�h=V���!���K%�×�d��r����J��� *���A�����&9C7BK�N����{
ؒ|k�@��8�[�h*Z���D�ܼܽ���	?"c1�1����1� &&f�]{wG�4L]�B�!mWp>�S0�+#�(z��FD�V��w�r�����6��S;U�ǃ6�zr�=�9�fp�"�-\�Q��-�!(V�&�Pcxb�(��+�T]P��;rِ�����ݴ�
Xc!�&!�ݷ0�j�q�䭈���09�L=���@��g<閻�[�Pؗ�M�7d�~�=�I,���I��xW��h�F�̞K8���P�Ś�N1b��Ƹ��=��$�۞\�9�\�Tyw�/�����9[X��)�>W��$����D&z؀h��*訷�ΆZ�3@�S���:)�ŻSoC\t�ȹ�/O�¤��̵��`5Cxh�u9�	��.��Ѯ����1�<�2Ga���)�EI���ʹ��qBsC6v�X��t�x���_��3��5�-|~>���8-��[�=�p�lӋmV����[Ala	�qq�/�K��f%�}C�b�ʃFQ\��G*9 C��>ܶe�B���q�0�:xR��c4ڲ�[M�ýf�1F8�T�֯.Ni�ߓ�b�8��4�e���|�|�=�Yx7`�R��z͗����-mvt�LV��"�-�o�4��"��isl�Z)�=	����X��s��3I���rG�F��d��֖��[u�H�?�����fv�w�f�څ!�)ӡ��hTۜ�����Y�Ӕ)�n+�DMW��N2�&�Q�o���LX4c1�@��a"0"  � Z�I۲v9��)�*�s=Ԛ`�E�_p@=�`�0� S�~"³9r)H~w�^��9}������mi�;��c�,����6Cѩ��b�g��'|�h�k�@�|~��F�y��:ao�96��i
N�=D!��18�/\`c4��qE�׌̴:��/�Q2���b[C���v�����MfGzhV�N*kb�KZ6�d�Jr�6��IV�(�00@*m�SE6��P�5D˫��e�U�n4Ӡ�\�D�t���@����cETaM�:鷕Azp8�o�gk1z��͉H*�B#��͓�o�<yQ�����V"5?S���D"����p���R�q�kp1Z4"d�����+^���U��&��K��N8��e�U��QX��ǋUS5���Fşk.�6�;�u1~�˯f��J̱kr^@�#bvm��zkn(�1�*U�s��CԬ7kg����xL'��)��2˟��6+WXQ�0��3Z.�����[���5*�(�-8;�2����@L��8A�m������It��UJn�i�\v>�5�ݽ�Ԭ_�����.f�����������A��(�n*��뚡3}�7�b>��KD	���-��
��6����h�_��@]���mM�fͩH���'Gq��8oG�a�T��9v�97.α|�Eb�����2�\���c�����HF$���ĐFG�Q FI�>��Ͽ��|��������0+�Y�O�슓E����Ը2��!DR~l�d�8������u��e��K4k���c�g�N�C���	0��ȖR.M�%�G`P���*���y�Xa�DWl3�t*.�Dg.�N2�s��Y��R��
�C}�#o�;���¾��q�����0��ڤ5�i�e�01�P�ܶ1L��T^�@�x����B�*���n�Κ�P�*4!z3�m�1�ɤ@�j�_����R����zC�P�X��v�3Ϩ�A?���{ޔ;��d-J��:��9:�_>S�Q�{��MY��K�N�a
�sf�5�m#Yp�+{r��2ׅ�4����6��:��9�i�BG�}�]0�<��-���*�t�0�#%oWwFOJ���Xgc�5.�U�,����Z\�o>Rbkb����v��l�L�3LEn���iD���E��^l�/���2��_���;k���_���ܔ+̡�|��v���k����v��CX�&������p��WOO>�|�2Ȧ2���q+9,mꗎ��kyMvWj,��7a]���}�J�(WV�M+\ΙY�}����6u�[3y�,�J��ES��e��#ݴ�[����⇒�d
�*/���=FHp+��;��	z�S-����x��q�B2l��b��Ί�aVԏ;��9r�B�;�5&�	��!8ceܜ�����I#$�A$FF X ���[��G��{��t��1>�Xe��{��mr�%�5e;	���+����|9�w�vf�ߑ{�\'��t+�qnK�l��:gxD�m�+ʦ�mk]�S��ם=��.��~ʽ�Ⱦ%����j9���B�L�)t�B:$��tRuϋ���G�[n�f1�ʧ+;vW(��C�I��w����1m�^�R��2h��_T�qo�ih��O�8�{X^���Ik2]gO(�Z�g�E�<���v�x'���Z�+�TDa1Y(��[z
�ؗ^]�������3̸�x#3x���3kʵ�6ě�#�b�%�{"rg���R�9����r�2���Х����kǧ��w���N�|��K�f���dY=n6���i�UC��v��t��t%�]��}f�|����~Y�����xg���I#j��;�۪��sJ��3;�
��E6A=�x*z"��/B�]�bW�#3/�Xv{c�׭l��zʲ�i[*CNk�ՙ��d�⛬#K��|y�� ��Їa��='}07=��S��������>���mV������j-�{yw2\t���^t�`���^+�3/m�����3K�)�(�V]����.%�uT��_&M��z�̫���_j��ZP�Kl%jB/s����S7v�Wq�C&�l�)�)X<����W�Ϭ�$�cH� F@`��4��_��p�W��GG���ȐW/D$�P
�Rμti�x���k#�g۪�1��M�G5R����+��2����oQ�����l;TΧ�!Ӧt���G�EZ�18<w�x�սR�̎���?Bf����=�}Cw�:'K���#@�y��ג�{%{���-@X/|%��t��"�/�M�ӓ>��L&��(/10����҄�\M����M6�y3��7��j�"ʓ����1G���]��}ʢ�B�~����li:���z`��4k��m��Y�ܣ�ܔ8t��͢é�[M��w�U7~�2�����)V�1�c>��W��Zi��gԅ\���V��tLÌ��Gb��Sx
ڇu<��x�P
�M���7>��z:�� �N��{tm�]�H=��1�E��n�S|�nS���:�-�f(��P�%Cj=���#���'k>���Z���IjfO�p��&������T�;c�AGZéq[g��y���+2��[����HA���f�P��2���)՗�c�s�O������F�{�]�R� 00��w���JH�QCݘ�`�o��&q��l���
ލN�,�t��(i�L�K����.��w�L�1R�ִt����UL��V��e�;\����h����4v� 8-[q������M�T/-��miY�L��g0�9��N��	����9��Y��Mi=k��<c��{��Q�%$tj[1A9՛W��f"wx�N���O!�nSIP]�4�/3�� �*T�U��g�sv�����\����+�o�����%@F�1�B�{ZD�1��m����̠�k��
��X̖&�Y�:鋮yC1����;ax�h�=�-��5�6��1��:h�h�ѹN�j�Ud�cS3���\7�6ŹJ�=�Ηs%�\�Hn��r�C���x-���������bǅ�TP���|��Ėa�E-��dۭ��t����ng$����.[��Jop�R���.el=�e@l��k Eb�:r��p+J��nkz��Y�Q�굆���
�_p���wk���o��\��b�&q�v��[��:X���\��N�o�w�uL�n�K�g*Ah:�%��V^��d�����r�M��u�7+'D�h��s�|[��k�e��f���nm�kq���XMe�̮C@�hҝH�������U���ƒ���
��C�q�r�b��ݽ'�A"�;�h��ُ�l�o#Y`�����M	=V��h�2ql��\�s�Z��a@����"l&slJkj�,�f�e�5>�y��{ٹ�Y�!s؃�X�f�h��[4�S/�V�IX�ˣ;9dZ��9��t���u�A����^�)YU�ف�mwW[rVq5�!�(�Cs�jk�v��F��MU��ѷ��#A�06$bu��3�)�:ټPD6�2%t�� �*G��=���!׵f�ξ �ՓQ̲�ZX��쭒��f^�"IPf"s�k�B��V�� ��Wp|�d�k��u
�]�;�%:#�Y��7�pl�vB[��'K�z��b�0���l���]A��VG<�/��!f9M��Y�+8����b;0�bW15��y��6�H�R	aV���L���WA���j�(�+oM����Y-�{��L�,����j��i9E-�_Vp9R*k�M�&��/bo���Z�%(P�z1�GSnR��y���Z�4K���f޵���AB�����k�l�:���{S7��d¥�s���vIQTr\ɹ!����d�fvY��XǢ��i^PE��}�ײN�j��d�h�a]�5	iHw��a-M���b=]yZ*:F4L�d�	I�o��:�[i�E�:�)Ą�ʭ��VI���s��Q�k>�S,L;��s�r涧V�8̚^nB�1�,���Au�,�*���V�ؿ�HID�MM�*����şMU|�^�X�IV%j+��e�F.4U�ٓS�j|����\�D�*"}6>��Ŋ���=�F����TF
��,e������*V�UF"TR�)iWMF��_�b�%ul�Ƞ#q�a%]6d�������@-�N�Q�ȣ[*V[`�
(*�oY�P��1���ȱEְ�%�-������5;7:r:�tfU�ز[N������i����cZ(���UV�X���gNC���ghUS�F;q�J*Vc&4F(���1��.�X#&�6l��~4�Q`ɉDY߫1�b-J(�*�l��V&�\����+eH�<xٳ�kt��`�Cn$�1-h�b��Teh�z�e��Y��ei��Ɍt�PJl��gD���qT;q�
-B����1(�E����dCMo�`�f*V ����¥`��4.�TM[EY��k(�T��e�h�'m��\�I�X�Ok���Qc;Ok���+ObP,�2���*�6���؋.�K�{��v���iw�2��yyv�]�d������/�?RI?#$����H �$�#$��!H9����w�=���Ո�A���ה���sZ���0�����1�n�Ͷ
����ٍf�umwqUv���.x??����0C�9�ԣс9��=y�S�(d�0���[��h���g�m�LxG9�^�A= IM���0J��C�-��kv{��g*2�dNv��k���/K�v���>��+e	�D5p�|s�s|��+H&<���#S���T�ۄ�Ɍ,��Y{�_˄�_x���M��T����0�k�}^���q8)N�p���{1��N{R.-~��{&���&u�tt�q|cZ��g���ƪK���@�ԉ�f�e�d[��#�t?��^�uY'�^Nz�,�[��W-��i^�1�J�-���4:��abz����/��U�;� ��n�=rT���ѵK�q{�Ui�r^����u�$)�5���g��=�qQ��Lr�h��w��������y��*��HY���q�r�Q�c�^S�*m�+R�8GvZ�Զa1��� �nϑ2Ҝԕ����T��2�>�D�.�߷�[n��1��b2��>��oj��e�iߠ9��ܦ+���'���J�ElK������
��i�{��T�{�'w>�@��s3R[��;3-wvh��^�Y"G/���M�e{+���eu����$�I�cA��X`Aff � ";3;G�����D�A�!6��H�z�kл��Azs�� ����s0�:����;ǟ�ev�Δ;#��ll�n�kQ�4�27�X�~ު�=u	�X�iw��ޡX�=�y�˓O��o�qk��Ԩ��2A�~��T�����i��l�G����.p.�m�-]c
	4fL�H��o| �S6���v�~�Aܶ+��.z�4Y�A����ه�9�a@���~⤋~u�r��朮�jK�-��*m�^��j^ PxƊ*]������	�ό���ik�iQO�m���OUS1�������߶�׶CQ����)��5��1�2�;ǌ��O��m~܉c9��{Va4H1/X�^�Q<s":g�\�V�BO;C�Z�_<�>Ո�hX�ֆ�B�_�!6�\���J1CuC��J���|�?p�,P7<�̷݈Y������PuL���T���L�����04.��Jp�x��4t˚�C�r�^X��t�V��VS��n�Oy���٭>tsF��u���g�\���D�ׂ�C�j�B<���R�-�01�cg��q�v=z�H|3�y��#��Tu���R��4Ve�f�hM&\��[�=�M�+I����\2.�3]��6�6�p�A������9���� �����)v���Brt��ZӉ����na�#���tc%�
vf�U��庽Yկ0�w���J��h:�#��-��|'"���h�GH�0*�:�ԒI����c A��� C B��"2`��n]���d((\GR~�#j�&�Bn� �������@�T:��v
���]�(�[5[d�Q�����H��UƀZ�D��Π'�<Y����q�E{*��H��T�mR��1�"ٌ�k�9Q#���	E�j�=r���$栩���}�M>��U�}�t��aު^gU�^����t�_I/#���݄F���йY���8�P�37�_����O��B��q��x�xY�`�q���y�c�k[�x�B���V:(�ͥ��sP&����8F��>��}as�l2�O75 �<,}�1i�ɲ��*�l%��eq��s^��U�.m�wu��~����܁�8�������O��@L��l1�蓏��k�آ�8�)Ol_Z�RjwI�{��٘�zd ��kX}x}+g�iQ���Gpd�8/�EOr3E�}{31��2,�MyG���ǹ��x�Y��j-9%�&�kO�u4�)"�x�@�M>�1��'g�+��K8�?F-gc��2uE'�*A�VnF�*�CH��2]����� 9�bڼ�]β�'�󹕭�=I���.��z������$q.�[� S����.bҋ�q⮧�t2T�!�+�|E.U�^M'պp��Kn�ʬe
�<�r����Ѣu��/C��{���j�=��v��ߞ��I~D$�$2�@D�2� ���,�Y�ݥ{�86~
N{Yz^��jZ�ܢ�ǹt_LkbG�@������(�>>	M��U���#�'�O�Jg��=�8�j��o���B~,�s��9�>�Qz7����n�ew�$�Gx°�]�p[�|]��2�T�"�RXe��t�r<� ����1z�95���o�r���v��p��� ��P��ՅȜTҴ�V8�6��W��#J����z�� �yd>H�U�_s����4'YU���<j/���bRٮ�vFJ��掂)��U�����XEClG��!Z���[����dh:,���x�Y̞Xi����'uT3��n�7�ܕ�l# ��!K/,����K��S�������m�o:ҝ�|�cN��pz�˒���ˉ�}��m��*�z�FN����r�*0�obW��	R��>}����8����fa��y�T�-�e�μӃG�]$�w��Y'����(]kG�G�%"�DY�b���[��J�����ϸ~��8�ˢM����t�ai�� �:B���� ��B�I�m�K���]`���P���}�i�iTE�G�u7L��9�w�N0�29���9tf�T�fPvyA׎V�iwb��U�v&'9c���L�����wM�=�$��0� ���� "a!���}�}}��؏=}�H�O�,�0�ъ�!�mC��k<�i4���~�N��˳T%�Ȫ[��C�(��������� 0�	��vq�n��" ��h:�
�gz�������uR�}�_^V��j�X��t�����钟pI嚼�UC԰OMx\�u�Z�R��(D5zvv�7^]S�{xb��40�uI���:L�˟x=�^*�mɛɅ���^zr^'��o�b%"�B��.	i�/��З���CU���!��I�-0��#�*S.�tO6���8z���]�dw�����b�!$��O�=8�zǞy�F�ხ;�mW0�j{�z�%�.�h^Z堽����AԦ�0��9��9D�&���C��>ܶ[���o|<��1���V"md�;T���&_�Z���n�� W	���:�ũq�%q�Z^���.r�G?)�;��6���CN��G�ݪ�U���ɿMP֞1m�0m:�:�y��:Ͼ�����;�]������S���sLYW�;w9�^ڏ��F���hy،�v��-�j����^��(f\�
*�H]Vb��eZ�����1�N�v��lnJ��-Z�J��9�'�z�fm�
C}b�N�qv�络	羯]U +g�=zX��(;�} <j���m�fU�z,t:��R����D7$�f�es{tx ���~Ȁ��$ 1$�	"	Ϯ}�Ʒ������~'ܪ#�K�^�۰���mrb�Ux��i�UE���Y��v/;��MC��L�;^
�~wantK�x�*=Q��Z6���3Wy-T9����6���V뚮�/��Ȓ���~�u�P��Cj��)߱�Ň�K�TGc��1����H�C��pm�@��6�}�D9�PNB���M<~�_��,�/5���:=�[
��d)b��ZگtIh�6o���z���)m託�Ո�l�B��@yml��*����9aJ�r��5�hu�7T�~�a�O׊q��
̱v�i����;�ǥ$D�bsj���C�{ki��v�W��-_����3)�p��E�\V7\��0zWK$���YZ?l�0KF>Ҋ��������k.yނF!�9R.���2a�T���tK3��3�չ������+x{�N���������DC>���-�,_t
w}_yC��ſR��|!�)�x�ե˼�o 1�1ʹR��1�}��Sl�u��j����ë�#Ԃy��{�UZ���'$V�f<��	��'Q;�^�u�3��֌��h�,�\1�c4��gv_V���D߯m�w�Sqv\"������m'@:̥��ם����.��ox7��-�Vu�^3�!<����N��Jkp>'=�][�]Q0�D[R(T)�� ��	�d 1 �0#!�# �k�~}}}��s�|[S���ಔP���ߙo��k�������xֆ�B|,$p��EFF$��u-|U6꩖Sf]���L��@N�'�������zP�e�_A�6&����+a�t��B@���B(t��}���»D�����na��0��l��i���qyyx�(^�l�;�.ٓ�EXV~ui�9師�lik���#C[P���MlD^�D_aҏk�L�v�˫=�N�N����>���Dwո������A�O��wZ�r9����k�֣�����\(���z"�}a2i�a��ő��{���O�Z���� ]*�c�u��$]������n�:��م�����
�y*��(M��hPCh�j36߂��l�b��|��yFv���n�"�oI��Ժ|�f��#_�9��|V^3mZ���D��I�F7k|���e��S^�0��x�fOED�P�t�'ܢ�!ݫ�=��Bkț�ե���:����Uz.E5И��`$��|/a-��K&Үe�e�y�6��K��x��ȃE��}%Z��\o&n.�ݍ���Q��&�}�-��_L��7h�2q�Ț����2t���;�\�=�4�^���2�T��<�<�r�x�K�ϓ��m]�.��d�snm���o2_3���I ��`H1��c 
�@FH0 "��@���TRz~�A��r�6bZ�pˢ@w��70!��C�㏫��ºVf?ų����5���G��o��=Z��{d��M:��ñ�ƀ~�&N"����v@�
��[�[\��ےO8n�;��̇�J�^Z�a^�G#!����(d�M^�A"]>f�����0�y�����R�e�떱�P�����H�!Y�rn���@����Wf؝i�q\K��>'6���E�E�~l��j��xl�z`����ڑ��H��[�[�T������F�1��'����<�g-��M]���U����9,��)��Tu��|v����]I�	���sԑ&�6��|{��Q˵Kya����(c�i`�u���F�<[�.n�Ѓu�c��4f�u̔�6�AK<-΄������l�4��dD�X�t�u�z�!�j���T1��M���3O�ų���I��{ď�{�C�ҳ�����5���g�4��^�H���ӆ�OC�Fey
�"�֊��`�_�%a?_wj���~pI��
�G�5B[��YrSB����8����7tǰ-�]R���f�-f}��ؚ(hg��7��K֭�EXj�9ٳ'w>��d�[`�k��˺����S3J�З��W�6	�Kg򪪫���U_I 1$#DB � ���Օ��Lu�_@Vz%ɓ����ޘv�<�T;�X0{�4�쯈z猈�M��S���Z�LL��/��-S��c���	ԝ�B�h9)�^�i�6>�ь�J�h��0�wQ|��n�K�ƽI_k��xa��u#���M�rsv����=�Ը�a���u/P㔵�'�7��� -�71���µ��Ndx;̶�y�)���yx��+vSLtt6��J���7�i|�<�ѵĔ�v��[�`+ܘS�$A��uSG`*��>O�~�̯������5���~�ou��'S�g�Ҽ }˂�,�S�u�}��C�<Q�ȨH�Yy-~{`:Z�KE�4�6gmm�=�����L�(�o���l�;�Rm�*�KЫzU�0#��1B�탇5xŢ�BЦ�^�^���S�/�=K�]Y ��0�T}~�)Ψ�\�T{ *7c*�xx�l=/�T�g���C�Z�����-xB�{���E�4��a�}	�?+_^�������̎�G3���ܠ�+C������O��7W�oqzǔ�h��0e�����~^�����}�7I��]z�`�о�G��8!X�ɞQt�ې����='\D� ڡ�M��������H*O��{wy�jQ���y,�N��H<���mt�׎��̵����fwA	��\��s(1��%�#�ݽ��u�>�@ @bI#B�H�$"$�" 9���׭Bb�y�tw�S�'[kW��dS�B���ý����O�������G�Z:5ȥ��nAg�i��h�x��ѤE��,^mD�@N,9XA.˙�GlX�8fw�<on��X�әP�]z^Y9�ޱ��+�I|�NI������V�x�G�p��Il�w=77j_(yV��6�"0�ߪ�1��M-}�;ύ�g�����`��!�vYpe��y�+A3+�Nd0������F��2rGF1�l��בey���t���8���_az����a�0]@|!�-�憸;"eK�0(VAOX�#�p�;�%;�����{�&Y6q��Xtp|����!;�ly�.�7�=�p��@y�������S�[�Bqݮ9����2���v�.��z��˯
��j�n���)�W��E�Fv�v�@��/��4I�q�u˪���QcN�	������bZ$q�����z��Q�������Ra)2f�OAT�UY��^��5�פ]άd!ĵN@Αjkɫ΢�wT�z��]�q��
�be��S�`$0�V���]	�~��81��(�did�)��J��n�ݒ'�`A:���A����o�St��ЋN���j���F���U�!l��J�B��:&Ծ=1��(z�#�[2���է�d���%(��7K$˙-V�hs\Z��,������;�a�=G'
�x��5�@��,̜�)������Z)�%h�V
�hRR�ˬ[����Ry�qlE{�w�VJ���\zV[�Z+�[f,��佥�CD�Ij�U�יj�g�t��t�I�r���*K��@��n�˓�{�*��E/�@�h���7c#�]т2�Fj��"ެ�p,֪��{T�j���R%��,nb][ӝ�ތR����˽��QgN��I�&��gcY1�6��`B��c�i�D��Q�Xg��ɢ��Ӿ���J�����쌛�7o*O�v*��~d���ş/%wFϪ*�k�)Y+���C��;�2���3D&��{�X��r^����o	���Y;��hN]!4wbvX6��{�(�V˃�Od�k�� ��L�ޣCZ7M�lg\�Pܹ9֧c�T�y�R�7����k�l�%�W�^�=S8U��V�܏p�$H�B�C:e���#x�f�Ws�A]C%+߈�2M-�M�2Fjv��;zV
;.�;7�c���RI�;;j�
� ����ٷ�s�����ԋ�5]N_gr�d2�`Ӹ.X�t�=����&#� ZP����,����D��6ghV��gϩ��3F�p�tT��k���6*�f��m]�ɬ�9�Fګ���Y׫7�r�3�p�'�޸�:�����3v�H�{�7�i�K�Kp̕��)����Ѝhmh�K�Ϻ�š��`�u]��r����뉨ƭ��
ӏj����qG�V��[��־��Ox�oC��3��S�w
}(�G9�7f޿������[eG�5��;���]��VHN#�h>��X�2�۪��CCr�]�ۯsm��r�m�Ƙ添�"����}%��f_VɡaΔ7ۑ>��9�6�u������b�e��|�A�vY������@ӝNpn*�`v����G��r���g�;��pN�]��v��5����M̮��m
����Ю�[.�n�nL�+���Ƣ���=/r9Y]O`U�ɛ����d!�h��u'�e���V5U�K=5��Y�m��o%��ֺ'(�cǦ,#a��٣1������V�,��-�������N��+��&Y�K�ιK�|W�������H�
�Z�������|B�-i%y+���t��kNqxÝ�wM�n�rw6/u��S�9�;X�rR�;��5��C'����o��{%$� ����y�[2:ɑL釭d5k��
B�;h�WI���-�]K�����p��W�(b�=tTަ��T� F�-��4٢�Uґ�D��BQ!M+ -E�B�3�2c� �m�	�,��`�\�_�4���	�*�A:lF��F�eK�˭�k[<�D�Ac%- &���n�-,q)�E�����'�''���Yi��i�(�%�dR�L�Q��Ԡŕ���N�l����8��Ɋ.T~�UNj�4�TGM�ېX�S#�h�+�B��[g�6vzrpI�G���6�)��L�����4�V�[-���vvnp>��-h�E��F�b"�eynR��Ub�*���:S�N9�mȘ֢e.X��U*T*�,��J���V��i�G98�nYF��e1j�E"V���"��T��e"���<p�HҁF�Ub�KmM�塉Yb
fQ1�E��G9!ƵVZ)Q6�9eE���j8�������PR��̕%�r�v@�(i4��)l�a��n5nU��e��hr�Kek-�V�
_�E�f����V�ɵ�YmM*���,c@Y[�Wg�tN�LU�l��U�S�b����޹���k�Fdǹu�mu���t)ƅBA(��R�����$�d�1 2 "��A "I	߿�;�~��S]J˺��-(_L�ڄ�d�:�*}�ƙ���t�^qC��2K�Ys�V�6<LTF7(4AU����w��f�
��q^w  7	��ֲ�D���3ϸ��'���t��h���'mf�g�:Չ��iؓ����7
^C�(I�>�"!��?�	����:!�(ɨ۟{rq^R8�n��.��I�sm+��b8�ߊ�-59�4���zrگ_�3���a������u)�	G'*#[���|��e"�l	�Z�����m絝z���L�4���]`T�)����ꖫ�	�P*9�l(q��&FO@f�w9��Շ�.�vY���i�
#�Q{,!���t�)��'��uBl�Ε��5I3��e��
�x���ڝ�[!�#��= T@E�s��P�Z�W�H�dkkTF��&}lʤ��5�C'�r��]�a�30���b����9L�[m�8�"m�ǒ U���=j�S����#wkwJw�{v��~ڤs �3]�w</�b=�̵�D5��Y���v�\"���\"�m;�,
,mTˡX���c�{o��)�/d�v��ٲF��܁�-���)R3�g	���%��ѿu��=k�6/�5���"��PY��؟�U�T���tM�މ�M�,n���Zn�::��f�v�cs2���.��c�}|�q�����buʯ���`�!��$" H�bfA`���2��,��f>vy�d��N4߆#�7tO vr���	3�|�ѷ��wW���M��h���Ϭ�Tf}�T��K9�zt}Y��6_B��x��U�!+��T`�f�#�p@ֵJ�YkޝA����
i���Bj=3�aܚ=u�,^7��m~	���v��F�{�x�,�oQ�zу\���^J�PY;�% �
�m��*�>��j�� ū޳ɴ��ܝ�Њ~{�<�f/�����c˧8A�|K9�v\H	d��򀚖���of��i�I/�$stK��9���؋t
������-��J�_7[��H�QvC5��Q�ބ`R�Z�E� ����o>5U���AV�<27j����V	LN.�{W�l5������OG�Y��)����*�.�(�]̫S�Y��K���{��,��os�Qʰ�CZ�`b7"۴8�ٖ�vI���u��t��X��H��-�Â&%9�3���gf�s?��]3:�~H��q̕Y��.��ysEj��
i��*��K��#���m}=/}P�1]�vƴ��u���՗iE~j��#�"Nn\	��,-���{)M�X1䗜�ǥ�v�t��o!��V��w�0,��yƯ�À��U:QO9�{5�yz�0��/����&�v)�O��ג͋�Z(H�ȫR/�pf�y���R�E���GV�!c�&j��_}_Ϯ@�a0��	��"0�`���x?�w._U$Ϳ}�����!���Z�G�yP�|��\]��Uݪ�#��Z5��ŝu��z`��\ǝ���N������2����w����z�(z�n11����pJ��l�h1΂�锜iFE�-�����Q1l���x���V�D��5�9��OQM���Ҳ�W!ɏ%��sk��>k`���C�W����O�w����1��ϣ�kyabj�#�6#iO���]�)'{qE�f>΀�����KS�[:zx]�Uw^�$��K+Y8��]�Ə{}lBuGmSW���񆺨�H��ڍ��M��f�ZJ�3����T��b��{����@MF�y���.U�f�˃o��?�y�?$���ePf��z-n�3l�Wr��넛���j��|>���߮�J?1QtR��굥��s��wl熏�����s��^��m�t+,N��-�J�ڟ��;
�a��/ֹ�ru���~ ze��9^?e%��c�@�x�FE+m]�E\R}�w(m��źܧa���S�8�ո���@��3�s�(�9�&_�n��=[��fM�[u>'J}b�(�5��Al͔�^�5x$�w��e��lM)��MV�ԡ��=@���9��x;��՜�1�o3m6��# 9�]2���t�����*�L9���>��3,�a Ą�0��HQ	  �� ��̼]o��Q�(|V��d��z�7钟�#>D��/����~�s��Tj/	UV>��q�O� J_� ��4b�����y�lUQO`b�e��G�f����ԬHQnK����}ݴ�^����06�ځvc�82��[��|d<�Ɠ
�R��m�r�G\��nx����v��R�m(�X�"c���h2�C\o�sW�E({`/[)a�4�Ժ���³";j��V������q쎮y6}��NK�/G:�ØM�]�}wJN�A��{J�Uܨˋ;�C@���禲����T�����Ɔ\A7Y��sh�˟]��W�t�UN�cЗ�3<ޝ�U��*K��i���f�N"�����ӱ�x4�V��6����C�;BnB\�ɁN��a7
3�����S��\��z�r�H�{ ϝ����=O[.5�tlטGSނ ���������f�,Ք=�u�YW�ˑ����y�	͈��������������o�C&8=�G�1�p��R.��y:M�T�t�2ҩ������r �=�bc�'\�;G):�m�t�vv��cN�삏m!�oZ����t�oY���]��ֵ�O.����0_U*��Zhv옦�u�<�Re�6��7"��K�����D=����!f:}ǯ,$tq��ho�ݽ����0~sZesZsL��nf��� �F$�Ā"D D�f`�w����'&bӸrh��C����;�6�7���%�c�j�"Ψ[��E@�����%?k��=nat�(�?{��g��m��g�;kk|��	�{����Q�>D[�vE�����4�_m��%�Fm����(��iQSL��aZ�&�d&�)e���+�cH�}���]h�m�{]7>�)��٫�Qs�O& t �9�lK�a����W��/VbYo)��h+2şzw�t�KC�E���|�v�:��e����&v����
��F��7���z��[�bӮ��4F�*I��ȋ��i+�a]�q�&��rl/}u�D1k�K5��]�#k�#:�ڔ�<�/~y�|']�q���ܖ�*i�dS�X�DFq�rύX��Tp��w���7�[�u:Q�#g����:;��qUeźRSߔE'ֲ��h.���Ds�_qǳ�S��w~VHr;n�B���վ���J.c�ڙ�@����GhEx�\�;�-�bg͸�p(���Ik@YVl�u��Q�����c�ս��}/�DD&<ޘv���������>m�|����E�
�%mb��|�u['gf!�\T�,��G��|��:�}�0���Y&�M�m�H���f�-�\���𕞕�m�C�n\��|�>D1���6xݗ7E�eMt�]�w9Z+��V��L��� ���P�>�ΐ�u��|ǝ���瓟/n>��	��� �c$��Dd"$� ����nk���?&(�����@F��QN_�0<馭�J�f�6%�i���Ĺ\J����Vx�3��7�8D�XlY��j��%���{���k��t(ǫK:q�UT��Wފ�šFO6�W�z<�ۓ,9e��Ny��>�]M� �Ϙ�i��w_BoF>�k�tI������;�=Ck�W��`��[G:�'�#�~\�T�T�NQK�7�9м�oc�o!�����_�M�^�/�'�;�e(t塶iP��3�C��៮�NK�ܶK#ɷ�p� nr�j�omN�x�>a�"�vV�1�t��5�=zH"��9҃��R��J�@P�;z��\n�H6�Z� �L�޲mo.�{�+3�V	�G띞��VG�#|���۶��4��Be>Ǎ@�j^���&�m�i�w�d3`�b6��q����[Z�YTڽ�(Wo�Zf~��q�A\?\'�W�&�-l�2���DN�u���ջe�v�#��0���[��l�l�7�v�g14��x�0x�FL6����^��Gx�s7���cR�X����[l�=��5��ĊMh� ͗�����TԺ7ʍ�"o{�z�{�u^Ѯ�42�B����	t)_H�����S;�Ȳ���fs�(ljwsb!gT���V���ܵ.`T��c�#D�v��k��[��$��BF0"2H����3��ܾ���H��> �c9�?I���+��.N��{^�V�Z��=Cg�A�X%Am�]:Z�sc&��$y�=9�~��\N@&�0�C{_�;�>�R1�+7Cl܋ch����/�IU]�������+�Q�p�&�
�5����>jQu�<y.�ԁͯ\����ϭT���c��P���|���$���M��~�')��h�6�tU}s��W{W�������}�h�K0��)��w!��W�����đp��z"q��)�/t���ƅ�4��z�[�����U��2c��H���S9z���<�,���i\L�(cn��L���0�o�u.}dp�Ь������(����S�5W��/ؑ8�[�5gu�u�	O#z;''9n������P��S����q�	����<�l��pƄ?y�s�i��L��r��Y�;ϕ��2�/8Er�N��&Ss�;!s{�n�υ�I�CIU%�t\l�l%��нœS��^�V�T%W��Y5���܌�48����RFe�����Mn���h]��ʉ,�qrG�M��d�!�ms��\��=�;J���|9���
�sޞ�~�'bK������.��k�7+�Zذ�G)t�-p�(�W�n���C+�HfÝ���TR�L�H&�G�#�}.��9�c��q�w׭��/���}�ay���$���c1$�BD`DI`Dd�k�ϟ>|���w��<�oO��v�ad6;灐C��q��Z��v\5�E[jy�o߮`/��̸B"��!���l:&42��E;��[Btk�Z��c>�
���ب��Ue|3�z}U���y��@�C�#iz�j�O�B�	����5V0��1d�?K�m����g���4��p��Yn��M��3J����0��kj������anPXUf�������jWkY�E�/ܳ#�H|�X��n�y0벘��b�\OE�>g��O���R~*�=�.�k׵w#sd �Cb�g��\�3R�.♰����*_���q��da@f��Ti�t�OEE2��I�wV�8ѻ֍wC�o��x�n`9k�J��V��ϧ�9�{T�93�h?L6�o��U���3!sqt�n��Xg;��<�\���P���q�A6��Az�<i��
���YN�-��J8������ds�xS0�Qm�^+QM!�����-@������V�YB�h���k_%�U�]���L��r<�-�g>�\!�)�J�r	�Tٺ��.��8ߖc��%��.��=����(�̂�^����~��F��Y���N�7f���d�_��40��$"�2vq����U��c|�S0�ɡ�s )ޫ���vPoy�j9���R�s&>� \P����A4q�CL6�c�i�H�$�WZ�����$����a2H� 3@`Af��2��v6��l��������jxhecђ[��J��T����?.?7Z�.���G�z��_��f^n*z�����v@P[�H�p��P4ɦ )ơ�����֪�<�q-�m]re�ăv�k��za4"w ;-\֡'5�ڭP!RD4�'"z(�6�lu9�mN9g�4��j�,�/��}�$�𷽸����
*�ӻS��1&4��� �������r�4��nK:�?AЙ�dW:�'�Ħ�I�P�A%ZG�+م|��Z��nў"{�,^�m�CTkeu�.�.�ndk���Φy���0*�% ��gȈp�ֿ�l矻�U��د.�f�m#?g����z�aZ�\[t�2�k8Jh�2mt+U�n^�X.�[�\+�K��i���x%m)��O��>q�2[�ll
)���b�,Ĳ�	V7�UT^��g�מ�m���<C�
ܘN�Q;��UH�b��w��� ��蓡Ŏ��ژuGN;���X�Hw��%��hj@u�+�E���x�I�?���]xD�^����ֶA����/O64�w=�K�tL��q���
�*��R��篰��x�9Cdfj��u<�f+L�W�皯~����/<O3,�[v%����4b+�vp5W9�� f�Ҹ�fc��ּ����k>Z�S��#�_k���o�O��1 �A�"0�1  �  4D��Gh����_�������LKZ���ئ�r\[Pkj���;��M����&\*w��[z�T0A�e���#��+r�ܩ���S���BR���Tc�'�?��j{10�����vU���
�4[�Q)�G�0��QB(��ߔG2�1#q�znm����tl=S���!i��� �:�&"gLzpR%��uSv8X��Q���/��<���0�"������%	��|��X��(:��ˋ��:ם4պ�6߰�3�[��	��wG<���4f��l�0�HI7�1��^��ߕ���O�62��\�<(��r�ѝu3���Y��iyw&:u_uCI�ۅ47�y�v��wӬ���T2F�����D>#|/6)7dm�Szzq�T��h������q������@q�@��})�5r��Ԉ|�1ʈ��{�(�ѵ���N���K�?Dc�b�Y^�nj�����D��ˆ3�/��������\ʝO�vf��;_�S3 ���j^�v|V�3��/��}������LE�`$;� x��z�]�Fߊ?N�'0p�����ȕ2u��j�i��<�p�go��6(�Rֽ��ޥ�s��9����Є�Յo�Rrd��f�9�i�C����!�|�ìb�yvfj�� ���h�@�������ӗ!b�ץSQ/t�m㕪�^!t.�۔{��t_'�Oq-9�H���h�����1��x����b���p�+��­
�����[���}2cX�J���0�*a�Gt;Na�-D�������jB4��&M�3�>��ԧ�}s����G��`ګ^�Fl�ӛ��//L���]��|�p�έM��{J ��|�v-߅����:6�w�B�*�&�3�r٧���e�&%r�S��ѵ�M��ӊ�dr����'��P�v�u�vH� ����ý�f�= �e�K}w��Z�kL�z�d<z2�{�z��	*;/E���Χ�q\o�������˾�ϟC�Z�e	[y�-�I�����LoSU�B�㇬�r2M͋l��V�AEK7�Mw:�`��Ҡ{]��^�W�c4gŐt��Rr�E�����J����c4J��tI�ҵa�����b���F2�*�^�n�w�����&�ʔ�Dd��|b�=;ːuZ���<��˭�x���s{Ge[�.b3���q�S�B9峪�hm,�2�T�v���䴫��[���L���[����.�Tݐǵ#��/�v��ڈ���:������(}p��c*]\ML�@`��1��J9��eh���뿡�����YVH�_F��6»��@��z%�x.3�9�QӉ�15�Ư��Y4�%��՗5%\�镗s�z��Rޢ��3:�J�+\eoL���iZ���9G7�黎neL%�mF@�k7
�J�K��w�ico6V�ھ�Y�g 媗���.�*Z�a�h+5�f�Q��S6vT	G�)������z"4�yǓk1�Ԅ�H*���raꢘT��t�驧'L��D��;�re�Y."ցw�t{z��Ʊ��NU�1��L�%�)����ƺ��"���p٭��y�Ë��Ŭ@��md�Y4"[�z����)�l���m<����Tv�v9�ݸ�����蠥��X;ˮ_Pq�d��w.�յ�G+VV��zkLt�s
�� ��.�ᬁRڴ�ڥq���Ɯ�4va_X�\��ŜT��� .8�5�[�doq���eݎ\��SLu��Z����hV�mI�p��kxG�F�l<)5oj֫�-bx�[�5�	AG�g`njw�Ne�8U���fs�SC'v��V�1����7��
���Al]�Ξ_̡��#
�,�y-t�_eu�7m"�3��9�_���/��aQ�9���<���A��Хib�J�e+m�(�"�+!��H��eT�������������Ta���+Z�h�YU��3�L�(J����Y�Z�T�:n=����Y^8�+b���WC�*�h��q�F�E.\ɋn[8j<���r�̭q�1�PT�6�0Yi`��Į2�iP��r�3&NNNNNN
�%��T�m�%��o��EP�Vӹ�U-��1�.8$�X���ӧ��hYyIU0���˃RQ�Q+J�8"��&`XTV�T\j�3�3E:t�ӓt��R�n5�[F"2[)s3%�֤Ҡ��ZZ[��
Lf%s�du��x��g	��gY�v��ʵ
-�KV�d��r�Î:��S-�ʎ&e�ZB�X1����(�Q:t᳑�)i^5KEZ���ƭ�L��\�ED1*)�Ȍ���ji�\�JcD��L��Y�3(Q*;�1a�~�ְqQj)�PQeVW-�5�mJ�3(�)r����%j���U��� ��^Y};\c���b�-҅����
I�ݧne���V,�QK��{^���ϙ���p�H}ăF2E@ D@��7���񛾗��|F�**�Mъ���_ǋ�k�͊ؿz�U�s�3z(�Q��"~hGr��"3�5�7Q�)�����t��EȦ��^mUР�c�b�O;����K��Z!� �M77a��ҮD�P+e孅����>� ���U~���n��R�}.��`]�yz�Ǐg�N��+Or޷�,��:�$܆��U��E��=�.���}L�^���� ����X����+��:��Pf{�XxR��*r�-�yji���;޾��}�X�#�SW'���R8���T(d�W�/�3G��+�Ȇ�(�����hsJ�t5�rZI���R��-�(C 5Ey�/�.[��h8Z%9M�ِ��Α;ںy;u��4T�1o�A��3Q=ѳ�Γ<��R<.���8�{�\si����}/��n�8�9��M[��Ӥ�z�E�!�Jdp�@�Ke�wv�TB�x��C�Wj����|R�A����OJ��h��B���C�:z��NT�����>���%��TD3�a�C\����\�������[�6
�])�(��	���o�_`[{4Q�r��S#L�����vpH>f��`N��CM!c�6+�9�\��ķ��کmla[�̘S֧5�de8�U��_>8L��T�,�K8ն5u����s�׽��{�{��>�1�c$b(���,,��UU�������G:�}�%8�	x�ƫ]!��&kZ�u�^�A��[�ϦZ�ޞu�UXR��V�>��l��ٳ�(�>m��U�Z��0�34\W�ؗ�i�
��c;���[�U]��z<Ĵ5�ݬ�=���H��
p����n2�D���l~i�	=�[�<�{�ގ2�s}ۉ�3��M�*˥^�Q5���m�=_��L��Eڥ��X��T��}�K��h�v���֬��@=����o� u�N�����0�SP��zv�Ww(ddE)����O;�^;%��6��uM���Sp�þ9ϒ�+ߕY3�_�.��K��=��@�t5�{:6ޯ!P��M�
����!��#j���f߫>�%'�QJ��f�u*��bZ����2,����	�>���[�4�7�/F�5]EX]uX����5���y,�M}
���E)�-[;]b�!'�*|Q[B���ra�C9۾���G���}��V�רK���^M�K�e8�dN�&�q[,�)�Zl�1|s��2����-�a��&m�Y��ǌN��ن�w]�S�9��Z+ege�V刅SZ�^�����#�*�j�����=�}q0�v�:w0ȡw��uΛ�(�G�����%>�(vT��b<�k{	���"M��*�u�}��ou4#���5��9f���~H~D�F�b$���w���{��|��m��A!d�'��+�3�;i͙���X�Z��L=j�`=��N��vw������f}�X�j�-��b�6�5��ԁ\�\�PԊC1�?t8�/u�lEq��i]�*5���;q�o��H�؆՝v �+���&��HQ.Tcw$�6�	�b#��w���!�ب�dЪ���Y�����Tw8�*4�|<c���K��f�U�{V
�X� �
_�z!�W�A�z� ��*����Z�$=����Rڵ����j��Ż�f#��^U���x	ŗe�-��Q}�P�Y�P�G�^�_|�~��A�G�܅����o4�j,�)����?h�	�(�w��R�����*>xE����£��,�|����e}<o�i��xeN!D������,�S�K=��������}���3�[�u.���r`:H���$��K�#h�5ۦ=���B��P�֨g!��M��DzK>]j�n��&�!5��M\�kZvE>r�o͌kP^2[��]����vSe�Ŋo���U���%�l7R�t���t�Ch��P�&�]�u���D�8/��Ou�j:�΂h��<�߫�U��W�x��Q�0�I�ogVEFv+�24�a�������G���v��.�]ّf�W�+9�����1 �A�b0�{+sj�����'���V}i�����U,,�MxKzBmJ�M��h������/�fu|8w/�_~�M�-��4ƨq-S�Ť\��)J�mN��2�gSP��V�'ar<b�g�K
�2�b�wGt�ȱ(�01�w���G�`�d�%�K�ê
���9�(�;�xR�\�9n@�i�s �%;,M:�$��t"e�X�}�mipaH�]�.��B~RK�x�L8������YՍ���iֺR^2;��'��"�[�X&*�0m�,m����<eTqtE'ְTsh���	ñ�Q6��:�'&nϪ���|7��?~��(~�3�-3ޚS���{w�p�8T�r�9�_�H�z(���or,����Su��gA�
�P�_�7��6r��P{>��rQEG7b���b�`�v�{�u��y� ���N}cO�Z�?�z�;��ń �:ڢ�w����g��(/߹�rv���v����Í��F/��(F����@���h.�]J��A�]įr�+d����ޭ�tb~;d"g`�����z��JrK�/Ã*����8��z	;G�B��yRtK+�b�����j�.kw�܅��u8���	OV�%� �H����Mu8s�]�r&f��"=����YX[׷�~��1��E�����Ͽ�s�!M�]`b�X[?��{��5��,�C�:�D�/�ӈ���0��gv���W�⽏�"�����R�U�GH.dck_�ϒ��rx�^v
"j��A2s�Y]�U�ҳ����S]G{��E��̯n���<�����(�q�j_�ή�%̕꫽���^<���_�9~Ze���MCi{��૵ɱ��w:"J��S۹Uub���7����cZ����ֹ,�S�؍��,��%�5QL6|�O��2�0���<m�cd%]�Y�{V�W�1:�/�]�񋈀'*J��5d��%�e�*��?\�/7��2�+���}uI6룤����h��cee
��ry�.���>cr%ߍ@��sf,�T�3�5g/��gloJ�{�A�."M�	���ؤ����Sx�}�i�t{<]���i0}]9�ou��e͌�.�kb�tc|S��zT�{*kh^U��ԎNC�3s�_GS�f�/Px]W6pb��{�4>��dS�25�	����!c�M�}ʫz��\�ҝho�A�,{�&��622�`4r�kr����lX��gP����ȗ�ՙǹDt�\��W������{�m�G�*ͫ��)���b2���1�i�j�K��-��u���V�u����`�c�`^�Jm��^a�g�Ϟ~.�^�?S�#Q��b � �C*���Kd`�ـ�9
߼��c��^ĺ)�cX}��Y�G��\�cT��g���D�u^.n�I�����kͻ�$:���(�]P3П�9�/,cW8����c�MgWY}�1հ*��eױ!��Y#�sǕ�x4[��tI�a�=�^*���U��x��u<���W0u�*E�<�0�����<�\n��|S`&U�;�.�c�Iz�n�L�J[�Lʊzd=.5(��I�/M;��a.��B�H}�3��u�->k� ���}ܔ��z�ґ/躾^�'Y�^�0�0!��W�m�̠K��'s�T;����#�f}�=��T�l�C�Jሚ�Nx��{z/RM�5��E���u�Y転Ngs>��C����n۪�BC"�ӍO�l��͖�t��J�q�$H'9Ks0��2����gn.jd�\7m-,���lt8��cz|�M�ؘ�>3��NAc�
xi��z���dgwc2�ֲ؄
�0�H��cC� �-��S��TT8���uYd��谝���Uʈދ�f�5'sېtm�y2�~�Ouױ�{�W���E �+�	��Uܐ|7MN�J4�k�V�U���=z:1Z���$h�m:�*�4y��|emG�u�ٺ���i8㥲�Սc^��F����l٫�}L5�V=�/6��x��T�2�+��Z�Fe�5�K�G����1bA�dDFw��_�[����5b)˹#�m����̼C�>J�\���M�UЬ�j�aMX�b@���{EE��f�[�.�\Ѐg8���"���!�k:jm�a	�>�R�!v���3x��"㩱� Qͳum�4�`����p�>
K�=� �0��(����WX�uL���|�zI1�]34�j�FDV����^P�o/mF�6��m��)zc^Yo�߲A�m���.H�����M�7�ɛ�z�k���Ky���*ꡇ�6&���J���G�q\�=����4�'U
���ک��mH�L)*���}��M��E�n&�熙��"��t�n<I��MQ8�;�n�.o]yOg�u�2�����wW�0F��ПW� ���4<��y�L������6{���L��1�}�]@>n��P�vL������=�.�,5	���h�9�*k]�2���=Wl�4F&��08a�.~�臾^���{x_r��G=GY���V�=�lJ|n��Cl����ux���7��.�`( ��|�,�G����g|��	�����h9��I�3�A{/w������)<��Շ���
P�+c��V�/��H&�;��EӘ�헝x������^���4q�Hf��q�	8ܔ]��_8�����^d�%�uo�wL�zfJ]�Ð3v��ɫ�u�}��Q�b�$D��G���Ӈ� �\���{��>?L��6&�1�7�Ѵ���NO*(i
Oi�l�uv*'b���N�Щ����o��VR��*rN��w'�^���S+S�d �ȈQ�Ĺ����`���oU��s	�E�9C=���n�!��H0��D���R&��F ߫/aoO>=���"f���u9�X�)�z��r���1�y�5�P��" BW.�3�b�n�p������*Z�}	=	Bk��c�!��xV)��5{���F2����c%���g�B�s-��m5�%g���0,��Mj1޴�q��M��/SEMʷ�3�r�DW���~p����U��-~ݪ�2î��CJ'Sȇ�y���y�k��&�kd7J�RcO���7��YۤX"fSv�UL��[�UM��T^L
����3�1�B &Z��>z�=�F諮YáXb�FP��4�uE��tU)�����Y6�D�ky2~*�\��#�S�����������h]����gu�R��ʞN��N[�6JR�����&�Z֓D��n|a��M��ت���l;-NylL���gw�
Q��s���UԜ��R\�W8��7���*e|/��2�"i��O�)WM]�<:��Bf�G�k+�18���9T�m��v��o^WQ��%�j�h�}�|*�
�A��FED"0�����{�������<{�DB|j��בo��W7�y<��J�O~1ˋ��}X�Bfa��U��c��&5�J�c��]ho�>ߍ�w7@Lw���<��|��46�uν�>5jf�^��4�j:�<$	dev@��6"�@{X��O�yTS�Ƣ��c�E)�N��$s�T?d֢ڼ�3�?W�����4�x�Fr ���������"�/ͅަi��D
;���]i�ћ���dY>�	=���\x�����oom���y�ٞr��9J�*��Nؚ�O{�Qӝ�V6'�-�8�����qt1d
6e�;�/6m��#5?��-y�5��6�ԫy*�)F�ƚlLփ\hjKVS	(��͵��>�|�m�0jSr�;_T�^�;ѻ)�k'�ڡ)0���mA�g�Ǌ�g���p�f�ڻS�{� ۍ5���޼����z���"�z�}�|-�C�;�LMP+b�3��/4y��PE��<7b���Kbs�8r�\���(%TͯC�Kf��a��	��V�|�����X�������M��&�\��0���հ<�����g�=T�I�pV�aKb�o�X�x���.���,�T�HnG^�>�XKs=��UXC�\��0;y��MCg:4s����_ƅ�.��M�9[��jp�vRT����%�
`��S�s�~{�>������5���bF đ��,� X�@k��ˍ�IS��6���ŨY�d�`��m�� L�Sp���p�Ļ�\���3�mm�(�f���r�@M�#�:%c��˞��ͥ���F�z�[]�a��ե��V{9�sgyE=�蚜D�sD� S�90�®jO�-�Os��R����S%�&�
Ul1�*s2tӆ�h��L֓�=#/�.�5��SI[��W�|%�3ݞ��An`j0ZS�S�t�z[�E�՝��~�)��۰rz�H�x��a%�>K���-�H��v��T
6�q"����wR�2љ����z/�1���X�����da��ɟ�X�����=�+�E��nn�n��h��)��4i�<�x�oda���bx<�=$��T��ӌ(B�秖���z�HNt��Wo��ŕ��T;�c���1t��G6�!�먌;%�Wh����q(�q�ݨ����9h`������B������Hƫ=!��&����r�g`V��c׋��9��Yn����H�9W�"��"`<��o#�H�\��b�����ͼ�E�	�-�x�rmЇ�E��:�[�d�:Va��1���@k�+`	�eG��N��y��`=P2T�s ��3�)791|��d�;�r���',��R|��˧�5"(��,h�0<�2��ҵv��.�:@�:��C���Cγ�;��B�	�n_&b��^�R͘[�|.�t�eF��dvɴ:��o+q��+��y���on�
�%�U��7�������<��Fê���h�MF�`�olt�;��<G�16����|�;�3&^�Y�щ@5�L*��w!�K�$.��]=�0j�ZvBwY��l^E2���������Pv��K�����b����?�3��ϸj������Xā�X9X����\��X)*YJI�ħ7/h'�Y9� �����ۺ�-��E�Aa�u�¸��Ic��*ިQ�i�dk��wBUi��~�k,,�U��\��̓n�O�r�Ʋ�uN�K!�����^��b��⊂��.1��p`�kB�m7���/%o<]C�	�rQ���F�"ǲU�����ֲ��oB8(��]�=�wuoD��˩�A�jc�g��W2͔�%y[��%��s\h:ۗ.Ff�ǽ*K*�Ib\���D耧�V}�B�-���pW+&�b�S�G�=O�Հ�x3R�p��]�n�u$_]7�/��s���H�Κ�ٙ�D�K���h�s�Tk2�v��%���08Xy�Fc��vVg}$��aCp��ڕ�J�	ɚa`��m�����ȿf�C��]�c>�w���?�?�#dفmF�^A	�+�A|��`��֊���3nMR�x�U���J�b�����I��1$� �����gh��b�w��)`p��<L,{���sc;\��k5j�Hv�Y��(�^�f�v��=����N�6{,��m֢�*��ep̝vu��3�ۻ[ڐ�\�u�)�l��Zwj�gdw:��'O9im=��ǙLݏe�6�j2��9�Srgp��.e	CF!\���(X�j�VIWH�lSZՋ�y��=�ɵeKwꛊ��zr����5��q�l��ɂӵ�2ޥ'4:ws�x�v���kL<����ǹ*���*��ʒ�ۖ�!�k��5嫢@��Gv�듗�)�9oP��m���J�D��{��n�S9
B�L�9��!��i����Ց&oJx��2��t�O{k�e�\uUͬ�ӵ#Ɏ�Te;�I���쬕y$���j���9�RD+0��w�Z�1�;3T��ms)F���?;���q��]Be�;�Yq!���#k���yi�p�{���F���gs53g5�~]�ʷH�x�3,uK��7T���|%�s����
��E�7�X4�(Ѭ��GY�o��I��sv�Q(����ݼvS��[�tGc�9K��p9���C[n�c��xu#�-&��1���'�C���)ogPJE����F̸��aI$ؒ n30�e@?��
W���-�T�I�EHrr��ȅ� B���V�S���5��8'dո�LV9KJ�im�j�CW0�6�fc���օ���1������J�-P�X��S�rvrrq��`��
�Q��!��Q)c[(�PU-*�UJ�c&am�Td���rr/�*W�\bڴ����[R���˪?����Zʅ
��ʬ@�'�Gӓ��++Q�*���PZ��Df��Uil-�0�U-+%eYJ�f��ɹ�#׌��QT��Rb�[*��Puk�XZ1�&��")�*�ZZ�c1�<p�86��
�+Aŋh�����s:�z@j&�Uk�L�Vط-H�*Ysh&<x�ɴ��()ܸ�QeE12��+\̋nU���"�L��%ciV�<x��x����W)WT�0l�-�eUV)U(�ij#X�YPD-��S�:p��ʣ)K��+y�,�j�£h�TZ��
�Aih,�l��q��h([`���RڥT��,� �#]�<�ݮ�3P^�:پ˚k1���\���+Yz�qُ:%�Cz��)�\P`�]��}��"co%Clh�uK�t����~�����(1��"0DE&�����Ϸ�w���_�
�x��C�/�DX�b'~(T�a;������6z_����V�_d�N1�#I�{<G��&��3���y��ʞ4���ܡ����cKY���㳜�SЏ��w�Vנ��2U���5a��x���mn�$�ޟ��2<ڢa�O�� X����R��c����t�\e�f,��j�Mp�9Bhn��^�)(Ήt1ҥ���Y�J����-[�=#�\�M�Fz3���΋| �N�.��	N��V��^���~U"n�S�X�۵l�=g'퉓̄4�;�gG4ƅ�,��{@X�}�y[Mz���a1/xb����Cs��O3�㉙��y]yv3`��Jݷ�DM:;�/%�Y"%��3�	�4U*��5���Х1W�o>K����[G�Ȏ�^٤�x���
}��:D
��T��������얨μ3�K5�<h<���GV���ݣ*��%�x��I��t>�Vn������O!��%�-z�s��t<4�TO%tr�#�[Y�����2�|
*V���m�����C:\M	�n;j���m|��s�*/�o�2����Ǉ�R��]6nը�F�27V`.�1���<�%d�v�^r����)c��y��sK�K�T`~���ǋ�۫r�s�������k�v�#p�Փ8������͕fZ�MNB�v���׷� �-����������y�_3R~D�A$@b�f�t�JHm�`k"���<��Ky��ɗ��s�\�sS&�������b�0�N5����f��1�5Am��L���T{bѡU�B�N1t>?x��q�A`�Q�V:f�u�&�*Yk�f�\x! s�	�r�I����4(3�p`��P£��kwa��yB��!;Yt�D+�;{�p�ǒ����']f�y�m��`>��
P�&t�Շ� �YƏc?mR���R�3���j�O=W��T���� �yC>VA��6q��ꩮ�������1n�My�8�*�'���������X������#�GQ1Sd�Y9�m�R�p��jz�eNˢ�T��̋Ȏ9��EoD�w_�qeX�J�9�;�j/|�ȿ��!�v9c�<쾵q톨���u�0a�Τ�x܌�Sn�����K�`�E�-l���#ZF���9?�Fo�U�T��Je���%4P�!6�5iJcAv�+���Dʎ�~�����'�n^y���B�xp�GE̱�1ނ��_/�nW�e��a+J~=����uf�˶B}��=�Qv뀩�vgY*��i�3jW�kL���{�W��ty��#�`��F����H�����	}�5���A�@��{�iWy*�e�/;wU<{�4��;�9w�4�s�$P$�>����EfNq�����Ė��wB�]¥��P�@�&v|J|�&0ۣ�N6b��������6zh����,T�=��l����x���/!�Y6�?�UM���t۪��4��uNFp�-��Z�+;!���nx.�q�-��x�ٱ6�@ű���u���^5��Z&p���g���|u;
�!7U�ցy�A댢ၵ<���}l*9�(V�әZ~��Ye�A ���x�ݜC��[>����)�Fޭ5<Ωi�����ѹ�(A2�D[j���Ι������}:&V瓧ڎ'en.
�C\�"@OkAG݁o�� �0��U�x�p�l��,o���S�&��c����J`E�0es�����5��ϼ��S�Ƣ��ј�l���8ŗ������.2Mֳ�]�!H���x/�P�b<�a��-w�P���z���䞜����Vsn��%м�p��zG7\G�ϭ�/ܾ�2����X'��A ��?�k�aOS�93j�l:�X({��"Az/�O�|����8pgI�W�c<��<�a�1-@��z��V�zʖk��%�Ξʀ����-Ln�k�n'%Ήh.�9[���с���x 낺G���HJ8��R�p�)�I�"�*r�kF��z���B2�jPv��,v�T���䫯��=�͔<	7~{H��Xu�%S�3��0b�MX�����b�co/z�Fk�'&�ۄ]�a5 8%E��k'�{f���m�Ťw-� �c��N���\Gq��?T�=s�Va'4�Χ2#_�3���-Q��_���*�k����O�әo���R@��;A��E���>xo����9��A⠭�*�_yg�O��ٟUo4��A��L��������3k�J%�UDG|���%^^z�{�.��(�����mY�tVWo=t���jNt�=�ɦ�K&�r��+�:7Ul<6��(�ی>xqZ����p��Q{�oS�d��B���׳g��V=��!;�yO���aEePK�����P����ͺӄ2�WW����e�ioktAY �=�U����/�%�MY1��P���B����pK7�pB���pO�wR�R�,]����>����v�\�����C�����+���%�i�p���W�M�6^�������x�����]%��ѹ)oK}[�̸e�#��f�3�ʶ��U��dnc����z�s �_X��s0Ьu��toJ:�6���6�����$M���s|���mh쭎���ɦb��RT�����7,m]���n7��
ɩ����5b��5�b������n�������Aչ\Ũ.�V:f[}E��q�y]a��s.\�q���迒x;�nA=y�<f�φr�l�H���E��hFp�f�k���KVr��׈S�urN
��N�T��t��<��eA0ݏQ:}�Sl�����W��=�ۼ�y�X>jN�d#@��M�En�Z0�hA�e�@����W��";��ڏ8�Kz<�X*��r21l~9@�S��ic�#���=O�:s^w��=B��3V�B��;=���+z���}�Ė�wNl�1�sk���x?m_i�^4���q��ܭ�t6��k1
̈��u]�eS �p��$�t����1+*��>	SB �N�jmS獀�tE��\��k��N�sYs�DN��Yz��7��jP���)�j�m�*x񆼼���kE��ں��N�Jt����*����Ƽ�FL��VG���~ՕF���U3A�@�:��-B��ʗSD��*}��wi�a�J�}���w+&���5��	�MW���s�+����8E_+W�K�>�ˑZՐ�bו��K�Б�,���3��@w\�.��ݵ�Ѿj*o�V���D��^9�Ž}F<��7���[vpӝ��G/v"�cRX��سQ��6T7��^ʿ�_}�����RW���������H�\�]��qK�q�ֶ��)�_TU��E�m��Q�������U��nr�c��E�=�!p˚��{s��?T���)G������%W3u���B\OT��צ?~~8��� 4Z믻�aN��(�u���#�.V^VPŹ>D��^�kWwNf�ȶ.څ�Uޝ�q����#�2T&!�Et�8��J6�H�7�M�D���g��혆R 6�c������F/�Q��Z�]x�F�]O�,ʙs��V�%��is�/τ���[XpW��{n���̢s</�����;ss���M��J����ܧzG��0c�Y݃�bX e􋔡I�����ţ�Ay{<�N��j�fcM�-���Y�vސf��_gz;��8�KQ�����洖;ۂx�-!y�����Y������DMG<_=
�%:�1m�c�kk$y�����5��]����v�u�r7P�-<���f��b���#̬�Pi���P#�.b��Ŷ�ݧ���)�� �L۾��HU*ȷbP���.Z#�H[��y�7�j�1��<.�����\��%ވ��/M�H�9b�Sg�8�s����I��S,ryxJʘν��f�f��q�za#16n���/I�	nHl�ZŸjT�K���j�jY�]Ms�N��K����`�M���DM�\V������%��ز7jm`r���kR��g���E��-}�At3���!|����G`�aL��ߤ�`��em�v�̪q�+uU�	-q��ʖ��;�{�=}��"v�[�q��rȬ��keE[��2�a~�"jE,5�o�Q��.��5hL=H;��4�4��3��0��lӋ�1U���^I�֏�  ��5n�8�\/9���n\h�qYX;��j)�]��d����y���S�*�|�p��l��NbV��P�J���}�,{��$1��͢:⯷�3������o���|��~̩�]�e���d�i�v�c������P�Ka�m�J䉶��Tg�3}�J�Bws�S&��y�֛ƅ:�]/O���-ǹ!ޥ������t�Oa��+�Vڌ�\A������Z�1+�̏��-��g���gH2�~Xga�+��~ WXx��~ڮ�4���W�Z��)�EO& Y��M���@�ؼC5n$*��N���\q�"9�����k�<��ZZ���YV������wQ�_�L��ZO�$�ןP_��?�{�ћ�~�ԃ��r��𕛘�Vh4M�Fqw.ґ���Ɂ�cx�2Oov4�w��������x�{�!�Q���#Caqv����w-�3&�Y�|5�ٍՖ7�ޫ��;��D�_*�+�Y���xL1$�BV�\�`w٭�4�t�1�@���$�f�i���*A�	�b�LX��@��bt�˛Yy���b8�ǔ��� ���L�r�x�k2��T�w(ר{yxU��ۭ�slZ�@�q|����O�U%\��=��n�0��}M ��m�g�dh<�`mx~�G��~�uږ�:�4#y]�M����.U��K��X��O+*�xOғk:�_4Rz5��#+*;Z���K�+}� i�i��&p����e�ݱw]Ɩ����xk]8v��גq�;7���sMY���)['_U�W�ĬH(�����\�fd��e�6W^��C����ٗ\�;�ZPj �P������m�������Y�t�a�э��e�`2M��pSy���yҲ=��-Rz!��
��7�Ց�4�k9��xS[��o��Upķ��L�;ාF�f��x�Y�q��S���7q@O7@p�\�n��[��es�z�s���w�I0w�s���oBF�9�2�~�=z�ί9�Z�,�J{,�hQ�FA��T�D��>պ��B�Brz��;�G�z7**�f�Hm� �<��G_����(���=�D����q�������>���� ���;;��%��۩e�z�����7��Kk�M^l�X��̓q4ǩ�x'j�Nz�oǹ��[N^)�`ʌ�q���cY��x��Җ4��	G��9}>��
\"�)��<Tq��/�z
ovR�ײ�M����}+�j������é�'d�CpN���@*��V5�NUnAǫɅ��ɲVA�8�����soa�WM�r���b12��KZ����3�ū�� ]���yٺ��7q�����c�����G���RӇ�%�N�S�dY����[N�GY�#=U_tffѦ$�w��0'�l��0j#d�
�@j�R56�}�<(Ø��wz�b�>��� A�Yy�/Y��/:���S�����zl�lc:�eV�wh��.� �{��~���$��z�el���}��i]�;;&�Ļa��Z_Vup�@u2���ֺ|�5(����aG��ۣ��m�N,\�{�k�Γf��o�������$\��_����P��s��hܹ�z�ҒY훉U��=����Y�%�u���ﲂ��J:��S���4&�2�"XK�%Zen�+d{�Yͨ4�>�B��:���W^��5}	��O�.�!�wd�(��8���ƴ�M��ϸ�g��ߑ�s���K1��π����P�P)(xzz�w`I�;{��1����!�gj�fvX!�t�p5�.��F{���zβ@�=�mTu�3R"r��bϼ�bw̞�0\��l,d�2��m�`��hT����.��w���V`OA�pӲ6��P�[�r�A�Y�9��3��C�[�e�]�o6i���%�G��:7�n9j�]�Y�M��4n�n��f��|^p��f=��H]���z؃�1�2��c����$�+0�Ċ�ߝ�JS��1���hh��Z��V+a�+Z�c c�+����^g
l��fHk�rۧDg�+a�՝e�< ��7�`<�'��yJH��k������>$e��o�y*h�c��pJ����y��\,�q��5�.��X�a�t���b7���=����r��NJc�������%{ς�;~{WuV�h�v,ż������;O�؄��1.��a�S6*�MH����Pc�G�^����f�ug"Jӧ�������5����j�#/� �\�k��#M܏��3��us��{^�xƻ�ᦇ�r%�9q���q�ǘ^��oh�a~�$-�:��/C7m���t���61����1h��M��nkrJ��)]mW�R	9w��;��߳A��1Ǝ^Rwtv�±�����o%gP�V6�z�q��%2�"����2���]��+X�<�閛�x�3��t�)o�[[ �3y2S���ɽ7�o2_3�M���Z3�]t�3.�0�Ǖt70Y�����Q]l����G��bʛ�i�<��٥Q�MW@��H�m��`�;z������U�gSk7n��cW,;N�/8t{�(Wb*��:-�|ɵ�oD���͐�r�Y�հ���]�YέBVa8��n��-��Y���U�A��S��c�n�og'1�^��⠱�j_Db�B��Ʊ��Ӛ�d[�rݛ�����v���{rn�a-JJ�nq�I�eӳ(����c��WH\�W����:u�	�}3�u���:�Z��R�����2�A⁣{G��:m@�u�
�J���b�u�^��΃SVz����Y[��sU=�j'�P�ZÒ�}ёɵ]�}�ۄm� ��,����}C
�����8��yǣ���AI[W��>���s�lյ�U�ƶ�nM)n��𻧖.��Κ��fΗ/�e�}��Чmp��"����o\٩����C�w9�+�PE5�U��^�1�X�hƣ�܊��^wY�Rto�Ʊ��Лj����V��
}}��&q�����x�������wU�'����Tc$�>R�^m�a �v��;)�27(�Y72s��9��^"�֬�Sª��+y��K��:�^Csk��,�����u>�2�{ɞ�*�^�p�4:��N�B���k/'P�s/�7VW��eRs�f�7�BNcVb�n��۩JUʙ��w��{s�p�ta76�V��su��֩�ET2�9�;�d��"e�J���4�P�#r�Q��j��J�1&F�����
jɌ��>N�xʍxˀ�@��5�J[2�dD�hL�S"��.85�Z[2nvvnrN ��Q�1FԪ5��(�Z5��r��+J�,��*6��;;;98N$��PZ��ʧ0�G)nd�1ED:�I��b!D6ŕ1�l�̞������J$T��Ps3�)m��F����D&2�ŶF��+Q�8p��x�Qmm��D�eIX��d֭�Tr˪U�*#3V�(��Թl��4<x��m7��)Rҥ���j8ƪе�5*i+W)�>���Q���f.L<x��+�b����-R��`�Km�qZ.���s,��d�8p�ÐN4��[�[�9�U��n��R��L��[q�}j��Qg�Y�h[
����r�~�����j��L��k)��2�b�DfaI�\��"�hZ��h���){{�l��}����H���prw�=��+4mNu���}�:<{z0$�sL��㲊	��t{ޱ3w��v�k���a�F����sװ���.�<���j��Y�!��Ƿ����o�]W�����p��F��9L �z��qhmJ`u���CC�Ƿ�\�7��C�?tK0c�&�c��~'dUܥ����_��!��(�!JǞ��3{w���WՎ���Ma��Ӯ�>qJ����C)�3�	��g��Ųe@䱝+,`��_�Vy~�>񣓂7J�.�B-b8�d=�6�2-V�����#!�t5�:�O��Ȃ�찬9xFF� �3���� ͖�͔YCT�vi%���+��U1���3�����>�s�j�a�KcZ[9�`�3c��1|5ȢWu�p\�Xыm�<=F��c��\e\�WV��)�/p<],���T�u!����[^J�k�fV+w�PZ�����^��;�C��6\�a��隊�O߇BE����ɾSK�ȧ�t�s�^�LAX7r��TZ��B�dś�
4��Oo��;z�q�PJ��GP�����nT�YAaK��M1��_�f��
ĸ��r���^�0�ӽ�X�+�G�4x1�����}�hV�2������++	���=2p�\
i���W��,��a����uKM�N/VV��/[,�V��k�uLA�u!��K7���}��丆\K/?����$=���]�;{Q��/>�����(7�0�g�@~�J�v~�0%nH����0�i��Y��c/���3�2�*�N��t�L�j��}�a������o*�Q9�-@�E���XP␊�׆�O�Ca��5������l�*rh��+�ź�Ā�Q�����zr�{H�٪�i����p\�fMR��"���a�Z�]�p�I|"��_����{����SumHj�[�^�SPi��o}�ݻR��H���(A�"�a��cß�w����3.�q�)n�Ycӵ������=���)b,S-�?"��0���L�|�1�qM(�z���d��y� ��s]=83������O}c.u-=�|��[a�)80b�oC�ಮ�b�u��F�ds�8����K�/X��l��7ܳk����w���8���yy���]pk��oP�-�u���8��_J�w��5�}Qٜ�kzKv��������s��n�N��8����HW�P�#h�q�,�5�Z�tb�Y �f�ʝH��c��^��-
��L*c�v�;+�˪��� V.��V2AQs��O�[���/C�*���c+�ݮ���{jR�t�9J��hI`��1k�s�+�mO�r�P������3	�U���	+]iS��-���Բh�'�nsL�|��f� j_j*���m� 2q���k�ī�'6\tu����PB�v�3LL��n�{�؝�o����|,�y;�.��"[7���Cz*�ۆ���[�gI��Q�|ږ���o�d]YQԢ{��z�-�AOEѮ��U�e��C�4��5�y��t��O.��硹@$r@|m��96?/�K�������1s��~�^ݧQ�6�DF�"�h��sz�R��I�����ftix驨ȽW��d�ZyO�/Ȱ�.���a���^-���Rݢv|���7G�jBͲڣ�Q~w7�Ao�E�ie[�U5��BJ�
�h���)=�s�����/�+�͙��z���uIh����x�I�6k�hESn{��!�N�wm��.�/8��&��83�t'���:^���]��j�6��pJ�7�󝽏Ayh���Wדb�t��l�o�Ǫ0G�bm�Qܕ���;�V��4�O�m%�-�ϨK��Ig�qW��־tX m r�(&�59���ے�t�NE^��@��������Q�a��Y&h�n��x6��p���>�*N;p��"�q�]�i��P@��{|ߚ�G�I�"�����e�T>Қ��Xk�Vp5��Q7>��KdMT{8s6N�2GsX%Q��: =z���u��f>FN��!�GC�ǊSUݵ���N�?�)���0T�̼��L0)U^�4p��6�R�������}g��lgbRжƐ�|)nG��z�M�������)���ړ@u~�|Fq�S�(:�ǿw�옇�ӱ��Tb���r���։����@��iÈn�H��X̸�K��g�R���LmT�m^$�NY������g$�M��������c��C��c��eXwQA�B�f�+M�ӳ �S�~;�6"d�A"�!�c����7��J:�QV��(�t��]o:��K���P��C�������to��,9
��cJ�W&��|�e�C��R��MFY2�	x.��nh�o�O$�r��P�/��	���\�ϑ�՟��������t���r��������S8k����r������u8�.�N(����!i\�i�mDv�IfT'nzf��o_����|���M�Z�G�(k��V�nm��.�D�R�Q:���[�ާ��DVY��F�r^1jG��ݜ��H���Ԕb`��{��:3qo���H@㛦��Ωm�q\"�S�e@�/F��K;�O��T��Fi����u��k��N&H��XB\�ӵ���ó� ��jM]�鵕&o"u���j*5�=T�F�w-�׸�/��VP~�zo`���C�_��6;]�gk<nǇ�K̳�L5J��/\j�F���\B��ۃ4����,}�|��]g�Mήqp�|����T�'�����U��w	V6qŻ#����f/hwz�2�d�6�=�R�%`��u|⩟�o��V�$��s�'�:�F^+�Z�~���Y�շ�ٛ�#�����w���4c���zf�`�J0�v�'�R���pן;����E�l��c�δ��UnLh���90��MA�{���r:�"�6��EO�9r��f��H����Ds�03i�;��Dky��x���#~�隢jcf%���|U�#�ҽۙ�#p�%���e��QOa�Ev;�A\������Bc�5��5�0a[�}������Heekkܳ0]��xVa���p��|�wq�~��ݕ}f�#{\�@�+��[9%Q~���۱���DHk�Rt�m����M\�\z��5-��v���R�J�ZST��o�u��?h׏�=�#����_|�M��=h_���:�E�og]�n}�ٻw�܃��9�z�%1�@$��k�<�h%~�}���T��_o*O��	S����Y��]Og�uӵ%_Q�w݆XfzDB���q��yr�sH~�1�gF��L���Ǻ��HE��ٲ�(2��f�-^u�p���.��L����e��3���0]��h#J�E�S?[6���֪u��
[Z諔�k_M|Y��cy�P��
���o�+�g�76�.+�
]��V7A�T��c�ӷGjwXK̳��Vj[&�u���Ya�	�<o����eA��b��W.���s�<-:�nr,�]:��;��tڻ<��yj��
&Zap�{����^�1d��"���As}� �Mˬ�-��8�����fr I��v�n�`,�����{�Ổ��Vi�	5�*�����w�X��}���ƅ}wWx�Y��^/��=�V�S�b{���80��	���mP-׊�������[�8�QYX�lR����+�uE�l�zzG�L�m���>�@qCIk�pU�G*u"�2�|wq
�H-��I��׼���"�MR��5��Hd�T\�2�V����f"���ܦ-�)H�����ƾ�7�^�m`�Uh"̭�
�ªCwRy};UV�'�*n9=�)�0���0�B��wPKlb�Æְ|nK5�
���޼ޛ��p`����us�l�[�:j��h�Ӓ��j\�ǫ�`��7]��������rk[H�<��԰�jv�!mp@OoL�f%�`���kq�=��������q��:'X�H�FD�ga���)(6��Y.��}���P���F�^�:��S�9�N���-���ŚD����e�Y`L�L.��y͜y9�����u�b���6�鼼|����0#��x8wE+�y[�9�+_��{��d6P%(�/03uDq1P�}�0�DK!@7��P�*}�{���$�������xˍ�e�Tk�[�F?�8����~��׾w���Z���.(�gsJw���{}�z{j����e�hp�^H~�K�i��mj�|,�)��zk�t�v���N��v�J�n6�=P�W��{!��v�7[�~�f�泬����h?���#�zZGP�a��\5��6(�]\��g��*;�9����ᦃ�dp#���l�3[�����&_| �h{�����:%�N3s�����f����������`��gO����E����nk�ck�Er�"dZP3]�x^���A�KX*[�Z����S,��j��3v�u��SQO ��İL��u뾁i��L��Vw~P);+���0�R���I����Ğ��5�Vedo	��D��[�M�"�ͮRyXX�/h��ώo�`��;�>o<�m��EX9_'�I\7Z��^#0�G����2�� �r���^�UsJ�z�N����ˁ���l'ǜ�=�躚�f�1����/p��OƇ��Y��{5":bgapK+6ȓZ����ηE�!�:������U���솻�7#/ERJ29�vi~X���ܵ��0�:����{�a�A�6l��8��;�:�֣-w�w�ql��b��.��ig�衫�};C_����嵓�Us�A����1���nG_u+z�j�,2J��r�e�D��g���/�U{�?G���%v�o�L�Q�0j���"����uud��Ǚ�����*8wM��Z���ir�^N�[���q}݆�3�_�w)!���ke�ùَ[�2z��Y����˾vʻQ��W5�y�6��rT᛭$Ț#�<έ�[��#��
������UU��휗��]���'1e�01	�3p>�o4Zf!{�ODn1����y�x?Eko%܊��E�E)h���W�:���3���s��i�l0j/��.�}�Uv�����ΐ�/>�nwS�c���i'`u�`��.k�8�(K��2\�,��x�y��z�}��������9������s������K,D�lIS��0A��3�FNo�\�Q�Mɓ�.2痽Y;{�X�<J}r���~rp���s7��9ld3d,��7�9�|�w2��6������W^�E�� �bҜ��YZ��=ڼ ��\g,-ww�}/EU�w�J���<"7��ߏO�l1T�X��g�4�1�N/�Fâ��7�c��W��?��`����_�i#&���9�ઽ�Y=�<ռN�-�ùz:K����*f���vZ��z҉r����>��ߪ�ʿ8�P�{3�5Ȏ�t'#�:(o%�+��:����e��{��Hi�TZ ����}5��̲[�X�lz�8�U�f���K )Y���b�7m�Q�m�v�j�=�<��p�Ũ=~�� p~�hwJ[`�H߲.=Ʒ��\�^��r�n���ye���j�:j��]cl(���z�g�������k6�t��V]Q��k�9`�pS@R:�����+0��v� � xs����OΌ����)�J�⽓�d����Χ>�jһ�p�|�*PVƚp�Y�6�p�urC1������L����^K]���8.�ȱ*)����fY铨ˍF1���ӗLh�.��+��9 ;xq�!Itt0�ք�s���⡄����Z�Ա��%�*L��[)l����W�
b+˼�yB����e�o��*5����.ǹ�B�����.`�^�{|3��5N��~pd��lh��Ȩ��q|� ��[2��%4��W�THrdͰ��җzT�f�h�12I�:���
��p:�Xe����eD��Q�ĢX"m�T�'j��Ak[Š�α-�X�����j\�}�of-Usv�Ƙ|�>�FX�o���r��^������6`�L�]�H%�0R��ͣ/3�Tr��2���`c';Y�=άb��g{u'N�*�6s@�*��%�.�(8.�-���iꦍ���I��'�n�'%mZYE��c�p�y���{���B�;oU�TK��$˜�1ۘI�g����t�|#�(��9=���*^�s`I{7�m��0F1���Xݷ��9���˺�b)i���:$����3���z���.�%��@w���6Ƣ��PW�k5N�&�1�̠*B��M1H���Pv�u�F�1ո{6Ļ37���vT��2f)�Q�Vs��.N,*yRأ�]����}U�7h�u�-�J�ڼ��5u2�S�����KT��ulaAT�����@y�b%�U���kg6G�M^h([�x��Z@�[��Y�uP�}__*@:2�'i��o� cr��u����4n=:���6�6�e�5L� ��p�r���blf�@��	�|�Q��R�d�z2G����l��b��V"73T���9@��ia[�T�e�'��w�V�6S�iM����W�5i�kuҮw4(�,5	��n�B�
���3�!��$jݽ<��1sQR�n�	z�V1t Ҩ���������m���iJ�*��(�8��gre�`�R!��]wOPu��6fnQW��̣�bɻ�J���
��v�ή�O�q�
�.R0ػ�����f����#�I�'�ܮή�Rͩ٥�����β�I
;�8rG�D����M�e�0�Ô�s٘��qA���{�8�'������Sw���54�F�Yƚy]���㮳b�:�mk9��=��ݺ~��GM�P�-|Ԕ4��A��N�B���μT�j́m�R���#Q'��Z�v0Y�$ ��}�Cn���ƥJ1F�{�q��G}u��%BK�v�]ڰ���P��</X�7�L&�\�"V2�wI��u��6�=�/������/��:k�:�k&��l{�R�o.@�rhwA�p���ͤK	�=�MRj0�[{�6��.'[�ۏ{(��hqVZXv�oe�Ssn;t�4�ͻѳw0˒~�h�q)�I n#J0If ��?B6��D�&�����UE�t�ލ\�d����kv�c˥UL�j6ڠ�ij���)h�emZV�ejcUL�pkAU�&��vrpq�X��6�ڶ��es)K�.6T���)m.Qh��K����f2��fMNNM�E^Z�+c�V���s�
���f*.e\2�fP�DD+\k*6�1G,�L������� %�/k��8���F �"V�e��3��AN:��ڲ�LJ8�E�p)e�����6V�^8e��Q�?w�+!D�#]�E���B��\33�ŷ2�&e�.(��ޱ�m�J�)������8���ܳ�+qɒ�D̩���*�������fd�J�0���k���E��p���8p�h�����\J&�\�lGK�1F|�ti�Dw��4���#���".�b�5��t���E��Z��0��|�n5����m��.��E��\r�����Y�Ym-����1ZϦ���Q泎�K[mfl�ÓL�qT�2����L�����Q������r�
"6�c��oY��*UJ��ӣ.�R�a�����m�e�v3M���m�m֊�m5O�P�m�V0�Q\CxU4��YQQUZ��S@��DWm�7���k7���|5M�T���m#r�&��\�����d]�Ӯ�q�F��ז͸%�C&�r`�`�Aݳ�2����3���-��AF_�f�SN��m�Gw�O+s�bF��:���˲ێ��N��ݷH�k��3����Ā�XR���)O�hte�*��`}в�}�]�eC��Xf�_��V�5Y������"�#k�'��:+�Y
Ԅ\�l��v:&��,KZ��y��ﱗ�EZ�������:i�jYB�YQM9�=�ZZ*�j����E�@[SW����[N�e���=��w<.Sa�mF�=S�;�/�����;x�ol��EXn���ỳ���C����Eړ�=�w���,���������̈́�3�<�6u�8��ê�EW��mA+���M�N�o��z.�l��[R��Sl�l6) 5�����()�B9�9]�J��]f���+S����w2�e����T�A��Ӵ�yZO;Y9Nw;e��ڋ혛��l�|�M��\���x��-W��3%�"ĵ�)�d������Ǝe���p�r
]Vw-P
�f3r;�Mˑ��)�T��c��.�	Wɉ��n�x�^Y��}hK����|��jNE��ΚP헓�=�j�S}S̚�R�Q�5�(�*�)�ZWeYj�=3��*�ު��ў3�x��O'��-Jj5h����8�G�ήM��ӻ�'4^e��/O�F�w��B6tmPc!q�]��-���Jk4]Ǵ�q�x�w���$���y4�BƜ�u%���� W�q�L�^-�1ү#xJ>ۮ���=���Q�Cmד�Rׅ5؂'�u�գX��k�F��t�9�"����E�)og�d*����?
s�����xzzk?u��b���P��р��P+Kg�s�����:R�ў��5q��:!�*2L*0��g>�fV��Ƃ�t��(�����}�"��G��	�tE�s��޵��r"��0Q�-���?��z�Hț�@�-�C�R��eQ�V���YD�m��:���iԭ���Mĵ[�� X,{���|GG�N��f1qgm)۾�gnͨ�G�����>����ƭp�&64��2�e�t��'ϯٚࣸ���s�uzL~:`}� �J���l�t�� ��6�mڸl�I+�w���84j-�W���zZ!w���6s�ɽ͛�p}����`&�ݻ�	ɓ0+��7�C�|���ͣ1�Å��h�r�_D>oXު@xm���$�s�����Vh927��4d��<0Ì2O�5��I:��?��'¹��>g��?_A|���hgF2/ܦ9���I�NCw����	��{�j7{m5cǢ�x�s=l��}�NW���5`#��0Z��ixe��ȍ.�G&ΐ4Z���*��t��sNQ}��3ky�0��W$��5m���˹P�_		#xݷ��$����3ЎwU/dS	�tLm���	j�H�u�8�\]X��;�7�`^S�V;Ƕ[c�Uˤ�*T,����������.�V}yu����f����M�g���lfS_�jR�ׯV���}t��^*YYWf�}�;��_�������J��U�����vHԶ�s���o��o�|/�H�z[���+vĒ��`�o�O����UYn��K	���#;�R��vǨOӉ薁�R�H�O�6/.߻c�9㷠֕��t�w�uoӣ�F�쏺/�]u��"�W^�ҋ+#Z�2�6��C����o��EJw��+^#��>Os�e�$�y��'L�Vv�z��fKE��v��d��,Vu�*�m���WV�vr~����K/on'��:��dƭ�s���=�3�4_��i*V�,��r�$_�}	��˟��38�#�Y��}��WT��Д�]�+�����we�����*����c<wVYGa~:�D��ẘ-9�n�UR��|��f�[xv���b��P�+(�tm���7�����ڛDR��r�_v���琜7���h�cr63�e������A�DU}왈7�-�xs�Sf ��+X +2X������ST�8a�<� �[�z�O�.���C6k;�C��G���}7Cr؅�<#1H̥� �l�Xa�6�.v	7ild���ܠ�y�,�s�Z�u�Ϣ�0[��IH��Uq�X�YW��/�r�,uu��4���7��|z�t6��z�sT�]9�4]��V��St�����oT�Ag�]TY�m�Ŷ�Q.l
�,������!՟;�ѭ��Zw�PYGj��tz���ez���q �i�2��	�`�1�-��3��d\zst���LnE<){�Ԇ��
������~�	�s!�{�T�H�K�Ӯ`˫ba䝞ڷԕ��:jM�(-�Y���)��n�F��`˼A0pՏ-pf��n"�i4�A�H��? �[l^�6@��0�"ө3���E��:����,�N.�,ɵN⨖�W3w��6�FYi��*���n%�V&�ʑ����*W,���m��q�wyC=ٞ#M?�b���O��'9�9-�K�����c'�e�#--���*�k���e��z��+��ܽ����Q�+T_s7mWA����&�Pf��5zj��qճ�|������$��B.zz�8�� ��k`"p����\�y�g�*�tb�7ڤvJ���|�Uv�9�o��f.�*Vc>խ7�S�ҔF.�W]�)��{��
�ܶ�?����ct;�~2��&*��l�w��N�pǧ�JT*��aݫ���SLq��U�ū��j��zt;���km/�dy�hQ��2.Sa���XOVcmu�o�h�zZH�#6�����P��}bp�}wg-d@yW��=7s��5-��[(.��l���t/t�ړYW��V�sV*qK�Ә��FoM=��ilY$���?���fug�/Jʵ����x�hX���^�{#�m��v�5[���P�&�[nX�s/M��9�6гo�"甽�>����R�[�P 4��tFڷ�˽�Ϻ�z��:~�o\�L��X�7���
�V{f�i���w���!�*��~�7�z�?�4�^^��Q%��ե�8��Hd��f�%[6�0�S�1��6�k���:�|ҧ�@M���%�e>@����d%8�����2mB������<�]��d�藥Ws�/����8��[��6y�``�;�ȣާ��d�҉5~�������B���7�8x<�>\��ig�g�3�om��س��U�K[-��˔�%���<dS��&=��ߞ�y>�Ar�J=��sF��.3#D�B�aX"��$�!5R�s3w�� ^!���ڊ6�ݰVB���P���6�)ݠ<�a�٪<�Ni�͟AM���j=;Ը�u����ܐ���2���Tȟ���m�(�{���09wzW-��̈�k�	n���Yuqk)]m�-X��.��K'f���]�o]��'pkl��d9�Y1dP�<�6�7Y�U�Bf�+�RޠLv�(Y�'u�m	�Eb{R��,[�������,s�:����t�B�*�:<*�����H�����LK�5s���;�j�mv?|
�W��hpݵ>��DBF��ޚ�=���zvF3f]Y�tW;jJ�tY�#3�0w���b��r����;.z,�*WE�Q���_�Ml�wQ���f��t����������D��C���F��X�äoqA��ՊFbh�'M��{N���<svw�5�T�aY��6-ڪ�Y7����| 1/B�)�9�Ά&���'L�O����3��t��Nڼ���9r�K��kͫ&��U6_p�Da%��
�to(��ԋ����rmA�xnA�}[
���*�����ĝ�r7;e�e��q>N�d�5��Oڜ�S� �5ySUH{�1#��H�b�w7E�J�t�;+h��ך��57���,w�m��h����Y�q]Žڏ�3�C	��T*�⡱���ک��8Fz�����tB��]�E=���m�ޠ�P���E�OS,�ڸ�e.��pK�u>0ivS+�tI�2U]΢bǺF�����Ws
�9d��6�b��j~�ՙ����z6�{5���TeQ�c�n�,��U]Q�!��ɳZ�C]�ץ��L>u�jȺG��t����!���_�n�XI�nⶲE*��7n�+c�+�ۃ��Qݺ���'�`V�+�v�Ü�);����p�w�2q���>#ynj_v7��D����Q9�<O��薍ҕP�cKKJ春�b�N^��pI�PS�}ڰ���["9oVo�ϭT����j�阋����i:�j�(��E��Y�_��C�;��g���ƪ�:v:��j�+}z9N��S�vՔ`b�Fty��͊oօk�ZvY��̠�qLA�;dn���E����v@�W����:gި���k���zӶZ���aS��������:����,��'[���J���rF=�R?N�P�?֞�u�h�3�
��Hl������j5��	�q'�\m��_���d�,:T	��Ɔ��W����c��[�Ѝe�r�7��;(']H&F똟]�b�]A�g~��ٯ�0�c�d�Y�_.��^}Z2�>����Lۆ-X��E��f�/��T��#|�#��zu.�1�W7�M+.$L�N8R���X0����Os�7"8cU�3b�����_K�j�*l_@�Ʈ(7D�Xpޣȧ.����f�{�_����-�jr���~�nm�ή�׷5��י{��c�:�3���P���j=L�e���h:�˩��^�/93�D/�� � M��8���:p��zR�G����bf��X;1Gt��SZJ�l�U���(�[EfPO-];u�j#��Ύ�j���΍�������,����/:�kr�N���f��{��3��ϴf�M�3Y�u�!�QЎ�ة��|z�����9��:'�� �Y'<��*����Sjx)�?�+]g��i]7y�Oeep��^����N��eg���T8�O�7����g� C��GAB���#,��eD<E���7�(~�)��VQ$��6oVf�@U�Q�Ǳ���]{v���o�J�t��u�C�Ҕ#7ID�[B��ʃ��ɷ4�q��-��k���Ť}m�d�׫��dVm�7�����M�PNz�b�}J�le̩���w�cW����f{8S4f�+w�4CdG/U��''�܌�@K�wG���"q�l��N���Uߌ8�"�̼n�d�1��w�f�5�A�z<�}K�ǟ:dn�Y}����S�ٶ�OU!n�Ej�~�x��
�7Zj9�5fEʏ>�}�O.�)��-캮�D\��Ǜ'�p� �w�Ey�Cv������-Q�;������D��#fH��{�Σ�1��pi�bk���Q��gA��u����8me�ܶ��uykh7���[�qk��cL�a�H}���	*�����w�N�h��A#������z���F}�-����IV��ה�UP�Տ{�6��9��!� c��E�=U�����2J�wW����F�V���*��=ғ�q��Y�Ǻ ��k�<�]���k����^�����R�ɵ�CF���&�'��FݍƸ7)��L۴�q��fQ����"6q��9Um��A˥�pk�-8)�xJ",Jm,��A����='?�.��k���1n�q�l��lw==����е��t�M������b7��L=�U��6�u��!�;N�SS��'�桔��S�������W<�{�U�k0�P��8��5�0$����e��S"*s����K��8�hΫűS�hQV��Qb�&1I�7O:�ejv\&d�}�D嘓\J,|D�nd�Uү��T�PB��CV�c\�д��p��\�4�ҕ���Wmk�|WQЕ끣IoR��ή�S��ww�����ᔌPԣ�kNsו��{9n�n{��ʄ:���/sylm����ܨu���d_e��:�m�n,�&��r��>%�R�BGFQ�t�������r�A��]��.�+��PY\rn���,kɂ�jP��	n�Dv�w�Տw�����Jb��۠E����a�#������	+fqr��ގ�"���z%��*�dm��No^.��ͪJ�Y��j�ǂm�BP�Պ�yD��;�:$��떮C��SH��j0�\C7h^�J�R>���uVn��(��9���;�ӮûSE��:/��-�ܱd��(��e`�cs/;J���Y'�6Vhb�'m�O\k�	��i�����W�vn/�Ǻ5�ic�U���,��4U=��|�J��l��{�f�a�lt�i1�^i0Vv�V| �i�Vm���p�	=u��NȢ�.\��^-�_��PT0�v.�ؐ����9cF8"4]�|�Y�5�E���-i9gv`�-�϶�'M���#�9��ؓ����+���;��c�|&;&��=Q�}�m˕��w���-�;�Z��=�'X33�a�4
�W$�l��e�3B7t/�y�S��0ٍ���
�&��.=�O�e�)C��K�1pUɯ����
��ܠv����*�ժ�6�z`M��^ٌ�V��8��Ji�?J*��sa��u���;��>�-'E6i�ѐ��Dc;���n]�)�E�,F�H(�ҨyZ�'w'X.��:��#�Y7�lo�6���֦�}]�4���f��3u��a#�2)6䩺�4�Lk�6�\l�K��R�nk|�V��)�n�oD�>�YG��\D��b^���;�aڡV0HYP_?�C@w.��-ʁ^òj�`�2�jK(�.�r4��Q[k)�ٕ�uG�r}7��NmniO��|2G�;7�Z�ܰ�D�.31S��Qp<��j�q��'fY����Ʃ�uc�k�\����I�TV��G�`��P0�;8�
&���ep-�h"⸥�s{59����:�����&�����`VU�̮�̶�o#�C^0��U�C�-E���/�a�Y��+r�`b��m�����Y�g)��is�B0
�S_45A��MQ!�A+jT�m�W �m+\������(P�'��998�ּ�jTfR�cc
�c3(�����R��0Z��R�X�R� �e̘�ɓ�������Jq�?YE`�S\J�a�qz��2��Qc�jY��Q]Z�3��&MN�NC��jdm��U1*3�C��6��+v�DX�Y�m�,*�h�#5���5�-�#Ư�kwF���f�NON��q�PQR�1ģYE�e�,�Q��u���E5h�Xj�%M4Qƥ�m4�m̹2Ռcm��X�1���T0Çs;N�ETY5K��A�*,`�F�̹�9J*��B��Av�饴ճ:t�Ã�qʕ�3�� ���6�̢#2�.T)F���R���:t��C8z��)�(�mƍf&%s����Fe����� ��*��:b�����B����&���jѨ�8��ZʣmYV�[Q�0�r�D�MZj�e���]5�pL�q�S.Dʢ��Z1fZ�R�D[JQ
ٙ�4��h�1Z�Ԣ���kV�wqM��s2�	��@v�߼J%���{�l�o��H�Kֱ{��]lH�j�l�RK��a�����5�ϟ1�(V��}QK��î5����&&����}�n�_u���vJ���K �e�״ձLܘ���G��;�ܽ5��:(iaG��Kt�",.峋Օ�'�am��3���vO7�P�U�gM
�wd�`["�W��n�R�s�ݿ��]YQԡ���sk�ͬ�Ó��/�j��.
�h�ʇB�E�*�7�b0��P*ko*�^�l3�f�d�9�@`Zv�E[�6���g�ߨK��;�7v���Qc��y��5�*Ȝ�;��n=��� �S�w����Y^�����7�L?l��%�}Gv�{��dSd����;o���v�@�m]���yл��|Cɍ��
�	�G���J��[�sGڠ8�n,��\��'�'��GMLIq�Ȥ����;���њ2^��
�.'��4�[�����|cg�!�:��3�;����w�)W~��fz�q�-Sd7�U���Y4˺��J����w:4%<��J0���;*��.���NR04-�̣�#�Xjb�GKg���$�e��i��7�L���Yf �V�%R�G"��}�｀e��f:���G.;�f#+`�mp��Ēa�u���-�/��|�{�Ǣo��2����}��0d���96�d�*��[w�xw���2���~О�5粗�j�VM�*����ծ�Lm鲛�7U��,.����B�@����<5[4j��fC��*�����!��
��j��7���S-Yz�a@dr��mz�؀�~��U�tZ�$E:����ј*����v}No'��Zr�Uu^s�ʆ�:R+c�Ne�J��!��K�.����pz8d
���t������M*�?5�on��m��mO)�Z�B�w�E,�ꂺ@�Y���z�9S�Rp�?EVE�=�yL���~���a�l�V?Զ��z}�	rfƚ�+���L�J'�g�w�/'hݴ	�${��d��>Y�W^o4f^Z�W�R{�����;{�����Q+�î��g�Y�C)��cU[�������]xp��G�,f�Y{o�hƆW?}~�����`��b&��o�Sw�yZ�u�5gRɉ��:/��ՑE���WB�7��O;g68c�"oh��K���#����RTl�^h��zR�]\���m�;�f����d���V�af��u9$.~�EPpFh�I�螎�w_���2e�eL����(�.;�W����WQ��\�]n�P�.���T�-;�\X>�N��Z�3��+o�X/�hLvf�5��+�5�B7�H�ZڋiE����3��H�P^6"w8���A�v���u��5Ôݶ�<���П�x8�f]�o�_������+kNY�^�'�/ŗ����ζ�z��Pb�|�x�ŕ"��4���P��w�*����ƓO��V(t��>G��$B+"83�}9Dv5>5��xk�9���~�B����X=69!�e�"F+f=,��-�^0A�u��0��כ�vb�Ɩ����ڟ
� ���+J�����)��S>�K�s4j�p3f�jI�c��R�5+�TX6�ej=&�mn��g��Q���OA�u�b��w�C���4��U�ʴ'V���G%-�.&2j��[f����d7Npe�E�>^�����Le]!��՚�/��p�8��܎m����k��k��`f�xX/���rp�W�C�\������\�n�̚�ݫ��0i�ł<O#�]���e7e�p�ץ1ޭa����m��Ɩ]_�{�|����C�m�u=��E
���iS�a�i�-����L�a��nC,�D�v�#�;lv+��wf�W
�Y{�g�NT�ˉ)�9qݥ�j�O2�����9�,^��m���r8Z[V��J�A/Xu��{=����7���M�#���a/�,q����R�����:2�}@�E�o]��C\�F5��o�����K�w;�KN�Rح���k�#�+M\�nR���45D]��C�"x�s+��w԰L���ԫEv2q���Ǵ�A5W�o��{p8�����|�"���/��m�����fV��껅����۴�O;u��4tg'�GL���cZJ`{2�un޹�1Uꗉ��9�H~�s�:��bow�5�Np�g�D�5��䍘lt�\�$����=���������[�Us��+KW�H��D��(���xǈ�O-X��"m�l�%��漓+�T� ZX˧��o�\�E�yK�B�É����(w#�Օ�ŀ:�7�WT3��K���Q.+{oL�Z����|�;�H�~����v�����]��e�}J>�Ö���[P|9g�7���B�,����=|=�Z9!ru�IV�rt�p��L��g�d竪j��T�)�&��%���;#��.b;�=n���h��>�L�w[�\����U���Θ�J��m-��+)����V����~��(=EvV�yR����k�桺%r*��"���ڛ��:M˒D!r2��mCV��Y��㊶�W�VC���k��O)��֘�ّ+�j����cd?��K�.���%�.�)c���uyvc�N�a��*��ou�GP�BwH�ϭ�j��0��_�IJ��+v�Y *��n��gӝ��sVǵ���ʅ��C>��@��+��n�Y�ƣ��KU�2���-.�g��mڮv�Λa�}�vt�~&�(���ޥ.�������z������5s�A0	=��-
�8��a�e}�h��h�29Na9}�4|b�?���:�8�bFw��mk��r�
Jȳ��;����׃!�]	�?�\D�ݔ.��G�y��bS�˛���5���غ��a��,�zR��*R�{�Ӯ/-Da%��e��u S�f�b���*�]���~u-�<�}Kv�Ipa�ǍF3�Y����	���8G�͌��md��w��%�'�E��_��=�Y�Q�
�r\'f�L�i�����r�$��D�$�z4!���oP��=�7��*F��1'�~��D[�v]Fp�ۍ�]��E�qn؏�ee8*�
�FF���?����쎝c�ׇO<`�����69���[�\Y8�S�u5
@U�ㅐs�K�[�ך>���de�&����*�g]Ot<{=�[���JZ�2e��(������ٽ�XFGr�Q�l�Ks�&�e=�t��!�E�̛�j��#%FvϮ�x�̢�'�$�n���b�~��U[=��	YX�&v��n�F��s5�e���|4�ڳ)PYy ���s\Si��!���<�$�f���%vT�[,8�PT�t��;uқ��ݖ�4���γo贸į@�s'�N�`���Gj~�U��t�H�<2�b㞬�4_�V�8�i�Ni����͇k��`���qu�[��2�]�Ѧ)�r�+����r�>��X�aƅnMy���{uT�I��xݵw$
΂:OT���n�c���kD�%� ���X
\��H���b�E=Ni�ّ��A�=$���?�阥Y��0��?9[d_����G�9Q����+~����#��&���l���������-�h����yvg�W��w�[�ܝ���V�[�!��>>��=��B�\y[�,A�lg���D?C�;t^8�w�:��)6��[$hv���
��t�7����L���#B��&��r$S�)��Ֆ
1��k>�,]��*ؿ5�瞶����F���h��h��y��J�+��U�P:�x5	��{�a�A�D���W��T?�I����@��MI�9���s�����~�>GK��=�"�|k�́w����KǑp����>�}�V��e���us����ʹ�-̨>>���z`��8ѐƃ@�k�>;��x��1e���!�������G[373ˠ��#�W4�k̻nb#�C��A,�e�Rws��eyw�"������nX���:t��D�uÛ���3�i����R�� %�b,��
�)��������f�:���9C�Q����U�q\�`��3y���Ԣ��zX|�*�IE,��j�z��.[Y�ga �Ž�Zi��R�7eKݳ�t����'[O�����V,��,�S8�D�W$ ����<z�H�l2��Պ�r{3q�<�Aj�x�^��\U>N��@��x��%s����Έ�G^<&h�ȯ�����i��勃���d'>V;�]�Q�Uo�.�l恑�S{��������|n$��t]�^Eޡ~��{v�2Ն���$L�=m�E[����F{���MZ!4��s�U�����g�â�m�T����޻�ġش���)ʥ�c���r}ch8^@����q�G�<����oƲ$���{9��o�l�������Q��Ɓأ�<�!%{B<�j&]�T-�WEU�d4�)�/���dR�#�L<�W*#O[�@%[S:y�V�[<j�S�sL7��/�]�`ٓ�¥�=V�Z���V�u@��N�Ԟ���;���e&gt�n5BQ���W����O%s<#ϰZ{y`��U⤶]$P�*�5��Q���MꝻ��PU��+�T��E����Tvm�*�Dׯb�b��q<�Z�%b��4��4޼�S��G�s��
��]V��#�-vm?�]��N����{��Җo���R���#��0A[�5�nC�ڢ�:�¦_Nl�l�7uͨqMD���COw�#��0o�\}~�=������t��C��i�:x?N�I���$�l��Ot[~��{`0���1CU9�lqw-#��97H���+��m���6�z�})��C���Y���R�ǭ]���q-c1�ja����y>��x������?gf'��/�O�]��n��h¬�On�#�y���.��	9!���}%�i[�����蛫��g�Y��{��1��e5���R6Xo�r�fB1�W����c��Tq]:Y����7pI���͔�l&vR�7�,�&|�z�1�|v���ifh#����xr�b��*�
��OЕ���"��� y���r�~�d5g����ޅ|�z3�����FI������Ɗ���>5�r4nfOb�أT�g�u�W��Tv{�BK�q'"pI���Gu�Q����k�����o���ƽ[�i/
Q$�ūkb�vG�he����N�m<y��
�Q*�"ܗZm={AT��!�7y}3��7�}����mk{u��:�" ]{,Y}�k{3^�â�v��m�2a��J�:���d�T��x�Fqp������k�w=R8@z�J��i)Yy;��+]�cyx��f��q��b{'_�B*�_��)t��p�빧�|��𼾍�E�65��g�r ouX[؀�ຼ�^9�w��:�:�{Z��J8[>e�
�ԼVU	N#�5W?F�t�:	�o����D�!k`9��w��c�U>�yD�,�<F9�df��O��ՙttY�7�m��oh&�lի�0���swEt�A�-J�:��`-W�����yeZ����L��a[6E�<�ff]�jzކ�i��H�~qײ)%�7y���NUkU�7x~Gx���biv={���$���iZ*� 3�Q�AP�����^p�/�{��7*o��q=��wyS�fn}��:�Cjb8���Xs�8R���l��
�d��3�����[6�hD�$o5�2(l��-��hu�/����`>����?˒]������_�`����G����$��v! �ٳ�D%����I �BB �A0C���B@��� 30!��q�������I	���5�I�!�@2 @�`BJd  �  � �  !� B	  � X� I  � !� ��a  � E� � @  �  �"D� B  A ! B� � H� $  (� B(	 #� 0�B 	$�20$��@ b�P 
D  �H�� $XȀ� �(� ,"� B"E$ �IH!�2FA�YA# R,�(�"Db2 0���AD c�A	D �B�\���s�S���@$$P		 ��"*�`-o����/�
����������-��ߧ�����<?+���s_�}_�B@�O���O����$��F��"�'�'���?����(�~��@�hHBI�������&A��?��C��g���������C���-��� �$B� 2 ����#  P� �$c  
@a$d �AA A`0�DBBE BI� H, # �@BH���I$�  1� $ � �B F� H� d�@ dI   0@" a�2 �a$@��	0�� $@A�2 �� �B��I �2@d@ � $�,�2A�� a b �!# #� 1�2H�@!L���I������B H� 
  � I�>��?��~�C��~��O�A��	 I	&����?��p3�?�P�xY����"�某�$���~��������	!$���$����~ؓ���I	K����H�N �g��P�����`=��C���p�&g��`P�$���@�?���	HI?hv
?��?pW�?hk�����������RHBI������$������r�a����?p���a����Mx�{�ÿ�p�$��p�3�?|,����n���^��>���O�!!I����ɽ$ I+���S��7���&�a��(+$�k>�[��l�0
 ��d��Iw��%PP�R�P"�ZҥUT�DE��B���I+MP������2�0���fR�B���U% �U$�֨jf�j�m�ͩ���PFY+X��^�͚�٭l��ٮ֬ضʳaU����bֶԭCb6���c3[5[�갲���w]NV��l-�����{��P���Bk�ًMQ����)4S@ڵ�6�iD֫�Sjikс�Ͷ�+*�2�$�iB�(4��1ikjͱYJU��u�
�֍�ƪ�  �>��aX�ݠ M�ݰ�!�t��������Wl2 ��̀�������֝�7P�iR]]��KN���mR��J��U[6�0%�m3f�W�  ׸��4(P�c��}�G��(hz({��ol[
=��P�CC;�ׇ��ݛ#���h��ւ���孵�+�[cgm��V��l�f��6�[Vkt�%��"���)ͱ�6���   -�<j��Q5mkM[-��ܭb�V��f���û��m�҅��΅��c=wE

��e�SU�iE�,K��KjX� j�z�U/5�&@im����M��>   ,{J6�[W��"j�X��k�Е4��ڥ�캊�)wu:�u�X�
;9uR)�q�UJ�a� u@�sjm�3[M�v�e�Z�il�
�   ;<5D������(^^ݹ�"�m՘�lV�+"[P��U���X�$��Tj�`�T�@[j�8��T7��jS7vUՍ[5�*���  ��Dn]Ҫ�Ub�UQQ�uUJ'FP(%�R�ӫ�.ڕ*�Y�U��np�nE��U�`�U R�4j�Z�Z�[-x  �{@*�rm��R��⢔��R��CK{^�I��y]��I]ԭ�J����n��"��{�QQ;��W��ELw��5i%[Zf��m���c_   ������=�w&�R��K��h��ݼ��^�T�oyURHU{�M�)@<�5�RBIQ�9]��������י�����y۬Vتٲ�m���F�>   u�
����x�/F�bwt�UPD=��)#�y��PECt�ނQ<�i��J��rw�J%���m��S=z�%�9洡!a��e��c�ʗ�  ۾�H�%+�{7�R��瓩�)E	���)]iTJ�z�<��UW��K�)%B��)A�<���*�#=�zT��w��*��J|���R� 2 S�0����� �Sx#UU43P  E?��  ��M���J� h �)PLUQ� hf���~���=�/�����MΞ�^���R�h�������`�������������ﾵ�o��1����cc����m�����@��m��������������K���դ�����U�*�@���ּL@�ť��oV��	ufB��, ��̚ԍ��ht���v&ںi��^m�&EkRn��Pl�Tۆ�� �y�C1CMx��L�m,Vea���n�6ij9L;�Q=�2^�gea5�
;�4ƸQ�~�Ъ��쵱:;P��5Ѻ#A�aH-D�Ű$)Ӡ��/H���1�H
/q�YkX��L,�[��0ݼ*c[j���Z�w41A��\Wz���N�o��ɘ�tiK�v��0Ex6fMϔ���JGM X�%�]���^�Y�%е�ъ���.Fi���;B���Q^@ �X4�g^	w�D�cQ���p��4,{�jH.������:
���^Ѻb�6���wiө5��䂄�&*V�bX�YQT�*�<�.x.�"��Z��,[��hF�:��9;̌�g4��<����up�2]]�Y{cv�"�7,�ʍ�y��M�Ѝ��mɏt�@k�Y$VQ,�0cW>QO���{ٺO�4�d�51��[��n�}ڍ�z�"�^��ֺƮ�ch�m��W�-���6/v�<GPY���aXh��X��겋�>U��fQ�
-ɲ�q�9v�8r�J��އ�l��!m��7i�f�"���
�qU�"a�q4])ydV�[pR���R��`�n�D��y�"��4c�b��N��C0n�.B*ֻ��Sw51"�����ZʬR��cF`�J)ąK�٭�QƝ�77S�4Mӓ5��+/n�i񡔞���������l9K[YKmD�c����xp�ONE����5��b���ʙ��`Y�h<��,Ս����yB���f�-�.��b�VƠn�y���qa�0�h7/I��If7ۆ�h����A�B��$�{��
]�'fU��E �$�һ'E�R�+t�6(1��������f+U�e디�90;u��%�tڣn��W���EGe��A��Zljn�k���n��b����jࡖ*� �f�k���c(�Ԕ�ڑ�wM��`3RCuú�؋ם�f�LKb#�طe�"[���ݲ��l]�)���e�Lm�Cb�
��@2&i���>D3�T�~Q#�m��S�R��D.�^�wXa�[ئ��Y��	*�?�!Y_c�[��Lՠn�fk�NF��z+c��{Of�*�4ά�ҥS��Hīv�m|�6[�8��$��d�
F�lǖ����E@���Yvw	֞���n6h1��#v�\r�"d�����)<�XK�Jݻ{i<��;I�Z��	=Lh(T9��VZ�U��d�e/�����Y��P�[��)�n�`�ܘ�CU����ʚ��Ht(�L�(�;wd:u��<9vW�̭��4aB�j�4ta`c�L�8��m�à;�ILոt;�Z�Z�(u��wR��͘`%u,a=P�KU��[��;&���;۽�
ݥ���SP����K�D�v�5��Uj��$��a�t/D&
�)�L��Y@D0�ou�u����ueS�v@��-��1&X0[�LGb�wu2oܱ���N�5\��(�x����T~�f�D����V[j�^�K�V:����+-Vt�X�%�9��K����1U�P�!
��dD�T���򒘥��#`���P�yZ���@��׭��F�И�.:�=۵5<8�yb��Dw�ԼT1)Ӏ����L�\��մv�6���D���(�9���Vb����+^��1�A&;g-�oj�)��F��hWmEB�@��+�s\ۺ��q�3)Ҵ�>ږ�yB�ˣ-�^#��R�=b�캔LmX�^+�o4,�x���%X�T ;d�,#1m�) �S@�F�Ґ������退FQ;0ܽZ�6\w,l��.�5SIt�-���X�����\���wX�2�Mx0%������ۣ�j%�xt��\w�J�H��oL���q蕁	&�0�l(��9J�p0��I��0�dMX�Gx1Z�Ra9�� e�NI�+Kֽ� �@����4�C����f�}�	p)��"��7Z$��ź5� �Yej�\x�ѵs�M�c!�Ǌ�ZM�Å+B8�ѐ
�B�t����@@r'x���nX�@z�
̀]b�2�t]� �xԘen܎���?A�I�/��^^R��fb��V��m0[Ҕ�{��>���%��)),���o h#�a�-RnVJ)4�V�ݿ�<I���S�ʻQ;�hK��0�R5&hQ蔕FN��x/���a�&�x���ñ�{�0O�)zvJ�+F�%[e3�5���0��jP�@��KVb�2�+����� �/V�C�XK� �bL��wSh�Ϋ��t���9�H��A䷇5]�%�n�y0�<Ϛ�,��li��^⣶w5\[nn[O}w��z�S+ k&�FL�t�%uĖ��JMԢ�σ��n�Z0i��P����W6�4�֣Zm[�Tn��c&�l��qfAnJ-��m���@�N�Z����"t�z��hS�/5��9kE�B�;?��+)�"�"���x���=X���an�D�[M0%H��e��ҫ�7Z���H�'���݂.�X�C����*�	�)!�.�*��vV�dX�'n�6�T����y��!:aR4j����7#�MKݺ�q*��1�k���*��u�Ff���z��	f
��nR������k����Κ]ӃP�[�	;����g#����yq��u
[��YJ-�k&VkY�E�[�"����n�%��2�Fڼ�7r=��1��r�[�7VRi�k4-�a�u�2�O�D��t[�Z��Ͳ(;ܬ�,=�.@���e����r��5y�k���h���s=�� 7S;P�i�910�mӯ���ٚ��8ҹ���׷���cp��;J�ݺ��l��F5J�F��u�e=��' �1e:ٮ�a�F�d.Pe��l�F���� Mf2��IͅEx&F�C)�[���o:��n汸�j�ب7��cd{�0��vѹ�3 m(��L���7�$�s0b�X�2�=2a^b�2�X�I��m�S%`��BSpTf	�tL�i"��n����A<z��mF�{��YAU���.)�Wy���o�2�}�H����^�EǣNF���"�b��~�=̼�X�k(^	�H�B���7j�y1�ob
8+2ڀ\Ǯ����hf=2m7�1-��pm)4�V�V˺�,���6dCl:z�\�j��G�VL����V6���!j�`w�a�F$X`MZ7[opu�N�үn�N6�ħ���@�Y3]d�/N�I`��F�`Ym`�#X,��2�TT�nՠ1U]B��"�r��Nm�yF�F��ņ6RRˬaF*���ыi9g)�mʆcx^Z�-�C& (f�,$h{�����+^��n !=���22Y�zf�ݽh��߶۽��TB��Kr<QbE�vlX������6)�rS���f�ֽ��7��!8�QR�[�!OJ�ۇ�4b�؅3�\��m|��Qy��e���mIt�̗�G��)x��;#�*ɫդ�t֙yw���"���Ŷ%��QGjĢ�n�U�4&�@�Y	��{�d�{{5��Ó��'Q�J���\���S����حn���-d�R���E�H1IK:3q�U&�q# c{v��7F�[��a�P�ZP�'��:�W/�v"�)�v`1�gV��V�&��5��J�O,�,X��-�5,��
F�f`#�tƲƨۣ�F�+���'XQ��d m��{�
�ҥ�{�$���%�o+H�h���1kSV��ңHN�Y���ǥФ�tD�t�C2�H�=3nY�1��~��Nc��[��-q�h�ʻ,lQ�03Y�(5<Yj��Y�R&�E��m��1+�X�~�"4��/���x���;&E�v@̈޶�7���Y����B��h,�I#B��=)�Ћ���zB�1�ߎ jM�d���"ƍ��h;Z�Ec]6@��S1�7!jT6sCI��r�dҁZ��Q�Tl��f^����-d������5��܄���'�n,)��D�㩹h2)��nlLӕ�&�YyK7hRa̖�轥�5��A_�� ԅ0��w�h�ۨ圬�V�Uu-5r��6��Ɖgu�/hV��4]:dMF�cF�<��neB����x	!,�u�t�l��ˢ�i���5ͬ�
Nbu��L[ǉ��d�P@T�wI��J齢
��V�͐▷�ж���D�p1�@&6-%;5�H�Մ��&��Ԓ�mǅ�V�9�!Vs^��̺QP�XE��2\7�@rEXh¨�TnMَ��eIj���v0�˧���5Vd����r"]ɵe\�����]Zz��vַ�F�9%�6�̻w��ERd�ړV륈V�W@,�WYnΪF9X2^��n�
�-$������j�Cu��zcǮVf��qDS1Yp��-��L�nSR`�qQ"���]�����8�Z6��{�un�s�$�nwo�i��i@��VC
�����3*�-Z�Ք�N��U.��Lԭ"�)[�h@ss�M��m� ��TC�k+`���,����v��%��/�e�$�K0�4�c4*�����YX\Š�_F�h_C�0~k�ЎM��$�	Di��;rv��zV'�po�Z~$�T�^�L�wр��Y\ʥłbO	�k�)��ws��a��N��n�p3��q��"�	�'��4P�D�e�z���fb�WE��r����ɉ�ḥM�e��IВ	{Z�:V�`ܡB��e��jAl|�:�k룺��B��ku͘u�X�L�jY�n���k.�d�������4�bBe��ƌY�*�/�O�Kq���� jbEɪ��ʰȄ���Ī�j��ֽT�ͲR_Xl}
���#�XֲE�3�
��"���	E�$����V���l�tpʺ�a��Ү���\���V�	.ڼ��ue%)َ���L9,-Ԕ�[��X�n��X�	|CUl�
sm3Ik�F��Gp �Q6.�7Q�%<FڳI;Ȇ�l<)���V�4�ބ��ݰ$�n�ّ�3s$/ݔ�UO�P��eB�-H�����m�f�c1j��i%��K�܋oTnI�
���X)�r*�wE�hPYGNL��h����r�.������<98i�ǻP�G!�.���G�RV�V�$J�bą��7X2Ռ�x^�F'X�O��#Qcar�����2ތCK�U���v�+����������h�襢͵�������Vk����Q4(m�n�SQ*�Ct�T�ASج���f�6��aV:�m,={�p��Z¬HF�;F��˫75���N�ϝ�1�l��Z�����ܫbf^K�@0,�ܫN@���"
�j�R����k��b	-"Y�v�.��ʵ�Tn��2Vd,�r���x��k&��46ZԎ,;Z�:h9�wbM�#>O5��z�%��� W�l�uy���Xt��D���٤rQT��IXj�ۡYz���m��W��×��-�}��3n��Ym�(��s)��F��
EȾ<�mD2[,�jZW����@�ł� ����U�KK�9K���F�UV�Ѣ��)"����Һm}�Ä`�v�!W{��Mf +]D�ŗ{W���ne"$u��+Zb��A<E��
v��Z�T�֥����l8���uvӻݤ�n}+r�҂�5���K�캿�ת�����pR�(��F���I��Д�����,:WW2:�^TF��6u���I�voa�T2��i��Ƈg%�-�[J�'D����r�7t�6�
nR��))�ײ�è��-�@Ig-�2���@ۭy��@ƫ`Dk Sb��#j a��ٓN��ybj������j�,���H�X��a5yƶ�b�&�0��-EMbĈ�1e@�XV�����o�����V��إZ��]������7�Bݣ��N}+ �i�;kRY���ťtoT*ѭ�[o^�0f≍�Ĩ$6�hM[IC���똻��D|�Q��DJB��*�p�N�f��-�v������o9�O�-���JB-�w����9B���2�-���nT�s��C#v�&��*Gm�ј�ɰ�#'a���B�R-�c��v�O�6V4�Rb�2�J�X+�Nf5�%�<L�d���Ŷ���fѦ�X��:"�˂���͆H�����Io0�jzA�nD��S*7$U�$�hPx��CM��l�Jm���p�[��q��:�T�P�[�-��Y/vmkx��5�a�m �K�͗V@�eD&o�d�4�(�a�j�8�å�4w�����-[`�)���4K�Y��A%oC̏HA���`����-��1�VU�͓l����֯��;���(���!�\n��Q��d�f=�A�=6(H�hH�W�E��,�l���ω��(���cՍ�p9Y���Zq蕒ݫuSqk׶�q]�(� A�'�_���H����#�e�ldͶIH�un�0�p6�4Rb���(�%�a4Y�0��艕O* �%fc��Z��x��Չ	o�i����b���r)�H)�*��j<i�e�)f�̧�[GFM\��Ȯ!6;�!�f���S%#F�Z���ڼT��aR���*Ω�IzK:ۿ���k2*C6����LRe���[t�c�Lhq1ˎ�5(�.G�xs1J@0�؟�Ș���.�����jAV��W��6,)Ju(�R4�d1��D`c���yW�ެ�L-d
0:�dx�1ۊ�L��:!/)X�F8�9�0�+����3)V`�����=r�},��L����R;�dѰ�D��\餠���YW��mx��U����V��X1�7dy��,�p�g������Kwd��N��Vɗ��8z\��m������Ή�y�&�]!%���W=x̫��C{<��x�n��Q�n���hdL� ��ʗ�Wk�HE��-���]]g������}�(�m�[��ժ�7B�U�_���@@�c�0K�s`�̚l�372�]����=�^��_9��"�Tm�]t�$vubN�gI���1������tM36�P�:7�Q�}m���e�� ��[T6>ݐL��冹�z��ϸnʹ�����?��%<�w�Sxe�p�a�|�ѕ3���^�fO<#��`�?Lr�܎PPqN�髖��$���ݭy��Yȯ(.�۶�G.�㖃�F�!)�0��!�YՔ�ӯ�"e55��\ܭO��2��ޗ¥�G�Ǔ,�2Y��Z;Z�ݐ6hk�G]����uY6C1��[:�^#�$�l�B䦋A�bW/�)�Aww:�9�q���:�Mq�ԬF�/E�A��9+4�� ˙8���x+i6>;�}�zm��@]��Na���qǪ��[���Ac��(��'�6�wd�/||���@4�v�V�����n')�{�$�0���鲎���o��e�`��϶T���&�7#�ou�wX��y��:�tmY���Ǻ(�&���o��{y�u	sT��б @h����ξ��b�تK�.˽1ʪY��-�����W�=��('�����;\�{\"�wF�5-���-=�����X$��a󛻈�������݃B��ozc����Ӊ���+�0��'��V>��I~ޙ4��T��f{�t[;#�\��3U����w�Ģg�\"�5�wJ�*Dౚf��e�����Y��ԫ��++ }��͗NJ�Mo:#n���ڳ�r�;H% ��&	�����tt�Zm%uk: 6���p���c9[�B���f�=���E����=���|�/p��u��vmf�ш8��b��/WK��j��hاZ�{Lԗ��1�(}�y��Ye��'a�uu�^�� ���}3%�*\y8t9-�)�9�G{��A�aZ~��Sf��������e�У��A��2x	. %>D�ͣ��\iJ gmt�XżJ��ږ�e��k:���{��%��x�5�o��Q96a��V4���J�q�b��uDi�$�6���ާ���ʔ�u'�hX�LR��έ9JU�7T��8��������13�.r��7�Io6�Ӯ��O� �X�*�I�����ԯ;T;�s,ʳ�ӝ�`2��G2,O���X'˂*2��U����D�	�Y��\�w�)fWV�n2`l��ǡ��ŗW�P�.����1D��u�Z��V�Yu� �)*d�7�����RK�igP���X�P�(��� ��n���Ƹ5鞁UV�wf9I�p��3�=w�7���6	s�u��@�}�FqgPt��]���*2(�}KՌ6�w��g�TxM�V�$C>�֗��Gk/�V+Օf��:�tD��ڕ9#-	�mi�L�*�Wu�ٚ~�q75۾nr�RLjt�t!���q�Ǵ���5θi��͑+NW0(s�e��棐�fJ㘚�=��:�S5�4�v<8ﳖR���ؐl��I�) CIۣ��%�R �m���֫RC5%��X}էt֒��0�����dj �Lun�bo���5� j�ɰ�9B����$�����g�d[�7��1z�ɸ��Zg>��g&)�5�E���qþ���"���'V�X�C�,�}��K�X������0ˇ!�,qH-�J=���J*dzn����]�p�z���j5o�-���q��4�죘��\���3J��jy�5a�F5�{u���yC{xiM�qc(��8*�ѹ�٢f�x�յ�ٻ �UA}�g@p:�zXHPR��|���N����v�fP��mI]SFo3�N�*��J����%�R-�w��r��ى.Yy07��j��z��h��׬)A玣.6D�T�$�����z�f�[��`sY6��,��ט�����r�>�p��-N	7�^�i`v�=�vl$n"1B��)�M�X���wr���YF�4��ô4��YG�3�#jv(�[0XA��$ha3WK�3�v
�y���]�T�R<K��H�sq��I���|ܗR�Sc#����M4�S��\Z���,�>��讻ճ��v[��_{7��7�˒N���떤�m�=���5�{a1�Ǭ��1<� ��y��E�(m�%p�����Z�DߦBWݕ�}�^�w�[�o���Ё��Q��e�Zxx����U�ҧy�ע�x'��J�]5�[�"t�րzrKK�<��>ܑ�C�gw�)3�m��\���w����Ȫ�{���T���
���6;�t!6ur�/�Ϋe��K��=�~e�Z#9��9.\����N\�Su�cI���ӳ�H��@��46���O���E�kF$��X��\�n8SU���z�RDb�ǵ���0�5`�O�{�	o;�H�\��G"|�Q��3w)�]�E.)����G�E� "�fZ���#8�8h��>�&woY�g W�����@GƤs��i�UX���-�Ż�bBOL�l�*i�\��\����%�9�7K�cS��{N��P��o �ᲆ�p�:�=Gȯ\A� �$��8J�j|�ͻAR�1�R���F�v��&7�<�M��T���=�"�j�sp�:2�9t�Cݛ�:*���B���i�R�CY��U�f{	�W�{�ܳsz�vv��A�^�����b7�DrYsM��i�}�2��V�:�hr�1Ӹ��==ξ[ip�3�ރ��Օ}��C��V�#|��C��L�˽�2�H�*$IA�ˊ��]���g���[ g���VF"ve�X�(ϫ�~�l�E��T>s�����<:�AO���Ӻ�龏H��VK=<���H�E��k���h�ް���6e\b:�� z-��Њ\��!��%�Ġb�ɽH-�]fv����.-kj�rV[�$ϯo���]�KR)}��^}�(�ܛ���s���ue�g2�ې�tg\I�9}�	�T,LYGh�AND��H\r�ݫ�xMނM���y\뫒Y�k��ş�z|��ѝ��t�\��n�v��'���}���6��"�5kЀK�C��"��b7��9@ɕ��b��ff��bS��M�,�8Wq�~��q+\k�L�R�Y�z�fŝ�LC:�$0�+V�pTQ���zu����;y���p6��n	5�)u��(v;�*
��mp�������2�}v3�;��&�˸�'��Ѫ������p��`��F�;��D�w��7�TZ�Z!����[��βe[�I��I��7�2xm��q?+J7��Y/������_W7޷/(���v�)�>�2�<�=��xe����EP��o<3�y>��b
��{��3N��L�K渁:����C +Yz��
o9C8����S(�.�Q��])�2Up}Ѣ��Cj���'vu=8��&ݎm���U�}٫���[��lY����*vS�Ⱦ�#��k��Pu�7�jXJɨ��3j�T����!}����w[������P��W��冭F�iV2���p�#0��� >�F�{�e�6k>[�}�VV��t�3Nv�W94"C
�8i8��J��Fl�h(
31eDF�B�hX*l"�ȳ�s��R'���h�g��>Er�]�c��w$����t%\gTA��@�Κ��'ic�w����-��-u���|���nmR���oǈ���lQt� ;кnt���\�ĲJ�Vm�6�l�o\�5lB��.�4'[?o��\�
�O�(.�fӒ��b�u���ܸ��k+-y��.� V�m��u2���#KoL�±�g-jYI�dr�pbQ�� ���}�M���+;�$�_�3��yb�&\���/,�{{i�]�e_a�����d��Ur�����w��>���x�1��Ky���fvu��,m"h:o�f��b�T�B�lϯ�Yw�Q��F�ڸn��3`�y*���lj��	�a��
�z���td�=nn�{��k }���l���)����Ȕ"z3�
��Է{9,��k�3+E��zs��'mv,�2\m�*���2�n���L��èS�v$�V0]�"�T�1	����kW ����\y�Ϻ�	OzNV��}ܫ\*Th���Vll����` N�|�.KԔ�x���o��֭��w��$��i�ҦeFi���]��[h�Z'[�{�ǳ�>���?W8A6������V�gGj��ys������uͷ<�y[�اM��*�yU���w�Gį{I\�b�$�Ej�`���3�c����!�Ѻc`�FH޲�]ɎR���sm�]����;yk"�K���l)�-��z�6��\6X����4T��֘�I���|�v{2Ļ��������Î�®��+U��E��Z-�@�r�7Z���QGeG����yX뺄i�珒�@�+��!��:.H1��M��s���/u�z�!�V�������K9���$+5�g(�:��	5ʹ_N�����:���]_��*�.v)����|1��U��Ե��*KJ�'>u.�˂u��f�&�*<b���[��(���a�@M����]�FWWT�3�=��ʼ905O\F���$Ieb� Wg/>�ҭ�� �չt��5Xv��1��j��c��@��q����?�Y�ɑ����9\6"ࢩ`љB�������+q��aO�`��}�QVzh�]�Q�5���b@&b��ʲ�ƙt��0���n�itb���Zo޼u ���u�S���v���:���Beq)�/x�$��Y�Z����Ol�Mo*�m_(ī�K	��"wt�����Hx���}�ݞV,׮�+'��'���-�ρ�oժ���Q��pO<za	�ڃԊ�UwF���J2Ι��HRz�3�4���e�,q��ʌ����q����%B_lΡ�6��dM�V;�$�����D»��y�ee��qpo!<���4����yf��Z����ډ���=E���;;��m�Y��&�_!��n�kL���,�S�L�t��7��_��mέ՞2�/u��?9y�8ﵚ�r`L���:��f�W����:�- �p�&З�u��5^/h��H�U�k}}�1�_Xn�>�ͥt��l�:l�A�M�K^w���N�xD��_�U�����8��G��#	��Z�F��˸�Jm@���'�%܀J��ҷ� 9y��{��- ���n�q=	�GOo@/��Ϭ��ƻ�V�a�Yq���G�]75�RD6�WG�x]l�n��ת���y�}/.�>tp�^q�.��&7O�A4���ĝ�R�Q���퍵դ���LZ�������w�-�����+@��5Z�[g�Vnug.V�F+ps��][�s�;[�����%�]��0H'f�0�E���zG*���Յ�C��	ͺ�|���Ѣ[�փO!����V��0m	Ip��\2��n۰j�S��J����S�&�pWm������̶�ѫh�B6�K����O�v9bv_3���z���u�8y�//u�A������Ɠ�WI�f�Y�B<=e��^GwY|,�b�:D��=�Ǫ�_��z�F��/�nj�ʳmI��έje�£�W�0C-R�g*�"&��Q��稛Ãf�D�s&J��Jv��u�+�Jz��y�Ԇ/3�3h��8:������`���[�F��g�F�|��1h�Ǻ����:w%9�芟n���v��H$!]_l�����*[],�{���5�|{j�v�أ]�Q-��]j�	8�ۖ���f$ rB@��inu��]P�%*�Wհ[ch��:��C�����8�qn�m�)Ul3F�8��i�ڋU�(K�
PI���+-Nŕ.m�+om�w���]{@���G��{Y�.��nn��.�/4���xJr[�A�N��4ܲժ5�6ܽ�||��)�q�O%�/[.M�w����lvd5v��hģӴ.�>�%̄�Q1�ѠQ�m3���k0�����3��+19{MqW:�M�Kɣ�R��+�1�d[�WC���ˈ%�n[����}ˠ-'qcFs
8����T+�ek�������/%��O�ʲ��>n��ye�Ǭ_4�|A����bR��O�܇wS�zq(h��{�QSPM�ɷH��#���
��B����U��Y��Hޛ��4c�I�2��է���Z0�6�%�R��8�>r���;}�F�1�nk2�����o9Q�Er�`�8<�@�r�ߓ�/�o�%H�c朘p�8��>z�M(0��u�>+��Б�b\��'��S���n�p�e�ъZ�[��<B��C������� Gע�s����B��ka]��.�ۡ���{�<R�,���Ra^�8�wLCh�RE���B�Z�}W˦S���[]=��$"�a��;$�D�xvT�x*�XwG�q����`B�[3y��H�z(�;)�]��M�4�mg6�;N]L�H'[�wMC�L�d��N.����ŷ0��m�떬�Q��.�M��x=�Z�&Weň��ܘ�Db7�7`�1�6ˏ��=�O{��㊴x�s'�Rݪ6+L�b���)�4��/:����H��ҤE��ޏ�hJ�Z@��.�Td��*��������}L��o7���T�S9S��T�z���Xw��;�3�����_|��}93¯2���9��c1�i8��a�Zq��9Hi�7�ڂ�W#V��(L��ɣ���  ξ��q�:[��|��ă�0L����V��rc5�����(�6����!6��q�b�Nr����z�pY{qF޻x����ĽKs"'�����Ն𛥍Z��?�o����{�e��Oa>87��܊zaNi�of��fo��-��}L����׹���x�Vyw/,�t�_�RH��_P�>�T�72�/"��6���;cp����p��R��ۤ����R��xqQ���O����?s�:[�ćd�4 �n����U��T�Y�W����-HHю]$�/2�uc�I���u\6�'�T�VG3�����5�:�a�Y	����.�9)��U�jU4���o]��p�Yw�� �0`���gMg|`��k�����V�˝2���tu�/$	�\�#=�m�a�	Ж�&����2�/D�P>�v��sE�1c�A�O#�-T�l]��7��֯'�b�b�C�@t�X����M�奬�s6�ښ����X�Dc�"�N��弮�]��D�H8��L�m,b�.N��5Ρ@���(^&�
݂�aE�,�p{C�[WF��4��=L|@v˙��Lv�w(�<8
�t��w�ݚ�f'0�R�B�Fj�6#�����Al�{�nf)n�X�{��ܱ�9�KE���t�C^h�&��@`���=f����ܧk8Wi�,��Z�>���]�e[�(㮺]�؜�$i�^L�IT�ޑs������+9QئӰ6�jz�'���=�s^mX�0�!�J����HV���
�+w�`���1cߵ����aP1e�&
��{Y���`��^�A\��T+�:��ծEκTR��M׽9e-�緵r��;�.j�����-�ϜN��v��`�Z:K�/�LLW8�4W����U�M�<22�'��+!����wn�7���dun[t�oY��/��L�@�7Ҽ�D�/k��C,�,yy���`�T����PoK���Q�e��_j�J����nZO�\ �ݞ��ހ�kk���B��;}zJø�@�h&bv&MaXwjUJ��S/DL���z��Ȑ�0o1)�t��/�sAf�f9��v�.��jYNɄ�r�����4ib�� h7�zV��.�wՁ)a��ϳG�ӏ��g>�KU�P.�9�N:1(�/n�8���;��4X�����_*r�t�R�Q��*�;���i�ػ9ob���f������8AK����6�Ln�=��0VځV�):������5�⾣�Y�o=��8kn��d��ɪ��{���|�}��s��4.P�^�t��ɳ��{�H�ۖ�,�e�#;�ԕ�;i+h����ʹ]rܯi�D�e��h	���#FJ�_U��wv�W%`�����ɝ&4���.���mA�~��Ρ6oj�,���b�Akk0�!#	�o{묔[;��V�qh�S�wy�l�$wv:q��!3Yjn􆅆�l�d����h��:�:��u��o��v��C�����Օ(��0��mR��d�\Mu7PM�ev�hP�t^�ˣPg6h+�Bf��j�* mm��Y�EŅ�Ңj����+�0Β�E�o;�NR���4�_	L��a ,1#�GA\W[��j-���ȴ%D��q��j�۴-�ld�%0i�fU��n^�m�>;��xJ	j����,t%�Ʃu76՚��K����:9�v��v��J�s̝Y�C�Њ�E���H��x�x�7j�;�wM�,M��|��3�ٜ�[�K�����<�Y�J8�,��e` V-�K��}��Yge@��]�#�\xS��>ç�l�+^�']��y�=y!4�,�ڻw��X�.��jSJ�89Zs�Vr]L�\�Ӽ{�zm�:71Th(-�I���x�tt3�_[��X�'.�y������h �[#�]v�� ͺ���^�nF
N���{��.�UpgV %r���Z9&��/7g��"��t�.�s�G@���IiMZ��qZo{g�N�B{t x����/�;�zE9�N���?{8HӢ����8�-I<H��Y��R�jcZ;�U�g5V85���lu���N�n+��j���\�#il�Zr�B�-���fvN����60�2>�[l�_�d�(�4�윖_+L㻓��B;Yb��\���⻳kw�w2��)��O�:�֣@S�Xզ�8�Y����X��ފ�����
TW]��YN�W��\t�p�����jTnpM�۵��}wZ�����)Y�Vn]:���0mԘn�N� ����b�B�i4u��R��:�ܑ��UA0��2t����»zK&�ގT�+���M�y���[�w�����)��o��q����,���Q���U�nj�.a�x毎X�Ń�ʛ/��j���y��kJ���"�8��������
Vj��cx����ʩ�̜�]˭YQD��S�@�y���Z��/Q�-
�p���w$Ҁ�r����)),[���Ѿ���I�>��܃rg�4��K��d��Nn㥄��
	�=�"�u%b�p�m5��	�;�v�����ij�F��V7��t%����m�����-��+].��/��X���(�o\����f��q[�����@�8���fE�h�W.���k�%�W'
j*㷋�ǔӤL��fC����&�8^+h��Wi�Eܵu^Y�q�yl@l�nI�mc�;:�
�>s���w.�u��i�6�����J�Q+}qR�Wl�x�eƯ�pf$���ò���u	��1g����Bcتt�opC�#��Q��+hYG{K
��|N;ʾⰒp�t��{Z����ܹ;/A��bt����qAe�����������櫪��Pa�/M�ZO�-�a����\۹�����(d-�M���hd�5��7��r��/#� m��kA���tyf�_c�3�0�6f�T�&3�ra���U�f�t���Jt����
(�j�R21�.-�|.Y p�t&lzt��ҶA`�5Y�ͧ�.�᛻S]�����yˋػ��[T"�����|��x�1��1��o-��[�r-J�g�v�E=z����@P6�k�m'8N:��/�o��"�}{�����Q�إl`�{P�Kn�@�ՙY˨���b]֟Zc����U�,�6X��5��Α�P�0M��S�`͝�n��l�� ���@�>�v�����<Y�.���S�v���N���8ű���E��_l�S<лA��?v�d��s�W!^6V�ץ��5\O�h���]/_*Z:t�$~�NKf{=�<�VL�>���}�l��*�t�&�
w�\858���USms{��MB{���|����l#
4���*���Rr�^F��6¡��n���`R1�a�K@��.�Y'T�[,�1���<��<�ݲ�� Q
v���dL1���:�72�ή�ۘ�.�Գ8h�i���Z��� I�T�1A�'�nSF�*s]�lLU��iu��=rz��+��Ʊ��mB�a��zo^Ҧ:�[�R���w��,�	�
�Bq���N;|�:,��V�E�ܲ$ya���=ZN�Q���ﻭ^wt�[N���Q�f<}�m]j|���k4�W�O碃5,��*�ۃk�9�Jڷ}��;e[uK����|��A��N�͖��ұ�2�N}`.�_\%��8^"pvA��K��%,�E�ȕ�͖����Ų
"83D�;H�]8
77�o9���
�p�b��{p�3�ē�n�Gg��v�=�{����E`�6.Ȓ��t��\i��A��ٴ�ܶ'L�������}C�y�Z��O�U5#�����>a�.z���]1�sP�"
�#;hf�T	�`Z����,����ۡ��2��G]��gQzΘ��W�Tk�YǛY ���@�}��3^��	��_��+�B//�*���J����1��༸.w)0�J�s��]�J��H$�+p3���wF�hmtՈ�S[C��:[6�^r� ��-_Jg�<˖9b��q�.h�d���h\d=w1����t_-o�M�n��i�e�Nd�q����G0SzX]t�Wrr�;K@�.���f�{V�����o"ﱼ���]C�8�Ir��/�z
G:�Tl�NjЦJ�+�ut����p+�E�tO\'�T�v�LkUac����6"����[!�p�S��&#�I����E����K�������ǻ//��1Ӿݯ��	��q���&Iy5���2�v3�Q� �����CM`���"��)��1�~�Tgm�=�s�w-��n���"4yT��Pa'N.I�z.����^E��Q���z4oN����p$��2(qgJ?]����S�Z�J\��s��T��_7y�Y�.z��"�f����WRV����fT��6:�g!&Ve�5+�Ƨ]�es
�B�ww�^h2�0��o.8j�����~��L'D�v5��U�C{���=i�3���wm��h���5��ڍ�{�K{G��{:��H����c��.�^r͐�U��uP�nu�D8��w�x��P�#�ֹ���򺷦9�ն+�mM�C,���o��+�wʙ�Q��9���Y`�s"�u/��;���zZC��Kv�ӣ���S�I�`�k�-<��Eim{���0r9�V֖b߸�N�Q+�4,�m'sE��GYS�H���cN������B)&���i�	��r��s���\M���tWp�z�Yb6�X��0�bc�oG-c�<Ŝnk�����km��Xy�m��Y5(����0��
}����V�:X;U��àf�(Չ���1����>�j��d�/g]�	׋��� $���
!����)w�c~�C�f���6o[��YՍb�w�&����s�����nk'.KOy��9�N��V�:��Nq'��8��7�;��v���R֤C��.'�n����Z�K�T���˸���pr�`���Fپܸ�c�M��15c��%�#��
���8'V�LZ���A�K��WJΩk�P_uKѝV8"�������n�3,;�y��w��iF�`�U��r��_o����['ސ�,��i��;����a��8��h	(��^7�7�J�����:��biǮ�������
%VH>�B� 5y>����v��
�/�tJ��}�ogH�enK�n ��嶽˂{<h���/UC��{:�([6+|.fԕ�Ft�7D�����)�J)��{�X
������~��]��Tp�G0M㊲�ܩ�(^���Vp�{��p��E@���%���.v��������ۀ���~�j����U <xZj�4��bݧ0=�/5o`�Rn7|GE�X��\�d��dM���}�͌�9��k7���zIǮ	wΑ}Z�1mN�P<��pu�_a�-W>���/�����t���U�X��/����Ǎ8͹ԯJ�u94N��D9V�EC��6�h٫b�K�g��/�h�a��A|2�=���Z�3v���9��g���áۈlG���窘�����oy9
T�~ڻopeI���B)Ov@Rz����e��D�3�Dڅb�d�Y[�[d�!�)\~@�Ӓ���B�_1�WTy��m�p�0��2QF\{�yg��β�U�	Y\���X�C�gRf��q�+.��¡�&��2-BCwK�4{v,͋�)�c��wyx������׽��=\ޢ
	`ҡ�X�*]%�;Oxt#��e����|����J��;r5�{��k��I�c3��3�7{K�مe�\���~�E�m����'Ƽ]��ıQǦ���R��>��8�2F�F�)�"�5v���$ln�/6�͊�1��%�s^���G��B�2����mV��=�R���v��ݟ�'}���m̝a�^�.�9i�V1��� j3�'�*r9"�-��Ժ�Y�9�x��)���keޭ{n���ԝĄ�M�������B�>��4�o�[:�e�"*&�ƹWSv��X���ǲ�ͷ��#��Na�X��I>N�[�7P�^�$]i$>p�
�j��U�,,�(�o��E]�Z�P������9�+g�0w�w.4[Y�qjaе��u���*3�n�;�P�9IY���v5��%��Y2���=.����Ȅ4�Ɲ���+*:�Ò ����n(,4�:jbb<,��p�Qae�z�u���ǥ/�Ն��ZTH>�fC�i��`ޛsKdLw*󍾺���c"��J.���l�P4�iV��n@��3wVq؁��l#,:�O�C�x�cR���[講��/�Ê���v>q�@wuڻ*���eǶh��GJ�ы�D�2AR����^ӷYֺ �w�]�� ?C���. �v��.��jӖ�M�`�Y,�Wn$��g\�j��DR����Vt�m_M�˵p2��Kx����Q�:H�Wҗ9)
�a�.��Ytg4��7s"�a՜#cSp�!���f���'9Wy�"��-�^`�O�#�3����}ȸ�5u:�R��(	0��Wqi����Z��K�n*G��7E� �T8�����'��nA{������:�E,�e��+o*J�I��x^)rK�p�(������{+e�*�Ja���V�
X2�y�n�>�6��]>_���:]�ۅQPv)V��ȧ_u΋@9f2Z�lA|9W�T$`QS�x�mu��x�ߍd���eӥ��kzfR��qr�����1v����k��FI��'����w�R=+#�c&�E  � 󦁸���{���ɝb}�T-��fo3y����ޣ��ܵh��x��!ݐ-մp+op��w�����i�ՁW�p�z��X�뮛Mbge�+]y)�8�^�4�R�VB-�6^�N�	�v���Z���Ʀ7���u���M�{���*��!�``U5hlM��M�]����|V}b�ZW�[�>�Txu
�^T�	4��4T���w7 �틎�O�W��V��nk��]u4
s�����n!1ï�ݻo�U� U}�|�F:J����hi6[���R(���7W´Vw4k' ���XƩ����ϭM��Ѹ� lp�Zgn�N�N�EJ���)eT�LQ�i�F�/�!���@��HOz��������� Uѫ��!���\x���vN��LZ�-e��^�V�����hdy\6�
�!�n��{��d-:����Ö/5�yn�sq��b����8B��S�=� ��+���D�5e*���O�^C�'P�`�;6�h�efk�XF���hc��ۤsA�m仂�[Bo�Kc��-l\���PN�t�H��Wn��Ӵ[��]���[�E�w�������ͨ���h��;Y��d=L�)u��y�0���<�iA#\�%������(�V�p��ʾ���YDy8h�fW	L
�7e+������vK�M-��\�gC���vaw��|�O�I[a�a�]�X�z���W��et:��G��J4hPPUz��t�5��Tn�f���]�[�&��������f&�	�89W��Eஎ�B�7k���玢��ur��V��;�G<AY�*0���C�$C2N�tHL���WL�*r��UΑ;SeiJ���C�azl��;����EF��C� ԩ�9�h��D�5L��ʊ��'uP�rG#<��V���P�+E�]-*J�(�䫜H*���%�n�EJ���p�j�13C"�(����.�^-(�Y��g���%��	:E���/[�e&��j�'J��p�+	3"��Lw;���V\���KI,T���"��3Y��HTI��Y��"��;��":�HQ�J��#Qt�4.k�{"���t��APO;�a�*�ݻ���R�m��}�߿G�׳ڮ��K{�3Mf�j���ov�=�Q�0#ï��n\��Y�VG��x�Y����|jEEt�����wB�:P��[�wv��n2=ZR����u�u�mW,����PƔ<BP�-�Ose���i���� �v�~�E`�t}��c�%AJ���e=OL�[}��c�j
3i@gK�uP	�uX"�+$��%f�sLF��A����TW❮R׀��L��5����e�.3��}��1X�pW�۸�wE� u����1�TH��	Juo1���}BD=�@�e0;��1��m�k(��ݫm�1q=��Lp���3����}bwV-��y�. `�5�@�[(	�D�yl@����W�*����2�^�L.By"��.$�S?Pȳ���:��oݮ�6�c���[��y$�F�!{@U���*,��^�ĬY�)�u}'���r\	�Vs�����v�l]mսE�bG'��w�NX�{�x���B�&�n*���ld�?U�|�NT,wA�gA:��qqː�1�N��2��*L`|^����q�^��)j��\9�ި��áy��.F_l�¡3�#kw���3w�8";�_d�C��R0�}Pt�z�LZ����lOٚ&�>w�����'��+�I=���ӪS�60^�V۵��޷��wpC �xnY��!���0:�H�.���c}ӗHӢ[��J��u��7g$����%�}fwN�pk���긎����i������Tu²��2��4�鳃)��"�^��/��N&cVZs���O��h�|ڿ���9ŀ2b���f�����3|+)�v�B�\\�7/��D��eB�Yq�EJ�i��p��U�ªx:�]�+�����q�C1_�Y5]4*
�x@H�A��˺�J�l�<�br�m���߽|�m��u�*"�tD"T��yPe�0X���S�s>3�@Vh�����)��`��8յ��\�dM������ߦ��rC�1�~CI�G
�/�ON>��W�_���扇�\�������jЮ��jY+N}u1�L�+�i��)f]fv�uU��a�ä�LX���Y(\B2\�6�I�z��y*�Q���]±qm�I�ŉ+�Ӯ%Wʾ��1�0��:�� ��,1q3���,2v���6跨@��Y�ov3��r�����8#�O��9:�2���f�����)��
�|�Vo�xi��>j�Kդv�ł��=f7U�l��hOx�9x�rtG�R��̓أD#n��nn��i�뻼����'p!G kF��7rN��9�n�<�Wۮ�n�O���WZĪ�z^�h�G�����O�:�Ką�c}��	�o��8+A�&��.	ͮ�X�\6��H�ܑ�Ɛ�����p��)���ڱK���B0P�~f��*�(ŝicڑg��b�xoLp6`mOC;�
E�5�薴�@M`*i��W��{fJs��`{�df/�0����'{B �'�����c��Oݗ�0n�g�����W���<n��4h�@j�u��[�KNN�](h�W�=Ş���6i��}�Kӌ���=�'�Y���L!���j�vW>�v�n�Y�qU`Q\@ϭL0�쪎w��\PΙc8+w��Ҧ����UfM
�ܻ�b�}�,l�=t��1���*Ƴ�|��Cq�CA�p�����8fԍ�q��n%���U�1qd�WH���0G��G���yG��(ɟql��r^���[�qf�	H��8��\����!_�e�a��r|� ������=�VS����=���G5LM�*�tn�t0�R@�v��0�T�����^<zBM�ܶ�oM�H�ʕ�.p��W��:�n`�K1�n�Z�r@�+�v���f;t��B��W�*M؃e�ï����B�8jo�K��Y�fh���kpn0�z�*.���9­R�Ef(]b�z7��g)��$�p�޸��Mg���-��G"���J�e�9-&��S�_{�n�`�ӻ]���go���I��] e��ުb�>\�ߜ��b8?���M��C�b�'�wq+w�.ǳvp�k�������5�s[L`��4��:L1_6��f�F̶ �Z�fGM7T�5]T:˂l@��������'C��I��)N�8Ʉ�Wt��ލ]r�L�o���d��p���&�Q�P�&ˉ����_~Py�V�J����2�;S��x���u�\��bvV\,Nk�!�:he��׽lٟ{�&�W��t��i�ޕmst �gx�/<J�ũ�u��v��v���F�,Y͌����K�f��K3]$��W�M/oJ`����#&c�F9���u� W�=1��t?x��AZ�=!�y�TfwX�4�R5k����σ��񖗅p�(U�.�����wL?��ܦ�Ue���\���Q��-+���R0o)I�Eg�t$Ns)�=�F:����.o��v�,��x/�g ���1���Ц���S�Dm�{���k>g�O�Rg�˅�R�A�����y[(]���Sc:��'M0:ȇ�.�EwH����z�t>�F���= �d�s	�U�I�C�r2̷ohw��2��:�j~LH��D����z��#u��>:rSK�ys��`Se푑ҳ�5c'^(!z�r+]y�����:��9C.E��ݎ�=:��p�Sg#K�q�҄K�v�t�VF���d��B��Z��܂�b�Ios.^�^�sk�-�mWw�p�U*L柰M9B�7NJ1)0P��3�#�3�.Q����3�G��Pza��wֺ�5g����NF� �.J�O�Z.����|Χ�վ�^pu��
��6[n�B�:
F������1p�hE|�7X[���4Ed&���� ?�xDL!t�L��ձ11����c3`L!��1q	�[=�v�S9�I�X��]��N w+�2'OD(O����\�G:�x���pT� �4)�$��9���!]��͵ 6n%�`�d��d��,F�A����Vq�I����E��\���'�����6(̽,uG��g��`3TT�nf|�F��ԕ�(��E�#~�6�.^,�U�v%{(P��r���@f���%NTB�9Gg8�̈́�Θ���Ӛb�P�7���uvo:�ч�8;=����p���u����D���������!�5��p��+���.˹�/c�Egc��ڄ�ر�X/!�*�C_��giQ��䳪��hˣwC,a�[B�ĳZԝ���[�~/��W�J9gv�'3�i�[Ֆ�Ԧ���o��-{����xT��hW:;p��JvG�ɗ��������*"<�uΪ`Ch?��ągU}bb�U���7PU�T�"���&��1��3,��N�'Ŗ��w����½Y��h�оUӃ�IX��|Ώ:���_��}Cx�P�%�O�c^�<]����W���;s�_n��(h���Q�غ��_A48���z��d�?(p��`ou�X�]QR��=�x+6PzXL�/rcC�i���-Dl�(��S(��6V8����U;} ����/&Xw���#��pdwM�/�«w���m�(�dVi,@X��e��nV�v���T����MY�V��֊ͼ�#�ӹ�۷p�꓆xP<����Ը֬�~z~�k�zɒ"κ�p����uD,��"�:�8��	c�h�Վdhːq�"��C�ճ"�S7#L�b�T図6�s� �����ד�5����1q36s�9�`�^�ue�V�h)��0ˢ䋎��P`����ʝÙ
gt����o�R�4������euo����T1p\�.NJ������4�_v����Ny������%�
�q�%^�OC�ݚ\�K<�*�����]{�����T�S���*T�ʖCow��{�(_h��)��`�ǙZ/�3^�)ΊL�urY�x��l��Й�f^��v����u�7�� �c�`5n1��oXڴç�'\�ZcSe�EE�3O�=���8eGP�u���\7?>7:� <��d�jLp��^ՙ�]ѕ�ݩ���T`u��&�1������A\�}"L(jc�RA;�`���m��(�\���ӵ�T\�W�Mk�L �u0�$�8��[/ ��A�F�N����K�����?�gpȗ���]�/�5�g�qb�|#�㒸�`˭ݺy��]�k��F��l�v�ܴ1DY@�δik5,�4�R�˭*���X��n�4jW 3`&���h(��ߝ�t��t�w-�U���D��'<7l�ឞ�<]ہb����;?<���oi3�v��M��z-���Ѷ���Îjo݃�jǲ@y1�EE��ɗ�����2���5O��<v8�
�M��b0=�����I��{�WݜJ��
xq%�Jk4�V�W�w�W�2��q/L\7.��o54�m���^x{y��'kE
���A���~P/�J����[_pV���Ћ�A�f+����<D!cWN��H��.���3t��ɽ�؏7 ��TDc�rO=mfq��{L#x�(��ӑ�@�T���I޻�E�3��y\��­6�W��y���x�Z�@�X���9�,|����p��{1!��8�D���
7W|�}��a�s���E3����+���n��}�n��$��E�\�+>$��������<���]�u����6�Y�O���j�����24j�N
���ȸN�W�@Hك���Ā���%F�խn�˥�#��ϥ#Qm+�'Cg���4GnFq�ȫUJH	��:�&��� k\�o�on<�%ũ�.J��f�<���[��S7�t�w�M9 m+Z��y[�r�/SS��;�w����V�] ���3.�.�1��ճ�Z��s�1`>"�H�����֫�~�]_U]��%�f�j�ms4���X��<+��?v�Wf���z��+8-F���ꡲlh�
C~��W�ɽ�)�0S�K+����T�+Y˜�W�%ީ��܁Ӷ�T�/f��]������0�\L�,�׫��[G�V]��sy�����M�;���2�|N��n;���l.
W^�d�+��H���.�oI�.��/P*e��Jg]���g�S��=�5���N����@2B���_;��0�X��C��Z��w��������PM,:y�t+܏*m���/�l�7,O}��7=�bKF[����i�[�1c|/���obǗ}�#អOZ/���|�>���'�6���n4��P�Z����*٨�'g��L���ԇ��]6�p�S�GW�=�����t��y��oeR�p7OaF�C�i"�����]g��_i1
��Tcn#S���тu�ƪ�ޘVh,o-�)�׫�O��T�zV���Sq5��u
����1��Ӽ���p-�ݗ�]6
ø�#��1����B�N�Ȅ�w�x�(	��DLQ|�:Z������y9��`�|�m���0�t��?!�o�東]2K�2u�yw`�9;d$�{�=�Lw���.;e�g����v��p���~��ܱ�˒��ĤK��n6'��5Z�K��v��3t@�z��\�y,uE���ACY��O*#\�/��[ٓ��e�d7o7���L+R,���
�14t<6J�`��;��X؉SB+���<�#]���f��X=��"�MI�{G��H�炤�^3+xfQ�y�Se�)�pCSb_oJI�� 77K��#C ����-S�n����<�X{���;L�KjR��G����1xr���2�����C(�V��*t���NV��	%ʦ�-h;׌�t�P��	�{KԔ�a�d�sbL���=�OgVu�ľ�A7�#�k�I�xm����
*8ї|�b'��(�x����˃���;�B���<����+��o,��T9]�D��D[��+5 4n]SaX$O�K%nE�1/�A����p���-���x��%���-��&E�{�fkO_r�Ϯ5Lb�ꊝ6�T;�Y�+�Y����E=WˬO>ǵ�)�;Y�"23�9(�w6��"��)��{4%�G�0��%]�kT��xYqa�ʄ*,�(X����y��ک��o�xP���F�j'1m��I��K���H{�+�-t��o���_T6+�O<��;>�xGk�M�XA\%K������8|m)^��.������gӒ����h<˗渟�CW����0oh���@�rv_6��$؅����+p�禾�(h�}��v-`0�%��.�zW{���O=��X��q������N���E��NS)�Z���W+9����P{� �5 ��"��7��Z�C�||*Z\�V��<�
[80<��(<=���zlG�
������ʽwxyr�B��.
��UHꙆ8��<�܍�"U��C�U���w>,����fVC��T�����֍��,sO�:;D�ԏ vg��Ba��2�ns��/����q6,�F���V�]�}1壪h��t��l�c��bԠ�i� R�aҡ˺�C���&��t��7
��Eeo-5؊9�`�f�K����7o@Ý!�-|a,n��u%x��с�O ̖��fYP�9Lb�͢�໬���y�����Vs:�Ok
��S�A�tkj}��>�t����53+�r.;	*�L��垣F�n��u�n �䅂�hA��N�	I�:��@�V3p�Z���Y����$wb�� \/n�}+%�+��Xcj�c�FWq�-�1pE"��7�]��6����.����L9��\�<;1�������z5B��E�(������]Y�U�+�m�u��g9m��*�pU�1 )�V����QkO.�t�{���O�6�-y�]=r�t-Zpb��K�9�-�e��hΠ���fl8M`G���P�Yj��f��v�%N��E�b�ͳ�5���YmA�4V\��R��6��.��C{�j��j��u�5�ޅF�E�#��YՖ���̓�����k^��SWeP�n���*m��6Î�3�Q�啭>�\l���Ot�>�7b;�M�R^�֚���	�F�m;g��8�. �Sv٧��ܚ�RҴ܌M�F;Ӻ�(*i�Qtz�:�rn*��kkvWv7
�1�|�]4ЈA�d}�n�c������h�I�X���AQ9Z��n;صv5��֐���2��0�H�e�!��X48��˄�n��z���W:h�vս�7h�܀ao
��"�菮���ʩ�v^x}�n��(��}�vS	����p:Ws�������\3l�rg���T��O=Q&��ѺmeZ��|�V�!�oV�>�Z%RVo��k� n����8����L����R9�"�{�;r�+zn�8����ҫ��P�7=�00��K��^�xeDQmخXS�.m-���n�k���x�L�& ��]��r���3�.0���˪즻4�]H�%��^�x��)�o9�
1th�K���c巄S�#k$��MݛVK�.�"�f���N|���n�h�;�+{�����-Bel��u)Si�Z�`���\��4��2.���W��Fw��瑇�@�)��{��5�t,@�;
�,�����w�Ώ����Y +)�9�β&�(�.�{}��{��O�j�9Y�}J�C2�Y}7��ϡkl^�;���[h� ����)F+g7b��q�љy/7�:���M��nsx��W�Hs,�)��-\�]��yiݍ����!WK�Z)�L2���[��*��x���s.�z���6�s-k��:��H�:D�a�n��{���_���`�ʵ����:�f����������,»%�'��N�$!%L|�o�w
�#׎>Q���ke��*�9�Z�q��BjN ��=���oI�h�}�%zaf���y����9�#3�;/]�� ���U"1UI)3�V"H��$�z�i�.w(u��U�4剳L�7<����
Ȣ+�!�z;�XsH��=ܻ�D�T��\�,�*�Ÿ�j"J$ET<�*Ke֡aY�-�۔`UF��,T2#+��yWu�͈�Y$U^��k0D2=H=wKD#�e�D"y-�j��Tik-hb(�C�DUA"�4T���ő4!'2�(�L�Yt�9Y&(�#��s�J�\D"��:U	U�wq�M5GG"�,��t��냺w	IL�2�S25P�SwsԄ��M�ʣ�,�����D��
S��(�D�
#6'T�ww+��'��9�f&"���W�"���A�E:���%��&Q8E��r�+�at��\]���3;"��0ts�3hR�v���u#�]ҴI�T��Eps6{�T�.��$�\pG{�翯�/��/u+'Ъ�@79ýib�L9����\��V�ڌ�޻���*.�ħA��[*��;�z���Ǆ%��;�w ��G��}"+�����G�<���D�_���q�s���S�z<ǔ	&�G�!�>!�C�F�C�?!�������J�|DDP�!;����1}􈅔z.�_��0Cq�{|�lB"0DH� Gވ*t����^O�|~pyw�i�~����}&}O����ʁ�\�����!��<>\���\~w������܇���xL*����s��Z};�U����l"p���N�I���< ���7;~;�zO)��������ޓ!:v����� yM�N����!;�ｼ�!�9��#��˷&����|q+�q��}C����C���i��<�'Ne�\Ʌ&�3�14;4���oi�9���`�奔�w�����aW��97�'�|��ϸ��y|8��ｷ�yv�;���޼�i	�����ܚ���r�_��۾G��o(CD�RiLt�W5�u�ž��Cs�����S�����|����q���[rSO�>u�traw��}����N�__�x�~~;��m�����������xw�r�X�#�6Z����?c|��DE ">8��~<G�<���׻yW{M '���i�Oܟ�P����Cۉ7�'�����!�5�|��yq?�I�޿}�$��Sy?~��<��E�������'dn�~�l��G��<��֐��|w��?x�����r������0�o���=��90�_��.��m�y���xM����C��e7�'�����	7�$�}�����?U!TF_ʷ(!��q�2���������ߟؐ��'?�߷Ϟ|��I�!~��i����ߝ�<tɹ���?8��oi�x���aw���}�~��®�z��xM�	7���q�C�1Uu�
��>�����]���� ?4
�V��׷oK���f^���?���������v��Y?�����7 {I<���ϝ�w��������Wo=�����s���xC�i���x��)���D���X�����H��g&3��]'��r�-�P�>a�{�A��������$����iޝ�Oh~w�߻�aT>8���<�_(~���%w�i����xC�O�{v�������O;ŷ&����co�}�����%/ձ궍�Z〙c�q���,��,�a��.&utby�_�L۹:��Z�w��8�Ozb�V}Q�h��F�u	��$����{y�B��:�i{�*�� shE�M>)V�zO���x�G9'-�R��[���7;���g;3�i������U��|� ??�	���������r�������q������=���y�����?''�������w�>;��~�����������������r�q$�G� }�|�� 4z��y�3~���}��4�O����l|M����M��߫�P�w�=��xq�'�}��o����{����n�����۷�����v��u�#n�e�0���n����?�����?�v�xM�	4e���9��y<��ԝ�x����7&����h���C�g��6",G���d��bn@�������w��(xO���g�1�<��Tm��L����������1A��٩���F}�A�����}��O	�>]ɼ�&7��<��_�'x���(Hy=F�;��7�����_}q��<����1ƖշL(�3��-tm�������i��|��O}M?������=&���My��דS~Bw��=x��}����wpN�}~�$���I��y�&�G������}A��\|IG���Ć����Y;��3�n�ސ�w'���P����!�>�������q ���7z� ���Г��=���oN���@�|O���É���`���)��>�?���}LP1��W�0d��w�ߦv��g��8?��B�m����{�����y=}��}OI����M����߻��I�!'�߸��9��޻P9'o�_|��]��H^���m;�S_/��װ�N���r�o��|��D�� @����M�<���.�Y�ݧ��P����U����ǃ������;�o�/�o?��a~�}�;w�ߟ����7 (���?~��zL/ z�������Y��~̵v5p;�"0E�D�����r;���S�i���7!ɇ�羡�Ǖw�Ӽ���<!�4�'�{Տ	��!�'�>co�O���?;y�~ps�����������7���znG�[^����ʇ� ���"�����_���|c�rzq����x�P������{O)��P�w�ߞ��C�
y�c�!���}�����y��(�M���<���7�'{��wX����y��K,�+��m�(�#h�R�3��ۚ��}�,���|y�Mhr|ɋ3x��{���6�����	�:H�h0���sv���/{�:�S
p[�QL��\��;,�ֲ����%;n�fv흪�9��
���F���@" ��uLE������}�������m�N��}�C�[|w+�'~����o��ׇۂC�����<&}~{���M��4?�z=��c�v�;5��;uB��,������iH�G�����s4}"!�q�9��o�ܚO��8]�:W&����ɽ!�0����ߌI�i�ߑIo��.?��7�$���������0}a���>�"!��ܙ��WdQ��e[x9���ޞ/�e����A��.�@r��=q���I���������@��~��Ǉs����^�x�xL*�����򜇴9����c��C�k�`?$����?O�}}����b�*^�m<��/{�������i�p)��ϫþ�^on}�����C�����]������yT¨>��q�>���'���!�9Ǔ�c��X�������B�
�T�}Bh��}�{J��9x�3s\-v�f�b���^�m��H.��},(RM�<oQ�<�ݹ7�'�=��ǅ N�{��<8�O��=o�8=!�4��>>�����v�t�>w�}��y�m��W{���7���T1�yꜜ�6��@k�CD�>{�)�>'&��}�4�o�`��9]�$���x�����w�����>��>�Ï��M�=��;~t����/��!Ʌ�����o_m�۝ݽ��|�Q[��#�?��� }|G�o��<&����ߏ;ʸ�П!���I��pH|���ygo?c÷:w�k�o����yL*�D����yL/�=t�|O�r�������{�_������y>�ৠR�(F�#�O��q��O�{C�z��px~!��+�!�~�ǔ�!��}}������o�H{�|{�yW������yt�y��z��N�|�	�����$�<��yQ@ G�F �5��}���u{}��B�����~{˂C�S����o�����'�������� z;ߏ��:C�?��x1�H.�����v��$�����s�ۓ~OG��çi_�燛��_��H�$]���X��L�;��׿?=�7�<&��O�#�y��]&�z�&�B�c�W��ɾ�|��}�����!��O�x��M�>�&��)��~��������q��������}�����C�A�U�Q�ߺ��4��og"֢�Bz@;�����G��	j�q�R߱vײe����Ӛ��R� �nڼË*f5�ٰZN�7��������v��p�;[�n1E7o^��Z'C�M�V���z�L�˳��k��7 �����,܈�ᗓ���{���׿���.��������w���A��7�9�G?��|��n}�m�<"�����{��7�$��翿|oJ�Ss�}�����s��'��������C��}>#������e]M�6�5�w�+�3�6�o3����Ύu7����y��)�C�}C�|:�raw�}O;�yO�r�_���q'�=������C�W{OE }I�>}�?���+�¨���¾p��PZ��[M�sfy��DH��8#�BS���G���{L.�i<���S
��w�ǆq�>'���<[�8$>���-}_��S��U\>��EAJ��� L1�>�0k��J��i�εc8?�5x�@��< �e�j�H�FC�����
�䑆pGh�H�Vqs�su]����	�10�����j@|TK���L�,��sLF��Pc(�/�a��Hi���7۷����}���z�_���|=����`3
�8�TK�(�h��`�����ÜN�6�d�a����c0���#`�� &"7��1�W\E�vn�X�����v��q*� �cJ�FF %i"8^}9P�YzP��	�X�n�J��7�<(J`�f_T����S]h�A>�����ͽ�Oi!�K����L^L*�[f� b��A���j��%=/PTK���}��E5u�C��B̢��b�����U}�Y�e��5�y'i�Q.��!�:[�n�.�әAP��;G�z�z��J�<�Y0�����w&
IS�����/��.뢮 h�w�۴��"&�Ň�^��v��R�w����A���!��Է�q�r�SUɚ;��}��]�l9h����˂��p�ƸCkv�}���k�x�tl��X'�D�sKj�}�.��N�ga�c��}������ϗP(���H<*jS��2��y�������<~��1ܦ�'UX@"��r�H�<��H��S�"�h��庮��m��u��x_��*k���]�¥���n�|F�@h)�8��_*N�UC�{H��J�Gv2��{ܖ���9Ƹ�fU@nO�CΩ*ᤸwǳ
ߺy�vg����Y|��>׉��--/��&�H [���d9�o���F�'�,��']r9�w��\p�o�"v���%�;�V�V윛����#�0w�Q�ܳP��}�r�������̪��^����gQ�X���=Zj2�s������ E:� �Ą�P�0X�<>or��x���?yF��Nf��}c����G&k�o�����\��@�o,
�u�9�t����?z�A3���[,?�����!��;�������Wʙ���~l�J���]41-;g]w�ǳ}�N"o�F�_�u�>��X�Qxb0�3
���A\�}"LH���ݗ�E71�9���� ng��D��jk+ *���<��q�G3	�<�)���}�N�8�t-�Fӌ`��=�{E7�^�uX�]ɲ��5���k��<-%�כze�;���6o._A�{���s[;�*�;�����vv);��:���� ��m�T�iȱ��Q]��V��^y`)Ү M����/(V��=�Z;V��ΐ�i��/�a�꽡2%�9)c��>�k��VYL������/*;B��Y W��Br�:j�2*�0T5�t��Pu��jYާ��/�{��?Nn��t�o
����
�ׯ/�	��C`�j6lr�`�F�y�ka�V=:%��=y3�cY������{I����n�}���Բ~N����׫Vn�Ե#0�4���	��a*.g�_�%+�f�g����c��(��9tD�壒�xU/�F����S��M��P�*��7�/�� :�Uå�G;��.(gL���E�[�$��[Yi���t]#�҆ګ�`6��t�*�߳�ݷ{D?	ʞ�-R�B$���$��录w�c��	���-����i��c Ԟ, N��F*O�`�x�Q|�:q=K�{U�R[�Q���+v~p��q�n@�F�N
�j�[uPB���	���wTQ|���(�P��,��6H��h`*�Á��9U:�b;q���B�f;Ø'-���%�0����$6`>�s/�DJ��
��D4�p�� }�C^��]hpȧU�e3RBK��� �w��<"^��fS���љ�9���'�}�W��N��ql�a��F���%�Qi+���t6CSQ��N���ۻr@��k��^��\�8P���+Z܊����ܹd�t�=f6+3��ȇT��d���˘�V0"ͦ�~��e
S~�;;�Xw�,���]Q#c3b4�pbD!<�[!3;Q��5g9�]�$b��,_D��zM�Nڷ]��a��,E�Y�^X� \�]&���i�u���x=�02-����Г�* �c��zq���I�3֮�۽s;��|�F�0���w�2YaC~o.���pʯQ��^fU#\ �z�O�{cݏ�F#9�:ߪv����f���=��\���1�:j[�������L`G��^H�����'=�n߫;]�2�Ύ1Xo�syҀ����)���4����`i����Sj�+�j�'Lb ,.J�s\��aB�2f�� b]R�.� 
x���L/��w�.s���ܭH�	���ؖ�F.`)�6�a3Z�L㖗�t������eE԰�k]\6ɵK�_;�|���s��Ǽ�/33�
�߂:,[�R�@/�m:����\�-]��e�'���bX���zp�E��7=/�\G�u��]p⤝���ݙ�e0�����d���&N{�.}"����A���N�h�@_^�B�Q�q۰6���=�Fok�F�)?�g�u�#x�~Y���U�+�w�co�x��������9�c��tƋ�Wօb�5�V��q!�*�W/�*�o�v�l��n�#�|q=�\�p}�0���P�[͵�Y�9|�]�]K��F�72O+������Cע����Վڴ`}�N�1�:[7~�4�������:z��k��rPq����
���P���{0��c�-u�h��������h.�����A�K^�f%���q�b"i�&9�-�����GC�A+�e�����}E�ȕm	������Jw�N�c��z��U��"��1�rKU�w�X���נ�LW��|���@�٬��xv/��D<X+��}V�n@��� 5׽p��ބPe�W�.Z#���=��u��ޞ=�0{�'�h0V	��0�9'��*��d���IL�ӊ꘍'n0�D^n���L%}kP�.�΢���ZL�҃��fgڌc����^�u�Cў45�=�M��PUjP�J�dÏ&��,_�C�X���Rq�p2�/�V�s �'@������#U5�V����\���+����\',YB�d��i^������B�s�Mc�>�'��R��ǭLӲ���'�CM��h=�)}�,ܽx����+�)����D���r��p� b>�O#�lX�1N�x�̜�����n�c��LC�'�F1�7:���M���.6��̂�y�F
���^�c��]�e���� �S�{�G���8l�Ӂ�:]\x���?e�y��g��d��[@������k���}E��hq�0�6y(
�.����:�v���{�h�Ͱ�Uә㖕�8�:<���ὐ�>os/)6I1�tv�`�����".���rL1ې���Q�P�C�]6�V�rë�g{����:ٔ;^H��6�ɔ~���3s��,%��\貑֦8Gq����.�uձ���H����+��q9 F����*._#	A��;�-�a�3<.L�>S޻���SʗOj�V�<�����%\4��;�ٺ�WO,%o����.�!��y�:��q��ԥm��F�q#�ya�k��D\��u�#�R�J��no �/��Bj_��.�;Z$=���>���"��*�2+�雄���𭫪�� �5C��z�Q�����e٥*c3�h�$1Y`���C�K�7��ѣɘ���Wa&Eⷷ<��?�������\�#�e#c�X����|4���ւ�75�r����S�֡tVA������V��"��WWCز����tr�߁����e��T���G���7�����9��O�&4�$�l����n��H�e�rE���=}��+�+���׹ƹ��ս����wND��ܙ���c��E�*�����SqDD���;�ނ����t9����]m�抈|��uV9��D¨�V�&3�~zj%J��庅\!�G�R���`$���^����fc�պ���18X!Y���<'|���V���r�Eə�0Z���Qg�χ� ���3�G��X����O�W��F��f�a #QP�2�zӗ��PGmT�.
��Ø�D��
��	:I���=�@�/M�h�V���M������,���==< � o9�4��\,<(_�����l�O����p�۶��1�3�Sͣ�|A�*����=V̞�1�~�z}�׏MT���l���w��x�t�f&���v/�`6��#S:�/T�`wL1���d�/N@���Cx��5\ ���t]�r�� ����V+�b����U����6O�������T�ꈄ&s*���񍼺��B��Kbjz����AW_[��3��*� �oxS*�l��s�Ծ�|�f��O�hϧq�c�7�W������7�HV��kx�N��8@׭�cVoEܭ|���}vj^����΄�p	�cǹS�o��Q*�ۘ�o�w��qS����FG^]85j���8.xl:���[.=:�<��D����b�rs܎�fX!��X�k���xeZ���(Z���Er�lh�ۭ�b��V';밠ޚ[����T�x���_T �7fp\8((4.)C���tᬎ�1[���Vc-e��<W)a�����PE�n�`��F�]WVn]g^#��!�kg���cǎ L���e���}lM����oN:2kTl���'�)[��:��w7��#9�4�u(�8_t����z��Em�Z�_�M���@+i�E^|���*ܼ�S���;Q������.�N��l���Ҿ"su�0���*\���������@$��v�H�n��?u���U,)�Pл֎n}+�pV6�_n����'�XN����U�Fy�jM�#��=ZP+	�+ik��X��WK";�t%]���-�)��oqf;�R̕`�rvM���]��i�u�X��A�tTK��v�y�����D������)�
���,CW��n����]5�-[Թ���^��z
Ru�j��g<�Ӹ#;\�n:�V��h�0��h��i#�w��j�W�G��Wv+��)m?
���vw�]�X��o��;1�y%b�����gg�*5@Q��i�I��j1Xj�azH����`T.%P��0�Y����� 2ɰv�#i�R�t��nQ�c���@��Q�㔖��2QU�c�U�Ι��b��h=�ĹL63�JNm��Gz,�"������)���A�9Z��n��v�aьuL
;�<�ʍkii��| � ����K��_fR�XA��O�3��d�gӫ嗠)�3�#��)B�Pg��!Bp�q
�I����W�$W])�:�oC���Ƙ�ީ]��}ո���=wZ����Su��x�GTS�`C����6��O
"�ڽر��*����Of�Q�V�x�r�Y���?h�ؓ��ߜ��8��0]��)��q��15=u'��c�K�ΫL��ǃ����"p|/�f��T��kB+ǋ����ݛ
܆��O��եV*�����w(ݳؙtRB�55�r.�%��t�
�������{�ܬb  m��9Ce��9q���%���L�����8=��d_rHA�uݬWS�4A�yd�rT@u��q�}k�*_�)�t6��IW�˓�&l�����R92`��B�_^n9x�a���Te�2s)\O6�x:��p tRV��3�+�&�:�����e�Ń�t$巃�'�I`r����Mt>�Y2�޾o}:f�P��)H�0�:�{yb�v�������ϒ�F�f�W�W^ �+s�����@��h���'Vb��E����&�X�UUe��L���LB9��s��U+�q�I���wOsv;�Kr���t�u�Cm�/T�̏n��A)X���q܃��{�����x���F5�.N&�Ỏ��[�[��Q���]��fԱhQ�{<�1Z:�/J/)�g#P�22�����r%����m���(�a]�u���,N{���JhJB�;�$uf����* #��9�'s(���)ML�R�D�˚��-(�Vi���s)ww,��F�S(���R,T�g$:�뻻\��t�HNU�9✊�jЊ¨J�3+eIft�3:N��qe�V�Eek�S�^�:�DE�M,��(�6r�"D��"���-��"�"TV���;�A�=���Y����sN�J�I,E�j�����'-U �B�OP�E�E��P���<ܤ�Е���p"ʌ�j�]�wu�[,�
���5IKHm:�y�7re�^ >ͩ��5"�׻fy���y�*n*)��Csfe��U�3Eu�}X�;�R��K��s�������ynN�܆;?ς|��վ�x�=����ON�� �{G�]���*z�tqj��V�����+�6m������oݤ��U`���������ʟ��_Y�y[�A�ډ`%oZmdԒ�F���vm��]B�X��v�����"�)�p4��ϯ[��B�������2��ڵ��چ�D9S���rDs7��>��n��VPƵ]���v��ͩ��mڎ��lG�1"`��b�5�)�����L�l���h��r0��Y`-�U�9V�6,�\�dݒ�q0�_�/���0����1qa��d;s��NJǚV/��Z��Z��f��Z�uFv�}X[�<W"��ߔ[��M>�Hf)zw 3�H�%R}�+�zF3-�w%9i.��<�>��1`:���������V-�f��>�>ǃP�a�9�j*;xm����\�sɶ"�j@n�wch� ��� �^����f�B��ҙ�D�)���2-Y��A]t��f[�T�,��a�wɲ�-L�,4Ƈq�/�H7�Hʲ��l�VKr9@����{�gZ���7]������ηw�0�4��W�U.*u�,���A�}�K�nӭ�]{�副"K��@�a�gT<d��9�12�����	��q���f�^��܍�c���W},�ʴ7��H���N��}'�����X�}}X:��z����j���וC�g�۫���~ƞ��52V�����]��TI�������[z
��3�^�evʉ�r�N�������3Г���*��b�����WY#�K2�u��]$<��-��ս�+OVF� z����g���TQ���n����U�,k<!7�-/
��j�Ch���$�٪I 2�'����s1Ez?���ǽћ���);�_T��u�7qs?r�G�w-��;dy�S�F�?tj����#�;�4ZW�('�B7�����!u�N�-����^�@���Q֧�\z5>�h9l�?!�o�r�T|東�9E���93��W,�Z=�����1�?
���5>�<5�)�k�xٍ�b�gG��g�� tl�^GBY˸�:_�4�cL�A��2���Y;�n�*�xk�vϋ��<t �Դ����\����f�adb�s�*�E"���f%�f,�H��:;ML�xyUU�x`CW(��5��#�S�k��|R�V�3O�|���Dv�{:R<-�\��q�}<��P����T�S�� �Y�z��p�mY�n�s}2Z�0��/@_]�ξ�B��#5^��ݒ.���h⬻��r��g6u�9&�b�������/7:�u�֌�<=�V"�>�������
�gP�Y$as�R}��Q�c�_[����vc�%�L`���1p�U��[�#�
 �o,
���
���'UQ9;Z���a��
hb��xB��To�+/*��u$/��`v����� 'ݫ����)[�����|���"F�w����35������L�%�\G�b����m�CV�G!q����S;�[ܯ`,4XB Vj��tmp������Ea�w���o��~5�u��j�^�JXWn��2_�q����0���p�� �:�Z-�u����C��@��(0ɦ'�)�����ow[2:p*{����	�[�~G�s���Pخ�X��L�}<|�����1��f�c�WA���6�c:�w��߽�e�^���������V��Z8=(EdC#�V�N��W�0����9��D]�;L��cr����6�=��*�Kq+����/�:t���
�\;ɔ~����SAq(�6��xd;Ua��᫫�<c9f�b~���^O&˸��G8�N�v�C�&�wmK�o+5\�Y�W�9xA�.��<|j�mk/N��6�g-`�85+���[���7�=���Kr�r��1�4���Ho�Z�qٍE~��ͮpԾ�C�un�f�;�|�>�O*��ꪠ�lܿ.�<(Y�����)j��\��Hr_#�e����>4#�9�2���N��{F�.������x�#Dp�����۪�Ʉ8���5;��C�BV�f�8��f^h�9��W�8�Zt0�N�6�|��:���u�#��)��/c6r9�OZݘ�p�d!"�:H�7(�1WT�_Jld,�x��U_joS
���1��g�E�C�d���x	j�>�ʩ�Ý��n��y��w����������v�I�ڌ�p��o:N���D�%a���}Q���2�fd�RW���J�����Fm�n��n�\�#�t�[$1g�F�� ���D®T��/�����8�r��E����y����.��3��}�j�dM�\�V9���&��:�p�-�]�¥����R�q�݊17?i�]d/���B��N���Y�fg�X�XN���w�.�� E��A9�Dqa��n�A�{�?��Ў)/i�Ku����yy[R�\�^V/��n�;�\_���<��t�6����e�������׸nvQ��t������WӬΥ�:H�bU�s)1vv]��-������Σ�{ȴvI�W��=�yS�x�H�ۃ ��.6�6_�/,%缣O@�i��\bTyի��UU}T������ץ��0�;#e�6���a������,O����pӢ|&�j�u��Ɉ⬎.y﫷Ƽig�㺣��z�n���|�����f�`��ݧ3�;�M5<��Fiq98!˚��&u�_ڤ#v~yj����g���	�V��iIj�Z�u��*�����r#��ƬWq,�r��!��2���ɵ�Ƙ�x|�QK��^WB�Y�u��R)�e>7�錶��?[�U��zu?���f��ʸu�[��#�V]1�k��e9Ŝq� ٰ�e�R�;=�g��S܇S��vTD���* 
ꌾ�{h��ds�Z�3+�P�9�#�����ϑuc��gk�47SlGM�EgĀ���#%�b��N����_�|�A �i�7��B���.��7 G#q�6+FJ���/��/�yҌa���㻖j@\_�a����:
7]qS��?G�i���1�86E�c��]���P�6޾�ک�}	��LL,�����0�.{\B�y���[��8�z.�"p�=����,�''mP\��^���2�w�x,��uO1�5�AV��2�򍁃��M7�nyt�[i��j҂�]6����w/^wR���p�OB�JU�� ���8�ː,��Dk)�]Dv��i�ɍs����j����	�a�'ZJ����x���7ó���وL�Ukޒ����R��t����M*}�$b,fl	C(e:�\���;j*b�pz����!��������f����/�ms+[���D[�d��ǲmbCgvlE��i�	є7��a�mP�
��A6 	���1P\�۟��⍛��t�]�K���K���4A��a3KV�1��u�p���C�(���YZ}�^���{N�%o�rgE'l6�"�7��կ�a��JUi�ؼ�׼���u�G�\��^w�k:�y���ɞ���}��5a�-�~-1Z��v�oؾ�:��s5X��?d�a���]�6k�W���T�A���,S�'LlCr�,Fq�*��Crf��R+]tj�pڐ*&�dmoGR�P��OE*�ٯyq}�dp�iX��Q�`RgQB���F�����v�u��ks��RSb;>�v��0ŧ�lv:��d�5�G]j��po"���v,x
�zL}�չ�t5R�n��O��s�Ƙ��7�y�wLh�WֆB��#n�)CUOF{`t]K���Ğ6�Gc�bVϊ��q`Ӓ�mX�O�jZ�C�_ X�:�����@�Mf<�	Ƿ�}�� ��M�`�"���f��,;<淘eҊ팬�ǧ�ʃ1��i���t��+����2�w��l��	��X7v�E�?�꯾����*�|���̳cյ4{��.=����S,�s�n���K��=|%�wo{3�j[�f��G��db���qU!�J� W�(4c�
xh���#�s/�T��e.�\�u�T>�pBp�Ӓ�lĤl��V��@��><��J��vϏ
]ud��f�Wg1m���g���s��:5��B ���&���0�|�t<7�+�b��_<ue��s'�x�{<9�ݾg��X����<�`�d!𪿎�ڮ� ;�
����\��Y�՛�y�F�p�}���W!,7�L���y +�n�����@1ܡ;s��:�%][Ý��_h���u�d�iz]�'�H�K�͖Ԁ���U�,+$��1tr
�}����V�:����1�n����W❮Ru������ϑ��K�<m���:��xn;5ݎ
���.3�P�6�i���ҍ]���u|�
v�[��^V��P��
7x딀K�/�9.�X�ol醀=�i�n�������|������[E��,�#�)S�vF�]3�ܮ�V�V����'��--�ѐc��@aZ��цvt�`Pu�؁�7g���6?wQ��g�s2�R7a�\��K�Y��7x��7r*}:Z����B���t�WA_���<��"Z�TBUy��V�m������~%����rg�q"���}�}Gj�Ӈr�D����Kyh@�s�k���_=�X/�T�}��>_n�o>��2���l��RK�Z������u�b.;]2n!��wq;�]pѐ�E|�ġ���;/��z�[���}�n.z�=?i�7�G�ȋ�t�_>�c�1�0kޣǯ)�%�����\��,8�h z|� �t�J�K�β�yyL��Bx��NS)y1�����2`daǶ�����z�P���`>1j��\������ɔ���ρh��b��4��R]fW�����z�΃�7��+����}����iW%þ=���i��7`���O4vә��oO�W��9pXf�p�t�7���4O@YuSu��e�-c<���meC�NrW����AϪ7���	��q��/����2*�nF�>ީ�Ң������C��Ov�v�q�	���}�3�mc�ٿ���V:�"i�AI�"�ێ�q����P�<]c�p`ŌW�ӌ���9�5����C����K��+��PقV����kx����m]Ԗ_�
��&�#����V�ݔ:����3�ۚ�ӻ�2
Ǒx;e�mBJ)(-gm�"��5dGLn��I��Pw���K��<�ڧ�Q�o<�Za��}}WF�׫��
�ުOꢾ�7)G�Ȅ+!�i�����jd�:�ޞ�YӒ�Y'�k|r��SkA__FP^���_w���+�p�3
�*0u}r�ɨa��(<�J����jھ��*u�K����2\�DsL
u�U���=��)ӓ���W�ܣ9ڃ�'k<S�w2�������.#�q�},2z��P���/�ۓ�O����u�3�h����dZ�0v�RS�5���7�Gpxj�˻���i�m{�ƪ�f�Ȧ�ԍ1�m<9�J]�&��6(n���d�C�F�E����7f�R��v}.t,�����#֜ḷ��UHG�QI,d��·&u�\j�"V��/S���L����-<�u�uƤ]�}�[��t0|*�n�������Ã��W�Z^��f$R������Z� ��e��h���^U�.�뫞�m��Э*��tހ�γ���v�9�.�SpP�j�˗|�mD��i(Xx�i���co�W|
��{�#tMVG��h+"ĕ)�v�`����<QF�TB���B���e�
�Oa���Y>�,+�9��Bݝi�*t��U�6ao��t�a ^(n���b������LXkr�2���o9n8k�QW��G�,^�r���R[;9�6�j�og	[���VH�L��ﾪ��⊋}�zT]w.p���R{P�u/�Q/N�kW1��	G���ͮlVI��{��`޵��`d�rs�e2�ڄ����$��7 G#x�p[�Q���WW*�T�n�؀˂�23f#�`�%��Y����YILI�a�#D�t]�Z�:��O^u�%��=�tC�wnLg�!�%�\M#X�v�T��#y��l�Ռ}͝c��h��نNMBs��A����Oq�K�T׉��!||.�&�B�J��جk'�lsٱ�
�|�ߊ��R��{Ψ^���ߴ�u�-����Ŵ�N\���D^`��]�T�Z��QP5a� =⪆3�M�Z��,vcVǉ�Y5�\y�[҅Q-ڇf�c��5ݙhbUR�pB073;d�;G��"s���Kx~��D2�-��(��pd�1�	b��w#��2CRt�L���c2�
�������q�eVr$ՇC�E�T��xV���ve_!�W����u]_��ם�ˡ�W:�mo�Af�g]ы0@H�s%��P���>u�o)!�AW<C��n>t�u�J�D�6hѣ):,nHk��A���ԣ�t�f`q��G�����ސ!���2�gLu.��|/�H�
yQ�b-ަ�iX:�ۣ��h؇3�*��0u�"��w��|��EME���x���Ν<��u�5O=C"=�{4����Iiv��j2n����-�O�6��\�<��ݥ����s����FZ�o��Ⴔ�t`
si9�fЩ��54+�ޕ���!݃sq�7�[����AۗZ��٤wAi�R,���I��L{����w>�Ya�G��H��7J�]�h��y�!�7B�JȺz��v��\:
]�{Ж_<�o���)�{�u�׸��.Z�}땋3�sbc�Ŋ�� Qʀ!�+/�W;���}��*�ôz-�7}d�_EJ��8����K��}ޙp[�܆�M,�r�����V �Uʎ���0��:]�&+���ʺ?c])�'�E�����A1cq�É��'96���wWhА�����AP�7k$}J��6�㸐��ˢ�YX���(u��Z�7q�����:������>T8M�lM��|�f^���(/�%�;ط��7Z{*b����zu)��wP�SNr�i�r�J�FN�{[�9��x-��<Ƶ�T�1�z2Y/,(z�ȷ7��Ek{�\ �����`�(B1�~P�W�p�����'e},���LP�ު��@�⺎$K5vÆ�wMe��'�S+*� t�n
�ub�%f�a4�۰�>�QU�>C�1���v2�6 �k�ebcB��z�-���bIsZ'꽗xၨQ�P�P�1�Y��'������܃�N:ʙ�G�Wճ;�h���rz'�C�~��-�� �>��T(#7Gc'H�j�P��Ţb�+�3zn�[r�{7��Q��w\���v�s�Q�W���S�{��hNN�J���Xi��&=fR�bO_/R��8���.f��P���jm'x��* fCn\r<ٚ�P�W�V/��Ŝ"��<����w�����Q�����|����9ӭ����gNB�R�}n�����vv��}�f҇[ʙ�A��o�!B�[(r�Iؖ�7���q���_Wto5�Z�K�gs��s��c�#n�]G�↖o,��gn��	RJ�t8f냌u-��XM��ۣ�"IßJ���3�Ӊ�x6���b;S��������P �(�	��{z$u�̜�m�<un+CW1�g�R���?m��K�a�p�=��5��t܃e\�,�E���T=��S���d�x��%]j��r�V����#�xȣR�P �M�_:瓎���CܽurH�H�*#R��ĥ"�В��t�V���9�T�P�k����FUi��z��$��%����*^V&��+�=w�'',D�[)*J���B鄥�(��d�Y�,#T�����3����V&�p��Es�NN9盪��gs���;���I����-LLI%ݹ��Esܗr,�Z��E[�㻲��w<OK��fe���ҍ�����Ii��:q*��B����ښ	ӫw[�Ts�ΐ��54Jk5\�tĉ-���SB�6dm��MU�OR���҉U�p��Y�G�]ɨ�sZ!�s�9f�e�9��%*�wwP�s��'Q*D�n{�e"�a�UV`a�%K���R��D��ODWeQ�fA�u]4)V�	f��w#��MY)$)A�S�V�|T�$�D���Ⱥ�0ojڔ�JY������t��f��Ү�A��#����O����7&uۤn��s�5�5>ͷ!� ?�����䰡�x{�p�ҁ��T�r�\_"a�0�I��T�D_D���yW�����ܢ�۹�,�}kxԴ�OX�! ?��a2�l7�Ú�(�v�1B2�f9���xs<ն9n.8�.t�-�A���i�Z·F2�;|r:���3�W��:5lL�_I���˔��&r�gi��]eC�B�W3���}�x+=�7)��a����?>Z.�[��Fv�EFfg_���^�ל���n(΀����>�[uF��kS뇐��0}���r�R�x�lY:�!�-�V�{T8���B��r��<�s�A�^�N�x`N������]�9mW��!�K�$YA�j���{�7NO���F�%��g�����*a��ɍ\�Vj�鉭jY���sK�w�`�:9d���FhDKR���bZ6`��T�LQ���\��
�m$�e���x��B�b*,�
��@w��0_��n
����MEc�uR����ܑ�K��^��e�b��7����1p�U����
 v�y`Z�HP;�FR�(�Y�B]��e������P��|��u�֥��r�-*��tFcMrk��0Y��dQ�a6O���r:�b�U��33X5���w�H��"M����u�*�z�8��ͭ:�slu@��R�!K��BIn>�����Գ�8������γ[h�.�;���W5��>���L&��\Zw���I��Ϫs�^a𕦠[�Х�ѣ�Ԁٱ,����jݎJ��)�c�U���u{s�(F��qu�U�eY�,���zO��ʇ�ZA���i���zx����Y�����@c-�N�������<)�/�U��W�4t���76�6i�΁آ���D$Q�p���i�1��&8]D�B����`6V1�d�Rr	���y�M�۩�:�;+|,W��m��U����
��	�=���Oٟmը�˳�͡�����G�T��t >�"c��&��{;�������~�IQGyRxqG\�r=��]�-y�i|�?�z�i��R����]m.ߛ^�u�Hk��M�%����X����{����ƃ�p3ҺU�>T�=Sq�ׂ��')�'KJ����*y�5"b��.���u�͐%��:�Pw�˗���f-W�a�丹�1W�b~�\��έ���pl�g�=�~a
�R�����n���᤿���)T��Y�b"�=���̂��F�2�5W�3��M�8�;�ը�6g��Q]���WG�xW����{tY2�d��D�;���!�Zݰwq�2���*�+��ە;jWfq�\/rFEh*8�=����9�,͓�׽���Y諪�@�v�R|���=1�c�_DDDG\�i���{�b=�vV��M���ܗ�r d�ݼ�G:�~�?w2^}U"<Fg>Ėv��Zd�Kz��Է�+��.8H�T��r��� `���2)�f�^x�e�$���w��_eT�^v�gv�%����˺�n%T6nY|
�Q�)��7ח'z�9�˕�ÒC�A"�0b���ON3�9��Xk�N�o�ޗ%���Q�L��w*�v`�}Y�)�=��i�_(�S�y�VC��9tz�5��J�7��M6�z\�d�eƤwq�?-7<� <�T�1���>iV�&�n�A�Qxb,T׆T�&o��궕A.�����N@����w�WdM=���6&~s7f�L:p��T�{c�o<}�Tj�S�v&�~`�t���dt;Q�Pj��π��t��o>	�n��K����l�A�9C�Y�~���}�^m{��JT!�����zg������)�	
:>���l}O~��+���/W�c�;�ھ��:K����d��������e@�i�.���\��I:c)ר!�.u�ϴ�`J5#�fA6��o��q���$�'��ɩg�l�z�.z:���SK�
�װ.ŐV�/�d餔��#����mr� 1O�֭�NV��i{��qv���.��y�S�x^Ou��%q5:U��
Pނ*{��o��u�&��?t!v�G�u�Ƭ�������IoR���.O�!�څ5�7�k�=_�'���|�[j��#���s�	��'#�ٮ�Ɋ*�7��m���/65�=��qd��U�M>u}�޾�ZW���c��-����S�
��+m*&�c$������~��'.�u��R��#������7xC嘨��p!)���za���w��R�4V�0�-e��\�w���X����b�G<���+��+^Xۺ�s�8��S2f�C�Vص+%���WZb�棥��\Y���u��L[���y*��s���M�Za�rt�5l��n�a�g��e��A��X=s*m�}в��R�u��;�vt��c��m���\%�)T`����.�L]�|O;t�Z]���[��s���GPC�����J�"V��� ������*�dJ���$�g��k�&Z��x֛���2�,
�޸o����=�4�ma͞�3��׈|Q���;?�������n��=��(�ٿ>�����oT4��- ��a�y7=��k�j�b����ޛE'�W��+3i�uڵ�]DcCi����f���^>D)����W����x:�'�~�_^NV/	��Q=-�r�q�n���Ќ���r^��𻞧�j��6��=�;���(�z��]�=-fj�}�����bѓ�zl�^j��m#T<SW��{-侞E����J�yܹ�������<���:�ί���}���|*�r�+T8Zg.ab�d�O:k��U�_s����Sz�=��y�e�x;��Rq��k��N���)2�_=W�h}�s�!�h�֤R���t��y� ++���uC��{��Ptlm�PbzK���'���qh��7f�^sӼ&�/&�j׻/6]��=]�*~c�^��;F<�|��WBg�coh������Ѳ�1�������M��i��%��Êl��K��7
����}�ʬ���j� 3��ׄ]Kܼ[����>7�S��c�&���
v풧�!�'~�	�����K���Mb�wG%��G����s?�ꪪ�����g7A�J{|���)1���0�T9eDOL�}w�\���=l���\J�1�n���0���Q�q�2�����a��
���Q4ǽX��{����%��4��ʝ%s���\7��݉�"%�.�+,�O#l�׽IE`μ��Y��f�.�U5��*�"������M�m��U�2��u�~��=�W1�Erf[��Z�-�)��W�]�uv���`*��eԾ�5U�U�q`9�'?ou��3es�ws����&���:��x{.m򻘄kh)�Z|��ޱY���� إ���*���K��P�T�7����*_[�;��Ti��\�JoL�<X��q�./��|�S��7�/�c\7n x���{_Ԟ�ǯ�o+<b�Ş��=3cc��8���C�[��SW�Opm�4�y��̫��Tչ���:V{ �m�Ly�ZE�C�h}6���oRS��*���/e��ܡ��]R]D���/wu�Q�K�~�-�݃T?C��.:���;Y7�B.�	�"a ]Z�	jd��-��tk2	׬��
9�����9�J�/��W�}TT�I{� �e~�Mͪ΄/"��T�
�������>�m��K�mU@;����u�,�qa*��6�TV��Y�a��:�hn�\����[o:p�{��R�Y�v�7����Tk��Ҡ��M>J����4�@�;==�G8����:�ƽ}��R�բ�cp�m��1)p�{b�{{���˯+5���޾E�x���ю1�ob8�KwS�=fQdy;g��y�U���GJ��R���q�z��-�<�d�r��������,�P��[�;1˫ .˿�9��q���u����ˇ\��If9wQj.}�!S)�[fOղ������$�����|U�l�� avf�η�.
܄��"�
����2Wd�b{��v�k^�����v�\���Uï��i���*��t�F �a~�`��ҷ�/��o��N[�i���.$�['N�r��D^c��d��xOK˼�EҷVӡq�����E�H�Ʉ�5ڀo�n¶��=M�qI��������z�ݸ;%o8���U�ŷ]�ՓƮ�fh��}_W���֚.q�n�\�^7�V�������aX빨sW���򹯉��;��q�ײ��j[Q�A��9�+�k��������6v������R�J{��';uc���E�:��ʌON�Ȏ�n�V�-�䒺��9��]�x�9�@B_��YrAx�SO�m.�����}Y\LW^�Ͻy��|k�&�Y��O˜άhڐ�^�⡬�iں�mWL��O^yB3wtS����
��7��V���q��t�M����U���DXx�y=<��<�#��=�����5��紦�&��[l�5��k�)$���%��o=w��y�ժ��f>[���J�M�\���Q�������Z�����7':&+_T\��rM��J��쯭��)�9�w����t����X�����GeIs�Zj�1t��I��7:P����9����-�i#q|<��x#����K�7A&�"�V{-�P:���/]YWz-u.�b�,�`H]0x!���_���-���ie1���+����2��+j�m��ԝr�_m�}K���iZ-���b��/�s���	v֝��i;��}3�����ꨏ�֧����ތ��l�*�%P#�T��W���/L�G�Ὤ��<;#��X���7x�8�p�)�b�☇υr�g9���v%����羡�<���ۜ��=N��������˰��[�)/g�������?iY�����:�y\���ơ����TC�2���C=λ"�����xʽ�<��hN�x�ud�QU��i�x��p��&�� C�f/R*F'�m�yPR��ዕ���sw���W<i��,>!q��C��.=uN�e��k.��ߊ>eb�߬g˨|��Պu����`.�b���.��,K�ܢ�*+�����F(��3]e�5�z�\�@l>�{��
;�'�Ӵ)=�]�Ys�.8g�p�9�<���R��A��?z���y�]�7�q��ܟrŴm�|���<�6l��?LL�٘O'�zT��Eyn�����+a���v�>���sR������գv����9���� ���G�1B�
Y;+�%�U�{�1j�^Ke'���K�Ŵ�.�-܀Ax�V����Y��\�/W*d�Ups��~�">���d-X�O�+j,�[�\uV\jon��q�u4����� Uk�pyљܷSs�j1v+G�Z�E�UuQή������>v�E��hW�}�++PT����%TA��P~�蘧�^u'qϝF���a�B�Z�����5�"�n�c�Vݍ*�*�d=��
���tKv-K�$����6�(��k�-qٝ�8�n��6ʸ�	GB��9�*��pՏ T��Ox���@��������|�8Ɉ�H�n�X!��������+ҏ���\�z��&�č��S��aގ��}n�"�p�7{;3�BԒ�q����bV�Cw{^�-��lbf�
Q�\U��U&S�a=\�`(W]y�����Ƿ_t����Ǯx�U8wϧ���L��������K�4��1U�3���7q��-�c��G��8&M�H��B�6�	��(|�2c3_��D�W�)b�ȩdO9��TRV�>�"���]�һm�Wp��Re%m���i0%�;\�U��z��%�����H}^9�/��
���`�˙�;�зki��:���}f����R�Pr����}�2�-�6��(&�R[(�O��ٹ(��<9��p=��2��V�{V:Q�\,7NԬ}Ѭ��=�qXo���^X����I�Cnﮤ�А<'dGrj�(ˬ��{[-9��2��_+�}�cq�ǉ�:����+Bs&���p�SV��KE\|��6Yoe�rD��PN��	Z �q��CN�tw&�5h��f1��WYη!�!�s��5n��i�/�&)��Uywf�����G�b>�yV�Uogl���ŝ���2Ҝ�Td���]v]�i�aU���N���)�/�����H$��
=ڒ���ʬ�u�gr<�5��I�VI֐�q�fa�mإ���ݧc�\r��PBzoq԰T���	R�<����a��\�b���ʆ"�}��dm�h[��j�-I�N�\x��`;Q�l�ದ�a>@�t���o˺���>�fSJ��h�}��i`�r�8����uYh��rr,(؜�e7�^��D�mM��i]Z�j� �o�N�ZWU�#6g�j�veD��'y�s����[s�)c��q�]р���# mnj�sSr�KQ,a�E����#4	�`А}�u���"��/��.�dt3v��8����͍�$릒W�j6�d˵�B�	��"�R��x�j�O�K�d(�y�|gݠPk�9�r
����W�`0Ɨm]6����DZh�(_3�z�B�*e�pC�m]2��]-ΛM_1�H���]�L��Q.����$qͳƐ��go��o�q	X���N$VT��NŌ֕���9�*թ,�}w�л��"��"��y�Y��7~O�aU�ٯf�ۈrZ��ާ����6N+��p,��5�����"��|�vq�g��qꇲ�C��0Ԡ��vB��C\���R��o8���������"˰��2��F�G��A�Ǚ[��ﱄ\!�Z�w9XCc�i��٩6>{8v:�P۴eA��㝒]4t(��s:X����~��kn�]yhd�vy��v��3a�zp�-�h`�࠻H�n�-+���{`<�23�7���dR�Dɛ�6���)}�B.N��.��B=��`p�J��oL �k������[�R�� ���ܒ����Y�:��|���I�Wwq��iy��;ׄz[bɥ.z�p��p�Q�ەt���˦v�fx��/�ҩq����VԴvp}�t�c�. 3�����v�^�!�6:g`�i�����a���9k��o�;�
\2��A%�=v�h�Ra'1�<�'U���q�"���`�p�+&�Ko����f՜_>��:��U�<�:y&���t{p�H�E��o,=��u�2��y� �>}D�6�H@�����̩#LT�j�Xn{��!V���Nd�Z�d�FUV��]�=�Gw\�$������Wt��+��zUQ�����r�5,]�I�'H��DLUD���UL�s�g.�IAVNN��zhNn{������$�-<���LV�'M�<�/t*=q��C-N���g����YBEG5#Y�̰�A��Zu�j+���u)5���<=�2�Z���n�zz�)).�N)�Uf��u�wg��去��s�
J�!��BK��B��⪅Ú��rGq)0��tTV�a���RXh��C�J''%m%�9z�1Z@�H��!R�J,�9�Xn����A�6IaX\/tQ�m5������BJ�U�x��%f���CB��Ҋ�S�r�0�(*����j�9Q:S�^$:���HH��*���E\�"�:*Y}�"�� �U�lM<�In��:�p�8����[{��O���j,�v�e��sRbV!��Zh4��t+���ٽ�����DZx�HT�΁bE�Q�D��ː�	z��9����^=wf-,/'x��O6�׻�t��%M�.�ⱡ��T�b��u�W��4LWc���,a����Q��G^R���s���QQ���Ϛ?5�������l����GׂԎNR>����Ӌ����>��K5���,moCW�=Rrեۻ|nbU���,lݍ�n�,��r胳y�{ق�nB�?R�_=�V�����kW��%}Ɓ6�:��v���u��LƝ������aRs`�1���^����5�݇��ؕ_�5�w��$MGnX���X<�;��pPi�L{���sg��3�w��v�aP��"�:�ЕNx���ܻ/J���i4b{�J{��0v�5�YS�{��Xb��EV�v��c�$��+�<��t¾�E�w�Ĝ~��Y���}�� c���#�Q�])@p�������[�}
ҿt��(���Z��	b�v �#�D�R���_>��;$�E�E�e���41�[�lG4�;3��ԭ��'d�]��Of���yp�F:�F=�'��VJ��m�Y5v�ƨ(����&�DkN�E܇��3{���	���`b�����}P���7��)kp���� �o�������?-�%5�4�
�.�&+��w��e�s���+xW
F���]���R��� n4l���n�Җ%�ѐyo�}b����w�w�{2ա�F�J��,�v9����'3��P�.�q�&���	[W}4@i��3���V��*��\ZJj7�cz��]%�ͨ}pT۸
����-�ކuR�.�9X��S�z�Z�ux��V���%v��]E��&ƴ^�ot��~�s�u�r���#�o:�j��}�鯵A��n����pfwe��ܶ�3�ƨԈ��ڵ:���[Aqӊi�*]G��Ԣ�~��BU�
�<��Csޮ�oz�l�rᴝ��w[w�1�qË��^�]K�+�@Ͷ�b��\�V���T<Ow>�{��znOm�u�c�Q�c��S_eZ�	'l&���y�0�'�����p�tmb�JeFŨ�S��$(O�^�Vr�\����P����	������2:o;OEA�mCCr
s2�VB��賷�K.os�Z�*��޸pq�z2�-R+J�3�%22�,�h�$��k�*vr��������}��}���>�X�᦬j�A�w��T<�������5���TstѠ�o9�7p�^m�5��|�EN㲓���5j�Jyx�wc���vl�P�z���Z!Lnw��d��^��Mo��;��k�NG��O�g���\��[Eަ��YU�����͜1�ᄣc�$���¢�Yx�b�iI���a-�*�W3�N*�v'ն"�?�c&"�5q�|8�ݷS��L˞��_O�$�)�� M=�{��g�f%���;��x�q���݉�R�\3u����W��yq�G}0���[���ӽY�6/_��;�=N��7��݉�R�Q��padI\�����*u�=�7ӯ�w�^Ds�)͛񟷘u	�;��=��!\:���
eP[��j��8<��s����~�Xg�x��f�PU�)�z ��U��5U�1.�V�k�����S�|��47ȣ̯��]�	��/�S�jŏ��c��3��bh��[uj��HL��:�J����*X��B�p�g�Z�tp�=L��1�j��(�[��{wK6���/>�;o���6�.�����*�h:+�쫴�[Y�v��Ù1�Vd�;{�2�U]K�V�b�]Y�=�U�����>���Fg6e�Pr��烱t���-eA���xnׁ�}3�e�`Z��o�ͥ�����s'��3<���ܭt�e��.;G϶���s�oV����_hR�op��d���w�w�߫���5kb��y���&a�C{1�}Ϊ1F5���sb�[�w>m�r���Y�k�g�nWWW5��]��K�ɵJ�=�������C��r��;[�*8�"�K.�j�,���]��=KYz1������N�ko�d�'#���v�nR)�-�9���}q/��n�� ���Aލ�|��[�)�ô{M�lYܤ{���N>텺��e��qB��%������*vCӴ������׸�?/6v{�hr�n5�}m)Nk��c����j�ɒm;����zׯݣ"��%�U.����
��LS�i�e`��"�h�Wm���5���5:Y��-��z�75׾]�{�/Q�Ւ�޿��5%�sxT�w�q�#��5W���Ҍ�qx��U���U�a}DLf��� ��Vu+\� �E�/�����m��%���9Ӆ��rHu�M��������0�������꯫7��e�l*�,��ڮ�≯	��;�]�þ	CP��sf���ٹ|�2���r?q��S��w�摪��F��|燶�龯�,�/)*��S������O|���xKc:2yeo��K���9��WӺ;���3��*5 4��n�9V�a�`}��T^b���q`=y��Y5���H�SL�o�f�����z����8޸��D��a��\����޵��6���@�F����ĸ���?g�9^��J�23���k)>g��ĽX�j_sUy9X���Tuʍ�B���kg��f0�4te���|���9x3�"�:��Tb�u�mv�b�x�-�Uc0t�out�3%K�[J@b���yX��2t��+���V�8���B�̙i��W��Ac;��-���k�\߻0%pn��D�5�TY�Qe�uǴM��g�^0�(����w::k�!9,��S��B���<B\��(j��q�G;p��o�p3 �c4�il�8��\r�gdA�§��P���#tnCn�Lx���^��TQ��ቡR)u�����O���U��^��� +T��
���v��G���T�"�4���GYp��ېޣ�y�}obU�5�us��{�*U��Q�d)�/�3ݧ^�Ҟ^8[��Fyom�uP:;�e�{Jb�e�z���q���Z���֥oZ+p���ڈr�	p/�p�o���B��2W�$��5���*��;P�sq��1� ;^P���6�]�+0�0�#%B5eD��}Y�]���.�PV�d9�*]�+{a_�G�%[c�c��ί��'�R�W�5�LEp1��ߢG���;��w��#��o�l��|�z��}����uD7biK<]�me|}c:,��E)��o�<:ͪ���D�+�j�����xʸu�KLp��_e�Y.ŵs�MY riWr�\�#8��}�'�zq�ɸ;H�AX�/z��X��x�?t!/PޛE'�y��c���w��.1���2��fl�m@>��N���C`�7��=�9��}8�thPfp,�c��{,�LI�&mT^>�O�z�rS�S=�:�V���j���w��M�F_^#Df��!��9��̝]ki���. G7�lc�3:�t9��K�7s����ufi��2�OF� Mq�K���興����� ��{���]�e�W���Q�u�w���si(ۘ��j��^>u�OY�z4�����=�~���6��jQ��F	# ���	͔V�xu�*nVjy�����j߸�Lx�s�Q��B�;V�S<�챎���<�o���r�njl_7}��.�n9��PHm�9��qq3ۜ���Z�5�8�V{���[jm����=��؍{��<�;R�U7�gyyy�(�UgN߈��'�ϋ��s�i�e71J�QQ��H5,��x���3���z��vT�2�LV�W�s�M>|q�D����`+ym/s��Ӊ��>�5��F�W����Q%��R�Q������+z0�h�m�Ku(��W���+�܃O�S��4�}�@�J��~��*�x��d���C���}&�/�>��<q��݈�Hu3h�y\9L���T�]���Y��NZ'�M�LV m�jE��w+��o7z��_\�z��F�}C�>8�p+��"��"����h4l�V{��������z����4���$I��B��=;����Iܬ�����gC�	���mY���Wug�z�T�����7�'���I�sQ�w�����;놞ü5u�s���>�k�y�t�Wﱵ��f�W;�:O�����WM�e�dix|s�W��7k��"�Y���rۃk/�xg9��d�v\�LL����M{d;S�}��JN�{��o�ѻ�޻�~�ho�G�ዕ�]�p��2n�8���7E(k�P6��S���o�J���TA���uy9X�D�׎�^^�ĕT���r�����K�Q�:��}�-�hn�m�}T�s_H6���OwH�N��nO|��m�Ϫ-�o�=\2����ŵc3����Zs�t��ݮ]�y
�e�T�kf�ZQ����ا��q<���xv�p�W�Ȗ�=Z�B�4��ʝS��+���pU}�r�7�S��w�!��f����R���۫�n�����:��c��~y�u�;B��NU��^�TK�>��A<6l�ת�M?l3�:y��	ܮ�ՁQ-4�<&X[��	���ʮ��u+��������%۽�.�'��;����*E�G\2�����ރ}�%��H�����Z�_1xFќ��;�ľ��X}�q�L�#����}E�Vc1�����GZڄ���Ю�γ�T+:�9[��>Y��r�M��ȉT�7�o�L�V$�˃���u�?s�;�|�˫�nTB�}���&�7-���\�������si^����-�w��W��в���ֲ��k-<�Ov\λ���Le��_.i\��F]#_5(�5�;۽�P띞��X�P��q2�;fGk���2�'˸����u���7.W˝C���-}�D�	m�y\.%ne��,+��]G6��ۜ����ˋ��׃�5�#��({办�C9���WvC:�O/��U}~�:PqH���f�����p����p�H1�u����.>aLG7<�w�9��|���=��>��8ۨ֜��K����e;��o�O��+���]�W�<t9�=��R�נ���t��������[���g�{Z���n���ia��X$�����6���d��N�P;��𺏋Ŕr7��ً�����e~�ǎ6@�i�b�q�� ���_	���wRnF]��Yo7�3��q'r}�j_N��p�cx2��$�gn��b'�ZkD/7��a3��ge��i��ߌ~ұj�1���K�==�J�����[�	�5�{#:]�u�	c���^W���u[��ָ�����>�:'8u�zT�/d��s�Q���w+l�	��d�\my�.��|�80v����[3v��j�@U��w"�ies�i���G�~�!u�=$��f9����q��8�c�F�����>�S]�p�>{oƷ�Gң+�p`���BoJ�Tې���Ϸ�c�����n!�Qj�Xв��Ov� .���w���oi�b�nZ�3܊�|�k���2�Z�n�ɫhJݽ���=�V 0ji��Bʉ$wh�k�\b�X�����֓��{u7
�Mv��%�:�p�)�+ BR#R��	��]����3׶���a�^m��A���C\'�-ؘ�(�CP�W�W+^X}�����
���v'�cT��og]�9ѓ��}f\״�	�[�oR{Y:�Jl�[�S�y*�	wd��97zM�Z�����vz׉jtX5����t�����BMk�ڄQk�Y���x֮ӶA�p�E��޻u�����ɍ�S��T�6*�f�v�Glkӎ�-� �W�������iq)�6u��{׎ĸ^�2XDb}[�*�m�v�Wiʚ��XI' ����q
=�s໹|[�^�C�$&:�q/_�l�@پ��7���)�;t�Z�7Xp�8to�.�:�ے�H��bn*�%�����V�'QK:�LS�{�{"��ou5n�f��i+�5p#�[��L5-�9sz2���2� ��7��*�����)t@�`9��S��"�CWa�����JT��U�vh-��9�;Yg���_J�
�����v����n�Y�;����Yx��J�2��ɴ`��4lc%W]OG�WM�y
���vpk��_�����<�HQ8�U�T�X�Cx[�o9vgd��}�%��ڭ�(��n�oQB�]�ҴI��������x�KJ���iέ��:�-�E<5��K^�y�H���!��C��S�������U�=�>9��i ��iJeޟ�Ĳ�i��Ӧ�g��N��kD�R��of5,8�D2���d~�9�s�}x	�K�U�z����SV�=�KS�c����;tt\�.����Z�Nԝz826�tז8�U����윴űܭ�er�����e��>�9���p�ըS���.�ĭ�kkEn!�#.c�P��ϰ�0���m�y4�vݾ����,^��0�A��8�\����ִ:�dp��0!�_.��Uި�C5E�k1�q���p�w`�t7]%g>h,i���S��zm�n��1�3m�{6E۩��
�qWsq!���+��ʳlB���_�9�Qٚ
�$�P*Q5h���r�0.�-��7���V!}AS��X�\�('v��y@І}v)�[{;��f�gs���ڞP�g]�wҘ��9Rƶ���nvtk;��z���7xz�NZ\p�{qI1�;4cO@����v��g�6^�2����1j��Zs�� ՄK����4F޸���j�wG�^p�=��D�ou��-�4�]I�]\o�>ݩ�mK�ܴ��)�|0q������Jh���-�_%x�h�TM���7�}wJ�:,9�E�Q� �������W7�F{d1�7�5��r���K�Q�)��GF�Ж��:j�tM<�W%3�ɜ�9�P8�kΙ�������F_2�˦��Gn�J@Ff�Ʀ.b�Հ˅=�l�W(����1cv*'��c�V�3���%�a��vA`Po�������a,ڰäŔX���]q1l��y���T�I��c�#/�x��ݖ��/i�Il��q78=�^�˲Q���n
=7z�_.��|w(�%\w.;$U�E%#(��VWH���D�J���wr;�U��L�"�;�T��˕H[JL�,*�Yd��2A��^���P.R	��%�k�^`�T��B��E
uPEU(��r�X[5e�TE�z㕢�	�K:k5
��&!Q�.�<�$��*�6Yi�1J���ĂNFTYXPTf*�]H��J!�e�d�"�zjp�Cg��e�4��L��Ԉ���\=H�V���U��K��D�*W�,�R���T�HШШ��i�
*�L�*���ԋ2��D+,���,�|v�z	=<ܮF�R�*��VJ��"���,����5;UJ�!�I&�af�T\�EO7AtN��U����qK,��t�3k�I�UR�:+�a��#5E�����S��I��f��{|B�]�vpl�N�,���\��lbc����/6��_���VmҺBN�«K�ʏ?����g�ɞ����H��������Gl7b&�+�+�ͬ�`��S�GJ���_7N�7��f��W1�A�r�5l��A�KLp��}�6ƚu��.�L�˫z�\F�;Zw�x�ד�AT.���OB�:�RU��x�ػ��z�B����<�/1W׏j5h3�UOIqX�ک9��*.+7�+-��5B���죊��*��r�1=5��[�-�{=W;7�}�T�ҐH܃��f��y�����UF�����&�B�*�MTgBnvé�	vj�3y�{^�m���9����r����$���y���<�'�g��޽�.�~Ե��}��f��v4-���Q:	���ƞ�ۜvs���5Nn�or&�)�S[����tzy�N�6�wR�ۮM��'�C[��=�;�,����c����x���)g���v��q��\V4����[��碽%�w�:�5��XQh#�4�"������ь�����5�����J�)l�2�[lҼ܂�q [�G۽��� ���FP�G��]�Dlmduϭl�V|���Z�;dM�i�b{M%�W����ˣ�e�r�﫲���gmQ����{=CJ�[�Mb�c����ҔQie
T�{h�u�	\F�P:9�����]�`8�K�br����/V�k��c��t��6ʸ�	}��왕s��{����`�V�q�w˔�sn�s�R����\�c��W_q⩘}�\puuo�e��<���v�F̍vht�r��e��]ϡ�S�8sw�ؚR�Xѓ��5z�;y��y��0�k���8�f�s�ô�M|�7N^BIr�Ce�5�X��z�*��>�
~��~Ŏu^wQU��=��hP݇^��i��213�{@v��.*_i�o��R�+�r��]�ٛ�����׏�m4��qy�;)�um�MK������V��I��Z�c��K����<����.;`��t닍q�.�+����m� ��f��u�V4(,wAq#�΢)� ���l\����҂W��[\��2�C����|!��x�q�B�h��"�f�N�i~��o�Zx���.������e�q�j�K�����t%�cK֗|���}*ӻ��#Rt+z_��֠lmr|{.�g��U}Vp��������&-��)q}B��s�����!�yvo���Kj����s�aC��]ގdNG�Z�b8sZڨ�b��K��lT<ǻ��TCW�z����sa�8�����W��7���ږ���Uq�E��G�^�v�Rˊ�j��u���D���ݗ���U���rt;(Io~Ρ��v�8���Se71������vJu��}��:yЦ�.5`�|�;~���c����6e���D�����\�j��o+�)�����8SM��Ls]]��u�`�[ý��/�>��ي��e�}˲�򷳱ͥq�;v��Kt�~��r�����)�懶B��Z,���93�]�;��t¾颟u����?S�sr_LC{;\%�P�sTw�o8�WL-u�ve��9w������:�F�����2��w��'&f��ʎ3�LS�b�������r�2�'�@W4燧�� v��;[J�.
�Ƽ�ĭ��b�����:I��;P7�H�;W'8]Y�9�YyS��T�t��7Z<��낊ۑ� (��{{�
�nͯv����	Q�yy*������g9�Z��M��-~������Y��f�m�e�>���V��g�+�`����s�v����֧����W�i=���[�[�Ci���p�ે
@�������]B	�[LU�ǝ7���ܒ^惉f�P�K���h���	z�A��i��I�5���;�{��q�<W=��Qq�v�Gܤ8�Y���CX1V�Zzt'�1z���H����|�����V-\��j��](�x�t479U��c6>^]�]]�,��ڵ�9[w�(.$)�yF:��6���:�:�D}{(���1�"<��I�:-�5ok�[w�md�Q������d�w�[sy��/��-�)g-�Y��ۇ�9e��PΉPkZ�܎]a2�jS�x��z���W�vB���y��֚�?7|��{P�'���ΰH�g&�)^\�i��ENíI���Z�'}�n�oiMr�6�J��cn6@� ;��Y�.�Ñ���f�{2�b�o2Rk�Q5���6�=�n��p+sup΋�[Q߭�,�䂶�q'Q�|u�4�!!��<B�Sr�)>�-Y+�wKWs��u*�H&����6%9�w_PZ�aN��&���g�}��i;��|�P�[���S�b%�|�\b鄱���4�!��X�N�.ډ_T�čz\���O<�jw�έ�M��w�{�ˌ\��uK�((��G�A����������;c'�T�Crʿ��T#�6�����	OoYk0�����[σ�
�%4]�G�7.�'��+]�4E���u7�{u�o;�ʛ�2�#��9�ws!�v�b�g����)\��5wWxkb�mq���/��f�)͛�m��K��C�s�^Ŷ��n�hY�����|5b|������mZ�1��k��z�\KߛP�#L�7/;*�eE����{ � ��/r��uy����j�wSߕS��\�.��˵��)Z�c\F���@�b�v���ھ>]�V-]�6�Vmb+�<��r��;����y^e����h���+����аӐ͸$�ң�fhƜ��$�ΫJ���"X��'����<�2Kp��١�6�̡9��f��լd��c�4�f��B�O(m⢷�On�z����6{��7�h�-7>�d�q��}����_�c���ĕ�.ˇ?����׹��.o+��Ǻ�1�u�`J�~]}5��M`ݸ��8�R�i�o]���y�i��8�8�X�B�{q��x�gD;�n�5�Ya-���SQ[:y�H��e{�ooi��:|k�M��\nC{?)��k"���dv�ք������5�j%A�֬r]�Ύ��}��IS!�;ƢǢ8�3��y��4�7��쨕%(��ꋞ֟3�n�1��S�7]C=�U�<�F���L+��Q��U������.T,p��;���q��#�r��	�=]NI{�W�w�dӤ���
��U��Y_OM�{jst�����f(��*ucn�&y�I]����q�������b�v'�R�[0�y�S�]Ի�3�Z���Ŭ'�e�ٗ9�I<r�jp��[��������9��nwR�
�8:�م����'��
�7�u�}N�P� ��i�Q�>bkn�⁭��yrt�ݳ�|�*W{�nk���C��h��!P���[n��7��`�|�aX���m�싓��X��h�u��MLGs�LL_2]���y��%�2���ǎ5&�><��/eC,�KVf\���e�ʶѽ��~.�q�xy4�3��nOf��"�l�S�:.}�%���Y��F�����	v:'@�*��\����!����S&�Ld����4�Q[�;��S�@\|�$��4�1T^3?b�w��N�јWW��8:�]��]�@چ��X��Ye����y�7�54:9[�Vj���9�3NX��7�=ݳԾ���-��v�v�=�ɧ�٦�ȯv@�=����E��8��z��Tdrz�g�wUW���j�d�<��M:�N�Ӭu���*�������y��عn�!&�{��=L]�؁�����o��OR7�h3orx��B��T��}�7��c��:��v��3��������;{�*��{�uk�*"v���W�b�ߞ�	�/���R@N[���>Mt��R���ak�=�AQ�R��;�Kf�-�Ia��<���[/�Lsi���r?/Tl��y�)��PY��T����Hr��)�k���D���V�T6���o��,�+*��;�S��d�Q���	���������H����WZ��������aPΰ�] �f�G�ZNZ�j��*v2��3*t�c��y�s8�Pʚ(D72������3�ؤ�]��39�{���[m.ݷ�?�����t����G6��awd>ݨr��g����
�eg��WI���OU\���Ǚ������.�W�!>�o8+�0��e�Ӫ�2F�����L:�5P!^I�|�O��"�{�W��*ݗ��Tβ+&;9B�J��`��a^�E����׊����__y#W�4��"rn�C�n�
h��Y��j��!Tv�w���C:3@�ߏ��]�7�C٫|�O&%��Ux�
��&&bP��W��'���_m]��bc��]wlUk��UK�l����x�����AWˤ�mA֋�
���m�6�U;��Tw.�Qg0os�Ψ�ǵ��\Gu6WIq���U7�{m7����O4kITV�p�t{�h/>}�bߗy���>�z��<�.=�i�J���Y����).�@��y5�T%�v�����:��V(�Q�l H`���bGx�,OO(E%�	���ɖ8����B*����C׼�Ro�#h�ڻ�
t��(�l���sva�QSe���+da|�Ѫ�FB+
���ͧ���X�a� �I��s�u�)8���G��VT�S�����ه��}w�~��7<[�0y;n���hlO#�������l]��}�̿yu*yA��s����Y��u�Y��T,�������ϯ����W*ܡ�����ij��s�v���O���*��<���%1���d��{ʟ-�����+��5�<����Sˇ����\�th��8;�����N�r큃y���tu且�W5kL+z��ㇻ���<�cv:�vި���;f�W��в��)p���/�]8��X����b�S�F&�O*�=W��kqg�t�7(��0�}9a�	�p菕J�j+4HϹ�>���7��TCͻ�u�q���b&"�0�5�aep�s��n;���N��>�'3No���j|��*��s.�*��Y�
Y*DuS��xm[�w�+�z�Z�=�9���W?F����C����_@u�]���G��.��9֣r,�f��AU���v�����/5;�Fh�tY{Q+��"5Տ���ȷ7q��ɂ���1-��h���5���^t'��|�����������x��ݶ�>�%c	 4���!�{�[����0i�z[���{�{��2�����w;�|�|��O��u3�;����ޠ��6������T&�B�)95��]�ԗ:�y���]Q}�y���,���܈�"(Ek�W�'������Gaޡ��s�wX�|]��~>]��w���sg��)�������=�x���ع�ΧB��3��B�pzZ��8k�|{������<����6�\L+x�g��>���{�j�ܭ�<Tޣٓ�2�&_�.lz#��E�U�1./7��_5���}��]�S���}�;Ս�"ϴ���t�,�n����*�/���[z�ۈz�nC���R�r1��l�P� ���twT-�U��D�3�TY䯶�ի�Ҟ:V�35M¤�֗K鷛��S��q�|����*;+�P~��~��a\���Z�J����.�.-rv�J���Ƴ��w���HWuJ�`�P�׉��n�%m7�ڵi��g(u�A(�Z.o�4�`9�
c�C���{ã��"�[�I��K���h�m��"�ZI^�.kֲ5�͛uy��� ɜAh��4�"�)�QP���kk;����&�N�Am��Wa��ڒyz�RT������5�"[ӻ�t�f�kT1ͺ5.��2�Pc�Cr�����K��K��ܣsˁv�YQ��Ħ�,P�a&f�Id��r��%^�W2����b�rl5�����1	��؞�]��<ju�7��|LmNS�x���XXF��8"Vw{\�5	��0̿��f�ۃ_�]s@ )$GF���3.��CB)�Y�U�C֨�Vך���K����b�R�X����6�F���c�����{��9�7��4�p�rum���RPb���4á��+���m�XW�Q�`�`�կV�RLά� �z}�;�Gz�N��lpQ{H��aʌ͝Y��	#�!�%��B�ΰ��֜��n��5/�+�4�7چ�� 8(Γ9��F���ݳǾTd7�t�I��}8�`ѻe�e�ɻi���5��M�{5��=TFK�y}��tXbK�5�S�v���:��r�ە%��x�ا�eK�6��iv��H�b���r���x��{��:0�N^ �����i#!%����fޭ����S��Khfh�˕�����9����tC����H���������[��ʿX�b���[l�$4��(���}owp�<����(\~	�W� [cΠޞ�iS�GY��
��}��oBV��N����w���w�me�o�	��v��`�l '`<�ef�|��M��>w�p�l��p�o�{��H��N,�iSkl����tq>JNF+�-Y����D�wn�f���o4)]}��8Fa��a��w��<xg�>�ۺ�pE�j���0C�6at0�Ĩ�o�Z�<y��\�%��_�f�!�I{�۾�K������.���Zv�=��K��O!��z9��u��Ft�m�x�Í�{��h��y�Wt�݃�D)�R<��m�:�gs��Ҕi�Y2�=�is5g��J���HX���q8��O=����u�=en����0}�!�{R��3,�'���V1�+=ذ����
���^`]�]Ļot���clT�|uQ�@%�r5e�y���l����Hn��ٗ�^�æu���؇��;T�f0Sl^�݀R�8�y��x�,�B�q�u�]�5<k(v#�R����� �������Ѭ�Y�c���J$h�x@X��r�^�ԡQw�B'Evf���F�r���n����Z,�x���Rp݆,f{!>��ʳ��*L0���L�ɤ�âx;ѷGh/b
i�9�+�හ�F��{әі~�x(&��ֵ�W)��s=ނ����҇v�N�	w`J�z��^f8����v92�8��+�u�xX����`n4U��]yJ�,sY��o   �_*���²E{Nw+dS"
ʞ#�J!U[*�ʮQ�*jz'��e�M��+�qr#�!3D4hF�U�#�\x�S�Z$��ZM*+0¥�D�t�P�D��dY&�j��4�,��h�T�:�A6����P���I6U�����D�V$�m!3.�����x9JJ�jw\���RN��f�0�D+�T|u̡�hW
�sg�w3���y%�e��c��aX�e"�Q�i��d\+�hr�t�J2�9���r*w9��W����9�:!{�]��ȍ�Q[�x˥�b䜯���*��ӓ�*�I-*:qn`^�p��b��䮎I��ETr�4���"�E�����b�g�rrNo�wn�o �
��> (�@� ѼG�YǙt��vF�e�VN+^RoJW\tÊYHh���K`Բ����
�*����Ý��xEz���6�"�_����9��M*�q�c��+�Asl�����o��ӻ�[ܙ����羶�5{��M.�Ek��_c�V�e)G��K��f��?��OT �W�$�f����{^X]�	�G.��U5�snXR�^:��qY�������=�B�����6�gs�èO��vyǢ�c؜��������q1��e�ٵ��M<3��j�'|fp�3�]��GPk8)��5Q�T5�۠�	��I}��T�j���Vn�^�}1���mk�o^턵�v�����S�
ſ�+��T~+��K��z[��sSO�Z��y�sf�F4�8;���;ZMv�:��|M5�՗k�|3yO{u�U�?m�~��eF�ڊO��ϯ�]	��C0�3�OHn�x��%��ۃםq<r�.�竨��f���~�^l@f{]�$ϛf���s��m5 s���޻�Y�o���;X{Y�C�}���y�i ����y!��et�r=��be�	�d���y�����]�&��n����,r.6��jNX�C�كs����S�狵(
P ��n�mf��lU:���p�z��J�S�y^����g�����7cO<��Ug[�UUa�iକ��E���n9�"�3R�ujy�+}���[��܉P~�֪�,�����g�B����v�u��W���4�T;{Jk����Y��u��PD���[�[�v������n��c�W�CAn�յ��Av�E��i0g2X�WWu���wi�`Y����F�L���mO{��Tl�8�n��&X������cu.������rܙS�U_O�}�@�WzM��hT��q5B9�g7����j$s��n0�����0���,'<����hQ����h�;�Ok�_��}p�y
�ؚR�5oy5��J�ˀ�a����%ڒi�w%C��+���=˦\4��-�+u Ķ
)e|im}l9D.��U��O�%}�VK��������L�j�W��%�;/�ۋ3�Q��3V++;cN��s8wCl�H�m�SJ��jo�rE�o��:���sK:M�2�tƙַ�[U��+��2:��.ܑt�r�ލh�y�w���-$da�Y��ge;�|Z�yP:h���<�竢��G�\�/�{Ъ#Qw	��z�"PS\p�t����Dbg�W�TE�*��{�A������\V44۫�/7sM�1T�>����I��}vΏE�Aq�>|P)w����*6���v���۶���@.�.!�w�����}^�m��v�8��ƺ��V�J�Z�*A���n��Q�^�.m{�{�g��>�V��lO#��	t�������;u�Ih�/:�y�ؘw��W�{���y>(�v�m�"���wS���^w^�ͨ�N4o=�{���;z���xT�5j�[��RS|��e�lo��c���܄����3��5͚����a"Sǀ�y_��R#�W)ԥ���Pe.|�_ы��h>��3�p��ܛ���+lE*q��[�Au���CՃ�;���F�N�oU����n���c�#�{�H��A�+emnu��F5*�nN�c�3r8�L�;�˛B��E��P����;ĺ��~��U<����>[�,�)��H� W��.���!���n3�v21�]8��i��N�{w��I	��ˁUv���E�ˍ�\�����)�4ܱ��+�j�r��	�̠�Bg2g5�r�ɗK8�4��O��Z��w����n�E)F*���,W��CYq�9]�"Ua�"�r�,�R���=<k�7Ư�x\��sJ)K<5���Hr��٭\�k6�����5�7�q�egPU�r���=P��r�����$f��{@q����G�1��{5�c�}�0x�(-��9��Z��Q����:��ܣ;��W{W�N��D���S+��q
dN��[�c�_3�Ȭ�n�:d ��9��e��p�Q��g�i:X���vrrn�9���q�\J/[�k�\�d}��h�@�>YyM4��Eh@a{0g���;\􈝳Mv�V��Y"�cń�a�E5�s�Sf�z�(�c��`;���(����@S��=����uy-�dNG�U�4�K��I�CC��nڗY�) ��8���q�־Mv)K���$�J���`�f��7�B���lv	Y�YJ/V �E���og��`�[�V�  ����fv��������͠6E��;��4���g#����Q��n�4�W�K/ou�Xp.Ѿ��
_cȣ�����U�ĕTk���Y�/1��>�Na=qU	���l3)筲zCeg*X/�w�2�%�uE_���^��ܩk�(,�ڲ�C>�!(u�b���a���`LWz��+�\Cb�M�e[D�P���n���+Ί�w�t�!!�|����t��=�����z��pe �n�b��|���	��{k]�Y��iw�}b����(�Se��V���h�G��t*�][/>�A�+��u,ON:S����Dʻ�����@[;�l�*���U��l�w�Rg|F���7Z*=�����&��m�=��,��9ץ���&D��lXQ�]��}��x��C��gGE�æ��`��(I��j-��NB�ݛotr��h�6١���5N����(��l�Χ�Ӻ�-�B¹�Ɩ�R�ԥ����3�gNTn�h���"���3p.%E4x���&&{$ȯ�f[�u��O)ޓ>6s+�����{��3�������}5�~Tĥb� �����)���~�f#�R0��4>y4&w���]�Gҏ�����^�E�����V�o!�\�O�lT!��Z[���m:���K�b��K�WCϗ]G�Y|i�K��*,��U-6��[c>m���,c��l���廭v�L_��\=t[O6�a��3��
�r�;n�1���"�[���F����TJ�w�vb��P���Y�q��J����`�ݍ�L�����K�4c��UM՝25x��0,F����:s��^���w����ɺ�
Ve���ǵ��+J�����Kj6�����W{!��ȦXf�i�4i�`��1�h�t��s�[y�\�ú6�k�e���s��3�<���KU� ?l�%}U����9�Mg��|wwytuy�]��Zz+��aՑUFV�<��do�j�'���4���f�T�v'�wY]��t+��C��	A=�,�}3�M�CՊ��L���dUe�{|s=�=��'�T�]��r��Xl0�bB���ǶZ^u�>�)ٛ��`L_z��]�}7^���+��:�0�b5tQ/��:Q��{���*k�3VQG����Hnܡԩq���;��˫3�m<�@�7�,��7�f9�SbU���B�^�m��~IK஥,��d��F��.#�]��.I��*G�T���q>�D���u0�ݾ�Ͻ�L_���ٮ���?Q��̢͈rE�."W;���w�M�l��U�2��z۪Tb��Rß��l�JN��^�����}(�3���ݶ7-ۈb�4:��� g������z-Ad�6^B���B�/*�=XV, ���]k��w���m�@]krV&C <��؛w��H�L���v��ȸh�ΙR�����yJ�\�	�D�n��F�ZuB�6d�>�O*
�Q[�J
A+[�{��CV��:��R�7�7�;����y��d�h&��܄�"��>*d�b�ofw#p���=n��O�޽ <��n��t<Z9�9��=AU=�Z�d&9k�Nr�B`�Ԅ��ɞ�pP7�r��]Qn��Q0���')���&k�A{z�:�}�e����dV��{c1+7\��[�)xȯp�R��R �] ���*:u�}��5b|��R:ja��a�FK&��qg�Kf��]�5y.���e�.V̀�����H���r���j �$2-4nT�$��k2�Sb�q�y��v�'�6�UB=��9/a*��4����T��tOT���0�` ���� W��K��ϰ�c�\ ��W�^�/��=�`z߯]���`BYyR��H���e�F�h��@#��\�m���m�ƀz��ʑŖc�.���zy�9J�W7���p����6ͨ�h�n��W�[���MĊچ�֕�U�*��bCW�Cꊌ�to9ZqH�!�+��I_Se�44qp��!	�����4Ln��@^�lH�I��0΃�(8-�Dٳ�f_S�X�Ꙙ�ǔ���j����z��q�,�a�|�n�٘37W]�qAQ�5j���Y�x�.SN\w���]I��(�}���S��5�V�eo��XǞ�y�}����W���z*�	���b�&w��2gȼ�wa��$�-�\0�BBY*���,��F@/��ȫ^�{�dw��^��H��m7L
<��L�ڨ^��S��t�^��D�8
R݌����Wk�V�R�����=��~��I�P�0蓮�[��4cP�a�F���H��~�%��#%&��%��!n������>=2�)��3t8ig�J��G�������^�;-λӑP���j���$��	�si���V贡�o)��Ү�w�d���!߸;>p��ٗ�b�6k���4ok6��ҹ��?g#xVd5�vRAЬF�R��6/�2��̹x��f�6wӫD�e��{�>u��ԧ��Xr���C�#eChFuD[B�g�d��Z�(4<�º��n��ˌW M	����p�c��2���=�٠9�ܢP�e҄�U�w��exqX���ؑ� /�n�
�oX�-���EKvS\��F@�1B����G*��Q��ev6��Ԁ^�>��@4=2/Ǡ�G�%ٖ;o�3O�SY2�f��8�ܖ�OUpq�4	�Ec|�u�ż^�D�q9��%�MeLۗ��nZ�`�""����}-^e��/�%3{K{SrDu��( �$�s^|���X��-��Lr{8��F3�	�l��R��X�6d�s+S�e�f8�2h<��_�ݘ��-���7*���t����f[�?]��Q��%�L���mָ+=�H���2�ա���M��l���V��%Y��6|Ȍt�[n����C@\嗔�IV�2�(�=���$];r����aS͈�S\s��ʊ��w���[<�\�ю��̯e�����B�ialsЏk�ud&�l���B{ ��w:�*��[^�!�i�s�{B����p��.�o�}0��ay���[���9���T?�t��L�7�>	�ǩَ�~�qcd�HD�~Ky���k��g=����n��ͤC����a)��nw�R�Z�o���#m���`Xc@)�D?,R��'��x�_z�
�_�}
r�=��P��(�tX�7p9�qF*=4uj�z�x�>�wd��SC����ez�*�`�*;3)�I�b�qy�@l� -Of�跾ٯz�����j�
��h�8\c��}���y��I������zUu7[!s����p��D�;�s:μ�v�������a�^6�g�[T����=�\�������5�le�{{쿽նa��VT��e!��S	Ts�e�R�v�կ�z\�Z�St�B��:���ܲb�z��p��`��2���)Ө�IT/�>�@-� H`Ch����s�����	U^�2oO��O+�~�z���n6\e�[ea�.��3��O,��\`�*x�QO��r ���@�=P�$|1ם���#ދ�������V�^�o��@����&�x����ñ~O�h�1�e�<7X�R+hb
�*J�s����C��U��΀�6 ]�e�V��(�M��EX��W��9��.{5��g���W�v^�%U���
lT�ʵI������.�Ό�+�t�Q)�@�����h�Pm�eX�\tΞ0���k�0���b9����vt@P��sH��̲�~�o��,�;m�o�W��qó�$�U� ��}�v9z༐PN"��ٷh�s�K�#�뛇�ׂ����Qv�i��
ڷ�$5��
�5�2�ur�s�b�=��k*�������������+���?0�|�/���+E�ފ�9��aՑUemC��u�� k����UP���UR�Sņ�u�z@M�'��nUϴ��.�Cl�s�&xa鿨���w��
�l�m3��m�\ի�*z�ږx�	�k���2��7
�l���K�2�}�@/m����U?s��э;˖��JM'�������4RZʒ��:�s:>�Ozk(�2���pV���*f�
\��\�9�a��i�[�ٵ�� ����{�
�"�#���1r�,�}�\�̞2���V� �WR���QN��[��u*w:!6����"�9�I\ZK|���HӴ��p1_r8��#�'��ֱo�6D�f�]�V�u�g&;��rn}����x�$�ח\�����CyW�8�,���䶟m��Շ�%�N2�/u����������D$ؖ*6�hۼ��$�*�L��Z�6�Jށ� '2v25d�1{��z���.L��
߲��Xz�-�s�t�w]��:�V6�p,��.�k��76�P�7�t�@:d��8�����m;Ȋw�]��UE��=�E���n�
-����;6��)0�8�5ӝ��a���>�䣢�׽���?^��h:m�j�����c�ב`����'H��%ȷhn�mc���8y��޴���v<]|R��i���ҳ�&��:��SS��r8v�RSoe�(��+;�w%�صY�x��q�L!�y���WɮG�ڙ*&�oN׸���3�������x�%����9p���F�s����sfd�1�j�ŁUW

�}�sT�+%��	ڙ|Vb�h��Oi��/y�ML\G��ŶK6�\3e=/1�3(6 R���.�۠`��үc㗏L"�kKg�ov�[f�uT�ۻ�/�h� ��Ѽ�f�t���� �E����r {wݯ ��,�K � �AA��7�A�yJ�I�����T�nl/V4/��Zr��9�	�u����"=`�qm�.編���_wv!0��jڔ̌d�X�����h�h]g>:^�^�Ki[	��)P��R�g������^�۬
�6��K��c�F
ʺt��ɚ��<%�[�+�)$>� �cmmE������:�9q�S<#��5�]%�kyY�}hy�N���;s�u͇V�@�Y__L����y��.���)�gS<x�Ǩ!�{�b4��% ��SM�������LtҪ�^R�IB�Χ[���;lscz�06tU\5]^���+�9n.����r��+Q�اzn��-�r�M^ �B+�'Q��Lw�np����S5uu��^������1����Z7�yWwK(a��a*T�������|{Ậ���c�Q�u��Ֆ�t��rH���km���
���=�**|�.�sK	Ʒ+^��\{Ʊ��h�)4�osHհ�8�0�XC���0:S��q<�nnּ<L&{��N���?T{Bγ�l�vDH���g%tjZ/����xM/�06�^_m>�� �E,���q�{��C�) 6�
�=G%�� �G6���\(����SC���u�[�A�ta"� P�T�(ՙ�҅TNURIT�D�eUh)�l�9@meb$�}��wB?:�Or4�͚�:d2Z�(L�(���0��0�]��hI	Ъ̪.uMKR���#�oGCZ�x�tȭC:_�>/W�KUL�5(�T��������%����(�ҊLD�Ґ�5��@�(��H�A"�@�O�NGUV&'R��qO�:�!9d{�Uy�h�U*K^�
"!D3�UU��"ZV�*�0�Q�&)Rs����r=Bְ�T�Z*��M#wK�f�̔�!\*L���W5l��
�J&r��D���-K�F��\���
ֹ,�6�EG�vm��WN��3��DȪ"��諩�N�ZF�M2�+�X��QM$ ̳���'�.�r���("�L�f*
Њ�S$��.9%EL�*Р����
�8�v�]�Щ�Ư$�:�
n���bl��˺=Y	�^n��έ�w�#$�m���l�n��O�~�N�;�UZ���w�/���S�T��s�㋯i��~)_�1�/.5�G�5��{���\��JK�+.���|*f��c�<�v����E)���Sl�J�Rʵ<q5�n�>-K��nGU��(����J�D�${�[(�¼^�m0���!c"�1���ke�\!��!F�wwmq��Kv�۞��x�=[5��*��+԰�Ĵ}�P�|��4
�U�4�����or��5�[�X^-Y	�L�lU;���]P�B}�G��{7JhW��{GĴwe�Z��Le�YrA٤Sn��N�Eϒ�x��_�l �3�d
�L�Q�A�m�j�M5yҰ�zYu7��uk�|�Y"�8��lK6o	eImR�>���W�e�Q�*N}5P��F�cH��B&�R-t�����3i��5�y/kð2�J�ô��s�:R�N@�|Q'v��Wf�NZ���zI�}u)��{%���Uk��^y`)�?η�'�v�T�t<0��ssN�bt�=G[J��m� nYW��%a��K��הHn���(�&y��۴�:V� �u��̓}���.]�&�`W�ilċ�8�vYl��K�n��K"��n;0�2���X�59l9YO}oY<�ٯ�r�҇��r�����}]�e��Z�S���r}�&����BD��- U5u�o�c�U��th��9tޅ8���,�OgB3��jP����͸�����̗Z�`�h���A��ֲ[��fd�b9�ʈ�O��n���K܆��+�'���Lܻ�e�P�ki�	e��/\��ze�F��OdSA�{�2�7���)V5@��wZ*wn���f#]�E{�>Sn*@S#�aJ�tR�W��<[�:t6�=���e�[!�G!��ұ�p���ё.��B��lrGz��)^�rۑ��d�s*�^,���i��':� |��>���W7�=3\A�W�u�gU?_�$߹t�{}��=���{��I���P� �¯BV<a\{����|T�U0&������^F�B���|XȞ���Y^�D�eb�=S�^�KbC�s���*Pc�S��/zG�Q(�5�St��¼^��P�ȔK;�dʦ7�F4�Z�11M�'�[П�}@`�z�~
r�/AʂPf⌅>h�q��\4�F%��V�������e����c��;��B���$�^iR�<K��d͘-�#�M�+w�Em���M�_YR���q��Y	j��h���H:�h�J��Z�]�ߒ\���z�|:�k�!C+v�mF)�d��lD�i(�ջxJ��i#7�Ԛ��Ƨ��3ќ�R�y�*�m�pW.�*�څ;��+��q��kge֌�}޻�7w!Em�L7��i�uӃ2ˣ�Q��g���.�:a�sy�F+n���K��&yݔ�L��^�������e�p	ш[�
4�l�Kfj�t�:fVƨ���ƵWn�
omՖ�����cѼ�Id�Ih驇�>&;�=�d	�a�[�4={yM ��d籓83vгeA��{�=	�-�+��L�-�HV���Z2�.[�5�!��d~�������X�]�U<�^�Ϩ{���o�)w���~B�$^�􁢋Ds���Y2�f�e�ܖO"V#Y�%]%����9n٘A��+��V��"�-x.�!>�M9�;U����,F���W>f�XD'YX9�n���P�7j
nGi�l
t 	[�t<ܞe�;9W;���R��4t��\I
�x�J�**�9�)�:���_Aq�JwE{��<���36_�O�����T�n��h�v	z}���Tυٜ,Y9㌁��9ڧX|�) ���R��@0�ۻ������n�8v�7���F����XO]T?�WL^L�7�>	��f:�{$@�ׯ�cW;�탮�����h��r�+��U�_��(r�}B��A)٨`LWz��)�1�l_��(
۪F]
���[�+�t��WGi ��j�����M�S"{GG@4P�h�S�[�r����2l9�wN����鰻T�6�{��Z٧����JI�V�����e��٬�;voHѕ.�v]C�j�/���;���TQ�x�K8�l���b�p�W��)��e�x[�V�b����;�<ٺ,0��8�5��<[5�2�Yev��@�Z�ef�#q��=�����o�3�r7��ߪ�~ܖZ�� 6MY&�֋`!L� {�m;��I��D�d��w>�aT<W­�[f;����&�u7m��+iL�in�ڸ��J�y�J�Q+�a��x�Fς��	.wǇ�O2�G* ;�yjg���Uof��ư0λ�=~�����VLL=��D������Z���')��h�&Xތ��Ɔ]lW�3�N6۹^8�y%Xs��"�=�n��]O�R��^H/�ʲ)��y�5�#p�h�k��xW��Ϗ|_�pS`����~�������nl��=�Ih�Zޛ��-�Z�	�w�X4�ݡ,���TP�%����M� ��^�����[�ɩ�r�6�6�N�֯X�����gѲ��4G:��$��耡��A�I�V�r,t��>�yј�,��s��=��K�۝���mh��D�ߵ��f�����w�w����g�������p.�t��Β�p��k�mAЊ�ɂ����q)���y˖@O��wFs���.�#ϳ��60��Z�<���v�wݨ�:�i�>�:�ʝ�*v0i��ի0of�&,�<�����-�=�&�wt�� 7���t;c��j@�O���j�׷�q�a�K�$�!�9�0����-�W+�p� g�SnղcK<2/���x�yz����#����t¾t��v���./9�٠+ne�ĵɖ������k�+�̷�}�J�xԤ�z��IZ�(fU����Z��̴��׸�3&pa鿨���w�F�:*�ޗ��^��.�*8�g���(��5��J�������J<��J�3a��V)r���:f�݈�#oJ�Y,h�d�
u���f�҈����*�`���cyƋ+k\j� lU�
�o���r�B�����u\��"�|�g6��r���q���m�"�S�2�X�4x��[xC�b9o�4�L�)�GH���\GqD�^/�
�篅�:b�{���I�\ɹv�!�7� g�;�G�B��yd77J���Q���RÐKGّ��5�uoL:��VM�a�Ģ�|h{�Ŕ��뎶R������G	eV!�C�ɔd��9�N�:%�o�����5�6��8�tO-�h�h줅�W8�m���;��Y꜑�#��S�r�bP5Lo��u�L'��tȫ[�w�7r���b��:y���_%�QZM���g�ȷ&�#���Kw*�k@�����l�Y�ָ�/;��y-�!P�Uԋ�� �~�������ٞ�]x����YF!���Y�y^�>�5DW��,H�ح��s�b�;�{�R�.o�t��pg��`+��%�y-�A�A�sB2��aܴ�u4J�O��b�3�f��k�r����kײhi嘨(c?P-�B[���ECW�.�[�3�l�32)�u��+w0�P6lhE����EK#W$��� a�."h�:�m��}�!Sl ĵ�=U��jvS��m]&�W��*��r����{^�V�+Ƒ����1��wy�I�f�z��d"k["v:�-S�ɘA�G q#T�����Z�@fg���k�_�׍'�­���;�ҏݳv�����ה���CE��VL�d��ze�F���@#���梢��t���ج�}��c	�f;*�x�w*+�>S6�20xf��E.����#u�rB˱���PaEd�eqw5Vc:B��g��\I^����ލ��@߳�'�B�C0O�.�l�t�cC�4��M���0"���[EŸȖ�aFL�7�L��O;��x�_?:�=�^�)IsA�Y�z���2�=Ĥz��U���^�,���ES$R*v*�y2�)��ژ^����S�y�7
��9V�_��&��t�"��:��s5�ލ��*JF�$�r�����;�"S��7�[�u��eՒ�甹�������VEa����/V�T[�{#���Z��xy�7����Ɯ;;.�[Xg�M��Ҹ�Lz�{�#�y�T�#Mlnv����)�3���N��]V����K��ޠ5;����w��P���(�P�LE7H��¼^�9�W�*�~�峼ZiNsRm�p䶦u����[�r�����R����͓�=��#ڱ>˕���`I��oپ�s*\&m��̲�-׻M5ҫt[%�x��)WT:Q�֙���e�P ����z�ű�g}[T+��̈�i��~5���D�ζ��d7 А{J�;�:��S�Q6e槬+m��0�_4r~hhn3[A�z1�i���5V��S;J�#:��!-�Ö��=�}�Cr�k���l*/�NJ'"&�����C���11MVѸ�>��Y��&��q�#�w��T�.�wZ
�0l<Hk��UL�,���qq2�e�\���!��d~��]��y���Q�zY�-��Y����T3�;F��(�,vi��7&�"��㗹SbUfI�켹Q�6�"L�!-�2�2!7w>#>�L$s�{��m�8j<��Q	�$).'���,�{M<i��
�Sn�}��&)���)�s�{n���m�A��!R�Y#@�fhg|��<g���~���gI�)�NVt�NCw�2���S'����^�Š�]$`�-��N��wdoC@����{:s��,�71l'��V����A ���� /��L���n#��Y��3z��hrWn��FT졮��s�N�,Be<��e*��4Z6�i�9�/6���.Z�d����cn"v�ˌ�Ү2X�:��Oeu0;!'�,�ܰz�~glI����[$D�C[�a�R�����o@uCw&y�Z�H�5�{�ɇG�r�$I��Q�^���2՜�m ��}s�}�hvym�a�	l�`jڇ�Q��'Y�ɟ��P~qE��3��w�ݍ���J���Uw�����|�=&�Sq5	��\9�);��]��zoi�7찼��E4��ٰt�-���^��оuj��S�Y���
ve �n~�\~n�����d_���k��w/X��	���+����)HC�P�P�b*GlG(��r#!�b뜬�;)ߴ"���T���y��3�e�Q�o���6��ܳ5�ކS�Џ�u팽�`l�Z����|'ةp0t���N��׆�p���M��e�d�ǹNjJ�(ع�����ݛ���� j�U?9f�~|�0��"bb�W�����Ǟ�*�2��U����KG����p�)�=���{2�u�p.%Pjx��𘘧մZ�nr��{�o�W�w�L��[ݕz�\.5�j�e�FӮ*�ʎ�ŝ5�!��suy���SǞbU��]�:��*
��y+@w/����5�"�U˔�k���R�>xw
�txA2�u+(�ya����+�pq�Ǳui=R,�xc`�O)�A0[.�X�w�J��i+�B}�a����,�D&�fv�U�V(��{&}#�c`�'۴%��UE
d�]֋�tͺ�?\�%t ;n70Z���!T�}�DM�vd�U�B'�9Ȉ��Kf��u�uPPֹ��C)/���Y��l��ce�;������E����O�����������{�m+d��8��S�d&��p���U���)�%��Ȱ˵�0�f��h2�ur�s�Y�"�C�U�w��I�R�|*�d��|�av�;wi�>o/_UF�>#�%���p���ɖ���Q�U�!���Qwי��a`-�ʤ!��߉���=�ւ�<�8dyh�.�x�zv(��
�Q�V_���&�S<�Ţ
��g�D5[U�,�k�e�qS�w���:��}@S��L	Գ�fO$��^�W�L��}p�2e(j����M<�Υ���;���[5�ۍ����ڪ��޿c��\��^��H�J�̰2"��s�[9Rǻޤ=���b�Z��W�/D���czj��iԺ؅*��d��گxJ^|�tޏ�)��]�9�<���Us`i�0���|Sv��Hn��w�oդ���ohj>i���!M�mcފn	Ծ����kWTJ�Lr��Z���-�����rDy�J��J�wU���ξ�JG�Ͼu}q�r�1��)ٸ*@[2G�&[(��+�wK	F��!CL:ݣ��VJk���u�΍&"�[{P�iJ�Nr/�2�"�(g�S0���8`;B�]7^��U�O�r�D�Jl�Z�B�ĿRG#��@��X*/��@����zdy� sɔdJh���ϫߩw��m�]���g��;�a3ɥq7��r<��.=8 ~�!DS�rE�P��6^%C(/�T��n�VtdVie��d<4�a�oE��'٨K*�[T����K�_��=�63�l]���������TL�C-��ڀ�F؇��P�"8mƫ�eLw��WN,��qLF�Ƴ.��6�:�z^}�w���ah��T�m���^���2���}ʬ�%HN0�i��l]�/�u�AL�K�Er�r��������+�;�A��MrHn�2�Sb�q���OP��f�¨��Z��ת���?�5r5OO�o��-x]f~�gא?/�k�r+��Lr�g�$+���
4[��)��n�;�f��4.�j�ʗJ�-�\�'�!��]��u����H��x�tc��1]�e �Du�;�A�����gֺ*e<��sڌ_ ���]ʘ6����z��XA�o^n��b�!���g8-}ۦ��N���j��xe���1{�Ѧip���s��] @�U78��@B0m�u����Ԧybh���Rj*4�Z��y�Ӝ&�ky7F65!��\����6;ʆ�s�2�Y7d�Y������
-Mtc���
u�������}y��b�Wl����b�y�$��-f��/9nDxS��I��b+����-vD��ef�NK���:ES�-��b���*��ʔ�ه���<��h!�����6���r�T]=9����1�Z�m������y����q\lpB��Aa�'K>U!�)��ʚ:���i�5�ʾ�ˈ�BjՌZ�Pk�v(ڇ���4k��p��:�]p�Rv��D�A����铬)p�aͼR�n� �s��E�r�ъ
ͻ��N��\�c
z��3"*r\:�&�gة�i,��o,��s<8�����#��Q
8s^�X�Ε����Yyٴ�pl�rʻ�Z��}�m,�|�M��3�ʼ�s���������GQ�r�S[���ŒK[�I�P�3��D9k"�,� β�jŊ����p|�f�ə��vN�P���$������ �*����6<Y�Ux�9vX�2Y�j��D�5��Ϻ�����f�*�c-�b[��� �=m���;�=�v����>����|i��$.��&n:5��+�+C��̍�i��B�.����E<��V���ٔo�:����!H��#hҚ��r����q�;}�pqK�%łI��4��*;(�� 5 m��ɺ�p�*�ĪA��fcF�J�}܁���BŸ�!׮n%�4�@3��J�8���P%{�f����7b�zz�.��
�!�+AÈ$1�������.�6�lU��$�X�� �U��U�>�;��]�!@��at`B�z�-�vG[�]��?\�j�% (쫸�+����p��f7`���'_k�K�O緮�(��v$�s�C*�u��7ȕ[�Ck2=��}��kH�%`��v��/�z¥���/7�2��u�2D+` %�,�.em�_�um��>]B�q�v�6y �o�C��q8u	Ϣr�$���oT�F�U�5�\M��	�"�]�,�i4�*8��C�v�r�]��o���%&���:z{�.��v���=��~�cWKH���5C^YM�
�:Ιi7���p׀t5��w��.g��9=�Vm��Ftu��6JB�
&�{�p�F���G�,`�os�#S�tZV��[��5Ƥcfݢ>/�a�0�+#@(R�DUxI\�(�D��rg*�W'1�*#�AB�
/$'%��:*����J#�$˦
�
Ieru""�\/3$U�,��U�4��Qj��9�q9t٩{���G
*�z;�l#��U9ʨ���,��Ȫ�((����	�*�9��/Z�DBe��"��DI;��#�\�Ug�QG"��z�"" �9uԓ<���]=��E�g�z!G�nx �=��K��1�g*�6^N;���wD������rJ��C��瞠E8s���,��@�wRڙ�{���Js�ԩ��Q䜬ȹ�\�8@��q.�IF�UV^㲜�$�E܎Tf�%T��dG�DWwqtHۻC�Dz��y�9z]f�e���1c��^Zp��Y\GL���Լ�<!�"��/[�䪆���yUG�+X�Q�*(��D�+�	E�f)s�=B����=Jq�5*���q�$�ܥF��r��-���d�7yD��u�f��@�x�c��o���+y�N�mY��q�%ou�;�g�~�,��ꎛ��y��������*�ø�j�����mO�u���O�N�X�7h��:��Ѿ	���fM��3sF �@�N2#_(E�WT5�ފhȗG9Rq��!�+��X�vD�S���T.J�&;���2�C�y 6r''�`Y�,�g����_9��H{V��I\@�Yy���!%}M��B��L�<6�y�c4;�(�lf[U
��j�V=����Գ]�طM��E��4n�JV��~}�,{��P����[q5�tg{�����W9�\h^�l�+��i�S�(�����X+޿_�D��,��CsD��� �ge�"��Y]�9q2x>
3n��4q0ݣz�i���V�H>��i���*�J!@r�ҫί��^���6�����7�->�0y��L��
��g�NdF�񨶕��D���;�9ģ{�x���-Qo7�dDs�?D��ɉ��t��s�:3��Zwc9z���R�Lf4���@����������m��Pb�����MtJ��;AƋ��Mr�h��2��	c�͌�H�@�Wق��`���	6r�w��4~�=CO�L�f�|ٱ�N2�L"����6�d�3���S����;��o���D����5[�'��#b�+)Ik�����+��o!�[�r��-� ��WJr�34�'�~�l]W�#�I�K�fl�(w��'V�R]v�.�����M<�gS����,�w�]HV���Z2٢�׮I��jr����tJ�%�iL��͒�������f��]�����#c�IG	c�L�~57���Y���R��F51;A~ B2܄�u�'�홄���)b˶M"�-x..i��z��y�3,�ʧ$���K����G:Ȋf������p�A޼� -����f���r�<^�j���h��2�.)c�.U�����ᕞC?)Y����<�_<�k����>������v�y3��p�l�oEw�>ë*��ɭ,^L��k�5�WCݴq,�̩�Sf�����i�x�6b��A}����<�-��=�-�s	�~;����~O�]��_��y�4�iy^�á7Ym��`�YҴb�Nu�j�̋�M��.H��TMCئt�3�C�������ף?q�F�f;��u;��OK��v<�>�Ϸ��)���^G�@S^�y�jI\�w��w��-�NK=�Fꎳ��9l��
{���0YQ�J��R�����x�p�L�w��3�L}����ҳ�#ݸ(��۫Q��l�Q�3P���n�!0��d��M@ݥW:��fwGS�76��WX�v�t͠m�R��˸�K`7��v[[Po��k;Y�`B"���Ov3q�6���%Rf�zG$w{� 3ǋ���R���G�]4M��ut��ݪ�Y��6cO��Q��Ϯ�{ ԅ(Դ�wnbD0���\{>>��y1-���*O�V.W�g�>
�ڴ&�G�z!R�����g�u�zs�l[�P�����,�/>D@�m�&&)�{H�2�&[����� �^����2�ӖS�R/�)@��{נ<�]���*}!��@���j[���t����sowr�M_L�e�ݐ&���oʯ�>>t�9�䮝嫩Th!>��،�P]��5��YZW><�@~M]&��"��8�fݡ-���W6/��x�M��� 8�Ÿa��9fӛ�33I� U��/�P�ً~�hF��r"�͛wmם253,qS�6�C���p|�Қ�kV��FٯE�m�E~'�xT�3�;^��vN��k���F�*�ǃ�n$���Uw{��绻�Θ�R���O4�E����H����n�����VbH��r���
��wb�Yn�Y���6���R�� ���յ:����u��d`�̷X�0ݥ���]I�Н�2���쥚�bK�Yi�C��o�1v����X�h��v��������w�e��*?_���W-�Y��πc<�s��4�y�Ɖ�԰���+x�2:b�o���j՝r�U��s9�>af���v�n��t�[T�'���X}ʵ���޾9f�r����9��2#�\�ú��&`J��:_��ۨ�y�2�\Aئ����FL��U�[,�Cp��l�Z��m�ы0C���ɇ��� ��w�+���f�]Rw�ΦUq��� �K�3`ޥ����p�r��%�7pU,�+��St��tU��)��z@[2�ʞDTEϑl�Ա��;޴<��8-�c�b�ЍE��@J�ǈl�i�WX^ݎ�M�J�^�����GQEHfH�D�eq�x�ͦ��F�q�$����]ym
[�����4W���*d��hSu����v|Q�/y^{��Fd�d�\�g{J00��l�W[�^�9N�J�\w1T�^Z�uC�R�7[�(}�3�!�魛'2՞�L8�ض4o��m��h���
�Y~� {jlm��$l[�e���:���ͭƔ�f�j�i����@�y�V�ʙd�â�P�;��Z�f�o�=�n����G:D��h�DNSq��=ei���wǰ2��pӟML'�k4����ٵ�fM^@�7"�S[/�8({H�d�d�ב|vy�y�w�YǼ��Xlk���ݠ��FP�b�'Ρ.�˝�E`�Mg�A|��+T�w�݇�a�B3Ћ �*����],��md::EU�+2���������u�f�^��9�K�Sʺ�z���.}��V���@��ωZr�|�dM�=���.�S�	=��I�M�4�P�w�gG^3¸�캦�.�=�$�l��!���x����-ʽrHn��+RF"������24�$ҧ��q���ԩ=���Tp+�y~e��3-x.��h2�ch��/T�s���iښ+LMg",�4�zzXV�<%z��'a��q�Ӏ��y.��`*S:�Mq�*��#ٙ���f��{��4��ٌ�	ܨ��l&|��N����䩷E2��i�������kN]��g�X�x�u��.-�T�ub��T5ft�tc�W��8L�+��UP���c3K�=k��|}������Q�Kdٰ{b��1s�,^L�8O�k��v]��eE`Ɏ2V��{G�Z��Y��V�*�`���ci6�h��DG8u<��hV'�=��z���w*���h����q�QtϺ-Z�|�יU*n�P�b|;�ך%����g[d�N����2���Ӿ>h8���=k)��=�يhX0�w��J�'�P8v�������������[�W���ߦ~T��O�%i��Q��(J�^v�m�:�j���j��&��h�
�1��I��.�+�1�[L.�b2�g|�.�6T�eP�����y\�`M�z�KԷ�J<^�N��E6�G�˻�e+��e�˿��{>������@�O����4i�W�z����Y�x�V�1�e�9u#��O�ln��Q��/�i���)��UB������Ӛ_��i\I}^�P}9Ģy��Y�:��9-Y�m�"�	�Q���I��|�ɉ��H��=� �V������C�x�/)�ڶ|U�w*��͘�줢
�.�^[L(�����n=r�hi� �NIy��ʗ>�/Lh��m��{�Ԧ���]d��S8�<��Yh�n4�$��Og�ùf�jU��~�>��uq�hp�BX�j�|n<Ի���NP!A麠h�hR�s�bqk����\N�\�B��r�+`�7 {��=��fzf*y�
o$j�`yGd2q⬬7�g�����G��J
���J�K�f�2b��YO��(�,���� h�n��P�Ï�O4��@�ހM
5�z��\IW	�=T�Ft�:�<��z���U������/��[,|�$n�qW��.<�Wq�G���$*φ�Y���=��5�I!@_�o��A�yv�\�lWS���F.�P؁ݤ�Y?#��}� �$=��>0+"��e����9e��-�L�8swB8"�۹����Vîb+�n�2.j��$q�����\gDV䳨�7p�i�G��4&۽>��-����k�<Rw�E��@����m:�=�m���2�yX0��|K��-��\=�M��9���?���+#��ȟ9��]nl�6e�����^r���gJх��|�t�k��H����ES7��	M��+��xW{}FZ���c\Cg
h:���t�,���Z�|zn��z��0Q���/�k27�yN���7'�x	��\�9z��e���xn���`�аa��/�܈�	�	ر��Gv��{�{��>�� 6l��z��D�Kgs��\)�RF78�=	�C����Į�4�K�Lې�Mu*n��IcL�0P{U*5�� �^9�l�/r؞���s��x�;�]e��j��ǌ�:5�Q���{��LZ������@k��D=��:��XNadb;�'��q3<c��М-�CX+�p����fA�ƠlD���d�M<�F2/L����+2d��rEx����
�O)��B�t��W�u��y];�u*�2�Õ)K;-�QS��{ٻP���o�j̇��0�R)�q�B[�TČd�]֋h�u�wm��6�1CEN�M�kx���+��7s[�m�@i΢��&�6sG�$�:��f/KQЛ��W��]�z��{u���z�@W|3����C���C�D�`ހo=��mql]4���ﶢ�{���*h���{F�Ĭ�,v�D��m�mhw�N�c�����[6�ۯ۽T7ȹ��׎-&Z�9�Z�l��CB��'�@��_�.O��Z��c���I�wKim�܅P��՜����Q���\��rJ�{Ξ��<�F�^e��S@ZA�릹X9��I-ۧ@H4D9����`5�4�{7��O�/��~>�v�=�#����,c@V7b��V�Y��ٛ��Ko��nʡLzʮڗO�ۊ�̌�����yu־=�-/:�nL���@D���^��w�j}tmc���
�k	�xTd�]1�U�b�C�a��6�=i�9��=�U�Z���i��C���@R���@��0'��\;ɔ�.2g��y�������_�DjO��8	��e�TZ�<�᳭.���Lm�,��uL�J��U0(�#>��-��Ǘ{և�sƹU����'V����a�q�yO�ܯTz�U9e�N�����T�KDw�ơ�I�n^�Q�I�|MZk^���W>&Aҥ�ϒ�l�b�
�zd77�=��H�����>��vSr:���n���`nˉ����vE��΄�}�����Ed����yMwp4�CzJ�F��,v���է�]���W:��'�;��$H֠U����ׯ�/̝�G,��{;�ǽ��	$�����i�_V*�H�̵Jj�3��.����%2�uG�\�zh�;��3�:�V��*/j��k뢅nT��۾�k ?Y���M&%����t�E�����M�줃��q��Qw~�Z����F�h0�Mu� M�S�ޘY�=>��D�����1N0�l�$[0b|�5
el�e��@i��??(�N<��s�}���nϿ��h���1��#����"�����-�-ܭD;�Wm���c8��7{3e�Ŵ(�u^~�w�Ѐ�-�ah�0�f����OAq��yY)՚��I�=�5Ւ������r�y��,�<�*��c+����L3��E��Ѳo�)%�.Q�<�i�%+��g��T���}L���S��./%�k��u��mm����E*�K�K���P�3j�ޗ��q��s����ˮ�0*ȇ)k�~o61�� ��"�G1��}�b}��Q�������������m��Gq|�d��녕�Lkn��4�rM�h�㓓���!�3��9鎈�!9<d{9��
·;��f�Uh�Z��Q���$���v��=�r�̗��H<��V�iR�~������)�ʞ���LЭƻ��������B���{a�e����N��;�3���t�b��*�J�t��)(��8�yup]z�l�	����(�
�I�GM$x��E��wOK�q���Z���%��NN�,���b�&u�'ȵ#c��8m�}G.�·�ׁ*�s#4^]��s�+j�ƿe�lL��M��e��<���x3��M�U�Z���
��e�VD���T^�h��'=8����M��4��5�O�j���n�/�V78�hgUy.�ApJ��v�<V�"��,��|��.���Js싑�V9
ZX�W;,Ȅov<�+����훊2:�}�@�FKGۛPѨx��\:��}��\F�'G�TOUs	�|�NƨM"�ʰ�c�҇u��@*bdȁ��Ҫ�s�sai�/�[J�mSY�9��@����G��ʶ��q�;��DM:�$��yD��ںD�S��.�m������e��lB�q�Edn��c�ɜ���Ψ�hQl�L��	j�޽��-���\�==�drt���s[uZ�"�,��{)	NJ�>r�CG)z��9�=]�|i�q5^Ed�Cւ!o1'���]ZX��r�L��G:ri���Jr����Lݳ0�%���L��l:�C�灢�y�oKK��ݙW.�Cv��<��b
��^Ю����5ݔ�tL"�(jrgj�p�u�-��Ҭ.��wZ����JҮn�,W$/�s��%�m�"Ӄpk���=�>QvR��`,�{ϻ)�<���nJ�4�v%��>��j���Շ��[�㠡4����M#��ѣ�&5ܭ�^<���q���W��0���N>���D"��Aܵ�
,]U4O,�^�:8F٣�s����'��skm.��oQi;�Kڋ�pm��B<h�T�t
�ׅ�jWe^�dg��F�.yݮ%N�5����s�-�������Q&�����2�U���6H�tƟ;9���ԑQg�U�Pϕ�����̟,$\���{�W{`��:`��oe!�:��"�ׯ�8Y�.n��n��/����5�nݜ���Fm`b�����Ru����ɼ�����}���hj�٫Åeo����5Wu���D� }�z��@>�i;����H],�:�g}v��H�ɕ�V涄|���ѓ��iX��jg!����W�k�:/	1�u�nd�o�{���4�^�?����7_[ǯ�\�0Q�B�n�j'9��kz5�}�c/�>G��������:S.�Rs`��1�.Ź�#˭�|�d���p��A����:��2�58K�ȵf:>��'t%b���\j?c��`�9�9r�6��1˪����E�oxs�9�
PX�s�8/Q�Y�WjAb�n��[�n�
㬎Pf���Jv7j�:�%��<PT,/�m4X�l��x���B!�%�3�{t�fk�`�OZ���r�h+�*�!�7)cb*3m���%
��ti�i_{�.#	�"���6Y�S�N������Ҳ�0�K�Z\*�'�h誛�͔^��:��St^b��ఇ���7L� ��흱��l�*�i@dB�ʊ�a�9�c
�&u;�T�p�;��e�DK�ze�3G��~���[����p�se#�I��v��+��GJ\��Yښ��W�!k�=�T�uݖ���,[�l=N��d���qX�0[yI�`����W�S�(B*Ѭ|t���;R����<XVY�,;�^[��+z'�����1l��:M�i:���}S�oy�J�=�v�f^�J�۷i�����sgU�����U����t�_f�֜A�9<t������P�ޞ��0���E��񩄗̩�խ���6�>я���ȸ�&B"j�Jn��Y�S�X����y!����":���D�Ŧ����N���Q��]��J�'����aAv-�ts�o�R�QK\-��k����z���]�2;dcw;���vg	��V�1ou�_�in[K[�s�9��bt{�XFK�$d�s-��^ �����2����S�27<�
N�\o��%��&�x��=�=��	���"'�/M��0����]hSE*۫ޏ�c/{D}%Z��z?�{�C��su�':*y%�wWP�*'=Gu
gs�WE���"���Bʣ��9!9�I�@�"$�OQԼ��c��x�����{�/+�-T=/M4ҫ̇	�w�����43�jAz�`�֓����{��Vt"�C�T��GB�r�Vaj�N�z�J!:��㻷-p����Q E�ÕG�/r��s�����4����Z�r��WGO
+�䬈N��NN��B�4A5u�=�v��(y�"':�hNz�9֩S]�f7v��.�N����/-a�����azYTym"�������ܽ	:�+��E.��9�xf�Juq��p�0��iGgsM�v��p����!9:�)4V9�#��wӪ�vQh�^wP)��<�QD�'p�W%B�����<˔^�n�wVPX��U������=�q�:E9�)�R�sn�/[���R9��Z��wtA�WW&�IҴ �ّ#-Q씮���^WY��㛈�.G��2Uŕ֙J]�����z��؞�D��_J|wܥ��P��5��3&U-�ŉ+�P���Mœ-���e`��D�nC���>�@A�kބ˖]��+T&+��-��
΢�ꇾ�$��2��s��x�{9]7��t���xۥl���q}�B�v�3pU	���/����u\�t�^��F����3�]>�Y���`t3�k#{֓������SF����~]�va�>U1��ZX��g|{o�xJ�Q7�cU�N�����-�) �A�+�|J�\����7G@�"�&�Ҍ��v�ɫ���	X�!p�3:��=!���,̳�h���;�2W\��BP�{B���.]ջK���k�fɢ���n駶���j�q�TT�x:QTo�R���Mms�$z�;�*+��Q���Nc,{��n��
d��X�7p*.|��٠ѾO�"���l�eh��B�5L��MZ���l&�W�/m�s\�d"-����Md��w#e�Q�׈�C*|`^��p��ʳd簆M��w��DҮ��B�@�h��
n"�Qx�;�r�s��h���j���QwJ~��7/��V�����4a\�K�R��>n^�
�/���:�~�®c�>�^7y���c-`|�m:���w�ëq�0{Q�&����[�۸\t�+��ɪ��/bu%u�MsOV�*����B�x��.�]0B{�Y]Pp+��럫�^�ǐ�(Ǝ��Z�~�UL�w<�אh\)�`���"c��!7�e�ȥ�Q��Ԭ̩��.�c��oN�Omf�uQ�5)��=�U���5=�|׫�i����ә�;����^#xf[<7X���l�
�wZ|"��R�wz�"���Lղ����ز%S�'�T��l1��D:�)0�
F3`�'v��Sv���]֑Aj�zߍ-��4֪���1~sr ��7�O���Y��~�2�&6X�3ZX�r��pg�*�o��-�#�g\2{4�
�UL���+B�������;^�����'Ei��?���d�B����W��vc��me�:�υJ��<׹5-w�"��A��Dsѷ;��gI�zs�:�sՒ���w�Ք�я�̶�^^������ ��Z���2�.0���0�墛 &�R�M}9B�T;��ڗO�ې��0��������HlVvᨲ\�C��K˭r�l�paStXU���N�{�&ND5Y�\��dr�̮�0L���>ǎs�3�W4n��c�*.�3z�+�;Y���R��J���hC�7u�e���G����<��`η�ޑ�ܓ3jM>H3�i�U�Cض��^�Eel�A�8�B�%�V�9P�2^у�gݸ:��v��n����ä�餔���u�.@.h{䶊)�{��8�7��ҽ-.�Ui~���\����w�7J�&�"GzG�=���|�E���h�ҕF�s�,��P�ʐ4��;��uGp��u�����0X�� ��B�j��xE�:-�M����\{!��vk�vB ,�#�2�D��y���Ku�14��t����q�hL������׿%��T<a)w2��['�0�ʬ4w
`9��s0}��ȼ�7����H�A̭G �E�}�S�Hй~��}	�lU;��U�IJ�aV�r��h��L{:μ���w|7D:�ܕb�	h���~)6�%:W�>G�Q�V c-�'�a����e�י�[PwLs� ��"�'٭������"���C,Kj���i�����u%��=*O���v��E��J��U7,Y�!��i��x�|g�Tz���`4�+����ܼܺ�n�R�MÙԳ:WN���)�ahۊ��Mf��\'�u[�4��Y�&�8���,��	�\_��OM���@yd^@J�C�;P����s�3"�b�'�%*=�/��Cՠ�u]̉߀珫ONW�c��ڼcr'����DZݦ���}hF��>Lu�f������o���(aڷס@,h	�t�_P5��.�gem��O�ږ��Г�=�}���=���юǱݙO�\��ϧ:��/��zK���{3.z���3��O��zx�� ���Ԟ۶fzb���f^_���|��m��HM��]��R����m���*�*C�q��ٳ8p{�eGS L,�`\r��
�a�Ye�K�$ܺ�����lXq�M�].24e�F��Pc�����ڝ��^���@L;�E{�҅@�`��Aۙ�]�x-�ymW��Y�ۮ��e7�����V�~U3�w����ٕ�.9�0ME��aB:�=.��C0y=���w��Q�{:Kg''늦Tb�渃�$�6#c8=J�+b��J�b�ڧ�}��~]AU	f魦3k�<a{�e���|T�U0'מ�Ye��z&�oR�䃃�����r9Q{b�W���î!��d)��;#ޡ딹���p�^�*�緊�|*%�<3Nd��Cx�v��e�7=������K�JT�[���&zc��+*��s ���r�Xd?M�(�qFG�%�@�d�}�P�x�E9�w�HE3���{ 
� Z������vZ鉬�znS*Y��)���*�P\��XZs#e��[J�}��(5p��2;5W�'�\[Z��5O>�gO�-���.}���\�t�zӅ���8m܆U��s6���[&rt�nA[��=�c<�.��Jr�{�S��Yl#���I�<Z��o���`LEg���\>��,6�G`��ͧe��80����ݮ-^�hܥ�+56��ܲ��n��N�<1ri�>��5WC���;:
��V�]�!��d�gꄢ2`
���1Qn�H
����o+��5�,��p϶s���voU�>�,w`�3�H	�o)�/�K���)�w�]HV�Ϧ��󽄧Ъ�%c�V�j�ޯGR��ܯ� I�5����ވo�C�W��ϊ�Dg�� Z�iO��y�ٝ���#�\��X�tEY2�^�+6�"X�r�R��"{Q��1g�+."mh�پ�^���6u�x�,vGӱ�t�ߥ��pSβ"����M�ȼ�͌�5�\��X�0��=�F��Rƒ4\ c!F�9���H�k����#}7�1�(=r���B�� =�?Gf[<�u�=�S�+�oi�����Ը��$z�.��2�&��|�x�ZM�{��)Z�1���D�ݝ.�����H��w�WE�C���Cܤ�	��ȉ9���:�8xR���g_��Z���D������[���yʖ�Ε�+��k�O[��������%�rU��y6�J��{z��V@j?QڵXE
�@<7W&;�:wT��Y�ԑ��3&�z�w\�+�L����_R���\O
�ź�[[��E�n2�*�'�ia�:.�V�>�M\Ư:��G{;�I�ڋw��n3�2o���4�d��y^.�KP,fO�M��f8	�Q�gxU�6!Q���m�:��CxvYF�������r%X�����m��j��!o�V��=�H��	M�`M7p*�I��CG[9m2�Ч�9�w�QS�(a�[+�d��)v�cK����n=W��F�֙�eHn*�z��D�d��w#e��z��D?vZ������b[i-�v��d�O+Vȳ�t�p��(0��^iڗw�6����!����f	G��U��7��R�Bn]w���.w�k��dV雅�pvv�+ܒk'_�d�a4pڵ�4��X@f�6�:�ޝО�l��q�q�ԗ~����)�,�i��Sl�<�@=l_3��cRs��;�կ=�dS1	�r�~U~9��=�̀�F������Q���K�� ��(����O�g�d?KR�H����v
���t���2W�w�f���+R1���u��Z8���U2�t		�ْ�W�1�G:�z�C�
��c��Z���|�Լvd(jf���IL��~�+̾@��[@\A��,ź�\� kym�SYhk����{VgB�]��ꕳJrAe�
9{�{�s��y�_V�!�lK�6��mf��7Ϋ\Y��l1ՠN��Ŏ�m��s'=Dg]�t3�Tte��+6��YN}�(묌C�tk����g���ux�ջeÇ�oW9Ã{���ͳ����h�s�U3�<:)a�y������P�7Vi�t*��l���rP�>��{���`O�*�㗺���:A\ye�B��v���{OK�T�+e^I�Xؖ�2ʯ�(���R�����K�q�e:���\����+e�+�ne]�ͳ�t��B~����R���n�\AQ^k	�xTd�]U�_�G!�-����@�Cٓ5��/v7`^e����IG�{�Qw6=uL	��øȍ�jk�:��t��&���/u�j��.��{TB܄��*Ծ�����9�K�2Qf�T����DW�>E�5ddq���[�$嚘��Xʧ��ܭ~gZ)����]tҦS{�)�4�
a�� :���|ޗ�u���Z�GѼ4�O��j���.�~lM�,�w2�+d��hSu����GD{��)2��ҭ��@��I�'��6a���f�C�Sg=�@������ڹ��4�mR�ݩ��2ϡ�!9� '�(�ϋ��%����܄���4SGe$,+�q�%�Ojy�#�LE�+iS�S�.ci�A��U(�u*�`�P�D؛��T�7���:^�qo8+l�{���eE�}��8�Qw���Y�+WB5{���w9F]1���xrܖw�Q�����p����Q�8�]���kdn&a�Z������2�=.�C�[C�}[!�l���w���)�e��Fs��F�68��e�9D���@�-�}�WN�������~��sV�:��C���1ܼur߰l*�K�1��-�����j6�T��jd�]l[GE��~�w�Ѐ�&��Շk̭lz&�Z�ߦ�ͼ��;o�=�d�:P3Q���r�%�M��FD{��=��mYO����_��������@�M9��y�Sl��c����>3���J��l� �T�I���\^K�Цo���G<�`m;ݗ�o
:_�g4�e�����Mfd�b9�a���:k����r!��Gb��e��u��$&��z�N�4�cߛ����A�{���W��f��7�p��_˽`c��u
���y�?~g����?,/Tw��+��e����F4\[���F�H� �lc�����L��|�;e��~�_�ivu?c��YE���l���=uL	��9��Cl1=I�M�]�o;qʊ�jlъ��$-���Jх�\��5����6�,i���c]�bu�O���3����Rf 2��WKm�4YDv�
�"�c��A[�����E�����{K�A:�P�Ý�vZ��Kf��9o�g�*��_��O.qS��3�T��u�x!hvN�[!n1r�ы8tb�M�Z��V�,敾�GgF�p���ѓh�__K~�ژ^�������-��[U��J/N\/,�{��s����Kա���^���5
�{�DY���v�n��˝Gp��.��Х�x��o`3O��,�U��T<]ƙ͓�=��2=Rݠo%�����Jczzրg��d�κ��ޝ�OcHï�5�+��}%�2f���*�Eϑ̀XZl�C%�}L��4��\VI���{���@7;�x(�E�GZ�=��8Z14LL=�VDӞ��n����e>��,��d��W��{�J��z#eCP[:�.[�ג�`�D�}~�D�q�r'�)M�vCS�;3�[��T�zI�j�Tu��`1k�h}���.�Y��uL꩝�R�2�8NqFc]��b�S�����MrHl�k���
s%9ym��LݻU(y�=���?ݩ�dNLy��w�5�:�s��t�)�-�[�,�7e�X+�; �2܄����v��[�"f$ġ�h���e�P}���v��v@�Q�pВ��B}"��=�O��9�r����ޯ�����"V��-V�B�扝Gji��7R58V�)ܥ�ıt���fǧ�� X��0V��/2�'�w���p�-0�+8!aC��5��o�I�˅����&Pb�yVv�حN��(e�z6�v�wS���"�yY˃郇e�]�Q޳���\Է"q��v��
�4%��] �|PÒ���g�p�i�\�ٝ��������f���x�gۅj�fJwB��i�e�����0[@V�s�n0�<ȩ|}�'�
���:<�|���@�^�u�۔�H�����w��\�a�	l�и�`;>��s{�X{m�+���X�}1�[�P��k����Q	��@ڹ��m��r���S&��}��l�H-U� �/Gz�)"�Rf޸x
s��l@R�_�XL�F�ݻ�&�O&)�r÷�#x�l:��^ٮ����%�(�tXM�
���r��hοu��R~������ЫL�VB`/�"�V�4��zr�>�2f�m�H�K����X�:��"��v��u-�x;ֺ�曹WplM��8�r%��u7M��9["��='���H3����Z�>�VG��#e�Vա*]/�Qs�gF���`򣄶�`�7��K˜��b�㓵��O�a15�KNA-�c�w2%�3p]����[��?DG�G����D|��� 1������m��������1�����m�n 0 �0co������� `�6��cm�����m� `�6��cm� ��m��������m��1������{1����
�2���4�P��������>��������n}(���HR�IP�UR�IP%@� $)*�E%IJ�(����P��*T��UIB���`� �����RP���T*A�Q(��%@E!G�I�AJ�
T�IP���V��cBO3!"銒�b�Y��A**!	JJRD(RJJB��RJ����$����JAETT�R�H��%H�݁�
!@  :(Uk`La�Q�30Ui��**c PڪK X� ,UB�j̪�H*�#Z��(%�  :�U ���B��a@*�5:�EQKp�袔QE(��[� QE�;�l�Q@��E�6�R�(��[��P(��QE;���(��irJ�SC
��I�  b�P.�h��kkiR(�ͲPŀ�B�c (6(V��40 P�f�EU��@
��$��R�  8UR�v"ƀ ـѪ�ұZ�֭�MUi�բX��MUTj�KLثY�T[a`�e6i*��JiT�0�$�IPR��  0��23el�Z���b�(SL�ki�
�ƅa�P���[ke �5�f�T���������F�jT� J�[i�$TT!
U$��Hp  �I
kJؕ�4�j����UM*���%[j�Ք�5m�kj��m��Đ6�P��Fkh6Ŧ�m&V�[Q��U(
��I
��T� H�\  Υ��Q �J��[l[m4�m`j�%"���6�k��U�ZhL�[i6Ȍ6�CF�C��#F���*�R��U ւHR@��   �Gm��k)��Y��Uea�U-�F����F�ԫM*�[2�Z`�UcUVh&�[&jխ!Jњ�5��!SCL���!B�T�p  ;�ɦ��mYV��&�Ҷֵ�ViV��������4`6[T�l5Z�Pj�h��
i0��-�ʭ��H%Q%*�n   7Ni"���h�T��iD�j��l�%[F�R������@�4�J��hm��ՠA�UHɃ@5�J  @ 5= ʔ��5F���@Oh�J�Q� P   s �	������`���`E?�P#&&�a�4h0� ��ddF�Q'�m5�CO5 �I eT�0  LL  ��vv�p�Z��8߳��Y^ך^iZ^�p�cp��(�5�׈�k{[X�*���~�2#TQ7����S� ��8����1��OΡ�}!� �N�$	��O��B@��&A��	XDEAo˥�Nv�V?�ݽ�ق *28q�4�gT0��&1�.>�@�A?~���~|c���ڜ�n����J�#s[%����W{)�{9�ֆE�$/ew�k��Ż�ð��57e���oE��\�����w]!H��Ko�'�?'�.]��Ux2�S�=��B�ɛF���V6C���u�yG5��7V�T�M�d%]��FAY,3D�(��-2.��ذ�L�Ô���[-�%��D`6��3Y�'��7p �� {l���wAk���f�k.��W�oב3�Q=8�#S�Q��7�y��`��d����E��'��R�t���[ӺfYn��[��O���z`U�6j��+Zۆ�iP/N�@� ��cvl�U��([�!�Y�5�/r��6� A	�4�_bR5wZ6��e���0�ŷXEf�W�F�z�Ʋ��z�U͓֡n�!f�C%cWP�Fx0a�r�-���Kum�G��Zc�V�n8-�N��I���MIvܬ��8�DU�t���y{r�nֽ�i��Z���ʈ�"�C��m�z2�#;�ĬS���&�צ��Vܙ��B�����.�=��:�t��nZش�|�����c��V�=�"[��a��vpV[Ѻc[@8�m`�ˏ#[ %i�g)d�|5fj���YF���v�P�O�j�($����y�³5�E$����t��a���;Y�z�[�.Q���4ӫ%	��q��! wL�P ��ku�kL�&X�f�z����n]�إ`���2�L"�I{2�̥�6���T��5ҫ���-�5��f�[{���nހ�J�u�b铯.nm�D�8aVŬj� �if����F����^Z��=�^�8ť�B�����v�����]#�nm�*�N>��7e?���2lB7�H&�3gV�܋e)���0-̠�㵎V����n�)J�3]��Mȩ [�@�I�z~`S�q�D��r�A�0��",�63�Y�����Z�^�V�*���,l�0+�iŕ��V�_"�o4J�0L�.�hw�"�t�Ʈ0�R�1*�WQaJb�4��a���qq1yh���r�+p	t�ً@���4(��h6(��[yn�]-u�z+"9��r%O4niB!y�]m��SW��9M��9��v&�T�� �E��̙!ǹ��dUq�,A���#�ݝ
�n`t�:�qV3��'6�wv���^r��1z�i�ͫv��8��i��=��JE�a�:46R�V�k6j���GSm<�ҕ � � ͢j]ހ��q�s���d.�koc��'�#z��e-�Pa�F5�P�?#bQ@�@�����1fَ��nΐ���6��"���30�v��ƙuwF�s6���Ĕ�:��۟f��K�a�n�3j����Xt�<�C⾵u���Ѽ�y�� ���Ӱm$3�lM/��a�X��wX����e���Su%��+b�x^���i�R���T��(�MǴU�[�w�d��Fbo3\G�WRN��Y�S%U���'VA�]f!."�e��yi��lJ��hr����֘	��K� �h�x���ð�G��iq�dq^�n��8�K ���!j
��,�UPˁZ���H�We:׍%@ǅE.�"��:bZ���3���0�m�c+n�t.�7M��'�]ʀF7I��N�F4٤E�5Tњ�n!��(�)J�̥�Z�6�VQ	�dh2=�����f�IHunbpV�dJ�l��j�ay�n$�S��P�+W�-�N�؈�W{�(h4h3z��R�5R+�0��&j ������%rUf�^��N�Ȩ6!Vozdv��d ���I%x@�yu�$��c5��P�df��-'IQ��w��+DIc�x���ՀQU(�ȥ�ڲ6h���م�;Wz�b�="M�WrV+l=H���4��-,�E0Ex��u��.`t�D��I/e�`Qˇc�:��Z�oh�/r����/r\�#��$P-P���
d[�0h�l�v%0�ƀY�V�;�h��5�㗶�Ma��������R��B6�6�c�Э'�q���V���g"��ՊF�1cU�i��+E�lRu�(�n�8pňY��D��F�"�cc4��6�iY'r�V��X,��4v�3i]=�+˩)+HŅ����T�s�
��	BY��&�&љ��T7FҺڒ�6ĭ�%�2m�k��*K21N���ʽT���yA5�J�B�^�]�kjM� �7�nm��أ *r^�m@��tNCJ�]�v��ƣ��N��]�n��Ij�u�*H���P^2�+.�۸�:��9����N'~ע��v�Ɂk��d٭'3bq��b�m�A"���*�Ce�yRٳ,b�yW7eM2�J�%%��Ի�l�2ވCr6�Xӹ�s%dukFJvه0��Í�E�bl.�q	@������9,ɍc@��sY*}��A
3v�ܤ�+tŢ1�7�B;v�<�v-*�c�p�Lˬ�3f&[[��6�Ӵ�~����-�5&�wt6[0O��T�7)�[U��% 4����WS[��N�Um�b��{���e�Iʂ�!1�si]X�B�GG/m�V��drVEq�tIˡ��»N�6\H�3��6�
�"���K��y�F0ɚ�\�O2���-��+U���ˣYy(&*C��tX@3y.n�v���Z������Ǖs��IY���g�qM���vb�z��m17
�d:3�Yn+�pn*�PM�9�Ln��A.!�%Y5���jЍ���]^��ܱ��l��֓��6��i"�R˚>T�"vd�k�ͦ �wǣi��(�ӊ��"���fɑ��B��LS5�&$���;�L�r�����i��+h������e
'
Vh��ߌo2�Uݨ��L��]�R�\��j�D�`�5�R��+�x�ѭ�nV���Df=ܩr�O���H���,T�F�*��If��[�S �D	p�Z���x��"U3mͩ-L;���n�����yy��`��ѭ�b��!8�_�7u�(5����7��1bB�9�\�,��l8���/^�6�,6hTe�2��b�B�S^��W�D8��CX���aa.��V֛a��SHh��@4����`�*[�(ZD�o+l����۬1PٔZ����m�(�2=ۢ�#K\�H�3���Ϲ�x�e����xMa��X�=p^��P:@O4�y���Q�4&�-]����	Y�sv�"�k7N�e��+I�e�·��]-H��j0=+#yv��/#L�90�ijo&d��A��GF�Ҏ���ݑ[U0ԫ�1چ�g��Y�h	�c�x��b(��l�7xDN�e�J��$u9BL�u�P��	��V$�<Wl�ܧ*Ÿ�n,t-�6�z��y
�ޤ૘��ճ���2�o���Y>}{b]�jN�b�t�TF����.
��	b)���w$�5�D���L�ha;���FY��X1�K�M�Ksr4ث�fe�Aǌl���i�Xt.Lٯ	̒��WI�e!Z��a�(�8����w>�^��FU���t�M���Q�	L%a}3w&�8�ё�7qh�s^�[p����1���0F�Y{NQ��A�q�E����c�7E�"��q��IQ{z"�P�*VU�˻b�O�u�I���]LR�
|*jx�X�[*3�Њh:�{Ww�dİ�25)hj�%�h��^���--.d(pD�'	��N���l��^�b%!�˖蓮��!���+l� m��l
R��ve)�BNڬ�ҭ �n��(3��u�*�]Z.aUd�v�QFVP�%2����Z˥9e�����w���%�16��2�ɻ�,��X�bJ������SOw;�;7����B�H$�,�Б�x�u�ӠD�E�Y��b�.Ah�m��Q;:�Ӎ#O�E9�flX��I�n��6fCoTR�K�����.�J��=�K@���	���Gv��ߋ/M�U�1�m)OR�w�/>ۥ�"��Ã��&��3S�j<�/�=	��誖,�2�*9tN�B�x¡���K/\6oQ��F>����{$��Bb(��Jd,ݷw��7n�M��$ܖ��r�me;I����;��n�Mh�f�1
��Ô1�#	�扉<Uʺ��:K�^*	�r9j�9Z���8X���y6���/v�<�e҂T��O&�T�E��m!�ݓ*�@ƅ���n�Z�4�$ܗ�3]������3d��*D-��l-;[Mѽ(Ю�iC��x兵u����Z�庑�k
ŬR�˲��6��L��{y�H���	��n�Uo+X*�V��>x�htt[��(bT�#us6�k{�GXX:��Dtnv��MZ�B�p��̨����@_��r������j��jYLZwy�7J����#ۺF��a)Y�K��Z��m��A���R*#��D�,u�,ϕc6�ɹ0����AYy��GLII;�V2�+���'f(K�3~���YN$x]z�ʉ�ܵ��Ռ1���ě
T(�Nu��ГDD�E��n�bZ�l�z�I�SY��*ڽ��n*=�ئi�.�����^� a����z�l�m9����C��rL�z#r�A��m(;{$�Ӗ-�n�J�"N8��6�K��j�n��0���\�n���M�	jfƳ�&U�j�/Pp��Il�nX1W�5xg�#���p* �.�"�,k-1N��A�r=&�:�AS�mG����Ք�M�*�:e��������C6S�Ws5�a�6�X��t/(%W����[i9���k+0�ٵ��¥'��Ż�X 2����eKD@dݰ�Z�%nhK��e*����Z�tP1^�*� ��(��v�^�46�<qQTݺ*�u��9�w�2��'1�Q��QM��96���D����f�ݷa�R��u�c�*�iڵ	!�`���g����,	d��e ��m�^���a�yM�m���LKF�4�,�w4K�7t�����@�����A��%!��-5�o^!H����hV�m�6��7)ۈ4�K�J�q��;�a[�$t+2��I���Ԙ�ɫoXQ��o@x�X�7��pŻ	�1��I&����iZ�r5&V3F��h5t(m0�%�$M��(�hL9�6��&�x���cH'5��`�i��屧S��j/
���WY0��l'�)/�I��`du�vͥbx䉗�0�,)�r\��^;��H��0e�wu���mZW�}b}yMc����C7$Z�Yل�d�pi� 6m�Ad�WYk)�e2����-S)�(M�	�Q9{*�ZR`C+0m��j�[6��!8hi��1�eP�Q�MR"CP��L��F�FL��L�+�VH\/4��)��W��t�n�˳�x֑�um`����ns@95�^n^�rJ�C�ؤH�3���ݬS7- �m$�Qv�ݱD��4&Yq����a^Pk6=�Â(�P�*��+n�Z�숐��R��ux���oj��QB�Rᔴ46��2�B81���
:��/+�-�.��Q<��V.h�X��ѩZ��RV��h�Û��; ��\nӔ�kZd�ج�I��u�R�n�͏X��a�g���2*,Vڈ���r����G.BXz����ڬo�Z(�Z�v�����e�cn�Q�U1+b�r��k �ڊጃ�b� `b�2�\Ԩ��^T`&������e�92��ϱ��ٵ�B;�0Vf݅��#���k�ο���S�]b�1u.K/&�ƛ�.�Z�ź�L�e-�������Rk�*�	-X�ch莤�Tw���N�6�M[Mc�V�#Q��@c��(�Fn˘36BB �Z�P�W��k��i�X�藴]$f[ �jnM�&��݌�f:��4��[�x!��F�*X6Q�i] I�d�t�"����"��X�4p�2��y[V��^Սk2�2Q��S�kWJK������0��{�����6ӆ���ڍE�Du��o!8�O�5R���8�]lZ�������dC�c$:����1�i�B�@�ϝ-h�w�	�-�p��]^&�����k�q��I�ݙDV��ٖ�㬷zr���8�,�i �mV�)�%ohd���p���6�M��գJG[B�?*jE��jЫ�1�\ݦHP&1�A}��i�����ff��J�����j�R�*Q�52n��t^�LĢۤ)h�vP��v�ދ�`e=T&�������BJ�blݣ�2�N0K�u��e�EM�uv��"�P�0 X�����؛��w���R��6�m2�H��ג�`�;p �QR �{�%������q-s ۬׃p�Ʊm�) �(
�*m]C�CݔĻ��!���%�<A��S旆f]$)��W1�s#٦�MC[���j�˧�u��j��v�-�/�kI�K�i8�ajW-\Jg�>��q�*b���_�T��7��0��������ﱱǟWt}������A�S��e�h�:����
���wCK�:����sX��\��÷z7,^T��ue�Nr�CW�S�ăU����f���of@�`
�޴�:ۧ����q����5�R��x7�{�Aa���i��^-tN�N�m����tӟ>;���ɷ5��෯��oz�H\�P�8�޴��vZ15eP	J�.�����KB�:7�R�S�BqY�%o��'�O ������R���z4���]c�ul���Ӫ����F�ĭ�����!W*� ɕg�XM%����NEB#}Dd�ͦ�3���(ue���p��wo��ܔ�v�ѺFR]�*��4m܀S��uM�8�A8u�!�"E� se�/�ĸ����b���V
�W�v���\�Pv�.��$]]a��MQ�Ze��ګ�b���4蕛�i�H2����tk��:3[v�������eXɈkV�;�QU�:�R2)�X��nJ�{�sZ��F��������L��[���R��dq�Fq|ے-Ж��n��,�!ܙ�wܔ|�x]�f��tÃ�%$\rT!`��¥F'XV���Hv]q�]�N��2v����qh�%>W���`���K�(*S�sk�pƫ�\�����@%�e�V>K	��k�r��N����Hm�.J;0���m41Y����sEyw���e��zc�Q�ku�{jp�v��t��������� �bk�@�Z���y��6Y�V�`��� \�����%��D�����}�VZ����A�дi�C��˒����˯�	��=��\y�μ�m�\N���U��i�S��CV5��d���f�r;����`�ۄh�%�=�;
O6:�O%v����˥�sq�ON@ �_	�܅�ٙ&T�K��]�`���]G�-� ͦ3�
8P�x�7��O���m�Y�nP���ٰX@o����;P4+�,B�+��#�Y1PA����
�1}e��p�6�Y6ɦⵙي�!�q�e
��o�ܷ�i�Y(�y�W#V�	wSf]�++v����J��ѫ�<L*��޽��ࣷ'7�A�Ѭ�-��2�E�i�@/-K�tm�ٚ�Z=��@��j2�T+�+�-��>]�Nʫԉ���Ic���p��ѡZ5���N��BS�b�z'j;�zzv%���XYƳ�}8ͮmT$�D�7�A�X����S�Ҵ ��7�I�l��.��}m�:�<E2���:����X������U(�.��mp;4��|n��]'8�I�W�n53��S[���O�p.7z��	ز�=��Z������� 9"'V���Ń�zum[�YM�]u�F�p>�[0�� Ll���d=�^dķ��;*FV�*h�7�+�ڼU;��*^`�;����R�����Ǳ卓WR}�(���N8�k�/��V����������
Ԯ�R����v�������z�97��/��r���:��N�%���f�q��>"�m�[�[%�K1>��jYu.����ыf"ge���[E�u
��pl]CAJ>(�OOZ%uu�RN��k:/Pq6�N,t��¯&.�g�`�ʉ�k���&u�	>��`;����h�����Sv7�K'K9e.߶����ˤ�}�.3����Jě�8���e6�u=�7�`�j�Z�,�$�i�A�Һ��Z�؅%7��F-�4i��;&N��0�:���ύ�oޣ�eb��7�b\�=X��y�xN����"��oj���I���q��6� ��y%��t�b�R�@)�.�}�n	.������]�ӜK�-�{cܿ9�)iڶZ~�n��1��z0L��CQ���Ye*5��PX���q<t���z�ˉ�w-���m���󫊯��·�xp[hWe��[G#{c�8W7͌�g��s���Y���oU��V��� P�Rԡ�����R9�To���Tn��-����/�]��V��2��nѦڮN�wm�����B���1�n�_	s�j^�4����eh��������qZ]�8f�
��N�Is�*3�[�q����e�sm;���#b�&;�j��־jI�ӹ�e��֚����*p�]��,\�F����i�h�d����	��8]]���b�
��c0�(�B�ȗ+����v��j�x���|�v�\�z�LҵTXd���+w�6tKцV�U����l戵�,_R��ʧ՜͊���j�2��+S�B�M޻���b��1�B	�Sm,`�R�-W]3�����S'R�T�{*�D&l��mQ㶺��Z�"�CRWS�)jD���V���Or���@���MoVg���Ղl!��v���g@:�yj��wa��%O0�^�Me�1���Onn�X�]V����X/�rq����v�Ol�V�p]��֡{¥�f�zb��Z�!٬�0� _\�[��P�;�w}.�1����7��y�������8:u��s(��;RN����k^�H�;��	&]c&�� q��ΡS����Μ=�v��l��5��U��Z�hH��yF�Y)Nӕh�c�H;�iS��ej=qh�B�3'��X�ON�)�Q����T���u��,^�I�=j�Q�"�Gԯ/�T�.�*�zʷ�Q	A��n�9J��y�y��:ۦ��o���i�-�͓/:�o-+׎�r�(��ȯB�w���ګ���MK��S�E�!͙iU�3�֗.��6�e�p�cB!�9�a�pֱtf�:���ŵ\�XvS#���1��CZ�{�++ks�Е'�5�L�K�����Wב]���Y�+~pө���v�Lz
yS��ʎ�]�4�ΡG�9�:�X:׉����'��p��N�d�3V��fZ2芹v��om����[g~\����6�Lwl1]�l��}vՍ<��)I5?�=�a�	PL�9F�ΉL��i��:CM,�qz��$e�+{�ha���Ç��Mh�f�I�]�,*!wgm!-����c7�k�K�m��B,-\�o���L�;PeC��.=\;�ʂ��G�J�Y�t:�d����b��G��Bt�yz���R�#��+Aъ���x"��ݩ500�p��S�l[ȹdɎhϥ$j!�6�MZu5��̡#�vR�5�Z�U��<�Q��9�g�+-l�����x�̻������R��ḑ\��.x�d�Nyۚ�x�!%Ly�n�sz?�!���r��z��U�p�w(V���M�5V2.��آf@v��γM&4╼3j� �GC�L��EX�XшSwD^������n�otl^a��cxkM�b�c����Aædp:�����t��
�+9��C|'�8h"��!�v�u�t�t�٫�v�`�-�����XJ��Y�ʔ�����Յ:na�+xƗ[V��]����Q��T�� 7��+�vT3�!ͻ���hgU�;\w÷z�r������]]l�)�;/�Z�۫!j��hN�9��yE�gm�:
����K�@�b;ч�u�Z��@�u�o�K�Y�,,IՏ�q7��E�E��� �����)A`";Dv�.��y���W(�(�x�{�Gwe�EO�d�2�я�B�/F�}F�5ݑi�&��.ї�.9ܻ��L���oW-��CFd�������i�/yٜ�fI�{�lLL�"��t����� �� >o7	������UwNN�a�f=��fK_�.� �î]4xw8J�qM�U!/���ck-��w�Ĵ@�*&3V���E�6m�1�������Cpo.�� ˭Ss�$�(�yf�]���P<�ǲ+C���e*���X��#;O�Lt���o�.�\-B�V��T/C�(�噬K̺���Z�n��:\2tû��"b믮ٴ	�q姣����N�7z�Fv�7�
����&��N���t)ү�;�������\�Q+}k��,D��K]��]�������6足|B�8��s2+�ZF��*T��v�� ��,�]�#EX<]��@(�N�g9���r��Y�L�����y,�����@�}��C��%'͒�#S�^����wsh��[�жF��y��K��1���raSV����[N�ce���ݮ*aa�t��a���K�D�� �4+������7�u�p�SNʺEQ�aG�zi͌l��<���^B�m:}>�v�\FKl�YiS���g"�h�`]���D��^�kjPڔ�U��+rj����es|\�)�*�����\�ҏJ�T9���D ][��U�ݱ9����c�B�;.GN�1�q3��*�2A�ono*�{Hl�U	��(��G�c�t�q7P;�.`�_ڴ���̙���jf�*sڌ5{�X�/2�:����|��٭���A�6�3q�%��+kmD�R�٠\����V��E���S�:�to'p�rk�ra���tt@���E@Ӊ���3����P(�J�V�U�� ��j8��O��C�e������Y:�*���<�W�{"�űM����w̍�[�|Gm\\<5��ʅ���I�.��b���5{�\�B��d��Y��s(����hk��Euϰ�ٽW��j����p��G8�:�7%��uu�s+�+:��[ώZ�i��Ij��̭�B6��u�4'��=�4
�MK\+EI-�-u!��k��L=��{�c�^�
�w�A��Һ�c���=�k@@T �i+7��K1}�N%*�jy uǘF')1��`���dRΏ�s�heڠ��t&mbc�]r����*ϱ��b��6m@0��5$�R�V����M�e��`�Dk�H����	���v7۸�����+;I�Rn��������j��3o>�KT����L�+�Sx���	��^e��En:*�+���#���&:<;�G3z20%%ӻe�iR�5f�#i�@��[��5ev���ˇ[�5�43��a<�)�,T4Jf��er�M)z�h�wO�����V���ٮ)zvX��H�P��E{��\dw�/vuc#������r:Uj���n(j�m�����4�̚�m�!Qr� ��L�H�I�.�)Yٛ�&�ܢU[jjl2f��=�!%�".wS_kV�ծY�`=����/:����C2q`�GM��,klQcˡ�C��z`BF,J^n��5�f���w��i��a���WYcM�B��ẗ́�5����{�q�ش�'�Z3W1��^N��ɝy2�=S�JŹ5fMO%1�I�yhW"�A�����W��θb�o�m�Twb��
�w��u�\���M��m߅ku���F�a%�����2�u�sX���җjţ��e�:�T���l�cη�o���o7�r���-�ԛAb�^L)��ʀ���l�F�t%+"�<є���O�m���t��R���Zgm<Z���t�%Z'�(T�w �QT��h�@�����b�5�.����N�Dj���N�s����5n�)���u�B�2$C��:���c c����tgzJ���a��1�<fHк���귐�#gm=�6��^V�-�.��'ua��+z�ish��a]�W��3҃�lF^ۣ8^'�*�}X��U�\�8�P^������'l���D�V����	�Ȑ>�q\ ���T1Z����:*�$^��/5'���.�l����B��̕�Sbc/j����K�J�(*��#�ZHe�ͮ�ʆTR�ެ\s������ܟNSU%t�pӷ���fҎi�*K*�+OT�w;m&�aɋ9c�� �	��m���)R�{9-ް1;}��Y�*��t]a��\�s�q�����$�n��)"q����jbST���ysY9�򸛊��]_� ��8�G�z�/��Ϋ
��2Nz8f�5��I���(q �^+ʲ��X�ty��ޥm��d]S{�_jFo[��.qF�q�.��׳:4�v�Y���P62�3;6���ԟ'�R���K���A�/��5�ݭ�Ч0(��Թ�?$;z��E�����]�)�}Yr��.��E���iS�,jgZ6��0+�4��ZM&��{���Z����mnCQ4�m��ܰ�+��N�;�fn�"�X���nFWb{��,ǔ�6�nn��dd��W��q
[[��ol�s���I��kV��d�,����u|;�����]��o;�]9'dJ��v-I.ܔ(P�����Ηp������7%QVu�;����;$���c^�F{�?^�������ߘ��k�OS����nݝd�@�[6�{E�݊�et��<�gt;4sIQƢ�x:�KU�6�c��]�Y����]�޲9|�����e�=/��3�?N����=����r>E�u{]5	����q']�}��a��:b
�<�9uO�H���(���j�ʸ�h<��U¬�ǜ�0�	�������p#\���Ռ�70vަ,w��u��[��9������5���ѣM)�\��( �-rH1�5X@E�rQ�`t0��*��!���:p�:�l�z�&��F��|�Vwkyڕ-� ���n�wj�RV��c"r�}\��kb[4�ȍ&%�K�ޙ�,�*�VI��R����4N�k���M��a��ά��t?�/��W]O1r}�	�ws)�y�ӃUv?�H�\6�.T�5|��+ݕ�,XY�Q:z�9,�Y�Z��vMS]#�ƞ��4''9U��ic�N���ø���f+�n���)��Gj��v���\v�A��z��u�"�[O��ǫ�*��I|��/(�q��e�� Պ�V+�*�b���+��Px#X����V���l\���8���g�TO����@��H.�B*�dGM8����V}nQ���]���^�븞�lj�<]�'MW����^��K6��f��l������P�6�qb�r�۸�^MgKh��U*�V��$����Z[z�c<X�͜To-(qrea0���Y���)�-:�6��Ư��j�)��Iee-�kg9Ow��0s}Z�x��;����"t�S,����B8;�3��oE>�����L͕�z���m�Q&p�b�ݶ�m��+:�;�/w�gup0�Ri�zi����+�6nޚ�ql<6;[��,R�f@S��L?N�����3B�aB٬�[��t�J�;Y��al��X��]g �blVz,�f��@���h�Xc'�*����
��[�K1srt���ԱS�w-���!9W>g��#���N���@���3Mڴ�A=��[�<���W<k����֮��z�>���毉9]�m��h���X�Qy"�V��I��Ė�ťY���{[�H�n,b8&�.��R7g���=yȪP��r��P��zյ�ծB����n�]cqWP�y ����ł�����30m
���5��!+�᝸��Ds
���}p�s�%ch]LU�z�LY���뱄���I4�Ֆ�ē���Ǖ���H���Ga\�AU)+�AH㛺�_G�F�̗J��,�����`ޗ۔ M��K-$>e�}�W�ۚ�4WV��1�G�]���=����]�M�V��H!`Ţ�w1��f`�JR%]^�Fƻ�i��.Fc���n"vi����*���ޘ����s>�ik9e"�2mg�J���r�XX�_n����:q�u5;Vb�Cq�H�h{g;��Z]A���޾�O`������Uӻ��T�T�u��,ᖶ��3*�1�Z�"����\��iޥ9�B5/���i
�I:�$(�����ð�ˬ�y�|��N�K�][F`��Wk�k\�ӻ�.ZK0�ޗ��:1����p�P���@9T%�*9x���v��ܕ`X4vV�CqF�t����W\��
� UvtHO<���(�)audk�\���M�D2W^a��1�~t���P=�H}Wy��L�pFjաq7M��L��޺W|X�W[]�r�0GcR2��q	*4��:%�L�]WC*�V�ʶ�+�N*}{�r��&lʛ�$J=Xrv�뻧5��iV���^R6��:����ܺ0�grPӀ���y
�O1v ̢8��׼��;�%�V�X�k�Ȫ�2򴽺bpo)��˻��1�37D�#�+1(�n��V>�[���;9X�i�[ڞ��4j�(�����z��wط�d2�<�M�N�w��v�^��6U����o;M]p!E�m�y�b�˶�\�_<c�7�t�t���77Z�nb	X	W3F��}��N�I�X4-����'i������Zyo:�S4�a/d�k�Rī.��=v�e��j�fa��gU�g�n�.��Y5��U:x�9t��-��Л���oXb��b7
V��v���t�k;2�G8��/��Ev)��D�z1݈�xM��+��c�B�ʀw�C�mH#3��2�ѵ�qr��X��U�o��꾵՜q�IM\�{��b�1�z�a�����΀Pg�`U��e�c2����m�us�Q��b�����'�9�Jbxx�/2�桺�ԅ�f�Ob����ڲ�-t�2����ۨ6s8ۤ��Ւƌ����W�a'B��R��Ζ��7�gk�ݐ��T��u���̤��}ܩ�ͦt�f&�e<����"��"A[cTX�B[�%�i�lGd1�Wc�''%��J�g�|�^�Ee�f��M�ݝ�x�DRslk=�l(.�ú"'��pX����G��軮�gR�%p�a3���M}�`�+-��eg,r	\U���\C"�5��;;��ݴ9rJq���y�B�S��9fX;�`Ō�
���v�Y�>��������YSM�B�"3�B���׉aQ_՚A[;�b���(�i[���A��n��!�2�Km7A��#4����(;,a갗�l�oP�(e�t�]�6�+:i���U�]J�]�ٚ�j	tQ"��L���vc.#�N�OV4�F�ל��[j�+w�@]�PQ��-�����=���Yd��wp��5Kl�`2���WA{q:|MH�[��r	��y����
�Hvl�4ל+ܡ��{�c�tõ\z�0��[A]��wZ��&�WYG�R��Si	�+Gn[R�\ź(e��nN�c*X2�i�Ϸn�ϻs,��V)Ǌ��Ƴ-�@s����-G������_^	N=���ؓy�f�L�t[�4�V�=���ɣ�����,��;I�;7b��k��
Z��hQiP�^�Z�n��܃����i9.���Ϫ�k�-glӶ@w���0f�C�����t���u��/�,K�����e�+�]kYqveֵ/�o!�-�� R�re��|���']p۔�;�8�s6��ʂ�5�̺�����٠��v�"��cʔ慪7͖�F�DY[v�bmIV����*�.ŝ���5�ְ�q���&8G���$�ْ�١Ep�[�h��e��M��uy}/���V����c�,\�]/vh�˦q�,��[ɚ(L�ĝk3�.�y`��4m�Sf��罴��SS�㈮�Fٶ:/Kv�3V��W���9Z�v4�V��K���=d�O-RS�������(��1�7�M��D��:�_�@e���et�gkv���kJ��`���Nշ�j��jѥ$W҄2.갖�a���H�IzL�/�'ڊ�*g]��VvGt�#	XfY�5P�!VY���[�i����U9D�]�a�6b]��Ǡ4W���S�n�ka�6v��0\���3�v<��\�n����[ݓ�t���:YB����о�jWoҦ۬p%��SG4=W17��e���`�I�i�|s��G�۩���	Fh�V�5�;�'�rq�{�st�kj�[���n|�����+/'v��`v�ة�,����0Mβ�a�:�ps�����uK'&�E"�.rؙg�~܅/��;����ݛ���(&1�� �Zw�靵�Q��$q�����bF�L �wf���Vz�t�������x��!:�vbc ��A].��Vn�Eг
1�����-�Ŧ>Z❶nJu����WLV���-�H��{8�e���h=�ť�c�./Y���ȷ+u^(�]��
]�r�h�-��`�[zU�xWWq���y�VЁulz�8�qk;
����6�ϋ�W��6�`n�@j`q�c�Mt����9���=�H���x7NR!�b�.�+9k��YY&VJ�q�����f�#0G��+©�5aF�ђ�S���`4��b���m�fegn4�QQ�G�v��-�\+ur)�z���HPd�[�
L���勲����c��
��Ċ(���l��@�ww�zscfEg�ܵ����ņ�6�a�9lDl�vK��-�Z�p6�[�Z��>���RhH��<��W>�;tk�E�fܝ�Y��80�*��h��@+�.C�L�V������ԾdK�bO`�	5'wna�t�]��Yw8ŷ$
f5�pi� ����wN�3wz�sj���˭h�cQ:��nƄ�`���5��֕b�}��^��a�b����{�ݍtp̯�T�&}�"��\�{d��7΄8�&�7�Tr&�j��&_��ՠ�ھ�{���	x.�A��J�j/��YT�k&RQ�SQ��u:%,�k��h��M�],����h	����A��b�r�F��*:ls7r���'b�m��>	汊�U6��;t����3�$�;E�R��ss5ȁ�1+Bs�эM��" n���LY�{ah��m�R�㙑T�:(>\^��B�*��%�:����)�S3�ud���:�Έ5�3���-�$����t���Eތ�]��R�i�V�
:���%V��n4
=mRsg��P�1}k9r���)*m���{X��f�ч��P맒w�_-��r	��=u��J�`�E9�y���lG���	�V�G��)�}M9�U�:��S5M/�[�{���jܢ����F$�s������{	��❼ը٬�Y�7~TOϗK�Rh�>b	��#��g��&�u��&��n�Sԣ鶄�-C\K�W<s��&���5�B��oDٸern�
C9�}؁���PP�V�f�uv}s0D�6�YMG�ݭ�]�d&�i�tN��ث7�Ќ)v
}�QE�3�0Y�Ӹ�2�V�$����s���j�ݹ�V��żh�ҽ�\���SS��M�0q��;��Ut{yM�ݴ���wFff�=���W��e0�����.��v���9�Y�^�Me��qv.)�+��������a:��핤����EI��.��M�6�F��b�իu�S��]�	��.ǘVp�֛�P.�Z�9�P��+m�qp+@	��N�5�ް�\�;�j,���� �Vt륄v��L�cy)�Z�[���T��,QV�8�a#�Ӥ�Nռ�P��f����jh|8�7�^���:��D���r2!|� ̙vJ�p͕����B�ԇ�V�I�Yi' �I�-�]�]][7z��Sk ���Pvk�oX�55�9k<$G��o9�"�cv��h�������X#�*�4ܦ�r�Wv(Gij);;�Y�K� ,�kY�vP�]����N�J
ʶoffcIe[H�����ԫI��p�\T��w�աA�opč���Y�m2�u	���5V����k}ƅ�Xo7
��OI7�"2�+����1ݜ��b[�:�l�3q���p_]�Q��5�X|}6�Nv栍�[��3^�����)�ʬ�]�]6�Uٗ7�:�V�ep)���tf��l���mZ��l
���K;�]uĒ8�t��$���l�]����e�Ĵ��H�x�����M��v�a�i�2�sD�̱pC����!��@V��]y���V��i)�pVc
.�+fV\8䃆����[�MصB�.
m᧝:q���l,ָL�Y�[R�$F�k��i	u��6�7�/����u�-�i���[ܶ8��oFh)�n��Us�A�ƵQ��vv�\�T�Z�bf��b���Y�z�xK��-����n+Bw2�(���WQ��\5g���y[�.�2WM]�()fw@�^>��
�;'����<�lgGSz�We'�o��+��'8�sS�7��9#��y���z8S�j�U������N�r�I�;��]���z]�,V]��wI����]z$���Tjb���[�"�e*�fG�c`���$D�V>�5�욹˕�{Kuv&��s�%�J��B��]����c3KF9�A����S�J��;���<�:WL��f[��C��+�(�V	h��u���>]�v���lj��f�n��b��aK�\)P�����q>FS�4X{:t���@�{��ұ�WS렡�b�tP�X�@
i��lVc�g`�}9��d����}��y����raKY}�����9h7 Ү��6�/��bt�q��s�G ?��7���2��ɸ���'!O�@N��o>M����Ԥ_X�Ub��L�����"�t���s�W*훴r�H,�|xN�K�y�^N@{X��k�=8d �>�7�<'��)�9���.ٌ�Ɗ:��������Y��q���a��k]���˼����DgD�K{K�+t�Q�9�(�N黎R��t-\������IL����@:�E�ؔ�z�D3t�"_9EZ����1��t�줾|0k���|3�
�WZE ��ßh�tc+&i]���qҐ����R�Љ1}5n}O�)j�wt���-�T�a�#e
[ױu�5���qC��dLN �,:o
/�v�f:�Y�g�J��enp0]ld�vB��/#���"u� ��pj���JⲰ���~P�5���j�/��m$��A
$�����U�qi��ܫ5�a��2�{ư%���ȍ���<�P�=���#�+l�*R�}@Lv(��Ȱ쳫�*�tsB��	5fuF ��0�Ȏ��(��,!WC��K��.�Wֹ�}�������";����;+��8���=Y���_>5�U�woV����L�S��{���O�O�	 H�,�``<b�B��������U�*�l�ԗ\��)��̔��Q�\8)7@;�K�\�M��a(�c��*� �xE*��;r4%�w��D�-t&�x׭�:�<vrB�������B��p��v�$l��C]�ܣ�j�]��L�o�q���F�Ɗ�X��\R��h�R�WWm�]�fP�s�o�KZ)Q��<}Y�m'W��K")�	�bd=��/�;�i2���l-%ӫ��Y�+\s��t\��lp��Ǚ��b��4*u!eF�����s7����_�拡{���ƴ�'(2��k��;�|��i.�(9�тU�Ki��ͺ.2��Gٳ��	�2�K��js���)���lW[:I��=��w��H��{�;bh���n�U�"�9��ydu��i�k2�z�rx�]�v��]��n��p����c�S�u�(
�;0�7�1�Jm9foQ��C(��{!���X9�*�gZ�(���a��E�g\��1-)m�YA��ô�W�+��2�PNLOq:e�
�M9ʻ%c��i��Cu��X��@(�Xnv�]+��`���R���ԔzDwiIu��=k7U(f������1f(��wF2��5;_P�3�w�%K�=Y�)���C�&)[p��Zk(�Ys4ͦr����qêB �2�d��qU�Z�xB�I�-<�Ma��]}����q�2t�G�8����E5׊s/}k�k����l�5\�7WK]���Ft����{b�-��"=4a�R�&%�U����i&a�\��[lq
��(�5��������U��Uc�Yib:��Ӊ1�eW,4�KJ"�(=QH��t�,��j�V*����V�V��&��-���TU����h�C2X�iQ!��������%\B�*(�,E1����*���ӎ��G�L�h��"�D�Z���Ku�4�b�et��L��s!�\�m�[\��q^�]J�EQt�-TV������jr)R��* ,]8�&�-�E�E%lQj�LEuA��rڔ�E�QZرTՔ�2��J"�����:�F0Z� ���T]!�(D����*(�IQQQ�J���J�Ƣ�R�����m�X���J(0�W��6(*0b�4����F��t�J�*��qa���'ο��X��W�~� Y���ә�[�'p�QwVi*��h�nQd�����6�]��- �@g$�Ґ�R��rL����uu)3����9B�t��p�P3�J����N�����wZ;�R}�o3�Oj�=4�}}�&R��21�p�{(�;Tە���a梢󰞫خ��*���v*�u*�Yr��0����zn߯}��,���|/�;�~�Ny�*lRo!훹�X�TO-md0��#D���_��O�L�]�=C�!HlF�^v��9�ɾ}9*�/��7BJ
�m+�r[�-
�����:��HQl���Χ��h�kB鱾{�;���d6L����j��J,����k���ҹ���P����I�5w��J$p�T!�G��c��ܲ�++e�R��BE�u���Uh�y^im�B��;3*��{L�D��[O*g�뜙���$U�+ټʚy��ޫջ�?v_�D��:���(�2�40{�sjg���Y�R�up���Uc��|����[�>b��I� �
Ѝ�9�5Zt�N�o��{.\�
v�̅��E��y��ŭ'���a�� k�۬WXv�&�8�M =���Y��g�w���ԑ<v�����>�6i�m3�b�=Z��:���x���K)��^.�oFM�k�uj�8�9����_>��W���tv��ں�ҝ�c�\M�l��wg6ˁٞ��!M����%q�wz�T��q�v�Y*��q������;p�ƕ�y@�wP;İ�nԺ._[�m��m����T�bY�5��i,��J��68N�����[8ޭ�Y��vYjA�ASU=�1VP��#�T����6�2LgB�^"��M장L!���`�ώ�����w��NyS�rU�-��Nvw���]��P�296���-��+j�p龱JdJ�=L�^�2��.�5��e�k�YS�(w��J��S���ڦX��Alt�7b1�׸��l�3àS�^jɐd�p�G/c���<���l�thçe�k�CT��*dd;�٢�Y��i��[W��[{B�����6[ȑ��3�
�]�h��[z�<�X��9kpV����N�ԋ�iʸ�0�U�CL<
�^$)��f�����&��o�{]��a=��Y����N�U���;!�*�0NNq�c}�7q7*W`��OS�f�n6
��D�ә!8�c/379mE��9��=^w-��8>����G._dq�k���rs��vĐ�]m�/�g[���Y\�0n⡮n�ǧf2=��Moa��=;jn=��o�3�~���i�p��JؚA�r_f�;�w	�u�8��sͰ�v)��zV�+���=�M	�L�_JGS�=�]�f^b]Ov-J���is��տyF��+ޡ����X�+e?)!���-�u�Z��\��W��=��}�a��N�����@��s�]�=i�\��E�]0;�M4{���ӧ<��\�E�0����Y8�891WIgh�e�:���B��2U�	t�5f�P��ص\4�;�/_[����Aw^٣�}]!��Nӡ��^����Z5���0n�Pʳe�Y���@?Z��ǍO+��,`ϛ	9*�����ћ�J�^��b�}y��_��R��UNR�y�uL�$���7�z��uqCC9a���
�;�K.iCUG])f��RQ�s��[,�ݮ�Z.m��o��w3��9��+f�қ�Y7JH��2�E�����-�-E$�}�Z~�ک�1�W�u�ħ�(	B<f��.gn^��cd�Ix�z㞰�F{�$��Pݝ���!��jS3Lٙ!m���<�dI��PG���ᚻ�P�Bd��a�7���P�"�k�Z��F�p��4k�)b�n�=u�)�(G�<LD�U7��ƕz��Y�vdH�&��p�T"�z�E6���)�7��K���.�z�߷#��WrK=,�Z{���#me��9�fc�Y:�4�zmZA���͊p;,u{��d��oA�}*.
��xn5���o^9����6P��5�AU��Ϭ>W�n��Bl��u�xh���{m�Ru�I��_��eU��zRe��]��Wm�b�*3U��6��]�v��=�;
u{:[9;�)��{�շ�κ�Sv������|G>�NK5b�R��;

5��Ub��m���l0	�r���d��w�a�{��LA�2�1���&�ќ~�ޑ�����/FK�p�z3
��ޚb%3���2/���M:S7�媚�5�].��L=�
Bށ�e��4��+�9������]����/g��9t-���Ɗ�.,��΃��Jۨ�5���FLe{p�v�Z�if)���ͷ�0Wb���B�t��ho�U����4A��Zd��6�!'�=���VO��o�dߩ�p-������T͎�:���z���ۛ�7���"�N`؏Jƕe�S���H���1@��T��]HA��N��~/��V㽖ɝ~��yJY�OdSY�q?s'x��:!�B��7�Ι��
z�X�O�4F�^�f�g-��ܩ3h1�n��Aߏ}�kAV��~��P4�_#p�n�@�c4�5x.�cK��Cbt8�o�ϖ�}�o�6�}���m[������xy����!	�
ɷ�XJ��>�͔o��E��N4�9�gW$�g�Gs�����t�p�RBS&q��b�*W>KgWglr=�g���jj�ѐѸ2�1��C���MO�_�V�{�i����Wu��l�68>�3�I�j��+1��M��с�}��E�-c�۝�_��ۯ���p�ћ,P�o��j��5]̯4.�eSVrOU�Y��,�s�\�6п�gʹ�7�z����÷np%{qt�"�b9K	nw	���!���Lϯ�nf{M\]���Θ]w=����jȉƄ�z6l��Cf�=C'��*�<��y>ޜ��2K99?T~��՞��	�>r;6�zء�S�Cb�b�m����կ9ӿcr�����-:^!���f
�*��u]E�&��U�͍m,�x.α����I,�Î�W�u��(N�����%�U�Y���v��G���Z�
���颺q)`9�>'mȋ6���w�1zl;���MD�;�f��dh�V�]Ь���e:^Z��<=�v��Ԩ:s��6�J<�y�\��|��d�cI��PS�؜��qscVV�5G.��%�� zĖ^⫸����bbn���\������ }V�s��ذ�}2�o�!�N�]�V�^[hj�w#�AB����jq\m�RC�߶e`��Hf�����LBs��S�Q��W�ҍS[n�:Xޘ�ߓ*�ӀBغ����}Wj�h�u��ru^v�^1{t\bU�6($�	LȄ%45�5!Vq�Jw��\t�mb�U��Vm�Oه]=0#�Tyؠ��i3�� �Glb�+�`���+�����9��WS�� �ja"��G �,5������*��]�
���e��!C���rP�����rxi��7!Ø��YF!ƫY�p�]�Nic[���o(\�YH�lVڑ��dGgnu.�;Κt�U�Zavé�M�zוQni���0cBm2pcSB�V�gwog^!���f*�ڷ坱A����b�i\�ϩ�4;����Cr��NO7:x�=���3�O����{~z�eU�"�FM���
"r�'�0�4��y�~�㳲��������]*�@"W�?u<�"k��Nt�Į����D�W�mMV�u��i\�y�Ȟ�����;q�JNRoX��>\[��Dgx���|�t㤚]��9��6�˺(FP�{+oUcZ�;͛`ƺck����T�M9��8܊ŧ�s%v����Mf�(��e�#�����j;OV;t2R�9^t�\;��+ʓkU-˚Qn��\64IJ��t@.w�%�'��u8�)L��r�i�c���Q��9�_��H�6|V٣·,������ڞ��Jު�:�J*S�i(��p}�D&C�4��V��(Eй0P켾涪��u���e�E��jTu��)�
��̦���Δ�+�:ޫ٨��NU]��<������xdF�^�O�pfS.{��e���7�ޡ�.��[�ł-Ң�'��
�N��v�+`�,�ۺ|�G��*9c^��T-âR箽���k�q��	�sR��Kl�j�k^�ݮv�3O�;��6���N����X�Y��@q�؍cg$R__����l`�v�{����"ga��ң�A෯q�N@cVTX%��m�m(oy8 (H3��Ui�7�ϥk�k���[���o:>���%��d3o�C��~��Js�NV���e�gFN��:�����K8����?#��_<;��2l>&�z�dc���d>$���ّ�O3o��׵���߹x����Sޖ̤>+;g�'�{'�!wR���`�{`G
��9#Am�Ϟ�'^i�H�����x��Kio���4e��6�����*�я5�������s��KԼ��#b����ʒ��6��t��)��w�s�ɼKr33��&����g�{�b��:GI[b�T�S����uº:/�9������1j��	-��YXp�u�#���yet��vΡ���8�T�w�k�(k\p�ĮE/t��	�[g$κ6�,�[wՇh���{�i�V'�J���r/�dߩ*�A�q�]�v�u�EgWm@]9;l���ט/���8�;RҞ����tu�`�YÖ�Ǔ�gnk U��AQ>��$�lմ��4���H��T�9o�w�z�������I\�F]�Ю�����J]ݛ��tNp�a\ⵝ��^Wt����`�ӯ�����讀C�s `�����ݣ4s�jZU�%<�O���.��ո��s�Kn�!H�N��yA�L�s8�m�Y����Ĝ��j�$^�!�:�q�u�%��ha��/��)��[�_n-��Cn���T1#pg�2[�<�"��U�Y�z[�w7��;޴����4C�Ʀ'��A��e�`5��ὃ4� �9
���������7Sc���S[��U���a�̶��-�U�"��(]t�t3g�{-��[�ڪh,y�fT�lf�(��z�U1/�������nj�����(M9����i�$^z�Ј�3���WGy�[r���q����ПL���2�3�l"�zSV�qU�V�[Ԗpx��`hVP��:�R>��k���@�=�|;?0{�=R��YY�D���y�;�l���m�J�|�P�yy}w �z���J��j6���`A.�kV:����������#��4�q\��++�Y/��f���T�W����s�6��7d���Tc��+N�ݔ���UcB�Ya*9�9n�S����Ce�_V]�Y�4�̣]�Vgge^P'���b�*���� ��f��)�F��vH�
�=�5�mq��I]���-�Y�Iܜ�,��vþP�K�sO~�}�f�5!��s��%є���9��:��Gf\�{s%�8�k��U�az� ��X0��ܡ��r�N���.���M3-����(����
1�'!(��,bq����hI}N�`e��J�1�b�hEz[�9����RΈiwW�J�B���Y �Iq�5��i�:}�`�%�mWe�V�3sF��;�:�&�e��&e+ՠ�i�Ca@tZ������W��^ʖ���6@lJ,Z��s5T��z���6�������Vv�A����p�nu8]�g�.��Av���ͽY���=�Js}�.�%�FQ��ǫ!v�Xx�ˬn��52��V>���u�:�v��ec�8K��ޙD1)��[�u��oJ�9ʄA]���k����qe��YE�$+x���la�w���(d�)9F\� �``�8��1��s�S������(4�u��0j�;bC����[)�$ �sKR�&�t�J�k��5`�o>>���MN��6.0�x��B�V�����V�U��1`�/�y|K��!Q��r���
�@-W7ܟǡ���E���.�����\#FIy�ζ��鸺A��裨��*�v;��J�6��uf��УvH�����OQ�ݶ,�Į�`���0���$H��j��J)�/2��l,�+e��,n�6 �FfeC�5�P�?;neA��Q�����	g�*��B
*j8�MG��0����,��x�G��b�����2�k�ceӧH�U��%M�6�����,Vm\�%�}ݡ�v�"+-���aTH��dX7CN�8V���y��+o[�Y�zo����4�� ����
{�Tv�2U`FP���*���z�JE��=Օۯ:���g~E��\�+�P"��Mu����B�>��3Z�X�gJ/@���	�d���Y��i�k�]I}n�bX2�_kuY0��v��3.�n��%G�[�	�Ѽ�K	��+ �"�.֡LFE:�z��֢r�����v�7]LT0�4��T�N�&���N����oc��[�p�bSR�U' �Yu@|bK/����_T�v�%��i����Z�Y��ft|���Gn���w��n����eo$�5��4���ܥ�{��a�����T�O)��~L8�a�bdA!1h���mh*��u�Ң �F(�"
*�����,Xi�+V�5�Z�F���"0QUQ�\Bŕ*���DDQX��"#�����"*�Ɖb�ƭ��"�Z���AAE�j�EDAb��ĪԤƈ����*�`�` e*,T�M5b�EF,��b��4�Ŋ�i*EEX �"�" ���PGHT�"�q��YHV�j�[E�J$�TQfZbUE���\B�f\E0��(.�"��Qb����TV�,Qdr�%j�ib�1*
�M2���(�+LLAQY-��J�)Z�J�)����J�i�RȪ�����J�&�"
�W-`�+1�j��ɉQWiJ(��b�u��ӈ�֓MT��CL,E����"��K&�դJ��et��k&2��U��QEef\��J��~��q�5ְ�_�Zw.��G(��hW���W>�f��aVCv�d�� �[b��(�,���J�బ���Yir}3{qzvs�6���-ag���kX}k��&�����9��56�֣�ͧ]���ctV�ߛfE����:(�{k2�-Զ.�M���]s�Ⱦ�Y�OOy0�r�}�C�#��^��N����%���Y�R�/wC�S�s���_�5�V5�o{0�li��	q���$�	9Fo�X��z��0�J��N9�Yy�%���$ҫʬ�-Fs��ֆ��-�E��ngڷ�=����cs8�ّ?S��3_wVM�QP+�L�A�.�%mk���3C�yO^�*Ѹұ���J�sb�y%\��@G�[+��HJg4\�ս�(3A)�3¯�Pjɐ��(C�±C��[[���e�|��Tu]0c�;�r��L)
�|r��T��*�,tqy�ݐ��Ĕ�Nmz6�ʅ��������c�f�p3��^ׇN�f�l��xCWn�6�x袓�{�����f��c����y�:�gn�|��!�5p�@��,�:_j7�:u���1�T�mL�v��Sv����9���R\�Z�ޥ6�%��h�./v��ڗ཯��[&�m��0��֦"E���'s-�gZ����nPL��|��������%��!�:�i�ť��9�U�כan�7t��J���="v�P�;-�S9x����F����Lϕ9�-[cܛ��j̚�-����y���"6�\�9�g*���2E>�Ǝk���P
q�>�~����k��᳭��_9�j5��E	�s\6@��W���[i��;Q�w*���FY{)[�N)Ui�z�F� �b�
\m��=���]C�I�q3=��y<��k.j��vGi�|lp�V���W�g�ͬ{�^��2G/yEp��K�i���'��F���$7
�4:�:�p�{(���|矻������{�oZ��VM���-#>L�hi+)U��l���M�PVv
���\Օۀk�3���Ε,۲Ðҫ�ѣ�Fg�	3�S��Ҩ��q��}�CW�k������1�K4�b�_�Śd$_9�gh�7#��f�.u�E�22���5�2��9�n��9}�ʂ����5�x�)8�l NV�u��}s�}k���V#��l'p#���2����Ƿ�Ք�`Q��LJu���/�e�2#Z	����9���ډ��.:���UЋ�h���;�#�]b�=�%�7��o` �_'�����=�w���j�Z'��q�Ī������5*�_��������B��5�D�&��j�"�z�i�]���3X��;�w5{��͝�RY�q<sTzk�fd�4L��U��w�͞mվO�ɜ���b
�B��l�Z�ڪ�;ĳ*u�9O��8I��P��s9��j����k�������$��5#J��sMg*�y�*�V���i^�֭��a���F���3�WR]�8�� ⫕9|�N����H�e%����!�7�Ugzޙ/&�x�{K7�c�fi�Kf��f�佛��""IW�̚�9�4�yؖ��ϱ*��S�Wq)�ŔF9.\;X]y�v�ZEui�0B�����vV��sV�_SǸ��"GA1�]�α�=�*9%��|泜�PWO{��[�S��#ީČ(E$e�����͐��(F��9���L�e�%�#=Y춳�{�g��zzw���#��C��|V�G$�f��l���q�^p�I\�yջ�"�̈́�B���ɻd�!��d�'�է;��δЙ;9���mm� >�D} @��r�m!�׹��&ӳVOPힰ:�2m�v�S���u�چ�<f�;:�I�2b,���IP�OZ:�k^�����k��QH7�;��F_�<d���0>I��y��`k�rO���C�x��Y�	��Y�Hm�u9�@Y�����[���=_l�N��xz3�§�<���m�䘋9�p&�V���Y'xn�'�a02��OY4�����y�>d<9C�x�m����c��{O�Kr꺾0^ݣ��5����l�	���2v�SﰜI�Laַ�8�X]��$��7�a��I�� |��2kT�Vk��C��6�GȏG��	��>bfkV����~ �8�ݧ)� )���8�����`v���P:d�C�o$8�Xh�జd~�a��	�3 x�l�V2J�9fOB�����J�.�~� {�E�d��I���d�.�ԑI��w��~�;�&��l�h}9��Y+&sy�RN2t}E��Ci�s~w�ߪ�-��>����A��>�����>�i��r���'O,��q'z>��M�y��VI�u7��z�C�o$0�a@�G��� �6��s�Y�ho\d����E���e�J�����+rK�|ik;yr�V�6q��3LtL|G%R����=��L=�&;[W��,��A�����5K8���ԩ�J��A����@U�r������E�׳:�[Z.7o�-ŝ���]��5���u�ơ1����<Bz�e �&y�M�N�w�N3�O|���Ȳt��x��8��'HO��ެ�L�v|0���7�/�)���z��|$����<��BVԝ��N��w��4��(q�<�2M�$�N2mOO)=I���Մ铌�7ߺ�E�!Ӌ���\3��>���l�#��!���z��Y��{�=d�uϵ�$��=a�'l��x�2x��Y'�:�h���&�9lo�<����n��3�7��ů����� }��xq�2��i'�s�z����9�'l�o��OOS����!Xz�2z�X���{��'����?dA��=��������}�o$��'o��I�9�$������C��ѽd���;��|������0
ÙE�2O��dY=g��G���a�j�"�W������jM�|!�:`s����5&�|��v���`m'O�7���S~s_3hN2xZ����3	<B��7���os��o�W��}wח�'ޢH�#̏q��Xt@�����jI�'S7�|�m�O(|��q��`m��|{� ��N��>�;Bw��6��Lf�y���yk��㺾�i�l������A �{̃_}���,���V�ՠz��&��Z���wI��&�Z�|����$�4���|<SQ+�{�+�x��Ow��:�7�m s��ԛC�LChN!Y=;�
,�hw�M�	�Sh��:- �&��	�]y���hw��� a�?-@��L�Y��}�X���G�x�y�L�$����2x� vu��tɈ��o$6�P���d�I��dm$�]�z��1�lRiyd��u��H,������{��m��b�^��]��`|�0hM��@\̡t�C��&=����!g&�!���-���n�[c�Sɳ`�\�a���6��4/GJS�[�����;�x�ݪ�'@��RNQ�n�M:̴�Y�҇��pZ�j�G+��U{W���(�y>����'IѮ�l��Y�����I��2d�RNo!Ğ2b,��4B�T4n�,�l4�'�'��>aS��^.�G����vs��7{�}�#�}�P������]X6��h9x�=B�Y��d�]�q��XNo$;d�Û�8�P���	�M�z�Z���������]y�~g&>$��f@��Ě2��IY����29N�q'Hm�g���2q57IN'����LOӌ��7�P;I�A��3�k�q�|��|~ ,=�xV�N�I��'�,P�2u��5�5'L�	�v�8�$�yd�&�6�G�$Rq>���zH�l�:#�u_}Ӳ�����s�*�;tã�d����mB�ŝ��&Ұ�x�����d�!�Y8���VM�L�I�N#�����>F�Ͼ�O+7����=�nǃ�������'̆Ӥ�L4�C�}�+�ۭ����n��<I�%d;a�Mr�2N��,�E$��~��󮳭���g|�T��H�ʺﰀ��d�}���}�	�G��o�	���x���~���LC�s$�v��(J��ꇬ=I�f!<C>�9���ּ��)�u�9�p�Ny�'Ȥ�����N[�)=a�ڝC}`C��y���	������	���o����M2t�s�Y$���&�f���1RaJ����ڽ��G�Y;g��C�d�Y'�<�xN2O���m�v���OP8��l���|��joX�H�$��!>��5$񘇝��Ϥ�ɳ�6>~�z~�>��{R#�b�+�iXs)zɮ���z����7l��,�d�ӺHm�I��,��f����Bq��>��o>������^jKS[ש>�`�+�w���!N��[��C���ׁl��n�ܱN�ЦVQ�DY{�\o�AJ�鑙jEܺ�;�n�2�pp{,8�P9qЊ��VMn��3qI|��m2z��g{�����O˵��o��WW�uO��u���>�='��}��
~�BͲM�s(�|�-�I�'���,&��rI�g�Om���<��L?cc�� ���ʨ혯�;f���>���p;�g�����8�Ę����$�
���@6�9b��P�[6��N�@�i<:�4�,1=a>fw�k�^�gk�����E/�DE���Ͳ!�8��� ��n�`i���s�'�:d�|����IXh�(�M�G{Ȥ�$Էh�wl��a���f��O�fA�{}�-ܭ�c���6zG���'��04e�2N������I����L�!���d��9�	�+&��
�	���,��	o/�}��>���V���]�[lQ����}���t�^d&���
��C��!�<I�:Ւv�i��!�m�u�sA�'��;��I�&"�kx@Xs���tvu�w�3�6�M}����;I���a7��+�'5d��Mu�H|�t���|�\�+$�>�'�T��!�i��!ĝ�H���\���0�7����:~��&�2��쇨�����a���ߡ�ԕ�SV08���0&��q���N�1!���J����.$��;~��r܇�D�{O������>�ʁ�&[oq��7�5$�'G�Ri�$�l�;d��|�+5�&��	�S�4��8������_f��~��l�_l��N��IRz�{Ch���A�2q��No�xɌ7��!P���+	�O�C�x��T&��r��'�>_7v{eeF�˗,����3l'��d�N�(��'��q�����4η��=�C��l�v釜� VJ�7�E���t��<��;�*k;��
��p7�WW2R�sg5R��M�:i9V����r�c�k�1�C������5R<��))�yح���Î��<��g����'�F���<O�#��¤���[�[|�]�ܣQ��L�ڑܝ;�wv�+���J����E� g��.�}=@?,�I�Y5;�x�l����	�G�}��� ��0�;d:������G����� a��)7�\����u���	P9=�;d�8�2��Nν��	�N��I�RMw��Hu凨dݦ�a:@�}�=x�z�|�i0�����ƪ�M�tw�\�|��>�����<d�=}���<Hte��i��8��Pdɭ��<I�,�E����2r�zÌ����RO��r��s#>������]��|=g�{�����������sTRl�<��l�!�Xz��;E�FR��&��
�윱�{���yyDx�l����]��w����x��O���OXN�Cl�:��;d:9�����!�:�Cl�����E��=I�,:2��&ϽL��D�u|��ʫ?
�z�N�u�G�����M��x��w���;v�&���f����	���C�J�'�=֡=aP��|�qsX,���Զmd{���g�c>HV��UY�H��8}�$���N�M�������ē�t�Y��쀰�u�3l������htɈm�}�@P�v*�>C�NT}_ӱV|�ōߐ�B�6����B��o�2wi8ɯ�&���I���5a�N����l��x����S�m��4��[�6�L����(a�3}�?�#�@�R�	���夘e��O-��I�t�s�$���'���h�靰4e�0{O�"�H@g��s���c��p3Lvܼn!u���i����º|���I�M}�8�d���Ւq�S��Rz��=aSL�����N��'̆�B�a��>lx{��Q��כ��e�wW�b��4I3��ݎv����ep��}^��͛I޼�uɱpH�^��	��c��_�A̾g��$�*i7Y��2gw�Np�k�״a�L�u>����;��\��6i��3M�Nl`�!*�nt�[�x��/�kh9�Gvw&�5�9eOw�^�˖^1���޳�~;>3�|����2x��t�I�La��8�X_��|�Ӝ0�RNw3 |��2h5@=ef�|�w߾\3�^m��-ش����]]v\w���g�}�Yd�=M��{a�d�'.�8��,n�@�-n�q���o��#��OM�f@���'�������}k]}�;�!�$���xN�{N�z��q's�L`q�I���y+ ���8�ݡ:�9���e�ѻ��i�=��W�A���u�7�k�Z���v�m92�i�d׶a;a���:C�O����]�;d�N"�D���L>�!ά�L�oxq��Yn�Y�$�WW��r��o�b~����� �ro���L`h���'�(̞ug'L;�Y'�'��1��Y;@�'q��:@�s�r��4�7�o�3��Sv-�ϥ�]��ڼȨ��� {�����N�!�s ��Oh�;`a�'l�m���4��z惌��[&Ւa���d�,�yI�̜�ٮ���~��3��sK��{O���q�|zô�����=f�vs�'��Χ>�Rt�(z��N��<Ր�2h�x	���z�O��${�o^��f�c]���_�X��v��'-:>�$>`q�k'�OP��m��C�o$�3{7�I�	�u9��N��!�Xz��;d�/���|G����"�!�L�ھz��n]1d�$��=Ԝ�I��'�7l��'I��=�$6��:7�Z��Bq'���>g��\�q�VMoX,�$�:u�d����6��uc���g�i��a�T��=I��'��y'��>z<�q�n�O(m���<N��BM�|͡8��@���c6�=�$�
ß��������0����!�ea���0;�}X����7l^��DD)�(y����3���%���y�T�k~��df0����趃*i��^;�	��-�i�wp]`���od{��C����&��Ho
�A龝�ŌUS�����n��w��
0�xd�	�g�<d�L�m�MsZ�|��s$���:����m��;g������z@�:@�=�>���w�����ka]��;�ܿ���3�I�������R(�M����d�,����'Vɫ@�'�{�B|���a:x�m;Փ�{������g�EK����|�I�_*�[��u� ��<��C䝡��^�C�LC���N2T4y�Y&����Y=�FSh��:�0�*z�|�`���?<�
������y��C�}�|�L��k'�ͲO��$<f�;��tɈ��o���%C�Qd�I�[�d��Mv��{d��g�q���e}7WZ~�|�mEm����<�%g�C�wd;g:N�^2O�ў�m���CL��C���8��LE���J�Fo#�$��o�����g��Q���$�����| ��rj��hc4g\�N2t�i�����6�x�=B��=�A�Y&=nÌ����7��[a�oq�<o�=[�g�����>�J����|�:|I9�dY<I�,8�+5�	�!��t�`t��vR
���H�q;�xE�m:�;�C��ߧ3{���}ý�y��2�*�cP�������m���)4���u��v�1��s\�4Ͱ�u�l:d�8�a�d�����Y��
.*-������ASV����߸٩Ev�7��Tsޡ�����++yr��N�������[��R��Wu/I��_^UE�������u��ۚ�
5��YD@��E,�]v �.�����+?�Vw�l�@O*D��)�@8vOS�+�u*�wg%w������2��H�V�y9��x!��"����'��j_J��}��qӈ�6R���D���w�q�y�!Ac���S���3kP�{x*	�J���a�dϙ}s�e=u���t�,\�W��57�X[����Xs'A8� `��i��:ꙴ���+���p�KJ�-�E�ĕt#U;"����l.z����R�^,��Fqt%1[�x���)Ir��s/xq��W##{�5�����Y]׽�>�"3qK�uݵ��R��vi�Xy���4brE�ygm@�z7�P��D�';�>��a�]N�S��tR�Q���D�D�7�p�Z�;��Z���s�b��3�z��w7�J2�9��/��qǷܹ��:�hm�QL���]Z4�X��o��k+C��d��S�2,Ew�2k��=w��s��m�8^�X�ʆ�W��!�g/��wՔr�ϩ3���d�Pke���1!n��u�R���<�Iصk+���7�k�/�e�ޜ:��p���m��:ܩ$W�g3h>�ʼ�������,EΕ�����Z�%7]]���;qun��g���l���Ô���s�j�n�n�%<+�NB�E����m`�4���h�\w�T����x^P���TgE���Z74�O˟%Ժ�˳j�V����q;7כ!n���6��ʶ����=��;�Lus��n����0#i�[%�u=�z���4��h���CS���]��Wx0ҫf�rRw2���Sb�����vҽ���DACn�
g{��B�����M3qҾڟ3�Y&��&]=�i�bM��m�%K�̞x�Վ��o-U4�4�m^�A��5����]�:�Ӑ��>\A$�nnXRa>ZN���lȄ��*ʥd7�A�B�[ȭ �˔�/���k0��D�O+%S���n�H-l�*7	��W2��ӼiÓF�JcL��q���I���i�C/-�j�9�d���F�c�\�f�����7��ˣ�R# Px�P��vģCH5k�br�n��W]�����*p7*T�n�T�5 ��N����c����ܿ��l�G,iգ�(��VKo�f�Gڵ؂�V���0����֬�5[o�k{:v��}s35�'�pwڝ�U/�$Ļ�'wr�َ�e��B֥�[�a��|b's8Ol����E�}Էxt=/Z���e���i�����>@k�oX=�7zR�麙�wV���Y];}Y&��7Tl���M�CP�yqr��ݘg^�F�\j[���r��������z �O��GmTbr�"�"1DCQeJ�G)@PF,�hUE�5�EX�kd\B��Ɨ)�Z""��STPX,���cZ*E%����V*�1+YQ���aX�����J�*���TZ�b9n�d�"�WN�Lk���Qm4���EET��[Z[e�Z�#"�Vb9�1q��+lh�VJ�-2�2�TU+*"V��s
�c�B�`�)�.P���V�%sTV��L�t��cZ[(�"��-J�`���K�\Lf��T��n5V�$\LJ�2�.��f��B�UQr�X��	�b��"�5���YZċ��U������*,S)Tm*��1��E�DIq(�QBTի-�J�A���0E����La�*$QciU
���D�Q�TR,D�+EDm�VZ���Ŋ1"8��ƺs
���m��UбT�c���T�n�B�U��V �D|'/���a��g����ݞ�̦��y�Vv��ڙqm��pz�+K�e	y�u��,�&��Y��lJO��99��� z-n����qY?[kE�̻��]k^o�?��>���Φ3*�{2�s�r�;��UTM��S�7���Hҧ�^hm^�X�W.������Z} (��}�6�T�p٤��#9��+�m��wy�3ܵ�b���ؘ��r��K�ռ7 �zG����vM��J���.�)]�]�"���Au)$��P���Oi��o#.IoC~��ս��Pū^�����U¯da�$�h���[�H���s�f�֐�#��b�&i�o{�����~Shl��j#&6���ki:�Z�+#k+�ԫz�%7;�n��$a2<FsFú�m�c��%�ݺ��u�ٹ�j#R�ڬ��*Oo=�A�NɊ�{��Z���P~�eV�Ҫx����gH�}>���8#Z��O!�_TE]����zB��q���qDiS�Ό�2i�>��l��ّ��G^�2�`/]���_sHޑ*��#�(�V{�;Q�
����P�#8:s[SuB-�vZ[h�s��bܰ��S3�[Y֮|�`̵DGBbw5`3�i������ov��vþ��q|?wdT��k��b�F��������;M��^�N�lo�)z�]y�3�ِ!a|#p�]O��\Պ��G,��}���ycO�8��O�<5�D�&<՗\3Q��_Vk�y�i�]W\����qj��Y9�:��z�P;��XO��&�A��j�˺j��ײ�f�k��.T�xС���t�����.}ݙ>G$�7)yx���9�z`�`.�v��i��\�s������{�>q�VgU^���ҽ��M]��%�����v&#�P�hn��g5���LN����S��"�!,�����t3P�8�:9���������,�+<�gi������xNC�|r�riE�[=#s��V��)�\���m��E�g�O]�����=��YU�2u�#�+*ǻ<VDx�3a��+	�����Y��I�<���H�P�.�8ЪU)3e!���T��í<�YZ/O]�����xr�ի�V p��E���P��e��,����Nm9��SNlmX�Y����q��IJy�6xgn¾�[� {�%�����f~��N;r�OS��܉P�d��~���f��Z��5��d>��a{4���Mm5ZT��
�Y=_APo�q��]L!m#$��ðW} �����[f�mw*�C�FS��{����qg1���;�����	H�Lʶ4�i��T_M3�̛����O�n�6����u��͊<���JhV�BZ�wٷ��1��� ��~倣�k��0�{�*��b�N2y3r��#�I�m���W��.�:m��O jby;4��2�+��qiv��Ox_��9�3�VdI�U�)��T���^]�;J�st��ܰ؊n+^���+��%��r8^*������e�Ԫ��Wjan�	����1��-K�Y���ʹ.@zu�+��Ȧ�T!5m3�aLbXb-y5*c��8��o�K��ՇeC���|)sӚ�.��Bқ����v�
���!����o�$ʵ��]Р~��鹬�L�Y\gs����iS|�[�|;���sõ�S"w
��\������D���.|�*��ዖUr�������R���aɥ���{z���ݛnP|*|wmߧ&}Hj���[��>�RyBJ��d�W��>��=��N��ּU��7��{fZ��*ަ�-{X��.=Xџt�\�)���K�6`9u��si��z�u�Yb���)��E>=Y.��)t-��>M��FWf˚�~����ͮn.gKhd���Ayb�zE9��gK��P�/b2Xf	鋘z�"V!�R�sW��a]t�/(l:˛ya�bg���8޾��m�>Z�y7�gZ��[P�6����@��C�{�	4�w�U���=�K�)�*ɺN�W�#>R��bF���5��ˮg�"rj&؈�u}^�uR���������bT���g:�i[M�S��VlӔ�EgH��A�oL����Y$<贞T��C�+f/k+/��J,Ф����kRӆ�)����:˻�D������=+MN�]̇�
T�;u��Lp�K
G��|4.��쾖��,u)>c֐���K���GkavȬx	��[���NPŔ�e���N�[���i*�T"{qg��xz/q��r]l#���
�`F��o�9�k.���L-ɩ�T�n��n�9T��qc� ϻ� ��5lm�	P%ʮ�n�7%��J�Nn�S��{C���4�˚|L5f}��wֲ��mNY]��ˇk�y���w��A�^�t���Ǵ���QY�ub�[������+���V��~(H��+�ٟu9ԫ-k�[�ˠ�Ӡ�%����엕��|��ρ��1i�����^�՚���t��tv�`\P)�^s�^�3�{��Չ�v�_%��L{��x�.*��9�u��ݑJ���H�&Aǔ�Ȋ�z��
J�g/ge)/V�Ζ�+��{��g��M�2�\�w�P�
%���v��ɂG�ü��5��9Ǟ��9��''/�B��9�cc�����g�]����}�]�fl|˗�v�C}im;+$ӻ���n��/j��]���	Ⱥ�߽K�<��m�6ߩ<Y!N�9
}��q<��w� ��.�7)Ց��1�q��u�;tPȱ��N����P�ٝCsT��\�ܖI�E{�������f�_����U֭;�By�b}Q�Ϳ+��u��:wq��?U�ه�[�?)���F���֫�����H�,��\u�pV�%��w9"����-��گ�է��EN�-��Y�j·��^��\$h�-.���2��t	�7eOu�З`#QX�w_r{XΫ��	L�!3�f�X�9���r���ٵ8"X�\�.�Cm�|L{W1��h�3"C�윣���خg�_k���9�@�K[;�7^�bt8���O�<4G"@|L��ᚍKˮJ��tֽǦ{ȥΆ\�Ym�Y��hjO�����x�����1׻���AcmF9�Y@\���4)3��@�UK�f�K�D����U1r�v���z�UM̊oh�x�jG�[�}*\A�)�C���GM0��M�cE!^c���F:a��F	����3�\���^W�μ�4����
�t�b�s2&m��C�����p����H�FԎLNY�wK�J�	 p�]�,)י�o[�nLy(s�����'S�ܯkrw=�{�	�a9s���㲾�Z�Wvdrːخ�ٷ����V4z	�ջo��j�8N96��iu�y)'�����?g��7�nq��^Ϲ�W��oV�/��	�A�teךp���V��W��ݭ{'�'&�����^h��]}��f��y�t�ʡ����EA��#1�4d�-|��������{6d��8�M�҅�)B�.8k��w�ӎ �j4�s�|������;�D���*������/Y�=�O�/�P�fu��ũ~�0g1�)�3�h{^����KQ>M�ύt�Zg����FJ���]�oe<�BR)�x-3jg��jR�X�]���w��s�7}N����I�Sa&n53�MN�M��[L� ���I�٩7��l��
[� ��-3>��J��KW�f��k�g;�i�r�Z��aOx�xk��م�,���t�DAqo�\��χ�s4�zk#��ڝ
���ygk�+z)٪�![� f9n�v:������7v�s��mk��B۾�z�}�)���<�ړ��ğ#ʳ(3�Ly��+G�3�)��[�����z��O�����{���56�)�l���F��~ɀ����9�b9;/��9�p\Z��s�q=��a����o���5#��:U�u��{���S��r���o�����c��;�ƬĎ����W^T��p�x�Nڻm�Q8�H��N�./l�^*���ĖT�/A�ה�
���[��̡���$d8�H�MZ����eM<������ٿ5�O�H-�ŏ��ixr���Yݭ�}Y@ν^��_��x��{������ �rsƏWW��P�y��g9�cd
L�$w��P�ʔ�vWv�o":�-͘u1/��N3jL ��Q��̡
lP��:E.=C��S��q��=�#y����[�.��h���yg�t�B�f۬K85���cuP����|r�?�W�����^M���:yMt��\�iS��E�f�]��-M��B	j��y����dc[�ת����BIa��V��v���6
c�mM�&��+�b�����å*��[���;�>��"�� =���oR�WԾ��#�����m�9�cзH�(\�M���J	���˞�Iʼ�T땺�%Y7IС�k�u�=N��q��$��#�A�~��e�BÂ5*��_��)���=vbTJ9�WJ�6�hit��'³����S>oL�0��aU�vOG]��S�;{��b+���J���v��|�����K��p�W3R��]	��<�"F?�5�FA��V]��yTm�	F%үu��<%��PW�
����lu��B$sxi��/��5e�C5Њ��b`��=�)�Ҋ\��Ջ�:[ާ���h,zi�̛�4NP/�%u�zsi̪s�ҩ��`O,Gi��L�Ȼ_a��6�y������ǳ��;W�R����(O�9��t5��ʲ�k��ݫ�y	����WR�/�l��[�A1Y��<��h�f�ov��0�dh���\ո��i^d�*���v(�zG6��:�kx�Z'*��mgTz"��73kU��R����s�PG <�oj�}�N��̝ٮ��V+]x�����9���6\�_)��e�Y^��w=3�Cg�M����^;]I��rtcWn��Ws�]�v����<�
��#������RI�щ��N\觘2���ޫ�1b�|�ל�v�r+tW�Ԥp����>C�L��1
3ݾ��%�;_��oǆ��
� t���@9I[g;�Fu�w�>���/z7�#�J:~�k;P�K͆�B�t3>��b��n>�.��7}�������[F��/	��{�9����֕d�.����GU�z󥍵ts�֍��Hoj������En��u��D�� ��+�nS�0��s�ۀ癔̻Co�%��{V��3�]��ɳƴ�����׫oX̺&�t�Pa'�h	L�r�;B�ףOH��>�.�nS��R�}��Y�\9f��Lo0�t3���9�X]{�[յ��Ty�e��)�r1b�u�q�4=˟��)Է�a�oq6�:{�Q�-���4i�s�[Y�%�ncv>��
˴e1���]tp��:rR��9�J;��޹2�+�N��Z��u�Yۇ��Wg=d$%�
.o�r7l�ٮ!�4�Gb��pٖ�Q�1)�f��@fh�6{2b���78\/�u�
���^,3q����j��*wutor]�ŵ��xWed��l��/���c��IΘΛ��9w�K��,KPm:͕z��t�M�4�g���J�N[�*^b���bP�y�-S�����QUt�$�m����SI�ܭ��|""��NP��L�J媒S:�X��¬b��+��R/r�f����V��[��_&���(ZWMJ=}��V��in y��Y֔�f��:뱨�9����,�ucFr\��:�傥X�6�\�����eI��[�ָ�0��r���j}�ݍ�(�E�t�sĨ���Ӥe�u0�jeQ�ɴ��j_�2+!
�3k�f�K[�,����p�6��)V���;V.*�6�rײ�D����+�;��a.#�����@��l�E��:Wo+�ݯ�7��,b�о]�Ȑ�O5������.ȭ�ұ:
�U��1ZP�M��1a\���W2tŷmh�o�pN/�MU�p��&)�u�,S���Q��.��r�;Z�Oz�ƎA�My������<�G�3�]��+��y���'����r��h"�s{Ox�FpC�~
�q�t�c6T4�ӻ��gs��wy�4��k��wk����'ui@�z>���"��ߴN��NiC�v�k4<�9��dO����?��߇�kQ��ޙ$�	�6�C��2' `!���v�O(ZR����8� :���|B��_r��lZ�S�b�6 P���NNYv�{���6��t݌�^J�V�u��Z+��8έ��-��3ɓ�
f��u�#��/�Á�3njʘʲR �N��iP�x�
̢��7.f�x>Zʷj�B�ӫ�R�<�����fo%��mŇKY�0��!�!p��q�� �|`�0��eb�ʵ:kt�4; ,���Xo:Ƴv�{�<퇵���#QvdX(�q��%��NV��vz�ٺѴhV��R'W��'�Mw�ee^����[W��!|�2�WP�&=]�Haz���'RvmR��촪,���n����1�a���W��m��c���D�|�B��6q<�,�n�v7�I)�91��G(v�8���V��ޑ��r1c��Ftᙦ7}�Dzlƭ�T/���D���o&�iۖ�M���n����V��S��Uk����"������VQ�*��Q`�
���E�X-KTKljGUb�"����TY�q�dĳ%���F#Fw�&��K[�Um�f��GIQ[U�e�cm*�e+d�DUPf&+1XbQU�1
���
�%J�qȪ�DX��LM0+�Teb�*"j��QLʱb�b�\J����3�]R�*�mTr�X��Q��,"�TՁMZ��)J�-��� �R�V�5��R��U� i!�M+2��ċdZ T�U�"��&ed�[\�!�(����A)G.��SLF��m��k(���c�b�e�(�+kJ��
����5�F�V��Q��eTc
�c"�Q@r��̷M�.��Z�1q[H�ӎ32�r�V,���Kb��V(Q�0���X�ţ�Z��2�"
�k4�Ua�%�+
(���ۋ�,�@eo"�;m�s��J��P���1����u�wa�������j+˸Q&����;T�w+I_�xx =1<�S������Y[WI���S>�OJ����1氵:�L]^]�[NkdM���meT�e��خ���I��rK�:������6���r�)��o*����L�8�b���[�=K3+�Bz��t�r�yՊ&o94�T!׍��H��3ٙmz���U�0��� Q�㚹$��}^����,Y���C�����D�r}m���j-_3W����u��!��"�F΃��ɜ۾Y}5��s�'��k�H�����3i��&�8���mtr�������A�D�rIe����@[�P�T3�u�J��1�+'�n�7Jh�����P�Z�dba��%m���wL��}.Fw&��o&r.ɫ�-Sy�'���;�mC23��͎��7��k�P����׵	ߎq}�<��<�����AYg������(G���܄7j��-�w�r��� �9WCz��\dj�lv�8^��^��d�goQp4�s���ѱ�m�709�-�pU�1���9������v�7�A�7-��{�����je]�W 5��]�y�eܚ��/N:;yz�>��E���� {ުc�o�����o8��Ṳ�6m�X��l�N�U��l��k�p�ޔu��>��k��S�	H�L�s���c�]�żyQ���w���3xR~�uR�ȍm�1���8�)h^��u����N����ݵ�f�oC�q�*�B����R
v)�pd6Ϊ��q�s�>�YorS�53±���frzݺz
�Ʀ(vBڱ=��>h;�}]*�
�����+=�u�����X�X�n�e��(��3�e[��xy���S��27sA�09َ�b����r�{6P����B�ηZ�S�E`�OuT�w������n^��)\�ϩ��Xj�n�\�����v9���f֋����79��-���d�k+υD��5m7�.䳺�sUQ,C&��ΌԍI�N��ڽ��"���So���٣rԈ�Dj�ˉ�@�",S�:ݕ�`9C��F�-��H!�j�$e�w�wE�p�A��O֓w\0��ww��}Ö;ZTa!w���9�{$��u�]��������}��7ݕ�.�E/����l�L�$tfk�<�S�{�B�Qbj%?v�S�y(���H����C�#\�4��:Z1*w�>�^NRU��{���w5v�<���2�#����农u.*Fu���Ƒ���m,o�ޡ�UnF�ٵ֡l+�� =~t�yf�<��UαͶ��PMzol��罩����ͥ��»�N
]Q̳o�z��0���f=D.�O,�h����yLS��u�R�V��d�7ґL�R&�͆X�S���_K4����y���_:����F�ۛ%<����B�4]F���N��[�����X<�h�{
w��V����N4�	�`�w���۽7�2��P���O�UK�����]t��T)H����r)F�>��wWwvK�hm�������w��3��0�20B�땁� �R�:�o��R��Z%OxĔK�����Е�����T��}y8V+��Q�@������gU��NY�;���5y�7�O���=q��pLb��H�i��/�RV��u�un��q����D׶�MYy��l����4'6W,'tN��5]ڥn�_�� ]���;�H�p�����<Q���3�*�Y�B���9�9���N��C#��iy�v�ZR����KPg�h���V�V)k�����*-��i��ӳ繑}��~�P�J��M��`�l��ŖIދ/��X��6'�p�h����]'��Z�7��h��MNܦD)i�V���E�Y������~��z��8���	��&:�J�͇u���A��ꀁ���ƩQ�,㇍=�iWw
�W�GY�*��7F�eņ�x��s�]	Gw���7=5� ��<S0;�U�b�>�0��a�=�GjG{ʹ[8�{bljV�ۺ.��J�9����*�>;qKJ �;�Փ�k��>ͤ;��yԩq�<8�{i╄����ם)W����J��g�
"��/,oV+C�bYE�#�LQ��;p��%�;�N\�V��SEz�����$t��Ny���PL4+A�S�"/��
�}6B����)r���>��0���,�|CJ��zJ��3��Ζݗ�F�i^���M.�7kN�>�y�OK��)m�v�s!`1��NEĶ�,��er�{L�;K�:��{���Va���h���7)��u%�<�*Ӣ�'�L�o�N��l��ܜ�!iWuA�ٳ����v�/����E�v�n�*�l��Pޠ�):b��zL��D�����M���0�����;�K��η���ʮ9���4p�U�T�|���B����é�<6V.E��u�Fn���w5���n�6��lf���?q����a���.a�x���g�2a��y*Ztk��\�D^\����3�[�7����X=�3(�ea�x!dg[˲�[p�S{�uFи�~8`ө��%��&��DLP��*zb�����Ph��<:z�8j�x�s�}� x]��J��'��ۋܚ(Xͭ,��0�[TD�J��i/]�=*)/[��1ɹ-X�Eg/B��f�Ƒ m�q%��f��"ガ.��N1���v��w�)���M�ݏ,��s�r{�/���guF/
�3��>����l1\ ��˦��{9w3K���=��-���V���LX-OO����V
�'�yg���^�[x�����-���=�hW|Q��Zx3ô�<���Ag��S�jb�|��a5�����>�/.��̌�W%���`;�7=����M3x�&��~��cړ����^f)"�3���̸�fD��|�(V���9���'7T{��f'��lp
��7Id'�`��ܞp��]�\2�9n��`�,)$y�����[�n��R�+�m>��\7�\����xD�Y/��ul��N��tH놌H�E�(���oV�O\pp��:B���L��ND�go:Ϋ�S>�ɋ��\<ӛ�)yq=1T�*��Z��C��wbT8�U��u���5����X���tn���W�3t"��r\1yN>mp��s9�|�ٽ�q�ߋΆ�y�y�p��'���p��*�0DÝ��Q@_U#bzm�8+{-�V���Ԥ���
T���E74dt2�H肍bH�Q�1@D"����c��Ӓi��o*�����f����q�w7l��aW�����6�lFʑ��%���.vw&�!�i�<Y�/_�a-j�_���Z��#�S0a��Ol������}f��GO#�
Q�vU�^��c�'\�Z�7&#f/X�U�,�݄%z�q>Y�"�����Z/�ʋ8�f�X�P��K���M�Q&��/e�M�V�T� W�t+@��I]�zW �xJFY{�V���x�z�·&Y�8Ά�P���v�Ð^N�.s{��H6�+5�\|!�vj̆��A�_1�-S�4��>Ţ��3e��ĭ�M�p��*�_�n���]u�Vp�Q�%�]�xx�|�i��3+q�/��Ī��t���W���Wu�u�kJ�����mׅ-��+z��n�Z���`�/m+�+\��3��Ag>�R!m�������l�1��x���bx�X�c�t�ug<|yз��+�z��5�ǪI諘{�7S����i:��rא�S�V뽽���z-K�l�M^N��eB-N��5�oU���t�G"������aO�"�<��=L9�Zӗ��X�<K�UJ��t���TW�S��j����z�aq1��,��P�+mU�`u{X��-��~P��s�,j�l��	�m�+ޜ�l���g\�ev�a�D��G�*��P(qZ)��U����Z	�����ļ�$8�g�bZ�O�������/ QH�k�5���J�$�_VT�	
�ξ|W�y�L�)X�}����Vq���t���2����x�z��u��d ��vIqd�r3�ztOY�Ð#����5���OdlB4�p%v$�)w,R��9����&yA��kc�l��Gg)�
>�$S3�]�/Jы{*.�A�m�2��$&���jo���[7�m�G���ݶ�B�i�j�;ň��}N��뇞�<X~��)��5��F�pͿ��t)44������_/�� ��E�SF�1+?y�;BT�Qƴ�Fk���*��`�,��x�wG^}� �����yE��7��j�(���}�'^�R�|:�#ex�W1�vF�]�:`˹R.�qn4���=�
��p�� ._���ԝz����RӉ�|迲Q�E(�*���5l�R�یm�;�x���`�B���4g��A"9�:U��FةF(H�l�{|�Ɋ���nd"�2�� ��v�RQf�04gU��0d8��!���q�1���w?j�E�Q�_/����Qugz��+�]X��� %n��0sr���)��{�{��B=T+�����w|�Kk��͖Xز�;�/�Mк����]���D]�PJy3��她M
>ݦD)q�V�~��*���>&�O��wh��N�'���3v�5�����ts�S~y,���N�o�QE6}N�<uB��Il���}y�^�Z��{�jq��Ź�#�J���i��^>�O�	T�;�>GE'ԫE@��:x(I�m�	�Ӯ�3��h2����Y�����(�6���L-�oz[�3�e�Ů�+9�u��H�_0z����i6�d7.��̉�TZ=��k0��5��e�	���U�S���9T���_{��L��m!�˷��{�{���ri����`_�]tEf�3�}!e����L�����g*K�h:��9gukM�]�u�=�k'�M�f Rm�qq�-
�;鬄U��"B��FԮzau����|a�{ v��S"���m����:�Y�A`�9.�:5��eduΫ%k���8
�q#�f��o.�s�;d����1��[�v��c	ߏ/	>G����q:̓ŋʣ��f;�Q�#z5�G�^z3����Yʋ
"F?Ht-Q��udE7~.Y�鍆oc6.����r�)�IOV��ʙm=>���Н�S|�|
����v:j��iZ�m�c��P�/���͑25P�;)C=��{��-��.�0�< ���ZM��IoG.ݗk7�⏄G�g.��?d(	����b���`,��3��3+3�"_w�n�~���a�E?�u���+.���NoQ4�Y� jb�׹;؆������g����{ki/XE^����ȼ�j,幷q%�,��RG����}�Q���7K�6,�x���2�h��a>���ĚXo�ǔ���gN牜v���`Yn�&kSjv��.���jsxhV��C�`�[�܀EbT�S�{���q�rh�ȟ�Mb��;౾Umr�-��=�xy��\�=�u���-�ڜ�m�@���\�X�U��Hx4�o��X��a�tA��j4�}������8�˨��M����Vy��mY0gٛV� �ڊ��.�!`��3[KU]Z��\iP�����8ߟ*�-���VU-���+uY3P��w�M�aA"�o�������P�e�vP#n9�8Q�H��+O�Q[��ٵvr4�17�7فp�	4�3�ѮJu#��j� �_��O�$������s��[�V�3��8�[÷	�q�{%r�XE���O%_�h���)yq=*������U�:%ЇЋܙŗe�$�AOq����S�'!�8�P8�AP�	+b��OJ�����#�����t��f��q����iq�%���dQ�f�+;�\�����dQKx�K��j�>0Y5�j�N�#K��9�C���J�ʌ��̋�K,�9 �"ВD��Y�Qurvd���q2Nou����Z�XکR4��J������28S�b����XJ��صnx��qkk`�˯N��n����/����k�/9�ה�R����C��io�U$;�|���/fZCH��_K��)�a-Y���AZ�Z�R*c��-!}���fu������}�J}���.ڷ6qw��ڽ�Ώ^8 �Ybk�;�h���)��9(Έ�"�in�w[���9��X���귌P�fF{+u����|� �)�w`+W9mf-�qs��#�5C�S��G-�z��e�x�+��.��'[�U`� 1�<L�DS��i��8��"e��ԍ5���(WK���`�$�k�RJ|H�T���3�Q�ep��*����W�*ӑ�F��8�*���@�ڥ��@�"�WR`�q�@\��+����ڱ(>������Z�6�nGKX�M4!Kᴱ\�o3w���p�V���-�Gq������Y={����
$��8[	��Gt����9l�4�k�zM�r��s����^�p����Q,)[��7ѪBaZ�\�BGc62j�TPL�}�.gi|�b�A+j���ebUǴr�5R]и��ڹ��x
x�.5��g�bM���.:✫��7W��g6���J��������G��PtL�7�1�8^�;3���@�w�yw���s�b�jb;���Uu8� �<$S��w��#�e��/�郜p۱\;n=Bs�k�C����7��J�d�jw;�Mk�@3r��<����Ի^e6?j���K�<1�L�QoN���@_`���ΐ)�B\ޮ�vB��Τ�1,��ڽN�Eq��b��F���wS/a�A5��X Wv��ݹnsS-n�,E�C����@a7X7��\us��.�b�wnGI!ﺢ6�u�^}v��6��������O�e)������	P����S�t����.���(��PQ\�^�ξ���76_f�ޞ�F�I�7�o&�cfE�ٜSk1�\�C����ܭ*�4f�ڳ�p&u����a˜�5unc-ca��#�r�! P��ڹU;ָ)��tD��	4ց�:�ٌ�]l|���6�Vo	�]� w�jm�h��c�'Q9c��U8�0��W��������$(�X��ξ�omW4�
|��yM�Fvf�m��b�R�oV�\���fA0I��q|�(�����`So��7{�����B��&�:�A����'�lx��M6�qr��L�*+:�r���I�4#�����ో$&�i'�b�$��f���aAr�N��^n�^�`=�I"��zgVT3B��"=K�wK��(�IH��f��,���]z��fk[�cFŔ��M��sKc�T��6��O��3��k��}��
p��%k�n���!8�U��Z��z��,NQ�iۋ���vv�d4o���ݳڢ���g.�R�A �H�<H�nd�6��QYZ�Y��`֫K�Y��14����B��P\j�����EVѥDt�"",��E��X�*�PDJ�0Em�R+h[h"2��̃��$�Z��nS*���0P�ʕ����@q�UF(��V۫GT�����j*��Q�P��#h�"�%)IR
6Ɣˌӧ31�V���*(���hYK[��L��[[�h��J��(�D�(�TX�`֨�ʊ���
�Db&dmmlh�����Z�AV���ժ��%J��Z���(�(V�QB�Dq3

ԥ�(Qm�LZ�JF�-����6�f3j�"ѥ�5aRf"��Ŗ�`-b��,��meU6�-aU�n����-J��X�PZ��iE
ыZʈ�(fP�l��m�FѺ׾y�\��t���J*e�����x�E��U���p&2��ኛ%Wr�C�b��0�e W $C��g���}_}_[K�}�[sb���?Be�=q�w�q�ˑ��J�a�X4Խ�)S0|�ι�(�')���9J`t�|"���'ҧ�(�FE��=`d�*)���,;��C/y�r~�N�˱���c(#�j��>�[M�E��8%�|����eG��*C/�f]�� ��,��6+j��6i�E�NI��S%�6�=,��\�e�J(t]Cpy"�m��C��W��2ŏx�/�@���Uw\&O�+�͸�r2�Mj\gY�ɼ�����c��AmC_l��+���Z�\�<�U2:=�*�z��^�׻@K��ٚ#j�K}[[I�z�[)�T-�-�鷽[ы���`t4�x+7wF�t=�c�T���s��
�4h_	�n:3e�hdiHŭ�E���!����<�nP�z�w�ZQW#�/%m���H�9���aѝOG�����F��%�TD��ˇ�����>�q9�K-�LS��6�P���SqLG�*!�8�<ٷ&8��&�����J����`�Gۮ��xq����:��#ִ#6�.Y�x>��*n��d~g�~2�$�U���k��KW��k�7%�GVr��ΉoΏM�A+��xN��Jv_uf��Crx�椋��"�}�[���9,�]/�xz՜�ۼWw���j<~�<]��؋'��؝1P�G�P�P�"��GN$r��nS�Y��ءM��((��R��{��-�U����xR1�H,�`�%F�DVʽ�F�R̞�X���0j�3 l@�
��1S��cT��TH�J��Xv�dJ�,���w��Y�k�դ�M|	s7�Y]�{&`��L<,c>mj88?�3Ɲ_Bk,�g��Ѱ�WA	�����GUi7�^��Z�Y���I@��+ Yʊ�)����#E�Z�Y?�T��U���a�#��� *f!���
�oԦ0�/�B�V.+��t|Bu'��s�ܾIvf��7a�v��8���$���].��մ^��\h�o�x�/������Y�\x<�&!j�0x�x�Sq4g�:�����S�\�dk:��<����r{�of,K�{�8�),�f�F�1c�:5���\CF,�p}pH^0W��!�}Ϧ^v?7�����ʭ���3��n���,��4)�?���
n_��4��~\&�x��kֲ�=��C7��JS����u��޿;�䶴���r֚t�B��y���oG*Xs�$O]}y�o5i]�EHd�V����q����p�,�Yhab[�]���#&��T≕z�<<��ŭ8�����-|E�S��<k1֛*P59���$����T���Q����MeL�Kͬ�W�;�^�#S��j�{i�
\n�Z)���@�e~ޖ\h�v��i��J�.*�.Hcu�=�]K#��;�H<�;p���2Ɏ�����z�I{�qrWukiD>ݮ:�Qi�a�4���y�^����Hi�-N葢�E�a�Wy��ݭˑc��`e쨇�QǞte�*g��{boR�f��p��BP)MǍ�*���)��{2_m�R���D:S�!���P�w�S(�ZdlC�踈��k����q$F�"��(/���DX���>�5��v}Y�;=-�PC�w"�8�w��:;X���~S*#;�����)�
Y���]��hv�;�^|[O���̡�-���C���Fc�V��^�Ց
xݗ,����;b�]��cJ辬X�^1ֺTk닿J�p�6�9�"�R0X"���kҚ�i��b5fyr�Ҽ��g�O�z����-MTr��Mո�\樳	0���狎^u�U��"�]�C{�������^�˘��yzi���h�5y/D�*�;�|f*���ԑ=w�U��;�9��^��f�ݣIl�St0u�ùVGr��c�{�ꅛ����;D|49gA�\h�����)��1AS12��#e�(�O4����{_/@3)��h̎�g��¦*ܣC�qy`HNDDO������ٜ3(�3ќ�UMF�O&�Η�(�F�fz�3�ˮ6������b)l��ċ�r��QZ�"��6�������O�v�B�,.�x|M;6L��n)�f�,�,�jIh������Y��2��T{���z���`���"�7���y9��_׉����]r��f{�x��Դ���C�OQT9�y�(�ԕnE5:c
Vfո��.3{j|^6�z�Ҙ@�}:f�.,+�.�R9�|���kv+<9W��!�)jv}�q5r�T+U�a��UJj�$i����LǱ�GUi����	�-Fk��N�ӓx4�T�ַ_.쬱���&��E���<jܒ:����nC(�U���lW37V^�XW��Y�ZV*�{][����K�S�(׭�#r�D+�Q�
���D� s��^T(%�(0�)����.�E,�^7{�kq_���Zu�P���J��#lf46���U^J�-ž���[��K�³:Gy�!���막�8\W��P��ط]wl5�m�'�C�.�t�z�5�)ή`�[o����/gs���m.zZ˚�7�{ДʈD"�B�R�&z���Q���<l�ץ�������Ⱥ���C>u���~�V�Q��S
�'�P��
���hR���w�ԸJ�+�<�{������������(�r/yU�ZR��;n�ȸe��tAGO�́�x�Vͽ�K���Q�T��FM\p�#MCUn%U�iՙ�t�Pr�6 �Ǘ�ʖ+'�`�s|\�)�yZ�
��iОcf+�*�qj����v��W�
W̩���R�r���%.tU"6��ږ�)R��])J�ۣaq~�K�w�׈k��ل��'س�,U*���@��W�S~�)���q��g��+(��^(N�ap*Vu�6�ֶv�cd0v�'�"�3Djïw�I����/|��T��2�`�p3���=�Jc�d0p�@�y�N���p�]�V���p��V�q/�6�	��GzZ���[�V�[�N�<Ϋuf�}S�Pyn>���+þ80A+܈0��`�[kJ�E�3�@=&�4.�C��J���u����xK{�^ݤ��;
�����ӓ#�]��1��z�]�^���O���׭�gHs�%������fӢ��e�ot!�c�\���M��-Y��M�E�����hr &!�.;;���}��UY�j{�=��=��N���GNK&�B�28�n����k��vk�k�WI���&�RN�����]�i
�����m���=KM[��d��ґ�
�j���y@歉�;J0������*�W���l��C�-�J���#|V�2�R��S���ˈ��T��H+�|�^��6[���a���0�!LX51�-�㶥D"�6��K_nVA'�R|�\�[֡�T�f�J.��q�V�<�*(�yU(R,�UO��}����Y�#��S�GeM���vH�[޼q��;�,B1���@�g��͘3���}�6������K�ª5��M����R�9U�΀R�w:����xo�X�z��g���
-����wV2O��L?����y���>�a�ҝ�R~�6z����N{w���o8�Y���W||OR�O��~z5��
�O�Բç���w\�:�=/�����Yz_G�+�� ԩf����ZO��|��T��'U1�uda|G�4#�{��.Y4^�W~�.�z%�{0Q�.��l�L�Ԥ�%�4{��w$�J��Sq�Yɚ*�v�=I�g�u����P�Oգ�MW��Z���p�>���`��ZIt���w�{�v%IM���V�d�1NX�C�;��+����}nk���'�ѭ�Μ1i?,�4�$c<銱W�od+���o�c�9��s���<Y!GOH3	���Q�N�"�Fp�Ptl�	��X;Os���ǩ�K'�Ou�c1娐�W'������m��4<ss�Rk���N�}p`�p�}�V�>vw�$�p�er��(-�-yxo�.O��OH⫵Պ���"IۡObs�,�}��t[>��{��B����v<�i��(�l���g$����4�Q��1\���]1��-!mu=������b�{i���O�h����Kk�^�.#��r1^E'����*���!�m"��,�8:�Ǖ�KnN�lH�6����k��%�����^�9䖦��+zYǁ��Α�G4��y�x��O��p+hخv߼�K"</f��mɺ����J�_�҈�R�=te��L��ȝ�V�ۺ.NY�`���{y͗*:<�]����h��=g����b}Y]n������T}�Buë9ȀXl��m����gR�zZ��de���]o7M�pT��m*��9��Y����]����,Оa7�-1��K��{���q��钔�����������Ñ��F��k��&Nr;ndG7�f�SVacpm.�}"s�W� yĵ�է[Cb>hm#~
�u|�Y�9��F��Y�5����v¯[z�hr�tӎN��MjX��Sf\F/@��p4!O�(�:���T�-�<�e��'�w���guQ�#n��W�X�F�E��#���u<&�.�d�:x�u��ckV��Ӭܾ�
~ܓ�v�u�Un,�r���S�������p5���es)�=g�f2k��*Q2�H��Ƞ#i�d��AN0�J�c%Q�Gbl�7/�w�g�e�0X�K	����pp��i���#�И����s`�Fp��IbF񞊕j��B%���x�+��l6�k�	�z=
��֠��$�LH������s�qP�c2]���	����(��u������IT���j��8̉(P������^D��uI��d��o]�[f��nԵc��ɯ(͆lLi6����w@�����Ge�{�;��8ޚW�Xܞ.-V@.�qV��)d��kU�5�&�ͫq��3����e�4lI,mڂI`moQ���T`�W6���e�x��X��G�v�Rn����um��٤��Y����B�[����/$�[�zl�}K���c����w{Y2�gdU���wm���f���8��T� ��Z��b�;������}��}�[wZE��@���@��*(+�]�㍦���9�\��5F�M.Csy�\B������sr�W�a>�X������-]�F�����]箆��٘����S����E�����:8eT�-9$u��a�s�t�3�����n��-�O��qC����#zD�D(�c���F��5�r��<qB�yoA���wz�|��=���^
�xcc8)3��"yЮ��`�B4�x�.mC�B&�4��zչ����Sz�����eQ+6h��3��<c[��G���'��<��|zo�/_����qyT�[��w��-��{�P�x�tAF��I"l`ʍ���x62��.�y�|N��\2l���fat�V�T֢�j�28
t�Y8h��V��6iRŖ����J��@Gj<-M+��Kʡ;K�zP�r�>�iL͑lj���u��C�4'�S! ��R�E:�X�J6�ʫA��w���|���C��$��$��b,<ʕ+-d��CM��ͼ�Y�i���blR3��_v�xS�.�m־"-�5��#�H/=���=ajͨ�G�������C�@k�.l���R�H�j�����qQ�xҔ��.ҵvN���k彶�[�#F�@�sU'$Ņ"�f�&�<<sb�H���Q`�f�gl]���/ڝ]��m���i��zvCהK$�h�I��g��aړ],����a/Q��J�Y��y1�r1C躍p,�czIr;i�Q�S���ёfk��Rʃ��d�E��$k�.1�V�_���G�5�cb"�g긂���_1��~��v���`�E.���dKiwgr��1��`:;���GM�1B�d k�S*�[��n�M��\��>���x��g� ��J��w
����6�M�'�xM�`�d��&l\<�B<�W���W�ݽ�SՋ�)�α��d���#|m�a�S�h�R���\E>�փ|�gOv�+v-Ju�֗~U����(〷1N�P��:uc�%�#<_����u�����L�ʀ��'�p\={z}��{a���u׳A�1"<v�U P�"��c�t��p��o�6�C���e/>'���n/��Y�������/<����� �7޳�թ˹	>�:��ه�!��]����Ou��ͦ��<�.��5Wa��ci6�`9spd%���C�ᬈ��:���.�Y�E�6u�4�{���Qm[�yד���TJ��]����[P�U�Ƽ��ҍ���u+�S��x3i�f�峍�=,����/����YU%F�K�t1�/����"��eH3�PW��T����� ҞӐ>���N�+#�S*8�;a��v�R隝�fJ]�	��k2��B��\e�Չ���S�r�+�+����N���y���Q![�D�T;���o	�`WpE=�Y��,^"�u�R�n��S��l�ߘ7K�N�؄g'G|^�]�����w�Ё"jcgk�ٙ�_AZ�m��3�&���i���,�P���Y[%��v>�[�u�5�/�,S;!����P[S//���C�z*㲃eAշ���m�ț�oqrWA��6��A:C�F���o�䩮�zr��A�z�y�S����d!!mRo��Ǣ�}0uN;&�Ѹ徖6�Y�0�c\s_Uɑ�k�z��%�gWq/
ט�;|�N��Q�h:��d�&�[��u2�L�V� ���s��%��v{bYT��ݹ�m�������W�n��sޭs���z�ΔR�B�o���_���׀����O��y�V=���Go`<�}t.E�'b�@�Y��Y�Vegj	hs;��c{Z��«�V���(�̗�O��t�B����K�N)�_@^��_)������bu_���)Aݮ���3A��ᄫ���l��~��n���A\���Ggl�!3ʳ�CJ��w����E^s���&�H����tn���L��GW7P�+�V��^s?Yb�q���(�İ��� �*����8J�Dm r��f�[k�wr�FEwS]��ڕKE;��Re�� � gL�t���@� ,r�N���v��Uu7�҂��*ʨ�	�k�
]��P��� 6=�i�ys��I$�.7�B��e؉d�o���%�����������}�S�XmA*;�DzE%h�N�4Vt�09.�?��v�m\׍-1�����#�n݄�U.�D�`tmZr$4�դ�4Ky���}��q��e6�s�v�� YWN]��l�/St��ʘ��љ45"�����gråm�����^ˊP|�.j!̫����7P���P�3Yn�U͛[-�+��5���=ј s�Kr9mf�s�����nHƻۊ�H1f��e@3����ͼ���ym�1�"��BW�r1�2�}�J�W�{��񥾿;!�;���KkV$�vv�fd���Զ�ou\�%��I���-���^[3f�$nΧ�e�kq���qu�5�D��/y�{[y��ݴ�z�*��!�S�:�,u����7v5��sŐdr�5 ή��&Ν.m�b��7�������zZ��絈mE8���R��|[�������{�Β����j�.26�ڊ�j�[mmJ4b��-�/�咵����U�+*�iQ�
�R�R��Ȕ+"2�\�1�����
���b-��Z��T���s*TR��V6�UkJ�f$�jZ�����Xֲ�Tɕ�`�4�b�m*V-ch-\��"kX��qD-�!�4��J��2؎-mf�c�2֨&R���lZ�
��Z����A�TDZ���K�.SM2��mT+V�֗T��Va-ZR���U-�r�+m��-�AKlFUq�iDn\-��nea�RڵQKW2b�qj6�LV���S)U��[*uK��F����0����*c��µ�2�-�[R�ei[p�(�J�Km�ХmFУKJ4̦,K�0C(�([V��q���R���Q��eKҶ��+�Yi�U�,[kը��q��eEPbe�����������n����(�v��4мG{rj!;^��w9�g*���<���G��WG�AYZN%�r���_������i��� �ޅ:I������K�����L�ίo���4c吮����W'�~�)����-z8�،���8#�;P˱S�s(ۋ
-��c��؁)�c{r���&���aT�W���
^�KI/-
�~Z$EW��c�9Q:���Ş����\Q��<����� ץK1^N�XhGD2�t�н�J�Aڥ}��I5Y�}�(�tˆt��SX*Y�l8g	5�R������f*�KN*��α�,�(˛ۮ�3��D=T���t-��t�0Q`��)��g���t�*9f9D�*޾�9�=�7x��	[�/ab��f<�u(ĊUn���3cc*����R8xBn���s�d�ժ�'�7"�F��'K��9C���yN��7&�����T��Պ�=���T�I�';W����38���b���"߶�K+���c�90���e�g$��V�>�~Ny�T��Ao��M>���v���տm2 �K���W��z%��
8zP
6�+����v�y�z�՘U�#�1V��U�l�)���A�@��(���巉!�˥^=��H�Ҋ����4;H](U��9���.8���q:�m_�qr����yb_GGU�ݓ,e2�pcR
�m��+��=!�9��}_x{�O��5��W�|TG�e�3H���[ڈK^��߈V��5
ڬ{��?`����>3�V�t�n4+�:\Ej�q��[��0�sJ���[1nĳ��*4���ؾ�Kxb����H~�$q�S0:��J"��(��Ai���v#�&�%|f�d��n8�C�W�!��xQ��ۥ���|�����thU�ϔ9�BD�ބe�;ZUnh��m�UOr�Yo�(8�é��k����/��ȱ��[�����[SL��;'�k\z�	{�^Te�p�"D��PpBw���J����5A\v�չ��*{=�'hg����x��Ga���<�ԍȆC#F?Huj���n#)�|"[��Wj{����db�S�<=e��=���U[�����7ZdXv혱s�J�X�4jN�w�ַ��7!����� �OV�"�J5�H�݈�M�6!�`6
q�b��l�j!e.v�d掵S0��0z%�ۦ�51p��^9���O��7����:�`t�I��h�F��MY�
����נ5wV6fv��e`W�U��qs�F��4��.���.�>Gү�����`�f5t����ϳ'f�<.����1���Ƥ�u��P�'�=���ή�U��u���k�Ù9��m�V2Rsj�>#OJ�(*=}K��K2�^�ЦH��ʎ#n7�%�g^/��"(�6�����|�`!R�F�B�d6��B~˴s���&a�Đ�nUZ��|�-�9]з2lp�Ұ��2&"��0C��7��	�y�Y�nm��IAԈ�On[N�5:�:�AGC�I.GmQ^i��i�{�݂�W�����1��3�H�N9y��S�zy��B�Nm��R~�(���wc�X���ˊ��֨�-'���\iٳ��s��wrf�S#ng�qC�e�w��R9��lԯ7��U;e�=}(�)�i�X���y�5W�;���Q3���h�WGE͗��n�t�)�����/6!���N3婋�Ih��ܒ:�R1�8�YE�C�&e���N]h�{JV.w*�S/b�P��+�Us�����K�R���ў/���{��V^��������](��>�[1�W�KI~�\+Ǝп��9@���.��\<:�
�݉�I;ݼ���MxAO���;y�;�b�qh��J�uzB���.6�7R�9O�M#��t�A��t���Ӯt�7Q��>7,{�]��������2�r.��mjp��f�0K�}������=��Lz��뱮Pq�s�͟�UY��~�ޠ�W�Z?)?3��u����R�t�wK7P�I��2�O��������5Mw6u�C*���	'�n�1���3�׳��0�ʰ3��w7l�Ӽ�U����d�(K��}�y�T�s)a-j�#�;P\#��Εb����r6"g����W�QQי���]ͤ\�6$Z�`�	xWP|}�h"�FJ6��@.=sx�Hm�3iky���혌B��zE�}Ȉ�u�^%��o��0��-�>��xu��eĜ�$��ƶ]��DIB��P]@`�
%�C�&9��aW��k�ۂ-/���ݼ����ND��j�8d��J�;i�Q	�DkFDڈ7�p�2�җ�� �z�.vg���?LڊX�nL�F��T�����\��ֲ,����6l7�jF�W5%;pg��a��Xȋq��o��˶,^�@�Ɣ������7�)�����=�z��������ʬT�m8�X��ʭ4hZƭ�6'FF��A���=>�ӳFx�GY7I��ރƳ	�&������;�#�U|U^�{{E��$_Dyf�l�1����>\�VK��D�[����O:��O��Se>���jΎ��g~��7^y
9_?U�{��f���r���[�S���yk��>.�&��c�^t�1ϕg��G�n��N�����y�C�C�sۼ�ګSZTC Qt:닾��^�(���t6Fl�P!LX51�y��Rk���n܊����q��3F�qM�Z,��Ɇ��:"��PU�(T��(����|�p-�Tj�b�T�
z!ӎ,m:gV�D�y�j7�Uq��)5���JzG*�uT�<AE���g�Ӥ���t�F��}ac[5L�W��
ϧs��{D�\�)xn����W�Yآq��K�ͱ"\��G�!`�����koG��27���$v8��OS�)���n�^�l�#(��	�ﱉ�\񜋧<n�����+��4� �X�y�ٝ�u!�}OgLF�GC�Q�ʆD�T�
LHXЮ'�S�l��{\�8�~NC�V�fob.�=��<g��Y�l�`+��:V�L�9�͒g�T��xU�El�X��>�-���%$"k@�ה3}�u��"�^A�t�A����"/��8f)���٢�#��3�А���Y�̔��V�EK�֙�l�k0]�����!����X����<��MF\��췷zk��/@��m��瓤V��<ɲ�����B�$����)Π�B�+���Ar1qʼ�X�cySQ1[�n1(��SU\��<��?DV��i�NÙMx��k�U�f�� E���*MyC9I�(dȬ�%����E�k�F�+��Z��]���N�ۆ�Yt
+C�\�����G�����(�� ��t� 7�+L�A"gݴ�T*Y})���`�G�!y,�xjK+�>�:Iˋ)�SCm}������J�xC�� ��-��V7/R\�jk"��(�F�"�;�"���{R��>u��<�;`C٧�%^����Յ{�{���"%V��tD��9}t���~�`.���>�xkk:�U��X�*4���N>Bm��!����p�T��ht;�ֻ���R�<�.yS<�lN8�;�����>�Ӹ̯+������x๞.�d�5+�~�.�ߊQ]1	�j�xaǹ����p��,s�V��>T}C(�h�(.s|'ȱ���l>틌�I�oU-c�76I~��yP�S:e�c���+��S�".�aC,ԊǏӐ��e�#��If	՛\�2[��M��t{��>:����^yv��n������:��jfy�ز�Bhl�j�綆�C@�]D����B���+�U�֓���|x�	�I���X�*���+�,�P��+jŭ�R���9�A�Ѷ� �2ȫ�Bs�rT��!�w,���R'�B��8��N�Y�����J��;�s��R7"@d?���BWVDFz��nS��r��r�ۘ�f�3b�N�
i���-�)R1^�d�=�/=�{{u����a��;�S�k�{ �2����n(�u8��E�-�oRE^{��W='��G�C��0{~K	��\5�>���B4�ʉ+��S�d ����ƽ�g��g���Ǵ=��_�GR��V�b��Ʋmp!|�>7�N�e����Y��LˎU�=����C�b��Z�q�Q�A�0d�'���oJJ��Bq��yON�֪�S�Ѵ�y�Qh��Y₂^�TDׇ:z`_��ݩ��0�I�(͆ncH��#��	Jcg�r�Z����c~͚(�ˋ
����w~{C�	��إb�Ϭ�,S���WV�gv;�ڛW���0h�ʍ�
b�}A��Í��!��ʰ�v�b�;�Yx�r�2�ܜap�:nT�Bʝ5V�6P#���P#\(�w�\�w��l�f�lH��^֩mҡ�9�*�2�+R��	iLv�]e�2�J���w�:ͤn;To+�f
�s�vK��t�h�v�<Q2Ч�� N�m�L����ۻݜln��м�	��n뺋<�໪�J�t_QxZ����-�����E�F0��I���UN`Ujs���y�h���Q��#H@*
��P�ر*h�3��T�˕�b0o�E7���d�Z(���%��!0�wbTgL�E�΅p4"��ڻ�����H�^�ަAR�&g�^�.Ct����m�;�G���%�wʹ�}�>Z��RK}���ֹnmm�]�%tR����ۆeE�C�X�+ȌJY����̋�Y�UpH�]�y�uX���A�
,4$�T8d�<:J냩�'��¬o�f�^�K�Q�c�}@*9Oo"r;\z�p+�T�u:��*"3\1�|�9�`��d~u���O�����(?e���|�^wj��6f�}Ҷ$]*f^��'èL>'Aaq�]�
Q�w/�z�X��}�d�B���B��Ah�y�_�Ix:=Ja����ϩ�/i����x���Y5qyp���8�%�$�!���"�ќ���D��k�/&z�_�2g�"YA�a�ZrwT����Y,�<�f��hڭ��ne�5�\��Yd�w5�ض9^�9(�d��L4.A2��Z��r+Z�Gۍ
�D5�:�N��dÜkHN������$���_^��ӏV���Ԗ��en�=�9���<��QQ��쌫t-@���|t�b�IS�gg"%�"���AZ��aV���x}Y��"�)��&m�㑚=�A��2��nP.�v������>��KR�r��� ��r�
�md>G���U�S�Uo( l���
�`ڬ��@�j�c]1��-M7�_(��ӵ~tA𫘡;:m�Zhд'�[��d�QbKN�WR݋[Ei��:Z�v7�����s�G�U�����G�V�2u-��!�1��"^7�5�h�F Pu���\��U���)G�Cq�C�9��-]vVZ�z���1\��GuiB�GZ��r͛���Z,㞭�x:'�
=w!%����Y�������4 �@��b�ht)�{ڧ^�gV{������/=�~V�`�y�oJ�5�u�S�
� ��t�s��#��.�B^={:�_b�}��5>���Rcn;6�\�0�[*�{S0k_��b:/-h�,��X�����9����Rѣ�@��Ӷ(�1�p|8���vC�����F�O��c���@���W=<$i�ةթ�Ӵ��;oE򧓌W�E-�λ6�N�v_p|��2�0)����^�ʑ=:��a�#5�[V�h,���C)N�'�}��Q���uz��u��Ũ�Eؒ�����(�L�F���'�B�ߖ�>�9��4���̓���8u�C���],��W���2�/
�kҥ��*3AXhWD3t�27q���=J�F��8�����da|n��Ϗ���OS_�R��d�P�L�4��a����/��iX��Ii��*+�mN�R��MC��X(���"1fa����7�V��o ���ѽP4J�k�[g'�p)���xg�m���\o�X�)�']�r�j����Vnʈc���	,����.p�f�*;)0�Κb,law1r$.�+le���|�;P{W�N�sC�؎daʇ� ޅ �"�)]Vs�ܩ@ٷR��D2-�ԧz�^���
$�Qe���n.��8�x�T��� Ϯ4�QZ>"M��gZ���|�F�A�G�t�Q�,�UVGs�g��UƗ�wjx%����)Q��Ow�	�TM���F��ه��4���ƩQ�;-n�H�~����֙���h^����\�����v̮�tk��c#��9Q>��5͡Y��	��L�Z���ۗ���6��Su�k���K(0P�l�e6G^���n�ۜ�!��5�5=i��C�l�V��G��#}XCsxu�2�Y�]�0W9�������^�+q,��:�c�q��"���ݟft���+a�b�X���f�����9Kc����]��29�� /؝N�C	:"��#+*��%1]�v�B�u:T��x�T9��&FE�fh6�6��8����6D-��.n
j���8�qͷ%૖8F���S)��1L�n�3��e���6����Fc$�\��\E���1��1p.��h,�f��5>[2ͪ�z�&���vx �����dW�W�i2/FRc�����6�Z�u.r.w[��Ա;5��2S�J	�__(��r��3���r�4��oT��ǈ|Ou����N4�RƸ=�o_�$�CZ�t��܃$��ޜ4"c�r��V�V%ry[�VQo��f �@A�{�u�,�1���@�aiF��P |Uu3������o�ʉ>�P�ɋmZ#,^���֔�u�#��3�s&j����A*^�2�EtgƑ�]$f\��<�g��C%o.���b��sa��]d�:�u����t�HI��wV"Wm�?@5���S;2�L�>qVT���m����a9��@���Ҽt�Z�a=m0�k6���XR�3ER����T��Z+i�:�sH(ƳHo63k��@N	�	?\����Rk���}����I^�fՖcY���ڷutt��N:4&8h���A�	�vi��ɗ�c$����ʻ�FH��l[m�3*�H�:�R��s)#�(hd�JJ��h#�~����u�lԭ��V���݀�v�M즴]HHռ]�7�����ј� CJ���إJ*l�bs1捻`Z����jI�a`��-�%]k��P0%ٗVKOP�U���.��!}�U�*���<��{[b�-d��J�V�Mm���A��9���-����5^%K1X-���K̺ �]Fh������ò
�4b������J���mea{q��9XjNCzkqJYc�Y�ƺ�=��;��򓣣�l+˽%���p����k ��8�`!;��6m�+A���hٜ����7���o��*�rFW*ᥪ]��T���T.�_5��jɲ�v��>,^�I��Q���$ �mT��M]Yˌ�ˢ�p�k��_W2�:��g��S{]�Dg�����C	ά�L���Tj8j��l��b�g;�2�}VhF�
ױh}�^j��=�K*ٜ�"Us��mG�X�gS&��Ǘ��:�X�D(�
�j�č�m�-Kl�m���q�h�F�T��+��kUDX�����1�`�Z�5rܭe�Kh�Ek+m��+-�D��[QS2���%W���-�[e���0J�iR�j�b�Z��R�UL�0��aF�iE%��)�1mr�Q��Q�h�r�mV[�[j�h�(�q�)�32�KTR��#����Tĸ[kLqk��iQ+F�UKJ��-ƢV��*V�j*��m��&9�+m����J¥b�ʢڣe�(��E�iKlR��ը6���Z�R�(����U-�⡉mhYm�ն6�֥Dh�Vũ[F��B�)R�j��-iT��6�-k\���UTjڶ���Q�S�Ke�DmX������>��Ĝ�q][�do[��.���ff�c��qVY@:��\�{�V�U���^�][���Z��^���2��&��m詶`�Gmn2�: z��-뉍�w+� B݆qH�7�
Ӏ�R����?R�w��R��L��z:Y�*�l����W����ޚ�m�>���Q,wS3@;����BX5�s���y��!Z��W�(8s��Sb��
�M�H������p�����Xu����|%y�����p��ph��mȫ��a�y�UG!Q쇊I�R�yQ�Tg�\F�@ShV�T#qg����|����Z��~����t8'˔5�}�aw���*2�k�N?Ht-Q����6�㓳wy�vum�vHá�����L��+ᒟ<�%��_��8���2,R�a���2�@�<�0K압���'b�T�t����F�(׆A"d�dTm7�:��6��(/e+G_{��Џ=�^�)k�Ab�i6�F�b��ל�h��H���O�n��X�N[om�[�!ýX[8f(J,���Y��(�B�ez�3�ˮ6M8{�lY�*�cLf�涘�XN��$���(Msw�����Ph���88Fl+"�+��ab�N�e$/[Z�n�1�^5e��bQ�%2�sv�֮\�G~�s1t2�r7��!O1�:Z���v���J�l	�A�aw]���9Ǽ�)y��JO�9�8>���O�w�a���q,O�I��ͭ,�l��ڢ%)x`hm��Tꍈ��jM �6^Z�I�<Z����Ι!j�<�Fl�`����ak��S�p�Kkr)���5L�ѬN��w�UD��ɥTmE\":�uLG0k6QQk�4�9�z��)��Q;kl㳾�/x�}�ӆ� ͇����3��b�(�r���#�(�w�o�^D��)��}�s�v~����a롳~r8%oR�e-L]��*z������JFfE�w��V��:4���b�a]�8�O����I�p��:B���+�!D�&x�Vꑺ��kܤ$�O���\t%�@��E�w�%Ћ���L�E8�AЮ�B��^e.��'^�B*���*�n\ۇ��Fȯb��}�r�=�m���U�w�]���6�VH�}���������� �9f."�\��E�x�7�i���zY.���[���̉�b�����Gۼy��&L0��{4I"O�����V�L�-r��|k�
�R�z�@M�I�U��P.S��r�����ܛ�nŚ�to��:E�B���;Qo�>HRx��kh�9�M[+}׸�*R��� (4V�.��ӝC�$$��k� "r����v[��X@��X�Zof�����!����C���Q��8���y|�XK\��B�b7^fXwΩ��-�=ye1�/NEu��a�z������N��BX�f���g�2��((�!c�f.�K��ۮ�$ˊ�9�)�ˑ`�jL5!Kb�M�"���9���J�l=�b�n��FvqP���]�qcDIb�I}�1�Y$4b�ņ�KZl<���Z={/7q�L,�z��^�u?�3��aS�@r�~��C�p��
�^�hs�؁Ow�B+�2�2cFN�s6����m�PdVVݠpp��~_G�F�m�>&��v�C&�7��dWyƠ��Ag���Z�yG'���LP���ҙ���v�)2�(�v��b�7����_t�.j��#	����6�Ui�BО4-�9F�Νz�l�$��t�1���]��������E3Y�y|����6�1����:M����{�t�7��u��\EgH��+�*�U����(〷0�t��mm+�,W��/h�s������=����B�7�t@|��A�����r�ٍ��^�g�͈w
��:�O�B�}u�G���V=����8����σ�.k�o� �k8���mh'W@���ڊe�}z�����s\���[���a_i�[����oR�c��ˋ���q��D#^�8���Q�~�t���Yq���4�g76`hpoi�m�����3/�b��P#��"p0�h4B*i��U���8���:�Ý�&��⁜�+��w=of�3�E3��,����, 2w��pt���룯S����|-�]Z����Z��-c����4��ϫ�[+����.��-%���fx�"��G�2���ʕQ�3��:��{ԗ��gu}�R��*�|���)x;�-%��Ь�~Z&�vl.�L�kF��EFweWd,j2˨��b5R8��):� P�%Q�	�*!��Sܝ5ۍрA�t���ç,�[�k� �R���鉞�
�T��� :\���<M^�g>�o��u��HSz�Ӊ��v�S�T��!(f(`�y��GgY�3y*R��.7t�D_}U}(�_e�8=��x��05���~4��	��ꕪ���8��/���5n5�Cۋ%�c�DWq�9W�������f�:]����t�S�lnM1��Q�:#&�8��2Ou1�4ȡe��O����J�{~�x`u�ɿr��kkN��"N�u>�4�u�VKy�������ܴ[~���ǆu,�ڇyjUy�q�ְu�s�ͺ4�x�>��Q ��s�f�*%b�d�ϐj��J�Yu��<z�R�����QX�U�Ĭ��0F=�o��K+���x;�<4-ާ����nk.V�e'K$���ݪ�n.��9��ǲ��O�A��J��k;]����c��N��D��7�<f�.#zpꬌ[(�M[�Gyα��}o�$�'�KG�f����+j��n�3s��x�J�<n�R���m߾�2�{u�;3��_�%I<�e�,'\��җ�{�<�62�k�F�)S�U�&`v�T�+��Y�����L��S����k������؛��f`�G��O\3bqd���q��@wӫE�Tx�{��!/��L�u
MKE��	�X�yQ�>Z,��x9�z�{VL��4T���[*�oչ�%�]�b�U�w��*����q���;AQ�I�����Ѿ�7�n��u�,W�ؿ�(2%����rs�r��º�{�^/�$���J	�t�^�H@זc�a��8�=&χV�%>x\)�[�8�8g�n���s��OI���p�!UV����M����.����;A���ռM�}+�I��\�:�Ϲt��U۾1�T��Y{�Uwv�X���Wtg<�����juoKZO|S���'���D�/:����٩�u��f�"��wOdǼ���;�x!*�T#�1}�x���x��ʺ1�3$*��]�i��|1�JU��yT��xz��mr�ntk���՞)b͡��Vog�s���'I������4���}\���5�K��ڸnb�o
g�`6ٜ3%`%���,W:5��k�
�Ǣ��w��f΄���I��u�Q4�_��S%���+��ZQ=	:��u[F��J��R\6:\+K^&.�-ū`�Pj���B����
	{�DJR������N50b_a�6��]�!�u#toK}���x����lR5UĻ��&:�C��{f�}.�,=��M����[��S���7#�
P���#���[N�䞘����#�]RQ����Ue��8�5D�"���bݾ�zBKkv+�;*��C��P��]OR��E�+Gx �p�NA�s����j�..�"����o�Q[�CeU�:17�bzh�3Ś���str��/[mM����,��R8�Jo��܆��PT��Kl�(J�KG	�Ve_X�ي	M�;1`�-tT��k�I�R� /�;��oښ�7��p�p* Y��X%_\s�ׂ�i��ެ��M݊jd$�]o�ۨ^wW:���/��Yo��_1�c�^w(��ަ�������jD6�=�B�o/���N"T��7��F,Z��3�C�ݣ~�P��tK�}ˉ���$8C�*�]K=|��cr�0*Y�uH�/���AN��Y���NǶX�ţҺ'�-vK�з6]J��	�ϰ0�l�D��Ըe-S���|�L��u{|�*r�r���״�dU��9^>wyU���u88��C��Ԁ�8l�K�T�\�!g�Uh,mge;�7���!ڻN��Y�mjހ�W{QI�)�0��bu'ir� ���.�hU���+�\_aT�-�Y��m(��T:"��dM�U`�Kؑcԩ�5�,T�hE�;���.Z�}U���#T\?{ؽ齱����@<o�`'z�&��C@��� :ȕ������{T~kޚ&�xG�ȊsJ0�f�^���{��#�0USL�R�ՠ]W�_^��`k����\�BW{����^�U���U��>�2X�%gm;�6S��T��{P�%�Y��ù����$we��C�Ht:m�㑛��ͪ@�t-ϟ9u/5��[4��Q�#�۫5ˬ��B����=u��<!�l��Hp���[�Z�Q�l�i��w�3��+8��7��N}Wl��u�7��Hɳxa�'A��g!�il��[�����;3�\{ ��o��SC�|�;��{�ս'��L�q�T�@<6��}���r�����0dvN�)�3��7�(P͐�Ź��V�Ά����}�g4�XJ��J{սuq��#(>s;:m��ÝKFp�E�w;ow}N���-x �4�b��.�s�ŕY=窆�_�ͱ����>��M�ɳɱ�cάU]VNp�(�G1�ˈ��E���@N�.�\�G�\�;C]Tu��Ksge��ܫ���
,�,	šw��D#�-�k�l�9E�u֋9�=[0�m�u$���6�e���K��c^�6�?��X5�8��4:��B(ӎ�,�g+$d�r��1���gLܮ奬ܫĺ
�2��+�V� �E���)�MxDqT#�;�0�*܆`͙ҔMx�f�/�dG����\�7��7ʅ�])��e�<5�Y��ODC�7tGJ4�T�n�S��Ҏ������r��w�%!=<�*����%�T��9��dڌ5׏4��NMF��`#"��(�ȓ����Hg���2�/
4˗�u�']E0��S�a۫�}��!.�f�,7��>��`�ד�o5��m� �p^Q�6�Yy�P��ķ_�J�[W�eX�Jv\�{P.N�Ǧ�B���W:��y"�Į9�����E�/3��u³���ni��Zuu����v�a�����l���~b�_E�3U�OJW��p�OA;��t0�l����Sر��Q��ɞ���"'Ք���E(�b�P`��G$�m��x��r��q�3:�"a[#�m5��[x�<
y�~5v�xX�z��^�|�Gh��d�̮g*�V��}�����s�l ��xuY���(/m#���!U��6�%o�����w��V��m{UA��)��M&�#7��u�L����ݏ�Z�7|��r�na���ۢ���Bsk�Y&z8��U��J�)�*��P2�
�s]=��/�j�ɉ����se~ޖ\_�W[O�}q}鼄���ii��6�-d�����t�3p�T8�QE�6��x�J��ަuԢ�͑�vE����u|�Ϋ���Zm���)�ЌtM�#.�X8w���\L��yf���b'�ʐ�wM�����퉰5+F]Ip� �J��<pDqz̑�
��<=�f�M\^0���s�q�앍��3r�����l�ӆ��ɕnes�SB�|�H��v�=F�n��]3�Y�P���<��5Ў�egq���:[�������S3>�I��_lM���;&cNJ�@�;���r�oqo%�*֚P�F��9��
�ބTB"����l+f@�9��!A���7�ܼ����<9���Q���5Q3k]�F8
�#�#}��{�MDejp���S�g�m��؏�9f��,9�
�Il8'˔���qs��*��d��޻�[�7Lu(>�L.����P���D�^	Mg�<+)���n,�p��Z׃�F͇�+5��u�z�*���+�szSZm!�6c%$�����.hTi���}������+��?yxJ�8z%�ۦ�j.b�����ݍ�<N��x�q�����."wX��Xf,�gˇ��/;I��k!���ݾn[����7�1�s��m=>�@/Q|@�Z��49S�����Qh�Xe�����-�"���W��ޞ��E(��{���Vl�b��X���Aa*z`[[[�-D��ͽ���Q�%���L%�=�0t�j�-Ɓ�4P7�(��*��K��ha�>���&e�k�݌�xZ���X�A�q49��1�'`���lj�f`������滏'����G�m�z��陷)�Ժ!���Z�
��_}	7�u-\M�}sq���ʲ�����N�*^@5N5o 6�=��̠�M	'��oq}ė� �
�G,�>���(�#�F�n�ˋ�^�E2%�MV5���]v�����z�:�}�f�L�H��[,J��R[��a�63�q�>�jm�]��>�۽��y`�F��A^�EM���Ӽ�������t����#�:��@�^�#XA����B@m�8h
��!�h�(�̷��jC�����2�mPBC�Ҳ���VS��h0jegjRb�hf�(���x�܍�ce뒞m�.�F�9���	bZ���C��)Z��}ǣ����^捉��@��RǕj
Y�j��ؚ�b�ړt�d����[�;݀���}fw$2aB[��%bZ�\�NQ=��ҡJ��qV�E3x�P�7&�M�{I%�[:n�3yl3k6�?1�JAܙ諧E5�9����Z ��U��g���x�õ���SY��T�#F����q�Ej;�j�Ǐ&�W���k*N��|��[�ȡV�D�B�,S:��ʝHpE�,��tlN�U�9�KV�!Kό��5՜=K:O]���S�>�,�ak��\�����q�*�h�Yz��#@k����Y��Z���Ug�P'{�B:?�p4�^U�2�ay;�NU,�0m,���(t�gT�W\�SG1��޺=u��S2�U��r�vE�������/��z�����<f�ݬ�'.�ʈ�k@6��	5��(X�M:�F�wN���BBG-�m�Luާ
l�6YV��B�'�����֍m��)$ei��2�^"�X RK��%��Wv����PՉyd%X��y��Cb�,kM��+ow�vF1��N��ҬUà�`��N�\��gm���ܡz(H4-�R  �N5gV,V��eĶ��iⵟi	�ҫ���&��!�dC5�kQ.�U��	G8�=�I�4)
�{�u�������*~�Вӥ��0�x&]��.U�fT�n�u�D�����Yz70�������{%��u��8�]1�:'�y�ӫ:䬥|ʮQr���M�Qr,��*�%��VHU��.����z��e"���F��[�>�}YJ�S��"�����pdc��P��h���t;��oUN;3�Փ��X{�-�>z7X��>�p
�Xb;(.�It�,��\��<����mV.��5��G�v����)d�d0<4!/��mR2P�,�(�+�跋�ƤZ;u �La㥽���cUJꗅGn5ˉ�\=�+6\u9�v7.ǰV���3r�ÖX�B�_�D�-o�b�dR�V�X��R��*Z�-eQE+dF��+h�R�Ĩ#1m�6�Aj�6�+m����+*KV�J�JUD��m�%e`�J1��*��U*(ڲ�J֥���XQR�֢�UV�-�\˅*QmZ��ێ*	���-�f�++(���V��\���+Z1�r�r�l�QU�\���+mb[U���
�Q�Q��J[Eb5�m��j(6Qm�ڎ0��jV��¥Q�D�(�[J���\LPf5��m*��j--
�"���5s*�m����AAU3(e�(�[,QjYj�%ZUs2c1��kA��[`��"6�s&d�DX�Ֆ�r�E�*-J�R��YiU�EA�JZ�*$e*��m��V��R�J�KR�jTQ���b,LJ+����F��
� ����d]�/�u�#���f��F"� ��<�������*S�#}P��f4;VdT�0͹�ˍ#
���]g8r�^��w���h�>��z�;��x�q��X��B:>��$[�}�j��U�`�,W���u��d�1	�-Nϭ��
h\ GP)�u�b����X�%��1����̕~�Sg�����?m<�zAg��S	҄�KG����p$�X��'���{3�a.��eJ�c.�=C�h�α���O��ɋ�LK �E�]r:���M�g,r�F�ˈV6E�hb�p��,��)���=�=�Dz�!�z>�ED��=���?f7����^S���U�]�W ��a��v��y����G�/n�6�]*x��G�T*0O(B����ۆs{��Qg�� �����cb�$��1|�̋�Y�肍�I"J;f	E���ּ|vy!�=�vzz�[���u��9Ʈ���d�8G�����|%u%.TF�\1�����6�Os������cg:.�*BzQ˪�m�{.�3�d k!��r��j�����.�F���F]ʻ��j�Q�;�N�R��T=B��[0\�c�8�(�ܕ��=-z ;��9ϵ�"E�=�z�^]��)Kt�]��M ���wл�؇r�RE���Uݹ�r�
�*i��#�ԝ�^hŽi��U����q���́�{�κCed�(�"lN\,��f��1R����C>�b ]{��k��=y Cpڗl�+�����a�KE�ʊx������%
�%�H`�a�CF.LDY:{��$�pbe��0�#at�g�1y�Un�*|^�ϼn�=R���`%˂�/f�~�>��8x��@��Xk.�2t�6�����H���g�ג��knh4}ڧ���]���m����U�۳~�,h~u��,dr��9��b/R���I>���5���kʵH _Ff@��V��9�˺��bv8��Y����'.54X��Y�zo�^9����O�%k#�(��E��cxC*�l=T6aU���VE��P��^-QH�ɋ�=�6���^��ƶYq�"�U<R��e�X�Ƀ|�jY�&��P�5���l*0�1`�sL��>'���>M<;�=0e0�u�e�֦�]�b���Y��G����4�<�P
�)��ع�<3����gRS�ש��f͋�<%3ۓۼE��"59�Nr�yt�z��-��@y�FZ{����ȏ�Q�'����iB$V�[��}��mj譳otZ��ݥ������^'ð#6��Ν׀���tZ�s�3:Z:n���W��֙l�1�H,�@�dB�$�GQ��*���<�ʧMm]�V�EB�(�b�D�}�.b�)��)�:����M�2��G�ʗ[�{��c�5�Jk��K��g�;���H�SvC�gm�肱���f�B�u��w���]aY�\����+Al�9�]g>�|є�xQ�ח��22O%Q���V�\�9b��Ю��#e���)��Y_Ut|>	�`�*Y�gK���6��g'������u�i�zC�]�%��Fzd�P%Epf'Paɽ���.�6�Z�c��LP2^��E{����"aeAf�5��[g#\
��<ju�^뼄��~�u#\��)��𹊻W
���*�dlT�P�DSFp�>�0w�,�P���L���t��橈.�wt��
�!�#���V*�k�����*/ό��\(�*Y}�g��2��<���z�����k6Qb�p�MtY}�hf�.��8�h�j��V�Q𥞝�uw�y�U�U��}�B�n��p�c�-�Wm�tΜ�k��[Yڞ��zǅ J��ٝY��&�����Ƅ�Z��%_e���ݺc�%����e,J�)�$���;ZuFwL�ne�aQ����..�8�6�d��w,98���q��Ӕe�#�`����uO5��Pux�x�Uy�ˉ�#5�2��,�=����y�t^Y�n��Փ8�E����ӥ�ׄ��ڊ(��t��G�g���ѓVRSҢ��TV]g9�E���ζbñ,�*0螚�1�O�!�fn*Q(�DW+��Uf!�)��Qsʙ�9�؛�V��Ye�9"3x�3�й�8��
.����Ӆ��,�ގ61��h�.�u�z��Q���p�F��J��q����Y�ȗ�����֍�cGS<~�T�EX��d2�7uQ3���6�� "�̸�^��҄`wCX�����w��<�5����uҒ�pO�(2�����0;�τTw���fhތȬwOw��BH~{��t�ź�|�H<��p�J��>�ΗU��P_i�u�SNau��a@��5�E�^+���p5�t�t��c�N�\�^�$N���Ol�c6����3/��m5�*��q�b��l�	Tj�D��G����Y��;]���R����}���of��S�wL<F%.��#V1�����l����(D�[Օwk4��
�Y��-��u�[�zo�u*�WF8�n%�U���tg��e�e>�ӡ9��t���7X���]ӣ��j};S;*Na����LFsNlh��T�3�ax3�����{K�L�v�>ݼ[�b��`�S�v%C�0���LH���>�l�s�pDWX>b�����z�q�LTT<M=>�8�NS�}��ꕊǇ�yI-.�"���D
�J�jIn6�n�L���^��>��Xo���'�]�����Ĕl"�M������{�h��)�7�����i__���5Wv��&�ͫq�Qe���@�0tf�*VglD��n����c�dL�cd'o��z`���v\�|2}�bjv}t���(q���L��f�wo^k�wWkaD3}:��;����WE�t6]Q���EdFěL�gsP�22���6�sr�+/��H�<�aN-�Qt�2�vF?g]uШ)��Z��P�6�^eVf淅�E�LN�6�Y�
!h�x�⥐��Isc�F7"\p鞈:�Y��;=�n3�!YBaЬ��ϧ7�/)���)���;y�	ض'����(Q�[��亍L5��b�oVw7%{���T+'�8�g�go)�]�*X�z��tC�l	d����{5�u��ei�"�'{�fm^� cyX ��od�LA�6�@�o.�̣$6X���}f��;dJ��Ҕg�R�^��B���Y�ֽaߣ��Y��w��3K�+L��O�ᔼ�f�,�w�6���ձ��}��FeN�E�F'�肎!�(혯D"��=Uצz���=^���F�+��������ʰ3����1��L*���|h�u:�x���qA����s=��$��i�-�U:S��h��T<���8%
�C��8�����yե�ۺ�(��Q�(�=*���yq��ņ
�7&(��M��ےUH�����$m�����L�͉p#+j�X6Y��$��E�=!��D�H����fؾ�o���������=^��^�U�K�֘ϼlXC��ƈ����_f0��|p��i�u�d�p�mZ��)��_�e�^-.�+mw	�s�ʟtZ�Q��.�ʨ�o^�x;vl�{�, ]y�X���o����M��P�ݯ�VF�F�YS6��8���N�z��vΝ�t4��=��.�,���~�Chf�����k��E��Y@D�_��a�k�rJXᓺ��s/��쬖���0>���ʛ�s��/:�s�q`M�z��]�Mh,�p}��9�ҍ*�V5��f�T�ܬ5{��};3*���V��� F9�#\{���xg*������4�V�,yu�> (lw\��)�r9¬�z�lū��j�ٶlz��;��#�n�&�Z��=�."��"ʰ�aV�/ .R�;f[�;���ak�}�ܚVyWJ�[�����1`И�lO�D#bu�8e�<-��D��k����S[�R���8_�ӽ�Zc�$��E
E�@�*E9��*�!������k�>]��Pż���d���8s�[
)�tAf�`�2!N�hDqG�:�
7W��Ft���;ڙPl�~���;(��m��s��|��<����=K	t��Y�ys�b@%O{loo���Er:9���	�8�u}�|�|�
�����&D��Z���ڼ��b���>X�++����Ьt5��|���8\Ń*�1t��<�9Zw�a�|� r���ZO�-�hN��F�lR���gLGKem�%�ŕ��+]!pmi�`KW�u7^���	����)h^�"�\�Qyaǀ�d�����5;' �f�TS��O.��4U/�J��A�k0����Y;�+�>��	,3�P���l��t��tY���<�GKxNML�:��|(�#+9ݒ���f,Ķ�}�ٍm�E+�7��C�(Gu�����ۏ ��֛�X5�����6d:��)��6�����u����H��ɽY-�DBƜ�d�v+�:�z����Ғ�9�U?9�I�
��k�]��.9�]1�0�ra� ����Ie���3�*��C�!�d�v&l�M��p��Fv���+)q���qۉb7cc�QY���-u���Ν��ك�����٧GEH�B���^O(g%�U�֜�@�e�3g$��vM����8���3�K�nko�g;���Q����1"��7�(���ކ\ ��{L��Q��l����&�-�u��ڮ謇��m���2�&:���r��F�q��ȱ���ޮ��U���DY~K���s�S�L����M�zk\�"���&`tx���Q��k6;{���(@���R���q��A��-�������(�����$����̡�99WGBC���C9Ȇ2FL`�L�t%B�b�x���Z�v�Y�^'�ᔋ:5��Q����9��������3\&��o��T ��򾞥]:��L�g�A��c eވ2��:{P�+�����n\s�D&�^��W>��9yi!��ॻ�	;����Q�u��܆u�A-R�T�PL4+A*8�FC�nʖoK�-F��1�����0�R����h�ReZ��V]Κ�="���q�g˵�2�-P��sQ��+��w�{�7lS9#It��\�mU��+��ρ+���`5�Mi��\5�|*}l�2&��5gp�sX��6��~���K��>����a]=h�#���P`�KI�xj>�N�;������&�稱��8��0���`�X�ٜ3%`ȕ����4BȺ�/_
�C:�Fqt���յ�2"�N�2)<�lÇ�$�]���b�_��1^jc"b*���s�������@�g9*�mF��Xܚ(_�p�^��DM%OL�9�7w�W8K!_BɈ�ږ"m�����R8)}��\���]\�e��R��3mޣp�:�闸^�	�C\7Ӹӹk�"4׻z�?{�ؼIոʍ��\2:��(p���ͬ*E��]R�n��Z�G!��c�r�/���n�g*�gM�鬇1�vءƻH>|���Z�4(���[�w��q+��V����eCT��� 8��p�*��T�ov̝K�k50��v� ��`!�ܠ0wL�"��� ����;�3���M;ս�M�Y�g�����^mN����4t�%#�vi��{Ԥ�'�>���bU�C��Z:�ŁU�Z�]ϝ���7y�'��y��
�M�tʩ��\М��6^�:h[�GVKF0���x����2T%��2Cwe�}S7������w(�|�1u���7���(���U�͖Io���'v%A�.q�B�1��+\��yN�ed���r�Z�:3��<g#���v��`i��WD�dWRM�%ʧ)�\��E7�G�iZNwƻ<����d|N�;���9��v�2"ծ�q\�k޼����r�sFEe����<hcH��قQt:B&�+�+ؾ�[����:�̎������SN�jLf�w�
�??��#��u,%�TD7��^�� �����-:!C�:�:�ft���b����C��m�lH�)f12�E���3xg{;^U+�r1��0D(s��Qn �q�LPxR,�Tڃ99Ů�{�Ӟ�/�')+9Ja��Z05ʊv�B�(�}����=� �d�k4�p����c/��Gfl�JS]����u��(������/��ف8l&�
��J�l%QYw��;T����x[�o��N��}�{�{h�A�g.�w5��&qV<�CJ�ÊU�YYNv�\�K(/$"��#32:���ƫ����E��0c��Ĉ�}l6���6d�'����)�n�Q�R�ǎ��i��;SF�ǌ��.0����c8�{�-Mc����uƱ�R�c�w�pf]5�	�k��#���vAE�`q^� ʫ�cx�ɉf�y'�;dF�"��i_H�5Ց>N�ZzE�α�o���u=޲��ƽ�*T�*v�^�YxS+H�d�V�;��ü�.C�%k��pvI�Z� zV1�����{��v�e�;ռƴi�Q�ďc�M��z\�v�9S2�k���yjB�Q��seD�v4WG3�rx���ۑ��֬��m`'1ڵ˻���L� �ڶ˹0�F�P��a�M��|��U:��tFUƆvv`1|.�w
Ŗ��\�N��=�q��K���GT|*���f	�\Ɩ�; :�T���L@և%M�O�:�=�.�'�m����&1v����3pp�ٽ�0�ui��ʲ,�q8��wQ�z�Lɪ^n��u��$��3}3E��gY=
fㄥ���5�hf���8�.Һn�*�ح9uلe�SnYu:�/���w6�C�wY���2��u[�(c�U�[</1R��T�ڛ�%;�͋�U��{��ZO�`c��,��-���Fo*��Uixc�1��4��hv�OA�P�y������wSp-����Bl�²+S;c�I,�wv&Q;n�8a����eV	ծ6��z�Mn�p�m�,$���˩�f��$�4��/��^��dh��B�A����:�jl������fօ����M�Q+��z݌�YS��k��ֶ!wzv΢7�g%R�q����L�S�R�+p��)e��t����|n��[�ҷ�Cjh3MA�&^pK-ży��I��`Y/2�յ����J����	V*���
�ҙ����7eL�C*�8�l��eYo2�`�����	X>9�m��kaI�J#sn��(�p٥-[���ǘ Ǫ�\�L���P2yV�z�U��v��6���l#��sm��}�t�B�oK�u:ʻ{%v��wP�\�v�仦;M��<-T�r���u�ՀӭP���������,�.�J����z-�9݇_j�۝s�A�����ĕ��4��`�ܗ�9���3X"��fN�3����b��ɻǑ-T;��4���f<U�{Ԧ[��ͮ��JD| �Pm�*��f*��*�k(�iJ[-3+���m�6�(�bc1���*�e+�ih��p���j-��Kh�s&V�[[m�ij�A\s11�r�̢�YQEE
�kYq1�
Զ�&P�j���QAQb��X���R,G�J1�a��"�(�(��Z��A2��-\l�q���mAAԮ�cE����ks0�˂��GA�*������pm��TY�U〥��"(��.(�1-\�V#PXVB���11��q��n8Z�E��F�ۙE��5��5�e�F����˙b�����2eDX�a����Ub���j*-)QG-B�㊁W32[(Ȃ��**�ceC���5(����m��EDV���V��V�LTX�!��(*[Q1��\*PQkV �-���*�_Mt:����p̫����ݨ�E��Q\w0Ur�f�x����%���ԭ/�&�!�d�[�W��Qm��\���B�	#��9&RN�2yI��H��B���j;���ED�=�&z��׾y֮�����4\KYpE�'J��qAc��2�2,S�'�h��=�w1����WP������q�%vy�xر�j ��D�����\��6G-�%R��h��|,i�e�{U�p9��9�y媸����-���5�
�uK��?tY�!V��]�tZ�f�$��ґ�W!�>x8���z�wTԉ�ݑ��x�L�1C���|�30��Þ��q���#��3M1θ�55�]�1���V��lSK�$S�ћӣպ�Uҹ�J�]:��Q���qV���qߵ�5�Y�圫�	Ϳa^IF{��޹|,~�cGU���66�:�ʥ�U�-xN��t�="�Mf��<�V�mC]H�I�m�
t�b��1a�,�,D)D��G)�^ڧ
�˵���m�ǘ��c��=joT��=��nEDSs���o��Rа��9�]fycepTx��:�Е���*s�z��:t�H*��b�di&�n
گv��h�=6�_06q�O4-���e��y]��8��x7��i��ף]ub�Omط"ri�������Wbޥ�G�^���-M��
�V�`<�w��k���}�ۦ�
�֍��85(�Lo\�29>���jv��2=����L:ǆ#�F32�-��Z�jWst�|�4�δ���5b��&ߍz�}�p��`�x�xpT�+Al�����:p�^>��X�Ʈ�w�O]��5����>�	ץ{��>����hs����|*�3�&�k���w��בE|2:��p�l x��t���U֖�N�*�u2xS�+8%K��8�K�����)�g��/��&4�Y�	��1^td�v�V���d,�4��'��]��U���*�7�٢��=���JȊm�i��0Y��:P�ٕ+C�Ǖܫ�h�f���=���O�g�lW�֯�V۫����0�E�3��s��sV+y�"��+lUag1NR�f�,_�p�M{�p����^Y/6a�D��8����4m����G%m;
�ˋ�QE���;AK^9xx��>���(��n�b��Zm���8�};�)���;T��@��N�:oz\C8���+l�*M�r�G�=B��<��f�e��M���Â�al.)a�ٌV��C[ݻ��Ǧ��b1$g@:֛�����_���(�ts�7�a�5��f9[9E&s`�.��wK���8�J��z�Lߕ�\�#�8�D��>�TY������io9�޹n�猌nz"}},��A�\�gB�܉iR2�wE�7�BQ�s�Bʸ����|�ܗֽ�Ǜy�a"�Ы¼�8tls�j�P�z�W��!��d��{hs<���Ĳ�-��òZ5��׳��B;���/PSs��u\k�*�&58���嗜��E�+���=����d�<�'��
�T�Â.�l�E{P|sޛ���	�^>d<<7�p{F>U�O�+P�ӥ��ux,�K3}:Y�[jf���Ok�0���U�_-d_�N.��b�}�R��p�!^�K �U����[5�� >	t�ud���|f�&%�/�1�b�4=�����x�M��/��C�b�����_j�zn��*�3~��Q���&wy�i�^l���Y�2����f�b�v=��/��U�S��m�ւ�R��p�	�!B��
�'Y�FD�:���y
�^��N���n���0�79P�,w��ٚ���f\�u�Cm�i�G_3Js��i�&��"u��N<0��ݎ�z�"�m2e��u�N�̒��Tısim��C7���X�v��捏�m�
��+�8�m�i���!���������WVg+�/��2�bT�t'��ǖ���`��>@>ْ'u��SB���ɵ[%X��z��K�b��k�q�'܉+�a�����#��T.�In+ٳG���e̥��e*�@����������(ڷ�z��^�o�l ��^9�"ǅ"z�1v�Fp��Z�}�]]Z��[\\L�z�2�y�Va>��Ч�S�7�l����C�#\��E }�������]AchS;�#tW]�g��i�駊�J�7�����]��r��,��O+�M2�Y;��h\�\l8$u�F3��M��x��L�.����O�b�Hy� ��e����%M&x�V��D+"�5�R�xk���E��*:�۵�����6�+뺌Q7̸�B# R'A�v��8td�|%7���x1K�ˬ�Ym��K���I�9U$���d��¿tN��;�\���hR�&�,���7���XJ�f_fwz.���+zM 1�~����2�N: �@bH��يך���z�z��U�;�׶ R�B�R���M��I�}��o�:�{��ڣ�x:� ��j��Wc2���P��ծ�<Rs��Kv.��Uw����e(��V��2�8^��y:�Jٛ\�gnRT��RqBNRq9����6�����D�a���]�F[f�ȿ,Ĺ�6�����F))^T\�����}B����{+5�#ד�.��Cb+�҈��U��<�J��[�Q����ï�9PF�,���g�
6b�p�XɣW���LHz�`��5�C���0����7S�%���0��-\身O��X�|t/zIy- m-���ռ9n@�q���H�1rc<ԃ!�6�5�͉�͛���..��}�Oʭ��$�{��[(�b�>����DcFE�������u�)c�?f��e5�9.K0��|�<��ˬ��Ȩ�E�m;�6��D�b	��a}��[k!��r:{�E�ܦ�����gB8^R(f�`�	���U8lj�|�}�:f��E��W2�;�yD����8��Un��0Kg��jsi�l�H¨�X;2�f�k���l� ��7�L���R�m
��91N3ճF��6��e�^ޑe_��+=mvEIU�~3RgY�R	̢�q��vԲ��R�c�y{ځ�9;�S��P�Y��MZ�����*9���D�`�,���_J�����xC@��㆖>�"�f�B�w8u�:r�9�:�>z+/���֣bs���C��8ɼ�y;8�Iw|���Զ��Џ{{�:\�=o�c���':�S�8:����n�
h���.Н5}.!嘳����wU��)�G�)NV�z6ra�s�(B�*���"��(�45+��F��)��uY[��}��QcT��k�D���k�\e�QH������gЧI�b���*C�<�ɕn3�/���#�~nz�wS0k_��h##4F#���x���n�VEu��ν���4r�h�g�gw�%!&tp�y�!fQ;v���!�X*!�k"Y�/ii-r�b/-U\)�6;(�l�aU:�z1hc5)����nZ���U=c.{G��4-@/��u�ާ��G��^:P�/����ƺ�ɼ3��]+�N�\��0��#�c���6IBT��BhV�7�	����9��dHxZ쪕��[�i�ۮ��d�;p��
���{��FR�
'�#�)NCw�4;tt��!sݾ�.���X��z�ؒ��\N�*M(g")�8e����,W�f�|��>�+:��=���ˣ͊��т�w�h:�Q�y߉yrc�:�Y�xrv�&Wo)���<)1z'f%H���������w�K���,N/"ᒉ�ם�&���;5��L��RPy��ubw����?Q�º�mG�v��m�� ?U�
֎Cc=�nQ�%���ܣ�|��W|�_�������k�]{�U��:�k���wz�Ϣ*_/WrѶ�u�&W�����.b��;Yu���e��ˌ�]՜���"��T�>�q����M�;~�d
��Pf�$�(�N�:e<d���{!z�'N'O=�=�%��޷j�H�m�|q�3aء���b:�K���bN�a��L%���w�ƎQ��:����c��v�"�yR�l7U��*F]IQ�B�,�Vj�2�D{���k��6s��bg���#�J�B��k�z��s��3�"�DF��:7)MŞ��F��de��t'A�S�,L��	������[�+a� -��8�m�M��+w���z�;���J��UD��+UwS���d���+����q8͌\���k͔7�4|Ϻn�~���z�{�]�^���
__�T��n;&Q��'����Ճ�,�b;kp������G�u��&E؍B�7U��R��g���㦍`{�4�^��p����.z��X�Ե�q�aE��aۥy��]d	t��q�s���᫤�n��ή߰*38m�\�I�ܒ��i�n����p�r��NQ)5uC�8k닿L�n-���S�24R�b��v��34*8��H�j�u��=������c�t�0c��v[�xC��l�ׅ*f*U�Yt��q2:�m���9%���_�����Y���T�����Aǳ�bf�w��;_<O3�R�!#D����U(����ղ��,EyA#S,r����똻�Y�s��(�D��"P���h�qn,Q��R�rh��,��Iv�������<�(j�=��"w'��~M���yFoID�K0}r�R�In+6h�>=��A��L�ͤ�R�S�8��eTV ��)���kTS�b��V�=Gp�W{Kuuz�0}�l�W�;��#��ԣc6Yq~Wx]�!�4����[�Xv�b�PF�=�jl�.k{5��6�E�X#TtWfgry�8駎�M���F�3[��R��.쬱��������,д'�x[�GP�J"�@v��(�Tc�pB��lz!r36j�X ��N��C���C7O=ҹv��{N���s����'-�r*Ȟ`�|,\��

��^��3�����ؓZ���it.�v��qM�V�Bي�����&n�ֺ��}�Q�v��i��[�L���,�R�De��gs�T�fr�^��-+Xi��c��b���<Q�[�hM�Q
(څP�U�df�
���Y����=N-!�R�j�p�*�v�gb�
D�$�E������:%�.�Q�8wvU�7g7�v.��9Q2��S��q�V���:��hR�m����K��+�/�dr+����{�z��6�V��"(gu3�m��.�肍bH�v�i�Z�d�23���nX��7Td�=!uԏT<���ouVT+N�ȗ,ƹ�q8-]��1�S2a����DFp�/��X�3ƶ�X���B"[��m�{)a��콱qOm�h�m%��P���"�/,Eб�}b2���)Cq�!:�Wu]�i�XE�koܭt�V��4�9�I;Ip��S��c>\��e�|�P�W�a�Y�����6��']���*���M�UۂWJ���Ӫ'%�O�/��������J^w'��7m�:zϾ�j�v�2Bqqёf_LƲ��2t����������}�l���{]Xwb�=��0]�=��H�l�眮�m6������"u�~���tUv�i/80��QHk�.��onrcP��)J[k��u�;L5��;���st��|u�ٷ��[�
J�w ��7�7zw+��,������i�T���`�+ �qF�s�pٳF��`���^��@Zж5^�^M͵��[v|��sφ�b�l� &zE8	L����b�
��K�����S��N"x�{�Ui�n8�`��$�'JF$�����`#:�^D%�L|tY]���k�s*Z�^?-$Z/���aͥ�x�u���Q�D�(O.sk����8�S�l7)G�Ɋv��(a�DD�8�Z�����o��V#YF\���n�U��X�(ټJ�qҋ+�v�bƩ�X�Wzd��"���lv$tu^&�o6�bGt(�/T���I޼Q�]q���5�,��Cی�rq^�^5�'v���C*��z|!V��;nu@x���"@X�\E���QL����C���$3u;�y.C����XZ,ς������N8ʾ�)
�vf*��\�o�Ys���
"�,_��'�K�D�pT�+>�R�TY^���Hc��HUN�F�.&\AW`��m[t//�L��m:��h|�u�}����N�u�x��e��m��۹nrG��Q��8�fpk�����Y�U7��Ȧf�$NNV�����H{ 4�Dg�c��Q�#6b���uvA\2��t�yZxZ���3k����&n�w6�M�܅ڦG�*�&��r�nc���T��d<R��w=0iY*�StA7vv|�ޖ�9 �p�N�m��©`WY�����h�$�e�vic��R}�y��ث�(��Xl;^ȍ�Xtu	|���t���(-IZ�-�;�u'%��]�[g�S�,FM����;�Zﱵy��@;�4����ȥvorT�CJ
�j��9��̈́G�����&C��s��x
�-j�xdUÌ(��h�[O�뫏B�tQ����i���/���ZX;uN��b�أ9+g���L�U��|�ټnw;D��ڙʋ����B�IB�x����N� �v�-��oi[�d	�e=zU���N�F�e��v���t���ΐ��f�nX�d����?Tx@��� KRjR)B��x��Y��&��i$�+8̖�#�z(ޅ�0�U���J�^`�}y��X��*$��iX�����]�}�� }�Z���C��Y���aeU��B���1SÕ����f���M�Ψl1+�ԆM���j�}p�z���v1J�6F��F),�;zut���}�[�:j�]���o�1qlG�8��jQ��x ��j�y-��27�_e��y�I��n�X�����|%�9�)��{v�j�r�tю_0���v��+�q��,*@�ut�+�(��z �mt;m��-Cq6y��W�a���n�h�h��V ԍ-L�m�m>IX3�Nx�C��Z\�+G���gRϭ��V�C�m���ۍ�K��-���*:���ų�:j�
�R�]���:
�e��0�
���๓0��� 吧,ȭ��/8�d���}�\A5���}��wn�Aw@˻U�k�N��O���󣂃������0�nns� �.��"B�n����N^�ԝ��&�7��3�z��Vt�S�@�L��+{��ɕ��k=��,G������9o`���ʥ�M5F���4�2�Eh��Aμ��nvkr�)B�kE���6U���:Ju���v�L��C���d�x>�5��c<+_y|�0�&���z�v��ΑP{y���D�]j�=���4�&#����Ue��<�v.�H��?`mgK3X�rÖ\�͑��]c9��6ؒ�O{/�D�q:��K+�d�7��6Ndm�u'�����n���$�IN���I����f���L.�����y������Ԫ�B���+Efe1cs0r�#�32�Sb*�J��j�S�0�V�ܹ���2�--���b��Qƪ�cXc
�
�؍˂�T����)Z��l�R��J�0�L̮UF8��ij���eEb"�VT��Eʸ����f88�AD�cF+iR��؊� ҃��K�QD*y�kEG5��2�B��f�ٖ\(������@ƥ�0e��̷.0����]f,DiVUt�f��j2:�c+YmEERc��Y���k5�Uʈ"%�����T��V�((�E�e5n��[JU+�f:�0����,WHi4�4�\���I�c���Te�U�)WC��LMj鈚�m�Z��麵Y-����SH%�Z�ar�8�mX��0uh��:���:sVZ�j,���ҥ��9r�Uf\��2Ɣ"��ue5hԚ�m--��-���:�¢�V��c
�c��mZ�#1�5i���˦��pTeh��fIQ�k-��]c�Ľ68�Q͎��ַp ��L��P면�f��v���;r���)b�^=}o�:r�e.�Uu����豾|[�G:��.�*	z��h�}uds3A4%D2�Jc"�9�B�Q���J;I�ɝ���զԓ������e�J��`�xK�:g����-8�>���n�ctD�2��ݎo�7��/%Q�K����U��A��,Jsg3�ޔE.�G��ku��ȋ� ���ͻQwŬ�|i��n�&:���'�E�����Ӿ�S�ϲۙ�z�뙳��CzӦv�X;��1C��Gc�~I�D+P�ۊk6o�T�<}h����ݡ��i��ng:3i���ll2�F�Iދ/���^
�o�Y�9)L9���og��m�G��{2��\����7Zlf�Lz�r�j6�?nt��%��J�ڒR=��,�8�wbS�9�5�#fC91$ F:Os���lo=�ֳ2�b8.��D_�C.����gHàrm�<�̺/:J�,OM`��N�[7�mo)Ɯ���!��O��з]C:Yǁ�E�t��
gr&�JћwE�2)��7tg�_�>S�rGҝ�2�&)��ܽ�k_Jۃ��r�j�nmt���o*2�+(Z�J�]99ǜk[��Y��+�.��x|F�������T1�œ�XE'iS�ΕE�WS�m�]n7mwnv>���
����tս��;���C�.|��8u��ɮv\�r�<�]X��]��8ȗƅkb.8��� 9s��S>/vB��g�����Ua� ��*Dp9YȄY�UHؘ��LuC��қvC�M׾c�{�|��^��sI�(
�#c�I�k�:�B��)�C:"�3~�zg�0�ʼ
e*0t!�{�毪�[�K!�U��˕S����"$����;gbC5��!W"3�5kwZ��΄�8kb��Z]�Un,���L��H�fHt-Q����¯��g�����o×
6��<�܋����0�pNp�R�`��<m﷘�De���
����`�~K	��x��hw^O�����*y�'6F,�=%h{J���\�.J���e,�^��\6�kA	�t�%�x7��b,"=����d9�g�Z�UپV���}]�֔L�D/�u����uIS�Мl9�8̴Ǧ+��;�������ד�l-�N��TD�mv��2e��٩(!��^R�v"Kql�ۂ��Z��=j�j�e�@���35��6�x#Kf�'Ul���sD��3�P��S�,:�tŅ�g_�^� j��]�y�5��-=/�Wp��Z���b��72�hk�5n��=7q��]���]Y���9>|nm��J7���(�<Z����.�-�:'�Yw������aW^9�uL� T�Cp����|�٭���BH�5�,��+�-@g��XE�n��V���T!���}7]z��{:��Uþku�Ʈ"n1^#tP�,�J��t��|�d�T���M�z�=}1+N�=�+!ʚ9�b4�ۢG�o��0h���w��H���r��e82�c�텩|�㢩r�us<�x�*����-ʈW�eP��P�m+%v�=�g���K�A�V�kc8:�.��� �e��D�\�b���,]l�c��u�)˴AV1���{x�㈫�x�j�N}����1^�ތ'��O���	�s��3w^m�x=��<|��r/o��EbT�T`�Y�N�r(p_T�@V;��t�B@t�^/�h_M�h�CΛ���8�VTW9�!Ӧa[3K�ٜڛD�Y�F���MR�]R�DAZ1�Y��n�Z�2>u��<*��nPA�gv[���:*ؽY��Dq�3�x�K��L��F��˂c�VrX� L��Z����㷗lWY���K�w�����[%�(lo^s����]kF>��Fe����N�bq��t�1���ײ�J]�Zh�+\���T��"U�>t�+��:t��� )�+&KG).B�{�J�\���Z2�Ѝ7<a�QQ1,>��%5��2��1�v8N��X�.P	K��B���ޟZZ0?�*)ۜ`���s�k�{��G���@�
%�Ey�9&(5 ���Ф�K0z�e�sR�OVF=�{��爷_i��x�YCդm�7Ox�1d�3^}Pb@k.��'J;�g��gRs�LW�k����dnL��pň9}���X6�lX�}�D[.�V~�Q���y;�ѳ[�D��#c�鯆�b���0)��x��[Њ�E�q�K���B���t�-Z�=t���痨;����x��E^���9��}���Wk�o*{ユ)�g:�j���^e#l�� �����V�<J�T$k�Usj�\�ص(q�7�����q�x�d����0ψ��Ș�-	�n�a��T#re�I:���Έ���5�R͛	�.��\t��k�1P�G���hq�CJ�V��+�p
���J�ҝ�L�Ua`h�X���I�f�I=��]mؼ�N��iP��ɀ{(�#��
WR�(s+w��(`�\�u5���a��W@R���Ō�_�V�5,��Ղ��������A��%r��=���ٽڷG$��� ꄗ�꡷T�8�Qn(c�z�Q"y>��>X������G�HyQe��S���Ap�I5�.�tǤB���m[��!��xH�[�Qs��b�dƾ�j��T�ݲ�!�]Fzx�p�4yh��L::�V#���`����Ƙ��z�c��9�Q��s�����0/�!�JdK5�K��%�0�h2+L��F��I�~��<���,��nz��!�\_��t�� ץH29����tG��o`C~�d��Yn��{���KT-��6��%h�5B1��eaR�a�6 �䁾��}�Fb�'M��w���<{7���ٍ��Vi�)DH\Y1:���a�ќ3C#!eAei���v�SM��|X��T"`��*���ؒ�xt��F�b$ד���3�ch��J�m�c]�	����j8�:24��͜�vP�^�n�̉b(di�S��}ʶ��='�0�N�{�_��?b�fg�ٱlϷB!{i�8_)��ڜ=�f�3e�/g$�-�3s7Iy�Ǜ�J��q�y�	���X�Vl�A\�x�v)�;��vf+���Y�X�j)���}Z�ێ��d�DǴ1e��rvޅC;����0�1r������&ƻк�m\V��ٺd�3VKwܯ�8��w9��Mn2�Z��;����=���N�M��F>�B�*���Kkhw��+ˋ9�ڗ�=uuk/8���.+��C�S<�U���¥w����k���Q�;���"�y��ۥח`�{���{��+zYv�vV����W�=�;� l�ΏB9��e�9�Ř"�< FV��^l���E�=,�F\N�գ,M�WjH�R�b1��������c=3�P��8��#u�B�[���!ӞP˕�h�w����0������Pq�T��@ϡ��2�4"�R6h�US���q�+�1���b��as楖��A��U�Ί�5�	�Ƴ�K(z�-L<�'���W�!2�_t*�,J�.���}���Z�nDX��|�U=B����(�����n�c7.��.[�[q8X��e�;��X\tӍP�(�N0��T�T3$*��:`t�	Rj�+)-O��n..]Gv]2*��gO�1�Ȩ�n�uX��a�������^0P]@3�u�t�����w��4s�΍����B�7m���y�Q��r��=}�>�ݷc:V롊f��gD5^������VN�����˝��B5T���ESp(�X����*��)��2�8������!
�:�7c�M�6=^5D��F���huuʔ^9��^p	��(+<�578���;�s=h�����R���t��Ô*x����r�<&a�^PH�5��b.o��r(pczV�����Sf`���^�����ɜlO���c�#�~�[�4�e޵Z�Z�(�y�V̑tӽ��ɔ�����XQ9��Lz=��^�S����Md��A��h�;p��)��u;���0����SR��`��W�5;�7���ۧ�����4֦lp�
��EZ�f�
��JC:^���kto��X�v�n7��nk�ǹD���9��T��P�W>�."��1GEu�zy֖x����U�A3;���H���/W�xwQvr�jb���Դ8��2��,Ҁ�"���t���۳r�%���ܫ,l�MHd�.�-�E	D��ߧ�<�����_������汋ets�*�>�]���:g��W
�T���v�П,Z�|<X����#(׭%V��OTt^�ȍ�H��8x���1,ھ;�;��Ga�W��戓�����J��TO8w�<^o�E:�����>��ַܝ��sU ^\�pU��#��<;}�U���*���E�1�PިCiӣ�:$����\-�瞳t��'`���V;N#Ҧ����W*��(R'X�)P��Go�=�{�u �����t�E�*���3�mՙ,��(p�3��3)��Fe�^�w�� +��@�(5�	�φ��'�휟�n�{�­pz��3��vG;/܅���c�8?��t�(׆2��X�3��� ��������=~Ļ\���t��)[,R�`�,�@�u�0D(x֮^Q��i}��o��[�z$���ن�:�*�'�K��,�E����\��v���;��|X�f1�M�mWLG�f
c��=!��D�H��䘠�d5��Pg����f��4z���;[����ݛ�����@��
.���2X��\��2Bqq�40��ᆲ����	T�:Y����v*c*�"�e^6m�T��wo�]qf͆6���E��m�n�ezŐa�v�!}����s���~�O��]Aٮ���t���>�@.��H��8l�n^�s۾W��d�-����cE^c[#�R�Y��u �o�<�]swKq�I���g.�Y���O,�:�[�N��ۡ�����wrYJ��N�ܷ�U����乽���P��۫۝K7���]I�o���v��WI����,�J���BZf��=*qH��}6�k��b�[��kh%ׯZY+������UX�e<���PS�>Z������|�N:�>��ȧAmt��jײI��yN��L.2{�֎T�s׶9�R�rm��h�ċXZ�
�9z����}�oR5�����^>��6�P��':���ù�� �!�~��89�S�.(�a��[F�R�������a;��!\�8m(�����T�uu�wٝ�f����RV٣ΨU��6��K fҋ��{�*v����}�Y7]$HIL�"��"�+a��i��t݇�ļ+p��cw�u�X�jY��`�)�,`B����x�-�^��g�u涞�V\���7aņ��kA:��0��Bgυb���V/3�������"}�,$(w)2��:f��m���b�`�G�o_IE��e�!"�$�.e�m�X�TP�}h�����}�5����sC�|n-w)��}x9Y��o��,��q�]����&oa�7V=�X
���R��+t.�����Vi��"�e�2ln�"���!�{ɖw7+W'y�T��X"ߎUД`J���[҆�p51��QXqt1!,\R���T��k�ݲ�^>�U�]�6�r�	lh��v����8s��\3��nm�W��eqdc�m���>�huEL�:�w���Ţ��e��UA㼰��̀ޜ���W727�w6�p.�_d�\�٩��m���Lļx�����ط�!�]Q�o�mC�ٛ������@g��w3��\�t���iu��!��[�<4����S�iu�e��QA�N�\�v��Ⱦv�N�9Qw�_�5{*lZ��:�T�C�s4�P_7V�}{�7��i�|R��]��kD§����j�yE�����%�Ƹcf�S
��p��1�^G��x���V������@$�&4�/��(/��%�ͬ��D]�&Xf����Ē����u�k���  Ѐ$C��H�2�k�D�G�(ZCHE�4��.�kmTF�fVr����H *� b4�)�l��쯮���0��<�I����R(oXiYq�a���$0��B�g�a�%b�=�-�\2DA~)��t�M{8�� @`<PAP_� n*
����������Ez&������>)�bO�M1�h�3�g�S�$��
�����h��Dvy��-šw����dl�,��{�� Y�kP��І�7 <��b1�U�G���s ��PX�Ѣ�RvT��"����늅2b�
ea���T�4����qd՘|�fx���[�x�_�mm��WK�>�j���qJ���1+��j��A^�C�:�4�<��ri�e�s.�b��=���S��{�_օ������f���%�w)��̿�dڶ��u��T҇B�|��k���
��{Hc�]�����&8�q�T�E�ć�GR�*f(������b��N�&%v�k�(\L�fX|˟ڊ���g��Q�?p�0%�OI��"(�,�$l`@���p��ۑM�+R�?]����2}��A���}�Պ�@��Arh����!w&�@T+��́#[߬��H���6�@�����Ԡ'>[�Me����q^��=��'�=��bS�I�W��
��:;m��Pb<�d�y���G� *+�`�s�>���e�3�<��&�������hK�0!��I=�$�ZG��C��<���D>���g��cC-����U�P^]���� �~�j�5.��x�A�'V�4< �C�L;o;�,C�,/va��T�`^������kp�۩��ؐ
�vvHݵ��+�[
t�Δ�t�A`A�$^��������"�(H>|p� 