BZh91AY&SY��"��<_�@q���b� ?���bR��   �( uT(JB�J�@����I!�((�B�EP(�
��H��Q*�IQPUEBUJJ@�I#@B���
�%"
�@*H��J(
")!*DUT"�TP���!UH�J��*�@C� �{�U �x��QTC"�$�\�ED@ ��p�*�
vTDJ*�w�=BE(R.{B�D.wrT��)��"V��$$R��    MOU*�M�����j�)�m6�D�kT٩4����[*��S����j���ʪ��F�m��eҪ��]��T�*QKZ�JR)EL   ��Ii�J��;�J�)�]��e)s�r���t�ԩvj$��3��\�J-�7!J�U�6���WM-�%�U�yJ���ڼ���^ګօW�x"
��!
I
�   	���T*�`��<JR��<���QU��y�T�QOx^��E֔��K�<A�����z�L�<z��W���^{�OY�UR����ԥJ��D)P�H��R�J�   g�R��{{�=�;�D�!]�y�" %�U�T��jB��;��){�o^:m0�K�S�x*T��{Ԁ��w���
%��=��)<$�
�RED�!�  l��z׳*�����]�����z�(J���T��+zK�zE^ƩS�{�W��PoG��G��OB�����*���=�^�T���u�JPP�QD�!�%R��   ٞ<���y�{�J�]��Ԥ�ҕ^�{�*����5O[jEK<7EDu�+�����EM�{�@�
������e=��*����D�R
�H���   ge�UT��{��!u=V��SCg:�T�L�ڠ�ΦQ�P�dXt��+i�9��Q@p�t9@"�H�J�H�   p��z1� n�7@�mc�Y�
r��+sMӱ&P���NDtr��9et#�R�	J�	J�Hx  7 �@.p��\:hh7U���2��� �t���@�����Ӡݽ��z�pUB�)R
�	<   ��l�v��c�� �&  3K+�
;��=t�P�q՝�܌���y(O�P   ��R�Q�  �b` "�ф��*10�	�0�)I�z�h	��I����4di�L��1���R��F� �& T��3UR�      I��ʅ*�0 44��������?���Pj�_�?�k��J������*�O?7=Û����9���כ���J�j%*ʪB�I�uܘH�]�C}Xչ�~o����Q�d�U��ffx7I��˪˞��2��^R���WV�͕�+ɇ��W��s���N�:2td�ѓ�Ό�: t@����'FN� t@�сѐ���à�ѓ�N�:2tIѓ���haѓ�N�6$蓣'D��`tI��'D�>:0:2tI�ѐ���ѓ�N�t@����ѓ��'D�:$����t@�c:2t`tdЁѓ�FFN�:XN�	: t@蓢GbD�4$���'D�ѓ�'D�: td����'D�42td�������ã'FD�:2td��蓣'D�|0�K&��|'FB��FD�: td�����" taѓ�'FN��td�����td�������D�'D�FFC��'FO��2t@�ѐ��сс�F�����F��4=:0:2t`ld:$�d�(��H	� :! l`@�C�@�D$�!�D��� F@�HH:�V�Q�*���(�0�с!�$�с�$�� C�BhBI� C�I	�I� ��	�	�BQ$��D��: 萁�� ��BJ!:2@:2: 萁� �F@��:0 td�`Ό���B: @��� �H$� 4ĶeTٕ�Hٕ�tI 萁с�BDN�$� `� ����	�!�@�H@:$ ta �! tatI$: HtI td td�t@�� C�# 'FD$� :0�:$tH�C�$��I:$�tʆ̪6eU�*0F̤:2@:! 萅I�$!ѐ!ѓC	�!!� � I:2: ��`�	ѐ�!'F�  pI ��� C�C�$B@��!'D�ى[ؕ�lʖ�Jى� D�N��N� tI����$� ��!:1-�JٕV��$�aM��ΈtIѓbN��t@蓢N�:$�N�(��'D��: t@��ѓ���'FN�td��ѓ�'FN�:2t@��ѓ�D�:$��ؓ�N�td��'FN�pz0:2`�ѓ��N�:0�N�C���FN��tI����:!�蓣�tI�'D�чFчF�â'FN�:2td蓂N�:2taѓ���Q'D�:$������:2td��ѓ��N��8!:$: taa�a9���3_�w��4�����1͙w��'N<Y1��@�Y�1�z[�[F�K�$?Q�Y�v�C��X������d���<��qSԂK{����+h�їE�s.a�lP�c����%Uf:D�e̼82�ʖ�(i�w��V�]�8��xB�o�olMr�ԗV솝m ]�����G7nM���ū,���nYz15Vڼ�i[�Md}-��[�&aئ����m��ʧC�j#��4�
�j��J�2�f���	"��Q��f�l!� ��j��Q�i+2�G:*`�,c$mm�n�%18`�3�V���夵���a��vö�_CW��E�h��7� �P��+�f��R�ٓӍ�ڌ�D���)c��+�v����ڼ����1۠p6+vե�9���j����]-T�O̈́
V1б(�T�a�82���3.򓫍�&ڦ�*�姀[�;��YA��\�%��hE�b�#��0YЩ���3Z�B�2E��v-{�Okp���ճIة�]�&m7G`'/$�WoR��"w�=�U���l��Y��������,a&gD�fCM�]İݿ������(G[�S�m-x/(3��_
a��U�$�NVImcˉ�W��1Q��/��u��&�eXm��XIR���k3%�����gsQ�]B��4 ٥���b��)fnO�q�
%[%�U�]Z +>��7mE�R��
�>{�rR�2;.����m�܅�][�7S5Uɭ�i��#��o�mnc����RV��V��#oE�ݓ��2G$4b�n�(�t�Ի��)VY�6�el�i�z�
H�SS�G�hXNR�Yjα*�r����jJ��V�a����3u{���F�Y�Ō��^9�k5T@Ve i:St ,X���:r�ҎV��:Uݧhmn�T-�.+4��X:q� ֢���wIx2F��%��t�͕lĂ"�=5��Qcvv�����%�+��W���,�)�|6�<S �����x�9�, �P�a�h:�D�t;:"{R�6��I�GA@;�ʇl��)Z�h86�.�GH�l1wHn͛V�9w!P����9�b!li;��)L&�p�G�ji6�!�����9�r׮�z�5a2+��30PXٸ�[R��Q�t���j������m�#h�f���k�d[�a��Re����n�c��/��k�n�Gi�A�Ǌ��+v�3N�����W7;��UA�_ƅ�5��i�ݘ�Lk��6�K���0�i� ��-u�Q�z���5&���4����:�Z�ك� :�t�2M`�z�Ţ
�)l�d��7cL���H=�=JA��@U�J��V�	�VU2lC4��F��MM�g)Ш��:�	��Q��"O��$:U�+Y'6_�1V��!6�'�	!0�ڊ�*�n����$�Yܖ�4��` 0����b���� 
���,��Z�g�˻�W)�AR �I�S6����-^ƶ�۠Q4D��i��[�eӵ���H���[X���be$n�7n��K�a8�.�<��++�P��A����˧K�bl݄C�-ѽeP�M�H��b���r����R�B:O���vX������ڂ7JZ�wh2��0`�H����Y�VU�JS�W+@�p0��Q�w�{�짲�Jn�soK7Z����zwhT*MZq�Niyr�ʴ���Ҽ�l�e��w6$�}�<��v�w���%�+0�Dȍ�������UۚY��{n�)0��<_rJJ�C��J��9�ڷ1蓵��Cg&�P��O0=�����Q�0�����e<v�I�T9��V����R��uej���ud��`�W�-���6y�%h#렅AB)w���n;nU���+.b��/�KiHS�VX���ظ��Qm�����"��SU݄�XB)d�l��\V	�W����`�:mK�e��2���i�ل6��L�-ԖҴ�v"��M�FM1�3��%n�n��̓���� \�b"e��/>���l³��IF��m�I�����.�bQ��Ne](���KYm�zէ�Zr���c֒���Z��ҤqR!���Xr3�!�4���	`^krIF���Q]�5�'�����[��դ�Dּ���V-�@)��{4]hљ����gnk��+�B��Lm"	�6i�U��S��"��[H��D4]�e�3kp� ��B�P��!G�^�%�Od�{u�!��Cw9h߶��h )<a:�=yX�v2�� �A�pn�Q��Ӥ��k6�*Gtʄ�2m�V�f)^����7F�^Sy#�țF�$6������r�#��(ʭ�Wz"�2�EG*ٺ߬���H��)�h!KU��2Q��7{��!����Oe�ЊĪ[{p�VK�q�f�6����L��1��sJ�.蓚��v��-� dJ2\u�j�6V�kh���AS&������T�7n�K�j�r�ͽO�"���l^�o\5a;�����ɉF��B����4�Sf�RC�JSt3{B@,��yQ���f�}I�9��t1tmM����e�QZ^7�N���'�v5��̵��C\�D��!������= ��TΖ ��M	W���Ȁ:E��+N��7j-��kA{.�n-�6�K��[�nYD� ��jaMKT�`K���v��(�HrS�v�52�#�ۑS�0-ː��M٬�B�J�f�P2-�>!��@�q�Vb�`�.����;O.�m$�n��(�m"�F��D�M=��hEl���2�m�8n*i&�"��v�4-љ1XD-YWF�Z V��� �uw�EEjo,Hn���Y�7@KY4�4�Z֧����G�Q��b�@&��n�KC/���RK[���\MiM���&J�Y��K��1Lmӹ�3�kM͚�)1�U��c�{*L���a�?X�,�e�U㡱	&�%�Z 8�G�u�b�
�$��v��tg�{�����r�֮����YODu6����pEY��y�,������ ,��Ti��ʚh����[i�ٚ+t�g[ζ2��-舤�q����@��X��b�{)+P�ZsU�i��%f��� 0��P�L��%�7@Э��nP���^�K����k%�4ˠ����f�H��51�ks(��Hې�Ż��!i�Rm�˻��д`Yz	ŉ)�`&䷸��f��Z�!#u�*9��L��Z�4��yV�B�1eb֬V���P$Q͛Q��f�p��A�DÖ�f�&ơI�k=+n���I&
�aot�u�����6�B�e�	�$��2$ؔq9#8��`�:�L�dܤ�"��㲮�^�2�P��ܻ��قd��LN�f���$K,�%Fi�����V^���(�U�9ob�oHUc!;B�'5D��e]hU${h^��uk EK�yX����CL׍�1��wx�����3hG�E3IZ��VQ��ܲ�GP�� �-�j������7V��KFжCSv�8�Xǩ���b׈1��1�1e�PW%i�t#�̆��� ���އz� ���^R
ܺ�D2ջA۠���yof%����ԛ��ʔ56,@��L<m����3)����k9b� �VHe�:���.+�����zB�%ǵ�):Woij0s0�/i�m7�Ƿ�����.�l`�r�I��婁
f��,p��9BU�wZ$������Iޙ�C�L�4���EJĩ�u3-�r�d�ʊ��;H���w�e �YA��9�IQ=� Y�mQ̥X�l[
ׁ�2X��d���hV��rRaR5�,���X+	�B2�V�P��OkAF�r�e�wb���[Vh��VV�fYs�V��kEF�F�6�7�j����������w[�̈́�Z!��0���I]e'J�S�����S;��	��]��h����Ei4�^���!�`e@ol�Y"��
���r�O��Vn�����Z�|� ��/�"Ѣa�e^�ل�5(K6
ӳ��+.��Z؇*�͹��^Pvv�*�3#Xt0=!]��L��ǔ���#gf��U�6eo)I4X���!���ôen�������S.Rr�Ņ3PG]�,��*��kFC��-V���
Zܵ�"(\�-ȥG�Y��dU���Dx³A�\��Li3��0aOp��{�F+*�	�(�0����Z��Fr�˰%:�C��4h޶��w��f4�ZРb1y�ƅ����%y�D��Z*�ѕ1-��k9�j�l
2���D[.b�2>�4�pmlo]�Fr�iJ@r��%�J��ɱJ����j<�%$��8F˦]�sYݢjEB�S��iֵa%ә�,�j���1t�[u
Lb�B�5�;�ٴd ,`�#X�)eW�V���n�EX�ϣ;iA`1a���w��m��� f���5Tj[Rf<t��܈n7b���Ӽzi�D� ݖ�NJ�
�(7�t� ni:��fժ]b���E��F04�n�#��70(�X�bh�0��;WN���q��m�B�s)��3$0wZ�l4��H89��Jvq���EϦ]�^�y�ջ�m@�JJ	t��U�*Ĭj�Gj;o2�]�"X�X~���ۧf�-��SQ\�մ��V�ؽ�b�����{�%�l�M[�*.n#��]&m�tpE*�*��d�_v䘓R���!��b2�VVj�C��[P�a���K�{-<��Etu�uv����q�x�;��u`�C!W;����n�m����O��}��i�˺k7��C�<ea{�7:�A��)�ܛ�U�@�l�����So���3�QI�q6�҆�`�b,��7	�p��Ǚ��k��ݒ���#Y5f�h]�j�2^��,�0VZћiE��V �?H]�XP@��鿈y/m�n�X���!��d��^���2SSj7��Ԭ�w6M��fD5����x��`[`��$<�0^����K��i�0���+�W	�����˘ȩ��0�-`Ej����l��5���lĬ��#�2�Ǐ6�Z �jN��4KV��n�B�*�v��[V�A��m_�{hQ�����x���0��Њb���%��%f=�Т(�V��S6�[��ѥ=`Ê��WBܔ���z���\m
����$1�-�u�<TۋcR��F"u乳���6S�W��&@�كA|�������iV#OR&*?6�@�l!�nn����cm#( ���.��)�nQ�k��f��a�*�,��'��Yl�l�z�#C[���ӻz�,���B�B� �7�b���d���n[�����1J�]�׹
%�H��E���i�������n R�3Y��Ҥ,P36n�t��U��K�q�{��ݫҳ(�"b|����%^�x��1JnAT�쳶*S��j +*�^ca�ZD]���yx[ߍ�X����-;V�!mh���.l2
ieG[o#��dY��n����D�ysE��*`s�yP�$���.�1�]B���Y�U��^�U�I�;m)ٳ��OA��GA��U�6]�!N���@ںm�[�{�*��IRBᔎ?�SEAgj�E�֒��0�G�
YW��6�5e*SB��k�e��cb�(;�2�nh�����R�p6%<�����9E�h��ٛ-��pe���C�P�
{�)u����h2�v��U, �I�nX��PYl#��wo���N,��B��5�dA�	�yP6�J�j˧H�PiϠ�a[V[X�I��G��VMJ�7tB��#q�n9���V%DjEL��ܻ�zQeG�&�P-�6�^�����*Yhǹ�r_�ڂ����T��j�:�L�b�m��$^���\w��5����?,ބ�u�j�ǫvt���3TqU��=�p%�n�-śNűxQ1�j�.U��O�ɘE5bnT�����GZ�wI��嬻R؍l$�Ϭd����e��{GF�kR*	���^T��ݫ�(m�,H��2h�8qZP7р��a`��#Vm��kZ�:�Y��/%j��ˆ̒�#V�M��ݴ��S Eaf²�s`�����U��s�t�:X,+^�X7jl ua2>փ�&؎��O'�i�\2l�@���׮��k)ՍWbȫR�[��%\_@�b8�[���?���E��-9v �n�����xne԰v[��& �/	K\��3p�q���#9"OufAq�!e����溎\S�x3/۽T��Cu!��+^��寛�d���S5�4cWxU�1��ѱ�hĭ�KhB��[�)B�{�
�c��U�"��haq֘I�:Ĭ��H�N�:u�o�LgB5,�Gr ��<0| N�[�O������E�E�[��@�Mсh��w��̼O���+X�\es��c� `¼�*J�໣� �q�,��Pz�@��`���#� ƥ�2�`�`�v	U`��l�CZ�c�>���&4X���b���������ý��
F�`��2�6G��4L}�Z#E�4A�0 E*@�-A��}W����x�]�j�cs�4�XW�t��uޣ�Xu���_��jf<eUk�nݫUZ�W��s7ۧ|z�zW������W��W�·�ֹY@B 0!��h����W� �� .�йs@���:
zu��A 
���������d+1QK`eA4 �Gvܪ��g);��Q7P`�N7zv�_�x�t���v��f�L&�Z���+A��Q4�XL� @D�@�- 2���������]6�:��^��e����������ׅ��~}K��/v&�1������ٍ���}+�GK�n47���T�l�e��=�|�gls c�{ӆ���d�YO&�"��A����uͱ�<��wDWI�Ӫ�H�vz�z��N��#�x�8�)igK���H�+xw*�:�{�;�S�Uٝȣ��Z�oU��ûեu>JKuq儉P�v���A���n����M+� a��1��(3�l�>�u�O��o��-��%dMz�3K�J��r�j�{�,��N��q&�(�)����ڽ���#Z�vӾ�/*s�J�=C\���|�9��>�2ݽq� $I���&�ີ�A��x�	�k���7������dr� l6�ܢ�ե�a�;�u��2�+��Կ�' ���q�����Yd9Jv
��S��k�I����g�cwOC�r��R���5w�<�O) ��e��B�����<N���2��J��͒,N�1�<�-����L��6��!�N�{G=��{P];T5��pٜof���f�Ӻ�~((��Rk,�S�gD�Y��y��;�e8��C��E�����k���,����{s�k��WG$HL�;YotQ}4u�3T� kܫy;W4� �UI��z�K��yb���N��$���hlٯ��1]�
q�u5���`�͑�������+M�婽ȧt�B�#3O-��x��2�u�a}��Z�r;YJƵ~u=��=�m
�W�斃�Ѯ�Z�*�)��׸W+�Y����u�g:�u�jb�5�(,��+����|.��2B�y���r�C������h���VzH�3N�-p���}�{�N�JS/v��쫛�d2x,�-B���*��զ��>�7_X��,��[Y0&���͖���zm�v���.��q�԰x������N�]�K�72��6�S���)oV��P�Ī[-l�2b�R�Դ�S����u�Gc��+]�>롌��Uy���������z���`Kr�j��K���Ś�������(����}d��Ky��'�j�����`)��|��f`�i���݉��a5����v�^��)��`�X�ܹy�8��u�ea�ֻ��p��`��`��X�wz7]s��p�c�� hsh��-w,n�Ɲt�p�&�V%��fVd�R�l[�QǕ����a���Gpe�|ʿ�l��e���l��\9���A&-|�<�1,\K�y�x*U}q�4���)Ŭ#����u �K����<��+�w$f�	ʗ���.'�
Ѷ��4�}��nix�(�Ƃ��4Md0"��h���[�����5	(��^,��H�xy���V��N���m�x�Mϖ��QU�b�T�!M��g��פq�n��4�ۡ�G9O�33��@�K {���f�{�i��ґS(`b��a�I%uyC�C�u���h�C!�B,}̂�][�*�3n�.0�Ye��T���)��;&��
��ӻjp��ץ���Ɛ{¶G��Zlj��Y�*Z�I�9��!��+�K ��*�,L��{KZ�
�#+V3V���_e��(*�-�f�>Y.��].�nA�j�f�U�h�9D�7�l�Q�t��/���ks9����//T�Q}���O���Ǌ��';��֛�\�5�-�=�j�s����E�������\�r���W v�c�X��i���t��g$��(�;�@��r��̮��^�'����ʻ!a�.���5c3yW,�,O��1[��`��u�gf'}(�%X����uxs���B�2�f$3�尝�sbJ�ݳ��.Ǘ���o5]c*�Q,��b
�加�sxۮ�6$�mm�*fT��3����/ق�4�����ҍ�A�{=h8kv��1i�Z��0���G���������X�J�2���i�w�f�s����s)�xW����b��C����.����d�ÍeζZ�}�_S�p�].�|�<���;I�Y:D��:�\�����+�/�B������.}Bc�ՙ}�gws�6��p{[Mn��qѥ�[!]յK��*Oy������ff�+�crE=��C�k60u}�j���L^Y�UR�� �
}���1�?:����E�,rP<6v=.Wu�b�od}�Ѻ�ьu��2���gZ����}�>&�|�=<�_J�3�'��d{-f����\�Gn���mm����J������l%ʍҨ�1�	��鉹����][Z^�z�i@�����+�MSE�|-l�Ѫ�Ƹ�8�ɶ{��t�Lg�>�j��>ď�5v�C�����R��G�,V�<um����Q���;���R5����lZa��Q����8fY����q��I�q�(��w����/`b��j�t��u F�橨-R�jT�,�<��%b��X�t���j!����=ܢ��)�Ьhˬs���Ն���S��� �ݥ3����9�65F �6�a�u�1>��c�tv�pnIH!\�-��V�=��4�Z1����C�mpW�嵵&�}��E�'�m�,�3�2�%���L�]�Ú(�b���h�)Jj���W�V$9�ձ��f����Uu��M�3�\�ٓr\N����c���WS0V��I_1)�ޖNK�V����Zݤ�����s�ѥ�C[P�j�X�R��a��X��1M0痥��eD����#�Ö�eL}Ó��H�8�#C���I��и��/����έ� �C���o"/��Ta�]\�Fa�;��Q�5W�6c}Y��y��Y��zWU���'L��y��[Y�|�2L�#�f�
�=/�.a)}��6���Ǳ,�o��8�"b�qV:�Y��L���9$!��s�P K�Rg�{&䩘2���^h��a2G�&tU�Ґ�ܫ���Ή,Ȏu�},����W�`h�v�S 8k��|C9ۄ��4(h6;0����[HS�ܠ5�ف��Zm���J��h%��F�㝗j�0���R���AN���7e�#K��!� ���;�Ve��.��k�j�w^�gn���5�[�D��z��.�q^я�L5��mʵ%v՗��֯��K6����cOt޹.�� Cq�2b�J���}ap��;}���1C����WV(f���|6��uMw�t�&Fn�.�p1nE��*�g �Y��_a��y�DU�7Fm7��b��m<qIN�g�y��j5�kM��VM�j!-sM�*�i���.�>�\k]cS�2X�l��%�e"���^oS�1mק9<�f�iꙓ�/�p�#�Q��xQٜ��@�vE�E7��^̤'H��v��rp!6�u��v.X�C���6N���G:u���P{��!�a0��k����uu�M7 ��Ͳ$׏-���W��C��sc��Pf�ɪ��x�b�9�ħ���!�E���|z��;;�`�:e�,.��3�F�9�)�]�`���h�l�D���ŇXk9wa�o�[��M2SŶ������R�e��Q�GN��F�Pw��o:ucnK5���[(gi4ѹoc0�E[`M�;t;.�F�2�Y�T9�����4��"�Z$�:��iKtF�0�v��;�+�P
e�:!���ߵN̎ʘ[���D]�@s��+n]c�s+��&�㹌�������Q�Q͇�B�VZ4� %L�}� �!��aW<-QwQ�۳�43i�'�Wݵr�z' �%��uuN�7�+M̭hc�/���j����N��vl���C�XǻmBӇw���v�GN+�ꖽ��9)���%G��;��pɯy(�Yj�W�IL"��Zv�7N�	hۉ�'ot�F��&�2�NLn�-���&��k�]ܭ@x-��1�k+��z)o,�Z9�����9�W,��]	K�y��<��n�Uo4i�
x����5����.���3���F XĆT�̍�t����pu��%z�g�59\\�)�ֶ�p��v̹���ܽ��Su�lB��eW[A�Ȝ��5m]ra( +��הO����Ds:�tj���À�ݮ�|.�yk���c}C��כQ�h�[� �Iϭ��Q;�)RՓJ/`�usT��t�7uv�rb�|&�� ��@����!��J��+�ky�]n�oej'9�Q@^K�;�bh�.��zJA��v�2Hj�ɷO�"ԝn��x���ڹ��Svs�|����jqZ9^�~�|5���6d[��Ԟ�Gr]E�����u/:�����ȍ�MZ��CoHwO*���k*�ժ���y�	��Hgv���������-d5Sj���Ǳ��3�b�����gF��P7�ڏKS�ʙ/:S�a���=)��.E{�t��!O���s.���}[5��I�4X�\b=�Ӯe�LkT�mҼWܢE�.��vps13'>6�l�u���x,��&ɣN܁T1$�q5��\�|��g�1h���lZB<yLJ}�mc���:�,��o�qo/����	������\n������*�\�C����p,���ޙ���#��#s�M���sC��k:j���50J�)���:�B���6�1>O���3���Ǭ��R�UEJf����L[)�[ѡ���V>Շ���g.��1m̱���l��ȡ���U�z�եD9���-���2�ge�bah�[����=�-=������dS��۽�hrS�?U�8f5%]��PL�ށH����}�C��%��r�� 6.���\N3M�QC+���M�:�	����m���1��Ar޽t�f^��4�}c�1��JY���k��x�廡��}x��u*pM���w�����^Yie�l�T�#Qm)hM�ok:뜩8�;rS]��:QR�8tR˳ʯ4V��\Jԫv�gC�'{�m�|���\�qTO{(Lu���+�&H݄�2�q�O]N����iI�M[�Teqc�L�\�n�]J/������6�=ə�x�M㗤%]�ե*�Df�y��{dmfVT�ICv���u[��^��O�b��-.\p�^#���ı	�JE�.�6z\I
7��͝xW4�tnq��<�3�7}�J�����{�mu�ӕ+A�9�D�6\���T��u��k��Z�\Uuv��51�w\AF����/�ɬ����M�P�x��wf�t���%\Հ��*ļ�ٮ}ʯu[�A�:^>՝)�˄�E� )7}ܸ�^y���Gz�����S�X�m ����'���C�ض8��gi!=��f]w=3v憶6������Ix�ulq�R�����B�k�6�Pޛ;]j`�4�OI[.p6du����ң۽�V
�Ǽ[�
~?sQ�ef"���^R�qZ��{�VڝL�˽ ӂ������s��ms[����Mn��P���-g7���ռ���Ě���j4>(+YN�CZu�<�`�q��¬��v]vV�Z)aǻLy�'�kA�t�"�q���	X�3V�;�l��-7DcI��/mPWW�s)|�����MҪI��r�*<#v�Җ
��e�5�ΎM�n��I��}J����:��UK����D0�<�!}�N}[c���Cir�o���#;Bb��T�bY�1]��u#;&�Ҥ*���sz���h���rU��N�-r�BT�Y�ԏu�)<�Z��|��Py�.�=�n�mS347�s�"
��w�u�:����JotU	7/z��l��H��\@�GA}|:uՉH��7B��/1���O��sP�]�(�÷���,g\�\�F����t/7����2�/����%6�1�����0G*�i6����y�J�ǖl��}��q\�Ҏr��μ�So𗧩��M^:t����tdw�v�Z͑"�U*�fJ+x%�:�q��lx���|v��p� \*_!�73n�1��%�F��z���8hg:�a&�
�Wh�p)z�#/���k���i��WopU��������m[�:�1��7��kN)X��ël��w	��ܮ�1�ݏ/;���u�e6������&F*�X�K�WtYu�t$'q�/��+���91ջ�Ӻ̈va:�kxe���ʂ�-Uku]�u���E�V��i�����+G_j�W��̈ଅ̍�+��B�1ͪɗ<u�m:J�S�d�\�W�v���q��	Wռ�7���u�q7ݶko"���R���#�ɽ��v����V���QJ�������l*��QwY����ְ��2���1:�׊����}����k�ǔ�왰7fu֛�� �]��l��Ytz�+w#b��*�ѭ�3vra#V�+�d\�F��m=��$�A��%�z~� �s��YOo6I�K��js�s��"f�gP=�)!�:�������r>��|�O�Ƿ9wL��v:�����$��:�4���6�N��M=��gNuڇI��9��s�]v/�=^�V��p���G��V��ט�Xhs��E��N������v]�+҇N���g}���o9z?�I�I*Đb�1��٭�µd�h�&@PA�"�(���}N�f�0Y� X(�q�J��4�Z�����k�3��[�ի�4ff:��10�mJ-՜kQ�8Oű��lqU�@Q&1L������EB`�Md#���S	��R�[,TwJ��A�&�V%�	�7�*��F�+X�<.�T���IL�B�U*I�p�I�IEQv+�,��oM>��P��$�`4٠�����f�H=h �t��X�Gb�f�	��1��ˋ6�*F�a'E�4HZ�J�&�
*��Y.��ҏ�K��2�i�����7I"�,K��|��rM�R2)�σiR�NU�B�[{f����S��N�P�j�$�P�*��
�V
d��;@:N�5(
$�)��i�i��r�#@�~.Z7�Ƥu����%B��J���uʙ�l���z�6�9)�]�aۏm��ꕪ�t���d�� I������ǧ�-��{/"Q埧��u:�G�B���(*�ğϡ��?,dM�
�7��Q9�]�jޱ���K��gsUA,�����pV�B@�S�S Rg^w-xed��,+��K�����\��u,״��(uCm[�\
����MQ��[��F�w,NF�겺��N]�T����r�QUѣ�+��o��@3U!V��6��rHxV�q�q���y�)$öx�t+_�f�t&6�J��@�\Ҽ2��̾z�윢y]K�m݌	�Z�Z|���#�Y���ut{oMZ��UD�4�
K'+T�y�wI�(1��4�\�{*;m�E9	��(Ў�j}���A������]�BE{�Wm�YZ@}L38M�x��A�����0>m�R�T��V�y�F�:ޒ�[lAXq�Q
us��77er����*�}�uj����9�G��{�y�D�� w4s=�1�j���"�E,і���q'����gi
�C������=E�Z��Zү��]_^�+qdq�n"������LlG�`ᷝb��nM	'8���'�**��BWZ�-&gP{���l�<Uժީ�2��},\Ѫ��,:�{�G6tcS��n��C/�e=W�x!�RR_+�Zҙ0�J�:�u��m��z���mc'(��\�%�/n�g^�7.G�bu�K�h$�|ܨ&�><x����Ǐ<x���x�┧��<x��Ǐ(�<x��ǎ�<x<x��Ǐ<x�~=��N>~v(�+;�WP�0+�Gd�
��5����\���Eֶ�Q `�U8�YK�ܼ&L�����*�Т��w���y�w 
��J�J����9�����Ws��^��8�|4v �SA\(��'U�Ih�l5��':B/6������)�D.wH�w]�����o����]eϴ���?�CY;�eu��yY�M��Fk�Yel9.�(��q����n&��yAgm�c�T7'C��qJU1-�j��3;{3��R� ����	��ͥؓ�9g'u=��v>ǺK�}7�����x]Kk��Ug.���f�r��wRث���
�\��Sv1O:g@뫨�n�o �����a¯e>�$U{F:�&���%:]�F��H��j\M��y�۲�@,M����3����I�hT5ۻ{��g_:k�*B�����F��]�Rۼ�_�i]X+���UN%i8�s50u�]*�Q%�@��ިBL�q�3v�����_VƎK�X#h�i���n�A�eZ�*B�Y�6���MD�PxM���L��v�o��o'*���(q��S}���i^��Ζ���[�1;��Z�x�*�<���S��$&):�^���G�U��t�M,�j,ۭݔ%��� ��(��%�UH�ew]��7o���}!�'sœJS�wTu ���Q:�W�Mֳ;�P����ԝ� ��S�N,p���0p8p�Ç8p8p�)�Ǆ��Ǐ<x����Ǐ<xp��p�Ç(p�ö6�DN6��]�(ɢlcK�u�;w����X��J�do,��(�rU�)���לt��]�j��\9݀ɺT{p˳2hƷfws;�
�Em�UC���*^����P��xv�yB-bW9T���nD���/Q�*ig��mJඋOw:vOŹ���k��t���fÀQ�lqǯy�#�!҇6*�Cpb�5��t�ۺ3y�֌��v����U�6�eo�5�*��5�� ��t{˺wGy)����-���iZD3�ݚ璹[g����+ ��Q����k�ЙYr����vTk���<{��;�
vHYK��UG�삮on�5
�����͜��&)��%�SP �
h;�EԔ���#��჊P�7Fk'��6"iJ����|k�m�GW*Y�r�%Ǎj/l�����V�C�e�[�
���ި4��n��Y3:�{��{�h�nR�S���6��22H��-L+h�q�U�N	�_m���Ae7Y�o����;%e����ꕖM��7�eF� k���wW�N��.��ӆK���x�eK�.��V�<|�z_f�z��X���q.o���6�K7�K�3*�t�K��\�A��1l�N���6�� %`����ҧ[]WF��]e��<'�<x���O�)Jx���<x��Ǐ<'�<x���OB���������֜�g?���E���-[�X�,�ʁVN9V��z�4D ��Ε�M�6X��iL�EMwK;t%��2�ۭ��9Rͱ�eW0�l���c(��e�f��f�E/�����[�s*�5)1�L[��u����᥎J��ٖ;��o���Z��X��(E��9od�G���n:�&��Q�׷�d�ɬ;��:f�jz3�m[�����c�`R���&���!��#r�۳ΡEcC��l}_R{wE��b�#�G3�V�}øb=���5t�z0��jp>
!�6;&K�,�Hb���֊��eAj����C&o���23��"�W`#[�i�˦q�`̯��L.:���q�_p��dӟ==OX�2� FS�4�s�U;rZ��(���rP�	���u	�Z�Ъ`���b��.}4啙���U���б�]��E"�Gl	�N��Q�k4:�wذ�qŀƨR [�q�'I�r���f%�8�P�U�zQ��\����[] P��]��NR�nl&޲cɄt�r���S��������Xh��(��]���t�ʽ�V�1�vU؎Z��m��o&�kawLs�| �-�UU1���69��k��]��Z[���kv�X��p��l���;^�p\o{�)���%+[`4���f۫�^�ҁ�ޡF^���M����h�����/xS�ͫ8��%}"���8p�٣��<l���<x�x���Ǐ	����<x�Ǐ<x��Ǐ8p�Ç8p��8p�]�Q��]`��n�l)\��f���L�{]��ZRQ��%ݩ(��%U�e�fp7�*[�̪г��[��\�2��
=)��� tѥ���$pǌf��Xyq�Acz0j�n�]ʰB�R5�뢰aeֽ�u���.���h_v�@.��S��F�G[�G�U�)I��_F���t.�[\e�)��<�O�,�͋��GT�N��m�Xf[�g��v����vq�C�:�0��:�z�_W�:�۬�w�D7�I�8��PR�ǥ��EeXv��t�+0��6��.����e���>�vW���#U0;v�s�>ʒh�̘G'ې�}�\y9*��戲�2��GKJŵ ѐC��jul�kM7�U���[��i4s�9�Q��i*`͘�QW��u$Q�مږ��U��	La��cE�f^���i#��a��[GE[���Y��3���:j�I+:��1��s����6���ޮ0P9�wZ��\�$�4�0ƭ��3�i[9�2�ɢ=��#g.�<�T��3� ���j`�v&�3�*̺��6��s�ղ��7,Dj ��e;����X��'��opө����ŁU�W�����Ac�٫{dQc�����h5c���[`e0�$��`�1ۙ�-.�ŗ�m�75H�����Kh��v�����1����ڒ�%uuu:��++���G�<a�Ǐ<p��<x�0��8p�Å8p�#�8P�ÇWWT������k�>[�q���H��ժ��κ��CV>\x`�_)\۽��E�1L��dY�'�WF+��܄����}ub�	N|�_��Y6vR�
څL����\�Ü~���<���D�5�~�gP��wL�;�����k���-��bf�MؕJߠ�M��c{6�:�:���&�oEue-�e+���ͬs@��;��Ʀ��m:���5��[c���s�J�5	|�B��>���,�»]f�'X*���}�Q�vx���� �].�c�
�4m���ȑ|�����a�<�ʜ���ٺu]; �oz�Ep���ylNvV�uf�$�
�ִ-f�E{���d
O�qܤ�l�i�9��*�k�S�k��	���R5�nb�� �������=�H�.^����+�V�ݬ�6D�C]�W��p�c�t�˽��e):7���jܵ������K\����au͚�hS��t�O��@\�'8u=}F>�7.���,$�FYr���EΤ�.�:�ʝ���T˹�5rZ�����"���U���9][�^W�+\���+��KB�Q�{�I�L��������;>Y6먥��ZQY{2r[w�fռ�˽�ZS�	E�(���ёU�n������^���Z*�^��>X�ʙ���y�ġ!��6yh�$�ч��ݝ���T�M��4p��E�8@�Ç8p�Ǎ�<x��<h<x����<x�ѣF�(hѣD�4hѣE�4Y��s3�|Yv0F���%Xو�@7E��L��_J���|�3V|�6+O74֔�":�C��b�P�vbY2�+U������+z�b˩7z��D��5
%U�("�^��K-n�Wd�^aV�"7�}R��U*[��M�ϰU�Ӗ�LM�T�H�z�
4���W�I��V+�����o:�������[���Y��C0oʃ[5�e�d��U��S��Vԛ{5�}��:�Wk4��Ё\�Hf|���e���#���뺚)["����WWoq��r��t��=�V�vA������p5�ۧ�F�2;j1���r��8��*�Ϧi���Jc�g�t�m�3��_҉d`�x3ɓ���
R��or������Z8E�р̽��2H%�rP�L}1 t��qQ�e�6.��w�VaEob�m��j�rKh
����
���Bus����U�˥�oq�	|����3�6��F@G�~����B�t�s/���ʺ��Xq���]x0�:�d��*nL��rʋm|��#�QU}M�Ce��w����:�*����-��l=���fZ̕��WV#@�-�t�%}L�q9������Ap�?i�w�������>����:�d�evF �0]��Ip�0�2m	'\[S�(�k(����Rf���cTr;�ۼ�#��d�D�������A,�3�._wj���|t����N�<SǏ<x��Ǐ<x��0�<x��Ǐ><x��8p�Æp�Ç8p��l���-�$ݚ�HP	GGk�ﾮ-JM\y歏nF�w&;�me���(�쬩�^'lvŴ��_\�	�1R�{j�ܧ�x�W(,��������j�:�D�9�,�*T�s�}�)X6��o	-�KV��T3�u�W�Ԕ�'�*���,�Vϒ��T��u�����u�]�dљk]_p���n���͔l�X�FA�#�M�[�]L]�uҲ�u�ع��*�/\LK@�M���ʃ{��9��t�w�q+�u�.�0�	�Y�lVՑ�QVy��Q����;�û헢.���8����Gk#:c��ťN%��6�X��tb��D��/�F�+�U�x+B4;���#2���3�
����73�Bp�_w�5%�½�)s�V/���d��T��6��b�<�e$7�����қ($�N]%��s��hz�벾nZI��\������K�!AN��
R׎��$�����k�����N�m���~Ԥyܸ��G�3Ak�Н,.cu!RW_`n�����i���/�)��iaM���7�a�T\��UJI��;/Je�x�R�Ec�4�B9ea����g%�Vf�G�؜��(�`c��C�-H)Z��/@�-��n�њ�R��(��M��_V�S��u��o3�jA�P�����*l��\�U�Oo�M�;��o��}ע�j<Yr�XqU��m���u3tx�5`�.)CG��<p���O	�Ǐ<x��ǌ<x��0���Ǐ<x�㧄���8pᣃ8p�Ç��ɻ���j���=�5-u�G-�X�7��[9]��W�m1zx�Qȵ��(�٠`��H�A��Kx2�0r�죢����Y��UھC� ��PQw�O�O�����j�G\1]C7g#�+�ML}���M������HJ@u	|s Z����z��,�ʓzW��Uv�ib߾0Q���;|7W$�Ύ(#ї���ۗP��p�u�t��]�WV'���`��g��z6�RAd[�bV��)g��Uo�is�\u}�.����Τ֋�q�\��N�0�A����8]+ .�ҋS}r�u@�ܣN><�[˝s�˷���r��)d�C�0
�X3�nDG����F
10�ۗu72Ո9e$�սa���w��L�q��;GZ`�]�9+�eI�S�dǜ����;��hM���)]�TX>	e���H���y�Z�"�x�F����=�|Sc�����p$�K2N5�av��n����s�2:�Wq0�X�mJEݷ�$��z��/�R�2��m�Na�I�B��21ؼ��r���Q�2�9��N�C�V(�Q��Nq��44�w5���ʑ���a/�]u��J�@��н��/���nw�FwUn������B�r��(��<*oWu^�S�oe۶�E�s2i̊��VK&�C���5vo�h\�f�[h�R4Q�y����dt:�ٚ)U���+�?��������t�݃�֞]�g�8�{:�ӅK'���L�;�s��hm;���=;�r�uN�Ѓ%%^�������@�f���R�c�A��m�������v{٤9�G�'P�O6�Ij�s���P� 6wLj��0t�uT����8���]nRXt����țJl���R��b��\D�՘��Zj�^iV�^�s%Т�}V#RY�f�N�|]e��3B��_�+�bf>��t�彰��e5��g]g$�gͬ���a����b
Zl�!U·Y���k8�m��!*�e��!]��k -����!�2��eᵕ�6�#��\����>D	����|���zZ�jm�]3�vP��̧U��l	J��s��[�,��:*0���It���WV3��$F�ʜZ���!V+�P*�&�=�T�*w�t���G]� ��Һk�
5;���qR�N�˸�ĨV�uI3Ot:����HU�����cV66�^1���'G��˖�L��	��J��#�]�K\9/Ղ�;b�n����ѫ^>�Fî��\Rr�/
t���յ(�;S��<����H�������;/�;ٰ�!��X���6k�����R�û������>��>=N�Q���њi�ÿ�W�m�?�[�M!��a[t%-�[��+�'u|���@��v�g�b�(.��6j�.s��fb3��@>��+ث���QWaE-I����+7T������]ݷ1fKx���]�gt��f�
?gL>|������b��ܧNzW�o��������Kԃ�|��Y����N9՛0msy�WK�/��5Q&A9Ӌf=��H�W٨7�.3����2��&&��U�
���H@K���!B���]���KP�߬$�.̢(2�`<jC�w4V��4)�xa-m��JP��k�x革���vŲ޽�u�j>�p�.��]x\����q���oml��S�G*D�gUݾ�Y|aN��P=7o�K�Wt	��+���[zf���b;Ss�	��s�h�v+l�?W���Z��q΂R�}����,]��P������/�Gr�֥V7��v�1�b%U���S:�>��-��g0Ş�r����3GNX�&>2��*�ۮR�����E��x�yr�n�mn�S��e�\��]��|�V�ͩ4��u.����[�ˮ����PW9s�[u'����vd�����ml;)R��,=����F����rf.,�����:t�������q�n�het��\�����b�����s]s��A޸K㢢%���G������j��ʌ" a�ʧB�l��Q�E�T�Q��I��
r�2�f��u�O��[۟s;�p��fe�is3/(PU].-S�Ʀ66�㍢\L�D���E0��C-�-�Tn�5M8�q��������cj��iL�p���`�j܆�Z�Q�Vꮚ!m1��t��r�LJ�lTk�T5�X�`��ճZmLE0VJ%�F�8pU���kDJ�R�֦���c�c�ҵ5�J�uqլR�9�T��J��j�ZV��Q�����8p��E-��.[iE%o֙��X�m*LJaL��쟩�p��T��%S��!y��h
8�F�4l�7�`�}���S3)��B`�`�(�+�m�J��5�-Xhp�-�~�m�]\ֱM���3f)çM����4Uq�Pֲ�5%�wpM�y�l�u�h�u���֣��6ڗT�]_f��xUۧP4(�[���L3,�43NWRK�f���3[)�t�V��Z�<||r|c�L Jex��W-\�nGkD�n���i��)!����4q�Б�+�0Y����/hfX�7�5�f^4d����B�i�u�T!p���� xp�?>>mi�ⵄ~f�V�-j*	�+2л��\��´%�ц�Zњ�	�:ӻ�*Բ6�&+M&:Y\mֱ�n�م����r�gf�c�ԩs�ݘ|x��������N�&�.\&j��G+�&9)���0��\��(�aj�~����=�f��q�K�����je�\�.���u���mE1��F"���^�4��0)�G�UY�w�m�Yۖ�+QKsk�5��o'n�9��q�©�.gF��up"���Z&�]\7zF��s,-�A@�
�do�>��OK�
��z��9�~3����~����p��G<��qgc�L�����f\�ޕp���_ۚ��w"���S�WQ/��C~X�R�)�nr���m>Ͼ�j�����Gh��I�\��|��mh�����Y-M�k�OA��e;Է:�m�}�����gf�Dֶ�-��<(?WHk���h.��~~�"�l\*j���z�C��;����9�}y:N��Ͳ;g�2�K�E�8̘�m��iηG_YS���Nzw�vv&���4;����";[a�z���R%��	O�3����
�Ԗ�������Gt�ݓ{,��!�C�̃��f��J���$�3B�1�~��ptvH���� �Ǻ�d@�����V���Q�LQf<}�|ף��ia	FW._vyq�5]ƶ!�]���O��I�*#IKt2B-�B��[�B�'��V.ޣ����D�]�(<�+)w%ܫ�G2'Xۻ6F���W����-Tzؚw{[�'t4'Yzl�7��U��$�[��+BZ���u�o>�.6ؒ�ݠ�]5j_#K{x*���W�U�q���Ϛ���V�(r��G6�2�EH9�H�fs\f?�x��j����}�+vw|Ѯ5k&[�ς���'F��63���Q��Ƭ�1c���=øp�osv	�yl���[����r��O`�R�9�_�ō�e�S{�w�����U2y�b���Ԥ��to�v�yW<	o��{i�HV�z�K�W?����^�2xk�-���}M��s>}��Զ�*&��DY��8�7x��xcx{X�ǤF�����C�S�o�9��IB�	�ez��X;^��%���աzo�=^��c!���/�|�*[���zM�6�XLbi��:����W�t̮x��oL��Ŝ�����l^m��	��<I�}���s:㩄�$4�hk{�3��)B�}U��_9K_��}ޱ���ݮ���c���-Hq	b���Y�	�٭ ��hq���4�@<�n����h��q{�i��J�ac����C�ֲ�ߙ��xڨ��k�{qpGi�}�-�c�S��K]O���/�N�oz��Q-T:��ܲ�\�P.�����b2�]MТ�:�:߲����5�G�c��铷ϋ�a�n�=oX�g�<K^9��ö�E����t�P�齼k��F럮�6���j��2�Ӌ�>{t-T9/��wyw�b�ۗR^ԧ2�K�NU��3"��2{ݎ�'�����ey;�ݜ��ȏ��{t����v
~��)�����tF�Ǩ�>��n��Y�/�X���J4d�U�r�|2��pˮ���-��#.��_dֶOg�p��}��\��i*�-�&�>
����렁y~�}����[�����B}�\���r�l�;^�i|B<����d�vkյ����q�rr��5ּ��	�DHy��ob���z���2T�����ʯgR?Y��y�d�E4����y5�TӲ��z�n�Mv��4a��t�2�s�^�n�&�vU&�e��ѦS��{V����iZ�����zۅ̗�f��q����+�K�J�����7Vؒ��V)��v-_��\����l��(�#��.�t����j�wN�@��8�Y��f����X-�\�]Ԧ��:�I��NR� ��UeUWkJ��h�ۜ��ݳ��V�@���E���n�IW�W��:�{�>��̩�n ��&����d�٫4�j��Uռ�9vNn����6��}���;-���t@�L:j5���v���g-~ڇ>�z��p�M� ��;�,�8�-�x�v\sj�Ȓ�}�I]��N�S������σon�o�6����㸷T�s,���0t��f���g�d6��aN8X!��I{^�}��2�pj^'����9��>'�������k���׵��A��s>�3>���9�,�b���T��Ȧӑ��U���(��>Ψ�L3���c��wb�;=j�����U�}��9�ٴ9�i��Q杁�Cl�����ll��6g���0�WggO��E�4���Y\��uN���	�׺��Ӳt�8e&s�m���ekC�х�V#\%tW��/�e��QfXF�V�E|/��5�AaɄ=�;��V��&0��6S��+]����f�=G�>VmA�N`7ݦC�}\�>+,_	��P����T��c庬��a ��}`��am�I�\E0���ei&ªp�ܧW)
"��t�����96R�{��<��!ݽ>]\�,�<k��7��閛�"H����dm
x�dN�8*���I��=O��9�y�b�OFq�փ����N�y��,tA�욊�������OP�����~���{�+�{Ƭ�=�+=&F�9���c��7���;I�뒡��чM{�'�����|A71�w�j)�4ԛ�ϛ*�8��KO[�۴��5Xn����8�mί#��f�I�=u�W8�3�b6`����;Uz�,F���G[�6�hgF�{|��y�����7sφ��oh��l� v[슶�ċ�{m�D{o�n�'l�iq1CMIzӆ$���u��0�V�$df������G���׶��ݗ2l{F����<�p�ojs���A���4:��@ �3#ż8��ە��l�ƴ���E��9n�T��s�%���������[Ƒ�vU��W��(�<&)�d�e_�U�P:�H'������h���T-wm6C�Y}|WQ�V����T]m'�5�'p��%�N���cW���gp����W�p6B�3�W�ן���G�����=^Cpd�V�p�45�$�ݕ��$C�ق'OD��ʮ��wLQ���S+������uķ5��'���VW�վ�8",���<�x;��mٻ�,�d֐i9}����%o��g��]R�uN�=�)�{y�3���5����'L����H\����>��Gl�=A�40����q���J�E D𥤗�7/`T�Ʋ��7�Leu��^	4H9$���F�n�b8�0&�̚�ɮE��,bʩ+�@6�K+���0=��?n����8ƈ��WeǛlW�s��W�/>�*�U�S��V��mJ�=�]��5��xa�����x-���Os�	u����U��fpfOD?eL�x��3��<z���E�S��K����w}'�f�׎���t^{��t�6Mȍ���1[ѹ~��J0w�L�׊.Vq[��Ȕ{�#���\]�QvTF�d$�ܗ� 'J3�������pf:V�1��%��3���;�v����ێ��\��9���DR�k1g��f>al�	�C���Z#��xfM�;���7r���J�����Z�Y�߫�V�t�Ҭ}�W����OϫB���j��JnC|[�0�o�����q�k�"�C~��j�����k�_�;W�ݝ:�◟nwK�������x���q7T�l�#�R�WLG��z�[w:6=�6���Ǎ�e�c�ct����6{w��C[c���m�\�ȼ���s�iP�t}��2����v'z����<���N�$]�Vs���`�ާ��B�/�n*�ը�=��a�Н��������1�Y�V-J�v����j�ﯾ�j���]HhW�?�1���V��st�Y��g),�ii������o;��Gn��M��ꃪv
~�M;ڇ%�������^�������~���9Q������p�5�5|(�����7Ch�5�	��b�]���\��q�=\�vN���Պ��:���3ǽ��4U���ܮٜ|Fj�_�|֚�c��VT������0iM� Ks0�9a-��3����k�/��L����VVg-���[���g��+!5��r��\z��=;����C��r����ו�CJp���=}wR�W׺{{To��ؤ|1�q{���v��d�w�յ�]�N��tz�x��� �:�vϟx�8/��P�{(g{�
�?60I�]��-�ͷ��{�ǚ�s��@D
 ���~�~x���g�	
��ĒyMYJ{�?<� '�7G�4T���S�z�q����T�QrF
-w�ݻ�遣���ꪛ�.�f������M��=��5~����W�����,ٷ��_1�w����5�q����hY�&`;W;>�i;y��� æ��=�k|C��9uy�"����A�	�z��և�ݫ�ִ���#S�n'�9���~�>��,���p5��#/^=�$�ǈ�!��۴d+/�N�zQ��Z�;�<}�Z!�P�3�\�َ6F�2;1�㌼���g�ݵ;���k���r{+�ط4��G^�<��&�g���������,j�gېQY���Y0��qu�ur��jx��[�Ǹ����uO�'�D��{�)�'���ǝ��U��Tpl{�>��<��Ѯ.���Wv�]��<��Ԃ�3�r�W\^<��wfpٜ�c�4����#'M���"�p�U$�P-��0QDg{��ok���owbG]4Ot��<�gmy��z_�{��{�!ԠG��vY>���k�Ğ�v�I�?W���D���:�9���g"��9zs�?yP{�}����X�<~��:����&��+��6��:�\�N�>�Y�'?��Sڵ7�E�^Z�׽=���wV=��6��;��|jdd��bP���P�����^40�Y^5�M�)��ѫ��lh���'�N6
���m�ip���"�m����Ծʾ_�t\�L�萜{���o���7��g��^p��X�O4xu�hzb����:#�WCݓ1�|��śj����s��Ǯ�ZGq��7�y����X����\cU�P �.ss˨��p��5雒��ct�� ����kHͨ�:Bg����P�/rs���eΨ�󹾲wё�A���q2�@�]|*��[�:���'_&F�,!��T���ot �k��l�Y9�d.��.�y���m�ֺ�s�W���E�p,ߝz�7�ix�Q��aD���+�Y�ݛY�(�i�j=Ś������VQ�}8Z�ժӳ_�Ђ��L�^j�l;�h�$��p�G�qJ�B$I�yk��t�6�g�z�u*�g�P=��	��`�f�t�u<DB���@/�7��_6�ͪ*�m/{ԕa�^���ܞA��^����/����<�/�-���m�>�L���T�s�8\�[GT� w�/�m.hr�"an{��A�;��I�x��&E�6���N5�Sר�g#gY�{K�^V/4��(��ٶo`�ay���5�t����}���li��-�=��t��U���s3i�'��{��2~��vmI�5�&�yB:9.ag�;��|:-���4X9a��f�E������+�}����5�@�1���3v��L����e��ͣY���l� �YL� �����lk�<�JE���O^h�s���=A�F�k�C�_H5[^x��(��s�}����O��=WܓK��CQ�h=����m#h7@��d�nt��@?�:~�����n������YC��RB�sӨM�:��Rd�h�#Ŧ.���ML���l�:e���)
4����TfV�.�pEGDe�_R��4D�q�f�weu=�h�p�j!L�!;��7Ӯ�ad�1]f��/kP�5�\J�T���1Mu:�܎�/sL�xe[y�{\�I~k-��F</[�9*��8�ݐ�!�j�zm�3���N$��v�־5)�Sn�SM�p�ֻ�s�=0V���;>X���TԳ�%G�0Y�î�gU�����R��o'N�1Ć�ޙ��¢����F�1�ڻ��47�w�mKsN譼<ba��,���ӫ���Yx��9fp���93��gh��4+ݵƺ\md@�bQYս ��Of�@Y����tk&�n=�[G��f�	rږ�ۻ���=]u�3��ޫ4B{��F��1�|76�������%�-Xח�VH,D���o���v�����F��w`��/�;�V�=Y3QW(x:�;��̼�N�m����0r��a�Y����Al"q�Pc3�Śe��h�;�>�&�I�i�v�n�٘��2v�]�M��s
L�<oh���3R��.��P��S\�B@�M����vP�#�=[������STI�,`�}䟬���{[Y-�nY��[)੢�r+Q��S�poSۤ����3����ݺ �}LgVڠ�]1�u��HY�O�;����e�7k�¿'18�<��YA��b� ��l�B�~���+1��/r3�l�6,U�o��e<g$���(:���K{���ղ�k�3y������s]����+5���1ע��csE�v5�j�:��5�,���Xf�[���Cb�;� ��z�B6���ᕰm̾��}
M,�k��KQuz6���6��=�_����8�ʰc�5r��c��c))�&Y�Lޓ��aG2ɖ��1c:�WL,���Q�n_.��1��KfP��#�)PD0Puy)�-�C�������6F��Vz��9�lۡ\f��;�oX�fp�;�V�;��e V�ʰ��w�5����u��z�FY��qww�ŧ.Ɩh��>���8�)��t2���w��n� oH��_dH!�����D��p���]�`b��807]�5�ئȆV����4Q[�e��w3\�QIF�OS��/F��SM���)�Z��R�Q�rc���#��d���{���e߃�Ua#��C���/(�6�)�V:j��}3�	�y�Z½�]�h������23����G*��hߎ��v�_�t�0Z�ECVy]$��W.Twq:듒���sj�
��WU�u�;:<�T+�-o5�j�ӓp���LN�,�6�	L.4���gqǙ�Τj!���j���-Ӝ%��Pj��&GWm��z���[|�P��+���f�o>�����k�V��Y��Qfk2N���݈WJ�D�5Lq(�e�?-�QF��E��y���e)�p���Ҕ���EX�[aX�.e�!X��EWҖ�ږԬ���h�����f�M�t���6|l�ÆsS
TZ��ܵU�+,�U���DT}aF�eq��[T��)��i>8p�ݩ�EDt�-�7CMM?�������jcmU��SAfS����m�R��0���gb�6��,�w�SXe�[Z�ʮ5YR=�juK�B���VQX(|˃V�5tS���E���m��
�e��3%}h�4�5h%e2���X�D����V[V!�3F6r1Um��Je��fJ��rʚ]]f�u���b�
[uf���L�f�m�V�0�����j�h�o��(��fJ�5�)��lLv�V�#�� �iTE+xp��g#YG�SY�I�&6�YT�-(����"&2b`��CV̹pu��O[&�t�Sb\�,%T��KeF۔�
bfkSIu.�-k+� �7ji[�g�{5��m2���z��}f��t���P����h�]�dsn�e�.����hYn��\�KY*� �v����'F�_�_���A�|7k;w?���HM;�O��IUVG�����z�4*#�m�k0�@xXkb�9�������z���$6�w{M3C
�bu��VPCLp�p5�<^TtK���������cƵAt��#�&@#�4�F0�6*���"���5%^f�e4���\�n_[�v�lؙ|��w�t0 ��H
�+��`l�!�c�a>R"��;R�n��_H�����8t=�-K�k���ي�#{;+Y�!���ۜkO�{~�D{ڮ����x|����_,.@� ������(Qɼ�ɓ�w��G��bYy�=��W�KD`Nf�r��kDF��[�0�Uk�J$t����[��ߑ�ʐ�*���v���F03�K�KbZ����Zo`Id��3mq�<����_O��Z0����ڽ=����q̽�͑i�}��x��>Y;v˖��E5� ;"�9��N�Er�����7��̢��/���h��ND������wl�zK�<���}�i=8�?�G��_��ɱ�|�ة������e�X��K���a���3#��P��(׫f����"���t|�G|���yax,��!ϭI*М���#J<]��X���JN�=Y!�r�$� �{T�4w7T��3�i��	5��4�Ł��"I��#�"/s4T�3M�O��8�S��]F��3FI��=O���ѷ"����U^�/*W����	9a�~�C4ćj�����"��[��Zވ��a��x�Ս��F��f�֮c}��y�^x��0����i�}�x�O}xe�o�dl��(�93o1��1�,��#,8�V��=>�W����	�����A�t�=�^���Vr�/��#��GK�B��j�|�{��
#k�δ:�df�Q" 9\b���r�_���U�m��3�ym�e���xi�LH�(�Ї�i1���遍��v��^��ЊϨ�P�1i�p7zo���깭��]���\�Tb�[�(�3!0=q�a	?6��Y�]c h03.��ovk��;q����l.*���j����{��6|kV�ˉ; K�h6$Uy��ۋ=�����7k�������ma��7����sA¼�����X<�,�Ȣ�шYMi��0	��3� ��=0�%]
/Lk�Mծ�C�	���L �[�����"����Ѷ��T\.�6Áz��j:��{2
�Y����AZ�D4���}�����R�`�V;��i���)۪`�F��o��mp'�Pw��)$vN!x�KK���w<����؍�k4�C{��Sf�\n�{h�=j�r���W���c��V��kܔ���ێ��l;�a�h.�����s��)��Vv��ܔ�	��9���;9�ۄ_e�gK���}H��]�V�(IN��b)��P���� ��C����Z��4�Ⱥ%�J:'rx����-�]Ӷ�����U�-�u����׳�/�s�趍qE���Xn0�G�w�� �:f�	_nҔȆ�	���W���Lkhլ_{����!�J��A�/N�o�r �cO��`��Ӱ%��$���t����K:շ�ʐ��6��fۓ�`/�G5yё���5��KO�f6X!�\.uA����|���{�7�e����^2��|kZCyq�B��^���E��چG��YU��b���t?_�)����+*��;]��u`��d���>ﺝY-���˩��v�kU��� A�˻7�l�T�z^wy�̲����	���7�VI�~�W=����To��lt��F�kEn�(��~�M��/����Z~ ,k�L�E��j�J�6����vh�8�e,����U׏T����/�p/�E
1
�t���=�#�K��ޒ}#}#0�͆��m�#��-����l3z&g�=�T�����?2W���IԷ���pT�Er�z����zY���EI�xr����c�>�}�s�y�gW�KZ{�爀kxOk��%bhT{(s�Yov�Zs��P:�����������*w٣�J2��X��Hr�p�@"/��X'����4V�;��x��d'�k�  Ԏ���rb�0�hN�7 ����5��#�"��������t3T�@�q��EXՉMm<;�$��կLm�c�n����/����*�X(3��q�髦/Dǌ<��:��`�Xâ���P�T���sE�UF5Ɇ�6x2��"Pg���
6 X���E0��Z�V�Օ2sr�:�t?0@zg!����oL8�=�5���L���!6h�˯���MJ�yuMZ'�6�chű>C��x��V��4�� l��4'��B`$;'�7Z�os���_Y�؈�f�-�럖�ӝ���	�)J�؍�ǯ/b���ؗ�$!fM��W҇�n�Q)T ��o�ZƜ�y��M�'����S�Y��Ki�آ�st���b���&-P�����r@�d<h���'�v�=����e������̋�K���E�;<��`p�z�H7;56׀ޣ'Y�u�]o�j�:tB�6U�!:��+��އU�[b���kM��3�c�i�Z���o�>��A�B���#ü[Z�h�hLzS��:�մ��2���ԕt;�����Y�B��w^����
�W�4
��p�]x8���Ijc���m�b	E������	ϧ-��+3T��(�4�%�F��{�R��[=����[ƶ�`W�0׃�:�C�Vv=ָ�<�"�IBc`��}�=��}����l @�{3E%�D0��������" мF�@A?-�1��t=U�˿5�=]�EPI�1�z9�)��ݎ�N�z�ˏ�n�Pز��4l��_"|����'֤e��&���f�~=�w9Q��FW�[bǍ����}���1ѵ$��`�ځ44t�k�
|���;}��M�lqUuw*�Bi1�ђ��O'�_�_I �b�$�-�P��Nĥ���y�v,B9R���gnk��@��ᢵN(K;��wJ������;����DPo^�k9n�q{v(�{��y��3�Y�G�μЫ6o�C(��X�"�u�z���{6���X*� �lŃ�7�q<?B�'�6�����!�24t31��WˬUOӪ��,���&���wt5�^�ku{��/���;X�A;YɄ��z�U���ycG�:O��\zL�	p���7�e?D͸,�3 t(��i7����	��g�Af�G���t�;b�Y�_G,��%8�L惢��=q�,��r&�$kmoK����|@h@Feb�4<;��-����.�:f��"�x'��m��yO�]���VZ�ɨ�B�Ц
|F<�r؆2��/*6u��Įc[� �rw㵴��ݽ�$�����V��"���[o�g	�(dN�v��I�YsT;Y�����W��a�J�ĭv��2H�S�P���O�ʜ�\�z�u��ٕ���ү�K�A!$	lv�x^�T�����FHxd1;�ڸb:@�j��-;{"�μR�޶�G\�W�#��'�u�D��MsX���أ��F@dG�I��\�J 9ܞ�$��m��5R��Ȧ�g���)����(/���fX�Q��<�zZ-��`�b6߄� �#ry�E��i9	�^��-?0G0f��Qlnx�69n�c�f&��L��d3��.C�q��DR?~�6s�����x�[����J�6]��z�	hB�F���Tw:lH�������۩��	�>N��c[P���3V��c�����|XJN[�O'��ʦ ��Ͳ6��yL3��f֙ȃc�7�u�)��z_ͯ��Z�a��1��~�=^��:�Ǐ�	|0u�G�`�soF�V����u���A��:e���T��,�n*�;i'���0/ĉ��oU��n[q��ح�ncsp�`��Gb�,b�R�JaQF�p�*�?<]�ź���;�@� ���@,Ō�x�i�e��jmȓf���R������r;�C@�q�1$JwV&=m�7���f^Ї��eFJ�D:�.��^)8*����v=;c5��M@��R����5�x���w��`\P�b<�Fu���U�	c�[{y������E���VJ�5�����b���n�&���+*	���'Pe�O5z(��v�5_^�ɇ�*%���)"F���� @���}������o�f؆�L�M����sͼ��	�#@{�d_�Us�����/���x)�n���xի�B�h:w�>��ӅP�M�Y�#5T���X� `��gzˬ���_;��d��/��U�q����O���>�]k}�� [��wCΉ��7��R��i�p��bkQ�U��*���%����)�X���n��F�ۜ8=�q�_ ��=ۛ�Ug����#�?�2W�;Hܗn�,頶d3aw	���o�Yx�{���������[�f�?|��N�������8��Ħ�!}��\#��� ��^L�myaB��=�8H�BZ�Z����,�@��A�/N�o$n@A¾<���@�@܁%�!��Mn�_�m�n�˯r�.������K"�xdc�#�WzkU��RV~�,@~T!uT��)��ȝY�e~[/g��TD7�C�2M
Ų\8�9+�Z�˔����������iV�8Y��s�8�io�18H[�
|B����K�:�[B̀bN��T��nʳ��HOv����2���-,ڨ�ySMM^	Tr����@ �4=��<�v�,:����('[��|��5f�E��2�+�Oo&�Q�����W�uE�s*������mRU��mw9��:�O%[����b^kL�R��3Bd����������_
I��
$DB#{z����~��V ���ϡ7S�-"F��ٛ���1'\u��]-(%�T{Xm���\9�����4�hTX�a&���# GĠ����ˡ�fg���C<�����q�ڬ���V��rW9�2�yʓ�]�-�ʁ]�"R��tP1#D2 (�a�����{���	}��5	-8����Eּ"�F��N�{�0dw�Y���H¥x�T�g�3��
Z�9�,.݃:­�k���W���@�e⻤"�BA~�ҏx")=\&�L���	X:���Ů��/޷����&���X�5nF6c�}}�U�B�4={#��	^j�������X���Cۛ�_af�>PDc���#��n�1w5��Q�����kj������#�B����Ty����I᧢�4jɞ$�����3���� �-�#D�i�ϟ>2Q���~"Y���S�z��7/�^����$�byV8л��s�҃t���X�e�%��HvO��uIkB���]�{ݻ8,ޭ�
���ɍueI`���B�b�`^�P��H"�-�~`pk\�����B��K���+�61�3m�M\���h�8(;���YO/`�..V�@���W���|��u��䯘�M�6n�֬�݌^ J}��#��n�d'h���Ⱶ���u�f�G���V0�|�r�J�+��w�i�DP�X�����F@D��� Y���V��d0}ٔ85x�I��,�^|v(�nY�j��T<�bGA8��l{�^��"�>�9�n�Q��!�zu�J�����]0FaI�)�>�wGGR�_$���nN(3׎�����^�=2)�ƈ��`3�����WxwR�����Z�O�a(,hj�����E�.i��������:C�*�D}�E��(G1�16�T�L���u�%�g�V�hl:��Yճ@=����lf�!=Q�xy&�dj�쀄�6C�@p�_�b[̖�F����S�±�l�m�D��*.�`��{��w,�+��<�Рz�Q^��-��h�����r!��2춊���ʘ�;���'����?O�}�{f	�T
=�`�:����[#$��w��Yp�u#�Ի���r	~����Y&+�㴬xJ�G�ݔ�0�z��,'(:c��/΃D@d/b�W*�>��~�������$9!��>��۷���c�����ֺ�n��y�L\>���J��'�"�l�Խ[ѱ�CZws��/��%T�5����DP�]���%�����'��O� ����8��읋�B�E�=��^TO�+ف��uwO�k�}=�~ &���VU�]�]Ӱ-T	���(�'\}6pMZ�4WwEh@��*	E>$Z�y�{;$|U�-^J��WG�������}���������H��Q�D��@FJ�H��������91na O�S��C�ڃ#�J��L�����]3B~�Y�Fm�7�p�3�;3Yv�V��^M�-\NPt/z���U�u�)(��|�.>��u�7=x��:��r�g�����]�e����vp�l�2� bN&��Y�\�Ɍ��c�U��Jp3�/ޘw������_����&�w:����#s79	���$��|�M:tһkj���J�����/j�0Wwˢf���"yٔ-#�nnGj:����\�Ȣ�su�լ�k�<�K��!&'�{݂:Q��a�!�O��1����r7'�	�I>y�T�*[�R&�M�\)���ܬbs��/�qm_/`1d�h�@�3��d{�:g���u&��Y�WجB1���LN�^;�1�ɷT��@�Oό����=��dt��G�J�H��WM7!���^b��F�����r,VF��}�Rǡ}_vF�g�H��aD1�:��z�d�t��q��k����u��
���@���a���B�7/�\��{������C��K��F	 1�kp�f���q�
3-l^4C���yd ����)����'YC��)Yal�(sP���`@��N��^�y�8�\��v;�p�9���`��'���uK��콡���i��$r{)��Z7uN�F�<��a�g)v��A]&�Wo���#�^��u�t��r�+�ü2���T6k7)�3��u��6ޢ�r�����3Fn��/on�'�˻l M���h�Z7(9�%cz�~�¤=B���=�R����.huX4j#�aj;�'y�]:,�u��h�l�S�z��6f�F���U��e�ˎ�Wtf�w.o�����řW���$rfP[�Xu�#�"�x4��ЬxF�6g3K�Yׂ�&�nuXД�
>l���kc{T��a�'��+P�]�[�]�y�c<p:�CypDZ�Vi��Tϱ���(�s����#��Q7���xVKʑv3��7�����CY��dݓ��i���G�t]b�=�R[�N�}Y���b|�����[�tN��c��̇�j �������K8h^�
ŹWCb+o�p�R���TM *TK�|�ɧ]4�IWE��V.�P"�uR9��To��C9���KR��׮�q��:1��ޙ���"���{���ݺPL�RN�i[�N��bPѱ9n�tpmu���w1(m^Ŗb�*�{�[wZhH�R�u��a�y�Z��ԩGE�J��R����/nۮk��N��YZ6�P4>P���1�IX��p�q�I�WI^�Ww�Ү"�QsşD�f�q�V��0ڏG[�\�S.'tQAS���Τ�xNv�$�ھ��v�roN���p��N�[8�����J�4��qO��F�қ����󳂌��-��{]B�\��7IK�n4���j�t��u�^�N��kv�/{Y�f%WmiH�P��Q�J���q]�X���û�h�Žl)�`�a�7Q���<w��YZ��Z�(Ȇ���q:5V3x�e�ڭ�ii�4�8RF�xn��`��/1	��c��F<�	3����<�yے�m�C��˭��	�#�Ef����\o\��-5�'Kl�2�,�M��->�dZv�d�h�6m��^2k����h�v�ݓ(s�:�nö��q��lC�h�u�ط������RbJ�wI�v�`W�_%zΡ|T�p�˭r��o�TKuՂө�q����`�4,Y#��e�Gq��p��ǡ�(1׏���R[Q�Ŕ$�o_"�E���Y���Ů��D��qt��l�65]����9�Qzh8�Y$�0ҽ��c3(�]���P��:5�&�ݕ�yg$��-�����-TڮƜd�g&�{"��W׀dW�\I��rG��&�[�>�^�c��.�79�y�����"uh��z���:rxV֥�M�7(��) ^�p*Ul'MӡIP,�IAQ!�F������{�J� �ێ�Z"�f��N�#D������T�֮���?��MҊ5�>qVQ��~����21��Y�Eb��S([[LV�2��?6p�G�%J�ar����c�[���Un�a��(�E�}f1٢�k.a�E4�4�(��ip���ÇZÉWT�P�Jbi�j¢i�-[AZ�ڸٌ��Ȗ����Oܠ�`� _�P�*-EKE~4x�Ç�V)l��4���̨���QKkhq���1հ�	����fQLu�1KaX�
�Yq�*0�ӆ�Kj[AB�*�8��V6�(,N2�PD��SI�8�+-��wh�m�%�:l���mk�a\A��DA���ʸ�ګ�J��娔���+m.�R�Q٣�M8)mb��2ը�m-����p��-:�d���D���m��m�r��Y���O����x�J��EPժuJc��D��E-��%E��E�s)o��*�>>8l�RT�x՘մB�J�AkRƲ�֢�ŭH(�h�V��4��KJ����mYSV�^�Q]k1�R��Y���:d���L�X��I�dŴ��E�h
(���[�l����J�}��q�I
�z�+]i��e��$37R�zEY��&u�=��J�s����I]W��9�j_��
�ai�_��C�@�H#
!"!"22$a#ﾜ����g:@���B8�������a��P2/�z\0�5<Ų��]6��ۜx�۝kf�����P4?�#��㚨J-d������~���/��P:�����=)�P�Ew[lb�]���˵a!���DqF�*�r`c%Cv�k��ēn�j��\�i��tv�.�.��O��G$�����j�P�¿��L����Bx�}1h,�7�>��CB���΋�����g�^��4i��������mi�Q�="���E!�����6y�-�Yz�ům �֡�*��[�W(1F-�Fl�*��Ϲ舉�" H��.z�Q��{}����L܄�r*ڽ�O�c:j��Y9���[J�eE�����W��H�~˳��e# "'�e	�h��O�5Q��v�tSN���)۪L)�d�t�O3��鍅u֨���󷗦^��ְ���}=.FBmrV�ޚ:il2�8��)�{�0?Ѣ,v��-��Ӕ���GN0�zh<D��Bc�l�_��}�ك�y�7�zxf��rb��m��2�He�I�ꋷo� Q�ۯ�я(]:ْ����Ó$��`	X]��v/��.F��nޤc�NO������|]�2ɩ��;nVv	�Z-%��-�4\;��D>s�n�A�ͯ�W���Da "@D��� +�[J��`r�ۤRz �h��1a�q��@AƿC��� �s��V���4L���2����ٓ�0K�Ͳ.���#i@��%�j���!A�:�a�pG�����@�(1�l:��-��Ȫ'uM��mU����}�'�!�K�;�q]�g*�Gd,i�[s���xh�(ulĝqvJ�­t��M��a%��Z�(�Ń���!߳�|-�	�8.=`��N`��������"����:�������o,#\�,�Z�g���
��`�I�%S�c�|K����u}0K���\G�jR���F�Ũ�������ޝmwv�#�á�Ӽ��O@�+��3��)@��xp�D����p��'�D�4h�v���ʙ;��=�5x>POyPޟ�8#��؁��	1hFz��_>֦���=3���8I}+�?�
%�߷i�fh�-�:+��PnF���V?qP��4���Ӕ�9N^��ъ ��8�#v�|��M]��9��xj��׊�"g�O���X�K�m$��e~�13��f6����ۻ���>�W;V�Gq�qǙ
/t*ʊ�+q��J��D7��ǵ�)/{�厈V���0�,5�������=2��_F��龭l,hs4�^���� ��xc�k/{%w;&�̰t2�t��������# "FF"H"D$kW߿�����?;���qEx/V��O)�fw�rEQ���Z�����S���X��kȚ���Y� ���.���*4C?a�����މ�I�w�3c�yufc�ҟM+�B��� �*ZWN�W|���1ձfyX5�!�\��ﯳ�-�ӱ~�s[{��9K �sp/	΂e0MJR�v#�x��ء���@��L�a�m�E��ᥑ���lC����@�X���2R��=[������#V�j�!���1=`�6�$Tj�7���o���u�Y��x������[jy2Ϫ_'�c���ӱ��P�M�p2�"�?$16W\nVob�`��^1�N�4�)����gu(qU�����z��ZQ���톱���Y��2k���h�:JK���:���5��>�_h�M?ӣ�	�Ӵ.�*��p�؂˛ v��|�ܥ�],��A�qO i�ʐQ��#�#�t�����z�&%�T�jexw+��yl�d�J;�2�_!�K�
���{W�ܱ�lYg�:5<#y"|�X+l���-�"b}�l��:�D!�/ģLDռx�FZ,��ד�,8�Ƌ����H	ك�Xڶz��N��-5�`U��;r�6�����,lKU5�jR:}��7��u&��j��m�f�B�.S�q�����{�����6w���9��}߽��|J !dHDBD@@d �Y�FU�	�m�
�m���I�����'{կc���R�hņv<ᚽ��}��&�G�|׶�/'
Z�PO��� 3f�����@� �/>�tE�n���
Y�a�H�D,ݬ����������}�x��P�����7�����a����e�c4Z�ڣ}y��,������YC�J�̞��Ь��O�V��v���t�F��Xh\�����M��t��=�ъ��{�ЀS��oUj�PdyI�#LeZ�Nf>�Yj�o�5���L�ӭ/Po��g�3e��Z���젨ck!a�P�6E%�H��O���o������1.�SnVT˼���4�"��Jl&d�њO~U&�����U��y������8�#�U���Н�����!
�U�^~��C�$�������F��CU�ԧ�rv���.�yX��^�Sĝ@�؟"rZC��dp���TĴ���-;{"���&���[׎�0z��.͘F�T�j�X�>P6�9�>����(��n�K��E5��}�Ma9^�|.
��l89�G��q��w�-HA׹[��������X,W��>�\=�����J��9���ܪfT<��C6A��b��y:ꖬ�=���郗A&��D�(ѥNu�nٽi\�ڎ�a�	��6�P>iW�D`�`$H� `���B"����_R`��z/�,���b�"Xb>���İv��x�.�&HY�'a��%Ы��u��ܺ���$(�.h�3L$����$8�!p�$���wFn�����5{�q��u�v����=�M���uPbCg:i#
!���vWH9�3.(�wP�b+:������#օP�{S�E2�d�5�B��C�r!�+�G�T��l^�m����_�g�Lk��i���X{d+��XX����Tȅ垮�O˧��=?<7]�M�����yEG�M�� *Pcy���^��:r�"%G�!�(��c%�>n���;I86#4$@9Y�g��F�x�~r�T�:4xR��V��	Q2#J8�b&.���Cw�a��h�BzK5M��1��f5�doM��nS�"���x�trB@��U�mGW�JP�`,阘m8TrWuΖv}E��ɌV��kB�xhE�'jJm�j�#(ͯj�M���K!,#F^�[���=n�:����-t���o�k�Ch��`��|�t�p���
)���a�[��t1���nW�[�m
����SI�e�Χ�k|�����n�\\72v����с��'����SsF�P�`����w,Z؝�{9f@����s�Y4خkp��v�.JB$޻��kOs�{���-&��f�{~��}�����7��	�20� ��	HA�?����P)�#q����L(L�����ơ�8'���A9 K*�z�Ƽ�=�zU�T>���"��-y ��б�ʘ�FG�|Y�Q��v��tS�;��)���W
��/l�]4�<ыrFڋ,uE��TH�~��]}0�3�tH�(S�ZJL���7�`<�y�"���c7�F��ƅ�)Z�qӌ$vE�u�������B�p����	\���0d��W�gK�r�^�YZ݀1��;;"��̌�;T�*�,�bP�!a�H�3�[1u	if�[��t�y�ʱ"�X~ڃ#2�����l�O(g=c�����D=�;�*x�T�����ɬNڨJ�][O��{i0������OW���4چøm2�n5�nʵ��nu:�ç�Ϙ?7y�sr|󮫨г`ĝqw�J�­��Շu�<��!#��	���uy��V�W�_֭�g��g���g�Ll�3�h1&�qn����.9]ηL�>��~��׋ʏ5�u�pV�6�z�}a(z4Ȁ�רL	�����d!����D�����Si���ėj��'�)N�&"X�K	��u������(2RT�n�St�5�'c��ܕfx���D�^���Yh�乜��艾8�9*&��S' �5�u�bX�we�B�p�>}:�$[�@���f78��y \��W�.����rH#	�HBA �B"���<=�Grr���]hv�5��������c���O�u,@�5H�U��E}��~	��m���a�g��c��ξ�2g��'���dw(�����zf���=Y�0�T5JP�@�;Wռ��|z�9�����]�V=��nb�*Ws�C�*>�e�A�ʺ&����lGO�[���U���c�`�!c�1�?Fd���W���Y�O����\��H �oA�����K=��}ݝN@�aT����+dP�����xYWUklNT�AS�!�_����w:��1
�F��9�3��� ��͑=�7	�آ�`�p��@�F��maog�'N�/���F��B�^l�*{�����Nmu���)�u�B�v�yP�V�ȥec��a�&C��f�U5/���z�L	�������%��z%�m��9n��-w�V�¿g	t*¥'����i o�x�w[T�5hѐߌ
�� �-�� �d�O>;bl�<�2/��\���.�%E˝��c;o*�]eC8K�P���������4�jVv�{"���>M��f�}H��6�A���܅k2G��~�=Et�2��^v�l����ȶ�.
<C5�����Gg
�js]�k�-�W���V�g[Lhz/���y[s��|:dY`䮣���N�z`I	�nk��тHY��kN�f�����}�s����{3�!?� �B"�A�"x0a�{�d�����O�,���[�a�}	M�&k��B����6E�:�Y����ZI�T�[�r٩Uŭ�
X򥥥�	o�Y��t�ϊмw&'������h^�f��;��j���oc0m��u�&=�a�ٷt7U ���H(�@A���#c�����$�e�>[deg5\���Z����a@���~*	{���8��&v����o�V-���^��k8��)ap��Ƞ�͜���1�'���&}:��9��K1�����Q�J���a�\�*�3}��ƤC�>'�O�����7��B=%�H@[^	EzB�šv�n��t�B�4rT$�	�0��1.o��W�������;���	��f�=e�z��w���&�.�����N�Dщ����F���|��b���n�t5Ԡ��`TMl��G�����ˠE{��p�~�j��6���-0k�2�d��U>�y���w���Su���&�K�����Q9c:x�nl�y��^鶫Z�["��E���/h��j i���Y�K'�ܭ�g'=����y�y�췵�PhZ�ͼQs���5k��k۠�5H��P᪍W��69ZY�en�f�[Q�Є����>$oj�K `�n1���X�{n��f}����{f�F�S�bT�|%X̫��:�kV�����	�$�0 � �D@�! ��		���(��8�""2�g�v�W;��!���4-��Nz,�v��j�G*�����.+�.v����(B��H���*�c�1֚a���&�o�%4��ԩ7��Gh����X%`j���~y�駥b�I?�z0#�u���!���G	ܞ�KbZmPӠ�"�)�jkB�"����k�P���u�u���lP">���I�Lh.@ܔC��= wQ������Eɱ���xT*��A�E�E�5x����}��l!#��4���?�����O���e�WNW�O��V��Uэ��� LZ~X�A/CQ25�I�l�"��8��ap�N�
t��B�*�w&m�F��e��\�~;+���&����7ʆ�0��:,TA��v��cR90kt��<T�t��t�Si�F�؁]�j@����������d���\�T��6-ݓ�k���� eZ���9�j�E@��&DyH�`lsV%�^�n�9���1�e�`�>�S<C��^��ɨ}��P�{���G�D'SQ�2��g���9T� ���������|��0Rʢ��J*�fo]͋j�ߞ�2qF�|������*�o;3�t�`��z�Z�P��n��]2�m1h���)nr�_x�-�=����V�.��h���e�M�֩ٮ�WM�y`�{�t�OTS������᪬e�n���X��_}T�KK!"$ Fa D=�7��  �,p1��m�C{�ò+ƫ�F&o�FB~���q*![���Pݠ��br_x�9��[ӓQպ׫m��Ej=�%/z-!=�ʵM���I���3�L6���f=�`�<;�U_^�Xկ�t�e�C�x&v��͖V��k�j�M����2R�t�xv	�s�oTΫW���f��r!�y��G��ݬia" �t�U2�Fp��M�Y�kt3!Z}����Ȳ*�n{�8I�"�w��b�*f��Sf����5_'� �}8VH��˕u��S[��U垹�
5�̀ʌ�����<�P��F|�Ƅ8��z�z/�E4��\�y�.��lX�60g>7��̱��U�Q��s�eT.#-aR��Eצv��v��	���%)�-�42�4��-T�o�H�!R��e���'�a��^$������&�	M�&��vCB,��}����q��o�̘i�5�?����gH�MW>�b6o�9J�d`d}mƉ�"�ʍh'#o���=j>!0�<�� S+�櫖�NT�D^z�"����l<�;O�ߙ��^�UZI-��F�M_:�[�u*gE�S�c���C���؋���J_e4�<�}���Ʒ7���f�)j���PS��w&V�Vd�O������V�=���h|2�Ч|gY4�擠�M���P�Ceޘ��m���P4.]�Ʊ��]���j�i��Ռ�;��j�uF��o�t�ʊ�f��.��BL��@�4�T�B>�n5����4M��V��^ڽ9r��۝��ma��lZKa�X�mmF�*dYOy�F�(U���e��`Q�ѿ�΃�ֻ֬X��%A���w8Ut������\Q@����A�u|&��v:���4饆��:�d�	:3$o�uM��3�o��w[��yR����:j�]��F�ө�+'#�Џ�J���㎚v;�+�ֻ%���#��Q����\p����k[�5\��
AvsQ�}]�3��!S[�Wd���vKu�V�-�4s��Q��}�2���v�f;�%�5J�������/�+�h�
�sV�e==�]n��Kf˹A�"�A�l;ͫy]z:��S;�N�1�\X�7R��r��$��Y����.	�*�!NRGͤ�^iNJ�M���I:��"��%<�#p�U��!q�v4f]]�_v7Q�|�GuT,ͬK���콮�oF�0)Y���[�T���)@ݸe��*K�]Z�J�;�5�T��K�����=7/�utM`� ~$�Q7�]e��]b#����d_yԛ��˧R�����&���5C�of��ZwZD���.уC����WP�P��7OAO"�����q�_v2��7x��q�e��q����TyW0.c1�݄6�LY{���c_c�u.3ls0��q< ��\]�kc1���j5�1�����X�B9���V�kz�]��ЎT�LKp����3�a��i�`;}����![s��t�{K�H̵�Tz���VOX��-q!�_t�����՛���<v�pj�����`��3���7+>i�敧u]��gzn�h��.;!�j��1\�Y	��!�����Y2�Z׆*��D�ƫ��ʋ��W՘�Z�M]�tnp�ȅg6F�f����mv���y<u�˜�K9���P�5։��n�.����S��y��p/\&u�7wM7���ONvtTÇ6���gJ����+D�����XUe����i�լvR�+:m1n�W$�{�2�V,d�d��YwFnme><�7r�`�p�x$���,�f�`i#O /@]�;N�[!�w��C�1��5�F"�4�۹��eZz����;>�Ӎ��X)u���)�)�*��k��Y����%��U)O����oknԶ믜`�|+T=>�$�/3�h�/�:��u��<]ъh�ͨ�1���T~�(i4,�b��i�����JkZ,Z�[J%am*5

8h�Ç
�eT�)E�AB�LT�~v�7i����k
�b�
%���Tth���Â)���lDZ�T�S(��iO�`�6���Y�3R�+��4|a�ÆS� =�PШ�F!�Sѱk"��QGZ���|IkR�UE(��S�c�&�x��gYM5���`��U[i�\UB�-h
�i_�b ����*Զ��*kZ!WVf�V�*�F���83mX,.�W��Q1�Ũ)R�b�Ы-�(�Ǎ.\`�V�a���8&[_ Up���2}a��@Ĩ���VLj4h#*T����aRҕF]R�V,�th��񳂸m�(�0de���Q���Z2T,��-.fe�����J�_e�mb%m�EMl��gN&�c�)K���I���J��Җ�PX�LűV���S�l��Ӝ��k�lLF՚�eG�J�����-(�kh�J��&���J����RҶ�(���z���/g��p;�v>e��#dK9C�Շ<{���gw;��TS�sZԝ��7�}����/z���s}�G���?�$� "d$D���>�����2���&��\ߞ���ȇ�ܞ�����Q�F��aTrW<��I�E�)��ۨa �\��l�yS�1�d���� �0���rBgdDw�	S��uK����,(Z��R�x�l���3܏8���,d��Z
>�>�G��d/2�]	���"��u�eu��c�"���Vl��68�6F�#���頖��!}�>'�����T>�	x�z:;օ�X��U�wclDBP�D��z�gbq{�	�W��'MvłyP���%-�����{WS�).�X�\ev7t�r�����f�ܒ���|	�c�C��4�lk���μ����P}�Zb�zsr��,k4#|�B���=3���3�|�� ���F]�l���l�;"��.�B���.+�@�"���	W��{#s �����%�r�ׅI�e��x�-�J׾�/C�}�LZ=+�}W�<D��6����+Q���*M�7�U�fS&�Wn6F�7THI�=�տ�6�q�����	>��5�&�%Mm8&	>f���;�����\�r*��4VA]N�9�^�gI����!#䚃d7F��=X���*����e9��_���+��O7�Ӯ~=��~t芌H��0�> *��}�l��:R%kx��`�WԮ�1��޶���kv�d��j4��gX����:���^^k#�6�7��_��?� �� ���0����`FIC���Y�6�Sh�7��	��`"!�hR{Tr����%_b�PgݓC�Q��%���gK�����,��7{Ln�}��頷���D������j������T���!�dh΋��ٱ�k*}����^{g~�LʷX�%�u��L�DR`\ŗ����ĥ-�3�^{������"��jDC!���7�u���)�\������آ�g�fv�T��9ۯijrZ<�ä��k�	���3k9���7p�4(����*�y��F��cФ\5�l$۪X^zu��+�A�����(!?l:f,G�Л\����0��u�E6r�Uj�/���@��F���u6��r��4��J�����6�@A?.*�2y�2v�aQ*�wBv�AUs[m�&��zW=����{
�A��m��l� ����������I��u����mqD��c/f��i�z�x)F��t}���i��F�'�tX(��]�Ųb����t{�,H�B��F	UK9\���3$3d��E���1�Qz�� ��ym�Ǌ�⃛�	��ӈa�n�ʬ�:c*,�$��S��s������2�&ʺ|�]����`bx��&]��s� ��=��g�w���.v&�p�*#8�[�Dzō�mH�{�u��^��I��2��Xڰ��f��O�\��e{n��k��� C�`FI� Da#! �� �=�����Y,�*ąͭ�`�n���p\G��B�K���7�v���a�࣫{7��4F��q��+�.�A�զ����k�Û�Aii�%�\�u^�"�.oݴ5��z]")����[!I�3US'w�g�3B�����zS~�j�M�2<��#L�g쌌��(���+X�^T�-�wݵ�J�T_ݭ�9��nl�k�eQ�3�mP�V��Ȥ�`B��>��\�,��Z��O��G��g%��^�w!)��NΛ���V��פ��T�����Jύz�xX�u��uC`�,.D@(<�٠�_�sW�!���I���V*F�SC.�8����f�W�)�^��|�+�(�F@��9S�#p��#r{U �%��.�i��D�0(:��y�L�X��e3�f�i���]��6�ܓ��\��(�#rz�9a��;�n��۬���KБ����خ^c`K�:H><;��_/g�.����ژ��jʟa���-vō<���0�Bn���AG"�E��j-#��a�`-��Y ��x�;�^^���'+�A�|]����:�K��F��M��KNͬ��4LB���r�E�p}�罼�^+���QNש�r7똱`[�C��R^/�%n�*Luՠ9Hi%9 �J���ц�l6W[�&�}����9�]��c�$�� �� D@�$"0$���D�C/kK%iŸ����oJ�i���k����|��H�r���L�C}�),(�k�ʠ���tb{��ۛ��lK,�1�BKv�D�:R(���?]��k��FM��)�S#89�[��i�՘f�[䉧PA_p\D�w)�|��E�8:|;MV�K�8Y��s�,5��qk;�O%D�̿vj���*X���	�}�iQ�8�B�H<o/d,Ϸh��Ǫ�t�@�������Z;9|�����Г��Z-q�<#���
�B;G�lxu�`��Np5��rTAUU���+��l,���'`��'Ì�yq4��ҿ
�T���i�<��Ͻ��ҟO����=���5ݬbcS����Q��w
.�@6�5{��i�ѫ�S�2�0Bw9�l�,td�_��Q���d�R�.�|�b�-BA�P��U�E�x���l�f�%e��}��:�Ҽ��IG�@��j~����7,��W������׍�CS�\�.:w)	ۊ��mr�U��e�E���M����
9�&'Q���O�k�����a �_h�њf�y�s-��j���h\A��t.��i��I���W�����;k..�b�YN�:Y{)G{���3�cO�_H�	::�T���O�q�M��}�������]��]���,�+n�)ug��iJ�踟}�w���us���=���$�!��F�!a"HA����^,�6��F�G�#z��U&�j,쪄�\a^�M	��8�_L6��%
K�!q��k�sދ��o,,�;�򆞷�-ÖЭ��"~܋0�l�D�C�O
�r�D�̬�5�UM�q��t8/?�%?<svzYzz���R'����>�.͔����Pn�Y��Qev�w��[�!k/C�/�&�y�,hv���RSՓ6Ⱥ��9�E�m�Z����ޓ�|cc=^ǋv�$vb�ōw)���1�pmu
��H�E���'����=֊�Szz����ʇ1J��,R�;D.= Dy��)��L�t����*��Mr�s5(�x{�<|��:>���+��CU��� AC�F��Di�&{����}�13]kHwT ߇\Ҝ��Z�)�V>���Orß:�"{lO�V��`�|L|8z4��vE�>x&�S�{�ɛa]sj:p+ 瓙�{�f�c���/`_�E��UO0(T.�\�hn�tL7C�Л����,8!�����.�zI��nRa@���	�c�@q����-���x�}�	��#׸�n�m!56�����_��
w������{���� %́�N]yߖ�kN�fu�"xځ/��|�P�GL�	���OY��^����:�5�D͆��.��p-�Pw��|G]gM<��A��=��\<yݽn��qY��-�9�(�.j�7����{�`� ��H#$�B"B {ް���t��Ů��*�~O����E��/�nQ">̋��{���^�=���9�)���Z㔢�c����/��̖ՉW�������QCo���Uǩ.8/̏n�38�T�u�<��kҸ��f�v�+ �DXM�1w5��Ta����I��W����%[��g�����l ʂˡH�:�����umD}4ҁ?Կ)�H��?L�[�5L��꾊���e�Psk�U,Z��	M����U�B�ߕ�vzs^��V�h�E�TX���~�R5����;-[��?<�0j1ΚX�z��"\6�g�r�H7b}9j���/�W��g�xg_��KĘ��V�,�� ��nOa�Ot�N��bY'C�YqJ�
���{����e��w��\6�F:/�F�91C�BW���2%�ܮ�?nErdXF�x��y��f�����-�P�:@����岴�&�E�a�>3!�����vNʇ�T4�gCި��jڳʶyT��d^� ^�T5�K��i�% W�/I��	��<v�'�W���o�pf�yA^R�)�n�~��0�����8�{Y^���Rx�t�R�ҥ�2�Z������O������׷�ǳ%' �^��U��YV:E�:���VL�3_[��(̖R��+�{H�����.�&����}��.�e�]�6wE I�0�e��ZL��!?���2�D`H� ��� � (I?s��{��??8���,q/3˘K|p����Adw?�[����<e� ���__ϯ��Q�H�du�_��nbO��u\l���#�헪�8�W)���pMhB���n"s6�3�}�[^�~�L'b1��ե}�#�����_�F����1�q�c��0�D(��b՝��r�h6�,4��
|���Mz�d�r}�(�_�Ǥ�x ���A��rs;���-�W�����vS�5 ��B�\�(5��ݠv~��F�cZDǌ]M�lٍ[�gC�*�	Q9N��p���(���蒘L���#�²کUk��!����y�f߸��X�Φh�fK@���#&<�ٴ�9�ӕ_j��.0h`p�A�t�{�F߅�7y�fmt�?Z�U?KU�ȳ>|���h�o°�ls~��f���4����_;1]�bEJ,���`�K ,?k�dzr���p�5��q�,��&��擩1l4�^<�B�p�%ۋ�Yŝ�w�9�?��<A���%����<�[ ��+M��B��K�a��.��C�)��b6@4���+E��(^����b�V%��ʴ6��{TU�S��_ m��1q��f��PA+��'o���#ĥ��ȥ�J-�>�;��λz�(GP�<��yb��y�\�]������|��ˑ�e�b�[x���3z��}�}����?�I"2B" �! F@ `�  �� �]듞I�.�| �6����a�T-bR1j9~�#q�=�y���)�{34��렮�q+cz�T��w�y�t͕�M���i�?H� ȄD��4/�?�D���
r��DHf����+w���p��5��:3�bӕ�c"�{�LYz�<�-�B��B}>r!5ܫc�a ��_]�g+#�TyplCnKV��3NJn���-98�A/Z�H�bX`=4¨��m
�MFx�>Ԯ �h�l����^���u�萮�,^HY#Z��Ju�y=;���)@佂p^�b#��7871A��!^�չ�T*�ف'v6l֍�mq�r:�ˏ�_Q:���ͩ�W�{�
���!�L1n��%�A����a'ʦ/,����tO���ŹV��6X�Y�8�|��=/o/eV��_�/�mGg�Ax-*Q�?B��U��V�(/V����w9P���)�!�禈�u�oEi㢗}��CJ*@����&9���.�G:��x����^�!-�rCc�u�*����b��(�BxE�mGW��R�lU�V�)[���W�������Zy��d���' �Go� G&=һ7�Gw�r;S'\��i�9�+�w����Sx�Q�V.�T^O\�k`�	��}����^�|�N�)�]����[��m��O�}נ��ok�E]��39;3���I?�DBA$F�I �$�C������_�>/�����-�����e���(�W��f��|-x�T5M��|ތ�p�zn2w;������ݩY.�,W8*%oǕT���$Yt�U2(�3�v�6'�*�f�ݝ��q�p,�SʈF�',�����f�w\�U�4�Xo�C�s�ۇ]��d?j�'�����mg2�؟	�@��&�N!��Q�9�ebn:��r�ϳS &s)��W0����O�DW'cP��x�>{s���\'k
�"8� 8�_	��u��FTsJ�nLC�owCG�����4�e�k�Zi��;J�q�0v'"�:�q�	���9�;z�cd�&����j(8B�r��ak��F��2��y��ܢd ͞��>���'��k�n�O[P���t��z��S �y�%��j}�RS�1L����Z�%ć��l��J=�N\���/�?�e4A�Z�)���������dUvKԄ��I�Q�}��I��/L�`�jkuM�fa ڔ��,V���!3�w��{��P�f$님*\0[��^---��u���{��,��"��P�چ:x_q�P�2ݪ|e�o�io�0�_u.#�ٳ>�k�8^?r��!�e��M9��L����Bz��&�]%)�39q�ɠ�Yz_Q4:�|"&��+�_m�!nDc�Ꮺa0p��o{'wB�y�}}��S��?�"��Dd���6$�dB��{��g7���g�0�0�2�S�4���W=�x��;@�� H��`�97�a��hz.�Df�U���Q[��&�Z�?v�A\Q�m�C�PT!p��B#�UGyh�QLm���	|���Z������kWjT
n���ӵ�ƥ��ǠYz�{�L�w&/f���U*��3�CX"�F��<E[��ܞs!�8v�N	���a�ׯ@q�����<&��3��TΈF���V�c��&c��,,k)x �Q���ݢDȿTJݑ�6�3T�a�����M�r3�Q��JOb����b'�Y���x���F̎��K�n+����"22��wvS#]z�$C{��"�ԙ���N�(��N	��M�"��{�Ten��3�]D�V6b��:;ou�i��n�@��E�Tˮo��AW�l���*yIL&l؅��&�0���Dvv�6-�Y�[�l�sh~BSe�I91+oaQ�~=9��4��Ԭ���J���@M]ne�uB~p]�>N���?nQ!�#qΚZĳ�X=Ӱ��պ�Bע�0>>�,R(�tl��ZHie�熃Z�T�N�V�)��pX0��u�ov1^^��~y��7���4J[7��pq}L^ֵ��}RhIKm;�1�Uhw�i��״�N*�Ӊ�;���=*��wѤNu7J=�9s�O��'�˺b�)����#յ����ͫk�Ʈ�Ep��L
���{c�}(����i�"�$�=�Gjwv��+X丳h]�7*=x���[L!^Y�Y�l�ycM*Q	B����|�)'R�%�u6୔+�8���@]hX �\�O�rܝЛJ�%�bJ}�K�:i��E8պ˵Q{�����J�[2�����6�\��f�p��E�f���E�nﶛ�ř�4�f��|3�W֢X2�IJ7��B����9�a��۵i�h!��GG|h#+(T�ާ�hb�;�a-�X���Ҏ��	�~-���]F�L��mZ1M��P��z� D�ӏ�4�GL�樮Y�e�F�n=���1լ{b������NGV�ae`8z�������*��i�'Z4�wH���oٕyz3:�0�U �k�:���2_sN��4U�m=�yyQ$E��%�ɴ�Ū��V��:\ۧW����]��.��l]��&�C�%!s�D��;.��f�Џ�ov��:��I�`W��c ���>ޔ���o�.�2�V݅�[�u8�;��qv�u��:g�}����):�7���P��ٚ�r�Mj�ui|ʕ-���
��6�?
YJo:2�s�z�����*(�4]5J�� (�(������-@�.p�4wok*��5�;���i��h�3@���2�}d���FmJ�Gz��OP���R�s���k��=��w�Z�Ć����M�R�������B��<�ǚ��^]��X���r�x���Ϲ:�7��<��1���ZU/^���=	-��Z��M���[u��4�g�Q�ӹ��,`�foh��W����(Vk���-�o��vj��{-]����ʅq�G#��M@�U��j֙*�=�#s�y�txj݅3;�����3�v�-�VsY���ɒ�ϹE�/��T���ԝLg�k��?���ӏSQ����L�u.�hO�Z�.�{>�|�.��d�-�6wu��4�R͂LΜ�ܲ
�V4�Ť%[�ȣ���݁��3�O�Um�T�y�|����*,�Ëz�Z�VV����
��l.�}hl���R�ɷ�3I8)r)�ǥo��6gt-���N���@u�h\Cz�j��ל�w�̉J��7c9
Ի��+�º���9�n�[����]��n�bFF\��1ņ�:u�f��,@��v�e���G��J��Ŧi��֎�ʟF�U�5�*	��h�F�V��:FM���T\�Z�b���B90*�{�wA_M�t�}t���V��q�9gs;ͩ�����$tS��0A��A:$��!��@R-�D��C��&@�m��@��P�Uf�$��4E��"�ʉ)�J�LA��	�E��gfZ�b�iYRQ�V5�UAeck���d*|�Z�-�d��+%bԍ(��ʅ�68&ZVĭ[V����������Q�ڠ�4T*�O���Z5%U�e�Uk�||l��0�XT+[�b�e�ʨ,b"��Y�T�c+��,��4pѳ�yKK�:��U�ӊ�*�Ȣ塃�څ�X�0P)lR�,̰U1*�������g�o�.�c�B�,���֦&	�-�������5Fҥe�1�f8\�j"*�0����ٳgų����30��O��"�F(�!m���ы�q��a�ŭ�Xf�1���3N�tҸ�\�E:l�ӗ���QEZѕ��J«�V��jJ˙�[U�m��ZaÆ͜��3�(Y�Md�Am�j��ƙ��o���*J�[[mekF"-�o
l�񳀫m�
ѬU���ҕ�˦1ի+
��*�7�xR��\J�-�\
g4`)�Z�)m-��1��^a��͙��:���X��v�>���=;��������L�����ڵ_R4�M�l��x-&��e��u}g�jN�"wm�iarõ͈ �D��5�]SWT��0p��ˡ��~�$�"$��D$��A!��� �Zp�R%�N��;�al��f�-N�	�:���2��=[Oآ�Y2�]5�TWO����rA�A���*��#`���C�_J�vF�*�ey�.�t�"�H]����k���E�����ƽ�ӷQ�NY�װ���#[Tz{=@V�񾗢]r����џ{w���������a�����y-4Д�}zA��!3�"8F�e,/��m�s��jkz������qi���n� �7S�wCu<CO�ki:2�ҧ���:��g������ϝ��8zO�1-�fy���8��OJ�Tx��{
�A��m�����Cs^q�||��ts}���ph�r�Sb4�Dթ�ٳ�#]3�����?O�}���l���H5U�\^�6a��1�#F����$c�9`�Z� �Hܔ_���zK��ŝ�q2j"m	ʑb���}7�"2�තO�p)<^�`�.�%(aq೐P��d����ւ����ڒֲ�L�ea��E����!��H�i�K�􍈨~���g����!�opJc��J�,�����c�.;ݥY��b��Ww@�[�:���vx3�`s*a];S��'�ܮ�e���?G�b�Z���t3(q��e��e�Hi�4rz��o2A����;7k��	�H�:�Kzfg#9���Gp*'�\��k|��{��x�L����!#$d� ��N����\q*V[����{,�����,1m˅`��V����X�2~5���m�\ �o��5��s�	�\�*�T�<���{��r��-͐�>�`�'�n=kռo3V�ұc�=���D;���y�.=*�&��W;��"Se���7�4��k��O����{�r�U�sN.��wԁC ? �ʕ�O~u�~�dL	!�V�"�b�oW��≉d�%V���ˇx���|q'G.vtӈ�Xt�\���G@�q<�Ȏ%	dF}�dp��'��J���s9�_b�e,�WKKݺ}������st͛�6�M�p�������m37-�r�l|��z���؛�[����9wK�֮�k���c�#M]�����h�Ba�[7K��Ik����g��r~/'L�}�0{;+�b����q��/�T�Zf�O�\������ef��3�η;:�="X\q����/i��]4�}�����/+ k)~	Gt;4&�q�׹7i�!Oܺ�����?���f0��vNU��luH�^��ƾ�I��#&�us�2b��.�1�l�4���h��A2�N]�{����&��p�L��4������:�fc�,�3z��ڂ�KU�5m����9�F���Eb�2�vmj�3\�
�U!�{F-Oz��;{�͹�B�S���W7�eʝ2d�w�*I�$@FI$��HA=�7�� �4��ʆ��&g�DbFB��lW������|�Q��s���<&CM\�Ȫ3f����-\�=Ntϋ��h*�Ͼ�
J���*#�9_ҋX�cEr[�e�+z�����A���pW����H�9Ĉ�������PTҎ����A`9��4�]�6�[T�\һh6���B(4]��b�_��1:"K�<��������+J�)�W8
JF�^�2"cu�=6!P�����hEx�]��d�C��־
2c!oL��!k(��7Gwn�b�xځ.�h����a����j==�����(��J�A��7�m�Ly��G�<�xE��L_M�V@��H�I@:X��G�RE��e��5�45��4nz��M���[f��21�d	c\p9�*���Xk쨸]W ���Q�fLN���u�U-��n��bj���8�:��`mѱ�ŧ��ȥB��amAe�5��N��xG���H�,^v��O�c�dv^�ݽ�j�q����8���-;���t�)�*���$0��b���q���+��~�9)n��V.6��/�H��6mlרVd�1Хj�u�=/���8�]�B�P���Ǌ��3~;���a�m�k}�DFw��j�}G��C���;�5��W��X)�ժ��ۃ"��ML�Z��{SY���oy�s-����� �$D!�"IOο��vU(�%3��q����r� ����ꖠM]&Y�0a�E'���@ߠ͛��[��W����3�I�2�C�t,7	�F�4@�o`I{�0���)��E�/�U=в3Y�Q�������7s��4��\�6X!�ۯ���L
6�aTsҹ�!^%rK�j��Ժ�O=,�}�$5	�B�!���	�H3��T�:]B������}E巷�]�r�.9{Qnx�lru���$r�^45Z`���SO|t�8�W{s���J�35Y;�c��j���(����^�A/l�����OD�7D����(�/��'��<$*ܝ�F߳27l��g-�O��:F�s�StN>�a�w��xsh�Yr�����'�#�zv��n����H������[b`�M�b�$�F�+���]Ȟ��f���4�]e�pP.��(�olE8\�1��JP4t	�3R0�qQe��{�'�ȽQCvGpJ���F:���Zb�=�9�t6:�2� ��n�tM�1���e��Bc am\��F��kN���������VZ�JN�l���<\�n\�G{�>������̽���J����l)���z�g�9� }��Ō��a��QlCv�٤��dȻ�Vn�3t��]��l�^Ns�͗ȕ�V�*3�d�ٜ����v'Ξ8�������}�ţ�mԕ�j��9����w�� ?������"F ��$7��ϕDQ�c���D6�8�}s�J� ��A�\z�46b�:袠`�",&БsXI�v$��b���^�.a�c�B׼0�*eЯ+Q�[�l&�&�\Ĕ�gǠ��&��RЪ<�=i�z\!��0�b}Rt��%����2��k@u�B�v�ya�P}U�ӗH���c�Yw�Zt��[Jq%�"}�_p3��4�%���-;���3N��h@�.���%7UnU+�ۭ��B߱��]R�z��]^�����O�RUܻǢO\mģ}b�-�������c�E-��)[RՁ�LHpNLG�z��;�`C���X��:�*�v�<{T6֗�!�nS+n�K*���hm�_��TXϑ8lF�g�����{]S��SWB��Ve�NR˺�Q�=/c��8՛������Zh4%(�@^�}�L�؋��n8�dA�~��j`��!ѵ1<�^U<�5 t���Q���	%�;���<��yR؈(Y�Y�ޗ\����H0j���J2<��_nb[�(>3�&u��a�R��PKܽ��i7l��r����R�ۭ��V�Q,�zzv!c¡�ơ3q�&��U��]�g�lm=�`I\��l�S���DW��j�:�y�~��{[�����s�d��8z�T�B��hBX�*E�\p�׆�d��6p���q�~���{3g�!�$" �,�$"$����C�?3�����?N>!T�#�p�B�__Џ�3�Z���e~ʓOO�L�u�J��P$^�q[)��c4�_g�D⦣0͈�ZhTtr
G�>R!O�r�(����ݔ\�:���pγ�zo��g��Άh�y���<tE1j��g�]����g ����W��v�kݥI.<��C̫���j���r�%��'�H"���ڳ�J#��L����b��Ii���g7*N�.���z�[CZwp�1��\G_<��v�B
��Sj�IJ}z+7��7Cv�T�g����"22�Lǡ>nE���*f�fBtg�V0f�c~���X���jfgٖ��sT�t<C���v��X��z2<'�ҫZ�.�UEx�K�M{�eMV��{��󫮫��G\{ϑ�����U�V�U�K'�"X\� V�:#s7:	�3Y��)����|�٢��O7����Ц���U�ԊV�H��D݉�,�[�8���s�2�+�jk}�W�x�>�qY�&�m���st͛�#qT'���B[�U�(d!�ex䦏����F�vBKm�������.��D�v�VZ�p�M�:�b��΍-E�u|)���u0b��vS��i9���"{�U�[ǖb0(ی:�o yNkVwB�j�u��&U�}�Ӿ�ݿvOѐ��"0<�(� ��������>����x�6}�.�$,�'��$�]1K��E*�q{�r��yI�9�r`��(�_]�9�$w�B�p�`{$N���#r8�T7��ׅ��#<�z�l�
�����uv"�t�t����âh<7A],��>Ѿt*�d�SC�C.U7�z��l���]�M�s^�Q��2a#��dI#uxBf;�"u>�ws�Yﻷ߅I=����p�����*��B�}5��cu��VH
��z��_~��y�b�K�d���[4�a��W�uN�T����E�&����MG��3>֟gxY��2���<�(ݙ���sW�}�L�q�%�=mM�%mmɽ0�_W�4�AP	e�L���W5�nZ��HF�+�iE�#|�����s�@��_��boú�s��#B1%ډ�b�Lpt=h1���S�z-���=J�n�C]ԇ%�Bi�Lw=C�Zs�љ}B(wNa��p����h�B1���+UͿv5����z�%Hp$����d�VO���6�/`����o~�Jw��/�t/(���t�7��YZ(˸e������P���ǵ��.wʞ�֩�X�`%P��J/�]�-������}wNF��V�o�4�r�4>��Kl�]�ɝ{b�V��e�<�l��.Q��ΣGc��n�ss�;��� �AAH�[�� ��k6�9M��C}�d�M�6�֙J�!�j~�v��7,��ȫg���e�5�m=Fޕ66����p��@��s��UѶ���B��Ja��
9�����ޱ
}錉��*�$���zd�##�p�r��V;��]}B���"��t+��ȁ*a�GdtDn����Fmɖs/�������2Hcr�u2�?�D�ڐh(�$��#�a=8К���t��Q8���}�/��AQ�6�o�As�(�i��;�Re�`&JǛ�Rz�D����5��ײ�9�Һ�t����¼�;��A�v��&�_@�=�a����E�u'p;�˓A�Jlv��i�U�����Mj������Az�S;#s�W_z�]��m{�н0�jj��&�m#o-yV'u�*-�
���P���!b �Q	�H��U	RG�a#^_^]T{��]���*���;�.��u�U��.l;�<����H(�<|wP8bkk���&�nיݰ]�S[�ĝpOB�䠗���9�3?t��j�Ƿs>�Ƌ&�:���U�ٔ��hr�B�q�^�p�b��?	<9|Ww"�����β,芏����Az�&����=�C~��뙀9̉!�}7�N쮧;Z�k�V��i�����)׏����L�+LJ��\vN�	̑�קhW;�R�E���KN��ֵn����&���\�h���$B"H�!���������>�ǘM��?����B�)�=r2�Hf��P7����$��yl�u�K�b};�9�=�q�S�zov��-�*�����Q� �����-��D�L�xM��;�r�L3x@�'��1�����-7!HEW@�juJP8t��g1.��Q
M����,˦.�_���G�֬�W�/av�!:�4�L�Mc^)Ẇ@%1�&X����}*�Q�3�>�ڨ����T�niٗ�V��A�[��9܆+��_��/���p�`�`�C	�+=�i���a
�w����C�N���L9��d-{aT]EI��"���2UBy�E:��6:�0vG������%C�}#^w�+��a#�	M�	��O���Tr� z/�1�CJy�ٹ�]�P_�Քtj�Bd+�&��?p9؃�0��|�tKN�s�3݇�-��C�����b�"��"���e��er�Jҏ� ,�|B��p��#s���-��cB�C(�RSYOE}=ƭ<آ뛦E-��+�w0�}���A6�!�d���2�W�1�\��yW��ܭ��b�i�(��ˀ�s4W1aɼN"Z�r�Φz�
�!�,5�)k�x.\=C����}��;�I$j���T�$�"�'��,��^�H��s��B�n��e������`��
�ȁ��+��E�J7Z�8Y��u����_}���� D"0B"A� �����y�+zVꩴa����/�J.�7E2�F�Q�� ���p��w�.� �T�K���k��:s��!���;Zak^6hV�[FH��q�O�`7{�9-?hhI���">��7�
d8'`�n���K[*�Z�<S��L9�H��uО/:��O i�ʐ[���U����5z7:�	���#c� F˪���[T)���aC�J�=��'��Q� `����`<�3є�����Ʋm�d'?9����B���f�y�:+�dJ��^5>	�љSS�g�דC���^�u�����.�f�z���	��1����U(�����>��P����麎�ފ�m���n�KH�����E75���r&!,,h|.&%M�<��a�<��U_QH�����l��`����D<M;zA}����,l�<!^mJ7��j��`�.��mOg�_@�2������u!ɇ`�{����`5��e<3��lU�{�����9�e[:"�ZG����U>�zq��RR�va5�T���� �=��x�7MeNhM�ܚ�ۃ:���l��<�7ʦ�Næm�캺�ѩ��#0�+�挧V����_ZɌh���[g�a�
�[_5��(���'�`�e�e���r���J��+2ȿ����4�,;g����3xM���0�4o0��)�Ǫ��[)�>��%��޴��w!�9���|�.�*u\�QCέ�4�ֲ�E'�����+�q=䳍�&�y�' ��ph ¬?e+ݭ�5�S͆����2��|褉�m6
��c�u�J�K�/EGxՂ����v9�f�T�d�Ч�*e�s~���࣎��F%��7!Sxc8[�5���ȯ�l��mX`Et�����%�J�Ҙ�{��du�f�6�J�H��s32R�e��F"OL��::�N��T��1�{��N�TL+{�pGy*�ʀJ�ԢM>TBƛ��Xc3j���X�Be3��i�i�40P$B�����vbA�r4��{�j�h�h�"����PZZ�H�N!�wznr�&��}��'��1�=(���63���c��1���(\n �v���G���5�um)���X�۳����T��E)�]��`�=|/~�Oe\���I3E"���ϧ+�ĸ�I��Ev�d�lM�2�SN����3Tt^�9��}�e?��~bz��^u��:3�kh)�=�hҵ{ugF�voPN�-��V�[G7��V��4^lW��gn�:��|�����T%�|���K~uƾc^�.�v�ޕ۸�����:w��U邤���N�x9vr��KЍ'�L� ��P�ɮE����T4��ь�b.��]��q2���p�[�y���j;vn��Ԗ�N��E�g=�H�e.Wͥ��i��.e�_=������}[���d�2����I�7�NiZ�b��!�I�{ �[u5v}��W]`�G�GF�=�|�Ү���v�t����R�Cv�".p��M5�������Y��8;�D��'���g4�2Y�*.Ǻjd��Ga��N+�Iھ����vcd�gA�T�0(�6�j�ђ�wq�������X�-\ǋ�6f'�B�N�¢ SX��d�����rs&���!�v=v�&̡M��wփ�,.)GpC�����]#(�u������YwZh!o�Ďt�u#�x�igf$o��%D34��o_�P��+���gK,Ž]�8�,���.;����C�]�ц�޻�`==K���\ɖw� ���Gع�j��*��T.�'J��}���
6��#���6�k�cpD�Ey���ʺ�����"�[��+�K�Q���{	T�K5��k�MF�>�UglR�w�u�0�muu6��6՞oC�ʼ�>�]����F��,G.ul�;��ŝ�KT�:�*/:���;X��{Z�'�ҐÔ��ޞ��m�l�V%�m��Ɣ~ʮS�kH�UFگ�S"��������Y��ڣ�j�m˃����a�\���
j�Q�X��-��M>6r<����hֻM:c�-H�(y����iVՌ�+H5�V�>8l��ݨĴ�D��VFۼ+2=q먢0��E��&&1��Z��,X�1gM�>8p�1��ԕ-h�w�U�h���VV�YR[jҊ��U$��ֻ¸ռs6ҟ>8l���n�ԪV���Q�"�j-2���̭��E�M9X�T�Ə�8|�W�*��c/)MUnZdDVզ%��0�F��F����Q��G����>|H9�K�SR��q��qeJ,fF�)TYl�US(f"4�aEQ1�S��8pQ��ŰA6��j��1YZ����)z��Q*	T�E���,�QTX �JZ-U)V*%J6��2�J�)��O���a���P���Dz�)׼��������s�E��,^GƐ[�Es���]��7p���)��g>���'����=���b0�Ȉ$"! �/9�k�߿�~�{��5!E�A�-(���yX���8�;��W��G,��K�5��c��/�A�|_q���9HؼLXȼQJ��XN/���L3EzdA]#�޻g�9q��;����ʵ��Q�͚nN�ĳs�'��YcU��JĎ�G"~��d4����|���"���e0{�(t2ڵ�.9nE������bv�N�\.���ûxO�Ƌ���%Y����sE#$"��_и���!�ۓ�L
��O�a1V�"�E�5]����L����{�n�[�(X_5�4�L`�H�U���-qmh�Mk�i����5~����{}5�Z��x��0D^�8rӐ�j
�[B���:d�S]�r�O�wr�ɘ�;x��}7c��jӬN�$#��3R�deN���!<S�&w�L��{0$���7��<�Ԯ�����Mm��n��F�@C3��ER�h
�Fꤾ'	4//j���B<�*��#G>�Q�Ì�Z#0�8Z��/��:'X0T)�Z������i��Yh�u�v��lPЁ_p�vy>1�����BU��u���<�4�����⣁`�D?�;���I-k�QV/l�"�r��V��O0IfIT�6��RȡI��s]�	Mӷ�}v(V�$��:��;x
z��i�N���7yf *��h�n�W
8wq�r�+��̫���WV2"DQ������fg���~~���9�^͙�l���}�����B��Zhr�\k�����(+&��++ׂ�{=99���HpQt=G�i(x���A��v�K�v�,Ť�I�]��5���`��]���}�(��g}�Z)�H��A�.��mT*6�X��Wӻ��]���A��[�Y����E�f�Wܦ�:�p4"~b,��l������Uɶ�� Bn5�i�s����j�;�)Hmo/^\��L�٬�td�B�V1��R!]�""��u�f���L�uXyݾC�U�,����^A:�_����m!�1P�� �Ár,D��9�/�L�d1�S�������q��T��^+�][���qk��ȀT��f.��;�o,m9��םPtGv�!Nb��0X[��-6�.Յ�-;o��v%�h]�8A��򟮺��O����oi�<�?D�f�(�dO�aۃvfȞ�P,Ze�c2�dW=�U����^T9�Ӣr#��:�Wj��zD�#Da�M����U�^nw�w*x�Hc]ϽEw�K'�f��=PN�0�`��`@�r�Ơn�]Գ��4έְv��!l�W��Ga�o�F�yӷ,w��ƶ��>�*�A��}R��}�� cZ�غY5�݌�\��ѽ����ݎ�-�:D^�Q,����GL��np93��]h��V��v7h(�.�(f�sEs_�?���F"DQC{ֱ�76a�y�"8Z���[�����{���{�2����)���T�{�ȒV����N��p=]U�[���E�����7��@n8�=�$5	�rc ��ڈ���jaOw�ݺ�X��y=��F��['\Y*K
[�t]x�����g�N A�O�&�a��Uv�AW�W)��k=�:"V�9�!��t���(�;�Ss߼���_�o�Gs_�۹eʍS�ѦG{!�/�#O�{�a�@˭#����~<�x���F8#�^�?���B�W��B���v��� ���^	� /[��7�'�fC6nt�LIz6�+#�����"��V��'ڟۓ"{�(�B�~�T� �@����d)V_{ޢDQg<�Do^j۽������(����K�����
��(�hdPc�L�"�	��ׯ{�{��l�qRluW��O�XH�@g2Yә����/��z\�5曏Rf��\)\)A���R3����ڛ%��p�П\([4��J�ʖ��*C�V3���<і˞�=a�*��W]�Y�ߠ;�+J1R���<ّᣍ�8�}tu�&J��ܼ��.����l�sǼ���-u0w1���Y��v]��F-j/I��<����RX���{�_*���&�w1�98j�:�g-����*b�VT��)��0`�M���5����(��""�{����]�;�������~%	����0F��a)��	���'�*9b�B�g� ����p�6�2�r�^�v����ř�P�i�`y���9�u�A�wD�!���u���V,v�.�Ƹ�)7���H�i}�>*a�}��B(}��o�sڪ��;�[��\�*8z�]c�X�ĝj�رi��2)�TG/|<���MȈd?(:Z)�վ�ۄXY�����br2���7n]���Qu�>���ָ��RDɿ�	=զ��[Y��#7o_z�+lS�$,��ʇ�l�����9buIw�'ݮ`*b��J����Ӗf�u�LZ�`�,���f9�7{�m�ð>Y:\�#uo� i+m(��f^M_z���A9p!���.~��!ڱ���{��b˾��"���z��w+���9bI5�Adj����cJ-����àG�~)�͈D�{6]��C]{E�]�'�����h�r�g�u�P�m=r�m!���+�"$p��ax�*�YG:�-��[���#�PJ2D�d�H+�ޝ*�c�[���F�uq�f�'�u�~shh�O>�4����gO�w��K���`UqN���M�vӥN�X�(����f���)Bm;�wE�z�&�&k�+K$��dv ݋,�{G|��o�]�5�:��$H��0�U����}�����������y�;+z+�(w	���:�;@ׇx��4��g�����unŦ�s���>>u��9n=�t�`�#�	HpwÉ�xmC��Q��/���z��P���iý�:��,��v���/V�ov�2����;��4
�R2a��ŧ�w>��/9O=�3�TJJ��0ɞŵ�*��ϸ�ڒ��/Y�����&��!�mο�Z�����f&��My�ٲ)(��O��L�sd{��ȯH\�J��Yb���=#dR�Yuco�2�E�D��"�b�U����.�(��"Xd��x<�[!=�WSpz.�U9;�W��y�Y>Fq^��=�f��r%}�������j���g��5=h�/	������Wnv���*�z���-�tKNۑE�7�l�QP0nEê��v�ޕ6�'��ؠ$�d"�O�ax�\�:G�v�7k��y3�z�TXsP&,����v"}��QW]����zc�p!�^r ��3��w$Iz�`�ָ��z-�!�P4��9}�#��%k������n���0[�o��o8��S3
���w��gK�3k&�.y�W IK��a=��Li�&�vlb�im>��X\�u�}�N�T�*�%��`�k�y��nN�\/H9����i;����(k��]�}�ҿ�uWVA��?~?���}���.4b�|��a�<x2�j�����k���N��:@vK��K(CY��`�-f��\1��^�������$ r���edI	�NB޺�>��܋6�P]���֕F�M���7��sܩ�:7�/Z�֦��?@��Ix�(p^"�R!ؼ#CW����+�3U���(*o9��X^9��1�����U�3� ��H��66����j"g^��ݷj�Ӑ��GJ6wɉG�=�#��}<��5�Dw;=��V�����Ɓ ��\R;�z�����$*9kЇ����U�W�w08><*.�����aǗi_y�yE��ӵeb�}�1�	�3=zkNln�H�3�BkúIv�w��ޔ<�e�
�+��s��9��0Ӝ��M�u������"Ȁ�,��X
�+�~ݛk���!C�D����E_/� ��p,���X?P���$��F�>C�����	�?B�TGS]��-]t���a��m�0��a�A�	�Fq��tm�?\�B��	a�k1�M���"���krܡ��WQX���o��Z�q����}���� X�u��0��La�r�2��V��H��-�ޏ����e͐��;�81��WE�c�C��r�Ԇм�I{�[�W����Q����.�.��A��{W������&&�\�������#@F0D�$�^�v�栟:��f'��Nh�z�lC	��L�}Hh[����-w�E���  k�7?�bC�y���_�M;O�$p�vInj�%3勢Zw�ޠ�C������3,�&�͚�7�Z�XQm^q�C�G9A÷��(�2=�"F�e�=���nܮh��<��-h`�<��PQ�v��V��� p�a��6���@�o`I]�a�q�E�57/d���LU�����#[_Zg����j�a���_lբA򰂢���_+���ݻ~=/'ג'�j��1����us
�����$�?6��PD��!�X�=�|Bgޜ�*���Ě���ۜ�LJ�Y_:��z{���\E��.{�u�'���CU �@���zvET�Yѓ���di�0��65�����hW�T-Y��� ��]�|����X�l�t��~����ߟ��`�<�V1�C|N������^\�݉H䟦�������ᠸ5���>XN�{�^���f����.,��	@h�
>!�De���y��Ng��렌�ˬ?ߘݧ%*�QX��nwoɹB�Z)��'�f����,;�:�Qs�v.-�u�z���i�:�i>�Br���?�s�J\�54�R�-���%�v�bg��\�'Y��F�y w]�gR-"9,Ϗf�z�}Ǟ�s�߹�����`"�E0`���ٳ�}inR��y�^���4;D]�v6�w��K4/>R��QQ����gy�"����z���4Č*w$n�C\B��F�xE�*���t	��_!�����;����%�L%�U�wh����Z����?fF�Pj�;��U�B���4���W��Td��𧄏�h�D�N���y��#��փ���WU	��T�>��o���un�KC�� �g��Zv�.�U����s7+so��qE@��}ca��9ao~�T�;�%������)��߯Vd�ܚSz�<ы��Ÿ�U�V��k
84TY�BM�B����#�O5�%4�Ψ��.��N���}9�ݚ�zCvKԥ*b=7������)ZP$!Ԇ�u0S�с�|�=o1��^�edu於���E����Im[آ���� �@�M�į��:�C!�yW�L;���\l�#�gr����m噃�#aV�SL���R����::֚H"h��f''�b����skAӢ0C�BeztH�5ڨVX�S�;l�oE���ņ�'��M	,N�D`c�ƍ�x�ˑ�v�V�A��w{e{`�\�b�!k�������p.��^ܐ"U�g`t�&Qv��tĻ.\C<��Z��j	�>J�݃���;:;�ۥ��w<��i���q������.S7!���c�\�S�K.>�pH)34h�ϓrƀ���W��"P@�?�H��dCo�c��\�'�K׮��u�?oh�rI�si��Y"�q�K�eW�T;�F<�B{w��ߵ�Dbb��K���ƃ G� ������$㯽T(�;XF����s.FO�"jb(T���nwkҮ�cj�eE��?z����<:D�2�+��o[��N���d�Fb�+\�^��ӗ�?���\{� S�(��T���O ���avJ�y�[g��ѹ��9h�g�"��H��]�F���z>�;����w�+�cpB:RS��#ooX�)��X<�0ɰ�\ "n{^��15�A�}�X��{��	.���/���n���Q�[Ggd��l�����t�U���h���O��g��g����=��	U!ɇ:���3�s�:�N�ڃ#��a3���
�N5�T�'UdZR<�3D�t0{�;�a��.a��v����u����(m��7�׳�a��*E%`�5a>SJqdwzr+�;C$����ϧGQǞ����KUϧ�U�#دr�KB�b$���ځ00͍�.K!���J��*���%����V���ZJ�Z������p��r<��@l{]�&ǔ���)�������'�Ĳ��c2��1����/��h���3��:���Y)I�ջ�Oڗio��[s��+�.�=��[�N�oG�]k�3[�|�s~���#Fy�`���a�z�S��7����C����<çB�8�Xk��ʍ��"�w�Mk1�^�w��)�i��cn;�~�#e�ծ�km�]st͛�@�]�X������.��/h�z�:{x�����H�>�͒f�p� zga	ݧM���6��#A���+�g�6����S[(G�r!6И��#s �E�v��>��mo*k�p=ũ�e���������M0%��y�[�
5��q"�U}�٣��t+!�M[�JxU`6�#t�����F�U�c.S�tr}w���"y�6y�{���`G=DUK۳	�4]f5^���[r;Ya�ƙ��[�֦\}�uL��E�LaH�x�ڮ�EoT9��L�l��޴����}l�����Xs�s:�\��O3� ��rW��#��%O��>��EP^�u]��͠�t"˔D-8�J<�G�d�����g�X;�b�NZ�/oP� Mio�����@����&&^.�0-��n�my�hW��/@ň�x {��Ӡ�\H�C���;��Rܥ����H���@GM_A�$	QW]�Ί�ed`���PE�`�<*�
����Cvn
��^Z���c����0�����7e����\-d�9�ɩw�n"7���O��6����K.pP󳪅��n`�����nd�v&8�.����&�
��؈��(��DR�|�� ۺ��'�����	���X�)�B%�������n�kiuՌ[ݨ�Iݷtr�L�h=�j_[��\���sP��ٶEN���
��u��rj���81[ �(-�[�4�NS�sGh���>-��r�8+7�ږq]��
/"�%Y��m������ҁ[D��)W�*7�X]�����������VG��흕��I��/0�Xc�����Vk�im�y˶�a�q�7'ҝ�_:�3(���U��3�I�9[Gy�f\|�n��>�;��4]�e�� A����Jv�jW)3��F�,��������}\�0�IQr.�FŔf�IW�1 ���חD<+ӷĒ�ho�7(�У�ڻ���T���5ܻ��Pxe�np�_�+�{��Q���˭=�R��a�s\��n���S���\�k@�(�Kf�aL�w{Ye=;������N�u���Nb�X����Í�jgb=6E��N/su�d���HvYt�۠N2���m�I�t�\�i�������u���AgVkf�T!&/$�o�{pG4+4��2�/�9j��
�]}6��Z3n�q�s���CzA������T|"���0�Gù�X8�W���Kg(S�d��5����)r���pt<��gi5ǂ����Y�C���S��g]V����.�i����G����6;�mB�{bE��R���D�tW-�u��}��Cz���+[�x �R�n�=�x��O���ؠ#V����_k�����u�&�C�-3�G��CE���:��5u{�>w��r�	D���An��հ[u{�i��9��CL��Z�q}�>?D�떶�=���������&�����Fw��૮�3��W-��b.;��G�;qJ#�t���ۡs
�U�)-j�Q�5q��կ74� S���-�}11Y�؄$���F͎dņ�5t��"Rw+4��o<╜��9�۱5�7���9�'[�Y��y쫱wIt�
�m����]�Rfͬyi_O����`˹���GN�yrw�r޼�k��<:��h*����[�`\�����\k�N<�&����6�o)��
x�Q�����8�=�s��]�WP�E�5m��į�ˏa���U�R���Mm��{�Y�qN{��[ɿ�T�U�A���tx����cP�bu�[�s^o#�^M8��ù9z�8��\X�k]�4b�WQV��M4�X���%�N�0�m"���O%7F���e;�@-*��- �4)�E
%ҧ�ˢq'u�[�I���р�% ���2��j���)imJ4h�%DP��h�T[Q�)������?�?������i��2�h�`2ҥJ�T6er�R�5L��Z"��ҵ�b�T�VԫZaӧ�9e��Q0[Z��hV%B�b���Z�fU��Xѵj4�т������5�0O8p�+Ĭ��$��UD��ZR��J�������b�Z��s-�eS8l�(���̸9���iQ��ej�R�eb-b��mDF��.�U�r�Z��>>8p�^[Zܦ2��юZ �[
s.-E�2�Lr�WGWr���Vڥ����8f��jT5�1�B�%�1TffT�mkD�R¶UT����U�3
��ԥM�8rq**��mˎ6Օ��m�����V��IK�0G*�%¥�MQȖ[W���ѣ��8+��E�k)JҢ[Uy�u�նҪ8���:h���*,�J�Ʀ1b�+kZ7�Z���#cD5��Z(����b��QQ-��1�[J1�LT1AB����!���9r;ٛ�;�֮af�{X�wZ@�+0hn��nw�Z;���͉Q�yv9��E�5�r�޾��a}��ZwUm
	Yqӭc��т(����d�?��q�ɑt��C�b3VS�H���4J7O={Y���X����d�^�$D����y�T�ߣ?�����_���j�_D��VX="��V2����Uϩf^��{ꖅ5��C����L�d/#4!B�849ܰy�HJ�4]�14�Uc�@��q��a^;�{��8�/���J�{`�2db�9m��|n�A=,�%����t�� ��b��u�&�Ƹ[#�j{�FdR��Ÿ�CȜ�ף�ёکlp/��eվ�N�1l�6��q-�N����u+y=�=�R�ֺ��G��::EБ� {$h܆t�l2��s�XH�\m�r�s47a�zyqcr�P��l�;"�n��p�Ű�_`.~��B�`{6D��4�O)j�(of���Ȝz*�T���[��)lV�	]�"s @c�a�!6�����Q��Tؕ�̎�8��}~��h��+��,gT�W����j��>0=�ޚ�I�	T��B�^)�]х������~6jZ��aT�L9���nR{	AcK���≥��F�:�� �IL�5�/��4��E�����r��O�tIm[�M�J�lX9J5Л)�d�u�����"6:�;*�f�IKj.זV
���Hp���9!��ls�R�N^6�]*�t�Ջ�*�����W��6{��)4�9'��R|��vT� ]ٕy�<��o�?��"�"���#7��f:J@�९�� [z�k�J��vN���*�
��̦º�����N��^]u�9���3�x��̳���7W�u�=_ܔ���Q�B��+z�4"x�����0*<�1ZM�Ep��_p�i��D������T��k�%ь�D\�|����(���Ƿ�#->�����UO� ���<!��~������-�̊	f�+7��5�U��33ѝd��,`�{��P�u�C�̇�m���cD�y�>@����S�ɮ�]J��藽�|���ދT׫˩�@�l�0=�˃�4�2�|*��J��:��w�gz��Ĝ���OFBH�.��ړ���dv��>Z9܆(>���z�5��\,Tv��5r�����r"ȏ�/yh5��M��T	���ڎ0fV^G�4�$Z��6�ȋ	�k��Ue��ٞ�����\��1P��Y��`�i�9�>�d�N԰�;���~&Bd��^�8j'F#q���u�?|����4|v��a|AC/HV.1m>N%��5O�m��{���gz��+7i��$�\�g;�m���ٹsN��[5����ݖ����з���۔R9zʘ.0���t�*��% �����c=�}��S�}���+��ݛK9b̮P�c���/_��]�E_git��wD�Z�B1ɯ���y�{���2���G��
�߂�'�C����9�w��^VS�4�)Y����[����C�s��қ�`C�+�	�I�1�d���T�5]+�q:x�}J�Y�3�|���Xf�7}N'+��xd9��H݊�ȿ�T�O�E}��A<��$��} �`cD�fM���z_�. �������shS��8Tg����dϡ^-/�2���Ӯ��d������dp�<��D"9���2 �k��:F��.��Q�����M�I}���p1�C24źMz�fi	���6@x"5�O�4�A~[sq�ڡE�t݄/;`;�m���N�LVu��q͞T�>��/j�A�����^�� ����D�3BC�Yj�u�7�������<�}A�̭�r����L���:�F@���P\iO|����@���l\K���h�+�'璁G'�=�l����ߵO�7�(顾&���Nu�z�#s[�H���H>��J�����N��c�j���px���"��QCe��YHS��G�����}O����d/��{\w���J����k�׵`��}�˱ֈ3�9Ef�����H��J�q�Lǔ�Q�JΨ�G�3��nǼn��oխ�^���Ǭ��-��x�a��jw���k8I/{&�zs���/���
> � �	��vto�]�Q�.$��<-qR��*�Wo����h�_I`k�]6�l@��ƙ�fut�=)	�V��Sj⒬.0k��
��31���zmԕ3��-#"D��2r�cV�:�^��|��M��}ϲ����U�+)�Ȥ��lpM�k�ȩ�p,hlb��^��iw{�f��w�'�-�`�O"Z�ϧ�v���W�1P�Ja��"H���-rO���u!��#j1Wy����]�%��D�Ν
kiY���k�뽢�-P��{G���A�ώp����ܗ���e�y�����Qt9��6#rEz����cd���7ћ��6��/R������X��ܢ���B~ݧM����6�uN���P�IٟC���,N9#�r�Llz~S���E	�b!7���;$Iz�a��	r�j'������{I��Wx`ic;L�Wzh�CdF�����aƔxj�����4݌Kŉ���6Mj4^�t�W!��}�k���T�J�ļJ��� �c�6A	������}�o�/sMY*���R걌j��N�T�7=c|;�.a逛B
�^���d����FWSN�[���R�5rV����!����-�Ty��y�4��Mc�e!���l�ۣ!�ϴZ亞�Y�G��n�`䧇w��KU�t�M�!yV�n�y�:�������6�:��U���|(}@P�G�����i$��~�}Nz�ݍ�m
���V}n~��2=Cb�'	G��nV�Un%o�<����aF��nKԾ���u%���k-{'��+��W����Dkg/U��پ_���������� W�a�0�}�t�^���]���c��&�?�k�W3�c��͸���>�y�܈����(qEp{gk� ȗ�V�s2U���#�
&'�a�d�xc)ѼӞ�ǤR�徴��O� ���-��e9��%�0����L6�k�ޟ��̈H��sQ9��Ӳ�;��#A��_J<|i��6�O(��b� Wo�V�]6�Z�`�W�7f-jn�!��q+Ԅ����Z��t��ñ�n���N���Z���iX��"������nB�`��&o���e���Lc�;���CRdᅉ1�#!�Y��&quy��zV�zM<�L�����j]�� �ܪ�+NV��4�4������$#n������	a �9DKy�����)[�9�� p'�ٶq����dbm+�j�l�]a.�I��dÕ��긞���5��nx��5��me����~�Pr꾻��8n�W�M��A����,�]������Q�Uj��R��ksH�]k��Ց�L6��66SC���o>��^�E#1��n����x
g�R7-����$����m���������5|Ϳq�9"��p���S�&p3�L�Ng1�b!�.�$n�d�n�OZ'�Q�襜�w^D��)LL.:�_�"�6��Kv���k�n���,���^�h�m
�� ��5�UR��"�$�q�x�!���^"�y���V�����!�|�vn�.��-㝕C�r�]����oY�/U]m�=۳|/�^`��p��~Ńpң$��'�Tɾ�~��w�ҭFLĄQD\}3�=�G��88V�����P�H�͠��6Z53�tr��l����=y i��j�^6���[��e�6�Kn�.x��jΗ��Uiq�$���#�Oi����1�p��]mMol��:%��~������=:EW��#��pr0Cq-EH��q �] o���)�~�;Fʍ�~�^G��>�}���#�'�u9���~�/�����ғ����m���{��hw9�a­퍺>_�t�ۭ{� �ee|��b��<���W�qX��cm�5n��|��{���;wb�#���y��w�v��O��u�іEu��_�����p�"�Xn�E�Ȝ����3�|zG*"O{�M�!Q��׌r�u�.��/��ƶ�ms��3������Tۭ\W�{�
��k����������.�ʺ�ĭ��H���P��թtdz1QQa��թ������.T���&`j�Tәl���pc�0r��x�K��cgT]�-���5؍�rk��U*��٬ʠ�}V��#��5���["�W;�ݝuL��冠wJK�]@-�>� �o����`f�O���/>�B���'8{��vP�M�<��I��ä��݁&S^p��O��;+3ql��5����E!���4�I��];�(sX	p���.naNky�½xy�|��+����9=��l߸��y�)�_w��iP��|x����Z��.�C{V����s�o���
ia�l��t�L}oz��M.ޙ�+|�����~5��x��ݧF4վCG���[�w�j �:s��/�`[X�w7�ZܷS��v ��������&TI�̚v�\pN���	ms�����9���!�f�V�����s�G�x4���Nr�62����ǒ&aI�<�	����!�������su��On�`��N�)Xzc[YB�y���kIS�8��#�!�=�ϡ���Q_��J�����o;�]�����.Zl����Op���������*u�t�M��i��'z�@��b�<u��-)�`�q0�gwb�X% ����Y� z�e�Ey糔Zr�^�Bp�,�si� \^UW�.�t��L���U�n@�?k	��z��Ồ����:c��������uM���8l�X���e�3��Yx�T
8ӛ4�(�}&�]X}
�Vx8�:��bu3��l�쨸Ш�(���&��G�.%���(0�]�m�wB#S�fqW�~J��T���X V��J�R�I�;W>�n�ө1]�q�E=���MU����g�}J��p�;H��X �j�J�W(�B\�����d�9�g6�O���ld�^jе�Op�3ZZ�Qk��C�苗�mC��y�U����b�w��yF�u���^ͼ��{s��|���FR�oP�k���ʃF���v�zr�vbfZ[�u���gR����H�5Gp�U��WDNN�'/@�w�ն�\�!�\z�f48�H�#٪��u�oJ�In��kh����"߰���dY{nB�$�b=�tR�#���U���صչMF�;�i����Sn�ԍ|��]�9����v#y�n�n�;k�]ȹ�j�����Y�3׀�H�IM%�:�c�.�2M�c=��Et�
�ݣ�.��7��%uФ����K�-�$�59"v�D;0�7�Дi����6�N�X{dR@P�Çu�ہ�iP�����{���1ޜ!g�Q����wo�_�W�3�9��d��ؗ�D��|�ih1Z���v��َ���F�M\����G �A��n���.�������R`�ٝ;�[	�V9H'��=T�C: `����U���9n��T�`���������� �E�h+mWh��^���*�Q��1���♎����\L��4�mt9{)���/�����LP�˘k�w��z��L��|��b��+J7������UR� �mb�J�=�Y��[|]m�ЋXm��gV�ve�7�� Moj)^�imp)�]���7��
_]n�}�K����J�J���H��ý�V%�C�B��R�/�GU�AT�\2�V�u�t��m3br��:����P*ٚF[m�
�u�2*t���A��T
;��̇��:$��_T��UWq{�����B�nê��m����tJ3G��Ĝ�<ݱ�oOۥ�.+W�f�&<p]
ȆHX��6w�?�����~�T��9w���9p�	���f��j�-HӁ�n��L��rAnmz�mTw�h���6տ�m����Ӈ�3�y��I7J��!�{]=�c�F@M��gs6�a����thđȒtx��}��p�Ҹ޺S����N��4�2�p޷��}�����)��ٍ=j;;�DѤ���w�O�1�<���Kn�j6#��4����y�5脧�� �eWr�k�B�ɐ�B�
�U9u�w�"�"��6�����R7*C�'�@��:m�wd�N`��aYxꅯ%���Ui1B�n��KV��\i`��w.t.��:����y.�k]q��ޞoEu ���x`@�� ��w ��w�»�F�scF�S�d/�k�8-a+�\n�Z�+�\٭"��z0ݺ�ސ&�a���ȡ�a���wH�$���f�^�κ	��u���9%�ú鋏o�.��dnb7 ®�g�'G��h5�]��L�4v�\ݢ���t/`T�0�u��&��!��f.:�%C��H�1r���qf�E�s*j7�ȸ����k���5�a����B����$�u�wC�=���Ys�u£���k]�X$̒�=/)�|!2%���L�B�,��ܦ��c2���<JyoV����_}���u�b�/�]n��� 1�XSu�$%��&��lƘ�ʋ�<+Lف�՝m�'Y���j�{qn��"����2r��h�G1�bzc���X��U����Ф(�[���Q�M��WV��rN�ns)�<�龫��e�O���VW,r���*L�m7�=6�v����rJ֡fk��w���SAI*���r��H.J��o-��h�g¯�t�w�Xz�#��:E�7ڷEA�/�^�VT�K3�ۨ�f�Ъ�V2i�|��̺<_:}��ܮ��ݧ��>�� �*�;�]ٍ�/�q��I7`fN�g]�m��N��AI����`JyC��;,"���:=o�o�J����{�¸�:zX���|[��(=����[\����qjs���}mW7MMວ �
+�bV�x��t�M�{{�<���K&���Ӄ�0<	�'.�+�o�Rɕ�F��<�mܙ��*��_ۻ��4�M���Q����m���i�8���c7:U�%-[}I��A�j�� �Mv�XWj��8i�����N��s�|��xN�ٞT��v��s�1�J�c�����ȧJ�
�F��ע��<Ď;��&E"�a	��U7[�5���ƶX��M�B P��c�}�6��:���b޺5|zP�
��p �w��+Hn�!6����� @�Y�f����Ԛ�lp	��W�紶q�໫r�3v*M}(�ĳ2����]eR!]5��V*�ieYy�S*�(:��/����b���8�m+�̮1�o;LӮ��$�}�헂�cm�'CB�}{���l�}�"�b�����
\�_J�*���\�M�j�«|R��C�Bb�4�w�������|�fY�lS#�������p�+�����%L���hZ�M��z=`�,��tN�
@��0c���B���O_;�P����a��le�{�G.�����
��NKS�\�pÓR�qk�����d�۽]2ٮ���qܮ��sq��9���!�2����뼝�b,R&\ʢ�2Ӹ\bc�ED��p*`�C��&�����˘U��*n�h�:l���(�+y��n�C�ڍUE�\�r�U�c��3���R��-��q'[&��PQ���L<l�Â����F&.w4"e.��������F�UL�⢵O˂
v���Jff6�a���gqj�L����.��.WXfR�̢!��]&�}�4�y����˼�M2��#iQ�N#��.i�k�e0���Â�T�ĮZ/KMw5�PX�e�-�������V��ж͵ƉF��6�)�]4.�:l��m��!d�PU�>F����R�Uwi���R�˘�fdR�F���1$f���:l�Ƞ�r�>�M?9s3{�1*"��mf�(�V�+����n�U���\�B�u���ǎ9���iG4[�nfbօe��T�a�S*���ESV�hѪ֣��J�SG8pU��
���֍m~q�M����.F�(��
��]_�Qb���ĵ�[V�����(�o22֥թ�2����k�r�Qt���[j�W-)iLK:s��{�>��n��aO����(�����h�nٵ�l=x�S=W�����!�=�LL�6��_>�Fѷ S�˯}_U��ζ��w��+c����n�h�Cy��	S��B��ymA8}�ɪ��� eu��'&3G;�p�c�.���>_lF�,7d+U�F�@� ݆hzQ0t �Pލ���u��i�\��������=������jy�tn���h���D�<KA�Q�/̺'�MS�f�Q}S�g3v<($���s�@�u�h��̼�3�<��TD��)~�y�5Y��4�q<c嚊xޖ�X.�Ǟ�MLО�3.�V^�ˑS�b��v���23.��D���dӮ���8�JL��U�WA�g���ۈ]M;y�;<&ȼ\�Zd���'(�p�j��5r��A��Y7!��5�d�ms�E=�<��_j�X��>b�Au`牔�%-�[�B��i�]"�/�C�.Tq�hG3���f1�m����Gt���%^['�<�3��u�GW�~�\�|s��cJ�p�	@�
��۾�sS.�V:��U!�\�^>�]J�9*>j��m����%Ɣ�����
Egw9w&���*=���G|mh��z�� ��p�et}�ڳ����3�("e �j�X�	K�I�����I�5\oE�!���;�<u�tr_v9$�#�:
���\6�!�rg������S���n$F����,X�x6�����7u�Pa�I=u����� JȀ/31��T���
�C��b�'��|�����!�U&|�����Y�y�^��n�V����7��N�S�Q�H,�&nگU���qv��p��&����37��s|��U���ɨe��7v��안W���l�|W]�v���=B:Ctn5'���!�z�f��D�0�e�]���;��1a�=òF�ǅFhQ���+ފ�|�;�
�	C²���0d�|��H�Ad�ӭ����X��k�c$R��S�/��|ITUɠې.���m�xc�,��onSB���"A&�e)�ا3��c�^jxR0=���w�`�5}����9��ooR����;�,#[��_�J������^Xn"�݄@
Uݽ0��5*:^���#��f^c��m��ETa��u[��� d�֊�}�+��t.�e;wvFp�e�7X֫}��W�bv�\�6�u˷˶�cծp1V��	����,$H�4��I�_��=�}���8`�گ3D���i#�m�%��q�(}��F�b� I�,�^�(c�x�]�̺X�,⨸��B�P\�%QV��W�M9�D6`O�9+2,[�.ˮ�/!�B3D�Mkq���J�2��N
�b���@��6ڟ^x�F>�vol��˦^��c��S�� v.�ڑ��$�*�w=>�;O^��物XK�\B�m�Jcv]�:��#٪7e��ٺ�f�v���Ɍ$TEIl����M�����Ó����@���r2�V[���{5{�������۲c�\�����a>ǭS��한ݞah,~�S��^{�%�9I�_�N��C=b��������D��O��ŝ�+,�X������n~�=����N*(���������eWs��w4�LW��59#i�H|~�S�2kb�xwj����w,���٥]8���h�U�g�T�9D[�j�ً�Ud�罘*q�Δ����V�}bt�|��0��++���5�n��\Qy\32�ҢFJ^Е+��b��<��o�Qm��F������{ƶ�,��sW T:��;�&o�� M��[�h�1ȱ/痎��|���w��$��-q]Ǭ�S�(UK�������@Yg'�.��*n�q�Z�����ی�z�$l�����BC�J��:��*�Y���[�bȺ�W�]f�9
 d��tQ�cy�y��<*��U�!�`Վ�UG����'TfZ���DH)��y��Z�Z.!���0�c)���c�5�]��N�Kΰ�5uC3"��|A��x�a��M�kH�Hj���,b�l���U�c�fS�J�3}�:���	����jx�Z��P��3ZmtVi)�$�gmR���G\X�%���q�q
�]S�B�GH�qV�0oo6;͛�Tz�M<�P ����6ւ�U�r�x�Q�]���5H6F�(���}� v^���1��r ����Ȋb�/?U���B���"G|�MҤ�e�vCW�̌ѱ��#fP�.��^�]�a�h����t�3��x�m*s���ҥ����`,���|u�gۻ�u�OYOD��ٮ�6n�gH�r�M�n7똲md����'d�I�WϨ	��Q�e��]|J�/�buԏ.���q��n�G)uC�k�.�M������(�T;�\�K�q�K�"�'�p���kg9�(F6-��W�Z@���~�u��ؕ[��h�^���������KF�E��@fÓ�U�C���qanv@r�b"���';*��*�ܢt<��q����Ź�)E
XP�a�7۾`WO��O�*!��?5�;��E"}<�ubЮ]����㫠��V�}�0-q�c����k�tBL�q�{�����"��8��9G�'���d�>���Y���3�'n��nY����v]�����z��$y�#݂zF�s t2T�d�}li��s=���)��j�XP~c���|ڼ��I�%��9�_7`fqa�D����͹�qχԤ<p؀F��DԚ�Cgu�F�4	�(���oK0�������.�J�|�x�g��{�%w=S1�sx�<rQ/#��s�¦l���ZS��oBG4�	�z��WZ��q�k:�<�e^�y,�{�N���/���ޥ�;�p��e����:^�-M�Nu���^���2(dՔ2&n�[w,��B�Tш��_f]Úzl��W�{[�!=��)}���S�̋�w"J��%D�:����<n�Vr�����^n:�7�U�˯�*��$܃�u��[ n��m����g�A^~���`��$���b�<���uo9�q
���g�*R��r���TDY�[���"���]q�W�8)�r
A�"={ӻ-��������El�7;s�v��Ñ���%���v8.l���{۲㔅aE[)W�r)uŗ�'&2l�����S��o������@��4q<[�F<Ԍ��y�=�ڼ>+ڋt�0kl0��#��Z����̮5���.�g���;��չ��xbI��i���ޏ0ޏ8[و�S�`�nќ���w��N�G=��_�q]@�ԩ�̤�>�0#�<pʻ{���j|=a���}//g��w>+��;��^�ڹ�WV_�������^�WI��Y�A�c!�ǲ�]�[��7����aY]�y���/��w�=�U����Y�S	]���+c�w���kEyzuG��D���s�qn��:iHb�i�zk�ST���e��c���ɦj^�^P,]]X�٩%�F�%��l�*#
H7IK�S����~:a�ak�L�ѝ׎��-���W����{Ϸy�$���k�w��#��h�~vh���L�f�ґ�3r��G1"J��UUr��E��i~�q�z�bR��y�#_pH1[[u�U�Y"�.�g�����S;�ѳ��U�T��#�h��>ا2I��C*��v���H#ӳx����^�Ae��_!�8�TQƜ�Wb�f�8�o��c���AkM6�j�um�:HU^��U�zJ	[���U�Ӓ.i�ǺߎV�tE�c����W@��g�J�� �ӫ<��7!*�2�$�"�L{�T�e�R�4l��_6���E[<�7�T"���ػ mH�rL�P�q�9v��m~��f�Gs	��P:�֗���e6������JA��G�"���mnw]�uQl�h�<y{�f[1�Fz�C =��O�r�z�ڡsavL+�R/:��R	���;�E�.fYs���[E�v�y7��[��N�i��>��~��Bӱ��Y����*�f;�/v�z/�}��!�:���Z��;eGyj�t�'�E��� l�.�vQ�j�C]As�{���:�ؐ�xuغ-�u����x�IMZk�/�/�r^)kt�h���פb3�xm��ƘJw�FXl�P�S#�lH7�'�ovC�Qȡ�o2��:�z����N]��g�c+�(=S����Е��W��^������]FV�͑L�|���R�0(���iW�8�x���	�j����fS�ݛ�sI�����i��#p�[��:6�j�]4Z������뮲w+�+��G(�;Fv�a��'G�)֭m�6n�oG�ʱ�mZ㙐 C�0z���[�6F��$�������d3�z0_/Qfl��c�32/���b����6��݊����ռ�_(|��YU�(~1�A�ԗ�؝,:���jEq�㔇�#�VGUm��P�@�(T���d�H9���?[I��՝}���K?��dP�������LV���+�ܿg��N�͵��&��w2I��-�!�}6�h;�@�H��.��Z�mΎ����1t���;�x�z��E���V�To.���:��5o�}w�]�"�˼�J.Ot�ӡ�֝yH�3:���T�& �=�k+'5w%jm�s�]��*<Ƅt�l��]���[j;1���b�5�J���C��"�}n���c���Vhy:g{��y��~Ef��qQ��������EJҰ�;�wq�1ע�U2�q���u�s��O5�A�Z��a$�c���)��F�@�k�ؾb1_�%?U[����M�n�&ےJ�t� �gͳ����1f��@������,�{�7��>y�CG_L�/rUҸ޺R1�g��P������a�s!�c�
�f��p�u��g��O@��4���tN�|x�3�{9�*K�͐�d�>���A]�������S.�'&�(�;�]B���12�S�n���t�a��|�w�Czc�N�մ��'5�L���ތ���� ��W�*�=Cdu7@�h�:��b�/�Yo/G&�U�ozQkV�<R���(����:��F���3u�Lw�5��M�.JX�g�)�v-��)Q]����޶����bfTJ�Mc��Zi��=3�	����)g����� ��ТHHX�pǊ�S��\�U��N:i|%�[[+l����o4���P������6٘��k�S���v�����j���v��9�b���q�=v.[�d�:�@���6�c�r�mb�:���,�����=b��F�F�aǞ�D���Z�D.ڥ닷7*.��ƣsJJF�ԯ<e8P��ҟD����3a5Ǣ��:њ�6��L���|�}{]=���;��=ܚ����/&i�D�"&'9�6����X�3PT�`+����戆�l��O��~��V*F�P�	��*eY=/c���@�l'R6���s�u��[:�T!dSI�ٖ�6���<���C;O��RB$�EJUA�y]mb0Y=��gwC8����>��v��9H�b6��BE {D��\ӑͽYy��5R7�1��w��������H҇�>[��ofh8e�Yx��#��m��Ak���/���o�E���� ��k����,�F��7:MxO��� �k�j��+C1a4��pd��#O3is߶�J�bOU����a춸Z�1��|�.)3��3����c��F�|%5��ܫ��T������Ι��6%�T.e�B-yJ�^BP�zl0p�]�w�����q�A`.���-ͥz��׀�B�e�����i�͕9�e]�bN�����V�%q^$hȍ������"�7+�����95�\�{�.qY�/���m�%ͥA�N��'��iЙ�Uf}�}�8�ﯱ�R�X1)P{��gi�c1h���[]�a÷;��L�;w-�^�Wn���WSE�iE���ھ,J����]h�]��Ǻ�rK�j����%�-�e~Qk�obwn���
��;f�I4�:��x���B��݃0M��l�ݚM�;+��YJ�}�9�xS��5^�X��|d������ v�U�x)tG$��O8]��g`lgI���\;-��M��곎��*��0
���&g�3�}c{��(�k>�|H�}{�fS�R���(�<�8�]^�ǫ���A}K*[�)�w�����`!�^�0<�jq%��2�=z� ���f�5��aq�{��>��n�6��J�(u�J]�˘CV_�W����Ϡ�񤰖����vR�!��@�N��:��9^�#w��՝�%ӫC��u7���lQ!��滶�7ܻ�/P3�6۵bh.XY
�&�z��O�<��:+Â��v�d��
�{]un��zۘ(4n]KR*	��y�+�J�	uRΏL����0��*���-�ǰ�n��#�.�v��ҷ�֩��=W�Oa��j����=�7�rݥ��q�v{u�>���V̭,h�]���-��ysW���ӡtKJ��u.��9�{/�	6�sg���bV�\�R�a�"�g7<��_:���t��Y,��ˈMvs��S9�nr�K���P���z�!���Y�@�./�ef�Q)�WR�}F�vp8��\n�S�V�W.}�x/�w_Pb/V�V����]�W�\�=��p�+��%|*�:�.����eX��tԞ7YW����Ň0D�p�/36u���R�����\6f}%�5���qUu�Vp�mH�zQ/_]�.XT�K��h���m�,Vr#L�%v,{ΨX�XƎ�]� ��V� �O��rv�u�,8�c���ŗYcWo.ՖXJ#p�5��CUp���2mEս9	�����ѣ��9t:��[|S(�,p�v���]7�+-�\d�.���ݕ�0n�E���cy�U�sW����X�3wJ�>�=����^h��U%�3o�e:��Z�Y7��)�b� ���m���Cj͛�4�; ʝG(w�ȀξA��Db]dB��@�ڋ�Ñk��ú�vB{�he�ŏ��G�9>(�cnV/�f�����ĕ�^�]tұ��R=;^u(�;/�N��?��i�{��	�c�+��{C5\Q�趐�l:�F�t�E�x>�%J&�j�d|�M�E
 �QD�EduPT��?�_1�!�mIӢ�HQT�w��h��mX��ӈ޷5em�U��a�Y�GWL�⊱�K�a�s4�0��8p�m�L45V���&���nTE���LTm��[�eW2����.b����m1�N�6rV�j��s�;����2Z�M�&,�\�&�MC5L��Uus1G&a��M8��V!�Z�Y\j(��~љ��L�(�ݦ���iLe2�\Eq\2�j�"�Tp�ӧx�m�LL�U�C�kT�ZV)V�3s4�N�T�e��\����W��>>>8|+*4�˖�U�|���9�W2�K�j�,�b�fV�ɘ��Wqi���Ey����h�F"�L�r�مkX�̣��+�Qպ�"�W.>>6l�<-��i��^�:�檮-��k����LRҪ��Z�p�%2��h�Æ�
���8�m�o.�E�mu�>��J#-��%Q�r�r�¸�4�J��YVֶ�Ub����(*�7-[�孴*4S9��GQ����z�:�r�87Ty/�D��v��&��C��m�,o�=%�3�k�o;\��޵��mF�bm��;�� 0���W�������WY��H%]%�������-�#aߕaz�V��e��֫͵I [7vi��
��9c8��`�2��7�0q���ߋ�k�"gk]a���ˑ�2dlm��uME]1y)�F�8���w8���*����"���6�v���4�?-�s�Ȋ� �G�H|��aq�}�L��-37��Z/A��(pep|��v3����;��3���Y��TW��e�&}�|�7-����+ȡ�vС٨��2�d�w9�p���-�#5�_M��nT`B�twsv	W�т�z�C(�B�9)W�U�f�hs�UfD�lT�e�c¬��<����+0!~)5��\y�����ʫ�K��<��g��L��9Ae��P��:G��T
8ٲ�
wݖ��f;�D^�a�ި	�6���|#l�q�4���\���.�N��9^�n�ꍥ�r�G�
�<Da�����3n
�osd�Ԯ�e-�z�^���o�N�XW���u�mh��j'����ܢ��$ܛ��#�>M*��
�z�z�;�{/Sի;�t��N��'+�l��o9K�]���j�t2��Η�;3��|;�yw�5�E�J������B�uO����L%�$em�/�~9os�q���b��׫��sU="Q�\%um�mi�jF�.N���4���w�C
��7��@VRZ.���~���t��e6�]y�A�w͜��:����J��QT�r��O����ѡ�2��94��&�)A�yO.���}Ws�x�EM{�
\�>Ůl��R;���ڦj�E�fT�ٷ37�;{DSHԄF�ʞ�ا�loZJR����c�vOӤ&���&"�s��@gn$L$$%0�0C������&��;*��J���2^`�"�z%�א�cj���1��n
2"��U��Ǩ���4͡���`Ym�P������mu������� �R�s7�r�}��u��<0x�3�l�euٷ�TM�gm�0df���`�<4�[ ��E�Fߋ�٬�z�J{�r�gYi�aK;g8�R�sp�MԨ�:w�m��U�[d���^�(�� +�����D3^�^�rU�r�u��u0���5sֵ�xYJue���l�.j��r.�-m����9&@ؑ�A��d�n���]awﾮ�2M��`��Z4�=#�q�Klu1����#��eCt�3�Zs6z�Bx�h���Q�|�݁R��;�\��9�!�]�;c�t�wP!�FW�ΡC^U{.D�z6�g�t���D�����I-��ȍ���b}��E+|�g��P*�OH�UYꍊ���|AqO�7�vZ�ƺ�㾭P��(�������z�/���_�ad�sc=ы�.|*��Mm6U���6����=&�g� ��~�יŃ�<�܈K�3�9H�=U���l���{�ve�$l1��"��-t�n[������*����f�ۋ�fCq��܄����H��s	!д�a���k�]2�{l	YqyZnt�E�[>�Z�˰���TJ��b-�x=����=9����o���4�]���$.�O��&�ĜU����I	�~���Gv��;�m�A�/hy�]}�5b�/i�`�������n��҈��c)%��N�m���՚4��,w'Wطgt�2�4����N��+u��<��{
�ݻ��v_*^F�Cũ�v-a�\�pS�m��׽�,����%��Ы.�(�n6S�,��-�OI2s��7U5���#������9�Ґ��P
�d��0��Fl�]1�UiS����˔u�+g~vՁ��w�#ܿz{hM+���-����F�s�Z&ֳ8��\9`l!�Q�L��#A>�p�gg��qf����I�ۜ����Me�n�h��@�v.��5�dد�Z�G��%�6]�q��"��w����*Y5�uDa��E���n���m��G# �����aj������0�H�h]B��hp������Q�32 ��	Bc�}��	�?%�;���T��e��:)��E��	C�ɯL�M�m)��ٓ,sN����n��*�n^�T��SU�ۚ��g�A���?B5<{��V��[������B��x�C��&��e����X�
:��/?S6�+��**�K�]� �ȏlu�"��֔�l@V��곃��¤�hY�L�V<���NE�s"�y�o�|n�X�l�Z��gp�B���T�:��"�|�VS}}.r��p��{���E9h�O����ЏL�:Ӽ�ks8��.�'��?"YI�.�PT��7�諾Ysݝsސ�L*R�>h��BGb�nAH=׉䪿o���!R��6C2%���}����2�l�����IbA�B �*Gt���%K}&��f>�Aq/���Rs���)0++�v�>�t��c����:�����#x2v�O��v��1U��5\rz@����M��^�#V�tv�Å���+70�>�ӹ|�r�'����>�[������/@��pӫ�Y�6med�yWս�zym�j�(¼1�썯\e��6'�NƊ�ئa��6oXt��H��>ٓ��k���(��UbUeJ}�{	��|܍�=M���^ptgPq��\e�z���l�慗ҧk�sr}!�eOl�Stӷ��{p�\ ��?sro,�f�,�-�h��K���,O	u�mÌ�jQ�+PgxC�Ǵ$��n.���Ѳ�6iWP��Ǎg�1Ik����<���±u`U��Y��S*g;q�ܡ3T,�޷2p�6S��~�±J�Ȩ%.��g�uzN��n͋M�"��ԟl:0��p�lTn9@,z�.���)J�7��D]f�ӗ;V#/g>�d��!�����ӝZK�qu��! t�p�gb��!��;��srH��k5��%?T��*�����4��vE��(�*�r-����y-c�.R#$nj!��x�of���hwj�{7�K���!�HjH�m|6��e2aٺ��Γ�3o#��:z��H��s":ɨ��Q(��+�#�b��R���@Vu�};����i�����UW"ժ|��[P*��&�$��"������R���`j93�
ߧ�=�yFBsR!�P7�v.کs6�:,�4c�'�Wf�z���1�GK��M�c���r��	�CR㽋iBɿ�/�z'�g���.c�2�!�)7J+�q>�-��z�a�՛��[��9F���BmxW�>�/�Fj��`'ص͝�!gsrͻ����vm����-����N�.;l�D]�x���˱��g'���ճ܊�7����mu�02�ި2�Y�������֬h�Ⱥ�"���7r�e��΂�]l<��.�
B��f4c��rB��JW_	�e�oe��u���u�P	���N��n��S%�(�__3B��.����Eٗ_���]:�]�|Ι|J.e��1H�5���Tu`d�b���8�ln�j����CZBL�^���p͏pހf6�,ҡ�ǫ���t"Çg�!@m��ywU�كk�H��T��#ﯰ5@�7y�\������oW��,��5�8��]ܓ�^F�$�1��zC�Ch�N��<������b.'sv�y�7Q�*���x�t�$�8$���26k���]�\�j�g�{������&������x�j��O'�Q4�`��1f�;��U��V<��[�$\l��0!�E͇�djj�r��GP� �T��65ug�����۬D\=7<�\u{����ꧫ�6y��������E;���3c��6ݽ�0-�(ٓ�'�D�U�(*�Y�mZ6)-�̶����Lm���B�w4zI�DW��4�4΁�:E��}U�1��[�	n���w�:g�����U��4O[�{�+��;���N�#��e�r�H��?2omj1pw���%�*�/�;�T�P����g{I�/���g#AV��yҰ(_:ˡA�,#*Cqֽ겇����vŪK(��O�������s���/U�6tj+�c	PH�0MS�@[��fYWȲ�iy6�虡�U�O���lF�p�$��RQ2�:��|fkj1s��1WG���3�A�䠆��K�A V�T;�뒩t�:�M�;��Ч��1y�n"���v�hG/��s�G 5S݉I��:Z�$m(k����`�"�s6}xL��S����'�5�-�=~�s=�{}�Ȟ�@�dL��I�3�<�r�j�{��B��oc������s��=/g���y��L�)9�
l�����	��%N����oӤ0q`�����t��]���b��8�����oiF�GV��ʊ����l1J`��]C+��1����!�`B&Ly�/k��c-4M���1y[L⩄��wؾ]����ͬ}��n�4��;�6&s!�n���q��\����i�Y�T2'���$x�4�/�÷�y�+���ݽt�G�Zи�	ĺ���v�5�O�z������h4>ef��3����\hj�nWV�Ya�.NNQ��ա���U��Ԧ)�bV�M�p:+(��[�oh���W#d�&�fj�����E�w�\���4F�ཝ� ח��9!0�^���̺p�����J~�ë���CL��G�������Oa�P�A+��1ѐ���vi���Q��ꍃ�Q�R��ԩI[f�^\����S��,��� ��8�[}o��C�C�J�������Fh��z�-���r�*��a��w�}y��ձ2���(@��Wj ��z`�K"Ug��^��ѽ�Y|ۦ��&<zB���C&��"=��{�%la'Ż=a�4oq�����I��^
��!� �$W�EmOl�˳Z��3ôm;y�7d��f��Τ�mrV�Z���� ��Lj�ׇ�/*�������v�G��;;��W��}��ެT	�<�:�����_@�x8�}�n�An<{�a�d�\���H3�PÓܺ4x�(�	�k�_�u^����J\��#�٘2�d:Gx�]�۸輸p��|�`��ݚ��x�'Y�v�qfA���-�(^~k������4`�Z8(�Tq����G��23d�>~���t�����7)����us���ιϷ��6����)�;ɩ����W�����]�K��=�7�:s�ȸ��n�ڙű
�6����P��f���:�[v�����ٲ/�ү0l Ϡ��. ����l�,q��[���[v��l���鋅&A��^�ϣ�!�{�0�e�F�<�AxO��̩�޽;8�U��� v��@���5P���}E��,>z��k���<�0�]�y�H�H1�,9��]�+o ���BLV�q���f�P��(�oZyJogic��6"�dqzZ�g�)N�#%�[�S��-��)�GR��Z�0����EV�̩T7.���!�J�QƑ�I�SC�`�˰�S=���f�D5�T0��s":�{|�B�	AHWs���0q�3sa���������4�"�T���Hkd6�S�k����MK�a=Toy
V�L���}�n���L`OMUf��POQU!��٘{��GcL:�y]��Ƹ�.k`]���j��J}���S!1�J�E�r���z��Ǿ୚�{�4��[��ȈcQ���rp�=� SN΀z��Y-�YϮ�t�Ř4��D*��{M�6��}����-ѻ�T��+�]��仕���F���9��`�94)]u�VY	���},�t�<�K Jp�N>�2�\��um��GKkx�e��=ܾX�W���X�d2���Pݨ��/ot�\�w2
�"crwg=��ؕ�:���8r������
NJ����m��v�kK�A�B�=}C+]nb8����d�%�@
x�V�Օ�u���y��I���>���Ǧ�t��Fmz��|�}��V���j���B+�� `��G6V�һt���U���u�3[&�p���`v�q�Gjy�u�˘*��v!������䳕vގ<�v7���r����WYj�
$�&z[������+���!y���^p놜\��KVw9���N�G{�/�qPl��M�[��X���op
����T�@�B�(�G��X�f_�����c�4�x��3�fbw-�3(Μ��kg4o�F����^k��W%|�P|w�;�`'���)wo �./�m��4&ݞ9�����e�G��C!�rϣͲ���\:�n���AR�������vZ�8V��k�CK��XnsM��.*��ε�j��X�2�]�NjkF�h�N�}N;���VV����+I�N����W�y6Dw�a"�Ӽk�2HѢ�H�� {sf�����UinH�:֮�f��*��A�ճM��qi�N�I'�jLo�3�#���4U�j��q�<ZW69pR�e�|�s��F<̰�$�.՘�S�uZM��(��������s��|��uǃ8����=�S��7�� �v
�Μ븎���z$$��\�w>Y���nƈN�7��J���1�(RF��ݛ����*	�I4!�֦�����]p�aů�+Φ:��R�P�W[s�J���e�����T���PJ�+p�de��sˏ�{ꅂ�wk�+F�VM.���u
�o�����8��XH�@]c�c��y�����z^)Y6�T�W��9�̕)��z�=!H�;�Mla0)�2Pי˹N�R[gh�����V��QҤtʚ�Z# ���'],h��X碈F���se��za֯�A���>������6�q��񱻼�)	*�9��t�,J�a�޵N�ک�r�4-�#�ŝ�f��xT�}��&��Ue�i�'s���oY��M|�h��Q0*�p���E+�YYٕ�<8��(n�2Y�zr!�dz�Z�����∥�;w���pZi�|�Ĳۧ�N����`�����n�6Ё�74ǽO��i+�N?�EW���3�93p�:�.z)�(�0��y-� ����P�Z�M��%1�^�tum�әx;\ʭqDi���p�O{��m�����c�����s;o�'NWw[y�&�7���[��pC��7��>�Ի���hi����4�P��kX̫E���Tc�0�"-�U�k�VM%Ka�p����Å{ g�]��GN�Z����[j�h2��ة�̘�kT\Kmn2fUVYp���Ç��It�QWQ>˭6��bV��,�-��wlU��EV�WT�3Z��M�:|l�UW��Um��s.6�Wi�ˁ���32T\[h4�Ȭ�
��o����2���:|lై��Һϩ���&���jTʷ03T��Kjk)�J��.�GM����Q5��eK+�4||p�¥$��5�ֹl��*QV&0�fT�kj�U6�f�P]�m���-�)�0C5qɆΝ8p���å�ˈ�ي4p�EZ��ك��.i�3����B��9j��������6��[�`�L�>>4p�ˎ*�8�%ۼ5���uL�u[p˕QE)iJ5]7l�sن��̟�r�V��˽]�����k(�.o&�~�͜.����r�Uer�.\2���-�0ˉ�M˘{z3W32�Q)����������&�[u�*U�2��М��[U��+�sZX�Y�L�r#.Sy���kW�5O�P��ѥ�21��PZ�1���U����G��r�)c��F�P6�e�k��(h�Q�64��r0w2e�#�G"^]5��	j�9
D8�.׽�5���EY�ם����&�J�E%���ԧ��4�	���9��B����,���b�i�X^t���q��'�.�l�l��5�8�̆�J�5���91�v߶�Qñ,�&�V�ڵ�|vu�Ym�k���������-%����Ѫ���OP�Sֶ4u�����c3e\\��f��'ξNё�8f���y,N/\�s�Ь�rD�a廽�X&��/Y�v�T�t�js�F���b�tI�9�q�K��-��7Q��|v?N���!���g{df�m�h�p]|#�b)5;,�U�����b�79#��P/��� �1�$�d1��/%�wD��.����>g�ʅ���� ���8�/��4<m��D��{"��e�����0GPI4m*�9�_r"ADp���-����&lydzRȴ{ٹ҂*��}Ai�BlH�IVVh�l+�{AŋǞ_��Y��\
�����ݩ�v�������z�/D|�3׾�m��8>ܺ�\4
��]�+��pe)�:چ���V"�&�>yr�ǲQ4�v�o?>;�w<!�~��=�Řܐ�a�@"�xQ��hЊ���x1W�y}���ψ�N��n��Qy����(X�(6j�lL�m}�}sIO��Eޞ��޺o�mA�QC���ӑ0�N�[b:�Ig�V�=��^u19}�*��f+b��Q�=&���c�K�_���cC	ChWqi#�5?^ci֙>��ȁ�v[RDI.(�5^|�»q�1�i>�XڍS�������Hl��KC��gF�H�7e#a���Ҥ�ETEN��/S�y(��l~������� hJ|�s��_|��V�k �1������	k�d.�06������`�u���V㓙o%g���ƭ������+2�׏w���D����p�d?-�+�"�D��+q����+M�eV��V��PU�>7����[#6nЋ��]�z^�P v�׆o!�n�&�%X��Y�Vk`�`�!y�0Eo��z��3�>�{�/�S��<�lo}�����O�Nz�f�m�Ifhނ��v��i(��O�����Wc���u;��v�<��n���x�9K��E�ﮡ�ʤAl0B���aįxy��N�wl5hLn,2�����'G5+*̄ht�c�����[	��;+���8��P��lWG�b\���+ǣ$ooi��z^�����-rV�R������
g��
��f�G�%	H(l�Q�v�y���[�;qOt��"�z��\�df��0�Q�"��c2�6��s�f+��9nS�E]Eh��>�Q�|��t6@�f�%^���]Üȧ悊{�w�0M�7MY��E�xHJ�-"�k)��;�J���e�m��X�{�=F^T�UM�<�^UX
�i����7R�D�-Z��7�� 6�1��fL�3l����Yd�T-T�ܝ����5sƌb���f�$��ɿ�a_p�ɲ�XՄH�]>nAH=�'�$.�"�W]rY^O��b�-��{'�.�_�s�!#�Z]�t�	N\w?gT��YR��t� '�v���hm��QX[�����4o}�������g�6�n�U��� [�:�R�t�6�S,N��oeL�*oԻld�ɡ��돕�����t�eN�Xn��b ��G�3z����D���v���� G@ʒc�����c>�,GWHk�S��P�<{��_e4Qݞ}ZLq�1�t��=��WƑV�H��>-��B�pY3L���e8;�5O�[к�ٝ�,/6�'��P洉���#;[}P9�:�S���S�Gi��\����;���(�:v��HW�'���6���{i����{�S�ó��@;㔸�R"����	R66��ܗQD�R�[6������r�N�vC��̯9Ay��q�b.2�/�S��l�̱^�E�ƋP4���ٗ��׻��Cns^�]lȍ�F�p�'Rw�ˇ��H>m��E��FW]��3�G]
�����:�3���9�[²8��s��ZÆ������*"�,쿘?r#A �8��,�ا�!��<�dimc�(�{�������:�5^R�׻��;x�Zv�E�򖼹y�ss�4�@����v�	��:�D��b�׹{n�%{Բ�a|m�A()
��pWk1V���U�X��'z�+�>Ø�\�Fq���]`̍�>�^��هZ�+��[�i�[���.�l1�M�8>�w���$�:���5�ۅ�GS;�ʸ�w	�-��5ګz������H�:|8��gai�y�n�z����C�m����zr��į�,q�����q��D,%%��!��&s�l����'*�m��H���V��X��R�����/��T?��7V�q_q�����U⌥3�j�S��g�]9�CsD7i��Θ�����8`�с�\��q&�t �K�R�n��]'#܄���4�К�eI�=Ż"��~�vS���	-n\F�3Q�%��M��e�S@z5��E]i�aC��>�6 ۅ#m<xm�����6�l���S'u�޹���Ʒ�%�j|:f�����ñL�<Zءؓ
C5Z�Ud�K����g�\{u`Ȭ����f��2��vX]^�뤓�۫����z{��'6zj�:���������oC���ܺ,�������_Uv�5^T��q��-���N������}��j ��Z�>��>$�Y�;pͥp�]o��+��>y����^|� �	�j.���+*;�o�˹l��#m�ɪ�����#�à��S�Sv��<���t��xw+���?�ҁ=ab��x���櫝%����v�yb}�t�M2w���(ߧ���$x���I�=7�4�y�H�k'���Ux��h�Pd�ͩ�46�͛�ʛ��C��)w���E����F�Q<�øq�ļ�:,���gdZq_��dL3�PD�`<!摬��'8r�X}f��m�[�bj}ow��q��?~����
�`X#hâD>��s9wi!ә�)q=�̮����?z�wQy���wK8�h%OU=��6ԩ
!�'u������k���ܯY ɵ&�Q��7�u3�����AP\����A�+���e���Q����tJ2(�5�<��^tK��m͖Q��&��y��3n��	J�F���/�@[��KAt����	��\!8�N�j�����Κ�|�P(�
~�� m�{��7$��J)cD^�G�u�@T���,�����s]�~0s>��xʼ�/+�ˤ�[ܥ�W�q�]�'l�6/Ws��vb��xΈ%�y��Y(�讥�j�o�n4�}Ӯc�!v�I\�ʻ�z��(�YzR�B�s}����K�X$�M�L�?��u\�X���$it���4�B��Sk_O{O���d�	Ř6<�Rs��h���#b�ʮ�$vIA��v�V0uJ_�����ٍ��5G�[d��0�0�pt=�v�6��v��L=��~���r�/�zXTJ�Kx�:С�q��>`��owF�����T��CU/{������<�w(S��r6}�n#m���;t5�g�3n�]=�ϛ���0����4=�4��W�]�l���LεkD^�*�n�t�iӞ�m��v*��;ڑ���=緶��<K��˙�����ݐ��j�2�Ms��#=r�@]z,>P�㧠���2��B�Zv�f�VFO�E��o��H�e�Q�l����\�M���N�e`��7�������i4�'�KA�Q�/��: !f�iRk��	-U&FUu����~����D*�!A$[=ӹ�O�;�6:l<D�ҙ��Z��N�a)h�`o(�j�d�(��>�YJa]�Oj{c B�#��R�]���Ѭ�g����fU�t��Os�[ٵ�c���c��������s+�V�Q�j�h�Ō8C�VU�ss:�o!|kMA��M����|!����v�k��d�lNrML��2�3�����.x؃�ݺ��s<�,�UP%ڱ�/wn��V�����׶�*���+�IFR�U��L���ʭ�=����V�V��}�lH�XD����� ��#{�}�"�]�C�a"��;�a݅��6�����v17cl��.��H������$��B�qE�?����ɞ$����N�X85�aBڞ	4ښ��Y�뎶dN�����o�d�F�W�v\��n��49zM��@UY*)O�1��m99`68�����@�x �؝�]X	��#v��tƪ��������
aR:c��;�����9:+-��խ��;���Y�7��&%��V�ͫ�|��%3�����،[��co��.�������fتѦqߣzS��p�q�8�f\e�&����Df�՚�nZid�/��pu�X+���W]�}�\�0�:���Uj�gN!�@l4��j�*�Xsb�k��3���#F�T��u��%��d��/7�pk���S䉁[ý(������"�ʕ1>
�B1"y-Ϗn������}����ev]�Y9;��f)�]�d@���´s9��d@WZi�'Mf�o�[�x�=|Ǯ�����uϷ�dv���I#�����xp�MN��45�l���iM�<��1�ك3ۖ���`C��o�*����j�� +D�?/ݻв��'U2; :�O7�n��/�Gq&�V��E�
�KY�.��Ӌ�x��׽�Dj�7E�޺����
��JW������u�RBk�Fj�]��#������,��bZ1�ud�����PWa�����Qq��WҘnMC�UCvE*�}ݙ)]�Hݎ�o.%u��XwV"�`����WF�B�7�u8�W��������\��JL��UΫuV�3�
i���>Y��P]�+����x�!b�n�IR��P��\�6z�t��lK��xW5���������FK#��úJW��ƛd�]@�+����ln?M�{x��Pg�A��A�P>�B�n֚Wx7��H�C��$�ލyn������8Ro����:���J�y���݈�e��ٻ���Z�H��b�j@�8�2���]1e�\
Su�H�p�d��I�4�}5ح)/r��;�r��飫�}���Ta�=�g����-�^�X�nP��l�4M.V���2��f
�쨩���9�Q�)h~����&3" �:������u����<n���(�"Q�s�~��qp�(��Wa��a�څFDF�&�E���槶�Pv�*{1��7��s`�	*<jr}����"lp���UӒ��&���75^���+����r��}[@�F5�c���� o���;}B�!c���vՄ�oX� ��F��{��K��TH�Zx�I�2=���(�x�6�HÜ�cvcY��em�@n�쳅�7F���nx}l&r��DD���N6��S_;HG�_G�h�pE�v����l����C�[z�U�K��~��+�8/���q�A�\�2��
�{��*�r��>ia�^������d�Oi�ً��8�Fk�^:�7q�ݛ��5q���۩�����{�v�'t�J���DW�����DQ���)�� fӎF)P��E����ĉ���@@ �$�A d�&�����B�@ @@y�h �  H �@�0(��J �   �    �$� � �� H    d $   �0� �   @�f  @� �   � �H! $   H  �@�# ! $Q  ��2  �  I� 2 �$  ���� 
F @@ d�AH�	R(�(F "$�� 	  	 ���b2H�S"U�����5��j%K�
d��2����g�����v��w?|�v������t?��~���i~���^�S�=d�U���y��������R���=%�-�ӓ�~�Mؾ�E*�>�������.'���n��g���u�c���� �$D @ � I$X �`�	0�# �� �#� "2I�# �D@	�,�E "�J3$
3*P;�QZ`@��   (@�" D� �B   , 1� $1   �B$`�#@ �$���$�$A 	�" 0��0�$` �H� 2H� 	��F@H�$� $@B2 �  !"@`B I ������"���S0�BY�:����̶�뵎��[�ФR��KV�N����[��v�ㅎ�\�)"�{�n��=;^ß���J��c�����H�]7��n�)V��g����������YKOv�W)�L�-f��H�\��v�k���)V�����C��m���z�[�~7�\�</���H�^���{$�U�Z���0�^~�7;Visx�}��2���o}��|$�U��̰��2^����:{���⺤�Uֵ���\��U�}���վ���A��PVI��A>WS��6` ���������;�R�T)T�@�������D�H�tJ QJ�@J��UT��%m��IA"���K�$��AT� �DV6��e�Yi۪��ZSk���V�,�+-���m��kEۻUvf���h�T��eݓ��M�j5��2ִ��
��sU��gv�Z�޷4�ԘeRi�Vj��ث1�چ����͌���6��f�Y�J�̱��Q��ێ���4ݙ.���6�kb�U�5m-MYKS+i��[�sl-��&���   �{n�le'^۽��*�������`Ub�y�y�[�z�u�fk��=�딠�{�{�Ww�Х^4��{��n�`5�ohz��{S@zm�*�OZ�SYF�1j6   mw"BE
	�0�D�
(����(P�B�
(Y�\:(�}�}�s�W�4�
6�{��n�ۦ�F:���{��{5w]+��)]�\�����z��t9C�J���֫��,�m�,T��   �y�h9��w�����9^��6P��e���E��w��ӳO�m��OuTt�ڴ�s\��u�w���N��kNj�ݻ�Μ�:����M=:�����f6i5*M��f�j6�	|   7^���ЧX�M�Wu
�=n�;����jںuSl�ú�ځ�u=�4�F��pQ@�h�;�T���t�Z̦h�B˲�l����eMJ�-�ke|  �z�Q���Ǝ�Y��
��;:��������w��[w�@w\�U���]j� :mv�$2͗����VlM����  �=)Z�tAڕ�P��tP����ֻ3n����v�n�����aT v�� �WnwXk�ųY�6�ر�Z���i���   ��i��P��IӗPP룳��@ s4  .�p (�c� wJ�  ;�\  ���m6��Mts��1l5W�  �|��+�,  �n  �S�  �K  �Wp  ��  ms� ��p  q�  j�jYU�M-��}��"����  wo�  �]wC@ mNp�:]p  ��  r�����@
�n  ��i�:.�] (��i����b��V����|   ;��  ����n�  �v�
 wgh :�� ��( �mv� n��  ��� �)���QP  E?!�)IQ��i���BR�   O�JR�  �{�4%U 0  $�TT�  �O���G���3��0g��f�����i����-�a��z>�T�U�$��܁?%�K�����y����<`1�����cc���co�c�m��0��6�������_?�ŏ[�`��Q�µ^ڵm�W�8�CA�b��C�ҵm,���I�:�@�w19�H8[�V^!v�TLԝ�qӼ1<�&:8q�_GB[�A�f[��R�,]j#+
I+ݰ�f\�aa)Q܊[Z�V�U�l�E���$�q��"����M$(�i��M�,����4��0��q,���tJ@j����:�-f"MVZ���
�b@�Px\��-Ll��a1F06��u ^	N�u�b������	�Z]�[�(�2��%l[q��ǑV+Cz��x1�]�	3{W�Z�ˇnmۘ��3lɂU�Nd� �\?L&�)[�$�i^�\fJP�ܫ6Ry��'6�����	Hf�`MV�wh�B�i�V����j�@A��	�tKM����kM�E���V�u
�ڥ�C0kA����ٕ���1,�3W���@dө ʗW��j4af����F�SL�,��9lF�+��h94l�ىM��`�.��yG(p�e��T��%ҭ(�F�89����p̲�{>t��p2�T�zE0���$���[tl����ⲕ!�9v1	BҬ6C��50��y�bH��,�`���"�:!�]�zх1�agrQ�Y.�b8�j�B�&���(ݡ���˻Wvn�7��mƾ�Y
�K^�l�z
�-!U-���13���бV�j[�
m]��n8F\�Z�8aچ92Q�J�vF#A�����NJ�J�����e̊�
�
��	�Q \�Wȝ�On`�M�ҵ�.a8��hV��B��I��ҋ^è�,-��3e,��Xׇh^%0��SM�nT�?�d���X�n�āe�w3&�{X�0i�Y�l�"eEr@�v�.^ �=r�m�:j�`�BϷ[)��4�c���V�������f��)���l�;�C!]H`z��Z�Ҩ+HRK��I4D�VF���	fh��'t@����z/f��-3p\�գW������6@�*���n��	��lgy�ʀ(hF�4k2�;u���^�aV��'91����9�HNZ	���M�J];�x�fb�1c����5E���
����l�n�!��ٳyH���ӷ�{-�x�"*�lh�$U�cnj�WW,Kki���4�X	.�YA�0(����R,:�xC��պg�S&�6�ܩD���yC��ʗ,c�e�V��3`	�M�zN�U���u��m51��j�\Ҧ�J:k�?��ӊ�U�.��e�Fjr����J�2�1娪a�Z�7��I�=qh�T�;M�%彰tԻ�1삛xcD �t^X�����a�X��3�F�7����b�፬Ti`�P��&�7�e*��͂�*f"�b)�[Z�ְ�<��e�֥����f�l�.'RP[>��_@��-(�A�h�Ef�BD2���ø�<imC���+̍�Q�-YwW�a�3M�Ű
?Ӷv'��(uaCZ` �K̴lS���5�QD��.�Vn����q|�׎܌�N�Z�`s!��-⫶�A;�sm�mb��J�JR�Mc��O2���
)!9v`�z�n<V#�a)G4B�[`�6�Zx�L�(��U�v(6lc��U���l7X�9CC�f�*񦆢��*Z;Z��n�w��)�w�b�,�Qɕ5�:e�'I�1 �����+XH\����mԒG��ol��zj75hC[�"u����#������&�԰��s@���_ѧ���ѬP8 ڕ�IL�$hՐMDf�f��"���	F��\	|و%�R|����"�ч%��V�EA�"��!���Їh�^4橠+F��b�Y0��/45	Og2���*�M�^aw������&��u���kyMހ��+w[�$p��4��m��3X�h=Wd$b�Fr
�\��[524�4v���n9&�Ę��m��b��&�l�e��P��fV7(9LH�-���,oI�+8�]�C$���6/6h4;F�e�©�	G�����D&|����Ս&�j�I�𗸄���ۄ�5��qq�
�rf[��#sX�I��U����չd�,�%<���[WM7�9�tX�Z�H����5�*�Z/V�F�4�B�L��*�(�4�sEA�
�݋�0Q�]X�Sw�
[&�X�;�]Q���cu4*�@d6�Ae�TS�ȝ������V����р�� ��s�j��{W��2��"�����@L9pS�c�1Uu��Uّ�xk @J��r�6�Hʬ�&��S�n^�[Z�kT�	Co���(Α!�r�n]6&�6�u�`n1-�Z^�)
ز�e4E�z��)�˴����SRY��Wh1p�`�
X7yX�A���U�w�(����6��{����zv��\���;��+&����`X�R�ql�d�jbP`HbӸo^R׆�%�'�K��`�w�X�N�	#�U���)���d7L-��_�OP5�*�5�wz&E�f-�e���Q�8�T�@��ƻ�w�1��JG�0�0��+������պ����"������Dgk]nĔŗR���YN��קrX:�YҔ�b=��،�������]����ͧOU8͍��V��X;�i�hf��L�.;k�,/�KnI�1�f�܄�aZg�dV+t3�ţ���jm�������r�t��	[��<��n�yw'$2�\	:��n�
?2r��MO��i4�����W����0�B�I����L�;�������V	��Q��i)p"]��*n������W���y$���)�Ghi*��Z���[��0��dw	���~_�41���2�qA*��IWu�ԓ)�W�5�[!�ܼ�e����U��3 v2�e(��@�x����N��l�(��m*;[��FZ�{�D�<����n��u&E�9h]Y��7˸]|�ںi_�ۀ���D��p��)<�z�)�0-c��P�+.��V��mJ =X�a���b���Pɧ5�:�xө�N��CN��5�7�9�5y��,`���A�ԓ�un퇥'r�&��Wdd��I��b�])�Y���j�i���,�Wm�^�F��W��Ȑ����o�Âa7*<�ASEu�-Vs��h����bc��pD��`&�&��d��*-мɢ��gth��-��6j���F}[�mM���'[Ia�5��$����Rfo!j^E@U��+i���'r���(�Y2��t+T��'(&��	�f8Q0���2�q1QWwX�F4�$�5<X{M�yn�T�Z$�J1�,¶��&�{�pf���C(��r�6�ۦˇ ���ҙf�vI�b�A��;���+:HThM��Ab����K��U��v��-˥wBL����{���q��S��d��jb̈VZNJJYA
�k��r��kQ��kr�4��7�e%ة�B�{wgE�V��e��V e�"6��h��!q0��ֲe�i��c(:{a�/]�@��Bp���۫��c�Xσ�����)d�k*@����d'2C+�\vЙy`M�Q�\f��HL+�[.��00މ� ��۫���	�x��¢��s��+J�v�8�v�Q�u6���D։�B���r���ޛ��lo�(6:1C{qJ�m3�,7�J��q���y���w�L��o�x��ؘ]�J+X�[�rSný����	k	\�W[k0-75L"r��wQj
m�*M���J
T�<�fFe�S��IN���L�
����l"6e��4�G0�;�ڋ^�b�d��2V�l8jKKb�I1;��[���J��4i��U ��2�*ݔ�dr��,�nB�6ǡ�b*�v�	�(-g��v�; 7�P�p[n�ց����H�Xy��0R3e\55� P�ޢ^���'A+
a�<X��%3kE�A^[�������b�ۤ.�]�㢓շ�3��Sg2�Z�ԭ]�w
��1�/L4�ixtҠ0+V�m��ڟF���)��O�ں�A(D6,R%�o0��5�[��U�tQ�6+�6�T4��������6��(�c75XwzDe6�2pݓ1����A.�Hh�R�c��ފ�v��m ;��f�n��u�^�c�Y �c�����F=WVҵW�kDB$f�8��ɵ�L���ٱ��ͫ�:�
�[�wVv�RN�v�A��ѕ�I=�4�!��ԙ� �o/��I���Et^�5�#*b�01�K]Mͺgg�"��Ӈ.d&� ̄��5�V|[ ����5B n�ɶ�І�^B	9������J�l�H:z�Pf��B4�:K]:ؽ���'����PGbI	;�jĨ�JN6q����7��=��:>�J��)�n��;ġٌb��D����7N��3n��̛$t�f5�`�_�m�9�z�*,Z*�l5��f��Y
����@;eMW��ʧ�D�q�J��e,�V�	��a����3ћ3J�8�J藐��
��u��&=�F*��b[&͒*��71��*��U�ߗ��p�I�v�6n��i���ЭR6�	2ۙrfQh��{rj�i�7���'WX�v�Z������"�ҋt�ͫZw+^��WD�P��eÛ@�4�����ܑ6(Ы�R�X ��r�b�]3FÌ�9� פD�8�H��0�H$�s2��㺕"i��[��S""�a��mCE���&�#F�G<�/��Eނ�Ѕ\�5k1�S���B����;Z�	�nZ�A�c*%.$�_M��r�P�;��n�) )С6��5[AQ�T���R��Z�`��z&�2d���1]k(���Qͦއ���Z��iX�%R3E�M�!���t��1��j�ͦ��)����'Ғ��A\�/l��A��h�����]�fK��ԏV�Zč�U
n(Iw�\�ݺ���Jw�\�������Bq NK�v�)J�*m��A�4ڼe?��ӎcU`�cM�mXSHB�-�D�T)�乌bͽ�Nɉm5�������h��Fں�4k�`Rm�'lf���'��m�ǹ�K)Jp�pT��w���5�[d��n���vEv+X{�(�`�1ǂ�b�-\B�ώ3Y��Y*�f��ið�4e0��ۆIpyv�U��m�J̵�*W��]�-˄Ln��;,1��6��V�ъ���k�!�t�.�bgR�Na�sax��TB�����ۓdǮ�����ϰ�$��C��o.�B��7�*�"�e+� ��j�9���fú�݂��샕�љW�[kwo$��kQ`�h���ˎ��m+�e�U��-��F��4����J��!�t-��]�5�)� ��v�bR�����Uh@�t���6�i��їqV�3+0�^@�l�d2���MfLNb�wn�2���2��w�1՜.h�yS-;�z.	�6�bܥ�.PoV�3V�]n�Y���m3N)ZG ��SR�.�=���V��^VJ�l\Q��(Y/*�4����V�ьG��V�]�e��̧@�t�Ǩ�	yS�a8.�v0�-}��i���׳t�P��A�o�d˹yYb��`'m�
�&�'{l-����&�Ʃ �h	���H'�kQ�CuEI�U�B��7|�b5�X|+s/Y/t��I,���E�5�"�� ��7�"6��x�Vfk�݆��Ϳ�m�&��L�"j���QP=̕#�����h-dm;h�[{u�m�ޔq#�v�ѻv$�<2-�e�5;�vkp��t+B��ua�4F�r�)/j��t�wyhܗg1�Sy�*!jzU��Hqg�g�%&�CCת��+*[H[���-���i��,�a�I��E�R�9O/����cY�E�iC��Dc���ɸ+�we=�utN�£52�b�n�@� a�:2e��N+N���h���2�̷�2��?LwV�����'r�lnn!f���wg��ϖ�Rg����T���Z�s+fe�,P	("�-nl�/�mӒ��36є�i�h��Mh�+!��0�Ke�"r�	]4n�u2T�Y�%�	�-��k�VZ��#�#��{V�e1.Rݕ7�M�nTӻ([����$�,y��4+r�=ohf��T�]��Z6���F8�7(6����ao,Ә4U�m�6�d���i�ѧV�-k��T	=����y���η����,���x���tI�1i:NQ^�`�:,�c-�f^!�E����x-:T���T(�H=��&bSH1W�[�4�"_�u٢@�n�j�ϓ�**qU�Z��d�N�[�/(���~��#��R���+���xD����+Ad�n�KfK�M�����/^���fc���wW�U�wf ���ʣz�F�Ќ�`Bj���R�JbƳ�^�-�0�4�@]3��eK����pȋ�p r�D,���D�m�,���Ok,�Hۖ+R�6��qݭ�r����i�N&�97U-ő�bd�)�N#>v�]�t������R�;�1lj*v/B6�͘a6+Gk�ӷ
���mÄZ�n���ً&��i��YzE�F��KmS�踨�02�J/nŀ>86�jbϙzq���W-Y��]#L9�Д�nY5��p�n镭f��xa6aL��s\�r�w_L[�Y|/Zx��ץZ5� ��j �\c6��%��>�0�{�X�����H���[��8�[15u����i���W��GiGO&��4F��8�����H3Zl��Վ��sq(�ZT6m$�X7��:��ú*c���-q�m��J�0:���l+��ב5w�ɢw���(By�@��R�E��!�[~�����؊;����g:ʗ�r��)����hG7s��Ҫe�lC�f�8�Ym�
�w1��˩佉ݻ��"�&6&�C��x	*�Jβ1>�Ie�7�K��Sit�ms�5��)M5�V�L��Mԍ��_��Zq<�mr)=���(3���A�6�(L�w�%\v&t���e�:b�5�+���{ Ǣ${2�e�o���`'B]�졵�@9e�9���;��@osb�v�cŒ�U*�ݦ>t5@;p�g0�պC_e5FA�Ʈ�.�NC������J�y�t�1�1uºm���͇T���N�uX)�rN��:Ev]<
Nr�Qʼ%I/*L@j}��Vx�����e,���K�q�@o�Y��mp�;- :�R5�^��7vue'��|-���d#z����x�Sg`�����������YZ���[�c��xU��lj�K!�y��"�ZI�뷇PjzZ̏z���u�&����x8��=���-u���tlp��t;�5�D�-@+���h��5�Z��6;s��y�c���&/k)���	!���|g-]�B�潴Y]����2��u�`��V��m��jB*��l��u���.=8*P�].��A�gE���9��KS�L�ev1K:6�fb��5��y�KOE����S��+'m-]ǆ�d�*<ʖ�='uNy[|+�qk������^��E,�m�مu�,�{oR{���ܵƶ�o0�5d�n�y#�P��;>����K-��Fa����Rj�Uԯ���=Q�t����I�9RA�w�K*s��M>�n��N���"�ղu�(1�|�̝�Wc���-}ܠ�*�$�|�h5����+q,�Nf�:_cѵ�%Cu2�hs�l��i�������)V#2�9����&�8�L���R�+&�?��4�^��X��5$�N�yD��1fo<O>w�[�\#�(3^rW����O�NnR�-s+ ��Y��	uKwn�����;33�b3`R�W�w7���k��<]���$��#u������}��{�ȥ[�v\w�����΍X�f�lEi9YC�dK�ձ�	Bj����1p��xv� 2�T^ڔ1N�5GK�cͻG�NƮ�9PL�%MhU��⾸�yq��A$r�.ƲS�#r�E�����eY.��Т_7��ܐoBq�4�.)Y�5��˾�ؑ��!���L�ե[�U����WP�9Ý�C���p�,��L�v�nK��ʤ*��w9Q�r_(0q�l@�D�Y8�ʹ
����K�S�_!n�v/�Cm���i�������u�e��E���u}5���*��t:m]�u��d�뗼�n���*P9�_*�j�,�&���\�ttL��s�2���J�^��)��$A�Rۂ�iQ:U���������z����8�TwsX×N̻�$h�Z;^��)��١݆�N=Z�s�ݱ��]mqG{�ҫ�еW��ڻ1:o��I`ѽ�i{p�i����%m\����i�oT�;��0��L��J__�z�һ��Y\\̪�WK�gwtJ^qĻ�)�r�Y��uCP���ٷ�=ݰ���%�|��S�켒��S��S�w�zwn���Nz�xL���Қ�!8�m�����,�q�ke���@8�LQ���E)�wX;�v���|)��k~6�z�4T�����nK)�4m6jA�y7��bڛ���i��էs��wàDc�4���渚e�&j$��\)��vM���%ݎ���b����7�-�����i��B{��������zf-�⸭J[��55�z3i���Y;��A�o��[f�#R��VJ�Q�7�n� \}���������bӦN��p������Vl���:$o<�v�����>V�] �����V�A|UK�/a��,܊�T��ށB(��+��;���ज�U��;��Y��s�GD�R�0�E�؇�]�ti�7J�_
gټ�|��}7Rp�Ns2�P���ٰ-�˱��P���N�08W��x�r�Ȟ�� �0ĒT�J�YD��\1��X�=.��r���X�S$h����"��V��;Y�ʓ0n�����;��`|U���8r�B��v���d�hG���*��j��Ӈo-��\��9ͽ���0�/���ŧ���|��� �.[q#����$=/����0�F.6��8�'��29C���Veu��S�G�ZF�v3����ݛ�UwZ���c�{)]�e�,p-*U�<w��(Q/�_=���MX��}pM�xe6&���Ҡo�Y�f���*
�sx�2�hҔ�w�����c�:�6����Y}��`���gNԛ՜m�)镽��Dv������P<��ٚ'D�4^9 �2���6���g#،z9L�d�8j��_T%��B�>-N�k�ck>S����W2��vkkvmܤ#���c�3��� E�W��V��άΙґs���Y��u��vz=i� �^C��S4l�nG:�\µG�|�.��2_6�N)$�%E��'Pp�ͨV94����=5��Pm2�z�_�?>w��Y3ihGD�ڛ�A{˹mK����e����9��S<OSc)7S#=����R��:M�p4%�VÜ%g^��X���|����eM&��WS��x��f�̌�x������>#/q���ܴ><ʚ�f.Y*R�jҮ�쨔�N��g;���\z�T�mӋ���G���rV�bLf��>\yo8��]Bj6�X{Xkk�8�R�"��N��XM�&M��{ܱ�8���	�":8����[�/8��i!t��k�Z/*�	�=yY�X9"�;O'}1�J.��w���.�u��G�,�T9ԫ"�:�T�_P{N���]#�G�nK5����1�m�ʲ'8>SK!uyf�^�#�0w#j::�x^��i��8C��&΋y3q�"P�mM5	�c3��V��}��Ht�Gp��n�=Sp��B�l���N��u3ۆ��5��E�Z2k��sq��5��1K<ސ�u���5�s9񅱉���8�i+�o�����2PW�D)�j��kD�kv�w �yȥ@�i5�ca���r�8lWMΥ���z:�\v�ٲ���-5�o,��6(����!Lީ���I�_��R�y��j��dz�m
���9�eN6'twc�Z:��(c7�N�>�uQ��M�!y�!2`ʽ��0hɰ;"�'M٘!NZgB9���7�a۫u|?y��|�o��N��ZU*K�䠃f-��q�B�"��eJ��y�cG�\۲���#�X�ь�!�wh�$�W��y�/u����M.��&S������6�����K�UC�i=�s�8�;
Z�w����θ���J�y�ĎF�[�Ӭ�����+^�.�t]�rg��D���V���CD�-fv!�^s��}RI���t�Ӷ-r��I�J��C�N�R��B
R.��pY�e��d-�X��\f�h����{a��vo�/��ǒ��4�tF�U��IX#���ΥA���Լ�	,�[Z�Z�aZe-��$
�ujv��ӥ�#~s�O�J�3��\-vb�����3Vk�,N޷�Pw��Р0�Zl���m��[�.e7H�u�]N���[�_J7@gi�uf�+vb'��=��]$T��p����Lk��Ҽj��{K��O+A������Vr�`=lY9��0vM�����!��{�iR��L�/o�[���]	���+���r� b����:U	Rr���t�4����Ba��ܕl풬f���b�y�s�L�a�E���ȓ�=,)j,:�rDu+�n�6����Ґ�n��Lm��B��_\*�Ұ��m�U�h�2�0ɶ�KN����S�b��ܠ��i��&�_#zvlmK46���D�n��O!������T(����G*ҝ.3�&;{<ۆP�I��b[te�ab��Ε��l�1�O���K��\����R�Ū:m�F빖QМ�8�
���@kl��_"���;�7�K�������Nf��������޷���B�)� (����� }j	VCE�(��nл�|�&�+��If[U�9�#��;�.N�l4�����d#k$����i�Y9u
Y�V�=e��C�qM;Ry�"��)�z�(9�[겾�Z$�E�T>��s�3s%�rL[X���oo�����<4�o$��lN�]:�u�6�k���6��q�pSB��s(:���F�Q���9JLYN�`Y�ht�F'��P�P@��tܐs+�Y�&t���t�:N�N��R�]���[62��e�&��:�2��.����
n�u0��&�V�f�q�mh��m�p�R���Q�P�(��ޅ�j�U�+o��]���������aj�a�=���,�YnFv�Xl(�"��δަ�e�U�������H��Ov'��W�+Zr��+�U�I9M��oNK��']�wqM��&�owmK��V��m�
����p��������H�8k�Z�;FWc�m
v��8���kQzV�(�&Zp�o]��.��T[�5/�ȶK�ZŃ��W=�ѵ���4Q�\�����Y�]/%�S�w4�;,�# Z΋�s��,Lsͤ��M��<�`V��o�W$�_���qזŲ};�CD����sc���a��&��Z�&]��<��b�W�H|s�q���(��B�nCd��y{I��Δu\:n�M+�ڊ��ZV@�����J�ع� �"h(�ï7H�-��`�����j�ÀQ����&r��W�zr����N3h�Z����B���<R�D32;�l)h>��3z�"�7f��R򐐸���\V���(o9��Z��IH��r��ner����e�}��X�w��MD�F�׹���%Jq�s�n��n�b����Y�-�S�{D|�!+�U�Q����u�ב]� �d�Bv��԰<t*'0G��1C�S�ӣ�Ź���\�r�՛TPҧ���u� �
]����b[��u�捵)5ƽ�(�S��Ku�*X%XV����c�"[�p�<.�Ô���:�q��";���YF��_7&F�8�V�|�j���'�U�cA}��M���'k+L/H#IșxiƖ@󙢑�2Z�h�)���
�u'�#h]#����LA��-�2���f���|�������ۣ#��V�Wrae�;K5.�\YdWH^_*��W	%���駵H9���9I�]�P[�umX����Ls"\�����E8�7J�9fԉh$���WV<D�ov�ل)��x��q�=yi��N�Q2�\F�9H�V�W§H�� 7����)�%&��m�젵�i�8�PΗ&bJ���K +��,�'b��v�P�D[-͝�[U0�N���w�Rg�"�����eC�;��|�S98�vܔ�te�opGy̎��s�4�6wVM�gm�!�zq���ܷ}�KWas��7q�����x_f�oz����6�=�����=����2�1�t����gc���s�ɝ����W.�/U�I���\�3]T����GU[�V��b�����O��n�a�R�m��oj���>�t�%�W�rJ�:��m6mӼ����m��]<;:�S͹8o!7���+�u�j�r���t4t�vG8ՉOsv�8���94������t��R�!v�+tQ�v�=u(v�k��A�J�IJۋr��Tw�Ï��kF[]�c��Z���c��f�7m�+��+5�pI5,Tr��Bo+��JHRd�b CD�3��ѵv�Λ&.bڤO>�A��5UvESʵxG#./T��&4b'K�z����J�3g�������'bjǜ-�����{�O峅L\~Ȼ����0M�w3\���PvP�<ԨN�G��R�[�Ʀ, ٝ�,��Ӽ�В��NB0γ����7���K�R#g^������L��i��g�}z,��Ԗݦ^ͧWJsx�R��w��<ӎk�Gn�B][�t����bn�K��Ǭr�������I�I˽=@4��ׇ֚����XW�f ;���q�ٓa�-Zs�u�R�\0s�֒��p�@�en�яn=�{`�qj}�Ԣ&�᧥k�燔]wM@�!9�&9��,�q�OFs�x������҂��S7[��������>�k�I�8��z�����%��pe�R���ߺ���N����<���ϲr�zJQ��l�,��h�k^�pMjB:�pG��Ȣ���c��-�,
v�y�gFWE��c@D�A]amU xmnbطbB|�]��M�c��t�Ҷ��]�����ކvQu}�6��{�j�Q�av�:V�T���;Xq�ۂ���bً��1�ۉ�/z����,�C��R�aP��׼��Ӫu܈�[X��q5Vy��\�7{>�Kx+{�#6�Q抗!�Kv:��]M��
a=X�#.m)�ea���N<��ߟh�7���9wU�.���< ���S�/���`e3��q�����U�b�-�ۜ�/���k�Nܭj墵�W�[;P���Nn�8(ʹz�����Y��n���*�����\���+�ڈ���q��'&��[F����Ė��띩�b�e����i	��Q��w>񱝵"j#]�`���Oz����2��n������ܫ	%��RX�t䂺�>�1V���E��A�Ԭ����}�@;�p�\���M�1�a�۸��[z��	Յ+M_Jɭ�,d��"]J�)�w2Ff��d��[eG���R}R����(�T^���uJ�l��ֺ������* 7�7�F.<�;]2�l��\�|��e��;�H���&�g=��D[�(�}��.��C�h}#�{��v�L��:mqn宮���~����^�|��6������y����]����Y�eP[�^�	��� f�8��1��`�e�X��bE��E͙)4^RWZE(&1��:(q����n�r�c��k�h�Щ
sk��B�e%��J��ݍ��O[`tt#T�,�
�bv�-�Q���Q���/�Am�޸B �JA�٫�⸍�{kmY\�ˇANgV�^�� �rK4���7eѕ�m�����"�t��G+���)�/F@���Z��A�ڃ�Ժ�[��y��(ܛ��X�钐U�VA%���뙽�]fF�9\� ڐ���SSy�0�;@s�0��M���Y{p�7��I��7���Nu�Q��=�fN�Gʰ�����}�0��r7�5�4\������V��n4��=����U�7�(}���-s����9wо�AG�+8�F����y�O-�J���8��R�;��0�T".v�$p��¥;zI�9�8�K��ʳo��;�+l]$�B��\J�J��Kk����4$��yPwV8�5"�:��9��9g/qi��F&l��֕iFE��É��f���vᦨECx3���/:�c8������Il�LLwU�r`�Zf��qʴ���t�Lפ�nwo�3e5��u�;H�Y}�3���I@	2�Ou�*�JWgWQC��+7
���s���Ѽ�oK�5��,�6���v��f}�d���<d�cl	�/���Z�t�ҁ�:�G��r���[��a:�k�D\�5�G6���Ѯ��ȕ�5�<��i�r��vұ�F���)�C٧૘"��{�gJ|e���c{*@�h�L�C�ѡ{���/��Cxi��V
a���K�ʩ��v�۬��Z\�l��ѵ: 3��g&j���H�$�݋I.ݧ֭U��R����%gFs��<�WL�zQ͙��iH3�m��LWc�Wh�'�Jw͜|��uҖxJ	���^�9+��v蹸�^���N�9��s��۷7�_b�y$uݜ[`[������܉	$��5�H�9]�����2�YC*�5[ut��}�\�@����-��;���/������љX�7�Gf&*P�Mu8��j��UN��x+�l���g-�Ks�QN�\���2D�c�����5���BA���ֱ/-moup���㱸8r��6�7B��z��Y�.�����h�i&Ym�ض�n���x��3��3O��K|���B��(��j��3w3o2�gwT�k �z�r��Bڭv7��!z�d���^b��y�Cl��0�ΣQ.������Q�2�(w��{6��cQ�31��/yN�M����P!��guLʶ�w
�6mۼ���j��p�|6-:Dl�%�	7��rH��t�9\V���J儇�r*��Qv��"̤]��K�ن�b����f@s/]�ɑ��Τ��lwMS��:Q��	���
WzJ��4���6����[��4�+[��%m�K�I���	��F��f��z���Q��t�.e��k#FY�.�c����\��{Iݙ�d�T��]�[nM���ʝ�h�F�
�#)]Y�b��9��u#�+���vpՀ�� l�E侴�F�KVu�:\+f0+���}*�h�L"�,ge�{X�Y�4
�)u`V)��mz�7z��f:�W��C@p��
z����,S6\6��D@S�[5�W-����YJ�nG���{!̋��т�n��kt�:�zQ��f�ۥ@cֆ��ZiJѕ�9Q$\r��b��p������\�{�f�l�N�K�oh�df&�[d���ٵ�/wA^^��J듎#1 �P��[��9����=qWt�:f3���-m�M�h	C���̕j���x[���;�T��Rmv��z����ee��\���ȗ2�o]�<����嫑LU9�Ȯ���R��p_xu�(؋�s��oM�(�NNgUԅѥ�s�t�X��F)tr*Zn]i�)���u�M����(�5v�l��Mm��k�]{z1�"�x}gh�z��Hi̦��rܽ��5�Iog�#N7����c$�+)��V�]���h��Rܹ�����];4T�*S	�M�f^;��0�Bp����t�:4suGu�9ZZ�[£���w͡�$J�շL8�v��Q�	 0{al�"�܁b�Z�$5�0_`y�խ[[�i��]4825�:#��ɛW��Q�\i��EYB �О�gעb��x��l���]ͦ��&�q�N4�*nW�2[5�E��oa���]��"'�I�v[�O�l�W:e���k��r���jH��6ݐUқV l�fٷ��i�A�� vc�N[WW{��Z���ة�0�X���I���˖��(;��5�yX����@<�oA��M�W�V��aj�����jW�m:d��n9W�ud�;�#m�MM@������:ڋ���	��/r:*]Z��c2õ��E/�.�0]װG/ŷj^���r�"���)���mU�M�̔Yn�+ R���m��ۚ«�G���Ճ J�$z����o{�S�T=]B������Lb�rAm�0oU�
u�D�ғ˵�F��h�[� �X��,{�����Z��V����A��vf���n&���|,����0��bC5}�	�k����������z* .7"-�"�bsJV���tt'E�7[I=�!nƃR��x�B�4^;Z���3��ֲ�\�E%n��D7�S�_��zctL�EH���㒅��St���YR��IG��@�g��-9|uo�[F�-��V]poa��+p��t�%�r���h����J�v��u�����k��z�����F6���+"v_:_M��$��j��77��#�fBm��&��fv�������G�坭e1�fVӮhK��:�]��N�ػ���
tU���X1Ӛ��r���qL�Ύ�n��s���M�mU��!�#l�T�+rR�]�Ff�V� �ri�)�A",�o9-E��ݾS]��qa�쎗��l2qB����j���}cT쭷kg%��v�c�k
���C�����Z����̮��k�;\=q_\����6[�|��΍�iL3��2����[�;�Z���:��L�#��=�o.�^s;͔$���P�Eo�7Q��$Zn�����k`l�ѽ/e�N�h�Ļ��E��&�[n��9�5x��/�����8��������$Pѽj�Ĭ�WֱD&72�(/.�9�e7lh�s�nM�f�.�u�!!�;u4�JJ���c��S����Æk<иn-���y���}�c���x3�5�.�vn�CDܷ	��%
ǨP��g	��-P��1�(/�x���o38x>�w�Jo�����`0g:B��pM���ݴ���R\�V�̑}ov�@X�;f��T2���ݹ�ý����i��EcZ�|.�쨋�:㪺�t�N��s����7]�Be�V�����)�a�[�`�p�sS;�L��y��4�aQG����/���e��ĎN��:���� ��v�3�,e�TK�K<`L�7�Ʋ=b�KP���(<z��.�es �'����e��7"�uٜdʶ�Z����\յ�6+{4p����ظ�|B��N��<�`��k�.��ѣKd:j�]�}�v��:P8��)�oh�ܾm��DӝYA�[S�]��Le:��؛&q=�z�}�e���p�«��i ���I)s�b�]��,yQ�B(�@V�I:���;Y@�O4��Z�']=��9��F'l�1Ne\��~�IW�lR�%��%G��4T+�/f%����󓢍o0Y�oۯ�ݣ[��]�)�գ��iE�0r��f����g('�)��`؝%���>Y+$��Hk^�R�l�r��ay)��m���u��}�Z	���Ѣ��i�ZaNV�|�UE���1#�Z3�7%'� �C'���F�&#�f/�G&�_F�Sl�S�-�S��B�H�.:�۬]�R+�X,c�za���s�!
Fا��G�����N�3m���qm�5Ĥ���:d�Q�7�L��gT��d P4�6;8&X�@}�]^���g���N��� ��;�k�]�E&�{ql�Imݳ��x���>\bx��*H5e�b�ݛS�o�˖���;�ѧ�H�7CW0����Ӄ����`^�v|�	�D:�� �����r��W+x&}��Z�;;V�\�ɫ���l���7�y�(�C�W,'hљ��Wn�ҏ�E��y�Fn�e�j�u')k��& vp��pʂ��ub�	z/Zv�"����M����7����wx���5D..�^M4�!s"kmkʵ۵ʤQdqgS�[ֻ�\���OLiI6�8�8vӑ�``/�U��]��:/b9���ۧ�o�o5�%��d�
t�d��0�� ���m���6JI�7�w+yoܢ��$���b��Z�%��,�B�х���n*���M��}8\<���ٽ�<i��-u	o]��kPw�g-�;2�V8��3WΌB����@��5m�.�q[�R>���}�{���s=tځ<��N�Ń70������w�w@N�RJ\�PQ�ћM��ۣ���b%n����Sjo&*E|��n�v�Ǉ�=+났�Q�>y�����.�Ƶ�
�l#❉���Wo�dח�B�����ړl]H���J�j��u�LB<�[mt�v��iv3��#SKj#���o��R����.vFw%q��ૄl[��Z�M��i�{n�кdg^�u��{�Ogi���]�\�ݕ4�R���2:^�WLW�lJ͉!v�%�=��(DՄ�2Ր6�L�MX�f7N��z�i�3ZM��⊧�Z���DhUwj��V�@wZ��\�ظ��r�փ4��޳FqQ!T�[���kUΝ�O�QVjT*���%��k���RN�����T��Y�W&+�Z�7[,k�Hkh��S*œV� �w،�t1��M�ǝ}A�
�z����ۓ4�])��؀��Ӥ6/����:���+?v6T�C��vA���5�B�z)Ք�}[��ѫ�0O]h��n�:k���.q��u��jc}��̬�����|��Y�*K8 �H]:��X�x�
r�]�~��iܥ��a�a|����Sf�����A�Ҽ��p9ʲ�7����N�wm���fE�m�Dఈr�-!̗S�;��]S~�kX�`�kTS��*���B���ݚ�@f8�}�[�6ec�ci:�Z��}g�)�=(�	�����7�+���$�(E+`'/s�,l��yJպ0뷁mu�//���9ʬ����W"j��σY��6��S�ގ��!]>����G�� �c봞�BG�gm'\p�8fe�l
���ݼ����m��}J���{l�s�S,��n ���*⭌�Il���=�:������S	�{Ř���u�tRĪ���f<��\Y�NѼ�a�%�V����ng����vk!�q>0���!-��5�f�ǳ���e؜�,�PV�Z�-�ꏱ	���Qhr��m��~�X���i@ꡏ+1>;���QѣfM�;\Ў�BM��ݣ���c���N�T���[Bf�Y��_n#���$����	��z�qA��ݨ���,�g����F�S��}���Z��j�T�������6R!��n��΄@𴚊���'j�1�Wu�ApLo�@���l톯k�b5�c��V��L��U�7C>��'L��=�9��+f��o�����&�H��\��H(΋j������ �׳$�Z�5WS-t���i�F����؁X(qgt�{V��K��;*nP#��5���7x�� <6����KӤZ4� .'ŖlV���r��X,w,6�m8�N��.m�V��v����
H�]��ۡ��gwz��6�&�
�V��:�fmլ��Ν��@V�DE(^B����yJl����q ��U��c��F�����1nP�%�%���4^�i�6����n��~�]��(nWg�OS��ŋ��c��Wy�+�q�����9|�J�݉���B�i��|�p��˸t�5�Vy���Dm����Э=ى;��kWF\i�/o4�я�
���P��u��u���];Q9ԩ�����W�RtWt�/iQA-��ծ)Y��'�W&6@фx*�4�� ���u�(�sq�Z��:��Հr�ʽ�(E���A������;vq<x�W=p�Nk:�L��i�p�S -�j�,�4O�];/J�f��-;�^�D!ϭ���~-uͅ��b���ø�8�g8�A=*�|r,�&g����!�(�tk0Og#`�9�I�5u��u�{�s�R=�q�E��b���3f�Jun�g8�'♳W0t�3�}u�aqÏ�e-�Ң�2p�V���uA�V+-`/� ���e��ui�-��.�h"�cR�J�J��g�D�94(Q�T��nܭΙP��R<��U���e�GTn��9�i��mnj��C�7����c��n[���_^�*Z�&�n�vJ��<Ŭ-e�V9+\	Q�k��Hprh���K�W�������>x�0�Έ���Z��|	G/+*�e�K��u�D��+ȃwk�l�\w�H@�ݴ��"���h���q�-ڷ����=��&�u��M8�}l`�V�,�6��9'^�*�9ʜ�7�GA�1@肁{��!��R�q�.�c�	�wϵFM�#�1�}�V	����7��z�L���v�J�IO��v��T�	5�j7�u*Ľ��S��e'f�a����-�s���:�xbe��R�]*$2�E ����4�c9Y���p�16h��J���z�Ts�m�Z�j��l�zf�X���~�W��>��������_:�qg�\9��+�ݔuǷ�*S����r�bŴ�N�o��5-n���������l�*�Nl���;ΝPɣ(EqwP���,Y�0kɨJ���g�����V��Bʹ��oSyj�T���f(J]uύu5h�e[l���_GZ�`���r}�*���;n�z֛䤣u#���Ҡ7����ۘ���ը�Ӏ!z�s{������y �`�m��cj%��!�$"\~P�{���l�4׺����;�`3�R�Nh�s�a��;�^r��3H8��l����mkz�{4bs�v�v7��/��,D�_	��L*nӠ���w��b��̹I>�M����9�Պ����t��t�p%�s5$��[�+~J�[J��ȴ�\;�9��E��3�z�/w��N=�@�f:U�+�w�lV����Q��7WZ$���N4���Sx͝jA��l7��5�4s��VN%y/�7$�#aJ��v�[:��Y��n�إuŽ}�c}��8pn�7��>��̦�Wb��p${��$K��o6r�<����-oc�[�:m6I�4 A�s������t�����x�fي�z���[�J�[����=z��ȕ,��=aؖ���bv�|�<�6C��( 1�����&ě*d��tg�z�U��е�>�^[���-�L�'\�E[d'��Fm��Y��Ƃ�}���������]@�\�ET�W�%r<'psÜ�wB��
J�#J�St��\���c��T�u�q���*G-wU=J�(�9AUQ��ۑ�s�HJ�u*�qܜ����L=��C���E�Ou�D)Z��atK�Xy�d\�1�u��p�r#Ѧ�<��,�U%�N�QRN圼R���f4��JJ�S�{��Wp]k�۝7w�I�F@������A�B��;��:�.y�#ԹT9��d��M�rIXEթ���x�9�t+R�qʼ��=)���Ө���i��HHjɥPp����Q���p��q�K4�%��+��u�S0�BDB�\r<wZ��T���]�$�螖��ԣT�K1H����T1Q�y+J̈""u9=3�˔��P��PCK�
��a°��]ww9��=�V�*�"[:s]r��uBȬ$+�^���
�.h�GX|׮�y���������n����w|zf7`��+k(u�:�V��/m��Ƿ��$n�vT/5�+�N�X���]4�����Wزq�]hi~K�_�J���l*C�V�������wL���k��֎�>{1��U���<��2��r��~�_��k�05��{�p�eB�<�SO�w
At�dɞңy�M��m��b����5�\�ׇ_�1}+~o��x�n�!4yx#�^�t�c���̛��zy��3�l$�vjw\��5Ńf�҉��9���tV�f��с��vo7gV�b���'-m /R�aD�W6��T���I}^�5���h��ԥ/�Oj���|����S�S����xQ���|�6'�y�ȗM��;��M�����r�q)��Yg�>�%�F�tV}UgI����'Ey������6<"�7$S���S�Y��R��ĸw6��aj�����GI:H�W�U}�f�:����\�Og���Z�i`�0�-���١.�Tr0�t���Y[iA���2 ��J=���g��i�;���+2Bx��Y�� �/zde�RY|r h�6���[��^`�P�����=�Pɤ�/�%���V�L6[?��rӽ���N���kp���qWN��Z���٥G��L�9JQ!Ж7o��Kq��O���!���[���gU�΢Hx�宼OV�W�#j�OP�L���]��t�Х:Q��Ii���Y�7��v�Z��ۥ$���S�T��n��r��Z�#�CRt��%����!h�(�AyT;���+��¶v����s�ct�PN�����bs�C���/J�7]��7tx�2�j��G�
W��m_L���"�렸�UJy�(V�]r��e��Z��&-���\���T��5�P7xb����.�"Dc#���4�r����>�����:ފ�M��H-�{͑cn�F���v�٦ �a�L�o�ԯ�'�����Fx�;U��1wS�.�h�w<��'k��>�"��)�&�t{(y��\��*��CɜPS��cͮ����l؎�T����+��ӗ�=Gô��ˇ����s�&�ˀvӽ��ٽ.��%���gl_��,���?.�]
4c0���Ӥ��A��A��>������?^*��u�# ��y�����i'k	V�3�s)0�������Z U�b�)s��5O��G9��^��;�R�3^;;*=\��ߛ��u����]�z/�����%<O`U 
�K"�]�^� �%��`?*�MJ�S�n��E���������O06����D`�o%���tmv�P�J]��z�ڀ��}�r�ۏ,)�E�`����kz�vWe���t�l�f�� ��E�6�g%iwQz�����b��O�,1�Z��J.�]`"'�\Cn�E��W�Μ�E��.��YZ뗒�_*�CQ��Y�=j_7���zk`�$�=��Ż��nxVm�޺��Y�����h�Z%���*N����T������:��]���|1�������n��SơQ���є���`f(�i��ս�!3���;�*r-LP4��[���0ڄ���*����=㐕웙�2̪�I�t���s���D������R����1��N�,p8{"����OHٍ*j���j���|�7^�?�I�y��W�1>��t�83r����r���y��O5|��A�z��f%T�G10"S��Z]��iQ���oݺ�Z�F?v��/t��h�C������K��&D�[�4����M�z;BM�^T���f��t�3�\��T'���71��3��
\F%�\�#�����i�����3��o�՝Ѫ�ƅ�*1J�}ʈv��*EK�޲K�JY��:�T�O����g��d3�j��c�����J���A�7jsS��v+��f��aJa�$�"hg�j:ked7_[�-��&6�h�򬧼XA��tM~�-W���f����
��Gm�\�9]��}ig÷��gβ��vC��2vYʚ�"�F������l��#6�$�>�����}2۟OU�h�U`�_V*�_u��\rwr. &C�l�	֦"r�5�x���i��=��x�஽6��~ϯ�#u҄>Ϸ��&�U1��f��EY�Uq�c����FF�Z�C�.��8Aq�/�2�Z�^�A8W����b�!�b�&�e����)*�s��*B9��\?np��Lu��p�f~����+*��EL��E@ֹ�tn^���K(�1)�\2��,�F1��m?�׹f�Utةj��A �r��s=�ct���>�n����*�S�e4*���
�CҨ�5�{װ�֛MDb;�F4�6����ݼ�j�#�(N�L�����3A����(V�Ǽ6y��t&ފ��'-r�R����-��ˏ��Q|~����p[K��EB�V��,����a�{$<�7nE�Wʖ�g<�ϖ�Q(�G@����Q=ƽwj|Z����OW��=�y|�㳔�|Ɗ��-�tCӏ���]���� 7��`
�U�q�^���ޛ^��Z�W�J������(ӽn��G�T���.�Z��i���Pm�]�/���^��W2"jF���to+a�f�O*ܶ�����+y�k�u<����ϕ���5����`��ur(�ɼu>�n��r�u 7�A�_2)N�b!]�G+�n�l��5v8dk�$U`���5�������n���V��B�D������ђ�h��YMZ�픗o�l}��c�����f0�H��f0EBn��׮�P��w�����=�vڥ5b��lr!�K���/�C���]l!��,�#*�:�&�q;Uyю��	��o
�T���r���D�
L��'>Τ�D0��?4���(Ue	I�}�_JW���|�����i����ʊ�պdC;yp�Tw<�2U�~aV*kqr�~z�E<[�{�p3>Lm�}g૗���?M,�-��;X��S�������-�ilO�;nZ���qϮ���� ��F�B{v8;��F�E�Q'�_M���D�t�J+�V7�b�x�.5�f���L<1p���V�;�*�tf�"����A���þ����]�O�V�q*��'B'/��`W׭d1��\E�Sh�%V7��F/s*t�\s��.��j��iؗn� �pf���fp�EK���|�>w�*R<��}�r��u+N�Evuu���[|�%�fTn�=����-�F�4Dnu=��(���h�l�{��pޏ��7��Yi�V3�1eԫ�T�ɧDN\׫��.��v%�o%q!����\p�"��@��G&ъ�S:n�!Ԍ�4W4B�nm徃�.�Æ� �C|�N���	��_X_�Abx�j���A���#��7=�����q�O]�O.k����as���:�U�$�#�.���H׸�%�bWp��T��p�v��v�df�fx������&aC�Lv|�/��l��tu�P=Υ�J�E���gB����Q�
�%�ZhM&���jK/�|4Co��3l�
* :	@^�r�IF]�/+�KNv������UM�v��r�ֻH�NQ���Q��b��ƛt�F�ɔ0����gzyM;��@� ƲE|K}9�:P��놌t����C��m*����ts�=x1�w��]�w�͘e�	�`򞣔cC�鄺5\��j�e�&�{�&�_�)Z���Y��j˶u��t<k��OD/���o�gw�x:��下�)�y��HWTG��ޞ)jy���~ p�����_+�U<F�bGe8���DK�.�	��ck�H����_֚�"�Jd�m�����K�$�\e�*�V��=�$ڊ�8�2]�Ys���` ��>2�ՁWb�Ĳ� M�֚��=,&v �j�A=xUޗ��ohөel��A�TW}��\^�ٓ�@�ЩP9�7�nJ^�� h"��k0mj�Ē��('6h�.1����+Qb��Mtod%�lۛ&��Bi��.���ヴ�u�������k��5��;i�ٸ�/�� r�VQ̢t��npW+YYSU	?�L0�,63��ZL_ٲ���l0Խ��N��~���XЭ��Ֆ�G$��3{3���ݿ���a�qSLp�δ ��P��R�j^��Y5�®��
yۉw�R^G�f�V����A�r�;�UL.����U��I)�{(*���l�O��\Up��Μt���m��ͮ�Vµ�u�=�"�<:�2V˙⾊�h�<�"�cPvJ������,�L
��+\[��W��|� y���w��K�xy��O�b��ɬZK#��M�&+��?tb����a�NS+��������� �q��8#�s�e�ֶ/�`؍�c+n��ȵ1@��l}q��1��D&�aU���b帍���~â�p�M��|����K��]�K�K8HRX����F1��=}W�B���j�
6s����j�`�|]�yQU(*2=$��?�<��r�8NhN��aOM�Y�u9�;n�E��4*e�]ez�5|���
�.:.�a�V��(P	���o^:� D���� ܁6U;g�0�}S����zИ
{;w@��2�$2!3�xV扙�t�k�D{�����
�XZ�x��B�hru!x��i>��4yTH��}�*�o�V��'��{;o*[��L�k'�ngD6r!��&�.hAD��}2�K�&�#�`�&0�y��\�|7)&���o�p'����b��rR1�p�q��*�)M"E+�:h��7�oZE��Φ�/*�}W�HXχa�����Έw�1P�vd�Bs��
�"��vd��^u�A
:����Q*��=ftł˳]�ouW�$�0�f��`&��kW�5���kS1�Ѵ�^'X�^�t��Qf�
���,M�U1�-R���C����Z��|�U��u�B�VN?���������L��}����5"wwU+��$��L��m:b9�������CB��������/��%��dk��Qq�ڴ�5�ޞ�(��Qj��ƮJ��Y;c�m_�p�o��`�� ��z�c�h�Dv8w�ܻk����5�NYGW����)�a��C2�q�����b��:c���v�Eat7lE�(��;�3G��݆OV�̠�j	F�oY�Z�'se��u;��6��v�gct:t.^�]�D���};1a�&V�Ҝ<� �v��ӝ�)b�� �8蕹���4+�2�PŹ/<�ɧ���d���'�?�m6�6��V+�����T>T҂��0��d4�k��z�ܦ{����Lh�e�W�eRfGY��*Q�� F���3Ԅ��w�4�+Wbn�c�0�3�j##��&^ܦx�M�$u�����uQ��2��I�W�h{�Fʐ�v]ĳqEi���Q�n�1��j^�O�����cn�N>�3����D��D �O�`
�UHWqۿ��չ.�j��]w�cQ����>�=�zo�C�a���ܑVݑ��ћS ���#OT�J��F�f�ﵻ�Yku�n�/��o�W�T�l�q��M��wlȵ2Q#{��M��N�E��N�,����"~��愣^�������	�VY�c%Xu�1I�#��Fi璷7o�q(���3X]�����-�Ɠ�9�����y��R�eD��nj�V�s��s*@�b�q��)����c�it�{k0t/C)�]t�}�5!#@�ݰ��{Ǥ�/�����K�
hm�g�œ� ���W����x���^�q �>!��tɯ���e:u�*{�ڗ���h���L��x�����Ol#�����=��4g�w�wyb��VI����"S[Q�vJ���_��8�	9�u�*�U��M��V6�L تЕ�{��M��RwQ��1c�����o�Hڝ��c�[��Nw��� ����f�{v8;��F�7,u�2~[[T�CYOz�
����Z�|-Ҧ�㑽)��u�F�i8�es����њj8W��	槷'{�c鑲�V.�9�����$�d�l�:/Z�c>�RꮌW���I}X�Ȭ�^�:������X��*�De���h��L��@1p0 &/��E��O>�g����#X �M�纟������o6#��ǉJ��b~'D*��<j�P	`��X��ѷ����1����j��;�xkyl��*.���u�6�֒t�G�]U�I�Ɔ� �뚗�8xȓ5Yݝo� �F8SӃD0��Bf���7Z9�d����N��`>�I*���H�y=˼��8���O�%Lj�<�=<Ԗ_�����\!p�m���(҂W�'�]JUl^�@p΃_��눮�l�;u��9c�k]�Z',�>YW��<�ĳ������ֻz��l�j�d�I s�҄(�놇-Wɜ҆�u�H�#�W{*7v5|;.���݃�C�z�KOq-Ǘ\!�q�E�N�PdV�؃:��Ʈ�=�;wF��,6�}�U��a�vb}auEօ_q�]^�/�j�5Nr���Y��Ӥ�{U�����	�[·tvJ�o���>Fb�g��w˜6&��
�{�)��w��L�"w���݃�X.WPƝ�CO7�p�C0[;5�ڂ(��]��w[����f��a�F�ˣaEԢ��t8��!����_4e�/�X T�h�6��6��Ƈ<r�^�ONr�ic�Jf�@��Qv�L���mp*�.W4��:�f�/u�g�����9���v���ԫZ'U���]��<mY��n�-`�h�B0�ޭ����p�K�q�n e�R��oj+ s�.n��t��Ķ�"��y#b�i��A�͙�+)��]��Rv�v��̦(�!���
��:ܗW&��+mV֧8���Y����yC& ۔F-Tv�K�dXvͭo9w�oḚK	�xz�a�6	MSlѦ�y� �2X�����%�B�+w*<������$��f�����S�!'e]��h��r�\�[$X���I}���m�*�=0١ӴeѬ����Q>oa�����e�@��]ǅ��ΒY{�df"vU�o�v힕�e�W�P�qƁ��V�Π"����Z����x#�t�,ݩ�Q�?�d�cb�yǀ/�G7l�����9��L������AceZZoT�Q' ��];XH�t�| �`�'Q
(7�í�؉ۍKZ��|���f�^��̡��dP9�˪Iε)����S=��V�� ���w���lᲴeΨ��1)�س���s����S�DXX��jv_wc����]LέF3�Pv��4��Z��t�)�ѩG�:+�۷��8Zf�V�Y�:R�2/������\��׶�wN�]E&,]�j$89�7R
V4MkdM����
�DuLGS�R��ĸ�q�כ�S����7xW�T��G͈ZV�b:��mub<3�p{�[j��h �1ee�j]M�tʸ�y�Oʧ!;Rn�=��laҕe`
n>Ҫ#�p�Q�;�������� ��@{���-�.�zȏr��g'n���v�ؖWgeI�j��l$�P�]m�:�gQ�0�,�ckx�ޫ�y��ӏK�lf�I�֪�Sz�N�NTܾ��as��|`\�T�8��b�۵%������-Vq�;s��<�9�صt��B�1���Yǲ������!���j� ��nW;i���5h�}���j*�.O���lґxs2�RГ�M����xs6�r)s�.�x�;6M�v�pH�Ĳ��՗wK1���b��I�	��gP�m�@�kT�:�k
����e��6]��m�qSo,�ۙ����� jy�v�����;�6r�+%5؃�	Y�S1�l��*N�Yޝ����i��9�(�c���q��V���vh<dɔa���J(�f0�{�|�;�����$�U��=�9�yJePp�,�քY͉U�8zbJ��i�������Sn��bQ{�\��蔘'�,���\;��S��'t,�Q��\/=�D����TY$��^��GJ��������.wP����2CB�$[H�
���=B��ZIF����������G�s���*�K��,0Ԣ�.N��K�T��sª�K��P���%T:e�����'e*Ejm#$�d�%�uGH��"@�ahD��"VV�R�U�EEt5KP�n��JlYQ�"���ny�A�&U�(�빡��d�f����YkNVI�D�Ȩ�4���B.D\�A*#2/V�!+�T�HT�*J�mi�U$XT\�D����ד����Ce�}]�ެg��)�t�{Y�S�����:Gfiޭ��6[KW!�W�B�&7ۤ�m��ӽ:X��ө[�jt4��+¾�>C��K�e}V �@©��c�BO�ro�:�];��9�v�����#��o?#yC��cr���7�����������v""4Aq����1��DL5��*Mxߜ�f����q��8D ��H� G�S?j�ۓ����ɏ.�v�z�?pz'���	8hߞr��|�W���9�t;x�����8�yNM��輻�"8DX�!)�@ }�5�sV�����N՟o����""�}�G�7�Q�~';s�����'�|v�ߓ{߻�������O��&����}����bw!�ܞS}|>.Ӵ��~Nt��9\��_S�<��5��״|}����̍���۾�������>��"�H��~���}#���|�F� ��~u`܄��}�c~C���������\N$��}߸�SyBC�ޏ�𾭹97;���a�s���z����C�>����yF�z�ִj��ձ�c�>c�7���om����|�8ߝ����^�}M��?����S���>��zq���&�~��e?'!���ۿ[.�ϴ��������9������ۼF��0�ץ��D�x�I�ذ�"0������>8�Q�]��@��N#󷷝��O'��P��;rr��=�v<&���v���|�1;��~���ߟ��0�������Ѿ<�7��r��4�������)�������D}³Ճ�nר����=��{NC����9�'�ގ��Uߜx+�n=�ɇ�z�c�e���܇��>�;۵����;zM�	ӵ����ϗ��?{���>�>�+{P�R5E�_o�w[��}�)�7������q��]����;�~��yW�>��='�<&�F� ���s��?����zw>�?;�S
���=!�7�$�O8<}��N~'�H����mv����eZJ�[�[���p��D��T}`3��D���~�&w�o���������Ą��}�{w�|v�z=����ù]���M���o�^�G��}M��y�����G�}�f<"��a��Dr��p�tOv�=��\���|B4DH�O������ߟGw���';y?}���?[w�����0�~v�G����$��?�����һ���{�'�����;^�q����'*x�mɾ!?��oϿ�~}����Y ��-wr�c1�V���9��A-�b��IbD���GL�2k�;]3��+���cB�yY���5Z��W�P���jZt�5CƢ-��(=ŹBh�G`t��V�QnaOQ�Y��o[��-�L�O�-?��$g�Zy�u��rR��^�­���y�-���a}��}v�F眻�����S|�|�}v����]'��{N~��s������\~C�aC�o�;/����|�L��}"�7L�Z׫ݽ��*�����rN�e�P�}����8�O����7?z����I������}��I�7�ޝ�0����>���}b8B!l�qy�"��yT�Ϙ���DH��O���}BC����r��C�����'�q���ɹ	<�~M����9ǭ��zC�a�~v�����|v�<%���~t�Nӿ��{!����ro��S��Uf{��>��ٓ�_�^�b>��#{O�~���ɽ����~O)�ߟ��Î!ɔ?����0��]'�����_�nNC�ѹ�?[w�h؂����|u���",G�(�<�{��/)�5uU��*�A��h�|G�������;~y��?�~��o�O�nN�o��B��c�w�������ŷ?S���Ν�7ל�+�P����]��toE;�8�����{tJ�Z��u�v�g�#��C��{�����������������?��/������<��]����}�ߝ�&���=o�}F$ܞO��<;s�c�<;rro��ÿ�9���M{�������.U�Y��w7�}D������=FDo�����׻�}�����raw�>����ߝ�p~���&����z����7�99���������>����ۓr���xy��9ϓ��jT�k��%m��r��}�"�}J��<�۴�������N��>uc��on�y���뿞M������щߓ_�w8��	Ʌ��x���zqτ9_q� (����E������O~{<�y�� N{�yS��P�H���"Dy���{�n�c�{C�aw�J��7�90��>;xWzv��,}O	�����~;
o�O󷟟=x=&�P�[���6��f>�>���W�I?}�B(G۝~V�+�	���w|s�Q�G�}�&>�"=�������0yw�k�����9�'��^��aw������?��w�����Ǵ9ǯ?;>�&_��ǿ�z@����+�w>C�W߅QKs���P՟��4���yw�NC��+�%�q����1!t��^��I��*�&�Ԃ�0$ȉiY3�� ����.p��[�\�)�����慴\���Fr�G-4�a��r�eg+���[�i�����1RYwW(h�ꛛPjw�\�������q�K�ݨ%Uh��ﵒ>�>��:����@_�w�i?&��|?������Hy���yq�Į<���}NNCۅ�F'}C�?�G���0���y��yw�}C��|v�=�&���y��n�7�N����`�>��X����|v��'�w����ۓrz>����K���w����zC�a��~q�<���M�c�x�ӽ8�G�ߐ��۹|�`��]��<�~CǸ����=��>q}�F�=tunǾb�Ї�D��=|w�~q�9�?P����xWe>{���<���<}��yw��n;rw���.��۾G�߸>��0�|O[��ǟ���T>�ӷ+��^O������{k{�pTz������g��^�����	�\
o���o	���|q���m������o��Q������)�P<~w���`�}v�=�~�]�>����gy��90��'���ޓ��rh�m�6�kӇ�;��|�|D����ճ�	2�O��x@���8�w�;ro�O��n�N��o�xI���#}?��ü�I�7��~����t�>O�݉?'�\J�X����7���|7V�q����u�y��\W��1��P��ԇ�>'&�/�{w�xw�9ǣՎWo��YL?c~C�Ǉ㷔�;ט���|~;s�A���K�������ސ������߄`��������R.��u�#�׾�>ޝ;˿~���7!~��O��*�S~w���|�=!��bw��X��q������nw��㟮�L*좞J?'�90���<�;þ�Ss���|����>�>����6=utk|�fv]o�n���L*��~>x����������:?;r��ǭ���(�~v�y������'�ޏ߸='�p)�z��v��'�çj��~'�� 9�]�}h|} t���3�P'j��Z|�o||Y�����w�.>�>b<>���F����%߻��� |߼q�]�4�q��~��;��/�|=~��oH�������V��ɼ'��<;õ��T>�"�>���V�cd3{ʻޖ��i������o����⏏����t��\��~Nq�į���I�'��<�������N�����7�?!�90����xw�}C�����\{Bq�������$��#/�#��H��i����Ŵ/-����ٛFZ&�a--K0���s&�� 9�OZ&akWL8���8��3q;�,�����۲x���ݨ+g6���C�-t鮮*�̴�Y��K�5���C��DR���05���ϭ��A�x��E#R�Ɠ�x�J#+/8����������߾���������܄�������<;˴�<�}O��N����o	�!}��||�p)��������ğ������;�s��v'{q�9�?^�����`�wQ�=����� �������|[��;ÿ>s�U�'���lz�x���_>;��k�os�����ە���>����}��ǧs������xNW��=����u&פ,[�<pO��F�>�DK?}�~���ڭ�?�Ħzv���ϗ)�P���&��s���[�F'}On;��?&��S��>��ǔ�C�q��c�ߓO�ϯ|zL?`�/ߞ�� �Kh����KM�\p��"#�����y�oܛ��x	ӵ��<���~BI���ײ��<;˴����?>�p�]!�>[�o���>!�P����q^��t?w@�.�p���gn�y~ػ�9���{up��ө�M�F8On���9A�#��nX��j�l?q�˝+���C}��
�/�v��\AS\$ⵕ�s���tf�"��1�8D��3��/��X*���rc�����	��p{��R�T!p�ԕc{:��;�"���f/��8��S�ـ3�>|P諚�T���`@LE����|(�g8T��勵]�K4o����z-��lGCc�w?����R��.-�`I���5 ��o��x�����r�طLB�u���YWݷSw8o������7�װ��@=���(�\٬�v7J���.�[d9�x�%���j���rЯf'�'���k�u$3W��+������?"�[r����`K��EZ���
>�ᛥ��fd<�괢�Hd]�R�bEz_}n��W=t����o517���F�J�8v����a��܂�}W۞���]�:�
��O���9xP�<��Ʈ����/�ρ�iC�����j���'3���س��'Q��(�q��ʎj�����ƈc:-��f�y�`�4�bmA16"o ��<e�`8'@���������L�;u��9c����Ga�:U����Ǧ��%ָY=jL�]VJ>�D2���k� 	�zľ��_W҆͜ڍh!�sJU�Ynr����m\7F�����v|'@�G|�T�e�:�Uݜ�[�V����R;_R$�}�Uv�8r��`d�n��v�$@f8|���&%m:7Eqں����d%ۼ�;_N��Hqo�F�'Pɦ�p-�`���<
��S?W�������z`��[�����ѫ��<�ѽr���>��5DZ)�'��@s��m�Œf:a���7p:���-Ė�ת������Gb�LK�u�]+����~d�.��(�ͣ�#��t��ܛ��NVxΖ����}bc�0���S���l���_�S�NF�u�[�%����u���Je6�Pv�5����WG=cͬ��T�~n�U� ��~čbw�o���+$�{>p=�tqAr�M�P�#�=϶��Z���]5.K}w�����-̙9�f넀5w5G��{$�V�ɛ���;�Yɪ1A��}���}����z:��{៭��K/�D��b�^8��� k�ׅ�,���*�&d��Vg�J���(�H�yWx��{�w?�e�B��^1�]��,�D������Fuy��-��-RyF����Ju��G²r��E{�h���uL��iL/�o*%�g���9~��za}r����;.�%�M5<��0���Ǿu֦�F[x@����}���NGz�X6���y�i�E�1��mL{�r�Y���
b����W�MiI��R#���E���z��˂v�ʕ�(�Z폮Hf9����2B �V�]�֓Q��+*7��,@��O:���C>U8��v�yI|$r�c^��sis*��5�E��E�vm����Cv���}��AU(##�@�}�����=/�Lu��f==��a%tK���b��>;��!��9�4yD�\ �
�H���L�x���d�.�h�b~L�c�_W�:H�pCeC���M�q.�A�2J�%t�}��ˑ<������5!Vhw��r��N7(����A��O����f˂;|b��}1���Y{w+��U��1�Ʃ�ɻVM�!m7�T���Z��Nk斏�6���\o]�����L���K�V�s/QW��odD�{��n���}<��L�]�i��}�ݍ���z�: �6"��824�+�b]NKf4A��Y�}�#��8H&�4N��q՚��o��A� �r���\��c>g�{��5&*!��ɸ��#X}H�L�����)-��-�\f%�LV|���T��pq�*���-ۿ�;��.����?v\չ���r^��.�_w�Q�$lA�3.�ug0|�>2�P�ٽlh�\��v�%i�{[s֢�8l?��p���36X��fӘ�Q�u"+�a�x:���(��6��E�]�i%X�j͊1�C��)���V�}&C�n�!�������R��/K�d���q���:DN�a\�����[�uH��2�(����j�g�d�1����r��Rٟ+U3��V����x�R\1����^g��=�i�IU���3��k����<�68���aý���!y�j�P�
�uEAl�O�dꠊ�d4�k��z��Y�;�ԫ5���Y�3{�_�醲d_�]�(Р7(�<Q\࿚]��<*G<0�<��_���mx�W�3B��A��qd�H���ӏ��\���[����g�����yfԱ���l��(�v�mk��-`L�ި�0.���4z�飔�"�c�qx�ou����Z��[:+T�f9YdJ�:��A���v'4�퉔C៪���G2z�=��5Z=	��2���:���W\������f����ͺ<l;��׻��#q�JȚ/�:�̹vv��k�!��}Do��ޠ��@�R0��巗����-�9��Q���U��SU;�Ù�;N7$GU�de�:�f�S ��Ȧ����nJg�z7��R@D;��������kgF�T� ��E�57P3[w#H�6So����<�3��x��4Es�j!W����ӊ�3���i�%��Z���5�L%&8�wYJ�Y�򱈙���w(�eB��]�K��:GG�l�4�g8=s���y���&�1�騳j�s��
?8�T�Y̰;��`
y�p����=j��P�Mw��9�:SM�V�����&4C��e���\���6X\##v~���@�4���}~�=BS�;����t)�.��Z;�4U��u�N�NF�@98$1�U�lB�/�g{�w���7�ކbOX�P��j߆]>~�x��7�n����I�k+y��W:3I���Vkd�gԍ{f��9�k)�c�*��^��u\v��^o5��Qh�����b��\�T��Q����?�|U���&m��M;��K.�ɉ�J�G%9/��C]��r-uw�9�R�)bo6��N�Bt�������!d;_��>�"nԍ|êf�A���Y1�4t����ꜣ�I������z�Cʨ������7Z�he�z��?U�,6���<kw1�7�C@f2�B��T�<7�Q�������m�5�o��T��ym��:gO��Wxt�_L��[o6#��1�d�����ꏂ������er�".yf��:�Y�\(C��P�y��LT���ò���ζ�ݭ$�#�s�*?����Y�5�(ƖF�ipP5��w:zcD0�Cۄ�\:T�b��"+��1V�[&��<)Q�j��<$���饧㦄9T;�	�I~�Ԗ_�����\!p�m��^��)��Ʋ�`�
�C<�����3����NX�,t��jN��c��v�Oq�oJ�{�gK����/8+�9,�t7�����E|O>��҄V'\����358��[�w5���C7��:�&��<dK?d#����w�PhV_�i��g������*��H�CU��d�"���A���&����lE������>�#-)�Q�C�7�3:��n�"�a��)��"Kn���o�i�YFQZ��C6��O�5�S�臖�K��|�:����gܙl�����ɛ��d�Kv��>�G�ok�}���t������|z��,����2�2i��v�&z��#�G������_s{�sh�{�w���*7��%�:
l� p����_+�U<D��;ˈ_�,��T�c���N͊u)��q�/��O���QjS&M��y���b�=�7u�������8��"��s�(p����^S0,;�u��Ϲ;�1��~d�.˾�3w]՛��}�~��O[<�y��Z(��.a��&0*0���S���A��l15O���o�L��6z���)�	�a���y�;W���}�@�t�~� �t�{�/�δ �4�x�Sfی��믳X'b��9��S��aG9��rj�}Q�m�>1�5�*��_%�.>���Eڱ��f�%�7���q�� ��ՑO:���,F.��5\!�����Qd���ea.8�}�1mb�k�M�?��W�1	�;.��Yd�y��-��+s�3n#���tܝyC!:�+9�7��ȓ^���%��9U���C�o� Q��Y��2�ۿ�ugc��¬v۶�F\u��;������du�^�<�,k�)qSo����]s�T<�͡u"��S5���C���C[�n�aI�)L���:5'�%$=bm[z�_Wg_ܞa��[q@�ǷX��op�\��v�*:�eK�1ښ��T=�"��luf���r�V 9����Th��қ�J*%�U���Vils����kyO
{�Ht
��T�@��kQK��f��r��I�ocL)�+��*��b�6V��T^9�!SR�2�-�Ūϱw4)��(�e���1�i�O����;���v����cR����1�Mݧ&�Z���=m��"�/4kTS9]��ȰcoF�W�>ǮS�qv\wj"51�h�h-0���7q��}su�I���G�P��vY�|&�屌������&Z���h��bIv�0۽��Ȯ�u�y@gL���Xzk(At)����m�9������@���>w{�q:5��;ٵ9GVZ��2�%&].�VK���a�Q�i����@��}��̎�������\t�%7�3bѨ�疴G���Q����Ċ�c9Q�807��ZlK��²���5`�T�:<�;KIFQm �[U�������@�x8�_.Ͷ�c��G0>��
 ̭�Xv8끊�]�`�օE�4�Z�+����'�w\��m_S5YNВj�8��zrU
ww�U1����Zn��e����ǘg��R���u�e3�1٭@����I7��I(�ޥ�K�tJ3)���q\��;�v�!�E�k���b�q�kr�N���W�kU�$�*ᔇ6I0��Ȓ'�+^��=΃��v� 7�6���s�%*�`)�&�۽��]�t��w���F��Z�__`GkhU��kyBtj�+��E�l����J��6�S�oXX���Mq��,��j�{9H��Y���X�X	/X�xP�sZ�53�f�h��(����#p�"��u����z�"�y�RV;���v�"/���}�'�%(e*���SFa�+w� �)u��ɔu2�.Q.sX(�XC���ƐՖf���3V�<Õ��
�-�a����gfG|��w\8_T=y�^(�s�[��hy1�p[{ڟQ�\���HjSY�A���@<W�yE�{~6�6n@�Vi.�g�����/fݶʴ�n�˫[��`�u.m��WNYz����^J�4�㊄�SV����4J׊�޺�|�����Y�������Y��	ρ��`7]j%�[�
.Y��R��`Ö�-�9��ê#����܏��uEs�m���掴.�y������%2�v�B�}�����B;;�R7[�iMw��X��q��
�&�.52��;�������p:����9Q�f�yH����uƮ>�A옦}��
u:�[�.34͜�͹�����@�"�՚:͞�Gv���V4a�ӛ��@c����:�x.����\C5�k7�;����Q
��)�2ӏ	A�pfs�*�*�~|{�����|���d���2�89:���Ag���!JY�*�S"Q"P�5iP��ZQr*���*���ADr�T���v���3���I!�*��r�Yj�ʒ�r�3*֨����DԨ��,�Ed��L"5"��;�Z	��DL�"�FiP�(�fj	!QgB��)"0�����TUQ"�Z%�NKą,EIQD�2
�i�V'�(���9G+��.�dVu��]"��"�:��ˡJ��f5�4K�d��e�T�UDE���%�"2NR�UUQ&IP��fs%�H�aQ�3XQ\�"�(Y
5�����U�Pj-$�
�$��)$:J�%FU��3%#iK4K�Q�RTij!�i�r�%:Z�aDRX�	�R5:j�Zjl�5
�iVeIUB�%��$M�$�:4$�N�*�R33P $�A �Gx]ld�y/u�}�k�T�9��$�6	tٗB��.���/����Ě�:o���+R�1��U�ŀJ�Tr��ΰ�ﾏ���۬e�l�7����«��b:I�2��tCƻC�[T|�wM�v]4.ۣr�;W{���A�����cI��X�p�v���@�7��(*�l�ee��n���
m��γs��k�滉�N�7/�t7Hq7� ڂ�4�J�� �V*�*�y�ʶ�x��Z�G��b��^A��~I:H������&�.hA�2J�{���o}�ŖV�uy�:_���	"�����ҙ��b�����s!�M�_Z�w7�]\@���n�@�Hn�30��s��U����g)������qh�������o:^'��l��Ѫ���Κè�i��P�줠��������2���� ��M��N����'���s5ܰ	�����U �K'hd�u��?T��7҄>Wl�za���7]�w�0V
&��P���fn �A����u�B�a����;��kԵ�bO} �s���yv�I3F��Y����C�i*b9��[������]>o�m��ڽQ:�&�U\j۩�w���P]q-�D���+�`�!���C(�QcxC�[�P�z����ZW��*��踐�\��o��aƹ6a;���x�f�׈��j�!�m(B���ͫ����Ed(��&S���E��؎(H���J?}��}+H�����6t~��_��%�����|0���p�T�2��1����x��#�[��Go��4�~���#�}qUY?x#1j�:�����a��C��39Ц|�ʊ�q�����v�S^Oך+�`�b���T�����:���fV���w�M���0v)i��]�
lC�r����p}�L���e�0l��30g����7h1���߄lS<�;����[�	�n�zZ{D=�����W\��#ĕF~�Q�e��u�o��/�P�,��p|n(�?WХW��RY�{$<6�H������@�Y��;��\���U���8��11�����+j��=�����!�":�-�#.�Z3ڞd��,��Vq7|^`�C��	nu�������غ�vD*v��^�E9��ʘ���o�>�=�)r��]�1kfOԈ�cQ	�&/�xeq��i��~)�u��Lk��CU�]֣�Ҍh�ǟ��/:YP�#��/�4ty�3�^U)�<�����"������Q �ɠ��u}|�`���l�5����I;�Ԓn���V�PȻbʱ�ԩd���c��oB��ַd���WV:P����|�6Y��զ%����v�A���o��v�6m^����y��G��$yI���N����}���o�1��J#�;G�MS%�3,q?X	�D�N�!a�6WV&�J�7�7^N�V�o��yӨ6���b�,�15W&�� 0�`a|��.��+g������F��v9�J�;�/pq��=Ur�6�4z9��+N
yRv��]��V>��Ze��`�� ����y1b8?��a���B����x�_�g[�����q8�.wpT�ܝ͖��պ��K��B,nŃg&���AZ�Yk�A�v+�%k�*�W���v�ԂS��pvN�@��N�}%�5{��A@6A�
����tԠ��i�Ȗk��z��Z�[ւKԳ�鲱�}�n��{�S���&@~b��Q�|��f{�1^|�v)�1r��V�\��1�*�7=�n��K�vB���uԍ��$�#�؜�@b�Q����sܺ���c��t��U�s�� h�\=�LÕ,o*���V\6�M�z�W~�������,|7]z�^?:Z�qc���z_��RY�p0BQkn8H�z:�VZ,��8h�v�y�e�}a���t�0ל�I�n��yF���}����F�{n��>n�_Y1<�%����G[5�0��9ԌZ�#�G9�{�x�!�n+��S�3U3�+&Cf��+*S��':��M�R�"EN�kٯgr9W*���W�}U���<�l����A�����O@��뎺��;u��C�8`���Fi�U�J�9{W^0u�c�P�9+����6W�v(�8���͂#֠]��}���:P���1N\t޽�1h5*�hՐs>l�7>n����n��L�H�EWBu&�w�3t�h�4��N{[�{�m��s�n.�=�#mR��a�4�� �w�,�����ElZĞ�3��<�mzS��6+#Ϡ��C%�<L� p��ª@�3�x7�b8wd�)5uz,��%�`���gh�oJ�i>����A�d�mH��`b}&��+�AĎ��S$���*�;z��R;ʏE�N�K�u�K����Ș�d�vw5�X�]ѝ.�lA������e�5X�P�;��[�I�����6<9�F���6�F���ŪpG����W��O���z�,L{F��R5ۗ^g�\�7�_M�gm��H� ;}P�2���j�9��43F��_S������́u���6C�]�6�P�6�ݕ���)q�-��TRw��w��\�ٍh|��|c:N]�;g�TY�"��j�J�F�z��r��u���ft�sq[t�J��P����M�����ͺq�۱>d;�	ku`��8k1�n�h圈��}�}���MQ׻���e�VD	� �䬋��P�9���&��[Y\5KVk>��`^�	�V���.�uN�v�p�OUC��n�b6v\d��h�/U���nxFm�;�4��2�#js�V�z���$�����%�"}ʶ�F	��E�VEڨ�C�o��<g./��Q��no��.�ϲp��<(��� �0�
��υ��~Qe�LS}~_t1��CTr��١ۂۘ�Bj��|Uc?_�� ��{"�&�$Qs���D�!�%�o[��t�m	6���Z0�I��X�p�7n����C��
��i9�_f�7��������Q�q�u��\K�QÜ�>;�Cuy�@k��`O葉�5-�H���(x���kA����@���ƾ��$q���}v��7|˫o0�j��L��E�8�Dw��'��,�`@����$�83�f��1��]nKf8C�D��4'6՚��z�=���j������֨�e*�]x����[#>�=�{O��5a�����&ry����\�JIF��������a�¾tG����q���==J�WhZ��&���W9���T�JTW���(��o
e��$�A���]
�{X�61izP��]��(��I�7�`F�*+�)i�4�����3bn�Y����*��_W��T9�x?Z�2}	�F��"�eْx"{`d���.�UR����^�6i��i;�=x�J,IϨ6��s4ܰ	��"~�U ���u�1Wu��~k�0����I`ξ��Lm���|��.#Ybڪb14<T��ǖ��T������q�6'�Q��B�tn_6;{�yt-���Q����;Jefڶ2	JX����:���&����y�27��r�Y�x�%��i������	CQ��u���%��y�_l�'BR�-�pk����kӍ#�]���M�%��?uL�����T]iuJ�-��{�q�=�k��YX%r<%�p��1��ӿP�
�tT@�)��Mlb�S��)�{�
�^�f�g�d��N�m�g���2/�TB�F������l���rW":9i�hT���I�6���S�}v!�n�>���z�}�=�(Z0�x�_W�4�q�wڷ;�;XRa:3�^E��(�QZ~EK��Ԗcn�N>�3����	%tՙt��ҢW"��z�%wc�PV�HC�lФ����H;c�v�̾ms��L�H�X)��it��u�B�h�{3z��CoxЊw��.���y��wZ�ˍr��xT�-]�fA�{o	DIҬ��b��	P��4�lB:�x��zpލ�c��'Tcঃ�������� ��K2�@d��f>H�頴���q@��y���>nH���쌛���zx򻳷�����$��F�t�_P��(����O�T�𽔋q|C�*��U�켷W�"j���u�2&�\Ƣ#���ӊ�2��N�8�����q�Z��1���\�k���,��]��0�;��F\��3	A�1�t92�Yj��$f�N䵙�����cVB��T�x̰9��>@w��~��x�GO�R3�o>��7Mv5�s�9b���5yq�+�e����7���健�SCl�?	�d���9�K޴;�r�HF7������)F0V�'w�5:ɿ��b6����E�7:S�;�����f�$��닇�TZ��KWh%f��s_��q�AN�qZʸ��}�+�Vi�Z�T�;0qC�K�pYK�]��ˎ��Gԕ�<J��	Z�ʼ>}�c}@7�S��5�q�:��CK��qW3{��Y":o�h�ET
�{�
�@xj�@�R���>�b\��i
�gg<���0Is��gQ����|��oQw,�,W:X:�V�Pav��-E��b�0|�̴��I��[�Fn�AReb5�	��B9	��,ԖIS�rS��}-�(��WK�v0x>s��Y���N���������[��Xh����"���φDK���u�i�O+����<n,�R� h��.�����b���:�]}��a��(ِ�1���y����1
��;>U��.���s�� )Z���o�Lh�k�CG��TE{���@,�-Wp���1�V��&b�Ҧ;!V_��}�酝N�Md��,�VkI�T0c��{�y�KU,wsV��5%���cNm�w:�sbk�k�9dU� �s6��lT 8d��<���uI��n��X�`e��]��ۀ�v�u)������'J���>��]B�T�k���F@p!i }7P�BzR�Bʥs��y�$�=����~g4���7]��cw�Ѧ~�`#�@\��h�\�������[�����&spd!I���z��I5hdC�H��f02Ss�l�yq11���Y;{5 Kʀ��(g�l��G�=x��{��Ӡ���Pɨm��!�`�����37ZB����q�$$뿼\r������WR��7�+�����50GZ�ɓm��Od�%�N8����t_�tM�B<�ך��k%.xs�����K{�������;0+h8"L��^����\
�"�z/�v��[��𷷫û��r�JɫaNM��Y+��N��ج2\R���˯�_���.��Q���Zc�c"�Γ��w�Q��f�gzq��/?�W���}/������v��VIZ��!�
��cΩ���S���iU�㮕���W�:In����vv��w�%�'*ۈN��fl���.�
�Fk�p.�I�����ٞ�8�\�=�Հ��T�H�S��CZ��6��d�/@�h�ؐW^�v���~�k2;���f�'�ێ EPz�^Ya�w/o�M�W�%W�Wʣh�z|e�Vx<�(慳�;���i%}��T�
���'�� M�VE�:��E���� ��ܲ�-Y��N^��
)��,�'����
�Yꑺ�h��p�Z:������p�f��m��ڐ;1;'%��_U�W��x]^�M"xy�KD�i{�[��4�/���qP������^�N����=�����Up�FOQ]QP@�T�����(����������N7r2�=c��C���s�����*����I���ꁐ���]�~�^X��&���<�jwm	Ա����(}'Yc���:^T9(�f��B<Osh�yO��ZCy_{��N�|Z���kV�X�J�����ب�ʗu��!XD�V5��+�Sޚ��r�8�Gh�S��C��K�
=�-�/J�ջN���+��I�=�i5�񍪴Ԙw�R�ҠO?��{u�o�w��}U����V��`-D��{���:��b}q.]G�9O��<4��`��(����W9�,��敠�p"n�0n ������?jN�,��Nv���l�'��h�������ϷȎ���s$�U%��0�Q%i��e3�c).�&ṎĞ5�n8(ތ�o���g��dʋ �r~$9j��E*�p:�a����+M�s��1i5q/�-{U�˽ԧ0�zL8�N̟xI�t�\�}d�i�����Pz�IOmF��N`��F�J�廸�a�%ۻ�E���Bd9���MCS:��d����߅�~;��Z���%�pm���絫�^Q�<!k�z��q���p�Sx�Ǌ��ǖ���Lsi
�0����1M�M��l�ؾ,�W�e4d��;
efڶ0�J���s�������Ox�{��,��ԺB���o`��t�T�,�z\z�:�$7�ƣ%D�5p�>�5̲dE��D;�%�Gj6��#�����_?T��Utةk��_�A��_sK�ඣ�u@%�����r����=�a�ior��<��Y��3uL{��p����k@L���Y� V���¦eev����c�Cl�U)l�1vF�.;�S��¸u\�:�����3`4bY�ȫ���0��ڽΤ� ��������.�"��X�b�b��ۮ�N��p+��!�(��Mu.�P��fZ��
��z��]򣆢��b[;&j6C��/�H��TM�+v�i8޸6�rnl�穚;ܴ&�Ց޷�mR��!�Q��\�ձ��I|:�7�3��ؗ'rw�s�*i��:��C�4��<���T�m�7O�p�X�[}����;N�U���=w�1N�o2Ȇ�,p��7w�hH޽RG�#|��S����:�I
��m,�5�/`�ڹ�M��t�h�pnV��U��z���P��q�c��P0���W9�o%��iIz�O������S�Y�B�������x:nIYl�����NXt��v"`�n�Wb�S��k��܄���JKt��CV�z�O��M]���z���Ǟ�gf.��:\9���|�.*�M���ݜ����!bt�Ă��bs�Y��T�2�>�Z��˩�j"���L��R x�kJ �2�;0Zr�o|�m�CoN�<+�#�Eއ<�㏫�<��� �x!�A�^�gmㅂ�of.��3\��gUж��<��N����3�D�}LA��^��m���	<�]+��v�5��Nk��k6 �g�{6�U�+�j5o�I`�7�"����t�Q���ӭ.HG���.I��M�Zk;�N$��j�t�w�c�ܑK\�]�.H��5����;�n�k����]NGRZ��Y1��J�E������M>y�墶�X���z��It�w�U�0���x�������<���8�Ў�t�]n��a��+8�!�}��^�6�F�dc�Ĕ���`S�k����ue<r��%U��wZR'2�VüV�GAE�b��G�Uʍ��9� �ڬy�)����iH��2�%x���pw���d1Rj��9�`G2�R�]���f}�8�7�rq1t�kn[]H���Y����U�`�YK�Z.9�I�������.��5;����9��OF�+5�i��)�i@1h�-��WYݵm�#���w��n�9+fˬ�=���!3b9]���F�7~Y'#(�b��53�{Fu<��tfj���p5eKi�k{g^-
}��IAsG-�n���"���
�#�j��x"x\m浱��I�5�d�ņ:]�V�ی��&���}Z��O1�0�%.��+��5���!���p<�qwG��qv�3�iؐ�=w�(�fҬ���D��<5��(W��*�K��JSq��𱙂g:‰�I�[������/Z �i��\
���EQ2VtL�gv�΀5{+u�R�����]f�	�w+�G�N�D�2�DP�(P 	�)Q.�Z&)"(�F�)
E�U���J"m���,�N�4#"�L������!ꚦU!�AF-$�#ʕe�[A+��]F�����"9AsPj�-B,�%4T*h�i�8�)�\�R�Y�p�!E+MB��D̢e��MYj$Q��L�)U�jRI�J�:i�r�µ��1d�*AX�Rl�ehT�lL��\�2�t"���2�Q��)k4�j�P�E��q�Y�)�-&]�Bi��PE$�AM-�Ι!EGI��,Ya��vf]Qe�JԤ��I�f(�Y��I
��I$�d��CR(H�ҬȐ�D��r��(,�"��h�Y�+R��K5�VAp���A+�gLCJ�)T�*MB̙V�D���
��EYE�-D�G
Ր\�а�)"|��]Ld�*	a�Jre�8Zs�z$���˝z.�j�I�Y�-����=�#��\'~cO\4ΰl
�}+���v���_}D@��'wk���p�ԙBx�����5zl,W�w�V�-��N��!Wz���}R�\�o��vu��F���*!�t�\')�ϩ�ċ����@V�?O�\�-�Dg��I�n�.�!ڷv!F�X�[��Cۄ��i���	�Bх�<I���+�K��"�߽={_,=H�����pt�`�B�OCRY���C�F>�5������K�'��wC�����`\N�r [5P�H�㯦���ڸ�Y�<�a���"5R��x�C��Vr���1ӫfo�"��Di�BG�t���	ǫ�\9K��IDk��3�n�vɍ�m�<�DҞEÙ�M����;�d_�d�P�H��$Ϧ��[,,��3�r��:n��Ls�x,�~�Y\p�,��\<���?]+��y�	T�Avt��"��va;C3���8��m���+���g��_4���!�`s�_`	�GJ`��P�,���)���I+׽��a��ʆ#c�屟&��� b�nX}P��}g���Tޕ5ÝL�F=��FU��n;�y�����zr��ݛW�P�|���F�S���'�V�s�Q$��r�LT(�)��*oA����"�	Bds�A45�z�b��ղ6��XoyFsQ��l�@m���#������� M��֯�Y�sE�/�׳xCD�����_}U[�̹�Ey���������6v�ߡ�S����z*o���eSN�ro�4���U9ȼ��ڴ���l���	�W���z��?r-z�Z�CG�=�����gJ�><��z}D�
k}��|3��,�SF{����p�a��	����×#��&ǁ�ܮ�m�ZΙ+1?b=R{wysgA)V��2��sh�D%V7�䯑��̩҄v �zU�x����YΛx�c���uH
�(Bm�i��K��ϝ�٦�O+�������C�1r���.U�{�B��<j����A���#���s�n��r���o��uԍa�֍L���^;<�����$���f2�����P4(�Z��dt���<{P��^q�s��N��W���]�pJ��:	:��
��R�Ωj����,'�5o�5%��+�jO�Y;���/Nr���Ўὸ�q
f�y �(� pt�ZS���T��n����GT�Ek���E�siqmIҮ2X�*%�!
�F�@�e��54���,�=�TD�k���k�%�}�`�v!��T�/x��kAt]��u�cX���(+QsljBW�R��Ԙ�ֺJ�s�:��A6�W<�O[�v���+�,{]K��>q�G�[t�gV�c���Rҵ�#���U�:��4~������o�,z�p�B䡃Κ���sJ��n����F���t(ᥤ(�p>6�g]_={���R���Ƈ�T5����MZ�D�a�N U+�p`�"�`�jPc�ӫϯ����R�G"��q�0�	��0�m��^C5�8 ��e<WQ��2��T����W�|�N#��f����o)����_К�"�ԦL�t2�0],,��8���Tk �q��I����B*EOa���+~8�����-�:K�CN��n]�ˌ8�?2jܸm;�/O2Yz(���]��S��/1�}[Ձ�;�O��<���;���\��hѽ�4��Fjt8��9�jʱC#�*p脤���@�k����sAD?av��+il(�.e����_^��!6�T�Ʒ�����_(�6�x	�硺z��y�z�R�!����`|��OeP ���.y�6N#M���5s������ÈȆd�aEˑ�,���V��ҪF�������p�v�e�ۿ���P[$�B��֢�Kl�����'��6"�/ �`_c�]�ETA*u�TP!�;t��,�D�筗F��h��顜���K�۰�����7�8	��/�t��ŔA�MD�]�댼{9�Ңueqλ�Q�����O�8`�ڵ�7��_ﾪ����w�[x:�$����w3�Iѱ{$��x('DƗ�U��O"��"���i�#^q�v؁Tv��٨��S)ӯ������FOQYP
�\�-k�K���̑�Z�)�=�A��5h}o��1��}P��Uc?_��!0��x		�;*���"y�'k�詧��ܥ-�g/�i��9Ʈ�"5�4.K�>$L�7#5�ܕ�IJ�ա���m ����F'�:w.�>:���m���B_n��mȤ�]%f�[y��" �"'Z������˺���t�ϜΈl㝬����-R�����;���ĺ��%���O�n � ���Zl^|6S1�^�7�yE�r��}��+�/us��@����D�����7�$9h�{�u�3|���
����<��[i��Z��ϲ݀)�k�4�`�Bn5�@Y��c���Y]���V�U](oo:ױ�R��m>�w	:�Nm@��ƺ#܁}�[����aF��JE�=���ԛY�**��e��7���]���7L)�:QnT�Eb��;� �XҶ�^��z�Z�w��r���62]�ZCV�)��C0�w��ŷ�\�/����ۅǆ��}-���<�u���I�԰������5�|%�ӯ�f{�ܨ��vF�������K���k�t��{Uvl�Z3g6h*����y69�M��So�%`ʎ�����]�I�Y�:`��|�aú�߻��F�|3*
��_M�T��끊&#��eO6�='[q_kM=�-楅���f���F�[�P�u@�|Q^r�ꖪ��~�M䗏5�-�L>k����)��ogYڦ;���_e�Al�Ε��+�b�}:��穙N�6*�������_=F�WYS�nAM���HF7�z��Z����)ĜU��E\B�J5��zǡ�&���o����g`����o����.��9�㸒�]uQ)i�R�_����{V�c�+��
1x㲩#=)�����\�L@���]����n�	��.�J|��9��ᡖ�C*z�@,﷦2�_@O����S�s�R�G(W:��>[jT4�iE��ac�8t�X��e]6}1PKHe�{a\��u*��#bҐ賓����S�҉r�(s��[h�Ԧ/�@���G)��A��ʜF�e�6.�7�!�/mvf��T�UXC!퍋.6ft}yաz�8�|�_|����&�� �z�k��_D�e ��t��3����>�xi�e�zכ��*��Z��������0�3H��
�nĄ޳��7{v�ul��;��?�r>���a�.5�Y�D��k}�&qY���ꆥ��˽I�:��<�v�mw<v��i�<ۍw�S��e����V]��vO%A���	cy��+䲭v�Ϸ��׵|���N�N :��/
s�gJ��y��j����c�[ꁘ���{/T��x���ʷ9+���6�MZ�J�ܣZ��C�繵�+�u�fQNFN_b�7� ۬0�Dob�Q�M�ie&%f�\󋂭m�Y��z�.�W!�_AW0.��i���r�}Ϻ���]�t.cL_$(���D�Ӟ��O:�:���:= �gr�Ѭz2W�OU��G\>P6Z�ب{��SM\K����@�[�׭��	�$�mq���0���o6�+�!g��%n{���v��k�+!��1m�dW�Z�K��r�h vN]h�4��\��c�|.E������.�9��ƬeU�ni�y����N��2�yir��(ͩ�u��a}]]����ǰ�]��}�D}�ճ�<�\��k�H_��!��(Z�X���z�z���k l,CMO���Į+V8so�PS@�*|�$�S�:���4��:�;m�m���C��6���mÛn�PS�/��} �����|ۉY�O�d����n�%K������|3��{.��ALw��a��� UȬ×b��5җo �B���rҶsV��:-����f����K�^k}��^���S| g�f��ds]��W�4�|��b�{]3@U�2����{L���+0j.�P�nV���:�rQ˙�m�l8�2j%��c*����]����#��#�
t:�ܜ�O&�9os��	�0z����<Lc��.��F�k�&9��Z���Ⱦ���S��P8�nM��_z�����m�p�[p6�ʨ�f�����b��H�I5���6d�S�D�Np������W3׍+���?`�����~ A�^�{�4��{:�i�%��
~��{[\��cG#�]1Ct�]}�&3����4�X�\�:��v�mnL*s�"6+ ��sf95]�zb"u>�PB�`���x���0���k�
��_}UG�k|�ob���u�nڗ����x������������<|�愺rmϷ��-�)*��3��V4��ഞ��G:�}�uF��]�v�=틔��uQ��M��큊&�!Py�c"%��Moic*� ���9�ڳ��1�E\�;��uCW��
�a�o�aJ�f�x��~F@ss���ޜ�����uU�c�}�l��"�cZz�2��v9�3���7��O��Ok��G�ec�g�Ӳ̃�O�r��iǷ��'��@�k�O��w��5��=�מ����]T@;����4]˷�tQ=�����j
_�^�WETJZQN�km�}V�cr�

K9�#m�\+A�@Vr�4������|�]_b|k�/��}��uE�7PW�393=���\T73[��ݲvKdl�}�@}�(swc�TF.�RzO�{�enoЬ�$B)����e�+a�F��mz�]M3}���4�ݍ'<=j���C2�eٍ��*�(j��7wG�]b�s2����oFV��w2�w�j�a����k�*+E���vHz��7�K޾C7PS*��Dū��9�I���ꪯ���ޗ7*��H�}�z�@,��h?�g���}���.*�,�_c@N�S�2�=���V�0��b�=H�|8�\��.5�i�涷q.�#f��i���n5¸�����aʩ�B�����g�紳��:v>����;Ч!��~}Φӆzq�L������M����hVN)k*�'zO]��[��}{W_.oo���;��F�U=.Ӽ���u��/Ʌ?ޯ�b��sX����W���yi=i�Okr*rj��E�}�e�ю"�c��_��UY^��Us�{¾���0�8��%<�iʡۋT����g��s����U�r*
�����Du{n���\6��fe�k(�0��LrԁIj���^�ׅ_�lͰ]l {�#�z5G�d.�)Cw��j1��=k/��W/��{؆�e����@Wp�\��̎�]^��ي(5˸J;�!�B��ˮ��c�4\"]̩��C:�o��t����J`7���2��jF�cc�Y���Q5r�J���62uK}mV�YZ����jJ�6�cv�p%f���e�|���'\�J�E�Ɨp�W�W�_T\�mӰ�@�@7�%��a�%J�kyoCYo^�ɧ֦�Hގ��;+.;(���Vt[��#�����+���2!ryp�kn!�z'*%p�뇬.�"��;J�O���GQ������Q���/pE_s�m�w��H��`����ζ��Y�:|�^4;��y�xJtj��A��qd�N6u;�sSyca66��L�ȅ=���d�5G\c����{|���oV��oMw'�|��1P�D���_p�ھ�|d�$�W�bu��[곗']�Fo*\���jL;eƸW�*63�g�j�S܏$8ut�Ŵ;��Kk���M���k�铢cn��=���Ld�jȘ����v�^aů�VW�j��I�ݧ�m:�\.}=�9�b����hjw:��F���w�-�D�ѷ��>�)��ׇ��v���y��� ͔�<��g2���m1y�E�:��k5w�t�Xud�}�u��Y�w�9�7�q[;�]�h��v:��f��*G^Xk8�lh�hÙbƟ��
���$oNv�X㽮�Z��ku��]�Q�/�R��le�, �}1ݽ�em�l�'�Ԇ�Rt�这��ڸ���<	��wĩn�5�d�/�mjޤa�v*�57�nd�xыp^��\n�y��Q����� �l����cöf�Z����1�m!�\Ť,����b�=��6t�r#F��O/]J��u6(��޾�q��"m���5N�;f��q�f)��Վ��rt)m�Z���w��ฮ����n�˭���E����0;g%����G�N3�7R��Ӄ������mk�R����0j���I�$�z-9�����}�CYw��ds�+�yuu`�i
��n�|#�R��jrY[�-;ڕn_�e���8��
;6]��Lr}3kmMit�Q��Z��f#@�*n��v-2��د���6N�bc���F��v�������l�Q:\��[O��̼��R��vV�~Ik�ܴ�_X7�ʆ<�Z���HI����{Ei�|��钁�g��9h��F�d�F�K���\�t`}���%���DZ�:,p��΂v`�Ǖ�f���'j	`��3v�O���*�M�q�7��ށ
��I�����;�5�����Y���S��ьV��;Y����T[Z0
=qLORwn�99�uՒʨ��m�����/f؉��[�3��R,�/k���Y��vNs��(�޼E`��]=��[no.�d���0�+�+�Mˀ��;�Q�%X��}[e�gZ����e\��C)���氍^��ݲ��8ڜ����=bA�:��AL\;��s�o��a+i�,d�ً2���r����j��#����g� �1���e��d�ͮ�r��:��*Z�R���c�f�w�w� <�lݑ/�+$$)m����ن;6�2Ax&��jQy*Ν��&l+^��읺��.�T�v�n�귕:.D�\�î�����u'����E�hPgO�p�b}������2�o����)}��&o7�86�uRS�p��[��>�O啻9,�Υ2�5�gn�K>5�?�i9��.���Pa��]Ԭ���s�T���������;B��%(��O2[���I�-Z�t����R��E�o,EJƇ'49�(rA�1�R�6ݎ� �/w���u�+}�`Eo-�K��#O2�{�J[�sj�
�y��������P�,r���*�!O4p�+_7����fje�"|�e>|n��լi+��r=B-WM��m�v
���N˟ٽ(!��R���v�}�.���ɕQ_bX
l]x�e6�{X<�ө�I�Uo8������6Ĝqt}��  P����,�̅FVi!�1"bHT$Y,��W+�eApT�L5A#E�"���YU�R,��"jHUZfDq0䈳�-:%�E�fl��#I$����%'4�RI9�T$qS	*���;S��@���eIr�-I*�K�e�b	QIʉCaҰL�
E ��N�Gf�.ZTJ���j�iӪZ�]��E9s�f*B2Ē�3-�p�Oh%�)5$:��*�)��GJVDX"*�P��da�t�# ��D��P-J(�DEQE��˘V����i��;��Z�y�@��*�.U�4��r2�w��EJL���Y��Bi��6n�TQQN,TJ�4��C�d�r�/\���(�F��N{��<S�id^�p��8sb8�Ϲ�[ԕE|�!��جS�2��������1�r�1�^8
�)�̌�]���cw#Et���������V�X&G9ܴ�kY�W��d5��uȆ������'C���y�г�J�i�R�+Z��j��YvWAv̵#�O��5�����{�.�2x㓽�_$4���K\�^o��γ���c�ͽ=��|�)q��P�1 �����N�j�kUsx����}�:�7x>5��{o��W#=n�Ӡns
��{Q9�:��ҍo����6��T>΂gl3���m��c�k�gX�U�;�N"J*�-����hn�5Ww��Wt^��ik��Ρ�yP�-�6����F���p�.��q��.����7�㴕/g\Ӗ��ֻ�0�%b�ﷰ����:��}Y��H?��O��O���p�5��h��lir/���8�|z/5��HiNR�w�&4������.���)&����8�o"麀Sn���w]M���U�j�*||^x�F�u]1�_�Ĝ����4������du�|���6SԲQ���[:�~<�ެ��z�'Q�2	�v�^��t닜��9>R�c���t��nb��&�|Ї���b�s�rW��t�XP���i.dl��DG�DD��{���j(q{_
NjV�F�:�o�K���4��7 n�
��-WXuΤ��=gW�*��¨l�G�
����}�ݬ��4*�P.�*� ��mƸW���6-l:U���]�$������n�}��)�|�Zp�jr�q��?	c9�S0g»7ں��AL��{��5��Ok�}�ίj��R��8unFW,��o8cp��E�Ͻ���juK�K���ڒ�gj�|�/�OZ��]Osg�_ovT�G"��F\ޜkFeAۘ���<��΋棞��\tf��[�b��z�]Ě���e��;���~8�����1��n����u�{m�{��w���&:�zr�k�f�5c9�G:�dɞx�����_Iϧc����)�}��}n��Mmv���4:����įb��f^�Ocgi�S��h\�	�1���3�Wg�1��jSh�9�,����v;灸�x�.v�v��oL�8s��^�k�����bf�[�q%�8�������lb��1Twp���\��+��;[W[$�h"sv���:��U_}�R~�'O�Hb���z����=e��=���ih����{�Kf�՛�4�ұm������ETJZQN�ko�����7��@�ʆ{��N�m����/������T_.�O�D9}�[��κ�6k,k�v1�F��1V-�*����EH�	�n��*�E���Ju�W1e��*�kzy�	���#�)��]2�\G9�`�3w��y�"��+��3;��X,*�sM�l[�<��R��^P3�_�������S٩�a��'7�s_B���*|ä��CI�Mƻ!;#gs�R����]���¼�\�s�]�Jy5��N�p����N�mƾ/�Aؽ��X%!�<��"�s�/#C���@Ο��:��F�ڽ�����'�[�v��=��ڬ|FZ�х�F*�8������Ϗ,qڝE�'/؄�c#G��bp@�39�����}z;���O�>�w[�/Q�um4',�K*F��\�v�dh�W�X��ƻ\��[X�*���k$EɯjҧG�=f�)h���K���.V��P6�u;
-��%���7x���E-�Ǯ��}�W�}���?���(�D'C���5�5�sz`{DM�T���T�!J���-�y=��΂V{���྿/o��{f*���:�T������Ї��Y��{�o5��TM��L[p�R��=y�7��^��cw`��ɤ�X&��G���*�=ˡ[/:���-�د����i��|��S����!M�����*v��r;��S�*�J��o����	��N��$�Fd�����,�H�Z��h���[�'��uQ)	\�\4�mpW�JSv{��
�C����T�|0u��]��Ck+�'��,A%R��S�w8+;�A�s^�63�"�Q>q�b/���k�I��k[������x���5*�crҶsU�{��cK�s�#�tT�Lߦ;��G��~��W����/��ri|���!�b�Ȗ��{>��q]���*.���_l�����E��5 ��&��Gnmi5�(�w,�䊟0n5|>W'��������V��LG˳$��N���(� ���):�cG>dd�j��9+���ĺU�+���0���77oW0$�]����F����kz?}}�f,����o�Nj%�Mf�\��-f��ö\k���__�n�7����s|�׻����enQ�s]�ky�MI�M�F�v���{�ip*w+��;O=������q��E�Wχ��zy�y���0�����l�ɒ�5B.���k�u�Lفw��ý���M?x��u����ɾ�PEi��tW�*��CeM�Q��A�:�ܺ��3���u���q%��TLV$�|8���N��Wnj���m���c�Kޭ���L�Z�nr��ъ6/��6:��+�߻�Pdb}ιK�$\�K��N�t�R:�;S�X֪6*��)��ΉIt����UP��}�GV��y�*Izs�v�s�C�6��WJ錁b�L#�hu�����'�
o��A/����(��GH�8��2���\�c�զ���dR�6&w;Z%q�[e�M�j3j+n ���[�'��$˹ݥ��;�#qX��J�O�R����8t�S���	���]��Dk&�E�k�o�]��-^�]�:u&t��[&4;�[�����oI,caK�wI��}�� �YIc�$6��σU���>Y�m��AJ��*����,����7��[�ʷ�GJ٥)�X֯�|3��ct�HY�o���5�A�yj��tm�c���P5��}��D2��Ʒ��ڗCz��\]�ܨsry�K0h��1�8�����˫I��$��-}�cU��c���lhb��+.uƸ���_�鸉[��Ρo���g�%�ْ�+��p�l����C/U��"��#��ڟ�c���Fr�1��s<VYg�z,/^�M0zq��L[�B���𹮇�m�ay���v�$�yy����K��m>�|��Zp�n>�̧�"�~��<���ِ9�1��f8��Sչ�+&���'�[���r6��U�	�H��oi����YV9�M��1��o�$�qڝE�'eK�p�ֲ{l_��}�b�CG��둶�n,���otfp��{]O;I���I֛�6�R�����٢��1�]|W?w���[r���B�f��h�+��QgTt,���	�#툞�[�:�l�o*�� B�me&,I���ӥ��[p���\����_}���,�}ﵾ�5�c0u_��6s$�q_4�:�iVᐸ�]Wy��[�8u%u��bK5�SWѱo�K���j��^ڝ[�C�U��Ųw��n�i��d8��m�¨�׼���<$��P/�ϥ��V7�3)�对G`*'�)���,��M>�uϮ�T.�����h��hD��}�{{XR��U.�WIR�n�ְ,&�ڛ�p('�PB���=�v.!ˤ��n;�-��]R��S���������p�&���������/���1�yQ$ń��Wt�Ƣ��gma��̙�hs���R����6*��n'��D)﷤�ih�	������-(ӆ�ꕹ�
�|���f�jf�����i���	���K�i�:Bꁠ���V���9���K&����z�t�����4�|�8q�Q�����q���v�l�~/�x�Ǣ�B�2�S�n��RF[�v����C��a���GR��,%�W���ݧ��V�'݅嗜�Dl캆���9��Oi��B�o�T��fK)}��{S2�TQ��h|sK�d�b�=M<���ΜO諭������Y�;�R�D����o�O��4�vˍwdJtD�!����è�&u�x����wz����{dg}
s�V隆6�jӆjq���nJn�O'x��0-��_J�8��F��ٮ�I��.�x�#b�+z��޸��J�������D'f�X������m�}<�njj/i:׺�v�<�˓�)j�g%s��kY�k����F�9�ʂ��Ѽ�Oxgi�Yú�j�v�Q�a�=�e�62%����c��[�g�8$;4zp<�tJ�<�ւ�;y�ջ��%CV1E�C`��.%%�"{�)�iy�xI�˧�x"�M��G�tz	�΢vUN�kAj-�����4}���,�Ǽ����uiy..-�-x�t��-O��/���TbT�kyp�5����"m�؂�seoZ��W�9��0��+����+�*����t�7^�~�O���L�XE)�[8�YX�X ٫�w|�S{�������ҟ�z�MӣjmΎu�0%��U�@-�w�\�ջ�.2%k�utw])��Jh���L�"X�˨��Jep�|��S�(�1���A��W7CS`�ϰ�T3{{B_����/&5iv���]���ڏ���i��x(؁�$wm|��֛RA�{��'!�=��k͚'�����Ƶ>���2��V()��zL3�K@yXڝ��b���o �8:�O�������͗L�!Lw˱˪pmJ����Q�1Z��<��5X��$ҿ�|�8�Bob���m�l���n���o,s�5��_�I[sy�.C+�2���.5��S�0h9�MN�e�t�����8r��j0
t6�ɨ�y5�w����G��z���i桎tOp<�3���ʧ�"p����-__/^�\�uN��뭹��Ĝ��>���ᚋn���*�0�׹o�U�ʏ�n�y�.�5�sכxk�Ɲ��h�x�kY��=�UF�1�<֧ۛCڒ�=>ާзOw9=�.#���4�.ƥ��Uf���9��c�]�~qzn��a-��bAҹW*��6Fs�0�#��9d"%kt50�ӭ�X;n�@�-��Gj�qf����N%m�o]�0���	D:�+4�{����
HYE�3�0ri5u�G���z����;�=wj*�e��L�}�}��v�&��[�>��G5Qs�SQ1|����^.Mf䍞Nw+�T�{�v�j�W��er�DK���X�
1���7����e��޼=�.k�c�o6�oUgYڊ�6~<��Q%��j�J��0�Y�t�#;���1�.O��I���]Eoՠl�P`>Dw[��ћ3�b�uݬ�ܣh%��5	���5��=�M=������D��T�dV��I�]9�18WET*[5
S�kZ�|3��n[��輋++���4�sN�\�;f�_@o��r�O�C��l��ϛ�m��R�w�"���U)����;%��k��KE���.�\r�I�l�v���w�s%LP��]\h���{ݴ9C����9��rt��_�y��f��^3�v@����� �z���3�8W
P�Gpq��k�}��U5��;��!�Fa�COe��J�M�.N�:��vEv�	�0k�Hd���V��8@�g�5v%���*���s7v3QRl}]���.�G$�ʗE��]���=���^�ro��`��e�ΥIb�o�/���wڸ]�Y)֣zl�N����`�Lj�����˵P[��]k�>�Xނ%�C1Td�h���0:[+���or����|�3Ec ��WX7
n�����z��c�$�L�hJ�.��'&sc�e�mt ��;��&��B`�%\�ʻ�P0�
��9]6@躖^
6�51�a�!'C���/�@)���u��v*2Sk[Un_X��F�Ù1���"��ɍ�Q2Y�<��+���j6xu�w�t��"f�P�\:�
؉�.d>�xlE��>�ذ��պ����c5
罄��k�ϟz����%�����uk-`��Q+�wHA]��yy�c��A�`^�^v�i�v��q� Ҭ�:�W1�C�Թ,�P�mJ�y\˫�Q����^�����p6���P2�c�������t��KT7�s{2�K ���h�+i<�Z�(��I��!1`�Rpq�u���0����NU�1_0�ڌ+MJ�|�;��{xh7[G]�c0�].�u&	�N���wVPs���U"6�_-;i஫ݮb-�M��P�Y�������Y|��	�9��IY,%:܄����w��{x�윊�_���mⓨ��%�)��+k��R�*���֧lr�z����d��m���N��d�q�!�}b=f�k��Eu���R�\�vu��VD�Շ�]�١���v�a:�{)�c{�er��͌m��c�IͭkGw�V���"��ΰ:H���[����}��g�gMe����g1�_GZ&J��TJ�fQL�6��*vC%)N?��d��)Ig&�e��I�BV��0��sx�P�Xr��ƦWl��r��KLP��j�lT�[� ������B�h�8���z���,��L0�^�W�X����cKfԓ�u�HՈ���s�V\����9��;yƑŏ(�y&�V�}�-ǻW�b�]�.�!��.m���������^�0��T�i�Tygan: ��ٜ[�Jr����C���#��B���OI[��+8G��N�N6�M��AS#�[v�5g:��gh�̲uI8�˭�]o�m���:�y{m�c���+sr�,��Y��coI\���۝ ǹL/����QP�n>u{������¹W8��$۬�i�$��Rކ�镜�%�s1e��#np��JQ�T���S^%:��K�����ԙ�����������kn�p=�'jv��\�n��R%��8�1a�Pp=���m�X}c1i��3�iI��g\�T.!2�d�Y.]�w��0��@����1so9R���íʽ�]B��+��YrO��O�|@B�T��̒<K�<���M1�IG	3��e�����)��\���uwO%�"V�	tV\.V��B�p��Fs�+��(�h99Nl�ɺ["����Z�����J�N!���:;��+b���a�5*�(��el�ꁬ�T��Q"e�G3�;�=�4��BW=a@f˴����0#�$.#� ��R�,X��/*�.��i�C��9��D8a�@Ў���r��IXeyN"�;�8I$�8��R��F����Į��\*;��xl�s�S��xw2��t�(�gI�H*�	H�jg���v�e̏E]�kU'wr�N���P�W=ΐ�b%���R�É�.VQ�4�wC��y�լN�ZW�"�*��MV��"|g_V���xr�}zo퓩v�H����f��u-�;����ۻ����z��G{n��B��YyuHW�!�����;Ė��$l�ѿ�>�Q�`�n5�Y��"c��V�_���Վ��5��b�����=��^v�wU����p�D6�m|�UDk�'X��x^���ѮR	eU$ƷR�*yk��T�?{���W?+�z*1%�d����T�7�9b��f#o�J����״�E�ߒz�	8f~=�9��8��˓�>�6�=r*��r,�Do�]΢����ݶ���FC٣�K���N,'�u���)�Y��Km���J��z���j��-�,�Ķu�O�-��Uٷ⯳��DS�U�:�8�Uh�r���xض�!v�J�{~���vZi���֦��YS�m�09r�rw�/���d.s�˔�to��=SO;�7ʴw�û)$�Y�m 2`���o]R��R�[A���쩩���z��kh�^�m?J��qw0��_�.�%�9��c��s~���!��	
��e؎���cO6	[飂�O%>5��m��Ӣ͵�-��2�Zv���Y]�����1S��J�4�n��!�G�1I��s�MZ���Q���of�)�׀�㙢��آE?�_UL�����_�5�V(%��Q�&* wM��_zI��)j#q	XkF�W�J	s��u�c:���.���
~ﷄL4�W�>��/�t�o��Kq�J����z�gpT&��K�j
c�.����`D�/L5ړyOs����P7UC�P�5p�����y�qE�3ӤWcU��⌷�Δ�r����'9>�\�O��I�l��
��0���*C�!�{yj�:y݆����rws
W;x�����ME��6�\��<ܺ98y����Z��J�"��U����,��?ET�<כ;�ht��Wٵ��(9�X���D�qp�#�	�W���}�H��3D���'����N�B<��{yJ��ŉ;A��n5��t:��ͧh�s�_�f*���|�����x��ނP��OՍ0�6�������Uo\��3�a�ZE���b���b��>5!�2����'ֵ�RZ���e�����#�'#`TU.�r�T���ӝ|lu�I�Ł'�-���/B���)����vް9�u�]Xڱ�4�q݄u��f�læ	��S\���ܝz�V������|�t)�D���N�끎���}�j��odO��>�4���� CT�Ձ��U����]R�'\%ze����z��v�/�������H�5�����SFz�>��Z�w"dN�
������1r�}o�V��˽ށz.B�ۋ��rq�҆�`;=F��BNzBR��v'd�^X��)�A�o�=zS��m���}�T�0;���:�dd��u�|�uG`*��ֹ�r�.ֻ!�ί���.��AO������S�%
=�Vխ����A��p�w؟mÖ����>o�T[ck�t�B!C�|���֑��sʕ��рV)Ok��F.8�I|��ض57���g[�Bz��ק��j.!�=@����Z�nMf�!�˙��㒘��d�B�٣�$º$k7��J�pU����fn&�؝Wl׽��{��ڷ�A�w�q
"z2�ۺ��f��!s����8�~=R����O�pOb�S��3����ClҔ��P6P�W�F���A�Y��ݠ��!���u�s�G��Z� ��+�3`��I�R�m�ᵊO��&��u�)I;�I�=�
U��|y>����3���������m�>
r�]�;״�%U��|vDzx�S(H,y�f���v7.�^���m�'�[p5;��]��:)oŶ˗�����y-v��r�q�ʢ����K���k5��{�_+a��&���X��k��;��*-�DIX2�TMcN�*^�oF��]��e ���;#�S.oNv��nc�����ILu�Q|������v�_7φ)l����j���Vu���ò����s����P��,ݭ����yf+Db�-S�K&�e����/�o��γ��l�r�P\#|�@����b�0O[���x�m>�I�����YU�l���˭@*c-���Z�-r�:��F�9���Y=k�����n�XS��9���Պ�vAד=�d\%z�kߣ���R�P�<k���V�e7M�eݠ5�1z�uέ��.�f�B-wlL�v�<"�K��\�w��0R���Ւ�;�\'���~�W�k|5��f@j���8�p�'��ʦu�u��pH��h�
�`��Վ���(�J�R��6C#��v�4�����$�۞ĒU����M��7�|��]�0Ou��Չ�/��gnD7�|�&��`�����s1X-�.��!�|����]�×V.9I4�N��R�R�D�Nw��`8�8GpSob��f���φ���Q���|m3�vs����pĤ��<Z,)�=���8ø!.:�ڀy��+\�Z��i�ۊYU��uOb��r���C�}'a����k��&5��j�s`9f�zR���A��lړ��˖�ov�-�%�p�|ہ��Uk�/�5p y����2e�����ӪN��ׯ��+ڷmKیN�"�R����m�J'���Ʊo�����P��	q�Gg��[��T�w���s� O%@�s�nz�_��$��y^�d�\�y�nu�ҋ2��cI�Tн��ݧoF�'i�) ]��[���U��3(���ި�8~dd�e����Mor�a���LC!�'�M�n�@���˔��������'��i{$>�b��� 7���7�Ӥh�Å��gtM��n���󥽳w�v��!��sU�5�ױ�ݺԺ��oNFs{2��<JLG��z؜AՖ�Eu�]}и��hc)-���T���"��TN?�p�6փ��)���h�ؘ�v�,�T���֞.�:Woz�����-�ZB�ؚz�s�S}P���(Gssq�gF=Fz� %�́����e_�IR��kyp�5��=��OL$T`��Bʤ������)���Ȅ�~��%-(�{�NFu2�����)i��C���)*n�PR�ޒ��I�s��ε=���,�kԮ���-@��qO��ם�O\0B�N�
�τ��e���R9৷��vg!W�{<=�|�jX��M�ؗL�!Lt��C��d=���sJΖ��[���J\漸�$��2�.j�|��!o�;x�������Ǌ�o}J�s�����%�MFrt�I�i0�q��,��+�FR��9�F�[�:C�X����y<�j�m}���6�m8e�{�T"��^(�0F��M<�֘��F�v:��j�𻮠o)�۽)��|K락�b}\�:gWǋ��ī�5����Qk�I`�s�,BL��l�Ƿ���V'ǂ˥V�}ڼZ/�2�ͻ�-+4{�h���؟����U�ک���;6ۀ��s�f�_�E������3��YV��'9뼂�J�m]w�~B:��J׼ᚋtΧ����ֱ�-�|2r/�|w���eX�=�;�}���e�˄�kZ�k����7_s�_�f/���H��v�=ݛ����׻��lb�k������sx�7�2��G!�����dPRD�X�ż
��
�_M�TD��b�䆞ԁIoB�͸o;�:תܻ}"���K��N�wW�:�\�N�J��V1�OSz�>��22��Y�e������Q�gj"�����I��}C�u��M'V_S��9[�z%[u�_]�t�O��}p��X��hU|=8��<�;44�m?W1���rE���Ɩ�>m�����-�6�HY��=G� wG*]9g���l���ծ���>�r�.!�k�ꈶ�TK���)�9��}��0�u���o�c��1[x�*n���dzn�u���B8J�ԝ������p���ro�>�G��3�-�S��d���d��l
u��ft<���"v���i��=�C4��1W�٧���O�cV�1\\7�⒊�-��Ml�Ux��c�VN�]̽s��Woo
���leP~��'�Db}�ZV�j��E�6��L�wu�A�뚛������+]��1qʄ�W����2��|�h΀�a�c#���QŞ��]CA+\��9�9쮜}:xڋl{��LTklOE��w�C�9�D��	�6v6�
ܓ��R��8��կoo�Β^zza���-��ڈ�dLG!���v�'���&$ש�{\{/��4�=������'����O+]�7���!��M�)��[ӯ�n8�[�+�m�ju�nڗ��Ƶ��uCܪ�Wf�Fl���Շ�����u2���F�앃/���>*^I�Y�y���и�����y�����Bc2�.��ɹ��O��
<���f��<i������=�����Y��vX��*���%�WӪ��f��Nd��f곳,������ܫ�Xs'c��2��u��c��z��k�5r�{�#S����8��/:�q4�M��u�����9"#k��z�|YH<�*����� ձvHvv���	����u�R�B���^KW7kէ�e���4�A��8�Y��m_�s˧�iv�h�]�*��>���f!盫��z��_��q���������I����]eUhݲ�)�#P}�������'rʔ����e�C���*۱at�S�I�ô)�`��2����(6��躔����5�vC�V�e��Qs�n�l�]��I�LP�﷤�!-9��]���/��}���Cec�o-N[��!�6�z����]�%-�Z��.��\q�r˝U����M���s�ϙ�	�������.��O��nd�w%X����ǝ��I�E�P�3M��a�Y�	��v�t:�ls�8��)A�X��Z�^wF�.ud�%��>O���&Bn5��1艈�6��Bd�(F��Z���p6���'�M^-�[�ѫNm��k)@�N���^�U��۳��:�֫�@�^���2����k�Kw+���z���$�X�����b|�HY�Ӷ��m��r��]{NwSo���Qm;t"���z1�5)h��p<�����י�'5�6�pt-=� �OwjU�Ɲ�f���-�H��{�᪅�]�53D��ټ������K�����>������(�Gx�
��b?N�bE�Q.?�;ʞ.���T�ɢ���e��g��_A$]==�g�y�n��~	���,�F��)ڏfP���o�zG��D`�p�y�y��^.mf�[՗g9��*��|{�M5�|�����j�(��
a�l)m�®Ͷ�gQݦ;�&�ٜ�P�W\����1�Ih놻�2ՌlT=ci���>�S|pne)��Sc9S�[�h�#�vxp[�yW�'��i�RT�kyoCY=]M��o`܇s�"�c�6�HX����*��_�t<�=���d�7s�����Tu�c}ᢇ]�l=�|1�o�+�邠����3�ٝ1����י�s�����q��63��e�</���0��d}�9D_%��or�R���,����t�`�d�,��@G/�8�����z&��B��!�[giy�-���]����P�C�fs�;=P�e�r�g�&�]
E:����XL�dbX.��t�8u�O:��i���nKJ��.�vQ�\�N]�M�D;��n	A<huq��������3�>?E��0]�w���	��(��v�#�SU��
骆h�n�	I1��wzݭV��r���hgF�7��88�s�»8sQj��b���n��%�(ʚ�*�Y8PZF-CK� Y����g^o˘��u0�k����u#�(]f�-%գ`��:P��|�gS�A�4]�QL;��Sc���i˽�&q�"���ǻ4��.RC�\iFb}Z��97���N���R�iU��MӬ�	��&���)Gk3C�˾u�2�Vr��3��'j�R��ކ;�N�l�lAƬgi74ӎ�h�k�WT;=ḁ���+�rU�Z!;ʳ�_�e]�m.#�'Mt4�{1G܆��C*Օ�5��x�RU��q�����moٽ�k%;�_	�gG[O�N���uC�õַ��:�]�pm���K"����!��<�P�̶�^ڀ�ćM˕h}�ao^WX��|�NCr]Ԝ�r�Bs��ȿ�aL� ��ݥ"�wo@�,�y��}AQw�Wp<ju�ztD��w���\Z޷N��.���w\��tu0_Z6]�.�a9��u����l�f�H�����e�4(۩G��q�_S���9�7iҥ�Z)��8�uۇ0f�~�	,�ޭW3�6�QVJDޭ}+/xr�Wq|͒��)C02���h�I�vo! �����I�֎�Qۊ�gNM�����7�;0cY|�@�Gu��<�˺��Inڐ���յ��yi�¦˕%k�E���Z{[yɓ��NeNW����\�͛����n6��SoWl(�xee9[�����I�&
�����K�6q��řzs,^�s�F���J�iԽTėb�ݢJ���c&9r�&,uwD��C����O�g\|f:{b���\uR�f���J�E�\��vR�;{���_�*e��5Y�)�r��N��'��Wt���ޝK:J��=Kb7���@�L��oi:��l����C�=Z��7�ݙ���* 6��FZ�Y�ŷ87+a���J(5��j�9Ri��/�)Ծ�҉��t����ɮ\ۂ�.�������ȸb�؛ʲ��B�<����Z;�'��c��K�]o��yǙ\��ڦ���uqۊv1y��Ε��z8d=7�-�rԚv^�۶�-��s�xeʆ<��\�\r�;��_P�����&%�2f���+M��.��*���|s�p�$���Zv��Y�J��{Ûo�%�H(�k���qF.!��%������ L6�3�<a�f���7����GB�AYB)[V��4�m�#e_���.X�eZmԅ��.Ĵ"�*�Ú�qԠ�ٻ���L����G+V����ܜ�e��㣝ɔ�\U��(��%�8wt�"��H�;���괨�$��Qʍ����ȍ.+��Cs�,Zy���MXFJ�Eg4T.Z�QI��CB�75
)�D�ˉ,�$:�r��"�����-̝�Ъ�YU�i�m�j�c��k*�YµT�PRuZ���]i{,��9Y��T%��qGi�q`��;��u̐�QFd�зGs��I7$�W#��LS�ic��8z�Z&pQe��!B�"9ܜ�7q�$1St���ZDA\�y�s�t�	,�
�^{�Ty�[B*���UpL'$'$Չ�%�*�6^�Rħp/<4@�A��Ert�9�J"��Q"�
7v������h��':t�  i �� 
�H-��g-��B1�R�R�u�r�����A{'v��u���]���d/��6�sޫ���FMȒ��Mh�3]y_���7q�{).��~�>���Բ�	����Bv%@�m��g�SfW�Mw�. rT��R\��/��gVD�)G�+t�LU��7���A��;>�c먕�5��.A�'�i��a�>�3����=���f2����nD����.Q�B��U����r"��vKS��s(W9�=�S�v8��5����dLG1�/�U����;=��{��������`������j"�3��{U��ֱ����N_���w���=��2�ѯu{I�]��8ֲ5����Hֱv��K�]]1�<��k��}mʞ���e�v��i�S͌�x�۬ۇ��vr�4�d\r7g�ns�.�`�p]��9��nr�K�����<��[|�o+N�Ѣ��=�k�)��mY��)��*��Q.z��P��i��cb�����|�-��ˆ[��ً��Զ��	���1�6��FY5�˃MS��8hҌK��Y��2����UN���q7(�K�����]n����ozu��I�Sw3OG�;��T�q��غ��]����Hd:���Å�dG]\�3���+�F����ʄ��{�׌�:ο����=�@�h���B?�G8
"�^B����f�3<A�i�yp�>�I����\@����|�\��*�j�b�Y�i>���/�ݣP�{o�Z�<��Y��?B�z`�N��
E����n�������-��Q_e�Z�c����y�HJ"�3^��ʄvW]+�g�w��8�7X���r���m�J��sV��;�lkI��5<�n��N����/�O�@�r��r]�.9P�J���Ξ�r�\]�����o$?��=H�|y�9���&��y��:M���uk��i�
7��8eƻ"b�?s�X3�u�3q:Sؤ���Ԇ�C\y{9F��d�}�9��G����S��C�7Dg܇L[P�s��vMm+m��]%�Os��͎���tbpͷ5<��]���c����l��|�aƙ|]��)U�8,t��ʹ��{��x��z�q��%f�"�:v^�y��\�3^.oe�۩3f=x���8����[�Y٦i�j��i����A�Ť�a�g~R����y�Ќ�P։n�ue1��[�����KVj�Q�
�7�ɚJ1'+0�ћ���6���kY��T=�z�ۘ�ݙ��M#zm�c2�;ј�&�ԕ�/�D�XӲ��I�WԠU3u�+�+C75���2���O.��1�_s�|���)����!1u	����麝X��N,'�������)����m6�p��p�pr�6���.S̾V������}�E��<��v���6O9Sƭʩ���]RmF$�k��:Z�X�����6�_Γ��M��*poVsEޫfW0��;�lt8�R[��v�wIQ�����5�C΄�ۂ��Np�&-���ʵ�E���=�0]}tYKN�O/浮��;�5��h  c�r��~�=��5u�V;Ծ�
(%��s�˫��ȕ��+���Q��n��"�_K�k�B��sT9�v�N����Y��É�^}M��h�U��aS�5H�nb�{2ѻ[BV��a�����>S�`vH�
�(e`D��Ջ+��Ӵ��u�{��Gx���I�+Tl�^u<����re�Ÿܦw�t��y���w��w:RP���H�BN�i>�b��#OT�oR��y�sXK��#\��L�ǩ�z����_Bob��k�D)��Ҙߏz^�v�)3Jjs���87���z��ʈK�m�i�a��1
P�����3_*ʪ�j9!�#��쒝�g=����_'�k�i0i7�\dk����fꪃ���('��'�0�s�x����_��ѫN�m���Q&l����t����]-ޘG��K�)�~K*�k��{{4��{���cyV�ga�Y��$)N	��Ӥu<�����!yӡ��"m�IX2�;S�C��	q�o*�W�,I�e��޵�·T=ͨWf�X̢�zt,���ח01Zc~�;��͠8[��L<i�S͌���Y�ٳ��9\�c2ǤT��|�{3T�#�Q/R�v;�u���H9m������Y�u��� qf�����gn`�]����-\l=[|�î|em�'р4J�X��w�^�Lhb���9�g7�{�Q�9Z-N��7p�/>��`�-���Bi�&�f�
�(�����U8=��XܘxDᚶ����'Fk%���Itlf�_;�	b�՜��}:�u��f<�F��7�c]V�t������Q�I�'_D������_Eh?s �=�;L��J�kw��5�����g6��8�=f�[���⾖�@�(�=��#'_[>jM,��ç�l�=M9�z�)�A�Z5c���}o�7-���T�LT�^��LԞ�y��Yٍ�`*��"���q��63�-��.�@.�;�5۩� +$d;��y��[��H?�㻀�Wػ��KJ��I������9�	80�W2k�"��R��}�%k������.i���W����6��I�����djq>��*�LǕ�����F赳W��\4���]ȿ7^'�f�"l�ϕD�^k2�^�ɮS>�;}�s��Q�=��|l�**%�n��+�j�n����rϲ��B_U�5�|��	>T}���~��>�dgz�AJ|J��pvp;�V鸭��ȯV�L���m��~7E>{���>�>����gП���P�y�	�~�p��g/���t<]�3�o-f�W}+�ͨ��_h��� ����ư��w�e]>%�|j�v�}nfΡ��W��Q��i{=���5^ӷ�S'��vg��M�A���װ�y�y�6((n��u���/����T!9���k<�v���òηq3ʫ5YګR씻ay�:��㑽)��u,ϰǛ�Wx��]�W�׼n<q���a�^���%�?�S��ի����(?T�R���D.�}{��.��������{�c{>�F,׊Ue]c��x�B\�zl��'v��e@�#�8gL� {��`V'lW�����{����>��pּy[�p}"���c:�t�,����g�C���H�s��5C����Emߎ��'���O�J��y=���)�<�Z��п�ʑ�<I�B��2��F|��p9��yV�uy{ww��źH=��*zs�'��D{���z�x,�Yh<�u�����yL=��x�H�9��z���?l����t|g����4��"|^�����p�#�Y��. �����q��}/�S�������w��u�W�
Q�����}O���N�q���ۈ�]�j4j�ZA�V��^`�>p@ݣ t� ^Sh)ak�!�z���ӽlv�Ը��*O��m�Y��K'����>�����d��ȈT	�`�OQȢ��p*�������;`��Tǥ�ȃ���D��'Vf��N�M`���-<���%G:��,Gk�l@7n���=�;j�N#{-��d�{vza(r�M���q�У{V����f�T6�]�ո��1�w��t�<jD���V��+2�vU����J�NZS�֣��h�{ޮ ��q;�}2���A}>��_�޸^>��{��[��h�H�_��jM�z�>� 7���@�T��6�x_��S��_V�U�N�����'hi�Z��/�l{��>��q���Wro�S�&���@w�����̔a��%�V4.p����X�7ڧV����E׶����|R��|����Dk�W��z|[���8��t�{�ׁ���s�.��}��@s�mhwS�:.):�{>ަ=g]��ȏ:�ddk�����X)��)�us�����OFG�*pޖN���^�;����T��w!u��x(�^���x��Ts"�}�c��5.~��p�z\2�A�wA��" ��WYU��*e��(��}�ޮ��ok��譂w���������#�m�T䞻������>�ET{�h��l��� �b��ގ�|�R!��o������_��Ͻj�{!{q����邏ġ��Gs�$x绖v��t/`~��S^t�}��w���d��
�������&f��ea�eP��x���W��Xq\溘�jح�ζ�7�qǵy��	���r|E=MSA����H�ֶ
V��V8ż\j�o�P�}C��=��̓ڑk	LN�C�	����q�F�p�n�ty��-�t�RDH{��3��wc���ޭBD,Q���o�ɚ�Q����+ T����yy8���޿C������~w���!ڡ�~ʮS>Ta�Ie�$�|Ą}-�ŗQ>�o8Hr�X;ϫ̯U']~{[��>�]���9f�x�s���7~����L��À�'>�W��
��q���`�n4�YeB���#ZA�h�zv�Ƕ=�C��zHޯ]�6�K��� 54}$O�-�p����O�ss��ݵ���d�.���ƣ_�M���>��OV������eÙ%�U%���A�������w�V�桩�^��GF���f�!Q�ڿI��z|���L��@u�3,����H����hL���8Ӈ��u{����^4."��5�^��/Q�~Wrc�������z�Fn9����3��&�����zx�(Y;���T���"��M\f�i]�c>O�r.1���v庥iI�qtf���Ft�����f��<���d�0��N�>��(�>��Å�^_��^Sg|n��Q��q��33��Г��7�z�x���ۮ����_X�����^j/�ȟ`-����c�+�o)��"n�vL;��a{+@�o��P�*$�Nuqڟ�mrJ$�p��-�֑��
�ƎSǛ��7שY��A���NP��b�z^�w�ҬҖ��>��LՐ>�p�$ػ��qy���|�N5n����8�4k�	/����,T�]m�(��[f���=j�3��W����|��/]AW���ɼ��:v�^����,��uxT
1��]G}�	�}S>�,�A�p*�q숗4�|L��(���%9ǰ�&tZ��:ǀ���ܷ�y]b�)��e]OQ�T��S������ߝ/�����j�{ެf)Q�M)t2�
��6Z��X�=ޛ40��3��b�|��s���dy���=���/z��*7;�i��kU�e���`{���3�YR���OQ�~ �bIH�uׄ�����{ף�������@ӱU	�pVhya�G���c�r!�R�f�g�*�Á'ʡ�Q��ŗq>'.>��\�#�v�ZǺH+�>��Zr���{��i_g���]�z���Ԗ������,�B�P��{V����^���r����ޯZG>����;��*�=�#n�V�ۙ� qP���6:&��v�W�_[{ຸ��`S�oZ�;z�1�M���&�����^22	uo���{��;�EI#{�C��x‧��TFwͫ�c=>V|s�;�_ށ���*����/��R�^<���$eeJI)�7�%��`}���ӵ�TO^�9��'U��x����Op�̽͐Z��V���R�bsU�2�]�+έd6���PyX�)Q�ﯪ�ݞa΃�8�S��yķR6����;#�O� ��r�5��?�t?~q�|W�z��/X��/��n�[5z��4����z'J�K�h5>��79�S�wȖ�@j��ƁP�w ���C�p}����+�j�n=F�W���W�t��z,���5WF�=��~��>�hoz�Aߔ��P��㳁�z�I��Y�-{����g!��+܎#��>μ�Y�~�㑯���z��{"�,Z>ɜ��Q�O���/���6�l������t/p�E:��:\Oޗ�y��=�潦1�Ew���]�^���{��?�۹^���1}n�~�|���M�g���Ф�*�;���W�y�����=�걽��:Ί�T�cc/�_�?$c��ʞ7���wo�3���?�b�kL� yt�}��\�/g���oU���\�OR����޺��9���*xݟ���xj�C�L��΀o8�X;�R�=�ՙ�;،��G2�N���\�C��.ʑ�sĞ5W�DUA�/޴h��ř��������w�ޯi�t���~S��^e���[<	=�,Ny�x=����=S��ml`�K���OEV ��8��/]���9�����/$%ʌM�v�.���^P	�R�+��]�OK��[�Z�J�������`��\�����Po�T�=F��:J�]M���q�78�Osl4���fV1�q�z����$|{k�c�ӆ�ǥ,����12��cZ��Sf��zc<n3/{��iJhV��D�� v���'�V&�Ǖp���ɏ�Q�J�->��V��v�Z����A�/Tv�FQ�q���2����G�3�ҫ�|+�0���i��"�Ot�V"{�L����vCV�2����p�m+�f�n��Y�Ǫv�;�_sD��;�M
�k�aT�7ĳ[y��;�{����$���D�@KkF|�kYn;T$���4��=˲R�&�7+ni�� �o8��iս��8d�g>�N��N!H@fwe�upV��h��5r建%���/����&�7cR�9��vr%!�]lGzqb�yB��fj��tW��t��Z�o��j�Q���3cL��[k�Q%�;��0��R�w��<1Dj��Fs�WDR�̮\z��T�]����1����ђp�[�����i��zզN��C��"�RpY�.=��b���cKe>l_6�q���Z+r�Ȥ���.B8��r�yr�3,7��e�Tw-�*�[Z_o��9Bo%�]*q[���2�v-��s�Bv}z�����]��ʰ[�T�V�7c�Y��]Z�A��c��JƤgV�9!V�@b�̬�3�#���L�<ؒ[#70v6|{B���p��娬�#�}�xnqc��`���Yf�qØ X���ki�S�ڰ��;X�'y�mq
Sõ��*���s��߽�1'�=M9 �զk�G��K�4�ݫ�3����rؖ�-v���3{D�ܷ"����i�VIOgi���Yf�j�>���t��ю�Op���;_J͸*�1m��1#�5S�X�MmnBVE��b�Gv�u�J�8� <�zR�LGG7�B�h���H(��۹;Z:E���R�#A�2\�k�2�N֢�V�M���5�-����,�m��#�0��ݘh۰�0'*�8l)�5v]����u��z�;�J�r�����i�o�5.4z�F�H�ILfoV�i�@����G'_�]�3�޾����xI����[�&�:��cۻ������^��!h���i����k7̹�\ڨ� Z�l�\�N����8���E��E��ɭ��s�Xl��9����R���gm�N�y��`�Bc��1���X�zg@`5��]lü�lDsTcݻ�o")��tq����Ȉu��c�FP�j�p�v!mK��ʜ�G!���3�̎���s6hh�S�t��`Iuݞ��}��e酨"�OFTx�T���;���ٽٖ��n򗯇��>y�Zp�DG:XRO�nK��/"��+�Q���:��%���k�]�#5��'<��AVh�p��%b��)�@�r�n���H�Ӕ�*ĕJ�۔���sr�DFh,�����哺9����I�9Rz�*�-=]S��4�JGH�(]<��U�\�����"�̂��B�]�YsB�J�gKQ1����i��l�QV����㎹�*���'�i�:�0�QrU�(U����ᡵES�AE�\�:���5�p�4s��{���EH���9��MQ	$աX��Q�(u=K�;��F%��TTRZ;�vt��n*	�c�9� ��SD��ʘP�M�9�I&�Z������ܳ��z�驄G����+�[��ݔܝ�/T�&�x��L����z!�YE%Wݸk4r4(�6���j$���G�R�~J��z�Yuڈ����ʟ�ɏM����V����ʿ�c�˛}��I�k�"�	��t��?����r���U2�� N�M��;`��{����wE����pӿqȏ)>/�}����P�G����`���\�D�w��˓�g�*:����W �r�]�zPȵt�s��B�>�0w�z�>D�������g����M��=�������9TA�=0}$Y+�ra-~�8gޯ;c�:���n�g��'1Nm/e�����>����t��K��" 5Qx���z�����
a��d�.<��c"b�٠���!RA�p�ޟS%�xΏp���.'�쉸s>�W �h�������Nѷ^�d���=��]�G���3�Tm��I���R�5�{ :�)�0Q�3�~3/��
�o�����[���7ݽ��z*y����<��c�x���>��^~��W�O�HUƼ8��p�f3J�$G�<5�S�U��t�W+N����^m>6���ϓ���~����O��~���Q�7�w��\��҃%zLyFΏI��N��Ϸ��\g]����vFDk���߇��A��T^,�/k�:��}�ﾟ�[�l�2�	6���9���Q~����w[ U���V6��3��M�Fk]���k5�6JB�h� 5��;�X�Q�P�n�	�[�믔u���=ך%�y)%��	��yb�YQ���6�r��%G�Gb�.E��!����+���st'�;/����d7��"�uGu]Vg
�R�u9�w>��T�I�u9ֵNJ���>���z�r9�ԅ���#.��ۈ3||��Ui����W,u��3/��/k�Q�� {��ȸ��^���TkS�θ,�=�.5NI��(m̼5���w}��g�j����N\x��@q���r�}���z���/n1q���<.�I=\P�m�>�W�S�c�(&�z"�|�/��P>��ޫ w���d��
�z_�����,��b6v�D�n<ڽ�?��>HΚD��e�0�b�R�uץ�E�V%���B��z�܏u����+�_p��Q��+=}�V3,�v�J�,	"@�mO|��'�M�	��F�1������E�Q��;��:U�g��ޯTy�����p8�\M��VdPѭ��(���g���ڑ{�FW�}�W<�Ͻ;^G�ޤ8����������.w�@H�"����萧��_m֥��]�=�ۍ�L�#|�F�~�ω�>�zz�~��>��2K
��6��uʬ���Gj��艮�u=�rJf��pڿI����'����9��i�{� �:���;'.��\}q�{e�v��:�t�'q$ hD�
=�q��Q�8*�q�dX8�~�~<���`�i�"�'/ktl�c�r'�e�R�gY�gP�:�"�ȁ�c=�f�z� ��V��]�w���GS���ƈ����$�#�����/|`��T�4."�+M^�|n��~Wrb���̗���Hb�U�g��9�g�cޗfI���z�L>�>��ތ�>�W�Lu�Wx�O�r/j�^��"�}��~�D���?^
�ʐk�Ī�d���a]z�M�J_-�~,���z�V��o��	�X��R��P��U�ON?uXWs"��s��n�>��"kQ�jԩ���~�kC͉��x�}/��:��3�%��֧��PU��8;7&��9�/	����}p++��{��O�Wн��N����d���@��wȓ=���s���;�Y�|�����6�N�po��YY��&xe	��S�:.*}C�r�\iw�oΗ����{�c�q����K��������Sf��ǣ�*Q���R�,e@3ŋ���7΃/>�4<�}^/������{F-/,K�=�3-��Y�3�G]K��F.ʖn,�'���
�:*e#q]u�.���{Nv���O9����W#H�^A�y��{��u�[㎲�y�L�%�*�qF[)�?x�J��Dy���;5����l������i	@m6�T���ۜ�lU�f��÷�b����P�iPj}s�e�.B�-g%��WIӸ&�=Y�bque��Y-C��҈Cw`�Զ�D�R��ou	�c�;E�}�w)�}zT�7������B���.�H��%8�>��\M��~ӟy����Q�RFt{�~�l�N@���<�w��;�0�	�[�\su�����_��X�9O��o��H���ZT{�t��3޲6�V�ۙ��s��O.n��+�F�l�W�@�ݖ���KF��C���0�;�����i7���IVа���~���fG�2QrH��DL��и�=�O����ۆ��1�z|���9�⼻N��ܫk��o�D�Tl�19Ϥ���^��`��Qآ��j�<�Q0�tF�N�l2��'9����^%��A�h�rB�OP2��}[�(����!"�s���7�˻w9�>����-�3�utq�@�������ۈ�e�(����i��k�{�o��Ǫ�w���]�G���y��^\,��w�5�����O��|��a\���>���Jd�dxsӽ�nf�axl��++�o�U�'��~.>ηq��\״�~���w{�g����}��{�1j��(uL�8�3㳤�[gG��(躕^'qu0*/|�<2%��x�V��P�7�zC��~�uu1��d�%�5�y{�%��CQ���x��dbS��T_���m�;Y�^em@ uu��Ǖ�x!u��Vp�ޑ-CnN��wm�WL\U�H���#��Ve��]��P�Tj� �����f����w�O�����Ə-Q*�{Fo���1q��:m�pfT@�"��Mi��]��}��T����f\���O=�vu=zS+��7��J����:�~��5�����:[�a�nN�%���m-��,v��B�{���"��/ޞ��Sy�z���9HsYR:���O�J�*����.��"߶oW(�%��\e ����y;��9���>�\?)�9���
%����������v�s�+"�_"������{�]TY������}�'��Ͻ�|{<����x���ff�˿b���짘=���ڃ(	�|nPϭ]?�����z�ў}�h���m+��tr)l�����9TVzz�v�(�|T 5����E�J��
XW��Z2#��lMr �C������v��?R�o=�����`�PA�aJ�u���*��r�]�{�{=����d�H���s�J'����_�:G���D�}3�����FD��Q��:b��b���n�[���SڍG�LTm���n=�R�5�{ :�*!�0iM���}�	^U%�0�p���?V�"��Mw1�шۼ��1��fV[D3�SXr؉�"����c��ɡ���1��Z�&���)�m���\6J%@��� y^��#8]�mY��l	2e>Ts9��I��tMB*��ras�EC^ɧ3��] ɕހ�X��n5O��^�c󻓌�%{ޠ;�Pێ�d�ً�w�����l��aǇ�ː����V��
�ͧ����.|���ƿD�K�=>�zv7�+���k�-	D�93��7�c=�}������U�ɏ+Z�O��N��ޖ<�λ���>ۋ�6���^FF�N.�n칧8&�5O���終�����Q;��z'tø��q��]h:��Ҿ\2U]w������8�z'�נ��{�/~����l��2�e��;��xh�T9ɝ4�؍o�{03]�6��{�w哞�� 3�tGJ�/zL�cJ����y�j���|J�/S��~g�3T�k�.�~����n�����O�8�O�����T?��Z�����.5NI�P>/3�w�=��^$עg�A,{"�Z���P._��oh���?K�Y�q�!�n[*��Z��Vf賈�� �X������ϭ��7�~<����������P�Ǹ|����^(�{Q��.��=�2K5�%Q��� x���Yu���Y"0�{=QX|~^|�6/�('�"q\p��w+���L]���K��+�fs����b�����S�So���í���t�`��I�M�De��k���Ĥ�/�z���Vc���`�;�X�Z"b�g��� s��s%\�o�a�W��2f��v�u՝�b��[N9����g��GJ�� t�G�~����L����\M��V%1Mϔ��D��K/f67�]G��q7���2=;^G�=�C��zH��S�̗5�" j@�A���a\��_�׻{����>̀�<��F�n��r=3�}����m���\O��e�K7#���f�g�&���'���N�<qO��"e�𫊟qѸ:_���
����O�|���8�~�:�Կza�&��خ���q���{�!ѹ����D���ZkT�+�${���L_���#gzniy�[���zˮu>���z�c��$��w�d���1Q-m�}��3i��J�
fߙ1�قN��zU䒽#5�s>�z|��ȡQ޺�kg��@Ʌ�'tN�إ/���8�-��y4/}{��kp��
�=y~�^��C�s�Cӳ��V-fT���Y;@�~7v�ݝh�1�<��N<K'��/$}�TϼN����s�ׂ�U�%���)B��~��'$����t�����j$�?�[
R>�ܱ묪�u2�J9��p*��x��,�N}��y�r�Fc�y����ӼST�j����Wt���гX�|���pΤo!��e��8Vw+���
��oK/Wuw�i$F�����ݤI煀8Ө�u���n���b/�[O,�v+X�Is�,���\��J��lW{n���{�$���]�t@�{��H�����rV?T>��ng�*�IrtlT�S�e��:���(R�������Η�~/�+����o�Q�Օ<h2R�2�T<X���7\�2��3C���k2��������.�����R��C��b�ʖo�<TA�~5U1u2�����qᲤ�z�����c�$!���G�3��!����u��υ�f��J�0�L*�su
���#�~�S������]���S}q7��N}�'�{=�G����Dm��]�z����K1Gd�y�u�kև����W���SC�϶cވ�z�9����'_�Dg��U�'��#��uqx�a<��ʀ0�@��?W�P�
Z7��HvD:��c>��[g��Yǽ��������bs�s�;�dZ�#�#ݟ@� ��q�Y�,*[�F�J�c�;s������q��Q��2Ϝ��������m���bf��b��z��E����U1���6�%�B����v�X'�X�{��[������@�������ϲ���n��5�G��3��F��ҿ6��z�SL+���d+��nk�3Q��:9�7r�0��i�FNxp�B� "����5
����A�N�q�w �*�1�vl�7��^�賈Vr�u�W�%ȬL�KM�[ļ4�ER�I���
�Nb�O�G��}ّgZuٷ]X�fs�]�����{���q���߆{ή�?H��_���fFo{.AGĭ�p>7�>]{��o%HO���м��>�]�t���K�yח!�]�ϵ������]xOc�e�G�3�g#:ҭ̃1��/1�P�K'�
>�.|=t{�)��/���F��ηq���tC~����+���Խ��������q��38o�����,~�:�NQ�u*�����w�z�g��|����pU��������od5|�m�ΝE��;�>E���kMԺ� m0y����ʼ�c;�R���V�>�G���0g������"���YS������0���+�H��|��������v����K�5A�`�zȿt�z{}�ǜ�����п�ʑ�x�ą�IF�������ӽ�¿C�qEz\�Ʒw w��}���~��>�>�낁D��"|��u8�ՁټK�M�M{�F�G��9�����q�X���~��'���t���+����ڛ3�/V�ȵ��]�>T_��Y�p@��������t�}^�+����}�h��S�� ��*�o�Z���U`>U�7��ᝡ��աk6���;]�#2��YI�i*0�7�{����<��.�������.cc��5�2����Y�::��9g�A���%:չ�/Sw>�:��y�|B�*ݛ�Ε+"���BB��t�v�x��{����+�y�_( r� z~��.	^S�K
���C�w��6qG�6]��3���Րw�=�޿߽�\M�����>�TN�2Y�D@j�O+��n(�>Іo����nh�חI_c�S�}^���#E������D���d��\ϯ�����27���㍠��[�v��������FF���k�l�CLTjj�%G��@�<k��@u�9�B�s<=1W��	��
�YEy���6}N
�|�E\T��z���\y��IQ�_��~���9��c�CG<���w������������_�Ӄ�R�藳�]�O������O�|c5�+�i��J���	ż��5Ҩ���YGB�6}�J�0Ս���t\Ru�����w�������T^f���nV��N�zw�Aו���fT�҉ݳ0�@��r}Ǫ]h;��Q�̌�=�݋m��� �_�_�O�נ�>�Jp�V9�.�/s*F_Ч��٘xh�T=��q�5L஘�ws��v�>��x��@�`
�ݑr�Kޓ�^�֧"�pY{h_ڧ$��s�Pڏ�A����QS���j�BY�f[6?t���kQ��+��Ы�z>��{̗�S�n�N��^K�r��i�!YZ|�]}2m����+߆��`t1�(Y0]hp��r����0�Y�H���wUUk��
5�.��Y�.Qi�5���N�\텍�W��cL;<���5�����:��Ѣvi�զ��3��q���H���/u����g6�3;�w{�'N7[|��i��"�h��:���Y���w1���l[DS�w�>�9(�[�uA��2�J9������b�/2K�<ٰʈ^e�wA}|t�p;��>�#C:L��U���nN���3��W�����Fɪ-�&��]��V������ɹ�(���Y'4%y8l3�YǄ��PW���\�l�DF���ۜ�O�>�33!Gs��>dUЙ.IF�A��r���ne:Ԙ�F��#������hU�ɴ�VPU�`]ԍ�Nl}�F��G5�)���G�k��!�J�����2�����(ݚ�=�#mW�vdߟv�*�9	An�̍��#��O8\n���1e\��:�G� ]�Qכ9[jH��pv)���Lbɕ;��м|)��H�	�P�\��1�J��.�7�tE��[���7��1@��9M��.�f�e`(�"s	�P�i5'̋�+�7�����h��l�s��r��g%Z�ٛ?s���]0�����Ү,W;��2��E�Kr����BW�N�ó�7#P�JS��kC���*��X�K�{FgN3t���E�$i�X2$v_9��inm��7�d�C�rQ�F�x�qtVc��ʜ��{�Xr�2�2��'%��R����b�[m9��;z�W�Zd�.�kj7���ße98�X���Y��řA*�1���N�7e�)���ngT\.��݆�|�!%M�W�����2���R�0ھ��Z�b�����{z�u�Y�����윑괠�d"j3���m�z��^�x뉴��Sh w@3d�[]֐� j8)a�ì�T�J����z"Ee7,k�=��H�.��VG4���x���/��{�1Flݳ�n�uN�+o,&7��C�_orWo�yF�\)�A��R�l_)pA�7����;���S\\��L���Q�o\�\y���F��yz���U��ִ�$Z�;G�HG�d=���:�n��3��d�r�<�GM[��� �*�`Ђ$M�b5�f�w +JW�FI���Q���Bi�RC�5u�&�f
��9|b�x8��y���M
���V�&�2�
�y�����o��������N���W�>�[}iZ�:O���trv�C�`�t$��7��냞c��d�b�ֵ k;����{�8D�Ƕffoq�A����̈{8'2��̠^�����)��J�d�K)�f=�8RM�;j�Ǵ%�gV�E�\*�11�P���Z�'r��+�ӎ)�Η�J����h����S��J�J"�=i3�\�͉']�<9I����T��)�@�Xy���=-��^���"�ӹ닔Ph������r�y	��ȡR	!3��S:w3��^z��Y�:�ӊ`f��Tj�(�g-��N��(稚�2�z8^��,��+����,�=wn�\�tS ��Ra�+��y���"��$͑*U9�%E��GR�^��s �Ē���P8jy�VhU��<+%�����v�!N��]����G<�۫7ws�s��7Ul����vQ&�w#��s���sw�w#���z9�ҫ�����r�����y�\���:8rT�13w;�h��g��h��E���rr"��t�D�Y̊�����h�";��)�'gT�=���F����"98[��,u%���q+W3Ԍ�]�-nD�N��DTPU
�E

	%Eu0N��צ�a�I�����b�?�=�;�[R�D�R�Ru
j������Ep���sN�/v��!![��+�9�{aʋ�Q�eTzze���@�#��47��o����T?���/n1�;���"��Ə)��\��Rlz"ܒQ>�qS>S\�7�頯ᮘ7h���C��y~��K;&/����'ˏr���=�zk<PVe��� �A���X��HOT�\���X�ޯFs�UHU�óC�������Ǹ9��Y���J�q �H�>�ԫ����K(ھ�^5�����-�A�=���d?uy��Tt���p��~����L��Á?뉝���Y����]>]�<Y���~:��'����y���'=�#z+�lM��� S�nEע@��w98�;����p7 ��G�֌�s~�ω�>�zz�~������g{�)R}���Ü��m��AI;�⤂�(VEK�rK��Tm���oޟ"||Nx�U�cg_�r��ؼ\�[�=�H��=7f��K��q�Zj��O��^�<����{֎��?k��67Y��W-bC\���>��\x=Q�Q��2J�ѓ�O��K[z2��M\f���S	��J=;y#vj��2�$Z����B�Q���޷���vU�'J�{�W�-̖�A�T{W�u�M
��|/3Vo��)�e�}��o��k_Rm���1["�#�X�0� ��aiY� �|����Fv�m�k����3���<��>me���k/z���~^Wr3ޑ��O�=q�B��R}��z�+��B�5�Y�.�V����_�ߠ�����m�W�^�_�������_�x��ǧ�!�����*F^�'``~<��7��=�෻��B�Gz"�s7S+IӐ�_��g[��}��7^�;�������~�"��I��C�{o'�w����&}��
�
�*��ĦJ7��p��yK�^>'b+Ӿ+�u�~�£��u���	}ŋ����:v�e��3�]O�躗C�r�^�p)��X+���MU+�uk�Z��2��޿\og�z�_ڲ��ş��c(���S>Fy�e�2<���5�E�U2y_X�ΐ}`�B��Cr����]!��j�Y�<I�3Ơʦ.�R,��y� Um��}�����F�+���,G������}�����[���8�)��L�%T��j�Oٹغs�.��_�]ĳq�\K�^���'�{#�D{��g���߇��l�V��y^
�.���}^ >�4�Pg�<��G")�\M��i����;��{~_�i�՟�xe���c���)P}�W���~��¼p���Ƚ������i�vt���=�K�[V��(�2D1v�լ(Y�4��t��:���\YL�j��lӮn�m�4��"\O�},���J{+�"6J���k�D��|w����90��k��m&73D�v�����L�ƾPGH���P�
Z7�R���ُ�l�����':8��ޭ��Yj��D�=�pzUS26�f�IX� ��42)�x�B3��+#��w]����{�B���C��޲�G�wĸ��@������bf��c>���7E����r���]���yv��^�+!��w"��x�dxπ�d@wC��>&?���G��E��?(���RT���(�v�3n�W����WF����߽~��9���{.AGĪ���b�g��oFt�=���Ϡ��R�p�l�-E�g^\,��w�>���s�>���ccd�{�՝�ur�f�������ρf�J
4�}����<r7���u��dK���ϛ�Wx�Ć��-e���.�m{�T�;�;��׾6�~3��G�gn&|?T@���*r���U��],{��%w�Ǽw�vٕ��q�;�������6{���H�M��'v�3(O�b�kMԺ�+�LPY�t�v_��(����u�A~^���W�^Dz������VT�>%+�0���Ps�jkE�c߅����ٷ*���f�޾ �%0.��(�{�Yzj�C[�/g�d�^�u:�E3�Z�'Sf�mD������7X�]B��ڛ;��:^�Vf7�55W�w!��5�:��?���=�b�q�����z����Eviͭ,�6�=��ڇw.�˲��7@{�&G�����{���޹c�׭�[h_�eH��O�n��s�`ܬ��U�V��>�9Q��خ�@>7��w;��*=�|^���_�ׂst��N3�y�K��&՟q9�r�%��<�=�2����G~����/;�����O�d�Iλ�~�l�Ť�W�{��c.ˀ�e�!J��r�E��㞿R��!�of�i�?v�vwH�%/;ۧ�{�t���uz�y�P��ʌ��[�"�^S�����GBi�ivv��d�1cgU1�N����R�n3޸<n�~��fK5�T	�bez��>�C��`�^?5�Ow���~P�q�Y#E�7�lg�ԉ�}3���?z����"o�3�FCFzN�)t8{����],�Gx�;7G�{�j��71Q�����z�>�� ;��u�S�`�F���y�gf��y�Y���X�>�
�+�E]O�v�Ʃ|n!/uǱ����_�����@w���~�ŉ*���͌��S�k*�O��S_�:ǧ�*V���*�i񸄯.B~���f'�dg�DI�^�Ȱ6��S!Ff��e?�=�����+��������^��w<f賉d�@x>R�r�����k@h�=+��е�V6�d��)��:C�a��n+љ|:J%��l���x�s4�#>J�ۘ�{�&<K��,�HJ�r����]���ħ���:'c�O���<�YG��͕�Ī0������tJs��l��;	{�=;�c���[n�ł}�Ǿ^���������a]���(��a=�N�9>�'�������T�S���6$��ލ��Q{�~�נ�7^�K^��}]H_ۙR2�O�����=��˿Y��J�B�Ez)�i����Yk�
�ݐW�{�]z�Z�~u�dG���rO}]��Wh{�`�T��+�=��˨S�v�}��|z}�i�x�2�}��q��z���z/a�׳�߷=9Tٞ�Dy�IB邏�(z	��|�."��.n!��W]0o�Yz}���ݚ����.��'�k���z��,�5����5���X<��J�'�}.z۫7�6z�mn.���#(��>,c�,�~w��<c�2K5�<ITe�?�"�>�����][���lQ�y�k�Gi+�5���	���Fy�y��Tt���RM���E�����8�)y
��{�'owNn��>�{����7���n=^X��O���RM�Du׮؛s%�O�׶}�,��B���ťc��⌲,�(U����Bl/B��JV�>ڊ�qˁf��7[��V<b#]�nϴ��mv�-�z�W�/XZ��Έ�]���d��O-!PJ���W:3��v,��⬸�����Ċ�_
��sVލkzĜc�s6�&H�LE��;]Xf���� _� ~��������֍F�~��Dzgx���g~�h��w�
�-^V��Y/�-v��s3�2J�O���"gޤ*��Ѹ:_��&3�m_�߽>D��CuCX�"d>�J�BW*�m����HT}=:faz��.{ƅץi��T��B^�<j5&��<�{h��Q6�;ى�� �I����l��Lditd�B,���L>�>��ތ���MHˌ�ۘ�Z]�w�{��a��������C�7���yX2����&R5ҊF��V�pT���V����н�S��弭��u���U�9�C�s�Cӳ��V/�R2�Y;�-91��գ;Od�~3����wY^F�}�����o:��3�'�����=�W��1��W(f��av$�&��I;�<����Qӣ�YU��Q��R�;�d����g�<{m��3ѣN����+�����7s&t\/Iӷ2�P��*}GE�.����`+����[��8ö���N�㺽�{7�΃=)��z���}�^��g�E���c*�,]L��#��$��}7�I���7ݧU^���lK~� �u^��3}EDr�`���h�.:w��i��t�R�W�V�G�l���}�_n\�t��C{�2�|WR˻�V��O��=���o����d���3>�L��|!�������Ѯ���V��[;1f�_b�$y
�+�"��=LnG�O�g����sX�5s,��$�A�~4eS��J��܏M�v��b�U(K��=�!��z�d{���s�D{���qsr�P.K5�%'{��(���H�&���k�ǡ@�UQ��X��%��o�%˯a�9>s��=��<���z����E�%䋼{d���З� Ց ���W��z���G>��q7�ZG=3�+��N�X��o�������|�U���4��!L��J��=0���g�KF��C�׭��_+5ٞ^�Q�]��yF	��Ϣ�i7��]z��C$���Hj�QW�Ж{�:��Go�R����c�x�X'�^=�e�}��wļ�ꍁ^���m���p&a��=�*_W���:y=gun�No�<����;������\y��>���u�T
Y3(fS����7�4˲q6��HI�{#����n���v�#6��m/m�g��x�@z}��|��q�ːWRt�Ʒg�vN,.�^�Di����n���q�;���˅����~�='=S�:�5�����/��&�
��~�Ϝ�g?��DĊȋ'���J���SF���9ӓ�X�rƧ�M4$��{Y�x�̒�R�4��W�(c�^f<�X�v��8����R�+��z�hW]kv_�X	cS��݇Qo1�ݐ��D��P�Ҳ�4��������9}>�䰬l�wY^qJ��>ޗ�y��=�K���I����N_�og�w8C�y:�=�~��~8�Ḅ|vv�|?T�NIѵ*����������Ҿ���e=X�M�s�`�J�z'Ռ�sC7��F/��ʝ7�wn�ʈ�X����ڱ���'Ϯ����Q�
`Vz��W��[\J��x�W�^z�����Օ<hx���0��͸��{��w��v����.�~��3��� �q���EǺ_�=��<�ԇ�����ʑѶ�Do�ؑ������+�$�#p��;Q�2��.g���z��#�'��{���ׂ�Vw��큗x/-��]�=��d�s����π��C��nb⺨�qIU���~�yI�|su��L�4E��8�-f�Q�G����5�>��f�9���_��
U/�G�ԅk�q�����^5}�>F���=�����Iү=냳�a�,҂*����o��%yNg��bD�u{صl�>�^���p�W����޶;}�\M�px�z�q,��x����c�EP��n�y�"������LV�8ֲgH��D��]�T���su<s�%Fl���K�p���w�F�]o�gצ���+0����^(;e��u2�ҡy��8OU
��8qJ�8�V�vՏ�󝖌����I�E��������S\�ԁ���-���@/Ό����_�����;c#��D����/ޝ���D��g�;�r���oH�ڰ:�{�U����s�9G�'6�x�&�F�j�&��R�����]K�-T���7�7��F���M��fZ7�S����R�v����/uǳ檼q��d�`��*���n�0:��Co��ɨS*F;G�����ױ~��b���w8�۫ġr����g�)��%�1�^��������������q�Ī��\���t]w���jAڵ�Θ߷�����`�}�z��C�{�3�~�ޝ�w�{z,+��9��3	��sL9���V{�6�o�=��G�>��� +�K�^���{�/az�r9�ԅ���#-O��{qS9�
$鼗���=.)[0��eV����X6��7d�^��^�֧�pY�������S�p������IG}�m��1�઎���=R����������L칆�K�iD��Ժ��N6��O���o���9'����z�&P���L�LO9�k�
ƺ`˃W�H���"����#[Y��.qh5a��<)��x�y���I)�wmh�'��Z���,�Fa���5�*2zj-NĎtLu,')w�V�t���n�|��fX��a-b��'�q�Z�vu�U-�3)�aύ�G4��� ��^(�yK�Y�q���=��,�_":+�P��|�p]>��yL��(W��qfS��� �	�o���<�����Q���q���<c�2K5�%��R$&�9�3�Ё��gv��[���{.�}t�p����y���G�*�=H7��~��@�>4ȁ��.R��B��5�U�{�CРz ��&���Ty�~W~�,C#ӵ�{cޤ8��z������3�oپ�ت��:/�`�� ��@0��������h��Ѩ�o��������ǧ�A��[5W�Z���{����~���*O�Q����"���������>B�m�~��*ֻeݺ6��	|�gޙ�����)�2E+�=7f�M��s�4'�a��T�����Њ�t�u��E�|E�#��rb���̛����Q�]>�$�"���d���1R�ތת(B����x��}��Vj���G����w"��zf������ȡQ޺�kg���]:�O{=�F�C��ի��Lo��v�����[�Å�ח�y�{��H���s��~�k2�f�@�����Uq�zZY��~�S�;m}/Y>;���Pw-����u�Gy���2�ڑ�XH�`�a�X���h�չB��մ�2��s�+P�� EXXxY�u6Z��f�s+:nnS�7^��q���eG9;�n^R�zuA�ժ9�T� I��Ė�;fmnƶ�^Ց$N���Uxn�m yo�鈎��k�t�ːu�b.��u�sKU+���u�9I����M)�Yv�:3�v�b�Q��z��G�N�;�ǩ`��⺯���8�F+{7�GZ2���'���v%��n���9�!�7
t�YtCͺ\X�$7z�n��ux�K��9��-k�\l�o��VVV����)�N�m���C:��8��[��xl���������
y\+��L<�Ά�[��R!8b[�
 v���%�w0��KR��w�T�s�;}ʚ�"K���f�M�L0��a���ˆ��n8�l˅��G��Fi�A�v:Q�Ȳ��[K`T��hHp�D+��,��!�t�S�*���% �9z�J��Rt�X��s�L�����ZP�Jա���k�h5%t��ل�WpIXz�|q}4�< ��~*Z�wn9/tܛj[��^�U�[��~EY� ��ג��5�cH�����nӖ�y��>��w���D9lN�ď��V4�30��
���&Д�T�k�*�ȶ"Kv�eu]�	,2���i�JpD��!ls�i兓���b[ZjuNa�}��VX<ת�����q�n��m��(�S!�\�ɬI$q���+2c�}u��F�%�=L�=�eN��*��)(hom�g���������>[�ۮ�H���:PaS���w:�S������|Hf^���ͺ��f�B��__�0�]����̷�s��)؅Ț��\�9Sz�<��3/
w�a/�@���e�<�T^�I@&�e���Ȧ&q��Cº�P�7�;L�);R�]�5@܆���V������BA�� 1�m���v�a*���5�-�������F�,q'y+�I�x�_vl=�Xr$�<|:� �_ju�ju13Cb����
�fu��a�a�2+kK�M��7Ih8j�@��C�3*�ʝ�>�7˨�n��G���!�V5u{Qw�䮘�n�X��*�W�h���ڈ$V!%D��*jmft=;T�We��DN(��e
�M�����*��w�ۊ�.�9�)�/~�7p�����}%��3$����keu'y)	|�rʹ�e�}��Ss$�"VoAm����/�+#	�*�l�A��U��wgz���ɥ���P��:1��t�W��,�nX���m�ײc�B�I���a�#�|,�8�C�mJ���e�LU�0eJfRn��-t����:��b��*����V�)�yNJ
���_[wڲ*�^�ʙI��ݶ��wG?�ia��_T���ȡ@ 丷]Ȋ����<���w=N92��**���pR���E��9�t��1��ܜ�wv^��E䞉�" k�z�H���㻺��{��EFM��*r9�I3/=�Ts<�*�ɚ�wuС�dTzEAS0�.t�4ԮUf��QXe.�U�:g�(���ww.�;�H�5(�EHԸ�^��sR���B<�W����Y��d$*;��h$U!�rq2�[u�i�y�wZ"��8�Y�(��u���Y��ȲueV��@�b������I2�����s�U�
"�;�k����.n%�Y�A8���yz�	Pԅ�v䇆�)UJ�RԠ�n{*;���E��.��:�2i�:��<դ\�8��Z�wY���8NJ�A\��wH�*��Θ���s��EK�f	��� �r1��.z9��PL�̪
��eduKP��=�EL�*	L�"%Dm
/{3[��x�w�@�|��VX�+4W*�Ҏ��)�7�X��Ϙ�B��Q��lSp�5�[��r�ch�XY������J��;����#T��t�.��y���"]W����ü�W�������1����jv�lgj^����9'.#g���+�N�VUq�W�G�����������UFhR�������:J��#���\rϼ9�:�Û2�P�஧�tIr<����M�ZA�a�߲ݷ��	�/SE���l��ڸ��������gĥpe��x��3�q�{%[��iKKڻ�v�(�x���o����S�K������fm沥��Ğ�3�f���4�=�T�����z*gY����<�;ެ
=�}��{��u����9��x.K&���p5�^���}*��<d�0�F}�]�����\K�^��r|��D{��g��Y�v��7�����t��]C�)#�Xn�@H���|\S��z�9��\Um���t������^��6͜��썺U~3ndj�TL���p0���u�C^���>�g��x�}�c���~g}3�M�z��׮�d\C�,ҩ!��u2W�п���]zo{��8(і�V[Wy�	�e/���z��̺=�!�֐m��V(ή�h���ofr�]���gkw�0����N`�|R��yt�2N���P�78H��]+���'f�[+K{��U�Oy���V�� �8�iN���*wIx�qCu�Vcp*�A�\���6r�h�g����������;�^@�F�������3�*�0��'��~�7�������{���W�E[5�Xk村�o��E���>����;����B�O,��`7n�=�=�-<��ϊʃ�;�~��v�6�񴽷��:�7���ޯ�������coTeę�����́��}����7������n������z_m����v��H����9�����Gl�=�%z7ݖ.�L���jO��:�W��R����/��u��n�.��*�޵?d��
�׬����N���z�
�~����\?8�������F!��_�֔�j�͜�Yٛ}�����O�{ dK�g�����1�s:vd�٘y_	�,m��u�	���5::�ay#%HFJ���Eį/g�߫����Cx����g�E��gם�=�r��e�����}�A�Q��g� y����7޲/�/ޞ��Sy�Cñ��dS��^��U�IB.�l�Qr�w�_��d�k�>f�ʨwF|����n#[����{N{����u����_+c=J��\��V+��Ψ*�=ո�껥Z�ڷNB�u��]l�Of��2R�m�V���[q�l��*��m�\�h[����MW��K��;hvi�ן^�%N]-�Xꝣ���fIڥg�*��"��U�������7v����rL�]U���g+��1��V_������I旀C�u�i{ʭ�fr;
�y߸�R����=ѹ;�:ʰ�,4�9��{�|z��+����d`�_8 r�2��
P4��2���Ӟ��'n��͝[�t�>b�]hh����w��\g�pv}T�>�%�P@�_��-������Q7�y���oR��ǯ_���3ӽlv�Ը�����z�[2Y�D��v�m��U����"c�JU�n(��G��Y#E��lx�Q>�8>~�p>�dO�#��*)������{�s���26T�2���/����p�Zbc:W�7���@�<k���/����ޘ�TN���y��_�z��_tۙ�fe���N
�բ�����=�ڏ&����D�7�w7���\3Ӣ|�2}��9ǦFoO�d�)�T��:�zpz�V���*�ͧ�eCs���Z�s�����ni(�'=�^W|c#}�I�@;�?^پ>�8xx�a�d�n��t'�r��d���cᶶ*|��o��gUX���ݑ�k����h�{z,\B̩�zQ;������u�����v��1t���rY��6�bE�4�$���l��6R��!�T�)>:b�v9U���<q����ڑ��Z�
�b��I����q�Ue��ڵQ��� �]��ѻ��-�Ά�q���.��g%���>)����q�3s$��h�ݼ�W�ƹE!�MG��B���|��"]z����z^�U�G<����ʑ�@�q��4Əo�<΋�Y~�U��{^�{�Zn�_�X6��vA^��Iq^�֥�Ύ���U����{G7�7'��xg�^zaO�Q��p<�A��q���|����xߡ�𚛻��x����*���G#�����{q�F���ȓΒ��[K�T��.�&=�Μ��{��o=��OY� ���/Q���C����wYk�Vf賈�e� �.�R
�Qk��vg�r��SssO���tƏG��1��>=o��ݐ]g�{#�Y���J�2��T�L���i,]9ڃtH�����ǗQ.��"�t�z2<���򓇔g�����ǲ���k!8\3wn5�sN� 5�1�'�^$x��:��%}���3ӵ�{~��&��z��˲���N���hz��N���=2ziSPHnx��g�T4oZ5m��9���Ȯ��
�<�����6^)���y_r�ٛs$����OI/ԅ]K�pt�|�Fϴ����1��wG�޿���VZ��� 8�m6"�X�����w����c#r#�xn�h�|�Ou�ĺT44ـX-��8�_^[�u�Ӻd�OtN���@7fu�SJe���u�l��	eG�v��ujdZ��>�Ĵ(���PX�9��A<�H@]wg$.�>rs�d��L��=��Oć�����)T�t#��^]��>+zk�VD�{n�J��۸�l���ʈW��L_�o�d���{�ب��Y�jd�a���a�2_��w�#m��_&�mtr^��r����i]����w"����������<��w���g��^
��6��/������OxǮ�n��/���+��qח��U�9��<f�=V==/�4+���Q�Uc̐����5����s�F���;���#u2��8�_��u��.g�Ks�IC}�5�qg�Fd��k�L�;�;��煼���>N�xg����+*��+ģ�e����w��ўWOFs����.1b�=>�t���j�{���x<���늬��t��2��.����ݏ������콤�H��	�2��t�Y����X�(�YS��ωJ��P�c`�%U��˔+�{R˲\}M���G��7��E����������Yk����f��'�bf:/�=�W{���|gkE�ϙ���	�<yb@�z�{���8�Q�~�=�>u�����2TȲO��ʘ�X�rn�7�^H��<�H�ZӪ�����(��ڸ�B�ǎ��ו+��Xe�mfc8�S	�L��h�=*�N�����L2d6���t/k���Z���:��fpXpP3F������*c�c�BE(�˕�FI:���9Ӧ+�u�("Nz'ʡ�-��.�|e���t��r<���g������p���G�kᜮ*�Fyz퇟d�� SQ%�0��)��ʬ4e�TJ�W�"�P����t�Gk�`�k=����*�=�#o��[3p�Ae@V́���P�
Z+��FD��]�ynb�$�/�]o�<s����=����]z��EÙ,�F����T��������pW����Ǽ3��q��ܬ��m_��+>9��/>�����X>���}��\��F�)A�x�<��M��7���,y4�~Wr<���?���4
�����1)~��
���2\/��eE}=պd6r�6���߆G����c�鿽��}X����yN��є�)����\�]>%P8=����w^��V���y��m����v��T�K��V޽맹]��`)>~�b{!������g/���cgC��إO����Ms#vgdGy�evҿ^(�'}���i����]���P{߫4�h͟#㳷>�·u����?T{���m?�(��A�F;�QA�Vlq�X�Z���X�Ar�(��ð�yE.�L��<��+�e|���0�Z�kq�w&wJ��y]�k�� ��91�,����5mַKz(�W];u<,����D�PH7�R��E��]�Wp�Q֖j���ĶO{}^���#�"]/d�X�743y��b�2�J�͈3>���6��"��*]thz)�q��z�K mxN� �w���W�^z���H\jʞ&�.�ݞ�.�\���xJ���_u
}2����� o�d{���}r�^�Z��O��J�����!�3����v&Id�g��P��3�o��p7��������I�z�{5,FW�w�Z����a�G-�G�����y�6K�<	=S,	U�[��ꢍ�UbP���z����k2-�4�>�}RQ���'ǯ<�dzk<}��,ӂ*���!�>nP�\O� �������W�����W��޶���'J��z���^�f�ʀ-2�
~ڔ_���fNr�k���<[�<Ow�2��Ԇ���2#ӽlw�=���z��_�&�fK=��O{�!g}>t�� Z�&t��Q\}�Cz��������"}�px��N����>Ts����G5[�5z'ޙٚ�F�I��F�;W�p�m�*:�5~�q�z�>T�I�&�x�t�~�
2��e�d��E1��a؟�jS�Lu�tѫ'HzLNr؆pw��X��T{/:݇sq�ÇMYҜ��r�]��m��vB���®����ኲ�sGlb]�SŝW]��o2]��7
����(�j�@�󙙧e�mő��}� o~�����ȅ7� ��Tਗբ�����_��]~y?CE#���c��a������'�oK�2}�H�s#�>ɒ�2�NKcӃ�+N��{^�D�l��t��n�a���y��1�~�����������Y�;�Ī��\@����������˶���֭�>4=�?S'���C��V<:<�ݑ��7�����=ooE�Y�8o�(��BɌ�n9M�>�Y��P��R�h��VW��T��w"5[ U��dK�^��u���^��yu!��(���>���ܨ˛�H�9�wl�v>U�ʭ72�J�LQ�� �J��Ϧ1t����Ց�-�lUo)�}
�X�ѿ����9'��ġ�2���W�n"�\3�������Z����W��\�]�S�k��M�3��W��\odB���rO��$�L��<�ϔ��\�g�_#��=۹��[d�!���^��|V�~��N�ܡ�b7�2��I��~Ȱ%�C��6�6v����Z�/p����rߪ��C�_���7=�|z���{���`�,�3	<�{�P�~ni�eݫLp6d1R�z�� �͈�O\M�M��T�;��㸲.qf4ޢ+�Hm�M�{[�6���x�:lJ�I�疱�1��n��Pc�a��MNm-�5u��[� �Tmk���YЪT��ٛ�O]-[��io�M;{&�b��<��9Ċ==�8��%���p����tG�W�[��*��RMǽ~��L�z��2��2q�l��7�ϡ�v��t	��\M��VdPѽ~W��zv��l{ԇ/	�|��C���^i���g��W�؛�S'Ҁ��@1�끰_fDP�֌�s~����f<DL�<���%�R���g�z�{ՠt���n!̒�B�-M��'��B���F��~2�p�A�5���,W���Z,_��u�7���㞙��s�3,��˞�30�p`���x�
Z��V�zwWF7����>^�<��]ɋ�7�2n��;�F�GO��(2{~0�4�B��]'VǷ��	�[l�����W��j�ͦ:�+�b~����=2�ޟ z��"�w���Y�. \OK��H�,>�W�9�v'tN�إ>��r��u��g�W����C�s�Cӳ�8�����ئ�,W��%��c���E�e���gv��O��^�.��y���>�U�&����ƣ�[٣����j����PUǻs����9t�;e៏�G��%��{�'����-)�J���Ǥ���)�?mm�$"yu^˪}o"�X�r����r��N0���9����+*��	]�R:<{p��.��RǛ�m��愑^}�Rޤ�R��`֟�S��x`��R��2��j���3��ucc鈃��	��^��H����Z�6	�E�}4�gkӾ+>���,�F��L�^��Ib�L�WS�:K�f��������;�LVϾ����ꁰ�s,�M���\od{׬��ʞ7|JVe����@��q��l�8�sk:{�CxX�EL�2܆Z�4<����p�1���O�g޺C�!�b1p�T��c�"YU�V�����V�&�f7H;>S)��b^<ybw�X{���s�D{���c�}��`�>�V�򫙞���f�g�.�ǠI�we���q>7M���:w�>d���;��{���R�Vk�,>�{��n����[ S�X�=��V9O��|�ci�K��U�|Ut��}���;��*�=�#g�L���dT�l���p7�/�������po�RY۾����oW�z}M�q��l�G�{I~�Aވ�]�ȿ�̖iT��t�����kʮcw[��ݽ�懾���܆e�q���ڿ<|��������Tl
�޿\K�TD^��{D3����R���_1=f+�J����^��_.VC	�O��>x�_~����|�z_���cm��0�����ckcm��m��0���8�co�cm���co�c�m��cm����6�q��6�0���cm����6��0����m��0�����`1����co�����)���1P/�9,�������_���0���  Z��� ��kM�l di�#XZյ�0Q�0�
J5"��V(��x��p�MMm�4�cfլ�ڊ+4Z�`�6�U�l�Z�k#FK3 F����Z
jl��u�f�Նl�A��j�նdd�4l��-��L֍��2�BR�mJ'���}���)OJ<v�jO`6�͠wtu:H��ȍ�h�`a�F;� �3kR/��^+Ky��cl�� :���w ���A� Q���� ���  �N�   ������X(9���]6l5f��f� ��=Q���-^����� ;���(��� 7�{�G{�� ;�<��b�r5Y�����7�PQ���E�����<={^c�G{x��Q�s@J��<�(�U����J�ܥQG���J��٭��+J�� ��;׻����M�����wnKl�w����g�z�ҩ�����t:��F�z�4������YVL�SZL�wx �(���+��׶���Z��{�����{D�)�{��%��`=IG{��SA���kk)���@Ѫ�x[kH�ڛf�  r���C�{���C+��z�o��T�6Ѫ���F�ݮ��ݦ5���N��w`���
��I�֙� 7�J�ogp�ݺ�k��[v��@ΰm�i� �a�,���uбܣNi:ٍ͌�Z�� :<
U�����a���j`ug6�U㺙Uݮ�w;�];���H�lԛm��^P��� �gw8
m�0�jQM� ��p�n�F(�P @P%   �xR�Q       ����(� �    )�1��� �     5O��%(d �h�4 A��a�z�4��5&��M#�d��3H$�I���"h���4dLM���p�W�8��N8�6�33���p�X�nTD3�~��Q�� �T�
�����" ��*"�+Ks��|�� �_����_��MD��80#��������ht� �!��!�B����{ L��HV@�H̇�������$�4.	ϗ����;-��<�z����33333)$U$�I*KKRV�I�I%�%Y��L�ͦf�33i�����fk33Y���3��H�I'�q	���8��B i$�� B@�0 q��N2q�I� 4��� d �!�I8� 8�C�@/)�@�I�H�HC�	28��$�$���d q�@8���$�q�Ić!2Bq���I8��	8���I8�I�HC�!8�$�BN$ �@28�C�HI q�*I'$2H`Bq$�Ą0�v�� 8�VBN2 q	� N2 qC�;d�q���J��B�Iq!!�!0�aq �BHq����C��@�I' q��:@�� � �*ZDq��3Y��L�&R\�X�Z���E+I$�H$���36�����&fffd�����ffffI������$�$IrIbIjI$���I$�ĒԒIi$�J�I$�A$�$�Ԗ$�\�I$��I$�I%�%�$�I �K�I$U��I$�I.I1�w�\K"Ӳ�K|ð��K��F���>Ȁ�Y�L���%��B��N��U�5�3�yjJt�#Yڪ�[W.V���;�l����X�]�w)�Ā��F����Ʀ���e�N�]8��m��K�0��Q�Σ̈́wi���B���i�ܯWG��!��h��4�f��nݺ�b�Cn��tbfU��x�L�䭎��E�o(n��řV1o�&Jʐ���k;e�����φ3��o]p[�)2��k��qT�&�g����B�am����-�������4��VV�X1��M�AVX��G�#eX�+e�
�QU�RYuIU�K;Gjo�]Ű-:$U�����b˶m26i���Q�j7#[N���,`����
	��eݡ�i>\��_+�U���HhQ�x��w�ʅ���ړ�V���zL�r[���ն�0�P�3�zW[[�^f0󒫠�im�+XGUmь��i���p6b���l�{kY���ůhb�ʨ��Qլ�@�a�����̗��P���V�X�t����C��ŵaVҳa�ܠ`�f��$��swtd�[;k�Kkt�wB�"��A�P��mn�U���\�L�T��ʽLa�ow�afn���-��rϑ9�k]�v.�C�[�K�����H+ǎlmU�H��]�DV�V��{˝�k�� n��f��!���fQ�U�&�M'uSW��+���uesd��3�ωrmwP�t �iRK��Pz�ކ���&�0��V��M\oH�kq��؅��Z�c*���
M�:E=U�w�^�ګt(��k�A��b�{���锱ز+������NrM�W77v�-I�PaNޤ�l�Ňd;-K���a���շ��6���73/�80����ˤQ�D�\635����9��b���WZQxQ����W���®������eh[��u]�Ҷ�9Ld�^%�K[#4ec�V�>85���8]�D@�w�e�`|�o
�Ed��YPE�x�k�.��ܙ��X�91�v4n�j��Lb�ܘ�ͻ�����S�M�,,�NX�i���;��!��ѵ�6�M��-i�gT;ʭO�=�G*h���ڨ�|�^EAa��V�֜/#���N��vPQ�	ȅ�ͣ���N��V3�*����PHݟ�WA�!%qݝa^�}0Y.L�1��Ņ�Tj�T������W5�:B���ʭfK�Goe�.F�c2�t��h����;B�7��fb�+^)yV�M��G��"�E�Qe3W�(�wyd�(룎��Zn�_�XV���@k3Uє�+5��a�{�EF%^Ht�9T7˧���ͳk�f������sG9� ����=�<=H���nʪYE]�6�#��5O1����P�5c���z��R��$��d�3�l��B)���)��G����X�U���)V`��q�0-嫲�SEW;�]��{���o��o)T�(��ӊ`�	�XMX{X���g�r�e��ك5��X�M}N�����]�������[K�9�d��VXQ��-�L&VMlC��D��E��6�k��{d�<��"�=)�M��V�*`*���-ڱ���F��~Sd�0e��r���n�e�V�:�
�џ'��oi�j��b��I�-�x�VsY<y]�
ַ��u�_�VpPy�V��=�R.��[�W�m�N��.겹b�;}���
�+�B@��}��\��1:E�hq��2��nm^-R���NGA�j��[���d�h��̥p�lm��	�<+4?�Իϴfѽ��ٹ��Ӆ��2�y
ב��n�ci)�]LjD�����q��M��M;��{�$�����)2�A�Y�%gbF��۬�T�mC�o�D��|�eP���^�469i�/�F`�l��ď-�D��V�VW5i޺����	��1��`&�P�f�3v�e��Fn7�|�U`ؾ}m��Z�� ���2i��^vS\����\�A�İ�]��j��d�e�o�]e�8G.T�y���fᗪ���h-e�N�sP����tE�yh�Ȗ���ޝ�eE|(��� ��νֆ����偮V	�U�[i��i��qR}���Uh��;�gq_k�]�f��I�[ch����`�8����*���x�j�<�2���EPя7o⩲*-ۨ戁�9u-[�`eɑҲT�w�e�
V��Өە{7T�����##�6��nc2M�*�e��l����[��\�0^y��/R]�S9�R֖��@�W�ص�����B�^;xwt��d���Q�����ʲ՛�W�)�U�Sˢ�eB`��)1��iq�R���vQ.��x���N*����,j�L,�1]�uh���ǚl�]�Tv��\.+�̛)�N�������Y$�)"�[�Te�����4��ڢ�l*T+j�y0�Ya[q'J��wf�*z��̏"U���7x2��#lY1�2b�u�`J�=Tk;b5�g4��m���m��k��ܬ	uB:�i����P���ݻ�F�7��lC�����(��m���YţP������_,x�1y��I4�����;\��ZC(]�`�O��4�f֫�S ��$Y�Ls	*��K���\���J��n�Μؘ�a�qҳH��8Uj�cV���zZw�&���Ð8;I�.b�����[�d�/d�PbovԦ��|�^a�+Yՙ5���!,�[AfV�gn�ia�XNv��֚yX�"��~�ʩyT��k],�Fk`�����S��[�bw*F8�-TCV�!�ʌi�M�R����Ǌ���V⡍	�a�r쓃05*�4�v@�V_!W�UX�Z�Yl��	��P��2��h�(�Uʽ��7I��ȍ���#QG'2��WV�MJ�Q��ݵ[r�W/lԠ�i7q��A�*kL�t���w*37��0un͚fʖ�2��7Xn�ەp)m���͇�A�m�6��!+6÷Lԧ�6��LIR�Qcj͖u+�]Z�G9>��S��N�Vk{@e�RzQ�2j8���,�.��@�F�T?^��;��]��f=�$H��e�p�%���q�q���l���=*��
�����2ބf�g���Y`�ő��&�Õz�ůvo�$��W��ܬ�FZ��J��t�u�b=�QW�b�
t}c���_r(�\-�r�R$+�Td�I�u��rC�1r�(c6e��+������ȝs��J��c�D�Èh�_nn�d����F\���p+�;�k`��UN�ӌս�Zu/)��z��.��4�Y�i��Sl�Rʅ���iBXÍ֋Z݆q�+���q9�Q�@����N^���95Bd�6�˖#��+��j��ZĿ���n�6�S*��Ȱ��7z�R��M�M1ڍ��$=��EmX��*����e���+�w��f�+�qU8FLa�J�օ���3qڷ:�K�kq�F�f���窳.�s{,붲�$8��!�O}�o*�Z{s6��ky��|R�Uo��Ry��UbD��lk�ǖ�rV��o�k�!���޼:�����:Q�qZx���ͬ�m�k�\,3�!�؈�A��/q>�\u�N��MO;��x���Y�� �T�eң�����T�۵�蠨o���.�Ĺ�O����w�ƽLw>��I�k�5��<���I.�i˲��t'V���kLګJ��2Yt�tX0�]TTfV��[��D��Y���/F	T�.\�+^�9�l5�o-�)�ւ���ۤ��"����a�ues��2^P�h?mjg��ά�i$F��H�H��u<�^�)6m��EUAY�+5��­n9t���G#mf^����cxN��Fj4U�$v¡ zƬ���UO+5�׃���I6�#���ۺB�4dֳ��oX�hh��;�H`����[�mf�e�s.JS��X�V�1f� �b�73[�bXX�	>����[�u���n6����Zϑ�g*�-�u�b�v.�WU�t�"�}#嚫
�/,�a����y��*V�2R����~1�U:A]KۑHB��XKM3n9J�%!M9R�ޠ��q�:�	�Jn��@Z��O�HF}q¤���T0�d��D[R(J�� �J�H�QITI	!Ow�lf4طF<w���Ru�@B�hINj{6���WZd&�.L�	l=Є������T&��T����mu�]e���۶B������f�I^P�۾�u�eH��X
�h�ɼP��W�NF&%��k|&qȭ)�y�I�ة˳�]��d̳����\T1G��\�Fb�q����Fd�ќ�N�Y�,Ԝoh>}#��8��P�9����c�N���qxw�6s��,�UB�qJ9�])��38��)�en��(8l-2��7��al�� �kzi�W8�EL�c����}���'�h�{���)%�]�5�ğ+�(v�Y��"��)_n:��w'�y͖�U�N�pH�6�2�&b	3%^�Y}3[<�����(��eK�R���
�<3��<;j��-E��Xq�<����D�:���p��YjP�Ii�ֻ�#!X}��W��|	,g�oҷu4$Oh����[��{|�9�K��֭=F�3"�3�32sshuj]S�M��A�P.�Y-��`��Gpn��������z�l�i�̝CA)8��o/f!����)�܋Z�noY���ى��Kb���[�M�����2��L=�`d9h�;�mlKJ��h;WD�zFh�i�|5�y.��3X������5r���Ak�,f��k[�QN�͕�.BG]XW��v��	ñ��].�A��um��(���.,۝Y�}ٳ�qjY��%^�1�kk&��B#�f�΅pvV��%D/�KC����"�_(.6����8z��N:��L�o��)����-�l���u���@����݆G��w ��Ä��W�]Qj����[_���L��(��gS.��7v9�:׊Z�'l����'�����+,�j�E>y�R�������B���5����]�Ŋ�%WO����_"9�.N�Ct�e��cM�v̐v��)]�ŹK��/r]��K";;}�T��m�o3���j���R�kǰ��(��b`�ir��4N׮��F��[I�cY�a�ɺ�:�a�G`d��]7Q}vCܜu0�[��U�|[�}!��ζ�˗)�0j�[��F]�۫bYT�Y	j�ivf�#˄5�y���b����WPW:�[>��w���%;�R��L	���0��\3�y�er�]m̝�=��Z)vM/��Dġ�u���4�*�D�Y��Cظ���⪩���nm����}�E�d-���2a��.�uص;���F
uwjEt�n4���b�Η�r�:T/�]�Ue�|9��m����w��I0�bai�3���k5�he�.]H������ e��B�Ҟ��`�X��8��qf\��I"c�a-�W�h��-���h�F��F%��f�jث[�W,�e���᯺�]��X�Ž`PFD��4��S;��F���=�՞���6 ����ǒ���J�\�>��J�Ɔ�Q�vK���u��!���ѡ;*s�+L��K�tz�ޥj�tX�f����ې_\���E^n�ǰ���.ʹ�n��(D��sXzZ�6�j��׷� "9��e�ø�ị�8�6M,��-K;{��-,H�
nD�ѯ]Ke�Z����Ό�w&�+E��!K-8��¬Ύj3��.�	����� `���Uܮ��9��+��44��eK��rB���[m\a�7]8#7U��i�	f�f=
��<0�Jr��,L�9+읷���z��l��nDPV^T�A����Ս�ԖVu��*9��J\8-r��Y*�B�g�h����X��bPMZf������� �GN��o��Ap�.��"�Ѳ�D���j�Qˇ9Vq�8��e���8����c��C��E��
����5�V��:S�(�q�U��^f�gH��W`�%���G�S�//�pxF�cr3���m��[�s���
v����N�!aՏv��)A���L�.	���aZ�v�����y֌��t$I=?�X{�p^��9�&.v{�j��#�k<���+l�N�¸J���;CmZy�A4��8v��������g~nf��
,��w#���z�e�j��l	��P��L����-�eG��b�w5 <w����{�2�U}���- 8��{��L*7�X�p,�P���p]��]��(n�'dPq+UJ�.�{�+�tŎ���'�(�>���UdV�a����KMB��7�۷/�ւ:�d%��qT:�4�٘���mt�NHV�̈��y����.�&�due�}��N�MY����E}������������At�sl�T�eP�y���WoN���D*�ə�c'�4���y/&�;c:��bB�5 F�"@�@8`jM2gl��Z�������k�Ҫ�	�5�ZI��٘*!۶Q��u`��+S��B��U�	�9���XNq�]r,�rŮ����p�&}�C�Q�U�rKhj���[h����Dr�Ȓ��mn�5�#i��jouG"�`�'���}����;����Y Z.,�p�M�ǎ�,�L�4�2���,��`d�\��^�0�r�ѧͩH�I�mwF�r��[\:6\�t�D��y:)�p}�{M��4�u
�\�y����W��K)�Q���M�A3� k�����Z8�9��E1Ɍǡr�/fuѩ�t-m�-�<
�-�"�گ"g����)"=�ח���l��[v�yr��Cq-ƺ����)�W����֫4��F1�m��nT���L%H<�'��ν�5�k�2�>�1r�f��mL�������ٖ�p<�>[��!���T�y�o :�7�y�|��9kM:G�8������wf���a=9�|iM�{+���n3 �a�����έrXz�2��c5f\LI	y#�y�jd"J����z]+�}�8��-[��棱K�C/o�z�PG����ɡjw��H.�P7�z��?B�Yʹ53�[i�8q)bG��K�ur.]>Ot)V�,�	;�!�.y�@�CX�TOn�Enu#�䱳�l�Յ�&3*�/���-h0����s�6�=��`�х��Ys����η��9�Խb�.�h����B�x���陛����\��z��Q^�6a�JQ��/�ɗ��$���9��_
��Q�Va��6t�cM�+�Ŏ�{$V�M��Z��[&KOfY@�ew�2FT��l��]�2`m����9:VQW�U�v����r��VX�һ=���f� �*�����V��NI���(��/`����\a&�e��7&���L��-bm�v^�6�_WcU��e�]f
5���FZ9�6*��2��ZosrIr��J�*����B,
�`�01���r%w���eacWVYZ��kLI�1��*(��3�o�t�t2�x/>=u��b鞧�|kGe�Ի��}z���� E���<��B-���0�[�R[��G5A1:��:��Q������ճ�V�<�Y�&6�
�zVk��ř�{��Ku�%�Z�w�i��(���0H��y���!��Nd�3�����rn=aVP��-]����#�I +XVA{�m�MG]���S�FN=�. ��qM�cހb]2)t*Μ��q�F^L�¶�,��F( ��`�v�ӪA/:!�
ٰS����3Hu��*o�b�d���Ӕ�85���p󚱳]����D)"�Uu��q+��V��#2;�k����02A���r��m�ѹƁ��3���GrRm��E`�]�u�Q�@s��a��9FVm��-�_pN�I�U��{3�K�cM�)�*t�����4����1�l���1t�a��ۋ��ᛈ�fJ�Xk&t!�)�[�Kd�	o�=�e�����G9Q���(+�d�R�A�t���Ng9e��:7��ՙm�-EWR�[҅�V+���K�GS�����o3�,[�����mӉ��2�ݓuR�S{:�`W�sb�}�6i_$pI�0op��[J�쫬|&�������(HsF%��4j]���<�%^�-�*�<�����Q����8�Y�88>Lmp��`�f>�R�����<���2�󔖇sM�������W��YFe3=Ʊө�s�t9�k����1m�܈�(6�[2��3�!@L7�̜ 䦛v�"���C�\�9TPP7�I�l���o�_�b��I��
��YE벙����"Y5NX���[���2��HԪ˩��momͬ-Ң�^5���nq�_%V9�[�2Վu�|yҚ�T���� �K8P�� ��7R�s� AG,�w���w{vE��Vz��U(�TK�7�8�Ò� �aP�ڻ\,2�I�Yy�v�7��<{#莻:.���՜	^sۭ�]��LO�Teެ�H`�m�?�eI�gQe&�ٮ]�5�i��Oy�5(�^��At�9�8v2�Y*���q�8�Y�U΋�]�;h�v���E�|�Au;jTJ�)N�o�M^aQ�mH���v�(⭖n�*��bc�w�'+�݋�T['3�e�e��"�+��U�h�F�#�ywۣA��a5%�]�\�F��꣑�U�45�Ώ��,�ڑʒI$�\�%I$�I�$��*I$�L-&;p�p,NaU������]
��v�T��ӖS���\'/�����3���2�3_�f<a�Gf�Zw��(�u�S1w�E���{)��R=X��mK��.����16�p��u�׌���TR�����rT�첰j3�3Ww3��FI���C�8$�q�T+���7�*o;&b�aS]M�p�A�s�2�e�x���ktb%o�͔3ܬg&���Q!������r���L�T-ʗ�	��Y�J�5F��*i�+���]n�.M"��*�*�X7��7�k3Y��R��E.;��j�wH�2�g6iu��n�+#I� [�'M�Y���F��-4��{����d��	��۴9,�l�1Z�=m� ��EA�X�	��}p�cvY,�Ź�31��knkE	��HL���f��[
�I$�$ I.I$�ʒI$�T�$�$�n����ꀪ�V�]�{wyZyԾ5E�e��&�U:����E'e�@�c\���`cV�ԣ�/��v��N¢�2��:��L@]��7�jn�ԶbT�9��
˨�VP:�0����u8�U�W�Xt�Z��ͩ�u(ө��U\�wshm5�z�ka��2�.�Գ�,��BkF�,����5�ҩ�S�ը�{���J�Ot724���N�����0��E�Ü�ݻ����o|��@=����$�.Õ/��*��E��>�,P�����V�;��3�GXRS�w��{cV�Z7j͘��;
&�!h�f���Z��a׊���������,׹GQ�enn^ÑWv�)+�r����q�Ο:�I�*,ɖpꃕ��M���@C��N&)o�q#��phà��%��(�k����Q\�IrI$�T�$�I$�K�I$r\�I&#Mw\��O"_a���0���eeA&PХ��B�U������K|~��3z4*�]�收��P)�p��o����u¨��g�i�4 ��|^����d�9o����*<�3w��K��:�Ҿ�	é<�is쐪��㽱����ac�o4*�SN^��[f>J#>!��WD�(�u��9��I��M1�:�7�M���;z2�.�#�ХW���֖1��5j�!�z_*�A��m�ݔ"�Y�z�;�+"0�x:�˚��s��i�>��'��w�:�3:/����yV^R]
Ӭ7�w0��tI}�t	�/�I*�R�E�W¢�H�n��-�H��[(��ֻ2����&�̔lm%�)tjt�V+Z���	w���V�ͬ�*k�ܝ$J�E%ɀI$�$��&I$�I2I$}{a�y��ti �b�f�������v�Cv.�|o��%b<��쫦UQ�#}b�)�s��!�����gt^�_\�DG��uи�rI�5R��d�D0�U�ϏnA�(֩���9v��v�Y����v���r�%�8�>yI��mS�j�{t�.���j�l%v���X4�VP�cra�$�F4��&�3Mc���ľqrS��.�2�k���9fW\ӳI��wf���Ck�F�p��l��Ro�^D��h]I�m���e�%��u��M��Fe<H��85힩���գ���˰��-��\�*��YV�B=.t��N3��y�N6ɢ�f���|6�0⬃3��z�eL���Q��y(�C]�W�Z�<�_)�$�$��rC��I�E$��$RI"�L���hv�����.8��]P:j^n4�mguJyڎ켶�'�����
��P�J�lᩏ����*o�*��Bn�ceJ������ؼ����oQsB�4;�Ύ�!3щ�+����nV�����Di���	nfr����P����f�ԛ�jصm��E����j�eJZP���D�������x8�F�rhV���PQ�B����k31	���^;a���;F�:��\�n�֗6�R�J$
����d���#����s�E��w�F����c{X|3*a6r�;fv�]Z�M�e×@� �W0�ӽ�2��+x�����O�̕|ԚɊɵ�g���ȫx�N�Bc�ͫ�b��iVg>T�'�Aً��@�W	�:�>:q�]�$�$�H&C�I$RHd�E$�I$�I��x��+A�n���F�֪��M���م�x�[��`vq"�p�+���5ռYm����X��`�����L�֞���;G�;gr�cC�qy�O�g+*�PŘ���YiF.���۰i�a�׮P��K�o�T@p-�d"�e0���Ў�咁����6]L��Y�������e[M�չ��3�d�ک8�V7vR�&�A��5�J9]�� �
3���T�թ�wG%v�N��pG�E�ui�"���d8T�ɝB�J�+���y�N:�"�J��|�pU��V�I[��k����qړ�M=��M�[Z�7Ӝڪm[
]j�G�Q�@_`�����RGj�˔.��+��U�3I���5�ڼ��'���W7���W�+jV�4�p���{g�dsr�[<��ɉ�;LE�6A$�)$2I��ܒI"�I$�)�I$q�������Ӟu�Hw���E�R�n��X����R�4���y��d�5�����8O��)�����u�� ��5)�GlR$�J�6�)��g�2V��`�XM�Ȭ�J� ��t8�i���Ҥ6�s	%c�UR%N����G�;�w���ū�ؕmoIu���ՍI��h��³��a����������H��t�%V����V�5��6I�[�;m5��٥�o���sLe�b��/�D�<�����٦nV�N���36a�>*Sb��q��IކIs5��[ouᗏ�u�R*�k����ⴵ��w<YYx;|YM�̬ǆ&���g�mw��p�)��:1wȇ�b�������ʴ4��]>6��t�����Ԏ\�I�$�32T�I$r�I#�$�I&�d�YZ![��W�0��u��S;(S��,�e���7	B���@)ݑ,DK��\�]P�K��v������צ��|Cмuk�����um����4���=7r�*巄�4F{1_v^5��',#*H�Pm�e6����4e���j���q�Tĉ�_�ud�.���=Le�w�*�$V�9ơ��!��̾����q�$�^�e��.��L�(ffʲ���2�k{�X+����>�b�\��]�c:-y�u�x(�U�v���`wª��F��W"��a�o�ޗϺ��Βz��z�<�`=d��K{�Zbbõ���a���#P��:�J��|��ЀR�u�-a;�,��Ϯn[��4�N݉�7`˶h<�["vYt���J&yC]���L�ڕM��6㺩�w����2�MT1j+��mXY�%���u,�t)�(;��!L���U��2���6���.t�^|�ݕ�6�b�ʀJ5;Qώ[]q�\�2��l��Ɇ�I�b,�`��+��9�؝�H������F3�ƪ��+6(p-ю�vl�F��
1C�6Rc5A|E���Q]�hٮ�H+[��F�7����vկ��J��9%P"�E�+B=�*U���j}��Z��	|ط�0ƲY�oLWƷ�FҼ��3X�s02��x��i���2VI;v��tk�:�E�k2����޸K�ۭ����a��m�9�l�Q�����v^������=ܘJYq6YK�
�f^_Yѐ�����/�S��Lw�"�,$��i�&3}�lyyX��{�0��z{�֡����r��R�=�\Q����R�42���I�V�֚a�r�U�UDD"F#$W�O���Ԓ����d�_�E"� ��8!�o�_F������H�6*GHjr�a�Hp��1��E��S� ����L�j
6��ޫ2�b��'Bk��[\yD���vSV^aKoL����8\���i����pŬ�T;��&EE�bȕR�d�j�I (��=�t.c��w/!��5��v�kxF�n&�y\���g3F�[sS��0�iwG=[5e �#�iN�E&eߕ
'䥋��r�S�zd�R���5�S��yU����wX�]He���q�[&�'Em�^��}�@d�E���U��2�	-�8k(�Ɲ�b��k�����r�ⵦS�)��U�z�5�݋N��H��u^���8�Em�)���2�6��j$�[��.�����-�·����4�\:�ڇ2�1%����8�\=�6��`��V\N�z�Czq��9c\Tl�p�J���.ղkd��jԚ�u��}s0�̝�X�-m�-��鸮�%EUƙB���{�jΓxUY�q�`�b�\��hU*)�-�������{A{i�[��"F!��"m��`��"�,�Im�]^	?h������?�-�"`�R!3"d`��I'�ub��Qw�`��e�s0�m*�2b��j̴n��}o�y�ְ�eTfF�,$B�A)!2�Ő�qm11*�	��hL��jܪ]S#DQ�Z�E��s7���c[��6���TL�-�ab�"�37��}Ssf4�.fIMY�(im�Q[���!��t�e��Ds0��\t�n�6*��:ˌ������p�Ns~}�Οvk���)dn��m�"�Cv�-��wl������tnE�|�$Ga~�?�����yS�P�˪��*�f*(@��?�m���{���e:�k:���5�1�`%Y���U���eE�p�\�CJ�B7#��=L���^o0�[^K޸=��V�Ne�sJP����\�v�f+�c����l���g�=aTF	�0u�䏆��i�܈CK��F�3�	��Nr7p���{�4������;v�w�lgV�1�$��*�:����	�!�l`��y3Z5�'M���#��6��Y�d�vc3P�`��w�D��ϫ�9�Z��ԬV�1�Y��C4��{�<E0�:幬v�'�O/o5�]Gt&;97U*�lb�j��^Y΢�%M�$��e�=����Fbbed�Gm�p��U6ʬ�������v��b�zj7�@9��X��h��P��D7��|��#�G�����AH3���{o�oP|�u��zb��G	�R|sP��[领D��c"7OmFݢL�@Q��f�&q�*7q�.R�9_^��Cu�������{y�M]���,eh�S=��;��}EG�m���o���}�˓���<���`�,Ah)��0��5=Br�Ϣ���Y��D�.�2Lˍ&7�]������7w5����ǔ�1)(;O��v@lbȮ�L4:7���h��Q�$ά�d���fA��'t��D�0=��4���a֔��Zq��s���-z���VҘ)�ow���v�A����9o~s�����	�6�Z�R�q���X!��o�b��z�Z�9��y�dێ��U�jU�Z���v���s�w�k�P2�*;�W�s�E�`��\�N��5 SچQ���P{dt�D�C���=Jm�o+����Ր�@B:��W�y���L�a��7�zʨâ;�*����١]���w=��2 �v�Tm��#�|[�����+^�����Y�v�X�{D�W��r�e�*S[�#�urS4t�An�3���Uk�h�2���U�eo[.���E��q��e�7MZ;Ӡ�
m�׻m�w3�$�xD�_ jp���8;���ӵY9��^�+t���%*�C���M�zx7T�8�ȑz�NC'@&�H�M5��*���k�S=�(�B;�Oe��&�߯{�=c)����"��8+҅w���0'YK�[?E��Rl��y�*���R�Ꚏ����SՌC��3�5J��d7��*=Ƅm��{;�7���ޝZ����i�T�/ݕ�7ϸ79/��{��O���K��u����f�8nh��	�,o�ɨ9/DV-�`%��A�M�}
Ov������"�~�37�R�$�w)Npz������<�α�
`����6��W�f*�ÁŨe�5̚U:�b+�]�w(�Ӛ;���)�^2�� ��
KT���&��ެ��v��r$8\��=������Z�A��'!9�ت�[ļKV�s�l�q��"MC<��8�4l�C(jU�����aH93�ɇ�o(��L�q��W#�U��}q9,�]�"�u�v���q���vw>ae9����ڐ��Df��=&�w�

�E���=]@�r�Aa�����{9�������]OQ[v��E��w�μ1j�E!��%�Zt�	(�R�2�p�|q�SUq�̕��/��M��/�h万>:��[�oqT��K�R�̒�y܇�@�vea;Z��D�X���|�Is�)"s59 {1 \�.Bg`^Ak�=�%-���^A�7=~��m��5�-���d������Y#V���Xts�i$�n�l�K��.�nTUKtt�=$#޴LKI�{'�i�
�]�<횷Q|"��.�h�_qzZξ���;:r@5�#Dn�"�p[��Zw�.f������Jz�"�N�����7�b�|��N,��qo\�e�e� �;Ҏ���h��Q{|y�yq0ە|G^���n�T�'{�8���䫶�N�pq{I���W�v�׎��e�P�.����a|�5��h�5���F9l��q�Rkr�<�����\��ޗ@�����Ȝ��ާ��[�6q��o��bs������3��F��1�3w���k=F��bFd3�9ɵ�Q[C�<�q��Y�9X��:E�T!T�	#:'�O2���ٹc8�����x��jtc�]�Y,�s+%?�7�f��k~|"ŝ�;5�&u �-OLط�N��2����"�4�K��$�d"�R��Fdո윅5�d%\Ț��ҫM<,U � ^+����+�A1f�oB��b��=��γs_�Gֽ��t��~��
|�q���X�e���_G�T�VX�����NoF�W���B�[�:��GE���z9��2k$�
�P�v���fqj�nj��7	�VD�{�6$s�7ǟ��{.�[j�r�Ή������H�Y[F���35B�s�aT���TpP�-��8D�"��e5��ݛ�c��p��f������B�,�e�!,��Ig}��D.y�ņ���K(휊�J��l���:)ֆ`m�gg��[��k��ӝ�`*o��{tўG�.0��ݕ5V��3/�A�o���<��N��v�U���_u��ܗ#;�G+���rpa�t4��͑o#�{+�Mj��D��i�tc^Bu�EG�!����$��p��2����a�U!�K�I��e��Wnüף�N�� �fN�,�'wXę\�n+�ܜZ��E9:�������B�`�j��W6�֋ʩ�5�lbH�[�&y����MƫRՅ&��M'��8���eA�qA�՗��7�n������V����h\#�`�O.�BӁ���%F_)�U͵�<r��5n�z�V�1;���\�)�J5y!E�l���Ie���;�m} ��u
k���7��u���h�T4���vO�����+�~pn�\<�����j�D|���Zc�P�%��s\��.�.�~�mf��͆��K~����鴋�J�PD�'E^�٤G�U]��v8��W&?��-A�2$�]%W�1x���v��w�vG8n�{��D�BF��`i�[������q4���W����,$uc���>��=^���CE�#���{�v�Ø�1�����v�5��.��g]^�v[U�2�A[ת�jx���Xr���"9:T�r7h`#�݉6O���^���8������=�a�NYR��#��5�>W�*��XV��>E>S��pr�r1N�����=|�P"3�u�=��ޒ^�dy>�a�x�A�o���z5��B�i�jW�!��Y�GE�Op�uD�:�����"q�Z&��/{��/����?` �j
d/e����z��j�3���\."�(��.�	K������Y�EZ�1ݮmv�2�Ou΄����j�!��;�]��%vl�a�dA�5�N�X�^]D���J�fc׏�V��J�3-�5�:k���,���(S�u#�w=���:�%�&H�԰'�!�ء�F��k��z�a��‱	1w���TٲM�V�=��f��W=��c/k�;�ѹxh�2:���LV@cV�=��I��e����4�\��
���x�R�Yt�k�����0![��+��z\��5��9yhЗ��2�*�:ؔ��d���,��=�D��(jǖ�:�e���Fgnr+��g��sil[S	ދ�;���捦D�M�X��Hb��p��*;��vp8S:���ɋ���C�e��\@�1c{G�~��{���cǍ���{��r�����8�W%��:g�]�ل��gk�,¢̷OBOdY��8�]�[*2���=�B��c��d�0:�e�eL�m��F�(�>����2fѥ�Uz_7ϩ_s?2f$/�2b���7� �X�Cn4��9`�N��:�	�Iüd�V[��]�����2&��zu�Q��Y���8XGB�YW��I���,�}�v�Zz��}`Jx��V�ۣ�]�7��)e�KJQ�-A��
��T�3�M*����1��)��M�pfC�٩`xpK�)�1<���0i�bL	�sE�T&���uj	��_E����f��_p1U�����g$�W��\[��.�c�0��j:ُw"����z�]w��C%�8�Ǯ�)z�)
zOm+|�b*�mKlQKlG��_��g�o��j0`��T��wq�"�(��Z��)�V8ե�����t�n�A[kE+��h��L�E�-[^����4�KS�X���(������X�m������i�-���DUDV(l�T��6,�6浧Vip�Kr�{��UgU���(8�u�u�[f	�LJ��-�5[F��{���"�JbQ.�:�`�c�pT�`�ƪ���֙l�o{��:��mfebm����&+1�h1SV�U1̵m+c�q��{�m�1�a�X\m�+i	m��q��S�6@q���J�V[LLKF��35���o�Jn�RD�h/�a�H��� &da� ?gh�$'k0��ua��O���O
�.v�B1xQ;�%Y�.>�\d�i��� AzK	�~>W����F�n�����ل��1�}��>��$�y?v�$ �^��0t_��^O�Y����=�?6��>:]B��qյ"�٫O��x?�������g_�u}��T�k�H�*+<���1v>���}��]������g�*��r�Wz3M��y�3y�ח��/QB��VWnE��1:L����_����[�y�{�c��8���-�6/[�`k�|ҍ�U�z���e����4z�\���*�y�K�(��o@��LS�=4V縁2b���\���C�Z��
r��ͮ�N�?���Cx,�w�l��]�B�l^�����s��e�՜0���r��g.�e�5�#N_q�-��)i-��>X��Uh�d�������_�;���o��_D�q�[�9��/+���/���i`Ǥ_��r�����s/�f�A�č�~o�;Þ��)�	�����d|'�ێ�����{�ù�q������
G5k��R��=���Ltt&"�N����5(�)b]gޘXPJ��Vs��P�1u���Q�]�7��l�-'��\X�b����o��T`��U<��#ފ�J��ؾ��w����yTy�x��=�s�a���u
��<,'˔_	��P�󡿿,Q�o32u6V���8#�Uwz�YU���kf�2C'��`�jkVƞuS�Oj�oz����>��h�Y�袹G��ެ����
tp��r��Rq�,���o��`l3ftj��������2��hf��=�E�b�l�W�]M�u�W
ofv�w�K�m��0y����� *�1��}|ϛ��BQ������վ"J�]���^�Ȉ��c0�-BS�gt�x��K^и�w�,/���a�����G��B��#[�km�<�K����<�?r���а���{��M��q�cҢ��`X`E�a���ze�uF�  ��T�Hr���J��zNF�o���%~��O��^	m��ޘ����c�|ʊ��U��`k72��#4XV�W�����Cm�u�a����^�rk��ȗ7��]�N�bלVn���^�g�n�q���\����![�i��O����d��OF`�B��w}�޸���g��!��-�D6�J��)>����5~����D��F���Ћ7g�3 jf����!���:,�x��aa����ͯ�3$���=H��]kY����|��2CǤ���t�x���u��@�;C�!��!ެ�z�G�Y'j�w�~����]��s��,���l=@����I.�wd�h�q�j�=0������ ��9�ֺ�_��uםk���x|��Y�y`��I����v�\�>I<�Ȳg��vɴ�N2MP���{7���{��y�yϾ!�����C�SI�'��ԇ�$�2u��$/�J��<�̑d큖�ē��e������;������Ԛ���4��io�O�i�L���OX
���1��~�J�ꘈ�/}b��?����Xq 険C�&��1 t�����������6�ӌ	��<a0偦N�7������z�t:�ÿx�q�q�U��L�N�.�;]Ӻ��0��b.u��%f�3�ԩ~�05��fc����L轢�[�
�.��7�����Fs��D%���-���:c�5��}�$�AH'���!�&j�2z��=Bt�8�'v�4������uT�6}>�4ɏE��)��) ���&��N��3T'I�CV���{@��22z�x�S�P�c�?EZ�RϘp� �}�~�#��~��$�S��2|���ORN�f�	��'��I��6����!�������}�]=k]}�|M���ydXa�<}I<a�x�䓦$4�O6�8�m!�hm� �v��@8������>ϯ��~��C���t�X�=d:5Bv��S��@��l':�@���8�q<a8�yl�!�=�n\}�k�u����i�>��3vLd�5��� z���;H0��I�&�@��	��I�z���e��8�fEm5��=3����F��&V�6�D�i<O!Xx���,2v���Hz�q��Hl��'�<<�����{�x|I�c'�t!�3��h����!�"�w�ĝ05J�x�֤�!��;I���Щ$��|��޻��}���ǉ'HwI�i���N�C�I���]ӌ*Ad��'��2v�=�����s�������s���OXl<I�	��R�z�r�x��$� ��;��
�gvN2z�ީ�C�l϶>�R�Z��Z�YWK�J�᫺������i%�Y�)��;
��,���C;wY��%��Pڋ��ڋQ�s�͍�@ې�giEm�D��6RNb2c��~�PE��Ψ�a��z�|Ƕ�BX(z�z��6��;I�Y!z�,�> u�s��w���=�OY;d�*�'Ƭ��@�t'>�+0��$8�����I�)'�0ea��3=���}ϻ�u�d�I'��Y�`al!���OYC��9���4ΐ:�@��N�<d�3t�d���x�Ru�;�ξכ��p�I!�'{�W�I��$��V�������S��$�'Gt�a�':7��C����k�������߯{��sߎ$C�P���9`t��&��$�u̒��&�,'O� m>M�d8�i��:�Y6����k��ϗ��_}�<��x�T&&�s)�!���ORu偶O5�t���N��a�I�-��%OY �������>�߻Ci }9Bx��	�N!�
�;7OP=}a>x��O�=I}���'I�,&3�VC�i��=r���]_u�}����B͠i$ǈz�>ꓴ�`,� x����m;d���尞&�$�VN ���ξ�u��s�C�<gl��$������1��!��'��Ĝa�L�=C�y��;N2v�|u�I:}I�^���s������
�O�N2l�$�R��AOY�Y*I�P�� V�O���'?R�����z�Qc��x=RVu�`�h��	B^jU���9gr�����M���-ڴt4�e������5_��KE%�(�c+)Л*�N�� +���BI�C�Ww��\Dl��O��2aՇ̓i��Jn�P��XN0I���Y1 P���AC�$��5�_|������{��C�/o�'�1��	��I�kVO�C��!�&<B���05)a�>d��}��f������}����1�
��$�<BY;OXO�@1�=I=C~�!�"�Y3t�z��o�5�}����O:O�2�������d5�=@:}C�,�ߍ>Bz���0�������z:�}R���Ϲ�IP�a6ɷ8Ì�N����z���hN��u���bT�׾d=Hzμ�Y9y���u�Z����{���6�M� VO8��y�L&j���O����	�_Jʇ̐�ꞡ<Hr��n�־~}�:���C�Y��$>��$=ݑd��yBzO2Շ�Y<Bu=�6�!;~`
_�ϧ5�+��w���v�2�ORM2}��a��2b@���$�PwH�m��È�S�Ho)��	Ğ��������3�����|~��}�I�z�\�������z�I�I�$���I�'9d�'��'N���)�>�zy�z�y���k�x�H�q�=n�>a�YL�vx�Y��=}I��<I�Hi�ޜI<G���z�MNos��ؿZ^�{o��9.ig ��l�f�g�v��3��»�]�e���~S��E]��l�R�+_侱ڨ��'GH�DQ�����G����SM�t���'S���=d8�״��!�v�a�Pā���L���d��ԛ�����/5��w���/��`zrȠ��MHm;Hn�� S=�8�f����5Ր�v�SGV���ԁ��=d��	��ѷ���׾s��:d�'l�Oi!�v�B|�J�RH��w��I���9�y|�s�@��Ƨ�ww�3�o�y��ol��S�OXM���{d���6����]��;��՘����&����Ż�sv@Zw���Oe^��?=u�I���Я|����L� Ӭ��+���s�&~��>�J�1�Ư��#���<��^H̵~����zӍ�^۩%��~�p�*w�tB��b��V	K�Y�B��6���+F3Y�R��t^pl��hd+67��]�v��s�}�կ�X:e����7�+-��n���yq����]��y�n�Ύ�ߊM�GQ^E`�.����y��M8�%��)+�����sq)�'����s�Ԛ�|l�^�*����u�P�lvc��{�O1�3�c�T(��pLP�X$��v֨z��c��Eȶ)���Z��qـ�����W�U��|��q��%��^�Ʊ���p�f��H�2��֎��I�Oc���lQ��1���v�)4��&��M:�9x�z)V����{������3���p�l"����w<m��}'31�^0�\^H	�@.�oO��He���g*l�L'ݷ|��__&�6���xj�M��٩���Ȩ�;�s��B���Z��B́ݚ�5[\��L:�W]��Xzn�-$�9���:�K�ܗ��F��T�;��b��4�m�,L���ɴt����73Na(Db�Y܊q�33?L��L���x{�=�*M�\��޵4ҍ!�
��E���jon�*k�D^p��EI�}{q�C6��]��13ѭ^�V~yI�5r��0/dm�I{���X�Ĝ=�T�f':k��.��
���a���3r�1� ��LU�H����k/ޮhBm�~�x�rN#q�P �P����^/��0 U�yl;�#j���j�ꌠ�|�a�ў�wٷ�c@Q�n�n�*��%0����P�2��N��U�nxI������h5�[����b򻹪�vH�}Q1�����w}أ��fͬ�P���+Mv�ݬa�� �*�*�r�ӢГc�XTR��#��.��S�J)ege\\�d�+�c��P�i�ڱ��Y�)�g�E)���na}i&�^nV��|�Y/��"D�Θ�
ݐ�F�И���v�eCW��e��±�3��X�%�T��٣ya��§-�N��@�
���F���(�D:��2�r"�'OV��L�Es�Tڽ߲ƭ]x-��r��1,���%�苿��[��^�]�TGщVR���p�t�`�sz�6k��]��'�$�Y�f�l;]u9*�Y�����EJ��d�N(V��{�#��9�2���ƭ:�8 ���<�ėj�z��/��Y��xY��n���wx���4��jua�l���5c.g����)��Tb$��q���\�	]�u��Yl��Q[h��Y $�(%Ie��%�!
��K$�A�����Hx~3õ�/�_�D�����;�UfPe���sH�RA1S�Y���5�]��s�̑\��/SxJ�I�n�ꩯz0�aMڦ�tC{�����:�qg�D�ɸB�t�WT��/V����B\lf�MqӮ��m�a���n|�Ž�nyLJ&I��7E�+ڸԭ�.��u4e�J��%(H-v� ��jH��Sp�a]ҵ�!�c?��p��B��k%�Ng�����e���,r��H�X�͗�	$(-�\��4���;+���v�o&&��\�71Y<�Emc|ɱ+�g�e�5B����]�ϩ��t�U�S%k^�g�s#Ğ`���=� =�_{Ė�	�w]�`O��Q�qw)���Z��dǪ5|�S\�'&�."v5j1+S%�ԝ�gbN�%~U/��W��n��-�q���0Lieq��Ut�!r���1�Z�.k3Y���b�ծ)���5K��5�ulV�3M&[.X�up�Z����������l�`�ٳH(� �LbF�[Ks�Q����0jP�r�[`ҫW7���+z�ް�Q`�1.e����-32,MYDQƍ��{ڳ��jc��e,Q�L��+0W-�)��
���c[�����Z�R�X�`�6�֌-,���T1�s+���������z�t�(R٦�ի���J6殅������(������n��
�n�WI���4㖕�5�ub��u�"ĩ��R�ﭯY���bR��+��0-\�,]9�\�8��Tˬ�n8�%Z�F�3)���պr&���V�-�>dyX�Z�	�A��nk�����u�g���F�2.�R���7�|�ε����]o����>b���,,��6W�=��ng7����gܪz5�����+P����%�+�9�^�Q�˭�q�Y�Xz��Pf�6s��z(E>w��̓�ػ4��!�C�X3S�M?5�����u�R��W��>2Fΐ^��&�z��������$�n��o*����F��Ž����J9�{��&�FF����y�r>pcW�"�ygo$�F�s}���	E��۹'�H��w�5w�qˌ�um�]�%"�og�<Pb��~��H�u �)ġ��W���I�mk�^�¯aC
"�I���1�y��w0���R�:���#Y���pw23#��Sx�^�:�=6�;��:��f�C�A$�H$��~�!��4���uهS1�n6�fV�[�Q���A���
3���Ѱ)�B6]�)h����U��/�dz�ZR&Wӹ�s����<�=uy{�i�\�|fI9�e�R��^�qX�V�O+H�k��'Tr�I�9pq�Ef���p+���mz�X�ÄN�7<JgKgg���h+�.*�55!ݬ���ˬY��#���#��`N3��+ x��%p��A�q���zo�*x��� \��Ai�쿮��=/c����[^�a��\^�g�ז�\p���eᙻ���'����e;�<���"�o�){�����گjh�n�����=���&�4���e&ښ;���w�?� �
AdE�}��7��?���a��wf���]r9}y�ں�(�Iƶ׭��KҺ0z���Lcޫw-T���ށ�T�*�l5��0�%֋I'5_�7bLN������+x12p�殭hmKP� -���:��\���dǅ�׊+�Z��la���:M���1�z�vˍ��q��^�wo%�:򍃏Ʒ�f�v����i�9�q"J5u��n#q��ǅ1�䃂i��Y�.9�<�4;��p��}cH�h��U��$:�N^8�S�������t���OF}&Z�oJ�[zU} �5x����Rb�Pn�[�p�j�y�{}ɋ����c:��;xT��ؒ�h�R"��Zz�ߙ��m��/]y�<��!�Y"�AIH� �ߺ�=�ߓ�5�}s�5���7�� �Trv,���'7�>�����;��ȯe`=G�'n��[y7�owW�}�'OV�[�n��C{�0�g�i��
^l)tE[�τ#���CU��ȝ���c�q\�c����b����ꋌ��k�v�l��;��s�S�0դ[l���Q�i�k����ۼ���d��W/aW؀�G���B�Ε��tf<����x��¦�o����4��w�Wq�Uz�ٙ��5�V���'���2P˨�Eͮ9`Q3�sa6Huu3&���ML-! ��/fZ=��}�=1^�o���TX��ɳ�����Û��ߛ����]o�<��!��A`,��3��L�Dm��{;�vb��ç�΃SV�0>u�q���"��խ�Pp?gFQ��J�͹�Y�C����+e'�7G�
M����$[ߤpf�x���;�E����)U|��ۜ�鵕�1V��ͳ�m�Y���1�o�����t��>�̻��q�]�Q��`�_���9d<�=�/FI�n�}��,�w᱊SI�$s%�M�<|�L`Y$\Ez�R����i����p%Z��cx��f�Nܚ��.:�����2��.A]�٠�[{m�۬^��a�����v<E�����u�R$����X�]�
cW�奸���W��Q�\�hD�˷K�V�"Ih��c3n5�oEn�T�1w�������?I��R,"�RE�)~��_���_��M�Эt��.��ۊ�r}�/�ݱ�B����jrsK�6�+��:�%R����v�&�7[S#,1�d�Gf�[I��U?5��i�FY~�.�^���[[����a�@�_UE`덍}7�7��oWF���i�Q`O �*o�[?����L�g^�qE�'�ɥ���"����ʉ�x��o�F{��3q���֘�,5��˭�ۯx9DC��|���%v�S�HP|Uۼ���A�4�ޭ��me�Z�f�ߘ����7�'T�@�ʅ�Z��yGD����Fʙ�ʹ��Zm6�"��>��{�(,�ίqit[�i�=&�/gm���� ��>$| D�XE���޼��~����s����7 O蒸�7aF��]�unv%̗��Q�OFØb2p>�����f��"��dW ���:��=uј8�9Ѭ�L�{���3�t�G��(�Ntz�+�$��=�ip��nz(u�Ε<�˻��w�TK���\o9TI��ܳ��˹�Un��3�8]�q8f7�+�����H�KoH�1��K��E�*������u�]�uD�ڧd���=��5�^�8�$T]l�NQC��d����u;{��+��`�ͺF����>�^Β�~H�Lw{Y y�m�wޢE�3w(��6�Fty�o��x�/�1hzm�7��5h�_����;Os�}�sίZ��7ם�����I�A`E (Aa	}��}����?��~�{՞�Zp�y�Od�{p#q҅(��c����yq)3YX��V�gs��Kp&��`h�S�����Ʋ�׵�~�ö
@&zi��J	kk#1�*z���l��Z]��/y��K!�i_l�
���^b�����X�қXq��\�X�<�%;�_�k���f���mX��G�M	|AaĮq��U��n^���Y�/=v;��bo]�Sy�1���k>�:�LZӠ�N{o�Tb�
��˦)�ߣ�wx;��ə�E�q���͂ꆗ�(T[b�kF��Z`A��d;k5�"K�W}�(fa��;�ivVL�N\Ff��wC�ZZ
U�]7�-jK���/�}_� �"�� �"��E�D�>��������y���]Ѧ���1Q����I���f�&q�l3�Y_�/N�{<�ϱ��؞[���܃X%�<���5Kz�]��$�N,�,�A�*��N�Lй�A^d����$8"X��t8��j�q�����9��K��J�X'�N�@K�����P�Ȟd���}<�⿏(�Xuh��w �qtN��N;Q�74"��n>�"�/��}M����������,�obĸ�
r��7�����.D���۸�pa�ܗ��;цcw�}W��&)�|,���z��yk��R���X|̢u��I�J��r�=ys�lg��V����v���+j��a�5���g��o�{5ɯ��޷��矤'�$Pa"��H,�R �@<��}��|9��M�=���<��;�7�,�<.�/}�?��l>11��;'�_we�9�	<H�0���3�p���ee���P�O�{{6�_t����(�����Bap~���G1Y��G3M�j� ���=ڑ�s�2U��5reN�iR��J�g����{Ӗ�]71���J���򼍬���J����(0���k1�w:�.��C���H��k{�k�xr"J&�&���U�*p!'����!ŧ��R��n��Q�Ѿ�<#�"K��W��~�~'~��&ughk�nd�ˬ��o)w	�Jv�^��F���ٸ������#|{$Y�q9p�Vu���[E�4gՓ5�Y=*��՛��ujP�97�^���	Y��i��R`M�l��0�&��@���̛��Su�t2��w�ntbY����p�8y��j=��W��[vJFU��R<VӉ��QJ�]=��G�I�U��PU���93qX�w�j�SWGJ#M�g�2"��;��xY������c�5�����6���S$�x�Z�K8��c5�RV���t�t{r�Z+����x	�����T��9{����w�h�RVҤ*ʼѫ<ԋ�)�5j��Vx��Bdy�Jc��}R��sB'K�ZyK\.��u���3*��t�ŧ��D�Y�"XN�Έ�J�]�f���Vp�h�Qs�X6�\��*X�;NRM�7��^��c�SCf9�]nn�����m������}��Z��%K|�rj�E�'9`�I�y��|f�Lڽ�/m^N�&4�v�E�����1%Ƴ�Hn��mᙏH��8�s��}Z�YGD�Cswy�6]�N�;��v����*ZeT��)��n/N�b�&��ͯ���h�G7�l��鮮�U��Opj�J��+V'n�j�]vN�l���'�Xp������4|u�Z�U�f���4�J�[6�C:��3�G��/v�;��B�R��1��$�q�g0w.h���`AK�>�2�����L�u¶9
�U�x::�Se�z�8�ۆiQ��k�%��%Қ�J{w\�Q�pK�\��樻O-��\�����q�̬R�2����8�3[��k`f��9�..��pNS:�z/Kţ�����8,Ă���Z�+QALuq�+SV������D���ۦ���Z�i���$HQd��LF�H"�޷��-��ʩ�FT�0�8�:eQ�f�KTMe���Z޷��V�4�ULݹB�L�0P\�!�
� �4I$��.���1��kmT�c6�WF�&�.�M7H���q���o���`cc�GV�ZUcD���̺\��#�����ۖ�fC2��ى�	D�qYR��8\��[Es[���Ve�6��GH��̀�`��P�bI	�s7��ٻ4�w���Dm��(ն���+-,s0r��e4�Y�QuV\��,���M�wcԻ������#_n�ֻ�?�cvS�Ǵ`�:ʝI٦(-��U��$H) ��E���'���"��V��
�Mtp�H��f7u���sAo&�/_�&�T^Z�1����䏫>�~ӝ@��Q���Y*�~��^W�W��]i��܅�Ln�#yO�b�\���sDT*s.�y��!�"�@B8�D�M��t��Z{�Y5xg�y������]��[�|7��;v|���|��a�3�W�X�W�\	8�̈́X�6�5�1Y���/E�7�6�2�jFh�V�LmU����c�B���t4҂�K*�������$�g�#}^=}��_h�� �qs���jx2��,���7���&%ȻY�����&Z�����4ȯ�#�Ǘ7S��ie'WlJ��H��n��矤��B$�B,�,�����!�}���)~���$NGL]���٘Ѩ �q?��"m�
23s�N'UQUQ���M^�Z{ԭC��%I[��qϱ��q��'vC�~�{q�:�<akT��p8���5Μ�+�;/,�����F�a�I�d��v�^�X�J�ɨ�G+vbs����\Y�c9�{��侹qD�
>\�y�͞2E 8��{��Ѝ"ŃN�SՃ 8��S]��,|^D5���A���Z
)���N�����}���볬����{YN��Rݚ�o�����#:U�t�cw�Ӛ铘���'GƳf^�4�w[(^9���[���Ҩ��`�j�p��:���5�Dβ��矀̐@,�
�!"�"��Ͼ���������������)*���޼wf�@��G1 �P=�[��s�w��|�昫��!M4��i��h�\�ML霎�C�K������f�U�z;�H��g~$E��`��2���.K��ae{k��߻�������v��}�����\��bo�au�;�7��f���(�4@��ѐ�=�VЂG\,���PN%J���$�.�:3"�؎X6�K���湚�8w�Y���6���r����7��|�,9�E.��}����ҟ�r��6�y����PsN�݈�l5:�4�f��l���K��1a���[W��&dƍ��mG�G&^_M���#�vՅ�ǀ�|�y�9����	!
I@�<�s�}��s�/��9�}���� ��$��
��w���_S�|�/��49�y�6��y�b��V��a�З*NM�OՠVB��rVĤ�-�+yO�=���\�_;u��(mݜ���ϋE������p�F�t,��n8�������OKO��sTk}���3ݼ�D�^;̫X���<�R�I�:���3���x��J���3Q*��z�2g��fTe|l�vW�6	�3��]�wۨ�jӄ��օw2C���<o�����9�j����=Ȓo�ƒ�Ә%�4h�G�6'1�z��a�VY,p�NҐ����������b��_xw�"+&�q1[�l#�u�W;��]2��L�Sj���}�u����x���w�y��� �RP RI���B�߹��������}x�R�T붚7|~�k\{������D~�xnyu�o+ۼ8��d=Ǳ�0�P>�Mm���<X��c{r�^�|������8��2��"}T�f��e���?8��x����~�G�]0�NR��^y�~`i7�2t��#Ns�LuP%�ٵ�~���8\^�������P��^2_��/Яe�|�3\����y�@-閙������������u[+��=����X��-!���Z� �Zpηܨb��f�o��%��j>�yS��dQ�����m@�ё����*��	��p�e�>���/�Ӎ��6C5�����w_����>dx5~R��������w��4uSG�f�ШF�UB����^�s+���#�X�E"n��ܬ5����Q�2�c�Vh][Ś��w^5%�''��kLt1�I�ba����}U���H���B) (YL��G�-l������F~��yo&���^�o�I2�8W�	i�ey���cM���͒@}�����	�5��z����J��<�כ�=Me�H��lF��zZ��S
r���٘4�1w��-<5������CVB��D����.2���3�}����Nߓp�e�p��!W�0`�����Պ�դ$���z�3��"��s_����B}��}Hi怲J ey}�ݬ���{��*?D%!��i����1m�'��iiY��S�_��=��pp�H�`�:������6���N�\�������sN�|�]:�L�˸���j�����ق�̺R�秚l�=��:|lr�ykDaq_g '���/���skr�-��=�ـ���"�(Ǆ�p� �t�n]���$)rXփ�0c��UL���
%��s���@�H$Ӓ�[���h�U���Y����x���^s�y� ?0�R (RH,��H$"�$6{��{��Yr@��	��5��d���ب7�7U��?.���V��l?�8VLH�9#z�0P���x�+ݗ�u�
���*-T9�FVW�����M��Rӿ�jȾ`%^7'��Ϫ�*�j/l��Ş#��?!-/{mvZ�W������A�_����O������f���Q�IP�R�1��"$H���$3�+��/���gU~_��7����?�1�x����_"t�+<�<u�ڛپ��6����U�
2�yF�ꕫ$]��cޝ���}�w�6���e�zE���44���~u�&�����D�� `�<�������c��0~^7i�#y8W�j���%WXǄem���F�;W9��n]x�;�EQ�i�{WV&jK�Z�a���E�֘�د�vv�@�0dyE���_m�b�7�N���)�ڪ��o��
I!���$�	@��~����d�ELl�����P�^\���e�qvؕ����y�ᤆxj���������<����Jb��S���m�Vz�A����^/Q<b��6��'�sxr����۪�F������5��c�w��Wj�~��m��׼~�:�;��D�b� �2}����x�֏�n���������^HQv�\�S������x�/j�[�S[�۾胛Ɇ�c�Unˮ��������Nu	Fj69ِ,�0r{|1���Y��F�f�)>F�:�)i1Y��_Bٝ��~�\yN��n1��&�^��$��ӈbk$<��WM��{�q�C��x���X}�r����#�F�'��2�����>Ri���;w��q�UgZ�d���徙��������ћ��N�t��|�6��;�בKx�	��/6>�ҳ`Q��iI{�'?~����E��XH�H�"�o��y��;�쉝�%m�R��Y��ω���(������o�ð��o�w�5�P�q"��帺��=,���j���wV�ŭ�M=�R&?
�TQ��P����K���r����~�����5��oNu!��ϒ��u�g�ӝU?b�ށ�A�%�E��wFaL`��e�g��zo-�����|�Upm*<i��W0g���st҉�@���K�Ȯi�S=���7��|���[�(������p��,[>�蔥}9ś��:rN�ګ������dTɝ���"HS���G��L),\ɸ�fR�� ���u��k����\9��<=ώ�Dծc���-�-;)��<�m�fOzd!��>۸F�X.۫<�yb�ՙY+d�q�8�3RLԾ�� l���Ql�}�& �n^�:j0�K�s�kE	�M��I�T��\����~a"�E I�$B,!=�����~��O�}g:���;��V�#��3���GO�x�/������܆�E�k�����0��r�Du©�^�8�{ON+��m�Wz�>���e�3�:�0Eeѥ*y����dxe0ΐ�;�m9��Ƈ�љk��ـ��-�a�6����K��*�љ���j����ym;(MtgUmYQ��c�W�4/y�`�M��>:�7��ڻޱ�m@�:���T�Ctg;�����K	�.���G��syM�~�Cw}=�ݎ�<�|��f��4�#0 ��T���n�H�ymh�x�r�F)�<|x�e���Zl��������SQ��g�W�b�YvA�����^�?�߈|~|���A��	�aZ?e]�ʮ>���ڕ@H!�sml�ooc�ǁ ��0��׃%i0l0A�e�kk�1[z�s�����ӅѭtUa�co�N6r�9�,{|���|�Y�7��Ǐ,9�_J�[1�m�O�X��t6"�Y9���1k�gn2�ZY�n����e�[][N�n��8��՜�L����D:�x�%k��u-��UC�;�eb�pb��E
Jb���x���o^��>��,έtŘ{S� ŸsDO���L���U��щ���M��'��V  �x���G��7ˏSpv������Lz0=w�A��L�{����
�X��OE
�H�<�C%�Ŧ�e^euX"aٍ�L$��*�,��RrT��z��*T��K�gR�+dچkA�u%j��rSg�3s9�u5�J#�Dy!ф�s)�x�"�������L�%�M��*2��F4�*$��I�1���AӊH�b6!/���UADg��Q�u���!W�f�����枨��u�р��dĶ��;˒�Rœ�$�p��Mf���IJ�\w6;�L�T85�Q���s��)�\k�L�6��ب�����$Ep�D$����a�*dM'��휺�5]�5�k�"�2��N4u�ڱ�!�{P�)[��#�g^�dʁk6���٘�u��~϶F��^�W#�����W�R��)���3rtc]'2e�����b;a�w�xV�l�{�>�#���Ҏ�+0�;�mʿ�g�v��t�7����,JAFxc����^��ioo�(�/E���R�+��br�j\Y��\�ٻ�y�:4�GZ�q93��'cP��ϻ;s�]�X��s��we���/�bP�������6�^	ƖVIMҎ���@��ֵ�������#��.
�b\~ʣ��̙�kE�Zu���E����]��QAݖ�7*��$��q�37B鮔��K��[�]�7XFŲbb*e��޺��m�IR�"���c��	��b��B��]m7�n�RԔ�qQ�n3��m4��������s1�7[뭥V:ك��mZ2j�+Q����9�
��Z��0�L�������۵�`Q���. �Z�a�,��%s1�ƢȰ���}Y��Ҙ�3�\Ȫb�*�̡��V���)Es�*�.��.Y��w��:`��D�ӊcq31L�3��D���D�
�c9J�F`�c+�1r�*cJ�����)�C��l�I�~:.1���o}�d�d,�B��ڐ*�9|t���	2��7Ie�O��@>d"�E$�  ),��� N���_�~��5Q�?�J�:����y̞�li<���8���2z%"ڿoi���a$q���%������CZI���'��!R���{x#	�䂭k�Ռ��BTqM~5��[��jsљ�LK�J�hR��{������n�HLUj��9�M�U��=�ו��Hߵ������d�_Ygs_�N�UlUG>�qx�|�(5�0��#wS�������s���
?Q������D�u*?y�x��RBr�^ŧ���z	�gen�ݥ܉��I�N	����A���p��}K�W,���Fͽ��Ë��τ�l�3�L��=B1WFfX��+�*�@ʼ��wDt�u$��c��Hj�N��$��x��g��Y��cN��z놡���~#��1�œٮ�>,� �%�ɮ��P�f�wS���N�q�L�z6�u�
�Y�3o�7$ѹ��U_���UwU�R��A`�! �������E�9��.<pm��E��l"�&v�7��kmڌ��I~�Em୧l�/�Sӱq���|Ն�#�{���'/�)�1Q�z��;B�3���O�#<�X���'����N˯wmY�ǘ�1��D~�������so�]{����!d�|�t��#��
�z��e�>�m'���H���#N�4���@���N-?xѩF�,�c������"L�RfeD�ƛ���~��UL_t<S����X����>��
 ���c�Ib�BCi�;��A�f씲S�S��Ž�-�Vo���a�q��%�>8Gm�<a➤=Z�1�o��\����ԃ�b�ĩ���o����J�������j���J�%C��rT1��8�
7���j����*�j5w-�����r]������A-�}&Q�Vu;ʀ����EU���Y�I�/�k����� 	|$�P"��@�<��~��C��?��%�Hq���R���;>3�Ψ2�U��{�����]$	u)3����������)i$�~�ɝ!���tXN`�f�ҷ�ρ7��u]	����ʂ37�Pw�x�����{Q׬x��^5�Z�B��0�e�j��x��k�ͧ�z��Y�-�&����uǍ�2�n�ָ���ܔ~�S����M��C�u/�ʏ�ڿR�Aս7�b�y�'����n� Mu�l�$_!�{�
l#GM�1�o����x-���&]k�b$�x��;�'pGg�2�l�rV�G6y&�
���Xr�;����E:��ad���&���������V{�Х�����#�r��c���<��&I�^�Ԏ���3��窾fh��-���}Q�hM�,Nz��q�RW[��\�L�襍gqqU� �m�7��lS$�!ٽ��L���$��%�?k�?2��,�R� �m��y����y�;�^TI�jcbjL��:�<��J��]�v�}�R+�SE�]�?��*�����_+����N��ܵ�ץ�7v��0�d�<]-!y���[�q2�go�f�|G��|wR6~qC�Zr[�C��u�xUk�_�}�CB,Q��j���[Ց�6v�3���ʹ3.ǭ�8K)�3
��� �o���Z���*���ܵ��-�*!�����З���P�a��j������²r��Q���S����/�P>!��}Lx�{Ӎo?hC�5]{�zy+!W^���\���^]7Bܽ���ى�I�"�c �
vUc��{G/��x�MB��Ԏ/�ܽ�� ��lrXDZ��Y��7Mң�Ldu%u5Z���S�ڱt����D>!���9ø�IG�F��UN*����`������Y�u%���i�R�su��{�ǒN~��W���)"�H,��a$��oȷ������/�B��w,�����v����w*a*��SuJ�=�	�pd�|�K5k���Mw1�!ZB���x�#gӭݬ��������oN���gǍ�,���v�NB��n�īN{t6�GN;�H
��a�iW�ߏ��>zz�)����?{~�\��d��k4�]��W�r
[�ռC�w=3���I�Dz��4�������8���%�j��`�&��4�vC�ה	f%�k<I���.��׶�J>��ǖ�!���	<�ļ�*cz8R�"��}L� ����@����hK��yjR����;~W�9�u]NX�+�W�6��B-�\�F���63�te�P��^tx釥E�k~���!U�]�JJue�&���t
�f�W�Rs{ү�Y����>��g,��0���QR�Q�y�R��Ԣ�Np��¤��������"��B(E$����������X��'J����ƙ�������b����|}:o	Zgb�7s�|���Iơg�|��^7K�)g)��4�������W�����?Y���L��Ў*��ͱm�)�%Į�-1��j0�5NW����ĒE��>Ct6����+.�ķ�އ��K�if�!.]>������I�CIq�s�vz����FCZ�U�ؾ��sK;˞��@���uf�6�d���KS�N��*�g!޿߭�B���*�˖ymF��mZ�v�pWg�{�%[��a��01KNy)��V�'�{��c-FP���QN�x$F!%��q�(Q#��`铬�P�L�\�70L���^UF��|�┸��B^������R�EZ�润��U�j>���>��՘bc_�79�L.�#ܒ�gme��Y�r���2�7�q�+65"Ѳ�X��Y��κ���ć�RABE���P��u�=����[�4^>���9��e+Z#%X���v���;7ƈ�����i����y���$B4�ù���L �,�ٟ�$o{�}�t՘C�E�x�~����%U�V��<����;�Z������ʡGܦ4�!�M_��G6�Vz�D�V�:ߌ��%���:���k���g�Zý~}t��n����`"��K!Y�Q��S�4q�KÏ�k,l�k���{Q>�Da�C�ʟx+�\��6��B�I�ķ��wS������\ͮ�s�QΡɐi�ꖻ�\��Yc�,�A�����?C�(���%�q�P�Ǎy�vT�,u�8x�fn��R���L����L	s3�;K�+#�Y�u����@�����#&Q��驊0�jѬ�5Rd�hm�u�ğ��[El9I]��'^ �Y����d�4`�p�岳�w5����z޷�}���~dR)"��Y"�ď��[�߽��5��a���4X�4�p��<�S�ٿL��6�?M������ޛ�x5����Cܴ�"I�\I|�;���될z�*���Ǳy���k�u1Mi�AVC�$Y6�=��{�;ő�h�Zm�B\z����J)С`r��}957���|OĪXp�b u�q��A�X��p�[�q�v��A��47�g�9�w�}Z�����'��\`�ʞ?�{��g��!�M��R���1�B�"���WRЎ��~��^�wr�]z�5��[��*��<�fo:�s��qs]���撹^�)��F�5LSy�)RZf!��<6�F�c�;7=�%�A�w9��O�%aTV��l�5���9ƣY;�(A����41W�. \�:����:J�Q���*]�|Z3��b��5�ojv�\u��}���ަ_h�v"$�XnӸ��fqjm7?k�������@B,�{ν�_y�~�zs%�Wz�>��2�B_���}�~�|J盳wk��
��y!�<���B,�;sb\�{��a�S�Q��[Eg.#�����T��6���H�ւ�#�f�k.rB�����N���݅}33;�ff wr2�!�M��^�i|Bf��MY�/�i~,b�VI�M���!w������䓜�2��[���z��Pt�����^j�w{#C��'���\�IY�s�>�%�����-a��5ײZ�tY���
8W�B����B��dŕ����zg�={�{(��}������{ȑ�+=��_��cf������*��7���:�!��az��H�0���Tr�RJ�6\Bm	TF�Z��ߤ�0;���Ju���]���ԍg	ٙ��QŒ3m��SsW��n�T��m�`��{�j�q\=ۤ��`+��
���_�Uw_|)�Y$XE!��}��x?ǘm��+��AV;z��:$)i�nD��HF�N�ɘLٚ��S�D���~������W+�2�?r��eEr��k'Z�P�͟:i���u[y�^�$m{'����dO-��?7{fi�����n�\./�"���&�\i(3�bcx����cc��|�?fˎ����/q�_�����O��F�#���f��͡&'eN��0�����m���T9}X��a���K�f�xu�A���;R�Vv$8��NZO Lt�E�*�ǉx�ff3#�:�Q���ˢ��	U���lXr.:}��B8���) L8E^�Ne�W�}�}�C*\d0��ʂ�ؾ���i���,.�C�� |Mݙ�{�ݿ��G�%�K3�_Mڵ�nf��ܕx
�WrE�;bZ��!��]i+�� %:�2g	a5��L�+��k%���N��f���+��бx$�!h��q�KȸB�,��YM���kr�4��d�v���8�%z��W@�)(B���qa�Ł�ת4x��E�N������gn�d7��蒿�Obӳ��G��Gk.e��_8�(�!;27��Fw�w7�Q�n��=6��ͮ8�3{���9�59OAѤU���ѵ��Y-4�j��Z��\���
��G7��YYN�wr�XFm�QͬՀ���qNoV�u��7� ]�b�e("s	���m��+��mU༇
ܲv�Ys�j)�X�F��b�s�ӕ�N ��������_&��+��(�#��Ь�tz�V9Ii�i,���LvPF�H���&��Y�o�s��7��ި7:��,�!�D��'t���D�5��}��-e�x�l�!ȕ�ռ=ޠ����9��fT��Rػ��K":eV��u͢���B�Q�����V��CXl�'S8���u�6j�4�uf/p^�U���eؼW΄��7�mg�[�|+%=,v�>��V¬L^^���Ih�5-���Nn(�~��d����,j!�e���c���-���ƣ8���-dޙ����YUҢJ⨗t8��-4I�:�{��4ֺ�ss^4OWb��
1�8�����Q���]Z���2��䶏En��Ը��h��$b���wk �c�Lg�7�)s�1SZn�tv�Y��1�.J��p��#�Yv����ZKR�3I�E���ßJ/"h(Ҳ�Vھr�VQ7�������Hl��`����E�T�r㖥�L�[R�Y�D�kV�c�Z�g}�{V,DQT�QL���aQ���"LB��,�2���#�M����"�X��:��ciJ�e�3Q�4`�Z��{ٶ�3��q�S.�r�r�hۘQ�3G(&7y��f�PD���d��2�bC%L�2�k+(�6������W�s#h��5.GQ�EE�Lq�by��a���̣��RܮW\���imr�m�UB�r��o}ov���b4���\cs1�-�ԩ\��o}ovu�m��e)�Qj�m�e�26�\�f �E�r�!i��U+F��b�k�ȃ�T*������9x+�w���F9^�Us��ǎ�دX�+�o���<�ּ�o~s��'�Y`�)"��߾�����޾��v��x��S���3�|��V�@n\����4g`����{����g�I7o���Ŏ�w=*KVr�j9xUcAa"�y������.#�6/#��7��ҡ�7���ٿ�M������g|["j���r�"�/j�����%��^���뤹ݮ?qz�^٣�A�<�_e�ָ������1�}�j ս(Ҩ�Fd��A�Pu�p%���	3�~T�����(���8��O��]S��kv��|x�+v#�BZ$q��eH<n`eB��1�]��RM�7U�r5���2����?<*}l3����g�ܕ'����ow؟ϱ�����Wڅ1n�+�+`�xJ[�0F�����:w�ZB,l^��v��Čؒ�f�{��a�A&��;YA8.�1�3-vl�s������M�l��p�fH����Uw`�R()$��s�}�o:O��.�фUQ��x��}���/u|L��W��@���a�+�Ց���uC��Ǧ�^��E)�U_ƤwFm+�����c�l�(��d'������|.��V�T)}/53#Nk	�
n]�)�ܚ�c�]�y����
�7��a�3ܛ�>��k�����ߖ��8��|��O>�����[:������A�.5,y|�򐻻(K��]�¡�Ha����g���>hV�������n�����l��i�1rs�Z%s�`�TgӢ�T9�Z�B��o-��B�v����s���Օ�<�(���z��rQ�]_������Z��f61]0mf��i)R�5��3��hZ���<� N�������=�eҴU~�B�!�Lc/p^�c�h��2u�ܸJvt�z$�#��L�ai��ה�p4�ޥ��Y�JqMV���F���<��9�f�&���O�矡?! �P

C]}��z�����5�� kC��>ei���~cqF�0�zY5ٝ��޴3��)�L#J�>;���#�{E�i���6]�K�hk◽�,��Э!��b��	����(ύG�� T�؃d���Kڹ�;��P�T��9�b�v�6b������⸦�v�m��}��\��bX���)1�ޟP��*z��ev�gݡ�:�$=0�ߦ��fv��{��W��L�nr宽��hSf�+h�hi-zz����W�R�VEF=k�V�����*��/V�!Lk�I5
����H�6��FY#�-��\XXp�q[bN�{Q�g+�	k�����í^���O<�ۿ�z�"���ܷ�U��!�4;��m�/Pm=* �Uzvh2�>\c�a�2A����x�f�vͧ��Ed��-0��7���a��\���P]�8�aoRͭ>�m�Z�"���k,(c�;t��i7?��E��dX(�Rk�~�߽�^n��)��Ʈ>8C�	��q���F�].5E�YQ�'g��&�>	Z�.#J�}����j�G����]�e{{�_!�*�(?Y���)-��,�0�.�4�ׂ���f�J5T�_)�7�!H��a��oK����A�N���w���Ȓ�
�4���`b:�HV%�q|I	���z�V콻���70���R�<���W/��א�Ui
��"�ݝ�y�|�޴"yY������f�C����濼�1����b$_[äD��������3-���碖u�R^�6����a���Qa�ť� |+���.��`P�t��~���]"���z��}S�p�D�&���z\��(uʺH1����Sa_�m�hwD��d+&�׾���/d�3yQg��U�e�����1WLX�;�N�#:���\�Uˋ��s�����껪���� �E(����߽�|C�o9�?�r�n��/��P�GXwDbW��H\,�x��=Ng٢\��J��X��P?c�331u'Uw9�3\��Ǐ�{��m�1�t��N�㧆�A�����@���a�0�|33930�]LI�iҳ,W�{ ��R�J�o\�m�uK��|�]Q=-���Su�b§HK�>!�@��s1�]��wλs��^h#���y1U�?:C��0CF;���7�Ggٺ���PKv,�Fӻ�t.�,R���=��"�\;+��D�:}���[Ip�$U�D�kׇ����d^���c�ӈQ��Ԋ�4R�2bT�sQ��w��Q4J��r^hJ���I>P�[ҋ�c�I�t$@6���{^?��wYd5�^�3���e#��}�t�|�W���9��Vy�.�&�,�W��[4N���j��rt���IN~��W����P�"�P�d�}�}Ͼ�����JVZXg?�y�?>CH��F�xןm�y�����r#O���uh��V���?�l���q�铮7R�O�/.$�^=ʀ�zg!K����l9Rtu�<�9,2�]���yџa���-{��r����'�O��L���?{�C�|�Kĸ�<��~�b��F|�B�8�Ν�ي�߳D>H9̑Qq&Z�����S5��R��;?�,��~�F
�b֐��8��1�_r����CNZz�|��O�:�~�g�#	2�Xv��$��ٟyn/Zɍ}36�]�,Ze�|�5z���2UT��)&/�T�~w�h�D��"�OJ8w5���ƾ��<�rӄ�kG+p�sq�vN�"磊SUKu��٫U�7F���Syht9v� �7�ң�7Cm�k��/8JU9D���6�f)��.ݸ����9�Щ?~? (
�)��Bk��}ן{���:8Giu�lyE���/�id��U��!��o���c��n[���I�1�8��8C<{�������z�f�o1��!f�l�'�S���A�zq��0h\Z٪nخ�=��$��W�h�h�l���Uty�ʼ�69��jY�ߦ^]r�}����ﵒ|����q�l��3{Ja���*Q���n�ٹ����r'�47�ԍ��MkG�Zs����]�	(���K���X�=�qD�u�'Q��F@���d�P���_1��3㖷P��^�`.�ǹq�����]�Z����1轨��V�4���	\/�W
q��W���=]d�w��a���������!�>����^# �8��zqwg�����%^`lY�K3�X����B��\�d�n�To-��Q�tMB�VE(J�#OF:^�/+F^�Vs��_i�_HgTM.w�~�,
,�I��ߜ���ǈ}���O-!�h�N�<��AQ1��]/��y�4���u³M�\mF��ک��4%L���{ 繞dW����vR"AN����(%�w�L�"��������A"ϗ���o�*������wJ�u����r�yj ��?%�+�*�+"|^/�F��H����˟��}r��`��%��#/�i:����G�������6fn����������ގ��RXϕ��������4[B��2��SqT&�l��4����rTe7bT]w���"7RK�P(S/ˈ�^�E�j�D����.�y�(��<bʌ���m����H��R{}Z�erʰ]�z`t{Z�2��XةO;��&ȶ&+?aڴ�H���z�W׍����%�V��z�E�]k:;n��=��s����AA@R
�R�y�����m���D��e�]o����i���/h;��Ϣ��E1����������!���]b������K��sf,�r�{.p������s2gj��K���A��|<�\rX�t��7��P��RdY'.:0Ć�zf.5�xS��go�f�D��z2�/ν1�E���%b���F��N<+4�9_���~��$���V�n{�J��b(��t�q2Ka.Χ�u�UT��QΜ�ͳ'6ܫ�V�K���l�����^��:����<�s�����o�qx������]��j���k��q��^AO4��+N��A��$N%�?�Fbւ5��`��I����ìg�*?�\�O��Aُ���"���t�TyL��0�2A7�p8m�ѲW�"�r�}׽�@ޥwt�:��z� ms�[�F=/:�ν���È�(�1�V�m�î��<��C�A`
H�RAI&~�耽�y��_��B�*jx�T�&��h�<BK�E�N���pg����Z�f��L]ӵn�%e�u_�dwO�o����f$<Ӌ�jC��~a^<`�^�|�L2��w��o�{��(+�愩�H��9?)�H*ސ�r<���u�#�3=����Ϡ�d�/tz|��M4��Q�ψSy<�Oݻ߲mQ�!��;�Z��#���.k&
���^�֋�2'랙�� ��u�D2��C��eZqI{=��wW�'�z|f-=�}��*�r�%$Ճ�F~[WiiI�&��w��jM~"R�}wU�JU�Hr�����r���%�ŧ�|B$�=�6x���z��=�63_���r�x��URkA=�wG��έZ�Ja0�8Vn�n���J����9)SO7FC31�J�a[ySy�1�v�9lk���-�y�q�N���/�����o5��)D�c���:�`8��o�T�^.���a.�ۧ+��FU�F���{��l����r�1�W���v�t�}4J��yG�N�"VS��KRv℁���@�nLO�,Y�=X��aީ��JA ;�
"��5"�"��y+��p#��6�#��6m��M�~A�aܫ/�3wQ�ު��j;b�RL��v�,.wLs���]��j�@Ј9i�ӣ��_=�!�c�Puj�,����^;\U��A�Y��b���t��\����ޡ�D�+h! y�f<�KV��)-J���d�mFc���k!a�},��j�IN�zn�-sF\"�[�6�ic���y[�h;�ۥ#��\T�͵aQ�֎�v�}��I�E&�ϔ	�Ϝ��}JBÔ�(CN?��3�U#x��V����o�� غ7�v��U�z�b�>��}Q�g5�m,RI�c%%��d+o .��N�B�%���榔/:��p6n�*p���E.�B���U�<��*Q����v��	67k����p�#� �;���&n
��u��v�g��b�pwi��Y�T����Ӥ��zyE�]�V(�7D_ ��ɬ/(�<0�e��Z�\���.j�u��tMo� �+N�J)�L��vZ�7h���5����u��[�����񪚝��hG� �6rɝ*VH�9��	4���s�/o����A�g'P��cr)�3Na꿁a��:��Vc
,�I�-s�)�.@��J���)�j9]s󹧤��ظN���ۋ�) �z�yO��lJ]���I���B���.��ݡX�P�.Z1De����Qm�fe��)�L�]����e�Vs)r�J̍k*DY��(���Kir����ͫUQe�wE��r�`�Y���s	V1H�j1���n���;���aJ���`br�L�Ȫ�3{���ݶؔ��6����.S1,m�k(8���J�\��{ث��kM�LA�0`���f2�R�{���\�4�S��,������W{��m,dX-Cw0q*�U�j`���ﭩ�B��[[b�F�2*�2�r�S3V����r�l�"ɂ�����Z��A��kh�;ʲ�7�6�p����GiG^�+���d�It�9#%����]��)�g	Պ�������?}�0�H�d�{�������~���:ZC><x�F=d�ָ���㢼��Μs^h�[�s�EO��J��u[�R�wQ*�=G�ʪ��mj�� ��C�Y��
��@�9�Ѳ4�y�
k�^&������K�߽���Ŕu�$o�Fbfd@6�V����|��>�M���\h�Q�^C��"5�0��?Z��a�������F��9K�dGkB�S�j��B��˚�|y&j�#�T��J�����ÿ��)��x�U%;v�W9��g7������Dد����4(��Rtr�)\�5����)����������L;A�� iw�|�ZD�@y��練�~�پ����c��*�&��^5��`��kX?�j��y����"�%1 Ci��I{R�h�T�хsV!v�i�VMr5�G��j��;׺3�cp��fLj6oL�TD;ZR^�i����o��������XH)BO=�}��������E<�b�Eo0�LS��(�ZV��/FP�i�'�޿��e�mǒ�1]��g6��7�m�s2A��G����td�
lCV� Hsÿr�ia����\_���]_��^�Ն~��G�Q�Ha�>˗Ye�W -ȧ�[��OO��%�З��V����#��Z|о�Aⶶ�0
����� n��n"�ڍ�촉�l鯒Y��bf���J��q��`+������c%��&��/�k���N&B��K�lw���tH4g���^#�-xz��Ņ�����Nw��f�s
MO{*]z��+D]]H �,���þ�%˥b�q�,����e�?��7�C�He�7�bJj������z=.�������^&���n�qW�en�(���d�wA!�0�/B̖:nh/�Je��Vn��⧛�m�X�Ňt�]6�sݶ�5;O$��U��("őH):��>�߾����D�<~�r%?*V{�l��@�TܵU��۽Ы^�a�l<G˧��N�Q'���@�W�ZK�۵��IbΑ�%�Lacˈ�u~��ԹK�3��/i��u��K`c�Sr�����SB����XEc������fV���瑽���{���g����Le�����f�^���~�O+��Tg��'����B�2~�%6ytCs�dB�ʶ�;�ق���G�*.���|�K��la���t�ɗ�羚}��;yWk��/��p�'*:0Ć�zw+�=A'�	Mml��S��"~��tz�B���ŅIa���z�����n�{��:I�1�⳰s���Y�b�X9|���-�O��ȉ��9��K~̡��V�O���m�3'wU�`��]y�zL�Y��,��:x1tn��Sn�R��ڮ.�"�sGt�v%'�W��U��R�b��C^��>�}�kG�w}תr�"DU��.a�2v���a�GN�z7���op������(Ĵ���戥��[����޳"�흌R��)F)/�}0�ㆵ#�Y�i�Ci��*	~5��ȥ�*��ɥs��+�ˋ��J������?@�\�3=7:���\�J���SZrp�&p��r�7�f.!o�R+II޾m��w�:E���E�ҕ.n�-�5���KhS�H&F3^�{�3��^~xq �x�p�*����86^{���gG6��g�����J�@����>Ci ���> �y
����_���O��Ui�Ւp�s���N453���*t��Et�U2�[�rg%�jw4}<��	,Z��U��g.b,�~2I}}N����9�g�.������r�Z��>��x�Q|����|.����6�f7(vFX�p��f�ۏ3{Gn���33Af��T���n�ffg��?��R��WnFK���G���oL�!�uc�겐���[܆?xW�m���Q
ޱ��fUqL
v�`���C2��{��޻����>3W��K�q��U���~6t���Gi�uI�~�P3ty���A�ik3x-N}�	�93��ti�Q؂afz��:�^�W�i6P�kH��x�393q�rWZ�3�U}���*
�XM�K|p�&"2��8IP�
��[e��{��1�(bg�Q�K��V�XX�h�H8C��/}ݝ�@���p%�ٖ�'��#<�r��?!�9�x�&�F���Zekl6��z�:��˸��?i<���	�ZC�6��;S�f�yϦO������dF�����!����zT��W�w�@#Ж���؅��;7�g�H���7ud�I���ow�$�n���w�u���%h�n��#Es��1t�X�]\�7���T�s�xz�!�!ak��ʓ��/�ݩ�4������d�,�FT;�����-�B��h�?��y\��][�{ځ>��7����':G�_#�����R.���j+GQ��������/�j�c1�/�~S�0�o:�Cu����k���]ȩ6������@�;9+���11e\�ZU���.�,4VuU��1�u\�
:k��#q"�S~�����g��R˽���88�]���X�hEk�:���ؔ+�ꮖ�[|�|��`����X�T�;���?s̽e�T�ؾ�(�e�_a����uFv,8ᠭ��:�=<���(y{s�:�_�{(�������`:B��%�Q�p�i���^���}+v��1�Rջ�G6N8�M�Y�/�* GzLe>�5�96�}��dYx1���+/$Z�9���]7��(MG38�d�q0�b3�.�r"���}?u�k�V��]��>��s-ɳ��Y)Q ��C�w��>Zf[��Z/�.�c)R�䚓���t�L?�TTu6�A�������`�%�8���~�����%�V�Ղ���gx*�	x2�h^]� g���*y���1?z���O�3臏���$�l�]+;��!*�fv)�C[�i��5Q>v]zD�������v��5h�����o�����So}y�<-�%�!�i&!gN�V�"EbG�o������&�"_Q��t�*0�𠇘��1o܇�����i�TJ������b��n}.� �V-h۞.�F��>��z���.�z�S�{����8�dM[)��aLs$޵^�ӂwwA1]\n}FqN�m���7�E>$R*_���qe{�V�N���i3�ا]d&�5���������:՗�*�J�G738�Z��p)z"��Ro�f�ڼGMttƸтQa���'f<�EE��Jq筍�)!R���Ъ��8үs����RdKD�TY�����|0/?{��=e�{f�^ܿU�x�`�W!��|,�_�:};�73�w�b�Mx���8��U3��`�4�;�\��P3wo;ڽ��G�#���ށ@�8c�G�t�u�9��I�p!E�u�k~Pj
�y�(�8t�"(����ؼ���������η�9a�t��w��,��VY,� /��ҹt�����XuH4x2�y������W�Z%���,D�w~��K���=>��d�v6L�� րз��3ʢ���]�G��}��w*!%�q�i)i��a!��z	LK�z׸�5}���M2�mYd.��.��ش�:���@X�YYM"U��$~!����D�1�YϾ<�Gudw=k�_*��,䤹�{�����Js9���j�T�Ƕ+�T(J��.~|x�ƹT�|x�����b��bי�Ѥ�(!����D9��/I>e�CH?��E�ߊ�M�w���Y:���Xv6m,3�����M}���^���
�8��f�L8�rd�)�Q�Y/��BWR��VUG��������eΈz��Jc��#ZI�ǹX�zx��t�b4��I�u��S
�0Ϗ�]�0ZúE*s*��I��:���[=*������S_�5x�x���������{��a]��W�8��AͩϦ*&���q�sY.c�Du�1㧷�=K�f�������:�!�0�E�K�F�h[�	��k�2����mWH����2nF�3���l>��$���l����T�1WC��}�f	��6�z�VZ5�c�L��=ewb̻��鄌���z�i�]�7n\�3�I�{��{{y�65D�����IV�
^��M�)�?�f�Շ���5��S��XsR5hi��˱��vw�#օ��A�̑f9}�F��Q�&zs�-F��Iy�o��H��xbC�k��g�*մ�cgߞD#ZE�ɖ����V�?xu�K���Ri�o�qW+��C��Yޏ��E��ׇ��<�`ô�p��#����� |��y��3�ݜ~&��мX�4��U���Κ]�,I�t�/c��s���^���	z�U����'H�Ӻ�Ȼ�y��+M�P��kpS#Z�Do��~c��&�V�㺑[��f��g�*t���o��/ӂ�tT9�P���SǠ����1ݻ0*�?^�(�K�>{�\L�o��5�fJ|~Q���舞��u���{����_
�Օ�U����ھ3���xe�AB���Dj˳�^��[{����(:��٧[�؋O��tre��4_@/v��x�j�u�)���n�U�R�r�f���7�:O�0����7ՙz�-Or���}��9�d��c�pU�����Uy|��1֮2�Wu��H7���1�S��fq�0C���nDր�o�+�Iu�^떏2�~k��s��<X���hḘٜ��Kz^�X7��E�j�`H��-�Z/F�6"��_^J9!YªY�c}f�D~�۩,�+`��b�ѠW4A��t4���ᬙ�G��yej0�fAs�EL���������m�^*�4ܢѾ���].'(��7�.ܶF����V8��0�����*v�}Y�)֔)* �[���fne٩*a(y�����~M��)ou���θfX01T���7e��!�K�^j�\;�j�U�q�y�5
6�]���2����38��p���m�6�
��NT����8:\-��v�b�-S� �2��eM939M@�3�� ��|��OpUɳ�-����̇����'�NrN�1��uq�,�*CdgP�\^�}ˎ6D/���\�x�2��&h��d�W�E��[CN�kz�D�L�p�.�ј���k�&��O\�G{��F�]hӻ�qfo��)��ϳqaz�B��������-h���@]���Zl\&Z��Z	'R�j�Z����*�5ލz���H�B:�S3we��a���Y��v���rt��v̇�Lwl�§f�^��G:�bL=�9�Sm�'+4�&�A>Ul�CV�F#'�&Nik\�y"�É�U���|1�|�����oΆ��yV�5�*�qp�w��`��J6����+b֪����qP�5������he+#E�U�1�q)D+������ic�ecm`��s,����V�[��M�j��x\h�Z*Z&U
�s
�Z"�r⫙��{�[J������[mDQ��aXD�o{�gT��1+�B��eLE�%�j�qb\����m��.8T����cZ��32\��˛���v��)Z�2�*n7DaW7��}3k������
�U�e.Tc�9Je�Z"Ԩ����Q��2�3r�c�L�T�1����{���.N�1�M�}/����a���Sl ��K�S�ټ	_�	�G��U��	h2��XqW�X�hZ��夺xz�� Z��)_�U��j��9���
�c��Ha{Xg�{Y�:=��f{��}��x��������+h��-2�5͠�Bi\s�؟��Ourk##U�V���lk��Dѭ��)�� kKE���3��Yw���,~��NT-�~
�0��6O>��O0�^�o�=�#�q�]�{�_-C}�+�������TE,����H!�_%9Px�p�ei�Ӱ�	����o��>8Y��?�o�_�$V*����<���O�>-.���ɷ9��LB��w���f��O�>�s�y�����8��a�li<�P�M�#i4�L�����u��Evz��f,b��"��|e�7��8��tք��7V��K�Ն�ju�Y�W�h���j=�FN��}q��N�Q���5ǉKʒ�_5<D���R�ät�Ii�Ɩ1q�b:�_A��*��W��{�\����HQ4�3��;�K��Z���Y���sI!���qy2���}��L��Ju+1�t�.otn�dgn���T���k'��ޟ1Ax�ȑ�&���{7������C}��f��52;T:xÕE��K%9���vU����]l�&ȴ�!﫟r�k����Z���QgN/�����>s�Aϩqg�g�_���_�j�y:�3O�� 7�wdK�(_]ߘ�-\�]7��9-e&�=�.V|$Q��ϐ�m�1�a�_���2r6�*Y���/�J!K�s�Q�(���W�ů܏->R���&:�[=���Y�;c�(��v��_�.ع0q��Z��(��5�;�F�:���}���]�[-j,,N�m�.���( D���[&qj9�y�o��^>���`�ԍ,�!q�<�$D�?9=��]�;��|<�嘯<���S2+M};�2+�TW���_��*4x�,gόL���ȝ%�Əz��nw�"=��MԲ����R�cˍ��z�p�4�{.��G���H�o�|���A֛#�Mh���ʓ%��9Q�%����52�騭7��u�Е:i/�'�8�S�.'��{}��5��/���/Lb��,3�!g�/��ލxw����+*Y��Q�^�����`�Ӻ�]�Rć�oZ�" ���B=Md����j���3n�� �qܺ��$�U�]Ş�=�F�AG�Kc?AS�?<?���҅�Q�-��J�g櫗��t�X���*�$���*�z�.Rp�cJƲ�}7�V���](^5�)ٍ�M��[��z��.;�A��%�)Dβ��;�ɲn�%4q�τǤAKI�ȮB�ws����S��og��;ｳ��a|~&��<s��pR��_hie敼^�_GI��+�X� ����G�G���ɡ��&���/�{�r�]\���+�u���L�:��+</N�w?�����?&������fٓ��
�NG�~6T�9�~�!u�ĕ�&;4S,��(W#�uL��S".NQ��⭸���Z���|��/��>�{�)���.��������q�a��|��?~h���� �@�����x�VN��x�twJ�p:��ڛ���S��C[=�,�8��8����N��W�}�z���$ׅ��c���NKT�A��k@`�J�f�ꖐP�c3Q��^n98��IG8��)Vc�ł6Nl�5|�����
}��yH�qL_e孆k�;Np�?y�����[d��E��Š����i�p�cf�
`�\e�j�'���zj�ߵ�h��3�0}�F݂a�%��qm�V��N�n��J��H�{k�OT}�!Ŏ���t쬘�y�;b��b���/B~���x�6v5z�֜ ��n���E��CC4F�t���8�n��.63�OHi4���g�#9l��u=��0�'g=���K�4d�r��{�,�eӆ��K۵�X=��	KF�Y�l��fK]	$)�z�����+9�M����E���ံ7B�Ep�:�G	�u6U❄��s7��d;�I����=8y�c�7M�X|�w��عr{�p9�NI	WFm�}G܄�}讧�y��(�ga,T�Λ��nj�x]nӾl�����Q��������w��M�TiqO�"�}w�	U�����ע�Xp�9�ϜHxMM_�x��x�Ϋ���u`�h9��}�q!���zEڸR��
)`@$�ۋ8��W�H�s��Om�f�I$�M�5>��Eޭ73'/��&�-q�Ѷ9%����qխ.`��yW���3�2_j�ye��x�"�u�\�BRi�8y��Ӱ�&+�]t��:����4*l��dtWW���vʻ��+v��Y���\+7��&��M��:�;LL6�r��ԊN��C�q�}��v�.�A
�z��]?��t��Poۖ������<��ՅpP��TLU`0F�P���kRۀ�F��6'�����4N�ȝ�=%�A,(�|ӿ^�O�/c�=���~ܽ&U�o��,O�K�^�6z+v(Tk�|�KI�x���E�|�k��ns��ݸ׎ka>D+N5^�7����1��M�+N�-W��S(A6!��(��y.�����'�e���T's.5�%�q����:o�b���������5hk>6�Bls�0c\nu�v��7$�&@�V��7�^Z��w���HL��	`:��&����Xz��r𗃪RV"�V��(_j%!4�AaK88gD���jE�8uvQ<�4KD���X�v�|�J_�N#bx� �z�y��/R�j,6��[��=F�#ɔ�Ӎꓳ��{�H�_C�J'���;�D�N1ӌ=t�>�;������js������kKg.�J&vJ�U���WF�x��{�2�Y�,7�.����� �MA��P����� w@�`f�@�r�db���=�zZ>un8]���1�Y���6�
��;�l�2���z[o�˭��5~�TG�׆0z�7�E��O;�~�~��0e�Xu��@�qv$�c�S�����9�*��봭XM<�ZN��f���E��r9D͜�E.J5s�}1�ܚ��7ϒ��R5TcQ�7S>RS�G��N��	�E���n�g7��Wc��ZQ!�k�������ۛ���ۧ1D�Qr�*
���r�K��Θ�L�E�?,�_����I3 ��$��^Cbq(�\Ҋ��%mOu����Cσ�A{E?j�!� 5��z��V�^�����}=�(p�l{��
	���#���q�����,�se� \ӍT9��uXɼqРEi'�����	s�8���ז>�k�����b+y,Y��?�HH�5�Zƪ��ӑμ蘋����Բ�DV>�͛G��7�2)�΀�2$����ݜP�c;ZR^�I��\Q���VQ�g�Mŋ��t�.s�B{��8w"͸����V7���G�cv�w�h}�Nܥ����q�6`S�5
��ޢ&�R��Jep�E}�4�
»謭�x]p����P W��%���-��9��8����]Ӯmg	��P3l�(��˹qЫ�B�l#��X*��t+M�{�P./ތ�{;ya����#�t�>�A���M_��w��(�deZvfpD��Q1����̟�D��}�0"�m?g��u��� ~��ӏ
%R������JC�%��,����u�#9ܝ mZ2��Q�}�; �Ӣ�E��;��L��U�]\!�{�<(e��1���2UpB���֫$�X�;oiXu-Q�g�$�ŝ@�|P������h1�S+<>�j]ai��d���]X��0��gyK�%&��w"h���h�f��np�+Y�RQ�7;�o���{O+�dۣM�\́��4��:T�v��௦6Ү׼l�y?�^���b�kv��%;WX䰗yR�CƢ�\���9K����p�ȵ��.@L�sŎ�@j���^�}xv��N�o�`KV��������^����ۭQme��9��o,�G��i�2�����N�<��"��wE����mo���GG����Ď.
4��v����T���4.@u��m���-g�c��xBb�E�W��[� �B�ٔ�	�+���z��Ut́'D��e��iˡ 0�R �����"���>x᳝L�Y�LQ	��qzȃw�R�E������&���Y&R��m����/�bc�*��F��43�K2�F�\L�ն��hn�-w\��b��5c������[�CWp��bC(^dز�%w,t��'Q`��Dr	֧���j+�EZ�y[�Mf��-�,�]Wjt��J���U���vrmPb :.t���J���'�N��Xp>�<4�I���=���qDiJ��[o��׋�8�#Ǧ�h����mډ�����|tr��KS0e�aU�6y�7;v=k�t�b�
���:�j�*�n$/3R\���3&O��*�V�~��������sr_��!���)�����y�q��՗�	�6櫬��zjFGal@f����Rl˔���B���Ű�Ӯ*3e�eL���L�ԭ<.��`��)m�����r��j�$����onֵ�J�	��f[�L̍�0���[E��s{������v�.n5"e�\KLL2�s{�[�ټ*��X��"&Q���ԹL���Di������i�ɉUr���VۉZ�3.ZT˙����ՠ����)��(�f
�¥q�-�\n)QY������)k-��\��V���*��&�i2� ���Ai���J6�l�L��i���aJ�U�bL-[�����R��Q�)e�p��f\i��1�R��JZ�ffWs
drեr��Pip�̴��e��s����jZf²
A$i/߫��(Qu���fp�?&�T:�����of,:�BYݷ#U;�$���ݍ9\g�;B{�`~�U�X(ߧ���^��<:7�w�M�:�5/���{������^��I*��D[,�8�|A*�X�0�A�ЬUko���y[g��2�hMG8�{2%P�7ٴ"�{��Dǳ��b�Whv4��L9Y�R�ˡ�f�m���6�&��p�x�Myj�V�P��-5Ҥ�ȩ�R���Epi��u�ӝY}AI��t3µ��VQ��f���ʍqvJ�<;�q�{^�甕���7�5�|몎�p�1L�v<�����=s+�8�g�(t>�=onrgc��ܙ��C�ۊaם��J�~�e�6�n�Q�$�F%�� �+/u)��HD���v�/�����jY��2LdQ���7M�ƒ+�U��y�Ɛ�#�V4-s��2c����S�4Ne��xֻ����5�|�����B�Q�����N\���ՙ���g\���˪iE5ez������E�-��"�v-t��t�$y�&�)|� ��SؑU'�����x}�(|d�]K���lJ2�".u�&�Q��ZY�MKim�8��o�Vdtag��QQ������;�m<gO�J� t�;�5V`׭��P�n��V��W�6 s�Q�Ցn�7���e_��n���(��l�Lu=�Y�V;����u''"I*�7!�ZQBV$8P|�H��wB_N�{�n=O��L�oo4�i�O��y�����������#�J�"�#��O��T����2{��=ȹ�h��7DVl.�'6G}�i��j;T�3*�r-��s	A�k����ʢ��4z�Μ�\z�&�.�K:b�*1y��.2	 ��s������?�Q!��U���5�֏��	]�	���?p���(uT�r6<Ln����=�.��v����u��3I�<�S����v�R���[������_�@��4��~v�u5n5n�eb����٣�;�\	���7�iǞR�����M]h��X!U�f��s���#���"bV�v�K�RQh��;W6�-��}{����7~�}u~�/7�b����ٍ!F%'a�`87����M?�Ks�p-���4%vx{��s^���1Y�/����^ȶ_nĈC*��@7��Z�p6�p� �Q7�zr�{�2:�ͪ�{Eg�7[J<E�y��|{�M���������dHr'����7�Tܭ��.\J�޻�u�s'�ѐ赱$>x<ګ�xy5L�F��i#�لT�k�oJe5�s��k<o����ސ���cp�5;����egtu��,�HBPu�b�6�G��Ï0�Wb�VՃ��*�a$��^V�[�n.*����W�l�)��-�.<S�a蘣� ��Pi��@'Ш��-����V����9���y�İ��-�=��ڡ�;�f�����u���w��ff�La
oqP��=A�e��q7h����W�"�|���	�q`��=ٷ��׾[0Ɲ�[�6���g�T7�	���kg_5�[��/�����>g�ˆ6H��*�'��7���ȡ98x�ǧPI2�&9^���<${۳�:�QP��c����+ǌzNg�>��|��A��;i�Io�¯�{mv�r�g��MZӼw��`�����uUu�`��v@��ǳ���Bʢ}X����u�<��D[}!!�����-A;��[2�9��t}0�I8����/=y�P��]]j�RD�I��, ���OCnw\�qb��fq���5��{r!�N떆���^k����<z��F�5�c�7Zi?��.P>��/�b�#tS>��g���JIN�n�}[�U��~�xz.���[�5��a�|}���b"�=+��oH��r�<������ަZ<�Be��ã
��#c�5k����9��E^�y��u1�	���ؕ
�X���䂇"��t��L���2�7��Fm��K.����CQ�E�������2��eJtɸ��A�G��9"��O&d����[�r�39�z4�/�_@4�MR���y�öK;�H�I�"��E��[���:�
��VH�w��@Ff��Z}�/�Iٸ�c!��+�uʮ��}�i9��@��N����1���$�_Jo�xYȧ�jޮ�`��眺f4PL�!�K�L����MK�^��8��}�z2�;��au��&)Ky&����j�7�Y^��Y����A��_yw���h�5N�q�`����{�dc6��V{ޤO��D�a�We������~Y�����g>�r�[�;@x|Zq��r�9�W������{�:�Yre���r�g�e~����sOe͎��N0$D�$5'�͡���FYV4�<W&�2�R�����7`�Ms��$�()X)s���ĥn�R	X%p�뉤���A�؝�w���-86]5oUd>}+aC��'��ۜ�9�b�a����W~��~�.0��n7����<�Μ�G@w�晱ӹ�n"7�HgYlmd�.|�i��*ɑY��򨽽g�1�����J�ѧSN�@Q_a�(n���w���X���[��4�3>�~��j��e����^�Ǧ��`�l�c�ׄ�Ξ:�zYK�#�u��p���|=~�/��{�9��=a=�s��5T��wT��/���}ͮ�����Bء���o��I�w�mZ��_un;D�H�ّw0M]q��Ew�y8�8�$���7W�[p�X5b�&fb�V��zT��3".X㤤�ՐhN'*C�&2��d�T.)w��luO�ϻ[�zw2�c����t�>�����1Sw�� �־��E�6�pF��ӂ�gE$J���oۣ�/���ׅI��W����R�t�d�{�{x��f%:��AI]�p�2\�O�q�3_*�J�k��z�pmbA/Ou	m�g�o-q�K۝�޷3�3�Sݢ�߻�@�{G�d�Ȅ�j���6��H�z�C�Ro�¼j �5�R���A�{O���7`8�,���VF��y�N�|��ʴ[ͮϹ]*�z�,������S��pg�����U�Q���$>+�]g�ES�Ʊfܽ����A�b�[M�I�QÝ���]�iaҮԁ�_�	�rr{>�>�
���=�^u]����؃��q_=��vM<�S���+o�d\uz蕗4c��p�z{`o�a-->�F\����u\�3�-[�̚��k4ϊ��ڮ�ŷS�}�/z���t�~�Y�UJjB:{4Q/���-/�Ed����A�t�y�3�4����+��Xw{����խ܃eM_m��Vԣh�/T<�X�`�w����	�꡽��$w���%��o����7����M:�ø;.���>�!S�4��Ѽb˨��)P;�aA3'"Rf���U"eou�Me���'�*�<|�Й�2���~����RK1��$���m>��Iھp��³����GwS��T�b�����L��;�/8�Khme+L�$Vsv�ps�,����18�w�.9�վ�x�[���	\���/b�"���
-\�K.9�5�tԔ�K�w|��kVz2����vSF�h�-�nO�Z�&ؔ6�Q9��S��ff�]�ݍ��tn{!]��Ҥ@���[	lk��+&r6�`9GL��x�K!7	����j����bU�j���_vwS�؜�J��N�K���O<��l��:�ܰ�0�i3̍���m�2�Ԯ��E޴U��:�C"N̠�M��V��X�w�Պ=�T!W�5�����)���}��j�+���u��zR��ZF+ؙ7;lv���H�w��vF��X�c��m�x�8�V��I��M�l˪��ʎ��i�z4>�4�c[���4&qu�cluj�([n�:Kۺ!�)V�N�$8^�h�ƧVjo8��(]���c�K�SWP�ϥ��%������f�]Z�x]^5y��0�8��˭�,>*"��!ؠ�8�1qt-PK:�;E���7�]��5fs�h�B�E��p�ß_|�<v��p�,o(SˈKܴuB �*�}6�w��9����E��:Ӑ.A�¹��ɮR�aqQ=>�JG2[��ӭ�S�ivj.��{Kt�oa�2�.[W��:�;��V;Nmq|�.�CZz'�Gi)۽���)�T���Ec��y��J�Wn(Uc�k{�H�����=#l��M&ZH4��.6*ʔȕ�ʬ�e��S�y�{���5ڸ
�2ع�d���)��� �_6[M�����z��p��V�f6ۖ�V�-\iKU���Sm�89LDӚ���Ǫi��0˘[*ܸ5D�Q���R�ۉs�{���47J��tj��[s3"er�˥��*��r��2��-�s{�[�W.;�-m��f6��`�WXWZ���1-����������ʺ��5�h�0��ٕh�W1k�GZѠ
6� ���"���e��i$�d8ح1��2�Ɨ)S� �u���{W�u�+,DE1U*Q-m�k\�pm�n��i��iƵjk3WFi�3mȭ��"Z���(�S?�E+bpw���ư�d�C�-MY�!�N�2�J�f����
%I��$�U�����]^���:�E�m���S�D72oW�=�b�vǲj����V�Υ�b����Pʓ�l|��#}��u�>�Aq��n6��t������E:�7�K;sZ�{�zG��z�k�{,(�n�������9�n��3[d,Ks��̬���$���ӛWV�z��pľ�{��T�kr�W��-d[��lu���$�6�x�yqZ�*M�^+ԭtl�ʁ}�2In�3$;q_4�i7��f�r���ݑR�7/�\�mv��"�TnTZP��)��J����W��G�w�>��C/#M"��Y�����r��ce*»$�{�ޞ2E"q�>�ti�t0�3��³�ܛ2��ۇO�ֈ�,2�mё�Oz�<�5֘z��9����RXg�T�����pW*��g{b�3�N�bh����w��t��k�����r/��xpn�B��,.������I�]Vt�NA[�:�6�K��X<B�a�Q=��0f��"Kw���$U���=��l5{�k963Y_Q/��
�������yVz�~�I�:+#����;���٬��/�鱊g-5E�j��@��k��}��sx��y��Ý�C.9G�%ζ-,=Pk/6Țf�	�����EDA24B6 ���M�������G�E ��0�7f��rl�qR�����g�$��/2��i��P�Qy�Q1dpg�u��y �s�I>-ŘxA�����W�ӏ����m����l}���nui�N�sޙs�T��4cِ�=u�''T���s�\mZm�h��o�|R���=���ﴟFT2gv�yv\H(>����v	q�6���ޞj-��=x���Я��3R���g�S��fs����M\e`V�r�
��D�vۇ'r7����r�&�k��-U{n���@N��0��d� h�ej�
�=���~T���E���v��C�H��3�sRs�P5t��f��f��Nд�\�'y��4�'��^w��f��vx}����嗌��2�����$t15wձW��x��'T�'J��+U�lL\���`������w�!V^c�(�� ��$��ɼ�G��U��g��u��\�ä�Ƒ����^���ꗲ��8�Uj�<!Ƨ��	����3G�˨�W����㱜Lm���#;9�1I����P��VX��U��{�$�'�8�T�!S�\��ˁsCk��/9�S�H�Gx�'D��B�ɑ��VO��%�Oee�Mͬ�v�?L�kW�&ah�.��]9z��V���K�N�Pk��[|;p�xZ���ZI���W+Z`�M��&I8�
+��ꨟd��;�E�Fnϴְ泈f���0��k&��Ti�|�����J��������}1���Mv�Y�S�e�<Gu[�1?oMqt��=�b6/W
B�/���NEU�x�[�U
5����I���I6��-�HL�o��-T��+���\�T�i!��q>�6-�lQ�q\f�S0 �Q;�������y)�@�v�Ej"�.͵�/W{+�<�i>���+&Y���h���z�tru{��Yb�/@%���[����G^u��*�Ǭ�Z�ȳ�0f'`rrE�y�=��@�9�+ԉ�Z�bcy�z��Q�����2�R3��v3!}fR�qW\�scJ5��~U�IZ^�xa���ц4x�l���(0�=eW�y"}$��eG�	��瑩�p�l��q�Vb���M��j��^c������k������E���֑���}��g�ӛR�=A:�[�8���s#��D�Gr����>i��u#�揸�C6��5-G�*������N���PH�﷎I����)�<��+C�w�o*�	������yz�FC��ok-p7ב�屰��f���Q�0c{v-A�A>Q�2����r5�D@��%|w<�]`W�+�_�}~y��(eK2��k�O��ҲK�����Ƞ]2�ʘH������Q��T^5oQ�md[تp��J&u����r��.D���=�B��v��a��Դ�3>M��0`B��e����#UE����/�!��\����*p��:Y&E\Y���O�6>Z[JxY�5�XW��e类7F<�5�7�������w��껌K�I(�![9���V�\d���r�Ԗ>-+�΍���"�6�%��Yr69�F��w���~�kRg�[���D/���i0B�&��e���w��	�啩�w3�QfϬ�2��nc�Zʑ�^�}���þ]]R�i���XuqDa��ׄ?�t�Gn��$Ԓ���9toVg/��(�˔��pv�T�辭�η�R���I��/=|�n����.87�R7��h=R.~\PWzn��rT`U�Z��v=�>]���+#c���Э&й- ��Ѿ �~����=Q/Z���+��T�Dz�ۼJ����L]����<����f��yӰ�y���ઞ�9��'�xa��~���k���K;��58$��q4��m�<�m�a���O6����og�R�*���͸_27w�SXΠ$�f+�Ƚ�_lq�]��t�$�}{��\ju玎�]���ٍw�o留6`����-�^������:d7�e�(�jn;��r�����u+;�:��Y�u�	^�0���c[9�X������R�
��#�x��R9nb��ͻ���G��:*�{�r&�rr�����m�(�A^��RL���jKȍh'����g��Vj�0�U�Q�jzm$ǵ�s�}3�B*!WZ���6�/{��,��E{y#��>�F�)Z��B����2Z�Z���.I�״��A���y�YEe�Da���}HN���oZ�Ίz�u�in�fn�V�;��y%/Mvtj��9�&��g%ڞhA���oMDq�y�oY��Ns��ē�MR�n�9J��*���,�k�8lg���3H��G`�����:�]z�1Ň.������bh��Z����˙�_p�'1��'��{x(	i{+שv
�ٿ� ����G1v�G�])3Ie�� �!��3W����7��;�*�1P �𭚹��\\=s��Y^��^v�`ǽj:GJ��˔hpUSs)��L���七�=��z��TI(��t���Sw&�a8=;Ԋ�����2m����O9#�[ׂ&��H�ī*�ׯ�o���k|y@F�wH7�p������y�;qW���Ͳ�z��^&H�t렄';Bmf���:J:,���L:py]t{P�b"2��~3�8}Vy��x�?Ǫՙ�%Hl+�SJ�_�i��:�J�>'�R;J�őT\��I$�@$���C�� ((�(9�((����������P���9M��0���������'[:��D�<H`�-�(BB�( @�I$0 ���  4
�JƁB�?���WCw�Sg@YJ@�� 1@AAP 0@b 1���t X  ���  ��  � 3�� ��  ��   ��@Aa,�u���
bB�'��B��t���$�����K&�d���̆~� @RB
E"�6�0�fa]c�/���N��_�K
���4N��_�"Y�::�%��Hí5!�d��N%�{��-a�b�U/s��00>=�A��3�"
"3��͏m�ӈ�G� (."�*
� 	�����	������a�a���`!�H�\�O���dU����t�Xe9Rt "�� Q��_�Oeb(���@�	�c��b��f�����b��c�JJ^"��*���{P���@��,)�RP!/���:�����=�.֬G3�G�0(���A��l�ؓ�L(��W��[P($$  a�� �=d (t�C��BH�!<�]�X�d�
��4�R�s��cv	��5�?"���@	@?�B�!��D	
��) R` 
���A5�#C3���|H�܉t)X���9�rC��c�7��|�����@�Ci%��=�>��ziZI�0�(l;�������dTNO��r�1{�����X({����U
���*�Sך���(y��	v��&#L��t!O�w���z�pT܁�d�?Q�Lq8����z�*hvz��'�;M�C#$�b ���m���
�"�?I �	��� ��|���!2.}P\�	����/!�m..WL(m�$j ��C�^��! ��l����"��p)��$C���M�B!��tP.>X���<��^8�s
��BIR�m"C���8 k�H�jޥ��I���0:Ѣ���冀��@Q��G�3�C��jy��<í Q��=gp֐��癐���������K�������~��>����ے� x��Ե ��;��xf���tL��O:��ltJ����:�@�l{ϸ� �!�x�.a��  ��R(������f���
"F�`sH1j}����;����D5Sk�SQ<�椘�0��	R�̳P#����ދ�	��(^�<��a�$q<�&�S����x�#����e��Dk`�Mp@D*r���b� �R�S��Ԁ�X5�Ȑ�ByJG��4M��#��D��HJ�Lx�8��*C����@�w����� ������zz��: =�O��:���{���( ������j=���c��A0ƾ���+[�RD0yP()�`#� ��5�����ܑN$�H@