BZh91AY&SY#G��ݎ߀@q���'� ����bE�� �         ���}0RP�����+L#A��*��T�BH��&���B͒�P*��(�Q)A)Z��R��62�Y
*�D
�R�U��;5I*(�I$UJ��RUR�T�-��R�*�*�	UH(� k@cQ(I)L mUB)Q+ D��S �Q�*
������(TJUAP��
EI*HB�����)PR"���*UE, P�.})   �z�H�� e3l�*� )��8aFݚ�(�I��ѵS 7o�WC@�2�.�
�*P�EA*�)�R  �u�]���)�x�������EJ����@r���ն�O{��J����л��j��W����M^��{�T'f�l^���!JB���$PR�P(PP�:(� }�����JR�����J�����y]d)m�^�{M�^t���zj�,u�z�h�z���zҢS�Oq�T�UNz��z�V�I��ת��T;�!T��('Z$����� 9�AJ�S����֤��Ǯ���U ^���T�U ��{Ҕ����t��UAK�;z��Q$+t�ީC�J��:��*	<{�T�vy��RJ���QT��$ ����UAR�y�9Bր8;�z�EUW���P�*wJV�V�J�z��R�l�ڸ庅

\r�T�+:��T��s�
��V�T١J���4�I�II@�}J����v>{�H�����$�J�t�*�JT��J��	�[iT���Z�INSe)U(���t�5�J[����4�T���u����*I(��� ���w` t������i�  wK�  v�c@��8 .�(:���� :3��"��H�� ��$ ��A���� ��8�:-&t���c��v�c� q�N  MXt��+p �����$(P�R�>T����|z
�s�  v�f� �]�=���n  u�� 	���P9ɺ� ��� ���A�rB%(;*]d���Ѐ��@��V�'p�fj ��8 Cc] Ҍ (�` ۙc���
  (PP	 @ L%)J'�`�1 d��4i�*~#��*0    i�O&AIJT2`1� ��B�R�      OT��*��@ h  H��H���S���z�a��d�S�w��?H�s3��S��?S;H���g(���^U�1���+��5��y�(��W�ϠW��
�@EO� ���� 
��mj#���#�?���?��~��O�U@X��$�g�x� *�i���EO��/?������m��щ�X4��-�m�lb����m�lK`Ŷ�m�lc���l[b� �!l��%�m�l[`��6���1-�l[b��6���`��L`�ض��M�%1m�lc�!l��K`��-��l��bŶ!lB�L[b��lBض�-�[�F	lR�%�b�-�[# �lBإ�K`Ŷ!l[bŶ-�m�`Ŷ!lb��-�m�L-�S؅�b�-�[��[�l��m�[0-�[�!lB��K`���{*�U���e�f�f��-�l�%�`�-�LKb��	lإ�Ki�-�S �	l[`�-�1-�S�!lB�-�c`�m�l؅�bƘ��)�[�!l�%�`[1b�-�l[`� �h`�-�l[`��SشĶ!lB���m�l`�[�6���m�[�6���m�l�Kb��6Ŷlb�ضĶ%2�4Ŷ-�m�l[b�ؖ����b[ؖ���b�ؖŶ�ؑ�lKb�ؖ��%�m�l����-�`6�-�l[b���m�l`��1��`�-�[�6�)�[ضŶ�-�[�6�-�l��m�l[`��6Ķ-�)���6��%�m�lb��6Ŷe�m�lKb��6��-�-�le�#��m�lb�ض��l[bS-�Lb��6Ŷ-�b�ؖ��BضŶl[b��lKb����4���-�lKdb�ضŶ�`Sb�ضŶ-�m�lBضŦŦ�b��-�[�-�#��`�-�[�!l`��
[�!l[a��Kb6�-�[�	l�L؅0Kb�-�[�	M�%0Kb��-�[�#lؑ�[0-�[�	lR�lB1Kb��m��HŶ�m�lK`��Ŷ�m�0-�SB�
�P�*�P� �*��-�!lAb([[`"[�ب�� �"��E-��lAKb�l 
`�� ���(�E��P-���@-��l-�� �� �T-��lm���P-�-�m��� � %�-�-�Q-��lT�Q-��lm���-���� ��V�(�[e1�"��؊�[b�lblQm�-� -�%�B0U��E� ��V���*�[b+l@�-��lm���E�"��V؀� � ��V�*�ؠ� �(��@�� �(���� ��-��lKb)lD�b [[blUm�-�U���V؊��T`+l b�[[`�[[b�)lPblm�lضŶ�m�hm�lKb�ض���m�l�%�i�lb�ضŶ)lضŶF%�m�lb[�-�m�[���-�l[`Ķlض��1�[؅�m�[�!lX�Kl[b�-�[��i�lB�%�b��!lB�l�-�[��b��FlB��K`� �li�-�Sض�-�lض1m�`[�	l[b���c-�l��m�[�6�-�lŶ-�m�l[`��6���0m�l`�ضĶ-�-�l`SbS�6Ŷ�m�[ؑ������G��9�֧��rzoY���c�ݭ��)w2k���&�
�c~�oq��/�sOcP|���k(�l����f����g.�A�s}S�{�*//�.I�a�n��aN�t	�J��d6�����U�NZ��[Y�!5JϝS�A\/C{u��T$��P*��Ey����5��/2�	Qb4V8ee(b�#�����C�n��Lېy�.�~��w5�8}mu��$��-�U�Cz=B�e,Vdݰ�4�(o�m�[�������M�L5�ʧ2Ի��{�m�f6#�ݢ�����.7*M���X^����q<�0%���43]�'�A�2m�����������c�֨.l1)��
�����gk��G�`����������̇���R��T�ꉚ��o�SU=�.c^�O���l&�>�z�v;�x�y{OQ��z��"��6Yۆ��-�G�Q�c6
���v{P<���1j����-yO��r����p%TY7 �j�`3LP��_.ӑ2߫d��怞ϰ*�p���כ��� =�O� v�v���Qx�CHἍ'f]�e�h*9�7�P�Y�U]V��#k	ڠҒR�cq���7�X^�y��3m!��3P݀��UX7�]K��G��v���#�B�aN©���:�V���Z*��+=�rkl#^<��o�$��u_'��xuQ�0��T�
�f�;i�Փ1R̅�uB��*�B�����Խu'&��\�Ӟz X�7"��Y�)2Kg�S(~�4=g�(7O���
M<4Ҧ����֬s.V�Dp`�6ɇ�Y9�]L.Z�ίn���n/R��F=qj9��+n}}d����e�f�_G�Yj�^x�iڜ�����e���F�A��cj�İE=�G� ܸ��&fQ%R̨҄i��!)
�V`�L5h�
�K|�S���n�����AĘ���BkW<�0�W�o�/�6�XK"9CЛ���6�N5��x��O�jH�m��Q~��1L!��|g�y�OIŹ�$͇*@�t���<"��VVZ@�ЧyB���X��J�rh�V�<�7� _�Q"\�����Y�nSذ��oޡ��<�Y���f'7I˗ �{,;n��Q�����5'�n�s|
ۗ[�d'[�r?;���װJ=�q]x�ힸ_�V�u�qX��J&-ܛ�wDb8��X�I�{m�L�8�5��<�6-*��R���r'@��˩�`�H�*�&�����8s	����ߊ�����O�y�W�i�6(}��s_�n��4��f6�H�j�Ϫ58���75��5�b�m�	њ�kԫdʥtU�hFd0�ٓon�K�����6ӻ@�	R*,�d���PGM8�l^wP֙#)
�k;����/eӣn=N[O�7.�m��u����l���w�e�]�f^�J�kɷe�z�%+4�kf�/�%���eֳ28rg�d:���7��\�Þ{wX	܁2�Dk;��k|��z���-�c#S�}H-MF��Tf�f��R���,��M�m;��b�M�.h-�����y
p��cı5�7��Ws6]��cG����N>JB!�y��,�l�? �E��R��Z���>(�u�m�/��8<[�!�m������Y�����F+ɑ�dU��i�����Y�.M����&��6JR��J+U0�	c0M�Q�t�u�Y�D�H��)��妡ńmT�F��DJ�TU�:����<���G�C}m�f�&XT���i��	2�����CRx�w*��.4h"�/[7��S�#��a����2K̮����TM4J���|�y�l�-����/m�x�M[���f=ǋ3]���5��-Y��q�F�G��;��8�m�2�w&�tIC���H�X�N�c>�*��-����ɔ8�z��֫`T8VmAf�15����c�`�,�-6^Tj%Y�'/o�Ś���z$��,y��ә�	j�X�h�m%�?+(�>��n�OJ<k���>ٻ�T�|�ؤ�
j�%CFW�J[B0�!K-n���Cj�w����D*���2����tX���hGܒF�B��a�+l]�$%�	���ภ�֗�lܲ�e��Lȵ��_K%SS#ȥ�B��zo�~����;5B+��S�&MO\Xl�)�70ǩ9���_�i?53<M^J�tc�����V?V"�MӀl�]śN���<�H��Ո#�
��p8��f�5wa޺X�6�r�Z�f�����<�8�Ȩt��ړϩ`~�dۭ9�=�`x�]�hGRαK=��z3|���x�'��uo��Ռ����K��3p�٫wҏi@'�3`�y	�������9�
���(*�J܁��[��:ʄ��l�F��_�#S.H�:|=JE_��p�tP0����ͺɮ���D9���cMj�4s|�S�+ ����|���d�}��d�4������م9�m�."�4�&�Ɂ�6��g34�˘͋$hd[��v}��*�ȓ�Nb֨�ssqCkDz��.X�חsM�x1�.��2]��rkIO��ɚ��חvjh��;�_��Fh�ׇ2�|b^��dBA�mչ.i���~>œ��P�9��i��^�ᾘ�GS��^{p&͘Į�wZ��(�n�H�
�@ӶcƼz�_�g��<P�"c�)�����4-dm�u#.	X��x
���h�&�n�[�nyX�'�[��1�������[��ERxn��v[a=��8`d-�;��~��6.'3Y��g��u��W�����zd���쯐1y�4�9VIUJ4�.�7)Z.IGa���㩗e/�ݐ�,���֟�xX�15_�V�<׮�M�X�{э��M��
z�kl�l��XG�2<�z��%[�a�������Uު�1�3�b-�� ��V0[�����J����ڒ����2<���2�c1X;*V�(;�V�X�V�Z��XrS�i$�^�VhU�eK̳lI�P�ӔBף,�r|��d�XL��tel�O��	T��%r=�,�3�Vi�4��0�R���ْ�i�mH�r��u���ZʹV�A2b$�2m��+X��'����.���S_�-E8�i�"r-,�@����وy�se�)����k�ܕ�_DF�NM�v򩕺�G�nk�i͐�e5��3r�-�hT�vÆ�/mY��aS6�k���5���k�;E{Qx���^z�8�y��$2���]j�
�]���I�@�̬�����p@7�Q�����x8��R0��A2������G홻m�Y�]�y0�t`�m�{uw���j���{R��l�E��;-Ɋݥa�����H\��U��MU�5���FS.F��v�n��P�9��e#�|���>�|��b��kx�_`�*�3�kכ)ym�W&�a��頠��p�TD�Y:u2"����y0�v�[C[��*�!��d��Z�,����Hf�GU2���'��g���<��vĝ,�����Pi����S���e`6��8�Mˤ�����75}'ح-y��YS̏��V�q�C������.���	�`ɣ'�Nc�[5����\'��[�E'J��_\�'�*��<v:�vC�m H��&�S�_���T�ՠp�(!��*�E8�7�����i�^�-���˦Й$hH�.I���!�Ti^G ��ձ�7b��8��c[�Ij��r�HV�;#
��b�ت�b��˩�f��"w�b�Sv�e��w|�36m��x�C^ϋ^�����wͼ��U����Z[�\�%�El�ǯ=��1=��!\	jȍg7<��9�£+m �Kl�{e�KeCI�`�F̣��Ѥ�Ƹ�r�MI/p4 ��S/�F�w���ɏ�Q��aŠf�nyXq�����N�S�R t�(Բ��`�Z�/+
ڹfUt*���T-��1*�xKAe
��!�f�iZ��=v9�`�)v��y�O���ExS�L�8��fz*�	��dC3Un��yUJ_�j�ʵ10��j����Jbe��4x���@��t�=w�I)���;\�����{#~�yo��SI���`�����{���Mٚ�Ÿ��F�1�o����<ߊ,���ޯ}5�Pwn	N��g�;�=.����D�|���@��ڶ��f*��/��paZ��	��;{0O��-�0�WŻ����s[̥-8�[n1-���=�Z�M`��n�!Lf�LW|�g����LY~y�d�FM0�(��z@���G$/����0g��+<�W�#���y�~N�ۆ`S%<̺�S�O3 A�m�6hYX�,�v�v���jS��$�B�N��ֱ��Iǐ��MPƖ�J	n��ah͟M~L�&��7���D���h�i٪2<�14��0����i�7�����q{����F�U{�l�l6U�F�l�nѓ3#�,�̰n��Q��a��2�{�Ծ�����6�i�1m�hm��꾒\�={.Wpk$�Lk��p� V�^�)��F��^�]�P�A���V�b����$@����4Úbp�CA��S��2��C�j&�&ʂKNe�R&�K���DŵGtT��e����xLMaѤk�`V��Q6f1�sB8Y�B41�-:#(H!M��x[��|�79>�=�#_��=F��F��7V1�q��tle��ߟ�����vM����m��5��{/���NZsn�����X�U4G�|�\fL���-w�̾9���ux�R�k�d zA����;�"���W�����<G�����̌x���KV�|�����j,�&YyV���P�Tmej��@�z���v�ڥ�lk5n:�;��k[�5� ���ǯA)��}���H�(��l��=�]�VQ�������L�q9�N��i���/�C/6΢��l��^h��^avd�<�����m�wѽ���i��RD��XeB��Sy�0�i�$�y%ڥ�Nˊ���8hGr�;��B4��U�7�
U4��v|L~-��dR�-̔3AYN��Ă�(��6��Ds*0���Kz�o�K�m��F��v���۾�a�{$�k���s�q��{m��n-�$�hg�e��7n�&n�0����W���z��8������$	*K	'+J`�;c�� ��Z($���|��i���x�K�k%�ZʧWj0U\��0�(�b����Q��I���@תZ�h��l��i<�����{q�KJYS�!z,�)��V����wF絠�'&OJԓ>�U�vmZh·]K���z��V���1�ط�d�5�(a��y�&���2�&5J�2�;������iD�[��K|eH;@>*'��!�M/���d˦�^^��`%)�ŭ�yFM���z��(�l���m�5��|�}��dm�w�3c��E�i��Z3m��f8��hF&�y	�1��yDw���q�J�7*���:kBV]n��6"�t3w3"����3j��\8j�4E!�a
K���*@ۍ���6�m�f���v1�(I+�^Y�r���cwkl�o$&0^
��L�;�E���R�>l��B��6�SE�K�*��iB���v�wR�����p[p�tq���.S��B���IPD7Y5ۣ7�Z��$�q�K͛���n��n��+��\�r���q�V\�K��KZn2�٧�G� ���7<����ܖ�u9��O���^�5(ܪt^�ׁ�B��)�O)�4y�M��^��4(a�e�Y�^�ƕ+���Z�'�)(�)I\�&��v�'��-wS�Z�]j�M-����S���C�2^*��jU��l��˅���.s{	>6�azo�|8z��N�s�$2'!��3N�O�)���J��Z�:�vJK���T����|0��v��58.f�d���u�3ډ��'�x�@�Y��d�m)����H��� ƻ�Lh��UҦ�+�m8�I냫�کY�%jj�K'��qT��!���#!�&d2Y������ІC���U"Ҥ����I�1�����a��6���ᔬ9H�q<wߡZO30��5�i�쯶�D�I�qD�I�p������+J�d�H5,R#��$�8KDxjͽ���2�G4�;��t�+O7@�Fc:���Y=����j����1��w�3�'�%��=��N�K���JE��;N"p�u��e����Æ?eG�ú�3�M8�H�b1��,>R�m�>k9[X�䜳�Ƣ@�$��m4��i�1m.�h?-��-r��&9j�6����0��&���ړDK����D�T=��H�Il�d9�B<��ð�'I�R�rY���N+i�-�	2��W��l���	�M3!P��M���s�2ِ�=�8�	�ip�9��z^I�4�L뛝fq<U.�&B0�/�a؇d�O�߉�T��aof��9���Y��]�J��#NB{��m�5܅onB�L�-�OB�=Jh�]˲��i]���\�	�A<�!���8�B+��0��ܼA%��<)�IG	�og0��2a�s����X���8t�8E){�ͽ.�9�و�\/��(�Bj;��ݶ����oR�\����2��-8�V����.��/�3��&N.�K�)Y'y�<VI���{�J�I?�xfI��=R)jD�ɑ�J�=���I��ҮN�i��lW��gT;js��m)�y�s^%���*o�qy��s�/$����Sr��M�N4�ā0�E��S�����x��c��I���}ļ�c=��ݰ�s6L�6ր��$T�ٴ��RQTT�4m���)ߎxu�+Q��^����$�%��O��&��Ի�<��L��M���@?����;�xH�~���M}��dU�N9gʺ�5��z�a��;��s��I9^�C�G�}�kn��07T���#�������Y�/t4i�C��MWg`��J�n���O��=;�y"�Z��tOY���g�F0 T��7�+���2/v�ޜ�+�;�9*�y�{�S~;gQx{��{�u��� .go���ݧ����%�Go�!t�
��w\�ch����7<(z�=����TE�t@��@�3��|�K�t���Ƈ�J��T{8۶�0X����`=��`���݅�WF��0�U����0���G\�S;:|U���A��vǑ�<��ɞ΍��]!�$�AY��@z�pa�kNy,&�Ce�.��?A���2g��0)�d;���R���D�렪�'7t�0���9�������.��=gv����l8�x��g��d��N�\z�U���]�6 ��DH�	������:�����褹wC�h}��-{�W\���7ЮT�]!}X1�d�a}$��>]��Ǟ~P�{-�yC��F��W���"��٠�7�=*u͑�zs/�Ur�o�,:��Z�{��������M챇��W	F�ۣ�!BKn�U��&p�z�A�[��]ܵE�㪅�i�PS{�R�L�6WP/�/g�t:�lr������V+d��=Gq�]�E3$�{DPy�w�/��S^��q;P+��Ŏ�0]�!����{�&r7h�a�V-9�L����2a'&L�fc���싎N�
�I�x:�1�>�+D����4���ިr��C#�UP������c�.^t9�?n_M�#*.����ॵi�>F>����p!/��q�>nqÛ�^��X�w�5�]�]����m�}�xj�$�����#��T��G��续Nox�F��M	��/��w���fJ�?73�oeU]�X���;�/x\�xXp��f����]}��Tw��m �}xB*6�E��#��w�d�0���Gۮ�҉˽}�5���S2a�1��o<�"�W��rb��0yt�����l2�ۃl�8���=�MU���m̼yy�l�=XݾK�ݖ�a��48a������={��{R����M�#E�Xر���2��"��#;�q����-�I	Q}xH��jG���ҭ��/0u�i�<Γ�l>dc�h�lK����t���*�2���Oa��܏�e�4�&;դw����D�Vn??r�S��1�tSL�Q�q51ុ��P�.�e��-���^͠�K��o�,H;}U�{�<�[��+z��X�Oc�����v2�۽'��mu�Y����Yp�Q��u�n��W��i�v���w��cny7^T��>Y��I���X:ݦ��m��䆞)��΅`�,�'k�=�-�������O�M1�ʸ�S���T��&���h�b:�����$ޝcxo��4N��#��S=�I���g�\���[=;�$��U<tX[a���s��Oo�H=�c�O�)�^a���O�SS���e�j^��6"�򺟳���|�q�[|y>�S��qݜu�r�W�����]�񏼻��[u�9z��3�{L���vf�yH�wc9����a�ڞ�V4jI�,���K$�c�.r$F�#��bR��+W�p��Y�í���IL��i��v:̕���7�-,�*_�T��{vg����9sR�ݾi����ii���:%�;���V�|+_V���h�ݕ�d�jz׳v0������&_b��(KӜ������3����j�����iAȸ�Ǖ!�ZF��@���ǳ-S��A��e�/"#݅-���ĵ��-͛n����5AA�ܽ�3����lDxUG�֡|3�U*��L�2�X�c�8����V衐=�J�a�Gz���-�xV�{T�9OP�����̌父�����I�Pe��Krj~�~ڄZ������!2���V��p��������G��x{���g��I��U�k-�n�����R��Q~,�9��=G�Q�5�L{�<fyB��ݗ�����t[^;o�����҉���̾���*��k3�~X�@�XY:���P�>��p@�������j��^j%���o.O����ڙ��t�"��
�b��N�!�����$�H��d�+.F���ג~n��#|����_e�l�x'd��p-x-}%~�~��g�����z�̹��B��PL�&p�]�o���6d��U�G�C�1(����[ӻ��M������S����'FG@A�X'�,��QC6��3Mm�&M����~��k�^�����d��E�7��a�sөFW��B�*��� ��\ϩ�+��
�nš�n�fN"̯���<yS��S'b�*f՘�>ê�= #�A���f�3A�"��w�G��{�ay�p�<r;�H�q+f{�TC�]2S&�����v��C�k�V�T�b��'b�-���h�u�>L��fKv�O����LB{(���j�^������[,qs/4�Yã9sN���K���>-�4���(p�<=���g�܅��S��~��;e��j�ܢ;���3�M�o�8���n*�7�[��dV2X>��ĞK�Sh=R�3z�U˫�K���k�}�7h��n�>3�Y��b�g���C�Ux����������8<�n�����1�yH=��ykނ.4,|�;���a�����r��^�
��)L��ٽG������~gx�74s5���FRB�{v{r�!�bح'|�C
YvF��Yգ�A��C7V�ݛ��=N�P{�]������-k��"���s���gec�B��%m�PayŪ�3��ua�ʝ�˒=]����D�_������7o��S�5.2���V�C�����n����z����܉`���:����{W�ŽWrN��������ϕ$l����Laoj�B>�5v�P��hބ��NM�Y�G�
r��rb��Gf�l����r����|`���l�ߎTm �������D�0�3=�oY�)����f�#��9n��{1��٭y��R����[�ٯg�4�Q{�{�����B����y�*�$�d���+wҭ���o�����2���t�����t7^t���?�?-�7�ۣ��_m��vrھU[TE�ƹly��E��m���b���ܲ��:��g}�g���/����Lm���н��%�#�������]�B�<��$Agz�.����U+�@Ʈ��0���{�������567���s3;N��퉑����\�\�}˻8��uL��U09�ʇ�p.��͚[���]QYʕ�����y��b>�v��^��Ӿ]Y\I�8��vBB��]�Zr���}���=0m[׏���
�.��W�z麭�W����;����&r%YcZϒ]��ݷu�9��bN�Y1P}�����1i���jY��X�%Y��Q�M��:��@숓 �'�%�&=/�n�[R�N���w]�g�HF��o'�c�t�.~T6j�0��y�e:�(��x��|�>}��2U�{Jj�֭�z���7�xV�I�^�G}���lմw���k�
�,՝��ݾ��e�ޚ:�r0����{o���u������Y�i��\�-�1N�q��1k��Î�=ޕCS6�r�j�T��H9��W���F���u���䗒mBQ��[��SU����^�u܆�gMɪ�ž�~mzJ����_���鹮���$g�)Tk]����
�˾$�.j>[<�c&z��k������vu��=�g`�q\����œp^P��˶�n�eM�(K�e�.��j��N}Dvs�!wf".���-��w�&��i�:t��t�B5��k|1�ޫw%]6	��:��XI�ͧ���s�c���"ⓞ��bx-9��}G�k�A�w��5j��U:�(���[��,s�^��ME\Ί�	0��+e�r�p�S)�rX�8���_����T���rx����oY�c�-��/jM�2���r�PD�wڵl��q��������Q�.m�3�w���gdv���hL�zk�;����^����옙�y_b�Ӡ�GtF�e,�:�n-Wܢ�i�Y�H�n#l1u��FC旗@읒_I�8c}�0R���t�ɏ�T�/�/���j�w����y��ڑ�Ƈ''1���Q��G�<g�<_����h�48r�'�ۮ:S~��#�g���U.��4I� �͓_���kk��Qg���Z&�5��];p�*{���� �{���>�>�Ӱ���oeM�;p��{=����"�JԒ�բ��!���N̐��=H��1��N#T�jcyR�(���y	vX��[������9�ElN�����4K[h���Ք��^�"�6���z~ձ�y��;�a|;�=6�A���l�??��s���]��/,E��w�n��b��1�f�$<M� �,y��{nSU�ꧮ�6q�9�߳�f�I�ݫ4�a�0�x�w&5ӭf�8˯<L�&����j��7�����)�'	�a���E������pv�[�7� �َ1��=��te�3�e���e��{������:V����K�(��"Ǜwל�{�s��5���*�u����r^��y�wDwS������9eÛ,CKrAe<�Κ����}�=rH�M��<�8�����|����v-�;yACb����y\u��#/�/�Gz]5F�]�}#�Niq���j3^��h�ֺ~34kSj-�+�UX}��浕�eg�7�����C���܆&�5�`����\�o��-���[���jO1��Bt沺Z%���P�8W	Z�����Ww��vv?]wS.�u[�}��{�]6���᫬�t��88v�z�]�|��쯘�Lv�L�d���~�lY�G��_'�Cs��7��W��%\�Gyɽ�v1����^-O�w�a����Cq���k�D�����^��ksC�u5�^GbQ�;����~M�^jw�܍����tb�zs۔��:�,��t$n�(��<t�KМq׽��yff4]bp>�@�ƶH�r���1j��4��X^�痉ތ��K-�͜���8�w9;I])�3��7$��{�S<=2R}�����֍L�<W3S��s=/��Q� ��6.�?,w'ծ��K��b���L�sh��ٔ�\S�^�d��	����^�3�,L�uȚ�V/>�2��t��Ʈc|3K��|�v�=��xW�����W3��&��3���x�3�l���zG�m�vl@��i92��X4���&�k���M<�=�,Ue���g�������=Ң�C�Nvz�:����[W�ɬ�Tn��ѭj�]q��%u�x w^���o����Į�n�F�nL�_��3{�F3�[o�������ÕhX�C���kլo9{y�zr���I;���Y�aj/j@���G42�d7xE^��ZD�<��g���$���9t��a��]n�U9[F�E,v�s�u�(�I�*nu�h;!���Dv3���.y9��!y�vӗ��46���O;=����^��X:�1���y�e��t�;�ٖ�_�}���P�:¯�[�:�s�3�ιog�|u��o��ڌ���b�q$w=Gp���kb�t	\�p[�w;o{��֮s��}�K�}_�,�eD�����'�g\��܇�8N��͜�J�fs;y��w�6�t���]�P�Ns;7�����Ue�/�������>cۖǸ�zk�c��pɽ�3��Xgv,j�,y���oz��\9��uѽ��A�ݺ�z�s�����v�ȹ�X���SØ�{._m�X|�XΣ����7�`��ׁ)�wwwKz[Î��ޮ�=����nN�7�{�M]Z\���y���X�z��>�<^^��K�*jr����O)M�y([��U���S2�7* I�+�;��E����nf�͐��{2\�uU:k�{$�S�Lߗ�y��j��yJ_wh����"h������2�)Sȏ��{��"�T��ӷ`d�Ԁ��מWb��3��w�����牸5 >�$�uڨg����R���b{�u.-��N{����/���C�zǼI8Q_;�V!���J���R ]J�h��Ծ�;/G�{��v��A�C�}�,u��@�֢�� D���3T�bdI�9��y ި.)�d]�����B�[�A9�I�h�/�!%�V���CȎ�^n��ז	 ��_hI��`�tW)��L��w��P������?���DPT>������	���� �#�?���C���O����������f�O�SWJ]{k�r��`U��Tr=9*uZ�y[;����!|7�[\7��-��h�{2�������Vc��h����t]��==��Ov�m]9��T�V��}�i�K��߮]��}ޘ�U9��:4_^�F0Y������B2�-~�}�BC���OT<1���ik�}
�aոה��RZ;��qф�%��Ve@gh��0-tzT���[9i��|.�-�mS�\�����PC&<==ӝ���CW�p�f/L42fd�+*Vv�K�(N���N�j=�r�sY�ﶺgf��Ӳ�_K�&`�Y6�Lh���#6�8v�AN�����"#���cm�1�3F�z�i�����{qķA� ����@X�3�7 ������d�{�����b��_PW��n��ܺh���q�|�D!r���(4��0����\g��B�.��q�B�NnO,}z �"l
�r�^��l�E�5��Wi��'��y)z]:6�YL˩]b�Ҭł�����Ϗ1���P�ӛC�c}�k8�2﯍X8���Ϯ�:�(-�p��|-F#Ċ��ʫ��m���{�h�w"of��&Vv�~h׃���e+o��rɭu�~.��@�s�����~?����q�qǮ8�8�q�q�t�8��4�8�8��8�>8�8��㍸�8�c�8�8��q�q�q�8ӎ8�8��i�q�x�8ێ8�;q�m�q��8�88��q���q�q�q�8�q�q���q�q�t�ӧN;q�q�q�8�8�8�q�q�n8ӌq�m�q���:|Ԭ�n�§�<ߜ��9�/��YX�M�>���)Vo�{�%t���p�s�pz�|v��5����R1 ��Uu�B���T]���3��+��`���f$=^d�"f�Y��)&�X�0.}�A�QB�6�ֽzGD�y]�&��1��`�8�w[�VZ�U�.-���P��	�&��]�y���eV���+���7�|���L��K����]�>�ۡ#ᇯ���x����ѹ���S+fu�u'W�y�=o�U~"���W�Q��G�!�g�G��w�%3��]s�!�h�.��K�
��Ӭ6"��L�٩�>���<����n���o���'&�·fs@)|d�iEX�[�AZ�k��m{$�)�N����o�lJ���PcW*���Q��5�o��y��{�Ɏ9���u�OGyUW�b�&?]C�o7���70���n��^���Vy��9M�zc׆����YY���鯘�.|O>H��@��.͝����Yg��0iYw��"z�vU�r�Cy�/a���A�\�JIUK|�a�g�_�eM�9���W%��)�bQ�C:+Y�_�M@�{���mu���׻�gS�]ic�����L�f�y�Wo�><v�8�n8�8ӷq�q�8��8�8�<qƜq�|q�qӃ�8�8��m�q��q�8�8��8�q�qǮ1ӎ8�:q�|q�q��㍸�8�<qƜq�qӎ8��1�q�z�8<qƜq�qӎ8��8㏎8�:q�m�q�t��n8�8��q��q��q�8�q�q��8�8��qϗ��}�]8�x��}��Gr�k�of���뱖"N�>�.��
�	Ur��y�(ǆ�ָ�}������D���їl�(����i�K���0|��3_]��@��y��W�x�^���s�� �IV��6�9�Do\^�*д�IyFd��{�!	�)X3#����i�x��o5��d,�|��� �zc�oT�o����.�W�+�8�O�S�ug����c��h��>�ܻӖ�Ϧ_+s�/by7�ۘO'�;��e�������s�n�U�O��A�*�o��뺩`���]U_�
�c6��L,�"n�bQ���(�ա�4����z��bu�!�V�ަg��S;ǖ� ��4�#x ds�sp)�f`�+1��f�x�^�<��!��=V�)��Uݷ���v%��Uym���+A����宭c����s\���y=��:�}2ּ��Ԩ�	3x?u��s"e:<|+��S�v�n]k�oY�y��]4f¶-* �Zl�R��P��
����nI�X�mv��p5ZUU]�4**��]��aT�z͝�]O��q���|�.��u��]��ZW`l�	%x���UW
�T��P�R�f��V�֥��ַ�7�ۏ�xǮ8�8��i�q��q�8�8�8�q�qێ8ێ8ӎ8�8���q�q�4�8�8���8�8���8�8�8�8�8��8���88�8��q��q�q�q�n8��8�8���8�8��q�q��㎝>>>:pq�q�q�q�qǎ8ӎ8㏎8�:q�8�8�=p{���-����$��6�&�E���>����F�������&�M�����q"��5qf ���+%Tκ�E�" �ᙑmmQvE�l�N�f#�����3�yS~�����1���5l�ayj��>��J�r]��
sc�O��Y�<<ЋA��}�tϷ �ς��T�����{4m;�^+-ʲ�"�'��3��<$��q���r��?ЪXO��t�;�sŅؗ���Zee�>J��<X��躚&�~��Y���}�����&6�z�wa��5���'�f��wΜx5���o�����Lk�g�)?�[��<�G�qh���f&9��*�p����O>�X��\%���3e�]:�H5�紆t�({�oA�L�2�f��U�n�n����*{i�!�L�����}��Xp�)e��&����9���6V��xnc�0�r��/�.V�׬c�i�fG���͜�O�
=��F.L17�˟@���=}�9C�o%��pS�ȾS[���ҔOn@Y��!�x[� ��=G)#JVyʹ��t���@u�C|3�yT�'�<��]=TV$�*��+������1�WnJ��<��^��'ާ��N������>�Q~qg��[�pN�U���е��f���T�+����t�5T�p�G�c=�p��w�K'���\��&�rL�Y�b#9�p�K�0��n%.�m��;dR�꺺(M�Z��o4&�p;��c�׷2�'�N���"�5����Cwuˬ�V���^��1g��W��*�s����[wY�'�D7ɋ�E���k��<	L��r����'��>�a&;��@����s%����$WE>m𚯵���l��� �<�W�L�Bg�x9�w�9A��Yս�e՝����ԩ5�Bh#��d� �ggdz�ϑ��;�B8h�v�m�`��{A�F#�F��0�'Gwz�O�������GhKe\�m#��J�5SY��A��wxpD�gSq��N�n� ������>j��"�p�:cJÚ����U������~�~[����=惡.y�� �;Ʒ��r��s�؄�}V��>��l�����:�;r�HΑ�����^�Q��̎y˔��Lm�^�V*\�C�a��xnW���?6�ga�
<�j�eK��78Hnn��f�$R��)?G�������緼��St!W$i|�~��(�'��p�`��9g��׽���nZ'��
���'�j�Gz�[��4��b�m��<ܼjm׀��r���� �9;|�l�鬾ku�vI�"����7���[[�>�=d$D�l��Lq�����o;J�WH�*�J�\xe� �4���S���<^���$���k�q��{3���P�7��8B�p3�X]�3z�s<�Js�Ô�n���u��Zȼ����z�>Ҡ�䬜�h���˛7Z�tN��!M�O�&:A����hf^�d��x�o@n����ΐ�����2`��{���z��=�z�^VT�� z��7�J��\�j����ݕtDf���X�rG�����Η�>zo�X��
}�B1�z���x��S��
�｝���I���p����JN�Z��q��6ؤ���/��GUW���U�u��2��7*�[�ΐ�t�����wc�xL����.]����E�n:G�T�h:L`5�s
�Y�=���[���s����=n%MW���R�[Ӌ�[�x
���ɕ�gz�}G{|�YnU:>S��]bg��p���7��p�b���
{͏��x���JE�}�-��g��`��;]�I�n�%a�<�0N�{���"le�p��;}�u}hkXq��9ct���=�Lb�i3���S�sk�Y��{�]�.6zUp�\.L�v�T6�`�	��{
+�r����P��R�;�|���k�.���XFqѬ���(�k��nQ<(򞙛_i��>J���D{m�<���A���$T-Vlۧ����7�ζ �goٙB��d�>�=��{*�qR�p���fu���d}����;���|��{����6��u��Z-q��]��l�����7��(I=s[����{srp��t�6�kwh�u����?x]�������,���Ӯ;�H�7ǭ�j������`�Pw��{���U+M�ǳIQ�>v�9U�P"���=uf�d�m9}��%9�f`�F�	2un2�\G�p;�C�$���=�����XȺ����CY�#ko5���L/3o{}�)��\�l.{�{��+xg��GTr��]Z�X4��Jv[����姙��z�_)py��x���'��t���h�U��\(�����TӘn�������r�6e/>��01��l�q���\ul;|ؕ"�S�i�Pr���)Uf!�nt��B������a&�ꓣ�}xa�lK�c�]%�{<&lo��e b�N�V�� ��z����,�(�@���s�~�p�b�&�����I�\x��̇I����]����B#��MI��V���ۘ=9p=�j�o����l��Y��WvQF��G�R�UC;n�����}�=�哗�����g0�}��G��¥Ё��o[H��Le�W8��:C��gP�w�,�,�F�j��V�l=u���q���0)�2DR0�I�L�z*����]���W7a[�uI� (�Է�us�y�Sw�>�7e�r]caޗA-$od��9�j=�CӴ�9�*�N.KSt�*X���v��/jA��ؽSjN�,ʭ����׾O^k��=��nnq��1�vsx'�M��>�s>���t��E��=���|X�}����Y�%}lcۄ.�8�����͘�"� V�,�:��gvM	_���W�q���3�YlͰ�Q�v�2��{��i�^���r�.�uY��oK�lrnKX�)f��]���q�$~/��{\����<�\8��u���ێ�{��h���<��n�<�Z�����U�*��ּ�h���o���lb5�l��kiB!���ڧϟZ��r�!��^�πh�U�����{���]޾;G
(<}��.��'K~W.��N1`Jr��o��x`����/�b��uq�+i����K&�����(�ՙv]8d�vGX �__=�u���$��;��}3CY����-�[�>SK�.�~�g��iU����2+3���PZ�ͅ6��F����(�-�S%�|�.<ɝ���E�R�w9�$�q\7`=�I��彳.0��l��p^�<e�"]��D��M����6��=���{kf��W}��r��d6)eV?MMk'	�*F���O��WMɲ��(M��򊹷ō&Z��+�L�8��W��wa�PֲG�@��9��د�Ř��0�J��&6"��F˕�ݗ�n��h��7G(ϡ�f!��&gM��W� J�
ɣ�|�q�R�6�h�j;ƏoMߣ�zA�«��벏IۚM-,ci�r��T�GKҶ��^tDp
A����v�~�ė&��|��xQ���}���x�k?:u!�:�9 �K��kՆ<,0�i�����z��#��V�!�q� ��G[D�\���3���G��b��J�ePI���đy='�ܮ��{���Tw_��<��g��>�ͫx�!U��T���)U�,��7C�Y�8)�z�6��Φ�ffBCx�}���܈<��}�#��[�g`]<�)k�upP���.w-6հ���}�8��?u��s}q�S ��"�=&�x۷/�t���u� ���u���]�b���u���@J0�5^�e3�f@���9�������q��������A���юKݑ�n��Ձ�]��K3�KT+eO���}.NO������ތ�O�f�y��v]P�Ua.�d��alⳣ�7RK�=��;�[ZQ���oXu�����w\(��tN5{N���yy\xs�b��� ��!V�>��"�y��(���h��w^GCe�uF��;�y�����2�N�+�Tevj8++�0]òon����`���:��m�v`E�ݾ�zW����*��E���[h��3���=YV�s$����}{�!}�T�v��R�������m;��+�$�~x�Ȟ{>�֯z�qz"�n7O�=UދGw�6��o�;՟��RS�gKI>�P��ޫ��4�ހf�?�[�&f	V��¼�[ޅ���=i�B/]�uwOe�����Ol�^5G;�m�O�f)��[Ń�S�����uNgr<�%:]1�׽2˥CN�ӗ:����r��&�&n&DwM�����' 0�t��|�w�P33e��]��1j��U䯅d���o���QV��Of�H"ZՌwh�,��c�wl)'�ɨ�Ν�d7�3����](&���-ٙ��t���;������\]B�C'���xm\�	��y�wa�z%zSb�s)�x�uQ�1�����ZT�=�+f��`�i@��-��3,sr	}JC/H<��ܳM�/̮��o�_�{��}�� U�����g����O�_���߿�?�?2_�n猈� Ϣ�H��*!#��IP!�C%}�ETP!RBdA�	$XhHAl����a1M����U �����Q-�,��$�Q�%2����j5!�	8�(�H��J���B<JDH�Q(�
,b���CD8_ҘI�]@crC
B�L�l�*����fC0���@�Ll�q���5RPi$� �F"J8���#� ���$�r4b��7!�) � �lQ�FQ�KT�A
-�l@�!��"�7�U?������ވ��O�[Ю��fY����u�z��6=y�Gv�k���������.��@n��g;|6e9��e�k~T�Ts��J�tG�.?���j��hAj��r�26ʪ�����{�������6��N˫Ȯ�_Ї�x���y�^�֤�����(�v��י�%��s["oP	�ۨ���_^l[����m��M�V�]%�#�:$�\i��Z�	�f%��k��psq���g�����`���כ[��Y�+���&�����q
�]Y��mf��8��j���`+��-�����+�>�S�⺴���� ����ʪ��_���׺ۖt!�d���쾹��MX�@}�V�]�rQcY�<ܤ�����i�S�'쀇*���^Yu%i;K�ʖ̡,p��'Ǜ���z]D~&���$T���&�=��H�����/ۘf�3�����V�ϛ�)ܾ=^+��.�M����UW�
��FT����x��-����Z �.���C\���Q�`x+�D�������H����{�G׃G���o]�{��{Ѷ�W����ΏS&|�;ʑ������9G��9�v�C����(�0��e��������W�#"���-���$"�(PK�P&�e�"3]j�6J-@��1DP5��K� �l�J�&J!ω2DY IH�hBI�A""$�P2��#D�LD>���%"%"ؐFL"L)�l�����!o�Y)���6�@Ĥ1# �t��)� B"��D*dP�o���! O�)$�[L��bG�!�wT�In �H�	��	@��a�"@�EzS�(D!6ˤ�F�U�AD�$�CF	-��2c�䑒Aq0�S4�!@]3#E��B|�(�D����P&�e�"0`-8~_4D��\i6����ϋF6Coe8|�((�≣T�K���iȊ���32@�Se��(&���¡*|�l$�I2Lr��$Q!|܆(IDI�jF\O�"�t%G�M�dP��h7�)
f���4�5(����_2�M��B��C�PB2��P"L(B�lH!L�����%"!� ��M6�n�$����HhyA>�ĺ���
�!R�IG�����7���^�z=z��8�^�z��:t�w��A���^���$�O��'�)��*�ۧn8�x��q�z����4��焒謪�宑>w��E��Pa!$��qǃǮ8�8�ׯ^�8�N��]UJ� M��,�#)\���cE%���5�Ώw��6����`أ���#��������u;\�w�W���.Wv����g�z}u���7F��˽�(�u�B��c�7���5n�۰����yr6ҕ��wMk����F;y��7����j��P�2��t��uk����}��wv��ܣr����7��������n�7�+wuӎ�Y���]�W]�rOMn����/_�{�������[S֏���k/ή�λgs�_o��wr��=�r��7��w3��|����[�^�/����k���v˟H��v�T��Ƕ�۹���^�pw{��]۾:�w]��O�k׮N&w2��w9N�uu��=�u������&���;�_5���]\޻��^����n��]K�B�w����o�	v2��;8�g&iۮW.�ND2���o�\�w����=��@�_6b0�c'��d41�J cp0�D��Ŝ4Y2�P�a�Jׇ�|�<����Z����uٹd�����سWoo����*(uA����\�ޭ���5�*�M�����Z:�(���$2Ci$qȓ(�%�p���q�AnH�O��4@�Q�"��X1"�2BS�3lFE�`�Qh&��'�Dc	(I0$n�p�-��8�M��!W�|~?�����桜Mnm؞��*�n�>q[����h��ߞe�/��_s���eɂ�\�yJ>�������z��E�Rz�4{kv�1U�:���Uє�kۺ�{�V'B4���cr�������"��aW��J���FḦ́�$@RL��f��X�S�W���]�ɴ.��߭�C��Sb�"�̄M��L��l��x{>�tO��W�q��5�m��ή |<��O� �^���V^wI<�o}�������Ps���GG��}��W��Y{Y����r�x^=��4�[�"ei}O^�l�H��"��%�0�snQuAKJr+��+,�*�F&�'KwB�0����LJ�]��4�����NK;4�
��|������^���N��
&���1z+�k�ڭ�Ͷ^��^�BO�����S�҉��^Sr�{���=��7��2����
�.���u��=Sf���z>�{ד�ʆ��-`��.�ɲ�ǆ��z���r�N� #��N*�%��V�O��w�O�q������
���\>�&]��^�����ɍpX�*�;��R_o���|>��W6�XUUA�tV�g#�Y�
�]#�R�.)TŔ�9iU��h.��a�F='}���^�<U�K%0�/{��y���;����;�R'�R	��	CZ���	�*c6���~��_�^��_Аk2�s>�oφ���&���̱��;�}ڡvvϟŐ@�G�����{)N�
|U�H�O�-hT�^p�f2*��t���Y�]z�P�}��)iʭ�8���*J��{����[�vBS[��1�K�n�%��P?�U!��Pv*Ya��o3q=[�sUqJ�(�x�JS�g��첱4� �5P�n��n2a� ����j-O�ﶋ�T
�)6U�n�Nǜ@'��-�^��e@�Y�暖6U�n�J�]^w�Ini6d0~���/�Y���W�&m����8a!�7u�\���G}�gKw/{���{��g�ŷ%�.%����Tw>� ��|� Q Y 7d�&�%�wj��wX�v���X.j
���j����a���RuwH�����k߾���g�UP ?���K��N��l�Q4�eߍ�����#��~���h�̇�ݛ�w���{�����&_&sfxu���+��~�t~���'��*�y�gs��+-(Kt���,�H��vi�k����]�׬��0[��F(��|���Ԧ)M���B|Jԩ;���ʔ���g�8b�$oo��Yw���7s����TD@�Xv�V鈗g�@'U��[2c#r�$6F{=���Y���d�Qu�9�12N�^wB�e犿g���{��v���k��w��߽��3L9n�{oO?���g�}����]������=�`�2o_^?�f]�[�܈l�4%Y_t
�,�ƪ�y�$�0j-�4cNA�}��Q����i��0���o�.�;=���P<�o�}~��y��߭�����=v`�G]��V��i�oV��\��c,��	C�ڝ�H���>�[H�I��1��z2?L�P?[���9ͻ�czH�u�qG>�n���xl�vf��N�+����;ҟ3q-��4^J���uNp�R���4��N��%,v�O�{����~��x�N:���"y��ZBi��76�N�'}<||@>#���l����;�W��J���N�
�r�|>�
�v�������wط�_f g���oF������>}��bU4�5�j�N��������Ĺ+�a����׵�*	*�ESm_����V��P�A��v�M��F/bP����۰����(6ʿ�2�W�n&ѽ�Gs �A��2�WN�KhAL�sr�ӫ �)k���.�NI{��j��RN�S��]mэ����,���ō�x��l v��IK����[T6yd��l�Fq�ݖ�{�CIڛ�gW�kK�Y��5�7=O|��3}�&�f��f��=�v�bR|�m��(�+_V�ewǺ��<��3X�lk���0^
36̛�m�%�5!��.�ך�ʠ��Q��h3�	��v���r;l.DT����S����^X�sݥ:���-<�C�s?ށ�B��2&����Ɏ������c�r�p"����d���
���V���Q����c�	5��ڪ�=�v�Ww�ܶ�kp��'*P�����|/v�*�`������|||@2�5�J���5��=��9��<�e�ʴ�7&b�ƈ�[M��d�I�DF,k@CC]m@*=B���c�jo8oؿ	8pn���0��d�x��D�N��$Ϯ���g@����.��Oꊤk�>gz����b��j�\�V��Ͳ��Qk��P1����5�" B�JZMJv8�j��/L���Ғ�'QWJv)�!���	o��՗�NE�V�T�%���)�^����Go�N~��kՇ�`��3�{�폇/���s�w���4)����'n��k����Ւ�.M[k�L��rQ*ϛm���eA"�6��f���N���Udu�yK�uy,�i�@���L?��с�ؿw�"V���z��m����M�mK$�)O�s���e��
�G����IR\4U�D�xů�d��V�Z�@6�ݐM�|�h�B�͡c�},B��%�W�]ۆ}}OZ�%Y)̓:�h��3þ|�Ȣ�M���J$y���N;������G�V��̋�����L�c� q�>@�(mY�"���lm����%պ&���X(���;f��b�{����K]Β�+G�LC}� �;W�{��-
����v'M-���-/���!�,Lmɴ�U[��ְP���ydӒ�6�;���ɯS��̟L�ظ�ʂJ��a�̯X;A���8�*3��b!G�3dn��0B��,m��䪗�M�T�F�jY�0Ѩi����dd,���bƧ̠D5��d\�V�џc �9Q����y�+c������A��3ff`��p�]�;�.ux�@$m��z7n�j� ��k�Fm2vZ��O񳼛�;��g��2Q��nq�9.��k�J��f{(�|�>��%�0h��z8�����蚕W�{�/�k�
�+�l��U�q�ݯ���3�{��x�d@.�!��Qp�1e-�!O��)`Y�l�VUB���f*��b�n+ڮ�@�g)�Q
��ZB�(-C"2a��ζ<	�ዷSf��^m�f��=>j��n!7A+�,ۘ����:�l�� iN����F�q�6�0(�v�厞3�0-���δKs��׆t��F�}7�{'�y����w�s-����;R4�h���>>�������5R�a�n�n"�_���b8�	�����s�����K#�h)�y���fظ�̽�{u�+��2��$��7�Ԭ�������[����T����6��:����k��q�85ࢠ������z_�������f�p?O�l���O�Ucz�V��wh�a>�6Y��2��L"Ej��k�&��c:�� �Q�*���l�Q:ij�S�,׈wZ�Ϙf�e6�Y�M��!f:wY>����2��6�S��4-4էK	�2�3@�i��i��O����e;��UB��x���ML^n��(�܁��/�p��!��:�>&����"O�x��7�i&|5�� lh1�nM{$6Fy�����#"S�	��������iN�/�>$�	���w�~Љ�fn��4:��S+v<<^�/���8���P棌Wx�ǒ�W{��� ���1��؎$�g$��C9K�0���y��9U�!*�(ֻr*�g�|k]�<U�Y��i��w�Ғ|��I����*��_����ë2^]�������_O�$�����9�I�c�)����pjp��׹�M�]�b�g��h�r��O9�"�ML�x�*��Я�����6����9�A�K���@�ϼ-sϙ^���yD���Ԅ0��gnbG�`�4!YJ}��F�8�`��V6]����˖�l�M�&�U��L�g*�����H�E()m1ʗ�$``ը,���6���J"�Q��2�Ub�l�-4����'n�l���TQM��4�9�0��'W0v=Z%][��]�'�$�S�EU>]��U�4ﭽ�[�	d�\ת(ʁ���S|Nh�Z�fBFƹJ�l��4�.!T�޹[�x*-�x��,���b�FȷR�'b
����D1yE^Z4d������''}�6е�"��kz���F�òŨ���@�����P�~~��V�Xo�#�GS��'�.�?.�Qf_58�����z��1��q�����������&B6�cq|���*���34%���.����D*�{�i� q#��ݖ+y���-;����o���w�����w'�6�1#`ۯY���_�=/s�Rpsǒ����UV�P�F�!Q�i"g�K�N�a�������g�}�3.e3[0��߮e���(��[�+ʲ, l��m^�?A��R\/���������w��f�����/�ӾujD�S�W��-5s�af�|=q[�������w�`�\)�P'@P2ҭ��[^9)#0SD���jFr��ao�ᘨ��bB�p����~^=���g�\�K�m��G0T��66P(�h�`�\d2�:��VhXg�k9CLfI�I�mG��ex��KY>�z�����EzK6�l�3LƮT��%������ylXJP�DUʽ�x�P�8c�����g���2����ƹ��g��纝�|�	��Tw�~o��oݜ�y�y�Xz���=��;���>W���v�IH��aJV�P��s�و�,��f�j�[L�.�����t�꡴m*	[a�Ր�g=}|�����ս�p7��9�'f�qn��N��c�4sj�w2���������{ô1ǻ�� wW�E�6��<�M	�{N��p�����6�J�� ����x������4�F�z��������
�-�Mԭ�z-����Uܔ�W�.�cS��ӳ����:`�մD�"�*N��tUk�ϻ�5�L���S䊖��4��^�zj�L>������IN�7������ڥi���h�a�����[O��9����v֦�q��r��흅�*�i"V���ە�ʀ�5"�EF����L/a�P�L�7 e�D����1<���u�Z̋��΅Zn�u��J��r�K_��Ȉ��W����iD�NH�!I�qYa+PN�3R6��9�"@�����+��6�g��\�A50_������}����޼���xOP{߹x���јS�WZ1ũ����Ɖᤜ�x��L�w�;�����w��X|;�fϙ�<����뚻�ɊZ�~|��ך�*�v�B�އ2���})�A"�$+Ay��H����>*z�BE������t��Y��uX�W��e�B"-@?nIo-~mB����iʐ�ͩ�\��%�=���6_0��\�W�� �m��z�܅�}ȱY�1�WD�+tf�G�s�6�}|���u���"k��Y����q��e<ޣnc�*�@O�qn@���Z�u�{Fw�d]�:�0��O{vS&Po��nў�/.�S���o��s�^��j.jy�ϧ���
�C����	��9Ө��5W�h8��C�uU���qN��`�1-�Z�Thv_H��.-w��`���1��]�L��w,yL=����Q+ɼ��Sf�#zb
�꩏��/���%�i�<��!��L���ym�\���oa�}�fv��h]vd�pu����E0�����L� y��x.�t� �}G�>��K�{4�L��o���6}��M�|3�\;�˾*�#1Q���kڽ\�
�5'�K�:�v)�m��oa����h�0��Ojޱt�"������ïh�aV�̋W�A�sVW1��K��N�5���M�.��O���Ҹ�?
��'��q*���;A�q^��G'�a�~�'f�";�V�n%�~�2!�*�(_��_K[�nS�7��(+�m^d����*!X���e��2/�4�ƴ%�I�d���n%�.���ue���(:@���H#��{^I"&�E���J>o��̟�/�9����f�����ly9��l�1f)�Zị�^�l|��d/�9��\�����c/g��U��n�&ك3��-t�W��8f�jw�N�	�]s�&&�ɥ�n:#��fq�JQ�ɶ����[/H�H���0֪��WZ�� ��s��z��5{=��!�@`}�Q�3�����C"��*���+.V������){;�ׯ�m�t��!�zo(�� �x�yVv:�f�KZH��ܮ�HB�ȝ.`�v���m�W���ovq=7Ε��M�y8��*/Y��x�L��-w�ĵ �p�3���Ι�%��Ӝ�ݶR�-s���j��t4��y�Ga,ocT8�xk/Kz��s�NE��R�{����o�>$�Ǯ��z�����n�BH�ev���i�r������Pt陾<�mƫ�v0]J1Cr��N�������B�*���)@�V�f�\����l^�/���<�dmv 7����˫j��2���e�`��LqgL�p��Ƕ�\k��M�����:M�|��_���W�d)��k��]�,�U�Y9�_E��C����Wk�����q<�y�5="1�X�w��:W��>�w{>�{}��<�,�?�W�uw@�q��^���>:���y�� 3�����݆�$�ܾ�ԪM\}q���cǯ�8�<x����붛v�F�QL��n�])��2Gۯ�rg��~|��ɚg�~{��I	)�9��#�${En��#���O_\x=q����x������m;v�A�I�����rM"r�}��o�(�(�
��*,�0f��_^>�}x=q�������Ǐ__]�m�o��	2o���wrH����~���Q�m�vӍ7�p��y���ׯ���%����;�ʏ�$M��L����b����(��;�w��@H{����� es�(^vF�ߏ�;JY,Q.����}/��K�[�{y�O޹,A`����c{�tO�{�#f��=�M���D�&���7��^��+�.���ަ���'�Ɏn�9�>�G��!����4���΀$	
�M���747�%��)��NnP\�F�)4����A>$���>��B�
F��{��m@r	ח��w,Vq�D�#�]S�0Y��=���EN�sKDx���8�4�CM44�����&Vwݞ�yo�J$���{�{��ؼ$������Z�t��- �N���-�>��5C�Ȗ~�Y���)uƴ�{�88a-��-������2\�׍X���·���	�-=F�[�i�L<)��mC_i-�����8���~N��TJ½�8|�������Ϫ��n�
���:~��dsM5�8��}��+��#f��nԅ�ɇ�5��ޱ��Ճ�]w�A�W���ڹ����;�4�\]��ڗ���WUO�y�y�&vh�Ÿ.�%=�8��Z��s��%h��a���cݿ���O�W�}\��|s}����I��݂P<����{f.A�^b�r�n����U}����՟R��,A���/���C�vu<d��G��@O�
aE�̄�����`)=��J~��)�G��
c�ܐq������n�ύy�{��W��	�g�~r�T�:E�.$]]ϊ#�����.���OI�ފɵ�c[#[yܲ���>��G���dX�R���C!��9돡�ۖ��E�����E�؞�{��hr� c�����O�v��D��χ��7Xe=a��J�zX�9�*���}ᓆm�=:���3��w�!� ��1Z��w���2��Ɲ�L��w���q�#;rr�bz��|{{ǵ���nz�t� %�r��Y�"��y����m.[�rv.�_�:��V<�w��Bf�����CC0]�w;�fa�!{�N�e�|^Q��c��������1�G�{�(z~�A�kG��>�q�O��TTD������q�m,�&
qJ}�O�2��Y�!h��,>�f�I���z�u�=ˠ�j�<<���<xV��`[g%"��D���/ݯa#>�z�zq��sĊ>�xK���?������m�ۉ�+�pɱ��}b���^-G�f��86����4�u&�7�|���w��9莹�1�o:��-���H~X5M�[b1�w�qv��w�q=����m�;�¶�vT���Z���yh�d��"LhA�2�L?�����u�Yy�,Ȇ�/���a��:�u��X��E�pCp��iO����^b{Y+���f�d5n���+�-��6�Ul�+Ǟn�H]��^ӎ ��Ũw^z�5���W���=�01��|�����"��;���xA/0J��D�J!Ef���!lSp����E��ί�K*�5���z�R�Ϧ��}��s�X�w�Y|�l�O�7������kN�c�g����pn��0�_)� OQ��:���%EÀtv�=%��v4�.�*O�;?~�?]����/��M�|��q���9�9���m���c�g9��o#g�{��c�;>��G�a����'l�t՟M!��ʺjA��C�X��J���8RfgQJ��uU��V\�~#�x�G���K��{h?��㫤")�\�wW��0�A�4��<;�i��:���}� 2��_߃���b�?��Q�[�����W��?_wP��\��r��h��Y����L��m�t��8huoP�5�v:"�35��g���a��n,�7p2ti������3aHij+�=����n;��=�e�;�<7��b��8tkO���� _��K��,���6q����n��xO�x]�Sx�x��~O�^7�����I�ԲI�t����3�����f�����/g5��<���T&xi�¨,�W7�SgTw:��L�����>oL8���.�|����h�q~�{#��������F:�=#�?����K�����v{n��y\�p��XA_0�� ��s�c��<< 7�-���ʄǆ2��*^�S��͞\�K�B}a��5:����v��KOe��ho;d�a�p?�^�P9�� ��}#Ns7hv��+\�%"��./�a��	=��d����0`��&1D
��P����-!���lFO�O� M�^׈�{�������{��k�t���)�-L�W��%��W� �F�Y;;���T��Q�u�	��;��&a�5�Q���#�x�L93U����B�k���W�a��ͮ��a����g)ࠇ��.%�A���N�ߵ���ޝ������B��x;�k���VNev��U�uE4�ݸ�P�_�?x������o7��C*�,�)xfo�֎��S�S�)K��h�<�^i�?�5�P'�����c�**Z���&ލ�:����_;0;`f��\��n������Z�]����(S���Ne���P߀lU$�H9�<x��?W�ʂ�H��r-e�Iո}6q���ҫ���n��bL�����`�01�b���p5�qMW_-�}�t06|�s�sr��P��E��ΨvM(Ex�s�m]���4l�z<���3i{������c�<VGNjI�mb19x������.��7�5G.�v#g1���P)ZP��վϙ���ib��D��!5��,F�����:��>��(�e�����{�/�[���anި�|\<� a��H;���˺����W���O^��
|`^���S�� c�ޮ� �V��"1p!�ٖ�ܙ�����?r�?��Ʀ ^b����]��˿�b�/����_t&�|W���P���N�M�\�W��x
��r��l�9�? ������a���g�Z���K��1� �\.ht�.zC5Lf`ԋŒz�;�n������RW�#!�����;,9uQ�iH�N���;��S�hJ_�{<4���j�/'T�������g�p����1��[�7�U���uY�BI��]��1N�)d3�|����F1���s���3^ߨw�r�ZnUY̲���>xB���m��";fg���ϵ�
��uJɊG\6��:ӆOx
NuԯG=��	����<P;�^dW�@��X�y~,R ����Dz#������g9j���3y�>���r7���o��u�r�܉���}�{Ph���Y��X�_�+���ڎ���������G�3;�8f]�+}����_p�ؽ;��;E�#c;�A�x6GlbP�j�mҺһ�>'��m�����&l���@r�~�G~k:c��P2 �
c��필J�jZ�:o=�ӿF�����a�_*�}w�=K���<�>�:��빬U�>�w]-Awח��9.��]��gxג�] ��
b��4y���z�q�����o?�|0� ݲiLm����۬R�t5w�����۴6 ���{gR�vO�Y�o|����#�����Q���mĞ��m��]���@��n����sU��+����p�=�v��O���Z5�,	b%�Ȉ�MѮ���y���Dw��	��>�	����r���Q��ѳ��{�w�a+=���/���x#A�f�M��E���9}��S{(_-�/V�z�LA���{�d�L�$ѵgm#�<1:Y���eϸ���z��f�s%�;���lx$�-����*�ǥj"�r���?yzc#������k�ϟ��hϣ�XEO�A����O`�J�H�Uܫ�gۀm��i.��h�#w��m8���W����.Cr���=�{'}�|_��	�9��WR�,`۷��j�Ν�ӽ�4&�0c���Q牋o���=<��'���
���];;�|�йB&���uڣj����� Ֆ�������avd1�aO�P���=I�%����'mk�F�^��Z;oEa��/���A��{��z��C�y4��C@��� ��P����N-��O�8i�7h#RF�w���ƞٯM�
��+��������ϋ�[��o�C �y)������b/A�+� '���vw�����"̊U�[�K>�c��ן����b���$�T�D�2���ic���g7~�;���GN�d�]�>�7��i�zp���%��Q��:���_1����'2�/�A�u�O��5>��l���qp��;��!�ޓ�?�E���~��x~
p s�׭eٵ�ݶ��"����6Rz~�`� �=��]7�k�w5�VsW���A����]�t�}��&FRc�?eQ�b{�ؓ�t^�2D�������P�ʧ�QtZ�`��m҃Nn��jC��@�׺N~��z��&;}��{8�[6bWz��<��K��Wo�\s/����Y�{�\����g=D%u� ��|=��{���}��7�<Nmo-}Ju+�>��@������^�o&�PU�j�*#��hмylD3�')�lF�s�_=�i��\s���$��|�;�b\zzx�6'�-㹲tk�gk���n&8�fnj]r�PE��sy�G}#�J����v����*.C{�~w��{
]�)��0�����W����7!����	�zPq���z^�f�h��ީ7�L�]����-�pD�������+�Zh-�4�XΞ��O!=I�3��r1�/�0�KB�7��]�P�B��+��d��K���>Xn�ht:z@Éi�W[����C{����eѫ����4Mwx�5�1�-�c������l�]}�v�a���v�H���ԣ�P�i���������K�O፧��Qz����{����F4�ͮ�k߹�7>`���h��C�
Q��]�*��`0��uzY��s��Ӽ�c��8��D��z���[�ˏ��6r%�]���߀�L�I�	�ܮaG!��G#�N�*���H>cX�Hs�8�l^�wוŷ�w�`�&=5�=/-�ʄ�|rJ�@d��ɂ�2[����X�5��iw�b���u��qQﴆ��]�TE�-�SCxe�~���Ly����s�w���}s2�U�>�l,*�h��[�VZ�a���âVc�7�wf��2���R��>�K��-�t��:��sQ�ia�]��2�c����|}���1�cLi���{��W�|���j5yȋ`+����9����S�R+��O�#<^��ҟ�1�W@	�[fpZ��;]��zU����֦����Џ1CG(�m�O��ベ�C���\Rjk2�X�ERt6wzܮ�
U��D�<W�l��<��C���`�`k����0��	�����4}�	9�'o-���݋��_v��w�I�LXix� ��; a��@���6ɼX[:}��߁��y�hކ�je�N5Y�W�v�4��f\S� ��z%)��C�D�r���ׁ+G�[��Yy��l�{y��b�oϯ8��������{���L���!
�hy��6�oCL�t�Mu��!r��h�����jA���Ao����ϕ��\��5�~b�ܥ�����y�P��ƶ�a�*�;��H���c���j�i���ƚ�9�]X�;����tM7|�w�^���w�c�cC�^r��g�%i���1� *�ZfR��<�ޡϛ�{�l��/��{�{�ܨ4v�=�t�#������{�û�j����O�{��o��]VV�J�������݁�L�����U��R�r�o=�2�J�*��� ��!�`�`�.k���ٵ���ᗷ��<����}ͣ�g�j�YȮ���,�d�yU�n;�p�\�M�w=���l�"�i~�������ա���Y<��om΍�|��Ǯ�
�O'���4�i� АEd@�Ǽ�c��Z���82nD"�Y�y7ÌSu{�W7�1e�=��=k�;b�s�n�sV�<Rg+���xE�`mY Ӓ�q1I����z��/-���uv�qx4@=���}��5�)�����{�cCp##���`6��H-�`GneszO�)2�=s��r��P�f�{Gw<�̞ʻ�c�������l�h��Y�>�����Bj��k ��U�c3w��;�:�=/��~�]�9�<��x�IC�Z9�8f�)&9�'����:�Ȃ�}������g^���J;�t�����W��u0���sܽ��U>[�}#`0`��ߝDz������י�\��Ҍ<ڻ�嫡*�4^7<�p#�^�(,����Pgc������o&�jwl˖ٔ9����_��ؽ��f�k��\�<�=-!/�YHנ�=4;a�� V����Rf�K�7(-���n��>��9mĈ���q��n'dQ�_|�����ɮX"���9����4�{{�J5��O��|!�1�GN�>����U����g����ڃ���a��f��n���Y\弽jX��1n�^�<��/5���X���Մ�x\���Q���ߟ��
������
�3���fj�o�F=��v䂗�-����Z{�]q�\��=,�f5	�s<�$�D���2˭�UI_B}4ƕ�1��1���"���2
s�：��w���p���[�\_'Ho)���A�~績u�.z��wuV������L�>ff�xO��{��@k�;�lDl^�9���;$��l�T����?�Zi[֢"�[��Rް����)�Ғj��O]�s|��@�V�o	�9 `Ѭfȵ�uN�8�/k�T�o{�o�B�7H�ce�-c��PοR�X6�(��O�EP��Xhuej��'��s��v��e�������ẞ�u�±�Q��@�^fO`�J~�.�
e]ʴٷ̟��w3x3y�x���������c_��v@�>�O���~��@�u|
#�7�����}�̆[qq��;��4�E'd�QкF@/�����μ?��t=<��[ʵt��];.�# qf��l_u��)�yew����W��������nƔ��K
�PKE��{��@�.&nׯI��>�b�ݡO�ɎZ;�#��е�\�_{�Ā��E��l�/q�9z���Nw�]�+���V��m�P�!����`/v
q��z��#�T������FO��g�vIh*�~W���y�n���yӆ�}7ݷר��j�-[�`ۺ��\��۞���fv�����ز��6��gr���,c�M���1��uu�`��Rou|n��=���޾��P�V��fo���ͽ�9�뺏?�=�x������'3�V�r��#�>�ȳ&M��WQ�޹w��`[��'�DS������2@1gkX�O�v�*û�ݹLYn�3ؽ���W���i�-wU)��7'����^{���p��SԸ[6y�r��3	[�AT�t�M#�z��{\OK쫩����3�vK��-�]rf�d?w��*��X���`ʵ����hҳ�2��x��LE���#!�H�/uw�v�;;�\�	U�.�p���7vww�;�����}<�-��!��}'���7�ȁ[|�}�l8�^
A��\�����|^DM2�����O#�w�-e���;�=ǹYvx���9 ���	��ѽ��?C%�����:�{�P��J�͢1��*����W�"֞���L����TJRO�w��1����.�.w���&!�bT0�t
6V
��ޝ{��?~ύg8+��~�<�A�����I�ϙ���/�M�wM&O��4�W����A�/�t���U{9N��pAv7Ưb9F������b�����u�:J����<�ؼ����B�������ݸ��\db��ܫ�����&ь��F�a'В�(G�96��&��/��x[7/�p[��}���]
�l�v�������������y���%ݻW^������mJe��׳��[��h�WOq�ا�/3$����y��ېǺ�nrM��4!,���>T̙X��X.�8VLyckFT\�A�Z�^��o{���j����ܦ����X^��x8�w#s�n��L�Ü��=ԖV��n�TS�H;�7�s٩����7Q��õ�^��k5q>׵U�nZ���t*UR�<
f��qgb�n��N�-�{���W(Ξ��V�΀�Q�|�+�sM�\�5タ��|fq�/L���-�k�#<��=���3�̠��
�˞H���mHqnf;��
�R�{�u:�ZtT�;f_\LzS��v�'Emә��2�U��R�����?\U��;0^�����v�ĜP3��h�f�>Y�C.����<͓$��w�v M��5�& ��xh������e7�3f�٨�L~G�>==!��G��-z���,Rɾ�˓4痧w_ �W�X�������ʊ�6��{w�.�D���!N�uʮat]o��SǽHi��	��wS�^X�˹��ɾ��8�ؓ\�;����{m��e�y^�d�Q��9Y�a�t�������?{���@�Y���H���+��do��А(��󢣕���Ϧ���7w�����׭8�}}}}}z���_]���{�����JF�W=݌#�w�������O]�CI��>��@_OV�^�z������������ǯ��ݾ�{���Ͼ<�	����(H�D�������Ώn�4�.�w>����x�\q������z���۽��o�����Ji�rI�����K]�1�X�X;�(��N�FNWiZO��.�I6��邌�A�Q�"�nE��ﮘ!u0�`�K���M��$��\"��B�C?���k���]t�YdK�͓H�}u�DQ�܌)w���z1����2��PspH����L�cg�WǱ$�E�/ͻ����4�d�!At�#�n��o/OA�6M��Q�( ���ś��ڹI#�$��	�ſ��$$�A#�3<N$�1�ZӦh��6���b
�BR�^!�4SA��`���9
�BD��cc}d*�s��گ���3�wguZ����Z�s
ff{-��Ѯ�l[�.Vg1}
����,X2F�.�z�j%�_(�%�I�Ï�Č�I��f�E\p��k�l�\1ƛ$n8
��0' 1�$�*���m�1>%��pC��FR_
��eS��$���>;c@��4�cJAE�o�
���Mo���c�����ѹe~�����e�ͣ%�=� �o�;���PT��r�S[�Y�~�/̈�/ݮ��I
gX	�}���wmÄ�VUo��3��l߀�F�_Ai�4��d�mO�I��plM�4��	�In��i�}��9EMޘ�k�km��,��V+���������G�)z�� a7ud�ǀr�xP&%9)V��:�"Dkf_Ci^q�<�ˠ`�����_���E=3P[�}�ѣ��dy��kf��2����3Ў�� ���@�¸�XW��e�'��J~/UuKO�`����6%���&�l��nU\+i�]����s��*�ѯ-²��^���\���>#'ƭ�8����$ŏ1ѳW�IJI;�L��4�� 6S�=7�S
��h\�ߧ�݄޸�;�c=( �1P�Vӂ���;�s��� �7��d��_�H���{d�o���S߰�	�_*��XK+n�gXl��eDg#�Zmx2����V{�߻o�Yº�X�=�:q�b��3�w��ެ�V�ҽ]��{�^��˼�@Nc�Sǲm�mD��S��{o@���<���~�(8o��h�+?b�d
���显h9"(d��Ʋ#.&\f9�f�Po�f���ݽ�q���_v'd�WZn����T ӧ� ��r�OS)��/dO�wD�]��{��,NCл����no{-1wu��\���S���߆�].��k�U��y��� SCBM((5��|����~|Czӹ�>O˭����P\UxP{�/A�����z<�ƴ��m�z3�4��s�ވ�|�g6;��!����ZNO��>�
nokp.9�iy^FO��
w�3��u�G�kZO	$�n;|K�1��pt�H�9<��+ԋ�b�#��(L�*��3���{p)rY/�}]ƣ�f��|�cJ�<4_�Z�j���iu&��%�龺��k>����ץ��giW{y� 4D*³�BHk~%��C�jEuxĔ�7s|�����C횔�k��:��Ke�F�S [p
�ĸ#+�}>K о��\Ծ�Nܩ���^���b��G�W|��vzl�a��6$�,6˭�@h����}͡�7�x��� %py��C��/gѐ�q_K&lR� ���	X��xѢ���tX�����ð<���hN���P������>����\N�Z��������[��qM3$qp8A��.���c�p"�W�z|�L���g%w�J�Ä ��ۢ��O-L6�E��1�vH�ޣ�|��޸v��e���fr���1 ����m�{�7���cu�ѹ����;�ɼ��~�W�����Ǩ�� ��O $|I�H�)�YB0�!���������Rb���2A��7|ᾒjKLrу)�8&��g�.�R�������>�G���
SC@M -A�DFEY
��%�~d��,p�r�����tO��[�_�%c�~�g¤Sgto�� ��eV������8)��7]��@�E8sqm�޹��U�:+Bjƿ h>�5Yw�·����Ĝ���/[�y��፨ �/@?� ���bOQ(��(�����3i��6MM��;����wk(F�yC��y�}3�s�oޚ~k��m�a�f*�qYZ��\�e��,�(��@����M�̍'"��3����kv\oH���֗%�{�ozP��L��;�s
b�.}m����F��:kgol���a�>�A����>�K�'�T�~���+
��oc&�O�Ȟ���P\�O����BP�0�= r�_���Բ�JΓ� _�F]�gt#y9�3D��?�w�k���n5@�!��.o���t����Eym��8ӹʅ�K�K����P�]3���5{�z��y7v�<�n1�����f��_��@v�}(�bA�B�><7Ŷno�����H8�,9#<\]	=��8��c&�F��?���]������w}e��*��M�7r���9u�nߒ�{��'������7���]�<td�:z)�NP�+]s�O ��w�<H�@��`�U�!�x�o8ඍm��o�؛��okjUp�[���]TW�x�r�9V*�C�5�������*�44���Ҫ�s�����/�dSu�^E�y�ʐ������y?��|������@��A16�?6�7ޫ���7���4��*��5�\�}�^��� �x���� ����RS�m4݄7aI�W[� �{�	&o��߈���5m�އ�t�BW搊�h��m=����/&'�#���7������Mv�\)����F(l5��Q�-O���1V7]��>�.��U�)4�9���.��Ѣ�q!>�;�i���
b���5n�x��˫*+��l*��h�z��ܔ;�pcK�Ú�~�`S>�M>�l~�5�s��P���r���o#;B��M"�z��ڻѓ%ʦ(�+z~�����tM7�=Mj�%�l9�zޭ�=[��Ýy���An�Z�fnʘ���Ë�<����|���=`i�e��D�)�@[0���:��^��м�[��Y{㷶���`O��K��1X�����Z}����.�,�ʹ����p���-f#���;�b�џG�H�����c��7[�xv\����ej�M>���>�mڔS�Ʒ���;��!����%
_�}�f�~�피�SחV�9�K^tC���I �b�vk�7�%9��6/%��'č��2z)�1j��0�-kF�6V��o�4Aݶ�f��1���|�Vt��g[�y��rj��w��%y�jI�=~���UhhTB���QE>{����Z�5:6K�]��m���N���~�6�q�1��'%����� �����YZ�2OI��<��o��:���y����̩];K��4:�̬�v��� �/�����f��^Fב�~��]��а��èB;>��yc[6탹����^�-�F���	�{&�I��|4�]�n�yW�%�~M,6Q�W/l�3y�>^��9� B���p���WL�N?T��ll��as��a��W�>��㴃�6��$�%v���/}��:��гh��*p�AV��#g�O=?�g�|�6�N;Ē|G��/!^���4�>Z�nW���y��+��=>1�;射�̿I���M�2���	;v!��uڛ���ҹ;�������A!�}�=(��/��]hx����&�V>�������b}�����w��4Ws�Aze��~�MQ�^�}��|Vb=�|���{�"��=��B��as��81�4sˆ�W�R��}�	���셜C�Oa�B=R�j��Y>{/Ց�TSE<���d˪n��S��{6�͌ގ��.�k����:�)��y_��,�pUa�2;pk漐e���/;.p�iIZ3�O*�ܾ�jUgr�,t�j�l�5�H4���|�������?pzL�ۺv5�=�`R�Sv��x����e�+,��ú�h������'�x��Q9���!\ߛ�H���iTi�� )��@S����&�{ϔg����z�Wj����\��4o�c��!�{@�5��͸�h1���ި�p����Jζ��`�0k,>}]b�N)�Ιk�������[ss}Yd�;*��\�\~�U]�%"ޢ�=�Κ߮dUk
������+#�@O��^d�߫ON���o�,�q*�/5n�zr7��(yk��\|�G1U}_:��~r�u�v����Ъ>}n.�z���wz�	-\8J���x	����4'��k��,[�|w�[(z����߲�~?��½���b��`��޹�?q��RZF�I�)��t�����W�+������;�29;��ڧ����:�9�7'��,�@��9\¨���j���)���=~YL9���I��)4S���
i��˳	�̑劣��<�B)�hN��������L/�R��X]Y�ZTd��O۴�������@����!p��^�Ќaٵ"��bJp�����7
V����r���I�:�z	�S�E�|�"'����(��'��G�|~U}��A+1V�J�[4[��x��M'��-�wq�6,�����t�.*[�+��]T"�F�ܣ��a�k5g��D��-�'�9�����{�F]�!�����FH��.
�<���gw��#S�?Y;�7����ے�؏�Ҏ�������J��&X�@|~���@hh@V���	��ΞU�K����
L�m��.�;^J�i[4��ζ5hP�G0��N{�WΠ�ez¨y7};Ѥ���;�x��s���kג�DS"�����<���\=��T��r�ozF�$]�#~u�ג�
�������~A�P�-�k�<1��do'mU�F������0W��Ё�}�jZ����9Q�_���5�l�]�S"��Õd\k�7u/�x�P�,?�`�$=��<��s�"�v{�cX�C/u�jƥ�=���̖��gѪ���:�-��͜a ���W��ۢ��b˱��|�}Zl��#�����U?\V���[����#P������/���R�LѲ��*<�!�����ʗ��5�l�9ɮD�ߠ;�xb��u�[`n��o��Er]r�+�~z>|����*z�;�a�VQ�@����M�}!
�����xe��������v�E.����իq)c'�N��.�����2�G0֘rϸ��I䘤���T�~�s0�@v�1��-��_�����ez����5Osە<?�����~��7�w���������G���� �j��͗���t��@|r@xPWv�ae��Q̛SG�Wk�v��4'n�u�<��-�z]�y���z�u�\ʊ.�� �}����UhiTi��*
ܭ���s�^Y�5��ހhC�Ѱ�|�&`���.���,���2�S��r�wy�(�w[��4b�=��&W���tj��0�w�|�>s�l	�a�#s��X�cbf��d6�@5*�*�G~J9�+˨��hON�����G_�?��.��m����
�jq���m]�i0����t$�/c�<!UH��drq��P��w�=iN3.�T</t�.��OL��i��S*�46����>�z	AinD�j�u�4D��3�-Mw�������~�w�
GNjd�_-�m��O�����H�r��@: 
bǗT�p�5w�{G�}��tRi`="�.u�ͧ�/��9!�0�0���I�1sA����Ʈ��+'y���u�T:��d�0΋](���������r��"��\��]��cT�	Aw�I�R�3)����O���Y�r�u�yV��ü=2$6um��^�����;�%Cva�i��r��;����+g`����~ˀ�+�qv�%)�C��kGicb�1�a���s�!��p9|����Oض��s��5��?�]�ٚ��w_߫�v�*�0V��#ʰ���t��4���k�����Ƭ=�n=Ϗ)��sZ�'iBU�9�Uݴښ�"�Z�Ar޻g�!��hQ��@Jhh���{�����5sY�vs��F�Y;ز��n�lHd��C����q�tX�d}ږ@���QÖ�KXe�mS�wx��`z���(By�Tpnd/�y��[xhF3�i�>[�t�&{{7N.�i
�z48E����q�@-�8�:��w��~�ܧ�_����%�f�s�6^�5��*��u& ��z�P����c�SX��̓鈔��Yh�:ږ�gT&"������|[Y��v�\?O�ϞG@Ƙ���O��v�z���]mn���/�i��m�Ih,;Ox7H�Au&�(��a�����Ѡ/�x=<�#�<����+�Q�3�����٦c�v�M��;���ct�o*���!�K���C>	���!b��s \Tk���9�G�3�=��},���1,�ٝB���V����1q�K׹��G�ü{ {m�;`Wl����Nh���m�'ܓ�9nU2%/CC�m����Lw<y�a��@_\�j`e�[�m��Vy㾗ɝ�*�%���Q�x�'�'��Am��w�}aD�L�ݏ�/*����u��;B��,<+��L�v��AC��x��h��|�莬�_��9�uߗe���uR��?�#n��y�}Dw�͎��{�r'�����显
Q'+��l�a�3i�g�d|kw�����w3��;���|���<��?s�]U5w�T5���T)��ho,����]�[N��ee��hն�L�����T��*44��C@��_��n����=~wQi	�&�'��1��`}(��Xi��և��F@q.ƻ�Z��͊�����/��3&�����_W���$�����`q�W75���vu��Y��݇[U��c�wF�P;%*�4��Fypުꖟ���y�o�`~��J��3��.;Xpy�ٯsq���C�3�N��	�4��_%���ej�׼]�F5Q>Ó���%��a�u#v�>A���e�u��^]�ı����6Ҡȋ�;{m�t<��Tt��7�'�1�.�9�F�T���3c�eOxa2�U���+/M<:g1�XS-2f�wDڲ(�w&�;j���x����7�{�����<����A{v�U�[n��8����DO9�^��+�]��"c���0��Z�s�(E�g�tZ��k_j7��˔b�]7���ԙax	�����.*�1Eٮ�d�����F�Ξ���iۄ�Y���Z� h/=~�H`UZ��f9	E7'����v����s��HY��=��>ٿO�T�'���m���ky�nt��x����q�Ӥ�ư-U�ʎ��)
��g^s���	�t����o��������)wC���yw��Z�/��Zi;l�INf�i� �U]mg�F&A7��Ph8Yh"�|����娌�<w1�q}���}A���1a�+�y��n_8y0��m�n棓3��MkU>���	 ~�4p@^����:�U��1�.�򸌒�'8J������=�z]Ȝ: &W��hgr%:Ue)8�wӖR4�Qaα}����{�άs��_�puǁ<�h@��	z[��_k<K�1���Gk]!	���}Po�IuhŜ;'.3���Ӽ.v��8L��Pe5�bz۱�1{��+y�~����w��l�Q����p_ ��R��F��+u�G_;)�UD�bñ�-~R9�y�<#>��w�������P�kE|Q�,�w�6���o)�Q
nv8�[�J�r^�p9�j۝�8����nJ`�i�$ �%[b��}W�q��h��t�DS��۬��V���p�+	��i�*|�T���x�1��C"�T�x}ajw��+Y��ןd������;j�{3/wdBx�W��q��p)�����z��a=am�,@����;{�%d���)����������T��EL�Æ����y:��keG��M�s_Xc2�g�mK�7YYR�z^f2�-�˃^�G+;�����+۽������o}$���q�]�uo�V5�����`�_
N�L���UL�r�C��\/Q<x�t�nG�6.��L���8l�n�S�������Jr�wZ���\-��¶��٫ٗ�Y�J}��S�K4���Ϊ�޺�m�7=S=���_��=��f���C�
�9Ĳ#�Y�GcҼ/��h�V��0sْ��l�1Ľ����D����(M�^b����)�S����7G�l���[h�*��I�9���0^���3<�M�N�g�k�Lo'b�գǾ��.s�i-��d�{�u������!J7��\���}�͌�ے�H	�|0�B]q�<��L��l�S,.y�ۜ�PF��Ƨ��\�I\yn� ��P���!����c�Y}���d�&d{�����(>Ñqlj�r�S5o��:���
��Cb�t.Xޏ�Ruq�Υ�0Z��Ver�}-��8���DJ#�ם<�S��{���[��)S��s�xM_
'׺[���A��ϧ��e��H�l��/������_�/�ӹ�Z}/�����^���>}���;�7ک��S��]}�����=�G1+}�������;'s�;ͳ�=牬�s_���T7�U��"/Po���$e5:�\
"24��뷮�<}i��q��z�����������_]ݳE$*��h��]Q�-���E���D�O����v�Ɯq�q���|}}v��V�	 H�ۢb�Rhьi�6��d�j��=�Kz����oi�q�����o��ݻm�$L~.��u��QS6J0k��F�+t��6�$o�w�u%��DV<��d����Q�����r*I	b���3�r����'��_j�I��W^�W�6|�1�@I!�$�F�Hd�`ť}uʊ����
B"�`��L��Ɍi
2o��� ��m�MI��@"[��?]n\)����E$k�p��,QF��L&�`�	%��ۛh�F���#&CE"b�����_�{�|k��'�ӻ8�M�<){1�ڟ���B�A}�ʥ[hO���!R���a^N��y�y/�����4(�CH!M
��!��|���ϟ3Z仒�naik��&��s�D��	�J/1���wBe�L0cX5I5�M��b�q�O��C���@���О=�Y�`Н��]������r��5��>�-X��nY���Vo�T�K�`иgh��a=c2��`��������>J�2�sc�S
��%�p)�z	F�Z�� �`C���,����f�V�ki��7:��K��؈󷞽Ʉ��Cm9���YP+R���lҞ�:���Bap-#ey��[z�yN���}�w���؞����S��TRP̱�+,����{i�p-�<�k˺��Z/����t���}��mF��"��g���� ��v�>ݑ����IH	vZ����]�wp�}Wꉞ��ϒ|d�1O�	oy�^�魩���6��P�j�;�#|m5��'o����6b��k�<X���n����D`����3v>�`l�wh���XiҼ�G�1��Cit�p��de�Mz���CcW���}Pj�����B�0�����crރt^��DV�1�L��fE���}x�vg��U��7���2g�_��o0�p���8yr�C}`ME�����uJ�ƺ�2՘���\�Dov=�r��e�4r2`ih���f$��/�[,�Н.�������V�>�.߰РSCJ�ǟ�{����ل�}����)��2u^�
�M�P���fRf(ޏ; ��K]�T�s�~W�`�JxUTy�Ux�4�D���\����i�{�k��g���S���Rɉ��*T	���fv0�E��:8|o��F0��g�4J��<��-�wι�<�w%0mz���uT�K3/�K�6��Ku?���zFxo�쎷M�^|�1i����)��7F�gC� �-�����NN�
���,��w����$��"V]���:y���d����uNK�ݦii�w{۫΅}��������W�{n���,w�.B��7�P3K4!- C�>P����U�Ѱ�CF��+;�IH�.h��V�B���݈���q��<� q����;w��Y�N&�nj$k�F��k�D�O�w��	\�{��I�^�Ȑԋ��a��3�X.��ޥ[X�����ֆ��I嫣�B7�<�@����S�^�PZQ�^�;:�5�Su�93�K��� =��6֜�����7��˝+�z9��N�������4��M�%s��|�f�h�c83��x�L��\�%�󞌼�x��
�������Z�OuZ	/j�:�T��E$��قLn���VN��B�k)������a�.����ԗzt�8��z�J-�  ���{�i��V��ߚ��y/��{�%yw��^W��7''.�E|EV'$z�����h�2�E�4�B�8H{�ך��U�}���m�5l!��]�/�Z�8�^��1��cGt{g>Kǂ��J5��+�ad
�F>�ӼL�Sِ?�9'_b��5B�#5��2_cx�;E⧘OuHB���}��s��W���eW�V�X�6	��1�o/8�E>��k)���f����m �T+�dhn��8Ú�ܶ��O��U�J���)'ao�zl-��%e�L��qU�-�0�ѱ�[����|0f�Ϲ�i�y�:}z���Eu�*�o�ݮO5�bT�����֚�:����Ɂ�.69�����>��_g\>��\���yP��nhr�;1��D��e��VtZ��Q���:ƕ�.�G�
�>�"�tM�'�����ypu�墸��l�ϔ2�-k5i���'��]�sp�C��?�(��'��7MF��r^���|��sUg,-�3��r�W1�J�Q`Y'��o�8�8ty�?6ؘ!��Np��;���v����"�ނ�r9�������^ ��	&
C�O�����/S�_��D��4v�N����v������0]�|�m+2�a7�ɒ*Zѹ���[v1�����^a�%����$���"!z͓a�V�����;�:���[G�D]ކp�l"c��,�����:"�/z��_e����C��h���
hiU
�{�r��No.c�`\}������T*�.�3k���T�e�}lwo2d���G�_��U	����Ǿ�G��!gQ�[�k�,>-h3�NWy��웮;z�pUR0�>�/��\;NT��<s�@�O�/���(��u"W����ԽfEu2♆�}n�Ԍ���@��uxy�6⫤������o��� -��ϊP}4g�uC�u�/-��sc7zR�|�w�Zg
̎����EQi�������Xhg)����k����B��m�[}�zճ6:���[��Q�)*�^����]�P[����^x_��D��`p[�������g��Θn�wik/�2<��en䀘�8��{�՟uKO�b%c��6��L��b�ѷ���%!�=ű�MǢ��->�	8�/s�C&��8���4��z�{ܶK1�t�Wzs{w��_�(։����F�B!��,��~6k��<���0�Û�^�T���w�����3h���B�Ѧ�|a��Ѭ\�琟�T�gM�6��Zﶵ��}��O`��
��Y��h��3e�������:ж�8����B/M��EvJƧ�U]d��t�&�	���B8�j&^Ɨ��j���y�t��vM�u�c�oHfv��p�$泷��T��4�SC@4<����;Y��o;����ޞ�b�t��{�����4ՊVS�?5��s��\�������?��o�q��:Z۔Bd];�~>��Qҹ��l�	�l��0��CV�F.�)�Wf~�͛5����M��8��k�Ix	��6H�[=.)X�Qiٲ�^�'J��2glER���T:��Tn ���5v}]�3�P��*)�?g����^F�3E��-L�Q��&��o��{�n*��&�d?r��5h?�F�w�z	�;g���ə�M��Йwqm�r�{xU���&��K�5��FǏ:�E<���~&w'|�߽��+p��:y�cnV���
�7�����g�U$�	^%��	���n��v�SmBez"���_�����q���Γ�)�,��-M$�`�"<��._�Dg �{5Hl���j]:���Q��W3E�k�4�y[@�Nf�����-��S�gS��hP��,�m9
h}�ʛZ�q`���zw����@c�d�I�̓�>�Sy��^�T�啘Οemr�ɫ����s�U^K�Q���;�,�z��2K-�˛�DU�n�긎�':wi�3 �l���q�knцaׂ@�H���T��?<nx�q��s%]!����R�V�m]	�;_�
�{�dJ���Zd�oU�5Ysr\����{�����)���|�U����������-�55Y�|�{�8���x�9�ylX<�"�^�¨c�4_ut��ma�v$��f0x����P��:�{N2-��N}1+61Y�^�p���:;[�����k��7�q\�xךנۓ�G�O���Ҍ����������H�Y��̹�}�X9\5�(����IA�y�\�C���3����?�!ug��frơꕘ���w{@������j�n�|���~�hR1��-U�e+3榏:<�*s����y�N܍M�.�8ވ�z���ͼ#[=�'��ݞ#J�O��X��+R�x�%{�`���D�~&u�߶��8�'%�q���B����Gk��Ys�yn>ʹ�s6�w��Me��[��.89�����"#�c=��2���'%�?0�����Z��E6�g\m�q^�1�ݫ�r^���=M*/G_�t=<hi�_`���rqv�b�p9�v��g���Ǥ���.�ˌ(r���X��1�����|0���T��9<6z�L�[�?"�O����r:�;~�{m�˓_�1�)���:d�L�E�Vk�Uy��_K�O/n�0me��^�79�N��;b����u���͂3[�s���z���y�&�^Κ�]|h~:r���^nI�+��4+M�Ъ(���K�=^a�����;��d�̪ҁ�r�A��[�En�d~�$�f�B���t/�Z��}ּ؞�l����r�����?������sӯ�~��Ķu	�,�gh��T�{�'�{p�T_�0.���5��M^����d=��F�г'V�����;O�Ch�����^�z�PZ|�Ȋ���NOsk'}��si�WXO��ۮ�O�.yX��-�m���>��O��`c�{�;����1b����K�T3D?6�����#�y �~@#��P����+aݠ�������R���ŵU����7<����뭄�,��ct�]���A��C��z��zI��6�i��qc�K����T�5Az�������S)��"t���O�������O²nC���A3@�]���S�ў��<�]�����ݾF�ޙ�z��ҤS�W�Z�Z�j�Fۯp��-���"��>��x\���^B��Tpnjׄ�;��
F3vR]H[T�Y篟}10���0k>���Аw�x��~��LP�K�O��Q-ӌ/����Sb�5�os��{�1:=��輕�?7��(2�ƨ1X�a���۪pt�3<�;���B��ۙ��Y\�!��>��Ő�.V�M�y�A{�mm�s;_w^KJw@��c�܎9�����w5��3��(��B�C@�п���ofl(���
/v��{g禷{1�y��X�/bԴ���Q���wMU5[S������S��\��$w5�_p1�,ǻk��F�o����Y��liˉhAn��g֜t���w>x�̸�[0�P�����G�ƍ`�_����Ã�!'%�{��c-r��=��+��X릹r�����!4�O#k�i�.�[
RScKw6@R���ގ���ρ8�S�^1z%��ۡTO��#���t�9��%<�A�R�6>ʆ~?����s�=���z�ܟ2c��L�I~�0%���&��2����z���gh-����E��n�魹�i>sC��C|�+B��ΤN�����}jEqw�4�kqx�/aTG\��̵(ޯ�L�y�w��y�F�;�t'�O�BD�~^ ؋�uTGA|�.��!�KY�=\K{�8\���Wp���~<~9�	
;��07¡F�i#�G��U��=�P�vnr�sF��*����/�R1)�%ɥ(f�{�������!�,��+zs/�*�-�k�s���;;V�ex�u�#�4�S�}k��ws��,o�n{D�JP/�N��������8���^��j����+v��6�����<,f�E=����M�V��5-�%};\g'�:�|����q�4)M SCJ������{�˒4�O��-Pj������zs���.�><��6�s�/6�jv����F�g3�8���"�O0���|bm�.*��{
�W�`�M^]s���!���0ɒ�ތ�FX��gK��x��%x1��_�W�]�$S�=�to��4�͍`�!��ւ&[��c�|5��¨k�!mF�|`����\�球Ї<�j�fZ�>UgD�Gۉ�/zU�o�'	�p9����v�mͮ�F��ra�Ӷ�++B��W����jNBo�$n�6�A�;c�Y����9�#!tt�qv���V�V^����EQ�/>���Y'�v��e����$Ҿn '�̺�Ȯz��S����.�Xv��#EK�n���q��n7C�l�5�Ctђ��I粢��ޖ S�$wKP��8�sf��U���j��Ef���% S�6�~H&�/�0��#��}T"��ԉ4r���O'�C:�9�U�Wr�R��":VA�Vy2�0�C	
�34�S
���w�[KL(&V�$�{��`s�$���m�O<�r���d�։ה��6~v��.q�\��ֹ��VLn���=�檊��|J�׫S�o�� ZC��l���������]~k�Dz�̊�s�:��z����`�*Օ^o^����;��q9�]���H������.kW	>�O�Д��4��"s������T�q�&d��Z�B{mi/N���}H;��~7�ᬄ1ùg����1X;��%s���{��9�F�Z�{b\0�#�����h�I�Cju���P.��DH���'��}q���*�qua=�����U�\&�.�Xh�2��o�př�U�e�8?#XBomm�����D��?��E��yW����P#�DS%^cj�}�\$�����%���hг�?��d[�g|w���x�ݐ��Q��M&ô	���1)�gzJ#o;}�/Q�G~�&}�h�hw��ՑU�4-Yb�uÛb�-ֲ�
9�t`�oV����W#$k�7n���W�)��:��B���/"aA��g��&��^�%�\��hnTdo��2e^��P��Fl�	��M˭yg�-�s��dI�+��.MDl�OL����>4��;Jk�R9���P�x�r4#����G̐�M�tw��3���N>��k�Cz�6i���xL��5m���4��m��3���d�\������y3�ا�j�����,k�̓\*R�h��j�o�F.�mq������xKF_t��s%{%jnɻ���%`��&�Ol4Xĕ��Jܹ�*U0 ��cc�Y�a� N�uw��|hZ��eǻ���%ܪX��j��.<s���~���Eչ��l�|^��.��K}�b��]������Ѝ
5���>�j�0&�ͥ�l��>��z�^k ��0'V�y��ާ���>�Ut(}���|���Sl_ͩ.㮱�c&Jw��q�jp���'>;2݇����o�u�]f
�-7d�q��A�ԠԘ��iɫ�-	Ew�軼{��*[W�T�dո�%��Q�*�������`������U#+r$:�˱�)�|����Dя2Q໴�;����;3��Y��y�/�'�UC���vyj�z�
Vx��oO�����1�rn��W�2��β����c4\�/X��
��m��.��Qws�eW�&_q�{��8,��	�����s�;�YGn��z��[Э�5��0k>>(� g�[g����
s���	����k��_�[�˻|�u�by��AL�����[��w����N>|�i���=&�t�R���r��86a�7�ewW`�s:�#�R'V��U�5�u28�tҎꠣ�_Nh:6b�;!��;re��4B�C)KQ(�/oE5�"�;�j��Z"�@�Z��H'���
�Α����#\�s���Zk���#��ץr�X�!]�mƜe��7�&�s�wJ��Pex������Q���n��U�׎k�]��#lq����Ј7EX9w
��N�M��}"����@�l��Ry��o��阣��0^��iۭ�j�e�;8�T��L뙗�7�+���r�l��%�W���{϶���յ��}i�v�ȫ ����=:��=��׀1{'4L�I&��n:P�VfiRl������wiK;��>���,ɥ�9��'����B���^M���Q�A:ެ�%:���G�{�^�g�d'8��&�4�r�X�U͉L;���{G�[L�=��=�e;q7㮈3���>]<u�Oozə�x{ tO�����n����{+���(y�ø���>�sO��B�%��6!���el4
s4�4��c�A�ۻ��!a���U��.,��7}�C
��K�W�O���^V&�|���:u�,y�\2o�<��zR���#�	P϶b�>�F��`fs۽�F�{����k��Iw$6�����y�i�1mg��;�yܝqI����C��0gA�]���ܮ��Q���y�W��ϟ���;����tIb�6IO��T�X�H��>ۑ#1`�W-������ߛ��Ǯ6�8��������۶��FJ*��e�ܓ1fJѷ�e]��������oǎ8ێ8�_\q�o��ݻm.3u�J$����w$i�i��4�(���7�
�@�$vۧn�_<q��q�z��[}}v��E�P�I&KF�F�(��E$Q���a������wӘ�0�ע����Jꛐ���]F��,�Tj0b�Q0�I21H���e�"J&m&
5�~��ow	��"W��}+����1�50M�r
�LZ(���*+!b�`�����cd����`fbh��(�TY"��$���͢�}5�����{ܛ? H4!BA%�!H�q8 )����e>EBK��"H���4J*�7���ť�a� �F؊D�~;��{�d�R�B����M)�k]��t[��C�Ļ��Is	��HX�a�������H�_�E�n&�n/�/�p��dDD�6l�Q�P��$6mB�i�a��A��&2������.D܉8�d Ad�\��ѷ"���~44�ҁ�|��vy�5�/��~n��结WJP`�e����\/	�6�k�V�/��������q��+�*��N���s���ݾ�H�b���A���e�M�`��n9�ٕ2�|�$t�7Da�5�}�ci{˜S�H�	�⪠�{j�le���݄z)�� �r�<�"hϴk0��Wэ<��'����ʹ���ٽ=)Ɠ
_�sz/����*��k����\��ߎ�5��DGՕDE�#_3{�]3�뇾	�;w��}c3WWKм�n��	z�dɥ�W���ot��$?]9ׁ�6�^^��p�:�1 15�-�%�zx��I�_��#�f1�]X<(|���EUp ��lP;��GWLh��+��������iH�5k�s��T{fĭ`<�72o8��2�7�T
 ^_�#��4=��ӟBsɿ����&���s���_u\}�u��{�X{b��w����������/|���.�G��a���\�P���'���(�6��o�v���4N�������H8EC2�S���1�c��J>;��r����}յKw�_)�J	g��&��,��3L���~�ҩ�Mz�������y�����Y�^�j���j���KĴ||���*�z��>֯�h��|+.E|'M�lIC�Z��b��&�����$�`8bcfDD^<̘6G�	����ǟ��p�F3gi*xzo�t�~|�thA�,4A理�.�E�\(��O>ǖqd���r�M`uM[2�7z��>����ꔨ����+���ݘF�����*����=O�ԉ}�M�d�E�^68ܔDq�ֈ�x/�U��������s|��zh:h�5W۽�B�B�_�,�ݼ�[�\��Z1U��V�Z:��L���ո��,,}�X�����ۘLm�6�`�'.���=>,*��q�|�ܰ����i`�i����_���4H�X��$�-S\��NF*m��'���=�Y�f��ٰ��N㶶��A�1en��2\��g�]�I�΃a��-ac���Ws��]lgº��,g�)���>�E��gG�����J����5l��96p�!�E���)Ai܂�/EE��Z�bf�O���ۆ��דXJ��7�hmn���&h	��P�9<^m@��χt��q�	kwVX�Ψ'l��ߔM���DGާ�v�:�����V	�:�W��϶v�p_0��qG?g��`���
��\�>���fS�,�Ok9�{�.��<K�~�q{�W�*�H�t���ӎ����z{�v�.���]�'u�6t�����6�}z�U�tcn6�\�:�[�luE�٭���M_7�r�.���?CT��SK�o�3�����k������_����Tm�BPze��(�P4qn��.���	/�}��.���Tew,��u��N���)�i/�}9A���~s��O�����_E��6�Au\V���\	��
�Bԫ�Y6�d�w�F<�����@���!@�l�x❻)�c-�d��<r��/	�(f4���y/~׶s�!�*���n�`�0Ν�v܃����)�ⶨ�W�7��̿P}��[�x��߽L��Z��!��Pu	����R�,7����<B�'��u�c�oW�S	�=G�X��OS���5.��+<aA�~svs2������\��-qL���P�9�����DS��ۣcz�لk�5�9˧]y���_���K�c=(8���W%�X���<�+���Оdc�2���9�;�k3�m����{��V؛]"�w&@�t�ԥeG&a^�oH�R0o��׀C�N(�eU>�>�3叧�W�[���n��c�P�w�5���Ǧ��+���S ���.��XV�~�Hm�M.x��n��]Sj:���1JȮ*�,�����a˻ 0#iR'���JH�Q��i��~vL�v��E��*Y�g��s��G���O�F�xν�~��>�ކN���"<w���|=��{㑶�=�2kN��=�z�[�M�7g��p���Ȯz��1y.}��QUw̷�oe&F����醄Zy}���A����>�T�5��[����t�o:)�s#d&�x��fė���fW� =�1�����/�d[�HsG+�U�^Z�67�u��e7��y��&x�ǐQ�ws�z��P�A��)�C������Ϊ���
8�w�����FI��q\U�/�Q~��E��>�mjOn���4�#F3�(��zF�%�3�и���\)���Wk�N��xJ	{hN0�jp���u�:��s3jx��	��y�k������k8b�=�k�y�����u4^��	��TJ�	�=tn�R�/Mj5��.g:����������kqkvn�6���4�P&%:Ṉ�(�̬��W��Bo+:�a��`�eN)��n�����Y�SU�Aӳ��H�V�3 �W0�{�1x.�]�25��d�,Mc^)3����9��~\����=�S�;��<7�ױm���i'�,-�}u��B���c⸣#}~U�^2�
5���b�ٟe�g�|
���}{�̿�����g�+�q��F�Ʌ�59t��t&<E���VneUo1��R����@�|b�ٖ�m���q�^�<|G����	K���J\i%�j�2d2��h�u��B����o]���蠧��b�T��������K?��X_����ߺ{<�6}g�:�OS)�}!׈/u
y���
��T�;�֦���.z{�u�dSG�O��5��a*���v�f�λ#.:;\p���z�k��kԕQ��ٽ#=dB����{C'�g4M7c��N��ЭO{ps���X*��p�݄^J�l�ͪy=�ͣ�~����|��'z|�W>5�!%�i���ҘsP�]B��t1G|�kn���L	�k�}��ҍ�^"����q���gى�ʇ%�2���� �ȰQ�-����e�b�,)�Yp/�q0���@�����_n�����.������l]f�j��sTư�ny��*�G!��ϟ���h�1h�����F4���
7`X�[5��.�?	��m)}j;ҥ�d_9k�ʇP�ݾ�M$�rz��p�L���]q�=}�X7'�h��{��0Ɛq*iu){��� wP%�h<�'�a�s��0����@�祾���a߈������(�͆v���OOk�=	=��8�U#/.�&�Vv�G��R��=Q2��'�P����9�5�;�
�F��>�7R�J�L����=;�{�sw��%�������y���`��j�;$F��vd�T,��/d��0�px�:k���VcD�_�{�o]�*��S�>_{����������3̎m0A�~�'��(<ZcD�]t}O�C���us=��<~s���j|f�m3֩Q��Mٙ"E����M�c	��7ʚ�*���lyq��������s�9�=6������>y�!v�ʯ0��-�P9���u4�������=B>}^����M�s��'���lj�L�L�ݦ:A���K��K��7Mr�8V�^ ���{�����n�ı�wƳ��{f����[�n�hT�����{�[	����>\j (�)gS�c"��d��p�͵�&��
Z�.`��AJ��nЮ��;��<��Yɚ���9Ga�w��]��W8�Kp8��,?'{q�c]ì���u	��<��㜽5��k�e{#�k�Q��`m�27�~VI�4k�����jPn Ʊo�Y\9x��kMp��%~˩��N�Cf�.SL�yP���F4C�[��<�����zC�c������{�M����M�(��];�~>�L��\��$I�mm��c�Y�v	+��IK�}�R�
��ݡ�f��3O�帤��;��2��=嶭�N6oS�ry�nI�m���ey)�	���G��҈�X�c�(eJs^w#`�����ȱڂ�5|�ȓS�dӵv7l���衋�0��Ɓ������~�������>wV߻�vx�I/ A�-���[���Y��ߙ!�%r�,RQi�����dd������߶�o�ރ`���w���}]�nAn�)�{�Ԯz�3zFׂ٦�[��ݚfO�5�a�p��\; ��I�m�ΡTO�P9��A.���h܈1\tV����n�&���
!�c�h�˕�z}� �^�0%��gi5��>�K�GllT
���&8թ�\� ʩ�N��`�}a����=	}l�S�\��t�t�٬ݾ:���<�{�2�aJ.u����G(4y�A����ZzQþS�������m���%�<<]�YpS���i���,�-!9�:j�{�Y��:gb�s45>�(ɘ����퉝.��0�$6<x�LJz	C2i�P� %�m=��Χ�;���=G
w�ğն�;��� H��k�2��a�7�y�8����s��t���]�j�&k��}}W��E��m�Q^��	���`<4���p�ץ�����C9������.�s�i�ڦ�Bo�8��s����NY��*Z1m�CU�t�~�U|��|%������8\2�6�9es��|�_������</��S7B�Y�S���	�k��FT1��P0m�Grྷ���ݿw%Oe�����<�a�ƾ-f�F�,�#��!��iqEy`T��+���|��S�ۢ�=�)��b��HKsoC������U�m�����P%�$k��8�.b��i�h�4���'�;><ѿG;C�ۦ�>�l:[[_���1���#"WOQaL�ű�M�\��z��eժ腳½��L�&��{���p�:lf���Y��Es��*Qҹ�؍�a>Gg;���C�5RܾJ�N�����c�8��)�F�e��vz�������}Z�λ��B_k2*���7or���2��sn0����v��pF�0v�FKnL{�����t*h��75SY:b��yݵ�#�ҫ����iQz��t��ߘ}ϻ��Vã+&¹��̬���v����<^��I�`���ji�k�?�a	�H�>d�=�y����Dk�Q�e) �����I��]I�z��n���k������� ��$< �!p�����[ųU���ر�����"�S�5�Fx���{h��ЍN�jc�<l�Kc���3Xc��翇_ݟ�rW�j�����!��?ou9xwv��<�������Fą�"3�}:`S�1��ږ�6���R4H5XD���syR;�	w�Q�Ͱ������tx�P;����g�Dw�S<;���F;߇����K"�m���v��滶�;���R�Z\Ç��m4	���Ox�.�zo7�U4L}�Sd}�{Eƴ��;�1���6__����h��["�Ҡ�N�Mb���3��$�l�K��2�`��,���zC	�Z���P^��6�L0��P̵�dN���1�<IͿs4h�GՌY^S��Ѭp���dPt���BB�u_)�=C��Pz�,E�-�v��q���w@�ҹK���;0p�W�v��	_^�}���,[�>��Q���Ky�&f��Q���hw!2U�f�^in�����זx��0�~uc^���&��ly��x����؄)"��M{�C*��e^JV�zݜa.:k�����~[�U4�a=�\�8}=�H����遠�O�Y����Ή�w�G7P���bx�
G};��o�oTVU%ܡ���;�֦�����+/�CZ"=~a	8�0A�ϺKS����u��y��(�z̞��bz����p��d�=++T�i8��վYB1�����$2�N��'O�YF�řEsM���]6Ni'��_��4�<��Xc�{��zǘ�zFDfH �I8���gGga<��J�\���X߫:��3^�q�J"�|�}�͛��A�Uu�5���J��<l���%w��ߛ�m���6=m��Oi��?K�Tan��2,�p�L��H��,��ݖx�3�9��M��j>�9�CJ(J���Y�{�Nl�}x����<�a��=/e��7�}��&�����9?`c�^��l��ן��z�J�-���zx��r������Pwy\߻��a�=B��N'�:L�G�|麜�[C�p��\>�񝡧t&�*�S�n�i$�C�CD?;C3��ν�e�m��¸r�Q銾�n��XE�-��[&�~�t�T�5�o�y:M��[���s�	> ��g�����-0����ˡ'�{끗\ǋ�{7sS�ս��e��9j��.|P:�����<ZQ')eu��>U�N��J�X�I����"���&��[�JO�%�3��63���i"{�Tk�<�#� �7ص��/�aN�-yY���_pa�S'q�n��0w�2z׎��-f�;@��
�<�:-:�j���ה��z9�5/���}�����^}���!dy�)�R��)�Z�q�k��>��r��|=������Uy�!͇G!��w���>B�}^�/۲�oLg�Q���ش��^m᫁J9�]+��4�^bz<�g�5�j�y��V��F.������ܶ��e�]�@^���[��y�\D�=�ue/E���Ǿ#�iZ=u����w�W�.d�2um�`r�ì'�{q�2,���I3"\ω�(W���T|(��y8���$����8g�]��D��]�cDO%�Gu@�U����c)� ���>0�;���w'9*G��|�K��XF�X:T��/�uFGK�/oZl�;9���R�ٚ1@Tz9ܕcY�U�bp�Qh����uY೘US:��{?#���=�;�d�Y܆A�����0�О�?P��۫��H��7�+Ob</�����8TH0]�*�<L��>wò�u�ܰE�����;�A���׫ʹ�e���v�-D}#��Ӓ3�J���
z_l�&oA����ɦ������_I��rl�I�ok��I�u� qZ;�^�t��Q@�m3\�>k�s�s���~����������t.p�/Of[K���(�O��ɉ=�y��Gn����2t�ܘ�"u�`�_�����'d𓯐��Z���p>\ޤ\t����c�ǥ�w����S�թ7�ݛs�id/T��2��{�P1��y�Wnz�7��n�g׫̾�(X��F�]�C�i�P)�򐵶�<E\�v�0'��3�Υ؏��f�:f�&)���.�p�Wx�6��7;7�X�*^<���,�1Z{����=�0��O��pK�?w���Un����UZ�-����x����7M��񴬋O���R £��Wj��o�Hh�s*�%��+�k�jh,�ΐ{}��� Y(�Z7�AS��#qz�an���չ��P�Cw�����$/ÈG�ְ4{��xx��"��.,,>ˀ���;S�ۣ�/	}J��ݙ��7>TcAl�'����8ǻ5��V�e\�X+Y��m��0j�R���7�w�mY�G\gw	(��Wˊ}#�}98��㋞��x���s�-뷢�Φ�c�R�Cj�<y:��.�a^T���0Z�'�[�2v��=4p����ϩ���:f��8/E��#��Uܭ������\:9k�7��T=��||�g�ڇk�Y5t�K��Lc:�Sk�e�)8�ss��.��_2.�>�_��{{q̃cS6$����������+�.�}W�n�� jd���f=�������*=F��Qkon���5Ŗt\�&u��5}�fT&\���U�4s�"�P�j�<84����=2/@����n��x��H�;=���or��qO�"�j�����mo�t��뺕)HlK+BQ�ER�ٙy��F{H:�@sL���$7H�D�ˈC�Y�Y<�A�^�ë��1>z�f���ܾ��kMN�oU G���G���Gҏ��]�_X1L:�vfYl��1	�9�S	���m�������w��=�b6#D@KDb�h6�?[��'�G���q�����q��}qƟ_]���y��h1;��E��,LZ�u��H1�# ���m��q��q���i��۷m� ��I#i?�tMQ�[�������6E�#$H@���O��^6��8��8���4���۶�dCq9�����h�Іɂ�k�ɍ�B���+ Ȓ2b5B�ե�B�Z�����ح<�����4X�a��1BX�RcA$4��B�Knh���+}���(���4Z��Q���ﭽ��m|r�&6bJ�P����θ� 6%'.�J4	b�c��AP��r�I �h�/��}�uq��yUL�c�! \����~�w��U���*���_V��0L���m�[{	^j�Yך��C��o7���w�e����N_�p0����}a,X]����d{�.w�#����<��)�l�Q���Ce�{�;���ט��O� ��E��.�d]�=�7�o�
p{�ZFң�\�8L�+�q�6"_��;�%�g�
�ߧx�n���
V����yQ��O�]r�L��U��h�Xu���_]��r�	�  K�U�mpqz� �2��4H�סk\��:[+r�
!�2��86��iW'��+�1�]Au��k?��`����7)n_'9�ތa���K��zF?�՟^�-x���9ί9���'M<n.�Z䬬�ݮ�_�cc�^dx7�GPvv�x/��ΡTrx�թ�n͔˱	T��=���Z8� �4���_����+{��*#�5�Cw�	Z�k�@�w��~n8:�9�;}�
��R"�:���9�V:��T���n���T�6��vO���<ka�ltCs̆�s�la@�z�SE�Ym�F=Tαm���r,#�Q����������c�,�ͤ��������ӭ;�}O,���f<� �XL���k-�c������3/<Ԍ�	�xr��&�υ��UEJT>��,]
��V�[�}�)79��]Hk#����h"p���%Sx����.�ð�Z������D�γl�+�O1�w�~s�V|�^�k���S��ONR�ؿ-�͚����Q�����6��e�|]�J&��������quu'�o3{vv�� �w�a���[q�n0q�媀�LRz�P̚J�aKe�Q�-s!���7�n+(�����7�2�����F�T4Gg*���_U�hM{w=I=��,1G�U2��4e�;z��Y����
Z�O�0y�4; ڳ�Y-�%:5��Agt��V��\�����=��r�ޮ�BG����u��^�������oLݙ�pwl�╡/Wk'�a���^[Fd����,W�0�ϸ��w��q�V�c3�������׎z������=Q@���[����#C{�ގeB�P���L)�#��e��=���1�$��n,.:���l�]G�x�-��=8`X��������s��	�qv#gMi���U��l���+�/F�!� V_��Ap��z���C=�7g��p��l	N�K��6��'�%�ӕ����z~�f<��&D��N�2c����pO`K�cFaʓ��x�������V뫴�OBGg��#���v��ز{ȑ(���1��'�'�Cly���G�,����o��~ws*������X�Y]��K�4c��9����-���g�����|��<�}R����|=��{�_ua�n>�}Qv0^1��YG',�aXdD*�*e�׃&�[�Yx%�-+h1�Q'��ŃP��>��ƿ}�r� ��Ҧ�e����U	ߞ�d�A:{K86�ۙw=Z<Y4po#]M�|��yk�庺{��S"jibX�!�B��}R=���OS^ ��O���|���A���理\�Os���Ra}�2}��#���������~���p����mб�+��]�['s��0a�X��,�@��bJp���;������D��]V@���o�-%ܭ�oh���+��C��E���ce�C��,9���jNf���Y�P���[u��kk��s����gss8���x֏0�����]�>����_Ja����Fa�wM�����o��3*~�s@��E1����w��r� GB�/U����}�BE���%seK]os=��F���d-z�Pi)K�����g��0N�!!��ԓ�Q��w���q��Aؙ��LTtk�E�qxj܄�U�B��[�:cP�5B�.��N��V�Ĭ�v�U�9�!�H)�8�. �H��a�չ2�r��c����-� {���o4�!7X᝛�l]�Exf'��F�G|�{�1;��Eicx8n�����YvH�B�	3��x�ƶ��	�d��#Y�LW����~�)Y�R���7���������Ux��+w�
yT3�����U쉇��^�<|G����15�w�}��p��Ǘ��`����������;� ��b��T[st_u
�7!i��߀U�e�m��Z�Ui��+(�����k>�$���Z����t�:歸�ym�����e��`��N���f��SB���?�C��(F4��g�}]��9�2��O8vߴ���׾	�[���~��V�Au�P��>ʚ��A�1z�#��Q�*MRh�Fx¼�c�����4�O'�@yn��lB��v��ޚ8tC�F�vsC���m��ޣ��˜��
��b.D��'qI��T_9k�^u{���ڄ/�as{�
`��yʹ�7�L�{y��������醶������S��[���@��pY���1��z��`�s���ٌ-3��lo�[�ڑ-�"���;E�=�B�I�\�����c����%�î�Eыa~݀��3	c4.�F�҃D����͏��@��Ufi(�����O�^���{���G���>���{��ib�("+^n���׶��og,6�I�6]�w���s��~��#����7�t�<��Q���Ӽ���-��8@-�d$w���X�y��&���tk�=�:�מ�7�l3ϓ�F{O�cG���)�:m��}"�Yb{�I���=����̝_���k8o0�?�T�ue�K9"�'�_�""�5+�񞈑�����)Z�M3��eW��M���]u�Êzn42Cd5l!�]'H8:a�x�
NDT>��\JC�#��ǚ��0Z���Z�#Ïi���W���O��v�V��`��HB��.����d`N��GU�T�s�;�{Q3>���F�m^�����IQ���ݡ�^{�0�3�*�zvR<����6��VI٪��z�����_����7� `鮅τdL�[w����^�P�l��@+r�{ыv�z�M��p\�o�b�),+�3Z�O��7���]�ȗ�~����5v����Ǣ���f�s�:���9D�'��|&��sZ�g:����J�A�~/�O�� b�d�kίn���N���hFם��qu/�η5m��Gջ��f�9 ��?g�a>���]���x7N�v�|Q!�0`ǁg��:��Xu�.0iWo�7�3��ـ5H���X��Zy�܈�����E�쫎�i��=�8�}�[T��+=;�C�w����� �����Xc��	>2�-�7!���<xV�#�F��o@�ه��g���*';�2^o.��n�_��D��緁%�^�,��~���<pE��'��p��9�fH2����'�rVM���������-����u^[..ꔸ�f���߇��������p�ޏl��ko�����s�.�f���	��'��g�{���uuݣ&�D��xGZ��pړ�1��7�=�2������I�VQ��9�ޫ�=?z	�A]N��D0�S}`���y�s���`���왨V�guU����T�I�A� �_{�EP4|�Q���C[�n��o:�.���>j��,3Ax��{	�W��kQs��T"ρ��5�����0Ǻ���M�}ɱ����<�z]�娶���npm9�g��jU�ޑ��������tv�,������>���F��]�}�[�����mm�݉.K����jxҡl�U����l1$�o|�++`=O�X�&�qv�T=5�q�j�2$��E���f�L�w)bv��]��J�0hք�^m�����}��n��X쬯��:-��]9���z�J81j]�<̐��w�a��V����V��_1��"&�N�v��cV�t�.��i~jk��]��Li#X�J�%�M�T/W%��곻/>ڼj��{ۃg\��!4��1��|��&� F�A#�����D3R�n�=4�xJ���R`eg�'����nRA�3�xD|#�}P�[���;��1`C-�ژ�;w%�	$���!b�o0�_�>�<�o|�V:�09�.�^tl;_k��3�|3�c�<Gc�Zws.�r�� A[x�ds����,���A����Pʅu�QaMA�j5�]�E�wUx6eNu-���"z=��-r�"�nb��3�Oz��ջ����jz(s*T���qSV��H��`��[B�8ށ �+�^� 5�vS�}
���&֟t����ZRo��-i��^���{�v��S��R�TFb�<.��O�po>bE�^K5X9�jUs�U)�8�^_r�f��v�6v�QL[ɸݚ�1+�j��+AQzV��{� �U|"���^A�"t_^):���&�W�y�8�oOQ /�7U�P���g���C���a!�BZ�'��V��o�m��Z<w��y�ꞑ�rJzkt��
��n�u�,�yY�*���� w+s"凸����w�����?X0�{��ũ�W�IOL�%�\�:�'��=��F�x��.gk��w;�<H�tF�_�c�0�WZ4���}�ݡ�Y�j�)�fM���u�����J��pM�p9��;z������&8���،�j�M�x��%�C�l���yuRY���Y��c}����J2hP��ծ��SQ=�;f���硐�<���h��0�?{����z]���V_x=^y��ʶh���vǆ|H�J�x�}�m{h���ŋ�u�L�1qg|��h������<�`>f�j1���u�bv��ОqW��=�������/ʇI�����T���EN��0/N"����u�'��7_Z:�AN��w������{���f�S�Ϩc�y>���!-�q�9sx7��ky;�J�e��L�����p���s���ڪj5��t�ŵ>���/{ǰ�:b������4/y}�WՑ"�т�=�Y宎-W젒�nsgN2�7���ֱ�kZi?<E�ms��J�65u*H>�����>i��H����X��-u�ك�vw�s�~�<�V��c���(����|�	t�picZ_P��:���UJ+:Կ�3X�ɸ�yȆ�^����3�x��m��x�q+OT�󶠁:w�0Lj��n�#b��v��O5�l�-*�Oa�;���-\�^[�r�aNbˆ����k�	�Ј�s�j󴭗T;Nk�Q����ݪ_?�M<���)޺��;��~�1�n��@�V�נ9yw��<�ˢ+�c}[T����G �B`kdO\rq��z��*/���D7�(�*�0g`��s�7��/��f.N�Χк����+���_:�p9W.��i��o�0�a�n!�P�\]{�aI/W6�����f���u��R�X�N�1N�E�ܶx{7v�(��rs�����r0o\�V������x����������/��h���_�!s�Q;���B���VT�i�R(���T@�o�dݡޮ�cf����{\�|�ח��T�:�y����s�|�@�Tp��n���X����œ�]�\i��l�<uԿu��uT���l6F��8hG��4/j���R$�j�u�����XF\̫���K��{�������������0Ja?��F�sʵ���ζ�M����M:�'])�[�.���۾����;7���P�b���v�C�37{Mq鳹�˺��؆����ľ1���3�U�!��A!A�Bzr�?�*k���a��{�+����Sh��a�}0�Z}�f*�^���.��"�e0��W�IwPY�wvN�ٓ}��[���ն�����2S��\P���ήc�^��=N��8�@� �pZu,S��Z��܍S�㱁n�����9�_b��>��
j}a
.��y��?_M�aݑ�;8�@i�WuTU��2����ܛ���=��~��e=zޭ�=�ѭ�_Xp���un�]L[��i3_z1��\8?�K(�P*�,QY�t�o���O��ԴɶЇ��\��n�A�Z=��ec���׵���G��`��=��v=a�������my|��(s�s�2�l�g�a��}�<��r�^W��k7�+�Ny~e�^�����1���.��ott�p��Ƴk�[}f�'����GlM�}w��\41YZ��|��<�;RqT�L�Βݥ��,:�PrB~H���]J�r�����=$���u�?��v��������[�+��8K3 ��~��szl��iu�~*�m�%o�,]t=Z�l%�rr��_-̈^m�m��Oõ���_�z����ƁUǲ���d�V &��t�����M��s�kq�܁3��/�6�s���?[Kb����@�q��Ťqǀ��e�{�`��[�@$!}�7
��WM��H8)�3�t�k;2��4�S~+�z�T�+�s�����/�CL3��U3L�i�ۦ�Tݚ�mJj+d��il�A"@�N���A�}u�|n�n�2ۜ��)S?wu Rk���&+2Ҏ-F0W��M�βr��#�៸<3��p��4�C�`�S㰤� a�t�>����	�Y�.�3���Oa�)V����Q&�q�]��.L�j|��L�3;#|��o7��_�M��u����Qw�y�t.PE�v���U�#�����`�ZoP0����œ�֌f�۞��{լ�*��FOl�Fh(\�H���Wb�_z��s�-=O3�R��y������ilO&zq/S��Ӭ(���2����S�eᙙ�ܘ����uz��ށ��=厘�B�{^�No��&Lv8!��)z��,u�!���R,~�OE��z�#58�2uۻة% C<s'F�B��^>~�yj|U�	�_��o�)���\l�r	Q}��{�Q��#�x)v�Zlp�2�����e^�kd��f?rK�?c{�{�w����dO?�`�-��w(*����}um�����T����B�t#�S�ۻV�y-���幧/F�F3o�c��һ��|t�6��\ih��0�����5;��9�KS�����sG)�҆�5&�:IۮAQWUV�Nk:6ꂇ:�X�A���H�`��X;	g3�j��&������K܏u.�n����:@wT���.��ll3�S��x:7R.�10�{f�,`����� �t���[sZ7������W>���X�}�m^B��TZI�<gUVn��Q��j֟Y/���y̹�P�������'�i�{)�T��}��3�Ft��e���T6���w��2��m�X�OO>��+�5���<�D.Fv�J�\�}e�zx֘��D���[�L���BaY�Y0��;��f���_�(zc�'�r�㎎��>�x:���v�L�;�[X��}�'�xq(�X.C׌9��;g�ֻ���|��o�ژVc|�5�q�s��]�R6]��;8�+���sئޖo��fh���}}�|۫=פ�wD뼳���v�s�>�Et�n;~V]BMk��8���1Z�d��*�;���gX�<�3]|�Pg��1�$�Q^g�\jf�zwq��bD�[a[@��;N��jΗzY��VM�l'����A�F;���R�����y��/h\��},0�P�%͉i�W������C(������L�e+�q���_EWǥ��p\s���i��L�M&h��3w=��^t��M�"�/qj8nq-��XNd�w#/b�ai�ߜ� \��n�zg$��T	�+��i�LX��U6�v�[�]��Y���zj���uȠ�y�L��w�v�b9%�i��5�]���9����f�\M�V���%�W�=b
=��%��Vo3KF_��~���T�=�7�v.���O�g��P����F `Yۡ�ޝ�{�wne��{�S*�3'���Wnݭz`������}}(�"�;�>�+��K�I�<�PT��㷯x��qӎ8����}z���ި�Qc+���o����ڿ���L�v�����s�q��o^���8�q�ׯ���N�ms�W�/(ϝ]6�~�.��d�B� �e������i��q���ׯ_G׎�3�b!��h�h�O��65$X1i"� l���$���W��c�nbЅ!�>V�4^k��E���ի��e��E|_V���E@h��EI4"Lll���4ʓ%F>Y�m&���n`��5s~��i^�4�&,X2j�Z�R`����H�ʈ��r��Q���r���'�߭�6�E����!+Ti5�_�>]��$��r&���@�Q"\P�L6�0��(A"	��Q2�(�*Z�7����,�f)T�e�['b� ��֙���{�zn��H�����{S�B�!p��/# T�o��&LI�H@H$2�-�
D!!T�����!���B���h�� �rE1��F���f&q�A)��mđ�B�'�vU���]J���5cDi�)	�f	~Q��Q�;5�x��n���'EXn�T/eĎ<�ßO%T˰���Ѧ�%7���'���L�l�~>����t�uy�U�(�s�W��T��:��o��f��a�������:XQ�(��o�o+fusS���t{]O����]�ø�u�7��|e�ݘ,����7*���Xn�c�d���;7�R.�M���T�i�z@h�d�q6��5�D�[t.*x{����Q��n�
�aJk�Ǖ	[Բ�f�pY�����M3��ey�.�a[��m{y솼�K:���j�|�i�6.��$ׯ3�ѻ�yo�3���t;kH�.dw�纇�q��f�,�I����{��ɴ6�h�t�n�ֽh�}���:�m�2�Gh��x�K�4��J��IVz9�H���e��p8��,�M��: <��RE\�![��I�bT���ei~���l��ϱ�2���Q��l�e�(��������G�IO������ﯹE~�x��M�����h'�=��+�\�㣯50��K=@U��E�̗��VKq	%edwku��=cf���=�g�e����0|�&�qBO��q�1��4�� ��ߚ��k�u���>��Ы��@+}v1u*��WV��,_��l-���Ff��73!uY�@a��zE��0T����(�����&MEE������SoW\c�B����#~b4C���{��g�.��8mWhV��.q�Fu
ֶr.J��Tr�[9�S���4W�&|��PG�S������{Y���6����5��'wԐ�J�	3����?����M���HΊ2�D���o5D���W�����(��B��%��ʆǱ�s�t�v�v�tE�=V9��wx0��2MO]G��y�¯����M>��h�=J3];l����V��e�tX�k�+��N)o���Ρ�J��#m�7#Sdmܙ�������d��}��i��l������]s��E��W�����t[��v.�9'K��ˬ��-�[w54�5l�Ǻq�]J;�?fFE�!����Uq=ꕘ�X�J����Όzx��}	���O����w&���\��q�b�T��5m����ю��v����$�w3���%��U�ͧ����_k��yI�����~���a>���ox3�����-�`�g�F��FF��Ȭ$�����^\@j��Qƽ܏P�]M^�ڸM�馀n���YQє� �n��=ۣ��+`-] ��:�;eJD�u��!��'\y�*ո���u��Ӯ�{:QǠWt{vOu��O�v1��Ӳ���M�Nu��-��7Z0�n�n�,��&�c����{��*�z���)���U�=a��b�eS���w>��D��h�p/�h�a�t�Ȃvw9U%�'�؝ֈ��a��%&ՄְA��z�o^�m3�0���b3����j[��.��U�ob�]Ru|�b�i*��9���+���`�xLVP��f�/C�0�8K	W�y�V���Nϵ��Ӵ0�+���8!3���אkY������U�y��K�$/v/ww���s��
��v�/�%�nL�]��;�8ޏ4u�E��v+hčԥ �Pm�[;�]��\Xf�kh2jv�f�����7�t�'`s9�OE���=yu�U��>��=��V���9�8�J��>���K�|WE�T�v�����M���T홯3�㘥:V#}<Bɇ���g��-��ߏy�3
G��r����#Lơ�f��~N{�{�|�k΅o�>z���T.�u� �!Sb������d�25Js=7��W
����]����Wۣ�"rS��J���W�C�����H^�3�쳊�����v���4w4L`����LWe4F�{=��xί-����B�&=s��2��PG2ni���qÀ�d����ӽun��#b�8�O3S�Uw��c����[�o�n1��z�&���}�� I� ���+��v&���ur�]ˤ�;pX]ډ,/{52r�U���K�]y�۰!N��h�GX�r�U�S(S�ܩP��}Zo��^�&=�^��mzG��u�#e�v �Y'�T��]&{��"*�so/M��<�yfף}�j�BL��Hh/��OF����ux�DM6)	n�G*�%D�^���L�ǀ��e��f�}�ߊ�.ni]�|nx�r��-d͕͜��	(��ڹ�D ���9& �}U���o����e�^�ʡ�	�<���Ŗ
�.�`�̬���U9gZmҖ(�*�m-�!�b�h�!��g��pP�瑀�3��I�%|b�?S�kr���������mz�{�����O.~=�Ûc�x{ �ӌ"�$�3���vl�>UЪ�F�8�!��xt`K���>5�4��74f��f{Kody-�^��D��4nwBfi0��yk��H΋L�H���ǫ�^���{$nwNd�)��b�ۼk�pd�k9��n��z��,����?��^l��g]g4ă;	�����dQ2����5�wN�T|��8�ڄ��+�C�.}�2 x\�\� ,��O*T.�юҶA]�y4y^�W�[���XQ�(���WOR�ŧ��Ι��{�zg����w7S��C��u��u�Q�����l��Θ^��_
Ӱ���z3������^��T�H�yѼ�a��1��7R�˝�>��10���p����O*��C
S\eG�J޼mor�L�z����7 W
�x�goG�ϣ���.�xƗ��2o_��7KT>f��{ҐUx��#���y�;wE��6�#_�~o`��߲�\��ʹ�v~�����5��L�dc0h�W���[[�3(8o��y�M8&`[��`i�^w��#��o���eC���w;
�Ng��d�.D7u��M=���G���|@��5��䫹<᪸a��'.}
�T��ߗv:/�7�Rأ���S�>�e[F�⦚2�~���*��*|�;-T�}!���A�t���㌇���~ ��'��n�-�	�����=��9c�0LpW�(>\T6�C�mzB)^rm��=�. g=c�l�!J����|�]����º�<�OdU�T��wP���P�o7���]W��WV��*�����7yWZ2��{v]s1{�ܜڥ��G{{���]����a��U�m���f 3x+��;{���㆗��Pp���0hƥ�������j̋�4�d�; �)�gF�+�ű�ag��P�����ٍ-�j�z5e��z7w�i�! �+����+G��XU�h��]�^Y�sw�Xݵ���>���z�I�O��"����U��m���S�K�sJ���"�������ń%�g�J���f�:�/n�Y�}��� ��?w�t	�g����ʙ(ӭb�Ù��挥cy��:ݰ�UZ�C�m�w�.����q-{FWg( !drY$~�� ��^\�B�W���ȥ�赳@M������P7�é���,	�Mr�1�n�4�L>;X<����;�_r�]�*ŗ{m.'nz�t�+G �dn�niԍ�p8o��&N�����3����/j�Z�So6o4��ҍzOO�n榜յ������Ko�Gg���Ɖ��-Ǧ�vy��%x�I�x�u2��*ci��\�.寧������6���R�BJ'���Y�p�RH�A�گ@{�S� ��]��ܳs7"��Dhp�@��h�ԫU&*��Ҽ��|���h�v����3��|ǚ^�p�;&4����ʃkbF����އjT*e歫�c��f�Þ������`9#��.r@����ir�^N&m�5T���,�Rlt�
����z��<Ê��4���q��$��DU�'��~�;��I��9_����c�`�����w����_���U�č.�b��;����k�9*#oSe�U��x��T>���N�"��k>�"�?l��n��!V�{�n�ј74wV�Uو-Ŧ+��M{n��G3}�8p��?����� ���J6�\/�\ipA��TWS��@���_V��P��<�Wa2mغg�P��E�:�D!wޮ���A}렊���#Fm-��6�Ӫ#^z�UZ+b�K��}������w�=����;�=��Hl��j�+���37A�p��d<4gG���2�����@��1:���H�F��d�`�U�,��)M�}7�3�����t�9]�7=m�7��EC_D��77c^�c�U��笃�/��_X}�w�`�ר>��\s-q��t�p>��<�Х�����������9�C���6̋��^��X����'kD�N�Mv�SnV�<���=s�5�'��,ˉu~��:�8�>T�ӭ�ڈ���]�=�[��v��<Ce*C�)��`Ywޠ��@n3�fmt�VZЭ[�У�p�D��+�7#�k��o%Ԩw.�Bw�U�7�c6���!��1k�2����L�E�!T����kpEb��ƺ�{�h������s�mb}���j��g�����	ٛ���@����?ʱ��w����t��5Q���϶׳��SS�)˧��* �2i�A��߾����_�՞��Hr?�������+��y�����<H|2ḿ��7N99��L=�`�z���;QS�a��!�7����7��� 5������mӨ����=�F��"+5��t��-�=|����'�'��e#͔2y.�~��"�'*O�n��8��D/^�m�6$���O|�voe��f�a>�m�}�$$0���lI˨x���5H����z��G^�M�Ua�A�l09瀛CH��m<�8��0��O�n�G^�ϕ�}�K_�J6������<��ˮ�� cz��3��8!�a��pߧֲw	�Vz�L�2M���U��rw�S��"���9����*�#݃Jm��]�f��Y�q�NYY1�ݽe$HC�dm1�� b �e��u���`�����Ɋ�M�{�I葅r�3ڋw�����&e�~�����<3����QŔPSz�<�~y&� �m:i����ݻ�۩u�D����3��Rɵ�h�sGN�hY�%2�9�B���ۃir�:C3�5a��u�ea�YO���
F�I췲��&4/���0�O�����7��y���FX��W,3/z/�j}S鄺u�����ݜ$gu��o�e�X�F��EA��l�.
@���O=�ۧ�=Sᖁ�EIH�hF���i.��T���	�퇺�O�J��~��{���1�S�4:Xh�:�j�wZ0��z�lƘ��X��N_Q���~�n
KЮ}���!� �oW�0��;ҕ
-3rzD��^��ݷU�5y��q$�ˢ�����f����t�����,s�˧��t#GiO���Տ˺��yqZl솪u>�>����>�}�6�,�v٬����Ӹh�5��-lm���3�(or�g��a���|����h-5Q�+)��q����C�?��+w�n{s�W��������u=#Y�N�d@����K<��?v���:&�I'�P��WV�%��0�P;��ó�c"_0p�w�C�D/-�u�VHP��ģ��5�1��������"��O9�YDpc���Y������N����/nD<@Ϩ�jvf��Y�L�u]��]�
�]Rbo������.�m�c�^Kw�7� �9}�[G�+����Y��p��}ƚ7��̛��o#v^ޛ�JȄ`nqFӮ��෣�B�i��c�/�v�;�l�OȲD�s���u�s Ƽ��N�I̳E��.ۅpQ�o�%@������;��߻�.x�6h�Ѿ����<��ho-`�]�e���5`�_oC�ݚ����Gϼ���#�n�����h"H徝N�~���+aB�,�y�{��a`�KS`�4x�*S/v�
u��>��0��u짖L�L"9�ǫ�r;jL����������8Wd7�8O�n]�=o��:��p�&{��E?@�?G�{0Wp*���bH�R����fa�g<�ɚ.N쯐�N�^��"}�5�+��������nӾ��ǡ�C���ѽ9Y�3�tҟ6���t���
�3��UM�ƺ�gFF�\��oh��򒦞ƨ�OX��\��_e��#G{��u]�sz,pt"��bT�{6Dֿ3�,oݵ]j��)��r^v�K|���E��wo_H�:���T`�U�r����#��K~��������5u����2�� �&D���.�>�E_��Ǻ��4Q��c�C����C���}u�+��T����MV8�OW���/� c����>;�/_z�U����R�a�<$���r�vռzm������f��Yk.'.�U�M��n0j��ɴ%�^i����C����&����#{$�Si�O�df�v{�\Zؓ�#��7ݞ=8�Ԭ\�8��V�Vr���gǖrŁԕ{B�D�7�vj�VU�5�N�8��v,Y��5r��T)�؋(�d̖d���i��A��a�mD^�J1�{ɏB�Qxp�CX�G�W/,��9%���sFݻ����ǉ�d�F��������f�tR�.��C�HfJ��=�S�����E=�И��X�Mk�:�_g-��5u���w���˽����p"S�7v���T�*U�q�ܥ6�Yc5���wõN��������Gu#���GN-
D���KZ�{<y7��+d�*Gb�T�pu��fY��t��2��IkkK53!rV�Y��Ẅ́Z����rwZ�j�S.mU�����)�OE7f���ȝ�T�\�wC���nג��Q���D�����<^���<�\��VgU1�L�n��,�^�_�b��=�qខ�y�^�ҟ~a>��s귺$�)t�&3`�s��/����ܼ�n	t���޲�Z|�?OA�xf���L9����C�3���I��I��$D�:���n8�ǯ�8��q�ׯ���N�I"ȦѴ`��sr�<�͞���O����_Zz��q�n8�����~o����+�snQ\��ܮs;�&�۩�������8������=z�8�z�����Ӧ��P���+u�W��7	+�s��M���\��cW���B��r�r�����&�4k�S���/6�4lZ����z=�
������tb�K^�Ot\֊�qX�M�;�EE\q�7*6-4Er�ھڻ�Y#d�6�[�=�\��W(��T���]"ž�5y�s�wk��Qsn�-\wm���*J�%P�%���9/y�L��~����؏��o<M��l�v�>�Tq���l�2s]{����Z���]���˃1� �vё�����Q)��7�;�.y� ��ab��#���g9$'�
�c��}���4<8�����w�������@FH'`�)T@�#��q��vr����u��˝�鲕!�̽諟2��ٱ�ǘ��NtNΫu;���p�Ǫ�%]�ٮ)��{�7��F=]<f%�!�&���y�+�E���v����*���<pa���m>��ށq3c�\��;�7���z'�f�Fu3�z���h=��p}P�^dj�K#J�n�lDQu��N�����]s:�������o:��6�����j�Y����.��W�P�R���݂��Ar+$5�����ޠً��*�5�m�D��V�8+��YA�ޫ�����)J�a�81���p����ǻ�J�����5�y3��4�P������gTk��'{}�zV��.�ڽL�\g$�X;��Z~�".�m��g����H��z��r̂�qr�8��ݞ��x�#0���q��o�|2r���;I�A��E��Q�������Ώ��:>�W������r��eU���P:9��>��l_wl���9�]��|޾4Čc��7�o�;�~t�-��z<z�=I��=���r�c=�W��z��9����D �|A�C���Oƒ�[�5��ś�Q���#[9����ϧ�m��t���e�R�#h;����U'EX�wJ�^��Eg��GV�[������x⡁Q����ι�e��Ѫ5�T�di�w��(;�˒����
���mq����0����pk�Z�2�Vf���T�El������+��h��9�1�!��tM�W� �W5�_-�\̂A���%��cӖ�ݕ��M1Wn�ޘk��8�x�U��cn�φ�y%w>V51׭�J�,�m�B�ӑNg���w���u�ݧW=_Y��Kh��f��f�y��F�Z:4��˫Gqk�o]#��`�U�#�����9ِ�����(&�UR��=����g�]~N忳�����ϳ󲚩_�zN1":��lE��uc����
��f������[��ߔ��`Н~���i���n���2g�{$��ٹUE�ݣ/���[��*`��<|���������ps�	[��W���������*��^-�N��F�"�4�=tNY21ݛz�\{�ìwm�w[^Wtݰ��
�X����yC��͞� ���)�pJ��V��Wл�)�ݬ�{�.zr&� ��j�(V\T�a��v;TUz���i�2�.S�k�^[��ɧ������cK�6t��3�ß��]f���?#C^R]H�3��n�����ٮ3���S`���T]�5��H�ϗF�3�-�{�����7�89mC�������̤�;ƒ����ѱ'?����`I-Ӷ�lUE	zb�>��Xyt��o�ެ{'<�%�5��97��ULrz����ne�z6��3�v(�q��q<q�����f�q����7V�|9!��m�P�Q�+ʩ��/�f:��_���Κ'����וt*��m3�Au�==�et�������n9 �nTv�_�=x��"j��I�ĆmL1��d�z�̀�;��&e᝚}��5\�g���S�<���B��{����f�`��S��uV�vίmV-�	�ˡZ��Nn�]�+cr5�ܮb�A���rb0�P3o'���㢾K3_����$}ð-����>���+��/���f{<�����^aª��P;)]��m�*xl��~[���=�DF_e�4[e%�M��ai}���!������{���do4<�ys�B7�\�gi�g���$ޓ#P[>Ho��1[Lqہ|u�p���R7t#	4�M7�VQ�eu.A�Re�\}�n�,(�ml���mP.e�j���`���ͯEs"��m{�cF;�_`_��Cm���u
]�OF�(Eh��Z:oRm��D'�)y���]8�r�2(�)`���z;/!�����|@�o��ziZ6݇� ����x��MP�сTH�jx��]f�[�C{�;)1'ԟ�<�u���td��6��/3/xv��]I�ow.dV����vN��,ȑn;�}�$��Q&!l�|�����c����fhNq�<�1���⥌�T^���~�V�c�9JWQ�1���6dl��U3A�ȡ����DΔ�n�|���|��,׮�)}}:<�Y�!�V$г{��h�Wa�s��j')� ���h�A>�yi<�7Fe�AТye�'qӭ��u���dT��ܒ�G����|>|>
�0�ԩ�e���#W:ʳw�=bT�C{���K��2�+���;m���ߣ0��C3PI��teN�F/�j���)���R�uY����6�r�����ݿ.㯾��"Lxު'� u�=]Z�s�l֛X��������Y�/a���BNt�cOJ����ɛ<��Sb�d�w�!$���=�;&��}���\8�a�m���p/)1W��OO��Z|񷢞1��-�JU0�0>-MYf�Њ�X9�M���)�O0&T��į�����7=.]tc�^��u:[V������@��xU�6V�=]>a8$�G���';�vf�D�������oZq��Mz�����\_�f��Zș:�3���DM�>���N���w������smzY��q@���UC��������-���:�r�4�Y\�F/b�����q�+����68�䰋j[��q�`8��78*]�VW/;�1�!����ܲ%ۇ	�T�q��)P�u�p�֡w0��ӽ:���{F9�E}5ỷ�'gQ���3�9�?|~��>}��gM2�U���Vl�%m>���sN��,��9o�@J�ŭfb�l��.�5z����I��C�IpA���ϹtwA"8ܭ����zò�z���X=i��~�s,�A�����S�lC�Y���uG.�ګ��~�x�t�Z��G�����;&{�u�N��3>���O0�*y�h�y�i�Gsɵ҃q/)3�PvLo��ǩ+ݓ�zyp�FYSH�s"X{Ӓv��(��� ������]xP�`Y"3���~p�k�qoD֝�� �l��W����eO�����*G�yL u�Q��F�w]>�u�b�Ӱ7-xO^�'�Q]�D��w�w>��!S>�?�L0��{��wD�dWj�z��iVz���z�J�ArU՞��2v��>o!�"GZ�y���dM�>4��w�n ������l�%A�20���r^\N��16,��]�w�_<���{LQ�2+rg�fb����ם]�)n>�f14�����BP�][�\{6%4H,�������6�oq-�c5TPN�<�͞?���yz���l*u����m����� 㪆�ֶ��5�� �}���|=��?5�c�{9�L�re�o.��]Teb�������vۻ��%����е��I�N�k��^��� �����{N	�I:W�0�T f� �P�֪��V)�������Ȼ杭��͗{VX�P6#���=���У^{�]���z�-�I��c�n&Gh�Һ{�	�Ee-ysy1�`�9�Ur�Q4Xuکj77O��aиq �[�;R�_u�-i�}#�MѲ�AZ��)#6�Sq,�����D�>ʟ(�R��ڷE��t�A����̸�S+�f�Slk�I���зA�vdj[���9C�^\��8�e5�{����3�V�f^�7�]o�V� �̪Dr�G����b��s�^�*��}|������kgf�]��W�lܺ���C���K��Y�"��xFm��L���UU7h�*�l���2��6���������Y��\�ֳ�fX�;T�q���Ǎa����<=�M�&���M[E�E(�$��י�v�o�I��b��Q���"��s|��Ȟ����{o�ޔ�ټ��X��^���Vv�5�{�Ƕs�8[�h�n�x�$w����y��z��2�ꅎ����S�Oj��}�k���J,EǸd���3=#k7[F'z* Pdm���ĕ>�<;�����]���=<���u5��*�s���I7��?�XW� �s�=���K�҂��۪(*�UXq�u6��n���M�<��
�8ێ�"6�G^ƭ���~���+��4�HU~�j�iP6W�딆[�����9����.�6��oԻq��.p�6�d_qM� ��A��=� ��a��y��������ԝ.��#���v�u�df;ҫu�ݝϣ�i,�d�z|�����gky���t33���
;u�.�l7�|�S+������
"0痟|`ڵ�hI�ؼSYr��W�/u[��v�E\Ϫ�QKhn���wu�l=]�)�C��X٪�v��ОGt��B/����T�f���;�>�o���3Ɠ��~����r�=>�xF|�^�/6U����u�ٓv���ʾLT�OHU��}4���7	���M��:����xg��+�Ɓ۰uW�=c�#�������������ҙ̟�g�����k�'�������Ix��#�ҏ_�~�sH>��}���箢9��k�!��UC/������;�~��Vd���4��i����w@�"s����T�`�Q�Km<.�\�L���ǳ��Eϣ��3�2��+�qb������n£~���svy���qR�ge��Nf:v�/���Ib�m�p�	A�X�����ۃ�-<P���i}�d���O��5�w[���R��K��\8�#��v��*���)��Ĳ|�9;���ETY�7w���\���ny�0�3��vDީ�x��haP�O�ՏOb�'1��f���36�k�c
A����q�A��U���5N��<m�l��w��gy�W�pV�rJ�O8'ó�ʪ>И�4�o:��&��ӵ^�р���ŲT�|���;�S�3ڣ	�}�PV@ ��vu �SQ7��zj�w���"��*�ţ �K�y�s��a&��|)��ɽ�1�B�ϋ�!}v+��T�Wz�;�_u��� ˴id�]��{$k^�{�=r�^1g�>��V&�.ܮ�e�gl�\*l˾rςz�1�Gzߛ��7�0��x?����j=iX�ސ�"7Ӵp�J�	�CI�av�۸y�[�Ak:���J�/l�`�������
L�7�{���L۲J�`�OO����?�7������ A ]��E�B�j|c�t�>�Z[Nk�,��h�|�.���Zx��|������CJ�c�S2z�����o#zթH���)`��R6Y�UL\��Y�naf/�� t"K�6�lf�@ՏI���~�J<�wqn���-��u�����j����Ūb����!���<�s�$:������K{��?�cV]m�g!�m�N��7U�������ё�¶�DЃg�����K���n�͹w�'�[Yk0�̈��޸TR��̨Рq�Tnϼ{�����K6F���Ǹ�⽝���>���Fp��[��k��"�!�݉��� �����5ps=f:.b�׻��������4c�O�b��S<T1��WqX��yS�����^�%fA�[���h�9�-T��ϑ�-�c�7Ʒ[k�!8�H��nҦ��4r�y/Vξ�7``�
wOe���\%Q4��5���q��{t�W����כf{���*%�VC̶�vF�d�����|ϟ�Wo
�νG9=��������»ѣ�s~�@tY�c\X����|���Zu/]g�z���?(C��=����(7�`}{��\��A�Vc���z�ϋs�3�O NL��#}�ȵ:��+��n��pr�C����GW��[)�Q�x���.��i�{*�U�57ڽeδ�����ھ��x�a%�7���\O�@�,�wd�yma�}�s}���]���{k�� ې�kn_`c�6�)�*3��B}���٬�N_��oyS���J>�4fr� ��^�S#c/�"�V�E�����8sv#���3����w������r�g��˱�g�;d+e�'Ω[$nTח��:��W	}N�+o*�R�h�D�ڞD4V����__Tղ^^�E���9A ����^ElaP�u�pۻdŹ����sC���[�y}��������M�ZIԋ�4Tk��;���h��s~��� ��c�
������5X��.��Ֆ5)�x�$����6�fA�Mf����;}%ͻ�
�#t6�Įϩ�V_UC��g�y%<p���0�[C,��@�v�:�\#�l��>�#�?����r�J���=+��զ�-gSm�P�������4R�G�\��,�V���3N$_�Bt���]Ԟ*�yC�a�Ǽ�K�� ��.�e���{^5��3�/��u��Bo>c���R�źuroq���W_A��x����zфnW{��Ϫn#�J�x�"˹�e�hȮb*vs�ޏ���|���:H��7�w��x�K����ǃ���]�Rvfh��
=^q�o#Gob���4�ѻ����YAX�yD��N�_{��q��(��֬��ۼF祮0 �/Et��pNz?�{8r��ߦ��<����[u+��y�����:�/o��=��,+/� �J�W�����[72�r��)��c���o���	�7�<3R��+�|���c~�+��!~u�bol�K�rT���{��aej�9e�WDӨ��������P�}��Y��Y��jɬ�ݍT7���R���RyX�y�un�^9�������GMѺ��cn`��
U�U�W�!����4����]Ԇ����;WY� >��S�>��ѭ�iMgt=S�����Z��:��sC��ݕ<b#�Y;�\Ֆ�>�3���Ŷ��}�u��y�o�r�t�x d$Z�ؕt�Ut�xƤ��BB|�\w�Au)�Ǐ�=cǯ�8��q�ׯ�}x�o���6�+���~�Z$�wh�&������ž{�7�}o^<}cǮ8�8�ǯ^����:h<�5����[�7�ͮ� =��y��%<}}x���=q�qǎ=z��}v��KVT T$�Q$���'v+}��yQo���+���+����y����=��nwUȣ___/_{�y�N���R׮��������|sF9j��弌����yͮbƯu�1��;�_?�W�*_�����j�K߽_�n�\���~�|U|m�r�k�ܺW1Qt��N�b�[sk�*�܋ns��A��h��~���^��_~s�q"�(@2��*��� *.8c��PDB�L��
tM�k�Vh����G�;�*����iܝ �h�x[e�5�z{��E��x
NM�!���^~�h�$��HЙ}���Z,�HTШQ`�KeH�&P$����EK��#P&QO�O�n"CYA�Q}*'I|�E�i �9!% ��H4ۄ�b24q�Y!�ۅ�C!+����#<����u�����3�(�g��ɲ�
`w�^d�}Wv3�.x�>U�w5w)u9t�W�U{�ܔ�Ng�����i0ò6CuA������&g����u�S%���5*��ܞz�D�-�W�HT��f��4���#��ykљ��s������撻B�f;�ղ���� ��ӡ1��J0fq�*���p(�H}쑯�d�#�+�F��_!�Z�VUҖ+0c0�H���ᢙ���j`u���|�����9 �8w����e�w:�I�0
E}�z���'��w��C����P��d��Nb��P�_�஑��u��/¸��۵*��M̢�>��h��Eɕ{��O���<*B�5���lS�,�X0�>�i�&r7�������ϗz��BU>�y6V�*ﺇrƑ�}"�<�1,�o���Ņ��Z��㨌��}�e7�v.��^��^b�Mtm�#x_X��x�n����f�r2�\�V"��??'�����Q�+뽳�N���m�i����Ѷ��Nx�M���{��5��+B�wUBe	̊+1$\l�%X"lޘ}�	��]���X���(��w����E������� �o7��b7uBr�<��,*�B:��Ll�5����R��Hؚ�����w������}������[���E�nE�6uB���V�V�uu98�^�����C�u1���t�#S�Q���)���q��RI����8E�Ob����"���[Ƽ��l�=�î���Ǫ��-�1�.���-&�^�`#���UǬs��y����5�1�V�5��nr"�N�L1�t�i�1���v�bh��a3�����t�'�7�ʋ 1}ѳy�W��?t���z��z�)�������{�Wk�T�W۔]���)�*�̬UM�o!�|4�\^�����?���{X*�Yop����^&�����$���Ӱ<��F�m��{Fy��c��@�F��ae��u�"6FC#K"d���/˙l�#j�!��|����F�����X�r]�Zf�`v�|���~>���ӈ���sqg �����MN2�CN�ҵU�/�;���_���GQ.����d�C�%s6k��',��k/[�ƽ8U��yk�ʩL��|h���f����^�%8��ܪtx�I���|||||=g����K���q��F�A�pI�cc!�p0HXR�����)�,6��g��������f��E�ҟ/��\s�[���|����%5А��G#}yWWElzu��
{�D�1 ��n�ۍ1����j�����i~�V0gM���M���*he�O>�|�ze�+g�U
���nsˎ��7�q3��:�:f6:�H�?O+�?���a��׾���o����}0�+ԯƕ�G���V�E4�M\��s���h���,��W�7K*��L��i��6^;��t�*�>_nS�R��!#'NNql)�oz��D��\u���3и�S��N�����%�a�w��z3z��a��\A���t27���ۃ���W����g���mf��Ȼ��̈L-�.�r����U^8�M]�^'P5�j��ز�)ւ�/�v����w$\�z{:�~�_tΜ�Ե��e���k/"(�*B=]Z�x"�۳/u_QA�{ٚ"�s�u�O��N���T�Nkf�٪�u�����������$����,՜�\�|�<���0#ߚ�w�v����<0���3����Yo���~�]1f 7����Ku73Lv�N�������(���^�iw�`��i��I0s��ͼ�+*cә�v9�����l�
ӫ
ݞ����*h&��{wve��FoW5	g���m��f���R+yH�\S�Խ:��-Ԥ2�:�����M�2��Hf�|Ωt���Q�^Jɕhz���,Nќ����_6�;w�{j}��J�|��^l��x���9��l!�k�b���s���`J��2/��(��M}z�¸xd_f���8v~��PU�������/^�{'�A;͆�(��H�g��;���s'��i���[�x�CngWn����6�W��z��0��ӒԻj�72-!%S��O]U#���F9
��}��#���|���[��Ց/���5|�jZ�؀�P��~����_�H���tc��~d�/��ܭ��׷X����������v�4m��YU�&C�ovUC�dL|3�da7o`�~K�W
v(	Ʈ��Q��NX)�v�".u��.W7���D+��gw5uR�6�0#�{��nh�G�d����t�����m�ލi�5Nٚ5���o���Z�y�8c��G���u;��1���L��gt�4+,���7�u���G<�'OlrZ^W������F��N
��x4T-,��O���)�k�:�:Y1�q��D��AV�ú0� K�gs��L�je0[�7�h%�Z���}Ü5����fģe�u�x2MWR��5*�	R޾丧;�S:�j0ñ����[Zl���{b��s�)\��{�nwU%�'�%���*mƞӚg���ڱ[��v`z���A2#}=;�9d�*�����Hs�ۃ�a=[���N%P+��,>��u	`WIbs5�S��áaA�ڨ%�g|�����ל�8s?�Y�%�;�=H��������]�<��t ��r���Q�ǓB��4i� Lh��j/���?s�Uj�m���{�Ww����V������OQ���
jL'�E�j.�3�d�Ւv��:��.=�%��~�ӗ���}x�ө{_7(�=y���؛��s���ܱ�W:����ѻ��J�/ b�{/t)�]Y�M��߿����o0��ovv�S���4�x$j�b����qڸ:k�Ww�ʹ��ym3�L����eU��,No�C5�^Ґb�NK8�k�"m���9���*�2�t�{�
�:}e_u�ر�ٷ�t�uN��k��kd�I���,%{�����>6�c���\8�A���+��s�7-���R4�h0@�P���_����5���Y�)몙�Rud�n���N]f�[ު�A��d���~�Q�y
�0��9Efz���L�ע�3�U�[w,s��2���N��Uܺ���X���jx
��"��)6�m�4��^A��Ύ���<9Uw&E �*A[��+U�xoì���X:/z�-�6�5
�A�so�{��#���>ǻ5�A��%�^կu7==�UΌ�n��|As���`�Ι�ؑG���q<o#��D9dK������0������0��/{�����O	w�Y��L[oF��(C�Ty�O����r{��U[1����#�t���B�l�R�w#�]��WWS���Kǧ��wVde�v?�|�X��m��Ny�]��5Z�ܢ��H��o���xd��~+V�w�����������}
w]x�K���uFK�]�N���j����𺫕L��!�k�P�dF�
Sӱ�b��V��.j��a8��rl�h�@��AOx�F��G������P��J�`n�Wo�"�X�0��{��sU@�Z�Ũ�e�=��gq���X�ս�\�����`vI&�����,_����jA�	:���,q�FH|���<1�f+��$�\���t��M.�uoFwR>]�Vx��Z�yeOv̜!m�wNs�q���;>���
�|��J�-��^!W��8J�0�jSw���Xl���j���~�e����=T��Z748�nx�b��fGVS�^4\Et��m��<<�l@4qb=�_'���.����ve�^�����@Z�N��<��4����t+�9�%U�E�"B�e�.�M����n� ����sp�S� �՜�;�+wb��{%s֛���<g&���W͹B���`���>�߬����α���,2�=�a���V� ����\}^�u6=`2"Y><^�������|>�ѳw+�c��Dw���\l�.�ܺC���/��r����L�ΟBQ�]{y̚�f����w��[��7����r��{����Hm�{�7��5t��g>�xb��O��o�����Fg�o��\�ۓ��G��-��3p�MwYQ�x�m�𼜐�4��^�'�q��.��7�T%�1)嚊w�ͻ��T��n$�+K����dy������hD.�B%�Q�b��;��G*"�:@]|d0d�zkg^��NS���冸`�,m��|\\)�o�I#m�7Uw�g�dwN���(���1�[ с���AH*P˞͉���'��{n����Ǆ�����w��)�;�#�2x"��ͽ䴁M���n���-���玾�@J
|�J�2��ok��t�L�n�����]nyC8�ȇ��R���X1����� m�C��f��Ȉ�PĳH�eʸ�p^^`��\[��%�Dmhߧ�׏�7�Q���zIn�욏�g��B���UGz��������/,������t��Q"\�d��s�����͘�9�ќO�Y<�u�2D5�8����V\��`F#g;5+s�Vjo{�ַ�����丒���SRY�6=��CZu�%E�VU�iH
�{�v�}BCͮ��{�
#�(��t��U�[^f&��n��.QoQ{���E�ң�I0�4�{jLS���5�!�w(��)�Saj�,1mC�AIʖ.1��]{�:U6ה�%�ah��a���L
W,�.7��|xK��%\�*����VWq��P�n{n�TӮ��b�Q}�9p�n�A�O��!���l9�C�����i���>K�H�h�r�:3��Y����/U2��x���fG/Wy@�EE��V�蘨���2�1x��nJV�3f+o;�l�k�[A§�T�
=�ԖՈ5��n��j5������%Eu�3ݛ�	�3���o�:�Gk�n�27�K)##^GEk���4�x����ӗ���{԰�z�O�xx����"��iU�vU�37u1����.�J0�1!^tHKvB�2?h/R^��n����o�'��/������]OL�_v�:�#��J|�㋲�K3��f]~&,@�w��H`���TK�r[��k��;|4w+y�b����އ)�W�V����s� ��*%�.��|�a���4(�ö�Uh����~ 	U*߇s�o4��7��b~�6>|Oq��*��s3r�zFU!.2��kU��s3��{�'�!�<�{$@ˁFT������eN�.j�4�<Ě���u�������-pۉT��4� +2�c��{���òmH:�Rk��[tr%�^B,�Y{'�ga"�Nq�FB=���������ttC�Z>��nT�y�-�2��݄�=�s�iI�eHdS���]��8Bձ���(�i�����[1N�������Z���Pfo`�׾sŠVR��Ndd�WLǌ52��:Ŷ���H.��T��F�㦩�.��qSݾ�X�3o�6XS�	�;�^��FFCfCX��X�=��fr�僫º}�@���4����4�a�s&}ܣ2n�W
��:�P��]	F�=���b�*�}�lm2�]�(����v5B J�*��������T�9@��@��.9��V�<�>��8o��׊��l>V̜�3�z�ؕ['v�=ݪ:�Uʩ�ucw��?U���K��N̦ɜ�ˮ{)/F�˼�RuC_~���ۑ�Z(�7X��ꮮ�i�SNW+�:v8��U���(�Є�%dx��KX�xfc]._̀X9h���o�M���{���8{V:V��UF�9��D)dF�spU��K��SWr~/���ޗMmξPh�e���H��Z�(A�{��ty�,�������� �7��rw��(�F�ø���C�f{3���z�|q�X���n��#Sղ��W�Rr�e���-��}�KB��ô��<(_A�Ef�f(�#��y���n�dT�qe��Æ�8����z�4,��0n������8qg:q����0�Suu��>�{Y{�n�~��g�*���\X
t�������� ���m�[�:e�_f����n��4:��Jd1]W�������؊����uK��N̔������s��y�0����=����-��.��+�ٓA�*,�O����Y�JCH��̗�3}�[D�F	ϧ�Ur�ǆ��k��i-����n���<y�F�D�}������x�,��4K�v.N���3�-�;!5e�:qޚ�Ѯ�<��t�V�J�Jg-���:AR��;��X�;��EM�il:��xn�b�h(b\�w!ܒ�"��-	�r�!dw�*�LT��<?�����懿��w<���vz.�]����C�WS
��fH�⇅HX��Г��{d����U��k���o���4�y��bn�6Q��� Pw��}۲�-ҽw�}� ����,�X�\�巽�����|���6�}ɚ�����S�#�\�;}۩mwQ����{ӓg�+�x�p/�h��b����Y����M]�K�h�Z*,VЫ�#��lP��=���yy#ؙ7�e�Iy���e��>�?n�M�t���n���v�}.K�FPݢ�N��L�5��V�<�X�֒>��qC����1�8�5���o/�`�o��]�z�]8U^3{��GF��eY�֦/5���ƞ�h�2�g��g�ϻh]v#�=[<��м|�\��Dn�Tn�R�ZK8V���Qv�L�-9���:9%=3�+<��������.w��K�mh����`���Fi8��MyJ�\�d�{Q�S���Jbk�n�/7}�)�Lqh�ηW`�k'Q�et�TJ���u'O���(N2�K�<�0L���;���g/L}�b>�;�7{��5tKo;:�9,�[�ws<�K�X9B�4��ϯ��t����e]ӗwh�zM���Z8�$q���eW���(�>�򖪄�Z�Q��Q��%�:��ǎ����q�x�ׯ_��v����͹͸S��}+���^�ZITB! H����ׯ�\q�q�^�}}c�N�<��.��Ȓ,a#P|�ĄK��T+n�___]���8�^�z���N�4yt�$�r���^�.k��)�y������wZ���U�˕�;����O8��u�E�]�zX�9w#���ů����{ޤ���h4��t����sW���\�Nk��r���|IG���/�.��]|����+�����j���h�˗qnW.�mݿk��z���oh��$[�'rI��N�ܸ�{��N��9w:����o]�Q��2���[�t�I#�q���sO����
�dxz�kZ�q�e��O>��>�}��؆+)�L�N}γ�Qv�L�<F��i�P�-���=���|=��.j��)�����e"*]~��*[i���ڞ���_���v�Kl[_��'��;է����q�/��Vv�����{K��<�[���sř��c��1��[o�2#m#6-/_(�}��L��ulu�kWF���^vh,�*��OC\7�ֹ}��#o�(���O]0҅BfؕopW0�]Sty���F8��E	�����a�â|��b7$B���5D����m:ٝb6��V����a*��[���}����i��az<�����W�a�JfV��;dq}����&��`�`��||��8��A�9��q�4e��ک@w�(e�|Y�g��Z������e������1ĝ��q�v㿿g'vg!�K�����tH�jI�d�"L�9w�Nk�;��]��-c��bz-�ҫں1{�.C50��+�s��!+˳Zlns���8��7��Dվ����;�h�@>t��&+sw�/�|��mG˥��u���p��5��/e�J���w:��ք��+D�[��7��\��n�~�3u�wy�Ne��W����;�|���p���dc��c�vaJ���d�g���mn �f��nw�|Ʈi�m�d�k|�WGz�j��Qh���GW-:�qv��w7u��KH�mY��]�X҉�\J��
Ѷ�?4�T{q�r=��+�9ə�zi����������Bޔn�/R���R���v�2d�M��q܁��I�m�8���܈tUS��k
~�cK{>�]�^ast���� G*�,
/���7��g=����ٹ�y�/z�}�x��U}�q��ϰ����p(��ݓڣ��b��Ľl��0��Yk��,1�O Gn��(�ɺq��m�xj���g3��l#���D�Z\��=�̘^�k�2v���e��Q�f����w�+���u��vx�z���D{�u\{pg�ݠ�w{6�j�纜7����T3�^�ViX΅�g�.[ۧ��N[���	�,ޣ�c��ˀ@q����v=Z�!�
$�:C(�5��5	^U�7.UUN}�z�#�j<���ϡ��7Nm��y�bЃ���8k��n�?{||����_�p��s���������e���~�p{]��.�/8g�W���"�r����l��(������-�����0חm��z��Ɯ�n��ƍ޺f�mM�ur݄��#.<��'zF�N�}�����; L�\�q�pg����c��$5�g!t>\�Љ`ɽ�$S��F�&I��ݖ�v�t�L����2�|�6���N�]鉊U�V.vc�w�ix�F��+�`�p�t���-~��\�7�л�x��8]�r���gtC�ƨr�e�nh��/u=��ϴ։��q�ղ��Ϟ�,��0�k�=�9�{^&�_so��.�C��͓�D"
�����R3G�T�湞ɇ�vh;{y6R�� o Fly�:�f��C��q��gB�w+����<=�zÚ�tys�E�w�S� R�[�����{����>W�]�3�1ܑ�79��އ���v�n�r�@L�s{��s�h�J����⊶U���ve�m��Y�.�z-�0�}r�
2i�.�y�L	�ǉۋږ:�ЧI�c��i���jZ}�)�˭��}���6�O</�����LωC_K��4��rʫT�0��:ZMԷ�����.0tjނ��9;�x�6��� �0��y�F���1�p/>Jt���ۂ����p���PB�v�����x��c*2���h�QOR�X����`��&�2m�a���W�3�b:*�9�}>�l�g���=���i}�#1����Macf���w0:�|�P��i�<d�Q�W�%-��>ΑœdPw]2�V�T� T
p���E)��LGG�0򴧗^x���_��]SS]a��U�We�{�E���ţ�h{���M����b�q�S�ɧ�j�M��u�]�Q'*:uY��~ֻ��C�c�p�.�Y8�T��mi��~y���b��,�&�2u _�|�9 ��u蹠ϋ��8&���X짋t���R'��s���w=��)	![bVKP�=����yឌ	�Z㓁�/*���L6��<�������d�5��;�}�7�e��M�ZXF�X�j��a�Y/t�ma�o����3k<A�|Պ���U{q9�o�[��b�-��m��W?g-b+2BY
Gq�����HYrnv#V�6{o�VߏƷ{�0@������u��*���޿ �
I���M^�K�t��4"���0��Sa
|x
�X�C�ʝ3��5Y���dl��T:��z��Gj��{��p�IR��v��N^j���|vĺ��?p,E�t`u�Uϟ�N0U�י�/n�wvr�Wr��䪣n���=m^A??S�0��Qu�5GNἶ2-��K�r��ہ�~Ӑ���M�3y4�nun��|�a�3�/���uʼ�*J�FN5ۣK�SVR�A��ݲ3{h���wm �uO�EP4������2�K�c�D��&�e�p�n��B��p��T�@�>��m��z���st:���_�\Vv�zݜe���a�K��W�����������G�ۇ�-��n���H
�� �8��3(��W��z9���
}v]9�O0�,^J�q����ʎ��{),bd��<���1��� >o94������4x]��O���_����EM,�s�ku.�q���{n7���~��c�g��bֽϨ..�c�1��3�#Zޫ���矈��y��P�Ǭ#J�����կ�䉥 [Y;M��o��D�H�Wb[/�s�O�\�:w�����*�[)X��C%/þ�G��:��c���O�T=_��l�:�gtط]>T�6
I�t�?i�5�{|J/{�^��8ѱ����/5��=WO����h�2����!=V �6��e��s�N���U�&��D��S��u�H��Go�M��}����t��qx"��O����Qf��\
�5�V�Pc��^ڲ��e�ݙģB�ƃ�yHH�-���Gջ�x�oc�k(͉�y�v��:����=ּ��!]j�FUKǨr̕4�&�63��sS�������r8�릳Ɔ��;�K��V�`s��[Q2�o�nMo�7���,l0`\���M��w�ަ����q� �o�̅����C��3ey�0��ӕ/�3/v��v\˕T����v����uR�z�"��k{��,�{���np��x�_mZ5�ɵS=�wтzt(�DO{���A��͎m�n�2	wGD��M��yW���a"[P�]w�e�3���<x�=�)��������������������j�?w7�ǽ��z�kV�w�+\}�~��]����%�R݌�Cg.�5�'�)���X�Ij�y9z�i����*Vx֜�1��}���x�0�2�r�#�2v�1�-��7]�gD�Wwq&ָ��%�y����dd^+"n!=�s/+�T����%�_o?vi�����y�)���oN3>��#��q��{K���
&������A�j�6_Z�6u*�U�H�a��������CTd��q�Rqx�w���u��W���5���HkpUA���]�j�(372F8Q����U�o�@�2NX�[��1ہ��R���"�Xf7��Y��?�8l�"�Õ���%~��$�!&2EAy|��v�p��=v�ݪg��ќ�d��3�1�����D�:���y}v�@�R�۳1m\��__�����\7#7Ru8�%�1�އ���.>%;X�D*3ԞD�S��>I��)i�a�Q�S1Õf�7ch�]C0]s�l�41޾�����z��L�19�V K���eHz��yrCA	�	�X�UfN�?�v1�b����L/�/�R���.��ŕI-�����.��j������T�E�ٽ��|.قMo]n+�[u_�WzWmv7�Oq��q�,5gQŗآ���Jf��WP:������gC�2ٟ�P�ծ�)�����"ˮ]��Z��_�}
�[@��W>��h�F�y�e����M�]W[f�����KiPu"�����)��^q���9Z��uc.TK-���������=���{��d&������qe��;�u}ϭ �nY=��A��mԣ{g�@�v�q#��{h#QZ���`�"���\�=Ù�T���ߤ��[��� �[ԛ�2�V��n�[8�>Wvٹ���Lt��+�.It��
���K��z��������C�h�t"|�'�_k�-�����(��� �Wf�+�����8�WN}�M��
�n�"0er�%������e��օ�DV(u�x�`�DO�N�A>��W� hW�@"E\��n������x�2T����j���a�)���Ik囃W1��}x�Kw:]�dZAr��'��`�<||������N���Pb7&���_��L��j6Cdf��h����1��蕝���9��8ߟ�j%P/>�$ӷ�b�������}��Q�`�$�JM�z��%�f�fX���t�Ԥ�����*s}n��.�1���\#v/w�C�@���w&M+ܪ����gǐ�E��Bf�<X����=�ws��[MwZ�n���A��{��1=鬎SXB������V����˭���S��a�u��*�ߞ��b3V�]ז"�3�ԭ|ڧ]xU������xu^E�?��P�с���²���g�,��/h1 �yj�\��;d�U�V�4�Ϝpw�U;�>�i)�å*�ud�go3u!Ҳ����ԗ �w.����\<�=�^��L�̌����%��ĭ@>CdVw^^kz;��uʛe��w��Ai��/��>�l9�m��蓹;{лt�Ή��\�E�#�PZ�,���5��:�zK�'��m�c���W��wIb���n=��9S�E��m�n�I�u���;���5�.y��Փ�D�M�<�wG"k�3!�O������y��E%3�*�?{���G������)���Y=@�������;ƞ�-}z��yB�{F���G��@��Fm���Vr�V�ʼŉ�h�˳���Y�_����v���DG��κ��'h�[3J��v죙�C�*�7k{�ӝ}�j�e���\^Gv�2� �ڞ5�ܩ�=$�m����d�6��}S\�&��TDNF]������󍾪Q�ݵ�eRKR8�G��Z�2��^��X�T��u��5z;܆��!�m��.��?��������_��@�����ި��ӳu�o�� 0��|�U�Y�yOp����,T�<����'�!��ߴ"��ˍ�zs#/��pQ�.��t���H{J��WWJ�Ve�Aớۧ4�1�]-T���{�Z�G�����v��� U�� ��_��� ��PAR����E�QѺ��c0BR��Mk2Y���������ki�&V�c5T�f֘����Ե�e��fc*ٓ��1�����Ԫ�J����SmM���R�jm���MJ���MKjjZ�,�MM�mf�55SSj���ԵMMjj}6��5SSj��������MMjj[SSm����Z����j�������mMKTԵMJ��j���ԵMKTԵM�ڦ�jj[SR�56�Զ���5*�SU55i�����MMjjj�SZ��i�V����[MMjmejjj�R�5-SRښ����SSj�����M�֦��5-SSZ��ZjV��ښ�i��(o{<�(�	��B6���55��j���Զ���jj�k5���ih�"�P�A�D0!6ںԫU-M��jU����T�+U]���j���U-M�T�5j���U-M�T�+j��mU-KXD@�-DE	jZ�KSmU-M��Z�j�bʭRԶ����T�6�Wv��R֪Z��RԫU-J�R���KR�T�Y�����T�-�T��w`��
�(Y�KR�,�,�Jŕ�����R��������ڻf1�Zd�kL�[Y��K)�ZX�m2YZ�J��f�5-[�����6�śjjZ���X�Vc��1��jV��Uf�V�ֹek1���K6�b�jYlͶ��Z�YU�3Z�K6�jm������V�����P$T#@R1?��^����s����N������:����h~��O������a�r��*���������?�T U��?W����""��ǩ_��C��4~������}��� ���������i�?�8��@�;�������I������
�P�D"A"�MM*Ҭ�Kl֥����jm�����U5��V�e�-�Բ�6�T��+5SKT�Z��KTkS-TkQ��j�����U!"��H �2��� (���U���Ȣ&�T��Tm���j�kU%Z��Z�����)[M�Ԧ֚Z�mSeZSZ�[SSZ�f�5-STե��f�5MT�-�Y�Jj�i�MRڔ�M�Z�f�-*ҳj���+*��j��i�kR�j��KR�-M�*�Ԭ֥DB �CV~�������Y�'��
2
*$��2 �H	>��+������@������@������?��y|�x����}0��Κ>��T U�����a�Ͻ;_����!�p�!�Ԋ��/�`��}�*�?��J��t6����x}�£��X� �?�������~
���O���������a���~!��}O����a��W��?_�@_�h<?n��H��|�ҏ�	A��z������=N�"s�Ҩ ��ܐ�<?bR� �������=_��(���
�[4��"����������)؟�����)��Dd!���,�8(���1!��p�%�V��,�S!�&���KZ�U�������eU��$kM�l���lʋY�mjjMcZ�Mb�4hm653�	$�66�F�j�e��`�F���%�h�DV��5&��Ҵ��͐�Sb�m�mm�l��ݓJɫSm&�[elh�iS#٪�3��lY�-[XU�[7��m�%�f�ث`[m�V�i��-�f+F��Zl�4j�V)��ʹ�ɒ���֙Z�El�m�J��l���0�Q�J�j��j��ƅ	i��   6u�۾�p��޼��E[m��gnڕA[G�]�o5��w�'ev�.kݻ����t�.��CgM[��z��{¦���w����y���^�������n��֧Mv�i �ĶX�A�����|    �Ǒ�>��M��(]ϵާX�)^��D��y�*��^�bE�]뙻p\��W������t�nW]����v��ڥ�M�k��ݦ���=v�6OU^��ZiR�v��u�Ô�{[��V���j�-���[j��   o���}��]ym�p�Z�e]���wlٗMZ����J\�wH���[n�m70�����t�ަ��m����]����گv��:^�5�����ڒ�۹�����-f��ʣ&H>   �z�Uko���]P�S*�X�]nWnV�m���s�H�unmî��n�����]�wR���x9ڪ�U����4� 'Xm���J(��T���  {Z��ަ��iU�up+���n�5Z�k[�NK�]Ҭ��]={���ͺ��i����u]Sq`vwZ���mZ��]QWlhśS@b�ե>  g�[e�W�n�wwX��:�[�j�lA���������k5������[�q�F�,�V�ZҔ3]���W��C�TUO,�&ƕ�S`�cS� ��Ҁ#�+���g�o�@PoC� �(�Ǽ�:Gw�n���]��r��3�G���AР{ڼzh =6�i��V�����ʦ�H��  |�B}�����(���憔.{����O[*w( �zv�� ^�����Y5���' A�U�@�M�H��K���Q6�J�m�e�*���  u�ACF��^ t=�y��K�^�  3v��A�v.��B���� ���{΀�vu�p�ւ���N= q崌&�m��S,�!lQ�  �>� �{\��i���p҇[�G:P +yz�l�������E�L{ 
������k�C���kn4 u�M�2R��H�)�FIJR�  S�b��   �~�R�   Oz�UP����I*�� 4��~���#��3�����۟Ջc�5�������)�El��8tV�LP�_���}�}_W�}���鵵�m�5Z����������������Z�ֶͶ��m}���g�y��h��@)@�[�f�bƍ9�m6 E�ې��
#wh��aIτ{�^a"jɔ�0���9{�IهC��Gu��#�� ��fM1�V(�[6� ���v�: |Iɪ�L���6�
Y��Uٸ�� 9yW���S���-����&��e^���d���)�[N���Q��QƲ�ô,툆�� �2Z�MVQת�<ʁCZ�EӃ`�e��L@�K�ɐ��5������r�z��9M!ô.�v�S�Z18�c���E�
��	8���FArfmDٕv���W5�@����]�;��ݽ�ic�	���F�=�D��R�n
��CY�X$���>�����%��3{v��kK`b�hcT6T�Ų�y���J�8*��DVӔ��(�$Am3h�jR��ݥ�hb8�S%df�ڑ<�m�p�132�02}1$�C5"fU�`#���_�i�H���,m*6nc��M�>�!{��GB���ɍ�^g�V���h²�Rk*���z+,
)�Y�b[���"h�`��i���j"["�c,�T��-7F��&�'4�XD|��ed��*,�[�!�q+	���1�b�=6옓�԰j�:i]���kf�LC@�41�
V�9��R�А����Јś!�ƹ��-�7nD����R�;��RJe�U6��2c	S ���3A����fX5d��p҉�[a��~B��u��y�*�)�w�{��-飢��& D�'4���I)���y@m(��R,Q�ݺ�2V��� �[�����q�4sJ܉^�*i�4��im3`��ڧnF��xS��&^TT��ڎ(zS�g�m�uY��E���:��^ě�S9(�vu6�ͬ���.5R0jѨ�M�W����c��n@k "1Vr�f��`���.�л�44K���b�j�P�s5�6�����SAl�Ǹ� ��YR]]�YcF(�A��H����WZ4`E[WN����b���ؖ�q"�������b2]��-"Ƚ�d�#�[ ��Zs�G3Me��8%Ѧ�ٶZ��}���P������d�����x�)��@��r�^�hr��K5�)"p����7�] �4*��њ�OQ	[�&�a$�%�PW�2bkk�̹�ԻA�t�D��C�,�
��ӡ��f�E�:�㥿&�B�]���Q���8��V��g>W���u�)Պ��r+օ��p)z�j�a�{�2mE��R1N�����X-�y{�j��lmc�#˰eFm����
�i{>R�dZl��k-֋T	���$�����l��A��S� jP����A�c��Xz
l�і�D�W�p�;�C�m�����u��Y��B���a���� �F���"q���CV�,e�&d�w�3d��e�K�t�@�f1�ֆ]��C	���BOMn�p�{ ��҈�Ohd�r&�푊�+I��4JeL-�vMi��tصaa�/���i�-�Z��6ҩNY%�a�U��������e�Z���e�"Z��'m����E�%;SYØsA�������u��z�.��x�nf�ۤ��!R��1�E�z�{�0���éQ8U�� [f�"� � ���G�h�@K��mXz)SEӬn��M���M����n�FQ����]+<����C�k�iP�JF�=��eI�'�'��}���eDR��|.V�X�\5�*:JR����H�!�#Or;��u."Ķdb��hV�35�L8E+��7�����=��fnFRm�2a.�k_
-j��˓*��D+��d5�Sʛ�!Vf!Wq�-�Z�y��3p2\�A�n�$��L7��ZQJ�`W���妦 T��^ݳ,f-���X��֜ ���o"
:�V*���Ԥж��^��	�r�卍�x8���H�Up�V�-1��ԑek�����G#Mޫz΋	�e�B��ؽq�ݩC]�Y��h^L�����nU������ɴ�AhB,��twHNZ�D����/v��ۦ��W-��dł�kf�BΜl�[SD�<kb��`{��e�ұo�V�54�la�E��S0��Ƨ��u�����RZsTXԡ,&��^	��t��;D���b�q�!�V�Tޝ��Ё���v�'o^cVȐɶ-�X��O@`�$l�0�b�8h� k��c(k��:��k1��n���ɴ�hc�\��v�$FJ�!���hJ4)�%X���j��̍���b��oݦn���Pjj��rVB��,@t�-e]`�v��[�@��e5y6<�76��#�X-�R�0�ʙyR��{�/a��Ԇ�ee,ҩ��LTJ�Ko6e�׉טA�@�G�aOu�� �A��o.����-���fX`�4�+ʼw�
�8���f��Gp�f�̖�[�MJ��!�4K'5�G�r��B���R�ClhQ��5��V����8�;�8)H$@���Vd�F��f��b�$e�6 ������'H�6��X�@�1�3j��0i�L3�p�~u�j��r�:-J�ئ\d��4���ESX18��n�^5Id�h���Mn�h��n�[2��u�B�%<,�-$��އV6}��ƫ5��I���'���a�Y��ɗ���%Zvn�{��41��6U��8���%�wx+"vn����/R �VU�z��]:v�;f,�v�m��EbsR��І��C��I�y�nb퀩Y(1e���Qq��m�ܹA@��Q��=��jA�6�ˍ����`��0P��rTYGv����B�̱t휷���Ҹ�,F>��p��2��!V�"�O�%�0^ڬ"�n�O4�5�1&�j[u�������ǀ\W7^[�X�X�*4"L^��BTT(VQ�=Zp�y5(Qb�	M�Q��V��2�-��j˼�����i��E�[h:M�!�d���0f�;7D=U ��j��Rf��Boj	/C�Ѭe����T�E���#nϵq��%�K����˭���ǁMV��(`�t ��	��SCn\{0�aƋ�윗��ѨH�Z�W�]�E9s4��$.��iј�l2Z@Z/絮[�ow�1���D�M �I�&�&en^�W����MѠ��u�oN-��%;ur���vj��ةR��?"�3���-�E=B�
veͣqd�j��ち�X��wj\�_ס6��f�֛��6(���-�ֳ+AsN��x�-���)�@�H�X%L���-�)�*]�V`0���=T�֌4S��.�t&Q(2](ɤpbk)�"�nш-�.<2��&*���#xo�Cn����.�I�ӳd��(;�����y-]�`�7�}.�v,<f��ɍ��w��O*h�Xn�,el�L�&�H)n����Enn����r�+�sbDE]!�����"�pU��)�	����L iʂ�9!�?]X�Q��Ṅԗ&�4�����41�偮��q��^�r�2&n�-�8��Us$j ��g$&5vnĄ�t�d̋pm�B�
)b�)9��]c�O0T��+"�lښ��,�<N�uh�� ��`�jIW���#zL�P�Mk(�F,Ųùp�f<T�:�Kra%�Ь<�,��0�U�g���]C++L�6Y�4d�ܺ!ѡ��F��	w�n˙�-T2�5��
�A�<���aMB�=��6i:�.��CV��ZU�����d�6L�;m�iŲJ�Z�MZd�$:2����s���q��d<M7v��լ�1��gKd*wYF����E�0�Fi�9DbN�!}���r1d��{n&��1VO�^l�iQ��5VK�e:��i�N�6��
�z��yQ�5�C���4a�d�R�r��3uChY�%n  :�%Jޕw�MĘ�d͆���m�t�	Z
vLZ2LzԻ,5B�EvnKr�4���ww0�I�SN���"m�-:�n���[�ҩ䖦A��2lth^�f�Zғ���~WGF���c,�CSE2t[����dd�l��]�m,�B�&�"�$�R�Ԣ �ۢ�ˣ/b���1,�i�:kr���E�1`�LI��C5�:�*ӅŴCxY��
ڂ��� �SK;�4��)���)�;v�d7	�gn^�k���'(YoF�A7��"̬1���v̹���p-���M[�zU�I�F@F��(���D5&��}� ��V�2j�S����*&΍�r�%#�S�Bj�t��`L�B�%먅=ӂ8���B��{$f�H�G(F#8����{��uP,%)��l�Ą7sB"����(CxUa�Sv�\4��/.�	�����v��fc�M��f�V�LRE������e� i�.J�qY�b�K͠K9
7`e��zY�bz��Ev>	a4�o@�YHͬ;
T�َ�.0Z/M9y��;���VR1��$fB�銅�`[%��a��0�)��6�1�����q��Z˚CߊZf^^9!�sp��v-+qn:Pǚp"�qʍ�� �[o0!
͑���D�Zr2s�)��+v�����P�Z5�ڸ��,a�/0ʂJR� ��мY
CM,Z�V����6�wwȭ�˸h-6��,�IX�[y#��C����"�bEJ1�<��L�]
���
cp�F�L��@h�0�Ak�P·�A`0JT1Rؾ԰kMd3V\����0][n�S����T�F%e;��#,�˨�AW��.��'Oٲ�҈1��
�&ܭ�wC��4���GU{��Ty�ۄF�|Uf�������SBRڶ�$&��T�E`õk{lT�-Ri֑Z�`�ݔpfmV��ha��h���6iϮ�D�i��*`Ưq���F��!�>2ȭ��̶��b3�X��x@���a�#�,�!L�6�$�
f�m9�%4���6�H �u�"�=Th�`��t�J��9z�X��׊��̼@�*\�6�Jy�X9����n�i���Z�7@V5��I�U��u�Xf�7P
�$���r���`����*��`x���	�U����[gb�e��v0���t0��!*
����r��Y U{�݆��թ.��+tYxd�H�У+���Qk�^Q�ŗ/5��b5���|`4f7x�&7ce�Ec���4E�j�t\ �������k�&�ܬ�H[@AR2� $�WeI{v@EqX�.=5�
YG"��:,���9H�	�j�!�u&�sf���m�׷�Z�')̸�e<ְ�ʚX���Gf��Mhĝ���*�L�4-�,��+��~Z��e�Ԉs?��%-q��+��Z�(e�w^\M�jжe�Ѫ��q�3�u�Pq^!��|pR����ŵ�!�n���P�/�����bZeG��)\�-ɢ��;b�bX6Z�qT�hAE]I���{�AZ0頍��Ơ�**�f��f�q����2+f=���a��YD����?#H&A�V)5N5+	ϥGR�zd�kB[{��hSF��%��5��U�8V�ݧk+K�9��Њ�i0˗i��y�K�GWG�F�ōҪ7E��n^X�vsN۱B�����rc�be�&��3&�a��f�VmƄV�є�Y:�@�nBl��3ײ���;&�2�:1��J�5���&�,&��o��������W���c�wh�~��r���D�I�`�D�!!$1l% 6�nԫ��NX�$""f��V���Ȱ��Srf	v��b�T��K�bנ�`m�Y$�s઱ԸM���0Dj�Z�V�X�v`�3jX;-��%cʅnۼ�R�C&�_ZfTea�:4Aq\VMnmb�M��	�Lٻ����u#�R�����f[�U0ue	E�,C�$c ��xܨ����4�2�m,aw�,Nl��w�-֣��m�����dLwp�WX�k�eb��AL�A$X�l��[�=�Si隤��[�є�d�o�.�%�9N�bH�8�b5$ǒ'[��b��æ��4F��M)-
bt2 ��!GB%�u�H̱��LV�M:ߕυ���	 8&����5j�i"Qa�z�;Z���7Ri#v]��o�Z�p<��ðS�K���v������
�k�&*Zǆ�!qڏd�=�OZ˟i_$YǛsqP	���y��-�KS%��:B�6��*�U��G��� Q��ֵ�[�Q.+8$ǌ7Wn˻�l�R�uy�ܧ̀i#[|���'�iy$��6�`e�E�����E�D�#�����,�x����Z�]``�kƖŮ�\4d�D�F��� I�+N�mZ�7�l�|bxM��Υy�޲bd�����Lf@�
�s	�$��J��$�%m��`T��%+��kL��)�_�jL0	wN&u�m:��i�UaZ�*j��l����lP[{�R��Eڛ%TYt�
=�
��
̓J;&�F*���꧹�K�D��G����y��h�է`�Q�x��/C�(���'(*�XF�I�,��ɛ�AI#ǧu��-��r�G!�5��T��,��#1��:����*TJ�[��j�^�)�Ė�Y�N��в�j�6�i�jZ��"!Ӵ�Ԇ�2n�wN���:
�/~l��&f��"�pǢ�9B��n��Mk8t�2*^C$B�R���>�Zh�7�Ƨ��1�W���=dd�I:F��z(�v�gњU+4�]�Fmc��,֍e��i��+5VKf�E�8)G>�Ŧٖu�j�f�O��`i�ݩ�/^��Qiя%��Ub*թA��r�v��<�У>�襇�����P[���M�jQ?0*�7�ֶ+N,4�Z�"���؅�N�({�\7���TWmd�}(T
]��{� ���1��j��R&�'��(D���ֹ
\�%�١���|�jZ��6`�ը�NC@���d�[��r����V���w�+$��(+����,!w�"��m>�m��-u�a��L�;� ���#F�Ɩ���@��ή
1�e��[	MD�O�Wt�áq5[�{;�v�-��+d.����ᙳ�{J�.'����'��d��+6�C@0�a�o*�l����JN�5��̭�}'���y��ɬ���/�Ku\{��A�lV��j��o��`���`Ͳ[u���u���v�e��nf����y#��m';-MTo3 4Z�@��,��t�2��U���R��]>b��s�����g[.u�Ȟ��� ��|6�x#��_I/�n�Ϡ���t���1��P�5��9�Sk��7�F{I7�')�hN������룩�����O���B�+��!�w[t]����.1b㛰��co�lԠ�G�R����T�|>��~Th]�V��|�=�}�
�U=+,����sՅ�eup9�J:��T2�b\�:��d�F����Z�C�k��%m7���+0ʜ�T��N�m;����E�0�
Pju�C��V�-.ǋ5o[�N�k�V�d,�f�7�8>��t"��Lu����O��6���m^6`�:�3%��W�3��P=}1���n��*f�8�.,�]���8�ۺ���ᆃc(��yƷ#bS1��ծ��2��+�}�vڙ�x�̦�!��f��#F�(��[y���{d���Qdl߆ԵAEe-8�B�ߝj�L�`��軷��E��0Nf̗�
�+�0�嵖�]��b4w�X��W�����c�{Yt��ݶE��+9�����ӍDg�x��$�� WX�j_���.XEn���nц�k��:�'5�|��l��#&5�T�����A7)�t��yxġ6�d���,+d���W[��*u���[g5��}pY�'dҽƹ�\��=\�=���hIC��+�.0��e)X;b���42C��e_c�Z�rnT{4u�X�7%�Cx�V�p�@������C�c��m7j��ͦ��Wvc���[u��ы�v�%�i�5y�dai��!�r��y4O�L�i�2��ӧ}v1���9!�E��rB����{E�>�!��a�=3T���ܬ�D+r�,e�2F���ku�\~�5�ZC���ض�L��k��[�������܈�75�{.+��tͧY��.�zM�ڒ�h�:뺍N۷QڒRiuq����V�(&9}2sF`�|v3��N�q%��#;�[.#'�ĭ����35���H��yQ��Ԗ���:�� �#��DrЌӇ{l~ι�z��S��)נ�*�2�`�o=�1�����&k��&7�!O\��b���c�}w}�ƅ�[�9��ܥ4�V �\�P��wx۹��V�t�)�Y������x�8&��ɔ��]���磗
�ׇ�W	$�v5ö�e�Ռ�:۲U�)�^#!�k�>+:���Ӄ�e\����'ٔ�uu��x��t5�;�n���=����S&'tܧp�ɬ s��$V�XOts.�^���;��v!��� ��u��5���".GX�:ɮ����t�%��V�łV��R4��5�}��t��ӥw�4�ʎ��;K85T��@܊���{ۍ��r�CJ/T�eq3�`5	�Y����;;�'|qwM�k�FN�W}	�Ꝗy�9+Y�B��ji`�[��p-�B�^��5|�	���*�����W11���5< ֝iaG�f�u䇃�����l$)���7�0�:@��3�wc�:թ���+�����]��{c���Ļ��H���ϡ� ��׋-lⳆ�!��N�u_c�L'b�7ZK�����r�in����5��]��;ܧ.�Q���-㾤�3�uӗ$yC*�N��ږ5�v��t��4&�!�"=b���S��8���X�f�$��%�/jM8(��H	wJsf��X�옹�< a����6�G���J��w�7���u2	:`�v'm�=���E�G]L����;���!�v��!��i�s��T�]���N�]C��_k�dt�Q��4i�ss��R0��7�5��=j�hn�w������1T�dÅ�6 �GfW�����X�����f*��Z'mo�E�vX��*/�±�TT9�f+Շ;�Ym�S3���yV3�|���Ӣm2\��)�Q�<�*=��[�ˌC\u�c�w������;����An����V�L�)�ܫ��D�U��Z{�����)b���Wά't����ܹ(b��r�FԺG?��+q�G҆Be�4n��s=��' ̑����[1 Ui�8t��we�yDS����F�t+�e+�_l�HmEe�8MaKX2���rFޗY�J2��wiB�)�z:��n)�VS
i�BJO$ə'B��v�=/!wd��kNn>��j��Pi���I[�s7���N�4�L��@��D���wE@3�a�ZӖm��nv滷���*]�ϐ \��@��Q7���&�=y\S�|�T7Y���|��hzc�b!��m��*��e r�����n4����u<�q_c��CG���3�r�TӨd<���`Ţ�y��G\o�&w�n_;���oY�c8VY�
˘�ڶaR^���z����Xw򹉌�8�t���c\���'��t��.��ý���@��Ӷ�hZUf�j�u�nu�I͆����U!Ӯ.��+����NݳEewTӂ@(�t�\ �kF�Fm�;t�V (ΰ9�浂=�]�nP�B��|�tłr�i=C��-�KfR=�,Q6ѧ-��J6ۛ�.�d�i��u���ᳯE_˭�M �l���BXq���v�1�]m��f�ϳ2v��f�ђ����7�%ew-՗$��B�u�k�I�f��F��2���4p�o?a�z�i�~���7^aX�D�5�Gs돻�mԠ/&e�ՆoPξ�x⥔�����+�����]G É!�U�"nN4y�Sn��^c�&��<�6�-M&��̺{t�U�x�Y���>��z��
������>kOn4�����4��p��݀}{$�5�-��%kvr�i�BK��3�L�a'�w�J������ H�'����:�w�٣��
�T�
��6��G�V�t�g)KF�O���Be_ w;�Vw�f�� MoՂ�/�he����U�Y��}��i_Q*�.��������&θzV��;��]uX��z�A��ǯ����#j�Z��&�OgI��f���Zw3�Y��ӓWvH�sF�S���q2�q���I�&yh.@��(r��ک�~��#P�o'sh{��j뜭���|�U:2��tD��wn�2�׽�']9s��Ռ�8EV�uI�J]d}���%@L�Y�ĭ�2])�.*�Î8-c��0c����by�%����0�+��}VEsd%�j�6��.�ER&I���Ы�$W�^�>t�������v��"�p��]g;[��+"qh'6�;�]��͠���opD�� 	�ZwMZjk�m�Z��A�>K����|���b�po*�����k�N�Xk��͡�o�v��Yw3..�%���ڣ��[3��/'g>o�Fͽ�\n�P���<��u'vޤ�Yw�0��vr|����iJd�H��,�o����vW�y<���dX�PK5�#:��*��6�P���\9&<�׵`�ۢ)XQ$�R�U}×X�-wvo�s���,��<#��o%��]L������++e����U������!�`s�U����5��jU�8,Y�d�#�"��K�X�` ,0H�t�s�Gz#�6�D9K'4�ά�@2�t��7�飰���6nP�
���r; �1��+2�&v���dm�#����,n��v�MA#��N��4�]q���L[�@d��	}K/�㔸aT.a���N#�顪`��o.��+Xh�KU)��a�VnT�m��K�9\%*w�6W#�Yئ̙7KF�S���5���,���Р���l.ۼ�wwi����n^Kx]L��P<��9r�۴qR�C�ER�r��e0� ok7W�&c��z[�K��MPĎ�^p ��ݬ��P���E�"��.�.[YI���ӱSp�7���V	W6eLH������RI���+�Xv�3�0�9*�|��	D��Zʊ�p��H���+ѻ`gLu��b*Od��Δ��� ����v�s���X��gbEI��Cn�B�erw�4�zV�f��u2�s�L[t�nٵo-^ρT�EV7�+��z��n�T:Gj�1�խ6n�n����"��5�{"����uD3�v���Fmj�G�e���	����D7��IV[yӇ��+D\�m5]�M���2\���R�<�lnm]v M�V���c/���ZbB�o��]{��T��i��Y9T�Q1c�����0ދ���E�<�`6tt���ڙt}���}�w�I��AǗ9n�r�y;��(}�]\���=V-ʾ��s�����q��vpǰ���)��}(|K��SMp�<^Q�'.�³h�z����p����<�v �+����J�]��Y���Ġ��#��9�Fܷ�fN�����qsW�xdQ=�r���}�Q����n-qȽ��u!xF��QEc�p�E�U��ʂ3Xz&�9:˂l��h�Ӄ{AἏ9�Jf։��4;�6��_aTƽ��j�TU��,��6
�>�-�D=S�F! ah�1��x��i Eܡ��V`b�%�gW�u��vS�X����̫_S��ϟh8��Â�A9��u�8.���M���qJ�ι���W;�M�+m͇���.��mr�چ�U�>f���S���e�r��h�%�p��Ñ�p��fdr�%G_:�!�^'*�3 %�B0ޭe����҃�v:9�5���o`rv�n"hu[B9[L�`F�bK��e�ǘ*.�{϶�ū֮hM Ǯ�L���ssf!!���\�R���o����ђ���{D��咋��H\�x�-��u�:�E]��S�ڍ:y����&:�f�J�:�C{B�_fJY�.�lm���w��|ٺ��Id�m�+��_l���0�(q҆]��6H[��y��EGRi?�Z�`+�t��	4�U����#����V�GԇK4K�l�j-})D�9����oQ���g�M��j��haܨƣ�1	�1N|�b��YÅt�\�Lo呺;rP-!Yc

͘l�]�La�Qe�u�%���2��#4^��q�^���7�a@:��&�}������V��䴕q�*��Q�����B�.)F�r�இSS6�P46��f��C^�F;���%�}|2.��j�q`�"�f�J��w07�p4H�0�˲:N��B�4�ʹ6����a޸��-��J�����YW1�J���5��r @F_\b�6��@Ó�W[H�wIŢ��u��X��XfL�ھ��沺<�Y5I�WIw7۴�tY�]�Eɨkɵ�̔!�W��38gI�ɔ�6}����m��_p���AQ��Z-�ST��¶#@,����,j:�de�G��nR�X�O ��$Ҋ��o��@94��*Y�
Z9Z�y6�]����s
ۅp��K�F�j�Ѩt�ݙKC]�c�-���>��Z�����Q��]�1u!rK����9�U����y��k��Ϭ�srpx
K�^J$�o�d�3i��q齝V[�]�8D�[�-�[R��q�^X�ԳZ�Y�i�����^ܲVX[�� �p���ʶ����dV#m�,��a�Zۉ\�(�Z��@b�7��o���WFL��{�ht����V�tc����'u�&+]�Xz�C�8ɠ�@6���ZyR������1�I;����	�
�Be���U��gi��0�5�T�7�,��!-S��)t�ǤH@Wt��2Ƣ'fK	��h���~�ϑ�E�J�:7H���ÒO��%�>K�m�����N�Nf�q����"ӭ:�]���E
_�f%tE�㩦��7*c�yN��'�{�-��o�bt�qnū�����%���:�ۂ"��
�l\�X� �q3k���2d��K�{G5��Z�Ĕ��dIu��T���g>�jQFØBx&��,n�JJ�%�aޖ��@ƀx����9��n�8�U�ޞ���$�x�{+x���}:b}-b�\����̩FRԳ�_(����45W��;�i�GM�}�F�ԥ�nL1�tc,�\V�昺�J(:�R5�Z���\��;�Y�S��]�'-��&um�캵���S��@�D;`�@�:�l�QV��[yٶM��ȸv٭u1�F��%�:��ѬϢ��ESg������4/㣫DME�knW̮��֙��W���$v *�0�m�(�u!&L��Ԇ�#{{�˴0�����	]rO��_'\I��^n<|MX2�[2��#
�Dc���]��[}���˟J��k�j"E�u�t��ș�wm�l���w"f�	r�f�{��`�N�t�wP�c�|�fwFV��BNOf����yEĨB�E��3^�s)$xS���:�'{z���F�h��*Jrcm�3Jm����
��\��3)w-�*kiO��7+5�j��<D�V�a���ܾT�ZOq)[}]HtD��,I�]S��8�7V3��3:��)���L��N��.��
��rL�]�t}������w��[�zw�;!چ�]��$�d�w�����$�'�5`��,s�n^�$�&+d�w��;�s%�����3337������7���z�t_+v���b��{��=�t��R�w�����R�<M	ʮs�]c�G:�-޻wE�n�"h�M�"�.�r@���AO/��@���Eޫ�1�\)p��]C']��9�����.�r����XQ ��{5��z&q����r���#I��}�mEwݙ����� [�V���x�d�N�r�����@�z��ތ�v3}:w*銺��ص8��&��l2�ߠε@vc ����f�0kym�unٷP;XCT�'/Y����U-"����+h�ճtR��e�r|QA*��mƨ4;$t*ucŏ:�Zz�u�ɖx+#m=mBVD~;�oxU���3��W�����x(=_ u3E��3��q�Zv�bG2&f��.��0�D��-lw�A�>�Z��G_pA��u��/�ӆo��]��8H8wml�k�C�+x�k�!���.g�r�����4�G�ĳ�ob�jN��,��.���7@��1/xA][fAw���E�B�!s�զ��l8.���ﻄ|UIB�  v�"�8-I�r�֜���aT�r�k=�E6��<G�NZy��Sy�V�Q�lQ�u�F�R�;R����+9]m1�LUgd�/SO ܭ�Ӽn7��	q9��\��jR�3�b��X�"�cŘ����*�r���T�Xt�gI����<�cPθe��r�}`��ʝ]��N�$��qc2;ݶ8V43��a�t�=+U�<̆�.F�wn�!5V���ÛB�W �ʕ�q��w�6e
���>��b��B�3E{H2��V1�jr��D8k�e��q��� ����@��[nu��D[Y�x��4�r�PVA�l� <���f���s2�nJ7�� h6k��r7���)������j��DԊ��J�*wNEIL2y�s5��7y�L
c�����lizb��m�K7��I5q!+�MƷ:�
�AA1n,*�QP����Цn��LZ��ۏ��ξnW`흌v��g+��ε7	8[Ma�%0K�g7e^.O5!қxw��duCeF�l��	��h�Z`o\S�Ga4x���ia[pIC�S�RNS/ ��oY�47��)�X7޵o}Ӛ-�͐Ճ�� >p�Lx�==N�2�����nfv��!<f��x�c^-�xj��h��P�e�K�I�:���w���l���+l�:�i��X��]�u�tü܌kh}dT���Q`ҵJ	x�cc�n�h�Ύc�H�q�6��IJ];���mq,��V�C�Ѽ�z�ʻ���D4뙦"��ו����\�gkW�d�}�\eG�&�Ч�}���B `�on��I�Wq�ϕeM���nb�����sm���"8�	�Ҧ�t�Z�	���pu��pz.ը�.yD Ύ��r��
�m��u�]�g,LR�
|�q�7*-JUhX�-=�M�א����_[���v:��
�͈��fA��M=�¥�-�3�NmJ{%��k���fؾ����}n=ڭ55]A�p���ٴ��2;R�ڗk�����{'nk��ʄ��j�������;%L�qH/��Yћ��:�h Qγ��ɄT��h]9���Å,��St�[�9*�>v}t�ŴbZ wX��87n�W<�=\�>��Yd&����Y�AR;-�6ۮ}v�[{O���vmr�m$i$(1��	�R�-P`�S��b����"��o�]��øp�O�ʬ�z�qD��"N�[�6͊��b��LfXBq��m� �/ w{�L[-!���]�١Q����b�F���|�a�,�jSq��s3��֞:������� � �����/9���mƭ]t �u�4��&����C��4]�vp�;��d5��oL���Fu��X�n��� 7����������k�9��F��F�K��m���S�o'v�zU)Ƙȝ.�.-d�ܭ�T��<RD���:]p
ˉ�c�����BV���x�A�	`?��˕�R�����8(�G�n幻�/K1ڡ��W!{ݎ�;�v����up�Xкy���T�9�7��wC�b�'ʛ�*��кW�af4n�P��1e�O����h�"��e^��8pӣ���	����jvTLgb�`d��3���Z���qU���;�h<#3oeN@FWZ6�u���/V�8�\iZ9$e��Ί���4Fّl|�*�:�Ȧ��pm�ΐ��]�eTi����=�,��+R���[x�Au<����9j��}��}%�oh,P�3��[ŀI[]���3�64�!t:��ЇS��{�ve������{��h��g�z]�[N��S��%�E��*�]�n��cXOc+v�
��:�0�Fw���[G}4��q̩E����pO,�+�\7#OPN�Jb�u&D�������m]w:�N��	���/h]dv������P��w�����JL��Y�ڳ>i�K7b��s���u*�0�2J�{J�h�\�����t@�fe^��8�
����т�yfr*����՟�q�BI]w�M(���h�
���͍p��.��'=�R�v�w[dլ{G���Ĭi7]cpsǽ9Ú-=
�^,�dr�s������`�k�\%)�ǀVu*LӬ�ψw��r�J��X3��wi]���*�$Y�#�*7�s�}��v�wi���}�fp�c#a�S6��.�n"p�;��rx��;DͶ���{�x��a�JE�#t��)R��e֥��!�x���S���"'گLYX��;1�P�����4d�X��F�����|X��=ίW3��ʁ����4�=����N��\wt¾�x�7����h�x��f����ψ�;�8�p�Q����������[��oVq�5kBweVԊ.�Zk	5´�M���^$�=͕8/p�-C���$��=,R�bu*`Z�9v�4����
en�b�̮��W�qO �(qe��b�4�19Zw�CnU�3�b��1�a���:���pj�����WW5�1�,'m�Z�.]m9�����k�kc�FVfJj85�tݧ�tU�p��]�t���ۊ�Q�[gV�:!�K/�^㕇��L�.����W�J��t��Hv��4�,n�*��{#��よ�=�0�!�b\��e�%������a���,�:|���仧gs����;W��j��!����q�o5�P�E�k��:�����],�;}6+���`�!�fcL�(mAY�-��Ĥ��YJ�A�ĎA�y�t�S�s�6�R�
����%mt��T�1�>�ǯ�m�+h�৔j��.ɧ��͗YP�v�wE�n.K�v�_4�õ,]f<s�̶V�o�2��V$�rΧ�,�P�rWDA/��R�uAf�df�#�� э��vd[Y����X��&�Ρ���@��)��W[�f�Ӗ�V�����p<�:�7nt;�7h<���1A}�{L諀3MZvW4�d�����9{iɇcᑜ�ڒ1HN�Ʋ�Uq;E��gU��u�r��EV%�
��zLQ"��g�dU4�N�is�	޵o����w@o`�2�^p��k���x�ᵜ33J:.�c�n�6;:�x�op�J�kv�W9���D�3i��Hr;�ӭ��L��k�26>��hTp�[��N��XpX���Ev݀m�W�v�#jp|�z&�A�V�2t���ƊVsp�5�W:n	3��W!�(Ղ�[�q��0*?p�씍e�F ��*S�c�Χ�!��ksi�Z�1:U�:: �a�hm��p��h� �K�9�_\���Ҝ����F��.���GAc֦���}�7y�i/f\!�A�3�����`j �N�w�yZe1���(������!k1.B��tYCU�t>�4\�V�i��˃E��Xawkƚ���m]�m��1b�8�7X�[n:S�3��>���!V%��Y�u:^!W��	R���6��m�S��_r�h�;)٫��W�խ8���/����]0)���򩙦�DM�n�8�:���;�-�f���>Ӧ)�ンX����l��D���%%��n�8qم0�W��`�'Fzg ��l_�2�!N�b�G�)\k�62mm����ԣ�Y'��.uǷdy�Rh�xt�X�z�G�㦐V��wH!#��!��'m�y�*��
ck��yw]��R#'ǻ��B�y�SwMÜu�r��3)�8M�(�>:9C6�8�j�1mD�#��"�0d|�e]��tP�'_>�P��
r[)�900����i�)�xE�Y��j�b�夓#z̭��y�6�M<�^�r�gHD|2,��b�*��}�mwsȥ>S�X}6����]J�0h�}u���4"���FKUDd!��%K|���1e��Y��{׫:�vH���YT�QPB	�t��}�n>�Va4Wk[d��<7�C��ތN������8b�6���1�t���6X�0���"ŨK��c�ku� 4U��`Ǹ4��徫֊���B�${��)�NG[uu�(o�� a��r�����:):��t �]�wu��w��z��n3YX.�.t�ƫ�h�4��t7�_ �͕�����w:k��U�=R�b�*��F�ԼqҒ��N�������Z�����Ӌ����2��c
����:�}>�N���R�ƴN��{#�M�!�ݼ>вV�X� �N �ėH�4���kbva��Z���,�o	�;JZ3���h<1Sz�sB^��^KG]�t���p@̄�J�,��FCHVh�A�O���ü�w�g:�2`<W�.u
�"X����0�Ԍ>hQZ��S}���x$l�48� ��2{��X����zn�>AK��z�q$v���#��t�� �n�n�wC��u0��>7k��꒸�ާ/
��;���CD�Wt:��ՕʂU���rt&�AP����O�=Bhɰ�����<���¶H�,O���n���%ɋz�W���E��3Jw5�T;�+�j�>ǯ�h���R���C�S�G�w��x��G+�����v�wGG~�@�GIIq��c'�6�'�X���X5��9�8Mmحo�lE!��oV�=�_!�R�<�7��2�{4N+��f�9���A��8������FkW_D�\�*c{po tHt{�)�	sv��4ߐ���ɬ����9����6qs"�i��뮐;2e'�i��!��v^E{����o����c�.�;�;��[��(m`���s�U&�e�Ϲ�5K%4"�o)maG�*(���06r�k+��FV����&�<]e,J�ܮ���4 d�q]p�um��]8��k{雋$x+a;2�֋k�;�5���Vt��t\��D�6�-p1jR��큱��]nĪYSI`��ܫw��%A����qΔ�M��QGA�a]t(<콻5ùΥ��5Ԁtd�]$HcVv��=�f�l\Q�p��I��.y���K�5n��H��.;Ɋ8�(s���#�z�s�PL�LS2���;�n��E�c��/��WL@Ĳ����-j�cs0T�5q�]���=�ءk��5;��`��:��O�w�y]V6nl��a#�ʋ����W	��K{|�hop4��@v����v7�_i�w�F.Q��oS�������1:��h�Z2j0��冻)v[$�9���M�W��eod�);�eL��J°\5�<N���WI%��[�@�ub�}�s���v�^�Ғvi�XI;'�:�[uғ��D�o�s{M�;]����J��y���HԸ�K���Q�*�vl�lX���ޛǬ�����%�+�	���@��AZ�;.�
�;|���ؖ����Q7պP��y�ã��E��:<��u���_f��8q��zZ`FcG���sTK�0\ ��â��9ǊQ�S�U�M�Q�*�hЋ5s�i�cT����Kº�p��R螓��Y�+A5�-���2�{�*�q�:
����ݗ�3SW-�3y@p�����s�V�R@&�==Kq�ǅ�gd}���]�b��ۜ�cTƲ����7X.a�N�e�D����{ur�K�Sa>��U���֬6�9;&E�ۋ/�<�{+M��� ��nU�c[�Ow*]P���O���M�u�,��	OuIY;q�9I-_L��C�5⺂!�07�9��]R�b����m�]}�]��m��w˘���}��AH�ܨ�n�A-.��z�N'DV˦}��ވN�(_s�uJ��{�k�����²��#����H���C��m�x�ٻ�CSzf��B���������ͅ$�V��vhhf���++�������/)�,��D��6n��elh��C*���}�5�N:0���t�=��6�1	�x�
�l�e���1P
��hor!aݬ���FP�UA��Gr&��*$�ۧ#L� �صR����Bd9b�c1�ˀ��t����!}�%.ڙr7\h�+b��ϰ 㹂r߀��>]gM F��4ՙ]�ᮚ�N ����f�_���kT�h��1�������r##���3�we�I跕`4Gu��j�H��aD���k��������-J��9�c�j2J�Ɏ;h���V��M��]D���W����+�������f,ݖ���}�8g�x3�^6�۸�ҴeEZ����PY���f-�#4�a��i�k#��yaµ���s6�L��u��ԟkJ��ff>�F^u!�<���iG��|�@�R�Λ�M�yXӨ,Te�ƕu�LN�Μ�j{��)۳`\���c�mB��aۇ���AԣɎA,�[bs�Lx��PS}�Ϻ��^6]�}�}�{��7���y{����i�~��Dd�Eb�~��M���fv�Z��r��"�n����X����;t��5J�>6U��ACǓ�c�ER�)a�hJ����2U���s@^�U���:ѹD��=������ø��t^\̥7n���Z��L��q7JÒe-�{�N�6�<�;hi��E���ҏct���O^��%���F�u�����H�{�.,�ب�u|ޥ�i��_f�d�OS�eN+���-�(i��2��x��ޠASfY�77��Ϳ�Q�]��<��Qbg�A��ta��'�*\��uf�rM)q����uP��n�$�k��E�e��\^QǓ��lKY0ӣ��b�E)}��m�7��P�i�U��.z�΅ �fg�|l���6��H,��]+~�rδ�7���ܾbg0�X�@gmnV�<�0xm�!�:��\��nF����8��v�����>Օ������zJ{��#\�"�J`u����D^�Lq�T6�\.��L�sYYu�d�}̬��݇yr��"�����W�L�I��v��%��݆� ���f�ǪAݜ���ד@-0tNZ���W%����c�ꔤ��3���N���ˡN��x_+����`��#j������y��a	\��'u)EiKX+:WS�LU�M�)`�Y�:��X�*r^r�r,��ut�������xc�M�Wt��pv;\�.�wI\��ӗ��ݺ�ܮWwr�����r�L"滝��77:[�7�gWuw\[��:]"f����[��n�+��������Mr�f����]�5�t��չ%��͜ݻ�W9w]�A�n����Q�n�s�����ή����Nd�ƗN��ͺm$nt7;2��.;��:��d˝.nL��wv.��wnwg\R3��C���˫��˻��ήMݮ��w]�s&�p�w\�$���M��ɝ���tӫ�s� �\�	�d�K����Hw]29t��)	�RF�p�p�fa��uӡ\B���t]�˻���NN�ݮp�.�fHNt����܄\�!�%!4���%�܎����D��Bs������;�h���'.1 �>�fa<2���/m����2�������83"�b��g�-��Ǿӭ]4F�ݘ9hԶ�ggX�1g�����w@�R
��ߊ�f�[a|���j����ѭ}�Y�����{�/�b��ʘ͹�G�@����f�ܱ�C<6�n����EĿF��ǐ�b��u�O��[��������}]�@zˡ<@���Õ�C.د
�M�����e�]���FPz��<F��veA6 Ԅ��שc���S=�w���TF��X\o�kƼ"��/���~���ir�J����Y`mz��n�'փ3��bT�D!�Y�V�X\7�z��D�����oc�jDz�N<v��>eT>��=:��zP�y*�vw�ۧ|�E��N����ޛRugh� �X}T�'q�o�/�'j>
������ I�{����W�V��u���S�ze�GM�竣ϕW>xDfa#��*?�5�X���𛧘��'~���)�p�Ӿ^����r����u�ϑ�����Z��뮙7.�������Е�O����!JD&ĩ`D����Y#L���A^�x��'@T"���y�p�:���`�z�7t����Oa"�B�R��^�[��jn��[M	AYҙ �T�d7�5+7�=J�\n�!���B<���[
Rcܴq_��n�r�L+���U�����{JY$�ʶY=Z!�=\�r���y��u�2��N���M�4�jظe1�W���'���ޙ��D������g��Nʰ\�)�}1e�@��Ǿ��g���� �X Tmt�x
�塍]����`�^������}p^5��}HJ�&�o�������"��s�M`�XU����Dp��|;���HU=��S�@U�+�8���$n��Z�e2h��H�;�3)ә*����f�YA�)��bi�j��lΏԐ8�x��VWy��)�]�C�}G�x'J��a�I���Li��R����&EK�o�x�n��`Ox,����8�>�C}{U��I�
{y�	S��>�y�,�5t���U@j� O���Z�_� V�e	u�''\v�&�zo�1w��
���<i����h1��l�Y�@�.�/{Ζ[�C�sx1���G���]|��=�����sj5!��E��dj�:}x�^�\�Zt箘�lIn)^�z����S�l��3:8L�UvGu�l�'��� ���K���~�i�O=*+e
WWP�!D�FiDaZ�Җ��'L�x�,] ����׽>���y��v.#h��tY���hT�@dO������j�w$�nv��wV'6m���čn�B�@��k�1�Һ��!}��k����o'ս$y��l�������N����K��2��SB�����3��L���*����r?:[�)�킷V�Ŵ��ə�l�x�h(5�R�L�=f��h���M/EA��J�rf�y����z�*���RP�6ʍ{i�z�)AvSN�q�!>���)�/,�#oٽ���"`�=I[�ۍ�D;l
S��c�/v̡���H�-���N
�)�%���3t���o�,����iW�J	E������j�Z�#+�\X�e3�m��z�X�{�:ύ����[@w ,�wG���)SMz	�צ1R�`"�,�a)�pt��/z��G�}U<��|��O���>W\@��}���A�]�|t/��/�pC>�&����uN���v�rX*x�yk�o���.�n�&x"x:�� *���>c����:�EI.t*M����p�X��E�D6�'�d~/@�+�c�*BD��t5�cD��_��YZ��/��Si�HiT>�7n�o��0I*������*^ü�U�"Vw�Gx����e'�w�{iI�&�����ޙ)ʻ&�iq�%s��:����ުL�9i��h�z�����Vj�=d#�[L���NS4j�*,�,|{�m�@rќ$���m���&�d�
xw�晹������D�7Q�b�脺�����f�҄F�y��__�O�\%�y������_üG�����q_`�n1�M�&��(��R���c6u�w[�^C����c��A�|��w��C�R����j���yJ�D��B�U�+ވ�6=���\�^�Ѩ*�;�"��E�Pz�|�V$,ba0�AR����i.x�z��I��~�!�?��*)�YRL���!��X+dcg����W�>�@����E3������Ed�ļ1�5}���
�ƻ��=�R�VP�:=OPدO ���	�<hO�z���(Vk���O�l�.��NS�:��c���s�yG�&'�\x[��?���0í�������	j�]aZ��R�:��j`_N�=��㵥���iWSKЮ WmbB	u��x3�W�]y�_�K��@�I�9�,��9<�$m�0.c;��_ �#��mH��~Q�E�����e!;p��NV&N���Wsx�����w�	f�}
���P���D�>Cø�a�qی7�_����z������������7C�ϧ|}��	e�#Zp�<\%:|ַ�ìJ2�����ٶ��臘��} ����Ȯ����#F8�uv���#�7�Oq�.W`�貝1�qc�/���gusD�
�-`bs�]�*�'>kN�2���x��ZTAub���Nt�m�Z����u���x��F�W`ew]�S��`��k�x���r�0W�n�3���*H5�8���بlv�jZ-�����>� V����'�qӧ�{�����%��P���:3O��w��t���J|آ�4�їX�-�c�f�9�z���0��Y��� �0�l����r��uG�̒�[!	�UiG�K�ԗw�i�&�������Vk���Q[��B��Dj�tz��5���x�K紙��lHXF�x�ݝZ]��3L������	��W���Ҿ9ly��՘_��"��ғ9��M�o�����b����s���F�O+���<�]�G�
��K���<�[2�ֹZ2j])�묘\ڄ��nEd����p55�ӈ^)��r>y��b����&��5�L�hN+����5������SSO�����b�V_�W\������oޅxNs���3AѶ���M�˯Lb��̼L|!�����A	;P�����P���zw��J�%S����AZ�o֍^s��[���f������QF�㰓=|�y�_ZZ�t�%4�a>c(��R(t�i�#��c�1����+4��D���uk)�Hss]p�����i��vZ]��VZ��K��-���t�t��;�WCC�����\#��*�� dn���Y�{n�+��tTt|+����
UXx�����:��=����vtC#�S�X�w��{{m�$�GC�T:F��]Bq�|'�_+Ey��X�\b��%4MTƻ�>;'�^J� ��ḻn��q�`$�Ihz:릐������;̼���^R�g�j0E�*��6��$i�ׁ�A[`Z��D��fmf���躧zd��� ԸN,�5zbP�F}�HOoL�*$c6�|�^�YP��[�64<Y�qw�������*�s�QX
� �tN|
�塍�wK���'��&���P%A`�ʺ/��׉����ȘgѮ��Xu��&��?��d�DpϷ�τ��5Xyp9����z��!>��=�睔�*C����]4�=��z�}�u5ڮ�yl���ض���-ڞ��]m��|p�8�5 ��~�S��X��~#����@���S���t�y�>��/Sd�9�~�{��}ü��`Oex��E������8���
uCF^�Y���q�a�8�i��Q�wM�6�m,L�R�riS�@��u���
��Â���zG�N�I��^��N��-��Y���e+�����S�\��-���
y���E�t��>�rb���sJ}b��ؤ��3���09ۜ����&ܜs�N�z�����vm�q�%�j��UP��X���S����@(���V�{�;|���=7�gn{�3S���xxER�c��^�Yް������\>�]�T�:�;.��{<	�ӑ'UP��Аױ]{J 2_��W
��n0�Z�aʣ�q��b�P�����!��v����ԧ�nՁ�_�B��_(�X3��\ ʫ���]��jr���ͩcz�[P}xd�=�pU�c���chVwC�`�Z�����W��y�.����s6�P�Ϩ��T�l�g�k��51�θ*���Y�K�x5B��"����P�RW���j.�ц^��}uCk�j53�q����7���y�3%�!�Ӛn�y�%^��t���XQ����*�1]z|�>���>�L�d�i���#���R��t�5i̛:���HAd� �2��\$������\�0_�/q��!�c�D��/E���a"+l!�cʛC¾��udw _qt���}��t�U�:�,f�e�ԁhx���^l���̛�K�+bYG�+�����{�7@A�1z|k5�z+I���$���s��õ�Vgc鑋r�NB.':q\5���X�B����V�bQ%���Xc������C��
8^fp�D�5���h��|�s�p��d:������a$�z�������#y1�:�y��� 8o���:
����t �\}=X^���87WR''�v	
v:��	�U�b]��x ��":�.���%[��V)?��o�d���)g�2��������*��A^�s����S��y%Vݑ��Ѽ� ��N�~��^B�1���
��O�$%�va�3�`4�U/�!�<늩J��B̻�ƅnI���(��[�KO��٘�������J�5[c���z�n*�zm&����"R���4\V	������}�s�!�X�oV:{,�,]׵��~U~�G�{ظ@�N�:��)v!n�p��)�Q�]������Lj�}��:��ƅ?��6=��uW:Q{F�� ��^��W4�}���3\���m9�y=���`W��y�?~٧��&��tH���!��}�IY+2<��e���������G�«5Q�T�ol��Dz�� Y�Ն�*�,^3D'�X�!�24�$�)�p����'E����<��p|��9�Cz���.�k�{�?f
/%s귡�KG�_^T�SU
��.X�P�^�g�R��iF��t%Ъr^�,�-�TG�7WX7���t���,͢�IQ�w`��/��wGzX�5:�a:���R�$ڝJv���w"��r��a��o
|��*�q�z�D�������ݮ���![=EX�O�>LS�\��:��i��F���ҡ Tƺ�^�f!��ppWgl��}@SF��n�r�QQ�Я���'���sĄ����#ֹɞU���/�J�!X��_�	h�X�L&� �G�?`ڑ���'��l������
r��>�_�L��6U�w8+�6K�W>Z�"�4`9:FB
���U�ofM�z��/��-�l�t�߆���ô�����O43�>=+�h"�u�;5�U�vL�u4�gNX�fX1�L㠔�<�^üj
��V�^m���<x>��k��Q�Y���x��v��p�p�Y�ziP�휾��3�Qr���A�聉,����׸��6�v�T���Ǩڒ����f�"=�jE��i��p���t:y}�yB|]xWE��YіVI����� *����������t�D��B�zt�]mk��^ξjy*)� m��dkY׉��	��N|T'|
�	�Nj�a�6���_�?,Wd>����o���֢�Ա�c�a`|�v2���
z�*�Ƀ[�;���V'���on����񼷍�b��l�E\vf*-���8ͩ�/��ٰooO2w4�2��o�0`\A�ظ��8R�ml�.����Q�%|�}L�1���eP�8r�zy&w�� =eО V/y!y�n��Z,���Y�MQ�
�^���� �cl�b�U�u����m�ӈ^)��o�-�2xӰ��5CN�57���s��0�\t�x����1Կq�ep��`�>��~��9�T�F)���s���,�W�k7����4��u�駄��B�|�xx��#T�{(g���8΍Pp�)���TG�i�T�J�ɒY�{n���'EG��/��K�~ R�< (���/�M��������H�97�]>%�^��sϕy��sp����t�z�8�g��/yo����$ȶ���8��ݵʢ��P���f���s�ճ&4�=w�[��Y�|)FE�8�I1j.]�u��hB'�U,��A`����)d�E �Ÿ#t�m7���$\�N�{ ��2�@�5LCi�hϢA!=�28����P�\k��d쨩�H�Ƽi���^Y˔��3W��<�* ��� �=�·mN<�z	��x�C_���ޛ.֣A��ɗ._^�y҉T)vsTg6�c��ϸ!�Q��z�-�zܻ���!�7s���B=��w9T�i��I�*[t��T�s�H���y��j��h�vb������9O�v����\�aR��O$�gb�;��)ohQv�k�N�d��{iMy`��T��g�Ŕ/w�)��i��73.(.�9�	���5�Y�dQr5ݪ����?NCw�Y��5˺G$�Qh�0uc�@�4(��Ѽ�&} �lN�b񮾨�Λ�7�,m��mJ��]XTSx��{6�m���cK�x�f�j]Vt�c�`AM�K�Ƴ&<8���NqrJ�B�#��i�Ŋ��ٳ���n�r�{ke�6�>�X΍�kv��Z]�s�L�<��VV0��:���fF�Vedvkx�P��-�Bŝ��Ҋ�3�ks&2V�/>ˢ~r�ъ�k%��+7聹W�u��	x[���]�FF��t��l�,S�cK�w�c�*ظ��{���|��s���f��NH��Lb~��Ս��}���o��Ι�����g1��5b�b�g6-(�����Z�n%NӃ�ì�[S�v�{�gh� K�]:�*��(��Ԍ��:�j�nL� 샕�j�y���Q$H�.�`��k��G
�4U�ܽ1I��h�@̼R����|��6�T�/Or\8b��*;z\�J�Xi��3N�c����#�5���Y��TDM�����#���,�u���+�X N�a@Mu���|����]�E>�g�61<c�V�h2_J��U1����r�%��ArCy��ր�=��!��,wf��c�D��40�VS@���gM0�#��8J���z��+�r�T�tyۡ����ݓgNޣ}���������pr`��y�`�ʂݎl��y�:���є��	,b��8��c#��`j��Ι���g�/��.|��S/[nŜhh�qNi҇a��0�\�����8k��np��Ί���m"}�m�b�D�[��p�7{���D�J��,ݑ֓���K0���6o�,6؃SD΋������\'&dˢq�T.�5���]�4R�k���I_V��Wn8~�=��N��s��J1PиA��<�i�QNӷd}�k0��k(��ܺ_Pg�Z[Std,qY�Y���1���ݕr��'�GͽXkoK-����+F�tq[A��F���m�d�s��S@�GWw�[��Ñ�ra�ASg�P�{!�1���ޝu�������xq܊���]�fksJS��A4l�w�Xad�=���*�	�]��J㊰�܏\enu�(W0)�$7��!:��N�lJ�]IH0Τ egv�rj�X7+���ۧ�>�@>Ĕ�}�w5��+���o���͉�q��Sk\��[T�	���Q;�Ouk��2���׸��҇te�{�k=���.�z�\ws\�z�g��XUհ��X�gv:(@E)�k����3K�λ�\�u΍���J�� ��ˡ��wrRh���ݻ���#��es����;��&1�3R��݈s��g7	9t��k�4��	w]ݹ�pr����˴C��vu�v������0ûq�wM��wk��.gv`wwNr���.��2�䂝ܹ�21f��E�9�n�g7wn�B0�Ρ2��˺�f��;7�]D�C��D����v�"����i�ܺL��.h۔���Q��N�ܹ͜���ܸ���fH�ے�!;��F3':a�:�E!�3$�8B��ù.JQ!�ʃ+���8;�1�#w\���Ȍ��"A ɤ��d��M�pE9��'q�s��1���C�\��Q9��U�w;%�\�;���$"�wu�Jh�2	�DNW#C�X���N�w;�k�]ӓ��� &R����P�wAr�.Lc0��	��wN�$�fK���wq�q9�r�Ӊ�@\�nӻ�}����e�X��}/�N�p�y2�8���lSYb���>|��F�0�f�ulv:��o���zv���u�{+zq#�PW��}X)����)�Av�Er�����W����ھ��Ү\����ν��r�}W�o�۾u���i��߷��ߣx�;3'`�LWO�������ъ{i�w<}��-%����?�����ܢ<���f���ϯ>}Z�o��ݾ��ו�������z�O]�=�U��ׂ�r����}o;W�ڿ^7��~_�_�}/�����*
� �� >�+�:��Ѻ�9�7�y���2��ٵ�����Kyߝ���z��y�}7�n�žwzU���6�;���-��\��<���ε�����}�������p���^7/Ƽ�o;ٱ�]���35�M�=�E {�sW���������x���_��^?Z����=�c����ww�w�2�Nއf�jJ%���鷏�<���k�������yo�_����_޼��r�ޯ�}+�n�X���eY������{'���Ϝ����ߍ���k�����/W_h���
��Ұ��~��S���Qh�������}��ޗ�G���^�"���{��y�77�����Wگ�͵��E?��z���v���cItf�ݜ_�����\.m߽_+��W���_�}�^��mʿW��������m����z~6������oj��o��_^���\���&���.���w�3j���x<;oWd3K��78v��g=g������#o9�9����>^���W�������~�����^+�߿-�^5��W��~/KA��������Z{���K�o������m�v�W��o�^�7���~�}�}5��"�%��M}D|�� �Էh0����?}�>k�����ү��<�7�ny�ןw��Z�k�j7׿�o������~u�5�ߕ����W�/<�-��/ֿW��ߞ��W���}z�����4;C�o\�vfN���������������[�/�>����DU~��W���+�'Lyݛ��0'����.�k����]�;Y����M�ۚ�����__���x6�������zx����7����xܼo��h�����O���C��k#�nb�Y�'�z^��|���?{cs>���x��6�������;os�z����^�w�_w�����i���}�<������W��=������6���ʿ���������N�ݘ7�ˎ<��n����.Nǟ`X/&M��]��Lk��71��6��RY�&N�4Xj�$sn��E�;	u�����0��#�]��b�/k>�(mN���a�"3���fbD
�a��!�b�+�z��i�Xy�t\�l�*o3�+�wr��pc���-�4I��f��vH7�?���A�{o���h����o]�s�s}~v�5{q�k�jv�8f0�?�۟����v���ok�^/��|�򽯵�������_��������<_x����������=Z�sR �_p����>�_����~-�x��W��^6��ky�j�[�����34���M�O�����G�;'oo[���;����|�1{�ٵښ2�<�9΍�%��a�Yߵ�O�hv�;�lC6;0[�_Z��y���^/���oJ�W5�z��/���*��}�u�oOm\�֑.�.�]����b��������B�s�?�����Q����O�v�^�,$�h�2b�&r�Ù�����;z����>���=�>���_m�}�����+�}5�{^-��EDW��ޯ;����7/W���o�\�\�������z^������K{�����A����ܴ��f��3��wc����f=n��������Yt_J�\�m�y���կKx�~/������}k��|����m�����{����ݷ=�z��j�r�{���i�o��߯L�����]�O*�۹�N�֮�I�uս�z^��|߿?�[�}�����վ����~_=y�~ur�����^��_M�����޷fiv��~�5Xo0v��W�^���<�ֹ�u����oo����|G�Պ�фΙc����������5|��-����[�8���_�⿷~~��^-ھ���z�m�kƯ�w�+���^���[ڼ^=���k�W��}^�y����o}.���꾖���0
��oy�f>Lԡ
�0ܦ�ާ����ߊ7���M�W��y6�nix?�'`G���Vz�������e���Z������^5�ޗ�G�}{k��k���W�:�*"���~y�����ƥ��~�G�f��-.�������=����_�����o����zZ7�߽o�x��ߗ�oC}���k�����\�W���o߿=_kE�+�������!���~�ހ=�yv�o^��3Ȟ|�".@~f��x�O�b%�����s�����Ӻ�?�����x�5��k���^���5�޼�V�^-���?�W�~_]�=�r������_J������\ǩ��vfN�����P͛�h��5�y�T/ ֳ���a��P|�Y���[��M�֧���^YW��u�͖~��3����}Xfʿ�e��+�^11���=D���ű�.��8�	f���#��N�n��/�T���V���Uۛ5��&�:q��]σ�Pfoj�;�Q�����G������z��z�7�n_��z}���M�ۆ���yOξ���}o��W��^/������Z�����}���W�ѽ��ߍ���^6���x5��[�]���c�'ׂ2�����b9��A�N�ݿ�~���U�s^w�k���o~����}+���j���}+�_�]��>v�W�~6徫��/��6��ߍ|�ץ^.��o��5x���x�_���s{o��_�>h�U
�(�����r�lk�?���>�k�x׍��_w�U�؊�����U;y�����3�Nއf`�2D{���Co��oK��_���ߚ���|W���Xlz��������N����?�-Сi��\ԭ=r�e���fhv_���_���[�}z�O��K�εϻ믍�wm��^�����6��~{����h*���ӷ�hv�8�����;s��۟�G������lv����k���;y�V
/4G����N�lZ��������lvhw��}�r�����;^�{\�m}]מ�~��W��K�o=w5��oj����޼������;x����w�x>�����׍|k������⿙����?|�֧ɍ���Uګ������T��V_j�^-��ߞ���m���_Mp�+��s��ߪ����үk�����o���{^��q���:����"��|xϲ�/��>���|��Lp1~��ޚZ�=��0v�y?���ܺ+�W���o��}|��j-�>�{�_����\�ߞy�5�{^6���x��x�k��sŠ؈�/�x������ӷ�ٙ5L4�����({й��M��	�ޭ9���������>�po{W�|���ξ6�oƽߟ<��r����������үk����|�W��[����W��o��W��ޛ�wv��k��L���5��r������!�+��7��s�_����T�}L��V�>��}P�a�����w�;sL��b��v������D[q�����tʦ�7�#;KCf�����~�s���H�:��f81�T㠔�y�dT6<�R�u^m�������ˬ��SH2�|;�qlD�H(����&{iP��R�wc�{��3�,�-�:P��*��J<��t���EKm:���Äa\��� 践t��eSx������<��*3���Xoi���aH��8���x��W{;�Sf�wܔ��%B��ȳjR��>����}wgO�� VP8G"^�L2{��Xn���.]d!��gg�=�|s_?P.eGS����/�?Ti�n�D{�����"��4�����dp��_vJƩ�y�fOo>����W ��E`
���>|�����Dj��G��^�p���$:�/.o�ůhM����;GJ�����)����Vkܫ�vX��*����{�X��PK6c1m/?3�L~��y����������'����y�2�> V���$L���#+�??ge���ŭ��G�M��i���s!�ƚ�e|S_%�Mi��J����^f�+%����l*н	��ƸmЗ:W8���\&:��\~�E��?���8��lJJ,��d����-{�]�/M`L�;�����ЩN��t�x��s��"��e��j�u�ye�/`�xgƢ)23��Lڮu�=��,�͢��4Ժ>
O��Z� ��N_n��ft�;Đӵg��S��J^�߽�>_y��q �Q���4f���eb&�|�Lr�-;ʊ�Ͳ9[|ü���z�cb�����զ�M�N[E ����|8�{܏7����}�z�d�J�@�u�u[X
�m�GV�J|x���R�TM�����,��T�pm�M��Y�c�vv�&}as�r<��tuN��Q�Ǜy��h`�p������^�b�+�S$j׹�nW˶��q�`$Ɩ���x�����������搂�0O�K����`D����#,�|Z
�c�z���x��?{�O`o�� �Q,
g\3�m���)��KB{zdqQ#T>^k�Z��j7fnI5[��!������[�8�7(�8�5�uOD�jo��c�/���`LL�q�K��;�@�ZNtt��7������B@�@Y��yXU��%�y��O/��Q���E����t�.Q����[����N�*C��h��4����SB6n���-87Vz���z�=�W:�*�	�$�\$�n�>���xb���f36�>�u�/�3��7o�Vx��>�x��7�|��k��ǘ_9�|�tB��x4�.����w��S���S�i���ۤ���ޤ;�}V�,�e��ym��<�r��y�k��/��]��n���eS�-���}c܍9��+�^��[�Bڪ
�1��5�0*]sưpyR�c���镛�`QW�e@���ym9��j���Kьg��0po��1�\lN�3G�}��I��w2�W��칥���c�Y@��f�L�o�Y��f���H9����q��R�su��bf�_-w������ck0e�:k��L�]��(uΊm(�tS�����	��o�,.���{���K�U!�j��WÄ(�x,�W	�О�Y�����<������6��ئ΄�a-]k���R�eW��d�*�����k�g��6y��Y H=��g�w;_pW@ꛜ�%_%\�	�}�x+~�E��E��q�`�w!F�V��&G�����3��@5<>�j�J��h@{�[�'��¼:3S{�]k}ɡ/k4�)Ԑ��$΂ϯ�^���F��K�[JEV�������y�.R	*�{\��ܶ���R�k����d�X(���`:7��x4��#��U�b�G����<�fW�;��p�=V|��V[�{��G[=GVq�֜�0�̭P>���Ү�POu���~�Iu�Xǰ���<���ZC&J��e�,*Ykh�S?�r����0Q��7T��Z���K�Zc*I�6؈�֕�J�=(�Z1$FC�4E��&8/y#�@����ܨ	mp0�s�Mݧ�GN+���,ݯ9PH@S�м�&�S$�i�TӴK1����4z#����5^o��dt�*k�@�a����\���������>m������z��_m:�
p��f����"Uw��W�)&k��kt�E�
 m]����6��%b�p��܇b��+�V���]׈�%)���6#2�;��]��r�cz87�nm�}u�.�m��d��P
��a�Dt>C�e�t�
�mt��,�m	�yf*m	z��Ԥ;���/�%�'���eQ�T$ۡ��QW:��.�$hu��`4�U֓V.��l|������0�ӯlc�{3|��ӫ�U��B�ƸM�/�3��n�%
��~�o����s'���G%淪�=�~��Xj�On%!]���|wF!�^x�]�h��,,%3x��"2&f`���֓*���-W�&)�V4)��1�cЍf�U-^c���>	U���{f%��i=U��T���s��
�O%�{=�nUCCղ2Xi�E>b�	�W�$DI�zf�d��C2שjL���銡M{t��[�	V|'�y/
ٞY�c�Y@�D�jYU{[�����3B��CW��+g�C�^�Vs��<���]ǼS53}=r"���ՊM�%� ����-�Ы#��`�</���#����V������P&�w�-��}΃�{�)y�Jtm�CV�H�ƍ���t*���'Ю WubB��T&W����Z�z�y����QL������ܖ��%I5�;kˬχm�$Gy�xtl�\ੵ;�㹾���8fl�9�m����}q��*C����-ή���Ş����5#w,\�w;���ֈ��z�緝Z�u�7�"k�3y�b���I�j�4��O���'��9}�1o��k6�"���YH���%���K�}�}���&��X�e�l�R�pR͒�m+ʰE�Hp')T�u�������W!��=��l�4�D��Np,���ɧǥx�+����r��$�}8��8�$!�t���]
�*�瞏g�ޤ�[��8-��lyV�����3r)F��ʐB3��,{�\نP�� m	���a��8/��pxϛJ���B4{�5�+/r_u���;B �o���q��4���D��:<����I�����e��C��r=V:�^�W��&�V���^GrP
��'}W���JK�R)�A>�̷Mtzͳ^�sʒ��(�3Ac��۹S��3P+�5ӇH'{����5�xFY k���C��MTa�+��"9-�٬u*#�uXj��s����{�#�x�Z��lf�I����<4�Ɗ�/'0o��̃}B/��Et���.��x���[�^�N�z�x��%�}�DFU~�Εm?L�k((aãC �Y� 4:���n	�����pd��8<~5�Wv=.�t�q�G�e���n��p^kǤ.�ǆ�u��t����2�G��:��Y]l�wKk�յي&�:
F�mD�p���м��bs�Me�9���ꇪI8����ꪤD�os]o;�L�,�^@I��Ƣ���>���LK�.�?l����*����н.���h	b���n�V����=�O�.��{�@f:7^M<"v�k���P�٬����ڕ������v���,�̵�ԣك}��_ɒ �0�PTuT���՝�7yE�ZN_�ʹ�wvZ��Q�D��)�i�L���<�}��ͬ0�;��b�&`�Gq��[e�2Eܵ����h����X���]AR�0��˃����@m��	�5c[<D7��_�}����m�C�t�AvAk*�F���FY>�����N�z��z�jֹ��3	z���/�}ܪ�S���3������F{T>/�V�4a�J�vl���X>sV
�}��}D	̨
�:��y@�S<�1k�_����Wa1)ʵ�j����,TѢ��J��{ʇ�����t�`3h򰫲C�F���+��A�.䰘`��I�\�����[�e6��_]�����w�Q��|-�J�sZ�gq�ͼS��nH>�QǝKy⼊�M$�Ͷ`&d�d��O�����bIC"S��O7�/^ �����6r�weL�ݑO���u0��SYS@v���F�y��]�va2w]n��mt��p�Փ�s�7��Wꪯ��E���,�m�g�c�m��*��eY%:�[ �x�@;�x�O+��ӷ��,�#���7S��<��=������s
�x��DF�.�(���0'����������������J�3�z�[���Q�}ʝKTm���j[sy(x�4�/�,�zz�����R[{=KR�zy W#Dl�+�c�u*5�`K�x���Cau{eu�w���C�{� g G���X?�Ζ[�C=�I�%��u��� 1E��@����[��j3R��v��Ϗ�x��o��w�q^�W�@$���Pm|��2���ZMX��w����}u ���|�xƽ{��w��Y=�^��O����wF�]�4C�M>��o�����n��Jd3v
�g����gFp��۟i���Җ/Kb�c���=�}��[�4��A׉�tN��4�]>@A��%�T%E�qȖn��7����b��%��)e<VNo�+� 4}��Q��0+�1G��Zb�Ļ�)�������m�"�tk��-`��ήG58�K��>�aR���e�L��ri�������؉�l��ӻ�ͻX-�T����Z�|�⭾:�s�g����4�v��v�tT�����ؙ�jg9Q�'L��T���xP��w�<9��׮aޜ4;�F%i� TpI���š�ҕ��^����=?����(���k�7��mz�;G�n�C �sĶ"F!Aa0�ݮ�4����٦6�篧+g*LT��5��K9ԶC��MEt������s2eA3��W`�cy���`�ѝ]Zp���p��2r~��eŋ)�lҶ!^��7~��F�Pl帞c1e53c��l#�����]IY�V!Ω�w)}�٢����:Znq|�t��eB��@4��j��Z7lX�4���oj��Rۈ�1�[՛��
:� @��v�h'���hl{d�y��I�}�^���7�݂֚){�ћy+�J�q�yMǗ�JL��vݥ��|ZHu���9om؀M/5֛�{��@iQ��{VPp&+&��Ft��Ý��,S��SgF�'uY��K�����i�2Cw�,�mmz��S��|�Jw�yݶ�m��WwD�9`�[,_���	E�9��z��gf��-��S���2k�&p:�ڙc3MkQ�9�:�އj_�)�t�v,L�d�K�3�.����YA=�Z��۷|.E|"�j�'�g�Jg��*� kh\�����]!�)Sz[����ʖ�H���u�2�1լ)��tks�{�y�i&�7Vh
�-��㽂�*V��D��6:��H���eG�H��WIhYp�n���]�Z�M�9�]%�˗��W.��T���f]���+�;Sl<�vM���+N�n�Fr[�+� ��āĝ��ܒa�����=WC�b�e����H�����n��t�G���S����n�Wp�TM`���۶36�ٷ�"(O��s;o��$�gr�@"
���o̩�U]\����鍧�z�ۛ�Z�kH��ۢzR�-�x2-���N��$r�v��+���E_\��J|�Řǲ�"5:A���彼횰�u�$�I��д���B�wˆ��J��s�.ȢɲL��i�W�W^�6��Jx��#�v�T����XqR���Q6�72��N$��u�&���LG1���T��7R�ȩu]c�vϺ�᝚vQ@2��ٝ��r�vPCM�{�I��ah���%��Y����/1騔�KD���^T�������/��g;HA��Ϻ�3��+xq������v|��W�ߏ	�D�$ۚ=ҟ��[���Ŏ�֢U5����k�f�Y�Z�W�-�� �r:+�9.�5�51�	+7���s���:��#%��hvi⤸澫��ۦV��H�X-�}�ZÀ��\��g#nm;���,5��=�#�wq=§n�y;+�ߟ��߿ۚ�ݸ�ݤ�2�Wv�.�H����	�Ae&s�n���(���L�`�wm�`9����B$���6s�.s�&f��)\�2��wq��ݜ�Ɍa�t�n�l�� b	�]�J7wL�"S���Rff@�И�dA�M���Kwk��"�e�4�1�+�J�1(��4��4�&dL��#1 I˘,�9\wN�wrI����,� 0�]��F1� 2h���C����B�1Mb$�B9s"(k�석ܣC"�9г��(��i��nnn�w7S��vn�r9�aݮ�����5�w;t�;�$�X�bs�����cD���9�H��������4��"���	]au�r�h+��s���Y���s���&I�*�!� �� P�5���y�]��JjjY�ӕw���%��ٽ�#A,�y�łz�̛'����od��c�����F�;�E���{���U$�I�5�C͊�?��q�Ⴘ*�:I�p��U����vhaZ��PO�a�y����Q%��\��9L��ŉb�S+m �����	�w@��e�"���u�<=6�ݱq�X�=R�.��u���C��#!�j�1�1�?y��|@��;�j��W<}�^վaORG�_����otO�nל�$2��dE��ɷ�C☗h�^ .]���t�S���[q}���D$]�0;��f�(:�z�;�p�t�"-�D6�'�dhN;�3Y��w6��������X�ѷH:��c]����0���дj|IT�wȵl)�Q�h���M�Ի����@ʝ���$EJ�Z�u�hYB��?/�~�˛�Cx��9=�ug�MlC�'��>���\W����A�Fl믃��uB��_�B��	��rw���Y������V\bǆ�p>�;gy�u�Lyj���=XЧU�1}c/�e�p�>���#���2�] ��ب)�C�UT��{
���
��3Y��z�떇��),5OW4,v>9s;����r�:�b]ǜ�F�Ҁ�ɹ 2���P<�}�Gs5Զ�AL�֔lc���p��]�޳�����GNL�^�� w �o`G����s���E[�P[���E���Z�E���K:8R�p��Je�n1���h|�߼���{�&����d��w�Ia�<��WmQ�Nb�xAQ�)�Z��M�c����Sqqoe9/Ԯ�����v�ܾ'���z+�<r��3�x�=���܅X���(��DQ"��v?
�|]�3묺����<1�1G��7�9����Sqg^!e�2���`���iPH6ʜ�*����}f����Ѓ���k�
�xz�t��?{��ٽ�����i׎�2{���mʯ-�\�`$he�y�3�i=R�g����L?NK5�����pw��ik&U�e�l����7폄ϗ����XO_ �bY�/E�(��3:wy3�A�=T/���D �4nZv �د����5����4�������{�r�|�T�0��3�,��v�c��N:��� ���1��Y���Kl8q�N�� $gU�};(:�H��� V�P�e�>F=�8/�7��T\��;x"��
��i-�phL�� �)W�YE*i�3�BH���E�3�i?�p��WRb��F|���>���@
�#���[��V"���t�}�6Wy��p�և�gD�^�I��9V�Uu{w��׆���7#�).�ԟ_vb�_t%���g���
޷���O�ϑ���BA�V��J�[c��Ϧ�Bo�������L�ĥ�V<��yv:c��@V�'y�dV ���>u�ߙ���Dj��ѡ7�v����cT�)�x��߫�UL5%��Lc]8yJ�dD�PMa�dg����d**�5�VN��/-����l�*AV�*f�crs�� �uܐS�K��W��ҫ+<������ `�w�	b��j�	����5e]{t2��SE��L��1lY8s&Q0���L�K;�y^�-o(� �1}���J����1�/������X>�쀎ݡ8aw�oӪ��Yà09��VV޺GF���M<'j���!C�c�ʕc7��V�K���-D��G��u[=�L���T�tV��z�b;REа31tN
���.V1�-����D���,�\S�j�wv�XN��3�D�Jz�^J^��sϗ�|��B  �w�z#-p쑸�e��p������v�r��%�4rFq�]�^��a��Hq�1�^�&Ja�Q!V�S��p� �n��K*��>�L�E�DM�K !OC�whxũ��{���86�6�c++[
y:�D�"'��e���7�
��d��泰�!��P][�Z�x�L1zqb�T�4wh���@��xE�x{��Lf���î�wY��.�wI��L�7��lT��\3���A��h˒Es#0�}Q�7����kho{�C/��2��G�����a��!�&=���ޙTHa�B��A(	wڱw�um+_^�\+���g���� @� S�:+fy�o �ռ��@��䙊��7��)|���߷�JK�����x�����`:1V�.r��!��s:{#���t��)���FK�Qs�2v��1�S��)SNDQ��uw�:��K�����k����Gjr���CXn����j�q�=�)c��`�!�q��y��o���+��-�~��D+����m�kQ��;�>Ӱ��(R�}V��͍P�$C����/h�1��1�Q�*���~_y@�K�*�5�]7�ݚ�����=��bn0,;����'x��IJ	�=ll�@�����
�s5�`�3Ƴ���6�J�C����h�3�U�u�|�!S�ׁ��:X^�cPϫ�d��~��2�J��WÄ>ά�#�<�x^)p�,!��u�\��]��;eu�����]�2�n�k�%�f��E�I�z���%��:��F��l��#�)Lb�uK_EXݍ�k:�<Λ�
h���/r�
S���j��C����n��k��]�y���yń�h�ԕ.�%������DP�:�ז�a��i�Mm˖�i�Xl�j�i�����oWCɥ��߽0�CwZv����p�{��شS��Z'��k;�,��Ns�U�o�}��uE}�,q��i1�UH-�>� C��A���vNm��ו䩋ݐ�Ʈ]9�"����`�A�G������%��T��Uo�<5�t\�"�(HTd�gP�Y�4L[$��t�#>~:.UܸQ�qc+�0P��!��N;�qW]�yz���4@�Nz��of��B4�&Pϣ$�L���#էpWI�t�C��U��J	�/Q�WR�,�}S�Df<�hP�ޙ'�CW�C����,KJ�^��E?�LxCc9����)?�y�fg�c;�[e�R&
���t����G~�7�Dg^ˢ"�Z-{�[� �g�j�T��>���&�B.Y���,��ݯS��j"ݑM�IL=ꩧhdX䈽�m|�����8�����p�w�#]����-�p�}�i�mvNYDY ���e�v�8tͯz�P(n�����!	#ұ1��x!\%����9"C�ǡh�r�\�QbZ�5�h]"�i�l��t�}�z�ۦ-�sr�N��Z�՛���u�6��rTQ]��=��c��:�N a����.[������uC��%��.��t9�2��T�'��Ʒ�%Y;+%�4��e�O��|t���`���pLM�:�Y����U}�|evv�S�;�����lIᩭ���瑱HϹ"*:�u�t�]`�\��ٮA_-y4cUkE�ޝ�ԧ�ϵבUP��H:���;��������@�z�;^x��<H,���_k�e�W+"��r�зk�Ԝ�U�w��W^Tǖ�x�[SՍ
u�2��C��\=�������oV�j�/�j
�T>�G��{	*�=(����ǥ�-e��d���Ն�9�w��&*)�*"���d٪?[��q�N �p���~5����q2^�h�H�
�rG3���G�c�^�5}�+g��=�i�3�	�41�����M�� ���3�E٬ۮ��5�82�U���\-�
��ߓ�!�^&= �A=^�W髨p!Zݴ�736���c.�*Lk�"��vڇ>�@Tt7�Q�^��Pr6h�u�#��ޯu�0
�$1��}�u���N�����Pnu�� �b4���7���o��{����R6&R1��[��d¡����R�p,�/�j���0Wf7H���=7�v |�o�
d��N2�~8.1����I�R�{x'�p��C�e!p�D���:�.,�G��<�D'gt� OU+�4�K�pfi��Q]+E� mN��)v�B������}ÇH���ѵ���O�ZkF��7��7���EP��@���@���A8�a���wIp�_uׇi�g�
�O+m�i����[�J�P��}�h"�J"i�ܙ��P�f6�T㫄� ���j�Q����OO8��{ �Z*v�[�������m 2|��.�*���f1�Nzv��([�&��uIMz�/o�� ��@ĕy��R��3�W� 94��Y���Hsi;l3Ǎ���>���m�rC�Z��(�d!;�P������#>�d�K�:�i�Z�Kbt��u�Ľ}7�zŭȏ��-}xT�k�7�;0h�#}��}8�Ϫta��60�R�U!�,���XC"�FFX�V�����)��j�хC������bQKi�c�l �1qz�4ad����� ��&|1}�y��k��7�x�y��T���oz��]z���as}�����w�`Vo�k��b��\���/�����cX=}8v�z�`�$Ւ(aa1��GT�D!�[Un
ap�.��3��SO��]|���S��զ+[�ͭ� �X����ڵܬC��2��r���D��/V�Iy�K��
�~݈���&��m9D����`�6�����o%��x���ȅ�]����+Y1�G�(�h#`����YI�Vp��e[6���o�X< ���yà��_|�����r��E�(;�a�.����D6ps���A�=�^?t��ph���PT��b�ulKju�=^��6j����l�=�����~n����}׷0�L�cm֓���{��O�|W?�5!t+�''�mV�`7���b��P��˃���l!�Z��;J�g��;牣^g'��.���t�]��'�)�h"&ʥ�р�������*�)ݹ�ӽ�
7������:��܈!�*@X>�Utҩ�ϗ�����f�e�Z�e���ft����5�s�*Y;*���gwӾa *:��y@���s��}6e�=�ºv��^O(k�Q�X��Ex7���*<v��f�^'��՚,r3Z�!7��`��J4^ُ���^5%W��?)�I�Վ�4/�ߏ�W<��;�Ƹ�ۂ��Cԇ��x�x��<���,�JJu¶BqӇ��U޻�7|�+����v���گu�*�Dk�e#��§<�tT>�ol;ް�U��x#�F�x��v��y��3q�w���6�v[9���G�8(�PIm�y%�z7J��;��XUy�a}�-�g	k�%9��i���VqR!�>����Y�ԴWO�a*�S�RB�7�N��po^�*�-J���e���z��k���L������y��V���K�ܻ���w�e�O��~.�R���a�����C��:������bҫ6\�Y�D�{�y�x�f*�c��@T5�#PW]�]A½u�a�/���$�dc3|�Ē`�j�ʙ� T�u�q�Ζ���3�d�T%�����5u�7�������k�ֶǚ��|4=�u��h7]���'�t��_.�	=�Iݔn��;̱Z�I�gLX��	��&}�,+V�#Sk��y�گg֪�6�"ȹ�[�3 ��͜��L�U���������۫SW���B�ͧp�`�@1�'J3��6٘��_a����tZ}����!(T��w���Յ�u�yFLt�Q��U�v�]8_E@�h����}�°���f=��G%(U��t��9�d����s,u�ǆ0gZe�7H`��u&�Y���V��l��ˉ`R�d]���%^��*R�`�2}��Θ���t��fH���E�y�9B�ҺVdj\�tB��&X4�|��S���U۱|nc��;;pA�r���k����Y�Pp�͊�F�H��A5s�G�R4�r���o�JuK��e��[����g<��]�.�f��-���y�ޔM)&&Gյ�VVѸ�N�x�[��ޫB��d�A֘0F�sO�dҬ���iL��<���ڻ%�D�!X���t���L'�s�m��:�qx�1֡����g��}S4s�=�^>��m��ku�Ў�����*yq�'�UA}�G?zi��q��x�(��J�5i�:����w�� ��k�YS��`�Em�=�=�>�H_�Kc�f6�	�N�ב2&�d%$ب��MMlک�ϙ���F"���I+��gU��G�y�9��v��3{�ཫ��Z��	z]��S�!��g{�y����+�6�z�bγhY$��Mj߻,�p���'$�շ����J��BN,�{��4׳��oz��N�l��lF��"9�{ޠj�G�����w��:��:�0Ym���:Ὡ23bbb�t=�9Y
��wΐ=A�Wh�]��Iܺޚy��C$��n���+M|2��^�ew���"�k��%I �P�>�z^��d��V
� �S�f�솀g[�L"&��������K|))K졡[̮��sO0�Ԡ�)�n�q*!"�� �!IwC�'V��8���~H7�F�r��$�LF���(K�:��θӬ��
�I��Lau-4-����e�ǣWѦ��̜2v\�D��H{���������o�;2��56�^�����L1��0A���ךU$��ɉZ�ֺ���#�+{;Dd�h��m=���S ք��$�����疀V�.�7+[��B�*�A+'G�$�����Wȝky0.�pyD�]�����s�9��:�h=�o;L�@�E�V�f*��J�ܮ�]L�:��`'1S��v�Ju��������TSgʘǶ��S��3�@�C	Y3���VU�]��I4;�T�"<�j�q�; Z�����a�V�*�>��a��vv�]�v9*��ŵ�u{Y�9vg4	}��It��\��L�c6���g��!Q�-f��k;W{�� uu�=�[F�������#���@�&7;�O�
�J���cs����7�F�P� s�}D�� ��8�+i�s�s#��f�.Y�'���u���䦢��n��ȶ;)gõMR X�igA�̼�kFt��R]/��R��('WS'I�H���L��Y%�g:g��+/0p��u0�1q�4��ƥn�z�I�D�5�ʙ3��1�ń0��1t� �sym�z����KN�qP�����P��+��Vg̄�T�Ab9�n����ڣy��>z^�V�s�}�������e5��)�N��Ɋcs�Q�f�6�i��L��!k�a|Tז]i�Ӝ����fP� :r"���ͬ��6�T�f������-�H+�ʾ���{�bzmt�T��ƥ�G�VT=�6R_3�"y�u��⽱�5�;��C"u��z�ďW)b��4�A�wwt�z9a���׸s��7���o&�y����b�(;K�\r��w��c�*�����T�d��' ��ɰ��wh�_\��fؔ�LM�R1/oJ�8PPѻ��0M{*�GU:����!ڂ�2�ӘJ�;y=ށ�'DZ)��C�:wVd�	�����D���眣�/���g6ۼ�I4.���*��Z�qM����*�r��Ч\�+v��j��$ӝ��R�ԓ`4&�ݙJeq����H�t����Բ�gKg"�jn�Ν"�eV%��oge(�[�gts;*�i�->6�f�[�ٝ�UC�1�2�L(�����vY��kn;�Z<�v�u6�#_WT�L�_z0Sզ:�����hT������}:��o5��rIK�櫹����Ue��\m@C�u*Jʃ�����G)䝻Ƹ���+TS-������������~7s]4)F,�N�cc"IA`;�D�8č]�(dD��&�$�C!�$h!2Dwt��s���3��7,(#j(�hR�iF���R�b);�!�!C4���RX 
JQ�А4��,`a��Nt�R�R6@(�"�$X���%�H��$$04&�ˆA���K�h��E	���H
5Λȁ��L��Mb��!�0�	�v�a��wk�ȦL6H�DȊF@�wu�"��CF@��l��ፃ)#L����J$�N��FH�	)4)J]�)&�MS
P�H_�z������vkb�mٸ��J��$�;�5*�T�xO����&9�D�y	�ٴ���K�ju%�I����3VW��7���SXd�Ze�&3Y��鉫&����*�uC���Q�WL�׎�m.eb�ՏBZA��D$�F@��$pKp�D�[�hgI��^�����`[nL�r�2Ĵ"�A�5��N��
c$���<�������f����ϰ�ZJ�e��U�9,�NW���lѮ��ٳ�}0���_=��Ή�U7�N�4�Mz�P�͡�c�Y�0&`P��f�[����`���g�[�r+V'H�saIX�!�2@:��U ө�V�cy/8�)�Ct�\�+���]1�cq]�s$��]�a0"���Zꐲ�+l�9⸟��]:��w��d��0J� �,�n�n׷5ԓ�Z�9k(�hb�;�W�������>RdgޝST�R�;�1�q-f���"Y��q)&�M������[v��Z)�SK��c�ׇ�]�];q�������%��b`�δ�z���t/�v��c�k��md���3�[��ݔ����}�4ar��Ö}�Rxg#�!��^�-Ӷ�i:�3���[=�ix���+��y��s�ooPW�x��B����^���z���S���(g<����f��
�gd��9�7�^��`������/�c��:�K}Cl?mI�~�_A&�L�n��in����2�^��E�wƣ�`�T���9m״	Q�ԝ-�_A'Pw�`�;��fع��{0�EG����S-��~ŗ6���,|�`���4TZy-XR�s���5�{�fr%\�^��KL4�jc
�ߘ�ݦ�{-h�mM>܃M9��K��*�&lk�7��>����E��nZ�N��)-�S���W�1C�+�ط�	~q��گ��Zx�@�h�?�V�������d%�i�tՏv�.kz��N�2��n�0��#�~�D���Ѩ1e*�Z�ڲl�+kl}[Us��60l�سr����-̱�s>�âf�4n4�g�m&�M��V�2�%"�N�&��lM{K^��Vu'�c�<O�V�m�x��*gO��[�)��2rwv,P�h>�VT�����ZNSó:΍�����Mٺr�ٱ;�L^Y�{k�A�x�����ገ�]�=�[��J9o'PΏ�8��޳\*�2,�b:/U={�U_&K�5���f�0$͢�4��y����t�0�.���[��)n[%�����e2bR�R�|�;e*��'�ڶ0��ѕ��g/���-(�fuX��v��,iQJ%��8L<�{�܈�=���ﾺb�ۅ|y�����q̶�Q>Ik���Q��X�1�����Lrx�z���S9�A~��h�<�G�����S���c_/S��{�<�s�$J]���]�_N�)a�:j�Lˣ�ҷ��Y�������1�Y
�sΤ�ּT`GShI0��������r|�fZ�����n�0�v�X�nA�"B͚T���)�-JP�J3T�M��{���I�oo>Kr���;�s2��WS��|f%b�b�6�e�Uqt�>d��*00�;'>��TWs׻ʎ�3�Uj�@Ʀ�Y��W�Z�M��Y$d�U�S��g����k�.�G�Qa�թ��������0��n�E&�����繈��k��oL� �&�����:��G'G�V肺M��C���cmKMZW���e��ƌ���xTmviѲJ�ld��u�ځ��>s����e���FHr�@B�I�0@�˲rgm��r�u=ˏv&��U�W��v<��Cԉ������fb˒�U�dz&��f�l�-+E�'�K(m7&ܱk�E��umx�H�TӮ�É��$_����k ��7V�����N�jJ����:6���$V9�:�-�����ޜk����wy�/| ~�G;s�J�t��V�����{��m��^7$^M�_��^��gM�#��R���׈����j�.YL�bk6�a�����q���W���x62^¶7�rr̂�i��&�e���g�/o�fX��p���F��:�~��i�=����]�����Z<�*=�_Q:�k�H[AT�X�(�hs��1�qD��KYW��6�/nhF�T�Bǉ��LB�E:�b�"�����J5�n>L3�z���#e���o7 ��W�Gx߾���{�L�BRM�������ک��3�ð6�j�^��@8��6+M�����)]���f�o��V���^���P��N�*����A32G�z�__B��h��0{-O�����N����ɷ�����Z��wP(Q���{/���S�>�X��٪�'[/�����ƻe�6�ˌ������3"q,�iT�۾h̹���k�h�����K+�IFK6��8�tU����y������BL_[ۖ�ow�.�����}jڭ���%U���uu5��Z�ӱ����=U���{����Xi�ƖF�����z��|���N�7o;�W��6����f����*������G�X5�̵]rn�ᵙ�E�κ����H�)�īim�D�a���5��d%Y�d�#6�b/X0���hf�:�[JHҝ[Ll�GӀE���$��O{(o�s������T�l�kj��ư�Sr��%����a��sδR�KszY�}4��p�(�$9A֓�Pb}d�Z�ٴ�%����t~;m�m��woz�/P'���O!��^04�4n$�M#�ۏ�45�6�3�Z��U�4ϩ����/vxm�i��KK>jئs�ի��K�v�A������F��-{�xt�~�5��tH��.��=�Ʉ Ef��ɉD������:�ݘ"����O�G��0��:_�xRƻ��J<S3�F:��2�HV�u��!�7���;zR4�|yt����=���M���Q�l�V��kn�������3J����R**'o��Rܴ�YZ,�TK00�w�a���d���w�4���*�����ۮ��>҉� ��z.��^QJ%�B���dVk���<wg)m��ҷ�)����-Z��湟�%�Z�:kE�I��(7Ǆ�է�.�on�����Z}TҨ򸖳p׊ΓN'�&�\S�C\n�ViJ�3h��R�՘���-�1�}{$���n/f�{5NՔ�!Xj�PM0r3�5G8x٣(o��V���Ε�Ώ�*��)���^b�lG���6?hٞh��Lu6�m�x�U�S-w��a���)d����6� %/E�"���
�9*���Y��.mU��X���Ty�MK]�-Q�8v�X��U��}��է^F�MF��b�v�U�q�&��1�2a�M&e6Kί8&}-	��Zm��4�Q	,*v�0)mE����kk�گm�9�Q��5_�\�Ϋcلa'��x}��X�'�kO3�ϰ�q�cn��J�]n�/s�==�@* �Om�᧸���C�>(I�H��v�ڥ������Yʄ5ܔݚ�ۋ�\H����hv�����_N8�+ow����7��y�!�bJ0����ՀA7��t����T��LY��
���y�,�1Se����"a�i1�γ��]8N��:�dizu�u�M��o�>��-�,����DB��rX���%�-̝w1��]�7�'��Psz����kގ&:}Cܮ��v�^�R׹*R��X�L`�}�{�f�����N/�r���c�wY���l��ʴ1D�J"�M���\�D�%N�+}�{,�*������WNr��(�gU�_��yIcK(��"}���f��!=�!��V����ލ�s�Tk$��zN��Qja�un�37��"z�^z���*�_[Ds�T}1<�Y�<�FI��5ȋ�9��׸�y�s�i�Ğ������R��<�V����G��oi��o�9�ϕvt���JpD���*D��&"X��5
���ж�ھ�$�W�<-�Aʝ.�[lǇ]�Z)� �swET+�t����Q"�eg��;B�]���k�ZN�Q�	�,��&ʄNo�e�l"�65���2t����5Bl+<�$��ԣ5����V@�Ų̩�9*��ȸ�I�pe�5s������V{ꪯ��VN�ڨ��^&���]Mm{vՔ�O�JIFN�����{�����_U@QՖ�S�f⌽�V�,֕�a��q�V�1�~�9pg>C�]��<��ֆp��'&���4"�-e�5j�^`cSP*ΕW��2��	�|U�[;�2��;��r���L5L��
���g�[c�Cn�M55�����h����&M!��(UyEa�G#ji�G*�{6��T�h�x_�)I�={�祢n������F��ke�8N��1�@�t���=Z������ot�uyv��Lh�n��,tn�c��H�sZw�-�K�uA׽A�l�Sg�.+�O�#�|F�7��t���������R�=9��b�H��r�fc�I�w��9�a���L����WN�Kr�{�hU�e�챝��d_�ߠ�H稅k�܄�N�Z|��
�cz�y��
&��F�-K(���}��5�kPr
`��\��8J�V��]����j���nmw������i��7��^���9>�5sFK��ĺ��3�_m��3����w+���*Ɵs�z�B�2霡U�g��X��<�`�g�G���a^�v9�I������}U__>��������\�&yu��i�:]���z)�9=����vq���[=Le�h��.i���b�D��
����~#��[K�d]�V{S��s֤�Ql-њ� �NS �1�ԫ*{<T���K�Κ��9?l�A��i�v��^�ZL�)��$�8�h�e���|�&�<�fp�o�{Z�z2�}
�S6���4۪v��BUʌ�^,y55�N�͋,��z��u+����KZ�g���{�Yu8_B�%6$��5Ȇ�����g�D��.X�t]1�{�f�'\�����S^Ώ�.w��#���N�������&�i���lز�U�W�Ø��؛ř*����������^�I�f��^a�3a��5ij$m���y+٭�31eȇa����޵����y����	��}��ٲ�e��:�iI�)�;"�{�����{Dт��⛅I^xw��7���[�:����^PY2ۦ�/�ĘMh�'��2���vAh�Y�e�����\�ݳ�)|n��t�d�w�9f'x��30�]�e���thq�y�샠�{����|����S���fga�˒��f���oU$T�h֝�q�-vZi���a�c�U�Ķ��kK^&�cr7:c~�|��T۾4
�<���Dzw!���V�ѺM��D��z���p�M8M��36h�����!���]u�C�nU��x���d��#A3�uc�zйe2M!n��L0lKC歊g9[l)�cB;[v36�8��A���9lV�B��eD�g|v�y�d]I�B�6��3op�eW���G�(�Ak�B�~���_�W%��я=�*���W����rT<6&u��M���g�N�Ik��lE魘�N��%�r^3�iZL��,����[F�=*���}���~��&D�N%�$ذ�CP12��f��p�)�[#$yZ�*�w-�O��»\�������_�������eU]���E�r�vԝ�~��T�z�b�a5�C��w'�fm_YcY{*�I�\�@l�Ьܐ�b/�n)�; �F��`Ὁ.줲�v�*j�Gz���"�m�n�{ԦJ���t����$�_>	O^����{L�� @��֮�Ed<N�cܲ)��FK���6�Y؆G���6����g*+�����hYyV|��V��Z���c�o����(�T�k�.�]p��7֐��&����u�!����:��;MG�xeىѬL���z����k�˷��0��c���mb2�"�z�\z�(,n"����C��,:�-gL��D�/Je�V"��Ì����/��W������2�9R��D�|�<��X�WYVw��(,7N�Kޏynml���۴�K�;75�r䩌�';ؓ��kU���SM�x�b܈�4�*�-z^������Ƒ��rXe�T�&i��8�@p�]ۖ@�4��B������m�<��vc��Ԁ�]X�屹�]=b�S,Q�reP���L�)��k"��d��a�9��+ϲ��w5���x��2�3wI��Ҙ����������-���}$l�]Lv��"(�&o�@!�K�Z�J�X*�sA|1Jgsx@��|/ Zu՝cS��,�K=cu�U{���6�.��t�;�k�sgMiC��|��v����G\܎�y��l&�«�LQG���n&��R�YCU9՚6�`}��79��f.�y`/cw����hU�� �92�uj�P�v{�74V���yZ߹��Ý���u��5ϭt U��Ɩذ������n�+�^���se�]�s̢v-;�[��9z���$UլU�q��G�$����qB�u�:� W��X�L��n^��P{:�[ae��s�w�a�jNnh��2�Vs�O-���Mя1�fS���bi��k���.p����pF�u��;��_Wp��ԭ�_wv����EΔ#�̼}���
��Zں`)^�����L��/N=��r���6�%�X��X�z�哋���|WvP5�Z �$�(�*u��4w2a��$�D`�0Ҿ�.��T��GNo|�j�ɲ֞�0&�=C�y[׵��k���<8]��`����`�<.�r�q���>�޾K�'����$1�Qj���F9ۼ�(��W�7�s���Qw� A��<�8�$���������ľ���O{�\�bX��^@ڤ(dq�.fV�>�k�Ҙ��<����G)���<�̡B���NE��x���&)���9������m<��W���k��*����jWLSz�;�Rn͋z�����u���	���u;{�����X�V�%[ﺖ�����V��hV�Smoٮ�� x�w$�izG)�8a������'=/hE[y�j�Fd���2n�=��wv����־��g w�&��݌-,l.Kd�ĳ�y"ג�]tk�w��(P��@�C��p�#DQ$�f�
g#t��L e0�b*h�	�d��\fPRY�;��3l�I �,&̄��㺸(�4��$3)$$"�.n%�����dlX	�̡%�D�`!wv��k����Nn��Lgv�%�Q.W.�r��"Mr�0"ٝκ���"Y��I&9]	˱` �0F����0�9�4d� ���뫛%N��Mwu	%Ν�K���Ƞ4Db�"Q��FF�Cd�"r��Ei�@`�(l����߿��"�(�F|�)Fw��N��k��]�<�D WͰ.�ou�[Ƴ����{���|:v)�)���p�u:h>�fo%;����9139����I��m5���r�������߲o���D/kE�VٹT�b^�2�9�����R�Y��Ow�o���0�K'����E�N����M}�,+N��Z��³�Ss臨*�s0�[[�.�o��W���U3ᦃ-ƴ�`�f�B����T�xOw.�4s��Y;K/��$9�#誁�h�5�9��uXz��8���5��������ח?X�r͕ ��ѡ�Α����_�k��:���/[o�wMVl��7S��J�����`m*�ng�]�0��쉿����0�L��cxX���l��ˉ�)]yGm�5��׹*R�`�G�q�2�)�3��MbP�lF��`���fuq����b)n[2[�*���)��� ���r)�NR�`��Rfu~+c9�j�t�i�bW�.�RX�ye��:�Ul�-He5­����5�ñQGk�t��+R_k���5;����&{{.�YG]������3��P�pa�6��:�ΰ}kv.��y��d�ȲwrLj2k��Fh��R�u��zr�Uj!`tN�bˍ'¹�������d_hy�����ꮘ���Ty����55�)��y-u��-�[0)f�s k���
��J�mvY�\��-��V׈Np2��UWx7c���'&�^��SCj�q����*���;�kMF��4�E�$&ݚ�e�E�iI�N��g��5�E��u�ӔD��]i��U�{*��ϳ����mg���6�-�k)��3+޼[�-���L
\t6#��7ۋ�1bן1K4R�m�٬�k��C`㒭�	��`5��_
�N�O:�J�/�;̠j�ȡcS浖�Z���ML
���+�eU;7�i�L�&V�Sf�2�N�fU��G�GW�u9���R<M�2:vU\�kL�D��CQ&���)��6�F��.ET;*��g����/f�5�y˻û�^��Ach�%��V�5���>� ��/�ӑZ��s����[�� }t�;}�;�����u�r=ßV�Ҵ�#�1Ƣ:��Ф0��/��oƩ^��GV$��7�s!�5�]�'n�[qsv7�U\L�,:|h,;�N�]��r���t�e<�N�;�S�M�
b�;����݆�s����6RX��:LX��Ŵ�af��W�:7K�VP7���:�pe�n�0�ZĢAlmd�{rހL��̋f�"����9*�YP�^�l0�5I�zC�c����hgD�@ӕ��$�LE-�fI�s'^�a�{J��h��Bp����:뺕[�C\����
&_v�Tk�b�n"_(�uO���M���x�7��!Ў�+H����e�ܬ�D���a\�h�Ow%�!�z�J����r����Q,bKhs���qF�Ml9�yo������q�O��[ �\v`��b/Me54j��m�=��?,��6�~�gsã����{&�Y� �L�I�i�����*z;j��#��6�V,�]�o>�Oc�:_Ѧk۪v��d%\�˥P����\ ����e�ekG�G?Vz�K��6�>�$�V��}7�Q���lʺ�_�-F�V%	x_"��%�@��u�[\0Ww�>�r�yҔ%�i����M���X��m'��1\jy��ݧ�0Zs����1��ˉv<���gj��b
��1�ÀZ	�)C���m=9������b��$� ��8�� ��P~����f�����j��t��P�3�?f�=٘����m�,Y�5(��k"F�iT*vfw�L�^*m�b˟Z����yC�og*��F��|G�VOsQ���jbZu`�Ek�ө��HߙMfRW���
���o<C��G"�Ӽ��{�&Bf��>��e��X-�u(2�*5f�Q��v�����Kq_w�>�R�w��@�>��[�[L�ݛ
e��RX��V��4��2�z�����#o�{�ӃΪ@����ZC�~hM��J�Z��DV�X���������7+��U��X�L5�$
�{����s�]�]v��n.\KU�p�5uh��k��.YL�L�[�W}:骫���C�]lx���S���	p���P�9~b�YZ,�T#���·�����zw�ls@�MfS9��n>m(�d�OE��,io�\O�W�p���B	@m}	dXׇU����Z��4kOR�[��>oiӬ����<Q���w3�U�0�3�ͣ~쉯�`��xT���O�]
*k�T�ב%Y�x���VT8��mN �9>b��ݼ*B��3�Y�����AXͬ�:Q�ʪ�����Y�M_o��ϙ�0r�Y���湖'TJK]W�M���|A��
�[4�ѥ?Ϩ������"��P�w��V��~�ʝ�*Ξ�t��F�c��}K��a��>��"�jk2�h[����J5�����}
�co�z��v���i�K%8��Yk����g�!]\{-�XߵQ��O����6{1>u�q�S��N=3��)}�����֦6Q�kN�EF(I�KeX�zVX5N�0�8��V'^��l��dU<��z	<����vjy^������w:V����=F�t���_�}�6��&T�αʭ���V�sd��u1mO9�m����3������'O]�2��½C���=��t�s/}\��e�t:���=S�U�@�
Ʉ���[;�]|D�(�����/w��G���K�o�NtD�zq��_���z��U��޾���	���V��R��T��M�3�ؽ����k>�ĻЂ}f��.0�PA=7�@Ҩ�Kw1WWhѵ��"����il0��K�È0��!��[���X+c��1s�<q�xR��v w��s��͕�"&c��+�Z��3Zc��<��1�ʺ]��\��Zo� Tm��r�Rh�eT`%]yGm�5�-z�)S`�G�[.!�]����'F��Y3Ŵ=��q좢X�DRܶKq�Z*d��.���N��A�>�}^>��gl�3���9[��6�M:�I=S��c*Kb�F��>m���*[�U��C�C�
�;�5ۙ�9�:y��S/%A"���?��'��=h[G����)D��9�|�8�-�ֳi�n�{�`$Gݻځ}��w������zk����T�[ekd�0;v���Ub��,�ԕ:Q��
�cuM��Ѧ��&���os���5�SCvHbu�|L���+�vU*���3.Z2�V+�^,��f���{W�ʯx��y���LM̗+�9�ĺ���\�C3Z�.��eC]N�X��B0��UҘ��נ�Է��Ǹ�=y��j�O}�>۲+p7t[�����;�x���.�=�Q��g�U����x�L�kv�^l�fQ���=PT���M��\�R�d�T�yKH�P�}t�Cb�y W����S�\�w�L�\����|��23l��Mr��7��j����:<�I��w׾:��o��>���-{W����wL;�,}�s��ӧ����nҫq�G��z�ݮ�{�/���iJ&�z3-��Y�6�����Fӱ#=t7��} �*���D��w�}�Y�j1�-a46�	E$��)յ�kR6|��}8�f�;&�2d����1?zl�F�	���S,tn�9Ċ�`oM6r��&Rh�*&-!TS��xB�3����i���ƨC0�J����֘��^��ܝ�k�y�7��w�����/�ڣ�9-��seTwh�[���m8G�j��NZ�{E����q��̨H:��0��+c�F�ax˛zPr]��u]T��8Ȳ�3��'
�I��~L���h�����"/����v�����9
�n�ڵ̱Z�2]R\�2�J�c�t9�/�S�-�'���OH�]j#�L��x�]X�V�ʚͅ�Z���WM�
�1ݪ�S30����Dj��J�u!Q���*�sc�D5)L�>��v)�ңӯb���Kv�؞�b�Z�i�#�����6�d\u��L6l�����9�KOy��Ŷ�Z��ځ5Qֶ/t)'f%���'MkH����T�.����'Z�]Dܚ�۝L�̬^��wM\K5���j��Ȗ��	d�b.+���T@���
�z���1N��`�,�g�RЮ���6���4۪v�e2	�ڔ�-����u�+TaMB/��6��P���E��UM�Ƴ��VV��V�m�0��GSa��m}Ժ#��?��r�w��{x�I�rά�T��;&�¨���Y�6�]�ao��w巳����>U~>��$f�-4�U��͖���N��Z���H���d�*�s3)eɼ�&��MV��ߒ�D��3>��l-ưZ6Υ)#L�T�=q�Y��ؗ;��h�3�z/�JT��͍�u���yb[j�I��qƦ�	�:�'���cnO}��@ �lδ�4e�-&A��U�CĀ^��v�^�i�wA�.���
e�4%բ�D�eԼA�2iT�Ά����R��B!��o���w�ʆ��Ed5'$Wd��y��̕��o++Ta�e�+3���Q�>	���Hԑ����5O+s�2CՇJ\�B�r(�2�����p�1��#�7�Q�3Z��>�䲽9AZT͂ܟi{l��3�e�iY'"Ԫ���g�8 E�����bk�V�ϙL�^B�I��lbX���4�N��v��zX@�W����ӊ�D��
�}ehZ�Q`Ù��jֹ�M�ul�Fe�+�����i��3V�3�(�Ak�B��K|����k��ov�3D���|��Ut�>8y�[�5�U�<W��uL�lF�܇֦ZgX]N1���^���B��L��Q�i[�k_��w!�tу�gT�&���@}���׊ǉ���3��|�1�s�Y�ҋ۸5��A�9���jQ�&gS"�m&@����\�TJ��m�3�	9_��{�ݿlO���@��J�=�Z�eH|�{���o��ʞ�_w����h*>�|/�
r�,�{��e�3p]b�+{��ꕅ�|%b�-��+=�T��<Ew���37;1�8�+��(�q]�҈jx;��r�~U�>"�>@�׮�)ׁB�~H��{57�4a�쮱�Ӎ�a�5��:B�b�v��];�y���f`�9� ˺��o��1C�A,�ʎ��N���y7s�tq�ݙՂ���p�V����Jw}(�Xzwk���{��{9Qè��,�Xz���թ�Tp���	�rZI��+u]��>ϗ�s��Ê��UK���/��*���s
��r
_-l�L����)J�*��86�:�ǜo4}ꝃ�x�+[*Nz_u'v�&c��I-��VP7��w�4뾾4��8\�{����%�)��k��2\-D4�YJ閺7Mi�$U���c������}4�n�/9��'�ҙ�"OS7	WH�;m��e����R�`�D���D�$�R�U��x�aL<��<��K��e%����--ǖV�S%��R�'v�rZ��}��0��<�>QNr=[��6�M3:�JnK�Ǽ�h�ݾ����L��m:�|��U��i�ޅQ绕}����􂞶�~��S캘�M���zN��[AT�LR�mv_%��ߏ��W�Ζ�$��/��Y{��8	#��u��Q��8i�/��_l"�h�^������^KT�����<{������5��j�Hqe ~�#�;��U��[e�u��Iw)��ة�f2c��V�ok�`�����+4Ϗh��� ���d�)�F��6��dJ��+���|�&K�e}�6�3+J�-\�m�z�*8��D�30_^�W2����h��"��${A�c�3Z��t�q(-�ڸ�[��-m1���x���W����9����/)�����H U�A:`��s����E^ޑÅ���c��i����W\+�:)@1r0v�zL݆�AX��fuH]��͍JXUٝ�:��+��#xuܝ.���;���!�Pœ���$Ji���О١ke%ە9�
i�O!����y�:������i˛P��`ż���gCL-M`M}]P���I��G�*㱽&�yXҩb�ARS=<iX�H�+zqc��,@�Y/uQH�&]K5�[���yݴ��<:�7}�
_E����.ۮ�yJ��(��˨1�� ���,69Y��5�w5��Ƅ�����RQ�++fW	�ҸX�J���82-f��]]��>����OTY�W��nWm��)[���R���'j[����$f �G��wzO2����R�F,�Z9v=ʔ���-n�>�����(3P.���ء|l	0l�8��4�>�y㓳aI��W��)��Ww{x���$+.��T�������6���l4������˝[�;-���逸���Pr�[Y����:�@�0�pɧ�h�n�&>;��! �uu-�`1-�yx�S�U�v'�I�@��Z̠vۭ�w&���������&���8�9�29[�t��tN�t9ҳ�7����8�c�ޖk2�gű%�o�.�/��1٧�;�,اv�o�JY�k�),�9���[yT�Oi����T��:��!@Y�n�Ri�,�$���`{��|�s܇=ԫ+J�&f��4a���w�@���Gs&QU;z���4s��5�̗�5)�.9��o;�..���� �X{Ȝ�r#�5+������ٵ��n˕.�p�av>�Q�Rdo�l��-��O6b�������N/��n��]�-�yg5�]��<X��:�)a�3uc��^�F'�Q�3M0�t���D�fw�W���[��2]�������"��+:_H٤�9���jd��.�L�͹u0U��0E�tWԳ*5I͎՚�c����[/F�jLurA��g*�O=��:�兛�:](9���e0����`�F�d���&bI���F����{�:��\����ѭчn����6�l�Vz3�JK�z�1��j�Q�q�kB�[Χ�Y�%AbR�1t�^�ݳ8�m�]r�a�}���Z��AX��#�X��vP���ӨKSOz��9di��>��F��}JRD��	24����L��J(�1�@(0Q�Ha��$2b�&0a��h�B4�2Q���)JP��́�iP0�RHQ3!R��Q���Q��Cd�,C$�%64d��C1̋&ѱF���X�4��L$�D�Y"Pӻ�Q��$HX��)���D"$���a#D�\��,��DI�
�6�#�$`I)dS�#R02E��ِ�0�Ғ!L�)���� �R����_Nue���(��v�WS&h�ΠÛϖ�ph�}���Y��(�&��K�w2�]gQ��6>V'TR�'*rަX�ސ5�KS��Z�-��543j�항��2�Uy3�J$f�sɛ���z��e�r��4٪D���^�V��-�5��Ħ����=;�vv�fJ�޽�}~��Y��L�6�-���	er�)��fur�XfY�콛Վz�YE��.��ҳ<���h�w�5���`u���|x ��/��[ig�D��%U��#��^
��vf*.}�e���Z�!CP!؆�e�Vꄧl�*�k�}5��cΞS�^wC K(��G����6q��Lww<��'R6ڛAh:���6����h�mM>뙯�>����G�nOi�ofS��gz��&��kf�!(I,,�V���H�TӮ�l�ٶ��Qװy����2��������LN�J��:7K�E[��Zȷy�'b�z�A�
X�;DI��=��F�Cԩ�tr�9�p�´A�K\$����Ԭ܃���2�8��b�S�֕%��OH��Z�:��޶�Z՛�P��C��	�.y#�B�&Q�j��ư���8�.�+f�@oϗ���ݕo�4D�2��f������H�F�O��Jc���^�A*o_K��;,$F���y~u�N!�rZNfҸ�N��Qk ��Q�p����"� i�S�ϕ�r�dĲP�[��E1��Q�އ>�{�z<tZ�0a����R�)R�ߝe��H\��Q'��Q�V��]h~~���lg���UQ�z��6��i�k�-u^B˚d-����r�NN�{�9��a6��x�ڷ"a���{�ωىbJuL�lE鬦����YT��c;�g5�C��mv_&����'�n7�m&D��d%�M�6NV;�P�C����3R�旰��{U8օ�RB��4YXn�hܞs�+20��"�n��/pD�>�r��񙾨R�P�~�BN_U�C�97�:�W3�������RxC���o��B^��t(XǙ��l=٘�����U�l����g�1�u�}��1N�޾�*m��eͪ��+e0TNT�I�U*���
�
H��D8U�v�yE�(�}�k�{�{Ѓ�->�D�!G���d��LWr�ih����YΝ�X9Ҩ)K��G��T���
Lj��h���sP��y3>0.��N�&Xx��.v�qNٝ�3�{�n�~���L��F���>:Z�2�oP�Ӯ��6����5�L�^�Z9���Fk�m�Q#n�N&M�P��q�}6}��[�`�m�J-�$i���F�,uTd�9Y��7��� ��3�Z�kyU���-�}cvl)��}Id�X��S5��[��z���~�]�Y읢�o� ��yiN@Zi��Y/�q�ah�u{�b�R&�'suɺ-���NPV�=9�>���׶tM��δ�WF�a��&�}�����V�16��j��.Y��5�B�O���l�V].rH���`���:�f�8��$M2�/�n<�B�ʉ`a�����U
��]Z�4U�t��v���z���n���k��Yyd�5�u͞��Of��k�u9luP��
����u�'�r�����2N��Ik�wm��̲����z��z�]����~N���zQ�iU[�k_��r偡]f �V/��E��WCyrC\8~gMn����;{gq�/�s���h�q��Y�����7�7<(uv%Z%�ne�y�ùG�,@+��o��߄�'n���˳_�x���� >��_)���{P�Y�*y��
�W�����0�f�Al:�1���JM�������|�U�mܴQ9�Y&���orRQ��ȑyIj����	��'�E�j��3~ھw����f!@eL^�6u>����1���M�*��,���Z�6мb����H�f�ھ�q��y�����zb���kMR���o�����o[���xa����=��V�~q�yT;��J�:���u���OU��t�zb��0�V��M��ɧ<XsLT�2W���%.��>��8��1Q��U��tu	l�q��#$^���+��Q�L���y��[�fg�]�C����G���;9���Lk���GoV�[(�0�Ki����͝�kӮ�1��i�{k���v��z�ō����L!>���th�c���Ҧ�ng�]�<��k�+l���޼y��N1�q,	WL���g�j~�y{��{!�5A�0��7N2d{�6O=�vy��7���W:���4�������^Vw�n�̂S5B)z�`0��N����CuξJ�ٳL(C|��ŉ��:�͜�6K��b�bQ�� ����6��}�{�=�7��S���|Ks����y��c����x��M/���Jw0��6����[���/=�@1$#�~�d��r"�0>�>F<��KC���+p҉#TmQ�P�n,÷��:���)[c(�9��s��lV�����9O{4K�Gn���I���</Z*'�-uL�ZuD[)��(�hs���0(Ya�ݡ懭���l,��{��7N�:�N'�&�LE�6&���J%�V���A	�Y{�C{' w|=�4��i��;)�!4�6����Y�J���y.��#t�.��y3�x��� OZ�U�f�>�7ͫ]�[��s�^*���^�'s%d���~��r���	tj�'/��U_AN�Ƴ��v��7�
�����#ҧ�L��(�Q�kֲ劫��G2�����p�3�oWM�
C�nF罣3T�b�ң��U�{��WD�̡U>�;=٬�uW�!�ճ��d��.�9sP�(Ζ�<����Z�X�ϲ����j�oA"Ãv���p���Y��z5�j�E)6���(���T���H�����N��\:H�����L��V�>ֵA������#�v���wV�{�c���-�q��mө���5yIY�G#i����1�ϭԢf���ܙ���e��[,�e����o$��)մ�֤l#�aM&"�Bł�&�w)��3�f��A�L�`�t�Yc�u�q"��+
P�ǩɽ�m� �����v��CӜe�n�5B�T�����E�:�LB��li��~�.��?1�r����U�N#h��C������*j�!�"ޖ�9XTރ:=���᫒�W3��}ֆ|ӱ�Y�
��-2��^�4�%�X��IB�u��䐹�P�9����+fd�����2=��x>���J�n����9�:�2]S2\���*���3D�.<�Ow����o��r'�v�l�k�X���S�A6*���/��̏ ���:�cԮ�z�^qU��>K���AW�n<ۊ֓}E2��*p���t�h�%�E�Ţ%+δ�;���GzuDkGNq7�.�oi�Z��l�p�ޛ^`7�ݍ�>�������0>-dO�`G��bȴ���n�fn��" ���c���ʖ�ݽ�0΍��^�U����hΏ�ҙ��� r��	����Ь}ꕼ�ھ�#�W���<�u}Z���m�aq(V�k�z�*���}\Uz%L�d�SX��ϭKo�ve�)\����^�Z���Ԥ�6"a{6J�S�Z�7�q�J�G��߶����p�n�~"��
�u�KeZ�f=�k��Uᱥ���{;��k��U��/+��{VI���2{T`J�=J�:^�3՗:g����Hߔ�e2W�oGA2%��Q|�Kf떗��SO���8���;any���:�\����"t��.�}M����A�1���wv�t���g:GѮ�ʴH�y7�W���&7�`���w"���`�2�]�cZe�-i�y��|��.M壹k��^ĕ��G*��zq�%�-���L0�����U��n���3��Cg_T�q�L�*�v�16��bk��-D��>�!ldXW�\�A����8D��)/{1s�ɷ(�f��b��N]3{��4`Nw�w��F�~�)ʺ޾�yAOm��'�`�uN\*�w-��k�C�R�t�����=�.��;�{�a&Ҁ%~}���"d��ܝ�B	�gw���_rx9�o�rTt�
[��ǻ�{4u
�)��uC�Պ�$M!Xp���h\�)�V�*6���JoZ���}0�����y���^s�[��D� ��!e�Z\��y=�u�{��F�{U�� ���v�:]��Vw��9�O'y]�J#-����)��_Qة��*S�x�(�hu��|�.U�nu֕uJ6�͐n�L�Aǉ�Ӧf����$ب���[Gݞ����ʌ�S�e_B�x��nw��Y�Y�3l�!,�0�J/Tg�PޚV�]X<���2{#�zo��n�h˹�os�F&�n�ʲ�5�Cj�d�UqSg�gs���͈Z���0;w��G&�͖R���8�J�Kaf���·r�k]&w�^ͫ���v�Z�9�X�]���~��3==S�	O���ƹl��,��u��Y�y���&OlU��f|�G<�na��z-�E�V�T|��^��-���y�ݘ�T�wi�WB���]x?�C7����yowo	�6�:�f���m&7/������N�T���O.Z�8�)(��fIt�������<	W]��s�󺶦}ը����tC���Y���gU�J�(szQ�oz�Z�ݑ�����N�)dsq
�B'i����6e�����}�v<�G�7��+@�=w쓇FEb�;XM�AQ�%��Emx����c]�<1������кH��Dq^�2*&Ob��z�W^Z��yc��H�sIk`�"�+��CYw�~� �F�и����]}p��m�bk٥�lH����>��eh��PY�+�-����h|�%��RI����i���U��[��������2� ��glbZ|�qE9ͼr��A�/d�Y�)��T��d�)�������'G����i�މ���t%<%%0�1�NI�_��s,�j�Ik���Q��Ryc�]�����(�5�j�ZfԼV�&�ˋUY�Ӳ'Ĕ�X�؋�^&��*TCq'5�lS�� ��귄7�;�]oi��vS�Agz�w�A��;��Elߴ��
��M��ےؔ$2><�RG�辺��Yk:�ް�T��a����#������l�p��#��E�ƻ��X��|��N(6�V[��=]I�+���!ٹ1ż�x���S�ޫe�+(M��MH��0�s�u��j`t�(��N�_R�U���6�v(7r��V���5�k�e2�;�N��82S^�;��4\+�O�XV��o�-|�S�I.�t�^�Q�KY�.�.|�}.ݺuNm�N�M��tX��c���g�P��x7���L��$e�)�6�=C�o֩+%��=��p+�5�u�o������hQ%{h]8�ꆼ�W�����kPe{ѨfRX1���T���ͥ�����N������T�,OQ��p���Ϋ���A�g-�"^�'���)v�ck�͛�%L��~�<�!zi�$S4�:?����!��=А��T���(�ɶ�ڟ�$C�q\�g7zn}{�,D6�#W�t�J<���ҝ:���V��׎C-�d:�\᠊�����w�{��q��:�6:Ju�p8j �Ck<2ʚD$+�\�w-�qy=ui����]��������0�L����D`
�C���5ݒ�zg�HT�!h����>��w[YFf^v`U�_4�r��}|�n�{��+�i	�q�3���!�Y(g�x�\suܵ=�@w~,�t�� �\�^,��h���L��;�}X�Un�+-�	k��צ+��I��>Z�F��G'��7eEF�iPl��E���+|�/�$!�4f����`���NN����=?GX�Bsߺ���:	��
���9�=��g_TYI�Q՝�pi���8�W�qK׍Y���hR���K�c/�OYIV���b^G;ql�Z���z��5���U*Kz�kp�	��*hY{��|+ ��ͺ��c7��j�X]��Xg��-�49j֣G/k%�Z%����CO��3����>ټ�L�y9�s��62�V��C�c���j�c��\&�U�Qs�X�޻�oc�xf�ؤ��g.S��5)���u���7�:陯�y�	%��'�ۥ���R�t�v�r�:MհV-����ިD�Om��F��΅v7���H�P��4���v��7ϦV�E�+uuH	G��«=�3\�#@�-
��w[B�(�C���a�ꮻ���=~z��M�Y�R��Z@t�_l�sb������LR�e;,�l��t6��-e���BTf��>n�
0�����7����g�U�Ǐz�b��2�Bj���b���t ���wvզ.p룦抳��wf������hԽڙ���g|�B*ɝ��PtdfR��чx(�zŲ�+p��<���nVg�Fs#ol���V�>����I$|�F"�7�%�t�[�L�%�/D�%[
�:=:�h�!����p�/�L��`a�3�M]�GC�δ���)n+1,u%Ҷ�l�6@�u��'��v�Ne[]�n��4����	8��^MHwK�$�$B]��{���G{Sxn+�fPN�1� �F�M��x�=Q���z���1�-�f�
����otD�F9J."�2֫4D�9KzF]"$�W,�Q
]i�o]΁<� iZYM���G�8wن�YB]yR����SVS���]��{�[&
yr[A$�m;�T{.���h���L륳5v\�*w���]��������νE̬�;�t�S;��J�b:��������剟]�K����]΁���<�&��X̀�][�]D7�Sp�Kx:�x���i��7,��Gҥ�f�����n��@�6�s����a[�&�ɺ;��K-�*ݝw���8�Gέ�ܮF�|�c�s2�œEGX{���|U��s��$U�g`��3��l֠�+���w\Dps
�L�7�b���vu���mΎ�jY�9���u�D�MK �{V-� u#�-И��o����=�Eu�<(��omq��BY�m�t�vU�1�����u}�ٵA�{�u�ݖ�����p���n^��I�r�
ܵ�0Z�@QMW {Q����Z ct�ݫz�$�E��)�2rV&�����r�ƋQe��}-P�V�8(���ˑuh�8b�B�Wr
�ɼw.���۹'/�G�}B�P���
fe%�I���CE��l�F �#&�b�ȥ��В��3�ff�*JP���2Sf&@d%�L����%��(�bI�@P��F
 bQ����PI&$�61l&�2Fō�Q�	�1�f�4Ғ 1�D�h�"�wnPPE��I�$4L��s���h����2b"4P�lF�F�����U	dō#%%�&X�	~}�z�?�=}�8mcw�u��G�Հoh��_M��T��^����}3~����������"�����3�D���^F@�NF���2͝~�B�H7
������������B�Q����g|����1�1�ɇ�w<�r�^�*��NmE�N��8��}�|%��W_SL��.4��{����6b�-��4�!����8MC��H�K�$�����\
�\�*$nsr�`kx~iw�Ʃg�J�^���)�v+��Gx�6�`�;�\��)��]��\j��*u�/���{�uǫ]�u��|�o6S<��#e�~�~.)�Yy]����W�u�kw�;�=s7&c�<#"fg��.�"�����+���vۺ���K�ESoK�!�s�|�uM7<�gw%��Cu� �,�Q)��P9�-Օ���J�֗4��x߾�~O��������կ�(�&q�h���^zc$kק����ᮻm��A���.�@��w�,1l�ʝ��ڝ�Yʎ^k�-p�뗌!=M��P��!;�YT\=A���jg��c7T��hAW�-Ԉl����r|���ۻ��O!��Cz�2�y-%t;��ZO����N�o��н^���z�r��Hg����#�厖�������3$���)��c����A��fc��j��k�f!-HDŏ��<�ν�_��=��Ƥǉ�k�	wJ�˨v��vtG�`�;�Qq�ʾ͗��gW:i@�1ģ��a���\ٯ�ե��W˹�|�h*՝�onb�Z0�c�B#��Us�7t^���9�@o�"%�A�T�#�����sϙXR��Ր��)�6���5S�����󩻌\�}�YEָ���?e^i�J�eqR�td\�̒�sX���q���q:'OX���͝��a�[c�8u���R`�S�wSKc5���W��8�؞h�����C@�
�[�hJ���%�H�m�|����+��\����vKp��}���xnwS��vy
16�>�����T��/k�sˤ��Φ�3dL�r����ݚkC��/4t#	l��þ<��}`�l��Ϭ�ç�+�'���k?1��1P��V���wX�:���u�E*i��%��v���|v/"Y�����X�ye�t�����q�=��ة�a��8�n��l�㼮���o���؟��u��A�)yoz�S��r��H�f�c�� �ܶ�f`w�A� WwK���!2�M�/����(��b߭�Ү�I~����O�8��敲^p�j镳i�4t���0���/����e��=gT�)���$�k���Y�v���a�
U�y�'Kk�-c��s�����̮�������2"�k�Mj�>�[�&�,P7�p���m���[9ڥwo3�)�U��îdԟZIM� ����+��
`�������$�����;�lj{���үa���p�Ⱦc�ϲ_��=zT`M�_��*���=���]/���t�`[A��v�s&�l����=:;�`�B��=���_�����X� ��k�|��J{z9rr�fu�mvr\���ę�Ok���]���W2���v�Cu����m+%��k\��ս�=b��VV�+��|,&��fy��wd�6ǲ��g)�6�y\�QB��M������i�~dD�P1]W���Z��R�,���"�*Y mWSf�r�OY�vA{f� 1	̳�k�OЙ�sKu���w��a��`���yc���}���*n.�ȴ7!:�:�G4A�{���̨}n.��0�x�c����+غ���J|�퐆�w*n�
s�u'�}�8�8��对��k1���,Dc�3����! =���˄�m��O sz_�i�bY�N&^8�̍m1�ђ���T�mg������)�2���-;	/���C�`g4�.�6�L�D �����+��i����t@��A��C�蠔���i���״�_l��п&�{M@��M�o}��cB�	1�Sc��g/	�t�L5�ݜ��ʺ:ek�������w�9�"�N��n�efV�h�^Q����.����-]]A���!���_���{�/:x��ƛ�S0��czy�j�19u�h��++gm>Zs2��t�zv�c���]H��K}���`H!qn9���޽�7�B�>��P�ˠ�����ꎳxh�Relc�|��s^[��]"��8���#8�!8�,�o�u#@t]��fؒ���������~���^�`��l��sza�j�52K�@�]ϼ��7��;�у[��8�1�]�N-
�s�E��k�r���Md'�c�V����9k]/��;�LE��#]R����+Z,���+ښ�?�TA���x�����?#��V.|yf˫���L��U�u��Z�mA/�9Ў�4�;�%��^\�� d��~!�!����!`+��m�&Cr��3v���٘���b�]<��z#�3o�V��ޥh��,s��P��~�IY�����dNUu�F�(��p�xk\i��I��E����9�o���1��D`��of/�I3N/:�rFuC�>v���Hצi0�b�'s���؞���.��W���o�Ո5g-� w]��eͥ��kw2k�4t���=s��^�1E4�tdK�`T�������o�K�IA��妚Ч�) }�p��ܿZ>��Β�kEe���?Jw��A'Pd܆Ҿ�VЊov�'��AА�d倡V���뫨7�5�������q�l�M���y���U�k%\��=��H���g2�r�t�a��d|0�UߥWv�O4���/���?(��R�9V��]:�h�~���k�iƛ}�xi_r����j�s��d�W�$!H9����n�Gq,�5��uRh�e��qۨ�y��Z�22�'��J(��wXv��]U���# T��ʉ����K<��ܪ�^�gT�6� �F�P�˖�h=D�p8w@�i�:�򺦐��;�@;�^�S��s�Jstx�D�I�`�?8��כ�Nl뫅Ԑkf轮A�e����ѕ�U�^��A�b1A��:<Y��z��$�����?�~;�@s��!�[<�������p��t�vdΗ��w�g:Yf�4���ى2(��O����)�#�5���̈́�:z�$j��Q�swP����{�i�e������M����t�,U�H� !�a��`��NC+�{+��X�mj�=�5��x�]��μLv�:��`�N�2/���g[�DF˒���/ּ��du����˴dF�8��&�A͑�����/��Q��nʞy���c��U�.���#-L0���k���/�5jci��x-�士^�S��x�#EF�^E��18��Dj�-� B�����z��fU�ʔ���e>�l=�|�r_&��L�Ibe�!�H���$�^1��4Y]%�k�+,Z�U܌��*J��5V�}�Ѩ�&���D���;�����D1T���s��c��~�?SR�P����:���6t�<��}Oo� �Ͼ��C=nj��r��_��y�1���8>��xf��NL�t��'����n��Z�gvn��u[^c�'Kˌ���������?*�d��w�M���ʢ����gQ���_g*��n�9*���:^�rY<��l�)��ݒ�_��Yy-%�C�l�O�k�{ɱ��季o�[:�eArTκ}�t_�dÓ� "},����EHL��<�V(ɸ�n#.���Ժ�!M=�B�l�n���y��eW�0L�� Ϣ5���YT��m��$뾯�7��4���~cq(MbU�8��`Y��mve�ç8u�p�gw*�?�F�P��NL�����W�ԡ�b;�-Z�y�J���YԈ��|����+��\����[���C�Y�-�� ������;���%�>����	/��{\����
[u�_v���8ؼc�C��I���M5�1!
b���þ��-`�~xdl�C��+�'�jPH9��˷)�R�'�Sܖ��� �hk0H-p�8�vWI3���v�s5������K��ݪi���^����{�3�t�z��*��8����L;�u�iox��S�����A(��h<;�ۓ�ad�x�Ŋ�-qym�Nr�;:��A6k�]D���;�x�|	�yc���z�Oܒ���w|(�^D?aJ�7x�X�8�5��̩�7i9ed&��3/�<�ʺE2����9<[�]u�)����Q�b�6)�жq�&R��wh��Uo�h�.G�1T2�&�Y��@��w�O���/��E?B��T�|�"���c��XS�'�{���<�^l��8j���4t��1)����2�9�*6׆9_�_��鮔˹>G�w�ŀ������m�����m?t>tvBwJ�̣X�x���6�1l����E��Ry�`����L�v7J��#�qx�)�ᮻi=����(�Ѹ�&����y�;�Y��!�61
}�WR��`��״ �:K\��w��b�Y�=�ߘ����ލ3�ۦy��]�\��.[=����缈��e��҉鎃,��-D�ff0t�������y�*O��,�6���oܲ��Ay� ���o����2�fƞ�7��y�"�4�pGX�ώ*�:E�tw~�T�m��"��bc�;
�6DT��4����a�3HU��X��3׈.�)��Wwǌ��C�":fpm�Fs5���l@ &��)�,
�m�o���_kx��}1��������:�*h��ڝD�����S[�篾�ک�*���I�ޗP��J0�
}�y<.a���O��L�*.�K����Ϗ|_�>_l�7�Kv%���Pәr��+6j��γ�����@���H��! =�V�^�.�~W����ҫ��T�f��FF&t��Ϣy��^0QU��z2G
��T���x`����<!����i�ب��:�R0�0����+�\�����M����UI滦GE ���@}�3��-:8l�F�fS].�۵fQ�u��6���+� �t^�����wt�t���B�=x�b�w�ɹ'z3f��<闛�Ǟi�����F��ydQ��Y���-�#8�'�t� �*:F����6�Mgv�+�h��6D�FƑ/S�pNb��/j�2K�@,�9�=\&�K)E�Z�k�2<�����2�x�0�V=ʎ�5��'�j���i�zk]/�
-��b�N�5�@-]�{��ӂ��6K>�� ��2���`eM=9���?�j���8�;v���~��8��	��T9ݓOӱ}�/�z��NS�I����*���GXY�U�_��KI���u����f���-�?� ��Y�L��Bj��bX��7�>x�Esp�?7Ҭ����V	��w��ZDNԩ���R	Ú��lP2U��Nsf��{ݟ�Wr�������g��z�r�	�뀹�����v:�v�ȫ6��e�x���zd�J��ЦV�~Jy�����<��ǥښyKM���-�~�`�kٵ��<v���b��ׂ0�	��2ݪbO{�Ө[.�l�پ�\ƾ�[1�C'|�ia�7v�6�%R�e����'U錑������}�S<��x3ߡuw��WM�m�X�CTnn*c_��8�q�K���PgI���<��8~3~k����¦w8�O<���`�����MF�?n-�����"�7y%�.� ���O~��Ezf9ʿ+�t��wU�����ӆc{8�͚E�{��W.��iu'�k_�G�c���7J#����+e���E�=�G�U�E�G4r�#�Q�:]֎���]U�ע0L��ʉh�t��X�4��&&�?V��9�F�����i�J��/�э��Ψ|���&���.8S&BU��h~OĨ��왰�s�h�g�qh�<ߜ-sg]\.��_�/k��Ѹy���3�g����/�*��7/(���^��G)�����g�K�J�������3Νtq��ۢ/��!��,�] ���(���T����Z�j�L�JS7�;���Vf�;wt�Jo�#���oa�=� v��ev�}�.X�{+�sO���j�T��r�5���] �N��Z��8�\	g
�������l]*TC���*#���]IF��"�%M�`rl,K���~��i0 ��1���j����M!���O��MC��H�K������)��1��I͒�����w޶�-n���_o�|�m =��d�M��\.u�Y`������X窩�z��33���M@��~��us��N!�7�)�O-�X����|�&�k��zA�Ny��N�J*�sc��WL�S:-t;��S�;m�R�G��"����㜋]��U��s�gZͣO�_y�g*c�����-'�5��;��y��_M>����<"�y����g3U����]�r�1�
�o�=�d'x��Opd�g�B��-�tO.��㫥;��\�/B���J�W�?�`���Ϟ0��7��C��N�T���ǭ�2�&�c\�u�VA.�Î(��T��e�%�9mI�,i�C+6GD���l�~s:��{��w��j������gyD�G?�T_��4+����jߪ �h�aYSH�"و;��,-��r�L���>T5��KG]`駯�Gu�gSw��SϷ(��h�S(. 2ވ�s�h�V��p���.heݝ�4�t�	E
����v��}\�R���3��`I�N�E��o���y�u5<z�X��*�wV�;�n�n�slɳ��G���d��[���:��5��Cx0a�R_$�?� ������ie%u%�^Kr����˷RQ����u,�L�Y���P���\������h��tiH������ӌ�����ü��*U(C3N�ܨ\CC��W��@%��d�x�v��6�8<=�J�_u�0���%4�+7&IZq��N�=��Um�ث��QL����O���;��yc/7�C NguRI������b��]�Ŷ�K�mNW�ʼ�*Ng��2��hr���tr'A��ٮ��`�a�ח���Z���xaQ�ˇj�T��<|�o+���8��j�{�|���(�;��7(p�4VQ��C���Ԉ�����9.�ݒ�\� O�+~;��o���jS?�ˡf�"���]'7��=L]��ʻn��`����څjd�$3�WK掰��	mn��׸څ7�V���5,ܢ��i6�F�ǡ���r�jV�ssy,�����QӨ�d�2��E��%�v���Ռ�۩7�]ؽ�qH��shFf���)�F����۠p��)˾�tt�2��c�К�d��
P�^�!�����BL15�j��=���y�k{3X�Ƕ�nwΔ��J˨`�]�#��W��e�*^}�&���j
�`���uw�1A��2�V���3E�,Fp�}��z�s7U�{l�2��PWթG�}]�U�����҄1�>C�����HV��,2�^�ߖ3��Q��{'|�fZ]�a8vf���u�_rw�i��X\J}���3����ܤ��>C,VG;�OP����]j#x�ӳ4�P"�!���;��#(�T�����fF���v��!��:_-�U�̳��u�(�o��'R2u�j󛾡2�£�8mk"������:�D�,oi�����\����s�e-խ��k*����Fâ\r������sk7���C��q����^du����;P>�]�i�����0��!�����soz�Sz""�0\Nj���c��y��)��N�s�����%�$X�}hmKQ�ʮ�$��z��˝��ѵa���w|��A<�]]��r��sF��m�S�ҠkU;���Iw`W}�6��KD�'V��U�#���Nˬ�s�*7���=��]pHʁ#��glƱh�Ѽ�b��Smi���(e��8�p�����̲��������h¦`t�djnWN���i�=Y��hF��kZ�4N���
�#oC�]�=pޜ��y�i���݊7vg}�	M�m�wY��;�0EcP�;��G�Xu.ƍ���0-er�Y����������G���F�fZ���� l�(��e;4��/.D�3z���z����_�_����	�DD�� 2�����hM�ب�RFb�_��@�"�)�B$���I����Vh�0Bf[��Cy�2%��� ���� g9&���FE$��LRFiw\�A@�g���dlXK `��VBC$X6aD�ᔘ�2Z"5��bCR�Dm�҈���PY6�����G8�0�v�܎�sD(�@Dx����^;6)7.W.�Pf@'u�$�)��p���3�̒���pd|��C��a�I>�.l�&��1�Ã|��wV�e��+��9M�zF�N�l�v�m��h왒�sW�1!�<5\JX�vn08-���a�[l:s�[6��]e�C�V#/��K��wS�a��p\K3�T5zb
�V�j����gR#=���gSF+��
Ռ�:L� �����6{�d�;�Z��$���~p�e�uk��4w*O}�Ϥ�qgj��3���k�Q�v���4�(�����<;�ǁ��r׆F}gn:F�"#�$Q�[SE����~1��w9O���yc���^�]Qm�i,��Ȕv�����4�iFg�5V�����%�zA�wIq����P�w��\��U�?lA�2%�;���+��KSsy����zctd���-�r���*�֠�+���y<C�oK�y=6�*3n�{#L�4��ۯ2+���ȧ�e=�Z�U셂p��+m=TC^.i�ݑ���R�E�Ԫ�!�f�h�������� }�&��8�`��Q�ed鬪�Ol��m��.�އ�j�T������)��Ya=�TS{`�f!����n�T����r��;�T�'�'S�N��:�6#.�����6�c+�Av��J�����gm����;�)]�Q-r�D����{Z�*��M�� MH\̡���w4�^M��Rt�.iA	�-e0��
�԰���lwwS���Os�.�M�ipfa
��]Ե��s�w�eA����(aa1�n;��j�f���1�}��Z�W)�偙LCz���n�����o>��t�E�8;�a�A�IA�L��1��K�=�^�9N�6ԧ '�h����=�]ڈ��앳Ry���=HsH�}"�s9�
]�RxE��d��*�l�WI�g)���4�̹�]��X��͙M��Ny�� L4pr�{p4����P�H���c��i
p������k�Z 5�qk�Oe�Ր)��wg$s����3T](�QM�����J|��of��g��8ޕN&a��xx6��9��#��Ũ�}��Z�yp�M��-�~�t��#��Z)������7d��̺���FH�L���"Y�R�>�3��ȋ�Mmrّ��c��DW4�r���Q�a��vt��{��<׻�GE ���|�t���unD*B޶v+�(�8���xdD�ז�R	�E��qM�ծ��7�j�	��F�}���E�l����Yd[�Lr�l�9����������7
��w�x>&�~�˥	�̆'�� e)&ag �u��<���W�2��K&OF.��PYʻ�pEȍKf,@v�[�o3i ��3��\G�y���]5��.\6;xeo2Q�/U)��`�Ǡ�&N��O���y�c����N�N��".��q䭥\��nV��r��:Q�؁�'��.i�'����B�9�0�3��.���9�z��rz�]V\��d�Z05��?4�3f��wި(?�{������;ڥ�����ڮ����OUC�kN�[�1n(BC���r�w���ӂ��%�w��L���`e�=9��B��~�O����Q8&�輬mZhFL����Fg����ݓOӱ~��-����^��g)���v��R��i�C���=R��̨�̵S<�zh����/�fV�iO>��x9�V�.E�w,s��QS����*zj�{��/��&tT���	�=g�7_�ozf�����-��o���-�ۡ��稾�'/9����-�Y�#]W��z��)�w3�S<�=G�=�WpY�+t��TUׄ���jw����ڔ.��b<���9�=���~6n�fΖw8�O<��3ܖ�s�	�����hWuO:6æ�n�%���7��{i�$Dr��Ժu7չU�_MN�JP&�#{_�x�}�mwR~�p�K�m!	�@�����dGq��O�19_Pޖ�d�|�Na�m�]M{aw��U2so�7�:}�z��[]��N���l�C����wLǢ�1	�d�t������ҭT�(��.�N���$�x�����U1.�)�*Fj���[����1���-�4f�B�Y���V+5��X���K���Z&Wp�(ŝ.�Ev��e�\��,���ʀ��b[s["��uK��̥
�����H�;E�YM!)$ +����{����p��I�^f��b}iwz�c���	ޙ\3�8=�^o��f����RA�V�A{ãp
��h�X�dIʡ�A�b�F�Xɳ]�?Q�b�l�~4�����Q�2�s�c�A�x�\��8��7���2E<ci���SȻ�x͢[��Z��fS�)�@tk��c�g�#�4�	���т�5G�<����Y5����F��܄N�.d)��W5�:�T����L����We|��j��7_��T?�{��A���P��T�wG5��~���|�C��l�s�B �S��n�pnO�䎣�&�kRgެ!h:5͍˫�D�΃��ߠW����w�M�ߕ�s*~Wc���5��,��������X�/��#_����𛜖FO`kK�w��L�����{�k06[�>�}��Y?p~l�9��s�U���e��qx#������m2}h2U��.�@a�~V�Q��ѿtyn��O>�S7\˽y�q�� ���fU����z�W[f`bΎ������v�]�)Gl��ǯ��l�\ɔ�y�{Şn�|�͊o�o.��s���[¥�`ˀ�gX�,#VX��6�me�F�s��� ��WՇdQъ7}:��q��o��Q�qu��NX�~����X]�ަ/N{UzT;��eIp��ӽFݪv��sYlL&3y�b0T�>`�n�������A�$7P���,�����w���Ly$�;��$Z�;�����\�)w��%tNWO?.�/Ϧ�z�rڇ6� @tE��,�����NB����E���{摬�F�m�K���Φ�1��B�.�ŀ�̠� �J�Y�ү;/�ʇ���װ� �1�P�+�Bk��~���y��m{��-�9Ä�U1(��R�6uϧ�Ďd���w�sĳ�J� ���+S�5	Q|t��h[��6�7����q/{�ƠL��h�365���OxC��8H;��<bm��}��Z���ܩ8/j�ɘ�ؑ�<�/v@�7��f='@�Φ��]M5
$!D;:3�}w=�`�o��s�ctf�΅�]�0��y~�r����@������w�t�[J���� E �lt�j�G�oF�lD���,����Rۢ|t��RF�Ewt�l�'��z�	�y]u�Et�g�@���aLQKii���J�?����`�V(oOYg>�xj>�=�U���g���ȉ��B3�u/�c�u_+SF��l_]qB�AE!�[��E��9�� $�3�F�*�1ݷ����n����hN�^���s�d2��Ç��m�mv��i�����H���1>��VR��V��)��]���L�V�#�A�&+�"U����!��qy��b�����M=��4�᫦W�=TC_�sO@�n��x����ʆd�m�{u��4?'�mR�)�@ ϙ��dc���`Ǆ0�d��eU�{�3�m,��̢��;�]�m���;�{Q��D��u4�]w*��� ]����ct���%�E�w	��5Qp���tft�mLN���S�9�OoE���1����Yו/�рfkn�,0�(��ì���"ç};��d���	�w~k\h=4'��)�|F3˲K�=�^�9N�7�S����a\K�v��Kb�g:Q��}�i�iɔ*Bg�)�g3�
]�RxE�T�@��k�喞���vA{�1e���*�1�z�Es&��^��#\��q���Tc�p)g����}���*n*�WT#
gj�蓝��;�H�����F�"5�<�OM0d�@�iD���.�|{f��)�F��j������:Y��?ͫi�߂���m���}���xg7A���TF�����Oמ��7�H[�������������](W��Iqs�ڶ 	����V�����x!�4������N�NK9�_.%�q*�ٛd;}�eǑ��1��8����ux�]�,�e�'X缹�ݧ)��LT��@[ݣ���y.�ԙ�C'dި���ۙ�*��D��&E�D�/̖O sz_���t��h��9[����)w��W��+�ZD�Lf�6�@���ٴ�M���Qs�nwI}���zfS����D����@�FS�Po��殖�	��0y��]��xe�Y�k�*b��h�2-�y���ߢ+��B�8�4.�~B�i�-Z̙������ D$|+E��8\%�k�*(�H���n����V��v}>^l3�b��5��l͊�#@n3�_G�<'����u���(u^(�@jIu�m���V�c@�|K�hŞWx�le��쫞�d7g��Gݯ�/�]֯t����~��`�{3�oů��:��1���񧩢��5�u�� �g�n�x�����(���b:Y��MqÒ̄56GS���J~nS(��.���4�;��G�.^����?��b�7f�S�ڻ$^�Wq��.��̌���8ƺ��=4j]�L��ϼ-�zg��m��뜑��S�4mV�p-ARY�]�KVRm�ᣆF:�������Z�n���Q��-��o��®=:D:m�v}�z�RLK��c��r"[4��Vm�k�4�����o��}1�]�y���᏶X9��1-���>쭤����Ѳ}�j��0���5�K�H��x�����4�]����v��e����։�����'�ggwV�:��v��=�b�%_�~gE�!�����s�>�rzOs��&*Z�(a\���I��Z!�Us%X�S6%�$K��B{g�LG:}�/ƛ�w��i�}�⮮�gm��`�/��{�R��%��6CWrڎ@���[2��b	���,�Ep3d�E�9��퉎ǧ]�U��k�p���k����hY%ն��� @
XCk<0�,��>5tDh�=qrǢ��ps1����k�_(�m���h�7a�|�]U����Z��ʄ_$Ei����+bF&~.���p��H�D�C-hJ��/����-����4��њf6Z��>f��6�OC�;Ƀ�S�}�~�g�q������gg]_�u$�/i!�����e4?s��/]���j���+�+,].l�I��@j�g�r��y����i:x���tK�?-���ک\m��iM�x̢3@��-�����ҠGH�x�m[#$#�5���6�<�Ni�=/R��g��Ԧe��)�;�s�qd)��|������H. �7�jZY�l���e(�R}x��n�C�5���΃U�>�7d��o���l��A"�����lf�[��)ûjj�l_��Q���3�ψ!��^+3yl"]5k]Ab��y]7�GT�w�$�5�y�3�m��.q��U������4(�>�ɐ�sY��غ�=���\?5~�O���Oe)�k�ߢ����rqx�͔�,zlDqN�t��e��Tþv���:��gpT���5Սl��e~'������vT���wT���|��b�!�EF�#�>r'�����_��\�e�ϕ�|�i��`�l�d�փ��乧x^t�<��ݜ�7	������>�6'Gܠ���s>|�u�c�4����N�u�l���l�\�������\ⷭ�$��|V�"4f��n��ʝ� ��_��Ao���^ ~�����D
ʺ�/�4WY�Ss3���i޶{�L�t,�}�mݒ^�9mI�.Pq��zzd�ܖ�DD��_f���9�2�}sM���N)=�8�������9�hWE�mC�j� "`""�J	�W\��W`���M]",�i�x`γ`駣��Ζ��S�y�+�趈�]"d6�Gd��'z2Ъ)�y8tF;��es���%fW��%]�یFpt0���-�1���F�\��Z�{���pB1�
,�H�w�sĳ�J�b
�jq�*/�igR!�Z{v]{3�9��T�Pc�nr�E��7����宦�L:�oP{��V�"}�n&��[��jv�q���{K���S����|T�9�ϛ������WP�1��G���6�\��@KG�4��+h���z��I���kgGp�Aa��y-���{E��j'gcK9lh��=���)UWV�-'�w�LC�C9�;�27�
�������ά�����R\����/���.��Svu4h���i�hQ!
b��þ�3�0S;%�tט�^Uu�o�����n�ʓ�� r����{�弫��~䗔K6���>�~[��Up���g�EYjm7�[��ʼ���]�%�[p�w}�Bq�uO8�3}0ǉ]Sݔ��/�a�o��e��<3#�lS��ǜ�\2E`X3z�Ff������P�|��"���P�1����_����f�I��.i�bߩ�z���y���p��+��D6.h�?6#������������<M���f=/���� hdZ��@��T`^�/Փ4���(�Qt�]so���W72=/���m_��餤��Uo�7�<]��7=���F8˜��g�1�.��#H�Gw��)��J�ql�OoE�~���8��yR�~�v�7X|0˻7��tG

]�̚������wz��=��o��K����Oe��; �z���>f>�?��4��n��Yk�t-�}]b�
N���'�l�MEn�b��&�κ.9���p=���yF�={V)�x�U�}��m����UA*�vO�U��5&��K���O�j��j�����=YX��Lõ�̽��-�i(���^�@ϳ���>��뽮�B�&F���O�ģ9����B��^��s���ڔ)mna�Z�`4t++�II\��`>[|x�yܷ�X�18j(���1o^v�)(���bL�:0.�`=M���m���6��qp�wkyu��hL
x�ߵ�:��ܙ�W%��s��y�J�3��Z`[W�V/B����y�P�����.��<&	87�[t�k��M��Z!�A�[l��'%c���+��]��Os����O3��o�a�˼�V���F�^a��}IT��+��h_eA����1�G��̼�	�t��ݫ�,7C����@"����h��v�3�gl��:��ԩlL�ۼGjM�~�d��'W68QVM��`��dۭ�&{*p�}��YB�ɶ\��ǁ��. ���W<yǺ��?��Y��~5�$*� �����|p�c�t�g��z�����a�Q[�o�kS��T;�����\��	Y;�]/
�#�T�hHV�p�Vn�Ϸ��֕{��7g�b#$��:N��q�ѱji�Ƞ:k�:/R��ԧm�^�O���0���M^�X`|9��;�s�ʹ��7=����yej)��`;;
&N�札����Za�6bb��|�����YSt������X!���5dng:|�/N �eg3��Pv��Y�%��l����9N鎬����:s`������iS��R�ٜ8sͧ�8"�*)�7�������CIҊ����Y�u��v+W��ü�t��fH�gEV�|m��;�h��Tɺ��u[Ju�&�Tx�����;Dջ��
�(4�E]���e'ڂms�K��
���\%t{^8��r٤�(����)�FI|��n��.��+�A� �SN�Tu��v��!��nvwu�G�GP�혯���� ^����si�]�ǀ��#/��9MHK9�f`����D��lO��]0^��z3z�ϩ�y��Fc{�:9Ւ�*"OwԈl���pS6�����(��dLo�m[q<s��y��K+�b��M-�F�N�9�+OoÑ�u�4VԮ�}Ň����g	]��.C��]w�Zm[�;:J�,f�sni'�j��;K��Jn��-W;��
�SYdu�%�� Rnm֓���କ� ,�ۛ2ȳz��'ُ�ZƄ��f���e�fm>��E7�\�3�ᙙ�v��2o,����ҏ�$�z�$fվ�P��k8Jd�;��d�٩��4΅|�=�̢n�����D�9_vT��7�	qàZ��S��̝ݛOEsvxb8,p9M�"���'�6�闫�F�:��@t��"��]�0��}����  @ 
 Q�N虮v`(0A1�1r���ܮ���s\��B�����7"���
]܈IH�Q��;��^w�љ.tc)p��6)u���<��݀�ή����wW+��w\f�κ������G�u�ۈ�h�9�ݹ�ۻ�x�:���'�Й�](�NQ.b�o眐���s�;�ƣ��e]�;]d4q���Ǘ8�9�u�^w�\J';&��\���ʞ5�c$�$�wc/.�뻱�nph��r��ا�q:K��nrE�w.���ƹau�\��.n��0�S�������FNF-�˒�㻕�gs�7NGNv�r;�4(|FjOC��Gin�C6ī�Yu�=����BR���5(�f������u��ɻOt��wq�L�� o%͵>��V8LIm��H��)eD?3��s9���ܕ�R�j��6�e�̕|�=��뢱�c����� {�	̳<F�@a�ҡʊ��q�3�Ut��tw�vh��
�ڰn���fi�0��m�,�lPtG���wg��L/M3T[R�uغ���U^��I�n�ɭ(B9=Fw�*n�`��7����ķ"1��Lǣ��\��[��F*Yh��Ž��pH�Ǘ��Տm��@�oK�4ݒ^0R��n�h�)�vr�6�ׂR��V(����v���Qb9��m�M5	/l����t��+��zfS�7t��ߔ/��:R�wFR5��O3
�;Q�yg��-�tʊ�H[tE��2-�wN;�7L�	4����tM����>����L��P^o�F>[8\k�-�F�EwG8_��3��Pm���ֈg|�8�<�����\��7�$G�������=�B�-����U��L��ǻ���O0�uTk>��	li����y=s���a�ЎV=ʎ�5��3M���
ۿg�Jβ�SEQ��j��[V���<�=�.��A�Ȧ�B��Wv�L2+C�3�������No1��#�ծ����(P��
M�$����]c�U�,����|M���{F�+ylvo)�|�
 =�����|he�c�6n��ÐZ�����.�����~�����ǭ�o6K>�H�q�m<fQі2���2ji!y�Z2�ٳQ%�xH��)O�,�ut^əDb�~��4�;�����˗�0 �qo�UMSA��Y<*:N^٣O�ͽ;8E4��0c�˭���,R�}��[;o��\䌈�a����e�{W�nv�w��ƅ�b|21�4���a3��-��bO{h]:���lبz���륦���
,��~�Rӱ,���m~gE�?!��� mԳ�z�q>��oF���+���w��؅�U�f�����ԑ~�`L!=ˈО�b8�iP�ȗ�]�7&��yj+;h�����w��#�<������	V�-�vLx�4LC{D�j��{�#<Z2��3�z_k�WR��k��N[��e��C�����+��h�S2 ��6��p�7���u䘒�W3H���b���Z%���ܠr���wZ;Cޮ������-h�/��Ⲇu
�w�wu0����Y��`�R ����e4�4%D�e|��,inΨ|��n�LkW�DMzH
��OkNuj�Q�ju=@���s'4���Uyc+��QV��67>���d���G�Y��J���W��:�sMyͤj滀��.��yϗb��ltD���o\�l��&���O�)�T�����tT�x$�V����Z�by)�SB�i�)g�q������vu���H7
�H)�x*��t=u�X��<�6r���UHK�B�Q��3þǜ1/o��X��u�5���V^<m
����<�1���1HAd�n�κ�ZqLOH�c�Ļj���ȘOtE4L¦QO�;��T�k�-���ǍT�2Jx������5�<�뮐\�hږ�{(TC��%7��h-�x:A#&��݂N��r�L
]�;��\�o'�yV���Oek����9������י��<dS�2.�dz���Ϯ�镓�D^.�~��1�9��R���&���ܻ�h�ť��#{�˸!�s��oکy�Y�u���o��s��i�����<"�����S��o�]�>��\�}V��评� ��>s���.F=4���d'xk��d�)����湫��Y��
��g��$!���n�μ��mތ�!�L^��������U����\R��%�w��i8px�g,�g��cuM��wd��Y2Aj4!�����Q�_�25���xׁPʅU��U������9��9��(<*t��@�;�}Iۨ�P�����gvoZI������Y���F 86o��Z4�ILLYi����Kˊ����<LH/��_��}��,��Zl����y�};���Ge*Ѻ%��ǽ4k$$��Z��6�>��K��R{�r�y�t�~}
�]7rڇ6� E��xhX�l�wb3)�_��e�3�9��Y\�`駣��Φ�1��B�.����[���yY���R� h�w�&[���5zc��l�%	�ī�q���������/�t�u�z�TN�q|����Dc�Ƀ�R#]��`�g䡱� ��J-�a*/�0�����gwX��^���GwC�4���ѝ3(2�p�)0w*XC�ǜ$��`�	�qT'�kj�*��\�
ޟ��W=�E�s�7t��:�4SuWSM4(��1Ό�þ��R]�l���PnX��i��c9�kn���T����@�f���w�t�[MyL�LQ"�i߷�Q3�)�Щ���;örEH�2i�%���[=#���\w<s��Bq�W]s�uj'#��ƻ�ݰ�:��n1��اcq�c�d�lo\�ҕT@�wK����uQ��g�w�{��Լ?��/��E:�#�[?)������O/�Vs��+{�b�&}�r�Ź�|#y����;+��Y���t/}�����l����ƀ7;�<Xm^	��9��-N�D���#λ/�>q���Zzf�o���.�GZG9��f�u��r����3�P�ćR逞U5��wF:Ҹx�r�uw|�R�J��m�e��o_7N"C��(ܣY�iuK�������n�{V�?(����+���~��j[t�3z���ʧ�;)�;��O޸^W��K,;�II~�Ӎ�L�T2���T�r1��ʨ�4Nu�I�SN3�[=t���U�-��ދm��/;fޙ�^T�_t���!����znh���$ň�DX����Iw{(�g��<��>#��%ͱ����lNF2�|O\�E�۹��G�8'�*:��C*��?h�	�g̀˼�='��(d��yWSf� ��ë1M����@/�~�ը�L�4<�O���ke��*#�KQ��6^�p�xgl��U�츰�βA�Ю�OK�
oEy(:!�����8��ƙ�*-�D��3P�/��R�%�*wvQ�5Q_\�P���B]ʛ��[�Ϭ�i:`���vh��z;��S^�WosF��N7^���}�s\�����uc�r�Co:]]�^0.����!�g�>��6���S�q���܉E�$��6!�X��*�i�#eШ�0�t���~Is���=<4��'�R�zeRz������ !������	�0q��v�o�+�uy�P�����)���#��ר6�(�f�:d]If'QdϳF��9j���{G�j��k�/��y������:��3�%'1�]��wci�U�A%��.�>���s1l�ɻaw}<�D|z�:g1���-�6YW�����tE��3�8㻥�#+e��.9�Y[[5�&��"�F��lO����c�Q�y�s�$漲�(�=wG8@�$CSq{���0�^����m�="��F��i�o	x}�pxf�C�S�����ʒu����̎��]ϽhKc.���M���Kh���1�j��]�']0GH�N+h��,v���}{n=UMk��"��9�OKE�l�yc�B�z�[O셪��c��㲯q5&}��pnsl��˚��n��غ_�W�&��b��_h�T=q�Vb�M�wfJ����z�9��T��Ϡ+�X<%�.����5(����x7��� �x)W�=�7#��l�]��Ҍ�jg����|\[��J���4��[ƙY�����N��Z:<�HexFm�qg�<U_
΋ɍ{b�cFߢ��q�i�:F< �c[w����,��SGW�J��3x��u��Ʃ$�l��vM^ە�4��k�|�F��G��e��z�1�P?�r�񰘚���n
*�>�WwV��P�Rگ�>��;�Ԅ�f̤b芻�=��u��Y}A�\��̭�%ckZD���W*N����tz��c���t���C�Jew#�9_^=.�[�]⏦!�� �Ne�0FҼ���ǣ���ӥ��,�\�m�=�_T���(���R4�!�������l�άzp�R��tX��C�F�[R���wU��v�w�v�-��O�\,��^�!������9]�eέ���Y���SH��LG9Bٕ�k&���(�o���Wa��]��ْ8�ŕܦlX��؛�4uק�	�(w|1-]��3�?A"�F����SM4%E钋�twcY=�ȉ�Ţ����ft=r����8B�0r�;�yҖyg�^)�{Ӯ��H6��L�JP���[�@�'Z2��.�h�n���D3�;�/��{b^�To�p�j�s�ɍ��ج�g�ܖ<�ʹ���hp�-�l�_SM)�� ��<x{V�Hz��m��9M�s�L�:Qcs"{�5�N��N�����|#����[��}ꞑ�D���ĩ(�sf��w�C�W73B3�H��\��-��I�5�G?E7z|���9�g�2z2�L�����š�`k<9��)�&sH���X�5,���Q��ߠWdsƔ�/����f�ӟ�fS�ۼ2�mu���iH�:�s��%oCk�3�_|�&�O�
JT���:��R�wqv��)I����f��2�[��%g���(t���X�0G��5�$��[�M����·T,� �i��ݼtWSy.��9�H��2>�oU��G��?����~`�ƒ_mr�ܲ���Z��6���v�2�z�BE�[e��'�|n�8��x6�}Mn�'���@�q�1��+Ꮛ�����ɺ�g���Aʖ�/�w`ų3����g���ub��<4緫p6u\��t`�!���4����W��<�~��P/7v��m)���̧]�t����[=��@�.�}��p\�rڒ%���E/-�6IUt;î�v���}�i��#�*��2s���*OtL�s�^����w-�s�XUXpjV�W��ɣ�h&�ق=�>�����k<�6�{�KwlGO�:嵱��^Sʫv��g�ܖw���1�q�}����,�� �����,�IXz������r빉��T����>
��e����a� w�PT9p,��iw�ϕ��DU�󬸖e1}*��H���N_��u"7����,.|��W�#�&�H��fp�w��x��e�Qw����,���%�9�{+]�4]
�����'@��h��V�:��L��C������Ϩ�MMcݱ5��n
J�^�e���(�DL�6�e�	�8�M)2k�w�Π�L����,5��=�-��Ҽ��&��$ou`<*>�ܬR��(�������]�5Ƌ�9��3�'����d��	�/o���c�a\��U� ��t��S���.��_�%Ý([-�;p��T����F:������TD@���*��TR�9�:���>��dT��a�mZ�ȣ= �t�|%���	�sX��'�)��� �<�8�J�Ch=�k�O�;ŢZα^y7Kn%�q��3¾��G���g��O<5�2�{,�M�I����l��w��'��+9�^���FW^�F�E�{T�����܏4���]�/������m��vKڷ��G���dW��_�\攟U���kDޭ�4��S�15V���V�^.��]�<'m���tR�ʛ�`>3�fx��źl�+��A�r�-ALZ[:�t�k��d�룵�~�*�ť=���/�_��m�̺��0̽���β�#kݗ�:؟�i��}���d�N�g��x����g��]�\��/�f��8>wW����:���^�!��Xj_�͇H�g�k������Zv2��:���R�ݸ�yh�\�w</}������9���'�*��<]C��yP�o���E���z!�0 To���/6[���4q'@f����B�:<����PpT7��S�8]W}0.΂�]��2�cGvT�7��$#r�(�7��Mv_W�Rw�cU٥���
��]Q������K�ٛM(��tL��3�2��f��7^pO$O\�l:0).������f�W�A�_��p\6�8��L/S1�D�������Y�UG;v�hx�z���緾��Ot��q��&���ݺZ�F�ͦ��w�q�09y)��Eb\	�5x�D�c�b �Y���_�.�{���t��ō���n�!˻>�;pa��޷"rh�5��s~a9.���R��6��i�H�{�#s�[�Θ}�����L#	��-�Ƭ�����;��� ��3��Ig�Z$��*b��h�8d[�~�v[�mX��x�l,~w��VDV���̀�����0�ѯ0ps峅�X漲�k�VwDD�>��u��-�@�#4��8�+��5(���g٧�Q�%呔B���K?C���[{=5���o	t9���Pr�Yts>��	li]/a�X��H��e�6�O�nV=�Z7�׍T]�`�n�r*��?e���͸��=��UMk��"�ts���i�M��,�D���Z�HB�%��f�Gk���#0v߶S��]]53n��͋��E3vM?NŷtH�߶й������^`ȼ��"�����R����A��;�Օ�� �]`�+��o=��T�%�f��w^0�=�={чV�X�؝]�IHV�F���o��H����q�:�����d��a��
p��9;{;9s���r��9�
��ӻ�ʑ�Y/ ���R�#�٬bC���CYCgv,�;M��2�����q���m:�;X������Jc�h�+;+vw��v�.���unue��3��jHAx�ed�=�yK��x7���� \�ǒ���()�xu�>���(3P̡j[�F%jEn7��1��߇7�������tK��u����,��lfLC�w08E�4�(M�K_5�a��3ui	�4Ӄ���x��&����^X�ch�A��C�M�7s�Y��l��74rd������o���=D���g#�F�JŪ�)�yp��9��4��jwMN���Tј<3��
Z�)�xM�m����'�{e�VڍV�ҦlJ������Z!�\�׉B��8�XtN��}��ʂ%���lp�=gq�V]'זK�"S=Dv]4r��� �˲�=��s<�I�S\��C��39�b���WF�T���yQ���彙/�t�WlJ�42T�!`��5��6^�l���V�9���*$kOsf�@Pџ!Lf��I`QEU:s�+=����a`]���8P)�".M���Ӎ�+�W�kj�W0��r��1�v0*��9m/�.�m�&��8ܳ�m?��w�
��D�{�����r�#3�Q^�aPړ���Nty4q����	
|G/;4v��؆G*��N#Ht�kY��V�����kS�"*�ʰ*,31����������0��0
Ԣl��ދ<�:U���<���d:ZkEu������{����\Y�-.�ت��t1j�ƗvV��0C)ؽ�q��Ir��j�+6�	傤��wc��W�8����y�I�:�7o�r�s�<�'��i�����߂����>uu��D�S.p�:���`v���R�9;L���5;	X;��|.S��Xu�=��̹
;�a*Zf��!���U�,W����I�Y�������=������f�u���RV���g����`	ҙ���G�;��&R�`�Yɝ:�����v�%A��n�P�R�j;�|'X]s���s��w�1]+�2c� s6�h�{�g;e|R����GwV�]��7�X�Ƿ�atw����8�'V)=0A�]�u��30�q}���ȣx���lX�`�em<���V��V@�=촣�,��(�T�(3�s���u��3JE�[�xaftݢ����`/��67,��z��=!M���ș�َ֚�Y��ѓ�PT��ќ�<g3H@Uk��"*�H�� �N��s����8�Mq��$47`z���5$��f���YW�]ws�$b�U7SqNWOGw8zp��6�O��C-���������Ͻw\��̦r���s����7u�7wu�戒#���˻� ]w[��ۥ��u������
#����8��u�;nW5˔��Q���	�w]s�u��.w\U�v;F����9�&�뮎�r���w\]�]�F�q�s��s��ň�h�u̻���cQb,H�5�t�t�.�������]۩;��nr��;�������X˻�4l������v�n%t�;�r3�Ww:���0�uv�wuN���u�K��n���"���L���2��s1G;�:R[���v��gwn[���r.\�\ԗ�wv�.�H�u�nG7	�nk�9st��k��bX��� 1�t4J�I�KO.� 'z3��^��Z�mH��#�Run�-�}�^K泗K�g���\z:�՛ځ�N���twtɜOK��?�U������,W�s�_}g�ZQϼ-��y��>��FcvYb�%����J�u�jg���>.-�U%�>�ڎg���e~�Pw��* iҚ���v�$��և{�6m6uZ�輘׿ٍqP�q�i�c�c��5�'rz���x�-�y[7xo���g9��3������tԵ缩�+�r��(3$�z_92f�G��5p/�O)�1�3K�~x�K�����O<�௪K�6Cw,�}i ���Z16�D�~:���{�כ<L�4�6:��b,�i�W�Ժum�����gl2��I��hY%ն������u�sϒ�sb���]��᭞<(��
i�Nx*3�Mw��m�K��^n�-��S��zD��ʨ�T&w��<�F���z%���9�v�H���7�M5	Qz�Q|��e�c\��e�R,�'��C�*��]ю8S&B��}�JY�ox�ppO�zu҇�d�Z��F��皊�べ����`owSFt���S!
���<;�9�{��
Cc��k��"���I����[��y�_L�|m}���=�CP��-�O�xL�6VGG���)Z�ƌ���})Z���P�^�h�T��=]��C��z��g����=C��/T,Z�]�
�;TW|��^�Z8���%�;6gR[kEN��-��ø�C�=�Ξۣ��5����ut����1ѯ<z�%��!6�#�{J^oz�w�^dM6G9������R�(�;�'|]�)��uK9ꞑ�ų�:�Eɗk����M���CqO惼R���b���<��ܦ	jQ΢����GZ/��`�W	e�Ov'���;Y;/3���~g�\S�Yy]����k`X0�K,��D^.�~�Qg��a��,ͼ���*S�'�hg��ƥw�� ��|�u���Xs�Z���4���}z-qO;�������h�9�:g��L>����<-�PFTG�e��1�4��5�F�}����U�<:n80�"����n{�+m��.��~��N3oVX����U��av�zX�9�ޤ�\����g���X��u�杍pk%;ŕE��=l��{eӎH��%���jH��a=�2o1�9��Y����V!���Rʧ&H���tr9�ζ.��T���t�����m�)9������c;�R�>y�0�+�#z���g�,<�[�yc�����T��^�R-�E�w�I��.ecV^������P�	W�6����/z�cf�珝Ņ�)�8'��}9��5�0^Jl�	l�|�,\����o��Q]V�s���T�&�a�\DunM/B�z�,V�%���tum�Q!����bJ��H�lN͝����ៗm�]o��eZ�I�I@P�νt��Ut���[2��&����Y��M(\��$B8hT9����eʛ�����!��p�F�ǜ�q,�9(h ���:wS�[yg�B�#��#)��������7a��]3���p^Lʖ����U.�9�w�Pz� gE�O8/�qV��BF�ߔ_Q}��:vu4h�uR��n�g�VsLR{���������_�NK����o�}gn9\�:���1�n�w���i(il)Um^F�f7�� �6�/I�c�j%���1���t��]"��K���8��!�S=y3��vn�2���w�f�s��0��5��<�,^u*=��l���-��0{3�k�C�b��qn�0�ȁ���}�x�}�z��;£���[�B���WN<�B��uF1�,�cZ�pD̦=˪�5z��T
]�^=R�[���� �[���z��0:�g�Yb�~�?;^�Cɜ��O��uV�Ʌ��غ_�+�+��u2�w�r��li��^�ՑO5;-T�iQ�X��~��\�<�3 v{*Mk�������p1Em�B��U�;��9��:���>|`��U���n�!��w�$��hb���NI�H�;��Q7�Iy�y�^�L�x;:���W6�4�:�<��I���ٝ���CoN�1��O?<�]m'��*��Q�Лz%�_��q�^T�I�m�D����\ߛ~<����7�{�n�T���9 k%;�z��S'�ڙ��auƾ�h<8�	�t:s�5
,�8�{M�H�=;>SDUd6�/%d�����������<���o.C9�e�X�i�Ю�WSfߗe��g)�� �B{���U1a�T:1^�<t��E�|�gb.6��KD�Ls?-5�øj�Q��aM�^8I���|�O^�2]�_w����Rw3(�}�ډ"6��{{n��O��!�R݄)�k�5 R�5�U`秃�(.��Q��l�Jh�R)���T�=j��˄�m�ܞ9��t7�ōf]]Mף$!')�z!4���(�xNΧ��5���w�`�S�mwSM4$l����#{�=�>������m7jߵ�Z`���L@��ܨ��<�vи�<2�'7i���Hp������Xlח�n�Wc���{\��z�h��|����s�^i�ah��~#X漲�f^~������ ���ʚ�J���`��Ɔ)��`�]HJS&����o?vi����mx�_��&S�r��%����y�h�ʽ�ż��1���Mղ���N�q�9�T��X�Ғ[r�7���˜]y��@I��# �c�6��.�Ka����b7����
��yW��F���ϊ]}�W�KǘK#c�
��c���8������>�7#U�]#� ��s!-�,�^ü���b�3<m�v�E0j�~�kT�]m����,~���c�����*�z����e����̅4ح��g�=t ��+���TԬ��ص�_6�y�l7SN�`��m��|yl��NOD���G{�i�v/���ou�L�E�9���)�]���۩�W�S�I.�zYR�����l��[I���	t;�Q{x���鬩�|��!��s.��]Qr/9Hq�(q�#SM�覐x�붙mڞ���3��o���i��zp�n�ͼU�)��~��a�'��g��i����q}%.��Τro�֦���؊�����m��,�l���9mI�,\'�g�:���ɹ@U�ut9�}�B0>�ti�*gy8�_<�Gp+�K񰦴io{�cD���n�9�j<��%�x�h��8A�x ����r��j]:��s���2۶y��OR~"�d�QM��Q;m�s�WI4P]��Ix.\N���U�5"��r���"������;��"GW6B��ı�7��9�un�Xd\�r�ʽ�Պ�=s�C�̴6�RsWn��{�h(j�u�<��eq�2�;�W"y�KMn��;�՘�M�����b�vj��#�X�lg�7e��"��P�W2�6Mw��m�:]֊�i�C���˸Ӊ���+\�h���ܨ���&X7�H�J�Y�*8;�(��Ux"�s���t���]�vuC�uM ��F8�I�����t��|�OAy�p�i������Ӻ4��*q���ʻ�[t^�ы���Φ���UW	z�2����L��ĺݨ�ӬN�A$�u��z�g	�}kj�����q��3tF +��������k�bzA ::327�+��x�VJ��wn��9"�rȚ��R�MOL�ꗯwt�:ٸG;�_���ye���hi��fC*�6ߘ<uH�" DS�i���?#�-KZn��Թ�L�ڼ�O���G܏L�ۺսy����ˢ�ڛ)��R�L����l[����X	l5t��OUZ��*ˋ�x�Vc��h�z�~�����=�Oy�z�W�N戸Ni�#SON>SL,`<m�h��Λ�ٸ;I�913<��db{C[gsN��x?}0���W	�m�22�#�2��ҹ�:5����k��������Uҫ��˰u�#���GJ(�{��n=Έ��������>��x�q�6Y�s�##=�K��&�Q�H�[���/���aԛ A�+w���٦Q�z���Ÿ�u�p���j_]�������NGچᩜ_ugn<y�̾'� �7F;�-�/�V�o%ռ8��[z�Vu�N�th���t���>=�;ftňpK�ND覞���Jw�*���<z���g�A]��z�]{9mIt
��<b�����d�h�5�Ua,��L�^��i�y��:�{bT��j���}w�DU�B���H�^�D�۝��� �1��ɇ�i�E�Dbn�=��9�x���5�K���Gt�����w��za�j��=�_m�e�Fv���1��e� L6y�zJ��P�����"oK�=d��e�/3u2��d�p����r��uÎ��R0)��Aq^q�C�$�s`���L��:�}�5ogjW>=�,�DcoC�5�i�)uW�ђ8S&�K�|��.�q��z��E0����B�n9�N*ח����Q}E�=�'@�vu4h�-8��#�g\QVU@k�[���K �v|<������0e���ç+��];ñ�F�]�:�2_�nݜ��t�糚g�z1"��c��dT��1�.s^Yg������.�njm��f��2R�ͼ��|�[�ô�A���2���o�n{�m?s(��?�W6�Q�|�E�+s��:�W�2��:&�H�ʝ����OtW� ��==��t�$��bP(QU�(5w��w�F���Z��|^�밺�_�����"�hHIӛ.Z!��\�N;�.�N)����1�b�al��zc���	��,�,�Х�3�;Y�Bl:�1�y�.�w���?��0���~|���uЋ���td��y\��0]�� ��U���e���ֹ�@\<f���m�|�� Y�m>N:���'��Q�J�*�z�Y����F߶�e�[��<m��t�DWdW	��h���*l_ a��|�Uk�ƴb��D�z�����s�T��^l����u������OoF����9�8�}+���QQ���~�i~W?}�� �l!��̆QQ1�A�d�w��y�ЦO�S<��.��)��~���<�S���4�����e|��s�6�)��qbDl���0c4���V�g�r���G��<m��`�ć�A�$��ٷ�����d��ռF��i��R�ь�����f���[`u�]���ΨC�_twm�i��0Sdw�8���a�Y��d5�
vQO�n'1f�eNS7��-�jQ/��GW=�k�'��!��M�l���� 'k�ؔ=u_��Nkg��T��{G��A�29^��~��4&-����D �z�C'�\d�cf�t�<�W[��.ᦐ$�f��'���Q=�hq3�o�Q%��&��C�fku ��a�]ݣ��5����5�O�rRK���r`R��r�:bA�~.��ǩ�HT�s��U���%Տm���ΗCi��K�
]]M�[������@m�5wʩ6�H�#��g�ᵞ�R��1�V�u4�$l����#{�=�zn��؊��z,s�x���ff�y��
)w*%�>��JY�B�g^h�9�L��HeY���m6�j���^KD:��cgR�}���@	��F)�w���M0�s峎#:�z�RZ�?7�s��SLC�M�)��n�����w�xO<��%�bퟟ��xN���3��[yo��:�ge�K�̈́�:��T�$���g޴%���K�w��= ��^7�]M�F�v��ف�ܛ~i�8&��	��M�9FfZ�~�����օ4ئm��gf��@�x���\��1�WR��?^��/EL�ɱL�;n�{}˫��OM~�b�~^�~���K66�&#�PGcO)��=�g5�<�w 59O�Ki�U/Y(�'�9u���g�m�<����9�}�g�����/���\䌾R`���-�~8L��W*�h��\�r���{+�b_w����q��MdޒS�aZ%4r���Δ�D+���9>��3������Қ79rC&%N��-�:��5H`�����M�*�:�*�v�o&��������c=� �����E��Ï����Z�s� �F�f��3"I����/��Q��b��}���p���]�1z#��u������}�[�V��옔�c��xf���TG�=���=�tٽ�d1�[RL������]*�/�_��1�\���f�$Kň#�C�5�.�`T�����Hn�/��)����L���s`yS��w1�p�LZx�y�5`p�<�l�w*�&���ʭ��^����~���F墩3�����;wC�w���ђ8S@D6���,��By��Q�d�p���i60�HHn��=Y�cw��5�W?^��2�w*%�k��CZD�_����>��!��:L�H���F3�#��׻:��%��1�
�`� ��)gg��^B�0\��~;zf��a�	~��'][B�H5�E�-̺�]�M]U\%�ЦBX;�-�}m:(�>��~ֿGjr���U�Z\~��3gjQ]I�ߺ8���Z{��Y���i���ϼ������ic2��V�P��	�� (���1=�U�6Y;���)��N�FZ�����o7�����7��o7���kkZ��kkZ�v�ֵ���������ֶ����ֶ���ֵ�����km�ͭ�km�{[Z���mmk[o{[Z�۪֭[��V�Z�+[Z���-mk[o�kkZ�z���m���ֵ�������Z�ֶߖ������PVI��YP�&A�}�` �������e�y)"y�II(�R�R��UT�
���R���T�A*	k*HCf�U%UI$RJT
QJ��mm"���L�F��hm03ۮ�k+j�+dk;��V�V��5�#`�em���lҵ��6j��V���j��
���eݴ�mm�M�USikfC��f�kI��R�J�Y��R�h��l�6���eJ�M��U#V͛-m5��@�ʭ���T�m��kf�V�f�ͥbE�aEd��К��
��Ƀ�   ��V��cy+֡�Z�5֦V��)u]�\Z�l�݇F�:7kP`F�c����U����8����wm��f��Q٩6�5lk5��i�d�   v�Ъm��M�^u��k[C�Ύ:(��(�(�����EQE �;�
 Qb��(��(��z:(���=\QE(�F�tw  Q��s�M��������UZ���|   �ޣlk���iQ�M�Ԋn�����Y wf7Whvgwk��\4t�u�V��V단�WAZ�ú7`u�v��΍UV�V���6m�UClSMx   c�)�Tk.�uݵ4.ն�]���X�Ruww
:.�����ӮnN� ks�����ۥ�n� ���8�S�M���օ5M�S�ma�Z�Ujm�(�K^   w�`W@��� we�]\�����h�nWj��7r�P�3�ն�A�ѹ�ܷM��Ӛ�ҝ;`�8�[e��������G!�gs���v��-E��)ٯ}QI	)ާ�ݫj�ݷ1�� )SGn�+��;���42�vƹGD��9m�nX��nwv.n�iԬ�t4˧V�]��hk���M���wj�클��C%S6�#FU[| �*��>��ۭ���CP
�V떶]����M�fw\���wv�iݰ �S���r�*j��r-N�mm�4�\�]c�l��Vt��v���kiZ����lkmJ���
�|(��}ڸl��n5��-n�m�����::i��e+��1ݢ�-�5Ӯpʮ���gg��T��nK��ۭݹ��6��]ҵ��5����e�3EZ����@��k6�&�ܮ[;��ӵ��M:wv�tvt]��A]�S���ұ@:4U�����覣qƗ]ƴѹڻv�]7Y���)T룛�U)65Yf�6[m�C[f�:�   ���i��˜U:i��lB�i�ғ�XN�wv��v��t�ݳ5������'sb��j91V`j��9UKf��N蕡��O 2�%  !���$�E  T�J�@  O��P   ���Q��P 2 1THA���?���g����?��������K��N�#{�Ͻ:�~ק��PTA]���TA\��
)� ����D�DTAX@QO��Տ�������~:�^�y�W���%��Sk,QZ�j��E�n�����ê��r��a�̖�d�u30C�����d#n�<�,4���k:���*5R�'^���dF��NU�F0ۚ�Hޒ] �=���ikK�νJ�!1+X����K�2��sT��fa��kY[[x�����F�a�G��Fʦ`�����F�3@hR�n
,��-٩v��LQ(=٥�T�\iT���Gy@|1cX]5��Q�ỗj�c��Heڛ&�Vt��
SV��ԏ%�U[FKcC?Z \?Dw7��٘��!cԫv jMP���Ɍ��T��O]dɁ��*;�� zᖆ�aV�� �\w��!H�El����ػ��Ƒ(��ɴ�s�z	ug�2�m���XJ�����Uշ����i$m��n�4�0�e�EB��:����y�EJ�"	s6�7&���%�6�M�fm�l�T�9��)J;ܑ�YwMnC7�[B00i�5�4F��ɩ�x� ��u�����!yv5�8$��q�V'�f��l�A7�}�KT�#[tnlD@���AM�&�b����M�Yw��*dG�����#�xM=#7�i��Y��Bƙ���T�x��MJ�"���Yn�����2�I��-4D��E����W{�뿠YMǲe+ڛLb����Տ2�	41�u;P�%+�KP��˥O��K����HV:�l_ȶ��p��+��)<�D6UҤt�̖t�Wbk�sn�9���R*`Ѣju*��+M��4 �4K�T��0�7�I��J˧J�ԁ[�YQ6��OaK��Dd���J��[,�q<Sa��BXmnEN;F��p䱕cT!P�ǈ�H�5x�C8����՛�ܔ�M�����j��P`Xʛ �ʸ�˺�(���)nDi+Z��[-l��"��L�W��yh�����ajGJ��;u6m�MdS��Mݺ�U��)jVS�3)C[A��$q�	3fh �6��`-(R,,-�P�D�@��Jn�e�P��t5IB�kQm��ʷ��P-Q�tr�bё�[Lٵ�LKEd��9��6�!�#�WE� �͒�XsD)�*�������H�#�5�Q/([ �Wyq���2��,���X��V	q4fP�� �U�ë3h0�4[Id"��鰯��V�l
���ı�
�DÂy��BV��HM�X��*��0�CS!�*�1J��1S$�I3t���V���e��,����7Ԝ�v�LSϤ��lv�F1[H�[B�$�ѽu��dc�0r���N�@, 4�c7@�������' �� "ՙkCz�7hf^� �oh+������P�6�� BʙI�t��ʗmCIeH5��Z���.􄮧�ȅ����L�*�!�#��7�xέ;wn�k]��x�����H"��=:�Ԩi<q�ُn�d�@�9a�Q��1'��YDң��l���D��v�9(�L��A����fm��n�nG���1ikd��v�$��D��ni�v��h-U�D[aV`d���Hj6�`̙�����0$i+m���l�Y������#ي�^�L�
�R��a�%���~����pb��p˰��]Q�a��t륬��K]�VtXu�a�$���e�7)+����f�:�Ay
5p�Eеm��j�z�	�AS��V���ݜZ��2L��nf��kiM8�����4���i?-4���"��ĞS�Ɠ�G@u1m�^	x�&�b�h�b��r�t��B��HUn�k�-`i�(Ƙ����J���>��k$��:22�"�(ۭ ���Hd8/UJbi�:B:&� �DӒ�:��b�E��7��(,�]*�X����Vުt�j���ᬚF�JVUf�D�Ֆ�n7�+vv�<v1Y4q�2��$�"T*c)�kc]{NԎ��);�P���i&^��jy�v���4��0�Jޭ���ՠ�ٽP��KJ�n�n��ٲ�Ǖ�Udȩ&>M��.Z�
�²8��a�N��,^�t��k4�!���f�sh�p����eJGlV��	JX)�I��u�5�k�4���Qy� �w$rF,bɢ�߬�`��2�7b�*@�%-��w���t�h5m*�^Xr9b�����z����n�(OsC8EN�l;'i���٭O*���6%8r"�e[�Gp��m�F*��E�V�����!��UĪ5�I�)⭸`ig�#R�3!��Q�-�4`��ip	WB�%I�fjN���)1�iKwohJ�օ�i�!�I�V��i�Sun��T+ ���L<BZ����aIim'y���J�U?��f�[�-#1�9SE�N���2� 7,I��Pu�ݸ�`U���Mڗ�4�]LX���5ܵ� �JV�ɘ�2J��Y֙���>wP�f��k!��ӧVt �-����B͵���.�Z��ݍJ���Z��4r�%V��x�p�Oh�[�4R���\®J��L��.�\2��Z*�*ה�W�nm����̛���E��I�x�^<�=jb���~�Ef�hR`]@��*]��ͬT#���cˏ1�z�m=�Ջ������Ym�F�䧆T��,�(+�����H�k	������\ �7Ye�,e��e��7O�[zD��^m���(ؼQ�C7")Re*��<�� ���Y�=9yl�ˤ�[�q���F�h��2���-�1���*Jw)��١��`���j�ر�d�TX��dE��&S�Wn}6\��ٻ֩�*]iN]1����z���k�e[ض��v�`���Y-�n��+g�Sv��2-٭��Y$��ڵ��Հ��,=#v�E��J�r1�^�X&��GtV�cQ�j�[���n�Ϋl�{{��N��M�����%�xX��4���5cTc�S�.���0�
af��\���6$U�*y(�r�M�j�ɯ��1e܈o/q8�
HkKۺ׌��5���]6�:v�i6�n
$:
�wHh�w��r��=�n[@:*�ŵ�A֙��"ݔ�VACo+FI��@��ŊWcJ�uN-.d4�)8���u��h˭$�r��ñ�f�;�]��U�tn�F�1�y:��t��C~#$2m�U�Q*I@2h�-��}���e�6f��p�nm=י�3jB6���% ^j04%��f�4�N�x������0�FnH�$2�f�f��6 t��GU�Ԃ��A�,�6�f�Im�!SXM�d�m�!ʺ֬�2��]QXoqb�V�Zv��C��Q��IJY���~���SS ���{�o ��^��@CB���W����ګ�j�kwa	�VQ��xY�\�Ɂ=�3"�u�i-F�m�S��8�6!�nn�U+(^��ċ���v���R!<�j݄�"�M��owo/n�Z*mŴ��[�Jw$$,��2}�]����/%�I^լ� �N��ܘr�,P.��Y���Q��k%e:/	h�l�mA'Mu�v`16[t]�u&H���wi[O� l�c��婨�P mV�fV�ȥ)0�6�keH��Pҵ�[Y�����y=6;Q�=���=����
O�H��t+J�-f*n�sE>@�
nU�(#j&gԷ+Z��o,P�V�x�%��[0������9N��i^}�@Hh��A	��-��·��}w������a���3mU��`�l͍��R�k�z�fd��"cFSjh.�z�˦n�&m1���4�5P{����uZ]d Y.z`�pF5ܬ�u�N}�*J��H�X�b�1Ǒ�uѤ
�]Lyql�6�(-uV�uwM��ܰ��%`}�䨩J���c������y�xf��@�$�X�D:�y��2]�0m#��/K��;��dl8sh*!�V��7Xn�RlSI���̧�੻)�U�R�[t4����Z�F��d�9�S �w7A@�#X��&�i��n��ͼ)U�p�Nӂ�k4V�:�X0�j��L�L�Ρn� �%�k��7�OtV�U2�@�B�%�:8�Y,��<Y�Bܢ�N�����k3�>�n�5}�64	�@�"5{ݰ�x�K1&�2�.;�����
e�����T��m�f�&"�7riՑ���J�t]�%�$���'-"]5���
��X�6I�&'B�V�n�"����6���n���1Z�������Oq|q+�A�Eإ�( .�W�٬!�.�����$�	6F���h�����V�병k�4m��CB�<P�s-��8裗O)K�~dݪr[��Zh4�k�OD�i��7M��n+M*�� �=�V����RS#�[dmԴ�Z��E�l
�F��X.�-�)yhM�*?��k2�1�H�MQ������x�x预��S٩	��<i+�1�ka����jH�e�WJ��𽔛��S[o2,�ɡ)L#���4�[���ɔ(��;���)I
�l�����q蕐aL�pE����7b� �ۺ2��z�[�d���e$@u+̺T��1W������1�9g6�`Cb�m�:Ν��M�3e���X13�
t�l��fM�iH��ee�Q��Qbd�w
�Zj��z����e	b^�ʄ��Ae��&dg��1T�����QS�1	��/J�5�Kj&���A$Khh32I_d� �|��,�G氣M^Q�,+�Z��N�M�`�1�v�&�J���jח6T�ۡք���l憶��#m���� )喫^�Ѵj�&��i�庻+;�Sw+V��8Ժ�/FY���������u�p�QJO+S���cw�Jj��>b�w
���tU��f�\,S&���H��W��`Ctn�,3TH�yn�5�Ś��m��X�� 6��6&������v#�m^P�r� I���Hq<���q�F�"�dbٵĚ @��P�@�c�J�%7��c2˒�qh+r����a�ZZ� Q X�@W�A@7VJ�*ļ�Jɸ��s\�*QU��D���q�a�,'abۺ��`�H_G-�w��+]���f��6�JN��.���Ê��[K�e!�y1��f+U�#�!�Z�l�� XN�:l��0�5�r�7#&�<�
��N ȭ����J��Di��B�t]��AKC2j��0��0T%P�F0��)��p��z6�b�,j�xN}�-P�B�f�b�ma6��-���Ь6ֻՙS��&\:�Uo	�1�*Vʆ$CW��m1V$j���X��ӊ�T�KI��.��w.��E|4Y9-TXV�T��
�lV�;g�&,�_"j<Ӗ�^�ql�n�5�
�vE"�Z�,��$�ߠs��ԌTX�:�0�)�ݒ��[����	i*V��""�3��YN�۠�����{����&�V��y|�-b6O!=B�(��֗���i�����c���m��jh(���7;�셓t�X!W7�V�ҕ+��N�ǚ��+!�>v&�qT�:��[y�ƫ�p���yg09�f
����	��ȵ��%)6�{m��岤v
kQtf�����6�4NM@�e$f��h��� :�Xڻ�516���h��,Z�j������w�tP#a�s[P<F�:�#��	����������M'#�Iմ(3f��ި V�i�8�VؙZCϠ+qHLe�u��i�����(�����]�5�V8�HQ��R�[q��$�S��A�u�d�h�V���B� Vm�%�)�9���Z�L�VC���0�,ӛb��pᘨ�R,U ���V�Xe�N�P�F��*F�����A�U�p��$56]a��d�=;�l��3����z7S(ѣ31����B�z)��W��y�o5X�"]��.�э�kN�y,fR͚̉��0�o�t�W�V�Ì�[���0�� ܻ���(*ܫuw�l�n��ؔ����2��
���򅥡8T��x�J9m07Z�R����e�](&$��=Eυ�r?�/l�X54�֡�D]rɈժъ�kR������W��S�X5,�ڡ[��`n�l���a'�,��6 2:�>2(f�i�R�څ�l�T�i���l�6��q�ꭐӺw+2�"�kBY�kP�����2Vjvʍ��h&_�6�m#a�'�`���@F�]��"���r�M�F�ee�)]�P_�.�Z�V6ִjkͽ�F�Zp5�_�bmP!>]�oǇP�M���l���-,n�(��aǐl�ze�Ԕe��O(U�X�ּ���7J]�.�V:ʔ3#�zPّ'��\X��j��RR�m�c:�o,�Y�b��)%,Ի�QԻ���&Z���M�f�lTT[kV�Y5�
�v*k]�]�ٳm!�wj;�a��n����ƹK�<�7��J��	E����u�w͢4jN�̍Ln��i#7L
��W��w@�cj* 5�U��c^U�ZՊ�ő��{R�G-�����u]�]���`kY�a֍�%��%M
�u�	C��孵S!gc�p�r��ȃU��gy�^��/�JA(�n��y8��)�;W�Z�a��f���PQ�{���n²ȝ�Y�d'j�ب��:����^�T���/j� [�mn�K�n�ߜZ��pS5y�%�V.�JѼ(�����
�m�+mM�7�ߡpP�P�u�֙���"�:D�F�7�<�d[�a�9GJ{n��.<t�Y�6����Xs,Z�� �"y�rfؖރ!B�d���kOfd���T�yr����?n�j�c.�Z��l�zݘ&q	D�]�oثe�0!�W`��{`�)RA�N:�Fp���a4n���e���;r�K]�V��ڬ�2��[�ѯTA@�p�t��w�]�#ưH8��_]�M���C���Vh�n
v�E9�ЅS�,� �u�Mr��xeq8�!�Ce��AC�ՑM��]����S�^�Ү5ʞ��U�n�ʈ�дG]!-�-�U�����_[�	�`Pg����)fzUWW
s�)�R�Ε5E�VE������SywdYVGzR����ѱ�l�8"�H[7S-eVf��s0�)�+{x(�WVdI����TTN���f3�(�SD�0ޓ��7"x�8Qk����@Mz��u��)P�ܺ�J�[��vBäs�z�Kc4q�vUoE�u��F�dlɥ��-���r�!�l�)n^G*f%����^����q���EU��^�C$�K'<#6Ұr֫���Ͷ\�nLǛV���e�"��a��*U�H%���dK2�	g#�r�oy����g*�{��P�@Iq��|�^���oL��U��9[�2�M�z�O�����zݷ�,��!WUrI#�9ö0������Lq���
��� ��U�U��]4d�nkvJ�l��e�}�v�S��XGq��-,wuu�˻e�N�Ŕ�;�ΎS[�{�+��s��X�n0�-Bm�2�1jӬq��.��	}8d�Ѱ�9,���2�w"��U�7@�y4`��.�Ӯ�c�2b����/�H��U��ʽs���+sO���y�����6�����U7A������ԑ��vI؏�2������U.��;�
�Ѭ����φ�m��zAdF�m[�D)�h]K����l����@��v��:V�.I�qF�fiox#�btH��RS=Zz�!��r��U&˴a��v�4�PT輰:H��6V�ng(^��C��t�r���l��8,G�Ȇ�F��A�3��@�ܖ��ާ���9r�5�W�x���O�K��u���8���+�1�4�[وu����ѳ���yԚs��ͼQk�q���`re)�Zφ��m��B��HWn��wuXn���4����A�J��V�ԜG)�a��U���'*_c �����Q�6CW�z��sxh�h�F���*�åS���X<�������K����!ӝ��yٗ��Z�����!z���m
QD��fvo6�����$��[�m�:�Z<V�ϕ`��f�ĥDA#����x�Ν*u�9"�����Ы�Wju2�<�˝QX�s�� ��
�+�ϴ��/�ݵ��4[r���O:�2�	��h�:pɚn�1(��BWl�Vp%��YL��δޠ�+��k_η�NK�i�묜�)����j�G1����Cq����N������\u��Y�vdl�
Į�s�����'�u����;Q���*5ϰ��.�,VFq�B���g=u�OI�z�#y��Ӄ��&����	�1x��#<���qջR%{�#�*$���c,���n������avyU��@%vVmb�7�zb�i
�6����1B�i��>�rB���,%9-ク6�z����u�Ę�9k����I�1u�ոó��'i�9Mޑp�j�?*�;��X]��-w��5�@ ;�Xګ�Y���)>�9n*�Ɯ�EA�*ݡ��'^�q�:�@���L�U!�jt���4��e؜�9]r�s71Sׇt�3��s���gfۭM�{��U�@�á��M'r��tn�{ft�(�Ò�ql��+~Gh�	&ʙ}v��:}3k�]������5l�P�;nK�wl_nݪ�Ũ���@Ym=ͬ��0�h���GS����"���+�m��vN3c�0	��wSn�2�/�*�6�m)0�늡�K3O�5ʽ��'r-P��Y�v��s���3���iN��ky�Z8�F*�����b��A��j�q V#���C��čc�U^́L�D�Pf�$�V����3��q�X�Q���+��A�w�|e=�X���)oNtߊ�uեX�̒��k8�Ļ�
	*Z�H�����>7GR:p�/G�>����]���u��-n<�4Q�e[�50�S�oSgY�]�f1��.��,[���[�+�<���ؾ�r5m�1 �>�}Rk<��w�q��mkR�+�B��5y�-\�x-�մfu����+O*��j�m�˭�+X3�Z1�����C2���V���g�������K�	����O���z0�twc��v��������Ν��V3���T��빮�r�'ǘ���*Gy�!s�v˳ ���]��2�t8��5G9W3ofuy8˚MI|s�J��U��K�5-�˛&s�J��x,q��vww%��2SA��ڠ��:L��V���^��up��{��
���iH)���U��0��d�d�n�VU����U����E�n�U��w8X��.�T&#S�@!�Ҭw�)�9��PK�-Lap�ř�6��6�R=�v(�� Wv��-���ڦ��a[ ���g|)�{�� "�U��v�f^Y�zj){г�e��B���P���,��H�ji��C�*���Wƺ��ս[�3y�.G�l#��ybe�y�3���]_a�*t�3t�n�7��nL �}b���σ��%pB��v%v.E���)�.��k>5*$�؞ٝ[�%W'c8��D�W��L�8��Ii��Zj��r}vHS�x"���^����\��쌬��)�㮝�f������#q%��e���>�[�7q<=�먲���gLT�;������˧	<��6��E��͹��;t�Ϸ�G��V�k���U+%��F�-�;ya�5c/7Y�"����z��1��D�R��~��e'�<۲k7�V��u]�$p��i���L| ��v�8a�΍7}.ٸ�c�7s-7Jԛ�uӗ��8:����c+L4�w)�$vJ�8u/��WK�n$mF��N�>����u�i�ˁ�~�8�8�)���[���kK���e�q��B��(�
mgw]���q��ր��K;�K���h�Y&��N���n�k�(��+��V��A�Kt�Y����Fkc5�"�K�)y.�ucE'!��j��	n�n�o��}mt K�C�\�[K��ȥop��L1
�ʛ.dU;��f&�� Ʒm��7xvX{&G�s��mr쉬�Q�J�]ݮn��qOGGvlԳ�*�vY�ج.�
}�;��U/8k0<�ۻ�<W��,^��CZ�ٲ���S:)+5d�#sE�9��C��t
�Q���^#�n]5�0iW�u�����с�}�$�c�)|0�X΄^%���7P�郜�(�b��7VX�����[�J�FItOWS�v223c�
���ۮ����y�>��X��ؼR�@9����لE����7~e��
�-m747g�	� m�k�8��7�% ��r�&B�u�b�e%W����QPY⚒�g;�T�ۚ�t�ﭱ�p0��&d@��ڲ#6��\��d�7S�C�y�P�\���s�pu�x�\]w�d$bt��$��q�m���3|'r8��qMР?��-++> �Տn����pp'o)[P���#�hjx�����rʛ�q��Μ���f�E��H�+sX$9k���cM۴꫇gT�L9H_J��Wd&�y9VVj,�z�,� �N��x)Ww���م )�z^��A�0*�����4��R=f��"�4.J���K�2qA�X0J+rcM��>X��z��\$�D��ufG�Ĳ�d7�j
���Z�]��Oe,�/�P̀�x�Zr�2z��!e	����gP��@�h|RpR��e��`[�N��7��$�\�AA��]�j�w9}��^�bn�vKZ�,*���r����~��'�b�ut�(�:�����y�͹�fu?�w��AnX��6%^TW۠Z�1�Gk�'h)�7�7sY�Y+��L68��-��X����h��Kp#�l�͔��u9�ʖ��K���Ml�A�kv<�����v�V�{XDوʶ�al�]��kOP��vJ���e\���"�W�3ݷ�ߤ?�=3�NI�6�N��F��:Zܬgi�\W�&�,J����m�L+0#�q,U�۠�����z�0_3=��bz��8{�	�'�n�\�Kr�GI��3`=�B,�{�+6���[�V�"�h$�F�Ӡ�l��q|�)�@+ӖG����5{������.�wz_dz$��
�`����.�ƴ��/��X�W2�u�N._	Wt����(���H��v�1��.���\�,�A3b���.��\�Э����g��h��͂��lc˴���u��m���_<ASH�\'�����ZVᔌ	ᘀ��S]�,�����y��k!���)]Xrƕ��s�:�KN�L�O�}\�p�B�NtN��m乵l�6{��� kok7�d�2�;��;�*<O���ih,[�R}��=ovho+(/�t�70a! �d�q�ڔ��]�8]�m��28���2�R�n�n�;F��sJQɗŔ�
2i�`C���x{�.v�Y�³yP���#��2�ڪ��� C_j�}ڌ��n�V�h������T��y� �ōܪE�͢�*��;�ěznPsJ��\�;9��R��ʵ��sqkc�F3��ɏj��갠�#u.@ֵ�S5j��4Sd�\��>�cX{[F.!�������3�oL��G^��a�θ[��ä
S�u����q+�uL�1p�ek`�Lw��{{\��[P��"�m�A�ݺ��_�I�!i��J����y�Eu:�p���i���"��V0}ʛ�x��kbp�6챏x��P�:O�Ym�+E�+�Z-wD�U���u�Y�,3�}�n����4��9���d郺��G�uL�7�Ӫ�FotK.m�J�)tϫ b@��7��w�Ӌ��׃��b�zo�o'.Z�pX;V�{�D�u�3���v�,�Kcf��6�kqn����nm��+�Q��B'c�TJŬ�K�H��M�e�.��
q�ޢ����<��R��:����y,ԫ���������0��ɐԵ�_f�*����#�����n�)bw0 Eqw�C[9��nV�2���ͽ�ެa��n���n�p��-E-�ӝ�q`4�@o:���
�v��KlSܺ�Ƭ_d�oU#AvPX�ܫ@�Y��^�_A+!�"�8�+WK��U��Be�Ԫ����QV[��W��JFI�e�Jp��u������j�rg��];��D�;Vp�Mp��X7}H��x��\�WՀ����^�6�����e8�����vڇ��}�œ�����f�.Xo)_,�2�QO��ٸ��|ZYՓ��R)n�A���t:hn��������%R4�ͯdhZ��l��c6��u�'��������<��MGs��܆+��v�-�fl��j]H��h�3���0ä�˜�*K���f�9a9��os�%7�#\�en>xH��̕=`�w�K���}��e'w<p�!{~�#ˍ�-5..�FU�:�MR�5)���s��7X:�|�j��x����f�� ޲���{/�nK���pʖ'+/O��ܢ1���b�h��0m�pnls��"�d]�R�]�].VFƾ�u�XpgbYX��%1��m�[�'��y	��+si��e�w����Q��d����Zo�<wx�)�ѣw���PJ�nC},i��n�p�[�y۬@��fq2�t	��kηD������vcu}��v���W�ր���w�rH'i��%eM#l���TͬLnӑY���Fm\d�&�/a��|���8�W|
��M�Z0��,�72�J�v��a�	S���{�ktpl͛��^�Y�	BY�nÝ������u2��z8D�@�c��6��(��y����s�o�o*#� ��+iXݠ��4���z�V�a
��삷����"�Y��X|��٫���-�{�-��f����b��r�L�)U�ӎ�����/�k
+�S��nG���'9`E3�3�3X��+����	��t�r��z;/3st�
.�E;���Ɗ<I#��,�W��'2���-���fǣC*�gΨ^�H�&N��`�KW̦e\���r(�{&��15y(ZFagj�5��S�7��ԩph:�*�S�MGWƅ�P�"G���2��<Ȩ��T㶴/��H�j�D���t���h���\�Fw1��q����;y�.v�qI�w0r�V��8`�=Rg/�%�y2[ԫz�~�oz�#�a E;n�Kd��:R���d��v]58h��u���.��H俯 q9D��jQ�xr�Ďhn�f�G�HnT:�B�M6)s���x�>�Ř2�W���s���I�8K�l���KY��l��漚�"ҏ�#SE��W�m���5 j�X۩��VV�f��A��\�6�YYm�ͼ���ʓ��e�c�8�&1C���ӫ3��N�>̆S���Q�+)��7�.�&U�ƫJ����Z�ĥ8s��l7mb4��r�T���or'Cfux�>��Tm[}�-Yn�mmX�6e�y�:��Vwgc�7��Kٴ�Wك��*8&�l�ܻ�3�F%�CKOr����p���=�EÐ��g'4'fT�����R�	�<ˮ�@1���w��y����*�6ـvS�[�lD؟`oVGv�3*�a�2��YC�5}�ƻ����}�u���~PTA_:�Xլ���;�g�i�o]_([5��o�J�G�Ń�d��(i��dӣp���;��1�6:�]� pF2��Y|�#��q�jI��T�(؈]Yz{B	�|1+��X����{��{�#^E��	;#j�*WImD<��F��	�=0����'\��4<�Z4�=N@�9���@�W>)ƺUPg#�:GD\ON�L�Er��VM�,b�y_}w��HD�TUf�mc���%����Vj�}�T]@b��	��",ȗ-�K�*=�ٱ)Ώz��a�5)e6��.<]��Vj�!]nM��{$ug>тͶe�[-;�87Q�i��&�빅�խn'���8�
���f8V�Q�%�S9T����S����o�Ñ��ʗ�ql���t��ki� tr��j�F��dN���ٔ�r�-��N����كY>h[�V֊�:�b�w&�J��ĩ�D�8v����1q`eJU,[+�2a�)&�T�j�v8�9����pZ��Ru4*b�వ�� 4�5�a|�K��Ϫ؋�y�+ڶ,ko>%�j�*��h��7�s���U���DX���=�o ʁ*�0�U+|ҽ��̹�.A��S����S�w{���lJ�xj���&�#7YK���ہ�+�Q�/�m�����tłvizW#��a=�#�h�]Q��a<�X�fc��
}Wn�]v����2��͊fQ�s,pu���+$ѐNf(�X~���m>��9�;Ԍ�m��vK�8��G����0���3y��-B��d}�Ⱪ�Ѿn�����$ݠh�1;�c�o%�Q���SB�;��jt��vQE�ց�x���DA	�S:�������0N������V��t4�J��k����םG��v[vqϲ=`�Ǳ�Jlr��a��Yy�pq��@�;�5֮�5]̶��t�6̹�+��0;`)�1��y�a_4)h'0�i�_%��Β�j�wׇ��OB����k����C0�S�2��FHt��%c,�:��J���m$���<���*]���Wr%��L9SCW���������Y7J��'6�Vcke<�^'w�s�SU�kb��QΛ�!yw0���P�k�۫KL���h��d�;G��wb]��a�5�a��(e�Rc�2]���_��13�X����M�
���[�AN�u��ꮖ��sxw8���b�=�����i�]��z�P�c	r��r�̬����4�|]%�.�A���ng��Wڏ5��hvT{Fؑ0[�r���;S�v��Xݧn����'�R�kl�9d�9j[H�Ҳ�u�}�`y��Y޹!�+��7�n_r�q� T)]�]���<��{��or�o�.@��nS�ꊜ��p.��u��!�#�̖,��	����0X9����W_�&��U<�9�5ø�ޗ�4���6�ެ�&E���{:`��]@�r�3z6���
�����v���|n���44j�o���[
}����9��i�� �Lf��Aٷ��ݦ�방���ɡ�++h�Y5&rݫ�+\���we
� ��[�\i��>Y�M"�����d1&�s^o��7Ȁ�e<zV�7םiu�b��A��p���:��]io�ºp��K��zp�[B��j�3ݫ[W��H(�ɹH�'Q�)�*����0�b����2v�"!� 2���j�ݒ��ᾚ]C�Q9�A�e��N���p%E�xl5٧BA2�� ���+�ƺ���(�x+��8�ɕ��4�#�b&�n�q[�
L�}�o��q�Gf���1m
bZ�}��̔v٥5�ћA�\7�U��蹆��ʕ��t�{o5��[s���ݰ��{
�d_hV�$Lk:ŕ�d쭠M�n�o"�K��x6�r�q҆f^�Qk�ǩ�Y�N-�ȵ��w]r
b����x�1�1�P�:�ݳ���1b�A<��oU���:x�n�(�Ѓx���(-��}k���_o1B�n �B�/,I�efu�Q���ξ�r�J��*��!G�̌*���i��V�(:�`�+/� -"��}���p�kI]�c{�q�+�Y�
Qp�Nf<".3������V�]��6ș�}�B�ݚ�fR��b�mAx~:�P�p⩤X������v��	\�RJ�k��Y;FSVF�J�Wewͽ�}�
��R���û���q�����U$�+2�ړ!��R�7~�X�N��S�YXzf�/%�-�u�|�4���_%�ƑfT���º�b�R�<�Z\��HL`B�X0Pޒmkn��[3vp�zW�"��U���'���R\9��̽=�-�=Ȃ��b�q���J��扤�6�G�M�zԨ���+�K�AP\{��x�-�Xzcz
������k�����toW�f��7MgT�\��Z��Ұ���5J��-wd0�g�lo`8�D�:�9���+��B��f��P�}Z{�%��L(fk����S8��^�h�m�
�{4���)7l���p!��A��<ǒ�r�����硲���9��{z҄�bQ솬�UL�6@M���`U' ;�)^�y�k���^�ʭ�܉�V�՘E�9ƍ��j�t�!�Ի�aJ�-;�{+}qh)�a�A$�U-��y��M�E��v7mlQܱKQۺˌkn�Ԭ�����n؅7Y8�Ævn:����f��;Ĉ_U1�h�:Zps�ֹ�-[����-�\l�+KPЦg/����l�˻u�֙��Ȝ�9��F��������0Y-�@�2�)�T0�\�VMt/z����� ��N�f�Ƕf���a��u�]����@z+WF�Ǚu���*i�т����BM���7!:ah�8cT�$���+e`�co��Rl:���B1Sh�X8���S������h�K�7��r���ޟ,fn�7$[�V����T���\��־�&�����\����@px]5gf\��yL.+�	np�y�ę�,h�O_]dm񚯤��ƻ]Δ�㕚�H�䥍N�4��C�,\��c�c��ձd���)�V�۽��nn�W/VD��{�%ࢲ}an�Y���"Wa=)�=�
��zp��AЬ���U֋pu}��}��h�ʏl����n��1_ao靭�r��]�cb���n7�BX@��ۙ�,[{��
:Ç7m�]���w�U�Aٷ���z�P��v�������J̬ �Ӹ#a/��B�K��z�:�c�vO���iEw$%�Œ�3S4u�)�Ӹmj���uW��fJ2������"l��ʳ{ǣK���`*�t�5����܇M�4���f^GB!�t�����Ff�����ݹ����ںM��|y��,��]}W[�xd��f[U�5-Y�n:w����Y|[N�)hF�ZK�J3Ue��������t�'x-N�[��ڰ�O$�NM'+���{�
C1��w�-
�$��7�J�	#�۠	�VJw��o��xT}�ͳ������}��)�mأ�
���N�x��N\��4��oq�#�t@��6����I��zHݽ:��Yt��nD��Cd
���J
҂��K��7.�ng]^�u�q�l�r�O/�q��%͍]̅\�$Ud�z�1f��[�ٔ.�e�W.���:Y�\�	4B��.��;۹�\ˆ�
�#usr贺��N��+�O�Z��ZûM1�\3sEQ��ni�H.�q���3��u�nսŮm�>;���J��Qzr\�θB2��;>/�̉Ho+��6�����4�����Rˋ7)���F�I�#[�@Cn�^ZU��7lœꭇ���b�At��9Q�0����[�gGτŘ����OHi�s�'|��wr�W^���8��Zf+��	��#�Ἐ�̧���]��[76��8��|����%�*��*;Z��	c_�viĉ.��&��y�עq����C�Jw�t�픥i��QƩ6�͒��j�(��ՙ��w#Ĵ[@���L
��޼��a2f���x͋�W�����(򚱮>T�<3�ߕh�Z�v��udK�T��1޸�8��v+�|�V�����Y��%o)�Z�8l���9�y�f.=|��L�6�N9B�2�uI�+mK Iۚ:�;:�Z����\��nȩ�����b<V�DZ���^�C�*ȣ�`5*Ÿ�� �腪ֹ��72�i��= ƭgs��3�%�4�1���Oe�*�j�Sg'B`.k[֫N4>��z��::Wi3(��B%ga���X�HAz�ZY�/L��k�І�0��w�[�K���h��s�r�b1wi6�PM��������
έHQv.�^�&i�a�_t=hk̉!3���X��o9n�*���Z�;�)��Y]�RЏ��l��2��n�� �+r���w|�J�{x��@z�Z5*�������.ʤ�a��J�*�&Q�]'���}�A6��N���Zm�C�:��5�Xb'���أ-K�-V�oF �ܼh�guƨ��|��L*(J�F����0F�r�δċ1�C���s1�z�:�j��Nj�9M�/k;�:1�c��#�W6�/�37"Ɏ�u�ȾM1��	��kZ�k�l�ْ�� �r�l�����7G��V2�u�9���o�wh !N�ɵw�_K�2�i��v�-8�H�ə��ӳg�B��'ݡA�,Wu �0���x�W���-���Nջbm��`GhW\��]�и8kҲ�A���&���ݺ�5[�$'&�tr�)���=*�Zͧ�Y�;{p�6�_H�D���[ک�=z����\jZ���p��]�dԅ	��F��o-2<#k%���
.J�&�k��^��[���>"�2�#��.�EX�z� r����� z� 7b�H�%�;��y.>�dTgP���x�u��pR�`��oS��o����Z�U��7�"�03w.���]Bpu��z���f\��J �a�jwn_d:�es�t��_kWq2֍�1��P��Bm0c����8��9�R���l]��Ҩ�.�"��]]9�.�oڂ�48��I��P��r9�;4e�Zb�0�ю�r�Xu��d�pL�m:S����� 1�S����/i}֎���}�#\NC�.�����=��g��3�O�N��y�e����8���`�[�#�[j̾�+��Rn�����ݛ��u�2��L�g��ma`:'��.��2H���������ffn�<��r�l
���WɁ/qT��h|�G]��]tu��]H���;b6��P�ULOmL�z�{��ա��p1�j���f�j2qc�y��B(v$U����;��<����{sv���Ӯ��cj.Hb|;t�*i��[l%h
Z�e�͆��Ɔ��M�'u27�:7)�b�@:����_�Z��z1���K7�U�u���P2]�[9���[��������3p&+]���l_Wj�էom[$ƴ�I�q;9.7au]l�ؕu26�q�J�YjK�_}z�w5d7�c�!so�e��r�x����c��T�ɲ�d��]s�'nm��6�2�hP` 6��`c2��Ȣ���{K�-�ju'XA�-CL�͙݁ȯxig*h�����F�^�ve��LU��7Զ�<U�.�eMJ���2�7���E��蘃WXFL�A����E�X;nM�L�;n�!b�2`"+��x���m6C���N�%�t��L�定�V;�U���-��{itQɶ��352��z軴�+m@�S�r^��`�U���αWV�[O����6nh�Ea���4��n/�����>M�s�n�=%�>��`n�hfm"��F��|GgseU��x�ZPA��F͙	Qv�"�	�W�=γ��ʬ�N(�ü˚I��fG\�=ڶ3��F>4�K�8\�:%aB��)X�vj�n��-�+�]�v)A�yԳ8�PV�V, LG;ڢ���H�{؍�yVB�z�bj��=�t�*�oz�b�!�J�&te�eڹ��[�9Y{��lw(�(����+Y�riw�*���dn��h�;��N����Y0�!&�p��a;����0K��y��3V!|�;7��C@�uM�j��x*�gTr@�a�&dMil����{� �q!�f�8BA��t5#si�����&�ƻ(�2j� 7�m����=�/[a�(d��d�����iJ�:4Ea�l�n�2�\Ԭ7����ue�����:'�XwN����Q!V�2��{}� �ù��(���O�����C��s�������:5Ef��@-*WdE�α�*��C��Z�7 �Ӽ����/��:���xN�Q��cwL�M]���Д�o�hn�I׶9��[��Bf���e
�9I�U���pC4i.�=�ә;8C*uݍ��a���Ew%p�γomi�c).H�=JuZ�:�\�8���c9�;��K��-�u{���avV4���H��B��;���ɇ2�,�#�VV��q���E�Jz���iX����We�=�&A�%����»�M]=	����z��SA��Oz��HwoF+Ĭ��i^��P�م�X��6��鯗J5:Pӄ#a�z�!f����nt����Zk7�U9�������Jر7&���Ss��Ft�w����O%\@b�K�"i�}"G����4�#��Ǔ]l;)�qmC��5�av�ƛ/�p�1�����j�T����}R����iL��w�B�>.`r��-^�����f�AQi"I&u�B	05��Lt�[WlZ��c����ӫ3�����G���G��\��]����e#��v���eE?�/��e�*¢��f5�]��o�66[v��e�J�ŵ �G&cκ\78�Ev��vX�鵠��̚��V��)�E3�vb���k�������gmNi��4���%��D�[/�f�ɛ/9:vn���y]2�ǃ�Q��W(�b���mq7L$�5��gsr��v8pG33���+�vc�ʋ)`t�������|-�&���]և{��"`�1gr�w�q��w,�R�Ĭ%�宀�.P��ZG�-��O.�Ӵ���§��I+}%Y��U��9�4��{%�u� �=�r�+s�1�d+�M:|/�'��e��KY�Ϋ_6 T4^(3�C�wy]t')��Gd:7:��o�I/&.�I'�.�r`h=������1���r<�7����������um��)읍�����	2�}4%X6N�o���N+�/,���m`&qy�x�-�u�}N�C��ڭ����c3�Q��_ZQ"S賠͝�a�ʲ�VB���]�Řv��ܙ���a�7lH(�/�&Q��Q���~��){-lȨ�y��;Yws�,2a$�Qz�!U�tl�5��)�>q�:����� y�v�t(l;k��Cط�#�:��Q��s���v2o)	�1�RU�*�B�>�g4}]�2u��ݾ��d)؆ܛI��fvIm���p�+ P�>��e�p��D6�Jb�a�ɕLfuN�̭$�]5ʸŕ2�5�gE��I��̖���Vj5���3Ef]a6���VY��F�6]�qlѵ�h�Y5�Y\�r�L��c�dڭgc�dr��,֥ͬҢ�K�V��2�CV�fgk4��ծ�KIƥ�-S8t���C9
��ʴ�-,iZ��:�T��*ҵ�f�٪��3��6if�͘��mV �E33Ze֍RZ�ck�V'WR�S5r��WV�%3�D��b\��R��)a�G��B�+Y�Z�#�-Y�&f��+#�%\cF0�NMQk�l��EZ���bڴ@�N�ͭl��u�+b$��9�migD�Q�R5K5�5������z�_���>��}|���||�d�B�Jš�9V��],���{�+'H��3.s��b
	�$��t�&��Ҏ������>��os�����{�ũ��/�b���+�o�;,RbuN-�s����)ŭq��&wT�ֳ�-/j�$D��HWά��gL�v�|f�y�ڗ)ϯ�W�A⧨)Yp�NE&����Њ�T!S��V\��OI��3��W��\�y>����)�i����.�6,�n`S5��T��3��P��(�w�u4�{i�c9@y���y��7-����qH�w�׽;3��/�J�*�s�b�񨳩ˡ|��nW<Y3��^.f6��QHP�ɥ��P�gZɕ���>3|��D�3�fy�Oy-�����\��z+Ӗ�����>\ډ��^e��מ�0��\d��"��}�L%�/�=�:*�V�X���"�nߡ��:�rF�M�t��ļ��i=J��8=*�`�PgZ��LT-N�S�c����yu�7\�Ҍ���B�n��Zͼ����k�����w�3y�!X/��'R��Ǳ�}������l���ҭ4�}د���utÖE6�feM�˹nA��.C�,�</\���,(������oh��;kR�WV�M��$�	Ԫ�cn�y�Ѭ\�F� ����Z����7*��u*�b��֟=�n̷�1�*��]9��.����yɶ��.���.U���W	�k#Q�W����L �c��v]!:��+�����'%�:$v�'�OO��rT婷W������[�������8���o���'����2ΪIN��Oc&_o.���UW\R�G'ȹn��OG,�Qp��r�b�����N'.f�� ��FMps[�ZS�·�uw*�T�2.ɕL�.�M���%���a�p����m���d�ב[W����z�R��/R�F�ud^��ŵ7��$l:�M���k"���@fB}��$gp��'�t�w\	GdT')�;A�ʇ>�?d���70�o�#Ɯ����[*�����j58X*#�d�t{�9L��W�����o
;w���0]�`:p{G�Ʒ�^�ɞ$�\-�Cfݜ�5����A�H���Q�1�5��c�*\�b�yl�]gR����UP�ަ�$�hf�S���ޙW���<�z#���Sh��w%�)pݎ|N������M��:����]o�n��%׻V����	�ШN֋����,90ژ�3��'wB������r�����6TT�\��:�-��'�D�A@f���9,mwli^�MG�~��!S��k.z/:uz�}'��.�+mOo�v�;:��i�����ד�Fa�4^��x��:9�_u㮕T3�d��R�l󝴜�\&�ܦ�_�f)���}^�^�}a�p�����oB��a���R�߂o���M���y�n���<�ò����c��3��1�^���B�Rz�|���o��r^��lm�f�7��SZ���zzU�b�<�Z�R�5
���0�ګn	�yiO�yjܒM��:,��(r�+ ���)vd.�o�r�S�}���e�>o�cu���$=
S�^}C���*�y���v��F8n�]u�)˔(M����iz�x@��/ccC�y�z��Ue��ܝX�x��	ڻf�����J��T�8�V�;�E��4of���Cw��ޔ�M[���Y���]q���.U�N�	E ����[e��1��T�P�6�vLmɯ36.�^�/[y�S�.���_el�,�XS"�Ҽ��sj���*۰���n�-��sp�"c8`T{<��<�@.ew��h]2лɞ}s/���fpU�V�Q��vEBoY�y��󭭝@�X`b�.w�y��Xה�Ⱦo��c�޵��	�0���<�b;C����B܍��]'iF�=׌�������Ҁހؙ��ɤDlZ+ZKT{��o�������W��Î�^����Қ�j��*;m�s��Hx#��Z�k8�ۚ���Ͻ�4�y�ݝk&m�Y����,��As�zve;c����j2�ue�jB��{�K6�Q��PasW��r���\)�u%�粡�w�T�:<��!s[q�5��m¬ͮ�5<A�s����*?t���uZ�5��)|�7|�-Y�o�����Q>�/��|��f���H�gU�K�SR�޷�K{Ӷ�[(�*��9���w�"�o��A���.���ƒ7Ux8�j�%`C�)�6��M�k��ŷ��+��AKA��2������Uۗ]nM��NSk
3!���:|�ء%�k�(ݵBsXJһV��2�vOjI/ǥ��J���E�B�>����_������kE�ܕ>u�9;�˷y3vr�����=PW	�Ma�}��J����L���$���}�k�Bj�Gǅ�{|�t�_*�5�;�����<w
�ςr��g�T��n�Ǔ�/vT���xY��
��M��d@]8�[�Z���Yا]y>YΜ�s���y���8O�ޥ��巨S��qhN��m������d�PM�E���}�b '���X��g�I2Q7!s�/��L��s7֛�����R��8���H59c�nS�ZЏ%�����9�����]�X�/��@o7:�(�McRT�y'�?j�u�󥏎��@�ʆ�j_g{7Q�{i�]��u�a>۲���Ov	nz�8K�Trţ�f�:6y�Z�_B�,^��th��-�Mf�cg[�+F��e,���֯ϥ��1G��*)mAET��%�Y�^"j�9;xm�$��}����<�|�!��^����9}��W�1_K���6��5�Ꮱ�]q�tu�
�E�l��(�hMv;9�:	Һ`�,]��7�l���Y���hW�Ţ㼞�)�K�Y�J+/��P��to��m���y�N������#Ͻ����z|�����q�̱�g&�y�j�o:\�����*B��u�/�{�ΈWD�zk�4�˼΁�]�u2�<޲���ٸգYprtv�'Z��_&)jtS���=��'������\}��_Fk�*��9F�T��A�LU�B�s:3nw�O7V��Z��Q���hY֛t]�^��-�.tNs�宏h�ށ��?g&XX�ڰ��=�mơ�I�4�>z�Τ�tH�u�yv_�D�L���d���p-�s��Z�^�ҧ������Cz*u�x'�f1�F�Q�u���c�~huI��^�	����R0x����#���M�����w���1�`����.2��!�=��7�3ɿH�p��s/r���9ڜdt$WL'Ϸb�tZ+��������ѳei�*+I��М�&oݱ����[�s-�
�Fq�ڎ��_j�y��b�'=u�(�E�g�*m�S�Fk��Ӵ�-:|K�t�h�y]] ��X��v݊ܙ��c�"�ř���?)�}�G!��V�ԭ�����y⭪�2u_�2 �z�j��ڻ�D�ry�n#dO��+\��u������(�ܪˑ���>{8�;�t"�S��N/<��B�{�[yq<�hV7�#kn��oC�o�g+%�3����j�a�R��ѳ�/��[�F�^ŷ���P�o��#�B�=�;c�=V�=���y��z�R�bZ�EOP�.��7���[~������׬,�Fm�����s�^������}~�<5�['���ɝk��ڴ�
���\	�_^tٞ�+i�B��*]���i#��M����3u��կk��*a��@�O^	z��z��]K^�y���S��zLp�ks�M��*�H^��iA"�W,v;sZg�3��<�¼�4_>	�����{�Y[�`�*�B.��� //�v�p*E�=��^�.=X�F{B-�1
��x^�����C#�2��x7+���죓R��t�����=S~O��S�hB ��Zfٮu$�kL�y�������Xmv17�n�Ʃ�c��,#]�zf5��l�]��[�:s�Pw�Rގa��=�a>OB��>���q�Ќ��tj�ⱶ�yr
X蔪T�x�k�ZЦ��R��Ʌ�g����b̢�[��)\�z�D��Tc�qA�tqK�!w:�|�36n�Ȏ�s�r�{�e���n�s��I��L��G{ao��L��{mrq��X�u�<ns׽���?-Ly�/[yО�s��ns����O�7����c}�s?$��tҀ��nr�nnE�P��������؟b
=-z�o��[X��V����vEy7�Լ�#�5tШV䖫ޭ<����Qz�����/�~K2c�޴�<&;�2��+S�a�vnf>��V�G�,�K�]���=�|��v��'�(Ш���|��^�@���<�P�<A�V�~�����_�̸nx�¶���߄yN*9��ݾD�n<�r����~�[(����Ҿ�A�٦�CO�EH��-_ff���ed�p	��Z�p1̍v�\���mm�R�=kft�g8���X-ܨ�(Vu��z�zQ[�#���ʘ�-48k-��e�4]��I����t)��,Of�vu���|a��5Ke��e�{/\B��M���׼{����n����m<�W�^�}�f�{�PVX��57�Neۻn��N��^k��)�\��O�E7�j�*i��X��s�4��
��������|
���Z�D)|�7|�-R��#gdin�n��B�]��X��ؗ4���HR����	�-�Ѧw+*ڹ=�r�ތ\�s�.˨6&���<�Mbн=�@/!�;oo6��˺-�m�[�l��=������r��鳆�Z�5!<��T��N����o��:�Yx��}�T=��D��^1�6�S�f���/w�Ժ�"�vz��gd;u�n��<���dsW1s[\�h���q����y��ϵ�eV�Y_7��3;��M���"���be�5|=��ur̥�o�B�aߋ��֜S�xm��S�Q�s�%x�܇|t�C}���3��K�a�#fŪ-�}>�@��PU�v�E�L�E��{�LE�K�����4�-a�V8��*��4a8*${V�耣vc�ҏAQ�	���u�E�_��oI5��tO���{7�����ƫ}p���r'/\���\�/A܇�
s���VE�a�f��\�d@<>Y�������nҺwl��9o{hշ�w�,��0��@��P��Q�;ٺ�����8�������Bk����mU�N�߻˝����/<��]tԳ�_��%Y���ɶʝֻen��~[���	�Ƃv�mO'��f�Ad�X�_JP�)���[�uN,i-��LVN��l�9KS�P��V�6��{�^�����˧�8`$��U�}�v]�����Ί�&���M/w����F�#���5�g�w�浹���zk؂�R��j*/�S	˾�-��iZ��VfcG����T���	f '��eV���g������9PNZƥ� RŬ&�ޅ�i��F�(E�~��˫1�q��U�E�]k�>p_M��iE��?L�b�^��`�&���f�e�ו��k9��,-��_^�1����,�C�N	���aJ�u<�7Ub7́��S����n�p��d��CӝF��5{ޤ���@
�<k�T'i8��6�K��ŵŉ��ˁ�2�貱(�����W�2n�-z$$�v��6O��D�p��dދ�p[�\N�l����H�{J��� ;ݦ�K=[]1]1�騱�C�s�V�tcr�ۘ+���vf-��T�#�c����6	�VkoAD��ǥ5|���^���$���	�ufj�be�Z8؍�JU��۴��+���mQ.ȉ��>���70�Fc%��n�)��G�3�F�_Qؠ\n� �����V��$4��fm-�$&�$5������q�(�meޏ����ܣ���(h[OjK�������1��tY�/�U����q�c>!G�vG��Woȧ8JnLt2��%���sD���V(.�*�t�%4��RgҝĚA�);*ھ�+��j�U���F�^V�V$4���,:�wAv*�U!�v��S�J̙Ҭ_o-X�����B�<3��e$і�.t��c*�Yf����gֆ.�M�ӝp�'p��ZV,A�E�uZ�T�AbU^Ѱ୧�Wj1|�_JȊ�Յ�6
�4�g!�W�m"6;�S߶\��"�u�ds�XΝ/$
��̺�v�TU�{�c��:�WD�P���f�]�kwRʖ�e6���u
����"����c�z]�%�/]ێ�U:�]�3e[ֱ�z,=[�㱺��*me�*/��*�z�;D����Ԥ� �}h_��-��Z��/\4G� E����_��_K88ݍ�Z�i�R���*�)K+%�I���>��:�Tǘ�3�*�ޤ'6n��
+�es��h��n��Q�}R�r�-$�u򳼚|#-e,�)n�N"�byT!�I��mV[�M�#��cM�/v;x���D"�]O����Q�+id����i�K��Jw���� �gV��C�عbY�{���ݬ0mv�y#�k8;j&]*>��������N�9��d�z�ΆG�2�a�kiaN;�Ywe�Iw:�.{\��ջ�!�b�an�(̏�
2���VP�:�� �p��-}j�A���N�K�ty.j\���SF�U��l��F�Fq��������J�\Xz�'kt?�s�엻y#�c;6�k��fganj�gJ	(�[��/�F�sg���_r)S����%�6 ����i�+��r�c�t�����K9J�JX^�Йb��x�ًMD��ꁽ�Nᘏ=0���ӽn�Y]7j$���6��є\Pv��9�rs�jsT%�$�.�a|3�C�\o�!��ܩ���5#t����%,�l@g�c��ru>��B�95�|/-V� ���R���o-(`�mUVֆ�Euib��N�Md�Y��­�����5��ԥY����U�겙�Me5s,�N��V�6�K79�
�Wq�gc-k:4��+r��eY�++�&15�cZ�*�Ltӣ-F\��vY�*�55��WM���I��֮3�V��9�чci����dܪk�Zͅ�N"�Ӄi�mlY�`�hb�5u�]�*L�*m&;NZ�5,]]v��֢Т,�M�2ƫ2��QeJ*i�u��MYL�Z�����i��+J�du�Xֲ�1B�s�KN�U�1Z�b̭͕fm2E��ƥ���6���YkI9e�as3
L���er���$9��̪]q�bEnJbV������w9WKYv�6��%h�5�R(P�_A�E�Uv�{g^n���ae��NL��.��\��o9I�5Vs]$�v��YsJ�y9�6�;��=��{�������1Zs����-���Ԟ���+������Bt]@c�Gk����z���Y��.���r�t;��+ޝ�O{/=	���y�]��3T���/^�Y���O���k�Tx�	_r�t�#P黫w��w
���)z�d��ܻ�����!Y���8�Rs��r�4���oBsR_jp(�\l�)Է6�ڭ��j���T'�s0�騕�l*��պ�{�i���b�b[ (�;6�J��J��Q9	�f��#dLj�?`���.ל�`�W4�J�}<�+|�	��Շ**�Ȥ�%;�q�p����̠gw�hR�]泴��65��E�u{Y��pg�P�+�2a;�Q�;Ε�V�*�<�y(�U�%�Nu7�~�����	�4���Ŷ�l�_3v*=]��h{��T���O�XZ��QQ9n�8�Z��C�WnnL�;�{Ge.�z�܄2��ko@��f�+-L��;���E7Y�&V����������U��r��B޾��
��6 �)��t��ޛI_f�iD{��f>IH�hn��RL7}y|�^�"QgVV/�ܤ%G���ʣɭǘ{�X[�?Wr��i���P�y��e��z���>(z��u��u���I ���n�2��1<��mp�}�����dK���O�#��Q��6�{��:V9���[�M�ڬ�HNQ�t_
fo�k�UR�n�^u%�s�^��'�_;���z;97�����;<��M����K	��ҝϷ� ��gW����k-hS�O]�'���Y���z8���n�����k�k��#�Tȳ�W	��&��)�J/o}=�k!��9�Rg�M{����=Q謝r��?h�ٳ;j���;�]'����q�W�t\��{Ȭ/ε]_^�G<.���O!�-��*�zu��6���^��K�v[K�k�9]�n��*OsΞ�����F���u�����5�>�Kx*jVᷮ�{|��������}nӨ}���f0Tԏ�t�+�rk��lh�-x���Bjonw��-�հ��+��Q�1�5]P���3��	)d�	lP:
���Uw��6�TR�!�<�PЊ�����grQ����5Yt�̾D	6hޜ�(��W�{�'i{$l�������.z�ȟ̇۱���\Üo�{Nn�I��]gr�im-F�{��\��Y��,�M��zОP)�0��<�o/-�ҫ�5>�T���4�ƥC��<b㰗�`f_���@w|�&��V�����NZ[Wp�b�~�8�M{�l@���<v�����.�g0�}��Շ9�{y���%-���O�vj������~����3���̚���f��*7;a�r�.u�Z
�{��j<�s>�����B{s���Q{�ݾ�ޞ���b�9Q�Wk�یi�Ȧ�nfX�﹇��M���j���=*��J.'[���HT-M�V��Z�ў��Q[��,���{��a��C��J�\I��?A�̛�����p�q!�y��;�q��߹S�N�o'-J�N�ηi��m-<?=Ԭ�+�P�Ԯ�V��y�g��R���Wr;���Η2r��ĿAI��r����e~�q�9���&���C�7//y���}�s$V��0}t@U�Lv�q]{3u�̱����*[+`ۡ�u���M-�H��u��,�{�"վ7T�:�@ %�f���o�/�ea*�Ƌ��]���ܓE��\��},��l.^���>��,ZZ(���r��;����U�������E=�?�d��e���r[���$w���y�����es&�>`��PRu�	�>���L+�7=�5J��ώ�:�7S��Fn���A���G�f#��]^��a�9��M[�̽��'��n_d�=7̣��^Ú��̎������������u'X������MȽ=���oG�<��C�����������j]��;�r�p�jM�{!�5�dո}�P���_d�9��z�{�+�;������޷C����݁Ի��Gvo5���<Dx�7��0H�_g�>�+��xO���O�e�!�Ԙ��GZm�����7��w/�S���<��z��'��]ٹ���aR���� {�">{�K��.�C�u8���w/���̎�>�O0ؑԝ��q{)��e܎#�}���]V�f]I�3�y�.�7������n�7��>������� ���{�ԯ$�y���b��nK�0�y��_�����܆��:��ܞ��a��{���s�\F$�>ח� L����
]n0G�z=B>nbǼ�R�yJ����dJe�|�^I�����W�k+K�0�A���>^ǝ`�r:���>C�q�x�WyuF����i�Z�B��D}�r���<@u�r
Wѭ�仂��0C�}�A�`Je���G2��2����5����C�M�j/g���x1����Vz�_{׹��y���S���y/r{����Լ�����7o���)\GF���w���2���q���=��{y�z�/P��އ7�=G;�^c|�W?��+9�x�~��z#������sްè��{=K�9��e���r/�nϷ��ܯ�ῲr]� {�}�r��ӛ�K�}לǞo]%����ne�7����]������H2�I���u˱�oA[��;X�����dIOvӼ�oM@`��R�R[���gB����X!ײ=S��L�"�a1���-D�`w*�)��F���;�|T�4�F�W&oỲu:�--� �^��[4�I��>�C�y�ՙ���Z-K�w�;��1==�9�z���w/g�_`伂���;��:˸�W���r]�=5�>"�T��FWU�]{�!�p���󿲇��כ���a�����>ϙ�>�R�;���8������u�C��
^������v�샸�����\Mz���h�Wk�[g~��w'1̛���>�M��~�/��+�C���ȾHnN%̞A�N�2�7���G}`7+���n^A�=��US��Wm���w}�b=s�����%�N�����<q���w�>s�(nmK�ay#�ٞy��Bvc��_���9R�;���"�v#�O�&/}YG�-^-�{��D\��3��F$:��u/=�xo쩉w'O{��������:�#��YCP�j_9�zL��;w��\��N�a�A� z.�va��Jߦd���)o%��:��b1#�w��̮�A�~���0�R����rk���P�������ja��0.�y��L��>z��S(�}}u��m|���� D{�g܃�'N0��Oy0.��u�QԎ�}/.�=�r�p�j�{�7�}j2��r�'v�����l
=���MV.y�G�"��d� ����29����K�Ľ���u8$w/#����'��{)�0nC��jo{#�]�o�w���z��^��y�}�^���|��'7���/�wy�2 �^�u�AJ���ޗ1����b]F%�8p�.�����zy����xMC��Ow�^}]��uׇY�ލ��5ϳ޸u!�wy'3��I�]���y��R��}���
re��^t�!�7�:\�!zO��1/א��~��`�#�u?bw�=Ƿ���i���V.:��ip�WY��R�CY��|�b6쑨��W#mcx���zD��jB%2�S�bf����Xw|�������n���
ˁ�qSɣ�ё�5���^M���>�Zq�ֳ�����ޒΞ���Q�r��>V����2�n�k��(G�B#���!�O��ܮ#}�����̽C�(N�̥��
{�2%���y��/!�y���bG�f�4����Ek�9̝���u�y������_���8u�}�����awa��y/pv{�y+�Ě��sz�yy�;w̥��1&��(|���Ξ�s.������\��z�Zֵ��o�{������8MHj/cǬ�L�`�9/p�MHy9��k�rG�1&ϵ��R���7���1)۾d<�r�����k�Ww8T
n����3����,�^��{��+�������{!ь�<�ˑ�XN�܏Gx=���;��p�AԻ�Ϲ�9'����R>��|���Nu��y�_{�;Ϟk�u��|�Jp�ɹ~���o(}.���]�Լ�̏�az��������_c�xNI����;������p^o���|߆+\�Xߚ�ߺ�:��9��j{���dܻ�Jv�'%亾�ӽ����7Ϻ�ϼ��f�ߘS��^�8w+�b;�pP���w���ѿy��{��ϧ�k������@s�/�j]F'>�C�>βn{�ܞcY9.�d|�3�C��};�W���}y�|���q�hG�z�O�=C��Cp�W�6lgջ__~k���8��O=�r
=c�5.�C�9.����w ��Yy�+�<1�����<�����u�ey!������=�������ͫ�:w8fO���n1.��x�n��vgaw羰����xM˨ć^`u'%���*b]��{�ϰ�$���r�{>�>�b=��r-�}?Oտ.�>g~w�}��s+�ߝes'���C��1�5��;s�2:�q�u�����8M˨ćG�˩y{���#�cЭ�#ޑ���?����wtN�Sj�Ѽ�?�,�'y�K6���$�U�p�%\ջ��Us-�	�׊t4'kܩ߇oZ�S��{�a��Jw+�HT��Ů�N��v�:�su��(J޽��%�I�ռ�l��'D�t�X6b���I���׋���wC����+���^�
�G��}��~��{��_j�<�Kٿ��3+�w���sѬ<��
CP}/#ܘWP�:���Gs�9.��=g!�ë�;3R��T��ꛩnd����GD`�|ky��.a��y^G%��y�~������3#�;����������u��������a]C���	�a]�n~��@��Pf��ڿ����D�1�Mc�5��o8C�$��W%�M@{�2�����y�yr��΂���\�@����1/Y�z8{�P��nm#7?/�n�l.Vo>�=���p�	�a]Opj^�z}�]�r�A���J���N���s�OP�:�y�}/|�΂��;�y����3�Ý��𭡥u�IЏ�1^gܾK�����_���w����0��={�M��yo��䜕ׅ��K�(M�	A�|���� ���}��X���VPë�Y��G{��Ͻg;��Wp�����3)�G���aw~a#��'g��p��A־��9#�vo�;�pQ��6~߻�q�q���GsUc�c��A���R��~�y:��>�Ͻ.|¼��V�W��nCP�{aM�y=�;�/�nd<���>���G�1D_5��X�wS_|��T���]y�}�P���MK�(Mo��_c|k���z}�}+�{�=�s��������=�ǩ��w#�{=��F������Y�S���P�-����`�u�|��>��|�{�p�q)�9��u/щ<�2��/i�{֥z������u�vkC��Xǡ�G�{�9|(t��=ە?5���/�y&�y�c�~���0�} ���"���z���W���y����ܾ��ְ���s޵#�5�Q�$G�B��8*�>�}UVv�����yU�L���	�f���/L$U�1�|R,YR�4�{���e��l��U����Z���k�U��`�@hK���Q������b"	�:$jN�V)�eK�/�8�u��$���b.��\�#9�[�Zi��Q�>|����?*���w��}ߞsz���n^���w8���nMH�w��R�
^�0�n^F#���:�rv�Y7��>�^K�����&�仾�Ӿey!�~����&J�DXm�[�߽�菝�y�����)�u/ӉԎ��{��P���%��j˸�ke��7��+�5����󻇛���������W-�ή_�!{�y�=�Ⱦ�y�D(~�z�{���Rj1.��s�=����į�~#2n
GWRnN$8���;�q��~�LK�>�ow��yҊ̉ɓ��^�6�ۋ=�1���B=�䏜�8��>ڗ���Gs��Η2r�O��'X����w=����}a9J��3��:�H[3����ٿEw՝kL�ؽ�ZS�C�cޡ��G}>L@j��W�9��{��unGǚ�$w����t9��{7�}.dԧx��1.���P}/#�Ʌu&��s`K��;SY��o>q"���z��ϓ�`5.���沆�9a�2j܎e������G��Q�w/5�G2;��w��
Q�1.����=�����;���sy�w�pC��G�WRrz;�}bWq�w��^{�;�r�p�jO]��>���[��~���2����N�ÞeOp�d)^A̟c��a�F+!��zsj�2�����"<���g��}���L#�~���]ǯxO���G�e�!�Ԟ�yC�v[��{��o��_`�޾|oa��@�=�|oq�3�ܯ>�����^t� �Z���bV��:�K�%�]]]�a�}A�I����}�r8�I����<�Ռ�Y:��\ʭu���?���+��T���7���_`���� �^Ýy�ܯ$��}�s������!ٜ��^]]�`�j:�������$|=�{�d�?��V�s�)ż�X�1�M�Af*�Ffg�Ԟ�R����k(��*YU�e=��Y�������� ߻��.#ѿZ��2[̏�:�o|�a�w9��L�^h[ƯsR̝�c��M%3�/,W��|�:�UJXBQ���G��6u�=�_����<~u��ù��[�ܻ���|�Pn_`��\Ȕ>����Gr���y����<5��טC�8˨|��:�;�>�0���p��Z��4P�1��ac�~�ﱹ\N ��d��#�[��w!�`<�p�8��\Ȕ?K�;�Ԏe��=�s{+�YZ/�%c=?�_���֪��I?B�{Fq�
{)��{?Kܜ��ac�wvk�����d��#�~�仌@�o�}�p�8��\�����^��^�Df�7�_�&��&�rJ�zGG�8oC����G����`;��=ǳ�y'!��/�u.���"���>�^Gr�����w��|�R��}�����u~{7��i�Fj�9��U��^�޵#��GVdz�ah|�/q�p�W��������:�pR�y��K�+���:�pw�e�w>��}������	�����G`��)�MK�w�׾ee��o܋��y���=���g �K�����8�����_d9.��C�x<Do�s���l}S�k�R�#�G�z
1�ԏ�qƲn]���7/!�Ի{�W����}�о�v�jq/R{%<�˸�83+��ް����LLM�1<\��g���[N"G��菣�{p�N#���1/$�9����<������Ϭ��}�/����#��Η0����'�v���wug��.�gDL'L���������uF�a9J���q�|��K�po쩉w'{�����7���܏�5eC�|9�zL��;w��\��M���6�2l�b��ٯ���D�!q��K��bGP�=:�j:�Ո9.��=1�ܺ��`<��S�N����B�^��NC��}��|������j��2��B�;��ܐQG�����pS��4U��3"!@,�~Q<I�w>pj'pP��Og)����b��{Z.*A�U��V�C�������Wx;^��sk�:�*mf�Sbg6DW v���Y���l�	N��´P#6m�J7����]j͉������G^S�z�����D�{�y�LzD@ �:��'���'��P�;�Q�ϦpK��N�����>ڃ�}dO�9'{�un2��~�z��#��<�~��뗼g�~���<ȼ�����R���}�C�(�a��Q�z3�7��pH�^G��V!w=��>�J{�rnC��jo'��9g�箹��k�{�ug�w�>����}/p������/�wy�2 �^�ם+�7�2��H����1.��� n��X;��_��0��#�;5׷9GX�~��W_f�Z�G�cގF�B�=X;�r��̝K�}���2�K���eNA����΂��=�>t��B��7&%����r�/:��7���~���Ǟy����wߺ��G�<�w!y~a5/��N�}��q���d䜕��9�pP��R�R�=���(}��|�^C�y��bG��3�������]y�������߿o\]^�b^��`@jz�w�����!��^�����W�5��J������Bw�e(7/��;5̉C�:ߘ�7�n&�ɣ�c�JK{w�p�zG��۵�H��r��w�'$5����f<�K�;�Z��R�}�H�$�X9+��X9.���ޱ���{˳�q9㹫ݨ~���7��mJ+*��O��׺U��j� c,�(�e�\��WS��	:�����hg�n���
�1MMd���]�U��'�;nm��o8ײI�=��{���jV�l��zǝ�j�+��.���VĶ�j�I0B�0�1i��[��i�ǭ�/6�m���i�z~�dW;;�3�������T�i�j�*�G+��WK7We7�!��%9��3y�)��J]+��r�X�D�ڬ����;��^R�VV�iB���o���j<6�ܷ�g�:���F�
X0En���c�SN 鿫G!�rM{��U��:[F�#�z�I�l�sr��@%�u���)�XhՈN�\E�fr��1�}4*|o�)�l]�9���V8p��d6���V��x�)�Vڥ�ʘyC,ϬD�V�E�e6�i��q�l��+�ą-nm�r�+<1ٳ�M���D2����o�O2�GYַr��$��öm��~وt*<�(ӫ�8���d���p�ưס݇���%�����i,}��:��ͮ��}s���Q)b=弅\����N�����^[��M�	XV+<Hx�W�ZZ�'T���쎫Wݕuv� �����^r�1�n�[�m��ɡbZ�-�X�^��L��^a�9��f�_]!�R7��6j����h�ɖ�*ݏO6���2��;P�D�w&�y���43~\�LU4�N�#�����K��[�Z�`�Rj�t�VU�2�jk&�)\�8��p,W��[<{���z�(�o2�,=6.����2�ٽ���Z��XU��a��Dr��X�h�lTl��0Z�K���sq,�%� ��+���=�¬q
�'������:�H�r�K4����kiW����><��8�H�ZnK��2%�4�F([�;g5�͋5��ۘs��w���{�1PF6�j�6�ˬ�t��Q���ko^�����`��h,Z��5l�&5��+b���G�#q��ʋE�y�r�����7��c�0�1'W4�����ذ��U�ʲ[���N���vMV�M�\��u��;{u���J���U�E1)(�����@�������9qv��|�讹\��_^U�s5��;�3�n�p�=b�&?���et�Ix�8�k7X�OdΙ����ڦc����Fk�ڎwfUY|a��S����f��fN����_pw
�+n�ߧ!����+"O�P���:}I�C��6M\4+ٮ�̙�#CiYi��P��`�ҷ��ޫW�^"��N��G�J�"��]�x,ꪆ��ЭORW �a�9Tj�7��y)4��=�o��70��V�$Zc��MU��m#�g�6�nв7x�jy�IKm�Z����;9�KZ�˜�I�T��gj�e�w�^=�a��U���)�����hR�/7Zә$�LVeZ��N@�o��r7�`�L��Εz�+"2��f}��g^L�u ڰ�<�k��i4�Kj%�-���λ��39ˎ�z��Fm��G^���Q7X�ba���j�����"���o^������-]u�Y�Y�S,�����h6�Ś\�\�Xj���JEs��I1S���j�VW]�\�53M5SU��,֑f$�j˪ıjfiN[\Z��5�k9uW\8���
���KR�jubQ�c)k5�KV�MU5V�Z��wM�vm��+j��Z�f\v�WZ�5l�Ղ�*u�jQ&�+Zj�Ĥ��V�JεYiZV�]����V�k.�,+\�����%;1k1fY�mR����u�6ul�I5�Wj��k&�J+��d��%���&��2������kV�Xij�\�1�lΌڮ�WY�1d�+�j���2f5ֶ5�sht�LF��f�Yl����õ����33W3h�3��V�]lM�wi��,���j�ԵA�Z&�eZ�D��e5i�ڵ�J��*ڥ.��:��U;Z�,�Mf�-fmfΝV��5�N]U%lv�I��O�G���b����!d9E����̐z�j�D],�[p*�N�K�{k��oI�n�o^Ť���8�y�W~����^�o��C��b�5���*V9�M>�M��*̠$7�
o�z�o�Yu8���鹙�)~+D�A��*"� �>�/��M��=�p�ݸ�x�,��Vu�s]�y�7+�OT���LR�|��Ц��	�Mo� ��)���egi��.�N�wv�n�{a=3���T�94�Y���l��n�n�����뛸L.��ul�Ȏc�Gk�1ʸ�/�Z�ڑ7��d^$���X�>V�t�ջ��e�=�����sH��ۍ�z�7���J�k��mb	_t)ܨ��;!ۭ��;t�B����1�v�����ԱZ��֐ٓ�ޅ>�ᓺ��mXr�9^8sp��-x�u�,�ž��d_����s7<����%��|}�umw�*FzDV~�2��2�3z<[掠�me!Þk6�{+㫷�}�u�^�Ek-�P�H��Lfj#}n�΢�&0E�)��r��.i��u����D��^�a^a���X��eN�w@',����6n��o�b�Fa��[�we*�:�\�wd=郆����	Z5�k<����g��[����:���������������n�lu����K�#����g,�q�^q�_��h;�{��_�sQqpe���Uumw�;5=M{XU<���/*�
9�����[ۅg{��t�*�s^�=K���(����E3iry�P<�÷��t)P�ٶ�s�M^K�e�W�A�K��Zж�gE,�ﳧ(Ɲ�_k��uk{T�l���H�0�S�\	��W����ޛ����l���k�CV��%���+2���<��'[	�M�B_�܅��/T��z'=���]w��=M��Jª�9*��Q��������9�����2�qϟ_�|��{�� 輁�b|�'UK��4��*��V�yܶ�>���[э��N�|S�;Kh�:&k����iN0ogǁ\�}T����'���[�kηV^&������?{'ox쳢'jnq�.�+z��|a�T�e��75�9$�GQ���y�V�ܬC�)Y����(u��{oƩ2��=͹�s�[������}{��1��^b)���2S���X«X��;�%Z��0Zδyr�K:�%*9�f�℧�yG��t�(�j�{�Dz=���5]ؓ�;ʸF���^TG��N��O�vC�[N�P��an�R|�������޹yC�]s_k
kFLjy�{6�s�~�W�<�	�rI�Iq��fSSg!yO�^|9�߳�QW6�2���hw�2�X�u���}/��XR�҉Ȥ��9�w��]x�sR�b�p�{y�u��U�S��@V㖁;��r�S��\��y�}sqS�^~��ǝ5�,/k+|�>��G|s,���@Ns�1ɨ�O��>�tj9���O^Mk:ݥ+/�kq��uZ�Nu>��}ۏy��XЯ'�E�<�n�#i�Y��3��A�]{�.aɭ��Um)���6TTNZ�ju��F��c__��a��+S~���יc��:ſr����/ާ��Rܧ9m����d�M��}��1��Q����KU0��w����֣ES�w|q����.����."���r�dj��m�{�'n��x!�z�i':nh[��:(:�����\�[M��KRKbk��K�Sa�/��4�yۡG��[4,���8jɗ�:er����cF��^ŋ+��YU_z=�zӺ�\5�jH'.9���Ք�m�̨��r�ܠ5�=9��cT��w�x�=1z�;�b�0��a5�B��ۨ.ˡ�q݀��3dg"v�;W��T#�����X�OM4�\>�o���M�k�H���u{j�4�O8lH[��yT���As�Z�-�J��_^�D�A�C���On�q;��nQ�F&9�]x�)�t����8���7zf5�� �Ve�ێw��}�R�k��U<���eD8L�Q�W[�ELS��ZP��c���*]l�P��4�iS��7
��վǳS]���6��nq|e\���1�۫
������RoY�hQ��U͹|�V��U�ɺ��j\�s�"�mf03����N;"�8Ʉ�z�Q���l�����m�A{ys%���^}��l�*�OA<#,s���+�k�'��ԍΆ�@��a����i$2����m�X��������fJx0��� ��T�׷�P*v,t5oux��qo"�k��m�6�wG�3��IM-kt��Q�C�6�vK]2޼:���6�v��Ŝӟ����>���T9��������Ҟ��УY±{z輯��U�o�&�T��p�'���߾�\�Χ�ō����QU�|����=Γ΢y��!�����l��zIJ>�.mw���)���?���W1M4�w'�����������9κ]]�$�x��R�ۄ�v���ͮ��YL6Y�g�=������\O.��lW�9Q�J9���[�M���F�aTA�̼r'q4��AS�*]A�)E�u1|��X�)|�o���}>齽�m[��M���q9��������K������O�=n�D�)e��o{o�=wm�yֻW���p��Y����������T�O/�g�v�7���@r��x�C��T�B�ǅ��^�����jg2f�1���Qۭh�h��������M�[���,-��4�`8�/jdj7)%s�U'�8����ժ�ޙ�q0����?{`N���Zwiݙ;"+-�����k۸|���g=~�e�[]գ&0e�
-� T�e.��&X9u=z�����=\���ռ�M����0L�ͼD#6hξ�D>9!�t���}�}�}�հ��ߟtv~G�1�p�_#���<��������"�B��d�l`��p�qw��Ԅ�Kܾk�N�{�⭫����b���Y{s��d[��a���݉h�Ɓڧ"V��g����A֫}aJ�Mmf�ي鵪Y�}Y���c�Q��#ٵ��Mo�w�O7W|��\��o*��
�97~�E	����y��~c�;��<b㿒�oi�j��*A���ݼ���U�n��j)<Z9�[�=�5���qva��疷��������ձ�ߤ�-����F;���z��׉m�Z���f�*�V�ٯ$����}˭e�'����,��`>�G�P
�gB+��wv�ͽnXS����%Zy!S�z�\<�5�6�U��{bn�˛{N��������[y�Õ�8��Ϥ*l�]�W�q8�#F� �v���s�a˩�{�K�O?`���P<X��y��:62!ϼ˩&�'[�xn�O�D*X�\���R���a]&j;��K�s��#���]IW�;���eT0S���O:ưL�wu��"�2�2J��K�e���X�GY!6�?|>��>W��;mȶ�n��r��ԵdS}��XU�㒨�eGdE&6��oZ&v����ݪ��Cf9>p�%�,��Te׆��UA:�֓մ���s�Xk�ZЩv���|S�:�Ol:>��b�	��.�띎췩-T�'5҂����}έ�5�:�Yy	���TN�����զ����]	��3yP�k����:���:�>Y��n��s�Y��/��>�Z�;5X��k2m��s$��0�}k���y�9�yo�ǟJ�_���.$�-��]Ӑ�=�7	;#=�pzrVϢ�t��f�1/Uf�vf��jD�ֺW��NBo5�Ӵp��:��;�\������;'!��~�^��Ug'4�(���ds�N��p���Ǳz�(���t��u9��Nݛ�ꬷ�Vc�@�t�
{&�>���Uz1h�3����R[����sl9¢�";�A>�kӝJқHId���6���<�ţ��+e1	���<��T���ؤl��SW�ƹdu�WYD��?L�=r����f��iV�H��%�1��5���M|�Ž(;*��e=!�Q��+5��:�J9Mo�����\��&����� �<`\��<��ny�nz'������T;�+�˹��Y��1b��쬴�f�j�_��n�׎-�X�e�U;��#�H��ZM��sk����k����a������O=�V#�z����7�M�P�ӝ̯w���oܳv��\�E`���I�ʇ���3ј�ʞ��p�������4�Β}]/�Ĺ��P����J�s�JM>���pbs�_4;�i��	�z�&�t[yv6�P���OkI/�K�R��=PW	���hT��i�>�Fd�K�{�(�ƻ�Jo(�1ў��O#ǲ���hT���c����5z'x�8��t��w��uP�S�1>�W+/���-��A���+2g����1L���qN�m���B��l�,�Op��<lT�T'�.0�s��2*�8�g{6��0�_�!D9��O�e�'u����]Lꛖ*4��h�;�v�-�������޿���x�-A��#m���6�1�ٝ8Rӗ3�'<@tFp���}YY]N.��=�\][b^ǽt�h���ܗ{aT�pZ/aΙ�nk�ވ�z==�����=�^����i����~K��B{(�x�o[��Ϋ�4��"��k\1�b�d���xU�a��n'"�{P��D=����f3�_v�E+�ԅ��t��X��ڨ�@LF�q�\Ø��x��.!�r����m����e����O�~��w��	�����cU��=<�?b�@쁕�*�y�N|�{K�3s�T�eV���j��g��sn9�{�������s���.VE��i7�tLc��Boa�Nj��<.�S񬪘�p��j^n0(4�{s[��(�?WTf����H�y(n����y��"��6�U�ٻ��Ml9ΜƆ�&Ud�Y��%eyU�/�prc�ާw�2��x�㶺�v9Ѣ�Li,��D̼����e�1���.�`/����`��+Z�򫅁:zX��aQm���=9:>y�x�<�?qn;��R��C?d�`�x�H^�-��X��/�-����_���D��x{�V��K^��U�iw��]�^ۉ�ח���Ow]�j򷂩��R�����G4ȍY�:���'iQ�br�jq�T��,v,{�E<ײ����]i��&�[<�f���	�X)a���1����=��ۊ*�n}�z#ѷը��徼�W�h̟S�ƥQЪ��V�Ω�\jQ8��^<B`�Ϳe��O+�\�{ues�3τ�S��Ԅ̂��z�z	�ש�G\D���5�p�Ƹх�������zyх����C6��71��g�s�J�J"�C�A�Z*���P��Nn��7�1�K����-�;K��\��r�]\;��7�M1o��d�j�&z�6$]_zs��D���L*1�&��,-�RtgyO3�q�1B�ܻ7�*4(`�������-�KmL�H�_˖�ixnU��ZM�Xx{5Z�~��1��ã�/6a<:����9� ���{u�m"���� g-s�o�]Z�xK40��dxs>�NO�.�w/7�����v@o�V�e6��2���H�ժ��x�,ا�%�&��N�i������L�}[רи
��P�J�o�����ahלˋ7\O��Q�/#e[�tY�+�Z�-؆�?��Ro��`z�õ|��:�\�0;R,��E Jn�2R6A}Վ*����^���2�ҙ�����C��q��|��s���Ч.V�8�9ԅ 7�9'^����0W/�uu�#�����)a�;LB���D�n9)��� e��^>�O��ٯ�2+��eal�
V���{�[��y����]��W(GO���$l� �Kӥ����_:����@ʹ��-rre�^ŗϓF�5:�mޠzW�Y�N�`*�٩vAÈE�z�f����v�¢4��ԋ͔5JɺC��_T�:�,Ҹ�j���!5A�3"^�GF=�.�4&�(@yb}@���w�j�k��q�1�JG���A��u�#�1��je�c��˖���ǟ-��5�[���d,�Xo{�S�.e���.J�_\�&�\؍�<�lH8C��u]3W�Ze!�GPp�?�*�.Y+��A��p�w�[Bnlm��T2���su�d�ض��e����*xo�'eK�9�R�e��sT�u��u95:�/]o&��V1.�N(��PҡV�a�Vz�8L�n]��Cq^��D#�M�o�2+�a��0��";}s�3J]�n_�Cu��pn��`͐#�����ƛ�@������s��ol�9ͮU� �+:�AkQ�ѵ����F��Xqk�v3*yܣ��on����i�@m�mY�}F#ƣ�[3ho�6�݌.B�ǒ*YP��9��s6]�y[\�X�����$}�:���oA�+C����Ҁ۾���4g�cLR�l��n�
ء��<x����YkJۖ��K����d]���F-�JţU:�jLΥ�l��Yw��e�#|6��k��r�:�0�L�%�Ȉ�N��K�����d�Ňt��#��/zq
ӊ��J�l3������˰��pEopq��Vd`u���p`�j�|�f�j�Y1��]8�{F�-���U���[�1b*�&��=ȵ}�c��/x��-�^�6�"�2���N��=y����������J�)��X���{�Љ4Jh]Z�6�̝��R������Vm�'Ewf��ĝ�]�X�ΗD@�oV�T&�2ѦT���Ь���r�em�H��m�릆����ձ�U�r��s;[����P���z���n�5U��Sӯ��y��1n�n�!o}�)�]n�Hu�B��t�`
պx�8���)c]�n���ȭ+��<��Ӭw3zem�ې[�x����X�u�˕W{��]��Ž��Y��'dt3z������:1Q��#�$S>;ۦ����9��m��U�GEi��cFٙfp\�,gPH���#3%�ܬV��+`WT�$���U��N�xVb�o*�T�,N��s �ޕu�5Nc!�w��f�9t�sje�f��֏�is�jRR�㣿fe�Լ�b����̂r�k��ÑԾ�Mu�,����a;�p85s`����i�e��Z�T���Y$��^��={�����f5�U��M�����`]M4�՝�R�VH�r.�9�mu�ir�2TT�5e�K;N�ir3X���dJKf��Y��M�\��fj���]��nk]�R��1j��F��e����6��5[i4�V�U�T�d�����5�aj�S�1�k����Y���Ke��t�j�f2�f�r��X�L�6E�U��%��cf�t��k��sV�r��vȻ���q��b�(�5�t��c4[R�̭�٘�ej�L��u��Z����죵B�ݙ�f���X��Z���(V�v7N����h�Bæ�)u5�K�Z��1��Y�J�-�8
�;0�j�d��duv4���l��D�*f:hpő735�j�R�٥Ӵu��̭��Vj�\6�Uc@e��iX֝wM�Õ�3���gk68�1�gN��P�Kcb�fl�KMĚ �(��u����� ���P��ds�v�<Aײ`�]4��6'�|�i2�B��a�ԉܞ^M��d�'k9�������0��
��]q,�w��q��]x�zB���s|�S�c� ^
��z(v�#&X���=\�k|�Wm���{t�E��"�'CdN͇�U��*h�cN���F�T���y��zsY�z�Lv~�����]c�b��|d(�)�;(>�N�e�gf��	P}[�s39q|a�]Mt�[�g�������Ok.�P_
�:��{��s���ۏ;je�TTef��*�����9��RҶ�0�^\�8�(m��>����u*՗^];Q�gX�����)7�d1P����N�������BR�����:�|t�{�HTǍe��]�>�֨[�Tȅ^�H�	����d�V�\�L�)�B)획[U<T,<
q�G\\�}�U�ָ"?�2` ��#��/����}�L�k�^�haQ�/2�b�r��|�l<Mwn��d��Ӥ��壢����>gEA�����oG���+���2oWy��ܪ�o�)ٰ�:{P`D���&��=yY�6�x^���=�(���Bx	�A]l�q	W>e�v�Iev�(a�t}��)߼1e�;T�Wp�����˗�h����c�}���*��^�����8̷��°58v>��5�ϖ�uYK:#����/ 3;��D/�r:����reԥ+NgVT�?}�����C"�)	}gF���X�"��p�� ��)}�GAt���J�NU�\����%.�<�D�B{���g�^ӘY�����N&��0�k��#�HЄu�}oې^�8����=��������;4�]�'�b'S�P!��t�f�p�*p���C�����Y�.0x1!�Mxk�%�_ر�	��Igz��B�I�#����m&���j�غ��J�ۻ�!����Ri��ח�NK��{�igF[��8��!��:����	���5�V��)�)b����E���o>U��|]
�}�xP�׏T��n[	���B�{�����i��c0�5:9�Wg�Y#�~Ci4!�(����Z�m�͎�tw=�F��up��vpd��q�S���fv,[z\uIc>�%ᄨn#�yC�{6d�9��N���u�^�"�f�S�c<y�Ӂ�ƪtǳ�V^��4wl�R���.+v�ofckl*$�	Ҡ'�Ҁg�@ߖ�f����'KK�P�(6a� Q�j���QԳ J;'Q�wR��WӤ�;����� ��X;��<���vP�P˺P�FHEs
y��^�J�MX�]�jã�M�в���͠�sB6-��k5��X䋶1e7G6ogN.|d�=��#a�0�1p'����ĭ@�:e�)Qt3Y����g��������:�tn�?��%�&x+�T̴H��0��ۣ�����t��U�Q�������įD��p֚�eц d��=��I�
�R��YVC(E([D%��1���o�q (�6t�"�^_k�*ת���6�Cg�EB�ÅmOa��T�z-G�-^Çk0�/G:�[��Of�R����\��O�<�p� T=�@TGK�M�D;�P���qV���e�l�Q��#=7�������Y�jU����ŋ�Y��8I�O�<ڍ�ڽn�,�y��i2\A�^��g�΍n��X�9���nu���cMs{���-���Knd��H�%�$���Q,�ظ��D�0�:��˺Ua�~t`�;=�1'�)[艧L��B���K��(F��aBŇG1Ȱ�N7y�c�3G�V�\�yd�[M�3Eq'å��Obb��k���+�w��7��R���=������M<O���v�=�6kùh4P�:,쩤����!�f�=�/'�ߊ~5*�`x]��j����B�O�%K�A#���BH��]�&���\�O��m��LW�m�{]�hcǶ��R�]ւ�r/P�����K-�EK�W���˲�p�M�>g��٩�'��չe�WT�-�8�.v�e>dw� In���okⳖ��VE�9����ꪪ��c��o�Tp���91l��X^Z�x������^׻%���goL�O�|���(����SX�%�i/��{U�/�tB����:��f�&�:c���th����L0PquպM5�TY<�J	�/M �%u{�te��%���LL�N���a2�����lO��3.\]�L~��٣{&LW
V]#�L��p�gp��S��W�ur�"^�G3\��d=m�Cy��s�L˔q���%d��s.�R��E��L6��J�i��T��[�VD�C���Z�YҚڐ��CxO@�xB�Dr2�c���ɦ�h57�M���-l�ں�a[��;���70=���s�"P�z�Q���D�����X2�{�t�n�
�z�%"��ŋ|�C��U7wf㖚a�L��Ftt�M�X�i�uf��'�%�|b���Ы�g��Լ/ֹїҙ�.ˣ:˳����nu'Yr󡔻7v*-�ۘ�MK�
������Q�pdiA�NDJ�ag��ci�w�,h�	4i����y��{ʟ�E[}����Rn��v.����3�f�E�+-ӄ��q��,� �H%��i�b�=���e���ъ�;�C������hW'>����nZ9x���K�B�y˔�\��{RIJ��V���I�*��a.�\������.]ޏ�o�lr��z.�Ju�\m�i���:<�v��*����*�^B�����45�SH�p�J�,���;�<T�E>�H]N�M(|P�x��U�k����ܼ��U������lа�	ĭ&��E٠�$ч�m�m�㍜1��;s���t�;_vq��a|��Z�m09�����g�_[xݻ��Y�!J�:��8֛����`���s�s¢����$��tEGs�����8�#��������¹����Ps��ܺ2z�81�3��m��٤E�'CdN͆�ȋQ���ܮ�vv�f�z���;=��=��7׫�n=E�gE6xU�߼]MLu	y)�q[H2����W~6�vV�G���ۨzb�1�k�bܰ��\`u�k]j��KJ�U�
���G�lk6��ָ]�haq<�T�����U-+b�0�)�Hb�P�6�3�]�I����=�'�/J{��h�u�3�!�x[d ���Nw�|'����B�^b��:E�*5_��#����;�,�t��`FY^7w�ur��ʶ�nZ��\��K
wU�a�؄@ T{8��i�s�H6��!UP�P����H!Dmem��h�-�(��P,�T˚X,w]s�Hmbmu)ǡ�L'Mi�x�� {��������c�t;jt+?zfx9$Bɕ��2��B�(�E��"<��c�8{f�j�:��r����Ē����#��9�(:�UA\�u��t�OgY���ȗSܧ0��aɖ��95i��O0-l��;n�GO@�[����K��,qR���*���t�Kp��n�ܫ���'���G�A��`��`�$,:�%qx���p��^	��3s�s��U�B.��e
�K�u����K��:G�u�]��gN��U�2g>#d8�'MGr�"��m��
�i�N&��0�k��g��(!g��;)�H�'t�-IU��p*�^�,:\�n��Mr�"j�P!�N��P��b�lJ�uӂD�^����$�nt��"��g.��W{xl�/��'S����B���p���Ȕs8½�\�ɬ|����.�^��t��k�O�.&�.��Q���`b�n�rN��ƒSq{���z�aUN����֝{s���zv��^�HЌ�ٿFl�P�򭗋��X���E�����Rp�_����Z��������.u��X�]kg��e6����}���%�	dH���g;�A�ɚol�L��Ԓ��^>[[{�muI���λ�Z�x��L`�O��*o�v�ڂR��������Kv�=�_GO
/�+#Lf�5::�Y1�F��R/:����>|�>��z��}�������.>b�GXp�O��^4�o�[aW�l��Pi����?"o�jʻ��fgg%�i/�LO�Lt�=
���Jwlg�:Zs��Ƭ�l{mV^�%$ڇ�Ǟs��ZQ�xJ.fXw�	�� �<�l�i���N����(j=;\�mu���G%]���0�L/�t��>^Lt����c�^�C�U�g�d�Qi�D�C��dM��]�E�4�\�=w0�͗���p]b�	d�D�O�Z:S\�	Kˬ�>\*&k���RI�'95�ս��Ϫy�y}O������R:���`y��.�Ŏ��U�]�u��h�_s���O�n���積[k���r/��<6�xW)�l��R@!��mLP3"��z&���N[��c��O�/�Ӣ�sf�ԫ;x�رn�)�g	#3V�=�9p�J.����D��t�!��"��xhCu�V��0\7"�T����o'|�ʳ�[gi�WB�niT���/��M7XV�pvZ�Sivt�!���:n�<�پ��U/��)+���G�Yw6���'V>1�t�Var�����Z�\�&�)��t Э�'v��V�������P�s6���t(��{��DI�-�-����Ur���6��E'Ip�E����݊��W��g�@V���c�P� �K�����ʲ����}�0꺨�a�%�PV�s�7*���Prs1��6�V�l�D�}��Z��@��P��I�\M���釐�{z\���LF�Y��PU,���(I�rs{���A�׷��"��d\�i7��@D��ċ�-;qW#6@C-�\^K|��S�y]����Q��q71h�"�`���7�i�����CS�EF<ۡF'[��N�a�6��4�R�~�AV�ٗp�9Q��S��	�Jx�㶺�unKC��AZ���N�\��'����	��ȸ�����SP�'OH2�݋Qv��;�B�1 ��..,�~�D�"众\\�])�/�K�b1ʼ�X:S3r�E�ٺ�N��c	Z��7n�d�xL`��Lƹ���Ԣx�����9/�������9�
�Ɔ:
}hg�	Z�ڐ��|P�7���LDt��Pl��~Y�UB�k
��je����u���1Xy=�v��iц�e�x�/��ȕg� ��&&ݩ�9�f:Z���GV�.2AOu,�:v���ȋŨ�jm�,�6oa��HVL��^']6�����z{�����]4���=���}_}UFM�[yө�����Py�}d1V�\�F7�`����r8\yu����W�ц�z�[�1���{�#���c������rT��{��������CL64��g�[������]dP﷉���NU���5�9���O��L!�s�X[ӱ
����ޗeъIOy^kֽTg/�feqj�*��0$"w�炩�6���l`��մ�߇1n	3Ԑz&7�1�]ݵ�k2���!������M<ഗ�.Z<�7�^P���V��� �c�5-�S�S��P�FQa8��_�m9�R�"��D����0�>5�H�O�W��^1,x�Y���Nɪ��g\Om3Bâ�T'��rFC
ɳ�Gd��{Q|����Vah�nwq���h���釢��R9D�^Z���go�����\��c9��2�޽.i�$�Ƌ~�"�@�׳������<����c|�Q�^��$�_b�s�]�������܎�ڹRb�yFVf�ڹGFN�Ⱥ������|�D��m�R�L���4gXx�Ž�a; ���c��|�gr*�E�.i�j����]%��3ʗ�ifb�����]��F5Y��𺓫��eN���>K���(k�X��b��A���!�Ew^���a�zL�z�2�!�dn�3���=�W�_W�r�<�K���_��Ǡt}�~S{�u�,�!FV��A��ͩ���rj�Y�
9������wi};ai�Ʃ���r��Yq�]�Ӟ��b��ԅ���8uVo$8�U��=�V��É��8UO�9��z�i[�o����םl��V(��D����u�P�.&x���<�7l�)ŋ�)�#���:�Z_��;/
j]TY�m�!�;��`���L�
I�2��Xml�k֗\����n	�tP7j{t@5,�3���{�6w���n��ɀ����3f+�R{:�puo�D����ܵ\M�'�,r���1�I~}$B��s���+�Os���.'�-a���YѲ�����(߶cRx�:�qJ�4c+zppV�_<�f�A�^��Ls��IZz�bPꋖKz�Ycm�,Z,��s��A﫻����w��gy�+H�WLmì���O,,bi��ߥ��;���ìM[Ϯ�K��w:�"�9N3 :�����p��uwa��4F��ݾ&ڮ3���V�RUرa��tVB
�oV���7X�F�n�*�ꜞ��2��i��/J�!�3U�d�u��c��T�N���`Ɉs��f�pzrCK��׊���& El�杬U`���N�&L�9����V+�L3U.}����Z�ϼ��0��2�[�Ҁ�Iٓe\�:v}l�}���Jl��1�p�
��k��N-�%g�,��td�r�tcJ�����vv��)R1od��_y$�4��%�-ӏ\琥�nfu�)��[Ru��C���K��e�P�ZW�v�&r��J���� ڭ5��m�$��e)��9�g�q#����q渪��T	�`�Krݍw����k�	�����k[�Kp�5B���aG�+�;.]�0;ٍ"r��[�NY��CY�3�Cv�ڍ��P9�<͗�f���"��^iN���Mv4$����܍m���k�����OY<��7[Ovos�%os�UN�8�J����k����>��gu���p��Q9�MC�v�Q�p ���;r���{֩�����.Y�w�|��[��=M��,��Mږ�%�d�V���W1�1 ��Laf.ޥ�����͆q1Ό���oT
��=/��.�U+gRZ����҇4�c'Ⱥ�/�$�R�V{a$��L]"�rݻd�gn��5
�6�h�X� {t�H��n;��sz�g`�\��V�Z3�ݗ�:`�Awj�uf����U�L���T�{�JpX����q8]컷���j�9C7`Ŋ�ZS�S����0e� {<��=qx����+Xux����z�Ӗ�����.)[7���YC��w��A�Ѱ�ַzNu�aQ�m8����Y����q�����գ&]��Gr��N'�j-�"v�JS��VÒ�YU��\�����he[�b��fQ�jz%���c�|��;�X7�1��h�ZA�Y�fﺁٓk9Z�.tC�M p��"[3jH^oI��;�9�.y8tv�8��:��&�](澺��Ax��1w;N�wv���s��tc\=-��mDWn�3E�����K>!�gI�y*�X��C8���dp���m�;�`V�Ko�'ԩi���s,9��(�ʙn��ʖ������an�s;Uz�nԬW�������w�Mdv�X�l%���h�耏BD�47Z�eȬ�7��.��OFe��p.\�T�06�v�Ƕ��)��,q[s��Nr��G��*��AGNw;�u���FwqE��U��༻�"��6� Ó�2-���d���?j˭���9�Y���!φP%�\T>v�M�=�wn�ʴ���F��'���9�*�uuIFNK��K )˺zP���y��s.�ptNԾ�r=ԇ* �EnB���!�WWa����+61ѭi�v&��k�f`�3M�ݬ�&�ʶ��K�j��w,[�*������6����p��-4�I�]k#Q�7V�:fci�Z̖q���L�9� +T��鍘em:V������̫�Va�����tf,6]�l�lk9���ّ��M9�dkN���g]M	�E�Fl��h��4�uGK34�6��S6�h�PI��[Ft��c���ܣ�i���1�Mkc��͆0�r���Yt͝��9[L]Rek1��f�t�1�f��b�f��	r��:��Lq�6��3�ͱ���ܭ`7L�18�͌�ʳ7*m5����	�v���Ν����I��Ԥ�*=y�����6=u9Mv��h7\�n�Y���5+��aB�w���	�}��F���m����PV���JN�]� }�8b��=���g9[*��1���sw��	5�X��'v�Zr�N@�]J�M`����d���'�F���{Vv�6�p��L�:�3��I��`�'P�D�YM���Q7����U�6x��G������e�@�!VdL br]�;�:���P��j�n��	)N� _*@�r�ZG9�7֫�ו8hj��j��pFIlÅ=Lu�ѳ�p����k�kas[4�C��������#Lfjtu�Ց��n*�F)����,=���F���Ӗ��B�����>��a�=SN5,F/S��!����5ca�mw�#�i����)J^��U P�8r,�B�&j%;�9XT��ݱ��6���Ьq�9�=�6���43��x�D��R���`��f������	��'����=���^�Б�Ӂ:u�8�����
��~�T--VT-�Fc'yD�dWe�u�'�u�.�71o����5��Yta��Y=����<Ԫ(\�X|��SY�*8��q��5�~|�����< Y���KƲcmY�2�f���y���6�k������{0νw��i{�wU����X�Ԩhwq]�#&z�,�c�-f��M*���:�R�:*�v%���٨FXc�먯*�l�ҊȾ����"=�cn/�=+�{]Q��6\~�s}b*C݊�1�n�� �>�J���%c�15,��]�5>�����\yK�5k���O��t�پ�y\.�N {f@�R@��ee�Xs�P�10���0�/�t�t�cV�u�BȀ�/�.��C�b��dS��Q��d�=w+w�Z�[d�Л$����p�<s�N'T0p��K35�rUۙ��Wn�\\�n������dV��NT�ȑ�w��ML��F�,�ؽ�D���i�N*s8FU��eM[Y7�� F@�E����2K

�R�nU!'
ãq�N��$�Z�ĝ��-��D��'�$@�'��@ʄ�&��Θx�{	eݪcؕ����g
�W|�l��o�aa�rq4��p�-jȿ�i7�ۺ��x�Yg��3Z~�i�r��ow���w�{����R,ej��1��"�`Z�o'��cG
����U��ݞS(;טc+s��\�^m
p�d���;T�������V��C�?�y�J���o��� �I:V����yÚi��~���Lp^�=k$��̽̿y�y��F���c�#t��%&7����F��-&��|o{��Ʒo���ɜx�m��Q�s#�g��\���ʗ���x�Tju��ں���kz�f�fmݔ��@��4�ǹ3�����}�m�~3V��������S��Tq["/,�����"Z���kG�벽�u�Y fc����i.�E(=��Oe��o�2`����F���砺��>)�7إ�m
7�tv���y۽J�!��q����|%j�fݿR̞5�V�G�R*�ѿPљ�3�z�[4��������%ƩC�"Y�n�C�Z��S��ԅnh�A�= 	u�h��^Ŏ41�tۨG�۵㞦MF)A�C�!����[���p��:��9r�h˳��}�9���<�#|Ӌ�!ǁCx��G�¯K��~��H�����q�?x���+�� �i��r�۱����+{u0))(���9��0�Ƽ����:3��9������l{�pfg��[ڡ��A;�O�$�+D�ѕJ�|b`%���O*kI����٫jǫ
̊�*�S�Y{��4���r���;�z�U�U��&�pZK\�y�o�]������n���4��������l�G��R�S���u��$��b^QC�p����8ƄY|��++)^G��o]xI��S���|��S4q��v�r��n*�lW+�L[��̧�L�V� ֊B%���ߨ���K�钥��*e�Wp�E��5Cz�ݺ
�ޛ���ni�]�1���cB��pBhj������T��6��>�S�$-h->��ꯪ��gz�iw������~O�-�7۶١J��	ĭ&��P]�"M��j�%�.���'{3��m�#��U�,eEڼg=�h�F��oyEA���e_[xݻ��9��$7��su݇�ĝۚ��C��]j�{6�T:Լ^F��p��*2���%�Ϟf���j�ى;�;j'�l`͚���=e��f���k�LO���{�O�;��h�Ɇg:�s15[�Ry�ZM:L�Ɲ�9<�L��X'��ī���<*ʦ��f�U��ܡFrw6���G珐'�8���cUL\cT�Nۖg���h>0iaV���e@󼽛�@ߦ��5��0!�:�������A�*�ŀ�Ňz���O?��xE�Z15S[�C;�3��F�I��=
���ȣp��Aŀ���O������M��&�{�.��{x��Ґp\�"���»#���i D�L�۩I���3���I־suyK���q�Ѹ(C]��\Mn�:�F�{��T>AČb�s��U'���pw�l��7��,zR5G4]KV���sJ��Ջ�"��%�������A��' t�n�
�8��K`j��=�t��G7��3�ryZ�����]wї�3�].E�V6��U�ɚ�j$:]�ka�O�j�D��cz[�R�09eCpZҾ˹�k�o�z���G�������[yy��;�nw���D*�۹�^��O`��Z��t�E��x��g�N�jQ^��=p�3�2�N�����Vn�0��1꺞� U���+:�y��O���{�D�y��$��ܔj;�{{ ����83̡ZE��6��X_��O9�<�ը��%!���zٜ�Mei���E�3D�V���\$_)�aC�xS�#!��7}�����hʵ�_���l�C��m/���o쭩k��b����o=����t�Q�kn����[���V՟]j�C�a�x{*L�9���*Ohi��hz(iB}k��d�-4j��Ӳ�ߟ�9g�
�?t��B>�0���(gl�#�Z#f����z��fG�l߻��K9BH_O5�����֫��{s���zv�.$�-Mu��v�����-):S��{�2�mj��X��kTE���+�mj��j7VZ�>��?�qV�i6uyOp�ݢaD����_,\c�Q�z��yK��`�9�W�0t:޵�O�w��F�@��R=�y���r�keg��x,*���e�.��g`�> 뭰��/}5��2���=��Ł�le��������Z'ur�45���ӆ)-gj�G��$�`̢�ﶲ�¨һk&�a�$����~�Dz.m�%Z֮��zeQw,i5�bb�a@�<�7�^Lԧv�A�KN@h���:0�����>��[���suc4�l��$�z?0�W��ϻ$���*̓�vJ�O%חi���/�	cQ����Ad'��OM~�<�:���-+�³�1uL^�9��EV+�E�$K�"mL>S�����P��lA,��^'���R��29_w|���Z:�q�0#C�ְ_lZĆ����)*eH�}w0"��&	Z^³���\�^©}��6;��.%K�j]1�a�p�B|�E÷O�C��w
p ��2�VƋ��z�UdNtj�K��O�#���c�I���O�/�Ό	1xn!�vv��-�ldf	R�jg{0t�[۱68I��$�'�e10���І���w
�X�/�ƂPޫ�+�`+���rʌz�Uo���.�ȍ�>^Z):K��,X��(&g2N��\��x۴1��#Wl���Khw"�8NF�O.��ڒX�a,�{�(E�YP�S�o����j�	7���-�v^�Y�E`�,���2xUo��^Ӂ!ى��ݖb2m���-�J��7wy�Ջ�7��&��׸}Kmץ��P�o�⃐�a۫�
�ۏr�kj}���ȣ����\L��d�(t���wtJ�J1�oMK�w�eL�C�r3���D9Թ��\�B���r�Hwy�jX��P�	(w��B{��k����/�n�Ղ�=y�=�׋�ӕ��yE�H-3:ݍ�7�dR֬�
�n9�>�{q"��N�P�p��%�ι1r+����������݈w+U@��3��x*o��c�C�e�)ְ�L�������ڕ�@��wч+P�RR\0�<�Lo�%����#�N�3 �Q1��3$
���ӽѨ]�=FM�c�{T�0=�q[�.X�sS��*� ���T���J�h�p�j���a2��s�Ue`B�XnNQe�E@讔��@��Yݺ�]j�j�ݥY/�ԄW���x����R�1��K2Q���c@���1������窕�f:ov`hq�x���(=�}d;s�Z�|%j����&dƞ�9ݼ���ʧ�fTb����H��WUB�U��b���!�����~v7��<ncݎ��q�:.�]��g$�L�ӓ�P(p#��=&z]v锊Ӿŋ|�GD;�b2��=}K�v���)�>�+�T����ՙQ���zD����>u�ˤHy�@��m���)��sS����R�`n���D�:oeB9�0+����ƸD:�մ�A�f�1��*ZY��G��F�G8��`D(]�{/�$���#�	���|9��n��IVA�����.����Mze�D�B3��aTדS3��c��o����*ӑƉ3�H&_��1B�\�.n&�=��I����_�KǖX&*�(q�'�y����V�.�=r�q�1�Xtv��"���ץq������r����u6_��×�5s��ާ�(�q���fu��,r2�	�� 0�8�UBFȘ}l�����Ɋ=���?Sv<-��ʼX*_�]�5�١~�����:k�٠���ekw1���K�sI4�N��DY�%��}��i>+�0�S~�@:�:�-v�[8ӹ_j��4;���@hp�ȱ�cDQ݈�͜��/fX|ު�.u��xlA6���ɪ>;�|��}�N�=鏄}\�~3r��]F�Ea�}�B�f�t6C��4�	YhT��i��m[�r)�U�Τ��Ɲ�4�i�:t_�mt���*�����Ƨ��tZ[�.3[[A@q�);(>���50�Ʃ����av;܍/ϩ=�Z�a��J9Hyô&w:N���:�;�3{U�u&T�Z��܍�����m�rR�b�-a�9�S�����E=�O���D��D�k�w���hJ���6�T��:@Ř���y(Yη0��X9�v����q�����o����av1�NB�ƒo��&�w��_���oӡ�_;�:��RҶ"�0�^\��59�DeU߭{j��m�]��C䱞���O��Q�Pd�Y�Q�[d!P���Ny�|�u����/�ౣ=R��X�z%GH�1%�ҚB���h.�w��kd�Qiu�Xg^�&��iS���N3�n��x!����r��RB�f�Q��9�Ғ����}�^X��<t�I[����s���������= ��=��(uJ�
��;�w*�67+����f�[��KQ��N����U���lh��G�A�P����`�9V����H�x�5	�Ժ:F<�JjN��>��GXR���P�"��p�,/����Yt�,s������(nιM�iw�pu<���	[��k��{+��t?X��m�/w�[�>����SY۷�ÈS���#�Ԕ5��9c�#�������T�/�Z��x�]�X�CukU�z'�~Ԭ�\��_�τ���gר
�P��k��T�,u������� �/�1���Ǌh��i�8�������j�;��YQ�˛�|`�ͩ1s���wP�c#o{1��[|UG]�q�;sݴZ)C�Ĳ�L�B�n�/ri�s�;�TC�>|��;3Fc��f6M��uv�U�sy�s0d�������l�e:ӹՕ9~e���=속	2�_�ظ0�\Y�	\l>����/���a�<+q���/՞�d�'<�B�:�ͧ<l�ȼIO54�w�z�����b��t@sMAs�����₉����k�q�X���n3f��u��qbE���Y�j7Ny����dpȆ�������=� ˋ���Hʖ�.!)48���/�3���.1�|��9񞩴��x������t�IL�o'vV�Ի6�8��Սș�=s(i5n&+�(g�f�W�%:�7ǝ-2-1��A�W<�������p�%W;�;IF�+����G�z� p��}؏�_����҈�#�\j��v��au-8�J�6p5�5�=��<����-"�f����]�ݩ��[�ڢl�j�:��쉸s�ž�Ӎi�Wц+Ĳz�]ə|[�*tV�g�f���I���=����7��F �6b�G�'�EK݊�1�NU��]J�xm1�iu��w�MQ�N"bc�D]u.z^�Lj�9��O�ȷn�Ǖ�Ѱ=x�c3�f?>̝�F+�=�1�
�8��V�P}��	�K��j�Q�P'L���S��ƻ�H�˷�G�+��'1!��QS�]�0.Iu*�ZY�9�!M�.���X�ݲUl���HX=Ɋ��`�ۉf���\���o�1r�[�n�uc�ZȺ`�ڗ�nn�y��7��:�T�qt�$���ݽZ�&t�8u�B�v�gȝ�����]�����E��֌L�Bæ��}�[C>5�FP�!�:�q�����U��)�;[�=C��Y;����<�p��u�����q�r�N;ЯN�6�,��bb����g1�̈S�e2ٹ�4`eKa���B�W+�c[d���^���8D1)�e�G�o��պ�C�D3���u<�:�-9��W�ܴ]���:[я�H�w�J�z�3�����k��٩4���a&���>�3h>+�Y������8����pO+-N�40hɪWkrY���W4l�%����D��5�����e^����:�q ۙq}���vq"�s��e���3��w��e��#�=�3ڶ���K�LFnA�'ؘ���ŋ�Xb˵�XL�J5Y�jY�M�g��'|z�����+�)���o5,.�߬��W`kX���1���ie>����n��;��Y�nyr����$�kv,��%!Ҽ=y��\Р�h@��&����Ў�|9{���L�p5X��6n���w��S%��-��n���|%phq�c�h�dԭ�$Us3ZUۓ�sM�bS�9Cks�B���������QyR���7�NY	K�֬]9j��ݜygB�J��
1��Hf#�-��8��;/9�o`blYy�i
�4����U��vi�x3����r��pXۤx>�@�Se��'l.��9��O9H2�å�V-�6���񁽧v�k���_R�I���J�Y�\+�v䦮�x7�h�Q�71b]��ul�A��q	�j���-��a��b���yR��"����F:Z6
�c�[S������D����Pn��k�T��û� ��/����<�� Z��:�/z3��U2��n��P�`X�L�{r��X�ujž��f��|鬩-�#��8���x^M�4�*"�u����ʶX����q�~ݨ���R�D�AF�s����6�e�u01��ݺ���B.Q��L�=u�V���;�n*]�%�}�η����הGIޥas�:��`�i��д^R���w�23�7Ifخn��㛵Ӭ�u��F��[mS�Y�O�A�*A��  Ū�lx��x��&DY��w�s�s��R//^P;�P���J�ڢ"E]�Fب��y�������L�
�NE�۔��x�rɁUE���}��P^.��LV��8��n«�=��};OgV�'/p�XS;�6���6�fL�1ԍPDՌ�(
��J��q��i�M	��S�4cF�*H����1��c8vn9�m1l��aS�Y�6�U,���[6v��(�"(������0�1�3U���h�H͊�5��f�N�*mW�����p�T1Q�q��T�a�B��Db�AEV1�H��1��������c<xq�F*n5k�����K��m1��ٛf�`�8x����fqɠ���f�j�bji�8*�� �"�0�R��p�m*��a�nº+��6guX�cclf�.%���&�	����lʷq��<t��M4�l�;�;���|����00�����աڻ�c�[�S@�|�J8�+�f��%f�`#F	�G�ʈ�s!IN��QI��\��s�7*���RKl�'$0!���ao��t�J�5l\4,�b��r���^���0WLc��[�Wj����d���GI%µB�b���Zq1��^\�15�%RF���Zo��ƗH���a��YŹʒy�:�Ĺ��ᬱc�^8��;�}��]���V�_u�UJ�92dY���EqƉ��/-��
,�����ZX����Ž�x�ΪC3�C�6��)8� �r'sQ<�4�{)����V'L���M�9q��Zp��l�a�*�X�w��#V�d_�´�rh�=b��%0��H�lLݭ�'zE[�{�Y�hUq̘-?P{v!ܭUX�2��cV�D�c�C�V%ؒ��
�v�{,1��|� ���0���xa3��=K����AYc�h���dՖeo��a��4Q�������Ǧ˞
�eV�|�+��u9���x�8<	f�;�9ݣ�m�Rg�����ho�t��0�Zs��p���A�7'(��\��r/�SNO �'����&yց��)f��@�@�zVe�NG([��;1�f�Z*�&ȥ2�@ޛ�b�J�g-|�q��urE������A��e-�Qťŷ�v���T�}�{#��ȏ�0�Vޭ��5�y��<�z1�ogvM}JI��R���\C�b+Х�������>�^P��jf\�덌(�P�u�5���V]�}f&����B�J&���!���-�hb�ֆC�+T��!'4c���ެ��9vV+�|���!�!#�J�:�WQ�P{���*�+�n�7��3�]y	�jo��_�Ih�w�l���̊��J"�8W��I�R��)�@�,U�W"�EԮ��4�\���[ݲ�U`���w��zi�3S��%�D�B:+�¨1�&��,-��󹗀�d^Y�LK���4ޗ���E��:ȨV�����Ig���c�& Iu��f�[ڪ,�Z���ynPp�zs��XSrrC�b*�T;G*I��Bx��S��v�jX"���3��J�ֺH�6���}��eYc��D�#�Xci�P�-NP���^���l���`(v�����Ƚ��O�1��	��lпE@�N%i7� t^�F��ScKk{t���M��#�j+�'��u���ੇ���m0��k�7J3���t�ѡ�v((����^�M��Me�K��;��*�|�+|�u�x�����Y��L˳D�6��|U'C*6y�;rc�h�'K������̲3]�b�s:l�W@�R��0�O����oi�r%���L��:tȗ�"�iϵ6Ǿ�7n�f�� ����\�8��o��9��{ު�,N�!skz�a�1;�/EE5�<��Sm['�t�,`Q�:�j��H��L��Z�=�(��-�*�zUbǯ]���M�fQ��,:�H�	���Ɲn��x�9�E��B�2���eV��gX�!�W[�79����h����L��%;���B��S]4����#C�3XFN�y@�S�1�W�&�1�T��X�V8W��θe1za��*|XF��KJطL.`eЭ�4\�-d8W��=/�^Kf��peK���Pd��Q�[d!H�,瑜窶�1�a���ϲKڹk�Fys����ve�='��X�I<�L�ꉕ�Є��|�ptw�~�B��jğv����ųo��B-���{w(�ARB�C� �����:R�yo�{�I#�-��(��zmw+�p�pU�|�&��N��£P�H���`g��z G�0Pb2)���s��Փ�'wyvI<���`�R�a�U\��pp�x��^C�Vl<���4)o��b'xE����O�i�Du�+`��^�&��y��M��]ء��|�`��^a�p�}Bًi��%�~�Ϟa^6��������7ź��N �xw�%��B�ۘ�1*+�Ks{9�>�}�\�R�φ𚬿�5��LRR>r=mkO����fWD�v�vI�܃(K�� ��01�{~q�aK��!�+H�WLk��J��B��+k2�$����N�^���\UC�Y�P�N��u�E�f9������5��Y[~���%/7��������TD#�`��|�������^׭���	5�X�5��8"o��չF�����Ԇv.!:E3tX�)ʜ/#��!��P{{xl�"�<���1��wY��o$�lL�B�P��:Ns�ƫ=r!8�6}>��ty}.R�D}���<+ky��#��ٮ"Ό���j1S EBwKA�s��mj��yS���9�Ec���ڻ!����ƒ���4#$�7�4]m`W���Y�c0�5:{�#nU�tQ;�հkٗK{�ǔ����m�!��k���Fz�//�߄�+8!2��cT�n.bq��X'�-[���4M�=�l��Pi���9����`�� )�J�1�Ԯy�ԯ�k��^��k��Iwyp�������f�QB}ڋ9��Ė�J~`=> 1���7��3��N�23�i�����mB�+0�S�	��HU[4�,�Y D����A��Y2�$^Q[��uZ�2�C�A&
�l�ǿ7��[��h�0��n;�*]�7�8��.�i뜻�S�y[��j`��l5�8�M�Ԩ�<�&MH��ʔ�FK�:�u��i�>���E:�����OM@�����ǈZ1QT�U�s��թ�d�#x�Y}�C�Z}�6�)���l�CZj�F���Oio�h�{*�2^=h�g^��\.J����xl�B.�m���b?t�9������{��B�[ͬp�L�m�WSY����.ʸ���랒��z^�.�����z�r.�xoW�[�y̹ն��Ļ�@�a�T�M�!�B���|hM|�i���vmyq�0XyF����C��$M�j�����p�а��X�3��<��$�'<D;a������:a�������s�٠�պ��skF�Ć>�ʬOT>.n%�nd�d�������$`G}�H���(ߓD�����o�N� �,0�̨���9i<���L����r��i�;�����Y��e��(�2K��D�@N�)��	�@�rRyW�*p���GIq��;��%=����;83�*��W���Qw,h5��^ZՑ~
�y�>�lv�:ϥ��8��u� �[x�u|�/VP/q�n���*��K���t��#�����mqᩗ�`�C~冕��:� ��,����x����#F]��36Ij�M��F���+Eݔ�"�d[|KK
W�E����尚ŭu�i�_��f�/���4�RR�ۨ9b����|�V�h�7��/$U�o����x{qуGq�!�<֊c���]õH?_�o��� ��9��+/��5:����Ry��Qn �Y4���mup��*4ƒ�.pm��:z-P]-��.`^9�wC�]�⼺����� ��~�up��:zq�L�9m��{z."���^ˮ��� ����[s\�~�B��=W˼M��b)K뇁K{1���V��3n���@��p�=�$z'ʒW�� ����Ph�PW/���)�k��{~��e��L�.!����~�}�+������R�a�UҐ����Hd��>��[�r/��cx����k'��[�wU���)��BY�)9(��P�^0c�L,���<JEaP;�q-�s�~Fzv�ħ�{�}��P�q!�S�<멁P��MD���`�����;��=��0>�؜�ge���ڞg8��vb���f��EB�On`RrG�yh旆�(K���r�	ϐ0�vnnއ-�'U13<�n8V4B(n��7U�S|Xy�m��ݺ����Un)��݅�FAg-1�x��˼�E|��\�	��Y��7P�'�L���M>���}��5�L�&�����r[��ǒxN�Qk�\`qr��\P[ӑ+)��Srn�ע��)׸D���IJ=���V���T�e[ݒ]iK�(}����3j�1Q�,u�SH���t��b��#"K�f��o�2�$��ا
'����lU0�{/i�ӂ+}��	��~�Xʠ(O�T�^��^�>�c���s�K����f��+�eł��x�u�'�x*��������?9մ	Zb���W��x�9i�^d�CM�4g��+���r���X��1/n,g�t�'&,���y�\\u�m# �c� U���~�n��F�E�د�#�@o�������.�{2>#իBDN͇��e�-����6��[��l���{0m��B]i�����;򄨛@F���h�2:��d�V��T/b�Zb��S];���#Fl�2pu�g]��]�"u��먨 *X�V g]8҂7�Ѓ�UO�S��~{ژ��t��.gR�<ic�Q�I�!��^�O�C��ު�� .� ɘ�Ȣ��C�|X����z�fHw���Zd���5[��\��ϛ���80��j�����@z-�뻞n��%�^��T��c������+�rН�S�}9>�1�5ڹr�e)bQ-�؊���`���k�νk�廸Rԏ`]��Ƣ�I!�u��b�\Ɨ3���)����>ο.�.̱�zN���-�!Z�����X�˰���k�j˥f�����L�/���'�j:���Q��AC�������UAD��V.z� �/{qU��Դ�a�r{rs� �-�ț��S�v
�z]��T��UK����뭡�we�s��,�W(F*U��U���lhv�[yJ��y=�0 �=:�_^�����y�t�D�����عD�|N��u�삫GXR���2�i��ܳ<۬c�!=��0l���xv@��p6�?Su�]�\�8^7�f9���
�2.���撔oVA��P��l��ʺ:a�}u�[
��1�����ow�UR�İį��(�
��r��KJ�@�JB;	�6�,��������:%�}�˴��P+��=Yy�-�G䨓Z�T��
���s��q�k˹�p.��ig���\��r��z�s�P&y�=����o; �*`����w���)��dXX+ ڒ�u���KV��!�����D�J
�
�b�wf�G�\�{{-�0!�Ӆ��F�;u�M�u�ּ���#AmpQ��)���Rǡt��ĳ���K�0ڻv�25�w��d$N�JXoF=���u������ù�-s�`�'�0>Y�w�����9F�zt!~�\}��o���qbE���F��7k���g�C-q���XIgA����F�Y���H�6\ƚ�B:��@��������64&V�;&��j������B�wSH{���Pi�ɝ��"e�&�n&&�a@�<�*|�������U��l�;j�~-SӁ�Ƭ�vǶ�e�\L�ٜ�'��S�'���N�	g{�/�$�^�{���k�oI�H�0�9Xz	CQ����Af��@�;%���[�SĖ��}�����闤�Θxn!l��->ț�s����ޜ�Zjra�;��N���U�=h�Bܥ���męA�T�,U��Im���	����aQ�>ʓ��V��W)��i�O��5��<�O1ˢ먡s��ڗLj�5��	�y�zo6����K�3��~�]�7�/	>+�)Ҩ���bz�|lGӸw�S� ��CȬ���	�C�.�L�m��������^	�Ŗ���ꈽ�:I<+Q��O\��N(p�qPo�+Lø�|���z*u�m��ws1jSx�v60u��j����r{V~����2G��d��%7 �C��wU���,P"n��^�z�T*M����T��Y=��S��\\%\�X���^����'>�V�2q���ŵe�_I�'	�3o���3:l�
2;�c���ȣ�p�C���X�s�$�s�9��u�u�Ҽ�;@}Z��S-�jtBD�G&��TI���:�������4�]�C&Ic��wi��<���[S{���g��,K*Y�3<�����S)8� �r'sQ8vk�:ʒס��D�[$�}}A���H\�sr*��Q�����,h;���ZՑp��hCm���jGV�\�.y�lz�}��%9�^'�<.�'<i�����P0��0%x+��2{&5�����w�MN�W��j��Eç���ʿ^F�/�%�	O/1�P�guO��6����"h���P�}6I|"(�x��KgF�9Ѣ�ƒ�.pm����
�G��/R�7|�U��c+��l��D��g��.��=8�&V���_L� c�;1gݓތ܏�՜�ڶ�7y����"F�)l���b}P�)of2	Z�!�cvUܣ�[YeI�)�k�{� �G���L�WT�p�R��Xx��t�0 �S�C"	Z��u��YfĊ (Tx�h���T�X�*1�t�u��&��)pW��j^�ǣ5��_El+�HV�&�F�x1�]D�D��k�����_jᲕ�Ϥ��|Ôla�=��N+]�;{m�{��A��{�zp���԰�T��F� �co�P^M4S���v�T��9�;�����Red�H̡�ʚԼ�qNak =�f��
�����|�H����*Σ.�����xʏ:�7���/)���f*\�5�*9ד@�K���o@kq���7�
�գ@��S{9�lԖ�/tpx��c����|����z [�Kβ����SY��a6%r�3��&���|��b�ځQ��W�|�+�oB�vI�l��!�]�]�����X�T�� �P�'6�JT&ti����gI���Q4C�c��p�Wz�d�N�ņ��leee+���s��U��ʻd,]�&����O	(�=k{��}֩x��v�薆���dA�v�!H��|�uݤ[�d8r5U&�3Wع�6�UbT��{����^g�*�$�$�!����Gr�t��h;��袼V�����[ہu X�N�W�>��Ic���r�u�<��X*a�M���jj���'���"5��oP�^eO$J�y���w�Rs� _�=+���K�8q�k��s�7�����\t�����vJ��9쬑V�h�-a�"��a>�ng5�髥mW6���!�Ҵ���s��ݥv��#G�����Ɉ�J�Vʽ�z�F��9#�tϱ��ջ�onS�1,x��Q}R�XZ5�d��%�ᗦ5�����V�_Ez9�]'lb���tx�cANB,�<��T�r/
=M�EA��K�;�P�]IWt��:�Fkk2�'5��BM�H���"w��a�ϓ��2�
H9�w�/t��o����Ȍ	V�M;hn�+t:��Ol��V�n\��z��״��Arr���a��&R�m�J�����d5k�-��ʨ���݉�����r�q_ZRQۜ��搐�F��]ݝAK��2���r���z�޻3�.i����av�p�qV�ʵ�d�_M�&P��ڒś�kcyG��6�4���Y���U�V���rL�
j���A\��g�7�6��q�7w[3`�rv�֓�̷��;�E��"�1�y/6�R��K��]�7{@�#I1]���3�f������k�,,ST��EY�j����)�U',��	D��xԉl���B�Ǫ�1������i+|_R�r���k��S9pՕ�}�[�r�H4I��ݬھ�&j�J�=$�x��)��\M�������R���#Q��{
-�y0PrXt��B��X���af;�OJ5gkz��n���в�J!%.�&ʚp���HD`?J�ަ]�#p_�5g3��Bv*�jy~��dGG;�.�)2Z��ǖ�k�I&捧��{#����cDQ?5����u�1����{���L�SKD��R44RSIM	AE�1%4�SMPSc a�"�Z����� ������"L� ��j�(��%%�,cE3DF'T�DQLEU���SAE,14D�Q�0b�M44�M��1�b��ff��(��5t%�j������ ��,�A���TA3MTL�fpK5DETU���fs6��aW1��V$���P�-!�$�"�ڬ8fpf0�Xؚ��*��
)�&��#3�j3�A4IDTPc`f5i��8�1����ycf��1���`�a�k��&�3����׿
�N�C�Ùϵ��u��j}�4�]�5K�P�o����i`�@�v�B|_%v����*Y�Я#͋+&�����9;wn���Z4t���x�I+���.�Y.ns��~���ve��O�MgV�8�T]���X��r8�Α*z�Q@�<P�C�B��E��vQ���9�w�ܦJ�㹗ҷ�`ߧo;/��x�y��:s�J��}=u*����N�B,.6 ս;5�W��?a���g�Af�u<6��9�!�1B��Θ���s��'����W�P#��`����5o[�N�~�e]̭���{�U�	T���n刯9��hD����X_�S�=��d��!�Kl��T�a�(o���9��w⬱Ќ���Y�[���.�p��@F�	�M�aK�(H+�Q�X���X�x���v1T�_�H�]@BR[�ڒQ�[���'�cYC��Y��jh�1c(eEۼgFI��1�������9}��=qPZ]j�i�v��םr!ًb�;P�3E��a��3�,n򇔗,��j�kkD�����&/ak�N3��,X����=[]F�E�UG��dց���m����ܷ|�³M��c(D��F�� ��M7���5�! Tφ���ӝC����3����MSv��j��D���˴gyFZ.�A��t\ux:���S���o3�e��z 7���2(3#���gZ���'�=d��(�s޼3�/�f:Л�x�Q����<�,�,w<,��U��n�#P��/w�v���9�C잓C	I�5�Z�<ݞe/{���ܺ�21�36�͔ɺ�A�Jwc1���/��v"ܰ�]��;��67�x�ުz���`jѫ�FɁ�4��a��:���("pp}2���S���n��q���'v�_�{٨������b�
��L�q&c�T��ꂃ&�"��-���x��\���&kj�]�{wE�)��}�~}h!q/1~='��X�I<�TȎ%p5;���ɳ:��n��O	S��!�v��#o��BY��S�D$(�P�e�
#$�������dō΃�߳+��AS�'�z�,��uܧp�aQ�9����ʹ|��+��;��d	-�p��qsĺ����U,=�����N�ȇ��ø0��[ۆ��\���x�\�s4*�+V�5YY�*"��_I�Q�����*�u�R���PxB��1���h>k׶q+�����}�>#�3��W^���HN�3M�8w|�!�[��k�i�v�DA�3sn �#������#�t�>�+����B�6W-	��XⲯLj�>jk	��r���f���ժ>�^��4�� �����L�W�k�vA�Fzt(V�gn�wh��	�'Gx(�r�g*,N�^We���2�P󡍼�nMM=�zGCǎ���g�%�*"ʳ�u�]�{F=b1�ǰ���]�ǀ�cd/w�.@I�"k�ځi�Gb�����,Z������:Ʈy�v�)r5������e�����D��⠧0�l'8����.�=r!���xX���j��9����[��g'l���4�����v�T��J�w��x�Z�+L��[3c��&��J�t���i��Ěf�d��ʹ`aj�:�l�3ܨ���7hx�E4 ;��-z�O4��4��ρ�B�Z�~Ci��\��Fz�X���VpOWaj�s��v�=̬l���~����{��z\t�3藆=F'�(g�e�͠�[�@]��Y�Y�ꗺK��z2*Zp4X՞�l{n!VK�r%a�-������P��^ͪ�mᜌ�ok� ���[%��_w��!�5���j	�{�J2��z�~��q��g^���s�_��Aߦ[$b0��-�E��~s�ž�Ӎi�V]cD8]���@�ޖ�5 ̈���;(!�Dl����B�C*��ǲ��{kn��\}����J��Xo=��s�ʋ�r�2�Xp%�u�d��KY�V�	KV������IE��U���O���m�]�p�z���A�����Q���;p #��ϐ��Jp��B �~�"pg_�;GY�g*b�p���F'5���Lӛ�Ty�+#�\�D�k�{�uY���`�a�/K���U뮢����Lj�9�����Ads��Ү�����f{�\�cyL] 1P�Q�H`B�ba1�e�vњ�?L�������oGLFUʉ��^t8���_evx�W�G�l��"��p�'���52�t���6m���|k�j�=��wT�-�T�[�]�����܊9�C�p�"��9ʒk���n\��,	]e�--���۽��F84us�f��Oqa�a�(������˸y�v��739����d�ޤ�m�|��{7�I�g�y��]��^�Bm	c҉S��%�����#�jk.�?W	��l�z�͜b�P�L�u��|0U�ţxr������KZ�/�f'S)�2�M�d�ʧ�^�H����}�%="b�x]��NxӘ�p�g�:����/�x�.��'��Wn�d	�F��R&�m!ݾ�4ph𑱏6�U���R%�	u<���B��n���G��5{�� ��f�D2�aC&R���لj�2Nj��u�\��J�e6gs��]� �;���_O
cڋ��A��Aڜ}k@d�J<�v��7i��4�����Ώ��E�o�39�j_z�WBr�yN���&���2olv��r�B.��;�K��ҙD�<t�q�]\6��`u���:��C)r�FG7Ժ�v���}#�|�����<I_^_;蘙:zs��ei�n�r���XV� �뱉y�C�fck-q*��P&�S$^)l�{LEyK뇑K{1��J�9�a�؅��Ƴ�����ڞ08��)=Q&cTˁ�mJ'a�C�!ۘ��AO�
QB�oI���譫��z'K�[RÚ08�]H�F\�vD��j1Jq���ΦB�.p�'x���^�Hn�)���>ˑ����I�DP(p�0c���aT��1l�����[(`�y�=6���0��q�\��#-�GQO�o��D'%S,r&��x*Ќ�md�'w[�&9��Y4�P[Ҥ��u����1A�tvdT+On`W��%c�2��+�[5�s;ZBtUL�N2`1S��(=��YL,���Ó�:�P���J�v�\%XX|�r���%��L5�x�g�ɖ;roJ i�RCEYc�DN%i��{�V�h^�\��[�n�B�1�Us�[���ԱN��;�eӌ*t�Hd��־3XS����suأ�#�OU��]���gK�s[z+�����z��oHpp�\y޴�ǝ��Y�l��W@)o7'
��*�j��M=��p1�9�^��n�ՉX��^�Kl�G����\��/
&��@7��۬�������3�h-��K�@mAvh1~S&�>#�vJ��}e��0�S���<����1q�*(�퉂ֻp.����;E{^uȟY���8��o�8�G����y�y����ty:��Vk������Z���:K0=��5mu��xV�<4@�T�NCq�W�8�4�E�O{5�^N�ȝ�y��[M۾���j�¡Q��߮�Y����ϟ���HT#*�	OS�ћs�L-P���g0z!6��E���&�(��$<���/�sY.O|�T��C���zc�L(buӁ�PD��ߕS��q����ʖ��V嵙���лea�n�]��` P͙�.�&c�TJ���(2lr(��f8�N�d��刧4�<���r8�O��Z\K�L'��X�I<�*dG'��'M��獷��>[��p#x���,]t.g�|!>�Q���Q�$(��3^�@svl٬��86j�P���{�+�鷀)|�Y�}=ԅk�M�`���������
���(�/��dA%!���K�Έ��=Q�֩�0��5��K�.P�U�k	����Snrj�p����:zu�������F4p��g�XMt�_D�k^�������N�{��G��y�@�瓈��Tu[�;�|ti��
��9V��ed
֟�_��;��~�`	W�����\�]�c ��;�T��/�+�����>9�=Iԩ���T�/t�`ŵ�Jbx��ىC�.Y,T_I�]ν���
]�����4E9pS�_�3A��|2k�	���)o��_����u�]�\�8^����e�{���
oY�9�t8K�� �8�c\�Pc!N�"��HC]N�C�2��g,���p8��]���{ĩƟ\y"S�����:E3tX�9R��L��u�4.����順#�-�dMy�ɴH8%�74 ��N�����8�H�6Rw7��,�ס��m '������a�蜞��v�". ���y��S E't��9�"�N!}O!h�����P~�(��}��ەe�C؏.��F]{��mV���G��"�u���Z���3���}�V�lz����M�8����c,�mߐ�_4!�(g��,\bQz�\Z:PT��ݒ����ݩh#}Ž�.���z9Y�}n�Kl���' ��QXV�x�yk������P���N������bf,+IGV�[�|vM�w�ˎ�orV�)%��#��kZ�]�"�obz�����է;ZV�Xʂ���l��H��U%*��l8�h�7�j����c0߻^�[z\RXϥ%ᄹ�T����'�\����o$Ʈxv�sa����)�1��-8,j�vǶ�e��ڋ9>J��I����PuҸf�^�s5�@q��`
�����Y��a�@N����P�rgC��PY�x��-��OKΞ�")o!�A�[�-�-ɝT�{閉���B�O�&���1p�OoN5��9���7�e�v�o]�c��,��^%i��I�
�U.\�!�"�m�mp��V�f��0��0�y���$x+��qY����GL��
 u�P��xo�]1�\���1"p+ם�7,��ܛ���:Cw���yep�S�P��"P.�6D;ʅ��A��Z�2�K|�$�/��ժ�2놇�Y�7.�ۺb�D:Ȧ.�H�O��WS�u����1��<����-o�Q4QɌ3:\�w���&�|�C�+���O���]o�e��9����Pi���Jn{ܖ
^�.tX�΢ӊ��M{�(s*d����C�X*-�綍.hp��wo(O
��E%�9-&���9V��7�x@���L�D�#�����HY�C3K�7ܜ�w^Eo����&ĹXt��e�8w���ҝ�r�ܰ��y%'`\7�m;�ًzP��	؎�T�FT�X�,�κ���e����I���x���ġ���*_fyk�����0���J �H���Tv�P��I]�tZk���]Y��b�L`�ًG�|X�W�z�:�9��E�
�{��y������q`��c<�9�kXO��ڪ�3�-?POR�;E{����k�����v�{�GF���R'J�Ǝ��X�n�q��%�	s�£�� ��~�|��rݝP<#��*9��U�S(���Lt��j��`x�oG��d�m�]����x�$'A� ?WJD^N� ����)�\��!�L�9m�U��b).� �{uaU�f���!
ˉ*��J���@�)�7�M��b}P���c!�F�KE���O�X3%�r[�û�,̾��Cc
u�B�����*Un)a��!�u�{#`.�y����VN��WKW��)�e�}^ͱ~��z�9�Ur���R���je�g�{#8��b����Y�9N�x�<����Nt�_O]J(��(q�
���~#�e�ۡ�ug��m�+���=A�ג�e3����t�S�>�/͌�DpV�K��9�.��H��N�pu-��*��Ag�vn�����A�m���:��Y[o�<v����ؒ�0��&ob
;�P^���᷏�ʶ��v�+��Zw�+�sS�o�'�ۜ��=]�8s����q�>3}t��;��7	�/Ϯ�'%Q2�#&�X��镐��w�t_lB9\�,vl��xmg8�.�P�w.�ì��~���H�}9T�]9.9C�Ԕ�.%�S,v��jx�P{Ӟ������Ó�"�@�0�d�y�T���cb�#�$�0x�G�ˊ�:�&�����f*!�E��4�^��k�$n+����9`����ë�I�ļ����/����Z�	C�o�soHln�*�.��I���\iA)�va��**BQ+I��00y�<8��{kP�M�j3�����ʏǮP��y���ڝ5)C�g J�*'N3�7��yDC�t����j�J��Y���|���*w��vF��p-t����&�9�x��ph}}T1dȞh�VlU��D�w���4�'�;<T��٦o�ȸ���P��-���ƫt�s�NfІ⫏TX�b��8���6-�&��A��"��4j�ht��l߫er��������xY���랜k��*/hK��mu*Buݤ�l�Y��	��N��{�4��ޱ�vvs&-I�Lh���s�����]�J!Bnry;���1�쩳zr図�.��%����(feqօ�J�:��0Kڍ�X)͆�y��qL�YSD�@snu�0�cBsv�Af����Wq��T�p�K���R��1��w��4��*&&n�B��Mq�TX��ܭwgN2�)v����3J�2b�5��r�$��L��SܙG�U�|o�M�8 �&wX���>Ԩ��c�t���x���k/Om�&���	��Mp�:�n�ꢼ�T����:���AN���D����\�A�d���S�ud�\7��q �kh����d�M6���Mb�����d=ݧ�B���TT���b�F��c�������E� ��Mɴ�̨�0tUJ�:H�V��]���Ջ�굊��S�V�G/{�6�k���ؤ	��QG/�Z֣ա��}9n_gMe�J>������u��_�VCA8�ۻ-O�����If)���k;1"����k3K1��*m���� ���e���sD�E�İ��ާ���wg�r:���;#��'�Whs�`U�]�*#�gI+hGY���#������{��D�E�΋�5H���x�zc���R�8�u�`�Jda�C�q��Ϊ�����������(��JQ�����\��/�����f����%�UMWܩtZnBr<7�f����cz,�-��p�ѻ�b�	�����kI�G�\\EA���Pڄ���l�U�3H�-������^�@�s��rma�`�2�KZ��V"�{ �8����Vo`�R��^�_9a�Hv)��3%MB�dðԭR>����vNe��MF]d��+�l̈g%/c��y%0��P��턬�4z]G6K�:�'sڗ�uܣ���J��/����l���\�kAR��&ˠ�I/*�9��Զ���*h)?��:+���(����W7�q��_r�)8"���Q�y�s���*�ƨˡ*�(j�3�$��>����P�,XD���J���+��̌*�,5��.C4_���r���7$�Ŋ�-o۹g�뙉P[]���ͮ�1�Ǧm̉�W1gO#�r��:����"�|m�Y�e�5E�SV◘�4>����8v[�K���u�[i.���_l_)�F7oz�ہ�쬮ZvwCel*���úgs���;�0w�u�it�]�����6<�{��X��ܿ�&U	�8+F&�OT�B�F��;������+e�����n�V�O(4��i#K�9_>Z �N=�[�f��9B�	�/�+Vd*��Y�k�ν�^ݬ	���@�,�G�Y�5�ǹ-�^�YS |6�[Mګ��hp<D@�=�x���R̥-f�}�SB"��N��Ͽ�_��w��ٰ��X�V1�6�SWM���a��
�q�V�M��ɬl;9�U�@g���0b�3'���8b ����$�D�sh:����ov����I��6�ls9�m��.�gR�b���j�����`�"b���#�0��RQD�Q,U�T�3Db�3U5UM�T�4��E��#�f��`k�� ���"���bk�ʰV�3�;8�f%�����1��	���)�`�MUDQ3,6,IQ0D��,M1U2b��QT%1�;9��'Ff0369�s6�3qR��lv;q�)k3f1�,4Q%AT�AUܫ7�&x�)v\Wrg(�TNsy���An�K�b�u+��m>I�h񵛱#W$[°,��j=���$��*5�OsK$���;::wg�3*3�y�vk�K�mf�ǕF�����	W�G�N��2>�`GĪ��0\�&�*e���J������m�avC��"��(m�gh��1�*TO�d�v&����K��e����l��dp�_r�=��N�@�2���<@c��L�Y��ٜ��A���e��1�Kՙ�cn����5���"�g��>����F�U(�RB�C�]l�Ow%%�oe-i
�����fc��AS�'!)W��J��
�C�"ǹ��WӽIU�ݶ��ـ��zAs�(=���xE���Kj����6#��|.g:�7D�=��2q�O$�ZT+��
�R�%R;g"���/��w���<�j*喜����yDI�2���׬9�f���%Y���c������p~�'Ll�5+���W1��je~��مe��Cq46.�^uwZ�4ED_]26�u�n�M���*Z�1��I�NE?l��{�����,Ey:��9v-:EC7E���@�
Bư���Ӯ��|���Zq��M/X�Y�����X�Ww|ɵs�,���e���WtɅ`�(4:�*� ��R�u�!�����E�vB��ظu���T��ꝕ6#E�����Ӫg>�a^�tRy[�O65��Sq7;��ո���6�^r{ =��A��
�r�|�i�O.�Yrb��s��95:�f�����9���U��Ӓ���٦lh��y��S Bu+l.�yS.RE\�>y��ǎ�dXX�u���X�D�,TG�e^&6�k�~5S=t�r��ж�P�����-%����6�w�������֚��Mg��ME��
!���ܩp�;��G=�.�_Z�xV��ÑB��1��Z����6Y��6hǀ��VT4;4"�N�fTfkYS
��OO���Wha�KN�
�1쾬��Go�8)��k`�s���.�}4%�&+g�x4��(7��t��C�(j0��ޕ0Q̪��}���;����IZ%Q<d'&Xw�u
��F#
��-�DZ}�l��1p�Jޜ4�̈�0b�vѵ<�,���lJ�8)_��uy@4v"�lk���˃�.'c#�ӲhC�{[r�{�fMgW;�C��4?3�ج����0���7��j�/���)�/��n.{H50��!bq�䤥��N�~�d^�|�Pu5�fO�&��Ag�Jp��Y��S3v�|�a&�Vb?�g)��ӝ.��������Rgawk��v��쾫���K;{�%,i�������֊/��g�mj���������!7�ͧ�kG�G-됩˳}+��b�{����$�7�ckD��LH��S���V�N��=�����1Vu�vv�[.dS���52�t�g��s�ʱ8E��ֺ �BbF�\�w :��p��ȴ��YŹʒk%9�P#m�)��S� ��
N�ᎋ5��	�b.��xuy.���H�T��v�$hx_�I�ʒf�f���8�<'���K�FJK�/��,:5���^�w�4@%��6L���3'ة���y��|siT��B��:�g�∪cY�F�f���>��}��q��du���X�����#���Y����E����i��z��ŭ=�z��˻�z���j��B�a�t��{Hv0h�ӢF+���2��/}�x��Z��u&bO2.�C��-��N�0l�c2��Q�[t�q�[\-�+ц0���j�N�7f�wfbjh*/ҥV�&�S"�t0D��W�O*��I���&{5:4�\�W���7[����� �D������.F]q�կ���������by�����嘅Ɵ��6���l�Y���c�D���*�^�NT*gc�J���꣚�c�nW"�ɡ�Not����]�Y#�}XI�DZC�Z�A�n�52�o ͮ�y1+�/^�t��|�t�g.v��p+�f-�[(G�	�)oU0���rA�[�h����8��0�j��{_�f\�덌+�(�43���K���b��=�D�]x�sG��ge͛y[�si��P@v�A��+T�[P��<h2tW?��/7Xua!^�	�Tv�i���һP�|�*=mQ���ġ���p��j)9(��%��(Fb���a~���`��� #���X����:��VǓ��7�����BrQ�u**��BN��s7RH��`p���0�k��c�gz�C�)�s�D<�:�;E	�NB)v;Ի���?OI��{$q%fXꋘLT�8*4���"VTt',gx����7`u��\�shvbRqOn�6�����+i���v@��T�VN�,@Ñ���8��N�\�p�<�ǹSV�I�0��%i�^i"<\�������u�^L%�-�7>��SO,�O�
Nx�4�/��
��Iĭ7�r׋�A�I�}�;&�F�Z�Ώnv��SΖD�(/��.�qK6���ͼ�P�������3z�R�@A�f�n�݃iZ��x+Hh���%Z7��԰t�n��yK��p���"Ú�@�ojY��Z�1�KO�T�>�y[)�"q��:�G	���Y��r�����	�+��˲eaђa�uTY�*{���i��`h�k�"�;1a�t�z����{�
}�]q,�V����6_�<z=q��**:D�s��8�}�t&F�-��5˚U�%��V��986���(�a���a��˅��4~^�l�`ɕ����ƞ�zo�jޞv�q�87mj,m��/��B���SB^/x�x�z.��?nCl����i#��ty��>ʌ�y�v|`�ͣ��<�*5�(��ϨKţ�t���4�ix�y��C��ӥ�DsҖ���βȍ����3�Y8FD��;���&��ft�����wd�*|X�����S�.̱�zO��<8v`�e4_9��=:�8���u��d�7ϪD&w���<=Ql�juR�B&���v7g������3q%jd"c��<�q$��[�Kܭ ��S��[uA�Vl���~�ݻDxF���j��|c�p�;��|C+�)��"\|�c�S�9�<�[����s���	���7�Y�`�A1ӈJ][	��h�Cx��
�vs�C���dS���*�
�>�0�^s\Ml��[��_#��IxJr�mu�qt�ꕜ^�����uM{�G	2�s�n�ˋ��\�1{Z�N[5C���ｋ΄b����Х�p�H휊��8�O���?�|��Wĉt[U���q��'���tk��l��E��j卸u�"c���'�UGi��%8jj����研w����m�Y�Ꞝn&��0�l:��/��C+!t��^�0٠\wk#�˞��h�b�c.W[cw�UR�~!	�	��#�����,Z���u߬�mb��o�[羓�|E����o^0�,\w:$�jqPk��(����9S�ǷW�S"�n�-��ݩ��8z�����fȜ�g�a�c����S GO����3Yʰ�h.����~OntиPsHgd(ׄ\����1��A�U�s�Z����\���v�"��n�Ntu��=o���_��Se�0��]engU�G�mK2�����%�]\;�]2�[t�fE*��r��q�Ƭ�_ze�&�!_#�Y�;�վ���
u�Ծ��z��n�<�i��:c�q՗�����R�;��������C�#!(�ס��u��\�'D�S���,#k*+��1E��Y�C�W�pӧ��jK��e���9k������[C��S�ʱ6�Ż��~{��aL�i���	�j� M7�!�zm-�d���;��.W���۹���
��'C� et��	ޅ���a����>����7lWA�6���#�.�F�A�8��͸d�t�E�D��S����Cޚ��/<��>Y�LP���^��.��s�0� l'p��3��*]/����C`MTf��D�_)u��y}1��!þo4l3	��R9�T��� ���W[G�ĹxY��f�ء���n/9-�]H[N�z��r-ۧ���p��S��{���H"!�Q&���'@���T�d��\GG<t�ۗLj�.�h��/�r���<�,\C��a�&3��%"�gPU�ᡔ:��v����/���a�[Yh<}��3�L�,{֎<����X�x����{X79��W�[��vD��u�0:>Z)?���X�����b�d3\Xa\T�ZrdvZ%�rK�r<���bO�Rw�艦������]/-O
�\<%<˫�d�Q*D4F��i�|�6EZY1v@p�% *9HI�\_=��AVK</S8S��'MW�}N�<ދϠ���}��M��vie; �~�w��Rt�q����W�ok�W��'IF��,�̔�t�}���j��W�[�y�	�vN,�X.C�^Y�ؾ�t��`�^�Ip!Mo�G�9s��D8��.��v���Z�jKvqf\�����"A{����\\@xV�|��^,�Y��a�0Yyw��٧.��b���v9�):<��n��>���g�/��m����Xwב�5��u*a	�����k�h�Br�^�tâ�C=���d�&ۖ7OE���p`jKf�.b��w}��jUN�B�:�债�Ε=^��`� ��ص:�w:L�3	��R�B���5>��ٺ�v^�꬙0@���gg��qmU�ً�R�6����/��L�!�<�ո�2�=7{0ڗ�X�7:�d���
��ę�s*���Mb�h��G#�n����niY�a
}hdC�+T�[P��!���z !a"�uT�}ܗ�|O7{�������I��d�����$��O��=9�<f�������駇��PUq��nN�*^�!��f�g��;��Qo�ȿ;�������m(_����O�e�&o{M��&�u�a�s��^OGT�v���.ˣ
[�D�5�zI���S+u��gn�[��]H{;ܷC��/���*����[�(�"��1jd�\c;b;X>X����s�vs2�۔j�^t��#�������B��'���VE�,19E!��˔n���·)�
j��Y���q�kסcO���7zqw+s{�n��Kr�p �{ W,u\�
���4���"%eGXN��9��0�{[���zcC��x�]mP�T��sDӬഗK��4�7-`��f��T}��N� g����z���;_��Z@a��UB�8EEF��5'��҇�z�X�fw.�o���8�(;��z�����١J��N%i��r�vhxJ�5�Z��t�d�t�a�4v�hc�Iz����|��a0�V��W{򞭣Q�ہ~gy�65�Qً*+���9��"Ω{�=U���K������;E��Ӣ*;�TT,t�L�:O0��>��J�4`�|�?{�h����A:�T�6;ѿLO�Y��)��;��j�4�"�g�>Q-_���;ޅ-l{�8:�
�z=�6ʡ�`�&��^����-���A���znq̝�3�{��)۴-�P���T�Nۘ�o.0��u'��]j��X7B+�y�~�sp���L�uӭQ�v���
�*�`s���O�i[n�]��p�����靡�*]t�!y���~�=@�Z�{):��p���=�8��]
�$ۣ���������3Y[��{�w#"8��Ŕ�e242��pҠ�p��^�x��K��H�]����W��e��R�U���Z��co��o��S���c���6ԗ���5�
Ҟ�b�z�ր��,�QpzP��z'׷	�_��!�t�*D����W[��=ܰt$�	��D*��������x���a3��C�<=Ol�h�򝣂FP9s���Ē����\��r$ ժ��&c��G��_��\U���c@9P������>l��*���̫5L@^�&K������|�G\S+�D���&k�O�+��d�M�c̼#�y�|^	�:]��:4)m%#�r*Z=��zlM%�eWvv���}��͛E>��J������Zn�p�,,< D��7�
�mn�c�#{�{�fzOA��O���ûӢG)�adT��FGy�1�j���8h�F�v'�
�����ޘv9�ݶw=���\VA�-��ODr�"��P.��b�:E3tX/��P�t5z����m�^����rJ}w����,_s�N�a:�3�@��� �6��f�9!l{�H�� 0�*��U_9*�p4�z��~#K>߷�ɯ %�d�����Ť�]��N�����3�ޭ8Smq1Q��8W�j���D�9,�t
^�+ck.Y�$*�E�]��WD�X�͡O�M��j��s�);���Vuc��^rO:�����+J�/��l	�)f={kg�3t�#��$��g;@�6
����S�1�s�׎è�s�ϕu�tm>���8�
sh�������P����W*��
��D׹r�\Ta�Ȝ�ʛ�e��ǝ@y�L\�t��84+Ŧ�̆�2lNn��YS2d��.�#-�Ҍ�g��G�jи�FI'o3����F�LGo0o[�N�
�B^����$�˛�g-�J�}u9N�A�.c:���Voe�7�h��w{�p�w�B��,�Ek��9J���u1cvՃ��y/L9s�e\.(d�);Kj���j���fm��U����Jؖ��� �ء|3sV�l���%��{/6�F�Uf�W�V7Q`ؒW����5�APьY���l���P1G�R��ג&:�nR�d<bb���Rݚ�������e�M�d�Z�!3z��G,���2g�P�X�<�y����ڙ]����Q��"�N��K�����͘^	Q���\A��֍n�CX�e\�v�A��W���ƣ"�C��;~R�R�UiF�ZV	=x����|��-�)6c+�'R��^tܣ�6�:;:�"���2��W����h��;��wk^ĺ�N�W>��/f@�K"9Vڕ���oV����nRuXEl�;���o)W�}�u��+2��$�q=}�UGYN�K�;v�sù��Y�R�-2d�d���EWh{*`�����{�-VQ['kVj��ѓ//.� À����B��D��<|tD z8`�PJ����e���{7z�s�v$R!pώڷ1��u��H;0eڸ�'v�Ud���q�2
u���8�-��ïa�c8�r�7��|�y�7P���aoGMVO������k��f+�WTF�u�ʕ��Z��g�d�X/�%β�eq��<\m�$�wQ�n]���S}�I�zT�Y�-b!s�0��6^u[=h�͓���a��	N�Jh��̻���Q2p�qX���
����k(�[�*������%�rW[Yy��bz#p7�Yv��i��yOJŢ��2Z�9
ySV��(���\�)ZZ���Kߛُ������ �Or�{"A��ʈ!�L��.a]A�iG�WV3�8�_s�m��_'J��:���c%].�+��;G(ʑܾ�8�1Ծ]x�[6pe�ĸu����f�O�P�%�t��f�h����B��X��*���#O��ݴ�Vq.S���t�4^=�M	�U/p���y\�ߔZЦ�S�����RRw:g	)QQg2gMv�o�̙���h�_<��p�Ċ���9�Jb^{�uՐ�G.[�J��-����t!�w��
��^��_w��>�Y��v���1]��f6����fg*1��E5TUbq12�TLFWNf�bUլa�a�3�3*櫳2�h���.�N�FH�`q�l%�U��Wi�퉦1��-hj�c,������4XZ��Ηf뫛�cq�I��U�FV��Ls*�6f�uA»������gnWXq��9�FWM��`�3��s�+�̧X����*�f�6��h�̚��s4��ek�$r6sU�k���6��-ʎ%���,�gfWFi6K8Z����m,�cW\�Q:s5Ns�3scB殕flfs����M��p���J�l��ޛB�'��v��
��S�ѓ�A9�y�9i�-���|;��Q�7�&
qu�)�܊��z�$~=�M5���^���=��B��Q��eY-�١��)�I�=��3|���UL�J��� \cڍҙ���g�_��R1M�K�ҀhB;)x�W�^_y�����Ӏ���Ж->c������T(?yx��Xwjy�l���p+�i��E�uZ1%5�i:���A\u{��O+�3ǝ-9�¸�L{/�Yx9b}�v'�u�Kti�����QrXu�t�WK TY��7e���L8N^��P�h�;�jc<}/�x�z7�V��������u||��;��9(G[6����y��"���,1�����NW����3�P��i l	'p��::��B���P�쎱���Q�����A�D�w���~�w�$�=ج����0��V/�X�_5�����HG���8��ͫ���Z9anz�MN�w�>W"ݺxoW�8!���hD�2 W[�Iָ�̙�A�9\�'�]�S{=�b:U1�`��������Ҿ�>�f����|듉�u�8��j�lr�M��e��wf5/�����+� �=���5���L6(r����i�6�쿰Z*�4�l%C ˭�X��o6����♜�+�+f��YMY�M���%V��$��T;�}�����;�����h1�=2~-S�d�C�/c����(��X�&�C>��:rj\�J�p�:��m�8�{����Z>�*WI��1��>�"43�E'�\0!co�qA>������P
��S�$8�]��kw�Y@G@vl}�Yw!�$��PV�%
�4��Vo�7�K�XٜZ
�<�v�/� ����,t�T��'�D�����ڜ0�D�%�/w�L`�1H��.h��$$���7��Kv�U�u��C�Sj�y3�P�����1�^�0�����c�跻Z��j�EfR�!��ߦTb0���&����7kE]{��b~E�ɯ:DT���JA�B�e��âW�9P��U�S(��j��;kk��e5����_ q�{��F��u����r��'��"U� ?��1��ry{k�*�8q�?w�(���kl�L�y۱H|Y�c>����	��b��K�b8u��3�XEWZ�f��|�n�#�&�Z��;n�d�P�Uc�:"���&�2��Y��~����n�PVb<���֨��h����kxn)���hI�Tή�1�.f��Z`����&Υx��_��γ\+��sF<)�����mi��j	�e��s�����jī����B"��;�a�S:�Ln�X�%cw���B��tGT'Q����Z�Y�=5ǯ\o�U\DB��n�$�N{C}��4�zf���j1�r!���E�DSs�0P׷R4(]f�����7ںI��u�i���G�{���
���`q�73�^��,(���\;��էq�n�HN���wf�[����M,�P�'3O�TxRzs��zӭJ��r#�t;S��y.�P�3=�uNk�i�m���y���Ȩw	m�
�rB&�\���t	�[T΁��� ��u�7H@����4�~e�O����P�:���
~R�?���4��Z��S~�`�����z.�4幯�3���I����YC�F58��\��\)�*+`������T�
�'c%��#7w$촏�z�HfF*�s��G��:���"M}#�K2�����{qs��M�hW�L+�SE7쫷U����'n�΀����!؋���5ϒTcE�9z��ٳ4c+0�6v��k�DW��TW�:D�':�b�9懶bD�|��]�u�����ꋨ���լ�p�*1.���-�2J��t7��࿺��]��7Ռ�6��;)�5-��]�Sѭ�1���Z�6_t\9*�s;'j�pu,��/3Ge)i�1v��d�O4mw2���Lf��a��R/���$�GO�L�7�Y�@'V*^1�qOf��a��[X��2V�wz�����bV+�bC��pz�
ߣكl�>��B,�SF��ht��l��ċ{.�Ps���q�<��WrE��M��z/I��*3�5N�yA���譪�y𮫩��Nm_	�s.35�����JߧB�a��΢��}KJ�t��w�DW�7��U텻��0�-����';Éq11�4u�7�d1H�,YN���}{i�_��6�XR�Ě�%jIIE��2IAo�dGTL��u�x�E��a3�ߟ	���{)��ׇy�QY���NBYU:\$(�P�nJ�j��.�:
�����t{��T7<����Eԥ]�҇*̞��t_#!�T��<NPu�գ�R��x{*-�]�w�B�n5RU���J�4c+zpB��E��Vn�0��>���̞÷���X.;t��P*�u��w������gg��aK��B��,fì��;�tH�g��٨2hj���%m(�!��"���%���٫wTz���xN�t�g
]��^b��s���ok'Fa�p|��T���v�bvB�h�ȯ�U�]0K����\�=[�p��uK�%���mS�0Tӷ[���M�Z�N�U�w,,u��Y!���:��59��C�Oמ��0���.Z�*m�XS����uv�8h�1cs|almCnz���IdvU^���|1�������T�_��%s�x�Zt���0�[��I����n�ĉ�r�T8d7*���Rd�׋<`���Q�T�v�`lg<�u��^�d@9�C�9�k�����.�U��^\D���C;f����.�
3[ǈ�t�+5�<� /ܩ "����s��q�}�qI�N
i�80\�F�#$�]K^���t�X��w%�Hd8��}~$�Bo���{Pݬz���0"ǻz�LK9�ؿ!��{�h�,�=/����������b�%��3k����Q�	�%z-�b6T��;	�p��5a�	=Y�i(�^��IF���Pc+��=U�F���y�Ӑ,-�vǷ��S��Y�����J�w�JM'��R��t��X��H����/��'OK��+n�9���ή[���,oqJ��D�=��<�@*������Bc�V�v�#B�<�j.7q�Zz�C΍D&��NZ�f7�V��sVbUx0�3�35��Y3�K��dL�1�k%����O�Y+���X+%�+ge�����d��-�7s�7[�-���=B
�ɒ��p�N�f��+~́C���x�#�&��OQ��[�+zs�i�Wц*	�zx�Ү$�qR�YD��q���ݑh��赩i\P�z莨���E·�4k %K݊�{��F�a����,t+X��e�ӲF;�zo�9ڟ\���\�7
]0�Z�=V�\�N]�����!���hD�*+�jy&�N|s���5��0����)tƭ.�h�MTf�w.��C�bźȦ�*9�RN�F��SM-�@q$�5��j B6�B��;5��9+�Ȁ��r��i*՝�Cz�"��ߗ�\R.n'��'��$i/�墑<2�5��	�g3�8����ִ���u�]ە5m���H�9���CH�I,Z���xmmR1f��p,:-m	|�u����ͦ���X��
K
Q(O��z��=��C�va�(���\����c9	E�,�lj��]����ezT5kV;+	�tc����T5
Ft���kgU䦮�'zy�O�/��<_�X�چ��z�Z�x���X��a��+o��$Y����=s�B4戋���L���	tDo.ʔ�s��V{Q�JL؈
`���a�{Y9�w�a_!i�B�h���� �J���^����nKN�E�������sXg!Wfv�,�V�A�վ��&0����7r��\���o1w��K{�嚊�r[w|v����84B��ʋF������Q5mS�!�۬{1�x6�e6�+�<9�E�Li=W::�gA�,/Z�da��//�w�1�;t���VTd�����S����!�>�ˊ�������T�;*�Kd�-�������b���޺uH��쀥���|߷�!����ơЪ�h��Y��@�[4+�NS*�g'����6��u	�pb�ֆ>�N5���D�@�xB{.�KF�zq��ܺ�M�_�R&�1Ks���b�����#o���{���9Uä+�k<�<��5ֵ��<C�P�Fp��c�]v�L�^���,U�W"��W�����1��Gs���XY�wn���۩�IIDP,r/�b���b!C}����z"�>�t���(C)�ӭ�"�2wk^��f(7r��-��o��'$"j%�`���M,&ì<=�� WW`U�2�����K��F��C%��;�"���Z{rL=�\K�yh旆�'�wCOmT�ZyI��y�*unl!d�oi l������Ce#K�*���K������a�m/o�.Z��h�d�]��n���Zq4�����E���
���M;��sOs���=��][b_��z�:`<j;{Y��Jݴ1�:s<���W}�y-0q��g���M#�<�MiXckΪ�1jp���B{�\]�����a���;���p���/�����̌U!���E�*��<.m�t�f��2lÅ�F=.�s'�55C�\��9E�^���s�v�V�$���:y�=Xa�w�:GR@_�R��ko������*CP_��!��>�v�|��m���������(��Q��_]��y��5wj�!�,���A�^��1�b
���H^�e��g�2'f��u�AI��b�-e�M�L�Ǫ���s��#�t\>��42�yP��/J}V`,O_d����t{�Mu��Gk�ՄOOr���n�i��j���m�z*�~�,/�=�;)���,�U�X��o.�W:��<:}��c ��i�zVۦd;�#C@��##���%i��C��3��)z�ƑS�1#x�j�"���!�E�b�S��<�O��;a��8N�=��nwo9.�) �ӎ&X�o�3��L�����hG2��烆��9f��pUU�����iJWDh�	�F��(K��:L��VBwsʺ���:(�V+�mz�mf�΍�~;}e`RmЈ"�(YX�e+e�Ҝ0�%S�Ӽ���7�[�P����!{�Ǥ�P�sf�����d�I��ēy�u�����Fz��J�/^G՛
�����ڜ�W�p!�P�f�&Cާwp���F1v9�B�����T=�!�}t3�ʞ��G=���>s�Naa�F�I�j�qD�
*x;����.g�-g�cU7qL�߮�罪.Ď#��A|�x��r���������HXt���Vu;!^���t^��8��o�, ����A��k�mK��B����b��XC�g9<�\����p镎l���^		�Y��PrN��<4tASl�ȀꞜn&�Ź�6�]��㫇3�hB�u�Z�[g�ciX=nne��Y�4��a-��p��h�}C�F��`��ŉ7郕�ޚ�����[D�Uj�T8d7������,�V�%���DfC�N�xKj'�O�i�W������-]�NY�#� d8�}.*�~V��O�j��xPWA�L[䙅02�T�ݍSj��۱X|-��CXyhB������؂�s�:Q���V�XN�<��t�F:��nE��ŀ,j֬�ǵ��~kVE	^��)Ϲ�<μXׅ:/^�8Y���T*��c��K���*l�OX�Q�oI���YI�Cо��u��M�fz��T��PG9O$:���i�t����;°���pB	�jW�o� �3\ZAd�9��D�]�<ӵ٬�Q!�W]�{&ྵˁ[��zk#��,�Φ�p��v�]j�uj�xumVWq�N��L�jۦ#r)VӐ�W =m8�ͨ�}�N�Ԯ���D�fD�0�=J��]A�7��|����ޓ��+
��ao�K�&��U˺1YwK�34}��w,J�E�����/.�0���g�@��Lؗ�@X��p��b6��ۂ��������,j8:2>tx�'I�2��:"�zS��^�E{�å���Y/leb�t]"D��!`0�L_��[Ӎi�V]b��zA;��+GJ���
ev������c��'�}��2�h�^���E·�4k $_��=�*�p����>����!��s�
�^�����RP<U���u�C��T��n��<�p�S�4p�����z:�%r^�g��$��� P��5��0����\��9у�L^�]�+����X}���Gg'��di[��q���� O9<MD��|��P���ѡ�9+���0M�h�:���Na��}Kr������.7
�)��'�#I�^Z)?�ᎋ6Lefs>#���xzC�f��R���-/7 ��T�P��ʧ��9�Jrέ�%��,K*
��U�7�D�������ь��ެ��\�N�|����+N+]�9v3m���.�TJ�VˋX�s,�oH�eoM ��C���^fu�DZ�A
!D�@�v��,�����r�A8Bx�����8i�|�g��]n,m�wm�@�#��[J��aZ�f��rt���n�� 6'|�*������t��1B�f ��9��s.B�e�y�U��[1�5-k2X��4{�
C���źD���aY���cf1L���P76Wck-�*Bt�����c�x�n�׻��Ǻ��ݣ�v��s��Q3��t�
i�A*�	��"�E/�m21���k��̈́�~Gd��:Z���s�l��c�PW���G���d|��w�g:}k5�W �Ɲ�֣Lz�bg^�ի8ۮ��;�%LF�
�2Q'\��nuX0����L�IP���@8[�&�5���8��C�"���X���}��S�O޾�^z%��dX����-^�Z�3�h�Zw� �j���\N�պ��l�b��̪
W7����������Q��Py%�Y���;v�]$c�e�[\{��4��t�t�6-Acz����[��{n8z�V�a��Sb<v�q���y����b�+Q��W��VZ/3���'���/�rR�;UڛP�o�%`�,��m3Q�}B=���,e�yo��``���>���U��]n����0:4�i�{����f�c�ֶ1�f��v�彋��'ŕ�D�:�Ι)*`�Y�զ[F��@v�i�G_.*U|Ugq�E��#;
Yz#��4O� XZ����{�����S������d�v��R���b��c�!'/Pmud؆�Ŕ��c��"���c�\k��HJ�y��$l �˷ۥ�JfR�}���$�#��&F-]�L�gI��� P��N5r�Yn���v�[ n��dyB�8o�x��7C�Gzޡ�%�h;��sT��������s�����i8��}��c�+�kT�q����kMr���[����u2'���!�}��\�5�`y�afqDm���̕��	F�ù�!�@δ��<�ҥ��T��*�i�{W�f�?�o��T�닰[���i�n��W��`�z�w@�9�\�|��,��nizKf�n���OoM�mH+Fi̏O.�sx-��]%�XF1��;�x��	�Gy��wWYB�w\�d�K��M�r��)n[걋^���!�!dg��H靘y����V�
�Y�vR�� M+s{ɷ;/����ӈ]�{Q%5,Շ�X�5V�epl�+]�:�<�sm7VJ����ţ2]m���'m@əԋ�$��j���$Ik:r5��6
i�7��
5[�WL
��0R;����|	Rk��%�`�e>�SY�a���ҹ�fgS���b��*���䣼Wӹ��U���^=��+��a����s�4�cv�ZYŃ�i��]�s	3c�eJӌ'A1�h��T1���a5Pj�V�K��pΨj����`�K�kub2t�:�V6Btrɱ���Y)bd�L��*�,έl��������Z̭;�R��s����3�i��u�mi��5e9�.k-.NZV�'(J��+MN�l���Ȫ�N8�%���j4��%N�L�ʷ2&��ƒ�5j�]dUj��J���5��3'*�Vڮ���5j�Tqr��,i��R,�]V�Vik�-lGV�䌚L�6���&��K��f��f֙F�i�`1��\�i�3Ef�-iE����,�Z�U������kK�ծ�J���ڳ�����e6Ziu%���5��e�jִ�|����׿�cr9mnG�yS"�y��Y��N���X�6Y�L�6�;���hޤ*�wս�����Ga���,t��Z'�q+����P E��'/Mì����'�WQ�-yh��Jg��,f�y��=�\b(�I�/��Ӧ�Rx��Ә�@�N% *#����U��v�5Y�������_�V6X��-��o`��2�/���oS�EB֬����ۺϗ�5�jy�k�fl��t��C�mo��I
�Ns�Z}A�؇r��ڍf�88�D��ᤱcVV�����s��h���6|=�)���m�����Լ�� B�)��ljÀ~��(}��_������}�\.��1쾳��1Li�p�������9���8< �V�qu�Wve�2�MD�s��-����0�Zs��p�W��$h���'(��U��P2+���*�Qs�刔{\��� y����5���)����4!�Υ�(Ş=��k8f��]t���;ו��=ف����5�R�7l���;�>���C[L<��CxO@�qլ�+b�뵴�E #Qu�P�%WQ�X{���*��َE>�>������]�1u[i3��pg���V�X+/bu���x����&�E̼����6!��or$��b�b�1�בż��5��w��N�����{Q�ݣ�4�Zz��坔]��:wq��L{8�8U���*���Q�/�F�ՠ�SZ��0Eϫmo=Y]�x2�� � ��q1�.��L�^��,(���\;��or	S�cn�^c�5[��dO�2�]u0%�F}b���b!C}����z"�>�����v X���r����9���f(*=GSЇ��]�����B�|c/ǐv	��I�f���\����o^��Au˕��d����n刨sqP�ʒcc��K�壜�����46�C�fo��(z�3��B�*��86��"�mC��#dLdj�lV�|��*�c���7�"�j�}�W�6脀��K��lи��^N%i΀�.�,�Ol.���b+:1Uril�1O�Gd�zK�*����,�k6�� �S�hl�Q~�0�k)���ZZ��b�/'�嬓�۷~��6Х~52�{����*ӈU�NIp:N���'c"DM0���G����1��*�ߡ�����B"��p>��B��/�dgfdV�u(跉���ݾ���Sު���H�z���Csȡ|p=��4.����a����x����'�o|{x�pnn��*���O(���ږN��bzY���jpP�;��m������M��ob*Q�3�a]�z�zUdW[�3�n[�g�����:����Lat�9p֞M���ή���xu�{bΈ�kg��͜�Ɵf:I������Jwc2!���/�t�}��U��K?E�`z+3��8��ss1kh\i~�p"yO@�Ζ�D�A�.�y�`MK����Yd`���}SB�|�d�M!HQ;%93APbƢɨ�<�6��b�|X�)�ӏ�|�I׹<���g��=R����h�:rU%��e$�zSHV���A�|z�=�r�������m�1xB	���5i��7��
��fPs�͎�%[;�M������G����S� S�ٹ�+��c��}$GS۹���7�Oq1(:�T].V;��W��WX!٥���>J������e���pP����yJ��<���jʝy ���HI{�s1¶W;�7��1�P�S�o�׳�
��65�+M_�Sp�,,< Fƈ������P�7�SSe�*��P��!,W�I�]θp¦م��=9��ؿ9�4ѓ1�Q��
��*V�y����S���#h禸�WfяX�e����b���/�A�Ϋ�1�[i�wn���=��gȒ���q�|����*$��Ҭ�B���A�G��/�bV�)��$UH!�V�N�Y���?n<U���-yw��6����3o/9���n�Ud���ueA���6p ��j��r�	���[簞?`Qɜ�Y�^{v�`:=f��50
��kG��d�׋<`�[�d����;���Vs��'��5�eJ��I�F���E��p��t��jT���a9.�X��o���<���|�ia�Ӏ��`�L	Ԭ�V�뉴��M�4�80&㒴5gfs��+*�κZ��/�2N�١�\V�},�k����7k'�O?M�~��a.n�=��ӻ���Z[��w2Hʖ�q	I���N�����:���	�M5(R���l�ͼ^�6#����2�ܸi���g[ ��d�p���3���N'�P��c�C]+g8�@�c�c�NOB�w'����5ڊ�݃C5��|D�@׭�],c�@�<���E�7�k���of�aGl�����g.Tt�:NًS)�ҟ��/q!jF�3"<�?#m����P~�ފ��|�/��JޜkMB����= Ҷ$�$�J��M��o�o^J������X��[D*�[|$*|� w�*G_�]���t�tU��=�䁂K��h��V�[|x�h'���`��ue�i����"��%��op�%H*���5HW*������7
�h�C��=����@�͘-V!�̀V��lWe���@R��8WLL!D����R��\�ݛ�.Rі�	�͏��h�;��}YY]�;�=g�r�ߔ�an�hz�����y�]�`�e�kҪxE�����셁��" �oW�Lr5��0����.�վ.�h�MTf��vv�Ʊ���-*K��e\�벆�}���h���N��
�]!�~(D����:a������wez��{	-εuw�j�46�Y�U0���^bD�0��/%�,k��qA��7�Ճ����vD�x���&`Ġ,OY#Bz������r��Π����Kw����77=�x��2�{3��Q��Wb���@
� e'�p�ɛ0��%a������q�:�{����k�v��4��ͳ��^��P�-j���i7�tN;ۉv�6�1��PWa�O��Gv1},�nZ~��Ԅ/�U�C}L��	�R�<�4��U�r�:�f��-�CC�b�u{yr��'�p�qx:�ߨJ��@��A�s�����	�WM^=+rg4Q�ZA�z=�3�e��P;?1L?�,\������k�C�I�k�a�{W���6w��k	�a�{�T͟+�:�fQ�%�q��q����<���6삟�1b�]�E�]��&��]�0Q�Q�M��e�}�*��y�is�k�2���5�f.���H8H�(�.��8^+:C*��S���5�������9!�-U�rt��0�Zr"ۮ�+�P�̤m�ZE�c�^5�7ܗ��y�g�1s�T���oϩ��/�@R��c�O��c�Uܣ��
�V<v�Ox\��+�˼]Ϭ���S�����b�{D>N��>��+T�5��&�e����2(����>@�OJ��)�.��^>��:>(����r7�J��P*����(����nBٮ\�E@(p�8*��1�.��xP�,W��ٶB�ք��Wvt��V#m���f�i�T��NJ"������B&+�¯דQ�(-�)�z���:sqk4^*��:���㐲]�����{�m�
NHD�K�
�1���*Ｗ����e�a\�9� %�W�޼����&sCh,G~!}�aB�OnI��bQ5.x*KFwC獎�j��f��#K%��00�!�VX뀦�i�'�����^I��� 6���k�
���iH���'4���a
�^��DUf+�w��C�:*y8��o���z��n��/p%��K�c�Je�X��}S�8i��#�q��8|��.[oÈ�4�Q�G�bDTS(Y����������:k�e��W@��Q�ֺ�;zL.��S	�<���ATR9:+i�"UMmH%e���	FD\��P�z�RR��Aj�.���q��o�)��.,����Pu{x�{Nэ�0I�Q0W'n�߃]H��WG1���<�0��,z�nD+��ʭB`���l�T��]r�}Vzc��5v�'<�@�^�=��u�d�q�%�롫&p֘��>*t;ۤ+׳L�ˮb�5I��۹��淨-!ҬqʨF_�m4^=W�u��f~k�J��ݪt�0br�{��e)ՙ{O��F���6y�u���Jd�^��1E{��1�}��^�U,�Pic�ܦ0Ǘ�(�6��u�
�*R�������A��T�(S�5OJ؋t��]ے��l�����5}�.Ce%l�Uh�Kԩ��`�<v�!�|X���-5BjB��@�8܍Ur�^�����1r���ㄱ,����DuL��9����J+�jw^Kjh���Ww�n�Hp���"�a��N�Y�.HQP
�%��T��Y�{,�}n��Q��1�v�wWnjf�ns��q�F������O!�0��9����g,� 5����:���V	�k�ݙ���S!��.Xլz!ab*b��g
�x�� t��u�<2����U�Α�]{׆$5Ãz��E�\�����>�ܮ3�.M@�Ip$t��I�ijw̽=/8�{X�$��ɕ��"K��9B�Ӹ��ntj�ȵ���]B|�y�wW��\={�'܇g��,��O�b�Hl��89�neF�����]��j�[��7
S>���<t'\������pڿP�`��)�1��^x�jw���c�Z�Ll�q��LvaNx�pmS^>�o����3� �u!�	��z8ƻ���Q�;�M�i�e�=�@�O5�]o�9��5�s��t�:c� V�����*�u�@~��3ܔT'G8Ʉ�sÎ�6��̈�:'��j�#[<��{Z�l�q�;K^���m4);Z/��g��MDrÓ]��n������u;�s�y��o�]1Y:�6TT�\�+�Zo�B{��t��-K���Y:<:s�{����l�Ed��Ƣ�9WK�I��m��2�]�OW��[��k~�m�̱4�����z�N����D�!�S�9�u���mܝ����M �ʕ�K���JQֻA�6��ת��e\Y/A��E{�zT���Z�&t�W�Jc�S�N]>���<�a�0���W˺cn��Pkm��UXY�K[�]Rv��>�>��zH��H�$���&���2�	�����&{�t�5��f�R��Ţ���iA�L_$][	�XG��$zF���SK����7��vu�7�r������K��kl�9��������-��b��a>OB���y9/G	Yq�Ypxw{g<[/Nn���6����K�E�6��л�Kx�{ܘ]P��זФd����]��J��٣_���s鱘�+<_]qK�s�|�:n�����U�M⽋o��7�&��Jި1�j_k�U�EC�ڝ<��A�/��[�{7V{T;�W����b!=�;ǎT޵sf�S\3u<��x�<T-r�Oq}AJ����$�b��ڈ�7
"��h\����5�M�r1���x�4's�u�S�}qJ��57�Դ,��rV���IǛŕ��=5���~���#��~�j��X��;�p�{�sb,�jHF5/,�&W�p:Vׂj7���(��^���^�job��*1v�t���έ̹�+���j��,�U��E�uw��W[��t5 �D���*a�нX䣲�D��9Z�A3��d,������[��ܪJ�Z�&�|n #o��/Pd�Y㕻�%����\��E'�E�8�K��L�D�3n5�v��F��$��ߡG7��Y�)gVƽ�z���Z��I�vK����� �����|��f�*�y=�C�O��b<��4dVI2w����9T��-R\��[Ow=K6�����j/z���M�t�9#��Q�˲�jGrz��o�d��WOv�4��{�nҭ5��+�퉚�7Y���Z�{:����'�����l`��p�-Y�o��aU�;��	#��{���)���)�&&�!P�.O�x'�ޅ�o�cssr	��b���]�z8g�5����Q\&�YkB���j!'˶m�:3˵��;�Oa����G�o����b9dWOQ}|wϹ磦ȍ@fLg;�x��'�I]��]3���ް}�����`�Y:��={�8��
��W�(* ��AQp��
��* ��"�
�tW�AQ���+��TA_�"�
��* ��TA\ ���(* ��"�
��* �TW�QqW�AQzAQ�
�2��K���'�V�������>�������zV��RP�e�Ը���뺷;c���\�*�h;�n�tͷ]�T�����ӭ���5�
n�
�n3��u��޽ɽҶ5�kjFɘ���ѕ�����3MH�gs�q%�kV��`Z���ִ�!J͡�(4}n�3�[���Q���Ŷ������Z5i�n�4i���Mj��J�m[m�f����k4ք��Z�f��͑V�����kM�g  �|Nl5}����=�k�W��x��6�7qy���ӯN�z�������z��[�����U�w��;��-Q�x�Mnݧv�k�k��|  z�[�v��w>��{j�w��uJ��v:�o{���ꪝm��U���v޽�ڧA�sݴ��n�#����ޝ�o��}���[l;�V��1�x  �
�Q@(��}�Q�4 _y���( x�   z��{�� '��w��ڭ[����]U.�s�فU,����^�{ַ^��W�^V4׻��i�O� �}j����<�LuU�m��UM��*�Xõ�P�����ړG[�Mζ�[�{�x�F{��W��2��U�痞���]��+emdl�a�]�  [�H���ܺ���Q��zz�{.���������� ˚w&��I�wkU���{w���gG@�1�4m^�YI���f�U��  ��
c_ovSM�QN[۠���\���z�Q���� �c�WZMD�ծXʛ5-6�MVٗ� �A_;4�SZ�u�F�S�W����gp{��x�S��4�s� �R�M0��J�  ����:޽�v6���{g��U���z�����o9���`���j� �X�vz�W���j[j�6�z��� {�>[`g��@w��T���:��3�ew�6�I�c8��]�h��u`�3v��z�MUF�jѶ�|  �
����� �9W(� 3�� W�霴��;^F�z�h����5��=y���|�    �T�) 4` i� �b)�)TU4`�d �L�����jUJ45jт` &&�M�~jT�@h�4h�&� i�@A��U4����m  Ci$�&�S�D���z4��4hɧ��?/���������7��Ow�I�~7��f]�uҧ��dy��r��3�λ����$	 �ִ���)$�C�?�����@�$�!���$�C$��?���?�48�gI"���$! �J��$! ��d"���Hr�������@�'��?˩!�:�ŗ��4�}�K��0�9�(R���?3�����ռd���n;����TH'�ֶ
XH8ժ:����+F�c�7Vi�ˊTM[��:��ԅ#��f�#y���8����am�;8u�@o
�!�z��n�o���H E�x���r��v�l���=O]�����_*�lՅkG��5��]�^5�Ս�j���OK+yX��:X�޳K8�׶���L'w��@�Qx��<4�gW;<:}�7�z�O�W��Ku�f*�G��OJK>9,�`,*�NQ��8�QaD�����k�~���7f�d�V�-�v6�Kִ:K>{��Yt Z�k��q+���cZ5#OF]@u�Z�m���r�sO��;���R�z��f�Ym�	K�x�e�TâAX-�5o�ܦ��GV���/GRo����'k�w�fX�W�U�`�p�Uv��p!a��>����b/2�x�b'�*�T�g,�]�h�'4��!�* 䆥<���0Z�X�ܴ����2	X-�Ť�D�� �rH�"ZX���̴C�̷�[W��D�ԓ儵���5u�C3����zлA��ه3*n��D�2r�E�9.2���b�]��*Om$�
M[�y򼾶+�Քr��PǕu����<*�'�]ݑ��7��R�v��)w��cY�u�l^�X���:�����wy��J�y��O9^1���+���+n�`D�=I��z�sv��dR F�7�N
E��v�Me͘�;�C�mcb�l<&��7d.�(���h2��]|�-���VWե�E��z�.�m�z��f���\i
[��9}j�2�sF ���D�Eઋ�2bo�Y��Q���	ǈ�nY���2์�h�>D�i0P���ֆ��e��w9a�y�i�N��+�&�$��n�X��2�6�jT@�iB�kn�
��e�V�W�n��y�����r짊�e<V��ސ�o/q�vhE���xJ�zV�%�LՄ�g
�{��S�CJ���0�a�_ݼ�J�[�i�;���)A�lV[֪�ggٹJ���yγ
�^��p��$2���^d�0�4N��ڤ���!�����x����
�Cw��gv�<!�]�#Vj�������_²���&P�q�ɢ���젇ݰX�V�������ct������x�X�Keq 󺵋CveҢ^S�ާJ��Hr�ަ޲�V�M�eXQ��.!�5��ma�$өt[�w�; ִ�Ի��F��XU�e��w���!���ޢ��S U��ZG]v��s��wH�U��Cz�Ֆ��:�JεI����v����uV�ˮo�+\0�����h= ee�ב6�:��{@1\����oFP��)��kh���7AV�u4Uk�r��<Z��'O]W�M�/�+U��]H��)P���Ř��沙��R;@_��\��!�E�Tl���4�Q�$�`V�a1&��bj�[8��݇�;��wi�@	ef�O��M8K*������w���*��}�F�wi_c�e.��;
#`u�J
t ��ݷ�5*E5�դX����e6��`D��
�2e��ʌJ���J�ۻ��U��;��&V���b��Ղ�_�Hkqa c&� 6��[����uE�@���5z�^��.m
�2Snٹ�S �0��ER�ز�-�|��j�këhgكhV�\0
��/���K/9lڻ�.�X67��5�t-rH�4��O:�apD�+1N�b�m���Sj�n�e9$����m��nŔ��+5�V�1[�iEi_c�N�������
��Npz��6l=w����V�[�	�{��V%t,�e[ar:V�Vc%v�y�z)�o�!-yoYL3��y�ˁ�![��t2R�}F����H�3I��^=T4!c��j|;�-O0WP�ܚ̴����2t+]݂�Z�A�Gx%u��{S����]�W^5�7
B���˖�۷��VA�ެ�j��1�ѻ���h��|v��X_.h��{��t�k��f��yj�m�}��z�Rik烃����������Es��giVJ�������¨Jʐ�CE㉨�YRp�d:�H5gyV���H�vČ���8�=��ore
"��ë���٣�����]�O���)7h�����l��v�]ȗ�e�x�Vv����܊oGtn%��{�]ð뫢.B�4�U��Z�<�lr5j�cփ�����ne0>�ԍ;���քn�i�OU7f���E �k����!���`==ǟ>�%[Ӫ���� ^V��\�ϙ5و
���;�W\N:�V�us�_.�7W]����'t�1|�`jO�Ջ��k��V�`�ǏB������2�4�a�hYM��6 ��
��W2�E�Gn���x�ߓ�����u��8м�J�aR���"�t)�B=)@��]}��#u.����aP�-�Px7����׀����� �7a�T�T��H���fn���^e�Ū9�7Z�o��'�.�>U�um�-���tVq�7����Y��u�n�_$�)"/h�x����+O�ÃM Id�Ql$b�i)B�I��ы�$SK�o��k~�qv2�</*�3c�c�[�ҷj�69[F��Ɔ�j��j�!�����eh�������e�Ov�4��l�A<@p{`����{�\�v]�K8-'Yh��4�Ն�[���������b�6�뀧��բ��m٭��U��w�ݏ}��e֒I4���Z�ia��E_��d�]�VMg+I_X[�ˋܷ����Q�sy�G�p�s�`��UwƉn��1i�i���k�լy��,��J��#ts����Z�{q���&]$��˲�ۀ��e	���JS��U�]�ٷ��A��V�pn���L��	��ˮ����o`l�5��ٿ��гkX�I�7�^�ߋ��8.�H�՜
)��,�� �m��⻣��=7���Z�̶P�wH/�bCM�3v�4�+��6�݀Z�M]+�8�%���z[:x|Mi�z]2��u�{E`-�+9��o��C5T��k,�w@�3���t�*+I�WM���w��ĳR���C+�aU���i{�;���4:��fkx휤���]6�s�{�k�['F��%���v���n��,���ٰ8�;�{�&)</�'a����+]�J����:�(g�7A��	�e��v)�cȘɨp�3����K{���Q�0����mj�#G^ ��ә8Pl e�*	ۣ���x�B�ڷ |��b�-�*'F�+N��*�S�,%��|�RD�̬�V��j[Im���W5ɐt�z�[��D�u�Ӽ����8��1������#Y�i�����o+M��N�-C]m�՘�|/�z,�3;1��r"��ޥv��t��nc)i��Z-A�+��k���G+z�n%t�h�u����s#�ʬ_ �3����]b<����s)02�kk�v�:��z3�i�j=B��0	����V�;�V�+f����Իֺ��b'/��u�X1��+��5S1n*�Cj����M̃d�Z5��hC+�b��>ӸoQYbŮ|��>������M-֫#h��y`^㺨XP�>�E��ۣ�%�,6�&��p�����5�P�(����[�)����W�X��&�Q�ɥY7)����.���*�w��A�ֹ�}j��!w��� �> �9CĨ�����h�Y��=	�t�L�|%���c-P��m���,���j�l�,�1l�*�xx�;X��m��}gq<���-//)m^��x��(��}�n�nP�5��H��[�)<�jD��C�N!,O٧p��x�g��i<ow��f��Ck�wX �ذO;w�5��e<�e����]���b�3ԵX��޾��m:�K1�k��C`��Y��ݻ�b��YC�#H��Hލ��c�4�;���v�Ҿ+m��*ۼ���{�Y\��f�����|@\l��Rk-��Xge;hݻެI�^4��th�H��Y�
�l�N�|��e]0�,�[afM�oqV�DV�a����;R:w��Va�5�IYueP��i�-VG;���e�<��Px�yX�f��v����H�_XY�qۢRz�@�?sO���߸�[��Y�YV�mj4��2�{H0Q�մ-[:KJ�3�t@| `2�Y$� и�n�Kv9����qB�-:�_�JU��Ho�2��m����r�t+@�u���N�\�2L%K�Э�-�u���Eyn�Cs6���R8�v�Ċt�h�xRb�_|� �,�m[=�os-֝�-u�³X�-�|�^XY�>/���oַ�{�i=k>
��;�6��ե��*�օ�w��l��nvm��I��kO=��ݓH;[�t�2o�VƚJ�R�]MP�$e�ܳ��i�\;Sϭ���;�C+�� Z���Y�P��V�+v��������
ˤ,a1�u�B�V�6k�]�XE�����]���F�÷�����~Y����O
s�b�&���v �$�rpc�vA�M���
E·l���!���o3e�ۍXJ��� g��M���>(�^�@�A�WK�&Α�{K	'���e0���]��,66�Y��}F���l�*/��B� �o�K@e�4U�!r����`�`M�+�[���	�Ǹ^Z����]{�<\������c|A?^�����Y��*Ѷ��慦�hǆ�-��v�	���-4o7op�VTt�1 74
z�w���&�qռ�Z�V״n���%wcN�n�44Ҽj�'���B�o��O�����3�91De']Z�� �0U��c��e�sk��Z�oubI���Ɠ'֕�V��^=Y�-f�����f��\�4��[X�+��ːx��=f�Ɗg�_RCz�4;)W�L�y��'���u�� ��d�&��S8n�C��LT0�B����W:�c� ���*�Gn�m]b��d&s�E�=���j�eЃ�J�NbɨR��M�.i��	�;�w=���g��O�5���ND�������B�@��H�_U}91U?T��ռ���-|KXU�a���+E<]@#�؛��Wt	��<����R�r�ƒ	j�u̧�gVnc��4�p[�أ�$�a����]�㋙b�ss�k;,�=���c`[�l��r,���>�}���t��V��V0�_�eyE�\���U=��[M���.[#�/��1�Z�C�רm.ias���2j��v��f��Y(�x��`N���)�Ɲ��E�Ǉv7�+��xm�n�	E*�y�-v�w����{u4����悗2j��c�B�<X�Z���_%�=GY�5��`���b�	���'	�7kH�R�yW"�v��;b{w�I�$R�s%ef��\b�M�=�2��n�{w9C}��&/H�5P\Sa��k	L)����ͽz�G�5-��-	N� $���r`S7bM�'�dQ�'v1�0侧YY�x����-r�o ����i���E�;�cl51�c�a<��4M͐R�;s�Y������	)7m؂喰��e�YбvE���fI��}�b��G���U�)�*@�r�'�q^��9�p��X:�mt�N��`%�u��$��p!��v����
8�#(��C0*m���A�]���WW�z�c�r��Q j������2�Y�}��1^c=�Y4��n��W�n�&P��}�ٚ���/x�%>i��\x�Y"����Z"�9J�e��뭂e5�,�<�g�Z�L���4�Y�H�j
��:޳�䮡B qaot،1�\�څ�彣Ye��u跱u���ח��$"��V�cr݅CA�t�հz]�HMH力��Ik;x6WE,�:��zԠ����/{�nnF����T�ύꘛ�r�X|c��2��aV�w��J�:6L�okV
v��5�V�U�f��Eb�����i���A�4	/Mk���ƫ��j�;�����qRZ�:(!�ܺ�n�p��X����3t��D*�>d�Je��Y�I'��<Z�c�O����m�	�ʺ�w'�j���II�+�2�5L`���\�{�.D�/��s}v���x.�Q� ��S
��J�Yה�!+�ܳ��h��+��2G+��.��B��P8�q���u��ᬮ�ѭN���Vq�ƃȴ0'��n_;w! ۜ��Z�L�|��`��'W��0#� �t�d�T�+CN��k2��38r`���Іq��-�n�ghݍ�^l �U|�r�WV*����+ov�J���j*���1{u�![;�m�M O�Ɨ3��<���R46������g�Qܕ�8�yB\��6���~�������L���Ce�Q�у4	Jv
����h�;i��[����%��t�>P��j�d����ő9��Ed��]h��} �J���(,����V�����f�P��[�HY�LmA�=�#�)ӛOF��k#]{��d�t囥.����A.��^im�Q�N,�v{�]!��mfϑ�χ�[p0q��r7Çٽ^������Ct���õ9�k�����ǰ;���D��0��zoB���D-��ŏ��۠�!����LoKw������\�r��XG[����.�Q�5g���.R�ĥ�KpWoV��B�9y���שּׂ����y7��\{]�B��oH*(�Z���|ً��8HӨ;���@LJVN�1�V��\4T�1����5fb����qwH��£KbE�3w�-��0����K�����՚�֪�Y��M	R��,����t&)�(��ND��2�r�mũ="��严���}P���w���v"e&�.j�K��@�s�=9����Xh���\3D�ۊ&���Qo����!��Yc~�}Mʺ��&uI��k���9��Qm9�%z-͵}XE-�v[2�(�Ղ�*ڵ��~WG{�7�Z"\����X��e_��V6��5����9�jI��bg�;S$���E�y��V"�E��k���ml���a,L��5q\���]m�\�������t��|�|����_�.�:�m"��s;Ii�V:�t��3���aSֱ�ZڧR�OnWq��L3JT��b�N��RH˾ƎNp��7Xv=X�	�7�G��\�.�� ��f�p'徤���u1gR�j�/���[�(�f^��(2A	�p89>��}y���cCYTr�*���z$���;�k��S1������詼���k�UcЍ�g;o1��KK~|-gaJEWH`��.���}F�U�����������w"�bWN>"��0.�ڏ\GZ왋�=�Z:ls*[l���`�]��*n:�t��u�;.f�ZN0ݥs�K���i,uvk�a��#�[Ύw3�l�❊�Pǐui9js(S��xw�Nφ��o��ȓ�O�a䈺��3f�+���4���K�ȼ�̣N��Me�J٧Vl ��!�ɵr�q���2�]pv6�#�Kǘ��aVP��ـ50�+(*z�Џ#Å�6�j��jP��n:|M#w��6ݬ�9��VR�0
���C���;Jh[�z�N|$q��Ȋ���4k	!.��Nh;}���ʆ�B��e\j��̫B֎��P(sT��d����ٷ�_N�E)c��>�m�o6���jr����Һׂ��h!����C۬ #!��T�7j�z�`䲆-U,�gU��Z���D�hL<E��x�-Z���ѝ�5n�^�S�E_�PZ
�V6t�t��^��R�7�0��]��9�D�#�P_g�ŷ�6�i�T�:����c]9��GU)�s2a	%��;uwX��4
�u	7)c�m]�jp �
��gTӦ�5aT�w�Uh����*��I+�����Z��C��"E�lK��{m�ԍwܲ]�@a�خ�a]�U��U��#a=����V�^o�T�L�;�.�t��ɽi5�gB�7��˹��R.�h���sW}���]n����%�h4��v�ǑH
�P�x2�u�+��ΪY)������Ԫ"hpȩme]F����j����9|��ōW7!;�ơ$h�֤����]��fثs�ll��Tr�'F�l�d-���<����pn
u ����.\gY5�Nm�ú��8�Kx�M�liz]�-�[��J���j���wK���2M�-�$3�U�-Ps���t���:�&R��h�4�P�3.�Jp���e,��|�k(ZEwk��L����iLa��m_�*͢�{ �lm��zw�b�/%!dc�Y=�8��#k;sF�=+��
})���Gjc$����GR)
��^`��3���-�tCG+�wv[��i<$96�ChB�>���n�7|y�b�a���S0�Yf���#��#��]y�_E�R�ي�5������Φ��jFNc9j$hT�)�3�����0��\���M;��B�~h�V���l\���Oc���Utt��4.oǂ�FI���o|Dy9��"N�<oë���a�e=���
U�`�uIq3��T�Kd
.y] �Vn�:|�tȯh�0�!���J�NH�/F�
n�̵1�p�i�Yk�r\�2w���4x�F6X��oo�XL������蚛�RuM1�3u&�䶶��ُr��7�/%��\�|�-�4J�ޘ�"u���5�Y�\4�4NL�:�=��c���;��w8�Oq��W̛�Yǭ��j覅�#�����z`΁�րcC��t������{r���v�b���-N�ú�4Z��e��'�Ge�̊���TkHEc�ibP��٢�4|Vj8.�ލ�*3�[\���Bݭ�x�V.z/7���8�㝍[�E:���V}�֊���)Q?geվҠ��:3�ӱwbnhIunq���$[8]��;׺Ǳ���EaRz�/o��F�d���tR��IX絹��0��=����$�{�
�N�ⱕ�R�6Ŏ�xẂ��bޠs6��aP��,w�Pճ�t=�lu�@9V�2L齄sם�w|զܽ�У�K@r�<�hh�C��w�,��+�-�}�B�Q�7c�	�p�e�ەx*e�j�<�K_5j�B^�a���`��Ձ�]#�� ��kD���4
�9�M5(UЕ��f��˻�[�"�ʇ�)�7�.��x%����}ū:>�$�%�3n��p �'�d�J�l�C�K�J��S��5¦$~��+��fD��/g+ɗ�g�jq:++zlvF�y�s_H%�����r����^Pc��z\zI�@�Z�x���kk`� ��u5�5�	1.��\#���*k��Z���n+v�%�EZ�y�K�۴zˬ�|ef5���v�����f+ g6���0h
�9w�j־h�7���ʷ��Cԟk�f�,��070>�f�6b̛6�7t�C0�yJ�'u���B����Z�
ݖZ�^>���K���Ho�ԫ�z��l��|�-�Vt���N�+U�q�u�6./��Ql��oM�t�1����݃Y��o����m7�L�g0P�ٕOv�9���OpT</���X��u8�y�S���nf����c�U
B�K���t\h���[A.W5I�i
��x����>�1C���\p ���2O�\��EnQ��E�]�K�4��}orђ���n�J#8��}z`ºZ.��&�m3� _p!�zws:K��wE��s�@Uԛ��&[�
}z�fBU��Uf`(�ޜ��[}ݪT2E:��K��z��Ҋ,�萖�ٳp"˒�qɒ�i�
�3Μ�0��&�z��qvڹ�v���rGFє�Z%XN9%dTZ�t[*�WNl�Z7����yW ���%g�$Z�	q6YU�R��R���v�J�R�S�C��BjcK��ԅ��^j�r��e�f��.��x)J��̃M=������'h<���Z"	��on��E������f��wݻ
�hTu|��ngHio���h.�zk����ʉ��@an�%�`���1��5�������.�l,��F����~��,a���#������	��Ox��H@��s������<=���?�X�>w�c��;&��:����ظ��#��>Tqu:|+:�)�����&a�/���̮��l-����K�V�u>A�KUe^A�:D��1 xh����{8$�9#�<.�Krbt����,rFf�cI��i��㶬V���PR�y�� &�ݸ��y�G��ܓB)��;��M��<4Y�pd_�i5�i�/d/xʑ�6���\�����z����G]�ӆZn�[��O)�'�E�R��W��u
�9Q;΁)��u[��	Q<5����R��}p�7\	p�`U��g�}��G��j�^+����4�U�r�*ѭ*��>�ӱ�£���u���t�n���%t�^R��.>q�#���~{L��]+8�A�D*�
����x�,�\@V��s;��Bzڧ����wG���t񖕡��Fպ���(27d�������ql�����<�,v]J�IFJ:,�_bd}�z�aS�8CV��Pl����K$Q�[o���삪mjX�_>�T��Z���ʉ0��]ۙӶ���HY[N�+�Mw����et��.��d�g�����[6�,/:�^�R�:8�ɺ~֚E���
4T�70^mt�q�|�_X�\պ�ڹ��R������Y�Y�+�u�m��o�wP���q_�%���(�lU��*��;��8*0{.(\ �@26��LV!�t8ւ�V�jԣ�%�ֺ���c�j^Hp%��޺��t�MѶx�K:�����\�����t��se�Ne�v��k:�p��Z�j��k�xNn^Eˍm��)�m�3R�)�ڮ�r����2dR�=�YWa�ŌL�죮�0w.������:�`\^��xR�7�N/�wp� j˫R��,;M����O�wb��lؖ�&)�7�Wtv�v�s�x	�ד�`S��PQ|A]*�q���m8��c���pC_Q˒�(p�j�vK:��w�0uWn�]�A^��yo�����i`8�9�к��k��z�:����x�� >�p�\ts�����m�N `�T�O��/���!b�+{��Mט)�f��j�u�9�7h9y5�u��mOJ�����QK����m�8�)"8`�������o6g\7��n�����s^�ɖ��H`���V���q])xl�U�jZRd�pՃ�ڨ�{�E�1�á���a�ecƹ��'$���ʶ��o�S�؛�_Z��k�k�X�Li���Dշ��0�m��.�bPj�ޮ� ��klv�o��7{��판�n�jZb��C�:�`�S��A�����T5��g[��m��!L<T��[�]�9��d�q�\��w�l�EV.�;j��sh���<4��a�ٙi�섊'��)�hlh���Ѡ�@��Nc#��� gO8���wmX�|�n�"���K�e���"��{~z��t����h�׺{�׃�>����#ie��9O �9��[����̏-Y��XAF��#�G�e�ٰ8����N�!�������b^:�WR����î\�8<#{�h�qmg�p�W�T ��a�|LDJXb�w;��/��G���Qn�����ǋ�%]{��Ѧ�\4sb������ր�E�OoX�����;�a�\�c6�f�TԱ�gh��S1�ATA�<�9��Q�Z%S8���7�[ͻx�/_��33mw]�g5Z*�r���+3�&	��[
r�cv�щtGM��Cw�LKt�5֛�[��V�hɒ�+�6���J<����D-V�Xm�^#e*vf���գ�ev+δC7��ό�,^��e1YcE�o3�w�'����Ӹ����M�BK�P,�(������ݪu�Xt��)u<��P��s��ᷖ�1����a^M��;��K����hBr9ڍ2�U�+����^��ԕR���YJ_�K�<܏A�V�=�'y	j�h�H�8b�Y�qyh9���kq�8�gm.W k�䳬���GZ�W��d��e�b��P��[�f	�I�9{n��⍧ٻ�$ByPu�h�u�5��j@bݪw����q�7�L�x�˵���Π�h�xMjm3�HQ�u���,$KW"�2ս3wp]���y��C�|�=�uoY�������T}d����+Ek3��Vn8����ͬ+�>����d}2�gø��
�A���n����6K�I�)��%�R�Z�Լ�RzD~��7��N�9,6sN6�q�[l�.���uʂB��cN��Qe]����0N�\��n�"��Z���]��E��Ż,hۓq��5>BUљr����CR��յhCW��g+S���o^�@,�4<�����s�Ǡ�֧!�����\���n�_m�gF#��m��;�`�������
����S�eɐ�|=�8R���	�������O+�Ɲ%��;U`h�sxݙK/$����}/�5,|!���B�ҮC��v�x�e��}���m�b[�r�'6�W�s�J`�2�E0��gB�{�(9�i%���q���űI��� -��]��ލB�>�A5B2�񭣼&�Yw�U�Î������H�_K"�����<2�KUѴ����Z��]Hh�	w��\h�hڲ�Ф�fU�$��%�ڱB���*;���l��9k�:��ڧ�39R�usP�rS=��T�|��MI`��a-d���f�mP��ެ�ɱ�L�0,�s�ʷS�[��"0	��MY#c�0�.ͭ����͟1p�Qr,��g,c�q���}V9bX*��ꔎf�ܷ+h����j��zҦX_%�B���H ��&���y!�N�:slN��]g`H��.�*U�v0�Y����7��s=�[�Ѫc)�z��5���2M#ns5s(�H%�{���W�4��R�)j�\��E�;Lל�Z$w���	&��q���PU#u*a�� �� &��$�K#�Еq�����&�u�p��P�a�}EH���ѻ�����Y3eT8T��q�!��N�ܤN_u����:�Ԗ�,m���noٹ��l�TA&�Ӽ][��Oh�m���I(Q� Z��	����r��_�=y�;V�Mr���l��<�V�͡�
	����W"��dcoҕ�W��ͺS5.�*R�P��
ح��D7]$���o�ki�B��1�������9�*������s�8]�Ky��os��!h�l\c�2̡G/�-O�5�� �)��۵m�����0�b���e��.A9��[�Gq%	@& ��OucK@��.ڨUo���X��v
�x+���,[8)V9&[ജۥ�m�����wsZダڒZ�h���5���O=Osz�;B>��O�g7��k����ͥ0x�[4�>+y 1�{�J���5;kl^�`�UvU]�"eKḃh��	����髕�j��Z�Ófu$b�Tc���H(��u�ɝGf��Օ�kyV8�R��9�o�w/����JfQ�A�u+_	w��0�''Jy�P�m���_ww#����w*Q�;F�U�J�e� ��O���X��l.�WCI��r�B�������W�����|�
�khϹ�S
��uo����;�ONU��6�i�C@|"��:�f�զ�[I���g-ſ3�[�+ .���X4�к���t�������E�/8�ę�w;���RhH�fԥ�[��j��n<y�/P�rBjE12���ҩ�uƬ�U��R	����'n���u[$�j>����,уE�.�I��pj��\�v�Ysu��N��t�K1D�T×�ӡiu!��]+����M`k�Nh�n�g��8���<����Yu2��Ŋ]u�KvZ���DYXI=��-F�oh´�i��*�XL�.�f��8Ԋ�A�V �L�T��o�U�n	�8QX�n]ӏdeat�k��^�j��������5D�Kb�j��oq��{j�j�cE���e�]w�k������@�5�u���v�uf]#v��6��Z�����3��n�;��Z���ҽZ~b�&�8b.p��z�v���!��4S"��'Z����lf��0�e_;�\ص8P&�%f�:fҤ��ɼ�sk����i���V�� fL���eS�����UaϞ��ǹ$����K�2!6,v��y*�9[��t��hp�Z��R��3:�>]( �Z��4Qd��k��Y/�-M�mc��qE�
�tR�e&�F���5*�������#E��h�E�����]Knvu�Qa9�p�ё&�]uہ����]��B�[� ���x�`J�_u�m�`�%�G �y+q����n��6-LM�4��{tJ�"I�|�N�|����C�߻U�Z��F���Y�9\t�x��m@�ȵ|q ���Zy�I���m)6�Z&��� � �}�ٍ�[U��֐�.X-^����W
�jT�J-*�qC�	48l%�Y
�[gq�ң�+uV^�?iaC"�Y�oo;):S8fx������wS36�-���]w x8�������]�Bg���+������g��1T5/q���)8���Ҧ��};zܳv�V����F�N3��ѱ�.wY�q:��}EQ��MF�J�!�i��fW_1@��<vݴG[6q��R�		!���_wP�����+3��v�,�t��wU������X1�Vb��ut}�9lj����R�s%�r',�
y;���w#����0�� ���h9�v����W��G\u�%[��6���m��p�e�3�TE���l �XM������RjG��(�&ŭaDĬ��gGm7kH@��[;(��u�s�a��#F�~4�M���jE��ǝ�e����l�T���a��YE�[��:ᇵε�\i7�g=U�S3iQ��(�4���Q`'B��R��t��Y\�y�U��q�e�g&V�A]�l�xy;�oWˮ՚�I��	Wz��At�ܵ{��j��D���*��{�!�
ȿ��d�>��,"|(�����R�?4o���,�=�U���PZ�.��˼"��:�I��i�ѥkze�J��u�G��n�*������QtԔá֗%�Xlf'{O`�P�5��y��PZ�xF��o`|+l�@;��f)��㘖չ��mm�XGs͖NF�������q���B�WJ(��PsX�gh��\�"Zi�ǭ7{N#�G4)��+#�(q�+z6Ab�GM��TA�Ԯp
�ٿ*T-2~W3,�^�]p	Y�=|���p�R��+��,�Z%7�w��D3*� �*MZ����f�2��B����Z2�q3���(�E�!zz!Y1�N���r�(Zr�^vM��8����7�:�!+>H1[���a(�����v����"�!�w��XJ�z���Y�s���se�����`��]��w��'�v�d�b!�e�mͽ�ӤO4��ڊ�l41�M���N�����Q�Ám!��̂
�'+�m��f�H��2��hWI�-��nk5���c�(�����0tخ�i[-ї-̥pq���Mfc��cL��QsT�65�q��ӦeK�4̕�rfcr��5.����
*�i�N9un^.G8��k��4�Ȇa\V[mm4�b��0�S�E4�:n7)p�Em����E��e˙i��Kh�6�����D��,�e�\�V�n��j��i0K#u��I�\f6[TZ�ƴ���*�㕬ƋjX�eE1Dj���0ix�kN8`��kW`̲�WaLVV�.ZZ-J�7.e+Kk�UˎV���PjTjڕ*�X4���ж�LA]f&]`��U�(�Km�ƶ���VZVik��:�d�J(�U��U�
�F�2��]h�\R�JR��5��J]9�5b�U�*��m�Q*QQ�Q�V�kX�A�X��[Z�X:��]aKR��.QE��(`�.�f������ؓF��&��t-�";rɍU�Y��u�]{q�oE7�Ҍd��3cv�7ZH۝��ٜ��b�������l[���5���2����ڏW?9��{kYJa;���\)�,��/+���!g�Ӈѫps�|K�L�Y��죁�;�$�l��Gy��!��4�fyq�.�2�gcMl�i�~�}�7�OƮ�0u
�#hH�|���M:��`��{3N �#mt�1����C5p;�¦Ɛ�h�,]1�*�Rw�Ǹ�{
X�5����ra�x��b=�1�s�c�6���Z]�z���N1HTM?l~:��K��H�N�0�w*�H�9v}=z*&{3u��.�\�#���y���X�=�)>WjOF"i.�$�8Y[۝�`&��j!Gˬ0�I���z#c�-�)�0F��p��@C��-���2�+�A��F{�)V����*��	N�=�|tS�����븓n��WN�
Q�=��Z�*S)1fP3n�mU��_=���fm��JфG��Ź��NtPsł��n1&�'qF>�U����V��A]��E��b��jtp&h�2t�!ݎ�3V����Yrm�Uz�isZ�h����^/*��ʤ��
^܌�+��8t�K���P2��i:��zK�pyZxm8:����Z)��±�-�;2���TwdK=rS���T�;G_�3��6#����jsj�;�؃�
�\�&ts�H�H-����o1�F�a�@��<��#���O��W�,��N)��2�.-NP�!��P���$��4��H�Xײ-��,���攚�и���jq{�ӃqƩ�|T �5��ķkvE溓U�6�`�^�攋�����]Ss�&�ը�1
��3o!�"�W��r_.1���K�#ҷ��ЮP��F��_���B �SK�'5fii���0�I|���|C/L
�@�N��Y�s��`���R�o��=aRBWNWQD���uju�}V�.Q�˖| ��� 2si��~0�,}��Z3G̛Ϧ�p�ьZb\}j�]�V����.V�=�AYH��	�:��u��Tf��V�ig/]�+h>Y٬ux{D�y�
�8%z�~|�Ȥc	\)�`�]�y��b �Zr�%(&�_��)�����{���6ḇ����U�)������H�����#��'�@Ug/;67���/`�tRky3�Pˏ�Mp��Q6թ6�kspiK�Q�k�r�HB�&hj�4���Gj�>�9ǋY2c��MjFZ��:1r���=,J���sW�du&��9�7��RX����O����F��ۤ9Օ��g�p�<pp��g" ��s�=.�^A�A�+��F�r��tG��Y���{+nd)uYY� r�x�ٓDa��v;*�~^�-��<��<�e39�fMoq��J�B�j&�规q��W�l,����1�c$���x��A^V9�K2H ���,h<b�Ƕ*�����K.�s��R7����m�\���'�	(��$gM�f�֥/� ��rW�F$\�.^ț�f���pk)9���F��rK�=H����������
��O��p�_�.�v��Y]��՝��&�����0��(5����NlϺ��rC��7���4��4wW�3�Q0�/pՄ8g�����_�Q�W�:�FMv�Q�G	b���dF�X���h�$P;�Zh�K����WbaS�u8�Tĸ�E\Ńt������}~��4:D;����f�*xZ�U��c�$�F�z�:�_N�84��p2�L�M�tej������o)��@�����@�O��d���@�57lEFm�vI&:o��1u��?;�1�Ҏ\'��^cWj�O�΃,UD�gk�ptI��"K� l��%�3�[����nYЭ<w~|e�2=:�����Z��,C9��}Z��1��c��K�Ɠ��t83y��C��F����뗺�y��̦w]���e:��66��xqn�}��:i�݁|����-��a�J�y���[��=[8
��f�(q��Y"�ɝ�d��ң�zՅS�[��iб	[�9K�]ɔv���*�hv��]�,�H�]V��j��1�Tj:�
�)Sͯ?*c��ھ�t8���b5L8B�^�=����u�F�8eq�/�t:Z4;���6m��i�@����!@蠚�~ٮ�>�c/ƀt�
(���e��������g� �;!��������?*f���o��u@��p�)$g�bU�@����������B�!A��A�"lL�+,�ƥ^�ڞئ'`d
y�I�4�s䣼�HBC-CA�hsy�ί��7��0z������>B�_-ZhhC^3h0������Td9��7���ˌ��/�	Zc��͡܃��CcH�N[�[S}y�	
H�� �4�0s�ywH���|�����9�}�N��Y�=\eot����E�h^Z;�EGY�"4� �]��s'K-��Iwt���b�bvh%<���K�i�%�})\�_K|�q��Nӆ��83&�;��^��X�����ĺxQqSƾ�"�#��'lPI����6�E�r�d(�K�ȦX"N���X�=�&�r�Rx��e�U��=�݊��z�v�Tn1	A��a
T����Z^���j�|y���M�2�F9.��<!>Ȕ�V���l|~A�X�Y��v��x�+�1U��V�!���3V��L�"NH�a)^�͆����l�z�8G�,��F�;G�7�WeGXo��#ϞI� �8׽IXk��F�6����� ���Q�6Յnbi�b��Y�E__H%Ɯ�B
�"����vx�9u����A0w�RՕ�8����bV��ś�;٬bQ��AP!��A��G;1���̻�[��I!�ح��B�^UR���$��4�4:�7�5���u>&�`�[�c�=<I�_�������cK݂�y�]�G�X�r%�u�w�W
�-�Z���I|3��)�U�r�r\	I�]�.Y��9v�UGT����y�ItI��˫W8ڼZ$M,]� �^���xy�_b�|X��#V��N)O�ϕl���W][�Jur�!w���I���1mN�W7ܤ��F��GI�V��71 (N��1pu����D��!�\��@���,qӓT�15�ݪ�QC�Z|V��ϲB�iڃ�b9d	�h�(=.x��=$�a�V����ᡄ-9X��4�����]�VJjsx��DZ���h!Ō���z���֜�J{������Nm_r�-��j�L�d�\S��,e��ZEϬ0�*���L�y%=��ٽ�A�9{hqGA`JxE�gy3:�rߌ�$R�VyTFV�n��J�����G���TWF��� 
�c
��.\�5K��;/��=�}�x����!Փ�񭲽�M�m}�_��U�K��M�^���LWY����T�F��O��k��7Q3/��"󖄬b�����^(p�17:�ҹ�fA�^S��)Z�]�V%(�F3v�V��'n�@�@��Q�u��c��O�F!�{c0���Gu��\�F%q�^жם�Gx��0�丨�"�2�T�|���Ъ���c�;��w�G/.�rA!�,��� l�mh�gF�Ɱ���t�&ʲqM
��<��<����:S�6�]<#�j�-����"A�m��;Od��b .FD�;�?����ླ8Ӹ�7P�)v/&�;�LÙO6���¼�:��m.3o(�듔�/C���á;y�����L���/|��*��X@�a���6�vK�\V�je�����c�8�yp/P40?!h�i����j+�)���\�s��2¹�Tb�������K� -:^����U�<�S}��uB�\�<#��6���4��_���^�]>\�G$e�n>���v�L�f��ގ�_1�Ж������:�ur�o��9N��u�����'�Ǡ��v���G*�ֺ1�=Y�0R���]�޽\'�}ԓ��WG������S=��:-����w(�wj��b����j	9����I��bLs�Q�(lۖ�a9��;j�<�����bd�`� ��9���Fj:t���p��A�e#T�o�8�A�7�l/^��"#̸�[�hD8�yIW[����ũ�Sq�E�jԈ�^��h~@��ܤBgr�mv���m�8��}��5}u�8��
�
w���u�*�z/G���px�Z��h�}�.�Ǆ�.�蕘���.,�kN�6/Y�
�P븞;��K�t���0p��:�t�Y�Go�U�S�1�ݴ��0�>e;�+�è�#nUN�zܘߕcj����g�^�}Lw�k��#=o��C��?=B"O��	B+�)�º˥g¥��6�����F�$v�G�D]�ݭ��	|pr��1I#��۴f��Y�jRWl�c��H�S�����W+�m>G�c�7ZӮ*m𚹬��iu���i���-�;s�z5�7��T�E��U���.��p�{�%�#�A�2��^T�����M����_c�|þ���şAZL�_{����V�׌���0�.*�y��ޅ���(�3	Zcdty�;�z� "�M������1��Hn��M؎�R1#�������R�.��[�@����
B�3�[��lZ��>l�8������}�@�H�@򵻧`Z�'{'Q�ml
�zlC�9�Vz�J=��Uz�+��E�ә��gtV��1�6<ĢwP1�,�Bϕ�*RGd��J���f�N�]����c/�e�2�.��<!v8J}Z���4����I �����ފ�[b����p#:��%�^��)��,VD�K�v��&�f�e���hr�Ԃ4E�.���;ʩ{s��x��W�O�/}g���Q�����[x]��{
ș4\�Q\����KO]��B���.��I������M���f�J�w!���q�:Ӥ]Dλ��i@��&%�%�3��M%�\΅�mSf�L�z���}�\��e;�7��.�Z��q�������ǻ����/y����F�[��3�mK��(�	>;W#�E
;pL����*�˭.�g����I]Wf���,���
��:]���{S*5O2�8&*�SMRp蕷��0v>[�a*=�X�7qYh	A��<P��ٳ�����p2�MJ�KOK��q]�Y��V�:j6Ø��İ����S6�(��ȅv�X�
�Q߯KYR�%iu]���VT��d��Ʋ�-�6��󛮨��TM
p��ڳt��HJ������-�*+��yn��n|����	�������ud���"YFv2�h���9>������۱�6Ѻ{]�p��w���J��}��s(LM_uI�l^��9B�yΊ��n�,;R�2�аje�t�GZgV�6pWj2����bM��O�Y��Tp_=ެ��X��?C�8�X��B٪ǿZ�ޜ͞�"���O�<e�Sf1k����=K�4��LJ��u��9�l����Ùu��͡od�]Y�{�2�9�%�a��CtT*K	-���b�¶(Y��OR�`���z��2��.�~uq.%m�eS5����KKб�gϙ�Ġo���ua��CT��n��u�kX�Q.y:��HBm8Wh�ֵ��Q�I�:�fc�B�r�+�#ή��D�h��^�
�`�M�N�m���q��>��"�u����x��u	��x�\�J:o��:�i�N����^E����7�Y�r����|b�U���œPdbPn�td������;Wx��;����D�g5v��PN��4��K��-N+0�t/D�ו��+��Fc�r�r��a�DYG�^B"�e��nzd�tWr����ӑ�58k<��|�Ε��T��GH����Z�kqӇ9M����ԍ��l��Ff��/����*8��F�j����SsZ�6(���h����|B��d�$�� �Q��hf�W"�upȺ�+1q�֍�
"+-�5�WQ�miU̖hҵˌUL�m*�V�90��)[V�Y����q�4�V6�Q�Lh��`�%V�Y�2ڶ���uq%pզ�Z��T�U��%���4X%m�����b�pA�-��ڵ�YD1m��[��P�ڙr
��2����VT��4�e)Eh���-2]9�k+Kf7,��DGT�գDUDjZ����(���)m-EVU��ն�m�Z
�*�j%V��(�5I\kR��,��.�"`֤e�ul�J��3(���m+TmcTc�P��*V3"9j�-��G4ي���ʍ�6�1�����[J(֊�kb�-*�[R��D���9����7?DdcJ���۹G�y\�)vd��l�Gh��s�I�_�{W�������V��k"K��S���`�q�/�Ud]m^)jΘ��1�Y��W�\���ٚ����Τ�%as���ӑ��
�EMA;���}�/�J�ohBy�sjEԼ���n�e9⾰�p0�P�< T���]H7�th��_M8�ϋq^�u�;�U,��R���^�do�!�ht	5<����6I�{���2	j�����_�����yx�J�i������GhV�0�HE�ƭ:麝8���T��!�;��/%˗��NQ�M�m�E��y��"���k�u�5�sX��[}ޚú*ŎZ|V���:9�%�
�G���˹5x�����C �)`7hj]�����bC�>AˌQ=�:Q.wwҡfz� ��'���DG6*l`~��Y�F�wn'!79A�[eȦ�J�W�4/���$u���e��ɹgY��E�KFRն���YS�/ރ�/Bș�o虱_�g��(4xM��+�'
�, ��3z�C1�A���^��E�G�а�Ӳ���G�y��}�-�ш~,�J�����ݺȆ��J�^�@�YtX�9�a�G~�#U��zi)���x]��<�>�~��PP6��z�>֬V��0�;k��z%�3�Ư=
���k+Z��z����S��*�b̰�Dd��B�)�^|z�{4���ɿQ�$J��+�������;:z���i����Ŵ����C���;��:#Hp�^k��m�^��T�\����o�j�Tnjb���/^��#*���0��E$���㑈C�W�놤h�z��llz���;Xu�����Fc�n����$u+���h5��uW���Z�����+q�5xH��0���\�k+�7���Y֠5�p�Tq/l�0�C>b��\Y�̘��d�m,��T��ø��bƌ �*G�8�9�EeB�1���n���r��+�s���5J�t��Ѭ��*��h�Gwt��'�Z��HqΣ��v�i����V��+�&J�5���Foᝅ��&xf�#�"��V~��t�|��yEgKoE��z�c*1K�P�ԯ�j�yp/P8�є�WbrZU�ׯwYҔP�ȥy`ܬTb�
v�@�̈́c�K�/Zt��{��]�Gfo3��L���]kr�#��[�p@Q��J4�a3�V�U�|��FCn.T�|���`�c�YGE�:�#r�<��z*��{u�>���I�F[pgi�5;���/�
��/ �U�������d�^f-^�� ��,1j��̨�2ݯ�����,IØ5e��zQ���=Rs�T(�9S%�U�aT��-��~�"��Ǘ�˷�ox�����U�����"�|�4�X���*�07e��A���o�_^�φMz�P�� �>h+�B������:����.SʮX2�̨��rۑ9%fP�e�dA'B�B�-λ�΀�4�>��@�mff<��b����j�}�ũ{�s�����yҳU⾙��4}&.�u�&��h"Rb�S`��rN��Uc駷�*�3<~��w(��U�N"����n��	�����L��ц)�KO�%e��_n���A�ۘ�EHReF����DM���i~41�A���U�ǰ[����j���i���v��h��W�u�u_-�;�^X��C:vC����_`[�"k�x��i�熢���B�a`w>Jy��$2��wSG ����h.0��姌Rc�|:�Gc�r1K�J�		h�ۮ4�m�lYhrFS���"Fb�+Lo?*C�4�^�:*7�=�F+ty='LV�d��c�6u<@�1��0s��˺�~���bv �ﯷn��xO1J/�H�qX����Ҍ�L˹
$��1�,9Tq�,�:�3"&p������y���*�I|Ǯ*��p:����"6�h�]++�-*�YbJ�RTV�����sv�V�9�/w:�:o_];��Я��6�׻��A�Rc#/.V�I:ܒEP�G��ߐԧ���k.�etw���:	�풬���bG���b�A����b�d�����˦E��g����Գ	���dWZ�b�ҘǄ&;"R��7�9Md��[9SYY��׉�\�A�z��A�Hg@Ȓ�z��`3\�g\�f��J�1�� ֺ�'�Q�]�ARs~��&��j�:�L�b;��4���q�Ǯ`��ɀ��$l�^��s �p$��窳�s���kH�����6�v�%Ɯ�B
�"�����rpr�<�gTr[�����"�L�=n{r3XģF0���CK��{[�4�}К<�W����C+�(�r:������!�BƇ@���r�Tvv���t�Z��S���=Vf��������7�/rj��_G�;�?�рo ��D(6��j�7& k�W��7?��K]��C��*D���;��Y���O�4ce~���ofk�2�=��m�r>k7H�-����b|�:�e�S	��;��3qΥE�*n�nI�)qhl_Y	m�b���0dw0�p��pO���>�$5�+՜�8@����ʯ9���^Jr&���D�O����H��n��4��`xl�$ 5s�"R�"v��Z�-���K�$2#�ɡ��7仗��.ӕ���4�1t���Ӵ�b*xꝍ�,uDS�3� ���u��b#��yD��_W'�{��H�
��:cB�V�;�	N� t��/,�_��1g��E5�����A��D#�J�ƾ��t�8��lY�L��۾V�epy�í���+Ǻ��ț7J�#'#_��&y�=�}���Nh�����iMZv"���h�S��˕�[c���@nʉf�%�
����|�:cWk��{� Z��a�
�!��l�r=)���A[���vj0g��s�g4c�~Ŵ����a��Ю���_�jQ�N�ո]������w��~���,���J\�����\;�a�G;ޒ^��C~
�*�Z
]�)����{��aǡ7� �o��>���AnS�2���þ�*J��NI3j��*�3�����ޯ�ՁC�]���a:ϔ�Te!qW��1��$߅��(�x�л��W��ا�>Tb��ؒ��ġ��B�QIF�D� �Q :�������������4�΋�������ۨ��փ9�X:�8sب�^�7��_��R�\ׄL筥<6�J��7�i3�3��FU��Y (1�t��W2�mF��'.v�>�\s\-���k�~^�e�̌&����ح��>����]�\�Ϭz꣘,�ܗ���d|����N��#I��)��{W�=�2b��P������s�M�v�n������p!(��Ɉ�O>�v��@���.	����e�nN�]h�u�E�x�)9�3P(����8�|�E��R3C����#�FW�c�v��H�:W9Fg,�Ge����!��P:*P�o7�m�3�Jg�����~5%�z�O==�e���;]���X��[�N��*iλVҵj���:�Lg�h��D�������*e����)��T�K�����g�3+鮭����,ɳkX�B�;iH�cO�U��Ϣ<�̾�ٔ�v�CU�7dtpޯ37���R6��
X�Y����hre\n~�Rje�%?8�ġ����͙�0��Fh=�:s�]�U�ƙiF�C�PZ�_.�L8[��%f*!m�4tَ&����6�/w[j�_H.�f�.����h���V�<n��9
���7qϣ��凋�/�1�@� Զ7��`�F,"���r���z_�0{��Iv~�H�6���)�V&+�����*d�:1�C3zh�[IA�c��׬�;H�.�_�<��
YSzؓ��[��.��F��kC�`}t����OƝ���QAićb�}У{�u�R�B�J��RB�������7H�m��t3 �!7P�uf��w'י2�8�	ţs��@�vuu�h:y�PtxF�b"fң&�]^�\�Tko���e����{��͈�"�M�>Pq�h���J�=m�5.'�%ӷeN_v���C�����Lb�������ٷ�b�⋮�ݤ�M��r�����}�QԄȧ�0s�BwBU��DJ93y� ��Lf�o(�gG��z}'d7�,r����"������͟S��t#��I�A_��(�BPl��Q�;+P{��*t��@[_2fV:��U4�u��<xQ��;%�EPVևl�կ};{`6G%��	M�9�B\�\t�tdIbנ�QB���!J�ks�\���;<� պ��!V��!�V�^ܳ~�f{31�����-��P��G�F��B,7%Rz���=+�_���3EM���)��y�����sԍP��;�\�n�&4��J���n��Ve���W���\낢jQ�|rP^�F����$� }��e�\]�4�F�{k��C~u�RӨc�9V����ne;���'J��d.25`�j䅤s��ZK�K.�CyL�s��W| �2�M9# �ӏ8�9�>�#r�ZZ4c@���4�b�t��KU�;�q~����dgzGA�G���A��t�
��jpFk�{���C*�	��$}�*@��>�٦��¢0N E��Y|���Cc���n������X�n�'[��*��(K���*��f��x�p;��Q:@��t_-7p���p2�Σ���U�ky#J����8����{��{��()ك����_$�7�2� vCZ9:b��x7^�P蜓��}�J�O8z����}�[1��(��q����2rn�g��g��V�ɼ�~P1���ٯ,ҪAOh�c֤<�.�=f�߶LH,�y<�E� D "��w�-�Do��_;�\a�bAk��X�ީ�$��+3�& .���L*oty���a}��yI��d����f$�� �>�P������n|���ʹ��������B��=c������N\I�TY�Y19dی8�2
A恣�����ͲbVz�+9aQd�*m�H,��m�i�P��Ŝ����a_��կp(sWB.�����~ѕ������|ڍ�,<�z��t�1@�>�ƕ�[�[�Âfq�OǙPWY֊��ns']�q2"�Q��S�O�u��B�ˣ˹ jVn��g5�Y���]q]e�=���P���J%�z� qC��i0���K#K*Aۚ����#Sd��z��qmI)^�;JU-�`+�7/ z��4ힹZev4�&<�g�Ӯ�;E<d����yW�г/����ˆ�{b.<��1�R��,��:���f��s�
��nNJ���;���
Bwh��e��%���p�۽�dJf�T��K֍�vg^�o����:-CD�l'&p�b4�>�����ySY��AX�"2s��]YV혮��<��{>�h=���z�uI��9��s���W0B��k����y87���<%���S;���[I�Z5�"�y[�(��_)Au����c�+g6����{l���X#
��\�kym�9G:���c�'�WB�q� �<1�\��8q�WS���U���\��l�ͩ��y�oJO��O^�����Ryx�/b1w�^v���55�[Êb�H�v=uz0��.Rn:���޴33sj��q��mv[R��W�W�n��`��D�4����#�-`n=S�����x�YI�}�����Z�݌� �q�oq���s'^Zh7ws�̀��J-r���v۫A�e�8�Kw|����znxl��)o|�çMnӒfѠ��=����^��-Қ�mݸ�����{kYL��u�֭j�;��Ô�~�ܤ�]���f�8���o4�\�S�)V�%<���� 0�ΥL�♷v�Z��<�-[��l0�嚔�A�������4�2���.7J'өP,�ݢc�M^��L�5�k�k�B�tn5PU����ξkh�!`����Z�[��3o5��ӑ�
�;*.��e�є���Z�fܲ�CIS=t����宋;������=ݥ�.�T��cq������7����R����zzr��0WNZ�;�D����#�{�(�m����()TK��-mmV��T��XsL�L�Ve��YU��9��eUS*��kee���e[Kh��Kh)Qee���EQ"#��Z��-)m��T[�IPU
���`�ckmR���Z�����k�J�TF��VU%-�B�Aj�R������ҍ�-��+�,̤�J1�cT�ڃTZUZ��4UFƖ�Z�\l�Y�.���2�:��%�PU&�h�m�Q����ʪ����X����U��Ym)meKjZ+jQV�C���]&m+�PS-t�LeDQ��efP�Զ�-ne�*(��[���E-�)j�*#n30F�]"¢�+T��k��[.]8��f8�Uehƥ��-���'�NTe+YǵQB���)X$oN{Gjm5��/9�F7RT$��#.���+ܒ�����[�4���xC+�8���=��%@�z�*�����醞�9Laά1�2Wl�N}�QH)���6ʐz�������B�PR=f�~p���μ9箷�秨
)��;a�����3Va�4��$+y�ᜲT����C�T��Y8�rNx�L:aY�';�Dv�S��b�ANY������OV�<w��ǀؘ |6E9�6��H)�j����N'�14��bv�A��X�y�9a�AC�(���6LI�Qa�*o�'\^0�S�9����y�;��́�XT7�&=�+6�Y���u�h!姈�B�ua�R
~S�N�I�Tyߺ!��&8�� �G��Q�r|*<m�DB��{� P+=T�ެ��',��si1 �sř�<d���WI ���4���3���I�d�����Hpaa�
���c8ߙ&��%q5֯>�[�x����}�潎QH)�M��l���XqaڡYƬ��Y�k�p8@Q`k���<a��r���\��i ��8��3�J��7q�W��M{���plB}ڊ_(�Q�{�ׇ�U�,6³��x�Ϛ¤��;k"���6��HV��|Ä��]�ӄq�&&�z�I��@��>���w��m
��~�����,<CL��&!ϔ1aS~�s���AaP��բ�Xx§��Y�tj�H
.�*)�Hq�����g�7� ���o^��w�=�;���:��a�i'$�.��
t�㏨V
A�z�a��bNP���+|�p��Ɍ��J)1 ��Kl�v���$�o2x�PR�L}�}er��8? &@c����P5�@��a�
���g'C�%|La���&�P<��!��ڡ^g�$WA�4���1�B>��π����Q+�/��C��U�0�� ��gSb�(V��g;{�X�g��Px�4?=K���N�6{*����v'���j)..Lě��k���U�ثf�21s=�^�VT�ZI�ܱ������ =�NX����m �Xb|8��H(q�&3�J��j����9� �l��p��L<aY�p����Xqi���U ��4z���8�5�!Xij�߾��tU��n���`xD >�����,Jöb��k,Y���09�ěB��l��E�M����� ��k�5�(����c�Xv��1�~j2>��E�6u�C���p{G)�B��;�Y��Lg	9q'[�H��Mo8`�R]sd�p�{��9��b���eb��ɴ�|�:�5Pڙۼ�������T���>� gvxɌ;��H,��f2�T:��<@��&'(�a�4¼�{�4�Y�%x�ɽQH)�ë&�O���{�r�߷��xuO��f���AH.���1E�bm���O|��1��V�H)��I�����vb(r��>0�8O}�ު�����}h��l����޷'>�=f�t4����%M V�y���!P�u}g��AH����1yߙ���0�bw��;2ŋ;OXc&2��
�{d���Q֦�e��W�� D��h�󬆷E�霝SI�u�N�4���<d����� �@��a�r�^%� Vz�CG~�SH���<�:��ֹ��7�n.0X,�ꁴ��a��
��Y�Ť�N�d�m�!ͤ,�&'}Y�$���%@��`���� NC t '�������P������9a�
���R�t�[����QH.�􁡓�T�t��a�š�����=f���恉�<a�8:�ă�S�ݜ0�Ho�<��.t�|﮼�9ס�+<d��v���L�v$V�G]�
ö��N�H,�Y&�ԕU%B�h���T��!]n���8H(t��v�Ȅ���yoy�qφ��x������y6zĂ`�6I�8\*��q���ȹɣA�;�Gu��Y8(7��*`Z֠)�nt��۷W�{#�+e#G�ux��Ŗ��������{8X+b�2L��W������4�MG�l���p?l�AH=ӶśOcT�B�]�����AaXk�a{�bAf���9��XuƲH.�5�i�2T���
�z��'����yߛܚ�A�a�0��������Ǿ�6��
z�ua����_(La���_s����S^�RbAa��Y��)+&���m�N����h�w�����I�R�0��ć�!�o>ROrΐ�t�x��!����'�5��G� q$���2v�T���e�kɶViHo3)�t��P1 ��W܆�z p{LCi+=d�u�1�W�ǝY��Y���p�a�97M3�M� �����d���/�Yƛ���;���='I�I�ظ�{�6�
��
T
�ä�:=�Ă�`��H);�$�Y�x��
��+5�;݇	��QM��ȉf�k7��~Ȉ L{��8��pkX=d���O+���R�1&0�7���C*L�9�M�R
x2m�[@�*<>�E�_��m'��g�l�@ʙ⤩��;eOQIXh�̆����Xm�H*�Y�J�*r�S�;5CI9d�uu�!Xc��d���]��	��/��yE2p�ɳ�1*;M{t�m!�S]ٵCI����m�C<eH)�c���D�Ş"�z°��(r���5M$8I]�\s��^N5�^o~���Ԃ���I��
Ç��i�2y��g,�=d��<�1*C;���A�&��L=g��<��Y������4wE�H,��k�w���7+���<�zܹd�Y�r�f�AI���Ԝ$s�����1��1��{�P冒�qݓL咤�t1��S4yt���S[� �,��S�����ޥ���2cK=�ͻ{(V�K�}�w�q�dئ�9Մ�)�pQ�uq4���3fd�fG��uy��vF�ב�F�o�¯5Ϝk&�c�d3v�4��O���@�ָ��}���~�Af��z����æN�`�S��g4�0�oPĂ���a�z�*�s�&�S�RVpY1 �f��a�
��tĂ�+�o�5�u�Ʒ�;�~q�<E;@���w�� �C[��i
�hrwt�N
h��&��7�Pĕ:@�'\o&�t�m�z�T���Vz͡�9eE ���u��w}3޵��w�[߽��
A�ߚ��8a�
�N옇�+;g�P��8�������&���p�0�8d�)9�gl�=I^9�R
v�S�M��{��u�M;�z׼���&2o�1 �L;O5@QH)�\d;g	�L/�JŞ'Lߴ� ��W^R�d��*,*s�{��L/�Y8���T���������}��߷���t�P�41�Ot�Hyl�|�+0�S�
�Y�m�$�TY<<�l�q�É���&3�|�Ăé�)��RT��o�Z�<�x���ӦLeOQI]��ă͜ud�T�sC;I�n�S�
�w�$�*G�B��6�yd�1��Y�<�{Z�� �� @�L�*ˁXEok'w�}�|�ŝ$��9�Ն�
���Y�<C�*)=gG�8H(%�Xc�W���%g��b�'A�<� c�՞�k=��1X�g�����1��9H��*c
��<@ߺ�5 �N5@�Y�c5a��a�{�H
)M�a�bAf2_,��=O�@��'�/�:����߅ǫgިE��0�w�R,+�(u�0��`zְ+=d��Qy`T�;�&�[&�}�+0�ֈ)<T���iQa�q��7�5�w称�4�ˌoTă��̰��$z��IRz�M�����=¤�nyE�L<aP��&$x�eE=d��'� �<��η��U��z�\���iB���r���he\��r�v���K���x~GH&Q�,�+��:c�dL<s�;��JSS��STiMt���˽����+v]�ޚ�X����=�m�u������	�?N���8Ld���ed����8�0���Q5�f����
��Ăͳ���b)+���$��rÖ��;�W�����/<{���[�RWv�d�
(k�Lt�������Mf�N0�+1�yO|�c+%M�G�iU ��4�`zԆ��WD+Y��q=�$�Ag	�|+�]]�����}��S�%La�1 ��8�V,��m��
N���^�1x9��L*ot{`V��E<I�+
��ݘ���Ě<�@Q��L��<j�h��*���<*f�ye!Xp��� �2u�:IӉ<J�9Փ�O\aͰRx�ov�^e�bVz�+5͆"ɶT�)��$�OY{�;�o��ߝ��}٦La��R+��� (�a�Ϲ8J�R:�+%��T�wgL4���cMXc:d���>�H)��&�RVpud��'�y�q���\�4k=���͂�Y�<M&�R�/��	\���0���$+=�g�E:E%q�ĕ�2k=�4�a�
�2y�����Tߏ{���׼�|��d�U ���ua�ځ�^�
�l�3��R,�YS��yCL=f q�`�,���<§,8H(q�1��ɉ85LE��T߶K�7��|�m���/���7"L}���������JG+e@��3a�=��=��+�pi�r%0�o+�O�M�e�4�c�A���X������ND�+���(j5��L�vT.��Tx�W�����@\�C�{���=�D.{�;#�E�IC��;�m�+�	Gle�Z��1|�mn�1��;k��U�Ϙ1Ig�*q�m��z�r��YXg��q��*Wģ6��{���e��%g�x  ��7�jvczz:�|�t'���HG�g�wEj΁�X���R��f��R*�9��d/ب�7�a)�o�J�v%�Y�q��NTT�����;^�^� �Wo�^�h����sW�͟q�e�԰�+��=�_!ơo.��?m��7w���{d�6�4,�EN>�F�XW)Ɋ�v� g�*�#���;wWwd+��pc���N��
lf(��5O���lUu1�۱��л[�[푰��~O�Ѧ0!��K�\��: SϹTL!1���T�/2���+g�� Q��� p�69�Ź��;�,���B�\�BEEE� �Z���4.m@m4S���N���� �\�]�=Qp.m���Z��r��RʛC� ����J��|�54y2���8i��]�Wܕ�љt+��wC�;`��p�d�	��kt�R��1��ʈ��2s�Y"gKZ�L���ۏ��[�(��ǘ�����4�"|����}�=�{Ӗ���+���=|�dʡy��Y��땅^���p�!+��S�Y��(瞅�#)^���+ϖ�r��(QA^!N��]�y����nHs���,�
Aųk�*c|�J!o/X�&odR\.(�>�꼌D����d�6E5� �ٳS��J����V,�p4�ii�:��7�y~fC3�b����͠A�j|���x}!^���{Ņ;d*ʳ6�Ӯ|�׈R\����@���{�qm]��JJ�:�-8}'(s�WL]��B�#Ors*v�C��ݝd���1sD@ޜ�$9h��aq�O��6����=m�}3�m�J����揕�8��H���9	�H�Q+Ll��>�.��m�����P�n��]�64���,]1�:��
������NF�q�7�g.o^d��_\\)��xWt��ց�E���ɼ;r��.+q<
t6b�e�W�U�C�8�6]HR�3�S*�e�x�ѧ��[��od�ո�;#Ȓ���� ̬�QlD\��m�K􃧁�C�v� �(bv<ؗOl\6��7X�<���ju������hB��Έ1�4^zȕ�R���ͱ�>�w���(b�ؼ��V��r8�1��	���!(6|�#X�a�&��܁��"s��"6=�r��u,l[�š�01�tj�VFu�n;m.Lo�PJ�zS�w ��E����2$�ET
��[܈�҆�`Yzm�A�[�BCTC�\K� P�NtA�
���/y�1��f���Y/��C,7&��5gL	^�<�0Vܾi���c�Nxu�>�v/԰����i���"������`�(�Sp�(����b��'��t7#���#�VN"h���:��ū��B�]��-�����g9L�s���5f_J�7Lѿ@��;G��Et�Ef�=���I�o8��@I����$�D^�\b��{&'fJպ��)��̽�Mٕ��X��_F+����'Ti�UШr����� +-���A
���Բ�&�-�=t���ȗ�7��t�|�ͯ(��/oIZ���,���$^��4�����	�zqum�o�jlK�;>��np�t>��Q:X>���<t��S�Ȓ�p'.%H�gE7bªb-HpŉXu��
yB�j�tB��+r8�"�*�pU
�w�dR�2���!�X�~/CJ�r.o{:6���b�O�r��]f�/�b'���2�:���˦k�DffgYr+B�rt�%n���d�{��tb'=kJ�Ec��f8�ܓ�1�#¹��UKH��R}_r�:�C��oN�۳��8�`\P������a���q�?3����b���[�n��>}�PW�{W:��*��Ns������*����N y�U��y ���,2��*�]�(_(���k�vT/}==����J�#ii���mL��$�T�Jww�])�,c��(��[�P�9d���cK�Dw���ֽ���_Y"*�W�  =.�6�*
/$���'`�}�c�V�>�0f����b�����oEM�gM�v�)щXn)�;.ݫ����uޙ�)�嶭֓�r8����J��6
#�Ԧ������u�c�b��u��M���f�6�
��cy�\����\�F�tzb%=Sho��6f ����$u�1�F.���*�1� Yc��~j߸N4��{�Wo��}=Y�X����¡�i	.�]�G 7�#i˺����o��`�NX殖��;�{�y�+��:<����e]�<i�V��5���3&͙9T�ܩ�����8�-���k]Ȼs����Џ&@ڻB}����7���F.]�%���{-^���/u�h�â�CU/@H�~�
���Z�"4%�~�]���.(@��ĉ��ʺ�nU�k.�XW[2"%G�v�S���/R��׸oJ�q���u��F����{I��u�w�:�,���n({�Od���*�\5%x�Y6P��aX���r���8��
�)Ъ	m�|�Ö�5���n��w�G=�ӈ�g .�kݴB�AZ��m��
�X[\�MD���{�� RC��]YIV�Ʃ�i`��S�зj�*�p���t���T�+ũ��(�Ĺ���W|��U$���Ƶ�J��C��i�c���;�ނ�eamn���.����ޫ�����=��94�jQXBZh�)�5��-�������!\N_^�b���h[F��/B�Í�����MݩL����mt!�O+$n�W�B�����v�[�V2�q�����6Ӓ�͉fc�ee͟>�v�+U%��:ں���SLٮ��#����yj���������W�L4fn�P�u�K��(5-�U�.!��W5f3��]I=ƍ������emu'@��N���srĨ�gӲ��R�w*�$*�6 ���l�!qJ�ۮi�"���:��&&���wG��3���xub�338q���A��jΔbQ`Y5�A��ԉ��U��� ��ɒ����Fg%s�^�����Ԃl��t��e������Q�^hM���9�e\uap��n�w;���Q(��t�zP"N��0�v
����P��+���v���	��Ӄ�
"�Pz��ŧ�ø0�,�'`���,tZ��`s�j����iu�f�_
�@T�/���[�q�P�v;�(#ϸ�1�Vu�Gq���J�� /�Z�ړ-�No]Ɖԅ�N$\pb빧q���eN�n� �]Py3)�g�1]�Z�]\���e为>]C���gd���ʺH��y("R��]!��]�p�ooO+��,3��QBm��{E�E�~ԑ��U�f��K�b����t��o�sT���.
1�mS��f��:�.ٴj��M����]*p����\U4�X5�i���u��5mm��:ĝ�>�]ǹ]R�f���#Ux:]Z�s/]�3��`��I�\iQ�*f2��*ʷZ)m`�-A�-�̨�Qơ�Yl���B���Kb":e\�L�
&Yr�ˆ[��b*8�5���.eTp���)��Eh�R��bQT]Z2نL���Qq�*��q���q�T*�eQ�U\n7*�jR���,TA���DPը�c��e[�P]Z�T�f��b�2�dG\)Z5(���q�ELQ����H�kY��,�S)MR����5sY����
�"�%��Q,�c���Q�]!\J1QF-[A̸$�K+
��j\��aLe4�0J"�*�\���VJ�EL�i[`�b�(X���ڬVU�LxGM�aM<�n{UG�ۂ	%W���h���m�or�>�W�y��諸U ��_����3��E��DW�!7�yNdq��/"�@J%Es�`)�;nI�ѹ[j�ǒp��:M���Ȋ��c�L[���y{��9ݭjn{+��Pq[6��N}aO�NT�P[B��>�>ŝ�=�rDl^ol���TQ�O��X}%�4`�[ ܄���T�� ჸq�ڿML�.[�=�%.hSXo������+��[�7֨�|��0������u��̡,��J�w�����ws�pw_v�����,#���¡H"��kƅKW[V)<>4�p��<�1׀)m<��S^��8>5������џ!L\7��+,�qD#յ�����6:����_��������,c6��6��)�ə풕,�1yN?��}�W�����^v7��).[
��/O���]w㞤��=�C+�k�8���	W��k�B桘����!lJII�^���xK���++{Ys���H��x���u���q{�%6F��FX�z.���T	7](>��W�xxz��֛V6�|&Cۚ� �ϲ���:��R/$�Qg�m�̞ݤζ�l��~��A�2�4�fF�:b��/ڮ#c��I�f�r"�ta%%];!��c�M��F��m�'�͞a�D��'KٻMn�FQ\���bA�2�a*�̍#	8n�Hꑈ����h�^����aOv+C���z1�s�_�1���X!5nlg���6�K�{��'�L�p9�!d�؁垾<]���T�]�)G\+���ݬ�؈�U쇆�ļbp�c�� d4t�3�S$����]f�<���,�t!����*#��-��_U����kEK��>�M���I�
5�Yhe�d2�Lj�t7��<P���,R].���@�m3V��>��8�ɀ]tIɶaj�d��sq�Fn��DR�����ƞ�O	#�Fȷ`�^)wjR�K^+��I��Yê)
�*���9LWX��R�ޜ�+b.^�ɺN�G�7�rc���9Ֆhڻ�ۛ�i��|�< ��iil��d��w�Wo�Aʋ��)Xk�tA~ۣ�� 
zd�)�
�$5*��Xj���t��DP��bB�]��d�*���͜GG7d8������@1Jo�*}n�nE��ehɛ������	�	� �hk�g#ݹ^1L�ۑ�i���=���	-�ҍ�V�<G6F�@�7����lL'��ʃa׶N��ky���s�kH�ۓKԖ��p�|TẨ�Kq[A�m��|�#P�v
N�������p�O�%�������0}��X�&#��af���Y.{ʀ�xȱR5M�}��5<��^�QS�����{�������J'�G!d5�dρ��9(�~<ᅐiA�U/j���	��,���q�-��a'�@"p�����5���Θ�E�˹T�����3PW�9]�<�.7�`:��uֻZ���BP��{��z������a$M�U�A�n9���9���嫺�R����#0� _9�~+諭���<M��2cjuH�'��>7�V��CN��҄|��^�{�|?_�^��{��>�k�
��"j!��Ga��N)���nFD���U,O[��C �k�C!A���_|�U�
�Y�pv:�P��)�:W���Y��H�#�U�լ1k
�`�8>�	��º��gA-"��LgXq`�C)FGA3������Sc��c,n���w�Z�\V�+Wy����n�.W�~���7��2�T㕍/N���3,�����(u�A�I����ToW��`.ݍ4ɻ��O{#�jfx�;]K�G��)B������4�ʄ-��y2�����4	|F.�b�Y))�f"@�C��,;��1QJ���Ϋ�%ϑZ�jX�؄�z�Pgw���p�Tr�v1c�1����&�_(�CN,���2��4�N��O�kv�mi�qQ�V����8,�C�eЌ���i;.��ΥN^�|��ɕ��ޝ;iq]1'<�Nz��_��xxxT��M7B�jFG�Ջ'e���ٟu�ۜ5X.�1AzB��u�n'��.�-%��ߗ.>~<x�OMʑ
��~�A��NX���Y�j��|��?1^��2`��k��LIy,k[���>���ü�����g\� M�G��!EJ� ��ŠZ�yq�S��{��es���št� ��0�)�8�^ȸ�S��6�	
�h�Tb	$��u�Ș� _[�C��D�q" Z'�)8�2�X�r�ؽOx�D���d���jX�k�O�>��T�P[B�Pڝ�3���ƽ:l"���i���m�5�=k��y�kn��yZ {��VD��-���2_LG�q���ԊcMZ�ױ��B8!;�������Yhq�I>���4?
�ܨBgd�Ls�bP�Q����	KӟU�n�c��Kb`�imF@�t��Z� ��p��;�N�d�Ag8r�4mob\�k�Y���Y1��G%m8�s�Y�v�Z&Wb�MI�d����Ca+�S��{����u��=��Aa�����Y��F���*��0i	��8P\7W�랓;�Y���=.�01
1S� �ٳS�>a.�J���kEJ���fؽ�������1��ش�a~5���)�JU��w5��*�1�y]���j��������%�aP����&��$YM_��X�"�
�Op��#NP^�������`nbE�8'[Yݦ��3���C	�L��-J�Z�>?�����R��$\��vQ�3)�8���:�͠�4��B@�H�VVq��ӹ�.N]?.C5K����64�$�C/͘իp =�'��%������ؑ=�v�0x�,�9G�g���ӓ�ҊԱ�-�o���0��=]�N��N�s�H�e��1�4�Y"�ή���W ����#�sE��}���#��bz�-w�E���r�W�PW:�Xn��T'gH�{=Fƺih.21V�2�3u��n2f��M%����r
�J���V��ɳ�n>��UW�+���oLJ|�����J�����+(T����r�Hi��*RE��*#cҏ�w�(u�Z������=�C}��Nx\�!g8J�������)�;�h�� X�p�N\�B��{�HP���­?1��<���uj�:�#ct:��˄i�i��2q͍�"k���; �����Jå���U��/&CW�[��P�O�P�tg|�Q��6�� ��j�8����
���7���P��C(�)C�
�ً��B�B����rH�p���K�Q�2e��Ӡ�2DtY�^�^�=�T ��n|�A�,�^���+�廨�
A$o,k�ĈOU���J���>V.�)Nz]�sb�q~F�N�ğ�tFC{��o�犜�z��t�u�Bg-������":&<�=�����^=ODF޵���7K�vZnǝt���Z���f7:WJ�/�����-Y�ܤ��KM��|x���i�]���nQ]wIW}�x 0M�M7nG�*uAo��Ϝ�s��"��Ul.���\,����~��1�`\�y�\�s5�H������dG;S������+���2��'u@r:9!�~F���*z5	wV�i-aq�Ã�����0�=�.1N����Nx�thv�b�,1r:u�e�S1Mp�b `~V�!	A�����L���r���n��/B"H�cn�DK�����{m�Xa
UKHF5P��}�h��ى���ˋ���Yhp����{W�q�8ɑH�7J�STp�[Ga��n"�+�<��6��ȋ����iM#B
��J`�DC�[�k���QβW�^I����p��dߵ��P��N�o��r;���'ǋnM(h* �f���ץ:1+Mǩ�yY���B�8hW@��zc� ��*�Q/���Y8��V*խW�Y*[���B�ٍ�v���,3}�G@��G��Y5�s9�z��nB�5���H�\�g��Ɠ��lC��9h��m���3�ط�x =��xW4��l���Ffԁ�OB�4΃hq������L6������w=�-lIǡߪ�w�g��Xaz�z���4�CX��11�����%�bOy���4=�*�P�9����)�c1�C�;th��.#�Ww}�/���@;QhqbWb��B�,sb(*�l�|�}\@�U�,+�(e��CEK�qP��1�s�����j�����d��vǠp�yt���EW����A�o�pC��^��B*e�n��Vz5��?+FS�@����]R���E��2�$;����=6��Y�d#K���i��$u;B&�3.R�97Z��g	�IE��[ 7��G�/��F�i���(�z��ع��U嵼T�,f[3�5@k�.够H�d�3JN)��nH�c^V�ڵ��F���#ͥ�ڻ�ʬ�1Ӛ-�2(�.�}���m�T6��M�&E[��Z�,��k��,��;37f&��sSɣ�.����Z�H���ݞ��W�xxxzn��M����u���^�AF�9`�	ϐR�ߑ�e� �<@g�u��l�u�1P.�u�j4*:����1jK��B�"n�&*�6���iw[z�0Ԙو�/��4VgU���=ϡ��h����6��N�do
q�A�i;��ѡ�T���gc&�V��ːf"']^��+���#L�F�j0�
Ah��8�"�l	P���E�q��5�xG� �i�~[e�\pǱ
1]��vl���oO���P)NnN��c���Ξ���y�{�7/0�F���4�̍N�s�sJ�Ѓ�yڣ���m[��>�߫���~�%�}�+ja�7G{�;\&�ͅ �$7J�$Bt�9^^��s�P.�.l�SLk�Ϫ/G�p�}t����;�H�i��H�]��.:b��@��Ժ���aZ��K�&y�h�k�^i��w�	��h��Z`
����}Clx�X�16e��:.oJ��[׵+m�.S,�TN�<�D����Xo//�����N�m��K��r��g쏺�בܕ_wSWݍuX��t"ݭ�)�[�.���-W��MT��B�Y|0R��5d�QCuz�r�PUݜ�[O x�LME��wt��b�Q#dtf�'Q���}u�gvjq�a���!��PZU�.�jW1��k;R��53w��'�oUF04K�3�c�5�X�+���8l+8�픅T�^V��}�NK&�L�e-`���kyK@��kW���VV��ӎ�eT��畷�;[�P���F'K��=��U������	q�s��)�f��It�<�+Q%V�������j{g�&��	�T\ξ�+1˷ ��G��:�;�U��De��ܝ��/�b4f�s���{X�rk�ƂWP��̨���s�ս��R��OHBӡ6���nE��Aug:�o/Z�cv�F2�R��p���Bz��j���C1,(�ŗ.�詐�C��s·z��W��/��Q��7�;h˶���䖰%���sEq�[5�Qo�@��P�<n��
�m���R�)�ᛑ�XC�{̃t޲򭙥[���Ekӆ���.m��.����}���̡y"�V�֝k;`t��@)J]�eA��((��h�ˡ�j)���ʻ�W�R�89	y(P��4%���Xn)a�q�A�Hw!�n�v�j'n�ҳ��������'a�ܳs[�&�Fv^��؈l�S9gJ����;n�6r��#�]�� ���	d@ѽKv�m�*�a�P]��8��m9�p>��r�ej�Ö��vyپz��C���U�Z���
�2vU�YVn��2��%����W��^qoR���H��/�c1Ē ��ś��Θ��N��oN�Rt��ҭ�H抳19�mL��i�Ğv�:^�+h3�HD��.J�-Zt.T���Fv�K��@$�	��K�����144T5K�10,m��Z�R"���2�QX��*[Y�EU��,�cU��mQؔdm�EAFE��U\eQV�k*���EQ&�mA`��& ��(�i+5K)��-j(���H�Ŋ�AAKlm��@Tb ւV�"(��%���]\f
(�DKbʊ��QEUA� �-B�eT�QaR�j�K-X�U�岶5���K�PS-�ł�T��ʣiX�,F"1EAh�AEEE1�֨�*��VұU@*Q��"��H�,TDAVҕ* �P������QUQ`����UV#(�[lUX"1+Q�Q�ێD$�Bc&̉ux�%�����/0'�a�,�K���ws�z�l@��9к*��T �=bq�m�>?�I�O��\}���׌�$iq�y�+!];�'��uC�Ҵ���;�z��$4��"p�!�:��sN���qF޲��1Yy�{"���P�b p�#!�c�������y�����a��C��G1�L_0�*�2�LML���u������$�^���T�F���X�'���"���Y�s�7)*]<�%����#r����[�S�L�0*X�X��h7)U�����t���1o�O2%*�6�<!����)�;�ih"<��r�\��h�`*o&=����W[��������!�d��J�D�wWݯP�Th'�U/���0�U�^�g���m
� �iz��Ci����i܀\�{����)���<��l
8FU��&�{	�*�+�8b~䍗���^�����b]Y���m���S���طk��Nk�Jc�^2�lF�E����U	f�m�i�V'�>Q���$�+�����P�SS����ξ���,���ޑ/&J6�*1��4����^��7��OlaHK5�codb��X`Ё D8@�CtY�+�Ŀa�B��mmi�*�湦��E�:�&�L'#(0)	
�����P�1
�fj�Z��L�Gtf6��]ϵ��7T�FiKr�X��`#c����3T|��g���9��i�~��^��	Y��B}���0��0��aw�<�3����j
ug�5hW(}�5.�<!i�Us��{VSO=�9����#UǗ
v`Σ�� H��"�1�>O�ʓ�i/8c2���
K�_������Ɩt�9q�ytu�����.)�Ϸ1{��`�40p�h�P3���@�Gv�`�z�zS=�J���2&�x\�,��
x��喋�dń$R�\D���� ���/�kyɢ�w�K(�f���Xkz�؝vj
ѕ�>5&1AF7�r2�1e]����x���b���$�q�P	��[����W_=�X�OE\/�TԾ�<�2r��~Nz��~�����Daz��f�2��q�>�Ȯ�ܞ�r��R��Oٷ��n�B:<�`H֬�4� ����]-[Z���r�3�ސ�a��^�vxU%*N�2J�fiOf�$Ӱ�[E�=�#���	�D#�Q��N�	\n��������."cy��yU}�RC�e-"F�䣐�;�i�v<%1�$r��,a���ح��䗻�hw�g����A}K�`���Ѩ����ֻ~gb�{�M�V�����4]��l�fd�m*�S>��螿n��X����j?�*+�}fq��C L"�؊U&a�7�b]�%�U�z�^��v:y��ő��b��=�jj��qGtf�^��Y��L??H��,�?p��<,K0c:�b�|P���}���w �M'����6[cY"����2j����d��y-уf�qZ�N���n�[����rI��������p�4њ2[6ȹ�*'����e+8�[�YW�}�	{RY��zmw�\	4b����0?Y2���0�s��WZ��ɳ�AB��:A^Q�:�x��6ƴ��´�z:���ŚV�ZD�^pH�\���lk��*p_S�B�労�d�L��>^+�]�IگK��'q�5@��\5���8m�A��x�fL�u�Z8�6�����Ւ�r�@'>�-J��;�[D��N^��D��"K��2�ɗ�U.>�Ν��.� >�|j	��1i���zC�B�o��W>�3�#̱�%,e6*߷�чT�fuS����+�q�7HE'�q��;������U.�";%zc��4if�P]!oWo

W	��͑�3]Q�@R�.���'h8��Cj��t��n��'LVx��ϴK�<)�k�r�4,٦)������U,VDɛwL�Od��"]��S0�&��m8�^M�g���T��u	O���͵ �ћ�tb<.s�g;����Qܟj�� )ۉ���PNH�^���q_x�i����>�'`�������g����S��2,�W��ϣ��q��տ�K�1r>�?��P5�N=V�Ł�*
�չ��C������
^��34��3wI�U��G��^X����!e�CNI���i��U��t#����"�W��8�7NfߐC�C-@h6�1ˎ� 8�2�[3]�1�Ր��'�`�`a�#��/ڼ�<-�T���u�oC�"Gj���,C�K���64���,]1���X����7/sb��� S����BQ�݌*����ǁ�C�{�x�k�LOZ��1v#���=����,[��C�y�H�1���.�#7"ԼT��;ܬ}�M����B�x��u�?7�O�Cg�]g�t�>���u�K��E����a
�$n/i���J]����^�l�]k��32�m!�kp�*�'�ue��m���z��.Ф���f�Y���[BY�H��$� ��]��*N�!��5��]��/q٣���+�������m�ٶ��o��R�<<�c)�����d���7)V����U/:�܅q�f����^P#�Q�cԇtdIv��§&b��LT�ծDL�W]�~m��ہY ��>�nog�ٿH�W�aF���W�\d�ӵw�'P�~��#�Kw��� ���Q�����lT;c��������H�u��0��3a*"c��#�Hv��HTj�x�ꏗc�S�Z7^Cq����B�
���d429١+�Y^1=F�L�|��Jr�@Q�Ʒ&�V{P�8F�6t:���ױ��2QYt��Oo^�qI�,���L[�PG5�q=V;��P�Dd���4Ҭ��YU�EϔI�1�?]�ӊ}����@�A�Q�LB��{J3�n�H����ܗˌA����;�cB�C���q�]3s�̾�uKٓ�(�v�K�RO��P���[Zqq�Dw��ɏ.<���S�������Nh���,Y���n�1;TAdO&�h��V'�e3����*r����mB��l��������wa�����c���7W%�`U
%]�7�e8󮊚EޒZ��������W���-9Y-�,>Aˌ�]�Ψ�s�ˆ�*�ĳ&"r@�iwmj;����Y���j�ʝOT�ۮ6,4��llřȘ�ƲU�)�c���Z5��"�
�R�%���L�����cO�g�;9���_��C�г���^+.<\���s�mh�X����<�M)u*:�߷$(����f���X�4������f�o��k&L{��#-mC�9�O0*��2s�_�*�1��q���K2�϶3`��R�Ȉ�F��7����'Tѱڏ4oL8JE��p0%Nf܁�OY�P�5�,�{�e�6x���g�3+�D �z�c�Ū75�YW��ר�Z��Chӡ�>&b�̛��xey�(�⳥�DMw�9@�m�iR����I�X`��Fi[Z���yÇ(˜��"�%bPf���E�,���|��Z����cq�%�Q+}�tO\��xN�D�}�ٛ��|��Z�=a[�΍,���(��śx�Rm��+�U�G�e/�qݨ�I+�?[u<kҦ��t�V5�Ӡs�cm�t[L�Yr���J7C<f��p΍FB$<X����VL��'Jo�e��L_�	 ��&e�=ٴ��Ū�shY�3�Ba)�#�9�$)�إ9��g-6��fO=���s+=
j�Lꃱ�&d=̬��J��vB�(<v�
|:P��-�1�ٕ݉�)�o�8.�����F�Oi�� ��5lߙ�E=�t���·ޭ��
Y�O�g�f|���X������ٸUZ����W�w�U��K5�3%����`�p�=�Q]ND�S<�gWK�� X���G�2)�N=s	���0��a[R�v56��K[l�y2T��~�Fܥ��k��d�.�'\9T�+�����V���c�^�y�J
�,��y}��.?�"3=�F&r�\ѻ��QD�8c����y`�0lgp썗4=��v	���U�~ɑZ��[+�=��q��GP�!�u�y�x�bK���dY=:�V����71�p����E�q�)D�a�
��\jٯ�d��pϾy_rz���Ŷ�1��/!D�� ��q�[�Q�Xm	�7}-�INMy��Vۇ�/�ODT.��).8gSD��ƕ:�[�V���p28�Pcuk�d[_;�M��jh���~��$��g���rI�3-o8;�:+��ˏjٷu���t�r��t�ͤ���M@^�Uw��JO�lFq*Ti�<�V�j���wvI.!������Vb�.n�ަ����>o�׀�gu����$ck�sa����p:�4.��;5rf*��8���1YR�Z!��b���r%��S�&r5��5>��r:��t��%�>ёkZgy�w���x�F��`�=��A�;����s�RA���sD�5�W�r�x�)Z0ufvyKŬ۴�w�|B���/�i��Q���7�����R��q�J�U�J���b����:�ߊ��1<->��o�6�Id�~bn��F��'�Z�����h����i�۷׽o:&�;x�bE(=bF�L�b���i�4��m�E�Z�XQFm�s�]�F9�Ж�I��}և����s�g了���	s{H�.B�`pƷ��qw�:Uڸk_g&�M�6�wh �x��E�ۥ� ѥ/2�ʺ��J��;�ꪝF�W]�on�s�Zn�ڸ8���b��̮<#�a܈r�SEh�V|-��2\`�`�j,�ؾ�Q�Hp}G��|��;���+�6Ev�uzQ%_qJ���P*Z�{���U6gM����]�����X��;��Gwo�+\� `}���0�,b*!��\��{1w��N�e��]'m�ƨwX��[�Nd���Ԛ�0������p��r�V4��-PU�/���*��6��x�/EÙ�[)��g�]Nf�e���]r{��h�5���ݓDĺ�
3RYւ��u�/���R�b�4�Wb�Kn�ڕ�^�q� G#ǥ1yx)�A�uęu�߮%�άlL�K�͂GU��	ʓEЭd����F��:�%_V6:�v���u���L{}5[���(�&ȡQb�liX�y��Ѱ�霭�QmE�����,*�7MT����U��esv�i�N|o:��7#����\[�����5���W�b綦�P!<d�Y�9J�]�x�.�����e_T�0Eb�L�٘hrfE��X�vT�#�ti��u�Ov�D;�n������xô�"�{�%��Zt��4�2�Sܡ��,�}N-H�"/5v�aqu���<�]�l��z'$5�d��c�茝��I��M�+�N�.�w��8ܢ3dĈ �N�"LC���o�n�ea;��C]�K��U:�w�x��\v�w��W�au�q*�2��:��("
u"V��lq�3NJǳ3rck��ⰧM-�!D��y׀�^̩��ѝ����(b�mb`��
5�ATL�y���'0�A��Tz�Ƕu������3�R�bWBOe6��Tk���e��p��<�T{Z�9KmP7�I��7��,|�Nkz�v���*�B���*Vt���X��TXQ�we����s;͋Kxw=�xox�V4���(�W�@�d/)b�0��� #�@eY���������w7hd��d65/C�h[Uᜏó�Ո�	iEb�#jQT�b-���-��leT�����("�DJ�X��#iQUQF���*	l��TEcҵim
��AV"�*�QAb-�ڵ*�=Ҋ9Km%,�R�
�b�Ŗ؊*�T��l�cKX��*�X#h�X�QdV*�+-����+B���UKhZQ��
�-iUX���Dm�TU-��PY(2�"���J(�R�ERc.YPT��F"����*4j������+D�ҭ��
�F�il��c[mUE-��ڍ�"1mP�#Fб��m��kD���ib�Z����]q�\��]o����)].��l���s&�M���,��\��݊����- 򝝓;�W�|g1�M1����ж��K!��	�g��k/��=1�"����z�L~8��*V�a���wb3f�CpnV���"�dõԐ�]a�v2P���$֨�B���w��69�n��
���wu���
X��ٮF�vνe)�������b�2�XI>��y9����#4=n(�8n_(����Q%t4�=�?}��I�u�n��)a�͍i�g6T�۬��yL�JF��J�DN�U�31�Ӕ%I�!�ɋI&�Ue��ll�Ym��Nm��F��86�³y�b��9ίY[��F�5=7�`2�*�m�&bJ���S�bsz�a����":Kcm[�7��=��C��&�n�|�4�+��DA�/8�Ύ��OG���m���)�$��b�7��feOx�+� 2�6�5�eA~d;��ʭ�f�m����sg�#=���ew]E�jKG�3���_*��]=�y0�.,Źv��\Ӈa�3w��W[�4�P����9o�~^������_:k�$�v ~B��h�x�t���^��7�}�h=������t��bk���V$��V�T�^dϼ�Fk�M�$�0��@^c��>�a�K͡)A�\T�V�&�u�5��щV93��z�U�)az��f�D�(�gt#��T��4�v�p��'�lX�$��.�i�Ҟ�^�K�(�:���gN�.`Cb�Q@Ғ/g:� z}��Ů�KOvr�����+�8�츙꫰^��CΡ,��3q=9�Δ-&�C���t[�A, #�91�l��"�;T$Up�%i����^���n*s�E���J_xz�+m�U3F�y�/Sˁ��*9���
�`�^�#��r�����W5���4��Ym�웁�/�_EE��<55te�����li���*�ٍB�DQisk#^:�|'���2��e�=�Gm�Y��h�\Z2�Z��7����/D_gfo��s�╆�&�;M;�]�XqG(��P�ojV@Y�����y�IV`c�ޮ�x��pm���]u)�mkk:Tnk9�6nr"�X����X{X��~S��!�	��G�[��}K���ҫn�EX�D���f��1�Е/���$#߄\�c9چZ�׳�nU���	���8�8m`Z�x"�����3YT���y�9��55��'����άnx������]Ҙզ��i,Y �ձe}i���օ����F��T�8$b;����+�������������g�`�/(hǹ�XEXA�n��҉�[��R)^Vۇ�gT��	����곍7'^����u�ӫM�I|ݝ��S��ZT�Q�4Y7����0xÒ�n�r"g_osl���f�"�d9����lU�+�&Γ�4�f�a&�X��YsM�c���^�T<�Oy5��{\9*x-�N�)4�SeN�����aa1 h�E z+�ݳ���le�j������y,P�5�:\��ķ�9P��u/s1�$c%�*̨B�4���n��d���X�{�+��q�y�uب�@��գI�����������_H����$ԍ=#bS���j���
0���Ҟ�� &��8eo'jE�3���������C�E�r��`L]ja����Ӵ�m`�*��[W�E�N��1Ԯ�ݨ�w����~�n�J��YmW�Usy���rQ��G]a����˙i���F�A�Oh2͍:�jA��)������Jt�F9Ж���g(g^��]J~Kk9RۯId#4R��9�D1�9�+)��W0K�R���R�i6���M.��ZO$�z9&�����9MS;��vew_�'�lE�L����3�vAUB�mX��u�\T<ZGQ˫��7���C3��RWX������&�*��+t)�)׭����=B9
%�nt!8a�D�Y��<��k,zH�[x
�;ˉ�X��gv:٠�خ�Ի����m`Ĕ��)Teɬ}�k1�*�3� U�u>���[\Ӽ�sWB�WR�kt���3��FB�+���J���4�`.��:�q��r�;D79-�ӌ'O��L���q&uz���O�u
�6K�z�7�3m�m��3}��}	l�sNf]��e
�lw'$#�1�mȞϬ�E���7�w8��^��[zЭL��Cw������oJKK�!�Z%��)��om���f�Ƿ>36�|�R�C(��\!a6<�j�*b6�����ܹ��:JnѠ���Z�p�v�;*e֥����kʜТp�i�uxlgO������<��M`�����7"���FT��z�W��j�T�*��U�z���C���O\���͵ͫAs�8����A�Us���E��Y����e	KaӀ'��y�_P4���2�C<�� ~[��_� m��+�rD���Ui���;op�"���ؗ�"��\���<X�p��<�;.k�u��P�}�����6��j/4������RUI�\iөX�'HҠ�n�Q�wI,�K��y,PIB���g�T~��żH�)9ĻS��6z�(+�ʝ�ĠH3�$@R�ޤ�ke۽�*
cR�)l�d60"��)�#g8��r*��%�R�\e���3<�
�n�4T,$N�W��Ǝ	���0M��B���[���7�wZ撬�v�0dn:V��5Dm:�l�S�	���o��&=�{/)�ڇ�H��	�yOu�m��^�0�E�_��8d�5��ʽ9J�*�� �WMl�yk������5�8�Y�qF�HNF�f��cn�C�mno������nb��M4�/q_58���N(=!HA�sJ���E�f[Mؚ �����m��^�n.�#Gԓ�vK�.�`�<\1�]c������_����}���roP�qIu-|�~5�}Dq>^�	C�'P��m��<�6n.?�9���j��'
M���Cۑ��:Dt��4��=�M|�ݖ[���nz�H��^|�}�n[㞶k�)����� u?���4y$5�$`�.:�[�Ή�`����\E\��;^��Ɩ]��S�3�OWr�ĞZ6"Qu���ôx[����N�6,RH%�%��7JJ��������'�}P�)b�Qa���-V�N�x�p���>"m,:��0y��ޔ_lh�����bsTNT�ֈ�,�J,�.��[ɟO4�����%�zP�^��U�{�l�w��o�2��{����*6h}�[����;GSV��s/3,�TW��qZ��<]R�U�	��p�*�4��� z��.䙑GùQ0拢Z��x��*�˄���'^�,EUq@�^:��	m
˿q���XK�ޑǾ�Y�:ϻ|p�7b���T�ẗ́m�!�Ľj�S��/�\����.���t:����8��V��,�r+�py�VS���д�j6`u+MeB����(�����e�
��� ��\�W,���]���Z-�,�]��B��#r�]`"����E8=	x8+��INV�;��ķv
1H0mKB��H�3��XZ�^I';8מ�Ig�R�}7F���f�����㽚��N���ÊR2�np8���J��n��[�Q;�wt}�$�Hzח����N/��85���Mf�0_U��pn����.;y*�˫G�#W\��!��=���yn�3��PMK]^��u �#.<���Oq4ڿg��O����`}CKb����]��j�����E�a����9"ڱ�����5������v2�FiA�BA{	
|��*e<�ȷ%BO+7Q~��U^�hBaf��2U��ܥ�$U�����o���ǴhLU/Sˁ��1ʘ�aº��=tz60�-^'z���_�R}�TO$z#4��-�S�;l��E��Ùx-7{(Pm����0�ڪW:HZ:�J�a`a��ٗ~�4������^���s���s2o��g��,r��T!ř��Ϗ����-������µmQ�/���1��&�r��5�fF��p�"�x`�6�-�I����bh׻� �:ǀV]
Ѣ춗t����"s��W6�ױ�G��.�xyS㶱fr�3�+ B�G�Ƭ;F6H�{-���� ���m\����&����n����mv)�h�����K�/��:�r�C&Q�8��)q�� ������R�)S����z��(.VL]��dmhJY���0#-hީo�p��y`G�Ȇ"!�֠���WA��cǾ���e�|���{�Dx�b�N�=�fd�zNZ�4�!V���O�d�Q�h&WT1��k��k;
�6�
�8b��)]M@I��KdpNX�ݺoq�[a��фR��:X�ۼa�<p�;�{j��Ս$����0S\2���t
.R�mڔ�,� (lg^˽�ϕ�sG���ײ���#����W`nE�Iε�si�v&�����*CG#vF�z$U��[k��1-q���*쬵��v�&w*>�v�B��k�(bȍ��; ?_Te�#�
��8��B�vЋ2�8I�����ںΈ-jQ=tx�t��"n���T����^����+�)���ݹ�!�'j�-V���td���%�5��4�qK��n_X&�U�pV�Y���۬�U��u��T<�8�*�e�̕�4�Fv*[;'Pɵ΢�7�Rx��J�o��)u&�C4�_\8%eToc�3~g���-��s
�J� ��--���N�b������yE��/��Wq�N-RsG����{�ݒi�Y��0�D�%�i���M�Hxݾ�s��ytr�����\�f�N�i�-��1���y�P����]Nq�����]t�dcގoRGZ��14>�d��iy�i����,�!Z�jkr.U���rv�E��r��+Ghi�lv�[�$�
ىKO�V�C�h�νk���WT�v�L�Wg���J�9�8A��'w5Yxhau����f�bKY�yk%GT����59cu�&��#<6��}�{��2�� �v�A����;�%G=��-n�ͩJ��l�+�(�QAfZ�Q��޳0(�ڶ�DE�m�U-�1b�DU�,A���F�ңTEQ�("�0F��Q��V�"
�b�K(�*
�EF"1TX���J�bYPe�-,1+��������ʶ�"�,b*+�YYZ�*��h�h1��m�c�+%eJ�EZ�-�"���ň�*�UE(��DQW(V�ZڅUU�P�Z�(��F%kưDLjJ*"����Ō1*��e����%V
���UA`�3(�+eX�c���}�~]k��IҔD+�{�ܶ�@Ӵ�;�$I�9�Os���+��U��b<��������i�����ƏH�tV�i�x:�쩔��ޖ|�4��\N�yԯ�o`�l�W�=���2]��kd��5bK��:�u��.��T3���I�R�O`Fi$�P�R��S+=f��R�v��fd����2�ݢ^3�R]I��Aӡ+�1H��0�se�Ѷ���Ҵ>�/|E����G��M�O^�Mp���B/*'�wXh	o��M�HI�yt�{)T5PKG��u���������g6Q�4��О����YĶ�+\��"m	ұ�[�<��
OB�P�{]Wu�jl�[c�툫�goa9���1����V�is2^�W�۫��r�4\���ɮW�@�^>�$I#����f��E\�a�:MO�@�w��2���:;�uXtb�yvpP��c��1D\umb�P�rK~�� f--&r7�k���嘚�<ʴ�^ӭ�ÿ>��˝(�e�iMo*��S�6��H�©g�r��ϝ-rК]�΁�5�n+���%eeT�K��)��YiZ�s�/ٹ�����ϥ�)}6�V%��^��f&y�rDc��մ(aU���F�a.s1�.���՜�Q��*U��:���v{�F�6�6*��8�������bE(=bF��\E�pY�&�Q�vorZ����e���Q>��jT�5l�K迮�Guf��o��|;X�9��m���FW޽�{}UgK,�I|�/Պw���H�+m�?A�6��;��s�U��U�e_��/u���@p����u��V\��S=�$u�.r���T\*n�Zd�2'�êF�I6�O'���mD�rp��"U�M������Iϵ}�z��	�Gm���fb�I�{g��\��Ĥe⾜��Y��ls���;��}���+�T7�X�j1�;�M)ˈ9&i�����sa����(ƺǊ{t�K`H���$�gV9:�k.[h��TLZwP�&��1c�Ă�0�]Q�dռG2��Q&��u%=�O)��H�;��(�Up��d��o:%���{H{v���c���^�jG�T��w ��V&�]ߧ:��^,e�CK�nt�I���I��������fxZ����.��[�hn'Y��"��6F����8��R�q������7*52z�h�L�����Y����2��y����S	=:E:p�o�l�ܫjK+�gs1:��\�ܗ�+.P{4S[��(#�*���"���$�[��g ��S�UAhz�Y{S���<w$�y1�>���SMEO޵*�{V�Hu(=r7"��{9�˔��2�E��z�+�/Y�[��r}Դ�;R�d ��m�b�շ��#�3����,�e%�w/{IJć*sj�Ծ�R-n�ÊV�J贬w��8�Y��E̆���B1���=o�[�F��xr�IO?L��&��0НjC�-�N��0�(���12ĝ�`�đ×�HR��,x���@�}��LX]ֺ���\��T����+z����p�w�6FG�7�4o�%�y��Ц��Wwh�����+���y/�YA�.��M�J_�XRe5v��k
�5�v!�[B��t�l�p�R�W�s�7Ji�88��舳A���uy�˪F>�{�mj��ӻ�Ѡ�4"kZR�6�����UF��2��Ե]�t��y| ��};��ba9X�.�y,��g'-n��m���л3/�6���b�L�y���`���-Z�3I�=I�!��d�����#/�j3ۈ��Mv�� һ4���爛���
<�H��#bOOd��3�2&���3N(<Hvoʊ)n�k!��2i�yr��b�Wz�B��D�7鵏ԇK�˓�`Fc��E��P��&���h��5=�2�Ь2��Ot��v&�Ϊ��*���%�Fn�|�����Ρ%פ�q�OxII��{���E���^�;wҊ��Ѷ�\i�h'=Q�e��-�Щ�s&�Y�,��|�E��[؉t}��83J�-K�X}I��,x�r��n4r��c9:=j�SPR�`�a��%�%�V-�S�����V�iJ��k;n��4%.r�6!> �}N�q�[{������8>K��L�^��"�ʘp)�$����Ѱ�_@�&�nQ%��"ڰ".�U�I���z��RkD��Sn�6�t�C�j����KVI\y3�'5눒b����bn�̫MU�0�ױ�ۏ�8?��IT�ʝ����5#�2b{`u*��ר��/u��U�:��87�J�l��F���Y��+g���\��'�7�]J���Q��)����<
�a%,�S͘�ڲ�/7����{�t�k&�ftf3��=���6���6'���"��'�ʡ���?n���֦OD����u�qkUuU��g]�"�6�d��\�n�����&S���> �f	m�}� �6RyR�#��.f,�9E�G~⑕�s��[�z�p�8tt�9o����d��� ]e3�='_M���|����.���Y��ٞ� ��6����2V�q��2��߽u�3��'�V��
5x���Q8����qc��^Ӥ��-��ėa�a���AW]t����OBȇ�J�MPŶr�Z�t��b{�rڪ­�&c1��o�<U�)�-�w��Uj�7W������Ѝ4]�.��P�'�	ۘd~�_�ZQ��4��Z�5D�N�FoDDȩ�'�E��c�t�9��Sآl�U85.�U�w�j�Wm4���Z3�[��H��z�h���Q��:�����W�1�V�ree�\��B�[�X����nwBt2����5'4t����vJ|��=W;x.��Y��-N�O��z�.�~�i�ܚ��h���[������g��{�� N�2 ��J��̶���c���dg&nF�ۙͅ�Ik)a���(n�9:-��-3���K��'� �L�{�{���y��U���ɠǵ\���JV�td.��z�}���QՔYk�+%�hQ�e�����WZ
�z�K�C�4ߴᗃ����n������,J���K!��vz��;|H{t$�2믵̭ڕɦұ��c��R��<�9���M�3��oFH�����_��-0�@��:pqW�mh5����[��y,� ��5;>j���Dj��ږM��	k�v.��b�x���ۊVɝǽ
8�Do��8��*�c�	�J�%J��NM�����]Ԃ��s'E2݌�]��G%ÞwU���Y+9^�GG8�ɏ/vjjJ~K�I�	!dv���f�\,m���o51�*�rW���6("�(w�p����q1��.��Ee�2�h�^��!�<5A��#Yݮ,�p[�ӡt5:�*�o�P"�D�J�3O����j�!�LFfs�Z32�7{(W�[c�T�ڙ��ٚ͜�e�b{�.0�Xr��ֆu�����X�T�4eM"'���Ɂd#�%.E��� �]�����¥w�J�Q1�D�	�h�5��z�N��u�Z�G�u��kNx: �{�Q�������ue����y
��8�½�eڛ#1�Y�P����^d�Ko�3F]0pItN��%5a�x;���e��W=|ْS�o���؃�M7�S`{D��)��8�b^��7�P�}�C ���Ν{p�{BF���T�=d�J�|����k�1���s��)�����*��������W��Ԭ�K����~�=����x�ίIu&k��z��-����IQ�W�X��CCJ�_l���`�C��ZӮ�#9��;v+%��զġ���B)7٤�b}H�\FI�(����KQ�9ge�)B�{zKL�ܶ6C�w!I&�A���3�
�Xp��q��tZ���W�rkU��;}sCw������M���k�2!�C�H,Q�tռY��Wl��ν���&����qr�ЍEB�,��9K�1NȱZ��p�`@ϻ���̲-�0cƍd��je$du��xV���ɍ��:!)_Z�&��Vwm�\�yU�����/`�;]@ֱ�o�Ӝ���Y��[���()�]V��7��d�(��k�h�x�䜻pF;E.g
�a��/u���Q�ʵ�g�]Z��to0���X�G]S2������1yQ��Mw3�nq��*�է���[7��ݞ�
�Ό���8
�]0�ɺ�̗�e'ȍ�&��A⎆�;3nլv�; c ����;����ni)��z�%�;/V]����n��Y��6�z��m3eh�b�"�2�\��GO�ҥBy�BE˧@.�*X�Y��
����}\��E|6�X���yo�+��"��_�N͞cnպ�4��D�ҳ����[�O6���ó��N��}CM�ɜ��Iu��D�k@6��3�\��ަ�yޢ�Y�-��lX��6����;��:�F#oY�����-���(�q�A�CoY�tci�J�u!�t`t���]y�_R��ɦ0�ܺG��.�0��ڿ�@�/���4���R6�mV�{�K��;ѹ��MS��=Mp<��'u]��}�\��k�P�j&3>�
��k�^2TC�n
��f����K)3�JK~�Ǡu�J�v����~U*Yk6�MB�DJ\��R��n��ka�eݡ�9�eb�9,��".݅T,nէM
'b7��f����ֻ�ܙ���L�P�r�\5k�{�$�Pf.[�K�D�R�.�t��=��n8%���Z���+L�u�h>�D�����5�YW���	H��	u�_Ed9��底��b�x�aʽ�N�"&q�d�Lkr��o������l�-��(��%w¹���1�wc�.
�Am��yh�n՝���2���ŤlK�Y�����t1гC3F{hS{���Mi�E��m�׭dd�ջ��Z,��gt+P��z[�x*�LZ��	r�Վ�<����Li�m�F��t�M�[�Z��%oV�ye�l&Ŋ����%�]rg6�׻��s>�r�[)�_�͡@Z��Q1(�F(���e����Qb�"�hX����̵UUW��8ہqj,F�h*e�(���X\�AĶ�#1��k**�
���URڈ1��� �%F�R�	�Z�q�DDA��[X�(��b��1Q*��r�`����VX��[r�Q�*�.,*"��-�E���*��E��ŭG�b��h�Qb�U�1amA�*�Z*#-.Z,AerሱX���U�KiAV�R����X����iDVڭ�,EX��)�QI�QKB��EEH��" ���Eih�AXe��*12���-\`�Tm�(��*(��	�VbV$|O��y�I$����MY���f�o^;k@�&%x�Y&:"N�ƍh���{.�g��/{Ѐ�I$q������R��g�{fEFJ��gw%R[�z]Ԩ�N���H�U�,�u���&j��ii��4�>���gnk��������µG��#���tޞ�i����V�8q�Pܣ�]�97�ho�ъA'Yf����4&���F��e��\;�#������gY���1H0m	"Y�SN�Tl��ak��%b;Cw�Z-��R
Pя ��鬜����=��4��^�)s���4���"�k�VsE��1m��ޯ:U'���]n��\�*7o������4'd5A�Mp��uɡFk���)؇kУ��Ni$��ۼ�p�Xn�v�SO"�1E����E.��I�a��#���*��{��+*UI��4ܮ����[gȽ�of��I�V��܊􉒥�w�"�q�,׾>wXZ֡\*L^��.�ˬ8�Y=;�ǚ�{��\SN)8n\��iq�ˎ�V�=�7��pS��B���=VG��idM�ގ�y����i����>R5vՊY�3����S��>��?V�ʴ��C-ҧ�E�`�ը��t�z%���w8j��Ou�ڝ��E�eK�(�=/$�%w��l��ov�~�k��Δ´�Q�/Ga�b�P9Ag��m�����T�^y�����=��Ŭ�v�!���H��q�3��:ګ�.^����W�>Z�]\1������}�~>���r�T�m9��+�qgrFo��Y�F�ai��J�bQ\D>��`ASb|�o=��4��a%;�7�+u�L䗛�)v����X��X�0Skq	I��6�3��,Ir�P��]l�K��Yƞ�X*�����s��V�,�;P�a��K*�A-̞gc�lOq��;h�ߠ�O=H^';�Rf��y+�
ڑ��­�:)sJrX��3��@�����3��F2�]�&ˉ��4�i�-��t-6,R3�&Rp��3"	M��_�5������s�ؠ��4��FbrD�Y�Wn�]��a��E9X!��3�`�)=	q���dyu��e�p�Θ.����{/�z(j��2Q��1�H|+��jj�fZj�i�7��Vp�d=��9���
��fP�U�������C��'m��!5���ު���Rx ��/����j�)�snU읖�;�h�`&����tH֢�A�,�a�����^�^\�,�UmDuqͮ�;v�(TV7)���/��~I�&�V|:�y3��W%C�(�XeL8}�<ֹ�V������g$5tiW�K͖��������&��ek�]�B/�Z����+>��-|�+�^��L�-)�O+;Im(�� ���n�f��'!?�1)W��8��+�R�e#u��:�`idut��U݁�
5����L�6¼t��;B
�{�~��L:ǉ����GM_1���v�l�Q+�N	�㦭fNOK'3�f����Μ)=@�V6�+��� ��띮1�r6R�w����f/ho�=�����r�6$����*�kt�F�;�]�Pg��x�[�%�R�*���� 7��\N�b��9�,�ĵ��J��k��h3���k1�#��s��q����y�ٕij��d9�B��!M:nI���sy\+���	o���G3=���m�b��I�����V\|�f�}�#��!Ό�PD�MԽ�y���%�n0�D)5����sB��Vӻv�qB9ɯZ��� �AsE�b�5oa���Ƿ�ݷ񳼜�U<�^�H�
�z��Ep����ȕ�Z���{�"���Y�5Lu,��}�5�8��vr�����4仱9�eU��nr�f���ֱd�����<صa��F�S����д� _=��1�R]��o�G)�}]����}h�q�
�3�YD����ҳ�V�Ą�=9p�i`j�SU������3�NJ�%�oY�vQ�@�ؒ"�2�O\�Im1�TX�:�i��jau]h��Mrf��}L�A\icJ&�ha��x��_�!�9(�=\�'g���^w����~H�(t˗�V\�*��c9-��l���
�QJ����}�e|��m}֋l�3H*.#5��Y��%�C��г5/�R4��a�1R�#I�e����Ź��3�?'���L�o)x$�8-u�b����y8`��U�7AF��jC�-�N�%�U,��i�bN�0J����$	MOub�R����e��5Y}�-���\���.p���7/5�Uo'j�v�,��b��=�]y�P�B��T8�phF;��iw.W�ⲃ�V���7}(P#TrGb.�j5�]�n�I��TcC�'c�̯[n����ߴ�a����ˋ���ϦЧN`H��D�y�hV�T,S! ��,�¹����X��-4 ��Um�4�;J�I*X���ֳoa%�c�r�T63&;]�R1����	�S��ո��}��X�W6Uuݨ^�*�}�����&l�K��!�Y��	�S����-��ub���-�b�V�һ4�݆(�]W���E�����1;�9�'���W����4ⅸ��H�j�x�:�x��[\�ܱ�k�=qnף8],bzy��T^_f���j�5�=�&�V��i��E�����ěj3S�qL4vJeQ���L���w��>L����K���//9�%Ԛ���v�kc*(�|X�X�饝X����kW���NHf�\+�e�eAǸՍ=wZ�K}j��ġô_��`�����&+kG�}U,І�yiM�5ۊ�ߧx,�99ENZ�C��f0�,�nzLS���V~�$r��g,U۷��;F�7D>k8��9��'���m�]&�[�(>�q�a茙�hɤ�w��r���X�r�v��{^����M�ܬ�g�!,���;p3�ZJr6qi��Ʀ���o�JD���W�'����?7����z��"x�Jk33-5]���FLT�P���L,��Jh&���'���:)]�`*c����.��W�>�^;1h�|�yi�4]�1c����{�̝ޙ�ż�=H�	� �+��Q�e������$�$��ոT�p��껻y7R �>��{m�8Z/�q�FQ�K��i��
p�թe=�!��y.ZȞ{PX�׸bEڑ����}M*�啊��ZM��n�t��eѳ=�0l7ǭ�����Y�B��i�&
��.�rY�U�������-&'N��h���ڏF�n�6�R��%��W���k��JN�xg�1t;oO��$m,�����tz�C䥇P�LM�ّk=��
�My�Xʱ��"�
5xώx��7F��Γ�[�[ulU�I]cM��m�VqA�B��F��IG�JĘX�BVT1m�����:ui�0�I]R2�;]̤�f66C00�����'Ӿ���,���랢�#C��AR� ��&ڲV������y��ô8!}�)�D)5��$nj��s芁{��LE� y�� �9��!O�M],�y�4<��UW&�WV�bȁ�
'�8�WYD�)�%�<�ed�R�2��eWlâ��)���j�M�?=��;�s�˨B샜�u�f�UAr���۽[�r����x_�S(�O�.��©w�Q�J���}�[i]<�:˗�/\y��c�ə��.�����5�rr���\�8n�@Jz�`ʌM��;HR��Eh�9|QKO�f)折�k+j���mO@�DŜͼ�JF��n�i���n2Tj''���u9��yq�l��#%�U�г�N�,��zP��mh���?jn�X��������i�/9Hz�n����6�z�2�nL��X��]g|��T>;��u�-����m[�GQ���Ռ���@IU�`�G��S��O ȇW�I�xO��>���Fp
�j��=s��9S�,lkӐV4Y�˹�p�IR
|F���W��"�:��W3}���9�bl�R0R�"7�`BŪ�hb����FF�w���r�F�#Ӳ�CaӊB:pǄ��]���z�Of��ma�2M��>�WJIG�TϞ.�:�&����vm��T7G"b�7"�� v���KQ��D�(�����A*�QK�vn���bD�:]�{�'c�z���ʰ1�Ff�w�E�]�˭�Ƴ��hZ���Ղ7�0�vZ�[�sl ���RRI�A�];^,	ݑ�7Pe�pڷ�ۮ�(L.�w�v����Tq*J儝�Q���#��sp�ڛƥ��留����c9Y{>ӽ�&oqY,<T�@��s+PQWZ��P�� �*xp`m�#l:Gwr���yM�ua��
�X׭*�EѴ�H�؟u����cɛL�Z5%�>�P�t���:�X:�&�!�a4��)X��=g^���C$���֪f��]�[����C�'�W�����8��3�ʲ�_V�EDdID�=���n.�. ;�]�tg^���i-�����5�t�;��)��a��5BC	�ֺ�!8$1�9��9�e&]V��.(�h�r���.Bq�}.!|B�@��6���D��.��O3�%�e�t�m��MX �"V�z,��j�s5��2�>xiX&���4]��V9��۲�U<�14���_�ѕ�+ +�ٻgȕd4��`��W�|������J�
A�C�T�G�������s։�b��pZЗ��+���U�xj�7Þ�.��L�ڑ�Ө�jax9�ɶV�m�W��:��X���C�SH����q�ݣ��N��Ģٹ(j��,��xj��.��5���u�T����.����N�Up՘�ٓ�	]�+��R�P{yNs0	ӷ���*�ze�Xl ����v�+�z���N�ĬZ9R58_˲����pk�;̤��	p�����sp�R���ƞ��^�0ic.��Eb�Ǫ�r�V�Q�m�rS�� ��� �Knd�5���O���ݼH���۵[F�7v��Q�o-�Qe��]�j����kY�,\��5��1`���tc�&L�{�汷�ᶱ��OYT$uxev)RC/��:J�bR��*����U��!F�Wz$9�A�>�wt疺aE�TTX�؈f��J���UVe��&9�բ���*�j�*#]3+.%ETb�Ub�tɂ.���U��cT�����et�Eձ@�Nj��IFi5J�te�.65�LL��J�ӃQV۫k�i֩���Y����Q�\W1�W5�12�XQ�j�Dk*�2�K�k��T����f
"�����E4�+(W�-�[uJ�jKVƕ��:q4�[e�[\Lʵ1�
�[X#�V"R�kmem��e��]SL�h�j�h���-�e���$��D��(Q@C�E�=�{��Yѧ�OP-|�W�F��'\�6.Ylɽ�Fc����ʷz��)+_S��Y�4�C�Ϲ�P��)�%鸏<���(�.����ڕZ2��CH�Q#�l��o����E*ȊQ-����cIg�{��4ee3{�;�F����ͽ�g�Ο`H���>~�Xp@Ss�b��x����܎&��(�i
#�:V��-Ry jc�s�;uެ����u�YU����\�}E��V����ĵq=Ԋé���wu}yn�+Kjħ3���)�v��=��u��,T��W"�m�a�zF�Hd��ɸ]|�gsc�q�T�SILg>�j:7�4vz\���Gv
��a��&s�����8j��4��Bu���g=a�W��~�C�-��z�=��vPU�Z#/tuZ͊;RS���a���á��)Ł<�r�97`�E��eӛF��S,��ֶ=��̹$=��h�D9�d���L����DB����M�%LIE�^9Ս��Iz����z`<"yD4[櫥�Χ�ޮ�ײ�XT��bP ��b�Ꝟ�ͫ�[V)q&Ԣ����\��NS�a����J����b�X�����m1��b�4��y>i���q�C��C�Z&��u81�Ѕ�[]��F���M�ڄ�*�'���gq+yY�V��590M1�O���:��4���'��e���MeL(���V��V��"��u�#Q0g7���i�S�����죩\*~�U|��[���q�2�PJvD��.Q{��9���4��v���G�v�*�kǙ�Ƥ�W֢|��6�A$��lJ<%�����
��DjF��z�mb�s�d ��%r�MtDű%.����G�ٰ���>��P{��=g+01�GL=����mno1��R�K��k����~����1@^r�N�I���ܷr��(v�f�#'�S�iF(D���u#��G8/Wx|ϛ�����z��ް�54����D��V:a�B�^2p^�눝���9�7�
W
�gW���ĭ��s�co��q���F��i��Ķ��Pn7�3�z�U�l�>�]a�.*�w�2{�-Mn�(�A��fpC���+}YH�9"�Oc֒��.xV�iM{NzB�DM�ds�Z��In\wnw�k�I���z]N��Wc�!O�7�@G�3d�1'��K�W[�zr��a�#�QF��R��S,N�e4�6���n�B͠������7r튊t��7��FQ��sQl#�ݤ�j�6�_.YZq���
9[]T�[�QS�/1��(�����#h��B��ۊⲢ;����w��U����X�[M5A �Ex�S=7vG���5v�z����LEg�i�2�{nt�&dM��|3ǉ�-��V�ٵ���H��fi�����%�i#�Q���-ފ�F�S�����C~{�![�.�Ii��������Cpvz�{dD��Z�G7Z5�57�i�4;vޜ:|БJX��S$h�V�ܡf�sUl
���7���!�6vQ�@�Ҏ�[Ȗ^����	��W��S������m�����e�V妛;U(3Ĺ�}0��m�a�s�Uj�p{���f"3�/�1�#9��V'p�.�� `���Z�������Ö�]�f�ú5+��v�I��'*&[����f�k1໛Ú��j��Ĥ�_n=�YE�}>rDOP;�R��}�Kp��r�b+Ѽ���rW`���%1=x�SykI�i�;>j�Y�j$�"�n�ND�1�]��R�,PE@�I:�:��a�}J	y�;�Y�lm`-��T2���N)�r��d���'Z��S��%�y���@���9�,�����
V�بRL��U~�n�P�#TL��ԯ4�7��g#m]�c�V�Jp>�Ia��MH&�J_��m�I8 ����)��!q��S����-C�X�HM�}J�J�*i']d��;�>F�o��=����[}웯&.w���:�d.�y,�Y�ix����J\z^pU��{����.ۆ��ͭ����[���I�����\�N�^�n5qsSV%Kk���M+��\��J��vA�؛}�W�Gj�g�����h��Η
��s�,�g}����v|�lmөHVU�QK&9�Dp��ql���9�lv��FUl����Yf+5�n(@ކ�J�S�NB�|�AB�z��a�I��ݥ�y��7F�	�;X�	cy�-|���;��X�#)8	x�΂�Iz͉[�U����:����Wz۠s�w���/@�}=z�A�$�]&mP�4;��µ�|��h:A�q6n�Ze3c�& t�MDe�*VU,��3�"�c�E�ʆl�� ��Fۥ��0��@�������Ml	b:qÒ^����*���hcoiF�	��m�]�P�^�R�\;Ȼ�3�.��T�Z�w]�x3[�	E�ς����9$ZUEV'\�����y\�}-&6��Z��{�k"���Z�H�t�˱k�(Y�9:=�M�p27����rb�(ۘ�k�����e091=Ӳ��(mAU�DgHu��"��$���e379�\8{��ț���BM�E+P����5�2��syY�]I\��"�l���ܙ��`2.z����F1����ջ�v��n���v��i�^E[ե�47Р>��]��v��N��$���U�N��[���3�k^��Ν����Hv?\�Rmr�lF��P#��a�t�n���=�U��I\�q�*��-�
$/4p��1JsE�s�lNH�L���{s�����@,��챫a�­fqx_�MqP��	��;x`������:�x��v�aĎ*X�<������R�	�Nе*3/&Feƀf����K9w������t�M�?���Y����~~�3h	=S3�[�l宵۳ӊLQ5��]q�{�������f��H��R�n���膟ъ��;],Q*+Ɣ��� �m�q��6�A�|��U���@�@��!H5�0&�����[�mZ������	�瘐[�a�s���V����UR-w��Pxk֩�JѶ�#�qF�TTd�:�[h�F ����7o/)��#)`�Ҧ3�sό�ӂ��R͊UƸr�;��r�^9�� n�>�z/-�L��8qGD�ħ&��>��ʧ�y4"ݦ�8�W`���b���n�)��1��[���h'*��#�C����l���<��b��r���J| �j��ʹ�Tqx*�X6122�i$e�'*n�:ɴ���':����%h).�����e?�.�g���R���j���Fگi��������c���5�iKaυi扮����l�vQ����ךQdؖ !q��H����J�;������V��6��ҋ�LG9ϽRQ�x�O*��9$�����|y��cwd�T���BQ��ާL¹F�y��kSbmc�V�Khd��AF���uz����{�84)3���T=�=YS�������r'���o�Rv��X#j�ݞ�g6c:}]���`�����#�@S}��*��:�r �.��u��dl��A�=X&�]�t��SwҁN�̜�=8M�NX=�A��;k�tz5�p)����-TH�]�^^mM�dlB
�h�sf��9DC^��Yx���z;et��X�[̻�9j���j#Jk�VĻ7�0�����n8��s^���7�f#���fZo!N���9cr��a��FOB� ��S�v'kR�穄;]�u'=���(ktnF�FT�"G+Z%h��yv�'���Z^���S�M��٥�cA1��6��zN�<78��{|y{Ŷ�Ϊp�j�X���`�#~�~󳞥����^�~+� �ނ�p\�ߐ�o��L� z�4:T��r9���f�O'�)�~���]�4u	rʳs(��Ɯ�-�V:��w�t�#Ic�+�AΡ%��0�4J���*��R|s�yh-!��q
">�N}lx�6n��;��|��&�Ѭ`9%����k)�ցL���`d�S�	'�"�,����+��.��uj��j(�f��
����w;;�,]&'nh�����Z�ʢ��N�\���):�V�X�f��`�0�oq�X@Dm�|���Y��GoVl�d�;�H�E����`vN��|w�1D�u[xo�ܚv�*�OQ��[2�%�ZA�[|
T�{��!�ee^�2Ѥ~F��NBVf����I:/��4b��$p��;ܴX)*5��S������{w�j+نj�Jd5
��s���LL��R9����iaG=�j 2D�8E5��s�h6�Z�"�.�Yu�kI�u|�v���B��ݙ�Z�`�ݠ�:��g��X[N�df���!u�*�)���S:j�ૢ�t�9
ykUg	����^H�sq�2��{3tt�c����N�7����\Ҝy�����P'x�4��#n� �(�k�ڲ�US�3w�����WP=7#p!�CCU��ՉbS��������չ�sr�@��uL�	(�x7������j�B�ȅ�y,U�̢�彲�n$.�dp��P��k�PF�l�*u�uY���k��v�pn�e̾e��s��L���S�X�ټ+_�����4ʎWfS3�m�Y����R��L�6�)"ɷ����wPvq��Pݔ����l�[-8������u�,:5J�Т�y�Y��̜�;�����Z!�ZkeY�6k���Ky/m����駓2�#Ģ�Ս�ùnD����2a�U�%x[q���%ˬم^L�u��Բ]h�AbJ���9������♄�-Ί�<��������Q�����OZR�L����ۨ~V����k��k�,�
Hk;ю�r�t��� �'�x�k��j����+Oj
�w}Af�r ��m�v��$�kZ��x��mC�KHb9�c�dV;FCw-�B��(:�v��b�T�-5{K���BUıj�Zѷ�ۢ�Չ��Ɇ�ݳ�s&��V��R���I\Y�lmM�[�d��G!�q9$�+e�n��ğM6��#qr�t��L��l�c�LB�ˁ��*��kPX�F5�k�-r�)n��AU�+t& �ʪ�[f�0h�ҫZ�B��T�9�4k)m�e�4��
����!KbQ��33-�3�p˙2��V�k5����qE\�n#i�fe�i�̪�q1�Y��Z��S�0q*�pr��n7Y�եZۣ&#r�p���a�SX���r�\�nc���m�q2�s.Z�ch\c�pk�D�ˆ�j��IEF")s��
�8ѕ�0L�2Tr�̷-f%s3r����b��Me2ښT�l��ij��ك�b���Zօ���W�j9���Lr�0TŶcY�nZ�Z����mm1-ŵUjS.�9]aQ��Vd\Kr�W1*˘b�S-5֊�\n%��sWWiV��F�r�.QyB��=��? �q*�^u�S�d�<��jv�o	�R�����i��%�nzW���%L��E%bOޜnnx�}wZ�	o�S�M�]ujE�Y���Y�1��H�d����;���OS����Q{���=)�#g:�l�t�D���\FHs����ő�B�,�Fv�U�Ʀ���cv�@TV�hE���O4z#���wڼ���"�t"Si��{��h��L��T�E{P�	4=@]	���M{@��#w����Xv,(�2f������%�;ͦ�e�r���=�}E(�yz`y����c�����1oP���Ԫ;^�&�S�ݬ�W*�jU�"�w�6X)e����)`�#���
�`JA�^���PhR}A�fc^��Ph	P���V��|r+W��׉�J���c.��J�=�N�P3c����d[�Y��s&�S�d���2w79�G[�E#��^ǁ�{{�����V����RgOW��pWիl`�u������w���=��l�xm�uh��SI���:���>H�N�P�5�G%c[CW�wA���9�+���){5ɚޯH�%��x�W���(�T�<��<�����k�Fu	=Bfau6�mE�ۡ!�˴`��gc.�]�bRЂ#o�1��s��"�����Z�hY��U`R�"�
� �i�!�w�x��OF��29�B��+Ȫ!I�Z�x�|q�>�kRv�c����O�	d<�o�5����W��X�G�j&�ڕ[��m�d@��py<�/\f�޻�yk9ktX��w^�:v�%�v톖��]�� ;����.�)8,����1q��;+��`L.a����Q ��]�[gr�Zr�l3fh[58�7F�Γ��,��SKc�	�y_Q��\

F�U� ��x��;���J{+ke��(}�D������қ51zI%c�'=��2�Qw��`�d� ���*}t�nN3f�`�:�Vׇa�83�Td���D��B��ʻYq�Z��徤E��W�d��xaz�{��C��N���Q���
gN�4�r��ߋv2��� Tm���P�``T$�F�g�rV|v���BƝ]u)����S�4���A!�OD��+�R"o�+ݠ�È��I59,Zxe�)x6��b�R�3 F��SF���mqQ�%KG[�t��M*A�4K�ܕ�rpFE�6�g5)���h�%��m����v-������91e��Q���97rؗ�Bhtf0��u����9�/�/!j�ĭv=�ޗ��})�����"l������b��®u�eK�Gp�5���;58^o6������m��۳��6("�[f�ri���"�U��;����S�F�u���5�7�e�%�Q�ٮ:�M�m[�[��Bp���Ԥ�fC�����^f#�V,��M�(�*��k�bhU`�7����(a�M	̻��c��3�!V�iZ���cQ��7#Z�SA<�^�D�S�.�l�kw
����hm��Fi6:W~4�݆A��!T�Ĵ�[��nPx�}�f���S+��B�ε��w�)�Hw�1_�Z�K��%`/o��WZ�x/�R�Fo�vfL�TE�88��l�1�ܮT\�5at�I��1,�/��'#����r2uu
錦�r��Z�7F��+5>�]S�^�&�����Zqj�f�ۗ�ne����g�[�@��ޠ%�
��Y5jc��d�Ґ�w��&��ATLtiA:�U.3���3��P]͛�WW=���*V�$�/s��A�,�����bUg`�U/���P���%
-\�íOr�-���Pn:�up����`V����5,�@b��z�����hb����"�f��FQ�)��L���>G"E�z�W�)�#g:�.6͆�g��r5p�f�-?Z>!�}~j���|����z �_u����I�d��lt�^#X��Q��*�z_��:B�5����Qk�c)�|y9����F�L։*ė�s[��x���z^F��oB�2�wJ{7�b�[ޗ�}}���au��{�C��LnF��9�|�p�Ź�
Ĉ�*�S�wr�6[i���Us诲2�-|$=4��C���j��;��L]jbK�GQIX�e��2���{���U�:�&^n�^��t���c%eeU�V:��D�>Rv	zeyzI�s�,�[n��zPV߼.2�͊�<w�7�/\�G�R1n]�:w�����덗��A_�&n=n�1<� |�D�>!�|U;{���$f�"�*#UU��^�U[i�ѓ����w�Q�=G#�ifI3KO���KޫF��C)S[CZ�Qm֍�nJ�K�:~R�y(��oPT��M�^�D�wB�g�i�Qx�u-��3��@[ͪŶ\	0�K8D�qm�����6:���������N��r����;�PE�Z#��]���5_e�-"6���)ox�����e���Kd���E��07�ƅ�{PS[$kfwe�����[]�#@�t{�8+q�ҷ�ԤQ�NwwCA[�f~R�TAPA��y��ýػ�m;Uht��3<��\2�Hnv-���D�y<�YS�����p�C��O�hÞ���I�k3Z]Sm��/�l�S�K���m���������v�.-$Ki���[���M)ʳ��G���V#�^Q�(�}fy�51���7k�n���-W��$e�Vq�Pv�V�ޢ1�
.���d��f���j�~�L��7Ԝ�]u�	��u򢶁T��x3;Y>~�'�+�ֳ���D��˹�Xz�-Knv��v��:XJ��S�r<,��Cz�G.	쎴�ז���^�ݨ��W2�i�]���l��;q��k׻j���6.�^��&�ͣ%[Kgn3��]>��ԾK�2E��]�Gcef���&N���1J�'�8~ُ�q��+��rP8c	��C��?�R��C�CU�gJ}�I��#"��Wd�O���p�(�R�P��r�Hpx^C���3�e�bn.���f\R�ѫS���G�uIm�(h5��S�P磶o{VW�Ԝ�j�͘�����s}�A�~�P������1g������|՘�O�X��I�A<��@�o���8ȹQ���aכ^֛��̈́a��פńDOGڱH���,�����*��Y*c)�[��`R]Z�^���d������S�#�B�D�W����)���-:����U�'�<���Ȱ;�=�jQ�Wo+#�u8�}\&g��\�%���)�c�2�E�-��63%���''���(�Th�<��չ��t�4�aZ�L���~1����,��b���g����<[�_b��ki��R���0QU�j̫���v�CQ���̋��.))������nl��V��̑��g��b�8��;l��h�]l�Y*͈M
H��zͿm�oM�#�Ѱ7�W
��lL}n�/bL�<�����8\�W0���lN�*>.U�-~���X,�ÏU�m��+��ð���i�M�`�c�,�:��G�CCe䕽=��RC�,��H�|����;��t�C�������0;��l�Ii�~���'$8�j�M��mz���4F�tzO(���� ����^٦>����\)C��1� h$H=1 i��S԰���5�ͪ܄�k�SQ��EB�
��4���7P�_���!C�E��͉���C��ب���:��vW����=ʊ:#���#�gr���%O���r2�~^ŧ�S�r���˞�.��0h��o#^^nm�z���^�k����b�����5�@��$OUfUЭֱ�`�g�0%D��|n�=-]
��Nl�f�@���wU	�g��!����J���:N��h7��y�3`(R�1��Ү�F���`E�K�d�IQ��u�S�,��ސ��:�*��#���>�G�+̑
�@�^�%����G.�s�E���n��<`;eyn=9�B�7�"+'5��Lwmw5j�/���Nr/�g� 9|�ܴ���H�D��pg��'��|t@�q^��;4���0dS�5����dT�Rʪ�	)d"H�
���� t��&�6�>�����V�b���bV���lG"Y+de��K�c^�M�1�"<��`�̐���^\�1zP��y.H�(g�L[�^��P�/�C�"�w)��ħ��t�@�e[\w�4NK�^��������\�ƕ
A���Lq�/����4f�vv�<��J�	]��]B�͝8k؅��\f�)��zWFf�����2E�bJ4/c��cX�Pp��Q�?q���?��~��J�TQ\��� ����B	���g�B	�@}𭀀l/#�~A��\"C�aACH~��$!�$���@�G�9B�� ���;ݒh4K��>���C�i�_��O�������o�2nHg{�?�Øq�ա�쀆��$���;�s��a�>my�	�8�qѮ�B!��{�?>o�?pB�0>��	��HH@$?�Z�,,�!���?D>�X�$�2`���s������>͇� S���� � ?;�0?��AP7�3��@�'��&!ɒ����'=����k��9�~_Q?W�?�S�����8o�$��̲B	�>0�y~:?<����$!�!?��2�*�y�)���z`\ϟ\�pO����6~�!��rNR�9�I�I���I����Y�d�~�>[�����RO��N?0��??��&?�p��d� �gv;'�~p�s�?���a�_�~<6vJI?_����}�����x}����|$���_�~����!����=�����������;���O�̈�	H���HB!��~�D��?jO�B��`��e�h?`xvq
B|N ~ß�I@$9��,U�L>_���	 d���Ѐ}G�9 �g��N8�K�y�<�2d��O������8�v��G H@$=0?���^�}p�	@$5���PB?)�� ������? ?�����O�>�0����7���g���}��I��������C?�������䐄C�>f���B/�B|�����C���>�z0�o�O�y�l���>z|Bf��u'P�H���}���C	��~����z�s��x������~�s;�>G}ӂB	��L��a��~�9�o<;O�R�����Too��NRJ� <� ���H�I?f~�0�_� �����A����d! C��	$�t�Y���0�5��>ﺓ���,��8�,�n�'�E$����(��y�9?�.�p� �Ƕ�