BZh91AY&SYS�L���_�@q����� ����bKZ�    � 
    �}P4I"U%-�1*�ZҒ�%JZ�$$�m	6jP"ڰ�b!+m"�֥H�(6Ҫ�D�VƢ�m"��(-�RC}� �*@��V�B��HT��*��UVʊ��(��*�(*�����T�fؒJ�P�&���z%\ �!-(��� �E�*�lɭJ(��T��EBR�-jR����Q*J%�ЪF�ѥ��I�0.����̢�"U�@l�P  ]���:e +A��u�cs;V0���ml��c����L��W-mf��s��3N�q����k�Xk�v]�[T+���:Ͳ�"����>A   \��O�ҹ�:։k*�[v
���s�
W����ZPv�*���E�`r�4*�uc��*�w+:gT R�n�� Rֈ(D���  ��wc�@�V�� *���{�R�	ޭ�7cT�w�<=J3N��TA�y7�TR�=��)@m�-���/A��=�T�ʔ�Im����]_�@ �w�Ъ��m��@��{v�[�Pt����U*R/n� OTxw�ޫ(h4oGz�B����hMnu=�� �����*�1A�U��:,D*U�Wϒ@ ��y���屠������ �^i��TR�
^9��B��{�PP ����T���p ��{\]�� t�v^��R� V� ���JD S�`l�+l_>R  ���@��̪�@��5BwS�Ю��(�MҪ���M��K�����U�:��`Uܧ�T�u
�
PJf �(R�>I  {�3�G� 8� Ms�hhΘ  M;� tw  wU�  ����@�N� vn  �p�i�**�H��$ ����а�9�wX p� 7g �wN
:ۋv����n  ��4r�	J�H*�UO>R �糫�@ �  7E����  ���` up�;��4 n��n�p Q�X `��F�H�fB�k*��|�  �| �� d���`50 )n��:n���àP;v�h � �           �������A�4 �~CR��  &  20jy2
J�~��      �2IR��    �II�A��L�0�`C B�M�I	� ��i��zO@zI���?�?���s�a��� H>EH4��rf��nw��e��f��6�A%������b��� y_ڪ�*�(*}�����%@W�:����g�?��vh�%�Ҡ ��F�yUW��D U��>��=��'d�D ���?��������dq��`q��fSe1��WLe1��SLe1���SL`q��Le1��le1��Le1��GLe1��Y�a1��Saq�1��a1�Saq��SLe1��e1���La1��La1��SLfe�Ld1��d1��CLd�1��Ld1��Ca1��Wa�	��CLe1��We1��q�1�e�SC`q��S`�dq��Seq��GLbdq��`Leq�1�&�@� ��G\dq��G&\`ddq���Weq�af@�\dq�1�� �D�� ��W\eq��Ge1��G�dq��Ldq��GL`q�ƙ`q��aq��G\fd1��G`q��Sa�q��Sc��e1��`q�fd1��a1��SLd1�SLe1��G\e1��La1�a1��SLe1��`q��Sa1��SL`q��a1��SC\e1��Ld&q�1��e1��Lfd1�1��Sdq��i��GLe1��Se1��q�YƲ���q��Y��$�8���#�.08���c+��28�� c(c#1�.0�����08�c#��&08�c)��08�c)�0���L�2���#�28�����2���)��0����08ˌ)�&28�c��0��c)����2�ʘ��#��28Ɍ��#��.2�����28��� c c)��2��c)��32���)��0�c!�&0��c	��0c�c	���;@�bɋ Y�d�4��#��0��c)��08���c	��08�c	��2���3�28��)��28�������28�� c�2c!0�0&2�0�0�0&0��28��+��0����c(c��)�	��0���+�.2��� c��0��� c#��!��0��������2�.2���+�.28��#��0��� c#���!��.2���+���0��0��(c(ccc��2�!0��� c*c
c L����8���$��0#�
8ȣ���*�"�2*�*.0(�+��8£�8ȃ� 8���(����8ȩ��8���8�(c*.0 �
�2
c2 �2�c 0�c"�2��2*c(2���D��(���(8���8ȣ�(0��8�#60(�)�&08��+�2���)�,�c+��08���.08��#�.08��23(c+�	��02����&30����.0228��c3��28�� c+��2�����̉��28����28��#�308������08���$�69��=���>�f_��.n���X��9f�(a�w��L�t	Z�m��e��N,���Z����pce�3>����͊Q���Q��xWxT��.�:���܆�cv�jqi�eI��P:���z�]-�n�L�!uD�d~%��֘��mֱ�YNKQ*\j;�:k58�r�r�s"+,�G�1�K��AP�Ɔ6�MGr��ͱ�,z��r%3or�ѭ	%�h&Ǌ�ʒ��R<�n]i�1	��ݽ��*@��P�d���R��m��vm�W6j/nSCN�رڢ��V�O5j�-��P�j�ρY��/7m�*�.h�Ƙ�d�),�n�w�93
D�ȁ���0;�mlM�e���Tl��*��͔0�՗��{ w�:
�R'���J���ڌ���7<b�j1CkΣwH��c`͔(��2��7�1Az���yR�YF=e9s]jW��w(Sͤq�5�fݽ�����E&�9�2��f��ƍ������+x��܊���[�#ÁOjn��W���zpG�b���`���]`����]�ـ5u����wq��ZIc2{����r�J�K7�7F�И��E����S�/�Ĕcӣ,�̦�۴
��h$E�e���f���R�Rx����W�1�b��kCg\tU��!1X4�wm��V�u����U�#:1:;���R�1:?���7q�ww��:�P��<�j�5e�I��ڵmǂ--��/�x�Mӱ� Z�dF������f%XR�{[V�����7!Rh;*������o@��mє��Jn&�����J��a�&cr����ඖ?��,�:��x�CE^3X���p�7�sQM�u����+M2��:��q����F,6�M��i��Ŷ�[��&u*�����L��6(������q�-�I̀*̹�b�j9um���z(׭Jz5</me�" ��!�eY�	xft P�,���"��Qa�9Y��pd1��Bfa`8�P���/)ǋl�w�J�X�@���n�Ծ��y%��FsLU��(fc7�V�k���P�(D.��j��V�,x���D^&�Q]�sn�n;]Xw6���@�:�:$4�yB�h�־��H�j�m��Y S�j�@2�:۴bWx���J��wY�A�T���M�QZ�fmM�4^�L��֥���gf�iǏ��#X�V��Jiel?(&��kic��Ք5ZT�&AeD$Gj��Y��+&OC#.9�]:Y�%Kv��Rލ�Q(�.�m��d�B�)���*;t�M��74�v$�b�t�y�^{�ځ�̔7q�J{���k���C֭���Dr�i�^�aM�ɻ`nڶ�a�dQ��z�;/>���Qi;1l3i+']���yY4;�&��c(�Q�]���v�f�L׶�i�� �Lʷ��5��cfT%�9ad!l@m�q�Ո��#P����Q��"��S�2Ğx�N:�����KMڢs�����1BA����k^әrè&�bK��=�/T�td�U3cm]��w�҅��V],x9��F銱�QR�z-Z��-D����j'���/.�L�Z�s���da��Ѫ�WdRH��Td�Ѷ�����Q��Pd���oh�t�J挘�8��v��n�i� Z��/Tg]�S�nT JO6S��z[0��wK+\l�k((�D^�����`�v�j�ڑM���Z/*�F�D	Z�Vf��Q�coR�"\ن���ja�{J���6G���s0�%��2;(HÊ���Ǌ]EWzTj��y��FKrTrи�RZ���%ةo]\X���YJL�N:�"��C1��N��VbB�a��X�m����x.qՅd��o~d�J`�N�����b�ױ��YP�Ǖw `Z������f�����R٧j��7�d�l7Y�^��*�B)�Xl��Rg��0B��I�v�7.�(([���SEY9�.�A^n��t��Qv�$ۈ-�ŵz��JO����lPSE����6H�5�Y�`X���bւ��k>�����o�*&f�ݙ��.��x��`�F��w�u��^��T ��5&��sqU'E��Q5a���p�U}����G�gCs�w���d��W�魎<�j0�V�a����n��[V���m�KT 
�w����zytQ���c��`��b{�u��*[��N�Ӻ�C�cA���8Xi<0CtSц�Mxv(�8)��L2-���Y&���j�7 ���3M�Rtb�6(nՠ\:�8�+F�Z�o43jS��),�nh�p�u�7Z��Niz�u�5�ePU��Y����Y��Z4��q�5����y��*�+�Zݱ��%�f\�\g+]����
7@�� T]�I��6X�F�n��Wr@kPC����l%Q�2õ ��kk01bKTG*GV.�eE��f&�,��eӡ�*c�2-�rm��Y�Zvu
1 v�;�%����Ğ!�X�YdS��%{����0���sT���r��oXa�X�Ta<�l��5eZ�q@��Xs��+�Z��Ki�ַd�ɷv(�ZET�6	XsV��SƵ�r��7mpQ�sZ�[xAA0iKm�9[J!�N]�Y�M��@�sw.B��Te�*����*����l9R�p��i�.,���#��X�D�BX-�t�֮�m7;۲�`�1�������@�5���J�5���h,�v�ȯ@���f�a�.k*���{q���H%l{�%H9��LkW��ӸU���Yv��ͫ��ɂ[�3S'�i�0�^E�HolФs(D¦��u�e@Ĳ���r*�V1�J���6*A
Lf+�6)�U ���X"6g���^�u6%,j�)V��(fCe��wo��ݺ��^^R�(�!��Yi��c���1�w[sd�g^ۙW�:vT8�1\�ئ��T�ѷ�An)� ���h�5
E��jxPy��4
�Y1*�qYW
�6Lcb�����Yr��s$;*�Fػ;����۱[6�i�ƭ4�
X�b�"���d$��8B�f��Ha����VԸ�"���%��j�[�#�ؗ0�U5�9sr9�����`qܙ� �R[#I�wT�Ө��-�L�i�������D��� 6r7
�-L�+Jv�o+*IF��㙩��>6w2%�)c��!��)pS	)�@`k-¦�7�I:��!ֲ�q
��Z���t���0H�Ҵ-b�� !^VL�4�4�5!��[W�Y5�wL�y�� H�)*����5x��P�Ÿ��% �]�z�A�l�&����3qᎱB��ాxQ���aS;�)wj�I�E5�"U��.����V4����!�P�J@�5I�U1o�d ��v�M]�U�#���^���F�!�S�	6��ڸ�*�V���M8�6F5:�Y��8턝=����`�[E�yeՆ���_o����|� pGt�ʛ�%�2��J�[8��pU�ފ�v�%"T���ۻaaģ�Y��-��:��K:��cv��XI�v���-�sT�_c�vJ�Ջ&�yEp��w��5�\���ŁRY�L�	�q3@:��Bླྀ�C]�4r�[���7R�,{[��[SF7v��{+\��`~l˭j��ެun�uQwYTX��b��T7��M��1�B��T1�=wtPÅ��T��,zp��f{�����h6��A"G*N��ӆ+)�:��
��B�.]�/$��l$`ɉQ���w�qcCEfk[��E��dN�1����Qw���y0��ї����v]e6�l�ic����^қ���B�Aem�1:���{Y	с�Գ[j��-�PU�^`�F��Q��!&��B�
ͭ�0�"��l3��=��/T�����(H�Q^H-��I��B@�������ܦ�I��[�n�Jh�@�	�%i�	�K/��J��U�M�g!�b;�M�t��IE���qIR�Z"�%�1cʲ��l�t.=�+�M|���;e�v��Ԗ<��b����-^<Twh�Qі&�����1iU� ��J�&˫;/pj��!��p̃#j�R�CȆ��k�E�gpG�����5@�e�t�6->7�hᕔ�MdXÔnm�K�a�mn\�j���Ӓ�p���Ջ��`kP���܄�ToP:%�v`�=Zv�E�R���^�1����+St��Xhŏ^
N�ѵ6H�N���;Sh��Ul�a��MB���P�c.�b�'�R��wa͙dȦ�U�S���n��M]�v:ge�wm���MXX��L�rJa�iՉ0mf96l�n��c�U�z��	�n����+K�6�Q����{{-d�E	�1o�l��Ɯ���{e�h�F���v̼X.��n��0��Aw��ɏo�ۙ�H6��
���w*�Ԓ�~؎,�/aGEL�,�Ų���Jj�B�ݛq�7KF4����U̼���ĝ��[N�WS/j���[b����>��
mՋQ]�ں�Z짙;N2m��FƦ���ti������!x-`tin�dBc0���ໆT��(&b���V1��w"���O#-�X�˷V<e�Qt�rR�����L��͎���@��9na��p���q��"����[#
��B[7A("��CvSeIOXG/.���kS�oQU���x���S�+-̡�2��,d.n�l��z^R-ʂ��#y��¨e�P�imVU�JXF����&UO)i�Ȉe[�m��L֍6�Y�c���l�:�)SWa-��#���+Z�A���3dy0,�#��ft��Ǻ�2â�5Usn�9D��D^���ǹ��Oh&��kqR�
��l�wN��7vcY��X�
s]`�KN
zn�&�"r��-�L�S��b����*���BY�g0Î��<�Gr��Ф�3�A�o�jĔ6%����Uj�D�)yw����7�ٮ�{y8�`^�-l��+a��,"3� ����X?[wS&\;{c&Ty�k$`���xh��j��Z$Za�N��t��n�N���}�"0$!��^V�{�l��bz0�2�a<��k�S�J*G"��L�+H`m�!ڱ�U�i
2�d����w�[m[7G)Ҹ�ȶQ̽�Q�v�m�
�rJ�2��X�1.�86�P�31�pC0��WR�:ײ��.�[�*�^�C`	��dOI[j�H�48���FL �t
�j֪�����nP��W��Au�k/Tǥ�.T!�j��6pA��L�x&Tx�k����i:V0K��ҫL��&ZvAɎ��\�ڀ�L�șQsK#\QV;y�V����b��;M55�/*-l��5M	��'X���nJ��E���!+���N;�3�h鬵����L1%���=�q�v*j�`f���c�)X��;i�-S�ވ�7���*�l�Go-��p[K6)�B�y�vt*����F^R	$Պ����-ЩTt7*l/v�B� ����2����F�6bZ-��6��Zf��K5.][U1o�)Yc1�^��8+�rkLSD��Ivf:�ې�8�̄Ř��j2�K2�T��ɚ]���f$��O`l 	RV����yc��'D�ڲ2n�n�w�G��.�m�˖3m��j(�ڕL8�ȶ�<Zn�wlb�43&F���2/I�2S̾4ݺ����WK�IuK  ��|nC�3�5b"楋d�K��XU��9&�8�Um*u�'�rb㰎dېS�;4t��y�Bb�е/"R���ZD�{�UbGzc�B$�۽��Iર^n�����P��$"�Z���YsF�{M(�X�S�L �l�豴��+����Z�ը���k(��40fȪ^4fe��F�6+EcKXk1ckv�nV�pd���F��ov�B�����zvX"P�J�ݫO]
�6M�u��f�,Kh��68J9(Q��r�Sw�[���ѝ���S]�-�hxHnMjcI�%խNR�ؗ� ~���-�/��YiQ��)�����a�L;	�I��^H�1e�֚�GQ��*M���-@]*�@�]�d1�����[�EI�+��>e�s���������oJ�t�m�
�f�I%�d�'M��=C�ݛ���aVw�l�<74�A��o�%�%�|�*h�V�$�E&��J)�BaD���Y^&C~o~ˇ{)������v���2����VpxZ�̢I�0!k*�ӸC;g��{M��q�\�V��ִoF��0P7���U+�R��.&�����ij�;���I)�֬��Iw.ɉ�_H��L�1$�;� 3Ḣ���3|Ex�;f�}�b�Aὸ�#�T=�L�N��ا&ъ�7U���+Z��T�Z����h��m��|򖧉�J��Z��]�������%#��:��,U��,��ݍ�"�D�K:���i<A2��h�&��0�@�&|v(6����ǰU���p�r�ERk{�)A#�q�
��!�=�-(�8������xy�qi� �I'	�%��Vc�C��Y*���_�a0�]H�0�3��4���t�F`�0�d3�zaa$ޛ'�Ho���L;��U��Q���*O���F����LKS<�庻���-�"b�喊^�<sO�P���Z&<M�ZɼM��F�&��E��,��L�M���mv��a��)��ĩ$	K�-n8R��,ԚV�E�*F"�rT��4�$�@�p�.@3��*ɡp�-#j�Ke��"MU$�Z�2%ɵ�装2x�,��p�<I�p�{M��o�x�g,�3i�d!mfGi[�z�Rmp?Z��,ړ�4� �[i��$
�%��+���[ղV.�8�7@Кf�H�C�	廖E���|���)�Y�C�|wH�p�oOP��z�<�U%��K[�wJ��NP�z�'J�x�+�'8��a��d�A�e7��&�҉��o�X�?���߱�����K����c���*n��[��u����;h+�K2ﭮ��R��{�d��
Z:{�͢�R�u���'{`�#n_0�5H�u�����=�H�9PgI|������b��/)��S�.醏j����Cw7Wf�N	�:s�n�-.�br)^��+~Į�v�Q�#���Б�Vu�+`3D,ד�J�N�g"�ǈ���]ǲ��g1��l�j�ꩬp��ΞS��c�Fu��}�t�7��9���1eҴ��q��q��Gb����7���7��t�u_�Wv������&�ib�<���7�����؃އ���oBȷ�cNd���;8�����ʌhݮQ�T��YW�����e+��nw�{�[
ŉ��˴$C��Y:& ��>yR�c;�n�BD�N�ݮ�����OkEӦ�2oNǬ��S��x��dN��I����8Q���jeV;��V�܍ɵ��6�+&�UDX��̠t^�kkj�m.�|:9��d�����9i��#ӄ�ܫ�]u��Ȇ�`���4��C����w]�nY�wξ�M��LAJ�eԖZǿj�7��a)c�rݶ9�dך��w*朥�aEA��ʌf��"V��/�[�/z����^�:�*�����e�6��.�n�aR;5wf�b�2Ջ�էy�n�ė:�U�K�R���_ft��˺�s�|�x8��ݾ��ۖvl�U�T�N@a:�ưR��ӝDr�n����r����#Er���+�Vk[�yW+f	
v���vÉ��B�Ɔ��e�̙�n��f�W:����v΂8lrJ�.zv=bb},fj�U5�f��>�M�.��8����[��_����fK�����!��@$G�RԼ ��w�${��.jL��}�g�m�M��Mn�H�W�NΚ+�Ы���T���od�wr)ڍ�V*��wW� ��M�9]؏XF��P_`ב5�e��ʺ´͡>ۮQG*+�;���h[�ו��%Ս�{��nG��S��k�pN�m����\ؽ�l<V�o���W�a���<���ӝ��P��r��61�w%��Z���.��֭c�T̙]�a=�EZq��Y�t�@��a��^��)t�mM���꾤')%��<�=Pv��ن=�V��yь	gV\�l�sJ�v֛n6c���ڭ�+����yq��2��VAS2m�t��U�ոG,V�Mr�R41��ʲ�@[�������Jy2��_P��5��l<�&3
���d���v�!�ٸ4ǝgl���"�vp�C�nb���J��2f���x�[��l����vc���ǝ)�{�����y8f���)�z�]UTGfm6�}Z6�a��\���hR�EU�(q��[%I\�U/,"�:{Z�t��%xiq=�$,2��N�m����'*8l�K+��]��P2��im][�4r����2���R:ڜ^����n�m������C�y/×�!2�X���o��D�7a���Jq�=�>o�0����LP4Z��d݅�֓á���S��V��8�̬�����9����W=����1��V����t���|BQ�U�b+9�țr��*�[��e��
7W���֞@���W%J�ʎ9���Ȭ�[E�n��Y
��ͷ���k����u�]���3
�pmN޳Nԕ�&�='jvZ}Ǵ�]��lAC�.��ܒ����v���Iì6#�}�o6�Tq�<��V�q�u!	�Ay���J,=rfr�˝�o���٤�$�5���/�m�.�����l9y���Y� z��x�j�e3O��S���xS��l�w�^OP�ی��G]n�����=�NtI�����o�V'-J��9I��R�)]��0pmE��n�%�7[z��l4�BX������19��]���c̨��Ý���>ya#��R�3��kxm�g�lWڹ"�=ް�����;��EWK�ݽ�}����.��p�DN�-��N��=��ݾy�ԹWeK[�8N��nme��Ϗ^y:h3u�D�����Zz�I��:��[T���D�����)*����Ni��b�lsOq7ymV+f	I�̈́- �n���e�8�wH�u�]�l�Spi�3:Z�nA�&���o�l�P��b�����q;�+�YPt��E(�t3ve������
�	�]�)�A���rא���kc?t� *[���qY��H�}|�%�՗���(��� �#la�ئ���=ٽm�+$��y�puf8��k-�Cx�^mi�WuL����&�����ӗc�7c����uf�U�����I�v�#�|�_�3�M�1,��m��x�q�^;y�Ji���)��;p=����v��n���S����7�aZ���*T����[�;nθu-	���/0��؃�>� quc���C�<�!�S�;!�zA3�Vc��/�w'VFo���'SQP��@�T��Wp�+4SM�@���3Bh�E[y��=���	�
tSsh��s�y��jiɻ����y�g�,��U	����`�HѹF�]]��չѭ��%+Uf��k��MK�ӫ��i4)<��amʵʳ�\'v(�jW��X��z�E-���%+u�.�r�z�TOU��#]Y㎸�y���J�D��Mn��M�`��rv웂��q����e�w�`�+�v�_fct���tƮ9�������#��b���QT�u����d�����������$�͞(��|�*i˖k�L�ӄ�	"i�/FMb�;��_;��5�j>"h����*���N<��rr`}�٬�]�P<^+�(�e�NU��D�κV���ևF�;�c��o�v
r����$* ƹul˥fm�gi�
�:xnrb�m����p˺�N��=Ah��S�
���2C��{��u l�\;O[�gbZ -�����,�Of�z��h�ʟ�};+$N:4e�cI0�<r�<����$[ǎE����w[Eޞ�
ѹ�d0����:c&��f�'#/����oRCu�:=���-�Ǹڱ�F�ŗ��qr�ϣWc�6[����)o^.�4��;8�Q�V�
}r�ݸ��:�����E��^�r�U�)�77tfԣƆ�ٲfV��E�����E�#nm��M*�y�w}x�N��@��KE�y�Kn�N�B�I�P���9fX����2Xn��7%ؒN����[l��W�]�O&��)z�Z��vwnU��c��NQ1@�i��h��<�8Roq�1��*an��p��/�X��QS�[�Uh8)�9/��]9.'�]������0��S����3���� �IU5&7e؉��#���4FH���Ҥ5��K�u����f���O:6�	�$ȫ]ٳ�+�<i'�.�*�uzm�<�����L��h�૰�s7�Z�{�Yz�Гz8Z\�ue�7nF5�����
����сmU�k����M�^e���o4�*��ݴ^��Ŏ�VM��Ԣ���+�m����nئ����A��aU����r��S��$d}�JH���ur-�<"=��3��rH��C7m�gu!\��+5�I.���n���4�q#��ז��N����v���[k
y� p�^�Y[i��/3^e�E��ﮥ��Mr�Y�uك"[�S�]�lq��u�V�2CA}�Nq�nn�#��hR���0\��𐸋�h��'S���އ�l���5�&LQ��M���r�W=-R��i�Kh���6���rf�;9����w�Q�x�p�0:˪�%�A�J�ղ��z����7u�Lfa����۳�e��:��ʻ3hT�
C�[2��ǕpۛR�[]۶~#�J]w��f&a�Gv�w�ֳ0�Yb���s�1�m�2n�v��J�N�עA�\Uu���:ieq�gl�A��=�|�ZԕgG�L��հ��҉�Mm�	N\S�����P`�laY�s�l��.��nD���̬s��`V���l���
��n`c]^�RrاA}�m�_mH<��n��κ]��16�R��[乸c's��.��d��^]���S%ӥA-`��=y玤��Ve�r�㊆v��u�n+�c�˳M�
��t���}s.>��mcb���o�͂������W ط7D�j�f��%f�Cu/����,����b�{�Mumm[��"�s���q@�=URm��b�ˊ��S���]5v��l�=��uJ}��X����&��]��ZymJ��e9�0(Y�7�7;0�1%�B�E�yѓ�U�Ԫ�X��
�s�i孫6v�M�x$�/v���s�;Ö.Q�z�帑��{���`;[싅�4X��N1��_���w��2�g"y8N���P����v�
����6ݽެ�x������з.fu�=�6��WWPܕ��J��[�Q�����C��՝x^&h��ohB�,k:)N�����q=w�b��Ԇ7��N�8d��n���T&�=��2WS{@D��޺��vnr��*���� 4�C9��2����^W)]�5��B��9e�rճ^������y<��J�u*����2���O��{� ��S��	/k^��涏P��m�D�.�s�g�݃/EQ%�,wj�f��[�1m�����U��Ǖ��`���
�<�g�Z��y'Pj���tk'S���WJ��Y}�𮓙6"����-[�w�;��J��ZǤ圽�6�Nf�1�.T�\���ű�,M�}����X���5i?;��K�޽�U�
��{��s	�����5|����D��w:����
�ғ��*f���ڂ=�]c��1wo�/,D�s2���F�����X��*&��9�v�4m�1Y�S\�P� �8�3!�����nǠp����$��O=SS���.EAvtG̪� ca���57s��y�Q�%qb�=���Y�L��a���en�;�}p����d�<�W�%�c��!��,AH��wՎ�Flۻ���7F9:�]�ݴb��ǆ˗�EvK�eԕ>�"}*u]	�P��g%�����(�ӝi_A!��mm��n�u���}�K=�&d�b��g�/�5/��������8.Z��lؑ��ng.��F�aѠ����b�����J�{�nk�/�H`�r�a]��_�S��ȶ2îU�����B6�غ[��g['4*�f�-��.��.��]��le��L�&��[r����+Q�j'r�����$*�E�G�^%���py:����Lenk��%9Ǽ�ɑo	�l�����􆁱$#,�ٗW�\��'v'�75��:����#1���$�[�Q<`T�ݖ������sʶ��x�wKV��.0�g
F�Z͹8Q.=;\!zvm������-�����-�޻V�����G{c+����v�k��C�Y�\X��u5Ag�X�,ӀQD�Ϭ1v���D���:���|~;��ړm�o��0�s.#��qkj۽ᙱ�˸hoN3i��t�����X��^�j��p8��z��KR�1�y���.�9з;v>iu8_��9�\M��Ƿ2>�b�]�Z�tʂ]΅��I6��jK1�޹Ê7Me��Á��K�� �q��#�3�A5|�q��g-�- rL�����ի�:�cm=�ݨ$�V�z��4�X�.+��xw�#�7��ˇ�`-Էڪ��63F*[�(����v]���eI��GQ!*��^UU[��+*ಲrn5ζ8��WJ �a��d��Y�W.ŧ��5l�=;H��W��WWj�(5e�&��{pt�a݈�r�!e�:]x�L�Mu�á��P��nN �Qv�L��s(jXnӷa��uL��jkj�Cl�{[���I�;۳}v��}�h낊+d��[�����*�4�u������l9Շz��ޓ#L cE��c��>W�A�~�}��{����WaL���9S5xI$�I��I$��-�;y��
U�Ʊ��g:p�:	�^�$�9��I9��I$�I$�I1F���e�qC5虣8GV]��=�No=95Rוd��8I$�I$���=�S{�r?3�ܽBu/�}J������#�X�#Ԡl����䇾���=g�y wrD���'�X)��=@��!��=`�xr/��@2�	߬�Q�����K�JܝA�_p��Op|�=��ʽ\�k� ��V�늟?�XP��c����� ^�߮��M� �S��R']b>�|��A똏|�{���`�@��>@�=��=ݒ�+���u�T�vG��S��� |� ��TDG�}��~=�����E�������>�QA�`U�?����������?�����Gz�w_�rK�mdL��&Z=����rÚ�ju�)��S��NgQ����I�p��m��jU��	x/�v�Q�y�2<�bg]WN����]X��6K���h�G�	
R�>"%�v�ݵ�M}�+O2�k�f������Y�j�*�Aqh]��Ëc�'sl}�Д]���Yp�ө�|)�]�j�]��)�h�32�	t�b�N�#�{���%{]�ϴ�ff���I�c�D04�B��c��D�m�<�vE��v:������*�<x����=�P�v3>�\�"�2��-�f*��tR�Y�����d�s�[�5ԧAN�t}mv+�̈�⊨C�Q����Kz�@̪�Y�]��.�=:�P�k�M�ͱ��UT���PM���q�5^`9r�V�^&�7�;(�U�]�x*M���7�[����q��ne')����i���Xn��z�iǵn,r��ѝV�[�J�˯����n��R_os�����O"�EXՃsI����&z�x
�Ct�=��e�bĎ[A��nȡT&?.�q���lK�v���]xCg��]-�j��&	G���mUC9��N׈�]���6o=N���)�^c�z�&k%>A�!i��p��� W,��&�����&-����ma�h:�påkL�p�8��ըy�,Շl�͹�EQnu���z�ޞ�k��G]u�]u�]tu�]u�]u��:뮺뮺룮�뮺뮺<u�]u׷]~:κ뮺�u�]zu�]u��]u�Ӯ���]u�]{u�]x뮺�n�뎺뮺���]q�]u�]}��:뮺뮿u�]u����x뮺��]u�^�u�u�]u�ۣ��뮺��Y�]u�]u��:뮺뮾�u�]u�]}:뮽:뮼u�]u׷G]u�]u�]u�]u׷]u㮺��]u�]{tu�\q�]u��]u�]u�]u�u�]u�ۮ�㮺뮺�u�\u�]u�_n�κ��y��g4s8�s#7�٫֪u��C�ݎ�fiM��tYRt�)-�wS�w���57�UP����,��SZݨ��lc�1U-uj�O�#�Н������e��0*�.޻K���Ql�}����zt��vԜ��Inkn�*��{�[-�Lp��]�jɖ�r�e��e]`�]s3�Y���Ö^���a��ʂ kt��gk�5�WD�bsǓ����D���˕�̫��RC�;B���u[0�DR���KZ6���-ty$}�wn��]���sV`��a���ub9S�(��y�c�v���0Y���6�*m�=p���������ih@�kd��]�K�f7�&Q[W�'8�Z����䉝"課(GK�a��YM�����gt����5�y}i������Lz�=u�Lf@����)���kQoV�:+\r�HT�)�����ُ���o"��@�S \�S	$���Փ�(�Ę,�[��)-l$�ԇ&㱌mn��ڦ�Y�u�d�G[|�C
]Ӯ)RnYy�L$��1|�Ά�{�BD �o҉rS�n����1�t��̛�z�ɻ����g��L��;ufݒ��rf�%6.w^��\)^�/�b�{A��(�s=���<UH��Y�qm��2���#0|�V᱃���K��w>���kX�^�GC���&>�Y����''�ݗ��3�G��ӯǷ_o�_N�뮽:뮺�u�]x뮺�n�뮽:뮺�u�]u��]u�Ӯ���]u�]{u�u�]u�]~::뮺뮺룮�뮺��Y�]u�]}�뎺뮺믷]q�]u�]{u�^:뮺���]u��]u㮺뮽�:뮺뮾�u�]u�]u��]x뮺믧]uק]u׎��u��]q��]u�_n�κ뮺��G]u�]u�ۮ�뮺믧]uק]u�]u�]u��뮺뮽��u�u����]zu�]u�^�u׎�뮺믷]q�]u�]u��뮺뮺�u�u�]u׷]u���*V%�@�ͥ��MގI|❍3g&ef���z�c���T)�̰��SF�@���g�
�.��΃�;u_w3��p5�����8��;1ɚ�`�ّ�y��4% (�z�S�.ۮ�}Q�T�7s{=¬8{DS��1[�q�(d쾫�.�4i\ڤ馕�n�\��k{����),�;l�J;��e�9
Ž�I8-Uy���R����Z�Ю��6���݅ぬ��H��;u�#�!���g	��x���7�\͢ތ�Z����A�ϐ��c,���k���jɹ/qr��(߾�}�1�ڴW�ŉ�ب�޾�b�Է�/ga����������`�{hbC�{oxt0v����쵯*RckV�5!Ƈ]	�2=�Q!r8�c�9Y�e����"��}W�ׇ{��2��S�^\T���[*R��v�Ts��E�]�0i�L��xD�Rz*�Zٕy)�2�*�WYUW�z��+�S���"�2:�0�.봌�.��������#le�X�,X�O���$B�v�z�x�)gY��+������7""��U+��N,:�L��ǱLwM��A�NK�ĵO)/{��V�Q쬻PvJIߞrt���(�@��u��o	�`ޜ��B��v�Y;����2֞���FeCYhA}����m�� ���:���<Z{aCMb�HQ�/*D�L��Ԑ�F
�����E	����V;Uf�3�Z�T���W�b�Y�/3k�&+�ݰ��Mx9�u��wv7`+[wIV��̻v�E맂����,U���c����>7��[{kmQ8%�v �9!O��S�c޽��I�\D��V�H-�d:�����8(��9�[T/ 
��	v]��0�����D������9S/�������of�܉�rV������ڨpɅa�'IV�I4�&��������YWG-K�6�;��oaOP> ̪�6��҂��E,�.[e�6+��c�t<�	ڛ��m�� �,������j=�JCq�rL��E[�(�-X��/��	(>��|�je�)s��/��y�T���$V�'�;��Vej{�5�{}6���34}��z�
�|h.���/F<��b(1���X�^�m�s��Oh�X�T�Ah�y�C47�۞Э�T���'o��Za_W��L���U��Nf�^})����Fp��J�����8$-�g
`�t!7_d�p�W齗w�V��4y��)E�-���ܨַ�e�ݧ���e[<&U	�c�X7�+�V�٬X2�U����JSg�9�/�JػW�9n��������{�{1��+�,lWmL�_`��8�x�tCc"���qvS*We�	4�v�ceoٽd�I��ۧ��*h�J
b���zsV(;^`n3��0���9�n;$Bv��s�N��o�3�U(S�z�Fa5V��x��^_^ݎ��$�u�Yc�;��mR[�}�l]r�v�!bq���ᕸ��y�j��UMCPkۼ��O&#�\O���d۱`h�WX����puZ���m�B�P��$����kr)/��:w/E��̾�G}=�t�_W@Y��%J��mud��gu�ٍߡ��KXo��־-�b��|� Ղ�-�Y1���G����]$� }�H�w���`�.;�Hݧ����m�KOc�;ifC�/d\�A��=>d4��Ս��B�eNV��a��Էw}�!��.�+�ky|��̥:���\)�Umv�%��s1o�,x��v;���'�ڹ5"�}x��Z�#�,pvi+g��p��78n��f��W ��3y���z�b�yShf)+�'��4WJ�s�M7�ؗt���wZ�o,�}�"rU*y}�Rʮ����q���lAn�T�$�j����v��b5�'�%>:�eE�uֺ�
�����)98s���cp�2��n=E@
b���aX�ix�kL'���T���@�H��[�Ֆ}w��VЦ)g_�B��k�G�w²�-�Kѵ��\��3t�M���ٽ���t��
���%��=��'�/�]f��h�ezO7V"���k��1Iۄ��v3WP�C+��sK5T�ׁ��i�@�	s�����U�/U�&� ֏D�v��^�htʫ���p�eh��&�y+l�&��ʻx���<m�p+�|d�x['\+s/*v�Ȍ��	l�-4��MDrڣ&��*�&�L84:�X�3`r�Z[Ke�ZK���:�=�Ȑ��������;�W�A��M'��Q�m󛋒J4���f�;����_\!�����!���.�FX���á�z$�2I�t����QR�]��K��^d�9�3_V� JzބNP���uӇYL:�ނ��:��k%����(+�e��-�m���V��xÜ����y"y��}L��y��ҹ���T����ihn�.�ig_*�ɱ���#�l]Hĕ��{�����fR���
�����֜�+m餤-�F�V�ޖ"�/�C�U`�% ��vV�C�v��'[����Sv��k2��ə�ي�>�k-��
iH�S�XY�a��E����P���oX۝:u��뻪[���b_ZT+�R6��ЩTt�I��}����sf�4��U��I9�/꽋�kz��?;�D��]�`�9���eIr��[QF9�@n�'ِ֭غwY.;��mX&�d8,�|�tX� �*-�+��h6��uѤ~�'@۱bh�b�xR��F�,�P��%�}45�d����EN��ﶢ��(�]m�Q��ۉV0�;��U%�K���E}�z'x��n��r�&^*R9�J�P�b�-�{��?��/Q��o��US��3��{xƝ�Չ�c�E%T�m$\����F����L�φV�4R�e`��ށցf�)��z]����qe*�����J���*gL�P�@A����6�_:))��om�uX���Mmp:fj�p��hl9}7� �($�WMf���G��i,���
�^��U3�B�k��Z�R)�r���f�B���bv
c���y���X��}ԥoAwB����o�;�B-_umZ�D�p���Y�UuR�7�w��7�:�
7J�sgU�Sr� ���I��5��v�.=��72�U:WyF�bv���x*6pB�^N��5�Fgz�+!�$��͚ۦ�e�1���rM�ͥ����S]�1G��w���>�٧%�B�BY�Nh3n8����c��]�ET踜g)WZbm��d�aiޣW��󗢯r����,F��%�ou$�bC|36����#�~X��j؏��+��{�a5���E* K���&�Ce-ٓ /Yx77%nC5���ǃ� �Rf�����­]�hk��g�� ]MJg5�S;hfkv�O���B��[��Т�T]f��yU|%���9���M����*|����Zp,��^!R�h�\�MmC.��M
P���z��D�z�˛�W�CKH�8I��3��Sg�z��6��u�,�PK�T��N�Y�%����|Ɂ��cLQU]�]��h�]X�>Ts�Fa�d��_��|q��m�I��DT�D�79}r��=�-��֕<����(=QoX��g�V����J�zˊX0q�di�Э�5rT <T+9�pBou��N��"���l����lZ;-" �;�Z��R�pqs��&XLAiT�6e��p\oo[#z4�6�46�6�`бX��phۼ��ۦ	�\���VX���쨘�/�5�Ǌ`VN�b�Ś2q�ƻQ$�iX1�F#J!�h�Q��<�9q�ʙ�1�4�ʛ�K��[���4�u�JK�Z��wa:+=e��B �6�[��u�����.��.�e7��lZ��v�����h�S��;����jZ����F�k-��w�z��������=�'Wc�e�̬�6jis��õ;�pv�j�0�܈�z�|�0�Zx)����ҭՐ��:R�be�W t��<���l&���\Ԙ�w�=��d\B���r(u-��TXz�+.>p�}��P<���0����J浫�:��a�g.p�&��E��Wp�l=7������*�$y��2�.�:"�Ϡ{.+��V��O
���խ�a�_]�D^d�o�}V�ˍB��VP,��׬�2L���r�o�&F���;���7�Q�U�bTW���W=w�ju���sh���ܙ@���|ɷ[�=3ٶ�nmQ�9��fF`KR�sm�������#��[Ů�W&�mc��&�KL��%`ǙV���z���S�5��=��3�f��6�iγ�2gV@Cݿ(�V�7y��n3���D�=Bיǣ{*0�jo�V%�Zɴ=}�N�S��QZ���mr�ڜ�=Z�x�p���93���E�$���u{�֜Oixؽ9˨������-�� �Ls$�<�3m�ehѦe$�Yik��dqG'or��B�gqK�)�6���ik��H��Z^^_Q�[Ki�l�T��.v�}�<�C�Zs���5V���LR�^O�Q+U]H�|�Jt������M�#�Ř���d���%o����\!�$����}A�q�rN�L�$���ͼ�s�d���/��av��wz�@C	�ov-e�#��� ��BP���"�mQ"��-���9���%	n.]=|4bx��ڷU�/�n��r+����W�*���U�j��Kuڷ�F0���.���t=51)vJ�[:%�v���z�FJ�f��rӵ*e���ԟ^V2c�w�{8�V��K��t�=4����!e�Ft�x_�an�ӱ�޾�Ha;�F��6�����\lz��}����4�P{vC���Zc�H��Z8Yո@��Pf_%t���Z��q-:�'/[yk�1Ԟ��g2C�3�Y�Ir�8u��gn�B4���%jt�b�Al���ܽ�G��W�Ŧ1x2^�X� �tX�9ePX��'�e��
y}U]>��;bKa�e���wm}��ƚR��&�
�s�8�:Ϩ]�0����׃�&�+ ʎ1�i�Zj�����̼
����v��y�U
�.��$#ő��/'e�a\��gm*aa�ں�v����ug]�1�#��g,CP��]���^���{�������P U��?������/���ֿzo����8���G���-�7���S�x��P��ҷS12�%����@I E2�2p�`��d����J �%Pa�cLH�-��#�0\"
-��Xd����z|��x�}��Z�P5�E�'D@Y����A��uTQ ���M%T��6����CQ�L��ԅQ��!"����A��I2
���h8��S:�%J���R �K�Ĕk*���܊�e��n��2�i �1躄����IQ�0'P*5LDAp��'C�(�Q6��`�8���J���x~PXѮ����'�n��-���������b]����J�w|l���g�T�wJ��;���]��;��ʂ��އ�"��PKʵ�賌@��Ǡ�W&Y��mD��q�<���z7,��7�k�Zt�b�Mʟ0 0�����z�������yr�wu\�z��L� ����)e�<t_gn_	�AsU��aD�g�5P`���Wz��l�u�F�M�Ӯ�!)}i_�{mЁꇦ�橕��x6��k��圵�Z��=���y�8�n��3f�T��'c�7u�v�rMP��E|��~N`�M+���Vd�;���njN��S���oT\��nP|F1(t�X��es�p>�W5\��nw�:����Ά�hv9�X�6;S��k���mM{��M@�r�^* �D���j�SP �=y7�����R_YӝOM���k36�����r�)$+�FŞP�ۻ��h��!��C�p��*pf�i�g�]�M�9�zQӦ֦����w�����;.:c�#�䲐}ap�KD�ٲ�:ܮ�wgw�g63fFn�d�넸�������fj�m���kk'V[O�ji���ۙ��ˮ��S'��t��b�LS����I�U2�g�#R@�^���{��w��{�s��s]����hBS�3�rX%
H��l>3P�ܷ����NÉ� ,2�,�Tm�ȣ$2���$D9!e*P�i4_n@��l\�k��S00�!�RC"0H�H��L$J8�m58�L&T>�t4�����Ǒ��'�.AS�$�HȒ�ܦ9E5ĩ1i)�8�(I. �f�C,�˅��Q&,�l@�M&R$�d�&�	�ը���u Ap�ʍHH0�$ �%����I��H�b!�I�#IC��(�H�Q�F&�p�J� ���ځ0�I�[MF{�����O�n���M�I���|��(�p��i�%��14C�T4����$�,�Uv�")�l�Q����L1`�\|aD�K�#�T�1P�����A%��h�J,F[hH�	�q��@�Z�X���e�Q�$-�r	�@ a��J"����"[0 �
@�L�Z�X���z��$˨��K"A�PU�ӝ-4��Y���v��u�㣮�뮺��Y�]u׭�����o��а�����#"fal�2��O7Z"uNj&r�B+!"�e��u�{~��������]u�]u�]u�]zzzz�����;���}��$���bZ툑��s"�����|�����
(�-�y�r"(>��	�n�*�0�l�JN�s��W˟{��fQQNI�B>W�\��+"�;�]b��+V��#�4O�嫐�����YIuB����d*���^8��
P�N������^�Urt����F��><ߝ���g4婔l��9�W����s������㢭*(�J/�����QzĜ=�R)�qw=�Ru�;��y�0��e�EGv=r �w��кZZ��L��MJ�ݷ蝏����uXnE��*���Y;h��ݦz�9"��x6�v�EDm��w^��8�88x��(��;����oⱾws�3ܗ��q����B�H�mF1"	O�fN'ώ�/�G	�w��+�㊫�sD��	2J+�� sx=���eV�pWW�:p�K������0V�
��9sMs��{XJ�ە4�ZR�ã^�v�0�咚��H�M�(�h��Q'P!
��JD\-��H!��`�9#r8
EN)�m�n�`��j4\I�،�"��&)@\��
N ��K�d{�竪{�u����wc�𻠏mˠ5vjв��W9�{�J�D��;CV�d��t5�)�ޥk5�M��~�쿤�_Wge�"N-6y�_v��ycܮ�f�3��O�D�w�H�m#������Tq�;w��lP�|�w-Z�+,�����A�sh��,���lwWq����L��WD�C=<]�U�Gvcu�/|��Z���5��ʾ���W{����W����.^5�"�}o����^���tU2/���l�r��B��4����b�1�dgtM��^���K�gw��Y�wUs3v� GQ�xz���-���w��; /5_t|�~�Pfyz^r�M�{���A�t>�y��O�o�1�����#{oz�XM��k����V�^�k�G����|p�U��4x0�:}%����]Wwt�����7�.�uċ��2��{��w:��Y�|ޡ��pGs�qu;�݄���!��v��Mi����o��h輾T�t�*˂wn]���`�徻/e:�B�U+ro>�Mq�\'�{���-szz�������ɥ@(�Z�_$�xؒ��;#�=�Q���Vn���eu�['q�ȯ7��s{��jv���|>rőq�����jǴ=r�J�.�����=������P�7�{�o���Fd�7�b�L���u�;����7����G  绸_H�wg�s:]J-9��/������C�qn��;�:�,Ȭz��v��;�=3d���ܙ����q�w���d�u�}�/M��8V�r^tX�~o�N����u?o�V�ͫ2�.�%W������'��}g-,��S}��ӗf3=U�Q�ok�����{��aT����͗°�Ib�ݸ{�����6
ݭ��8��?�b�����W��ooeڧ�\݋��_>��z�vx,��}r�!������ѧp�wgF5���C��}���������=����b���}v����/��n���>v��U����g@ncvv3ǭ���Ӧ�����?a^��\u�d���o�,��CJ!lӬèTk>�c$��G�G����V-��B�&Ð�jc7���3u�-l iׅ>���ò�M\8f%��m���ӀQ�q�F\|��{�}�6=��(ۋFj�`��G5��&�E/�ʡ��|{&�}�u	\`���غ;<�+������4%�9�^�Oas��3��ǡ�zb�Df|p����ܰ��5�c�lf_7���{ޓ�*m��ϟ�v�'�L�K�B��N'}*��;sd����KL����7>��}�7�F�����m!�s�e��=님�|˱03�&{	����>��}��crV0r��g�����G�#�pX����Y�����^�A 䓱�T���u�b��!2{��<�ҝW�=���T�%�/�
��/�'}4t[=w�oǜ���rO's�=�OۀT��e�s|���q����꿧�9�.���Ǭ��<�;g[�����5���^2}�����0��=-h�s�]f;e��ﮂnތ��͝�@gh��}����:��F��rKϮ}�5g	
�?=ۘ��͋���;{����u�������+9�>��:��m�ޙ�ɭ�K	txN
�r��t:�V�'�n��Z{&V��¼)f���6�$����*��T�"��=]4�SD�y�ytΙF�_N^��`��P����r�y~�l�ǅ{��O����6�Ok��PN� ��HC9['.�'�s��ӽ�\�����v{j�ݙ]mMF�S��e�I��f�T�^��d�-0Qx����h]��������z|��M��/ѹ��s���2��Ol�$��}�eu�9WMI���P�{�Bg����������y���O�߄��H���]�A�*A�J�o����c�;�[0޶�;E��'o:M�Od�GQ���9�<������~��{o���k�^�����<n�����-�mo����mt���\?hb3��r"#f�����cޮͪx�^�M{�e�}����办��sD��%t{���(�a�Vw��5$�7<Mtnx�f��+>Ö�zr5��Nt��un�Ƽ���=~���.|klI��s�$�Sw7wMa�gb<V����V�I}��{[Ҵk#��Ye�Me^�-J�)w�m���3�3]׷�4"�<��$�(���D�ɒ�QF�������P�Hք��^��
T<�V��o�����;{ܥ��B.��^��qr7[	W}�;hV���v�n�[�[�O9�K%˸�eC��	g4V���0yp�\���
�mn�����WԌ��U�6�q@�����3������f�?i���o��S@�w�9���P��$7l)�H'��f�oN�o�:�@8*<ϣhX#�[��S�����E�bQsط2{7���Փ��\'x��e7�F�U��5��;��c��{⧪y����f�<�>p5���m��J�z{�f�V)�2<2X�������[�wz��Y�x
ޑlf��;�!���tq��0;���i�l�z��h��?��@�&��8���A�c���O�a������Fq��x_.�����f��rߞ��{ӕ�^�K���o.�`�5��=����/I�%�ER�S�i�o�g3��ɖR��g��������Pw.ۈKW��i�xvG�%�z��wG��=�v�ve�͐�Ø���$���JAd�kF�Խv��ld�zQ�e��S��75Э�b���46���mB��	)��y����X���/,�k�g�|淚O�"p�:���|�V,9������_Q1��";���)ďWE�:�nU�O���}���3�w��펟W�m���5�C����@�tW�{�>������F�i��}T]u���mwow�a�ߟ=Đ���z���M��l~�F����8P!{C��#˄ml���~c���)��ݹ�W��ZTa���Zߡ��.��U	&yd���>�Ϩ.��s��mni�,+%��Z��v�w�>}Ѽ��'���l�2����X4���Z��}s�F�|���6��C�ͥ�.s=�{�,�K�㭘�g������`<uu��5�yr�ofѮ���� _���t�A�%���g�`����~<��/��mE���gc���,�|��g����~��=�/O����S1oR7�]ݜ�Ǻ�ڢ᪳��>��@S���v����m����-�ng����l���^��/�D�z��o��VqGxp�z��u�5�4�%��@��B_�Sg�u���t#P��Ů����_\�mR:'8"b���;�DUS����7Ҹ��%�=��������3n�*=rX���7�G���Sew����l��0�缎w���o�e�]��A֕����}�:t�r��5 H<�d��]�x�|>S�*R�yxo�c��>����[_TҴ��{{j�����8�� �)pOzN{*�;�g��-{�����Y�'�%s�w����"wO=�Lc����wwU>��~�|�\��h��75�u�YD�O?�Ot��3��C���8�C|}�t]ﶨ�kF;h_���t��p�@�UJde?e�z=�=�jz���zy�f����zd��'���uz#�,�<���d^�9{�v�2�߸�/Gܟ�,~� ��k�?��Q>��o�v�ۚ�l���~�;_e�������p}hsx��=^_�տo��N�mdg���;WI�E�yvU�I�+�ʯ����yA���jW��;�m{
�������>����(��q�|b�2p'p���^��x��m��ñ�5UB�U���ע�:��8�m�[�dި�:�n�x�BW+*FM]�\�gb�}�i${.L��1�I3|�^�����,/#�t�R�:��u��w<��vu荃���l�)ھ�b�|||�:�/�o6
d��h������6����Z�2gN��[ޮ�/�n�9��'6����a/
�O4���"�b�������;�:�Ogo�5��/���j��g��Mm�o"��n���q������w�rt�Qù�H={X+���o��tf�C�w4�W��pq������-��m��]�+ך�GOq��|rn)�C�W�+j����7�D���rs����{��=g��l��'���O&L�۹٧�3E�Q�xFd�r9=l�r�X7�<_�c
��G%����:G0� t�wUQj��8S���y��W���֟W���� ha��݈��ݍ�ݷ�Fl��"����s���׃t�G��CԥQ�+=���;�{���t�d�ooE��oo�2sݜ�:��������̹�b��;������i�}ozs��P�z�m�E!�-���tP���H����U�K{~C��m��ǲ$�����R���F>f�	yf�S�����-�q��!���#::��f���]IU�EǼ8�*���7��ۺ��'C�/!�U^Ҭ�
�:�J^�wvW_̟����� �hr�ӂ�Yp�����=u�P��g����vͰz����Q�_Ik5��;e��.�����\�����O�ޓ`����}�B��/�G�OhJ����V%����Ґ�R���d�ƙK��牪:O�o{}�Ǟ�P�����=y���s�x@�'�h{�!�v���]��&0��_9�q�ƝR[��3ܗ4hТ�z��뮡��]x�+f�{�[�s�v�|��43�{Ѽ{��}ϧhk�<5���V��G�,z�S���U^ћ�T�;��D���C�S�y�w������o�b�:��,xk|�$V�������l{�O�.N������bb��~��d���;��W�Y����w�x�6l}w�*̀n��[�l��_���"����g�����;�rv�̳�^oӆ[����ol;�Y�-�4uP��{����۽/1�t��Hn���T�G��#?�X����lj�gt>z�HآoCɕwN�<5g�/ ��V+�:hz��FBl�B<���YY���ã����y���Q1O�)l�9vY[e�������v&ɚ��Y���o������w9ۏ�2�����M3�����]�;wd�]�a����:*ߨTlK�����׮͚��yW�3��C���G��/�P��;v���Wx)�����(̞��K�U��g5�ev�Owt���Z��@�@{�vЌ���������q���=�t7^����=͵���:MG�y�;G�=���m��|$���o�Ix���s�~��g+�����g��{�=<fW����&y�i^x�g��<+`�L���mwn�/�پsד�g��q3{��~��O.Mur$��������7�5��":�l�w�k���T��o�>=�޾���{�� 
>O�Zǆ����LL �_=\O��j��������ؙ^�]6]�:��}]��@�� ]�"/bj�{�7�l��9쾡�y���33�d��	�E��X�`��xx�1��ö?=Jh���ؚ�m��p �y+w��W�'=k�trN�-�I��]���S˔�0��1����ev��[`���/����h�V��Y���`S�=GY[Fe��|�Ue�_Q�q�J���|8vV��1�����RzZf�g#N���@�w�&��z媱H.o�q��zʗ{��L�l-|��7�9�W\������^2Z������$��;�[T<0GM<�N���pa�V5:Y9�q�j�D�.s���Iۊ���O��G�7Տњ�;J���_U���b�ڧ��j�}��E;n:�ko�{�[�ۖ!y��m���{��P�!���OoF೨��v<�l�RMeL�k\��d����=���D=�)҅����y���yYו�p�9;�f�9���V�a�I�p���PPT���]۵jT���)�z� �[��z���B�\v�܄r��+���T�o,Ik'4�_|��jȃ��W�^�[>�;���ڗN�˛5����_t�wg��a�$	��/U�ò�ܞ���J�-2��{�΍I���w[ٖHn9f�M�u}
Ս���/14�up���Vt5�k-�V3@u��$#\�s1��岕�0�1wC�}���d���]��=B�)�W�jH��n���[�M2�e�}��ⵜ6:ё����Z�إK�ڣ���m������,�a��9r�#�[oO#-���mْ�4�$���_�V�I�D�l�[�i3F�]�`)g﫾^�ؚ���cذ�_z��;O��B�� tM���>F꯶�j����l����+19Z�,B���\�Z���:؏&�x�XȢ���NՏ�S*ʿoTxxr�#��N;1���ik���4f�ȓ�2�q��u�Qkk3n�h�Z���8�mQ6cZ8"I���B]-�;O_7ٰ�,ޫ��&�}Kج�+�J����q�~ά�q̺�X���ƛ@�y[s2�N�0US{���:(V��\�n��a�0M��q�W��]v+������`���TW\S�u�h�y+V�X$l�p�X�����ܸFƮ�:nN���
�KfvnD�ۺ�)v����=�:[YrM�Jc�QЌ�k�ػ��j�36�n[7��T�#��ͨ�!�WwICs>A�r� /^�R�o��01��]'��u�MSX�R�r��<�x켬�㔳5��@�L�Z�*������vK��w����ݤYJ�ݾ�Y�km=Z��_L��٭����x�V�|L&��4�:95���n-�y����i��-��p���,�w�b�����ԑ௄�^O�K�'r鉛�|mTY��ޥ�gv����=.������3:���:$ӝ��*�wwWP]	�a/�+ ��������KaXfdC]ŔW�wz��K�[�dD=��I�=>�|݁%����	8�Y+ܝ��NK8eY˕3==>���~>>:��Ϗ���뮿u�^<x���{�s!"D~������'KHf�����&ILR�޷8M�������f��=�%a]ơ^z��=vOLO��P���m`���{������v��>�ߏ�������>>>>>>>:�tu�]x���_��Y�x��0Ȫ��Ī����r��Oy�zQ˛'���X�3������_/q�#\��^��v�]������'v$�EC����-�%a�s�*��ݸ~tw�[}���9Y�َ��Q[	�� ��](�~*����h��>*<�t��y��D��DDN�}�z!F\��$�"*�P��'�D�x�C��;{'Wd���(�.V"UG�('f2�w��'�}	��.��E��eO�DTE�K�J���&�Ͻ˗̞d���^�9TS.���F�׏���H�TU$��>;�`�[���u�qp�<�)n_�v�\��L��Μ���Dߞ�n�(�)G��I��	!f*����u�rI��/ށAN�U(�"��#!0��v�{�s<�R�~F�_)����Y�ק���.�H��{�׹yP�}��,�o��MN���[�h����ǟ������j�J�f�p�����.�u��9V��[��@W|���ԌX-rct�� ���e�n��z�uN�=a�2.1���z��z�컣B+vy�W+��<�-��I�a��16�P`���/1F����P ��8>tX�
������vy��xD�ϩ�T+�c�&�{�[����"+&
��H�a�����{�mL�`Kyڃ
ea��b�Ҟ�wh���S����r��M+��XP�O8��me�16�;ޝ�.o�U�Ui�U�P�|��x.}8��d��&�%�-WWGe=|b������H	Y'��i��R�'6��Y_��ZL|����/q�d���k�V��i�����G�O�1̓��JuiH�U�&��ﶅx�d:�=��{ի�d��Y�כ��P�q�����`>�;pa��RO�ИVT������z���r��K)({b�$�� ��}KH�w����~5������������n9e/��-9�e>�"q�#�QΡCS�wU���8�=o����g8g�s�����5ô7xU�7���L�z�i����N���Z�"�}��\mOM����C�����u��_F�9]�2����ǵ����,�Ԇ�5�kQ��j)wV�V+��r�E9����a�K�/�l��#9t�gr��]��oc4��C���?�͸{w3����s�k�^�=x��9��@���Be���_�	��#�J������R��C�r-��4��}�:�x���L˾�B�U�	����=��5?n^�m_!�ǈ���*�@L7�����c����9�-d	ĸ��� ��}g��%���Ͳ��li`��=K��Fײdd�����<x�0�� v�u�w7y��0o;��`�[���8�<zV�
?0�oǖ|yq���z��ߨn��67��d�[�p�:�m-�fT������� C�?��^}���Z��?��~iomV�?I��]��#.ۧ�k��j�F�^�(y��!�P�?��>5��KO�2WG�����,���q�:/�����н~�9��x����	��I\���z���8n��e|��o��Ly
�����q�T��~�v�6��J��ݮK�,0���j��%>��z�8�E�T?V�5i��DE�k����k.���!��!	�l���{@}�c߻�2�]B��UsxSW�\[H�vb�|�?����>�_�
:�sF������K/
����z�S�+�yφ�R��Х�o�X:GL�Uu1֤H�53�T/�`��fd�|����ņg,io|6�X����7�M4�@�ѵiM8*x�'�d�K��\�_C���ȭ{:��_��y��vv�e�S7�o�Ȕ���ʮ��$�u�:"�ѣC.�Ь���Y��0��$Z/��}<|�����Z�!1m���w8�%��="����Erѱ;n�p��ҳ�Nf!����b��F1����dܜg�:�*5�i܏�5J�,e �L�p:.
�p���=���}�x��lYۗ�!ޢn�"���@#'0��>���,���n!���@CU[�73�&��)aE��u��m<�	�o<�� I}�ڼ��0X��2׆6����}a���~�ć�|���2��k
����P�[&�kJ9��U'���F�><��ly����/���c�[7����k�^��ꀞ�PU����ܫ�PY�4�°+�\T=��꤀}@�|dvX����_�m����ؠ=���G1�LG�о�
T�����p;��{J;��K�����Y�3�7d>�٨X���!���*�0{�gɹ�Y�=S�'�~��5 ��c��k�t	��A��s{�m��u�j�o�@����	Z>u����!��K�ր��$�[�Y�)��=�tz�i1Z�ϐ���s���q��H�"ڨ��:��8�s�<���q�9ʧF�ى��՜ݐ��O&	��A9}7w8Z���:EZv���rWY:{�L4.N{�@��[��S*�um�|��	��;h-Ƥ�y]��7�*�5,ٻ9�o:R���-��Ѵ��p=Wy󬎖�<���W�8eΥ�򷻺F®���y..]yY���y�a$}��ؚ� �@P��C������3�:���@�;ю��2���<�d����w�����t%�8��{hq��^�O\�BT���o��=C�ז~6J4�9@7�g����iC����� �n&.�წ>��[�����WAW��oc7��f�03���0#J�K��6P���9��S��CG4�q�s�%@f��}�ɮ�	�]B��D����ٓU�_8�����f8-��E=��L�F�k�qL��������ӭ^}� sf��U<�i2U��q��zy���J�8Ms+�o ��Y_)J�p!e�����<���6�.���e�n[��xy��t�Z�KIP�2���Oa�U亓x1z.�!>�\8��-�0Z�k����Jg�]��ڼ6�jA+'�䘮t���ΰ1�`-�u�����������6�=du��-����n����^pDsm	��ͩ�4�Ĝ�2����� suy�)xjN%��쨦؈�J��\uAj����l�R@ψx�i�|_;U9�����.�r�����SIP%�@����}ڼΜ�i�j�S�75��n��z��ӭ�j����3u�mW�z%qr<�c�ӒE��CuD!��2+�Yg�ݵ����D΅�%ǹ��ft]�o��*�ݾח9�+���c�h3V��rtY7&n�؄=�8���צ{z�������?EI<������@���8u�[�/-��ȖR6c�E�* E�h2����������+O�����f�,��䀂���������ٲޏz)�� ͭa��ڽH{:���_s�-|���X��xg=�8'5P(��	C���/�1���O@��4��h�g��n��UN]v�g!�f�)@f0�y>�x���Dx�M�={D�������+�[ú_�L��%q'/36���郒�*��~�� -�;�^2��!3�T=�Ǡ�z�Fs��A��[����9Mz�J��4����{�xCG�(,�ǿ,�jZ��Xȏ��:
���>���
�w�V��A˺9vj�4s]N��W��jZfb�gC���o�ڿ���ז�щ*f82�d`c��NƔ�Z����,3��!�YA�4	���l�"�X�Ur���}�Q��;#�B����|�nU�n��n����P��xpϢ�� �p2j����t[�?�f=��z%�-ٝ��Kx[y�quY1y[Ts��iC�9��2ss��%�{	t�+�>L*�����E�t���ޱ#�M^F�v~+I� ��⡂w.[�52�l�{���{}j�`�g��������˗�i�=�Gt��n1�������t��ٖ�l�O�-y5d���ĴL�����5��f����#XP^��$��wN�|ע�c���z}�����?aX�o�-��>�L���!''�ӘL���JuiH�Q�IZlk��$kd`K�\�Ü)9����j(y��E�֘&C��7Q�:}�&*@I��&�?�c�BW�X*vqs(��R�^!��ng3�`����-|Lc�<>\���(��r[϶�7 ������?'���Y�:�6��p!�:�e��!:a��8�}!�7��s�E>/C������e�|D|v#z��cx3�vef,���Qx́����{�*.��⒝VQ|:�Bڑ��DxF���W弲��nr��{'h���JN9��rz�r=U#7�3]�=�K�T�6�U�5*���[���U�|91��8jR-�wJ�|"��{}@k�FV����7�NmqP��ekήW0�l��`�r�1w>�i~��XJ��C��;�MM"2OR�_&Ԍ܄���sߍ[�8׷���soͱ��8D6�U7%n�ɯa�x�e��ҏ�y���:�yd��!��{r(P&'��sS�VtE��J�y�8����g���@{�<I�e��ސ#���ߗ���]ѡZ�(z��f��ە6�i�r�C�ت����� �|/M����షƞc��n���������-ŝV�>���QK�]�s���w0����>,�j�*�e1��[��&�������_A5���d�Efr�))α�TXp�5X�g4�4Pf��{�����=�@ޓ����}-��ꬎ͛&���{CGV�h=5�y�٥����F�<МEہ�b��pjߔ�JrׯE��:��Hf�t	��[��\��zz1طuV�Пh�nI��ū��fnnU  �׳o�U����zw�c�Xe��'��E�I�/��l�҇��kь�usmTr|ka��P%���K�;WGc���L0��&��!�B���lE�Ź�Xw�<��O>fɲ�%��q���3�#d�Z�;�қ�t�\%RaM^G'�0�	��+:p����="qó5z�)�8��oB��q>���F��w	���w8�<'I���Q��a�l�_	�=��\#gzhX�z$8��8�~�TkӸdI2�2Y�2v:�_���R���z}>��ܸ�E�wwP��睄������"��ƾ�z�����k�
xfn:z\u�7K�C���p�̜��I��>��<ɖ����h�k0h�/��!���"�i'l���	�^��o���~�rV�J@T����|�e&G$^Z��r��Q���UCx&wq��n�6ԧ�Ycq	i�9�{�kB[��_=J 6%H�����ʹ� ��eV�����k%�޳�L�ƌճ�uW���<Ӛu�GP54�j���q灈2�_�s��=g2�]�)r���0a^A�=� X�BY���]a@�����;:{e�J��Mu��􌹎� ��ŝ�y���3��U�)�ۜ����=��@����|�y+(���{k������}~��|1O�e �O8�0��Kғ�y�ܵy� i����Z��lR6��� �B���}�:�gl�@|N��حѕ�H�ޡ�9�x�׊���j���v����\D�+~�]>�+��
{F�J�0��0}��#'@�s:,m�+S<[`�V�����d�r$�����[�{�g�:><�B��R|=^H��W��e�'9х%ٟ����;߇�S JY��)�}�#�ʟ@�ǌ;L�xn�^Hf��@�N$ō��/�������2�7h.；��Wؠr�R���z����Z�=�3j���{R�&��v�3���JG0!�8�sE��	lĤ,{]�H�`PT��0�Z�2�q��$�^/���a�}���E0>Y���|��QV@,�n�	�x�U�V��V�]���[����Ù�6=I�.p{��Z�L�J�,xy�HN&|�;�)��mN�#Q�(Cm[4#ݥ_X�mׂ�����)F�c�S:yjo;`����|����ԝ׍��V�2���cqV��8ygL���I��R�����-:
��������)�|m!�A �O�>[+¾�y�����y�\���m���"�/��^4��b�^C6lGNYtũ�y��f��{M�NA�{;�b`F����g�  z=�=�{֣zt��C�X�Z"[��8|s��̔�}��L���~�-�JS�~B��~U��1�/��?�~�=Ļ�jr�Cŵ�7���7!q�����b���W:���ޖ�]����^�eӳ�k�u�;��)k;7��`�^��!����o�y�"S��f�@�Q��(��%܌(x�|�{�ZXʃ$�����@�u��_=���Z����M�r�}��� ��ZX6F�]/^Y�Mܨ�hy�7׉O�;k���l�Cϧb_�9t2���%\�D��m5����2	�,�6KX�CR��^e���d�n=~��y/���u�p uT���l���>�!����4qi��{j��zVȇv|�l�ܛ�if>�]3����<����&*����m�9�
��M�\��y���啱{Jٮ��"oOˢ���:-�U�_p��ݿt���m^YX��?��1��?L�}��`��ZH�Tx<j|?G�z���ܨd��9@[m�\�;���N��)ǵCT�H��Ufa������~^�yxxe�.�>4"����v�8��mCvy�7���B�O9�b&�-�/��]\�¶�5�@U�:��C�� 9��;���c���C�v�X�d6�ꊲ��9��ƍ��u���C��D��}�]%@ֳghp�ִ�-9ٹ�_:��'o��3��p��6�1nr�k�Ï�KY{�jl>�� |<}���G���xx%�o�壨x�۸�z>���������D �~��n�^k�WiE�Tiߖ҂粨���=\���6�[�z��zFN����|���C�X�F@� ��Ql8�я��M�-�Y)[�C�3ϗm�\�t����<'ЗN0��0z�oո���v|��w{e�w6#w�]��x��u��zb��u�>�	�wD�/it�(J|'|����t���2�)r4��"'���Qᳺx{�\��ИL��"Nw�sߟ��'nxN�S�L�-���#�d�i�C�-��T�t��헨y^����!�r��X)ܓ$�[�'טM��ȤE��W�kYQ�q{a���t�k�����=�FA��:ׁ�Aun_�`��e/o�=Mu)z�;Z�l�O<s� �-!n{��W���@&+��D�A>���5������ſ`b�K׬��7�Z�
�⇫���y�H��z���ԇ�JuYD1�����E��i�d�0ö��ܞ�oj�!�å�L	e>Rk����7�
IOs�s�U#(lZ\uW��8�888 B�׆�n���?N'YR���ͧR���f�B�J��٧X�rM�X�vK��7q�چ�0�#WY���#O0S�u��]��Oͷ���P�ε�1MWу.b]�Í�mYM-�Wo�����v$��	ƛ����X�a=�8G'C��l)��v�lї���V��� �Y���A�A�v�,���ǌi�=����1-��b���T�q7u���Ntu��7��o�TviB��Q2I�ǩ:�,�I�N�����p�f7qN�R[ۻ}yx��B�u,UE�*�R�i`3���뱡4�7�do����4F�UKh�o$��vb�+��ת�RR�h�v\��nNR�9״Y���.Ҹf�z힍��桻�C�|�Y�M5ӈ�5� ��]���yZ˷�d���M��lk{��9�;v�l�HfٺP�3�ԛ��/m���	r�̡�e���Cip�ܸ��˻�
�8V��u�u4��.���XbٹJ�˝"֛�x�fV�ku�b4��Y5n.����>0��V�c���+y�|��.[y��r��R��\L��:)��(�^1�w_<�A�N}%��:���9���.12:�.�v�.��sl8P��+����ӫ��� �/h^�F))uo�M�F��m�{�x�:з�e3w�8�*2��f/Dw�b��K�ݛ�'�F{R�Xwsͺ#�S��
�	�`�.Y!��/%�L���\��ܫ2!Xh*����49P2��c�	T�2| �ެ�J���$4L�;�8�����8e�/\�*T��RuBm�w2UA����W��'�20�q��]�b���w�
Z��K��Ђݫ+5:t7���Ol��]���Km&�x�i���
�F�7�f�2��A�V/a9CU�]I+�yئ�����j!�Ɖ"�b���]�JE!T�X�r���ح=�z`��:�����2�PYt\kh9.�%gvq�>N�Mq�*M����Y=B�^��;�{�5<�v2��z�I�75�����I%(�si�VK8f�mu��X�pZf:U2�_e�8���WX��VpC/�S����lZN9T�l_�̆��d�FC����1�����S���wp$�㌣�NwB���|�r��/�q Eq2﷭�Kb����m]�s��{v���s!!:D>�X6
��ad�hdV]NX]Ribȹ)CǺi�)s�uu����&������4H�ÜR��Z��ݰ=�y�%%m�_V�v-����®���+�-�{�T�V�Z�l\��3b�}��bu�b��V�T�U����'�w|=��_���r9�-u7*���J��M�
ݹ�4nXuH���!�5�Ґ��r_Q�ӝ�5'wu�]���������|�G���EBY��(�5�wJu ��p���k*�2J"���8���������]q�������������<x���=�@QO����Ɠ�*��
쯬�ա���f8�R�?ǏO�������]q�]u�_������Ǐ>?{���".PQWEa��2�/R�^d�t�"������A�
��B���䈲�B*�(���ʨ��?=w�p���Vp�	_^7D����8W8_R"9EUUs�"C���E\9�Fd���΄��#;:��Bv2s��U ���"Ν�99I,3�Z�"����7-KP�ٙMP�(|��UQQɔQK��=.*%E�t���.�D�r�����r�Z!�
,�.d��
B�*�w!�A�\-��*"�uB3�Ų��Ƞ�L���8PTL��"��RO��w��ȹA�����D�N&Mw��]���.*SמȺ'J9Tw�p�T:�Q.�IɔI�wѕ��8NJ�����|\B����$�Q����i9��qr״sφ��^w��}��޽)I�$%"f����ى�Wf
b�t��n�bs8�fjw+�w��1�°�|z�d܍WI��[� S��6�cZ���3���rU���"�#������z���޷��N��`�/q����S��%OuϹc�<��w��嫑�p�Ԑ��E��a���"!�\L��-�d㈰��pps�W:�1�<x�B���׽��<����ۭSZ[�''|�}��n�E�A#p����НU���i6���"�'W�a��O���ZFiZy|?b�o�9U���-s H�|}���}'�Ф�Gsx�,��`�� ɝ�o>K�>O���I���f�Wp���%��DW���.���C��NYZ�`oC	.*���C���$e�)�|@���|+�N_P�by�J`<w]:����:���HѬX�����U��>�Ư��,`� Y��{��?_�<�w���� P�ʐ݊��}�x�-b�^�T��j���z#=�<=�])i�z��WG�����zye�%��irn����m�=����d��+ �������^K���b�`0-�<��x����c�����J��8P�S0}.�9���	��%AO�x`ըʒ������8���~�ΪJ�[[9g��!�oe���D�B�q@<����)ŕ��Z��&T-u
��sz<ŭ�jc'���f�w���ݟ���9�e1������JO�8`�'=�C���w=����Р����V-��8���B:s�����o�ׅ�C'O
����{���Lϊ�!�����3�nq�2��;b�,+!�Y��.�\��E.@`��6����]굷�Ĕ;�����mɯ�VCc��c�ji�Y��W�$͵�mmDp_g.�����vh���̉N���x�(;�}���V9��]�^��;�����n��Y꾕��ϧ���y��{�xk�ps<�R�.���� ��������R]�)�Yz�]�0�f@�cH�I�Lxp/WlB��4��Y1��{��,!���i;�I> �Sg8	��y@q�/A����� �c���6��v�:\�Cٷ��d;�8i�R�E��J���;=o-�P���=�0�'�q��tR�k�QQ7U�:�3gv�[xj�`��b�!1�y���I���<�^�ߟ�,�Úض�i~���.j�Nڬ�� ��p��1n�:n�LQf�Vݞ��V�I�9���Z]?��I�ώ��B��ά�E��%n9a7Q��I{#'�xc�8�����Ph��9S��#q*�	HYU5qQ]u�N����q�����&���������P�`��>��8�o���'�ڞ�Q���y����%c3vv�7���[揱W9�0����y{J�TH�P��΋�����ɭEso>0^P��oqQ�̿P%��H�oK��hki�ǡ��8f��hM^�������!h}��| Pm����ThZ��������r��,��4�t��i�wH�ֿ9D���uT1�W���Dv?m�d;�PR�'5���TNm�Y����3oW*�c�z����J3d�Ũ����'�,�^GĂ>"����b�v-.oL��7u�mNbCE�XM�o4��y3fǱq��ܔ�Σ6��B�\S����f�������O�~�*�<g� {�βuab�����ENUES8`�3�-Ο�(U��P�/|��s��� �T_R�mW�Cu�O�qLN�:�;ˬ�C�z���#���.-<�5QLt1e���o�i/I�?���w�)� �e����PםkI�;Z������"u�N��N��,������|ǟ'4.�Y	=��}[�;����d� ���p:��0L�)�6s����i�x����]��,�*�/���ٙ���}���Ԁ-��tG��U��3) ��Y+�a9�,H�5m&^������3��M
u�P��V�����Aa~ׇ��b����O�t��T�u�b�Rޠhtv?0P���O�p&2Ne��x�b���9����mzc��͙��'q':L�{� ��%�m|tie6��'�s�<�W�X�>��|�^=��t<,4����m�ӭoܫ����m�qE*�'6I�z��~�@oX���i�}��x�����E�&%�Der�dl��j��=|�ֶنx�O��O��|��:��c�2c��lx)� ����:����lt�[��ᔞ����%�s�j�ɳ|z����6��Z�xWv��s���smݺ=O��]s_"H���0�=}�Fh<����:�dZE�>�G�a��L���n��tz@�X�gFcp:Ή��2�
���� �9���ϸ����x�AQ�μ�wן]���O�ں�>��n�=CK>�7��^�~��7"K�gc;Ϡ��FK�����Jf�WW!��t�k�⨏˧�w��o�,�����C�{�
'�T<g/X(�w�^q���s�uvga:���>C�l#�f��	|>t�l�6��a C�;����< t��S�ir\D�Wz��o���[�K����
�A��\]K����Ow����ߨE)���f���r*����`�^���}�YeP:Y��j���b?Az`$�����[���}GQC�ے1���SlP�]��dOC�S�|���D5a}����X��h�_~��^�F���p�L	J|��BSZ0�&�Q)�%��^�馞9�ݚ}"f��Jx��m|�Y{=����@I��5�A�8s��`�Fy.�es��R���Z�Ӂ7�p�e��6�����3�����F����2Oo�)ե^�̒R��O&!r�z��P�1u�eF$�c���al�� �SQ��q��T���&妘]c��*��aN��'�� ���p'[mpF�c��{���B��[+j<����g
ꕈR��v�\�S�'�p}H>���S�|�h
���6�}[�\���2�6�>�����(�l#gt�f>���9.�ڽȩKݮ�ݗa���ܾWDq�<x��u��~ss˾e�|��gw�˿ܟgr2<��U��T�j�&�;��e�~��r@U :�o��|�g�|�����}!��X���kA�]�/������%�/�oi:���(�CǞ�%��z.y2�>/Ky�]q�a$��-�������{Y�jg܈�Վ�0�9g���h�Ad��C�Be/IA/I��q�	�X"�C\�Q�5^1��<���v���b׸�л�T�oK�gi5�	?� ��OW�r3�=w#h\[��p3�K�,���,'N����C�6���Lii��_������l�#(jx~�|�3��5����vě��O
c��M&���f����ҽP��Æ~ni���z�d���FHܔ|�v.d
a^�;E�nU�Y��Qyy
�({u����Fua�]	�LhzQ}a��ֶ� &J�2Cc�9}^\�r�z뼮ص�}���{��kG�̐���P�d� �B!��.H��O^����uE-���.'!������5�!�{�bR��+�>s~،^xo�ꖟ�d�ty�y>A�{������lV-۴J�}l�^��隊hѥ�7�dܪ82K�4��m�q]�����~��mђU�������8�_���=��z��X�v��Jk;��;��p4�y�+�2��ɇ���3�c�-���f�'ƀ%�L|����ޱ�3�(�x��|Ǵ�`d�I��G)^�R96�U�Yһ^�$�t��CY��-�{Y2�j��� �~3��c�x�%�N�����^3������oL(Dz�n�������p�'��j]X�]k����O�I����맶�7 �3f���t7��+�?.���E�0:b��}�cu���H�S�׺�w���9��{�	���b��Q�of�+i�Tl����s��.B!'�.�6�k����Ɣ��&d\<���嚇��y��������F�0�nE�*3�7�O��@N��`82�*6��ۨb�:��S�P8���WF=}��-�L�p�!�'�%�qA�Yvk��n1���K����r��������99`��n@+ʆܘ)��Y��L~ߔ��B@�&�;��1�v+��ԇ�y�3��E�`;^7e�4p���/,}�r��P7R*����q���ͽ#�O7Z��xx��t���2b�9��|^y�zzA�rO8��<�^ƷR
�X5�
�~&�l��i���C���C�I<@��=?WXk��A����/f�)�q��V���D0�=���n��}�[Q�'�7 kQ{w2`0!��68l�(��W�n��m֧ئ�V������7^�ҥ�c����H�Ռ���	�V2�ا>(J5X{X�{9�Z�I�7�ҵ5��g;Ϋ��cx�E��[hl9sy���i��2oo[ޔ���]{��k�͍S�u�f�w�Ê˲�1c)�oM�j�C?���u�<x� �>w�|>}|�������x���18�%v�u�O��A��@N ���` ��Ϻo�jI�^U���k3At�t}J���S�|���y�=���P�������G*�cN����W��{e�΄<����N��)�f8���=y�J^\
<D�zxn�q���dщ�\��wn�_x���1'8,?�p+Y��;J�Z�p�ϥ�� �z�r��>���엧�-��G�z���tDy:�|����>0���=d���}�+���r��ߛ�5���^�˴�mn;��W���������
�y\��>s�Qp���*���,��7��È.��<���5b����L-��CEn"P�����!2�j��->	]�+��c��o"��� C��0���t�'�*���˩�[�x��7^�R��;�N��oλ�R�����P?��J�4�V��9�����&���6��;����y���=���>�2����ɹ�S$���,��>q�u�,y�"Ow�M1[d�i�<X!��l��\&�zg��r:<LW:o]R��1�d��2�/�m�a9p����)�L����7NU��n9�ݝS�<��|n	~�Sx��啕��_z����tk^��+�uӳ	�Yb��JZ���|�.ua�믦�aϊ�ڱ*BbO����U��n�� �דjެ[/]���+�SA�9��NW9��<ޏG�� 	��}Җf!�lז��6<;�M�?������M�fD��;�9�I��zNZ��9�7n�'髚.NY<<q��~���<�!x�� _5��=+B����[0[�����^e��K�e�Fe���$=��330l��C�9��U�n��-�o�J�����������Z�=���c60p�I�Ӹx{ku��ߟÏGC��N��y���e�a����`pc��6�xʈJ5]�C���l��3���V�ʶM,�ϛ�>�~�,�7"F���hi�lmC�;CDO]ͭĮ������!�^����%ؾM�f�rs헏K�k�tE0���M�!�x�s�RNi~��
?V%R��J�G��@��\�~���X�Ր����@w�
؎چ�z��ӄ��v�/lZ�%��\(�ȧ<#�8���Qb���/$z�����&�m�ni�����jF
��	�|�w�X��'b��� �����s��}<��,~�w����%��=�Z��V��'��sw���|��RdS�zËhs���ߙA�a�oti��n[�e޾�����k%��ˣ�%�X��5̪�f�CF����Uv����F��̒�����e����]�q�w:�ȰX����"����]��]��:�� ���uʑ!�;6����zg^(<g�9�μ��fg���gL�s�s�ZWў��D��DK��R|�p�>����w�s�P��~�(2j����W���8����O��v`"��m����vʖ^�����W�S��@��E���2}lY��s���P���M2���uA�ƒ۴��]�LZ0��mS<:��#�Rx/�t%zS	�y��)[ל�d����a)t�ܹ�$���������JX���Eê1���ڄ%"a�eO�nI��iRN^'m��h�|�F�Y�l�.ι�St����i���{����E>����$/�Ǽ�DZ�^H8~wUEM��:�w�NʌR�=&�̤Y��f��v���;"��YG���gݙ������ꕷ�,�a�f�����Tu�Q���^쐙K�\�������񭝅,��5
�y�f������탌��)?0%�A�\�`q�O�K����}�02�-�3�m\,���-��'d�ă/@@�p|�ƅ}Q���ʄX{}V��[�F�װ;����W��dDc�X`&b�aؔl���B���p��b���\�.'�������\#��m�6�v�9�V����u-u�*,<�L�~��g|��*��>UT���F��*ʂ����/YF�2:O�H$�l7��w횎�R濡��p[��er��M�z�
S�z����'n>������o��[��K�W�iۇ��g�e�/���|x�d,�<]�<���,�)f䐆���`�m�qx��cS)�C^L���M�ko���,���3y;N�s�W;2���D�o�y,oC�U���a���#�N[bc��,g*9社+�;��C�wpϞL�[ϋ�G����W��3����mt�H�-i���n���9�r:�}�uK;�{	X'1���$�'�B��)F'{�1�r�w�=����3m��0�;l�0DU�Ɯ��{���N�p�09בv����Sg�zR}kzO^���
e`$�Y�K�S���ZL�޻p�GM}\��Jb�'�����k�hn�:�stmqj�j�W]��Y�UD����>���G=nϢ����(G7�GO���/"����)��e2�q�05Jզ�[f��2s� �y[y�=
Rq{8�|7 hTg�$=�y:]�%����:���2B~m�����_�{R<�5��F�sy��n�c"��]�)�Yp)��ᄌ��Dc�KSS�֮�[3��o{ U�y���@�T1Ɏo��\�<�=!5E�E��5���� 0h[����RL��mQ;]N��x�
uB��غ�;�������a_��6`���)�ε�T����Z#giW�Q�{v�vK7޼�Д/Gi@�v{��R������cH�X/wJa]p&֎��O�E��2��@�[�qz*w�vA��j4����k�렷.������fᩞ{I�>���l챥�s�@=�ͺ).n��zz�h��4�,��^ȭmc���e�;�[um�����G�N��e~��0��̾/��gJ���k�U\�(���5��P�Zp��PI���+0�7��=غc���(|a�#�Fm��ޮi:��3R�R�Ll��ݪ�J9���S���ݝ�5ml�eN䲤Q���\�e�1��Aُ��k���\��.�/3:�[܊;����*x2�^���L|���8x�� �v�i.�%�ʕ�Յ���G/m4�'hb��Y�x�Y"-�tV;P�ty`���h2�P��*�����N���Ku6:|B���J=��>��{����ړ��78k+̺�\i�;��lg�hk�i��/f=��wWj�tjN����j�;w/A�UX����Tl���E�s[��e`���2�b�:7�&_FN\���t\ ^�p�u֕+��+{i�L����45�
��la��r�D�9@��r���b�#E��)r+HiV�j����X�z[!��gP%G�i!�M]��_��X*��gIB�T�_�캾��*��E޻�ܠZ03a�Z��<l�)a����jܑ��=�v
x�7���BuV��ȄT���ph�ꟊ�UG���l���,��m�VUB�w�P���f�,S7��q�s�0�����RQrm�vV5Z:��eM��T�N��S��X�����\7.��ډ�,JGhښ����՛GWn�+e,����Xb ������%�0b�����nd4�| ]��а���8蚇�{Fh�����["�f����}��� �����\N�[�d�ڥF��5�ٗ����[r��Ar���z�I�ø%��;����������"�k�C���t�����ݷ�L2��un������ �m��7y�_Ku���1	����+%�Sz_d�i3�c����ŵ�u��JQ�7^�1w�tҮSr�iKj��M�{2u���<�X����������u���%<r���g6U�1�Tkv�Цʭv�j��֥,;��.�z�\�V��ɀC���i���<Y�7 �/�<���^wt�r�K��}��t�f�aY50�{�5��̡;��KDSY/���M�4��:0�wE��׫����W��Ĵ@وR��x�	<Ds�.���_�#Ի�aTr���*��+���r��!Di%9p���P��K眝z�9����ǧ��������뮸뮺뮾�u�O<|}7���8�{�G*(���jk�!QQ�2�)A�vY3�*�d���<~=?����Ӯ���]u�]{u�u�_OOOO����hk�d�}��<�!�J
+�EȊ� ��}g՗���Pp.˲!��I$	pO ���É.IA��q"����+!$YQ|�(��Ô���&'aE4	�J��٠��IP.��7س�S����wX,3���dI!A��X9]�PG*�(y,���rH-Zv���"�{�9L����RE�a�9Us�#*Ԯr��]�48�rR�ZpJ��vSN���	el�zz�q��eەЄ�ie�@��D̈�����
)��S��PUS�©V��ʊ�9BQ�r�I$HH"GZ�$��"��\��v��˝�(X�����Xv�e�Ԫ7"�;��~Ȳ{�c/���c�"��q߮u����}z��r#�zg�Lx� x{��������*��)o����7'�LiG�o�¨�/-�P�����UW<,șи�3�Ԝ�]G3
ԇӭu@��~8y|hi�U�|y�P8I�~�U�+��U�3���4�5YӶ�������@c�0n��>��8P�B`c)��|�GW[��N���˦Nvv]N�==Omj���7:�U����'7�|<���Nu@�?]zԼ�T��G[f�f�mU��`Yx����|�X���+����k�Ĩ�6C3��:��	�4Ѭڞ*ig]��`��PZ&�\�\�s�|��V{�?``S��l��.��ĭ#�s �&�g�z��� 
fop��oVk�Rr�"��vQ"D��f1ܦ��� `���.Q���l:� ]\���3	;�1o<7/u���bM���𮯾N���r��/z��y\�!g��u�����g�}��Ԝ���1�����/�s��1Oq �x!�/�A]��؃��]�`��[v�^�ne�D�5�\�R�x���x?^Ԍ@.���z͜a \�C�lS>���L8������&ȧ˔�����qh�&[Cy ��wg;T��I��Τ%��[�-Ld�8�#�Y�����K$��t�G�̻�L"����]�E�3�7)���q��9yO�v�REP}�)������j�K5���ř���\��ѽ9�c�k'N�y����޿7��+��<x��R�D:���{�ל��������B�:�|d����I�WO��1�U�j�39�}(���00�>B�ˮ��F���YG4��O�hVgX
�Jj�)Մ���ɪT.�g1�ok�:yjwi��SC#lB ���u��q˸g�΂u��0,��0�W����7��I���2�$�0��8^|�1HFSО��S���w��]{�<��	�4�Ct���r9��&+�0�.�\� c����̆e}�U%c�'4﯆��{�w�b���t/�X��N[�=B��HNo}6"�ԟ��<kneUU��G>7yR�7���֜��!��B��?;H��xcO�C��^�ĴqŝQg[r��b$3����SmɗK e4�^��i����#X�ã�I>�D�|��W��W47�Cr
Ms
���Q��ObUτ���t6-���`��U}�Z���ks6�%���� ��뢎�=U×���o�91W��� �����3�=�7�;uLS[�:������
{�╁��՜�Q.�-�m���Y�q�����vs��_<����=e�f[�Wt���]5P�Pc���$n=��?٧�ו��(~#�,W[�	�@��)�%�4�m����LB�kjJ��<0_R\n��6�*��y
2:l�$ɘ����Q�Q��IqK�됳h�mͺ��&0 ?9��縸����D�Ai����]a�=yz��[�8�I�3�I� �[E�Y�B�HR$��c��>�A���oCGOxۡ�G0�P�Ox��/����*�!��X]���� ���:��nɄ~�g\�n����D�<e��l05���̜�^��l+L�pD\���f�i��	]ҘoL���q"�.}��y�fuB�����w�����m�G>窵Z�:�'�G���	�̨r�`���s�ƃ������h��r~O�8j��E�~�>�<�H�o�����o��W��0u�j��OIt�
c1�ޢ�y��`��z_����|����b]� ip%d{S��ÜWtK$���k�
�m�c�k�W��Xv{3;���WW�j%~pk�����33y�����l$]�ׯ:oBd���mk6&��p��������{ՙ�Se���3��6/�l>P���0-�����X$vz��y\l�gڴ��Y�6�]�����1�I),��v�{ز�|��y�>;|�8'MҸ�Q�C��M�U��l��&�òY &�����̤���F���s�� �Z� ���w�~�W�2æ���$ت��*��k�QE1w�	���3RK߳^��R�����W�>�b �l}@U4Xk�5ۍ��W��wb�y���2�R��Nܴ)KԴf0�����V]q:0��/��ޔ�wt��3�9�>���q��<q�
4 �#J1 �x{�Y���q"�[����K��=��O��%�쐙K�[� I�M���H(����>�n��}��m/�|B�w:n��}0%�vg�Ů�%z�8��Jz�s�U#v�����5[.]�3�H}I���x�>�~P4~_yTX{/�Xig�X�;���̵��"�)>=�fgo�>��\��>X,�pb ��ŧ����&<*�;��k�tO��f��bx�;�\�Hq���Ҝ��P�BK��O�=!Aw�}խ��͓�ێ�/=6�.��l�A�����܀RU��G�?z ��W@4V� �1�\��oI٣ْ��ɫ�ڼ��m���]|d�^G�`�����\�11�0oވ�,6y�Z~�	ތ��y���߽�y�g��hp��.Y�˼�|t�`I�/�z�71�Pj	t��ٶGXs�Uv��5�����ד�N� W�X�^a��=�[QM�� $�`;0�z�Y99��5����v����sb�X�y��)�;�ӵ9����.�"������z�CM��~�4��U���7;��+�y��[�z��J��³4\�ve�3��n�ޟV��9v�S����ᢴ�	��.�'�!����NX�zD�r��6`���
/k��&_nq�6��@�nN�Ƞ�{����<Tg�x @J��d�#f�����0e� f��
x���q�Ư���Kվ3��ޅ"�z d�-��Kt<X̄r_�R��[7>��^����	�$�F��F�]y�Y�oFЌjN���r����NoۼR5X`>�^X�R'�ʤ�?HM�����>��Ͼx�f=S���$�U���ۺHζB�����Ͼǟ4�VѨiܩ)�)�:�����\f�����+�[�k��������~h��=���1��y��z�@o4�)0�����ݓ��ZO�(Lg��e*ݻ.��ϊw9�l�P�
xw������y�n��KԀ���\�z�Wl���ʀ� V;���Y���rN.k�n�	�ZAzJ� AC��!k�|��<�%?���`:�y�E����=�cP:d�6��!�g��%�l�,;j1�{w%�
>��=1��b��JS��5%�_}[�f�ح��jvxiV�),J��1���y��=�`���*zd��
��b���e�ε�c�^�a�k�z|��cp�a��}=^�n��q����z�.-����WEa�K$V����:)F,�}g!��OO�g������{��Ҙ���'�4�-��Y=�q/N��������ʌ?Y��)\���c9!<�8�p�E�^��|D�34�+F����IN�0�⺳��J�};Mm�|?�^w����p	�?g���Bx�Ǌ�D �7�<�^�؎���Tk�<��;�O�ѐ����K.�d�
ߘ~}�!⋞{�]Z�')����T��>����r|��B;|� *��f�+�J_�e�����7���N�[�������kia֪r<�E:H|�_|����xo9R)�8ї�b����En�4o�2���2�uwOfz8�ka��)�V:)��X���G�j��{+O��{��.��P�z<��=~v�1L-u
N��\c1�[ռ4��;G�趫�c�ۧ��h��s3�y;�P�W�S��=�:�������~J}%�`$�1����<��w�h��n~�ϣ���D�=w�g��&���*`ry���������ct,��+�l���÷E����v��G���4�Tss��	�5��l��� #!I��r^y����2�Y{I��˝��)��;^l�ܯ+mC8�U�5��Ң�|��C��r1���ճ��@���[��ѻ�,��g&ʳ,M#/Z�\d<�su#*�y8�:����� �@���0�ΰ�%�mpj_){*4��a�z:+i;ԣ{f����+���wV��Q������qҍ��k���Ҷ͛!R��F���5�X�=5k�&�]uI�jJ�>�]�Y�Qܗo�9��N#�kkP�y5os���9X6j����0�~  y�+��� �x"PA(*���0rE����eN���;�z�����o��Av�utݪ�;nh������;rE}˪z�,�{YM%@���i�x܀��k���[Ӷ���#�9Z팬��B6��ĲT$H�R��`OB�!(��¸S/b�n�`ո:�`�d�6��={}aׂ p�Eۻ2t��v�+��P�T4��|ootzu��)��#�ߍ�wy�+�D�!��Tg�"��(��TG���`�|�ϼ����r���e�+���YC��=��>Un�u^A�'F뀼�[cPb�^�d�s�%M�r��6UB3V��z
.n��^#�iE���=ݞ�� j�l��o��魮�!L�!�_�ޘ���N\?�ha��e���F_Ob��Є`��o�8<(g��y���]�h�-39�
b��A8�B�����{����]n��N7n>������4�{<6�����F�U�o<�5��e�����Ο����(H/�ʥ��;�Nnwft)���"��>Qm�fU�W�{���/�ɭ<'Ժq�xq���#5��U�l=Gk��9�N3�P.q����>�$��8��y
}4�����A���͐8�{��a�6�/V�;๎��ȣi��+��e;Y�{���Y�i7��M� "݃)[ʰ����@
��4�A����/�P����\1�����g���/�	}g��ٓ�*�������"�zo_3}����|/�����ǀ3ǎ<��R%
�
@>{�߯7�{��=��6�mY����9J�`>a����x�"�$�=�"����M��W��ܿ���svs�]q9�Q�'��M�T���A�&��q}9�> $z./��Z�TZ�qdiC^����c8u�i�vf(w�B��$��r������9���L[AG�?6�r{!4���=�&��^R��By�#.��g,��wE�((�[�#xİ�c��Űll��Ӵk�eV٬��1C!��;;-{�[hnp*�Jo��	�R�����}���'�yyx���>�ի�jwt�W�+��E��ߟ������f��[	�>P�%=XW#ϥ���:i�������s�Z`���~� ���9��Gι�K�e�xJ�bK�^5��L���+���XV�I�긋d�C�m���3�!1gld���.��E�K8gg"�ͣg����k��
	��[y�>C�)C`�<u��7�覧���M�-����BiHnu���	�OG����D�#z7�Ҡ1^�52�'"a}g��|`s0��WTֲ������s��H&�4�*R�
�5�[��jn�h��^!��>�M�N�w�@>�Ҟg;�t�*rTk�][����-^�(:�U��No��);�t��KE��'8��7]Bdyٟ�W��L��q��<x��I�R!�y�սi.��X�Y�3P� @s}��鬿X���ҡ���8���vz���Z�׋ͼpcM���V�C�t���Rh��GP~���"� ���n'K�:.�y�/��<�Pd��t�k��g.0ksi,;b��eMT��!V3��*k�s���E1;~��[4�	���}��i�Ag����J��3�6�.b�ֿ���N.�Ÿ0�^S�&�[�VJ�T�G&ּ!���-�bv�u�YU��JĪ���j�y��xB;<��􌩄���p*�D�M��lj�'��2s	����Jt�H]
R{�5��0��Ш��	l��ېn�1v]#�i����eN��m���L��d�1�I���S����;ݼ0�xֽ%:Yf�ua�U���2�����q�l�4�T��X�e40�P.u�4�	�-/#sTpfq�7�KzWH߲soV�zx]��wy[�� P�2AŴx���_���5㔘Q���zn�);��d�X{6ms�f����"ji�]V��^8����<���6of��A��3���
�_�B�wqA�����?MeY��/�j��Z4v_�utT�ß37ob��n4�ٺ}-�,g�>½}}�\\��R�9,�D��b�ẛ;T�⦋�л�^��|KA�=�aM;+s:s��̽��E@^�x��}8�x�ǀ*Ѕ W�� ���';)i�R�L[�Ԛ���g怩 �P �Ӝ8W
_�~����䶹�[/�i�gM��9�hk��d�$ek�J;���Aa#�߫Z�~��[-��ziM���}�N�W6��d�xZd��./�'�4����m�l�G�=�&{�i� ����^��	�m�ݺp6��X��z� �� g�DD+}q����w���7s���y��U�1��q�;:�����#Wۧ2��Ω���c���yv��v�~Ύ�Bn���T�K��k�P�5�B��]���ۙ��?
�vf'Ky�u�W>1'�ߐ���&e�n՗v��¾{I�輈�wr�+��1^�s�k$H�y�\m�j�}hg�X �?����'�.#2��u6)����s[NOb���mz��_�C��������ʗ�
�|��,(��Mʑv�eN�Z����2��.�d���|���]Z����(P��m4��)흚���Q��R���T%K!�%�D@�!O�4m�֧��]�)�Q�t$�]��c��A���3��˖w���`�kB���sp�c9�\#b����y�:���o6��,7�m�"�[ݮW�9Zʂt,6۷�]�+`�7dZ�:���pWp::
�-�w�jөg�'V��{i�R�X!D��2�Ҧ,��bfM/>E� �WT���C��+����'��;���`pJ`#��ktrv���2���;���=�(m<�q��"t�Wq���mP:���y�ʈe�N��9Զ3���Kr����tr�P�����n�00�[�q�!�ďa�C��s�uMB�6��9�$*��m�s)��"������b�Ŵ�������͔:�d[��Ḿ����37A�|�_VS֣;Ϛ�s3��ךo~�'R��_v؈�������ze]�n�u�ve]�Q����wY���\F����'�Z���onWQBAއ�Ҽ���}��T�x8q�����{�ֺ[ת��m_55]e��lNv�Z�ܻw��;�cF�G��Yz��vn��>t����p�s#��0���`�e�������S��]Lp�;v�0<䖽}K5�1�]71YߟR�1^Yv������-�s��d��Y�[/��ۏ�#�ٳNZ=�c}�N�]ƮԙJn�{�o�.���{�z���֗U��7G>�}d��8��u�ZX�����۱�M��.��:�M��Vs�Nywrj��ڝ{�;�E�]��%3�v��-�,2ݵ��j�b��S8�͉�E$֍��lFY���Q�^eTp�hR�=y�ʪ�vd��[��[}滙��-�z�+�\\.�ϑ)Vv�4�]�Zڗ�6̽���HH�޾����7,��L�Hj����@+f��hv�^�Z�T/o1�E.�k���x�w�7+5jm�)�5�oc���sαA��%Z��<���W.�
C�u�tmv�K�w/����Y���71���[�O��q]'.�a��
H�;j�l�i;pdz2�QQ��N�Y���Ft^.�&sx�'ח��l-�A}u9��F���%j/l��Bt��]Fͮ��Ԯ����2u���,�5%�{���	�����vмYΥ���%�6�^N��4)wBaΆ�h�;b��Ւ�ff!I��\��	�Fm+A��G����k\�|��Tw'Df�}���ƒ\t��w���@��� ዂ%��TշY���v�'S):�]՗ӛ�*f3�r)j��A�2�� 7�2�S��J۬�G`#��e�ovӳ�&W�fu�����eR�ŅDqW���Bp�]�@�����,�;y��^*(�b�v�A�|�8�voB�r�s�P�,}��P��;Owb���a��h��~�ڳk�1�ծ7�8���O�'v���wt}�����h�N��|bЭ)a��4i�U�����PW�$h�D#�]&KMXkǏ���n�}:뮼u�]u׷]g]u��===>=>��x&{�>v��J�
�D
�i]���TrH�@S�MPUG02��<{~>��o��N�뮽:뮺�u�\uק���������}�s@(N�����T�j��vQW��*<����AIIЂ�Mi�Y�I¢�t�v��Ua�9�-6ʕ�� ���I$PE�´L�؜�����0��;H(�� ���C�NhB�9jDDgB��wC���r��fAfUP]���ʈ��;rr8�D@J��N!$�()�#�\֐]�����9<�\�TUr�����N_�!ȋ�/�5M�rq����ije�8��J"�z��"�I�����vQC�DTU���Й�ӴL.E��ED�@OE��}�{���q��B&�(aED�h"Crb��#)Bl�R&S&BH��}y�"���ޡU/�N}|S��
��=�.�D�#ͻ.��Ȼ��^�&��$�u֢噦�o�U�4�,{Xh�"�%�b&B�0؍@Ka�9F������d�[i6�d�!q��)	�0Ѣ�%EF����jB�n�_t�����S��ϼ]��Y�t��}��N<V�x�ǀ�B� ��p�V��^�ͽ��Qj��wv��s��'8j�;B�$lV计����A0P���x��_�Ya�C�|�08�Fk�uzA3):�7C�]'�b�]4�M���DY5���ޚ�`����h
oW��k~#�\x����<�r��|
9�M�@xbCW������;��؃�Ž �����]��PQ�r!6��M�,ȞW�q�V.g�Ύ2.w
�OK�Qi�XJ9�P}�~N(�{XZ=@���hX~Y.u|$����;�fs泆v:���_�3HYʅ�)�~#YM%@�X�4��l�$D�#X�J��mdk������ד��}�1,�L�c;;E�ҋ���T�.���5�M���m2z"����;�2���,:J��~�'9�<��FO�ejy����'_��lD�m4�(�6fP���َ�����{����t���#nW>�C�ψx��R{{T嘉��J��><�	G��4_5�2�r|��^�"T�=��%�;-�6�c\K�Pb���{X;-���S@�������#_��0���8v�.;&I�N�ݐ��[i�kCV채�>jW��íҶ�Y��.�e��;{6pu\r��o��`��Y�Ȟ�����|4��v'B�H �O{�*�csw&���w�;gea���oy,�0l3f�ۮ2W,䙜��)�=��@��'sB[��7��/�9ϊ���O8�I�h���T�ɞW���l�ς�=�m���L��Ԅ�w�CT��@QN���l8�Z�9[;����cy��ǣ^i�*f82��X�5��Pz͜/C��6�*�;��t��;�NYa��d�����w�q�R��v�J�	8Jl�2�&��R���Ћ�3��*v+-���Wo�V�ʭ���L�H{O�GJ���8s��I���s����}�ٚ����'6����Ξi��$t	�\:a`V@�;s��1����d]�ɵ�l��k�1<�}i�cXIV{��[D����p tgJ�rgi��p��S���Ϋ�0n��\�p�T����r�3�J<�s�wFkן#�^oM���|u��*���U��'pu�)�H��>�2�>܂�/����e��Z�ʑ�bXa0����B�jUr��n�0e,�eB�/��P��������������쐙K�PK�|w�wf.jW�ٷ��
Ծ��D>�=�_�@^;�L_���m���ZɄ�y������1M9Xbg���i�Q<����}��7_�h��k��.����pL#6臸� ��糧4�ũ����[Y�Yf�2��)=�/��U�^�D�g��z/3���wW�pF�6�ӺT�gp;��7�[�M�ƽ5V��������<q��#J� ��{���מs����}ζܮ��ݦ���AC��<�C�|����n﷨Zˉ����z�f�'��­��i3��5��H�żAXЁP?��z~�����d8mD;�-Ϥ�Z�9��P�x��+e^�c�^�i��mx��x�O�����m��0�^IG�^�N.��&e������LO= z����� ��/^׶s�!�be�of��rѫsg�4m�J�Y�h��8��5F�z��p�3,Њ�3��J�v�}kO�G-���K�m���Q͵���̽�`L�"�0��g�V%�J�:7����P�x�s�^~��H��@!��6�q.��W�߹�Y<Z��I1c�X?|����ȧ�=�sm�'Ƙ�]0�o��:j�k�+��r��wV3�A�0���$��a�X��魓N���l�ү�F��w}~R�⦃{��P��)_�W0��{���8<���x�5gq��|x�5�E�X��b���uu{�G5z�'@W��Ř���!�%:K�.�^��P!�1��Y���g������X�[�^�u
�"Y]�gN0⽩��8��"`�M2�8tT�vPr�O{�n��n�}Y�6�|n���L�$���}�J��_�UI�����CɞM�����I��	`s�6�ͥ+���Фm�yÑNo�{�hg�ۏx�ǌ�+$���`7���2�;G&��p����bp�&:Sp.9����t�{�W�ŗ݊��l<�4R��]�w�����
1��9�08�[�e#l�3n8�)��)�����!3r	��_9�7gwK���B��>�vW�q uFk$1f���a�6�@�|r�
�rx���z���B^%m.�6h��u�܋�L�О��|yx���dD�^���>�դG�N㬒M4��5�)a�ʕN���fsj�}@���Ü8E!���u���!���:��長yڄ1J�WS��q]�ekϒ�綿*��x�Y�S�x�������hפ�n;ۓNJӔl֖vgeL���<��.@���s�`s��|v=�++ަp�P��g]i�[����H�|��.�L�S	��7�Fؘf)�����T��X�I�;-zJ<.E�˵�4�@�J�tɣxޠ��\QV��L|>a��Q��)ӳ���f��2��2��ܮ�9��f�z��}�`vt��nWh�	\�|Ĝ�w���ER�3֬��>ﯾ�a�r���Z}/��rjp��/*d���7B��)v��F��+p��'��_.٬ N*f�8���N�(�wI��b��UU<[)�g7��Awu�����+�n,0o��@���Ы�t�.�p��|����^��7ޜ�X}�ғ�n'�<q�C0С,�=�y�g7:�����T�[��[C�]�^�Cv3��I���d3��N�/�^l�ʫ��6޳�G��Ԟ{�B���q��=C޼�ň,d���q<�7tͦ�7��v�-���M�x�R)�zE��A��H���
�|�DK����J��'��ay���ʴٝ�Fw3�~t{m�>}�%5�	�Z��Į����{Ǭxl�eG'��6��:��nqdˇBf���1L�>���:���y��%:�%<�3��|ԇ����L&C�w^\͗ͻ���gUsǖ�Q�R��F�-�u�Ǽ�-#lפn窻���q-��U5hu�t������m�_ms
�Ƴ5�����s���	�1�Cr0��T��C�F_U^��DU��J�|a�0[��b[��z;���mxw����@r!6И	��;m4��:�ݫk���v��vQw�W���=��!(��aC� '��d4x��ca簧eۆ]Q���9���x�$'e��g�3O�Y���5/�#YM�����sLC�p�-{*��ud�o����;7Vz������^p蹡1-� Cu��a ��װ�;���8����������7幇4�o(�;��I�,��w�z�;��%W�&�K��F_U���桙/.�h�g�[C���xeS��:v3Z�0\Qv�"�w��`3Wun���Z���c�ڬNr��f}}u��.���8}��Mzq�O8񈠖R� �3x0�Or�U5���&\0j���}�_�=�9Z���}C(jy�������u���dnA֮�3d��'1tyЬ��9�*�o GG�*���k|�q$�� 3dxm�/��nPw��Ȝ[}t4��>��h1���;�����h����"�0:��7�r���P�ݦ��2�����8�:���0y�h'����E��(��2�>2���d;��e?o~�3k�\׮�/I�r=U&Dh���'ǪG�y�B���F�i��ƕQ��G�·*VZ�����%�->Í�B}�Ѽ�
�P�6��K��߷'ɧ��9���m�.8�4��T��S���,:ב=�+��ьUϜ�%5��s0iA��<s�����=�Z.j�ǻ�2��#��ު���8�������8�����`��������>{)��Wr�:�.�b�(�@SL�R�Iͽ���`��֥0���k�.��u]����]?�;iMk�vQ���:��=�Q/�	(Ȥ����$O�Eé������5�B����w�Mv`��;칧7�b�n6s9���E�طi�ECWج6Yݭ����@eDm���>�����u|Qk[���,�Qئ��ݧ�GW6�[����S��$��lӅ�L�J�dohbG�.�ŵ*MWR����[�ϳ��8�*x�Ǆ����0`{��Wvi�Ux}�C��`�d�8�k�'�?g�7,�t�R�U�Wtg;c��l[wn���goU��ްC/'"9���m×�ޗi�YK��NV2����r���,.m�m�c�)���î��Ag�E�����LKn�:rQy��	���Q���>82fgF�-s���w	s�-,�8^c�a��&D몘�����k�e'��D�W)ɹ��;܉.3����UH�طq�`�6���]ٹ�?	}l�}"��إ���j�x�n�AvNu�&���:	��7���;�:�#Ϩ����~<Q���{3`�mt�5��49J�'��c��J#��={�0ym�V)����N�P&xL2��sج��x�׸p�I�ϱ"r�ɳ�d�s׻f0��+��@8"�ֽ���I�&�ء/y�7	Þ��0vX��\��zk����4"�g��r��I].۽z_*i�����ȟ�\t^�_�P�]u�KE |+���W�-���u�{����_�ή~l�OЫڳ��i����:뱸#˧�Hes1�Y���kʚ/:P8��b�sSR�SA��2D>�:�S�lΪBM��ZK������j��E�tP��ﶮ��r����:,��ᦋ���El<Ѭ�:�.�����k�h��xQK,��M#6��@�Y�GU�_"�m�qL��^�|�����#v�\6Ƕ���o]�[�qCFޮ4V_�9��uj��}���W��t�j5�@���|��O�"�zE���y,�{b���ڍ[C8`����M��n��V�o��b�R�U�)��rs��:�!�[�:�G�*{�O�s�{7�r��~�/m�mj��sw=��%:K�.���6q���BIY������[u۵��7�A�@.���S�ٸdI'ԭ4�p�$�m�=��e,ضڴ��I�\z�/-�N��H܁�ޑ��xL��C-�0��ʒ��tS.u]�W�=��x�1�$�ێ�q�r]5�^w�a��َC"�%���P��r�
�5�����ڝ���Ҭ���x����n��P�3�����i���6>9���_Umާa�~��(�[���N�ar�aK�U~WZ�>�B㤱B��13�\8�������L�E��|(��Ly@�@��R��=��,7�εx����޾�T�߬~�M
���J%��6���Ģ��tw�z�&<��^l�ځޙ�ˈ|`3�-(�n��.�☵`zhF�[��-ֻ%�\�d�k��_V�Rnv�;G;��H����n�C����J�9ҫ=�7��Վ�Я�ٙ��ǌ��Hii�
�a�T��U�O��350�t_*�<�����}�(�����:w�X1��H{,�=��̹����y҉^�?���Y�q�v������<<�V+�k��H`sqn�9�\O-ǽ�Gsz�_�
�T�_XO��C�o���~�`�f��ڮ`K�>��;v����o=tD�lY|o{g	;� &�S]{�cG=x����$��
�)F���QY���HB��C9�^���F��O�Y�44��.�;DY���x�?a#禬hy�#��U}N���s���Oj��$�6d�-�Z���\���!Euy��n�����זx��,d����f�ڝ�q��]	q5"� Ώ�{�P�C���c�:gZ��u��x*�0�{�N5�ff�`����O5C��M�V���������&~��)=��\c1���r�4ת�һxb���`趐��k�"t�>�Ѷ�Y��so��S�	O0L}���ѹ�	͜F�;�,	@�w^�����{w�>-��s�K�O@Y���H�7���ٔ����u�����]�n��|E-w�R���!�+��GL�E� �D4X]!mOOa\܅��<���[T��՜�%���[��%.�P����7�-�|���X�<lbA�Λ������ > ���z@2��5|�7 �9}c�x��u0�����J���*��O�A��K�;7+���c�\{�=u����?O����!*�a�Xm�W'�%sz���S� �*��GH/�m�s�mx��'�pt�l�k�F���7��s�( ��V��ƃ�&_��9b�n�eC��~�M'`=4y�^k49OW�4���>�����J}�&i�gu�S���5��J�/^ �|����;�Q�W��W�����'�0���Bb[L�e>�� 0�T�� �w?]�+�j8�&�� n�3m3(R���2� �ٵ�\;6[����T6�^5>�S��S[�en˹�+�Z�I�i�7"K�n�?���>Q�⾳��#�h�
�V�z����k�j��L�N�UN��=.x������LZ��ж%����F�UM��U�#�[pduG�S�y�g���=w��mBO^<�@��.�g_�F?�lEÚ�@���v�m�Mn�+$_s!�����X��H�J����z�ߝ��k�7�u��N�xh|n��P�T��gU*Y�|he��G�ק�?��S�G���e�2�Ùy.��=�Ț!�u��vm��[���+�=�8�/�#��X�>�C;�����
|΅۲+T�:v��ۜ����/�t��Yf��զ�W3�Ȳ�hǯd�ʔz��r�,;�Gx�Cx+�$��E�%���`��A��o,��K[�qۛ�[�4��E�� ���=�{h��Y+jN�1e���TD��Ღ�d��<��u�[=z3�M�+B�g+��9���^'9V��"!v���O9W�@^�xI|Y�5S��}B�	nƚ=6`r������Ю���c��7��{1���e�Nԏ����ɠ�&��v:�pq짹�M?F0�K%<֓0���+}v�����o�̔��TU�hH\Y&1iN̜�$2�]N�]�(�I����Πi�$��&jI�4�h�6V8i����M:�OS�[$!�&��Pʚ�g:�KVh���p:�����	��^_�n=W��;i�qyhT�Ơ����jYC�݆�늞g��ڷ��n(�V��ūXw�Kb��6�pSf�jՄ#�N.&�G�q3b+�_Ҩ��\��O�h+��p�m�� �&X�eގ�1�ۦ+q���ȏ+�*��]�ò����ʘ��α�� Ky@^K_*�\�m�8�V��ց�e>�1!� �ܹILr�B�6�uXۭ�;5�"��$�;lܚ�Hex ���N���Y���%��虘�וE��޻�p`D���:�����B_���،9�ו��<1D!�C�%�wA��43\L#��P�{�I���d�=� �i����:0�Y��Cvwue�����X�.`U�م��/����2���5k��N��|'�ۢ����m��=θ��J��YAڄ���`�(vA��IVz�,�O�hw����$8�i����c�F�R�ήF��8���:�t�9ǃ�!�#��Z�/x3�̃�rr��S��{��uAZ
�b��玲��Z�<r-{l�71`�R��m�m�Uf��"��o*u���4�R���Kso�2�$͛gm��ʱ:������瓎���][y.|ɕA.��LU�}��M�Z׏wfQ��ZV��n��w�i=���9{DA�o%��iJ�`ޒ(;�!KAY�9&�<�Z=ܬ�<%U[���1�w*�陷��4]�R�6�0��*ː����]��mt�%������:�-�r��\��9�7[�y�Qe�7#ӳ
�eh��k�(oU�	�����S.�G����M�P~YD��eríWP.x>�}x�[�T�u��k�&�0�B"cU�i�s�ZE�\!��ӏ���ۑ��Hk״�P`Av�n��d��;�T�3��O`$�
wa���wV�ek�8^';�ȧww\����C�
T$�^�xRD{���	P�C�EE:��G{�܂&QQ��;Zݾo���_�u�]zu�]u�뮸�OO�OO���M%�2pa5�2N���*}���
"�(��U��3��OǷ����]u�^�u�]}:�:�����������|�(��|�Qq�UȂ.T���.r+SQ';�)�p��y;�DS���#�	'�5�Vr�Q&PAvS�9\���Hr8�@Rt��|d]�0�^K�E\��]�EE�%U#�Bq""�G��
y��gTT�e�
Q+��]�(�������.���#X�?����$U�����C�v�G$�\��1R���<���<���84�����U�HP��"��Ҿ�ϞNj@zVI	*I,�����tsܪ#<���Es�l=�J�Z�EA@Efy���נ}|G�}+�+���|��n�=/�r��d���ʒ:,����ӱo�E\��oc���6��e�HH���;��}A?�<'�HM1z�Y���P�"<Z��c�>H2)�,8��a�u����s�����q�1;W���_��殧^�gŵ��y��̴�Z- J��9,�(��ǵA�@S�X�-� 8����uoQV�	�n/a.���R�T������><Ҵ�y��~B�G�T�ɝf�z1��z����(��@?w�3��?D�I@�E%I��G{��k�:����8[b!t��U{Y]�5���C��jw�Wl�q#����7 `JJKb^���#ϱ��L�?'��v�N_C4dz<�#XS6υ���+T�M�G3�����+C)�����b��0R��+^�/'Vf87��^�|��l#��i��ó�/�ĜT(�qy#�Fy:���i�&���ϳx���[m�����m}�eǺ�B�@��}#]d�>�4d���:6Y�L�l��^��.����}�e�y\��`e��w1�+�a\/�f����ʢ�ڬ�}�)����sk3m]��{�j���	�[���2�aU�0�����Y�tFr"�/g,o^�k�"_�t�;.Q�[D��B-#z�
�C���ʳ�!r��s7�T��}����Ml��\uo�Pz]^���Q�Iu���7ʬ��+z���Xt�e�uz�c��8]譗��q�����x�ZW�o?�����G��<��<�=��M�#�ׯ�d�=lA$�ĺk�5���{�#�����zi�<
��>4�L��o����pR5�>�;z�-ge��@x�n�`*�Hlx9}B�ݭ�.��>3�����w���'�}5i�T�'t�^T�Ș��+��{dK�!�z`yS�+j�w���|\�k�y������U���zb��.��Y�sq�(eo���ݞ�Ǖw!���3�"�|V���|�� �E���C�	�����˪�wzJ��׵���^Ͳ�n�SU$�c�1a}򁫵DPvǶ��~�����kv�E���|k�s�q�b]z�w}�(eE��x�fpP.E���N��u,e*�{+sNƳ��,�^O��س���!����&~��+IŁ�-��vu��Qp�Ol�a�5ְ�갩�_��څB/��k�)��>�n�nxN�29B��]���Sa$̔�q�w`��ђ����o@��i	�8�~� �;�D��T�w�;�L���E'�Wق������n��i�A�����ۅ���4��s8�n!���PӹRS���|/*�e�K�X ů��3�7��k,Y�1N����ks9��׷�:�5)������*��ν`3I�:��y�=��TVz�T���{ܨ��Kǝ9�|Ғ���{�k�#7�S殂C�\|\\\@~<�幻�����m��f�����v��F���#Î��ew]�؀������X��}�)���h�/8r��{h���r�.���皈��c�n�kx�}��&ysW�y�,�\�Q�ȩ�ø�nC������b3̙ˢ�Y^���h���������	drq[ܫ�R�%�*��pa�K�c�������f����v�/8��ژ	��	�0y��+O������V{�N��Q=V��%f�?{�����#������C��RXsN�T1���qL�m��/�A��`qqR3<l���3��;p�^^"q�;͹�f��n�pڮaD����~ԧ�O>8v�����k���n�`Y_)�Q'χ�#��S�dT�,�a7����%Րۙz��k:�� *��x��G��&v��	_1'��8{t�;�͖���6�ѭ�6�mW��0�nq��z��A�]^i�6��1p�����h`�a��������)Y�����
	�ױ'�$�ȶհ)��>�T��ھ�<�"���j�ٝ���A��	͝y���y�5ή��E�g �UP��%]!���<�m��/�uṟEx_�^iz�yY��G������
K�C���}q�9�+�:ˎ,�G���]�Vs�.Z�LC&.�Z�����*f�']�=1ʾ���WB������<�8��z���Ր;?���4tkL8����\{�Gy��Q�07<������=:��ꜹqG��t.9�٘i]�4��*{gn����Z� wHK���B2�Z��	���S�#���`�:rk�dT��5��c(��q����l��On�[W:�ʘ�2OC�B�����m1���e�[�l�^>�1�e�h�2IJ`\ŗ�5�"�׶}$t����D>����Uwt���WF��pz�91��.�N��1+��X�2�����N��?z-�	�5�*��n)�a��39ݸ�)�HL�<dO�\�;}�Nd����C�$�Z���ݯ.�,�ek����*s�W=������QX��zEs���}��^���R��\��[*�5�Snmޖ��f��.�n�,:�(�y�����lT&D��l��Z�9/T�):�-L9����F�Zr�Su#u���`�+�0<y@����U��:/�eP���1�	tI[]�,Qs�3�a\�?���d������	��/���˟X���^��9����������T���Nr� "y�9�@#�'��慪�N��v�⍋���#+�Ǽ�35�0�b�Çs�e�$}���^9ۯ��o��VmjIm�ծ��J���kDQو�b��5�cD����"ҋ�;٭k�{��*@�7���? $s�[ѹ�|�|�[�	e&+��=-$�(���)����89a�p�^h�>ܺΚ�5Ĝ+5Ժe�0	�U�G1{�7ŏA��#�\ģ[}p��QO.r�m���A
e���2/�^��d������v9�SͣazL:fc��k��+���smg<2�<��cKJ
y�/��Lzȧ���<����`�\��&�3d�q���3��'kZ6�e�H
_:~��[/�C���6
I�Y��uς2=3��*>oi�)���h���T6N���(+�oy�ފ/I)��f*�V�ʀ�C�������Ϻ��9�4Pu�{F��YF��d��	<2N��nR���ߔv��s�:zkw�
'�quh�nفK�<������l�'îN�Q̓�<'G�H�TJ�g��N�:��ǻg ޺/�;��N�|�a�;�!����A�S���aĝ���<��,ܬ1�H��'�sZQ��ڨ.觛S}ի�t:W�E�0S�A����>��kT�M�e�C�-9X�Af V�n��T�X[E�n[U��Q��nS<B�����j��L�a�αpfi8�bo�V�=C�V�ˑ���������� �	�|(�h�(�Z���1c�k�����`>n��d�X��}����yJ����9}�Y;:Z�K2pw�w|���^��|�����{�xy�:�J����/��+�D�>��G���Q��</Y���*�%s��f�o]�=�3����(��*�x3��y���('�q���YD}�2�_j�|w� ��h3��l�L��M���X��lQq��d�Xd��\�1��;H>�
c�f������,���m�5�=;�v�(�9Ad������y<?c�{g/���VZ�A��a�h`�)�>�V�c|�k/���YC�xfO��/F���89��L3����Y�#�3��L� >���9�)-�����w/>eP�7���cO���|���OoR<W�O?I��?~�mD�5�|��(��=&�k�k������v0�?���E�*/|���^޾]�^�/۳�筂�g2�}W�l�7��
9�� �+Vj�O�(tk}���5n��V��:+>��Nfz{��D���8�+q�&875�Pj�]!�b����j���0Ņ��5u�vG���m�Oe*��z)�1���]5��	� �VǞ ���'�1P�C���
��\����
��ed:�FJ*�V��H՗w�]�,>��yD٧tg�]X��=���~2�5�]L"oK}��iYٜ���i}��AB�Y�ɶ�k�a�Z�gN7%Kt��%�|�u����1U����\����5O�\�@s�����	 �H۽
	�+��3v��q=�ML���N�����D=�Ƌ��An�kUz-��u "#Ϩ~?����-t���v����}�O)U�)�ux�CQ��|z���ȷ�~n���d���g˙�����bb=�([����M�}��v{���:�b�
�JN.�j�., �^f��]���R�h���m	�8�����X���"@&U&X�2S�l���+n/2���������1z/�]�D��Ϧq��[Q�S��?A���S7O�B6z�Su߳����ܒ�<����y`�<~g�^�m^�	N�M(8����E����H��c�J3w;�}Z��[4^Z�e�N��w ��x'>M �u��FP!|s�ic�x>�=�'`�j(��OI�&B�IN/�O0�,������{mi��1�謾�8���nn��
�._�8�a 8P[!�{���J�����+^�Q���\����08R��3��ܿfh�}�i�C��gH4��aٕ�	�q*�:�U���&.�5�_M�;��n�6��C�V@Ɲz�FC3��<	���p:��{�;�g��s���C�z赀�����f
r����/�EI�̢2�e���٩V�ƻR��p��ꘌ�ہ��e��Z�x��/�h$�Lvcܼ���Ѿ��s��&��q�+AV�l���ꊺ�#N*�fr�4l�Y�n�����v�����K�|~����0�fӉf�I���p�6K�q�
W��Ҽ�֒c�<�P5>VC��.���:�?N�vY�ӹ�q3/��O���X�1�h��#�g�;3S�����2�_8jކƆ��e�ZNھ�kB�Z-�G��,�Q�F�v�ɚ�Gs�g��n�����זqQ��F�C�,�ۛ�?�$Ӊ���{��E��������Got�8zl��k*��q��N�l�M��6^��d�<
-�i��=�Y�"Wq��P��)9��)5�k�ڽ�[τ��Z�v�Ui��VQ���9�6����������Vxe�˺�0��=կ�I\tӆ�NW�J`����w9�[~�gO"���0���*`$�,��u�÷���YX_)N%z�#y�2Z���>ytS*��I���<��¥=�\<�n�2�D̆g�Opu�����!�d@vOCω��LL.t5�-��;���mxw�h�=@��ג\���ѽ�H���G6��G��-O��Y��t~���(��aC�!8�y���H+"C�R��7��2�~��Zi�啲N���{a�j��T�l�l{3��u��Q��s��z��Eܬ�r�k����"�K�*xn�����Yז��;��y+8_U����ie�%-�K����N�t�C8��ȸ'��Ns[���y������@a���sU��a����lǥ|V��W&�F��(��].��������	���*/j�p�3�YON�\=#X/�yísBb[zdK)��,(�(��q����)�(�on䕼�N���UH��u� ��ǝٱ�(vl�����Ku���2������CO>�S�נzO�:�vc����&<�P�����.*b�2Ǯۣ՘q49A@f0�'���`��$�/�ۤ$'+��PHz��g�������������A��L���߉i��z��΍Ǿ]�C��S���E�4���r�1=�U��֐n�,�&��t�,(�v�)ᦞ{FH�4\Q��<�h�C�tq�,Ԟ��Yo���u;�J��E<643�}hn�{�O��r�OMT(Y��H�QVTFp�噷`��E���;A�ٳ��c�?A�RV�`��v� ����g���d.����ѱ�ܽ�(2j������%v�Ui�P�+��a2*�cڷ~����}#@��T�;t?Gn��9���ij�{ƲX.��|3{b�
#1����=���ilOy��������$�8��:��ꨯ�el���z��%��9��;E#��K�.ݼرlWt2�I[�af8b*����w]a;�#@�>�?��8 Cz�3��j�v`Ç|!u&�0�q���9	t�+��ŧ8��^���y�=@��j��P[�.�Vқ=�m���	�tpu�}��=�D��+JE���s[[׀f�&FX��G��Їq#��Cx?��#%Y���wa 
��Z~ނq��ʸI&Q�2ۃ4�*I��r�����4�bC��g{/�ˠ�<��$(�?M�0Cl���+T�"ܲ���Uc�; ��V�C$�c;���� ̽}�!}�Ѻ����<>xc^�(���g2ԉ2ϴ�e���Y�R][��tϕ���r/������B��Y%e�@C,�����Ǫg|�����&�ޑQ�k��l-��;E��J������UA��i:�>D��A�3ZG�g�:��MO�UY��U_���Ժe{V��4�>��=��7a����Bp�����{�_{b�8��{�w��w�=!-l�D��O^�_&�ʆ�;6��3L+�@���W1�9��q;\/wϕ,�g/��d�"^��������ؘ	�����LO=�nn`��u����������?Ww�7k����d)-ݦScY���:Lҝ�V�.��Sz�q)���ŘC���0a|z�!u+�a���s��u���[5j����6��U-W;��77�tB��]��/�����"�z^�]S�x7�s�r��=pM��*�W[�m�롩,"a	��=��r���YS����u]��2��d�$я"��ԈQ�H��s�ܛ��u�."R��n�ucͰnL�'�B.b�%-n\�VNU���6)�v�Y�i��A�� �޻���hhS�7v����i���͹´�7��7U���Rf�MR�lQYVq�ҹ�"�i^iub�R�=x��U�U̲�Pi��ξ�����V� ���d�=��샐ziգ��r��(�V�8KὫ����O�����Vm�@�O0�o�s'c�	��C�&ӈ��2�$�o�H�ի
�#��M<��t�&�4�.����;D֞ܮ��Ύ��� ��mV���k�Avs��̄���}�Q�zI^����,�coC���z�<\��KT������9P{)Y3��mͧ9!G��x�R�='m��%o�뫮}����i��X[�k.�R���q���d>�G{�V몮����K �����]�Y���u�A�U���y�/�k�V2^S����k���̼K�+=��ڣ5���l�(�z�K-S+!�n���e��X썦���A~Օ8���pIU!71����A�(�n��JuBz�S��V��!�LRV�^�p'b7	�x���������8�����և����O\���vS��+FʚWg#�$"�iq�]-��z�\4�I�����o`���' ���I���-g��p�v-wQ�У�A)l�/�t��Vg}�2u�_b�k�J��?�-K´s�7w��o�7�y��f�+wܶ�����۷�B���GY���H��es���<�X�.x��t[~Ďs3f���pYM���Յ,�˰���rP����jxs���x&����6gg��=��m{�ky�]uGk�vՎ!�61��T�#X��E��|��~�ە�n�F(��b�ŀ� ���zgt�`���J��{Ei뵛]cf�Z���k]459���>X+r��9�Wp��	�W1.s\\��H�����+���-�q��y��ag>|e�u(��.�g(]_]���yoku�Z\#�o��E }{���_c�t��Y��i�w�.��  �xKL󵄦~���_Z��r}|��<�3�e�7%v�;��F�"VlӮE�+Ӥv^K;қ��M�}����kv�;�ʝ��r�V�.�!���$�N�tZw����]���]���7�N��[�݊a3nQ�=���=8]'���"�3 r<G*�!�[==c�P�J�IIc�<u��{}�x뮺믧]uק]u׎�==?g����X|�>!2�eP�2�;�A�\�f��|v��S��9�nַoO�������]u�]}:뮽:뮼u����������Ù���aa�,np��;'!;���P��y2�f��W.�����H|j��Gdr���(�8��.�8Qj���r�|q �)�TAt#���(̯�Ur�����Np�uM]��/qa�J��Y-�b�7���OB�8���:d�"�Wo$�QAq�N��"")R"�/!Ng��)�7���
f�*��xqLwq#�\�/�:�p�B����0��RW �^�p������z�l]�xʼ�T�p�Q��w���ܮS~6O�!�9����E�ϓB�I �a�����8�x�����i�����N7	q.�*8�I��"ICp��Y!�#E�f� Y��(�����)�ue�/�.�Vk��x����tP=�/s��r�8��w9r�p9��qk�qQz�1!
i�F��H]q�l���AQ�2D� M��Hc�^����:;�빙�^��D�!� �p&�(�q��M�P��xd$$�'�I�>���C����>$�x��.g�!Y��UC����ӻ��n�|]�i�L�2�eՠ�L��Ii��ȏ�W����U��>�Ƭx �:���H��~^����m�Z����{�Ws�q��ߌ�/s����Z{C %ty�>�|V���`K|��F��-���~Y'ej7�U�:���>K�z�R�6�Dg9�g�Ź�P`ü�ړ��0|�������(����R�.����#9�n�6ks�«#wni����*��A�{�+�hU^;�H�h�*�q�>OG��\C�U������u�AB�)\��b���n��V��/��̲�<zv�Ɍ�[��Kn��̑|�lpP+H��`n�]=7M��'��Q�u���]�65wq�S2��Fc���#�c�Я�*2�̸M�i?j�/!��T�����ڒ�}�8�&Cp��K0�]�
��rn�;���m^Y����#N9�q��]%I�εC8�g	G�I�����j�6�Jxm&p���Ͷ�F)�*���{�f�nu�rﲻ@L[hŮ!������lH��۵�y��Tk2�Y��� �
��HJF1-H:�{j�'.i�kn��PC���W	N��b��G�x��>Ӿ����h�A���I�'ՙ�۔���*������������ ��R�ň�v�9��uB�eW�r@F�N��<e���8흷��7����`ER`�����_B�5��8��7��aQ�7Hm1w��K ��y�扼,*���"Ǉ��O&a^�N05^�+q"G9��mL����.��3Nb�̓[}�uq�v{z*�����XF�Y��/5�=�;j����g�ɳ������@�w��|6Пto�t<*>���ﴶ���^b̊��	]�Fgt��sgo�@ח2,���NهR{s��Dc�r콾�Y�>���tݞy�]%U���M7�8����M`�j͵��ن��9�����ʯ)aSC+��:�{q��Z׻�y��ޣ��t+�-��_�U[�&YЧ�� 9��*ѸB�;��"C�������}�7a�>z~��R*��u���?t ��m�sh��Oq�?	\�%��!��1	�:�ӷ.�|����w����k��F��75>2���͡Dꯍ3���	��:E�rY%��m��i�]K����y��s2�S#0�*�7�t���n/v��1����:�/��qqqs��<�˟x�(��{/�g�;��?'I?�cn�Y\��Aķ3Вqɺ!̊����`��gut�0�#����R��%��;����2)����G�	36t�M�^VR�Η��jF��`��R�le,��r�76��C�����Tv�7{3���u2�؟KU��(�"��Uf�h��t�N���W*��X�ف��nNN实�r萭���n[�`��g!��Ǣ��Q��Ln3��L0��i��}��|K�i3�T��k�z��i�7��<:����xޕ�7|��q�zb���Z�d-"Z��͕f�7��χ	Q�ݧg���i�8��ޛ��XRTe��0_�7߼�������g���`Rk�=�\ޮ�پ�0;E�>;;ż�~�as�;k�b"�y�Z�T��t_w�|y�=�X��ݸ�{��L��"oSc%�6nr*iE�?r˭�ǵzh>��D��V��K6*�p��1����ҝ���(ky�.�^0��͉����m����ۋ2���ẋ�oM����ܶ2$���_b蹯�|�Y������?�����gĮչ�E����º<��\�OUߞ��g��
�Y�9�sz�`�=���N�߭��������[,�pT�K���Xr����� #f5U^�ᛌ����CN��<{��i`�edz 2TWD�A�&U�I�hM��"��n쓀%�X�:}J�=C�⡧2@���UA����u5>K5n����������}���c�Q��UB����Um���ܑ������Z�r�Ѵ�Cr]A�wWr��R\�e��6c*�s�3*k�v�ݻ�׈��<^^v'ãr:sV���L��� ��瞈�7uo/�{x��g�KP���g�Ѱ�k��y�-v�-���6�S$���O�ڟ5\���\���v=�_��Kk �����]6��uV6F�֓o����d�&�՚b@�IMy"d#���tl0F�Y��u��_���<g6��1������g<.�[P�K�_{���7�B〥�t���7���5���Ӂk�}1��v���o>��#�)݅������ř��	��Vg�eȳ7���;j��Ew�1�7{Qq�d����e��;�fS�||C������2Sht����l�z��ܽ��W�dv����)��N� v�䉇z�U�D0�do��ԃ��ǒ�ޓԣ��e��l8F�t��Rv"��������H��\ѓ��t���y� ��4����Y�ܓ�2v�1�����H�뷪;���m-��=]öGq��^���fx٩ު�a�σ��Q�%X1��~V���{��Ʒx�k$%�u�;L�!���/Y�Px���[�ar�g��ֲ�m�̏n�K�����|�B���@5�v�L�y
Y�e�]�᭲q��Dא�v�xt�T�������ж@c����Uqv�~�Dd��#7�vS����P��\�R\4�7N���)��Zw����t�y�� wh�(@@���Ժ��٣��q�ƹ�V�J�?6�f�J���5S�&��T+�� )�a��|�Q�pw\3��˾aQ��.��% ���%����i�.U��3��z����6�t�+�����wr�?-�@�[��+�`�����w�����S:8�,���ت�0>����l4�R�gg5L͜C��fv��enWw(we�H|�x�����Ďq�V�z�fk��͚l����wن�1�,��
��}�E�\9��q�f.�b��o��or�W��4e��df �eHϣ��@���;�[Gv�T:���uq�z�R[ϻ�ɟ0�^���y`�Iy�<%vU_D��⥷ޒ�;M�Tq�t�D�;yԨm��P%=mz'8ᓰ�9�l\y߻?� ��P:�����U���ȇ�Ρ�b;k��,�И=���8`g�hI�"�	LOg����W�����RsP��h�5p��5��ة��n�HY�x��b`��� n$J�w�q��zK�q;�E�5x��>��P��'G3��x�5���F�Ҫ�z���8eX=g-#���s�w��6�3a}�T�V�y�a���wMo��I|`�����pIO��Go4"��2&�!������������0jAbZN�*u���W�m&��=)�[�k��#!�1���UzU�/p�����v�9��!�vy�*RC�Lv�۸��]�;(d�'4�
.�h�r�͒�v�u����=i^��縀�x�����x����6��|�$i�t[��]�?MX�����Up��i�����[ۋ�'�>����Ub�C8��At�b���/f:7W�t���2-LvS�QɜD��wn���VZ�=sO���T��t0di]��"y��-1��.�b��ݬ�+�ڰ�j8��r*[��"���Y�?t|+N>(�˺�4`�'�8��Y�6A"�ݝ=�ݩW�%M�V�)�v�wo<�ڴ�����s�D>�����;�;8O�
^��
�7BT�zGwr�9�4�n��:<�����˞�{y�9��¨�Ւ ��ck<bF��q�=�w��3�ǻ�����EN+�[���)��@�����)������Z��*5���j܍ʾ�8�Α��E�B�<�)W�v1�w�Ggq����B���|�}}���1�w���b�4�0�i�@�N�)s��Ո���-#}�t���#V�Rj�)q�����ụ�+ߝ�j;����ȯ��W%
�V�V�<��#��ƘBDD=Xvf�W���˦��{,�ɡ�;�d��u�GQ����0�Zs/Z�trw,4�y&�d���=��G��^�?�0����3(_����h�/�^ R]�4�K��e)����	q���'��{�s��Tj���v�n��}]Ry�{0k�e�h�?05&�󜆭�����3���
�q~�G�G�^W��k�N䨺��:+<h�<H8�����׽�3Y��6�<D������Qx�������@�n�I���-,}�n6�V�ol��������=c�!u�<�Ed�Z��z�0��rwKUFM����GhN�a�������	�;�y�0�\��z�.�<��Lʳ�bm��6o��2
��]��������fڳ�u��8�w5�E�۝/uf��=U=-ڝV��98G�]qAH�=��9�.i�� ��v�z���
/��{N�Z�(�0�pg���J��T!tϻl���*M����NgM�Ȃ�dp`����V ���$���ܯ֬$�z5�|R�y��N���\��k젴!���(���rֺXSخڼ�@�vN��r�	:3�v����Y7�Av۬ȕo$�\bl��wS{������Qb���H��|Q҇MF�sy���r�̴\Ü���Vd;�� �g?%���z�$6�x�:��n~�m��d(v��)�-^�I�UQ��U[���n;[��ǭ���-�"�T���	�RK�����i˼�ǝ�;���q%��ُ���C��21�ѱ�)�2��,�"��뜪�p��:�����U�	���X_��X�[��>>��W�����������]��q�}� E*�)��q�����sa�8���qTX�md��9x�1�|n��@gܾ��B�Ͻ$�^W��]J:�$m6zd�E�X�T��޽���p�`���Wg�TF��hմv{���q��ac���s1��ڙ������#����d
��KKO�x�>;7S�=[��
��¼�/$m���ps��5%X0�w-��܃s�j�/7,��Oqb�f�8/�v���:0_3�>�Q���3M3-"n2j�vt�)���'�ܸ@ţ�m�0�O�4X�B�2m��M�3�v`>E�|퟈�@=�^5�
����+N纖I�uk�l@0E�q���
|&>�{���{�9�ͨ1;��ΐ�<<$�4��2�(6���|��=�r�gZ�8-7͝����<j�;Z�72��{�Gd��������ܜO�~�{������y�����0f�ָ��D�^}��Uv���)CDVJ�V�A���tc^�-n�4�绕��ݑu�ʯ���W)Iuϟ���z��cSt�6f�"�MKp�?�+�#���;�q�K���z:H;�4��T񪙻��~��%𜑹h�9��O4�#�G\�QDe(� �3y��Ͻ<U����C���������;�{���-nS�9�$[��ay�ZA�3�Z\���R��'��{��$��eO��6�Ϛ��Fc���-y/�s63&=e�$�W�y�J~J��ܜ�G��_�(�@�G��u�.8���5�����#��#I͛]G8�뤩"dv��*�+��`ugp��;��}���˴�D���0�Q(�Xk�U��=f/�$�ͬu�ِ"!�b��_�9�S}*\立>�<�"�7~�vu���%��CX�)[7)Z�m�VTD&���K�SIl�M�M]��E�Z�\X��ӷ�1n���+9�̹�>��ԉPu4��i*�M��Ȳ��6N5r�:/n�o�Z)�!�ݎ�`��F�W8��;�q�1<�m�feX�G�[קdљ6�{;}��v[��-?-��$�j�v��3���C�I���]���E:�����.p��uk���[���f�,+��X�Ak�2k��X�y�.�nM�r�M���ym�c��������t��T�o*��`��7��zl�ɣ�3V�C���άHVm��aM�:M�g$��s�vu�9�z�K��ypg2*���\J�E7j�����Kɕ&�{��j�N�뺦�(u���KN(�Ż�d�����O5J��^��P���B�M%˽0�l�<�������G4e�
�v.[��D�Fm��>mh����ѥ۳��د>G��;�M��:0@"�M̤����3;x'���U��$��:�j.g'3��X�7a��ۀJ±��5���{
9�v�:c���Pސ_ۨrw,��33Kݨ�=Ji��.��#F��G�I%�®Ί�O:���8j*�v�<;�����BX���7�pƺ�ռ6��wVΈ�Z�"ۦ�*(�z7��eYyvy����,Ve��(�� �y�rjf�;���w]�^���Ch��
�&
:��V�| �Y��wm/q�p���C����J�C�"��e3��<��ђ'���]+�HP��+�wx/n�!Sp.���)��íNQg]c\�k�7��o����#-7wIm;��7�YU����&�\��[w.�}�}�8���k��-�@r�s���E��6Y㵘�l�E��se'W3pI�Z��|1�ܭ����b�{b�;jghY��pmk�V9�>��ų��9�dɻ{���a,2r+vz�R�NӽqV�r��]( ���ܵ��5+0�����V��Ki&0knd�RS�3_br�"��x��E,n����a2���1tT�na��b�Ŝ{UAU���XӴ\��/�!���m�>�ΥJ��L��6ѹ}W}Ka�p���9�LB6�t����q\ͧ]B�	S9�z�N3w�b�s�D\s�S[]J[�Ҹ�2�����2���˺��m��U�X�e��"��!�K�;7T�t��f�ڰ��ޤ $e�ϒ� �ٺ\u��o�T���+��]�v�����S�`��j�-��n�Mn�I*����U��ɜ�\��7��Y� :̩�ӹ�ݹQ5E�g7݃���)�.��ﺥ����N�w��c��}�ݛ�N�ږ�H�c/�m��>4 }��\��L=ݎU�����"-�03�3Ǐ��㯷��u�]u׷]u㮺��^���>>3�?>��Ƨ~�H|xUC���?D������}I��9*ʪ	8�������||q�]u�]{u�^:뮺�������Ͽe�O�,=�r�d
(��s߰�����U�*��\�y���q*BO;�P\��ݼ��C��z�e<���mWwt�un�����>m�#��N�o�9�$�&u������=��)ե�tB�P���D�Fl"L���Tn�\ȯ�����{��Mʕ�X�4H���)=�pꤚiU�NZ�B���sX�,�I�U���MԸ�.�IeUy��*y"��^᮷=D�A�� �3�|�������:)I��ou��5&#��I��Y�h�=���)�n�;�����=�k���[�S��^�<�{�>q����o[��廒
�_��kdu1�o�h,㆘q��Q$�뵋5N8K.��U�^��͕�g+�0�8�ȟ9�6�iG���;�C�Ea������E��}��2��_q��[\�נ�P#kj�e��ϟٷ�{�(��'��X1����{�=Ҷ�yu\2hr(��Տ��ޝ��Fvi�#b,"��\MI��v��oqQ��o�j�z9�,f�m��G1��ͺ��E>;MP�r�O�2��}}T�WW���X+�i��8����;m7��\�za��P]N`�
Ґ.%��rb2+�4g.�F=b�J[B��fn���Λ�4�h�8M�ɰ%��� �)Z���%vn\���x�̳�3�ϓ���wrꄕS���2� S<i5�,�T֫��ܫ���pÜ��JV���G��{���Eߨ=/��A�śu�P4�C3:�홫a,|�|�����
�s��Z;��)-�x��3�n��V�[%!��oJڹ����@���٩Bd����f���-)�9Mh�Xhe7�Z�d<�ph�ic�������H���(ʽ�I·�Mp�����^C��������v��ߔC�/s]��7d��Uܭ�zT�;o����c:b0�N�^��U��n8'b;'�V͘R(��}�L�Ox��D0�j,�{m�,����a���~����>X�f�~N��+�MT���[s5�񓛔tф4���ݐ:ў�}�r��C�zb0���K,� cL���;����4T���oz�ż֔*�82f�e-�4�~��z��a�y�$�� �q�8��4v>���D���<d�m����9���m)��7�Co�#�~�e�S�����@��4��	�l��ɤ�5��M�"$�:�k47v�j�$���贯|ق.�Ϸ{��tN�`jƄ��Ӝwr۽6)#b��Fy��;�)*�U�P��/ԮsN�����˺�ٽ��f�HKG�+�b�ϲY�����>�����{����>+޾�|���isczb�W���ک�]Q,Yf�kg��J�;-Y�����Δ8��n����䳶��IN�p�r�^ϻ�E5nͽ:��������Y�{�>T�ߴ�Ky��/��q�9nnK�d��j�C�{<|��������m>k��2�����A�tf���Y��i��9ʕ���֨��7�����l8su/á:z���SQ~�<���`�Wʒ�i͵7L��-C���)�Ym׀�+�想y�=���ԕƮ�����

��{�ڮ9�bi��O(a��(�IZ{3z��z8��E33V�*JuPK�T.��~^�7T�\�g����smS����Lj���uf���i��c�ܩK:I
9��rۨ���k�����G���|S�@�I�U9�@�5�i%L�����3�k��`���l��(�_h���+��D�)�|�k;�t6>�2����E�1oJJ�V�c��aa,`5��`���{n�o%��h�5���2P��:�π�;m%4&B8�;>[\yf�6�ʘ��&ٝZ��o7:K��NH��He;;�5D�{�zs˪��L�!��k^-^Y��"��`�8������t�؏om��7��F�thH|nj��o���R���4�u����{Df�}�8����SŘls��C�gGt��p��r�'����5�y��Z�c�� ]� ��R��h۫��:ڻ��@�\&��1�8\�����t���Lo���;�2�������=6��轈`�}~q������(�l̯�Pm��d+��!Ŏ��d]p6�� ��'�G)�@Y�4����"w�r�2^ϥ�Agy�\�U�Ÿeí��s��f�t����z|�ڗp8 ��2�1���]U)��|���N�å��{��3.�w�G 8@�-m�1o�,s�3@�y�(qs���G8�M�q�eR�r7�6;��>y"8a�����|��<���΂p�q`�=T��FE��Uw�t��*�$㵝���Ei������o1��Wz���Zg@�b;�T�E��T����)�{�]����3�ت�̟��>���L ��Ғ3)`�j~�3��h���tшf�5x1��{��UA��z�;�'3$[�jK(B��
�v�k�.�~�;��(�.�c�DZ�t�^6i��n^����)�4��}�b�[�cWX(v�R^��$>N���'qWi��Ih�rMWn��XnE������\w@
ܦF��+Ź$�}�]޳i�2���F�-�L=w��D����إ�9�tp��/Y�oJ�ػ���ü1c ����?�߆F�<�q&�؈f}������#\�6�e��Ky����Xbw���,�k�������8���S���k��q�����$L���*�Z��D<p��:�f��NO��M���w����Q(�XOyTQ<�W,�K"gh��6t��B�`l��l8f�a�H�Šz�a3��&��C<k���S;�:���Y�'% hǇ�4���p�|ڤ8W�bo
~n�L������<��5td���/�����G6�����3�݅M'��/)��}��@���}�ݞ:7յ�oӰ|�S"f�Sg)�ܓ���Wx�O7���s-�n�� ��'��D��L�	~Զ7V擘����Gz�?�l!k�-LT۪�j��zo��yP���V����v��wn�*�S���"���]�;/iu�}i��N�����-�X��3u��[�e��O��l�İT,t�re9ZA{�y:h|ƞ�Eu�8��q>2��<>XB�κ���&��������E�����S;Vm��ʾs^:�W�`�]dB5Ү.�w����\���z}^q������՜����A �M��o���74�>�gB���`����URV(�.���A���OXʠu�k�T.��SO�:���t�K��4MB���y������������B�뷸�^��Px�����Ȗ��,�1���{}$���W:u�p���8�Jۛ��J������kX���c����t�7�O��1P��cGqV���R���˖��(\�m*c�@$ '9��ٵ�vi>�7�
l���ɲ<�ㆯC���ղ,�M�o�2��{�s=�G�����!�����/J}�9][5����k7''r�.HTJ_�;���5W�םݺ9��.3lKz���y�e�A�^k//j�i��ϥa<�%��t�L��n贈� �M$҂x��y���l�q��1~d_A�vN�_��7���?kk�,#�k].��v����.9�1r�PZ�ދ�q�~�Ԯ���:^����.v�oMl�n�V�k��\�0�3�]�d����Z>��ʒ͌��R=J}���z�Y:vT�ss[�9�G��vl�:�� <8-����X�<ٚ^WFѤ���.������Ǐ����r�g<1��)��K�=�#�N�/9��+*6T��]��ȄA;Ԑ����Y�fC���k�Z��d�rI����1�l�.�)j�M��!�fz�+ѝ
��{M� E�}���xǴ�6b8t�K�8���S�N�d3�wB�9IW�[�=B�h����q��+I����RO�G��[\^_�/�� ��8j��լ�kkL�W��y������G��zW$�����^m�zz��]�^6���T����>}Rovi{O|PF�t�U�9�s�����ՙ3b��֞�8Gh�+���ޖHl�z�����k�:葒#8K�W �;[�k3�u����;zDJ~�]3�� ��������7�[*_�r��gg<띗�̿_J~��uz��B�zLB�8�p�Hg��b`��2ϔ�oY��t�l�qD�gǽ�A\?�F���Cm����l/n��)�Y>�]v�U K�P�(�z��EluM�q
۴�}�{e��d.�Y�]�tt��hH����  o��iN��s���m5�A��K�!KUp�ǐ����,�ǚM[yזfc:6�{3�N0�����������;ߎ�[k_~������M�M7l����i7���"�T�
"Zl�Y������@D{g�iD��FɾJp$L�q㝟�mu��D��]������O�a�e���Da�B���4JJ��R��Y��î�i5+���&����n�0��=�(qˤF�t+�����Y���K�t��%
�Sl�����S�o�o��1�8���'�v��Y��3� \�b{v�M�����'��@��i���Jr�(t|���Ѩ)!A+�Cގ���Vuvl��M��3�� �<ޯ6���]1݆p�Do������/��x����4��]�y�O�7�{'���h���xk�����Mu�Z�q�OG�hE�;�!�iYJ�n.�r����'ek���Ǡ���B-�/t���e�R�B��w�yc�C�}��O1���VK�o�3rf�b�=��C����Z�qk�{���X6��]/Lk�����⼍���dҕ���&����O�{�j��*�S��gg�}�:�N�%���f1Vwr��ҙ�w��v��N{�qqqs�Nw؊�G	�7��)����r:��s1��t��f���ZPx�z�U�yu�A^�Zzy����3OL�0u�%M�&�;ɞ�Y����K���;\܏+e	w���?wU�����G2%��2��3�EGQ9�x�F�g���{�I$�T�����Cg��b��Ma~c�9�N�$33b�7��X4��l��+�#�%��>��tL�U4�+,�ãx6��R�q�+�gl��o�bz�*H�ݩ�U������	�ӥp�6@d��}iw�v�U0oz���oa�q�w���`���x�J��|�f�l�8��l��}Hdmh��{:4��m�8n�44�II���4���~a�+{�jعˣ�z������:�HY��9���0�ý�:�t����Ƈ��+�ɽͷu��D��r��.�Q���v�H��S�(4i�f�ǧc�o�Ѽ5�}o�m�c]cD76���zD8��n�౒�ֹ�/1,����G��L��N[��kHcN�vI����XC�nI�^�o�y��}3׋{+�|0�@[B�J�	��y�����	�~l��x��]u���q�m��P�'��$@ѯ�h��=���=�}��^@y����n-�c��*���YZ;|�|Hӊ�c�}@�.�����e{L��j�5m}�y�v��&B��zA�x�l�X&s0Y/�)۬	��Ψ�����I�k����m���7��.i�@�gB�.�0gx�b���o�mF���8��IZ�N�wm��~��`��qp�8���^��<�<�?i�Ve��$�D�W\���5>m^AG�D��}�R��6�X�e���!�'z�ŵ�����!lovLw@��l�r�3�Q�ж�Z�]I%��[K��yH�t�5�2_{X8���țEA�xݿQK<��-w1,�+���55g*���;��G:x���+	�ϧ��r����Ws/X!�����M�������1IF�HX�/Tn�D]fU�Eh���(t���醕4�׭��a�U���~R^v_U��Õ˱&�봌���:e��Ω��J��΍��c��X�z�2��7v�,�j�7	r��-��2v:��{4k2���q�:�T�{��Wc�ތ�x;gv���s��10�}�/�=YX�����j(���Mc�l�ٹN�D���jتm�;��&S����+M`��0yp��n�0�Yyr��{��<'=�_R@���Q��#��E�u�5Q'�3�5�gkY,L1�]�ӭ4^6��t�t�JWmn��SY�9`�#Tm�����~��z̝.Kbw�m�]ɬi3�e�['S`�;m��;/g(���F�뷃�v���"����Nv-��sڷi���V��Z|�{2ƺː��1ʡh>��%�����ӑ�Zl�Wݺ)�I#x/O-{��q��i,�f8#`s&^���>�6Z�T�,0����R<̘^wF8�&3w�q�ٜ�X�Uv��s�\�F�<����P�4#�UD4���V���`鵇w��4x\W�O�D9��u)w	�#d�|xV���׊*��Ut�\��2P��w ����U�0vw�K�����75u��X����nD�[ޕ�9K<+Z�6�
���b�n���愧����~sx�<Z�>V�2�)N�]x*-%��䛌M�M����ʤ"��OVgtch�[H%|�0��`+��+��ν涥���˪��ObЬN
��5����zf_��/qO�G�V�a�yn�
���>��t]�*7UT3pp'T�uf,r��%K%r�� Q^r�$GtE�zf[͍e�b��E�6�E������x*����1���Q�5����!�Ά��7��Y�#�ˆݫ���u��9V�<���gjs�K�u� �*����k��DE�q�3#D�c7���2^L�Vl
��iB��&QD6��|9��u����o���WF?���d@�<��[��V�c#�u���ᓜ܎��sx��o5t�;��]���&R����W�jl_S%C)�tӴ�ܭ�Mâ��ݓa���q� ~JՎ\��c��ݥ�iFʮ���0�e�[���4~�}}�,sšSy�3�lT��D���l��Yu(�� �#rR(�e���I-w�tah���sk*']���P��ޗ�n�Z	�ӂ��2P�E\���a�H�-q�ίT�pL�*��zj��L9�R�R����s%��Չd�i�:���g��X�gT�x��v'�۴�>9Y�l������RVĭ��o9������o���Ss���,��?�˹~�~�򧚵�����	���f<�2)z��:i��x�}:���u�]u�^�u׎�뮽====:�����Q�vG,�3�1�(���OZE��F�G��r���EE��}>�O�����u�]u�_n�㮺�OOOON����o�%H�����'i��&&da$�˔C�m3L��ey����䐆���_w9�=ez�.Yn��su" ЊR��V.y⨙*ԋ��$�~�֓Ш��䕕t�a�����O=�R�DO<ww
#7uȼ��Luڻ�)H����/�x^>�;����V�r�S�ZRR���E�y{��OW	5U��(J"_6�T��G*=S�i����=YQ�G�μv�D��V�9y�0�?;���P_�˺(@�J�V�^4��p��2{�sȞ�:=��ӑ�}�x��y��Q(G���m��-H�lH"����=y]V��k���T4�V��1����.�R=�{���^�@�Mh�c����yӪgve���ע��$F�M�T��!Rq&����6B��G8Ѕm	�>�:��OT�����Z�!��n6�>2S�*�-�#�w���t�����仇�r����W�ɽ�?�0a�������h59ikˊN��orKW:�o;��Zv�%��L�b���f�\����9wH� ��:�mF��l;�a·{;�_VY���9��.�W���޵>=LwY�;4��D���2aR�����DwH��|倞E.钩���O�֍�|���1)S���$�ٰ�&{�n�^����S�������흮��rxB�fش�Sf�t�L��3���Zg�Y����q8��W5�Z��I�����*���9���8�������q���8L���ҡYQ�14�v`=>7�p�%��8�8%k˝�;�F��E\�ɤ�7̅\����a����u���j>����s�Eet�Ng%�X1�0׷v��a�V	g�w�Ά`Ϗ�!A���{z:@��pTz�G��fڑt�5���M<3<�c
vn����
��{�W�E[�{��PS�W�����۷��Ϭ��[�oӓ��}�K�5q�m芙/�e֋�Y5ە�ٳ�9�SN�h�c���`��GW�OXb���,n��l�UG��\�]�PV��sk��>`^�*����^q}:��Z|�K�Y�ܑܷ�}k�t������r��q�{|}�>^o|:5w6�Vj���,g���}���n(K%�����I�.��l�Oq��������˹�W
�[@I�lz@�ѷہ��.`�q� 5\�{�=w]�6�0pϡ�p��2�ʨ9��7N�z[%��YM�S�p75�!���s䞌�K����n��c���7ݵ>lǍ�+nzl��qk3�٫���|}=Se�m�3]Ԋ��aa|;,E�SMp�g��[;�����T�!l�!F�ڙ�[o��H�q�����v�mYM��ٕ�����vh��#�,o��i#�T��I�f�cMa)O��zk�2"c��Ҏ�BS\wi~�6fg�*����4���q��S���_V�;CV���k���ܒ}���Ǉ�a�ۂ��Fy�0��2�ÿ/����pn�l�Ͷ����K�O����s?�s��Q���R�F�/L[�\�'��;g�uB0J�w��g�������G{J����e����t�w �&���Re$�'`ۘh�b���:�e��nm欭��\s�J*�*j��à4d0NW���ܣʒŶs5��N�כ��ˌ?��<�x��p �\��u�!��:�T;aH&���v��ڏ?H�gƻ�$O>�t8i���4�,��,��^k6����]���ޡZ
�T[���Ri�SG���ѯ7x��
�=�'���S�C�.ڽ#�roW	�D[4�Rb�3'_�3�15�:��i[�-`��r��RhE�ԕнC�5�Q�G^$���fk������d� ��D�H�g�A\X��;�T�o�ve�W�^i�k����ݼ�<	�k��5�"���̓4�&��aG7��ܖ�
GC4W;F7��ǆ��|�	PK����l���D�D��q�+�WS�rmv�%*\/�gu�v�)%leHK�τ���}~�����o���{����x@���z`��P�m�ۃ^YƗe�ϒ����]����ȶx�F{�0�Gy��i�A .�4�?���W���ۦ:�pmDȳ>+�Ӷl82���[��g��56�|{���ECN�c*j�q�QǨ���+:�Wp�7�f�aG,O��\܍�GGo��̎q\h5����9Ψ!]�ܜE7*E�K֫�����eXX?�������p� $���-���Y��L6�e6��_V��g��z̃��)q���5����f�v�+N�+ʷdu醑�Æmy��a��\�~�L����NFf����4�=Ǵގ�iX
�q��8\o�Ag��	����6_+6v���l��p�s��d����/ǺAʇB�X���}�zl_���E�n�W�,nk�&�6N؍�s���ew��E�
�{���®y���^m��h���=�����kj�]Oӄ�5�;�'�Ȩח6��B�C9���D{�U�u�f ��]1CGU�6z���ݣ��I��8���Êz)���wB	C��T9��Ů�2Zɶ���o_J���iO`�6���鹧��g����h���/yq���lޚ�ӊ��H���
��%k�]r;o��4�b���1��o&^�i����Wc�b\��:v�)X��^=�N�it��E��;�2��8b5 ���֖���n�e��%
�}}��#��,,*R ����Z�ޑף,؜�}����_\�9-j�WP�mt�gZ6�Mͥ+�p�б�h"'c/ �Z�y��y��p������g�%��o�s�t��s-W`�١o2���]U՚]�D����_��} ]��>kq��qpoqJ�(S���)��M��`�z�1�snY��Z�#���g���@!Β�.�ϕ���������P������X84��~�h�U�|�%.\�ӆU:�*��[�_���I�M��� Bʍ[e��m'�=�V3֭rn��D�aY�oGtv��#>Pit�%�y��x,�#e�)�H��dtnNV���h�jR�uw.��D�n�Z^oul��8������&�+�ם�E�qD#>ٓ;f�ryK�ťK�����[Zz/:��6��p"����C��06�V���������v��^���pēuE�0j�5@��sJ���`+�k����\��V6LF��*��8rH����/�ƃh���0����"R����#Q����]1v�^�^^4���J�U�{�Ub������/(s�`�t6�<v������[������/Y��9C�}Xj9�oO+|_w&[s���;^���X�Ί"&9�0�8�l'6���!��N�x�o0o_
�����7��窕����mO�����t�Cx���;�#!���:h9�$�t��Z�V�=�M����9��Ջ�{}EO�`et�b��K=�
_�Dj����VnNp�,0g`2��УdU?�r�Z��N�%��3mH�e�5ު��FFM����-�,�K����3*�v��૊�GOq�@���m�˷`�f�TĹ�(7��wv`�⼌��z[-����Yq-*S=�ْ����k����s�ߦ��<����g���m�3�;Vr�s�w���~c�67����spn�N�l���8o���4^�%���
o
�/���:vW ���<�z�+�xlvwhwg��^à���Ԝhӳ�jM��+pT�� S��{h��u"���/�o�J��&.Uhs{�ԛK��̣���'9���v����鑶�$�%4���,�È�������}�L��x�}����u������MǕ�s/�]��6n`P�*(U\�h9Ef[ǵ���X��.��<'��	��O�:��v�8I�7^�q�c�RZ��p)ik�X�ے��vco��.�[�";�9�2N�׽ja޿0�y��Wb��_�3�v���?U7��G�#�N�ƚ�JJ��o���ŷ�T�tN�.�����3垷�����.�ۊ�S���Ih�'��]����þ�K�J�
w�qb	��๛ݝ�-��h���M���եx�'3t;�oq���!���Ϡ����[)�ő�b&�v�����oxBY�0c�u�v:t��p;���� qٔYz�$���s�o��z��i�t�&�O�����>�r� �4r�]��yՍ�[j�;�q����`��=�u<0����@�Ӵ/H��2�$��i���Y=�s���_ۡ�n�F�s ����&=�P�K�N5%zv"ΈǶ�u��l��B0p�M��6��f�YzjL�ň��K�e�K�A2&������c)z�׏P�ҨB�ުG0��E��t/�(����x��*�a��_Pj���״����k�����[P��a��ħ���>�C����G�j��T��"'ش�4+���;���B��@���#�f�˶@^(X��R�s�Ǖ��OYN�Lѻj��_���{<}�/ue���,�s��{�un[b+���	@K��n�ݘǵWf9��1I�u*��4���T��"����+H�����Ô�6;���Z��[s3�UwVN������f�K���>0u�c�ǫ�m���%q�xbor�r�y׼6���9~�*v���`�CK�
�{�Fa���+WM1�0XMK��<���tn�v��2\�$���R6�e5�a�֕�G)8���hR,��j�li4vo��Aa*k�V쎽 CH��8�P�_�9�ŗ�3&w)���
J���s$�n�;��uq��Lc����,2�{��²͒.9�{z\ED�gs��s@z��{� �v��t��wHn�)�pZi�]ʽh���9G�6�@*�P�]��h��;���޾v��ʭ���7e��=kd�!��3�<+ꊴ�`�wE�w��9\ҳ�m��w/j%Q;�W|�mkM#l:.���"L���]�}ڳ�7�����]�|Ⴧ\6�h�E#@:r�W�
gS�tժ57+�I&��%�s賏L������(��['5}����w&�����U����b�trp�������Z�_U����D��$пN}$�qwR��c*ഩ@�n�E�e��%��.�&���`������� �������$뮼�͜�EԀz�k�d�9������5e"b�6|��@�A(w&տWc�o�[��M�{�OZUޠ�����my]�4�����Lb��5��p����Rk׻X°�Ty)�q��nV��M?]�m��a�Y�33i���`��)�T�i���m�ø�$��$�t�'�����d�a��8
�14�\{$J(��m��	����mW�{z�/��3d�8U9�-t�U���m��7��j.%Q�y}�7:�-�(�o@�7)K���+�G�a��� ��E�n��|�<��#<�s_�5������_��dv�豅��(�/r�y����?No�Kױs�	�D���\{�t{r�J2 �gq�y��C5����X�{uxLS������D�wfd�,ݪ�ܵ*�r�t��vD��«M����Q�ϳ���s5�zD�ˮ�j�^=-��5�x����ƕ�����a��
gB,�] ެQ6�u�y������o�.��T>+�p���߫#	%-)wT�U��j�2���"����{���;���(
�U��05uz]t-ux֬ތnK���"]d���D��;�}�\��n�٠��]}�p���-v��T�1����hi\�@o;n@Ӑ�ޣ �g�;?c0'B�
�=�1�J�2[q�mQ�ӹ��7��y�'�noG��A�]>ȧ8�@ �Q�I��V�Y�<�S�&�����ϜS�s���=��w�Eet�S��t��-�n,8����
v7����e�C�6��H��G�-K��fڬ}�>��-��'L7X�,��y��FZ��[�இ�O��yWxګ�T�|(P��s~w�q%�]�D�/Pd:�P�r#�yb����#_xGo�\Kt�m�p��_gl9��Ҽ�R�ݝ�X[?�uz�����|��?��ٙ��R���|-������U���4#�ߏ:t%�"ZG:Z�-�9�<��w@�7���Y���RTѲ��Ʈ�����BvWOa�{kWT��X�!���w���zv�$z;U3��o�b�����u�
������6�0���,�V�����V8W yZ�A*L��v��E��>��I_dUd��{�U�#�=�J=
�v;�lk-���;GC�˫��>yWF�Zh�Eɑu���n$|4F-�.mE�n����N�<e]osʅ��ژtK�7d�1V9[���qBRN���i"���|�=њ���8�!��Xꐘtgna裳� zK͛�ʆ9��Ejc8�V��u]b��Hl��(-�����F�La�F��Of��[�Q��!����ʺ�4����<j������]b���:7�GMiL�9mbj������s>\��$�x����i)��2��.;iT�}���O�\BٍE�9[F���Klq��e�|+��_t,os2�@v��*��B��ɬͿl��o��R��.�5k�sq��Za���Ci�aY�
T�8���դ����v�#Cv�#�=F��=v��v�J�49F���XEZ��/��٦�V��{�����̝�܆�1��kO`};�}��2���a$7�:+r�"f��`��emJ���T�n{w���6Ic%mKv��H��.WB�z�$���ݚ�t)����8�vj�~�nX����^������qݪ��q��6sT��t�1J��L�1��}�w��\2SQP��W��U�rz��V�(���>�?˓��V��n�|��Rn��˺o:����b�d�ֻ���Zގ�p�z��H3zv�T3z���;&ⴂ\���;1Οt�I�u��'��E�S�m+�y>����I&�YE��=#Q���F��W��έ]�B�Z��jV��������J���U4nv-O�]��q��;S�Ƨ_Y9�R�J��-��0<��:��33^h�n�=�Ϧ�]�,���ϳv��N�����Dt���OywW*�P�o�f�-<M:�:/!ӳ$���W�����kM�;{��E��r����u�X,�}T��Lu�V0�_u�>�"t����nol{���{��-�h��И��h][G]n�F{�1պS���U5b�p+K�0��㶡�Jn,��j,�vūD+��T���e�S`܃M�'J��(��0F����Zn�!�Frk�ZYl:���9�(���^gd��9�n��|Se�J�d�ͱ
�cg�m{ڔ���볫&��m���u��)�����o�_v��^��ؚs������SС���\.jj���9^��޽{�'
���������q������룮�뮺���\u�]u�������~|>LFLM%�f��k���*��&DO��iY�\_�ݻ{~o���w���뮺뮺���u�]u������7�����EJ�4H����s�����P�yF1��1��MݙEZ�y;�|��P8}:"�JZ>\�J'P�R�z��+�sR�9n�zDLҪM�}��G�B�TT'��TAEf
�ԁ��l�Rl�U�ܨuZ��s�1�r@��9���px���]�ʼ�Քf���ۤ�*�k�9�($��������!�Us�L���f-
$wwVf|��N}|�(�(�T�z��� ����P�b9�׻�Ϭ7'Ե�r�#�S����c����V���{L�9��p�B���UIP�$��ZE h|�~9����%Φ�U��Ş��������h�������˰8S��N�)��>���X���r��٪y2�y�����aV��)hbd8`��7_u6��xw}����m��t��l�T�����ͲmU�l6��|cvr�� �==�{�����ͧ��ٌ$1;u3
����@�9��x�Y*{�Pl��A�S���ε;�h�ΧN�8u�y�뙼a�j�������5��&�)���3*vY�N�s�l�N��T��<٘�����c��2c�z���%�}�n�$�f�ܓ��%?�KF i�o�a#N�Dm�B|��B,Zy=��)��k����{�_�j3d6����f��]=�K@�u���Y�;��R�Z[c��vϻ�l���&��CF$�hz�v��Vu��gp�5��JK�F�]����Ǥw8$��c���!�34�*��N9ao���#�e�U�Kx�����z	o%����'�6��O�۝�3(*�h�vng�eq׽3{�L!�]����� ���Ĉ(ѝ��oY�@鱜��Z�6ʮ��ُd����c�L���᯻��v-���u�n�wq�,�
��Hi�w��}�K���y�v�8�N�u�B��$h`,�+��v����^��Du����]&�霜#4�ͣ�:�����V�&Z�7�$�0tE�weB
��".�/CE��.����E�R�%�����}Ce� �,G �n�J�u�9��ۺ'#��F�/Rp�A��Ƒ��UW��Os
��� ��2�l~F�1��6�ޭ�Ύ������'͑��Ý.���T�쵻n�"L��3eVfU�:s�\5����GT�O���R�jK���Iw]=��3�VL�� VG6ө�q�d��4'�ǫ�I�ވ����{��h-p�[be���7���ȡu�	��>�i����
r/�f��+j�>G7H�yR��r�L��{M^׻����e5y7����y:� 1v�^+K�)4�B���0ͻ�Yv�[d��:��T�U>���Y��p>�~щ�+`����LK0z2+`c�]m�`����+.Z�0P��ƚۧqd+]�X��y,�+��5OlI��	JB�K��D��b��#�=̮h-\�q�6����)H�Ў������w!u|�d��2�%�z�Zp/w���sc֎�ܨΡE��ڜ,ܜiAH�*t2�:9IhU���-�LL�w�vg��ʕFoe1+8�ye{��W�]kdcG����ǜ�>�;۷[�/��.��P�M�Ӹ���c$��w��UL�ݎ�J���5s!�h����^�r��qe��Jl[���D�W��c��w�vK՗�s�'3=ZY]�v�/�<*��U���tԧj�n�w��i�~�v@�80Y�g��~u!$�Dּ��Yg���<�0fJ���<��s�Tt4Vtm�Y�/��nǎ�z�M�M>�� �<�q@��b&L%Z}��'/8C�	�:��k� /��ݦ�E��������MB�&�ʭjӻ��P�!�������[�W��p	��J������fV��{㞁�o�mB����E��Tw@X�x���:G]�R����Ul�g	�ʍA��F�t	���r�p#�]�vz���k�ו;q�4䅧�k��T�"�8�{�(�5{ʆ�U:Z�yuu�ǭi֦m�o�CR�0�ݖ^X�!�+wv��4X[�G[�,�5׏#8��`Q��lJo
)�y4�����Ҝ��Ok�R��ے��/h�C��>��W���r�t����T�ζQ�.!ĸ�a�[^��GmU�H�q�q���_L���V�ZQ~c*V�Hd5{�E�	˰ohZ5��Ӵ`0������fo)(#���-o[vq��~��ա%��;��o���5��uMV���e����I��?eG-���Uܺ$+�gOq9Kxu7���y�[�����&y�(��1�z!G�FJZ|��`��VΦ����~�û�������T�w��
�8�d@ˏQ����y���ҿV��&�-��=��3�IC:�ʾ��=���sW�́��ǯ2y��;{")֩Vu��7}�sg������r�/�4�;:ƄY����v���&���L��]'�u��Ҥ�y�7�ױO<<5��5B�¶=Hxe�[���E�������O8��S�=�Zev��΅a�ŗ�R�2���i�J�A�CO�I��rZ��/m������L	�aR��T弓���7uɞ�W���8l"��N�6���.qy:3��x,cK�;~���w�d�i�\�������|�׼��gj��˛�t�m�/k��x&�N�^���8xy��G��r�o�ȁ`�Ug:s�N3���
A�J�]�ʍ.B�#����p�l�ڭ�톐(+�`���]�V��w�Z�	L����깮�ӗ�/W�P�s)O�ed۪��#�}`,t��d�S�*�duu3G^n�4-/<i.�P�gݷz��U��^�(�x���[o�Ě{~5:�cM���w���1��c�;�*I*cV ۺ���:�龧v����'o����
(n&9-b�P������lǦ�60�����l�������?Sm2���d���H�e���{�,���UtL�d���x�my�C{�^�`�nDB�cv�g��ě�-;%�ry�#w.�Ѿ�e��qk����q��+@{���}�"#�n����%�U(R�o$���4ssv{�G��Y:)�=��3@�r���e�4���$ƢB�Sbç��|����;�r��7��9E�ܛ�iH͓@[�x�`�ѿU�D��i�1�%eq>���E�ɷ��nؒ`�N�S[�V�u\�m>�I4�۬��B_p��5�_�+���K^y܎�K�1�nl��t�o���='�3���x~�+)>��$gS��H1Y;A�7������x��ul��q]z㌚[g���w����a��Y܍�]���ړjz���67n?w��v��6�윳���X��8$�+ML՗���<4D������c�~	е��<��{����˄@.F�<��.��p�����~�{��H����W@{��s5R=���nD�_]:ޮ���d�׮=X�H�Y]>�n�g��($j��w�M�}�0�}��gg�������^�dW)U�ݍ#�Ew���46Y�
�?p�,�ȴt��&�7��ܬ�6hT�H�TqU\cٔj��]������Y��}���X�����e,��Wu����)~���U�.�vR��ٷ����{�
�1�y������`���l��r�b�W�2��&�ޜ��ڽ�YN��-�����#-'�J�̂|��j���1!���;$��"��^�Q�x�Ky�I��C����ˢ>�B$B�>�I���-Sr32No|��+S�ޱѷZ7�c�Om.,���%]z��81w����\�1���#����z{��'��ˌڽ��r[X��K6����j�#�PYl$σ]`�u{��ö��tō�WB��1��*��5i16�*i�r��_l9���:2��3�4�EBj�B;
�=t��a�{3MX�R�zL"d�VOD���Go:Nո�6Y3{ >�%���ɼ�m^�a�1��N�`�xSq�XJ�9��|�*�hQ�9=�G��5��w�rr~�s�"Z"fs�3�#���绎ϖ��7J���/u�m���)6t���;��=�-`�2�77���h�'J���ء9�uy�d�4�A��g�fg�;����"ſ��wW��P�e��G_]G�`���q�'W�����t9�Ft��_P���62�Qd�a�m��vY�"�9 q\'����:EF���e��<�}�)nڋF+q���N>��ʸ�������T�܈�w���SL^ڣ�.��r�zu��8�Qu�
���Ń9��ZCYG���.�k�J�ܼ�C���m�ە\�^AW�yU�íק9'Nu��<O�Y����޹��{(��Z����Z��6��˛b${�SNqv�-��/Xͫ��=Q	���j������ze�w+����A�g(C�L�� +�zGMut��m>���.i�Գ:��C�H��Q��ѽ��O�}��&<��� %{�)�w��k�T.�{a��u�}����w��*k�S��R�r���>׹,��W�=��h;S���.���,�V�fk�Q��O�s�~���n�vO�(���>8�6�)�V��ţww��^pm�=�o������:[)�}�P���:�|����<����y��I�ޣ��;�{|��+��1�-�P��#��L>X���w>N��(a��_��r��6���bI��.���WI�ڱ1�����}��֦`n�ɘ'w;���wm�hv*�E�jZ��նWL����:w��ƚ�`}�}B+��:��{�fL�=\w�u��g����nuF��g��$ƛ:v�*p	�RR��/���{��A$��%r>9w9�}��}��_,Br�}�ɁV8J/(gBw�8)t�K_����w=�HT�Ցj���%Ț�ju�]y��r�m7�W�X��ğ2>�b���U��s�
�r��e�Z+���L�>�ˮ��(���K���׵-�s:v��2Խ�颠8?{�||�|bt����32����T�	F�����M������33ƿ(��>���[֢�`ߙ|Q���` �c�	ӢM�A�c��	�sʦ�9t����{�k�8o;��fž�'���#Ǜ�x���s��t)|�Gl��+r�Of�bk�����g�����gUw��l����q/�"��ms_���C֔��σb4'U�P@�5O�)���%�Ú�L��S��;�v�tx]6��8��,w5�PW�"��pW�9�;9s*�z���0H�ǽݤ�˟K?_�2
�P�>�� ��[C��>��+:�:�����$})t��P�dg5ުu����s��X�we�B}6l���^u�3��T�u���.]LZكg��u*��\���z�zu;��حn�9m�z��ݻ���᳈�>&y$��A��wg_��}�i�/[�Fdj���m`�u�ϭ
�;a�(�:{ �h;�C�,��o]�7���"[ٰkԜ 9��&�2��{7���v9�˯#֭�ʋOm�;��#g:G0:�u�K�}W6��WNT/�����W�}Ps[����7ۻ=��3OL�u � v`��u���T��U����a����3��	�4�Ւ��`5ϡ��-�A�N�(�Y ����+�[=]n��6f���Y�8����K6Y��R#�n�����T����\�&w"�|;d�?`�7�U�6��1�7�f��a�.hh�H{����]w�_{�L������}ݽ]��}5̡�}>3�Au���)��_>5{��H��w�h 
��嫟ew��v������ӑk2������n�f��o_�t[p1�ϕ���K��\uҐ9�f��H%�GV��O���Q�e
<*���!���,��h��t�'�@��	�c4�g������z�V�AYf�[�c�<�_��h���U��{_*�2���mj��f����=����o�>�Ώ<���ÿ^������/��W?�Q�����?��D?�Q3��8@"`z�Gy��0�� �+� C*�ʰʰʰ�2H2�2�2� C
� �2 B�0���C ʰ°�0�@0�2���C*� �0�B�� C �0��C�!*�"��0��� C*�+��+� C*� �!"�
�*�"�ʰ��ʰ�0,!(�(��ʰ�2�2 C(°���C*�*�*�
�ʰʰ�~�����P!�a�`VV@�P!�a�B!�eX`@�U�!�a�eXY� ʰ�0�0�� C ���!*�(�0�0� C�(��°��C(ʰʰ��0�2�2�2�0��°�2��� C��!
�*� �2�0�� C*�
� C
��2�+ C °��L���	�qUBPP��T `UBP�� aST��@9�rE �� db BA@��U@�E@��P3� dAbTa� `Qh`had!�D!��P!��P!��9� �a��T��H��Q!��HhdRP���p``B eX ����`aX@��`e^s�<� 0U��`eX ��``XV9�8 C*�*��2��+���|�����EQiPT�A
�?����~������|�������s����}�#�~����O�v~����o��G�ߟ��� _�@G�����
/��*�
�������@�П�_g�O���}�� ��{?@�2?���C�A����~���	�3�����~�
��\UUDbP!Q@e�%QP�P�A"P�BB P�P�BDP��D %@	@ �!@@ �$I(��2 � H���*� Ȁ� �J �H� @$("� �" B0� H� � $� ���$�	(2��� ʲ��0��J�0�"�*�~�������ꨈ��"P �P�%���>���?�?�(>�����?a����@\߁������}�����?��H�`�lN���ʀ�����>�O?Rt|�W� ���?2����?���å��<� PW@��������}/�=����00?���N���z9<z�* 
��I����uҠ ������1?N����t���?��?#�|���	?��C�C���J���?C��?��* 
��~ãC��&/_G�?0,����~�����>��J����g߳�LP���?W�8��|_�|_�@AE������� AE�?����wO����O��PVI��T�C���V` �������7�>�|�6̰��U!�Z�Kf��жZ��֤[Vij�ٱ��ֲ��M�0l��kil�U���(HI��j��ڵ��f%Z����H�5!kd�5�Yv��di�Y�U�5Z��f��Z�m���V-�kc��ٳjlښ��I�jm���6mI�.�ĵ�I,���Y(&��zS�o[��m�mV-kj�ZZ�m@��mm*kf�j�Ul@ֶ1��(M�mZ�d[*f��-1�%e�f[a�l�fa�Z�m[X͖ʹ5f����t�^۴�`�   �^���]�s��κ�mҫc�潷� ����#�5�W������՞n������8Wi�Ӫ{����u�iVv˽l�@�ݼ�n��=zR�Ým[m���ZՒ�lլ4:�   �:(P�>�B�����E
(hhQB�qáCCB�
%{�ۏ�S[��ٯg��c�:�lol�o9�ڞ�Ӻ����[���Zq�z��m6���q׽�����M�҇Z{�����Bm-mje�f�f*��m|   ����4��s���A��9s^�y蔧Xk�{ۭ5�������z�r�={���ݴ���+ս��Ҵ�퍡�²����vޞ�0��˭��H �%�U�h��E�Ym
�o�  W�o� wޭ��ppZ7{o-��Ѡ<��#�t��8
�WZ��=��
z�ѻF�NW��j�Kݧ����Ƀ6m6��ՒA����f�   w��l�}=��=+��0S�.�k�b�UV;�Kn�:����P����]t�v�١��� Q�\���;հرQ�V�P�&�[/�  ;��
�7I��u�0.ڠmR��]on�7+����r�����=U֎�]װ�z�z�M]���Tw9�=u@�"]L�ڵ��k[-��h�a��  �P  竸 ��@>��o#  �X �畇J ��n 9�p  =��  6�  p��Q�QM-�*՚�V-[�  !�@��}  �^\  n�o  n��  v�\ zw� �f�w�pCA���� :C  ��1&e�Q�+Y�����  ;�� ��� �>�<{�  �v�  M�� t��Y� �7  M������  ��u�=4 ��,��T�E���f����  n�t V�8 ��kp  �`�N�4����� ���K  wl� ���u��5wZp  > �~@e)J@  O�2JT�� �)��	IU ��F�O�JJT �����  $�RCJ @����o���~��_����7_�:�p�u�R���d�a�\z�N����??7����{����������1����m����v1�cm��c�����6��m�������?�c����yG�(/�À:�x��AV��[�ټ���1�;N70YJ�{r��'5���b�1�~7�Ls/E֪h�0\�P��w����51{�Q����y��̑FՋSk�d"Z��(cܫ�A:T��#��C�3�K���U���aҷ2@K �X8�h#%�=;s5=�t�1'2 
FJ#rD�V����T9r<�o-�6�K��	*��Ҳ�BPmQ�`c[�pP�B��%X�$y��\�6u��n�,b!S��nf'L�Ylh-�ͫ��t������i��AӅ���V�u8�,rk�cdm �q��u�y���j����ʽN�N��ԷYE<�g�&⚄�]���VN���Bn�؂S���ě4.�aL����U�2�[��q�8���uxqQ��"`��7J��`V�6<�u�~v��'W�Dݺ�:�ی�,����[�6D ���)ާA�r��F�]݆hTX�Ӆ&5�ț-h.�B���6;X���T�KeM�h\�3)*Sõ��2�(����E+qSȎ;=P�ݭ&��%:b�e�@����˄�M��R���ݝnJH���!n�J�Z֥@�c-��Ȕ�)�&Ѳ,�FI��<�i�.4�m���*Q�X*ff��d=U�ӄӴ4e�M}w%�I�4����A�_McAf֊����ɹ����,�5�N]	���8p�1�֤*H�R;W�j��� �kh��vGNe<�K�'a������������V���r�%-�H24������U��Ђ������0ڕ)mȄ�C�Fȹ�L�Xv�L�E�*+0�n 4�[lٴJ�EѶѭ�/���!��wP�Q�n�]�7L��CU�M���܍��VՕ��+5���1{[� G]l��<�a��Y����R�/K�Ӻ/F�^I�+�֍�k4�mS��cU�(e�.ֳg(�8�ڻR���^6�D�z�̷�S�fX��ee�xb�ث���MlkrVpn
���nV�� 	�K�r]���� ��V^'��A�G*U&�
�%�[�W�!d�`�l�]����ӽ�c[���b[�es�����t�.�sE����V��`��@Y�лr�R4r\Y��G5��,w.Z_:���x�` U����<.3�K�՝�4F@\�1�LX�H"��^M��T��4�cQ���9K!{#����Q����[1
��w	���4Vb��fhaV&}2�'t��]�-��q9o-����;TK[/v�V�;��1�|�M,�MâL6h��.�-Mې4r�;o,܍�K!�ܡQK˦l��,�uD�b"�c$W(Ya�jI�Uf!�-(ՆU�l$5@`���F����4�&(Fw2�J�GΉ��07z�K5R%�B^l!���-���2hU,�����6`
[�6���A'e�D�8�Zm�j���+�,TU�����N#�ڕ����E���zQ{���P3��L�f�Xvtxu�Q���V�Fe2�X�,$�c�v20�Z�Z��)�n
0˙�M�M�;	t�nS�,5�o/a����,`q�z�N��V�ͻ׮����im�D�;rSf��b;�镭���<�{Є
df�N�#I�m����#��R�{4��E=��Or;��n�U|�;�k��ai�c��ir)*��GDbହY��r2��4 i�u���WTr�ud&�2J��=E�dT�����hB;�m覥�rI.ڭi�u�?�^Ų�J���R�
�V@����SAQ��'	���e�Gق�)��u�`��F:��-���Fm�F��{�II7$���@c��-[<�D��J�m{{���ɨ��-��q-�:V��H�����qma46	��/��!�;����Gn#��4�t������HJk&GD�4�#,m��(eMJbc�a'+$r|�J���q<xZ����Sj[[�(�]GR8cí"S/��X��{��x�m�7'$9JE�oY�7���z�:�Ŭeݒ�ѭT,�";Ǥ�C �O&Y���-i�����b�Z�[*��h�� -�n���81���eD!�W��%۷77iq�v�b��cnl������I�cɚkY����u���P��S�)���!���u� ����r�������c݂ۖ��A�UB(��ϑ�4�� ���ǻ�}:�Mj�%ei2�<6�F?���FI�1F�)TX�[Sͧ�� ]�i��X��-l:rj�1�ۚ��:8ڦ�9�e9)7&�Z�w�m˧���r�̒g�~SsnW-�#1�V���h�	�M�h���-^=�sR���a�Z"iT�x�[6�V�@���PzD����d�l�]1X.���/+���n�L���dk߁���l��ڷ� ����ޭ�Q��^& 2��12,S]h��n�(�r���sD�p���E9R��ǹn)�D&n棿:� �p�ykaQ������抲�d�n�<Bci�(k1\�m�z�Z�P����;��i ���of)H�!Ć1WF[pY^�e-!�Yy��z)\QnA�.e��"�fPi���:��#��Yq喠�,;V֪���`��m�`,vQ@��,���5m<���&���&�%ǅ;��[d*�:�ۥ20f0Bn�$ Vbm����sL�����scЅ��@3&C�8ժyN�H}�Pؘ{�
\R�m�O!{� �#tG���^����aۭ���}[V7M7`_ثM+ǎ[�{kC̡v��yW�H���V^[v�P� ӵ�5Zc,�$�Uu��λ�!���U2�F���A_Kv�]91kM�Wwf�SX���L�7Vˈ ̥(���t��aK�t8S`��WOZ�����2�I�r�!��lt�43�흧B�n�wRL�/D�GV9m�`K��][9Y���;K(U��R�tǬJ��@;������8�m50j�Է�r�6
���y#ʍk{{�e�DB��3 �n͋!Ii,�e�F壷/]d��,	wg%'�E�$w�$�fb�2���e���Stt��CÐ��oA������]c9#�A�q�Ej�Cj�UHvf=S(VV�LVf�)���h(�+���=�*�w`#|5'�fb6DnAae��ݱ��K���]*h�� ��)�
Q<��#��f��֘M���,5#��%���Rd[d�n�nQ��촷#wQ�jf	AM�f��X�e�ܠޡ��Q*yZ�0�(�G.
,���od`�AIM���-�t��������<�{�BV��K*�%�1��P�{R}�%��&���G}{"��i�~p;j��s`DS�ଳ&b�/�7��� �E��Ɂ����o\�[X�����P8���I�i4�	��EF����@�B��Z�hc����3�˛V�\rА���Z,��FQǺ)�{��2˫�(�2�H�õ-2�%��z�����R˒�=��^���f<t6R3d!۰f�j4o*��f!t�N��Ojh�D�L�p�9(�(�k���$�cIT�pћ3Co.B �b[tk��]t�$��x �#g���t����w.RGd&ӻ�eխz��s0�4F�\���p9*�w^���3l�)��Z��B%%&����[O^�p��9.��`;�i�]�*�hU��5h7`
�˚�D�mn�=z��*�7��ŭ��"Y*Ij���[��b� a:@�m�p�Ӯ�����5�r�y+a�JՁ�g�4��kYo%3$bmk˴�h�u0�(��R��-�F[���j 7#ъ��Ol��d̔�).���{n87-��V�_!i��h�v�T�ʷ�n�lȞc]Un��m濥�D�~�Cd9���ch�����a6��ō�țӃ 9S�54&*��1*�k��s5LwA��T�m۫��T]��ޫ�NFj2c�z��0P�%�y)Pq�A¹�*�j[l��q��M���*�&� �	� �9'L�g%��ҷ�ƈ�Qc�nZ���67���1�ܦo�"�����A�{�e�ut̫� T���#�`����N�e&f���/�8-�w�%]2l����#	�g{����O������nKI�m얨ۡ2���qH&��R�V��h�	�G+66�PMؖ�)%h��ۺ��ڏi�d�`Zs�,�n�J��Ű���IÒ��y��ÇnZ�f�W٢Gב�ܤ�����,x�ss�*��p!����v�݃�r��jE%����Ӓ��H�3b�]ӈ;`􋭲W�㎅;X��V٩����]�Z0�ÖoY��l$��,�����;/^� l��ǁ�9��
���1̧��uf]*���8�R�M�ܩaJ�τ�K�Q;�oP�6�ZU%页����J5p'u��Xa�ւ�fĦ��(TL��^l���0�j�Ui5��
G�ej��o~4�݊�n��j�k�A�M(Q�Q�)уsm�E��i=q��7N�FiMC�A6������\	�I�4������F�����b(q�%�y1�h�X�QّjQb�M�����dJ�7���V����SK�j���>$^�v�^��!�kC�z�ټ�h�4@�6p�*�:b��Z\�.ɬ��T�Kz�KU���[ǚhJ�j"��u�!�'�a��16�$��qf�+M�U�[ǡ�5z�R���d�t��yo~��yK7n�%G��q��Jy�h�8��X[��-��ISh��\3q\9��.0�Q��B0���a�e}�Z���ӱ�6��ٷ�w7-dkD��v�xl�]c-�l��r�Z�D*5w�*\�ZƝ��YQӑ����u�6��[�Tv��"�0\�MU�D�ڟ(ۃ5[��b
�,*�z������"}/e9�
���+7wi�p�����V��[�3i3�0�d�h�PnK�m��g���/��˧��9KE

+3c�p^+��v;�JV&寶H���r��@c>ܺӮ���͡N\�b�l�0����U��oHv2�XB�a�l�6������ĵh�yf�j��	V�	ZE2�h��b']���CZ��z���V��F��efeh�^�K�z@:�A�R:�m�U�/4�C�{[(|/`n�U�@�Z:���܅n��J`�Rܐ](�ZÀf�9n�]� �݆R˸Z!q���Fi���S�2�\:��5�Rn�b�xv�d�
%�7)�N�8.����	)��i��a���lV^V��giS��Ϳ�Tj`�nώ�Ÿ2�%x�0���� ̆�E�wu75$"f��:�Qـ�h�,8��i��+I÷�����Mt���&TTe�mX���ɪ�f[�4��/Tn�Xv��8�ֹSз<Vb�m� Fn���[J���&`�*�*�Ŭ% �C�,�oX�1ۢ&��#�SŖ�6�yJ�
[,�[�.�R��YiU�{���m�0�$�����5��3yN�/3fCE[�QԈԂ��R�Ea�aL��# U��[;�s0�Z&nӏ�	�1�����fcz�iQƊ�FC�B�p*��Cх(�AP��ɠ�Ƕ�۽���^�B�4(�N@wl7Y�y�Mj����Kz@>��ģ�P�̒Y�jM��Vi�"���b���f(՚J	Q�d�wq��X�]��ݩp�,X���卢�Ç4�u�`��z���r���ѭ5���v`�W5��㻧yNXw[:`tj� *�ٌYIԚ�D'MeX�$�lK!�9��:/�5�2���vsb�犛��(jK�l|�P%(��y%�$C�k���@���@-E��-	x�A56�Jqk{�O�p�ʷ�F�E�uxmэ;�f����j�x�Jvh���{R�?��چ���b�R(��d�wOm��Q!��mYd^`��N��N��6ekR�1����CFV�
 }�풝@ٷVԗ,f#U��%�E"FD��ј溚j�qR�m��
��tkB����K�!�
��sm�:i82�����XϲëpY����l������i��.�5�n��q������.ؔ��@:�^��/V漼��KSe%ZU�U0F�EW%0r�|)/�5���Ek�m�䳿@횵��������rk�5�YR�֗
�D9GK˗Op�CV[�6,�"��7{���{�h=�h�5�gq������/�W�v̬�T E��u��7f��
w���}�[s�?2�(�j�^��
	�����,a�Qo�r�B�4ǚ�]�A�RL�Ͷ��tq&��l늅K��w�[��Cv�H����f}z񹦣[q!^���@�ݼN�;��x�;Xr��4
�Zvd
a�aMH,���M �;dL��fEz1�Qm��C4>漦C�F-���sͬ1Շ��ڇaF�yN��1�d����v�����ܰ��A;�W- ̹��n.��OL���6��P)K[��o!��BA�[4u\��T
��!�7^�s^]��T��������2����{M�۠֙[-�ݼ�,�1:`F��KX�[��YxFp�+1��`Ѧ��ŷ� �r7W�ѦD��L80�Q@�UL^&�̏E�aȉ�l���h	h��q�t��[�vd%�A+�T��/1藕n�5���+)��j�\L��.��>�+�/1�ۊ��Z�`�zuBj�=Vf�Yxdq��V:n�Wܻ`Z�������l2��L̻�R�e٨j�0�$�z��`e��gE������2�`�"���+�#n[�jB�'W�:;�f|�K�����Q.�ws6�u�v;��BsnV�����|�u�՛�������;D��dd�sҭ�/�{�'�Q����ҁ��aͮ�|����;��v�ӡ��|��'W �%��a�/�W!U�^�B�)Z�EV�ӳbu���e\uь�{g�9qLۖ���F��&9�q�zP6�Ť�c2��zxХcz��5��.�m����G9�%75���tJ���]V�v�J������>�e���p�#;��a��h��S�P`���͚��{IV�L��Ѱ������Y��+�8_i��=�G`�G;މ.����}g�8�ޫw�-�s��m3)+�c
�J�ey������+djnikM-�R�J<��]�̫U��: �3jn]�3f�l.�%Z��EDK�.�-����:5�2:]��&:�~y�%̖ɝy&Ad��Ҽ��{(�v�J��)����7©5��s׹i�b;�ρ�8�$k�v��&뺴�mn/L����o��Nu��=t+4��'{�Q���:@�����Ζ�y[��[�ls2��Oe䣗�m���9����ۀ�8�;9�Β�ߛ̓�,l���n
�%����c�թI����peMeݎ�,=\���poM��v��LL�8H��G��$ű@.<���ǃ;w4����g��\v�kz;/:S+�b���G���l.�v��z�>�$��/��j�KK7�#w�{�Q���'r�΃��m�fJ4`���8@�w71=�3�q�;gqq�s�LHVnM���F���7 dsP�)N��lRyq7��eq�|�K��kK�>0VGv�;�����)�ȼ8�!���vk�����f��/Fv�eLu�0�ç2��%É�m�v�՘OCku�=k�<3��EqȆY�Z��8�yQ�x��;�
'���_e�n�A)t%��D��Wpl���v���^ube��g$Y�Ӻ���awd)�z�}��[�nԓ�O���x��F=.�X�K��C�%N�Y�c��^I!g0�t⫝̸��5�
�x�\�w�
�u^�	^d��9>ȸu�u'�ӂ�͒D޸(n�v"6��c]�ց ��j>���Յ�e%%���Z�)�P�u�\���F��]"zC��sh�|�	�9b}D9��k]��v�<0qB�]��Ӌ����\��NVf�OK���{Hm9�� �c�v�^b�Ψ�����@h�Ɠ��}��s����0*������d�%����iX���v���%>LS��y�m�=������R��8�v�,H�����D�u�B�n����7j�}LpAN�G���H���=v(�,��
��N�:λ��'W�s:g�K��nr(po�4��:V��@rUѷ�+2��<����D�'%Za;V$�A�YbqAGu��vh͢:�m����I,��k[�ܽ��)�b�V0��ޕb��pX[=}�4�غ��ӳ}�e��Dɹ���3K�؅Ե�V
oj�v� �ݼ5��J��@�#b�OK��-�7��n����u�ʖ�&i��)�5�|9�lΩe;�ã�a�F�H�v��DϦ�'�.�7ʢ�宍Y��٘��A �քU��'V[�{��[��4ő�W��kp�5���֚рGw�.Ün���O���x�5���@ݵ���q��4����M]�`d���`Bo��	��ј�8�<�c�z��F�������i��]��m������n�Ҷ�g��k��r=��f�M�H�Yj����'6댫�9�7խ�(N���Y1[ݺ՝S>�-tA:��*s��x�	}��$��OI�µ�s7��iޫެ�B˛��v�f.�-����Jp��A71k+N����:R�ܚ�j��1#�4�uŜ�3~�u��]�Ø�4��/����wZc�(8�O���p�I�O�,��M���r����;��U�[ Qv���ປ���\Y���y�4�\���+��[��LsW[8ը֝�˰���fR��6�jS�O�:7��S���
�⼧���8%N<J�$RԖ����	EC7�k�%A%.ٗwd낺��S�2���d��3��-�H�����d��=-�Re�f#َ%��z,�-3�wq�Ĝ��!wp{�6�Ӳ�wC��X�H�p��ڝ�Y�-<�רX2լ���Vf�KF+9Fn+wn�6h@ö�P%�B�W�s�süZE��ϝ�w��KT�®)����s�p*S�t�pd��vC�8�v��4_g>���8s/8٬�%˔���q2yר�q��n�tۜ���X��w�WY{���qZ�n��mc����3:KW�i��:�y�^̌�ޤuѩ�뙔��3
w�*Y�ٓ3���	�ݮ�M])�|�;����D�;�I�6uY�K]�I��臖H����;��3n����۹(����䂺1�w�S��J��3#�f쫔�Yx��ੋ���b|n��L��.���>*����y�a'mI���fw_�f��ܸ̺uɾ�v0E}M�g
*IJ�]�T�}�1榏`�hd5�ML�K��X��ɽ*��l�g�L흕t��f���u�'+�u&�M;T)ӛ�\F�����9�f�3-�+���# ��O����c�w�.��ʈ�D���H-��O=�+A��}2�uKlm��th�d��f�*�Nx�l�*�yǻ{�h���0��e���P��^U�.���ɗa�8�^�Zn������e�7��.u����m��pK���NR^uN.^ή�fl\�f۵~�=,��^��~��r0U�\��fp�!3�J������K�D!,����R�'[8��5-+G+Vξ�:^���[f��S�0U�wGv��!)��d^|�v;�r{9[�LۮJX�sd�m+器��BU�X��D��Xƻ/�۬l���c��ț�gރ��rz������{��Xk�5ܒ�S��o뽘.�ӴᧈӔ��3����7�Y4gbڗ}Kh�ygL�I�!���:�͍������.��i��i�F� �y�0]�rk�˰C:Nu3�{����5�z;�XY;Z��òz@`u����`G�"Ӎ
�q�qU�(H4�����s�%�n��k�t=�I*b,�N���d<�����,�����P2�bp.�9����K���<�]�o����GVXÛι��!�LP�:;�Ը:�%n�w�9wc//�P�q}g��:NT6.G�Qeh�J�.Ń7�G���2nt��O����&D�oE��붲�|VַpwL��ԧS���Cז�ێg���<������7�����o�o�\LK��r��7�G;ë_	�����#:���i�f����N�w+"*=�}����fgdc����7D�ÎA@�۰KkP��u[��{C�JR)�e술$�xt�E�ŔkE�z�HNO�z*^"�5�2./��Hܫ�.�w�;|�}.}1��r��H��Â�n��rg�J 5��vu\�x�OjP�BwS,T�{�vJ��ݒ������/����jj��VcT�����c���fp���Y�*]a����y7(�܋*�&�0[�C�k~�����X��<Z���:u$�����������ozZ�	�+
ܦ�?� 䳲�c�f�ux/��ÆT c`�ι(m����v��䮡ą�u�'���y��S	y�hVX�J���T-b�g�i��ʎR�m��81�.1[��b�JB2J�Fp��#�F>�e�kg~�A 8!��Pv��K���_ue����>W ��9&ne��ʳB�k�{�_��m�z/��9LDx���Z,Y
�&�(�Ne�7�R���S������J�^�.�%��"�U��(��v��8��KA���$'�fS�\/���:�j�_���k87��xkS��}��<�E�,]<�ξ�#��'q�-do ��y���[8޾ŕђ���֪��S���dLa�*��]�橳��o��n��锯l�;;�m���,��+��t� 8��$�7���Uz���[.�tO{��[}��԰�\� A8vId��Nokn�O,���5�5-ȩY�8��W(�Q�w�f\�^��署�f�GWA��ձ]��Ǒ�$un����:N����Ko����P��-���rѕ�)"I���+8i�M�=j�1���k�u��KM��T�)�5XU���2�W��������:�q`#M1���;�e&s>WΒܠ#�.)NP��js2��'W�kj��u���zQym�E��x�^E|\c������w�y����[�S+r�Y�)&�핏#�ƣ�vtb�	(.�;���ḧ́D��')b�-nrnelΧKu@� �*��V+z��xuvց{MY�s����>��f��<��c��e"󮭽���7�+;R�a�	C�s�y����Ө�B��KW�a���8����&{]佹�x��ʹ�b4�*E=l�)�3���v�5ywׯ[���ɓ��d��uݖޕ+x["Ֆ�;�0��@6]��c!|k-�Z�4Cn���nTB�*�7n��og�e�j[ص:��J�쮠����B��'w�`��/��M�iƛӚ�b�"�ȄmBCvR����Pػ�#t�8�D�Ǘ���D�-��Kp�t�~\*
�u�[�J���'4���Tý=�V�x'�܅��9Z�1J�ܝ\�[|�h��Q�M��Ϋx^��N��΅�Ⴕ��9��0�%�ȨY���H���z��|Ci��.��l��]��S����31��^ �Ǵ4�q�-雈�S�C6�GK5�y9vY�ز��^�upz�f�t�$�(���L\�iv���y�����7��J(>؝z�g��o�vSC�Yݴ�.��IܝG���Y�.�Շf�kfG�sZ��R}e�i�zs�uԹ_��`��x��=Y��:l}��^O2��}�6[���j���5�����r�}n^D��`�k�v�ml�}�8��\�s*:\V�.���R��2�Mn�ج� �o)�������ּ���S/�^G"�\*@��T��ܧD9����H��N�:�����Eۨ,N%\�֛VM���pA���v�銘�X3q�ۼ�[��J�>O0;�ۢ�Y���d���-��o"����!��4d����}ҝ����l�\�S��nݗ��ɲf.��%H��Y�3�7�;��H���)��+� ���b�6*���Ȳ��+�],��i�1J�ux*���HX���{Z9�30!+�hg_6��Uº�(ʓ3}X���O�H:t
�W�\@��"Zޝp��b���[����
��m��N�o �b���+^�#��uԫ�����UNS��>��ÐE�z:�Ֆ���|k5����@�Z�	����\�Z[H s5���=�*�'���nD�p��I"�Y��0��9��	����'8�%u�S7�+�N�=��6	5�^Tko����!X��ju�-�s��h٪!N�R���K;�&�΃�n�q�Ei�D:_2�|T�:<���ys�j���z����^��Pc͙�GE-6.f�q�/%D�6q|fQ�Ru�T�]͎�1���L�IS\�O����g6���ۭ�'r�rp����&[/Q����өXN�>mmZB�2Ėh�t#k�Qs�Q���p�f6�ɜ���7�9�M�K��Y��-[��;8��R��t��e�֛�c�(o:���E������n�qt|/�u���U���d�'j��"�Ю+�x��8OZ�
�2�l�(�u���}����vW3;)��e�s��.��R
�s�ӫ���\���b=�h�rnVUãn�����k��t�iTՀm�l�O�U��*{��X��i|�6V
�s��2?��P��a}��F�sL����H�W`��v��&���ܭ"���K��;x���-���c���o;�綊�L�C,�λyA�����k^��Ԯ}O�\�j��T�S�8��bTM��p[�+mSڒɪ�|��8���2��V�H�5�K������!�N!X�B��psk/3PC�m�)пw��-�%��Y74"�ڸ9ζ�m=�����<\���'^2�ܟJ煋t&g>v�޻����t�o3�bT��'����hsk��;��v,�.9��\v���H��8Tֳ\jq��-��E�������t˝��R�$�)k����=�\����{� �tbT\wU�ZZ��e��-��w�:�f*����I��|o�r��Yw7G+��I�,�����9`t��[���_��{�����=�v���2�>.��Q��\��XBy}5���E{{�s{ϭ.��
ks�lΪ2fLӈ��,e��}J����.�
��额�p���##�ݥB��z�Tnl�)����(c���o*�ă���z����*nu۵��4q
����1�6�m^��K��/uc�O+ ��B��lǵ�t���`�6�A��i�qs/ ���D-U�� �n�M��z��9��e��D���A�Z��g�_a�k�2������a�F�=Z�:�����]B���CjЂ��ˉ��'v"�����:;Pn��tj���I������`̗�;�&�2����&z���[[K�ICW�w̼�e%R�g���->����`v+z��oF���yu�"�h�K�������E屮��	]Y�w�6��_R}� ���+kXn��:
���W`�c�S�l0%f�w��p�ɵ:a��:���v���	$�}���_up�+{_�sk����PWú��B���e���$���QF�X':����>��v	}Z�7��A|�N>�R���7\��૖�C��)�*�Q�vn���&�8��.�λ7:s��{�;F���,V�Nu���HI��ON�+V""�*�Z�bV�Ԯ�bm+KUB�%���}[u����|�����-�{����7�ߟ��}_W���;�7�@Wg�m�?-����LU��g`���e�?����nK��������:��m<��.�]�[�4>rpbL���(i]9Jάf˜&P�ᶉ����>�to���w���h��'Z�`^��U�&1����"pV��]����P<t6�Ɖ����������i��q)V��Q�A��ҕG�t�F���q�盎a����ֽv��U���4�.Qng���#Y�ȭ��bٜ���G.bolry�\u�h�������7w(9�E�(���Yv�K{/Sؗ1�t�rQ��?��]a��6']ܡ�hVF��c��
Üy,��!R�� D���Z ��,IFa@I�S渉V{-<��+�R�+#t����,�sr)��U.�����3m�xE��0��r�V7
� /�'O%v�n��Zo�C�u��]�"�ƶ%�M���W�M���nkN�t_咳��E�L��[[�* ^��ے�n���'oaE�t#�]R�SA[W��y�i������N9Ɵ�z)�2/�����a�ز�n���]
����pE� �\��W3w�ڇ.T���ܦ�ǝ4�t�k\m��:�+�<QT���6T�k.���b��e���$���U��Q��Wm�,N�wU�rvc
�PJ>�:���vc&Dbƴ�MYI�F�+q��dX�p3�������|�5�A�6�4�yq�(՚-�m� �'r��z�o�a�n�ݽ��R=���|Z.�����9��'=�cm�(>������v�j	���|�:oe��1��1,�?YsA�l���}g9f��b�.��V�o9듨���<ɮ�3�Vɇ�m��Y��\H&ެ+ns��(����/-�LC�3_��s��m�����2��G��r�C�j�L��X�q�g�Su|ke������\��e�;F���X-n<l�L��MշQ�nV�z�,�s�� �Sh�<5nu
OA�}�Z���hl�.�g[x4q����p���7��j��Z)l��#��]s��8�Y1��u�-��le1��.�4��K�.��R���/����/�c	������w��Ƌ{��udTz�۱N�`r�9G{��f�{F1I�Yo�%rs�巣9o
�t��"�>��M{u�(#�lQ"U�s*�:�E=䇢�mY}�)Mus@�1�<���hL�*R���]6��9w[t��A�kti��%����ܣw6�n�8���=p�qI�ǑJ^�{�.�.���⏱�L��ͬx�	�	˝�)d]�q����J=y &�C3�zt.����oVwe�������.�ۡ�n���=.����pנ�b�TQ7j'�g�A�++W����$�(�S�c��@EC�u��e٩���I|�R5\8���.���4Ⱦ*��Mq�([{-=�U�+���\{�|6��KӍ�)n23}��s�G�z���l�R�.�ZCl�fho���1�\%�����YR�9N��WR�ܷ���&��� �94�<�%�L�㲦�5�qR���!'*Wv�V��9*}�t�����F�f��*Q[n+"	d��c����;�X����� ��^��q4�o�k�;����$�7�J�I�w���%����ά�忙�q��Bvr]C�o9d�GoYkz�;��������������xY.͝�E�m�M���+K4���㲎Sg1G�u�L�j�}�S�n7��*nSQ�1��7�ǣn�X��6�^$��ܲ�T�LCp��ʾ)J.����o\e�dT�6�*��"�[[�v�.�2I�D��
���.��G
B�!ʹ�7]�ň��AiN2\�x_�N+���R���IF�v9���ͼl�r�ku���j�V!H�OS�ʦW\|� ������Wi��)�u	׼��f�Э��4k�r�|C��;ݓ�p�5
��S�/���E�g��N�[jO7n�l���5��s�1+J���zQdE��S����K�y�+������%e���̖)�(ו����,F��m��V2��Ko�TM�.�.��-�l����9n0M���]���7x[���RԕE��`=TEh�s:�f�
�c�@���]��*/BMy���*DMCpQ�
�%\�q������)ьܰ-�xd=n�@�J���O�++(o�`�Nnd�t�-���L�6J=���r�KoH�:[��9K���L�]]���n>�V���	B'�,�J\-��߄������o chJ�t�7�/��L��0��A�
JK��V���j�$`���żݎ�͉�-���L����9^�,jgf�5�`�P5��ǒ�A�W���=�e3���̭;�fq��[},�z2*r>��]�K��t�nqZ�S�K�!+fW ������o����t��Iss���n�/; �MC$��G��jYu�u��#=�����v*�������M�쭴1�\fس�[���.v��{2�ݷ,Y���M�_*��ÖC�YNi���:�Rm	α�5�tf2m��h<�7"C,;S�e@�1D7x���V�$�o ���-[A`]5��۵[�q�K�i�-��J �m�/Jfm�;j3z�RJã�`����ȫ�ެ.L�j�%�.��{V4�y�����4�f��Ҝe�;K�m�K��VScVm�f|�s�\�t�T�S3��G�_$Mf����6�L�����\��s�5�kN�ݳJ��X�پf�<�Ӛn���_^6Qh�eYBl�]I�:2,��R�7���yw{������4�i5�ĹD9��9Zt�W�)<V��ov�չn�c�ŕ��^&K�{*jĔ��g��.��O!ٚ�Lک����eVZ�}�Qg/A�W���&�K�aY�ݫ��72H�:U�Qy�d���sr�7���J�Nȴl;F�Yo\�]�޽1����q���3��;/�{9֕;(���+Tr���M�H�֢d�=�݃{hSɄe���7�SŽC�u�N��]sZ��̡o[������<�>Ǆ,Y��w76���djc9wR�Fa��d��\#�E��'� �"��Jd�'j�1�)�6QB�/l�.9�x�1AY\���s8N����5����Ot.�ʄ���W$4�͢}i�i���)�8�-�`�}V$�j�����p��R���sgkq��K�,}�V�hVη��+I.�$n^4�{< ����m\9��˕��mJ�c��/��M��js�oL׷2�,ns�A�4�n�b�}��@�<���wZ	f����l�q���5�b���2��11v��EW:B%<w���F�{�s����*��b���[kj�*t7jTc�ð�l}]@M�����W}���/WU)��R�e��gC��.�8ԧ�i�0#�F��k�ձ�fŎ���{mc�����7$Ӡ�j��]�>�v�����f�d��]��/ygL�K��J��%O�+U��[Y�#�-Hj�-;C�{8ku1Gi��#�ni��F�ʌ�dqz���C���d��st�bαO���"U��i�:^���5r�3ݔ��4��S��J�Q+α�&�k���M�2�L��o>{/�T5ԨY�u4�n�kR�:���.[g>���/��k�w�F�S����͞z��ǁ-;�.�����]8�7��4��C�7�t�:�;��f �%�b��ڃuWp�ԍ��k��x�QYLW[����29��S��!��ܹCZ`dP��}���P� 

�g��Ɋ9�.�s��c]>��^<��Ne�We*]sذt:���zL0ao�����:�վ�u�ok���4�a<�i mCɛڂ�8�T�U���[����>t�45f�úi7t[��+ꅌ�;C�Δ]� Ѹ�CGc��ŕ	CjX{fA��d��L��%˾h�Ҳ�e�y5��SV���McK�8�v��=��;m+28������J���%�jP&_L���b��(%��a�.7XG�:����S��u3{G�ghÈ������Ȍv��qviY�ñ|r�*�+ċ��ˈ[���4��剆ڝ����j�����*2�I1Ьz�r=rgj�if뿜t%vv���"�k� �+�l-�t��[\��*]ފ�<��ot^2�_`��lc�f�ώ��.N�֯�y����䋩�	�+�d�EՎ���A�H9�q|F�m�4Y�I��:�4n���ȍe�;B��m1��C`�Suj��\��,�����'>�=�gY	��<�<�޷��.�ˣ���SY��݅�$�2u�2v�
'W4�S1�i�*�ӽqlL�M�����m�Pu�0#�A���η)�m�UJ��s�/�H�FJX�6.����u��v�+�V�Ʌnn��\L�nvd���q�}�*Τ)��cKm�;w;�)��Z�8 �o+S���闪T�w)O2��<S����I����J&Q��}�%@����f��4�3�D8�y�_.Kjbۚ,:�.�>gfp�/γZ�B4-�gu��,������O.�B{]��w9	���������6��t:�l �`o;V�yݪ��U��WO���6���㦉\r��;�Z�[H^�!����If�'fw]򙔞��0[���Y�t�im��*�m�IV�g���+���N�]W{nl��T�v�4����X�
�뮻�Y��4���k4S�+e�+��c�(�eMvq���J�R�v1F�3 �:��[.&-�R��xZ��cG�ƭ΋����CB;V>�ҳx]sI�ʗu�q���
�r�M�����Vs@��ތ��]$�/M�um	9J�-�ɶ)�׵ft}���]��S�W��ax:�(gP[97z^�E`p+.J����;-��A���|�\�����v��)�� J<{�3y�K��N�%B��s�e�4�L��qntA�L+���[YǺ�GJ� ��#9�9�Bs�59���m�ot!�i� �yR+F���jG���Ğ�3��k�qSxtΗ���2�Ef���Q�\�n[0ø�������d�j�9�v��)2cb�F`{D��˾�ҳ��Q�꡷�	�]�!��c����d��,	�k�+����lj�)�� ��tn�<n��*��i��}v/�1֡,�y�^m�ns-7���(r��qFȂ��-�=�1.f
�IoI6���{�Y<Ŝר*��}����>�q�yP� sMJ�v�J<�n�38��P���%i<f�)��O�\��ݫ R�6��t�����^����M'�ӑf�rm��G��J�x�s�[{M�%-�w��w#�o�.ﶀI�a�Y)uu�(��0WAl]gl��L&.M���M��@b���I�jb5��bh���Nh�/��d;<���Ẑ�{�+1W.�y�a��M���7���ơ�SOlD���}H�t:iʗ���L�ӫ��ޛ�RM;��)�Lu:��ʄE0�V�㓸eɜ�\:�r��A@\����<�O�x6geu��clL��m�trX��3�I�5Lͦf���޺ͮ�+{�hUj��r�:|�[/n�f���]1�ʺ��L�,]��O��1V>�G5d2���O@Rͺv5Zy[T5�A՗��w|ә�V�_��W�O�krµ��x����E��o�Vv(�r\�f�"��@��1p;ih�6Md\��+�Ұ,:=u�>s�,]ct�w����Q�tJ�$It�kT��
���E��qq�kjӵ�	��+$�J:Kto��nɫ�V�]�����*�;��U; ����IN��GJU%�o_P}f���yu����6��VY�1rKY7Ȍ�4�ch�+:X�G�|6��˴z"i���{��̖����#�k63�\�5������㹂�s�� �jy�'���CY���7z�L�އYuf��+iY g���7�h����N1v��n����FmS�Y�t��D�795��p��[�hM%M���J�v�#wabuo/FК����,(���3��(�F�]�dS�/��[�-�s���
�ݾ�x:�a�ڇcv�3�+���1�'8�y.�d�&�=`Kn�Ϋ`�\��p�q���2U��;l\J���d�4ަ�#/�:2�a^Κt���˸cc*�f.�Ң�с��u]B��� ��:9^�HnT��w�n��:�i��v�κ�/��՛��%v�lӠ�J{G�]s=���]���
<���xeձgj\\f�o.u�^*&�z�c���h�Jه$�p`����WGn�0um1�@�ڸ�1�޷O�QP��k�u(W��6�;!i(TP*̨�0����v�6�X��]������]XiRO딓����)̊�u�`d	l�JG��)u������ NP���N��w���I���u/�l�W�v���J�u��Jⶔ�n�}��Y=��� �|-(���U����\�R��
R��s�M:��&�b��TA�=�εAV��ә��g�'�� ��S�w;]�1�E2x��]L�kk�O%˩u�l��N���;7mAK$:֌t湯�j���s�2��*/��f8�smd�# ��MEG�j���q&�������*ģ�u��`�F��[�.MQC++p�$�:BZL�1�����A��jo�Kk����8��k�58uEl��9ЍNwP�[{�̐ww���d����&��y��^Vp�'Gd
C��%w�kӃ0�h�GQv��Fˆq�DȞ�K�뼒��/�EW@f�!s�Hm��ձ��z��<�����+E}; ffK�)w;LK�\oXR�]��/�Q�n�nGY�ˣ�N�ȇLOI'v��W!��⭢�o2�t��p�\�����O-�ɭi�q$�Qpu�0�����j��ig4�!�S�:����]N2����ۙ��8jZ�N"�j����m�5��X;�q\V4�c�����y��o{��&�D���<s��=s"��<j,�&�x��)q�n.�ج�vp��U҈�{aL�캎�ς��/���+�{ҧ�$��\��.T��Lg9�i��&Ю}�#F��Y�]��4�69�g�䩕yZ��j7I"�H�/'�����Ǫ宦��f��ӟ8UvwnK�!v��ėҲP\��G%�s1�呌��I�>��jQ�i�D{<��٘��-nq�u�ҰS��������5.��u1�>�����VL�v�F�������zn�5+&�ct�����;)��z<]��|�e�5�G���"$��H�:4xv�z-�J�󫤃޻�6�댼u��	�ĵ���}�������\-̓�VB_R����u�H�5�LJ���)��wN���Ŏ`s��*U�AQ���Y�.œ-��#����9�<�;�5I*\����9�7�u����7۫h��6��p	�/���7�'B~��n����_.8���<q�s��k���L:dt���ure@]}з]I8���9�3�s���+�bm�G'U�wv����3�w{�����6�}�ou���0A�	m�:�z8W\�\�;؇!Y�\%H��t�Ve.y��s�p}�|�ډ5�8 1�K�\�
��g��6�p�-�J����������szJ��*7��h�訾q�n=�4�h  �x�8ejj+R��$�ED*EXrD�.hg�Ux����'!�Z)f*"�b��k��T�E@�B�έ5!0*�����#UR
�F'M�y�' �E�+��FV&Q%�T��e�U��*n�A'����UEf*`�e�H�F�qRx���*B�+ �Im4Y�I����
�U�)Q�+� ��Z�Jl��x���p�Vs��S��
s
�$�-P�G�v^�ET(���DQQ:
�G�.dR,�B�W�D,�#J-4��y]�%F�r��/WD�)3$����ʲ+A�B97,).(�Q�Uʉ��$\�	*�QgH��ATEErI-�䅩��jf�QW*(*(����%�<���&�q3"��(�H��A�nd\�yFD^BQ��*���� ¨J��a����U���t�e�9�a����O�I�랱���jDҜ�k/�1^��ӆ�c�î���r�9Wܘw9.�Oj���|��]��F|�p�u�PR��ܬrYXa6�k8l�mņ-ʂ�Q�J��<ÚeŘ	L��M|rl+�[�B��>f�d6+�
�,I���:�;Ѿq�Kl�n���.���޻���o�5�P#���_K^�ʵ̖s�n �(bȳ���2\F����L$�tw؝0�,{ʘ,��>&�ѯ_����������^�r9��78Nf�X����*u��df�˯Y����"���9}��k���6�{�T�T����7Pb003��|��@�uu�u�i�Ok�Q\olQ�ct��'7�\��7��<�����ഷ�5�P1&;�ss[n��M�ˍ�ی���
2�"
j�dG>YRk.�e�xԔ�����w:�X9�kp���'[�j�5�DX�5q��ĵLvv���O�0c��C��]4��x8f���y���z���JK,_�1��\!ngz�� pD�*��>Y)�ZF��'\0�v)p�0j��<L��v��ql��hB��;��}��_[�������v��{(-e�g^q�h�3��G�S")]gӐ^S�g6���'����_m)9��@V�3r�7v�j�����tb��'O'ay�196w��{뙌z~<x1a%��-��[sB�f負˳`��u������2'��Z����S}lW���>��)gKF
I
q�f��\U�gl��2�8u�����H&
U��Ƈv&�ݷ !I5hd9�f.��bQ�k ���Q_�-ɠ~��ғ���*�@{M�T���og�'��
Ҩd�bzn�%z�Jđk�_k�]��q�c���v�S6�cA�~9?L�b��w���L�%vY.=�knmΟ�M-In����j��)�&�t8s�`�����8���4XHퟞ�T�N�r�̝:Ԗ/�e�ˮN�؋�s�%2�NjwCn��EDq�:(�`9)eh��I�M饾���H`�����ï�hXB�z�ddjtW��:�D�o2��0��Y�����î�[�y%���Z��v�r]pU����(�7�>s��hG��Uu���߽���O/�gHКa2g�V�<~ՇRy��c������u	�Z��AV��V'}�F>��DŹ�Vz�i:�_uv���Y7�z6�+�`�����(7w}�Ք����*���a�M���4[�����x�R�ge��FAP9c�Ͳ�t�����8���Jk��0��N0%bvg	֫v_s��6<�]�+�n��S/k��7����v(/�Ѩ:/�K���Ժ��Ш�����@��ڝ�M�{�2��m���|�����+b�|²��jus}z�XD4��/����T��x���#�Vv��}���3LX�:�Tt�E3^��o��^T�h�5�8^��X�t_��17�ֲ���N�Aꤝ��v���ɡ
�鏞�,Z��v�W�9^q���������]Ϻ�2H�����$��1�2�*�$�<�XC*��-�-���gn��w���y�����[���g%	��(������0R�+�.R*�~ѱOn*�+��)�оq9],wk/�;�>�W�f��l�(M|�Qsp� !#��@�S:��0���Y���o���aq�:!3�9��nvG]:�$��J� ������������^:�^M-��\�aTr�h㙎�Ù�J�k@��B�y�!�H�����<mV���������H7`l�v���ԘI:,�s1��ȯ��d
�yN�o�~%����%��U���	r����8�����_Y�X���6�8k�Rx�O���W&@QSW#6�5�����kl<��t(θb�̸>�)v��z��:q�FVD!�ؖ[}V7֍v,��pv�]�l����x�����A�7�?w�������5f��w��܋	��[, �)�*��/>d���<�7C��I��5RA�?n��E{m!�������\blx��=N{Y�q��C3�^|�b�)�HTȇ�����n�.��zdF�c��>��1{���t���c$�}^ݠ!���S��٢��#�6cG����ڛ�¤_g��_��死2�ַ7b�L��f%p�m>p���^U�q��.>Y'��?"չ��e����-�*�%���F���eKk��y�3"%W"�*X�ۄ�xž���*�Hm���u�CV��r����U�࿜LQ�q�11��j�>��2���&Fq�v}����釬���5��4p�C����@R���kua>e��b�6f0^,xHP�`drWK�Eì�	�Y���
HorjH� 9։�f=���L�\�M]�9�ݢ��!�l�mQM��Bey���Ҭ��@	ɣ @���xwL��< ��=�k7�������kX��?�f6o��}+�8�`�Z�t��j�s7,Wj~�{F!�5���e��I*�ue�n��@�BPi,P�Bky��u����������� 㺹_>��S�_L���[/�"�������F���^��3��^>�#��t��LF���*��d%P/Sz�\��C^#�E�s�H�r4!�Zg�V����c͗�!��_<u��ِT�GT#������o�H�9MAX+�hK0�����:>T���rՖs�F2i�@t�'�c�Ū���e��X����H���(M$X�(s4��Dv������M��^C2��u�㗰�4OZ��U���STu�o�P�l�tz-e
�>�\+w��l�v�Vn(zJ�#J�s4s�	q��0�%��46ˋ0&�d�>;fø�m�9�Y�X+<j4���6/���B�n]��G� +/�v#�X�7Pa��,�����TK����-�6+^^�R�[�;s!"r��؆�^�J��]S�tm��07��!�{�'E
��$.sln'�mZ�:�S�Z~(�7��H֮s3c�:�rM��u�4�H�/g�ۋ�[�����s3�]�c뇇��xn����g8ߗ4�D��g���x�{L�TeE)���
���7��:�2�ϨJAz)1�#m:�b�!SC�T�T�ڷ�r*��b.S�G�P�EW����W,�:UE�� �ʑ��:u��$V�;���d�U�!�z�'d�A-��U��\%C�-7u>ǖԽ�N����!AN�펕���8im�4,��~�$��>
O��C_��qT�缜&�jhb�%�خ&��Z�m�xG5R��/�+���WP�D��X�>�+�oļ9Z�ڞג��tg�3�O�#��N�3�c{�U��R��xc��=u��W�s�exj~@g�w���>v�..	c�[g��ӑD1�ڸal��EBRA�5N��:ec6���`�[ً�����%_�(1���ijN�3�װ�C�4�B�:�3co7jv�/�u3�e�? [魀P���Z(\B�������n�������Z����q9���ko��с��"T$R�&��cC�j;n B�j��s��¹��ά�fGl-�5��4a.u�\KǑ7dHB�� ��@4��,垅����®�n�˛�!L���_J̚1d��T�y�h`��c ���7��S�Ǝ��l�Y�K�[�%+����>��\f诫�]PE%)�&�7@s�8�xE�h:�ߍ�
t4X��]pzym�W,x��Zz��ۭ�(cV�I��da�#��9��#�wK�|��v:4�<�VˣF�����t��s����]kB�����Z��N���敷�[��y �x�ۙM�XsT��Aʫ�|����K9�=S���)�n��E`�4k{;�~-��2V�꺅��ܘ���ȚN\	ۈj�m�Tp�5� ����Q��eJYcg[&bSXpTE)�b����B���>���[�@�qBv�eºj����z'-�>񄻡��Ctב�3��s%67.��(�7	S�.{�)k��V�^=�޻�a��{�4$�L���<��Kh���&e\ _M�~�e��]��M��ڙ�������NŽ
�{��?����?��`��6FK*i�*FnA<l6Pv���W�E�q �u*�Y�_1Ⱦ1�'p�Ԛ:7��VOuA,ζ�Drڞ�o�jPtì�4QɄ:�:�]0L�r�YM_܌_NP�f뤃���"�l땞O�z��(T�N�$zyN�b�>�[���0چ���g��F�[׭cur��z�
�ꅒz�` d>ja
�&g�<�K4H�U,`����b���Yٽ��AU���8�<��(�N���C����r��h*=���z[huR������Of;��Rz{��:`������^��L�����}�햘��K��V�%��(YhY�Z�"�zr����YpFN���6ױ��i��o�5)�P�ɴ�\�kd��V�17��]r���Ǵ����E�5zo�zֳ��%�t�_f>`�s��lۼ
u�Ẳ�w"2W�Q���M�7�  �����@����aqg�!tv��mG_gP��KK�a��=<�'.-����6\Ђ�SJ�T��pHG3�9`o��5٪.m���ڕM#C`-/�:�.��9��\C��'��^���y���tC�$GF�J�}n�{���Q���L`�A��+��ޢ�\jLRI�g�F���2*�d�Y������Y)�H�+������N�k����,W����N�!L�X�k?����w!4�j���B�B�OF�}�'p�Y�9�QB��,;k�o��Eu4jL�����܍w�]h�,�fᩡк�=���7Gu�[��6�`���<v�.����;2�V�=ݶfh�L�� +�j\-��4_����
|���������L�_���n���.��^�sNϾ�U'��"Ms dIcY�n��ռl1�cE���.em�.�}ʙ.���f>Bw�ꤼ�z�����������9�C"Ur*Ky����Ӏ�S��o���-ØܦT˯aƶox�l�LT�3GG�>ze�� �
v�en���j�3�n�1.�|˥]�ο���$�4qwf���.O�H�:uk��X��YXnV/�9JW.�w�L��F��J���,�V��E��h��]�C3H��0�d��tY��Va���&7�ud�����.(VR�e�11�[΀�-�e��S<�����-�����+�c���YS����ǹ(צ��EҐ!Rڠ������a�.�KZ�ONW��OH�oj|��G�����w���@)b܆ڒ7Hu����xJ����h�VA�Y��P��+���7Y��O+z}�Y=|��F ��x}0H������ڃ�Nc�n���X �V�@���k�gވ����؆����Y�!@V��U�`���WM��1������ztE�#��9��;l�@9���cw�D��;�d2Q��u9Y}��u#L�wM��2�C�#�Gʒv��,��������rN����K�
��4��zL�.����(M*�X�7g�����s�y��uľ۩��	�y�v�yԬ��"0史 ��&��2��QQ���ц2k*��t�`IjOD��O���9�Z, EBr���)��\Y�?5-����c�R�0�7�(u�7Ҷxn���o�i����T���;�j�(�*ڴ��)ۨϞ�n���}��Rd���mL�D�]����ש���Ӧ�����ז���J�5�O6�ۻ�i���s��JZ���˭�5�o�e\���͂���F@.����B�t�U�%�T[�e���h��b�s���N�ro�(I���]�����Qk���"��R�->bfĸOY�y�Ik�LZ)��%���Պ��{�<ι�'��ы��K&0\���{�5�g,�7Ơ�f�����	��߀��Z�`��kN���}47�^��m�X"�eY6��;{3��C�����a�X", :;�"�y%�c<�7����9�������Y:=�[t�a�y���D�R�ࡻ��5�?�b WAQ]���}���}�-ɧn�����7*{o��&U�I���YQ�D>9!@�M��oGte*鼳��Ko��1�H���a�u	�R�1ثo��s�j�	1��W���7.,���mj˙�x����M�8H3�c��CRYzr�c[U"m�����RA�����b�<r]�p��/��]4������_)A��Z�#�ԝ*�q�*!��!�������d5}�;
-A7E@�� �=��)�z�}/���܆븑�}��̀Q��Z,/4�r)�1���(.]ێN�jU����� �yK�ʝ�^�T]-���|�퇈a��͵V��*Lfuw_r,�K�Kw-�TՊ^)Fn�O�km�Į��88�WJv��s�W[\F-�>ʐ�!��oQ�w.=����G�N}��yD��6бr�[�"��N������`�vc΁Wt\Wu�S�\���{�p�KXVP�Ớ�z,�7�)��G(��ֵ�uȻ�����[w���rq�*.���F��)(�n���t�/� ��6��ᣌqn�hc/WۉTH�}}��3Y}�2g8���ܩ�<4@��1�V��@S����$4���{l\r�������moq��y��R�SAVѹF��j�bV�t�;m7K)�=-��+cǄ�7u���b�lI�`��w�gL,�4��ٙS3�Y�ḝ�]o�>��w%J\=#�9g3��v��3�a{�k��2�KK���g{/����a�)ɪ��ӛ��haR��e��F�u�ϫ�E���7~uE�H����T/��遫�cO������p�۫�x�p�p���1��Bޘ5I�0���D���4Q���u!W��8��:3�
�������6&)Ps�9�{9��`R��J�Z2��ZU��[��&��tc0��BW���[A�u	X�k�k��}FRGk�jZ��eY[5����0�'F.'��+����]���o�d%wC�<p"���:₩v�ڜ>��"�X��䬧�,(�w�5���a���l�M�]R�Z���7�{P��ː��k�d����{��������m-�2�h�|*�0�-�`�=�v<���8�a&˱�#n�`��歡8�7yɛ���.p�0Z���f<w�l릱X�F�|��J��f=���1�P�nSR�'H�Y���z��؝0D�skl�b�C�n�ɧjK�����N� �8�_v�G��:���n���9W�1���h� �e�4�r.��A���.���r�T�V�o��ө�Cmؓ;mgF 8sj��Q���
%`u��Wv�=�Ք�>�ۥ��:�I|x.�P��]k^h�`�0�*�[�V6�@U��}zf.��ɴ�s:G��K��sh��
�)ݦom�B=]aތ�^���Ծ<�Y���Z��,�:k:���_ډ��v���W{QK�|fn�A��\�S�V���=�w^Q5���<��H����1t������f��bE�T���U*�V��Y��qN����gT����x6�g�ɮ��g���7�֪�=�"��{�C�?*�˜�S�^`�:���|�u��=X��ì��U��39�J�동�ɒ�i<�h���ج}�޼��I�^u� ٍ�OH����irN�X�A�J�M��5�:Y���}z�� ������:H�v,��Zd$�
��f��!$ť�N*�ĭ+᎐|�����j8���"�������\mũ���:�F� U
$����Ȏ֥PGJ�P���$D�r�UjE¢��DT �a��8]2*�D��s�\(��vRI�A^��
�`P�(�2jкd���jfy�p��V�l��<��Er͇T�Q�Ӛ��H���g
���Α����ʹ9	\�Ε���\IeȎr��JҾq�(��T�G���&�RdDO!��)Օr�6\�kU��N�I�E�E���/�B�˕E2���$��6&�,9ȵ�ip�(�:Dʢ(�B�+;U�)X�mg
�TT���U�N_U�
�a�ӕ_)r(��D ��>''AG"L�iPT�"Ǒ�T��$�TJ*(��.U��TJ"��VE�H�( ��l��*弹x�dEr�eEw���I�iv��C_I(U� r��͛�VFջ�n�ݒ�A]��/�C�l���FNx�eM;�ޮ�:��a[y����]´gFK���6�}z��Gm���o��x��w�ޮǧ~�&O�lr(I�M�
�];�����	'o�O�>[z���~tnT�v����<L?#��׿��N�ē����|���"�Az� �F\�x������;~�*o��vS!?�ܝ�|��яN�v�w�?���]�yؼ��� z��d�=�ϭ�����\zOi�'&�=A����r&�B�O� >���=� eR�fO�s���/�"#�a����׆_i������<w�k��7��w�������)�P�w�ϼ�����C�|���~���|L?�nv����z:?�x�Ǉ_�=$xG��D<�V+�|�-���kܫю�r�����,�;����瘓�aW����zM�N[����o�rs�?�>��SӉĞ߯�����$'z��e}X$Ӽ����?_oN���ؓ��DG�F����}8.�7������O�N�v���N���w+��y��ߨ^���m㾦�yǯ��o��L.���ϼzq��'&�~��͔P���;�Ͻ��m�N��O�����N���~�c��B��J���=��z�?�/�~*N��
{C���q�Q���@����^w㴞&���;}NT=��97�'�����ׅ�������}��0�������y$�>�x��І2�/���_^�<��?4;y�������~��O|NC�i�S�r~���raW8�����ra������=�r��;���~���>$����<p)�!'��y����N��x�������ٱ��+�G�`�B"=�71N��+�{�����?�zW�_~��O��C���o����C��!�G&|C����\'�®�y�x��	7���7�99�����N'}�W��~�ˉ���*��r6[}b"4A}����z_�	4�n��C�k����<��������B~}���w�{v�~�{'��oN�v��o�sɿ�.ps�&�y�ۣ�'���n�=G���ӿ��?��@֟eSv�s�}ٝ�>`� ��O�9���`�ݲ����߆�$��=�����m��>}�&O�׸��x=�ɇ�?����������|OI������~�p����ӕ'i7�'�����ի������d�G�aƂ�v�+i��,iM�0�\�ev��9S�4�N6w't���C�g]�̠#�-��|-L���V�-���[@=�1�%5kb���eZ8vҴ����Z�k5u��g�9m4��!�H�Νi�t�y���@����w�Vǃc�=��{�����Q��ϴ�0�'�n���N��~��8>2o����zL5����]'��}N~��s�'���篼�0��ߟ<쿮=��_>�� �"�x}�G�g��:�ɱ�h�ޟG�>��w�|�?{L�@?P�ts�����睃�o��o����x�����6��z�?{|M�7�&>;~'�Ϝ{v���{Qa��v�5y�1�X��)����$��Hz����7!���=n���8�yw_n܁�$��&����z7��x��׻���Ϟ��v�<K���o����;��w�o��ߎ�˯T�<�����e3~�B>��	��}>���1;�~�������S�0����?Sӎw��߅���������l�O[���ސ$�������|����&;_�߯�����a�z��)ހ�1W�'3<|�V}��>���}���o���ݾ<�����= rO����c�r��۾�='|�N��~����O?��Ν��~$�X�!�>A�0ѽ���'�o��Ͽ߽>��f^�1��=�L�S�#��#�� ��~����0��|����q�v��|���e����������t~|��]�9'{O>���bM���<O���=;x�����ߝmΝ�q�����������@���N^��!�x}D}U���[�'!����B�s���܇����$���z�>{�~;돉�߾w���&����|�<���N~'���z@�IĞ��{zO�� x�}��7�8'y���\�麪��{q`���}�#D����G��ӿ�G�x�v���;O���^�]��~�ro���oX�����щ�~n���q��'&���>��w��?w�8� (���_��zL?��z�����8��K��ڇr��1�#�D{��w�}�m�l~��O���V��߈ra����oJ��i���r}v�yޓ��(]�߾��~&�P���Ϟo�FQ������_}$��"�}��/%��9�~���w���C�߮�m>ߥ��L.�~��z���A�7;�s�O��_��aw������7�raO[����������$��?\~��w�_���P�� ���G���fIw����έw/!G!��.]aav�Q�u�<��	��(����D�T8�<�5����CsLz��e�s�a��v�0D^e��.���N�b�Ǝ�Ն���[�wJ^e�w��t�P�u�N�囀K�k�6x����UYj����<ݛ�m��
o����N�^���;Ӵ�x�>?�>���W}��<q�\~�Aɾ�'!�Ǣ��1;�����'���w����9��J>�G�"��l���"�v�2�|���c��o������n߈�q�y����;rϟx�	4�l�����>��^�����w봛�����v�N�q�9�]m��_���뽼����
�A1�w� �5w>���ۭ�{�s�|\|w�����~��Nq��NO~�9]�P�=~�����a�m���㽿Sr��.��}��q�}���O�©�?����{C�?/�_������k�|UT�X�>��>y��η}��!�������H�?�>�?S�p)�]������w�b|O��[}}��_���]�����^{I0������o`��G�8N��r|w���o�&~��~|���?�!#��ޝa�z�VD���u�C�#�%Ǵ9�kg�	2�O��� {Iߎ���܁�'��]��N��rN���_�;Ӵ�S{K�矉�Ӵ����{���]������s�����z��7�j��m�����w�t���Ʌ=|���w�8��������BM������Ǐ�oHw��<q�}}�s��V��!&�巠��Ǥސ����~���6����|G�N����a�w���1�k����v��ޝ��?��m��|�+�M���?w�]��={�N���ݏǜs�';z�nw�����x�U�E8��{C���G;�|~&��^q�����?}0��h�{D�aY�t��k���i�aT�|��ͽ|���&���Ώ�ܮ�q�}���$�]��߼{v��'ۿO��?S�\
o���������,���N�m���' N��P~j�BD} zY4�����eǁ'�^�s�H�,&b$G�뚨���8}#^�xo���]�~w�<�'�ߩ��Ϝx���~8��~���:	2�OG�߾m���N�w������;r�߷;���~���� ��BY���)}~�Q�u[[�~��l�t��G�>#"<L ��� �M�]���{q+��7��NB�o�>�1}��_�~��=�Lh��:�ۯ7����X��:�eoS�ʕ�n�z����۱5��2�V��7gw5�_M���!�z9͕'�����o��H��ݎ��<��U��\�����q ��j��Fvl�:�n��u���.���#{���Yq���zw��&�@*�Λ���"��V5����� m@)lп�L1�����I�d9j�9�#!��}�/�9���X��5k���SEtĩ)�@�� kh0y�i���\<�l�8p�?2��:�I��KN �̫�F�Y8���E�?���n�=���E��3^�2�s���|;Su6D�A��K��5�$���A�9�`iy�SCl��b���s܉2)��*s������)\��_9U4j���yS���W�&�
 V��c.��bW���	����A�96e秄_/Rw�r��d�Ǽe=���za�N'Y_k�bV}:6�f,1ݫ\|�y�l_[�b���4�F���X:�q�8M�gR�/Z�`��kN���Eaȶ��wA�)����ܘk�C�%�4��Z�i�v�¸��Bb�lO4��b'��L}[p��X�<Bf*�����C[\/�kn��8J�~���
��j���<`/"��'o�5��@=��S[n��p�`���3_mԺ��&�X�>�]Z]�1�ܢ|��'�GۨD�wc�ǥ�I�2���{m�K�.��"���{N��G���VJ���G�y�� jo�b�EU�+k�����Vi�D܊�y�)��\�3Pb�Ctt`�ɴ��g;M%S�j�\P�7�i�6�9�N�=#bZ�N���*�����e��W���Ji�*��9S&�!����f.%�bg=�.���5l�I��K�˨ǭ[gͮ���.����t��P����i���,�9D1�ڸb��2�4��� �Mc�ȕ���D��#Np�1u3��U񯔠���⡩8m�\�ʵ��+{��[�k]�6&���@��
�:��yT
U3�E�R��g�C{H�]:��c����{u���%��'�Ѥ~�n`3_" 5_�Bt�cٔs���r��ê�t������8�5;I�b0Y;�n�^�e A3�h�� �8���C�������-m����X^�W�5��^C5��/�c ���6����������tsWc��t���+z���\���Y���K�<�td>��%�t<�
���sA�N���Ô�-%W�u��:��R>�Aʕ��u���9�u	rwrb��������j�l��L�t�[�.��I�Ie�4VnPU
�,O��������u�΀"������{w���8�=uGe��qm��)�Yb��=,T���Q��8��`ֽ���^P;��2�.ۇcwbW�r|��s��
�԰!hܛWԦM�$̮f���m�2���֌�n���r�)�v�=�H�s+$�׻�E����.��wf���2���9���{(I9/_]�0f���ޑ�:<L��`�k����C��ƫ�9���vdѹ�n����
)�픺�`�2}�U0�j03(��%����T[���6��X&�������3D�s^A�*�����-���^�PJ�;vk+���r�.�Uѳ�!�me'&]�%
����Fi�����X~�u̳�S��A�̈́�z���xK5��A�^�6��q�<e��	`�ilUS���	c9�u���3�����)����U^^��ݵ9S�������A��#�P�IG���唲hB������t�3�*�u���+b����A��Y��kQ��M�*�J���>���U��%�}t���^z��K6��Ui��CB�0Ғ�ۘ�p��۸yr�7��9I��)˔�˪�G�^ʝ^kȊ|�2�on�\���z냥9O�������#+��4�Qsh�>`��[�n��M��3�ޏ�=F���\j�_��I��膎}v����	%
꒺jM����jR��[;:��S�4%��nE��ή�6�s�n֏�59����R����lI�X�0�N>wp7�T3|���� �V��,�r�l����A`Y��	�W��=���cd���d5��jre�FWa�01���iζ�|O;���u�<�3�}_Us@�F���~�TI|P�q���*���,��3���ցP�[2!I�ɉܾBj�tP�d�sښ�=��(;�xׂT8+Z��V)kƢ`i�ޣ�n�f�w"��������q4�ca�
�yJ�J	}��8�].˨.^��ƸI���'F�B��/W�/��L�<��!%�`�<������1��].��?5�!vxW�������v��]��/ܕ铡ƾ�bt���ANͧ4!�Q��p)r��LfKmM�`t����t�{�Ԟ��wY�{�3��<~�	�' C
�1]���T7�e��p�A>��lݞ�	�c��^�w��q��>n	�WLD�>�x�k�"K�g���=�>����X���|9��[/ԖcW�t������ꎮ�A�OƇ�u�=��+\�PA�����p�7ջ=Js��z�-�P�%�^@��)�1Mre�Lze�j�>ۻ���}=�{f�)QN� �"���kn���b���+���kc�8�_�Ov>EQ
K%�eR6��u.z���y<�G�]�֡� ߴf!��6%CI�)e� ��7q�f�nڻ5$�ˡ���SVx��Q��+C��ڷu���Y� �d�ljs_uZ����;v�4������x�!X@�+.�on�;�"k71���´�����_}�9��{��֦�����p��}�N�|kf�>�Pi: ��0��m��7Ik�ȴ9�&C��7�i%j�w/�~�R��(8l�����S�����L�E׶ ȍw���qΏ_�%٭{w����A�G3�Wr��2�a�Ja��>}$GS�r2�Z+!��DSv���D]3�p�u3#D���&xE���{hy��c �zr!����Q;�����"D�d�M]�Y�zd�p��Q|������^t���?��|�rՖb��m��ղ��B��
�]��'���9��i���$Gu�	�T��"�a�"����G>��&�QG5�WL�6~�Sħ��DQ�LBt��U�F�CЉj�tzͳ^��,J]Ϻƨ�3��s]0C���c"9*�7��健�23`��Z�d��~|j͏%�Yp���{$=��7:Y�;e���,���zf��F� +]Wy��Y�&�ׅh�(j��\g-��^�r����%��}���#�&���G�5C��W3�ꘕ��h���Y�%� �������a��ڏ{l���kOZ+nq��xU�Na[�ۦ��ÎI����*8��p�w�2^_i��dK��)��W�j�B�-D��p#�>嵂!J#t�u��%c�My�
�R�M��<���#��1D�{����9Yr1���ƃ���1�a������~�S���R��k!��uX>��k'w(E�h�mn��s<����z�b0�H�/�%�Up��xJ�ڸW2�b�P��Z��ګ̔��<�ee�5i����"��%>v�Κ�E��x�S����>
�C�;�=r��K9���-��?��~ԫ���,G(u\0nwezo��][T >�lB�+Di����-ޓZ��
;����mR:d��D0�۸L��-S��o��9&:�JW�� �+T�!\f�'v�����(s6�g��e�Yx_�D1��jዅ3��=w.�s����S����DA
��P��w*�iT�|��JPc�Z�#�ԝ*+�FgƷ�jccck[���n��8�:���mA�0�k�꞉�P<)}3�C\�_�l���ғ^� ��a2�D�o���a8n�������ti����|���G�@��'>&4;�F�̷D7�z�_H��֥�`4���s�����m� ���"n�W�`� 59�5�Jca�Ap�.�ݣ��yxE	����=�Y�̨Cy#O.����W�9��7�n���r�9�=5�.������jv,�mlP��]J玙7	�%NT��VT;��霬�`=�;_V[7��A+����i�&oV��x9:�3�2��/}��}�w�Mnbj������{4T4�-��S�kC!D'w�n���5V��S�8ӎ����l�s1�m�ct�+�n����T�_BR�2o�M������;Qt��$+��b���w���z�����Oa��:�W+N�]B�N�L_���Je��Xa�ֵ��sk�	��K8N�&��5UPj��j�5�`\g�A����z�g�}!��Ec�g����z�ԀC��a�\P��.Q��΁��P9��L>52Pcc��G��ũ�P��=F�GA�T��3"��?5wR-��;��Y�>���Z�w��\}^SM<�M�^�U��� ���cUC�(1�W�
�Ń�����?��`�.�V1�QW�9��Gf.c�źuH��b��� '��u̳�N�a_���N�
z�Q�c�{�"M{[;��ߺ�,׾�t[�%�"}m?  u��^�g:�0L�7)�����B=��̧�շ���m8�v:�}UڸR�>�� �|&�2!
���uR�N}&�+鏭�t�?���TG�Pz�`�� ��*�όP�e�n��\h;�$�fW*{�j����7�11�u;�M���97E��r�i5� �i4����Me�R�OM�����ݭ��v��kDK[c~o/��v}6Q���P�P�[��C-��g�fܮF������u+G\k�nLY���Z�ᶤd�Y.��R@wz�J̴�[���:_V�7rf]�T�jV��W{\2��̅0�rP������m\qM\��M�ϰHz}�z�f��X�t��|��ãWn��I��E�ym��*�SO�\�//��,�uw=���ZѹX癪�rFLU�&�9��ʶ+h�"�F�
9͠���U�sc;]�"c$�¨� &a_�o�u���˜#V]�t��<���=��\���wl>���+L1�n���O#�8���B�J^ͭ
�3���wnuc5��]P��>�<���nS�ؓ��S��v��ZbZ:=u�J�Z��˅��˛��CM�|��2�sq>΁�wb"�n����v��I~���ۗ�[ܰEd�˨&qM6��\{�.�&>�dU���q�P�L
WE�f�@���o������̤��Ad
ix/���ގ�M*��X��.�v�W;_6�dOb��s����\Ķ�X�v�wr��}Ol�ή{zE<�����B�]�P�TfƖ�ِqԎМ�zaI���uև$\S�f��/P�V�b�	�+i�Я���/P*�j��9%Z�ft�|�r�u%��tC;��˖�d<��H��u6�3�w4�I5X�����Fnl�K�f�x0��m��V����Mީs(����k�K�R�Ǒ-A�cAv��-�م]N�xc���)�V��eDfG�Tۮm�zI������#�/��{��1ʉ�-��s[ �.Ѝ�L��L�)���^Tt_n	ϫt���],,{-�׸�C*�C����-�l��+](��w�m�����#��Du��^�L����7`�/�MV��=�gI�5��23afsa���M��ǃ������-�����yJ���&���Md���%��U'L�,<���c�N��U6�mERħ*ҙ�y��g y�gIJNq��2����U���ֺ� �sfN�ټ/k�!M��|��b�m�۰����4f�Ι��(ҹJ�S�� A�W:0:糺+<K�}J�.�;��ݸ�e7�yR:�j����(�f퀝wn)kbZ��%��$�����y:k�Ӱ������ �Ư��yM��"��,���YM�����%uc�L�Ff�r�K���i:������[���l0�?J�t�e�|��bveI}?�ew�5��Y���;x2�L�u`���a�Y�����q�����!Ҩ�r�rS��t���R�zE�TeF�땬�ͳ3��ν�۳ͧv{[����ٵ�INp�VЯi���xr�΂�!��C]�p��u$u���!|h�@��]�g��޽���Ju,�TAb�*\
�!"�9'YjQOI&:��P\.9�UF�IFja�0�¢��3+�G0��v�E2"���+P�*֙�
����9ˤ&a��	JUTʎF�\�قt��M�*���T]P�]Yc�Ey�!5XQEZ��젃��G���h\�UUAJ	
��.�.Tr���B�5�,ԸPGq:��J��nH�S""dTTvDd�eL��D\>3�Y�2�DU2�"���(�9Th���4#�(�O,wXDQS$���i�+"��.D�$�9єQA\�J�SH��
�9ʧ�'��㲢��J�ʮ+O��*������z��ED|VZ���(y@���Su��W��*UD�O(DW8NFRUp�+#�EE鲈(��+�N�K*9UQT�QEQr8�"��w守r9Q\��ªV��=���;��ט�hm�r��)�y�Af�/���=���u�:��oo\[
�_SW!%oS�l�:�)���}_W�UOY�#���4	�%��y[��+��	< ���Ү�KF�|����#{|'2�S�Xh!�#�Y�sn��ϸ�l}�����P\�T�":bEbn<����}�^˧u]At�)��n��m��E�Bj�.o�@�h�tӊ�3��E�<o2�Ó�&�����t��s:!��9��o�ݑ�N�A�����p��ꨝ��+�g4�.	�rV�3 ƾ�¨K���f8Cg+�
���mN-���U�Mr�!�ꠊs$>��`�H��ƛ7�e�G�5n�I�t쨊�Uf��)U\F�j2+�����S�҂_m�Mv]@�/Cn�p�}xS�6�,�cw���v�g"�!J�� v�����������9g"����!WI9.�e�q�SK���Ť��\F'A�HS���
hU�a�;A�i*�=s���� ��k!�9������#��^�zjt1=�b����mA���|�ͣ�k	��*Wٔu㏹wn�Ǻ�GW^y��8��j��y0����z����'=���{s�и�R�F�+@A�����ﺜ��q�Ѽy$p:�CC��f�4�|(P�U왼gWC[��Q�r��F��z�1�:
t����sH|���rn�N�֬YG{�ꪯ��،���s�\�!�J;���t�V>�jL� ?����7w�_ϫx�,�z1�����J�ڃܶ���9s>b/��GF�!谵�sP|�������o/ t-c$��ȋ��W�a�a��T���Zx[�b�.C�����5\eT��O>n�w�w+�R�edE:��DL���ۮ9`�?.3z���|e!B�[����Σ���k������L1�i���ٹO�Kh�S�<ǟ��tŰ�q�L�su�j�\�K�cG�3����~Z��^��c����>�;e��4͓�@�U�/n6���=�^_N
 ���h�5FCf���q7e�iL0��Ϥ����t��O�^��T�n)�N�G9ā�AY m��@1���Zw�և���f2͗��!t�K>;�fV�	Kj��y�J�̖w�D���žU�@��ꨴ}Ϲ�8&@�� �٨���2oN� �D�&����M©�F�d��Oty��i]E���$v�z��Ɨ�*��n��6���[�06��\y�5�k�z���V�ǁ]��:����G����+\�EWy:����.R]�Cĝv�ͽ9C���Ӊ+��}�(����G����g������&�[��-�թ
���\�'OMG3�T��Ps��s�]ג��}G�{u};�[������Bn���̰9�`g��R��q����tz$ ��3��-�w���u�C=�=Tp�q�F�]!˦��Sr���b_+�5���n�s܎��r�Z�[�]^O[It�0ri�ʫ5	��H*��G��]�����n�@b�sa�!iW��D� ����йs���P{���]������װ�.���q��U{Mbq:ʍuLJ�U����%&��B�+���Pxx�yF�j�E;S����M��ׇ/]���ڂȆ���]׻i&��j�;����c$P:�@7fa�&��ϩKT@��*c �S���K��Q���9���Q��Cu���E�k=�a=���k������pᑑ�SGo�cJQ����T��:���t�'3��ls���Ʋ�vCZI�t�q�>��v,���վ�$�CW|�Ln��ed��s�M�4C.�L��T�gʶ�ZS�a��Μ-]n���[��7�q�L'����eZB
��C���!(�D-v��RY�c!��\!gHU���3xeb���P���& D�G��T[��f�,�l�n��Ǆ��[�qY�ױ��N.���Ӧ�P�]6��׸UL&�n��s��}`��9}��>���d=A�1{���B���;A!Enq<MCW��e��d�M�kjN�)Y0^�=��y��YMVj�h��q���;���n�@73��|j!J`k.78����N-Ӎ�Xr��vhS�F������1��>7]D	Ί� k�꞉�<*g�
 ��Z\�}0'4{ޝ�o>�;��q6��O�4����e����((������R-޲��]��J�rj��;\�c1�	�mցr��N�C@t6Hg8n�?r�;B�i�9ʋ�/N�����PҘd��AHNh�)ݰn%V9�����dukՂ򳸷e�x��Ҟi�c��Sa�J\��r�))L�6��9��ր�"��@��^-9�[jO7����y�a�1�¥�a����n.�y�:����F����&xUV��f"�Ng@�Hʕ4n�u�Q7��U���U]�0]�5u��aA�R9w>(�6�v�=�&��j�"��s���+M����Z|NX��d5�״���j1w�A� w9��t$=ۨ�qe�ҧ�mtK��n̟wUL=[2����d���~�P[��:Z޼�m�;ܺ.�6��&i�8%�;��رNɗG���
��3���e�A&�*�,�d��o.J���i�zw�Q��v������u6�[�f��@v:�+�� *�N�J��F�
}3�Ҫ���z�Y�H��m��ݠ�d��Q������33x����3�{���p�PU�[;_����`YA�}8������\F=���0Dϯ$�Е;s�q����u{w�4�܉.9�S���t.8��k���kˮ��	�C�[+ie��\�!'�K���k��tN�cK�R��xl���q@���7)�}��c�(���S�C��H䮎��!Lf�NP�fx�{L���A�M�N]e
�7����5�3����}��$8^X�`#������Mj?]V���tV�C��ƕp$��᝺��O6��Mua�uO�h���gm�p8j�p�QF����* H�~��~��c�=��B��h��6����J�Q�|�)��n��^�"� �(M7T\�  ��OX�y���iu��F�z�^��~��������R�"���7Dl��F8������О��AU%�J�$!#�+�+K��5��%��d�a�h�Xs8�5�ҨI�m�)u��r��Bכ�!$zo�]�_.U����a������!\Ƥ�����9u��@TY(F�飺����2�b�+Yޮ�v8QVN]�%���:3o��,n��h�W�Qj��P,X��$��s���
ԁ"tʱq�l�Ν]{�/���2^�6ؓ�j|+˧�!��D����E[-�s��c�%���uy���fW��3{��OWE�V�����f#]�Q�P� W<�EA?v��b�mF�R�՘C��z������%�k���w"�&B����S�
��-#�tʠ�����L��;�s��R�.{��)�V�,&`͞v*�:��()ٸ��T4.�Eid����� �N��J��Ż�O�_���7��*#f�̽�2MBN��̱[��vh�{j�W�0V޷�U�l�!�������jng
i�ڡ�o���S\�X�y���U\vTX�;t��W�w��}[��h�0��d�9q��Q��4��O��WTup���Sƃ��ǟ��inԾfM�ӂSY�}i���y���V
��`�x/+~\�d>�@O��kf�`��cR�3 7��P��)��N�5�#8�&��E�:`�Я���*��>gvT�Q�=X���*H�ʨh����|&��� �)��훔�aA��D�<���f�c��S-��cl�:2��L�L�)��76{A�_\�V�'���Sa2D���^ϮI ���eթ0A����}LwKP���o/��w�	ze�K9r��x�M��jzn���y@���R��ySp�y�n�Z���1��]1*�l�0i�8}�Yj�X
Lz2�Vڒ�s�Y��m|��/�L��L�}㚖D�⪪���V�h�[���9�ԏ ���Cx��V��&W��0��>�#���gF�KR@��T�����y�E8#���6~	T��lv�!_N?_�z���9y��"tD#«z7�\3���0C��D��+�d2Q� S��g���|��r��.�c�.]35�9��FQ)og9Y��p`qҕ�r ����EAv�&�Tӣq�$%bx�!�#�U�f�~p�C�v�pko��ї�Dp���\K�fX��"0忯���Ȁ�P�[iWv�d�ٙ��:��Q�w���E�ѓ�F}�������"����M����+� ��#�G�Wݏ�JmS�b��1QC˓���}g*��
�,�z����xP6���rk��׈D��'�oK�O��*-h�B/��@�ֻ	Âx�^_��^���I���W�������ӛ-U+����6�|���C&,C��
���~(�7��H֮��j+�}ع��q��n�ͮ�g5�3�Z��Ld�B��4��+�x&T2���=o�uq����iVd�/�m�5V5r��b	�V*�VUk�u�ï:Hh���H���ј�F��N�s[5��[�����z��r6z�:�c��f�x��)L��N���k�eu��)L�f�,W<�5����EZK��7��v,EƜ}��������t)�� ~�oA�y"]F3��٧���k[t�Y�Vٟ�I:#�Os_l��/��ۉ�曩�x҄7����6�*2�r�nkm��W�G=���ˑ�<I��S.M�a�"������� ����}:#Kj�Y�2lh�7P���P�sۂ<W�L�{���vf����	;�$u릐����N68.+���膤�����	�PT��e\��M��]�8s9���Y���$�`t�4Jb�f9����JPc �ߘ*���鬑��r٘����Vs��P�W�z�M��}D	Ί�*� ������7	_`5�*M�٘�����^G��w��N��ɹ��Z$*�a�R���vwv-��Ԧ�	�&;{j Ca&��;\�c1�	�mցKǑ7dHB�� ��0ț�+0-;T�����nJ���ǹ�[�jP���[���BwlU��z�Ƭ�u�vm1Md�T�?���?_�m1WR��Ҵ�w1_r�6�ɒ��� ���:��rQ���7�R�d��rB�k��U����OqL;���o�+�[}(dry��]�����E�.^����Cw!�H��^^��C���@�ZhNǬ�M�z�8Y��ڰ�u+�(G������7b��S�m�i��|�UW�W�����l�_�<�?�|�_O;z��U����r�~t������g'w&$��x�5L�Z�v�w���qu����t�o�h�b�y�U_ƽ__)�O�<&����Wx�һ������"ES�p�S���0��ަ�+�2���81��.����n���K*�M��iQ��*7.���2΃iS�9�7�ݯ�̹�:N��EWa~���-y˚�M���<5?��4������S3Pc_N}�;�������;vj��A��\�T�[SZN
',����qJ�L���`� 2;�s,�S��W�ؽh�kX�my����x���R�#�*�i��o����iz*��  U�+9P����GR�v`�}�Ȼ^ɾ��
��>�����!w�
^7��P(W�p]]�o)]���exD�>Fֶܚsܬ�5�S�`3����)�G��4؎�$�@���1�f�ח��4�^�if��X�pЖ�[�,�7n�����>�Sc`צ��OX����	2b�OnkՎ�v�W��x\m��ey����s�,��EI��ny�1
�g)V�WH���vA9r:�`���MTLlx��޲�f��y�Wh2�ީ݂�F����Z�D^����3]2b//gWvt}�%�-��z�R��X��W�UU}���K��o �Tyz��0g��u��Pg-�C�����`���4�Qs�)��͋oo��n� =C��#��S�<��-�H�C��s���nȑW*�#�O5����j
><8)T������+K��$��*�p�;"�u��e��Vzpw���w	�����y��TFD��uC]��W��	��w��Sc#��J^�zge�u�wJܚ&��\ՖY1�����8@�r�=Am��y6Q���s�Y���K����rTm8g���������ȁKjZ-����{!��;��r�ݻjɬ�[�s�8f��#�	�����k���>%,�u�ө���Q7�_K���s˝\$�k������ӜǶ���-h��8��r����̢�3M�TD�_v��|��3�,�����z�k������E*�n�W_8Ǚ;kes�ʕ� b���~�T�ͫ)�\v5}��oh쫵�]��]>FRۀwes��'R��*E\�ۡo&���v̡kK�k��i�m�p���,uz�ѥ+oT�x�_)h�d|��wa)���eMO��9�;�*V�1���ޅ(c,�z6>ĺe�u�ެ�W�koxH�ne�L�����{ݚ�X�G)���hqq}Vo�ڽ̱��Ԋ�萗�SI�{,v�r}�nȰ���=�u
�0�I����N��X�\fpp�C���>0bZizبf���s�ds��F�'�Q%t�cco�|�=��	f�d�v�P57�e�y�*��')|�[��s��J������4��M	L�hmK�*I��8�囊��Q�hw���B����Xᔝt�拙kk����-��+Ylu
Y167L���a�e(*�$�A.k������e���ru4� [��-���3��3W_�
���O���ӽ�t��֞=]��P��
��o�
��ق��d���jْ�Ry+	�u�ò(4A>Wh-EVT�����VѮI�����e� ٭s`���,A٭g>Z�L]}�U����y�V]07��[;�n�E�{E,l똞�h�;��a۸��kmR�f.�e�8LR;v�����E�㽭ϖބ�s�b��Q�qq��3!v��|�dདྷ�^7j���� W:yu����\Agy&t]A2h�ҸK�%ss��4����3��ki1̈	s"�q�w�f67��S%�Ka����p�/c�G>j��9�=@�hN�<\rR������-ȭ42뤩3w� lYS�߶?�����<I[/ж�ށ�>������a٤�\Ou]qb�Q�����z��C�Ŏ|.���?'����]M׷e�0.t�V��&#�Vq��{&(g8�hPwR����
��]3%�%�=�8�u�A��#�H�՝����Q�k)�q������f��I�0iғ�R�e4�
{�ܵWZz�.����q9t�%I��u]^�om�S���[}HQ�難CD���;��|�E���V$9��.�7q��v��|2U��V��)-������Ң������vkl���M���f�u�Z�*�P�^wB�#��5ٮr]򆜫�cz�f$���Rj�V�]�>Eg.Mi{ˇ^��[G��j���j�>��<8R��޶{N��8[��·!�-�CA}ם%��X�k`)��Z�J�H�u�;�������ۑ3[ب��Z�-"h�2�%k�J 2(�%��j���΢�s��'K4��bG]@wU֐�๽B�Q��X/Bd3R���F�����]a˕$�yH�{�/�Mڗ]K4e�r�ZȤ�#M�s�z�ҹn_m��y��?(����:�COxm��ۙ�I��l�{�&��r�Msq<��SlA�z]gGa�K�)qOg5�Aҋ�M��1X\��af< ���q���bL]�!�\F�/����X�����{�^�����AU��YUWYPU\��(����H�Q�9�U#2"�YTUW��s2YY���z�JĈ��f\��$PW#�E|�W**�D�����\��OV��"��T��L��8QΝS*��U�QYŏL�VT"""�"�E�{�UG*>S�@\�2�#Y�ޙD�As�ttљ���\��Eh��\����ۑQUw�G*�*���Dʪ*��G(�93�UȦT�q���/2"���%09QE�UQE\�ZE�S �
�L�r�͕�K�%�aT�Ep���GQ�.ab_^A¸TPUE�(���*�(�hҪ��9DHN�!<t"
/�Fr�tNˑW9�J�D]��,K��8A�Q��.UU � }B��@}n>D��\���x��W�o/�u��zGvd�(ג��):�c*u%w6@����s�&�~��p0��4����v����W�U}e�Ž��󅕑� ��%�m�{�U���E\�;ξ^Q���'m1������X{��sȥ=���/_��}<�W-���%�"=3������Б�yx����+���)F�OV��ŧ���
���g�Z��B��ݥw
�Ӷ=_4	u6ک�������=m���Ͷ�=y��*��T-�O<�ٱ�1�:O~ݖ�oT���R�.ֻ!����7;��dn�� ��xyĪ�l�T��?�J+��l-��z�iJ����� ���v�ܴ��ډt�ARG|���J�p�n3qqغ�9���R�!?�\��_3�T6�(�f�˚�F����(����uڅ$*:�S3����*�2�Og���s5��q��G"S�(�f�������b��������'�����ky*5i0i������"�؜w���[A��W�Mu<}vGX޺�۹S�y�;����HK%+n��x�앏+u�^��Xړ�#5�/*<YC=u6�œ�I�F}:$��B"L4�.Ʋ�S��}�< [��:u-�m��m' :���P���9��b�%'�qjtg~��꯫�V"}��~�Q����m���c]�O��Y���9gz����VM�ş=�P�{5zҋ5_&:`[��f*�^eD���2���{r���s��&�f�y�n�m�b�*�t���̻�zCxIgڄ�i�/��I�X���徫ϸ�(nit$�c;+�z�\��n�ce΂K<�P������i�|��]�7�s��� wD��p��N֥y��m��E����ty犍�k���xy.�S����nT�N����gr��"�i�^ls�P�a��Cjf⪐�\�Яw�X�8������-��kb����O�Z}������.��ʧ�m���Ϟ����/� ����%���qu��>^Xٌ|26�:o�{{&� ��nq��.O�`��U'��RXk:]!4MV½����
yŮU��nr��>��StފWܧ�BQ07�K�����9k���2��s�j�s]����r�n�a�{j�ilS��N�][�F>��P�'��q$�����5f1���³�:9��9��M꬧Z���vĢ|��N�9�yK*1u9]��p;cjzu�wFb�uu�`�]�E�L�ɽr>�L�!��G=B���U�U}��Ջs��)�[�ǽ<Wr����xΗ(�7!����j�ZqY��Д��us���q۽�BM+�s[ϙ����D�}ŹU��·^��f�p$�8iI[w��ж�[|��q[|/k��ۇTҪ�
�X�$<r��Mb��aWܺ�I��9ݝ4h���U����q�j��9�D��TO+s��Pے�2�SɬY9�i�[L�]4�����^��(�p�C5�n�59O����C9��>�ڥ���U�"P��س:��	e��������r�&qCR��S��|�U�tv�^n��Q�y�)D���]?eֻ��V��'���=ow+��u��9�TU��)�$���'[9�f�D��Kc� c�����L�=n�����5���ǸS[~���FNw�?}��㶨���5���gT��ʓ��K��{��QL�M�ㆍzB�	�T��s g�q��ic�\�g()�l�1�И�r��p�3��E�����dd�KwJe�7N�-�S�n[���Ԥ6n��n�X�u8*�kgub��*�yЧk�R�a�g����㨕��f��a��W�������2���UEg�n)�vm��4�I��l������}cl���F��h�S����'-t|�>~��ݫ���P3����KӞ�8N� [G���<>�iv�O1ܮֆ�އ����9\i��p
`�ϑ���w���qU���m�.����2����1󮃦��צ��t�c�}�7X'v)���������:퉈��R����Ww#��!��Oʏ��9S�1�E����|g�}�Li��O�5>Y�檣޺��8c���`�����T	���zU3E�\G�Di�jV����BԹ����9ng��ө�Lr�h����w�7L�R�q�mIZ澕�5�^�����U4r'$�H��'{�M���l\O���\������Bo�N4��N��\��e��&7{�Tk�N��k��)�£!�'�V�Y�]�m�>�U�;��W�U�,!�E�Nױ�]�o+)�8��H]Ω���j�/�_)\D�~�]BP������M��+&,*�|M��bB�(������<4�JΙ���L��Aw��8#}��r^�����8��K������+��z�����e��X��דYV�y��؜3V��Nv�ŚQ��6���wm^[sB�^8��m�x/"3��e֮%�N5,*w�pY���­��4�uj�7��P_Fb4o"{�3�lEc�)��f���oi)G�������3��zE����4=�Rj�n	�v�y+�=�^7���貚k%�m�	�W�V���T[.{FZ����:M��IJ��:wo������(�Ϯ�Rk'���3����!����ݓ�c�"���N�撸��ݽ�O�OyNr�ASfg���t�ݢ�ze�Q�,o�l��4��/��+U4�=|�����,�7�p��dcF.K3�`������J�L�]S���t���oS	Wt�U��Y�]��N�^?�g*U%l�t��0cO�(��o>���{�n]lc �VA1cg�����r�W�t���n�s�f%}�һ�o[��a&�*�p_J<��g�Lb����z���]��bnT�F'X�-�uy$���ҥ��v�Ru�	�Uh,�WG�h�qi-QT�'^cz�����耣��>�[�_}_}UEH�܃}��xl��?zx�[5HU�ﶇ=���2�۴U��:��05�;I�W]�>M+����loͽ��S.xтTla�BY��\������#���5�����ܹ���2�]�#�?'lQV��y��X5�.w��;Ԏ�ʒ�IN�1f�ˤ�I�M��p�Ge���C�cZk%t;��46&����~�[%���s��o�|�jw��6�k�gzsSQd���FT������^�����>ۡ']/It�	s|��󤷚�%c�����gy�=���W�G<e�y��o0���_O�1T���V�;[�:iw������pCX��^�m=w�^�>�{vo>��2����OY��Φ��c�%�绫��+��d���@���<}�����X�O_�c��9��s�����S���&��^�C}R��c�ss��W�6��ڝ��˛ݦ~�v���%��ݑ��F����o�쳚fJ\��L溎gL��V���ǒ�;�ز�GӺ��S�����j�(�-�D3F�&�:t[���	ܤ����o��)����Y��f*NT�ۂ,�AFbk*o~�y��7Lm6G(~]6��;��J<�tė�����lT=嶟:*ЛwJakDļC�M].M�uc�.x�; >Dw�O)kyp7oj�P�Wfv���IT���{p��6��� T=��<�J:*���v�)��;�����O8�|�7zl:�}�N�	A�8� ��0F]�r��h�*�X��)]֎>܆�EC�t�G!����#*.i�Y}���͞�E5���E����c�B��V�kle��C.�f���N��k�fe��s\R#���0�[�	�vhT�3_6�;giK�=�q��9������ǜ/�G����K욌Y1�®]E�,��U�I�И]��v�f�w(�q�k���nz���c�ʥފ�C�kEJ<{{ �Z�7�n�ֻ��֜#I�;MNS�dO��E���/f	$ԭ4�c[Í�b�:g]��v��$9L�;�1���� �o]69��z��{���{ɧN��/��F�`�vK�^��4W6�����%s��K �ev�2n��,H�w�L`f�-ޝ�|ƹ��_1�;�J��^����:v�~�����w����OUz7r~˫{�oF'�����.��!n��*�6�[�\�z{m��|��!�.%fԬ���u��镢�|�\���r��82�V�=S7au���̋�T�f*��<�h����y���7��t��1�i��/!�W�k�~����`̢��˜�P�1Gh��s�ƅf���h���yh�Y�=<�nm�Z����V;���D>ȕ��xV�p��;�˷�Z�0���7�i�����l&�]�T}P3������Gm�ۛ��WW�z�.�\�F�]���[�������-�����h�E�SAje4m�1���/H��),(�{�k^���W��z(,4�"�w#�9��i-f�G�N��/.垘ܘ]������-�������2�y*���9�9<���\}�F�?�O�4�K�O�`-��7U�i[9��%�~��iH<۴���:���������GF�QR����#�d�^��͖�
m��t���B���YOc��Pj--Y����.�_clYG6�u$�8�.��S+#�4�^�te�OM�{�}�i�j��G�57b����U}_Ul��S���ގ�:b���q�<�ODy�P�SX�:sW�=�sov�wJ̚7�8���&.�G\q� mIZ�%vL$DR�`�����5�X�ld����Q����q���l\O;s��/�h�j�[G�r��;����c�J�,OvN;�v��Ms�_͸�9O���VOs��S¹��)rӱ��S�j�VeD�=�{�ky�tbp�[�v�9֡^���X���Iv�]a~��m?lz����K���i/q�Ui峇G(�i���t�T������{����?���I�k	u7�}q��a��7����|�l���+u�|�n��Ϳ��Y�75T=�i�t���Ȧp�+�'�}�a�nh	s�)�����r�ϴ̼]�@���T��iLk�K��o8���+��'�ss�SM�Q�_&�z���:��D�Ux��e�=������;����e����F43�e�8�׺�vi����>�;b�_;��=hfx���da�������iw'�[��h`1��$�]��5�k$��eU��,m�Nϋ�~�՘��#���(���:���YG{���">���1��w�����*9�+�n�!�o��%�֧9>k�`�U�5��Sڞc�_
k@�; w2�/�µR�<�|�zت�㈚�1.�`ʽ�U�M��6D/���Drk��7˦�X3|C��B8]��A�Μ�N��t�����%y��Z�qe�-�͊[�y.Y��<�������ڗL�RG|��=�X�7U$8���j�jiN��=�|�J���lkob��j˞q���B��1�f�5�Q�^\�}���4-�e�o��sgV����4T� �����WT)-��mO�nM})��b��x�)4���q�K�/�b�b���=�Kf�_!p�)Z)�@�u=�R��b��:�\oz�<��j71�e�>�N���rʍqf�X���b�y�`�������ވ�`�"���9��)��N����������x�m>�^�u�:�>��IH�;�[����8ۉ��8�Nt��}r.%�����3D׉�u3����f[��E��s9�R�ެ�KO6jPw۹S��g��'.��8���i�+״�ob�vn��q�h�K�Tƥ���ΝZ���c|�N�׷!������&�]����-]C]�EwG#V��jX�0�>S9����9i[�J�f��i�j��VԢ�$Cߔ6c�MJ�:3y�zm��aQ��1Jd�U�],�PtR͡�ֳ�Xu���'ƺ��v����cqյ�E�8��"joM����K4�V��kC��jD5�a71�5n�K�gq�gK٧��E�=퐇|@Ǉ*\�3�U�73�X���
��dvx+W�ъ�L�u�*����dM�dix�s�13WYN$F��3v��L�|�1C���q��^KoM��8��ͬ��4�k/�⺈u��L��M�͒���Mn���vF��m:����s�-^@v��%w1�t@�F�WSj�ѝ�{�ŀ��qs�%n�l�t�a�)$h������/{���O�)x�.��Ӣ�,Lb�׃d��+����m�Q�J�W:�_M�q9�8��6XNݑ@��3W�4)n�u��om�8�+N�\�'�]����#��ހY�бݗ�I�%��G%��Nub��)�� ���]���b���+s�m��[��Nswörޡ�+8��Ò��!\�nh����p)��7}(h�O0��sB������B�#�� ��/V4q�Si��2��u;F��f7����t�������v$�\C��ъU��̼�;�:˚�v{���4p�&>�r_dW�MS�W��_Ge�l��}�2���̩mN�s�:�n������36Kw��c8��+f���#�чe�A͕� ;�D�SgY�1co%�\��A�][�1�������[�a)�.�aw۽�ѥGZh�8˱vB{��;U*m:����v��:��n�s�c'T����R8���6����W��gT1$��ow;�wvzh��=q��f���=3v�S�N֜�{����PG�u�;�L�EqI`��.�"˫�[wM���Qwf���B�ΑM>��K	=�`��l:&t�E�9��6�E��_1�\�ۭ݇�^W@t�Q��/%��Ku�3]�e�U��a���y��L��]Fe����.�KYύa��Hs�V�!r˲EЫޝ��t.�;Ẓ�ӊ}-�ب,x��CF+.�j�F�Mq�hq��>ꛘ���*�C��Zg18j؛N���W�_N�æ;�鱑�v�"����ڵ���]qS�G3��Lp���}0�sxWP�g��1�;�d�	�vsu.�f�����p(��^<�w֛K`��L�Y+�	��ɚ�E".t]�oZ5���;BJu�}7��\w�T�L���Ar�D����ՔEU(�D@y'*�UT��P�\���aDE�A������r��r�ke���jkST8g��"�P*�J**-H��A��DA"�9�UR���Er��E�$"��t��`r��r��p�B���r(��X�W �as����(��� �M$.TQEAEr�aW*;"��Ep�(��y@��U\����tp�TPUF�*"2B���EE�B"��0T��*�
�UTNeʢ8QȮr<�EG(#�DQ�遒���EUQA8p̢�*�*"��EI#���UQr���@-NW@��
(��s
#�UT�r&Q"(�TQ�L�քz$Er)���*(��0����y����TUEw=ܛ��*'P�EI�ǽ�?�����ށmf]7sWE��^�\�*
C�_2M
�B,v��+�]:�ؓ�#��]{���xz�%¥�w�W��|7*�oU�ie����u�q���<�'a�Ú�ޗј�m���v�*�e�ktM��xK���/��R�_�=w��{ϱ�6_WA%�w����^ݭ��/&�Gn���j�.z������|�৞��k�{���v���F�<>�Ú���r��9j��fU.�GC=Q��_IѹȦ��]���uݠz\;sxds�\����i� �� _]#�t��_5��	^c�իu��N�:���_�R�<�:�釮��=9�!>��k��f���&��jl�8\�z�6��)��#M�K�C~�O`�m�p����H�r���IZ��݇�w�ֵ��g<�z�7��_jGc�h�����4ɴ���d0����ǳ�Wr���;R��{3N^��C\���Vn�G�g��j�[�vhU	4�����߲�/xW�߷{�e�M��,B����[����zU�m��[u�Vr��:[ç��1v�7
pӕc���;�S&J�L �z���^������Y�NِvU��H2�`�@��ï���T��J�s���U�[D۔o1��c���Й$J|�����o7CT��GwmVȀ�B���l'�V��{x;�Yp������	'�8܊��g����.7l,�`֏o����b���L*)]8u��K�6Z恤�k�q�⣝9�N:j�L˪]�Mz��uC��&�8�%�K���ڕ�NM��jr�|,����g:��G�f�6����l��)ެ�˫w����ᚷH����5�n��2�s�1p��

��O:������o������˭W2�$��}.z��G��[q�*�&�{�=���=�$����؍�ϧ���{;�L�)���p�˕�z+�JUJ�θk{��,�|\���չ�	��a��jod�V��[]�xYYa���}�iꧫ\|�H�=h�H�:���u���%y��T[��m���=��6�}r��7���j�U�"�>��g�-���ֿU�s6�Ӯ��u�WN�s&�,�ss�z�zN縩�9-;�a��#�Iq���gT�#���B���gQ8ђ�]yڶ�E��j�L�<
���ud�@�qL���VΌ�F>jN�b�[�&ٻO0��o�����
y�:y�>����̙��!�����+�kwp�7�C�m=�9���aWˀB8}[*�,�ɺ�q]kG��-�Iͨ�ܮ),4�<��[oCלm�k��,���2/B���9}�`��E|]%n���JWu�8��xl�Ln!/3�N������;�3Ժ����t��0cHK�O�b���H���p^F*��R�']�C7/xe�	��-��#�!��
�'�uK��E�t���6:��x��Sz��	����5�
�Șn٢���Pژ+\���vS�j&�˝t��j�L�������jL;����r%�q1�����e�d(�"nGAKt�(�pw�
W;�����է��#j�'�e��W��nR6���S�n�VeD�{q�&2���:�N<_���J�鬮<�f.��R~��d�W���i��}�����\�*����ꕩ�Zh���-����^�NL�g���O+d������t�g�l�t����⣏�$�Z�J����,�`����S�͞��	�*���n���:�R���o��cZ��RRQ�*4x�a]���$�+s�ɦ넰�fұv�b��j1������Փ�}�?Uw���S�����3���{xf*�������9C0�v�^)t5U��#g���ꋈ+���)��u="�a�G�޴�n�#�J�4�����*���R�}�=����Y.�n!=�z���X�*�~�󦮡_��T1o1ʟ�*v�a�a]�Q=����i��_>�9Ԛ��#&�1|�,[e��7�^ �w�:��=S����w��7�S��Z|������W!�������cj�`�*�JU_+�j��Z��>iyR%���g�o���<���p�[p�۽6B��ء�'�ү��w�RXmqUb��ì3U5��o4��Xi5ڟd>���-fǯ��r4��T�]�a2D����x�JV����i1x���*3����>����8�}%b�^��<�y{���wlGf�I4�!���3�W��د��f��ϾsD�]�(�����,�bWk�yz�<!��Xg(#f��c��w���V�J�rʰ�,0��u��٬��#/�w���/�9c9z�({-��R�ᡧ��ھ�ZR�o@� �R�7�yeևm�`�auZ7L�;F�O}�;�MY5�;Fw��}U]�W�r��f�/@`��jV��b}���j|�.5�#�D�>oe���3�#j�U]A�U���ѵ0V��Jy5�~�x�9*5�M�TָA��z6j��e�����W͋�TڱO�۩�����x��o¼�a8%�����,��B]շj>Nr�Ś��c� Z�������\:(�ʦ�
1U��뷳�=��u����g9ˎ��̻�l���A����a�ks+�n��^�N^�W�+7�b#-s���q�^��f��cG�*��uĩn�~�n�[k���v.�8��x��泪��R欣Y��<�紺yՅ�j���dJ����_Q?w.ne��s`�����AIU���,�����\� �/�TrA���-t%3k�4�����h���>�^�K�YgL=t��=9�#Kӡf��j��O:�Y�G�{�O\]\��(�ˎ땍��N���]��j�f�Ub�7x�bD�5�ks��p�����ɧ��R���z
ti����X�2���.�O;�M�+��|O����|���w�ak��߽�{�Pe�(S���D}�Kn�S��C����o�M�P�6(w�{x�1�_0o�g$sS���ۮXQN������:�qʈn���a����A��mr�}ڷ�zp�� �Ŕ9��jԮ�-�tC}�����}.���
�M0`X;���U��_w}��KD-u�l�١T$Ҷs[�gpSӊu�Q��'=�ΏAV�|�J�����I[w	��	.f���^93P��h����v�D�ݱQS5�.����K�Wn/T�o&v'��ؚ��H���}�0Sq��������}Cn`�̴-�W��]7��Q��N�{��w�)�Y���"���NS�dN��-nWI�D���}{�n�1�.'3
ś�'.�^����n���l5�lg�k�57ks/�жm@�F�l�X��֮%`�I���S��Ux=�=y�r9� � ��۝i��.���f��R��_/�+#�^i�]�h��j�'�8V.\��6`/6�P���Vv���o��N��#+��7pd�m\�lt�d�
���	'�Y��&��L�3R
9r����M��{-��UW�^s�q�D��^0�꣭N�MK��bu/�{|�-�k��2��Ϻ���2��t�J�{�f��l�]�����Zc��uz:��Q�n8(�r���)���_�r�O6�{7�hJiғi�6��rl�!v�%q(�D���%*3çv�tO݌�-����/=]����BTo3���b�\����w�¹JƷv�7��=m<��'hc�σv4��=�q�K׻<�eA��_IL��RXj���km�{o��XX��f�)�Ė�Y��_jg`��~*���[4�w\B8�jY�f\]u;J���R���r��H�Cr|��#a/�=��f���^3�RO����Zެ9n#�ry�
�m����!���4�}%k�b�!���C����������ZgW�9�9K5���m>�0�g)޸Yev��ْR��zlf�r��4��;b���̙�M�t�vTv��F�Y���=殻�^̋{2
�x�����7��������P�n��u6sIZ�^��0��.u����9m��vv�kZ��[���(���"���*�[){磌�s����o#.������:2�a��#�ب�v�ݵ�#Gp�m+X6�#eEӂ�aN�cLv�w�Q�Nm�>
s�{:;�ӑ�Mb��o��hmz���B�.�G�K�_˧��EQ������EL�&�+F�V�>\eJ��8�Nv��5_k"�P�U6�`ʌ�?e֫�l���r��׸���7k�58{.z��ܯ{��w��03M�T��s�V�ʞ���G���f��>�Ք{��]�1��=OH��nUj���jU~
��c��D��4�u8��ځ�����8��.�6!=�z���V;�]��7�����>>Ng1o���o/iJ�Z}�z�M�nr�j�uϭM��q��lk|%^��yG���q�S��̇�*9R�JƷv�7�Sג�\�Ê��ں\��碃ߗ�w���R_+W'���R��*�����AK�cq�wN�<(Q����Ss4�w�u�����3Y)���X� l��Ƞ}�u��F�g��n���ʐPV�c��v��9�շ[טuwS�(|c�N%��Ƨg8�Ec��.�)��c��W�/�}}�vf���CE�\z-��smޛ
�܆�|;����Sb@�Q�{�E�&:�]Xl���ˎZ�c���t��͇P��&4����e�:�כ��w��5ʥ��صۖ�������v��L��H]��gP޽���j�p����nK�|��>��Щ&��/���q��@tΒ33U\Uҕ	M�����j�%m��'1��Wܹ�m�w��}�>cG�F�SOK��%l\r8��6��$�sj��׋���b�޼�Q١R9o]�Y�wz18r���v�X�Ѵ�'�*V9�ŒF�16��MkH^J6�[�u����8f�ہ��s����U��E�fs^�i�m05���Ҝ��3�^��]Z��}�Ƶ垸{3ݕq�f�+/i\����c���2���V�����R�[O]��^��{�s��=m�����k*28�.�2�9C��7�����ĲfGi��K̤�~F*����c�����M�ܬ��tlt�{�19�ܤ��RGM�>2p��e
��\��7�tjP�-4�ұ��|E�u�Iv�V�t��3-�kg���Dr�34��~���Y���M�ƆO��by���lv���b�Py�)��o7��ӆ4��~F$���:��*�➼n��P.]/)t��+}Q��Wtqun�L!�c2�a\���*��*����\L��:�"K⣖��i�d�쭜j���5���{_ɧ�������ޚ{*���!\s��d�yy�R���.V�v��qڞ_σYoCچ��m�\�;TJ�Ӌ`[���-i��C,0ޑ��ԖR�\5�v}�s�7�7M�⫉�wՈ�+�̼�7o{�[���?���$s}7l�=�R���ې�h���(����[��u��ȸ�#_�l�J*Ƭ-��Щ&��9��
C4S
�Jl�Yh\5�+���{S9�*�����i�/Et�����k	w�w�>̲7d�.̚6\w$��0и�퀥���]Cj~+\���%�juR7Yϥ*1<�YJ��ZĲGbP�i t�$�Ǘ�w�{+Wt��W{�Mq��z[r�o�����o��;���Pu��!���3���L.���3#ѝ���;V5\͝uc�9�c����3W=ݘ��R�$�]������LrA;ܥX��-�[��M@���H�j ��Z��zd���.e7���=�8g_!>�'>T{�*�N��8Æ!��/Q���KY����[Ҝ����<_L˰yp��l���;[�eC��3�1����٬�la4�s���+���9��kU�E���V�����
�6Z�ݸRĺgT6 A�ՙiv�o�s���I�N���V��-0�+����N��^��p\	R9)�رy��k�`'�9(zW��a��2x��k��2�Yz�=������9B�qV�I��rG$B4q��]�"��夁��4m���95��0��}u:���ӎ�_-v�aC(VWrK'Z�� <�e*�V�^���R��gդM�wSs}�|��@�85.����Ź��I�c�Ky����c�c[��N�SӮU[��n>Tk��>�]G��.:򦲰��xYv	���:���@��A��+���E����䆦ae��enmv�:��l
ἢ��3���G��:ض�F]��ˤ�8�T��8�wZ��l�]�=M��J���m�;�>�؇z�4�fEt_�����0F8���W%n�ݼom*&;�>��8��-g^(���ܭN��nViLP�|�e�b�w}Zu���i�gk9N�wĆui�P�qv�7,�G�d{�7th�*�-�����vܝ�5�����/XO�Ύ���u!�ӻ����x�wC�s4�6��l:�]x��U�9A�J�g���)O�:��mhk�����O������k��_C��˅�v2l/�uwD/N�,5]sp�s7�B�\�������m2�
u�|]q1X�����4�����Xj�u���Os�c@\z��>�ٙ��z-�>2J�8������t�#s(���\��н^�1����7)�ӮC@ۜjUї�DCz�����%�!$t���x0K6Y����뷴�)�5.t�/����f,}]d�:^���z�CX��Z�ŷ}�owDʐm��z����q'�\�[�^Zn ��38�$�㭘����a�l������x����[���fc�s��ҳ�S}�Q��S�O�R����*���+��JX�d�At�f�Α�Y+E��u��H��ȅ�喇-cb�gJ�|&2k"f�"�S���M;���m���ꏎ�.�bE� ���-]��Hՙ�)�v�>�aW9��}ov���+z�x7���f���`�l!�5�w+����N�*+�'���Ɔ6�!�aK���,gN��r�`�e��{������} ��fe�L�(��b�n�u�f��;�a P{[��\���w�fN 8���ռ�4��+�^W� ���T�r" ��#RT.s���QPy���I�~!Õ�T�A�D'M�"*�\��s�Df^YG�/E�EwS����[�hDTEU\���*�N�'0�U�&Ȼ�C�(�Ҡ�i�Nd:�Q.8�G"2H��*�r�����ʊ(�\��\�щUQ�r>6D|�L�DE4��AQ���+%�S�ĔN�U_)�\����Q�W(��˺-�H8rW�"����ʫΜ��E�L��2�ZQ��J(�A\��.S-�lJ�W
�A(����օp�'�&ETUȈ�9	9*���&VE�dU󻚅sRI*�(�(���w��(�x���)p�$"(�s��"J�\
�Ḧ�;N��$�r�Q\(rW*ߟ߿���6u�sVJ�n�]7�L&����&�������^wcwD[����N�w-�j·�KtU�� C�ޅ�R}���jE��m��c'�y���˨�I�I��c��o���z�����m�@y�&L�k��ͭj�,sݓQ�3��}���p�Gɸ:Ѽ�|.5���dC�Q���aN�IL^���V=�Y9uj���}x�3Qn���9Њ0*���1���J�9zq�?}����V����w=T2������yO:�n�q��M����U��s�Z�JxJΩ~�|�;&��d��V��O7�ηw9�.�Rz�'���)[��z^/y�2�R��"5��ݪ\��%<�OS�g���p5!�ђ,k�\����P��NFu@�]�{nm����ϭNuBk%�pX:lG+���-V�g`-q'U}2�ڹJ�kwoCyoC�m=�9�`W��;��Ӹx�v��W-L�;�IH���R�\4ס�˄iؐh}�7+&dB̕�U�n;��T{��o>jߵ�w�o�v5�Xp�y4�=�']w�c���#�;��t�h���*O��㕢��A���Cr��Mm��C慜����=�T�A�:0����E����%Jz�Z�!�_<� |^�{CF���θ�}�dL.���)�Z����l:�_r�������G���x�r��~b�Rt��ig�n�S�|��Zp�Ψx�T�F���_r��dO��]����b��r�8��N�k��:\��B��s����a;�`�W�����;6�&�4���3�+�r&�j �f��ƧA�q5� �������pw�jZ�����
���RL5�.5�q�ظX����w�Ҟ���OnR��L�Z�m��y)��b��ob9*5i�5����Q��nKz�M-��q�\7D�@��2�D�ʞ�7ٖ���?���]6�d����.���Gn���Ś��c�[�������|�UoF4[����=����b]�S�we�[��Q�3��2�>遘���y*̼�n�\���j�R��z�)�)�L�l-ǎ�wV�*ﻹE��Ft&2e�n��i�[�x"�]�X#���w����g�7��9j���լ����gs��WA�!Mk��m�/�
Y|����5q��VX��vq�ֱ}�{���4f��p�A>s�̴X=Yt� {غ�W�c��Qّ��%/���tf.c��x�-��ظQ��.
i���y�	�W�VU]���]f�jW��p�gnAN��=R�u��Ob��"�j��\����:�M�건�gi5z����U���} �!�J�Ue+��C��|`\K@W��t�<�s�5|O�K�L���X��?��:G��N޴qW�	E$���]����c��l�5�=����o���m��aR�r/�{�tM��ƓU؟��ɽݓu݆�WbXֽ�3����+fè_NTi⷗��(���q�Z�q��v��َǮܴ�!�׹��x�Ժd"�����˗��H/^�f�~I�q��sڲlvhI4�/��g�m�d.�*�F����URjiQ)�5�!���[s���Go\���#U����"{��p�y\�o6r&�(�f��֏n&�؟�ؾ��gW�d��֖�Gp�SP�ｵ���NZ�ͭ�ש��@�Or�����ڨ�m)��|��7޾�J2{�Yc�j�+\��ӄk�-�;��t%��\9j��b����.H�e�w�2 �ػ8v�����s��Pגp̲���j��/�����ZT��Kr��L����]K	(�s@�ɸ�qN>�;r�S�n�'�*V9x1�΃r�uцa��v�x�.��ڕu�'�[p6����j���](I�z0eG3�-�0��:���ՎoFTF%9un������;�,�ӭݞʧ��N}ih��2�v�<vVl�ڗ�3�n[�x5������}�ͭad�x�k�sz�o�xg0�����MF��:Ԫg@'��Q�g�S3lb�\1]dPކ�g��w�{�ު���늱�P{��z���T���IP��z_-|���.�5n�6�犞�=W�u�:�K��<;[�V]�T�Yj�����tO`i�6�_���o�m���郰j�� �z���2�߹%�oN�K9��r��ky>c��OQ���6�\�q�z�-dFVf�����qsk�=��,(�{�Z�>��T7M�չf�Ҿ%�ے���˭lS䓮nV��8�� �[-ΛR�����N�+�Iõ���]D�&{K8�v�%>H.�*�.M�x��ƪ�9y�\��FUԠW�{�ln+�ru�����r�[���z�O�0Z��2v,�K�D9�!�Q�s����0w梾Ϧ��ǳ�Wr�9��n4BN�ֶ�l�Ԝ	oj��X[!�����Q!cV�f�I4�z{o(�[�J�_݋���֎���Av�$���.�	���zmӍ)��|(�.�te,�K�K��l��Ȗ퀥���]P6��5�Y�`w2x"K���x���	���\�N�I�_&�]�Y�����۞�O���k���bLv��F�WxIY�Q]J���9=�"ہ��S��Cٽ��Rns`!J�iM�lc	��R�
ǘ������/��N�t��s���T�gp4�j���-�xEA�ؓ�����$�dw��R�e[����?vի�}��k�fOy��� �cӭ5�n	�,��"Ѻv�j�8�l�8���=|���[Տ2v����c�冨H91���|���hbsٯ���yt���!6ތ��e1���'+�����3���]�׎�c�.N<�]/ڕ�ݨJ�.�Km�HQ�si��D���ݔ�\�K�*�Z
��*���7i�1Ծ����R��)�VS��z��Mkqu� �{����^�������jT^xwF��3�{�8���u�y�	ꧫ_�V;�
�bb�[j��,ls�t#7�ץ���(oR�b-��i�������K�gup>O!챻��1��sH]�/�¹J5��z���z�x��{de`&�q���:��ڈ\����TIH�紖S���ք�c&c�9�ǜN�F����n��Aj�������!a�Ɉ��VGa�x��0�⓷xRޛ&���-��!���a���(�/g.�0V�6�;�v@�[�y�Y]��)i\3��a�q˦B!dt��6䪻�b��CS�Y����[�����G5�Z\��2�;gL\d7l�,։�]�Z�	ŭ��T�ȕ�5��oQ��I�\. � ʡ7'�B��sC�»sP�tm_�ne�Jy5�c�㿖�[��Փ"���h%W(���ZuΟ+��;���&���S�>'U�c1�fiO�zB�����n�\M�	0�+��xuL��Lgd��]�TV���*\��GK}bpN+˝7����םW��>o}�ַ��pEY�a����ډ{[�ޙ��U�|��4d�U\g~r����+sᖫ��OL�辨��W���-�_gf��&��]պGn��qf�5�����'Z~�K�������Ѭ��x̦|�}8I˜��/m'ޗ;��n{���/��߆�C?,i3���z�.�����6�{�X��u�)뿡9͵��1�N���z��n�lsp�>�eɘw��G.�R�T>�q�v.�8	��%�m���$�"5U��%�!r�]<��U�`U.x�]�2_F(�ZԿ���*(F��쇏d�.�������r�u]��m���t������s]�A���i��>+�d�J����.�n�q->F�ti���v��)T���P�o[�qěͽ���e�p��.bzվ[p�۽6���vḮ��s��9�m��sF�8�on"�aEu�%�vC�OʗI_�6=�N�o���U��#�6�!��u��:+7[+���۟�ga���(NoV��3;�D{OYF�n�]����/�o1��V�\ ������g2�P�ۘܥ�xw��E�t#DEc���jGѼ+xr�pCN�b��ao���4�ȱOv�~<�4>^����ݏ[-&/%�<gj]3����+FTJq����pO�������א��P�J���8�u���kQT4��A���:AV�9����j�5����ps��O��aGzX�~X�W)f�5��Z761��F�g"S�+⭚�T�+rj%<��1b)�{���q��M�[���d���4ۍp��>�����co�L���Ƈ�"�Y|��ԦK�ܩ��wd�mZ���u�/C5m�ڄ�+���wO�!�5�]�W
a^��yx��q;�_O`�����oK�N5���3+�*��D�/�y��m�ۜ�b���FgT�ډX2��Q���^=w���n
��Oc�������onke����|�np�;F(��>w=��A���M�����wL�^�۞��lM�؁p����Y�`-<�=�������[�X:���i�����0o�t�)u�3�暁�(���Oެz�.����1�ޚ�g���z�slu����D�+���;ga�hk�ʞ���GP�Չ̼1�
�,|��^��ܖ뜽S���O��R�od]�_V%�֔>SffoO�)���]�q�T=X{*�U�֏���r��sl{�{�h۽��*;_)޸�`I�6�\����Vt��Rm�4�eZ��gl�ۄ^z&w���4���������i�6��aD�	P�[�������U��v�S��=�$jdw=�KB���k��zl]Y�橻���d��,�\�M���); %y��޷�ǷR8�J}W�UԒ�:�J�[�����m��J9�u����c����T;�Q���ꤘ�~��]Ӈ1�q�M�����.٨S%Tt��#a>��[�lFVr�T�ŧwy�m����9s-�|�0��r'��*��!u@�@B�� ��3͎�֨j��r�Ǜ�.[%$�5	��adN����۞�Z��Ky�T��y�I����Ex�:if�V�#M�P����\ q�֛w���7#�f�Y�,l6f.�b�J�ԛ�;q>�N�,1���r� �v������Y�W8�j^��1Le�+
�.��`�_�2��[�Ds�I�ܞh�2B�SF�x���`�R�P�<��}^O�n�r����ވ�C1����ܺ��^�bpȜ��a+A��'2�UU�q]��H[��?mI؟��A.�w�Gx�.�t��]���������6ɻ�|���]{2{͗>�$��4=:�R�o��u9��2z���i0�{7��8�)���7�ިǙ:�]��\��d�N;�T�$%wu^)����)g�hI󋂹qN�S�P�a늱�o�H`����@�x�������Ұ�hΥ3���i�ľ}p�;tek��|v����ʝ����_��"�"y�24�;�������އ���U��:+qG5t�?��;�M�Q�Sw���Q'��%�����b�2ap�y�Ż|���m������v�`4�$�z��5�&9���%Z�y.��e�N�Gn|�Χ��K�j��}�Li	E�A��7z�Y\��`4�m�Fbn��p�v��-�6��M�j�\�4	Գ0���:�������Җ�\�	�Z�u��9�6%�Tj��Ù\]������7�[��V�-��kx����CKdG.���ۛ�3h'%//4�V\!�Ԗ����xѼE��R��N_N�L��f�����~����^u�T� ���<^����|"۱|���E�hTmM\-Rl�φ��rT�����o �7��Vmo�z�Fm
suu�o-ڕ����v�m�v����cܝ�h��WSs#͹��î�c͐Ûc�5��ͦ>������:�,��Ր�[;b�H�4�O*:v^�=���6_v��<ɻ���4�h��KF�rpw@�J�i��N,/���'SF���Z��-�{�^`�/yl[ǲ���н��b��MZi��BTf�'W��v��Cj̖-讐(��1ݚ*ݵtg/�%�O�S�mݡj�C2C�����}��U��w�A]vNEC�nJK��bu�^�x[/����R%��h��v��d��M��U�ۧՌ�U.դ�:to^�p��J�]\��{/[>3&S�.� +n�2}��M"���,�Y�rWDz���|�Ԝ�7�)Ӻ鱇��V>ʆ:�{�����ɵ����j�Vh�:|k���+;��v�8�gg
&g&�X/<fQ�����qu�FQ��"�s�����d7�u|�{>��w���-f�z���[G�[�wգ늤�F�jm�m_uE�Rb�S3~��3��g-���j��r�Ҽ2�`���q8{���b=���Z�6x�َ�1�q)<�W�C)f�u;D���ia]aWXzsE�\����}�ph���b����n�c;��\s!��;�ԥ�ENμ7z�^.��Tˮ���9��ۘs�η�ӫ��,�\��[�n�:��B�6��pt U齅�����=gkI�8���&9�� �k�����g�1*���!Kjcu2h�(m��Tv�����M:�Ϟ8z��wIjl��ו�K(ʼ��,����ԝ�C:�s�ƴn�ۉ�t��A��<�it�� ��:Վ}C� ���a��ܦ��������tNout]0]��1�lV��޾���Y��[yNޝа�x�R��V멥D��J��T7�Ә���L@�n��CY�-�	���9jv�ޝ$����u����i�%*�<�D�5�E!�þ�>���!�枅i������- ��SA�p�|_N��R�Ӝ��y�l��6]	}�^�偉����_�[]u:�APS�y[d�B���Ҥ�wc�T�e��wD�ù�Z�Z�����K�'W*]1����L��B�Nf�d�/��!r{�b7�ɝ����EN���F9v{"��+���ĘO{k"qvm�yy2'}]��6����q����/��Ye��k��}04Ť��ls��;����!�x��pY�v�������hG�2��"��UC�[wD��&EDS��R���G#�5af<B�]Ͳ�*�ӕ@�9r&QE�$��dEV���_.NAv�L��$�+6p.��dQ�|w ���dr���rF�\ ��2".��[�H���N��Z˕D���.Yб�xYr�R�uZAv�Ȁ�O�9vPk��'q��w2.ȘP�TPR����bG�q�q�@�$�r�\��*�*�L"
(�PE����pH�BIʹ�	�3���BTkb@]�c���[�0��]�rc��JӅJ�4GM#�^d�R�$fn�<�u>D�������9!�*(�G*�!��;��~�����S�[�y ޭ�����o ��of���B���%��\��]r7��:Z�7�6�b{E)��b��Ck���'�0_W.֦�T�l�f�-+g5������t��Y�:�b�3�4��� �5���j%�ˀ�~�Ы乫e�w�0����ٌ�{ό���W�17��N�"P���Q��F赳ZX�.VC	����-����:y�����d�ʯG�Le��^�Tn��s��L��ѵM.�߆Bn�M���փ����V�����>�����=46�ї�nfV������s��;E�����+=�=����*��e�7�-�>��w��:� zK�=t���Hޅ�3||
='�\�r|0�l��~ڻ����T�G�Ǹ�WT{�M{�d7����Q������w�t�3�����
��ؓ�_��_wᾡrT��r���u0*��#�R�@Ϣ_��r���|���7ٕ\}�Q���&0&/37.3��o�>�v�f3*�>Y5��)�W��`-t�{�p=.��.}63Mg����[V���"��T���c��ۦhY)��7^�F��_�j���rB�Kޚ���P�
�"k�K�K�Y�ů7�=Q�I�f��]�����G�|�-z7+������_VS@�|��K�[����u�W��vZ��y���jn�q3k�L7N���}7�:�{0����뗍n��\�+
	�}ː��T�o�+����e���{6���C�A���/��Ag�(��}%�FUC�|��E�L�>�a�ϙf&Vb�k�f�v�Ԧϩ�|Ԗ}����;��m��p�qP$�xU�e����b��l��ټ���H�dК��~��)>/�G�O�^y\>���x�>�87�ug�8*/D3^�3����g=���g��-��7����[G|��^�TNO����r��F��^�U���wo�����F<�@~">�ȀX微��lg�z�;}�\MǷ�
��GWr�o����T��.?ԿR�gK\$zz���ؾT-�!����J'ԟ{�Ŝ-�O��p�j��'������{"m�W�n�Z6H�}G(�;W��?��T>N؛�U٫Pr�w�^d��I�%�`�#Ƽ �d3Z?e��Y阵2|��=6��[/�h�jw9,�%�����.�l�Fn�ǲwrn1��2}�H��uCoʎP�X=Np��+�Ӄ�:�P.�O�D�lg�[���pz��q��֫ˇ���hƿD�M��}���ێ�3f���9E?;�Y3�c�	���Bg�� �Q?].B��J��uI�J5M���4l����L#�h�u�Z�6���G@}x���K΢�T���副VN4,wTݣK�*_d�ͼ��a��q�@"[�`�ԩ�w{ŉ����Wtu@����[������_���t��L��/������>:NaC�r�ʼ�5�Gz_�o��eg���)_w������zB�9z�O�x�ۃ1�tǶ++�n"��;{L9~�cS�>n��5U���c�ox-�"׹�+�X������ۑ�t�ۃ0���w�Zn��*�m0B֬�v�yW�Y���|�E�=#�K��:���y�!�S�.�����,�-���gH~g�O����I��F��bW��0;�����x������y�q��/n1~�[%�$�S,*<�KnD�tW�:��k�Ĕy�1謐�mt�/ w��,���/�dW�ǖ9�GYXe�����5���;�-�sǅ��1qU-zs�A�����>��7>�Q��y�{���ǽ�gRG����CL�h[�(�� :HN����<�CfIA{���D��Oף�g���ʎ��X����=
{w�%�?_\{��e��1�n��=+�V	�Ƣ��*�5�r�E�.���^ɬz'���n�p�}�RMǷ�#��v��{�G�l�<���u���>�zc��YS1�ysNfE��r��T������`ʹY9�$u
��I��y��7�LYL�qϣj�����ٺqe��o"��P�+4��V7�c�4m�=�(���[Na��k�D��̺_W3}�V�c���/�"�����x�_n	OZ�#�?�n׎G�w��|vp��|�ߌ�:��Z��@�ԅfn�q=�UǳZ�[���z���=>[£������ȟ��;�|����Y�EĻ�I���&!�8�c�3�4��.��F����i�t���e鯣��C��ܘm�������b��B����S�;x�mu����z�|.c�������N}��e��Wx�^��x�A�߽> ���jpvL��j{��&��z3��1��ωT6c�bwL;�V���vX��r���3�+w�+j㢟�W���%�X��>��Þ��y��Ο� ��7wj�ey���7_�r~�vEH���NR�͚ބ�Q���T�����x�yUxR�wf����N�)�t����P}:�Ui���y�xU{R�M�z��Z'���@�Ԯ<���D�Wx����*�5�}�<�6&X�\�}�/��gǺ31�c=S�,]t�)�;>F�����x�ϥ�eK�Fo?_3�(������sq?yM]�׻Κ'P:/�,�$��HeX١�5�QY��VG�O�O�p�=��6BP�w�bZ&avV:����߬���h.�K}O!b�ѝNņw(��`O�k�[�x��LV�S�/���/C|��'U66A��^:��o�)��b*��t�8��c�/!k�=��m��XU���If��1�t�Z%��\�̑���Rq.�/GRJ�Όy�ۤr,�J�1�hʦ.*e#2|�ytq��X^�>���#MEmw^�{4�dN���m �Qf�D�Qc�I�wF[7�L��i���ȵ×��W��.O;]O�����=�{��q��6�=�g�]� '5��Cu����)�3�rodn�e:�W�>��Wp��E��+J���W�\���[3~�P>6��]}2g!t�1~�#�%>�f�� %��� �5�ޮ>u�l�zw���{I��Q;>���]Qgފ�����=���³wR8�o�@�ۚ�w�T���گ��ώ}��/<j6`�}�}5z`Ϳ��SJ��5�7�#��OY��}��7��j�X�B�d1p���6���ʙ߯�!2�S�9{��@��xe�N��f��i^��,�I�5��5}s��LWfˏV�����j�}���J����q�@sC{�u�nfz���};�b���5��׶���L�g)r�ɻ��~iݣ�����g���~���2f��zO�����E�g��d3��v����oQ���B�I�����q	h�{��S�+�7�-{���K}s��vvM���^i�}�0ͅ�V��S�8�<��wܯ�;kv�I�m%s����6�k�FA��+����m,�i{Z����Fssy_y��T��Cg�r��تk�c�R�Ͻ�^�������㓟��Um��}�_��5UkA�G��l�ۊ����>'o���*��#�R�@/վ/�Fo�^�4�o�I����d0oɄ�&��G�����c�QR,NӱN@��\R���2]y�Y�2��7$��c;�\J��گ���	��Q/@��Cu���C�L��N@j�T<|5�yF2gwB���o����p��5�t��Dz�����Ae�$�Q%�PeT;�>F�	�xx1��.�Ҳo'6κ�%�ޠ���I�����N}^u�m��%�	(�<�;&P>�������w��L~֦?}9O�G�P�_��#�O���'�Tg���Mg��8��������̲ c O�o_Nm���2|@=�1qS+ޜ��D�����S��<��W�\NϪ��3|u�8R=wt��x����?�@�=+�k>�[�����ͦ7��R�\��i����t	�x�Q�S�\M��h��"�|$W�����Y�C�;`�B�������wQ��H(��MpylǺ�a�Wg����I켹�q�WJ����P�iQ��'/Y�K��d�W��fٹХ8Օ3�Ce��e���Q���nי�4��v�¤�6�8�m���nX�c�,�x�s㌶r�wq;t✲u���U][s7xO,\�O���3��?z��g�&�Uz��%� ��FC㕱��/�(��Y�o"s���H�/Dy�R_�(xK k�5�?]x�Y�D�)��`�����
�ݩː�m��z��(<9�0��]ɸ�/���� o�T6�ʎ�6=NE7z�^ ��g�jng��5�����{>Ӫ���/]���9��w�~�qޡ�l��nWy����[��H�	�|Ǖ����^�^�'n6P�F��3�ydf�P^��}5�+5�W~ͿmI�˳zE{&�=�{2�g������wVW��9�v�i�&2���*�|	��w@��#�*��X�lO��t�����H���n]���s��u��(��2P���`��ײ2�s�F���ޮddK�����/=����Y8JL�4g��e<��31�7v����S�4�
�p5P��x����8������<͢��$�K	�H�}t��W�w�����l/EL�L\WH~�}5��0;�Y~9�K�Y�y�~��y��a^'���j3ծeZ��(�h��q���N�}/y���J�ɮq�X�$u����̰M����.�l����#-�gb��3�=���l��;i�g%b���]�:��2R҉��R��gv(��⩺ʓ�5.��'N����at��5,0��VgC��^���3� v�S�B�Zs��h:��{<4dyS�����;�s��ΏnxK���+�6a{�QF�Q'�g��R$TA��n�P^ϭ��"�?^��>�2��l.��[�9��Ѳ�;�	��W�G}�!:}��G���C"tf:��
=+�V|&[�e�oYܫ�=T��`]�W����O#��'���H��S�{�G�l�<���P =>t7܎{nG���V{wMsS�z}��G���|Nq����h7�z��Vx˙�,j�-M�B�@�ڪ���o#բq��s�~b�/N��}�P��G�!�~�q�O�>9��w��!��*=��.%�zIsѻ��}��+ڑ��t���|����5q���w��&����o�d�@�C�ϳ�\��y7u��e�s��@�̯Q�D�J������g���j�X�UV߹z�E��3�~���K���hΫ�	�2�U{ ;���~c*GK%T�}bwL;�V鿨�>�0wۗ��V��z����{y��>�>mP��Xsӏ�C��.E�O��<�̘}W?iRv�m��@\D�}OI���YE���>��b�n;��y�廻�u�X7�Muړed �ZF��p�4((lK�*���or5�;H흼i�U(wId󙙰����6^⻠9�3��ѕ��oQ|;��Vc_�U5��Lq����&���2|�ZK�!k�#�[>42������n\T���N7^��g»۷���['s�:������t>���c���=�ZgVx\��)�>��O�@�Z�Ǳ��� �N�����B���*xtC�:vVoi�ox
h��2�6Ź����A,���2���X\�w���.�+>�������^���髥�Z�w*��(вR����$��rV6hyg�]�Y�xR�z����B�T��p�W^���kx��ʯI�c�ѕL\T�Fd�&�0�|���{TL�N���o{j���.��h�Y��C�C���8�i�r�6�$�c�)��e�$��q6�P��Y�+l����Mua�D��]kNBr|��u�7�TF��^_q�%� Nz$�����gH�yxqe�?_y�fAL�U�Wq�9��\wޓ�_��#n+�lϽ2�C�w��]����^�
�NI��
;���*��ޮ!׭��޿3���'��D�DW��d\f�D-6�u�|2��M��>u$5	�>�4.)�x�@>	oQ�m_����ώzg|Kf�\����mh�IoE���ʀ~��zD���5�j�m�������f��y B���ENt��{�bw�osKrޤ��[��\����r�r��f�۠�k%]qʷ�����Ά��(��Ն�_��(ѐ;���t�*�㵛�O.�p�y<�����&�L��p'��K�����\F���+!�M]�һ�7'�v�e����x����e�����=�u!{/�n��o��QR��L��ѵO�˩�����ò&��M{�iUɼ~�=7��~�����w�.y�LʁA�l9��2����tN�\�ԍYѸ}�yp��������n#=t��?]^�s5�>9>�wzOzޫ�W��W��z�J��^����Ʒ/�*��ϛ�R���UxR�/���Ӿ3�d���=�^����9T�vqx��Mzg����ꜣ��K'WK���#�R�@ȗ����hoS��hӓ3Xm0�?������-ۯgIݳ0�O�X�3�~� yX�`R�hq+��;�����&@uPiY��<'ԮW��X7�}�ԅ��#�g	J���L<�U#t��fG�}�7/
�p
�����o����v�'5�~�<��hx,u���ʠ�\�J5%�_U�ϑҖd�eK��V�bQ7�{�U�q�3���{{���r=��g�|9:�A��]Ô	*���};�zV�+8יݱ ���ȓ�+s���)Ky\3�^����-d7b]��!�l)��mW>w���9]
N��7_oQ�����U�]��0�� �}G���u �$g��V^�q����P&�,�4լ��շ��s3���5L���/�wMu��
=y�k��`ո5� =˙��IF��zT���,`\�R���M�K��&�[�O�ךe���`��H�@���`�ЕDM�C6f�-&����Ua�ygSfG���$�VG���[�}4��5�؊E��*T�pK��ବ��C}g8s4�z���,��S��u:y���ܽz�^�Q����|�r��I�7M��CƆ��J9�&j˫ug>��C0�:�J�U�)P�<��]��J��iK�w7V�7�}��nIۡ�n�h��e��;�[�g6k:G8���}���V��mߖ��,(n�M�g<�[j+��{�����J���u��P��O���f8�6���>�(����nE��B5R���l�.¤��唲K��]�\��O�S���D's��Px9��X�@	���&b�9wͺ�7�eY�]�{�6��2��n�vw���k�黑��3��{����83l�@�����/���plZ�����1��!�xzؕԬ��2[�u/W���zU��Mԋ)�(��)�z�m�{��G봰q����4D��N/�^-���X_.4�*���q�}b��wEk۫_wQ��V���ζL5ǻ�rp%�ժg6��mY���N2����Wd�ݲ������S��.��K
a�o�����4Ԙ{f)I�[��8C�S �oeld�]�*�u�К��]'M�'�$�)�W��^wuuŽC8t�8nغ`M�C��*vɽ}����$~�x�~��Q�7[!�\�]1���\46^>Z��s���/��-�k-��塔�^V���t��²3��Я&Z��.&E�fmd�	���G�ʑ��V&��"0O]2���v�+���,
ܽ$�#���p�n���vgާϋu�o�Z�x���v�*�ij���z�����
ߜ:$�M {�m*-bu��e�u���a�fK=ѝ��ː�%J��nǏ�0�Yh�D�U䆹R��%J��M�<�G�S7�K�A��W����a\.c�<�gCՊ���1.6��u������titor��=N�9�s4�M ��0�l����݄�ל
����Lxk�w���s:n��]�pu���'y�mWw*w�{ݶ�b�� �#���'^�\=}A<���b���T�A�'3A�S9<��<v*�x���IdV��v�
2m��b�4��uj�;��)`Ô��3���,Xɏ�J}�p٘����\q�q�L�hR͕����K�Օ�n��-�\�f�Yj�W�s��q�9����1��y�{֞ۥ��4	 �ps��ri�.P\�w�<��"x�=B=��%L�^az	7$�"2J*�UM�
�p�6Qǎ!�/T��(�$\�X�ǎag.k�T�d�
(���19Dw3���+3�G�EUE��wq
���^t��L��]���A�q
9�9bȠ�!У�r��9\�.���2N'.�H"(GX�[(�=�C�,B
ri]�_!�r����
�*�g+J���Q-��v ��9�8�Ay��'@�t\ȉ�W�9�VE"��&t�1Ҵ����㞖���PЦ�&�<�'V:��:���;��I�
��'��rԒ�J�=�rXUӉ!�Oq��2u��*㓄ᜢV����Fr�=�\�`-p"tδ��[�ӎ>���&�|�iY���eZ$Zi����<��e�ws�c�f���V����W4���o�����*�����L.�^����#�'ǯ<�x���q���}��j��=�lN� ��e#�A���J~�JpKt�����yIү���͜�^�=����r:����fy3�r����A�^SX����G���Ͻ;���1����qQ+�7a��w~�'���'�ӿ\M˚,�" 5_	��z���|}�&[�Cx>�W���>�v�szV���h�L�dxΏq�z��g�&��W�P$�x����F�㴲غꦽ=F_q�����=�Ga�v����I^���� ;�ցP���n��~J��?�]��x�ؘ��5^3���Zݍ���h�i���eC��ܜe��*=�P�s#6<����`�9��a�{��iuFO�����O�8�a�*^�Kk®6^��yp����c5�+�o�l���]��DZ��[{g�����^g��]}&�������I�({�7.�1�}��~��7Tu�k�u��2�<��˼3��H���r�G�yo�wL;��q�s���0�_��V!�#&����M�cF��ec��C���;D�ʃSq�}t���e�bԖ�]'𽟯��1F��B����\lP����<�b��r����ԚQ��7s;p��� ���7�곚�w��L�vT�Z�3^�.}M�yYx�zUI3�^e�e����nv��Vs&�E�d߰G�%��ޕ�E��ۑ�03n�϶[���p�I��׌e��a�.7rԗ�����<���r�/�.�7�v=�>��C|�(�8Jq2��ꅷ��G��ߧضf]�5܌���}��p��P��������y�Wؽ����u�P�RIOr\FM�D���]o���	�
�gT�Ґ��3���T
��Y~>�~=>U��⻶��{K�]��S��]�#8}�� �x#�T�Bd�9�MV���#�z�܏u�>�͙�W �mE�U��]�	��[�=��(��(���,��ٺ�A{"��.?^��,\�.�}��B��o{p�{�t�l�8{޿\{#�Q�d@N��@��x����� v�{<�]�Tه
�/"y��Þ��X�9��=��!�߷�#����~�Q�� ����Ku;��+��z��������	�Ɩ�v߭��zgx��c�ՠ�{޾�՞3:�����KR�o��&:}@��#Uw�����W�T�x��xT;m_��{��O�zg|O��k@��z�ďF򛎩���+l���Q)��m�g���ee<�f�<�}�r����.V<"�??T���H[[j����u(֮���Q)^�fd���gvN�+Z+�m���,&�r4�<+9f�+��5�t�eq�
��e�P4�� ݝk,0r��+g6+��}(.�sS�;RzZ}�}�o�O��GM�xП�N6^����URa��2S.��2Gz�ƫ�N���@ײk���n��){)QY��=�*%��N}���7UU�7���=�ǿ1w�u6��Ef1��B�¦}�R�={���<�T
��*�l��;�׫t��E��g�Lh����/t�l��9>�I-�>���U4u�G����Xs��do�eȷ�t���py��P�"���*Ԣ��2�s�ib����J�(�>�w+�áUW�����^>S>��wf�����;�t;q2�4���z;}Ǝv�5�q��m���u\n�D�ge��[�q�x�S�3����y�#{�ݩ�Lg\�ʇ��}1�Wt(ksZ���^�ѕ�c�T�NG��,�5�
��k�K�ʗ��˪��=&��W��<���1�Զ圳��f|2��,]L��!�cf��|5�QY��U��Hm
g2,-��דL*+���=5�ſ=���(���y2��%#2|WRY�Nҟz*J~�ڛ ���w�q֦���4%��{��u��Ǹ㭤q�,�4�ɞ�[�����=yZ�
��a�����Y�l�]V_>�Y]�;ۧ�:�ۺ�8���r;y�fK��G.��;s�qh.q��ލ�9s� ��w1�3�/H�_u8vΥ'G��k��݇�xE��>��Rmc9��=e����O.�YVP�����6�7�edZ��g	����F]�+�{;���#贶�o�N��<���g����*#n=�g�]�� ���x������ԗ�7��r;�����n(�Zn"���\�H�3�+�ǽ'J���g}^�fn=�|N��٧��󧑔�u�ߢdO�� ��B�Ɩ�py�m�ȏN�����i7�z�{��S�����.�R�:���#�.��u$5�yM�s�;��*��d6�x1���9���G��|+Ü:�w>�%{ƣ`W��z�K3�(�A�0��z���j��c˕����V�O����k�fM�B^�O����n4
�xe�����&�F�=�/�t�Q~;Y����>>��oUͮ�F��ٻ�ᐛ��c�����q�|�ێ�e�󛙕��|l��l_�������û�y�x}E#�s��_n^\<�^�G>���o=t��?]���d��O�F�ˌ����i�i|�B3<�C��O�8��{��Co�i:n4��r��⩯q�o�K�#�uW�,�~�ӞpK��盛��)Vmm�7��Ӟ�3����gng�W�gC����Q�9�X
��#�S�@/վ<ET?g*b��fvt��ո�B�AF���6��X@�XWf1�wus�3i���\�S]�9/�LasW��ɰ9����7E�M0�)�F����o���-+U��+u��᷉^gs��ZR��F�R��C�m�Q�%��n����:d���Y5���n�J���G��1{�ۮ8Γ�fa�	�,\VMi�� y\�|��Ko�������,���y��W���~�B��n��8J@ó�z��Ez�������N�ׯ��uW*��M��\�ߐ���B�Kޚ߯�ǟ�����-~{t\�J5Z5UC����zmb�4�4�y#�9q��U0�>���I�����NEyׂ�u��ϸ���INs�������aw[��聞�눩��*W��"R�~��'������<�dzk<}�h�q�V�q]��y�yg����n�s2��-��.]!���[G~�A�������}���D�}N�L?��8 'Pd����yMd�T-����W����Kӷ�i���!�����R�o���q���ܹ�͢ 5�^��t_n	��6=X�_����Te'�nǾ�j�<}(�?��n=�WO��:��M�2KD /�W�ת����yݹ�j�L�z!�{�.B�ɪ�����@�#Ƽ �dC5�S�_���Vz�-L�)qB6�ҵ�m��~�Na$Giև�,WHMa�-B�n+��$%j����&x�I�[u�([�Ѽ�Q�qL�f�_M�ӗ�6�Q˔���|��t7Y=�tc��uom�k�\W�����D뵹/t�p�bY����})fɷϟ7R1\CGfm.�v�y�vu?�~S��ʵ�v�Ɨ����wro�'��_T6�<����r�Lye����؞F���O�ς�Ӄ�R�迩�xU���֫ˇ��v�f�EzM��@�����c�-�-P����M=��JE���gĪ��WkCv�a�����b���7����҃y/��ǳd�V�����.�Д�2��u�z'0�1;��Y^�t�Aۍ� ��r�0.�|c��̚�ie��DuS�"�/N}ޚ�;����ۑ��9�f>U�*��[��c��S۞���rS�D ��Jȹ^����J�{k�ϼ���9�*����/v�%>�~ˊ���V�^�c�9z2\Ο}G�y;.���I���;���y�q�������s�k�bՉ��Κ���Y�l��/�#�L���򘿫���|Z��ިd��}��W�ǔ!=�B��.ixn�ip�U�t}�^�G-I�@�,uJ�&O��fC���0{�z���~+}Rb�y]�Y4��M�.�Mo�{8�m�I`��)*��u2��[y�Eu�_zY�eW #?�S�գ��gG�rk�n��q�Uf���U��6WǶb�^׶ܣ]nRڏM>s6���śCpS�ﷅ�X�>:��gCOة��չ�e�IH�W`�\���5������!	�idҸ<[דL�yjݳ̀Of�sj��w3O.U��Ǿk����*:UǶ��7�������l�	ј�����Wgύ�C���+ϒ�C��ܮ*�5�c��#��RMǷ�#��v��{�G�p��j	ns=�^�������st��s=� �:�L.+xL>�o��ȏL�x匿A���|����nUIc��{� A��)b����-Ϣ	���*��Ѹ�[¡�ͫ��x���q��ր���V��f(k��mMy�#��&���Q�C'��4.�+M\l�5��!�ɫ�16�fK�ny�p��>��8���U^����F�D?P�'��+�y\	�1Q-m��s�5{,n��:q�`bW�M{��f�7�iP����> �ǞEi����<��5�nL]�����'a�T��$T7��P���p�~�#�������C�n3�a�N|�4:��rFg�>'j��F���uT��y�1�(��S�7z��'�^�w͗J�{��� �7t�/�ʫ{�4\G���w�:v#��O}[ӗ�̪� w�����qYU���ģgg�)o�ǳ�3� \Ju���m�,�F~�����}&���R��P�Pe��Q3�D}.r�ff�0��N�ׯ��p�L�nc��� �;׌�I��r�TCyI�:��F�Q���x��_pw.����Vh����>���ֲ�ww*� �Lt%˽��0�{�DmZr��q�Q��ʽ�Z;�
���	Þ���O�S�:.��)���\w�����L����T�k#r�-ŉ���Ai]�Fw��F/���J\e����ē�v)�e\�Y��p|z(	'��;/}�p�mدG�/��Cə�c���x��P
�3F�ʦ."�R7U>	�8�W��>����]I.�hP^	;��x��Q����qs���rYl�K���@��P���W�N������|�y�p>9��Mç~Ӟr|��G���*#n=�dq�%� Njt�~���֣^�kb�8{��:]�D�2����n��s�3�+���t����l�i��{�Qq����l���� Y�8��@�u�~�+>�[����u�l�Dzw���x�2��6��&6s=����QF���y�H���P3�������!%��hC��ϯsE>���9Bx�����3��g�F��{=q7���ID���/��n�[5{,z�ٚ=Y��W�-yJ�ǜ���mT�Bn�O����b� �xe��^���dy��TUR���?��&����w���X�����!����Op�|�o�PKh���Ժ�N� �]v�"hWe�	�#��xA�E���Nא%ם�\1Y����\�х��w)SU*v�ח+2�\��m�q	������8�Esԙ�4��Uc��Uuy{�m[ir�Z5^�Q�=�)��ԗ�����z�C23~�F\
�<�&eX6������jb�˺fRQ���ᐰ�>�>�_n^\<�^�G>���n#=t���Hވ^��7�8w7���+xTĨ�'{�v��Na���6��n~|���
�~%��\5&}�9�E/�=�^�߾�l�Nn�zM{'��g��:��c��Ι�Q�C�rplR���`t^�dxd:��kpMV����EY�t���9�L���9���^���n��3��� O�b�kM�9�����������(�l���r�����+Ճx���H^���4,���0���g��z���y��Y"��w���24o�����MW���<|�-����Yr�(��Z;���<2�$��z�Vm���u��E�7ze��|;��>�|}���\?)�9����y�p��q�ӿQ݆<�g豾��`�?%����g�j_�.�ԙ�y4&�Z��9�'����I���+��S�R����q��jJ�ɕ��8
7� /�_�J�71qS)�rۭp��2�[D�ܟwQ����u|:�� ���(�n<���.8�;'+~�6��l-<^>$��}�S�w��7:�K���kT��H��b�8���,�뭠Y�H�^���d�L˫�q���n˽�d���m◼����X	���v�ܤ�)Ց��G��LإQ���"�@��W�G}�z�v�ݳ#�(�� '�@��/�Ҽ��:���x,@
�z�P
�0P�������xm��V�k�.'����^�\M˚,�ȈP�8��9�Q|}�N�7 /I�'<.Ӵ����я���O������>�8<OG���.}�ț�U^��FIh�g
cMB�T���boal��H�:2�mG�W!1�M_�߽�@�<k��3Z�ׁs7�����y37S+-���z��e��C�-֊��~;F��5�ۇ���7�9~&Mǽ�������X���s=�V¹]�#��z�9�c���i�S��/�����/]���5Y�Hv��ۗ���2�M{ N�R3��0͛��T2a������>Ӣ��;{(z�r�
�F}���#��[�v��q�5Azs��׌��\P���.Y�>'t�a�e{��S�z�1�W�E]-�����=�� �n��ϕW���n��9ޚ�;J�_��ۑ��9�f>U=�c��ޟv����Ey��Q�'�m |��"�z��.|3�+����>�7�r�_\�(m};�O�+��aV~�/wA�N�U6�7�`ʕ8��e:̂�[�O4Ҁ]�/!��čj؝�w��;]vs9����&U���9t��m�ؙ����8���\�oϨ+;s�"�;�ǫ]c�o�}ܸ�=�y(��77Eݳ�*K�H�X��yWR�7&�(�d�˲�h�p�.��N���|��Ytx��U͒[�QKZn��k"�h3��m1ƢBf�V�b$b|)�V$�]��nK�p�p��ڗ���{��n�k�+v4I���������so���h� �c��I�38��pNA��s9GC͛�Dǔ����c��P�ǥ�L�1�j�+���:lS�Ò�Е{n�=�_],����?�޹]��v�TSۤ��[a��];{�w�D�R��mM}�f\������7�vݭo���AV�� ��l_����t/���6�[�8R.�����sIuiw!���x#�F�ΜVmd�V���`޺ᨸ.�CU����᮷p�ھ��\xnI=L�X"�QLI����=�&�X˫�� �3o���x������1}��+�m^̫��亾����S��Zp|&�(qr�+mYDc��m���4+@���M�xR�6jUh*d�c/n��YV~�d��Ϲ�P�R6��+�k����q�p.�D5�1���Č��b��u�V��5�о���Ό��Vn]�tm��ZM1Y˯{����3�q�@�oi��`���Ujήh\�[�9
��2�\��$����>����)u2�M2��g1��k478�WU��Q�tF�ӹ�"�k�^\���Ӷo#|U�&7j,f;xE��F�#�2�\`��un4�d�!����Zh���D���=�uc-������K9"��2�{y2�Q�w�*���֚��G�����0M�,����m�͵Z���.>Ș�	����*���g��� MJ��8u�R]C�!��zw�P�J��m�y�^��Q�n��@�6��.�9����4�\���ԗ�o��"�V;֬7͞�̨�Ԯ˼�*�!
.-C�d�)�-�����+�٢k��zs������^��y	!�ŵ��j]�Ц{��p��F5�ܛ����a�*
�귔��uL��Qcnh5�	 �ڷ4)x�ʹء��y�^,ŷ��w��}�͌t5��Qb��:�Ft�u����8r��Z!��u���T�J,���u9M��5��7��=ѣ�c�ywu�'lB�w�M9�2]:��3]�^Ks�#��n<�Vƕ��WSc{i��Ak����v��kſv(�(�d�8��|���ͼ�iVa�E	��I���drj��T��
�&�9�&ʾ��pl8���E0Ղ��WWk;��1�T����M'���/.A�����J�@ǑA�L��*��!2l�U�a��* ����-:�h5���yֳ��a���q�����賻�����,�[+��K˚�l����;��IQ��( �}��L�u��E9�b�M8����Es�{��Aw�E1D.Ny�t�9E�넇C�%ʩ�:��xTEP�Nr�0𓸩�iHsA�<���r�[���gq��廻���ww�C��KG:T��g�`^Dj([��r��Rs�,���9G�s�D'x��<a	\��җ"�r�̇:�nyW�\�׋]㻮�gu8�B�M��������ȲHH�<�i7eyh��k�y���s��vAj{��Vy��i4�/7e�&��Q�N���W���s�)�#֒�q0�,�X����˔���u,%�iqW"�/]Ź��uݧs�N$��T�
��[��%vh�-oNMȋR���J�x��L"L�ft9�Y�4t��n�J�0��[^E�Z�>VV���V�o39F�aY[�Psb�&�v���v����Nu8�M�ޕ���-�� l���:�k�����e��3�����{�8�*�e�8�(u�zϠ+�����'K�ձ~�~/=j�{�+w��Z	�S�Ol�ʳ����rIu(*�3��S>S�'7��^@�T
{E���K�P��;<sӣ�E����]'	�=5�ߺV���RAU�~ȱu*��>NzMV���V��0wRUw�?cHh�X��Q��C�|��=��(�2�.�� �H���l�T���x(�ӧK���%Շ�$t�V'��V�Qү�HN������9G��d@N��1�&t)�8�ё�}4�ϵ�$kɛ�@����+�5�d9��=��!��}27��lO�2}<��Z���{�,jx�ƕ�}��@��x&=ơo
�ߩ��3�}㾞���_ }7�2�E�kM��
��Z+\�w�����R[���:G�!W/����{�*�j�&���ȟ�����O9�f�x��rA)'�J}w�)�H�D��I�2G���R�h]zV�������C�M]ɇW������>��,�2}���ꍊ�� T/ez��sW{TK[z%�a���6�����`���=+��ΗVF5s�_B*�١n�Kl��7v��T�1��YySGp�F�����72bzY��L��ְ��j����r�d\���zK0����\��u����(�z%����(��r���,]����{k�N'J�3(FA�ג�.����Kt�Ə4��c�3�֮'��T
��*��>��a�z�O�1��|�&��<Ȝ�~IW���2��r�h���C�o��Xsӟ?M�����>'j��A����F�pݫ���q^�u�d='���n_[���9ׂ�������q�ml�����[�{Л��X����9��·qYU��&J4r\
��wϝM/��(�����y>&nvz&��s�Ok<�9��~�4Yx��A(9Ȱ����Y�k�+���%�^0+��˔oTu�;�����Q^�}q��w�ǹ�J*����2��,]L��!�p6hy8RX}Q0\�^ĭ˨r��ԦϠD>ҭ��~��҇�9�F-��׎YD�Fc��TĒ���v��^+ݳ5߿U+ʺ�������,�s�X���s��=����.rPk�.N+���2g�N2��ٯ}��~��ϸ�T����K�^��r|��D{����߇���.������.�z�%nn� �@J�T>�2���z�o�N�9g|W����W�\�_P=���a𨵽��Y�sp*:�o,�;"����37���,�2g(Q���
�vJv20=��~5��+Y�<ۘ�����oa������z���й�N/�t.X45�+�u�egK7q�pE]��F�{����I�,�O�C�C+`����SwGe$����k���E�Xn�@��B�|V��jz�1�zw�̚�����k){�y��u��}����u^26"]QeI!��H1 �)�t�w P���S�_�w�6I�wot�ɢ�h��[����/"<j6{�뉿�Mz�!�=F��E����)3��=_]a�5��h�Fv�	��ۯ���b� �xe���Q�FG�s��K�F�g��J1N�X�=2;�W�6��j{o�uro�M���>σ�qތ�ss2��G�2q����R��zÝl�D��98�N�M�Z}ǃ�ۗ�#�������o=t���Hه�[^�^� ՛xo4����L�Ӡ�0�-����Y^qR��7���Q�}p��S^��)x�랝Ь�R���*�n�����_i�����t����DL�
�·u9GE�)�Nު`W׾Y�S1]fnEsKf���^"V8���9�M�׾1q�ݺ����a�@�"��Mi�r�cLT�([̉^}��H]������_K�?KدV��ԅ��#�g	J���L5�>�|0Dz�5 ��0�׏<г���r�\�y���Ԃ�ǁIh�7box��2�.kZr>���3l�/�5}w-5,L�siͱK.��o U�\TY�ԅ�; �.�ȡo9�!U}�wd�%�x5t�i5��ZB�6��w�3���/r?��@�2\7�-t�魿S~�CÔ:�B�~{t\�J>� Ww������g�R.��Ϫ��n���nU0�w��r#�'�ۑ�~S��^	�R�	O��q��w�+Ý_�7�s���g���=�2�����9&���U��<���9���SP���c{�
]V�	��Y����|o���0�j�s�L���n�M�v���F��U3�C^��oc�}�Iҽ�����l����p���� �zW��@,q�R��\'�7ױ>�0�{ԝ�x�W����O����7����K�,� 5W���ps��W�Tsk����ڔ�f�v�oa7�L?�>�O�<gG����\��=�7��(Z*�Ǧn:gʲw|O���#�MG��-��7G��\mB�\�C���M�ޤ�<k��C5�S�_������@v����o�U1�s'�l�ب�բ�*_�����w���n�N2�L��z��|�O��L�W+s�&��<�N�QՁӜ�s�t������
[/Mj�������Ϡ��t�G$��o_��IJ���;��-��3�FW�S�5����� �x�>J�tU2��kJ���X7
��	���Z�wk�v�,�/���ܹ���Ӑ��Ɠ��c�o0f]�bR�b��ܢ�\�ڹ2R`7��N�қ�Ͷ,��KP��T�r�z��}�f���Ī��_�kC����Nt���=�{�<���Ǝc��a�t��>�cѾ��25�����k�VG�⇽wR�������cʠN�VW�����ݐ��7�~iQ���W '/��1Uz����ӑޚ�;�Eǻv�k8N`0��yZ�j�����F.CW�%���Q�%\� )kVEįR�����)߽�<�н󭢭F��� nY�[�no����^��5]G�L��Qp<��v}_�]Q	:^>�����s�Q����$���$k����ԫd�����&|	�I�Br��׋�ިd��l���Yx�;f�+=�&���E7p�zkQ�}+M3�����<��_Wk�yO��X�����8�x/2�]��Sg��A׆纏�_��=���=��(�p�$��<��"�>�ȿn����g��2��կh��K4HR�X<�|�z<��WG���7�_�=����̈	ј�޳������L��v{�����z��0���u�_��C�y؏z��n=��q^�bn=�����2���ll�P���O�a��æ�#T��6�zL<�M�=ڴ�AU�n��-��	]��w.�-ѭ9��y�c��Y�gd�z��7c����dXY�{�"�X�q�v�'���~ym�:���ם�*Y��l����_Y�*�f�b�F��lv����1'�W��q� �/�H�Qn�W����L>4��C����|Nq����h6���3��޹��]g��i]�Y�|�N�u%��@�ԅ]K�p�KxT;���O�|��8�ߍ��i��lz��ϻILN���<H��]פ�)���b��xП���;���nߝm<}�R���>�{�G�&5FO��}��Q�]�@�^���.c�Y��koFE9����n7�T\�+{ˡȟf]����,~��n=���#�"��y�>%T�}tï��z�V����û�g7�Gq��S+�����3�+_�x��g�Þ����{�#3��5�s�/k�N�H�|w��z"���7���WS
���ׂ��*�
Y�����I7^W�֤���r��w���t��3�!b��M��Q���R�;�d:�^ d�Wx����lǠU����.+}�ʩ\�ޏ;�m�Mڃ~�E�O�hJG�,/�.-x��ճ�9��9櫶��xY���.��ϫ޸����b��nQ�8JVe��g�O�ا!��dz�{:�F_�gLO1Oר���������V��к͝j��į�+"�]�nf_]	b�S�X�8:��o*�/=�{��Vs���~����{���W]\�ĶJ���g)��R��鑾�={M�˳O:k(1O�	��(�b热�yt�;�,X�����ԝ�?p�����6}~�K��^�<��F9��׎YD�y2���F��r�?W��r��g�>��p.ϖ]w�V��>��t��Q�[�:�A��Ͳ�/��i�<Ʀ��R��q]jGР{㞨������9m���Ν�Ny���u�7�TF߽w����\1���m��G�'c��7� rG���l�Q���w�q6��G!�����������D���Q�[����)SXg��U��Y o@n�W����Y �+zx4��ىj�<�����~zޡ���>�3�K��'z�w�"�]QeI!�L@+�h\S��܀|TO�GH8���.jϔewj[���n���O��������Q�=��D�3�*�\	�0_O���lp�<��z0ݔ��5^�SH���\��/��܋��^'�3�;��h��2�T/e���2<�}���y�>����s�w�p��gj���]���\��~�=7��~��9��ތ���ۂT�	#�^��I\�L�@����]:�7E���/MF������r#_�I��]1=��_
�x�$�n��GeaKn��� F���z
J�
^}t[��Vqz[HBA=Ӫgd��&�G
��tc��k������,7̖�"C${C���ys�E~�5��_&@�|����L���NЗ%o���e����5����u�YO"y�R}��`���1�]ß��������ۊ���мy�L�mWZ���R��K�(������c=�1���T�,�߯��~�;�:r�vv��c:�,�w���u�~�O"��/"}�=W�]�6{ѣ��\�}�}��47���_�v�3����fT	�,_ՓZK�j��;W���ows������Qڭ
���Q.��.}63O?u!�yT��8JVf�\�5래��w|sv�c�^��:�7] y\�,�����k��MW��/Upc��p��۠�un�m�&����K�����w��Z� |��2�e�v^��ǵ	��R�hM�d2�t��"�����^�������Q3�L@�w2���O�3�恥���R|_*�N�Cِrp�N��SH;��w��Mg��#��,�8 'Fx	�)@���.�S��Z'���=5��7�7o�a��=s�#�Rt�o�':"�v�?������A�:`�zW��;��y���j��뺐�^:��y����<3�^vǎuxj�z�~�\O�z�w�sE��D�H3�^޿{p~��\n���N�S��9ŗp��枖��
�,�&�>�F�6��x� ZA��&Ĕ��koa��vF2�z�v�[79��}-��v��r�.��TZ��uf+��gu_F��fVsֆYV��wN�e�۷��[w'p�[��}�cwg��/+pI�bj��R~���/�n	��!oa7�Lx��_����n=�Wq>�dMê�T�5tFw8�;Z����i-�}�}�N��c&�ʇ�Q�
�Bj�'���|�k���+�	ߟ,!��z:��Uް|��1�JSǦ�K��W�K��:��m�ϡ*�q��d��b2���f�绌��`jp=T6����	�S����(�c�+N�{>�/N����D!�Λ�$���o�kԳEe��j+�}��'z���w�a�7|J�0�d�}S�:.��;�P�S�q;�xk�^��4�>X��O�n�hī�#5�����k�VD{�(T{ٗ,��c�b�~��d����� �;�]q�9��_y��Փ���� LF[���T����ӝ��S�J�_�v�nC�'wv/Ž{��z���}��v�n+*��Q��V6� ���d_ҽK�dK���=�"<�����_�-:�����\����@p�X�uW�7�����1Pܩ32�=�Ϊ@��o4��]���!�s�PQjI*�e�P&x;��򘿩�NnMx���[���e����r�t�;*}%v\J�"���]�'�7�P��女I�Skc�\X#r��S%*"���nO�'�$)ňwY9����p ��?u�=��]�92��1[fs3��)T�ضA>nV��˩nV�&Q>��(|������X���pݟ�r�VDW�ǖC��_��QjH(�c�U!uS���+��{ѕ���mʮK���R�0z�7#�Gǯ�w���o�{#�Q�Ɓ�Bw�9��f���]�
r��/w���>G�T���h����w�W�[Tt�����޿\{#�Q�D�\���`�������+���uǣ��y�|io���X�9>G}�᤼s#}^�b{}���zAO}:�*�"���)�$q���P(��>�-�P�>o����������������Z���u���m�~@z]_��z���B�?��O�����|tl�з�CmW��}}�ߥ�CV��V��gY>�����<H��u�(���uX,��	�Xk�МT0�5c}�0�M�[��_�ˮ�Ŧ�fM�O�w���6+�B��>��\Ǖ��0Z��S��P���so,��'�o�*�*5�Fz#z��w"�����z|��ȭ7�2�Tt��P6a�)���b���Xcږ#U�G���Emn����ί�t��*�#��C�o��XsӐ�4:�<�rFtDY�~6�>��	´��ó�7T�!	v��Wq	m��I��I��O9�M����7��L�W��V�z��
�)v��q��Me�;��gB�m8R��r4T5�g+{^�\�F�:����}w��`�<ͺ/w:P,��w/��b�&E�	Z��#�;&vV�\�:�c`�v<��g>���d��@t�M�,ݼIn0�9�����b�u�o_i�ѷ�9���_G4"�C�H��YQ@[������}͊�=�V����]����jV9ɡfER�P͜�uֶ�,țǘ�}N�q�f�qѲs�*�h����fY��wd���$���� ��)Nj�ͧ8��y5�A{��H��I�OZ)=wpM�׳,:��1�6��n�֛�P։79u�
,�C�e�:��kbh,�\��b׏2���ɢ�9��Z�3�����ev]c���8���վ����7ے�h87����9��<�`c+�渍kDͬ�M+�8{3��;����{�u��[��.t��V�c�T��趝[������j��2f�g�[�W���
?J�#�����SN�[{]g
���e,=�ns��W�����-c뼓d��Y;��{)�.C��޷r�6Ly+Z���:n'���v+$}5��XB ��"]�����w1ɬ�Co]"y�����\�n҅���V�N�%8z3xG={�r��H\�t��
�Z��Lq�0=`�4C‼�B��k7�(�#\���F��t�l��a-���ulza���oF�:+���HR���Z���n��� w�00��c�zk ��i7F�9yƻ��"i��)��+<����[ʥ��|�u$6F��mvN|���us���͊�9X�0�iK��v�a3��G���6&Ea���*��ၪk��4�]��\3;�)CG&v���[��Τ&O����Ӭ��
Oh`�`z�]Q��s�G��l��m��Yw���X�r��y�5��eG��u"w�T�@�_b�j�Q9�䁽�=[նO ��9�����H�J��s�uԟ>�4d�rӵ�w2��!����7�mn���s�29C�����$b��͞Ù���h;��K�ۦ�����HX���w&���b�.�<��[\�^�4Z530SƳ��{OEՕέG2��NX�f�L��]1Wӟ)�{���]w[:!��Jѯ�<�l�R븹���3�������������w{���/)0��zeӡ��C��9�f�[���[���4���V��=�X�TX%e:�z��9p��)�v�}�(5&�nи�,����������M3xѳWQ�Ӏ������v��b�M����7ƛ�a���$�Ͼ�lDj.�X;]��]��Ӊ�Kx�t�B7P�p��n��Y�z���F�=}��{�sV��ֹ*�Eĭ]H�3D�K��/�����l���U9D)l���(�:�s�<ss*e�0�����ē�<�r�y�С�<�T���=��vVVLO+�����ֲ�':Gq9	�gs31��������Ȣ�*�Չw��x��T]y%N�\n�yҪKR�r*S@�)2�"�r̅Jo	��:�
�N�HQ$�V�N��[���U:q(�� ��X�)K�KTΕ�����J�P���	;�6mSy�o�M�]UJ#"!5e��%dkNIФ�e�P���v�3YY�0�>q�rC>:��hUd�-�<���Y�@�+�_�*�*�Q8���t�K�TH(��ec-�Y��G�s���j�ԡB��ė����CBT�I�43T$D��PxÔU����,+z�矞=׻���&oS5(,SOb��£s�7	\�]�=��u��H���m:�#mm�T����}7_�sr+|�#z�4շ�%�>�s��n�C���#t}����w+���UT���ü_�W�'^T�wmq�#~溍,��XՓ�sЧAӷ��`�t;�ʮ7W�F�������ix���+z��,�ȩ� �]Y~��L���or�o߽��S���ך,�K�h�;m~��YR0�:�6�����A���6}���T�=�~��~�f���9p���_<X���"w"dL���M��~R�4���5\ ����J=�~++ԇ�3���ʯDYD�ye�v�l���(d����7|5����-ґ��߽�H�^�p�x�G���_�l{�C���ϯ�j|(�ԙ�7��>����$�0�x��uї�$��i���*���r|��D{���TF�ؼ�^�����Չ�I�rY���8���Hzj$���C�ِCӱ]�\Mçi����!�1«�=KT�u:�;���r6�ճ7�P>7�8!_L����<�(TǡoW^x@��%�W�g�i^�X}�c�)�o�c�=�����'��w�"��nI_�@����㿌n�__�v,ǭ�1�� �A�ۈ3uԮ�:3�yB�i�V*�t�EE��t_�jv[��{�$�pF�'G��'�ɬ�Ӗ\�тvY��������
|�m�B]#�s+u�.��:���wI���^W�⁌�ƕ��.��G2gZ)�s�P=�K�b�[��h���ip�}�d;���1�����sĵ5���\K�>��)���ckZuBUo?p��
w���:>��f�g������j�Cn|O�xπ�1Q�l{�.�ר��s�t=���V��z�z%�|w**%��9E��\mC�P��~	��*#�M����>�hlk���Q,��n��Ю{�To�R����lw�������7E��]]C\�v�F�P�pE;�W�cF=7��ur���'S�����t�jO��:��d����+Ʒ/�:̾�m{r��.��[�K�1��QK�#�U�K>���7���������i���(踥?��p��U�fVܵy�`��=����H��=�� dG}K����mʳ��,ʄ_�Cu��X::��B��u�W�\ɮ�mB�譐7��H
����^^�.��/~�V��ԅ����9p���P�
�3�o����+����eҪ�t�+��C�F���^��ߩ�<��"e��#g��`�UK�[��ˎ����\�K$$r��]�7E�L���{��c��p��G��j���W���2�a�Qw�c���*E�.FW3�s��p����O���[R��)m3G��ζ	���)��AƗ�\g�]���Me����] ��o�.�^B3E�$UA�efL㮸ϋ�mj�'%��KR�ζ���a*aD��뽔���*��#	�[y�cwpi����W���r�%�\@�w2���O�3L�:�_�F[��3Tj��5��z��M�Ho�g�y����{�7��gf�p@N��?(��sJ~����'y(�Nxm6����!WZ3�O�m�):U�}q;>�f���8 '_�l�����)�7^7����r��hד��|�R�|<3�W�������z�q����_�&�\�f����]^ܺ ��G���p�h�|VxLyTB�����2#��D�#�tx���\�>�dM��n��L��wza���ͺr���*�@����s�����^�?�\�C���O��@��׀�w��"0a����u_�	]0|�Tũ����Q/�E]K��7^�����<M����%aќ�H��>����2}	:���Coʎ_/VS��ς�8=%i��Ok¯e�JEH/v���ڝa��}�[���WhƿD�K�l���H��P�6o��T2a��mhw>Ӣ�7ꞛ�w�N�J�Dף��Tn]���>���P^���mD�;��}����A���p�a����ި��;�ю�k�Êr6&���c��9 �VT�;�s���Z�+gSz���(�����c�:�G�_3�*��Vu��8�E���s=}������TS�MEC�ǳe8�]�Z,Շ���qɓ���e�]L�ۛK�������8~�5k������v��`	��[���8�yzs�4=�w�%Z/ݻr4�=[4{3#�LZ͝�#�'+�c0��]G�+*��Ex�@�`�Q�K�>��mp^Tu�{���Qݲ�*[X��4�h���Pۙ���B���H�p<�|v}\@�@W�:^>�ƞ�1#l���^��q�TW��}q��G�c�[%
D��e�P&x;��|�.����Q�p�xJ�U��>���Qh���+���֣o�i�r"ԐUA����|ۜ���f�-�̷}��O[��#k�[=�=Lo�O��y�{���Ǹ\�zD�_�<���S;'��3�������@e��T��n�H����ϼ�����\{i	�~����r���Ss�5J���w�����c�&
T G�*���P��qW����:�ޤ8��o�G>��b��lw�=3�ko�����Q�� y�A#�n`@z|И|j�m��.=3�}���H<�*�S�գ���W[�7Z����ê�,Z�-M�H~�*K�6~4��C����6�; זE�\��X��+n�é��[r�B�L��˭���С�#�����_��J/^ՙ�w kX��\�l��ub2_n��K$�X�M�D��L|z�6��\���e��о�x1�J�Nq�^=Flj�N����3��e�vwJ̚>�>�)l�����g�ց^�g���J$����b��xП����rf��Wػ�h����j�L\6�fM��>��Ϡ:��)4@^��B�<���=�{�%�Rh��S/7����a�ؼ2󛁌�����ǽ> ���Zo�!����+���@߱��}53���d�%��0��t��ݑLh���c�ϸ������z�9�����h�]I���0'|oB�=�r��7���v�F��G�'��xN���ۗ�����ׂ��"�f�¦���N�u�UH�{j{x=�ml����0�c��������+�o��1����U#�g)�[��y�O��
��yyS���c��ݨ6���ϩ*�?(;-~������>>���'���wv.��ە�ݯ.�*_�3y��E}�YkL��N뢸K�V������=r~V���B|��+diW�٠�������z_�u�C�֣���]$�\�pdL����d��N���G�\}}H]L�7����a��z�g����L{W����rm ����2��U[�Bl�┫�W��v�;>C���k��aL/�Q��X��Q��e���Tiw�^��)�dU/�� ��`���>ࢫҢS1���YiYpf���06�_s����j�P8�ֵݼqZe���
�#+�h2�m�����d�	ד����$�1�tǲ��n�|�C�Q/�{y��ȏu�+�Z��ь�;��-�N���{��}�9 '$p����# ��=�TKt��5(b���Yݝ�T�k��v�g���*���>�g}��|n!����:�;Ǆ�@+N�`Ί}J7sd�F��-��r�>���o�3�N��{�p�{����]�ȹuE��@j�H+�4�Ib���'|�n-j�Ώx���!��z�����3�&�ꍁQ�g�&�Mz�!�/���Vf�o��f���IG�G�;մn���iCܹYQ��!�>'��|y��޺��(h�\ǧ�e\�[��Z�h�#��35��]#���C�Q��3��\��>�z��g��B�{îz�����{%P=�V��7g��V�/O��xj1^\<���C�_�M��Z����3��y�߀�wO�T��w�d��O�F�91�2p+��W���T�'M��x�;�]� dZO�w��Yg�~�M>1��)x����V{����ߊ�������1�C��:�E����ch��L�mi�HjU�5*��H����~	3�����?V,md�0ƶ�g�b<���}f��W�W<��jL6��N�+z�;���A]u���&�1�^���ܭ�bG�Yg
�L��{�1 �7#�݄�:�B���5�v��&�.IO�5�T��Բ<1�z�_���q�hod>��veH�p��3���û�གྷ!��Ezi<�׀Z�;�^^�.��鱚z����=�Dیq��/y��1=.����R�"w�f�˨�Ҫ�,���j<��@RN��5��c�=v�t�x{�����f�ymo:Z��<�.Q%�>F��:�3�7E@�nUx8�O���I��F��k�uÇ/k��٦�WO��Ag�m�8K�r�%T�S"�Q��g���Z��Y�Y�~�;��N�6}H��,�\{d��+�����q�� O����70�2]-��P�QYv��#��}J�4g�����Rt��mA�z��~'�@��1��r�ka�w�Wr/4�����Y�(u|���.�hc���v�Ը�����q�5���f��6zk���]UW�+;w��@o�@�	J%qy�a�|���-�;c#�=�����ޝ ÿp�sPﵒ뼮�z'Ϊ��2K�pH�>��Q|v�ه�_-�P�W�7�z�>����}yw�P�ȉ^܁�T�Z�ds�nOJ�g�C��
q�J�5���M��km��u��Q��t�k]���V�G�Q��o���Tz2(˷��K̾�r:����dc�a����n��Hm�`��IF��f�:����s+R�k�A����?~��כ��U�$atu0����t������w��f������;n�7��Md�D5>d�~􁾇1���dT|�X=Jp��+8*$�K��\����;�
�tfdMT3�m��>̼��}�݈�~�rm�}z�~�q�G���U@���kC������N�̻��W���tz"�i��e�_n]���U呚�C��=4��C��
��̹g#��ܻ����P��T-�r��:��j��az���קA�ڏ�u1Ъ��9�yz{�G��vl5>��V�����0���}�}��7�K0�n��Ex����|�.����u��S댋�*1{g��w�����.7����Ɨ�Ur�He#����^���@�^��=��e9��0���}N�x��Tf�m��ζJd"�e�Qg���򘿩�f�s�k������Koʊ���|_�{��VEz��jk8���4�DZ�
���L�Xy����p����d���.C7�z"�q��2C�_�p��c��Q��y�{��h������%>��)�vަO�t2�m�S�a�Et��g�ѻ��'��sWS�YcEq�".���[{>ÂB`�&񃯧v�#��ĝ���U��}ZCP�rgQz��"Ù�:�+�,�����u>T��Rs]Û�ۘl9���&m��[�Հ��Ճ1��WWn*��v=yFt��ͻԏ��񊞝�$��7x$8t�z3�|�g����m!:o޿\zP~���b�+F�.����^��l	��GҼU|z��*��X�9��=��F��Gx��1=���Oy%Sڼ��wz&������ " �_�@+��>�|���~��k�7�L���߉�[�3ݧ8�����4��gΪ��B�-M�O���d�>��z7vf�[�ƼmFSz����ݡq��O�G�wļ����������2CW��}.{Ƅ�@�����ݳo{�9��J��Ͼs�5��5w&-��"��}���lW�F����+><�*c��߿!��Nd����z���M��9zj�f2c;ׁ�^�����f�ޟ��qZn#�e@�f�O1$�U����F�a;��	���u�d=>��CF�]FDoz��}��<f���Xs��U���̂j�ή����Bilװw��"��+��ѳ�P*$�'�^;�ԇ*����a�~�k���ۺ.t��.�ĸ9���������N�93�b��"�l��n=��~m��^��n`��~L�e�?�����W�ϹWK�Tʛ��µ��Wff*��K�R����wp��8��z��[�Gs]������z�3sUaރ:��b��`��=D .�V�L�\�q-��ev�w"|Et�r�B��I.(�t��j�2ﷆ�g�����D�Wx��z���g�N�O['N�L����R}'G{�l��O���w��Z[�)^��Qڮ^��}.�+"��7���EG�e�Ow|eS�����O��6Q;�h����y3�;��x�4φ��+�Z�~��?��C�֣�*�vf�0m���9���7��^�OzƳ_��$�&���a���{���s�Q����#љ��{�y�:W��^��Ӕx�2�2l	��WFP(�/�㨚����"<����Ƚݟ;�W��������*�����=��p�n@	�D�B�ґ��!x�W{��2X*��J�`��<�P�-������*��둷^�g�6�C�u2Csx��<5C��P�<dq�e�>z}��C�}M�q�޿x����'���ߌ��K:�T	��x��r�V5�:�t��O�\ДwNx�͢^�}E�zg|M��Tl
���\K�>��yd���S3<o{�l��G�rbP���u��f���޲#y�	*d��e�֪0�G��}G�o���6���6���1�m�c���q�co�c���1��\c�����6���1�m���1��P�1���c���1�m�0c����6���1��<c����6���1��n1�cm��c���d�Md��*��_f�A@��̟\�"��� �HI  
	RE ��d �  ))E(�P)Tm� �� �(  �$	@f�"TQ4������fb��m��6m�ڱ�YTڦ�b�Z6Ѷ֚�ͬ��J�mZ�el���3��1k5[���4(Z�2U�֥b�{��kl�Z�Y��U�f-�V��LF�ٔ�UZ[%�(�6�mV�Vƪ+X3dmJ�Z���R�5���-j�jح�ڭ5��L��c-5lw������twO   ����U�Fz�{1�[:�qOGX�{�w=Q�es���e]��q�ۮ�\�qݺm`���UN��@�]��(�ӽ�mU���H��H�kS4�   _O����4����n=;�ϸ��  P  ����EQ���zEth��(Ɗ(��(������(�(�;�ǼQEQEQ��g�QE]N�i��j�t�kbe����%|  ��|��������ɏY]چ�z�8�J��D{���@e����M���:�kX�=t;����@��gu�f�f�kim#a[fŦEVV�V��  ��jCmm�}5��u��{ӷ4�څ]Vw�]�Wuh����i�i]]����Sݴ���k��y�Y�6�<�J��g1��ow{Խ-m���{e��r��-+{��cM��C�I��[o�  �}��m��^�zv��]\կ{�q�"�om����=5�tp�G��m���V���[n��U�[)wV��r8�8�ۮQ3wn۝��Z`V՛ݽ��+km���֔ٖ�mM!ݸFն�-�  ��!+Z�g{�r����X�^���veۧ=sٯV�:ݶ���e.��G]�7R��f�Ww����n��ۜ�n�׵�έ��r�gZ2Wno*�R�۳�v{b؈U���k5�j�hW� ���l�=4��.�m��g%�6����5��:�F�9u���v�]���vQ,��۶Mz����\�۷][���-�l-w6{��{;L�Ӄrc�C�/YJ����m��f�u�  ���a;[Mv)���i��۾��җv�wқ޴Gk]�n�y%%=��v�g�v�퍳N�8�B�R[S��q����V{ծ��]����=���]-�m�z�m2�V�l�Y��n����  /})tj$�u��5�7X���zv�w;�t�޽������^:��lh�;�ۧy�imV��x�׹֑u����֭ze�Y����Ug�oYǽܺ�:�jmu�A�+iB�5�lVz�   Ϸ����E_z�u�Qv0���=s�^�N��z�Pִ�m�ݵ���f���Y[v��˚�����k�T趽�{���7wt���o�������u���<�ʒ� 2 S����  ��S�&�*��`@� ԩT�0  S�i��#�  M$SU ��j~?O��~���߯�K�Z�w����t���ѽ�������4�{����HIN�	!II! ���B��HIO�BH@�$��HH~����o��Ʈk�~�5�&����b��Nr�ܖ��Y^�w��ƶ1����:ۖu�K U�Jԣz�csu�ަ�A1�Ly6t��y�7��jY;t�@(��3�����mՠU��e�tt�o� ��>��ч���'�gg�>� 
MR:��mԳ���n�X��5&�َ���ʊ]UX3��)�`�����X(x]h�w���f�OY�����8���;w��b�@F>����omU�r-������X�f�d����v%��qn�Ȝ��.ݰ*�wf2%��M���xL��7;��ߊe7�;�"Z����`ǑjoE�[�$�o5Pj;7�Xm8�ʸ!����2F4>��k$13�C�Cu�(5���ܵ]\4�j˖�`����<ᬁ���L�E~|_<�b�
s1�E+��eb�&�
:Z�Q��^��$8.�j�[vޝ�GdŒv��H��[;V�/���gr-Ն5��ۋ���&�����kk\*�S.ޓLl���@Y�a<gT�G\[نj�����+b�+f�4�W&�L/r����9X2���D�i�h���	+X����UU�9�+v��CȌ#�2pq���{A{L�yI5Lo[ŋ94�N�VV�:hm7�&F��Kյ��� kH��6���[�(W�E���ܵ���oa(��J,99
C:�m@�:��rي^��!��U��[:�Qlk*���Z�������]�.��h8���ѹԪ6�q7;W�zr�uIT�.���6M��޸�ɯs��x�F��ϩ$-Mꗱ�V���oM4Q�M���P��r�;�{��刖�ìQ���g+pn��`�l3�8�^��rݹ�9�����7� ʏݓSX4,�!�K�� 7@�1��ˢ�nA�<�K�ݮJr{ݼ4��JG�x$/��Ό�e;���O7+S:-C����q�Ȍ�Y��0���F���v��s�  !m@�m��x�9_�qJT2n�-�q�8���i)V0rɍǮF���8��gR
j	nFށ#�BZ�AIL쳰M��5�8�IҢ���Ag���n�̘��s]|�p��ɹ#ǰ����I�{����8���$�越��92�n���{h{��v��J���w1�#:N�4Q.I��MD��w5��KE%�),Qwu���5��TJK`[�bcK �ةt[��S��87���[�m��r��1�v~�V��ƥ�DX,�*B�k�k��m7��l�A���_�^�"�5�φp��9�nG�n���Κ���m�((���GB�St�YpA��KU����W�`�)7\���Z��!���$�B����4�ݜ�c�O\�Uq�k۷�-, ���';��ka�ze�1� Ә/v����a{(f��bCY݇�Ю飻�Z:��r��7�=.��n��H
O��yͣ�\����b���l�
�.� Ǜ����y�vJ��Š���-��CC�����bE3��&Vbt����������f]&i\�1�ha�.�u O�U��������]6_=v5���|Nw,yns��jR\��1��恮J����y_�&��3o0Tp�M�%��Rv%�S�>w����\�bK��m�z��U�w-$[:l���F{�� ��hǫ�v�R#�f�]7���J"k2c��5=�srl�<�\��%]��XU{���E����7tT�e� =\8{��}@�)��aZSX^u�{9ϳ�f���Sc&n֩ekCѻ&Nů�I-|v�ۏ���n��w���77x̫{Ov'I��A czcS&و��k�x��y� Ǥ��>*�ww�m0��&��I�Γ	�tލ��nn��V]q�LĴ9�7���|QE|u�3�B�6߃ƭf��z�R���0U�ب��2��02�m����f'�L�b�i���=�6���!����P�����!����^��H[���U����ǝ��wn�oU;�B�,�e���Rg�`�+ƙ5�,�����\�끓���粗wWf��.�{M�}6j�&���Vv�I1��Ӌb��ѵ`x���5�v���ŀ���z�&<��Z{�ܜ�Rs4 ;Wha�#��]bi�Ϟ�Gy���j��u�0Wu��[OL/Om���V0٭
§H�!�f^�
��L��:���<
@����n���ä�<��)�����%��i�GL����ٺh,Quخ��)7�!�5%���w7�$�7`/��:˻�+lj��A�P�C���P�Z��յlubx;o&��W^xk.;9��sqh�v�Z�zP�kp`S�;�"ݫ� ������ph.WE���qv>��zN��ț~=I��J�B�M���۹��5��	ιZ�+1��:�sF�3�E��&�)[Nun��7��O�]f���9���L��W��{f97T��<&9����x٫��)�Ӈ�؆�+��G���:v��E��E�k5P{u�`�(�w��>Q.Ƞf����>�FT�-�t��ag��m��^c`�o� �	<hg��p1����0r����në�l �M׸���Jo �mA��z���u�O��U�(Xqq�\y�� AC�aӦ���m�q���HQ2k�� ��\D����ͯw�!y6)T�q&9#����j���c��Y8`e�n��`6%�<6�V2#�t#�V3Y2��=���-�iΑ�NsՅ�0���{-�i�x�����^��ڤ��]�Q��l��٪�6+W�����wo-��ᐬ­�����J��8}�Z��{��M�S�.Y�ӑ��vnӵ7�ciN�f�� Z2��ol]�ֹ�ӈ��݅�����dX���{<H�}Ⱦ���yj����E�c"�ml]�4����(�GÝ��ֲ��ܝY����뫁ͷUoy���䞝/�K�c�f[6؟U3z�z*d�m���د�Dɴ��y�Gu3%h}6�`����uXnN��[l����Fa�{������l �C�%��gV��H�Gm4�W��:(9M�*��2�1��f�J�k�F
Gn"��<��ފ��^f���d3��n�А�r-<��lս
I��v�����ln���|��Gmmm�v�&w�m8�h4.$[�ku��}�l3�Om�`x��f��uR��I9��iO���:�v�5�����,���/N �g�4i�K�-��z��ʆ�;�f��N�/��ݛ�=�6�FUù�q�84t;���������y�/������d7�[c_&\""�7�R��=�H�e ��m�B�؈��y�E��9�O	�M�+w1K�U���r��`�@�a��e��Y��5�7�p�׍�������yh���r��|�,�A{��W��pc�Uz�7#j�h�2eX �:�֮��Nu�p���9q1e�v�cVJ�ѹ���cj8m��ʭ��f�}��[���0���Ʈi���*�����"�6t�DU�t;Ol*x�ANG���77y־����dEv�2vtX��ī�P��]�2`a���T5�i��wyKAǃ]��e}[�35�%yP���wY�>�B�.���yr��k��=�ő%�r
Tˀs���v�aEA�1��hH��;-���-qh���+C��*&��\�[~�P'�v�J7a��Hh���3�&�X���(mf9u�����"��V��+�JQiQK��l�;{��
iŰ#�>%5ٶ� +�� ���D8�wAݹA륤:ѕ0���e���trl�'R�n�H,�F��j�̩
�Ʀ��A��jwBIV�	����$z�*��Z�{.�]���Z�x�����ʇt�1��1���)C�Cc&���^oy����5�bZ!�̱Y�n�RF�RԪ�5�#lN��r�B�]޲X�
��+-���%V��Nl�8�\���I 5dm�!6+fR��6	���B�eZ����s�W`� 7w(�B��m�l������r����-Ĥ�g��]+#j��� �YSDZ;R':r۪�&.߮�(疜Y�s��P�Wu�۳��+�@��\����kOaɵ����\���S:蝹r�Nj�Y��3�'9�����GmP�u&ֱ�{����x����S]�lÍj��\O���k�[&0�\]�����n'#(�����A��2]T�#���[6����6�ˏ�X���7sN�7~Z������
�P:��[�G|ӭ�S7���T�����2��W��,e�Wu\�qb<��.up�����@6�7��ѣ��Z��s7�w&����:!(+�A pV �}�]��!_P+]�-S�IQ���Ս�%)o.��Fi�;���0������d�~J�0wyir�}i�[��5�ec
�&�V�ӻ���5���'�vr� ȅ�=�v`JLQ�@������z�®�x��n��(�^ӫC�/n�H�"*#,$��2M�(E��l�m�I.����A��#P��r�\_�b�Kx�8�IeWst���𣸄���e�n7�r��f+Ӳ��%�鑫���k]�&�<�F���}�wM�K8��E��c�bދVwV(h�������12�M�Yoݽ���B�)�R�y�%�f�o�6h�l9�di���h����ǝv����Ep��.Gbަ"�R���]\��<\���hu�o�]w��~�p�G5�s4��JF>�N(WR�F'	��w��Ϭ .G 
�R�pd^�B�����T���n��S���j��9ֳ+���"��Z���ڶ�����9�>|�x񌯱ذ���q��Y��$�Tv�w�%��#sco7�g�^^WN�L���Dqqz��:�ۙ(p���\�h���V ���חI�k%s2��vEн�4�0]ӪL�܁�.�l�9b/ZG:#b�[�8 U�w@{q�'�;�l&��A�pF���SpnW�[�t[|�&f��j~C��}2L��g[�gv��t���3�Y���p�!���xP[{O�wڡc�&3r-=�E�sG874��A�{����u�̃N���i��R��S�Ɉ^0��gF��orG0ŧ�ח��F�e�I)3R	��(�OpN�JE�nJ;Rc�b�n��M)��2�(`O��� q�3+�ӹ�Κ.�%�a�R��/sX�	jI.A/H���x���̮o9��#;9��3#����a��4�XLɂ\�aP�u���L�w��+���4���r�9��T(r��i�L�Q�F���%u�f���ob��/S��n�2#�{Y�m�D9����"�x^1�Ł�8�����B.��o��S9�#�[+��q0f�/O4���b,�M�6�ǻa�,�y�A�	��sLa�j��^�Ä��\ݤ��U�p4�͈�7vc��r�MY0�g4ɺ_#�q�
�(w{�Ž2���o%�p0l��N-��]B;�<Ր��sN`�,VǍ!WN��e���k��Ĭ��C�q�7�;'�4�N��x8ʺ��#��{��'�RrwI�bO[Q�TӇz��U,<|_��[_,�ޚ��UǕ��R���7��R��P;^{ǒֵ�7���C�����#x�e��I2����~ٽ7�����xR��˃kx'h�#4^���Rm!��dh�0������t��|�%��/WW��8����wIP��P'��K*|��$��N���+��
���~�9L]p�vԄ��մ�.�kS�觖�rٸ���Z���D=�;�^h|1o9�y�6v�:����D��ot�)����Y˶��Ϗ���H��C�������:hѣ%EDD�W������>����l� �W�ehC��CTJ��Z'iʬ�@�ќ ]w.㨴�,�p�C�	��*p�nt���N ��r�э���zE���E����:b�l��yh�1�C�׺�p{��z���Dv�c`��80V\L����J -n�<��F��^o��\�['*V�-����7�93���Peֻ��u��V\&�n�63c5,bǫj�¾d�����3����ٛ�	������q&rjyҌ6�ïAh;yT�r�o��=���`JMF�[S6@�;+ �J�\�X�y
zg�UyG53�h*��m�l�)b�� ڦ0^���HӋEF���8�ܹ�D�7��\Ps�9cGZ�껠���n8퀊5}#�*4r�i���4}�TD +����I1�t�LcSNM��{��59��-��Wf��p�ی����ge�r�r��cI�;d�wNvH��31�Ž�3Sy�a�S�I��楅�˰�{	���?��:�	'6�Sx�db9U]�x��a�%9N�"ƫ5@U��X.�t�X�F*],�0ɹ���d�L��Q������Ï������O#܆w`���;�.����B���Q��dG�L���'�o;��RY��yzU�+厊Y
��^�E�Nu��jmn2)է�f�dԵ�˄�Vv���	.�ݷ�`6��w'Ft���$[�ظ�����{'��׷����j��i��hy�իo����Z�U�.R�i�##wCP��&�v�`��mv�}�6�ў��sڰ,�b�O �V�7˄[����X��(��Sl�)Z�hZ2�;ẏ=�d��o���e�F�V�G;�v,-�]c�!r��E��m��^�1W\6v�oS$.��)4W�3k�<ާz�+Ό+*f��Ns��$�>�K�Ƨ^�a�8�WԖ�lB���oY�Z�C��}�Wk���r^���ӽV:�����ʈ1l	���G+dyW���mGg�63yJ��U75S�Օ�f@^��SwX�nN�4�aMj;�D	��c!�鋱�]�i����TfQ�Ҷ
g���w�������8h9��I2-����ARi.���/��TM�'���v	��M|���Ԗ)��K1����۽�fF@�3�5+vh���a#�?�r-�k��_s���b�\-Gf�mH�TU幕�)Ԯα9K�~w3:��(��ܻ�'���cs���N����!wo-����\)@�j�a
�q�\�Ve�i�`gS����fk=N�GG��ѻҒ�4P�v/\����$�H׽|�\O�9ꓞ=�8�ٮ��_ �S#������P^��ٸ�J�=Tq��t���g�jH�?X��LR�!-|Ǘ|�E.{���*��g�=�_/n ���nvТf��xi)�o���{G�|��ƫ���Z� f�_P�Z�X���:�w���z;V��B�{ҥ㱚ֻZ��?i;mu7S�gJ�>@pWA`��ǋ��2��6�v�S��"�2���z)6�QZ�N[n���i�˞�&�z5�HF^�|ޅmmeGp���m���8��<;���˕�L7[�Mcx�W�{K����B(�ai1U藺2��gb�@�c�����]���KMR�1��t,����+���6K"���W�A�>��p�tMW7:��I
���@H#G+�u��;��Z��P"o
�%ٙ��@,|���-e.��H���nab`���^ag��|��ؽ�"q��9��tj�����˷�\�q��I��C�ػ�_@y{�� �4~޷z�{�J��R���4���D��yCQ]��vtyd��PU��ͥ�0̇y����d��:�:���ڀtx�˚vGv̅�';���u��W#��W�v��'<��rE������Ni6�v��-�wd[;�׹��⢙6��,�#-��L��d����O�X�"䀫�æ�@���+���4l��ش�<o(EG #���/�{y�X��{�2lY�D�4��v�Mr�s�C��^����۷���2�V���7�d�Ò��+X����+8'x�{&��8\�-�Ӻ�z8	�Hz�t��闦�QyI���[��gF˄ih�s!5{ɤF��ܵE�s0e,�+$��\�Z�)P��(�G���oy�ϣ�2ue˷�U��,�)�˗�x�v���YX)F-�r��2��#��X��T�Vvw$��'1�*L�z��p\>��M�ZaW��Gm��Ν�΍ζ �/3k/[HNm\dB��o���f�Z��ŋm<��[��YP��������8�u�Жr�V��H∞�L׹Nq��&6��F���o�ʽUq�`*��&���.�,b�4A�\>��w��݂<챥�Pg.�u�9-�Շ-�����ҺT�ݴ�����紌�c�>޼H�xe��l�0;6{O�8��=[^F�S'\2���<��>��ҡ�s�[���6{Iz�`]�"��2¥H�˷@��2ܦ8�u��~rӂ��^��u��)0�B�c4ɓ��\��w�׼�	sa�Ǆ�V<䖌�/�T�`���0v���{���ݒu^���B��X1�P��=g9�!u{�H&�.c��X�]ym�2�*��H�3dc;qk��B����&�����=���1�Z�6`R� �Ԫ�˝���Y�5[�X'7EH+I��}���s���*k}]Y]��o��t'�m����Ec컫�M�s%O����E�-�8�pq��=*���ďV��՞��Q���1�K���3���Id��"V�\�+pI�nC�yoS=_��ܦ7��'�U2�,�6�.�c�\����[Z��U��]'/���;�eʽ d�V9�{Z1�Ýo����-�GP���ԩ�Q�⎾���b�R��[�R ��T)�^�6'����[Wn�gLݘ]���И�CWF`kO��[�z�u�B���BS�4�᛹R�u����	�plJ�9�K';�o�j3���]>�Cą�x���a�8���"�#������DR��wv�{Mb�>����V�p����{h�Z���B�Uq��c�f�r ��ap�-���� ���%�c�W�����EE[;Y�;�w�s�f��B�wv����2
�����{��ܕe^s��]��o��IzWj�ԭ_1��;$�,��~ԛ��71�
e����+O��al�N����cg6V\�����Ng,^���@�#�/y.`u�]wM�<U�؈ ��(��4�E�j.yh���ŷ��8mѹ�\c���oXNp�.�Z4̩�+r�3"�B�����P糆CJݾ�Y�	e0V�(�>=�.sf��:{w+-1��ٜ��guS��k��ϖzЎ������Uo�ў9��@��6n��%�9g)�����x��F� i�`,�.˫|=ru�5�$��gm����|��A��}rͤ�`O��Pm�.��v�#N�yi��ԏ����ds�*얢b��-���<C��݌H��7�����y�q7�uZ��7]lsd�jf�<����fu#Syp�S[��	%��h�]�`��|��<H�.2�a�����:�4wPf�mݍJ�sV��5��L�p)�
���ޓA��v��q�	u�K�p5� Yuܩp��!��o+U�G�������m��i5^���D�q<_�Ofz���1qxGR�u>�a$�浂H0n8ِJ�wR[�P�c"�{m*��9x�?�?�v*ݽd�b>R�}����GK�G�j
\�%C�=��*Dwv���i�h ��m������GO�=a����������,q�S��{����n�.aȥ������D�YW~30q�����|t�u�gvn��7fu��41(F��蚛I��7�=�4����>�8�v(��}'K�l^�{����9���R�9�{K�rմ�I��ɤZ��W!����/�%햺�:y�Wqh�X�G�0��ѓ��V�g7�ƙ��[y�q'vR�j��z��,����Ddw�f�<�o4�@�ڻ���n�<��7�ڨ�IZ|Eܴ��t�ʽ��v�V�+xojD	k��m���m5g.���x�DrMԫvY�<�,X՜�[���ثD�	C�31��M��L��ޓh�l�:nd��A�ڋIΧ���+�j q�]��zf��]�b�V��T
xe�o��A8�:�a�-sŧ/Y5����'�~ z}T�uG�q�e�5`�K�跷�$>��2��X�m��D�R�8ƹ���.LW��[�j�� ���D���5�w�7 �y��1�r+f9���1+���W9V)�}1d���B������9��1��Z�r��nG'rc�C6�f8�w��U�u�^(s_��c��GC�<Cy��) E�n�]b�t���wQ����wJ�%�Ҧ�N�N�w9�h��^Desُj\�Y��ɑP-�ռt�A���sU�H�iS��"������3w0 ��(u�H
e�Vi����Н��>y_�g�xn��9ޗ���.�S�.�N�\}�R󯔂�_.d��f�%�G�y����u�ɋ2���jr�;Q�B�����O�����a��ګq�*]� Ӥ�G-�ä���ζ�©��G;(d�Y���P��1L[w�W�f܄��]�ù��$"ʶ��Dd�
�'Y'{Ũ��c�<h���L����J!��#�_TR��S�f�Ԭ��%u��R	k�DX�&e��쭭�ù*9�̶s����.�(Ջ�I���Ahl�U8mpLX'h�{��h��{�۫�d3u��[nAOUկIW:֩��,y`�w�.]�L�{T��M���sWM��-Ւ븲�)\�h��kP�H�W�Y�Ke8��y�3wg�/�:�����J�N�!��-�n���n�gA�7�4Vo��өm��/͜:��H����\�ח�lT����8]+tҩ����u՜�5�Ws�I�.��<u�Ό4y?Y4��aeOzev��.������(��	=e�;���R<X�ח� �بn�b�A`aU�m0J�N�|]��w���וɞ�S+.�soVWnPn/��O�����y�Ö�h�B�!��a!�5�w��Vζ$���+mόʜ9�u��N�Q��������d�'.Z:њIU�r��RD�:wG@^!(�zf�
�뻒��De_���^ʂ�l�f�G�6�XM���Ot.ķ��46�c��9��#��-mj�Ђ�ǯ���a�Э�j���7F�qt��Ռ�f.�i���)i�����n/7ច�=���s�syC��d�2v�,U%kw�E�x��!nV�3�w}�y ��ո��𘱹/���`+o��	��y,��\{���ފʧ�b]��"R�x�� -ق����OK��S�x�Gaw���p���[��N#���|�#�����٣�Y�ۑ2���R���͋��J����]��[��-���Ӗ�'{�x^��󓮀�� ��n82%Cw���K�jvۗo��@e���/CP��ƃ�� �8�{X��R�k����*��&މ��,K��d�g�u��K�-��n�d _9�@�b�pZª��moh{Ş9W==w\^��8�ޖ%�t¨~Xh�ͅ��e8��/]��Ɯ��^Φ��8m��+���E});Z�56YǥT ��r@*c��b(�`Wg[��!L0�I�j��r� QH�U͕<�=����JLkڥ^�ж�0����2�n���c�0�0���M�L�.B4��F���t`O���.��~	$5�s���̸YJ;5f�N��cS�(cL]��ў��c��e�U�`�\ioϷ3�Xt�b����Y�R�R+�#eV�X����y�+x�x-`�H_O��1Ts,�BWS���;�ZF!g|�Q2�AR�q3(˒���Y��#��:�d�v̍�����Kd��/�Ge(#��\/j��s�R��^]-�ea��"�Y �_1���dѸ�כ[5��3:�ބG=�嬮Ft���4:W���T��­3����X�cf��A���Hy!��E;t���:��F��Wzu)��V_j���[{�e�*iwF$����4g2<6��UwFS����ӄ����3�"y�����k���|�����4���\p	��f�X�H�E��1��J�#��`#ý����>q�LO�&��'3��W5���9�ʵ������*�ܮĴ�O��{W��[��=��:�3�Q�[}4*r�<�?��ݼ~��o���	�	��U�=J�b���?3 �݀�����EW��aaN�]uy��ө�vGh���Wi'ټ����	Vt?;%[�=����=�o�8���y�z|6�>ݚ�bV����{���2b@��B	��x=*�A��5z�wW��Ir��$<,������3ۋ��sOlvuB*���ӫ���ݭ<$tc�꒲��X��a�ss�M��07b�(kZw�S3ke�� �Ҿ���#��Թ��N��2pS�^S�]ӂ斻�9Y%�C!Tа"V7�nU�X�t�HTm�ӈ>�ޗ�R�$�k�\�!�+�3��B p0]���AQ��I��fu7��D�v���1w<Q�[�2�\#.�@�W��(����8i�{ӈ�%��]b���V��4����e�F�YZ'HE6�(�P2j74�'S���.n"��o.�n������$����@^^ [���wt��V�E�/;:GO�?pN-�]-������"�ٍ���X]�w���O 8���î���N�;�4�/�X���^����S,k6l �����8��/��<�F�.�����F����gV���v�+��{=�{���{��6Mx�t�F�Z�Ym�"^�?>j�����:e?y�}tJ���vC��%O/�a����Џ&���D�]-q��B�C\\4zk�/d����S|��̀�\�J�])i{&�o����!Z-��	٪�0J��ѝ��ۻY��B}7P�KT�,`+�}�5ӄL�N!<[�#ֹ�1h������D�,�����&�u$V�1��^�i��3���给Yv�d��Q�=���؜@�}{���}��4<Jaz��}���6�S|.ēK���oZ�%�*��.��������ԩa��}3��k������yz���J�`����%k8l���1�S�e��<e�Z"0]�0o.Mr.s/����Ͳ�H�4sb��n�+���2���yzAP=����7�I�����v�A3f�D5P��nU�ɱ$�;Z�ov:�A�g\��C%��=�o-N���M��~�=A����]Y�����.o���厭�O���Ζdrtُa��'n�X�vI�8I��-�����f�	6���F@y�}���I���BH@�w�y����y]���0b��ޱ�Q�Ffb��5]gj n/n?~/k^LXlz��'V3rX5�d�l>" $8����H�4
R��N3�R�Z�	Y�%Y���&f,ܦS[�
D{w��I��_�e�5���qˬ���P�r<Z�Z�!��Gf�L�qu<�މ�P���ͫ�����A;�n�h��!�k��Ǡc�J�Q�)�7g��Z*\�J�]�{K�a}=�́��~C�wmk�,q��5w��rW"v���-�t���a�4���WF����� oU��9���+�]�+�����CO$�ۣ%sN��	��	#�񎩝�ϗW��6�9MB�{y�O��oOܤI�c5.��V���R^zGr���z[!9zvD�F�q��|��^��c6�Z��6i�lΝk耠x��hU_Ƣ�� ;�]�Nsy��M*�@��j��y�ļ�R�=E����X�����bB���J��@�w/g�W���ל��8s���ߘ\fQ��9���ۂ���:M#��k�X!VwcWB�H[׆�\��W�᳹�Bקּ��.�$�����&�b˂�2�����T��2��@J7K��݊�5$���v�΢ֽ�_X��[˦�K�pt+U��j�sc��F��5a�śYV�(q;�N5܇:l�:�������gI�Q/M�r�Ӳ�x����X�j��9���/4��\�����I(j�	��a���9��nqu�_�תfwj��m)����]1W��gk@�̐J�}� ��bT��LZ}ͦrV��)�F���s3g�]@7�8�6��ֽc�7�Nc�V^�f��]#P�m@hq��|�U�=�؀�z��n?5�bQ�ygwT��h%̾=l��;C4�K������V��d~43g�����6WkΚ�����a9s8��w$�L�*-�.vn��j塤�X*;Q���Z��P�*�oj4(��k�����3���Z8���b&
z�ݕx�z�l�3���*�����vΘ�r��#jJ��e��N�I]��7.�"T�w7ɪK�Ϸnpq����� �F3n�\�fF^x[w�^ls���ŋ8�of�ֺ"�lv��[�v��Č}D+�=��cׄ3B{�r�l�d�
�N�E�"�����Sz{G�#X2N���n���T ����Þ�op7�/�i��j^	F���<�+�~���;o�S�)�8��f��sSj�0d�o�X癇 �;@��'ݸ�,ُBI�r��O�l��A��A�*�Բe�9q�5}�e�Eyj�#���2��5�.yW�T���}w:a��ޞ`wR�i�»-a��ۺ��D�P/K;]QT�Ǔ�������-8iݢ�����=�K���"M,��{��+��ʳlV�OG�5̭��øVV_c�k <tF{5ܖK�,���rʨ�*���8y�6��/bq7{�?o�>�B��W=H�珄u�l�{2¾�6��E��8/o���p�ܙ��v{���Zs}���L�bo'n̼���8���e��J@uq�v�o7K>ۓy�ͧ�a��s��u����}"�R=��3��gi�Bn�t��N�U���퓮��+zI/o�8�hc2"���'P��샜��T�R̈́J.��GC�}��k�b�ۄ�Wo��\G���w��O8��N�`��:qX��q�>֘�R��L�7X��5!D���xji@��=��ǯ,1J�����2��7��#hB��K�x�5�Zyǅ,(�]̝�1u�6�pkFނ�`".�K����7�tC3�V��`�"_:Uj%�kbB�a�c7�K�f0(������3o��y���x?&4��E�\�yH�՜8O8~ol��vJ�o�)�y�ouݨ��YKq�Q�ka.us�c���ϝKVvU���!v.JǻG��{�ǭK�%x&vy�0V�;��¬��vML�hQ��m� �&��2�,on�|��u
�p#wq5�io\'S����r�e��Λrq��i�q���+�C}�ݢ��f�xG���
V�"�,s����Zs��c�ɋ�����+� �}~�|��{^͋�H�{�}�n� ��L�a�Ҷ(O���+���Bʺm2��kg�:y�Mk�a΍��Wy�M����t�l�"��6�7���҅���݃�����]z��U��_�x
��6���Ƈe-s+�z����nE(��ʨ��n��GG���/qǛNn4�PW�&�8����r�,�R�T����c�5���������.�Y;}�3,��������}񫣸�f]�Ib/@Mћ(
��w:��(�\�PƳfC����&�������瀰�����8,;��-��ݪ�.t*g<�˃�� ���{^A��<��쯜zvٓ��e{�f�1��u���x�W{�*+�R:K.��yY�=�����s�yV?�<=��1����g���Ҷ��گ�$˱�!0	M�v�3�jޞpb��uz�e~�Md��SM,8�_�!�<*5�K�Zj���ַ˸�Y7���+9���f� =���9���I}7Um�wGu�Ovn#[��G+��0��jN���.����Z�g�8�82�b�	�ʄ^���(ɞ�Q�w��c=W>���NK�J����cmYfω�u�v:tb����y��Í����v�����{C�;lCY�/8�W��� �;y���c��}�2�M���u��
�w�\��[K�aGY[�6�5x���D[��h\�U}'-�=~�m�;�'��5�'lIQ>�xK�U�dGЎrv��Q ٦in�ѽ��=C��W5��:74���'����"�)T��.Kەg�j=�7xnW8��tG!��i�.�-���t{B�d�3B�V�������&Q',x�㞙�mv��!� �}/SW��",���|V��[�M�k�[����}W�����3�aK���T��^�����a��n����6�}���0��虘}-ûΗu�ڝw`W���xg҃a<S;]]0�vf�q�ԕ#n�Y��>$vÑ��>82��
��r�ݙ@�W��.�PjK�cR��
��"���������=�k19?dB�I��޺�X��5n·�h��١Y�l�=X$^U��x��Uu�#b#.��u�O:4����e6�Ngi�k��T�7sLTYn{�{�~�"M
orN1��/�匾0��a��x˵a��.�;>�X/��Y��8<�:��纈;ON�QƍH�n��w�t����9=��6 Oܻ#�.b��czˤ%Ы���˨3� �3�~�=\�D��<'}�v.�4I�y�Bg�޷P���
�m���f{Iů��։p�����[����U+v=�t��A�rScj�F����j��HX�Ѱi���-�i�����GMy�$ҭ��.���=U��y��"�*q-�E[{Z�em,C/e��A"p�d��$��ñ�v�F�\�w���Ɲ�rvY�o�}����*'���;K�OW�:IOx/o�珠~��"���ʖ�-�s���(Uq�ANim����I�����Jŝy���j�U�ʼ �I�i��8�%m��p��s&Lt$V/6�~m	q↊��u�%��<��]��ڻ}��ag�g�+Ջ�uu���8|��SzZ��f�j�;�ҁL��I��jʏ8�S)�Hk�Q|����0ʋX�����A�́ ���o&杹d+��i��+Ydu�ă% �U�篫�KJӻwdʡ2�[u�[�X��q�p�fɫ��|�qN��^x����ʅS���- 4��� ��u�f�6�Wr���)�ʍLc�.���^I�|�h�bk��]u*�mu	��rt�(t�/T�3��ΒZEѭ-,c��z.^1܁f�+b�h}4�	P��8u��0΂�]��Ѭ��Μ9�A�Je�A�w��*�yë��pZ�3٩,d��\�h�AΛ�ׇ}����V�o�=���޸��F����%�;���e$~g�AeL�ikK��:���mͩnz'�������:���R�mv���Ǧ�X�Mw�k����"���>0�u���\Qx���ܨ�s5�u��T���,^m4R�M���w�!cT���Û�ץ݄�v��c���e�"�|�r��\2�f��9\���s��gF�$��v�0�ddC�`�ئ��%7���k��ؗ>ڂkyQۣ|���6;�A�ӫ���h;e��$�/��laE���tR0�MO�5�]�#��K��p�N�oP/��LE�[�NoB�(�Mug:�Qc��K���:��M��z�{�0t���Ut޽!�x��{�~p��힟-�.YǗg<��ss���7M�7Ѵ*ʽW-��ѝ#����BՎ�ю�Hk����N��t����k�G���ԩ�'z�7�^�y��2���h�!��� x��i�M�)���X.�h���"�6��^b��iΣW�@#y�X�7!�wbA�A��VTՀ^�:�'sxEǏ_>�m��@���� ��f�u!QvwYX����@��˧`�fƸlt=#�R�r�ݍ'�M�����keڰ���ѡ�u>
4��@�K����c�V5T��_;�Y�E��wxԹ��/n�[WYy��U�	X�xJ��������/i=�9�sz���+H bF��k�󱸖�=��b��̵xdk��m���ܓ	8�F���N�4 U�9����ڈf��,�Cæ��/i�Syqҗc,���kӞ&&[�M�����5�����9��YҟcvtS�o��s�[DY6���|�;fC2mԱd�R������z�3l�\��Z[ڸ�1��ze,(�+�d��솟/k:�rx��7��X澝	��+��z�x�C`�KLaYj�*"h�o:���\x�f��z���M�m���|���1g�3��mJ
���*f޽ȭs6h❙��D3U(=ǈ9��n�SE`Ё)���|���
]���:���ԥ����)U�bb�Vųo�e����b'��E��Ε��Ȭt�T��F�}2���F�!nΝ��3o^�{Ku
4������^l6P4p�Ǯ����ʱ֖@z��A��U�k"��0��q]ny�� ��L��=�A��LY��d�0v������Qʫ������:1c#��4��[՝�Ǧ�� w
�f���]>��*<8m:�r�e'`4�ξh.�G
�ux��7�]&������L�r�X���ĤYc@a�;m_#����{������,fo1���+%�p���"�'�J��E��W�;54kH}H���q�H��B��;5�79:�4�m��n�pH����;�}��Q��.������+)�FV���o��
;�7-��3S�3����� 2��lpWHJ�-���ݘ�c������y0�H
�y�p�b�n����;��������;��1ci���	�����z{��:>K�ϕɋ;q�%�g/VX��b�Uꨟ����р����"����ݘ�Ͳ�ӇR�]ζ��*iSTc�=��)K��4RCeb��:B3��a�&(�<�PךR�)�v<�Ήv����{i��]�<����vr�f�2���\���b�ǍX�N���중�A5�N[��7kLJ��X��M�ti÷r��yk�)H��e�[��m�$�N]�*�@ԺD���(�6ht77Q�C���=&�>N>}phٞ�Ӣf�)�]0�w��[��ә����7��+ww�@cyZ9L����:l�ǎf�y���b�lV�� �˧7[������	S˨G��C�M�I6.�7�g��ꥁ��[���n���p�ru��G6����Z��)	hp���H�E:���WV�oX�X����U)��+x\DC��vr�:����W���"�Gv�.�'Yלw{)��ȋ��^����\�k��{�x���u5v�ⅉx���Y��s�MM�Byl#O��q�)�!m���p*�˹u��A�y��7������G�nB_J��Ah�Z��	1-��6��%��7ܛZ�];�٣F8��h�t6��|��(X�cekY��Љ4l7g��M���=ь{.=&��K8h��/��8h/<=��b{&���̽ͱ�� U3hs�i�gu���fenF���y� w�F��4�i+χa��g<;�/C]�W��O_��� !��m��n�fƵ�(/�L�7B�0u�L�0E�3V�+�i��F����ou!T���w���2��Nч�U4�ܦ�M�:����j�ըN�x%wh�5 �(l�k4� ��s�̓q�U�L*'t2Եe����YW���,�=�W�tE4V�������%Yq�|�|���h���L�{����T:�x��W�ˇ�x�x)��O�ګS��+ޙ(�O$0=���Y��Ί�v\�]g�i̘Txe�|��;�cGAN��i�b�8t��>�=�+DZ�}X�5�ŋ©;����J���Qpٲ�Z�c��Z�fS	�x\0<j�RxS�z�}��+�g_x��حR��l�6�3]k���ct�������哓{�:t}67� ��+�Ԯ�����+�Q��B⽃���EI�{c�7Y
:�DӇ�''5o19�{�da$B��J^�=��l�)7�tS�e��j������������������	!H�{)k����x(�J���ə��s\�9f���r�ᅜ�nզ	{�J[o�rx-nuȬ!�V1*�ŻԢ��w-�+�����n8k��1���+�Fh��ھ���67���G��G� ��n�o���n�wʹT&Mef�u�q�jb[�Y%k�������m-a,�p����ǰ�eg{��ș�zi<��,���{݋�#�n�{ܹԟ�9�>���
��\�	ͷJ���s+bz��8k"�~���'X�<R8X>���W�e���I���U�}��5�X�il,e�Ku��ұ��h�<1#��r3zF=�S	��Ά;7���ޅf���e4�������yB�9��uw�o;+��{��Fu�db�i(�y[��i�*Jԝ�TY��Z���-�:����%Ϭ�7R�&��+;m�{��Ҭ8UbᷣD	�&�������k�Mv�S��-�z 3+��w݌����n�+y��}��#�l��Z�X�w�f�ٮm���mݭ`�7�z���C����ɪJ����m����̺����Ncl܁1+��?���{�y����DA0�9�!��=�à�C{�9n���)=�Av���5�{8�ͲW�c�2��EN�Ks�*�uƸL�I�*���ɬ�.g;����i훱�z�r��Τ���x T��]
�����'V9��Ȩfgd��(� Q%�L�F�Q���խO��ƭ��؈�*���lb����V�J(ե]9�	YJ�Z�ֵ*[kR�JXV�bڡX�%T�ҩ4Uj��8aEE� �1���-cV�YJ���j�iVѫEZ���kiYZ*��`ۧ[�bT���jQ����*�"�"�4TV�-�8�j؈�j[[V��Z�D-�b)�DLf3�Vմ��mDm����m��J��Ec�aJ����:D��Ɩ�#m-U*���j�QU�t�G,*��V�Kj5m(�b��FV,���EKZ� �#5p�E��-UUX��*��Q��F�VTc��Ԋ�h�"DU��Z��D���R�J��+(��%,m%IU�9��e�1�k3U�%�ei�EL�����(�-���QE���TF[X�jUTUF*�J��1Dk(��Vږ�TX��h-�PD���YU��Z������£HT+U�X��9J*��U+�ؑ�[F-l�(*���#�o_�_�6)��VOK��su���2��w�e���W�<imE�b3���v�'�i�������L��^�b�;�N)��'��m��l5�����ur/yR�z��X��,��c�fv%�sG��4-J���+��kB��[�U�D"�s�[��9 �p���1{<�z�Z�:\mt���1HeTf��9[W��e�'�ڥ�Kū���y�_=�%$��+T��u���EZ"{����ECadY�z����x7{��5����u,\a���=�WJ~���T��t�Y�	��F��l�k�O�.���/n���ǵy]�I���]f)Y!&���ǵie�R2\r�3i�n�kv�_NP���	��[�u`^�<���0�����U�?=�V�s��ZЯC�{����,GҷfAE٢���j��"�p�$�J���n++�{�V_&��{����s��j9nL�\Z�U�3O�2����+Ӄ:�W`LTbN�S�q��\Ci�K�r���n�����g�!
Uf�X�륒e��2�){5��)�A�:=�-Zu�k<^���Z�*vR�wî�Ͻ�$��F��������A�F�vR��P;�r�6�Nݶ9���3S������U#cik�465��mYS�z6�f�\>1�l�&	�S�V���qy�Dil�����P�9�k���F�7�]n�d�o�ײ �?<��`��Ye�Ӯ���Թ�z�!�T�Cw�ޙP-�ĸ���'m�m�qy���T;ݯ �U=<O@�Y���zދmM�0��&e�iI�����e�ޖE>,P���d"�Cc��ȱ�
����f�6��vݏ�I#�^�eg��bd�~�+���d�V�������ns�]>z�2�5<삯:����l�St`	�!�5N��=��<VCc�x��[1l)�>�X�}~���e�G1��n���]�*��{^*��4F���k����[���[��E��U��G/��_M*��t/E��L��ћ�(.��S�.��/�1�2ko��a�܉2��\��#��5��Z�L�
[��9���{T�/�ީ)ˈ���B����1�ߙpZV���t@��ˁ� �o7�7SLyE�;�2˲(U�򳮸<��^�Ķ�H���P��n�D����3�ՙ���ʟx�*\nE�+��f��+�xGā�Md������v7�c�}l�nL�7[Jm���z��أΚwz��c�P�-�K�ٯu�]Ln��|0�urOsܜX��VKW����֧^ZЧ�۹�
U��|3��Bu�ZZE&���^6}�?D�J����G\���4�9��]ԋ���u�7���÷v����7�^��N�6�
�4�ε�z�鶔���n��M�{��p�)�~m>܇ov�^RBr�ܺ/�҃���磛� �Tj�]J瞥6��_;E��y���SAW�����A;�j���I��lYR�����'�����qB�O]��\c��~�x:����3GT��u�s��|+���:v�4����̹�mt��	;م��yO8��[��}��*DN��E�XA�k��ʁ�v.ơ�)�M�;��݄7v�F����w׽g`�"���v�9V�^���L�3 
�T4Uʔt:KԃU��<:}�ݸ9T�&EE���n��Mo�|su�k���]��q0��4��x��8L���8�M15P��Z�vegU����[�ܓ�545M�FwMٕ-�y�R
;2�]	쳱�ڽ�U���B��'�oFjy�˭[̏uU.b��|󷴺̀\����̡�1
d�騕�����}"�7�J��Kڷ��V_�u�q-�Au�z���֪���\��n_u�ze��� ן���ܭ��r���Q�e�V�L�M�������{��9~���OiNz�1��r���C%��ab6�r�Ҏw�t���r_^\�.��二ע������X6�8�+z��G��9��5L�����勏��	���8����z�y����OM�V[�9{~Sѯ,09��$ݱ:��v���ޚ2������P໲�����������-=�Z�P�܅{��n֗޽ꢰSwx�v�R{U���������������Ӷާ۞v�n^R�9F����f�Y=�1؜嚠r9!�.�9��!���)|�k1������	\}wVnS�8Y��۹l�Դ�YB�AIF�gbd��O�i�{W���PN���2�4��4��jU��c��-At�B�J���陉9:v;��%�c&�S&�9 �������*�nw)���p͸9XȃTguv���f_E�{��!��b�����K�ʟCA��ßG�`��e�TOh�[8��MSԷ ��<^�	o]Jw�O�{��ϩ��衶�a���]��S�Zek�q���C�1��xc��OQ}u�'��لBڹ���eC��Nu����NV*{��t�����)�b�=��r��/*ܙf����W��������zzx.���z���q݁&	M�,�)�@�X��)�X9���c�iﾯh�M������A��&�弨.�RvG�Eok�ҙ@����P���H��Ux<��2c5Q��B*��6���U�,���U,٫�'�l��t2��"��i�*�K����֫w��'�s}G�$s�K�V-׺:䮼�Nb�-e���d��?�N��3:�y�G��6��qP�-憽����j�b�9�[X�o&���{�n�Y^|�N�Ig�sZ���x^�����)����;�a����vl$�8t�.*�h�m/o�f����_��s2�$7���.*��:Z�,DP�gVm-�x;1�����;��y�nI�{8�U�}c��'�T(8F�t�8Ffm�R�Z{���R�*|��E�¡�Z-���������|�z��}%���᮳���2�u��ѓK}[p��O1��>櫳coK�}�Y\�D�j�����Jj�V�u��Mm�mk����H�n�_s��o<*d�5�
�/Ӄ:�W`LbO�t�>��ŝ�����N�ƭn��y����;�JQ�l�u�$�yn��fP�J3w>ҷ�3���rIr��:z!���G�z��\�/�䳕E��6NUܐ��\��9`�3��nu�P���Fa<b��λUk]�q7�d��fP��)5�:�Yy(��/!�C��c����`C=B���WC���)�M�ʸ����>�n��!�`�Y5۪�)��f*D?3����W5����t�	�sS�'��`�pg�,4�����(�	/;����B4��	�pa��9;��e��W��fE9�]v���F~�����:>��7�v�%��P�HNA�^�97u%KB�b���ɸ̦�Sk��b����]�"�y�x�@WkmݫT�ϟ�:�����p9w�j������X��S� 5 ��d�['w��j���P���u��'Pۨ+\��u����1B3�ũ�jI��wOE�䖤��s�U�����.q�f��=[��m��Y��0/�^�~���׾�Y���g(	5���mT�Ю{v~'^�5sU�B_z�d+^������R�����ac�ݬ��{{7�`J%�
���Y�T���[�*�N��xTte_��ާ��'���(�ă����r�5�j�������U�t}�|�S�)��5��_�+����7���c�����G��{�m��mi�g6����'Z��La��pQ�ɍt��ڀ�p^ҸE�[i��;{�j����4��Ǻzi�b�>��.^�"k�А��)|�!��vknё�hܨ*R+@1f��&P�	t�%�]���NcA7�p���s;,;ʜ���b��]�?.��d�Jʸ��k>�J�Q�E%�r��'T�ҝBR9���k�8fV��d��2D������M��j�rc�ei�d����U�JED�iA\�d6b��*w�ȩ���!����(S���_+�p�oѯStś櫥��kr��n����l%�u)�e�t��`�Oxԧ����rQS#6P���v��"�ݲ(���!�j�
<�����t�ꉛ��z���/���ʧIUCvc�Ok!���/g�;����5�Q��&:gKv��Է*[m�g��ٔ�B�:��S����»k!�N̆�y�.�.]�������<�be�W��e��b�-�s *uk��	�OL���oCR�f��W���V��9P��m�T�P^v��R��ۮ�Jc�)l��u�W����漝(�����X��t-t�/f�1m�S����z-ӎ��}yq�˥q�/5��PW�>�yU�����a�\�K���a����ǵ�+�\�y�'�/�⧋��1Jy�� }�}2��K,q��e�z�r�U���wd��\��hNB�?8�T2�-�?��󛕠��:f���[ľ�����Vr�7w�Gb݅�ξ��T���,��9���ϥ_P�&�u;�b��bY��;9<��pVH�MV�;h�;��=w��u���!����6_Me�U�yTV:�Қ�Pg�ٍNZM��/7j��)�i�ۅ����6���{"oY�k�9��;��wMIR{ӗ��<r��1�\����ߡ�}���ګʅ�rj��ouN=�[:�ꀴZ)A�֢�B�t��A��cK{!���*O�6f�ؽ��L#$S;�N��Q�I����	G'����f�
!9�S1J,N�o3ԛ�P�d�������io]Jv�_�y���ξlm��X��Q6��O���H��`�=0�u�f+��Z�[�j<ӊ�v�mt�>���3��I�������Gv7��J#ϋk��r�o���ci�^o��G1����d�{$>��\��.;�0Kq
p��V׻Ӈ�4���v��xԗY���_'�8������:KaI�P���2��N�f�W����,�75��Yy����v[h�����i���_ ��lA)Mھ3N�1GQ�W��pz�d��{�xך|V�wl�����Ճ�w���RM5�"�k+y�t�6,˼|���9��:¥7�R�贛��%��{]�V�b*d��	�'�j��/S�����o��J�lNB����L�댦�:�mu���`�ֲ�͕��+�����[�v�6.������o��X�����7R��usW^_�9��W�,N�U�ő����,|�r�2�QP�-�=���X�^ؼ��/�K)޽�"m˭:��M�׏�z�X����T3�ݭ��>���X�]�2*��xѸ���Xs����LVJy��FU�\�n�[�纡��u�frWFG�&լw� Jǫ�Q�	ȟ)N�ެ]7�y'�/=mi�@L��eW:9݅�SY׎#kMe�K�+�(3�EG`LV$�N��_'ޱ�vRy�s��}"}����кy㒀�To�S����.͝�%WULÞ��m�Ifs�����m�Nh1�p��䷔N|:m*ng�꺺��M�zS�V�b!B��5��ETȠ�9[]r��3!G6���ҷ���ن���%���:�k������U^J}0#zs��h�汐���r�`�`]N���@�gYtzW+}��� j��?a#Yz=�s"f��v��1�)r7�qّՎsh��*'Aa��鎳P#�͍`�K����J�!�셍��+�KF�%��0K�!�Q�`ʵ�݅W�*�"Bo��ئg��-sI
p�yz�	��S�<k��t+����n�,C��YkE��L�$Q�u@jV�m�I��﷫ٷC{N$jQ���p\�u�8���W`?E̺Kx'�g{�����_:mW�姦�V�	tU����E�����<�ylD�mKxxJYE��Wh�0��W[RX�4�㢏j(�L�Fe�2A0���8�4��F�>s�ycx������W/pR���?X�՘uwj��t��=�^��<S	���ףw��f��;��[���l� �׹�&��N�p�4�ꌃ�����֢��H�6ˇq��}�G���^�`gRA�)>��j�& c�B���,�}.DW�Iׯ�֠*��I������x톇.���{�����!3R���?x-����'<3���
(p�}a�]V���t�����0��6憰�����r֓�ĭ���z���0�cl�ZYʈ�P�]���d�]�0����T�`�[�ɓ� ���W0F�CeA8�C������\�+Un�ѷ��.�{w6]�L�hNV:�bHW� �C�_/S��'�į��X����zq�GJ y�m�����Sc���D�H�yː(JS�wi���E����M샴�y@�� �G�SYn�V�YT��-�\�%*�K����6�[�C0N粺����TXd��oE�Ĳ��[�#n��=
�e��b�Y��-�}E9A0����,��m�)d��8�8e�PS}�`9z�:��*���ʓf�ZHZ:�ݕ�5-��H<�A`V(^��%>LL����NyE�������hA�b˚wwʦ�\�Q�T*�����YRUz/_�SK��6���3k�����S���"����;����s�_6�}Ә�d��DK\�az�RN�0�L@��GȬ��������8^
@zo��KJ:�2�]�G">>�D�����A���<���.�I�#�̮1����\�����G.�H.숶�!J���fw�@�����;�(㩆6o��.P'kGâ�^Z4l;o��R@x��6�e�{�=��,{no�l�(M�b��K}/��ݯ�e�2�@�^��&\J��͇��B�R�LI`ܶ0L��MG+��^t�1����� ه�S�<K��������ժ�sa�1݋�9�.�n]2�Uq4*#�+9��͝H�}GG3/d��h�(�C�'�Z�EKhĴ�,PR�VѲ�iKJ�,+bF�X��m+��TT��Z����*-���(�Zժ
���
!�TDUAE|M9Q)eJ��QbŖ��Z"�cڊ*+-���ҫ�eX��J�b��ƪ0ZYR[j*�cU�Ujj�U���RV�IEr�ej��U�R�Jъ(�F��X�D�1Ke@TAb��F��Q�ke�j���YDCML��3%�UE&YcYRQLj[*9ZY����Ze���(�aX�
,`����R�
�PDKJ��������2ҥh��#�У-��ƊE�Ul5���
T(���J�,Q-ҡFVQ�Ҵ� �hԭ��U�E(���������D�TPR-kkA�UQ#P+*�XUJ�J"Q*�H�TkU�B�QJ%""����cU�mXĶ�k�R�EX��DI�U�ت��*���(営"�%��+~����zĭ��唧Jr��6��v�kɇ��"�t��9sm��,�[p6�Q����Q�6�;���ŦA���q�R7A�6ˈZ'�y�W�qy^�cj<�A��k���Z5��̺gb���\��+9�����rO1�s��iI�-��{0���Ȩo�.��xg-���Wk�ϫ�TwP9,�m��t�st��[x��U��n�q�{f�X+�c�|��]dx�σ�(�)�;ٶx׸u֙L��;�U(�ǳ�[�⛪*�'Dg��oIYL%���Վ��
[�ey'�9l���p� ��ED6���hI�m׊�%uM��Ω��l��gJ�39X�5�'R�km_��������a���s�S��rX��.9��޾EkU����Q��MECah��L7u5�-K͛���A����Y���{~��R���碽��ϖ>�-ݳ���T6��ĥ|���3T+�l^L�YJ}Y-\fʌ�z�b����Z��s�ker�W}�Q�2r�˛R��`고��e�o"p�����sɼ�8���^��E-$�+o�LY��a9��-n�M�!��w���ʇqw�J�^~����F=���}�F�V�.zWޚa�9g��kSKǕ>n��%>t��׽&���/6��-×v��sUӹx]t^PX2����x�d�C�@�`�ƁQ;L�k;��z��7r��v;���7��{}F��Y݊:1�b�V�d�#�)
x7MQn��}�����ov�^RBr�ܺ�|.�.�'q[�	�:�m�<|�L���7�N����Y~��m��)����˩+���ӘS:��QX�ZT,�ð5{�H��3�}��w�f�s�>o-+K�v{5 [���XO:�K��+���'�ᨧ�kҞ�Cq���јp/5"�{ӧ��u�0�����U��Q�K�!v���+��1���-;iF�ʕ�N��T���8I[�9�pU��v&�CDٵ���ӛ��X�V�K]�EN���]�,u��)�����v�
�5�v��n�6�,�/�s�ޅ9��� �jÕ�����p��4c2������{j,�1�H��i�,nz�\g��:����A�*;޻�����=$��a�V�ر��u,�%f����R�nm-<]��ɣun	��RE5.��Z���V�wб�K%��2sÓ�`�`�ΞEM��]�p˅ԩ�uI].WM�mZUx��V�2�[�^m�DT��1S���]�]>�<��)�+�ܚ��s�"��E�"c��NTk��m��c,���}Nn٨9�����_G\�ח*K��^�k�^�Pr�:6k���.��P���I�|�t\62a���X�꺯*y�'��y�T���%�_���u�yN![���{�ylc}���M��Q]��V:�N�k6��ϟM��/y꽅{��*ާ8��O��W�Q�m�6�����^s�0�]��s�=����>������U�e�km�}��ouM\9��!j
3&�i��.H�eN׊�4�η�!Q�E��Z�if�#ϣi�¥��.�9��٧��!�G%�A:�%GO�11�j�'�n��Ӝw�yg-2��m�X�4�p��ZC�=I�o.2OP�lՇSL��yağ2�4}�:���o��=��'���FX�n��L�ZA��8V�z�z{�}�DT�; ��F����;�*k�6���蜔ͅTj�]͑��U8	c"��i���m�T�X��4�{�:�i�]�ս��V�})�7CE�}fn�lCs�Q��nގ����#�J¤��<���"?}�Ƅ!1���R|��a>O?sxJ�xΞsz����ݧP�� �Դ��z���I�3h|��>y�y���E����M�ﳐ�ɿ��gs�N�q�9�@���6~�<a1�s]�<x�����;܄�6ɹ�?h���<��%ABk�q
���Ğ�|���o�}�z�_~\3}�y~߿S�O�=gN�������8��,���d�O�xg2�����$�'�M�$�m��Mv�|�$�w��N�Ӿ�Ԙ����߆��n�=������*N2��P?$�'ɳ	�'��n��8��z��2{g:���g0���	��'Y6��v���'�,�НC�N������.��.��}�[�w��|~�^��>C���1*I��ԕ'̬�'=d���	�SS��|�F�u%|d5�8�bu���#�����({�z4DED�sl���5�?s�����3��m�h,��p'P��s9�d�a���RbT�^�$��~�72����uӳT'&��6��q��Ԃ��Hh���$Ĭ3����|��[�?Z��O�߿=4��	����O�Xw!P�'�,�y�*O4��d�a��+�I�~�O�X�I�O�~|Oڡ8��j��ğ�q'�{��������̹�=���݁�i��w��2LeCG}è,�_s�q�����'zʇyHT�2w��L���]�Nr{�)?>05l>@�OόϝiO-�/������~�w�����i���a�?3�M��Oǖ��N �}I?!�=��:��14~�d�*��i8��T;��O9;��|�is��J�a8�j#�{|��tk���^�����y��O�0:[0����I�&��1��:��'�c'^o	?!�6s�M�OY�9�d�T'|��N�y�'ݰ=d���4o߷���}��[�	�!���l�JFN�s�Og��n8N^y��:�M��J�^K����u�0�+sD���X��rrvu�q�|�R��g[�-9��
�n{����g����8����~*1/����@��n�KR���x\)R��K�Gb����铺����D{�����o�����'�0�O�&ߙ4�e�d�%f��N!<��2q�a���d��7�>I�7��q6�<g9N�ph�xe�������I�3�{�֫����'�ԝ;� z��O^��x����=q&�x���'��N���2OS[��I�hu��,�}���N����8��.~o�-��WG}���><鉦�;���N>0��8�Ԟ>�wvN x�Ǽ��IY<`l9C�VM0���4�ĩY'�u1 �Of���'R�"�b�a�e�u��Z���G�G�x���rAd�O��_�N��y��8��~<�>I��'{d�	��u�IRu ��+'�?!�XCL�M̦2OP�h�z)�zTO�[����\��B8{ޱ���|�Ĭ{���'<����d�M�����g��ԟ<a?��'��O;��d�����%IĆ�B�|��﹭��T�ɸ��E}�n��E�=����蟒x����I�P�'����d�'|�߬�d�o���I��w���'�6���'l�=��B�O����m����߾{���L��{׷/IPP�9g�VO�Xj�=I�O��
I�N��v&�N3yC�N����2q'��xsXC���o�?2m��}�u�d�描Jx������?=��=�#�ӝ��Y'�ny��%AB|ΡY>J��$�'�م��'SF�>jI�h݇�<|di�R~~B���{�S�S�
or_ǕlbW��D�z�z�D'I�i��u�	�4����$��jLJ�|�aY>J�P8��O�O�a8��h�aְ�CSv$�����з�MQǘ�>������,z
1C�ē��0�'�<@�w�
��<Af��$:���3��,'Ro��I�RM�0����6e����wT٫	�O���\������O�]�����u:��\z�T픷����M=�/n�ES:����yA�݈�tC�TN�;��ţ�Q�G*z��|�5��C���K��(��ނj{F�����u����ݳ�\!����ݥh4q�S��s���o�z�S(�}�'�U��^�q{�s^���į�'�?���W�a���I�X{=�0�$��ܚI����!P���w��I�'�{�Si'Rr�$�z=��F<���߯�CE㳮��z{�|�OY=I������ٷ�O̟!�y`x�2m���Y&%a�ϰ�$�9gRq!���*d�+��B��&�����M2]㿽��k_�j�~�z����<�s�^$���Y� h��8���~5Bq��S��&�q����i��ny�u��
�s��$��s�:��VC}��8��V󿟺]�׿�R�w������5j��i��?d���u6}dR~|`j��$�����q��x��ԜI���1��?O7�O�u��y�PXOP�������\h��r�����\H��A�}������ԝ��'��w��ܓL�<���ē��"�o�4�2�2O��a�a4n�3I8������:���޽��J�� aq�X7������G�D91�Ԓ~C��ì�J�o�a�N�z������ORz��|�'��xO\d�'S�Y�&�yg'�SF�8��s5��A�<g�k�
i_kW��t�b�
�
�*��ܓ�>d�V~��q'P��a�m���fd���w�����'��쓬Rz�[�O�9C�Y4��VC�0{��J�}��Y#>�?]��9�����!�
I�_�������'�s�0'u��N�d�a�N�q��}�L��ORw�N�O�Ӛޤ�8�r�Ƀm��6~�v�zT��G��=��I!�d�6LI=C�bAa>|7a�O��5��Jì�|C��2Ad����:�㙇R|�$�ğ�?o�>��*>��ۛ'/>Q���^I�<G��N���%a�AC��>Aa�i������0�$�l5C��I��'�XyC��d��{ܐY:�}��$�#�\|o��~��w�T��Hq�S��N�M��t������-�7|qT���*'D��uoj
֯9*)��e�L�q`�-�n�t\���J�b�2�r�+�(�:����J�=�3΁n��_s�/����A�L�wi�������f�Ym��IN���E}��W�UY�wgyv���Ĝ}d�����!:ϙ=���|������>��!R|��`|���O,��Mn���	�o(u���A���!�#�̱�l9ɑ�<#�%�Vη��@�L9���w��:�d��o�}�OY�M�s��XN��u�T'���!Y>Jɠ�z��o$�'Sl>���4�[3V]F�#c��~��&������<z��܁�I�/�Y6����rN&�=I��7�	�6�{�$�Nw���&���J��VMzLD1���!AJ��"��Rk]�����M�z�����'��I_���Rx��3�~I�I��p�'x����:ͤ�����N��&��,'Rl�ޣ�x�G��\��7������H��=w)>d�'ΓO�=O?P��I�6~�ԕ��l?yN0�Ρ�����Y'�8�����T>I�7;�	����i��ʣ�:��a��s'���{�:_h�����rE���������lՐ�������N!��`~N�m���gLeCP�ܝa�I���o��@辞7�;4}_�N����?z6���!Xxɣ���l��?N~�/�$��E��ha��?>'�Y2C�i�z�������u�� ��V�����g~���؛_*z�@�bvs�|��
C���N2x���y�+5�k�I�O�d��N?$Rm����q�ԟ���m'M���N��2��}�Y�?M&W��8z�y�������=�XO�9��8��l�?$��Ԭ;���2{;��|�4ɹ��'�$�M�R)?>2m72Ì'��~��o���@�a/*6�t|�9��==��?&�8�ɹ���$��7������:�d����ru'Y���u��Ԟ��P=I��>a<`{��'����Lq���4��U+�px�:#m=-.�<O�L}݋�»�1�D�	��X�ަ�"�Z�³����Z(9{�w7H�V;��~���wpU����f�م!
���ڃ0�1w U�9B�y�"���f�����)�u[N{0�v0��Qm�C���ٮ$������x}��������d*q���a�?$�����>a�[�L�Ad����d�T����a�ϰ�m�x�ygY9���p�'Y>}I�d�`z��������^]w�n{ǜ��2��C�O�ɦ!���L�egXO���AI=5�Y:����2'8�<�����ï̓�?s0�'<�����s�]�����}�N�{{F�{�<�y�Dp�p�5�%Ić��䬟0�
�x�I�xe�I�M�Xq���$�+ϼ�T�d�T��� �q����������F�;e.ZH��y�G�L���Oǝ��<}d��|Ԝa8�Ӻ��+�%d���i��'�e�I�La��I��Xq'̬��X��˥� ��l�M��{�(��ޡ�`���>���7�|��c'ܧRz��w���q=dߝ��T��y�d��̇��P�� ��i�������|Ì����7���s��u�}���B��c�>�=�ލ��Y:���<���P�~�<a1�z���O�4���!>M�{��+	�=�ԕ	���B�|�����<�߳_||�����{�@�'=N�I����n��:�a�'Y�8���g2�����?$���M�|�I�o�	�6�}���:��>*�7S�dN�v�s%��" ����#�G��I��Rz��Q��'�����q57a�J��h<�':���g0���	��'Y6����I��'�,�>8��Oe�W���Y��<�E��Ү� ���l�jLJ�j}x�������'��:|5a8��k��|�F�u%|d4y�N0��a�)��I>n���g�n���/k޼�}��2m��:s�
��<Af��	�=dٝލ�N��9��&%I4�$��~�7��d������8��5���N0���^�io߹�|�y[����[�tn�+����)��v�况dn�3������d���Ь^`ӣ�/\����rJ������ۏUo���7��o((��#.k	:��'�c ��mmE��}��=5�}w���j��u�<[_��e5�
ǲ�U�_�z"=�u-J�-Zii�H��"�=�a�N��M��m��,��!P�'�,��a
��MN����N��9�$��I���,�~�52���$��������/�|�|�T���v��D�=�=�<��=C���&2���p�$����u��,�$�OYP��a
��MN��F�M2o��%2Nn�OϏ�;��&/>��3d�t����~��&�Y�P�'�����q�l8�����N ���$����è,�G�a�O��7�����=eC�y�=d���o>cޡB�o��9��L��{���.G����w�"���ì'��y���i�1��:���'�i��/���C�yϲu6�=g�{�Y8�	��d�'G��c�w�ά}Y��n�չ]����BN���q�������N���	���iY�I�Vi���w�4��M��x�Y:���x�Cs�d�m�x�#���oR���V?�V�;�H��`�{�w2q���xw�@��Ԟ����=`o��=q&�x��(OL�M�d�2��C�,�{��N �}�%Iĝa�o�T�N�?_в��ڀ�#�G�x����	����Y>|a?w�q��=~d�;�$��=No����07�2�i��o,���N&��=C���D�{ꟺ{�����'.�\�Ԉ�"�<J��}�T�I�T��d���>�~I:���N���	�K䟟Y>;ܓ�'S}��%IԆ�C�VOXx�}����1.,ï�3����'�@�?Cd�C��SL��C��J���0�'Y9�{d+'k���	�;>�N���	���I?>2l�
�=M���%O1�o������U��˥��A� Xv[�d�6e1��N��a�i�|�:��A��8���9퐬�a�_RLdRz��ě{�I��>w{�NT���jʚ�^��CKp[��p�t"N�Ԭ׼e��i��\/�L\t�ޘ�F��K��������Q�1;w�J�?<�sl"=9\y;��ױ�X��}��P�Iؔ��\�ѕ��gS�!l��~S�:. �?\�C�Ep�܅3/�Y��Υ�)���DG����oC�?z��cߣ��	��|�d���@�ORu��RO�q5��L'��=d�������I���C�Xw���Ơd�����_&�on[�z~�`��zǢ�����M�l;���u�w��PP���!Y>Jɬ�q'�>eN2u<����'�����x_p��<~@����칌�Q}�V��+��X�y�>�l�I��{��6��?��u�l��@�N!��jLJ�j}N���%dє$���SN2z�~��XN!϶�}w���/w0�A좒V�#�i�����$����6Ì���0�'�<@���*d����HuY6gw�XN���oRbT�׌+'��<�'���aی
��)U����zy���{�v}f�RO���$��6���2LJ�^��Xu�s�nM$�
Cs��(|��;�B��������N��^~ԕ+	�������K���w�w=�s�Y>q�d�'~}LB|��zn;2~d���<gY6��޲LJ����$�s'Rq!���T8��V���4G�>���^\Iߏז��2~��G�zt<��W�I׌�O�y2Ì�����Bq��x�d�N0����d���gXOP�6}�Ad���d�+�D�X0*l������bk0��ѣ���N�T�2h�ܓL���I_�'Sg�E'�����$�����l8�h�<M2u'x�������I��������}y���mP�(@��z>�M�ߤ�v�Ũ�%j�����G�M԰5��Ω��d��OC�t�D9u���ͪ�m�ڛ�s�;ty}�����̆�֗��l���Q�r���Χh_8@99�/w&�F��e�L拗]?��0p���ͱ��p����	���7��X��xX��R�l�D��n7o.e�t1�똂�y��	C{b����t�-�e���e,g������w;0L�	.Cz
ӻ�,��u��Щ��4S��Z����]N�!t��qpX�)���տ\؆+���d���]�í|5m
��Z�YJ[�۔
����G�|8]M�pZƇJ˓nK��gv�T���⽣q��9�ͤ��)�.�U�9�`���1r�r����-X��Q)�H�yթO��4K����j��Рv���{0�xUfб��UX��M� �2"
<�<�v�7��Z��R�f��v�������&�ź2�L�Od�vCg��4�6�K�Y7+�3feΦ�jz�;�voM��n��jH�Q�*[n�Y��錮��ߐ���O���4�����(ts�W��D�+���z%n7�xJ�C"�]�`g<��9Y�7VM^��Y���� ������Pq��Wn^�?	|M���I��W\��7u8@K�be@�شk�SFjǛX
6S�Μά<��
��h���jQ�G+����K��7�!���
����J�u�F��^ao���n7@�@��x�K6ţ����]�w&{No׏g5%��=��q�����V��="��O$��oN�%��tD�����p���+�]�ۙ`��A��+vvi˜v�>����O���G{�r]m���d��J��.k��܋!Q�M=�;-뛝�N��q#���T]д��v����\�
�x8>R_ʳ���,�F!s=QR�&q��-����\f�x'�x�ޤ\ۊ�:Rg�fq��f�<}�Ѭ))K��{��CH+`��['�8K6���;+"}��݂��,�\�	 �wjr<`��w��]���d^�������N�{L�����mn�In�t9�)���x2��"��L�/q7y�i=����F2ͼ��b<�j��:ѷ}з�1��R���io*�m�j����(�=�����v���dW�����,J�)�`�s �%YW��][�Iq=�)������c�xM��r�o�����/s�Au�Ԯ���|�]⦎����bb�;q���.����&��;6H��8マe=)U\2o_CY��긲�pY�+)ΰ����hwLɝH��z3���ͤ�g�B��fV�%Ŋ`��p����6������=/���)��/��͛�ե����4�R:��cK�)�iT�zq۩�g\ev����mc�$T�\#�o!������	JcGo
x��gd�V��Wy��f�e�'u�I�� 2��Sk��y�t����U��k�0Jx�e�84=(� ��c����E����y@s^t�|��ŋ��+Z�h(�XȉUmaTV҂Ȉ�Kh���
[J��$���d+YP��K�V�z˕EKVB�1s[K-�TUF �"�U�
�m�6#"�Q�`��ȱDDuh��(���*.4�1�(,�*
Q�
%��Z��UaDW-E&�QCMU��¡DU%H�fb3
PPPm�l��*�YZ��PX�TP[k�Db�eJ�i������%��*�c�"��V"��YZ��̶��T�S��DU�UX*�:�+`����ũm5cR�`���b(�%Ab�j�Dŵc(��
"���J�ʕ�F(,@P-*�2�A�m�Q�EW-ƭhȪ�D`�6®�Q��TLHڊ���mUD�ň��)PYZ��3�"�,\�y��߳=��헃��&C;�Rr��Ƃ���z4�[�E�Z��F�Ϻ�*mU�{��
X�'S��e)�;GU_W�U������o����\��1s�x�q��[i�睽���HNt�ݛ�=+^C����]P��R��hTv�E��!K�p�Yq�;6᷎��sD��\;¯��d��cO?��.:����b��I��Q��VԽ�X�Z�ǯ���@��ؒ���^����)�˙~����*ǎ'\�Ѻ�r��\K���Nk���t"y�k���U�<+*RDEga;V2o�Kx�t�Խ��7�dP|Y���6��[�s��.nz�wL��7��靆b龼���[�l��iى�8Jː����'r���Y��N�l��}@{d��'�7��*<�.����'����EZ��Q���j���9��N�"땵p���d.�6�5��!v$j��c������Q�:���ɯO9��t�"/��������e�r~��s�
:u���O��l]L������pniF���Dv�ڼq��2il]Gq���e���s�'�A/( �:_+ݕ|�Y��ޔ��̳z������8��BQb���Gx�"�Ŏf�|�xy�'��;ݮ����ݘ)Uw�ވ�DDE�[Д5���~Ln
hcu/!X�]rW^\�2�\nK�8�s�B�֔�ʵՏ�a��2��T7�E�2^��GX�]��fM-P"���T�����q��QY����6�4*_1��7���j=�+VR��#����<��n�aQ�x�TeZ��6!kB��{��v��ې��X&Q����8�\�4��J���LW��W�*�Mbz�6+$�O�W���<�u��<���;~�+��)D�q����)�U����ռ�t��ݾiog���UaT�rUA:�ң�)1>�	z����e,)������b�7�������fߣ^$�68v�'Uz\���ɨX��j�=���{�|7��q�����Ǧ�u�f���fz���}�\Y���]O3Ϲ�[�j%⹶��Pv�C�U:5WP��i�*���QeV���co�u�q{$7�ǽĨ��XF��A��"���3��y���{��71���C��*h��kU���,q�CB�O�u�.��:,���"ܮ�z�N�`����]��lU�r�ESy�tɁګk�4�J��G����3���͍�����s�LV���gaX�����Vzc0�j��
�z��א����48a{��i���>��GU�t������}F�<M�z�w��tcUl�d-���7��5^_:�y�{{ݔ��;<M:LobʛL9���6�9���*��f�5:�Jn۞�;0��H�6���۔�F�E42[�w�[����]y>�oێx̋�.��m�Y[����c�QP�-�ه�SQ�-F�*/n��k�j�ܘ�}q4�Ւ�ظo����Pћ�;L�zɅ2�ֻ�q;��K�3/�v-lVg�k�m)�d��TvU���[kZ���IˬUs�����r��5�QչYxUz��X3����T^7�P���J��5�u�@�|{�b�g'�n��������6,��tE(3����LCm�.�9 1�k�`����{�� wQ-T�@z�y��$��U�)r B(r+��Bu�������'ܞ��	N�;�%\A�aB�C�j:�_K΋kV��c�wJ�UbVCH���Z�*��q����(��Αv�t�k�7D��坄_ϫC�r�/����z=��3ս+Z���6�t����\6�󧘦��.�
�u�	���9�
��n�5��i������y�p�ؽQM����׃�A��HV�N����Uwb�k{Q+@�r�Tð5v�/Rz�9`z�0��~���co�"��l#$dX�c�TΧ���qI�>i����]����i��k����W�u�÷��Y�b�l!�����l��_t)�n�UD��,��}g���oN\�yUΤ�'ޘE>,�]���B���nf[at�E�[T�\�e+e⠝_z,]�n��G����Â�7��79�����T�R{}<��Uy�t�]��M
{-�9��.��#DLjmE*u��ܯSm0������}6�[��}��^�i��a8튆�L7t�X�s����f�KBH�a\��O9��W��5�=��j*��k7���f��ɋ�����!�fP��c�V�%�6�]o�5��rSڴps���Z��恄��'#/��B�L������_w�3lY{�{Q�8��u�[,^!�D��6N�ʝ�)U�s5T�G������_(��z�>��ٙ�g�f��q���h�]Mu���˓���N;�~�~sM�_{i�x>���V<���{{5�k�� *u��+%��>I�+/ҌC�L�<���}�ꮝ[^ZШy����W���������k*���q�m�噧ȭ��<��ν��.94*7���wo���mi�~9�(�/v��F�{i>��Ox��JY%g��ʠ�|_e�i��y��W��fB����7�4��*lf2���.&`HW�'P��"�\c�ͨ�K2;sr�'��@�k�czWN�٠��ܯ�D�K����{Y~�P�)=k:d�0�#�����Mg-2���z�uy���ýڰ�U�
�>�Ğ�;�u���e�޾o9�F�T�~􃝍�]��,�ŏ�XA�u�t5+R܃j��9)���X���F��wR�R��:3�G�����u�>�!·[%��i�)����Q��۵�rrscnx�:ũ����v�}�%��m¤r[�H:U�����z-����Ϸf����a�.]��(�Z��H�(Iv��]�v����e���d�5��*�J6��"��B9r�F��"#��{�}�.�?��1{��F�%�9�삲yk�x�{X/�ږ:�LB�Aav��N�=̩Sa㋤��
t_{5=�*ڰ�{Iz���[[���r\O3^�T��(	hh�A�sQ+f.�����z�^�mXr�/�v�m]�8mb}϶ET>oDK�%��yFn&���G�ߛ��B�R�b�˂�X���=K��	�������±n���0W^\�.Qg��	���ؓ<�6�%4֊��82��7k�C&��{�Z�������\��v�2)�U�5o.__�%EDgb�Gs���M
yoN	7o��Տg�Q"��2el�^�B-�Jmn{�~/��t����QQ�j�:խ���+ݗZ�j����(���Z\ɝ~��/z��4���T^&;+��7����vn6`H8c���ڞ�8v��vb���m��up����XH,I��|�1˔3m)������4U�y���ٶ�fX4{?/Q����Qw)�<��S}A�#���Km�=j��}7bXd��m�n&����=��"�(I:�J�|5�o���C�wu�R��:@�.Jy��F��u�[
w&V�0T��|2�hC��?�}�����lUNJ^�ӫ�y��>[���ߕXQï �']DJ��LbP�h[x�')֐��j4'c���,�׉_��t8w�VA:�V^]��ݪ�}r�ީ���O�{���S�5���:1���*�����J���f��Iۢ��^@-Ӱ��k�{ѹ��b��+$wc{K[�(7|]��ºߤ1R"}�,Q�vr��}{<v6��G��.Kt��WjC�X��;���J�CwKl�!�<V�x��c�0�>�e�{�oy��
C�
���]�ZS�M���Jy^.�'Ds�QM���0��iC� u�M[����,6e�V��R��9��.�ߡ"cP�\�v�H�j��-;=m*�Z6ۍ���%rsP�(l+�hd�t��ty��M��¨�wen����ۂ��U��3%f�7�A�rj����*d��F<�&,�l�;m8o�-��VL�ڇ���M|om�Cg!�� ����5X�*�9�f'�*��nW"��*(�;��>��
�K�=��7WP��V��BF�{�$v+�Q�y�C}PqZ:=XTb�L�5v96pѾ���YϽ�{���VU����GE�^_�iLV:W�*+������kv�T�j���Ԧge�R���\N����U�7ε��{ך�bs'y���z׺�1�����~��9�ݓw���߶����G����QW��4����]�u9�ʷP-�V$�/C���og�ǌ�ү�G��Σ�(���4����Y:���~hr�	����i�ez��q��������7j.T�M8�N�9�;B�7��	��F8���^sA�9F'&o�o�]y��M�rv����ý��P�Ԟ���^�����n�K�9����oiy$SΠ����I�ӧaG��]������٭GS��*��ל�i�{���c�װU�;�X�]]*�u�rW��O]E��ZTf���T����]0.;�0K��(>,�3y��_S�.�)ʔ�5�y�,�u���o��犃Cۭ��Q���X�}k��H��:�ݰ@|6�J5�����N��F�N��c��s�`�������{��A���s��lc$�C/v{/���R]6N�6c�Ŋ� �,�J66����¾���z'�����i���>xþ���9�ٔ��*z�]��Q��m�&�X�\C^ʮf��h�35��O�)�6'�6�Rİ9Z5�='��B�l�kv��K)t�D�O��ձ�W�����Bq�
!��=;�&��x^�p����M�`*�rV�\󚬵�����Py5eML9T'�)v6�aA�1���u�U��0y�_���J�]g=/-�}P��6ڡPZ}¼�-{[9�.>���������+-��e�7^K�9�ťjT7Wɸ�ZШy����SW�Yx]t^Ux��� ��t᩽�9����9Eer��Yɠ����W���mmi�6���4FD��$[q�>���讋�J/��r������;{�6��蜧��-(fO8��nP|2)D�c=��I�B���k'�������6���]�&)�|��+��e�;��[�ƾ�&̕ ʷ�n]Z�Ta3����ʓf��um�����{Q�5��e�w��5�Q���ۼŢ���4B��Z��p�Y."��c�G���c+�,�,��5*��:rU���D{�w��Ϛ�1YrY^i�ƍ��?��5����=2�T������m��w)5"���\�N�,�����,��(��	>�R����=����`Վ��+�T�����8sOy]t��} �{0��C��~� �޺�Xڹ��7)��{�}���u���2k���Ӧ�)�T%a�c��p��앙9��=.�7z9k��H9�ה9���Y>����*�H�]��qP��YV,���S2i�X������"�T�"x��[�犀���p1��ye)��e7��P����?kk-�۹��m��I�4��3/.�w��\s���^*�¢�uq2.�Bts+��|�^"gCOQ�(C�U	�&�)�XFq�t�/_���NP�^Շ���3��_W$���-+Lи���+	֨��9�A�DY��u�D�;6d!
�\�U�t�s٦�|��m���K[�b��g�/:�N�t؏�,�"�q۪����1q�[�h�m��hI*yŇn�ǡ�b5t��t"��%Q��O��Eu����]+���>,*�u��Nݝ��Q���xWd�K�5�f�1�닚ߠ���n,V]���駲���]D�qY}�-�*ݹ̅�Mjf���]3g*�71"��ӠG�ʎ1�W�ٮ�L�+�<��S+����)�pŲ�#���6&��r�v���R�&��8	{�G�Č4�e�
�2<,�؝��$xS؂']� ��ʽ����w�甹4�ǔ9f��E�K������3���3|�箯�: �ki��v!�r��ID�LV���uo<K�M1��7�Z���]skq�0(4�-�Wz`g�;B��<�j��z�m@���,Ț��3�X�-pJ�[* �s`��<��V_d��q3�JU�9�i��ȳ���Ŷ]^S�67��;z�^|�#}����ηt%
�{&^ď?s����ff�/Q3{��Цt�@�vr��B��tnJlJ�M�XlM�3���}5 uxU�Y9���9e��T/[�2�&F[[B��>TC�g�ׁ[�Z<�fu�֙[P����Jnц�[�Ӫ<ܘ4�7)^7��0!�"*����t�T+�Ua��^��i
�\7���k*8����9���V����&w {�W{l>�H(a]�㷻���bt6B��U&h�Êf�Z�H��]u�F�n��c��R�g�pN-������������(\+N�h����I?T��,�sT�ڠDZ8��VA��grRL�R�����ћW�J�M�	�G��A%�5nd�뤉)u�k�vc�ʉ��쾃��$�x��S��Ŏ*����������v0KX�91N�wY�ʦ��Pm�]�{�EV���c-���7��מ�3bo��^[7Ό�����iAқ���{[*�j�_͂\�7�P0�go��.�R��R�:���íP�m��˘I���3�s�Ӏ�}��jۃ����0w/�'�)��	}�.3���Z��QnF��b�/uD��$.q���
�Xi��ޣ��?s1�=�^)���J�l+��'4�Ku�8e腚������=����8rZ*�l/���q٨��:�mMh����W�Gn{<���0���y��r�����T�H9����"�C��e2�����_1$1�m�9Ҏ�Y�*�V�����#�qV�9Z���__#s�Qu��_g���gXtמ�Y��8&d�O�@s���Ǹ9YD�fRq)�FHi8t4���[�]AL��8Z�R�5���77cUݜ���\�7I��ь�s!쾍䍬�|�5/n��A�t�`.��G��D�x������[&7�=�T�;c�5lR��s0���;��;�"����0u�6s�+��>�Ĭ��B��
���n�;y����t%��oM���$I7��>K����� |H$�N"@D���TFE��b")m�[E�AT�,�FE*��iQH�m�)Z#@V"��!m��+uJ�r�`֋1�(�r�QaX���,��k�AJ�(Q?�Ve�b��f��)iUR��+
��\�T� �4�PF*�����1b��R�EC �q�KedPPPP�,Q-b��I�T����G�YY`�[*ЫiQ�-�DE�Kj �R"�ȵ�]ڐDU�5�]R�\�V�ʣҢ�����X��T��dU����b֊�Ub����ڲ1��UjJ�fe
�+PF%��U��Ȫ���Delkwj�"��[b��r�"�\e�X(EdTk]����AuJ�##]���E"�"
?Q A�����y�d�ny��Ok��{
�����8��w�����R�i��F���ˏ���WZVܫ5;�U��\�ޏ{��D�.^�e��+�(~��A���p.5N���qQ��"S��x�xpo�g]
"v��u�CEk�w�\��4"+f\���t�^�".#'Cd\m�|�m������︉n�b�l�;*�[�Ke)�E�jt��V҇őZ#ʮ�W�:�����M�n�e:��GA];�;���׸�h^!�����z�n^`���Ք�hZ�X����P=5ǐ����go�7k��j8QS�x?)u.1�-=����y�1~(Js;E�c�dD���W���gy���D.�hز\=��8�zP�x����ט��SID:�`���O<#W��zp}�5%̨�覯�b��s�89B�f�A�v*6�]�(iݡY�\���n��R\�.�X��k((e����Px��]}6� ���1r���xD�3�U��Y���fO=3i��4�6��Z��֡>v�Vz9��G��������:En�K:��-9�b��R��@��m��ᦒ=��\^(�6��z���ءn�U�]\���75�M��ǳq-SK�9�^X���#�����"pZy>x��[j@����P>��c7E��M�F>Al�u$=:u�O)��|�S����b�NT��-��O���J��;MeM�a�k_uE�7L�Q�$��_}U�VE�������w�똴��9r��3	����L�>ff�WC�����.������>�0��xHz�юȀ������ظ�a���wa��4Ex!f����@&ݝ7ӭ��̾���pLx;��w���q$�%,D�T�krQظn��^�X�,����͘��T�<�$0���Mp����L�V��{�h�S�N��C{ָ�}Ĳ���j&"���k�6l�*d�P{�p�@�;ϯ."h!X]6=�4�����Q����`@��CvA�/^:��,ÓvJ{��X�*��^P�9�B��5_+z��ڨ����5�mA� ��ؔ�E#�Mv�殒.z���\�9^�k���)���S��|7h9��y�uI����:���W�T���¡�#q�h�<�tI�憮�m]�2}Ii�v�N�9��v����
��Y��!3Q)ݱ�.���Pc{[�����M�u�n��5�j:��� �����6�J��WK W�$���R��L8NV������[P|6��i�v==b���Ǘ'6�\=xɰ50o�w���6y�9`�j���<�T�L����ѣ�X�B_�|ߥL僂X5|��;��{�y��i�˼+��Z>��L��wս��i=2���N>�	ފ� f���k�#�4�w��j�;��U}���Q�e�a�0,��l��s�A\���)�s-�
͢Qi�D�)�	ﶱ�1H|�Ɣ����Ҧ����@'`2{K�3�]J��˕������t�N�gN��O���>K4^�zՍ��^l�@���	v�����W/Ⱦ��2xdk��\�~���]Ak�5�ԟ,��<5���.��a�|R$�#��P�
�Yx��U�MV]5�8(�����XĽֈW�(^,r�߆vC�*`�r,IRik8R����ػEzn��C�>!��h?���C����ꡇD��x`��iK{)VfV�Q��eJ̞�1	4I~NHxn%O�X�40*��;6/��뤭�a�]�9�J$h/�7V�/�;j��9K6���e�<���((
��O�ܦ�5P��_پh��J{�9AX���b���]z�M��
nH�^�;�}��u-�a���)U=T��rYQ5:Ь����ڷ�o��p�����:�b/԰N�E|&�೏��; t}�a.96�!��j�4}s�u�d,�B�л�k��iڴ�{�`��[g(�u��WS��l�l,]��WF��"�]��I@�/t��ve뻷>̈́Zkj�}F���N�CPd�ѳPM�H�fopGbR����V2���KZ��O�����-�����}�T{��ɞ���=����;EE��c6������o8I��,X�,{e��L޳�mTX�i�3}�_�x�8�z_�f��|t�޻��v=�t\��K����Az�b�n��V�r^.Gov���������t��>^�X�x �
�<��d"�i�&{H��3�7O�����-L����>���Vw�������$>��&�?�t�R�.�n�=ޙ|e]�zڙ�y�Į�ޫLׇO��0��Ы��[�C��P�B�ٜ�Õk��YQ�9�H��IcB�/�pVl��BIo�	��8�*�A�ta���������k�	a�An{U��E�W"Y���q(u��"����0��`���:�m.U{�Oz�(��	�q*�=)�Gib�*���X��uG|�
b��i[�����=�ul�%�gF�`�\&5���/Ӌ��x���iqzȪܳNȸ����w�e!Cgw���9	uK˄w_7���q8�a��*儡��7�ܺ�]YE���s�W�q�kx��גA����^'�˖B��~����*ţ�em����at2��M�e뒆���0fv<{8�6:�e�9�S�u����s�*���m�ܽ)p�Yɪ�3r�B����ꕥgYvTԳ���r�|W������������mb�+���,L��B��ƚV\<����z`��CZ��vi�+�dBz�w�h��,.*�'$5ڎJ�TD6�	�1�~WK���.��cٷNjoK�qF9�J�9K�%��'��W7$Vpk��$5ږN�vĬ6aϹB4^W����k2��䔄�b}�A��q���4����@p�4�zY=�͊b��Ʌ�3��)�ؗRov$qP4+ٚ(;ڦl�Q��*7�J{8�)�S*��4�vҽ{4�"��f.F]�Ɲ(�;��B�f����6���2#B�h���V2.*^�s�$^ďil���[�ܝ�����B0Ϫ�5�頠_�g�N�=�v#�1R
W)t=�'�����K�`�.7S;�3�r3W�>��i����R�-��y|䘵l��{͙u�=jR8�u:��|X�.��c�Z{a�1ݐ�0�ٝ��L��gL:�á��W>��V�>j�;��B�|X�.��q>ͿF���X)��r9��<���֮�6�#��wH�v�^�,��Q�Y�fS����HG��G�()��=�;8��M{����{F9�p9at�\�S*lww����>]�%�(2u(n�ٱkNŲ���I��5�ۭ�.�����V����d��Wc�y?W�W�WΣ]Q�����Z~��:�S"L��&^�!����mW	�_��b�����(R��&k
�eQod��,��� ��Lڪ��1�*���C1�׭�ț�:�r�u���R����'�^O:j(��{�����񋄺T��	�°�Y�-����s[g9�J7�ذ�L�o�:�}%�6�Pp�I��&%��co��Ǻ�v�]k��J������Awx"����iN�ۗvO3"��ʺSS���sYs�U���̷�8�f���IF��D��Sl�B�X\*��
uK�0��H��x�N7��X� ާOD�%���~�����W��$�uB*������-����u2ƍss"�J
�YR�]��[���8��3�MA�w��i�|3|�2w�ҞU(O㄰����j�ƿY�ܔ���p��L�b�b8e�4�1}yuI���0n�U�Ϋ�����-s5��VCu��T�#UN`-��6�+�ۓe���cB��F�d���l�Q��"f��A��T7�6�<�|�!��]6�HAw�2��H�-�cW>�J.���omr4��Ǒ�Ws0��t#
��G�q0�N|��=�Bgo��k�ZCG]%�9�k�J�};Y�l�ѧ���8���4��5�B()�ٸH���Hs��=�K�Uw*}h�_x�44Z֬�{�7W��\��X~j����,�Rƫc��9)���tԝ�w�3��V� �fVR܃�fv��gk���M{q�ʩ�mM�45Wo�S �;��?eݛ�=m'��S�^��l?R�,�t5)ݱ���i�e7���Ub�b�jc/�V{5'�܇ɣ�<���$�K��Mu	6������Иz_j��R�a���7�K��{��3���J�. �NḞ���.d"Z$veb�DZ}�2�u�Mݝ���Yn�vr�k��X7�l<�J�8�J$���z]ɞ
�*U.\�(�b,���K%Ɗ��ޭ]o��	p۴$]7�4^���g��l�@����.�A��(m�gE:�ܠ��M�S�|\�ƽ�5���,��n��(Wd*1�`:��7���'�ט�3��z|��z��[�y@��w��/H�2����gk-[.%�S�$%�r��p�P9����NꨳW%*��J��q�<2�ڽC��ϫ�`~=v<rJV�2K��نa����=z�f��h;�v�f�-���Y�ۮ �jKA����36෎��8�=ۥ�(=��{������_[JV���
/#�Ǉ���V�Jr�r�il�u�+,n��9J�M��U���l�(1ݗp7���J�g8t��%N��z=�����OC�1�?>;l���Dv�
O��X��V/٪���,0�����	��m�-_�>�"�}�_I�Q��wB�$��u�.xf�7/�yj��̼�4��Zٞ�!s�bqQ��	@K�� W��"1׽���݌�}Kp���n7�OMJ;/r̄�5�gtIt�&�v�e��\w�c�v#�x����@M��g>�,�ږ�'��<盝�Z���P{�|ʼ0�*�����.���宑7�Hwo�GO	켩Z)���pk|}$~�����R��T63n�9�����v,�`��rW=.֎�|;��gJ
[�4�{LH��5ũi`�6������/x��Z< uX�	k�\,E�ӕ�Q�v8��N�n�x��:�����E�y�u��P2�S$\-�8划�Oy[0�#�����\}�m��Wv��{hC�]��Zhx؅%TI��qT�p�Q.�-V���'[z��"�`:�Q���/�����>m�إ�a,��du��|��3uF]��cn�=���1���,s�.�#�)y2[w=�d�@�s�o-�z�!�T�AHmk�1yqD��5�S��o/bbLm���q��a�7K��Zǵ���5��=���]���M��sޒY��� �y�o�W4�E�|�,��ވ�C���yV��t�}���衛�L7�G�F�򜂸�{C]	2x�l�ϭ�9Q���cr����g�A>��!�K~XuܻV��Cc#�-B.��Ń�����Z�+	����=���d��>���D���Q��>
���o�:���o-QhC���r�ĉm-f֪v#C��q�9O:���J���O.`&HD�t*QLud�}Mq8���)L~�z�T��͵Yy��'1��r}(KL��E�b��z�&���(�y�7���W���CZ�d��]����۔�oi��ڑN
�ÿ��NHk��;bU��M���x]#8���{��M�&ë��G�4k�����q&�m�h_���T6%i-I�+�s��%�E��c���dmz�����D����:*T�9�h�f��'�DĬu�����������A̂������z�wzT�-��Yu�XY��YP�ͻ�{km@sz��n�霖	���0`��/C��]�jVbS�C��]��Z��SĲ�X=ynW��/�x�����{0S�D����f�m��o�n�e��t/�,�gk��9������.y|bQ���2��3�)�\3�f�O�*'�Z�bo�"�թI�b��2�m��Վ���'V�
��5�`Le*���*��5!j-܃��&�dGuaK䳹�{�9����{׃+Q���MM���t��{��}Zw҅��ȳ�yUH�����]J�u;��L=.J[~�ݍ��Y�xt�چ	��u1C��	��ӂ3W�)z�:1W�B��A��[�a|���禧 ?>��� ʗŎ�Q����i퇔�vC���(J~��.�bf���v#���g��=��ym*����%�o�����#��}�z�C"<�?��� ��xn�go'�B��a^-�T�g�TC��eXhtSV�b�k�E�9�q0����W��m���{$d[���fʒP(s70Puj�"��<믦���`���g�ر�.`Ύ�Ӟ���O��S���l�D��@gOPtb�-R���'�xU�=��*4�_EEtg����F�;�v�`"X�a)�M+�ښ�߲Y,u�7��ÊB�`�MVi�˧؂�á����^��\�w*f��H���ʺSS��a:�,:����W[��~Z'�Z��y�H�Sl�d@UKK`��jv����uyZ: |���z�U;4��6���q��}d��F�V�o��g:[��{��sHz({�Y��gE;�_� �[�F��9s��
�k$��r����,���7�&��&�=���o[gv{���{<級��-q�rNw��Ƀ*m�w��}](��&.>��E�N�C6X?\�*-�0��ƠƹI%��펜&��iQ��ƖV�l�Px4_:�^"�I�lԮ�%!J^Z��djV4,���۾e�vyn_����ً:�3��Q���m��f�D�R��;�h�j�]�RT��2�h�\8�prgA���������B�r����\�0��b_<�gT��Y�}c�����!|���5vP����|�٠�����q�ك���4w�+��Cs�����	!�̌�C`�kH��@�¨_]d������L�Q��n�g�4�zt�Xso����!��3-$z��FF3SI܈9ʞ�$�j&����]j���ô�e�gG*�s��BM�*�{�>P9�|�Vny㈿r���f��؇Y��f������f��5�N�x�b:��8̠��(ff��U=PX{�V݌k���1��{
9�g� ַu�����RF1��� �Rz�t��?L/C����Á(g��k���`�^��\P\�Y��45�,[B*��FYs��u)jɾ�9ҷ��F�uc{�(@+V쨸���K��b��C�1V9����ƄN�\7k5��UwL�.�)K�3�M8x��_8��1�w�/k{��ʝ*�aB��3��e�w1�7Z7�I:�9Ww%p�o�	���;6\�b%N{�������f�|g�4J��Q�0`3���;�Hj���޳S�
�{��;��5O>S(Z�%�(.izY�u�{/���!6�l2�C\΢5� A���$�rę�Ϊ��Q�*�\�}J��*�����}tkSe��`j.���^#��/v�x�2�(B�jIE��A�-���w�hC�CUt9G앵��p�Fy�ɛ���w�iN�ˣ?������n�9�f��<���V�|�W��ʰ���gzm���0v;��>�jL�ʍ���.��B�G����Jj+����n>]�B��J��H�@ݭ���6�}��)𢣐���o��9�s%@b���<��xO����]�N���+S�zs�<|�p�{�农����~ꂫl�2�ٯ�a�ؚ��c�U�F��^b�(f�Qܢ���Z�`8��2�45$��g{�dRӌ�#�p_��ۏnb��2�3!�7.�L2v��9�OwBo�ӏ�|R�}-���J��zrqМ��北@K�?;������ˢ3�h|]�� k�Xkq�S�U:�uO9�0����`~�9zbΆL��:��u�*�]nv;>g����;�_�{4�E��]v3���!��V�:I:�PZ(�� �,D�Ԩ"MP�nڢ���Yf0�(�(���PU(�Tb�
�J��X�DE�""��V*�1������Օ��D˧�EQ�j�72b
[A�-��%�QE�e��U�8��6��b"�b�ĕb(��1AQ��رTTDĢ�PR�DX�E��J�F"�q**������2�5*J6�*4�m��j(�EU4�QTU�Ld�"(��bj�����(b���(�Q"��Aј�*0U`������ �%B��DU�U`�dc��EV0R"�B#��[s!��FZJA�,�D5lDD���U��H���X�b*�U�ب��+"�DWT+�b�%�����3N���z��]֍�+�%���9�cu)�o�������2��*CgD��|.ye~�c c�Y���y�""=�Pn*r�͈�?�J�n(��ٸ'���%�I��WK�d��F�%be5��Y�`s&�C�ܓ�ې"Ą:�\T�,9%���&�8��N�@v�GOF�xd�_f��e^%�'�>˺Y'��4׊�^\M&�]�27f��kc�O�6U���M*@Kn���Oq�5��ѹG�暂�8V�F�FIlκ+��2bm`�ٽ2Z�-*[C�ú��!H����؎M���S/�w�>~j�ߕ�;��P�����\�!���V��uN��\eO�T�����o]1��a����mM�45if�;/|W�K�3C���.N
�-+ g
n���(��\Jwldt�Zs̠��<�=�����Z��x�l;�^6B�����b����ߩ���`
�d��8�g�7��'KHܗ5I4vC��\f�jt�X�.B������v�y1.�\%�6%��Hp�L,7�U�3r�q��K���T
�C>�+ڳ�6TGJ$���idjU.%���i�[�dk6M������j�h^���V;�SKۚG8'�j�s`��621�h�3A�N�߆�k�$�I�Vٯ!��եZ��^&��V�2��$��R��˭cٶ���D�����g��[Ok���dT��eXoU�qN��U��Uvg �95�B/�'@;{\$tR|�E����E��3"����TA�z�szi�h�L�z��"v{��Lj�5����fX��٪sd+я]�@�Q#@
�����)�b�4r]�w��9p�hR���x���[~���qL'o�����Em����I�i@*���dC����Mmx�9w,k�U.�G#MOB���쫚���i�}U
�ޝ����tI�RGa,���Je��k�U�͍��xH�V���5��]z�2f�$@���Ԝ5���R�'�P�3���7)�)S/-AV<�c�&�k�Jy�~��逴v������椌n梳��]l�c���tq_�o��v�u�?9����QVy��;���^ZՑl�ZM�TEy���4m�Ia;y�G޹m^$1��C$�+�Z��6�q�-���C"ߏ@���䘛�Ž�f��f��C�E�X.G�FV�O�S�\��S�����Eʆ�n�8<������]�h]%Lt�q�ѨX�&̓�c��␐&��祵һk%��'�_�Kʺ.�l�)�P��j�D��&L��;�ڊ̯d^剔�����?I�O�\��/�z�d�	7��JSѺ��񜙳]��,��t8VwbN����B֐We��}���f���ѕ�7��������n��=��Nb�*,զ��뤰m�Qh.�0>^�U�G��	��;��r�ӫD�.X� �F7{�fv�${K�:5U�p�eD����끨�P+�d�Z%�O���m���[���Ĉ�"}+w���m�Wk�8��!�M ��ȡ��]�Y��9�a�cw�q����Z��D��P[��Qn�C�/�����9�h����'�)޼���+P��/[ȡ��UC�K�Lb(<�@0��+�qNc{'<خ/>��b<sf$����,�v|���-�u˱4a^<m!��:�[�-w.���C���s*�R�ڻs/��p���w}��"�8]t`W�����9���-�8��L��K���ŞK�߲�63b��w�;q�K؅r�,.�K��Bx�	���;��9�*&�����)!�:ފ�o2�kǕ7�!2Ϥ�-0j(F�b�t��oi]u1�����<8=�y��(D��s�����̄�,+sH��+�smT�"��>b������8��6�4J��vv��CNkT����a��a̼�.©S�Lu�����<Ս���8r��)�i�{���#�流�񬟍��=�pvwyA׊^��	Z�`��9�wQfP�rG4qu��;��z+��^lHH>�i�I�ٟ�}��%l��f���0X���q&��m��P)�+I�j��hHca�1،o"�;j�{J�䠪H�ײ�7r�&}Hh���|��/��>\$�4Y,�C����3���)��b,4E�@<l�\�^��SNIp1��Tn'H���/&��;yN�v��1���P�X��Spm5nϴ�j�ϭNyt�z�iq���/�u��e�A�JunRޒ�+Dc�� b޷}�^Oq������u��7񂰯����LJ�Z���;�d��)Fx��p��r�y�.7S;�&{�NFj�`��4��\VN�"w���������ЇiS�{�Pf��R��c!K��q��3�xI��#�Q�|�3rx�ޭ��-7�Q�&a�J��PXd�Gd�Q�b��E�bԺ�u���;�<(+OfCvs7�2EXN��F�g���~���L��y1��Y9���*��Tn���{���P��G0���y�&�H�Ҹ��P\e�3��$��]}6�}f` ��
�����Wu�x��i�VA��A�����W�����&�Q:=ǓM֢D"���l��=6Yq�Q���+�k�m	�zJK�"S�m^��݉�:�AbG\�t��ue<�`�H�����z�oT���ҺAlw[�u�0$v�V;u�4�3��_V�t�I\���ӱ?S��(�1�u!�ݚ!=Ch��Z���O�Z�X)�<���&�.C��Ռ�G\����y2��f���%��Pp�I���T����'e˻�剮��s}oI�ӑ��yW���]��
]�5�K�3e݀�1N��Ɋd�~�u��������Mԇ4W�t���ձ_�v�j�՝��T�� g��vpDG��z�}d�EAV:�
 j�V��V8����/����HO��]����P]��fMn)3_�kJ}S�.�$1�r�R��ڰ�6v�Τ����OD,ҳ+.(�ңU���S�t��rx�>˺$�w�3Mx����<^�}��!��X}���;�:!X%��qK F�u�硩�7�k�^�>��5��K��Ь�m�����9|绖³�l���9�5kVE�yM�S���.U������qޣz��sG���q��9p��B&��@���ʞz�Yѐ+M�t�nC�Ѻs��:+ BB�7+���}�O0�b���X���V�u��T)|���a�4F�ʲ�^���?]_���~��'c�e��
����67X�MnicJ/"V�v���B��/�����+��5�J��Lu
kd��x�o.{Y;yyњ
]7����(��DG�ZV��{<|�7�?)(�ZPi.��J�>U v�=�B5)ݱ��t��(1�8��B�7�hd�a��
|�K,}�y�P��E�'B��Ip���S���DH��k���}4�6.��@��{�{�Q��yoϚ�B%˰b�Է�*U�E0�)�s-+�D��g:�厝V�s�V�rM�
����`{V�4�T x��a�|��.���d{�4��b� ��MM��~�;LFf�׭��]g�pP���H�K�g�`�]�G�T�b�;7�����[�ʊbй��֏S|�,e�Od[�,: 1�� �ˉ�UQQ��h���-�D ��̄/f�_��u`O��
^���sg�Tr�S0!
Nb/4ٶ���k����CY��$jJM+��:W�v�B�:��S�MA�7J_��(F� ���9n��T��7�V�O�X�`��p�S-$�E��R�b�������E�� O��{�������h�nz�v�i����`���b�ق{�޴�88)���ߛ��2����'g�
�s��ű����mbw�L��3巪�U�{M$�g;�_-�==C���e<�u<x[]·��K�i���� �}�+|��)�d����%�7�Jw��Z�!2鮅>�ͥu���gM��7Վ��}�/�M�ѕ�z==O"OWt��ģ�&�A����Br&B���N�}&U�yK��o�ĩc6f����`f&��]�4�5s��k�'�J���h�ݳ��ǵ,��K�{t��u5�δ�{ͺ>��w��e�@��꼈Xͻ|v���Ǣ�z��l�Kݾ-��,��.��{�>9��c�i�E=w�	q�wIxi.����/P߰�N���yK��]$y$|���`y'=Z�ɳ�-����S �փ�4�_�A�u}l�T�Kd\d�`
�T�Y����ɾ�8X
�-T�F��M���	�Ӟ�y�엗��AK�F�����jPO��"�;���&-�m�����-i>�鈥/�#-l�Dk�[Ӑcv�
�
08��%t��o�ȳ2�ˊ�2��;��gf���~����`:�CL9�q��]���G�KH�i�`��%v�MY=U�;��#���FĈ�+��ʖҰ�q��ɇ�G�G �C_�<�J|��C��l]&��ǜ�T�&�I�`�,�Ae�������UܻV�چ�G�Gʄe���3J�o���u=}�0lR3.��ۙ���̌�1���6잗l����d��J��P7����;.�7[܋�F����{��]�ʰ뛑Sp��L�A�\��3^�K`\����	��z?���y�:ì^t�))hCxW�=��ކ��[Σ
��炸��h�r[U�P\E[48��^N�9�_[[�5~��V��M��K;�ۗf$J.�˸�W���BrB&�\���oßب��'�Z��ps�y뭷|��f�ʛ��3T�c�tz����B{��i!�SK~��e��,dܽfS#��-�R���{޵���wV3��+*�
�� 6
�6�\Ȇ�&#S��g�v����TGU
F&�����;�e�=�l���`g�
V��-p7��jY��GlJ�f�iӦ�M��̕m�Ҕ��[�$�:�v(��N��&75�i7�*&��P�� Z���PNݔ���=;%�b�X����=��ځ޷��լ����h����5���V��B_s�6��^O�A޵%2�Uz)�7���5Z��<�ˤ/L�62t6AO��2��NΒ�}1�~7K�7>���&6�OShKk�-G��
l�XW��ůJ�:��8k7��y�.*�@qg�;R��N�;Pɲ�u��~=� �����������۳�Cj�KB�>��՘{(m�ؚ$f�F�4&H<��^�a@�e��z��JjD�P�K�/���I�P�w'��^)�c!ݧ˕���a#�a�.�:�[CL�nu�<�,\L[�{Y��z�"W���/v��L.���BMw�2;�W�����=��G��^b��A�+Θ>��<���\�|X�.���Zyܱ���0�*�_9�O�I�����Ln���f_Ȫ�G�k���d�Q�@!ބ_.��s\O�{di�]�u����:,8�����.F�\\YUL̺�\�dtS�l�����r���[#ݷ�oϵQ�Q�Bc���]��H��;��:��
����z�Mq���䘮t���μ(Ԓw�`-��Ţ!֬l�GX��@��rL���B��\��C�z�EP�:E��Ў��</}*�;�=��O�I���%�,�E��sl E4Z3O(�Cf���Z.����j�o����jN���odw�� )vt`l֑o��O��
Ǻ��2{��;�1�G9��l��Ȫ�UGq��,['Nƹb���Y~��T�Q�jv��[��r��A*�x��+F��X��|ճc�R�'y�H��xRu=w(Vܕۮ���ή���I9����W{b����e�(BF�J�w��g�u���4H����m��W�%n�&J�y�l�o�خ[�b�B^p��|���S�:���g&��d��#Vr�{SO��M��pP�q��Y{ݦ>��[ܾ��%ݾT���8��L'���,u/�U�դ U<��sT_��_��E�L{�<����z�0��興��BsQ��ʋ��:��ٴp���=�vĲl�y�]����	���]r��@]fԸ���W�H��0'΀��T�P���r��ժ���8X�4�s9Nڪ�w8�36��/���?�+�����6��=�ֵd\=����e��w�/����q4��������r��X�U�� G���<L�8��o]1�wZ7O�zV��D���]T�����Զ�%�삂�ʥU،>6�����߆r�q�ˊ-����m��N3:뇱��x.r,��Z$�^@s����D��Db�>�ۿk�n/jZ���+htuv��k�CQȆX��`3��;��!o��[�bZ^�������I0�˵�O^��E�:Q2���b�>��l�׃�ltTD$Ĵ��L��~O:=�9^�Z�S�l;gJ�"߽��uoo��O��XTk^Qq����G@S�T���V$��W�G܎N�N�q~����iQb��	����h�D7�2�7.�/[�,: 0����o��ZNIFKHM��߸�Uz1f$YviЩ́\��S��ۊ����9�]��cF��kP\m*1n)ݮ:T���6淋�c�y��xehO<�vhD�V`=z�Sޘ�y����]k�^��ʑ�)�(Q��>��{˥m�{ÖG��Nwr�[]�m��#:��e��;������Qwu}g�&Y�z��g=�s^��{��TE��7̼�m��Ӡ҈�t*�}�Pi��]�M�Ԭ��Á�wn�/{:�v��b�=������*ۜ�V���hF(H�P���r.�A
�M�Z3E�f�f�n7����i�i�I��2K�g�ɨ,�gr���ce�.н�8���Y�\�w��F��9��M��z��c�Z^��	hR�ۀ�S�}���D�D�eM&/�5��W�0�Zݾ�U�Qxs>��vs���cp�х�������&�y`�z�{ة�,��k��2��0{;Kl��E{���s���Z�X"xQ u*�؟d��݃�2���W>�������j�E9�%��*�Ҽ�[�>M�U҆�4eXuT�a�7�\Ӭy��-;5Д�ۖ��A�⬭td�{�oW����̧�
6��x|�ź�Xu��%�=��"���wb�ts,���c+�w��k\�j����{/;��*��*�Hw��Rϰ��;�j�`���w�RWZgLW�����oe��r�k|^�'ZLt�Gչr�I��^J)v�*�v0��[� 욆s��HGD�2.��9_wɻUy���K�Mق���yQ�2�,����.b��i�v�& l^"u��v����o�>�"��ݰ����ICf�SŎ�"����5S$�!�N:x��}w�B�^P�\���Y��֬��X�]���+WVJ�f,�F��ۗU�a܌aJy~g�߽^rZ�c�X;��*g�����
�]
Φ�+�B1+r�t�)%(P|UՊޗԝ��V_�vIj�p�аh�1cղ������M��7d[䀥�,m�U�&�
���=�u�Ώ9��ޝ��E�*�9j�?��#��#�ę�{�WWN�Q�܈6��j#�0�92�u�22R�E�GS�X�&c�t��ﱍ���~������띰�z�f=���/��q���A� �滽}�K8|}x��@\��`[Lqe(޽�ww��O�qdh4��VD7Tȥ�񧓞�4ܨ;Y��I��,��ER�q�3h�]��ϳC�/���/$U�����WK[��5�P� SQ��滝~�ʟ��xaΏH^�xM�'����eP3�wp���X�U"�s�����ԏ1s��#��M�R�ܛ�h���x�,;�Mj��GC��?����EB���L�x͘[�Y��N2H�����Z��Oyڳ��zbpv�1V���n�%q��2g�n	�����|h�!
Tl�ED`��`���V5,��X*��_mDE5kKj�J����QDAF��(��J�
*0U�cR&R��"��T�����A��QIc#0�f&5E�\��V(�""�ƌS+�Z�1DQ��-�`���UV �Dk
+UQLj��m�h�*�J�\�TB��UĦSN"*":��0dQUUDb��+X���Ȉ�օd�[`�-*V8��8�
�����1�H(�DQF(���Z �����(ɖܵ��
&���V�T�A9f8��T,G�l[[YF*!�P�����h���`�eQḬ̃JY-H��Z�r�E0��m��YF�r���V�AF�����)m�|�K�L��z���{�;��0ڤ�����{���x3�G?_"7ܓ����;�J[*�˝�@�85��ʤ���ڝ<Ui�ޏq}�q�6�0�N�&�#N�P����|�'����h�~b��G9Vv��Y��c$�13�����ǩz�𿡲H_tG�iA\���A��Gk���R��l��m���5|[��յ�E��9T>7�w��wD��9#�ߥ��P�40*�gf��9���n�ˬB��KI�%��;F�@�N@��M��^o.���I�%�^\3q�)_y��f���^���͇�h���$��E^�
�6% *�2�ʸ��6at��H,��5Wt.���]����OU8n��3�J��흈�^=�N�F�&��1=�p0PD)IY�\��DT�\�zkı��&�����7�v�����f�pt?���oۮ�$E���$�wq��4Hpԡ"��;��w�4���b�e��:!Ez2�9��w��S���j=*on�X��ζ[Z'���+�N���#c�Qh.�S��x�x�w�	��qY�*�Wڀ���\,�.��&{N<uñ^^���"p�I�.�]p5*�χ	�����z�h�m��MD�F_t�oFo/?Yw��=ź�]���n�]%E�r����K����1`�v�	v�΋�e�Z�}l��x:�'����΀�4�oڋ���-z2\I��8Ƕ� �R�k�\��#!���Ss�2b�V��މ�]<����O_>|%2n1�Q�/�B2��k���������x֘.��,�/.�\Y���N<�kg��C,�{C��P��И{��^�Q���ֆ�+6W=��I_h��n ����������x�P\�u4�r�7�0�ld}�r�~�H+�/���{��'xͤ��v�E8a�\#���t��!�W�w*"�+�Eb�{yR������N�³p�
c]I��<J�c�0��]vQ��yF_�9cSO7b��*��i����7%H���%LB��1`�qP����
NHD�x*ڦ:�`]�AM��1B<�����A�|^��YLw����(KL�B/�,X�e����j.{��]�Gy(�`��Xd]`�/O�ws0w������FJ�DC��M��ɭ�
�oW��~�.qQ�}H�u����~�;���l�~��M�ZM�TF�b�F�9]�:�ͬkJ�#�E�uGd�D�;6d!{v��Ӵb�]F�}�*&��T)W�>��k�OݰU���g`�:��bP�wa�<0����^Ya@oδiA�Ͼ����'7L8�<hl��bL�˼���"��}��OQ
S��ތ���o�p��2B�rQ�b�C��Q�y"ߡ���1���� S�^뗶�El.̥z#3:z��m`�,�Y�:رb�G�Y�z�o����i�(դi�=u~����!�}�lP�'g%5g-I��Lx�ϱz�0��]X��{�oS�!\��M��#6a���`�~/ �vF�m�(`�&6�z�Xf�ci�v|6���>�͹�8T\id��7���/�p.#6S&�n�j]P��:���{��K��y����ҲH�2x% QQ����.�890�zal����6�b��P��X����=�}�m�9���J�*\�`��|���EW
)J��<J�Fo�V�,"���HɈg�f�t�-\�i��[�,��X)����*C�ʪfe���W���6Q�N�-�۬�0G16+8�돴�t`���#	��Wg�d� �̘=�UAS��������=�Wؤ�S�f_�xUJo�غ!ֶ"Gh��@��	��\%�P{�ڧ�������id����ke�'�צ`��x��&c7��}$��Z��s�����EQ��f��,�G�R�v��c4���;�.��y4�̕U�{�R�?\����(nk>/���ׅ%���nu��ћ$��T����ߍ��]���������\<Z�Q�2kM<�{Y�5XmT��8b���ޘ�fO�} �QE�������zx�7��t׷�{{ ����:3��ZE�:cn]�=	k�<i^�EL�4��Z=�4��v�B��_���{ΐlV�vT��6&��)"�Y�HN4����,ܭ����+F�!�P��k����
�t����wM{��	�#Y�0>��<3���װғZ2KGM��P]LG��LT��SPy������g��f k)�����>X
�[}��B�I�#��5'�몠��/�@�5O�/�AJv&��R�,.�z���|p,3�=���;��5���X�S�m�V/�ה9�{Rv�r{AXLwy��0E|��R�mY�7/ǰ⳧+��H߼�Se}=pM��.Uj�s�Z����J)1z�:�NƬ��S��X#qYu�_U+:0&V�����3�ν��z�.�Fs}��dϪ�k�ϊc7ꭵ0UC�X�(U��R�
�:"�S'l��;�Ю���ų*�E7��~m�v/�Q�KC��\<��ʮ� ��! ]������	.Q��(�=xs�qm��m�b��&�e��?�4=<�=���MPR�9��%>��9�D'�@��t�_0{U�t�X���wV|2vmZ+p򃐻9O&.,�b`��)Z�Ʃ��N��V$X)�2�л�O����ݕ�Η���~va_�t�渔5��Th�'p��b]"�K��ļТ��X�v��9{ؑ�Px��z��+�>��l�׃�ltTD:�0Iz���%�#gI�T��=E���xn�b35����qI���XTk^Qq��5��ԿJyY�iܿi�!�>K9u���uu�P��xBr�%kG��c!㧆���pqH�=��Ne������%���d؎�&��]�C����y1��vx>u��1]��Y�9(3)N�/p�ٓq���,�L�
�*m$Xr��(+�
�o�Tʵ�S�MA��7*f&����5�h�ŕ7p�LŇɣ�JS���ς�i'/��Ȥ��C��.�e���wt�ʮ-����D�]%mC`��ΔH�lIK�Ğ̇�eX�a,�T)�����n3�\�������f��k����a��bP��#)�����8aI�u��2�s����F�a��ࢬ����P�,s8���	�Y���5DE{�c�/'���t�|vZ9�^V��Y
yf�[�����j�98}T�N{�l��ܢ,�^���8�r3��9�[&�wxg6�d�"��`�Ii����6-v񉊈n�;��v��٦�o"��Laݐ�F��dw��S���o;�ʝ�"1�X��ޗ2gb�ع��:Fjd���N�i�^�P`�ev[���87�NT$�Q���{gU7��������p�P��YyR�ٻ��M���ˀ������/m��T:�R���t�b�eF�ǉo1�ugWf����R����A\`>>�*�_97��fH�щ��( ���[����Zr	�Ӟ�>���}$4}�ρ�IHkj�K�����'`?[����M�B)}p���c5ĭ��1�p����c��%��Om����~0����ʻ� Ϯ.%�v�^Fw�:�6�d�٪�V�{j�J�x帼���3$�`Q�	��E:�W*����P{��`xf�v���]8�ۖ����xg�RrLšz����U��9(�p�8*��C���&�r�. ��ݷ�zr��t����]]2�ys��;����-})rWU��<-�hl�F�l�_J��SRe��SOR�Z)d��s�o�y��ᒦ!Gʘ���=��ґ䮼�F��qU���Nw��',2���W$���&�h=����%���qwz7p����u�����Oɽ�:���y�ou��'��UP��]��O+�n���L *�e]Χ��d�����>�|�wJ��(w�\9&�2<��pCK��0�	��qw�,`[W!ߢS�=�j�<�8�<>�oJ���Wp�}(KL�P�Rň:�$<7�4���S��LT����9�.~��&���FmME�ʲ°����a�}v+�?��1�u�etL��dm��D��JS��]���/_���`�`=�� �\�!�Ԣ�LY�?]@�_���n�!�a=�"�N#�j�����o��^�����:��)��G�	���Ә�9���n>��N�������1LN!�߁�٫)ځ޷�쭝��E�RMMγy[G7][��A��t�����Nם�0��(?��ջ2�U�ME��Yn
<�<�V��
��U�:���Y���֌r�f|�����0M�Z'������-��dZ��BT�P8봌����{3���\:H���P/ٲ�7�H;T���XaD�q��'��3�oc�\q{i�NuW�|Ԣ�{�аPj�@B��8�A�A�/J�����΀x�%.��4O�n6�b�(m�gY��*�S���\ �9،0��,C����?1�VvA����v���6CgI�V�}���/���3*{���:�~�<bDoL̿�(���z�>z��ڲ-���ZNwQ��v�P)3s��Z�[�3�Z��N���V��.��J��e`^IO�5t<닕�ar�=0���Dr���v.𵒯�E�.V�Z�gfV����u�VbeW���!�@��6�����+�S��0�zmQ�ț�o$\�[|���IK:��/�}�P�/����14bG��L�t����;]\6o����U���m%z�mh�����e�o�qB:�S��]�ۦ�L��\������2���E���ӱ��;�PVz9��G�D�a�.��/�``"_ޖ"��ɋYS[�`o����q>��x���eD�����������=S�|5�_��1�Yٍ���X�:�@p~
�-��j=%i꺨\k���{��t��:A��~5��d��E���U���}�2��,1���1�S����u� �5���/n����w��K�߸�d���4�;�k��z��Idh�u,\,���(d:�]J��o�� VZ�Ī$�H�X2J!5RM{[��P�B�^Nq'!�<_]UY%B��_ک��{�^*�]J��gݼ̄��3vi�,-��`N)`�n�h9Oq���\U��,uݎ*E�De�7[��ѕ=º�ഞx�]��E+�ݝ�R�A��˓�[�K9�}��[m(z�s�J�W`|���u`ܜ�f���d���%ev���9��w7H�Ǚ:V.g8�]0�6���i�y.�6qK*��h�צ�r���Ι�������W4�<y���P�3B2Ke3c�=�8O>~�#k��6UO\b[��<K�w�<���)֏V�R�����Z][�)>nP�<}]��NJ3�`&V�\'d,hNXq���ᢰ-kZ�;V"ۺѺq���Ƭi;%����-��oQg��tFnd]NԄ��r�F����-9���y��V/�E�����Ip����O���ٵ:��P2���i��j�6�NB5��w�]-9�%���:�׉�w�\�Wg���eÕaq���K���泷� �|�����,�'����(�P�6
z���J�!���0f+��S�.�H��8��Eʳ�]1�Hk���H��^PXTj5�ՙ����]z{���@�|F�A-��/-�B���L�tC|�,c�O�lH�X��n�uOjw9L|� 1�\�<�'�q�B��x�u`O���K�Rc�7VLW��}�ns>�+w�6h4��c8�8����$�]�x��Ⱥ�\�Wg�p�L��^i=��%0�f�<f��=�� ��,a������g�EO���v�R���+Ϊ���/\��V��dty�Fr�J�$�Qoqɒ �{����{�w��&��3|�^t����$��������8�tT򥆮��Ɠ�;kqkCJ�e���E�]��DB�y֮ն��j�����U/�ɣ�m�>7�)�.�]�Ga������k�����1K�X�GN����0���Ӑ#`W����˸y��Ib���6�=���Q�gT�z/��
L��¬Do%Q[�d�B4L�MΤ}rz�Y�����0����}������b�������w�{B�c^�18�����ѱ�Ց~g�Oγ(Vof�޼^��EN|�}0c�_!��g�~5���6J��]F3q8:8��,�UW�n�R�t(�O��A#�T{�76�y���%�����zߨ^*:�,m#Z[*9'c��ڒ�0o�]%s��m>S ��h0�3w�t,.��9[��ݾ��XBC3w��sФ��[�����Wt��a3�q��W���!���S&9��jy��#��nT	�l�H��['�����e�����Z����f��R����n�Xߪ��婡q���;Rf5L�6ԢV�����׭�haԂ����訩��T���&���f��.:ܾ��9bz�Wr[�ir|�Y��q�����%ŕ{(7c�k�uhU|۠�TyO��箨43���T��9�ڱ!�Nu�a���i�tBt��^�2󶶛�U^��Y7f��d��)�E���v���f�����c�u��X���v���z��w'n��Rʭ��[�|���W�A��mX�Ⴗ�gC�����i��D�%�U��BJ
mܻ�*d�=.�;k�2h�t#�gwq��-��v��裑B��p��l�6=�u@��r[]��T�ȋ�fX�����L�nd��]i��}/6��"�~||�}<w��Jg��<5k�Y1�[8��ʼX�3�@y�%��A����+s
]R�'s�D�N9��̮��A
X�I�&L�[�O�8,3ub�/@D�(�oV'WGX�IP�ie�ņX��zؽ�[�:ںh֌iyv4Nu}�<d��5�<Z�A��$4w��h��Q��ꋝ��zB\��z�L����F�zz�"7jW����"˙&I��ܝ�3������+ܡL�<x��f_Sw�($r���l��l��yn[�la}�u�@2�5݌'ʥ%�a��<��pc���T:'�H���~�k��N�]V�&q������ǁu�h*yϔ��v���y�Mj�ў���p��/t�����[�}�{�#D2�vI�j�H�oo�:�+ξ[P��sl��͙C{��r��{���6s���,�ݱ rn�Dd�ʇ:��i^�d��}V�cQ�����vfR�ϞI�9�m�"R��,���)��+V�y,'�!Y �%l�7��MMzx�ɇ!���ua&%�OG�|7��mTB�l8������Z�����є� �u�IC�U����³|��1���g?bCy4��C�u�����n�C�Vb�bdKu-&�=o�n���9�;�f� �\���j���ȷ�V ���Z�3���"�K��sHv�D��Q��%�2/:�q؊�8E6���[۟&ଟ<I�uޱr}��������|�m��:�(D[���d�Q�#!7��qS�g���pWE%t��h�z޺��:��|�x��zeE�3v�N�D�d�O;���U�;�a�i;�����Je"%2�@u�Jb����#�
׵�-�@�(�FY�W�uj�]��=ݜhCI�����;�E���t
��I+�HHq+�]U�.c�έ3������]SZ����]�J�a��$����5&[K�m%�!�)��J���27����s�沸]=��z��|�R�_F39��ܗ!H�3�k��S�BMp���?)E��/
Π�����=��vjv7��:�t��2m�u�7>:�[4�ǲ݄d\�����;�'"p.)_3��m>\�j=V������ڂ�
 
�>�[2ك*E��V�HQ��X�XT\�2��S��[IX��2�$�E�̪�e�UT�W���q0XŒ��eh�b�Z��ҭUEX��`ڤJYZ�Ĭ�E�XQR,hUc+4�#lU*J*-a�1!�h��AQ��E\aQ��aR(�媪�iU��c��1k1��V�����R��D��b����R�QA�*5�YF�X[d�T��c��DX�9��+
%`����3�AUV�Z#[��RҡB�Q2�-.5�bc�JԨ�T��*���PDF�-Ȣ�Y\T1��X
����-���T�Ŋ�X��U��Z�J����AJ����r�����߼׷[�ӡ;�<��]�;�g^wb��֔��4H���B�Uzg*}Bv,�"����ݩ�������F�w�b9��imq��Ȗ���r�5��߁�.3|6a0���(�ǔ㧫�={���v�A�T/�#��6M��ȃş|���Hr��4���{;K;v���V��k�^�FI;(��PE��;��i`�/]р�(��c�����l�����W��ͣ��:u�QJfk��s�o�y�Ӗ�ىN]��&��4O"!.���(���g>xx�y��qU��P'j��ئ��ʇ���~�����P�;��i!�����)E�@ɥ��R6+�|PY2�Y�,w��ښ�U!�VXW�"�%i�ѕƳ��ֽ��{1*��|�	��?$y��|a��C�yx��u�Z�$VD��A�*�%bw5�2E��:#Y�!�DY�Q�;&�%͙^���3��h�R~�d�N�2=6���K�u����v���i�P/��CM��#E>κ�XU"�P(<�ʹB�j�p�k��U�Ý�ج��zv^��_/pX��L�m��<Nx=:)�u��;%�����g-2�vr��a�E�`䋮�1�HRr/������O~,��Ae�>�p����c4�l���@��٥��QB�~�]���{���ڒ�P�w&����vG1B�v��Yy�$'o{:^�͎�������V+c�Wu���%3)ks,f��1-,nt�,O���u3�f���4ȸ�Й�X��P��BۜPϦɍ����x��V҇����ظI[ۨ�Zz�V��r!�#����}4͔ɿm��S�������:�'���Ytd���9u���KC0<�y�� ׅU��8��X6�Q��a1a��نL��{���~S����YHwgטC�lL�~�1�
��L�IE�`!�z�<:�PhP�B�����A�j�9�}���:�L_�����2I���Duz&g�W��ᣓmY�{$�X���D.v�9B�lq��χ�15�JG���3q0P`�^N܂���}�w�oU?3���eɵ�2>�m�n-�{(��阁��&Mu��S4��9: �y�7�=��C\LN�\�]z�`�<�a������84e�w³��b�����8ne�V�z3 A��J�-��
����:Z�r���f`�E���5�+�J뽢�ga�����;�rWf�|f"EԙW�)��P�oC�nN��1#}�m��a�N�Ze�i=g~ ^�Hy3�b9l��S��2](��[,��P��E�5�Ζ��t����{�[�-�sv�!��k����K�����a2�y�w�ژ�-���	��;학/�2��@B�֙���s��h'�Μ��j��陵o�����Hf+�qޮA�k��?&&��A�ؗwa��8Y��Z0o�B��۩u�O���hݬ̖�����䖓q$�JX�n�@�䣰ܑ�C��/�r���,O�g$��+˳!w��������v�Τ��N*'P�TBs��9�Õ�pv���X	�,�ޞn�>w���	���B��Lh_<R���"�U`��v� ��wKAƧ��j��I�y7J���.�������<t:���-��[7�٠��6�̌Z���a(�!���F�˝�k�.ޙ2��?5b`�ub�5]!�n��=��;jfv�k�`��JL|�'4���#|&^���6���ém(�T:�@iq�A���0�Y�1Q�j}Y�z?v�t��{v�B�KN2��-�m��x'�o�hp�K����j�9��n���ҧ�R#, ����!�o�{(<3Ke�nf9�t��Y���j��؆g\R�zN�.`�+�k�����*�H��4;�܉�3��P��0l��=�EB�4!�!sb�7��lMUU������g���ɦl	9�t+�}��9ޕ �O�á���w��a�}�SU�n'K3�R�}����ԃ�JfH��ƭfO���dp�k��g^�*���oN˶tk8�Qu�s���Us��-C�sR��v�����c;�},�N@�	�v�&XrT�7��a�R�K����&w�&4xu�{6J����f��oOm.G#y�`C�]�g�&9T]ug|S�5o�֏W��cX���(dL�6^��rkl۷L]�1�x�6��&�u��P豔;q����{��zL��L���[=i�����(^)��c;!Â��XI��W�|*Y�\��]cYJ9��ҋ����i�l��r^;����R��Ib5�0\8�ZJ�r�~YR�zӡ�Bx�.S����Y��+�͋�j�&���be@؄��ܜ4�]��(��4�5/ M�sԦ/��(��J
ߙyk�(`�9�H��`'�U�@~�P ���6�U�s]��is'*)�Q���;��܊�"}[1H�B��O�3�,g?v�н��b�.Uk�ifd�����{{qB�eC�C5:&�e'~4��n��:̫�-�x�;qg�v��1@�z��j�A��ڤM�q�ݾuÃ�E�x���!��҃Iy*ͻ����w6���D������� \�o}}Y���C7n[�	�u�����v8B#J9�k]��h�>��Vg�QP�.�갤��Q� ���Gt�#���`ҕ����;����Ǳwl��K�:�����0rv�C��DM�a=�����x���SҊ��:�hۧw�)�MC�Lw��PE�A�)��:�A�ھ�
�X<�w�F��Z\�o����C�N� �<�yU�Ȅ]-0�gp�x�*����D�вu
y,��r��y�c�Ů[+nQr�O���E��-�~�LE)}p�kh{`��B}�^�>W�lQ�˵���(�^��V�F4Uo���C���+Aa�k���t)}h1�&�)��s��mf�Y�-=���$1PxO@�%��D>V.]���Z}ˌݖL>��H�+1�I�����GM�qNc�'!8�-̴x����.D:XAz�t�=f��@�d��:��8X�5��ip-��U*�(��S�
�'%S,r&�!B�V��t��S�	[�N+��\�����s�2���5"�˳r�*wSa9!}��q�̭
�(�ݬ5�g�8r4��t0�|媥YL,�j��s�@�X��u$���њ\�����Y�$�p��My-�����a��:����і|%�'^�d�l�=�vZ�r�m�q#�A�c8d�j��ѣYL��l�v^-�(N�������3.�9��gb"�`Ҫ�b�0���ԇ@����,��bv!�w*���!H��đ����}���:.��l�`���Nn7s^��j�b�n�3�w6�+wf�ړ5��B���e��]u.��G�u���-yᴊ��*ˏ}な�u�"G*H�(u�����Y��I�ɉ�%�#�!��7�;&�J�9P˧V�f�g����Ng�i��r�I��YV�ҀŎW��4>��,E�^�r��٩35u�(ҧ3�fRl���)���Y�+m@s���-�,n{�rY6�ɢ�e��SpkV���j�e�+	�B�9£Zx�2P�S����"�'Cd\m��]���m�(d�1�1n�/kǽ����/L��]�I{�p�5"Ǹ�Sg�a�U6o��c6S'jP|�ݍ�uLX�.7\�,��
'[��ۥ�~]�ټ��4��Ԏ���!����,�PF��R��a�7���ne>�
��3in-���㚥��Sή�c�P�6�KY��*�SR�s0x�]��	|ǃ��@�K�=���۞�����r9�'���C`�%eD��wS":��G�s����-H�X/��"��"+�n���#�����Mb��T�����v��V���S�����7&K����F^���{��۫^j����Ů!��fȁv��e�w}�W���T^='y�(���$����ɳ�"�]���$���h��؍Y�SE��襓][J[��GU��{��j륐��i��:dކ̔���ԍ�1�5�T��;1^<�=��di���/u����KV�$u��3>1y��l�7珃�d�*�CG��D�s�0QS�t���C�G����R��gi
�l��|�F3�����݋��s��N)���h.;�Q(q��k{���2�e�gB�:m.���o*�M󚼲џ\�wva<p��NR`�}���u8���/��:C2�Fi�1��峗���,�6c�u]�"Cb���D��g��(!f�%u7xL[�ʤR>��l����6^s��V��Ϥ���*W�3��)rрIh��X�9S��@��8���g:{��hՠ^e^��篈��L[Q��9����T������:NT#J�����Xݠj�a�=�u��X����e��T��W"�����V=�	"����q��'s��\�Q)^�.AQ/2�>R�g]A��q����3c�|�W����kVCir��{\�}�j+kt�,?W�r��L�"3������[��|�Pz鞦	�ǝyX�G*ົ��\%A,�/i�\{��"��k�V����8�n�p�#5�k\�1��i��P�� f��SE���w%�U	��W��e�s������J�<AΎ��ǲ���Y�j��b�ԗ]�2Mu�y�x���]ӱm$pk}�����"{���QQ��yo@�!fw��խ0�]�&˄o��Ӻ��g4�n%���/%ߩR|�PS��*��㓳;9ҵ"8I��%�h�z[�c:]-, �jyl{nX���ۙ�H�L�r+�F���Y��d�����w�x�*7$���R��L;�]-9�P�8���s��;�T\NMgX�M�m�'�9�0g�Pj�	���"h5,�DXΏ³�}C�O]x9��f�d�o|���Q�^��Ȥ=D�e&3�fx9*J.VR����!���#���Li���[���v�v;��XC�}�����K�D}�-�ゝO,�t�ul9�E��9�r�o��v��鼰�OY�n�����;G) !��&5��0�/�t��Yur�z��[�4�.X3l,
pBa�U��r��dZ�,_�`�pE�#_9I�u\C�dq�P;,c��B�_%垞L�(��5}j��	T0�JV�2K�0\8�I[��öi?g
WO{�)l�IA΍W(�ؼ�RMqa��ʁ�ܑ�ܜ4�]�޵���mp
eT��F���'����]T�j����{%dd.ڑ�K�)S��lř[�v�{jg�zh�ܿ_�ےq����Ѵ\��;��;�魁���"�����koOu��'���zy����)c�m.��s������9�Gg�֮Ma&Ǻ������)S/-AV<����{�mE^D
�Ġnn�)��xӖ�kH��N��c8j_R�&���
T�S����3���p$�J�����	^.�\#���dDTǎ��`�R��3S&ǓV�T^�B�h���Wo9�{j�-��j��#ch���NQ/.xn�u8W��2�d=��w2��^�,ka!�<���K__͜c��u���J�̩��`� �.J���k{��~�t�چ��N��
/�9�x���rP-�ke"/'C VT�G��.�.���a3�s��ò^^��+���욓���X�R�Mu2�@]����R%�����OU;hxl����p��*�q^sW::j�y���q��)
T6U@Y���v��n�&p�cL7��rq���^K9镚q+zr#��=�KH�YL�I��˰�SKN"��Y����V�n6㮷)>y�T���\��9���q(w;���b��&�!�0pf�p��5&���sJ V��VP���ȋ���m(z�&�U:X�P���:��]�=��F��b�᭻��~���ӘsR��ܜ`
��*0�-�;H��hȴ홖���������<��	>��x%֓;XaND�q���O6�Ӟ�G���܄jC
;`������β��ia[�r-ܱW�we+�:�'%S,r"cm��]�]����5�<Us1�!`1�K&�zX[Ӿ�:6����9�r�ċ�.�Ļ��~O.`] �p�/n�f��J���O��(#���4G���a����p��Wp�J�ʄIj�g��1ɝ�+si�H`�夅�4�����s�z`�CRګ�����N�y8@�)d:V>lۗ������j�E^�lC�
��z��J�2�Y,vW��LB5R5�+���M�J5��Rv {	~j��sb����GdԞ;UXx,��j��~��;g���R��s�-�ɪ�%���,!�}Y)�uп@�t�9@��g.0IЇԫ��5K��z��Z��B�T��qQ��"S��x�N�}�t.=�;%V�*n��e�mnz9)~�<:�.��2ȳ���`mL��[MS�ҢOq7��v��E��8��2ft8ܧK�y2,�<�.�V1՞ ��D�r�v�ݍ�0��Ǡ=)*�g!�c�kx����ש�WR��s}���{�������N
=���<�O��Rf�d��'���&�ӎ�$ѯp��oV�w6���;5��A�tW�O�2�4���T�V�41n�$ִR�S�mko b`D��3�V�}�8ty�W���`_K�tx��m�X�,6���e�ZΙp{����qeҬ��#��6��(A�oV�5zn������i��<_N�$Ε)U�5.�ξN]� �k;��I�@�j�Vpu��B�/Q�d}/�;�[&M��_���R�I��t����ά���&�_#�f�9N@�۷���k��e�h/kz���-���a�3
���D�Qa#�M���T�ӱR�T��@[�QH�=���^�z���n�~�au>�QU��N�A�Vn�,?��V�hc�z��#w�NI}����G�0�������?6/�~����l�{�W@�U)[Vȋsn���rl��լ.v-+- ����+7G.�<��C{wK]����q4�2�b���Bj�0�Na���(��yϯ4���tY�6����c7�����r��m��+r9�uڲ�"��b��.�c�Ɋ�0�j�N��6^Z4dw��k��Z�5��iU��8vJ�1D�O!��1�J���s�T�{�y�"���D)�X�"�S�3��`=���G���p�Z�0��[����Q��rb���34�d��x��f��b��yɌ*�qJ�&X�e�kr�n�:=��z�񻾾AE�=��;9V���L�\i�����i���^pr��t�1���|�64��ה�#U賤µ+�G5ᇥ�_
�雦m	`�*�4<vK��I=��N{w
q��p�-�R�V�G3���8m������#a�8��v�-zy0�7&��*&�}>n�.�i4�޵ٍ%r��ǝ1� l�g������v'���V���^y���ǹN�j�QmɅu�X�ku}�����Sx�0��uԺm*�2T}����P�ƭ����t:w� m�kb7� Mt��zv�<ʾSE\��5[K�Y�_��Lc<�v��^9˗ew�y	��#�l�u�E)7�c�U�w�\�eCEE�rU�R�p���~ԍ��v�K�P��P1EP�����f�Y�p��_>��q�hs�ڰsM�9�⢭]`�tF8pٺ}$������1�]T�O�'C}0|;�wU�d=�qŕf�[��&=���&wIz�	m�W)��7t{4���K,�!�=�%�%���O�O��:)��	���K�� <��й(W,�&sސ�]�s�ww�^ً�~s4OR���L����Iv.ۂր����E!{��9�S6�\B�GTKhΩ�$�;��WB�_u�5�'u)T��}����{�'���q�$�ɘw#ٓ��M�U�����I�PDTa�¥LLA1�-(�V�-�KU�B��[�TGĸU�ڳIr�"ʕ��l�e��ЩZ�Z�V
�qF	������jۧkfM:�-F��"��H.d�+*)m��Z˕B�T��Q�D�[s* ����؊E-,�J4���LW��JP����ZQ�V�"���l�!Y(�#Z4k�"����5�F�Z��ʖ�*���5Ur�E#J��Ю8�mZ-Deb"�-R�UX��ʖ�+keF��+Q�E�f�嬶�j-E�EZ�)�)��mĊ�2ն��G)Eq��ؔe���k-JV�DU+\q�)lbV��+��h��4ŵ�[0m�T��f#�f�ШZ[l�T�i�rܹ��ť�4�TaPQ+E��Z�Q���P��-�,��k���*�**���e-���*�L�jc��ZF��-�Z*�#Z�QK���U���#�(�(�,���z����aU�k�AGd���πy�A��G�)`᪮�l���2}�u�I�Z�r@��V�	j�m�L59�Z-$���qo�=�&5y�Զа��Hp#+e���(#�<Qn�cX�P�I��b7sxo�WN�=���O\-��FF�ZϮ�U����c�c������*R;��PpɲӰ�_,�\�Dk��u��A�X)����* 9����s^��wu�qY{�(77���z��S�j)��(œ��|�|�`��_��ݘ��)Г��1�C�<%<�ۓt;=�
�s��h���}}6�2�][���D:Ս�H��*u��j�-���H#'L�t��Os���txE���K8�<�-��`�9行�4��f����yO�X~����J�.�����_��ʭ�Ys��n�;r��ݿCRMe\7ֵh�a��iJ���Cb�H��&R3S�c������JZ��Td��bVSw]I%��$8jm�yU-8ؚ�3}.���P��G췇����;�x��]��d|���9��w��I�R�My;�ے��rF��.,k��@U��D޸��]�i��ڕ䑺�����xV>�;���K�L��u���}�0'v����6�ʖh���e��C싫�e�4��VAj̄j'�t��z��+�#�z��M�b�"�$�\���@�~������.y'�2�@�J��<3՗Ȼ���gh�q��I��⠧0�o�9�Y+�f�E���c7p-Y5z�'-W���s�yD��� 3ş/�.�*x�e�ݚD_�c��`Mb� ��:Ov/��M�lǓ�y"vϫ�%��K:�V�͍W���)}�<6���	�<�
�Ɋ�%2�Qv��djɌ�۞ի���5�2F)����.�AO��3�Y���v�ѶۗJ�W�^��q�)ê�:!2��R�cwZ7O��l�j��EVډC�nA_=�k��K%��ռ��\�GnP��JwlgK��"A�쇖Ƕ�X��M�L�p�}�m���&��(t<��U=`*{< �$$b��@o�V���7�2�:�uPꐌoj�Fٕ{mk^]d�-Lu��K��Ĵ�	��S{�����g���}�S�UO<�33�U�|6���z�ѓjȆ�i0m'� xMj3��n/?
�r#��� ����mܠ6w+o��+2�0[,:5�y�1,�{T��(>���qMLG���0�:c����cS�"��k���ܼ��پ�z��>Y�4��jn�Y��^����w��)4�C������>�d':��*���O�"�Q�����]}��}2Y�������V�3kd��>1v#�N��ƥ�O6I��¯�S[��ob����a�ao��6>�{�2÷.ͯ[�.�]��ǂ��R@ �:��(tW�����������7rwV*jð���B�g�Wb����p�L}$�|�&���!����>�$nU�m�qs�c}SC�ui��n��X�U&M�sIU �@��!���x���9�R�'�%Ý0zώ�764K�>ǛP.�# Srp��"�o#۝/mCH�V�v2L���-yp�����Pee�Y�h�,�Bv{e���X�Y���"p �#)����죆�E�On�<*��u�v��x�uG�D݃p�U�f�N����0E�ڕ�TDO���P���
�f�A(f<��f�U�u�/�^��z(��h{ä����L��X�i�t�K&�����,؜�!��C5]��JG/�y戹Sa�T�ԇ��Ρ��Ջ2�~̤�2��<t�q�,���ph�1����C"˩~�x%�BE�Oj@�-�g ?eOq<�� �aQ��g���\:;+�ߞXJ�p���o;Ӧ�ϟ���E��~|5.|G��xB.>�z�VV�z}�(�ob��
:י���#���\������k�S{�e��,��c��\���~��ܽ�?~����ޭ���Nˌ�k�*���Ióivğ+��Ao�ۜ�[�!E��8j"M�E��*�+�2E��-����<ÕN���o�W@��Y9�֍=J���#ƴ�t�
�{*�����ήJ��5�l�a�)�i��|9�|�Ѓ�<����=�h��aЙ�	,��	�T��W[K��t��#����V"����G�L&��(�C^S�W�Z<},�=җ"|���]<���=�*����b�����q�?2��ia[�r/�刺�Q�w�`�/��
NJ&��`��N޴� �Z\*8)8y�k}����7�ҋF�]�p�1
8ʘ��C�G���fx���<�݇�T=<���˄ixv�"k��CQ{ӊ��X�S�9;�Z��6�k��v����9��W���&������:W��B��j��=���wfi�iѫ�����.l���DBmK�!��M���~WK���w�^�;��/Lܭq�5�)I�73�9ݩdIp��h\E@��ĭ&�#Y�!�\F��K^Y��6t/�йN7�wvmhUz���y8�����Z�d�^����������Y�D��o����%ni깕�������C!�;V���!��\$��5{{>�P��̔� �E���Q$�a9ն�O^��s����z�'BW�hیpэ��R��Vk��9��m���0�����>�d�IՕy�?o@�p!��#��uи"��(�V�t�v�'��jr�=����sj���ڀ�ޭ"ۂ��g%�kܚ^j�`>κ%��k v]�noK��&��E�IGle��Q���/n�;���m�����Z൏qn]f9�s���=�Zs}[Jɑv�U�܊��Vxҙ*#n�w�N�n�.n�6b�����w�v��B9����T-�L������)m�y�C�
�p�q��ٛ�R�	e$/#r�U�PD��(d)u/R�����y�1e	Cn&v��4+�A�}X>k;�[Ԝ��Vqd���1XT"��pS�G5��:�� �D:�L_�����3�Y[C�e��O��l��vp��O.�[�i
�K��j��F+9���/��P�/�є��ۦ�gR;�
N��%����Ǳ�iѝvy ���mh�hu�|�&��r���£}�W�<�3T���&�b�s�O}�t�ϼa2�\
�bPvQ/nxF
<�a�Zǜ�84qt0=���Ve����D'�d:���b�G���X,gGU�s�y�u���u~��_b}�+��7d�&��~T���X��z&l�Uz�~�D�ɶp_�ʾBnU�YB�g���ڂX���E�"��]�P�j�L��WW#����<�o��)ʵ�q_m��3�E9���N�t�"�4Һ]��+�Ϳᕲ�9N{>rJ��}(-��*ɦ��Or��O�˳� 6kH�t�ܻ� ��*�#��}����N.�B���n��ri�GVN�H�.�(r~
�i���ز�Q.���P���F�F���o����K� �p�.�!ʶ���SN3]ēȱ�ݨnJ:2KGM�2�YU�Uq��9q�����G��k��=B	gQ��bv�g��yԓ����N�@�Nq'�ƷS�<Q�F�[+�_-.d�P�&�D�˟^dVK��n�".6c�w;qK$�VǬx�6�gg�7WX�����f���zd�w[���/N�*����t+l�l�Q{u�C��'3�º����V�bR�L�Jȸ{��#��놳�x�	���Rƫ�e�"���{u�P+^��ɽY-��'����S��+
��LF�Ѻs����5cs�;G�w���Q�R��M���K�og����0�U�Y�J��N��K��A�쇖Ƕ�U��~��4u:�J��~�l#�x�8-�Ϫ���*w�h��֭�*����89)I]���Ůa���G�oq/ޙ#�w�*Rb��F���I�t$����:b�<�'�_,�X�9ySF[�)������4Kǩr[�[�}6��w������xd��t�a! {�h7����`l�Z�P�����&��P\�23ʐ8��bO�:��J��.]�ʩĊZ&�R�O�&�X|���M�B�a`�Ҟco�LV�K�Z*��W�d�
�{K��<Ԫ(\K��Ժb3Q��3�)M[T�h�!�>K4Y��p��E�3?q{� ���e��xh<|*�3���Bǉ���8<�	�̱����y����{
�D@A�(��G�\ko6�m�^+��������V'���zGg�P�X�g[����K�I�#�ˮր�B�	������y��@C.��6&��jwez��xEv<z%K�D�#X*`�P�sg���3���=���`�d�}<���E�/tX�Z��b�cD��=�˾$�G����L��LH�������O6���e�<��IB�AXj'ˆnSpRe�*Ǒ��4��`%�y���r�1ƫ��"h���� T7$e{��t�ѳSk�nJ/Լ)a�q�|k����u�
�hT����v)�k�nt�8���xݢa�ʬ�i�6V�ʋ�S�ܵ�F��0����Z|�������q��aj^�,��eu۬`�g��jq��m��8�S�{WSt��3�[aeB��Y�A1ogu�Z\q��{�`'A�9����Q���TDO���P��P����%ǓV�H)��Z9����+�o^��v���]F3~	��X�"n�!��4h�e�C�U�f�s�R�9�$s}<�8�O%ڸ�3n�8��������.J���[[�y�.,>+e�����M�]�mg���(���(:���Ҭ�M[���	,z��ua�)��Cüc*׺@�f$�~�s�*y�j����!�5&��ە��H�R�8�E�BS��y�v:.�vm&��Į�]�r���ԏ�0]!��uҡ�����oݦ����)�T�Sx�o-� Sn�B�/�pVl���=�ZF	�`�I��!�r�4>�7�.�f\Ѱ��9�v���i��Uk�G�&_��p7ۄA>}� �"`���O{E���9�|k�#�+��iw.���wFL�F^�f��
c]I��$��̮�Z&oe����M(W�r@�<�C��6z�'P���N��)�sM2�Ď�9vgw�	̐wUj��x����[3��@���y�ٛ�C�!�ύ�x�o_Tֱ-.���N�H�LM���~�_���{�8�(kW�����-����9�k.Y��"�[�a���o-SM�=�e鸄"�M��\>��\��bv���lx�;&�Ia>ւ�����s�WSԹm��r"�yp����U���渜l>�Y�3T�998[.��j�ѨO�_v���+��B��ԺH_�ƚW�u1�t߇:�z`��CZuy�x���l��t>Ǔ&�0渁~lJ�.P�lT�"�M	��~V)s[u\a���a�3��[���Z]c��͵q&���4/��P*������sb�	B[��WK���?:�k��̖�	�M�W1���e�O��;_I�ʼ���XC��#Ey�uи"�	��gtx�4�`�)��gNE\�W�L<�����դXn��3���������+ӗ��R�}�bE[�\��Ux��E��J{4�á�2��p�P����0.�(���9Eιٶֵ�v�0�<���pe���z0���(F�Sf����q��7�H2`R�#6�%��ʞ,�[n�j&ˍ։ꅿ	��ӓ���[hc�DL(:��Sq�L�0�2�KZ��Z��1J�B��<pz;�NeC��ڑ���V}*��!��T����^w�c���+���1���`c/�`Lq�V��)k:�N�	)u��1͹��ʈ���܋0Wعt���G����r�O7�σ�>>����Uv�l�ֺvX�f�]�ʒ�K��Cz�C,P%�A>��������lv��;6�O�Q�	[���d� �_.
u�渟g\k�A�X)��Rx�kn��=�WN�k�;�gN田s%&v�#��2��l���x��p#��9�+׎Oy��f*T�@�H��/���v{*��,'��ka����,���]�v�d\m*6�QƯκ��9�·Z�9D��@����S�R�έB|�p��sD�{f��r�MM�[]�����],8`�3�g_b�"�D��A�#�[�P�.�TK���:x��i���m�#y��ܓ�+e��P����f���tƗT�PRe#5;�v9����5�L��V�'�)��4n��J;�bF�j�f;�Zq�46auTJp��0������������:��bL�V&-{Q-]VǶ`����������-$�tC���]FW,�������I�㞈
�Ps9��w{x&V�g��{�������Y��^b��a�ݸ7�hsӊ��5�2틩��\��.�_^Zb�z�[��/U`�����_R5,�]��C8������px�'eY.���KP�Ty��Y�VE��M���_M�>N.珣,e��S���ܶ�C$��z�@�lc3Ut�|�Le]@@ѕ}F����V>�mI7��޽lI���=�l��c��eh�l�b�5�h�3�K�p�S|=c���}�Q�#0��37r�j�ap��E�&K9f�'Q �;.����\sY6�!s�E:F� ����<��Vj��KUG��	�Y+�W<^OLx�,�cs�Z��YԮ��SJ@J�e�ǌ��9��KqM��j_gF�N�7'T|�{�k�GM3m���JN����7v,Jb$����k��%Ej'w{�
9X��&Zըš%T�).�;3��P;q��yF-x���`\Mͪիb̹d}��(S0HvWkt/�(K���L�,JNN|�t�S�����Ϝ�u��o��pk����+�	N���,ߢd�}|�x3���Y�̱C�=ԕު*[�eډ����Y�a�L+v�D�/ �e�V�Z��A:J��3pL}}�q�ձ�ҫc���OX��H���	��^�<A���A���`�ࢪm_N�J��}j��8�uǮuc����a�����r�>0�v��"�c���Ӈ��L	���6�Z�
���9��9�uu�v��|�n���۩V͊�kE�2�|��(J���;����8��2�{˕큓����Cy����A�\�%.e�;�%�.ʁ��ը���r�
�����]{hź�E��Gb�M��۾��H�G�X��LgM<@'��=�U��Q�3�U#�u�	M�1��2�����b[J�Rޫ�s�?����M�,�,0�zc��͙�E]�خ���ʌ�v��7+O�)O)-��4���}�)Yگ��&�h�S�D��ʠR��l���N#$���jP/p���%�`�]'	(��1�ɦ�j�M�KMKX>T����77h�פ�`�|2�)e�p:�^yQxC����}�@Y�����+G��85'�9Q�M��o�^��������jgot/�ˏ&e:]pN`V��tBF�u�^z��J�y���g�z*_[���:�}"2=��Z�`յ�.���z�I���v�̫�q��B�uafǫ��� ��2�1��(��7��Q�&M[�n}b����h���[����Ʃ�37
�oj�k��@)����p>����heڱ�T:rT��q��	vo�[����]ܞ��nln��IY�5cR,)�hQwe=�l
�y9v@�7m��t�騘*[5Kee���l��~sZ{J��M���9N%�j�$"T�^����?��ֻ��Gx��TX�GR}�wO"ni'8äG����YW6)�_WU�j.bU��=���/!�U.eJ�\w�3fl��ə�+ɒL�B�R@
$
�J4��q�EJ��R���c�d�m���`�@�TD���j	��T`�[e�V(�-�V2"ԭ(պeLJ��\j*�GE�����)s2��-*8�2�҂֨�h��DZTl+�曅t�2�R���i�d�k�ELVV�J�E��TY��E�(֭*Ⱥ�Z�Uj�QE�h��f!�&T-m����a�i�1L)m���V�Vŷ�b�N,S)�VTD��T�m��PEeBօ[[T[j�
բQE+\�P̱\)�3"�U�F���j[(����)Z�����H��ҭ-����X�6-�R�qӆ���։Kj��b��(��Q�mcL2��c1+Z�TF�&[�Q��`��*����U�ґ��n���V�����іʢ����E�-1++*��˘�uk�)�3M¨T���c���set���<Uׄ<Y���@w,������VV���|��f�+lp�x �f8�ct,��s�|/���ܬ��)�B���{q�U{�!�r��}k���:k�ؔ�mY�g�N������oZ�Dv��F�Y&����^N�x2��G�Y�,j�������#�Z銯�)�m�3OEeօ}T���
:b1T��-��A�W��j��X{�ǯ��9�*}'4�W��A8P���b\GD�d-JXT2��X��uX�\��[��كJ�<�d14p�<�#�:�0����B@߱K�L>E�Ӛ�P�=���lAa�����}:!��h�Na�N�A���B��!`0��9z->Ȫ6;cuS�t��ݿ9��:=u��lvJ�T�p��3����B�.P�Z��w�j��!���9�u�F��g5#���5cg���4�	xˡC]����o��+=�!-�:,}��cP��y����]��y㧆��n���va�ǂ��H�gt5�i���5�6'��T�#L�x���[Չˇ{T�"�P�N.��c;!Õ0\0�_c�F�g�p�]&�a�2֛Vz����{7�Y�y�w	�A��y"��-Q�rX\�N�%�3�*�tf���m�s��C�����m^.�q\r}vM���(m�����1yv�ǐF�ul� jn��ioF��Gu����#-���'}\�j\�vN���?�ةg��WXYU����w���aߺU�$�5p��y�=x�g/f7���l��-%IH�eO��CD���gf���g�.���궤�rad�If�|�^���}�wu��c$�J����IAI�v���̼��!]Yk�{앏l'z�}0(+��D���nu#��O^iZ��MEᛍ�Rf�1��X�n ����Ԍ� ���)�h�5���^Z����IjH����/�eE{H��8;od2m��]ojk!E� �_"�?nUG��!E�ţ�	�щ�'��R��4h�>�*���wO|�Ë�t��E=IF�r�E�S��D(쪄5:��)�M<t�qW����� T֎ת^t�.e0j]vUx�,+J���[���e��Us�jw��^�	��^��W�m�ί#��{���&{4�b�J�K�Z���]-��-�7���w�k<�s�r����r�h;P���[1���^����y��(A
b$�c�U(���4�Rp�l�����B>~�+���w��3���Buv�������@�>��3���R���>�D;Ɔ.5ι�ݚ��w|��e��Ԗѡ�o����%l��Q�eoU'ң����]�S�&��%$z���W*ݞ��/EԻ�˱V���o��n�)��3��("�_Н ���haԂ�q+]x9�;Č6f�6�#���݋����f@,���{�oT�LS�U��@�X{��b�I���n
�吆���M��^�a����c}����(�9t��mjM��ŵ�}�j/�zL��C�l/3���:6�&�ј�rGK�,�[𠸊١��객����^��1
5,�M�UK�+Z�^���It�{-Pu<����yp���:�TgI��a���v��<@��{w����y9��9�-0p_T"Աt�mO`\KQp���X�@��r�9ں֧A<1�SWy6�$�ڑN
�ð���lJ��3b]P��&6Quf3���XBK}o��¯��d|��<~P^<��tVD����jτ�GlJ�f�q	:/�s�qd��^h�1kc��V-H`���}Zu���6�e:N�;P-�i�j����B��g���nٕu1f7��Q!��:8��{kה*�.ﶶ�7�Hn
�-��I^��.��?h�6���:�wmsɶ�˱د���>�	��*���u�`s.�5¶tԵ/�ܔt�K��:��	�n8m����M�L�7^ʳϢ��u�^%�e���&9����D�����#[5	������^�ץ�2��4cγ7a�j��α;��v��S2E�Uzd���!ш��(�wSâ�i�á�/Ѷ�z�ѱZ�1���� _e�E7݉�(@���%6��^>��P���R�1\�s�{4:�6[50�[��w2i����u�)NUi�-1o]>�ד��diɍ^j𥶅��	�j��m-��_�f�Օ��+KS��]u� �X�m�-=�yLwc��!�P�rK�����r�u��	��,���,��r�&��<��_r��>�M� �D:�La�m�+�*�R�5�����7I'G"��*��ȇ�g#˳��89B�l��-��{��7�<�2-�]�n �!x!��E���f:�Q�I��>sO{"Vfb��M0���Y�9�-i����e(d�@�ih%�3�W��߲�+Ǖ,=���-C]�����I��]��rT��e�1���}�"�D��`�)��P���
fb�C{�aM�(U��������}i�w���K�� 6oV\�w*f���$�G�`��a4�D�������݋r��י��&��Ʋ����0�2�9��p����k��9+/���MP�U3y��5��]�o?u�-�댗���.xHP��(�1�r6���8F˅Q��H&Z�[��"G|��9H0RrN�l�Xef��4��h\�t�����긃�뷫��� P÷�L�ub�����|e��?(�\���sTF�/�&z���=�$�B4Iw�ȓZ$�|m������T�!��2�ei�6r�+�9(L6�\EOQw����,����V7������e��(Ȗ�[�u}�%�+��:j˺�N�����U������iLsL��SV��e���d�vMI-�E��Z5:)���\,����4�}q�Q�rZ;��Jv�3e�]L��j���q��-��P��!�Lf�sî!�K��{k�.���S/�Ոڴo*J�Kh��g"�8ɕ�"���eօ~��vt`L�O1��u�t���kLоg2k9��kV����ᴺ�
<N%Ũ�V�p61���.�|uu?(\aw��2m<��<���}E֛��>f�J���Zo�RfX�dзP�a䐐7�X��øE�Ҝ�ͭ������MsS�:��h��`#^'	�6�c��W[��z&�R��D�fx�Oi�S����f��I��Y��z�s�^����EM��n���t-���� 9�=��=��p��=:��y7:e�u��uʂ��t|�]�N��[��R�
�f�����:�f�����n�L]v���-F�y͙�%Zb>Μ�}�%ח���_9��EDC����\���JL���e��]��F=�e-MD�P�m���	�,�-+^Qz���#�O�����ɇ���>ff��tW{��L�AGl�<配V�W��aۗf׭�p^��ϩy'Y qL�wڏ)5y+��&��w���:cPs�14_9Vv�֭��)��S��_(ņs��*�A�M(*���dC�Cbh�ɬ1����w��	�����q��ƿ��i�UB��N�W�˺$�$�b�)�q�
ϋ�՝��J+5=�馜� ;�d�Y�u�5�B�(N$E�mN���Ia@VK:3�2�LQ���!�'�zV\�Wm�w���6bii5 �mD�0���椌��&��ʸ�__�w~`ǆVQ�z����o{ln("�O>[�Jn�:;gemx�̟u�^X��J�,����缛���!�{v�We��W���۱��TTT_Tc6���O=�C���&
��={�&��7Gm0��״�R�ë#�p�nƉ�M����n��[�d{oZ�͖7����p��ڢm�ch;����y�Y�#O��z��=��ebN����%}rwDZ�����n�2�A�wc�r�9���/nݗ%�Q~�2+��8ߏ���~�q�D(�ʨCS��؂�Dמ:c���3s �}h�'���}�����C�-z���mE��U���E��G���W;6�Z�=���X�mRsZ�z��=�����_�g�Nčҋ�J��q]-���[$?V�d̇��V�@Onwn��Q�V��a��W�Q��<`�	t���R��$7����b�m�b��HѢ_�	A\b�BuE� ��+�Ӟ�ܦ$a������fa�^��K7���(F��0��D׆qa���j���7�s�ġ��C	���������rU��n��Mp�>Aai
V�ͪmM[�mCc#�Q}K�`�S�Kr^�&ty��Om#��yhԔkı�ߦ
\,1�&�zc�d����<S;|��v[&��̔�X�)��D��O.`T'$"K<�e���P�Լl�5г��{�x@���i\�3d���кgs�u�����bÙh���(�y�~��fC�xi�.�(�#��T&������e�Y�Xmb1�B�ӫA=�ɺ���f�k{���9�j���b��u^c�,��N�b�[�������Qv�uf�Ԥ�4�����}���Js��m2.�d-�w�>U��0#$9��˓;�{���;-5RtX]�i�ĭG%v��vD8:������OT����)���42��$}���R��x~J�;+�Ȕ�
~Q�}��0r6aΔ:��n���u5���~�
�dp�yj�BǶX&��*�L�r/:��Yܫ�u!�u�5��m=.dԆ(Sq8��I��y��V��
�q0�:�E
�6�7fl-��U<�ֱ�D�s,g���i�#�j�r�<��
�^�3q�Cd\m�(�s/2��=��(�"1�'I������}:.���x~J�eS~��W������@�4Z�i��ގ�3{��cg�,0��}ӯ&7S���|j����*���;���7�Kv)�s���D�;���n�A�ڄJ���Qa���]���������E�Q��6f"ճ��N�F�R*���*C������9��Ⱦ,YN��՚�bS��{�i�}yC7�*F�ϗ�5i2�`��f]Q�W2�4!�,��+Ώ(�(_/ ;.W����F]ks�ul�0,� 9g#z�$���&�#fhλ=%�P��GZEt����Gt2hwEp�W[+E��1%*D�3��<��+���vE�0�f�%{ ��=mS�`���=��	�l��
��	)ʌ\e���a>K�4�]R�.���a����3�Pu�UA\L�Y��S��|�t�Vn��mJ<ZT�h�ؗ�u�V�؇Z��H���z�Z�陂�p�Pyծ`�]�(h���7&y����9���#�.)�|+"-ҳp͊��B��GI_#�v�.i�����ׯ���#�Ɩθ������-���ў��t卿K����O���U���{&9�����m{�b�8{y׫ڦ���U�rCb�mD��a�Z��S�U��'$�"�EĔ5Tߨ��]e�_�Qsw��$��)b�@Ȗ��K-ͮ.f;����h�uH59R"F6�\T�u{x/2���I�K
�3P�o7{����B���Fm��M��d�{�4IS���x�g�V�~=U]�j9s��X��w��V�`'��/�o��׮��bb�����E����Y��4w梆U���#�ݖ��Q�6��1�kTC̘�)���Z�vޚ�~R1M��Y�T)%�=m[$0�g\�����klg�q"�C��Ǣ�v�Z�����������������5�9RvX�|[��)wl���`�V��QM+�7��5QX�2�s�ѭ��Cؚ�Q̗�fH+���Qs���T����e�B��U<�\"��!S*xE�⽗Z;�](T<t�f+��<��8�]j�È�Z��XːM�d�=����c �B���I���g2�Ǉ���f_���D�*yDt|����DYۤ�?G��_�
�& ��d��7�R�x7��)ݙ�JpLZ�yҷ��a|�P�9��`"�r�Lu��yyTgБ&�S��@ʞ�����=�i7$��d	�j9���B� (i;�]"�u�י���P[U�p��wa�{LFb�!ս�.��!��k�#����!	��}�}��g���Z�lA�9��i�ū����fXǎ�ȷH]�f�x(2��۩��u���S�� "���V����Zl�58!3E�gk=jر�h�3�M��ּǁd��(�nRiX��:_qۆ��Z�W��+�ޘ&x�X˰TNL����ݾ��jL:Ȫa<�A��d��y��|�RiA���i�w��g�}O)�-�����,z�O�CW��u�S�/g^\��қ����R��o-GG
�Ήwy��C���c�[b[�3v)J^��Ef���Y��>R �[�ko/sf����nv*+����R��ʰP:w%�/�%�4����ͱ��dN[�H�P�e	˾@��세�G�fͭ����t1��;���-�5:�� 9�F�i>ue��{n �:ђ��{����^q��k"��k9�z�����M���ҏ:&�rP�V�H#uu�w������^G�<Ln�_%�x}� N�nдw��4;�Ֆ�-��!��3X��T�.G�~Y2�;=̢W��Ti�YxP�Tк��x��{��U`�(�3U��tG�]�-��KE�
��P�U� �l����?_>���,Wi��m���5��&��}�����V`=���.{�v��T��u�O��bɟ#��xs9d�t�@a<H���zs�q����j�ϖ;Kgx�����_Lܴ+������o����"Xv\�,}3�zQ�ɷ�zp�H�) Ev6��o�m����P��"�a�F&�/����J��Cj�']Y �������'t��Zн��d���We)��b�@an}y�cd]�IZ��a�o$��qWK�Y�,�1eԤ2�g�5�����{�S��b���x��op���"��B���J�9�wh�����q5��X��oز�e��xn����U���|4E/�I�Z<8f�5�psۭ���͵P�5��|�j9<����w�r��1"�pQO��7�i��#;��x=�!��%D�0���!1��{-9�mP��ҳ�+���w�G��嚤����Oz9�y��Ҽ�ڠºV���=qf�}�k��Qb��k��n5��w�\~b���>��W�$��"��v_^�<�:q�<J�7{�FAPv{gU�߃���ٸ��U�w�J����g.�R�?s�TX́b��@u3;�:��� =P�Ź1ݢ�º�|�����8gb�ePQ�+C�]�ZK�#!�B��Cm������n5�w�V���y��1z��X󹙐܅�b�ԍV����z;39�W&������+�wFa�6_g��1ѽ!����nk޲%p�J���p�dI����۾z�<s��9G�eC�h؏V���k�-*��Ͻhq�ɭ�j�\�).SM c����������OtK#��4uSU���.�sK}v�oP�Q)�+p������g#a�R�M��ȝ��X1�u̇�zXj�}d@%����a`���.O�{�K����+���\px�|y����6l'�6Z�o�����nZBqiq�I0]�o�}G���P��0�z�{���k��/ٴ@O�R\&j�m��\a��/>�U{��l�Ƴ�v!���cu��6��7-N^C�+������U�;O��c��}A%wIPU�@���WF��0V���ql��YU*�Un1��a�r���C�T��`Ҋ
V�ԬAAUAmj��2Īڥm)jXQmJ�q��5X���*Tm%EE����f[
�-T�9�r6�c�+EjĲ�r�3XWCV�[���.1֑Tb���V���*f���\n�TMQ��EDƵb��ֈň�9K���i��,eV�ش��i���E1֮����Y�DF�]Y�#�fe̊��\(ʙn(ղ���8Ֆ�
�4fcAˉ��J�[��[5j����Xe.��cZj䩀�R���s-ʦf+��)R�Q��Z��cA����i�ĭ��e�ŕ��d�U*R���b�ҕq��娈5˖.TUm3&0`��V�
�h�ZѴF�m���!m��Kt�JTDV,�6Q*҉YF*�-����#imm��m���kX��b�7(%(��V��T̵AV�FҬF*��X��YD�V�-��TU�����"妳QJ[Q��b6������ߞ�z{�kP{N�	�:]�����g��ޓ**�`т�� �.�P�AU���Sz#Y����867s\)�#ǛG#W*l�6p��˶	)�l	+���3��ZJ�fKˆ�PReݨ���8��8����Ģ�	��i�S+�q&��H�Ğ�R�;��(s}��)�r�)�o[1�|D�)�n��:���.�����I������q���A�*��l��޼��7E��	A�dM[1W�P�l_Tc6������5�"���0�{�����o'���]�B_��v�g��/ԽCp�O�l��n�	���ۼ�Y��R��ږa���\<��p͌cKʯł�iV2X�u">Za%��ܒ�Ә��1*X�L�8o��;�y�_�g�N$n���ұ0|-Ԉsٗ3�x�]z�糂9Z��p�Tx��Z�oNx0���(Ş+�Sf1�K���Ί�}BoNmk�Et
T�k�K� ���ũ}hg�\Ok�=C�)�K)��ky���S���
��m-�T#@a�UG\��c8��L7�N�z!�)�+���#��D��ep��8�/ݗ�C���������6ۖ/M�/{�%{s^խv��/u���~�M4�}Z~�N��²`ө��`H�ƥST,eF��^���3kFwL�Ph�����/5��ۣG%F#�G��ׂ�r�	�8���9*5(�ަ�-�Gz2җ6���>;n��gq�H�m&����h ̰�!JV���M��Kje��]\�_LW�a��o:L*.9��LNJ5�����-�8��L'A�kx͔߶���-C.���]i(ޙ�/��ى��n�Zys��5.x+�c��s *:Nl�W�9�ǵ�Y{m%�ͫ��*�u��-0r�B-K,9�I�4�\��?�3�*��z��Gv�rNX��S{�!w��¿4�[bV�na���T!��6EE{`�Ek�6�r�LdTj�)h�q�qT�{\/�}V�$�u��ᖸ��j�'R;bV0���F8fn�(��GG�V!���L�̙轫m�,��
��g�E��T��݃r���ྩ鷈ќ�tEE��6r��9W1>�t����.��6;�P�	i"����8ԗ�i���~Jt�%|<��3�GJ��f���և�np�^�3xt6Dd{ݏz�re��9/��y�ߍ�:��ۜP�+�O�6��87rvK}2P�3T����,U� 9�	�f�;�X���o{ea�P�cL����ē���g�j�5��dw_�q�4��>:6f�xw׬���aB�=��>m����Y��W_XG����D`��V���y7_T�v��*'�onjw���W����78�_�զ�x%�����F����������t�<�ݸO24:�5������W�.�G�=�����qy�X���\y`�e�\0�u,a��x�Cuü�#����KjN�Ȥ�QsGt����v}J�!@�1*ܤ�Y���-t�8���C>3*�L,y'r�KK�3����LJ:J���qS"8���q�	����7=�yS���z�=��u��L��T�j�F\5vx�HU��h��q�/䫬�觱<�:Ό����s�g�q��Y.W)�,GI{(�C%��4�	�3
�,�3ܙیB7h�s�,�i������3��<��m�
�[�f����Q��@× p�7pNo��K�x �f���qu������h��o:�vw��G�i��,m�]�Xv@�0�1�[�����ʨ�.*|)quT7W�����'Mo:��,�B��-#!����,�^�n׷/[�s%D���VY�A[e��ˬ������c�0RV�\�|Dz=w��yd��!e�2�)��Є�w�_�ڜk,R��ۼ�潬����+x\t��׆��V�u��9����]:��]��\���bP=b�k�m���Eh������Y���xe�=��3�/s�a���rwY�Fѵ5,�+c|�:�v�Ht�o>{Mj�KGM�f]C���Fc�E�����.��_��,\o:�u�ҦDw���B�4�wN����p�Z&��7�t/�$�w��*}WsA	��vx"�ڄ��c��9I�j��`O�6��!CwKAƧE>���YG
i����e��O���J_�Fjˁ[g����մ���S�ݤy���nxu��Y��ޚ�f�a�u{�����x����������#"��/]۳� &P�x�̅u�t�r�yZI���C�#��ٸ=��sF�Jg��No�b��}(2P��G�;�3����TegvLS5�8�;���âŸwH{-Ջ���V�*��Y�&e��ɫu	6����˙]Z+2�p���k�G�V�$:{���ȆX�S0�����ؓ<��B���y�k�Py�6Fm�(�v�J&X�$~�>���Wk�9�+�lW��@t.�h�ٶ%nLT��l�+2�b�ݾʷ����<tn)B-��e��q�9}{N�5�)�fb�!��)z�!�e��kɼ�Sn�7��u���4]�����$�<=ɝ��֐�;�):�Ax�~ЂL����s�C	n�J�gl�R̻*�	�=�#��Z1.N��f�#D@�����Eb.4����֭��f5��.�d��X�����髈c}��pF�f�����r������C|�,d<t��9B��0�gL�v�&\��8�9�d��I�N�!B�4mO->�w�)zk+�u�vz�K���@Y�n�py������r^�|/�l�U]�_�A\��B1lTPӓ�c��9+�ь�"�^�7xμ�c�ŗʏ��MY�L/[$��#���K>J`�|q0�8ZG7q�ɽ��ӦKg�ªP/���*�����Ib���.xm��L�r�VGm:�}��o&�L>.��UH5ܮ&��D�@jH��yW�&���o_V~`����*l�lRmS���0o���PBo����n����LL��z�	��/f�@r�q�1���Ț�b�{U^��:c�ptW�:D��CKy]�Փ�̉٥/_�=`Bq���HO}�f����g�o[�����S�+g��b�G:���N�ީ|�Փ����g�yL�����kK^�KGY������O�_شx ���~P	|��֟�J��Ȩ����[V�Wcb]˫A���5��j����]<b�MG]���n��(�7�<yF.t����Ҹ4��VW%י��d�i�����E��Xi�ڰ�%n%%fZ������u�I8����f���Yl��i�qra����Wڀ��/j�r9;|phL�����r�x4V�XZ6ϭG��R�v7���zk�{��?4L�k�[*�Tx'�*kf25�|�(1��W�Q���c�*��L{�*�w�	��W�ރ��䯴K�;�u�/�����9�{L<3d�)o��q+�/M�������	�X�v�ii�(f�fNwE��S��Q��K~s�������D<��4f����!�
�0�5����o�H�1�XV�\�����u�����B*uT*.5�/]р�(��F�
0�*���<��Ȟ��ɬC��͓q���)%{W�J��)��'��]�)J��L�
��O`ך�E�^X�]p�a�%����>/\�D������	KA���,X����5�_�*�.��d��^�j�_d�8Y0z,�ʚ�u!�VXV�:2ZE��4��dB�"�����m^�\�m�R�QX\��_�� yz�0E8���Eg��
�#�u��5��{ّqE2ʻ]�@;,���r��G�WQ;lۻ����n���܅��}J]���z~r0���η��<�i��#:�U�9��d����6���aҶ�Y�6Q�&�j�'$ю�ؼ��h�\����c�AWH-�q��c8�Y!��}��JsvF�<��^�X�4`�Ռ��W{y�u���N��t�rv�nz�nB2�3u5*�3ZX2�/�����v�бV#��8��YN���ǳV���h�^'��|-$���lM&�TLJ[ZO#h�. -:+ϳ���Ք{MV��ŏ:[�3]珠�z�m=��D0m����MT�\C�u�������n�mtM�=���-�^"���s.��
��=yȍ����e2s���:�����;P�6\n�OS-����<j�USzik�K���EѧN�Ǘ q((0B����zW�lq�+�Yc=��0\Cj���yLw��K��e��T�}��|*��EB�����5�QF���b�����N��â��M�V�+�zr��J��{/z��X)���n����K��"�))���,��(�c�7�����6�r�w�6x$o\L`��;m]�C$(�f�fPw�����1P�d��- �5��s�PPLۥ�~~����e��]c�1a�I�y36�q�4�a���6����#+X��X޵c�Fл��Q�񋡾YMy{���&�<�Rnr)�\7v�99j3�l�}|�=1Z�Y�0���QZ2�̕{��0��іy4����rwZ���7t��������#�d̈s[����r����L�\���9�b��xyL�j�8,��&x߲_bϢ�D��`��3�X�j�y^�������(�+�a���������1i�2+�x2\9��a<f�%�W�{�j�#�]T�"t��4wLiW��g��wӽ�X7����^��9`��*�����ݹ���[�L1Z�|Y��C��-qv=����TN�=�%o��L���'���5ޮ���9<z.�4PwR��NT���@U�B���\<���L�վ69����1�]$d>�{Յ�|�$�7�Pi���ܔp��Rt�CywB�d�.�:@�%VdM5��j�ۇ	��7{��V��x�6��j�J���k��$h���J�u�r��ͮXQ����|3�����]*�f���!��t+�o��ī۬㥀4T-j�{��[�p�,����,,�Ǜ���uf}NƫP�LVU(�Tte�q�N΄D�R�`�@�kj��&nO+죚��8�Yo��Ϟ5xg���ʨu+ �m��(�₺fC�]��Gk��-=�U���� �G�B�U�eY�4!������Ѻ���7��.M�S<#}�Ā�	�7�2'�j����tV7�<�zU^P�X����Vb�C(U����y{�-k��s�������,S�x�G9���9_nh���Z�wڏ����םQ�� X�/3�U����*��Ҧ�:o�1)n�e��q٭��SAW����R��u.9���к)댴��H��Y~�b��p��q�m��v$�,X����!��c�/8�m3z��s��bc�'��:{�})�f	;0���7�ki�.�^ý,C���u�d�P9.̅��rʷm�]>�Ev�A��չwذ-�9����'Ƨ�X����(�+���̾�=�V�z�;q�^˩�.�X�p�K�^_;�|:�i����'떉�h��yS��s�ۜ�ݸ.��T�� �r��o;�1��F^^���Q�&`[$j_�d�2�_�B�$��.��&k*�5{G��c��xI�ǟ��{7�14D��4�(���M��ѳ�����ۆ���+���+Rj��,<�1H�� Z��hw�6Ƒܽ�b!�ř��0Y�]���i��f\�K�m(a�\xw�n���	�幧v}��˵��;В����\g�sq<d��?�tM��9X�aE�*��Y�i��8��乆��޽�\j��m�o�٦��э{���|m��a�n,<�-���)z�_�U���N*x�2ʋ�k��ױ4%���C�e[��Տ���>�����+$+}t�+%E^5V�4ic1�9@]c,���p�B��{��v���m�qz����J��_eξ�Ř�\ɶ�4�O+���Y��P�>�v�Tլ��p[u3�Q`���`���ִ�j9���{p&)'1��\qK1������
��[�7��pH�e���c%iP�)���
y>v��~�6��J3��s�iF���d�p,w�P�:��1؛���t�N�|��D:������Mfi�Z�c�;.�,P/e�U�v�������gÇa:׼���>����;m]MK:�y�=���ϳ��u�ߺBH@�����$�����$��B���$��	!I��IO�!$ I?�B���$�	'�HIO��$��BH@�p���$�$�	'����$��B����B���$�܄��$��$�	'���$���$��b��L����m6�p� � ���fO� Ěw�o�!@%UR= h��� ����R���T��QZ(H � �PP�U)P�B���BQ+Z((l5�R
�AiY��2TJ��%e$�����P��(�Е!Um�KF���F�U[`�6�/Z���
�R��R�B�u����T���RR�m�Ҵi@H�kJ�lȤJ�!
�B�*P4��RZ�%(��1��Hv����  ��n]�E�XJ�ev\cv;]J��[T�wuֺ�wIT�*�jW2�mӧV�r��WM��ͬ���֕�����M;�m.��w]mu�j$IQv0���AK�M�  3�ZT�ʭӫ��wJ�ڗr��m]Η-���u�R�;���у�ݵ҆qn��V;�w.8�٪��sn�t*�j�[n���[��V��ܨMPxt=藳A!���U���׻�   '��B�B��w
44(P
��QB�
(P���СAB�
 ���(P�B����
(P�
 �K���(R����v]ڮ��+Kgm�]5��:U����R�dTEE"�R$���   '���։U6�[��[v�ݜ9����wC�n�]S[����Rݺ�gF���\�ܴ�U�v�[I*����������ݭw!J��8�2��Z�R�mUM�o   =��k�ú�]eK�lf��Uw9�#wv9ݺ�eM�ہ���b첍��ݩ�RV�Lն�]i���%twn��ZktU[��Ü]�W:�j��j�c"AU�TT��x   v=�c�m�v��٫��S�U��Wr�;�*�pp��m�:�ʷ;�v��ݴ��nwsv�wum;�]nu]����:��mp-�J�����ݺI6�ۈ�4�V�V�D����x  ��UUvն; m�����a�wr��nK����+�b�wv�ʦ�LÍ�\r��AZ���PwWt�%a֋7K����Z��l�J��  1�����p2v:�(�+ 
��اv�\[c���:
j�:�	UWN9Y�H�tX ]Ҋ!J$�� ����   ��*���@�wWU��!�jAD�6Սs�@7v��桠�e���9�Uصn�W 9�.��Z4*T�J����Mo   l��u�``Qv�9�gl ��\�5ج :�nj5P
6��WA� ��m:�RT�s.�N���Q� 50�*�� ��)႔�@  T�4Ґ����)� �*�� `S�&4�� �&�$̪�4 ���Y��f��9cxz�5M𢺆����HA�v�U҇�ųX���9�O��}��M�G���$���BC��IO�BH@�g�$ I)$ ����|a�1ŐQ2�!	
��]� &j�`�.�����C�wY�2��/�WF�6�����l����b������+wu�b�h+U�i�{�Ձ���tii9��n,#Q���.	X]	xF�V-���V�+N��9�	`p
�Y�;*:DY9����:��)�ӊ���-��PZ���\�`��^35<*�±�
�(�0sV`C]��줋O:���Z
�ӁoC�b�4]b���s~������� �G7.��
�"��Y{6���.�QHѬ'3^^�I/kM���]�v����V��񅐸T�~>֞T�Wgh��TȻk	(��ᕷYx�j���0���Jֱt�iGT���'��1Ԩ�Xz1�V���3)c�U����5rZ���zIzw�z#-iͬzue<=�=:	xVv]-��i��3v�5nfۙ*KTt�kK��9]ǃ�ҕy���+^�t���d�+V-�n]�v+���EP�;��x�'��G�R������\k2�P�t��[����4�l��tH;��P㍷L*�V�  �Iӗd�8ƫ�v���kP�͒^��Z�7v[tV��k�xgו�g h����{�hh�K�lW%ǳy�Ht[���j��t>�9u��Z(�wk653u-L-"�j�]]�4�	�l�7J�L6%�slP�̴[��7���9e�T�ݭff
V�i�B��J�A�q�� �M�j)BԄh��]M KR�+�.`3a���L%6�f�'[ǥIM�@�M���T�3%bkըK�:,5�u�Q5�i��cvnV: �;�{0۰1�ԗn��R.�*[�Z�w�{M2��Kk�]�S)m�^݆�����Ӂ̴��a�YA�CJ�,R����ܕa=�ȱ����i0lO[Ӱ�[���96�bEC(�d�ú �-�z�|^�s2��V���p=L�r�C�:�ac)���NY��@�
;����ޡ�5njM���uP���f�,n3Sw~�Z[���fk���Z�KGoe�@$�X�R��P�������%m�'��Q��5Գh�`�HD�jp�Ph;j��u�2P�c�[*o��)��6�S�s.��E�K&�ͪT,�"��Ό�^�tt��7P;1��J�DA��w+m� &�+BՅm$^�ZMXh�L��MU���N�-�^<m`��CLh��*;B;�k�x5c�V`OoE�wD�fEV�B[v��Y{33/$� 6$ĉE��l\�{,��o玹�!�x��t
zB��Ǎ/��ݣ�#I6:��J�8��}U�G�9xqcr��r��Se����7jV}Ֆui[�Z�DP�Y�z�&��	� �ie��J�#�]�mEl�ɠa�P��v��0�m��Y&l�0^����0�x�yyB yJ��w,]^�=Hwf��M�]�[��wJ`�i]F���m7�m]f@r�z�.#� �X���Q¼�[����Q�5���
ۥ�D���֛	f�}�B�t�*�c6T,�T�Ҫ��2�w�F) tFi�sMY�Ye�^���Qb÷&]F�u�i�WR����Ҷ�U�slѪ�3ik���R+on^P�Pf���2r�(�Wb�# �w$ǡ��$��*�Z�B3��ut�F�E�b:���n�n��%�Y[���x�wi�i`��}�Q%u*��Qμ����"�ώ4��
�u>ܬ��*_6��L�:��=X���r��w>L*�)�-0�t����'w����F��iI����v*���Q�4֩t]2�G���3��n��1]-�32�U��i��n*��;���^h$�c%��6��t�bzM�]@�,�!���)4�
PCV�������[�v�Ͳ�[�[��:�ѵ�F�yv���(9�5W+s�f�]�&��2Z�Bk�N��3��T�Nѹ�Y����m�c�kx�9l?������4+;]�><x�����m���X���t�6�a���v;�iVXY��)�F)F�"���\�f@�řz�D����<��l9`٘�����Ҳ�Z�sj���t �q<ُ6�9��ş#W��n�
j�,Xd*eVV[B��2��O.�G/S[zqj�5��̽���h����LLŪ�5�,�W�V �(n���qZ�KqkRb���7*AC$�{�
�n;�r���_jK]�<hf7�M_4w(V,�cuD���0�T�w��^Ödߎ�q�HnW+|k8e2/oS�@�ƕnꕍ"�¬����
�z�݇���`�'��fnr���n���a���$���{L��A���V���aY�6�# Gt0�pK�mC��P��m�ӆ���M�i!R�h�{���X�*�f�ZS9��^V:U�-"�K
Çn���(ܬa�	%x�V�͹tײ��n�R7xj��ѳ�h���0 ]$c�Ԁgn�2;ˊ�5'�$���4fBO�l�X7<��BH��~y���5���a;l6�̺Վ�mY�Rd̏`��J5���l�@{���v�1+�'^$�lX�ƨ��.ް�kD��C�ܖ�V��o �iG2���V�t��,�e��z(�JT��<VpP��U-��ko4w$�_�vJT�]+L�6
qd4�tBV�'/c�s*�PX�X
1�O$O��Y#tM�Wp�z��R孕��wf���86--�;�Ѳ ��U�l�z�fJY�P�����U�[_8�I��7�*Q��jaX�>J���6��,)x!�6�m�DS� ۋ`�-�ɓ@
�,Jfl�+A����Z���'0����S��wX̹�y�����˵t�H�I��	�2�'����9�[i[:����H��L�М!��i�k~�o"Ӗ�ȒK1�lnP1Yd���nfm	�)�*P[t�
�=�l0���3t�a���	Q5�os�Q��`����vZ���5�D�<��Y�vFekVjb'J�p0������E�p�+�VP����r��t�܋w�'h��cm���褰Y������ѧ34�����@Ԧ�k�?c��ˣ.ѡ��8/c��9�!OAbnհ\)�)fe�Y������o��UZ')V��k��ֶ����NU�M��Š���3��c?&�f�]"�f:L!�	��B�Y2�ǎޭsF�N��ަ��Ubܫ��R;J�����`��*W21���:�S�n��T�2�ŵljL�ދM��(�Ȫ&���FRf�Zy,QJ\pbH�ӢF�e#�1���xyZ���U�\�PA
�ޞ7ݮ���vh����Ƴ��{X;r����i.�{V2����s��o[:�����N9twX��c������VP	4�MM㛐�t���h���6��p��qћ�
�х�!S-��j�=�Q�x�R�ŹW��h�Tܢ��J���tK��*���U�����٨� �v�]̢;�
i���m���)ut�KV�mZ�Df���k�E'�ʣʻ���m����4j�����M�Zj>Y�ԟ:q��:ҙ�[v�Ls26�oc"$ܰ��`g7q&�8��^]-˄�t�d��nm<�X�N)X�o/�@b4���A]֌�`��pI򻢪i�P��AW��F�����>��7I����l�D��B��g6tR�6���H^#�h�.zA:n��CZ�� �zn�U�m�����c*#�Δ��t�UR����I����I��.*�4�wZH�A�&�4
X�1�ҫ��Um�� QA��^ma����D60�$�uL��!Uf�L�l�Z��mEtJ���>MU���;Սm7�qď[l[�$&L�N���u��t��T�1�n0Y�M�B��0/�f깖2�#t�/-+��7����QR��[Z�LS�i*����`;꽼4U��B�^���4�6�ѹjJ;w&c6��A�U��n�oh)�D&3t���&[�WKM�N�;(S�\Ue,�������q�4�êȷ{�k��`�E��r��Vk������O=�M�	ܽ�2��u�,]�˦��yV̽	�5j-�oi�l�ؓv�TL!;�j�K��p�W٢���^Kvj���#R!G�����W�*P�Cx�U���ec�J�s)�plɑ�)V7-^�v����e⪅i��aA^Z��Nţ�w��qJ�:�բn!L�)Sn�v��T�"�B���Ӏ3��
i��eQǙ5��Vvfe�N�Neʎ�p�V��������Nҙ!����QW2��,,U�(A5��r��2CEU�!����9�n�����&���5��k{(�)kZ�e0��)��.�廳��e�mk��=���7׆���TѠ���`�1;�hm�Q�ZH�]�4�\IV�-�v:�WX�c�9�5�Y��,�t�yz�T@m����+7l�:���o�Y����-�OX:���Ѻj�Dܫ�7/1�*��@{uM=�*U��dY�@�x-Yx�2佑,k���ц}d�mGrnm��h-�� 5У[X��5�FE5�5�:�he60`��K�X�e�475�ڻ�/]J�6f^+�Z�:���m0l�Z��s�渐Fe���^��QH�5x�a����sKяB0hֵ7����ڵl�$Q
�Z������SŮ������M���E2��w4U��R��\���>�B�ܲ�uT�&7H�e�T��h��!��U�&���QyJ�҇SGCW��h_u��ā�Iił�I��kX����:
Tsi���`�h�
Q�H&�<*�y�^�S�Y���+���֨v-�L,�.V�����4��	�Of�ϲ��:�5�����A���@#�uS6�S��oay����n�2�n��6�j5�m+�0���OZ�T��F��F����)�wC�Sq��G.���V��8�az��CGy�a[���̮ܪ7���M2/Of]Eu���2�:���wQ\���g�hX}��V�V+������? �kW>[ƊN� uw*Z1aA�c���.;��w������#T���m�QJ��/R��s�'*"M�e L[Cqn��;���i�D�E��?�k��<'S����6 ���-�8��X{y�*�˔�j�KS̖�kD��Z�,��4U6�4��3�z��M��I�FQ�u�oc�Jx�Pv�J���u*P#IzlmCZ��@k���y`�Z.��Fj�nA��4F��d��|^S�V�W+�m�2���d��{�,�j��h66�-��հ��F�-nZđ̼:�+n-ט�5j�jVc�� &�Mb����]��1��ܱ�e,-^�d�����.�C��qY9nU�8�o�Lia�6A�*�]����E|oP�-
��q������Pf$��U�HG��٥�-��N�S�X���}�i����FV�-T���ۂ����w�am��b�F�a�k_!�m6�l�f��#�0����ZW|ͱJ���d:ׯ�����Sn�ŭ�@��2�u�;��.d%���$�"X�V4B;[7=Q,�J&�6镈;�Dl����h�M�ZĶY�Q�*���匚�TA��@DVH���BHp#(V�̆�8A�a2�&4��2��Ss7�`�B�hld��F�Ur��L1U��Zm�f� ��Ù�mՊf�RkǍn��2��g�Q% 񍣌g��`�*��մL�6a��-V��ߤn�;�f�P�A%�̲&"&f<#uݚU��-��5n����F�$�<��W4q��bɓw�g�6��f�Вh��O��l�*��[M7� �̧��R� �Ukq6V���:�����u�c��yth3ؗ>�XB�J�Y��qE2P@L��Z�� �Y�r�E.����kK�!qP��U`�Nh`���U��L�	^�����j���ֈp����Wtv�I)�~� ���U�i��F��\f'x]�AQőeF��n��x��(u��q	K��&#E;%뷺��Xkn�~
���7T9X�U�̈́Ч((�@E͑T�(���Q��V��C���"[���V���2�P/f���7�ѩb��o
 ���Hhw� �G�x��޾u1̼�m�ԃ75m�N$��f��(,��L��]f��{SMZ��iP�V��72�jf��a�F�3�lzRt��y�Sj�(&Dƫh�-�� �Է��%�O�����"	"�hM�Vl")�h:/A�@6r6v�m�H�˹6;M��n����,�uL�d9�n�D������$12� Me�כZ�vv�)\�]�<�r�Ѓ��	ZY�Lҽ��5Սs6Ƅ�o5kJ��٩n�T`qe��`���)��z�7����w�*x
���-Z��o #*��L,Ij<�謵�iq4���v�x�Jj�l�R�f� �k+]IZ�*�\�J���]�CRi&�
��b�{5���`;Yq�j��J91�)�O1ph��G���Oowd�ڡr�mA�c�w�_oK�XB�mWc4Ζ043,�Z�һ ,x�BUEYOk1��;�ʺ�m���U��U��R��i����o�;�d�b�]R�� !0i��T�PC&����HS����ZS0��E�5�eKV��V�8j'P{j݅ti@m� ��9�Msc�i�7�DO-�J�u�:��
�)ׅ.�I��h��Mg@�A�R;�R߲��+h��̣�5S�5J
)��^h�nd�%,,k�ݚu��5���:�7zP�=b����p�6f�̫Y�����+3Lh�#Q�0���k���(���r�i���;����ܖ�LV�y""�̳lX�N;�6~�-�̼��l*��lf�e��¦݌���d��oG�)�	�2���+�H
��ė�MD(j��d��G��=�g�l�KZm$�im	]L�9��wPQ��/k��Ù֙"�3EX�8�r�j����fɷ�/w��
�7��S�S[һT��O���Gƒ����Գ�r�1[9�ҧ$6u�Fv)[P�oG���W�\�G0�����%�J՛��>��*Ŗ�=�=t�%=��bO=5\ȳ���P�z)^�+�9�5�:�@YkM�����e��լ"��M1��ݘ��v�[��{;�ҁ��E�Qj
R�b�̢1���T�)���*2�b�5(�*k��W����r+�l�Ke�P�395FQ鷬�OC3����YqX2R�|W�(���Ɯ�..L��x%>��θ�%\"�����+�z�����L秦����mI�p��C�%�?,�� 0���\�����:֠z]b�dN�[6�����Ç,��p��N]r�B�I��0J+c$��x��:ae�.�.=#G'ً�P�����ð��L���}��:oQ�
��0��b���N�Y�U�^)*p�Q�m���oSڀ�c���ÈlS�8@; �B�S��b5�	E�M��,9SE�õլ��{l��L&7[t��SP�"�[�x��7��c�r��SՖ�b����4Y�]}��Pk��v*��u�Ng'T�ǚ��a��{�����0����YI{�hw\���W��7��Y�ԡ��Зzn�ĺe�q;����5�̥�wM�=+V��n>08_6�ݎPu8 ξ�hs{���;W���ͼ�;�)���q��$�N;s>�aG\5���oJ]7
[�"ޥ�H:�u��#�6k@ �y+3�� ����W(n�5e�s:����7�Nr�8,*��zu�b�훀K��:��]q,�)05m�朣��w��dnjSQ�&1����߉��b�bD�x�^�SG	��7�Oy�,�%ӱ�E �<�M�7��iK�Ŗvy�20�hz)L;�k�m�W���v�X��lҧp-���,��+>�mJ����Z�77Usx�"��2)�ۄP�٬��[+��fn�`ŴC�/L[s{��Er_>)`�t@�d��M%�j.�86�q#8���qZ���+�Y����1n`�W$3u��6�j�E+z8�B�K�E|��m0f[��p.��v.ɢ����έX�&���5N�U��;;�5�2�S���|n��^�Y�ͺ��VνS�|x�>�(t������NO.��������3e*H�k�­"��W�ܫD[&��X���^$��vSr��n�OE��j�;
��kr�ǜp"M�ޭ������`/�
��L����U��n�����I�^~(�"�>�Pý5�fnR�O�O��OK�(�[����w$�#U�[[�bܮw�#�3�w�N�����N�tWzht?,9E��7`�V��d()f��R��WC�1y��F�v�o�+�v�;!7jl��rՅ�iRᵙǍ2���Q��듔Ӳ�:��y;{��C3��T�I2+U(�l�wv���\wk{r��� �lU��f!+b���斬$S'�4�LOq^��락����,0З���Q�}i^p�ӂ��ND^�v��Jٌ���� �h��EX@j8�f]@m�Y˴I;��$�DRp�y��N^�]�f�T���Q�Ԓ�}ʸ� ���.�1����N���	Ҧ�P���ʥ����d��Bu��θ0>k.�tA�����!����v�����3�)�X�GE*Η�mD&�����yq=|w0ݖL=m^�Z��e��7��
̉��d�2w�¹�GRr=3��]`X���E�鬈7
�r�:��mN�. ��3~I���1�CF�����ܮ������D�V�:�
���w��gK՝�u�ؽ/��Bʋ��iTE6٨֑��ė{b�F�az���*ξ��gʰ�.)cl�8���74ԉ�P��§tN4q���kUKl*��p�'BحUIe0�oX���Qj;�8jL�K�wcw�*f���ƾ*�^ps�p��*5e�vi^lJ2�9�WN(%+�+�����t�"`ܕ�2!=UQ�%������4���T�rt=�[�r�;	WwCl�Y���
��/���?���+�W���.� p��0�u$v�رs3y;���B[6_;��AWj�7���2Tx2�$7��H�ӜE9 �-K�ҭ�ٗ��BP�g;2�j��Uk���䚲�X�H��֋_ei���֕�+2>]kw�����om*h�VS�ܯ�B[C3nٺ��&����E�2�QqS��z��}]�P��^�Nmy�.�2�V֋`�d�O.W!)��wO+��JQcК��g��;�(Sy��ɥ�>ވn�m�v�gY�M���l9|v^����\-�k!\����]᷐�bM���i�k�Y�^C�A�J�Q��f�f����ڝ�Sv*e��4��%�e�x��j���O�f7��9�4�[L�ZcS��Ù�᡽w�АP嘣����w`�o X'����̎�]f
�f0�H��ᖍ�j��+�\5	*�,���#��/�-�,��Y�c��A`�ׇ#R^A�aŅ��ofEo�����yE�I3�PRV�p�&_�M�u[.^#���t+�p�l�M0ޡ�3%<�V����t�{t�9����R,Ep�)�!����ǯ�w�5�x�~Bu�N��Gq˖����<��BL�0`}�)<����MxTT��: ��e}wcS�X����մ����g��r��G2�5�t�����%Z�Ħ�kT+5>�`Q ��w�nł��(c�{��I_1f��Q˵�5W�������獜y;=�V#��!ո�5x�)4�cѤ�}����������Ŝ��Ԡ��K3�Ay�5D�s\�|ު����Z�7Y���Z����-ݒ���9K �v�}[���֍�fn�LU��yX.�d���՗5�z�\8�3K��Z͏��\�,Ε�͝g5r[T�8C�����.`iv��+�B4$���3.�BD{|$������-A��QAk��zA� a�NVBTh��,�8j���m��A�!�s�5��"��@������t�Jyvh�ΥA2��ܘ�)��4F�qzk,��w�]�7g�j@�H�O^�X�+�̰R*/��R�� ��3��͑�t��"L���,��8�櫣�2����W�;���ц�s��ňs2���d�=N_Ŗ�u�[{KqVYw�7Wq�5a�ka�;-�aoXɏ�e�m�O/ƆU�O�K�w�Y`�LD�����v�X��9mT�7�[�wH���e�&z��O�d�����n����:��,�ݿk	���֕d_4
��u��6�:�~��yMB!���Jf�C1Fq���OƖ��;��Hbk%m&�X�9]��f7�8�����w�-'k�M�o�Q�7,mA���b1X�%�������r6��c��c�+P]��'ew����e۰����T�����.ʱ�/j,�2�Kv�+x,cF�є۝��k��O.=9h�
ǜ]>f���q�Kԍ־�Mj����r�*�����ky���e<�����]F�7r^����c-ܥz�����.a)�:���v�oTQNs]�eu��v7��oV���ܿ U�����i����p^X�9���4p���&e�Z+yY$>� _Z��V��Ô�LT���`�X���w�)Aֽ�b̶)������^���L�0#��:�F���ٟ3�$Bs����6����3�V�s"ϛ5k�f��o��U43u-$,;�z�]@��K�]�h�:��gy.�y���,���Q�K�U�ۆ�9�J��}V�M� ��)�Ge����"W{'3*U�����odŜ�����ޡͩ�	5 Z]!�V���E ����u��=�7��F�C�  D쓉�;��R��٢�@pK��Xr��Ѣ+,Q�Y�]Et�eޝ`�L���WQ9)Q%ޚp��{�Sm�O����ۚya`s��b�֝�̨�'�d��nq��'D���.�6�K}�;�����6bO����@�K��6�.�u��M',�SYX6��C.���<<fJ%�Z���d���lz��8��[W��Vr��@n�H��؀�ud�a��J}�#[]��h5�A�"��U�����M�=��˟}ͩ�j�����iP��ua��6�����̛����w�G2�F�69P�VX��=�=0���N�cF�ɟX*I=j���fR9׆���ZWd\7N]gA$��0m�N�K�m,�gέ#X�2���������@:sC7*�G']�u���R���G`S�K��[/�[�yXdڝX�b��*��u�a��h*���*d!��H
�آ%��BW�E�M�ܩ�d�Z+�8�o�⾃<����^>�/�� wk5���`�
�����f��!�U���F���܊��*��js��S�N���Q��0�`5���5��{��:�b�`�(����=�u՝Vl�Y��ܠ�"���p
g@	�eeՆᭂ)`�ra�8�Y��@s����d���)L�h�o 9��[g"nn,�v��Ҍ�[v�ٝ���]�)4Hi�Ы���
U����ջ�wv��e�@Q`��W�XS�m��Q�#�8sw*(�$�y[�^޺��٬��!��.��9���­�+X�]�V2ˬ��=
(z�E�u��0��/�xi-wO9�H�q:o]v��J�?.�+b�Q#/S��}�^�;x	��Wg���:ވ�
{���x���X7 k�m���3���XDo�)����.a��*��Vۘ�ҫ�;�D��z�m���V����	â�#R�s�*�%����3���������ͮt%d��@�k-`�+��Z�����a�ns'��Z���/����#�{)��18�,��~�B�r�l�*w���p����ƛ�1\$S��� �����?-Q��Y������U�k~��2*fH)�gR�GkM�|���e-���W�oPt�9�Ɩ�<⬍�xj��#�����.�i�<[�
Em�6�vզ%7�!����6^��v�UB�V���Y�v��o�ا�會o�)Q��1E�v�d�;�5��#o�or�5V��^ ��������|�2�#`�Z�d�׉:{�r�
�$��>YH�mD�TծC����vv"e��m;w�6a�4��tƝ��b�cJ1|ݱr��t�ɫG[lL}��`vs����E<�r<�-�3�n���)Y�T�re�ml��TѐdN�S����Q���r{0ݔxv���yCt�O1��	�m+��T����Ɖi�v���+���NvV��6����WY�[NI�1��rgm��}�P�1����w�Yb��h�|��s�U��YR�._��:���%$8ߌ�f�[h+j�d�)U��GO����[�s�j�&>�z�y�S*��-�M&';E�\&�CJnd�ۛvNf��I�i�
}7�	-"9^u�c��P_l��� ��k��#�8-B��;�c���R,��.itgLJ^L�/�b<�Pȕe��.�E:����Ă�a�նЛ��	��=�֌ss�o�c �3�׵I�7y�"
��fn�ç����t��[G��&j�xN������	�FuA���#����Tx�.���B&��R�o�P6��I��(�q�ouI��a02�����if0!�BO��F���Ρ����v"�4Y3i�.�8�ӆT[Z:����.�[�8�����ŋ�4���4J�y�E�x]���7�O���J�8�L|�t���]wܵnd�J9�A�U��k���W+Yu I��c�ͭ�i�V83m�Y[9^[볳q>jF�+�q̥��+L��Ԣp�$�g `��c�qК35���gm�Mwv���;�ՙ:mW�{�e�}���Vg\�7�|���"�m�R��
�Ի&$n�9�B�aܳ@�<�ob7�[4����X޻P��CT��#�@HF�U���S=�PHe��%ʵN�ř�^�Te_�`��M�o5��o8Vtm����ى�ɶ���ը��C6�}\o������`�f����ջV.K�I�ȉ�]��.�f�W�Ŝ��3V����l�`_�-�I�IZ�h�bk^���ʒo��D�cV�F����xi���ƈ$q�U�֒�&��OZ)��ڝF����*]teLv(�
JKMg,}�!���&ێuu҉��ˡl�Ip^��ς0�d�)_M�N��%,��\��u�Y�۠�;�;R�OMͦ���	�P������Y�#��}v�vF��s/�g^qJo	&"5�\U����í�[�x.M`�����C���+v�.�Ֆ��*&��F��Y�{vs�P�-�T_U�N����ux.��.H����6�6�[�vq�@S
谦������eʶ�B�c�Uə���@���7"����w�GV���w ��Qk��ӭp�k����G���;��iХ�@(kY�C�}E����v�Ř�.���!78��C8��T07��f�Ɍ���C1uВ̜�֪@V�j9�ˏKWZҫ�����(�s6�Z�TN������%�5���q�:I���c��b^�n>��2��+�N�%)(�=Chn��̏5j�Uғ��i��*��6TPh�]�9�p�sI��IcVo��G��ۚ��^{���I���BH@�~=�՞q¿/�
�F!�U��[��+-�}��.7+�ؔ��;&Q�=k#]]��i7�����[�ܺژ;C����n_݇"���3f�)�]�b������<i�@�R�����,��x{/�Ԩin�d�[���L}�Q���M�����a.�-��'TI�J�y��]Z�Tk y����8�:��n1n���No�/"����w������tQ��L���q�]f�b�o�r/`@v�wW�ރ�d�qV'�k=s��y���}����eC|�'�%��fӌ}nd���W�z�� �L���	yA��m=&�t�[�7��8U��Ɋ6m�#GHp8�`m�y�t�1:QJfYׁb#��vU�g���H��w���bK�:�fd�Y���4��M�wLU��/:�K�|ɬ�}�T܎lH�+X1�I(��d�8_Qt����Y��e���m�ʰgi$�ǜ�6�슳��R�S��Yy��:�.X��_+�q��Y����0k��H�o�w E���.�Y,�
����Eے��g����oD�R�>A�^��g*�teq�^'�t/"s �RA��5qJᮻ;Cp��C��x����Z�X�H�x��(0gK��)k����)�[mV�S��+r���#�q�䴴q�	Ti�{tu�;-�9�i�ɏ��w�1V��5�D�Z�O�-ӷIg��ݦ6_U���2뺡�YS�V�h�u�Ԧ*�tF�Rit5jngG��� �I�rN����,Hz�����t[�Q�Cd���ZM�$6�f�G/Nhc�����e�ʷ�=wIaY�ҹ����I�����;��}���U�̓7�譾"��YZ3ss�蕦�큈h�,�6r�h��)�Y��2��'���|J�/��<��:J����9��d+
���,�r��Z��AvWԲ�Vfǘ*
J�6�L��K��`��^uX�笡����hu����3��-lN�S�e����nX��f2��-�ܽzw[q;�ٟD�F�B�COS�
�1wP���;Z�Y�Q$䔫h,�d�k+��G\o�[1T�;�n�sF��CM�G`��-Yusm������ND��%ܺE�����5��Ń|��o
	}�gF%�\5�����A��QIP�%��/7p�r��J�[[
�t+hQY@:��2G�&#!SB	w(��:n��"ۛ�j�5��]v��Mf��p�0�3i��ܴ_|ܾt��%']��7�)���L��]�f�s]u���\{�8Vљ҈�gv��H;i�B�hqL��7���t\�k�� 1��Zu�q���h4���M�/���6�$7���/�M���L����@ނoV��+�:�=5��ԓ$�S���;7��a��w��A�&����)I��񗕴N4L��$�̓Ľ ��!!o� /.���#�rf�T.�e��wʭ�y��mފ�4Y=)ij����a�HͶF���jGٴfv3�ER4;��F�v˦�K,�]0��G;k��\;t������ ��&�}.��^�a�m��-�+8٭1��;x�b7�~r���iIB�r��P<9J��Mu^�Ve��tDR�r�c359@̫���$$Ѹ׊۪�؍e�ow#5%֜tN��q]���t������dz�ֻJJ�^�Է��}O���5W�$DfB���9�J&�gk1���%ˡc�v�N]}Q�삸��ՏG���b�7~Y�G]9���0��B�"��us( �D�n�� �=�iQ��t���)�]��,��CC5�w�1�=lN���c���J���g�����t: S�q�9+�@�o�,$ֆ�d����w�&xK�L�(_�ζM�ی]��kCV�SXx�<kQ�0^\)Xs{iLz���'N�X�ޥ�dTث���tt�T�˭n�>�嫾�V��*Mw��/�V����eu:j��<ڙ���B6���!�e
;��ŧ�>��raS\��v�At3�$�����"Yy�+�XYugq}����ME[j���ԫ���7�5�t���E5Ҧ=�����\���"J�ݸ�6 ۳�&x��)�f#�<�V|"|��N�(�f��u8���,�V�+�Yȩ�f1��-ַ�q�w8��Awٝ�	͂�	&�R�W���u���'�j��ٵ��Z���Nˤ5���+`�u�j�[�Bp�
��sM�� c�a���u�n;�a��fH$e��i<��C0���'�>c��]�\�x,�Vl���&��K��%8$:�M�:�;w7�:EbF��V�ʝk�"�fǵ��3M
QR}�R���Z���Y�}�%�LD�*���� �>��%H7���Q�s�.Fk�sޮS/Gi������x-J��(�4f�I�l��IK�ƛ�;HR�(`kr�C��r��z��3��v��=��Ļ��4��S�5���Gf����Z"���D7�$�i�TYWʷv����G�j��Ė�q�T��GG}��,����O�
yY��n��H��Z�#5V+6l����V�+�wկ���U�r���a�Ef4�A�V��؉�����k-
���4��-.�
�S�ť�V�eC.�Z��V��89WT�R������VD��7dv�-k�Эn!$r�n[�WnB����@�v˺Wsc���w�\ǲ��l5�Rƪ���$3,N�H���ʏ �B��;�H������+���2���Ʀ��j�'2G��eؓ�Nz�c���"�+Q�7��[��*�eX����kݳe=/v@�Q�jZ�w%��iT�z���jǽ���Z�uXyzy�τ�֔�k�Fpb�-h����qQSla��.��Q�;�XO�H�B�%�!R+n--ԁ��G�u�5�0�Z�9z�N�ˎ�1*ˈ�Y%�4(��W����Z1[}�h3���ޑE/�]�RpXGin�۴��Q��&n���j�[ˤ�'���w8U��n��v�I�i���ܮُU��� ?!"R�ڤ���p]ڡ��r�����U�r�ZGX[����ʳ��=����o
J�U���;��I<��lWq|��9@l��ӆ�Y��wC�xsZ����]�˜2��B�@`m��WN�h|jU�����, Kn��"2Y��ߕ1j�]��)�ز�����f�8��ғH�kI��hp����� ���L�ֱ��TCTsZ�X{�L_���	��n"7�J|�����:�`ÂQ6+�y׉�&��PweC,���2�F.�\��cn\��nh8��B����t��ND5�v��E�u�mKl1Ty�8E�ӳ+jR�ƻ�� 'J΅ˋ�wf�+.�⚓Ky)殧\�`g�Ὣn��ݲ�s��e�C[ڹ��1�nB9�a�ln��PG1ȟ4愜:�\���� ���/���t�����b
C{e�-LF�e6�{�P%wCE�j�yr���^��ŕ���-�[����VM��	�=���%��\�]��]����q�N�-�7�n+�}�V�IՆ��s]�7q#��kf�+�$ �36�6���'L���6 �W���Ş7�+��u|<y`�3ki�ȶ��Ɂ�&��BVԵ[�nn�\�9��X�-��$�)dV���*f�c4�/�m#{12K�T��VL�ݡ��r���JE]�$/��{2�b�4�b���)d�����.���P�-�G���O�⬜��cV<���<U�{��,de�ş+N�[*AY���J:�m�����K�v�/��1$c��,�\�담�ۤ%�b�v�to�4����GN!+3eDUL�֫ԟ���[М�L6Шj�F}��#r�o:J��C�2w_�ާ�O%v+��|�R髧���9��W3Y!�.��ۊ�Ғ�t�U�s5�ї-�c�O��{Gl�G�m�{)��Z�ٽr1�VLn^t��=DZ�� �c�=��q�*]MU֠dEt��Ys��te�eh��8u�ǐ��>���m)�i%%;�ͻ���2<��R�B.�z�tB����K��Uu�)g-��f?g	Gozj%�M�`^�X�a�Q��(f�@;�SM�X���':�t�M �b@��XEM'*��� ˒�J�K7��)���;#��n�:�q�]�;�+b@֪tuMx�V^�ox�uj�[����2���wn.@��x�c}t�d�`Tc�b�V�� :�b��6;9}ہa�ޝ���z1m].x���Z)�Y4hg&�O8�f���\��v�f@��*+mĬ�0��4�=����#��0�v�X���!�y��{.�R�u�Q9B������Ђ0�9�a���go���yz�IJE%E���r��3���?����LhJ٬UC�
>s'"��sP���Ul�gkI9m�+�Q`�ή�J��kU��8�rWC�c���VU��N��k��R��ڒ�Fi̤̕r�\��
������l��ٗ��'jpԅv�̂�f��hp[Xr�%u�]�Rp�\��j_c�y�r3{��0^�R(X�q�����ҡ���Z Q}�b�3��Cxs8,R�pL����"�Z�Ե��C��6��u��^�C�(ռ��W�^�������2��x��<+7�o嶮)�5>��7
�yK7�Eq>8�b��x^N�6V%�KAT�wz�̐�0Dڗ[wX�Gp�t�t�a̫]��6�;Y�D����b��ɀ�G��9�[.�:�M����)K&��e������S�J	�kY�[���ڝK�`��鉘2i͖e`�}g^!��Z�gN���)h��ˤy=�Qnjb����w
;��J�`b�/+�u�yds��8-X"�?��+t�a�\{��8e�]�d���n�����h��X�a.({��VPx�n�=}s�I�Y��f���QA�4��}L&ҽ]�q�-�X�/���GA��ǜ�q�A�6���;R8e�f���R�r*Zl�y[|V��z8Jx��C��[4��_��Q������R������AyV�{z�i��q�9�+��j�� 0'����x��$�WƱ���L�k�ʺ3nP�Ϻ.ϭ�to�)�m�9M#�4�f�a���9�NɄ,�)�`__#Z+��׊h���:�(h��`��&���`�v���]n�K��1�ʼ#�@�7D�p��j��;DQ���|YKr���וyf�=����}��w�H6�9|����qZ��F�Ulj�MNLD�����/��S5�[�N�v���fڤA� P��TQ��e#���s�b�]gQ��!U�t��%G����z/P����Ev�0�����P���܂�݇w�� Z�=�̕��/6U���w:ʬ�urC��b�UɋY���á��m�#��U���=	�e]��8*_d"��\W8�7������X����R����:v��^�����1},v�|87w�t�8���-��]^+��X�{��&���/�V����P�B���ښ$��j;cp���W'X���{d���g�LZ蟁GU�<_Y�ۍ]KyJ�n,��0�?q{([��̤���J�q�)n N���mt��br0Q��\����0V��x;(�݅ݼ�
-_D�*f��,>Cyc5�y�w�f�;�6�����G�T;�=Ú�d����V\e+^� �ooV]����61ۃ�=uz�S+��Unk�(蕋�.!W[��s}n��g9���Q3�nv�f�N����{�W��Khq���t�GZ�U��P6:%��$�:�9(=�k �G�������rHꔌ�6���v#�e�g/u�嵃kS��vu�#wʠ��J1z�XC�N���Fm��DX�B���C��b�KNhw2ZI�ʌ��B%��a-����ջ�ot6�v��{�l}5L|�q�p`�ݑ�QU�D�o���1кKp]�\�J0MI]r&��V���}���u��y�%	 ����]�/����7��q2�2���=��k��D��[ܜ�m�Gp_g�.(r#��w+e�֢��(�w3nv8���Ѣ�k�]���G���A#W����eZ�Vܔ�?�5�GgĿ2m_��aѴ�9S!��_Y31��/�bfGM�['������0#�39� �s�w#:8)�B�Y����)vqm7��(�[K��xԭ:Ih�[9�tލ��y�b��,����㹔f��Sh�ǆsK���\�w����sd�{�7���(��j �
�o�[ih�|���j]��ݙ#�?&m�[Ϛ��XJ��u
��&���Yq5���E��c�X4����ʩNR*sF%�dڟm��ꛈ�m��/\N��B2	گ���[u�s�Jl���y��aq�q����n�PG��`�Mm�x��H���*^�=Ϡ uu����J2fF�cǎ#u����M���uZx�{Q�w<�t��H�utԫRYP��!{��F�ن�6ܡtÎ��@���P����^��d�syգ�����t^j��p��geS�w���rWGc'k�ػ����Cb�}C�wjt{um��14�=4�#r�����h+�^�{���eä�o�i�I�2����a-^bz;�r�Fhy���J�aC;+/�uZ�{S�#$�aɔ�:��Nv��v��Nݤr�����Z�q�3��4w7%�A�H�|Q/�.�%��vw+�}�k�����}g��l�vÂ�j҈	��bY��u�ʗՊ�x$���h2*��::耳3W����Uq������X�j���^�шF�����gK8��Z��̱�	�
��T�$���_޷Y~��|y������$�/�s�N
�{\�AX�;`Q�U֣޷n�7P9x*_X�bc�3����|���* _�a��s�@���li�۵:M�t�����\֏i6eݭ
:8 9tr����}��XbX�n�w��Żq�Ʈ���O[=c3������4i �]�P��)G��ii�WF�c�8G�&�@��ܬMp܂�s�ٍ��[�Y��sJy¬�ɡ��v��"�Yu{u���v���W�4��]�ۏ/(�̧��$e�$%U����u�#��Jiѧ�u0ܻu䧎Mz�
���e�І�Cͻ���OW=ts��&Lʷ4�dq5�wt�L����v�x�^,Wu���5�e3�.o1P_^8�-�t�6�a�d�|��bv�HpY��T,�8�Z�1����F�\Xb����ز�$;
<gMm�0�[�Օy�x���ɿ��w���g^F;�����Yd'M�Y��������HL�9e����HNU�v� �ɮ�2c���nMjT�]���Ҥp�,�yXv���'����(d�Ӂ�9N�t�g�p��`	��t8�y2���Է*u���F-���[) ��+V����;��Z�7+*���v�i����ڷ\�Ǒ-[v���_\��R���C��Pn+@�=����"MK���x���b��P0���
BUF��y��^W����ۥIA
ѵ�l��-T�1���V[Ach��[V�0��T(�J%�FԴ��-YEV���ڢ�mR�Q��-�%�ň�bԬ�hō�TKJ�ce*�-��-����+YX�e���֭(UV*��iZ�PF��T��QDZ� ��T*���1TF�kZ�FEU+D��Ҋ�������Km���eH�V��QTF#Z֠*)B�T[j*�Z
UQEJ�QPX,b(�����TF1J��-
֪�-h�[[T*2�R�ZکkmeQUKeV(�
Z�V*T�ւ%��ֶ[V����j4*�*��)l-����(�j+m�b��֢�l[A)P�ETQT����(���FZ�Kh�+Z1m[Q`�FKA�%�J0m��F*��j%���ڟ��%�kP�s%G#Z�̩q,X��T*�c�E9j,�X�h��ie�*�U�Cd�ΦRf�}������H��a��;��1�n���!�u)�57��0@E�9��YW�8��;��ۯ�/7����+�Pu��4�?��'����ņ2�c�N�3ѱ�1u���~�5��v�)N-�O{5���y{���t��tn����N�{K�����f	�B�Q��L\Ҷ�'��]�X=~B�i���6���x�ܱ��Q�'a�<�t�E���嫚vŜkM�[�����x}k�����@�č��#��>E;�}��w\�K�e�e�S��q||�z�\,�G����Jk�
ZF;v8�V��la��}���x7���}[�p����Ï�5K����j�W�ƁLv�����.:��&�V�]�*��-�ꞧ�t�B϶��\u�M�ù���d^��S{+��vۛ��l�n���۞�3�}4��p�,oO��©9��yn/=�x��U���wQ���!n�߂	x� @3c�=��������_�k����}>Uc�I���K�9x��⑙Qi"88��n�mm+�{P����f�ҭ-�`L�	{��j�rӡ�{���5���D�Ξ�AL�"���KgU��L�9�^�Y���L���
���5���x�8��v��5�˄n;�F��1usP�m��tFm�;
�ֹ�;	`d)Rl(��W}g"d�s@|g��+���6n��`�ݾ:`sbK�7�w����m�NI�*���B��yaތ�f�A�dl�=�*����c5X�!ޖ�j��.��L���Υ����HB	���[��z��r-֜ڳ�3����\�_]�EGF�!G�^�c��{Y,z�'�2����N^[�}3���,cN�x�Ι�:=!j)�o��+����j���M���}� �V��)�ҏ�h��f'��$�*�hntbf��CE�;�͒I(���65(1CX$@k��7������W�dc{�Z��[B/u�Ė�Ѱzf��;U�ӌ�����`��|���[Yp����=Aw#�%-�*E���W�x�N�ed��L������A�?�f�3j�ޝ9�=����YrZt�o]�E��\�������_{����3�b2D5|�\]+4f�n[���>��L~�J3�Qr3��ʋ��݅����q���Fy��
T�6szU@p�;�/&��O�\<6��tŞ�@j�5�k��U��b��t��,9�S�|jm���CD/H�e{{�.����,��N�B-/J܂�>CoA�c��՚c5��"�R����ab*5��5������gd���LF�=�l���|Q��t�j��4�)��q�n���[�"̧��of�����C���퇤�ufI������T�Z��٣ܾu�����]q�_o�B����L�o�I����f��g���~�t�i������Ĩ}�3b��s�>�۱�Y�v���=��j�=-�yo�8��>�0+ú�ĺMv���9#���kܧ�l�?q�s�Ӄ�36C�W	U5a����p��T��m�>.�.�W��嶳ְy�W�I�����a%f(��9(�b���o�A�`n�B�yH��1G�������gH�o�f��*����o�%nO.<�Qs�0M9�]K$�赞ٰb�:�����&�[��u�:�nj.L�]Ot��Ù5����'MX{E�"������K<�Kk�.��gÞ(�7l�O=g�[I�a��;����GrԷ�4�l;���f<��4L�si��
�oV
��2v�S*r��>о޹��Xꩋ���qĴ����}`�a�@h9((t��ƞּ�V_ⴛ*�����8�0X�;S#Z�Qo>�k�#�O��2~�a6�����]�0�����]׸�w�V
�~N�=�P�r�j�d0:>N�S�CWd3]r�=1�ɲ��@2��54��e��M�r`Ϋ ����nr�2�����vrN�A�W���_E��w��I�"3-�.�ˇT��5���f�\#�9-.GK���1b��|�������uwӼ!���(|/����2��I���u�|��M��9/�X.�V�QY�5У	׉��Jn���)�@Mx�[�~�\X�\���.�F���~7��z�#��p�@�^����n��Y�Z�y+=��ml�����B����`�9�>��#j�z�C�*&/e���O��q�����a�&^��kp�P���GQ��zs��T��o$]�#F�w0䫘�:w��3raM\䟞Ty����g���F�uA���ψ�п��|jஇVo������S81���r^�]re��M�n���J7�Ɓ.=!mp���S���]����B�Y�b�� �~��m�FɏpZ_�J��~�6�YKܸH���Gdv'i��I_^�d<`j7U3բ���ԬO;r���ݍ�qў�B�`�G�bܔݨ�s�p��L^��p�%�/�m��v�*�1t��÷���e��6�fM��Ձ���ڃ�&���:� M����.�*&�:o�g]L�\�R�|L�p����������P�c��3��bFb9\��(����v�����^ro@.�m	�wV�T�3j��6Lv�a���c�NX�[o�؁�*����\��uJ�6-e�od��[�l���z�s
ĎqW��2��u��-�\�G�2��:}VW�1�W��%w8�%��Qnl[4�����q�scma��V�,v�*��������+a;�1ovzy4v
xRԁٶ���ٷ.@�$�B�<	�p���F��ꆕ�*Aa�)�FUM����8>�� �poO�,xU�hz�w-��]сfƼ3 �v1�:w�Nm���5��s���\��=��ƘV"�
te|؇�+z����Q�1��*����yOG��/��S���;��l�G�9������/��2]P�<�ia���c�W�P��T��~;�5����1��a4EOS���8B���P����4�q����m5cS�x�kEŴ��R��a�2��wOs`�w�$fˍ�J�t ��l��L�����Kf�
eK׮�B�g�t���S�����<�År㧪�5ӝ���CPȵ�`��r�-s�!V=]�3D�V����R��k�u"�N��<h�i�Ln�M�}���/1w��]L(��}9�{:����w�>:�Á�j��M[��"=�{Z���Y�Mb`:9���eҀ��Ͻ�be�h�as6&K����@�G�4�̚2a�b|gf��UƆ`�@��]�5�����(gsH1-ȥj�~��j���]dm�U���8�^{�㑞*�Е=�о��f�)a�����,3��H�Y4χ��0M)[J�=����';���9��Q�6<>~�qر�Y�{ˌ�Z�e�wr�����4%xf���6 ��v�ՑS�1g���}仕��L�9/����nQC��אt7`ŀ�e�c�(9�vN�5����L�g;�M��Y���.���P�S�E}q�!�Q�k<��F6ltfF��o�P��V�M���87�N���~>;�(�G��S����BS�Un^������ZpthmY�Z�E�5v�Oc�k�EΏU�\����tpp�?>d���1c'�=~s�uM�����Zŭ�����V�@�~KTX�k�$N�4���r��^�!��')�?E��&�y�Ҏ�}M�7k���J�Ȱ[[�#�!���JP�H@_�%Qu7ӄ���hd��d�(离�wi�/Y���~�)��-L��k��Y���T��iO��`��*�r�Ư8��ј~F���=��s����`�ÞI�b�h��Zz�����FI&uūI�̓����jm-_s���NF�s# R5�h�X3��75�o�]'^C[�(͖_��ۮI;�"���1�Z��"*�n��s���:�fȻ��9v��,�ْ&�gN)�"��6aތy�i�L�\��ī�/w>*�L6mC/9���Wt%z��ζ���N�`�J�՝-�t��}Z{_VZ�ú����r�Á��8&ӮQ�����۲L$Q��j֎+�Q}�����*.B�A\�L�2y�ʄ�j���J�$ͯ��>A8-�i���Tj�i������4����DW/Nb������X�9����v����{*�~�CB���p<�A��'�o#b��_U����{/t^h㦰N�}�.�yG՜��[���<�*}�d4]��T xCI�w&|E�Ҭ�u	bk���c�L�qJaT����J7�ƀ�{)�c��Ĩ�����4kB�XΜ��Fp��>���c�I���n�h����S�}�q�������Ӿ��U���� ��EWӀx�^�\�~հ-5د�߁R���*�Ĥ[��y:W�<��"���r�q�8ܝ�hf�KW��^�!���W����z��l�1`c�(��x�J-ˋN��7�+4<Å��˩�6�/�z�]���9Z�$�Z#��n�r֡y��������Ɲ3���Fv�".��u>n�VU��b����;�4�)+_3&4�)Á������'MXK��
}Љr���m^2�����q/4�;���[����[���F�.p������H�՟
�D#�uZh�3]��o����{Up�|o4�\ae�%{����N��;�TL�n�TF��0���1I�9��j;�V�+;q����)���yMd�B��Y�|��K٘1���Q���t{D�v�C&R�0���rk�(���eB6Ӌ|�/rӽ�Q!|��Z;�'��8��O"���bRi?a�� �a���J�C����غ�N����x�7��ע��ñ������eܫ��U��q���%7���]�t(�u�s�!)��t9�'[ww:
�ք�H�JYR�l�E�	�Ȭ4o��HUn;9z^r�ϯ�m��!�Z�C�xB���5Fϵ�}��5y0`���
�zCHڹ�zhd����nvr���f^��a$4�.������w�lN�>J;<?#ӝ4�\T=�A�ńx4mlt�P�d�G��ITa��{5~޳�D(���#U:����A�C�'��>�a���@T�x�n�-[,���KI���v��澭kt�P-���k}X�k���e��TLYyN`���u�ʇF�a�d�:j�Q<�m�o���X:���%ME6lA�h�A�t��j��ò@��*h
V��r�o��#w9h���J#f��MO�O$;,�s{��6
�i�nt�yC�,7A���bR����%?vW�ɷ��b��2C.�C,ᾭ:}�pZ_+{��b���p�;��j;#e�e1�V`[�J1��(3{�Ov���^��4,��U��|l��PP��\~�k��e���T���-Y�f{T�E�x��h�P~�P��[?.)Z�m���Zm�"�XC�XD�lֻ߲�t;j2]^*��4����3Jv:͈��?y.��3��U;�z��Ø�h�9e���S�7�lز�@m��t��u@�ᱲV�,v�+�1�����5uyʔ�\�wK�{%r6�p�~ɤ�=�nT�*I�!cv$��k��lO`+J�`�d��F���r���P�����&�L8P��շ:�r�@Y�xfA��c�+\���0��WۼW%�wX�_�ƘV"֙�lC������9��{��Xn\�d�ds=�+uc���+�cņ{ŀ�}�O}�b���L�	e�zϟ!88=�^�Ƭ�{��&z���iY8�&]����r3�tkv7��4�ƕ�!�9��7�V�^H��;Q^
h����0��3G:�A�{��2�/��՞૕& ��em�fԐ��^G+=�i��C7K��v�5U�c_��LXk�8ݫ�;<��!j�*��Uw���a�ș&+�+;���h�^�V�z8Br�w�ySG(���Ռ��&�Ft���T�iFP�g��.[�CN�OS����ua��?S�ÝR�\̵��{������P�qHŹ[>���MLS�r�q�S�]�\,�>��5�ӫ��S��fl�3�dXkj�����sX�'oG]44��I�c�c�C25K���#U���~�ƁK;~��i]���_�N�v��
Ŋ�W/.��u����G8�^W�FS�ؕ=@AD�P^ô�p?1��]G�=����z>&��4�Ү
�������Nv%�w��\%eH|�Q��;�g��^��c�z��aΌ�����x6f���V��Z6)��U�	9}��LՈ2�_����+�Z�W:¡p���W�;-�f�ʼL׾�V��C0&F|��z��y)f�X_��ӱu$@~�A�XQ��WM��{]`�u�U��Z�s�A�ӊ����wy�Q�;Aҫr&6�C�����V�[�a9�N��ޜ�b����L�uav��&Vh�]a�o6�h���7L�)۾��t��E�,�����<asOmq�\�*����g�%��8F�� wwiv�(^_����j��nE5ֻn�3j�i�Ψ`[ݚ5�Q��v+c��� ��,��`@v�S1�ĔKS�j�'�B�7x��� L�y
NI�.4�mv���V�]�)�2�����[@VWe���x��ݒ�7]�{��)en�5PŜ��	�m�'�.�C\�މ��۠�Jt�u�C0��(�0��Ø���Y��+9L�����^gwҭkd��F��vQ���@Ϸ�f�ޡ�8��u)���˩}c{k�ˡPdtCZ��.�63�g7��.f��V���f�>u�hI[��Q#��t�@�]�Έ��ڈf��d�s*di�3/�}:�)h��jz����z������v�Wkp<VG����P�mP�R����L��l8@�f�V�(���+�$���xo.���W�bjA���Ǜ���a����n���L���jR�G�k_<�T��n�M��$��Wv�+�KwiM�Nm��xc����]���'�*���\���[ߋ7��q7�@tè���P��Ɗ��Y5>w��A��f�}������K�N2sPj�o]bf'�7Q���rAP�i���=b���q郈mu�d��AᕟF���yB�av�w.Wf���=��헜29C74�*�$��\�����Յ�h��0���5��6������d��ݖ��g��3���f���v�Km�\�2�ڴ��z�,�,
�E�hamnGn���$�w���U#�M��X�a5[S��m*P�;�mJ7�����m�[z/F��uq��n������#��b��t%\�+�6��7ѺxU�sen�Y�,e�aOS�}�)
́L<+��Z�IX��d@h�-iו��c�WҒ��h��afӍ�6]o-$��n�;5�
�v4o*<��-�+{c�_��>�y:�c�jf����<'�۾8T��I���LYFd�w���t��N����y\K��ܬ�~�x[��86������ڤ,fiNP�S���0�i˭#d45�NB�Y6�4YY\U^:�hM�Ԫ�(�N]	hr���Q��Z�T����{+B4�����\�yd���f�#p5 �`����u}��O*0"��7���s��"p@��"�j�n�A�i������əP��V�ApV[��9ZH��V֎�<N,p�[6��KKv��iӮ=Y�3����5^.���щ��?1�m9xL���_�b���؟Ƶ ��ݫ�)|L��jK8��̙&rY�E�r�#3��z��(���a����D��q�l�t� �ը>��-�2��p5��KM�e��v���h����V���fo�ytf�lI�EO��A�ւ�m�#l���ETm�"b*���e��TU�UĪTb��KE0�2�kbe�b��4q����m�Q�TU�0�
�TS-V.Z(6�1mQ��UU�UmhTZ����-��ұ\nYG-D�m(��Rԩmq��kUH�̘���*!Z�!k�m����m1�QƊ+KU33"�j�����(֊�̮%m�h���F�+��kF&2�k��-�Q+AQEf&"-a�c��m�QATEcYTc��-�J5Eb��ۊe��-iU�kˉcl���ڢ�W2-�DUTDb���-E�+�F�X��Z��J�K*�V�*���P����Ecc��EZ[�PS2�-*��+�Jbe�EƉ�UEm�5�Ek���
�UDE-R��QrҲ�Ū
%K"E�V2�Uq
���7��\������5�epr�=b�7�}&��9tt����mNV���G��+�:*�*��2ɻ��<�[��"�*��������;�lϏ�3JCo@�֞5�!�Yn�-��R���Oz��e-7�J��l�Z�\OM�a�8p�EE��^�~;c��zO*�����8�!���o98�7�m���D-�ы	�W��3�l�&5*k��, 5�%bo�T؞�������i�%�v���&)B��`�ʤ�R3�A�B|�p;O
�\�x1���4�C�����{m$�}�S��j�q�ѳ�ߎ�:�)��|���+�/��W�2��r(�����{���	�N�:���
L�:[�r�]!o<�;�g��ژ;ŅP)N:�.������oV�Y:�i�Sp�Q��r�A���K�W��Y9L�8��%�bfk��Y�Z�dݎ�樂�jN�4�:@묨Y�_W$�~�ѮR�Q�JNr�c�LŜ]v�]�6��=z"��E��@w�b��5V��~6h�/����C���Nu-��=,�J;��n�E6挡:����u��:R4�t���@}�S6+���!���6lK���L��~f�3h�^�w�-��`�.��@7r�ڭ�]�fg�q�2
�2J��T+��j$ l#c6n_5�KEvW�r&��骕�ħ��Ә��ț:/���sc�d�ŽZ�������!9(��Eu��Y����jG[ݽ�Cy��j!Wn�ų�{)��{fKQYSl�����s�"�ma�V�:W�&leo<WR�p<���ú�ch*���y�p�K"���W�{*;�j�թ�k������P�uv�������2�6�^!g��x�zӵ��V�
n�]���g_sI.r��Tg��i�o�������4��?���=�oe������Lj�trL�c�s=�_�?b{a��&9١�TTA��Ui�=�+O���'W�[�.��9�zLS�K�ٙ��^�+�����z��F ��w�t`(�/w��0���%q9��sh�17 ��!^u}��Xꩋ�#��~��T c_X#=�+/�#Aڗ�!xVț�����`z`�S�:g�b�.t�A���<�U�-#��0j��w
���2�y��FR���<a��8(҉�a��g�qQ���uN�����jګoj q��R�e�l��+{iTdj��%��ƀ�
.��B�q�r�HJr2�r��=�>������/D*CO�N�#���x��U��J<��}[��ȼ9i/�������5tb��'J���V!z�Te�:���nuj[�9�3m�bD,f񬶧XaC1��X�.���ؽ�&S��V�z��V���)��o:�"�|�u�l����ʁ/Ih��8J|��Hˑ���:=���.7X
��V�wA�lΕ{F�S ��#�8��/=���v&���K�E��x�<k,_�����ՙ<���F�1�O�L<��N�f
� ;������q���}K|_ȼ8+'�dV^5��H�?�������4�ܴ�����5BuA���п��|j�v�U7n����T�͐{K<��;�s�67k�V�8��%�cD���R�U���l;��w�����a\"k��w_���ܡgϟ�n�A8ֹc[��t��T�:qKWZyu�w��2E{|��wJ��xPe�hՇѻwo��}N�Vc���u�Ba���W�]�Ď+�e��F5�8�1z���ǒ���_8�����e��,KY�n���H�?I�+�{��\�N�㵝+.j��)�#��Չ�PPQP6���Ը�)tn]_�$�7�t�_�Mz��N�
.�n�;V��g�|d�jv�T��*�A�(ydWYZ7�(�yo��v��[ ]��)h�>㬻���}Lu�;�0C�1�6�9���[�֣p��jz�I5�I���[��Y2�;��'��a���,@F;�ᙙ)nɍ�p{ʪ����R��Rģɘ/�Q;�k�ddQڭ�h"N�(*�� <'���szr:}���G���2i�͛r�g�E)9�Xǉ�q��o��lYX����u�����$xW�5��n��J��|�7$Z��T�׆d��q'2���:��}�I���Y{E_�gT4V���ú���,�Q��׊2�gҮ�i�{�Ek�[����dl{����T�}�|~�+OU
�]P��,0�L��Ď��Ky��R�!d���0��{�9��hfEd��J�N]O?Is10�h=\����x�;�'.�zM��8�
/TWBs��Q���ñOs`�n���?S�¨@�έ̋-s����;f�y2uw��Tm�+Ԉqh�_�ޟ1���%)�y��I*-�{�k<JEy�)���x﷏�����#��;
3�M�:ɋ���2��(�9Jz��2�$z(D�	�W��� ����T�~^eM�)ϫ9�T�/I���쫖����4�7��l�YK��?(~i���*��!v�lP�W��k�qj�6.����[=��&V
�/�<�n+�94�5|��{W�^>FW\� O�6ѯ=�.^p�/m}�����hnS���S��Xiٰo���/Y��~�Z�<ј�Ϭ�&�=�8��E���S.[%�ǨN�;(��н�:�M��uܴ���v���{�MF��_��"y��q��n�,>Ý�n��^7�fn�U��͊��jFÃ��%��n�k	J�)A��ӯ�\�u�4�t>�rm׽5�5{3de�p��8�^`{�{z�jֻ��dCO�����ާ���b=�H���>�C��bN��(Z/h�^�;ss���y��)㨇��'�b\!	N��/Aw�x�'"í8:24)�칧�:-V�|6�*{��+ydQ~��UMl=��5��H����h�����e����Y�����E���b#����ӪtT`I�'�*/�@�rt4�S\��p��ǳ�^�V{d\�>�y��w�W<�DE��5�q��=�m�=�}�P8�H@X�(.������x���������w�gb�,��`޻;U��q�#<���`��%���o!�J��y����M�eѯEY��V�-0�}�<l'}2�����J��t�x�p"�"o<��QI:Qra`��7E�������n{��@��[�=N�g���Ԟ���~�a�q���wi�'{o��]묎�yֵ�8�{�&(V�t�8b4Ngvq~�v�_`7]��Jz�?����Z �n��`)�s6b�*��NVDY��eW;��]��2�s��{o8��:�2P�>�Ej��N�Xn�����{�ײSom>D��P�T�DH������Lz�>��ѐ���E�[n�ɝ�(-0���w��oU컧�Lo���?�j�'֚tō���珂���M k�{���|�TфC\y,ۘ���T���^���w�b����'�~6k�ܾ���9Ҽ�5��W�Q�Fl����b[H����:�~�#MW@X���?��Kr���!L���ڥ�%q��^� t֡_]�3��txN|Q짤U�������!V9dWOq=�h�ɵ=���]g�ޘ*#0���\K�lg�����Oy��{i��n�Y��rWcʑ��t��o�9���c�M���V��=����m����׈B��"� �y�q0&'bg~s �<S�	�L�����y�\�?+���k�����Z���g'������}��F�/8��K�z�������s�'�����S�ZE_4瞻1p�eY��0}7`�)A]8E�ĳR�q���9b�s��4�)>UD�@��z�4�l;���A�u�uLNZ��<�ʉ �טz*+M�rf?�.�K�5�q�Hp�+}�5\w�i_53Ϳ�
�o������4k�oL��tG�,��V�6���1|坕�C 6�#sV��,�}�N�y���y���)ι�OxzG�?� ����p�Ǝ�}_yM*)�H�d� u��2�S_�6��oJ� .d4/���g����߭�RI�ðC�v&����JNI�Z�ab�,�L���F1N�w�.z7�6:��«��J*�Bw2~Ӥ(�P���C����Vt��'�E���T��|9�9<���^N�d�t�|'1EH_���
[�U�^�
.��Q���!)Ȍ]D��?E� a�𑣔�'��y@���ǅJϖEA�|�D�
��{�,��YY.g���j�I܆B�E���(z뽒]�9�����Ў����&cgV]�r/�E�\�p�g^ԛ��Q�1fwe�>1o��;�!;q�T�1��{��+���[�p��j����w��]�t���N�����W'W���g���F���.#D_B�C�;���FF������it%�
0b�Vo��gOnצ��
_��7:
7��8���2����b
P��QXqɮIVU>D� h���k�n�u�vr���}G��oQ=R�<�|��6+�I�vE��U��
��u�j�xX��x�B}�Ċd6ЯN����[
��r��>�t^�!Vw+�X��K=�"�ι�Z���\��}����a��ĳK�j�J`��CG8iɸ.P���F,"Q:��''Y��8z�p�»�\n~�ﾠ�{+vZGOd���@�u_M^5�f��'�������컮8}��3�8%ܩ=���������T{�j�0ζ�F �<�=3����ɛ�Cn}Jhz��b�]���]�>��L��f���0�xt��w��U杬���XasW�i+ �Ԩ��41�u��o��/e���ȋRz_�U��lת�'͋*�u�9뇇66�%kS�§c<�fחWP9ɺ�ܚ(V�b�6}Rh��ɤ�͹P3�R�����;�Q�m]�>�hN'�Hk�n]x��^w�=:h1����p�J<a�>�J�W�Z��,��^K.�����{w��%o/$7�P��U��"����b-�.������.�g��x�%�H��O�ba5W6Z����(+��7�T<�e�H��_tw��l,U
�]P��}̻��p�qՉ*:�A)����c�;;oà�*��P���w|��4qB�r5�s\�	IPz'�&{T��{N4��7<��b�wOs`�n󄍇~��rS�`��D�3�v�w��鎋�]+��t:������Ť�I��f֊�UIZ䶓�;G��sBT�7	Ú%x��f��+�9N������+��MTFr�s����|d����U�.��iwqYΓ �@�X'WXR|q��;��qP�}٩٬Fu �UQ�����r�M-c>����)��a�J��*�O���m��͗%�K��R�\�H���yڲ�G�����)W�C�����C�M��?���r$�d�E���"���6��[ұ�Y�b QB%�.���2=У�k,����������Ν�~5z.��7{����IZRͩ�����a$/�s���O�C�Lv��*�1͞���c�q�9*D�����K�=�'&I���!<�aG�UP��9њ�ᚼ�ٛ�#բuΊ��k�n��C ;�T���`���~��IOo���
p�yS�b٠�o�ޚ����͂2�i�!DwG�2�d�$#�W�Tش�����c�*z{ov�g���$�<w7S⟙'L��q+�:�g�m���oD<Ց<P�\`2/cu˯z���'!+%�]��wB��n��~��s������4�֊|V'����!�@z���3���ܷ�������!c�i��ܯU��N�,����A_-i�W�砉�\9v�Y�3p��d�5�C�F!rk�<�*�7�.�E���T9���gH�/n*���p�y���W-�J����OC[R��8�WWLy46���9:�j&���GV�ۉK�G���ˉ��ٛ� ]=*l%я���p�1y��Nj[ѹ��Y�ڭ?{��{�%��}2Z4Θ��Mr����wz���6А��d�H@b�s�e޶o;޵�3&���0x�����W�e1*���gj��hh�i|�J�䭿!G��d���H$ �v-͊U�w�p�r.)0����w�+%�ɨ�1+�_�k_r�<Of�e���U&�3t݌�
��:[��@��[�)�l��+K�]�2C�v�I�7�q�TXp>*�$B���JίZ����y}��x����-7���ǥ�."b$���5�Npr�	����P�A8.�Ӧ,謪�}˥����Q�X;�"U$�r&g��j��"�AC�eX/á�Mw��H�B[~6B���;�����&�����W�+mK�0Kૹ�*u}g�'I�JF����U�罭`�~y2��mtͷ�>~dF��
��V,���:�h���`Vo�L@]��f�m�N���ܰ�0��)��!ְ��]�<M�2TY��w���LLN�bM����?�����[��#�ݡ��Vk���Z�5#�càlG)?'�d�'�$�*,�J�d�����B����6ý��R��M&3������AN"��CO�?!��wg̟�a�a'��ά��Gw�n?ͬ�.F�)�_\�?6��j��%�Ǥg�5��8�-��L���3eЬk"[�s�x����ۓ���Z�v�i��游�}��O5h(8l�j��-��'���MG�E��@��M�@i�He]��Z՘��4鱹L=�h��+ �ɽ+�#��B�Ú�r�pқ��S�ǨI�N�<
=ͷ`���i����wf<��ں�'^-��V�is��VF�e:��xo�2�;l�{���R�60��3�c ^ќgf$v�3�w* ���,�9L���ԧ-f��d�2R�itM�o@�ehp��Y�I*�d�#U���5H�T���[�j����:uj
Ҙ�z���[��W ���3�;7�ևet�j��X�B������D��
.�.*؈q<a,'�d���f`�R�jgV��K��]�<���O.�ϕ���t*�̍j[�ӳ� վ]N�]���q�����H���})Ϯ-�ۻ�@����L"��ܫ�ޜH|����zV0r�Dn���7-#Ih1��r�f���[J��ʉ%����#e�Hp���ۧ�&��6]7�u��3�ܱ(���՛K�ݺ!�yFܴ�X߆A0e�����-���݄�zk�u�b��C�(V@\�{r����h��v��Sn���͊��Ɨ.+a�#���H���ݹ�Rˑ����"1A:�1[�]ft㔑���!��^��]'�E����]I�{dpC��Y�  -	.�*)� �j��;�N��a�:Z��xm��AGD�,��������9I��PL�˩��1�\�&������e��bN�5�T;���5�D���Cu��^�ޥ�Ә��gPn�RM�t�RM�]xխG6���
������t1���L�*gP��F��Ƹ�.EoU �)�̏��;��Օ=�G8��5��eʅ�Y,�l��{��2$i��ǩ�����(f�6.$�
�4�4����'`�Y
���c�.�"�)��r1a�ܶre�`�V�e��в��(�&P���rLV�$�V�F[�X:L2���΋�5ZZ��Jb箎�]��QZ,�������*�Ms��ø��B�"���k�ɫ�3ΖQFD+�|�����v
�[��mb1����
35a����g.�K�&�r;k(˖A�A#}!�9+e�ӏ;/;$2�d��+��x=�r�%��}i*�Ӭ��!ͱ�v�����{��t%��#���u<��\/�ֱ�"���N�\�Z�U&a�]:dfʇbM�f��F��*��$x�2��W�,����*��gue�	�B���nBs!�t̅餁��ҍ*ݴy�=���F��[�U��d�r
j|s�^�L{�WN�TZ5��"�44�����(h���DI󳴕��<��c�x=\�,Bc-c���Ց ���q��'��$UB�J�m���gs�S���f3��|`lV���SԵ�6(*E��QQ�+�̳0*�)��cZ���.61Vڢ�EĪ��UjY�TEEU�r�ʌ��-�12�$ps
"�V(�EAF#[J��m�±,&2�*�J1PD*V(��b#F+�c����IU�*,T��,`��b�Z�"��QL�cb5��-�PU��Qc2�e��cU�X��9�dA�*(�V[\��)ff*ZV,F�mm���-AF�Tb���q���Z��rܥZP�A�.Z+�¡mj\s
�H�R��Q��[(����[l�֍��b�q1��2�J��L�mQ���[Qc")��V�D��" *
��ܲ�TF.9��4��Q�Y�fR�([�U��*+��Z �Q���PĬ�(�J㊢T��kJ�V���f`ңj�#�U�G-1��j�f%�[kC-eK�nc����n\�`��\6��QLnYS2���*������+-�2�8� �Dih�UUQX��E.f~������5����RB�LE�Յ�+��r�>�B���ǙL�mʸnl��{�V�&�d�oe��9��2�[�+���<ka���G����2�L���t=� �R����Wi�'�{�����B������Y<�4���1��Wl��wz���7�'� ����'wa�B�����Ăͳ�y�ۛ��=3W���ߏ{�����~aQH/~�m���?!����#凬1i����z�a�˦�������E&:x��b~C�M�rOCvi��+6É�����2T��M*��=c�>�k��_=���?��o�|��=I�x����p�)
��u3���Af�����x��TR~�I�Y�i>O�w��~�V.�M0��P��(c7�&$Ĩ��;�'�ݤ�
�l/)�>�y� ��C�3Ȥe��.<xL���14��Qg�ys&�^2u<���@�?!ܧ����7�B����C�R~N& ~9�4ϒ|�M%G���2c��Z/�T��&����~� |�8�ѕ�ڞ{��{_>G� c�"�>d�R
z��a4���1������Շ��3H%H}i�*Ɉ
)�|~�ω�
����&ӌ���C��>a_̚�4�'5�i�2W�~����_�����{�}������t�"O� ��Ձ��|�Vg�M$c?y���*,�\M3�1>C�1��<��E:w@�T8�=�M�Ld��~�i�Wǈ�~���ϴ���۽�����{��y��<f�5�d;���=aY�h�Q� ���氩*�N!S�ydRi�q��̆�HV�>��u�LH/����8�C�*,�|�4�0���S���x�yd������q7�~��؞,�>1��  `L|>u��v�����`iaS9a�f�u
���բ��8¦$R��TY�������w
�@�6���Ԟ����xû��u1%/�7߸�sͽ��D}��xm=����Dz�{��x���;�S��q�s�!R(x{���a�<���Sh%f���t���S�L}a�1Im��;�'��H*C7�Z�d�
)�f���\>̾���:��/�qP: x#S \��;@���a^�~�5�,�%v���C�(��;��?+*��]�?e��
�o�,:�H,ǈ����E'졉Y��'�8�_��c�ɿ�a����ׯ����qz�X����2����U���Ө?�<���}��\�'Vͽ9����i]�]І�R5&iޭ
��oT��3[�g��G��V+��9�Wtfw\*b�Q���ms�r�;�E6]���aY�� �����5��+�83� ~�2| bT4o�&������ي(|��x���D�+:��}���6ì+<OZ��m ��6^��%UI�]�掠m'�ӌ�7��!X*���k��D�.��t��ĵ��<>f�;5Lf�~LC�T_5`bV��o�q$Y?y��6�a�w���N�Y��LG��§Y��r$�+��w&�E��u�������2�;����%W�$x����(��y�%M��
����z��B���{�O���i��ğ�I���4�ALd�o���*A��?}�x�0�l1�C��ҳ��ܕj��:⻍��F�|�� _��]]Ԯ�mN��^Y�&�a��T%d�߲:�*��0���N VoV~CI���v�L1��+�'�����Ag����'uE ��~�6$Ⲥ��4�������4��;|�w�fH�5>
"=����q�����i��TP��4�g�14��	�d� ���6k�QeaP=J�=��S���QC�J�����O�Vu��o�!Xz�c�S�R��?&ME���YzJU���G����9���%UI���i? T�g\~�p:�|�*N�<gS���Ğ��g�=LCHWa�٤��0�bo�S�4�P��,�q�2kW�i� �����ӻ
�z�f��jx�ZR\E��;�~�I���Xg(�q����a��d��}�6���;�&��I�����O�y@��0��>�M'�� V|�CF�"�S�-�������5������[�}�"��!X��I�;�'�t�&�6��|��M (�h7f'I_�|�� �ϙ9�|w�:�h����svu��y�kB�2~q=@��懜�{���.�@���I���_o�߻&�|¸��<��>a��4�Or�Au2�@Г�ʆ�#�!ܰ�塌�&0<k4Ρ��
�~�1�0�����6�|��s�m�G���������~�]}����&W�����+��&3��CH��%q���CĜB�x�}�+�W�TXz���e��*�O3�O�*Lf�w+0��+�gL:Φ!�i1�0�be���)M���}�����.�m���D���>*��T׽���K��=��2
���P����G0�a�������s��Ʊ'�Hc�am�H�����y�2]f�N�AmL}iT��a�&!�dm�8:�" �|YWy+7��38WGU$'�#ʍ�����  ���:L�x��}��xt��`�H<���ClY�u�0�wY:�I�
�v�㙓i�a�k�q
͚��?Qd�>�y m+�M����2T��d�M�+:k�=~���߻�='��Z�������}������U#�&���x�Yԝq��
�S�����.!Y;�3��0�h|s3hJ��S}��Ă�9a���q��r}�<#'�=�����I*�>����Ǿ������1���d�9��̞�H>�z��N:w�a'�=f�������{a�O�'�%V����1��}�u���;���T2�e����}��+8�3�N�k)�q�&r��i ����CH��*��8iRW��L�>�i$���5ܒ��
γz��?a
��w��6��9H/߳ǽ0:=鈀9h�P��9k��܋�ߺ(m4�RgO2.�q����Vz���u1=�Xq1{��AM�Y�u:�$=?}��+m8��y����B�ϩ���x�Xm���&� T} M��qj�!z���e"~���E�N3�9��6��WL<ްQg*��Ʋz��@��Xm۲~e�$��r����u6�Y��{t�hT��z�:��
�y��P�Q����1<��OG=���{~�1*���oS�IR6_�J�E%qw�m ��0�߰|��
��W�`{l�%f�d�����<����!S�'��v��4¾�}�y�x���DW}Z|���,��D�:���{�d�w�4��D�*o�ͤ�9��;������0��rg��f��i ���4��C���E�aXj[?%C�J�:��t�B ��=�Lq��>�\/�/�Q�@��!Y�,��0�a���p6�q�<>�i��T�%W��!�6�@�w�m�;a�����{�l<gɌ4ͽ��Ag�11=/�)*AM3G�,���*=�/�U��ptá_�^�ꢗ��}�ş'� ~J��+;<��I���~k!��h����Xm��N8������^����6�>d�6w�<d���d���~Cܲi�t�(a��U )?)��Q͘�+��Kt'�n'I��A*�dP8���j���a[�]���9���&�2x�nT�ub��b3�z�S�83!����F���i�X�E����aMl�-�l̈́��,Ֆ��m�\�i����j����Y���1䎆tk�J8�8,<]�������8ɏ�~��}��)�� ������J�CFf2u��<�?P6��e�u@�*��L⤨
l���AN"��Ou��*Aݜg7C�,?0� ��<ϔ{���f\��w����߿s�}��ɴSl��i;��M��1�,]yHV���鬛�4�SY1�'r����I���2i �H^�T+8É���3l�Ρ}>�� \{��f��|����p�r߷����tS�����7Xx�=aY�Xq4��+����� (�P�c] bO�W��,��p�Cz���6È�&!Y�%N���Rq
��L6@��ё���\���O�qe���[����_�%a�x����ʦ�6���w�h:�E ������~N!�?Nk!����1>g�� q*M!]�Q�ɤTXT��$��0��,�5���TJ���^������_V���ȖIϽ�#�=�>�!2z��a�=̚I��'���e��a��o�p>J�H,�<�p:���TY<�̊|����<9���&3|����8���Sꤨ�o��~�a�J�I�҇m���`DLw��q��~s$�aRs�x�H}l�O��6���d��Ý�I8�N'�܇�B��7��6���T�����J�ɬ��s0>@�����9�[����2�_DD{ xC�{�>���
Ϙq<��Y�qf�̆�H)Y�d6���1Ͻ�_�:�f�W\�|�C��o��Ԟ (��l�p6��$�<�ܬ������g��똊�ߋ��ڑD�*<{#��EH�{�%Laܪ�O������8��n��gɌ7���m ��^a�>B�������Y�u:�3���咱g��ɾ�x��T�O���s�y�s���w��t�<ݓ_�CL4�j��v��P�auE��E�0��r鬕q����Q2u18�7I���ɠ��Mr��<`�0�'S
|{̩>v�Ĩ�������쮏[ʸτr��f��`d{��tm �@�39����u+/l4�g����{��H)QB�:�$�E��X|¡�i1!��}��&M��N T�B��>ۿ0�y��`��a������WQc�u����*�a�]�n�ՙ�7s�wW��&�����7��;��Ao&E��Px����u-UƷ`�_=w�CI�B�6M�,g0�������q�W�f`�5�8��j�l�	�jq�^�T�������սݹu�������!�<х{Ś��8�#�`31�1��Z�q�~.�����'r�s��8�D���f�l=��{�ʅf�xw�H,�4�l�uE �uQa����=���|:<*G� �_|	�f�~�?w���y�{� bT8����=d�4�	�o1&��d�8��;�9�aXVc���h�d��:s�6���:�혓Lی4���n�a�i1��0YSI�G}��~��;�~�}��翽�݊T8�E�SL=f!�z�:`_,��7�|�H%I����l�����4�l*w�O��������d:�²k�牷�J�6�����_Y11<���˞���������w^�<��1�`y�S��9��e!Xm6��'��Ć�'�=q'�Qg����2u�<�� ��y�i�{a������m1�T��=���)8�}�x����5�羙��F�%.䳜t�c�۟�	��'���[4��0�@QJ�G�»L@�=Cܥd�;�=՞���'���~���z�]�o��B�S��RqYR�y哻��Y�y��^��3˳;�:���k����P<"<�����&��ͳ�<O�z�!�s�a�E�{���=J�0�r��& (��RW b���u�yܓ�vi��+6É��7�>d��_{����*����z�]\RTǜDDd06=�����q����)
�l�g]�8Φ�6w_���=B��������i=O�� �d�]n�m��?%Cg�P�o�LI�Sa�;�=��u�];���&��|QԵ/��1X_)��d�;a�
���M<d���y�d���N����@�?!ܧ����7�B���P�T�����c>I�4���D4�2c��-���9�t:��긳�S]��?�1߬1oCwHJΪJ�ՓH)�h7�M<a���,���N�È}n m*C�O�y�&�S����>'*N?���N2z�i�c�����z܋�X���~�͚�߫��Zԗ���%q�c�)8�FQ~VT��֬nÊ�frÉ���g�;��q�E��}�4�gb|��c���_�:�O>�,4�Ĩq���<J�z�_������x�調�+3`*k�*]V�!�}xqF�,��%*�{K��rs��U�( y�̓JU�<�����Řp�`��>v1�)�w����Q�X�mK�	��΍�{���e���.�����j�̓�"��˥T+f�
�i#6N�v�U����x{�]���$��Ld8 T��>Cl��Y̅���+1NUR8ɮk
����>ve�I�u���C\�+f����:��_/�<a��!Qf�d��Y�u7���ὐ�-���ZM� xA�z`}����0��|�̇�m��d�?r�"�L*g,>�d�N�Xb���Y>q�Tީ��J�8�5a��M�*q���kRz��B�����?]m�C��ŭ�{�t
�ｵ���q'�|7�H)�'\|9�?���<'���<a�V��)��ҳJ���6���SG
)1���7�L�~d�8��H*B���ދ�5�{����G�0 ��5�z�q���eCI�'��;��u�z���׾\ ����nk����S�;�x���3���a�B��0Xu6�Y��QCL��E&�߷���2�~��]��QE��&<� c��H6Ì14y�>aP1*��&��Y1�ϳP�%v��o	�Vu�y�s��u�g�浓��AgXn^��%UI�]�掠m'�ӌ���+�'�)������G�� Tx���:j�Ͱ�1P��j�Ĭ?3�o�u�Y6y��6�a�v~�6��V~�����L*w�;���+'�;�|���:��Ͼ�������l?�|�<> 8����M�\C�>�Si�
����Y=e�!]���n���c?�c?$�ě?~�H��Mo���*A��~�$�<a��br����gU��<OX���^}��w�}�*��n&�I]�������Mj��㐨Jɣ�duf2T>����N V~���O̝s��a��W�M��sG���W���;�)4��>�{���ǹWaF��<�#��|��T�%g�����LH+�4�!�x¢��}�i6�Xbi�w�<H?�1��TYXTR���Rc�u�oVb(~I]�a�nͤ��gY/������;����矽������+;��>Gt��Y��O�UT�O>���'����p:�|�*��:�a���$}�Y����
m�3��S�4�P�2ŋ4�a���{��7��Y��~g˺��9�,��u��yw^�mc�vX�ҶmFԼ��7����4͝u9l塍�l0�1j�V2r��l�R�������na��8QR�&޹|��b/C/����������Uj�rӺ�G��0u&���\";n+1tA��0�(W_�=�<E?�����sϽ�6���V}�Z�(��?�����O��<?o!��d�>g��a��d��{��M�(�O�!��=@�<9ߴ���/(��a���I��c���+>I�!��N���9��{����>���E ��勦���Z�@�c}a���& i+8�~�&�Y57f'I_�|�� �ϙ9�w�q��<Jó��svu��}�݈���� z�޳w[�&�^_|��~�߼�=CI�M9���&�u�q��yM�|�z����QH.�_�qYPݤ}�;�|�1�a����3l��0���� ����=��@�6|>����O>��4;;�\qaH���1�0 P>�2�0=1�zc?sY"����x}̇�8�f0��V0�����uH,�,��IURxg04� T�͆w+0��+�gL:Φ!�����}�3�c����Z�}3�y�����>f�x�������a���g�|��$����6Ş'Xc;��M���f�C�3&�XV�_���Vb,/�Y8��a�J���Z�g*��^��c�:��G��e]F�y/�����p ���>���>e�'�����;��&�v� ��:��s2�E ����;`��d�l��6��\��fm�P1*l�U& (��Xb~E%xÎy����?x�|�x_Rg�޸��=�,�0�%g�Y>՝d�6}�M"�d���K�T�!S�N���;�6��_�#��
���J���:�̪WP��ahim�'��ۖ1�V�j��L�������*\f���n�D�*2�Ё��j,.5�^5�W"n.<�!ZU}�+��)���c���o�^�CRG(�t'����$f�(��֤қ}v8<|��3��8���U�a��;v:�3|�<L}�x<��-�1�V|�zr��&�w��)[}���X��N[�2�\��jt��h��(�j�[��IrU���j^O8�8XY��$.���O�7�"����@��am5&��!�*�ja�ښj�w2+YL=����u��z���,�\���Y���U��� <<!�����S�w�^I�����0;M
t;G���8a42�j���qe���[�kӯU��y\��}řU��7�AS0n��a4/�p6�8|M�`&��U¬X�������)%��W�z㿝�t_�,s�KzV)�y����9њ�3W��ِDzV��gG��ϟ��ۆ똭�j���T����p����'`ųAl�>��o�*"V� ����'�3Ά���^�8�殕ܴ���� 0-w]'0nq��oސ>�����/�s�����f��/欉�l�B��r��U�'���U���%��oݬ+ȵZpt6�����;��ر�����5��!��e�wZ����s뒑�r5�3d�!c'�<�L❍�|�B�}���֙�n+������hC|xk)�<�鉃�\���X������p6�``r�X����(n�_8RV �|�n΍��N@�H�r�
�V��<5�+���88f	jf�]���7N2�D�Fj��3HTCϝ���M�k�c�\X<i��)�O�y=F,q��[6RN�e�2�+n���v�3��>5*h�vȳN�l��tӐ���]_gRT�BzMNMqnx2ǔZ׬{���tt�������F�WŦI��߇�=�xiE�o��I����V�.�S��*�P�|��W�L.գϾ��k���z\�H�S�j��7d�g���0�.+Pcl�P��Vf[�{
���Ζ罎���f�]�9s�^h�3��iEkճ�χ�u��g*,UAP��2D/���)�^��E�u���Y/����!bJԷ�U�"�C\cis�q�����s���<�]V�?�5ca�� ��rWv�-��:I�g�mi��v���Ѯ^��P]���,6���.���q焇Ci�z��D�)�U��s�o����i���#�
��2�W�{��'5o8��&���};ʸ���B$[�
�������c!ũ�ڸnto!�.&���D��UCӖ�H�I�s/�E��m,�h�*R3��­�۞��(E�ח���A�g�nB.
f5�՞�;o3ǅ+����^�������X�KNV���[�*�su�Oh����g5+�Ҍ�X�y:W�.�>���B����C�k��G�|��"�Ϸ1v�Jmno"|;�}K�V3��J|IͰXV�{�X �`P+�+�x;l��� b�4��h�z�����%o�{����*=]�w,� ������y�+��<����A�8���N�Xt2量����uy-��tV� {�xwN���SC���tvW�^�j1�ŧB�iΊ�yL+o���h�7*j��nG��v��h�aGsj.l�1�ۧgMy<�F�׊�dN��*d��������}��9&�l�&���a�Wz�b���I��N�����W���Ⅾ�t�^3Bl�`��*��<��+#���oJ��c�b��aW8D�m�G'�㐼X�����G�w7}��HwG�ڬGՍu�����G?C��⪗.�~���-�#0ܗ�雒;�k*��<7�%��ڶ���(��ʸ���|��%7���P���DqUs���VMR���V'=����C������z��:�X�@O�Em�qP7[�����yv{�t{��./LW9z��z�B��L�7cDX����TAP��|��rϻ�sd&.x�v#��\L^�s�3��rɇ�wɿ	>K�W�������k��w/�I��<�\�o,V,#�4mWs��?����J��+�W�S�Q�8���ڋu�]�Ǩ�X��[]|(�a$��eԾ����ս���(�aj`�r��h��M;r;v��U\/1��j2yPe�yv��s�x!4�g%�1�vw[�x%�\�$o�,�J7�4ґ��Z�eJۼkNY#&�;d'��:���rM��A3��)Yg_�U��b�JWSܥu�T-����.��]�hO��pmG(;�vsjnY9ͭŠ`�(����1gK�-�	PSP��Hz��x�M�;�q�03��#�++&[��Nf�͵!0�{�(�u�w�dW3h�=���A?�g�	�,Xԭa>�க&P|N^����R[X5�y4V%�Y;���Y��&��\��6*D��I{%�LGr�Fj}�,��Y�P'��Ee�y��X6�f�M+%k]��
�Zޙ�Y�H�}��Ed*pnݥ�l���PQ�y��v_KQ�u&��iG���ŗ���.��k/�8rw9������-=g!����Ob_m n��9rn�:��X[D�i#��΀�У��s0�}2&�ήP��S�m�cWaOZC8�$�ݻn������n�a���!�w�cbb;]5�ͣh�t��%��n
/{� 8P��Nr�Y	�X�q�dv)�M�E�ݲ���ĳ�,�m���a������K����K�]Q���]����>�.������[XoP�	M`U���Vt���Kw�C���3���w�@��bBk�����ңF�խ�ڴ���W(��Ա|��U��vN=F��l=���f4����������l;���],�P:�fg;�CZ�
�V����ƹ�31���6<��(�Ή�8�pl�����O3�h�]��K�7�c����
���ut7k�mԮu��ջ�.X���f�Y�5�b���7Eoj������ڶ4�ۓ�r�J�7!*\���]��Br��滨��v��=�f�l	�b�6��C��8͇�QeB�c�T� K����3�d}]���eK�簽�^%�v��������I�,��#t���-����M���PԄ}"��l�lʖ �Me�<�f�Hr̻)�Y��D�X	:�Ü�]�����>��hr47��;f�;  v�Vs�|����u����L�G>a0`}�j<�Ca���j������&V���۝[ZX\�|{S�Wph�E��:��B�r��&s����y�����Et��ܕ}�Y�å�b9Zć^6[���B���T�vY͹_VW";�8~,�Y9�Ǩs;Z	jvP�8��o�Wu��LS�x�޷Wͮg�����nNP)cRS`�P�e
�˩�5j��!:Խ8��%P���R�v	�,�Վ�W\�+�:���7s@�!͝�Jx��z�1���.����{%��b�U%]����nZ�)�̢�J���`1r��D�[J�-1�
ŭ�$E"�Q�̕cV-�����Ш�R�����*ilH�"�ED�EE����Fڢ ��Qh*�)b�QD�Zܴ�TP���TĪ�A�QQZђ�Lh������b+�Qq�-h�K����\ˀ�lj\���f�ţb�A-���1F�E����Ѷ���,���T1m�5�,\��.X���%TTƢ��d�1X�8Z� �Eƣ�s2䫈��ZՊ�`c����h�B���""1PU��`��P����ъ[b�������Y��Z���-�ES-X�������R��G��̵�����+QT�*J��R6�r�(�H���b�e�V�-Z�V���d�`�E���F��ԩZ��*�VԪZ-�VҮZ��6�J���`���i���ҥj��RեB�X��R�h6��h�K\L*�U��E�ʊc�����媌ڊ1U̹iZ�`���y���<��t�H`�Qcѕ�!Y��f���͗�R�U��fc���;:80��6���.)%V$#G��ܞ蹥��  <��ZE�Z�����$Tdb}:�q�OC��_�S7�ݯ���\):���3v�N�����.I�wヂ��-�>���LJW��H��,�0�#�]��kEenؒC5����┪��D1��\;�j�������<�M��<��FŪ�A�{Z�5�Wt�a�Qў�b�wS�$z�1�n�&���1�P��d�uEW��:_H��-�_g�-w$|T�R��.�QV��ͺAIү!�܏�S�};g����^�-��C�f����QEF̿p�ey
(RT�W�z�P�plز�|۽��ո;���[3���6IZu���뜆vjU��P���͜_5l@h��+�'"������wo�0MiWo.ƭL�������Ak`0�v�\�uCbx�Q6'�cM����Aq�8O^v'�л��ѥإ)�)�Plk�2t-Ύ}V_X��/�Ψh���3��i��te�e�]�)��P��x�4w�J�����OG��8&�sME8�c��V��ھ�Z��w#7���Au�g>9���F)#�)k�Y�M�x��Z��LR�J���oK'"�-RehU�5Z��왼��w��]�!{�L�aWN�&k���E�|,���|�m�
�v��5}6"�2i�{��y��ʞ5�e����|�%u������bՉV�#�B�����0\�{�8=��4/d^*P$D��^�i���o�6I%��>R*P���u��!F���AFV
paߩ�l#����1�\��E"q`�cc#�8B�Pl��^�O����}��^�)��xM�D�u�"�c�/�gwn_�0Ftx�wH�w�
S_xR�#�Y�L�`{z��ex��`;3Yi�����%a�<{��[���#S��ƁN���N��8A`��=��OQ������Mr*7b��V,���*��AEBt��s�'�?4�|RCC�zk�{��@=D�g�E:�﫻�+1�ƛ�Gu����q�m�E���/�sJsޕd����N��R�r߽���KP�c�
�6N���6f*���|��1F�-��CMv�-V�˫�Y�
�x1i"��h��|^��]�}J����z!
6Ճܴ�ާ�@f��*N�(э��'a�깤�jထ��a�%z+��A�|��OƢ6+�B�\`2*�#�l��6��W�^���"�B^����h.��M(�B�����]w��|��1�v��ka1ӂ�w\ѳZ(������	����vv��'Fno1#�S*���U��6aJ�ٷ��95��xGZ�����b�2p����'��U*oE숬�?x ��{�M�MGJ�Ϲ߭c���:llw�VB�k�"�~�k�������B��X��λ�M{��*X�W��s/fxb�<	�[�3�t*�Kv�`�5�:���f�c������eGF�LX�@���`�RvTD[��b��6�``A�<����Kv�5�%E)��XOJ�:�L�L�~��F�`�)���{�xp��2rȗ�&w6n��ʞ�y{�%�4в,��!�@�<*�9�R�Ez��ӎE��lýǞ0��0��󩳅�<����0ٳٷ�W�]ˊ���lچ4�.�+A�H���]���ԡ���˜�=`�]�EwDc{Vw�r�������B��UFH�P��y�4�k��&�8򘗝����uiFJR0� r��t��㍗w�07^�
!Ȝ�f.���w�㊓7O1���� u�P�j0�6�9TŹ�'A@�hXx!����X����/�=j���J3�N��ZjX����Ux٠E���Uz�˵W��挜���C�ɦ<(����IĜܞ��uM��M����^p۶bnK�WX��}�՜Ż��N�u�smk�cӎWww��b�����׫�ݤ%��(�Q����W7OEV%M9�|HNVL��,�D��)�Ҡy+��f��wop@�]/.�;�\�{��U�WԚ��w��nn#M~�X���'�X�d?b���ԋ�p��F��N&0�w"N\�꿳�w�_ge���ߺfҊʖD�;rG1Q�*0�o���)@C {�L������@��%�X)�s;�{-�	׹�x21�|�NV��c�mu�=f��s��9܍ "u��:)s�����囪�V(����X�|�vԭJF�:W��{v�Oo^ɪ;TP�1�ƫ�,�qnXiпZs�ku�4]x�6.�#��/a���ds�ִ�zf��뾋����p�'��F�v��:kT���P4� �j���s�
�i���OQXf\P�Z��0}Ԟ���9�Qg����}�ӎ���B�Z$rF_d�f\��ff���?���T��}�Em��F��줴ś���U!���O�w�*$.-5.v��PҘ�1d��A�QB�_r���Y�-t7ow�7���Ū�&�<
/��L��f��5P�SÕq\��p0��M�����{��][[�ƅ��\+W�v.r���T]5L3�7����˒E��=C���'[���j�ք�{�O$7:�1�.�⚪2!�)�V0��ࣥ�7&�v:[�`��Um�����z�3[5svkI����;�5<�Ք =��+-sr__4���}[
0�X���BS���C�瓭����6�S��Z�+���^�ޙ���ZO$맛�O�4H�G���Ti��-���]�\�~=��h����^O��.��ޗ����=au���o��+�x���������:�'|�2���<og\[�����%7\?#�M��^�P��*j�a�W]�}�*'B��V�3��U�%z���zL�G;6�b�
���_����@��O^r�J�U��:��k��bǸ5��j�nq�8R�����!�K�+XR�U��D144C�Q�|��.�vp��M�f��g�xWn�I��aZ�U��"/�kT���jF6�`c��=Ҭ��@`YG<JU��;᮹��-��_�b����s�'��;��*��_����:��[�� A�騰��L�۝0כS1vnnIbw��ɼp�[��ӳ6�'AW��a�~x�gF&VP��?x��G�&uy'�� f��\�fmP_y�Bȶ����te��0��V��۽�i�%g"Hqk�4��>ڞ|0Ny>��w,u��]�gp�{�a�V� G�I�}Y�Zdqt��wN^m�V�R��XƜ��s��vɳ,��Et�:�/4����#IHV�C)d����!� i�5pO�`��X�R�J�as��r�eݷ6��&Z�"���xx��岒�ޅ27'c���R�\*���_El@h��<T�-W(F��W��R��t��d��KŌxxq�����W�6,��P��zt����z�Q��
z3�����gq"Q㐠�Vo��.��Rw�#�v1�:w���|\gT(j�bݶ�zH1_BqF�
�������x�-�}*�`nqOG��gŷO&��6�c�vBٔ���"�>^`�+.ś�j20L�(����J���;0p&{C�B�E����uPK%ێ��v���Q5P$A����@4qCA��+�U���!�+r�o1,h��[�"�&�Y�t~��	�=S���ָ��@�W���8����bS͋^񗨊|Oy��f�{{��{;;��_�:|�ǇC���G���־��a�U����S|�dn���7��P�If�G�J:S5/���i��h�i�N�h�>?a�C-C��F���-�^���Wt�ol�E�bł�U���8w0����.��>P��m��;���:Fʾ#���mv%�	0Q8OY�A|�}2W1����)�㒯�U�I�Y/�̉N�Z�y��o51���xp�����Q����Bn!$8i�7Ȭ�2�hfLPqG�2���0
����L7���w("���V;r�� �%HU_�����央^�-D~U0n%���Mv%�~Uf9�f���ͺ�>}�:3[�3W1�
<�vۻ���3P�p0��ޤl�,1g������Emuʘ)���j{��Hqµm�a�3�)����~�o��s:��X�K܄>]*�i��pB��
SǗ�����MS$�����Xw��C���I��*G/�f�:�<�'�T�ו7��;�3�f���KUV��W�y�a9t��l�E�E
f��)��P&(x�t��#�KR����a�P�f)K��Xǁ<q�tΩ�T`I��D���s9��4_ft.^l����ҏ���	��RL���7�f,������39ynm�g��-��rD-+C�0�@��DRJ���1v�1t���bL.f[���������k��ZmH�};wb�����v�B�S��Z���~4�}�G�=�(����ܸo;���`}2�	Prj1*��n�M�"F�2��U>��1���`�wc!����5�ށ��
1YFƻ7�v�5 �Hޢ��Q�������^��n����:.l�Ы�kΕ�g�q�׍/=q,}#�Xq����v�"�S���;Ƚw��F��(�=a����j�Ov	'��ý��^�,rM��v�=��:P2�ن}]Yk��hNL����UFH��~�R���J��qVʭ�/pѫ��P�1�4L�Pj�j�r�,��wC���@j�& ���!�O�><߮\˩�4����![ZY��}\|5��F�r��(->�\�X��\]9�^;�5.�S��'8���?`��~�����#H��x�U�}��%�T;�2����G[S3�5c1�\[��h������b�@��W�r�J����\C�L�.��yVNB�����]�����7Y�k�	~�/�H��ig�G0�S�g��@�˶��o����&OL���_aF
���`��X"����2�"�t���4�P�qqX��fˠvo���ؾ�}��d�� D�n�D�ob�\ꞼX>�=�:u�Wџ/���]M�%�ǀ)zDw_�|����W�QΧbg�7�^9z	��bӠ�M�n����ߌ	���2�xH�Y]հy:�ȖP��{E�#Hn�������W�鞜/����> ��q=���7P�!����L���	^��/�:�Dv��Ԡm��==����/��`�-�W��{b "(9L9L{�I�E�x�w�Bcb���tv���ش͚�Z'����G3y��b\2�}+^2�7ʣ�q�t����`�۳Z:��묕y������ԟJ�ɒ�{&�|U9�i���}N���Q[��*�������!^f�h�*%��Sx�>X��=��xuV�:m��zU���>�A��E���[eq�a�ʞ�<��{��z�C�)��s�2/]�.]mK:&O���;h>M�
�jC|����N��Wr�C���
S}.�x=2��7mz�T�*�s#T4XḒ'=����4w{�����&]��3����HJr0[��q:�<ͩ�jw�C �`f��+1���T�ܤ�)/O\�E�s�j�{5��yˮuq���CK��y� q�<�Y97�]�]�Q9�4�l.��m_]P<��[�Z~1H�ɇ�u;q��9ܮ��;5[e�nz�#8�������=�A�ł�|�����:P��/	���K��Q�4Vl��71L�C��|��_o��`�i���f�ݟ�p�8�؜�Q:ɦٜ�,��9�N�Q�����^���D�hh��چ�v�"^;{z�~�s��{k�#��=�U+�Ε�����o])�ՠ���G�0�FLGOw���kh���:ȭ;�9$�7�T�W��r�ݒt(�=-Չ���������X�u;}4�v�R�q&��K�ca��?��ꯪ�(T�RzJ30~zptg�����E��k�>� ;Q���:�OK�'
���]�6�Ϊ��=s{B��^p���wP���б���q�z�-�j�6���1�5�L�<w�Z�sy���H���fvL[�]����f0m�
N��!�<��k:,�Mò�"_tt�oIX{wcJ��\p�T����,mw/Z��O�I'͋*�!p��VFT3T��ަ��%{x�0�م2N�x�f�o��c�����V���R�����ߗ���+��G-N@jE9�Xǉ�p�ݨ�:9�eg�z����6����kmq]��x�D�|bX����nt��-HH׆dn�9�;ئ��A�w1e�ų�9�u����MB�Tz��j�v����*�?�78�xߵ���N�lY�GF�ŭ^�ƒY��f�oJn��>| �����U�.7ŷF
}��j�{UVj�ޗ*�7�h�H���5#�㼱��h=T�P��1���+�C�GéR�-к'�nY��߭�;`v���	�G�S!9t���	v��_׆����с +6���S���Gm)��4�3�A�������UL��O7M���VQz�ċ���e�s���f���E��}��KY�ABl��3�35;��d���ԣ]��1��	H��
���ˊ�#���`�9���c�ʳ�nv���y;�h�uh�tha��E��[B�uE���7��ɞ�ƽ�C�&��ݚN����7����ܓP|-S��Зz�jp�޻,9�u���+�ؐfͻӘA�)���]i�5��)1�*S.�
�{^��*�U�lժڔb���I@
c���,%��w`���+�ݰ����|ĥ�n����ӹ���	��P�&�MBU�����:���:�æGZ����jK�c�)�����{V�Xo��VN��>4~��U��al��S~kd8 �t���/GS�&��;�Iޤj��Fr��O{���5�����s��!iG.�,���olƍ�s����W.O�=a�~����?�v�t���v��q�W�A���6��yn�	��B�.�H�dmag���/(*���4�>NX[�ZN��!JB�^�QSm�4�B�e�Z�X	ї({2�c
��e[���y�}}�N�y��7K��h�B���Rn�w2V �k��P�7�u��acm��{�ee;�{4��0�8�t�[��fq�VC�P��}�8Yi�w8"']*}���awN��o�ݴ�ur缳�V~Z��I`��!Rs��Ê$�r�������B�&vr��:����eZat�6��S��]�ݽ�r��L�n��5�W�Zj𙕍���Ĩ�u��e��r��*V��8�>��d�F`Ӈ�9�n��Ֆ��cn^�t�� Y)s���Z�X��M4!�۱%m�)SM����@�����/��U=ww7qм��&Fl�����w>�w`�H��n�8�3r�Z%��+��t�o
;BDq�z;�|a��S��ԛ\:	ؓM-a�gm�.Wj��c�<��J��V��m�n�V�`����e
T�t�"����qKk�J���* c�xT�=�R³58ˑ,���%w�R}]D��E����`�J>��|*����WHmZ8��m�n������(�.���D|�YJ�/�W�զ5#�s�g���bkz��1����լ�v\W�TtC��m�t2çAo:��s.���Q!Ks�qI��xB���J�Rud V�sn]��caW�CDv!y:���U����Q�\�&3{ۗ�X�<�.�%�WRT�V�Ғ�[ڂ�w�=�X�BzJ����!��*�hE�k��"�|ݬ�;�� �2�]J��K:�:u�nz��J�hT���]�U�D�q�-�˝��^���/HBQ	�7P�v���Jݒ]彂��|H$J��$S0-�B���kS8ڔAѶѢ��b�0���r�5����[)K+EF"��U��������q1��(*�,m���V�����%�Q\s+h[[D�V����Ԣ�Z�j9h���9VUh�A"�TD̹-3��j�Wq��J�j-T���\�32��2*��f%ZR��4J��qƋkJ*�Q�5*%��Zֲ�
�X"Ķ�+mAJ%�E�V�*V)q��R�R�U�R�s&dj�Q�Q�m�+\jZf*娊�(�D-
�b�ejԪ�(6�.9�JZ�iV�eX�ʍh�����VZ6Q�h�ʆS0�8�m�$EK�-���PX��\�J�R�1�T�e��rԹpLR��ڬr�T*Ը�l��m�\̦	�i\�9QbZ2�9�U�*��Uq�q�cZ*R���9�0���ra�[�m��R��B��eDX�,��U��)Qe���FU�ɖʶ��m-YUJ�������e���ʶ��f%m�^R�X#�;hc���i�>F+���Z���L�.��$])P�9s%^�;#]�i�X{0�6�ͺ�td�����{��*N���4OF��w6:��^���q��8*�H��X#
���ůx�$����Ȳ�T�e{{R�Sn[qJ0�~�%��q���T���ߩ��1�WVe�<�m��̯]fΓ$��w�������I���N�7~N؏X��K1B��#�3w��7e��R��y��Iq��m�]d+޷�8�_*� ���7BT��B�� n���Tz�×�*^B6���KZ�$��ҫ�bǺ|��I�b_��s��:�
�����>�{0$�g'�J���7T��������+�mY=�x����2����\ �u�;���#v�ɧg[S��#&���#;��|+ӎec0&G�K܄>]!ܴ��8�����uAm�ufqPH����YŇz3͛��4C��VG_TZ�b���ʝ��y'��(5�R��CJ���2Ar�r�UjYu�i�NE�Zptkj�R�3����\�X"��i��|4G@�A����i�k�]��\(����S�
"%K|Ōx��:gT��x��$��H�\=&�6{�E6���ӓ6{�[��^�L�n��\���{�\�Qx,��Zoђ��]�M��n+j����r�ۆ�bZ3���1S).f@�;�$,�Ջ|��ҙ�d5�3��n��eh���B���J��1���d��SvH��7����u.�g�%
�~�њ}>i����!�<����ǰ�v�k��47������-N�We��Λ����51�P�|i�������J�ڂm��������!�T(B��ɴ�ܖgwf`����%..� �>"@����|����Ƚ��p�M.���A�Iy��D�L[�����ubS�q�&}#���W�1#jB�ufn������56�ħ�N2���f����snT�-ᇂ��ϰ7w����PT*�$B���L�3������|�1[�Q����\9Qr�n���gqƉwz#�@�QD��&w�3�L8�=�9���U��]$B���C���ډڏ�dh�)�Bhc���V�t�d3f9{=�&�\�ȫ���|ߍ��}X�Uw��Z�,In��i$ӄpjӷܖ<S�_3�'I�4[]�K�-'�ܙ��J�8�����V��<9�
�G����G ������7~関n�^�!��"�Y�3��
�p̵�?'~�P���j�v;�)�m�QcJ
��Z�}�M���	۬W^qrfN��I�uqA��4.:k%�$�:V��彛ib���#J:%(])�6�Zd�A��ѕ�1�W/�}��yX⇕�ZT�]7�\��/3�#���e@���ܱ9���������*s8�<�v?7(E����U��R,�\b�1V��9�F]b||��ww=��؏ΔY�ަu�J�s�7���V�%<�[ǘ�ϼ�^񩆓����C�ٲN��J���˝�l\���5���i�s��W�^�j1Έ��[�9�4�:h�F��fr2T��]���E{`?p�qlM��R*�]��X6U�ڗ��x9�s����]���:�����:�X{�Ծo�2<;��@�#a�-�FM}��W��S�Ҩ�#8{��F	=����X����G'T�\DteAU��k�b���8E'��ֵ>�p����B�k�K\f��J3�C�P�gTHP�z}.v�@PҘ�1���ެ��rp*N��}�����RLͼ�<��.r�Q�|�+��,'����џ_*`���_��<7ӄϼ5'��yz�`*��L8��]
0�x���	NF[��q:�<ͩ���Ev򢈍���de
~�̪��$��r��+���J��+��;p��d�b��v+�M�Cژ8��;]cx0��^��Z�{�&mm�f"���3|�4��[�_R��r�;�X���0X�,䛓E*�����,PP��llE�x]6-� Nf{޽mj$�H{�η@�}b+�f�7�7s�"9�r���t
��T�x�r�l�b����'ka���7`�w�0 *	A@��	W�����{�i�C��:"��E��V���p�	"IZ�髩O��k��76�dyPj�a�W]�1Q2.��鱻���ck2�����a�\x�w<'y��T��A�Я����}�Ɲ��:.w���J^GB[�͢����U��NaS��b{���s�*�J}�)Wm"+@�æ��%ݹ�i�p��M΢X�g}�j�z�_Rz},7L�B��U���`�wu����P�O޷�6�L �<<�B�s{���������q���c��Mc�juǦ�myѝ����5I�j�"�g��+\'[ ��*��㷼��y_�:�,"�Go<F�K�d7�{L�үS��8u*�{C�-���32���P۷�W��}�kGvp��1Vbj;BͦZ���ո�T�F������B��P�l���l@h��R�v/k�/�EʡoJ�k��F[�R`gH�'9�<�Q�K��Z�#1#��祉?M��R��FP��H�pq}��[��9�4�/ݵ
>�Ve�� �؏01ep�o3Mf�Q���Y�����X͇��v)���)N�h�QX���gD(^q�hR�Q����ˑ�^c��ݠ��+�ϲ4]�V���7�������r�n{i>GTz:TO�L1~�vܗ8���xfA�݌s�ӽ�z��@��E��r^O��a�(�rbDX�L]\�
=V]��k���~�z��S��z�	�rr��pf�볹���,�U\�fmD���|�D%�b����w�U�C�yW�էr�Hv�0Ɲ��ǛQ�����+�=� hN|��-�A��h=T�P��=AE��+����\ƶ��v��s9��TM���߬䎬!�Z��ZS��w&S���.i>'�Ԟ�4���,x�Fm`#S����aN�P�ܸs�V�΋k�"}�|���7v��	� ��V��������w�\���Sf�<��;b=bX���X��F(�$�2\�*#o2Vq�-ީee�FޛQQ`۱�����UL,7bT�^�˰{�i4�ٻ�l�_���v�=�x>E���Z�c}>o���=-Ş�BIU���wPCf4�j�,�[�=z�va�ª�j�x6d��Z��N�})U����q/x�C����f����n��o0�XE�uu�'�s�I,_ve�o�0dYE�|�7q!x�Y.��R^���L���d�V���OH��us'xWtJ�T{�R��)���.�lt��qR�B�X'<�8��-ֽΝ6#Z4�H/���ΈW+��y�o�#�]�lSX��ò�5�U�CG���K�Ꝺ�nL��n��⹤��g���ťV������Xw��Cc��Xĝ�XU�W��F'�!=��z����akIh���Hg�}�����6�JH�r��߭�v��M���1KC9�����fV�
��k�0�添Y,yr~����xhq���$.>�����q��+�qX��a�`"����ycIoD���^�:dຸB�Y��؇�NS~��ڄ��}��'����fo3X�I"��AQ ����]	��2�iX�^(��`���3J��_r�����
|)+>��.u�������#'�F v��ʃ���k"{FƻU9!f�'�D����ѵ
���-0�&xzJ��w>*�@i���P��̸لִۜ&��U��zoQJ8��Q�k�:S��:P2�ن}N�gͷ��TX�PT*�d�N�řr�ט��%}y��l�LQ���>��Ǽ�r�y�� �vN
gq��]ވ����ͣ�~I60ɣ��KX��/�"�|��fZ�=XX��/BWE<�ίkKv��Z��:�[.Ҋ�
#�:�q�g�4�����k�)�c-ɯ{".�ʹA�D�*WZN!�w�J���^��9v���Ut��OQ-�9�O�؟lvI���=�\�s��Z��'��l��г�U�>�|w�D�G����B.Zq�9��;q�v5��$J�L	��5[��r���B%F��_h�ux��]�/��k�.S܊Ȩ�+6����d��_A��*W���o�T�u,�P��*�Nv%P�|kg�s3y�ѓ�q�GPqA�~l�B������r������Bݥ�-�AS�A�FT�0��>~=ˈ���Ī���9KA����ZϢ���e�E?������0�jE�3�zyA돻/z)$NJ&��E߰߶��@����!l�~��8|�ϥ���i:��b��b��2�6M�%�<�Qs�i��R�:-��j����9��.�zk���+ڸs�b7zH���"��Ms7��Vt|�g��,��ԭ6�,��p�Y�e�k��p"|�:91߯"w��{����P#H�þ[�t`5�_*4L�siҜ.�	[�䫵��x��x�=p?�\�C9�k�GM��ҫ��~�F.pJ���?3�ʲ�<�����r
�w;2!�:H��~��Q՘�m��5�+���t��{����w2^1�*u/��h'(f���LZdw�&7A����<۶!�ɥ�qE�$��R9�X'Gx�{�<��:�&^{
+�����#��ξ3�SWA寽���X�΢^��@�Y����Z�xo����ME���������H�<�ؙ#F�Ǔ���oN[I�Ӊ�B�th��.FF���K��e�L�}��h��=�*�i��Uܻ�.1WS�V�-#�6T1Br��aE��PN;NX�	NFt9�'[s�ʐ�L�d�y�2��n��X���V7h��BZ���X�\z���,Лa��,�n=���nW���h�2��9�A�@�M��T&<�Eվ�)���"�w?9;��֥Yh�@NXX�CeC�|�p��zs��@��=�A�ńx4m:��;ٚu>�ZՋ����٨MOu����#/���NpZ�B4F׸/���'R���מ/zg�}�g���\���\�a�zj̓�ݧ$o!�\~���"�o"&�M���V_�^��(Z>NGs6��\�k���|+�<���^�ù�C��vGbv�.�n��fWD��5S=Z.���J��R6-Ul<�q�vб��n<�ǯ��Oρ�{}�ѵ�U�۩'���x*��]�Q�g�6�W�^XW��Z[�䢡f��d����m�Da$e>
V����y��$W�7�{"��J��̎PL��"�F���x��KDg(���K�a�����e"v��"��M
��7��A9�]W*������-�2�.�pvP�i���uEV����>���T��[]\wy1�Wg��i;[{r-Q�x-q�_'���G�����f�[%S��[J�!V��e=Lt���7JfɌ�1��iq�K%��ضkBn��L�C<�͒��`v�*�%����
؂$d�TL����ֵ zm�M9�n\"��B����	�(�$:��=��Q8$���y��1k�r�e�I�[�M ����,xU ��}�ܯy�.�@Y�k�2t-�t�b��ژ����a+2n�˝r{���\P6"����}V]�?�ڌX�~�z��ܨ���Y����Y]g$ޛ&�إ'�qF�|�B������%���qW��G���`e�A-A�����k��"��ѕ��4��w�y`hↃA�r����!*�o���e��!��^�p�a�V
pa߽Os`�W�A�q��)D�A�>l��^�R1w���g�����z���e(�ck�s�j`[������fR㋪�5�ӫ����C���lʞ���}$�c�S��/o��ks��W��#�g3�W0L���{A�ޱ} � _�Jtt��:U�㜅�v3E�u^̥�2LO���pw��;+���J�fβ�!��lv�>��c�L���MC{A��ٲ�t�De,���U�qX���m#+z3�uk�W�y�7��Q��nY��b�'lG�C�5�b��#�v�l�<�Y�央Υ��X�5�zU5�������9�^�=��8W��U��+)0jb�V�ܭ�ZerH�Y4����Y"��Pq@X��F��'(/��~}��Q�o,-��]�]�.�$������'���NP�%t�ţb�EV<��D���x�рz,<��������[?�hv�-W����t~KE!v ��4Ϛ�U�=o�<�"���w�6C2��5PBu�aތl��1��2���㕌�c�tM�5U��z崗#x���S���~�BS�Un^�~���NE�ZpthmY�[��zNgT�Z���h�t?(���~�]��f��i���:hz���E������?W-3�^$LC�8�:���;��%mt	�W�F�5�A���`��(��1y	�gMb��TD[�W�:�a�{�S[����t�YD6А��`k����^iX�^(�.�.@�Xj:o1u|��4T��k�{ZRC�MY�,vl97���xj��Dn�n���/'{tt*]��m<<�GYJ!�hAʹEl���Rz���$m�����)"�� ���a���Z�O{�Zh\�2w-mZ�ڛ�t7X	���|]M�oy�1Z+SUW��,U�������l��F O3���r�)�Ѫ��X�Ӭ%�%uY}u3�����Ny53:e���/7#l��ɼ�CN�78�*l�ET3%v}ī(뒍-�
�;��t��Ŷ8R�����hR���ezޥ^h޷�VU�Y&I���/����3)�x�ᳫq��(u�}����BI��]df�v��u�ien�k��a�>O�m����X����&��K��V7(m'9�k��z�@��F**�v���4�@;�9j�nmJ-��,0dξ�j��+�c�tޓ215d,dǫQ�ľH-%���'�AsD�����r�K��̷}�H�3�4P����9��0�Fi�� q�Gf��+���7��+�rR��lB�^��w�hB
#C���G�������C̎�#��%�\����p��7�	�'lA���pvھw3��2�!�`�
j��:�݀��:��-�y�q�-�0������WH1���_a���GAL�t��@7+N�Ul��-
�8��h��p��G��u�MUcu=�<�+73M�A��f���j��ULᦧf}1$`�%�6&Ǩ��E��pYg�VQ��nB͕��Anc!
�,��.��9�(%Ԩ�e+Sz�H6�F���ɡm�"o*�i��"�I)��wtw1P��4��A'6�Ұ�����'�v^��I-X�'�c�1Iն;���B��s.�&�p��dt�].�݊ǆ�J��#�PV�As5�܈-l�����)m��|�/WN ��Ұ^���v���)1 ��i�\ބ�@���ξ���(����qh�;S�.뎸�k	�Xl�Ѻ+S<*�4�##E���m���8P�t���ޝʺy�n��Te�t.�xN:
�æg2k�hm�)�.�J�n2�㫣�]�n�|���k�)�)�YY��:�m�]X]�pT�dc�3���b]�R{Qֆ{�g ��������t���Sh�-[m�s���x�Y4�mf�}2�#xrn$�+{:(�ٺ����d�4s����Z;���f넥[β��,%X�r�m���\��a�׎�R�GU���-�c.	0m��� ������Y!��J��*5Xv�G^��!�Gz��V�Z6��a����	�e3�!���t��㶬\�{�V����t;��8�,�V��>����z�n$eՁڕ[Uo�%��}�tX�ݼG}�h�ٔ'^j�'!�EI�t���f?�wF��8�]q�;�¶6���ݕ����
�s����k�h�g�6_F�?��}<�fEU�5�J��Ҭ+�*4҈���j�DQKʣ֨(�%�B�Q�*�������b,Q��U��Z"�h�e���X��[B�`�#mE(ʫZe�����Kl��eb�U31r�aV��r�
���ŴJe�أZ���R�kYP[i,m�Z��k,ETZؖ�)Z���5Q���j0�T��j���k�0��FE��m*����Ʊ*�2�Ĭ�[�J[lm��h��̦ �B�2Ֆڵ��QV�UEkmR�+�0q��-���eXVRڪ3E1�1�R�mJ�EҨ����QQ�m,X�X��h�j"#)V(��˔��ۖ\��""�X֬m��W������Q�R���ڶ�TE�i-��J��.e�J�E���%-bV���Ɣ����FҡZ��KeJV��C�V�(�1,E�6���̙"�b�m�kq�kZSm���6�le�I$	%IfMB�u��Шަ��
j�3��6����R|�Zy��Z(h���5`���ں�x�N�*��U7���'&B���r�r���N53�vv��R3�H0)zDp;O
�\�8�$�OWM�kθj��K\MR�z�L��ѳ�c�	�L���3�0��� 4�ٵ�}���Xo4u�Q�����3�=�*d�_��n{(X-ᇔ�|�VT�梂���t����:��o%s%%��
��.���iFd:.F{���T\�N�gW���R����clc夻��{�����P� ���æ,�����Y���@��Vr!���*�QM�%{�TCG&���͡������%.��دB�o�ЉQ�g�|�c������r.z�`5��س�X|����V�i=�\:O�R4�}�KP<!����Ҳ�^��j%갩��������qFaT��j�)���0��������3a����B���/�sh�LN��'~�c���Z�Öt=U����P�A��9\i�'e�!?s�*�F;�A�g<�{�0iO�\�~�[�]���N��� m�׈B�R)��������^ȫ>+}C�)������muvom�nkU�h,���>V>ln�&�̎���DU��:wNf���!h���(J�F-����*���Ħ_9\��v��]뗭+�9׻�8hM�w���B.�nM*��g����K�w/�x$+,�Յ��1��_���L�/��T���ka린>�e։����<}{��9�zkH���{���J��y�:�+n������=���F���7���Y籀mӀ�'ɋ(c5�\w6�/�+�Ș�k����qD�#�b_a�;�3G锞��B�ݦ{�vI[of�{�ݬ�~SY �{��=f�%�v�^�����#zT쿗����>�m��t��8ˎ-�%�%���v�I��U�F{x8fs��z}��Ƹ�d��1�oa�#��1�oH�{b�I��Q/�>�T`j��ބ�(.zeA�ojsڨ]�E0yɖ2��j���	3���M��dE��Ko�k�5@������.�	NFt9�y:�
��Ǌ���(��Y�a-�Q)]Kl�E
T�O)���K!}V���=��/9u�:�����u�o0�!#q���uZƑᱬ
;�~(X5��� �
�zCHڹ�yh�y{\w��M���9y�O�(���IH�,�:����GQ��ht��^���x��h�Q}�-�-rF�yc)��v��<=ǒ�����
�"'p7�{dȂ��";�4�pߕ�ۍ$����-�T\�z}��z�,r�Z򰬲�_NV�X�'��%Pq��wW�Ŭ��mî�P��5�Ů��;-�m�Ѩw7W�k����3a����g��I�íYJ-`�|8R��B�>�>�i)���5����W�=H�ܠc���	)>��)�s�lnצ��p*��7:Q��!���o�)[y�D���+��g��^��}s�%�H�F՚��)���Fm��Xݰ�_�,kvԌmV��B��sP�?7��(3yN���X�0e�j��ݏ;��U��Y+1�}5�Ǳk��-զ�j}[�q{8��w�I!$_�@�x��Y��;C3��Ծq7o�����u�Z|ӂ-�o�g�2�^�U��A��o���	�}t���u-�Є>"��OS0��ڳY:�2���%9�g���Di��bʭ���[��g�|R�R�y�Q7���gݎ��#�)�PWNOs�z��M�0H�y9��\�B�w ���x'T����� V(�V�AB+�n��ےn����,1��?5�J��J���r�Pl�r7c��u��P�e��Y��-��{�z��Ua
Tqb��Rp]\9����j0��f�w�J����(���{u
qd�
z�Q�S�蝇U^:$��+'�����bCήfj0��j7�mt�hYQ�*\c�ІB����2��:R�U�f�����'�avԮ):� a:�S<*䢪���:^�pP$�`�*\�U��k
�+���j(?�!8������F��������E`��{auC�Ns��;U?A"HG���%��.R�tXY�UZ�;r�X�*ЯG@�\��o*4qCM��w(xQ�\�rl�i*�iFP�`ja9.B��8����go���<|~��p���]����%a���Lܳ�6M��-|���e^�)��ۮ�����C���FSN�+לy���&��>}�+���W�G"4�M�I�p|��p�Yȳ��!����@�s�T>�'�`���M鹧>����0�k��v�qqc,����`0[�*c��E\��{d�l����9��^�����i��\�cޟ7��Rs�*���O����$��tAk[��#�n��aΌ�ۚS��J�X�%WJ�Z6)��V<�~W��;o5������֨\ �u�4�t��o�6j/����2�pͺfeK��tO�MC������q�z,e�/M!g��Y�z3͚t�ݬbN��
��~9b��|�g��~�Z�%AVP̽\�﬎�`��՚ճٌ-2���E�4A�܉f�
�"�ȭ���;Z���Gm��Ŕ��&�A��$���Z�0$�r�Jf�xN�%PǦ�7�tp5�1�LY���m|f�L�o�d�뽚N����_y1���b��r��߭㰜��8:46��+�M�6WWyo�7KS�ǽ1R�
�z�>�>GG��k��Q���B�鞧Sҧ���PBo�(��:��8�f9x�.����G|5��W�}N��$9�\5�=��;��+Yn��,ُ޲�>W��XhŅ����vBQ ̡���A"]%C�ކ�4�����e(Z�꒖��E�j���LR����`��m�ﻟ4<"C�!��¨W#�b|�x��S�G�y!�I&���L������o�����zQ��PuS����@ 4�[�Uu�~���o�Bb�]թ�D�������nmʁuN��r9����;�糯h/c�V.��&ɰk+��_���(S:�޷�=����E�T�+�}��h�՗X��U�2M��7c�xM�P���ޛ����ʅ���>�ڏ�5�Wa;�ڪ|�#^o]��w��谁����}����|�Z��٣ܾb�������~����XHz��Hem!�(i��(z��X]�Z�\��\pǔ����n�O�bG�x�����P�9������)�a$j��}���j��uǙ	H<��,!R�Χ�W8Χ�L�[�X'�����l������u5�)�n)�G���%�U�є'W�{ǝy?��5Cx�.��t
��d�:.v�ڗZ'�ǌSh�j7�(�#vj
�
7�ƇN&(>�E9����_�(����!���>�����"��3�%Α=��ۂgWG�Wr�`�������S����	�_:�|iDz�g*�����fܓ#������Y5_��n���⮡V����1H���zӵ��&ZۣPyC��I�H8-��#>_X+��v�ˬ
xjxZ���/�d�9�_ۯ��ڪ���f5ӄ	��m��g�ЪoB�~WYb����E�t�!��ׂ[\+op���"Ulo3��Q�٬s��C�n3�:]�b7���z�4�A_-�N��k��)Y��*��o�I�)�����鯴�?`��_zg��7-tH��oNwҷ�񫥴`�K��d�[��ˣ��'ȩ�Q6&�فgjԜ��Z�ab���:�B�i���}X�4�S�bե���WV7ͤ� ����Q�iD�����Y��S���]tʌ��{S��J[�u���Vߑ��}��nWCXv�mg%v�Le����P�g��^�AΒ��_q4�4W��U�Tne�;�IxJ����10��T�ܸOEWy�Mĉ��+ x���զ���o�������]E6���\�vJ{H\�Nt���y[x���M�yƃ��Z�P:���}������m/aB��#fu��xF}{����.����.��i���ҢƘ�r�MG�3wQ��7`���M���]���nƈ�T�hFPuB�m\��y?(Q�3��JN��:������e�e��b�Y0�M����@G`<���Nt�
��U�H�XAX����+����]={7�Wu��O���(!���#S��~(8���׋�q�:"�ؖ:i�d�/��0�C��&w��zwg�J��Di�nt�yh����F\�U�Tj�D���G&j��ս['�s{4�GW�b#k���^��c�U���w�ݠ�w�ֹc|ݹ�;0�J6���0�.����xH�|A8^��4,���.��:�[��a~.��q�K��KK\BG��)m+Q�c�2^�A{C&l!�6���a���b��]wV����H�����,f��W�J8Ѽ� �4��������^��p�T���!���B�i�����TF+�B]Zo���K8W/��5w��]?P���3�;�ZУ���L��ef���������
��c��\N)sn�!�9��B)�Ԭ�!2�9�Iuy�Y�0ӻvV�2q��(��Z�08^n��L��m$��iV��[iI�c��5��k�b�S^�B	�]kn�;V�P;=R�R��Q8p��Ê����^j[�8��תg������[�i�p��Q�u������k7�̻��+�>0�`ck�����At(Q���>.���*͍�r	j�nMlW5��Y/�I qp��e��_�Н
N��uAG��]����Q����W�?t���\MpWv������Rc�ƣ�bۧ�OB�q1o��!-�o��FF3С���ǹH3�5��$��Bɷ*%7��)��׍���	���弑8�D-T,\�;퇌������6C�=��`Xg,�4�P���go���=k�����@�ʼ�vD�^3��/$�ojr28�?(-{�^�)�)�O=w�p�\`�w�u�W�x�)�fQ}���k���L1`U��:�3�]���y���*��S��>N؏��x�y.�Cd�$�����B��z���F��O���_��鳥9���{cDp�2V-3o��f�^��ܧ�Rپ�g����<3��Ed�Ye�7w1��4)w�����R�����b6V3m��y�o}�G�h����Ie@F7OGP��t_h|�L����A��wu�%KH5AV�HJ'��$TI=W��\��fٌ�YW^1��/m��M��0VR�����X&���\=���I������J���ۂu;�Z�(�a��q��n�Y����շc&A�>�Z��v�����צNd򷏱qJ�)A�0����u�"�v�=	�1l�[7��zj/W�h�3dj��<z�Y���1��w2!��O\؂d���4�B�0-g���6lt��ht�_��D��s��۳��ΐe"�i�Ց<P��EᎭ������Zptv�4��ʥ�I���۳�<^쯏
f���N���5��@Pc���B��R�1cۊ5h�HY���x�${�<���S�������_/����M,�ꆻǴ��8�HF5�ך�u�W<�DE��D������Bz&5*p��,0�!ұ=P;6Iqh����l�ZM�0���������<%��7�vv��f��"}>B?�v�^����B3�B����6�(ע�'g��hهz1��;镂\��į(N7N%�gzT,�����^U��N-/$��)�[41�fpR:Ǒ���%�J��{��5�^�yz�Ò�Us���Fp|����;��F�U���z����Zu�L%�0��aL�Cj	:�U�W�5-��k�-�XFm�éGLޔ�V>�v7Cm�s:=.9#�7=[�������ԟZ)���x���QG���!�uYS�V���3O�m�Ȝ��՘.�\���͡�}R�	(yo�J��R\�N����}*��Ô�s���$�~�w�x.��}#���<�b�4 mU����珂���J� k��k��;�yA>J�6%\���Y�6���Z;>=�`�}�Ц�w�b��v���v.�!
������m��3Hʹ��%�]����=�yד��H�T7�b���I�w)73�X/#�{z�{rq��z�2Y�~ݫ�䮫����فx�t͆����1k�#E3�n>�P{76@�^��b����T��9J���>�S!�e�E��%��h̬��y���Cd\��U&,WWc�=`c�m� m�B�)��(�r%ޢY���-�h���NxD=�:�
�����qPv�ˮ��]hs��>��<|,Su�^\�lt�}���$w�	�M�9�7��t��~0(5g�hU�=��fg֞��.�ի��C�[J��2F2C�t�tH���S�gA�M�;SVΜEn:�,x��v\�(��o{�:�o�#����L%���]@b̜v�����{1�����p����eܹO(A��ف���ƆI����J̥۬aZE��:�uuL��v�:�gs)��H�f1)��)`ٽ�$|}���=�\0V��+(S��w;��@�:u��BM��k6���=��a�g6�vh�i �g7Ge����]��6��2�Ko4>��T/h�q��d�wxzFm��1Qu�)f����ոMwX���̓�����( i�N�>�x���9{�P�t6�u�G�\KC����(�4��z�nK~>�����s�'q
�a����WJ!V��6������d�EY;(Y���d�ᛄbD�;�o��-�&��fr��\9���n�W���W³
���P���.Zّ?�%�N�T�o���9�[	�!6.�k%7W�wW��&Q�\��{LQ�7p\�P�RL�ّ�L�N�"5Y��3���
}�WX�'��"��QT��6oG�A��goA���W\�6��{����ʺ�i�v�v� w'=ٱ9��6$]�ӕ���:�T0�Z�Ӣ��hX��|5
�n�g�wk���3w2U!���i5���m��vt�n;,bSv��"*�h��)Nn]����E5���z���Ǉb/c)V�g��2�Qc���qU�k�)ӗF:'���a�e�,dGtuV�x{�FS�1�N�u�]uӖ�#Ns�2EE����[���Ȱ�B�0�/l����g���c�J��Һ),
d����ٓ����k�bh��N��!������/%��cKr��ָ��Q�ӊ��n��3}C/Ek�>��6��>䷣���vqC��������\��;Ar�l���52Y��5�#����E�gK����]��`�I�;�
��r�q�:d�G���#��>��<[�γc4�0�+��Ʊ�rI6���Mc���Eu2!=����� 	]�C7�AF��F�%�X�B�Ƽw�k�,�S4��'�S3ԕ0hu�b�����uЭKw���u=<��'����i]B_��7����=�.�
t�a�qs��e%��]�S3��v�8M�˵8��Ι�em�Z�D��[)i���:MUmH����x�'bur��I��P�ʵ �4N����ԁ��_v�v�w"U �^�����ˠ�stc�����r9��&�,1j��Q��"/{���a����,�/K��uX;���1]�`T�D�)	�y�\��_R52"~�γ$;{�5B�`AJ��س�n��kX^	,|�J��/��I;�.�&&�q��̛������6ԉc,OR�r�TH-?�r���Ŏ�Y3ru@�7M
ʻ���6z�Q�-�}�j�5��H{؃��p��ѵ�|�j�]b-�J�n7�G�ږ%nZcX(�`҅��Q+DZ4XQ
։s0�+J��KL2�����*���l���eEdKV��Ym�Ŕn\2�QE(#R����2�[-Z�fd��R�hT-(墉���Z4T.S2�ڍj�\J�[h�JC�Q2�ELe��a�cS-mm���!Th*�m�ֶ�Yr�E\+mk*X��e*b�DQJ�kh��DeV�bS+h��[jۙpjֈ�*W32��\��+E�.f3-�eE�YD�8�X�Q�X�����ܵ�)kܴ*b`����[�2	Z(���[�XP�(ֵm����R��9-�c1*���cX���2��re\m�EU�lh��6�Z�R���70�,DQ\��"�����ʫ�`	�P!� �IOأ������Y$��9pl�-� ���➪�^=*(�."m�3f���D`�ݙaѦ/WWp]и��Iά<�x�n�7��yMy�5·��dN��:�������@�#�o�р��^!�Q��<�$u#�jh��)����cP�65�Q9�k�GM��#zUا*��i�>56_
=ɥ�)��؋���+p/�]E�V2;�=�39Ć�|��+��V9p#�RE7�<��:�kRQ�,w�:tO�� �a�
���܇�7��b�О��TE�s��aN^v��m"�WMt�(��qŨ�a�k\a�5`�7oӼr�0'�|������i=GvA�eV�x9fmNjw�B��|�*h�9�)��p�@�(V���5K3�IV;Kqm%��q��C�\1iv�۟wP�k����A�H��6o�����%����e����<�op��a���A�b�Y0�N�n3Rî�#@t��^�|U@���_d�d�d�w��V��*,#�1:ޠ��1\���q_������5Bu@x���п��_���0�U�Ϸ������[-�ѮS�;�~ݯMv
�9����yC�r��r�n^H�1�j��r�!��(�����y.Q�V�j��'7[	�t!�HF�e	�)>g�:�&� �wIc���,�p�:4�ښPkt���^�Тcsy��r��a����c)���e�
E�K�׎m��ve��)i>h����H�6�o�D<��4�\o�n�u�vr����ջA�Ƶ��
�PZ�۵q�s�$e���r�t"�Y�+�Q���ڽ�<��R6-e�ñ�n:3m��gv�yO=W�a�}�A����2ۣt�{5`:}���c�P��Y�D�q��U���ޛ��
�wk�w�c�.0��v��������tg�+&�:h�:4����J�Z;�z�Q�u����~�R�E�=4f��lר\��ٱeV�۽��v�Ù'c�)Y�L҉/�1�3��,�-�g�E
��UFϫ�h�eaR/�1����u3����J:��Z��>h��.'���c&����n��=*��5�ܯy�.�@Y�2����1������I[ӓ ��{W����늾/�ΨP6%o͈~�햟��,~p�Bڿߴ)Q\�V{p������,�=7�������QN&���N�K.ś�j2)���(tEfUUN�2�ֵ*:�#7�T.o1ق��B�E�T�H��t�_��[��\��5q���^u����q�e��$��ڄ��RR�B�&�<���^#Ed˷��p�8�[�#K��g�[7��OW�i̠($!���
T�w�*[N`��I�G:LQ�ޏ$	��x�B+���1�W1_t37�䎖�t)]j�FP��5�#%˵�zp��G#�%�BS:h[�,��
.�80���n�D�6\lz�
Q7��#1'�%�%$	�uQ���A��uz�F�s�i��jsܢ�aN�G��d��.�D���H��ҫ�����C#�M|��Dx���S;��\&r,�{̊Y��U
�5���#�;�G��"h#{jxA(V	�<�uW����Κ�S���壾��kEg�q�{.�'��v�+){��0�����*���6[�w��Y����zy�O9w6M��s�R�Ű�����q�m�E��s���뺇�����þT�*`�uޝ��G�>���#��ޯ\�3�u�"�nڇ�;��o�^��^y�ٛ#(t��g�Z�II�ԗ^��2������8ʔ h�AY�`ZŇz46:��Қ1_��t�jl��L�0�
����k�[VD�C/��"���r���s�����F��;S�J���Y+v�;�K������gC\m�:x�����ԋ�����4";x0%�u�=�-tv]s�k�.W^!L�K9�>�e�:�@y{�cͮ�l�o
N�2�%|\��p�mi�>[]&㩝r�N�D��"M����ǲ�n����{bv�/l"|����������ϰȵ�o$�yes��f�/��x��Y4�*�!c�[�3�t*�N7�&/��悾[�t`����B�)VwS����+`���E�A\鉾�r�"�ߵ�C|;��G�Bo�&5*p�a`!���t��ö���d웲Ux,��zv�1yj�̦%BBZ��c���V7N2�g����!lE坋څyǵD�u�܂@w[.?�Ցxn;�(��֞�w�Bw�+%�ɨ�J���l��ǌ]F��f;���t`���tti�k�u��T`Y�Ζ�ҁ�����w�>�Ϻ�t��duA��3�4R%�p�n(X��*�$B���W�ίZ��-� �v�Fr��*gT��p.nJ�ii��#�7e���R���s���<�p]i��;���YP���įo�h��K�r��&J�fy��h֯	�B(.����_B�j}�ňrE��o�Γ���O��Ď���VoN�E.EFO�*����;)H���4d���`�y?t�i��Pw��I�</��w�kf3��7@{E�w܅�g�nͯ�/��]��KGB��[��C��q��]�.x�Laλ�c(�\�T����TYݮ)�^��`'W�����U�2�ux������I}׽u�B`���E�8�,gu��9'u��F��Ri\��w:��.���t���(nJTx��*qv��-���a���6�̆R�>5��9�����G��]�Ơ;����Z��"�����yڹ��sI�����<œ�����y�n*�<O����L��'2��`����T�[�����X"��XU}���a8Z��}t��˭y}�2��Z3� ���9�oV�j;VN����"��]i΁��S
���E:Fĭ���F���z��Q8v��(bJ{ZFga�:�:k��<��_zW|U븮7���z�|F��0����c�p#���_U��7!�x9�P��wNyM�KL�@1��yߵ�P���b�	6���)d��Vz�v�2P�k�`��R�"J�:1ځgjԜ���C Ψ��Zj)s��W,w�^]]�N�-z���#�?��1��;h>Ir�\����->|�>���fi�B B��	f+���fV�G^���s ��"_i�����o�9dS�8����F�ゖ�_�*ӊ��k��9�����s�4T�'�"����
����S{���������W[B�^�ꂄiQ�s��C�5RU����7K'�'RNK�9V՜|.NX��l��}����ˈ�)=�By�D������MV$	1O#"I-�`i0���N1�.q��3|2a����Ɏ��������%��&�WEKН�z�B��g<p7cDX�Of�`���(����X�$F�4�'1��R�b�����)��\�c�!;q��K�W����?w�F|����0���r����}���7z֑~ZG��+%C�TN��q���g���F���y�c c��&�˵�jN�o[G�W��f��B�
x�&}jv�L
��B���[1��x�~f�)�\^J0��\���{�g��5K��~��%��#F�jvϳۂ����o�>'�U�7D֫g=�ᴵ�ȗp�I�y�ע�ӛ��q��0e�F�>�ݏ;�ဴ])y�r�Į����Vc����:v�{��i��aA��U	}QU�?.*��	�h�B�x.z��5O=a����Zo�t�v{��p3��<v��+&�:j%�Y��Jχd���Q[�G��F�fVK5
�k�rDw`ٱiV��~�J��62��+Z��?�=k=�����q�gu͕�w��s8�j؀���'}�NL"����x�êx��9����,z5�wn�hs+>��L�	���6i��(M� -��jMuͫ@�㇀[-{�>p�@�z�{|�}��-�bW|hD�[�QT�ݨ�Y2#�tI��RA7�Ix{/��-�&x`�r7�}����/4��΢�q��#��:�8����|�fP*���B����Lc���Q�U��4:w�U)�d];���]��O����U5��3!7Bܐ�%`3~���1~�:#��*tz˥�A����\�.35��Mo���|1ީZ��ܘQ㏬L&�侅�s�>_i�;�T+�a��N��y��/Y���INTg�A���slc� L�xP;"�R�"/�ә��0牆kh��K3-��K�[
L?T�St���T���AFT�0ȧ��u�Α��q��j{b��9Vk�̤P��c(7TqiD���o�Ϲ^�C�r>�؝uAq��!�����鄻ƇnB����IyP�+�~�1E��\���.��T]Bqgu��o>:4#��Z�w�ͬnh_\���~����R�$�Q˱�E�'
�Cm�ɶ���hEQ�q���%!YUÌ�sy�-"�%l�Ucv����nK�;m��x5qL�� �ĲypwW�E��4���&�mf^�*�z-[���"*�(��
���ı�5�{���N�ݑ*��Q�t5�z��!Z^�f��<�r���%)��nܴ��;��u��m��]ѡ��*�ý�]�e`�:�$�a^���x�Tʆ���M��O�>���rC}�).uԉ��]3� �{���K6�nt��\u�1���V�Zw���B�*s]�B����F�c�RI:�i�qH^֊��+i_�O[Ab��歺�U'6�5h��sR�{B]ޫ��l߰ﺱzp��o�01��=N��V�����j�i۝:�'��:�l}�U^�v���t;����d�N.j�<6�r��[Z�'eb�1�Т+�%�Z�����ɳ^�wĞQ�V�L%�A:�Xm�<��+�a���esE/'����O�����si�i�+�L(݃��5��[(������\KEQ�%��;ۍ���V[}6�M��˫�3h��m=8�2��z��oR
H.o�_D1�c�}��Q�6NG��Aͽn���X�8��Z��ŰU�Hm���,L�HcQ����v��!��nG�T�;�Y�+� k�FuӓK^ovM�������Fmqq�z��㛿f���؎X�w>3#=��5(�U�퇮���{�U���HA�"���T��xdۊѫp� :֩�9m�8%���:(9�H����,�f�$ic��L&p&��A�g�������9��ܥ�^zz�ڮ�]����K4�_�Λ4�9[EE;n�׀C���QS@���n�$e���N���-.kO`���5j�X�m�+���f�#Y"iv�>[��ᾷ�y�|aM!F8�++f-�o��!zu�䱵���x�W��Z�,�̷��&�ȡ�#��8ݬ�����7u��Ek�sa�s}}���]U'B��Y�4k�E)r7��ZOئ(a~�;�s�n,ԕ!x�6��M �PON�w��>1@X�!FKz���X��t�;�Ե.�aNբof��6��L�Ν�
='1^�ylnVQ�L�0u��isK8�F�,P�7�*MgJ69v�K�-x����{~^ӷ�?�#�.U�����mʳ�k��ڃ>g�\���n�!��FjZf�fQ-��x���88'�Vmw�l�޴Q����޳ۚ�]̋r��r� � -b�M�z��SV�}}��oMxS�L�s�I��D9��,9�ץss<���,!?8�!�t}��:�����.�5��Z�r�����������y$�T�r�V&)>CB7T�R�]vY��g����<hd��˲-2���c(�{\�J�c�_}�)�k�P;��g=^�v�b�x����Y+��o���Vs���PZ�ܣ�ըGH�p<�綁���@q�}n;����if
eܳ���H�^���Ζua�]�{^YE��d�nƘ�Y��	��i����c�mծ진c��Q"��R���<��e#�O*�/�Ω��zqlN��
�u�ߛxj�e���&�9�.�j�da<�U�+�зj��m���ӱ��V*^�"�7���v_��A*������KU$T��k�؁w�®�B��WŨ(�浐�{=v�w�V���5��Z�Z��Vo_�̎����*�7�ܬ����ȴ1wTR�o%�	[8��{6�7��b�Φ��^��z�ֺ��xN�,�¯޻�b���.�p����k;L�kH(����9o�^�5;�YB��:�p4���G`��#u|�k Ld,�N�g;���NW��m\�>8�Ӏ+��y���xt��s%��p���K�B�;m�̖���|�Z�N��֝9}c�j�5)�p���Vw�z6���Z=}&(�h��#V����¶���	�5��&w]����1����l.PFw@t�چ�;u+#�<r�8���J0/7��n��X���U��َ��C�tLՐ�Q�Go{��kgi9:c 
���r�]���׌���h��RM�&Fvd���`�W׷.���N��W&����ڲC4lw�S켒�����i���uo��w8�9:��i2��$��>3�#Sd���	5cY[��f�؅ƎrJ:x'@�e��zVݣ\܂����ڜWN�;-2���ݹ[W\�+���%���˺7C6W%x��G� ��q\=}���6��dZX}B�pm^>�yՄ���a�7a�}K\&��Az�իI���gkRD	-����_k��׋{�l��\A�S^uq.�2�76���$9�;¼w*��4L�q\�r�u铫�p�z��jƠl+��+;*��ʙ���.N!['f�4���o�/d�76�[,�q�ӆY�mE9m��VJtE	� �
:�.��M�S�{Q�Y�4f,�8���9�88ܹ%�ͭz99h�h���h���]�wmάKWC�{pȻ~�����������d[���G��tī�J�Ԣx*=.ۦFW�y��iV���7�F&0Fn�i͢��nm7�̵{X��y�R�.*ݵ}{J��&b�â�>5�9���s~~?��Ů�-G���굟b�Q�<�l4P�;2��ɮ{,|�=XI~�s4�L1�^j����u��ƐEY�6.�J�.k[:cE��s�_�M'p\�Gv�]��3l�(+����&t�B�XW�R^΢k��)w����:ؙ�B��@�=�w����&[h���	Οv\����*:�q���%Ȍ��b룽��Kv4Jʹm�א����ԑ�5,-"_Fy�]:$��=���bP|�%�^oSDV��J]��k�;�m�]����ؓJ�"*��Ӆ��>Lg.v��έ{�[,�bY�l��ojq�/�X��2T7/{��:���cP�#�.*��ޫ&�"���!JII�K(�7�*�1蝖^�o��T�$�皳i����u�6���:&C�F�sm�Xd�{�G�Z��G�cw��j��6��h[/b������[��WqQz#���� ��3��N��lɳv�C�����O��U�ldz�,�:=�5EKwr?A��Z�)��X���,��m�ڕ������e-�Ԫ�EU�A��S3���2�[KTm��j�֤TV�6�ZR���[ce���(����-����UP�JR�.f5�J��dmKA\�EUA�*���V�fUQ2��33#�C2��YL,�m�TX)Z��1pLı���%̸VQ�(9k-���e��011�DJ�4j�ZZմ*�V����*�D�FYKV��̵Q�V��J���e-��[\�+�kV����0kjZX�%�aU�DDTl�Yi�X�PEB�*�U��U�-jDU���le�2�����R�JTX���h�ʭ-����0L.Rb+�q-Z��j�*�ңR5,Kkm�J�ZZQ,,[R�c.
R�m�Q�&&Em-�*"(��ڌJ�XUV��UV��FV�ikPX��C�r�o��|��4We�|%lo{s�T� �C�U��5wV5���y���DYkJ��$7b�hgn%__RN+����I����Ps�*;ct��m3�ٿ3ks��9�^���q�5���YU4��\���y�ʫ����ct�Gi��Y��L���*���N�uS�d��^Mz@�x=k�����Fe�&wN�s��E
�0�̼���»����G #U	�B��j�J��NĖ}�[�q
��O����6H)A��h)c���8�D�^�x�@���t��;�+%yW
c8���G��j��B��0l6�㜄mYt��[��]�
�*�E�X�G�q6��y�x�&���A����n��R$/ �&��B��ө��<H���c��Y.��f��.���O�����q�Tb���{��̖����lUlr��{�-+�l�{e���Df����x�[m�'.C�1AP5d�5���F.������,������~� �x��R��y���qVl����C�I�.���u�L/�m��n�����Q����c��wfv *Ԫt��+l��n@�t0��v%�evl��{� ^A{8Mo��>��;k)$����_
LF{:Z����T.�.��F�c\{R��giFH���U�Ew��aAň/Zw{�9
~�W��b�ڮ]у7/%����QH>�E54�[�ŀVmnj�>��9Դ���,ʖ���E1~nx&��7:�T�hEW��S��=�l��؋Z�rV��
�ǆ�Xݵ~㭌����v�索�dEE=��%,���#9qh-c�vr<�\�9Ⱥ�.g���R���#��G"r�N�T���N��w]���k<��u9cck��x[�+]��f��E#x+i^OW���U7�̹O9'w�z�ݾ��d�S�{C}����b��	�v'��d��<�g��՗�ĭ6��r=��3c
s��v�N�I�9����}2D�YٽQ��T�%�:�abj[Dt�9�Bݍd�k^'eb�� N�S�����tӳT:f�a�e�E$�Hiڻ�g���wR�Lbg;�/���:��,�z .����0�r`���U�����Ku��o�ꉐ�;4�z&��xMx���S��a���{��7������v�c�
�݅a��WI+BWܒC�1(H<�i�Q���	��sPu����:��Mfaǔ���}�Ka����!_���k��7��9��O�[��Y�U�1C��H��ET�W7�S�T$jW�n;Om�մ��U�6��+2�΢��ی;�W��Ԏ���r�#Z�C��]��+�I)-��U������w����
�W��S�n�$im��:d��52o�)FK����i��j����M�5QM�;�1���q[VWR9���D��b�󜽷W��<TS��W�C^�m�����^.=���8NW6x��-�ݠ&���f:�U������J#w#"���ܞ��*䨩~�"��h�kkf-���v��:��x边����������G~�W�U����*^8OX��x����җ�۹(�LGS�׺���Ԃ�����E���T�":-ҋ�
�R�a܂����I�VV��'�a�f�h|��n���0L�t�ӧ+NЏR�-�ͻ��N�D��G�����_�	��)6m�Zo�]�ne'x�i��q˽h�7�J
����mrt�{��駣B�0R�:�emW>w��Z�Ё�[Ќ֒�i���V�V�ڠ����I��X�J֖��:�ԫ�+����\���
T�'��6��mc�i�s�p��q��l�%7Y��E
��hL��qݠ�kJ69v)g�-qۭܬ��]O5&Jι|� {dhꔅ	B}L��m�x9cXaB��ל�7{��,5�s�^��&( ��S�%(��ò�^���q�l�,�|�l�S���C\�J�8q�~S�]Q�-^F�͸0�{ ;�+��|$o"�	27��g;��07�*^�^5���	�Tv�Vr�yu.%�WpK�i�l��
eؖp�w��'�/���R{���ry��!��ar;���Lu�P�M]�N��F�F�������ݓ�MP������н�8V՚p�!|�ef��	�h�ќf�E�����̬�(���zxo}�q)u�� �Eؒ���T�i��md��.��&h���}�ߚ�w����M�����@�m%���H:nr���VCr�4���l�hv�ǔ�sB���y��9E>��5q�r�Z���ܮ�=%�cǨ����xy���V[��~⟟'z��c�7j/��q�K�'S֖m�eD��*ڽ�b4""��Q��Vm�;��oJ9�a��L�g�U0��~婆�}G/<��ӯt
����2>hS�Ķ0���8���_�����7Su�	��,�׳W�(!{�NV4H�JIEv�rd�h�ѻ�!�����_I����>agLVuO'�޷rv͖{�� zº+J���,��I�ۤ� �Ý�x��܌>1�@z{� �'}DS��ð\�Y}r�ؒ�8���ڎ*���ȫ���M�8�Ol�����%��}]$����[���QA�3�-�\�F��r�k0l6���F68o:�Jո��Ŋ�NV3����&+$�z�p��SXʼɗ|�7g�-��&4'1yH�<0�[P��<�ۚ���Z�Wx9w����MQU�R�6��	���ª�Uo`�����ܫ�b��)k)��o�����JI9�t����ץތ��ӌU�Fy.��U��K����y������m���h^1̙u|�\I6�J�)":�BK�o���3x-� �M��G���r�e_���wN���@S�1�.q�U�)]�+��-,�e��{�5�Nޙg�+q����*�=�,R)T$k�#����n��Z�rv`;s2#��B����; �2O�}oEwޜXPqAzU���
~�^˚��*�ެf	�K��.��'t�:�L�B#��kqM��$b����E��iw�[mr*2xԱ�J�TS��&�o����QS^�#W;�f����%�-�m.(�Tc��u�L�:��ۚ}g{�Ӌӭ�:$�Il-�C*�P��zc5����.t��Ⱥ.g���qO-h�p��������4f�	�+j��B��g{M+���Cp*�-6h�F�Dd�����wny�@�E��o7�}����3-oEmӢ�pfaL��w.m���3�3R��̳���&�v}�	��f�OsG�"�՜��%v[�CD��w��F(0k��P^3��p٫v��3(`�X_Z�nV��'sT�ޑ*�i�A�ELco+i^OU�X���Y��iLVd){�(�x�6��v����5�^(U�����t����N�	��2�����4�{��	�nt��'��bhvБ��2�59V���������S]ܥ�GM�������׀9;+�LP�ZU��Z}Y��%p,:�|��z�GQ����J��7���s��ח^mm���-5���}����]�Vw�\�ɾ��3�H��X�.�q+�c�ɼ*��ۊ~*�jV*�xO��hw��Z�.�=ga��0�[���ͻ���G
IZ�jGe꾼=M�⺞i5S8��%����!e�(�!�j���X��A�CMzwMVC�yb��+a�y_��%X`���j�]Q��Uў��P�Ze��WF���·Ǔ(]m��ܚ��Ӗ^�`]�����ZQy�Q�Sk�/V͈�7l�>*f�*\S�ٓ���He�l� Pd�h�L���)WNX��L��Hod<�͎��b�C��I�[�,a���/�c��Q��2�5�`���5{j�o<XQN�nhc�u�9%�L���꧈涏�alU��5�M��V�Vl���7�������|�=_g]���̈́b��l��jm��[c)�ݤ �u��z�����-u�m.k������Az}v�R����{{�4_j8���]t��A��M�\���i�N�o3�4�o���+'_OV�� ^��������;�TB���Ǖ��v�������|b�]���ج�NT��|��2�o�,��j�cf��6��L��N�G���H���l�=����i���ܣ72V���\���8�VQv����9wػ�2n��BM,A�б�t(n�ވrƖ��T�i�+U�|v:�
8����x�� ��hF�S�J,�޻�4s�6�8�)7_������vO���X������u.��N��O�`�O,3�]곂`Ps�^^o6sK7[�l��OM���g)��7��q`�7XL�0w�ޚ̹ܚ���O@J+8x�p�s���{�I:l�ĺos�����w��X�B����U='�+\�i\�\S�_����;y}e����Գ��Jg��~=��"]S�D���舱�?��2m�kH�6�?(�:v��\]+F�B�zc�-+T˹gu��'�/D���Jt��Y��Ey����P2/Uz��c�g(vp&�妝�J�w]q�L>笤J�,#�6)�8Fa�ۜ��{��(��ww[��?<�2�m�t���m�@�;KO8ʠ4di��U�+�b��ԟ��ߪۋ�f�u�(�S��8/���e��� �Q��VkiX`��F�ش��S)*�n��:���>����M_�Ȯq��`�	ps��O�H���T߀g���>��m2�6���&���1����+~������֐��
t%�X���d��R��rs^�X�B�!���L���bG:���%X�(��"����9�Bs�/�*u&H7m���[·Ї�5Sc7&���^޽x󅊕 l���k-�б�gn-��9��/�Y�;��`� �f��۷��I^�ء*��.5ǒ4�}/s�x�]-��[Ew���jq@!y^"�	�o �U띯Y��%�m3�5<�f+^�:��Iv���ڒ2��6A�N�'���W,�M��'�fg����y|K�XX�-ߛN����=��S`��ޯKB��SN��ʛ�a-��g�"£׮��)�f��<r�g��:$h�"76*��/�N�I�1B�6��w�)�`w��96۹y�"t�ՎsSZ��FatY�wɖQ��X�5�*������K��M��_���ϋǒ��Kڪ��%v�Q3R�ax�&꺄�w�|����Vz�am���6�s��kl�ܬ*��/dJ
4!ʤk�H��a��݁�:�a���᧳*�B�	��s����F�s`������9AȾ�ni��x�V�o�͚��*d+��U��aЌj*k̅^#�zkqH�{{�m��W��j��^#�2Q�����M�!�p=nƞuwZ/P3yL��R�C-a�W���{�U9M��~���m�R�*�ּ��̭�YrY��`�[���&��G��*o^���;UY���D��UdҼ��x���sQ��#{�Z��V���OSt����1��l��F�^�hΥ֦.o!N�t{��\x��j��;}F��(�%�C�ڙ�}\\��]��P��`ԭf�C���^���;K�tA��yжwk��ɠZ���I��.P~gk��Y�:�x�;PT6��	|�2��Zh�x��)�ݥ1��@���͘4Ѥ5P}t�`��u�j�������[:�;1.�\#Y��)����@�Q�5�8��nh�ٺ��̣Ѿ�%f�D��"P5��4��Q�~6��ӛz/��č)i݀6͊�#o��Th�c%�� n99�G4�JFv�u{}S�թ\��o'm��/3���M��,U� �-�5��!�Pʬ�ұ s]��-o$��5��淽3g �멋�S6˦J�|����yN�C�(�M�J�7%hXoX�*�|p�#i�k(Ӆ�Wt#=beKwL=��}P��Bt���ʌ^�pԡ�ڜ9��7����Z�<���:J�x�����i��J={��qه�N����HFn��i��t�$�1j�v�T�ۚvZ[�h��C�Xn�v��%n���:��8�dw|�Vv*�z5Rn &ɪť�:�e�[�Mm8��qe>���e�U*>kq����I����_:9�̵p*#�À��q�#�;$K�a�5�+��W���`�n�˜���xD�Y��P�#f50ѽ,�V;��#���i֋�k0�)�x��ܱA��Ԧ�.��oi9n���2t����5&2�.�+�<�AAy�qv�M���E=u����,����:ق�_'1�o%Xp����qHZ*�l�F'8�֊g�7P�c�Ju�):v��r2�B@���p	���ڕz8_��XUJ��a��{k�7Y����υdXv�Δ�7�:�ew Ι@�Gx;����l�ڵ\�#z��쫵��>f���-�0���[tU޹����ra�U�|y��;v�u`)m�e����è����I�xD��۬F	}���`��=��j0��=��KZ�C.4��(�4
�}[aQ��'m��k�Au��Q�[��C(iF�����y�C똠@4�p���	��	m���wr���tۏ�I�l�������9�?�B�n n�C���(��pη.ȼ��f(}��?IFƮ�)��+UM��K�@=&��w	u�6���*b��<l�,꿹��z���^byQЖ-��Rvt��f��x�z��M�|�H(����X��/Y$������	Ȫw �frA��gl���opoLg87p�����Gz��Ë��&=<b*�K�t�΍U��$l�H@�B!�e��L�m�b��J�F����J	m��V�P�YQmJ[`�KQ�B�eeE�UjRҢ�E*\��Uj-�e��$��b�R�s	[Ze����X!PR�kX4`���Jl��F�mj*Q��s2�*U�J%Qb�K��Ze����PQ�Y��ˈV�3+\p`�����+b��ai[C0��TJ席��JZ
�A�ie�����Q2��m�j�U�Z��nZ���8&-�(��h����*+n8)����\����2��7)DR�[+m�[h��1�KmeK�G���*"R�m�
�b-eTT+Pm4-�TƦZV\�L�kKD�q�����R�iK4�JRֲ���ګ+32J�U��l�
�-E(��Kb&8���Kj�6�
X��.!�eb3�1��1k�1�WFڦ!�!R�h��3~�����sw �5��MN��c�yY�+�9��eh����#�M���Y�^;�7Ԭ�$��x��X��A���Ҍ�t׬��qL��p�46۬�j*Z9{r�o1����-,O����w:�o�6ni����wӭQ�"8�+�v�\WR��i���}��<7�A.������կؼ�B뉭�I���~7��J���K�N�Zwj��<6Q%Ӱ=���D�x�q�o���y�g�%k{YΚ����Q��X}��`�&�s}�zW�5�ZT��F���ۤ�s�{[Β���{@�U;M��﶑�Z��u-K�ړ�2�Y�I�V�v��8������,7w$�d�����꘍9r��I��M����cYK-x���v;'VgAN���E2�%������ahRB�t��7��aa+��Tl���	����#S�ERP�I����Ў��ץ(����;Z�J�PQM�������襪p�	�W|��k��C*���QH&S]�f!���8	7f<����J��hr�.�el]Mfk�vr�a�G��
S32M���Sv�T���[z�%}Ї̍�#�P�ѫ��ᡮ�,�;&}s*�1G��;#����-�C�ⷨ��%r�9q^~*�2{���G�ػ�����|�rKx��l����}�3��|=:���d�/�1�Z�u%����{����)F[��~���-��/r��t�xP��W��<ͦA��R�JӶ�D.������0ij�\�Wr�v!�	�4�J�Dt؀q���Z(d1��Mn����Ҭ�i��`n*�hkS���1�3�.qJ|�<�_���F��k����:-ګ�m���9'��Q��4ZH�=82�u��f/6:��tf�>�q B3��4R�[\-�����vhi.��v�.����+��;�=�k=Z��p���T���UC/x�
����$,���,�׳O�\�"�l�=�+�>�,H�^Gw�Q�zrX�M��r���o�O���I��5YW.{"[QQY��M!�F�`t��WY׆���Ӻp�x�M�:˂ ۜ�v�ƈ�9o���Qrk�փ�]:�-x�m)s��$�,f��4�<�Tˉ��#O6+���ܯ6͢3�]/`���c�ل��s\Ѽzh��ݲ��A��JHRc�'EW��h~٢�Vӹ�ae$ܣS+�4lS�����nظ�b���v��<n	�:ig�i��ЁB��v�./���F	��(�`��Z(�[J�cw��fuwW�ی�ھz�����X�9{/���U#B3/%(Yݦ�;��Q<Wh�c�o-�5�&���lk97������?)hK2�訍�5����-qF;��%��l�D��l�O�s���Ȱۅ��]��G���-��>]�o�V���pc��ZYYl���s�ވ+/p��d�\��p�8{m2���� b��*��ؠd^����i����;9��إ�����Bԕ{�׷=m���̍w�/�2?���c�՜�]K��.�թ���Z7��w���b��E á�T׹��t��0փ�C��R��N�n[��Ju3�	����@7W�s�$#��:��#m<���m�(��Զ�έ��j�\�ͦ/�\ Q2H����N(FmM鷺[����edO*��.��*� ��:H����3H���٪�g.E{F�	9�r#�8 �=�〉��KE1mĂ��J�tb��T�@N�swv쳼o3j�Z{��'������5{�����3͹��m�y�N��g�.��^ͷ�9��ւ�'��oW��R}���x�6�C¼��t9��O�e����m�)-�/(!F����m��R�}�m*:0�u(h���⏡n���z{+��ٿa�x}Zvw����p�x�0�7ɶ{;��aN���IA�zD���s]��.�L���R.��^��%�J��)�pr�ɧnt�Pvy3.���f�R�̽��f�</ ����kS����G=�[�f���c9%�R���	�n���7j�x(�n���Oҁ��'�j��Ħ�w��s��r�TV^em�w,}{�K������N�����Vw��K��6�Dʊ����e�!Y�o���E���m`j^��}7�y�i7�!����K���f����W��,�Ev�j��{37�����(���B�tj
�{
ǌqn���a�.̙��-��:`�)�>����7tޔ@�����h^n^̚[���H�oN�`�$������
qA���J�	n�A�g���m,��N;�ýo'�X��ǁ�ٰ1u!_8!pdh_JcP��G��ǌ%�3�<�0^��m��X���ܳ� �^���?�\�;��c�!D�P<v+�sSؾ�-%/u�0mg�E2��A�P=
^���'�A{q����F-[��4L����C9�_[�.��*)�n&���Y6�T�e��*"4�;<���E��v'�ͯǷ��n�d��1�/�固�v�Enhma)"U���sT�Bwmg�b��o��бۨC���8&�{|{����$d���xTAf����ǃ9���ۮ���!��UF^.I�W����o�u�
�7K7��N����nÏ�}]���`| �.�T�ag$��O�vV�V�;NÝ;�������\u��q'��(e?dѝ�c.
DJ����T�����:�z?N��v��c��'`yӷ���ј_Xm�,uHP$��M]t<#�ЛW���sV	;$�r��)E�Qr	��!���i| <�5���F�*�V�k	o��h�e�γ�Ee�\����|:,ݼ+W�)�mw|+�W�o�_%���k;N��աI�-��� SmԘ���mb\�(W@�N���urM�Rk:m�!n����t��O"XGua:k�SD���d� z��BH�������m����"=%v���k�D���h�a�ÁK�x�^X��n��Q�[�w�39'-X�����ǭ��Χ���+�M�W+<����5+F���`�.12j�U��6`�F�F�1�
{m,�����Y�w�x�ȺI{���r����lOQi3�ǚ$���]�oK5DK8[��N	A�:���ym^���Rl	U��sz�q�k9C���-~��$��MU`uQ[^cksj�8,�F��y�B��[���3J�m�j�,<5�d��֊x����dߑ��.�τ�k�Vnb���Uzm��E�47����k��;7�wwTpBe@1=��Tӻ�o�h�]��~�՞�\ռC5�o���u���,��q������hڜ��[��1H��})^��٬�[��fb��]�թ�緫\=lR�7��J�7q:*�{%D��!����9y
����hg����|�߽�U'X.Ϭ9G�#[C#m���Ԫ��C��Iu����ebu����`�`+����zW�/�m�g��׾�dd�I��]����y�(����"�i�� �C�����"ͮ��)�w�+j�3~�Av{�����UO(��M�.*�S����8���^���Q�c'�r$��ǁ�`����um4_a�R��x�l���X=^��6P�<.I�饝4��W���ז�F��/g����%9X˓�ٲ���0�SK��E��÷����ϪJF���%�,Y�`�m7/e甘@�"���95��W���ל����;h���f�4��u���Jj\P~D���u�KoLE�r�:u��%���|�Ǳ��D��l�O�g;ٿbW"7�� 7{��5mL-�걯�2��t�́�*�l�����,�����<4��N�#��գ,=��Cù���u���� Kl:'��۝a9B��S�L	��A�b�;&�I�;h���n�H��U�/[}�f�X9�\@�$s=��߲��[�k����9��iee��K�;d*T��v�����H�`��!CC�o}@ު���)~�$';*v;(sD��c"T��J6 ��wq�Y�����tNW�s�j�3��XfzB�8	�΃���R�h�Z24����=���q�iO_��"�%�f��l�*)��q �2��f�1S^DEQ��^�a���J��h�Y�7�m����[sO��盾���DnM�sW�qV���.4�fH��P��'���xo��]*4w�ɳ~f��
G��1,���b�o�9;	B�����/eq�[,M�0�{�d�~.TE����� C���RH�zF�(�M_��R�%`���Vҿd�z�&I2�&�]/����(�y����;s�{G��z{4'N���6��{�|")9�q���]a&^笫�P��#-'���kjdJ�:~�a��7�.��jz�w��s&f��D�����?y�����S�e,9�wQ΁j#L�8�&^��	A����ξ|��涡�=	U��]�����	jƨ.�R��S�o�oJ�<��i[tx�i<Ż	�aΝZ����`�H�zh���PB�5�����.*�6ShJ���Q�i�x���q[�[��E�Z�[Ǹ��#�<Q�Z?[VE���^��N��	|��t�J���R3RX��/5�-�Д��g���������k�׼3r���.P{�ͨ��o�&��\��?r���Ta��A�~=��3ބ�"�Ec��[�>�ån���Ro�lhw�X�#B�!��U���sv}Ǝ�(�/ˠ��ȼ[m]�gsc|ӁR��CLN�ґ���Uona}�(��lвW4����؞���O�x|m��༴2�� 5���0�M��}�����z~3�VipW��*�J3.�lR��fS���i�焫�F���4���4��nt������t�\wh�]��OGv��κ�ݻ�XS%J45�C��ǳ�,�{��
�6E�2Ǔ1BԠ�t�a�C`�kr���VmL<[=n���_8�nC��(�6+$�i��Sr��ϩ�Id{]ELw���A[JkM��gf�0����2ߋ���QsL�� �u�;��V:�b�M�{��s\����Q�iK]<�jGh�wY�;x�:j��E��:���v��s\/2y�E��R8�z���>)*CEc������ok9�W��������zu�w��#6u|��}��im��(.�V�V��ӷ:w�7�'��J�KQA�6���W�^���S9]J�K7즖t�x9�x�aΝ[�'���\��3�%�Oy=I|�#Q�B9u�6���G �-޲�S��7����S�l����TC�"H��W��gm���ˆ�T��XJ�7�q��
ƣ� r�^)1K�PЌ��)E-ܘ�K�,�#Y��A����v���Ұ�W���%r�ˊ��U���-*�Wi"ܵ׬��Gj�؋�ieg���Vs����E�J��O��\���(�[�nP\���tp
U�"v�t��lK{h�`�+!;��W�N��n�ʹ�\u׬�C��:���#v�]����Tx��n�YnA��ޖ�Cb��N����X��!Z�夫s�TPj�$�;b����iK.$z�!��=�q�D��,+��z��S�7m������.���*6�2.�;����Wu�kS�~d��e�GZ�� u��֖Eq�]G6�jY|o��d�v��uh��$f�/���X��nT��=b�ٓm�T�N���2��B��PW��j�BDH^ʽ�o\��{z�ދg�}�f��7��;�*�-��oc1M�J�=�>x z��F���f>��Q([ܖ�j)�������sO/�̐�k~�َ�ub�mfP��P��r�Ӝ��f��U�)���xrI+��ڑA���p�r���fq�kI��n,Kq�ݫ�&�Y�_��X��v�,�6:�)X�c�u�L�8�J�M���y��Λ��Hm��"<-�`�Bt�h�6��[���N�GT�C���OjDw:�}aJ̸3��j�iR�ģ���m���5�Ϸ���6��Ѭ#�#�4�+�ծ]!Rsi�K�-&�&5�{�G����z{�ܼ2=:�®�r@,_D$3��.M��F�ັ經��YB`����]h���,:���S�#�*"8�:�S�&�az2)��o/+����/o3�`��S%j1�Yy��N����Q���:���u�DW:sp���+x��99�r��1U�kP�Q�*�U,�ut����Cf/[��A���j����T3!������Xi�'�=֔��3�"�>�2&oq���Y�]�*�`2�.�a��fQڼ"�k��(�������}�һ�ū���1I���B����t�3��͢n��h{�0Ӱ�h&-� z��WL�^2T��9;mU�`�h�1��
7X8�����TgAv�R�@��s��vE���F���mh�Y��E&r��\�?���4��kY����[I����ؼ�y��|���G&7���wL}��h2x�쩒:X.n�᫖,w�[�ȶ�)g�ohN��X��Bո]���o�]��ԩ���e��GuG(W8VH��wF8��nRN'=�뻽ԵFλ�� ��5�0��X-�WQ���wYBƽ���B�R��LBm[����7�PV�q��򱛷�D�i�[5�v"��9-�z�1J���}{6��;�{�{��%�Ly���ۂ��#c8�']�V��f!��+�8���]�!Xn�����#�i�OPjk7+QP�xWJ���&����w�&�;��є�jP�5Ģ)Xw�{:��H5c��s���Ty�����5NQeh�P���A��5�d�A��o_�0"?4,�0ײ�Q���{��ݵe���K�r8�-r5�0�sdi�M�S������BV#�͊��mج��8=��ͮ"��_ P��lY�1����h�R�*6���YikPZ5""��%X����Ĵ��k�-�V�Kh"�ԍ�ڱ��YT��6�V҂�m�Q*5,eR�,JZ֬h�l�liT���KBԬ��Q[m��Dm��mF���ZU�Khյ���4KB��Z�kk(�QbYm��Z��´e�PTkR��Z��bQ���ѶШ��m�TQb�bִZR�B�[VZ6��Z��e��K+j�kkQ��F�R�mh����E��D�����[e-,AQKE��m�A�mR*���m�-Z-T�D�[Dk����(֢*-��J�KEVʅc[m�j6��R��h�Yh�Z�kjШ�-�����h�R�Z�Z��UJ(�ţ*-���mJ[J"��lm�����Q��hU�Rն�V�UZ--��5�'T��z;��]a����ҳJ�3��%\olp�z�5AҮ�}Q�E��YX��ǭ�k�[�l�A�뒽VQ۴�H._

@���r�i�l���j�	g7z18����pr��}��ĥ�d1��7]�3z��z݁������A��F�͠�n6yX�/RH�An[]���9����bЮ���:�x��n=; �
��,ڮ-.���E��ʺ�Ǫ��i�򫿽蘮���+�����6�Q�=�9-�d:�a���*�	���h��W}ʮ�i�\p������ؤJ�2M1�dq�8$��Y�][5�dW��wg����{�fg#ڌ�J�H����T����G��	��,���{��*·u�b�i�=<�I
L`�^�Vr��Zf�R�r����'�y�2K�:���)�s�����J6[�*�M�M��+k]��hvL�<��u岒��sXIX�Ń�1��!t\�`:k���_x
ޢ��$��HM9�컷��s:v���{-�Z1��=�����k<�$��R,�����D/rW�=T����fͤk0�*-ѝ�$��+z�ч�0[�m�]�%K�d�+r����'qe�O���⃨���C�m���GN>���~>��Si�+����R��z�h�ЩF%c�]���ˁ��D��j��(�5�6������y�hF7N�����S�]���L��;��$ߎ�7��3I��_A�g%�RÉ�y�r-�#���޴RGɛX�5�*�A�`�3x-�Wy���`�^���fb�<7N?/�3R�ix������w�|�i�l����]����o����յK������Ɲ豅실!�6}@ȽV5��k�e�ȼ���VZ.@o���'��~
�u*.�]�c�³�+����UҤ�Po�F�a(�\�_'f�����-1�%Pѐ��BO�f�{�n�}�R�ˠ��5f�i��*)����h��w�����1k�WE���@���AK|{=Y��w:�hq��m��v���MC
P�j���5�8u���:)�S�! �v�%m]������.��6B��i�N$�RHɋ1ݳ]Blǅ�Qd�	+��V�2�̔*N�-��^t��K-�B[��*�l���z�2G�����XG'P:�u.}�$�8

m�e�M��;κK�F�n��F�r�P]�����t7�Il�>iw�����Y��'�>�p�'-�󦒸������zq��V�[f��҂�̝��\>|��mw$�u�v�5g��y����u�b
�a���;r����6�-��.�cmE�ǈ��+�G�N���i���2�>1B���N���gˤJ�}\�GZԏ[
O_��Y��I��M;t�Ф��ԛ�^����Y�,Q�,��n����&�t�<�25�-�n;$Ϫ�D�2�fVգ��֤���	:�$HIEYj�~Ʈ��O�a.�A�j�xMj.;�<�$�R*��7r�)0��-	]S�)EY�~q��-��;�dCn�fd�KQ�8�WC�G&�+�~m��Z$jV*�KwMJ��d/vaao���y:�$I����l�{g�����D��|�*��]kvrM�6����]�8br��]5:5K7A�eff�4�x1�3-�c�#�$�c3���/Zy�T�>�A܍h>�@7B��� �.-y�z�Y)�VwJ�N�:!ɐ�Fm'X�l>��p��}΢̋&�h���u��ڔu���ů5G��3Wr��`z�E��}ȼZ-��K8��������N�v:Y�k��Ze]n��d���q�k�K�Wއb���C#���Tq�Vs:J\�C؝բ�hbsB��X���QL[p�45��D��;�c�$J��:DKk����k1n:U�v���Ĝ���¨9���M#y,�ݴkg�Qrȉ�F���Xc�ŷ��S�����U���g0�:��h`3�,%2�V�L�OO0v1�8ݹa�G��w\H���oy:����-j���!_i���Xn���s���Ey���Oa��w]�`�y�v�=F��+h߲z�e��9[g�5�i�Ӛ����.��ڠN55���q,�\�
4$�8(ҿd�~�igM'��<Ӱ�N��L��WL�-�����v$�����1�J�6�~��E"}�[�nwX�����=��YY666�mNp�3�q��خ����Z돭�#� ��~g;��C9K�ǳ���@�����90��R�fa�l�{j�d]��Wj����;|tCq���m���e���Z��-���9��7�Uj���M	1ć�]�A�EI�@�H��$H(�m+mJ��	r���}�q��7�BZ�s�,^��&+��B�y)B�0.#����%�6���	����J�}
Ƴ�c�Y�.)��F�0�h��##�ש�MqE�I�K����ie`��}�9�́�܉J6�J�6��_^�%�d�$����Y7C�Ug��9�-,[�m]�,���D.��9%�=�M�eq�҆E ��7]�Aީ�^�`�m`�� �����R�n��"�5��͡���ߑw6)�:kuH����[��;�7��k�������6f��1�*�CXsr�L����u5����e��,o���6&���n�>�8��qτ�u%Z�Z���4\a]�>5]=ؚi�={�ϖ��ߪ�QޢzW|���E�3ª.Y�^��z�#��]�޽�]�"ַ^�xu�AX�V�V$z����Y�����;�*@x;��=q���5
֚�{\�T9�nv깘�,��jE��k��\Wb��uCR4��R��l	T6���{�)�Vɻ�Q����U�e�4l�C&T����`��u�Nb�ҴFJ�J�����~{^af����Z��CC�T~�(d^Pb�N�y�ڶ�e �+o+x=�K�5*GOc�x�DO�T�,^PR��nL�=h�%Gv��4��2z?E�$�����}0��8���U��5��!bxй&��C�pxR7�ҌƏE��+����[��i��@rv{J(X=BF���%̴�]"�b���J6a����So9�E�8�9�i���y�&+�va��3�&j��-v�7����n�W��W�5`�#y�X�g�J��65��mܺ]svA8�ŋt��ƍC�yJ`��4%��<��3x-��琓��[1]��ٹ�����UKI\�	:~.�bS=�u]��zc���ʇ�qV`D\�oU�h��rw�E�b{"�r�H�z��[�KS�L4�����k�E:Y��Gw:6��Ye�:�-@fų(�7c3��*�f��`�.���rث
b9fN'�*��u��j'�K}���1JW����<������b�Hvg3�]��9��v󘾑Q��.��l\�i���"yĄR�m��y5v%�x!�	�����kuey�4�\Y����)�-4�J2_+��m`�� �U�w�W����vG*�1��b��Vc�{��.2����}n��g�E0�õ��:����Ӕ<��i�f�e_z�ݩ�k=Y�3ۭ߱�CN6m��v�j�Fe^磲�r��<�kU��"�Ə������� �J��{�P��\�җ��j�2{�r=�^��W"�c�����6=���@���Ll,�9t*���ȶ
�9�g����g:i�G!VŇ��w���쵫 仆/D���0s�Fy�of�mSA�v�N��ѕ��U�������[�h���%�6�?JJ������D��S~M;s�V�'�秦K�4�mL��� =�����ު"�$�[K%4zm�!n��6�ƹTƅ�`᝺��\Vqh�ɋ@�<z�A�n=����:e�f�Z"pH-]���s�<��{qa4�����y���vƗ�ɁP/*�rk6�c�$_d�X_`��Rw������$O�J1���9��D8H���c'�ӋY1��=�Z�})�r�+��ҊZ�~Ư=o>9��K�QGtun��eշ�������K뗁I���-	]S�)EY�`�3tI-��'��F��iOV�QH�����ĮE��?���L�n��ۈ~���{8�]�XƼ)��[.��n�o؝ȱH(�!ʤk\��u�J�SY�D���w�c�r.ʶ��,��C��
������S�)M�;0�=9ܻ�C��aY�7�h^��"(�q5v%���9SU�6�T�ά��h����,br�&�^Vm{���W���TS�$��o%f'}����b�)�a�hD�#UMcx+6�b��V�7*��e��I3}��K6��Fiu��n�l54Ȋ�F��=�h���.��G�3�=�& ���Fо�`��k��]�5mdp}��:�7o�����m6�Q�ߊ���)�xGG9�:�`]L�G��pJ�N�*��5Kt,F�f��W�N �=���.�Z�]|ken�d����YȠ�!ŗv&���2C[9h޹x� c��6��P�s;0�,����9x���Ca�Rkf'#P��R��v��D�k<�y�W�.�/o�m!Ƴ�K��M�sRｴw���C��E��-ϔj��&�c��N��ӝ[���Ӷv�q�^+�Z��E{�>P�Q"�b�M�J��t����;9�s�x�Ř����籗�QKc���o�2;���i�a�-i����\�3�ͧH��"Эo_j������/+�������K�&`�Ҭ�0�@����z�����P����⮌u���p���֙�9�ڭR0�P�gTHU���s�ƺ�H�N|�c��yA��L��\��e
���Om��MD���FF�-Vt�О]tʌ�jڸ�*o*⫙����nP�}�|iܴ�nIB5/�ᅈ�����NY����C��9�3jpjw�C���}���g�&ɱ��SF��}L���j }*8i��/Bv����
.�3�;�m�cV2�Q�V��(X��tH�APP+#F���V���}����y��:wU����P�s��o�"f�lGQ�v�����3��+�������0T�K��K�nevV�c��(cX}��Yb��ݩ�˿��������Re.[/j�+�.vX�f�YI̓y�amZ�)o|��\�[��+�rE�$��Yb�	t�.X^m��H��r�#�$��9�7`�5a���W���x�R��/
������8��^�hk�J���d�f�ȳa�B�_;ȹ�]e|Gi_+�5��<<k�F�΁s�$l��s���h�Z�o��CHt/}�f:< \~����#�7	,�CD?�P��Z~��\�u�ʓ6�x��nq,R�{���=R����r��t�Pc�b�bxS��f-M�D��X��l�۷׻rL �=���H�/�UY���6б�.<�m��)�0ͫޗ�Q۞T7�3����3��J���.��&+iF-��En�`�AI�U�8�y�m�K�	�a��$��r7�߽8�ل�Ԩ��C��ܯ��Fz���w�tM����{���Q�u2��v��Ho���񭝵
��n�/���N���G*��y��5���R``�����x��`wj5΀���x�Q7���(���P�ۣh7c�LnH��E�ֲ�b�j��N��i��v*����pJ��Xf�x{��{����H@��BH@��	!IHIO�BH@�BB��HIO�BH@��	!I��$�	'���$����$�	!IHIOB����$����$�p$�	'�!$ I?�	!I��$�	'�B���PVI��r���@�6` �������&���DT�+�2��T�EJ�U$A"TJ($J�h��(ш�46TU@�������)RQ@�EJ+U�JƑ�Ihi���n�X�R�-eUl���k&����F����Z�)�L��"��kYm��YYT&��Z��Qfm*,���z�$�Zմ���ͭM��ٕ���5lf6dm�BE[j�6[kF�`h���jh֦�eLV�mj��j�f6L��6��B���Z�3g�˵c5�j���  :�ݰ��kv����\����h8N���vۻ�]���.���;�Ɔ�Gn�6�U�[������ݱ�K[Y��b]��m��]�t�S�K��kuY�JV�3m��)-�ʼ   7x�(q��6:۶�J�we���Ν�[]���k��:�SU�eۤ+KjS[��is]M.ڎ8�b�δ��-��΅-�k��RabՖu�R�BRԘՒ���  ����gs-�N�uN;+��v�v�m��Ӛ�ӫ�CnӮ;��nv�m6�t7`[u�ͮ�r2�hP�e��(PP�B�
���(P�B� P��9�(�
(P{�{Q�f%�Z����+m[�  ;��4(�
�w
��
.��B�
(z7w�w�P�w�v��i��.�l-�6�u�C�Pmt��k�5N�r�u@Rj��5���X�iZ�ʆ�  ^ �l׻.��t̦A�whEK�έ���\P:WnZ��k���껝�u0*�u�ݺ6�@]el�*�E*���m�  s�^�ij�����h
�N�@;���G@9�s���\�� �� �;�n��U����p�M�iT��kBe�jڤ�  ^2��7qp:�%�ttv��P���Y��ڥl�t�-�:݊��-�Қ����ua�i��\.u�(�+i�f�m�V�m*U���^  ���ZR��Ve\e�m�E݃Wt��UZr��uwA��w-��U6�:�2���[a��L�ٻM���[;���GwwXf��vuZ�s����jۻS�`m�4d�EV�I[Xm�   ��E�n��U�[wdiN�l���]��U	J�wv��c\�]�+��[VNh��*ۻ�ga����w[�Z՝u�n�;)P�����QL�I��$٧�  3��v��	Z�u��h�5�Uݱ�;�TW�wm�ڲض77Z���3���IK��l�ջ��v��r]f�3���ӣuf�s�it�Z����RR� 4 E=�	)IM�h����&Hh=@ �JR�  �~CF�R��  M$I�T�z�`��4��+�Z{�DcA',DM�$\����5=W��5�v�[��w�IOkԿ���B��H@$$?����$�B����$�H@$$?���`�g�����g�q���x"8�Q�p�9&���/��h�J��HLӉХB�I%GF�'H�A%�`ՙ�*��:�wO\,�96���Hbu�qGVrRLN��[���x��:/
�I�Z�4�(rRE�����H0�z�ff��u�,�%NRP�35���H[{����eV�)0L˸�b��6�`Q[SX̬��k�h>�����Ci5�M#��1�AT�9�ȑeb�h�+hh.Q�j���aĦ���H�v ��1Pm	Y��j�谰�d��f�*F|U̺�ܺ��J�*��>5�c{�Yy�%��"	�vv��dƂY	��Za���4�b�WSj�`�Y�&��Q�f����x�YB�M��0�/ncNƫ`���p��^nW���	KT�)*ڬDU��������V֦�آ3m�w�s7<��,� �%X�4���r�0b�����跴̹a`A�틠3Uܘ�=�wJ��Ł��ڟ&M���^d���H{�6�PUl�H�cz^���+F�{�0�7,��[k��'koY�۹ܷ�Lp�](T�f9W/3���jcY�Ū�#�x�5D"���e�x�[Щ���XXؖ�-�B��1���z�c�t�	�}�u�*C����Y-�W2	N�:F�̧y>wk��^Cr��)0�7�։,�8F]K�X��B��i�k�p<��ƆYG.���y�HX�'9 �s1+V2H�iӉ33]�/�XA�^^Sb�u�|A/L�f��� [Zp�!U��Y˒�6Hz" �ۉ3�
)�t�{Q�뚆�7ѵ��A6m�p�i}u� ����"�Ѻy�W�	Q�.@����߅���I�e���k(T0���V� �������+�v�S��Kt�5�(����=�
��+�M6�Q"s_fD$��m8�jKmژ���$^*�B��y�VY:����C`�h(��kL����&�,�M�vv�E�Qz��L��̩wMX;���y�v��4���z�kU���I�X �R֢�;����Q�d9G�ۄnGV�sj^B�8U�e��j���kC5J"�ݬ���u&۬ӮH��ۙ�񫨤k%k9�ձ��n�ȑɪ�i�t2��H�>��<T[��r�ű�i4�	�����4�V�KF�(:#�-#��-��ko`ʴ��T�L0��`�J8h8L�`�
�CYv[:!��f��{H�
�B��`n��/��`	�w(Ȁ�eոݬ�)��m�����s��t�X!#�^cדF��"�'A�e�â���lkc�C��*��$�g32bP�t"���a#�TT�l�qe�-�Nm[��&楶�l�y0=��J6�Ih��0��f	�ek�%���ӲUf�������#��c8��S�˾8.ɠ�́��T(B2� ���%�Y� ��G
���A��6�;u�K����cm��2m���w��Sh1�RF��L����5B�llfN���e����RJ��q�*ˆഎ�YE�ڥFZƀ�Tz�6�ɎBܱv�έf��r�#`3^յF���Z�fۄY�3��z�mX��-s�!-%Ye�XQ*�I2�V	�&(�kb�ē���z��L�5Y�4.�5�V5yr��FH]Ы+��W�m�
٪����C�m����Z���m�o�vX	]�@���cB��A��lX;��p�v�Kյ��y�Z�$�)�+�R\ Ԧ�.�q9M��F�՜['�;���Í����:�,�9BL�t4�(�v xF���K-��׍�N���̆���VԭOA�omB�!AF/t�]�A4q���,���ײH��W0A��-��RU���虘��7�b�V�-˻z^C[�!�ej��1v����6.0��bks]K�z���f����ń6����O��ei̒�ToQ��A�A�A[�v�Ę ����t��D��,�F��k!�P�ʃ^����0L���eG�bB-6��Z� �c�T � V��Qۼx��%��K(ޔf:)鑑�A[��*f�������B��4� �D���U巋]Y��ojak��R^���V� K5��R��"��N�4+�WXP�T�9tN��*z٨��I��1Q�N�����6�j7kaՁl��Ĭ9E�.E��_����e;�*ZF����e�J!Y%����1=`�)к�x�MK@��@C��^C���J���mJ��V��6�ئ�[�Gj�9
@6�ߑj�N���4JIm�V���7*P�YkHi�2⼘e�ņ�S�Ts��Yn��V�!GM&�s3A����[bŔ�x���1%c���%Hἔ��H
�,�F�+^!̵K��qˠ���c&��"�4]�dk2;����7K����Ԙ�v�WQ�Z�-��*Ž"�r,H�t��i<Xa!12�a?�S���8f���f֦�9���XkrdnT"���>�xeK@)�h3I	X�i���0#)�kNL��E�_�2��+&R��[���T��(���RP�N[�Gs	��֓f��W��X�Ж0�ͧL#�Y����j�5\��5l�j��kR�&k,eRzoh\5e��n�+L�N;j�q�l&��,�X��ZUl�pIH��&��1ݻ�*��#j¦v�]�nΑyܬ�OvX�wd��qR+N<��H�v�֫�k)�Z�j
ɤC�F��a�8��&�k���t�]�	]á�e쩙@
�AV)\�z��@#����[��E]��W�Ti�OlZm��bP��^\4
���JoZ֚ݥ[���ȐrVy� :6�V(ޑF���*�U�t���{��������o���J�ZIOZ6,�B����S�`cj�JG$W-���r���n��e�yf��n�D�	����0bT���yb�]J�,��kE,����]��,s�k��0XA FZ�<g0�Uu,�F��։C�j�7I�Y���(b6�kS�B(q�R�R'Y��+�	?�XJVՀ�
�&F6��j�(mލeKf��@�w6L��) ��I]�Vsfcӗ
��亡�H��ndn�9���s<���cbX�8v�
)�(�g��0�@�ݺ���R Y�q�]=.%+��wJ�@!�ղ]�@�	gۥ嫷5씨!�,�Q��g[���w���2�:�{{�`�Y̖�<P��wcXݺ{�Q��E.�H]�N,��"���@D3/6@���eC۶Dt�+eg2b�˵ Ų�!�LÑ�^'%A(��;�j@rB�������a�*o,�LL ���1T�[l�FlZ���am��٦�1�Q�`,<�!	��]�5�v�K��{m�ߐ��ʺI�v34Q��
 l��%�n��8,T�VT)Ӗ1h�r�452�v��7��[�]�R�ս��V!�%��ʆ���Z�Kmi���y�E�y�X���b��ۺR�A�r��R0�eh[��*iy/&n�ɺ���\��ĳr��JHaZ@��3��X�%�D�$( ��]��#Yjfd��u":h�r�A6��04����@�ܼ ]7�>����3);{2G�H[{(�p�tn�޺1X�2�����3[Pe�t���`�p��s7@���=tr�m6,�j�dA1`8��(�m�=��x �of��t��"X��B�W�z�,�N�Z�����^�w�8�����,:��FSI����k�N�[�uhb��P��m;���|{�1Lظ��[؍�4��,�Tը���7m�h�W��͡�[u��8�0�8G�:�[֜N��j[s
L�n�"�\#.dۤɬrŝ�`w���&Q2g�Ì�ֲX�8�k%<��/�uB����Jе��LL�4.���%�ҳLE�vUmh�Le��")�O�U����X��
����ͷ�/f})-Yc���SÀ��?����/2�J�����lh�ӕRKlmb�V�vn���B�cP�d��q>G�0�YO�U�b�����[��n�0����geX4vX��iJ� Ď=���i�7N�v�NY!+ˡb�76��:FZB^)�iB��h�i	�r�+�1*�
�@�\p���9�2E%5)<9��csuT4��g1;U�1֜��)���
���,d�fS6�	�dam ��۔.�4F�w�QI�U�,_Ck�i�惓v$���f�*/뱙�ܻș%�o&�5�i�Y-��YcX�hh�a���]�kr���Wi����`ԕ5����[d���@ռ�l4�nۼU+��h1X����)�Ů�]�h��trn�
�iyM��m��
�{+��3�2�Y.�F��y*��:Ӈ7lf�۷��MTK7`9-P7P�����Y36 ��Lf�4ic���1+��XUn���o~L9*�m5^�b%��ى}�
2Ľ����g��S��6-�J%Ll�Q$��I�JR˭o��*�ڊ2^Z�NE���5w����M�D��RF�Jv�=H����t�{�ȱ��"�{F9M[ii�Ԥ�xͭx񭺟$H���$�ی�cl"t�Y#r�C�k�b�
/e=��*W���8䱀8!-2/+(��a�2�8.D��ܑ�f-z]KLIj�M[VM��J����.��Y��  �����]X��`��O!�N�]�:�4�e�r-�$Kwts�"P��j���R�z��/��f*�Y�Q1�7dٔ��Ӄ.|*�ԭ�ExC��Lۣb�B^8����8fԬ��A���B�T� H�[YejR0a$�T$�r��6�G��-�7*'-'Xb�ܷf�
oU�z��4㿚�H�ˤ�mU�� 7�V�ݳb-�w4��)au�MD(�e[$�
��MB�a����׆Ҭ��Dl������4���6M�N!��m���H�kw�ue� �RK�d��dLe �
 ����d�!Q�2�j�P+X����"�K&c@b��(EЩgj�V��v[l�����Y�k�/H���a2���;�?�1�R¬��sl��\�s�\��%5m��&��d�F��W2�V�fn�V���M�Z�hl`�f�Ӳ��6<�H��mǬ˨ό0�ʲ&��*Kh�&�\QkVrŎ�S5�,;�zvۢ> �CV��EPk�rՃwX�Y3� �M]�iZ���W+h��� �n���)�,�S)B(f��Y��*�u���
a0��"�T�M��jZӢK ]
*U�ܢa/������9��ݵ���4��	��LhXZ@eح0�6��Hf]��"���&�-��V"X+/ZZI�M!��HwD��h��kS$�)O#��WwaEn`r�֘0S�lM�*:��HeN�
��,�f�4�Mc����B�!QL/�*�5��Qx���X�1e�y2i�5j(�cN�]0��	�u���M=ˀ�PK5�f�.���m�z�[��;-�"�8n)���(6ޑ7�uMɺ�t򵗃��w�u�.��r=@��u�{��CZ�d��#&T,Љ�c[�J:a����z�k])ݫ����T@�����vko*<g��l<�-���#@���:ۍ�"�+V&�w����l+!�1��6�/���.&�ay��j�8�ia�	[$�(�2��ojQ:���Qm����6�^ko\Ү6��m���Ǳ+�+
�0��λH�:��Q�+*�,�e4*�6l�zJq;�ulm6�o(;�¹6ҏe[7m�C-e�=8�n]Ҍ�o��a�'ɻ�aa�R�m�kr���)Ha�Hl��{YD�y�tѤ��U«�dɭ
�Y
���w�fd�J�`��]�mL[m�݇Z�TfE[�y3[�˺N�TL�i� ͬSP��i��%;�&��*����m^j�RX4�=ǘ�xɠoU�ѰG��gI�+\K1�i��n]c �6p��EYm�,ϡ�5�չv��L��`���1�8=6;Q�� z��{�Ҷ�,��Ə�튶�j�ѥ���X��X�[/�K5]M�X.k'����mm�nG��.��������J�m4�:S5��A3�R�V�GFJ�j�u:V*]��2)a(^Lњ�{Z6@�u�B�VC���rT͛�(h`�����-V�CT��ҥ�0f�� �㖷>f%5t��tSJf;�ꦃ�ݫ� %���5�7X�ȁ�`9�h4�GD�GdJ��e�h�&�{��yBTY@dv�O��	m�&��%n�[r��#giJݳ�wdD��*�c�{����V=�ke޽o^�l�XU��v6�&�L-I��[���Gq���Rz�����є"λӶM�W��۩��񥚂�/-ǴZ̬X�*�Du ��f���k(<--k(��t�ԫ1��7p�1��n�3�iH�%A�nb�hl�̚�7	����n�Җ���ti+�ӢڑeĨl�x̺���B9�ǫW�A�% ��b�4�{�6�lV=�fSG*�1��-���v�`c���i�x����S�f53b㙸u���\�q�wu��F����5 �]AM���^Dq�̬��O3on�� ���ւ��w�w�[&�t$�QR�3Wt�Q#m�'���pRm�XU�
�w)��J�waQF8LNe�����z6]<�)��mm�c���I�@fÃT��a5�H�c(�f�����1�6�N��L輲gҔ�c���][{��a6E ��a4�}����آ�dO(�����#�s��>H]�bru��%w۶�v9�=[��9�c#pm<�4�u�PvГ��}S�DcW�����z�	I���hN��[��;��f���*=V˜�W,<Q�A�z�조�j��Bm��+��1(���ȸJP�e��is��n�{�ħ$�iWM�j�nf]3��K_�򴫅�K"ծ�fV�N���w-�u)��2��SAU��Co`}�U8�8�ۼ�W"�;���h��m7\��H��-�`Ү]SA;��	k;1ݬ�֌!���RN��Z�{F<�i�YviRz�nL����j�����%���`"�׮���#�A�oD�Dd����-ow4fc}C[�<q7cl�]��j�-�R�\��K7tQ��߈�K����y��{��k�fq��9m�Ⱥe�<�> U�H���pǆ*���/�l����h(1���Q��0z%�ް��u�$���:x�F�mj���ql�9y(
�Vjn}/#u�/��9��3|#����.z�z�%>�"�WtF�}r�6h�U:^d���B����tH6A�\�D�������	�F��Hκ�e����v�'�jѸ$�TtBw�^ �w65;ձ!'J�F�Y��+ ���u��e5�m�7�R�ٮJ��ܧJ��$jR���R�r}�&�����q6�ۭ�&���3�;�t�oCWO���_'��H.�6��Ha���uרg�f�Lwq���ei�&]S
q`^��U�
D��6B��;�w@����x=֩��$��S�r#�^r���7(�;��1��W�;8f�Y����@j��kI�"2h��gA�R�5P�՘�W���ف�տ3ǯX�K1-��،p@���J:��5[R̂���9�1��(�;hE�Ǜ�Q�u�%j�q�/�ֻ�蚞:ua���v���D`�K\7����O���U\(u���<�]��M�^�H�@�9�\�J�ݽD�v�%�A�hp�d���w�`�n��d��5xcA5َ�V��f�Q�̂�MJ�o�I�����+Gn�W!����/�u����3���VЭ�]�+�Vn���*��c9, z�,b�4����r�*6H�,*é�rػz��ݜ��G��$��Z��(���곎�m������fG���MM�J��ٺ3��y�u#����Wsׂ�H�t�S,�"�.�5	Ҟ�� �y!�ۤ��Sެ.��Bu�����ɜ�c���Ќ}S^�6�D~��*f]+U;w"�LBEֵ_G�tf��<tB��pd��]��Z�nn`��h���+svR�V�mt�le����q���Uy�s�/���X��������wm��L���hR"��&��{�'u�U�8u��goۺ�k[�1�'��ͩ��(qk����f�X��x���l-Y6�3�Sv����0�a�n�\7	��2�	4-�ҺJ�j���Gq��t\�Pt�^v���&v�V�ݲ]�ؔEl���(���M����@�@�'i�ti:��T|w��5\�]�f5{d6*e����s��a�ť˺p;����_k�P��w�1�x��䛢�l��52��(]gY6�51�-�3�S��J�RE�5+2���3���r�[0���Z��B���C�9F+����1��a	eB��.R������z��'W#!��xB��r#5QӉlA��gV	Ԇh�,���ǲM��=���՚E�x\�LGk��hZ阨YvK{����	F9���ܜֶ�t�8rE�Wy����R��G��Aq�gz�K�1�"���Zv����]�����M>���]��xǽij��b�u.�2���5��d�ޘf���X>����j�a�V���2�U�����'M���}&M�;*h�-c��M�U�z򜙽ΖR-L�[���{����s9�x��yBU����bEY&����t:m���C]�(s9�J!&��'B+��( O�������Ψ�w��v���.uخ���"�:[��LVS�d�$ɢ�*=O����+aK�\OIC�۫��Ζ�X��!�1&y��%c��9�<��d�R�Gy�\]Z��8S�Cq��������֌�+Zh�[S�=����Jc�������z+�*��#9x����KQ�xp6���7��6]�/���K�������M�u����Z�5���� {X��O�͐�)q*/(3�z�;��K(��ս¥����	����f*j��	>�"0^çݮVݼ��:�ł�.�xt�2;��i��I��ޣ���������h��p���\7�K*]�9Zs��x�.���[��$�}����)�ݚP�U��-M͂��v��=��C�6����M�ܡ%/T�Z�
j��V�M�꣝N^��#IzڽG�w�O]5�o>$��y�m�|�¢��5�V�C7no���O�o+���\�`�^��uA�3&!T��|��becªҝ�Y�$z�3-��D���{�zSU����S#�Esxh��:z�NRs�,}z{��Ѯ�/�%Q��ZJ҅�j�㧟Y���(wdK�Z�㬽mՉ�M��k�x�u��]s�z.�S�D�3"�@�:��TD)��r�8J����`x���Z�T�z(��[��V[4n��WC����JH�\A��+�偂X|Ņy�cvv\״un@�K+{�Q�I�`l��2gG2�x>�E��D*�c{���A>��Q��u��%!����7<�z���-���`[��4��ηy�zfS{!�Mٛ���!id�y�)����\��K������ւ���M�|�gma�kCB�Gr�f�ti�5�ā����k��Vӳ����k)]���P�����	C&��kh�[��{����8l�N3�LJ#[b7T쾪�xl쬵�����ו8��D�J��dqn�+̙nPI{�Ӯ?���(:�Z��4�ӛ�g
�Xܲ넺j�S�#�Io��u��mM�Ȭ�
}��hp.���\l�-�gjΆ��x����h��e�q�$ӈ+���/!Nu�;Ӻ��O�	fp��i�{6�<�L� 뱱*�A�V����eV��9ƹV�4���H.yE��n�кky٘6R��Ʉ$�u%� ml����P�s:
EM8���`�r���;�?��l�oWv�vES���eG�]D��{�y���囖���O`q�n�t�����X��ۧ����׽�����G���C�������ړ��vP��/wt"6_A�S�^. Rw%B��۱;���5���Ɏwť!!�{�w.>�]�t���X�s5�Α�8rFnR�����6���g=y|\������>|�c۶��tr��=ʄc\	��
��nH�%�\�´�|��F��(�2/��ݽ3��v�^�(�V�T|�V/in��{7�-�=}; 8KJۏ]@2�qSꁄ��p�kK	)��d�UΞ�P��U�jFf��9�W�gL�ڋ�:�
yj w��g��^t�I�ͷ,8)�5�U�L:;v�`ú������O�lǂ��m�kf�	Y�KK��+���9͡.��[5�L��	����z��ź��T ;'�P�R�ԠE��i�&�=�:�q�)%�iV]�j�m���G:W[P���:6��R��6[�j��8�qp���e�|ƅ:8X�.t�ږ�{���ɮ����&��F�ئj��=ԸӉ3c����Q�֖�U9��7����3�����gn����
��N������c�#;�"`��)�L�>��5��N1�+	�5v+��r��u���׳s\���h�8��K������1�8ĺY���<��oV�&�-T�s�nQ���s�q����Y{��[�EX�vŕ˃��M5�S���c6�L���? ���Ԟf�m��'w�K��:�������h((�mH+���I��V)GY�TyyV(V0!�r��h5K��*��X	,"�!��MX�i�K���3�k���P�ۅ[�O�N�?wҬB��]<�|[�D�Ju{ړX�7z�`Q5l���vJo�� N"���l�O r�p��wW�akW!Osl��
��Ό�Gra�Vq���v�+I��:�S�v�i�j�:u!r�M*�Q����P��hq�����<N%���(�|/� ��=�9��\a����/6��I	�
�n<VٷZu�ֽ�ڈ���Q�K ����N$��� �ɧ���<��!:�G+mL��5�pP��:E��n�oH��:
;۝
v[XF����c�r�1W�W<�)ض��m��7����$��Bol�eN�:`�Ei"ttxW[ �O7��J�4�˴��5�x��:�.(,�P6i�!}(����âS��>�8�wN<WbQ�zcz��+Y�hwn��3-RYv�|����ޭV�\�wN;��mi����q�	��>}��d;5��;2��Ȥ
���a_Le^c�ꪎ_�1���;����#�r�tψ��C�^gқwS+�J���w3$���]2�m����m���P�P���s�K&���#t��Є�Վ��č���ۉVe
����7#�2�oFt�ut�'~s�����c����MI�չ�P�L��j��QT��T*��;,]��6�ZX���U�uf�h���^��S	n[��]�V��f���4i�����yn�j'Ls��y�"���x�7չ��
Q�˃�2n�A`��ɕ3Y�P��N}Y�ʤ�<�Z�V�Y�bv�{%��u:�<ј���v��'�+KOS����2=��j�id��s�w7S��\��m=9���J�������`�ΌԻ���.�,H�I��`�V���fsX�<�����WjՖx�n]�=h=4�d]fW#⭓�����}�J��SID����WJ5zN��1K�-\[x)���OY4C���m
o�ϯh՝�cB�f6�ǻlN۾�pc�aj����64�D1�:�.8�̴4*Մ��zy�#o^l5ٺ[���`���6`,Տ�}d�ﻄ��&�-&A���I,�=�ѥ
V�f�)�_�2��f�'����4ƙ�k�@LV�	�Z�rL���2m'k����8-��Gh�K��/"Pp;�k޹k��a�7u/Z������g���!�e�,�њ�"r���e�N��]V�3����H[�	�Y�P�-���iF��v��{3N���5�o��</kan��
TUZs:��Q)�g�
��Y�Jϣ�#���=�u��-l�4 d�b��mB���-��[��9l�������NU]@q��B�(넝g+6���'K
��>��)C6J,,���{w���ݗ-UIQ�HEh�Tb�tu'ۍ��,���jPz��:�=�ϱ��E�Bǚ���a9M�r�z�,ӍN ���ke�D&��pX�|�V;M�٢�XL̉�"����uұ5X�n̋�s9[ʚ��,E��V�q��&��u�Ҧ�E��in�Q�`����t�]	Ȋ��zjއ���yYQ@��ն�l�A�Qz����aTb�K�R[Bt;}��+��vj4w���)��C� �0�Zo`;0���V��&h�� �empc-�u0ʗ���sv��aS#鴨�������Y·�� �= p*�'�J>�/�R�l�f��ic�WDMuX SU�.����f��pLT�Ս��+�.�+���ܴ��B��"�V��ќ�r`�5�֞POxË���n]�,���k�����|�kugb��d�{q�(���u�yCR�S��F�� �6U�����L]�
�q�ʷX�z���M��FV� ��29��)J.����4����SM,�;��{�<��;遜�� �ǣ�epo�����S�(
�q`QG6Y�׈�׫k&�����1ԣN�����%o�V�;�h�B�G� _EMx��7�|u��Oj^��)�s{tm�!�
,xn��@���|���椘r�%,I�RH)`U��ͣ�r`�J��9�)k	��F�\�uv��C��^Ж7vt���)�gK��:���7}������֛��u\$1�=0�ޝaA���z^d��z�)��sh��9]a�㘅:`[z��Kt���)bp�ûfs�>��{F��F���d�qΈ�+j�/+�>���[�s�I}̺����D��m�Q�u/�$��mS#;e+��0��δI�2e��,P-���U�ݻ`��p��pG��� ]][�V��vE�F�k�$¶�ی9k����;(�Gv"�v^�Au���ep��4v�d9�(����h�������383a=1ӫ����B��L��GQ��K��V���u�̮|;l=b�*L�UN=��,��qM��֞{Հ�[�H�^�\f̃�X�v�Q%|���f��c�<���������EB�+�ô��8��"��
�<ܫ������(��qV��K��rђN�up�4���6����ٳ�0��aQ?�t�N����O^�D�7bg�c�97W�R���AwCݠ812h�Krim=����[�ۂ-̳�D��.�yڤM��]������pa��d��d����:��s��}8�*����+8��]A�7��r)�m�{�6�%1q־�גʚL'nӾ]Ĩ�ΒnD��;',���֗kP�C˧t�]ݢelz�>��eʉ���'e��"wA�Y�{��!���3A.s쎲`�������I��V*�]���G���V�:x۝?�|> }	�H@�_���_~��瞣�<�����-�{S��}5G�u�f6�ճ�m�R��m" ]�N+�Pw��я�ִ�d'L�A�Ấ��b2�$��&���6�[�,9Cg�x�}�.��2�Н���\:��''a�q�b�Tdi}w���*��R��s���V�N�)S��ZtxbA��Z�ʼ�2X��0L�و��r\N꩷��r�Э/� �ڕ���݉I�೯�
��i��_ئ)d��Pc��S��Ej�X������*�ѽ㫊@i=�����.�4ɫD�k�j�N�������[�=y�ٺ	,�`���x�3{U����rT�v��qm�%Mn��^�4�S�>��]u�FW �f�Sc.qP��"�fKJ�q)
G;Р�_[��A�Y|#�SVs�;���Y������]�v�k�f�P��JH����H
;o�sm�oU$]���h9/��(��˪��k�R�KҜŶ���<�`�/i�ܒ��U��|�@��{��ܕ�{�ݼq+�mj�i`|T&�<���(㋆Hųt��Ԛ��s��3z�N�v7H�A�h��R�^�o6�t�*��OFv墁�*1���{ٯ*{˻^�lb��n����� �ktv��1�;vN��Q!
���G��B�6�F��U��ژ�H!�ӽ��ʟq��d�4��ż���O�Sb�L�v�C{�A�+Wu��_P�*;̨��K�G8ӎ����Z]Af!YAv�:v�X�2ޮ�a��hHe��@c���d�-��t{x˩���ћ�9 �t�r�"��ARl��B۷Or����8���U�ʴ���y�0 mcE�v��+w&��Vʔ���V����h�����������9�Ю�fu�"��I�e޺�]�u�悙zVw!���Se���P�ZؙGi�sgQ)��hoCYڝ��aO����}T*@��
��"����ŭ�kz�K
`�1����1�+Ҷ7u�;ON�_l�V
u�f�L���lG;YRm6h!��WS��\�v2j:�3���Vq����	�E0�L��o5��07o�_f�8�c���&�:6��a9��� ���(u>�0��	�F� ����lF�p\[ğF]gQl�X#����]��t�^�Oj\8�9����~��p��:�N�v�'V�\��Ҍv���U��"�>��9���Y�e��k(��&Yu�QԠ�jN���J������R��v�=��ΧǦ����a9�:~釰p����w�Q�pT"�#�	Z�s�\!��
�9[y��41���i�
*����1n[F,�W\���1��m��+{�P�ls*тɽ��K^���\dn�/zv�t*�gl�m�T�sd�CQ�f<W��F�K&Q�or�h�w Э�e�L���Ğ�Bu���F@�a�T�򭜞Q{]!�F\!g,�*l�űұ޸�n�꒘��f���+��X���DК"f���
έ�i��j�o`����H�t6n��Y:�,�/��u��I!��:,�Q��F��wZW1D	�WcE�kj�ѻ� �8�7f�1Ug%�m��FNV��6���-h�ECH���bFNǝ�ok��� CE.S�w� 6E|�udN�Vc��
�'1a0���	��$�mV�T��随��fe(.s)�m�m��Z4�:1f=-"�s4M1�����Ճnw ���@
��g�]iGx@��z�8{��[g>sf�+��k�;Td�pb��ʳ�d��ɒ�Z��(f�t���k%H�����,��f�t�a�(��Qj��w��9H�I�S	���3OE��ʎ��[�����]QYSt���T�ٗ����3���o� *Z�n�����E`��n&7u������l�n�sdh:�Y!;�.�q��CUH��I���|Q�D��+��zaX�q��QGՒu��C:q�8��s�X�����m��j!\��|6�&�x���%&t���sCw-���5l�ڝ�sH�U���y���(iq�'4�G��1K�X0��Ή�p��veg$7d˽�㬡���W��=�Ļז�Y�G&®f�����6Jb��[��ډgCKW=E���5��Y��4*�d��[��#cYN��!�#[������	۝�l�Dw� I�Tu��ӅM��L	�_rb]��*�Em�SU1���쪺���{y7�Q�o s^,��a[u#�|�PM�̃��"��z�a�ukN��(�I��X�=[y;s&L�Zެ�`q`��T��(�6��p�ٲ��+�h]4oܫ�'�\���2���di�c��|�\������VN
��Y}�L0eVU!+yÎ��
�/F,���{�\��D��y�����-�E���F&\H�ݺZ$1Nm��]��^�oK,w q��L�ȗ���`R��G���g+�M�t�v=r�aP�w�����#n���2�hۧ��n� �P��)�ɝqg@��S�_3���Q�1
�u��v+:-�6Oj������m�zbݎ�d�ܱa���ۈ�#�,��VaXOṰ��:3�ͮ)L�����{N��8p���Nɢ�D4��[g��xo0�'�ѝ�>K�.��I=7{s~��S�Ύ�Ⲳ�Cu�Ts�^j�n��mJ��*.�9��3��)�y�ד�	q�QY4�o��t�b��q��'j��1m�*bؖ`�Br�2]$N�萁r�$7�쥝�a�{4��G�do#:u�}����&�.0���;��E����T���9Ή�y�Fq�'i�*n8a��9��z��o�&=ޮc���<���.�剜9�ka��h�=�R��}ڨ�A5���&�L�q���i��m�Ԋ��*�S9�õۡ�:�	/=��Cr�f�s��ao6�x�]�c��g���D����m��l�� M����N�x����z�o�˕0���W�ySk*�Xj�jެ�*d�n=�VaA�%���䥍f�W��E9pE�U#��N] 6�-����")aj$���ؑ������o�%q?l	�M����L���a��m�9�P�,-�Ӂ�n9k���;��4�=�Kh��^g9��hi��%���[�v,N�B�)�A������ǲ�S�"ݢ9�'4AO�=P�7�f+:�̧%�_umFw�o>o�L��,��UAP��i�)Ty*�����N�5mIX6��U(I37���k����� ��MS�GG�j�����@�+B�2�;�-�m:L�0������N��A��BP ��w[�D�/�]gq-R���6�И�yJ���\C���'�N�jiw��F��)�z�d��zv�Z�;u���ν�5Imj�"�(An`��L�/��t�s���@�b��ӌ��U_dZ�=�k�/E�:�_T�-�p#��J[t(�6*zќ��w�������#1��X��հr���:��9U����n8�K�}�MilX0��k�M�ޛ��ļ�5Y���6��#RPˇ\M���ι.����M�ȑ.eEc�v��zM �E��^flY����Dh{����j�����Ǻ��q�t-��\���#�O&ݤ&*�V����}�1^28`ً�����v\BY�ܹh��#w�ن|@VD���˳0*�v.�ޡ:��x��;�Ȩ)W1Sw|I�0�Y5���y���w�V�趕f@;�3n�ZHέKYH����{�hCXFb��e�+N����jr�&�H��2�^r�V�PZ5eǣ��A�cK�	ה�v΃��8/�}�aC�sYGsz�K*L�E�*=����g1�l��̙՝7�U}$�v�i((/i̳H�Ga>�=d�]��i3C7�qP�>��)��ۣ0\c���+5�����I4�[]��ҝj�Rn��M�W��F���������D"���NN��l*[�{��Y,h�5��V��v�f�Δm;���E���\�Ž�v��ʬM���1�P�)��w�B�N"N̉�'o����]�u6����`����d1�tg]�]��SJ&G�9[Ԝ�z�Z�����sBr��U+0�f0�����x��n���o�ҍ��	������'CQ�e�jZ��������$Fe�2v��	�6C��л�T���ș=���r�鬾Ꮀ7�R���IO���Q��vs��5�n=J���^��}��!��W\����NJ҇���:�q��`ɜj8�Ǽ3-Z�o��N�sWIN������CsK�X����UA�_\�	���2��Kb�޸(^��֖s7��b��n2 ��>�8�WԚ�DV��u\��.��'�d6�u�Lʵ&�#��������Xw<�];!f��y��j�u8(�`�YP�V3"�5β�ܑ�f�d=M�/lZi��9ŢX��8���n�ܩB��&�izӖ'���A�����^�F1Y؅:ޝ���ӄ*m�+O(x�� [� ��TΓ���ƴ� >�@U�m����-�hb�yb�j��gs�l|�o`��q�{�k_u�+�X{�q���ݺ��v9ǉaC�;�Nt4��NV+T���A���n����c�}����o{8��Z��|���u�0`�p��j�JUDh��|�{�q��z�Lc�-ɄX������L�W��4fɃ0����)��n��@�6�7�����u��M���i1O�*���׼�)���D�kN�U4�Zqt��ÃE�LV��[���%g�[�Kt\�"���D�J�sQ����</qP�z��hK�#Y��;�rΦ���at�K���_ج��f�Ƅ�rz]��&"�6���렙�.>��`�N����ea]:s��)j�����o�f��F�i�/��p��Q����[��E�P�8�]Qm��ٕ���"@��w�
#����E=�(s�;�F�� �MCj��x����)����ݡ	��[����k�B�'��6%��xcpgnt듧�D�"T���jos:q�o�l�J�o��V��Ģ����c�W�e��M�n��f�h#)������\�,:M�S�kK,m��}x�wk 6��S���s,��f_+�p\�-&a���Н��vf�\�
�Nw:٨�@�\��� !�(5�y��Pp�t\��lfܾ�0�m�Pضq�u��Vm���:NVn�/s;7�I��w`����K���م��duH5�W���o1+"0�|.��G`5\l˴��i�θTs��2��uG��ܪJB���ސ����-����8!�x��X�Z��d�N��Dd�Nމ[��U��[�[��K�q�������PV�+�#8浻�����Czn�w���՜Z�%�CB�ȝum�{Z��g��'�R��[įdE��\]u�s�Wv
J�J����b�Y 0wԖv�ń�:�y�}��ӈoƸ(Ri���Xkfǹ>�=S�}���+�]�шع�#X� AhH�gQ�{mG�TV�TUh���|���u�l��Mt�.c����B�]r�ܝ�%�\�qֶ��!]��[��]��P㵼9'�������
�A��\���s�AJۣ��r�� v���*�7q�I{�;朆K�YY��n��m�F�B���c����.M��P�ڄ��7��xv$*�Ur�S�ΰ��;��tPmb�7N)���;�cE$-�K����8|vqN�Ц��:��c�8h@f�����5�VI'[,&��j�S�&}�Xޡuv2�p���oY��+�����A��tp|m�qV���wu�d��"�����\r�i��[>�gr�����t(�Ԝ<MLq�"-[Iw#�/vsԐ����Dp�O�xT�#�&7U�\i�{I��y6�:��{H�墴+��l��:WB�Џv��¦�Rp�Sm���P��qӉ�*��ئ53b	ٌT��j����.�Hh�!9���"��Ar��;���@�[�Yh�ZlY��1��(df2���t��n�x��uw)�%��l�`ʇ3�!��A[�֦��A�vua�W.��H��c��C��[�[!���8��I������������4F�5��nb:������zP�˩�a�nK̮}|�N��5`*����p�����>��Z�qoI��n�+v�>b�Am��zӑlU^��]eV�hl8�P�ug-��u<�Yڙ��o�7���{a݆P}�,�f	b�0Cd�ǧ�őۘY�$�]��]�K�X�m��TA�.��\Rw4�ۣ/;4�7|�l�rHe�pWVfC��PU�-p����<�y`�n�C��]��]>T�s]�*��������|�OB�x�CD��'[�9N�V�}��j_d\yai�V�N>k�۹�B�mm"�]�}Y���_QN��(yJ^�Jn���[)^#��c*;;�iS�z��{Q�4(�Vt���e�]��I��-}g��	���/�uMN�v���6����9�I�n��
[��{B�;wzs�ͧFޥ�r^�++V�o���ٺL�-�tᘊum�]]{�
K~�\� �)�d�����Sfj�r�%je��ܼ�H��3�����&�L�%�$H|�R�f��k�:�(�I[2X��n�`}�w�r�T`o(��4��jg�R+j�lQ���p.�Բ��1]�5�<Q��X��X�h�A�M�׏�/r[=ʰ6�v����i��F^ق�L�8/v	9�;�^������=T����W��=%G۴��K8-5�$b��u+�a�y��g:��HCk��JDX�;.
\ч��GB���L�1���s2���>����=�g�w����;g���L�ɓ�l�Z�p�c�]�+Bw�Htrv,�9�J�o%��6����Q.�5�N3ٰv7{�{uZ�u�����E7���6�5���lv�(:��4�M7t9�M���Ȯ�;yP�Z��PȺ�����5MٔFݦ��zu�u�5�Ҕ��FD8��֮�HS�f*�fږ�9E�vd�c}u)�8��U-\�m�㵎|���ZNu�����W�#9��]�¯)�M[�>G��Yڎ��	�Ŝ��zO(�u����#��I|��ܩN�nW2ٛ�{]�9U����Kz�<X����i�ֶP,Wx��t��z���	��F�U�.0~Ǫ�Vu�wz/6uQw��{g���JD�_c�J[��kC��o�[�M�|E���S֟�&Wn\�[���9fΣ�J\�q�pe��:���=v/.�Wc�����ֆؔ9	EU&�1��.k�˾���n$�eLwvD�v�׃F�+1�W}���K%��Z�d�5�&���u��E�3hv��B�i�
4���0�/:_:,JPM�$ܼa�K΍ָ/�����'f=P܏8O�uo+~iZ�������k���ޝ���_������d����yyj>m�U:�s�Q��1�ﮙ�^ݾ�8k�1Ѽ�q�,݌���yN��t�㙝�MT�ܺ��U��w���D�oxA+���[H��[*��Ԣ)mH�YZ�m���j�+�3
�PQ�U�#1%I��-m�&a�������)J
�E��QU\�j-�hڊVT(��Q�J�[YX�TusA�u��Z#TEP��K�*�b�F�Um(�TTcZ�VA0X�V��`�ۙA�t4Z�Pkc*��V*"#5�n%�R��`��L�\Qf��F�qUE"�P�b�
��m
֩J�j�#m��jڨ��F(�(�m��q�,�#iTc[���E�e�R��ut�.j��Y�S\��1"Ŋ���2�u�T��W3Z:�9q1$��UUE�pƶ���R��R�X
5���+�)4�Uե�c��iU�.��Vک�V�**���Ƣ��PեJ*��8j�1QV��SL�
( �
��J5Z�im�,uJ�T��V-q0AETƱDPkc��9]5T�ֱ4�-EE�b �����c @� A�}�n;5�s�hN��n��FP��fWٖ�}����x�pcy#-bWNg^T&VM�r�R�-����B�v�淞CY�Z��g:���SH�@�_��/�R�f��؁�&QߪúϮ����ڸ��ڬ����p�TeX&���8qaL�ѳl�	��Q,��:(6|�ȑZ:1LL�K2����kʺ�N�E�O`��)^6��!��<�#8ߖ��x�	˒b�聇��XW�gJ�Y�[}��F��Q�u3�lTϓ�U����
�;5T3@Y���Pp������[����*��o�C
�_-��Iq�~�dR��3�MZ��9�%�7�罷t���8�s����}_.^i!@���6P��UȨ�G�S�\S��8�ӽ�-��i?������5tD&?4?,oE�
Z��Ɉ����˥��@輂��A��w��(��{�SYDU�<�y���Q��c8�*!��$�aN�X�多v��];	e.�+�ؒ�_J������hLPޖ�gr�W�F�X��j�{�c��m��!���~�ُ_���fsNv��s>!��[}��(%J�E�2i9b)�huΑ� ުO�ݮ�i����$��L1^:�B�K����3E�V`�R�To�\�^V̪��;��V8���BBVU���qî�.�#Ô\A��l�R��gs��%h�o��;aQtٛX�·j@�GڧF����#S�u�oQ{�W<�c:��Nr�������Ca�a�2jʋ����΢��)�&�D9\hHUǪuՕ�6D�`�C��LC3�b�W��R�<6 +'+(s46�(������v�/;ʻ�2��˓yd����è������koh�u�C������dlds'(O��-�9��kl�����Ҫ�=Դ��M��0�tg�uNx>�q�*�զ�`S�5q��ӵԀ�'f�������-�P�&�lC�D��Q�2�p�f��Zn�F2���;%_�Q��c���kk�.{��;��V���ιP�����tۜ�Y�q�)�p�=$�3��*�!�V�F�Ťk��!XԒ�1��+����L�9��Jy[
:�v��$���<*�"���JJ̡���=Ez��d�G��B��Q�A�&n0έw'm���m����qQ��K����:J��KT8Y��m��x�.,T�g<3ru\�_k��`b ��ա�>����qd�K��D�8 9����6(�r��D�u�"a���-"uO���=c�f�P��c3�h<&d%��{K�>G�Y�2�z�T��k8�-\]2�:��i���&��ޒU��Q���W7ٽm2��5�{.�Q5�Vc�Q��Em�њ5~u��*w��ÔUO99^�Z��ۓ3a�9VT̞��.rӀ';�:�K�"�J�x�}��#C�!BOM������n��6ok����Y�a�t� !��,��m;v4�6��8(LR3,����W��M7/u���.�^���Pͣ
�H�f99�Z�	�(]���d�<�I2����}�֘����}��ѯ@P��c�>�F
�v�+���U��S���~�v��Gs�g���\�D}sLt=�y�5Ȱ��A��8.�+�q�Y�5γ= ���}��&L�J�KNUVD*chtD�����Z�	�n<zz(K���"�\g�bV����Y�1TQ���a�/|a�b��N*��!�7 �nh��V8]�Ҕ���c��9���<�@"��w�4�����<��L�z�����e�����(FP_��Z�)ɝ��r!b�<��I�b���K���T��qP�꽌��v'NW
u�NE���;Z��!&�q�.��d;�P�!�J��d�1	̅%��t�.ob����^�c}�#���/�Y�^�Q��cL��a@F�^���u+f��=8�����e�9��M��iK��Kk��GgJ��kW9ݩ]+v0{�T�s6������gl���D}%�}���4����CI�2㶀�]\�#�W�bg���eǻo�XDW�|���U�Yj#H��J'��U0�A.��9*�c���OUP��z}�}�4]q�������RMseH���
��{<&: �t��$��Va����Yohi4�<eV���9�RS���(q���ї��pey�J7��)Y'0�V�EF9N�f{��=�K���K���{ڎ)����;�tۈY>9��6��K3'!~�������Ƞy+P�I�v7<���.�/n����tu�]��N[�X��0j��#�D��)�M���Ak�����W<�pFFPN�ǫ�δ�2��e�\���.�U�f�Ζ���D�FA;&zV�b�	к�B����']��c�0`\߳ݫ}YJ�g��$@��n�T���jV���W�,mv���h�q�
�\ۢ��0���/;�c��g���n\D4��k3W:���z�f�mlnT�v#6::���yS��d1��j�UG{eto���D>�1���0'��}���1��0�r0�>��1�d�������3
�ŷ���&���:�IU,����W���w*!{�f!�r�um`�Y���1�����6�D�D�����u��O4gy�������[���^���̾� íef�(ή��q1�N�#ob̋�&�֧��;mF4(%�}��U1F��@�!���:6ͣVZ"$4�aG7��!��ul���̚;`��h-b%�BK��X�7,e({3УUU�zC�/�å�GA�wy27�%U;y5a���f����{]�Uٮt�xe3�$X�.������/��X�lwf[��+�<���oo�9̻~ov����}\C8�+U��؀�j ={��@y\�2����N,Wvm%�G�UdnI5���%��y/ME�Je���C�ހ�w�S�W����շ���������"�2R᲼�n�z��'/�D��`�)���L�#کΏ���;i8�
C���n((�*�ҥ������J��
Fq�-���'.I�����Rd*�i=姩����.ʋ2��L����t���n/PU�٪�������p
KNi�������CU6�N\v�/�H2gʄPd��"b��F�ϖ�k���s}�m���<��w�Ͳ�	��J���;�h<�!+2#���"��3t��E޾�e�e7�GWz�����}/�wV��l����3s
�$s�z��P�BңQ��"�6�+�M�8V��#�73Q��H�"+D��4˚���V+��]���`b+w'IS�R�W;G9%X��mk]��^g8Xnt���bW�����휍>zܗ�����*����b�����߀�1$�Ź�LG�&�&yt����k���'���{�Sc������~{c�d�%�C��ߡ���pyNTC�q2|��'��j�-�R�QFy�9خMO#��'�����"cx�J,�b(6��|�X���m��W�ʰ��0g��ZPܡp����=+��q����*Vj/��I�^i��"�hu��)�#烫�秪xe�i�uG�B���WfS>��+ui��f�M�@R�_j������h� ]����r�ߓ�US
G_�6��{"bNݎ���U}�w�^�r3�%�V ��r#�+���οP���\�	·=;; ��ʟ!$���n�!^�FVьN��Ìg<�S��EG<�ɑ`'8ڈ�C�F��J�Z���/���)aٮ��8 = ߄�G:��1��i���X{֧d��./i��v����j���\{�ߚ�<#�md�H�V"�H\�M�tۗ.n�q�
VD*Z�ͻ� 
S*�M�>7��Z�L�̶���&.с�ꯐ`�\:��VAbZ��5J�Y!�,N�����SSlw���0D��j���d=z��r�8�j��ٲ�w�8s	�=ϻ��w� 77�P�ArR���{D����\�H:놝�I�ڬ�ޜQo5��!Z$��S�t���6y�Wb4��r4�R�y\�>�3Όkwڹ���xh�Zyy\kh4�Ģ�.��dytx�P�c:�:�w�0�}��1Grj!F���n{m��-) L�%��Y���e��x�6��@+�-��3��s�2�^Ӛ�;���+��R6�N��Ɉ�� c�A��I�E��z8��vpލuk����3g QN��� =8���n�ؗ�p,#qQ��b���=����G=�MȺi]B4<���O�
r�����N�,�9�3H�Nݍ�sX�fĉ���.��Lm*�}����(�L��q'�\�
��0�t�fc��%�@c���I��#6k�����T�nj	���Eə!h���["c$�r��+��D6;����%ZT��'994�F���S�obޠc����]M�S`����@��vc<+�㮳��?v��zZ�~i�S3x�p���W���+�(�2����#5�=p�!�z:_V������T텶�J��0{Y0����6����-Pɐ�C�vNNlԀ(���ok�ֆ&��+�s�ͮ�n�Ϭex7����W�A:4�\5�Զ��_:��7Vf�o�u�QO��ȕ#S/�j�}.�f\����_;{A0fR�ᱨ�u�RM�����P�Xwݲ�ڧ~s�ژ(��g���@k�jǭ��4fvͣ��=l.ܙX�:�N� [A_T��0�s���E�up�&59�;��>�gG�v{���$L���xV��(�x�����X*b^�Uko��*���V<��`�j4���FkBf��&�:Y�3Z�W���R��:�뮈�Ds#��l�96��c��b�h\��F��cG���m�tE/�
zYX�̯j�j%���y��d���=��fNzosrchQqV�h�rۚ/�G���F�T1|B�F{���2���NT�pN.Y�I�;q�Xr**ڢ��hk�90y�)zF}�4��!IK��h��x�y{��ybd�#{���棤�W����ś�BZ������O�ķ�L�~f��T���',�5�6���'M5������g�ym���at��'��N��r���]��%����P���:�B���,wI���-�mmB#���{kڴ����yF���hH�-����b��RE5�66��W�&rǴ����������5R���@�T"�}- �z�c�5������'�k��l���c�G��U�����۟�g[~�~!Ṙ���a�2�v�������S�=�m0�U����h��ᬘ���L>}��<l'7%�"�N���i@��p���8���P�%�iwK�1
���$@��n�*W%<֢��@!�ؼ���X�,��e�����irE��0O�wF�8L����E4�d80l�s�9�>>;��`��������`�_���&}��7�XF��ݮj�B�ޒ�S���� ��Rw*���R�{Tr�S8�ޠ��+_l���:޽�u[��c��t^�F�Ţ"@iX�0����'כӗ�Zb��p��Q?D����J���*{j�Z����C�/LªP�T���u{Թ�HK�����V�a��1�=��b��sq�3�wćg�Yz\l�W"�i�R��<��Ǚ�-�UF}��_�6=������F�!�@Ȉ�ND�(C�Aor:�d�v�����1Us��UN2fhInz�%\�>V<�\���t�{N�Ԟ������9T�Sj��i�P:�*�Jp���n��Vq���N\L�7]���5�FG����]�Y�H ���w����N��Ȋ��T�Y���i+`�,�o^���ai�84��eX掁[��'8~j�8�w��H P��:��ݬ
dF�3�u\e�7k�dڛf�Ɨ'��r��;Q��� 7Ҹ��ƃ:H���.����7�!Z��,�F���%������
J��҂�:O��N�.k�Z����H��4�D��)���/�
�f��]�UC4���U�uc��0ݮT�AwW��E��I!	�$��H�]WpVE-��� �SV�R�P��jurkȩ�z#�%n&.N�q~N|Y��D%G�[B��вU���r{H�7O���j�f��q�p��><,Xuޞ�E���@�'^-�DG`��$�].:C��Zj[q���Q��Č��.6
�ļ�b!�_����+`y��H����Nt푾+��p�jf7���5������nИ�)�� �b)�he�$dEs��G{m�9.��1z���=ө$���`�3ۓ����̕z�a�	R�Q�����M#@����j9���N%�E0�9����جQ��
���n����T.�^(p�fqbw��[�:N�c�e�@����;�DPm�7δ̬(a`��Qb`��7C��n�$|3нp�܄W{:��^�	֫�N�g�DJE��;\��['e�����;T��Y}]K����ҪQ�aHw���5���^^{�yi��a��R�՝�Y@��a�cWfdf�ޢ*�sK�^-h�8�в�^�`��s���p��J��� �ol<�z����U�iܱ�ʙ�1�]Z�y�����T+E�P���z_�f�t�S�ea�&��D��!�wB9e�Ǝ�Q��L\�.gn]�L�÷���Q��%��pd ��(M�7������ �p�KgY�Q��j]Z�Z�+z��5kU]�\�r��Ja�˧&��i�IJWBY��>���ź�8��(�4ج�$��hm�s3�։=���Ge���F����]�tԊ��:���$]
`�ɘ-�|��e��P��hP[�[�5�n�v�E��SI�+G.�/j�����Pk�曌Wt�YR���Ѡ�,���ɘ��9����o!P�\��}A`[��@+�����nI�;6^�DڃZ�ۼ�e�;��̣{�1�|��G(d�4��]��x�%�=�{����[I�E:���J�����]�>��ƈy{���.� ��aW;"�OF�]X��&\���2N�=ɢvk���\0�k��EV�|����²�86���=��=%
i�v`η���N������=/#�p֛��/.�w���]� ݝ�__@-V+yA�1�J
0{���6�����t��Y��nn򎮧M�WT���Ɖ�� ��0ԡ|8NF���]����ՙ��gAmk�3�]b�V�h� -D�i{��5�1W^�h<1�`7]rt�+����=��'5�)���T�j]�9>V���]��&��dmM�a��Z�#�{�ۻ
��S���K���5����q���uի�np{Susaw�՘��'2c�<u��Vo0���v����y����i����Kc�=���J�)�=ف�8ɿeq�L���v�
�L�};�лOGl���w+)��R*�B���O�.�Z��b���X��킎�&6C�[`���Qћ�[���\����QX�2��UwK F��Okդ��ٔ6;�j��c:K��.�(��mE��R���ܛ���`�V�Ȉ%��j'�]�,�S����W9�^V#^}�q����{EG��j�r���e7]7mF2�2͛��&�A��c��-%����u�V.��Ǽ��M�Y�p��1WL|���ERk�Ȗ��9���M##Ս�m�\gw�&����1�;B�]�j����:�+�,��wsx�9�Y˙z�DZ�f-Z;4���b7�մ�,L�f�Ͷ�S�FLgD�e�:A�_L��\9
7��g�����G��B�.�7/�u>�w:Lp�;j޾hXK�,<�}��5��V�"Jy��k����
iJ�V�P���UQ�֢�,++"�U
��b����,ejZR�|��P�̕����DF���#��V��M!R �J��DjT+*EĬ5b"Ƶ��U"ZU�J��F ���*��X

�l-ƨ�(,Qm%VYDU�am"Ŋ���l�KJ�QVm��e�AQ�,��Z���F
AQ-��V,TU+F� �\�qE�c�-m�,QjUKed����R*��lL�*[-�
�(���L�T*�Yb1����1D��"� �KeJ��Z�b�d�Z�,���#@��Qt��bQFV�Y��Q�ʈ�YDU`�H�#�-B�
�V%�H�6�EXV-(��+����$�Ub"�E�VTTbꁉ�k"�P2�A��UAE*��e�*�ł���UE���ֿy�ΰ�N]�X����|\*�j����Z�u���<2C�K�Ω/=:�݆oS����n�P�g<�5K���9��|�?|��y~�o�߼����K��0N?��.�,��`t�����r���xj�����R�C��g�p�H�瓙2,';���1�OBNY"l(5�{���r�����,D����z�I�C��q֛��c�5�=jvJ��%ґ�wa�݈+W2se����b�O��+]!s�*��(:u�.����¨�Kf��n�RW6�(|�r%�U6U�x:I{L�S�Ɂ��3���f��l�SI���"�-k��0e�t=��O���dq�^��CA��X�-P�%�&��<o�(Y���#Ȏé����wM�R���e���(�9��'IW�Tdp�7�C���2�q��n"7ϷV�v�'�zቼ�q~�-���b4յ@�y��F�q:K�=�P0��2�����7��ޝי�ܪ$��x?S"��R���s�o�b_]����AF�q1�� Ň�݄�f�kmn��N��hB�xL$9;P�����.mNݍ,Ͳ��k���(E��i�wv��ٛ�Y^
�b��w�P�v��9���Ldw57�=3-c�˳AR,���j�p��R���<F��״18�}��IT��v�pb��/〡�}�J�x҇fЃ���NR��h"�e9Ū��cz�1m;/�sow��2��G8"_�\B?s���!���e����Ĵ!�xN6�.�v��U�ќ����[�&���|)Qg;n�D�a��?P�ۣ(��Y���Ώz���oD%z�^���D}�����5>\���]�;��*B��*l�uq\5n�1�p���o]D:�ADA�����"��3�!�CGO@��hdv���r/�.^nԺ���4U�vIZ{K�8�s�ڛ�s]74\���3{��wZORQ�nvr���Iqd��doh+�T��2:��8�i���@zs���^s����V�{n�Iѽ ۉ����i�r���ʈ��6��Hު��tC�����'<�6k��o��8�\��B����^��	j��vE��O��h:艱%da9��ֹ̉�۵�Iꮜ)��,h�'��Q��V:����j0�����vy�ح�CUP��3 ���O_�.���"�����Ӊ4B���j��km�p�t��7-�}��6����(����}�]o*g�37wx�if��Q��((�����M�5��
Ѽ%��y���}�e�g6ӌ�������՘66{��k���56�s�oU��m�ybp��]�2�M��]Jp�̹�\�#)�N�IdǾ#�={zgh�Y�Ag��VUlbrZ����g�(������V,ˣzlLղL�sQQ�*qz�(�,k��"�u����}!�u���u\�^䶤�gxC��{v��0wL�g{�ڷY%ji8���ΰ:�^F
y���m��}k5���}��Q`��z�D�$�1 �ʛ�t��ǣ ++�k�X:����;��\kλq�f��6*Q��ܖ�*	iF����P"z�����4x�)}�m5d1Nj�z�A�>d�=�¸���i�ܮ�cX�~SU�ה+��:���C]t]�~�7wF�t6LSr�"��5����9ל��z�����+UF�_q�ؾ���L�џ����Ub�������<��K��^�jȇ��Іn��W7=���^0����>Z�.S��:��w�^�X�b����-
��z:�Qж{Z兦��K(��dNa�}g¢��o��7���mՉU����'o�˙�p����Uˆ���s�o {r��Pte*����;R]���*\�����uӼg+3hU�#�[�*֍��z�nϝ�
��ܻM��ldP�-�u|�ѻ�ns�n�Af�-^r����j��k�Ad|2gq�6!��js��If6^�^���ŋΈ���诟^�<3h�g��7��F�����������G��ߚ��y�_'�y��X,h�S���qN��U��ߚ/�VGk�#Iڇ:*�'Es�6L�j��u�1/nئ'm���:�qUS����$��σ���ܦj.Je�5\EU!���mߔ-�����>UjR�e[r������9���\ kK���=��D��J�"El)^�c��
��H�qX�Q)�a�_e(�)����m+O�Y���hVu<N����|#K��~�cj<40ꔩ���;,���"����/R�������X�=���M��(0>]���|����_���'Q��W|�)'�g.��Oܪ#m�q1ޓ�TZs���D%��J�Q�P�z������ܵ���3�G-��^��q�o��!�FE'n�/����A�s���6�c�F�l����nvY�=����q�#�',R��y��,ֆ�c9�9Q����W���葂�M=��w:��{N::0�1L�g5#�^����Rx��F;nľ��٫� �2�fl����mΓH�j �L��>庙u��I�4s��=P�֩���^%�*���u�5m�t�^��Iӏ����gnw%�nP�O�3�,�'o�ᕍK�A���o�����qȰ�[67���۴&+zS%�e��ѡ�rFDEU����fxt���Ͼ��� ~·'�%��y��lk����5)�&��#���鋈��)�M�h�腗zP,�s�E��'ܮ�&CӘn�����ZC4u���cA�u�:�<mg��^B�9UJ M��e���i�7δ�L���p-����LI۱�Y�H}ٴ�ٹ��ީF��ea�}���g������|����f�^X�Z���5�T\��w����ol�_���<d(�q�q��2�}B��s&Bg"Pc��Z P�6!0E����N��>�tUԀ�װ�H3:�Q��4�q���~M�ȼr�֛�́nr�9x�Iƹ����
���3�q�>���ޔ8��D�m�:u�3m��6$�u�=(��4�>�\)a^<�ʡʦ�����(�%�ژ�<Ϩ�iDܘ�Ǜh7�{#�ݞX�Xȼ��1��/L,�dtRr��^9��2P��	T��9G%j��_KN��q���e��:�اK#b�P��uXb:&��e�n�u��U5�:�}��^Ԓ�h*u��o���Ln8�e�ݖ�
�_k�8�ގ�����3;S���ғ��7R��L���U'8��^�_ s����$��M$�J��6>Θy"��L3�{�Wnx��5�B�pT8:�R#���/њeb��N�����2�����qcz[=���i�j��gb���t��LD���z��g+�E����3	��7x�]�S��NwM�blK�
*"
/;3p�y3=�{5�G���d�4HD6�%�iϬ.�xLv�$�B�r:�.mNݍ��|���y���oa�b�t���"
�cݕ7�B�C6�*��������l1{]���f��1S����B��<�F��w<���h�@P��c�=��,"7^".�����3O�Q���E]Xj�¡-ˈ����r�X�]V
��z0o����Z�xM��dFe"�V�M�l����Ak��}��_�SWO�"��p��u���zx�]���p�<�y�T�RF�ʆU�VzK��X��=�qL�Do�U��t ܮ�9�Wݛ�I�jSDDk��?����k���Q��u�Z}����.g<�i�o]\u�]�i��b9Ed]R��Q�.��O/ �n����[%��D�^+w���������������t���^���$o��쩬���VM�ruoGU�8}��":�5r0w��ɜo����'"�&�4�ݭ�'�����qd�L�]@����<�Έ���ӼD��JvN����s�(���vb�Z���r�Y������K���^9��p������χ�b�%�����:\���|��@�غ{{w}쬿j��%�(�pO{t�4:r�.�v⡒�"�"�Z��3�U�Yj#�f�[c�O����1�>��M�o��W����g�'-������_O?_�p�T&�<[�S��=�Ms�IW��Z����w�\TP�TQam�y4�<�*���i���
J9~����/�o������`0 r�*e�q�)[��΃��\�	�u�����W+.{�������5'$W��t+@T�=��{��7�������n7Cc*���UX�.��¬��~�ӻ�1}�׌�#B����@����[mA��ޛ�%�}d��zGoT"G��5�.-�7v��\�"�ةF�sr[ȑ���*Z�GF��L��z=,�ڞ���js�3F�a�]�7�]��7^Ŀ5���W}D��v�l/^��[
����}��3��u��^�B�j�hklX�%�<�C�5p��^��/�g��x~�=8_s����:LG�1�aǍ�g0b�W僎�׋I�[�]��6GbI/t]f�OZ}%��(�*����%=��Ӱ��ڂ�_2i����������~����u���;�^�����_�0�q�#Y�8b�:�3��Fq��Q�ǜpl��L~��͹�-z�'dk��6Dn�2�}�PZ�||��K��T�)����Kb���uwݺ	��i��9�s���^ګ�CzC�,v�N���F���Up6���e�]� |�G�K�h.`�i׈�Q@n�ZX8usn�_N�����߼߄��+%>Tz��2=�7�w�#����]���xc;�C���G1����bا�Y��6r�W3���� N��|������
F��!�@Ȳz���Oy�L`�ip�k�jz�ӫ�=;�s8U8pɘ˲��%[Gr�h\g�yX�ٺ�F^�]��f{���H�>���hg*�pwܩ�g���=Y�r��d0�"bs����7�
MބB�z�%�ҩ�+C���c�_;�(�qO�`(M*ё%��=53�]MS��`����xF�qD������ᡇW��-Ruܚc�&hf*+M�Uy���.���%�րy|�jӘLm��YH̷�ۦN�x�$g6��ҡ'�k<�4w��A+mp�Տ|�	>�f��tC����*�;2ЌS��o�d#�μ0�m�2�����7sD�ӈW��cgw�{�)[K�1Y8'!����A���[��<l-�!+B@Հ��3斎!X�mY'�[Y���d'ݙ4���궄a��ݽ��>��v�:�|��ΐ2b�y��<C�ȝ�;jް��Ӹ+b�$Tr��F��^��������@T�x�� l�H��Ӕ����aj�T��Ξ�:6�$:����R����b!��V3�r��x�t�=���U<`�U�w1�#�ӱ52��X%3{�`H��7�2Y�\�F�=�cOm�	�׻=ͥ�,��Ǚ�y����ҷ'��xrʌ�5�ÿ%J�E�2EU����f:^.͔��蓢��@�ob�BW+F��=�i�fC��Y���k���
>+��~1�|��{ʝ�v��o*�A�yM&�DW��9bo�i�W�#���к�<�&$�����K�x��9���1	��ԇꧧ'Q�������[{��	�s�Q�vvR3)sB
�I�ܛ����N\��6���'����ÌguN�.����¨������ⱚ�e�$�]���*F�sgz�]̪�Z!JջjMG��7���T��.ՠQ��j�͝7wgD�@�f��gu�%�f�tvћR��y.�����|���V	��K��^:vE%��2C.ª�F�&N���*����;������m��H{���#/F�ܦ��M��t;�ޣ��i��q�n�Ft� �4��+cyC��II����Ո���:�gJ��G��L@�>x/����9a]6�T�+�@�ڇ�D�3�P�x�yxR�>|��*�B�:I{J�v�XХ��s'j_��^���7&2�^�М��__◦�����HD8�X�P��W����|t����|��.i�>��lg�����N\a�Wnx��iC�Ↄu����4�ީ�����#I�@٫mp>�L^j�ܪ�b4ж��3�H�q:K{&"�WZf�H�qc-�u�ث\[�9t��M��
 �]�
����NwM���}��P{]o;RsF��SR` ��q�w��ش�ڬc�z�=�u������g�$�̿M�=|os;,o��ߐc�Ŋ6"�����&e�y����aWH�f��7G,K�Y��&�a8�	�}.ۚ�B���R�R
,�t(ϩO'�a���oL�:�B�
��ڞ��hX4ku*�����6Q7�t���\O����?bt}�}	��<��Z4,a���($�v���2x�S4�#K/�

����L�z�S�h���ܗ]��q`D�C�S���p�Z���f�ƹ������t�	+�
�(b��Cү�A�9�����盛�dҜ�pS�u��hbv�'VsW�t�u؍d��	�u�4�J���ZY�0���mo|��@���JCv�>�m���lmC�]e�P�.��U�|����)���Ѝ�:�U��U]�/{�4t�M���s�Y�T�ٝjl��ᇎ�J����z�{���,A�f�����Ѥ�]2E�jpz�����墻w�Y���t#J]z�O���꛻����_B�Ҧy����Ui4t&`�5'͍}h���5\�~IQ���0+$e�@�e��7��Xخ-	\�m�j��3�"'e�-\י�\42�,BUv��
���Z+��v1�7�D3)����ږ��4�6���SಋB��A0:c|���S_4���nv8%Τ�j��4���\t
�Q�k@ǣ�J���� ��z��Q�SX�e���d���90����w:�Ւ��l�]׌�®:���9t��:�e|���o�m��-�����EA���S�w�qh[�Ԯ�q�øe��c^��㔔�m�F�ǝҋ�N���c[H��a̜�R��w����u�Wj�WRfS�]pPk݌ɽ�����헑F��J`R�k�V2�'�ם�s�o@h+ܸ�s�������Pǯ+9��Q�����ꗯ_9]�
3��B��ۡϹm���#K0���Բ�
��%q]V�2�e�q'_l�4�L���<��kٓ[im2�w�E�	���H�޴_J�2���Wj�'};��-�|��+%�L�kl^���E��o8���R�\�]o5�s4��[�r�d�L��t�/�ӥ���.���rZ��0��>���W��-5�"�t�CEZ!y�����CM�q����9��	hSy��Z.�`�1;#:��a��+��Hg ���ִ������'��j�+�ŨWe÷�6�B�XmrH(*��
�S!�pV�\��m9C��m#�Oe����y|��ۊ���{�>�ǘW �|�uRbѫ75��)�x��d�})<��ׂ�W��J0E9��#��vԝ��=�|��DY,���ϥ�D\ ���9/�m]��wQ���@'�[��R
��ި�������u��/^����1�z�XԻ9G���G������*����&�ĩ�h�s.����Q(�xur�)��UM�ۀ��N��Zʔ�$�h�}��٠�N[�� 2�V9�hK����4_�����~�����ɻH�m�,X��YT�AH��*�%�#Z�%�m�J[D�
�L�F[AE��4������֍���,U�R�e�(�B�1��,(Ԫ�*ŎRQb*�����t���dE�(��AJ�����Tb�@Z�E�ԅQ"��Ym����D�*�Q�rʂ����UFآ2����)+*����B���,+b�DQ]!X�L�*�Z��
1DDX� ����mQEej,UV� �X4�U�QU�4V
F*�Pժi
+"�*��@�����
�E1*��B(�1���,)*��Ȗʢ*��SV� �ZՊ��1�h�" �"�3��2��	�UR
�%b�H�Ѣ*��+q�U-`��3T���aTFj�*"�J�+U+
 �i[V�Z���ikE[K��dŶ��
�JԪ�D�R֭���A|R��?�$��7����Ś�jFj#��;�Ӊ�H<�l��:VٮGV���s���|�ż�:�Ԭ�Jo]��(�PD�r��x{�xx��oiܜ͸
/vj���T2f��ԃ���Bo�y��@}��z uH�9ޱ+�*�l�c��8k�c.��q6F��f�0<�p ��� ~�Fy�d����h���η��U�C�۝탊z1��p229�U�VzK�c�X���ڧ�DC}7 �v�[&��*ش��R��@yеa�W����V*�S�릵KH��s��M2'f3ֽ�ž��6ī���b5�&,';'nP8�[�P<1��;1p
�`��{9Q�W�"9DDӘ���}�����9�Т᯹��Gk��p�\�*����~lS\����7oB�zx��"����ٜ��wꤲ�!�l����q�豉u�vTy@�6���Q���7ʫ"cjՁ�J#Y�FxTY��'{e�
�Kd�ϡϹm�ǆ#ҧ��/�Uh��>�5;{~�:f+F�̬҂��;
���0��̢&��,���U�,�9��Nv^��U�S���&�QADnEz���`ֻ�����^���
~�t���{ʶ��Y�$L���1n>�>�B�u�*}��Ì$���V)�#3r�t��\��	��T���U�5��۴wu��Z�Fe�}&�R��{��f}��`o8h���7���-���yR?�Gx����NK�oh|-ڛY���"�o�xx�6�ﺓ�.��u�l�_���t��a��|X�x�;v��n���aĞ������+�T�c:\N�푉�f��H��Du�)�l-�Bsu�����iw��Z��o�xj��h�3�I \^�;��i��l]E�Ք�����Q�Ꚅn�vtŢb�/ChgN�в�I��(���&�b��Pp,)�u=&bR��q�����Zc��q��_p~j�[��?�B�:���4w��^ ?wc������(%ӱ� �J��Me���s�V6��붫rx;-e+�@�s~����P�F��$4�"����u&�\stW
sW�<a���BwA�Fפ;�"Q�w�J���Wx��h�b����+�q[5s��AE�G�@���4��"$7Ҭ���YC���A]��Y�������ڮ����\�i���<��������l��_�O:�Æ�j���P����\�o
�Fh���b��ah>�Y���W��h�*g�ફ���N���w���ۻ�v �z}\C$�|�8�ciS�@�,�'�^ӯ_e���Hx��.�@/�n�x��lw.�ok��8�<�MC� ���eZ�a����ݕ]qC��Wkv�u"�q�	ꢍթN%���s�-޲�k3��M���7ja`��*#X�E�g��p= �l0�`��?}��UW�H�-֚��W��Q��h1!�A�u�����c�VF��5��i��zj+�-v7gr��C�y����>��
t�oB�k3^�T"�q����n�"�|��=�|K�
��m�=V��DÁ�Pd��s������S�Do����&u�K��W�x^ys!�-�.��p�b/I�ЙRL?� ޞ��cK��_m�\��h�����T�\�w-39��B�0�z:7���rɴ��	��/T��q�T٦v����Uj��S'�f �������vո�1�Tjs�� �H����|{���M��������qŵ��-;��a�]3�0�>^,��́=�ʋ��n0E�@R��4wL�8�Ԯ/�������N��+«���e8���	�!��T�/=F#~�D\SuX�	�d��[��K!bb��r#(��>�b'�1ӱ53�r,<���04v�	�ޔ�gr����T�D����+�f���J�{�c����< �0vZ��r��Wk�J�<5ݼF�[���]H蜵���\�uq��Q�}��x&�[�޴�)�!ʖw\������2]����{O�)�|&Sjm($ӛ�&2�1.�L* y��BgH���eNr�����pU��1]�փ�s�^���%��ޔm$L��=�
���%�5M����������5� ՜��"~��(6�MuΑ� �q���C�n��V�כ�Y��3gv'C�뾌|� M��4�`��<��z��0���B�Ji���J)�𶖝���A�mHqC��ON_TB�K��o��O9�o�<v8z�tx�Gv9����8ʺ���
(	-��>b-셓�AGA��'T�c��s&F�*��=C�ڧ���VE�"xb��m�j��]���a��zj8:��1����O6p�W�ݕ���9�X=z���m߁�#�V�y��9���t�y	ޡNT���KSo�u��ꭜR�ԫ X��8�r�N�EIB!z"��z�&m�.X�Y�3\�uRMDʾ2|��q6�$h*��Y�e酝,�6'�Ԑ�p/��X�-P�ŝ	��B���G���!��].!E��<�c�'֧.0��v��Ԧ �K
��AnZ�q�M��'����n��W�|��^����u��]�ݣ���mH1���F�q:K�}銽���t�m�8-XF�~&��F*&F(h�*Y�r�m�|�F��s��c��B��|����+w{�Mn5�ؼM�)	 �r�~�<����杉�}:��zv�%��u���^U�E�#�N�e�8T-�zCYMhe���O�;B� �F�퓴�� xz�wn���UXb W�3$Ez�7�1�lc��	Oq�T��<��~�n�ިW`�~*��-��8T l�w�
�д�-8,.�`c�zǧ���#Ƙw�[0b\�ʹ��5zX޷cr\�y=LX�EE0'h�B?s������;~�\Ah��;�����V��,�?^*D�� O��P��k �U����5��g�����7��,+v��ӹ�1��:)�UѾ.2������刿s�u6��-	�턞o]�v�f�}N�}ʰ�Mlv�(�W��,6M��u���ڪ!ՇADAMTF>�l�\�3m^��'OV�|�3��*SPL>��puK��e�PU�g|]U��=%��b�{T�舱��U�s������B��
�>@�e�+��w�րlU/���L�}3��ԯI�8c���\��3,M��Nv�>��~�cG'�����,��xeS��vb����Bo@qЫ��1�5��^;��mU.S�\5~|�c�؝7�Q��*�:Gh�U�*b�qQ52��0�s�V��TI�IZOj�k�)i�;쳸�#o4��:��ۜ6�6|�h�6��a�̓y2����3���+�[4�����5	|������d�(�ox=���J�H7L�G�$�E��49�nk�����}�Wnw����z&k��N�\G��zb(7#�K����xw��N�=r�#L"�_�V�A��;h��s�^�v��Uvs��\��gK&�e��	8	]�C�	]�ш��*źq&�"���ksw���CX�Y�2�{�¸���0��̢&��,�M+U�1�q���u�V�&r�1�z�3� ��"JES=�s�n:�)[��΃���%	���l�fʅ���r땉`o;�p>��c��2gʸ�MD�ɟ�-����˗vuxF������1D�s)_��p[v���
�l=� :�� �1㲠T�;4���b�8�yZ�:��c���j*0��e�22��q�.m�aM��S5%�Dq@�������L�ҫs��f��r!�#������a@�N����D��7TS6�o�SW�؍��nD#��c�������D�;�g�ˡwC�0�hK���C��G�r�"�F�/��0�؍¥절�m�oׇz��>�Չ�x���ǃl�w�$dP�p�wF�etn1���*V��4��UK�ٗe^��G�.3��ʲ�ݥ}�8�B�2�M���Sw<��z��4ι��B�)7����ǡ��̽��ns't�W��P���gYa'�lQDy��6�rwO1��s���
0�ZmtB�7y�[����6g;��q.�b7:T p���j�?|1�<r�T�_��j�Ot�8+�P���廅t���Z���E�f���+,k�2EC��`R�x����>�6_r���Y-���ҍ,*� �ȸm�z��t�Ճ"�{�o�����]��ҳ��+�XN�^'�����RM$X�z����r8����'~h��Y����R4��C���w[׃!c��;X�������q(ר����H¢"{�s8��ÆL�����9/mm�f�������c���]�Qym2�U��������X�T᳁��n2b�dg*ȉ�~�5�>sfټ;��U?/��'_�k1=��+��1"�Iǎ��,�������i���<a��i���e��s��Ksz��٧��0g����<H,��u����s�ӌ=C��Ow ��C�2�>J¦����L@�_7���y��4��R/ݡ��6��|�������.>�6`��k(����!Y�%|�ȧڲ~e'g��6���$ߙ���0*��klu*A|�V�l1�&!�=�i�E*N>f�Ċh-�ԕ�Jì�6}�j���
�g��uT��9+=;���=B�%C��m
�u���z�AH������'��>�r@�_Y6y�h������I�ǌ
�Nw4�1�bM������q��ˤ� 
&/B��"��'b�,�*�;��ͩ��xU�g�{��(���4,~�����S^!͑d᭛��[��ܢ�����e�ͨ���V��	�L%m�����n�b�h��t����2h�>�f5���QŒ;Σ}��.�΃K��z��Q=uV{��gts~��?��6�ZŇAO���ɪ� |��OXx~�
O���}�Rx���1��>3�����%g�����s�� i+<5ߵ'�^�*Mr��=�=��d/���������� �S|���2�W�P��i �a�c�O�Hu�<�k���T�򟐩���;~ɶ,��/,Ǭ>C������Èba��LD 2�N(x>7}x�Of'�}�fs[��z�}d��u�FЩ+���&����S�l�AH��jZq5�!Y�5M |���+�,I�u�>��!�>��]0Y������LxLy��>��U��c�ي��=�~���:�ƺ��vs�h�m ��y�֦ ���7>��'�VwvLO>�i��B�J��I�*�>�~t������u�����$�����u6���:ϯ��g|���z򶦩BF���i4g���2=�1q�|{�M$FN8���{��:��'y���Aq��6�_�bAk��d�����a���������,�Ri*A�޳Ԙ�a�g��c�~I�Y[�}ګ�=3ta���Zw��;��6  Ƕ<?&jͲb�~�d�����>��6�����CH)�M>�;�~H,����sRg�x�]3��p�}a���g�2/�
�ϑj����S��D����L��jCsv~�#�Q�c����c1�����A~a�3�i1"�Ĭ���0�����~>�O�m
���Y?>�ěB��]l�ځ��;߲&�HVi��wh3,��Fwھ����+繮9����*<�1���e�P���凎0Y�VOƬ�|é�1��U �dR�yN��m �C�_a�m����֊��V~�9�I��B�';��"��6�����]�'����j��aG�� �߾�H�M2z��gp��h���C���������i��q"2u�1=?P1�dm[8���\I�{�_{�������q�"������������k�WE-�3���P=Jϓ���C�R~J����i�=I��z�~�!��i&<O-Ċ�Y�7hf���9���:ɼ�0+��8���U~f��&�R)�5<��.�������~Y=�xC�:)�N���Gd��FJ|���[q��-����h�6��P�� Q���yw��`l���4���7���73`�1b���+�*��s����͜��ǩ��ԫ:���V:i.��滐�@��p.7��~�ץl�:f���#�Q��ȿ�������<j��~������$�0�q4�u�&��^}��~C�ć�;�N�X�L=LMr��if"�H.�z�KM&��P8�f�a���&3ɻ&��+�XU,��馾̳����v��{` D�_�X��zw�a����|氊�d�sjm��Rq��3��OP�?�
��X,�+��CL�&0�^&$�E/�0?'�m �p;���*���|����Lz�dx��j�&�=eg�Xm4��Ru
�?w2)6�f��$�_�?:AO�P�
�8���}�g̕�_;��'���C�~¡��LLx������FN.&���Sf�i�U��2�
���G�=�4�>v�H.!�C�I9�d�n�t��S�]P4���V~�0���I�V�a�Ԙ�����p� ����g���(���{�.��&$�
+�7詪j��B����=������LB�d��y��|�hu�� ���f>�}�i���5�_�q>M'��Ԛ0*��a�m��1���d�?!X��=L�9���P��`o~Q/�y�R���ue�}����06�J�@���EaXTǬ��J��I^�ϭ&�T*
ah/?X�µ���g��O�ud��ܡ�?3`T�>��|I�+������6�)�|V�b*�|G�A��d
�ϰ3�&0�w�ju<H/����h���bA��k�E�A�%f��%d�Vs�xZ@�Rz����+"������'���s�q*u������!͓H��'��Ngި��Ǽ`ϙW�'���;��u�2bc�=������~�M�x����{�ש����䟟wt1�5a��4�
q=�������̜OXm�J��.�}����~�w�9����8�w<��������zʑ@�+����~Y�LC�C�Y�Lˤ��M��+&��z\`T�h����|H,��l4�d��O�̚|`Wu8��|{��p3��X��ӿɟ��1��VwW�T>C�c&�1�!X��6~���?!���g�bAx�=�'P�<J�I���8�aXT봞�(J�I\���p<IP�w��.l�T�P&���K.��W#�}J�G,�}��I�)}3n`��#$m*�r�`<T�JʗZ6�b����)C��r�fզq�:�k*�����jE�3J��<;��MrC��s�6�������yQ!������g�J��g=�Z�i�,TuvG]��BZ�$��}��� S�壥1uw����G�~�q�d�N�?e�����٫�|�'�Wԟ�f�Xx�?%���1�0�c?&���Ax���&��z� y��i�E�����&�l�ef�e��|굅W�����  ����t��,�Lg;t�Z�&�>��M$P*T�6[Ι���c���'S�>7t��W�&&>�� �F<�_Si�C�Y��q���y�w�����j�^�Y�v��U}0 ���@����>�E�AO'}�h%@��
����"�I_Nw i��I��{O��Aq�'���YR(vj�2]��&'��N&��L��<��i'�Xs���y�����m������t�v��):y�h��箒
~;��&޲}�i���B�0+�O;�t~C�����i����=Lg�y�V~B�g����A|a�xZi�g�bA~�o!�6�J�C^.��d��z>9=����l����(�OϬ���z�
�_��v�ĕ
���H�v��'7�i�a���;�4ͲT��s�?2�0*y��gω6�~C���m�5��K�*A�\x(i*W��r��|�M]?�L��x��bi��bO7C$YP{Cg�iIY:���}�&�*T7>�!�IY���h6�^<d��^ �P8�9�d�;g̕��3'��jÁ�ͺq�?�1N�f+ITL�?4�B�d�r���)�-�$|�7a��u�1���qĜ�X��3g��*Ҥ���q6�N0�Ri�s��Aq�I���j d��Չ<	���v��ԗu{��xʑd���SL��r�$���@�Vc&e�P4��*Vj��~`Tj[�N<t�w��d��'ݦ��J�_����q<C�+���>�Agc� P�0�3ao�ξ��˫�'��\ཁ�*�;<��C�� �a�{���xΡ�ӿf�a���"����0�*q�Rb�P�Y^~�1%g-���lM��E�0�g�<�T{#�1�@��,lӬ���n���-����5���+��z9��ϝ$�
���ܓh,=k��֧R�c���0�LH/��R)�4�C��M8�eA�7hbJ��h���L@�R���+"�!1��]���u�~��z�-n����*��O�0����L㎟n���+��f1�)�b&��4{�ec9&���6��7u�)V�7-��ZcV�vs��wF�0� ��������H*]�w:&�m�q�\�ͭ��'d�^X��"+3R�n��'�������ҟS`�n�A�[&���ئ��������"����|�]ak�J*��On��Q%�@�P�nc"Zj�޺Cl�/\�Y��ʬ�-͕�� s�J^P}1N�ZǊ�TY������=��!6ׂ�uhMa��{}��N;�����V��a
:��\��F���f�,37���C�o�ӌf	�r�Ֆ_d��W�w}�`�1���f���Mr��S2����wPU!��V���G(0u�sxZ�uH�2�.�s��8Cˢi\��(��6�e����v1t��КO`7��d���W	Ke�2�[��u�-�YZ]{�ab�[sbY9�-�R'�1a|�u ��]�
�˩v�X0�[�Y�X��6�fE%<. �,lr��n	u����3�=	r��,c2Y����,๱/��a���g�����3��f�v�Q[[�"]L��da\rb�o=[	�5LorO�)��2�;6(Vt���S�TggL�l���3�ۺ�#���Bԃ��gp�7�l�N7oo��6Qb�3��Wu���=v�>�J؈|m�\ޢsA�|0v�3�Š�j9�E6^��r{����nb%Ѯs�-')�JNɉ'7Pd�o.�b�wJ��9Wؠ�yԵ+���j��{P���+�8�����K0N�R�&���d��6�T$�g���]�XX�Ʈ���ӎ!U���_E��#�ܱ"���y����or�+���Id��v A'M$�>���x��z��\z<����dcY��n��܌7]�g�+	*���^�u��;��<�5��:-�	&�p���8� f���Gz���"�f*��#n�xqf˽a�H��k"���S�]����^�X�8�t]�%o}������fG\6�{�DfG��3���R M*���ۛbM�J
:5�$�K‽�"D��}�1l�e|��ˋf����/���-���j�35A8H�F�ǝK�t2�A9�3u3��ά��mF�c{
�Uu;����b�rv,(>]�cn�Y+i�ٽ&c��tVsb��7su�P�m��vr����^����g�
�� V���v��-�cv-� ;!g.��A�����N
{-^2�Mk�y�)5
����;��N��jrr�+���g>�t�
Ў���[�q�GlQ���v���n�,����#�R��}̌��[�jE��EY���*��)�v���c����WX����4������}�R!Q.�#K�u\JfV�J�z/�wh�Ȅ�*H����K�L�ʬ��e����u�Ձ>E�z
]��� t�$"���H��ђ��U
�R#UX��U*,/��%J��j�+F�*����U�*���[V*��X
T���(1Qb�m�"��$Y�3*���Ƌm+UTDX�J$PU�+F�J2QUDDTլ4��2٫,�1�k
���QTh�UQB�M$*��TjV��-*�V*,��U��-EX�clV"�F���,-�R(�$Q`��ѥq**�**��c*,��
��2�AT�*��V".	U�i5aU�"�EUk"��cX�+�ʩTTU����UPQH"�r���RТ �J�1UV6�F"�*�R��KJ���C2�*"�"���Q�0c�X�Z�T����T����m5�Uam1�&Z6�A[e���m(�UDAA��Y���.'�a�Ɖ\���X���ep�D��:VM\B���������7V�ݝ�]wHٕ��'V=�zj���������g�_��&�?͡�AH�~Msz:������9���~d�c�=.d����M�h����onI�����䎬�x���;���8�����I�q�}��u�s��|���|s���x�@Ĩvj�L���ĚE*A}gX{����!�㿵��+�T��s��|�rΡ��ɴ�Y�O3���I�;�d�W�
��sY'�:�����}�Y�}[_[[�V�T����T{�_L��^��g��m$��x��|ʇ�6~��q
���aS�{��z���Cy~��uLJ�p�sHJ°����M�~J�+���U���/m�֏�/����*W��rm"�V�u��f0�g�yl�ͲV����vOY_Y?n�I�uĞ�_=��4���Y��1�%H,�7�u<a�6����sO�u6�c�J{��K&����jtO� �@�G� ���l�@�Y6w�jm��d�
��ʓ�Ĭ�k��x����~�=v��d�S�O�3�K�xO�N�?'﬚I�+��I�l
��3?w��pn��wwIs����P�z�L���8�ݓ���l���$��;͆$�k��AO�TJ��rOɶbi� ��������O����<g���"�MRq4�.Y�5翯��G��?>��o������a�%g�x�j�R|�l�W��߮$S�?=tÝ�!�m��d߇}���������=OShm%v�w$�1�Se�&�1
��g�����6���W|�R��Kr~ �(�& ��Dǌ8�&%f��bR��<�u��:�=��m&߹`c�7�Ch)�l���<AH��8�������%g��S�,�e}a����I�~�﫠Dw6�iB�75�qQ����Cĩ���C�Vg��6n�=dR����{v�^$YSG�g)*J�����m�vɌ����m'P�R�~;�h�B����9�= �X{r�+wUu����D=�&n߲��޸������6��WL�L�3�$��'��I��ALB��~L@�h����|���?X��!��O�Ci�/�8�
u
��ܺ@�Vq8�.��O�ǖi�A]�S��c0�/)��&R��c;B�ִL�Y��79:���;��`�!i`�7���B����MÍ6�hooT��,s-��l��9�] �W�|܍�HgvK51;$=�C�	t�ΝCA;��U�N�[��'t�!
{�{�  ����&ټ��1=H/�'�������Oӝɧ��&;eI��@u+4�r���H%g��l5����xn�M2U~`Wz�)Ԝx�ȳ+�O(_�<"2 6����	U�C���]M�}��OHz���{��2������Ρ�y�E��|���9�i����|�'����4�&%w���VT���8����i�,	�g���
�"��j�����#j�|�~�u�i���
E�aٛ��HVm����"�n��+�~���m%g\I���0*a����Yԩ��X~M��|����	��q8�bAx�OŸ����T�������_{���^]��g7�%�Ww��G�=l��xY�@��+�T<ى6�H>�q�����=�d=LN2z�=O��Ch+�&��4x��Ri
�k=ԛLx���s���ɏSo��4�dm��:�=3�s]��z|~��RP=q�Xo�6�Z͖��H)��f���Ԭ�z����<J�^;��u'��>C~3�?��Lzʇ��*���vs�nu�� T��W��~� `z����n��~s��{��|�f����Y*�d���m"��׮��1���3V�}����?0�|�C�?]5�PY�*jS�4�Y�~��lY�&2xg2i���c:���z ��qL�:b���52��������� �c�}�z����L@��~Ѵ*J�vx�	�1"���4��g��i�״�f�oT���Y?2�w�@�N3�!��8��)��rz��%`w���9�[�k彏E4�˯�<�� LxL{ ��g����o�抆��'��jb�J�S��$�ݓ���6�I�+Ԩ�Rb�i�Y?:AH�5�q4�d��<?~�4�į�4�e�w+9�}����b�ltx͝=�m�'����~�M$FN����w	�u��M����Aqs��^$״1 ���O�ALB����<M�i+:�'�l�Ҥ�=I�� ���������ۻ�{�g�"���&<�{̯Ol1�Y����Y�L@�+���:���g�}��m+%WL6w��R)Ěw��_�+%w;�jL�O�xw	���M!�6������_Wˣpߒ��1}���3]�"S^�!�\6�,oQ��
�Owm7G�U���w_/�HF��J�sn��l�������L�w
/U�Y�SA�:�:�T�nX�)�az�k e4�(��t^N�4�*�|�A#��6���~��:�k����� t	H)��1�=a�c����c<|f������M$P8��&0���&0��:�B����s�m&��)];����"����=O=�+4����|�-`��7 � `L�{`F�}`T��8�e��i��Pvk!�=JɌ��&0�x�5T��J��:�����	���6��J���kEd�+?vɟ����N�^%��q�l����v�Fؗw}��=��������M:AC��?%M2~q�9�̛@į�y-SO�
������i���AH��~LM��c8��-�}LH.$ֽï�=�Ho?u�E�1���֞+�����q0@p
��0�J��V|�w��<@����p��z����0�?����>�(%g��hf���9�4βo/�
��!���_��~��
E:��s������~z���V|LT���X��>�4�]=�OXu:�C��O�
�Β��LC�&$<9�ju
Śa�by�`x�Hc17o�A|a�yi��T��5��'Уޘ�����'繃L����	]ya����i
����<큈)p��a��R�|��@�s,�9��6���8��3��OP�?�+�`��6�CL�&0��o�xD(�����g�u}��/�_/�t!���?����ԕ��f�L�������1*O�������B�sϲM5������@�S��3�k�%@�W��d��oX���CO��0&�|v���b=9���@�S�!"2~v�8��ve��ɴ������d�ݘ�� �P�M�M |���0���<J��~�i�:��|���<H-g�1ߝ��)T���K�f�-/<��`��g�;g1'}�
�g�����t��Y*��̀��S�P���AeAe}d�����k�0�|�O�:�O�Aw�Ì�!�c%�������KxҾz侂"����l������������$L<�~�x�%H�xs<�XV1�&<풦!RW����i%B�������,+Y�&{HT��Y1��(l<��4�x��U��]++���٬�=�������G����uL�G0@����LC��J5�	�sYջ ��n��//0`����X�C4�U��f�(��1%�S�fNծ�*�VUZ�_j��*��j����㒮�tn�6ħt�D�i�|�L/`��k�zX0�_UW�}����֛ʚ��&:� 1��#f|�q*;�i�0�c';�SĂ���]֍��:�$�u��m$��s2JɌ��,���J��R�JȤ�+�l����=Ý��5����;Ϗ/߼�>@�T��}��l�J����N&:`T����~d�Ǭ�/p�H#&���U6�Y�'�=z��\No$������<��v��8 �` t�?�z�]3_E��o3�=��'� i+;�&=g�1���<�������m��P:����>dߖm����Vu�2�'��M��+&��z\`T�����ω�>톟̝�4��Owgi�|~�{�����f���!Xx���̚BT<d�d��>ty�����lLf�'ɣ��I��p��2,�t�p��E������]�T-�F�U��d_�m��Ȓ�]��EϬd���g���|�m��*�O�X|�?0+��g��z�}I�cm`�ľR�0�c>?Sl�6�^!�ϲi1��b��᧩T:����}}�{u���=��㿹�o�s��4�ɤ�'���Ou�䭺�y��w��?��Z�x��Mp�r}��=���
�.�]�|������&8=��+����	�X�O�{]�`��P<1��:�X���[��Nk�4�`R��:�ej��2���8�j���{u�>0� �.�U�sI�o��)�+��op�Nh�+@gK~Z� ?��o����$��Ǵ��*��cs��as}�d�=�&�"r�U,u�m�G��K&��D+�bL��!�+�q��L��4���v��;c;}�؟{�}����;��Qѱ.�Xx`��;�V�Vz��:I��f�΅N�ݮ��+u�Ӵ�S�G�e����WqY&����	��^֓H���_2#�i\��8ىnF��}��4kG�W��R�[6b*+�
������g3$���ȿ���
�Bi�6V錿�p�4=��E_*(��m�;��X`���m�g2淚��/H�i�W`�!ID���:�JD���}f�R���lH]���Kg+��3�b��|� S�:�<o�j8H���Eh�?o��}��k��$u�L���>�2{����p�E����ثr��Db|*Y��#�,1Syr�Ur�����ֻf��(H#2���}�K�F�̽�21:������J7��ܖ�8Y5:��CJ��I{��&V���, �]a!P��p+������!�.����C����<
N��x����ʗ�5�r�cX�~�.����U������C���=�=#���g%�\�^�f�'^SC��Y���V���Ja�k)^�n�[�:/��y����FS�|$�������I�O��t���YDP�t�h.wD�l�t���*�k����`��l���l�!i��t^�F�Ţ"|ұ�b��5�vA��&�~��h�b ������u c8�\D�[��L�	:b�p�K)���>]���;Ь��H��w��ϮPB�v��٨��EqQ��r�+GbP�Η���cl2��]��#���`5a�Zi�gg��Of���m9�9dc���yԸ+���������=K�ErxvcZ����oG��subVj�g��S~Ε�=ٍ�7Έ�=����m��tK^�q�nF��:�lQl��,[נ��X�'m[�tf{X:��jL��^wSƅ��q��`��rv����!|����2��洉ٚ؜;.�Bc�j\�i��[�[;b�P��j�%�J�}����`n�M�+��]Ƕ�n��i��ɓ{�z?x�9�������tgb��W�����q2�?^�57簤&��]�kcc�f {��Ĕ�F���+V�-�9��VI�T3�f_���]ƃ}M�\w��.]+_OUe_�F���ym����#y�/��4{J�xʗ`�OD�N\e���[���U@�~3��#yԎ[@])<�n:����'L�;����>�ڢOV��}QR��[�i�-ߠq������3{}�{L�ӓ���5j��u�]�m���4������5n�z�v�%�����2�1͐�5ݡԄt�a��2å0Z��r�I]��dL6j��9j�?���o44w2���y\;D�fK�:�]b�s]q7�cN�`�<�C����}W���ߣ*�L���{��q���#�>ð��t�{6%�nw�Ծ����9U�5.�(w��>��ܜ����չ��O#4w/���w.o6ũ��;:�uMx_ �y6$4�K�89�t^�|�3V������nl]���q�<y��>ɧ[ζ�XsO)My4$4��^A�.3�-�5��;b�j�X���y~�q���d�/+y�oK�y��bg��j���n�) n�w�p�bGP��^����X����N�闏�n4g����>��~Lb�3��rw^�3XON��Y��ܕ^��Q�~��<�kH	�ޥ�tqa�2g��4�7]md��a�wB���B��5c������BX���SǢ^>f�6�˷p�:�};b�0��W�:���F]$�$U]�'����U{�V%�Sܭ�alduَt��N�L��Ȁ^���gM�f����g�����V�G�g��S�v�׫�/���<y׳�o^�|�_/����r��w|��q��z]����_��"�ĹbD-ȋ�"ǧ���kd=wkq[����P�V�/�"K�D!�(�}Z���d��P��j��8�.gG��hI\a��z@���Q"�v��<"���kY��M<�Do4&r�^�����/�4��O'u]>=7j��6��'�Qb֚B{y�Y=�.���~N6 �TG��yԎ[B�}}�
y��m�E�]�"��E�1�yofR�_��w�lI�n�q��|ui�{\�P%GϜ�^��mu�~��҃}��'O,��`#a�)����L�\�5h����-�^�^F=�;��M{��w�lO>���XSnk�KM+� �B��[��or�A˽`Bf7�S�ǋ��tv'��1/��Ŭ�J̝ѵ����d�:K9���{�#H��>�Ee�T7]m������m<��J�l<���X�eP3�ݠ����6�O!�\�2ֵ��k����,�v�����OKy�Ck0��"�G�[��eR��^��] zJ�p�r)�"ǂNYH����\��m�^�K�.�s8FW��M�q*
��jX*9z���I�G���x�K�~��v#�����fvb�J�!P�&�)H+&7�;v�uv^ks����î�����";����P).v�X�3�߀�����,��Wd��7O�>���~;���-�;4�<8�]k:����8E�;5]���+U��+^'mX|�1���g�m��Z���v�-�d�֛~�=S��b_!ܹ�SnÚ���P�獑;8��˶4�S��곾� ��%u	A*]�؊5�*
{�������<y��2���|�<���W�T$�P�iX��-:�|��x�p��m�����k[��٨L_w'o�����q{��Ϥ�]�υ�a�e4+x���[zxgj@�S��~��lw���oc!���X&7��L�_����v�r��a��X�'���qn�}��f��$����@��s1<j�?��E���V<�g��ϟ>��[�y����=F�Q��3w�����k�͞�UY�b>�� ��!:�Z��9>�~����{_��%�vT9�,\�{��V�]Z�����=ɤ^�~[�^�VD)ץ{�d��Cpg^<�Zf�H�<�c��1Վ����Ԝ�k_
��t�Jn���#xk�D[ɎEv9vK@W�^nf�͐#B�Z_n��0�FՄzЉ����=�E�_u�U2��d~6懜�H�B�%��Z���fs��Ď�|m�V����v��e<�U�ꛓ��c����I�2�)�e���j������KYXv�[3uf�n�i~m���Hm?+S���x<�5�|���q��a���sM��I������:B}�w$��K���iX�1��<�������=q�3���T�Ycz��}.i�	�ٛ�B[��mS�J�{��1w4cB�~���O8�����N�镍:|�V��g!��MP��������o��v�≯<�ӓ�օj�S
e��0��9V�s��K"̞~���ƶv�,*�]�T$��(wW�K��>�-࡚Y��f��.��^��.wf�jY�ݲ��ى���y��L��n71f"��$x��qi
;yLbڶ�OaHM'bP�s~�x_�O���*�<�Lwl��FT��c'��3v_)E��jb�}���*�֏�åun-�\��P-��Ve��(]�m�E���4��􋃣A�մ:7F�oժפ�,f��9֧�t�eu�@�:��\ĩ>��:��l�q
^�LyV)��Z�a�[5��l<r�w׵5C ���oKU�Ym�!��逃�r���-�Q��&���2�P�Q��(d66<� &����y�n��8����	����ũU�v��w
˙�[��6�<�r�L��"'.����5f��[��r��@�͜ʻȶN�;[�dUل�"��T"��M�aj��b�ʉkl�e�A�8ލ!n���WE�7��i<G�V���wE����>�I�׵��,ѩ2jڥ��J�;,ۮ�Ų�ǧo���ۯ�f��	�wVxMuU�<�i��J�� �.�Z��ۙ�}nr�+ 0&�#U���Gj��3�<ߗMi�嗣�h�ʰg^�b�0�ˆ'�N�6�Ġ�����Y�լWRxJصvSY�ھ:�ZF��<)�E�f�.$���V$UN=�XCL�ף�����	��hn+�ԓ�q���L������՞oj�t|�\��l	�p_<���.�P����\��bw���}d4�omc[[rs�����v��ʾn����lJ�|vV�M�ƫc�,Д
�}k���C�=�]^���k�z��E�������'��л�N/�6Z���a���X����G��&^S�}m7CX}aC�v��fgV�M^��,�l��^yǔT��A�t�զ�ܔ_*�uuc`�Ivv�xj���� 7�4��icT��@�zͪݴ���,��V�1f�H^��-q�lw-�y4N���jʙ9-u��94�;p^/��;��X���U���3.�.jr����K���灔�l*��57�\2�0g
���)�*{R	�֯mE,��Q���!Y��R�x�1�f���	�賴m�u͖���i`�[lv�J�m{��{�&R��CWэ���g5�o��֙�cKC?>�h�m�h�y��(�})�c)�}Q����rqt�oD�Qq�Z~�;�eeV������*�h �k���qM�w�c\��&:9�w����i��Rٵ�S�@��R�Ah������Wجm�Z�nLBT���@)O��u0���<l��\�9���7t������h�J�-5�Q9�z���:_.Ҍ�_j��tXX�-�E=�ͅ�|�����ރ)�	'�Ү���le�6R��x�8�Ե���n��c�"Z=�3+��;!V)oS��uܳv�8C�����K9Br�+��)�䗝t���{t/
3�9.��e�i��J}Õ�\=�	�6�9w����p8���g5��˴��u�1�\�57E,]p�O*����3Z��k���v^�Z+�8/O���/�W�U��|�}�e�=<Ͼ���.5�|��,R�`�E�AQU(���QUQ*V*ł$�U�Ƞ��H(�Ve�P,X#"�lq(��X(*�-J�E�*"#Y(��*�E%B�A���QV"�EU�"�DX�(��hk,Օ*�+YPa�B�6ʂ�*X���c
�ȣ�U`*�b��V(����TX�(1��PZ�.�AX��KiT��*�Q@EV(��Ӭ�QQr�uq�2��P�T-��cPD1+UPTV*8����Y",Z¡Z��*�Y���UkE�J��,�Q�T�YD�+Q2����-f�2�e��AIU4�E1�V*1
"���u�C"��J�*,����m�2Q�1TEX�%��"'�A��1�y�K�e�we��nm��s�C�9�ݼ�^��N�ѿ�#o�w�D����J}7Tjd<ءr�@���b����Ο�<<6�^�O���4��N�L��Vp���H��h7���c#����NrU�"�5��	�E�"9u%��U�̍廍��O��^���qR�v1�ؗw����Pq�ڞzG-�����
����ME�
W�.�mn�j5�}e�T���.����8-4-rU���|�V<��*��==��kB*�\[�����78�l9��)�auT#;���Ps0o/Qk�����˕�2�N���>�l���%��$�V�f[��JdԶ��>Z-�8j:��ܬy��3��i6%�b|�N
�<�<�݈���.��n�.�CrwX8�,O[�WfW�[}�9y*wɡ-#g݆y���"ۢ��A���0�����0*e�Sر���~fwꟍ~y�<ز�U���H���(x������Y�򹶗����ު����82ƾ.gF��go�׻/9z�����ۨ���Ά�u�*�#��)=���Ƥ�ax�����3J!W�+�S/z�Of ��]jp��p�i���}bCo�p��8���ť]18n��w	+�aU�m��f�_Q�1.ru�����ܻ9U���ί��'���a�	�к+=��em��p<�gȃi�r���p�V��;̴�4��or񭝺XS��0s�R����c��z�7/�Xw����휐-1#��6��˧л:�~�ڑ2��
��OY�j�ܝ��[��bN������=h���${�y��.;{:]ԍf�o��R�MWb-��]^��zKJ��k���fgԻ�ec��r�%��px�O������t�(Y��CJ��N�WH+��o'ܩ�%v�=�{z����s��i�ӿ'�@J��=��G-�n�Z-D;@ئsvaf�)M����4.�q��ڷL��z�U�7P8�Xd��1�ֻ�f�V�����L^FO'��j�N�C4�k�S%/i�X�a�p%z��$�,��,˯+�Y��ݺ��hCby�]78��ۖ˻�4+�>0&;�z�)!De]�+K���# �9���[���;��F���X��P5Õ��أ*,��cZ����;AFN��ˎcW��1�WvsY�1%)Κ�l��3���˓:���Ն��a���'.�U��Ѷ�E�,7�mݧ�?}U�վ��3�չ�At;�Ƴ~��#�x�&��E޼�l4�BʖF��57��UK��(1��hP��R^�X���Y^ɵ[���PsCf*Y��#�j���v�t3�K|l�����7t��%\eg9ɥU�M9��x�7˺ʚך�+e�y����b.}#�Fd�o����J&a�s:gb�s�k�Ce�2�D���K��սwA�n��ONס�]Fr�}�b���O�]�a�Ւ_j�;?S�>3%k���偍l�K
st�FET�<��W0��
ʞ�X}���Or�mSn�sY^����q��4#��`��7w�n��=~������aw�g�F�%
�����*����b�yk�=���"':#��%y=|�^lyW.v���̨�����MG[籑ԱT�0Ҡ$�1�f�>�3ݳv&aIʉ����F��u3m�Fƪ�NH+9��w��b�V���{��Q�r��,D�M)��.�/l��{*���a�O�]_0v�Ɵ�pKq��k-��e-�R����c�
+fJp��:������������N�ҕ3��\�����5�{�{���.l�;��2}O�����d:y*����.��`]�U��}��&�p𤗎��]��qn�o���L�s��=מ@nyH�������mX�+�x�vH���Ϻ�
���+���ͱ�s����*ﹼ�٩���>�:�@�L�[�A9��=��r}��g��vc��Ӹ��v#;WѯzqŹ�<IKbv}\�׃-ew�ܼM2�s� ����m�pv�3�Hm|M��x�}�$j���R<�k��@��iE�����R�sO�^��ZBC�6+^A����/s �ފ:�s���{|Ƽ�.��okW�R�M	�K0޼���u�Yت��Tw��f��]-�j�9��Z�ر��$�ޗ� �\�U�5�3
�F���e,�i���~�躌�Ss�(�C�-�Ӫ�镏v�xUF2k�Kȁmu���3|$nlޕ"&�{�K�2V_����3A�1�7+���c�����<&8���ī�=>ݞHY�y��j�$�֍�C�P9����*����雺3�gE���I����~�[!=�q3�]�)���jTy_I��G:�g?�}��<Zd��P����ח=���;qc�ίM�u�'��5��X�䱸z��a�b���.�V����j�%�zP�X���x�^�i�2�~���y��*���@&�]��1>2��+������	��+�bUt��أ�i�v"���Ri;�9ldw�>��>�z�}x+ey�f��� m�8�n��D���F��=����F��D��Ku5����eB3=��[3qۙb7���H����W��]��:����<��x�z5:��rV�v�z��{bm���$��g[���?�EN}���V�l^N�w���i��\����Sh:n�%Sqr���Me���v�:7^nq�FÚ钕��Bce|1BhB:�a^��HF�/|���ښ��p�c}Ϣ�7's�4:d�S	ޢ�Z���?\4�Ƀu�5}��]�MvD��CN�.T�GV�=nW<�Ì�um������گv����=�r��lŁe����,��b^m�]}��չz�Nˮ����"����|��5��)ȷG`��Z�hh��HqL]b��?�}��^�����AL��k+�}�1c�;����f�a�c<�N
�<�9c�(q)Fb��3Vo_����̿OZ�W�ɥ@o:��9���MN`��{K��)�$���=T���������*�+9�N��~���旅ˢ$}�v�9�7�vX�����"�G�h��X��^ϓ��
z�z�z��ɻy3������v���=;BE��h����)au�7K_P�&��WDwg1�)6e�y7�x��إ�W�f_�l�� ��IŽt�v^uxV�����Z�
�v�۸]�i���H��u4+é�qn��W87�'z���a�;�|���K����f�þ��Ʃ�܎m���Q/u�]�瞒�zKJ�U;[�[w/k�����R���C��4A�}7�r��ig�Ȓ�}�lH�w�$�ў�)m�y4���m�*�j� w�K;�X��J����vM����u�ɮ�ۢV�׆�༆�%z$��򅑍B��D�6k��ÝZ�1���u�c���*���9�-� ��bPܚ�a���-��{��ҥ r,��M����Q�ȿ�U�T����OI���_{�ɧ�ӝ�i�à�V�cw�b�M��2�-�~"�ܷ�QYSl�p�^��޷L�{NѰUy8��Xn��U������n�=Z�nny1#2@��#�w\'��������`#a�)��(	:�<n�V�����^���mf���s��0�ձIP8�8�����t�s��z�W�f缨e��1����bq4��-�[��d�,��L������V����{`ƨ��~�>�yo԰���v��e�=�[��vm�������AK���6hk�<魍��y�k8�S��^�}��0$V�JT��9o����s����mf�"�C��t�{�;S*u��˥�8���[Y]��t:ee��|���y۳6���C�r�;j��v��.UKQ؆z�Ɨ�zekN�=Ylc[;��eR�E�N�&#�.�k�S{��(nU,�ۅ�n�	c��{��ŕa$���_:�$SA���~/
}yݛ��X�ҁ�5�CIp���;�PY�	%��ЊW�Vc���M��^��d�Ҷt�ZΗl=�)u9,��Qӻi;�� [v�R�ś�pmW�e��%�1��$���T�fn��]j���ɕm�bd��C�9��p��r�>钂U�ϯ��E7k��]�9��[�=Uj��?3�ֵl���H�L_*�����J��|��0���rQ*�<��v�w籑ԱTxE�L9�ׂ�/�5�]��uL���~�g�+S{�X�}�C}N��Cy.�ʊ��tիZ�mD�nq^��F��C�^9m]����u���󝤞�]�m�ꍛV��@�T� 1�(G-�#�j�.}��W��<�	�õ==D���]��Q�W���`�'E�8�L�ynX���B��f�>�S�W�+�\�tgD޿����|'ܧ�ԏt���'K�n�vc��2����61զ����w�D����n�I�C�9��/�D�ܼ�]5�K��{M�j$By��隳:h������SС�Eٴ��	��!,���>�__�w{�E�GM�]���d���ɹ����pI|%����e7'xPӦ��E3���N¼��fP�s��5)�5�5Nn�K7��iX�je!�
�� ]^!ܘ�;���7���� �y6����lW���o�7n�R���Y��՞٬�b]��z2iV���v���SI�!��lk�9:*����n]x�*մ;����Iv��������^=+7��O���Rf�\�s�[���@�nfz��u�z�.�ÏD󎡈z��\J�Bv8���қ��z��o/���y$����H؝��v�؆�ʗ�i鞌W��r���\�j�f���%��mK:�%��K
�!]�U%�J̩z��&�y��!'o)�z2��m����ԛ�wM��U� ��o\������Yk�}�WEO�g{��\��U؊r�&���gZ���M�r�y̳��;/i�bzz����:꒴��]�8u�g4��������S��it�&r�X݀��xX&U'�ߪ���2�yn�c-��q�ڦ��k,�kz)��!rt��8ri��3�wkf=$�Ҧc�T��6p'��0������Z8g�oAw���eN<6i{]-�6��+{k����Y{�l��m>���a=rX����Ď�p�'c5�����n0�U���� ����n�Me�Y��ςx�<��8�	�פrڼ���2�Ԍ0���{o��;wk�̡���{NѰRr[���G����3��B'u2��W�jVLc�y\7�����f�E/�H�@�|;�۝��`�'F�|o֮Mr����lt��Mo7�Ϣ�7'x��%����f�TN˷��c����Xy]Ӿ��wT���Ɔ����86Ǳ ��^��+%�]�L��h��X�ooVa�{ζ�ki�)�r��e��\���N�3��qb�»L���!�d�������\��j����/���UT�_{zT������Eȇ��f*Qc[�n��-�}�^�#4��s���FV�O;e����o]з�9a=;BE��ntX�.K�׬����׸-�Yի�I�4��os�Υ�U#�61��l�bm�#�m��o���WC�ʵ�}�|jY�v�L�Y[�=5�)]�8�T����-dO,�l�JͫVu ���RP�f�z��h�mMq��:��kh�4ӽg._D5m�P��fu�!nUw`oViО�
�g19�)Z{�{��0v��[�Tu��A���S:!T�'�Օ����1�x�m�d����#�U/G�A�|��,jsW��C��f���?C��Jz�v�f��ِ������XQz@hܭ�+{��4(�98� n@�	:���6�a�9�i���&��<`<����#�onAv�+��\оc9�}�˔åW; �*��SrF��ȞF��sG&eV�+�t��Ib��ӏ�_���J3]���ӝ�7�S4���ӫ��MCc�Xۮ��-�ivͻ�	l��k��}�\VN�1�����]]�{�ft�tB��8pޒ"���P�c&e���jiם���&�G���~�SmXX��p�#}��"w���|/ ��[����UǶ&t�r�7���_��%>�І�>u��.w%Z���%�t��;a���h����77'Z���sc�a���`�$Q����r����Ӷ�m�ř�8k"��nu�W�mrgb��o6��o�1P�����lT����R�ԼVy��ӄ&$�nm�;�	�!y[��,�:ezle�3+{�2"��q;���s7���.spCdY�q��.��S�z���w7~�:�XYa�!��X��n
yq�E9����f���}F�ѦΆщ���|rX�YP<*��+,�J�vt5�E�H�׭Ei&0<�j}ѻ��zr�H]gfL��x[�& k�=B�NWs�U�
t��y��o�;�{��n�W�Z�xЎS�s+5ݛ�Е"'3����X��Ip��٭��S�=Fٽw��k�#b��'J���wv�7]�Sx�I�����54��YPP⯗Wa�1�%� b�]��R�Ƅ5rfZ��d�n�!f���&��\k���T^��I�N)�6�F��S���Qs�fK��M�����%X7b�ViL߃9�"O�a���fq��ï��=�.�h!�:O���#�����&ë���̞(-�pѣ�z�&r�4nd�n�j.Mv�i��_vs�m���V��;�U3�)ӇW]BEjԧMoF�t���7F�Mfc(�M�ر��X��Y�N�*��Z�;%,ffJ �&�+����O]ԣ/�{B�>Z�=�9o�N��ۖ6W�2�G�����ٙ�-�Kە�Z<�CXT_3�H��ۇi��$���o_%iXN��7і����o(,5�s�ғ��ٷU'S�4rsQ�zv��V^����1���-�1�fl�=�TU�:^���IT�'U�]]#b,k��6���4q��DSvT�^WcRJ��G�$��YD�J��l�m�D*,�
�ŔE�2�e�֎ TY�I�Q-,E�("�EQT��0D�(�Fj��A��$Lm�#��U32\��\�\jT�P5lDU����H�QER#QAb$�\�[h�Ea��ETQkP\�UV�J"���&e��1Z�A�ʱE�Lh�����`bTX����DPb��@E5MaU����PE(,U�Y�Q�J�5k#�U����a���1YYPĮ%��,�TUPKn4�Qb2��%J�E�Z�YR4��b��kUb����J�Q��2�*�V���%���J�J�ATPQT4²1`���i҈��Q�Ar�3)����!BҊ�TH�-,�Q%s#lA�p�r�3�F���ƢϾ6U~ ����ѽ�IMːB:��Q�v�Y�q�v�i�ސ�U'X��r�>����$�fZ�d�,i�3�w��t�����~��'x��t��s�'���J��'݋��M��n�.ΰ���;�uZK��}m	5\a��u�	/�PJ���_:�E���nel��)��.���ڞ��W�lgFGRlă8P9��),R��-vN�3�7���B�e�}�]�ڠ�wy����du�3�hM��7��7��ns�}%��W`F^�y�U�o���w`�2i�4�iZq���D��ox���'���dbI��pmc��
}�!^���j�3@��h�*���F�8;e��ؙOb�U�Ωf��Ϻ�'��C�A:yt|��W^Bf����������-�w���v�/-�{��\����9�[�� v��a�X�n�e���y6朣�b��i����o����i����5�So=�]�}RQ��z<r5�i�u�~L��1����|�y�ηjv��
�@=&c(��v)��(p���(:��M��nw�wJ"WA��ו-�:�w)�R���F��$b���f���Jw���������KWS/��ˌ�d�G6��x˙Δ��)opڵ$̝�$��1��&"^�ꕴ��@JS z��c�t��xoOnʹٜ�5[yç�<@���4{���F�����WQ�6""j�	�����ldүs����9ߞ˚y�Ck0��\�G�b�_�j!���av�������Z��VXާ�KV�yٓ;���˫�:o��i�9.���hư!�6w'�u�Z�^�镯<��>{�of����˾U���a0o�BmU�w�n{/��E�2zx�{ޒ��$�[=��!'/Q���&�v�B�
�F�����eϫxWDi�����i�#\���On��h�=U;�d�M����|��Ouze�6\�j�"�v,s�{{�������2)�Jl-�S�{"�q�;`w�2�s�~榫����-iT�M''{���/��ԷlbE>�M�;{�vO(�Nۺ���.�7�M�~�b}���tc{�pqŻ����9叱2�j�vr3ʱ.�,����}b�p��� �%3�]�8r�܈�1��u��򺡗{�Zиw<(S��:i�-G�<���*��+�칯f-]|{	ޘN��	D��O{ �B"��fq\���I�CZiG����a��"�d��D�R�Ģd��k�Ϫ������V����ب�U#�E_H|��8�r�%�e+�SJ�6�����Y0��U�f�u��p8�A{��r/!wk�k�ب��ֵi��7t�-���:���v�5�% w-s@N��;d�<�Ov���r3�6s&:�&[i�6ĵ��7'x�L>��2��Dmj��z�%�k�Q���sn���T���M�i	�ء� ��o���PB;!^�yԺ[�3��g̚�|�$cO��~�g�T�B@i\(Gw!�˭y��������#nz3$�誋�|�'z��y~�]��奲�h3Ӕ�Ĵ����ٛN2}c�b�	�ڞq>������囙V�~�b�횛S��v�}�z�^f�zv�����rv��!��]��ВXs,ֶ���s�9��{5�N姢�j�!6�;V��b��R�B�w3���[�r��X���Wn�/�[��W��}��ii��F�۱��^1�_oq/�'O�m�6�Dq����T�9�>8�մJ�����M<�}���;�SSj�54�o']�a:�R`N��4":�JCu��7�)Ɯ�{���Lgcq\�v�v���I\`l�9�}[�����+���d��w�	�g�~��zm��vY��GCX�L��%�s�,��C�]��%��-uW��f[�.wT>��:��[�*
�y�<�fo��vД*�
�I���f�js���[�v]m�c����~��h��'��xD�#��R���>��2^V<o�#ok�����4.��y��3^/i�6
�ẁ�XcV�+J��!㫻��n;�Ν�N�.}ɮ�	�0�'4��w�l9D��Z\���q뗑�3��yt�t3`��s��4!�Ϣ�78+����
ص5�0��սR����7�$�ܣ�����l�lKH�vY�}�32�����A�a���S��2�*�*���+������F����S�9~�a�q��F)��[��7o���#�(uj�om%�k�U�a�VE������C�f�7�7M� ѷݕ�Ba�sd�¦��p��⸬�׃_6���yə���fD�˧\1���.����v���lNb��}�~��٩�v���gp��٭Y��z3'��xUE�s£|p�C�ֵ�KKVU�&���9��?K���a�ks�y33ƞ��27)+f�1w������1����J�
�CzV<	�O]w��M��Bغ���xڑ������kLa8z�G��W�)�N�Zos��V{�v�Wp�ͼ�پ������VVK��H�\��Sn×mu�N���҉�$�-�}���qs�@�d�����Mr;F��Pf��HՕ��t��9���r��b��z�f$B�>��c�ľ룷�h��5;���sۺ���-�'m�\jY	G��#��j2��A���/*��N�z晫W|���k4�'��+N6<���`����8��ۍ��Ww6��ݯ[���ێ��ݡn��^�s�Rp~��߉�$����;0�M�Ψ����Q����ɽ�!q����"m�dP�����˶�N���]���F�n��>�Ɍ-M�]4�J=��"�X��I{N黬��Xa���'V�'^���u4;��6�r��ڍ���v���z� ����͡#�}W!��B��C�����s�:�~-KS�G	t �]1q��O�ȼ�>��5��;���2��'۹�vefdy�����~�rz������yj<���#{��E�{l����Wᯉ�'e�9U��6�y���^���h\s�����XI�=�i��;=�g1_<�sA4��}Ƶ��o�݇�|<���(j�ֻ�_Z1;[}��V7�޸%�]W����n�g�|F/�^1Z���q۝ȵ�Ļ��c6�WL���|���R}�3D�h��k�Mȵ�4�ֆ�pf�?F9����Y�������ek���n텒3SHbR�kg�wWݬ�9^O
�wB�z\�(=�r�r�OOe{L����'5����rn�٬����%��J®�U	/�҇�׽d���^�qE.7��i���ڇlv�͵u�n��"�;w:;"�j�*�2(ȼk����d��s��c-��|��y��YMV�B�Jξ�6dvL�U�FJ|�v�Ct��){:���k�$��c��ٕS	V!�ૡV���9���$���I��Y|2��\��olr[*�6`.��T$�
�VJT���{GL�#0��rm̊ގS`-�)���"�k�0�ǆL�JdwT*oBk�znc�X����WI\���n� ����a�d9̣�]���W�Ou�l����3�53�jFv�lZ�j�4��K�/��U�}PiU�3��y�04�:��3�H�WϟpU����N�!�cޞ�ki,����S�!��)9-���FA;��PNo! 녭����Y<�����N�;�n�uA��`#nx���'f��;j�g.��V�h.B�w9c���N�q�m�q�nN[��z����n֎�'�����z�n}��fU]�u��S|�)��B_i�����<����]Sz�bfj�Bp��������f�k{}�9���M'�Ѵ�^xkV���
؅��v��win0˴1R�=Z��kY#{�;�@��v��q����z%��	PK������'m�{��T%osFa2����bz{G�n'Ckz���}�E��ɏ3{�M�EJp�ꕙ|T�R�"e/�������Gú�~76�,>��d�5�m	�E�?LW::.~+T��/lc�'���a�z�}~q�1o���	�hx��n����n˫��5s�v�g�������Ö9�ڇ�3��9;BP}7mA;Үn�Xn1�۰��>Ij��I��䲽k�r�v�v#n�44�ٷ֒I����Ѫ�K�_!#�8��N]�}�7�^��+-ޞ3J�t�{�۸���+��T��M��S��HM'a��t.ĭ�r�c66&r�s8ÍEk�=��%s��2u�χ7�������4�趹���vCu��<����� %@�>�}�'yتs�o���GD^��I�C�����g.��!���/iXO��T�!g�߈�Ν��l�˷�"N�=�Ψ���wR���O2��a�F�Tx{΅mu��}�t���M�I���.��ј\o1��w�z���Kw��t�-��嵭�X�8�</Pܾ�{v��RnD�vH��%�&b�s���$r�dqu�m��:��������k��ݡx����M��3{��ݫ��2��w3rT;���q�{O��*�cp~���o<��潄��}���R3R��'���N��nmߑ���I��e�H)i�=Υ7����ȳ{u��lm۞�N�by�]78"����R<�dW����z�`��yW�mx�Ĭ�k{����e6a~�R^N�w͙���Le����*/�Fԗ��%[�b�9���\͋���+����O+�@�v���[B|���w�C��̅��U�P�����Qsq����-߼Ǻ� w�8���s�����a�b.D<���O`�C'�d�{I��>�˞�����`���NZ�����v�'�خ�iI+��j��N\��r�O>�B�Ń�U��v�>��ܼkgn"��LtwG���o�5H�U>��	S�'��x/��\ʖ�˾|-���{޺��=,�;��~�];b�10��(����{�_8�p��ץm&�VÓV�X��u�ڹ 񨘓Y�Θe��;Z���n�4S��;+�I:]�7��P�"f35r��7S"����]Y-+��S�W�fN钵��N��e���̮�[pv���L�
�w@��3u���`�(��vS;���M�Y�ٳƭ}�ܬ2��nM�����'�Ht?gc��oVIH�5���ԃ-�ǌ9	�7m�\jY	P<_D�i�f��N���*w�n�M���=�gd�W����M>��{J�q������-n��{�3!	ʺ�.��V�j�r��@�����pOv��5�������L���ӽ��Ӷ��]��#��=6�t\t�s�Z�����{Y��\�}Y-�j�˫�o�)�Kۂ��krS��R7��'��:]�yy�q�횖��u:�vt[f�#Nt���8%<���1��-EJ�Rp'O�Fv��M_tJH6�}��s�<d��Fԃ�u���t�p�82���S�c}�ջ�u�s}U���M)���f��#���݌�ʵ��>��u���Wٱ)Ζok��c�{C�S@'�Ck0ߵ��Ʌ��NO;I��`#&Q6�l҅.��͗�^�N�T�}�;���R5݋h��'�Xl���ˬ)2��d���.�0��]��Bԑ�:Wgzc�Q��t�����f_0�fI3�#���8u꾑^YRQT�,��9{�hV`޼�"T�Dr���K)٪ҙ�^�(ov,:i��WОI���T�T�cU��m6i��YN*;����D���T�E}!�1���j��u̘v�j��8��kaqInp��4qVm��m��b�Y��\�� V�v���;u�@��9qus�	���f�Zj�sYvY�DKr\�/8��p��!%>|���g�g<[�؋���|�Lt�W[[̳{�[K�% ��}��{N��Y6�I�G�b���yݣ]�`O%I���*\�`���0M���9����v'�bI�]���ҕr6k�.�u������59;K2���Y�U�y���9�\���۵GpR��Fhq��Q���h'm���R����V�6z@��x"5�İŒ��>ͷ��9��zP��j͜���j*�g����68�+Q�M�F-[5[�$�-b���e�+u&��d3[��`p+-��	�4��c7��ڮ��{��Y���Ԙ�<�nc-�4�M#q-�Vi.c4�Nc�MȬ饕q��c����j����^�c{��1���.T���yݺ�-���
v�c�V�Q���+8�[J+����l7��j��Z���M<*�Q����Æ%u���I��,�����Hw#�[��!�OB9�K,��	+�'hN�[����>v�'��ݟ�ᑽVu�ą�)�zf��W;��ѡ�!��8��s浢Η�fv�7�k�FC�,%�v_	r��`�2mz��N���И{�{�gSæ�4u��]B�l{�^�]�Fl�+3�;��Zi�(B�s���ţ�:0U�w�k��/ �|�r�o.���K�w��oCH�W>̶��@:Q��O���8)��)��P�)�y/���kS��Z�okQ��ۓ��rd� YCD�}\��gmbg�ܱj�MJU:�8�2�7J;�����y7-K�K��cI�۬b��H�Y��&t8l�t���&Mr��
Dq��4��m9�f��W�5+��3h�zY��&�ƾlV�GY9I���%�s��#oO,{�I,Ү��]�+qY�\���B��p�׵Υ��u.{�ڸw�a�!{4<ocM�h�Q
��4����|O�7U)�*՗�I��S!S���2�|��&ì{)�uޥ⭽ l���{��^l|H�&貹>���v��������15��3�d�i���j���Gt�sn��	
f0z�i�MF����4� �SR@��t���}{���B���fT�I��3�%�opS)Y)��"��欽����������y�-�%M/�J��Ƥ��$�}�*��TY��DG(�B����V���+U�ȸ�e���0]A���"��V�q�Q"3���4�dEEr��GT�,�qj�Kn�85+Ek@Ub�X�Eue�J+QZ�P*c�V�X��JXb�����h�¢,PQ�*��(������!P����:qUj*��"�A1(���i��cZLJ�lKje�ID�U4�dA�U�Q`���V
���QAQ�t�@���$]YX��EDr�VLj,D�XZ�feִe�U�E2�\�p��4��ҥj�(�*"[��R��mDFТ"�Ze�2��iT�T�nEE�ķ3
�(�m,D���\���F:.d���33&0��Z6PX�
��AQAD"H����6�C���8M9�&��{z�q��Kt}���]�;0�r�YO����T�����b�*�5�E_L��;1�k~�}}��s47�}%���2�-�t����>x�]��ELБg6��\�3W��,%�jE����Bzۥ(��<��ī�e��{o֪n��xx����9�K�-��;j�;z�̔��"��2���}h���_>�)=���N���{/�J|9z�����TT7%�cy&iZ״q\�uI��~š�,��ۿ9N���Ml��x^U��3�[�|�y��\�jJ{�I����g{lQsjgս���i��őQ���'��Ɛ�t��i=*�����������W;Գ;؃�}ƛ�x����k)le6�M�tf@�~:,�	�t}ݻ��-�o-�j�RQ|���j��G�.v�:�m<�yH4�]!{�J������A�� ���W���5�v��fSt�۰���'E���9	���f�G�_��4�Kua��f�3�e��a����m�_f顁�R.R�nN�£�u)���N[j�V[#�h�#��sk����Q����J�yV�FB�������nD=�\�d�n:�P�\���/�����ª�0U�0�l鶄(f=�ew�|��������߼��w�v��Ѻnq�F��L��'gе�JU�SΦ[�v�c�ri]N[�#�jw��m�q�nN
��t��1܄ڽf���cr��Me�,��v�g�]M��lKHH}��( ��M�q+l�W{��Ln�.�:|��n|���~�fז�!����p�瞕\��}P�N��
�љ>(��/vx�-����$Nj������*i�]���8��=�����O8�Z=%`�-���p�9FV�O;�s/o��u癇/���R"��;���T�QN���v�����׸�F��Ĥٕ��յ��K�˟-P����Z�kd��Y�B��|�Zp�&݇.ݣ�ٌ֛獛�S�1��5�o�5\a����=7λNW���k���#��e�IG�r��(٥������|�=�Ud���j������Ė[J�m=j�ڠ�*�b0��u��Yw� �١B����ْ�t�5�Fi��_����i��ٹ�n[�����d����7�)���=u��v
�b*{3Yܥԗu{���ё�]��t/\��&���EG��P��c�O��[8$'��M�;{K %^�~}��;��*�Q1ĶD)[��*�)53�xm��n�c&�3E�+�x]��8F/㾡��^0�۲'��g��V���f��O��+֝ާL�{N�6
N�@�U�����v���RM>��=+/;�n
�s��X����汹�h�s�f�"y��[N���t�UV{��;L<�Ӭ�;�淓��+e�N3�5Z����W�;�sNd�~��\���ߗ�mT�sh�xZ�!�M��j�-���:/t�oN
�G:/`ƨ�.����uQ>��l�"��֭o#9Vj�栦�#)�/�٭y���#2|V<�%\gI�]/���l��Y��cNY����J��5���A�O�Y������-����2ߊ�{�JLzi��57+;%��u��[OX��A��#��#5&6.c	3z�����9	�{4t$�Y���̉:ϒ�	��||um 䕹��T&h�b����%Z�{�Ȼ��Y&�����.��D����X�=i{/~��2<�-��axJ���O�7Ʉ�&�N�_�ŭQ�v��i��;}�VӃ!���b���E�э~���7;@K]�g�lF�Z:e;	��	���!��G�f'2��u%$�Þ�6��o\����<�H�\ͅM�J�L��a�h��
uD�{3og��j���_z�
�K�ú��q+	����l_P|���4^b��r�Y��z�M���|�OO�}���=A$�s�i�Go)�����or�s��c��2:��J�&�H�-!������{����R9n����]�'ݞ�2E>��V�8�t�Y$!p$l�L��w��Yz=��~�~��!���#f�y��z}�<�}�鄜�e�w��Mނ��q�j���q��Ϻ�-n�ڝ#,9�#74U��j��#[w׬�n�̓<��p4-0�އ�_K�s��]OsT
+�g-��� ��H��]��A�G�x��X�ԫi���G6�T����D��==�N��\w!$�X�8�������XKQ���x��k��Vy����m���JdFoq{�;8U�l� ㏁�;��u�[nj��w#�'����3ë��z��ߓ�w��Gb��ưHA�K�[Y�W'2��{�5�ӉM����pP�h�/�ѵ ���ty)0��v�����Q���W�owT�s^M)�!��k�<�����l���;\��cnw�>�.�g)4�oK����SI�m]�׷y�>�UYڅ$������ܝ��%\ec"ު�L���|���L�ʘ�og6�.5�U��07V��xsD>��������0[�K�K��w!,�R\�5�㻣<���m_��,cÔ¨v#{=.a���DC\؊2є�=a̬��s��nk).δ�w����a��X==�cp����pq��78]ſRcqw�n��:G�m4�o�//�Ciڳq�o]Ji4\���1���'tzm�oG9�-�)���G�����S@�F�,��\�4<yt�K^���O�o�準�]��ٴ"�gR�CI�|���{�UPu�c� ҥu��Y@��g�:.s�V��x��τ̒��mrWO+��%��&��ѻ�k*�J[��U�ɼ��^;C[[e�eQ�]0�m��ºe���[zC^�5����7���L�x���le{dDIUv�\�t�����Iپۦ�T�V�Omd�G��mT���j�p870�y�������*�d�����.�@R i��"3�Hkj�9���Z����a��3B�yvӧP�ڊhN�~��dw��L\En�}��p���
��d�����;�W�tn��v����)\Nɹr�a��"��s���3�s����c�gC�ݩ���45��7'x�'�������}�[�&f��Ľ̼�yYw"խ�3��i6'��]r9[ӄ%J���S�ʼ���>eTv_\i��w*��Ւ2iP�u�;Xr�y���ط��&�3Nk`���y�%��o��ߏ����3�L.��Pu�[�"��]fܤ�d��Mk�j�=�4u��ٛ�1���nt����Ȫ��<���nǧ<��[����|s
͔�_Z!{e26.�>J���TR{���Q�4r���q}�Ҕ׫^))�l��m���3*g+H)c.j�=���%ҋ6�϶M���)�<�!]�&��Q�ܼJ��ƻ�5˒�^1N�2�JpעA����|�l��X����t�0�xscUЌ�9n�+�f�m�[�}�N�T1�obAת�e'�ky+}�kglR¦b��%�{����}���.esVׄ���v��7�v.g��ݹv�#��KD�b-����'fזI�+�<9�wΑ��������s��Ǟ�K!�0�l�q�]W-~V+{I��|�IJ����=>����eč�=/W�d���%Bw��R�ܹ��a�duyd��1}���F�Fx׆��P�ei_�V�#��q���E�(U6�0��dL��$� n�#���	y���&�����K���c�
)Wq�n����v�M�}wѸ�(�q1��T���u6�[��~@�k|���{H���������t'nƖf�k��bo�ؘ�x�����т��QE� 4N��#�;��P�fх]#Y����� TR��T^ 9��5G������t��jT�B�wov#�"�m�!�]�ZZ���4Asd kr)�Cs�����]ޫ�~�:�)rrL6Ҕ�\��o;��ARlљf���̚i�"f�*�tm�6�D�9~�Z�ʬ(׼֧��݆�;ܯ�间��P��G�nn
�
�t�G�n+���w\g@��YL@x��n��L%G&��e�:������ۆ�	[�j}�@�Դ0E��E@u�Aa�WR*e�����8G<a먇V|����#7؀�j����	��=5ۊ��e�|��u��v�b�t�����42���~���l� 8��_E[����Y �����*{�It���<W�Ş��������OM-#u9�sϦ����|wH��Z���ϒ����u�N��tnPX+��xc��;1p
�V
}�#GUR�:!��N��$4D�H��ݧ(�nhњl+5�
�U$	a���اU(�s�N�艿���Bϣ���a�9޼]�8���vb�U���w�W�޾TEe����FW��z�s���B�m�O�=����7ݾ	t��^4(���)��
{/�B���ʉ.%G���4v�d��ц�<l9�B32x֗ft�|��&�P�SJ�A�[�,+�X�%,Uq*`q7\ܦ^w�.�Π��t̸���̘��'����{�伹*'�v/���;�&s%Y��Z������+t[gfr�,Y:�r��V(Z�+ޠo�	�]��D�w���Nז�uQRw�Sc���pq�`���˼ؕ�|?m�g����C���6&���B�u9�7BR���8�9�b�}�&��sϤ�0�[��Y|�Z���2ٗ"�|���sqǒ�
4��n'Cb�ˀm�wf��Vyg��,���ȃ�*�F�"{��*4M��E�C��X~���~�Ũ�|�'�^4Ur�v��3�Eƿg]�����E��R�f���!�;&zV�b�	к�B����Qt��<�5MrySYD�/(/!�C�D��ꃁjf�ԭi�ܯ�X�����U�ջ�(�'Uʤ��/�s�(:$u�wF㡲a��#CH�E�f�s�9�t׋=b6ns{>�S�?~M��ݤ9��[�����q��p�wG����@iLF>�1e�A�I�[��#YS�(v�L���~�^��p�`�8�gJ�����v�.��\jz��;�|쵏p�0n�tqG�;T���ApM�K�x����<oG	\۫5W����َ�]�:��z�7���ݻ7������?6�����g|Hug�Q{�>�W�]k!�ƫ��g*��ٖ��>���5��<���%��a�W"Z��.�E���W�������Ε��.<�gU�Oc��lm������b�uVF�5�1������k�q���ǖKټ_.ut����r=aԗq��M跍E��EO5:��A�n4��{���?{���.�����)�������h�����r����7=�'?Q��0�&Zu̩�p�y��Ie�gN���Ȟ(���O@��V]\'o�f7׉����:K4F��,�r�㈇�S��y��a����Qb���4�;�r�6Ws㞂$�o�V2SHV��5��(Q7Ν�R*\Tl�VdgiDt��jj!�'Z~OVb8 =�y��.�_S)'��
�t�����AWGf��rZ�Ơ9�*W����n=+پ��`��k�	���� ��4�E��z]�'{�<�GeK��V��f����ʢ6ڧ�;EBgŞy$BW�@�3h�x�x�QiŞ�o���}��YB`a̮�˜��8��Н��/��t1Ru���1"К������s��u��C���S�� lO�"B��Aq�/�x:��tE�y��g�D:6"d�*��Nh̖\t�ɼu���̿k�-���o�%�czLݑ1�ҙ,�,Gѡ��@�Y�������OH��k�*[bd�Z�N�]N]a�������s͹��h�2�ԃ���L
̋��tZ�P))	�眱[�t#����澀ڠݙ�n9���u8
`ѕr����V>A�ىK��&�T8��W��AE���KSw��F�ڬ������+��ae�fJ��b�� �$"y�[]%aJԵ�IR�Un�#a��I�b�4$��"��/+��v�(��@�Aa&K�Mr��J�/u�N+.(�Y������3T�Z�=d/��.�F�>'Bp&3��ݛ��܌\�v��6���.�4M۔�wĹ�)�T���<���H��٢P=#:�5"��3	�B���ݗ�k�"\;4��fg�-mv�&�q}��� 7�&�XV��"m���&M�K�0	V�d���RWFn�j�ʠ��1��G���|�On�z��#525�S�WdV��e��9cB��%L���j�U1j����̮��U���k�3���Γ3�Ҕ�< �S3��agr;:�l]/x�]H����5Wz���-�[�����(b����P&F��
��V��j�f�U�MCQ>�48�vGU��<8�;�|&������;G4����\��[Et�R���?�
:�� ���	K)��U�+&��дh�Y�u6���waki��<�\�Y�/#*\;�)}�˹J�rq��]G�
������#g67&R�ݷ�����5���Bj$��*��m��(9�݄�@uf�lo:+�,���K��%W|��{hI�+2��r�u����̜k��'ZM�g���6z(�k'�6,⤝n�?�7X/��#��'�{V�]߼fO2I�ܾ�&���Ę�^���+wYLQd�Gr��	�s�e���$2��xK}�d`��
��^�N�劼�[P���d>��4%e��Vn򌒍�h�)�c[������!0��F�#S��]e�`�ƣ����Y��f��W>;�t���Ԥ	��d�{e*�=yWV���<�EfiƢ�3ww��{rC�rq[��>H�l����s�_R�uلUA�wj]+�kgwcC��Z�V#�w:"��ꛏ��n��rs��Km�u�)�O�-A�ws�ö7"+%b=S�7y����C�{�� IܧV���E�Քő+
�&lg%x�Û��� ��O.�����to��8z�W���ͧ:nt��.�qSG���\�8�J�A�Zul畕��>�mӠ�#Z+V����B�J�L����  < ���Bݓ3���Al��@�`�Wo�r.�ΐu�: �g��pA:��T�\(HE�Ssb��)[�S6:�c�׭.���;Lq�+B�ܗp��OӍ�L�T����v�|��h/�Ӳ�%w��	p-=�v@��YJAR��<R�<��t6޲؜�_F+F��v�.g9�Vm��k
T讫��X��A/�%PH�J���*ե�ZU�h�>�J֖[O�2�V�m*�ʢ�a���4�8e�-F�*Eb����i[EAXV�5�����"�h�-sp�(�-��n2���f��1��Z��u�YPZ̥��L���"Źk�b��uK�kF�*.T���ֵEG�bڶ��m�Z-hUAK[Z�-̫kp[�%b�m�b�u�k�&f8��W*��Uim1�r�۬��t��u�Jc)�GZ�q��+R�Q�9�kV#h��j�+FT��E��b�t�q��ƣm��p�-s
�.2�-�U�X-VT�4��#�mU��ņ
1WV�k11�am*[ehRؕYU-�4�&�QZ�ˍmn��m-�V-s`X�*���
�-�U*�Y+�Z���&2�nd�mˉS,)�(���ڲ�+�h��ڔX��Cj�*�S�Z��5��[��N�{�R���S����]q����fg%ԣ)b�}��������9b��˵�j\�z���(��yc�5�Trv�g����)�>�.^��o��a�J����)�&�r�P[�"�;W;�=�.��X�w:D5�"�e��?�"��6��k��]�N�o U{u3ʵ��=�����m���1W�i��"�G,M��i�Vp:�m�&����w�������\�(��B��IXoͺ����zk�:�M�Le���q�-����N�U�_S��	�t�񵠾y75����[��x�8�S�q�l��W/&Bg"p�Zȿ�&�hy����پ�dvО��3��L- ��G:��03P�݌�ea�0��L)Y�dsN��P�k��P5`���3�>@V�_yM�^�H\�J�m��Y��"!>���Y*�\C�4l>�\)a^<��4�Ò^� ;�cB����o���"�o�{�O'ǎ�G�ǎ�;]��:Ynz�IX2�_P�-P�%�&���<�����y���}�ݚ���:�_�3���Ã�۞/�kR��$(h<�����=ջ8�攷���{s[���Nf���Hi�F����j��+{3iswjI���٩7�e�k����A���LJW��gG_��ͥ���Nvutٹ�ldesʂv� ×��7���u��}ˣ���ތ0޺k�)�J�V�C{+��1wH�Q��v:�u�&z���u�*S��1,�)_�w�쭵Ng�$c���Bڠ`=2�pp��{F"�>�m�@�S���}ү�1㛣�M㜁^)Wq�T����~�n�ؗׄdXIQyX��L�����Wva2H��It[�9s�FX��3�G��sh�NݍY�ƴ��;g��;�w��^s7�ױ]:A׊wJ���
!}���P��0��k3��/���uYm���Z��v�֢yV[�r��	��:mM�F�)���Ga߈���"{��	���מ��r3��4�A�<�MЎs��*��kW(�x��G����VC9�3�����B��#k�]��1�tD�j�h��8L�sp����E'��Ȟ�^�;ԓy�˞ܣt�\�t��q��~��~'�_E[�����ƺnfȳ�PB�V��Ս�!u4DF�C����*0�������L�#G���3��7�~�y�<y���7q��a,8)�h�v*2���%�)��;+ �V�u{e���E(��ep0�V.�N�X�-�dx�.��V3���َC�>
��N���½f�U����;�b�lx���b��ފ�{z��E�o%r�o&gT���fM{|�p;�]���noM�9��' ]9�~��]�AL۸��7���W<�,�-��9�[����W֮�oIXke?6)���[���y(���,focUW{C,��<��:w���0���,�����/���lJ+ܷ�P@C��)�;��݃����yWTE���T�=~Q~S�}
d��n�iY�@�s��z�����˥��w�I�����\W������򢈛hSJ�A�[�؜��B�J�&:��K�£*�fc.ث�pE@��ȡS/�囎�)[��s��湈O��߃}'��d<.������SRq�E{�Ѐj����/LW�����v��ȯJ�(�N3�����Fo_4�A����j:��s��H����m�נ�t�Xb(� ��7����T�!�ki[|�V]�#�Ű�q�f��6*Q����t�b}=+H�(�j�F�+ZP���1I[�ܚ�(��|s�y��/!�C��b⛪�L۩�����d��v��޹֫=n$���=~����lpGveU��Ɋˈ�qv<0��|��z���QGV�x~s�zC;�
��!/2h"�%wt�����%�w9���r���Qް@���ьKmP6�`�s\'|��dr������t������W:}��l�J��-u޹:��}X0یf�3]W�ޭ]z�&��KmKN��r��q�[C$��:��7�`n�3Ꞹu�u�i�tfȏwٖ���>�����(�=�t�:эKQz��@D��a�1uw�A<��g�cA^x>����̯1F?S�3اP�8Ů���]�~��M4$�P�G�f�z��.��>x�e�nmWt	wa��m���c������٥9^�5��=T=ٍ�>�:#��������՟Z�$Y����L{��t���Y�g!��U̹��4�ˋ���|�!ۊ�)����٠����(BK����!��N
xvoxFs�P�"/��3�US��@�%��Z���)Ȕxx���h��c�1�R��I7�j��bH�4 p�ư�5��E q��*p��Sp�՜p'/�FGl��(��]�v�{�I�Ё�X�|���4�h"��|w����3�.+�Q>M+E<�������}�7��SG�����=�\ ��xJiw�K���o�7ŋήz7��u������rzz6}!�y'}؍�Uw¬ <{�4�p�2�E#�ڵ�[]���(��nX�צ)+sT�I[U��7"�4�w�^~�ej}���� �YK�9	��r��X��K��+�rrY��v��֘�����B
��λ;��@�eٚ:s��gr��/��ݼR�¹�׫k���a����w=�;0��L+�5��#jڷ���ӟi�	Y�d�"�t�	�Kr��"���N�8��0���{;�J|�X>,�s�죒���A�'^-������X�1۽���}aj�T��=�X5��^��%�"��tE� �V3�r�ݨJV�f��ŷ�-�~���}�5g�����o��`OnИ�oJd��,E6���VhsYwz2����K��\�3�$8z�!���Ǐ����<�ϡg����u��L(�����H*�E-��4�\���1��&<�ݝ���5BګP�c��r;~�w�^3�~�7|U�-��@R�ս���{�ܥ9֙�b�Ps(�gʉ�č�z�=�֔�cb�$���/�ʢ9�]G��οPmm��Π��t��([0���vϢ����2��l���`���
4q�q��N��͑Q*��Ȱ�ZkR=��W��1�ݒʵ���F�����P���buޣ��D8��q֛�����ٞ�����F�=Y�+ls����0{<Aݶq��"!������pq!+vѲ;+��EU[�#w��I�s�5R��oE�t�vh�.d�&=o����ٚxu8����2���V�w�����y㺴o�6���9*P\���N-��E>g�ݠ�UrN��Z�P��q�F�Xc�n{D��)����B�"x+���7�a�fB���xeV�!�9���S^*RV*�($+����ϟ ;�WP����j9�H�t�&�UU�њ�Od$h:���K�K#����%`���XV(�Q@L˄��K}{E��{ɚ}L�6��j��#b��@y�ӣ������5�LL�!C�ŝaMs�Zx��1v&�.����f���}"�x�wX�b4յ@�xC�H�q:K��b %���`,�WW^hHmX%H� ��Q�o��J��� =9����n�ܾ�WfR�c���u��:gz�� ��q�w�h��h�o��S������ڄ� ��K.���鞮����M���S�q��W����F&e�2:ͣ
�F�12/9�٧f�u4+�&�a8�t�)�P��k!9o=k �WHL*��6�g�w���N\M�*��Z�w'sn���tCE�=���5 Ǳ���ε�ک���EtXh�6�m\O�˯%{2�XF�{.z��98k������UoX;Y�t�~� ��W?;�Q9��U(ǵ�����h�Ac&�5�7{u���q�7��J��[�����Q`zkG���K���l�2n�8y�Dw��#B!�
�2o[�uN���7�q��+nm(���!|���<�X��ݙ�v�'�>��IS���P} ���g�C�����ԠrO��<�w������-{r�ҽ�F�����������W�V�"|ڬ�A���:^�1m�sw�K;"!�,��~\�����6�C=�&���3��
�3|*�7R�q_��4��<I���5�&9'7����vٛ��t����#$l��Hy��d�C��ӛٞ��5�[�^ ��^��XC���1T��Xke?6)�@{e�{n��S�sL��i2�̘��5��[/;��r�aE�}uJA��B�\h;A_���Z�ڮ��F�������e8:�3Ψ�c'���D.�$�]�C��/�Q�Uۧk�*<>�5�L�ݽ����!|(�#1<_ǅ�F�|��%l��y4�<�*���NA���mQ{��)p+���(O�(q��P�����u	J�ftw�1i�X� n�c۫Ǟ^<������Q�Ez�&N
�� ���}�@t[�=l�ˤ�aГ�ӿ ��)*�G�@���+g �����{�k��[g��B�(��U�ZS!P��YlDu�Y�e��=��ӻM�;2F��[~���mON}a�X�R���݈:��Qܵ� i�F�żᗟhO�:��o�SJ̋.�B��K��O!η�<�$��7�ivu��3�ll<�pK۶Bx&Y@=�G��� ��6������ٺ)h���Żz��{7��n�0�t��Iݸ��6Ȱ��J6�ܖ�$B2N���i85�鞥,��C��c��$svNzP�!Òb�uA��3~�?Mͼ��@m�^���Dsd�y]�W����E���S�
��2F`��$Pn\DSH�E�0p�s�9�5h�K��|�L���_RJ|�(,׃.��-U�f
��g�f}�����<<){����&�(��۞�s��ȴ��+���`��Az��X�O˹B�U���=��[�"��{5��GG3�u{cu�`��Ռ�5�"�����^��|*R��\=i`��}Osa��^���u���1���qQ�G�3�7Tw�,v:!��5����xTW+C'^�[�GU��cM�\CɴTXUU��U{^y;�F�緱�_u�vyH�t3�.0����w�Aכ��<�%n�;L��ch8�."$w:�T̸p��@�Inz�S�������u��:��4��U�nK��b��U�!�T=�EFʴ�sx�\��%J�G�ҙ����IW�=�/�^��b-�(,��{h���zY��̷}�J�ډ1�=���ܱ|{jNwxynA\�ۆ��
UF�tEKK�QLK�i.�<읱�n��D���.ѭ��W�n��g*�@pyK��u7��*�ƿ-�������i���h�:�Q0B5	�}ꙁ�BHiO�;/���3�.+��Lt&�uUr^��p�.�p�EB��b6N��^D�N����'���/�қ�G�b� K({1����͙��I��;И�P�Y���Pp-�eSRH�AEI���E�U�ЏX�bN���Pw��/.�!\����
Su�-�q0cd���^!.2#���!]��Y3,*6�%�wM���A�̕n��5�7M��z|,xX�������g�و	9�nv9�����췉5偞�<�4�5y�+FT���Vk�i_Ñ|\:"⛪�cr#r�<��V.OQ�Z�Z=y���Uy�����ܔ͍�0$v�	�zS%�.X�pXR8]���mx�n�a5 �y��f�������k���e���cݫYc��Z�+}�G^�g*a�95^D����4y��	����ѡ�H}�2g��L<,�Yf�?J5�-�k.4pf�]��(Z�J��V���d�mm�k�6A��;��z�WU�k|J^�WYagM%���Y����E!�����IDb��u|�uQvR;�NcO]�1�WRzI�(�Π��V0���	�+_A}���:+;�8z�뾌|� M<�)���i�X;ת�`(ae6��R��sh�gV�j�=�\֝����MmHqB:J�cy�G<}u��^���Ѯs�C����ƊΗRg�s�mƝ���\�&�|�-�bzh(�31�N����*$r�d4�s*mvmS���HY�*'�ޣq����=�� >5�(@ZA�:�Q��4�q��8㋇d����P"����/Q|��`�^���G���#a�יи�[�Z���(i��*PQ���M����_,Z��W���+��)a�>\��j���U{�\�d�D{��OA�U5UbN&U�繦�5�Cf�t�C�Ui��,�6'�ԕ�e����1��l������-��)EkS1*a�CmT���i��k�rx_�,'�@����Vk�b���m�ݽ�=�u�T�h�+ט%��l���#�xձ�Z�b�=4�����
�!L��V�K�wmE�'�v��՟Z'�V?S"�J��9���t�;v'=�BYz��W.�Z��Q���%�;D��\��l�F*}O�ɰ(:UB3��o�[�\�uA���;t�<[w��'0:(��E��h�r�����:c�ö/zD��Vd��#CgjU�cNP��^�*��]p�<%l�W{�9W:�(f�-���l�O#˜F�]�U�׳.Έ�-Y�s�|���Wm�[��`�ȭ�nRI.�<gs��B��K�G��󲼝���{_�j�A%+�"Ö0��[�����WL
<�X��^
�#JN��1��^�iֺ��rh&�Z6g:Ŋ;V�6���:Z���w4���+����M�X�K)��P��޻ȳ��CXN��9̺=�i�T�M����Y��k����Ћ~w�w��̔skBa�fLGܥ��Z6i�%��0壑T��y����m��wa@3Ty]��-���@�4l烑Bㆃ:QweuۨQ:,�zɪ/�vJp�}�)ç.ԓ2�H�L�gpd�v;̫�[��r};-P�8l�2���5�U���ͭ�5ZB��Ұ0����-�ԔK7�䲯6��3�}i���Bķ�W�)b��pK��u������3�n$2��m��#�a�����S�s�*<y#w���UK���ӓX�R�l}V�זD&��]\wy��q�Y���d���s��`㖞��7���bm3��f
�����X{���{U*Q-�l���
?1ղX/��Zl�l�}��3dP�Ŭ>6��ʭ�ֻL�q����b�$GP�Xz��%hN�M��{]���V���<�ȼ���rs;4��i�8c��w|x7�A����ɼ��BfWv�%�/	�i���v�����b��ZBL4��૦+&���ApqiK�J�!���ΦN-q����	�G�p�pe`:]u�2�]�y+a��M'���Yz��\���Lqd���G�d8���p��p4�v��Q�\J��;(� _�D��\\����B��C����\J�ٶ�b"��F�-�r�����:�Sh�3A�hY���Q�RK��\v���8���Uč-9��O�Rn��;��.�)����g�u��iԀ��eNx:GQ��U�P=�ԽS��ob�<�g�A�_3���S������kG��>Ҷ�e�[T�̸Ju� �����J5�4`Nb�6��7l��9�'�� �5nk����:Y唻0�8_:���qS�أ-A��&��ii`�6�k�]0�2�1YʖNjj�)��l��+�s��]=/��j�,�Ҫ�*
+s@D8�`�ϐ�	�z.��m`��>��%N��ˮ��Ag���H򱥱�|]�Э^V�KSk9:��`b��G��[�ep��;�U�T<���03�T޹��wx�*�D�\qj�rM]��r\��ET*�>=�'&)���\����6{��a���9e2gc�0V�4�s�{+�0��򉇗�I�S���1��R�fj�Yn��+*%j(�Z�%�R�B��ň�UPX�A�h�s+l��*�L�m��e¶�Rъ���Z�k�X�JȰ�J+mF��EFQ�ˆ��
)+��hTPUTT\�ƋJ�e��GM���lƘ�k�-�"Ŵ�TFjأ�6]e�[@�KZV�(�e��+PU�[lm���`�P��[j�crх[KmZ�U+j��a������TQZ%�ZʍiQ�ʥ��p�R���[iZ������N.R�-��kUE�KQU+32���(��A��kj-Zڔ�,��q���lƨ�V��c��Zʺ�9s1ժ�dЬ�i.�&[+R�*Z��1��-A�P�L��hQ�U*��ha�(���*媍�����P�5U2�Z6�ұ�.��Z��X5*i��Yrڴ�V�.e��D�.U�MS0�Zѵ��f�"⭖�Z&eŕ����:Ebe(�Z�9���.f�iB��V���3-�Me��d�i��-���e��󔶝��gv]MU�$�X��b]�1�-c�LξyK �����2Rwd�[���V��峨%�E��{��\�P0���4O����Ф�-�``S�����:;P�C��S�cu� ��1+͞wFpM^���v7%�c#<�1H�J�I���B4�c�C�m|�ϯx�5D[����VH�3}<Jb�<�(]�浐T�:<<�jHV �lQ[Bb���0ҡ�b�nS���Ժ���^�J�6#�d� �8�j��K�9b,s�u6�n%�=+:���p]� �[��Ú�
�U\u�`P׳<ج��`y۠� �j�)�dV��g��㜩�ɼy�]:�MA0�����[UXug|m5]t#�����xJ�7�9���&����}9;�w}F9����Z��5�2r(K�g��F������ii#�����.�T���S�7'o>��&�^���>庅z���>�	��D��;�R��*"FH��
�Sy9S��w[�N.Բ�fE3��7�>�Rݪ��w�,W:�H�Z���\����'AI�ٚ�7�	����2^��nG2-T�^x:w�̨�QmmTk�D(��[��U���E�,�v)�-p�p�V~��N�qyr��{���f)�YU�,[�<KS�����Q.p�/3�_Vn�ܒ>S��i���g6�����S
�8n��c�7u��o#����p�L�\z����]����3�)���G4�wp�$)��%]D��v]��S ��A+
z�����Tl�`[�l�����6������j b��(��F�H�F����|��%l��&��̦G�)<��:����T��~����z"`��R$��+�n:�+q�΃��?e�o�����l�[�{��Gg^��d^�Dw��d+�5+�����S��;�8p̞b��pӘ�z��4�;wg�oH�~�.�{v�O�(=���Q=EF�:�PC�ͺ�0^���M�}��j:??�ءk����Pe�T���dXSb��sr[�!'`�1��t�R�/SU�ɣ\�t�$*;
ru�^u��D��s!��䧚�kL.婭��ݹ;��ۆp�(��
2�]�8��ݻwDt&Lsr�!�f�Y�8a��>�ݽ��B��}��?�J�uK��˦��e����p몣�P�E�p���Cݤ����̴!e�lC�����y]��{�cAZ���L�{��7Z�W����w�$�9�m�����������*X~�Dxe�Q��J����Y$v�;G�Oh�̮�s�fCf�wo4[<�	A��ޱ@��Fh�1u�J�ɲ:zͮ��)N��Y������)�ɼ��wC�l����Ѣ\4�T5L\�	��3��t]UT^��j�Z@���G �;T��}�.�i�t�^!Eecw�������L��;ϫ��SCڪ���}5�=X2,C[�QW΁��C�(@�!P�������k�����a�ȋ/J���EU^׉ߟ^�d���lf�'+�EAI3�	h��n�=�K��8>�����]B mo:�p*�p��@�Inz�Z���9Vu�˹oj��Z��n$�R�E���e�ˀ`.9�5����B(d�r��&��#���Jգ1r�������m�����Pl���D��h׻�F���T���/�V�L�'�{;�K�ﻬ,��+I�x�N\�ODHo�	M.�>i}���ۻr8�� �n��J��6z�U�ٮ��z: �Pp0}�.�,m d�(��4�R&:���u���W$;=;��.��	'���Bӭ�Fp���Ł'h���Śy$BV��!Q��s��kb�UЇ
�7Aq������ܘR�/��e���OD"���`�p�Ls���[Y�A^��9�����ޣ�S���G��t_Py�4��ӭ�[�)��f�w(�f�U�{	=�\�����u����zp�н�S[�����:K[3���$_�/�ln
xN���	��^Ն��{���ZR���a�ޙ͢�E�7t�$�|߲������� tM�HU�A�T�%�:��tF�r��V����uR�vjk(�h$>��^|��չ�;-gx0]F�Ә�,߰[��7�6�ܵz���N�\!�E��>F���y���<>"a��\�f��y�x=�JL�٠x��㓷�+=vj��M�M#@�uΑ�9 ���=�1H{ٟ3�|�3&(��ںٍ�ʌ�4r7wсs��4W��Ҁ�i��o��|AZ��5�80�ԩv�&;7flwmo(s4ԅ#��67�Ds��Q��ͬ��Z:�vX<__N*�Tj�j]���L,=�܍�y���F[�
ę
({LÆ�yy���b��>�3�d��;{�N+ԫ۫�=���1h��V�ƪ���g�/�ag]�9�4�q�׽�j�SD_6�w���Q6�]A���/�X�J������y�� +l���oJ��ǽս�P�%Uw���KˮJp:u�t_�
V}��ȗC�M�!\Ԓ��������u	4&7���t����!���Wo�]+(^Sm��p q����Ҭ9^�祚���Z=���Q����K<I��Ҟ�30V�r>����h$5�q�`k���_R�_dԈ��:��M��]5rJv�Xb�ssR�;�_B̘��D�m��+�8Xț��Z̀��i��e�K�Cf��Jy[
3ѥ��yz��(p%�	���T��c�{��8ˮ�����w�L:��ک}D�S�pz�s��SJ wW�R�t�q=�q�*�h�⮁��\f!���+dT!�)��t#
���zi`��mE����!��
���%0��
�<�w�[h��X��`)/�?����
���8�1\�>�5v��w�����b���DS��D� ��'Q�hB�xL%�څLE��}S�i��b*��p��7���ܗ5��lH��#0L���B?s���b�^k�R�ɿOYW���9�̛1�d�Fb�uİ�9�u'��xѺ�s���5�0:=������K�O7/;�6�"��=F
�v�+������2ɚN�E���7B3�k�+��{�]���{��-��|��-,m��=�HVpD�
�뻁~�Uܯ��W{�ڨ���Z<����!���ywTr,%_�c��#N��]�#L����ԅ�ퟄ���J�w%�[�=�'��ʕ�sy��1��SVƜ�"}�����ۘqa��{9�H/�����A;&JGZ*��(o7�:��Ŵ�v!��r�f�s��Uv�#Τ����P,������M�;pю$�ەt�l�s�9�⬤)��.b�=[�굜��&�$˻&V�>��VU��z�t�ԧ��]B����{A_����bR��^_*������UFgQ�3�?=uqb�&/����=����]��|�N���{�?f{"8��7ކ�p��B�6�e	UQ��{���,o��a�����M�	a��)�@�o�Fv�5�i44��g;"3_��"@�L�RR9�j���:w�̨�P�����j��0�WYŖrU������vr����1��^ui7���hc��0J����8���~������m�SR��RQ%���$E�:�FW�"��2�C���TQkhh&��_FcR2Ll�7i캒��R��D�~n�y�Z�R�^�T�[�W�]��3��\F��d5���K�<���ݶ&��q��&�1	q���AXC��ŏ��?������H4=�,·S��j��r�!��v7t6*ܸ���!��^X=�����F���tRvl�q�OA����X~���\XS+�{de��z�.m�aM��o�9�-�H�uc{��s���F�u(�B�Y�CH�� �~�WO<��X$݌,�^���<^]��n;����j��v�$]d��/a�J�om#=l0�`Ʒ�
�r{��LW8�B��jagm�
�A�Y|�)�g*����N+:��k�B��8��l9�	�=&�霃��P#]]a!W�v
�t��!�tL\Pn�8�u;�qf�"�/J�oݜ�:�L��W�%�V����C~4%��̵�3�yx��ʰ��j�
�31�=�N]Iuy��)a�x���k���k�pO�-U�W^g�fUn.��E��cCgM�-�'�!�+�����]4L8Q��=���Kխ2���{���mU�T����(Ԥ�m�YuYR+Hy�R�a��5V2k�2F�b�m#�R��*�;]�ӝ�(\�c��[T�E���d^��q�������ݛ�ް��>��!�'��a�����{7�ݖ�n�S=Ć0��/K��\� �����ߚ/�VD��C�e0����55��/Ѓ��G%�L֫�ׁ��bMBOw����UNg��@�Inz���gZ�[�p�M���JN;�ؔl��ˉ��`>>B;MĲ�r���85ʜ6{�ӝ�����{��:�Z�_��7�^�ħ���t9C���)"8�HzJ������p�Xq�ǵ��(���*T��W^:	�^����f��S�V��FFw7���&tCz�K"��]��n�F�Z`Jz�<)��$�<)��2ל�Z{;b$� ��Ί�k�9�/uT=���/��ɳQޜ�s���)O���7sPS�����mG��"z5ӑs��� �g`tKiXj�+	�t�*I�=4��4�������ŝI�<����zn��`�_?Qbi�o�����c��:4S�{�x�i�\�M���A@��4�n?��N�v#�^j�j�O"�gcb��	��۞�9N盨��[V�b�����O$�H$�E�L�q��^�\ڸ��ӡH��H.�P�
���*s���3���@�[��
�����{�MI�
�Un��yJ$C��4��z��
�7�!oH|{�e�/!��r�u��2�0����|VI��{�������������W�w�]���]�3Q�1��UmCoOt��Q��G��,���ё0��o��3>��Re����%,�z۠�.ɻ���ӷZ�����5�|ɤ刦��Z�"4)�'�ԟs4,�ڛQ+2c7��;��^�k�Zx�=.2�j�E�o;���b��5b#ZG,O9�2�"�u����ҭ�l;v�0�6�v����b�r�P�k�RP����΢9�]G�������]UBr��h�Xki��[��vqv4�"L��FdP�����0R|��ڢ�ُ��G�,���7��M�۾�F������:Q���PF(+_\I֓� �1��>
"���vU`٩M�+5�:�����H͔C{��lJ˝K	����<��k��R'.|�oh+L�6{����a�%����?�g��J��%�]��5�u���q��.�t�XjFj��zg�]�n�y�ly�}MkQ�\,Llk���Xz�� TP��h�tx�D���}�6\��J�~s���%TpdC��Dۺm�N�<��	ˁ:m��Õ=��������������ЦS��8��L��b4��C���K�K#����%`��brs)�cetgNL�tdlW�ga<���ut1�-N\a��~=��֓�D\\m<ѻ-����-�Uo�EW�*3]5w�eq�	M��]���=��<j�����sy�!D��������B�vy r�U�w:�(�ڦ9�R�〩�L��q�K����j�dR�&}1�R>��ei��@w@���+@���1�`�&!�3VT��J�u:�YSYGn-��P_��Fӷcr\�y���n*(Ɇ��B�畨���Rw���C:��k�����*��(p@�~έ�c�h sv�i��V��_Ě�D��K��cJr��l�xC�%)kޫI�6s}2�����R��Fbɥ�4dpwZ��z)���Uo�粙N�sy�\��>j�J.t)�Ug�N��w%Js�Ԯ��4F�5��'\K���(]�5���V[f}�4k�(`��=.�͏]u�������W���{�e�z+�����Ĥ��5 ǐ}�,E�u�����q'wWb�Lѝ}I'���� #�졢�>���
��nrϼ�W{��{��l��n�|����6L�Y��GV����mTa՝�un:�#����@q�'�-�����}+�v��lS��DCjn����.DG9gz�F�6@��]���p��c�W�3\C�����i�o]\�0�����r����s�(����P=�3O^����0E\(i��YZ�������ώ���5�C�@л�V�Ә�
���r}���[ug�9Ɉ�c)�H��b#��[/�yʌ�����DT��}�,� ����'A�Y�C�Q�F�E�	��b8v���Wt����dFZyQ��&��y���f9"����T�i� wN��{���aqQWʊ"o�hpxg]�(&=�w�g�)>�A<]���������u�ijl�e��Y�ST���tZ�.���[�"t.�]tJ��a�D���?��i�䫊V�35�Ϊ��4>�R�e�f�̀�K\-ꝻzD@��g�:����0^e[׹��;�SMp�3�Xz�<�
j%&�״4�>��Mi�5��-}�Gʌ��U+�7��pj��ZZ����K��7��w�TԶظ�e�=!�{�2k�pF�/�1�P�fr�p�@bPe�n��<�`�ׂ;&�_�w�]�;����:f�s�b�^"�. w_J{��U��Ngq��(�|��:<��'/�F����w�N�3TڔJ�%�Ա��ԑf�u �ϹV��Gn�ϵ��y��J�7]��Gk��ԝ��̨X��ә�Lg.�q���]٭�W5ga1)Ĭ�.����dp'�<6_h�/�ޏ���S����qAS��J1[���Է;����˪ZF�Vz���l#�9��3�שf�R�h��
X��̾����K�`���n�eHv���9�y���P��.��Ǧ*����|ˑf\�B�;R�ca6B��Yt ��U76��V�̧��0�o���A�{[y�	�֦U�H��]wE�Z`Cl��2�5mr���f��w)-��v7��h�&�J�yyaly[JF܁R;|7��}鮨�x��5�1BH�B{�.�]͇����]��+%�D�Ȟup�h��,�m��R:z��{[!;0�J���f��8%Դ�D��v�-w���Q��6fA���\�yq9ץX�ٓ4L��=��J1R�g�<)�*\ͦՉ�����:��i7l�}݇�g`�f����W�S��Lq�X%�$�ǽ�F�a�Jd�U�.l�^#9Cm[ұޱ*؛k��Wז�LX��q��7��gK��]$�����1Q�͝��.N4g8�`'j���+����m���:�A�9����ogQY��i��_Jns�B=�J^ӽ܉�k3:
�(ΔƜ=B1ۨ�Nל�:�툆�.��7��zՊ�T�f��$=]���y�n��ک����f�+"]�Kyّ���m�wP;iРxNg�S�7�<�0ˈ�ժ�uS���^`9�ᥝSy�xO7B;SgL̂��:3[x8�"�}�].�;�p����,��9ua%�"����U���m��P���(��n�M|2�(u`��yw>�ebAT�K\^�
�VpM�R�oQ�J|����:���L>����W,�aXt��`��]��oJ׋�P�pS�[����;��R�)�w��uȶ�pTv%���9VN��(
;SJ��,>�dv�1!��!J��"7/���GP��U.E��k�;˔X��*9w�L��͛7��J�'<Dq�������q}�o���Ѡ�>*w8�`;-ܹNf	Ԇ��w�z�A�<����8�h]�EB�A�XW(��Ks%�հ�t���fZU[
)-kh�̵J����!KQq�*�����eQ*�i�Ӭ��k���+��D��UU++mh�V�P�t�G��h�kr�r�թ�������6�ժ�Tj����)���Z�T��FT�q�)�EG
ۤ��TF�eIV5*]9���i�ijU�U�����KB�UF��V��2�1TQĶ���0F��Z�(�3Fd]e�]&
:�7�h�q*c�R�S���*[B�1��.%QC-kUm���+�V���,��İ�LV�,��U]Z�����(c+%��1U�KkZi�Dt���NdZ���f��iX��l��F�����Dcj����E*\�b�DQQ����ne`�b�m����j�R���Zf�	u�cj�%EVѴjQk)iZ�U�R���c̺޿u>����#�SwS�4΢�;����9�����;4�ݒr�g-�7���@R�N�)]z�!��z�-�fC��8A�},n��Dea[�X�%�r��)Os��q��n0<���j�0��UrZL�ب�_�L@�S�6}����RԈ�(�8*�h��������܎�����b篣c�+)T0{6�8�N3����e�%�R!�T�od�j�����[s��d�8�ѯ�Ϻ<�ʐ��V~�}�s������Pe��ݸ��6ȿ)�R�f��sBY�r1��}���bsӜE�5B�	
�Ӱ�P�렼�Y�.����(�֛�q��K��ޣ���=Sso��.1��j�[��;�Uۘ�9���$?���7�^]��M�K4�0�ҁ�y����1@�v<5�82���^�wtj���׮�g��;a-9U4!Q 0ڨ����\d��>�^�;�"Q�w�Th%
�������Twf���a��4�qh����g�(�CGhݒ:
W�� �1$��S��8�Z���oG���ub���_�I���̪��s�chC�v!��^f���f���o�zI0�1=���?��9��ap���:�T]����@{׎̼�Ax꘣B��:-A�Eȵ��x�t;4�:w��>W�j[��tM@��n�]0̺��6P�A:�;{�Lv7��u,%-C0o<�ɠ��ot��q1s�l3�Х�}T��l��0���z\��T���*��-W�~��˾���,1��9��]�,D�kH��G�+S��f؀�iDGs�g�U8pɘ��c�dÍ}��b9s9�T�����ݪ�N煺ؔa8���@{�����K�u�Y�ol��4;ޒ_l掷h_cPWJ��z{��X�~^C�(%��"�_Ȇ��#�eZlk��'U�U.N&U���gW.+�Q!4�<FFqZM�ǂr�"O�n�E��Yi�OA�&$��N1U��Ѹ��n)�X����=�����"�!,M8=�q�ˣzP��~.m3Т��	;ݹ�r�~�_g�x��KmC<�^C	2Fy<פWFo=E�����~2!��ݡ�q�A�7��E޾��J|�_�Ŗo���Q\�>������N���3��@�~������c�N��l@V�`�f����ry��M�N�Z�t�tgȽ/��jy)�+��<�	���!�<\��V��<���Dlک�z�U���}�!ۋ=��rWD*���L��{c<f���wo6��cKo��Iq�G��v�D-S����Ỗ�N\e��Y��{G�y��.*�1^��rԧgbyt�,٣����p�nq��5�N�������!)<�j�R�2�3��vb�f�ü��g�!�d^��#"(s��F}��<>"a��\�g�elu�AJ5s�k���JOQ�n��5�>��6�����NX�i���#|� �wS�z�r�G+�2D6j�u���5���(�*/J��2jˋ���Qi�yM&� ��nR��.JA�4U������i:�5�-R�<7���C���
��9���]G��ΰ�Dv��B�Ҍ�-f·{��3��P&�T<�2���M\��̜�'�E����SAE��aƳ{O����o������ʅ�<�ɑkզ�`S�5q�t�vt�X@hb�t�Ǚ%ƹ��gT�I�4�Ȑ�ܤB�55B�㕦��;%pgOF�Έ�Z�!�o�I�7ٕ��H�SǶ"�r9j�9�N���S,R���r%�U6��P�_B�7ݨ~}���h��<�Θ������}��L�!�秡4Ul(�����$B4foL���s�:�4��Ηqw84C/(u�*�:Ixw_ѡ���SP�U/P�q�P�e8���{���
�^�j弧�1rP҈ۉ����٬4i[B������>ɂ������,��Y�g���l�W�p�~�ᙺ��A�����G`��!}u87J��q�U(�a+�U���'r''R�(ѭ���ΰ9ҍD�J�}!�����U<9�YdV犭��3]<��eq����]���S��OmZ/�θ�ۋqSZo�9�'.���j5��N'Iw�b (�����TI���?S �]ʪ��l�~��l�6yugM���Hyx���&��(�N&!�b VFx�GY�`�.��כ����=�9�|��D�wo�C��_��F�v�n.kؑ1�E;�@b�xQ+7�
+�"X�E,������ltu�i~�/�lTo���y@�}.�sZ�*n�U5$(�-�-u�ɯ'yxt�OX�b�D���2�;����Y3�:q��n����[�*4fOL8���#^�jޥ���p]�υy�q�Y�5���w�ڪ!Ӑ� �)�U\�!�v�5�<��[AZ�Үό�}�ǫ��e�PU����v㮔#��zO~A���:��;���t+����? e{��Q��@�ϕ��j�\��n��d��$���
RU׸\jz�W��U��3���\�t>;�LXNvN����������I�L��m�$;�{륕b㫝��d�vy��{��-��c�]����#U���H觺";Vs��ߢ+}r��_@CF{�i��uq��hu�S9��٥�����s�}��b�����M��S�.�=�B�"��T/�s��t�;S��psilNA��p�vE+���>�R����qpվyѱ��;��
2ES���ѬEt5Z2U>\욺��1Ӫ�@OLC���Q���PJG2-T�^x;�3�P�~�e��e�j��o�2x�oh�����+�j����P�ui7����]�P���ϡ���"������mK��WݹiQ�U��8�
�
�%ں��H����l���B�T����nvD)�[�3�D_���,eV����w,B��U��C�����.껽��q�Xc�`'�='�Ha�����85�@��Bu��g<�N��Ș���,����ybpUR��x��f���k�_�GmdP);P�|	�v7��^�./j����m����.�nV���{�kC�.v	,�7r�|z0��e����8��6�F��6>�Us]�ռ�,`�Tܞ��ρ;&T�"���$*��p99�-C��`�$@�d�nO�$��m/9}V*��y�r�%�c��8�h�Wp�W૝nd��;ĉC{�^���q�%�EvMU0�� �2�T��WT���J�Vu)WF�"}�_�B/��^8R�V�+.�ȟ��u<��#=v��"_�6�^��t�}��}2�ƙ*	�^l_u	VV��\'^���KC��7��%>��q3��ɒ�����Ξ�;/q��v/t�=⁲������|vP��v<t�x��j�p��� {��3w��+��l�
�p�*����p����09ԇ�#k�\���8��K`��s˕�ۻ<��ޘ̙�9H��)ѷ�hՖ�����(��dNa�h<c3K�X�o�R5�P�^��l%��쾾��q�C�-��:��E�ݪ��tm�.�)�[ӛ[{��5sGA� >#��uZl
<ɊTD���qs�\�*��<	Ͻ���vD���� �,ž��%%���5-���ĸ�YZ���6���n���o��{5��[髻�OT)![����U����9�\eV.PK@�!�@B;�4�r�/v�Pj�K��+7}{���i����y+�b�}�y{K��\X��%�������r4��ZVu޺��i
;c"�Ŷ.��.\V��SJ��
Fq���x�\�	����`�ߦN{}���n5'SK��M��.9���tvU՞��M���2�d�HZ�n�sLI�j�g]Xi����L]�QfA�������=���O{���D�\Ӗ�w.�g;Z��}P=ܹw�}R�ǁֆ��n��ʮ��]-���a!�r>�}����(gXՎ�R�Ia��ž(�7v�A�P�S^1�[�'a�{w�v!7#C�DH=+���ƁF�I���`�´��#k�ո��I�*9�t�/�>:V�i�Sw�(��"�"8��P���v0���ܸ)O��Ŗp*I����;����M���o�@��������$T;'�%���QZ���S�^��O�\g�GhI.�곆r�9�q����n�n�[������ !N�RW�ܔ�3]=;lt�8z��̞0�Bb�ܦK8\��42�Z5`o�gRHxw8{-|0礬�R��:���^m����[4����o�c��I��2[S�BS�s��}Z��%��3}���>�qӺ�ּ"���FPɫ*/y��b�Qi�yM�����'�}�!iW����Q���P�<h1[C�`"bNݎ��C�/����zn_ج�����jl^�+<I��|�ڿOYKo��������i�s��k�]~Ґ3n&B��I��U��XުP��.)��L��s����ȹC��ճ���iug�m�zD��=�^�����jp�s��0�22-�&�.+ �;޿B&�=H��EBW,���\]PWL�����x[�g�pnp�^����]q��V��u�B�X��Uc�_N7,%͜+\�jt����xE�V/8�QV@Y4ÝZ�Ipޜ}wZ8��ނ*�Z�V<�&=SL�&jj���+Mi�jvJ�"��1�s�%��R�9�3f��Ҩ;|θ���>�N�`!�*��.T�{�ޟWyxR�)��K�h�^e6<)�K۹�t�F�h�K4Ǩ��hR�w���e3I�l�R���*�g�c tF�j�v�����*j���!�����24��sDhʾT��jj�ר�G`�s��=ż��T2��C/`L��tUmf�/���e2�ׄ�ֆ�]H��)��G���w�����S���t��e88K�=�@~���s��=:�?S �܆���ʹU��{٪�9V_��@�8��c�b_]�Ϣ�J��Ɖ��$"#@��|���6��o��Ӹ2���&6�;P�#�8E͢�:�汑��
�0�����Ca��������4��_NT�/.kȍ�Y�aWH�f+��%�9G>�m�k ⬷F�5�m�];eo>Kө�ݣY���7�i���xW���7��N���{����I*���ˬ����5ظe��4u:�|R���BBŇ�l�R�<��K����j9Hx��v��c�ű!���#���U�[.���`%�ty�GE���<��4���)N���f�#��2��g"�g��~�������uju��nS��(���b�z�l���8-}A.���c=��r�:�y��^�DfS<+Ϊ㮳>
�Y��T�s�h�JD3����H��D����w\Cd5u�������q��C��x1b��|w*�*T��_=я#�s��e]��k��gK_�U�U��DD�� �A��\�z�t�ԧ�����;�;U���"�x&0�X-PJL�#c�O3���\�w���"bӝ�������.)���t����h7�̀s�t�����R:fV9B\5o�tlf�؝!E�J/!�C'Iֻ�C�qs?D�#n�T
�1��J"ry��R9���\�����;ړj��;���ނ�$�b�5��)�tV:�e{Lg�W:���y�ɾ�tB��$-�;�\����x�������G�ǆ#�y�"�. O���Tg�أL�s�e��:��S5mY˪�2��� �m�c�)zFi�Wd�
J_�\M�=�3���,l$��O;���U����Z���8�:�@�}�&��p>��~f���%�5�j���ռ�B��2�v�\�4�,6۾�}zl&�:���H��de�G���37,t���{:-�@9��J�zC��pp�z���x����֝N�{�HܼCR?s�.���z%���aR�w�E^H��Ӑ��oH�[� y.��i'><>�n��75ji8���t6([� Խ�D`OEK/I��]8����Y2��޾Cj�#\f"�vv;G�_S�р��e���ۏYsl�42q�a����z��)�>��TG}uAP��1>����XH\v�t��Y8�>�7b/����x��_��ׅO���kL.�tK�k�q��vX�_�Ƅn��6��T�%YR�k�/j6��H�p��.Ī�@�|��z���`��X/���X����c]r�����ݜ��gu���b��D>�1.�����s�r'��X*^���x��Fvңګ��B�7��tl�hՂ�>+,k�0(C�(����(���խ����G<xT�y@nU�u���+�ub���_�H=X2/���TWM��F�7�՚�|����E��XF���ʭL
)0��/K����qUW�瓿4e}O��(֗jw��]���}�orٮ�%ѕ����@,4��-p2á��ظ�'��k߯HIO��$ I?�@�$���$ I,	!I��IO�BH@��	!I��IO���$��H@�����$��$�	&�H@�d	!Id	!I�HIO�BH@�RB���$�܄��$��$�	'�B���PVI��G��^�Ec���X���y�d���o���o��PP�(P� H @�U P(   �@T
�� P�mIQ*U))*����BDHJU	(%B�J
(R�D""�HU P 7��!JJ�A% �@��%J���RP�H�BPUDE	E)UIU	(��'ݝR!U  v���5X��%`)55R�[Kj ��4�U�Z�&m �R�D�A���U� इX4m��� �E��0ړjՐ`�&LٔTh�I��֍�ST�J�"D�M� �ѫm1��,�̬��P@TZV �2�R���)#e�`�Vej��T�m�U$$K� �) ��Pj�-�$����� AE�p�P w�( �ܰ�P  QB�Ņ QuT�����L�R� (��� ��Y�KUV��k@����٠U6�%6P�lET&�V*ڕQ�e�҆���Q�f�4��X%J% "�  ��U3jk��сmU5I[Zѥj�6���UVX�UA0�e
Q�m��c[+f�E��֔�Ҁ����R�H)� �*v�Z5+THUbilC��چ	�U#T�n�Y��U���Kmj���lZ�.�
�5��(��EI�  g:�kR�&�[Ue��UAA�dUm�1�4�J1�� 6Y�ڍTM�il+A�*�V�i�4A*U*�*J  -�DR�13Z�V���*�4̛j�6�Ҡ*[%�P�6jJ*����J�,d#YJ�j�CZ�"D$� p�-Z*����ڔ��dVҀ�lִ�Ԙ5& @	F�·�|��4�=������щ�& �10S�R���@d �  i��#M%<����6P   4S�A*U4&mL@a@h� �)	�� 244MM꘏P�4b=4�H$�H2T�a0  �l��q���33WkQ�X��ô�=6ޑ�^_�B����8��QM'� Z ����AU����2EE(�K��#�D���CX"A�(*(�!$����C��HV$�����/��4c_>�y�"��N��s�/���c:����1��]O0,�iq�un����75�[�Z]��Z�-JV�,E����%}���++v�9���e������YVv�wA��k���&�RA�{"����SbE�M�H�GY=V�u�t�����8,s�u��ŋ�l0�*���Gf�٢їx^�a\Jk�[ר޵a��4n�0)�j�F�����F��w�_��I�.���Re1.�pi��4½"�����q��v2����R8/�{�+t	�vw��n�&�
L�)f���vy�˷��B4�7K��i&[&��m<F�t��[���@��ǹ-*M<���[y���qh%�1[b�Y:�Z���NPݢ�ځ���A�&��+�-k[pZf^c�,�i-�W��B��xDhՀ�4{��Y�¹u�,���y=�f̓JR;e��n�%n[.[�F1sA�f�3^ŘfA*�U���ݭ�L��'�32n2��W��!$椊�� S ���ev�4����>�/s/嫹�t)�aw������*�ۚ��k�"�ӬL�Ќh8��n;��P�[4V�ɶ.�ٖ�ĨjXYc���v�����?*�PV�݇V��ώHO����0}B�-��64k-���[Y�a�y�
ɘU݀u9NcZS͊��oF^nӘ��z�Z�1`đF�Shm1)�X́W[�ʶ����kq��G0s���
vn��J�ܢ.n�/]5B�Qh�Qf��IzU#�t^�̌ҹ��uaVYYR��Ǖpf���;���3vX���{r/b���kn�3E�|h���eq<�YF������f�G3�CH0U�qәbmʴ0����n蚗Q	*t��0ѭ��&Jw�g]�41"Mij+�*�Wl���B�ֺOl�)�4Jl�i
�����������6���J�D<�KYkc�[0�w2��h�jI<�6���[�l���c�����Gk~�eL8jG̱���[�*�b"�nc"��Bi��ׯe�L�f<�OS�h��*�*��9�K���I@C�K`xŔ2�a���X��m��jZniȋ:��Ȕ74���w�ۙs�t�˺�V��A�k�Ee�Vda�ƥ��I{{@@w(}/q:²�]=��빉�l<�v#0��X�(�":6��٘k.�[�/wr��D��O3KVby[M[@���F��M�˩�t1��+ְ�������c[υ�R�̹wi�n�l�`�iU�YC;�.'t�;i�R�ctVV��aL�e���u��ѽ״��x��h�i�>�"���sp�mM�z���H��<׆�	�`8r�:���nD���DY*�V7�hj���s^P�騀����,�Vʓvm˻(���A<��P�ժ��w,� ())h��!%�#�u2���"�܌`�+��t�=�V)婃'ch�Z�4��5��U�� �v�s^muc�4r�Z�͛	Y�y���̓G���m�0��a�*�A
DVӻ�FM�!�����o)V�f���L���Z.�	v��� A����{j]�H=+���Lz�f�Z�Bm�+�ɘ�%I�+J��5]��հ^Y������ʴ��R�����f6�F����Д�U/f�B�'����kwV�yV�Xp7���Ga#�#9�S\t*[�s�*��n3������mV�]��[�rd.Ԓ(��1�G�kq���4VݔKHO�:�Q��el*RRt��dM�7sb��&�Q{N�h�ɷ�hِё8�u/o�V��b�w�V۔����3 E�mLF����%��jP^ު��lS���qo٪���8�����T[z�*�dx�;Y�o�7`��e�ӏ)�p�H��e�]��
zu�ʹ[�\`���[CC.�"�f�͝��ҕ���١1XLʲ�`5u���F��wY0fLۼ76�k:ƩX.]�jI
�%��PPֆn`E�����/#Kte����ál8�n�gˤS;J��IdR��/��E,�4��
�I'�>=�;�!��`T�8�,�U��ᴁ��+��`<�
=ɞ�W=��Hu��R����ifŭ���q��jei��x����[�U� �Z�1�^��,v�ٱ�ZR������TMK�«�Zcv��;!֢2ɻ�����Fxѫf]="�ǻ�[���X�.�1�lP�[.�Õ.V�Ǣ���L�7��� ͭ��YI5�DNeq���ov�E�ˈ��7�y{Z��[R��G��z�It�ѵj�{E�J$�V�!���r��.�|�Q�kpe��J�
l҂$U�84��'t�!�ĭ��u�BŐkw鼩v��(�ج
9H�l�	U飢ֱ�`*��4����Ck~�*��ɍ裡�Gh`�`�-e��D�j�PE�,^�� ��6ҷ�ه7�V�Nԗ�&��
Wf�:�5��St,1`�0�!Sm���ʌi����6��:8E֌;�Ժ�暜��� r�m.�������r��qK��Sr	J��^��[9F���f�dR��7�:��T���	�tňh*��Z�7�^�\^�|��YE�W������i^��z�]4�O�
o% 2͹��[;�[ѫn�z��N��Q�kej�ҰM"�(�)�å���f��X�f5%��n�ת�^�AE;��:f�G2Gm����6��Lh��s�W�#�%���I<�@ZB�AdyKnC�9[mmj�Q��Z��옛�Ca��Njgktf��80�N�c�[��ͅ
��c�\+�؄waS���kr��1V��I1S15�Xp5,�4�nл8R�0}��̭5����tLǘ�X��%u/(<�wV��{�wV ���j�)��5KmR�Ć���y��t��.�ج�D����Vm,T���+��Sʻ�/-�4]�2��6إ@�l=��K���V�����˗�ZH���E"�݊8��Vu�n��j�(��	(�����/���#j�k^d�1Ov�/wLdY�R*�"(m��	�*n�H���=���/ieIQ,֍^n�U�V1(���c�LƷ�N�T��Lk-D�EE,Q���r����Ɇ�HEQP��-Ê�
btʙLڂ"p�w�T����m&v��6�I%<�%�W��L;$PZ��ڎ��9j86�%���싡 �O-dh�ݬT.V͖S�H'ګ[N��Y��_6�4z�6n���[e}�wY����*���Pm��Lj̤���կ[�Xgu�gr�g��Z�������C(+A��2]3[urUt,�f�֖��\xj��JXޛ���H\Ea;Bn��{Fe@jL��0-hբ�t��'�VY��d�"fu�J�cݱr�mc����{X���O+	���pJ��Y�͚�hK�/����K㶷lĨՅ���kfŊ��T���w���VFjq'W��|8+�|�>{`�ò)nX3�g$Da[Dd��P�ݹ���h�M�T�V���ݦeo�]m��&���L
�
@��ZB��-ߣ�77I�ͷ%@�G�.U�{Vu���p1����͇s)L��M��2KҼX �+ձi� ��¶�B��#/|]�����"�;��*dE"����"�U����"�knI�(�0[Lf�J,��̙m�̢�DU�ʺ�:� /��& �Z'().�3tb˶��i��S����Ռyv����mj�%����g`�eV�V�릩�oW՘�-��7��F��05��e+��j�]�N�0��Mh�Z�vm6�qGN�l�����o�#Y�S:��<jָ�r�x1�.�5�cQ��9�fܧ���hˇ���^�[D�����\��8��ѷZ2k`�6�T�52�R�w�!zJA�lL��m��ؤ֥MU��Hi��C�+KA�.���E\���e���`�q*�c+!�(]۲[�xuX�l��.�k	Ӹ�!WEʕ �Q�����`��*�-���q�U!a�siҳ�������������L�M6��L�A�����W�4�L�r^
��hEv,�5AZn�w-ּݒ��W��嬕1,
�wX0�΀�V��״禎��]9.a{�:�n)Q�6��,�u7H��dv�GU�K�J�Lǖ*�A����(��n�c��le�sSw�֓�*��6�6T�f��J�����j�l���:�
�ۢ�q%X7�����u^Z���凲�����*�KѲ�*����['6�p"&h�e��+96�thn�6CYa���f[�2̫ƍ �2��ʺ�野��&��R;�L�9M0>n�*0Nl�zP��i$���L�7z���-U�ّLׄ�z�{W`�l��ɐ��7j�e�D��4�݊�ѡ<%�B�: mjߛwV�;�(1J
h4g�b��%�m��6�V2�Xv���4[�1+��Itl�ZV��X�O-��Hl�Qok��5�+mY���l�M�V��ų�9��BPÖ��B�9��ڳ��i\�U�ȥ��y�jB�Yٕ2����ǻX�����q=`�-`_���R�Ų�j�z-ˢ�[0=��B�GL��+�NbL,;Y�o×F���;���*%a17N��)cV��eC �Mh��3I�օ�l�ā�G.^�ƫ/*ཇIEKA�F��(6V���{�˰e`l��6 X�t�_uq4o;��G5i���o:5e�njCH��F咫#��[hh�A
��қ����#,�v�b�&衃H����8��+*�r��D3. CY���c�� �.��U�XE`����ƪ¹4P�#-�kj�̿�F)� �֣2+�Qf��k �x0�8=}�y��0^:V˗2��P<�fQx�^�U���;D4/��'z����bzt(j`nދܸ��F%ZM:���A���[o �n��a��f��9��ǣ�V��͂��ݾ�>%fU�&"U�5�Y8��"	U��%�f�+Fe����1�wm�W��������4U;���aZ��%��`&���9�����&�4ܗ���9f�*�ɤi���J�e�݄ܛP_vZ��/>D����e-�=�.�{{p1��`�Q[��nJ���]�;�f��Mw{�<��[@]J��گ3`H���v%��.�6!�`[�&]�)�b�z��w�FLM㵎*6�t��jV��[x����zN��ߣ-�256�R�i�����bdT��wq�����A}7"��2j�����veuu+!���}���e��e�@Ϋ�Y���ʜ����/A1�*��Nq3vW_T�8�Y�匾E#��5�����#[yI��́�s�n���!�-��<z��*	��\݄��2�G���V�>�u��z�	I��(�������C�7�=*_p��̭�7�Q��Gk���r��x蝛J@��VKYéG\�&�]s�ڨ�c健O2�)����+ض�LU�c�I��Y{RFhwE{ë�أ�pj���
:uu����h�Λ7�-Қ�x؈X��鳭�H��.$I��׊�g0�\R�Ok�lDAK',�	WֺR@�sڸV�cKtZ�Ų��(l}:���!�è�J˿�L��s3^���+c����V�!U�tu���(�;y��/���$Tw��Z��s��	"�>�7F�Ѯ��W�ue�Hӑҝ.n��[��8�	ڈ�]֥�t��XT*%2�.m��h�.�.���]\�_���ґj͛j�o2�lp�n'�S��63{{jݽ�/[a-՛���-�Q9��=�g,"2O��;l����A�Ǹ��E�앙@�(�������r��_8_gZ��v�!.l�B]v�>vV��kZ޲�])M��Y<&�򹳗�٧>廫�c�]��ʞ���+��DV���	Zu�۩��=Ϩ��i�ƗbQ�ێ [�U�tc��vѼ���@�{�'������>�'���L[�7���:����R�/(N 1�tB��v�|xE���ȴ��1N�Y��Q� WW�qǻ1�a �f�`����m1��ᬼ7�bT�X)��G;�Mʏ�y����Gz+f����:R��y���6gS�Ȧ%��"��c*;����/w���]��K�9�]�t�,黛�-��Q�˦���� ��;v�,�I��T򴳮��'%Y��
(���Z��.'Q ;]�[��,[����/��u"-u %s<��=6���!�GTWٕ�wL��6��x��нJw��a2� �	�%-���3:��).�<I�%�vR��]�׳j���P�շX��@洶��(s6�>}�X/�e�/~��KS�A���e5����)h���z�s6���`Lke2cåU�ݠ�M�)Ҳ4ˏ$�(�v9)P�h��lu��7;���&Q�8�G��'2�>�2B�sp^4�\�k6h哝�A�B�g;��;0�Ɲ��9������2���)9��6��f�����M|�Z1nq��1@��\�-.:�V���Ec�T�iKl4�j�NWg�C�{�p��b���E��N�+읚��Ş��\"`
ad?Y����h��{(Tl�t�[��Rj=����R]0�	��QK����H�)�ú�u��T4�N�O�h��wQ�a׻�_V�'��̐<�ԧYI��t�'�kI�<��!���n^@M_Q@4(�Wui-v�p��i��*Q�%��	��o%�]�g-�*C/me�{9:��Gem]܏[nŬjD�"n�;�M��G8fT��܂�7[)>��i�v`2����+hw	öh�^j�$j��6�eO���4��;�w�7�U+e�-L�E���
d_V*��n7t�y�I�u-��e'�a��2Zk�%���'����k(_<�!J���
��=�=���t04p���=� ���鑌�m�oo��iR���&�D�e@�ӹ����.Qd���z��U�}؈���P��ms�ǵ�ݑo�7ݎ6�z��(n,t�8.HR+&L��j(��j�h'ck�ˈ��?0�5wY�Zl�x9t��F���,l�(EEsm>o$�u,�${,f�ܡB���L{���cb�wi�Ц��W��H1���)l�n��WC�=Y\�����}7j^����n���Û�`T���Щ�3�MlYݑ���t�`�yS2���}}�q�;����2��a�R��KO��Sv����"�:�
�;zPʱ���y%ʐGr"/Z�3���!��"���8Kvj�a˛�x�w�3�U�z����GK�S{%������t;������'����T5�m�O��r��˼���IK/�5 9����5��T��R��1^9|6�|(�n�#���WA����:yA�]�6�[wD��
��.#t���Ǜ�s�9+.��G99�s������̥#�^�uРn���#ި��8t�eP�	�wz�t���CU��ܡ������~4�J��5w]�nC����/��eun�B�w:=���<^��AH -0�-nq�N��J�w�K�Tͬ�Lv;�r�*�L9V�����!.Sʾ5r*�ʼ7��+B�%��>Au0`Ɉ�ʙ��۔��\6IL�Zr;#��`X���.�eL������Qxo���.�7��th��ݳ/.M�|3c���w.XyXd}���}��#뫖"QWQFC�$��fo+y��$u��Y�X�P�Y+�=J��H���$�i\<�ʖ��ԯ���xIȊ̤�͕��s�²��<�`$�ud�Tp�u�+x�b�h��n���ܝ�b٭�n�6�)J�8b#�u�
����c�k�ܪ��xt.fʼ��I;�%p�F����]v����r��;d���i�λ�='q�FF`#6���wT
���^��*�͂�� 7wu�b{de���I��3n�]$�A�{l)JSX!3kn�r���x
4.M�&>+�
�9
�d%���e8�H;
��(r��x^�7m_�R�E���쎴u�x
ªѱZ���v���@Z gj�iV��5����s)���~[]M�C�V�,�[#T��� ;�\��%����$�@(��Y�*1Sm���Y:ę�9-�l�u(�Rǘp����bR�c/�m7+G�E���G(p�8�	�Ѓ3�WB�RE��:��_e���V>=��Y�&��
;q�ة��c�}�X��R������"sP�X(-R�<{����fZ�Q�0C���Y�[6�/]��d��4�Zv�ݛ��˔�9ك��T��1ϗd�0��.e�)dG썜�3h��ֆl�=X��8��.���Sd���W)��l��J�u�:\��x�\�ا1N���k�E�.�ZI�gR�6C��;r�v�Ϋ,q�֣�-���W[�j�^e��R�5j�쥬st�-�j�E�p՗�.����N���H�L�,
<Q�tnK�(�@^j���*�[&��d *�Z΅pn����BY���-t2@�Y��ބ�[
;��+����7y�'V��q��?2��^��N%{��])�Y�ܺ�xM9�1ȻHy)�r�8��z2q���A{�+�&�[��`r[�e�J/%,�I��Q���\�*�q�x��pŮ�[�P�U
N���A�6J���Eaw�}�^��2T2f������J$�q\�-K��O��T�no���`���~��^�n"����V���v�V�0�����VM����C�Kz� /s�8���	��2�p����>��K.�����H�%��!��ǂ�v��q�z�mu�R�a��p��AO��4z�t49���䜈Zl	9�	�|�6˵���1�sv�0�y�5Q�C)�n`�����o����ia�Q�=��L�B$��yX ��@ⵛ�k�d.��{Z�Z������&�^<qp4 L�Y�G�M����m��V��a�%o�r�V��֑й�*'Y����ا$9�vwu��o����(k[P�����Ee�f�S�H��HJYVt�̵@�J�ucƸM�{�"���r��B�S-��%A�VP�X؛98y��v�e� SAV\$Z��d��{Ë5&;�mRcK��/�G���Ci\�lWv���yd��KC;����� �θ�{z�V��.�e;-�b��>z�B�>ǚ)������çv�1)R	S�:{u{r��R�1�ݘlnL;����]!��{�	q�L���yR��>��1ӫl��.<�2���v�송شk���j���{�p-�ȅncr�V\< �u�ޠ#4xԭ���\�u��;����%^Z�'-��P�j�=-�"�f®�z��+��
AC���ьp��{`���f�e�x�$gg<&�+'�v�6f�8�W�2R�l�܁0�9G��:+4�S�LrP�C��tڐ^;<��n�?�=)�l=f�*�te�z$�7�{�;b��;���m��V�X8�(J�$��gB!�2��N�{F�EkL��Am�	�km"e��\[�a�H��sA�ټ]M�Qɚb���C���5՛E��t��Y±qƲLz&ϊ���K4|x�ೖ��rg�,*5{NhH���Y��Q`��v.�
\�[T*i�sp�!}�aJ��]CI�l�v�[���|�N��.�^G��d<X�a��=���6�y�Ҍj�H�T�<#�F�\Y���U����[\�(%�\�r�����/�Xt����"ʴ�gDEIq���+�Gs���uN�Rmq�x��>�� ���,���co�I���Y�i�w� �5����=���WxB4��M��*)e6-��1���u,�S�����)�-��C�3V�4&��M��u��8����h�C5��ͬ�3���R-&>(N�J�j�8����P\��+K�<N�k�Jۊ�u�q�tf��s�*iN�,f4�5��L�ຍV��^ܩ�G�̓�ce�-U�$�w++����[�Vk%Cr]��$�8�IL���R��gr��h�Jn;�IR9���1v"S(3�bf�¹��h%�Ŗvmt�\uԚ�{���49&��z��������}��*TǇ3��H �����P�Ԭ�9\L:�Ե"�4D�*iJc��ڋF��^Z{�\��Gr�8���d�Arw7�J�5����B�e]؝(Eo��z�^��s,�3eG}ʓ�����㻲U\�3R{+���
B�s��I$�I$�Ŋ̒L\*�t�s0F��˔qu�J)E}��:o��닫'� �n�m�uu-S��\J͋wV�h�^��t�&tbь���q�#�#q��;n_\72s�B�R�Ra]�x�δlޱ~�+h�޶S(H��#-r��Ӯ�Gml�u(��qD�I�غ��,�k��[�8�"��sf�0e�[L^�K�k��iz��������Q8S,��B!QL�$��PDK�[4@�6�f�1 	!#�`MvRu�K�cY��k�y�t��j��v�mu���z���a�*Ĵ�wVýU/�pR×2<�ю�iwK�NM���Eahy�r�M sCc��;/�On�� }1!��F=���s��F�KZ�d�wH��k�%�T$���jCT vu@!	�f˦����v֕�L���=�*�op�ʴ�m����\o�%�٢ӫ�c76�.�v7i֝�
�"{�'��y��J�ٖ�4�M�Y"��3{�w1�$o��F=��
J�b���Z1^`7M�G5P�*�m�M�ݙ(��n�0ep�T��#����&���Y�箮��Æ�Ԯ�!�^hE��ҙ��>]lqY�\��FԹoBX*;�;��
�6Be���<f�<m�.��GG*vOL�+��P��Q��B�m),�3.Wf��X�ú{JxAki�jo�|w�H�:r�Q��8��lצW+���~.u]�yucp.]�@O�5�ӫY��.�����$�͎[�wh���P�z��a� �)iܩ-K�E���]Wsc��z~�>���.��(H�9�sX[�iH[I�A��۱���;	劤��d�O��o#%�*�C�S0
˒�Q��Wg�N;*s��0]i����5ʚ�>�{H�clod�<�{�흦��{*�]�B͍�{q�Kz�a ��#�yV�XWt��2[+�)6�4�ً9F�e��F*v��ڳQ��q�Ư1�Bt�סgR,�[�5��0���
q�&v���満ŗv�wYՎV���Y�@*:e�-*�w�e'�-��w(6w=�f��NlQ����[�8��{�u�j*����t�?��f�8��s�xk�紗p/ح�1u�X���b��+�ڜ�U�/\U;,q�	���г��łz��m�N��Y����V��Pb@ޠ�dW��8�oV��c4X�[�S�+%-�����[A��oi�]��1$Qg��[��*wm�4��Y�;5.�f�1E��w}���K㢅���X�,T4�e�q��<25���P�a�3�X�.�V�J�1]e��K�N��.��y��$-�m����@
��*e�Cn�O$��G�����1�Y���ݖk��tc�b��x f�U�^��]� ��<J�.��!T��+�n'�6�u�Z�.3	$�K��M�vi�yh�ӝ|}�ث��iq�\.L 1��V��u����N�����;�E���7h]����1 P�F�)���GvB2����y�ځM�;n�d�s��P�7xc�"�����>��A5��+�A		����%r��%���նsv�k�]+�:)Cs͏y�š�yt�-3����EJ�Q��pʺ�خ��Wj̶���"���H98�W�	��M�GiF�����и��#�sx\�e��U�{�n机�����[y�(�; y��@N���tAG�r�դ�m�"ƴ��풓�	k�\�aO� �\��M�cG+s����Z7H�o��B]']p�f�����X�}D����˚��a��9���t�����]�}�E��J���m��g�.�:�+�[o2�Q�:v(j�o+0�ݹ2�]��r�T`cBr�a�+��J����Y�u�^�wR焲7v�f��7Q�g+1��|�p����!AWi<�pp���9H�Yk���$�7���֕�:��]\��t�uZf�� �x�@k�}K��Bl�InG�O(�VY�u�N�+*�q���1Q5/� �P<1X����e�iuv3n��G]��
�Ed�4��:�:�܎�-���,�ؔ�@e��̶;)��e�cf��E\�i��nR75�͏��Ե<hF�.vl��Mw:v'�����C\�*X.��[��3��!=���D=1Be����v�Ȧ�� �wJ�+�|Z�ד)�9��hu�J&�zL�NOb��%�h�zk��`�5ŝ�V�f��s�l�V�"�x�l�&�X���j��ab'/j����{N�.���!i_ ��?�>�r�}q�@ٷ[�&���bE���	�W*kqvZ���Ֆ�@|mKg��t
FOm,qK��wF�
(�Y'_i
�8�()�*�}�+w�(+N�4��s�6��B���Y|xi�Z�3s��PZ�/Ed�۲- �U��h�x�Y��,F��.��r���f���[U��P���K�Ν٫�]��L!k��)�v�/^��,u\2�<�NSuT!�����>���Uý�]\������)j��ή���.�ua��XԐ�|����-p�Z�W[�6�i��j)�8ὁԘr����)��YEp��6�p�Ű^'�
2`��*D��aG��Vɛv�
Y�����{���wnƪ�GV�6oS_+yB�m�9E�o]�Da�u��m�yt���x�uVz�M�' �3�lip��ZS�ck�3pS(e��{�',}w-
e�'�i�U)U��:*�A,���V�l=�ܹ��$�-v�:�Sj�PΛ��FV�]��`U�{�8��h:8(��.M��6��a��q��zBa����5��"0ηu)�i���i<��䲷ta�#6�@�t
32 [�Ķ���.�[b��K~�A)[\9�
��푡�KN<N�fVx����wv�cWro�D���1ؘj����C:gu��"{��uj]�R�L3(5���.���S��PT�!Y��0o�t(v[w�p��2�|�TͲ�72�"�ا������� ��m��2c2v�(X��tu^�L_H�`�Ps���b�8P�u%�[��K��h�ݨ%K�3��F���I���)���[����B����.�+��AT.b�$}&nJ��0��j�tp٣�p�z&1J.���u6��K� ��rѫ�)Mp�b�nl�;�͕VP̝"�s`����z��r��|��|�g��}F�9`��]�u��2�4ls��"�X�[��9�	���C:���D��j�;Au}1��/;��U�;��
���X�mYU�g�(�vtk�5�ަ;����*ƪn���|ن��9�l��*���\�g�]�]�J���m&@����Vp-���ѭR���j�u��Q���UڛE@���.�v�R���:)ס�|.mEsG'��(�G;� �㴜r6��; ���Ի��w@��D���N�{��4�qc���a��Ljs�X��挸1�uY��j���;lpѕ�|2(��#�I����/id��R��u�X�\׏"��b��*�a%Ӷ�fi����Ps�h<� ݣ��eu`��)+��_6)2gU���S��Z��+�6�os-娖����a�
sJ�Ump���k�L|��0�3I7ʶ�=X��Q�n��^t�� �k��"�{�M�ws���s}��m����KMwuE�@�7WY��#�;��wǪ���	�	ۏ*:;��r��瘫���'	���!��F��Z�[�j��
S�
僉R���Ù�!�qH+�5N:@���0�30K�O���c��r�*[�:#ذ��ݭ�Z�W�}�,���o8ѻ���*���3���,���Vυ������ 菕 �=f�h�ιdV`���s>R鯞�*���촱�ܽ=�p�O[�/��<˭rPHYi��|C���N�y���#����gu�=�e�7�\���o�v��K�g�aRD��jh��2Ι�Jn��e�Kz�[ohH��+;VCV��V�,-����}.��˺)��A��le�9��G��ȩ������ߺ]�]�x���J(9�\��!#g �V�Ѷ�M�O`�U)� ����}�����3��.�Hnf�aAE��×Y�-�Q�Iʇt� ųn�p�U��j@1凝rb+N��[C��¸k(�b��i�wv�LV�f�,�I��J��:��D�_����[��ӧ\��E��C���/,����\��KE�����w4�j�&�f�d*�,�WLϜ�.��0�[��dmi�\2�� lr�*q�7�*ܼϔ�[�ih+:�`;�p�����8(*0���;��  �8-�_<�}!�#f��U��M��Q���fEż6�;���a�e��f*\�uAj�a�j�ՠ��ֳHosQ�7ۦ��^��N�n�uϡ��u�Դ�5j���u)��A+�#�ɕ����.l��������·6���Ǚ��%��)��T,-�c����r���%�\4A؝��jZ1ibeES�#��S2^�m�y���N�$e�<�D]Y��Tm��5i3�͏eJu*�d��y���kx���&��	�� �jPJ��%�ճ�;�	�[�|��	p��l�:a���2�;j�w#[��v�i�� �5��x��%1�P�rm�23
	�a\�����2Q��͏2����>��)^ok�2�	��m��9s�Q�X�o_$A�~�t�mc�>�Z�添V�gQȱ0b�{��w5N��J�=jм%z�޶���ù{f��㮄�M���\�r�em�0$V����f7ǥ�l�p�Y#.��$qS���:M8'��G�H�����K7�ϖn�v�gو�C.��e�"�f���V�Z���cxn_&����EA�95�鴻�q�E����OE�u�U�٘(_ݦ�(�S���q�W�^*op�gNÓk#J�f�ڏG�In�X��Y��ӗ��g.�����Zk(����M�:]���t
b��%o��v����d�T�����L{v��#v%ʄa���5u���{�fQ�s��"�R��z��H`�mW9��9�Q��ӃWv�s�6��u(�+�F9\���8�������j��]%+����Q���j�$����%�.�Q$k}F�c��[�u�����J�f�[f�+��V]`�/�8E�be��T�E��Me�#N<������ѕ[đ=�`clNN���*0��°�6�r�!�c7R�=J�Ɩ�k۹�C��b6��Tkd� Ll�Ë�.��ic}���S,������B������/]�����vԝ�MGw7��`�81p
�u������嫄TGY�g^�t��3#��m��1����7�����&���.��[z��v��[���k2�R���� &��W9J'��`�7G9�H�-�D9�Z�ѻ��ov��~@�*Ezd�;�2=��� @������kF��o^��C,.P�]�FK�[Y'yK6�bQ�P-:�åܶz�ƞ�
�`lђk��8Q�#Y�.ﮉr���J�o5R�)��S�Ή��i����[�t��r3��&P�g�'�;��js2��t#hS����nY}�\��0��U�k���ow'^<5���$��^Jy��G�Y�娉=4��L]+K#]e�
݊5��F��]B�U�o��u�Ef�u'�(Gco�R�av�{}�7(>�����zT���n���9��'�'<5���k���YF	���Lx�SQ���L�iͽ�Y�ß,���2�9oob/l<�}v�� ʺ�wSp����t5�_�֜vD(�V��Q\��������s��ۛ�:ӥz��m$'P��.K��$�E]ׇ�`�mӡ�z�^�l�4I�{��
WuA�';kT�����	s���\��+V����eID�[5�$\9G7;�t�$&ɗy���i�fA}��FMk��{�v�u��y�N��<��TUH�M�"�����UXT��PN���J#�Q��"c^��(�dE"�J��;�QAE4�D�Q`�U%j���b*���(",�+,\jf%FՀ�A�Z��A�X�$kKeKm�Q��ьgM�]!SV���.`bL˃�B��TE"1ml����(�ѝ`U�J"�+tѶ���R�
؂�PEPƙIFDEPTE-�(��l�TTƕ���(��ʆ[���(,E
�U+UE�����<��@s��6MF�;X{������5���.<��:�~�/;��gM^l��:�N�����4�w�����hw����:#��#*u8�#����o�&x?#~_��OuW��\d���=�sk��o���OV��Ї��&1w=yǅ�R)Ae�����L��}=j���y@�4��]�G:���(����p�u�.�s*���
�����a)B��5���^���$�AIP���/N=�9��� ���E�.��j��K��0ڻm�Q�_��U$�jnzXɎ1!i���]f�����*���;�iE9z%�+iz��Qͬ^�h?g��(r�nQ%>�F�LiE~��D��"���d5-ʸ��N�������d8����| ޣ�E������6V��&$����
ډP��Wf��79ΫDv��v!\�>=�s�FP2�)re+*��Ɨ+MՉXF�P�eZ��vɌ\�0T�Hތ,���kj)~�U<�_q�P��2��=Lk��{�nj]�U�ۅK��1�qU=#�V��rz��"b��F��:a���&��1nc$х>�,u�"���h��l�I�m�	��]���1��JYD��0��ta��{���I� ��ߧ$^>����Li��J0ҵaI{e�5p��iP��w�MNUf*��ol�1��ά��R��t���^o�k�KB�y�@�m��L� �{Ġ{v�M�eqV�{�~I��9@�2�;�X�#]s��T.x�f�^�aV��Iנ����y3O��y�pk	�o'h���&Oy�~��J����~�ٸ��r��(j�gmn���b$/��;�N��ô����Xppn��pfv��oB�Nf��z�4�.J��5���ݥ!�PwA�Z�t�ufS�4���&.I� _����"Lq�O��[ڎ{�[�P�f��U��w�f:�5f7�G>h��1Y�5ps��n]V5�-��xڸ�1j�$%hU�'���Q����1���9�w���z��/4<�U�*�P�㡎���X3&�/��������+�F�x�Ve�J�A���{�]qz����}����QU�"'-*��.��q��u�����ck0�F`u�S�z+t8�X�_E��_f�+>��*�;���<�'�M �7`��9{xL���{"�*���� �F�ӊ��U�E��n�:YgR`亮�B�	I*RC�������]��z��z���2+} �܇���]�t2�s隍|;oe@P�bw<C�w�x��F��Fq��NS��c�(=8�ׅb���y�N����:G������4��U����2�9��+�nV�z�7f�*�doQ�9�1�6gU�X���"��ᜤ�l���<��*������gO-�>CA�
5�q�=�6¬�X,��R�d���I��Y�GTN�-�K[�Ɲh�ڲ>Eڝ��բg����Sx�f�QF{��=0���`�<��j,5g��N�o���\�ؖ��I7�`�82GD�j��_<1|���,9}���/yo<Tz�H�2#P��noq�F^X%�ktw�ִ�jً�*/����)ڛ�S� ˁ�d�^��
������Qq�a)�7�v��J�����^��T�I�=�Y��`���\V���{n΅����(�)s�������>�SUp��3���=���Q��ɽ�~�]�7�OX�$�:̸�3���d���Ҹn#�Ij�CZtX���}����
ݶ�L_I#R^�c���WFC(��m,��,n�`u�8�L�����;Y���ey;[V�EKMѧ%^,���<��|PU :Y�P�*c�R2�ol�뺱�ܦngi��8�uV�{��Eю�x$��c:�j�\�#}��y7)����ӑs>�n��[T�=}#0�CZ�}<4+����Ӏ���X�sxc5%�-�����F�P�7�C����^>��CQ�ܬ���˻�7���s{c{�z��&�]E�)sb��"x�Z���v�aU�_�ŵ��/k��Y8=�36%�nx����:�W�z��^��JI��ڋ=�qB�W��%[��.�����v��|K�4-ֶ�i��g�NC���x�cM*��VA�[���}����\�T�}K�GMZ�Ǜ�T�����f�.�;�T�hM�rC���E\a궪޴��kmUN*�۽��6u&�g1�ALq��z���̍u�e�	�P2�S����������E\R�GC��Y~M+�90f%<|�w�鐌��Qʎ^���5�|��Oi'5�����ڌ%t��5S��'��C(A���y�}���yOU����*���L�P������ܑNٮ4e���-����yʱ6�$х�X�F��ldoe2��Q0
s�Q8�S�Ef+�Q�%&�W�	u,�E� �F#��"�v^U�Ƨ�a��9�uG�!wvC�:TךA���xi���űؒ�驺3G�
uȃS��1W1+F��-v�,U�}+=��q�9�;���Z����9$Sx]�<�JlT:fo��rF53)����T�ZЯK��o�x�龼��-�EE��vg��:1/���������С^�Qɀ<�^0��-���wv��<cz-\Vd%/{.fo�b�,d��L��H���ٻ����m&gy�S���{�u<I��e�����b��"��e޶t���;�b��R�l��[c\�i
�q��o��a�{�7l����,qq����V��W�1���4]���,�F�X�����j�T#�xGO�q��-��]}6�񒂓�z�=���d}��V��K>���i�X��r�u�����y�/9��5^�U�+}P��@+��(�����Hmu���!��i�%W4����L��]yn��m9V�gA��o8�,e��v��0���gT�̝u�2�ح��Z�QH-����A��Ӥ��N}�1���\;:�.Xh��m�r��4�:���;�]����B�UY�t�6T;��cj�o;"�u���V�}	�2εv�7�Bܲ���иC���L��Mzb,��,�2��䶡A~s=�.P.�iN35.�#���I�U�E�ST�9I*k�!�Fu�f���5D��+'v�Y7�U8H7ϖE��t��X��o2�{J����\U�
����_B���$Z�)��:���y��65����N������ g{|b�����[��Sf����!kؚ�	�*�^�V_.<N=����]h�3i��=EV�G� �}�sN6��vg�ms޸µ��$��S	���I����vǃ�L+$]�з]�}{�g��p�C6*6T[�]�R�ٷ^F��oh_C�ޝ*�G	�h��;�/���- �,ɮ��� ��|�|5���yN�A5�l����#n��0v�w�g9z���&�W58����U
�4�6ѝӽ��oAor�dH�n�g�0�yY�j����2DO��6���P#{�e�ۀ�n$�o`�
S� ::�J�\[�:�E�"�45s��*#
�+619�뽝��:"X׊>����6�?L|~�����M�1����iC;Q-$Q*8�Hu�1^}�z�i�J�M7�s�W��⦭ٻݵCIׂ2�R����P���b�0�ל�z�j{��������Ҧդ�r8q�Z�o��f���G.h��7�/�H���R�tf�KI
��+��f�Ѽ��ʞ����tu��1���k��B���0f���y_��-d�V�[�h׮�|�z�U����<�9�L3��85G�0�8�e*G$j:i������lQ
��V�f�.��pvr5չ`_-���qȤ�zyJ�.z�G���I���#[�Yǒ�Vo4�;����3�e&:�o]���5:�[�VUqJ��i���n��F��gZ.�s��{�ء{91��ԍ.��M"�9T'��؞vC�I7�R��t��z)3SY�7Y=1���qE5��گ��3�:ܞ�/W56�g�Q��& =Py�Dk��7M�v�5����!�3�;�r/ː�&�A�V�s�{r\�Z�Z���l�H��4�.%=%�>��=CJr�������7ڹ8R�7���σ	:�]��1�μ���W�������k��=��qC�q��7*��Ǯg�����}�b{��f�I��7�7T���F�(LՄRV�[��m���q���5�Ɏ�sm�;(��:��D�(��U�A9(��잝�aڛs��7!�r�H�R�RpX���X�l���/^�W:Yp�
b��k��an �Cf6l����n�gErD_e�W�uN�J��rG؝��͒���ӻ�Gv��Z��l�e������b�m�eՖe���[W�M:��(�:p�%cT)Uv
���#g]�m�i�_�e!���Z���f\tr���p�_A�M���֮��	�9k���J���m��6��a�ټ)#s	�ۦ�"��X�f��X�Wef�a�Vf�˥ՙF�����oP�aM�r���X^:��6jC³�IѮ��g�[�'�ګ8��w�J�y$Ǎ�}`�MG(���B��r�ݼu*���D���佭��zF
[�[D�Y�`p�3n��z�wX\ӗ'BU�J��:L�뮳gE�sh�o���ZU���zh�����&���m6����)�	�l��h�tΧL!�#d뱛ADwŲ�OX�e��e����@��3�LӶ{Tu�r�/��#���>F��	�H�P���W�35n�M�闧{�kp�u}��v2D���PKokM]B2!:ţ��{�$t۝y`��%��H�W9f��i��6l1�8����H#���ɑ-˄�<���3��V��Gg%9dƅ�s&�e|�vTY��>��)A)e�f���+��7h;�� Qic8��Ba�`j�H�M�B:�f�n�D��c6��];zl�ں���x��f}a�E���B[su�"ִX8���9�m֧Ь�����T�9F��7$�x�1Cgfm:�x���K�	3/�
���`c[��,Ɲ]�m8i���2dR��)Qs9��y�v5��	^�?z#e�r0Q㔑�)�><�������/������)�P�:�Np�k2��}n�i�9Zб�M�Ar،[���6�F��5p��oʰ�j���
���q�k�I��L�b�o�]�'0�";lٗ�d�nB'� �����osn��dw	%��ڷ��`Tpޞ�X�!wѡ^�^f{�|>?��z�ժ�b%k"+Gl���U�(���dUX�e�����cE#�b��*EX��&*�� �kJ�2(*1E�
����+P���*Vш�*�aJ(����C��X*%lA�([�j�1�R����(�0��j2�D��YR��e�V"`�e�̌m-�Ȋ��e\���q�mU��-*�����h
�2�X��r�J�ӌE����T5lY#���EH��FDT˙�!R)m���F5(�5���*c���
�Tĕ�+�b��i[kkY��8�U-��Q&fb���1\b�U��Km�7���f���~��.mv.�T�Vs��n֊m�E�v�ǒv��qy��k��v�ԙ��R��r&b�]^d� '֧$׌.�p睞;X���\mR=��� +Y9�S����3呶���d�|$_����ݎt��<3�����{��ʫ�Q�[roL��ξ�f\:���)!�`�^��ztgvg�5,���ڒ�i�wGȥg[����p��b�d��Nj<��ˮ����S�!){�i37�)+�9V�,��ݝ��ރA��K���Ԟ`����fYl�$��yݎ���TLV�z�Sl�}�rʢ`�r��)��E�oY�(�QMK��*出�Ҡ��d%-wP�]ݼ��T��c��������G��AP�_5������5�O2v*���T�*m��u���%n�������Qw�����Y�A�S+VI��w����Lrg%��u��R�ޒ����dr��r̰����WY*t�6��jK�?*�z��0lˍڢ��17_g�f���+1�)�s�h��.7��Ưw��F	�򥾵7�{�r�T1�+��N^�o3�f	1I���)�Zd�5=��\�����@�L"bq��T�sr�ux�km����s� �fZ�6N��p�n�.W\Rqz~��3G�WGr�a���@��s�?��OvƘ{>M��T�Ԍ��U���ht��Ys	���ԕ�w۱{�L����pd��ץr��������Q��k�dv=�T�V6�zt�A�%�F!jS��r������U厱�M�E):t�3�p񧻵b�V����6߽��{6����1�na���J�2���zx3kwl����<y����
�vW��~U�c;Kz�=t��cW!z���+D�Yf��N�ps�,��.���ܛr^)�������yF>���y̃ٗŇ����.U]�x�A���kG[޻��Ӟ��|v�M�j��Ǻ��.�m.q���ο2̵�H�2pv7�F�g�t7ۥq%B'.����F�;%$�)�@�ʎ�"�=�)\8�~�^dj5��^/z��Sh�H�]��ɹ�EϷ���y\jgyuk�O�-S7rȁ��Sz�����פR'ںO^����K��	����b�ޓ�'��(��z�E՞�sU�+�V��\}oo!YNM��8��S�^�J��X6����M�Q�]	�8=�ik�
�S���9Tqc�Ì>�����y�s����2��)pW�d��:���������x���2BH�c�(���ok�f�,�����m[U��gȎ1Y:1w,���uk&�r��3#Gmq������6����8��.S��sĿ9�1b�0���9�v��#��-���'������asܮ����M�'F3�� >ގ��z͝%��9�F+���g+@ǳ~��tG8Fl�+7�*C�}O������7���ӕ=�U���ó�2��$�ou	��_B=̇��Q;=~z�b��yų���!��tO�=�Wo�z��-ڽRL5���J0��o2��۾ڹ�I�iY~k:�g�s�]C��*���>y;lz�6j�է�3�z��Q��d<��uuU�����H�3(8�ꁳ��#z(���E�E�%Ϻ�m���e%Վ�ݢA����L@z�y��}Y�wx
ǔ�T^I�.^�f��ʰ	I��/���|l�Z��1���M	���8�.��]�{��'���!ݚmQ�Zb��p�tj�M��o�r�mG���@2�6��7#s3���ã0�?�̼�Ȯ&�EO;#�n��5,'�r����:2%
p�,��5���E����<�L�ӊ��oq���.��U:jL�w��P���gT�P�g�V�nW`E�awX��x�T�
�9j���.�P�+�rm�/�(慽:��΄�(��*u�/(ґd�{�����W���Ef;��Ò�fh�|���[�u���y�1�$�9�8���؝�+ =��@�����	O5�j�4��^�&��t^��ۛ�ˁt)G6s���k�K�w���-�Qúڮ��"f���_!��y9���d�ԋ����]އ�jq��,CƢg�M�w��35X=zp���i+`�_�N���4�7�yۄ�����n�zϑ��(|�J��Y}u�*ͬ���ś�N0�G�B�#��1I�[1I�����9@��փ�)e;|�ک=�2`���J��½ϐ]^�v�}2��+�ٽ/�B��K`��닍���^�*H�4�r\���+�ݗX�ݭ�b3X�m3k���\�w�*X��׆��H�����b�y8Vr���/���U��~��q3Hu�>0�
Sݾ��G�|X���U3��V���\�7�(Ӑg۹=Xq+�+*9�g'V|$�HI�!��z_	�Ү���&�5LeF�WE*�R�9ڝcf�f1�>l=�\��\GXF�m���f�+�7=mus�am�;���)49
]v�~eYw3���6���>ʴ�L��w�c~�a+�����<T�(.�Ι�X�Z��7�)��Wn�����.���ܐ܌ƓW�1��TN��q�.�Q��f�nѓn�+��^���J'c���┗0]�1�*o�Wj����iŜ�w�;]����.�]]<���4�EG)%JHf�����g��i���G���np��qQq�J�~~�U
X���g�#H�{v#�/H0-�&ˬ7�@<����΋��9����ጝē��k(�t�1�+0��f᩹�{.@|��k�Uc����ʹ�z���[EsA{5;�=�y>)��H,�v�^���9e�Ӝ����{�μ�\쫇{���7��{ǶRM��3�+p����=���������T�~+~�{j����gX}��۩��H��W �N���P�_y+���:K�f��*�ByVS�,ֈ͂j�3�o6�Ρ9r�X���/,�T�\�s;T#zՏh.�WVNl�x;�#M����9pKWA�hr�l�kE�=.�پ�or<�x�]� ]$N9�&��Vk�֯yWVbt���M����o�G_��.<:�1�P�(��Q<�FaX�g%��*��x��]C�.A���3�6��i�7[����Zp&�;�j7�#bg`�(w1^}��S�usp��,��)�n�V��؋�l��,v �wR� ��h����E@)��zq��S�V��e'F2:�Z$��niW�9E�r�b�m[a:��w����^��/u�B<e�N�=��ρYC����Q��"WlPwuى�)�:�T-}7�òb�2�M��޵']�N�sz��̺���s|^㷑�xc�l:�[��Q�=�P�f�W���{{-
�Q뾰n�tj
��y��r�.��e��)X˯@�1��O/�oD{��P���]�ڐI8�SN7�aE�\Y]ܰ5쮬ݹ�k��9H��n$$Wc���d��f�'J��W75̫S��ꍭ�m��/GhQ��=yΡ�E�O9��\�d�Z���Z��T6������p^�l����f�q�1�]���j:�L@z�y���2r�.%�N>�T⋯7�7	O�P�D��'��W�3,���t��Ӊ�P�����%�>��f��m�V_@�N/�y�t��%]�^�5&c��(B�y��w�#V�$mH�]��k�}��TuH����T>���߻�=M�~��T-�)���*�d�Ƭ��*n=�C>)'^=KՁ�Z7�eZݠn�9�&��c����|ڭ���7��,�Ҳ��K6�f�J}�pv:Uw�,�ٵV�#/���Y�0yC�Ĥ�T�z�c�7��7�4��elxp7��{�6\۬"�D�D_M��'�t�Fr(�_�{ޜՇ�7�ٿc�p���P7�7s���^R��f��޴�+ڢT0�qS�!P��#N�ΐ���Mi0��Ou���}���U�5>Z�R��k�Cu�wI����>}3��7>�':E⺆#��z��D�m� Z;���|��}9��aK���=�����iÁ��s���.�{�ZOJ��ꋔ�"��Q6�.�]��]S��a;N� �z3�K�a�P{$T7YĤ�;{Q�z�~�yM�Y`�86`��Z|t{�f��-	����qbLֵO�P�H��*��^�֟q-�/8����[F{)��9{hCyL�wu����Iz�vfoKg�5������V��v�.�ƃk�8N;ޖoX�9-�_Y*�]lw�ԡ�^��g^Cڂ�	�uo�M6lM2��n'G��{����q�x�ѥAq�킞�٦��ϟ&�ݻݫ�u���!Ks2�� 95l�k�nvm-
�hbw��/&�E_D>�ol��c�i)�J|*�Һ���f\׏R� �ͫ�B�ʚ�䜺#�q:}�Ь�=�>R��#|��5n:�Xި6���V�
�&�uqN��揟V�uR�P��rE] ���0�ם�VQ՝��)��wr������<Xt���vœ^��C.�������jT����6� ��eX�goL5�(R��W{ ]��$ZiNW�rj���Y�6qP�ݷ{E��2�I�]�i�xsis쒋�&=:.�]��z.�J��^�+OH�q4�vl�@U���g�O�I�"ˠ���]�'���Ec��*���s(�n�!���U�E�� wp���=,�B��L��SD�{� Aq�٬�:�ؾ��㋶��Ի��ͫz%c�!��Hʵ�߻"�9z_�ȞLjb��+s�d�ܱ�V����b��[E�v�	>��#�	�$�e�����Wb���4N��� ��<�u�F4Ix��k�ל����ru�2�w��bi&�C/ZV 9/�r��f������#�l*��bPU4�jQ��wG]���M�׈��Pl����'49,�*�4�m�y��h\hT���;v�<F���gu�/(cu����ثX.�=�#4�(X�+f�u�|�[�-"S����eN��q]م<�����d����Y�`Ǣ��W{��n7�׋i
hYVa�b/5�+E`�l��i1}t�}P ����z�\��3r��Q�lL*p���Z��Y��Ƨ�L�"	����X�u���;Bֽ�b{պ(�Vs3*t��@��Ǻ��J��y����Y��C2K�i<�����h\��[�Bs��1��\S(�?En�Zɽ��b:6s ��!]C�LQ����;t��6!=@m�4�OmN�gd�w�J�d&�%G(�������6��gQ�/����옥��%qM	�aeV��S*��eMe�Ll��[P����e�B�Ym�6�����Q��hR�V����W�Eb%3.U����V�f8��֮&[Um��Q��[D5n&����.V�fLְҵ,j\he�,Uq+L�k*jҥՕ%`�\�y���ң��+m[lJ�YiX�kQKi�9�T�Tkb[VѫaQ\n5RQT����J�P��Y��f��Mf`e�CN�r���Qe�b�QbƵB�H�*(�c��[J���CI3�U��(9a�i��-��K1*�l��Q`��ej�5*�++Df�Rc%Uc����E���(�b����2�,���ѫ5�pQT5�`�j��D1�cR���0���w�.c�y�|"��������8�BJ(5�v]�`r��':N�ެ�u��23��G���l�s>Ŀ@��*�bw����ܕoVyk�3(��Z�em~�Ui�[��Z�_�"���u�R�Uܸ�����N�C��*!���@ۨ��Τf�o����մ�k7�r���N�Cl�.��5�B��/I��ȗ�[�{����5Lx#.)V�lmR�T�4[<���"��]]v��:��S��*Ig� �>�i��b���y����q{�o(��{3�9y�^T��HWS��6^�Y�iɓO"~Cs��^΃°.��U8�t>�^7������^���C�.�F��y� wg�?>.�u�������g��O?-��k��	�c����832��ؾ�����y�N���aś�d3xڬ��㘕K�PSJ͎+.�[�	��>g�Aq���::"s�wvWY����9	�3�c��r���YF��z�%*\����Wh��7�\��ɽp��-��O=6��1D���(��9F�.�حE�Ov8�_�ב�&ЎX�*�Ċ���f�	�)��j���[�������25d��sS��8�`�@���&�w���W�UR���=�Y!�9��|+��q5��Z�gD�:Lu��W�wT���Jq|�8����P���j��5�ђ���i���7
Vո���xyT�%C,|bڧ.0q���-��.ˈ�Q�F�4m>�UZu�}k�z��A�����O�Q�1^�k=�k�V�5Hg#���,�V]��5Fj=�1�:�M1L��t��x��5J&��Іn�+K���G��i�Z�Q��-/��-hV�p���0��d�,7H`��� 4f��Q�w�d��!"t��LÍ,��7%Ԉ���pfV(s����B������R�K���@���t#{�/��m6�wp�,��s��fC�yo9��8{Xs��o>}��]��6��Amt��Y1wE�aS�q���
]x=�r�3�p�^e���Q�8�[��;֗���N�����=�z)�l{'��3~~o����j?c��8�g��_� �J�VN|��a��=�qǝ=ɚ�Qh����m�����7��j���x"���8t^���H�ݸ�f�L6��@�[�����d	Kj�M�rE�YN+��e=�脦�
D�'DEL//1�Tl����7��]�g=�Q0V��z��5fU�o�W���`��n]u\hͧ'mb�"�����M^�;F�ե�2��e�7:��@kI�*g	��WIj��;�f��,,����D*4��)=b�����(�us��6��-�\�~U}�c��\��?�5���s�k�!����u$'������y� ]{�� SU���t>�*�L�9��n�C��r�W����֑��3�O>��m����7���~[Y�=EY�g���u��<�uq������	6g��Bg�j'� �ܠulf��AD�y��qj.���-R���1�JHkX3a�REe:����0p2��J�4��*�a�7�_Mho3[�x�������,�������bAD��4.�d��^=��w�J���}7�ٝE,Գ��#���洔�������k�oZ�`�0�����gz���HmM5z��rp�7j����T�l�1P&:��|͵���)�.� �nŢV<aŦvT]D��4�`���̫˳�̘�Nʾ��QlXP�]m�םȢJ����{)m�}���N���v�SWH$�@�R�3A�Ӱ��$P]u�3UE��s޿an��6�1�	�xyp�9��@�ỗ���ެ�/[���}j�$vKY����x��E�oJW�jgx_3+EAޘ���j�m��(Vy����*N^�N��esd�;0{�ڡ���Z��E�"�L�u�j"��)��a�/n��l�uQI��C�km:ȥ���;�%�-�3j��L7��� ���px<�/"�[��/����f��I�������`�Fᘞ��v��9@'r@�j�7��t�\�0r����-�^�X����*�vU�Tl�v{2����N�6k�90�ƨPVa���{� ��^M�B��˨}7x�(�i~�X3l�
��v���:�����f���-��fͦ�jNr�9�U ���)侏{����؇F�L��v�~_�O�?K�u�v�\a+���|y-�.�ZzZ��x^�騙4��#Q�}�LR�۬��/����^ت����4f��U}��O\��C1���m�����o��qv�3���u��(��O�/@�<�rY��G+G��2�ʏ�G���i�`�1�3��hb��;_����E[5�G��O�2������M��A��v�=ML�[�Ό��05��-�F�Qʠ��[���(=̬���V�w���HMX<�S;�
P�!��8�J��H}�|�_1���7�l;�#{7����K_0�qo��
8���V�t�?Y������~�S�����<�5�+_r�8��dJ�7�.�1�2��a1������ol+ޗZ��q(����s*:S{Sڲ�M��)�����ͨf����-���qe�U�u�އ1����_}UX�i��f��ou�͂�:UU(��r-u�y��=-�\��#k0*�3>4�Rc�e�]��X���>2xJ���B�����ʧ [����k�ur�d�7Ŗ����v��=cmM���{#*�Dr�v�[^�%�כ�ڎ�R7��x���b���^c�6v���b�S��"~�{���+(vy��� zHv���w�ս2���FH_<���Z�l�~�yx�V�s=i�*����K�O��~3ώ�=k�N-ܫ$���Us�Ogj'U^��l�Ҳ��r-���hEFTpf���/Y�nKtp��sz�0�ꑑ݂4<��^^�rm0:٣�$�����m��o��`�=:9�|,߅r7X;˷�H���/'Wq��A͹�-�����X��pd��_=M���ʾk�qw�~�V�j�+�������޽����n�,�ɶ��RL�#�t,������T�����3v$���WaGS�m���7�����#��,�)��_7
N_=u���Oz{�M�����B)�غ&q<-a.Js-�{~�����*$���E�3�d7�R��b����{���i�NK0i��T8s3-$X�P��"�FJ�g���Z��D�B]��9}�-�ke���]^����l�P�϶{+����{dӐ�Ź����1P,�˼�����ݒmN[��8MP�k�aTė
��j'��"O!��PF�q�o(ʾ�X|�ʨ�u�tźQ\�#��I
�X3W���'�<u+˚:n�gl��<4��$3� �8J�{#�����k�j�k��Ja�l���$��w�t���:̽�Լ�~ȸTHe�n����r��=U�f�U���	Z%"�{ވ���q6�<?�����į4�"���Ш�T��<�{;�8Ͼ�cXn?�����+���Ε�%�ENǏ���9����Z��E1,��+A�E#�q��k���}�f^?�~6��5�mb��Lݎ����D��,�gk�&�Y��r�j���d3���2EA&4�ܴ/#�,�W}z�*vUüJ���-�z9�ao��,�5 ��'a���w���op�V��L�)g<|�^�l�<c{�7�����~|Km4|g��YC��Cw�{��!U�u�Ӯ���>�=B%&��jy�+9���+�d]eiZ�/��\D3ƄZo��xI������e�Ys��6E�s�y} �Y&jT*[�w���
�+�Czᦝ�R�Xs�z�{+��h�����<�O�s�dA�+�L�Fh��e�;��S��~�{��G;5��U����w@����ۯN�p�܅��'�,)(Co[�R9�te�vr�4���֖Jk�^�.{��۬���2|�t;A�8Bh��:���8jq)���u�;*��j*#�ڋ���w��͋U5x3T^�cP���s5֝緡�ډu��8�wi~�U�����Z5`���5&�<DYP�	2����ZS���,���T3+ϲ!�s�����1᫠me��B�M�W�`Si�Ƽ��OcW���YWV�[*�f����8�Ǿfɟh��~�}�j�����	N��.M�����k��:�<�����ax�ez?�soq��c�UQ}�]��1�{�Q96�q�w�n�L�%*�ǲ[�2���|���3��eQc}Oqp��s��Ϡ��P��r�ҍ��u�$��Dw�M�ydV�gR1�������w�weK�1җGy�
(�h2�v}Ք/�fq��6��|�[o���	���S��;��,��8,]�@^�1�L��zB���Z���(�7\�yՇ:��G��D�uѭ��m,�����^�o���}aU�<��]vK��*�щ�v=<��5+U�'uݭvLjgI�r���-v�1�w�ڼ�__'5ҵ3��Tڣ�Y� �컴-Ԣ�ݛ��l˥&V��5,7F�r�CYm��)��z��ch\�ܫ�PD�(^?�Ա9\n`�Y'[<��k�7�O�H���GP��u�CL�']]Mrb��o����p��g��O� Ri���s1�ًR�UȆ��5ˎv�ťL绺�Z�s�=�x�/p�K��(]4��u�P��bt��Ro���`���2��!6tͻ]h��݉r�m�{�G�Hq�
�=�%e�f�,QH�(;�2���lD�\Mpߤ��-�cw穷6rs�I���d\���[�&���a��/�ɫ����n���{�"/��m�F̎�ᩣ'sZt2�֣�-��ƚ���9�sI�1�r.4�i;�Ӆ�sPa����%����Ky�)f;7�WM��M�v���
��
'd;�q�6���S`� ��۹!q�zp���S'j�%<hR�uj�&��v��8�fkҖ���sg��j�]q.�Z�x�.*���/���Y8��z�<�Yt�rXI�d�5��z������4zlR	b��F�4�ۧ�̭˧�ݲ1cY�o�.�rsg[�\S%��k�[�C�'y܀����-t���c�@U8�f��C3�P�pu�7�ŕ4�2�cp��(uo�7���ds|�E�J�ʝj܋M��u*1ڶ^�}c�E��x&����:㎼@����'*���$U�/�c�2���H�j�1\��;>V���V�m�f�����-��y�2��0�y*oL���m�ծu��}+�K[���+z��ut��~�CEWH�ʚ!�Qd�f���DJ�C5�5��ji��:j��GY�ZV+XB��L��Шb�2�����±k�.Z�Mj�B��"���%F.YYU+"�Zf&4n\q4�U2�Z�F�ư�MR��`�Ra��±���n��(�R��nT��
E14�:����4*��i��e
���c5�ʗ**�2��2
��ul�
I�������E&5�@�
�aqi�d�+4�2Lj�T���XTM2�t.���)X�-�X�Y#h�+4�0�<�Z�g^?u߭�K8��-��톷d_ɗw�����^*��d�w���\�-I�}�}��"�jI�56����*�f�GE@լ�gQ��P^����g�p�D4�2�͟[7p�ٍ萚���6,.�մ��sЭ��O{��R�T�M�ш>��ͮ�6��av�L)��:�4t�PV"UYB
;W2SҚ���IC�.\V��;�i�9	�L7++���h	��(����{`�=��[XJڬ�{�sF�4�~�7���c%C�._F���c1�	��F����s�u�<%Bݎu?�q���-l���f]��;��e�5��/or�CpĝH�f3������h(�6 ��[;[�҅��e�qҎx�+d�2�ӯ�^�x*k��g�L쳻K�U�4z�[M�5gAWt�ET���Q�w��yoT���T]kk�WV������Nx���F����Ct�	2A�L��]�ȭ胐���v��VA��6���D{���"�.ߢ��z��0��J���k鳺���-�}ϔ��/�P��-u�j:qr���Brw��E�T���OB�i��g���Wp��ߝ����r������y`dN�kkj����8������^���3�z����Y����ךXJ��YprbM��E@�>ތ����
*7��ΜҘWUH���.z��m�Hj�:c�^9Wѷ�VsxYq�[Lv���>��~��ޞ���e�n�u�6f-�G���=Lgp+h�8�����;�����B:t�xY��I�t���ը��W��עC��'��.r���/)Mt>LE��q��S�^��#/��]�3v��1���#n��2����6���y����T'E�:�C��:-��>�J����1m~;X��<n�z���H-\2���Y��gDⲬ�{Z��R��G���d2[�_��j\�qP����7�l�WBі|���i� �w4\�2�
a=P4��0:�v�vD�u$��e����4����q�'�2��(���R�ʳQf:�;�`,�W2����2��.�ASb](��IIR'v�LK[�5�4/�.0���o���9�Nt���I�^=Zg�,,���u�����{|x�Cs��s����z7p��|L���i��C�U�������O�_N�qw4���q��Ĵ��k�&n�I�Q*��;�܌7@�,�ұ;�gT�A�F���GF��\���V�7����s޸����mb�0g���`�U��/y�s����:�eTbv"��lA�ڼN�s�]yb�;�M�Î�3ޓo�M�C�gF�;�#�T�&.��(5P]�͔/H�f��鎕56s!F;�[	R:�_�������������>������i�z��:�ln�Q��&n�\�ԡY���\n��M*3̢9z��}��z�%�7�_�^�}U��R��i��'O�O�w7���<��&u;�j�=�0
��V��M{U�Rp�m�c�x3z���*!�v7��s��w�8O��.,�/D� k�I�>f�)���2d�g;HCg��6�K�d�&����H����e�������ԕ�@�Ld���&��	��֩;a�m��I+*yݒZd6��&�
y�Xm�PāϜ[�(����>���m%|a>=���q�V���u{�N0<��O��C�VC����8��XI0�XH$�N0�!&	����}w��B����D|�{i+�	���
N�Y:�O�I��Bq!�:�v�!6�}XL`a�z�:C�����g\��־�|����ibN2t��Y�=a�6��o��I�'\�x�Rx�ȠC��<�M�+%d6é�!�>Hy|�On����λO}ԫV|\�S����VQkZ�j��,u���L5��ʃ=ӡ�e�'~���K9�<�
�yqwK҄�od�6d��ԭg%�M�\Tu���;����p���/��D{Ҵ�E�s�z"�~ɓ'O���'��=d�'���!�'h��I;d��0�'�0����=M�n�t�v��$.>y�}�O3:�zsǓ�:d;a��$�Y�O|�yd��Iǌ��P��l�!��C�0�ް��I�'g���J����I�i�7��׽k���_�ϤC�y�22ϐ� ��Ԝ`h�0!�k�_�&��I��!�!�N��)�>CyO�N S��z��9���s{���LBz�n�c&����5��!��0� ��(���i�݄�'���>|`=��O=�͟!������2�{��z! ��ϴm��a�d��5hM�l�-���RE�<`x}d�'>{|a8ɶl:��I����Z�}s����t��|wd>a�q��$�u��t�:s!�+!�(�w-�$�O=�
H�q'�;�M�z��}׻������}��_�L�:���'�u�6�k��$�+���u�N2�׶B��{Hm&�jء�2O\d�tW7�^�)f�FK��G�X���c��'O�(M�>OP�	�O��ӦC��`�''��ӈCη�� ���I�O~�v}���o�}�}<�x��d���55d�%{`v�hI�Ĭ!�����O
�o���z�=Sc�IT1�=�k��7��u��˝[�c
��"��l���$��=�x�m=5d�%|`jwa;aS�����1 d<�(m�ާ� m}���V���;P�溭��>Y��c#V�i�ʓ�u����h�U؞�;v٩�1K���������5~���x�bgJ�s0N�I;�~= �+%���ܧ�lR �Dԟ���ﾯ�L/�|��C�I���=`,���!Rz���,�zɩ|�M�k9�u�$�vY<d���8�*T�$:jd6��ڭ��]���>ߚ�BbI�0���l��4�����Y1�|C�P1E��B�6�k�i�VN2�u�x�'��Lgg�q$Vk��L�,�Gs�_̺Y�C#�"#�<ǥH/�:f'*T��M$�T�r�=$1�9t��$w@�I��i
��/����dR
C/N�>=���[
�����.���#؅a�T�H)�8��i�O��va�T��I�R.�{�d�!Ѻi��$���q���*}��1'����eH)�S{�߽��7�����I=@��m�t�PR(t��>�󤂁���M2��̆��J�a��d�+�t���&ЯG���L�2��{��0B����������N��|�澈C�B6����i+�y�@�ACYg�Ұ��[�I<B����P�&�{dӤ��]�㤞�f2|ʛd�>|C9��sz�nm�����7���ϼ}a���>���IY6��4�YSi�Lw������I�8���՞�g̕����OYSh��I�8��ڐP�4yf��q��"+qn�%�'�ϧ~����X�@����u�{b�Y:�2w�&�����CI:B����i �ٞXi'���T*J���H)��;�i��T8����5��o��浾���<�ஞ bOY�U�d�R�v|�L�OuC��&$�3�|�AO�=9��8�q �*C��*8�P=�a�Jʐu�z�l�%B��>ε~�1�3���;�c'L�_�1��Rq>�|�Y8���b{�!�N!Xz§�u�!�J�����Ol
�S���q�X
m:-&$��'V�H(z�~���.{�{�xe�+&-�qU��H5g.֣����|�6�����P��L1L�+N�7^�h��/�E�,�\��tqHI�n��b�r�Vssz�K	a[��R��'0J�8H+�"�D{��)o6����?,�:I��1�fXbm�n0��=M$���06�o��H|����i��T�i�E'���t�������zf2T�_}�|���߼��v�ɶT�E�P*N�����=zH(o��&��q��'a�bAv��Ժ����LR
ü��|� y��I$���U�1���6yW�Ot��?2�q�$�*MwCV
�n0<j
E�^�d��k�M?:@Ĝ{;�L���`t{t�V|��z���bANٯh��I>a�bM�N$�^�~��^}��=�]|C�1�3��'Β�&ӦJʀ�>a�ĕ
��=ee�Vړ���Y�%d�tut��3�=ya�4��G�6ǬD1��d�/h����]} 1��4�Jʬ:�� �M�wa֬4�P�����VjA��jt���c;Փ��q�Y�v�I�f
=��ڬ�J��+5��_}��Y�}k�����=��c:d�4�O��t��V�q�d�q%z7@\g*IY+*q����
�l|��d�
o�`�ӌ�{t�T�����<ä�DD�i�S�LuM�٫���}#G�Agڲ{���bN�g�H)*d�d�*Au��a�N!P���q�B��j�q��c*o�q&�{@�=�1��}�u����y���s7�{��Ϻ~���J�$�}�R
|gy״��g�vI�:q����0`q����c%eI���'L8�IS��i �q�Ѻc���"9�\�v�����IB��Ld�>���0�<��t��V0�ў�C��a㧦d��U`j��
��/)��H(x�a�`V�a�1�Ƥ��gέ���������~�!��&�g�t�:H):�i=q� }�ۤJ�W�);f�;eO�]a:I�+'SVc4�P���Lϙ*u�=eM�l11��߿.��1��;{�������j:7��!�n���+d�A�$^CM�86n���Y��p��'2պJ���I{�s�u�ң8=��+���u=��F�}��:4�2��ڨ��)�{�w��@�2��7�s�ֿ�L���D;I^2x�韎Y1 �C_S�i�AOw9��6�����S�c6e'n�
M��8���j�zϘcb"GDH�1�0�g�G`�o�i=�뿉��Ag�vc�d�x�$��1=����8�ya�X(q%g�h�Xx�� ���l8���S��d�=f�a̰Ă��k~a��H ��%;N�n��|��l��X��H��d����ĝN������m�/�+m}'�CL���זq�a�
�n��i'�<B��Ci*{�O]8��8n�6ʩ>�{<~wz�׮s�n��}}�&!~ך!���e�Oz�+Rz�`q�6�ߔ� �6��>����Ш���I�=q�|�����VOS�ô�$�
��;���>���w��m�++%C�|[1��Y�#i����@�P+2����O\@��8��d��מ�H.�]P��;H)�;ꆾ���(r�����>CG|���]k{��y~�iuM!�LeI������zϋq ��
��)1���׹�_X�}�C�+����B�l��z{@�IY�tr�����sם�������޾8�a���A���i'��ѻ&$=N�O��5ý�
�����*m�وTP���Y�\IX�Y��!Y�%N�l8���D��>������7*�?��(G�����阜@�x���k���Y1��UCYa��
����\�*AzݜIu`V�l���Rs<Ι�AN2w��z>"(G�����w�U�'⒁.M"�|a�}Շ x�3��,�ed�=q*i&$�;����%C�[��mg�Vi �m�Y�@�*gS����6�
¡�J�삱ͽU����.��G����j=�i�AO�;�kt�����ćv�'�����R�a�VM���J��a�8�7f�!����J��S��H��X}�����ܾgG�|�]i5t_;�,blEO�9��:}�>5q.�s�ͻX�PF�Px9��lǰL�r�>�eD��6���"���tll�6VmeeF���U�YF�=��K�-.�ElqԊ�G���z�4�]r����1%}v��i'��%�=�!�J��'O�R
O:����H�S�&3u偉�XN�jEiY*z�AJ�l��
s����q?M}�"�z ��2�����%d��t���#l�2��
�gx�q
��y��|�P��M0;k����N�U<d��
��b)�z$DGY?e�v��R���D�,
�`,�i�i �����8��P�gي�����e��HJ�Fy��'Y:5�M'��LI�<�XAf�*t�I���%�y��������:��x{��Ă���T�z�R�^RiM�m�xrɈx��a�S��$�<I��A{�s=@�)=q��E!ա�g�4��X��M!Y6ʍ�����|�﮽�{�므�x��c��i ��u7f��J���<��}`Vz���8��{gi'�Vq���RU�$��R=�y&�z�t�����I�9���fk1;_+��Dz �@T��#��vyI�Jɩ޲i ��6��I�T��wa�i�ĕ�_P��M�Y���L�ea���=����Y�}PǣP��g^�G֪���7Y?z$@鯌�ZbAd��׹���V�P��*MP�=I��:�Y�����G�~gI8���q�Ϩc'~�P����ۙ��[�w[�IMR�7[F�<�G��H����]T:1��"̮46��d�wVU��
�\8�=�	��6� 9�5�Y�H�Q���^���j�6	�1�wŞ�i��yG�FD9��}��T�I^��<8�ѬU��D�W&��]	�FeuU�t�A����x�	��sC�uD7�e��ڋ��[}�<x�,�N��%��Тa�=���k$E��Օ�[{*JOj�tk2����]`]wt��2G'������ԛ��$�϶�w1�,_�i��Sc�
���xwH�J��}���W�Ѯ�ǝ z�bi�~�a����ߩT(p�(EV���f���eC�e$����y�y\�U3�ӫ>�>&�_]ypu�b��Q�Y�o�"n�{9��.JƏ`�
͌�^8�U�,��(�xG��2�n��P��H�C����R#!�ͭ����X<� ���כ⟚^�l�r���=�(
sΪ(j�S~�T	�1����xp��\7꫋՞�v�JN�qt�+�!\�4�
���J��x�}@!�'��WDl�|�7z��| ܖ!i�ޮ|+x�+Z�]j��ڻ
��ȶ��z�2���u��O*�K�������z�_$*;��¹�C����6�%�h�'����H�D}y����b�WP9�߯��Y��1A�px������*�q=����5���	���6���g=/F����ZuU�jlF�v�B��A�������+48P�n�ne�
ݫ/l&�ne%�nŋ>��m �z�Ր/�J���Z*�ۀ7@e9�Q�uڳ�j�v�tX(@1>��U/�٬��g7�S�m��o���|�~׏y̆����;+&,��n���.�	�������Yvc�٩�Z)�-7���֕ 64�'�b�P������{o+qt����%m��νw�䦱�b��h�ʑS7eL#�.YĤ�"u-X^�o�Ҳ�X�!�:����Q�8����<�gbr�+%ǬV��&s��F3���c��41NT�b=Cv�m�)q���e
��T� �Y��-s�[\]��%��Uso����8���ث�h���xu}l�KF@7�.W�c��;��M�R�j����-�{����	��^!��Yx�\)�*�1�Q����Jg
V(��/s�nv�	����]r��L�z������n���щY�t�������O~9��P�ۖ�-Q9 �O,�}i*z+�m�r���ἦ�P��%8ᨦK�
��J�5՘k��؆��zksgd8�6,d4K��V����,oXw\=�Y71VH�X=��âl����2�
=��q-�Ipu��ua�P��l^�'V��*Y�s!��={0���}�������xIqcܭ��F�bW��YT�*bV�Yڐ\,��k�PR�OJ�v�N�&벂b�	�*z)
�Lp����vhN'q�#K�E�݃gpܾ-�:��+zk��7x�W�l�ڃ��N���S�;x�g����v�RoM��V]!�Lx+2.	^&Mt;�k��F�H5/���P��WWê6�[b/�������Zp��>R/��4Rv�ڧ�ٰ����&6�,�	H���p�J�V�:���:%t
�Q�yD
���b+5=}��v�� ����)���O'1;%�بz
��7����X�j}-wb�GX�.�r�h�t���{0�jq�I]��iܮ��W����xơ`�0\�����P˶t�n�(w7z(pJ�Fk��R��f�ݒ��t�*�}�Rw]�x�1�X���*�Y��V�V�RTU���+�`i*J��J��1
��C.$�f��aF�L&�̪��P1��Y��4��(����Lp�
e����r��e��P�i�E��Q���f���`�c��Q�CI[Z��E4ɉ)�����E.P��E+*&����5�,̦:T
ԕ\eI�14��b��¹������˫d��k�.i�a�XW-*T.�m�L�LJ&5(���I\ն�h�kC4%E2٫[LI������Ʀ&&�5���
L�2�6��e,���Lk1U��je�i���M+���2��ֲk,(��GE*IZ���iUR`�	*�?|����:����9��J+Ә���s��N5ڨ����n�<P�v�X;:�ϱ: �!r~��ﾫ���Q��7��R9��*"r�̡=,eC�C���tV�[�}�̼{�z��=5�Pv�第�S�[�&��V�R��*ָ�|�Y�.��0���S�K�MM)��R��OTT�ܠ�3CJ���[CeY�N�W��^SYu�p!��ګ��%��ϴ=��.�w��>��4��%Ss�3��Y�E9`�\eB1j�G��4��(��f�G��$+�M�ˢ���}�7y����^�*�خq��Cl�ϧ�����B|���A��=q`�<=5Z�{k���yf�~^�x`�}��Ts 0S �	F	�bvuOKП9��qae�P$8R�*!_�:`q�#�È��r:"�:� ���w� X`K��*��ഁ�$ma�k3��.���1�.��J�8i_��.�6@`W&�z�qB���Wi�~G\>{���G;���z��������!+��%�n�xAB��-N�X�`�׊%������ZƜ�#�������>޽�x���R?��)�P�@Ţ�t� BRD�<�vxB׹R$�X��}J���0\�����\�F���
�i�)ͩ�@^U��
�ԃ�%�M��-���ȼ��XgJ��؊��c�ڒ rI�J�\7��K�|]ok�a�'+z�!����C\:�������c���,���j�a�^��sݝO'��ey����c��g�y�;v8!�o"�I��ꈋ�c�Xy<� �aPo{|�)��,����Ȍ�ؤM�$���u�u�\�7�P��ti�.5Sv��A�����mM�/3)���F�j*[�`���>��1�7i���Ɗ�8�O^�xJy�\�ڽ 0? L�$;�[��HSҶ�����Qx�6�cl�^3�0�܋J���TDđ]1��A�����N����;Γ.�]y�͕��d|/�tF�Ž�6�h7uc��6¥N���2�

�YZ��h�	������*�^���ia���w�]3(��pM��s�@�{�lo"�+�����l��bj>�I�*����Ʋo2.�� UXwK4h�*#_�X��-�ȼ!N�7�Ǆ	���ó�#��<9���No�ZU�L���������Dk�ЅT7�ҍp�g��(v���hTw��#��.������w�ݯ�Z���J��˔fb���V� �JPj:���0[�^�e����Pp":B�0:.��ʌ�͔&gD\e+C< ���f̩4��q�C�iR�6+�=D����)[�զ]`�y8"�d�y��B�9ɨ+o���+A��Γ��p��]-�k��ì�W�
�d��ޭ�0Hj{���䃠6�G�r,��8���]��~wԹ3}��|7F'��T;�#�f��p�7{%�ڳ�2���O�ćl��nl���B�C�}�Ç�&4�uЊ�P���� ��Z
��w{�:����p��7y�yD*bWbM�TJ�n���ɑTݣ+�F����|.�m�O���ep��e%��X�]*l���M�͒�p^���F�4�E�n:�*켧@�fFT�G�""Β�n�z�h�E|&4p�0pb�ܪ�-�p�S�=>Λc�o��k�o���C���V���T�Â/*G��s��#���U���c�w3��fS���3�8)��2>	M��T� t�FC4��(#���^�¸�O�L+T��!���b�̌n��(�hOz�&��B���5;b(8��6�b7���bӢ&�GV�ʤlt�vs��Iv@��ǽ�+h���p�~z$�����U*�eezf���O���8@�/1��:[��g�=g	�����
�}�`���9���t�U���0#grЮ����ٍ�W҅*̣I�{����x���=U�F�
���"��0#kC\����x_&%��Fԫ��-�Xa�W�à�r�J��'���	�1��D�r���U,�~Qg�c��̔�m�?*���,�Zw��>��R�갠��=��40Q���T��>6
xV;|D�Ԯ�a)1=@ڻO�2tˆ����U�H��R��[շ�W2"������1I���,�4?-xZ>= �Pܨ����`#:@@���!q��Egۇ�Ͼ>R�dЫ��C�� �6I٠�+�b��,<�e�]���E#1x��tq׃V�T�t�V��N��xW=Ph^��w�T��[z�ԃ��S���B�cF�ڡg�V<>�8Md�O�CB�B�p��{JnΈ>�d���dl�U��i�}r�ͫ]�L�����~�����1�7Hf��J�U<5�����$ �7��&�c)�5�wXK�g�
��L�X|(�<+��V� в�1[�;�sR9�ehS���D�#�P@�ޕ��q��j�F�C�v�8L���ܢ)��Ҩ�u�r"e{�눚Ͳ3�n�Nx1P��ACFXr[�P�FC�D}�<Vv��w�a4�\<�<�狮����i�&T>���M��-񈞯F��ֽk;��Y�ເ7���=B�'9��LY�P�㺽�ܝk�"�*�N�����N��g�M@91R��Ċ\��z=�ܼl�w����t}��� 0�cE���=*,����)�.n&�ىM~���^*2��y�t��uKʕn��H
��_Q(h~5,NȾ�=+�v.��R����q4+d:����4w1Gg"�u���n2�r�n�#�H`�*1֊���XPѴ8]i��Xx�����E8�W�yrСQ<ӷbbS�ۄ.+��9/��
訹p�}�
<t1FR�p�k���7;.;��(+^��y�#CS�(��x�#�yt���_��k�eh�:��G�"%�^\�ób�8 ��(�=���OV���#�4�7�׽�������hp�(.&�]M�Cs��s��W4�/��j��������0���P����r���FS̗YF�(�\���^W;����W<:��B��f�B|o{}�j���Ƴ�m���5/�6�262k���L���7t*Y����*��L=p�e�u�T'V_n���`�\��'�g��j�n��.#�M�j�&��I�]�7s�4=���	�&Ƥs������t��W���."�����o�U�0Gi�/U1�]��4C�&r�vkxkY-���:xEЅQ���`Z�
ȃ��,�LQCy��+s�wk��Xp��$ k�H7cDp�z�N9V�p��J��[�)pK��w��^���2��T��}ˉ�h_:���;�H�56�y��W.$5�FYW�Z�����ƱM�D� �t����k#�(�㈥"��я&���Aߕ!b�xED��B;
.܉}�r��Aҳ�;z�?��
��=(�	�#�=�A!uT
�&^9Ήi$V��fh��luc_E��m�^&���.�вB�f�A�vo7IUY����q#$+FG���[7~R�J�G��U�V�.������ ���T�tV�YԈ�T+|�E�2*�p��|z�Iq��~x6����-�)�w-��b��*��t*������O��c���y���"�۾���q�uٲk4�H�;��E۩��ob���)^�r[�O�3u��gw�rO����[�y�':��wD!j@�J����ONx�L#�Eѵ��l�2�"�|�.������8����@���q����UֻF5�=1�,nuh���OX<T������TO2�~9�K%�0�u^�f��
�W��&g�;�4^ �QC�G]��3LuЊ�U>��H0��
�
(��ץ�F_�ɢݛW���)���3�U2��{&��t�v9���X�����ݡ���Oj��Q=\.�V��E+�u�J��-��;�QM�܊�����a��GN��*�����j*MS��k֘���]��W�L�qQ��]pW�O�F)��:XƮ�[�2�L� Gv;����� b,�%*YС�pr�S_�*ỹ*8|��59���^<�B�3�-�w�}{sD;�SX�nn�@�4�
�m�q�\
=^�*�R�-m9{�i�<m�t��7�n�N��I�c]��]c�4Z�s6<�y��_i���d��������RN],���H��mT����R��}�E��)62P��z��Z6���k|]6p�vx{&�Uu���A� ;�:w��=�2�8� �� �htn>�����ʳV|�.�s�;1���6W&�e�d;��nAu�v��Ȋ��сZ�,��X<
����ͷEK��ŅRdML�s�@^��%H_��r�>P���4����������ܜ�k�$dm�p��P����*���L[���*�n�~����+��t0Dz�zy�R��A������
�M;��G�Nn{H��f�O��1*����V��NU�V�ÔN��x�w3w��=9Xu]��^�du,][T���ו�:?c�)�w�9<��On�&<C���m・Ȍڮ��T�.b�up�S:g/[��6tX��5��,4T��Y�t�tsub�MA���+.{=��uH� d�l㋌p]A��.�ڕu�u�.���g�{	Rm����ϴ7��Ӏ/�PY0�l�
�yVa6�.����iM�Msz�������3�`���G?>���Q{� VO���t�VL F)y���5Js�@+`�,���*���c�<z�xv ��(B��;%�8��8��6��������
�N�Jfp{	��!dv�)Q��0����TT��?/�X5*�Y�^^j�Lp�Ww"��p � 9�n���A���9&}N	�Ήa�gf��u2l��U���!� a�T�ԩԬ�W�u ���7"Pw�Xj�[�ø�t�b�yL��%XB� �3@�<#��V��J��x����m�>�:8V`�`S��[f#�z(����f�L>��L_K�F��h�3H���<Mj��`��{����Ec�u����QN0p�j-.^<�`i����}��JkP��:�g!(�İ�'o�9� ��N��)�"}��Y���B+x�1�Ow�Q���e!���͒�(�}��&T�����mޠ�������WN��-�y8��q�-�u�om�Ù��N�,�����KC��|���w7
�{yj�m�d�Q_���C��z�аksa*J��̒�r}�X=\�Xd�39��A�X�3���e�{-vSc���.����f�$ ];��d�z�A�R(�2�nы����p.QU�֝ٔ*_1�F�*"�t<&v��a��[`n�f���pz�?9f�ǳ"Y���b��P�`.r��2�ʴ4V��,e٢�EKc��JRc��ܷ�;7`�Św�)`�i�C��x$�B���@�kI��(�]�hQ�<{���!�sb����(./c�x�e�=�q�L�:*$�7�O�NP	��rt6n�de�[\��?�jXD�p{��)�4qg�J�J��.��0�;��2!�r�F�p�����`o�eb	(wn�v��|�q��K��`��}(�F8N0G�,xr�d�M�$H8�K�YN�L:���']ݏP��`毜��NHyL��䄻�ُ%���#KX�ժ�\nK��8����o<.�RҲ������!�e)��7�0��=Y ��;�M�{BE��K�j�oU������}a������=/�,U�DR��c�f�Ɣ����hT:]��Q�T}���(�G>S)Mx�9�Nt����VXU{�R��P̢/�֚=�u��ۏW���4!��WB���;�`�vIӒ���s��8h��s�9�%�c�uI�-t/6���}���]v��.v3i���\��^^�E�����Ckvޓ��yY��6u��>�r�!�����j�ל7a��b��ю��]�;��D{���˿t��ʸ��w>©�~z�������u�!ҋ��;�ך�F��e,!n�&����VC�$3H4Kj�.���aur@�`<}�+��0G+�Yn"�Ȝd-�uyQT��&=.�T��}W��w"���u��S�"]��b�Paؒf�)$�3[���6rl�J�Qk͋U���ߝ׾��nl�V��ObxԶ�j�2��eJ�	��!�b�JV)X�UˎW�Th�B��311e�2-0�mV"�
�)V�,�2�U0Kl+�h�mLa��T\M3Y�.�q���Z��bU�a�bQ`T�V�QT�r�P+���Z��J�\�Ʋ��8���fZ�
��ʅ�P���(�JŒ�°�QS��U-��RiәJ1[h�b01ċѢ�ŨE
�E�mej�U�Fk���V�kkh�ˎa��̴1�c2ڭC2��1��C-�E�Z�*�-J" ���-��[`6�(����3 ̪�-�2��qS2�V�UJ���Y�� �\�uj��PU�9Lej�����a��R�-�TW2 ��AV��ŦQ��ص���EUH��G�C�����Q��=~��������)fǵgrW7o*������C��9�,pŃ]=�qȤ�����Vr�����1�A5#����oD����	١���,p���dƒ��so8����r@H.X�-�B}Q�6V��i��Ce?��__'{���Ǫ���Fc�8��aS㑹�P���m,�TG�z���Kg�x�`R;��l�^ʮ��tm �r�����3K���Rc3�_fnwr;>&�e�Ҡ*.x�L��P�i��Li�hq�H�5U��nj�V܄����U<lr�[P��}q~�1�)H]c�U�;u�`���8���{�o��D	!�7J�����[��T�6�r��aJ|�^�6���t�b���:�;܋J�ɁwLp70�́���Z()�4c���q�:]D��#N�0� p=&bb�ȯ�kg6Z��TH5801���,gK*B�����A\hF(�͛����
%�(���dؾx&�L�b�SN��Ӄ���N���͍g}����N��e�\[g��q���^�T�s���U�&�������s�m��u7�5&F�+����q�.܃#螻�]]S02j�yp�5�a��GgڴsJ�t�j>�����ceh4ܩɖuײ+�r>&�`�m�@��#�SS�+�ܿ{3v�p���44����
ၜZ�z�A>�r���V��c�H���:�,}�{�*W��XxW�H���Em	�au��9����t��T*���
WLZ�R� J��Id��}!�(^8e>�o9�������Ǖ>PzW/��&��eq����~Uֻ����#f�	��I�e�ʀ�u踊�/X0*/�e���]g�d�L�s�\��1Q_���ܑ�Uz���	��tGC�C&c��]��P���!�
�#H|�����ɗ/�^��`���{W� �����7�^B�wM�d�oA��I|��ҵ.6}�Qt��Yj��L����X���,wwJ���!J׎�v��6�'@�\��i9^�Oo��J��
�48��E���`�"�Vŭ�n�g���ɗ�Z�A��p�K5�}�����F�֥��tj��f�������F�\��z#Эȶu��#g��5�������v�UP�	��l�I�]�Nm�����W����u�|j)�.����k21�s(1J��2wi>��l� A.�!�(1҇E�1q	�j��k�{���ۮ����5��!��C�I��^x�g(����y�*��bƲ�\�X�][���]%���8<�=iԁ��7�8:[��l����D��.�X1��G3��]b(!�ɟ�>���ܱ�.	����|#Ńe5�՟��<\�ʷ���,�I0Ԏ�p��P�C��~$S��Q�Z�,��'�F�3��ޡ��W���/�D���^K� �A`>��e.-:����7dy5X4O������Z[^y�H۔$��'qFz���g�wW�<Y<3�A��D��T�T��?
U[��}�֘;��/a�U�B݊���?�P^//#9Ѹ=u7���uΌk�S�5�敋e��1M��3#����v����o���m��e��֧#�tu��E��u���`�F���3�v�D �H�%�=�j�%&��\��;�AyS�]>��E�n�§�}��
�����F�L]o�(���wB]�Dk�V/�j4[�f�D�\��6h�}���~�����ҹcs��6�y٥ӎJ�Ӿs�;׃!/:#ev06b��p,^�� oZ�efij8�U�%�;%�l9��Y
Pv�犺U:���MA۴��:�6�l��6Č ;U�yQ�)}(B*{�k���*� ��^PՅzyy��9T���2����댦!猘p{,O>o�87���;|ʚ��<�d�J�\5b�yw]T�A�P�Kj��;�0�w���To�_1Ō��t�4Dۻ��u�N�h�3�Wc[�R��fO��d]�e�W,.-��O�I��"�x
��X��!� a��+B�����,��bnr���SP���u>�P��71#8���� .�h�@Zp/�CF�Z����>a�NeC�������w�\�ԯ0��A�IFW:?e[-VW��õu\�8��y�s�&/8�lHM��k{�q��q���R�lӁrXVL�X�&dծaH�����+�p� �j62͎ã�J`�V-Ҭ�4s����\�ά��u�r*�\D���4�(h�
r����&��Z Xꁗ��3�Q�eihl�3�e]H��`<�ŗ�Ç��>|%x�>f9���n��-�T�)���#t'��P��[��>68WE��{�b�w=P��`�ۑp�a	�dS��l����8�5i��b�@����N����Ã�?mF԰�L T�3~��u�U��D�p�z6��mS�Nѧ��ap:2�6c��T2�i��
��S�O�F�*�g�b�Me��,L��e�v�E7�4�4}��U�_D�V�ݴ��Ȇi!k7"-B.�gIK\���9��`�����U��)���ɘNa�4��X�Q�v�����M;A�QB�Z��N��*ƃ�L�/�a���1��:".�]�"v�-�)[�¾^]����h�ҀF9ZN��H�okZr�r�C�"W��%>Ō��Q�w�q:!E�|�n[�:�L޵[˂��ʻ1��8_v~�㣰Z%"�ދ�ծ������S��Hhm�b�	 �	�� +��^���v�]
fz�kL,�S�y
���q��3��J�&}ˉ�hTh�U��Ahq���x��Q�6��{��k�z�t���u�(Glb�/@ p&{�hC��68��B����G�!���Co��j��"8@#Ԅ3:�tye_3�d�#Ն���e<z�:f�3O�{*�ΑR�	��"����] ����d1�P�T��+/踚��}��$ӻ��/Cu�*6nT&y.�)�U��!�Ϊ��"2B�`Z.�=�;���(L��hڐ�U�RT�êV� %�5����B�T�.e3+m�m0�96�+���������m�
p!c�I*�%���E�< NS	mh��h�S�3���Y+f$M5cҫ��à	U�wU�Ƴ�~]k�*tn=���;�2�$& ��Q��v �o�u��Y�.�-���GrQ�d^r-��3��Tp�WhD�����]2�D}W;�թ2�V�Y��t��M����'i�jC�/��������N�E9H}S�:��VT`^�ϕ�%��nW|��vI��׃
���9Q�@1wE��¸eD�6cB�ӕp粁�m��{O&��( �֎���9:8]��h��"�+�<f��^CX������-�gi\s�o�8�3�G�k^%r����H8"��Z�Y�OJ4�m��#.\d�V_g���Y(>��a$�3 a)����u�b���)�t���{\F�!���B�{�Lqu�,cWq�ә@U�o�����x��G��5���ZՃ�F��7���0��=
��[�j(r���%�r��7"ԓ71>�r�S"3���핣αW��X�H{�g��&n�8�wL0��.��H��.������^���p9�}�B6mU�GTQA�&(mϹL��U��lN塗ح��Y;��q�h�5iU�5PV�w9֥ۨG��x�8FT�>�l�,0A+�&�^Bh��m,I�3���X�K*�շ�3[��ϝ�t�aSUpi��v"�єy�u`��j�]��l�!K�%}���R�M��,8���H2�א�#���dE��p�ڂ�S	k��vew`�u�=W�AQ|b_k�@pXC�ʣ �ҙ`25ڬ�&3���{0'�	�o���'5��3�t��R��
���4���z�YC�L�{D4�|ŌrE��Fb�;b(��׈sYJ����"wr��/�,ʰnOM�Y�zټWD�1�u��UO�����1-�=9���	�̠(!���F���=Fvc#�0Xv������wgx��T3�K}�`�>��(:�5��V���3{1RԸٹ�l��w� �48ʮ�h���>Zk���WJ�Bn�ĝ�&����*yc��W_	 Ⱦ�u�TpJ_J3�^utC�j��^�T�:��=�֧�� ��<z��S��A�]�G^S��u�a��U�z$|v�}��,�q��tu�νj⹉�2�6m�7�G��7+i�@,�	CN�x_�����@dh��qr�'ۃqk˩/�]�o
N�]4�Nܙ�3ä�<�-��I��
\���׮�y<H��Luq�)Q>����)oF*:���sۧ�Ӧ=S���
�͐�Y�h�@�w�=�ո�s���`>�/a����*[���1v��|�U��HOP}�Gʄ���=�k��'(�9���H�/�xe�_��W:�Z��mr�V�0P��@�</9�*RoV��!��D:������Z�-(R�ܱh��U�f�+§Wv�A�S���`�&�/O�GN��	�
�U9XI����xR� s��°gaΛ�rJ������D}o>6�A澊)����R�>|%<˼т�l[M>˰E�>����Q28��۪��Y��58����V.ߎ��"F����Be		+�m��؁Lh(NMg���j�m�\�]�qs����*J�3m���N�HV��$�I�~���U�[u��u�7*f��0���ɀ���xqֻ[�L:�)�׷V���{K��`�5����3A��|����3"����)�ݜBd��>Bم���Y���]+��L�����'\_�OXZ$H��Z�x��fc���O�>9���������ޏ٢�!z> ���!ʮ��vJ%C4�ȘA�őJ�fnO@���|ES��N��!Ri;hSG�
��0��*��z|)��Տi�h�m�ݮ�[$0��7",�P#C��V�]��[�v��"�^E+]T�X�R������Ƌ���$ hI��Dp t��$�ʢC�:��P���Xo��Һ�!Jk��K.A g�`���+S���]��'/�I� ��ƍȔ���=#K��]3|kބ:�� .*cg���U��)�{�u4k1Qꚱ	�����T���Lp�������W�*�zJ�
�^����kB�m�,^F���<+ʅK��e藿!��*a^<�6Z��x��_hT{�GN��ΆGT�K���� >�|*��ަ�7~�M>�l��,�۵&\Bn�حzrQu��b]5��w&���-Gwsl�G+'L�WxV�]G+���*�Vĺ-ݣ �3X�Sa7��Ӕ����5�������X)Py���q|�%�z[��q�n�������K�#[Ե�z��MIywȓB�gqЊ�e܋F3*	E�&�J�L��\����v헨 �[SB4��'r?a�ݕ�l����;���qSQ��f�(�۫&l�]f0fq���6�@T:zZ� p�TLT7����U},�Dgt7�>e���Dc��9>.�խ�)-ѱZ�t�ݑW!I��Wa���w\����+�����2�ӪE�*��9.�y�U�Y8��B��9R�ֹG��-jS�v�]
��x�6g/4���{u��uz�k�Q�F`^M������v���fur]ThV^�F�(kyX�ڸ�YG{��cX�U�K��"�͢�b���7Y+wou��yޮ!�wʑ�Œ:�r�����|nc�_M�
,L漋��٭�S��cj)rK�mm�"�����PH���^�w���/R�{�c k���,Ve���#r��:�dNк��{\�M6��R��Y	W.�e�,��p��K��t�C}�
αP�g�9�I-%.7GWvD9���89�\�1��$�S��WHlE��f�9��
7;�gX0�{M��ʺ���K	Ȩ_!wB�5���pM�ڠ%5��n�8����ԝ|�[�9���-)�gt�-���\.�]�ʸBNᩇ�ڷX_ �m�X�ҼuShM��:�S�X��ʮ�8�"��+e�R��	T��gi>�ma%��6�N�Bh� 7�1[�*���v�5�G/&��o�!*+�<-5T�X����A�w�w�D�[i��.YI��,u�[�gm��3�S@�->��3�N�+$��FN�7j���1;���Y˥i][<��\y.�s�V�Z�Q��aI� �촜�m-��r:�27W;��J5B��%��n�yA�ٔ$ҍJ��k�OQ���^��`����W
�2��v$���'�=
��7�fn��G�b
ٚ;�s�n�6k����0:d��[TQ�[��5Z]�U%El��E�Q�Z���R�[J�1��Y*�.�0Ƥ-,Z���ES�&$�j4�eB��&Pċ+Ps2E����2�)�Ն+1�bT4�*&��N8�*�m�+�e*T�0�*,�d���@�*hb�e���P[h�-*�*�
�k����ح�.X��+�G+��*9aL�I��Z�p�3.3.aV�T�6�LE��8��l����1+YXVkY��K"�B�S�R������-2��1�33S�#-�Ҁ�9LpeJ�j\�e*8�0�,QEbR�����©R*��X�Uբ��F�L����	�$m�%Q
 򔠏���=��L��� �׾�eyn�L�#�r����1M�3�W��x�Nlg"�%�Ӛ��a���G��*�$ph
�����с�š��>���Q'��4�{�{��I�4kW��L%�G!� ��@���C���"��~���h����)V
��Z�4yUEd$�zr�gL����i���T!�z�]enIܨ�M������/��H:oD#��'{�%k֒o�A]��W���.�[�"��8ߋ�U�Hr�k�#�PX�3	L �/����!��naU<h��P����>����EK�IƤ��wcWw�C��`�r����D`�¡�+�
����:&+�e������Xy��-.�����pa�ʙ�0((Z��^�g��1!�VE[>���lU�y�;*l5�;����\k6P}1�Ӂ$킪�p&���f�УF�o-���s�I��釳�	|j2�Y,W��Ⱥ%��&�j{��~غs�NC6�����3;7����M�P�c��e!�|�uM�,0�'�,a�xn;��Xgf�mv��h���UQ��ѹ��&�E�59�O�f䨷�2�a�̌�?z,��u3Y3��L�
��U����bx1�(;����w�ŧDK̅'�EԨ\o�/��{~�ְYA����Lx*wܭ��L���wP�j�CǶ����&��T,��|x|��Oъ�?����õ�����˓p��n��.puƐ�~�*�*[��u����D�htnZ����%���s���zW7M�Տd�~�"��U����c��~�R#énJOv�Iy����
,8���w88m_"?8���� �<�ʅ�<}J��<B�:�w�=Ew�/|`�K*C={[���m^ۤ<�PhCbK.g��e��Ļ����/��e���H��H�(�Zt�(*���u�xB���wv���]4-����V��1�u��U(T➯��bw�yy:�?_qPr�F�P�P�pk�h���N,�GJ��Q��{��/�r�J��{�`f�کڸ�·T���Xt�:�m��e���,���2-�v�v��:.A)�Z�ws;�<s����L�<���}
��,=�`I���/՚�$�ZR�=]�RN3�}�LϮ1W9�rT���9����ĝă����a�����W6'��݀$��Aʮ=$A��+k�i��R��g<Uҩ�n�Z���Ւ����'j:v�m#��}��g�^���
r����R�N�P�W�C�6
>#��г�@@�@c�!^QyLB�i�Ν5���thO+�sW���-�1�����c����ڈ���*1v=�ͮ�WaŚ���B6��"jDp�@��jE�{M�n�U9w�Eqz�
O�?X<���q<~+yV:;Ą� *:��@�n���Cj�+��@�N2���QMo�}���51#T�U�%X4q e�`J��?���b�pvn��z}�����+ }��t�d��'�����=�W��:̤}�������^9XI�[�
��O����F���}�H+������vT��{jQ�1H����Cjvgf��C�unM�Hh�+�&�c,��+�Z��THC�P\30�l i�2���{vj/�D�Pdb)K�z=�]��{��F~PՄӮЎ��#�ۭ��R��<'(����(�&��8�[}��à!�"E�W;<�d%�;q8�����#�����lqwɹSn��R��Ԏ�CL�"�W"ʑ��=Hqg=qB��{���kD8�"*�F�I OL T�)�-���3�*��W�k��EQh�yYT�`qSAІ�I����AWJ�S㑯��5�bS͜_��R�����v|������ Q,��uk�Y��\9 P>���[�Sډ��lFA:� �I����"� ���~Uᡬ�lN�j9�}�UfP���$0���r"��P#A�.x��+NQ����]���f7���1���� 	 ��� �[z�;��Ɗc�,3��YO���WT��![�ׇ��e��@]+���-���g�=��>j�AsLۼ���;�N�sB���O���h{4=+��}����E|]���Ύ�]��6��6���P��x�cm��L�edt��Ywb�l�:��W��{�E&�or(���4F���)�;:�k����K��u��5�oBf��pQ�{y�  �.&&7�$,�ք"�gdM!��ÿ*A��`����r�<��{�~�[�S�\k@���<~F����W��}�2�B�Z����/�4W^XO+G_���Q�0W����sQ�n�"�4��������ޒS��D@7!J�Q�8O���#�V����K�w
/Fv)c⋋���{$LΈ�4�xx�� ˙�Bܢ�s(�;L{b�_��7��Q`��8j
UgB����p��K����U��z�t��g_�y
��3tyEp�4E�P{��t���� 5Pz�t�cg����X>�R�V��PSmh�#Hhu�~.�W?�e��s�u�z�y�cE�U<�3q6�˅�/�U?�j���b��7�D�
%Y�����{�3RGZ%n0H�|�	�.PF��\���r�겲���)��m��z��zb�u�].�f�:��Dm�ücV-A]8_+*�z2̧fZ3���v��;�"�\�^to>d��=�Db���`���Th}$0aJ.5��R8`�HO�WLP81�S5�;�s�p{NK�ʯ!p��\�잟g\+!�R�
n�N�UO	��Uh9W�J���W��`3\7�ã{'�Of�Ug����I<cUT �I䮵��٫���d�5.'�*U �Da4�ل	����Q�c�����&g5�<�M�`�+�^@<��rR�y�/R�&����������B�i�A���g��Ns�ļ�u�+�6к����T�[�:��M�~5�d�#��I�P�GR�@�T��=eT�e#��.o�sӴ�{o�ޞ�-B�C.@���$=�r�S�ܱ� `��ܴ+k�ݽ%��U������f)*_ay���X�kֺ�v\��ȦKiڀ$��ⶲ�\X4_?]D��Z�఍>'쯑^�z�H�{�F����S�h�P��9:[e��^��FnD-�j�g �7�1{s�7>< �j��X����jjS��]����ՇC����ع����T{ݙV���9R~UW�Vi*G�:M��6OY#��^���C6��m����0����;|Y0�P
�Q�Xb�&'D�۔Wƃ�CD���Y؅�U6�Ӊ���y���e�=�k���˰��Ȍ�zټVO�pD��Z�4�h�ٽ\K�����n!y����z�����X}�z���GJS��{�vֹ����Q=�v;3�@�@�x|[��{h[��𻼷P"���}�=��K�yh�P��q�\zH�[Emd9��H �#~�� �m��Ȝ�pz�S�*������h=
�7p�2�i�tr�{M-]��W������S�=^�TT�`0�.��:�����Y���t�yw7sY$6���x�,+���`@r��F^�!���k�e8G*!Es�2�A������͐�u�LV���Y۵���El�Cm���/ə�BJ�����^^ǯȋל����yX^�+cY���W���Rj����fr�H۝��A�l|��8�Ktr�ʐf��:�d���-�����������Gi���Ͼ����T�������4�S"̀3��==�{2��%�V
1�a��Q=��:�Z��*nm��{�f�q����~"�(`�+���o�J�\V�B���u�wo]p���N�ı}`E�;g�,�tE(tX�^���N��U�n`f��Q��%��\���ڠ�r�k�	ֈ��Q�Z5��E<k���ة�-�<�,��Ͱ���*H�T�G)X-�s��Q}���Q�o���}UN.��X��a�Zx�%r"᭹�)��x���or��0a����4z��ƃ��T�Kpu@t���t����2S�2�b����	D+ e��o����+�`ש	g��P��d���',�'yIxQ�z�k!��j\�Vx(�
vpV:�ì瘖V�~�ӝS�A;��wX��$7F�';'X8�+�2�K�'p��5����s8Vy\0Ey��7]�W��\$du)��b�j�u{r� �0�x۩�rڀ�&��`�״2;��9��}���ܺ���*7��j����5�D�*�|(� O��.%]��k�����P�����Hit�����ȋ�$Dh"\��@5x:1p�L��F�q�q�G���LC��cCo-� �à{K㻷�#�W  s��9�A{��{ں�ny
ڀ��0V��NL�:Ϳ*�O��j�қ��bpWLh���đ�l��.9��1~N�e�`$�q�}��-��u@�2 Fꨐn�C~����XjP�q�'�	�4��	ftC���;"0�@r�"�v�_�������2�>�����"���o{I8��\��hm�!����]ɐ\;."�+��Թ�"�SEl<�W��eB��6�/i�J�w_.������E�09�/�$��D3����osOt�|a������5��C�+�V��ΤF�����M��#U:� �]��
[`eNw4e�ow�&�C�5�`r[Xk�y��u��CH0�g�9r
OV<�N�,^aS/"�b}E ��|a5m��gs��\�eŧ����%h���=N6ʷ�ą=HOOSb��CUcC�p~3H�h�4}��7��o��^n�C�邩�pP��Z�;qR	ꃧ��4 ��N�^�nn�\o�=��]kI��l�ťoF��S�j�����m���W��A���< ��Uzj��$���r�+Ƽ	om;�ٳJ�i�Te�ˡ]B��
�b��^�I܃��.G X��g�+�cL�O�F�߫B#{3�^�����g�?Lu�G��k�|�_*@#݋0���ݫ��Cԭ|����޷�ң%�pW�O�&�1�zN��Ğ�=f��j�Q������zЖ�1��AK��� ���nD�ٻ�R�C=3W�c���S,B �0C11�$Q�$nާ�V������5�3�6���V�_

�1�N�վ#�����7�쥅������Zϭ~At�]iu�:�ZL��&�*Z8'j:Iw�5ݩ4�.T�hE�J��R��
�k��[���:�qJ�!��/�"ɴ�?�{t;2`xd��C�[�#��8��WtR��ڛK���j��z��Y�MF�3pi�Vr�=Z��[r�tN1K��ϥ*v:�&�~�یօb�CO���sѲ+�,�����(���'2���B/5�Ħ��'�r�򦱽�ȶ*�a����4ݧH��6{`�Nō�m;��M��t��*;YPVp?hx��yV�Ӓ �G�r���a]d�;/�t���}҈m-԰ګ5q������=δ�;OG $Z.��P|Ι9f/�z�n@��O\G�V7׃s�$\�����a:�Z��frTuQ�'��.���(Q{&wVl��G��3�r�mǆ����Xh.���'3�R���TU	�X�����ʸ��7@ѣ}d�
�M��΂��m��%�{��O���\�k�'ܚ;�h�SS�_hB�=Uk7/��y#��%!�]��b-��{3v�pNT9[s�e��m;	�&tͭ%Q����+.U�4�M������s��j-�vB-[&E[�\��t�Q+n�z��H�X�l�����3�&����Tލq"���]ލ��c�C���F��.;��c{��� ��s �O��T[F��$5��z�f�5�]��[؛n���v�/8-Z���Q�nα��ve��<��e!��WKF�Y�O��|t�7���nFu���E��yu�pS�aA^ Ó�ƙ�y���͝ݻ�͝в�\�mb��,'�!��i.��_5����K�@���T�drgfI�V��+OV����;�Ug2gd�3$���jIʅ\�z��EN��׷��A���n�R�a�m�S�Xf��[��8�K�}z��4.9z!��ZM��Ԭ��4��!v��7�ِG�ڵ��.�R��d������sv���/-�\�犱)K��,�K� y��	 E��u�|�=�Q|�VsM�	�5O��a�쥙g�w�W��gY���6�^1>bc�-�rXt1۠&���1�w�R�	1�Kf�i:z��=[��P �D��B��AV؋2�-�T�[rʕ(��kc�TJ��C
Q��TAW)�v�4&e��1Pm��T�ċ��0r�X�J�F"DC��V�ԊV�cR��X������EQ[b�2�bW2���`�2��E1
�k3%"(�h��,APT`��5j*��QX���D,cb�b��$U-�R#"�2S�[�Db�(1�iQTU"��̥�D�(e�DD[j��
��-�b�ŭ��"���Jʦ��SI���DEc�DU�*l�QQb#X����b�#YQb��QDQ#�*�D��"���F#A����*�+G}�����}{��y�Yߎ��]:G�����ش��#�)������Ё�2���T���}M9Y�_�{S*`q�8Y�=Qf�Du�ڂ/�I��f�N���w���}>��,�i�u���H/�ץ|�Vf�/Ǉ����1�u׍+�f_`\Ed�������/���
�"��O>������{Aœ!�����؝�1��랫�[����T_A�����u��O��������쐷P'!��у�\(���xq�Qܗ���Y>׽����:��j�n��8k��O�b���̋	!�e1��s)��B� ���>5ʵu�;��De�'腪�b��څ�,�7��q�5s�����@pBU��n���T�� �����©5�v9kfl��,b}�~p�����ľ�p_�猭��>{�c<����yXNd
m�J{�ܙ�&�bX�5�4�x`��Hs�>�K���Z'5W��ȍ"��oP�Σ�B�Œw���� .��1� e5K�y	��h���3	.�j	���t##�r�*E�����[�w��V��D������ݞ�Nb-�#�����V�I6�}��O��,2k����x��~������xd��⑻٪?Q-���>9��u�a��OW�]z�x�X��GvM�Z)6ҵ֬yŪ�8A�����";��lLmF�� !���hK�)¤�p���ͤ6-�0��sB�Wr.7#�� ��d�e�d��+a;����a���`1�ܦ(�L�Ywo�b���־�J|i�y���ړ���
��zkb��^��x�V�PnL�#�3���R_	�u�@�h�������h���1+7E�ˮ}{͇�R��47�P�]��4��(p��6�+j�3��qa��B8̌�:Mz�B;G�T-V��|Y~5�"�T�uٍH�u^2茅$ EÒ=MM�-��{گ��<��__-k�V���,W�"��:t"�YP@Z�����=2�&
=�N�)b�ۨ��rQ��]_R�qɉ�,C7��kI�z%0>ћ��Ó�F��#��۰ ���1sٓVb��+aE/�"�4yO�ˆ�����Y�K��p����%r!��/��7�R����J��A��a�LS���\�� 0V��a{��T©�im�[���(�2d�
��X���4P��ǃ�?jă����x����`V��j�,�wO�����U�R�o�D��%�����!�a���=��,���~ޯ�ȘAѽ�ƴ\s5��V�-規�1�i�0�|�_{��1o�Q�r�v�ج�~�!ph܈#��8U:���F������e^ �cC��}7�\\���,C=Q�$�@�I�z˓��r^��c  �!��{�jKه
ts�S��VӷBv����z�7�&=@�C��1�!�Y���:�k����\��u�;��!B�i�%�Q�ׇ$^�#�3���A���C�H{,(WU�����*9��� >�{\���m���V�Z�PRD:�I����؁'�=��C��5A4bڎ�b<Q^�V΀��u%z�;���Lc�ׄ,<ݘlU��9�����ȓػ����U
!Z}��9��hk�/#HPe��^xn�K���E���uQJ�.w&@atˈ��!;{�����i�f�5�f���(�6F�u��W$44Ob :0' �&Ono� �<���f��tUCF���(}�6ꣂ��gq�S�Ψ�Rs1��\-b��,!!�6t/�5��� Uh}�SiD��읒"/��]fK�QRKu��: :��>>��:�,,x�sD#� �N����ê�D��8��AU�jQ�*�&�{����J�xzMv7���*��:@A�>&s��V��u��1E�ٙ{�Wr���q5"3UC��a`��]H�����W������O���C��Sq�^A���K�~VC�t�\��y�h�t��"?N�PWc��M��Q�wC=�K-K2�沒�F�\f�WJ�݄o�n�B�e��z72q�D�DҺsJ
u��d{bU�9:��KV(��C3��ʇH����̎i��"���+D��&P4������T<=f�.����y�y�(��,��)��l�D����!��T�t³O�C|����3��L"�65K���d7.e0�L�q� b�5����>�#�F�^�������](6艸U�3�
�- ��C���}�|Cѽ����M7�5�ߕC��v)T
4��(z̀:H�P@��y�*�O�=�y��,����@�%�.�4��}zU-T�3X�(x��v�"��
$8��#/��Ƽq;?_���e%J���W���y��h�r���Dɑc���˫�7(1�Ȃ���?j�P)�ڼd��ٽ��0�~��$*�@����c��W
j,s�`w�h�;�sIt��O�wG�K��;ڨ�1V��'��EU1<p]CHJ=qf\�����yB��M�_A��ڊ;ٲ�����������оkmu�v���>�j��&d��oo�|�d��緆YNMΈ,"�P��E�B�B�]⫼��D�y#Q�+;���o-��S��Ɩ��H���z���ڂ�9�0�)6apݨ��v���{+M�Q҄+�X�����#;���]샥%5���i�J����>�O:������>�x�Zbpp|+�o�d3�sw|��D{�h�>1V��"���F�V���:�Im1�d\sX6��\�{Y@���t�tsu.f:��q(W��P���0-�`�%6髸�AŚz�L�i�����$��z�^�^hr�%��=��₻�o)�s��oi������X6&6��ro4���|�t�I�[�qY�FE��-N�sE*���~�PM򍌾x�Oq �^�k�+k"gǶ��=~�NW9�U�*�����ri�O�.�H�S=s�jVFV�}H=5�>��;�q��H�*���DC(��3�Ҡ����+&��{^�m�+h�17uϗ�]k�/Qcr�AB�5�\�ש���Y��dr�1�%>�3Z� i�k
�鏦��h �H�sb�J�[�x��9�6�"Ƅ"C��i�i
�B���!O�i.��U,Bk��^�ڀ�i��iÂ�W�%�VwL�M�D�m��!��a�B6�k��cO�#�D~ʳZ5������YL���ܗ �	������$.�����SGR�[��6��( ����2U���ƣ.����l�R�|F������E�VT�ӵ���yÂ3�X�����V��g�H�c�5.� 0V�L�9\T�T��3;��KUĺ�[B�BX�򷠂7�>�ăq.�t�*�n�R��>���ω5�������0��ԩ|tJ��X+J�����ns%Iݡ8���!���!�
�ƭ&�e��
�힓u�}p�f%���\eT;Uq����c9QH`�h܈����3���7�|��3�b��qm�Qu����N�P.����ΰ�ʥ����V�����ф{ӌ����)�sv�6�'%�M9W������� h���]1	�A]�,���. É�8A�*M�}qfczo�i�y�)$� t�5���S�|)���@K��$'���盕2�x��`��0W�惓q�oZ��{�3�z�-'�5�8�U�ʎ�� ������V�y�evR�W�>��T��4P0�B�����[B��+G�WS���O{��x�g�D82ø&Ћ�(X����W��u1z*��Rz��g#<`�lhyp0�
z�s����0����sV���~�h� ��䰚U��V�RE�#N��V�HhgU^�<��k��}���"q�J��>�3�S:	?k
Ꝫ"�o�N4��-/K!�X�D��k1h<|;���P���K�� wM�l���)TM#�;8�atyh�mR-O���_S�J��yY��Wa����p��",�=�W�9�&���З��^Z>$�A9��_`#=r�[�;Mէ�F+47���Sױ*�]�P��.��m�Zxpe���+��Wt���YʵG��Ҝ��`Sk�g��g����^�5b��򷁣HR�E��)z����6>���_`��GI����Ab��S����K�P���SSbl�>�L��y�l��c��Tj�B���)�* �^��N�����c�+9\�o�UPz����u*�ųPoM��=}�VCn����SPwY3��Ng#��T���Z�D��V<�Z����k��/�W:��Mh	�趸�z�!�uP���EI�*'��"ܠ�`��a;EX���|�o32���3~�A�w˙ !D�w !����#|\�B�q��E�$8�D[�;}կ>�j`�H67�C�Jc��zVO)GwkmFMVܹ�ZCިB(`�Ƅ�\0h���@�-�͊J�5�[��C��P�,�1b�!�$g��̙��6юH�b�e���R�ev8,[o�קpVnv����˫�:�&�b�����­f �f��f�\㷃:ڨ��>�#.R�@,#�rc�y��;ALnt�mIғ���e��I�N�!�p���/n�)�������x,��Y{O�.�s��f{��K�ୀ�0#k�y8v���ꯑE����ݝ|�Y���>�U2,�J��/�'!���0%��)�����PJ�/]�@��h�{}Ζ*���@9�#q5ڝ��>4O��*������E.�Mw�ަ��3O�c�Y��}����}���뻙���lϱ��ׄ��(��R���;�u�צ��!Z�[uꅮ������zOYh��� ������L���/�A,Ϲ�f��V-�������k��[��j�E�����EzR��
w�������U>I�nw���V_�K�����[Yj���Qb�3v����������8�G�^���)O9��+:��T�`���2L��d��f��/>Q���b�i��w��7��u�\�S�*��f��k���Q�8�F�^R�7���yE����,�[���%8f�!k�ԟ�f���.�A���d0���7LL��jS�S��"��;+��N#�27��2�ނ�w�sP?43��t�Lލe���ތ%Q7éI�b�R�[�l�'lP»��9J� ����n��c�t�b��a�=���vV%0]o����U��}u�;��O3z��#�Aۍ��$����9�z��qn�wM����gk�@..���^�h`�)1B��t�;��t1�BA��d@c�/j_4{�b��w
-�k�� f�EZ;�>�w��ʻ�y�[�2>�r�W�A�$��`x�rVҺ϶Az��d���c!{��ok%�甖H�h]w��9e������]�0T�s0���9��+�֑;7F2
;c�;A��n��{����l����a�/{�Y>J[}:`A
K4�����p�xqT����T��m��yJ������ev̤S�bݝ-d�{�CXm"0Ӕ1e&�m������U>ɐ�i����{w���4����m��J�S:������֫!�15!���V���;�sQ<�|���l�̈́0�jΪ�l"�j��	��k
��weX	��ñD�;�u�GF���hQ7��t�l_5�r��r�$:�%ԛAV�P��(ԗ��q7ks(�o��ٰ��%�v��b��/kYlKNMc�a�6*X��+x�P!Gf��bf&�ե�ԂbLV�κNXai����ΐ�}j>���Ɇ��u�b��±-��M��R<�oB|���4����-�:�ۤ�$�꒻��s��w�(�`���uh>9��N}�6��
{ۚ�5ֲ+c켿��{t�wv�ܚ��duf0��R���k��3j.6"ja�n��o��9Õ.q�D�u�rY�U�ޓ�0ٰ����h!�6���#4;�����;��̵v$y������ֺ�7���	���̃�{P��D_.��m�^�0�cttwHE��K�vB��WZ2QQ0;6�� ��� ���3_M��dw�[N�BZ�*V�E��u���t���C:T:!5G�,Q �DEQX�E�XQUDTV�Tb�""�U��6��(�墊�TUEc��Q��UB�V*,q��H��[j*
֌EAXZ�TTT��UUb���6щl�\Lˉ�����b��)Z(��"�U��EQDQb��Ȫ��h�**1F"
j�14�1
�&�YTXe�QX��(�� ��(�*K-E�(�h�2�e� ���KiQUF*�G)�� �
�mb�X6��"ȰAPE����b�L�]d�U���A`�(�E�AF(���_���t���9�G�� �W<��(���9ܦ�7��'JZ����WvՆJF����&H�&�7Rf�gѕ�\e!��[Ӏ��ڼ�s�%�bcr�m(qE�U�ą`@+�bVwO���-�^5�lg���UR-r!���^�T<�,^Z�ƻ�B~�v뇝n?���R��*���s��{��!�G�����|�X�i�m��\=z���<��V�ZgƤM�N	���Ay�&]:�f�C� ���,hb**X���H<4��(v�m��⪅b(D[�D���lF@�Oitn:hӇ�¼+O�o5��םɅW�m�Jh `!B0ꁸJf.'+*}�6������(�[J
�;=6]����g���-@Q��G�s��r��j���/wp�H�)���)97��uȴeCSōl����0��(H3�����o����2!�P�R\�1u�b/g�8PY�G /�!"Ž,	�˚ʎ���Eh߉��In_:]��I�w�]of�՗Y�L6���=�AV��.�Cf��8u�8�X�vc=���^��WW����'`�v��ق�)@�.J�JC�X�G��k	�D�h�%�jއ�"����c�H<��������{ч��,{"��ʙ��0�|r'zL�z�T�H�(kU��6�L��$���`䮒���]Tk�����RѿEwCN㿮�ꍴ6n�Pܗ�P�ơ�4����
�wEV�+G���3�7�޹@a��=`p�FT������߰��b��w���1��y�_w@����j����� ��{��¸�O���VHt���/��O ]f���Tx�}b�࠯�p����8>���~�=�&�����@<�,���U�WF
��C~��$+Kv����Ir��!#Tp��[��M���X4ڮk��j�
)E��L���D!��P>頮��"`�`[.��DL��XPoe98^�ϕ�Օ¯,�6��Qb4�1u��']��5�ϐ��%�����]���~�>�/��Na2aj�t���$[Q��'}�ZĖ�w����B��tgoVvm�E�9I&�mF�]qU{9�zSZM*�έ�(�6F�x�Uy!�������J^v_^�mȰ8��g��o�o����C�EW0��&Ukmv�5��:!��dh��� ��vSP1U� 7E]�~�������`�4}��9\j�yh�f�jx3�Yy�:�j���������}�+��r�N
~�AYd��b�]a��6<צh��uE�]���q�l ������]�~^�Nj���c)�GM"yx�R��z�f�Q1ǪDf��-��B�`�V�H��]	ݧ���2�PT�X���.%���kg�:Ր�\�ݷ���YJ�W�lx�_� 0�<~�tj�a�^�﵈��;���:��2ܥ�+�u�Bm���
�S	M��ED����"�~�NЫ�(���z�Q��=�YCQ�͵N�c�˺���5�����P�#��9|1�=^���Y�mdVoZ��ƆAr����3n��.�--���b޼nٶ��k�i,Ŝ���nm��O"���v52����mfF7Ne !���6 B�����۴y����fD�l�qn��'DM�����[��xwH���\�#�'�����X���Y����W�?�W�!x�43Ɛ�fP�E� ;���]��ʀ�N�nF�N�B�D���l�l�g&b�l:V����
1���};S�_	�~�p�C���x����)(���9�W��N�Ԍ-��"9�v��0*6�T;u|�0��kxη|�P����0⪈�23Mr>A�KUp�J)�so:���=��=K�aT�
�+�<� �	uD�&��F��y5�$֬�^R7��| �Xb��3O�^�Y�^j�a�üP�$�E�{s�W��RHK���Y7錘��Yw#:j/��O�M�IV�=ç��̦�N��@��V�\<�n���`��әQ�D��Sep}� -C��WP�C�"�ui���[�B
N4"���U��lcT�cNW;����K�;����l�fU����F���M��華1��,:����Ǭ�xUb^�<�+$�˝��UG	�+JO�����#ЁzC5ڗ�xS��/�V:Q�X�[���ɿX.��N]�!�W���A��<�ҩ�����;h]J *x����2�zPy������
�BԼ�c��1�31�I���z�׵���W�d�7�Ys����tB��:�)�W����wL6�ǵ�G@`�t�fB�׈���5�ze����Ͳ)�1ЧG<�B-UH�=.؞�t�W����Ǻ ouB����>=q�3�휮s��^^FK<��'Ȥ�Dk���Bz�
�֏���#���b���G�������j��m�ɩ���]^���H0 F�<)#�a�xyW"���~�;w�G�Ί��V�壚U��.�8 ��������\�8re��o�*������@M���*�]�<�*!�1�E���
�j5�BM�X��{W��{1Tv�$]W[V��PEΖs%���u���
��x�{n�;��B�X�)9V2뇩����}��xR�Mr�$5�\L\"*NT�w.��ɮ�)��[���A�e��+��l];!��!����r�+
�ǚ����VF�b?uBr���.���Ɗ5VxR�|F�[d�Z�6�{���<�)�(�h�8�(U��p��:� ܫj��!1s`V�'\5ٕcG��^n:~�XK�u�+�%�t�躚Ά;gƥ��z��>J��)9���P��\*����+��+�f.gT��%g�8lͻ\�Q�l;�".:}7('9���:7��`��1� F"��Ի��q���;��#b�3�\J��T0Eƚb.6X�TC14B�ѹ�&T�9�i������p#����k��[�=�t���uSW�zb�S�z�mL�ZK��W�  �	`����	��-�O)Dt���³O�'d��b��E�>�6<<ܣ׼=1�KB����kO-��q��>�|x?���*S2(y]r�;��.�33�b��^��X+c���\�uT1ěd��7C<"��Avf��gti>���O�O+���0&���]1j��纐}8����V��e���ޱ5���-��/�5�y�MT*úY�F������ I<���L���Ё:PVM�P�9LQ;P��	G�����3B��¼>VG�u�G4���0���Դ�s�gy����ꚻu���iT0v�R�DU��p��v�QE䨊� ؔ48��.�ϐ���%CF.z*�eк��j�L��yBݸ.ꢼgD1�&A F��ǡ�^��P�:4�VeFϳ{���âũ���M������#:B�#gj�971#�6,��E�/�fO�˻8)���a��N�=zp^����dm^�in��v�B���+8[�����M[@�x��!��}�V��W��gN+1�wVB�*�����Y�#�";u�Y�7��ŕk"eS}���5����c#�]+�1v:�n�Fv������q�3u=[���<	�&ƤsR��vs�P��J���������{!D�B�]OIl���9]���5��XӾd֕�gc�}�
U1�ǒ��O���;M��d����}�-���oG+<�j���VYƓ}
P�IW����P�W����nU#�S
ꝵ^����u��@�j�O���U*�)jh�魨���7�%8O�Yf�A�17���K/����3�Չ��ӡʎ�^����´Lڻr�޽��g�[��<e]�֧�+6��DtR��#Z�D�� �^S�YM�`�=|�|��7Q�n�x��\Rw�R�^�pnX��9��� ���'���}�����8Iqč���͗��h�L���Q��d,��K��"�^�jv���̤&�+Y0V�Yܼ*8���V��OT��$�.�;:Z�cH�vwQ��G"�����O���_ЯhcuF���Tu�����~'�cVa/説Vb��H��<�ꁰ����H�ze��9��eU�QҧLK����I/q�uf�C[�sw��ޫ=Fp��皻��.�(��r6�J�W�,,�i0k�Y����)^o5w:d;�4�6� ��V�'z�fV�",�5��3s�7<hl$T��Msrvq�����Zfsz�q���PQ�� 3k0�Kx�e�\n�pY7�W�<�s�4A�_��2N���\ɧ
3"c5u�vk8�[�gI3#����\O{����c'�HO�����n��[�U��
����9�3]am�֗(�{����k{�|�-310A����C��F��gƈ����n�9]��C���-���ȸ��4�X��S(*����wm����9Nc<�r^	~��m�����3ɕ�����%���Ӭw��@���ϥ^b'@��>ʣ=����^����͊HV��O �D��^=02�ֹ�S��6-����P�u�n$�˨�X��Z���w�"qɈ��q]�x�n��s�z)�C���u�������U-)ڱ2���ˬÈ�IF:ثS�f�2�������Q�P�;�ss+vaciS���(��ux��0�L����_W��3c�#N�v�u��q��I���{�zb�ٝW�x�w�r���n�d�r����X������Eũ�~Vz�q����6J��7�C�nSq���jS��Hz�0��=�R���F�/���i���bC&
a��ifC��\���;y��v��y�#�.%���X����r#Y�b��VHV�N������;S^��u(���_�mN�,�#�_1> �=�U]n=7��a҄��s-��tZ2���r^�ʄV��MKq�]8����Aumuvn˵��8�ܾ�#;�ȗ��{A���-wM�]���<\�y����ɬ�:R�Pe����(n�Kn��X毭���e��$p2�&m���$�U�۫����N�s�������:�����:)���<k��P�B�mcu�sU�t[%��+0T��t,�S`��qe��ux��.#��`ǆeҕզ��>ޏr��{�r�`�=W��}�6���:�S�� *�Uwu�b�;x���wd4i�[�)�K>�~¾c�%cQ��f<��p/��I���\�73�+�7��O΢g�&�5����� n7;8$�����6Η[�*}��bQi���E����5��/i���M.�J+T���Lg��糧p��(�`4���P��/��8�"����e��֭�e��"�zn��G��Z8I���Kf��aY�#�2�]V��ɳF`�uo��z�N�t�7O���M�������VT�ʖ�Fi��X��+x����e���-�ɴ�}�:��YՒ��]�7���:���A,G���G6��M1�+$�Z�'�)^�U�0���E��]�=��E���1޸R.h*�G݊�Ɓ�`���;Uƛ�ō,RM��'#Y��2���֩O��T�߬�#���x���b#t���t�W�/T�iօ�/'Q��͛0����k�4-y;([����m�]�N��ԕ��s炒}��V����'H��&⼦�<��JQ�ݼDv�4*en�-tt�E�<� k'<��vޛ+�����0z��Y��&�k�i=RQں���r�(�
Ƶ���]�_���<��{]�P�t���q\u���-B�o����Xvd���1�Z�9*C�-�W�8̹R�������MG�����[�^����ôD��UQJ���#{lQFҩ�Qb�I�V#E�򅬪��J�r�((��U��
��t�T1�4�X���R�D����X,U�eDA�h���V�""��ETݖ
�5�ر]Z�X�`�1A#���
�,U�R�ň�1�,V8�b��H��EL�VTQdEE��1U��Db��� ����0Ɗuab�1X0P`��V��PXň��bAQU���PTQ��h�B���b�
�"��UX�H���$�A����}�����p����r�w�D&' ٲ��<�{)�CXR�4$�M��%�o=��<wJ���/(b��>���.�fw�Z��z���yڵ7O*]nԾ��W-�8^c�~EѦ�o^��{�ۙ�7C�F�j�p�y��|�L��U�K;Y/h�V>(A�M����O3Q�K��L5�2]]�E�F�$���@MX<���KW	a��-Νo�-��/���h@���fñg�9�x�q�[Le��/��AG%Ī��QDt����e����ᙅj�pG�H���FPbʱ�>�-<���j�}=���ڌ��L�M���Bȋ�K�F��Ea���YWz���}8�3�u���>�x'�"�Y>`��۔5�	�$�HT8��љ�n��:=�mv�Y�����e:x���U�������� T��š�CڳՆJ�+Z��r�sS��ڲ��C �v`��E.(QQ˹.��Q�)�㺆�q�5�:M*��}��Xt����个�Vb�)$I$e�1�����^2*C0D_����f����'Hy�>�a����/w���9�T��r��o���Su�11�+���X�c*�{,�l������*1�:�3�GL�+|^�u�~m�n^5�>�nޏ�vf���t��1�[�y^�M��O���U���
&�-���&�]v[!s�'�Ź9��cY�M��%�7�y����17s��l-����ڢ���u�j�@�j�Q�זY��ć�Cy`����M�i�Ԧ,ЯA�2Q�;N�T�����%9x�>��h��\�R�9��(�HϚ���ma����ʺx�e?���&��|	Y*m�mie[]�����Y�+�y��F��d\0�`���l�7�]�Φ�I��u.q��c��I�اoִ��G�9{hJ�+l꼂/�&�p��$�J�k��c���]��jy�sWu6�'Yd�	n��]��e�z)��Z�GdXu^��Sy���e{�٠��Xe��Q�p�gD'f�;xsRH*�$�&���,�.�e���u�)OʤWk���z�svI��A�Ga�}��Z���ζx��vV�_�t��S���Tߩ��Tr�*a��5��W��.x8���ʁ�d�Fc�����"�%���<���Yqh�==hV/*2�L�<u�^鲈�Q1Fg;��n��޾Ĺ�e�L���Yk]�:�p}���ꉄ�i��c̣�^��um�w�)ѭg/�uF�x�G9	W�w3'�'�݀�(�	7h֘��;��Z�����]wL³��?frr�nלp��F3�,ᱤL��\�'c�"�E�.q;��a���d���<٨�u1��;����P벢�׉f��N���Ҧ�#I-���8W_)L��@�j�QsY[��ms���ޙ2r5EL��>%��\^����>�H��F�f��z�o2"��Ok|y��ut	��:E#���Zg���	�Z�no���t&�e��}*��7�[�*���M��dЧ��0՛v�����R��,��{��!{8=�>�r�e�}��ʡ0��!
��<����t�̺ʻ~����'7|����T�d�t%EK����!o3�+�7}<@�=���j����ݎ���T��ʽ��a�~v�A��3�rGoۓ��XR��/�Q!�a�Ki]t�(��><(ˡҶ�_o��W7���t�?���;��f�gTs] ;�3��æ_�{ ��*�Κ��{F�" ]$MI��}Y����j�{[�3���T�k�a肣�ߥ����ȭq�KHf�Q��NQё]p�u���o�~����C���RІ֍QZ0��H�g�by�q&$c��Tfe���x��������-}7�q��Y��!�y�wH�/h/h�[$�~r{{�h�ʑ�8����d޿�ީ�W��|�9�םp���v�U�{����-q��mLg�7�r=���9�/!�dO`���u��Q����I�42GD�լ�f5�}0;1�(��~����V�$�`F�oy5R\Ω'3��v>L)9o�]=�u��>���B��-L�,��>��P��S�4f
�>݁](�-���*�W��c�j3:2��#;"��G��+a^��fR�C�3f��8���,o_"H���i&� ;���Ǘ%v�MC:+q���r�]���M{	�zb��%
R7k�C�M��Ox����4��j9�+Tk^M�5�tU(��-��ֲ�$�����V����S�靉�$��q�����?VH�TT�DY���&��/��ؠ�G���6�7
a��_y�6?�5�;�i�������,Ҕ*�q�S��f+��.	#-΄��=}��0���Wd�_�o��D�U"ml�KP�5�6�˺�%�L�ƖP/��Q9U�k�J�7RWCy`�%a��/����H�2C���.��>�L��N.OḲ7p3��f+h��9~�H�V+Ѓ�}��m�~�c.��㒐s/�����	�5�{�zzj������!��������v���q�t�C3y��O�4o���9�.g�4�b;����gD릛81j<80��r�[�a���Հ&m��L
��۸�]�{�~ax��.�U�����+�,C��e�oq,,�qkQg��ǉ&��P��� ���[ǼP�W"�+����y��q�|ڶ�$5�jg��SD��[��dL&+�u�v�O��6h:��\�=��U3c8�w\��^ܗ^�c9�w��fa%�Һ��kܻ��Wn�y�{>�b���wo��/�S�����E���q[�7����-��o;��p��"�G�2���aޕ���#����m@��@���U��Lx,���[��K��fa�G���չ��������J��5/�oޤxu�V�`�N���)9z9��[���/�z,BH����wt��p���/C�YC㳹i�`Rb�t��\8�]�K7s��<�r�Wp3ru[h��_H�EC@v�u���g]�RqV�vM�ha�̊'5�z(ee[��m�^�yyUv���J*#���z��O�,Y�w�9ؽ�q��r�1U�'y�)�Oz6iauXWC]�u�a�qꇯ�,��FQ���x�7��Nh�=5Q���;�\_�'�	K�ę��r�>2���zbe;K.���Ҏ4�y_>����[5�թކ���]k�w�=xS��P�t��S���'��r�������'7u'Y=,oW����xz��=���Ʒ�*TᖳN���Z�aC87z..���(g<};��f�m9}��\w��vUZH��Ov�kL���N�N�_�-�Vش燍�ڝ�j���\�x}So=����a�C+ϩ����U���n���嫹f��lN�!\�舵�nM��oo�I0* ø5g�܎@���|�ɋ$tj�Oe9mm��nR���q��׀Wt7�&H�o
I�PN��]�ѱ��&73\�k����VǬ�{���\��+N�8�s��.!��K���jD�u���d��T�ɮ������rȜ\�Ґ�B�N%�iȗyqY���1�	fؽCo"�e6�P�c�8=��{��'������1�MuJ�J��wn�T��l5��Փ�t^�Ou:y�m���m��N'�H��a�g�����s4����TWۋ��؆�ye%'uT3<� ��xm-R�TB{��ݜ�S���N�IŤ���؉�gz=,��& ���ݲ)�{5<�3�/=/��WUAZ�W`c���f��X~�8��ϡ�0�&��ܷ���a�p�X8y�m2�V\�,U�V=����ڼA�-��7�tbt���vL��`��v��އ���
=�<qU��A��"q�ƑNŃ��}��m����oQ��"���3	��ۈ�z����)�@�V���Iat������{ܷ�Ʃ�n�@���/���}�>��0�^~.0�#T	�Y�����,�z�g�r�e��yn�sk��J�K	J��J1g�ڹ����fp]����5�*��0��`��d�SwI՘�L��q]�X��`uv 1|�P��q�ZN�f�(��VGGr�es��)����"l��"/RER�2]�S�)�v�����'�	����_�ǢQ��o�]80�Ғe�Z�$�U�_��8�`\����q8����DDD�RE"r�����2nEE/`�"����&s$�)��;#��h�]�=l�'���$	!!�а�$����3ߩ&�R�wC����$E:�H�#%ՖX�aO;��zgg~7�XX"6Tji2�+�S�6eh�WT-�,���(\�,qY��+�AQO�q�x݆�� 	WR*)�7 "��ҌBIfs��	�A�>Kb��?�s��a���X�������2���D��q!f����;"Ϧ\hرh��Vp��I��<��6���}�Q�7M��%���w�EE"�E��r�C����EQP6B� n=*��d�����~��a��P�yP�t"����J����rfvh4��=h�%������	q�b�w�wrY������/���a�D^9^�¿x��^��"�rD�F@I�<vn�6����!�v�C���.�6������PTS(l���X�>]��R�[fG$���� 
��cc��;�H��,��d�&4��%�����$)��{��&���U��q1�f̈�%��1
���Ê	%��Vn``��vv1�k .�k#�!���؊R���PT��s�7p�]	��q̇�
FWvU�	�{pOm������D�3�͝��c���m]W�;��)�C�̓�сh{�EAAQMF�r��v
o� ������G"i(t�Q�0׉Ю���jLC|�*@�2��BdIƉl�ԻM��W�C�៫��E[n
f#�AQMC�rѷXS<�����d]�ҝ�X.�a�Ɛ��@PY`X����Q_�E�0����30.��=YJ�ב�:��`�W-4qYDd�\aD��U��a� ��I[��vR��.�p� L�O�