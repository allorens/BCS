BZh91AY&SY���;�_�py����������  `���}�Cc}SFڢՆ֪��Y�6KZ���Z��*��     � P(     w� h *�T{�4(P 3�'�P))vwȥRE;���vT����leN��w�kh�x��m�
6�5�$ۉ�wp7n�ڈd� /�x*%;h�Pۅʮ�V�l��w`qʽ��q�^��m��Q]�J�q1R4�$� ��� 46/+Z%馁p�"R'n+��Rt� �E�m���Qp�u�J���G� )LؽPz���\�v�u�����KzR�C��^��\��������ΥN�a�x  z1�w��-�,���J����+G����2�Y*��H����u�����     P    ���kf  �?I��*�J0M0LM0&& !�#L�S�BR��� 4� d  �B	��	�
z10���i2I����@��L�J��MM��2`2$@%J���	��ha0�Q$�TBh�z�14` SLFk����jn��4��R������+͘  ����*
  ��
o@�*��s�)_��+(>$�C	X�Rx�$�MS���V��2�?�t �ڑ��'��Ql�I$��)U �!�>>�$�z|=}_�����!�.�龓�<w�3�It��ȐPZ
�DK�P/��=�-c�i�u[}�J|֚�)���0*���u�g��}H>�Xl5�ȗ����=(%x��,��������Ij>�/q�����*���V9��'�e�w}��{�q���M��`�cO@v��ѷ��ɦrV���C��m�#5!Y��.o��wD�.�_D��7g���hZ�֝
�&�t����^��f6�m
Ɵ=�/l�g��#<�~��Vo��f��i=f��9s��D�{��s��׽ޗ�����ËjCq]�uw����a��<�g)7KØd�)|��=�W�F�+���C�ο2|��}�}�N{�v�X��;	6
�g�}����!W��%�|�c�<�T��*Y��X�����Vi��~�Ǖ���r�k�Xfa^þ�x��'��ϼ������?<h���AZ��8ͤ���ga^��⏃��,52�����ާzμYk�gѾFr9��q:�f��K�UVeQ�����K��;�LD��J\jԱ��̯�$�D���7��S�؛GY��'��]��n�Ø{�W����I� �������c����O;6��.�&��:��@������v�ou��]zu�0��n�w��ln۷��F�Zh�gƮK��y�^zR,�����;��<��~S�މ�M�u^���u���u��[��$#۩_j[�K��{������ܝ�f^���I�������mkms\l�GY����x����E=�u�zS�K��ʢ�ڱ�r�*��u�aU]*��:-����Q�:����qݛn��6u�μ�c{��B�2�/d���s��{�������f84qqv�7֧We��/��'o�����6�-J/�^�������6�L�U#ɿw�������*�z�O,H	�$ve2�a��^á��E`��Q�*�ҫv���cf&�ec��7�z����z�Fx�A�.-qJ��W���Co�l���UQ�u�fS��8:A���w�m*��O�[L��^(,��6��c&ٷ���ާz�յ���ETg�^��>�#�$�|��/\*a�<)���>'ŪR����-�����k����v��`��]�z:���u޽׺�k�_��m�664�U����k1�m�ڤ6��7��S�؛GZ<��|�֏4u޷��uٮ��:�i��7m�~o��5�hӤu�6<�U*�z��]W�=N��}ןu�����~S��D�7�u^�~⽦����sn�i�$��.��'�K�K[K͔�^
G���<����mu�����[uN�����0��]�W����sȯS��w�O�e�6TUҝz�UWJ��N�O�U*��ֶko1ݛn�}�m����w���)j[f�2��c8<����}��x�!�XT�1���xOy,�+�9)�Fh�M�w�h�ܝ�er����'��Rϸ��aU|�T�M��J��N��j�h�X�x�X�|gψ�U:��Ӳl��.Bu��v�xΙ�ɣ�~9���~99h������~;�{�t�UO5��^�(u���5�uK-�S�{Rs
�įa^�+�[�ʫJt ګ��F4�mڻ��]:�fI�jN����sL���;]F�^	Ոo�����`����Ҫ�S�xڠ�X�ڣ��`���ٟ>"�������q*�R��uЬ*�ï.���GX�m>��xi�6��i�m�3j��uh�U:�CB�]����U�
ͪ�]���w�1o��Jt/U}��I�)��$��R����E�x-({�k�v�[�TeVҳ]Q�u��K=Jᛉg���%7��ExmI]ES��:kN�I٦W;Gh��~�p�F�pP�R��z&��1����^6�5�!^�����/��W��}hj��>��P�Ué�t�h�u�գ���{����y��{�M�WUo���h� Ѿd�0k����&)�C]8�k�t�,>�iK3��S~��`�����b���b��V�>�qW4�pl�v_pk�u�������b���y��}旼���~:�<7~�Q��3[�#i�O5/\*.K��}��<<G}�!aTG�1ЬڬF����B�޽:�Xz�O7����E`���A�R�}��18Y՝W����vC_��]*��:6��ڮu��uV����Sgg�vu��S���d'Y	�I}�XUg�^]�Uގ�z�}��y��~�=��:Nv0����p�m~�5k�q?�HĲ��HZ���������Ҵ�qkv�ş>�3���Tk|�S��D/;���k->*8��}�l��;���I�������<Gq���.�1s�bx	��WII�z>z0���Ѱu����[�3��U�.jB�&-����z,{����Q��s搶���q�MD*�Bkާ��ur���-3*'���R�s\������)��+;��et� �!rgw�,YI2�@`}q�A��h~���}7�����D���	#7<^Qӭ�IG}�Wf��8M��{('L�B���hG�=��R��sC�b	��4�D�=	�xv�	BU�j�3��YrcG��ऱ�s��7���H�)�eNx�;՚H��f��m�ZC!m�CPн۞�>�3���N��^
�9��>y쯝�FΑ�w��~`��|s����	�W<���!��i�i�:�ҟf�������L2��-�b-�G���V�������5{�ƕ�B'7:�g�k����}��>�ddj!���|�!=���/�&.��+)�6�3f)���e8wE��v�ǧ��Y������NL���H����{����>=�<&Y�=.qK��G���������$�$yk֍�mz��#�qv�s�E�27�g��$��������V�0�Z֊��wV;W-������S5�K��7�;�Jř]BxQå�S�s�,�xS�-Q�nl��Ybt���]����uf|������=k���+	|�C�I0��Y�<G������.�n�n,3pY�oJA%�"�K�~�hZ�+�����|T0��� <����r)0�w.q�����M�[0�	�L��<��gZ�t��~>'8b�'J$��K���<���Jn�;I?�}�]�[z ���i��{� ����hf��^%��j�Y���gk3sq�h�e��yEGM���8X\w	����i���3<�w=��:5��/7n�vf\צR�2eC�=[�j�a'�qVܵ���/�p�H����ƚ"���֖4��N�L���x��^OG�������s3߻y-/(g�\��.[���"���8����Ǹ���;�<q.~�L���͊J���ޒ��w3YU�y�6�qY�B�pb��{�*�Nf,�e�.?ovg/CsUK�&���b6�;������6�C������{����{ǈ;Ϊk���=���=���mX�ی�#�?�5�[Z0ˆJo����@�F#���pY���}[�5z���&����+��~���yV�n��e�&/W	�K~��l�⟨ٯ��7�_����)s<\]q��:�,�ޒx��_�6J�9�2r�	ӥU�$(H��FfS�>1������x������=��>�����������W�8�6v�>7#~���`Ȱ���k�0�Y���b���j0�,���V�2�9|�n�v�s��ػ��\��i6���5c�t�nj<U~/������ggmN��g����3t��_qM��o�y�'5�D��&6�W�m$���d���	������+~���6S1ڷ�љ!�2E�n����+�A~U�2��O����q�KNO�ě(�'������o�y��PD#{�fY��{j����������^)	�{��|��~G}U�d�'W{g�r�����>��c���wcOؘ�Oc��>vn���QzIA�����F�7KGݜD�c&|�'W�Á��)׶�Y��Z���{0��
n��w���q��̸�!"�bѹ*7ƅ����=��uȹ�^CI̫:ۚVO���̞zaZz����)�L�0��i�p����y�s,9��GE�62���f%�=w9��1�QӐ��\ݽh�#���ϴ�'3�fG��]S��M?���D�=�[�9�������˗��G:}_��a$������.?�+�L�ۿl̆E�<V�'=����<ףK$����J��iiܺj����=���Ş�����9���
���X�e��!�C����.iKa4��昨���POF����l�`�p���R�n�ӫ܋Sr��^�	����Z?aZU�S�g�׹FO���h���3�Hip�}Nz<�;�g�ә�7sa�4F.8��^��&�r<q�f\�va����Ƽ��o+P���W��^���v~逴��:ٿ�o˯^�x�Y��=E:t�f2t�����f�>�+E��9N���^���Ɏ��;�î��=��GOKVC4X�osϓ��G$-�Ǎ���?c�N���y���b�|zs�ׯ�'��<�5���e�A�Z6��qÜr�Tj4T	����)H�U}st-�4�Y�h:Gl���V��,����o�Ii�K��Q��v����v�����RZO�&��Yw�]�a�ק��Q	�L��ժ��(o���C�����y���U��̣E�S�_6�k���2	��o�gX5P[\�ꃩ�Z�P�����W*��l�J?�ܭ>���J�W��"i'#�hH�캊�Ld�\l]A����������w3�u�_��1Jwg]�3^J���?:��Pn�)i�ƿ/�uho.4^����`)�ߑ�7o��?��5	��L_���m�F7�ʮ]�Mk9�0�w��̿�k;���C�������KX�瞺g��Ho0K�cZ�׷I
�	�eJ�19M8ֆ���[V��Z�B�P���%F~,����H�)3Z�2�m������$�
:�-�����ɪ��?B�u�PTZ�5�A$�$�8��Zx��$���n2IP?�P-*N�>a���a$�Y�>?:"!��O����Y,@�O`xb�"��Ɉ�*0��TL����v@Ԋ2�s��������A^��D��P����28�s6�N��$!��"���~O�P���V� H�@���B,�D+��)�$\��a��fZ=!���l�0qr-��w�Z���Yuy�˦j���c鹦f���f��2IIq�1�YL�bJve��iٛz2G������3���V�i q(H�0�/�_}���3�i�6(�Z��m��Ib?�Q�!z>Y�I�d���g1�jd�?���X�C�1�V�ss. ��Ț$I��
M�3nq�����u�?�''�%$���p��Y�}�����XcKi��
Ϳ2"��2M��{8�1&�l)�C��Ǣ��'���
�	-�K�=Y��#cY)��d��8E-��#��_��11|�~�����aˤ�n��!��n������6&_�,J�8�	��$��x��5�4}�͚�50eЊ�Hg�nQ�B�ϰ.Y�} ��Z���2� �$ѕ� AW��2aq���(Ē�"���J.}!D]�A���z�Y��e%	m���\H0$A�/vMEb?>����PBp�w��A���I25��)�/D�蛢�7V;,�F	�c(A}#8G���E��2IG>r�5�Z/,�M���v�E�jO��؃K��	�0`�n`�������7#��l�0�gU�������3�	�]�݇�����0 ���O���H���#��;	'�D�Kôs���CS�~�C&�D�ƶ�����+� �� � � h A� x@ �p� t@    � �p �� @  B�=�_��z�w���{���AIE�;��8�@ � @� `�p 4��  � 4 �    <0 4@ t� 0��  ���{������{b�\A $D���Y��= �  �@ h  ��� �2�� �( �   Р � �p
 � o�^����8����"�D�J�H�����y�3�( ���  B� �8 `���p � 8  �`  � 0� �@  {����� x` ��%�S�䖴�� ��s6�`@ t@ � 
 @� `�`
 @�` p 4
 � @��    `�o���x  `r��}�mr��� `�p 4
 �   �[ @�6 x` 
 @� `�p 4@ 
P  
����{� � ӟ$���|�,� �fn*��$!!����~�~A��S@�qS�p
��ASa�f�V�6鍶�޼m��=v�Elٳf�W�������m��6���m�lm�o^6Ҷl��!qR�b���˨B�.-Z�b��˨B������/.�X��M���nճf��Ɲ����m�i��b�lٳm��j�m�����* �s޳${�ٜ6?g�-L�����
4;4�R�,�֬�˳.�p����7� �22���p�+�lH�,d�&��\�c8
�2�*�D�(6}`_�:������Q�IƠb�{Ye~<ߔ��/�v�d��!ϊDA@�'��!t�)��Xe��)�!q�ʬA����uy�-�&��
f��ղ�D_jc��r�N�I��a�P\T��m��c�j��S�Y���AD���[)l׾��L��2���Yp�WX%˳,pL���]��I�	�d�&*�
�O�X��*h���E�6�!�5f���`�r7p,�ֵ5u�ls��a4�l��J@��Co��Fgч�:O�|<�
�d.�Qh �* �8�.I4�eI�|+�g���N�į�/�I'#�L����7Q/��}��&]��������r9$˻��#uI/���&]���H�9��|�$̻��$���10��c���9n3-�+߭�߈m��hc��Zj�jB�iF�B�#(��s����	��e��e̺548h�����4�(��	XO��&'���ǎ���	��?�NϢqN�qVI�/��kG�Ys�%I�=F�������QԚ�7�f��Z���[
Β���CdЈ�!�
+˓ٖe��cnCI�4��:�!uEJ��+TesI��n�4k�������=����Z��xXa;L��2q��o�\I�d+Tu2M�Đ�@�|"&��B��~�ѭar�\I&�pN^�J��*ӎNt#H_4h8]!��.Ead	l��N1�cL$N��p
��)i�-�x\�-�WL]W!wS���	�O��I'��Xï}I��5��tDL4YC�ı��8��j��ݛ�&�(j̹HçO�fŧE_Q���o&e�]�n�&%�f�4��9~M�/G�.�#WD��*�}�5P��2����lA�% aZ�W�S+�n�Q�(�����F�ɣ�c�Ut�0 �v����?֖�=��X!�Q���3�A�f�]v����6��A��Z�e��miU�J���0���v�������hO�q�b�@�"�F[&'"2N]&Si��M#0��9%U�`t�+Y���/K�6r��M�2��kF����NU�2!��ؗ��I�N(|���G�UUj�K]��h����/�0Lv�ӛri:��u=N˓Üa�8��[i�c~k%��,�R��ж�d�,�H�M����
hێ�.9��I!�GRRq�;nӣ0��H�{�G,�!
'���K��ܬ�3-��rIY1`ˣTe]Dh��C���BWK�.����F`&�E)E��־(��� B�D��BY�M����̲X�1�q��y/�N&�a�u˔���	_�Z>�%Z:b�eA �������I��wI� Ng��.�Q �B�.M�m6���0��d�hz�qM�a�4W�4�M4�{�����O&�$4��4��B}ྀ��G���cq"*8�"	$�E8�N��I�&��SN:�n��xJ���E��o!�i���l� ��Ӟ'\^�AMI��ΖYe�ckX�X�E
�7+�F���]�2�^B	��du5f1!��U�~b$�%MT��[1���֯NF�Q�m�8�������B	˖����3�Y���U�ڐeˣ@jV4������Tf���r��۔�p�.S�E�6��$���ه5�r��9�S�#�@�>I~\��(�D���E;�t:�u++�%-D��PV[X����,��>��%��ˆdI�����P��D<+H���}Jh�v��3�Q\D��ciהs�!=N�H���޸S���ʭU��/.��"\s*EQW^��;]5�Q��]6�Ƀ.܉��{�o��A!3$DЉب�|5�
?�
5�k��4Bxi<A���\^׎���q\^׋�⸺_��p%A��#���Q�5�H'���	�#����Ê���W��q~W����>WƉP|(�����x`��|;]���xxx�9��,<=&}$�4M���x�:'�Y����O�x'��'�6?���pOH>���'�qg�I!��l}����d��|(���|C��|04x�ߨ��}���w~ם2Gy�PÝ��淿�x����3h3���=J�և�\��oG��{ù��> ��2���Oex�,����S]�A��8n�2����x�� ��G=���\ĩ�=��>�}/&dR�G����� �����g;/�k�\ӗ�o���hD�9����D���ϻ�k3<{�����$�&e��=)�4�����w��S��$̻��)�rrrI�wqBS�������fx�}��yab%կ�<x��,�z��(��(�YT���ȝY�"j���F��=��1)L��t$WI8����$x�0�J���1��b�8�	�6�%�@�0����p�|;K$LbE:��$��M�)"�H�����<"�b< �O�׍&���5DYdՏ������x�<���)�v�����M�,��,����?i����Z�jգ��f�Q���&�1�r��n��W�FG4QR�S��$�~�Q�����":<�{Nm)3l��(/u6�&)5 �ZP.c+��wM&�$�����t�H�ܧA� 2��,O�=��=�ڵ������'
J���b=�P���fB��!���$�1�V�o$���mt	��e�Yf�h� ���:�K�?Al�]gX��
Q�'Q�K�j(���� �F�hHP��T�&>��&D�	%�Y2��	H\S6���EQ@�sQ��ӗ$`��,-rH��]���]Rj|D�%:H��RD����=��jQ=�n(��{$!
mȌL�%>xR����G&p���J��Q`kt��H����$t�PH��ar$��D8u)���5��wrOd��;��F��Qc�<�D���F����rv�2��[rb�0b�����{N� �pYƿj2,{E�a���(��!��e�Yu��5.jlQE$W)��)���wt��Dť��)[���O"e ț~!I�&(z�4�F�b1#��*�qӴ�� ����4�Kcq)��.,s ���T����km���q{�sN���,̌�Ը��H��'b��fQ��#��r�5��Č�L!�m-���R�$F&����<�
����X�))��a�+L|C���,��Q֍'�I?fW�
0����6�"|r��|S� a�!J�'cYJD��C_4�9�9�DPI�Z��Zd���me2Qt%K�G�����˻w�ue�����Ӊ$y�IJlbm��M¥<��Yeݥ�fu�j:�o��
�`���=�J����b[$l�K�����P�}$�����<�$����#,�Ѵ�k��`>4B��!d4���,��Ҳ�����"aj�1m	cM��)	���Ma�$$$i[�,�$�1-�P4;�NI|y]���7�:W{Xdˬ���-W9C\��T7FQ������w�}�4-
r���U�G�6�`eS���a����|G[n݉ ��!V�뵞}��ױ�x㑣����LR�p!��e�Yf���w��$��&�0�!�U|Hi��7�l�^�>��p��5d%�Be
���`��@�!L1mZ(�㈈��(��SR$ՎK�r�e�!q���ܗ$������(�;�!�;���{�Ip�ݧ�>F��d��l�u�	Ԫ�i:�&��@d�����>�"�t�d>3�����_��>�e�s {��&Nf�h��XH@�hP�I%?|0x ;��7J�y�l��:�;��4xڰY�l�e�Ye�!�'�a�Յ}'1:Rq.m3���y��uz�b��̧-�|86�m7Ú7�a�6��p���9`mئZ�}�)�!%=��WiO"L�`k��K�m�/N]�Lu:�*�;5
t�1$!$<�ZI)�K��~>�4�z=RnI=�Ϟ�
�Lc�Oͱ�'��d˴Ly���HX�W@�wѷI��>�L���|����2�� �S��V��.��)@���dK�L��w`ZG��z����l27��0�F^$��&S Q'pz�Q*J4�'Sŧ �D��;��N:�%���&�ƣ�V���ƛ~!Y��Mđ1���#�^^6�����Q�x�u�����қLr�Z��AӀf�_���4M�l��f�(�7N����$-;�Z̀p;ȝ�w\9 Cn�%�����I8���1w��Re�o㤐��f��U8�ݫu�>>�|Tx��;W\-98qQ���V��uQu�����~�����6a���Q��v(��#��D`���L�qU_��W�X���1�W1⸽����q\W3�����M�!��p|(�Q����DE����į�O�����{_���qj�\m�+g��8O!��M
>|!�0�0�4z<�����<}���xN������6;��!���<a:>xgG����ɳ���C����^,�|~~��N�����2p�6?�3�YH>���|C��|>,�45�zq=�t�n�*o{�c茻��ˉ	���|W4>�f=����C�ӷ}�=�E��۝���	�\Hc��Ɍ����J	j2��ʊ�S"��D�f�xV�tIJ�j��
W*ͯ)L������Z+Z0$.0����(_0��9ﮜӅ�����g������S�F(�5l�����X��{M%�,����z�L:LvMT46@e�L-$}��d����C�F��.#��$��)�Idj4�H��PhD�p�ٍ�$��,"���2qz�me�/((�l�`P���y��i)�:�Y�A��e5
���������4c4I.%# ���a�Qt�t���K���|�0��Zf�2Yi�؍$�C��Y�� �29!E�]�X�(�@�~0F�`�,�w�0�5��%ᡡˍ�c��W���D�˗�ż�^���E�N�䓒wws"��C�NI��̊�9$���Ȥ�T9$���Ȥ�T9$���Ȥ�T|�\qXV�c4�ck�>��9�܁�D�A��_�2��!,c��*�Il-nРr$�Q�+A�r��¤0��8i��>$0&aT%A�D��ˍ����4�H˲�E�6�Є<�<� +{�7w.\��*����`q/e[p
�C�C��&.���̼�>���i�١ɨӤ�a�
� �c��޳�(����$�[2��6����>q��̹w.T%���x_�2���|��SG+�g[�$�� ��<i�$���k(�lА�!�͞!Y���/��x���]#vUť��2�rܼO�n�T'i1���{S���a sI�?:h2FL�a)�f�n�E4�*vb~/�&N%�鯨7ߤ�����k�R���$4�)A��b�1>5{��+�Y���i�C��`M��S�e�6�oܕ]ƹ����j´�����BX-C ��V�L͒$M=v�G�T�+HL������q1i� �>�8YQ L�UԢ�ѵW��Sd�˾F��S%YwjF��$L���$�	d�$p�"si�a�eӠ#^Hi0̙���7��d�̰��RM��@��y7�*���h�KO����	Y�>���#F�E�E�lH	e��B������������f����0J����|�L��I������7tMW�3�j��ő��#X��Nw�-����	Ԧ����D�Y��WL:o�@q�rC&Im��>�B�6b~M��&��K��t��t�L	��h<V���f���1��NI��P۹f� �����AZ�q8�E(������~�J�qB��**�a�q�kҢmAZ�_�J8b+�˒$�C���8�Ep
�t�щ��b�˦-˒$�/3,�#b\�d�7�p̐զ �m0Zy>N�
����X5��ݢ�	�����V�I<��lm��6ٻ�(�	j�ږ�6�;s�)+Ʉ�y�o f�f�s�n��?z�z����-\&9y�X�W+���6m�y6�L�e(�����x�M�=r���vⰫ,�>>?u�s��)ij"��.��	��=�aĆ �h��&�� �x�vg�$���@e���8�m/���Ā��I8�����"`�"���� �]����W;�l�,Q��e��V�li��>.�x�pG��z�nR������v���{�=qXV4�p�b'��g재��#d�Q��D0똺�#�x�&C�9fiKL%��=*�wF��9�6��OA
��Oױ̖.fD�p�]�9MF�ǯM�u�w�[�ո���-2��a��KKj�h���-�3�1٧,ٷnL��L']Ǐ���)OZV�ӵV��[,�]���^1U_J��qɧ	ܴv�v�@>�����ͤs!���G�\N$j� }`e�>$a�M��ӂ���:d��Oe�<���i1e�iF��>�m6��(r�ȓ)/�Iu�T�J�]��H^�nn��[!A
!g�!f�������A	��-��m4��+���m �`r Y��mTՑ�����Q�j9-����RlHBE!N1�|�kZsĘeշim�90T�en�9|�����H���H�Zk	��Mp�g@h�׊a��d�]I�x������i`{0�Si��'Mn�M'�0� aʛN[99U�?=w�֮q��z�n\�p��m-�d�$�b'N�i�c���:0�ڰ�V�*��U�Ok��5�_C�#�$����nLBL�ӳ<�yC	Iǹ>L�#�.���5���%��8���PJ<�v&��W`X*D!�o��9G��N��	UR�M(i8�f)�ݸN#��&>��Q6�k�S p�Mu!�a�Z0��$�ٌGtNQt�	I�e�`�x"&��"p� �Q���Q<a ��W��!���'����|:Ǭ��8�:gmx_���̶���qj��*�g|�g��k��D��c�d�OÃ���'�j��:q�k��^.�˶b�t
>�x����J&(��OD*����^YOi�^=ge�m�]�gn3k����;��������d� �x��d68l�<N����pt~&Ჿj���_�~/
������sʇ�x~��3�T�H��;��x,s�?w�d��i�uJz�|�����y�S�Y��K�C�s׆Ħ�wE2f�N{��Q�n��p�^��<nǽ+��1n�{8��(0T����}��˹��~���9$�3���I*�y�$���܊IU^rI.gww"�UW��K���Ȥr���K���Ȥr��%MRMRk�$K<"x�\TZGaG�O��(�op��L������`S�LL�K(�X���r��Hg�$�"KY�n��(�&뼫��>�~U��}-[}�}N�c����6��z[�μa(�L�Rn^�I�=�T�߱.�� {N�)�دc��+
�i�V�����^��J��*�R�`�;�(�9FVQ�G?Y�������f6������-Ʌ�ٙ�[ �BJ�+N���W���Y��˘��h1��e��1�VTͺL�<�>L'�Ӕ�i�9���b}�I!,�Cq���X��M'�O����#��87���4c��b����8eW����:���b��K�,y�ra%]Se��j����b���q؀�󊚓p�)B�������3i��L�a0�>e�F9�"�F�j˛&^�"k�Q���v���J�QP�������Z�ĮL��ȏa#����	�xH��ހ�|���%TQ��L�>}i����9)���Yr��i��i�vg;���cr����G)��KNi&��7��k���|�L��q!�,��l��	fY������d2�ݖl�4�}@^X}�=�&v<p�	�s�.+�N��5���ϼ��MjI!�I�28�R��L���]���h�"	����r$ڕ���|�L�M'M���:�!��q��C����aӵaX�ΕZ|���ߧR4��:�kC3�G����1�w>K1I�!#�Q��$��/=���jZ3߱��Y���5]N��}Mr⟬ڙ�bK�&0d�d�1���j�ƶX�	^�8}W�O��L&ؘ�́ྉ& �4�i9܁�����%9X� $�%�6f���^۶���a&a �s:���$v��'\�k�z��F��������|dr�,ֆ󂊕TɁ9�oyu���c;�S	�������,JL9��0�/1�eÐi5CO_��r�����I	-�߉	6nN�=N�Zm) h6hH	�K<"|t����I��AH��驥&8~c��e�	�����n����J���)�F��yv(;�C�1R`�)�Sp�e�ї�g�|(���3��e�C:&g�U�����jH�ܖ���*�z�t��k=G���%?���?�Ht�!�>g&��;!�e-�|���6�t8�K����ߤ%�N8		.�fR��Q(���tJj�wP��HK��]���UJ��e:�~)�WP�i��9��]�n��$�p�,���n~T�j�H\�|�4��c����o�ܰQ$��o*���si�� S�Ž�L��M�u9̚r�(�4oy��}ÕTJ�H�)�|�l��0IB&��J�J������6�X}Gfx�Mc0����8�q&�t�����$"q�Sn��:pH	��O�n�0啉�f�w
�&Jq�ǚp�y�����'i�6�i�I I5���&��y�V����+F�]e�B컖$Lm�E�Q-7[��k�D7Z���1�]�������JJNbܦ�Li4�sک(���N��HB.�]��m%!��6�%�ͮ��	����:N���Z��Kh�m��4�`ܜ
=CMsɔ��%��6�FM%�?۴۴����>�U%Q*��7�i6��gĒH4��y'%��	����&S.m($ve8����Js�B�����$��H�C�,�RQ�XQ7�ؖ0`�U�x4��Dأ�i�#�D�X~"����OG�W�'��pt>/�^9��<\|C�\=D"z*>}J�|(�N��Q���#ب�D�Z�	�?C���+�#�	������z*t�yJ�(�Q�׆�6x�5G��OG��O'����&�����Qz�U�F�qjࢡ8�^O��qM�&��ֲ��'��>>'������w����`�l}k^����������~_��s:���aϪ8�!JH�?̇՚"?l�`j�\u���]��{�&@���3|��)�#�va!9s��Ä-�.��{g%/�7��[�
���R�}4;y�d�#��b��.����t,��f(��L̡��֥"�<��_wK�⏄����Xz����_���H�/���ŏ��Kϰ.��c*�́s��C�-���z�=�W8����;���!{��Y-���
�Ȯ�y�7s�u3�S�A��D�c�:jd�Cz:U��,u��Xeu�2�U��F<2v۷"P(E�RȨa��9v��^"�d�P�k ˙�kK�{����vn����FU���c^D��߽��M���롋�L��o"�h!Cd��Qy�c��f[���IIfAd�K���Z��8�"Q"ڪE%3@ ���|�&����p�EM!����J�$���W�"I��p��Ҝ/��ò������I&Tp2"AJ�-�RΆ�%�6�?���E��5��v-�E���}���̾9O�I$����R9O�I$����R9O�I$����R9O�I$����R9O�I$����R7:�J(�����J�P�<a���7%�י"�+�b�2i�`��&�$4iTkL�ⲛChX#h?�HH�H� e�e�Xq�"��1��"	r8�68�u�Y%�z�I�JxIycpyH�P֓�k�D��r�O�&0�L9;�`�����Sl̄�:�g�r�Q�7���K����F�N�@��<��5zHXH���/�UV&9&�6�"�ē��x� ��d���e�q=a�т	���!p�^���d����3X̕x/\�N�Ԥ&�ϝ�N���=��W$��"dc�|��`~M&��ZNZP�(+h�?U��3�=2L%�2�fe-Ԏ9F��6�;�6m4�2�L10�~Q�i����{����M����tڱ���r�T*��i锡�GΥ'.�!��q3i��D�aJL${�FJ�	�)Q��d�$����_r������a~N%��8�������D��T7�gOƓ�$8�-"`r{�R�5<������b�1�f(�\/㘻*�&�6�����I
�{���Mi�D���1¾�LC�8��$!��a8�'2/�,~{�h�0�!�7iTPh"c	w���p�|C%��o��u8�xk)�5��D��:������l��(~z�<�!����L�>z���~va_��g�f�j��"Z�p�#��9Qل6F��L�kQ�M�P�CJ�����3 ���YNV���d`���
�}��, ���$��$�'�Q:CJq=`��_&]�ZhL�,M��,)����y/^Fmƚ
�e;Á��i((��a6��!��,d��9x�\����*��bT*��n�JLW�ռ����e!�w*D.��^�N>�69|�6@��� �!�D!���ݘ��e�%L�d�� 窻�%4L	N����O�\RlOq۠�M��k� ��Y��h��c.�24�v�I\�oA��|�����f�����\ƃA�!���^BR[#m�W,lh�@ʔl���Kr���D���&C�Uӑ�	$6�<EƓi��Ѷ�]`!�� �"CF�B��e|K��Y&��r�z �6p��Q����^�6�MI�ɽHt���,>�'Ӓ����.e>JN�:t^��x��tB�>L��[�6�u9��	5�O|\�F��6��m("�[�ʝ䪰��dA0D��3��]��YVB� �v�V�g(,���}X��52]��۸�7#T��{���Q�z��k�Q�pH�뇽2<��C۰��Ə0��R��݄xVSyi��s���Q���d���#��x��'Hp�C�k�W���K�]�HO��Pc
�0����YC�+l���L`��T��|Bl!mM|�RI)�1�O�1e�SE�BG*c�0c�N2"�]�\5f��@���:�RCp5_Í��R}=2�ǱY����|vĪ|N0+�g|M�O�m<V~r���Uz�r�iY,��$'�a�Q��x���.�ꝺ��8O��}�UAVF\�F,^\K�	�8���B�Mi4�������
<@�HpMO��.5��22Ƶ!�$TMK/%��Z%ⱉx-� l�!�-����d8�ޒ�&�f�ǻ�gk���4:H�O:�0>��ug}��$�CF�۴�^�V�őg$����؝�Q����Q�{�I$$�L�I�	��i�|�24y�$��[M0��s�Q0F�"t�?�pQ4(�(�H�Q?
'�$�#�O��?+��{^+��q�+���:'��a谄��D��G�\����O��G�>!���<g���������qv�S�xt|K=
8x�H(�Q��,���q�8�9�l��4�/��g����|4C��|p�>����W�����|t����ڸx�>Hx��g�����p||N�c�qp�0|6>��Y��|����<>~���_����M�#nC�[�#���^{�B�׋X�*���ty�{w��ч�A�-�k�߮^%R5�&�����5-���NHDI�^��\�ա�2����B���c!�8��bc0f8:���Clb�^�z�� ��d�9���Q>>����vk"U�Fk����5�T�l��y�7$S[ǞԠ�ay[���}�5���;h��X��t=D�\G}���vO|��y����׏_w���!йӣ�k׏
�_6�<�i!�����5�u�#N;�={Y~<���L������&fww|��]rI&fwwb����L����#qk�I33;���NI$����R75�$���݊F�Ҋ*J�&�i�QUvq�G9̬Vvr2>�m��v���ٴ�/�:u������R����uG�!�>XO[-K����nʪ���61��<|u��68�s`t�d�0�e>,,��I1`y��9�a!��S)��Dp�&����a�{yw�:/y,��[!	%����A�>��B�ˌ����$|X��;�L�17��U!^��S)��څR`O$��a6|�-2Z@���Y�qɃ��2n}�����X�.�� a� �"CB'���z'����A1�!"ሟGT�B`jMh�Ԩ�S�4����	l33��6]���9�!"�.�8 �R��,rĒj��Ic�7D��آ��kU��Ȣ~�C����0�Hm��aI'���s�$�Lo��J;��^<�y��0|{���.*���鍞M�Tx��52e������tY�(CT~���ڶ��ǳC]��+�V?*�a�#�2���eT�A�D�X0��&�YĬ����|擆���#Mm0�=몢��m$�f�	4�'Ղ�$!ww
*�)�} Ky��N$	�&YM�$�3	:`�q���as	��A�DA0D��O�}�m��2�j�M8%�rZ��kl��w�b�pƤ�9m4�Q��):����!x�&�)���S'ɼ��A�q7.U_r�s.T�3!w���DZZ�����z	�I�\`.Lzp�	�K	�5�-!�ԝ�� XG$�Ƕ۸�{=�^��V;Um���IZK�/mc��i1�r�#�0���'r��GI�Ǽ�	G	mE��c�ar#aYF��s���$��z
*������=L�=h0�-4e>O��Wa�&��0���t�[H������*&��(VO���	�8"C�����Cwm���b�p[�+�&c0����0�D��0A)�1Ą,*X�[k���,�	�8e(����#�0X�0�NF$3( �5"$�BRMݱ����u>��<UN��'u����Fm�|p�KA�}9��4� �
H,��I��<�>HYڣ�ߙ���De��h�BH1��[m�B�%��J%%=��_J�k��<4�m]*����Cӷ�������8e}���UT����q>��H|m���%���I	�����Z��,i-)8~ M~\J�5y,B�����Q`ٔ�d��0c.��t"W��/��Ų���F���P]���1��> ��$>6[4]��}��X��Q��k�����8�:�=���$��HZD�8�U�y/(h��<��q9ve5����H5�V�m��a[�=�U>7�Vx�0"D���!	�����V�ګ��z}Kg��NvJ��H)�!2fOH.eީ�	��.*��3�@�{�J=F��4sa�{��=�n5]���t~��ó�Hm2�K\�g�SIv��a��|!�i��-a��\��>�Hɷ9	U֝f��N!��lM�Iu���?�5��Q�A�DN��`'E
0z(ׁ?
��W���.>!���l|&����+�xzx�z'��	����l�D
'�W�+C\જxy�/���2~^����Ǐ�~_�2pOO�������	
��U�+�xK<O'�g������'������p|?+���b��Q1�T!TB�+����oÃ���G�<(�>'����|z;!�qp�0|6>���h�<�����8r/KD2�e�.�b�ؙ��"<Mb�������oٻ3|J��mJ׭yV�Z%�Nd�����q	���z!���>@O:g.���Ҿ�K�;�!Dj^K{�D�8ZƁ-$���Ѵ���ۗX$�#�'S�|�B���1��Lȗ�Z o�,�J�Q�#9��3���Y��b��4b��m�*("�p��lY�mDg-݃4�!K��K�(T�c!��8R�����YM1���7�����dh�O��c�<�G"�؅ �>�T��?^�ok��.'1��p��!�eơm�Z-��U�΍�o���
+�!�Ⱦ`�L�q�'�-U�A�XX��9,����H��$�0�G�h3���(P�-)�tGr�&���w5Op�X�Gw<��*E�����15�n�D8�*��?V}��CN|�e�e�OL/;[��L�o1�����4��uR%R SQ�5�(�!A�F�G�F�8�l��E~��n{��sDF��$�ffwv)��L����#s\�K�����c�Iww{ؤnc���ffo�=��<O	�<$A5$�F"(h6�ЂEM��!��P�S	�E��j
~M�m ��e�g���`�������F�u�>4�u4L�KM�J	
xp��v0_��'�9DC��ei���Ge|G�P�`N��Ɂ���3Sة9w���0�`������
����PR�,6 �&����Zqy}�z�U�Lt��2K'��J�����G�P7G���I!!'�UB���D�����"�����+t�<��s��y����7}y
4���ډ��b7*Ҙ�(��ϴi�J����N�#�Gq�RW�'�Q���'��xt�t�*��U��.��ff���I��iS�(�fK���(W�;���H|�7O�ƒ����R�1�˻����3N�ޭmMj�ܒ�%T�&�.S�[GR���,��e2�h��'�B|}��M�M�>�(��v�3�h�FQ�� &�����=}���F�i�dʙ��z���j��ԕU4��<Y��sȦ��r�̬�1��'�'��/Ha5E�Le<f��2S~I�HL&�]�$!�{L��>>�[2�[){������#ﻣ�L'��� ��#Δ�)����m��ns]�4F�H6V��:)��$�Y�!��c�8P���P:H�BlfT,٘e��i�KY2XҪ�֘\�ba1`�����S�B�$b0�`�V���Q��:~�#>=7��26�c\�k�ƣ���a��㭘��6�F.T���>��z�q�,����>0�W���_��p��Uc����y⬯�Gҍ�)^)���z�VW.�Z9bUP���|��8��i0�J#��^�M	)�{��s�����$cq"sla0��>rg�f�,���ߔ�?�Tef�S1��`���/�l��M�KN�'���`�O`z�}����V�Cg�Wjq��c/�2r3g��[�+�B����U����d�BQ��2�C<'�<�4��Z��KM�&Oe��D=��WW ]p�!2��8�|u��I�$e��I�eNԪ��~�4/��5O��C����X�
}|�C���5�dmc*#��g��w�DzS�S�f�'�$$�X�k^�	(�!%Jk�4h�k���SRy��䲌$2��	$>�L8Mh����I�	��R�B��i^8�e����ID�)�a2�l�XK����~!l��ל�eb���̣ZQ#��ܡ�EJ6��3���u�H_X$�(�m(������bC L�a��(h8�O�B���>�28ْ�Z��]��f:ִkZ�4є���8X�(��"Y�K������$6�X�ם�B͐��q�@i8����BI	��#�FSG��}s	��z�RK�����e�Ȗ�Ōi!�?	�$]��Q���)���x����B�.ڻ��"�s⫤FQ�7�n��>E]Q}Uk�9��L��M8M��psNo��V�	N�
*��(�f.Q��&Q�owܖI�-���r��7�ˎ(��I�=F�	A�	���8���gn�|��1�q�p����+g��T��+M
Ѕ�b����*Mlٳn��n:zzzzz��q�t�n=��o��;m�lٴٵ4!
��hX�-B]B��j��km���x���6��ͽx��n�m�ح�6l�]�i��޽m�m!q
�BBV���&���Bs�����A��@A���Z���=�f�y���ݿR<�#H}Xel6��0�#K��s5B��^�g�����S�~o<1��خ�U��",����V�yF��Gs��Y�y��ް~-*��yg�T�b�Z=�[�*Yԣ������ȍ�rI.��dR7qI$����H��$����E#w�RI.��dR7qI$���ؤo��j&�Q4��*(��$!6M%�����P³j�9ڪ���\t���Q���#��7G�v����1󙗍��U,���酪p14�4���u>�y�S;��9��JO�NUQ*O��NL8$M����7\�=ĳ.]i$�F)����ÒGFR�=��f���Dr��(zK)�#	r9���RQ��HMi"i%&F;��$fa!����Y�!'�uő!��S���I�ЉrH�/�u<~w<�*��+�Ut��a���ަ����m���3�Fg�6��L@����?�F(�d2SdHdQ�M��IɒD�^|-]20�`2e|�g�X�����M<tYi�&4y9��˵2a4k\�;��IHCm=i��?P�;~s/��Yuy��48�Wj����wӹUiJ�U]1�(�o��d!�����rN�2i8�$�BS�e>͟&�>�#>o]���޽��s���'h��j�����Q�&�˗��]L�J4oU���n��<�-�{	uE@�_i�<cǅ�G�AE|WiԮ+��"A؈�!��˖(	0e����ˁ�zZRG�i���<ui�;E�ې���0�9ٽM�r������NDHKT��A[#B���<)Ӵ��^����p����l��H<Kl�=#Yv�<N&^�Ɵ�G�v¾UW��1�vB��11��zt~��9_pn�F���Y�qʞe��k2���K���$��L�N<L:ќ�8�)5in]�Ƀ�2u;���HH�x�#�rj�oؓ)�?'
ODр(3�a�)�舟�C�o�K�[�X٬�ở�e��W+2�[ʉ������	f?�u� k�1��J-@r�S}�}12����=hDJ?�	��	���C��2�8\�V�X[���Z��F��	1�!!��_ť{[���Kf~�JO<0�Ǫ���e?�"y<�N�Qt�����0��e�y1��M�Mo<��+�͍4C}>�*��̘�y�wڷɦ�"�^��ì�&���mApCB!���g���7t�C�:!Y<4�z�m�&�%��II���(�$����j8O%'S���bS�F��}F��>5�˸2��0�d�xlqx�]�ʷ����p[�)O�I�̍3��n�;GģWD"'	�>!��KL��������L��Ep`L8zd�HtJ���k��-�Q���}^��r%ŭ�!jɄ�کz-�t�Lr%��ׂ�m;�6X������0�N�7P��=*�W����8���H��R�2f8�dHO��j�MQ�ho#�����y���wD�;V˪�.K+�����R�&a����'^'_]{Β2�;����$8�<����2{��M5���Ϗ�l�f�x����t�m�m��|퍪�lٳm�ÏOOOO��\u�x��=q��|��f�fն6�M��,B�u
���KV�+B�yʶ��;m�o^6�mi�+f͛6�ݴ�v��M���i	b>�![_ew���N��^d~��T�['���+��mGC��2�������v��İ�����7I��͈w�;��\�!2�O�i+�V�KL:��Cy���G�D�]��v�8�~y��y��ٿ����'b՟g�
֧��0$`ٔ"#1�۲T�5�	�RJ��Sճۦ9*��JU����h

H@�c��$A>*Z���!B��_��Y>[�ƌJj�Sv�}dya�:�1��Bt����f��%s�&�$�I����sh`�((��E�3*v����"iX�-hmF�z�g.Mj^����Y�$.GM�{�`#9{��&��B��ΰ��U��J�G1�Es�m<�.�+RN7��C4��#�ԕЂgm�YyXf�	,���T�U$J��A��H��>�̒�8i�c�h�
-�!����*M������4Xh%�m����po���������#lDm��W�XT�X���~,Ly#7�*���B(!C��J�N��c|j���TI��iU�O�,�	뻻;��7Ȥ�]���R7Ȥ�]���R7Ȥ�]���R7Ȥ�]���R7Ȥ�]���R7Ģi��RP���!����k�qK�U��5e/��Ye �k�ƅ��Ё��X�:��,4RRH�?�D!�ԍi'��m���~b0I���(Ez�fA�!<�]�B�Yc�領�1���Q�n8yV�g���?ߓ	��ʪ$���S���s_J%J&ͱ#I���T���2�z��ɝ�(��їD���_F�^�Cۖ��2�d�d/2�����*��4�����:xmU�c�U|��7ަ���N	�U�Q���.�l*^��7$��;	�8Rd�H�z�B>�8�\�nB�:E�H3^�R{����i8��F@����UBT=w$�#wW	�����N%�h�-�d��ꣵ��59�B)	�VG�cG�V��*��1�g�7��3/�[}
k(��;G�ī2��ڔ�j�nL��'l�4r����.\�I)����>��H��;G)����h��4h��~�tG���s)��#���vBZtu76���Ն>UWlx�1j�O�����B�W��?��QcW_��es�$�3&b���ē�"��e�u)��wNSrI	'R�:�Mļ�����Y���$��2��m��TH�x�>N�N%�'�C.� C�"p��BT��'��F��FYl�萵�B�i�RU�%�"E�Mt�$!|�*q�#vJ[�U�F����0��̕�U�JL�S���a*L�D��|���0	\��x�:dϪa5xO���Y���sV�)#d,D̻.d�H���7BJH @��8C�!���w�Q�ƢP-
�Z�mm#[a3s|
���ޛ۲���BN���BC':2�hND�|C�Б�$d-(w$�d�-Q�5G7�;R����#.�hZ%c*�
E��ۈI=X�%L�����a�:UW��c�����~֋#.�2`ڏ�Z���T2��'{��Q��j�B@����q2[Vw�y1�4V�Z���.���9sF��e����T�+t5�ں���i�GO��g�����	$L<3�i�u/ې���sHU4��q6e0�CAd���!���ίn�N^jFLbp�t�C�Ry%�L�	Gr�j�6ݩY%��=����B�$�a,���5�)��Nz�UP�&��Sv�borM}���L&�m"S-=Io����pDO�B����m'��J���m�c-|Cl3R�"Ju�J6$�����H�Kf*Y$�7V(m4Y�6��ȘR_"as#Y,o2��#�wj�X��tg4Fl�*\d,��D���u8�:�4�[� y0�d�)�Y	g�k!Y~�t$Y��Z0�M�]7�%�|�L�ˍϬ��
�TZn�1Lj+p��Fg�[�_�������,��;0�1ꪼc�0��������:�u9z`f��
�Cbm�综�$t��M��7��'����z�)�8v'����i��L'q�gc��ęys.A���G	F��ڏ�Tj
VI	6��4�M��I���n�<q^M�>1��͛m[zkk�[^�m�m����+f͛6ڼ<8������\^6��8�q��V͟Um�T�+B�b�yu^V�ūW!��>z�o�i�o�|��]���m�ۥlٳj��N�x��ݴ�Fح�6m�ڶ��m�{殼�ғBD�ƈ��.�6{2{�{�����y/k�)�N�V���^l���y�@����SǼ���fp��O߅%�{��s�w���,�]A�dSd�[[�!��G��J�=C�\�Z���×�Y���N��G�@���b����d#�<1�E]��AIF.~��E�3��8-����c�Q�uY�6�7-�ճE�
���hyt˾��0�m�`����� קԋ���e�ԍ��ݿ<(s?�/O~�K:S���]������]�ܞ��\RI.��OUE.G$�ww#�E9#�{Y������ C�"x��B�j�Źe��,8tG�Y�}�I-0�0�n���M%���ɷ	��s�ؘ�L��R�j9G(�~=�9�=KA�}����BG��e0�h��)�~H�x�Jw�Fk�B��
��ۨ�6���1⪻c�1���;�{�ossz���ʵa�6Cc�SF�#��¸qR`��u+�>�ӣ��Tj2���C%�L/.]�+�w�$����`�`�ZA:��6�8fp�[�Ȓh��|��W�#��FQˣTY������ �[䍨�A���2j�̙+7����kwInX�q&�M�`DR�E��\EcNMTX[%�KЙp�*7]A1a�w.�ꨳg���;���4�L/w}	�L���	�y<��HI��� v��u����$�3g���<dTS�=_p�Ο���W~I�Y�I�.�]�W.�Z-��������T( |@����B�N7 b$����4�gĄ)8��[���F��f^9G��X��cŪ�&�t����o�lv�g�*�(�˻���]�\�>���"D���r�$$$$�i�)k�I}pF�^���G7�H�¿Q��tDN��B�u�I;\���x������}�@�LV+uE�0d��8n���ѝ�ӝ�wm����#2L.�r�k�I�ZK/�x1.��_�^C�O����y�a:�b�	ӛ=r]�Qe�KnNRe��c�����D4C���ؠ�j4��q��\Y*�d�s/�W^��,��	"�@�F��������i��8�"�4x���h�;J89�D���V)��L�pJ���2�Wz�q0y:`�em>Ǔm&ͽ�d���ڡ!�DO�>!x�뛎���{�"�@rSb:G�$���E1
}����dI8���"ӟ��4(@���,l�}z�%0����4�4����1OS-'�i2A`���P�WAtKd���&�'K6ӝ�:�t���GU*�eeJ�3욟� ��1&B��.��!E�|�a�Ĵ���e)t @��D��.t��^^���Y��cQG�X��"��bם��[�-e��d�m=l�ѧnw��#h�m6�2F��A�'�I�l�e2Z]'MOQ*����˪0�����r�U�h� @���>!r����Ƃ:��J��բbEX���^5%�g�]�UJ��lޡ$'+g�z��u;D�H#xK�UWYYCG�Yf��wvd�FE&]^�r�&��i?ri��z�<��p�6�nIR�U�r,鮝9�i�:;;a�6�����!$C�i�5�M]��!���E�ВA����F�P�n�mR��ϯ��^.e���0̨'ƫ?V땪�=n~�c�:a�[��u��^I�Q�3'�9$6D��nzI��SF1$�U��&�$ל��� �B$��I$�UQ(P��w�y�1,|�I�G߸�Y!�Evf� ��&����蔙�������%(��	)�\"�R,��DR,��T�H�B�,�E��X,Q �%Id1bL%�Y!E�QdT��QaY!EDQREYE�XE$RK"(�(�"���(�"��(�(�(�)%�Y$QH�Y!EBQ`QPQcౘ*���(�E��EZ,Q�a��Qb�E�)E�,�ņT�(�E�EQeQf�j��,Qh��YE�YE�,�ʑ�E���*Qb��T�Ʊ�����ҪyGt�J,QeQh�E��Qe�T��X��,Qe(�E�b�R1R�YE�,���Z1I2QEQe(��YE�Ie(�K,��,Qb�(�I,��QQE�X��,��,��(��T��Qb�(����QEQb�(�E�X��Ie(�E�X��P�E����(��(��X��(�F�Z��YE�YE�,��QE$��YE�*Qe(��T��d�e(��YE�YE�E�IeQe(��YEJ,��Ib�(�E�X��*(YEJIeQeQe��KR�J�*X�b���T��eK�,QeQb�X��,��$��YE�,��(��(�I,��,Qb�YEJ,Qb����,Qb�(�EX��,��IeP�(�E�X��J(, 0H1�1 ă`�J�*X�R�)QK)b�Q-*Rȥ���)ie-,RJR��X���--��,R�YJ������e*�Qb�Qii%E*�(�J��X�E,Q,�Y)b�JX��R�R�k�%�X���)d��K��J%�U,R�*�)d�E,R�D�K%JX���R�b�(�)T�K%,R�))b�JId��X�R�(���)T�D�J��ZZX���(�Q,Qi����*�)b�D�K�TR�K�K%,R��)d��X���K%,R�KK�X���)b�JX��U��C"�)d��R����)d��%�Y(�K%*�)E,R�D�K%JX�%X��Ub�X�%X��b��eZ�"�UX�Ub��V*EU���UU��VJ�V*E��UU��Ub���R,�b���UEY*�X�%H��V)d��b��U��X�d�B�Q�`��X�H�)AH�JEH�
����JE�F�H�X%"�JE�R*H�P���T�:�FdE���d�H��PR)"�bIH�JEDR,��r��>������4�^Q����Z��H �`�*�$��!�f�_����f8i�������?���߆������G,:���
X���(_virPI?]9��$4>;m[�ѯ's*c�؟����M����.�?Y��EU�9��������~x� �BK��TO�
0`�����1�KG�nazB�}#��_��`��a����t�F�;@��"��8	�<>0��Kփ�u7-_�`���ҬNt�}�tJ%ʘzmh�r�~��@�'�o/��:��%�t���{�L^�;c[�0�P���"�X��DF��!��n �� �%p,�Uh�6�%+F��gu��ے|�ca�d(� �B�Q�L	-R"$�UA$%w��ð9�0r�1|���ORK�0�A�� d�%�/��?N²�]�(��Q8�
���^��Ã��|�C�<���.��,�W��>nAx���ipQ.� {����;��G����<&��=b*���< �͋��YW!O�ٰ��z�p�.c�@�8��*��@�^��#��+P?6�(t���р��M$�(~��҅E ��i����jI*�`�BU�(�#��?���I�;I�ĳ������JhO�hBpr�T����-��\�x'�ǀ ��Aټ�'OٰFq޷�UD��!�"��M΢ւ��z�;2a��=tM�PL��դ���
&���Ր��<�<�?G�}��A2K"��hQ��S�0 ��B����`��8�{~a��8�תf}����hb�:^�� ��H@�ذ!i!$�b�E�̇��:�v�H��9	۴ �6C=�	S���j٭��k�.p��%���p�;o!d�(�S@t��Pr	�Gp�V��)�&8�S�B�^X.�7l	����?��4N

F)��o��xޚ<�"��j���2���E�����D�qp����S��y)D
�"e�0�ݿ�]��BC�LwT