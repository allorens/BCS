BZh91AY&SY��)��2߀`q���#� ?���bJ^�     ��$�����*4����h(2Ҩʚh�&iJ-�2��2SMX�mX`�jڲ�m���Z�3f�hI��[I��ٶkMkJҕl�l�w5�Y��YFM�XƚVŵK@֕�Fժj���k}�l�\ڔ�bkZ��֥��-����ȍlݝ�Z2tT�:˨IJ��mu�5��Է"���<��Zl�M��,��m�]6k��gV�L;��Z���nE�!�"�lM5�썓[ZS�v���VZf���f)Cc5l�ZҒѡ��N�)�����Emkb�� �ם�dR����{�{{�z=&oFս��v�ڶ2��[��������W�vݽ���ӽi������u������c��]��������U6l�=��ٔ6��n�e�z   �|T�b�T�=���{�zӃ����W��Vz�jHV=\�
*�K�-�
��׽R�c٪U��]�"�P�t�J�JW���[��ݴ1UW{����K�V�Z��J�   7޾Kaݭ�UL�y�!JH��}��}Y�YR�>>���:���&����:��'}vܮ)V�T���ٵ��l�9�|}�ݪ��S}y�}�Ԑ��+｛�>@�UK����u�6�n���c:%�|   ��ꔥ�ն��ﯯ���)��}�Ҫ.��7��_{u:�|���Jھ������>���i���}�J�%��{�J��ʔ���rʓ��W���}ﶕ�w]/��fYZkeU�U.$o�  ���+픏n���eOb�}>��^o�>>�֗v��n����*���/����jS7�z޲��u��>�JS�N��RT�V�_|����N�����ꨊ�'|��j,���˳MU5Q���  �w�m�R�=��y��:Zb�^�^�U%UJ��9��ԩK��=�-����R�j��\��J�����P��gB�{Ǥ��ƵON���EoW^R�V��4��v�M6�ͫ�  ����:Ԓ��'RbL�gJU%#��K���Q��{m��*��h-��{�R��{f��yHN��v��Δz�h��L:kJ���� 6��ɭ�]�֪�ئѬ��t��    {�{X��+UAU�x{����{{W<��U]]Q����WW��%��/k��V�^�{��Q&�=ny*�U�ڞ<l�:"�e�K-V-��mjٻ>   ���Z)Gw�ہT�����v���Ϋ�J�p���`U/z� ��Ӯ=*�ޫ\zOY��A%=��{�T7w�֙Z
�j��U���­��  {��UU�{[��օ�����z�Ow�Z�����6�Wr�U��h��M]��yѠ<=�g�����B��  P  ��RU(h ����2JT�      S�b�I��� hd  S�&��EA  &� 5O�MT�F�҃@�  !(���L�'�z������4�����G�'���tU���Q�Wz�_R�^;{���ۆ�c7gMg� �����3���EE| AS�*�������TQ_�~��X�_�{����?�}@ TV몬�
����d�AQ^���?���&!��.!i t�� t��#�G��K��@���+�S�/H��$zJt��� t���G��I�� ��!zB���#��/H���@�)�:H�8H���+�@��W�/H� �/HC��G�/I�� x]$q t��t�:B$N�I�t���= zH��#��/I^�=!qt�:J���+���H^��!zG�	�C���t�:@ĝ!^���8J(p�����
HU��$:B�t��
��" � !�@C� 'HN� � :@ t�@� ��� � ��C�*Hz@ t�@��P�I N��t�R$@:H�t�� !�U^�( D:J�t�W� HP1"�%:J����I�"%P:J�t�W�
�!�(!@:J�t�P�"��A�I��$�Q�(��AC���IEzB��^��!U� �IUzB$A� �$U�"�H�*��W��H�  :@�*I�! :H��T���S�/H^�=.=!q t��+���I��$zB�!���/I�= zH�:H��'	zJb��H��!z@��#�S�IN�=%�$@��#���I�� �� H�:B��� t��+�W��H�)������1��"��bwG�.E7,��YNt�P�?�����j���h]3�UX��#�B%�f��J:$#N�"�5x%��YL`v��.�*����ٻ{���60��	b�v��Y���(��-��,@�*Ց,�;ƍ]� ���om=2�
�tb�A�F�'!��A\���%�(��Q��l�����'S�VRiZ�S��M��E��ڼ�tl	)VM�ҫ��Utf�=�'�a�l�6q34J�����O0����,��w��f-t�e(�Co~vT]%K`��g�AT�20�QG,m%S,e�M�2���ɨPp�B�S�z�.�I�*�H�E�{�%c�'*a��f&�鎆՟��jn$*�U*]��X�\*Ŷ��t���0
Ȳ��XkĮ�fe�S���TMZ�*t����aB�����]�X�ے)��u1� �⟵�܋��us1%J�X����')}��TjG��y�32��Dv�b:��2���v��&�m��4���1o���c&*­�)AWxq�
�ʩZ��5�̤�ڻ�,�h+sYE��X��9�NW�j̭�T��Ll{�(�R�3rԦ�7t��dę�X3Do*ݝ��ҏ$���*�FTG	���՝��lT �f#��̬Grƻ�	��xi6[�˳vt�"7M1Z��Hu�v���tA+d2�mt�8/AgK�	3�ر�2��m�
n���N�����L��y���[4	�c�o�P0��G\��p1
?��Îb�4��9p�@�]��.� \TT�Ȭ�������� ]�]^J����P�ո�'�ޓoF�[�H�O!�':��(���XՊ�7mݳN���q�a���ɒ��&��cS0Hpf���nY��[�7��Z��cf�T��lց�Ś�ZА"����w��\F���1<si�j��#mc�p��M&U���f���ԩ��hYE�Ίڷ���t���ݘu,��H�YSv� �U�ku���	r�C�F�c�Z�;[�����M�+��K),��媺�.��
��W��Q��n��(�l"��;ۚ1Vf]!�!ti-��=�8S:P�QÉ��2��+K�y	�'�Cu(BjT�TpGI����
;�2�7(�J�,��Y[�-9&}c4�vn����8ST^Ѵn��Mؐ�]�d��d�i�:n�O���N��ڻl����a�ӓncF��y���"ά+E��`i	e@)�%=4� �Q�̡B�K�D�԰(��ڷI��������m�Gm����R�5U�
��q��VՌ.6.���3E�{Mk$�f����&��[���X��#y���]���%I��Ц�=���4nV�,ܚ �!��]�S���eH̑�V�6����ٖ�sf*7�跻Ysr�t�������7.!YNQ9KD�E^�q�suho,�V�	{M�{b��]]ꥲ��6��5�A���U鿤FH^���V��b'T��V���4l�ǟ]�]��Ɛ��vw@�S��K�w��\DRCZ��6vN�F�;�mI��ՖeZ��ҩ*E�4ނ6�n�ݳ��A����1�H��z�ɦ4q�����9u��*�)f�Id���h�*b�f�̕�Ad�e� 7�2�@vCJ,�TN���m��ƛ��%���Q�c���)�g»TD���q��6�k,ZK	�/[l�h�d}���4F��Ba�ib�O�a	K����z�(������1Z�e9���|��}��wPb�0�P�l<�z�5w�Y@e�pfb(2�I���0~-� ����P�BAz �-���B�Z����5��C��0�V:S�m�����**k2�'��*u��<֘3M�li�sX`#ӡ�G��4 �X�+�e�p�k3nQ�2��i4+�N�cB�fL�-r�2�Lh��Ua��lݳWGQŒ-ib�m\A�ܘF���U�!��JE���D�-���a��sm��,B�V�r*t�5M2�щ�~%X��U�)-��,�F��&(��b�B�dY�6��iۖ���QWib�1 ���oEx۪ܵpc�Z\1P�ۏS����
��o�1��W��v55��dZ���n`v�RK),���XR��6��w3뺑%Vp˹P�@����5SYvaK���̻�v�+nSjD�6��q�,��2KD� 8��:5^Jo�+2 cw1�w���\n�&�T0!pS��4�7z��W�d��&�Ur(�P�n��n�C�?$�� �u%�P��Z�(��ܩ���,�FDlQ81�Z/RxC�v��ۼ ���BL�$b��ɋ+BWyn����Id ��.XM��	`̬�.EPj�N�-5d[М���kU ��6c��-R�I�ڽ�e�����nEOd���V�J/�wN�4rݩ�����h��J�2��.[���ب��6�����q0 jn[f�R��[��N�Y����|�.`�*�a�X6L�^�`�NP[Z#�
�f�5	P��+��ܼ�2�J��u�0i�RT�y�[�S/uX�l�{GdҶ6 y5��T{��+L;�+9�.�5��É�{�J����\����d��	����*n�t"0�Z̗%b�Y'F:�.������'11#f�na�)�:i�n^K�M�\�(�H�C�jY(���-³$ܲ6�`��G�W]�ԕ���0B	ӑG���Y�X$#Kd����J����b�Ø��;OD@l<��gM	0]\�gh�qI��s�Yd�U�}�4����ۂ"�ʒ���*|�Qt�^lN�:���BV12.�"�e5.�[�h�fG+jŉY[��=E�u�=��.���V�0���B��Q�T�'��*�]��*���:N��7�}�yE��Բ9ر;�C�iҤdk� v�h�E��Vֱ�՜&�[�T��6+jj�;������"�d��!5E�Y2����b�n֕�ᎵM<�m�ո�e4����5��@j��V��29�j;��@Tb^a�(���쩐`Ʃ�	Mc{v+&A�&Z܁�tٴ��A�o2:Ǽ;���w�<�F�aݬ�56�� V�uS��Y+\#q��7�.ؙǫLF��F�\���(����[܆��C��d�:,U��l7�^7 :CI�/�[Y%�A��	X�`ynN�"JU)�[X��%3l��Հ�]8]�1<ym�ӭM(��pLX�"ިQ�����=��;�t zn��l�Ⱖ
��nD�v��S�xL�w���(�դ.M/9
�3T����U퇗O7�T �.��E�����q�r
?:i]*&,�N���{ER�X�Leav��dN�E�5���Xu+A%��
�t@�y��cS~�Ϋ���ͫø�#�!�dɑU�֒����Q�*�޽��h:F\،{%�xj7��d] Px�V�u��t�Ȓh��W�i+hK�lŔk+-�:��D 7d�hh�n�� [�e޺3o�,ݽ�ԕm�y��B�V�nm%��Y����,�bD�cS!4<&���-�m0��2HȻ&����XFc�-�b���憧��0��8��B��zn-P�7�/�Tٳj9Pmh�p��"�R��Z��-��ݙ�B.��4�:ոѹ�J��<h�Y�vS[���&�2��
c���r~;Wj��d�E��Yb�Ty�Yt��� ;�$�惚E�QюL����eVQN��,
7y��T<�p!..�������}v�ɘÕb�|��J8N�F	E�� $���V|N�f,V�d�f�fh���Cb�1*Bb�v񭖀	��r�eeд��775\B����*�f)u*-s�Ր ��6<[y�L�5��z����\9t�-ԙ�C\Q��G@�B����T%^7�����V�y!�#`]�+CWj�b�щР�)M�����f��v��0ۺ��0�dǹ���7"1��tV[s����J:FZv�h�wcC�r*�I����Oҥ�/����o�@e�]�Dn�F)���fP������R�l:-�5��we� "a$�	�w.�Xآ��0-���
Ӽ� &f�z�m�w�t�n��lkô��M�6�/�%:��0��1�w5)%�R�e����[j�Нh�dttVZ���#Ene�p��Sp,.����5�Z�嫑@ {�V��h# ������L+/�R��o!r
 �K
;V��i[�&0�tn�M�ʆ�
��u��n�Ʌc���[��U�д@��Ei���0J���n����!"Y!b�b���[84V0J��XmaA�kB�/]��a��[k�Z~��*զD�������f�j!2�!wo�Xd��GF�*˄����f[B������2��O"i�X2��]0�5�V(�+%�ި�Nk�8�V�t S;x���)-�+Ș���X"�KS�t}m#6^�W�Q�
i�Q�O5�G �*�D�n��&Ű�	n��.�ްΠ��&��K_a�.����H�,��d�J��p�GD��JY&��e���Jr�+f�2���s(P���.f�h_�f���󩄙Q]3v�27F����������I�g0꽼	jB"��1����/�,�Em8ag����8�6'0J5-E��{��s���5x˩�n��Qx�ъqn�+V�*ܷ�Q�ZB��#�@�0���u��r��-]��2��-T�·i�vw��[��f0�XjPSustD��A��M��nHԺp1&�6�x̥�*�e,���L@ؤ��2hbHP��ȵ`�,�I�V�� �IAz���wZX���JB�j�g>j���(�oʱ-��J�����T%�z�ǂ\Ȇ1���V���vKƜ�ᥓ�E�䨰9���&��r�	�t`�j9*�'o�����U��ì�A����[��)���C[I2��[�f�MeI�e��.m��n�%��	���9��@�Z�����-t�w��JE��w6�A�So �f��Or�ք�� 
�ȁ�gn���m��A��zƳ���c	��j8��Xd e�i���&r�IF�p���ؽ� �!�n�	6����3$V�����q�iԫ��)D����ϛP?A(�s1��@܌*��kA`Q���Sq1E�2�n�C!L�ɹ��M�֩�5�XYO�ou�U�]/��P���b��ء�����mniٮ;��JU�j'������b7���[�v%�('I�����2^�(�4L��D���+e���-'@�R�X�N�<pF�Ė�W�V��z��r5�����N��J�_rع����mA�r���6i��ye�HB�`�4nkpf��^��9�&k�N�y*�c){�VOY���U�V�sEXT4��i�76��P�M�C�ʂb-��Ukea�͙��TnF.EH�m�ӳ5���9�ܐ��3t�i��-їb
��P<G�`��ہ�n�t5]*�V((����Դ�ڭZ^aР�f���B`�a]j��e��[&�V]��R̷MY���ՠ��4�"/
�eVZed�6�b���P����×D^��mӳ2I�)q9Db
�jj��a��o����[���ch-���ڗ�3U�P��I3�٭�l"����P9�՜˅:���g4���U����m��,P���*�`���E0�1&�6��T h�ct2�LYl5�Pś�*�i�j�ĥ�SA�SюgdU+V%�-�yv��L��`NTAT�$	�a�~���E&��xdUu��h%u�fX`[Sd%���krn1s&(rЅG�M#n�PY%ˍ�Ed�\�����^}N�V����e]:J�E�ܕj�́mG��X=o����W�<�z�F�we=6��2�?7�.d�@���!�����[wA���i���۷�킘��6ɂ�{���/oaLءpZ�",�jէ���53?bժ��ÀsWqG��F֙t�Di�:�у @�,i�u�-�͠^Y�jԌ�,�"��S��#EU�6Vx�ohn�Z�K�rלxiO.�e`R֛�T��CU�{�ǗW���k��m�&I�+�R��B�����,��fӛ,����J�o}�ya�oYթQ�jM�S�%jh�m���K̎�l��$˦��8fb��42��
���.�E��P�^=+ �2��S*��+r����nF�! �,u��f�C4\�"`�+
U��[7�@a��z�̣�pʨ�͕o[ b}��ͣ�5[��rJ��`c������XpކD�Z��M���Q���{B�C.�=�5��P�D�,���-����w%�˗�Vڣx������Q.��J����4CD�"�m�(�@�(�'FV���nS�<v��!h*�9�6�e�U �D�J�-TSLJ�M;�x戣o
��N)��6Ĩ� ���ucFا�)<!ъ̽���`������; ,��b�j�*9�c"�WCwH2��cu��Q����`�ʈѵo+�*1�	�y��Q����T�i���,�Y}��:�5��7L\���V�:Fc�9���ͺĕ�{��t'd(�'&9���H!z�idl��mF�wq67$�ؒ沩�
��w&��/i	b���F��,��ּ�N�4 �p�ǖ�.CkJ��ƳF�f�4�L�ZU�r5�)d�@���b�;E�	[*����֊.D6wF�iM:��u�	�]12�	�t-����:�V�%���7	ש���9���8#pj��	[��(�E	/Ml-�eK�!BC�{W���R���K$;�MtӖmZW��z���e������]��y{���!���~�_]���7;÷�o:���ޫ����{	h�p�}ll�˘0���6�;�f�9\"J�h���(5�0���v���Y+�qR����_h$���]\��.�N��"]nfG-�(�leR���a*��vk4����r}װ��2�l�GU�T��vK<��c�4)�s������`�LU�v`z�g/ٿ��a�����o�;����e�pL��h,B�����JS���öt%DQUx�$hަ�S�i��w���c_"�(�I]#ؕtz�P�A���WV�+���ln*�l��6$�]5T�ɬ|)��.�ft�&�[u�#i�ڄ�[;GM$j��w�d�tT��f��SPڮD��f1�e��aMǷKM��I��9�'�
ݭY��v�]��=�O�*w/�%�~�e����;�D����W��*�u_[�Kw*��v�:)AY��t�u0$����v�{3&��L�5��(-���e�ծy*CCJ�����J>������c���Q�e��]�����?[��H")��n�oR�+��c���amm����v�o_D�v��ڷ�r,p�8hc�ٔ�I��y��]=��-��ΒpW��:��4�2��չ������:��v��2��x��SVu��I%�ʴ^��R�����⹍ا��G����h3��RT�7_��s.T�丨)+w�#uv��燨>����^-~�<�tF���n1y5s]+l��ie�^� �q\�:�]��L7r�=Q�C)W�YRs��0d�����f(851���N�곫�9ARÃ��-��`;7\�gFS�[�t}�5�����*�?�{�dI���>���;�R���j$��ȓ�ޙ֯�n���fKj�r��8�{\�.Z�Gv�`;ز�J\]A�ʌC:�ձ!P�8�LKgp�+4�y����KV"����	�]���-p�Bk8�܎����eFnq�ٓIQ��X;g�݄CF� |*�t{L�SU�]1�6]�;!4�.p��ک��\H;\���D����wS��S�FV%s.��U��C{]��*��F��í�\���$�g
]�)ЍA
�Є�4����x!��w�s���#S��댖+E�9mQY��I��.�+�՜Y���+��n	)�]�.wS�kv5qI�*�Nwl�'�x�Ĥ3��]cэ�S��ol���ݘVû��NQt%7����n��e����<μ�.�{a���R�T�K�L+RG��`:h���0��ra}�Gu��iXDr����c.�����K���+������Sy���|�{�9�d���LjvfV'�XαZ�6+��MH�a����Y�>q.y�$�t��'	�z��f��]����}��8�4��t«��j#x�P�ӻ�Ğ�gұz�z�76��U�'����TK7SÈN]��gG���VKE�]Qd\�{�h7H�se�@a�ˎE�K��:�	��r�V��u���Y����+0%�M	��]z���JR?Y�bR����6u3����P�D���D9L�6��� &­��2�Qg���!k5"/����.������[�����f���z��n�6r�	�O�#1)��ٷ9���1�|8+�Azↈ�u��ou�Y�I�:���'S����-��w@gO��X��vO�\�����.�=��9k;���]�E6�u����Of��Wٙ�*K�)�/L5/\v�A� ���`kke6 ��tgS�t�}6=㴣�2�V�8İJO.3�h���)V����uG}�f��!�l�-D���5����gBWjSx-5u�Di��}��]#O5�1gݜ���]���L+����p�v)s�+x�r�v�Ď�`
��Y����c�WFRt4l\�p٭�ȳ�ٵ����s�]�����Fs���Y�e��V
��ڜt����*	��r�ެ���E�1\�]�\;y*��h���'��e4yp��zjm�\A�6��Vo��S�h �5dˤ7�v��r�{�e'������J��le.�:Nww�CSm���{�&ˍ�V�t�xf�X��8�$Ƽ�g��v��ِ�n_f) S�4�90�9i6�Uu�KQ�Df��"��|��nXB�e�y�\�Rl��5�&�u�j�X��;��K'.|�Թ{�NL��Y�}B]��ke���e�EXi������u)�2h �M_lq�ֲ!^�헂��Yf̔�[�rd���>cn���?���&s���S�6����h�3�5�]�0����7��Oo,��=�[�.:�T�]��)�ov^n�˺[���γ40���U�[����I���)����C"ש���[�ر�0���
��jՓ�1nj -�2�X,���k��s6�*9���kt�9���E��X�S��L4�ԫ�U0�l��nY��7�.2�!�t8*ޗwJ�)L�Lf�h���*v�jVo��������s��\�k0�*������rܛ�
Hn�g�������r�I9,Jj`��m_l�����G&1��ƪ�"S�8���`�&.���'���B��u̍X�-�y����16�]Kox��3������A9Sfa�uIe0�D|9�q�ϑ���u�-�4�:)�Y2�,1���eD���X1�˺��<�g#8�E��GEQ"lVSdd�{#�}��5:�j8OT��և7�]l��A��VgS�Sb�Z�;��ݾx9�Z���Ռd/�[�`L���븝�9�e���Тnd�c&�Vn.��A�*dR�
�F��͖w:˒���5Q��rG�u��̀q9c����+|�})$�O!�=�ץ2���ȘF(I����bp���oc�m3CWj��C�sP�\�w�������x"�f��p���,�Fk�fd��m��b9���h!S��Yկ��۠�i�sH��i�t�9�[ԁ��v��r*�p�N�Oܼ�S�֯�/�.\0[��4�3Y���++(r��dF�S�k��Fm�h�6w.�`Nc1�$�dbY��.ģ�
��u�b��'s��X�V�0[��}(���\,��A��E*����zm�J���䢵t�k�6�Sk��r�G�J�R�3rҗ��=0[·UD���qDbI���b䮾9��|�.iG�֌x̸$�Y��T�l���U�Q6�2����޾�h{�Y�F���w���{���}]y@���rƁ��7�>�<�㴍^�V�Y�I��N9��bag=�ʼy&��<WO�rnڶ�dd�j�WLVaf���a����WQaaP�;��]m0) ��͘��ľX\|j
�r�J�8;[�n�ܷx�P�u9��4��/��E� �@5��spd�;%N^��0*o&� �Q�}���gXf�o���2��c�LC�sʼ���;Fհ��h���`e\͆�C��ǖ@����e�y��O�5W�Q����C���$�H����0ВSlѮѠ.�х��PP��tqn��ųY��s����ک��
�"�̖�䳺Ŝ3�`^[�U�є��Aq��=��9�{�(�ϯP�Nq�J��+k�z���<\��+���p�� `X^���:O���D��c�
��D����]�\N�7y9���kra)L�S���.މT���*�Ȱg"#��-���������nNЦC]�.��(�J�N��M*��eu ��"j����űt^
���/6�3�E�+�`Е����a�H]����T[�7gA��0W���tՓ�M��]\:���w+8wB��hn���vD!k��Y���|~�bJ�soot��U���&��]R��q#���[�J�"J��MƓ{���ؖ��y(q�ʊ�
-8���5�%�X��|ݚ�b�4���l_y@�2u���S��<1��k�����|�y�"���F1���E�������˜ٗ�L ��w@݌-�׵|y�po٧�/�����!o�������ٜx��|�������.���q�x�����=V5�w�O��̄��1��e-��.��մ�j��^�F�C��+{n������� ��:VU|�t�+�xj��ŭPm�lQ�&��3\GK����Q�s+9b�B��]s7�7;މ�]^o�m�^�B�.d�mX �?]�Dl�f�2��߳�t��K�3�<���j���շU�����齺�f��a��N�L}�U��̞Yd�\�%z�,7n�f��R�J�3��U�#Y���Am(zJ�@R��*�豌P����N���J>@bI��J�}۽�y����$0�y�pT��z�\'��3EnT��2�\4��>[&��5�]&]2�ε�T�uwVƦbٕ�.��+y���]b�:`��YU�n��x@�.�no�m�l5y�t.��vE(-��,ıLDQ�ګ"��3�ʒ�:�֋�tʡ9ۑ�7��/n�f���k-Joq�<QBo�s�1�]w�M���$`����3��"��i�%
�����\�*�����w���aWt�W;*��Y�I��MX�r\)�Eʷ��Ŷy�$��)��Q㋻9�����M��[�@�u¦
u�	2���L�V�X�2?D2�U�u^Q��\.��7��*0���v�[�í����E)����)_({T�X��ۓ�ۛ�V0s�v܂M r��߶�2��ܕ�+ �N�<Ɖˡ��mp�f�e�u�Eom��V� ,<��`�]w�o;�)΅\x���i����+����s[CL��N��.�!�e��*'Kõ}ё�R�5y��I��Z�2�u�c8�\�1�%�;��X��W^�r�z�VS���b��p�/[)��u{���N�gm������\��g;t��c]sF�8=pn�)h*A��`I��-���l��c�a��X��ݫM��y�Υ�e�V�;���g`n�̀؇EWMW�'Y�.��<���� x�mZd�u)�i�f���
�*km�S��ս��^!o����'c��]e)]�m�T�=���X�k��G���/n>n����RXQ�.ѭ�/F`NQ�z�e�r\��$�R�yT���4bT=u�9�n�^��}Is�PV��3%��5r�����r���caF큵�\�+n}�n��sQ׷��%;u| �r�-|*G5���e�ý�(H�#}Ք����)���}`�4�-�s$��^.L<�]X�gV��8�����䜨�ZgvZ�2�7:��#P.}�.�Tdv�Bh�k9����2�=�s��Fc�2L���o9�Ҽ�S�V݂�hu�3�}}���#ٜ��2�$�,�F��x1N��G.�vs�p�6a�70M�7��
ɫ��-�w�p��q�xWJ{��(d��t����҉9��.�'��oM��/F���X��YQ�Zha�v�X��x�X6�#��6B���\\�T�7�OYe�y �wx&RBZ�֒4�k�{�`+5��M��:�S������A���j+��0�����v���_(���n�6�B�R�æ]-��f�����.�tA5)ۻX�N�v�dK�Fe�+Q{��=��E�$�l˪�ā�r�^*د�^�a���`K� p	����:ĈT,Y�n��}̮��J���^]���l�l�i%2�pd��1�;	�AF�ЂN�_X5�1؎��Z��]K �Ү�q���G�8u�͋�[Ĥ�1�9��#+AWV���_�QM�9UЧ����L���l^a�E�n�DȘ�s��퓱��A.
�\�<ڽ<Kn��}@wF�b��q�H]'��u܌ԹP��:Ky��X�*]6ƌ�6��Cy�,��k���y�t�Dt(�|����Q8�ٗwD٨�SSbR:�v����4�?JE�ޔx�C�����IX#|�6ּw]�KQ�ɝ)�<�Ds;`yt�pHL��^t��l�o���뇦9��������'����p^k҆hL��}c�j䝱�+"Z萘Tt�u��������A�479jT�L�E[-�H�|���4[����Ŋ�ou�V3���`��
�ഃ)���}t܃�x$��̋6��ʺ'�v�nX��L+��V.�o[�7L�:j�5�K3��k8M#座on�-)��p�f�}n��PPgM��m�뮠�K����o
�W���;�Ѷm���]`�be��h�>�R�]m��r+e��]å,���7�VgwSY��p�`��N��V��v�U>��5_+͸5�8���b�3����t3�ꕖU��&���9F�)kUfIr�饄7F5]���%��Ȍ�t�ݝ�3Ep�n�Uf�ռ��gu�+�		����[���JjЪw��4�t��bipq���=�s&��',C��H�^�V�-t������J��:&��x �V��z���slI-��,�xTK0�]��Fv��;�<�˒��b�+:ޭf���4(-i��2֊�xZy�6�MΧEm�ǲ��Ŷ�>�ٚaƥ�ko=}�-��uis	[�|��ye��f��0F�wY�.���m�:m%;�
z�[e��mbm���{��s$��ٓ��1�Rw�euom�.N�b	�۷L8)U�I�m㓌:i������b�z��4��܇���Kz���Չ�=}g�1���XUn�p������AQ$&B@[f�՛l�m�����f��IB�
"�&��t���x�!4C��:��JH]��9�٫
�P�E1@U5MV��@�i]�;���hݴ���T�.�Ux�A�AR��iiRHit�� s1�B��h#@%S��f�+X(Ր�2�(JZ'�)g������ю�� �Z! õM�UD �:©���1�B�� �J�@Q)Qj�j�
"f
0	$!aq��>Q#�O��A ��}�~� �/�`�������q���??o�����'������	��AQ�`:�^�b���-���^*��9���1��vK�{@�����R����-�Z���9]���//K����l��K+���eͩ������� Yc���7w�M��u��9��:q[i����KlW�Q$A���u��eO�R)Qפ�'^����Z��C�ː%�G/ ��e�1*f"��%ק�����YV���p�jR�P�Ͳ�r�"p᮹�aN+dGi\�δ%J�ѽke\,.{�ǹ�I�X�#�V���O�]��@�Q��,��5�����Y�k�C��	��+�[K�*I��U^qJ2'�u��J�����ݫ������T�4�U֜��1&2��߳���+{R�T���B<N�èP�y/-^���B��n���Rq�C�0*p��(b����+PۀC�$���u�w^�<&ޚ� 'i�T�A���Vau�wu���Q�S����<39���
]�.���>��́���Թ�`�bv!�*���&�E���
�F˕��݃��f��*�w`y0#���31�,r���-4;+<Ω;)!����(ޛ���r��M.O�7���aӕn0���;j�'�K���{�t���|y��C�k��f�"�_.�$���:˲��8�I�c��-��u�fp�w�,����Ө�h6�	����� �0�`a�b0�1�a�,0�@a�a�0�a�b�!�̵6��^m�N�}��(.�G.�X�&	1,��x�
21��ĭ7���u�j�Ó�'m�FԻ��/���w���C����=F�VP��Zy��WO�Jb��k(�l}���O�}�j�Ov*�2�镵�	d���^�EB��K��$}�+/q�Vp�JIB�K�A���=��fcV��}kV:m^�Z����&����V���G+-��hfcs�-�f�A���
.ÚK�	�����ݴH=]���]֫�"̜4I1]�Qo�³F��5�["���;�XI:{#J�شhlfD
"U�D7iY�n�t�W��=�5`��P+qt�w)�^Y,j{��M��y2];Eх�oj�Z�߫g`�8��;��0ur���6�ww�9v�lÏ:+�W��v���u݀P)U��|�rw��Q�6�Z�ٳ�4�:jb�F�M���w*��:�@��Z�E
(J��)�� ��y�0hV>�.�Ɏ�g@MD�m��t�t�ܧϠn���l꘩v����6bT�[[OV��X�p]��J"�іf`�ss��|]�]�l4E2(��p]9��2a�ŵ�a�_vd��b"�;��d4lL�9��Y�>�z�|��t�NT��b�G)�s�abU6���F�V����`I�>�����g]��ux��ScJ�p�	��|�q7k�Uet5��m�[�[�:s�<�f'�M��lZY��!��hb0�a���1�$@a�a�,0�a�a�0�a�b�1�l7Oe�V�^ӻY���+t�8��*,f�7�)L$���H`6�����yr8����r��Jĵag��ńq(F�oiRH�IF��g	IK�E:�Q�!=�z�3e�Y2ZP%Ѱ�4��X�ҳw�ݳM�YRs�":����i fn��'Ʒ(���Ё�g�Hզ�<�	��x�/u��1�"��j^ϖ��9\���-��;r\�zgt��t�c����*>U-N�1��Xt!+�e�P���Ȧ����POn��1�m��V�nB�@�kt�J�buݶ��Pd�i�N�ۣCEv�Ѧ��)�8�0���+s�B�ۙw������V��v���A��C P<�7��r��G��;
��~%�k;
JN0����+
s
���S2�!�?k���Ǣ�D*ɧ�*�_0S� �^q�o��y׹���]׉`�l��u����t�̠�hk��j��/=eK�ϊ���l@a��h��˖��ym�K�╪٩1�ǎ�ۏ�[A��tʼ�ڹ\"Lj�
��Jcp5��i�����-ъȌ'�-��p*�v��*�[j�^r8GN���3��(n+�*D@k��9:�EP�Z��=dX�I�`�v:g���V�]ҵ���K1TݥO�By8���'o,o7R�[���5���)uw���W:aX�yGr >��7j��*�ۆ9z����(R��DXѢƍ`�a�b�1�bH!�a�a��0�0Ɔa�a�a��ȿ��/X��ׂ�p#V*F�.�	��v��
*eԶ�0V��[�isV�賅�[�2Ѹ�6�A�W΄�拺X�
:|�f���P���>��8Vd�ѽ�Lu�G9cȎ;-8���^eH������L���T�R�P�L��[e�V�r��l����K��n�f�y؄�[:��F��˸4�2��f�!Ȱ��Q�.�\*�e�� I���m��>/6��?h��$%Vm�k;�M�/��_9&��6���������|��b��2N�i��L������.�u�S�գX���iy�Qm�,�[��1p��]�7=��~x��RsEi���[�"��FQ�׉�)A�9�:1�,U���z�WI�a=�9f�3N�o oh��������'�%]�vY�Qa��Н�f��<E��	���3�\�!�q`��TsS��46r8��u�V����AJՕ:�iS�qĈ���X��K��\�{(V���XG�wV��X,T�H��v�!��W��,W|�8
e�Vl��E܀�"��������V,̚c�^�.��SCZ���̜9�8T�X�R�Df͏U�ʼ��w��X�
S�φ�Blj�	5�m��:���غM��]�
�x�q���>�BPA����Ϭ��4�Ӄ�,�P1͛��x���W�4Wu�#k/�'+(41��a�a�`0�@��0�1��a�a���0�0�ha�N���J���1b�N�f�9�����uG��T: ���ܘI���ލ���u ��z��ܻDe=F��ct,����s3zEPU�ʂB]ț��_t�n�P����+N��s�R�U����K�'��m"gf�(�/鱂��6V�
L�&�m�m��vU+2K�u�z�����ݲxN$#t65:[wm���`%ڪ�Qm�)i]h����h�uZ9c�.���tb��.t��LV� �數�Q�of�2\��]qd���G�60Q�1��������7���ʂ�֨�V̮ ZA!d���F�=�%��C3�]�2�^���a4\��MI�� b���˺�c�:�5��/��	u����48\]�EY���jB��}x.v���ha)\c2s��WTO��<�R�K����]����X�Y��������՜̑��e��J��E���b����T8���Ֆ���V=�� �� �f�ӝ��z��}".u�ݜ�SW�k=)�Å���oFZ��Ju�� �hR�ZV�*X8�	N�N)�z�kn��ˮk4���'b����2c�Gx��ʽq6��3(�t��N��35=�q�k4��RRŢ�A@Z��ͫ�P��En,�B�e �VV]�\3v�j3i����pk���(Wu r�<��(ΒVoU�w ї�W�XhK7�3�r*MRP�X*��>��96��z)�v�q��g�ʀ0�6h�(��a�/���*�/C�il�y��X�qV6��͐�s��1={ߊ4M�I6l�բ�KL��R�3��Zn
.®Ί}�;>�$�7��l�ηb�,}4b�ˡW(8Yt�J���K����g��6�[W.V�@y��--��b,�*n>z�'(�2k4Vp.�i�J�
���Ɠ8�e�,�r�vQ�}{�֥s6����rd��]��=��L;�qvhﷅ�>�pX@18��Е5N��͔[:�yPNT/�p�gdϏMpl劝qr�}���"\n���hQ��N���[�+qD��0rX�0��X������!�)[+eB���Ab%k�5���('Bf����������ԝMtu"l�"�4�*�!ῖ1���!����7��a�եt�>��X}����1cӽ;�\������1W]���4'�����w����2�%J��o����5�֪oL��pu�f� ��û�1�2 g_����"��<�b�L@̛;J��S.��4]��&8���Y�?n�p�`�(���I.<l{F�� O�خ������w��;��J!}SO���z 6�GX2���PR4 O���9z�T�6S�x�FK�ӕ��F�����vt��o�.�a��IPW��z���dÄ���+C��{��Y�;����]�ۦ���Z=`n謇�鹀.F��3�^������BF�c�`r�P��.�g��t��q�s\��u��M��Rۤ��cY�wB6$�:�x4z��Y�s��X,�U�ΎG5�ݑ\
��W�9��{�m(*j�ut�f���k'���M�|:��X.�haO�W�ǯ)�z��e��f���>�fwS��p`�`�mĖ7n�6�+ȑE(9����!ت��|x�Z�\F�[���ꘄQ�˼J3���[JU��e;lh�u�]j3�z���tH�qJ���,O���p��s�/R����z��8�	�	R�F3U6;2�F�|�Y"���̵q2�+�p�A��r:z���.j�/3�����y����6�D���,�҉�ͥ����|�"��噏J���4��Xtr)�wq���-O��r��v>���+B��P�&�G8Q	3xx7��9Xv(�6\Y)dht��Z$��[�re_���iu2	e ��.]���{1��2��%���Qw�����
�\���CJt;1����5,�C�b�S�n�GQ�cɡ��vl���t9�%w&7�[�W)e��E���<�s>��Y�U�f���(<0��oPi�|2��'��C�z{F��Lٕu���]zb������X ��	�,-����V�`�Kܺ��&���O]4h�����K�|)K�퇛�WV��ťH(�@|fA��Y�OV�3m�O��+���80�;�"��Tē��n]�����#b�S�Y0�L����h�ј�*� ��EYR���7@�X��PIKe!t���\�[�I�w&=���c�S$���$�$U�+�OEJ��b
N�̲��5w5:;	F��Y��ndxӽb���%]/������眭VP��٣�X~�LA�`�'X�:&��0ܱd�	�x%�Q�{�Cv%x��T��ʾX#�S�ct�媉�X��Mn�eBD�.q $2:Ǔ]�V����*��:u+"r4�9O5����:�� �aUې�.�ܦoՑ9�cG,�7�r�1�?NeN��O��X����(G�*��.bY#�n�e��c�x�/F(�.���P�
����9i+�e�z�FcZP`��Yf�咄;�4)��U�Y�0�.���FCM�ݫ������в�3�>��U �I~i�ڑI�iⱙ��'��G:�|���}�d+8����^9���m��m	'u��d��77��$�G���T1�)Q�m�`Ti���?k�2��3Y�p;�:�&E�8q���)�Mו��B�SW���q�)��`��גt57��Y���*Ҭ����c�q'}(̺'d㚕����[����Aa7ʱ�)��L�H�	-5��z��׫���Kɸ��_L��P;W�r��ήsp/�Ծ�R
*R�	Z;�uPP�q	f�5��wk�[;2e�)�U�9x�n���ڮ���vv�������G�+yW�:��F��-�]�쳲�0�&4�"eh+����T�7Å��*،���ܜ=OS�++Ly�\�@eٰ�CZei�#�!V�1������@����F=���Y���lǟ�e�|2�K/��skQ��㶦e���v��ֹ���x!H0�xED��������z9�3Uv��f�:���,�v8�ՠ�K�l��ؼ۔wUƪt���/���E� _�.�x�;�w��E��p�`*.f�:"�o�t��%��F�����̣]��L�!���X�'bZ�gq��,�z<��1ǲ.ɑ�v��j�*-x���2�^n�����f�%E�-�7M�ʛ�ef�{%_���9Mdxrمtۓ�+]��7��N	�Ty�_lW/��itL�������|��ҵ|�Sj�P:@� ��R��b2]�jv�
ǆ�c�f�ӯ��R�C9w}&5i�� =ƖAo~?-���Eo'N)SY[�U؎�2V�!�a-�;��Xv::
i�$�:b�L$�C5��p������<��Y@b�o���݂��bo�G"5*�:�_[WO���.�9�������{an|�7��(���ڙ��R�&��t��.5�r�:�?`uԫ���,�W��>�nr�rk�|���k��([��z1�a։��N��Y4�[���Bh.�N��WSIutsb9iwr��l��a��In��ut�Et�r}�t��٘w�qf�	��WM��X�ܖ�e[�Z�{x�v��J�]*Z��c�|�U�VP���M�J�]��[/	��RV�W��P9��f��+�B�i@5���6���K,�y�ӥ��bx��T�J6Dqh/�Yٚ�ahk1�7S�n�Y�t0�Cf(`;{�w�S��"<�p�R.�5��,dmaU�j���d�5�f7J 0Tj��A͝��)n�M�*4]��V;G���)Z (!�Ukܺ�s^����m��7,��=!��7Pb�+��tue濭�XPl�R�B�IK��CJ^��T�ee�I��K��G*���eW:�BO��7�acw�/���6�Y���ÕE5i6�����2�TI����C��U��a_�����lc�nvRӮ샡�^ܒ9²C�a��Nb���i7m���엋CW5���I�!]�C;V�F�������)��&�V�M��9$%��iRssl.�GEd2Ӻ�\�N�2i|4�ۭ�D���Q��Y�>~~<�y�������UE�A�������/�������g #��o��߹��s�`�4n�O��e�«QFb�ArPΛw��bH���A4eZP�m0\���
�}B�jL*����u�h�H,�ڒ~����R��w
I��)×�ԷR����1��wS*c�;)��q�����nS���["�v��n�E�bS���..��s��<j`�:����S����I��&���;��-.�>l�� �V6%�G+���sX��0Ǌv�w���h^3��nV��˨	n�q�Ѻ7ĉ��[�[��i�?p�b�{�X���Y��M�m$�Ǜb��FJ�r�9u\r�W�[���ϛTi�+pj���@��A]oz��Y�|��V��3V[��r�a1��#.w_bnjȰ�Ʀe�{���l�f��f����`D"���9l@�V��B=|�<�������ԕo3y�iB��Ř6A�;�L`��ԯO=�)R��Ru$W�aJ��n�6��\ʗD��m(�v�ۃ�[�Ok���2AS�@�N����I�3	�3�bȴ���	�<�77�["q��ݷNP4E���y�\���O`��h,sx�(�m�$��m2�WҐiG:��i��K�M����#5���j�y�k;D��p�#��s��|�gY�<S@�&N���Mfvw
'��f��U# .�.�EQ�o��ӡB]�N�tE�h��	�j��ŗ�0fP��@U3D�u�6'��&t\&2�j����� 	@��6�\-SD;�A��A���nh"�>�����=��TG,Z��UM5EP�TLs.��6�5�+�w9�����ǧ�����SE�r3T�̓b��S30b��[gQr�4�ͪӮD�zzzzz>�6`�b��9cEA��2Q��[��U37OOOOOJ*��ض1̜.G#�ŴMS[b)�5LQ��UQUM�c�l�ƹr�r&�'��˕k�܂�ڪ9�\�b�9���p�F��<�.p+c8�xwc�5AQ�˓G,Z�;�STTF�4s��'��9�L�1X�3�9�(��T��S�4Q4E��[a�щ��F���#Zn����r�fٵˑLUG1�;�UDE��1ݫ�y����ݼ�ԤՃ����\�Kc��\��m����Ǚ�:�r����������j�۞��~�./��[)�7�]ykfT�3��_�OՌƶ/Uc����':*/Ý��eW�ȼ��=���(پs�c�����ͪ��%��!=���e�j�v���ޒ���`�O��s�[��y��w���\�{�xm��;~qm�o^��7�"]�g����~�k�wA�����X9銌�Uv{�so�^�[{)?�+�Y�C�C�,О�1岦�Ǖz����&���8���ȣׯբ�\���Lh;�Fi�{h�xf~�<Iۮ��c��=�ƃ;Xwdq7���ͳ����Th�p+^��.��c�y[��4a�0M�`w ���@�l{���k�]k<ְڱ��z0��m!�t�/7��7�t�O?��7�U�����S�X'z>�U��͘�oH4&p�E��ͪ�'���O�-��y�^�jz؝�#f]9��*s�`t�߶�3rO6��{I���ز���t���ʏ��)�)E���Z0�**�:mݘ5ee]Ļ�Q�r賲���v����V:t�k�1�ؚ�3T�NT�w�F���-��k{�8/�G���
ݳA�И�u����m�}=���.߸�M�M�\{HI>�̥�;ޘ��n��1�O޺{���Nvf>�PO~ǁ�8Yn@��r,Y1������@��r;Hͳ�~���ͼ{)z�~U�Ѻ�&��B=���9��nL]/ɿa�rwA���{����<���b �E�?S�l��z�ޝ�&w�X�d�����}K�Γ�.��"o3|�w�.;���>�+��<��,���O��g���_�k���qO>�Cn���_��	�7x�|3�a���u�돾���A�UP]sTb���v�~ܿc�z����~�Z.
��L
�'g$�S�Z�m'��W��k�ؔ��X��Ƿ�:��¹Ҏf��+\}��<��|}�r	���ȼc9�a�-S[$��݆+n�f��h�q�f�i�t�g8��z(iy3]9�VкU7���3��vއ���������g鼷B�N'DK1f���o;D[�}�p�:I)6E��ݡMVugA�8y�5C$����]`���P���4b��/֖Vpv���W�m�H��_%P����\]��Y�z��ز�*�nʐE���7��S�DnI��-��F�X7��ct�~c�k�����j�l��?toTNH��4*!dC���ݼ�>��ήu��p����7��}��q�����W�ؿ?/^�]=��՛v-;�>ں���o��p��;�W]k�5��%�8�\����U{&ؽj��U�_�=�D̙9^*>�����U|����B�bH�\ɼzn7-�;�m�b:`1����Nq^�}dGT����Z��X'���cg���@h�pUeYtG�6 ���|�g�ʛn��p�sk��j�<�<~����g{G��J�㤔�~��G��^S���Σ�Nێ�s��U�?S�,�,E�n�=��������b��]v��_}=�lJ+ڲ���)E�j��u�����[Y���_Z��_Z�S���a�ag�o�e�_a��	0CWw��
���E�V_j�H,�2�oqfu���Δ��1�yo6���z��'���_'�����Ĳxq��g4ǚZ ��I�b�Oc\Z��������6� '�h�Y�&ފfv͝��6������Ů{Y�\�@/����	ȳT;�Q|��k�=�2���ww�G
;7}���k�����>��{�c�bU=	�C�RA�<�5���}�,?$$m�]g�����������x�Y��,��7q�o���lSt��D
��ζj���n����D��ó8�s��e���fo=F�(���9�!�2t#u<靝���|�+_ǸC�������'��	�tI��^k�5۔o����i{��EP��I���A�l�i|:ٝ�s��x�?I*��n�s==C�ْ�{H�O5U������U��=�guu[Z:�螹�t��{��}=�7GI�<z6Ɩ��fp�`�|�l�&�y�0�1[��mwow׏�nz��x�5�n�_��}ڽϏ�����L���ݬ�C�ݣ���̏�7]2v�s�Oz����u�N�5ڏ�b
�~͙��iK{�hܱ������.vk�F��[�a4�#���/e��|�^�EiA:�r���H��*�*�w{ݡU��H*�1���M���Q�V���i=[�q����	яl���nG�P[HM�%ɬ�ß�F��;�$m*Jŧ��V\��ޡ(��3Cp!����鞏���i�7�6���K{ǫSF�G��m=��Ah~�"�Yn�d �+de���l�y��5�&��}�|&��'}�ɟ������N��yM`��'Kˍa��
�L��=[9�.�=�{gC�l#���`�M%�<X�l,�M}ޠ��Վ���w��ה�h*��{ެ�Qr��J*��ȁ�v��ܧ�4��̟������Gώ���5���k�{r�څ��-u�����E\���>����7�|]s�{�n�)���E[��ێF�ݜ�'��������v���Wu��*��o��>��5�ukt_��T53\lW�n���U�:��I;�ܧ��9�}�}[��ۿr�{[���w�mg��5?mrqB��;�ƶE�~���f��,��*�Գ�й�לf���1�2�6�iN�0�Nmu9����u�Up;ώk�"i��Aȕ�E���H��FFS/dR߫+.���Tu���i:��d\�-�����:%%�S�ƷT���|�c�u+�v�3�1܂�`!q=
TB��b�镄u+��2�PwwfiҶY�b7y�<��n�t�7�2v���5� �V\,Վd�Yߴ,%Z����=Nh���S{���߯�����ވC���ه��Á����J~Q��^��Â�nl�����T/�y�̂wN�9<��6��[�p7i�������1���}�>���<~�]�h��t��;>�e\M�2[n��T�����6L�E�>�k��g�ҡ������=����p�⽵~�ٵ���^5�|��e��\�NT:|��g��zr(�=rx�G7�l�]]f�8z���	�=�1��@B�>h�S�Ez�M����S�{}cfF�$�s5S�V���]�l�p�f�>�l5&o�_�|��~��Z�ڋV�4m��=x��4��,�$�1l�X�(^�jznt��o��8z��P�uFv/�k	���$��ǽ�iG���z���>�BT=��KT"^�[��1�7�	Ɓ��f
Sl�D��V��P�*��q�d�tg,�N\q}t���Y�����OB�Mbn�9+
�W�,��V��V����CJp�+�؋��s�g5���M��]k��w�Ij�.�y�~qw��twW������F�h��n/N�Kީ�Z�7��� ���eU��W��>�����5*�+�k��]iї@�	'p��1d����35ߋ�|mD��N��oq�O�ə��8���Э�d�up�oq�=衠����t�L�3w���L�R'���[�rI�0|:4��\2��F��㣍��9�Ot�'#ʉ��<��2|On����Fz�oH�dA��k]�34͈�<e�	{o��:��+��F�=NN���y3S���ќ�ε~�ϒ��}��7��*��U���7���S�dfOW.�z?���{lޚ{wo)��=8�tL`���׫J���\���+�W�����aޭtO�ʡ�-���w:��[��E���ݹ�GI�:�LoY��=�Ü����t|���/�����@�z��De��t���O�&��d�2�R��rE�[��9�"�E�F�pK����4H:�s��{+��\ǄZ1fvf�6_��}CS���^���N�����mvc���M][T�E�eʋ%w ���z0��y�$zג(S}	������yE��r�.�;(��<�en��8�t\9��)��f��ǂ�ս����/<��x񠧾�_�Q� f��̍��=�H�7�|��5�T׷����}
1N@�m#++��a7}�R��y����@
g�/T޼��Q �f=,le�)��j�n[��{հ5"�Uw����3y��o�S�@k����i_?;���X��z�^��ȏ���^+�:m��������&���u�w��:.���tƴ����޷�9���d�Q�-��Uu��'���o��U��V�_�����ٙ<v y���{�c*ռ�R߻��@�NBgr��s���ܷ�ģJ�7�)si.�gz���vfSBD}�:]^�Y�Q�|n�����������Zc#���x��������1̯C�:b�6��g
��E�W�ӻ�\�=v�:���mt�[ӭ�
���+e1���:d����r�Y:�j��M����<K]ٖ�vs�x�����!s�-a�y��"���g[��F����vSW�beof��`% i�\k���z�Z@�2�ۇ��ϗ��	3��}�w���V6��j��]i�p�Ž�s�۬�ױV� �{=�6�p����T�B�i�B��G�|�簵a���u�fy�`��˻������̛�}����v��˾(a������������eQ��ޮ��{�޼�3��9|�0_�Ȓ�{�&y��������f߰SP�>鞏��w5`�c�\hf,��=�t�	fO��P�S�L}~��i�'�ߥ�����%?r�槗m�R��~�=`�Ӱq��6�����6k��_����n��'��o>��:�\��(_����c l`v2�@}�b�eޕ�^�Gm9��t�}���zn�s!�k6A�Fz�� a�h���/y^�Q`=j�x�Sc��D��;{=W�����LN��^��b�f�A57��@�Hcܳ��n��=	�Z�Ҧ7/�Z��H�N��Bbҕ�a9����X�G�+E��Z�����;6D����f����ڒ�Ӊ'v�mƃ��[3U
�Wq܎���p��0E�������-�i�\kQ�S*���;�=Z�o
1�B���νi%I���n�RJ���Y^����JC�=^f�x����v���~>������	�73	�Ƕ�R�R.�ju������ۯ[F1�?jK��s����&�9�[&琉U�]uHk|�k�z	٩�5�k��?ݵ��M��=�;��`���������[>�C�_���03�qg��{.|����2��:�Y�����K'��M��0�h��uK�G�x=��������ts�����D�5�<~���*n���O�I�vHk��3=��ݣSݏW)�\͙�¾F�K�B 6�H�����c#,������q�9�b4,(��Sv���Nt94�u��5���J��t��~5���T���u��K���Y3w�ln��P^�����շƻ����:�߸�M���<��g���p�q�ԥ�WL��s�=�3�q9U9P�>}���}���x�=u��A���1�ڇ���Vz+� s� 
Q��o��[����׎�T<)ZaZ�À
k�K���:��i	|3;n��Rfȷ�
,��r�UmnX��i�C-�u�����U��tȝd�Yz`���
��Ⱦ�Z�d���`x�.��Ma��ֹ5��'u��� ������kB���I�U9�rs�JMԘ�����G�V�Ǝ��cF�!N���.��(�F`��׮���nci�P��b<��ە�A��u_#��JܩgzfT�IS;]<y���2(Y}cL'S�y����]m��s���ZDkb`r��e��a�oe��N\��r[�,o��̔��DN��ѵ��d�ٳF�Qb��C&mc;�a��vՇSC(�p嵮��>������|+]ݣ�F�|lo��sdDK�Y�롻uf�b�ħEg���7��aW�*F���T�]�Ď�s�y+q��f_X�0vM�CY{B�1�O����i��$a��q�h�5ǣ$*]��ЛM��u�D�:���'Vt�l�K�W7t���e��ͩR�p��n�Q66D^d]1#Q�hELGnl���N�.q�T@�8��$�Ѯ�{��4P�uؘ���uz믜J�v"�������@����H/��7�_U�驓����X���77D#ٙf��V65q�i)��F&;�d\�Q��ۅ��0�a��<��.:�ƹ�)��M� �\v�iV$Ӯ�����!J[�5�W�NՍ���@omTZ���S^r��Fe���YR�ȯ|׷~�d|8v���xp34G!Q��F�wó��ں6������]v��ʵڷ%���=��(�eLA��R���SJ�j��t�
l�ާ�����x6�E-�evsu�]��!�Z<Ji� џ�笁�\^��a)�ꕢ�����p��D��z�^}��A�d�Z����-VH�eGƖlS��u��G�+�Kn�e�Z9%,7l)]V�s�:q�������Y�t���*&�:�� g�����ky�o7j�͠*ga���#���.]�m����`����cvk&}��zՋ��/d��������m:��jr%�b�#�n]�N���_s�R���Hn.;æn���-:]"p����n�����K�@��q�����{�U���=cpʘ�+� ��VNP<��
Xy��U��M1^l�)�u�Y�Ł��\�9�2�V,�;E#���O*Y��2����ɕ�0���Lo�O��ˌ�ܡ�`y�l����}wC�>��X.�B������F)�Y�[A�gi�o7��C���Vs}.��qoV�A �r�3��E�������k([�i��1����&8�v������B�k
Q'^c�32�^;�b�s��;+���x+A����7�j�eH�����������{�����Ӎ�;λ�G;K���-'�J�|lL�}�εs;{v�Z'�M�C�N�b���3yq/1�疋�#�nX���7#sE弼y���F4t�H���`�	 �"2(`�"��2j����";D�,Gyǆ>q�����;��2V1�^����[m6.G=��p܎<�xt�===b��%�{��[�y���1�;��Z;w���W6�������3�9s�lm&���"6��5[cù��ڳn�����1��A��69��v��9�׍d�g�Ƨ'vE�Gy�\��;×s�i�q�q�w��zzp����3�lr�;�j�ہ�ˇ79�-kk�9ǵi�����nj71͸]���G1�w�6�q�gcˉ��TG�rLs��s.�8Vi�V����6	+�4�7,E�V5�����y����v9;��zF`�wnw[�Vع6"5i��j���9���Qk��*��+��Վp0L��x냰r�
^A�A��Ū��'y��^Gno7)�֚y��c\�-�c��r�Ӗh�gQ���h�EU�4DU0W9�Dr1DDZ��gn��UWm����@VL#w�h!��5��m���ܤ�<q��}�V�=�Y
�&�+m&�=�V�a&-9̲Hga����5�a������쟧�O�́���|N�����e&�8��haF!�M�3b�m�zJ2���5���*L42��K0F1ޖ5��h#��Hҋ�(;@q0ISi��m�By;5���s�1R�-���z㼕�%$r����L��>�����Uu�~F�x��L!��v��Ũ���ԡ�M�_2��>=kӾ�|�	� ,�Fb����}q6C����ް+�z~�-���"�4rT���@;�nu�z�9.�qE�Aiw���C�<�ʑu�ɦ,+����&�����λ�O�i���6m����롛2j���d;+�lo����傐C���  �z60Јt���➉��*�Q�7����H����xV�	�Ny�ڢ��P%����=Y�;Mf�=TlONh�����[����ݷk�/��}(�&<�dЋ�s*��%�䮑[Ji�1��9��W��_7���+�� Ls3�Æ/��<�>Λgn�J�-��<��I�p��x._r�5�:����n�#��b�<�8�V����W��k�<vڄsq�I�z;˻�zjt�����83u��/�����s���oȰnj�!�Ĝ��6����W������'�\�r�EZ�EV_�Z�h�x�s߸�8�Q���urJ�,M[\зC�GUѣZ�Ճ�jV2	�7ݍ���Y(8��?J�੫si��GT>�Cf�@���q�{O��67�k��H�L�ͮ��%Ck��T�~��q]�����<���R����,�'����� +�y���p(�Y�J�3�4>Z)���7L�>�ϟ���ܒk�xt����?)�^�*��2� -�hR"����&�LQj��H����a��v�Ti�W1Y=�.�ZP��݋��uxa�^)�j2-�gzD.����E�t����ѭ4���p؆;MU���Zf��{.�/fKT��uC#ؑ�=�\�P��m޸�0���EX���I,�����;�6�X}I��A���F���q�P���>�����c.��d���o����H�����"��ܝ4�(�T���@�RzByW��T�4�����a~�Y���:Pj�{'�έ��UXc=����;�|��{�YEw���9��N�W�Br}��ӎ)���OA��،��r�e�Wڅ,S9P�s��P���� �9�q��#6�=P����
�l:�wk��vw�>Im��gU�@�Q��T�
�{�������j����a,�[~�Z¼ں�}���}���Ľ�7����j�Y�ľ]ٕƢհw4]��=������,=�Uf���݉�p������CcZr<����Լ�˕���ޖDN��u%�5}v���gl=�N���s��Q+��l����RJ�H�V�v�IQ� G�C�c}��?��oR�<�􇌖j��Ɉ/��#�h��t�\�j)>��{iV닺�<GU!з+y��ع������#���{k�~���q���)�M�fWӬ[DgQ���\�`���۱G���tT^�OC7l��\��-Y��׷}�̓ _��><�L!�^H42�ǔ��
��y��ױN�z�v��~^�X*Ys�$��гt6������|DcH�L��K���^��*��?�Gb��]ٸ��t�.��L(���;)��]��|T�p����>�ٹUar��D��$��C�q��v�F0��Y"W�Q�i.~^"U߷:�E��~���C�Ei��$0���u�bt�a�|v�y�n��LB}oT�w9�T{�ݜl]�U)q�����m��� ����F�[o��B�^��NM��oc��8iH�X>��;��TQ�%����7�+'�� �mv��3�/h��o��x�Ƭ������P�~AXAj����c&�s�ΏG�5�8��K�|��%Wi�3��wy�W��l�^1ba��m.����FDJ��j{�kH�
�z��.��u	p�8�j�Q�_P�'� ���[N�Pr��4ѥ_�f�p�!��e5NIySC�|D֕A5��yf'�X�i<u�4A���	Mc�mM�H���p�P��Ͷ:�(�zf�qmtam�;��z�4t��⥨wp]*\�t��㌆D�}L`ag�\f�URj�wT�Y�˿�a�*p��l������i�N��gqi/<�\/fGC�9N��.9�0{��6;�erp���'{z�X��3
���ʌ�w�]LOi���p*j,�c[+�ɖ��{�=�<�3�!3T۸tj]�=w����M.[�r���4R'|`w�кF�4�c�{�c�(�M
���*�6�c���xw4����q�7>ﳲ�N�#���K�� t}�BtU���ȟ�e�����I��ce�D[��;�T��W�z��ֲ�UYQ
����Y�~J�b�]���C��ܸ�b*b�SqNq�TK�y7L{H��˘/WL��w8�2.sT�u�2񅂣6`WןB�K|5ܣ�By���� �k��瞀x=�A&缟��<���<[�
�ouZ"���g!�v.$[���_���3�����y9����]��Dk-�ۆ�;�2��JJ{���_�G7QR���Ҡg؊}�m��3aS�؝�.�^{לW9�"9q�,�Z�dK�b�o	�&4X��Lq���≮���֠�~y�����f��Nj$���x��9��[�bٴ7��{�n^�8:.���=n��I�	c�J�w�SzVun��jU�ͅx�=����X;�!��:4M�Ɏ�ۇ��v��t�|x�[0���K�h�K���K`(�X��LI��E<��b�5;��cO�Ʈk�IA�$�hz����DGwS�m�nj��٩N��6n�+/3��O]0ڛr7�$�f@�&��.�] �r�h0nB��C����k�J��F��[a�cyQw�a(�$�޻�U���Ħ�q~O�i�j������0nc>Z�5�|�n|/D�K��s9J�Z��ť�J���F����=��&�A���?�ƃ�������5�MdF�fHz���i���izʇ���T�21�=��.�44%3p�^Ƈ��Y�8գg��kΑq/�}�SB�"�Z��f����_D���y�	�_?)Eהr��H�%M���nCLv�*�^kp�V�1JXIG����=�%a������Veߡ�ov�*Pm��<��<����TK���Dx�����7�K�c�K������Y��MG��E��"O��n<��r(��+���ӻ)��Ls6?sG;��t�΋����J��b>�q�hY��R
w�B�>��5mN� ��fvΠ
�Q;�y�C&��ɷ�Y,�m�����N���@=4���W�����:�"���ǖY2?�	��p�&'1J��v�|�+-C���h�����U�f��^<�v��.��B^'.��w��v�X��.��/��
�=r�� �+a֚��d$����q�^]���J����!���jDv�¥	���k��95D`��)�| �yR�U{26����TtI�%�:���_�4	l@%9�~����/��.���G.�/sl�����Ӌʗ	P���ޗn�dށd�0����Ut������j���N2� ��q�u�Ի�� n������eӻF0�S4x�pQ�.4x�gi����E�k����)��4K4�}�;�9��k)��+��1��x\���j�;mB8��I���퉝{������Ӹ��/3�����5�������Ϥa=�=�0ڣ���-B����l�xTZ9���OVr�KT�=�.�R|�F����o�4K�k㻶�44y�{�qBT�T�dr�0D��v��B�Ӫ�ͺۋ����TJ�a��4'�͏E�N��?��h��.��a�m�UI��d�[����XaK<~��1k�8�QX��}�ƇYs:�n$hcZhGW�Us�����/�Y�,X4��1�}�v������:�5�a��`�"7$ux�N�L���:�S�G�v�R;9cy˾��lX�/A<Ј�a�6�0�:/^�!�^�'�����N���|�I�ܘ�R�����R�����S=��I���:���s8��W��NW�V�Z�_6V�.�n�
{� yO'H�ޟ,�tb���e�P�ԫ'n��R�Ʃk{*��wm#`V�ɷ�Z��j��-ՙՒ�ov�J
��5�k����[ <�Ġ�Kn)%uM;��Y�1u|����jR�P
�9�@�ܞ�z�[���xj[1H!�&���ϫ��d�(3����<L���SޛK�8�j���y�ّtSIO7��Q6�V,|���yq�M�ջ�P���A���YL#�u}"M���J{�iA��B�侽3����]����<j\�y���佑VOԄ�zɋa/�Wk��o(y���	e
��*���<�[a�㊭�lC��lׇ�s����C��|��WG�O�1����x�mq�^Ί����{(g���-R����NE�f��/�=�Ud"�԰|������iC�$�����/}*�mZxv��A�.�VK�^��b��Y̡���z�ޘH|a�&J���xH\�d���	urm%�"�*ǔB���ʥ���iө�NBy��_J�t�U�T�DSL��*&0ȅǚ�^���5;"�A7~j�����99{8�޴��f�T��9���T+q�?92�b����m��@]����r䷺�ۋ[a�l�^Ǟy��P��0�M�V���O�{��;!QXk�pQFM����AU��}r��&m��W2l�Cy���}{M��9����׳\<�b���Cޞ��y�w+�Z]�ռV����4�j�}��+62��^q9T��0�3n.|���+;C�Ð�;�)�鳖mG�T��ڢ=Y\���K)7����]f��0���&R�h!GҖS��
A���u�p� �A �;3.k{=������b9��f4���t��0*eyf�'����,����Ukt�Ωe����s�g�S$fD�\A0&:a�1�����H쮲޿��ZSѐN?S1��^�D�����mU2j�Q���$
��J�!c��M��S��bwS1:��=9gT��t�m�����Lq�3�UO����p	�)�$dDla|]����*�5A\����]���5�T�'�%��+�B���WI���;���x�5�3�2$�D_<�=T�~�(�8>����ͮ.�:���r�����!#���(ͳ��w�^���B=n�X���;�,֩�y�c	�(騵qx��ջR��/`��)�l� E����?��b�n�Ƽ%�L�Yެ�
we�0�-�*�G%g)u��4��.u*�Ƽ�%4W�HM��3�B�ٝ����jO�S��{���g�Q�.�������6�:��	P؟&�US�w�������]w.�����i��U���̱w����\֥��TB=������pCS$H9���]7�nմ�v��n�8�6�����ׅ�nɣ�U�����:�³s5��8>�ǻҮ�\-�s;�AR���}���ҳf'Q�5��<�u�k� ��lrg�l�%�[}ϖ����u��)Sn�\�S�̍��7Kn2�br�{)��f�}��9�]]��'X#��S,Xsr<��E0)�f�uq_.�_d���p����Y���Ko|(��}�D�k�!H�����O."�o]q'eS�O�Oc���5�����m�Ľ����,LfELVM�7��z9�>5><p���i�eҢ��E'���� ��-&33[\��J�}��O
��\
����֡*_�dK�U��v�K���B�_��mB�sj֓"�o{A.�Z��U���8�����T��`��^��w��|)L5"s[�㪛\��a���&:&���w��K��@f�*�&�)=���PŦz���3�Ż�5ob�q�Vդ�I���-W��A5Zċ���L0nc>�͆��Tw��޸����p�{���X���z���yS�5��,��3��z��1>�;ф|:���H�����أ��7��;��0P��85�������F�6.5�rBN�44R���b,40/VuE-��t�|$Ao���Y��� y|b{'�	C=�_b'=!��FCy�('~Po��F*�M$�*�v����#xBL�kV�GE�G���]`�03��a�8�-��0v��6ϲ�\�E�����F.�t;L6u�%�T��,�7��p��]Fa@g�8]gW@����2E����|:�E����f��^�sf4� >`�޽�}�d�N��_���˥��jR�J80,jN讟r�:$q����m�{�B�|G�X�k[_g��p��"�����3�8�����ӰA�d��n��r������N���+ޫ�mx
�HQ+��GlZ���nx���mr�12��+>6������č�=��,b�c8�g7;��0Mf'���|Wz�\̥Vm�MI�$�e��G_6`�=�Cy2d>v}�+�V9�~vE�u�~��A�v�Zn��=��N���N��-��%���`*����+�锱����k�P'��l�����j
��õ�=}�����"�)%�y(�-G�C�p��FI��P0SB�1����F��9+u}t
�x��G�����nc�(��;��$)���Fl�J����6�P%�Z[C����7�>L>8�ʏ��W�fmA� m����G��@�۬���u�q�i��ANl3��{f1���L�H�{`{D�mWҧ���R�;0�����;��=:�R)��ч��1˹õ��
���중�D�����y� 5M9�}=P��w���� X�ϣ�h��G-�+�%���ۃ7j�D!�X`�,��k��2�K�ծ\����@�Φ�v�h�У����'R��6�rlV��^$sj��\��m��:�%mp�HW�nZ�2����U���nS�]hSS�6�c�]{6hX��#c�{)�{�npF��ؖ'�4A]�҆K�\j�g$6�B>Վ^aV8�O�e �&V�c,�S���V�H����W��uc�u�`u�μ��{R���h�s���f!X7�32ΐ����L'�7{������o}!m[�.���쥻��E����7*r�m
�x�����)>��S��u��Sky�3$]%�*��	�16^��������˻�#6�KqIM`,���T����ˡ�͸�X�XhKC���ٚ��u�W{a�ৱ���r7���R�$�Ew`�ԝ�1N}Qt�6�=�8��t��(��5��)Y�S5�䱚��*��^2���d�h�+l ��{}�c�H�#�L�j���OdϱZ��>z���v��ݷL�3+�5��������m�����l�
z��>W�u��Q���;vv���$���}��0J���d(\[G��^�EQ�&ֲ:��YK���]�R��fv��L(w/u]wP�s;vv���[RM"A�;`1B���b����rS��
�]��e���̬�81��;�'R­i��3�j����ڐP,m�1�x��������j,&�&f(h�&\L�Ò�bh5�e��o1���X3v�����	�
�1�i��I]#{������ �
'b��c�)0p<���Z�ZB�k%��"�dZ6QJ����&�`�����g��L7wb�v6��գ�c�]�+x0t��Z�'kw:�����!�c��u��8u�$�ܝ�|h0��n;�)�D��"�)����s;1+�R���v��<�`�ˢ�Ab�+���wfvM��*�*�ɺ�:������Y���h�������/g��p�ҫeA�{�%�D�cޢ��9�V+�-=ҴJ��U/�Z�R2!;?��Ah�Z��ܳ}per�+y�/%I՝o�Q�ޮ���Sf����^�gz�;K'=��B�Ô��:���ݔ�:��+��l�S_����.7-|9ͣ���+�����V�]ݘ	��k�@�;R]��\���>z/w�R]���U��p���������H��9�{x�Z�s%vjrlN���z��:uH��ϭG��4��u���q%7c0��3/-�d� �yB��jɦ�Xݰ�ݠ�%��Vk7��ϭA]F�W}�Jܜ�ާ�hv��L��.f��r�\��e��.�GY}6����|Ԭ��ڼn���|�嗯2W-�J��8r�5�d���.!WJ���o�Hd�X�|@�s��Vw�k;���WJ�e�PgL�آ�^=�X����o
m�uGK�B��¬2��+4�I�$	���&�ZE�F��T�X��T�=F՝RQT�kUTų�**����Tm�
ѩ������|����[6�U;`�
��+�ƙ�b��ڭ�f��mS�M�cI��==<<=}L�JtrLE�`�%�7��Uv1�հj(��3\ƒ*���.AEr4�������MZ44h֋kZ��(�֚��α2�:�5�{�\�(��zzxzxzǻ4�4F��ء�g2�cg����ͨ�G$�TA3p�k����b(���\�.E3kU�M��m�f�5�i#`��N����M�ű�f��[i�ֶg���M�n�����r��K`��U����m�Z�E7"ۗq��*�b4�
�d��5�����[F�5h��h�ZS�e�ۄ'*�Q$PLs���-���8Mj`ӬI��qI4�:3e�����6̓�3�����DD�!F�  �1%�K���¹���Zf��N��y&��AC%�*5��]A��YYo��Ʈ�eR�A����+,��4�dX5l�T�,�Q�_E�>�EG���7�`�`����R�=G��1ᣝ[�N?��ȋ#$�L����1˳c�����l,+�aMky�ޕ;uW7�{�b��3��	������5.;PǤ�:yP�.gS��F�1����_�p�z��ǠD��f�N:�{o���Q�D�}�ZG/�ؽ���Ρ��yCYYIz�f~�c*ؙ���[�D{"+P�ba���K}@(TC�A��c�!q�VI8zCݯ���w5�{���>K��{پ�>�z�K	��`�g�Bb�-	����ꗁ:�2Ȅ��qe�{��x�U��6N�^>м�yMCqr��Bf��c��f��WN���'���oɢ��<�X�p�@���MFDgћ�g�W	U�Y�ܑ����N�He��K�k#Tۻ��f���E'I2E�a#EW,�ӋқT���],T9��.b����-|Ѓ(z��'��'k����9�=�i��b�F���{4(�^�"a����o�b]�{���(�G4qǚ��N{�u��sL@�4�wu���t`�5���چ/!u�6���:hO��P�ZLZ�X��I�ӊ��*��y�h��$o��k5Ɯ�}
���8�����p�cMa|�`A��x��kM��;�hĻ)��+�FrŎ��.�MJ`L�n�t�� �x�b����p�=b��S���[��
�3�1� n=�K�R�y�b[Ê���q�c=�Nѷ�
�9������}y�|�|�� �	b "Tx>�pR�]�j���|I��/^�^P����ߵ��SK�H�*_��	��� ����E;�ϲ��[Vu�U���m�;��ˠ8����`eȹ�S�)���s")�r�(�2!q�6{�,�U>���ͽ�2�mY�]�3!Hy�+��M�b��S#��TX�P�Ĉ\%��ϑ\�����9�Vt?k���Cb^��y��=����<�9j���d�Y��%l=3�k̵ι9�Y�z�]�dǷs7˩�������1	4[&T�7�wg��R�7}�c��߹�>�g��wP~��-�k���˄5���NA}* ߋ ��Z���^����P�>?H�IX:��xtS_U��J��g:��E�5T��Lc9r����1�
_�"~��̠.h�.�L7,��7\'k���q�\��M��Z�f5��Ij,L1��ͥ����Bvp�=0�l��������۪�ɛ����Θ�����g� �Y�ql�U�f5.ϜIZ�_D}�<��U?x��S�)ff�S��'g�
���V'`���A�c�>Pe�0,aSl�t��B!�!�߷��x��u{7�Y�Q��fH���O�lU֮++��Pv�$�n>C�\M"����2��*y�{9�z�)�y��{)�$��w5�9k9�]��:�y���WN�:����f)�|g6殖����u���b�s�V
1�,>T�:�N#@��Ka�l��>��	%"!h9��������������~I�uC��Dg|���S-`��l[^l0�"!�4$I~���:�����6uO���'<���U.���91�9����~0:��BѮW�����&z��Z �2���u�NN�6�X.�I~�=<3�j�};e�U��b�0ŝ��O���s^YK�C�U}{Úk���r��GEıʾ���K2��-���ZĹ�s2z�rV�z����SS1�����Q2;I�wMנ��<��n��+QS79�"��=�m_s%�o,A�k�#���G+h�U�u��H��1)�	`��n��[q�A��M�+2-�	7>�2<�)��3^m���\c��3�GMK��� q�o�B��\\1�%;'���_[\�#�=lu����z��`����*�	�O��&�����O;k��1��P�7��b�Q*�;�w�t[��C�-.�����W�H<����5@y4��4Q\��L2%.:� ��*-l�m���I�V�����N��Q_{���:c�Gi�Gh8�(h5�p\�<!�O�����1�]TEnH>
��{���5��e�� qU�omKtw�{}��z�u�r�W���̥^(�5ʚ{A�z�e�Q3���-Gz��=����oL�T5[�9-N�(�>�:�q��R���睤�m$%����"��\�]7�i3>�n���H�D	��o��p���������<��}�M[iJy���Z-�O��	�֯FKσ�0����h���r�xHn��Jee���~��
	�Ƭή�ˑ������=e;쬆����y��Z�Q|�r%��]͂���&爡~"d&
l
A���c�:G�qcأ�y;�24HS4�+�B�g��1�G��vp��_R�rA��2c�<pJ���]��Hv�{)�ls�-���
�:����qs����6E��ɘ'U�0g���3��?V?�f]��i��J2�1*6j�:����|�p�K_��g>޳!I��t�3?%��	�+ SLh����76	m�˪v��Q��W�à�
^�*���<O��̞������նE=�D����SČ��u3���[r>�Kwz(�b�k��H��
���MI�bIm�rݝj�S���n�b�H�Wt�j[�1�؍�i���f�1H&F�����Q�T>���`�cEg)��"���s׵��H�
o&!eGUV{uՒ�.�a�XPb��]�
*]��82��y��)EŇ2������Ǯ�ƌN�e�I_��n�Y(�x]��ŪLެ`��n+ɺR�����h8�Ɗ�/�ϰ��f��sNS��hv�o��lV��� r��l�Qw�vu����&�����I�2Ɣ�1.k���ĻnW9K�b�u�E�p����m� ?	(�nw��4)Y+_w����[�\E����<a{����-��N�sr����\�͚�g��\�R���7�r��=�r\/��M�G �n���=sX%xf�2f�50�����n�e����d�%�-@��ag�e�b�c��^���q%P:+?k�]2��c�ԘkJ9���<����9"s����cg�A�ܨ�<���W�>Q���K(�%$vDF����QC3(�b����B��X:���=����8Ȭ�L6��y�:͏Eo���p�^�0�3pv �ǳr�;Uٙ۾C�/%\���aS�q�ƥ���<���\��B2)�^�STĈ����m�.�Ӝڷ�)�@�^$<D���Ntx�=k�#�������{!�
�s��'��O6�ț�9K��|FӞ�HP��^S�)(�@�G�F~��m@<}ْNR�|����]�<�n�O���xq#�B;\��T�$�3�sƂ1F9PJ[�j9��zt�ݗ
aN�O�{�3�M۷F۹ψlf^U�_����Bfǭ"1���vtb����:��"��>.����(i���'�]jn�"1l��wb����<����q���WL�}sLY}�ʩ:Z�ĵ�U��+q,�'U�v}�ZW�Tׇ���P�5��Fwb�ښR�e7ŋI�ɛs9dO��Bu�{�k�����
VL��gw�����C���x{��{�³���$��ϧ��ץ�[P���ٝUz�C�B��:c7�	9��%3"}��j3�� ~sq�n�z~^��Ǜ����7.���Xb��Lc��U�W-�ݔ+^���!���]��~�(�̕E<�>�:TTj_3	W/r�X[�bk��i���՗�y�h!Ng�SNsnEbF�\]�[PE�Gx�?n���]�
��`}L��=�3wf���T^:Z���ߨ�s/��|�����ګ��=�ke�X��)�#$HH�� ����k�]��L�1��S�yڄC�vC4��(����X��J�^��%l��8���	�~�E)軳���:ծ��nO^�^E����SԦ)��Jdp���J�!G4;������}Z�*�KǛ��#O�1	�f-��YEΧ�:���N,VZ�ai,��:E�.#ZB]����|�J��W"�L��>�1�#��w/_�s�O��0j�U){�g��uԠ�����q�&}E���n�ۏ�{MDƦH:�@� �A0F����o/]E��׏ٿW��[履^kՈ�Z'RvyU��"]hޖ�v�����h��ĸ�XyU;���nIK3KPda�O��qm;�1��Nsh��	���k��Z��z�uOo��{|X�w
�|��z�O�7r�G[�zy^�s�qcv�!���C^mb�G��
a���\��ҿ��@ \������}�>�^��ʔ/��*2)dsE��ml�3�,���P�	�B���H����+qtx{�γ H�UBmY��XŪ�
�Nvi�'��y��y����)���ʀ���>� Ļ����n�t���7y�WwT}��"�*;;�Zh8�t�~P3�W�	�
�M^nZB�tK>����Aሌ�H9s}�����t���4�.���4�x@#og��>y܆�D�'�M�d�c�<!�T�젱�*���@$^�+˶ab����b�S�G>�J�~ł�ݻ�l�0�
�vk;�{�Qz|��/����v<#{�bA{�U�~a�Pr�+�c#���.��4��W��H4=ɧ�;^n���VB�쀩��b��X��ZEP�Q
CT�lٴ�lЄu�=�������))�]>:��7��3����\a���4˯c{J��Y�j!���*r�YJR�g���Q���{l��n�{{����A�{3� �fSJe�?Sm�̬a@�����x"�-�u@�6�޽�<+�(�	��j���by�I����yq�Sſt���v����aϱV���l`���l���H���)'.�^�z���V�iv��  {�h�&�2�ޥ��
7c�4�G�T�>�
���,��"nhFF�M����p�I3B]�/�F*�B�7��u��q�{O�g
���v:V�w�j�&c��ߍ��>O/_�S�BH�B>`���shę���Ze��1Ŵ�D[O��v֯J���l�-!�M�peAN|�)?7(y��j�U��1����Ǜ��^6'����
�W�=s1�MK�����k���|;�
�]�F���cș�{qv�d�����,s�]����t�}�	+Ue.+�4�<*~I|7�[cd�|⫥%�Y��"����~�ml�*a����o�����2;MI	k��yɐ[c����J�`;�64U5T���Zg�J���/j�]�8t2�k��5<굫�FK���ᝌ�`3A��^t8����jS��x��	圬�[	݋�~ϷxZ`F�5�T�:l�]�D$������C�-�iG��"�,�my���?F���` �>J��4GTլ^��Ŧ싷�f���y����je�d�<{��X������ٰώ�e�m"��8M{����ٍ�y����M�	z�rƥ-$���PpOt�XƳ'�Ϊo�V�	e-B~���/�i����G�'4>�F�ݦ���T�yRXˁ)_�����L\��S]%���l�A���hcVJ�qj�����9%���E<�u���u��PXqyY⒋�=Y�����W{m7�}O( ���k�wc.v��殡�.a]�m�Y��F^��V�dJ�?By��
H$R0�>�}���H��X���}���|}�����ʠùx�}��l���^��,�C�*S6����f������'�ɞ7H��ȯ	��zk�V�o\�jp$�	��M�Ht4ĭ{Ѓ&��ɳ@K*�o�mk^��x7��3���dښ�{|��w����2��wkN_V#b�:$��1I�>j�OE��h[r�LBYX׌���s�;����F�<-��Uf�.���ʒ�s�v�e�#:�S�����Ԣ�ⷧ�.j^^fj̺7T��)
i�)U�Ʈ��x�Ϯ(;�0r�=~��XP� �v��y����1w5.�R��{ة���ж�~�R<�9CoƲ������z
��W��W�-��&��+sN�@2�ˍ��H��ơ�s�Z�<NĮKt߾�]�j�����ױI�\���屳iR��fw�;qp������[/��z9r�Sߒ2Yn�,g�|״���崁ԑ�q��3.k�{��Q�'ѱ��/<位��w�h�I�������Vl�.�L�6�K�UK�������o���0�NDF�P>��J=ҟ ��C���9#C���
h�z�����Z�w7^Qo��v�v�r�����:uFI��*�F�G0���76	�VRu��X��AD��rP'GJ绸�<�Cf���%M�͜P-�>�y�j`�����ے����㔫^�,��R�3�^>�����H�� O>���;�6��Ԅo�N�c{��h/��74yݛ����ؠ�V���N�,�Q�ybC�������w6�$�m3�S�B�&53	o� �<�2#bک���&��lyOx��	Ȼ;ؙ��g*���L�Y�l)\��M	���N��N���"7I����MU��"2ު<�D�c�b�G��Șh��I�pN����J�vyͻ�mQw3tos��t`W��WI�$d\.}��)��#�ݮ����tx}�ޜISvS���5��q������i����ER����Ґ.)��ĩc��A�<Ҋ.���ɠ�\�uZ�sǻ�Э^�XSQܗ��uB<�r@+־��R�W���\h�Eb�sPvN������f���ަ�u�f�(8Ԋ�*����nXcK.�~����BW��"׉�}ޅ�j,秛��?��5��,�Л�9�\�S�M��/U��>��U�Rg�����X��j	kq��+f��u^-u!���A�3�۱B.��:>c�\�S�F�i����4Beb߾�>�{h��Ao�s�nT�d�gh�|0f�i�y��eՑ
����Īe�g�'
�j��'P��������]�LCr���}�[�ST+w3�$����O��3Cv�N��VGV�Ia�Q�v5���"�WuL	\*�ަ��aO�lf�TpL�Q�����ǎH9���й�^��R��˲��S����2�ˍ���e0&���܇������d�?'[x�ƣ�ZT�^�����x��7r�8qXde�`}��wl�0���dF!����Y69ժ�`�M�X;�J�2^�p;u�MK���)i��sn��;X�]\��H�_T�/�	��/�d�f�#���+�l�����򺆑	&`��Y��"�W^V��u��+\�ʨ��@v^A��K��gtRh���V�];X�b3J݇[g�V-߰<]��&����:v.~�a;\��Qv]&��=�^�X�U��VV��Sx���Ӹ��R�;���lm��jk��lf8����j���4�����Kr%Sv�ۉ�_V���q�D�ru�uMK}ٸ:�9f=IB��������%�[�f��C��αCmt��CLN[�a��M�\���#�}��_oݻ���V���<xsw{�8�go`��X��b�j����a�v�r�c��BS���`x��]ю�+N�2��	ǩ��\��X/�K�Tj��4�P�4�����\�h���Y�8|���tu�Z=(�FĻ`|�+�4p\��T�[�6m�Ȁl5���P�*,"#�'ak0��x���7�����ʙ}1}ּ�����X��^�xp��[҂ű�E�<��F l�ԥ�ٵ�+��I�i��t���69Nv�9��t[F�S�����Bx�YF�s[��o'l��$L�'2�6�b7&j��	���=b�2F~Z�P��x;X���'�T�ɩ�C�i�2�Mu��_(S<����Wn�6�[�@v.�pFE�m+Ͳo�r�9J-�BE�����G(i6�e0YgN<�k:
<�<9��Io-G4�Y��踳Һ�l}J�]oG��+����0��ùܥ��<���n��XQ��)f��z�p��e�����H"b��k6=�r�*펭՜:=�2�&PRS��SY3+V��C�`��ز#���N�+�3s3; =���4ԭ�logT}�\��U:�s�J�f�Ꝅ�4 7�z�Waɠ�meH�7z��Z��t��=�w�R�\��	�RK��2Y����Bs5�GR*V����Z����X#����-,5z'��"h��TӕمVO��(n��-���R0�O1���;�0��/����kKR=������.MJǋ���š�ժ��bl|����#��f=s���6h��u�����yX�����G��h�T�F+�h��`�k��R��i���$f�{��<9�ք�Qky�S�1Q�
k��g1rѣQEE���U��1:�zt�<=<=.k:6ڣA�{�% ��l&�"t:�M4UEIPl�5��'!Ѣ����j�����p��Yւ�ѡ"�b���E�N�u��Ѣ�Z���0rSzt�����y�G"*
]:�AFڀ�DIV�K��vE5��DAI�4V�ӧ�����ME4�Dm�mT�Aj�t�v�RPybJ8l�ATm����Ah���m�X1��E-�ۜ5\�yh��l��6��s+@U	m��E�A[m&�ѩ�AF$����)(��Wc:&��Tۆ���à�wn�+�h�b�m�kmf��ֶ+i�Hh�%Sm܎l�UE��4�E��m�u�rkF$u���Z�N��8�x�y�E�c��TjmUSc����9ȃlV�F$�b�*I�ۜ�3��xG+�&�Ţ ֪-h/�{��=?c�*	�f�+\z��Ǿ*���up27"��Â��g�;�.�c+�.C�^�g�4y������!'|�__?^}w����Q�+�Ҁ`�����0��7u7�-��K����%�@{��i��LS��2��n��c��PmR�
v�N��Ӛ��0��/��q^U�ô%G��08�*�-K�R*�φ�8�Jy�%���Y��Ƴ^O���\ξ�hg%E3}��XA%���K_�D�$�_��ƅU)q�%�#��r���kƹn��=yP��{zq�Aa�Z�gM�:�(`���覫��^��e��JxS�����]�b}]k��ޱ����ǥ��TVD�SkP�3�����H)@c�h�#}�U��g��scu����ܵ�3L�9���5s\Y1�o^&��^�����D1΀ͥ���:_6]�����q�u�}{��\#��b�F�(A�V�E�rU�O���~���ާ7,����)����5pT��^u�Ȫ[�\G�D���$Nd���v��׻�s�r7�D�r�|���E�K�oz���>���wL-\��>���|�3=a����V���/C��2�,����/5�`m��;8�3����bAH�]"%�#��r@+ܬ?��#\ki��l�w|�����+���2���:��ή:��A�ɱ/*�^`uo�iV�:hYT_+�纟[K��i�"oll�R�� .�ʦ@����%Ck�L2l��.흴4t7G���7n�`)��c���ꕂ�64f;���Y��"���1�����bbbDT�ןo��ןc���/�~�N3��C
���r'�cH���>���{��<�_�E-�;��t�3�ns˸�'��.������fX�;j!M�K����1zk+%���w"�!��/0ҵ�Y~N�CdhhGh�%��	�Lw�d\��6�^Y��(���+���ԫ1�4V$r��J�}�r�T�g�W۱�s�T��tC4',�U)���U�m�n.\PN_)љ���;�����c7Zjt���F���o��/�H~�(��4���8�s��T�/ֻ�Q[	�)����@0�?-�믒� ����������ǽq!��^q����!��r�5��ޑ	jW%ۗ��򁺸s�,��V-��@+�AM���M�����������V�or��ܝjk�f,�����{��F(�ҵ�\�|���
�	�ν�|�L����j�[����֬��֨�4��ΰ��%��j�aމ��$\;a�s���cΞ�m�u���!I��U(����U�h:��Ss|��z~�)���鯹3�yf�*��!vl��©����pִ#�Q!%w�O7_�JJ�S"��U��)��-|�t�u-�v6J=�05Z%%�E��s"��.ft�݉N����䫕]�.��K)���f`�ldO��VI���d[Y�U��h����+�����V#�
?���s���~D��Ĉ�"��  yx��
�wI��c8����>NDA:9x��=,�my����X`ksQ�'@v��w,!Jjo"����׭�6n���	�d�q�P
	�=`ǲ=A`�3�;ｲ,��hmԝ���]L���v��}���ԌE'��ɘK�8��U�g�ܪj0��H4D�:J����c�S4�p�l�aA��#�����/��K��-�P����Z,;�v��6��X].N�Q�ܚ����0��ͮ�D��ղ�$b�ɘ�oV�_5�>h�nǞ�&j���ё�bXU��K�ૡ�Xf�t@�A�M(�M���g�-�k�8���hx1�gsW\�=��5D<2 �[�5�����2��h����٣����<�1E'ᝡY�8��jj�Uxy�ж��T{��V�cMn
�>�Ǻ�0tlH1~�dPO���M�lx�P��f�F�������z/ܗ+��&�kI7=/u�_�X+:^�?�y��\�����X��΄�o�{T3���Y9����Q�)P%�,��nC�zFK�88:�{�B�s�mדlҫ�@����<u�3��T�Лy-V�=����}o�e57�+�'%f�(�K*����Q�%�Зj��ʋgה�����s���zp��'��kw3M�r�˜7�a�W[�s��ߛ�������� ���Ā�� �}}��~;Q��)@mo�<74�x��>�T�nQu��{���m��X7�09��Xc+���	=F�����0�:��)xE�^K�C�;T�l��\���2Ynx��h��J�^D(3���N�W�t�[���ZH��G��"�a{��k���U�C�4,�)���hO^Y��z�����s��ӻ'�2v���k�jXH����T��-�u�Ǟx֫��q6=�a�j���?R����G�a}߲�&h{D Y���]�k�z|jWb�/�*�-��)�l����2 �����]/�dfzf���,L5C�R���;@���+�c'b�6�
�!�@c��Y�nd���8�:0��&Y�4����^J�/ԗ+�*���}��O���v�e�S�S0��^�?�fD�O�#�B�G���+'��?w����bk�\����p�6�yȺr~֪B�Bڅ�|�U����PC*�Kf�O�!��"p�&�4׸{;��Y6�9P���2R*�E���Q��,1(X��2�FR���M76���y��8H��5�ܤ���k';����T�	�&TL=J�mZE>���M�r��/�,�5��J�0~����N�;IH���u�L�yè�lll#���s�N�ʲ,X�q}���l����]�Ҵ���3;���	�[����~����~C�@���
�oxy�� <Q؃)о®�K�oe
ҰR�}��sm?jZ5���es��ژ�?���/6_�Į@��Z��o�u���x��킫u�������v]^h��i��j�)�GP�^��	��C�K�����֯���GJ����c�t>I=�X����o��U}�Rg�p9s���u���s���erY�W	\�ݠ���4u�/~鄝[(�\��O�O�Hݍ�js".3",&;s�\��rT��q��9H��+�\{�J�-��<�ߌ�/=\EjS��29�<�N�/�'M+Rӷ/ݫ{�f�_,���R��exu�\_��c��y�������>���̺wJ$�]�D�&?����f�^OyE��!��Z\%����OG�
�?9;گha~G�5s�Q<��ܢ�>����Tr�����=��7��kDji
dtoD�t��v��Yq��*4:�w:1Cq ʤެ<�#��AˊY֟ߛCC���~"�yP7`鿏yQPA�Zd��������"N0"�#q-�w���W�1������\ѯF�KP1bc���*�:�����ُP����nVf��ک'�WgI\����-�w� 6_N�투c��ۈ��e�X:j��uvfM�f�3�l��+y���ۏh�ܱ�č�5����;�-���0j�$��֧��8,����s���|�|{��(?�T�A!� `��������J���y�����	v/�/>7ǅ��4��g��_@?@�g�u�}ז=�a�+j�F��DV-���;��ĳ㪈��lR"}*p��[�ֽ�>±�k-A���fz����j&����Z�qk���p�`@���6���g[(��U����[�<k�8�>�ڦ���@��h���UѼ�q[\=�؀�$NP�X�mܽ8�uC��
$삳���԰J�x�=-]ER��×|�W4�eU6���Ri�6�R����=ϲ�.r�����#���T�H{��y��F��(l����O�H=*���K'��4��ا�U�
�����Ky9˦u�؜=��K}~��J��,�<�x��mq�%�x���p%Tȹ�SmԳ+M0�7��#P�SYkoub�����k��
-�>p�kϭ�h8M��Hȋ��0Ja�}ݑ݅B٤��]�V6i�����^���,4>�
����1�tЖ#���~0~�h/p-�1�O��ҟX�f6���:���rq^T��g��tObf�z
-	�G�EZm����|矦��c��$i~:QR1��
V�E7���[��Y>~��#����=�v��*]:R�gtPND�Y�-.7�Ub��y��uȞ���:/�k������.��֫x�"�_w\����µ�;lϷ&�+v<�r!u�)�\��^̖Α��߯���_���Z�;� �P�D��

�҂ �;w��s>�k�ܡ�f�$G���On��^Ϻ.�j�+,�>�������C����c)�����C��w�����wTƽ�%��۔�㍅�sr�P�&���h�Tt?j�n��=����(���R��`�ӱ�h���O ]%�*�y����l��c5͏�,�Ұ*�}��� ��D
'r�\{�J-az�='��]C���=o��g�s�l�R������5h�5��ױ[Zw��^�t"�LB.Ϣ���nz��U��G��Qs#[�؊z�OuusV��=)u�P����P0F�B8�A9�0�`�TP݆m�]{4�ʧʇ�n�i[��a�nn[���6r�T�AP�].HS�KL���mA���S�JuO%��̬��7�=��-zRg��32��'w������ �f�5[Hy�:~iwա�N�lS��0��Q΢蓞t1����{��q2-¸Ī�"��%�8O*�w\���F�踈��y�DGg����΄�W^�_p�y;"�P�<���kLJ��t1��Y6߂YTի� �����/8C���V<���6�.�^��Ű-�OB"�O�0e�e�X��#э��Y�e5 ��f��@���ɠ�G��9\�3�'��b���O%-�WW�魼l_�:�>�μ�����d��v�I�N�3_�}_W��XJ�@
R�B*�x��g��6���R���xi��2#Q�Hڈt���g(ƣة��\ןK�^��]p��n_V�2�i>~�E���-��v_5�]hq�)�ڽ)K������W"���}��Ϊ��Xj'�x��ۼ���3Ե����_Z�a��''%��c�t���h��2}���鶪�^xz2\�����+�
2k�e�*<��JGs�Khu�VS��z�2Xk޿����:z��h�G�'�?3��H���7&%�=�8Եw+�`�Q�r�`��g�s���
I��xn��@�*��-n,�
��Ne{��ǽ-���*�|���M*��,��y](����"�=���/RO��jH�b'�!r~[��k���5?9���yt�c�K�GFF�U5ܿEw}���{������j�TW�,(0��L����o�C��ŧ���QW!1~���Q�/l᪫G\^q�l�Αg_=�,4��0?	�
��D�G�}!v/#��-����ȷ�VO_/t�|���֡��S�0Xa���&�yw��"]トb���}K��ߵ�!�H� �$Э�x�nJP��Юtp�)��L���f�4=*=�ٞ�/D3e�c��&�!b� ��F����<g+��G�bp㺗I"��<�M�&c��T�o�j�и{�p;�@6���Ҽv����x�+r$@�ZI!�o�  �@����� y�{� )Op��]\V
F_��m��ln�د7���{.��5��r��E�'�yw�&\3ͼ"YG	�X�!���ȉ�%������0?��fE;Hݎ,�PY���wrV[���c�k�*���\:v~��~��NMyY.�yTu���a�.�Uγ=v����<����N���xg�9gDnͩ:v"]�~�IO�m+�%����`���U}p2W�}P�B�;T�բ/�[̦�У��9�0a��d:����`��[~�Zm�#���0�Q�_HjR���ܥ"�q�|�'�^�ެ��Rܠİ�Ƶ�Ys�yO�1-���1������C�4,�}fp�ۏ&�? ]�Φ��3��(kZO}{:|j�3a9��ϫ���5R�~\jJ��Bu��7�)��ׯy��bj�9H!D˧�(!���a�n���3):�6��E΅���gC6f�[��6�-���;�s�b_Uaѐ�g�L������b�R3�Y��${�)��9�\�KUṹ�"F��Npx����8��|7��D�[F��	QǪ`&��1�{Ȫ���2�_r�h@�W�_���xmB�s��\��¡]հV�w�n�E,�|W��{�>��!o�����զ�gZ���hu�4�e*hUĴv	�mħ��͍9�S� ����!\�
�i�v뺺�@"��6�[��b*��%{c�����ӟ^��|^~_�$J,H%A���=�����<�mޙs�kqfڎ����{�z%�r2V�q�&壭����k�M����o]{L�ϖ�XOm!k��0�zy=���
��ИX� 될h�S0Q<��~�p.(�s\�v���m�t���*)��=I�\NX;|��ȡ��t����ɜg/`��?(S�zs'��;o6�����K�p;�G�>5�u̨wZ���f�&Dw�x��=^H��f_cĸ��f߂��w.�$L�]�"e�5_J<��ۤ�Z��0���ag%ųa*�M�D�9�|�;���\����V�%�i�:O����%\���YSPf�b#f��G�໌�Zݤ�su7�� w��	;��6;�e}ɈKWh���r<B9�&��w>Á��-��f��i{��V�~���#[��r�>��	�5V;���Ӱ��q��������(zw��6=p���f���٦��U�cg	�iH,�+�X���EW��Q	�K���**�>^��RѓD𝵬�8T�i���nu�=ܥ���j�����*͋�U�2��`}� �c�K�=}����՚�DR.l�A�Ǣ��.���Mi��nv�J����sh��2���(ړ�wp�ӓ�\�ț�Ż�$���8,2}.���c�Ks��2�m�fֻao ���fJ
�b��6���ack{�v�h�ᬫkU�e�1
���ο����q7�v,�E9��Ŧ��]Jb��8X� �鱷s��"��/S��γ�ۡ�ޓ�)�nNQ���8�{�ۆYN��r&>�����r�
${�Q�����f�v\�W%g-}N�@P&"J�h���{̡N�W�8���b�B�E����'7mu��4);z���Z�X�R��f$��vP+0Ve��n�A��{�.�YO�Y+���Ԫ�_�H��9�[7nA�"�lot����ea�쭾�C�[��MBY��.ѫ�q$�	��Nv`b�H�!��N�zԵ��9��1a	��ێ�J�}��jN�ՊRᎌ�̊�����7E��Z���6������"�p��4���u[� ���N�뎲��*�C�cB�W�H��i���&üٳd�u���<�=��v>"��`{�>[j��ި��;�����by7�E���h␛@mn�{�ΰsj��r��&;�QUK]��/�����iU��gI��r�͙��ul ?)�5%Ԁ�.���ͬL<��6�PV�W"���a�k�ۮ�
԰�yu�d��ꙷ,�zq�� �a{���f_ej�N4��	�P���P9�uѣq)��.�}����bP��k�U�M��Oܻi�c���f��۩l��������xa��6����}�ӝRhۡh��g�-��A�}?8�6��N������R��{�v�A�Z��m��N�Q{�v�bgRn��i3Y�=��Kڲ���#{����3X�ר�w\��;�s��B�Z�;]{���  ��aU�,�}r�Q�C�-�ӧ�|7) ���p�}BgXƒW�M�o\չ��Z�_w>�㢞�Q�Ӣ� �@��u��v�q����U\�p��X& �5�Q��w�5MïX�%���9�`D;�#YE�;��xw�P���M����"B�QZ�b���v�^�tR���R�X�ԭ�Nu�yoU.AS��q�6�!��㴜�	�uOI�uːe���������A�H�}�=�D2��\��OS:�n:��!sk#m E�:Bv�E��}�g-�)rJ�T�C�wDR��Z'zڣoFpä��Ծ�|s��$r�K�ނ$4�\(fj9��}Ǻ�={c~є���j��O5�s�1��b�����Wu�X�{W�k;t��]��jYo���I��3���2�ے����'�B#}����Z��w�NށX5�T�Uy��_�'7�Wy�;��Zwr.�h"��U�+2��Zfa�����m������;�pt���i���p��|�w!|b�'*h�`�����]h�p�|
D�����߬���.�O��x}PkDZlF�Ͷ��[0N(�j9E�Tm���P��SE����:t����o6y����O��
S�4�b��i�#MT����b(��ӧOOMɣl�m�����Z��*6�$�kV�O&囖b�Y��ZWM���WN��:zzs��ؠӪJ����J'd� �ǜ��֊4���&��mZ1������ֵC��ڵ�s�Z�5��UZ��"��m���N6#�7"���1����si���cVԚ��Z-f�S�*�'U�Ej���N�4訆�t�ƵM��5��AV�ѳb�6��9bm�����j�ӌcCS̜"���V�F*�+a��X�tճK��l�SP[h�6�����Fٵ��6ՠ���أSm��s�ͩѴm�رSMj�SM&&؋[c��j���[E��+A�[F4h"+�t0F�:)�6���	E���~���H���#�Df�|���S��)��<ko��C�2|��֙|O�#�S1Nq��m���q��)'a���	�`N�`d�����"Z�}���\�;��=�=����!H�B%V!F��F�Q��B?	�0b;���y~��R�fa6U��W��.�X����<���n��+�\��{�o�T�B�^O	��y�����(�L<�^g��b3������<q�h鎘�7p�Nz��}�V]�z�K�i�V!J>J��J8jX�/�ߌ���;��/}fmL���]fo;C��=�atW-;ɝc�{7=�T��V�G�Iw�M˃��J��D�N*�9������oQ�=6"�T�z]��S�Y��	#{@H����?��'���-�-;�]��E|/MhnMmc
UAd��n[�O�L
(�@�v��{Ё�K���߫��*�rmgҥ�T����:�ͷ���yt���>f�&�[�ݍ>p�1
�¹�j2�of
�k���;2���.�e��U�)�ˑ��s��ޏ��~�zUh&w7&�Z������������3k�vl�2���p��
0�c�9�R8�0���og���W�x�72��@ζ�O7�2�w(X�U����^���j��(_�<T�{��/�xT��HRD��cu�^�%�ˢ���9�޷Rp�sH)����V��M�8.�/��♴k���jU���e.��sս�䏪"up����e	�q��r��w��{���bqM��]�\-�l�%Kݥ$�p� �> ���|(��"�Ui �Sϝ���N��5��U�ia�n�^m��$`�t� ��M�r�ԥ��p��+j*^��7u��
f����X]�|�feT5�۴�s���j#��\�Y�T��6�T빃�|09�y�|�u�}
T0�x�l��+� �2��J�7=��l��)���{�=��2YIΟ������U��h~�kW��Q���̹�]K ��'��UC}�r��T��ǟ���v�N���(6A���/d�Kґ�=���dz����/�sבx�"�e�TLۯj��N[O��i�.o��mENc��ձP�yz����RVj}Ҏ�ݖ
�&"�������md��k1�>�p��2��(����5�U�X���]�u��$AM?=��8TD�h{��-	�m����q����gT3��%E��T[����V{�[#�+�m ������V,���=�����5�qChh��(x9��ȼ�:��"���{���LkiF�cT����/��ze7��.��U�~]�6�(m�K�~6*D���R)��ɇ��)�=����M5�Px��(�姨���Yz��y�@�3����1B���װ86�|�d�����I,���YhT)��3u���fi�]q��%*'ެ3vC�g���E�J̝7r��gUe�a{Fm����>Y�h�4������gqRM4F����Y�;c}������b)b�bR�*`H�h�T� �R�f�^l~�$���?{���K�Q��fS��9�<�6��y�E��qz:.d^sc0i*����gۆ�㑏��j��Z��\�u}9o�Xk�
��C�r"0���Q_�^4���Cr��]��2��U�-F��v��e�jG}�#�0�SUzכ���\�~/�C��}n�Cx��z|]�7.�pv�*��ޝ�^�֬�F}�������9�C��z�&K�'|)}��9��@��Wh��{/���*��A�Gp��ty��NS66׻g��~�Kl5��/)6{�x��E��E�z�X��S�<��X�|�'|��"k1m��)��9�6׻�:f��B�w��*cމ峔^켭��W}�6�=�B���/K3ʣX����xjUUɿ�i����1�����˿َ���y���_�%e鴾SޛJ�n�#���K�J_�d��b.�n��iK�\�)�g7�{Ü�\�\��S��,�[>�"�ܕ
qܣ�_r~z���q)V=���Q�j�Ǚ��o�)v��&�csZ��K�r��S��j��au������o��~�'�>�?Fږs1[bއu{�<�&��F�n�W��� >5}�?s��)�@r�X(X��z�!^�J0���[����:K�����%�sg����3��=���b����o/$ԝD��X���PrM�a�
���2-FF�f�� �~~%�@���%)�V���ޭ5r�;�f�z��_�8�|f�ZkX���4ZÙ�_p%>D�Z�g=�䍠9ev�;�p�ٶu-{ԥ�jp�¥��K�/��CGa��=�Q{s3ܻEi�~}L�x<g�PYz�\�y楠�w\=
�!+�a l���]��na� [�y�ZX3��I�x���?T3#s�2�V�m]���}f��Ӽt� �3	`[j�#���C������)T��U�%:�F�Dܿ5��el�ae,��'53�W����q�x���GS+ˏ������T�/�q�oi�,��fQT���[�	������<D��R�2A׵4IL�j��]T��m��B�j�i{[�!UD��9�b`�or8�bJ$�E���RU65��Y�_gF�h���0����A��ѐ��v��D>���d�q��@���LώD�3�ɪ�ӱy����f��՛�k,��v@%�D�=���FHX{}�u��3�xY՗��6eLI�9Uqټ���2�M/\�";�
k�8:DC��@���r�GP������O���ێߑB�┏^��i`tK��(�k0�f�1��d�]=i:�7� :��m;4���x��i?����z�m@zu���y���Ʋ���M�mc�v�of,��WL�f�<�R欥�c�Zu���QSw�R�˄�#֯9�?y���"��h(R�)*(">? ��ޚ�ռޢP|�^_�#��}�H� �� #6Ξ�a��DKl��	�T��p�f�3Cպ�9�X���4<�hmnc�b�H��U������B��#ε1����[+�k�yⳐ�OT�4䙧^����q���mk�"SE�9�w�,^��Ȫ�ʈR�%�7O�����fE	9���4�ދi�p=� ��.���t̟�Ĳ��X��+2şx=�	�=��{�!;��3]�&�:L	�z�R*�6S"��g�u�d�ݏ;�}}���Y��~m��ӽ�+�����W����;�n�ڽ�<�,N�|����]�D�����_��k<+5�8�N��>�O�u�'�J�B�H1Wt#� �#×�`Q#C^���N��|gg���u�W'��E'�Q��B�f9y8��Q��\��n"o7}��".�4Mn�������,�7zὈ��HVa�9.������-���;��8���穟nhR"�c� �C"~��6��2�;��=��*Bhd�]BO���L�iZ��n��A+lK^!���������*mp{�˩d?mC���0�`u)$N�;�S���XLb�	��t�I�a����s�z��(-�j��z�;�#��ݾ���dE�h��U��X�s��y�GT���^c��jr]K��M����l�o8�~����0�7�i"�%�db��& ��>#���^�〟o�P0��) �G�P�-q�Rt�κ���W�������)zmq'}��$ԥ�j���q�<7�J���A@�y!��O��v;ʄ��yP����q��Y��f�)��}�6��Ӽ�y�l���ȍ�%�}!�I��X���6�僶ၲ�4a|f�H�F�U���%�T�k�|�:htE��>t4_��7^JPB��3��1U����ø�W���ay�#b��q1��;σ�G���W��ڸ�qmf�	��+�NX��G?��@e��F1�1{��3��DWN�)�锘���5ݖ2|[3&a�n��b��x��Hþ�2z�r.�)'���9�y֒����(��q�P��uи�a�0��P�2��(L����6C=�=��B�^����?���6J�e�J���Cll
73ڮ&��GV�΄6l]٦�h]�5�[��F�V�]�����I�=EP�ߑH=e���|���k��x�G��a��o#n��ι�TRsc�m�%9�v
�m���vWA�}L;��N�m����ݳ�5nkÊg%���(��o�+ed
:<r�L���T�X�](��U"��:�^�:6�H'h�]�����۹���������`��:k����3�ս�sŢ(��_t�Y+n���"l��0 �1�;�ܫ�ِ�kw�J����3��o���}ܯ��������(��h�H� �
B���V <��?f�+T���a/�(��9�]��E�'��j���rc0E������8�錼�DoM<�v������\>�?�:����*-n`"���|�J�/V���$[f���%8�g�Ts��K�#Pb
�X|0+���P�|��I�<oҋ�e�Fg�O7R�R��u����`;�N�c��U�xLIAZG[�=R��R�����k92���.x�,z��iD�Hg�J��kv����kF�.x/������ԑԴɑ�GC�*Z�+�M8~�I����n�����\7��r�ٳ�]�h{aY_0N��H���y��f��uOtZ(�=�ц˯e�V2��2��P��s�lГS�\b��*�Ȃ�+��"��{�vR[n:��)��j����:�����z���^2]��h�빛.(ŉ��<���/�q	7�+3�{��F)ַ��
Q��#��K��D���S~���_���Y�i*�1V�LM��mݕ|����JY��`,��]O�+NR��fd����qB����ڎ
!P���T��d���ڐj�LG�C�F��|H�g��E�����O��7���r�׷�yDQ8#��R,`��hi:�%��M�+4$\}���;��ft�]4� �Va�:���n�aZjP]or�.Ku�R�A�o��ګ��tn�'���x^�[�\�������3L���4��{�E𮫤��k����vy�ۺ��6�.
Z9�/@��j��Q�w�fz�Ž����VE=�@�.��h=O�Lf��F}�	A�Z8}t��{�VL����v�Ѻ�+���^�[UM����$:T�W)�{�t�����~K(V�a-���J~u�g�z�ƪ��
�b���F�lnfӡ����1��Sy�5����^tW'c;(Z{�u�ɂ7��G{]����zE\2b*�f���0��·,ժu�o���kfQ}J<���۵�ڻ��;W+�*k#MU+x�2��Re\}	\:#����
T�f��2�S.~H2t!�v*S����YUw���}�w�ٹ���ő!�]*Qfj���[T1O+�G����x���tU����ʋ=:kyԱ�^1ot��x����C>��F�U�~Q]J�/���Jz^K��v��M���h��;�3`�\g�ăv�XZ&K%�=<�qCS>�}vD�&A���b538�j��&}�j_7з^Ш��O�o�6�P�/�eמ@����<C�+U=�
r6A��oa�~��>绖�J6ٍ6^v�I��:|�glKY����)"\��-�]\-V�K��|����'s�����̬ѝZ��}��n̹Q������H��g�e�WS��u�c���We��g����&�c��1���[J��;Z{S%k;�6��c�W߀���dd*h""Z�*�� � �!"{��ƾ~{}�������2��?B/���TS�ORoP�uX���������݌�����#ՉvO�������\A�P2�vHA��E������1cC�W5;Z��Ɨ�Msl��� [��$�p�c���c���&�:A+���R�<=dlg��<���!�V�q�J�8�`��v�y�xd���a3�]q��rR�$�^�">��:��Ӥ�{��4�.vo��N6�"�$���Lݏ��]�6/{���A*��Q�gO=0��f�'�T�.�.��q87�qV�i�W&|m�ݪhj�X��*m�r'5M���"�P�:`[�����d��~�dH���8������u.9��%��UM��D&�jBm�%t+�5kH��,��~ܬ�5#xؖ$�/2:�4�s�=�2'��X�r�O�1M2��X��Y�,n��Y;[t���P)������V�/4��R�3y+�zG����G�C����2�މ͈W�I�U@����<^��5�b����aEE���^4Rwlk���l�����^�roVxY�����b�0�I�s��Eu=B��/�C�)06Vl�y�޶��f2Yٜ,GĴ���+�����m��ٍW_A��(����F[�9ܹ����v~p���ɘ&�D�;op¬9v�<Na%ebG�o6,9�>��D�n�2���� ��&�!"*��Y��7��s��KVo-���by�U�{zh����x���PYK�Y�1W�kg��&��k������k^;�ɣڃ���
���^@�z_�^����gX�J��J��<����=�wd)�y��1�����Zc���Pw�z��!�Q*�=��]�Q#��.�nj/���j��ihM#DZ��]X��x�T�"#�z��T�^�%��م+��c��	?7,��♩��v�E�}�;7�W��x��.�zA;�
WzB����<��%�s��6��O9όf��C)>�f��I��V�3j�mRlNƅ��35�?
N�yP�Z�,���X�]>�y��gor��u��:���}��G:DmI����-�������PXL>�BB�.���oZx3ӫ�GD�pN_���9��b�e�I�(�/^"�CHfb���!����{�7�����}W���G������N��A���^������AP��G*JZg�lC�ym%Nӑ�j�}�s;❨3�� H�_���G���L�N�4�T�����V����+GLȤ�+�q�������k�Ӷo>�ièP�3|����"���}�{��t,��T�"�����K-֍;t�I�>�F4�Q��j�Y�T��fqO1��>��i:<�V~�4����ñN���t�p<f���8�2���0Z�Vd�ͱq[���:�ʽU�eX�@	����7� MBq�@�������s�x�&�~�"� P��&F����u��u9`����N����T��ajZU�������2�����f���N�y;~���i�eh����Vc���7ؚ鵼��f\j�,���*�^�.���E��T�1�T��L��܎��6��Di&�Gy}B�M��΋��Њ��S+����G�՗@vK�X�fW.]t�2g4X}9A�Ց#L�8��U����{Õ����"z^�yO��[4�����F�VP�r�� =*ҩ8%�ks���3�)#�NY�k)��o.��T����2O��\E���SF�\�4t��U���e�fm��9sC��JA]�{��X���̘9]=����j�&�@���
��T�����a�z.)z��X[� �?5�=Mۘ�;$W9T�j&��5]	�m�{sA�W���'�t�JkA=�ȣ�V����Vf�	ϑ��)�(�R��(V�ιp�Ar��2boZ�tgUJvj�4��_q1sn��Uy2ܦ�C�$�2����T=��K ;�땙c�+;����&���f�SSm�U>�'���'Pմ��[�_�y��O��5,���˷�9�8K�&�C,�����Ո'��wnb�s^ aC�s%��ue͕a;e�������v`�)#��u6͞�eq�.Y��Cowq�����t"�b�0.-{Y���Ʉv�(�ll�x�6��Xl�C�PKCI�M8����qn��v�&�`��{��zPJ�����=%�{4]����Gk�;֢y�/zlb]X�[ΊjE��kei �y|+g_2��{�j�C�nټ����	]!�.SyVUB^^�̋���M���ʺmY2)ְ_q�!T��'�J{�;X�.�'�"��U?����O4���ܺ�h��U�[5v̖@���G���mjf�1"�緼s�J=S�|a�h��٫����Srwخ�����e�3�X���$m�w;POJWN(�g'`�"p�x~���*�`l!��a�4��U��Hؿ`*kukyC��l�4vN��@E��8n���F��Þe��\N:ճ%�h9kaNT��nX�������t5����Zꊠ��c�:w���O#�Ѯ�f���e�k�$wY���j��G:��Lz�'9�x�͐�Ń8Vf�yPv�DZq�U�F�kNױ��u%�dxM.劊�eb��)4�)��3�M��cm�s��Z�+��|�@��+�s�4����F��Zv�lN��PPR��<>M���"(���:-��l��[h4�֨��%.�4S@U�:zzt����-�Α����at�cc:vƬX
LF�===<<=vJm����������I@V�li�[e�b*���gK�������l�q�{:ND�T��5AV0�Z5�ն�7����ڶkTC@�!9'*)�9m��xZ���9�mm�h{����(���эn\�4U��S���N�:(�5B�)�ZMP�M���#;AZf�Ztbl`3Dւ�ALl�#e�4�Z�IUBV�Zk[b���j��\�Z(��;�����Zđ��)E8�lRRU P:hU�ӣAT�и���׾}|)��v���e��WR8K����9i����Wq|W_Y�8�b�^Cܳt�\�������}?�?r& "�"X�	?� �� A�u)�&Ƚ�_Nw�TU=,�E�v�t�8+�ϕ_��'�����+m�C5Y�OU�v���I}��Dg�DE��+�f#����n�m��e]c�<:�U]o�eVEn�w04�a3L[s�&[h���q��,U�ɓc��_���|���݃��GI�7`k��Y]��+��F[�y.��QI��M�U�����^C������M{=q�Z��|"�U7�ہ��2v��ph�����)E�:�_�Qi>Ϲׁ�Xά!���b6>X�ۗw�Z:"c�ֳ�Bzc�h\x��q��:��-�;�T&������Z[C�54Q�&����w7{��+8�b���U�.�sO��m�ö{o9]5�P���(��]4��D��,��`<���M��^{n���IZB5�=?ڟ�O'����އj�MVvL=�4�u�KA���sk��t�r!�C>�b~��JYCcGR���9��qx!�Oާ��l\��ی����UY�{,��g�bg�זl�.����������:��$нʟA�g�f�]��c�W�f����Qv�΋]�]��c��`�ȗ�3~�����^�)�8\����7T����]�l[t9�����gKB��j"f���ӌ�=����r��P��H^Z��n	�cL[�IX���`Ʊa"�T���$�j�����I��H0�y�7���h�V�Iݏ�輎�491�N3�F�5,����n/A��|E�3G�)�a��}��}�J���_D���N����`�7�<^ǳlv ^6��g�m�.(ŉ���^�,�KYW��� �����6<d4h�LVg���ݯwa�n��޼L�`7y����]ۛs����];���@p�"w�U=#<�J=�Pw�(~�m������eJ�^����O`��铞�nu��bj]�ћw\�mQ�u��fEצFW�{�n)���nL��h��-)Ge};C��^�/oؗp�p���pm�'Tۻϑ�w��j���P'DE���a��S�37<�h4޾n�i�wIM�=�ڡn<B�}�lwe
��>�"�}�20X/�*�v�!g��;�^+O�o#Z�k�[�y=[�Liu'������\�����C0=�E�
��+ݷ&��P��;\'cK������g��mN�j'��5��I��S�M�m��{Ř̪�C��6"w��y�jõ���BN+�g�u-V%p6���a�3Or�^�̤��:��y�N�15���T�Qj
×@�{v>�S�̂?���*��f�^�ʟ�[�|����5|Q��^c!��\L�w�� �|�̕H_�CQ�J�](:�$j����y��N��ة��
�m��܋�INsnt&��m�GMc ~-6���~�
�$~I��E��ysܲ�Hm���o�y^5|r�\��D��W=DF4�2��[[�)�9�Ƙ0�鎃�����^�������u�>5+C��$���{��R��j#���vD����{��5N�R�fNV����ݩ����J8hˊ9j���d�X�0�b��}jh�D�$r����gU�I[U����/L�O׶�x����P���]��/��鯚 ����z����#�j�8Qg��akЙ��
*)�	�WYoW��V7F�c�E)�lm9>��d�T��ȷER��A�(Tt�?�"~���x�Cw��kњ��L�2�e�95v&����إ���a���	�-���"'���('���,E�V��[x�*C��c6q]vQ�=�{�9ʰ<��5���K��J�hD{@�*T�qBk$���-͓4qM5���/��
��hw�qfF�܏�>4"A��4�f�;'����DKl����;������+�T��Q��br0�sfN���r�s_	�7���n���ôP<U<���kd��6&� yCZh�z��=�0�l�v�"Y8�}3�e,�^G���b��2�se�W( ���7����R�VH�(z[��Ŕ�X�U�i�٪>!V'LY����)�oU�_(���T@�w�*�?�?U_�
��8L�jh�~NZ�
����i�T�27��t��4�M��Rmt)��N��Z�x�/��f�^nu<�%f~Jʹ�SmP��=�P
g����ԯ9C%��'�&��_T�A���ˏ6���~̕&sؑu�p�E�L@���&?� C@�[@؎�,4�[M���j��]�݆�-i�b\�Sm�2q����`U�:�c�����7�y=V�)�?m�%G�&��qtm��ӥӘ�酥R��<U[:�^�^�S&�H�R
�}�a<"厄���r�ќ�y�i�L_��R;�"ጩ)�u��ƨ���R���X���*~N��p��w|�e��b�y��_�{D-^���U�e>���=���	U��Π�G��K�ۙ��N�oD����w�Ԋ�@�1B�6�	�	q�_T����{8���:��؆�C�^txXkػ�22\�v��[C��ԣ�����nB��	R��'L}����:n񼟣#���S��K*G��l͞��2Q~D|�ÿ'�
~�w�|e��U�z0_w^Q��	�����g��º2oycV�Kg7Z	<ĨXNqưR�Of��D�2/v�7O˺�<.�lr�v|Ûسa��� Il�ڤ=��Xk&��W۴�2�5ţ����LU'H���%]�o.v)/��� ��ǒ��2k�}�]|��Υӭ7\�@�C���7�p%��{p��k�~�0��'W�'/�[�����]Xu�;�f�~����ǆ|S�
����4�� ����c�0��'�h��-F"PB��Fu�@g^�!� �L���>����13�>4%����{���n,�h�$`�T�p�*a:ܭڑ9e���S�,0�ޙxk�t^D���5�,d��7wn�i2�A`̹C0�+��;�,��Nfv��@�cWN�jfR��N� W�~���%|��&�tr��_d�Iq|sTv�0���7)��������Y��}Ig�����*�dѠn�@~S��]�u�jG�2�t[��e�弳�z�%-~�m%�M���I[��Pu�:&�GYt�Yv�త�f#[q^��B-�ǻ��ՆFH�����E�>����"�k�Ncݕ;�^͇eT=UT3��{K^[d�V�(l�v%G�{����s�#��҅��J״�ӓ��_P���NNK��O�b�<�l�	31KK�/^�3�0�B�?;�~f�nuC;{�)-�`"���}�	P�����g�e��k��yQAF��ڡS����qk%8�]��8ҭ��s�m��P����S��gIw�fһyu�/��m���Q^Dv�N#�s}�3(M��w_m��Į8]v�;f��7��:q������gGy�b�S���%��rwG�6w�${4��G����wm��U�Y��Ք�~�|���"%�tSƿ^�=?����Z��E��bQ:'��L�ee���^���}9�����IAZF�G��PکSˍ�R'�}ؤh���L��f2�&�6�sQZ���C3��8g�ކ+��)-��RE����dH�C�w�De^{m�~�C4�f�����g��*��_.͏�u�)��²�����F�V^�Q4r����n��\1�<��\�M�gS�����^:Dm	UZ��,B��"_|>���n2�����p^KH��rB�^���zCݽq��J�Α��l�.�|��U��D�4{<���Ӌ�JO����mT��N=ͯ��%�Q~Jy��bUJ���V�c�Mۗ:iz,�Xԥ�"�U�T��চ��3(���3���+|{�&�!��藓�ׯz��g���ਜ���vy�8+!��y�D�y��EМ�r��V!f�/xOD�{f�D����7�BUz���eEB/�Al�����	A���>������u1z���:>,͹xba�C�W��s�m57�8�l�y�j�f��<�©�7���\����+]
F��?n>A��H���31���Y���wBξ��칚��%̚�u�/0i�4N�כVXP�,�K2T���:J�d���pb���{���f�\�r�-L$&��~��y1L$ek�t �����a,�[|�^�f�VJ��-]'Z�~��Vw���m���4�}���d�Ux�/9(O1�14����D�Bl���Ŕ/l��qrEң|��WZ������e�������4cO��"��)�]�T��-nfQ}*<��X*J�kG��T��H7U�{��f:J�mF��!$�3�D�U��ξ����l�{Ⱥ��?�[�9o�n<�.x���T_S�\��{euP�js"(s�e�QH�O5@���r^�#�G���K������!�ҕ�,Ԧ)��Jn�8������&:��,�j�FBTqk����l8M<��U����َ����T;q@�U�.�4Y-��0�Z���֯"�$0���3��G_mv�hR���?%�s���-53��Q���a�Jm��P��Gs��%���}x�gqI�y�LD[��Q&(r	4��+�&�OBf4��L�v�YA��Jz�XJz.+���y�U�~W������d��a^_W#�W��u��?@Zm��>�ԫ����U[�zJKګY����)guK��&ͺ�5�d�K%�0I���$�B#�����u�|�Ⳓ\�bT2���@9��K�?ϻ�*ͫt}K�N�=X�otv`\+�@[M57:�!��%{���IvKn�7O.n j����.���~�'�$�3{�f���_zS*��Z����E�^������|w�44���'O��@r�3��{Ԝ2�ڏy!qb�-����PՌ��dw3�y�X����n��P��P^�)u8��y/��9�3ӞC�Ȁ^`�9Q*�5��2]x�'����N��܆��$`�T��f���L>���m�5}}�o�o�]�j�j��;u
��E��t��ݴ5�]1��2��H�����)�EF1ְw=�f���Éز��(�����j���3E�e��g)���	�*�6�wf�ܩ-=�xb�/�>����.�M�����
�8�g�
[�>-΢�uC'ޙ���[
�Xݓ��{X�ϋ���y����m�`�w�D�I��}�%���K�h��E�;d��og���o¶#X�*��s��۩fV0���`P��:��|h����9_LX<y��rg<���v�S�so;T�͑*3��
��zN�Rڔ���ۨZ�����|b-�-��}��M=mVr0�PuS��f���Dk* s@�����.�\����/́?7�Zӽ]" ��,ۀ�+��?{/v�j��-E��a���L��tR�f^�':�}�z{.	�'�/V��z*4�
^��t��k9�S�<���*��Һ����r����tO�Ui�}�SV�M�;�+��L9��̦rN�A�oe����08V���j+@�6�?��	�N�k����Y-�Kȉ��O`9�f�]�w����"6z�uM�w�Ǹ���,R"���+�AZE��M�`T�l�����*���FSSi�QUCL�d��]���:��iZ��k�d"�� ������T��R�鑳��� �@Z|N��~?7Uw�����[X�apV���>&���.Ļ�:"�p}4Q��*�Z�%T���>��Cn�U^�wT^���N�g��u��8�lǔ�a����p	)y����DH��{��kf(�g�o{��WεN7�a��#����|�A=CE3e�a��؄q��󈞡�]L{4�ѓJ���x��v(��>r�J����S��o�H�����M��]��T�����gua��t����L9I��x��>��y�t���~f32��ԌW���w���v$�=<!]V�u��&a���i<n�&e-�
�@��>X�|�6Df%5�Э�L.�Ȭ���Moa�ccb߲h��F�E�D�I_$str�x������{���}K8���i�	�L����R�ض��9�$a[��^C��I\;!�tw�T�uŝ=�:�����n��fH���U�-7��s���uY7ef�s�6��냎��7',1�Qi���gZذК�'���J��opĨ����ƁqR�.���{x��R�_[�j����}B���x��)�N�h�f?�΂5��M�䓍��~�Bc���ͅU޵�0D=c�O�K�@w��u������-�����S�s��Ӭ��(����1�mԮ�?�:��֡Ge��) G}M4吝�f��C_(�����U|��t���f��[kQۙ{0�_C�s����˫��]x���@��k��h�޸gj䤳�����u����N謆������@㡫���YN�|�n�F!��TsT%xdZ��vڔwL��u	�TGG���ޜ�2_W��Ę�Ɲ�������P
�0�]�=_J��	S��jD���\���7u�f&IL�f���Bj�]c*j{�H�e�����3�a$k���_�W�
?�v���<���G[U�
�Y��y�
zO>3ƅ�=\F�ݲ�r�͟���i��
���u4�͜�l�(�6��[�0�RΙ��40Yѣ�ϻk�����q}了5�"6���zb�Ax�ջ;(�֙���F��l�����"f
�H�]��}!v/b���X�{��e�KS�d��6cm.�B�P-��Y�Ʀ��˿�(jd78�F�)����N�`����n�[,շ��E��تT_VҜ��n��i��i�]�v�T��6��׻lDDD�D��	�<��DT���T��9:� Wd��t�p�j��7s�AH#'ۨ�;f��ܴ�UgOR$6�n�͈�� �xj*Cp%D��@�,��)�ڰ�c��ֻ*nB�j�����a@�FF�G���_n��ދ8j�4��V���q�ɷ�s��C��("���o]��T^�K.�ŝ����tar|jN��[�;gQa�3L;�g*���݌�.[!�7W*���)t����Aڐy�88�5`�V.��r�����!�E�L�k��uk��O�-c���Rx��iU�&�^���Kp��Ʋ�~�{WC;���0c���A��t㛖0.0L�8,|�`���%��pv;cw&Ytwbf�qΝU¹���c#���P>�X�\X���2�.	#6V���+p���J]�5�3��p`\�	��$�+"%
�j�ky��a��U���q)�)7j����]{-�����+)��Qő�ХM��7@0V�j
D�q%.g/���VH���T4�����*[9j64^������.�-v��"(��մ���+��PUv�7I\80�uՃ���� w���V؈-1�s�+��
�]./v3ԪN�2������,�w�)�loQ��۽t~h��:��,ո$��+WBȤ��H���F���&������ytB��q=;�����:j�E0Ғ]�O!4VP��(C��&_-ۑ��T��N��Rq���sٷ�%v�^���20�E��8g�d��^R��\M�%���{1J�Wۄ����N���9����U����=�9\��U�=/�s�����2�`�;��m���2�Pz6r���D���D�D�S��v���'Nn�wj�nv�{���g5x;+�.}"����Ҋ�]�
��ܙG7w�Z�͚Į��E|�u��{
�ӧ��AM������G3�+7.�D��)ut�Ԕ�*tm*��ܭ�U��{_D�}�˃F�l�t�ki����r�o��}Y@����p��th�Z�dĢ]�D��h�AJ�G5Q�0;��3r��utT:E����� Y��$;�����w��#���B���L&�^������W78!�t���i��I�V_Q>����*�l�?��C÷o�OW�0�n�Rف(nlo�V���v����bD}���OQt4�w{4 ���\+���J���X��Z��Rh� ���ͭ�G�c}Dc�T�M�lc��ٮ�T����)<Gkj4{0�y�]Rh��2f��B�g�	�Z��4���:�ʜ�y�&�Eg*³�ɒB�����)��.�K8�k�Um�Bf�(hR��ܩLH-qC��`5���Ӫ �Ν}�t���H�[LbV~W��m�)�q����NG7O:y�<��h(�j*�cc2��0�1��:\Z5�4��i�v�p�'������ER[%��EkZ�Ø��3�*ء5I���y4�����㇧����J{!B{���+Qys�"�:kli6������F����=<===�JZɥ���5��{����!J�:�b�T��:
X������1HQ����4�h(-����k4��Q�DQkESG� 9R��`��$�l��ċ9�sj�:��@Ci���QCI�s��6,�T�G��TF���o8
h9�\��UUr�PQUŰꨪ)4�V�H�͉����i�喃U�J�F�-�M��EA���㤠+T9���clPU6ݞI�܊���S�5ʓδ�-�El�`�+m5[h��HbU��mSh�1�Lh�m�������2Z�HPV�6��֪j���#� #%J��v}�o2�Ѷ�NH���!����-�Jv]D��$�v��7�;;A\�!���;����L��M��،g3#3��_��W՗0�����-�d�ʄG��T��J��+�ɛ��ߤ7r�����������Q�OU;��4��d%;�{��4���dשׁzFyR�碝&����w-5�\6��9��v˲�;�⑏���d{��SޛK���B1�U�E�ANDjەoR�*_��U�v�n/��#3n��k���!����l��q���e�X���Zr����ѓ�?-񮮔)D,�uo �M��0��P�~s~O�f��"�|;{j%FJ��������hu6���W�t�����;�yAJ�cKEq��qǹ^tW'c:�X��Q�LD�R��{כ�(]��"�#�����h��.S8�r���zŲ6MgPXĹxY��-�f&��7]p ��+�X����n��V�Ҹ[j�h!��X�������H&����_W����7+k+���.�^x�NBye�x�+ƅ��Iw1�ɜ�J#�ǚ������`�=�$ș͜����o�}�L�/1�a~3	�{�V����IJ���'��"g\)�_qT�iQ���Ye�v��W/�ԞU�mUt���r�l՘q��qヱy�[{nQ����n�mS48�߯���8������l0���a�7�+����x�y:��F>�'������Yv����&up���Tԯ�\0"�����Z��nʐ�Q�f��U�ЪP��q�+�~�f��r+��Ȫ�a�.(�\��FK%�����L��Ϯ�kCS/���;����6�3 ��hM��~k��q|��t{����qT���ިO^Y�2�RXm�1UE
��mR�3k�s�>Mp� r$��O�[��QL��h��q:�C6��Fl&֛i��y�6*}�ΟY[�UG�yY^[�A~� �/���L�<��ǫ��t�Dp�e��gj{/qWU���1�o@��z�KW�X�c����c�P�DO�F�ҟH����r�s1���;{����<�� bŜYg�`F;9WI��nY�s�>�Կmg�#<$ֽ+������w��rf�h7}�C���5cQ�#�̔gv�j��6(�8&�`�������t��=���X�D�11��&i�t�-(2�`쒁�Qf��>5uږv�/`������f^}�X�X*s+!��`o�7�0{]�yȎ¦z�I�s��2=j���)um�[U��-@M�=��m�-���ǫ�ݨ�J��í"�똇�{fjjm���x��gƳ�W������驪��L�f{�'h�g_�-���;X��^X0A��T/�Zv
�b&>�۰�����ٽu��f�����]�y�-�� c���Șخ��2���.�f�EC'x�A+u��2�Uu���Ͷ:���afN�J�]�	���Kn�����
[�3��Ƕ�uϾK1JTl�	��Ϗ@�9�t5�z��:l�u]�.P�Mk��/�p�b�h�n�YX�ɁCא���M˶u��vcٸ�Y�W���|+پ��ER^�����A�GE��bS�	p�M�m+�63���ŷC�q:��%���}�1��Ǩ��������<pf?
�2��S�U���R~mO���
��!�+ZPr��i��p��0I��W*�YEG�?D< g��T6�PȖ3��Pޑ�LP� �\�è%�*hf¥��H��j�V�S�=��Cȴ`�W�Wҡ���2��t�Ѭ�w\{�{U��o�nL��K7sq\!Ѐ&��L�-Ak\�mt[�A�܅'��T�k�J��8��g��,��ټ��M_a������R��O��֢FK��`��b�q������~y��{�3����m~�@���P��{/ZL�u���Rצ���>�����@�OU�e�wW��A��b��P�r�zGF'�w�:9H%̌mk�F����A����a��O�qח���o�b�$�ȱ��e,C�4�`�B��F�w3n��"�HbFg,<���.צ�7ȋd��u	s1:y�s�~�4�����Qq�m�JI�����{IWw����[�.�ힲ¾���yYM�J��o>��yI��k#7�w�wi8�W4����#�c�k����gO���~�f�Nտ��5�c	��	Y)��n�g�hcgv�f!�5�"Aj;�����Q�������������'@Lq������}���d���ޔw�:�f;��N�l����h�=`��$i�oa��P�cȸQ� KP���.`�/����Z5�Y��2q;m�ً�z�+��fע�i���i�N(����\,�ꐹȺ�2E�v߮��yX���;�ڇK:5�b�:�5�dԞ5�9T�~KkZ�F����Fz���m��+�Lf>��f��
��wbP�#�uT�eBLJ���.��TRs�Ȧ��o'�N7K�)�Uո^�n�;�!�NG#���}������m	�f��_.R��eQ�I�?q�_H��/,�4�}9�����6�D�.7g���"|S4z�>Ȩ�h���;H�Qk`"�6����Mww:�������6���@��Z[C�ʲ�41�|������ �eT(x=�Y�3���v,�9|�����,�\�s�2�r1}1���X0��ZFG`{��%r�'#:������cF���b��\��G#J������6xw�l5�lk1j �~Hݿd�#�C��)0��|VT��i���\�yn��5�`�[]��X `�t>�=xa��i�qy��u���)s����q�T{�W��a���]�'�� �T��U�Z���F\�ݺ�d�����0oz�=FRY��o���zE5��.SJ{	@,q��@X�.�[;"#A<�OW�+��襕ך����K�}�O\�:yP�T�|�y�	�l}��M3c�
��~aN�%�W�}��4�f�:	�\����E�O=:hu���N7�C�@}�5X���-I�w�D���Ƈ`3k�Y��'`3�wi�Ijc�����C�L�;��N]��{�d7�?R�ϧo�~b���hP�X�j���Ԡ!Dtb6-��B��#��y��w+Anv�QZo���mvf��Z�Pǌ�z&Y�4�r��ų���Y;��US��y�uO碚j��k�,ۘ�a�������U�p^u�ʮ˔�>�ӌ�\�>ylۺB�g��!�Q�@�n_C]5h���МM_��
���^�ŵ]�3�f���82�����"[,^��w��ۼ4�P��7r�VZ%T��1��z��ZW�FEP�5�2�<�ʛa\ac��J��B|ЖP�c�k
i��t�	�3�UI6�O�j�ך0�־<�)��rR2D�u'�{y�Y�%GY<�Y~T<�����V:No͊M\Q�/�����/x�N��rJ3�dܳ�@b�]�<���K�G�چk��ii��2 �Y���LSw��
�c��1(rb�,��#:b�U�m�?	`�#dA��g�k�3[$��9S��7�u��f=3�]��V�sW�{jH��z�E��M��T���Ndx?-�s�c��j�L�������{�����t�����c�yCoܶ�^��Re\��N���Ջ���]��W��3a1��fRu�e˟�����]��T��cL�#�\y�zv��Y`�{93�I���!Pm�B2^Fa���S	Ԧ���5)�Ή��J�*:ĳ)[k�Ч�K�v��˶N�o[�l^��Ƅ�-�����؞����쮖Gs�}�H���h�7ޠ�Xv)Tt�J�>��.�W$8�"���׌GBc��� vq�w��C��;���lo>6lf�%��d�K���o�u�w)`��T��H;��L�az5���q��QG�vWYo�E��x�l1��۝���r&��e]:�:k�W�8@�H��)���	�$E�w42i���83O^O�>���Fg'e�/\R�Ʒ�<я��Ij%4=|�� i�?y�uO^x�x�Y��zfw�Y>�9�ώ���~�a�.+Y��xY�ql�U�j1r�곦���{c̓ö/+������[�������U����%�cy��LX�%�m�x�CMռ��|c�sL�u�tN;
ƞ��^�@�C.�AC(
��+���+��$_2�����3��[)P6U.�{ohl�"<���n��S1�m]T����	qؑ�j��s��x� >�gN�
�NJ�&�O=붸�̗i��ߞ�16�#���4�6ΞU#}�:��s��y�N*X��T!�
Qg#۴n�SC^�c�*<�mBD��=�ㆌf�}���;ػ^��R��*Q���EG���#�A�}S4]ouQ�c�0��B�s�~k#�.4^>��mH�]�i�U�vTB����J͙	�ٯ�	j�u����Z��<���'O��K�=�y��7���wa���4ˬb�omx��c�Cϭ��s׮#!�S��;��:g���y����Q�;=�ߩV�g@�� ��M{ ��E�{T�u_ea�x�Loʄa#Ⴉz��\���v�ʾG=0<_�L��[��V�Ir��fa���-�,Ͷ��ӆ��E��d%;&�[9&j���BTVh�}�@���p���i ��i�XsJ�vO<������ʉ{��2
��;��w�oq���	��'l��H��ZhK���ؖ:1N7����*�:���h)a=�d���^�N�_�p?zfܵ��(���P�P�Iq�1w�ί=�t��Ob.�*b���ϡ#�4�s��N2"�⭤�壆��K�-�3{��lN�J��f���Fv���]E}`��,��نվy� �g>`�y�~_=�E�c9�>aC;��*��7IgMӃ\�M齛�tPuĆ�N� J�=Y3�D�찺Ow��{͸�bc��`���z�S:�V������.PX�:j\���v�����h0����?*�T��`�����V7"n/yoG,md+k��`)O6ߖ�4Y����3:�H�v%�71؁� ?��]���&}R�ݮ"�4{Z�(��ܫytt0m��ز���5 s�FГ;#�2}�{"��ɸ�R����j��>�V��F`v)0bU����8W�h�O�WN�X N`-�Y��9G���O3X��f��T1��h��mxs�'k>��A�p�!�LV]�VR���s��qT���Y�[��E�����mȢO*�2���S9���5[4i����J� �R��`��vF�M6���V���V{�`������IJb�[.�+�#������T4Kõ�32��գ��IBsc�s]E��>�U��Ԫx�ʬX��y��}�~��uXլL�׸��q��|^(���_��v�[B���U�[@%����l�y�.�����EĆ��5�J���O��$����Çz���[Vf������k�Ŕy5N�{99@�V����	��J ^a�]݊&��:�e=͜ V>����l�L;g˲�ɔ��0W$��Ӗ6hձ17 ��S&��賤E��?�5�a� �>"��?�`�`�0o{�%t�~���T��h}�-Y6Ⱦ
/��rQ�0�
�ۃ�Us�hj�Lm�k(����8i���ʯ3� �5Ȃ�]ͩr.�GmU$��>1�O:m�����y��{�+�'W_G��,�#zn9},��Y�������ĝx��\�n\����+ӝ_���b��|��w���sz�AΌ�kE�"������5=����N�#��n: �2r@�����|�O\n�,G�Z����>�B#�P=�]�~G�p.eVd]��:���+�JQpq���I���m}o�9f��;��OC�ׁ~[�	�t���4�*U^4˝���^ﵴ�G��O��G�hg;�Y���i.o5��<+�65ƴwU9��=�C%����f��'��z��?�'�#o�@EH�ru�r9t�`���m����������X���$>���`X0���(�l��/Ϲj�.�v�O\�e�O,�_�`����ojN4�+J�m��,QX���Ӆv���5J��'(}�1^h<�[�C���8�ۣC��/h����;۝Ғ��&]��I�f��f�9DE���D�M�� C�*4Cm�l>c�3!n�}��X�u�����[}C#6~3V��U���Z���j���/5���FN�9C~��ʅ#�����:�f�4����KM�L2�̋깘S��R��C���+h"������0�%�hn�ٻ��U����nS��pʌ�2� �o�~}�t7J]��wxB��h����5�QkĜ7cq�
��}T��m�$2E���K�S��6��<u*|ݼ�%�4�iH�6v%Wg+���5!�
l�!k�}�y|s:�M��V��q���M��.��n��|WH�oh���v�]+-��Qc����r^�֠ �S뎏WXN�79*	Q((Kq�5u$!s��6�e3!�O1¦�s�����=�tn�O�\�f�����qE��]��	;�T��e��5����l�g����脍I���A��_^&���ع���Q�K��	�I��h,�Y(f�.Dc��]&R��Ī�N���v��'��:`ҼFct�טW(�)*f�c�!#J���}�8�Ma�E�x�{P���m]��z=����-e]�j�蠄�,���i���-
9q�e�ÂC��}n������۪e�(�2�m(Һf�;x��ڭ��K��LqT��������%� 0�ZL�0���s$��rd�&�Z7�v��Kkq)[Y�kn��F�9O	�+5MD6���}��5�X�h=��]�kNX�r���9ri�,��\]�Kܕp�y�b�<�y���pIsT��8�DD��6�*�D�)�2z�
fͽ����F{%�s.���&��_	<)Y�T�U�rWɾm�M��X��YA��Uq.�֎�f���t�2�C���%Ӿ�6����&a�JԽP��`�N[q�:�CnQs�tT��aE��+:��jX�(���ASN����%oK�]�'V<�/*c��쬬��S#��(�g�)�|z���͕��o]X��s�փQ��rC�h�)_`��|�tvڢ(vf���9bƸ�7u�N�.t�Jx	�Ʊؚ�,*���C�<�r�wo�(��۳��z�J�{pq�Ң��w\(-�W��j�X�赕�4R&c$�뾌���4�/[2uc`�
ط�}*�v�~1rN�k���΄�f�Z�E�QZ�6]����+�q�t�mf�;7w�u��J*��C��a�ۛ-�7��rm�-n�]��Si@:(1d�o������L!A�Ux�����	�e�1��1\�0�T� �+�uhbͬN�٧�,�̺��ŚX��6���%����D��eHgǚ��V M���XT,�������(ND1B��u�[]�^��+K�s��U���B�W;^�`S���d��z�K.��WJ������oC�Du�t.��аgo6��o�e4N��	n_%t�w=[k��l������b����೸@	*:�M
�M���D��������R
����cE�Q#}	k�Kv��͏x�]�:��������3�d_1"�pk�y��b�C�8������1��J9I��E��d�/����EΨ#y���|1�Y�i��g\�Le��+�"�Ɓ;3d�2��W+(P��`�%�T��욺�����i1���6�w.%�,���	�����<P6p�i#��'���zw�����Xu��g� *���,p��%�[�`�k�ec�r�1دa�g�8;9L�/��s2So���G��q9���2�+Ȧ���ӪNA�E�t����v[�l}�I�+�[�\��j��r�AMkcP'�zXKm�WX�p�k��,L�zE�`sr��P�瓪l�\��W}O�_5Yΐ��15F��Ϲ)]	�����/ J_v�j�7��R��t3�2���̨/k�.L�=b��N�v;�3kD[���ӗJ��`v�N2��2���g�w]"fǕ���U�m�TK��4��ȃ�TQEV�UPRST�U�5TbU�\�(-�5HDcb[�uÇO��==h��t�E#[c��DG+jN������NMQ�բ;.�[�ǧ�������p�*�"(�).�"��KcDALE;cF���R�٢"�(����Dm��8t������c���<��9�h֒*
��()���mm�(�+�0�:
��j#Z�S���������L�-��X�^�h�KEC\�S0h����AM3E4�Awb�#������;:i���ֆ�&<�MW6�)�s2Ts:y���m�ֶ4�U���.Ɉ���Xą'9Ǎ�U���f�HsF5�6�4k��1��lT&7Nr^G.s�q���V΃sr1�#\�n�"��%r�s�h�c�9^t���b��ۑZ9%3D���IMclŪo6�"*�\��Qs��1���9���ͫDX�;v�v��C�8wh��rB��w���Y��s\܊Z9b"Jy{�|��rh����gpŧ[hb�s9yh��w.LAM4UW	Ѷ4W783���Q�w�(�)���0���/�~u�v�4������"��5��n�yG�'� He	nl�B]��Q�Q�кE�Zy��`��b ���Φ~�5�_$�a�=����:��ioy����:�~��v^/b��d����i��oxi]-%���z����l�� �lȂB���!M�dZ5�}�y}'�&9�of+')��Ȑ��z�4��q�ȹ����J��ۙa�m�i}�`n)�:}��dgD�nX��|U� �S��q�-�.�]�W��)�*N�"&�V���w�uѓ�X�ʓBq�X�x����ՇTն˶���|+�l�_����z�J'�� �V^������J;�#��]=��n��e��l2��k3q�R͝OJ�w�n�K��Qج��ȥﭾ�����aȉ��!��7*k�j�ȭ�Mw�a��U����\���q	U�;^�kh�U��m����Ϫ��M�4�zo���v	ȋ��&:[OpT�g_��@�,M%+U��Qy/��~-���'�9��n���dj�96�m������38�Xќr�`�)��3۶�T�+�^�Գϰ��n>u�l�PLHؕĪ��]Xٚ��ZNwAdK/QV{�J̷��
�4N�Ĕo(܏���X<�ղPB��Ȗ�O���6��k�e�7kD%�!�wf?�{�VJ��b�n���v5 -.J��-6Um.��<�3�I�~ʾgʚ5�|z��]K=�-��Al�_+��}�Q��C��Go;5�)��sfw=��6N��),ᾬ�/�	�j��ƹ�|�*K�z4@������4�['w�r;wv��ҫ��sga7��ZȐ!v����e
B*.��J��|'�z糵��AIw,���,il����`��У�{U��1t2WW���5��1��������m��6������"؟o1��m��?-�D���$ۻ6�/�:�5ms�,�Ov5 s�dA��4�4�e�NEe�PU���_ӄ8��kS�:!Y�g�gs���Z|O`�G"�E^�,�i���.�X�Ņ�*zB;��Ьȃ�P�����q��c&�bބ���w��ޗ�X���)t��s� 5�J�f�Y���\D�mD�U��|�h)�|���+m�F6�۱�xt�������$@C��(�_l�;��[!7+@�H�R��7��'�7ձ�&ڴ�̼9n����ǳ��6����R�{�l�5x�}�A�t��]'j�:/��;��w`�0��0øoB�P�j�+��ᨰ�2��g�$oB���f�k��Sj���ojb�c����ݮ���AŎ�=�r<�U���	�A<��bSx���V�됞_$����A�!�V��a��|��U]	;gڡe�
�R����%nɸ0�]�wLU⡩>;?��������Z�r�k�d����d����*�k��qqewS�2<wZ�&3��[nσ-T�b
h�'u��c
���et,�53;�U�"%���R��U�NO۵>l��r���������TT�"E�l�6N�D�I4h�o\C����2�o�l*Ivvt;<�iɣ�g�V��e�d9�������]��ix��z�����.WϺQ��h�ɹe�������)��'�oVf9�����f�{��%�ޟ�|���:�É�}�����L���R#��Dr5<�oMP�Em���|�v�r�F�����c+E�e��}<s(��g/G��ܝ.�3&��(̙�9��٫o�v�N�b�(�R�x�ӕ�(mt���	��[���wu�M�)�jNy����`ɻ��6%�I�W'@�ܷ�&j�9�w�=Ǩ�k��.Ղ����xe4��'v�l����>�h1���=H��Pl��[�uf	u�E0��VX5�#�Ӿm��\�@�Rr�����9�&[��h{�^Ԯ���5�8�u�|��p�]���'�m�V��!���1�'��hw+�>HcN�֬�޿����n�7�_4 ORm�[����Yx�!e���C������������+T�9CړqH^{H���}��3��-8�K�X�4����ෞ�����^ɾ�>�o}Ӕ7���
U�~�_��G^EZ��Yc�5�,	N��~���������j�v�ho�u����Y�N^���ko����׍�z�g���-H������S���b���7[����-��ͤ����mԋ�\.�ic�ق�k�ީ�Ϳ1�J��]�����������s��H���٥Wʪ,=[���,�*��'�֕�?n¯�>���!��S�eD�i���y��5��7+m��`��W��?	���³3~��.�?��"�*|wYzdP�5�r��������y�Ev�V�{@s�:U���� ��rNy:�%��M�̖�9���W8��8����˫<W�Bk�,����I���t�7������1����<T�Kn�D��'�a��p�/\Z����$��D2���vyL��SS}m3rj��v�j����������Ƕӛ=;�j����RS���'��s�nu�/��-�s�~���t%��y����RS[�X���7{�t��i)�ڭF!-��6緘!���"�T����5�i��g3�=�<k������)=�}�ߴ���Š6%gz�T+��?��d{*������q����Fȓߗ�ݱ%���4���t��m�3-n[�ݛ�}x���N��_NH��lZ���G?aq�|-$�	*�i�:���c�V\u��0�Yx�f�d��!�x���:�OFn�����C]cبX��E��[o�/_n$m�F�l3�5L�f����7�@5�)���n���ي��ۅ��2�~�ϲ(�8/�����p�ņyp�J���<(�]��Q���J쓝�+y�P.�uB�X���rt��N���q�qזP�}���y�vs�+27V.r�n�T�u8-qz��ǩ��e���Q~zFc���;�~W~��M��9�;W"�jY%\�V��T��j3细�R�&�C��]�Dgb��r7d�}�;��~<��]��fUb�x�j��aL�r2�n�8S�k��8d\l�t%���B�����EfGK�
���f)�x�l���l���-T!�=�u��Ժ�t�*]�U�+<R��B����r������2�h��ꑫ#y�9##��{{b���YPjq?6�������U�����^�7����!�����Mz[\awS���c���!У�x�ތ�U�x�3�܏2�"�7���՜A�W�8��F�7�hx�Lݶ�_v�
�o:���0ng�v����|F�F�՟�{;�fx���S;��=�\�x�z�Ԅgd�m < �[K[Z".�e���س��v���u������틕��Փ}�U �#nΧz���Υ�FJU��S+���Q��ԣr:��d����_d�4�(N��Y}.n��-a�(������v�D�����f'N~�Y&KY�E4��U���t�4m�J�B�����tc���,�����B���ؤ\���/�KwĠs�-6#�Ҧ���3�)cn��U�3T��`�{�n�CE��0T#�a�v`�O#��Q{-�#�֭ڃ�n�oY��.+'��O�d�b5�|����u�2LF+�
9\�gk���.�kt�f7n�x�k��
�#ʗ4q⌃m@�qT����<�ҝ�k+8�t'���(E��O��hF�O���$�������5�݌��*���Z��9�g�_�BHd���S,�n똞�̷�E��ߥ7&gzP������E��u���_���*�oGWNLdNC}W�5C1�Լ'�`�7<|��\��ހ�
��-�,����U<M�N��~�op0�(|��s*��U�nyƚk�4W�Y��$�E;��rϐ�+�������?wr�0���~oޑH9��&��ئ8|�T�
�!<�:��V���ê_0�Y45�+a�t��t�]S�S��b��T�ᷞ�ꍍTUo\m 7yûQ��Ć��]yi���7��f�O�����Ǳ�|���<���9�'���O����h^�c]J�$������vT4�k��m�Gp��ᨒ�+�-��5ߋ��s�#����h$3=	����v�˲zdbG$���i�O��� �����e��9���A}z62`�*c��K	�������U^�%���.��:um-j��7ϨLVg�33���C��/Ff�BZ����v
++�5ԛݼ�x�<%��۩�a�����v`�-L�k����u�F�T{���zh�f;�����UOov�،��Ӑ���o0�
�="�RB��ʓ���S^Qm�{n�,l�}o�(m�@Ö�Xg���c�O��xM�e��v&�/wF�h{ <�u���f]���ר��~[d�g�,�޲���-���5G	��>�)���ff���Q��y�B4ʢzd��=/M�&>=G����>���{]�i�K�w����V�Ȍ��N"b]߅h�(g�i]e��T�����熴:�T���˰�5����\��f���1j��Rʇ��!B79^�a�y��]/\]�:k�ōG:4���ᘔy�����:\��W�2e����R���ַ9A���EL}�A���one3t�p�e�C%S��i�(
�����n!8���Z�_�:g#�#τV��wӿv�P��|j��`(b���.O�b4<b�����!���^��}y���)]^���J�����p��"ֺ��㼻K��sr3���ͳ��y���E[[*��ԮjϤ\ȭ��c�rϒ9Ѳs%��ڂ(�g�%�H��+������O�"k�����$���v�<ǝjO�v�q\Y�hrT�#��N�v��EC[��f�3}{���Gb0���<�0}[��pz�E���H�X�nwM�5A�l�ܸG�v���#3�;C5�	Y���WT��#*�>�VFD��g�ڞ姦7{�y�x����%�~c6�:��?DoM4�����w�&	�=����#��)v߂D����}�N/}^dF�ǉ��[��p��VNڡ�U�������I������u����&���J>����=��JS�> +C Y;��<k��%]-�Q;�������g>�|�)�ʹ���{�\vw#���%��'�m����G�H�3k���k�u5�ŷ�b��N���c@8�3zO�UӜx�W��ݲo�崓ϒ�i��#Kiֶ�RG5kS��u��8�/ݮm���&{v=��z�_9����%c���n"ķY#��Ζ��
&���(��������<ú�^�<��d�57~O��(m��m������`pt�i��r��ʜd����O�.a�V���_ޙ�e��<A#U�#-�g|�'SHv�.��MX`����2�s�{z�6q����4�"�qvdZ�}��a����c1����Q���goB��7z.0�܂�R�;f��)b�#�bq^4��Zr��������4��C"��E�^V�8�2���H���&�Y��Uo*ac��ڞW5U���d��cBFt�H����N�����w4��yZ�2��j{i��S���5�Y���\���/q��eo݃q��z@�i�6���vD�B��db^��Űm��.�����:C]˻+�{���}��8��H���XXR�ͷ%��;,��O���d@���T�����ut ]�}�rt�<l��S�m̲%�Q�W�W��ͭ�;�7�-�T��C��*l���K5��n��Ǝ��:pUZ\R��O����z�+��!����vV��`�m�ѭ]G���GL���LA>dVM'�c	�b&%Ѳ��ε��+��G��q�1�]|W��=	� �Nm6��^�՝cu�֬���{/#�]TVo%9WT[7@��`�ڕ�+!l�
��WŸ����s+�U����m��+6W&Nθ0
���3�]D͑J�V.Ï�tG_ly)�g�gQ~vs0��/�3qwD����T�57�y�>�F��)���{��&�s�޻n0QǊ�U&Z1>=���q\nk�s�u f�v����-�5`((2dv$y���6�1�`[V�A���o����v�y�y��^�7�ےa��+�����`Jg4���"�L��WQ`)d\���y�#;Fkft��/�����xM͡�e�X��]:fw`���E���;��s��6�ؙ]]t�sV��\�y8g�tso`Tn3�l+N���/�]"p��듫 �r©X&�9�������v�{��x�U�&u��y�z�q��Ң�.�m��Q�̹S+j���w�VIY������"wG%3!͐�m{�e0�]���e]����R�r����Db�e��,�z�rQ3������RZ��ofm�e^f���x�h�+�u���F�PQWDl��:[MC��7���E�]o���5��v`�)��8�`]��\��W�� �ΣO2�:[�#�^���g���Z�>�r�s��Փ]���1�d�t�tz�b����i�=J���*V��!�)X�H�luvj� X�k���}��J$�v���VɔQ�؝e�D
��9+0�'^�}�ak�_M8�#wp5g7�ś�cC#+;"�a��1t��W�j�P=w; �'x�������k��һԬi�uei��}�q��[�f�����N�fV�(۝G�ġ7Ay.o�r�})��ب���;n����|Ν�}��q�WW8�]-��^е�+��Z�Q��yPc�]>m��u�.�9�\+�RQ {�h�{�׎])E%�_�^��[�� J	�wt[����(�q��(�nkt�i{r�;�I����DoZ�%�ynG&��'�x\���\�l�d�e���׌\�:��Y�b�ƣ6�ӓqv����<�:���Į�m�n�P�f:���>ƹ��Y՝�olTd�6��J뉛*��Tc�k�����1���^���lH���*��oy���������f�D��tH 3G�(P)I�(�N�H:t�������F�*�9���EQݩ��MSTP]ػ�6�(֎N���ᓸ�F���#'m]�nETE<8t�����y���Eݤ����8���-(��NmTrLTm�8�`�Ψ���F���7�t�����gE���"���Fk@�j�*���`)��(�������*d=8zzzzEUT��5Tגj������V�w����U�"�*���5Ff���Q�:t�����{b
ӶtP�<��\��T1�EN��C˓���r6�U�ACDm�jƋgQlQgU4D4�E'(����+�PQ\��6�q�}����c:ti�m]��-�5Sj��N�=�vV���%�j�j	�cUG��-��ӣZtݹ�>A�8Eݢv�R�[rw�S��lUhѱ���m�T��M��Jֈ���Ѽ��
��m�L�^B�c��"��"�b�"m�V6����R �t�#�s�Ԭn�͝Ūv5,%\��<�Y�/p)�VF5��eA�Ń%:`��!2W�lYHdD]Nˆ��umWmsuȯ�8��{�j]���V��"4.^��C�3��o��j�O�����!v�6�z$�"X���M۱�l�a��Hw$e�R�8�Fd��_Q�3;nC,.��3�SǪ7!\A��Zy�v��i�֔*K�e�p[Kj��'̼����=��J3��!��������x0+&��Ո� �れ���W�LC���w���������0⟨�ʍ�;��/A8:����TJTն1�5��Y/S|{�.�9�����7wH�F`,9�4���vokٖ�[��uo;GӺ�lWޖ�.���P�x���?"�I�/L�g*�C2�Ϥdpx�7��7Ne�ae��X>J����@�lL�M|���ƻs����צcf� ��L���ݧ�-�+���,*��e����ۋ�kf���u9y�e�(6�.k�N*��
��<�b�2�V�	sL}�����^�8gdz����΍%Z�PR�[%1r���t�G�Ȱ{�bT�jdyA[G��ʼ��f]��2GT��L{H;�:���e��VwM[�0��E���A���U"�=�ciֶa����{(��@Nf���-�yx�CE��9�J?O��P*�0vR�)`�j��왣�'X<V)��s���8�K7C���9��Yx���p��<��a��f�yӘK�D��U��eP0�'2�H��k�BB�"uf�DվA��<�[���w�u}9��p9Y Q���2$����B���>3�u���y>b��n���I�Jq��[VVP��uC{X�R��l����V-[�c}�uo�׹����Ҹ���л�� �X0��2��`��U^J2/&��VT�����Z5Wļ�t�y.�o�1����zf��[�3+\R��9�-�l�5����oG�#"\o^���V�>�,��b`gt~��y?w���l��ki��އ��+��F��Q�Ʃڝֵmj4�zt����9�b�|�3�i��vXm4l������u���e�"��4�M�T8�
��t8�!��R>�s|��� ��ۦa��k@]5��\���I�npP��%/#���c[���+C|ws�v�,�k�!�N�;�c���_b�!yӂ;��i��\'_<S��n�����G�� ]zU(�n1��h��m�������A/fQ얐;���ZC���p�?,ەӒ׀�Ň�hl���b��!�"��m������a�I��n��K�;��!l}�]�};��5��]�:No�+��ۼ[��Fl@*�A�m��xTu�r�d��xd��;���tV��r3�}qͅ�U�J�C�������RۺL��e��s����=��=��X�*�=�k������b�E�ܵ�k�?e�[v\��j�������Ϊ� 9:*���NMJ)����h�v̚���YzM�̽Ekڒ��wUgH��C]Ƕ�<�p.j��&:i��1�d�C�;���)��d�I][޹��bE[I7�l��4�j�"&��a�`���,��ɨrFX�4zV�⺩�މ����ޖ����Y��c�T�g�u�]���%�7y*�4��2��XV�r�1�;Վ7[��s^��˶g���ex^4��Ky�ʀë�u���9���-�r�Lk�����%�g�a2��C|�#�艌Ŏlԛ*;�	H2X/oyϕ�s��\!�(h"��fѮ41+z�s�<��_A�Vd��S�^�}��:�cl���GO��-�2���3�W�K����{�X6�w�����}K���;�������֎��/s�z��w����s�wS^��f�|�xy��9'u_c�������X:��gq�^G�*�_�7�!Vuq��1=[9��b�K�戞���t�w���D�Ȉ[�c���}ұ&-�H���sѰr[vѲ{q�5��i�����s����������z���R������_��{���<�f��L41֩}|$���l7OxTyee�7���Df)b�}��u��%'�MsQܣ���}yu{5���bq6��6�saD���hi��PWA;�=�z,�:�ܡϪ��X�]�-�^D��BE��d��tzC��~Q��U>$���J�#e��̜�����@G:��W#�[I]���Ӝ�"�M'5g|5��x^��VT5_���6��:1��y�+�T�+]Z�SGV\m� ���Q���[���`Ⱦ/�9S����ϳ�ٱi�y���7:n�+9��R�i�@���KgV:�$�����D�z��F�Q�<{�\�	�oKYIJ�����=�V��4�sn��[@u����%bŎ3��W]����.���'����^w �[A��,�rdb�{p�cbM�['9/3xٽ�$u�Us�%�RqR���q&��R�f����]�;��o�O7~��o;�b0dq5/�g1�y�7��q�u ��T��tt̎���˖��ȯVL7q�Ss�{��4�}Z�s��(0�dk���Rݗ9=i��e8z�)lY]�*�\�u���0]�q����r���ۧ�����0�+̷6_ZA͹��5��1��j[��0�f$"mLl�fEi玲�w�D���mr16k�=��鰡���\m�g-�!}�u��,;�^�e��@� 9@��Qcma��8���g��wD�_ۑ��Z�f:��fR�>����Ud�����nh�rw0��`M^��c�H�A�}���<�DgzcA��e��X ]^s5x�����j����'w90J�ww���cGf��M��4Wfȱ�.���g˭��g�l�7CpYɔ��Cq�',�냯c��`��pkW֖g=�R��W���u�i����E��b�Qn5�ҔE�ޔ��`�3V'�.�R¥�ZI��ς��.1�3��"��U��2�)�z����	�*��V��:��G	3�R�˩�@x�k�隽�l��Y<4C����>xκ�̗��Z|Q�+*����.������~��*{����B]173m	�=��'(V#����j���Y��j���ws2լ��%R�3/#�h�}\���P�mQg,f���w�a�ѬZ���I�"s�[ɐ1�Q�yɻ�.���������>�m���6c��{;�0k':��m�T
ǁV�g�\i��)����j$�s�aW�֬�m�ʻHdq�~k�r�G��VH�Khr̉ �Ԁّ�)��X�Lɥ���GRD��G$8��t��ܑ6�V핱�+�+���t��&��v-[�R Ӕ��/�}��w�뫾��ʻ�o���WRF�7dn*fo;.$F�bIr���E�n㎅cnטM���>ޏ��v���;g�fC�c\o���������_	}��,±�[�9�9Hw^�%���s���R�=�e m7�����\��о���u�1��+&bԲ���.o)`χ��]� c��G���'���������UC3�z��R��6+0���L��b	m?|����7�ۛb􈄍<�۽7|��҄�p*NuR��w���r����A�9��:��` �A��؍d�-HQ@�l5��E���{0�f�`j�5�!�F��o�8@m2����N�3۽��m�}bǪ�:��g7���[���=R�ݧk�l�/A̋`�C	�~���N��aM۽tgG�\w]
P2��:����lD�,�T�ػf`��bh:���������ߌ,K�R"o�����w^)�r4)3�=�q<��C�ά����βE�ETUu���{�a/����u�5T�m]E���H�S��6#M�k2�!��rdC�h��d�����Lb��-��p}��0��(��	��6�@[���j��_xr��^T	S���7��V*�n=
C)n�&Ɖ��ܝ�����)�N�k��*�74p�:�����AC@裝w��+�:�½Ou((g�~�8�=1f�ɥ����+�BWV�˖��ob�珷f����G9.���+���c�T��&��x�_N���������xiU'�~����W�
��6�ot��3��ݙ�+Br{���Y��n㈍,����My���]���V�ʼ����������l��*��
h"�Wz�~���6����h FN��(�]�֒�� un�]���V�0��0��[Q�t��i��H�E녹�)��1�Į�5פ�Ǹ����7&��@wY"5oW�A"N'ْ�*f�7P�s��3u��@�>)c�@�M���3�[���\tUB�/���1u����^��We,�x�Iݵe�!-�8g@|��r7�S[C>=��jՉ���m^g}�DF@��P��{J�DeB`���s@��Z��!��#'o1r������Y����m�GM�w��W�����^��_�=�?v�8�6�k�0홀�ؾ�Y�s����ﾞ!`G�\��!����*�ۚͬ3�����p-���/6�]�N�Z�����k�;�D.��^G��!<�I`Վ�NB+���B������^:����̲:�D�V<4Q��������dA0^Af�*��v�Va��V��8S}�s��ڐ�)𿮁�[?D�Y��7#�pٷ�B�F�ByK��b,�/�7u�Ե�[&��f�o>[vWȽ�v�@���8�n�6�GCl `E�ƛ]��nǱ�����2s�����̚��b#��r*8���d{U3@�Qr6NzTd���2�sl�1ƭsgsNLI��wpq��!>����U#�z�;�R�a���*1,yz�6:���޻�6�Χ.�1�8k�P�AM(8M,�Ve.X��k�lEn���B!z��T.��5$���##g��]��IC]A�q�I�kiz���y�ុ�oH�=2#=&���kw|����6w���A��6g63�����:����㈝
v'���ݙ0@i��4�kV{ݣ��WJ"U߲�g�̓�x��}@q��k�A.d7Vϙ��>%Ͷ��idu�|��3W��p0����[�C�Xa��ӓ���8x��M������)r1C�X��q��ZT���ѯFC��Ky���^u���u{��M��í��
�1�Ԅ�s%k�j�𠌨�ck'��Ff2O'�9�7ӱ��fK��0���U{���*[�ҕ5��Ǫ�p�&t��J%��EZm��B��Z鲯���S��N�})�	n��a�����=�޼<A�;�-ǳ8�k��۲��DjU靏loU{��� �3�Qف��ts�!�+�4t!8E�X1�/Y�s?�0#lȹP>��k.��F�����
�	k���>�~���z��ξ������n�;�I�}v�)���w��ח���s�"�υ�����e�����װq�����pnTN��f���VVa�]���6����0@J����]�`ւ���U��ƫ�ޞP�,�}h�fK��m(���L���'B%�:����/2:kyctM��{<���E�WWf=|Bt�K����*�dLg���͌}��+�3n���=u]	�ĖW�P)�����mDt�
m�^�S�Odq9T2����v���}]��|��ᘱ7��7f�쩭���?�t�i8%3���`�+��᎖����Z�B�~h��b�� �yBw(&�Ƭ#���E�ƭ�M��w��M�Ok-�����	f:n�q{��aq�|;�K훏J5�)�F�q+^s�]9�gt���j�V�3�Ȩsw3�ide
�k���Nx/�u( �;l]�h�28��pmvű�Z���f��lYI�X���*-�h/�`�u���`��A� Y"�w=�#%)X��}!��u	�y�Vު��m�4���t�l1
'Yy)f�P�ˈM�������/P]����a���;��u��a߫�_@>:c�K�J�G����Ծ
R�W'G��h�"����r�M��B�\�a-�+�u�
1W��9ʝ�2�����h�b�	�Dc=��Z5�3�پ\3{�cܮ�+Y�-=��n<�W�G���5w`��njU�'/��2w>�w���:tFv;��H�3]mZ
�Gv���We�n���Y)kI�lfX#�V:�d�T���N��VXK`RX�ɼ�����b�� _P�J��{��]G(�P�����`��b���%qV'���c��;�������-�F^(t��aS7�9n��S0�T���q,)q�G�]�ܚ�}��!�U��;��y�����q���������օ	��A��e��VWp��p0�F�W�x5� ��3��_t��z>��	�O�\1�������6�mݝ��R���#�����;%8u���R�
T6c�a��H��ӂ'f_��IƂ�&����ZA�ΊR�<m�N��Ϊ2_c���"<u�q�ҏ�p��?��%�)�Oe=!\/gf��E�l�De).ƞ�v)�*j��[��
ua�(���b=�r 8Cwx�o	�POu֔��x:����u6�P`
�p�:���wf�{(�n���2u�Ӎ1�;Yo�pr]�������\w�f �L$tnb�}կS������w�ܳi�}��`�Ԭ�E���������w���P���wձ�5��G-\7*
����J��*�xm�t�.W�>�i�*��������r�P&�^���#�j��˱/e��2�G�D�6oh�7���ķc�KW,�Ƽ�^ �!�}2��J̻���	N�:l)iǂ�5�o<��6�9���"dQ�ޙ�W*.����Q��m�Y�.�:K��%5�]�gH�l��-��꾁����=pi˅]�s�����+m���P� u��Q/wv�\�{i�G�,�&w�L7%��<N-��8�0��j[r��.��֕A�Z��t�+�O^!o���uvJ�*ir��K�k@�������N�8.{���B�)�PѮ�|E��s.e#Z�T�Ap�pG2�#IY@Wm�'d,|ֽ�&�t�Y/�R�s��h��K��veZ��Kz�)�z�cqGwƸ�P��A̫�V{Ҥ�*�k\�wtő�� ����?-T�6cU���b#lMSTF��6�mEl�4X6ˈ����G��{�D�5Mm����j ���$�gO���Ag#������T�MT�^�3Uh�s����*���TE[5�(���c������퍵�j����S����DQ5kLM9�0EA8zzzxz^D�MA5E5Q{�EEMlj��ڊ**��b�[Z��ڍg�4�UD�m����`�*&.c5ˑ��43L�IQ�cs9ǆ�FƂ�`���{�-M�4�F�A��Rf�9sEm�7mE\�AQUU�ƹr�������D\ڙ��:�Eբ+���r8r5U�L6�E��l�PE��H��U��-�s��AZ4�#Q͝��:9͹��"
i�mQDD��$�	�ߪ�ꂱ�z�n���z���@�(27�KT�id#��{0=��>�)�»g���GU5�=j��J�����U���ʳŌX�iWS�ݟ��=c>�*��X�*�l���k�)���ež'�&ڡ��ѽ�+o].�Au׀��G+&��[��wuq�C=�\8Jj��5)9�]o�P�1M�p6�n�Ò%2��el����Ӗ��Ø��-3�6s$5/>� GR3%M���r�и�	%����w{���]��zD1��dܲΘs�!w����U]�ě���	�{��65;Z&��UU���;���J ��j�xb=ޱ-nf�Ў�ǇUy�s���b��I��^���j:�ׁ`@�������a�hfP�["fvwF����)n#ʊ�ؓ1��6�_��_fNrW}��UݯZ�#+�����;��g�+���s>�S��T<�^е�+t:���7!x�(��2$�p�q�� ��H�b*=}]��e1�s�!�S�ȸ0���K�����>���Ŋ�2��Pu�ݾi�ȱ�u-�7�9���,��Fu���w5W���.S��N���d1��;�7{�X;�˴*�B��N��w:�����s�V���Ԇ�7>�3z��Tۋl�տk���|ϰ֞!0�"f�Vu�����2��)�L�F��ȊSd��@���4�Si�<l5�{*bk��oda�QDMs�>n]�+��9�����m
2u[`yh}�y��R�jc���z*#D=C�×{�թbܑo�P{4w��{n��ݲT9;���^-c��?*����1��v�\�7^Ԓ�R����J�����uy}o�En�LN��T����|,V�4��pX�S�J\��jտ���ޓ�&�ߓ	:��w�<�����8�O�%�,�|[�$3�(���zϷ�5���UUF^kЭ�vvۡ���!�8�K,�o�Y,��Wh�5��x�M"(�n��x�=��;e�{k�8�W��P�t6�UK?@wX�����y�ب��b�=�z{�����ή	�c���:�VF��7dz.K�P(-�i!a�ۯv�0��o�L*f�����6=��*��`�+�� �oX/CgT�3�T�ˬ����e��R�A�
"z��z�4n��D�tT�ewN��.�xli'0���{��Z+v�i�+E\������K�caa� ���{d h|h��7����ѹd	F<���Y�;�,�Fp��f��qy1V�!ꥻ/�q���";d�����8���c(Z�ܭz����ZL��Kŕ�sb7�4O��� �k��m�ܨ������')���FA�x�%���8��n�;�� m�4��I26���ߠ@�;�nv����ja�gK�;�y�SUr+:���c�DƔ������?`E��*}b�{I<b:��,dB��T7h��綺lq�֍��m�{�5wH�S9�5
F�\{j�.*�{O0�~>�˷z���r!�d^)f�z�l�2w�9i@>�a�m��{�3<z�"T���)�ϯHO>�ג��V��$a4��5f{a5r���Д�M�2���"�����m�AJ~$�ʗ{����@��s�q)�~�RRU�i�zԪV��$�(���+F�/!�=yKAT7l�Cs�T,�xyK���֓��_����Iν�}o2�!�l�D���Ff�SۚSnR�t4f�9tx>��t`с�����iN��`o2���^D��(<E�sLݍ1�7\f�!�,eZux�jZ�D&�x�R�;����f<�zO�����K���T�%��;SQ�ᡱ;A%<�m�y#op�n�ճ�ucuQo�RU��	������f}d��[>����S�ۮ����n\i��VWt���s>g�}�W��!�>��'B��^اk/�g�@�������^��,��>^qW�y�$�_f`8c��v��U�z������>���Ll{l��V�~�J��r��·t�of�O���6޷��p�[�m�w�:��`�����v9+�hlmuEc�ؓ>����y�����,��6x7���":�ܭ}:2sE���f*�,=wy9W��W�6���ƃ���D��e����E���N&�Nb�;ot�l���C�ue�'<b�4�66:@q��2cL8_�S���+��WB��k��޼�V٬z���%la��{,�M`A��W�LK�i4�V�!�?wQ��]�Y��6q|{u͙xEQ~y�tQ�:����p�!��Wb|&VI�Ys��lN���d��֮57\��Y$��f���t��ޜ�������u,`���r�D�B��*W��R��0�G���'M4��w�t&�x�l�����32^}�Z
�s��bVͮ7Ze�U;��En��m4/�<`�4"�<\���ZU��!l��� \�UcZ޽����I�I��}l�q�|��g3a�T�f�ӪDǰ��j�7�����F��nx��Ȥ����������S#��]�v�+<��00�%��W2:7-]vp���k��⮇o�2vʜҳ*����Q�^K5�mq2# �M.���������v�ʀ}(ט�9~H�웟Oc}��ڭ��DM�(I{�����N�#�E�YH�;��"�yu�
f��%ua�=���{�9ƬOò�m��Y{!/�@c�7Ժ��ɀ��
n���%��(K*[��Nb�h��۲װ6�i���G�&�7gL9����Ƕ�K���҃pu{Vt{�7���Q�'��^�y�}�NHxJ�=�1�W����T%\2X�Nz��}����X�>f�z�e�B����`�2�%���]h��w�(��s��a��>^6Xз7pWI�*՚leō����sR�*u>�]$���кȲ���%�E���5;�/_�äW��!s{&鹕}�#�9U��ӏow3���9�~W�u��c�h�?��Y�����j����m̙���v��o��HO�y���>�ƶ|ft�n������nZ��-�0�2nwS2AW�|\
�.����/^W�Q��Ӧ(���C�A�ʙԞ�������%�S�__�#�]�}t�%��9cM_?S^7�r��.��񾵜����uf�o�{=ݗ��-�'8�^���Zչ��������S��=B<z��mZ6Y����ꩻ�X�h�MStN�s����[���s���χ)�^��<�4rΏ�^�~��w��t�������lf�݆=*����rI��Ê�n���_�ߥ�G���@)���ڠ�-]��Sb��Y�,"ԕV��H*�������++��<�o��5��� �Jy�L$�"�qZ�׃���d�M��Z��N>���n�Ni:t6��ܽʣ/�X���2`�o��sOC�I�;�G{�#b�l�s��1
X�\��8 [ϸt�2C��Yb|��r�gW$�+�se�[)t���ų��W�'����[�Z&g��وq:�Gp����6�pJ���P^n��ށP�m_^D�V�T��.lt��{�[=�cҠ<���DzĤ@�+��g���Į�R7��7q#��;�䶣�����,�Q�OW�J���b^���S�u�]�
Vj;@m���|#V�Z�Z/LS���L��s�ي�\��A�zGs}����en1���r3;�e7{���.f�OU�w7�%mnZ
O�^9�{�%��Ԇ���l�rl�(���9�7hM�f#5���Q�ܱY:�<! �s�LdT�ca�{58z*��ub/k}�� 2-�jU��}r�����@��&R�u�ӣ�U#*ʓ?y�#=X���Ge�S9�l3���˅f�v�-6��WJ�@5�Wn���S5:���&��
�ZC��m�� �]���v�1"���6��$+�F��Qz���T�Q�2��g�ph6�SR�Mt22��κv�f@��y��+<�1���ę��	�ӭɭW"�k������X&@�'y���Y�<�`Ю�,yBq��/�(Sӽ�f�ݝ|s�� �u�!�}JU�t)�;�WM�L��:��!]Mz��P��f����])��MI���|�A��j�2�x8���;�d�9�=n���߱���.1S1�ece���cq9���A	���M�3NȄf@��hZ&nE��{o�G��f}0^8,�a�>�y��Ww>�U�-j|��i�r�\�SEa�Я�Ԡ�QhsQ�Sa�g-�U�n���2����Am����W!�5ϒq��L�M]��N���~6�^�q�^��=B��Mڢ�f<��U>m#K�Ȥ��)���κ�8�1�UB�y����J�wX+���u!�E�L�U1sނ飡<�����/#g/�Pζ��y�q�sGR��Q��<�x;m�m���PA���<$�d��u�C��mӘ�Q~��P�J�A�i��U�g(�P%�qT��u�q$��v�ԧ�Ek�1���U|�~w����������q<Z��φ�0sx�-���Dou}���ƺ���NR���f�q�F�f*��i�Dǆk���M�{����Y�ݓ]c1
kQ�ì�����'�r]^��DxG���!=Y6��.5�2�x���;@��tT��R��B}էo�:�`W��K��.�����%�λ8�_Z�x��Qn��k���T��gem��~��!�1Fc�ϳ)N�|��e;�|򛳤�~��xH���7�f���{�ᅿ�wH�Fb9KkL�ik
�:�vs��QYۜ����_O�Od��!��69CA>mVs1�d���q�b�ȅ��0b���q�y�p7�# �)/.��tNiΛ9w���=U��"y�3�d]ʧ��V{3!�ۤ�b�����͍��X5e���xt�nSh~�k:7a� 5*�"�H����|����!8=5�$�Y�1���w�V��s��>}�*D�F�?/�WL�S�S���J�o�fb�z�i���xAU�R��W9Edڧ{S.��`��iR"��N��<����јٛ��j����e]�J�1�l�� �ʠV=[-���_���^;��SF�b��ks���i�-�g;�$�c��{�ND�YZ��$(��cdHkל�e�0lw��V�uû��k�HA��g��D\}yhH����/zL�G챨]<��Rŭ�!XӗV�QiZ؇�i:�|�2�ҴC:f>rdɌ�:hW=���a�V&I֗V�6�i:���9|y��1+��z�-ړ�g"U<�x+��/aw��ئ6�}�!�$�1��en5m�m�x�\�[���f�a�O>�}!� 9[>�4ϮQ�� m�����k��#��Q��X��}��fr��&��Y�<��x::��.3q�6ҭ����_n���j��[���rt��	�bacKd����a�f�-�r�V0��Λ1*��c{k3���ĭ\��Ve뷣�h쇤�߸OR�vM�F�12%��D�Q9���p���~V{�e�O,�,���	���0-�#�K=Bh�����D�m��"�H�h.j�ǲ��~f���߿n*�~���]����L'F��1	�-�/�v,��u���g(^Lʖ��M�ű;x,7�o���d>��˺�b&�VqweϼՀ�u��Mnmf��F��/��c[��9�\`EV�����������  *+��(
��/�?���P���������=�� "H��@BD��  	 BU�"`$TĈ&VUV@ �@� 
� ����U��  !U`!U`   @ �+�UV@ � *�	UX(! @((�  %Ua�@ ��!� �	�P(�H�@"� ���"(�%�"	A"
!��" �`�@6S�DQD 0J �QD(��4J �PQv  �z�U`$  EV ��    A !X	W`��!"K�:�o�AE�Ȣ
D���^o���?���ן����oo���O������?������?���i���?�����Ͻ���(���O�?������ 
���@QX����?���T��?�?'��*������c����p!������|��q����?���B� ��
%
��    R��( P���0 � ��� ��  JJ���P\!
� � � (   B� ���� )*�	  K  I  A *���~�,����?�EQhJ R��$��������G���_� ����M��ˇ�|^���'�?������� *+��������y��̠
���UW��A�o�E'��� *+�ß���?���'����������N�~�^G� �������~� ��~�a��{�>���������_�����` TW����� TW����|^4�~O����������������O��0|��@Q_�>_�?����?�������?G��9UE�ǯ�x�| Eu��~����?�� ?�b��L����	��� � ���fO� ā��|P � (�@:h(����(k@D�)@�
!
 ��@���PQEH*�h�	4��)� &�V[}:��Z�Sm��S)m�:��m#kQV�֭�ݪ�����llP�n�WlѬ��J�1[�WEd�CU�Q��6R5Tb�%l��F��gK�����EEM4͚�e���[6�֎�Z�&�J��Vͦ�Vմ)e�Қ�e��ٕl��fej%�Y��ikԍ���&�j%��N��U��,���  yT��X���V��mh(�J����)����m�V2ڕR�m�4XU����V3����-�[]i���43T���l
�R�9["�*���5������  ���P� z(6���=��C@ ^u�СB�
(P���w�
(P�{j�{8�Z�FY�Ҧʕ�7q�T�26���:[5��*mdh	�B�ѫJV�LH6����;-fl�^   ���Ԓ�g�h�-��k��M��U��X�TQKM��m���a�Ԯ��*�ی� �u�U��R�m�6QX٭�,S5-d4�0�mljCm��۲�5&��  ��V�
)d1��
VնU�4�[k+V���:S��Sa�Ф�9 �J���w@����Jm{�E@)��PQwje�R�[u�VJ�*��  ���P4�zwCD�u�U W��*�lL)�j���w@(gq�P*�	)��� Km�w[Klڍm]i@hփ �< ��%B�R.v.b���E(ݷw4]��5VT%��)B!8j�V�T�U�Тt�Ԃ����eURf�-X�
�Ū�Y�5� �[zhp ;u�*]2�X*�ږ�V�
 Vc"J�tV�QTU1a@
K��(��p  .魑�`Ҷ�*�;�\��a� g�  ��u� ��� ګ  c��  f� l�� 'We� Pm�4  :�  ԕWcRM�4��[�͞  ��  <rX  u�  �0  3+�� �m�4 %6  �` @���n� @�ֺ�j���6��hh<  ۯ  1X  w0 A��΃@ �u΀���  չ���� i` �7]ր  �~@e)R�	� "�)IT5 ��)�#R��a )�A�J��� 4 j�F$�  �I	⪓  Ԧ�&`V4 �I�h�,��Fsr�L�Z����,xXA,Rj�?�U}��_T���^�	 BI�!$���$I?�	 BI�`IFB�BC��������]�*Ԁ��z�k����v�i�]ep�j�Vsww�e3x0��'w1��
j�x��Q�45�]�dⷕ�;)�0�[yL%!�=*Z0اHW z�^������h��F���
���$���Y]Vckr��S�If���n�ɕ�q��@a�MVZi����I�4�oF^;�`M���'8�����˽�㋛g���pBv�H5��.�=Պ�u߶�&�JΖ��7j<ӢK�!/�4�Fk�{U�0�j����9��^fi:�,���*5�j���<�_vU/L�y��Jr2��U6��v�F��Z�1͖`}���ef�ްfv1��l�ػ
�gVwu��/ �z)gQ[������p[����B��z�k���w�V�8�����B��Ƕ3�//��Y�6蓚M�W��W&��kr��ۯAfҔɸ`]h^1�l�B��@�4�]:D��;a҄��1�$Wɉ�7_n�{�}�ͽ�VICAu��!�b��!�vu�E�L�-'8m]��N_,ۀp�ѭ܇�Y�_ݦ3����BX�Ö���R������y���jٻX?3����FƋ
�A'�n��7p�K�ڜ[!�鹼�fi崕�4ƾ���������ܮh�JF�$�o2X�V��{��8��o������j0^k������O�)t!@p���g%��Nv�D�j��r��T;㹹�5��v�F���1��[�����aڛ��z�/V.���X�j�wBE�9��-���9��Zx��O�p�A��b�m�[;�^u��a{�;���W&���!�����{��epV�Ó�t-���-bE"��ެ9G�ޱ��C(��W�ƭ�]GWp����7Ӟ��T�\9s��f���� S��	���i^�����p흋{�ǌ�D�t����I�;��v
I>�F��Xv鷻��v�z8��cz$ԭKh���K9�����/Y�y�>s����&�5�&�`��Tz�z���Fm�nXw��E��q�f��ӡ�݆�	G̯�0ׅ�͡d���S���os �Q�����b!\�	Ӹ�˘��3N5m>�cw�;о�	�|(tۅTJS���]��u��p��C�CQ��&����b�pߍn���-:��J:�o.���9��[)��w���Bҹ+1�N��V��j��p�b��W����q4�(epOC6@��P����'�L/����m��a|d���Ӵ��w�c��D��5L#|7��[(�}��,�)�]��,�2�٠�ň��n�<"��D�=��>�F�&�;���#ʃD[��(�郷����'J�:ӏy�����2Aĩ}׍uv�n^$�*�a
��Wy՚�b�:��s<u�PI���Kt����U�f/_3��_F8vz��Gè����"��;�<�è��kz�ϵ�B,�����ɸ~2{'^�j���Z�;˻��Pj�欣vwSģv�g�t�9���jflu� �Ej���2�Dc�D�V8�<׊(�,��#t�;�>YE�?Z���N���U��xC�<�\��$�����c7��y?��fYݏx%�ͻ���"T�c�\��Ӟ
Z���;5�kZ恛��tJ�o�]x���A�ʷ�6Q;�)4�5eB�4����
��2�s�x�J��X��CČ�ڃ�	ۣ�;A��7�I�Q#������B/�˘Y�z-T��*bzKEU]ћ��-�$Y����D��u,��Q�&�0�α������+)�����}oP��w/�slf��+o�lq�� �yEno`�G̐�F����Yظ]���C(n]�d��i���!��zp��P�`�f���ʾΘm�vU���m�+T�F�}8��N��}h��	��œy�֗r 6*ݰ1�39�$��4]��8`)�`Q��I��jߥSz�(R$���uH:�MG~�wwY�S���l�-�
��ǸQ�\6��Id_=�Nb�q�sNl�Lܸ�Q�[�j�F��1���i�֪ܜ�s7+_%�C�:f�Cj��gt�7Bdj�tH��D�U�7���t��8y��&��2�g��`=&rc�h˹�9�h��.���^�5ܱ�5j�H�t^?Q�e��s�ˎE��R�.�9�	({�K����Y�|�jѱ���+���/�J���!z�=o\���/5"��)ɕ��z��Y�,I*׹Vw��5Α&�ߠ�f��i��K��ga��rM����N���s�$,���@Ɇ>,u}Np��ʬ��ɀ\��mh:v5;���^�� ��9^��͟ �EВ2u!o6��>�7�ux�ќ�H�
}�@5����7�v�_#�YǪvD�U�����n�bv�*�Ղ��4�`�!��ɴ���4�U����5�f��:�u�@�ZY�7��Iq������T�Jf�,o�G�V5G��g I�s�[����C^��cLS��FkO��ܯERJ� ��JO'ߖ��ԑ!q4�P���bmg-��sGd�c{����v>�����˔�9a��
����3A%w���t�}�r�^���C3��G
$��/e�|7���GO�_l��R1kFe�麯��{I�ؖ.p8��U�M�X/��J��n�u��3�$�=�[H=��cn鹨���������a�wm��4�w��%�}G�����P��8�	����K�q�`<��	q�KO囎�<&:��wh��s��gRZz���`�u��e�Mu�t_fCcKoSX¸���1�7$�,z�� y��^G�W����K�G���BL�F������ޢ+0���8�+N/�C׋�h�����-krtbΓY.�E���܆F8,������wٌ;pk�'�i���^�'B���$���)��jQ�j{q-���oG!������l8���� +�v�2ˌ��ZԆ�	�8*]݃�X�X:���,a�|��~ �V�N�X��1�zv)�oJBF2��k�U����/R�
�$k�A�!��=�=�d׼j�f�C� �� Թ��T��Gg(q���S�ގ���ݹ��+����,<.�㕴�䲷�Dͤ"����wZ�&uW���l�8I�Ձ*l�+B95�.�.vL�v��ݲr vb�#Z �w94���dXf}k*�o�����L���7;"��\�3 e-k~���,2g�>�&V����$<�Zr�];"β�8���wV�KjE,bܲX�3�y~ۏ8�~��qh�#o�ؓ�]E.��U�z�K���,�+k|K$��t�ֆ*�tu��ysp&0>�Ӏ����(��[��r��$Ü���;h�oV����D]��Jn��IH�����:���q��ַq� �S/z��-��W#��x{��@���o8�#R�gU��+���]�j�򁺴��~���ª���m󥖊$۶]g���:�N�8e̓;-��GJZA��v�Yr�I�jo7�n��f����6l٣7�&7^�MP��}:�o<%R߻� �����gL���4����a�ƨWeo'�Esx�� �=n�\���Vu9�ʗ�@~3�;�u�G����7���&�=6�D2��<��eO��`�9��g46�k@޺�7�] ��˗0�7�plpY�+we�t3���bq!v��j��T�*f��K����l���zy��#4��#4f���B�n�)xA�IFm�N���9sh�-<���cH��-�t��3L:aR���}A_N�e�'�d+:-2աz-'�+�ӛE�cQim������Vv�Zx�d*=�&-]�c	^���8��!;����t��|� ;���|����jD�V�>/����C��q�u}��*�~	m���o`�F�&�~�vF��3X����n ��73CT9KsXt������M�����㠧6io��Ќ�U�&֜;�utl��L=8�}���X�ڔ���ht�9JK�լj�"���]�u m4;i[ꤛ=�S�2��^ˇ���7�B��K��K�e�nw��a����7��s��^ںe�n�E�� 8
IPMT��"���Y716(����O��1�����4�r�0s���Vq �-�־\@-�i���ͽ�{�1�Nfami��(W`��1A���]_�Jʳ�ǯD��R�<���l)��+IF�ɓ�^�1	��^�����@�ce�FJƚa����z�%Dao��tr�n�uio[��;sEYU���m.���s~��7m��J$�x��n�p�s���jCb�wN���^���˶�y��_QY�<ϷWkC��K�E: �}I�Opr[����k�0�K�<ޱjY���31�,�I��D��2�/)�4�ނ&O���)g'h�%f���7ܮ�M���;ywJ��[��f�Ý��N�R:j��^�Xi�Ŕn�F��:ã�(t�q��7H����.Z¼�J��X=t�6�]�A����S����-��[��z:�]���y�X�ҷ�2�q{�����dٝ����Z�s��(=U����nW4v�G��l%+L{�h7�]�y6�1���S9����,
�!�,f���a�wd�����Ŧ+I��K��6�%��W��`�y��E�M�v�����(�ռ��Z�ՠG�V���,���N(�!R�v���6�gV��U��ł�X9�KT8�U,�@�Z��4�uw�js��=�R)�V��{-R�7R�2�{�rK2�ҤU_YA�eށ�\Ő�R�@���e��L��י�|����+�1��.@�w�۳�+R�_"*�=�L��O����L�]ks�+C�26MpV��ea/�S��m���f8��)P*w��2L�����s/�j��%�hx]�I����vDG0dS��x]�^ƞE,u����/4�,�">�z(M�Kh�@�n��Ϋ<&v���Yi#ݪ� 1�����]t=]]���{Z�:������C$M��Clm��u��v��N�5h���4Һ�,��z!�94���|q0�s��q�VL?5A���v�+;��e����� ���@�{XK�·�e�U4�Ź��2�'pggur���-�0cnqӧ"��1�K.sPG��Y!�r����݆u�M����l��vs�t5j��Nl]����n�K͹ �滫Lu����jX7�81�8ү:j��D�"�9���Ǿ{�i�!w��a.�oH�wux�6�ӥK�<�b1��Ȝ��Y��&�Q�KV>��1��NP7X���j�NP�eY+ o���(��0�R?�mz� +���P�\�,���T(�w�Kp+��=�r.��tCpp�׵D���֙!�9�+z�d��x܎�;"}pk��c�x�ːe���93y`<��z}�U�C��db�ξ��V�D
��_�1p�Y�@l���WNq�ߢ�'s���|*H|�섛h\��P��,5vw)�ʹuuu��e���l�k���ǆٓ�콜��"S��}*k87N�
Z,��,�y��Yr���c�"��;y��I8L���&�\^n4z��z�8(�}��_�@4Į/�pgK���Qk���;s�X2Kn��n�iq���
n�� 0,�w��7�24đ�i�H�Qp���c��҆���烊��On�g���Һ�ơ�.㹏J����I���r�GV��lS$���+�-"�6N`��(�OnՁN�[I=w:�r���1�VB4v��ܩ���1.��oM�!!�7f�!�!z�"�S�1�O�i"�e��i`�P,��6A�A��6���M�6�z��e�}V�ň�sa�V'_ȣ�^C/��h>�w9��.�o��c�?gIYǬ���� ��Y��t�>�_�6ESjD7�����f���8���ss�90�ۖ[�V_m�Mrݽ��DAH�ԅwo.ѡ�aF�q�3YAf�ܭ�L�xG�;n40����F{�Jo*O�9�h�a�Yk�8��G�f�GIb@U3�YCT�.�{���C]���Ntڦ��X�\9
ܨ���� ����tM�
3�q�XG(KLt@
�At��M��Dؐ�s�:3�7:24;!�p���2�uդ�{ʬ,F�����&�fM��������R�ё`�wwp�bJu���4��zgVw<��+�.� (v�4��]���a��/aY��s2�:N)��th�.θ{W)�{�*q��x�������8��7�rl���f�6��/��y�{jտD(1Wl87��Si]�X~��i�wG�y`��|�����=�ނ*��x�ħ��nMjd`]�����e��w�=��tV���-Ҭ���J��6�^�SrpEa��A'����?�rJ��y1��]�V�'�i!R�+Us��j��"�R�%�t$�9�4  �=3e�P���A�Z0��
�����2Ż�R㋮�r.Yz�Yυ��4�Ǔ���5D��o�@���]�h|��_��]Ő���j���{��s�d�8�b8)AQ��^��N����ō"��9sb����%�Oo0'wQp�rNu��1P\4E����Qx�:�$;x0QF.$��,�A��L�;���Pg�έ���:����w��Rai22�$��%�9��ɳe��w��r�g@��`��M�C��#
0��\�T�Į���m|e�b J=��>�&��	2�C�wW�����{o�e�r���q��	\ ���잶N�da�)�0�oN���JAѐ�v\Kw� ��+����䯱<�	䨼
���T�R��^���
7F�������&.�m�ނ�s`��Û�o�y�Z��7���Q�Fٕ��m�}1�	�;�^d޼�]�he����SE������T�rj��Au���[oVq��y4����,p�T����v�;���	a$�B-β��V�v
X�Y���6�PXn�F�ࠌ��Ӧ�I��e��%n]^�2�7�v���~1��q:�-]}t	�<}�+�褡k*';c�����?m�Z�ͦ�{���#��C ��/NNc�����\!p��p޴�	����%��0v�ER=`��YO	��/��-ˑub:�܁���()�0���͖sp�_Nc|�?l�UR��ܸ+~�b�������(v[AT����۾��濻F>�E�n�����0Bpu���vsߧ�S}��-��V�+}�p�2�A�S�D:�q�֠鵴��+�����8��8S�3����҃���}�l��S3g��Ƀ|�5�{;�W��U�x��T	�tC_�o�]�Gr�=SO"����P��y�{2(�6�J�����޻��y�Z��?]+;F���s�=��-�S�{|��mm�rai���!�Ծ��AT��*�fv#՜��:_f����t�Edyǟ�*��Ή��:`�3ge���hݩ�k���B*��Daj���[�8��(���/K�p�o�.H+�ELY"�������M\�`���w7��S)3��v�l��[�#).�ҵ�7�h�oM�Q�R��*� �u��f�� �fga�N�sH�1ņΪΜDx ���A��������J�vM�V�9��d�-^�h�~���9k���%ʡ]��j�s.�յ�k7�Rˡw���P3ZÝ�EK��1BQܤS�ה͇�kAWcQ��f�XX�ӟgO�%���X��jҒ'U��h��/"s��nQ������~��1.'5=�hx'\[g���0��j�2Z�\O�A�b�ZB�VQM�X{V��oJ���f��i��^)6o����󵎮K�l�jT+�8��=���S�Q�Ѣ�W،�������2j,�F�Q�VA��Y4�^�����z�[�nr�c�0�X�ïLƫ^أa��5�i��P:v�u��E�㾵�u��r{��G���0�F��Bt���AX�[pfpYӶ�뤃�K���q_��7V}��T�,�n�]o�)E)Q`7�0�D�x�[5��p�Դ`��	9�����Q�]�pSx�Ve�K��SG�s=���C��TY	ӹN����;��*!���5���J{�����̙ý|�=}��X�f_b���|����D��7q[�x�t�ͨ�VN�A`�zNZ���hj�Za�:n��v(�{/$��r�>�<�3���������_Np�`������s3�x�W�q���C�k���#���,˼"e���.q�7�I�J�J�B';�{x�wEjU�PT���[��kC���oS�� �VuƓv��f+�=B�♽N(\ݠ�ř��"en.�:�X�0�[�n)}b��&P[�r��.^��Ļz���Шm'`�6�I��ɖ�ˮ7�T�x*AuL_]0�W3��q���}Ut3!Y������*�K��0���~�^ߣ2""������>q��h�Rp���nu�l��!���$�a�{k|������xj���pW`%TY´�����0[�y�1� i!�WZ�ݰ��e1�Q�j�G3�57�M�-t ���;D�?w�9���YN��|^�^�9#Ի7GI������gZ��i<���ۉ�w&���P�ތxkqvc�s�Ri�A۫*vn�W/��!�њJU�P�|
���-��e�ylyx�e�����p�g�G�e�ȄY�Ӧm�Q*�`�~��u��!�S�g�����D�r�7N�I]�Dfm�%B]3����ɯ�'d��+sb#�ʧm���ie���D���הId�+Y
��M��'ve,8~�uk{�uRI�rK܊�ܷk4�,ҀY��7�2uh@�1�IO�U�=�eX��eѕѓ�v��]^]�1�:�k�C�:#ˇ~��Kxe�k�)�k��a��&��k"�Sٝz�6��z��WǓ�9md��k���.��*[܃mKh�[�
�}om�(�zg��Y�z]�qn�5f4ǲ�{4�t��I�ږX���� �M/��n�����a8�F���f-2���6�wU5H*ɘ09� 73A�^������Gd����pV
�͵c����+�v��؛���7s]�iT��xI���Rp8���ju��3���Z��w[2�W�ՒvT�*� ��!�Sⷢw]��8���2v��R�ɗ\��R�%��HS4��J*�<1���qi����ww{/w��%JC���E�ne�̚A�+�KlC���..�K2ڐPr��fnb��1��3Q��޾������+��4���g]����ppg��E��*^�Q\� �9E��Ʊ�y�Uh��Ηơ��:�_;'��G{K�\f�m�m^K�Aխg&�T��]]*Ww7ed�*�J�����.�3���NŃk'A�J9��	-6��!��TU�n����5J�u͙҄�p;�Q�]�01�-�7qv׼&����{.���C�Z�N:4C�!��1�n��ʏeޟ.:b�h��ם�6�f���CGg���	��g���CjeЕ�i��2lԵs�̌4CG����.$��E�|�%؊/��s�B��Κ�i��f�Y�/�n�O:���Ŋ��C��� �^2:4��1���)�����.�N7|�Hu��՛����z�h�д���@`�X�Gi7a��c�^" $��*uJ���s�
(5xo,�uu	\���qMj�ig�;�@�-�%R���}�uB�ߗ�6�؅�-���������5�4��ˇ��Ă��@�Ә7l�%��SG.sX�V������[��+�Dt0mkY3���ٕ{@<W4^��tm:@���t�Xϯ+�ܴ���w�|�FF�Ӝ�y�s+r4+Yp�����Tt��W}�#V ���k���lTV���y�n����>���P�l��q��P,�X%�H�X1�g�F�y����E@l�)�Z��]�%��ݽ��h�{�˭=����9����AX�%�.X\����Q�r�s௣��؎���[\^eЬy7+MA\�:,h��IA�F��}�g����)��!��r���p�*] ���@����(��]��^�0U��5��qiУF��ӷ��J�b�����ZWq�k}|�pW/	�4��9�i�����M�fz�=TE�˽�۳��ea�ɑD(q�+px4����f�}�1�{ ����{7T������w�H3c�Ltq9F���X��C:��L��s��G]^�?��ux�^����Y��]�u��G�8a �m���z�^��S�����D�4����es"��z�ԡ����Sk�9�V{7;rc\]AP��*D>j�&*�v��چ�k�(��4W��J;l<�-����{8�$v��n�7�l���2h>�V�˧�-�k��<%�F���L�J�A�e���)Z2á��y�}����^D$h��N^��oy;G�u�*��g�9���3��5��0�;�,�W�����Df�F%�r��i�+y�`Ѥ����uf�!�^���ݧ�w��ѩT������b���/z�TՎ��<&�k�ST.ƗMBuf[���:��`R�B���1��S��[��p��S6�t��j��X.���������)�0<7A����H蓓3OO����M�U�9	��G�޲G��;���ehvZn�1�K�]>Z��q�od���d9������F�^:Ĭ��}�����eȕ��uM�M!�źrK�#(�����C�U�!m�F�u�+�%���6,�m����W`6�z�]�=���y2��
L{p�6���q��EEwj�b��}W3��t�h[[Zj�˹1�¦�VÂ����[w�Q�㚚��.v�b:�U�R� )�	���7���1��5������U��GJ��s�S�3�4g���ݗz�۾l�؝�L��I7	b��oF�{�^YC�3��K{�ܖs�#@10�2)��son�2�ݞ�jKHUU����}�/����hXں��
����f��Ss���9}��Fn�����m90����rwm�[�oSrqvKTu>h��/s5��Ԭ�+��H�3i�������
�8��r����7S��~jq'����g&r"�S�uG�����yٴwEڶvw<a^���Խ�W�SW֭gy����
�OyH�儕�z\��"0^I�;f�M���
�0.8rgR)�d����I ]�p֯W����o"��S�zݬɳ+6o��r�6mѐf����=�h�Ok;�Z�Űz��b�o\�d����k���`�u�Du
��r���A�rR�Ǵ�n�@T��T;�6vf9!�,F/5F��{Ǹ��+'���pH��8��=Y���N���2��x�j
v��5��F����do'i���0��03���ʫj2��Y:�&o!��Aj,�����5l��I@���.B��3��U�ϟs�ߜxi4��y'K����C������tA��"��7���h��i�j�Qו��P��+�u�D$���6��F��7�R�!��-A�E_\j��	��^������j�
�J�i���F��-Ε�A���y���S��Օ�����SZ�.T~,�`궵ʑ*�"�P��{7~�N	��S5�%�kh�$G�o�Znl�6�6�i��#�Q���v]�\�LLy]8�=�g��-/ʦ��So�a4�s�J:pu	�5��5�	��Cs0j�.�c;l�h��R!�ŽPfg��͂�%�׫�r�1�6�U���Ѩe�7: �V�=`IB-��+�
Zb�����`ߚ�^��)��{1�s���l}���-x-�(Ӱc�~]�9B<��7Y�}���@;��k7:�.���1Sڈ���w�W.Ҷ�1���*��qc`�ɛ�����ͷ��$� �a�ZR�i��mk&�5d�g�˖�;�Θњf*T�A)�4U E���]��R3(!\7�V�3�X�C�����BҺoUJ[G::���֍t�
�n�s�O�,��)۠o,Nͮ�ܬ�����Pf�Z���De�Ѿ6�/�fq&�V�Ԣ7Og[�f���1�����Z�a��X[ %e�{k�v�,�M��k�D�f
� ��k��+뺁`6L����p�i��M�Y/��:�ǣ�j�~�����w�O=���0wPWr8U�I����K>X���3^]%�٨-5���ܶy�D ��E�����y�2�{��%�R�t�7¬�Y���R�ƅ�����ؐ���2bve�r^���f�]㥹��`R�]y�P�$Z#�CF��M;�)�krQ��8��R�,�[�=�2뻝;�}(���|7�o"��|���YN�%g�W{pH�:{q̎g:�a�K�}N� ��q��}�V�I�ִ�)\Fޜ$;q���:ACY�%P�2�o��#�L.��T�^�5�ɡd����[jTI��9�'^BO0�t��u+N�ѥZ7*R]i�y6�ʵd�Y��b&��]��L	�پy�{�|���[^ �y�ʻ}��#[�N�8�պgX�ȶ^�!k�f��e��2L���k+���=K�"���{C$��g2��}m̽���̀Ң
q�%����Z�#�Cu�C��՛��A����@��+NMW����o�ǔ��+^H��1}{�X��݋<4����K`Je+u�L�+�r{V��xE�kW�,���ҟ���us��8�*�R�ƣ��f��N��{kkg5�u�����S�ʳij���
�����j�+�^��a��w�V.�ɿU���h�Gnu�G�cU0<ht���>&�ڥz�^�������{��[���Xok	Q�΄7+!ǚp8��勗n�I+!�zv�`��H�'&91*Lyb���ᗓ��wfu��Jn�V�2�΃P�E��;�y�0#��r��V.7'm�'B���/�%�J�|��e���l�H�u�	�Ww����Ƿ��^ŵ+p����2�Yf�L�ɏU�E
�7���}��۾���g��c�zX�J��_ě��(���^"e��{ah�egb�O&���+Ey}7�O"ͰI�sC�/�|en��Lw��p�\�Η�rb�X���BۘeY��t\Cxnw��f�ڬ���eװO��e�u�r��8�4����E�z��{mk��t�9�2��뷽��;:�����b��d��҃WrM��a�*�h��^��g�O����'�/��&�!��
I��o_a����]ީ�	��733  qF�WV;�3�HH�K���gɽ���D{oq����q�YQ;G��;AZ��ԳD�+�k�c��}�M���5׫�����:�H�l��5u������$K�x�i=I����SM��fuq܉�>u5�O��O�i��7qŌ�.�3�/"���(�5�k"̦3f��\��JS$�t�,� B�����O)�~�]���?k�~���$!$���G���D}}�p'vC���&{��={�Ѻb^���&`��v��J諍�Z�w!�9n�<ܱ�,^�Kت�y�����w�ڥ�qe�<�p�j���V�[ڄ�r��m�GF��h
���b�{�S��-"Հv� ����M��)�_K*�ǷGx������^/X�e~Q�.z��nMs��!:�C	��\��Ѹ��9��SP�RX-�e8����vz_�&�3䆌�ڍ�p;�iT�ù�V�59%lt	u|��U�'b=�.fp��Uʆ�}:cS��8�X���v�kELt�nD���^٬bNp��RǕ|���4W�@�왎��\,���2��)�Ayzԅw�Ooot	xc9G�{n�ov[;����wπ¼��	3ZK?)t���0����5�anT�ݬ��@��Lļ ��L��E����[�/�ʾ�𧂄|0�����@�GU����հ]�hw-@��3+�!j�L���p����V�ͮ�vS);��v"�R��]tG.��я��[6� �ۺ/]�]c�J�k��wu@��Zo���_`�g��e��7����O'O/z��2v3t����+:��L��x`�a�aj�EzW;������{��·ΰ��3���^�<l�x��3�,����V��F�ZvM���gE��37����
��O#�&[ՊFF��<�J�7u<*W�o#���ԃ������<X�T߅��	�Ձ<��SƯ�g@���x����FJ�Ȼ�4�fκ��x�^R	n8�l��Ρu��ŷG:^K�I>/5�r�mY� u"ɰݑ�j��;pX���HmI�E������ʆ���\,2c�e
�tJ5�K�*�ԕ;�.�i.�˴.�i��P�Pal�8,�y[u
+��ێ��S&�u�OK#4ɷ+)D0���³!/_qݧq�b�w��dL䋤�;�7z5�WA"\��(��YX��ӏ�/k7Q�[�����V��������e���+{��Rʌ��$��_x�=�ᢘ�δ��}r�V�Q�@k�n�	�<yt���X�Fj���c��1K�vj"4�5sC7xF]��PP�z�N�ܙ��Fj�����Sv�������0]J�Y:�9g$�W)01�Xs���I��OF}�G,�.k��cF>��Lg�U�|;�T�ޙ-o-+V�G��[f��=�
s���
`��]���p���F��H�w�U�A�ո�Q����Mٍ\�Ǩ.�E:\feڼ�軅H���Q^|���[���CuA�>�[�ː�f����5d
�sh�F6*'33-9���o�|��7L*�ו��kS&���1m��*hR�rIN�ae�C�o#�@�u��B����
�V7�˝ǵ��W�݊��^��I��2\V��#˝����5w��}}�%���7V����=�+F���p��[�=���˔X�y�g��&�6�\Љ>�U���e_��gq�c����B�{����z�è�T�:�
I%�X�V[�o6"t���GMܕ+����n>���2�	��k
�����X}Qx��l�FB��9y*!Or'��1�w�Uu�f��D��x�+c�e�,G)U�e�N���a�ʆ�K}�]idZ��jQ}�x�Z�}��ޚ�n>���BL�_"��hJ\�Gd�m!a~��-~7�u�pT��%�̎b�䮚m��L��au�q:w��7,ϏkMPj	��jx����t	S���/9��6�Gn��9�hl`���,�y���*���i�C%sp���{Jd�A��8�]�F��Wѥ���� W�߆�op�Iڇ3W���8I��}2}����X�*[N\%�N��.K��b���G��'Q:>��Qͩ֠�><;[����'F!݉�:�\#�a�Y�S��-v�4�����t.���ر��c�M���c:������!�4�������㩾��=C�5/2����)f"x���-o�zQ2�T�-Qv]k�Ԟ (��^f,���&�&	��d�ܒ��w�����W�r���ё����5q��z�2WS�G9��x��Oz<f#��1�A��M�KE�G�`�+b�D9ʆ��	䑌T���'7LmId�yʤ��f��X�c�=ެ9S)���]�	Zcel��v���4�4�j{�ŕn^z�U�)�q�����ƽ��w�Ѐb�����P
��.������p^�s��Cl��:l���̬(<v�Z�Ϥ��ֱ6�Qc-4C�7UXz�YD��t�erM���$�Ej�eÖ.u�1L�ۂ�a5ڲ��e����f����'Pιw��ʒ�+�9*�$,0z,�x��+p)��p��A�|0jӽ	��#�EE۱:]'���`�Sb�+��]��ټWo{������_,X�-����|�T���$�<.���E��>��`�\sGņ"��
1��0�Y@�̚5�D���˕��7��vQO_{����D^9�hي��b��ۙ�<�ij!E�(m���ӔI�a�`��ZUv�jV�r��U�|DN�e�j��̇⢼R�+����[c}�kl��V�"eve�[
//�4-�����;�n�Z�ݰ��WRbwP�$v�J�/�]!�K�b-�K�4�YMˉ:٢�������}�]r��ZaLCi��b��P���r�\��˥VΨ��p�*ބ�t���-V;��$yV��*�u��0n����X3e���^
[J�:����jצ��M��#�^�u���*G|�[�q�������b�	�w�\K>���G�H��z�#�@��f�X,�j!��Vi�S���.���3�V@F���@Ȩ�����C�׬���H��ra�ِ�5�v��[w�ojr���×NR��ZN�c�W��ÅK�N鼭�0ux�i����#.-(��>�0��T�jE�#��g"<��B`�Z�n56�ucu����E�,s������q�$����4`2��X��'b���촽ӶU���X����H��ۈŁV��m�N4��R��J��fq�������+]ҋ+�����qY�θ�r.��k�h���#�3��K�5E�NiŻ��o@q�Ѹf��7tk&SK���)���O\�w+-�P4��2���Y���0>t]�.�B. �ٙ[��T1��T���}&�� ��{qɝ��
�3�U�mų�]�]�Ǝ��>�	W�XZV���yfv���uI�Wp>'C2�[7�����NCa����G�	w��q�}4k�s��9�
�{"vR���^l�0�\�(�ge�1F�N�w�%�����B��qgu5v�K0��#w5m����$�X]�T�����<�� 5٧0��"���,#���(>�:��V��S��γ�����1n�l�j|^�ray�(��N�X�]G��\2��@�J����h� �bޙ49v����RS]#N	W��En-z2�q�a�M@���x�` �G�t�}�)�:�0�W�o3o���
�Cm\d���s+S���f�˙{�w�yk�L�O֐��]�e�yb�}u{;}�]c�b!�!�8Q�f:�������A�FZ��7���.�d�!X9��-��WN�����w{��V����⼟���&b�d7���y����yG]vu�@d��%8;�T��L�qs^w�vN&󥪺 �U�5���	�6m����O;4��IyV��+IY�W�d�N�U�&ݡ4Y� oy��
w+�B�S������Z�7��fq���B�c���a�.�פb�!śj���70gK�c��	GN2k8Fz7:�R�2v!!������/�Q{��
Siy0���7�͠�[ۺٛ�×-c@.�0iw�?t4w����q⩱����,�����Y�����[��l���x#�y�ĈWDN�RӸs�c�Q��&��X�Z�������s��>��s�1%|{"<p?�
C�vr��"��=�Ь�.-���j$�\�&��,�{[��i䦄{kq�C�'�Nk��k�&�NE���Kz�.�S�$v@4Z�w=�J�k/jr�dc�N��Ւ�����)Fzi�ٻ9ow rC��B ��y'.쫷,��=D�UkO)�t*����P[�q������Μ�|e���LY�1���	���ga1f�^�:8^�<<N�����]\�Rj�S��β����e��`ʻI=�\C�n�Vc\������ԲBT�$�5�Z*�obwmY���rg����	z���oR��ظ��� ���8{ͱn:�0�B�|':� R{���G�����l��UKyW��E\^׸���6�j�W<��z)U�;��Ts���z�
��x:՗o��8�X:n�XL���+�f���I�b2X4�D��8�Ư�y�ل�t���Z��Wch٣���Rj(m��)�s�X��ʈDgJϙ�6��Xodn῅�;R�ӑXƚ����o��z�f��\GhCg�wġ��d�;��7���*U�HƖ��0uՀ.��b^9{�	z��M;47ĝ��nkxM	�9B��h1��2��*gP���
j��v��N��މÚs�����h?�y�e����B�����o�����{�3���ý�tY˭�-#WU���Ū�s���rك����ý�y�%�l)4s06pNff��r^W\t;�%m�0�df�f�߶�M��a1�д���-��n�N�Z�U��Ê
�f=�����z��n��0�`���B��ӯ���E��0:�*xݸ��v�A��eq��vda����`��k����嗮�
cB�-j���9�:�By�W3��S�2;_í�y�������x�'��-8�k��w(�Ǳ��V�a~ܪq��t�{냆��jȑ&�/`/¾~�Ln3³�����Z�,��wg��fѬݫ�u�rJ#6��L�7Obĸ����I=�n:TgTli��`�`�>N��-��@!@^�K��d��؁�7���6�gbb:��]���V;#��+ZѮ�h>z�),��k3��3hR�H��,_iǭ�"��$�Ae���������M�ǳ4f�.+�YY�[]���[f�!�V����Z���7������T`Ơ�,t��?kZO����ۗ沖��8Ѓ�=���,���u�.��:/2}�A>O��-���*3��f��X�?�V�t�yY#���yB�oP\�NV׎��%���Zr����{&޸�() �uu%ڭ��kK:�}Ҟ�1��B�r�oq� �%bm�a��IR���r�!*���m�vU0oY�F�T��h��C��Ow�,#p��.�t^>4�a����J��̈.ˠ�őK�jtt�дk;��al�L�1��u�c�-P2�ky=����1. �tE�*��{5g*�3��-�+Wd��S��oPo��Sb�^=���Tri�J8\]�Ս��z�������7�j��L�y:�*�s���dݔ:f7�q�QM��[����@`�]iψ��g`��#��fpn�����2���l��{E�U�I�k��&6���}qܩI��
 0���+L����zv2��6r�Ɋ��эŵ][pg%�k�J�)һ����0`�� y����px�����;�|�R�Y�7�qn�4��U��o��2�^uFh��jy��d#��㡫7On8�vxi�Q�������9T����5t� 6С���c���..3�c���9S9q�6�T0䦵�4q+]���V�0��퍊/��n01Y�r���Sa]S%rF=�X6í�V��y��ȟbw�+P��#��m3�W6'�!�m^>��wY�$4��0Ƙq8���5�Eڧ�@'�A�?sYr���2z����7���^�5�EC6=�Ɩ��7�R�Pۚ{�KUKAсU��ʼ�w����I$E�F������[Ŕp���ہ�70�mD&X/0�.��;�$�{Fm�a o�;���cIu��5ԓ�g5�!*������ɻz��|���4�B����䇕3�{��F���/��5��6&.U\�g�]g�+y^��	;F��0q�N-i���o�0�#Xۛ�F��r7��f��_cҌ�n��vu�kU��ctȁ�M�8"�`��k0x2�N�]KÛ�N�[XG"�K
V��G� !���k��:Ֆþ�<���������$ޫ�,ჸt���K�o*ܬ%��2oQ�+6��(���]˂\�����%�n�)��37i������vK�[!}[1�dl;��RABc�V�Y�ND��ފ���R̭��p���О�dgd��W���8��岆5yxkt�qp(H�i���&^qe��KC��NH�y�hT����J�q��	}a2YБ����܅�U�������˼<V`�v����+J�&���p�YYɅ�<쎻��O������n6C�Aj��C��f�l����e�e'�h�.��yJ�a]���M��/{��u���{�=Xb�^�]��k�ƌ_e܎�0 �X�]Ae����.��5g���FM�F�vr��x���	M񽇴m�ğ�vMΙ����-��V^�\��r�-F���ū�&^��l4�OP�W@���9[{�c��R�o�]��^ ��4����vV|r?v��d���*����qN6nr����{B�7)�)e�3%N��.Xj8Y����aN���g;�s�:�n�m\:��u.�k�k3J�E��yƝ��҆C��$�9@�uã��o���׼*lT��}U��D}}�V����1���9�{�:$q�]���ݰ��;�W]xx;�נ큰��d�A�}�Ima����Eە���5�,����V�.�)�f�wu�#˴itv�
0�BtR����g�~	&zL}p�r��=j�xw�L����p�Ղ;qoxW�ߞ���77�,���-l���hxӜ}.c�.���lZEk8r�&�Es*�{Jy�I4���4U�pM`)�y�7n�Li�����ܙ]�X�s{������ye������S�O:�c���IX��yCMϒ6�ƣu�E+-��^�k7;<�e%vt�p���Epݽj�T\P���Ǻ9n������z�H��o�>�-��&:�Cvi��8<Ьm����w5�qn����Vn;t�ic1�l<�BÔ���W:���*HMT����h,�ë�K]�K���Ҥ���f2$VJ�/0�`��[k2}�s%��I�]#5��3D�LV3������E�ڋ�9���1���fǧ]LB��'Xv��,�wș�dl盺�I�T�p\�c��כpZ"�N<��+�:�z��dc��e��,�����l'|j�-�ҫZ���'��{=��K���Eh�ww���|�@*%eqݼ�S@yZ����J�ލ�çDc��j=h�0j��⋞o]@W�B��h�
�;�L���M}�R�;;T�|�9�j]h�Wo^A�b�Í(���DPU�F*���#"��PX�B�H����`�V"�%e���0V*DT`�2T����*���Y���YR�²���A���#�Řʢ(�TDFED-��`��V �*��V�Q*(�X"V�1*+�0�E�UT+W3!�m����`�Rج�������UT�UU��Q�cDL��*���*��9Lp2�e�QDQUUG �"�1\pUU��(���"�e̘3)Ue�����*�#���V**�(�"��AkUY�TUks3��L�TUr�Q�""����b�`��*)F1E�11�UX�b,"(��Z�Ub*,2���֡X1V+�*���*9J��0�%aQX�b�"�6
��*�+�U�jTe�"<����ٴ����;f�3bN~�S�=:y����]���Www[c�/&<�jW����ٱ{7���h����Y wN���Pn��\)�v���S�T V9�`�9�֗zlL�gp �.�������̯��x��~z�����R E���Ȉ;�f���9!�ܶʭ�h��qn��������+Ab0Ro}x���x��(4��-~�~�(髁;4��&��̿���b��k���p��@u�'Ê_Ƴizn�zrN�ç�e0�h��x��*�k!�����s���U����L_1=���q;��-�2.Zx
��-O��h�p� C؍�@TGLZrE�7�h@�N�u�W�+�M��<XW��;�@���ݒ.�����+8*;��7H�+�O,}p��&��wr9�{S@F��!��Z��wY��k�}_]�ㄡgV���%�ά�x�׏���t5�q�m�Xc�	�{<KԜ���|������x�;��@��b��,%c��&c���p�5ؔ^	ٻ�,-c]Γ�(:�n[)�1����U@G��@.-j�L�#�X���t�:���/�/Q��R�T�ufT�c+CR�e�v�L�#������/�����uK���&�ߟ��+��{���8BU3^�
��K��d�Ua�̝��Q(tA��S;�}��Br\DH�jR�������&�l]Ňpbr��R�d;���ת�q���������B=�2�����;&���� o\��7G��Rn�9��d�8a.,�9�]DE':$o�5_τ��s d�o!�=�o��d����������鞓
T����=����)�I�*I����{�ɕ�p,�P+�n���PU��F!#?WM
+i�#��W�Si\U˨�v�D4��f����>o\��B�`7��}| ��1��B.F҃�3F?����9���8L,"��Y@E1�S5������5�P�ٛE�Q; u}��.�ʀ�誜r�V�W�Dtk����'�f=}3���c�ג�W��)RT��&~zT���$�9rV��1�k骅�L�:�_P�%e��0#�R�I��LOݲÿ������S�j��v�o�`ŀ����y^	�K+%���<K�=T���r�v�*�^�h*ֈ ڮ�a�S6��`nbD����MF���8����چ?�^��cxUj�o�}_U��
ٸݴ ������4ԧb����\ڶ�z0���]Μ땫����/��&�z:K�xB��k��.��Z_��왻Vl�n>phɌ�����r�̄�A
�t��o>�d4��Ʋ;a�7h�^�%��ª����D�Q��W��7F��_5� �8����r����7u�W�f+����yջЪ�*�V��^�H?�u�����~7T�A�X���A��[T}��M��B$�!xq�$u���s��U�����۟*�	�w�p}��:��3������'<��X��V��5��J�L܄a���.!�l{=�d�e�<`�/.ׂ�]7�[4^!Ԁ;����l�_K��կWK�1C�J�{�6��阐�gSg��6��OuF\7�,��#��wnԼ�
q��F��T����<NAt,���M4XϺe��8��	���VW�� ɣ���<��EX�m��}�T�}�K϶Ny���V�ˮ!
��}p���8T)�LnͣǢ��[����^�͠4;ۨ�4�_@!t��F*\�$x�\^櫀����뽾��yp5K�S�do�ٽ�4���8�-]��B�@Kf�`��.bD�/�_��6�N(r�NK����������TI}NOC1�8'36S�@�n#	�F�ƩWy�V��W�O���ǫ�TR]к��,ppzw[0�Trv�*���<�m��uCypVK���#!�k�fK|S�(r_tt�W��۸�͌Ԫ�喫gGK��a��+(M���	Qu���Hd��][f���	��P���i�5�� 2�m֣PJ�[Q_�F���m�m�_Éɖ��Xc�ة��ct��6��,�ғ�Y�!GhJ��/�LV�Č�,n�J�ܹ�3��О��G �9�#�d�����-�y���W�m���XƎ��Q�����5�sK��	Y�/�dB���6���Y��uoM����4?�� mG[�+�2Z#4[�
)uAEw�
Ǵ�d�f��Y��}9=���ל��Y5�Y�?pN��r���B�e����^V<��=W��?rT��<��wg��N�P1�*3��%�r4�?g<����62�)�ɡ�y,�V�9��=��tr/���q=���0�tE9�(N�Ǿ0V�6VW|���ܗ^{ԗV\��Uk)D�=��0�{5�ɘ�P1�1_ڞX�]L@ܼ1(�Ğ�Ȏ}{2�ڬ�my�y)z#h���۴���Qb�gy[w򸍔(F^)v��cE���#�:��l��<�M��{���>���Arh��]'��u.�t1ͻ��D*j�������GX�ܬ��ͿE�F�1ko�m�����hV�D�Eh�l���)՞�_�S������Z�;ov��Ѻ:����Jm{�]���>g�h`�-$^�����y�.n�(T3���x�-Vk|�oS=�G�ܩ��[�����vfT��W4�זiV�,@�JKhm��D�b�ǒ����{����u)�^2P�,y�<�)E9,�G�L}=������!�i�{jQX���7��w@"�S��m���Bq$��y�pv�p��E��4���d4&r h���ܺ<)���-�NLNɻA"�R�݄\����Gp��b�1S
���9����{_�{�묻�R�F����1�c�m̽NE�h��U�M*gG����X�kW#���_3a��	ހ���{-(�Yv�����B�� �!�Oq�@Zi��r��n�L!	3X.�L��� NӺ������*��1�Ma�*Ӣ Tc��3�W�����nw�"�v
�iX#��l�ؼ�V�"� I�*��Z�s����ϫ�L�r��,F���gו�fD�E�T3�5\c.�F���_��g���F+Q�p����v���ԕ�*²`ɵ���!Ֆ�:�a�)b�<��S�u [�����]h���4���[{s�9��^�˪l�\��<�Ǝ��X�����
��p\�����`�׷�w�-�Nq�u���un��*�`<u��x�s��mʺ�4İvl�1����XXt]�%�2.i��=uٳ�Ye�	��z���a�V����oc�Z6p풐$_TO��\��00�e�Itw���w����t�Ջ�[[��eqՅe�i8�R#�	��2�7T.�}�V�G��e7��*g��m��\���:d�:5���7n.�E�RWNf�R�PPW����ς�IxaԇoՒ���:�xt4bUkڽKc�6�|%�*	�E��c�%��5J.5�O͐D��� W���U�C^�G7	5K�Z������E�}x' �^�+J��:�u�p�����֠+Β�E3�RΪP��Cܥ��4��<8E<���;-�{M�/���X�0�m�Q��}R�1��7·�5�Zdw�]̩.	�8��<��]dD�u����7�p��s�r0�+x����D��l>��⽨�wgp�k޿�ͪ�V��}�Py�ß�ۃ�j�
�wo�1�VT#�6m����#F��Q�⺘��
��Ɇf�a�JC�Y���͊�kO���\W��>i�ܑ=��e�+b� E5$L#!Nɸ�A�0Pu�J;��Lگ�7DBs�a9s�"츌zk�]0�|�m'm��-�����J��3z�������؎�ym'���������_ZA��H�/GmnKX����u�)cJ֎��N]����.Y�w�{KpUb��$^�0T׭nL9}q��^�!��ǩ��&�ysF�ypjh�3d��"����Z�:&�f��Ȑpk��	��uN�����Iv��^�L������e�g�}*T�f2d5���t�0��*_%L���s��q��<���&�d�7cGE��e��I1p��U�D㎨���Ʉ0��(;J�K�Sڡ&*9�|��r�m��J�׸�E�l��n�j��2��זTk�k�@	��a�IY'���z0k6�x��Ԍ�+�Lf��7[�x�k�����^*����{� �/,���Zw��*Ǖp�&������P0З��w�u���U���]cۦ(�ѫj����jl(��X��ꪤs��p1G�~�_p������֍��Fa��Xh����*�I��m��;��F�+�zva�wHf+㮾�N�(����C(�琉
����Uкo:�f�:u]��XEF�f�&x��ʼ8;K5�Em��1!tD���	�h���r��yG���gĮ��U�6�A�R�B�{��F&(1��ERjw�&� ��ȗ��\t�.#K�	�v#)l�.���)p5G~$lg�-�.�����y�R�&��<�ݘ��T'7P!�~*�{yl�*YX��iR��[��ފ��w��si�6�e�V0z�q�oQ|&����Y��o*�.�xf��"Lt���u�YӅ�N�!�/aA��>�����\��^cX���..f=��-�gBO��]��@tK��󫥛�Yrvr���k�ޢ4T$��E�vM"������^�I����<���b~��O�-�k��}5�<~�ȶ@��<��uP�n��j�F�R��׺�!�\�x�.1��f(m���������:6�cDpL�+��ȥ�J�'>�4��}�hތn�է�z��!U>��P`�����q�2��O$paK�P^R��"9��)e9(�A����<�k�3nҜ�8տ��	�O��Y��P�ٌ�a��ճ��P}9F �n�9iܞ ����Fue��y��2<9�^CIϻ�w	�p�e�L_F��v��dp��>�zu��y�˱"ƈ8'�\�U�-�K�
+��<�u�mOc��( 7߲1�h���'ù%�O��7UPй�>���aa���^��i壿q��v[1�{o,�>�U��e��s�Q7Ł��^u�o'0�qd�
;8vX�N�cg�Ok��)�5�B�S�K��6F��(��ED[���O=����uV�Mp,��bvݧ��uf�w�w�{��a��צ��s�E,[��G��#١�9����6���6����B�x�y�t�[�v��X��M�K���0Ȇ{-�g��Ԃ��\�7@C&9�tŝLsD��^��N�������cR����Ưd]���ʼ-Zxt^%^� d��{,vC����zc"�I��f�*��YYkJ��P;#F�;��nLX�&8:�7L���eM�{��������=?n ��?w��om�}���s]�J���	��-�b��^�S���]P�"��^��wr͏s ��&_L��Nٕ��~.�w8.�ƅt Ҵ�f �qׅ?��0��p�0Mo����Ń%Gf���"鳃D1�^�#��l^.fu@�P/� 7����6�-]��0�0�}����@p�q�ƨ�1'I_4&r�-�!�å�B���7��FˬBz���K�_��9�1w��x��Y��Ó��Iy�eVxm�V�!��{'	h�^��o鉆��GC�pJ�p:Pw��Pؕ4"��8H���ܼӃtӃ����}Z>��",��ӄ���bbium�f�:��I���������z�d�M��N@Vz*�OYdg�<Ƞ�xv?���Ds��{L��{_�C|Z|�S�؂W�О�Q���!�%{��n]��Xޫ>�9OI���+D�w��ac�"��ӉjKEy��\����!f!pL����.̫�s��࠰l9`#[^�-��L|1+WR�P�͉����3���US�9�(�^����S,�gt�.�.�֖7 {[����ˣ�=K���çw��8I�9rV��U}r��M�
�B9<��̨� �88̾(>o3>��
1X���On����pSʻc:�#�KǙ�����ko���9V�3U�
Q�,Ʉ}�o!�����Ά�w4&�>���y�Jū�%��k=5���EɄ2�*���P��p�T;�e�%9#�byX�cʳ���9��ƛ���O�3l��t��2uSX�����u ɱ�?,r�*��5�^�\�Voj�\n���s��S� �_���Ù,b�]������g��káu�V�vfi��z�G�Ҫ9�V��i�\K��5(h�zk�f� C�ܪ@^��y��w͆5.�N�;��ٱ�&08�h��N�<���9l�v��U���=y O�v�o#g�OLML�Y�
eH���KBə~��|�̈́)�(<=�J�X�5´o�؝�exe�b�jr*}�Y'T��0�Vy����V�Ei����[�쫱u�}�����w��%�bϘ�i`;ղ�|�wo���'��i�f�)3������S�b��K��mνWssc�uu"���S�+-�gl�eR�a�s#�m��\}+���B,�'�:uo�T���;H�y��`��s�֕��:p�"ܧ�3���������2fT1(lY�}�l;�l�\cYb�*�/1��\c�8��ғ�7�[�L����^c|u��ޭ��+	�ft9�����Q�x�m�N��˂�n�Jb[Ϫ	u�r����^�����w\<Y����(,�k�y�:�8զW�ُ��mZ�v�/mI-�L�e��t�
�]nK;��H�ꔞ 5_�S�tDUj�=��' ��i��q�c>SH�,�������tb݈�(�8�mwL�=D;F�Kë⛫w�~�ZԾ{��,��Wd-��K��9�r�;�3s����W��{�^�.�q�r��h��#���:��eL�IV3k���b���u�m*�FKn�SyK0Y;t����;�u����R�;{6/�Z�)'[��.F̠ͤ�u��/r��H$�f�^Ä�U�x�t�K2�n'W�ŵBK��@u'D����ѥ�wz�Z�f���MD��8!M�R����q��T�p�A°WG�rgkK���� ��a�Vv�.:�ޥJk��D�;��K{��R���2��(S7t4���u���]��v���,V�}��-�9K[`�7v�m�}�$kH��b��y�|���B�WBv+� ��C�W��{���m��:��ǣt:��j.����:l�͝up��۬�l�Em�y���+�E��uV��Ʌ�[;�4�N�+U����j�.t����щ�+TU�K�'i}w5�a��$���fyI�byq�c�-��܊�mj%b[��E�g>��w.�1%��igDqQ��j�u,Ư�Ug��<<L�';�ѽ�7C�{e�&^�7G%�1�T��M͑)�>�=ܸY/7�:ܽH	:*����*�(��]�;j�TqDJm7{-(��w/�VsZ��`�Q��qD���{γ0P�pr{Q丯;QKJ��²��^\�W_Q��$Ϙ����ǯ!���n/7���l:���=�R}���+q
�ub�ʾ�ro������V��
O5�moR�'j�-;L-?p���W"�Y9�6K�>;k�ˠ􍛿B�h2�B�],:pM�7�-	p}��Uz&*�Y�9�U��?k�_n������5�f���1��2`
aԺ��D�0�������ﮗ�AveZƙ0h��E	����r�����~��5��(j{./�<�TB�j���U	���6I�^ewLF�/bu�Y�F� �+�Qz�#I�}yT����U{�.�^4��n #�n˂UL�g��;`���"�b*��x5��h�W����2tC��8hɀ�]+ �M]w2oe�d�S$M飍�i�Ehb��]�Ug)c��	�.خ]���f�u7RUmڭ�Q�Ab1E����(����k0JbU�TU�#iQTX�L�0�E�*�UTUPr�b����,e��,q�X�
���UQW�,`�-�TT@G-�TV"���+�ER�(1q���T\L�1E���m TR)

��PQb��a����d�ŨQ�XR��Z��U�`,2ܥX*+��H�73"��A�8ʮZ�+"0�9B�(,��j�ZUX�
�,��*Ă�%jR�P��84V6əAE1�TJ��h��#�`�2��d���(*Ȉ*��E�E*fY11rŊb��&2�"���+ER(�c*�mTL�Q�e��QmS1��d�-Y(�f5$TaFEYR��TKd��UDƱQU"��T���ڛ7O㮰TX.r!'c2h�Di��Q�n�Luj�'���*U���=$5�w-!A���#��FR���&�Ոm��Y�>��M�z�Y�������N8�
��ȉ:�A�1��P�q=�3l<LH/�)�u�|�!�)1P�
�C��<H?�6���+6��bT�D��>��1��"=��cp�Q7�7�_�6^�!�<C'K̕'�V|�y��L�%g�;��O��O��Ĩu��?'��U���q1�������/��0�>LI�P�q3����s3Ă�:�����������;Ӓ#}c;_o��"8G�,�{�ً ��c'�5���?!S��o�?!YY*���hi
��f�
�VM���c1�]�TfE�q�<2�aU���W�k���c�'�?{���a��
�J����"GЄ��p���}f�~q��gm$a����I�+��y�>�u10���$�x�YY�������2zv�VT�����Ax��3t�W�O8�P��/�|}�}��3�~��G�3*O^�b�dۊ�t}�����u#�&!ĕ���O2��Y�s;I���A}9�j$�c=��$���������i�&07ی�4�'�O�������~�n�y���_k���UXT�wT��8�3J�RT'�u�ĕ��d�����\�o�CI8�z��s�h}�`bI}�1��Ag�y�i*�������U���u���ϯm[��>/�������W�C�>��>�#�z�La�=LCVm3�;��$I��{t����^>�P�;�Ɉx~���O�T�Hy=�"��V����i�I�*zw�<a�Y8E�I��P�kco|yd�n�w�jk/`�T����hY�%I�/{�1�Vϧ�:�������P�a�~OM~�Ă�$�����wCĂ���&�|�I��1���~t���g�D1}�W��=�r4�n�yr�v4D��C���<Vm%�&?s�=H.'̙��~I�%O&��I�g̕����O�VO��$����������J���a��z�Y�{�v��P�!�׌��%ޗLਯh�'��c��0*vwz:���Ld�_�V|͡�����sԂ�m�M����At��V|��l��4�$���&zk	�4��.Z��bM�YԤ'|￷������:����<����D�5�*���.�U��gI��3zEj�7��j1�ѻ�gFX͌��	���-�جx�����yaZʕGz���+@�ݣ�(��v.�)1�Ƌ����5�]�㩭[�X���T�)��uK���������ԇfN�%�}�+6>���#��Q��
�~oG=J���g���H)>�0�xì+�>�x��bm&�{�g�~f!�w�CԂ������CKWl*6�&"B|~������;�}����I���Ӛ�8�P�,6�~CA�$��N0�_g�'�mO��4�m<���M���C�q�l��_��W���k��}b�O;?{�^5X��y�{��~�٦qH/C�E1'P�j�/Y6�ͦ�L��V{�~v���1=>�bIya�ϳ�=H/�>9�h��:�4�t��k=d�����ECQcы�̼�W39u������U!_X�"�Y��8��EU����d��4�Y���4���ĞC����UH/4�N!�m�&!��&3l��O���2)��][�����>�<=��:�%���s�*�������gV��T�I]��sxz��~Iy�4CI:�g��ړ�sbO�eaǎ�<�c6�R��b���H(jӉ��a\a�a���B#�����𣃔,{�*oݓ��=��$T<f'}��
N��N3�8�C?v�0�,�ę��LI�?w�u�ORx�eONw!�bI����y�'ɧ�ՊL@�<+ԅ�|E}�:X�фs�����������k��Y>f0:�?!Y>f>�w��x�u�=��u:��i�~jNv�07�4��*M�S��c��&!ǿ{��IY99���3��8�&!~5�1�������1�O��}�����Y���ER�<M��(bL@��H�m�����Xu&�>q��̑I�+�|é��f�|k���O{M$��Z>d�):�C�L@X>C�s��� ��6�l���7|~�͞����Hc?0���
ͳ�1>gM_P� ���٭�b�u�q��Y���{�C��I]��a�8�C�73�_)
��W|�Y5�����$�]�I����w����3���t��~�V|�R��:}�iI�T���LOm�q����Ci�?'�����Cl��0?'�1 ���Y�?&��}a�T��NoP:�'�/9��2i'P��p�f�n�����j7U*#�>���=~r�����y��˳asnt��B��֤�J6r�j[�l�ub�Zc�dO�yg/$V��]���p�`35����3��j,#2�� P]�g7�U�w�v?{��n�_t�
��*N���0�+��>�}�z��u+�d�E�����C2ɶb��T�B�d�?e����q=�P���Ă�>���wt1�l���*LC.j��߼�Ǔ0L�/z]u̅ޏ�F��sh�1�X}�i�g�Rc��kxT�����w��OP� �N_r�Cԕ'��b,�k=a��8�M�z��� )8�}g�u4���q.���|��<��鋬ƞfR�ѣ﹘��G�d}��16�Ow� Ұ�^3Ԃ�'�;��6�C���;�eg�1<?g��bAT<7ߵH|� {�gl1T>I|hJ��W��N���p�g�{���9��1DE��x�U��R~g��L�%�����}N�j�?=t���a4�2T�m��֏U'P���{�I�8��l+�P1��c��ڛOR4���%C��}�{�ϙ�Ox-����%׸G�|DFb"Gޚ�gԕ�x�j�@�T�����x�ɉ:�}�P�+�
��N!�+
�����x��~v�x�����_{a�5�'��f�9��O�����5ғ..�����Y&���{��`� ���C���Ri8��S���J�'9C{�VOR���1 ����a�J�Ͼ��3Oc�>�|CĂ��~�)<C������'ݳ��G�}�5��uO�uyT�V���>E����sĜB��=��x�'�WÝ�Rbx�`T7��ɛ��7�1�d������ �5C��x�^!�X(m8�3�<��tz�X���|�}�����M}�Z���"!�AT����
�C�1'��`i�a�͡�}���C�J��{�l�������+I�Әed��@�2��++�]'��3��*U�c� G�_��O��;�^���1?&0�ç;�X!���l�6�$u�1����>ъ���~O�g�{�q�Af�;�|��%I�~��c�LI�R��Uv�_���1C�#�#��� '�R��:�o�Щ��T�=Lv�QeI�n�m���}��I1�L�M��
���9�_Rq8��~�5*N>$�hb|_�VO���}�!�Ax��{��U~>�*��]�T�Yo.4�xw8�O6���Y3�;4p���b���%������X�9w����r�JsT� WK{gjW6��f�̹�í'��k@���N���%��;��S[��Z^�:��[`��dع�J��Lwye3:��8��Ճ�]�Tm%^��>��#�#�G���
�����'�b�Lx�d���&?e���Y:�z�s	�N�S�=�������s�]�q1���iԚvɜ��w?d4�2_�8��{{�ZlR՞5�wچ����G� |Bڏ��<H/��1��1���V)��ͳ���<N!�bAu�`~aS�|�3ܲc�6��'�x@�T:�ӝ�'1&Я��N$��X
�s����g����)V�^�}�:o�OP�������k��d��/��u�Vm���$�m1���՚k��?&x�:ʚH,��06���!�=�a����~O���$�������g���3�رvz,H�������qS笘����1�aU���$�*w�y߼��1%C�u1�J�*��'P���O�V��_��>I��*|C��|�"G�o��tXY.�4_������{����VO�Y�;��������é�1=a����%eg^$Ǻ�!�$g/�K���$���4ɛ���t�Ԩ�~jx[�%I�*l@觪k�=��.�r��?/�A � ��� m.��������3T�m�����s��|�U��o	1�1 �o�|��16�3��!�x�Y�o���1���
¦��sH��Y0(�J��z�����,Dh�$;�a4��T6��A~O�1'�I#�d����F�0&9_�<1����mg�}%��:��%��ݙ^r�i"�Y�Pm�i��`X^Dy�:�>V��p��L�:@:�&{��Vֹo�z#�X�Ob�˃<�w|,��[��q% 1j�G���6Ff�ζ�Or���}��e�I�����j�/<�fq�J:������Vk<y�
ϺS�(��{��A͑AG+�`�@[^�+�)q���׋e@��6~/a͡@\�K���j�WGE �[��/ ����jZ(�R0Sγ]R
b�&��\��ȥ�Ջ���=@�Nɠ��'������ۘF]��
,Q���Y0Ӆ�K���M���v����<L����w��jx��߉C�ٔ�&n�΀�`����wqw�;��;r.#�Շ�
e��U��[�"�까��<�]a�;o�{�WQ��[9`E9��N�I����Wв�C�i���KGC�(�8��Q);��^�m���}R����>�����6_���C���'�]Ӣ:![�-������������%��-�{�tOWi���Κ��>H�:����r����=� �yp5��[]�g#屒=O�J�ﻶ�"�O���	G'Nn �f�b5�@[.�A)�޾�)� �Ê�/���*���a�w��0��su��D'| ���R)�zMD�"�0Ptx|d�u�Q5}��(lQ>n�ӎOU�x���L����s6���$���5n`q$��{�U�0�FI4��UU"G)!TX~ǒ�oåJjL^�Nnb៟��X��qƉ}#h�+����=��u�9��H�t����X<�xj.�]��Ԗ;�d����c:U���5�W�Vt|�ok�����M,����A��G�Y�����鰲�M m�W- ջ�iv�����`��%���R��[7�ޤL���;(%V��w�!x4
X�R���X͖{7A�Ίq���t4��	c��(������2����x{o.;�3.,-k���a�x��_�堧n�n���dH8}~ooĽ���H��QR;�7⽸���bڃQ��7�r{�{~�7��q:n��.W�{F���@
<t�9��g��Y��-�?9�f���9]Y�ǰV��N����z�=#���ZJ��Do�,e|��&�b:�vۿ�T'}t���p��9sP�]�{W��e�G�{��*�|z�-�W��1Y�_e�'l�t��;���4�+��׵<f��ܹ���"���)vAV)3�+��~��Y8��Em�Ҫ(�M���壙,>&)�+'���Z�';s�WK쒭Ŝ~�Q�4�7 T���7�AT,���M4XΙcl��dn�J6�����!�H��q��o�w.�d���HU5LF���q89��6�8WVWfvn�OG�y�������:�ct	�o.Òx��B�% �T��BG�=�2�OZ@�ڔ��*��r����~����9�rDr7�N
�嫡O7HK	5_ʌ�z��rC�%��On�(���{n%J`�vewyX��K�|����,��r�jB��4������v�>��a�p�f���q.>2���ݚ����͍7HG�}{��
�k.�2^����j�R����1L���4kj�&1�Z��r���������<\�b�!�s6[6Ҩ�����j�8 ɼ+����QG%������K����g��2���kcD]i3�9�0_��a���s�\�V�������ڦF�	<�����x�G�k^���䘅h��et{[d�����hv�&#��dR�h��:�vaq];R�j�\�]�aQ�9��d&'���zz���]��~؋s�k�(C���DgeI���c����wC�2#�J@z��� ��%�3c���څ�/M^��F"M�tV�
�1���Tn�����%�*'G���x���f8]DL��nL!x9j�IwyW�ډ��:�7X]3v�D�e����"��NF��z~�ZVs���߆촃^s[;w�3��
��V{"�}��:��Z��w�F��$�0�dOLԦ��ML�5�F�4a�p��;�a���!����S�к��*ۧ�,еw�1˴ZD���Wa�>1	l���̠M�	ƓSǨs0;K'�|���MDj׵^&���[w�U��QNT��=�B�s3eU�
{�cN]v�tN\(�3[3f�ג�kt���&�\�{7~�(P+����|��5�b���⯢������k���]R#{@�v�2�ę��KGn�5
56e��x޴���%,�����{���f:G�*��ԍW?XP���"zjJ	I���u�+���x��pVg];�c.���J*˅ξ����x癎u,`1��qFEk��Ί�7�Ꙁ[�/�/f�r�b���h�e��\UØ�x�O�"鳑D1�n�]/X��E@��Niq�Nc%�̋Rr�9N��T��
��B�1жH��O	�T�#㥳c`�}P滠�e��UaY�zX^�L�;�ecx��y�]|O3�s���L,j�<�7��x�z'�����oƭ`^�vZ�=�XΣ[�q۪T����&�3��l�Ʋ�(;��G�oP�;)7׊�b�R&�C�AV� ��y�E|.\�d�;s"�������`���I<��f�y��TP�'�G �[��!�i��i����U`���2���E}��G���4s�)�>��7%q�=E�1�R
�ԞNj@h�7G��Keʜ'�F�wX���U��}a=��i�����5�t����ژ(�Dc�:Sʨ}^��s�k���+.�9�A�8�/�X����]Y�\��S"L��h�{��W���Z�X��7�ՠ�����p�̷�ʺ������}�`���x��ȅE�,@oQzwi����&�r��\�i���֬+��"�[�4f[��;O�X}G��4s�hK:W����#zi�PK80Gk�/�h�mWv<�3�;P�_й��B�[ݏ.\�N�ЎѸU?#����\�P��ְV�;'&ȋ/J�� Cܔ�LZrB*&���ˇ����K��P��^����^���M�0�%��G��D� ś7�퉬i��T�W&�m�7,2^�Gw����<�lw	�k��ˉ�0���x:�w�*DD�4�cJ�9$ld-����vx>8%��rt����1ے�f�jP�kڞ=�J늩�kH\\j�\�ٗ~��*��^���5�ӫAΐtH�9�#��j��%7��"���!Z��nP�����.S[�F�)�m]zz���MwBr��������ʠ�f>z���#j:%ѣ��˓��M}g�[��nth�i���cj�^��m�H�îT�n�Cy���|���Y]F(�	���d\����=	����kLp!��L��� E��#D3HȤ����C1�!#\d���Χ^��׸�Ѥn�z���N����Э�7�#��8:�gd
�'7��vJz������v��d�W��Eb�s�;�e1JR�I��נ�F1Fբ�
�eJV�a��d��LI�*������2���Qٻ�Ϋ��Y�*�%N�mdSތ�����F��(�d֛����*#�o"r&a3NUh=���\�@�;'�P��
$�jN�d�\Z�F`��r��`;�t���f����b����b�u{�d�~T`h�~�n�P�=�u�����ܹ�YL��Figpt�7�4L]B]nrc��RPw��I�Ĭa��L==�S��{��nE�r��M׺�`�׆��Uڠ����nM���øv�{�م�R��̯Rg�C釶��z��ˏ��i9P|v���{U��ê]ڭ1�}�vu2ҿ��Ŝ�n��F�T���� �`�9៱��[���������t�{77�-g��ΜWR�U�Ku�	�t��|��ΨY��ԃ��#�G:&�;���R�۩��qz�λ���qΕ��و�u3�s�M�0g�����}��LM�{h�H�.�3��xw�y!��޳�ͮrR?���.k�L똸�t�;���Θ/%2���4�+��e��ImW=*JY�Ϫ�X�QX;uM�����s8��շ\uTPQ���&飪>��l2�gk��*����j�2&�↟̻_c�.
6��AɄCG��wA���/�{�v�a�3�Ȥ-n�&�$Uto���B0n�N;�G
I��{�ޓ�o���w�H��+z��.���߭�B�Ɍ��)Z6�f��e��ڤ�Oƭ�;x��R�X���P��DW[ʶ:��CC�ϋD"�'vf<7eK��4��)����7}q�!R1������uΡ�p�C��X�(��]�h�X��!�32R̚��r������.Ee&���T��nu�����t��H�k���Ӓ�V�O�0�,���wIX�\gs����i���JSK�*]��%� r�*�AX�E�3��KG�5y�i�ɔ4��L���ڀ��X5\�!}�cZ㢄�C�H��(�C	�E�8g���� ��&��k����c��>6v�n��3�F��#�B�Q���ּ$0*�,��8�7������=�j��<�ΰ�tw��7�%<Lwmᥩ�9��<�DS�dZ� 7���%�;z��׆�$6ve[��eP�Q�:q���!��tb�Z���g��s4�V�������U�T\*Q5Ѿ�(ر]�/�gY�*�`f�6�Cc�FH��A;�n��65v�?<E�LKb�� [�7}e���ٯ��'X��ǃr�e噳@�s��j;|����H��$@���gj0[��J�r�MhYv
k]�̵����3�:������n�j��q���ѽ$2�*ሄ:�f�X��Y�(�9в.ے+]�v�/.cї���7V��e�o]l�قn�X���+Ō�j�{g�:=�.%�4U��M��M
-|�q��^�v\�y`9S:�nOi�W"��98䋈�@"k�z������5��Wu��Cx.
Ȕ�n-��-��L�p�!�wx>3E�NM�Z�:��hdƵ%y`��v�T��4���{@�rҾ���2u��e��R�W+�|�����G@�Nc{�����l�9� /���î���q��!nch�I�;�
�9ލ�C��ˢ��VR|p��x�_�G��Y��ۨ��;���<��9ண5i��o]�]IP�e_l�2'0B�g�+�6%�8�l��I���<k��Y��F���-�w;K��Ѻc��t} ���q�.�B��Z$0�;�x��PRU�)�
kE���^b�4�.�@�,Ƕ-�;�eXﰩ}���Q�b�nV�f���HB��y].I�̾��aͧ�rbc�/ϴ����}3L����][�\}H�ǹ�&uI����$eZ�+71�L��k{@əNd��L������Ѿ�˭jk�&�����m��Ᏻ���Dޞ|�����1pO҂9�ڊ�!�c�FA�i�j<�a������w�^�Q����mv<JZ��3�̜����6�Tt�b�B	 ��uv;߿�=�ٿu����Tb
m�Ƞ(*�+
�"�b!�ɂ1@�X�Q�"�dU��EH����RbV+mA̸���±b�X�-UQEX���U
�%ekQUVT+-DQE��E����+�iEjU�*0R",E$\��b��+A��CT���T��V\lP�,� �9b����RV(��&R�3DXe�(����R
-�(��)P*
F�Kl�DAE+X�H9H�RV�KV(%���UcZ"�U$Y[b�EX�QUjT�T�� ���b�XbV(���21"�X�@[EP(�	mH(���am*UH�*�)U!PV�����*JȪ

A`�"�E �,XT���V��,`6Ud�,���� ��m�1��<������i�~Qu>8�B�v��,53��Y��.ѳ����[�V\΂��Z�]�l�Q�Ϗe�](d&��w%�ٗ��W��K>����5�2�e�Cf|(�S�����@LT�M�H����M4Xݜ��K�lL�+;�'Ԁٜ4��ϙc*eވ �ʳj!d�o�/�4�|N�j�μ�)
"yZ�[𞽱�U�X��'P���J���	�COQEX!)�����?^���c,L��(�(�u�Wo�Q���?"�w������yrC�J�� ob�j�w���%;F�C)�$)�ā�q��v��L�6�x�y*�\.y3�mK�Y�W���4o;���d
�3đX0ѩ=}d'&�e�a���5s�7��S��VK��찯���IQw���1�YW��b%麫��x���2�V��k�ҧ9�����ف����2{},�]_o�����ap�.��# u�5}<ٮ�e�ۅn�b�?m�j8 �&��]���K�����E����Ɇ)�ݩ{�$`� ����(�7���n�-�8�Z:���m[���;�l?;��h���q��rܶ��t��#n�|�����dn��Ö�^<�������U���R8*�L��܆�U�Ȣ+l�n��#Ἲy���;�����ݾ�c|��d	��__&"t|�Y�cZ��� ��q���jM�1P�Ny+�ᑲ��� ����'�=o�ˎ����G��6�y����q�҄B2�UU}�T��>��Eu�����GW-'����i��^0x9�2�v1���~=�< u�q����k��q*vɄ"�q��1/�j�x<7��� �u�N��8�3�4琮l�D��*�w��=����^�ah�W��Aj�<0^%^N��u#K�7:A�ⷢQf��\R�o�i^l�k�"[?9�2�K�0}�V+_�T�t9�,������odۿ;�>�g�V�ثn
1��վ9��Q�q��u�����/�ej��`�ZR�mGJ����l�M���Wְ�Qg�KG��/�9H�:�0w�KX�[4#mH�tr!,yp��v��M���S� zTh���}jb��P�뇈�l���zP���v�ڔW\f�%�Fд�i��#�rw�;�Q�*.Phŭ�8.:'a$��Rf4E����q�������>qw�#i��%��h�������9���T�x��F5c{�{�U��q�d��,~�Q��Sr߅,�T�Z��]8���Wz�&��gG��+�e��A�}�3��8���g</ؙ�m:�I]ld���Ze�[Z��/ʲ=.\�8,�7Gh����*�ծZ\Ӿ�xpn4��#Y�`A�҈��ހ�f�Ŗ�I*c[�in6����e)V(j�u��mh�M�)x��:p�!�Q
,R������ct,���d����V"�N
ϡց��EY��L㶐K�K�s�@V�Va�������c��!6e������.����� :��dU�D@�^�{7�i�԰u�S8-��\5�4�mPDz�"�_�k���s�w"+6$:ji������:m��6�]��m��M�5b81CT^W�Qs��d��f���9�7�Z1h�ctt�{w�r�R�$A�ګj:՜MFud���ԗƝPz�f�`b�d^:�P[�����gf��Lж��+dI���W��Zj�X8W�X��P��� C߷) 2(��*�M�S���V�ed���B�N_c���ņ�Z�;��J���aY�Q���ĕn�n�Q�y�U836 �r���tɶc��Z#��pѕ���]��.�(0�g��l��q0�{������ͬy���뛔z�o;~c��1�.6�+T���Fv�p*M�(������T��u
�FKf=.h8u�	�g��6^�`~���{]B�qVYKzW[N�,�3��m
�.f-.��y��ȫ�EO\�Ѥw������9˵�=*�z�"BC���
x7gl��MC�)�\��{�K�����8�ǵ(.6퀝^�[{�V����^ãul,�C���__p����֛���2+��8�c��{����;dtW,� C%�S���O!-���:�8�p�.{�V��m	<{����Kt���{�������4T�ԣ,����Y5��z-����~z�n�|[Eu��A�'�ۀ�� [���1�{\��>P���%���=�0�5��Q�*�t\�*�ZO#���I��@��𑂾u� 6�B���}]4�OvFԥ��0Χ�1�S٥�=�u���M+�kΧ��[�{*z�OٍU
r$����k9т�o�tSY�m��"Yc����ρLaa��3_V��ϜͳRo����Y&��ÜF�pmNx}�~�*��s9�V�S�Dy��?Oا��#$�/��nb����#�������Y0\�.7����I��7S�`�|5�LM=0y�#�|I�pͫI/q�GRd#sv�b�(Oc���2��H�s�Z��j]b�iu[堨�zR�F��\أ�aQ z�����T�����E	����k��ɏ
��
>}��e����.���2{�̳�~>5W��Z)����V���K�x�)Q�Y� ��ȧ���-kY��Kw�ĝY�	�^q(���hg�+�Z)K�)A�w8#W�v�V���B��qN�L�5G�|�j�Uk��9�*Z-������H��ϰ[R������ogo+˖/a�3�vt�0R,�	�pF��p0�iy�"�������r)��ۭP"h�K�4[��)çq�Z��f#�R�m�vɱ�8��|��£����xcFTɚiSr�u��F'}2�p���:9է��X��Q؄5������ׇ�l�%��Qy\��G0��	n��������,؋�k�S`��>�� v�O%�p����c���=�)]�;;��e=��Nu���[�V�yFx����F�/�{�'M�[���a�#��u<E-�2j���e+�vź�:=�t�Za2��J���A8T���)
����S�e*�W^�tv���JZ�����	����s'�P�}D`���T�����#
c%�p���-R�ݎ*F�O�\���47O��.��'$G#i�J�ZuQ!rάs]����h\'��G�vm�R��;T���.1p!�w�֙\��ˇ3#��'L��yG�'Θ����f�@z����#\1�U��o�pׅ����j�!��!�.���N�D�Ж�����)*�(���#!	�^
/&]�ʜ�l&�'��n�_��%���|_F�*��U�+]���D��X$�@��Ϫ��R���̜���U1� ̬�i~s���)DY�nF[��m��v�ی>@,/�-uD.��i�wP~����S��VӉ�+tϣjb5��ˣ��2�V��>&���H?�/ܪ��5L�r���ܽ}X���2#�J�M�!��(��ALsf��|v��\en��_���c���e�U�����S�X06����B��@>F� �z�[�+�%�y����֘���J1�p/#U�o�� �]Cg�n[�3���9��0�T;G*p�~���y��W��AiHM����k���	x�����Sq�1�����"�ߓ�ƣM���T� ��(Q�h稟:^�F��<��o��,~bb�ς��#���mׄZS��#��(Bܭ��y����:���|}�����f����jK��Zx`�ī���@�u��c���RJ�xM�mt�54 �k��|�pm�e���Z����
ChՊ��U<X�`��gf���ӣF�q�4�'yk��Ќzݾ:�1j)���o�p�tu�ȞN�������n��5��^e�z�,��]'��5���{*��j����,<7�R1���Uu!��"6��<7�F���p��֮�];�K�]� �ƫ:%%�Ԑ�(m��LF0I�un�n.��$鏮�2)2`	a�H���h��kK��ԉo9��Bw�*�d`��(],ORt�˞�_���n<�,ߦi;��R[��r����i��94����
q��rQ�����y��Y�O�.}�Ҩ�9��b��I>�xT�l�ن7NC(D�v� R��#�Ps�5��C�y�`@ޕR6
� U����GQ\tM$�#�T��⫷���g}1�wF��t�Ul��~��1���v=��c�3�l���[,*�}Ox1�h�U����`חj:j'J�u��OOy4"ʥI��#�11��GC��6��h��yzJ.�u�o���D�V"��N�q�rm�� .7�2�V�ſ+o���bW:��!]��;�d���ሸLN
Oj�Ϝ�6�J�@
�̲����VW�1������Q+,�4�����$s�U�t=.�BS+䤈�N��@|[�������3n��R�b9��A����k<S���r��ٙ�C0���G�Trl�F�{��'Ns���Oi�U2��έ���Y���S�"�)��޿exX�*�R�^TI��F{��ד�X`޽3�j5u���5�R�P;>����� W�{�Km�4Ofq>��h���u��}��ˮih�r�`>9i'���^˭�-�m&�fn����pH�	q+A%��q�C#�O��9_
f���#�x��x�Z-O���:�)]QWU���n�E񦕞��՜��M�!��<	��d]���=ɽ=w������諭���_z����+2H�5�h@�86���Eb�X/�N�!Yk���c!7qV�(ksw�q���� 3j5۳����l�#���W;|4f�����\0�,�����t
�g�$���i	p���#4��r�r9U�N���a��T�oE�>���;���ת�&�]�<O���^�׮2eb��]Q,�9��0��y��Hƌ��3�Ӛ����C���9�1�bqt�Q�PMoy��
uSA���-:�gs1��J���Л[[g
�Q[
����)��t�d�X��1N�q69���Ȏ5/q�ڼ],M��Vmb�ӷ��Xp��n���N�����c��;)��y���+T�|v�NCB������Q���W���*S���J(��F%	˚�@�ck����uw�x�%���oOYd�ws�k�+��}0�_5�A�P^m!*���#^�8�>��\���Ǟe�X����pP�Ĺ�9�gt����Qɚ��>�b�͢�⭠9j�b��=��.�^�m��2��V��]�ga8-	�i2��jҧ��=�=~Öš�ĨsV�e��v�.��J(���`��98Y��2�-�5]��G��}�Im�ח�ȩ���e�ْ�l�ﾏ�>����oV'�a�z`5c����l��u����:�1&� ���XU������)=ƛ�d��s�9�is�p
�$�Y=�I�Q5P��*0+,l��!����H�v�	�*p�q��������&+�W��ʐG/^���#�+W}�eA�㞋�(Qk��JޮWW���R |Pa]�Ru@v�R2�׏�[�t�3�m-u0ګIxݳ|R2�H0��t�}�ʰ`�[�p �qx���U8��:]P��A�D�7R#�v��qcg��r��9��V�;�J��f#�\���b;���5;��q�9Q��|mN��}Ϫ*b��o";�Xt��xe�[�:�#��쿹;`�:l�1���T~�>,zyJ.��X�C���кo:�|����*�^<����ָK���$~��Ps*��oB!M�����݈,4Or�ϧ�׏��Q�
�{�'M�5�|M��H��X6-�=�ߴ��L�T�u��z�c#�X�q�{L\Br��D��
�R"�DK	��5���I!;�p�PF��Z�R	;[ӭ_T!̯�%ܮ�n�u�s��M ����z���E]�)��֦h��R���q�tS��K6����a��[|�B�`����8d�0�k.�/����=�a�*n�Rc�o�h�<�y�?�*�8�G�DDl���9|�AqY�i��{P�9�D�;�Ց���C�Et'-{��=ʊS�um����8ח��g�����W��q��R��rDr7��e�bk����|�p����@�^�Q�:�T�1{�]
�����獌m�I�L�ch�w�$�ۧ]���Ow�26��{�d�;��w�[O�C�����.��!�놷0�V���j��'cMگP6w��5]=n�Y^gI�#!��[�]Z�4��t���/ԝ[��Z���yT2E'����B!䨁#�lL�6gA��n&�\en��[f�1a���w�x�*�KE�}H`�J�0���ڠ#uA�`�^Uܴ,u�>��n٠m�p��3�.�q���q�r�;�-�c>n�Y�*����42f�v�%}+j(V;�2����V7�%�hׅ����k�gT�.[�N��3��+��q���27]�ޖ���h��W��g�V�k֞&�?��ku���k��Ȇ�v��N����[�/��h����ju�Mc�F�N�m���ťx�p�W���;-+#���V��t�!n̩gx���n�f�Mz�.��ռR��/Ec$�b&œ��f��r��du�s�N�)a��	Y�։YL���U;6c�̺�YB����x��������ν�Z�`zV%o����6!��=d@Iu�*�����!�c�}a�C)�O�8^r=����^S*�v���L�V�p[)�OM5l�ˬ����a��R�0��[9��chazX���%�se�^�ܝ�f�6෷cچ����:�[�/�������3KOza�+]�Q5A|���b���p������Ii�w]D�djjTv|_X{�$�X�E��c���&��WN�ۑ{��|����!a���{(��ak;�0/�ڼ�G�����Nj]۷�Ҹw?���՛V���^�wC���6�`��X��~}.���
.��x�ؕVfܜn�M����O������������ו%�>��|�<vL��LWvëuT�ty�+w2�*RLR@7Q�����6�7.���p)�� �Y����:�_l��p�w��6������n�X���X�coo9���<��ｙ���*��#O+D
��w������c5z�&~3��L��u���ڲ�L80 R@i�����&9��
����t�_4z������_1�Z�W/��7�lJ������@(ݎ�
��H5Ʉ�4]
���>Y�� �]c�����÷��d^�܂esZ&�'�sU�˲��NY�x^���H��[Lk�^AE(��ӛҭr�>����[�}�^
��<�E�4� \|�t^n�����v���/.��2x3yz�dՎB�������E[	�ժ۾8-��Z3V"�f�����{��A#�>���}xq�k�:�6lK�`0Ѡil�(��m��0�'te<s{��l2�G�ۘ�� ����@ 9X��!L���7�Vs�m�|�E�X��bm��֮2𻥉t9��� .+L�W�o[���99��`Н�ct���Y�v'� Q��H	�~]��Ȍ��[��}-2�|L�{���c�p9����Rk��k��'G������}q_u��k�LTW
��j�*�҂ ����$=���_�#n�:�������2Ɋkɜd�#MW��2m�:������T�]N}8V��}���օ����8tN��Lv�����D��b���mG��=Օ�c�#��Y��*�����]�F��7{	l�����V�E鰸�[X�5R���:�NG{Y���UA�.�	�l�hei�|��y����ގ��r���⥣�����D7-�L��.�a��כ��8�8k��o��UTX)��m���YTPX���(�#++�X,X*�2+Z#+X�UEE��"���J!�fR���,�Qb�-����6�E���*��
"#aZ��$$�2��T`��,ER,QArؠ�Ra�PR"�؀�UPV�T, �X��U�����Kh��UQIP���mE؍j	n!�X���P�*Ab�ª��DA��#*Ҫ���R�0�[�Lea�1���* �+X
�b
AA�%�TTE��X)��Q*J��ĬX#(�
(Ԕ`�r��@���E���X,TD���P���G�����q�P�F,X)Z��%d���`������������F�z_7s�J_p{��"�`�z�Q�&�����{���	\��^�|�q�o*�+3��1��2���W��}�<}�}���D����o���ȑb�����Q%|a
����bU��d d�R�u3��xW�c�Ut�	�SE�l���xm��ò;�j��
ChՊ֕OC��k�EM���O�B�`T�x��|����DQ���1�%��e����\;>ؙ�Q%��Z�\�ݫ�i6G��*��$..�m�&T�_`�V�#%��ᇶ�F�i�Yfꕠཇײ� *����(	�UEY�R1 �ԟ\<E�g>!��oe�bd:�˄f�Pa��yi����[�G��@�& 䁽t�(@��A��G�D�%o0�E�����0ޔs�7�6U� h���C�txd<�?)=$gl����.�0��泴4��w��sQ)K3~�S�s=b�=�*_����b�&;`A\v�&9��&&"���9q� [�YIb�Fpư� �ʓ�|�hCF�rw�;�w.�W��2<cv�,��C"iaR�7��i�<���S��q�8n�@�!&f��}V�.@��� :�<6EZtDE�����goI���l͛��쑎��Ǵ�Y`L�ͨ>���U�N�,[uy�\�N��B׆��jt�l�Y���gM]��`�aV]�F��� =�\��J��D����zE;v�����̶hO��ڲ.�"�_1ȯ�=�a�}
��YEIy���F(��Q����""��o��� N����!�E��5�itR1�ab��	;�7��é�?	��+p����!�j�y�C��:��*
��s�K9���.�����\50Q�M����ō�,|�
��Լ��}���yWlgnG��a�~��3j�+!�*�@�o]��LoU�~�����t��^��<����x.�uH�t��=��~��X�sw
�u�M\��V�NbӒ-=� s����"����ؒ��3�	c�D�[x�b隣j�wb+T�3H�S��D,tɰ�=���|"�;�4f�_>'�Ķ*��HU�-���o��q�B�:���}7."B����9�a�ܖ#4�5(h�������*{f���W����ު�Q0p;m�ﮥ�L�Zل��Rw�s��l�;mڔ����ۺmR,Sҿ,��#OiL� ;KP�|����\ ��!����|�+�>M��~���%��e��7���S=u]f���J2Π7��2�&�j�2���R�5v�؂2�� �&�y�,�;)��Y�~雔5*w�/��{���ME�5�P�����B���fF�6�%�V���+,8���![���ˀ!35� 8�Fw5e�d�x��λ%�;�}�P����,TkV�,WCg6���:�b��U_UW��c��A�T��]��֛ϳ�{��&��������>H�9+����4��/*��E��S�!���{��V�������E})�q�oi�H�L�2):sp��C1�g�=e�YsS�"�Dt��|uWa�%#����D&�����-M��:�;S#z\_;G�C�nB\���� V-j>�(4S������̂Bgt���&k�����3h�%9QX��m2�Y��^V��@S��$��@q^㖭�N����ّg��Hj2LV��VA�rp�V�]���m�����}����XK��x��)ᮩ7S����׆��A���a}�}Oޫ���[+��LJT-򫒅�jb���z��ߡƁ��vFq��k��r�MҹM��%nh�/���v)LC�qu�Pc~j�V��s l�QBEs�_V�:l��"�v���:�M_T]�~^L`���vwi 8gb�N70�=1H�x��H�ؽ��t�l�wg�z�y�9���a��N� ���A�V�`�S}W��2T�u��E}�ط{YSR�a�ٖ�ti�����R&�DNV yYhj+j�HlW��o�nw���ݼ�*����m�h�g�6�;ܢ�cT:���}'W-�����ܜ2 ��"�L�e�����a���)�*���*Gʍn�ؑ����">�G�5V��ޫȟ�P>�Fa��#����.�u��WZ�#�����1�1�������EIN�l}{ְ�Sʏ$���ڰUк|]R��Ԡׄid��{o��t�9�����4�;�&8'�s��m�h��n�7H�˩����Q�W��m��of_�S#����N��4�_�X^���eK�F��9o�)cE�y����b�5*�1U�$체Y<���Z�+�=���t}�b�ۇ��B�z%܇�F�N���eJ+ Sfg��H�0�7����%�81S��eqy��6�G�NR,	��Vt���}�[�g�����`�p��LE�H�*_��a����6�&��L��QEE�����һ2,E�N�q��A��㈌�F�kT����ħx`���b�pC�fj���c_��͚��gGZ��s��fᘎ�]�R�a�_�o�uk����t����x�7ɨ�zҨo�!��C��e��X��:�j�y�\	/�lM�.����0�!v{GU��[v��E'H5%WW{��n�s�{��g��=j���QV�)�O�\���,Q+��D9����B�S�ً��#'_���ژ��c��F�d�N��(m3t֡����u:owGuw�iϱ얪#1 �fKO��0V��Zh���u/��ꪯ���Q>�QGO܎�����=,XJ��㌈b��`5�Ayv$_Ä�	���re^�oѪ�+���3�f�S�.�(���� ��+�c�fY�t}��ww0l�U�E����[�q�gq��!�2��uHׅ���z��W��?rWU�]S��
��O&g�"[o��'V��8��V�����g��'<�e���=U���w��P�_m�h��]���Şoh��]P�!ѕ�J`8oҳ����-7�)݌��IB\�75�&'Gm�a*��J������Ce�r�ū����}r�e��"(FtL�f�u�	��m�����ǌ��
[S���;\r#[��N�땗��=5ô��-��7�	���^�.C�y?����p�K*��p����]��tQ��,h��wZ�u�|l�v��=
�؞+����1L��J�����VD��R}P�.�9��n��Uz����Z��tr�ܧ}��^���ᇵ������AR�
��1p�H��
�[���[D��x7�{1��ιQVuքM405c�Z�����|��߷,峔l���],���v\�YF����v�?vu��ʻ��bp�[�ѝ��!�T)�zt���ixu�_lK��r�j�ڦ�-�Ys1]X(�O&Y�ŕ2�ǑmX��hSɈ�y�U�UU}�S�yX�ē��{䂤�C<#E}eP�]�L�EOQ�y���+%Nx�����(`�\�P��l�ϏW�Lv>�\�i�=�~�g�ͦ��<Ckc�]"a>S���ۗ�g�B]��Z!��|Y;�2Ö��$x��s6='z�ǹP�s ����W8���޵Z��0�Um�0����"�rsz2Urn�!�)� u'�ȗz�Uj=VM#���_�D�ȡ�5�1�_h�x����]i�|�ȫC���N͛�5@4^�Ug!�"�̲�fV-2��Ͻ_a�I_T��{p�+CA���*�(i���A�6�w���N���.C\�̴���0�QS�)�|�T�4��ƙ���a��)�E�W��X	�_og%�S��ѐ�u�����c����֚��{�k�5����(l�m��cim,���)F�"�#�c�)�"��bJ����/��Bѩ`�܇=;�J|l:ᝨ^�Մg���qtF_N�ؒ��U���"o଼H�8�?v�yf��j��y���o���i�+/�vP�mpi��)��5`��ª*�]�����iT����5��<9h�z���G9V�C�5'��-�e5gf�]�f�,C)M�t�(V蘲�07��Na��m����b\���s�������~.p�Z�#�}�}���&���r6s�2�2�`��U�}V��pm#����x^�ZRd�Q���^��WhPj�y H��C�۪@O׮�a(�s/�Շ�fj�ڱ����ܔ���Ӽk�h�[1oU@G�2@�'H�@mN󓇂�,���1ۥ��t�Z�fR׮�L��ູ�Oi_2����큂;\#�F�}$���;
r��z��1��j�w�6u�����CM+|;����彎8ʱ	H�KJ����l��r�8��-����7zb�q��u�OPy���r�e�1jI��,
������nQ�n�d������wve�qN�M"��ގ��&m0O@��Ko�S��>�}���!��V�_�<���-���{O38Y�u���Y��]��+3�t�'d&4aY��j-�5�f1c��z�CwQ%��-�nO^Z�Xy	�q�p��J\)�u���_mD]Qy��ޔ�ℱU��_����
���@���+ks�FB��Y�bű����� �3p��4��%[��'��5�j�Ǟ^f�]/> �F�7�+��b�4�+Y���R �e��t��_j��U�|����ﾵ�\.
�:��v�ۖ�Zڂ��yN��'�p:�
ܣ����_nH��9֓�_,���b�D�Svԕ�����g���cow9�v�"q-Ϝ�7�]�ޠ��t�x�FV�ȕՎ��#Y�݉f�o�^�`�^-Ԕ�O1l�؄��44��}��Q�}�)�]M{��%�tb��Y77��������}�C��qw�Y=U��_��w���q��q�w�a	�@�kr)��6�,�S1^�<lo���l����3՝�n�xz`�*{h�r>�3f���J�\��M�}�p�}�; ��R����J7јVƧ+�P�wv�W&_5��(��B�����5��T����a�oJ�8���QT�\K�}|�-�����ZW��_<)�bT�f��W�����:�����a��2�V��⎘�]ƾR����>�����Q��HN�*>�G���s���z��Ll�Q�� ��I�Na�o �%���vr��b�L�o3��\������X�|m�d�.��L��ѭ�g�n#��F�ahl����G7r�WDJ�[�/��5��]�7��쐄��xr��u8�p��S��R��	mJ~���'��&�����y���˨��Aw9�(>Jq��Ӏ�B��%.�ʹ��.ڃ�\�6/���`����a.M����=���C7���r:�<1?+g�A]����гZ�rM��+��2��ݐ�%drN�5Tp�q͞��<)�󋼩k�To*p���:�Y���.{IQu�B��>���;�p��k�5��(�uˠR�;�/b�����w�+�*z1�_<�~v�����z�"1��A�z����O�V~�ϸ��}������[_2=�G���Y�IH �����~���'��"}�g����4���Gݜ3�SF�4���n�۹L�J��O(�x͢�^���~�<�հmP�%vf�x��pW�Y���L�a�ؼz�j�¶��D+ͨN�o^�����s�S�~�߰�u�p����e�_fi��`i����v��U�z�E.��`,i���Eg�*�i=�]Yno.V�g%�s�/�: �=S�x��ۺ8*�����>��Y�6�.oqO�{n.Lo�m�z�{���u ��g��^���}��}��]Ix�������;Qe3�A��Gޯ"}����~����xN�q����D���2z/��ug������w[�iv�v������;�K�nSA�_u2�mt����������'�i}�F98�^���f�bFf�[�k�x�hK��B��s	p�M`���\�K�t�b��dy��,��xC�ܭ�ɇt���U�!)�BR�g�Ϭ�VIW��K�XJ�'\M1[z�J�6��uuBk����T����T��]�9�1=�6[9&鲐��T�rk. %��}��/�����B��V\��PnjH�{����|�"�?t��#�g��/~I���5o (yP���t��7��U�N���Q��y�8TA}�^Վ�xg9��Z�����MB���u�듊�STYŜ<�8�|)/=�/��/{ﳣ�1�x�ɀ����֚MEa�Y%��=;k�n�Iv>�O`��q�a�9n=�J̊S�3�Vs�g�E$&"�}�Co����a}�iH.���x��þ4�>�δo���q���1b�A#ivI�]AW�pe�*�[�-�M�9%7o#�����tw��pV����n4�WW�N�-���(���Jf�N])N��gj���]2�*�i�BM�uJ��6Ћ�@��hO�P�ϘΣ����<7���r��}��x�R����#�<��Mڶ��6韑�_�Ui�R �];�m��RДq�7f�Y^.�n�=��;�6rҟ�u�ֶ-�+���p.��tE�V+���3\M��5l��Y(�9q��9�q�N���j�B�o/��{8ԩt�hKm�U�P��kW��Y]���g؋Z��k�x�e��E���y>�ݧ��T����������=�`�!�a�8����S��*al�8st㳅�J��R)Rů�!y�AH����2��0�%-oo��ʮ�I{�ϟ�"7�w6�l�:��j�2μCz�a;�d���7i����j��mS��k�{��r���9�ON���"���8�m�"V��
�L�Z�����^��<��K��a�x�	O�vח�{�^4�(^�
{��ee4V^����'i�JRV��'��&��Y|�9�דѾ�z���Vn�$�a]�s]�N�]�7f������>��7�{R����2���"40���=B�A1��6�&c�;.Ԍo")[���^�l�E5 �\�m�z�SJ�6cq=cܶ���Z�\O�^ܫ���`�*�U��fcEf�r��:@˙�	���p.�����%��J�w��55n�Xػ0D�+�óqJ�e���� �po���
/u��(�2��NuīaYa\��/��ކ*�}M���#�_QYN;W�u%����u��%f�]��ޣ�- `��.�&;�g:N��)2��L���Ǣ�;�r.[ɺ�15�p��l�Z1�E�F����,���RK������t`м�~h�+ܯ��Mu�n�4s�`]�͔y�W��*��C�NU垫�4m��O�;��zn$ʤ��5��m.,���H<<3@n����F�B*�x��g���]R˕:��\ǚńrk`�7l�v_ݸM�i3-�ST�2��,���ɯ*f�y��`�������I������^ë����h���o�f�B�:{��)S9�Rv>=��}v�!�/�8�����Mo���ד*w�\�JBG1�u��㑗M��p>=�nl75w��Z
���ú��[ԥ�LVV�ݰ�mvc�#u��k5t�WyXF��,ٺ��|Dx��<.�����$���� +��Wv�ߟ(�.�����[�Y_;n
�⋫�Y{^�|�aD���#����CT�^�3�|L��!����\�AV>�Rb���ʁ���iEҬ�3-L�u�(ED\���Lb��ekY�`�
���T�Q�(��dPR) *�KJ���E
$��+��֒�k��[Q�Ƃ�+
��A�
Dih�IX�Ab��ZDJ�P��VJ�R��ֲ)+e@�,s(�J��̍*Ҍ����B��b�X"(��T�R�b�V.R��&0�EE
�C2��[-(���TE�
�%H[`���V!X9HT���6�`���Z	JUV��PY"��eH,R
�-�EUQq%AQQUb�Ұ�Q�(
DATZ1�+"Ŗ�*�� c1�5��E�P��+q�@X,D���� T�J�,�E&0q��J�*LB�U�<�f+�G"+z�),˰$���j���v���J��K;1Z4G,��<}0���q���t���vBH�7��Vw�����@z��{�z�wW�E�������7��q��c���V�ΪJ���2/S�qNWT�/�t�������˩�8�|7���e]سpԅ�b�dOJ�n�s���u�a��ت~K�o��	=�M�����&���Ͻ�OUo������0V)�5%�
�|�{!ں�>(�K+}RP9OlvQ�_KS}J��n9Y�YɼXך5��v�o`�ђ�|��v!�ZP�od������k>���-��:]3��x%u���\�\�ܞTs�D��N9&�)��{>աu�d����A��*/�Pc"��=�l��y��]���.�Q��7�[t8,�
ddoW�Gh��b��)�X���]��ksw�![�jZI���{w�{���B�eݕ�[g������jr:�D������壩w��o8+z2~�t��
�]۹�{�A����u��a�8i7��zn�Р�����-l8Wv���+l�� ��V3z顫�y���I�n�C"�s��{�1�z�vɄ�#~'37��{���d�}�\�\�A�-q�_�%\V{���;���գ�i,I.*7�ڻNK7�M���W������$p1����������w�O��0��|f\GN�|�T=N��Ј���6+���ckj=�wK�5�ç�3yф�Jܼ��g{ɝ&C�;�N���.�S�+4���u|�D�Rc�A]�imE����,{�Q֕a�FX��x9Ҿ�_ڝ�_ɳU��]��66�|�����=����U�mx����g�b󯒢�%kj�<�p�:�u�[��]�q5�����J�hw�V�Z�׋uh;X�z[ߚ���!8�_<8:bS�w���NR���i}� ��O�2��F�-X�R�f���_�w����T��ac��{<'}�����X����z�/P��eԛ�
o|Sj�ܛ~�Lt]�n���}��CL|��*9K�LfVh��F7Wek�6�[ow>��P�-��^����U��QZ��z��^��۸sz�%�^�q�w�Q�&`���B�6M��t�&r'��Y��Y��t��Y5�˲�^�*�J\��`'��9�{�龫K�]���k#��
=�G�՚�ĒыFÏ%�x=�}^N� Oz�Ft�츸�@���]�#4�&<o8cr��������w�c���OS[��m���[-�GJž�U��y����u���&�wv֟yVcd��yE-{�\��/��o.#v��*�;
�g;�Y��� ڙ��zܞsn�u�ĵ¾��֎���-'�Q!�����<�-�#A����J ����_j~	o��
��.1GLR���o�On���ȵ�k�`�R��]u�.1�t�2�p��BY�t���컎��Q�Bҥu��9�V�W����9�'��Qϕʘ�٦9�p1+^H�9��eݪ�[c&�4�J�=z�i�}�}N��o���9_'�U˞WmZ�v/��n����6����jz��������u�;�T=����b�Lsg�������a�;�jF���r��UkN,s����T]B6���!M�jNJ�<z ]�w�',���%V�dG�9ΠL�j5h3i�r�vԕ�q=A�W1�K}+̆�����۽�utO�w:5���WZ��\�hB�����*�'�����[X�x���ޛt������騭�GҩVs�s{���9Q���)��n���z�ش[MHrƱZ��bsE�Өq�����=&�W\�J��Uf��_U}�2�(?��.��(q0����E��8��������{Mn(Qi���7�ɜYvkt����&�7~fi�Y<0���A}���uE��ލ�S�訠�"��4��t����V*x�����0��b���'n�$	=uxm0ʧnwV���fq�oHu�tc��:ێ�l\F8zG����G�ۏ�뺣��ׄ���d�71O	Ϩa�}�S8�/���y�\�T}�m��m�X���Ӽ��ր�I��:ǿdo2P�^�1�)�7�������kP�<�T+K�dlW;�^�B�[]U+��>�=|�c�����X"�8Ft6��_���W�յ�v�u��BS��ި�0���YWgy��P�#Ӗ�'�,��[�mKJ�jT��<�g�r�+��r
٨�Ut���twCY;��[֔[Hӝ\�pJ!��_<�*�O_�m�ج��;l�z�urt,�Ռ����]^��Ux���w��7O|��yS�l`�T[.�w�J;΢TYF�~��ͫ�=1p�a0�b�aS�]MN�vž}�u�|�f�>�+������J�Tv�ngn� K�#E3�8_V�܃p�Sc����� ]�F��>�>�]
�˅����C�:�/�2��6��i[�q�mB��6Q�$":�8�x1á��Pc����nN'��9e$�T'���T=o�j&ě��t�{��W�B}�����٬4��E��<�R��&���d��ہ���W�%���K>.D���{,�ڌ���3��mo|<�)���:��E��ٙ ���6�Ug�=Ã�Kc�3G��
��|�8͌��Ȼ���S��󁜽qԞ�8�hgv����>�cr��<�&}zS����J�x1����h����ek"z���?$�*����ј;7����G�窎�K]j�du~�ɔb�;%�Z#�qCGsչ�j�s=a7rN۷��1ݎ�FXֻ����tm�+:�/��v�9;�j�ĵuӥ i����k�v��V}\��r|���`t�ڞ�2	gF^#$�����VD?]�kB�vR�Y[uzhzA�����Vu��b^���P���M�4�XK�]^M�iy��`b�K�0���~w�c�(�VQ�7��\(��d{��6��x�z�˹'6�R)V���Եca�yt�޾���W��B�p�(ic�»�,��5���s!Eq���/w�+S����|�IXϯir���z��9���|Zˌq۶�ڂ���m��L���G�@������ 9N��b�}����_4�|;s�9��[��̢>��nU��r�3q5Q���*�3.����	qU{�i>�o4'�������H�Y��8�ژ}���TJ~���-wave�N���5�wHmo݋v�2���}�'����W��{0���K���ʞ�w�"���b�]�jdB�����I]���F�uƥF�L��n:�ȟ�1¾+��-��a:�
�ol��
�V8�Q	Ѻ�&*�MC�S���%�;.������9�闷��/�L�<~�n�%r�]�;IK���'}������^�-[q�&��Rm?��uD^gU��zڌ�m�RV��6���²�F��#Yr%���)aV���\n�Y�t���?Z��I�u�[� ����T��#���Z�]=�-�-��b��t�Mʳ4�m�kk!ǘBl�4��鐭8+���丯A:�o��X؆����%V5�,m@�rm!d� !�?}�}�}U�M�T�Sĕ��r
�u�WQoUE��OM�t��{�p�ؕ����ɷe��T��ȉ�^v6��{ �a����<����q�ƕ�m޷;:���K�H5���#}��x|1*b���-c�g|0���CR�q�}V�깉��O�׸��V��v�Yv���m}v;��Q*6��z�^�o�2O�F��X��Fƞ~)T�cYp�kr����쿓���q�� (8̹X.3+�|��.T�z&+WTvW;�/���-�F�]��u��:�%�aur7�t[�����`tj��R�__5����I�A����n��b*��h'زjھ�ͧ���p!)	n\+�c�?$�7���]�z����{��O�h��r���s�9m|a*�a>�!�x��'F�e-���[�!Y��������,īF'�]�9�s"�Z.����iiw����j�"�(��ʰ��vB���A�L��}�$Y�궮�<�2]�����k1RX�r�S�.ekwvM=�.b�2������f�LN��tj��J@d�&BY�껕����HOW��d�ġ��	 (���WZ�FY�C���}�>
-kp����;s!���5��)��l(uy�,�y��91Zo2	����*�.9�;�5���YIQ�N_C*�p��&�@� n��6��p��7��;�Pkv��<6��\��+�l�-�7W%��׹��2G~��<9qվ5����ʋǵ�A���[�Y��Փ�I�L%�Fa�pɍWN���,^�wW�uy9��E)�M��10�����urLZ���Z�l8����I���7+��+���G�ٮ��c�:YR*�#�]T���nx�^uQ�SM��y�U������٨,<��Qjw��9�Z���V�������벱��#d���hr�%Ҋ?`�mu�+��|0Υ������Oq}M�� ��X��Yٻ���r�SH>�q*�Ug��[I�|����O-=��x�qlN���.�ኴ��'�!]���8��p����g��޿��e$���K8����2��r���G�e���ٳ��>[5r�8�J�tN�$��)q�P���fQd��m��/y������hR.Z2^\J��X�9��}��M�n=���>����[Q��U�d��Pz`�k��%&*�G1�񡛺�aSm�OD�����o�u�5Xs�����ڂ�;��R��%��B\2���3�-����C�Y8� �)���i[�ܞ��wI\�U�!)�	wGpR�K��3.�Sdk��w;��^�O>䭜Э�S��+��5.��+����m�����3�+A�z�����6�����C��SUuY4/<���+�=�mIp������0�i�[�V��i2�6���X
����[:����ȭ�u> �c�Ak(�ڋ���<3��o-�gDU\8�^<G��6���U�>D��l�l���vѥז�/@ʕ�u���pP�Q�{�u�WnѵQ�8=p�i�U^0��죉�dN�"�ט,��>�K�Nsb2�O��ݵ:�d46c�N��e_�hme��-����3O��SeO������5՝�Y�9>޽�M}�܀⒃��"�X�4ĵ�w\nu�%v�}��Md�Ž{�8�c��c7kcǦ	6����X���*󖹚�V�Q�tkn�4~�@x$ԕm�r`�ź4�C=�G�r�f̦o;�˯�S���eu#)�'��Qߙ�_����7�B�
S7	k��c�b�iv˵k#�kg%d��Wd����V��r�i�e��0���<�(���VxZ��?_R��.��*���6���N�cEک��Q&So���������w���R�ֵQg��}�]\���l(�'ݭ�*���v��Ko�S}E_e^�]Q�zNF��-���Np�:j�}��
A������w	�/��CݾL��o��(R0�Fn��T���qǝ\U�wh��b��
��M%�v���U�J�u1�N�v㘬D��b7dl$x��9���K��qu�k��1,�I��F��ڝO8kΧ5�*W�`��J����]�|SM#B����x��mb�Un��ج�G?�a�r����Pa:�lD��'�S�����5j�.��s}�
vw+<�B����Dײ�7�~͂	��s�.� ��&$+�0����cR�i˽����o��V��S@W�='7a���8#��CQ�)�[�J����Չ����eZ	�W�p�˨#'��6���]Y�����Γ��Z<(ؚ�+S��WNv0S�跎��ʲ�3\��u��v�ۃ:��i��.����Z�a�����$Job�#�h&^雱��1�k%h� �I����p9H+X�҈k�"�C�/��#��&�P�ث8���K��ս/ 2�����;-�Y�n��(L�n�W���5�l�3�wQ<Z3�=��6���j@�Y���]��������n��D�}v�ژ̼B�f�3&��c��H�3�b�42�kȃ�V��C U�j���\�[����2�pJ���S�����Ip��T�]֫=����;l̌o�+���P�y޵3�)7�܁�>��O�ϯ(b �f�'����ӝ}I�]x�̮��F53s�.���S���d�E�y��V�@7I-�`��]�Z1�S+j6��n����j���F���t���*1*pf�b5���/�������G�	�}9'oĂTc��4r�mI�,S�n��ܺ��~X)8��Zy����˭`����\�[Zr�gd2������̌*#7���2����[��#�6�w*3�j�9�b�5'کQ�y@���4n�ώ��� �W�]!��h�,j�v���d?v�2��+�:t��S�����΁b�A�)�2[�e3���D���*vY���j���`�vpu�c�a��B���T渹�9�PS[�5�3�C7��hԦ73)O�fwM#8T]B�J}�R)�LC	�(��bu�]�St��E�^Y���u���6�/���gn$�O1l*�6 2���($�� M��7κ.YMoλ��u%偰���A��d�ǌ�9!v�:g��*<U���7�'/�f�Ź}��ҕ�R�Gؚ���+j\YA%��B���+��}�������r�k�]@��!	����_e.�ڔں���n�m�8mۙ���������	�Bb'���9 FvJI��N:"��z#u'�������'n!f�t���U��(@Fӫ�n�=��h�{�3NVt<xq#��p0a���8�"\��mnT�e�vl�Ṽ]^��А+5��E@��*�n�(����M��5���WBҎ���];�2��|�l��2�����yץg#ns�}W�mݻ���U��%�y���Et@�IPf�&]j�A)s���-�5Ǉ^V�˄�W��2���'���(<����`3��b�7���xI׹���Ж`E�Z�J3�E�-�`X/\+�'l��t'��*P%X�q���tu '˫���(bw�9����Y����*��bm̖�m�ٸ�vf��l��ʽ�*`�lX��5�ב76��9������������]�&آ���'̨`�E�H

,�@*L�Bba
�(A`�d�Z����`�� RT���%q��AL��%�,�ԅ`)*)+"�c	m�BT��VH��l�b�b�Y�V
(�72�ŕ��J��*\l1�DQT�YRJ��YB��Ȳ@�*���X�V0R�aIXB�(E"�@YYQ�"0 �
E��,�IJ0RJ�T*H�� �� �X�TE �+!U�d�� ,���Z�j���˪˫�Ǚ��mSs��j�=���5�[]p� ����n��:����!���$\OI /$���~I�A �Vb���U}+^��������;Q�[����OGT7�?Rc�]xim[����gV��aPiku�e��;l5�	Q��&*�MC�9��c�b�4��̓.�(-�g�N>x�i�X�'_%E�Ol[j_���<A��fv(�4�qr���+-�q+�uo#��n�Iz.C*c(�-eU�3|�}�e�,9_ju�Q�v�u��bzi[L�^o�S�;�����O���{�����T/�$��VA�3�����TQ��D���1} ��yws�)}@&G�?�G�|œs���	5G�=��[��C�iŨN;9��}���h8���E,��<[k��c��*��ŷ�·m&�Zrkw����Y�w9\�#eR��kZ���)���޸������a>���l�Ó�љ�u��rm�Ծr�ޖ���n�ɽ�jK��tRX���f����d�KM�.vM��΁*��������?AX�(xu��S>iU\8���M��t.)�&�۵����Ba]�c7�t�]ə�a���R+�̀�c�����kM��n��'�`oV���������ܸ���}}]�ѐ��7��j�����s##]D�1)p���ksw�)=h�����U��Q��u-��7��{�����R��~	W��~	p���.1Gc�YH>����[�����8lw+z2]Ҕ˕��U�&�ڞ}�w$�F^����w���'��C�闚q�@��8�B[�c�&Ηײ��E�^o30C��Yp7�,s�Mg��!��n!�GT'�a\��[�>0�P<�B��I����:J{�9e$�r�I�j�/ wH�ęs��,[���=Gn�T��}�Ǿ���:ޝŎk��i*.��VI܋Z'X���(�ꧣ��a���:�#՜���.Q^m<2��Ǫ�W�fP3��53�+�Qp�l��\l�G��/��TA�u~�xoԓ�[6�6��]���.9lK�M3�F���;�I�ʈ�7+�����޿��y��j�F�������D'�Ĭ�/J���\�i=�ư��Wr�b�����Onm`���#��K8� &`�����6�(ַf����pu^Z7�.q]7y4^[<�c�UxL42V�9+�8����5e��g,�Ԕ��]�\��'���Z���gw8u���i+�����8�̏������S�/o�Z�&�М�fŽ�?v&*-c�q)����ὢ�uc�4�=�UM�o��9����aDa�a��!�E�X��K��x4}G�U�[̍f#��+�w��; ��[�h}:�a��SS֥�m���8�y�TkegbQ<�@Í���y�p7�/�Ԩ3�TY��k�Ϣ^H+�3����|�&�n�k�oj
�V;
��A郱��A�Rb�-����0#D�4�y��.jw�)���9�ڂ�<������\�wB���Z�|��B��A��ˇ��)v���W�7�����=�������̾�p9��:�+���9�u��\����F�ή�� �sUD<��Z�����J�.S��j71\�y�vg@N~o����;�m�S�4Ὕ&����b_f���_h��L��8�f�9e$�2�Ď����/X<��{7��Z,F����&���c�F�����K��2$qP��i��\`�y�rXGRu�I����'ۇ��?O��睝N����1M�HL�
�M��1�;u�%Y���rE�*���S�Ϟ���H�ii�E[
��	�Lp��(�ڈ�O}���꤄�⁡;+���oQƮSp��)�P�����+�����DKl4A�;v9����G�:����UM��K�qIU��'��7Z�]ٻN�L����,�xӵ��<ڼ��L��m���b��ti<9��o5����/�/�|}���l�����2�����i�OW� E�Ӵ70� 8r��t3h��ͧ4uY�Dm�ʃ�\Ue�*����T�njB8K
��V��R���� %F�">���-uk��t�,㯠ێYs�g	��N����jU�&��4�r)���bۍz{���u��eg/G�ԯ�-��5��T�}���.�>��5���W��,냳z5���������D��hqk�|������qk/v��&������V��$�Ǣ��ţ쥚,��R�%����Yvn�|&k�qy�/s��;m��nuCn�BO-\�Z���=���)����n���;_֝���h��%�E�T�Қ�{'Z-^�ݙWZN[�|r������<����s�|з��.o�}��d��脅�\�:������L.�o��Z:~���Z���w�<g{�\΢j��� 9�P:���{FBU�09��\�֎��B{�D�j�W)+K�gB��G]+b�F!�����˕kj%5�0���.#�q���/���>G��X��`.C�.��ҧ��|x����T�)�u-tF�U�Z���sڜ�R:����l�{-�6���NGSy��PWeDZD����ygoU�y�T.5��}
���b�5�� a�;,�-Yk����jv�#w�w��*�Zg�xrz��=�ڃ��<��e�P��ooN�{]���C����#e�	��>]���*W>���rKwff�������"=x��옇w�'�^�:�#=U��:x�,�e)R�6}��Z�p�[�8A�}!Jv��Χ�b���X`Z}�SBܕ����<1m'�P_}d�],>�\W١�<�Q��]���y�(V�wL�e7*��T��6�E�ѥ�úK���ӑg�]m%��o7�Ij�� Y����Y늡۪���QB�R+��T��a�=�)h�+[�j��F��{��M��C�}���SNM���[P�[��)��u]LY=�Z�~�~�>c��ĳv�r�l��z�(꧞}�O�o��=���y-���1叨m�<�c�����\�}/�1�Dj�{���K���-�s�DFʥc��>Ƶ�M�^s"�-�>/kW$��iĽ��ny��C�N�M�:�{|����SKc�1Ҽ�3j��5��z�ȅT��j��dK�E�X�wRz��6/.O��s3}Z�0�U��8�vIIcj��o~�3�E�+8b��u��1�_KM��Y�-B}Ԙ�OE�S	���	eDJb�nZ�Qy�&�N0��̌˦������:��9�����\����m�\?mf�K=�z4�R�/�k�#��$[����?g�gy�g����t���[���kX(c�:�n��6%vMDb{���E�yH:�?�y��s8M&��x��)KW]�V��c��]�Ru<c��N�x����k�i'˦�t�����`�e7��"�ba���A#p�\��R�9�d�2,w9h�C�ih7+o���S��1I��dK�|j. ./�aL9]���͚����u�:�^W������
ٴ�m��W&r"���nHI~G�Ck��������zױ�Udg���K��FoT紹\��%�lѤ�oQ�=N1(IK��l����-���:��Qx��h/B�f��aAk�Bi��gyx)�rWy^'R�Y���˂�Q�u����ǳR*����LV����\lG]'q�W4º�����o��O}���l���0qk�fg���mE��qocqF��ژ����;͍yƱa�4%�3&T�e�6�:��E�/�����:��1�-aN���K���w������fɪ�a����&w�\}Y��g��ha�X51���"����E�{��	%�ސJ@�ro�EO,lQ�{���X������v�����雕�Q�3���-|��I�W{�����]}*ғUY��Nv����Jz�S��v�m�4����`t��+����*��ݚ�j��b'�����-��jiu�J���aR����ˮS#�w�7��Q�`\_F�i��ތ�T3]�c9�Ym�wCKˬ�&:�.�����"�C�v�ά#��P���w��`}C����X��Ο'78�����]�$C}֊�����M.�P�J�E'��TP��wZ�e,��"�A�2���v���5L�K��.wp�����s��=�<�B��p���˭6�B����?P+)Z<�we�1\%k���2�w'4����D�:�珬i�䦼���x������n�0�i���ɬOv�,�v3(����
�,�;�0L��>��A2S�S�Ԟ4��P_e|im������iA��ia����WS|A��k�ۮ�;�L�je�D^�{.
�.R;�@P��O7�t����O�ǀ�v�I]��]��yN�7�uHsp�䡮ܝ�x}]�Cz=�=XL{�}�͢%m'mۥZ�lC�6��M��n�'ww�����l�����(��������/;���b�[�����;��XO1d�db�g.�2�S�́צ���*��{]��H�}K/��`:!�G�KUZ[ٜ��#Z��۫��ƪti�&-�Z'�-:��KhHl�~��׮<��xzӛ��%=�vd��3x�m��*�ΫJ�bܼwq]��v�'B�^�Ȥ ��+l�vm���H�H��3��|�ՒƵ�U|㳞��41:���>9����Y[��&��cO�>��Mbۍz{�2�r%@�7�+I	�*o��lץ�^*N��t�Ᏺ�mvS}Qұnvj댃ڣj�e����қ������|�|���i�q-eÎ�ގ�Ŷ7N��3XM�b2�D�Z�)����Lwh�\�\-���M+�û{v魎��0F�v�v��y��dRm���zf>�\�h���q;#�����r����'sBp�R���K��5�a)�������]�יn�啗��Sk���,������	�'�c��.�	����dA��[��褽^b���di���.�6��ʇ7
�A�S:W;y*���%�8���*�;ç��������u	1T����=�!����zy�"3��	�w����ڧ�o��ݤ����(g���LW�}U��h&��`�aրE]�j����O�|E�u��X��\�bS��_\,:O)Z�9�L��M7���U���/j3r�d�j]v9%+'r��Nq֕��97�X��7.t��䧋:�Z�q���M931�X������-�ŀ�gbv�P��6�O9��{7r��]�����&�in�����|�WEnQ�uy���k�f+oKuUY��z�ɶ�-�3a�o�J�k����ŉʇ��<��[���۸��.���W��F�P�*��~�A�Qp����VOd�0u-�!s���W2xG��Խ�\׽}^%�}���<>�1d����Ŋ���x���2ڻ~�\9��Q�9Tl�ˍM��ۇ����zC�|qq��z��q����}��,V0:�zo:����]��_��M�����ƅ.��67�`�Wk���/��H'<�{�<핚�o&���2����Cri�����16�Dfk��v�g+҅0�YQ�)p�j�hⷺ,
[�̉SzL�5�sL�GS��n�ѓ�7c��b���U.f %����/*��EF�S`�=׋/����*}����@kG>]su�ۖ�aܓr�����yDj���r�*�sc����͙���v*i�_��,�U#\mdR�L�Z�5x\|�Ƅܡf��֤Y��<�v�Nm7x�Z��Y��͖Z�@d[�^Pzٹ�eeLm�U$P�Y���He��>�����xQ��r�˳y�+�q��*]�,���B�'m������z����`�tF1o�9u� �ke�%������ �R<�d㙡k��9�x?7[V�ox�޾�|����u�Ύ
�a�7}�O�'�'�I���3e����޵g�X��O�\q7Q4B�z{X��4�y�c*d ��Jh�z^�dd�6̴�FWZ5��X͕D`�=Eg��瑉�����z����@w����E���}9̫���)m���ؓ
S�P�z�n�ow(V-�oI`v�����L�CQ"{瓮��耼uvP�`�bb�-~���AqHB��yx��΂VL�u�wP�(pc,�e��ֻ��.̲^Z���J�6��']:(��y�71Q2�뾤y�qN�����:��a�n�f��1E��ހ��N���9���q��<��M[�7ֽ�f�ŭX��$%-�v,��{G���u]�c9�.����(�"�mm5ԭ|���"h7(K�u�n̡|��ҕ�M����d%��@��x)X͕n|�ʰz�/��4����]\��y�Ò�Ҭ^
L��b��INp;�%ݕ��f�2m�ޞAV\J��8ҝ{��-R� ]]ao*�rBC�2Ę�;���v�{qŦ�g%6���)2d�;{uyC1%Hp�/�-��vV�H䧱(�x�6rUAv��u���o.tY�+��(7�icV�ta_}n�#���OX˝Y�y�)�#l�Q*��6fxҶ�ڷ(I�q������e�zE7yvMM�7[c��e�KW���ik�5��B��V?O�z��)(��棩����"���6��FqG����5�v��DRc��ȳ�s�M�%�9�����{�E�x�ɪ28��ج2n�!Y��5Jr[{��˷f�rR��t���2�^ZwL��{[oL�yaէ����S�������$���M�Źw��0�`oU_����7x��f,��fՉOo�;�L��_�5�D����%�Y�	:��On�py�;@��'qj7��r&���S��	�&�5�k�{Fڪ@k�h3紲���`=� -L������A��ЊL�b4�v0<�1VZ6tu�̱a:��j�zP����W�sN�ф�s������I���mI|r���s�E�I|��/�W�$�ԥ��&{<��gF{Vݷ`��'��-�-+�s7;= m�j��'�X3e��-R�}׽f�xLK��@^�達�R��ɵ�J��zY�[}��Gx=��70`�z�haAS4N�k�Ԅĳxw*�M������]^�Nw��ɺ7�待��ȭz�|�~���b<O �dΝ�[��mW�}�U@}_"���)*�k*�U��F�ʬ%eaQ`�`TR���D�)"�"�a,��il*�D�R)Uc�a+�Y
���D�V,���-�kH�Ĭ+�m
�H�QHVJ�"
*ŃK��P����PmQJ2�XQ��Z���+"�F1���aYF�Q�#kl�	�\(,�)X���*���*(��HT��J���[j�D�1��P����@D��f0�$�Tr�Hc
ʑB����B��ԩ*B�F$U��m �XV��m�J�2��r��R�QH����LI����F�E/�p&�;���u kX��E�Z�`HNq%׀�#&�sq��-Ͷ1��%��J���+HT�,mv���+o}�:b��n�LjJ!��wJj�+�L$��u��\b�b�����l2�k��]���[_[H�9�ؽ�&5T<�?+�1YB�c�yȫ��K|G�9�ﲏ���l^"��V��s�~�Ư������*���^Դ)w4�p�Zt�f�հevMb{�:c�Fm�]<����*�	{8�v�n����׳�������-��η�չP��gS����Sv���r�x�i14N<�__%g���<G8Y��nQ�u����h8Y[ۡ�u�!
����B7�:�%T�IPތ��5��Yq��8�+{�n��9�9�A�q�r���k�ek#�ڣ���"�/_��Dܓ��@�\���M%X}���H��>�篾�꞉x<�AX��K���;�Z�}%��-����4�g�
�W��[q[m�ۉ��W}�feH�CیAZ���U�*蓗nP���V[S����^w�ށ¶cy�-�S��O4�/z놶(,��A��!�t�57ua���9���2�*�G{)��2�i*n`�a��3�Y�u5[�v_��Wlrt��b�I�MA��	(q�ZN���l��Ӿ��vL|U�m��lK�̞���B�Gd�VNL}<��F���έ��j��OT�xѷvXz�z�j�W��4�T;{PUr�<҃�r5�J���= 󛌜:n�3���G#-�N�s�'�8��A��oj'_@�)X�D��3��v�q�&��yU�QE�K�Zk/壦�i��W��ܮ��t�u�r�w�ح`�θ���JWL�����jn�9�����4-f��]^p������"�i�L�d�WXt��-����+]�뾁ɶ�gFE���b���w�]Y�Tտ�ޅm�+v::
�f�2�'̌�Bӳ	�S���NU
���u5'��7Q	�B�x�Ɗ-e[x:c1���{E�i�Z��-wlֵ����1T���������3���פj�e��f��9k
ۣ}� �>b��;>Z�?>}�n�4fN;��ͮ~�Yf�R�G�l=��{���r��`喩s)R�)�D}����
�:�Mu���=��H�R���'I�\4x;m$���ٶ���Y+UH�d��b��j���N�+�n�J�mA�j]#f�r��j�GHz���&`�f�%�^b���L�Q;��G�hh�g�k����C�<^�L`�)h�g��0w��^�Qo�A���ȫ�KJvng�t2[��;��W���E��j���V�0�C˻�+�hgܮ`Hf�+���������i8R�#>^X�g� �կ�I'�CY��h�S+Չט����U���S�Z����d�+��.)^�8q��Ŭ��R"s��}����N1��&��oz
���v���ݬy����}��u~X�x���)��5?_Pr,����q�[�����7�,mTܬܩ�6����z��~�������H��{�˅����i��Y���Ѭ��YwΩ�|���D��q�&��[+�%#a*�{�o�
��V��ٹ�3ws"t}{��8iE/�s�2q{�^����p�av�Gz�:�HGWt��9�Kuo�r��X|RC�W6DY�p�X��aVY�%:����e��E(m�vթNI��6��`��A4ᥢ���+h� �綨+�N9v���m��K�z�:��yc�M3��P7{?;�4��W�0�q���X���}��l��LE�l�f��t��j
����	�*���W*x\�!8q?5���o�����9v\��ⲹ3��}Nٴ�S���K8a�ޞݽ3k�x>��	�gu���9�a�mE�N�&��7m��ݜ�Y@TݡT�};/�RO�����:�yfц��{	QuI���]3�ԕ����+6&k�<��^��V�}���u��(�7�>�N��3żN3��~��'��U�[u޳{��h��Tr[��NՊeVn���;P�/9�����0��C��)D�XiÇ���{���v�*SZ�]�r}�:�*�����ź�Q�M9�(�Oy�iq�1d���z<�×hO��{}6�i]C����=�W&Ŷ�:)f�By�zUۿ���[y`�j����FX�\�:V�dri��Ep��s�9:�|���7,J4�xp�tq57|��4'���LKV]|/���{����X�2���C+�t{;`̊��E��p�T�#�f۠ў��e0�_f�%%��9���ۄ�r�f�����h�RR����a�|���Ow˶ʿ�L�Ʋ�O�|�@�x�4��"\�oQ�K�����õ�k;�u�Óu�\�|�&��Tp�� �nb��Ȃigvc�7�U��V��	�z�1__5B7#A�����ѮU��9���ZK���x���f�R��`dpfm�f#�˙8���T4z_��2}M��ޤ���轇t��*�%��Yӕ��c�*���Q7&�#Ku8�����]�'V�5����
�%0�y3�1h�g*�Z��]��<�0���p1+^\��ϓX�B�n����)�֫`��r��lMm�r煗���&��>�c��Z�ہ��k�O���=���u�g�v�/�i���4����xf-c��r�Ʊ;���1'u�e�- �P�����u�[�k�E�,f��γ���d�Τ����H71��B���I�\��3^[�R��K�����j�w�i�Z�K��^�֭���������;�ֳ�u��9m�qCβJt]ޮ��'6��a���\��`��q�he�k3�>�Y�*�*�V�&�2V��,�g��	l-��� fo5R����ɾYk��y��z�J�Tx*4P�=��W-<꼜��2�L{§�Gf��i���:F�Ҥm��~ɆQ�X6G��}X{�}��>�FV�jzǋ7��q��[�E��,��&�VrEPU��z�뜘�x�(���֭lLf�k-E��^�w=gS�<Y~8�w�+�叨{s���h\ş*�����i췃gh.��!�{�=��nk͆�����y��A�q�ݱ�6Ϫ���lY<S�pm=�B޵�-Tl�_N�K�C��WT.¶��;�7kh��VP�Y��_�t�I�o�Wo�����|���S��53���v��w'Q���k}��G\T$��2�Qo��������I��ׂ����En�»�_U�m3Ȫ��Jc�c�V��oLRo;龎��_� �Ǫ�wV�yc�!uK�v���$�3T��^���[q�CKI��vd��<���B� S�Xf��2���)�5[e	Ӥ2��b��\��51B���9�ձ���;0F��׃��u0zu^�~~����m'|��E�ӲͲ��MF	Z��8�ᒮ�2��.ڃ���wve���4��ZG�o[�{��7��Y�_�!��-�x%\��+�1Θ��H��뷜;�ڰ��M�ֺh90z��H�w򜎤���LpW{�x[_zF�ߖN��1g����8z�(4���{Տ�{n^�1�;���h8�z�@g��;� ~�{� �9���֧�Nu�RU|�A��\��E�빂v�c����?Y}���u�;�OVg�;�)t������ڼ�M�
ft�T��Νo�L�Gi�]�o��>Ow�ګ�e�P�:� %w���/�"n�8v���œՐ{�'oh}���C���20H��l�ff�i�����*.�q6ܛ�����:������y�^~y\
�֗u+��\��gUe�n�-���T+���C�叾�ݫF��L[�1v\��U���Ue���5�YR'�>w�v�SY���)+1�v\ĎnE�v5�R�NHL�厙��T��:�i�U����U�`p�9����#���kNڵgp��9��fit�tvG)�[4�΅ڄ��JN������-�����U+�nC��ķ.U�B��f�S��7O��u���'
^J���1W�W�)���;�-�8�Ά-]��z�=�cg��zk�g����]<�7�g�3�Jx��J�}�Q��|��q�Kg��]V�n�%��W�ۮ	>L�����޴8\z�^�(�`�SD�	L��҂���]9�5q�{B�^d�"����o\O��E���}���_{-�?W����AWL��^�Ǽ~��LJˣ��zp�@<;MǹS��7Q������s�G�!����˕$\����u:0�׵�0�NǼ��O������F|\�N�#,j~�����ǣӔ�3�9w��	�~�Z���h�Es� �~���,�չ�b:�{ٕ\rNb�=�1��N���hS��M6�zs�7�דG=`o�ːE.f�����C�����kNMDj�</��׀��O�u~���×���.h��֞]��:h��蒎\��ax��T;�7�<��3O�������2�1ƱQ-�j\K�"����gN^�B��ɖ6��Kt�;K��T�ӺG-PX�R��o �f��j�$K|މl����|7���x�N�S��߮,�՞i�|���+��y�v�����b+���{��M�gs� (U��9��R���q#�o�o�/e�3�c���������r�e���b�������G|.���st���Nx`��l�
[�!3��:�µ�\JyS�QpT����?^ƚ�<5�ϖt�=q��
�=#=7��`u����֣�+ޮ��鉿>Օ��#�k��U!�/�z%~?}�.;���ɭ>N���\��ꡖ�y�1���Qn�we�ל	3^~Bf.��#����ݍC_����#0����__~~X���۸O#���{�xg�m�&��1�zq�N�Ŝ�헺s��L+�O1�ު��'�>�ꓨ�}����e�ۺ��N�9�.s1	�2=�ܶp���]oNC(-����q+�g�mK=�@�@�M��%~P,��j����c�o�j�~�\{>g��Ͻ�Y�>ミ���mK/�_���tp�=n�Z鹜��ei.2P^;��_^��n��c����x�3�w�.���Z���}0o���B�Uq�}11�����:�G�o�S�:bTz���~����r��O����v;��zMt�QR�0j���Y�F���ų�2vA�y��ԭ�曝;6 uCX-.���v��O���׻�<^W�j��$������Oe#�U��oi4���A�K�Ne)a�v
L�r���I����N���K<����l�fL.�{�^w�T=�5�Gnba:��LM>�i͙Ố%Ru�|3���䞙�����Fp��Y��9�ю�\G������-����ƾ�	��)�m�K��1c<6�ص�ۨ��`���o+34O�z*�r����~~�DTy��&�|���\f�*��l��V��y�z2�T�$6=*�x�$�#�y٨���n��	G>k���㵤�2��,o��=U��J��:Q9����K�ў������f�[>�O3#�s2�=��^��^Gjp�̽?�
�>�]_��]K�}�{����2V�d�;��z7)�Q�o�<=��Z�
u��}���]�q{pU���w��#~,ǹ	ZnOx�يȹ��.3�Zu�3������H�{iq7���L������3�s�ױ?��Ƿ�H���j+�V'0�I��3
��������r��~��{�;�}�r{�x�Kya��G�R���y�3�gE�<Tŝ��(z�λ�y3�����:$���V����3�t}��1y���}>�]��v��?QE\l�*�����諸��<�+w��y��x��0q�(e�mV�<�h�ʲ��Mܿ��2��G1���b�$?���5E<������4�{³�Rd���+���wU���w���NL��z�Q4��%��nu�@�
-d�J�ҋ�o�,���Ծ04�c.*��
��Hr����s���:k��5 ŋ4)��4���<\��\�^Gz(1k���1�.:S.�NU�X��1�mΎ��U�S83���w��K����PGHe�wZ�5k^C^��p��}	ɽSz�BYA���� }��=�^��垹�*7t�^H���u�b�s�:b&	�j��
V�z^sF�N�
yf��=vEl��K*�[�͵���W/�V,Vk%`�Vw2n����$����+�t��	�Oh	+[�/�TE�XY{Ϻt�2f@:� �����C��W!��F&��@��Ա�YHN��6��޻�\{�.paOW�
�m\��c��:���'sr��]bM��@���<�&,��g˾�EY�5�.ty��bķ�u�oyܹ�O��r�(�Y3ky�,�(uw�^�_mY�Y��e4�;9yi�}���MYEU����.�귺\�vZD��9ph+���=E��M�d�!8�ڱ�4�Ø�i{���ܙ�q$�������!9����N<ʼv�����^b���n�s�r��.���.5(V�c���T��8f��;�Ūh�ps$�]�.�F�|c�5{('��sk���3AF8en��v��v>�ww�BA�edt�Ir��8��/a87���d�/(�T*_��vZ[C%�2�!8ؼ�y	�u�V¸��0��	�I�X�}���^81��bN��`rjͭޮF�~����!�J�b��e���1�,��F>@�9���svY�±����(r|���z!�A٩��C�ѡ8J6B�؆Si�.ʹ}"���q}k2�
w�J�B2�J�iI'����݊1ӻR���R�!��v�t{��0����8�Λ[ڎ���%�?�о� �60]��.�3�|�����/hQ���U�j"��U����w+<U��]�3~�mP��*�l�h�=��A��@��'u̲B�>������=:����+x�0z�{��B�3oF1ǕҬ���y�u�u/�1MX
����D���2�$��B9�sfT#M�ǟ�ݫ���y;u��6ܹZ��kٷ�bmR�h֙��;�S�n��N���Wu�H��u�6�o�ָ쮦��������Î�Ў��=۩�������;`���x(��f?��U��f�\�7�S�p��d��p�s-w�فٔ����-$�H���}ݡ���>��,�h��dQ��+g�"KA��m�aP��\�4(�ƺ�0!�6�����9k}��8���T���D�i#nT#\�]ՊA�Kl �*VE��#hT��j*2.*TR,-K"�+m���d�Y"��B�V�+"�	U��
� �J��m����Lb�h%H��%d�� ��"�V)���DP���jЩ(¥+,��Z�QJ�FUҪ�1��p�`�Vҥ(ֵYTj[am�-�IZ����m���(���Y-kl-���U�PA��V�P�R�����%bȲ�PƌU��H���ҡ1�\��TAB�V
��ł"5�����YD+Y��Y �YQDE�B�@U_~�/��FZY�P���}���e���%Zh�!�N*)Ag��eh�mZ{cRw���e�u�tPi�u-�*�tv���������e)C!5�^9�1��xsޕ������GC�,�Ð'���D��:jF���@V+7��m�w芯5+�����n�z����
|�_��봿�DO�����'.�fǀ���l_zY�}�_��޸�t*	l�o�>-m���؄��,8�	�������ٻۧ����ĩ�p��n@�٨&r��|W�aȂZ>���¯��FA�����%�������-�MO��wu ^{��ʙ�Nn@!�뉐�E������ 4s*����٥zbnsNzQUA��{�P�L���W���=�@��Q�IC���0P��H*v�Ïg���]:ȯV}�q�9��7	��m����,{Ju����䚷>*M��p�ᑳ�11r\���w~�����ZdTo��93��q�ύLwя�ǜ�RL��tw.�o����N���{�\M�uE�`���zMGs�o��Suc��>��yP���Gz���
��L^�7]>C��H��THzs�v�z�LU��M�5���=~�Uq���Vr�d��-k�!O�п���5���75����, b�V�������K��gT�-�N�,�.����ńaŠֵG���WYV�xjmb��nu�]�K]y�d�M��Wy��>\.K��r�YK^��t'Y�yM����/`��f���E;���,��<���_~+��ُfzai�������[�,�k�����Ch���j#� {�D�b,���Z7��Ck�����t��^��#�n�\)��V/R�5#�y�>����`oNw��E�{0jx����N`���A~]�C%.p�'�P�^x�Cc��lJ27�3�1s���Ozhg'>���/�i���?b�}�E.}�H>QF�h��j�=�x	��S���G�FL��t�Ϻ��q���~rі^�����ʒ�̺���/�~��`�v$��uL	��|N�L���{�^�qc>���yomyFέ��)�&ցt���W�\��+�=e\,�!T�<z�1)Wq�^�>�(�Λ�6�	�9�%f�T��{�S�Ͻ�|g��4S���3�;D+% h	N�^�z��y�f�}�2���v��9ޏ{���9
����#q�\9��~�B��~���\�\F�&

�/�z`ԍ����Ž�Q����9���O�m������o��������۷!�ˢ���`�T~-x�v_���W}c9�2���+麻�mn�ހF��7b^��V���@��Y�L�t�P����� �j����k_MۙE'4[��k3��r�VR5�&�mS[	ι� �3��+e���4)�5 ��{���I\rcp�;�u��3�9�;ԥ�LBvү5鉇1R���N�������F^���9{��f.#�W�}����D���U7���o��g��$w�lM�>���LO�Ӓk���
�ۆ���o�aU�{�~^�u���e��Ղ�¯�t��t��r���(�8��^V�y��5���U�����sꎻ���3��$��u�#�ޠs#ý��d_�$��2�h4�|R��+�<~~Y�m�p��+.�=���L����~�e�g�T��ʠ�����=��N�(�L���D챙!"UABr��-Q�mD�y��M���9Ł+/�Nwǉ_}J}��~�q6�5���������̱}sc�0~v�j�Yyg������`u���8���{��n;خ'�����Nk̚c��r3���M��v	zn$��|/c&��q�;�s����}v5�2G�ޯx�:	��S�z��_%���[�v��F/0JD�Y=�UC�WLa:�*+n�<�f5����I�|`J�k+RЈ.���*�=���E�!�_��H*Hc�T�0+�P�2S/U-��>ڬ�ߟj!�����V�/`J&�T:�	���y ��8c�3%(����㚕I�p)�`����sN\#�A#�)8D�Tݔzߑ4+r���w���܎VS���a��t�sh���I������
�R�id�����v��g�UC�����euz�<��[�����%Q��7XnV���sQ�ɝB������E�f����\{�6s�%�����}�����e�e�)-؇�'=�����9�.��_-q�Ǚ��] �-��7��1��2����_{-�8�4�24P�>W�K�^Q��0{�\LL7j�a+�a͗K�v:|E�Z�{��H�����3�Ǒ�UFv2�8�o���ofD�����,�Z=s�(�ȧ��9�����~��5Y��U�>�o�'o���ow�Շ�l�p/!{؀�F�Ɗy^�@�L�z����bi�m�w�P��/7�c��󷜢���m�rF�>3�ޟP��Mh\{�l��~�����[fl1כD.���0r�=��ܨ���q�/�ҕ��?Y�o΀�9󭻏1�$���\�L�.>64�q�!��yK��X�Bu��N�5���5��7ٙQ�UO�.5N�o�wc&l��s�c��/\/��8��:��Nׇ�3kG�2tV��s���`TG,�G�}�\��/P���x�>��[��xH�(��s1/͹�.���;+]�����W���E���֤B4��b1uZ��}/��C����ΫC�z�|܂��=x�aw$`��kt�t�+����x,��m��&��Q�*�����R�I�[�m��r�s$��)Z�h��Ro/�L���b{Mğ#�f�W���g��@�_m�+��z�$Z��}��9�����p��|����>j�Wʐ�o�֋X't���uT<5[P�=]d�1��=5���ʽ�+6<����??z�MǶu��^��e��;�i�̒��L����(��Wp�u{Z��n�e���G�m�yoO�ԩ�G";�Q����=ҼW{�e�#q�;��RQ��z�����B$��Aj��j�X��d�Q�ɖ��!����^�����=���G�}���mu�(���C�/�ZxT�d%{)S����޸�`LT�����6��G����1y��ΏC+
���#$g����T�|�_��������uWV�}F����Q��l�o
�{���Uo��G��06�h�+�>���].��u(��³���������p�����*1PW�aωh�2\]�+��z��^����Q��[��v==H���~��PϽ,�z�yK���QjhTA}^�1#P�1]��n�8������u	�y��>�^+�NW����=�CɗJI,v���c�ϔW�N��a��9��NLxf��{2�9��X!P�@�ו�m��x�e�C%�:402lg9n(z�,+�����6EJ���� �W��Q;&=�'
X/wf�Ց$�Y�Kֳ�����Mdңt�Ô�:eME�=��?I�i��r2�sBuM`��dڋ�H�G��3�#�T�)��{��ߎo���I߽[@;�Lӟ�2����Mz=۷�\M��M��H}+L��;�Ћ��7f����~t<�"\��� GFϜ��8���ݹ�c�zI��rV��>G�蛨���/�I�s��ζ<�sD�W�p���W�p��{�I�~��7ׁl|6t_w��7_��v�z�L;�6�Ǽx��`/���\���dY���U��G����r�9�ꄌ��5���x�̴t�ó��w�U�մ|<���ݮ��;>N�_{V��;�̣ި��:�'�p+'t��q;,by�w^k���"�m�]��mg��+��E�G�;(��s�}��*�SU��0}?+W����'9v1Kw���伛je�]���7�'���L\N�	�Oz�j~���Ǐqc4��w/��4�b�ks������q�[%��XwŇ�U/ӲP{.�(��py���{ͭ�yM�b���=�Uۜ>��/aOz��'s�7�al�I�*n��1S�����0���yz|>�O_�a�]؅]��N�,�ԗȎ�GavklU�4k�,�72�sw�T4gb�|;�o�ł�F��v���Z|����������ǵ䛗����5!�w�R�[&�-Ȉ�x�ޝ�dC����&�:��5�9�����pvD��biF���@�_RH�G<ǵĮ=���u��b�
��;>rM|O޹�bb��M�^/k��H��ST�W��1������zR7��>Ϩ��_����Tw�!�������Y��hϥ�?I���wg����uAE}Ҹ��^��C��S9��wB���E����I�q9�ؚ�%�8�MK�ź�!^^����N.�����ȓ�^���q(���/�u mf�!H$tk���z��߲��>��{���g�po�Ҵ�B2��'�adO�_�3���/L�x]��&��u�<�~<���"Ec�Ǚ�����0{�elSU�o\��B,gC�yGGt��Zu��{=Z����ϩ;"v}�"��}�w �^��ϑۉ���[�����_iz}O,=x��{p�:��;���H�����3,�{΀��s�c��+�蒎\L���y���o����aL4�j��)�!��g�P�i<��m�W��$o�{.�m�=�Q��e����cF&L�Q���t�^�^~�
�'kf�J��7�v���=�?W2�C�s׵�ʜ=�Ema>�`U�Y�����kkѭ^�Q�:�1v��U2��g&�s�j�UJ�OTa@;ۉ���szm\<����*�z��ITW��3�U�Ix��PR�ȫ���ӽ�9�m���{{\bp�5C+�Lˆ��k��;+���bŉpW�iW[Z�%��90��٪ֽGu���d(,wl�$}������K�����/�/�_��o��������7���_��� �����Uy�lߡu�#��wM��,��2�kKN���5�s�X�}^� ߙ.��������m{p羾�p�����b����,�ڇ�X���ɝg��m�'B�k]�O�w��=;nY��{���v<�^����G�و1���a�bKM��0+�P��Ꞹ��Y۞�+���9��Ǒ��y\{#���r7��Kb�~.%�2 ��g��*���,GsK��+=�Ǐ���B�|��GٳCQ���=�B�6n#�U>-��>�D�W��VT���~�1��/�M׀Z}r@���#��o%�3��Q���m���
�9�#~���G�Nz��w���~���ǟ�� �T�GV���=�bʞf��D)C+�U�x�T�A܋P��$�߬�����B�����j����baz���}�Ih��TǼ����>����5�sҊ�Ul�r�I��q��"�W��9��G�dƯ�bb��vJݟ���,���]���4ù6�/������Ɗ/T��N�l����W��@���\�Ĭ��?3q�~�hk'%�&�~��ŋ �o}�b��}��1޶��-��תe{��Z��UGeC2T�]�t�e�Q�n���g�׍��t��� ��M�V�Et��6�*Ǉu��V����~}�������^�&���]�)|m�5��h�)�}�n���ԓK��/r:eI�jn�ǳ�;�^#��s�\fօy:��l�i����n!�ˏg�]Ә�'O?;��J��u[���$��/��u�Y�������D�x~����:'��5�lW��:���N��e��t�{C���шP�;w4'�G�nt���n"KGo�ڇ�>�٭7�@�_ݶ��S�p�\f��޸�K�-������');���BEF4kE��N鿤�>YP��FV�<��7W���p���o&��TR� �ܮ�uǷ��n���l/Z	z��4���%��cM�<��[�+��3s��r��F{�2�N���w����>�O�Wl_�7��>z��<�d	Z��Ξ39
I�+���82��E�W�+�Ꮾ��|���N}���9���=��7*�����D{#@��w*Z:Ƕ'�,�C�'����T���^�y(6n�H����C�O�ё��q�pe����-������kW���-�g�c�v��L756�R�K�S�IΠ�ZC&-����w0l�{h�r7�.{6�
m�8�>5�>s����ɃjH���sPZ+CcZ�s���2��A����.B!eM!���Wf��W��֏��� -�����ǤWU�5Ke�y�/�Q
��А_q��b����W�T=�=
r�� d���#� ����@!��{T��|W�a�%���yt��vg�qT�*�,��ח�C�=Ž�z=�F�e:��jy��L�ٴdmmI��-P������O�ze#ݰ&=�Q�%qE�~����=Z w�DO��t��a��Ϗq�1�0+(\o�u"}�?Q����wNAR���1����|M��.r@���$��O�=]�g�`�^P�k�����f�����H�\�2*#\�`]Lv5f�m϶�.9��)I��wu��8�V̯>2��`�F�&���^�/�����+t�>'��:��=�������=��p��4��EeɟB�;>OjǱ��w�VvK�;P�y[��׸�w���Q���zTmz7�b^�]WG� �F��؆�{�S�'>�П��b�����t�-�90��F{����{Y��9r����x�=7��-�~'!�y�qz�i��uȿ��Z-d�:K�?DO�麔���u
��"�G�1��(�o?fe�B���Ѱf�p�f=+"u�E��Ď$��X3"��<��:ݬ�vs���3_ܮ�*���Q�4�{V�@�]<�r�71�)BDJ3r%�GӜֹ?��+.���.,c�L᥼7��2=A��X� ��4u�)��6��Ѵ�Zc����TP�bK�*m)�7U��~|�*���)�V��G��7��O���Ȟ�
]c��h�iZ�\E�W}�6r��69�*q1�>9��[c��.���u��08>�Ož�Y�P���aF��z�KV_r��1�<Y��r��۞~�e��Ӝ׋�[�Y�ŀ��"�3��W��鞵{o0s�|���M([h�]��}�9�%�꽳��p��|�*bSǂ�KJ���? �]WP��Y�#[[�H�I!V�]GCql��P:��8�GN��l(�`�C'-)�w�`K��Q>���%��k�G]�k��)UCv��F��`F�I/-W_�����ʱ�ՙ���3��uh�S�]9���5������7�z�����]�ꖁ:��t��tnV8�yA~#���|�L��_�ޢc n�r���ܸ�f�*���E�|��1'�-G39��}ۣ.͗)���-2n"E@�qJ=���+x�G�lY:�(5�L��h�����D�-ݭvn�Q�k�:aJ��t�[])]�^;�X+o�x.�׺p�-%�V��G8��>��^��&���qdm�����
�|�eɽ{mE�)˾.5�ջ������1��}�˗ݴ��~�O8e�*H`�Koj�Izm�fD�|A���̘e{��9h;tՎ�k�i�x���uiSP��<m�k�Q�|��	b�ofD�M7&^ht�N�m�*����عf��x�qbKw�p����{�Mf s�f�;���u�'H��k.+
�SL�cea{��$�m�V�`L�r����f\COQ�\�6�f�o���V'[��¬�����A垉�-+�۹vR{ӹ�|mvhx�����V�&������ԩ��\�X[��95%Sm�>l����Ų`Ed��W5/^�o"/2<�ʛjdv����ڇ���͈�]3dZ��sdu�|�V��-ʊe=�m�w��t��g�,]֌�ǝ5�/I�J�z��Ӈ-[�n�+�D�d+��!0.��hήp�{�Ĭ��(���ӽ��^������Mx�N���u��m���~�oc��0�[��M���������j]<��4�nP�N��.ˎ�uQ����3u��
hS\x.-��a�F'�%��Bw� X{D������g�Z��
p�	�<t�/��_�gS2�6�2�a���훻��~�xĴ��X�P�PUAAH�O�UC-�e`�����+��Q�Yl�+m%����Pm�
�Qa�U
(�J�e�m�ciQDaR�%J�
�ڴ���J�UY���*
E ��ETU�R��X�����i�H(��X�aT��V"��V%aDZ��jQE"���iQ���cJ\���#QDAUEV,fYPE[k#�q"�-�UQ"�*�Z5E��E�jR�h�T��X�Ճ� �"�Z�J�iEP�1d���H("AX���,X��T�����(���**�aYX��d�m(�����3�+
 īlm�QA@E�P�Z�
KZE������F�*¥B��������r����)��[��x"���U��Y��,�����6����IaH�����hf��Y�gF2z����=GhE�C:�S�����W�.j{O�o���|:�z�M�s)w�p����F�Ѿ۞7.4������0H������>����\�.���2kO�#&w�\��Oz�n'��7�~=�b��fcI{}ꗐ3vrnoGl�l\V�Ϻע��uύ��R7��`M�x�����]�t}Ψ;�l�{E��=g޳0��ܹ@^�9��~�q�R|cn	ҢO�SqT���G��aL�{w�Z_���{'�3z���}4xy�;ё�%q������� ���v9��'��_�P��t�{�;=�>W&vcX���]�j�^{�X�M��	�]��#E?_���^��'�nD��Z��2.{מWr�T�p�u��H�낍E��&�׭"�J<��D诽����W��X{U&F�J��@�+������D���FDKG0����n3��I�V�@�'�~���ڥp�VV{'�Vx�w4���פ�n$�v�ba;�NS��чҴ�B2��'�adO�_�B���aw}'��ս�Z��&}�:�� �<�ID�Ih��M�>���LSS�q��#��Z���]���m�ܓn㱢�kG�+�x����;`b;X�`r�����@�U�u㽯.4��E�f� \�ns�3���)w�3�{x��[��p�'�
[�Q䖛#���*����Q��VLV�>��$�GjwJJSyW���!����ej;�*UAf��Y�Nij����o��1I��f5�dT���}Rx{yU��])rpW��R�� I�9�M�>���==&����ъ�vE��TW�3Ԏף���ߚ��������:h�^�(�����^*�ǽ��+ܙ�:�Ϝ��W�:��>�f�����wu���U/��yT;�e�{�����r�'g�#��Ǝܯ$ng���蝝x�C���ٸ���8\��^��zuM��i�_TM�N��^�Bs0OO���j��|�%�(��;^FMiW�O�i�r7�v����<�kQ�s>����bf��=�|�d��������ʞ1аN�/�ES_d֖/���t�~��k�
��u��Z�GW����>=�\�U�|{jQ��%#q%�=UC��t����\��KN2��/c�U�w��؍ȏs��#}��=�Q.���
�D��,r����ܓ��V�C�󻃸5�~�^���~)׺��^¾^���{����s,� k(a�m.��a�]���w2�p>�����X�n��#�l�K=�=����=~�q�����7�ᩄ�A��Բ���2�9,���)��zl�7+t��{D.wQ�pؕ���b�]��#��o![2�<R-^������_FĮ���v���`ǈtfR#pS�U�YXޜ۩׭��1M�CN�!���x��}
-��Y^ƾ= s��t(�h�,y�Zݐ�9Z�?Sf/�G���x�_b}g}�'�T�ˤ�<4���q��'��0[.�ba���Q�%x�9���s��ʐ�����}f�^/wv㦽\X�����#�Ƿ2$T<�7
Gzbaz��14���	h�ց��5�9�tLc��(���_�yc9�+�P*� }�����Ƹ�l� >5�`d���{�U��bF�$�n*��P�;�����g?*� {S�����M�_[�I>���YC7�O �퍏4]�ċ�$/[��Z}��R/O7f�n9�d���P��uQ�x�I:s���}76r6˾�����_��n`�F�ࢹ_����cL�B�c��fG��:�s��T���ʚ�e���v�M]��8^�v��^'����x~���댝�κ��m0'��#°6p��'���~yuU��^v8��U��u1Q�;���lN�<��+�X�٭7�@�(�w}Sy'%��7㏂'�t���>�������{m	���`��r^,����2���Wma5� ��LƲ�+�ss�p�h�yR�º�����;���*J�¾ܺ	�^�&߅�[�)��w}���)\`ֶYӍ�Ļ�K�g�&,�#F�Fx�N�eispw���9(8�觼�RQ�í�xL'�����g��u��t���;_���{'}�������ݞ
3��2��W�@�K��m�Øg����7w
�&w��r|=.�3����Do��+��q�o�=w�;�R����=��s��߯��G�e��A�U &/�øɔ���K����~���||=ⴿd��\�"��%��t�|�_z.���U�(�N��*�S��p��P��G��Hy�S�tZ}�0�K��޽Y��n��������g�=�mK1��]�S>�g�xW���������6jϽb{=���H�л��d{��elt�����g���CsD�neI�+԰�����W�"c޼�
�p)S�s�����29ש#��u ^{�����wB߫�p�9ޙ�>�=oUf�V��ܶ��=�����Z;�G�}��)O�׎zr����q�Z*!�S�&,z(��u��e�ZR��>��(:�tD�^�Ӹ��9*|s��G_���L珤�*�=����F�q�wS{ؔj���<O����;c=D:���E}�wǡ3��q��x��T<=^���~L�V�~�͌MP�lg�hz�=��Dv���V����ם�YӶ�'}Ʈ���n�G,_k�]�d���L�0YX�ॊ�?n����/
�j{��㵕xq��fb��e�/R1q��#�Cj��zun���_�����]�r�i,(�:��՘y
�úO��f�I�����$����j�K��|:Mk�k��ǧݪ��s@�G�3Mg�3^�:=�qm��7�V<�L�7��	Xn$�;N�/\FV�f׸��>������Lݞ�
}G������w��3/d��*#���H�^�Z/���9s-���xv�xQ��ΰ��z�&���i�=7��{��^�jND{�MF�V��=5��IӶ���y�A��"�◖���������ۇq�����7Ӝ�ßz�M����{���b���:>-D�Ks�&s����J7�e�;	�`��/c&w�\�S��MO��V{���B�+�N�)z�ŏS���juh����y��VQ)�N�,
=�����ۺA�S����]_]�{&K�Y�ݝ��I��c�*�=�~�"]���~�Y�2�I�*n*��O#�n0�[y�^��ߪ�Nv��r*\+��ؑ�z�g��v�{��Y>�bhڧP�!�u h�0����Ox�>��ǃ���F[d�h�ȏu�E纣��6r=�|�{���~�S�Yy�!��7O7���Y(.�gq��T�7��+����,�tOu��K�k��׀��|�^�鳗>���2R��cO�x 5�jQ�.��bk�o��h�緮iS�Ӳ�_f>Q�X�nc�F��+�ؖ�y��P��_u�oP���d!�oS��j��r?���M�Jc'��s����ĵ^����:�gc�pO޿g���c�F���ap�CI�oM�E��P\����2S���I�S�^��%v��W�ᝓDR�B�Č��&w�L���j�ND��0��H��s�:4�V�P��s�:�+�ᘮ�������Ϯ�c��V�s>��?*��פ�7�����C����û�n�{�:j���N��zEz#�W'�n��#��yND:��R^�Dϑ�S�+t�mL�ׁ�K��(�ś�Ǒ^�(.;^�˱�3�B|+ΪY�{��}η0xlzw��d�{,v��9
&n���\�_��\P}y�a�����|x>&z����w^��T��ʠ��{.���N����"�q�N8��g�{�M�N�x�C�����K������/O2��͑-x���w���^��sk��5�YS��Q=��҆�N��t���
�q�F�o�Xk�x��];뵗���;2�S��b����7j�{����`����L�vg3�7:�w��~�%)Qsc�qv�pŲλ��WH����hd�λM�˕�I챣^v��wU�pǲ蝺,��|�P����U�'ڪ�F�j���N<����)��h��;-esҶ1)����s�k ����.�e�9�&��l�uU�rM�a:#��uZ�L�0��{Č��}�S�P����u�1q�%#q%�=qUƣ��+n}���p��m�K�}apv;��}�*����܇޿q��z��z�ÔK�CFC�Af��$0�����FEת(�q]���J���d�}o����:��q�{NF�[)lC�d��SWT�ҫ��܁�SxEH�����,��=鿨�&)��7��w�}x)��~W��H��>=�"O���Yn�<p�b����#w��zN����; r����M�<�b�:�V�p߭��et΅������BI�ԢD�4�'�yn����^��D-�0a���F�^++�2#]x5�d}�5E\��GWV'U{>B}=I���7퓥\G�.$W���,�Z<`��J&:�W���n'���c$kID�.��B��~���5�9H���;���O+�hZ:HMd�����j�����oS��=�O����wz>
��m����y���z];j�TG��ȫ~��y���ǝj��9���;Z������͢E��5������٨ێ~�f�~t�ϝm�z��_�g����ܾC3��ʚ �3 T}���gP5��]^\"�-i2:M;*�Wp�!��lY�١F�G���gp���X�tH[���B �q�ɺ%�(��1l^��E���D�Y���+�w`�)�E|�˪�
����:��=�t�+p���ܰ�6�;����c���ŏSy�ϛwu郒0�50}Gk;��j���>]�q-I��~eaI�;Nׇ���>����\�k��`M��6	.r���+��o�]]O�G����:k}�bn��L_��=������v���W��y�Z|w|��`˹���\��{�_���l�M�?_�ϕm��>{��X;��gܢ��Vl��@ɝ�����޸��_��N�Ϊ}���c�z�MǶu���� �{-�{�!�J9�h
e:��Ϩ�k��B.}G��خ�^L��r|9N�7!����}⺦1��{���f+}���3���Kr֋P�4:Ф	ue�_�L	��ø��N|2]?>�C}ON|�>�h�׾��d�����m��c��6?	��)�c=��۽F�z@�]SjyzM��H6sjtz����ム���7ɯ�ã�x�h��������eK0�'�H��Q��l�p/��z���z���Z�M��^"��m�~t�����QP�~�����P��~�t7uJ�o�k#�y���g��D3P�Xe���u:�40�d�\`ᣉ}�h�^;�T5(ӵ�]��>qϗ�=&�x]�����$ڭ
��W���qr������:4QS�9��h�RV
;8c�V�����t�r��*���9WQ,ƅ�S�:0
��J���ȁ�z�{�D����:�R+��@�~XG�߯�}��w �)}C�ǽ��7v�"v���^�yRÄ��p:����QG�]��NW������۷"�P����x��s�1Y��i��m��mt�L��n&
ԑ����wN/M�O�q���W��g�VJ��S��}~Kvx
�ٻrME���A�#�t�^z�u���"��;����ݛ����ע��6+����~���o���f�}>u:<�̓���+ND�#�7P�N�v|6J��:
w��R�+I������WP���o�h�]뗑�r�/:��gjA�xJ�q%��څ��2�L;�l�&�^ܥ#�_�}g���ܶ ��X��<�����9�ꄅ�3���x�̴v=5o��1�#��7ʹ�Q�{ʡf���/Ǧ�;m�)n;�9�̣+��fG>3�}.�7��
�lۦp/Ǯ6�i�����ջA�K�V��]sN��x�u<�K�S��7Q�jp�5�μ��F��-�R�]6׍��F�^X[p~x��_ؖ����t���U�ϓ��V_��`^z|J��	�ڪ�.��n�N��=�=��S���z�t�2-~+q_)��0]��R�#���X�I��X�p^Vn�y+m ?��'�kܺ�:��Y.�g�(��Uk����uf$��ZT6�F+����.Q��Yʂv�ǐ�&:�u�x��f��J_�a9��nSב���pY)�s���U0&�X�ķߖVݸ=����C1�Okr������s6|���I���8���7+���>0�6&Q���3,	<���[[�.����~�Ώoж�<�g��>�z�dF�%q�~�������v8�D��Ǻ+�Bfr��*�J@r�z:�o
Gې��O��#��>�x�����@`������G��<�F���Q�T2�]��K��}�8���4*t�������AE[J�n!׭#��%�F�'D��;�K��m��-�qw��˩�p ��0j�P�.|�di�ޗ�W�&�[Y�={���_��8S+�y���?!�3��ۥg�T����JH!������E�&�����;�#,mtWC2�[��Hg#���6|���+s�)zg#�;\{�pjW��nKGn&�d���j���\w1V���u�!ʡ�3}�^�;�jN���n<��'�"���ǎ^-�K�}�_�u�1j̞�4$l�s�˺}1��3��JMiZ}W�W��۳^�U,���<����g���Q�߾�[^�w�;3G���%�)EY}��ύ�;i����pu��n��]EFVgj�;�����zoj7�r��p�u#��fV�z)�z��yr�س#��`6�m.��yk�jӗ�Kr9�4�ڐtY���SҢ��])u�p�_,�.#
��-q���h�e���1���Z��7��Ԥ���g
=�.���y\�΋7��4�f�!BS�V�
{e�qx0:��ΰ��.Y�>�,A��uca#�@�9T7{hT|2�o>���f�q{)�[<a������*g�Q�ynҭ��Z�n�`�nT'�����0qS���J��(����(w�NZ�3pv)&���V8�_mf_�op���S���)˹��1�!W�<;OT���jf̋�ˆ�$@䧔Ɏ�u�0-�:F�5k-`����-�[��t����jU-ӏi�-�6٘7cܺuwc���H8�]{u�=�j�4�*f�S�]ޝ��Xmh�5`���2q���pb�"�V�T�q�]���n����n�R����96�����+	�%�8�Oi�ݠ3�	sn��-��R��1 _�[t6��ӝ���G�y����9�aۇ����.���ő�A[S��l��a���t�S.`��2��n�yݓt��w������yF��9�wSѕ��o+y�iM����To�����a˽2TǺ�4;���u�֭�W�,���Hƅ�yN�y�U��<t�{�8� &���V{�]��q.��Q�^�ȷ�D�^.Uw��a���)čN�c�NkD�p�"�J�l�lU#r��;��:��f�%�>�ꘔ���������k�⾈0kA�4d�m<�[��]�%��x�x܅�?���ƣ#�'��h��{�^	�av�8�ڻ�+�d��M��/2�=���Z7KAg��n���9N,yk��k샓�qf�,�Q4O5	�Ϻ��{�I1Ym��}L�T�F�	6��4��} �������#Z�v�A�*
�kb	(x��1�j����2'�+6ahr���$��V�������r���9��\HfAt�L�ݜ%=ӷp<z��wf�Rv�(����|L�U�|�����n|to4_a����ݽ�گP�i���!�ȫ����8�n&*�`]2^6־٤�ܬ2V��E�����i�ȼ�2<�S�;���	�d���GEg!���'o���lػ����S_P���.]�]/�f�&��6�S�J`��,o���p�
�ʷl�|�.�	��\ k9��ɹ7zy�G7�kϹ9;Dy{x��G�{H˲�1������-���Pw3E{;w�zEe55����4��HN���Xޝoy��u5R��Ihq��ٴPT��g�7J����oʳQwV��{jGF�maUm�f�1T��ö�����췕�FRX����pn���̽h�5أ 9����3j;݋w�����\������ �Q��T��U�*J�V�# �dPcAX�U��5*�`�
,��ZѐXT%�"�(�U*VJ��*6�XֱUV(:�+��Y1-�K+X�1 ���dDREDE`�H�"�*FՊ
(2�P+D+AH���bE2*��U,QTU+D��c���X�TQ�PR���Ȣ�ij��)��V
#b��&X)kW(�QEU+*"(��Ŋ�X�#"�"�(��QF������n\Ec�ATAQUF
�`��#DL�1��QUL����UV�����9A�U`�(��L�-�EEE��V��V�b� �Q�F![DU,V1���)�E��ܸ������`�"5��QDX���$`�Eb�TQE10*����,Dm#h ხ͞+�rصT��.~B��z�*����egt��9J�[t��-��Jъ>���}�9ۈ�It��[W9:=+���g�՚-LR�W���q3{P�S���nfY���j=�ndJ��nH+jLP�Ȼ�y�Q��%%a؝�2�8}9]:���e���~�e��W�2cޘĲ㉞�oN�؟>�����NGǧE��Pۈ��2�&���'´�k����w����q��<�U�mM�P>��WȠv=��n9*��{s�-`��Ix|��������d����ߔ��%еx|�Z36���k,w�}�C�=��߭֎���;��(������'��~;�KT�[��u�����Ү����Ee.̉�u:1�����F�י��
��8dy	C���:Ȭؚ�Hm����x^m�z��F����ʡo�+ž���u�q��8���7��J�^K�lNDّ�����]z�x���r����C>�n��[١(�o�"qz�7�>+�s��8;�����I�z��'{}�2!l�/�_A����ar�7�Ǚ܈�@*�����z}V�tϷ�j�,�g*�LǗI��t�5�p���E�����J��V��o�}�3O�����V~W���:�vpj��]W�/^wI��G {_����݆��G;�2�k3�'gXt=g�j\��V;�3AUpx��{�V)x[���r S9+r��z��1d/��i9�:C���
��)�ͬ\_��fP�`G>E5KO$2��t�m�#�s��k����2���>�Ckۙ�x�B��h��10�r������{���㰱��|�8��i�=�w����M�>U~9��@��~�������D�G������|�T�2}�&&+�m�>���
��o�pt?*��S�<��?3D_��W6�9���{��$���͎�$z�9%f���(<=٨w��l��<������
霵�.9N�z;��jI���I{�|���l�}�^_l��eqc���z�����3{�D����LzU<n>̏h��7~?�zr$�����ד�}�D��s���y~	ibc�/6�yL��P�!�Ӯ�9�w�4'>���L_xOi���ӳ��qc{��Y-P�£�ׯ�.��s>�7���ٷ�#���h������$w��օ`����K�}wl\����~�>r�C��WTm�*�7;�^}��f;!���O��=��WQ����G{�!���R'=��r�5;�[�z&X����U��=q�;鸜��GS��ϓ���}��x�����Gc�����$A�xp3~��*t\���+tbv{�=~�W�-��0U� b:I1�!+]gEȉ�"uv(G���FS�0����_�¤H��A�ڽu%�޳Ѽ��W�3i�j�숪X����U@E���\}���knL��S5u�ݵ�����dl�(=2���\;�ڤ�ä��W������:7��Z{�g��~JyMJ�w����"R�����Yy��x��ڦ������A�p��G���W�1��R3;��^i��u��t�����w�p[R�s���ǤW�z� �D�G��=1[����x��?<��Hp_{Θ�I�ӽ�@m_��y��_�F��O��J},��>����Q�Ϗ�]�"	H�1��U�[���u�H�{�H��4T{-����7X��<����(�j��z&@�j�Я����	h���T?^���Y>V�ߜ�*����j�Z��	�f��뗪�7�Fw����Rng����TE3�r��(�zS����I�w�i�Ə>����0W!^�='g$��ے]_���J�ڷ���g�G�U�������)cn����~�'ֳ���o�WZ�����BT�2ǽ�u$�>%ῤ������k��^�z��n&;./�ǥ���>j�w�5'þ��=�"vW�h{��Ԃ+�%a������B�D#�o����D�����}�Vv�WHi��K�g!���+=�_�{�e N'H�O�6���EZ��w����b��`��0F�#|�_bۭ�tD`�5ԞE��\��1�n���� ��L.o	����tbS[�����h�/��ӻÔ�Y}�j������p3{L<���UO�N|��~�]������X{x��W좏�$(UA��l{��ߢv�p�guG�fp�x��� r�w�r��G���g\�*N��������$�è�>c�$��3�������W��sN�}9N�;!��M_�8�u'$�X��-�I.Q����R�dNC��*�ӃW�����؞�]b[�U��1<�w�cs/ނn��l�{�u=�R�Z*}`��Gt�9�<U��\�xp��˜���7=���οL��o�*w�[���@��C=��{ j������_��7/����x���*n*��J�p����͹�����'C��*�?9�#���^��D�=����� �AZ]�d9�l�U� p�y-M-�)��f�R�"o
�z�����������.up�Q���� {���Gk�m��+=�ez�PO�M�zhQn�7�MwLj*�W�ԑQ�QL�����^��>�U8�l{���~��S��鿦�U
.|�d�Ә�����n�viҔ ��E�1�/N09�1=�{{N�|.�k=�yT�s�"6ҹj��S�����n�]��R�`m��)��&i2�(ܨb���6�׌��ӈ<�ô�wD²Qx��~�:��+�
����'\�%]�0��XGgsr;0eDy&i�'�&�q��P�gۇ�3�J9	��>��n�SʧECGzbaz��N{�F|}+N����o%ڰ��v���\��=�}�%D&z}1�����}' ]����(��-����^&�g�z齾��^�m�W��������7W'���K��.N��ːE|��H|�e�۳B��ʆ��r
��9�OL;�]&�4�O������ׇ���� {��P��)�DwW�]u^u���>w�q[*r<p�67=l6o7j=y��7��3Q{p�n̿��x���۰��˻�(3}��{м�T��J6O�aS��_�����Ɩ=�=���{}�齲ra��G�6=��]'�%#MouF���s��O�S��fj����X){m~�78�ܮ�1af�yׯˊ��H����Q�}��=�{�޽��
��$;>�T�VMi`r�__�릳�=�㽈��Sv-�^��|�
1�"�W�t������)���w��"]��ⷧ��N���� 9C����w�3�1��tӳ�>��9��y���W���v���2�02��Ц��2Dm�է����H�<z���Q��r�`�(��0ѽ��^cOL��=�3��;>?s�n�o������5�Tߒ9{�J�ܻ�_=n��Hu��9�.�w���y	6��y{t��_z,W�Y�p�%�ah����'�7�Vk�!�<&����u�j�w>s�(o�����+�aL����C��9�����l�ȏgg��59��}��ܢ���Ƃ;����H���C)��7�d�]�����q�}M�9����N]����\���;�ѽ>�}~�������٣�)�H��p��q}��[�f�+{���a����X�caN+L��>�g�=�e����鉆��Ш%x�<�����ș��A�
�a�|�0�3�؛�Ur(?l�����w�ȑ_<�7h��j�2�0`¼sE��d9&=	�����o����D?RG�"|��sζ�/`z��PC��փ������c�ޑ�y�z�m�ߦΒg�|&&�մo�/ǻ�z[�ʯ�=.��38 S�rt7vO���b��ﵪ(�����Fm�Ӳv#K��7	u4r	���4f���o[���33S���O]�������d-�ǫ�c���χ#M�6p>����e�2it����|��w�r��Qsc�Li|f�}���\>U<m�n���N�2���s�k���mh������_�}�ʡ��:�?ٖ%"�w�jSE�ZJ�),��̠�-��QIl�Ttz����ޒ��fʹ�־�	O7HVG�(��ֽY��z�u{ΐK�+�����/�f����OY��*�[Y���"2��1Nة���U�MlB]��w��������E+��ʜ{�DX�h+��@���ױ�㮸�_��p��:b��{M�%��;P���k�j��g=�ʣ��w���3��l
[X�$d{�M�/V����/�zkB�wW�ª�f{���������UG��V�;�]f�}@k�^��}��7��w�]�]�Hh���zL׃��Y��p�^X�Gd�v��CL���+�w�S����_GS��Ϲ���7���{�<���)8�U���z}�=��;��3+PF:K����߀W߮�u�S���O�!W�Ǻlg��|ҁ�׻:�"I���JS-���F��ۈ欲�#d	F���;�,���7��g,y�U܋�K<]o�r:��/�K��`>G����9�����/=q�Ϡ�,�\8�F�����g+�G�f`̑����Y�,�D2����Y
�߯���?;c#�JG��Fs��#�
�M��7 ���� h�v�7��j%O�Uz�Q��aω�>����U��������(��F������ɱ���pw����ϣ��O\��SB���a��
a��=��*�}ּr#ӕ���>�m�8��[�<Gu��-3AWċ�fh0uZ9���G�aFtR����M��-�S�m��E��l���5��>�8`w]�)w���@W�֜z�.,���I��RG�݌𣶛G���Ƙ��o�$�9��C���)�"�W<�ٸj��U�<ܯ_ +���vL�R{��&��QN{N���ӐT�7���r�c�j�]��7�};�HT����s�I�)T?e�5�ĳpf;q7LvzH}+L��s�=1��)|kmo���g�p�w}R=4}�5q�L�����tz�g*I�����$�����+t��Ǽq=�]��x����{i7ԇ���>۹�F����mX���7�%a�/���誏&'���(�ʵ��R���f��s�k��`
�~�9�{%DyQ�]P���kF �O����Sޯ����{�~Z��n�s�y�Zt?����`�]��NG������A�J��L���WS5y��l�A^NvIӷ�φ3q;,fN�.�=J���7ӟs�}��"5P�;6}����Y>��T��O����?�xS�'�h_�k�P�Z�q��C�gK�ɝ���!9}�ч�����^j��A�`�����Y�i�k����(ՔJF�\�=qL	���ce!�Nx�T����כ�]>Wu���a���:2�^g�/��K�Q���>0�	G�O�STɎ�ќs�3��3�d !)3P#+)�R�Xʗ�'����|��o�y�m�n(�賱7����b1'~י����z��ـS�M"�h�����R���7��'�̮�r\�[�zCZ��B��ڻ���gX���\ޢz��Q&x��vZ��~Nk�X��~���M�Gz�:��H1qaw9hݸ=qo�}�5x��f�u�=�D�?�2��a^/q��F�����~�ϸ��4<��޸���I���7y^�~�G���sD��צ�D�d�}���f��5O���M��쨲}��y5ҷƎ����y�����Ϥ� 6��a�U@3�oAai̅��IӅ� �̧p}���odl��O��V��s9ģ��x��=�r*U:(����z�&&�-YN{�A���DS�̊TW��6�{<�2��*W�Wީ���nA���(��KGo麇ל~=L��s��Z��r=$ǵ:Tn7�q쀧�n����o�~9�t<�N����.A��H#}�}b��7{yk�:jc_������I�������pݚ�5wL��=����T�D��ݓ%N���W��|G��$�˙c�	�̘w��*8�&k�ۇ�q	�_�y�K<k��-���cۉO�Mx���V,�T���ӝ�Q������c/Ӂ��WM�������`�^H<\2+���d#J����Kie.�B����[�>c=3���E��f���u�LT���� �f��"�eq���i��=��i�/i!���Vd��Ռ%�1e�8Ei�tz�`�.�� T7�X����?v.��n�ݐ�av³������ϣ=�p���i��}Q5��J'����mk�ˬoD�_��o�[ޡ,�]���֫�<Ͼ�x���=��ǁ>�����PV�^C^P��,�㟡���W��vwr��t��a���F�U�������$g�>Ӫ-֎����;}����	H����*}FZ�2.��������_�*��5�+�/&w���p�t�xc����w��8�=���*�z�ތw�.v��C��'O�/}
D��,%7��0&���%��?����=>£}-��f&F��}f<үm�X:���z%Z�ɖw����<zn�i��7)��hJ=M�dx��Ynz�_f߸.z���p�����2��O�߆ڔ}���@��_Ar�7�Ǚ�A�~ZU�j���}-º��w�؛���c�)�_�N���n����K
Θ0�J�����>���/��h�y�<�=<�{�W�hM����c_�3�ȃ��Vz���ӛ�ρc_�fF�Ddx���T��{���S&+T�9�*�I�GFK�f����	��<�_�H��	 BI��!$�X@����$��	 BI��IO��$I?�IFI$��@��� IO��$I?�	 BI�@����$�$�	'��$I?�@�����$���!$� IO�H�}H���
�2����0����������>������ǧ���UJ@I ��UB�BJ�		D}L�*��ҤR�TB+fU+m)	�%P�Z֔QM���<Ʃ5UF�B�b
	$$��� $E*��({p�R��+6����`b(Z��f�����T��B��T�	�.ƅ 4 ���
A�  ��T�B�hc6 ���q���QB�m��A�ۡ��.�q�4�#lB�*D����������MU۹�u��K��iٔ*�����J���p��G(;1�#��֛��a�wp��s*����A�wn�ә��;� �D�B�vp���t����*BWf�v�4��Wv����KmG]l�������P-iQt�ā����8�R)]wiӻ�*l2�P���U6��Q��Y"P��m�AT[H	�!J�T�nI+�mI)[l��R��&��ٶ�M�U�ZQJR6p�U�H6� T���Z*�+[f���@��
�   ���)J�����d`� CA��S�0�����      ����&MOS��S	�h���T� JR�~�� �SMF@ai���O�56���~�d���4�CLL� ���	*�F�� � ����[{<�|q�g�{5ƹp��R$[_Ť��ED^G�ajSz��G�*E�7���٬x�"���+m����������H�����T'PUT��E�L����7��x�N#(䲖b7e$�S�������`����?���_�_�����m��m��a��m��m��i��i��m�[~�o�M�*o�F��o�o���V�R�����J���UV�*���*��U�F�o���o��o���Uo��A�ClT7�I�Bo����o�&�$o�Y�o��|)�Jm� �6�i��m�m��m��m��i��m��m�m��i��m�m��i��m�m��i��m��a��m��m��9�����?g�T�O�}���-:a��[^�Ve�����Ǜy����|K����U����gh�xJ8�hmm���W4Y�c.cȠ*-�h֌Kfv"#td�T�ZtZ�fj7�m�͠�r�׉*��	V�D�.��lc�E�1P�l�5���`��U�r����B�����P��dD�����o+��� �6^a�H�GN���[�e��Zj�D�:Y[�.�VR�0�S5�F��D��{2�D�؛����X]�<���ۣ.��1 0}6c����%fm�7�#X%�,���Z���v��2��5N��y)��4�z43��0���U��
̄�݅l�f�#{�#�4��R�Q��� XT7��Q�2�dʆ}fh1!����m�墬�l[ʊG��ypS���k�^���2���&�JX��A�v�,��24��m�/��1�9v�Z�7ql�fJ�s$�*UY{2)D=�(�>��ZV`�-�AJ�&*ٛ	����;�I$������D
K@y%���:v���+6PM��Yj��PB�W�Å*	F�&�ˣh�R��f��"��m�8�L�]��'u�C[L�9�c�5k�5t�y㴎cvNpt>V��	�N#{2T7���vHZ�vj�!�f��M���r����ԡi
+.�Ķ�bBŖ	5Q]�/F^���Mإ7B��
Җ�m��*�2�0�]i2��v�^�L��	���$ e��b�1tlC�*��,޴�gUL���ݴ0��m� �H�c�ϐzĔ�;W�>Q�B���g^��Rw@�f�d�Y�ʲ�Y/��q�J�r�t�fA/w(��:5�3����v�m�'��ӵ
���V�٥���A.�]9�)iBb�̕���=un6\���(ᗌ+C�/%ԌZeK#�	^��X��ݽyWx �m*d����^ޝ�x`��M�n��=���[�7*�J��R�=��G�+Ԇmbʅ�Tl�X5 Y�oq����v��?��1r� �ij���k�Fh[D��Y26wTe:T^�N�F�Y[��kf�i�5Do�N��NC�+ۏQ���r��YB3lÚwY�X0²`,mY:52� UV�un�@��t��l0��C�`�&�%�-G�=l3\�J'�i��ѥ��A��Y "�_�\c���C�Z�����i�� ���v�+��B^PΪ�L�b��0b��)n�VȮ͡��'0�ޭ�]ռ��1Z��4`��A������o3
`ӛ%D����k,3�Җj+n���h����xDke�杄�����0�6򅐫��R���΍��VJ��ƪ8P��Oh�PÛ���VLi��h��kj;�4I����k�{4�Q��_3T�"P��T,[ܬ�&���VǿLub�"�Yׁ����c&ldKM�j���9�!��e♗Q��Q�Ɩ�܄R�@�2�V Ũ��)֊=�WbۭC5��@EZ��Oܩ#s�d:�6lGbSݸ�c�/7Q
��d�����n����ө��&�R��Oc8{����R��U"�'!b������Z�VU@��B�0̘슼t�z45���WzK�+�-���X�o>�%��]=v��[9�lva#d7�֖�1��1w��Rј��
1nCj0e�Bղc�ѭ[w��S��Z�.K�v�E��mXٖ�)N�4nɺ>sh�0YKA����A��a���f��-h6�	���x�02[9W��WP;0�� �ucm2/����`��m�D^��h�#t�n��E�Z�;����7VcKv�m���*�UE��&�7�Z��Ϭ�E��2���J����激�VU\�ʖط��\)+�g�E�l�s�/^d���f��F�-�ՙ���y�ҙ]m���1�JeU�-k���e����(�dD� �m�ub���u�Q��V�ybSv��&�Xp�beך���Њ�Xݴ�7�^
�zo2�L�0��X����T���NJ�U]�vCϭ�-�7��g�u<�㽪�(
ikl���H]Z)�O7�L��ģ�W��3��L�Vr�CV���!�0�{�ER�c�-�MSj�ͻ�)J¦�Ķ��6V��T��rE��$����
�����g-�mf�F�f�edڔɶ*݋J�w26@I�8򕏪V��y��4�Zm��&�@A[�d���%[�)�FbFj�&i+2B��xHV �m��I�r��ݗW-�"�8L���J(�It��X�[��/+�P,�U�^Q/B�՗�ʹyu6��+j8�c�#(�-l[�Ŭ�`��"är
���{��Nئ�`�W�tC0��u���ۼv�֜��N�F�)�����e4k��6j��[�	�N�t-�*�8���۹��+nT8H��h��-�i7t0e�B-к�m�L7{��E�z"��`���fY۳`�-�45�PE!�8�ј��Zj&��Sj��1Y*ˎ�T�=T�Wd�@��%�*�lr�6�7r�Cm�Wj
V�����z�E!���61��q2L[Hd+v�W�5`	9��e�qY�v��+@�9HN�V�;V(k�%fh����<�Ub��όA`�FV�c	���F�2.�6!;�r�fV:y��ߨ	Ku�j��y-��&Cm�wLu�2
9IF��;a�-�H��`����VFC�V]��I�^3��k�9����� �hk̥)�݈]C!E��US޺�6Wʅ�6�m��U/���)�F�N�R-J�����ho.���rCX��Uԙ:�7�tX.2g�H�θk1��m�,#�dPZL��2�%���I#_���6�A��r#�T;B]*�C�?���/b�����Q�h�˧�W*T��+�9,5'j�;�"�A�гVྚ��S��{�r�Ż/@�.`��J�A�;�lc�����q���&��Yv�N���G{9S-�����R����~��_��X#��duq�i�c�5�V���C7w�	��õú ��
�j�Q��í	[t�|(���Z�h� X��K4r^�h��}*��<�X�7P`/v���o[��&��V�x^"\��{��1�n��������믻Z�����7�;fd���b�9��K���Sѯ�wՓ�'�Q�z�,�b��5;�wI�#.��ȍ���%[�5ʶ�A:=�X�BUL�b��\`�"w��e�A���N���dCF��:���!MU���s��Gxv쥃ƐOE���=�&<�=v�ంä���3��r��F ���Ec��șw٧�o�ҟoU��):��w��+��Wb����X�+j��m�����M��N�R��J��_ƩN�m`}+ZUKͳ�}|��܉K�$��1��;Y(�N|*NO.�f�՘�u�tnc�,c�%�ov-Y�ʁ�D��r\�Õ�X.�Mv�k�j�B����Ş�`��+�h��Mr�d�ڡW�fz��y�'^
*T�Zu�(o:I�3Dz.�g��E��]BqT2Jy�#�r�{�e���US6я�W
�;z�U�� �}�[O��3��J�.6�<�K�Ȃ?���M���;Q���TOM�������r��M
���l�Wl+���;z���q���+���b�7�;�Z�0�w*�2�;�D�]��%Z��v�.%�j��1����J�jpW���!��6uٻÎ�״�M�'	"Ռz���=K��j��ޝV� '23���)֧E{�����F��9]���t{�)k��V�a�v���I�kQ�=�H�hV>�o��`���Ԝ����)���vl�&<̶DNE#��N-��#.�����r�Fݚy��f���y��Ӯ�N�ѻ�z�Y]`�.ws���މ��P��.�JԹج畒Q� !]m�z�����Z���Z�/��×,�=�'gY�#T�oI�ʃ�ܹp�'����t�i��茣�IH�;xdtl:��;_o�;*Gq}Q�;9�;��ʫ�x,gX�����VIڌ&�h@U�5ݨN%\BY����k[�Pw@���d�����Ũ[��p�F����o��-���-k�쨊w�#�]�y�wq��g�9���ᵥ��X8*}��� �+.4�Y�<�9S��wHCxÕ�_Υr�ï�7��Qژo�,���eK�92u�4��I�㏯ ��j�-���V��$jy��LL��w�r���C����ٍ����uXʐ���i�μx/q��Ҫ�v��Y<�RsW��F��qR�ɵe��� ,t�bUmK���Z�DVZ�yNM�w`W���m��H,*[�9ݝ��yw��R¼�[3{�ù�,�x~E��w�7�e8���I0�<��s����]�Ѥ��J�케^o��H�Q�E���:Z��:�%t��nK��T�YB����?�&�%R�n�yۦ/����llhQ����������bzc:�(������o��,�����VBt��'.���;a{r��X��G��B��Ó�����|L�_u�Ȍ���oJ��s�TM��;ΰi�S��X$W�ݗ����KN��Dz���qB�k{�!G[CU�L�9��*�;��}&���v�X͇y�r�e��J)7f�Gn1��m�]��؇!�(��:��5��Qrf	g����LB��Iv�LX;uK�Ds�}���4զ	R����4����vNj�mu�)S�`�o��^
d�Ca���7m�����Ee�����gJ��p�-]q{�nVP�(�����OL���3��
ͮ�X��ûЧ�cl.$�1K�u㑾�M���+(���	�H^��S�Jvh�ZVܬ��6��%���2o�].�c4C(���@��{�N����s�ҝe	)����V�Q��'0v2�r�x+k ]�w�ÝѴ�mE's'zy�
Dl�3�@�棊�29fc�	�p㣻�&p�����[7�X�Yyv �ܪI�*^�I2P�ۚp�2�����rf��7j)���udXoxٝ����>b�W��n�s�4T�z�Ma�	��o.�h�#�4��/��[`&�x�H	6*3Q\=q}�I���3.��;r�W;*��oG���1�`÷�,�� xv�B3���W]!���X5��0LU*Eأ�˻�y�]��{"�n��q؞��#��"���FWd�.�����ҹ�̔�����§ϫT�_w��C��v��@Ic쾂�Ft�#6x�y{�.@�z@�u��t^U����:\·�-��7GKr�J]l�Ew7ݭ �N�j�P"r�;]����xZj�N�ϟX��M�v��q�L�����k��̐��P܊�|i�o�u��Jq��4�NYpt�v�;:�1U��]�L���S%A�n9�wyN�;l�;�6��ݵw*�bTV��q7܏�y٫�:�$1����gd��E��x"���Ҳ�G����\�W��k�Y���=�9>�4�Í�
@�+'wD0F��bc%��{�"��I���$��Y���ܨ�:r�a�꒻{��c�)[�q^𠕇��Eɪ�TgF�T\>�ܫ=�����m���j�2�;3�
�<�h���FY�պ���JЇzV�����R�������_��������H�O������N������6��>^�]z)vq�����U{��ûY���[Ҁ�Z(:`��	�:"��Q��9�{
��B�,��	wXɝ٠ʊنU�X�X����H��˱[j�Ql�U�]/��Y���v6A��|��˭��c�\����q�ה'��Y�u��!�O��9|�Jڰ�b�}ɺ3^���T�9\d{cD0��lp�]73v���5�n�T�Vժ�Ä�C-Y�77�7�d��r��:GU�]�Z�ZZ��KWzX�$�ʖ;G
mn"�)G;r^��-����7K� \f��]ʳ	v�՚��"��b�/Uo*7�=�
��$�H%)]RI+I$�$�$�䒴�K�)��oEX΋��-�X��bOf�t���q�W[Çq:����{V5)+v]F�Y��dR;���QvD�8��+5ú�W�_�١�u�T���pn�Z�86�&���W�}�oZ˅��*4
��xAں8�[��.��piw6��Z5��x��S�cz��]�9T2��|Ȃɬ.�eN�#�~�'5�{��۸Bm�h�v��s�[���I�K{��w�������Z���7&m�s��lԜ"��=�6�.���|{�%i�|��$�i$�$����̴�IrJ�I%�+I$�$�#3�~����]�F.�m\vc�1\숺�5�=�j��������ҷ�U�䫈���f��ʮ�mM�R�gVީ�Ud����O�ѭ͛�u��R�Zr�t��!�Uл$��3�Q$JM�]�"@�c*��N��5�f��/[�e���ۏST��lP��m&9�6nt��L�q\uܭh�A�~��U	z�Z��Y:8����fv�u�tva�ֵ��,�S�yJ��V�'/P�o K���hY�Ҫsq�S���q9b��IWGq�p�v�h�.�}�$�%i%wk%$�I)$�H�I$������-2㭘���Y�FdaL����[+�ЫMv�5E�
�Eu�b!�BNuj���n0�̮{ʂ��<��a߰�Z{~닲Eԗ�8�^(��X\�d�-EV�1<`X7����b��Rru8�wm�ᕋ������2vP+���Gx~�eR1�y�
YDYg��7	�HC�|-���U���Fl��L�ˤ�;�-4Ψ �y�͙|����$onV��ЭT���V�ő�q(�ou��)ī���L`�E�H:�(�I$�IBI]ݥ)$�E)I$�)JI$�Hc���%��Џ'a6�����/��F�Ur+uc
�r�0��pgQ�c+���f�z`|n5��d�9gr�q��xV<"��+rЬH��s�H�r�4�7�!Oe���F��*��٫4�w?�5A���z�ّJ��DEf�^J���0�]�ɏXj(�fCf4;��Y�������b�34��Od+"�	.���9*ǫ&����xXBT�W#k�f�i���&���'*�h�<�upZ�K�wQ��r�ɺK�n)v(���G����sI�SZ!�õ���%�愻����Zѹ�YZ�L���-	Xك6��Yysz�$��TbPrm��z���̀�FG����a�k@��F$����Ŭ��̤g)��qR�A�7�M��C�P�2�:H:F�Fԡi�T%)U�w�Ow�[F����W���ű�Ե�y,X��>�a��dPiˎ��y.�$�<q�5Z��5ҔM�E�ˬ��}+Xq�N���WȳywY�4��n:X��V�aQ	F	Eۧ]	���	�.�m�i�9���pfHf7�or!�Z�p��<�N�*�;\��u��t6݉#H�%m^�3|�qY�}yb��^�.��b7�&��f��#�ܡD��NB�QNuL,M�/kn�ܼ�˾8E�E,�Es���Ó�cVa�eŒ 0G}�pv.l�ds�{�u �Իd�n�.�I�hԫ��*���7W���r�B���º�S>���淚��U����]LbM�&<:�R�ck]��'dϬ��lJO�U�P�r�g7� j�nY��/r��BمR;�O8�̘u��v�<�֏b�V��وt�|w�Ѝ�[|�;ڕ٦�<�Y4���Q��sC�����G ��Z��ˤ}�/NJ�󋔋�K�ǍU�$�N;)�8�t��2�`Uf�[��u�N�ŉ�lXsF��*��G8I�4K����9�;Ѷa�0�I��#jr�\�v��E�b�ɹ7���c�)�q�*Z�	���W'���3!������{�J�f!sW��j��W�B弾��P����c���[u�Q�rk��.��h���by�gX* ���τݬ�q���k0��'@z�i�ԋwe���Ã�.wJ�S"�@ʈdxkS��;� �İ'�ɩyX.�.f�F�1{�Ѵy�:��B�����t��ss/��ª������ �v�o� ms�dl�����'����WE|��u5��Sq`����.��hV2����5�7d�#6����V��<8s#�ov0�����'
L��uB��6��Y˧WB�U���~aUE%N�T ���j؜)��h��y�0ѥl���զ�T�U�:��+���fhAqg[v|��C��������]�������w*uѾV7����%nP��2@i N7Ip2���[JS�,轇+�N:B��`�_To��
-ŷv�Rjk�9��[��'p��x�w���]�̑لܽ�n:�{&Ke�H��X����C���F�G��!�4�E��.�����I��n̔�K��y9O{F5�F�O,b}�2��vf]�5��x�>{��!�a"�i�viT'���vtr�M�Nr���4���ok�xJ�YN�D5��������'y���r�]uqқbv;��NA.�n�FgQg�ҽE",��������~+N�'�n�ұ=���������f��vHj{���������	#$~�#�9�z�V�	��^=�t�חxgY\����b#8VrfU���|��H��Ɗˌ��G.=�L/z���muU���<9��C���m�g����jɮ�<����̢)���_;l�sE��TnF�u:B�ՙ�6��50b vޞ@�n	|8IodYB��/�{݇��ϕxH]�fǤ�q�˪�W�v�ې�ɲ��t�@�	�V�o���J����(H[.��@>z�)L�)����ӱ�H��,�v�v�.^
�d\L��#��]c�Ւ�Q8��5ڈ�}�ʎV�no$�Bܾ�Ib�.H�	%�ܻy�or=�9������gY�%1-����b�WM�4������bTSLZ�U�k�騎���QiӋ�Ƶ�lf�Q$��R�Kqa���nF��"&�-��H�-����M�UQM$D�#���!i*H4�*R!lRI�E�Ci[[��#.��nJ�c$.Ԩ�ZH ��$$$Ym��^.�EF�-�A$��D!��/�=�<�mN�.�%b��=�G�%�WCnm��+��5�$]F�Z��D�B���C>:v�E��j�;Q�Cݞ5�<���դ��4X�,n�ob%�SK>E:������~��t~�<\lW��r&"����{g(�^�΁x ����e�2MY��·0��,gE!;�.�A��Ll�˃Éb�|��)�R��W����>�UX�$�_����
&o��_�4{�"�d�����=|�~yf����J0�[V_��R�v����6)����C���3�Bb0�\��+ $�J�
쬪_g�P�����T����F��ڷx��U��dԹ��
w}����UwJ
5��o��z+<�ݫc��d�l7&4<u}�F�gZȎ�x����w���/���.ͱW��`��n����dք��P3��=qQY��k��;��xjAq�´��8���C�2�VU6z��о�5 ��y��f-���\��E���.��/�c�3��mI�x��+�gw������O��pu�VØ�s��TF]Y��ik�6�y��H=b�@����{����P�O���g������]��j��	�|w�t8���Z4]S�ױ�u�+��C�"���y�98k��`:�=�q5!�M�K�/o�kh�,+Ħ�����U��`���!a�F�pP�CϨ+
�u�o�۰�;�t��n��Fmg�k@�����,�����3m����"õE9u�ww��:=��r�;�We�ovl���L���"��@t��8U��Ѱ#
��{O���%4R����"9Ѻ1�eoջޱ�[:+��b#V�mf�
]K�G)̥�9гDe4ٚ(��h�s7� ��W�4Ӯ�z����kv6�r9��
�'� .ߌ����T^5���b�±���ѾQ{����f

�^{�����;$��ɝ+�J�������eI4�(3�;8�q�9� �E���q���wu�[>�.H̛���9[�.R�4a�[:p{Nqbjmv5��R�~ŗ�}�
E��93� ������(y7e�Xcc��x@���qއ�O����a�,��a5��I�Uݣ���Yyq�G>�su��5��o>r��:5�9ȣd'R:��݆�7�'�o7�-���onq�~a)�S:ŁH�nZ�Ćc�˭.]`��ߕ=W�k�ׯ$6r��d[#k:��'(�{�
��H�JV��s_p�ݱ���dT��Y��:�R�IJ@��Sr��������W{�I�7�@��ǿCD��}ҕ*�{}�.fo�s*�*�s7G�&��hX7_|�����d�]|K�������Ԕ�0�� ���E�P���p�^���Gk�W�̭޲0o26��_Z�IS��y`un8�D\t7h�kk��wr��
Tm���]*���v(���3�;�vM�GQ%��,�	��A�'�,v3���m�e���V���C�����g��4�p��K�$但y�F�ս�g ������4�NljZ:��Yz��:^���H�H �k%��bQF��L�[��n�l�N(��˲k��2#�R�wV�y���f��g�{�QWw��ќ��z�[�ʃo��	D�Zr�Y���8a��*pD����$�'��^�ׂxM���ǧp΁�ݪ��cmzϸ�f��H�{����_m=�Lj�X��%7#ȥVFS���^᧊��`����o��nK��}m�{�w�o�F�O����|d�x��坋2�嵩^�����@9�g��0�����Eܺ����9�̻�ظ�L��Gt�bf���mbUB�2�!�7�������٘�9Ga�O�*�n۴���~ʻq�0,Y.�YƑY}I�7v���:��ȭ�z����I7�5
+�R�1��$��=$gqҲ����� :�r�ճiգ��<D���縆$3U������=Q�=:�v�ˠ�=Gp>�QP9�uǏ󲫅����/������A]���/�a�����a�5���� �	�s����v_L���K�wv�Nђ8C��@p���UsM�i�Q��U�.���׮l�D+����n�;��c��4����G\;FU��;������^d�;���EJI%YҹԞ�@:.OX#s�s��A����Z�e�!�)�J?�;K�F��{�x��1���t��إ��̠��ł����Z�c��T���H��((��:��ǝet��C���"�oQ7f�(_E%�y]����T˃�s�+:�c�z7V���{h��*����G.��`ӳR����j���-+�#A����w��L��n6}o��JoO[1�8$�����ۯ���m�ޙG�vS(5��u�����pދ���Q�*%q�ݫ{�5�D-j��[����Y��<0��B�������A������2�D2���i��ĳ���,�a�4W�R�a��T�{���}{��Ķ�;�t�ΰAy�ɡª;�He��������P�J�����n[BV�X\��o6(�LM��qA�*�-ְ��ra�Qum�\ �]Et�?`�/ALݒ���y�q=����ȷ�j�ÎA�F�K���ێq��m�
�9�m]��FjX�+t���z?��?}c�MњwKW�H�m:� �V3R�4̥`��nb0n��hGsVI�>�l�U��k	W1"K`��LBU*�3-�-�
�U)F�j��hYe�2�B�B�Lˬ�P#�C�6Ik(��g�p�b7E�u)�-ݒl���#>֚߅:� ����F�93�E�@�1�j�:+l����CJ��,�-2I_Y��;�V��E����1]��d�aV%*˵4ĳv�# I֦�s�L���^4�kCSxp"���=Z�˧M]�4Z����F��iy)IH��20o���|B�D���$$��[���R��b�#	REF���Zֵ�ZUL�iPkW�kZ�Ԋ��#Jh�e��@A��DI4����F�nE"� �bF��	#VĹ%�rȴ�ȑZTT��k���lbҖ0č�a�!��lHf��8߽�����I��̨�fv`�D��[:�I����ٚҨy�LV��!�8G�����6�70�!<O�@����x�����c��:���I��5.v�xM-y�0r��xk�x��F���^��*=(umCڶf��[m�:�=�N��C&�<�u�u������v�C�=xE}[�Nf�9�0 ��7�k�]h�{��U_�⽨���	J���sw�<9��sk�m�$e�Q��Ɛk�xJ��/�Й���*�L-T�?U��]2zu�W��΀�$,�h�uU��ե�!�6�%}/��zb(Ž9x�7�5ʊb[q����I�Ψږ�o%}f����Ѩ7G}�I-�.g&M���=x���Mo`�C]��oᦰ�ޏ�c�zt�L�{�+�ـ�8Y�W��I���;��5a�7�cո}^�J�����sG�iGݧ��{=�Ӣn' ��T��<w�f���G�^D��+&%\2"�t����w��sN��>h+�6]��k���Jb|{�2����a��dl� %Tڞ��&b�N�RI�OL9i�v=��SI"��׳E� F��{R�C��0�ߪp�̀�/z��vwTl�SQ��<�^F�y-d�7:{�$��~���u[>���}��>�O�{2��S�{
��0�@�GH������Z;m��������w+K͛��84��?�
��2^���J��N8|���_-*8dt_?
��L/%�J^l��Ѻ^��*�%�5�N����t*���H�*���v��3F
fn��*ll`T)a�M�BL��]���o���!�1OX:7v�ă,M�O�ܛ�dp'��|���(Й;�$l`V�=�]��ٿ<hx�yR���2���#��)pb�)��"�C-z`�F��ϜI��Zn���	�g��|�s}Ŀq��u��ѣ۳UD�F~�J�TQ���Y@.}1����[�h����@��QF�N�GZ��]j�5GP:Ѯ�ʢ��F��ED�q �O�0�y�c<*����u(�VZ�iF�(�i+����*�@�T�������_9|��geV��m(>J�-mp	U�;J���wp�Ug�@Z��ʣ-Qցh6~k���vAAdy��i-~�	pC�`��s����Ǻ��9_Ꮖ,����0�D����������� ��v؎y9�r��X���7���\���-��ך:�������U���⎹W\�d����fgg=�kAƫ4j|�h�j���<c�����(:���i��U��E9
��J��ҍ!t�Bګ@���IUį k��{����+(j��ݰ��TZj�,��̭���FNXq�]�9�U��k�>ﾾ�Q�ʯ���	U��:�Zh8���Tj�ㆀ�FP�iƶ�-a
����z�=�>ϊ:�Z+MP{=����8j��LB��]k�UP-Um�5G9
4u+�A�s���3�{]<�^J�A��>J�-WەTC�>@�Te%�@+.ҨǥQģL����8ﹳ�U�֏@2�U�ƂУ[��,��3���v�N2u�i���wZ�s~ƻ�6���U�>j��j� q�����E(�T�Q�(�A�a[h�����,w�k��ZPm�%Q�J>J8��TZJ��W�eUh���*�%m����뽩/o��1���#�tJ�,V��U��XБ�7��>hXĒ�\Jr�:����	8��7�c荘�?}~3�j�y�8�_WҋJܣ�]h8��Ch�����Ѵs޿�s�޹U����2��3��|�4F�Uh�AփmQ�+��@��V�;�o޷���z'׿�G;
(�Q
�TOJ�����P�ƃ�|��,�5Ui����!]j�7�s�(2�5֪��i+�Ua��:����m��Ҳ�Q���U)^M5T>��c����MR�A@�Tu�:�Ԣ�'�Em�����Q�+MT@-���4�w��a��~�Tm;�T
{v��+�J��R�#EW 5FR��ij�Ks�:o�L��=�ڣ�(�i������ZP_ y
,�0��Um*��M��U��>j���*���-J�=J� �Tu(SHQ��A��>��WZ+�B��UiA��>������t>h�(���F�4�]@����KA�B��抮���T5T{Y���]C�3�^5�uTe��Q֫)mUJ�U�6�D�F���m �0��GǥQ�+iTY~��0N��ēy�x'��̻%h�)h@�Z�\�vNE��.�up�J%�"�)�W#
����6��"QN!өv�-Á�EL}�s��'WL5����nK�#VUY@��K@J�+�6�4g�Q��˖��+�+�Q���h�*�mHU�Ĭ�U�ң�y�5���9�w�@�Q�Ҫ�p����i��������4x̪%m��ڥ��P:��`��5�w\���*��T{��W�g�UD�l>Cǻ��!6�k{�/�:o�r���n�22�n�6\ت�<���ML�r�ΐ5���t���p��fEI�|�c:!7�z7YB��ɜt��Er�l1��� Oz߷�_&E� �����x��[+*:f�ٮ�[�@a�\Wj�;3mj�C��ޥ��������I�6ȱ{��_ QI8��ۧKѾ��
 P��JԌ�՛�P>�������}�ٞ�0�}�b�"�W�0�&�ݜb���g=���7�Ju����y}��u/Ӷ!x�@�X�����J��Ϝ�wt�t�5��}�{٥慚�Ѫ#��8���"牰���WYR��W�O/;[G-T9
gY��E�����L&��ը�}詭*f������>1��9��b+/�}]`�i �jF�ɛ�!)v��L��=ĕ�m6ȗ����9����+o!G�O�H��K��E�
&^�9d��'�'� �3
,L�o��r��e�}�Ǟ^��9$�͐���AR�T|�;�h�z�W��\b���y+{{�<|�Aׂ�x
�ک�Ӊu��W�L\�ncz��N�:�Q���x���,<�.0u+�}����
;DFSx��xA�R��Vj��l���a�&Xʋ��ͳ�=��a�y�v{�����J�E[�M��;�Ea ��N!ն�o�z����5}�޲�+ż�����͎�δ���S��������l,�;�r'�˓9̜�|�tv�m@����:��:O6�",aD����/[@^-�V)h�wPM���Xlp�9��<5ú���Y)"��&}u�I��/ʣ����@�Oԡ��'�O������i��A% <���?�}�DUD��i�n�~��%e�DH�n�M�DL8Gt��.R�J�7���#�ot��q�*�2���A��7�#[_t~�����5
5���4����]ܘ���jz��G)��oQGv��X�]s���R#d�6���u.��-�_�;��Br���+q�g���.��nvIS3��(�B�K��6��D�R�)A�J�ݤ�|��+���aMg;w�I����:���0- 9�Ҽԯ��V�M#�����V釯0�&:6�X ���Ù;D��ɕ�J� )�7��D�hOS�2�8��9�>:�1��8�$Qr4�2I�(������ݾE56š�R۶�R̲�΂�A�/-�T�̂7�fa7k,`U*�M��U^2����	D�)ǅ"[D�eL�s*�V��r�F��t*�Սo0Z˗����'j���ST�
���L�:�-���A�Q�1ti�wPd*O�5u,Ҋ�0�W1�̘��.���u�%5022��wZ-P$����j�@����a����f"s�&S�U��̌ս�#N�N�e����Z��̽�h���a&ƶ���� ]�t�6��Α����^�}��[ι���-��������u�8q>����E�LbD[m2�4�e���kT֙$U1�T�V��Ie�kzֳ�"j�]2��H���n\�gUv�"R��Ͳ�q��H�i�I��wU�$DQ��qA���4��)i)Q�F1�QwmP�DQ��%0�#q��$"	l�[��#Crі]-��!$8n�d���Y �D�V�4w�T��t�%�yd�>ӫQ:�t�Z��',�Sbx�^���67�	��7�א+�ώ�i�)��k� +��~�_��E�`���sF߾�����as�>��h{�f�4{��O�P�"��]�6�?_TC����L����ym8�.�S�>���]Tb��T�>�j/��o�Bu�E�u�,5�=KŪį�~��ʺ䞯Ӎ{C�������'|P�j7�q~�*����Vms,GwA�$�V��(��^�ә֧���N���Q���)T��$�?��ǣ��}��tonml����F�Ԯ�?��P�Yg墼��^p7���"��T#����ۮ�h����e� �����jw1(�,Ί0�I��nߩ��C����⧨nGhr+p���w�q9�oC�	�qu\��3l�nΧ�5�KVU_2ИPxnl��G	*9j�)��bs��σ!4�R�������x���r�褘Q9fM@�:����x�}7d���Z�S<�,�[�7:0v�1�D��阙����~�ɨ�O��3 Z�u����NFVUW�%vW��"O׵/u�^=p���O؉������0�y�^�)ɝ*�F������m�Tjr;\'��+ck�ԀP.4��3j+�\��a��Dިt��ϠǺ��g�5f09�E)�������$�<a�ݝ��xn�É�֌��&��I�����Ҍ��G�.;�d�5j2�ϝL��N)0���g�nM2l8�����4$-gV�&�M.5
+ �J���bbf>�=�~���_^�?��i�z�^/Rlo/2yV	��Wy��E{��6R啇�F�13\Ʋ�U��$���#f����y�6�r֒�N��x�X�l�"�M�K����G�wm����c����������G������ڠ�z���x����ZAvU]u&���%	lXG��;����	Zޙoo4�p���}b����� ��<Y��Ůjt�Ds�nuF�\�֪�D�
윑E_HE�}�~���&c阏����~������fTXe��&��u����X�WL#ϲ{&�ȎDꉂ�r�~���)F���g����� Mdc��T5w�E�,j�'��Y����1�]*[3/�c�G�7�aR�f�˳~��V�:�azϥv��
�wжŁj��=��/_��3]�c,��axa?��~z�EI=�.�wC[����Y*�V��Q���ݨ�J��4�G*I2
�f�!�mŀ����n;λ��[�;�w�G�Z����#�������'�/�~h���9�:�f��p��q;�Q�,v���b�%	�B��]Gs�cY��U�!���셶�r����Ł���?vj����{�m��5���Zu���s2����Ǫ��q��e�b�W`��C�Fx�.��nod�GK��u<3�|y]^�8��B�)ϋ�x��,�/a�#[�Xb�r�,ִ����ͥx���9{[b�������pw\n�dr#gU�#�G4�����[�{����R�)UU��>%��?W��k��֚?��R��M�����v��yA�w�߾3Y	pū͊o����>q�H�]��r���uA&ַ���'��4U��
yϩWe��'�nn�JK;�E	�;�ӌK����R �:�=N�i����y�g��e9k��提�;�:���50�����R�@�w�㢬_�#o�:q6�i��F�9�Ԩо��2��0�۹�s�r�~ѭJsN��ut|5M*c[qkūB�����?
R�@Z��/�}���u�������{��r�
]ǈ0{6t��W3}�^�N�B��f��ժ��Wp�ZBr�5�}�M�~�{�;�v�>vo��l���#���W,��T�9	]��s����m����GOF��w:�0f�N�/�	W݆�&7��'��1Wd}ʦ�L����F���~t{.7��$mm�oM��x,w��Zھ[<"�ʛ���ǻ�w��Y9.��Q�*��j�	�����Ո��O\�Ξɺ�m�9ar�{�r�2�5����$Lyڲ�V�ayIWg%w�wn���<\�DΗ�90��#��e�ع��Oz&Q��(�^��$+�6872E6ʠ�ws��ˉ��x�k��Ӡ����[f�E�f�;�OK�u=14�=�C��ß���9�5`^�zCww�;a7�9��Ԝ!W�<�6��i^�m��k�%� �C�Ie:C�\�e9s����U
-U)U@{�����O���u�b'N��g��8��LYxLwr�ƺ�oҜ;_V��g�C׷�ױOg�����lu��a���qm;�:yQ߶)�lFV��j>n������֍���V�7I~�Ǚ�ԇ]�>�l*�I�$��1OBTM�̜EU�7m�,u8J�]q�����P/�r��\������}�E����}9�8_�e^��t�t�?5���zIKw��5P5�U�#W���뽷��s��l�;[�
�Ks��q���Nf�ݍ�݃:6o05(��MU�S^����/���� V��iw�Nǝ}�_#���3��t�[�ۚ���;�!q&����Ok4�C�͋X���M�@����]�N������5c�uE4qn���A�	��3hӣ�rB�8[ub6��NYw'U��>m��I��W�Rtņ��온�敓X�U�Z�;�a1L�_o:�u�>!GۂAӬ+N����	P�`<���D$E`@�B�tqmn�ug4�X�i`c'e�%K��Vc��%��ْ���Җ,7��a-�-c%˭[t��Af[icn��T5;���U����XV�
6�v�ۂ`�"�i��l�U�,�EDj�Jb�ݲ��U�6�c�xS3 #��X�c y:����];C�'i�ʼH�I�M7����m��)��z�n�ĝb:�^s�e�~�'+�h���.�X��_Km�H����\ֱcR[c���d$�qx��J���ht´���iK`��H��m���kZ5%b��F�BB\.�#P�$�	5��Z5q���H.$j�ܑ�7�q1pUEF�]�R�IB�J�`�l� k[��j6b춮�H�F5(E�"HF�,DL0q*bZ��"���h�(" �EZ�.�ႍ5�	�����:���]��1f���t��	4�{6k=�_<�;�����- ��G�}��~��{�q��g@�^�a�������Y���<c�ڹY^�m�A��	{����S�"���^�WaK�NG�9�gc�T(ߑ�i��݉��S̮�z��T}<�-/Ε#�<-�:�x��[��|�����7�
��OQ�X�M���z���l�_���RW˰�w}�%"x�B�Ȯ[�G��q�W����]Fx�-{l�U��1����a[U�]��[�Ǻ��A�Y\(��Q�:w L��H�+��U��j�j�@��w�����Ƈ��N��X����P��5�A��KE���P&��-ݭ�����u��}�aÜ�f��QY-ԅ|�k� ���3Z��N�W�`n��e���nZ%���锗*!��#�����p��]F��%�aJ�o��;<C��N�ӎ�ݴ;��n:�V�U�ml�B=�,��:��(q�5A%y�L<�;���S>�X�؟�_W��_[@-P�TUg�o����o����d��ι�u�������0�Zb�r�	����s�K�lG�mr� �
�@�λ�=��%�F�Rq��Rq�V;�:2����d��Pf�Ҧ*A�dYy�z3X^�]|:�.x�|�N�[4=�:{�=�b67���m7ď_�4�2��'�>��}1�F�L{�2�){��%^�Ҭ�Wh�sg��W�B�MA��-ݴU.�ǒ.0�q(����8u}�'B��D~��>���J� >�^�������f�n�5��dd��U8s�5Mч�Q��<T���G�
���?�Q#�Q����
ɖ)EY�n�)�9~^���U}fe�}Ko�7���ٍ�U�tm�Ε�d'y���z��	b�L�yvUd���b'��{7M$����Y����ďI����W��qVP%���޺���U��g�B͇�+0J�����p��ն�j
e\��)�DV�
�0O("�]�}�;����%�P�P)@Q���}��{\m��fr��_�)F�zc�I�����y ;6{��ڊ_w 9kKϞZ�tn�T4Fq�b�M�0�&C@x�R9��`i@�P��ko��ô���`���ƶ*\s�ŏ���"ͱ"μ)>�țyHq�*�sN�p'�]tn;6/g�;���Y�2Hu�q����֎B�א���S�|g�����Cv����@�H��r�-`onM���p����|���h��<t�+�+�8sX�����`�� ����Q_��Z����*���O{���O}{�k�#���_����|�����!1����V���m��9��[T@3�z{���Ć��q�� `���%�V�4���ތQ�hHa�'G;D7�F�ti�]�8������/y�:�Mm��ZV~��F���U��9+Й�n�1R��us£ �Z�u��S�e��X5�Ûv���cf�5w�҉I0�!ش3˦;Hͼ�Nt����_}U���hj�Z��7�g_s����
����k�@p����x��p\O?�uᓃַT��{�r
��T�Zw�+q�����B����o#+�����pѲ���V�\_a+ �:����#E&YG��i{P�N�{/��nv�v�?o-3�,����_v��.�]�ae@���v�=NoiJ�|'f.xw�Â���ߩ6,�g��J��u�7��㇏9��{����*ܧ�R0�д�霙�������VAh�����|bo��F��s�M�+�<�;;��p�-9��罥���iR��7�o{�;����--�@׏���?j�	o�˄����m��t�^�����E�#�(�<|~���߼��{���=�o����TP?Q~��̸緌����>N&װ˵�*��[�̭?�3�}���&l���������,�C�7+}�$@;TxS_^/���K��4���[��^W�~����,S/��(a�z�t*R�B�6�>ix�Qơw�j��kk��k.%���j�4]��aD~79��B�F��=�o�~��N��;�ۤ��`ө]ƀ���j���j��T�8˗r%�hP�g�U�M\�� ��@X�I�s��]^�Z��|�w�����P-U-U-A��������Χ	��ǚ�f�p�4sn��2�o���D?`#H�ˑ*c��\�� S�(%��'`����E%�Ӷ�	(k�C�:�ۮa߼���,��X��!�O�̌YؾSG���\Ζs�0���l�t��,�_!��D�umf�OE	�	����1�����O�r��M'a����hv���ȏ�\=����{�5D!�{X&��<Ŋ�0$MLu�f��l�=0�9�Ց������Px�s!�@�
`K���}�]jsj��ǅGy.�:_R�F�]�F}�G�.$�I^T��PQ+z+R�(�qK'x A_����-QJU-P{���wB~�~o��,�E�~���6��=�������F�{�{Uy����R��3{���!��}��#�\x�z��a������ g�Ä�Dn�j���}�]J��}���H�r�f�di��/�W�ײTI�{�?�><_�a'��v+?
�������~�8~��L���,b�N�H/"x̛�0lt~n ��̉k�
سҮD�U�z�f�DD��j�l����U�q�]�gFF,�r��9�#��������*�MwR��x��~�d1��W1�˧I���~'�{�|�Q���w^��p�7�擡R�-ԅ\��d��S�����v+Czw�G�dޫ�B�@�g"vv���|�����Vآ���종Ane� �f�y�<E�6�$>s��YW�gGlN7���w�����s"���5Q�z�w9�ht�4�M���J��kp�Ӫ�1���S�ur[�b�u��f��V-D=�ɗ�/�F���c�Nt���=�oV��D����|�A:���������_Q�{$�1�ݙh�K�.[�U��v�1;:ܝZ��C ۠�m��b6�*�j@�S���g�!��S8T&y����7������+�]�;۵R����on�H�h�!�y�1�]9Gdd�}��k��H8�F+=f�Y��7��+�"�C�c�2���v�q����YH�� �gLɣ�\��4f27x[�����x��j�h�d�8���J��y't����FNù�6.,��v�;v����jL5mC˷`��Ns1Kʅm��}�8��WM�pf�4kY�FӒ�un>���v�l�4�[��	.�����.��fqE$	I B)$��0���H2����=��o���'=r�T���xI/YƵ��Y�	W+���"V1��Z�,�F����&1e� �-��VV1��Z�ub�iE̒�	$Em�Q1&1u��69��Y�(2U2*�R1�ش���eb�%���*��LFˌ-��)p��Z[Ī��1ńKp�b-4�a!���b��TIwm�$B����qb��S��m���G��L��a}H݌�FقU�-���-B$&.���,0�@��5�Gb�|���ft�{�U�\^=���Fs�L'Yf	E=��_ 
U(P�W1���}�O�Qnę�ӿ�ș�)W��g۳�Ow��]!n_�rrͧ\��C���lӭ�܏N��{"i;�F$��>z��2�ͺ��[�N<L���rg���K�9�M���̗��"�}DZ^?>����d<F�a�e�FZ��/ˏb�����q��}��ɮ7�稤18N=G�����?bx|O�i��,�K��Dc*�1�24�cت���$>澲!����a�H�*�O�i��@C���(���Ⱦ�}�?��_�6/8��(��Ǡ�En=�����ʆ���i�-.�7c�ռe9Zc\`����\�;��A� ��E^�~�۶}yǡ9+N�&�T6�*&���]�^��?��Y
��~�_�z�gg0+,�kFv��l<��/1r��#N�7�r�MŦ�w��{zng$��&�����=�:3�
��h�1ʔ��n�`ʓ����C�m������R�l�/����3���#Ix�w��:w�������]�~����5w2�Rp�>��w���y\�/!�k�]F�j��uQ=����G��5.�8��8�aa�,��
��1�Ӆ�����~�����}�@F�_���^�y}���lV���޻Ӻ]N��Vr/�A{�HG�
Z�8��"��Ǳ؝��I��U_����*�>Î���(���m��][ˡB������i{)�}xG�-�G��r��a��Sx���wU�=����?h��653��}R�OS�T��B����>;��X�|r��h�Q8F��}�-��튩�#�ƈ�7��#96F��>���~CB�)�:ek��W��h>LurouJ�*���Y?
���3��}�T�p��l��f�>{�e�i��Nݡ=a����;E��m�p���f��t�g��"��t�p�!���"ȳ���!�z�=R�6T�T�ju�[���v�m���Mhʸ(�1h+%u:V�b8`Ѭ��3������@��Z���(�g�}��>o2�'ܹu�����i�����5�4�>� 4�Ulx���N}hh�t����ӵv4��}�,�/�l3<���	��~�e�o�t�|�2�E4�3i�L9��"@��tt	Șf�ة�aE��8��Ӟ��g]a�=�c�C𳺳�DYA��h�Ff����<2�,�c��^5�x����<�������f��!j�T}k᜾��΃_{�w����q���uj�"q��w�<E
������f,"E�"�> #���>�}~7V!9��,c� Uk�y�{k���o)�:���l}���˛�w�
�]��@;�IU7�p�G��c�B���@���>�^=꿧ɼͿ���}ƾ4V��N��5���Y���u1���4�A_�8�?2+�+ݢ�_]�Pÿ��Hy�a�"�i�~�Š����]E6x��>?JA�}���ߘgOˎ�J>����/y�mC��	�M:N?!�:��<ӗ�X��Ǝ�������,THۍ,K�Ĉ��ST����5�d�DÉ�ȧ+7z�l�r���ŚR�iv�DY����ҹ���N�1O�}������"���\:���w����S�k�G|�b��_��Pt��{�@�b�+������j�{�k��s8sd�����8�>�r�-�ۻ�7����������������}����S���p������͝�8k��[=Z;��@2�,�6t�`4F�:�iAd�_���u��b��h��.Սvkτ��:�mӄ��m���B8�;�>�����p��ş�zp��(���~��Lw\MI_�z�Lz�T&��7�a�/�٧�̰o�7�w�_0Ӹg�.ܛL�眞M���g<{�A����Z�U4F�i���i�5;��}�gs�;���^v�2��"w9�{{6�=�Gھ��|�b�D؀T�b	h^e9��1֑ն
� ,ڎ"9���b�z;�F�N�D*�w��Y�o*nx�]CW)'W�]U]�T-P�UU��:��̿���9������8��o��5�J�5�f�<f:�OfV��,�5����[/7���w������L����Ha�<E���Lf�{������V�8�~_t�^�-+ܿzXDx<p�,���x�!��&�/e�5��;p֘�8쯱����>矌��Z��I�ڂ��Bȯ&l�"����"�;��}��'��5�����N�YD��z�W�E��}�t��f�[ _-8E�1�^}&����l�����<EEgM�B՞?o��u�^�ts3^�o}w�Y|~���܂vr�D7��h^H���颺����2\�M�΢��+|����(?5E(U(���>�%�?C�{�&��K�����I}������6k��_X�w��/���W���L�\od*��H.~�./�$ZB"�l^��_u`���#��o�#�n_��_���e�[h����7��Qк���<x���Gu�������Ǿ��t�[�q2�z��R�J֘32e�XY����7G��1�ky
�2xc��8�<ׄ�7�ӍO9O<��������y�����w���cDv�p��{3����x����
�>5�|�7m@��͸8�R���Gk�k�9e��+xD���F��+�;�S���x��������A���
)B�����d�����+��{5u9���Y=��0���T��7|Y�h?/��x�1B� ���**Y��+P�G�8G��Y��9k�ꐧ���h�#-}DQ�dD����իH���׋�g�~��Ӧ����52��=��b6w�H��20� �
BdK]�N
!��
!��k�v�6�����U�����tj&�p��u���\|���̇���o���h�~��hU.+�!����@���V�w;ֹ�hY��X��� ��.\�����j���F�C�U�*y�L�;"��ʃ�;F�lUl�Rh�Y��İ5ս��&�pWP�i���~hZPR����}އ皇�!��ի��JN�u�ߵ��o�S]����f�H�6²"�{KpUol��.�MZ'i�k'O������x5K����g��D:lB�C�����gN���c��*�ge��ՖG��C�V��Q��}s;w�j�A�������e�ilC_��v���V���_ZA�(���F��$���V��Ǿ�+�oAdl� �2	��J߳��ﮭ袳�x=�J_)_���w�	��'�{�!�)n}��5�c���8�f��0+���6v�����N:|���dW�YT!�.l8II��w+ |8$�Cbs��/(X���C�����I��v�Ֆ���}�݅�iY�:Nu�$�0�Lg�0����I��i[��e���Ƿ�1Yr�����R��u�s���JpJ�>J���3D^Z��MK�+���ش�J�#X6	�/t"5Gu��%vSG_mlo�.�n�e;�,�d�z/U�D2f!�G��+\�̱Y��-�N�Ìu�=f�]9.%m^c�U�F��+�k�j�:�9k7��V����VZ��٨cu@�m�ā��_v�=�w;��Y׽�w���ǽr#�V�˫�/��w��M�H�|�X]Kwi	Co��D5����w�l���̫olp<%�m�3�儸���S��x����]UH�S�Z�,�e�����}R��9~��ԑڒT�5uWWB�!]���+�
[ ����X�z����"��v�`�s�w]!�c)�:�'�RZѤX���j���ӎ��F�ܶ�N�O�f����7����Ӑ�ݪ�|n�4+(ѽ�(��\\��֧��B�M/u�ٺ��:V:��䳓���	����)�H͜��}B�vq㌸gK�9^��)b�iI_)Z�P����-ֺa�ڬ�Ꮖ)iw���L��$SR|� �Th��i��."����gBL�`�q�`��R+�01-��ZI[ӝk:Ŗm��lH-�X����Z���IpeM^u�k2���Q��0`�ĻIS)T~i��?(�	E�q�!q$�]U��F�$_B�f�("�J��!eطU�	�)n	,��.�v�ݠ��Z"A��Z7*"LFZ�%b]F%�H�ɋ��EH4��-�*�.�Q���f5�hH�l$?8����(�A�wh\%���qd[��&1�BAp��IB�*\�P�UA�	$"*ҐVH����~u�n�~����{�K�|w:\@sy�x�ZF�!�#�133?}��s������Io�'�ʕ5fps�,����̩序K��x��Z��O��8ІΚ�^�������QþL�C�S��0� :q x�o=��������~�>����tPc�BwSY������4�G�C�N�:||w�����Mm����G�O�_��1��^b'���[gS��l���F/���fRf�>T-}�;v9�:@�����G�=LB2��%͙�ՠa�9�����-��-�5��o��o�=���0��_;ms�����cU{zkk����f�m�$*0)�B哊-�G��"5�Fo
9'��u.��2�u���a�w���w�~j��j�����>'�>�����?>� �<Q��4A$7���~_o[s�a�Χ�U��M5�n~;���w��!־�sKK�d>����!������0�Ԭ=N�R:��r��4�Μ_[λ����i<۴ҤO�}9��>ބ���a�C,�8A?��[�GM�a��W����e���!<9�x����!}t�á����t�X@����kF����\��*^=!��╗��ay}�!gN���y�?IyV*��K�x���j�y��g�n���;�Pv�.bf�}�ܣ
�o�+���o2��Ќќ�Z���<<�/;�WXy��=T�<܁2R���Sh�i-��������_����*����������q�.�Ȧ��_:�.���ֳ�MU�g;��^�G܏+0je�?-C!ּu�W5���|�{�o�#O$� A@DG]�����V�"lzp�i�n�rgЉ�����N��#��%Gق"�C����ƹ�;�$�G���ȡ��}e�!��ۧ�O'o/�cݜ޹�ƴ�p�6�:��۴0�z��D��+`�l`Q�,�m�yvץ��� S�v���	|�E��F]�9}����a���iF���?"_�]�7�)N�}5�R��^y�k��/��z糋�=����+�R��R�s�g���tD���MDַg�Oɝζ�"�4]~�}d�����/�?����+��dz�}|y���Jo2Ѹ`���KU�9�4s��e]:�Κb���"��c�x��a��Y��P�4�{�uF��0�!7���.O��FhZ�9g��z����=�����o>5�ʅ T�=3#6�b�D��4�ń�S�&0��"$v�/�q��Q���Vw��u��
�i9x�5�(�:����'��tcO�HY��G,j�t�Y���x�������x�g��������Ӕ��D�p�Y�}/��)	Xk�:?��q\�$_�#�1���L�-G��}��ɯ�z�Y2�C��K�J�(�g�w���I����X�/���&YD#\�����ʟK�X�������-"�$9�Q{����>B�|��\a9?N��'�tm	&Ư^<��Ҿea�@�)��E��(�g=����nd^#L:}��� O�D�����ۣԬ�L��v/C��p�hA#7���8�HV,4-������3̌!d���{{鈑��Dx��������C�cѤ�{(���N*�?~_�P$�������ތ�~�0E(�M!�9�+�P���o�vo�ks��6y���೑p���J�|c��I��_�
��U�����?��Wni�e�o\���s������{�-�i�F\4G(|D��Ĉ�gw��o���P24��
"�����g�F���;|�t�?e�����ɯU̓����ɵ�R���!5�2�}�y�zĭR韐���c�g
=�|ȣ���=ХgC�ĝ�G�?i�R��:V|l�&�8������5n�54AM�w ������w'�#da��4�äup;3|�![��&D�jW���c�]0.Xo�Q[�V�2��܏;Ρw��qV��W��v��'��|q��eΠ铺�y�]��n�`����iqu;Q��;��A�>�9�������A��_���߰����K��a��/�f�WLI����8��x��7T��~�R�AU\,N&��>?GOש��9�A8E�c�eY0n�l�@q`Ѳ/���� N�ӧ�?J��Xç�Y��A
XG������3�'�\������#�$Y��\݆f�D�for~¡mBwf&0ӔI��5�78��`I
XC��C1#5|���±U�M�e{�~g�D:�������nrFb���V�����aIDa��r�C�*�b��5�ɧg�֍ ��G*���/�zu�vn�G�iAJ�����>NrV�ن�:Lסn��o�5�y�w�s�����G�y�n��m4��}�w>���#��ȳf��'�hC����ٴ�cCd3-|͚q��G�k;��V׳���.� ���? �C5^#�� e~G�ժ�h\E��>jQO�BZ�r�v�'���`����oVB(�e4��ˤ���^']�����:l�8]�CRk"ύ�bh�����S�s������C�ӎu띕�ޥ/ι���}�5��ht�5�W���8�~v��SH}hxt�Tr�76�O�i��i�ѫ.v�IKg�xg��)8v�V�oY�/��{�y�����T>���i#_���5h����I���D���N�fW]���9LHx�ƠsP]Wyf�=9Wֶ�ȋ x� u
0��/S�S��ڼ�}�^�4/����M�,:x�T�����?����?.!Z��|����F���[�M�����ev�е�t:��C��0�D{�5D�j)i�!g뛔��nԭ4��2]P�z��+`��"�ͩKn�����M���D/���ϩ
�*~퉪�����c�:�#�M�j*��P��E`�����������oL1���f�4�o��G��3j1��it�Q8;�+�G��&b&~��������n��C\�����N�K��[�wou�Ng��oGi$=���u�[/�c�1��;�*tU�:��$�4h�G)���Nr��(E^�{t�4@��j����+�5^��9w	N�����a���/����͐yU����s2�ϴ.<G"��@\�Ҍ}U�6���y}��[���g���%'C:T��>����aBb������ <��Яo{4����w��_c��!�~(�������?V�x��X�� �q뮏:��T�f���D��-�m���.��1Q[�7r6��녛����G9Q�}g�;��.ڮ$�y����o�6�Ym�M��2��!��dc�\9v��M�Ǒj4�zf�H.�9���x�:���"4;K�ae���` �U:��Ac���KITZf�۬f`͘.�����2d�i�<(k����N7\�^��j��'�uu���ZuR�em�PwP���㝧7C�,UՄP�vs=�$S%w.���'��\��ڦr�}"!U(ƃ-�7T0�_�Y��8T,���n��`���]���e�}f���qRr0� ��d�!1ڭy�LXpR��V�I��C2�V��Nb�3y.�̸*�,�.eK��l@�����1f+��%�n�L�:�mEx.�V<@�;�)0ۉ�t��m�X��h�/�mj,�mh5p�I�y��e�+	MC����MٵV����Peˤ���-T���Or�`��I��Z��tK-�gX��@�"��]��������������E�m�Z�Z,0,RG*���k����v�<4��7l3M��"�^e�\�maJ����ea$�S"tP4/&�0���R1���w���D���VD�"Ȋ�?�H�|�(d���(��H���m�$��4F��Z�[�cZ�z�RK�ԕ�¢�	m��1t�������_6�	�B�i�~�2�l������b[t����Ȍ����l�.ۄ�!rU�8�Kb4#B�w�1b�q�L��ZKHܫ�-�m��(�c�^1�[ĩX�b]*\�*)p�h��/l�$L1�ى.�*�ZT@Je�ۖ{-�8=w���\_3ښ�S�1�Zc�|h.r�\Ớ:7>���.���q�E��-Z��[��ࢊ3��>��2���5��!��`�ej��'������c?_k]���:���
4pװg��.Rtz�g�F�<��B�lM2J2gf��wPZ��c�1��W�ɜ#�k�x�Ɔ��nL�\���I>s�Ymץ{pä�'Mg���{>�Z�C�U:�2�#�\훓�w��,vc�Sf�8�m�%2e�R�������3Y��2'��]�~��2!�y.^�L��f����0D����T&����Hd~,r��%w�0���~Bg��u
��=ʁƺ�a�������I�Mq�0
]�pU�Qe�E�k�����(/+��}w���s��j�����w1����f����1k�9�k���՜���u�:�(��� H�3ƽN��O.9�+f;�P�!��A�C�ܟ�~�9�/-j���ϯ/����g0��m:�C�GC��,��y�'�&����8�h#+�B(���p۲�g���R�V~�h]�/�c�_m �%��"�C�m�""8aЖ��5Z�*�շV0����L���+�E��!�~�/W����TE�����fr������ٝN���E�ثc��a 6e977u�:��\nAū[����5:��\�y��[�{��RеKUU��o��������GᔙP�9�9��������"4�dx�gᙗ,V�s�3�iu�!�4�'O�bDQ~�̥��_L��D��PH�?9�iD��'�����d�'�D U�@F�h�Ծ�"p�է'�w�X־�-��D7R|��D��=�7���7�=����Qq�t���h�-��_c�Q�ő�f�,{^/�~�B�ŝ+74�į'}�{f���ι�wjmX~�_�ޱ|���&v�d�I�U��2-��iӸkaj��yu�=�ya����<�tV�����b�tx^E��������_�ZD���{��i��%�H����/�����,���!���ˢ�<�Ë#H�_Ax��(r�
�6C磌����־�VY�$��[6t�!�r(��/|��,#8p�*%�	�mB5��|nr'>5�6e�N��k@?æG�������V8u#�U$D3�~�x�)����|v*a�a+�²���,�df�9��D*���,�.�`�ћ��1��t��������]4� ^ܨr���|�(���>����$��/;���Y��S�l��o�\�����έ�ܭ	3�
���;�ߚPZ(����|����{��w�j;�\`��=��o���M�~��g�ѷ�#���Y�U+yf����]�Z�B�)b��Jyǎ�f�I�h�B\��b��ӗ��6wKG��D�{��a����!���Ùs���\�1����ɧXE�#v��ْiL� ��}����|�%�AW��o��B�l��l�K�굷�'60��Ի	��gXW�/6F,�x�{��=�N�=D�ZZ�ܷH���	�bv$};�����g虈����k��|�N����ɇ$�T�)�+�<5�soga�6`�q)
��z2)����5���^P�5�E|�9�[b]�(,��s�gJrR�1��
�R�ݜ��w��$ɶ�i|L�V�f��^�`���DEnO�q�bu	p{3��ĤR��=ᔬ�$k�y�wg[�3Muqb�F�멝F8Tq�)s�E�5$�[��k&���c�S�!+�ϯ���"oIXV�@LXJ�w;޻��[�;���W���~�߭�n�]�^W����m�͎����p��o�����1[僷ѶntEJч!����)��<kƸQ�]�1\>�)��u��
>4BhP=�f�/^y>��E�h�$nttkȗ�.�g�9L��p�^&g���(���x1{�39��j��]T���̷�d�}�ЯE��	{��y���x�0r��y����@U��~�Z���}r��(��Y�-(ѡL)Y$��Q0�YۘTe,�o��y�t�w��;��~JZ�����o�����߫ ,���9J�=����u��y�'F��vd�����]}�\c_��r�Mnf�����2�ձ3����hM{xJ+�mo��µ�$�]8�dF�ɣ�Tg@��a�d-��2v�sϪj�cE���J��ٵ}	Z�L�F.�ȝ$ϳ1]P�g���ݷrA,\���y�K�f�b�`{�:.>Z��*��Q�̏r�ڶ��+�.��RJr�DP�;�]v����M�}-g��"�&^����Ey��G�
R�R�R�1x�������N�m�!	.jn�R�%D�{����:?�_��~�������H�vdJ�fU���.i/��T��e�s]�E�	���{P���jv�Erd�|zR"`smʢa�si�݊Vn5�P��=X�~2���0��(�i�����<a�yfV��ؾ˪�[k]�gl0(b��=.<B�N����4�;Sۤə�i]w1��X5����5�:�LsZ�|�o�ӷ�λ�o��W�������?�j��\:��
��#[YvXn����hq�f;1��s�eQ)�T^��k�3�+�t���w�y�Oc7�#A�Rd"��b�>�碵�a��l,�MGa��p�5�����R�~���:C@ǝ%m��g��K�u)y���&��[�_�~���F�^P0f��W黪1�~�%���_�����RBP�f�2�5�̤T�fU_겭�Ŷx0Au܂�茝-]��j&�����r
қb�YޔwE�CǶ��O�LS_meZ@�v�}��X�nt��Y7��q���V�[����C�kY�
����鶤�t�2t&ƕ{��5�^㙬@�V�3b�i�5(L�T3dB�'��胢��噘���dlh,u�\7}ۼG8g3�ӳ��[�����՛�w`E�Wab&�����u�@�
^��.���	�:�9�\FSI�ځu�-�w��-nێ�2�'>4շ��z:��{f�M�mi�F�6��%M�
ٳ�m`�5�������
��F�����S�Y�����p�fԊFE���p�?�2X�&ŋǒ�F�t��}�P� �o�i�S	&���F
��aC�͊��GUճ��z�8So0�l��ZR5�J,.�S�:N�&��A�k뢚
���ß�2�$�I�%?�cn[�+���72і��a��I�8��:/i�)�bx^�U�d5�H�B��n�BPm��
��w�����0GPS���m�b㴪�ۼ�INa̰3S,�k[Ku�eڼe�t�^� �O�2�Q4J���T�DH�&0��Lqr��]�d�ۺ�3�i�e���r˖څ�[,CX�S"��ur�M�QB�A����L�]˔����T�`�Zִfe�TP�"e[�5 ��Wuv�Espӌ8n7.�"��B���r�,G	���"�����KE�K�V�I.夶�uu��xn�$���b��E��!j]�h]%�cK��ld.Ѷ�q� ��I	&.[��nY.I�#�X�rTb(~b���Y��D���d*2`���p��2���!6�e��"�2Yh��@�N���f�L�E�� �Y���!� �e9'N���q������q��?:���^����\-"�?B��#G����wh�<VX��]��5+ͼ��ػ+f́��^�rG0�)`�TT����=�r��Ȿd�o���u��+m��,��l��)�B�wE����<�d�)S�C��||[���dq�6�@	�.xcU�t���\����EG��6o<��q|��@�*�-,��wb��S"�!��O�;*�Ufʙ����1dfb\�Ft��	*�H��&b�N�RK���_��k�����zz��Y33��pt���	a0�N
5������/;9��1˒@s7�D-�����]㭸��]�ӻ��F�
��k���m~V�w�d�}�7��Y���)���(�3l�;�[����_E��&�W`]��s��5RE��|h�b��4��H�)�w�6���ږrVy|���vIz#���%�8��:��ӟ,��>!��s3f��kZ��,�\�_P�I��+��rU�X�xt�10v�8Po�G��M	�ۗ�D�A��h��goک����K�t���kYl����jV��dsPM����yV��|+�d���a�cd/�,äW/^])��:f�=x�@��-���X�5��~�mЂ�m4�90��2'E�	�Z!?vKQ�*t�ّW1L�����Q[���[~�]�pk��Q@�U�)�C�gD[=���`�K����n%O�&�q�.���l�LODI��p�El2mA�_	������hCϋ�S}��#+f�Ɲ��Hu|����(��0�gV^|��;p�f�ݾ���gIJ�\�1�{��yƢ�c=ǈ�gz�\a��zr�MĽ�������\��"���c�:����<ؐ�mh��#"����|�����g�,�i5��ʽ������{Ƌ��zm�հm��-��<G�����Ww,p�ug):JѺ�l=���A(ԏ-Q-.I6��S��M��4�
.yԥ���۳I��b9��{�
=�$سY��]�7�r��5ev��v��ϫG�ֹ`�t����n.��v�R��ͯACF�^2l�j���coF�S�]jS<�篶���.����� {}[����z�f7�΍�0o�M&�z�U��Lf�5mv<o�eD�~Ć����'Q���s�%Ms��N)����r��;�����.��h�<��*{�%e��4�S��s��pm�ж	x�6EF3 �����������Ƚ��Fb��p�?ү{���s}w�lo���!�]�-�闑v����X���o�a�$KV�d�ͣ��(�]�zK	���;'"x0_h���P���m��k��F��o�{1]�^�ўY�U��=U���+̮��������t9b��*�[���Y�1qs|� ��#�<;�8]�i���q�Ò�nt�U(����J�v�}���z��9���u�ѿx�w��w�ն�Í5+f�Kk��"�5ܸ��dz�l�����;�;cKL�᱀<�љ�9�4��S�Z�׵]���?t�@�7i��U���'{����5j�g���V��t��R�E�U������I��͝�/s�OO�06�N�����d%]X=Uִ:��v��,��t<o�Y��l5}Ը�Zs�e��Mβy���KJ+����WwN�xR}/�[�R�&x��:�z���8�b�ؤm��$�A)ኆ2@��m�ufk���NhB� ����'�Q�jگ�%�� �H�=B胿c�I=�K�n�玮�]����x��L$��-O)+�����኱�V�ff���k�g�/j���2N���v������|��w�y{�g��ި�|��w_�m*�<��@_��A1��Z���)�����l�l2	v�4���Fm�f��5�4��f�\ksг`���r�J�,+5��6imΛ1`>��/�o��9�
-�����xpN�5�MY��������^,0���Ws��*'����3z@ў�*3.�Ÿ ތQH[��l=��/�oru�!r?U����S�p�����Ge�m�q���ʞ{���m�h�5"�Qj��Ӿ9��f�WM�Me���})tq� bc`�l�d�6_9z�έ�C��u���q u(�6��Y��9D�!�O
���u�X�݁e�����?b�fbc���kϭ8�����T�P���kt���jO��3g�ɱ�r.�l���Q�y�GU�=�ک6��+����oe"Ɍ�s ֘u]���1\��jK ���b9�a��خ¤r4���F�z
���JHJ��[;��yU:&�d�S:��]�Q�xǚ[��U���`�Ô������[fZ# �P�G�tZ�w�꠯9�g=�����Y�����ѷI>�ǥF��7 ���F�2�aVv%�����vu�E�q4ڢ2F�kڛWN��wO{YF�GB\[4�l�K��G��)W��	�9d2XBJ�vee�d�	�h=N�@�8$�<]�$�)R/OK(X�mG�x����k$T;��F��&�Q�̫��u^�8M�n��s���麜�j� ΐ����3x�̾�M����.���G��7�y�3���$V�l����3����|Ո��Q=�l��Dq�xp9VJ��ȭ��.���2B�7#���1?�Ɩ<��C���Y�:���^UY��!�C�ol4h
%h�횶����B�MB��,�m���L�5�P\H�d�x�QT���3pQ��V	}�QT�X,h4ki&��-8)Y!��^�T��wwyt$��C+2��nX��LU8vެ��V:��i����e��m4�///r;2��XOYc~�	a&S�7��X���%�q$����%�^1�y҆$uusX%��Z�vŖ�2"	L$�M���Q�գZS6�H"��K!��0���,��g�@�CQ���k��`��l3��i�E��m��-�B��w�h��Ij8ĒF������+"ˉe��ˍ�v��w�lmcW�x�%��-��T��E�H\E��t�FJĂ��qrB%�˱�jIF1�� �X�ÌH��QR6���m�ʕC��X�R#$��F�nۻ���vb칄"�%�F�������+^e?3xI�]��Ewv�Or����)	\��%	JԖ���:9z6�xRU�#Aq]�;Ҳ�/�T���n���ܤ���[Zǒ���%�z668�vG�����E�P��c*��\[��ș�u#��~Kyx���z0d�7��(�P� ��k��/׶iѭW^d�\[�y����"�|e"sO2��Rp�C|+���
��f@.5�.���c4]R�S�601[���$��}{��^�w�W��J��P=o��w:�a��[����=�>�j+5�z�{���Ӛ�P�7��&kw� 8=�5�g��0���~��:�!��L��&�9�k\�N�\����Y=����[r���y�ڵJ��sU�5��G��]	@Lg:
�t24Qa�Ѝ�vm���V�����<kΓ��/;��Vo~���lP�(�f,�;�޺�����>���Xp��D���Γ�B��s<�
���C�^L*��V�9R�N��v��E��n�v��{Ϸ�^�9m7������a%e��,�qXk�+f�� &��:�8��qx��c�t �Dɼ��KS��j�b��<W�1t���e��5����u��ݫC��({��ym�������r�5��mq�P�lF��Fh�W���B�Kmnn5�/����}�@�gS�ډ,Y��݉/�CyX��7u����$I��/X��k=a���xp���=�R����3�tq��U`�+8B%J�����K�R���z�&�66Q��Ï�F�#�T��:�z��k��Q��˝�~#4��ao6�j��	T�� �����qsR�[Q�uѝ�WY��z}�u�2|�ǈ�⡓!�ѷ��T�n��֏AZ�8;�����iq��Qb޵d�`��=,��|�r��C|��"���I~s��d���J7	u�{6��t����*���dCF�r����ffi�A�g.�k��7���Qh+%u:nQ)Z7�hVr3bx�U	����A6���D$ ��i^3��>P��]=jH_L��W^ؘ��x���#�c��z0[��PIݭ��miS�|�ɨ<o�)s鄗� ��~��!�U�c������u^\�ֵ3Wψ��IF�k,�޳Jk3Vi��f��x]$l��>Z"��'�<r�{p����]0��9ʣ�"�J�x3�2/h	�9��6�
p|,D�wqW���;��-	�����+4u�
-ox��������%�F-����>�9NUJ(N�Ԝ$��WÄ�;��K�T�gѵ:����6~oN�R�؛��vk�i��w�ڕ�B��1�������n������x
�/;*t�Y�Y��hs�{���w�}����wП9��W8PB�Jg�0��05f�u3ǚ�t��K��zM4��a�5��b ��Z��`xQ���P��S˺2�d[�i'O@nᬤzH���;�yJ���ۡ��������
:�J���fs��ޜ��p�`����>�2�n*����\�KXS���&�$�s���������F*=�6c�]e��;=����tn���R�^��ϑ��hDh����"S�����j�O����gw��H��s����{��,��@��p�{�>�w����܋�ΓH�>�V�V6�����QN�#:�/{�+���D�����Ԑ��ܢ�FMvt�v�>o��j_:�&날���Y��/#Y�#I�I&��U�Dx��4Vܵ��ޚ�j���6whJ׉b�q:d�����"x��kݓ%f\��J��-�\���a�����v5-KI�U�y��Ȯ%x���Gz�z/�U���s�e��[C	"�+���/#N��6�N��=�5hs�����Q�̞���ŬQ{X9MwR�a�gp�� ���Q����"j4�C�ё`/O����U�	�'�D���JiT�:	3���W�*�*9O_�iW���vG��=q8�1;��y��n�cKیjV�kд\�l~;���4�w��~���&��+W��ނ�+��9��xg�&�s7�&���~��г7��������|�@'n���AS�^k�@R�K�����)Y�dU4�a�a���@���q`.gU���E�s�E�I�sлQ��3���2�^�d_8��wqt=%��M��.yob��������f�]NIU����z~�ywۧ�ҠJ�L���+͙=�^i�].�;g�~�ַWY7.�k�˸ķ�\VPŜp�'�鏲��p��9����1�۫�z}_sk�uarHs¯�ft��yW�b�ဗ��ukx�W��Ye��8��E~Ot���*�mR�W�K�D"{b�mK��Ws[�+���}��U/%���h��dC�ژ�I��29�%d;�E����)�r]ؗ:$e�����:/b�a�Ju�����uu��K���FE@l�CI���mY�MA����V)'Q�sР,�"w�q�Z�K
r�yr�oTb<��-^�Y�>�����J�������Gs8юwqu�[�ɳP��.�RF�!8�y��ȫ�f�M;�sx��z�0�����h�� ���Høz�냨��V�ޗ�,��
gR���ͷ��Kn���n�`��O�ۻ������;&��2��{��#�ۡ����9:4�{�V���,��;.�E�sanV�s��L���>VL7
�ҷ���U�f����V��wFH7��|�����>�B߮J��/y��!q��m�e�D�zևW��ϴi�8��<g�78���^��lG�������\�1�z�KJFU����N���q�/�ޕ6��X��k'��z#��)�	#������<�HiD��,@��^,���;��z�Y�b9�<����8�h��hGD�	 �+*������YPq	X����!x��z�t��h��)AiF7x��6�m�H./ִ&�Ri��˰�˺f��hDQi2�35������#�e�]��P�ʲ�1���(���Qicl��$�˻-H#"�*���d&^.˄cDY&����ik%��Z[���"�(��KbLb��.ₑ��e�p�S�f��_���x>��p5ս���&.pWP�i�ӳ��I�q���P�{[� )�7�k�y�
E���iB���Z��qxZ/����I�ޑ:N7�5ʾ��1�֟aA6g��Gm���-���~ϳ�'{h���WK�X��7\qD<)P�*�<&�:p��<�D�O{a_揤�f�鱳�jm�{����'�l��5����9����>˗C���-�D�F���_�^�f��N�'�����|�cג7(?]�ݐ�F���÷u��{8�T�P�q)�����O� �7s���-X�7�A=���#�W{�o\m~,���w u�V׻!��ijM�����i\��&�(FֱS�f��o���.A��,`�Y�Z1Coa�ђ�'mn�ә�Ę.\py��ƿVc�;+:��o����eũs����<� �Ҧ�����P��C�{!����{w8�\�l��>0�/o�Qlkr�'�;���J�Nw]+��0wul1ut���HF%=�)p�^
��	\9F��k�`�ۮ����r#1�LȅYn_�U�m'���Bq��e�@Xg8��Y��)������U�vǜ,�:�j�F+ �����-L��4��v�Y�1�S�����:GP?K�sJ�w�+3�̶�y �y}�R22�F���K��,԰et�|�.�ݗU�=t�<�1��;}Ku]Y����^ɁBW[�/��+,���b�bQ1Z�R�p��PS�(���*⺱�Էk�_cF&�_D���!�����
p��H�a���Z�F��>�Ss�,�[�.O5��Dĵ�׵�l_:�znmF'3�N�K�l9H)���o<Mq��y
���*P�&��>��Rӌ,�u0t׳���}�-�]!@�R�Ȗ�7ٯ��ƒ�a/a�n�&��K�D�F�gc]�n�_b����7��{x��gi	�"�S3� Qvz�l���R�V-��cr�A�������(����ʸ��g�b`m���ٮŌ�iNb�䋂�.�OD�L�r5��O$��d��c���˘zʥ�� {ǫ�E�F�����'�oF0t�y���9�z`MB]�Vhؒ#=�]ʮ���<7��{=���΁_>4�n�g���7��sj���]������[q�>�[�-e�)��Ƽ�ud(��\����h�r.�)��v�$��%G�1oN��m�wЈt�Є�QZ��)$�.�G_��{��
�͜T����e�E��c/%_]��R�\[����]]��Z��+cq��ҏ`u�	2pC�i����]���BG=�G{:�y�,�d�X�hç1���+��ќ�+pG�?z�kdW��ّ��>Ki�w�1X��y]t�������Y��s��o��	�RY��X��y��ټ�W��@����2�J���U���Z85�A(���x���{��ZF*�Nb�Q�L��g^R{��V]z(�Z��,����q�5TS��*�GLN�n;}o(�}cI@PD�ꍭH��#�'UQw�:j���n4�k��c��k� �y���d9��;��q�Ӿ�h���@���#�Kʁ=Ԧo�#V�M#������>��o>���9SGs U��?J�ހ�/}Q�~�̳׵G[-9]ԥx�(Fo�7�.q�s6��}vE�D�(A��rͅ�(� R�;������rȈ�M�Wc�}7f��:�����,�����-�f��,]�\jb�=;o��dk��C�A(�߈&�xg��/�-����w���hh�Vfb�����_z�S��2��9F�n��tc�{=A�ro�*R��VM��?*~�$�>����gϟm�V��,�d��'��YѢ{Jݬ���kDu�je�z�{#�ξ�xg]vq�*��\�8�t��I�
|��{��e2���u�Aa��ccWX��0p١ޗ����b[2�T�:�/��¡�ۣ�/�uX̥x�y�m7��kJ�q��!��9ш_u4�	��H�]\�d������<6�@�k9UZ=��p��#�g�@�GPr�o�O�ye�y̪n�^+J�yru��ފNAW�z��4Nص��V��ΗN3Q���䦪n�°R#��V+Uک���+�q�z/M��
 �6���-�˃LRW�ӯ6�h]��&���99f�����y�Z ��S�����ݏ��Q�+����~�ie<}��`�v:��*�}�)'�'��f����|�u�썔K|�Z�R�f�3�p�E.��p���������	��{�
J����{�b�ү7�O��F����_����ѯ���S�K Q���?��O�#�ZU[�IU"-����I~�Қ]�@]�����2�~+m����l��l�s��������³�8��<%�Mb7��5�TkF�֍U*��Ԕ��UL�Ԉ�ѭ@��?��3�23ue�DAA�@DC2�(4� �"
��	H4� �5H(" �#T" �� �"�H" �"
 �"� ��#m�6F�4��wV9bk�Q���-�Zfk�C��+U�j��f��=Ym��	2!�f�1��xY�ׇ�^]yxr۟i���&���޸:���cg*���y�n�Ѻo��v��馎�l.�K9P����6m���RXY��N\m˝�]aD_ڝ���w^��׸vk?����*���uTE��Fa�c#R�{ǭ���Ļ�����y#�3�⻷�������e���|���3��>UY���t<��i�m�����d�X;�=؛�o���S��瓆'Kb����Z:�,7����ݩ���Zm��|�N7�k�g8aǋ��<O^3s�����.S�[3�~����jH^�M]�N;4��6ϳ~Lo4`���URq2��g1�V4�0 -B憖��h�V@�~!ƚ�������-����<;��8w���xSE90�	�)�)�f�0�a��7#�;��ӱ��x�������5�2�_��j�9/#��w^�<i�U���ͫ��n'�����O�[4��9~�;���P�.uheմy�~�r{��O�<���sO����s��a��Sc�ا�����ϓ���=,��K�r|��%a
Bpq`F(��BYH���E�m���b͝�_�ڰ��{�����ٌYhw��oDі�L�1E�6>
��_%������S׍Y�O&�s���[�׃&�w��rw�$�����2d��Z��եa���I"�d�j�_n��ay�gE{�;]۱�2sl�֖'�h|�t�ߗ~Kxs���L��i�.˜q�v�,3:�57\��h���>��>n�r�씈��ϳ��b�;}W��OOu���������y���O{Wx����<V��ܧ��=���C?�ߌ6g��X^�q�L�|~��%n�ͧ�������vM߽�������×��<�cg�5�H|��_ڝ�/�)j_�!��1���O�~c��{���v�Rw�El�O�}9�'>C�XaΌ���}~.7c+6V���_�sOS=���/�S�,���Gʝz�6>���fr�~��ok��l�o�fg�����)l�Ǣzӑ�}c�l�y�h��j�s82:���4�~���8�/Ws1w{4�a�S��ɧ���ގ�}�3���v��%��/�,��m}�a�}i�٢��?��=wc���yJ�������1s\9���r8��F��zڎ]6�l�F�p�O0��F��L3��/���U����.�p� <�
