BZh91AY&SY�OL9��ߔpyc����߰����  a� �               0   �@     
  @ ( 2�J������>�����  �@ �`筽ǹ�q���<z��m�u�۳�w��w�]���B��s94]���S���=�P^�Ӡ�z{��x<#ȠU��F���`IV��� �P��P�<a��װwz�=�6���n�^��{nl;�G����i���Ch1k��t�x�w�v�w� ��if���pozOg�u�����@*��c 5�U��׷K������{n���ݵ룛��S����0$<Csmf��ǥ�zf�Nٕi��-ުw��떈��ݺi��T�X�7�]r�ԯm��l���w�^qݷc�1l�J�w��ǽU��ٚ� �{��1����ۗ������=^y��c�\vt��Py�TT- U��u:�΍Ǘun�C�Z��흴��=�m��=�1˝B�#�Sgv��z��r�뎷f��R�^���f���l��(J ((      *
 ����P�`      ��f��E24124�02M0�?Ј�R�`FL 4i�ɣ L@i�R�
P �h  2i�@  	4�T�a��FF$�@�4�4�
yL&��54�@U4�b�J	��F��� !�a7��H� �
�"�21i9��9*��kPTQ�T�D$Q��i�EQ�A6���U��0���_�Ȋ�5�� ���������-LL���
��I"#�H��"�0K1ao�UQ*I'ɹQQF�
�1D� �	$�I$�>ȥA@p�g��Ɍ�x'���?5c�!;1�s��ᡫ9D3L8x()�:2;��Ώ���gWFxe0�Y�_(��1�c=�&G�YC:�x��Y�L�˴�C��T���RBGN��L��x�	���1A}(f3�GE�.�-./K'��ä�#/!)1�"_�H�W"d�Å҈��<�[<wޅY�VU%��u��1��^	�?d&?/IE�"�V0r�c+�@ڢ�p�PΥ��2P2�D�y�t�:�WW�@ɩ��Й�p���:Lc�aׄA�FH�C1�jI��$�3����(iL�Vx�F�c���'��H����(~\`�!��$��L&H�P�Be�$+?�i��i�4÷�iB$d	�� c&�N�}P1�`�x�C��e���1�=	���w�����2`vW�1� fS�$d����a1�B��L��x��(���d"�x���t��%���=p���0x�d$�K�ESzy$w�i2�2�;��������"�ID5��)�lE�L��Ba�N�ay��һt\� ��C=�H�L�2�)��#	,�%%.�Xz��1�ag�,�PLt��*'�C�q
�aY#<?	3�*=	�|c8X3S�����P�!�B��
:$Όw�L��~��,��t��=	��Gm2		q��0��/tc^���+ ~�&`�aix�ɗ�:?D(#L&Q�ǉ�2�`�!a�0e�!�1�&Tu,�C��H-.X1��	���20eVB���p��u8\�FBL��wdxcy
�<���t����5$@�_D�gF8�&x����L��p���m��:�c����8L��i�L�z���X2�爁�Y	�6�������P�c��e���1���q�.a�1���2��=*���&!��<3�>b�.�9L��c<[T6`Q�|ȫ�y�3ŝ!�#�|B#��0t�%�!2:�
�Mz�1��,��H�)2��<Ym"�a�d0�є1@�^8TY�� f'�J�ȓ�y±�^8M��~���:{�(�P�0|�C dE�2c�Td((��9\�`��c�B�xP�� c����(��n(}�,<G�.1��P�к1�fn<L�2i��xc�%�q�?&IcK�gG�t���	��Hc!+0c&����$}�Le�xr��a%*�7	��x�X�Jc��Ldk����2�j�Ɉ�@�>�&1�����w
�c��:<\d��Bc�W��1�:�GEΖ���G�g�<��Yޮ���Ь�Qe5d<�Yg�xg�?)�1���:2�(�F`�I.��H`�,�1�I��c��ɵ#�j<A#�eg�(a�+�2���a|L�KIWC<�C0���F��X��>6�Ē2G
�$c)�3�1*:0gP��O2�(�����2��8�����1�����1�3ޅ1��b�Q�xc1چx��ПWDI�cU�f>��$u1���1�׈-�1���(�	��c$d����C$g\�f1H�~Qў$s�8�9֢IጥJ%�j ��nTxg�ڎ0|mG�$gp�*$��^2#�#�(��D3G�Oon��b�g��#�$�H�^�c�3���:Q�j0d�D�:u�2�S�X�x������t��,}Ȍ)�9U	/DI�O$�GJz*Gw	���&�0���L~�L�L��/�xHc�˴�1���c3�3�Y��1��-"��P�q��SD7֨��LD���Qu��3�3�����)�t��YC�@�0�����ɔ�������\ac��1���9�A��4.1�Q���C	;�q��3�(븏�ηGH�QC�QC=)�c,c��4�P�)tp��b�`ܨ�C�(�Ǌ�m��#��_�8P�e* ���9Lci!�*ǉ�>ab��C�c�\&X�?&1��1?(�6�bR3�tc:�(cB�ZP1�;�):3�:ڈ˄8P�I�1�D3�QԠ�C!҆uڋǊKј>�C(©��5ڕ"G�1�2]�P�0�WZ��P�`�1I��.���D1�.2F�˹P�KW��'ń�2���y��GZK���ã�C<ՖI#�&ŃyQgFX�X�Q#�$�5��G�:�,d�, c,beP�1�%Zc$|�1�я�Q���X����c0��C0c;��G}#�RC1�x�ӯ���p�A'iP�k����FJL���qp�c<�tf$���`�,�0�3�2J��(g��E��藆x�.��]D@���{x�$A���1G�
�[^.�3�GK�!����"E)�mP���ȉ$�%�Fa#��'�e�#jJ p�Y$��2�*R��k��Z�$aI@�s%�Q1�t�FQ��`�Sѓ��I�,)�0����w��Ȅ��HƲ!�IP2qq�y�GeM.�dy@2<���&X��D�31��Ę�~q1�DX�X��bL��(t�:H���3�D�G�;�v�c)ʏ>1��(|~P�(��c��||]i$2!1��Ǌ�Lg��Lg��}P�;Le�׈1�P�y�Lmt���X�2�SP@��%ʆ2Ov��>Y�X�t����`�}Qc,fb��u�^(����E����mE(��(e](C,f6�t���"�}QC<>��d8���C�J򅉵$�:1�cVA�0p�c���Bc#��c;��.F:L��0e(��ʔ���C0��e��rJ-U"�NT����TY���MC�ܓ��-�T�wX��M�,$Y-�ȹ;��۳��3��H����v&��e��vf�vr����&9?�2txp����d���b�2�]�]YNc>��$�{w˹M&d�dKy)���vf�w3�ٙ�޻�-�g4�g-���})�����~��!6n���U>��9$�a�fK6H9&��6�2s�p/�r�5{�ۛ큙(ɕۄ��Ond�3w"�ၜ����8�M�6�,�f@YNl�U~W�v���;�9��)t1m��3����=�t�\�ղG���S$82_"og*ř���6~vH9�r^�X���'����r��Ou�n����w�[�v��C{2`����G����ߦ��N~�~�>�%�Ⴗ� �fL��8+��My���O@&���1�zr�����L�Ž���\/.l�{79f'T����{��-��~���p�>��\����鷐&�S����>�z�3f��ᬼ�]χ{�Y���fnL�gᄦ�w2�_3$1�O��]}���>t�?wL�4IE��E�''X.q�k^�����9�ӹ�~fs2��)0X[៲���Ϸ��ߤc�L��w������57�4���Sݞ�gF)=	yӪiv�t�S>3��7�`�{���ˇ	ᔛ�ܒ�ئW��6j�������b=v�~��|�_�ۧ�1�ә-\���7����vd�w�o9�8��{��˳��L��r����"^���];�I�ɟ�]��S�u�{{�+�'ԜΥ���*W�0w�j�xOc׷^�h��t�Mrj�m���g9�q<t�忸�}���?s��{���}�6+]�m��k��/8��L�{���sV\�����Ι7�i�϶t�e���y$��>~唐���W���r��SMY�ɱg�s�u6w;5���fI����t "o��t�s���՞���f�1SA�)=�������L�7�&Js������]�rLX�?77	+q�n�7s�����!�~�c�s}�������������a����$��䛣�n8���&6�՝霾N'w)z��vp��i�[��`���;'Jq�w�gh������d�h�u�>
���+25n�t�N�G?OC���wzm���S��&�8g7�Y���=�Ł���j�y�,����ә������Iw��t���ۄ�;w7vze���8��`x������zRP�ra��$�{��>f9��&z{��LJҪ^�a�:�{.� ���ˡ5�W#i�K ��Hu�O�'Ӳ�K'�d���7 㘹��k�29
x�V���5�N�(Y�='7�ڔ9�>ww�vw>7w���<�1��������n����������9�2�:l��Ƀ�R哑Qm4�<�ec)�7� O�t�۝�}��z�vy77�mgSs�ኹS0'��o��Yz��'���~���{!����̛E6䳞�����N,fܘg������(مI� �v}��.��1��?N�R3nN;WQ�a����4�$�g�����CM������a���I�sx39��?w�����{�����|�ܖ��5�z�](g6=�&q�9̛,�e�[��qɥ
:�y������ǐ�ݧ�	osܹ���}�&4ޘ~�g=�$�h����O�f,�/}�����~��I��7���/�&�~��p817/�&d���3a��ö���m !s7}8���y5����97o.�5�_� ������u�D��a~���~8F���K'�{�P䥆q;wGZ�eB��L��`�f=�{�����fvH��;,��;$�'/&ܗ:�U9c�3��l�F4j�~��9��8֔�ovY��Oyy���h�H���>>o3d]~��d�O;gd�9��>�E�c��Omm�Vק��(Y��YS����Ε��9����f�x�qu���sM��fy��vC{w�\���|�s�!�����;��G��,rk�/kݕ��d|���py�:1��̜~�Κ��4t��ܗ'0yj�aa�i�{{���o�'��M�7eV��!p�M7��O�O둹2wNf\�9��/ӿY�r��ώX��p�1����� �l�g�GN����#X��-�y3f�3���d��s��9~��n,��%�n���gg4	�5n���rC�s�.��N�!�#�zt|�=�7=�����M�4��Lg�Nr�*\8w����c�&v��N%�>!���K�gϒs�7g,_��>0���A��i��0�q�o��� ��F��nl�w��a�l)v�?��糒r].[3�ήhm���ɳ1z߽��8~3i�3��M�`�8��;��Y�;Ǔ9��0d4�B���Q��O�f���� ���p�9�K�/] �c���nǴ<W��+45>���0HI��wvvI�����l�}^�� n~�V��nd��(^l% ����d��l���/�F:��L�i(Ū��Q9��(�a���I�4�цs9��Y���|���Ô1�o����r�|jN�I�OW4��٦T�;�y�{��>�g��P���G�ɒf��3�gϳ�����$)C����n�y^�o5�4�Ϲ��"sG��'��D�Ϥ����;��իgM4�����������\�����y�9N_O���}����6w	(MК���0+&�8�݌��n#��nY���:�n���'���s5�0�`r���+�ɟl6'/Nnl�uw�8��!�6�e��٘p3��y{� �����I �n/m�廙�{�a{t�ɜ��a���w����x�Q��I�m���9$�s9�{��>��c;���6p���C�&��l���~�����7�7�?g��v�iR�|�(���,�ۿ{.i��/%np�!�w��)�N�vA�S��O��ra�Sϻ�~�\*�!6NI6I������<���7�f&�@�'�ü���o2I[�3�O���@8s�c���-�w{��5��,�y��a$�{&Y�y>Νü���>�f�W/gg9�M�>j��������磟o7#����B��y�/�!�Y���~匿���ل=�d�d�񓑇pd�nv�'�y��~�xswL&�߻���s�\��ɓ33SZ�]�0��&����lM�rNuq�e�^7��e�k��y���h�6���������������TwG�TC�	y8p߿v�A�3R;߁�o9�����<	,����6��s^hbp��_��z��_�S���mC,%��j:4�Pe�	L�1M��ؔ��i���K�^\E��D�Xh�277+:�j�v�bu�]6݊��-,�Q��V�����j#�rh���ֲ��e��̲���ح&w�����$ϳ��f�BE��N�5#k\���]�"v��UTp<�5��Ow�$o͓M|m\�n!ƚT� ��v����<�Z�YJ���;Xhae�����nv�t��~z�{��{�|6�M�έ.˰KX��Ou�z%r:cfKZ�*����&��O=ۊ��~�՝�}�~|�H��W1o5S�;$*�;<^ր��qp�.T��$�<�� ��|M��q�i[M[b�����OrC�(}��s��Z�p1��\\��B#�F5 i�8A�<����2G�W�x)�:?��ޞ�)�� �+3�-��hb�H�H��ʫ�3�،���ڧ�Sh˥ݑ�.{�
t�N,ۙ�-N����@�,Bq{͂���6�5�U��UI��B�Ȥ�yE�zx�~q 
u�����d*ؔ�i:��r��gLӳe�Ǽ���@�)2΁�?�� �<���W h]��g��|���XKt�R�ͮ	N��1�����H�}��=�S�|e�r�-X�dQ�x��q+>�3r�Ǡ���@���x�(�wV����"�k�4Ɓ�@g &�%�䈝,����j`������/��uI�T��=���ﶽ�����ɼ/C2�9W����p�5��^e�Ĭ�����01�����`�S�GFP���FN�F�.�����`���6��@�I�?0Bȫ�%��&B9< �3R�u=��e�����Q$s�h��m�#�u����!��t7�Kж�I�t͙��c��"I}z�f%��	Lm��qIؤ�@�'XB�C�K�֓�Q7%�qY�g�����[�7�<f���U�y|%��d��'_�*�|b�?7=$lJ�j����6�#���O�ҋq>���8�7,^���ybzشJ$K�4�f��vfu�3�m~ ]�[�C±�U\C$�G���xx�ڪM�=�~�ff9_�3�(�s�rf����l QTn�6I5n����{��e��*��}�md?���=�˝�x�	A	 H�IdU�FDBD5������^�/���m����om�鱾���v��m���m�m�m��ۦ�m��1�۪���۶�m��1��nۆۖ�o�m�ߛr�m�m��۫G9�� )�D$	Q$ K�8	9� 8�8p�qN+ͷM���6�n��m�6��[m�m�m���lm��m����r�m����z�����r�m����m��ۦ��nm�y��om��
\��\��H
���2)j
HH�r�Jm�ݷ���n�M��m��m��-��6�[n[m�1��nۆ�m�6�m�{���ݷ��6�[p�m�m6�o�ۖ�o�m��m��oԠ�IT���Kǽ�os��{���6�o͹m�m����m��6�m�p�m�m���۶6�m�i��~=�{�m�6�m�p�m�m����x�m�m����v�r���BA�	Y"ȫ��$8Z) RVIQB@	I��6�r�<E`�0�#��=_�@���M��?��/�[���Ӈ�u���.�˥�0����3`�ad2���@ΒQ#:"D0`�!�3H�2�xc,f6,3�,��3X�c,��0�Ktd�c�ac a� c�H�te�fe�0`�!�2!�-�L��ѓ�N����ug]$c�3�d��1�2Ft��1�b���F1�f��X�&3	�0��Yc%� ec�3�C<1�fY�p(a��ι?���Nv�c�Z�m�[��l�]��E�4����y��Ζ�B6���WR.�	��ĚXK�fИnѳ��3�OK4�z�T��ٯfU�Q�;V.N�m��M(�f��˳��7B��-.ڬ�.t�KMn�\:���6�11k�c-���GE-i���hF:ٔ�a\Fy(�eF�S�\xf,�ѭ������7_4���˳I`�:���Kv��O��앉�A�4 �����fҵ4�(� �v�5fq��aƶ�+q���3W��>�F���E��m�����)Qһ:R�v���Q�3���JzTv�-�bE(Y�n�����[@Y�)v�3�A2Ci�Z��Qc�mM�jKc�)��6SFjA��m�K�^ҕ�k7�ް��C�ۓY�!�kIcZ��6ͺ�*�X�-�j���;m,�[�ڭ������V�Kv,t$�����i6-�t.$q�
�j�j�bilHK(�;XMv���v.�JћMv�2LS����;5����9�Y�4&n�%���KdJ�4$[mAՒ�k\��w
�y���'���;mıc�/j�V��33,R����EE��U
�:cGjЄ�6��&��TZ̞���$�sQq���˨K	�&nAI���.f�)M[��r]��J�J��λE���K=�����2�έ�MwY�^�iY]�kvAHL��^	\3J�/�����u&��֡j�.�[��.6e`wm���c��#�6]�p8��n7JfXlԓkvЮ��ˬ�k6�Itsm �M�M��f�cR�̋JMԘ��h�,Ԇf��ֵ�&+11��Hѩ^���at�i�K3+��,͜���8B�Jgb�l7V��m����	���K]4���[R��FWnbX�e�f2Y��i�)j.�r�;hK�!�[h�V��e���R�JY���JY�d	zʄõ�,n-k�P+k,m�l� ��[G[5t.��M���|��kX�t�vg�Geu%89�NO�������7��V����n����9������m��߷�s������n����p9��Q��M0њY��fxg�2FI�V.���uf���i��Q��Z��(J72�l���PYv� ei�Z4���9(�f�m1�-�
,]�Ƶ���aJQW).�.�kfl����3\@A�:�!�+pñ��A��G�#k����	P��-Gj�:��ػ�Y��� �hg	K�Ha�KXd��˪����g�i-y�m��h�sCU�asٕ��m/�,����f�Q���^	Ov	���3 ~G�C���m7�xE�Z������&[}̎V���a߃��������C��;�s�&}�.e2����/C��e�9��4ɞ�r�T#������aNXl�0,3�����M̀@�F/*�D�@�Z�z����#��ZV��ag�4�Ɵ<��,��3<3�#$�
0�=� �{yC�f�&飁�;�CI�6C'��jw�N~��n�v`S��M5:��4�ٳ�WN���Vh�-����~�eY��6��!Z���7֎ͩ�$Ӯl�=������Iv�o�1Lȑ��4Ӯ>1�ac��጑�a�.zFH���3Ǻ��	un.�Y"����Hf���kE�);��kb��RS�3��8����&�(D@�T��t0`��S���_i�c\<�,�����dd�!�p���N�>��۸ma�d��OO!�SҞe�gi�4��+�v�S岔�,t�fe�X�ag�xc$d�aGnpr��$a��T��=� bO�*���T����RV�Ι��Z�賣D�R��P���zI[oH���u����=M��X�]��}N��t���פ����B����O��rEe����/U��4�QAE3�1�YC<1�2L0�8��L������]/�+ ��1i-�16�Q�c"���1�TPJ������S\�e�ݩ�!Q7�\�&B���%��ؚmph��SY�VW#�BJ���1U�RQ�l��cK�w�
���%"�#0����m�Շͭ��l7Q�.�ۧc
z}:04�鍶x�!M+�%>y�}�i��b����.0�4�K�7��{/��q��[��߳������U����z%Y�j��p����0�	ã��!�Է��q�l���q�\u��C#$�
0s1F)<Δ���=⬡�6�����B�M��#��þ���,>�C��DOI�֘۠d�⦉��寞g�#�a^�^�˻`�ji��RA�3wS;��v�ek&����~�v�_�WL[O(�z�u��/��Da|�2
:t�aE�`�a�0fP��&Q��fw�H3���#Á�;�S�L��X�v$|}M4a���ۺ'i�NK84���I�@����S6.ԺnmgG~����z2��O���f�)3�L�P�6�+ ��0W������1V���S�3�����Ə<e��8���N�u
&ޘ���w��=T8�5kUʸ���s�x&�KoA�;�!�A�S�0�|8*�YW����<���u�q�\u��C#$�
0c\@t���[IGKW<M%z dR&�T+i�!-v�M&ݴW32:j�g�P�I��=�V�\��+Z�xDf���(yڽN��.����oΓ�x�Ą�Jf�]u�X�ܧ�ݥܹ1[�P�d��)�6�G̴�κ㎘�,���&Q�����JVz9�F\ǯcێ��&5#Wl�y"p[�x1A��I�5W�ץ��)��^��·�k��+j�)�w�+����z�qs:�MMWġ�R`H�a[j��̾[�Y�n����	��=ҽ��8���3�J7�X��,��ǵ��t�.ru^<��w;��K����C�*�a�J.�xʢ~x�1&�39��3��ə="�MzeA�#��7��c���;!;�gE���g2�˖�̰�rFCӸ&��{��c
e9���M�	����(Eo����yu���yJ���D�Y��a�1���u�]a�q���8��F�����Rҭ�(i�rRA�ϧȳ��)�?yx��==׼̹fhQ��n/�Rv%zO��d��C��:ڵh��e���E�x������.���)��]��~y���ݻџ�}'|^�h�=�vW�^��<�����E��mxN�O'�l�O�F����'�M'FF��C4��F�
��%b?)�E�/�#�)l�c/̲�~'���.�a�<^ZF�G�#L �`�dH��1i1,0�4�-0�0��a8i+���#��4鲴�4�E�0Ӳ-�F�(4'E��H҈�J�������y8�x��"�O-v�'Ɩ��(�4h�|T~��~)~ak�_�_������K�y�_�חǘb�̢�O'��/�������ǎ�/��'�Y�&M f��f�'� �H�]�h��d,#L#F�dB����F�I6V�F������4ZH�Y�4LO�s���%ɖ��mp�Sd6HK��|�་2Z�[���W����!�y���ʝOr9��ϝ���www��wwows32��n������̼�n�����ffe�4��c��4ҍ5�^e�[u��;i$�f�]U��J��!�%�J�uD@}��&N��4dDI�X����A(��BY ���2%�x��B�E򔪧GF�L���U9���s�WD��JF�X�ԕ�[]��9	��ၰ@0;��6�pD��C��Ō��+h���MP��" �U�V�)��+�Wz|'�!�'V�«���@��Q�@� _�d�!�4�Fl;(t����I�4N�FHw)C�Fҕ�V�%�=H���Xe�ο<�`�af�t�I4��0��\Agʪ���A!�3��Q�o:^�� �����ER� C���?9���pS�c604My�
ŏ��RE���X��0��K�57�2(jb�@�T�GФ���Q:,D\���~2�M�(NwmK��8 ��HQ	��չ�.�0:�cD���ARL:�)?wߏ���+SDB��!���9��A��O��ú�m�U|:;�
��=BbpA-$J{I�b�GU�Q����6��:���>a��i��Qь��}�:�%5�Ժ����X)�	�M⎊AQA��H�+"�{� Ɋ��s�p����`L$~�%�(t���|Tbn*�cb.)��������:�r��T�3Z����� !X�o��[(��;�z��Nq�^lT��@�Q��,.���Pu�)���d�z��s�9�1�soqN��;NY�I���!�JZ1Y]+U����u�OD���!���VHuԧ�E,�	��(�����q�F@�Y'�d札�80����'� ��(��	�+�Dm��7���F�ʳ�E���`�Q!��:���:�������D:�,��4&$�S�"y����C�����@�f�.ntM�ބ*ftp'̒a��'�$`���aDa1"��%W)��Ī�y3�m)�O0�q��3��i�i&�tc<29���*�"!1����2h!�h�""T�Kd7��Q�����v�d8 z"&0�2Tؖ"�=>��vJ"'^R�/�Wߘ��멡K��%m�о��hx�a≨�����B��*�~�rw����O��	��Dad��t2o��ہ�m#��]B���Sr��%8�N���i����j�xǢZ�\�3.��$�?2	紑)a�e!�Ʌ9?}�u��L�;g�	�L	"[gp@�҈���5��`��pJ���\i�����8덺���/<��2뭺�����$�!�!4`gͽ�v"%@��х&2��AO h����B�.I��Aa���҇2�f�"DaD
��"CFHs�ÌbB�:�3���u��7*�~�B�;����Ԍ��'d�1�9��C�S�'��@�`���%��d`��Ȥ���):�ȈQ9����@��V⒜���$?@��G$��# �>>�2@�%"��%��pDN2N	c%�O�`c 0��fDN�F2IC�YUR+����8��O���:��:��dt�I4����ʿN���"0��ȓ�Oǅ�8�t���A�D���s�8$1(����"\�.�=�.�l7��/D�µ���d� &�������
K?AH�&��G����{4����ߓ�(�A��"�'�KE���4$������bK�� �L���'v�(��B��5��pE�BT�L�~0����B�E2R��,�h��<ߏ���CF ��#�ό2r	��E��'Q�ȝ����+�(°�f�|����:�n��o<��0Ҏ�g�|}�R�Ga"&*�Rb��I���ϢE�u�I�Fe�1
��xy2
|x��Q;���"5����ڎT�$,c��,N6䴎+(�"��  ���?.��9��j��6�~ �v4߆�6��w��L�m{��g��5gW��E,?	��H��BT��K>�?	�BӮ�~��Ė%A�Me$��tTO�����Y�H����-�!��g}Q�"0�r� I��=�
!�>ȇ�c��������}����w�w������L�u)���dM���/*2j=������S�n�k4��G9�s��d��l�y����o_��9��:#�8Q̹Òh�1�t�A���`
�*�I��U�>G*S�ό�6����ۮ�[�2��<�.�ۦa$�_��KJ=��}������'���!dC�!�d�f""�&��?A*�O�3	*��"2�L�J�R�D��L�	�i'�N��ޡ:����Hr��F�������Y�)�jid���p�!a�>N3�1�!�r�J��7Wz&�V��i�(�E��)I�# ܠ##JO�NN��F�]W�����%���C��������g���N�>-F"�*<�Y*>JH�\9H�lY�>>0f�i��i&�tg�G��'_*����dd>��5�����ꓵ_��2���8��+d'y����CD5�Q*[��f�͎����h	z{,LIדwa�	P�0���Y	�	�g��j,�i��������9�k��Ŧ7����{���9;*'���!����	4C
t�AL���^Ǭ����V�WUƖf~K~Eq}L��匐�5'N3���<pN�;��쓯�����	P�``���p��6!Y�A���������*�==A�DHpa9W\$����['�~y����0�Ci�i&�tc<1�p�I$B}1�7�,��Lr!��A��Œh�Ȱ',���o'W��uc;g�l)� �z����������M�^cka0���S�8�El��*�Ҫ�R�6�q)��n�	*���?�Fz���
��T���(�,��`�1����COU�|<���?	���n�~��)���4�d�~����O�M��其c=(��l�����0�.�+#lB����b���~�M̝%���2��%��`w��h��<.L,�˴�����'��6��O/ͼ��#4�4��tf�f��H4L�4�!6�M��-���//)����y0�����1�y�������虰���C��A��J4��K#L#Eb���L&��iD2,�$��??1���~_��<�O2�=s(��Iӥ���xZQ-4�tX��������h��+E�j��D�����������iI*4�ZF�L��i$@�:F���5)#E�J�di�>>#���4�Q����#��Pa�1h�Pɴ�#G	a�`�4�6��x"�!E�I�iYY���	���Ԭ��>�H�;�6���Ϡ��9X��F�����e�b�f�Sѭ�󋸵�x�M�Wx��&I�q��ed�ଳdpo+���]�-�!1����^�Y�m��٘���ۥB���3����)�ISʩ~�j����Ù�qe�,i�$�`
!�?#��'�$���?ev���V8�{2���g-/"h���ʹ�_O9���Hͽ٢��=q��i̊ޑ�l��wT��Â��$��Z�q����T4V)�ȸGW�&��8��d��F��وEN[�ݖ��)f������W�OZ]4��R7�o0�,-%w�}K�y�M�N"*���1֢��]�����]����JP*�~���b&[Kn�nl"V̺�[��	Q�Mm.K
B��ǔ�Z�n���&�<~��R]abSS[u�]�4����.��w;-��9���e{{�I~]su�)x%����_v�ڱڔ��#08D�e�&9���0���G�Wff�����fff^黻��{�������n�3337Mm���fff_4�Cƚa�4��x���4ӧʪ�^�^�OZ�6?�9J�<�^���Fj��JY��)�C<���lC#B�UD�<������]f:ͩp����\�F�M4e�0�%�+���Y\bۡ{BJ\�#�p��TZ�rvyͤn5��H!��m���k�����OK5e�mn����2ٖb&n!�+jϫ��}-��-%��#f44ɚ���Ci����,؛d��[O"&
)![(�\ 	\��E�H�m�4��Y|�F�1�`�hʡYV_�����-M9uk��r�t)C�w�/����N�a␩�L@|�`�Nsų	��$8R��'D�AH0D2#A(�-i�oŇ�Oa��=6N��*X�D����LC�>��=���0�""2u�E�c$���G`t�d�J��C��0��!��4%՝���h�d�Rq�oǟwg|�D�e1�����[�������/a��z����2��X��k���f��]|m��~y�q��:�<�̼�.�ۯ{7�W"��"%<⪨���ɽ���A.N�q6D���ȫ��)a���{�:
|ak{��t0�G�������c��t~:�t�����*��2>�K%H���Z��/��︶f��LS�$����Q�����-��N̒xv&'<�m����4��a��$t��(�aџ|`�<P��F�i�N����̌F�I$����uWz���g���Ҫ)�?vY�0v��5�`��I.[L���/�d��?	C�v�R��Ta�.��)	�x��I\�����Ƥ3������H�}վ�[d�J�#)[r��5&�a�4�6�f(�UjV#�u9L���O���m����Í��[wu%8;P�$J�f�ױ�5%�\�4��[y[>e��??8�0c�4���!u�%TB�s�W��S�FE��5�,�q4Ҭ����'s՛�GQ�\Z�s�.����
p� ��,���{~�${2���=�~�p;�4Ã=ɁCɅ2	C�����,���d(^Fxj����:�)�T�9U�ϷM6�H��Ƙ|`�x����4餝���S����eMF��Ey�H��^f&L�L �7k1'dMS����NMt C�{�X���12���7�˗�!�I��fL�ZUmpp[x]�L�͖�SgGm4Nu�� ��ݴ�,�a�[2���*�C�D�&�.ef�)��cz��7�٭Uo7�F�����,�в�w�9���ٰ�����9��`p�n����r���C��x�զ>I�r`o�~3�y�pNÓ
i�R�o5�%�m�t��S̚"�N�~]���)�kROW�O5X��L�^��/u}/�8�q< 5dNLi��#�ڴ�o��vS�N#���e~f��w3O<�#oϜq��]m�C��4餝��C��g��k��v-�]��g�>~�.w��~G9S�  ��ђ	�Xa�Ρ]Tv��kD_V��|j�$�0��/�}t��0�hCJ����xbW�:�O��7%J��u�y�+T����&+��y�&���S>\�]���;)2:xy���̹X�~��3̓a�����QA<4\�H�f��D"���L�����ٳ?{
t#���̷3��]4���8��i�|���u��t���̼�.���a�nI$D,�0�3��Nd��>�a���mi�m%U��j�׫�}L�C�{o��g�6cz�R����@��Ļ�`ֽLm8�*�5L1]�k�/����G=K�0�P��C򩿯��X��>x&+"������Z������ywU:���5�k����b��:�G�G����o��n$���Y�]H�a��]q��6�_��SNW*0�[�n���0����0c��t�N�������1!d��?y�p������m�"�m�\����\`�r?�����]ҕ��V�"x��S��'`3Tx0j踄�Z�u4%ly��3��~����N��/za�+&OS��}�.�R|�>]yuj�ӌ;�'�Hs�>aG4�O�S�#'���w��~��t��)ՙ#2]5K˚J�f��\m�|����:�e�3M:iӣ���"e�z���L��JjZ�Y�?K0yəTn�ʞd��Q9���bLPI=4��V�9�F�p��X(�&\kF$A�nն�� [r���Zh�)�c�Z~]���1�kJp$��9��M��;r�miW�'F�N���t�=���+��op��iOdC��Q�d��|Ċ�%���bw߲��.��ag�� ��O�V܇gga�:S�v0�H�Ǚ���~\^��#�*z.�ن�zY���9'�����7�x�Sr��7 �8��,)2%�ʻ���N�v�Z������}MS��ç��>0�L�0c�4�M==:;R�⪨�
~�~���F�+d��6��u�u�S��;�f��(|� V�#�x��
G��w��*$���]T����������ͽ+$#����kT������j��,�_�b)��n(����+�G�J ���+�*$�m6R��ͱ��yZN�궟U[�α�?I.��$n�#%UQ*��.d|�O�/	���˴Zu���o%���"�4�E�L&�#"M�Jf�����|�&��ܞq�M-�O/)�o.4�\yzy�<�fK�<Q��dh��4L�L�#��Ţb��H�4D3H�H0ZaYY�ؼ)4�z�)#ai�w�i:-4��,��G�W��X��O��s��&^_�m̵�����a�J�<�-�0����gŚ�iDt�N��~)~2���Qi$i$h�F�Ɠ���)����x�ic���y��i�:z�>�H��e|tަF�B^4�!�D� ���tdtXiG� e��eqi���4�*4�,r��MKHb��ۅ�G8�8VI��DE���ē@�D��CP����3$��fe��$:�@P���ē��ZB�$�9I��R`�BC���,��"�2�@_��k+t�Y�����31*�3����;��������*O����p��g׿}��ٙ������������Z�m��fff�m���333�ҍ<#M0�0c<P��C4Ӧ�4����UU�t���Wj�'计��W��7.n��[�7_S5��u�w����2	�Nó�L��֔,��j/5��	�U�m�����I]��d�����2�\��0�[��g��\g��g�\Y�^��X�4Ԑ�$�΄��K�Ŗ�9OVY~m�y��u�m�N����/2�N��U�^��H�+8I��˩�bN7*�_�d�����V{�5�����k����j��0��/�>Ny�6��ۉ���Ϛ]6��F)��uU[m��l�߄�*U��q����N���3��R�|~��RVi��>~��Wk�j)(�DD@�!D��O�OHæ��-�0�??:��8�m:u�u�_*�X�Z�d�|���1؟���@�R�&�+B��T����kÍ�Yǋ��~٢zc~P�n)PTX���RV��ka�;;k�l�H�jZN��  �ŉ����������`��x
p��W$
�cĞ`�J��S��	C�vT�� �(�h��3��Y�|`���,L�|~)�����wOe���
�C�
S�{Pf�ӎ�3K����&�Sh�\MV�۔�>�yt��g��n�)��!�4e��3#&+�<g�#����:��OD��$N~�R�HI�a��<Y�`�0c�4��O��Ad��+�
H?���QY�B�(޲2(F2E��# (U@c,L�C����E$�����'J����P��AI"0
""��f�yu�j��ԧ���v�i�_������t�C�xv�:��z���è��� �#��џ�{�'{��$X���D��R���[�~t��+F����ˮ,J�߻e��tâ�(6��9X,��� �|w�{hEi��qov�X&�&	p����f�#R���'�x7�r�D�a�6^�~�<屏�䆣l
��7{�3�H�=���'�FU�3h0��L�H�u��Z]��UU�,B�-Hޅ��)k<�A��H����)`�POT !�IF��T����w4�E9Zp�B������T��Ǘ�n��Һ��b��� �Y�KZ%�:��5��f�+R���ɖ��l����2��i�������P��r.�`:h��E<kX��6�)-��ୖ�Z��.��mcWZ��~�5M�W���N~��z~��q�������W�Oǥ�xC0�L��C1�Ӧ�|p���ڪ����g��i�r�X�#&�_������~[�M������>���>*kTU2�ƎR�m�ݸm��ӹ�
'���~�i.=$�)�Ϝ8��q���֮J/�m���Rb�+�m�^���|l�6����ܹ�I��VYr�=L/f��Y��,��L��C1�y��u���߱RI$Bߘv�~Ft��G_6ۏ�n�"g��쯮T{�7��9
e�W8S\0Z�Tm�'A�O!���N�C}�w�)*,Q�;|>���A�_7�8ˌ���2gh�$�&Yf��,��ǩ�j���I��yq�ȷ�A$�I ���߸1TB��3� @�\�p�8iF�D`φ`�0g�1�f�tӦ���>[��c����P�"�m��낍)vl��D՚��<����6�ո�L��;�l�U\t���TiV,�aB69lt-�	����,}}�y�Ey�� !'���|f���ñcoV�7��6���j"��E>]r� �j�4fl&.:n�f�K�mrN�
��l񊊙�-�㻷�̛i�#G�Z]VQ��{�������kF�����71w���V�!fi�����<y��7���SM����]:�qkot�+����au���xq��F]�[͜D3�H��l�T}��1+-��4�z͹�!��7��2y?n��ߤ�a��Yf�i���x��C�M:|zpL}k|{�CޕUO�4�'�'�l�+0���0�=>�!�t��� �|�l|��Q%�pG�\,��C�"�_;���H
��h��K;��Z���Hys#�c��<�[q�.U�|tS�~:�8u�q��ߔT|�øo���.�M8dJ#eӴ���o���:㎶Ӈ]G]y��y֘t��ofI$�],(���`h��}��=�tF���dL����&`��ߧ����		n���_/�rTC�N�T��]�N�D���{ǈ�3�K��>��Ø���*vp�g���$r�g���RN�u��v���UθDV���TG��Z1*s	��arq�g7�ZC5nkW/U��O�m�So��[�0�����`�0g�0�1����4e�I$ �Y�i��L�#�?�x�~�U��4���%�ESO�r��[Y������zUO'p�{<���U���+�^�y��4��(�||p�������p�SGz��tӁ�,���a����i�,�L4����o��k����av�Kuh��-�?1�%�������4Vi��4Xi���'tL� ��/��I>O6��m�'��<�[^
!F���#H4�,�t�^&V�e����h�ԙ]��D�i�;�"M*V���=�F�i6*B�����i�����6�lZy���<y~Z���4���ߘ�O�����r��.<�-�0���ˏ,Չ��iGA>��ό)��ʪ$�$�$��H�-�����4�l.i�<�����GIҏ��Ti�߆G��Zl/�����d/F�bZC��E��bZ2zd-#�B�Ҵr����(Z���҈�Q�ʳ	�H�h��(��o��f��N��&�L6!L�Z��d�B��Y^��wq��nS]m�.n�W���f[%Қ9��g�q,Ў���Io�Y�����"ˁ�*���k��7��h��)|NCƣ\ȩ�4��j)�J*C�}�1iNbʝXH(��ֹ!ׄ
ɮf6g�#x� �c�p�c`�2��6i���X�]̶c��D�������O�Uv-�
�
�N�q�#�r�O[ŮM<�D�A���(�h����=|�|�Q<���h��-6��Y��������4�����I��
�*�E�ޞ�7�jO%R��u���sl\�Ōod*D�ƥ��~�<���w���+"$����7&VT��c�|�ҳ��v7isl��0�e�	�"�2���ZY
�#~T����\ۦ�J�Ym�:ѴQ��PZ�g��*���q�u�}v�S�<��k��i�J���[������]��MfN��R�Z�R����v�Z�Q��|��L����1��_ٙ������˽����[����s33wV�m������(�Ɛi��3�1f�4飞�������IN���-��%fs��m1e�0���!�F�M46KlM���X�e4��[�Z�0�]K��ۖ��F�ŋaT)L��6ֵ�*�HoO�1��ɸ.x�KX�#�.�ʆ)��mc[1��E�#�&�4��0��k��W6୷��X�M���8��X%�n�lسm2�� %(V!�ѿ���`�N�0��2B�ͬ�l{ޤ�S�̥�oԼ+w-��ó�sD<���E��Ϻ-�~�GA�a�;�g&C�Y�ǉ;�Z��>C���}K~������7.�|�xv��� �҇�m/$��;_7_>W�Q�dޱ�����ɸh�������i�K��!�o�z|!��3��:�̼�δ�I$��IRJ���W;���U�����M���	0�vaN�(��D	� �Z�C�>���?(S�����[Zvp�&	����x|tP���_\��.4P�HS?v8�'�����w�}��6��>�G�^�����5���dܑ�!����ꬵO��N|��w#�G䦜�/��0�φA��0f3�bיy��~��{�R1��$�r��זּ�S��,?���m��4�{�[a�u��HH��E�A,��ƾ���+#c~H6TT_٫M�M��n	��xtx})�C:$���j>>KlV����t(�I������0�A����Zi����쥏S�=��������o�p��F3Y���a�<Q��!���e�_ܒIXZ�\:���V�z�f��Պ`���u��/1&�X���p#	ygT���&��~��:�����o�ny��nT����Q�}�+m}H�s��I%����a�����	g��lzQne:�Au�.
E��Y=:tDγy��\�'�ǽN!��6��y����t�њa�<Q��!��M:h�bS�\��<����J$��>c����i�Jݞ�P)j`��4��('_E��3ƞ�5�vK0[m�b�N��P���� I����?b��PF��yG��3�f�2���u�r��ڷ���\.�S�Ȣé��;�
pқ[������$ϿR݈�2�L}!j
k��K�$����p���=�w�p;�ѧ�~��<�'�ن�sa��Բ��O�e�_E��-���>�q��I<'����8�%��j�<�~�?C�6N�ؙ���s0��<4�좏A�4f�`�`1�c$�N���oYYϤ�H�jѽ��~��j��r�)�i��J��&�o2i�ے�-��i1�r�$S�̐��{Z+��$�m�1M�BR�k'�_���J��
�C�d�\���C]1��s�Q�N�L#>9'r'f*S �^��w�'�?V���'�b<|�Wb^(�&�gi6�ێ8ۄ��f�`�`1�c$�N�3:,S�ED�UQ�������H�m���LS�a�5N���,v���é�(��3�K������ ��z(J��~JI�<k2胙��wa��hlD>����v��i_N�\�	�9 �	^�1s�s�>xq���4tI؜~��S-���j��]�+S��ͼW&R��w��tyo]e�2������O�Ǿ�K��I���aߩm�b�j����6ɕ�C����8�ߞ~u�3�b�4Ӧ����g�I$Cч�Ӓ֗�O�?C�p��OХ(r~��Z�SU.��n��ێ\�Wa԰��u0����$G��5���?S�-��1M.�n�SߪO"4��Jx���z�~u���g�~���z4n�����a|��c��$U�#�x"�
';ٚ{;�$�e�LS��-��uź�μ�x��C&�tљ�)�]��;��5i,ܳ����S�b�*����c\��3ra���BK�����{7�kB���H�,�~ 	n!-�9Ӎ�QI��{��x�Y��Y��CF��7��^�.%�-���#]p�����T�&jݧȳ���-��]���=�a���'ǫ�ͩ�����"�Rw�����L�b����X`�D~mY�ъa�^�6���!�i��4�ߙ\d�=]�2����D?�>����n��)3Vƕh�i���d���0���>�m�Xg��Y�> �M�3�b��M��RI$�sdL���r�3V���{2%�?2�꺽Sl?N����L4�АY*��cI�3P�-��u���2h]<��>9��M�Oԭ����ڸ����[�3�[��L�z��O��]�Өɚ�c	�WY�b%h�2�)�-�5�%�ݮ��u���j���M�F�������#$�ь��������1�1�Qg�xC(f:1%!�
1�gIΘ3�Ό��a#�E�����eg�x�чF1�c:3��:`2H `��C#ьc-�]|�]y<�<�x��0���ͺ�V��[�un�뮶c0bB0`�2�єP�xc4�M�4�L(��$e���X�f,d�2�a��1��Q12�-����r���5%�S��׳q8��^���bi�֚�u��������G���mG��b�Ì�nv�8�s�so��Z�<�Ct�*j���}��T�ǵT�5>����̏o�}�e���������/s33wv5��e��f����y�{��0�OY�3Fi��F�2Fi�F~���J!2��ul>��1xqꑓ��6�?���u-Ӳ�����ro�)O$�O���`"!�bR�r}8e��˪����evA<(��Q 넟#J&��E���wn1O`�W�|��?a!���vm%A'�a��u��r�:���y�P��-��.�=M$�G!	�����$�3>4��A��4�x��C#4�9�Jy�����UD9
����qk1������(�yl
#� �m	����#�w0��}��i�K?���H�Zf�����Sߤ��WM��6�0�L<����?}u%꾪�Vߖɜ6�(�+�sO>� �J�|������#��/��-ӫm�e�<�&2�4���Fi��E��2Fj���3�ߟ�4%��6-D�m+�J�p �j<�]B����Q�M�n�滘ߜ)۝�-�Z�Z+���~k��-i�ή&� �����qU�s
��0�#��  ���I�o�aٚ*�lg�؞��]a6��R�.�m��Bz"���(��G�OY��g%���O^DG��B�x<X�I�������A:{S����w��+���"=Qp43��oǚ�i�dGk9\��L��Kl�[�7��3L��L{����]e���ى�TS�`m��mmώ�O�=������tx��a�f��F|3L0g�,c�H�:h�,��DAI$�A�V)���G�:�$�|�ϑ��`4��,QO;���>�)���g���[�����Ƨ���,gI�Z4!fNM�|0�J1�q?�3�s��T�=������$����`}4�(����+j,R|G(�#�ң�a�DW}���ɑU�UJ����WP��ַPo�.y�#;���>�mm���C�i��ӂy�P�gQ;2�;����QK�=���|Ag�h�$��f�`�X�!���t���6`��Dq,���esf<�Ub'Vxd͟)�XP𓳺t�t�6�I�(\��Gx}�oL��N�i����N�b�v
b�\k�^�N(y3|W�$O�/��4>2S��D����N���VMN��6�������7ϥ5�B#U�_$h���ߤ�4�#�.�_�)m��[.4����i�3�1�c$f�4e߻ܵU���ǅX�f��A���9�I�{���Jaci�f�t�8[j\Ů>�t��6o	�d7��u&��žF)�VW��+�-�et�ϟ0O�i�+l6��8��̮��m�I�4���j��6�%i�h��R���Ut�:bi�I�
4�	4��L0g�� c$k�W���Y[�H�`6���e���Z��b��}|���զ�P��
b$R
�ޖay�g��������ƷD�B̷gT��II΀�ys��\̰�ٳƣ�m�һ����r�].�އ��z_<�/�hw��ĥ�[��.�N��ǲ����z�Eqe��1Z��DG{_s|�+孲�����>��;��~w���xɪ���|�����Um�M+����ۓ.;I�X�'"1O���3Yy�ԑ��g���~�DR�-�b�f���I���t���5Q*\�x/p�"p�S�a����k{=�k �
,g�>$gƚa�<P�=0����ӱ�O8��`����p�#��{��b��ɺv�H��+T���Lr��H�=���������"~�2z��MJO�C#�s���⃥��p-���sS>ҙ-��6Ү�m0��짐�0D�هK��v{�m/��Nħ�Q2h����N��f�wlE���&x'c+�:YE�1�Ӧ�i�YC0dd�Ӧ�sĄ����qZI%H���HI��w�Ć|2�\��	��G�)��ΰ�8�kF�}�}{
>gȁF�܎�p���_M�ã�Q����Zͪf�R����ASʲ�E���QB�~_.�6���"��w��}��qK��ދ0��N�Gb�g6.��s%����W�:�M6��2�Ƙa��3@�H�4љ���I%�M��ө�-�*z->(��h��~�A��X�0���%ʬ��#�BW3Gr�nTDZ�S�=<<���O!����"�v�>?d6{�t'�|�$P�J7���iU�QBϏ��F���ks���'�~�Ķ�$�N_��J�;�g^��=�VY3MUQ���̢ߘ~-?�I1��A��ҳ�,c0f�2I,����Ptd� C0cΒ1���d��`Όfұ�2Kxe�b��2�"�1�2�`�t��$���1d�c(c�:3�IӫGV��:�&YDd��ƒ#I��3���0c0��$c<1�a��f�i�Y`�3aC,e�tfX�,e�(���H�bg�YC0c,�F�N�_t��	!yB���vR�rE���4��)`�GQ�? ]��6���e���7�S�{M)e�hM�r��$��͘l<#k-���{��6��{Oh�T�j|��U��[pс�f,�J������G��L�m�Ev�H�kw)[����*�Mk&P�i��RB�l���ㆴ��"����_���L,8YwڭE"����d����l%��u�Hk�v�gMn|�O3ơ�S!dʈ,h���Q4=�9��[�|�×�9�u\�4�	▊��A<��Lm��qU"��W˙�
�P��g-B����Vl�v�v�&�9,�R�rк&�B��.���[
R����ێ�.ĥ�cv�}���LnE�K�Ɗ3�Il��$��T�m����4h�ҺSƬ�wj2�X�����=(����g�o��I��v���	�Ӓ��Z�pR��jN5h/_wټ�3/����ݝm�̽�������������ݝm�̽��(�Ǎ,�Ft�M0�K(f����i�<,O8����f�[f�Ve�ks���T1�;D;A�Fդ!.YqHKa�!T5��s28�5{Wb���uٳ͔�5�vKx+Jm�Bݩ���b��֒�+4���-33]���)�������V ��	Y��Y�m��V�Y��e�� �mp��Uf� @n��$�����b��4�J�3�5��4,��Y�;� x!IVYt�2�V�B	�Tױfy�!"��dخn��S��#��5��`��%��R��W�<h�L̩]BP��J�t�..QZ�ny��<=�=?l�4N�⣰�S�0�m��n��5�ݒCl"���s��:�~:~m�|�N�����-[nrMS�0���S�}.��{@���r�ԢuTE
��.�<R�e$q�-�z�f�o2{�i�i��L��M��3@�$�M���$���(b�2A4x�H��/��WǛ�S+�Q��"S��!��@:Kn����]����<0����f�	��:4��J'�����pţ��z�*��_��R#�aB���s���Jm*�t���|���N#lb�%�Ȩ�aB�Aѝ(����h�4����q�y���J�nI$���wf���^+�մC�n?0��p�x�\۹��,EUQ";���6r�r�DF0ޮcq��W�c�к� 0Cd��X�����a$�r�����0')/�,�Z5K��|�z�ӷ�6�9~{�N;����6~�<3��C��D-�Q��"S�ݮ-o��e�<�/�<3,fd�I�L4��� )2�W��Ub'ǰ￾�GF���%��zl>�Dӡ:����sUp[�G�$l���v+	]�y���5�$�#>���0�~�"ĉ���9bJu���',��mimr�JWK��~)�l:�4ɓ�E>�&f/�ͣ��{H�oi륻YagU�,��;�<�;�E���<X�4��M��32L$æ`�gD-P<�C,r>�Ye���S���~!#�"m�1�
����
ԮQA��q瓒�]o�(�G[
��:�����7��[��K��: \�9�!����q,XY��S뚦Ҷ�'�bn�T��Tn-�q5�&�Dn��>a���2�:���WpO�`�����\n>~�a�G�w)��EO��[gYmf��}=<E��ÿ.��B���_�o�<[�n'U�Il����;�u��2���T�/U��g��m����P������իW�B=����M�?q#9c<X�Y�4�M4fX��0��i�ڻ��d�����	�k���:<N����Vl8"~��2����	�&2ÿi+g�d��o~x�<0�m�=��1Y��h�c�Y��$�:Z�j�	h���%��ʘ'�<:�wƸ���_$�Fӑ�P�n�0�Y�����0���Gƚ3,fd�I�L4�؁JJ�0�Ȫף��)�<�Ӏ��������߭�!�a~��7"�/���F{#�:�xOݔN��~��6qj�3�ZV�^��_���<�ab�\/��(L�>�@�Bx|a�B��9P�YX���K�W�1e��eb����N,'$<�V�����Ǩ�_��,���2`�)k������	kpKA�.��%-�{�xra�&���@�=��I;⤗ro��P.;-ғ,��'�u��b��z��1�&�[��y�s����k2Wk\���D��NG�cc��e���� ZN]
�2�k�~�/uE��%' /OfLC�S��"�-TƘ�imT5�[�߿s�xݲ��	UT (9j�k��y�F�>���k�<!m�-�6��m��b��<|��1�8�yd���&���FLg����PZ�[ʚ\�i����o��vY�`�ֵ~�g�JX�aZ���e��Ր�i��Ok|++3��jF[�6=�z\�n.�G<�(���'!����i�k����4�?/�n��a��_(��h�4�M4fX��0��O���ŀ�,F"@X�
��)��a�/I%@b@�(2���(�`���@E�J��C&ud�&0!P�R,֌�����B��P""ȰP������T���VM@;�V"u;8���7�?��<=�0�"'g����Oٮ��s��uRݗsF�1�r���k�'�S��Ε�ժ[ZO��3�,��G�M��u�
w�e�Zi���v����J'D�}NS����.�WȌ��L�����w����
/�X��R�#83OQfi�i�0��`�I��t�L3Z�P9}|� ��(�T)|�KN���B�qU���@����*�
z�Z�U�r��)y�6nV���q���H����ϡ��Đ�#|3G��}3H��Q�5��U�q?(ѓ	]�N�ߏ�V���`9���"�)+������ R�I�=aa��(�1�����]?O�FC�e�MV�1�����FQ=��5�F�J�[�~̩<��|����&y
S1�Ӣ�׏�W�~�഼�wTw.e��;'b"v%�C�����ۍ���O<�<��u�q�<��]I/I%DyN���yf\|�s��Dz٬��~�b1d�#y�~��~���ARMSMqn�W�����=H��x3�r�$�E��艂�HDѹ��転�����L�S���j+���tQ?h��S&�}������L�WWY���ken�ya�L#Ǐ-պ��u�u�̶c0f��`�.R��xC(d�3F_0��ӧ[un��Xu�]u����0fь�FX�gFxe�2��ђ2X�1��	�1�QђH@���2X���u󭶷N�d��:u���PGCCM��#I��1�1��1�c$d�ec<1�3M�4�Fie��,fX�0��$��X�<Q#�Ό�N:��q�\m���U7*��Ȇ AN�C~����q Ԇ���@�����Y̦�����XV��c$X(q���ٮ��)�ʐ�}��L'��8���Ԅ��@���5 t���gV,3%8���b�	1 (�#��-HUjJ����&���*$��$<� �V.0��;Hx�FAg�\��JU����D⿍�s5Y9�^f]�fn���[y����f���wu�f^�f���u���{��x��4єi���K�:Ì8ˏ�]r�J��z����qD�9��tΰ����w�>�ȏ��(����ޙ4�fS?�3	6ɮ;�F�|z~*�::�s�<���q�o��т'�Q:aR2z5h�(���Ii)�Җ����׼�}�èw<�N����:`�B��:g",�(��(��Fa������<;>(wUEx#檬Dp����S�P;7y����[�����~�!�{��`��~�6�q���u�.�S��vaO��f�����⭥K:��a��^��� ���q����`�>���%W�f��a�J�b���y�,��G�Zr$�V��J[X1�4��̴�矚i���K�&a�4�!(�˚B0�j�D���o�ѦL�"�
�V��گ�|j�
G��4UM���~�Z>4Y�YWRҏ]6�5��vS�/���ګP����+��.��	���-9ew�h0��12M�kQ-N��,M@�
Y� o�B��-��"6���/K�}�r�çȋn�V^g�6��)�)��Ϫ��x=fL̾���D��4ri�}��&[���J$���\|B2=GE�����h��З:g�x�\�m/O�>1�Y��sy�1����$E� �Ǐ0��i��4fX��<0��ó�:�������~���8Qc��F�~�0O�E��?�Fh��"��}G�HB�(�$!�!1޸�!�,���TW\?��2��C�k��x� ��>ffgzPӝo9m��O�
p_.��t�U���$#�8²��b}��%#��d��T��-����
)��˰����u���W|\�h��[�|0��bd��e�t�K��B"�9����(�φ|i��4fX��0��Y��/�B%$��e0Jj;���m��v%�|���ø�Q)��0��"����â�Q?~��?s����;<�9�֔���31s��ͳ�d:Jw���h�ó~+嵻����R�;�3ݫ�|7���!>�"m,<w�s2�}�꒟S)M)6�4�0��m�?i���0��X�H�0酚w�K�����byItS9q��w�R�$����-m��~�M7\��S�FY{�À��U<�S�a{1�tƺ�̷7u�Ʈ۳9?;4D�xR߶ղ��Z�0�b�ah�>�l��oԑ�N5]|���-�7K�]�0�|��|���S����KGy��8m�|�~��"Te�ki�G̶��[<2�|i�3,e�d���Y�y���b�['�RX䂤hry�*y����T�j�b�E��<Q����V�����Ee�v�d�2H�M��y���۴S jѳ����n�5�XB��� 8B�3@�&e�X�(�m�mz�(�/���������>8|�}�1�nWK�����0�������J�"��������~?"�	aL�b5'��Tۈ��������~��|�%#KZ!�[f�Ͼ����Db���<��B疭��0�^
cʯ�������[	��5T��4.x��o�����G1piE1��0��X�H�0��>�ԒK�G��y��9�g�^=&�"M�""���r�K�&��H��T��Zc5�m���<����'H,�� tQ;+�"���{��[r�ǫ�[W�#]�
�l̻kY�+�u˗6�;�籬>�I�����_a������u��<;;)O�B��f�N������>)mSNrp��tQ�4�����2�2FI�L,��V"zi�Nv��뻛N�zx%�0�D��O�j�=:0���6t~/�p�`�:=�����~^�G--�P�!��鄖��^�l�z�3z��'�=�rT��V����'o��F:|�s/Iw_��7LJ[�y�I�������ʓɳ�]2}^��Vk����i��q���Z3,e�d���Y�1v` R$�|��Ʌ;�?O=\��b&��>U�0�{�m�>�r�nfQ��c>[}SVHR����R���+'s�>F����C���mC��:0F	��p�&'�qxQc5��^��DW��_̦R�az[BR�}�'Br�ͥ�,��a���U�[�v��N#��FV���� e�0���2�<1�3`�0fIC<x��2Ftb:YӤ`���HΒ1��g�2ã0c:1�3c0e���,��,g��1���1�1�3�@�0`�!�gF1��X�GO�:�udt��2�#&��!1@� c$c�3`2D0`�!���3�L�����L�M4f�Xi��`�(e���i`����Db�tc(c,C<3<3I��KUܒ&����Y�#�ڮ��Vl��d�L�g�,�Z58�fXx;-���p��ۣJ�\��!��}l��"|���k͘�:�d��ՅP[��,7&�^qsjM����&�>^��iTc��=k<�&Y�q?Y��Y�r��G��Z��7yr��&�W�0W_�� �,���G���٤��V�-���ꌂD�D5T��B���U�6�\uۘ�Ne��3g�6xi�&���5�{�=W\���JKHԖ����-F��M�oZ�]s�E��+�%l��r��`��]e�-q�Ĺ�]�t�U��&/{Lm��\sr9F����îv��m��,ЭGKL�\Y��!�a��qV3p[���n��
k�-�b���6fYv�k��ZY�z�*	����˧[���m�߿zn���[���������www������ww~��A��(�M��h�4��1�2L:ag���� ˵v.	tsnc�ڔ���m���\�EV9�JXۛ�[uֶ].�B1us��¹���]f�Mt�%΋6�b��GM�X���Yv*����k	�@Ы�ԁ�%51˴J�]fbKp���bYa�x��/���x2�,�;��&!)5�L�hUD���R��j[�5(jٍ��$�T��I��<��IH�ml#K�Zr߿ �������7�� _|ݫ}^;Ĭ�q��0�o��g�2	��[�y���Ѻ�q���r�7]D������a��<�7ϑIN�Ftt&�`������8���â�ã������<E�&��\(���Y0�O	̞3�"=����L'gʌ2`���?m��s#(����Z�ҿ~��1N��mʑ��SM�Vmm�Ӎ�i�1�X��&0�E�ƥV"'������>;0N�j��	gxX�V!�i�q���#	���U�	1
��Jt"~)�����������$�JYم7�Q�i��)e�*g���Lz�;۽�قl����:����2ŝ�`���(���e�Ej���(��(��Ŗie�i��1�Y��d��q��*zI$���v����3�9��gG!��U�a��[o�t�gEaن�p���շ���fk��h�޵�j���H�.<8l<��:(���\>2R��M8x~��]Xz�̢b�pD�|�m�gƜ)��^�N��a�0矛f�G_f���j�4��:��y�Z1�Y��d���Y1��B���\]���T椒\B:iC(�d$����=ͣ	�PD���1Q���c�Mdm��9��hB����A/}������/����W�y���"��?r��z��,%$W1�S�򷗾yUu�/�\����pc��h�ŞD��g��G����9�-��Q�駫)M|���tn}�cv�Sӳ��"���ahD{�$��u��>=H�4ԒO
(�
4����h�if�1��Quub�湤��u���$��2�w����c��ı���蘋3��e�����x;m1����KK�&�lSK������xb�s� ��Ƕ��51cr7CR'
�wε0��~U7nI1�E+��]�U[۪<�m�v�qmj,��+��z���}>��C���<�[[ѷù0F�LV��"Ty"e���na�J�U�Xy��J��h�p�+���>�)��9�}(��f�x���hgB�{a�	*ղ���S��ͦ&���OgޞCOR0��i[Fߖ�$�m<��>tf����X�H�0^���:���j��*�FOK������9�G0�9�2y��m��#��ˋZ.�9����ɶQ��׼��{u����e��j�')��IY(�й�ľ=��h<�H��pq7x���a�Ja�C�F�)���ٍ={űlz�>D��>�����#�	rMa���Ǟq��~y��1�Y��2FI�X��$#>UX��`�2\�����N�TGo�<��3[a���<��0��Q��ON�SD�9���ȳL�c�qÇ���s��oK	Yku�O��[�:�n�8�Mj�F	`����q��ɭ���o�0�y~~*x	���ɻ<���;ZU�lJ�wS��1��,�[(�{��W9%��%x������/��~����8D6�׫T�8���ic><3F3K4�FH�0;�xn�oʫ<=�����𝉡d������m�3.Z���˙�n�����8������w.��[��{���,��G�ڿI����!{���ԈI�XOH�V������t����Zu��'��C����p��NfFt�$��4��i�1�Y��2OT]]X���'T$�ƙ�r���ԣ�v��_D���[/�z��@����=4n���^kec���yA�D��!V��\6��| Y�4�x���v<m�2
/�ن='1�|h�9�Y�-MdOǑ�q�fA'{:<�f�mn�����y�����ҳv�u�m�����7�:6hS�þ�ij�3�����ibx`�"rti�����A:���\H�m6����WNe-�G���ɪג���̾�D�r���W�?!�"�����R�nrVƋluuu�q��%:����{�>a�a���4�M<3F3K4�FH�02��$�
u$���\JFt�f��`�éfr�=8Q2�L৐� ̧}�}t��{=N	�d0��Y���"vy01
�W��l-�ݒ����ܗ�>T����6¼��*�����|�B�L�y9>�����l�'b'�rw�j�VC4�?r�_�j��t�.�E����8�����un�$c:@��(E�f��37-�[mn����/�e�ӡ�F��H�2�xc,f����X�c<xe�b�c<Q�(r��1�X�H� d�C�&@�3�0c,c,gD0`�GVDt��O2�#'�<�y(�d�c�`�$0`�!���`��<1��O3M4�0�Dx��3
�,e�0��Y�(��CΌe����5z�N\|�g�1�]\�e72�#��)��gS� �6x1�O-��\�s�H�Q�C.��+v��������Z����{������������ݭۻ���J �Ɩi��i�1�Y��2FI�_B�ʫ>��ɇ��a�n����DOK2f��,�3��N��,�D߷iO��M��S)sn�WU��Q�r�0��ֳ�Sӑh����H�~m��-Y��w�N�y����.Å8z���*�%8�i�a��]�M�����a�ܗ��l%Wv�������m�uҌ0f�|2��4�ƌ��a��*�D�O,�8~���{'OȦ��矌�^��S�����8��Z�.n]$���Z�q?a�2���%b���~��,�r&�|40���NM0N�܃N��n��fq#oMc���<z�ز#��Zw�x�#o�-�oi4�,�o>]2�L4��Ӯ?:��Vh�Y��4d��(��FX�]G���'�Y==]uZ$��i��=�+��,f
�{���پ_=ʻܐ���v�lx�yTUl����^4&`��isn� ����Fig� !	��JOXБ�Ġ.[.�&�30�/�loEz�Bf ��s$~�k�P�'&�0���)`�]n����v����ts!�}:00�Wߗ换�1U�j��%I'Ya�a��(��C���i�iQ���::��*�SFڭ0��wT��I�>�J5U;���iINN�yD��]M�76ݙ�)�ER���X�!�������O[�<��|�1�i��#$�
0|�5$��"d���J!d�'�,D����R'�fO'�a�~�-���4��S�h����u�IU��`,^_�%�x�ŢTSH��<��	1��E���#�|A�1�Oլ��񈰙X����z�T��u�O��	�iхǂ�س�P�><т�N�	�P��'�g����7j�Y��n֦��a����d2z�E�%�W:�[F�@�X��%1�a�I�VҞ�7N0�Ϛm�ZY�,ь�M<h�&Q��|�K�s�����l)��\ON�av,��%aS���1	5��~���R �hY�����8S7[|;<�{4�C ��~ȥ�$�%�s�Q�%!|ޱZ4�e:�Tӗ')��G�W����jH��^6K��YTD�W���[���|�34�ƌ��a��"U�jJ$#������O��}�5L���t��a`a���2�J'ѧZs6�f1F�_(�;rGdU�W��E�kz��0���y�57���˚�����0~�V�~e���ȉ$������b~Kl�v��gS�OTQ���PP"����ɿ_.(P�HI�W,�%��
$e|Q�φi�,јY��4�FI�g&2� ������=���82��ě��$���G�E���q
.bx֊*8ۘm��-l�*�Z��Mf�+�8�]6)5��} !.��c\
�Q����,��V��BWD2�=��P�J�0˲�SA|y*63븛~�����q�љ��X`"8=��p�F�b�ǗX4�r;r�W��)�;��ut�~G1a�I�~�s��K�W2$Yψ>���/BrH�U�4��**@������m��3.��O��Ӈ�4�"����6��[����<㯞u��<��0�8ӌ�ҽrI$%m�F��<���ӄ��pLFd<��M5��9��1/φ�ԡK<��,A\����_O/�Yd)�NV��ۥ���[�Teej�V�!�|�,�=]C�}����b0D~>���ԥ�S!�!��m��\�M�s�p��aҌ4њ`�4fi��5�XqƜu�^�Uu��&�W���Vn0�,�Yۤ�,ן����_���u͍���,�xoyj:�3�����^��n�^�%-H�����9���A��l0K��tӿ�6�vu<��0�L�E`��t�:]<�Y���,��|dў��hw�,���⟩�U���~~y�_<돞y��a�q��xJq�Z��6�Q铴����~�z�#}�j4���ƶg�B�XL�O��'��}Kj��v����S,V+Uk9�����'�y��0�;L)��!g�G����PN�3����ЕW�,^�izjld`l�;_qΒ`��Ub�"�				J}oC�=(��&���#�u{�b9�4э(�{D( �2����Œ�&�d�$:H,��;��
؄A)�T
�% �J�!�]!%!BHEBR�BUB�	HEB��T%!R�Q	P�D �0A� �� �D�P`�`�1A`$BT!	HD%!R��%!J�B!*�J�D"�D%B!JB!*0@A �@b�RB�"	HD"����%B!�!*BR��!	UJ�BR�T"�%B ���A`��bAb2 �ADF"D"#��DJD!)�BA��DdDF!����D�0A`��D��� ���"0D����""	"Dd" ��������� �DF"	FDH��""2"D�H�H�A""	# �A#@FD@DH�" ��`��0DF!H�H�JD�����Db�2#"#""# �F��0AB ���A� ȐDH�DH����A"#DD�H��(�EDE%"�!��q� ��dA��1#dH �"1F"Ȉ�A�#D@H"1DFDA"�D���$F�AdD��A" �"A�$DF�0D���H0D��DD�#d�A"0DD�#" ��T�p�H�A"2"�!	�F�`""	��dD��DA"D`�dD�ȂD`���DA"DdD ��H �D`��A�@F�0DF�H � �#A"$����1 �"""DD`�D`� Č`���A�� ���"#D�AF1DF	#`�b""0B1DFAF�""$$`���DA"A�""1F�0" �`�"#""0DFDDdB�%� �D`�#"�H�#dDD�ȐH�`�� �# �2""#D`""#���"""A Ȉ�����2$� Ȉ�DFD�DDb""0DFDD�#H�#""0DF	DA�Ȉ"#D*I`�#DH����"$F����H���F�"2"Db" ��DDF� �#DdF""�H0DD`�����DDDF#DB2"�#F"DdH �D��D�2"�� �0DD�Ȉ#A#*IA#H����"��H����1�$F"C��
 �#" ���0D��dDD��#"A`�I`�ĂDdDD���� �FH$0�@�N�*bJ��fb��%�B �"	!a� �P�
���Y%!)	HD%!pY	P�B��JB ���JB ���"	P�.���A)
�
�*�J�BRBT
��BR��"��Y�V*��D��%%.(��!)BT!	H(�X�"� � �D2F�*AF" ȂF �� �0ABr�A"�"�$"��B*���B!*�A@��A)
���!
�%!%!�JB��EBRBR��J�B���D%T"	U��*!J�D%!�J�!)D� �2 �1A�g7F�d�BT"	HD"�����!B!��B!*�JB�%B!J�!R�"��%!JB!P��AJA��B�B�%T ��!�
�BUB�B!	HD	UBUB*�P��!*) �DH��T%B��D!	HD% F�bY(0AA!J�D��%B ��B� �%!J�@�B �BR�B�B!JB!	HBP�P��J�BP��!	HEB�!!	P�!	HEBR
�%T"P�� DAB0A��0A�%!�%B�BA"D ȅ����B*	HD"���J�!J�B)B!)B)�!)B���%T"�BT!�JB!��B!)�BR)��!�"�)!Q	HD��% �J@�%!*�)A)
�D% ��!P�R�"
��$�
 ��T"���D"P�*R�BT��� ��! ��BJ@�"���B	HE@�� ��BR���"	HD�J�	PB�B��b �1g6S�T����!�Ȁ�"�b "�PD"�JB!)	D%!%B��P�%T"A`�!$A�A�!!J�T*T!��!	HB��%T*!��BR	U��%�PŖJ�!)�!)A�D �2 �1da��2 �2 �"�"� Ȃ �%T"BR��*R��!	HEBRP���B2 �DAD �A� � ȂDH�"A��$A�b� �b	b � �A�B1`� �D�0A�A�J��JB!Q	PD%AA	JyQD�OA�f��Nlu2kp��:4�)�P�����9�
$b
*����	 ��a�5�&߾�a���ݧ���6�����' �����q?��������r��s	M�v�l�JR@�?�g$�I���]ָ$���j��"�Ɗ�����?���җo��E4v�S^T|�z~�W���y�D��L��b���5�H�"��ۊ<��.��琇�$0֌J�e�A>c`�+�8:���/zCk�S���AQ������}�A�����
@xc�([����1@�$�l��L��z�RR}I��n��4�[�rsC(����<·>~kz]�hB1�'Q�Q#s�CT�Ѵ� R#qE�X(E���A�"��P�PB�@���#-$�SNP�S`�����W����`�:�@Z�"H����B�R`�@AZ�TP(+ B��  ����LC���A���+��0���=.8������.j;P/��3/{�����z˦/q�DQEN��f-�����p~�q}H�z��1 �}+�jV��/^h�t1���F t�2jO�'�L�H���Hpx���[��i�yLO3�z�Ew!�b35�t��CQ^Ns������}� �N|��q����������(�Ӝ}`1^p�n���Je��Ca� F��pJ6$�`E�D�����HȐ$&�X�S��`襝 ��$%����a[�;�	a�+�^6IK�JB��pP�����$F�.,/����&2_!=Ò���`|dd�Ok�!9qWdEo!z��ow"�m@�C�=���A>�npm�#`@�M�&�CԜ�x����$���K$;���x�;Q�nQ�P��S�v�;��{Er�)�yf|�03J����;S{�h:����d�� �eCNB0 @��z2�� �I�
�f;G��)�`�E.H��R����Hہݝ�Y�}��:ļl��m5gИ���(����0n��TNa�nh���.J��a�9��5�9&�r�(tD����F��6GC�wJ�5��	D������%�ގ&T �O#�b8���f" ��%�Ph{�K�ц��s�9�.�ǰ��$a�J
Q��b�������.�p�!^��r