BZh91AY&SYX�I��߀`q���"� ����bB��    �)cUKfl4l�F�ֲ
�TZ[c1C%
m���e*�4��k%��)-E��
�TٶB�M�(���Mz�ٵ��n�AK��5i�m���kV6Ԇ��֭��E����V���J���Rm��j�6���V�(��-m�֦�*٣J��t<󖶌�V6,�U�
�Zڶ4�jY��e��Z�b6dE�X��ee����˪��5��6�@Zͱ�d�Y�i�3ljZ�e�ՖC[Tُ=×�5��,��  ;�o�Ыb����mQ�@z�JS�@�ݕO]��C����c=�q�J=�];�5�W�<-oz�tR�eҒtԴ�i��wk26lfF�� ���*R�M)X᎔�S�x{ҥK�:ӽ��=�ʕU7��ER��Ŏ�+�U����U*��+���R�����U�Oa��wvה�*�}���Y�j�mXZ�ZZf����  s�|�ARG�ԉ*�.�k٥J�wbr�kMM����R��m���<�Xt�ԫ�^�(�Z��{���ӏtC��q�]+J�JΦ�UU:ʗ����f�6+T����j�7�  �H5�8�:�*��ױu��O��)��sҡC���_w�R�J����J�������ﾯ��ږ}�=RU)U'���UR�+m����U$+�/�wakV�4ِ6KZf��+f��   �{��J�}�y�R�Z���|��HJ���G�>��W��]�ӆ]*��Wb�$*w��=J��lӽz�z�R��Q���{���j�W���
R�S��΃�6m�Vmh�R�U�m�   �������+�����K�%*3ϟ{�
��5[��y�T�����R[j�4�{�}�^����>�Ǟ��R��^��V�ZUJ���U�N�1�JU{j_{�McP� �i�f[Zڵ��  ���m�6iS�r��!��������2��`�����m�G�-׶�K�T�{�T�Gzuv���Uǽ�z�%Cr����Giu�t^�M���LPE��1�#4	�  ���n�};xw�PQ�q=�@t�������.�p�N��thWE�cq���=׵�����������\��liޗm��ɂ��UHj��  \��Z���WzP �Q�
 {׃�5����(�޼p��Á�-g=�w�H=<y��(��t �^ɪX��T�$مUZ>  c�P�  �uW��*�󋞊:h����ގ�G����=����ִz�{��������о      S eJU F  A�0���*P�&�b``E?&&�%ST      T�U%       �?LUR�3P@    !%H�	��L�)7��46�M6��z�b������у��~P�⊯������~��cʼ���;<�p�3��s� �� {�����{� }�T� _�T U�Á?��/���qV��TN ~X>T�P��+��?/��=�d���Y͑��cف�d���ek x���>2>2��__� ���e|_�_�@���d�������G�G�@��|p�0���<`V`<`P<d_vD� C���م �W�T�_Ef_PU|eU� �a� � ���_ |aU�W� �@�W�_|dy�@�@� � �W� �_~YQ|eVd � � �P�W�DC�UC�AC�Q_�|`OQC�E�@�2"20 �2�2��0��2�2�0�"	�(��E	����P��">2 �2�0��2*�2>0� '��3">0 �0 �2 �0�0�0�2"�2��(xx�"s ��!�x�2���'���L�����L��L!����2��� x�2��x��x�2���x��0'���+�
��'���#���0�0{�>��!�ϳ�#�#��������/�/��/��~>C�������}���>�"k�3�'`�fG�����@a�`t�(�����_�{�)�E�&�bC�wq��dΝfi�OFŻ�\��v^���H'O�wV��ƭҧ��Y����Sz�YNFEh�U��l����Y�K�|���<+8^3��9F�)]O5ō�#���,��Ģ���J�����e7��׆٩�DWV�M0,y�]���1��^!�B�OU,^��㠻�oqB�X�9���]C	��]Y�h���³��L���5ߟN9��x��3N�1�3f���zZE�P7wv1;��+O.��-�jEG��sʄ3X��2<zU�bR\z��B�Y&n�ۄu��=ȝ�	m���V���!f�Y��G;s�y�I퉮��(�'؈��"
n�G69($�,ۣ��Z��N��Yݹ��%�@B��gG˫;�9GA7�f;��'�vs��Uxɥu%���E���7X{�5�i�<�mYB�ʺ6����V��"��	�;l�1�	���f�'%RA���jq�Q�ʮ��\^2�	��X�5m#�=��M&��5,Ӧ�sV�N
���!�!��B���7S���p��56�u�]�yHYA��EY�V�М�����ߍf�����NՊ���^���m��|���[��:������9�+�=�������o��
������C!���.��t�ݡY��X�ho�z��hٻ�S�
ɯ�nC;X"!I�ߠ2�Ʋ�����ɜ�KJ�T�:���8�J���D�Ĳ�ŦHv<��l���,t���^j�{jͅ<�@iW���.jI��^�E����8f��a:� ,��1��s=��#�'�@;-�
�g{�Ҏhv�V:Pm�,S@�`����um�q��%���z��O�5k��j%�n
�e��M��[�鸢��`�[�FB��C��l�<w�gu^�����P��qa��JU�AԨ��F^Gb��J�iD%ޠ`�x��Fl�5�FV�;Þ�g0�T��V�]F��X��Ϲ��p�~8�Eۂ�0�e�n�a�&�4yG����8
:��|�8�fgK;��0d<�p2v\�wAIA^��Gs�֩�4�u�K/�v�Ni���	�z��p�����ΐ�LS�.�qD֙T�Q�s��;E�PT[yhʎ]`��ѩ�@:j� &!+3�w���򱛊�YУ�D��Ywj+��c���	�ϵ�D}�
�g�8(8��G��[��N=^*n���ħ��C�m:f	����jH��@;�l���B+��a�Y� (%�
�^�n�D��b���,�B�am3� �N��jєo9*f\�x��*�E��p�2�Ѧj֪<���>�E�CNR���C`2��-�N�v;(aʼ�˚�hQD�{�ۙ;�H�T�8:*�
��6Sڵ*��ܱk2��ka�!`���),��HQ�*�M:9y��0�}��;�y@�OV��\=R䢤	-Y~�@��s���1�{[dŢ��T�2�1
�kw��6�u�68��!&�N�n����<�t`�M���5�gZ�0���tB5��{%��]na�9���e���+4;9b��Pbö6[��(r:�jS�;;"���jx�<2q!��a���t���+�vB-xl!*8�)V��`�5⻆NX�Oaj_,�&<[bN��l���^��e��I�^I�YG3
Kn�u��V\�z� U�B���(Lm�ܛ���FM�x���ֹ�°��n;G7���,��/�W0�9�]r�:FTFc5cs@Ë6��mlD�w��|5!�S'�5�oӴu���(�[;��	�Жo�0�a�&��&fK�ޒ*��v�=����ѻ�J����Q%U�,�QvB���n���s���:Ƭ��9ƺ�����XCKR��\��
��i���R�QXP�Cl83����tͱ�Pe�!�FɰVN�'C���v�x#�zl� h,є#		��b���$�g� �Ci��V�,�IyX��t���ݨ�">�髵d�G`�d�t٩=B�zR,�h����`��Dz��R��Si�3^��8)�2�ہp=��2�K�;{YjV�q`	7����Z�Eݏ�^��.�iٕ7�{���g+A�����3��X{9�I���Y�
f�<z��`J��������x�=�2�}t�rw0��iw�2crlf�N�X1��ܬ�j�A2�BUÙ�D�����lӂ��5��ńn�%� ӈ1�n7�h51��¥iXJ���w��5�5�U��K�si�cq��-4����(��YE���	���4uUt6ƕX�Pq[�n����Hٛ��F+����L+���Xz^Q`93t�[�Pd�<;��r8�ec�|��J�l�"-�zNu��=䠂���hKͻ�����Γ�W���G	�T6���[r01����{��6�QqP_���K��@�j�<��&��K�Ŝ�yS#M���8��RAAh��v�a#L�G����bi�K7$,m��t��W���z�{pC�Bޏs��qL\�]���,��Ȗ-�ZyܺY᪵�ћCN�^�Ch�:J�`����<�rٌ��caK��9�O\�H��z]�Z���ȑ�pƦ��x4Ӎ>ȵ(��ї� ��<݃H�p����p��q	
A�c�Ź-'�����
ŵ��j��R���
9p������S�:�Y�`��E�H���@p������ �O��}��˴���[d��e�8�@�h���(�Zp���B�}��^7q�o�4)���kt�v�"��%%b�S4�rF1֕�25Z� r�ʚ�����"�\���Y�Iݣ2�(��+6�C&P�U1��b*����kכ��_��4-�5L\�������s/�����2����.w]&��l��^�P'	��o���vX�+�:�#�6Z��F�g�Ӣu�ԙ$y�0ڒұ�R��Xi���a�b��͜�����Z����^fiL�GmC	�[PY�^���y��Ņ��5=���$���vC<�xv�,�ʙ����5߬��)��}$Ĳ�i� Z �mgwl�ҧ��d�Wg2ΞJ.jb�ղA��c�>su0�Z�"Ѷl�;N��v��n��m�t�N̊�Ri���$:8)�!����&P�����m�6m�GLm)J�9B���>�;s�{��Rt�e��H�+�#��-ܛ5�Sf��sr�gU]�b�rM�����`�XwgKVv빻��(��=��M�oK�Z7w����rqգ�����}t���q��g��5��wR�w#�$��zŽ̜e�Mv�)���^�j`�Gd.�*�2����/(-Fe`5I<�#��k\>=�8&�N�N�D���-ײ:�m`���H{�At3f^��TI��L�9�����G^��v�rˣ�p`%�m�6l���ť/*��	ݦ�{��tmhv;�8��K��KM��N���ceį$��Q��];.�\��ffU�zJ�wu��*sE���z�8���f���CV�����x\�z�ef�4�A�kmww.I��`��c�n3	�rD���o&��.vPC����U���Z�W�װ+������re�t5�fƵ���K���7�8Fu�3ztC�Ƭ���;E�g��Q�LǬ]y����b��kb�?U}�ʻ`8_ �'���&oe�z8x5̓��Q��0��W��F(`�{�5qb�� �3&I��3
7�0��"��W9���M(s��Εڶ��0�"�n���$�罋s�0�;)�/��к1#�E�=i��~�ȲfׇdC��X�ɢLv�p�]dH��,	 ��F���+ �7n��V�|���qu����&-r���c���5E"�����L�%m<�Of���E�Ap��'h@ӢTMUHT��8j�T�G�-I7X�� ��FWAC���ַE�R.-+��λ�2�K�y�����n\��!�66�q[ш/	P5�V����$Մ�׌lr$�"
e߁C�Vwۧ-l�ڲ.�s�;Nu+��F�2�Y�D�2	v��L�ҭ�Xhh��L2���n��3��9�識Pz>�:��xz>��0�d��!g��Rp;ێ^��Â\�Z�F��)�gt\X�pF�T���kb�@�C`C�u� �����,�E�owo`A.�0�N��i�)]�Z��n�[��Gr������h�90S�#�8��Ε�]Wwj�]�*�y��:�V���ג�&[�4d6Q7�2�7�'a��^�$�qh�����r� r��4�f#�rw�3h7i'm�ZS�T|�oR��;��Pȁ����hs��F��)g����v�ڸ�<_od�˜ɚI<�+��	��}v���$��t���Ra;�G^x6O��(��ϷP�G3v>%��r�n�qPxn�h
;�K�A��4�a�I���=�CǧS�΢pk��3Z����G=�q�&���ΡA�8L!A��o��T@l���ql��d�Xz�}��,U���3S�����%lP�֠���u#���#��׆�фƪ�I�9���p�z)r]З�Ʌ����M��oq#�#���6�X���R��P
H����g3�#�9�Ys�"^�����$�%Gu���!���+�2-5AWv�rK��6W��b}{�'7WD�2p'��^�Rԯt2I��I
*n06����QōCV,{5��e}��F�׃���5Lw�:�ƃ���D"5�����U[�+η^��`���ZG���Y�;�ʛ#��)��O&�����h�J^��aF�j�Ƿ/]����8���3��lY��B��%�0%�!�l�`��=B����zeSH�g ����A������AfG��5�+ɡ�$ni�X�j6���[�n�NJzɴ ۍ��[>��x�LBV�@X���w+fD��P[{o`q"+e��ԩ�Rf��D6��(+W*Q��(֍SϚ��=�����|�ܧ|�kq
�!��)`W&j�K�3XCsf���&6Ӳ�ܨqd���Ekv����3/dt(fQ����-t%�5�,�T��\ �a��&��S���B���xFiJ����m���vm�y�|]�,��߫H�6��,�����-]���*�K��ڰn�#�a�C����ۧh�)���/=�z�.6�X�v;x��D��^ �K�W�+�8�q�Lai*�>���t��q25���*�<��ʙ����Y]���h���ej�f�e*�oB��I�� \�m_nS���F�)+���ܩsMGR�\u7�gŇէ��n��+3�⋔���f�Ot�,핢h�,+%�=e�5|X�󢴵֩n�ɮ�o7V�gJ���1���V%+"��5��!ħ��r3����˺���8�C�Q=�h����jlכ�\|5�V�Z�1��7Ned¶���-��5���6�KBSȍN�N���=�Yu��ǈ˚^9�&Pn��P�hj�]-��%�	�鼦��[���V�z�%�t_W��y����nv�eJ���s*L�Y�̷(*G)R���c��L�ܥCE�{yZp���T�LӑF��,�l�Ƴ��L��S��[������oE1d��I�A9���ݳ�Lg���	�&��sD�z��ϧ��{���Y�W�q&>o��rTś�ʻ*X;Mou�g#'��B(��������(t�Q)�\H��u8�7�_-�c���<o7 y�3��1�%E�N���EGJ{0xkz�b�7�,Е�U�Ҏ�	�2� ��zbŝ��4�����Ɛ������]n^a���Yy�,�q�DZ���b������Y��]�:S��.�՜O'���Q�iR��@��;ClBe���j���YF��+�RCXT�`��hcplι���pkT&�Z2�1e7��0�X��((�f���<�$ߞ��xO>]D��<�wd�ټ�5� h�$Ľ�Uٽ���8%I�s�m&��B6J�7�Q	@�i�׍0�vL��KE�7��E��wZ�٫� ��Zm匥@��V��q�ݮ�9�Б��pf��n\�fh[�hy��oSd���zG�u/v����=�Z�6W){x��1���W�����yIH��⳶ݍ���R��Hn����%;��Տ u�\��:8Q�c�Z	�����RK&�;�$_�NќJ��9�Iy���H}�]�uŵ�+�v��0U=|�w�a��a��M��lj��/haצ��}�T]��*��FE�=׻)��,�cȪTT�4q��'�؎��X�6.��Ӈ���:*��V��b�a:�}@f�����m7�g��4�.ǎ�P�ssu�����G���Է#�6�nS�M�3�-u�P��h�xp��p�e7j/�ե+��LY�t�ehcpA���;g=�kK8%]�=��K%1�x��t����3�o��#Qoҳ��7�ͯ��#+�u��93K��dd70na�D͵��� J�bE�����c:v�^,�N��4j19�7�sF{��ō�ƙհXJ8�AX����h2\�wيlq���1Mнx9��|ș0��_5���}I�" ���,�A�Ga��7㉷}��e�`�c�f���+,�\��T� n���̅)�w��.�ͼr�2��+�:�)�Z�ge�����;H��� �o��н���<�~� %|3i~̫��Z��k�G�V�i*%O\�X�wY��N��fsMְ2ړf��̸�0圣wū�go&j���cC�+hvɝ��+��R�+�Z�l�f�u�o$��9-�n�;Y����OD��vYXﶊAt�´T�Y��'�P����҉�H���iR��K�*�m�Q!��uL�V�����e���5�!
�rk��W����]t9����8 D���;��t\�O�{���a1�{�]���x�9�Q�k
6����ő��y`WR�z�����`w��8B�5|�zw��0p]��{\>�f��T=Ț�x�Dr��9>�t�NdX�t�[��&�sNv�;I�����T��
��9�,1�!g)�. �?�_eថ�{:�5�$���6�q�Ջ	�NyӋ��yh�3ˬ,�
�]lY��"�Û
��[�7��LG��7��BW���}ۥϐ�2�)�1��@�e��X��4ݹ{p��w݈��d��9rQ!gi��5��bFU�ٷW��:�zZk�����Îj�Xƾ�i�L�d��4�]hn���# v��e陸�"��F��Cj�]3Z	��knkӘ7e�L�CK�ޗWi��9���
��f�ݖ��n�KM�mR}Zc�LxUm®���L��,\�O"��'�1X��u[,�!p��2aY�2�
�|�I�;��]02�]�.�3��y���Fخ�%^��42tN\���Vl��qU*{croy��)���IZ|�H> 1��zvE����N8�~}��L�Ԉ;�o�[�/��M�1�����cy�vU����n� 6���:�8�<���bӸ<(�Ck+¯\H�'���t�m��������vF�*���'C�җ�M�;Miv���ບ��E��9O�kr��={��>�p'3��]t�=��^�P����Y���oP�K�c���΁7Evm���r�r����M��vO<�$a��:�n�{O-��v��Tް�VĮ�I�Z9�9�S�K�	���wG{<�g�",Hl ==��P����4?z��w����ʪ�-T��T���y}]ܵ'F�E]gS9c��pѨ��F�&^����\n�[ZU��j���];�T�D�k���ު��Pw��繓���줗 ;:xK�����`�AD����̃��<�&�����1]Y���;�t���
���F�V'��8���ђ�����t�0���彖�;@���&��;M��ӻ�-<׺�c�S��="�ݲ��J�$��hT�����f>ӌ$2��1�vN$ExnK�I�7���4��+����
}�EF��=�).�1 ����7Z�93W@�d�!�au8')I���R�P����Ď'�%B���r�)p-�:�MhghV�7� �z���ss}�������W�k����}|�1]�lBrt��7�:��#o���^-X�ͳ9ŉ�&����s�,G�2[��՘�ҙet/��x5wI���yL|ͳ|P�%n��m�u�Ju���-�ç�%����%G9��3���	�z��P��X�W�ҕp��׭�^�9��#՜xmGR;���6d��!���l_�a�6� ����5j>�O��b��ha`.\DΥ����rmS�����[��:�e�)��#��J����Wg��z�4:�6��9�5�T,����k�ϝN��h�ű���O�m&)���i��R�ql"3�>i�t�`��L��k�@fH+��i�ț�za>��D��
�
ɧ��/S�Y�>��RK>�Kaw�����&<�߇5r�;ޤ���h^X��9�q��ţ|����_oj�����n*�����8�� �9�z($�I���kz��̘��Q��ׇu�t�͡�����yX):)^X�y)��ԖcК�E�	}�'v(�"��ug,�u�$��/����lȽq��]���9�lz�p�wرMuw�o��DJx>���2p�8��`Q�l��T��R����ˊw��M�\n�*�Qn�d5q��c���rĒ�[�Qo�}�`�nu���v..�K�;��L���>����FX[t"|3Z���Z��4��:�ڪw�^:�8�5�wv�!���(c�]'��4�"){��
@j�8��f��+�J̮�taCVN%;ȥ�f������f��܂��2u�X�4t3I�'���#������7ey���6�vr;���l��7*)4�y!�gh�~�=&���7Kjp�je�
[l�wMK��T&�Wm)���OJ�V�rr�����Үi�2�̬K���:�.�\l�,Pon��9�����]u>�� \����Mn�lŲ��cy ;9��5|�������b�a�?>���^��A�7�8oj���=s��Uˤ�|z/dr�\�u���Yͬ��L��un-F��Ѹ/�]�iJ�PfH�|�k^��6�q�����K��^��M�3�M��|7.�!��x7<r��T���ǼgտL��{~9�ޙ�*z��mY��x1G��F'F��&�˙j�R�t�H6^�1G:N�^e��/f*�Ju��^������M��Y.�G��'�ͬ��I�Ȼk��/+��F�޳SN�Z�"c�'�y�.k�<[��k�ڶ,��Ғة��1�E'��}t�zk
�a�=�)��1^�L�n����[�Q�r�Zz8����K��朚��S�j[02e,�<���ْM��&� �)��,^�����{T��y���ɭ+C�"c%/�+��'9b������.靹q`�/b�|��o{o7���&�<�V��2O��[n�4�)A�ά��5�W+�1�C�aʍ��b��D�[�n�w�%)�F�N�*$�d[HĄ]�Lʷ�CÐR]� ���3��8Yp�6cO�s�I[m:��9Y��]t�̜k:Q�n�[\w��K�}�QB+�%Ƌ��.f,!�5k_o}71�eŘ��&A��7��N��#tLv�=�n����Z�ÜU�lr�7&?{�l������m)��ar����kbR���4�\�T� ��~�MU�6�X!M�t�n��Ip�B�WM�l76'.�n��I�v��H�8�j��\���s�2�J�nK|�Z#×+�Y�d��$�uFXYK(����s�&"� �����5�K�0�,s5��c%j�ڇE-��V%|S�����`�N�I���P��y�z�k8V�{���+����5���&�ے����=9������k8)$]� H��v�R*���՝����3C���^�u��9N2���;H��ww��y�͜�u�-��\e������M�����R���j���D��s�Z��ݴ
]�i�M���	���tx���6���|h>��r���cT�=�}���Ӱ�U��85Źr$�1������7<1��?<�eͩ�;s�iSo���`����D�@g�d��6��6Y2q*��a7i�h��F>/��&J�y-J�M-���+����C\�=Pw:���a�6�X�e�P,>+�N��L�Y����	e�lc�]}�<'�`�8�yb�Y��k�6����r�� 놂4��	$}��U��[[�f�����-�g,�6�aXp�4S{`��/�<��&����sz��/�%�`G�kp����(��=�|Z]�`N�-��'3e�]q�I��qj��_���+S�(��	 ֔��"�"��؅J�Ikl
+�6|:M�4��;6��5=����R�hcx؈����Sy�:��a�����û�0���?5�2gsE�nB讻�r��d��
����6�icϑ.ھ3b4�鄫5i��J��ӐL��`���r˓
�]C)on�1�Oٔ�8+h7T�a��WXӋ/^�X���@f�����%O¬����׶��L��P��gv�I��!8�YP�e��^ ��{|��'؁�//7�U^ca�8�PG@�h��d��"M��)�8A� ���Y�zE�Vj훯hNบs�	e��s@�|�B±�w��]dA*5�=��b��6�Hx݅Oʃ��3���GeY�ʣ|+�}^�Z��F�zx�)	��I�W���6�33q*Z�]F<r�e ���s�u��:�ٺ����6�h`���^+�����\����H#+0=����Cv� ��h���K��y�SX�w����9'��8�4	��������zQ�o�p]U5p��E䤬�S�s��X5��9�ۘ��{�|
B�Nڏ�>str�S��IGWrE�v]�Gt{��t�w0�#�h���s"��<���ʘ�ʭR R�l�͐)�WH���w�:�{�ek�^��]SC�ǝ\U�B�Y�v�vC��9�s+5Ld��H�v��Y%#��X[��oI��[���$���q)�$�A�t�2G�Mq\��D�'��8��,�STYƲ=U���ec�	"u�B?K�3@�͈$�p�dLQ[����c�5=��F^�w7~�!~�o���VT,��gߠˈw��(��t0&�n����%�>(�$���o���3-3R�PN�#nf��[��l	a�����15��cI��c,��{���h�E�WϷ��Vd�+e��]�A��	P�AE��u!Xq�(���O���|8r>}0O	��jI���b��]�3۽���C<�OS���.�w[�!��#4.�Ь9��e�t��#��ʗf��j��Ղ�y���V�F8bS�Bu��5�5ڍ��:0�KVM�9�*�I�蒴�:ـm.i�'��Wn�����'w���@^úzVT��s������)&���Y�z֥I-��ץ���}�S�z��)�A���m��l�t��f�]�S����{��Ltշ�@�����^��g,9}=�rs`unP�Zq@{V��`VI��;3��mS�(mA�x���8�M����ֽq��8�,��v�Т�j�SqQ�egI�(�&�W��8;��i�M�
Ŏ�E���]=�^��-Ցj����zOt9b�QX�ט�Z�YYn�ַKv�ӂ���PI��M�詋�kJ��Ɖ�ԋ�}�L�x���1�j��4���G����u�f	�P#�Z�d��h�]e�c>�yy�l;V39f6�kl�Ɓ)��:��v���fW���&r%,Y!N]��Aބa�ܚ�upFf��G#�CV�}��2�o����Z�Nb��uj��/�e��
=��&p��w���1n�������-�ľz���?nI�[�����+�1�&D�-᣸ȋ,ӡE�sSK(�VM���5a�<N_J��nݯ�{2��;5e�9��k��]y��F\�q��i�	X�XD����OnL��� ߷�ǉ�8W̭��]�o���ys<h䦫��;g�m�����v� ��lk����'�2M��a���u>(��u��/��A`r�Ŷ���=G������0�9ǾN�W���Ifӧݪ�����t�HQ�JQ�k6��V���R��{�ZG��q<>�)���_n�=�9��w�,�k��c^t�X�b��Uo	z�B��b$���3!k����{�~:�����p� ��C���b����-izkY�t�Z��Φ��q�\K�n/o�3V���BK2^�7+�u:�R��zN�֖�;��F^Y�6���
�(<[��,��)�W-=q$t�Ke�>�ʾS�O����ה����R�p+]GC���]�A���7.���c)���;�-�#<�#:�l`U��d��&��$��Q���Y��AM����� 4���6%���rrCWa�����ܱ�.��Ȗ)�d��3�W��eQ�}::|JHc��Z�0�\ ��q0�R�	�ؕ��8 ׺G��QQ����5��]�5(";w�o����t��GQ����os5�l�7of-GP%�,C"S�.�ur+/��b$B��bE(�2�ki�رrk.�n����n��0X�7	��h�#�K���4��JX(ӓ�'}��ϱ�VV-dT˴�eIC=�]��t*Ε�����"�fv�ߑ�P0��}��4RoD(+��;���j�儖+����ǈ�����8drl]�p���ֿ���W�Gsb/ke��];�u�0�gJF��Ԋ|2���)�5��Y9wD��cFN:@�(Rۤ��چ���CJ�]0�Ř`�v�"��
t��b�ee��p$�l�5�ok���BBD�C;+�� �����y������E��ז��v0�>���ax̆�T��dm�7
��-R��1u7���c�<�.�2rj������]�yL>j�US�{�Wr�jZ��x��f^U�,N9*ӛa%�;�����d�Mz��v��y�;ϡ�>��J��}+m��}�`8�bO�K��{�*���&��O*;�<���xV�Ihm2;:��+X~�<��7]è{V:yԞ��t�.���0븙�:���.�@Ҙ�b��Jt��]�o��#$j��ƨ/+s$˫^lp��;X�q5IT Vi�S��wt�v^��۟b�M�ͻ��i<Xe��,�8��&�W�W��<{�H�5������Z�-���m7��ŧr.�!ǁ�G�]`��,��ŭ�Y�*^��a٭fJ{̸kAC1EBb�Ύy�je�ٲ����/������=Im��Vuռ�nӝ�F�%
h�4Qh4�!p�E�HT&��Ut!-Ӥ�- U
(q�C�͇" ����I@�&A��
!@m�LS-���0 ��A�h�,R�i:��D 0T�,�E2[4i�Y+n��(���`���	m7A�{"A@5D�4�"[�X��L&���λ�$&�RH"�F�]�+�$QE�������A@>��������>
*(������|�g��ߗ��^���~7���|�
ʷ����"��=�WMu��6��������<�xMy�)0b9�
?m��փڥ3j=x.�B�lԣ}R�x���펌e��{2��GUw�i�rK�R帲(�eC�^�q�rnR�m�6w�C�δ�"�t�'P�?-9�8L�Y�y���^���}F�;���/�� B{ϓڷX$�J���-j}8v�m�t�m�
p[�eWT���ԜQ$�{\�f�Y�|W�P�^)3$+��f���V�h�7P��eK�u�5 C8�E.ZM�X꼣a=��U�Y:ne�8��N�ӗ!��	u��V�e�u�3��]���d	�iԣ9�r��,M���-�f�fJi���}0��<�t�HV=�x$r��O�0݃��W=��¦�\����X�/-̜_�����+`,�s���t�K��f��kV��)���@��)�@+��V4GtR瘋�ɇFl��������}�oVbr�T�����y���h:Ŷ��efp���1�y|���4%��aR'Hmo�"����fᤠ훙�,>�GAo�W��Q":�����q���?�g����� ��@��`���0�EgU���η�4$��h�1=�uj�]���lcj�G7~� ��t�wx$@VPko9B��خ�g���w0��j旋�v�Niњ��2!���u��%�����p��Ѝ�K\�.H*f�R}�a��'����\%�gsX�XMq���n���}:�$hEЬB{��lGw�=�bX��۝���bs_e$�(�&����G&S�k�NZ�ڻ�/�j�M.��N�4o���2!1f#�[��b�w�R�ٟ(�80%�[t��-R;P� ���'}���>}�uq�b��r9(4�uq�J��"\�Zp��N�jm��C%�~�����kjط�H���wU���XMު-�bw���Z�t,�;���,Xxp�se��e����O&r�O�^2�}���y>����yծ��yhה�]�vG���?e͏���Y��W.�
�'*D��3�����Ǖ'+�D���:�I��?_*^/_��F�+-����l�lPo\Z����G#����r}K#����j�8���H"�Ç��u+;�!���ݴs�f�&**Gs:��U���o�����;�+w�8i����8�����1��K�2芌UphNR�����X<-c(�:�/�#�2�VZ��k����G�2Y��������<�,����KR�C��Ƀ�,dS��LD]�#�����������P�ԨD�w��*R��'e�A���{ʕ�*m⼵�FI�%+:y�	����c�!yE���}���x~�.v���c�7���o���q��ZN�?,����uR��[�4���0<\��"Nu��G�2��$U��0�]r]���+#t�`;��)̬�}#�`�W�v�����!���BjT�i�Yԅ�<7�
E�bar����ֺ���#�!زgpQn�����]P��0|�+|��Չ\�����xo�c�����A|��du�n�_u��ŭ�J� �K]����B���U;�I��s7�mq�q�jlM���f���s��ޙ�f�̒�:�kb3j�����'{�}�7"�UY���Y�1�4r[�٘l]���)������:v��i.s��MPu��֍3���<�iJq����?w�Y�,yd�8}#Iy zX�)5�=�#y��sӳ���o�İ�!�Մ���m{#6j���2 {�ڼ}��(�Q��F��3�n[ �:sy))9.l��+\�����w��G]�J�Gr�F�*��|a��0B+Rt%�&���i66�(�j��ޙ�]�h��Y����]�|蚼��{{F;X�Хg�e���cT�q�@�Q�	Uok������s�2�-ct#�Т|=/��L_ѱ?knv{����@A����]����V �iX ���-�l��{��j��\����:���ǲ�t��:˾R�Ǉ1�ό��������wf�����K`ٚR�J^{�z60�t��á�w���]H쉠�9d�+�
�b�^R�0}��Gc�G��^v>��N��
n\X�og�!��Y7���:�s�Vjr� ��D𼓶�.�GO4���n<O�1���M�������7�Ǹu���9 �|�=��|!���E��`I��TK�qT��-;AȌ����Xus�k���,�l���ܐQN����Y����z��]�j��{�K��+�0����.'�5�T�����ŻH~�8'>���U�Ʒ��{��`Y�=\���fJ�YS�E�%r��>F�������c�h�O@A-�l�{�c���>�6���@�V��6�ؼ��y�����וd��8M_Ƞ��`�ݷ2[��J���L�1��Y�i�<{�,�`�\�f�Q������٩��.vc9��.x e�$'7*��f[l{�ۜщ��hj�������ux��'��^�Fx7<d�r��E���c3�x�+:�+1,�4�<�wP�r�_ 2qz�IgV�т����زr�<<��lP8{�8:hQ����F�����{����g�ɾMd=�h��՗�{��ݴo$;��`�7V̢>���o��nYCt�<�m��ڊ�K\���_g"ܐH�;��ZW�:1�q�Y���C;F�3T��:�L�������ۊ������kC���e�V
�Qk����YAv���V2:";��52NJ����{ʧS�6�ַ(�Jl$�l��ݯ�.�(�=Ö�1�[p��Ma��-l���b�P���iU�n�{�e�FWN�W,ϐ5�xs���1��c;�#�� X�y���y��rb�����"ג���H��!=8���۞�G�ý�CheO^��ٯ����J̋��9q�B���-�|t	r��Ȟ�]#!5,��DOt�}�GC�s���݄m,y��*�D�f����*��u5]�`U�s��P���q�v����*�5�B!����r�L��5�"}��4��T�������f��E� �}
�K�o�h=�+&p��m�Mq�0K��΍j�����v�ά<�.sBV�Z�ճP4�<{�c�9�e�e5$����8�R�r��ם{���������]�L8񸧸�NlX�x;�b�9�1�~A<�=�	���U����[���l�['Rè	���[Ѓ[����
=F�@�Qݵ|�������0bt^���ԧ��VOO��cǍ� L�()p��G(���x����s6伧����º�ν�ӌ]� �KB���FP� J��`��L��)F3�+(�C1o5(�������m�j���S�o\Q�J�A�d�g������:�ZM�+x������l=��<>��5=ثxaGw��F:e�����*�,�|��@ȃw�����V����Ub�E'�[�p#�^�b��z�0��u�t���&��ѭ<��Hj �h���U���
լGN�R���A�b6�⮉7�jg-�+%ޮ��UȂ��:fn}�f���གྷ�k�{>��RL�
�P��t����!]$�����5��c��!���޺ |�Q�O�T�S[w@K����YO���W0V>{��՞;��~J�*�0b���OGHL}���hxv�-�3��e�n������Z7:Wvڻ�F%��ce�1L�:�Z/��%]Q�'�}���H�|��V�P����ի{y�:}ʞ*J��`)I�삒�棱Ng�ZA��������$/	�&bn�+��w!��j�*�ț1<��p2�]�A�s�^��}V�u ��ȯ��i2&�X�����EN-�ytq�ݒJ�Nr��R��N�Mygc#��"�}4a7���v?����{�Ή������W�6��}:b�g��]!ע9����CM�s�[�Oh�>ɂ5.��^'K���ɥ|?&4s7d5;'r�7[���]p-+< X�Gν��+�ˇ�uw)2\#u�'����_(f˶��:"kx�["�^�I���K�Cj@�����ܲ{���+M���[i3ϳ2���Wy�܍ٔ��a-��V�u9
_=��aХ�c�w*�������r8��M�����p�ޭ�:/͙�ш"2�fg`��p\3l=!۱ף2���I#7�im�ܮ�z1.��VUxr�i�[�]���e[�^���U&^�5�=����.x�|�YȏHn7aI�=�����y1��3oބ?�*Ż�[��-|H�4�Y[§]�t��*P�-����!�]!؎-k|����R{H��aqu�l�͑�K��V|RZa�$W�1���(j�N��[>���5Շ9Sx�X*�Uh���N�S�N_}>`��'�慡�+Ioe�d[���Mb�-ۗ��K��v�\rò2D����DPV{���|���E��:�t��SU���V�a�uX�q��^��Reo����}<<���ذh�=:�DLY�P�],}��^Cy�J�'Q�/�UK8\b)��2�[��m:�L8���f��\qdh5�0���8�yA����퇩�A�N�v�܃��x%���9�§V[<wҺ�h7A��뾗�sĲ@��5���Z��2�Vs1f���-�fk�ViP�ʺ6�Z�Yɜ4�m�x�F��3q>��z�KG�΃��tc=n`��:Ė	�Ċ��s8�����M�t�����I$�@�բ{پk7�l��Ώo�' ���zd\B)@�h$�M-Rc,'-'e�ؘ�Jd�`qH�N����L=��}/��|�	1��؍��>�x�|����{�\�������,�r���vI)t.�yavGY��cW�mص�Xns��s�L�{��G�i�j\��Ș1b�x�!Ev3��q�r��GkS�X7Ww��)�h,7)�|�Df�ȓm�:�������
���F=��Ъ�D��d��:��l��55\��(@�l��+h捆J����A�*�)�%6:&=Y+/u�V�
v�5�W.�|�t>��	B��o,���S�g��/�+=�*]
�6�h�2g7��r��}0I*p��.�}+�;j3�%��T9Z�75����	6��=�]+�WA��"N�bI���]�+�j�˛�J-��[�y2Gu��G,�ܙ�WV�Q*V`ltb{�i �"�N��i��u�C&J�w�f��--�Yց��/_3���<-X�ӳ��H��*]bچ�<�t��	n=�RbK�=�Yw�l�{$�FM'�x%�[@���0:r�s��Ε�4C����Sr&n#5������C2���SX~���L{�g��r�)#�
v�/G`���uU� ,Dd���rHw�ۜ�l�<1H9j�z�2�m=����w>�t�+��b��lkz�O��Z���5P�E��JZ0g:K����/�F�^��;)ې��2J��W(� 
�T�E���Io�\�_Fn8 �z���A�{�oz$����]���3��&��5�wqU�h7f"��X���]��s1�'��8#/�{` I]��g��G�
�ֵTq��v����t�ȶ�����u�0Bj��1z/xSI(x�Ǆ��1�Y�o�Z�ݡV4s��������L�p��/x�e�=.@RW7�P��S���p�ڌ�V439����n���Wq� Ԉ׺ ��ӭ0�\2��&�	�M#;�)�릮�̢���p
��n1H�`S��8(�X�]�Tk�o(�����b���fݜM[���u/�n�<8�6�d�[�;K|��)�ٖ�/Gb%v�J�k�����l�z�ee��u���t�яyA>�<^�U�\߸y�\оqX��44(;�F�9����4]F��[�U�)gm*����0���.�ᨫ7-�%;��o$�l6@��9��ܾ���_��vnX��@A�ٞ���a}ޕ��5,����B�S���~���ݯ���X&�f���C�ML]yvV�h^��4Qp���VKz4mV���2�0v��q�И��m�عS�U�qiծ�E���
3H�Oi�z�Ӵ��E6I;yi�u��`�k9��:];᎔� R=�V3�֮ �;��꩐I�(�ևX(L4DpI�'��i��Ef�F�x^�:����O �.E	槮��p�;��!Z�N|vì�׍n��}P�˚hd�:�:�XR�+
����#�c���E#{<�c��!A��C}�q��!�����-�Bl�k�WXR��c���fV�*!�в�(P�ʗu��X��_4����zp�{�%s>C�T��pw�����R��Un�Q7$�!�"�W��ž���lg�}Or�%�A��;��ZMQ?a�}���IP2B��v����z�������&C�jn���u��3|=܋��'
VHQ����*cVuT��ҽ���<1;ø1c�]GX:��/��M#{f�+%����S�Qy>r R�FL�B�����}��u,-J=Ѡ�����=gp��\cǧYM��rא�yYeiw��&�S�(�9q�T�d+��,�5�P:ug^�9Gtz5�wφn��b��@��J��U��3ٝa��k��?����"��&��U��(}f��ذ��eBvn�2�ys=���;�j�T��/����Fj�z��@V�ԅZ�i��e�r��X\_3��M���sq�PMYؒ*_?^�l�1����� �<��X��Ko��uZ�VweΛ}����wD�׸�^	^9����z�j�������������@_ʃ���?������/��g�G�W���}>��W�~��?���_lco� ~L`�!3$8��;1ySё�Mi��~H_&�k,��Aj��8����-Zg#�\%.��_Ϲ�)1W1*�p=Y����%Yȭ'Y�٧i��î�@�c{�`�Г�vPӼBT&~)�(Y�o������c�{ݳ�1v�H[uZ��Ň2�oo�2B&���6�y��\rV��8�W���+жFY�5��H�	C��J�c5���MY`%[��C�W���Ǣ�힦9��o�2�Q����x��ݭ	\;�����H�g�bu�q��}s�3VY�W�s�ջ����x
Ռy /DԸ�1}+���Љ����88+a�u��r�*��}`��:�O\఻�$(-پ���Qs�G���9!����̺�YI�f�V�a�n�ĵ�R��Wg�����ݍ�\.4m_�m�e�e�8��R�m����-n����N�i��F5��(��.��B���Yq��Ҁjg`��R��}�͠f��dy��c���q>�(,�W^���w�o�����p�Ɗկ�P=k�N�g8�utN�Mǎӕ��Ljv�)e7s9���N�B m�"�s�A��ǋ�-坨��R0p��Q9Lغ&t�ĵ8&MGkn�����	]8��^�B�=}���<��h��F4W��%M>��`X�Ȥ)�&��A�	MR`��L6C0I@i�{���M�ABR���|�t<�n�����/FՍ!H[)H�Z
M�E�Z)t���4Qv��F ����\Z
4&�ZCM��ŰTAN��Ph4ӈ�h�i�AN�(��œQ]t�RL�CF��	��Y*����%!���]qܴ�a��(+�����h5TDcb�i���'��q���:����F+clh�l=tZ��H�����M�*�d6��V�q��!֚b:펷n���vN�3��ՌDS�-V�vN��F5tPq�ص�Z(����Q�箢
(+����h�i:�ض�OEQM���ӣI�u�:��t[wb8��UF�Q�A��.�
n��ւ����=߁K��؃���~P�6�7�~>^N~�^��u�8̣�5�Vz0��`�ԕq�S�x����E\���V�2�w_(��	��{v}7��g ^0��r̰z�o��t�/{�]z�I͸�i���}'�MU39B��z�p��^7���&�씫��ԅ�{�=�v$����]�OB'7�=K�弧O1Wzt��U��u�/�������I���_��Im�[�Vv��eU6��Rg�3��#�P��Z�����הR)��8l�b�ȥ:��{�L��;ߞ{�-���V��~N��c׼<�&���7�iu��غ�>����-�k���^�uS�9��W�E�������>�j{���Z��C^0y��:��V*~�L���[hV��`V�m����t����s@5o*+�V]'���W���wSt���;.�ԽX&��qe"�+�3�
�mO7�hzey_Z#�&���d5�����xpe�u���3��mn�����I��3�����~���c68��vXE����u��p�i�s+�mo�qev�_�P��ga�<e�\��Gߑ�ƌ�u ���-�oz���d�y�y�Ja����J����+W�X.y݄c'��Y<58o����e1�C5� ]wf�$$dq�Wb�u���3�C�f�����?�X���6�)��w�5��o�^���{�V+;���g9�_���7��/��w��X�{��Εz��@�L�sz)Iϻd��Ӯsl�s��c��8��sG�q�9��ߵ}�y�dC�.����k}�X��L�}��gͷzⷰI�S�k=���3�Z�*���2���N�9d�l��A�=6�O���I��ާ�N߻υ�~���<0�e�%<o����-w��CZ�3���{�}+<����+��W�Or�#SV-�w�n�}�4��D�B����_��G�߷�O�/o�=^[�Ǡ��~���?%��>����$�<I�A� �n�ڏ�3���-�]�o��Em^(��|]Zrwީ�Ӿ^���w%W{1:�����#������7�}e������S�W��y�{S�$8h�UB�k�r�^Gy]�%���V�(�[Y�����i�Xx�rA��̰��+Á׳=���t�����{�1blh��󹏦-x����uʢ����%���jV�v�v�N�fe����C�^ӓN�[��70�S�����[nܚ��심�S��Τ���S�b�$[~����
f���8��3ٗ�ĚsdA�ٸu�kOU���}~>:�YB��d�����b�s�	Rz{�����$D3�����	�'���ެw}loҔʺo���ϰ�2f�{=�@��ޭ�/��徬�����PxC{e���
�\w�՘�3�H���!ʠ�`��$Ǳ�?��N]4�������&5�������w��1]�S��l�������G�Ǽ���<���=�~����DU�x��޷��nu%���x���=���W[�>��|^uߦZ�>̍�~�{���N7��[���K�~4vkN��mS���&�{���׀���|�̠�}ɥ���~N٭L=��lԟ:���HKU��OZpv�<�Բ�tǝ*3[^�8Gs=u��Eb�f5}��=}��j���ww�zkv��0͜;Ws��C�U}�x8Mx���&X��d�E��Х�p��O;��EJSP��6�[Xxcku���淽�V�^���{�)���m/1�Tڍ�5Ӓ�qZ��]^���WGn���s2���Boi�}��~��+�Ε�VJ�T��%`�(�7�����)�k���!9��Od��$^!෼�W�S�9nل�Pd�$�>~[�F�=�:$�Έ�e��t��{E�Iw��)��� 1�\amsV7I�gϨ�ȿ��n��o�x�k*���g�]��yr�<�����'ST�}=�;��;�J�0�����Q{s1[�ĳԍȻl-Y���@�'����`��n��>�����c��̲����l�Ճq��M:+}��yD�ṙ�a��,�W�]p�\^��醖7<s�*�y��Zj�8޽��8C�ѳ�γ"`�_���7�6�����=�'a�u���ߓ߰&!�Pљ���InMbi��������W�k�wn�7��m�S�3�
����;@o��r��]�OٞS�w��RC�j神�ϫ&�47_uߖ��}݄��^�:�E�ԍd:���*�?��g��($Ot�kU�>��?<>C߼u�)ef]����	�͂�Ca���'x��y���o���ŝ�-np���Kٗ�/2:|S�9��Wq�Ă�ܤ;�n���������6��~k��e+�o9�W�:P��&�R����]�ug�~5�w��^�\�o��5�6j���t6�{�
���*G�'ck�Lm����܃1�6���.���nB�㡛4�H����o/Vש�sf���~?!V���+�Sߟݜ��a՝TZDZq'J��Js�a�����P�q��뵖{�����:K�;��m�C�{ϳ�f/R/(�Q��ݯ��c�R�=`o��X<ꭎ�c��l����z���;�_�����}K���^h��n�n�=f�޴_S�W��oǦĚ-V�嶲�9�92�����^g��ϊɕ�j�V�k�`^�c�6�����mC�=g�wo��$�Ў��s5��� >u�[*���y���?�g�wj�p._~�1o��Oaw�k"�n�a��=���ҶU�'���6kߟ/��u{�5}����:\�_���f�ǥa����::.�
g�S)�2�t�ڧ����308T6G�6�
	^� ��8$������L�~O�<�d����DD|�
Y������.ޭca{�
p_q���R�80qV�$p���̢9躎��ݠZ���{��:;s�D���c�?AyEzJ����}^mmT���J���l%^v�Z�<+M�����lV����w4��a�o��Gw�v�T��g��{ͧ���6��T���W����9��t�=�����_f'�P����WU�I�/��]���b����izYYW���50�_�z�q�Y�E���?T��z�͟9�S��k�S1�	��;���0��նgL|����3{��k'}��P�Z~Q�-������Qo�(���ӷ�G��pϺGv^c���m'�K�<���k�qnǜ���%����K�l��Ҭv�����ncF�cms�N��i�2��Çg���h[�ح��̥�(��i�ǵ�,��2��O�y��5����?0Z�K���wгޭc����[F��D�4�lY3"��~$[oAwY-��z#����^����u����o�/4��T��{����{'��q(�b|��G6��]�jaZ�0{>:����J�V�& ��I���V8�M�uu����1�=�3��[F�$�A}]���_G�&���N�1������J�by���X��߭w�]��|�z���2�8�~���n��P$o F���9�C;��v�u]��Z�n�f�o�?*F��~����	�o}�W���
��'�y,*���So����i�;f_��i>�*�^��S���&��ڷ�d���t\�v{3P~��~�����>\>~�.�E�"��~�랞��ď�'{��ǎnwt���}Us��B��_г��1+^O�ıw~�S�����V\<օt�߲vc�"h�%�)ЫG>���;�w3�un<����� Y�ݝz3�W��t�j�ҎF2f��E��@���(U�*��o:K=�k��6ն]���nq�sY�ߧ��گ&׊�TVo��4>�Ӽ��Z�Μ���߆z���s����!p9�3Ϗ��=�������.���;>߿.k�r��������t��M0C��'�Z����<����ez����o�>�ɕ�[���=�I˻����ףƥ�0����@:��5%yEu�{�hΉ���
��]�7N�9�*�Ӛ��Iʄ�H*Èe�|����5h�L!�sB}߭%�ex�%��\��N�U#76K���o7X��z�8ny�����;T)��w�b��4cH�ٙ����e�h��Ώ���޴�{;�u՗����e0�<���	�+���{������	[��`��v@��T9�T�]�x=�C��X�[�'bf��}�;��5g�����H�ٺK�A��~j�������׺�"��ʝ,S���׷�C�{�ıB1��Vv�z��y	9^''+NL��}��ҹ`	���5w�O��̽�B��������Ͼ>�>><��K��=W�PO%��H�׺�x�H_{g�����V��I�3�����j��/>�"u�1t����Vxl���rW�R�����{�y;T�X��^�7!��ٚ�^�G�'��ǧ@9������{+��c�����)��i�������ǈ���3p�/�*vT�2���P=4�^R�w�3��"{�٧r�C��Fl}�AIҥ�ܬb���̡n$��"Q���3:�%�g]]�	X����n4��!��	M��N�ʷ�?#�x ��OJ��y�S����bl�<�M�v�Kv{����wODϧ�tO�]����<�<�Y_zC7�ukw��>>�)xw}EŰ��{�O�<������P���N��q{ޝ��ˁm��{Ĕ���1T˝�{غ�����S#�3��ڟ8���o��#��ώ�~���bs��w����W�=�z�j囃pR�S�W�=R�#Z�=�M٥[{��,ް�ϣ��M�{�.r_S����㒇I���k�&��=��:R�o��2����\�՘v�������9���1�Hl%�M&��z�46�C�y�P��_�x�i���T��9����Ȭ8��u#4�dؙ2�}��Y�_]��(,���+˹b��_�?f�{����]��ߴ<�/h�G�Sf��R�^�W��% �����j/���v�[�����9B��y�rA57^Í-�&3��oǨ���Wk��D,#�J�@�w���k����l՛�s��*կ�BR��9+mH-�\�N�-�t_�$�l<���7�w!�Ԑ�J�O��,�z9�&�r��9��b7��W[K�j�©qo��u.ޙ�дq��qm^S(V$�O�w�9ٹ��]��KY˥�>��5	�F|�~��02����yw��gR��9�M"��ry�r�'� o ����;��v�T�]��7%"/��|Q��Q���oQ'6v$����� T��ζ̈�=R�`lz��{=�<��O�����Q���z��6~��oz'Ր���c��=h���e������.�/K�L�N��?uA����$��׭/cf�L�@�h&N�w�":�Gs��&M<����ȍ�y��Q[�����#��v罴�߀n���}f���zs��LQ�1�8���[��i��N{�a̳Mq�χ�Wo��S����^��Y�I�|ߗ����I6�:�>>�C/݂�,�~�^�x���ڟ9�-�ϭzmVS3N�5���{_#���T����4~��E}^P-���{���@g#�`���^�o������^�O��<}�>7�߃�� �U��쨱����t�
y�W%A����UX��
X_s������ؽAy����i::V;����"7��0=���Lb4�"��\���K7��Mm�B���G�[��? �gܺ.8�+�x�ه�LȻk=RV��h�����'�I3!�M���*��8i�yč�r��!wI���0xaĖ�Wޞ��U��x�Ggt��y��lr{��ar���4��C�2E:�8`욪���8�"+X��Ky��n���N��r�w#S��,{�+��^�Y�%�z�E�����2�w�-�`<N���9���RM� �DӶp$4�6�PT�l��hnS�x�w����(�&&�}�0�N��9�[���ʚ3��p�+zf�,��T ���d`MǸ��%\@��o�|P��~����̕C�oէ�e>�X���fچ;_thA�9��N������Z:O�D:�D��[��v�[����ҝ�r���΂98cN�jkL�������5�yt�K1��v0{��q �2D��9-����˞$'���n��20��1zO|�_�QOV�@�<4�s*m�Z�;D���/[�J�=w;�Z��f�1�CF8v��v9rMQ=����ѧx�P��ՙ������`Nc�u��6ԓ�l�Z"}FҘ����c&��2��-�7y;1�j�aa�s�]]�=��N2qa}|�f���V���ղ�Dզ����ט�y�Ņ�/o��}m��R���l��1���t��)C�9��.�����2D�j�~��R5�� �R��c��n�'Ԕ�6�NN�eH�[��Ƶ��GT=����e
=�<3n�ȭ)�w[Dh�E�޽H�-hn���}<�^�����4����H�]�[ض�b���=X�$S��Ǔ��$���ºtDb}���a��L�����A������Fe���H?M�3Jb��7��(a'��X7�T���-�'7T��ݩP�Kgu��$�V6ofR�&����4u3�J8�0��K�<ʾ�ۼ�e!�&	m��T�)�)
��&��2jXv�*±$�J�K��@���i�X��������F0����D���/d����U��3ǧVU�rv],q��Aj�.�^[u��ʬkz�*]V�7��մ�V���ԓ�'���V��Ј���%��k�6��/J��,:������=�ڸ��e�����	sDzo��5P�2e~�=}��.s�ݞdp+|�ȥ:A���X5����n>ڐ;VQ�K�jM؋�f�k�*l�f���ff�8��RFCjr@��E�YݜV+Ġ�ջ|��=
&p��l<qV�f�v�soj��Q�v���f<r�`��7��Ұ �R��Dn'm����7�-�dK��VKp������'���^�����ZMy�i�B��"r�72Dhx]ꛬ즔���q�-��vm�R�:v.����R�@��}0f��|r�۝����q=�;�����Eu�i����鮈��v�lF�v�d����k�\���h��k׭\4�=]5�i���^��l��ۂ��n�`�ڌF�k$���Z��ژ�LU�޽w���3֣�ID����=i=F���v��%>��h��(��ۻ4����6λoDճ��z/U���P�յ�=tQ@ⱎ�5��g�Z�Ŏؤ���k�=lzݔ�Y���;��=���]�:5��n�o]�/[V�o]��]�wv��]�K����� ��E�-�,��(0B	�AP�vq�[�tm�����uůW�7`�d�����6��Z����ӈ+խb�k���]z�k���=�P���=ws��V�4i�����Q݆��������d�t���ڛX�ӈ��z��n�h�F�}v��X5�m]�����S���4Pt�lM�����5ӬMTl�:+��CX�mX٪�@�c�>J�����߿Oߺ�,����"��}K!rݱr�٘���<"�.�\[r�\��H�S�d5{S���򯗒�{�^D�1s���̍d_ u]�dX]1�[�Y���M��oFl�J=G:}~�n�mz�ז�K=�[�N��/�ȴM���#���s��|�D�Si��3U	���7.�Rk�����%�=IY�g Mbf9w(�8#'����/2�X
�hh����\��ŷ��}X�F�]f�c���:�4n�Ů���d&#���F�rp���qG��%5�2�ᇍ��\��R�p^������2r�K6��Ǡ{%��}�ʒ�S�j�@]�)[�:�cἢ�d��X�]U��^���҉tA���d۞W2�@��ת1���&M�c��BE���y,���HG��%kv��z�������tRuϩ�?b�޷�	N�v�vZ��ʫ�r���x�:�1��J̛�J}��Y/��

Qqa̪<��i�'5P��U�5������K���ҙ;w���A�oٜOH��#����wLɶv��Jဲ�AR��	P%��|��˹�}|�V�_�R+���k�9r�:��[�9�د诞��E�y�WcHӹʥ��2��<����6z>�᷷���o*�-�!qT,��R���$6#;S���WFckheJ��Y�)���@E^��,x�Ӆ�^8���!�K��~2�d�|�0i\󂔬�BV����a���ǡ�;��� V�tZ�-��7e��Lm��U���d��R�Ƭ��Ǜ�e�?����E���ѝ)���h��vx�>0�e�K�sЗ��lT���U�lG�z�V��B��{�BA�׮�t/v`���w֟�h�J����/�p��ux�z������1�;g%��{��phJ|w�dR�i0�[<�^�Ǫ	yXv�>���@n�g�
?PȞ���ޛ�{F����\bQ^͋�#����E8��3�lj�8�nUQz�!�Qv��p���Y.%V5r�㢮� ́���>)MBC�9�d{�i��Me��1���8�0��6_�x�S�t��I�^:�zV����P�z~L#�"���$�?�������Lc���]�p�b�tn��Z��:�f��1ݹ��zh��s�^��`3�}s��MQ�W��d]���d��"榘cN
zr�A�PY�[����ROt�+3������8h� ֱ5ɘ�$�m
�M�9ա��g�9�%Z�&ޯ6Hca:��]���)�J7�G�]��e5����ށ/�o�	Gm���Ւ#i��{�`��Ry�e�E�K+¶�*�Է��}툽?�����4��9J����K������:�池;?�ث׾S.m+ӂ�ܔ�g��� ��M�;i�}�9g#a���~���N��Z���YV�K�g�f�&�/�֫�B��'G���cR'�;u�ۋ�]0�m�M�BL{y�d6�����u�JۑfX�b���̚��f���>���38��1��"�h��2d��6����Y�V늣����Y���|�[�UW28SG�K��ʏ���qB�i=Y:|�ӵ��}��G�{Q����p�<�,��.��M؆j�.�elo�<�/Z��a����� �dσ4���(	���Q�9���g˄[�g�:���1���#b���U�ݘk�b�A�R�N�ׇ���f�f��Ar�aC�J;��==��0��Gy|,-+�	g><q�9;�.be�;#���}��j��{�"��|lÊ;j��,��I�p��K�A �=w�w�.�Q��ncQ��8ئ#��̺�6*=�;8ػ�K���Bz���q���kT>��Pz��쬎�W:3��{"x����������1#�[
y�Oۺ��B��)nu����qP�{4�Q^��L9nwb���ǫ�O�sJ��ao�ψ@��]D�`u*�s\s�LJ[c��YX��M{��2.4�Q�dƙ�C9:� {T����I��?B<�DAQ�_W��埙�DLk�x��>3Av0�Y�.}xim%�&.�<�7��޺t��Ҳ�i�W SX�;��,�0��++�[�7&�z<�٥�O�𗲂jjڐM�չxk>l���WJg[ڙ�oe�{��o�ܛ�0�h��W	a�p���N� ΓR�+��>�K0{W�别�'�F:&x��0Z���蒼�[���|���\��ûK}�-NǗM��E�G�Y�y{�oA�� wEc9��<�ߗ%��o+�P��mJu�>����<����
#'*��b�cە� b�`��I�l�r&�M�����=���?n�
q*8�1Y8}�����N�M�� ���5]��p�7J��U�`��D�R$�Dېz]��+�lĕ���5���+�ia�2�[Q�)J��р����2J��7��t��鳙����a��e�=2+���e�n�k{��.�Z�mX�i{����i@JMn�S�@�_ז����ћg��0͜U��E�fu�p��E�j�n�Z��
�ɁB�\S��m4n�1Ǳe��2���>�Q��<[!�b�]=D��1)� ������o��̍�j�~�(�|[�q�����Oy����/���t�����Ɔ���W!Vf�J�V��w��{k����N�my�{TX��t��g�t�BXdF6��-���(�/u�r7zs�庻4�3��{oy���X��n�E}gm����[[�	;���6,#i�:�QV�X�Fk���+U�y�{|���Y�r)���&�-nq��F;C��u58������@n�6�(�c�ͬ
r�wL�Sk��Am���%��	ê��K�/+9�F�NOh��,I!bA[�6~������e�A�sU����N� �yO�1Sї��V��oRʾ�����G؁>͢�h#��.�����������=2�V^Et�|�H���Ѵt�L��|O�]�����h結p�C�Vl>�>�n|/Ϙă=ʦs�e�uvD]��ʑ�^�ޥϺ<c�L�odtԘ�H�R��`G�c���<�wήc6>�54a�1b�$��@H�I��*��k9P�&F6�bR7rw���"���H(�^�E�gyA��
�)u�¹���1�rY���a�v@&�r�9����c}u�P�>JN0��1� ։~ˠ�v��3q�Wb���_5u�Wɘ�{�@�vz����Y�T���.�A)A������X�5��#U����`k�Č<3)@Sz�K���t��bT-
,:{�DK�)�"�h�O֔ק�/8E���Η�6'|t�wO�Ύ'�F�\���ȏ��6�ء*�5V�-�.�I��jy	PGW5a<(�6���Aj����<�5ډd���{��T=�晏[��%QO�ҳ�����e��VM~�|K!���}�������k}=�?�^M�X+�g�s��$�a>�#5�ny�f����
4\�fM�k��\�,m8w��s��@2]ҦYE�2����P1}��Eu1,��q�;K����}ck�o�@��g������L��o�y0��B��1���@�x�mVc�]�ܣ�/��2�tU�_����V�.�*����ا;�௕Um���v���Џ���:0�
QqneQ���ZruH��U�5�g��g�y¨�MpřS]�^��O�� ��j<�^�^K*3�t��;z/΢��7��L����+cm������}����m�#q	�-�"�SA�n��L#e��<�J�z\B �+6��Nz{aX?o��Tkٷ#:Đ>"��1�0^b�_,�1WG��J͇==�a�Y�Ω�5�����I�����,��[1�\�s��G���������M3�����|�s�HP~���q�8*�xm���	�Z���5�^;�};�=K�ټ�C��s��)\��ew��Ŧ~�:�ȵ<�<͑�5l_!⌋b��FP�U���4��{��m��}Y[������$N0VjF ��<X;��2=�F�,�ۑ��0iމ��'����fj�4n׌��oct<��LW�P�N�K�)����oαL�z~�&ɑ۵��3�����6�&���2��[֕=;��֕>Z֫��xF����'t�Ǻ*�礭W&�J��X�a�4�"��������m]]���"�N9y�
�����
z��j����/+:V�ky�%�rm����sκvWi��q��]Z�d��-xeج��ϲ�!.�A6{j4���XZ^���8�z`8������WTӔo^E薐Q}v�z�j��\�/��7�g��L2�gE5��4B?{�/�Ul���j�c`�h�4��Ym����)�=Z����s�A�s���E4�B|s��� Lw��8Uiɴ-��ļϭ�.��>��+���P'���	e
>�*��5^�>ƹl��h�o��őSѰ��g �K�X�)��y@�~8�>4l{�W�yz��Ez��Ũ��S���x�����C	��G0*?W��Y�x�GI��u3��=��=4�����͍���XGXg��k3���d��d����C��.�g�=�wO�MQ���_а�cO��f�&}�oޘ'�KYU�u˶R�={N����<��yc����i��$�d�s�>[�xva�=�ah9����	�
+�S ��{�bf�9a�W�xZ�^oZafa1N�c����Ó��w����D�^sh�g*-g ��Aڦ�$vp�e�I���?Z�QYI�]�$�Z��6h�Z��,w�{43E}��r�lJ�F�?U�^,*����8�e�%�E�&�i/>��5N�*>;/,:d�(MA�Ɩ����L5u�ε�A�GW����
�՝��i��:A3�����wc�R/�����n�Ҕ�i�:�ӯ���i7�T@e���I���Nf
ѝ�?�
sݯ�g�L��M�1	��f4��Q���6/J�2��j׬�p2Ғ�ޝ�o5�B7��a�V��l*-�9��c������S��j\�Yy:|M��T��f�FN�K��`��j#�B�̨UW�@Z� ���t_)�A[�!'����Ʋ�;�ӆ ���8gW��%�����$�Z޼MsF=	5:g�r!��1�}�Gɮ��ޫ�yx��G%�u��Ә���F�w�$/��:��S��}ɑ�u��0Z���$�s[g�dH�7h��1FS�K?V���V� ����<�Pփ�|�h�}�<䃜�Y�COς��g���u������GA�5�E-gk\�4c</������]�A���#�6�O�����4#'n%��{&���h�M��?�������k�.����} �c8�MjBmP�����Ht��r��Ԏ��I�'ZEPÕ���n�-훌[X�L��0��FD�|^��V��pr����ۮ���i|]�L������Ve��[-����إ+��4p�*k�cA��&I��{����}�~����k��:�P�!R~�i���Tf߻�����m��H�l��f7 �L&�ۗ&a���}YwKᜰ�|�tOs�%?dȶ�_wg�&`���i�N���nL��6�Tz�����M�������n]���5/�'1������o����S����ގ��;�S-Ī�8*�7�6�AQ},H�k��J��0��Gۣ��aؕ�O:>Y��Ѕ?�i�l �7�C��5(��9q7��N�87��ёf�H�"����	D�x�-Q����5F)�N��8e��8���flv����zw��Xlr���Լ]��
���U�7��z%��k�S��^^���O���
�u�z����Ur{u�)P�h#Vo2K.���ہ^Hp�]���G���o������3���ON�7��\��=���ȇ�L�j���ѣ����3^�;����j���#�ǁ�@<�T\dE�>11^���^������-�yα�mX�or����(Z�g�V�F�p�;:�8v>lx��`(>}�m4�^�jjț���oJk{�\�=���`t�'�1�}��2������Oz0����F�4�����\��������윷��5��Lw�m[��Ck�xᐵ�%;�"Ľ��#[�Yu<�Oy��;ޕ5pףj9W|�81afDuƙ�/yȴM�}��c�{$�4��4@���gOl��ֺ�l�l��1���{s�F�ߪo�Bw�U�o��Q}z�r����ռp�(x���8,�߻�E��|r)`����ͭ���|�Ѻ=�pwd�������H3��S.�����|q,W��#�yݐ�������ێ'�㚍��د4H.'����U�1��(<�~��t]�G����KB�o�BB�W�: vĊ�;+��y,���6�A7N��]�ڴSK6�����e8�t���{��M�!RN:�M&|�׃ס�y
�O
�.���pnǻ҈���6�b��T�կ��ށ*؃3!�i.����E��-�pځs9J�[� Ɉ�ɕ�i8۶�+kMW�<�1� {%T�P�VWM�o�ޝ����H�<X��H�=�9�yw+�6�`��!)��aN6S�Y�ff"=N.6��9��=�}��P����GְY��,P��0������Z�_-��j1�G5�SEn>ŧ��V���99/^[��셼_���,��׮�9}Ӧ�C�����W0VUeqTMeZ=�7�a���~��1�^ĺ�ܣ�%�o@|�{pf^�:��DO��<��A2�B>k*��~��ƙx�����;�e���1%ex�0y���%<�0��A�<�Lu��b)=�����#�߶��y+���N�FZ�_�eBWYpRG�|�[�o���}��?�������?C���G���}]o�=������s@MDڲ���n�Wi^���^����Z�\x7�a0�n��$����M	���7�n��vU�7L5fV!�-����u?q���1g:<�=���$��r���#�zJ�B����Z������,Hy0
y�vA�%
Yx�����zuǜ[��^�]�b�|�S�悼�Ǹ'Ϧw�8J���C����N��ul�AWC����˂��kh�w2�����*խx4���C�ႂ&�ju�I']�YE��NI���񘎟d�����F��٩��g7s��� 䴷<f���+ʖ!��+�����n'�]�T2���d6��Z9Z敵}��b��#9I�֬������"r��}�D1?l��p���iם>��(ל�\��]�Cy�3�Q�Q^��^&�7��њn*�Q�#�x������P�=��\*rW���o�Ո�y��zV,�57�@�jƫ���-���R`��$������\d����%_[ʘ��Զ-��R#z�D�����mmpڅe��e�Q�u������LW��ÒR|�*�q�:��v=�y^�x�wfs��=5$�mY�l�ou$R�vU��p
K_b���}���s���R�/3�j�s�T9�B�w�5N�x�n9ҲZ鹉ädw1�T���Z;O�>rk5�z��ao2�60���K�
���BF��g������l_hn�F�RRP�CD��mk��ܷ��Osz1�'X�d��"����'.=�IC
��wo�����T5H� ���z�8ta j�N܃o�"2P�g�;f��M	�J'(7�1d������)`��\���Klݢ<��c9�-L{�����:�S�S��7���^,���y\��}v3DU��F�ɤ&�^���˭�J�\s��ꇦ(��{j)w.�����X���oz6ˮ��I���EE�J�M^�Gpj�
x�!��pu�phEr��6��_,�5���e0�c�9�0O���xk�1��i8��]���p׋m�MP5e��Ϯ�./�ʈ#��L��}aL8��He�X�n�(�XP�IZ39�2B����Ha������wJ���Crd�%~�f1�D����:I.�ez-�^�sD���d/z�cɭ��n�k�tH�삹Y�띢�>���Fx�;X��%8_n:�|���J�8'*w|�$��<o0iX/�7��vy3�z1������ٻ�_dՒ�|ON*�􊌧�3iO��Od���h�O�!�az�{� �/h�lѻ��d�N	5��Z�91�J�ּ��������� ��%c�n��x�UY"u���/{���s5{�$F���9�㽙����>�����ڼ���i��x<|�2��c�^���v��M�:��w���)�<a�:����,�a��7 ���-��X���3*s��tF.��T�Kl��N]�t��6��>t�k�k�J�<��T9?���6X��֌�*+ʶ1>"��_na�s*TΣXW�'�v)���s�S4��v���f@E���X��������}���=����դի&kF;[lUG��k[`�A�3t��jŴ�ۣV�C��g��N؍�D�F��1F�[���uֺZ7a銴���V�Z�[b*+Z�n��SM=�8���7c���j�*�؈��k	DΝS=t�Tű��]hm�3��*������:�ւ��:4�d�uVɠ�QCA��-�Kn����lS%����ą:Ӧ��F��D\�+��AThH��ƋYN�
��Wg7a�I��ں]t�蠧Em��{`(�E4Dz�T���4t=��Pm�G�1j��n�5N ��U���ݻ`���;h����-�Mu�$�k5�����"#c��.��MoC�����޻ׇ����~bR��t�e~hF��	�)L"�ܑ���ཀྵ�=����wo9vk8F�v���.:��]7��♢"_�{��4D�l�h��^q������1�hY*S 2���kg�tL�|Օ�`G�:(�<��iLd?Wl)[5��O |��'z��!��?S�f��[�q8��(�Ơ��FT��{��BDA�дp����K��V�O�ԋ5�]km}{�Ρ�V�z�_�]�O׊)ɽfn��H�������#8<��'�w�	�XZY��s��X��Hr�d3c������%����;�[�K=�ږ���R��&��7�8���S�o�	�����w�?�:9�3�/%M�z���q*�$��c�qZឿ<�,/���#8:&uK*3������8G�*���O�=����:�o��5ǝz^��j���L�z�e@�(7X�6����	(�M3l�kta�4��Be,C�2�/Z�-�U��2��T�s.g)Z�3�P�-t�~Œ'kܫI�1Ia�C}�Gݐ(Φ�;�]��
�_@\�)���%�'#�O��>=�x�
O�q��\q:�eSL�k��̴	D�닽;P�o!�u�oi��l�)�M�f��ZŬ�4[ޞ�HB�8�����yB���L�H�s��@X��i�%���s�h�Y7�*�2XT�TMِe�������?�h@2���ڙ!<�^�n���z�$����*]]�ݼ��I���k]sL$2�����\���Ym�����..�E�����M��y��x	:�agIn�4���>D��b���3*�_ܲ�^����@{���Z�G,���4T���<�&��'`ꨮ�A�/�鄝XOǟ��gz�n����v1a�Rva�=�6us���T���^��ǴR�(� Va���g�Q5)�|uRYth��-q>�����]��w[M|�=��\����Z���~/>��Q����.�J���sKcOu���w���sӒi��r�c���Ew���
ݞ��a��6/�[t���Lػ�*���������Г�|Y:�|����ë3�w�7T0^�k�OI�6� ���&?b���m	�Q�m|w�J���m����h��OTU��Ҟ�>3��S��A�()�f�������wu{�{M_W��P&YS���w�ֹ�7_�)6p�S�lƙ�\�gg�#�R>Mv�|b1���U�d����qy�>�4�G�b�����+$�¤n�D�uO�\�k��pW��z�f��ѳ���:z�i��\_��W8�}q9�m>��<]��l��r�C�4�SM߾��yr���� pg��>�\f�"ԓ%�2�P�tz�Ɋ�q_>�ġ��14=���lr�������^5�#YSw��oT��HtT���D���f��R�X�4S6��L��.�O�9R6�>F�o7%�]��o���'^��v�^���J%�x펣"���|��݌��N_Ϯ~�� �`�@�騳�`eF7P�-m��XӦ!�r���<@����&���d��kr<��V$o�Y�Ѽ���=�MoiL!�dR����WLZ��Ϡyv�n̵��ɪ�?�-�����++_U"�`�8��2d���(����u�
a�����qSؽQ����湲���$a���cr+'�ޟ�u�
�/�-��iv"nՄ����}�9���<��#�r	o���G���P6D����*��9�j�n�Z���rrc�S#_ZE�nb�<�����[���ggy/��m=�����R��s����Kwb*���u��ͱ���Ͱ�%�ک�pdFT�up�-ـ�a2#ӓ����ꀠ�H��4���I��?6����t�W�'�N;��S����/P�Wy�H����`�K�1,�)��YԌ�@�n�x����w&]��A�۹mf�~�[/|���k���t����J1�`C�����S-�7����ު�U�tp�݇]"/1���t��q�a����PLw�ʒ>�	�y1�^3������wЊ�;?Ɩg��h_�tlj?iM�	�=��]v�n���=�~~m�s\h:�!�䰳���hP��{���eL�{K9�*�q�*R9�^uJ��=  (6�bU��s�*�u��Im�ڏt��H-Ol2��GC�.vL쩚ژ��i <<��3xxL�
��cBu���jUm`q*�<�����Z�S��3�n��8v'5�N���q�]Գ�;�a���qw)�8�}��<k���x7�c=���"Lפi�h~j�������ߨC{�S ]��;w��xAU���FC]�$F��?Z6���l����8j26o�bG�؝Pq}g�=f�}W��讀Y�G2@L�g�`G\i�!{���l�zB,fm�>��1�D�������=�f�1\�B��V �lL��H�	x�L�5���ydK����^���O՟x׊ұ�:��͉Ⱦo���s$I��J�޲)��R�����[a��S����z������.�h�,%Fr����d�!),���\��]���#�s��}�)V�n��blgv����bOI���&xx�BuuD��������\��}�s'�n�u�[L��6�0LUH��q���Cz������=#d7D��X��p��y�yv/r�Y�b�M���=�u7u�즁3�+���]f��Y�.��z��~�9J���@�xE�a���
�~��ż��b zY�J�[��AZ&K�K/F��X������T�5�r�*�Qӽf�YJ|�{;ܲ��8n֮���Y��8cJ5!���\� �e;��xu��֮|���ɝ<_���-�}7���a�������Х�yC��y��m(crY����ҽ<��`� �8DG���b��;�a;�� 7��ޞ�a�D��=x�{+Y�Xd�z�N�'���5�J8������-�j�:������R�:�1����q �^�-�ЮD6b�An���b�A���3��˧i����a�5T��5,���YRզ�X��;]���oo�kCV
�Oy�eg9+���/m+�v�\����"S�n�k�\�BiO�,���,h�|���H��;�(�O�E9��_5�ˮ�8F�/	����<�q�k�<�|�y��Z�{�L�7��0��׽�q��f�S�o�,�|��oC� zv�U���1�)ܓ#y��k�^FE4��3p�DUa`sy�×Y��u�s~�~�WAq�0��"m�D<Ԍ�ts�HA]��^�^,��ohpD,�W�ٖ�
wl��F�wJ��=̙�E_.v�}�H���P��ik�EyV*���Hܭ���a1�hS�m��>��/!���/���2͒�U>4]�~�	{d�yF�(�8����u�b�{�Az.O5�b֍�wusPc�y��|M����eg9k��x�+�)K�6�Vup=]�����e���m�l|��t���Zq5���X�7�Y�Z��u��pn�ʯL�DN�W�p�V�zn,ۧDn7�oT}d�r���W���O��R�&6����1�̊��+j)RL�:���A�|���Q9�Қ�F�V��!�����{��Lt��H��M����S]�?����^�c�(z/K���l�S��#��L峞q�4N�u]���l.^Z���d	��u1p�U�9"�GyP��榹���ߙ�Ǡ-������x�NU������"V\&��ڄv&��b_%��)�<���~�OD�ƿoBeΣ��C[�hK6#��(q��Nc��[P��ݵ3�{4[p�H8�-�4V��,rqn�����6d���~V��Χ�J|��K�8�w<��s����������w�IA܆[e�48��۸_���f�eIt$21Hf�wt��̢��1���Ԏ]3��V,�%��>��]:[�c�G}���X�^}.C"��%��6��gL9*�b�T�G<�<�EJ��Q����Αw�W�
��[�O*��]�oO�+�������~�M"�Y4a����XH�d�-�#*+Pv���#����ʊ��QD�$yx�o�k�o��>��dL�ޥ.6��Bz����L+��"�nnB�[(g}�D}݈+���"l|��	���Q2��LlTS)��-�� kJ�{5�vpR}Qϒ����3��;��퍏i��YCo9,=�{QA�,�\�ʁ��ͅ�SL�ϣ��]Mh�o�{�R�y�g".Nd�������Ǚ]�,Wba��F��[����xvx�3i����N����)�}��dƕY�/�������d�+�ھ��縢��_�jO����ZH9��0|�k
A��#������+<�u&�d^'q��=�X�j�_���.Z_|	�l��X���=} �j������G!OG'Y�|/�����p�mq(*9��� n��^���}�<j��Ik��pV-������c��f�T��^��R"g%'&�Qx�>Rh��z�5,V�}��}�D�̓�m�o�It��e���>�t��^�Ɣ����Z�+�y�.��j�@�ڦ����X��J46�ϭ�����n=��Rs�8:�&ҿ�ݨd]CF�~N0}�?,^��pw���} ��	���z�RI��f��u`�_\=?gT��/���{�g�'�&����<��@(����D5R���X��ҡ����!}9X�7��~�SL��V7��̱w���w:�`~��Hm�mWO9�YJz��R�qᘺ�*�4�,g}��3"-)�\�}�m��k+QQ�0*񢓾��S�6�S�w��o�Y�@a�v�1�1�k���J� �1)�T��Ī�hZ���=�mM����A�Zkfr��u����'<��뼬F�����0Xnw��q������ݡ+Q��=��4��_Wh�Yw:���o��KԚص9s�������R���7�5qX���:�8%�L��x�JĽ����͏][6rc�d�j���e��x�mȹ�o4z�������=����r��_�k�j��Ϫ���DW�����ay7�mS����E'�F�i�Q���p�H�~㛫w#���5��G����m���ɷc�Y>�?N�����oӚ �-ɿ`Bܼkz�'`�C9y����w����v<�=Ȥ��1�_BxD6��!�앏m'+#B�!m׳��{����㛍��b�9�w��zg��nQ�XDq�c��dy�^�b#��3���&#r���"�^ʳcǹz��Uz~&c�d�7��B����i�=���ʎ�Ѕ*��G��S�f1���}��@�H��I�^aE\�:h:�4<5Z��ży48�W6q0���^�"��d��^t���#c�"�*��2����ʄy��C�8���\m?u�>}��D};�鸂���1���
��d����4/d��p6w|6���V�����7n�3�+�:�����F(KĔl�����³�b��į�UwD!\7)?u^q�C9u;BPCf�am ��AHم�)J��CT,!&�r��5���M�#��聊�����'7���Y�c/�`y�n�#m��)���m;��qv�!�1~u�ǟ	�\���?b���!{��1�s�wv۬>��[�9�:��[�ɻ�ǳc�;c�{�d���L�%�0l2��gaFHo6����[�b�V��U}��U�ޓ��`���45�	���f�,=��Y' oG�#��M��zQ�[u�R�R�=�W$N+4����un��]�HZ��&��c1S�6��;ʯ�]r'������	�o�QB޽+�}��l7{N|����W����(���Y)��qu�V'��b��.�<���ȣ�B�����9Y~�n������k��5rE�����R���>��0�!�����k����NL�[Ռّ5[I�V������DY�ˋ�#|��%Y�1���� 0��䲏�`k]��+�(>��3���~��r1��l�v�)����~���c�v��'ا�Zީ���P��D���V��e���8�������΂��R7��6�0qW��v�7��E�"���s�y�o.�T'�Gb�M@_0�˔Ҟ�Q��p9�G�)^+$|&�{Ǹ�w���O2&��]a��&	=K�:/:�ϣ��EQ<�0�����-l��L�1t���ڗv��s���wɕ�}a[�%�zTܴ�;n8�Dwe��q�Q���Z�pg�4Z��ӑ|W���n�"g�b�9�:��U�O;\d:���f���A���g2�����N/���Ԏ��������L����S���3�2�dٴ�+/����:�����3N|�ǆ�5�2�f%�Y�F-����zz{CL@�������y�������4��v^������>3���I��6�#O�KL�X�v=�wy`-����ș��.��7��4g}IN�a#b+P���=XZ^�|�Ʌ�"��@\w�n�&A+E?S����ť3cj�U���T��]ޥ�ɠoz���t_)�%��y@W�#���'R݆���FŪ0lj�D�7%������9q>Q��0ʯ�Mî6�~��܉�7��A=fo�m���>��
m	5(n�_���y�:�[�!��%H����8���y��[Qww~;1�ճ}M3ޖ�d���s�L��m1p�R�rC��t�����Q��]]��pG>��i��k��>���EA=��=	�.��m/�,p��=��c�(�67Ub�`qi��7�����	i�G�m?f���U��ߵVܰ�ze�.�m�;�b�;����Kxۇ�;+c6({�A{�C����d����b>.x��&�����̹��s�V|��j�b��Z6h�Λ2�.����������8�]�Mk=����\�f"��J}�H千әP�����}������>ϻ���ϳ�?O���s��g<�¸{�My�=q孷 �Pn��;J�w�is�0x=�q��N���<�p2?��+��Y�9��۰�ā�'׻h_dBt/y؁{!��n�J�X��4�l�<f�ʈ�(SuB@=ǇD�#tH�#��̹��&��r�1'��5����wMsg��aN�#��Z�D�	�R���&�7����f=��u~�����p#���M�����]n��okH����c�g����R�I�����إ�Q�r'�n����g��l�vH��;BDrd��o�ȇ����d��-TTyM�Ft��ZF��bQ�Or�֫T{��9;�`c'ep�����mM��a����v�ᒶ��d����9�$����[��ƨAɁ�~]�qy�;��&n�p�]��!�ȳ6�ja���4`)Pf-Β`���*�ЬHD���sKk���ʗ�T��_h�����[j.D�s�s����ҪK����jN5��0}{�D�p�j��;͘�����/�٧ؚW��f����w���3�WJ&�����8�U�t�x��5�|Z�u�t=za؄��=﷣ӕ�'�p��Y��I��f�V��m�Yϛ��Bd+���i�i3�G0�i�}���V�X�7' �{���+��oz�^�/h>���oF	Ϲ6��K��	qao/1�{���u�F�_q	�B܎n��|mfZ�Eċ[�~L�˥�f�JLj
d]�,x!�*���f�����&���e�G��i��ӿӼL�V���܍g�{++���,���m�x72l����eIg/�&�֥:PM�ˬ��E*^�Av�S!�IVҧ3�Jv��֪���7��WC����"i�a��G<h��O�`u���:�1����j��3�w��+���Gp;�P�������.���Yx�>XA�:�Ӊ)+�͌d8)�r�	�:#׉�V��ɗ����:�0��&j�X�G�t�ے���>�	��&#�Ql��b� �B�h���5�Xn�4-���]:#3VM˼E�X���&*If���Jkf��-��( T�,,f�]�5*��0�-3�Л%֨�8�6�
���t�+\*���f
�ڱ�c�D�{Q�V2w��]c*�3LeC���d_sqY�X��<�C����gMj�u_6�4Ч�u6����[V��2T��g��<��Rȯ
,b�R��/��%aT��MB�~����D��0j��`��+��9r����Z���PP�3V�t�/��f�O@qړ4�yQ��[\�oV��|�=��av�I.)q�x"Y��ή�,J�qÆ���%�(`˓�o��ܤs(qq���厖b�r�`9��&j{�����b�sE����f��-[Rr�d�a��:�Cg�9���Ns`��A!��R����u�]���ĥu���mt티颊��"�60E���u�Lm���X�E1V·N�bk�5�cA�mک�;��vO]�&#���E���]m���-b.�m���d.���뱒�j����ւ-�SDkj��
��;:�����h�AX�kZ���
j�UU�k��֊����tj�
")ލ��mQ�;'ZTUEI5&"&��\P������wcOTD��Q[h�*���S2Pi��{��EhwY:M�M��홍��q���h�ёщ����UumF���U�^;.��gMۻt��4khi�-����F ѣX�=�֨�"$�m%Llf()���Q�tn�4]�`������{��{�e�*s*�:�$Ʃ�%��/�\L��ߩ\��^u8l��N�-�[�����1
�Ҽ*@��n������X��]�� ���\.b`�����ֿ�����yO7Ť<����LSߝT�]���S�RR��������=~�н�^��~>S�)h�2�t��e���O��B6z0���Ýy޵ϵᙼ���t�s�^��8_����y�d0�~��1���j��!�+�Q�����*����onю1�z�W:+��ĺ&98�JK	Z�ӭ@�ޟ<W��
�	as�S��~��<�v���B6�o��N30m����Ɣe�ϯ�S2|sT��ڈ9�L�������mM<�eʜTGf�Φ֭��m}�,X�F����q�q�kz&���w��y���:�j�/4|���>ΕSx��2����FEb���(*9�Ho��X�*F�Ot�\�k��<_�g
d�-�
J{��W��c@q�����T�������8�[�}9��׫���D�}ދ��C���?y���&} �� 5{�LK�����9��z��N9c.b$��0��\F�ܴ���Jh�j�}�e@��7f҂��6���#:S5`��FC��2!1b$���&���>��d���[a`Fȩ��wj,���N{jn�2�F�r��7��2��"��J���3�zrvr��dR�^�9͉��A!�L���3�2�. <��H�]>���\��.U��~���f"dC2�`׳r۳>z$�v�-����}_U}_c~�o��������SE*�n�R'��EP�D��NDذ�|�Dk�7Y�{g2h�F2#2�:��i�9C���SX�R���)�]cc{k���an���c��Еڮ�^���V`��U�y�+����b{�#�_l�:$����p%Tȹ��l��\�ʪ�9wR��"Zɰx{g�^�݆le�U˶W�2��!����V��S�UIn�	U��:�f��:�3�ו����p���1�n�|���xBn�	�����wEŹ�E:�����m�k���W�f}�	���v�5z9�eB�Rl|����,����g�a�{;�Glr���ؘ���!�]��]�����|����E0�� �����M�B��\��J��	2{�Vچj����c���ty�c�-�KG�5��,E?,�e�ܷ3I�]��Y�q��8�b+��?�~PxO��0Ͻ�
�s��(Z�3T�j���d�71P�E�`�iA�P�-�+������^{�E�^�9�0ώ�δ?ܹώ���c=����3^K%4^Aj+r�U��b�k�cm��3xDo��g:z���7�2�D�G.��J���������4��w�Z��8}�s����,H�N�u��o'Aύa�u�6�SƷq�f��jn�"ŗɪ��v%!]O�p˞�4N���3���r�5Cr^+#��y�өĝU�uC����� ��A�A}ϟ����'�Q�v�C�~��ݛh�,&p����Q4���#!g�Bט�b�AT�����S�z(/La � y�o'��&�^�j������9-��
=�R���[�X������'�Y���p8��/z+�S�l�>T1BXa&n>*������"]��٧:WFM�����u�W��)�l��L�B�dr�`Z{)@Q�R�a���LG�lI����Ě[J��߬jk��yצ��u��`�TO��2|�H�f����{ղ�$U]2[Ȱ;+�,��{C��Te8JOv����pD�1ܢ�`d�^��+��x�&x��M�d�QhYn��^M:*����޻4�<<��p����`��H�p����}�G3������N&��I�h˚����x���ֹa���ܻ�1�Iح5�����R�����-�,Vta���B�����Kt���u��i������"�kh&�����]x�4��^�xL^\]�e����GI���De�(gmӓ���EE�QE�p%@��Z[C�J�Ӈ�d���xO�sǼ�ЏQ��W���[��D;�L*�9C,7�+(�\��&b�W&�n��zq�l��� �#�m��rQ	b >���5"���	�>S��MA�:9��L�;�C"�92F58�j�(͐�k#�[��_V��U�)��������{����f��f5�F����ž�Ɨn¦X���PO�a�����}09�ex�1в�36a��p��˚�}	�<4'㾩�#�H��|d@��iOe,���}cE;�ut��&3T;o�u�P�e�F�7���/Ё�T|^.�yꞵ�4Ȭ �I���hNE��;������+�w���O�zյe}>L%D�m��sV�b�Z_��=#E�뾬��m��}(,sW-Ϻk��Oz§��f�a�D-"m��HųѦD%�k�Ĩ����po��VНM�_�P�r���t�xEkq�V:�O�u�Q��`�00�~u���,����˰���j3�A"6�_U�<z}�fk����-�v	�cz���n��#%�(5���p�ҹ;�[2��ٯ�w�}O�4Վ򯅅������҄��'�8)&�uL3��7�=0�z�
���{����?%�x�>����u���|r�{�w����s/EB��r�-�sJy�n�zI��*���r{]��i��j�Ho��D�[p2�G[ȹ�a>ĥk�΄C�ې8%��}�J�޿��¥�֮b�sa��4ˌ����e�m+4knf<�T�6�9�[tby[�;��Qy��4V �*��ᛸ/l�mU��s�W2Z�}�9��Y�F�����޷�y�OoT�,��S����+���%����5$������;Û���s���_��"}�JB��=|���<jW
]f�/�w�}�N���W1����Q�����'�L�缢�0�nԱ��ˤ�ё2�h w��mk��:�a�O׋(^ߊ���&m�;.m�4�m�\�C����P���w6���J�]��Y����-a�����Q��')X�zY�Co�Tj�-y!�7olm�q��޿�|t�Ryu�~��͡���f��ʔ���t��>�S�G,m�L�LR����л����.=��Du�yro5G�3��-ǔ�/�Hy�4�W��LS�T�G��������W:���7m8^���|�&�����!=9"㚤Z����)@a��(���ֺȉ�C;��a����Gy�+�qy�K��4��؉��ب�G�8ؼ�$�Y�j+v��f'����k��gt�uj;�e�%��Z�O.g�,�l{�s�S��U�LMJ{͞��1�v<ԣ�&�����(;p���=�l�k��H�À�>L,�
�g0(k��������Vڵ��*�aVQ�>�GuW��TefG���F�i�5Ȇv�V��_i������;p���|�Ym����e�R%Ybf'Yj	`�>D���BӾ�I��6-����j]2KR=�yL���.udDb��99����=����1�ܤ���LS��XM,��*���}���e(�m��|{>��Ͻ����}� ��R�Ъ��U�i�[I���ȉ���ץ۟XH���m礟bed�
߱:,Q=�J��	���ȕ��v����~�����e�%��/�s�LM�򯼏�b��Q���ߞ�A�4;��a����v�?]#���D�$�S���kdy�V��V��mеg/ވ0z��ʹ#[E{*�CK�Ze׎��!"oT۸{�,��h�����+yQV�S#A"|Ȃ�nZ��'P�,��T���7��н�!6ׂWB��ڵ�<�CTCȾ�w��E�џL9^�fٱ�N���o	�{[ԉ�gf���>�\�ǥ���SI���8��fX�v�m����E(�3���n���eu�&��k|�O�Av�A�#�K
�L�UL���N*ۯӟm�\*W�m�O�VA�����^�]%��/?��di�Rt
��
r"��%9aeT��Z��3�y�]*�W/fV_a���-��bں�P�PV����ބp��{�c���Gٛ=���ƻ���0����/��'�k�b)?2����S�Xk��5�������q,�N�����`��C��}̈wXIu��hQ����������9Y	`�<�5=ލ�{�0g�NـeǐpZ������Ռ#�9�:�a��c
a�_F��c#�����xu�<��zU}O1�+ݯ��y��^����;�����r����{�ㇹ�8v�0���77�ϾQ��@JhV�^���������_oo��0P���]"�����%��=*�`r���$��0A]�5��^�^Y��3�Mo����mcgNL�Y�Z����he�<��sÝ�`\r�~��rF�Nlë�m�'�����yv>�w���/<�Cc(�궾�:��Ah�S�iD��٫�\#��͊���k��{�+�8c�lak6�yq^��<��FX��P͏�����q�̔Z�}�n��������^=��|�'�V���X��9ީ���n2$�ş^���s�0#�r�I���d%³dX��Z�nAdG�F�Bd�<���ޛ���7揫o���f��-�5|��V ̀�ö���d�"A���].ԌP��$̓X�����\��|�x�/��63{C����W�#�ƌ0yQ6o)f𶐺�C��:z�){��yOj�g�8GEڪ�r�D�oZ�/��q6ß���O䤳'��$�{�(��t�ǧe@ ƕ���V�kJ�w�^(^�.�I��r�Q02~�T0���Ѓ&�^Ĳm��U5k�kBk1t��#X���?Ff]�[a�2�!Am87���6U�f���>7qs>ES�p
� x�v�m?w��!���f~����Oz䭌���9ӠSH�+P��m-���DoK{��[N1�������y�)�f�� |�  �=��Nq��"��sW�;;"�7tHw��n�!���O1Ư��m,1�.ŷ�I�
9{�v����N�2��[Js�����~jWH���R�";��H��S�n���D���#s���&�Q�	̚\��Zrpj�}^�X�X
�''%�?���dC�0 �����#5oc">]�)ODR�:ƺ	��e��L/�}�v󟒊/۞J�/V��땕'Ǡ_SDc���{ƣ��a�*C��%�L�=I�1�ON��!��Z��>�c>�O�9c�F�)%�}~�]�*�>�#Ǘ���R!F,��`F(Ⱦ�F�k֣j��s߸�,�Ϗg4⮘�1�J+���G�ǩ#��~�xD>w�k�%L��1c���j��.���M:��~Uo}Ç|�^_�}�oMsW���?�v�3��I�$ܴ�Ї�\�ιH{�#�Z���y�OQ/f�M�0w)qq��
;^a�F��#5�/V��"m��wf��2�2#�F^н���
�sn �������w(u�1t�D�a��3e�B��r��0��B?}�XE���ȱ55wJ�"m(*"���+����/�Q�z�/g�li+/��N���RO9n(���6xs�F�u�R��A��,-��y��\���.�+ɺ���
�����ru0+5R��[q�ۋ��� xH�p7����)I�u������o`<<�����kt�8�_��ʲY����z{��_��aw��1��G��qB^�v�ըıЎ��9|��HT��"'�ҘLL[��}nQ��<҇r�m{����u\�Z���Wu{y��d��(��4�Pm�Z��G���WhQ�*���fe�_�~�P�m��-ԣ�#��f��OW]p�V��i(�M3%�]-�L�@����b�^R�����lE�*9�oQX�]��n"a�^K��+lU�)�b�mFKG�+7Jz��(J`s�[%��چ�6p>��TtN65��.{�(���e���^ŕ/�h��i����C�=��&��f'g�깜!�	�}{:ŨGJ���*�iF|�[B�����啲���,1%Д[]m�Jg�NG�����`�7r!�*C4����;��]`O�lK�Q�F�f��嵩���xA�G���:����t��ݘk�⟡p9�E�O"�K�|0�h&�7'c0���&�z��GE߬�
gg��~V�G�b�&.�yͩ	�90��c�j���~��d^�P�� a�k�Π��}�5SwϬ�3S?��߽2�1���͊���~��N�@1e��;��񎐮J��K嚕^Q��Xg5��]�Q��\K�3���G��գ�=]�]:����a� N%�c�m��6�7OM�ҝ[��Ffu�*x��t�=Y�#����?�}�}�� �KHҤ@(P%A�cY�IU�RڎT��=)��3�,������D�$r�ˆ�����[�>��=H:�]	�67m�b��f�v�:��Gs����;�Z��A�ϓ� ��ط�B����6&�b(��9�Y��TS)��-������n~�x]Ll��k��N�i@�e��O���U7���N6�.�H��_U�1c^��VZØ�qD����k�1�I�-@�	�3�R��}y�����yZ	�.&lGE⟡^">���W�|q!{�u�§u�'��Ѱ�4��7��[��s���^] 7���Dt^�����^�Ћ���o5.y��9�f�mGT��x�YNM��բAlQ>�E�חHm��m����K{�A_N�e^��>�=�Z���\�SW��2=�_��پ�$M��X��D�����Rh;{J8w�%َ�x��d�B�f�M����4�>]�:n�F��lnA�A��ʼ�Ь{խ"��i�	��b<s�cU��Y���Q��2��QOy�Ȼ����}g3��ʭ���oiThV-���@<��o�������~����x����7��A������ڴ�q�y���j6�
n=�t8�oB��E��5EC�غ>Q��z�x���\85ԉ�f�@W�$�73J�u"�|��iM�52���Հ�n�w�ǳ����k�����||׍m�̚� -H��Uֽr���%D�z����cL۱�
&a
�7�f�8 J��euZ�w�m\m�s��J�Ҷ�����jj1`��VQ9��q�_��"�ûe<�#���{85��^�e�4K�hpK�8���8��tyA\��)����.ҏ�@���zYg��ՕfMC06��=؇L��Z��.Q���3oxyt����Ү�I1�Q�}]�p�o�wS����$r�Vp��(wWVm3��)l�Qi�<�\^��a�VĘ:��	}.s+gv�|��1ə��}�^�[;z�yPv�j@����M��W��,ѕ��)Ʊ#'ilcObX�=��w�j�Jh���Wd��}�DwH3zP���(^+2Vp��."O�@�5�d"�4(���u⋆t<���P!�dX����!{�+|�ɺ�]h��ƹ��R���{�s^��<�ڹ繀k�.߰�kg���x{�P3�Cޫ���=�)V�o��-��������<�/T4&_[[Ƶ�L�\��"Ou`�/���4�~XW��HQ��ۭ�x��ysO�M:�=�0m��EӴ鬆���(�=b�\�Z0q�U��a�<Ƞu��7������f{�ʢ�*6��s���F��&b�s�{�n��|���@u�&������y��Q��� ���\[��S�C��X}�F��ק1ڋ)n���Q�k��;8��o!v��Z텺녘�����YkOIxʱ%�W|��f˰���Z�����]M	��',Ӭ��/��}�-�CDա������K��UC\)�[�k�J�y:RҜ���{U�,#�:���*]�gU�۳:"���%h�s�A;5���s�Nޔ�.Ƿ���n�}��^+�).WX#R�7�"d��#�.1����n_S�s�2����;&��a'؜�N�8p���>��x������(LZ�X�>o<g�a�Q�J��X]<�Y�<ٳRS��ɢ`V�G�,e��-�^v��w_u���y���{=C�.�� G�-�C:��D";Q��}ܪ�h郉�X�Ȕ�p,����Ղh�/�p�t� ��Hn�y�ݞL/	3؈�Ɛ���nv2�ڪc����j��!�i>9V�*��p�晖���&���{	z`en�y�hڬE�:��}��_Z��s�5��g��<+Z��3q��V�q^n��x`�=�՞Xr�������nםG�����h�z��:B�9G��]��cM��m��iZU|�@��'}20:�ы�j�`I��5�6o^:�tbLU�֬�(]�nv8 �sL���c�H�/6�1���[�-�ax&M��S'�H��c�	{��x�x*�Œ�
�I�����h��I7(�E*P! L��	 �LSg�$�g�c���P��t퍶�f�����QGY��h���jў�wX��{w)�&��Eln�E&�Ƀ�nڶ�EF�P�U�J �m�����Y(��v"6�Q�h�g��kQm�b	�f�1h��΍�1�Z�D]"��đME5Im��6Ŷ�\Dݢ4�P[f�1:6���4v�U4h�kTi�whۻ�����km���u�����MW`�Fl]8-���Gn����;��m��Eku�) ��Sv�u�1�ۡ�1m݂(*��Eњm�֚:.�U����bkX"(�,[��ۣ7QMkE�nx�f�:��⊫��g���RQ��V��Em��΋v�vઋ��S��#V�������5�mE1�]kv�탣Uc�wu��+F,NcN��Qձ�(��*-w:�l�ͳ��:+�8�=���:�v��1�mrF��:-�`( A � XB���N�;��k�˕�jX��͊y���dp��7Au�;�6A]�s۔�ʕ��k��|���w�糽�7R$|#w�q����0B��M	 Я{��y�w��[�=��Hl���������W������Ǯ��.^J��s�T�q�ΣwuUXlJ�uQ����뻆$U������G3�R*zZ�i�(�{�H������v���f��w�W�����նՙ:��v|}*���)+y�f�`|r��x6��rM��#y�7��������FGj�nyx�c���ְ�t�`��O���m��z��F�S�6���Y�pdgd�VسU;z{3�؋*y=:��Ռdf)�vp��i"�zs>Cw/�)ڌ�k���F�0B"5��*e�=�h� ��Y��[|���;����G�0[z��iJ���+k^���A��C�I�^y�CCk>�M6�O�t���,�;V���K��LaA��k"�u]����Ǣ/�0���Pb�S����<��w�e��e@���4!tV)���N�}�n���'�}�l�?�=!^��*�D���@�F9�g���)���~�c�l�X�~�N�WP��\�ޭJdW��7�uȽ,��zY��~�_ڷU���x@��Y�[��r��'8�W,M	�=��8��G�ʺ�ǣ$B�SqZ'֟���EA�TP*��2-�-�U�?q�;uuی9-�p������ϔT�Y���B�-P�a�J�ٓH��&����������wǿϿ�o~����>�}���R���
R�#HP3IJ���ϟm�k����U�i��7p[4q0ISi��0�X�	x�L�|UbgzL%�,�)A3�R��E�M�i%��&9���y�R����E����sT�&��@�\���~8{%�̮ՊMק��VV���&����*��`��TW���Y<R*�7=����nG��]��=K�ML�][5���<�,�!��:H�I��iSR�q]KEc�x�&x�]q�-?�>�	Νk�gvO1�Wv�u�z��r�EUa���H�8�+�V'���	��i!�Ӻ��k�E6�J�_��궏T�_�f�J��ބ}7��U��Gc�|�
Z�D���}�4�p�uWC��R���E�'=���Z�a�@������;!o�˧�)���&���L���)��\�.Ψgm⤷9���u_w EXI���W"�Gl��se������f�_N!}	���p�����(ȼ�@��]`	�܌X��l���;���mK�՜��,S�|)$G��@����?"y�H��|dÜ�M)��'�_�*�k��?,o���Ɠu���
��]��&0�̛���gM�U�{Y���S%"��{]�*]Az ��c=¸�cẺ��ɫ���ȆЧ7�<�|h{;˰I`���4r�����ͣr$�!�X/�K���k���ej(���q�bu�^W�_�|��a�3���ߕ���Ŀ����߂�K�s6�����<">z�T��F.�t��Out�߮�K}�J��p/�[R�XˠOO����sP;�����1K�
�����2�َP�����͊���i�v9�*���1z�I�h� ;����ʾ�v�#Q�"lbF����Y��BcwL�f�F��r�G���N�涇[6�@���(��%ꑊ��L�ˍ��u���������4G���甘<{j!=������iz��q����{�(�t_*^�=�Y3��q����S��K���g�ހ�GF��sR�.S��h�țj�)�3k�!��ұ�C��m4�z�5;j�b�Wk�^֋�_+�����)�(��3M���c�K��t�W#��#FI茻��{ A��i(6)�k%������!��b��/%EC���.�ꃑ�YS���VfJH�����QI�@Ww�T�t��2/�P2Z=�]����б�Ss�}���q�z�e.��ɋ���ɖ9��p܊ħ1�����Ƽ����g�1��;b�WjQ�C�����-C `/a� ���=�k�A/Ev��&.�J q��"��M��@���a��2�6T�~U�g���LE̑	��\7�8C4ҍ��0q
�ur]�7��m��JK�]���ěf��h��V�M+R|~��~��T)
V��Ϟ��w�y��]2���:�q8��v�3����V�L�}�T�gV׼����*MA���f�a��+���YB��<�u�
Ԉ~	��@!���f��(���E�y<S~J=���6/�e˪���'4��N�~�P6�w�Z�o�|��)��g�=8ƃ��[�y���l�L(R�����[�J��iẕl�j��)��oJ�!G4;����n�NI8�}q�W_(�[���X�u�����\C��u6��Su�&Q�{�-�">�5Ex���Q"Ɂȿ�Q��A��S��8��җ����9�]{�J��J\jޘOI�^����-k�׭Dd'��ea�z��`��[Q�>鳚�����қ�I�cq������'�	[�aq�"�x{o�y˭�F{�|�=���ep
��h�"�Q'�v�Ku���(�햁���o���X[�Í�&�RrK]��謐��{`3v��GɅ��;�p�/e�ɾ����Z9Ŗw��N��i���3�M݈S2��<��r`���I~�C<�:5�T���T����P ��bFf��Jb7)��yE���p�5le������G[�.aѷ�.��3�%u���R�5�×\� 8\n�ي�eS4[�/6i�(of�U:�'��)X �i����R��M�nݼ�rS�1_dy��օ��'r+��(�UW����� �0��C u3�pͺ�Iw/��6�P��R�`��Sm	��Ӽ6kd�@�5r#��m&��r����+�t!�hCf��S^�e�ADʼ9	{�h�}q
{£Cӓ��ؗ���������`�� �������X�7R�*����3���X�6���+_{rEW��[P1JVll4+��u�uT�u�9oL���{��l׋P�S�ܡ��{�.�b�oiWt(�2zVkT�6ɷ[wf!p򤰓T�h&6���H��xB���,sx�1c۫�v�{4h���ػ�˛"w]�b@�k��V׶�6�����Cv��Ӫ�=��t��cD�f�If��,mAy`��Km�L�e��u�\7����B��-�W�������j��Z����<��=M�NC�o*�qniQO�Q����9��eR�-bv�y��
�@��i/���S���H;!�ϱM��8������ksj�b94%�*�=��{Om��b��g��L1L����W]j�e�+�?��칈>��i���� �k���ki��A�ӈ\�k:�����M���_e�Ś�~Y�o<]���E�M,��\����3]k63�'��z�v�|#ۙ��P�6d��L7���ɇGv�ʣ[ɮi��cr���+�P\�[��D��S����!�p4kqn�a±.��>.!&NW^�[O�wwt5>����0�f�-�D:���x�@z�qxh�M������궿wr�Ӿǧ��CW�F���ӝX2�U�)��9�^��</����!2��BL��@>}�D#��;K�������\�|}�j��bóYn�qo՗K�W�YՓ!��P͘-i�/)l&|9i���w�m\���s�75�E�Ip+l�b��p}L��ג���Չ@,�m�	��\zY}�f�Ds.��	Ջd�0��Gy{!�:��nn`(f��z�i��#z+�S�R�H�r�6Y]�4��7{���Q}U�:ux���/���'���R����
�7ܥ�[m�9�t��x�ԈJsl��R�U����LF(ZĕK�8_d�S�#'�މψ���x;��򟻪$���Ǆ��]uNn��+�FҖ�N�I�J�o.-�5@�V�_PΎ����޽F�۵Orj3]W.���ZZ��U6���X�!3$硪5 �@��"f��,Wz��t\,�cou�[ٛ�Iu�QE�>���?b�M���=��/��쮵���l?��G~ӗ���G1ς�^�&��� q~5<\�x��Acϊ��[�b���%� [�騷2��nd�v9L\����i���¹[��d�aT�W��1�������4S��������h�y�ێ����qwI�6�%�V�3]���8E���j���� ���` f��cܡ:���vΰ�tt���ʮ�I�?q�B�����֢q�Zc|���
vA]�qۖ���(�n�*�e��l1~Y��L3������*,.s�ޱ�#uH���ĜTV�N�Sf+�k�xz���I��T������9M��ʥ��ܢ�'�.�!��h�\n�B����U>��E���ēx�v�%��K�~6+hW=b�->�2a��.SJtn�'���M �]�{0^�̆f��}�\%X��my�ּ"���y�E�S�=t�w�Ș�Rs:�b��/�;iq�О�Ǟ���j;��@���@�#�
�u�ܑ�e�����pq9&�6�T)[��#q+�����"�^1Q�ُ)��z��D,$Ox��PΛ�[�$��Iq����K/H{N��a�g+�����cn�	�>��xW��g��@~Z�J�G�mcʷ1��)���ar�Y�>�HXkd_�R�ё��ʛK,�ԣ6	�cz���$*�u/Jl���MOA�V�]{�]�W��}�~"�:9���<�ĳ#�y�	�|O��=�tUmuNtӛ���⪥����R�K�M����^���`q�sG� �9'�T�MC�9�s�K]��J���5�
oM�����ݘz�k}繾�'7�j�$�f)#�4�cJ
�R��� �`�{�7�ʷoM��5���R�z���V��x�c�����:���w����������3x i��A�4B�
��޺�y�Þ6�Х�W9�b�G��OЦУ"���W�P�}�F��Y��l�1�m��܂W�H��N�W��9	M�m��D�"�7}L]Lw᫃89Rr���E\PB�Q��7{:e^���W"sG*�خ"=��H.��[K���=�Rz���>���z&1<�Ի_���SkP��˟�}�Qy�v����Ȋ����n�+d蓪f���q�M�O5z]pq6�+UkQw GI��̢��O�61[5�l_�3(jWu-ȇ�EZ��TmB�\����*^��CG���m�R���"�3�}�~Vj�����nq��_n�r�ӹ]�a����aKG��1�P�2���W��R���3�+�R�r��ίLA��^�nJ-Z���&G^9�J��A��hK�-��>9L�㚼^%3���j7,_nDN;�mG^]9�OC��V�D�n�[Gy)+��/"�HY,~9"����5Žt�m�؊�T�3k1�z�˯8ؽԩq���P���s�F�P��������0�%k�W�*�a�^*�=�fE���.���w0��}O���;�[��-��Wp���~��xo�J�X���L�}�qV`�5�}��(��a2Jp���u�*�N��g��0���2���eSLZ��Nvw$.�K�$�L��tf��u$��{WX��@F$j	��3�����}����zTu���mڀ���_y�����*)���ޯqX�*K�P�/&e���4�M&)n���lK���36�7_� ���y��/ɨ��g&���Z��}��N�b���!�<@f�|r���w����!��!#�j�P�p�"1�(�uY(*9���V1�+#D�ݢ��a��*0Ҏt�M��ⲍ�ٍ���T�C�Eyj_x^�1泥ڃ���}��^��h[�ӓr��V�m�3r�Y�y/~������J�Z�
� �#��y��6oh��V)-�ɨw۶����}�f�uA���^;
{���Û�m�,��h��N��<�R�MRo��Ȟ֫��W�h"�Ҕ!�3"b$��}�'ƅ���R��R�o���V+���`�N�Ȍ�U�W���ix�&�c�?d<��'���V5��,��b�e׊�����:�^%拇��?f:/�¸nz[QJ��R��m@	I��䫘�lWz�OH��"8��8Z�R4.�X��fd��-\� �NOLa�������?5e�j����rFQ���F�탪e9Ӷ.K�"b�b�mN�kn�����Gs�tm�+%�J���76&�x?B��1��G�4����������	�-��99�g�ḿ^啷�|��;������b,Y�j�%ZzFF�<���m��d�27
�������(��*(ifSϟ_[������{w��#��sΘZ]t��
i�E)8�sӍ��5
3 �Fބ|^��ո�1ܠwH�se��\b�G�"���hHg�9V�<��c��ގ��_��c?�ם���JcK�\ͬ��;t���e>�D�M�oH�&(EUr{��G��C�B,�Ӊ,��-�9��Ij��=𯏱�	�x}�72}"�4�U�J屆ڎ	G7-��kܠ�`�������b����Nl&<vG�@�~y�~���Р��{"Ng;���4�;�b4j���eۑ۫�ܽ�U�\[%�N�Hx���>�"�z�Z�Q�����F/���2���yuOOe�/��Ϻʑאȍ��>͘-i��#���k�a>��0(HQ��-�Nc�Q�'b�hk[ٓ3	��t����Y1|�^'�`��+T�nAk��h�M�祜��/��SqJ�W�b=3;T���Fk�i����v����l� ����7P�qd�tܟm�e�Mڿv"���Chl0�Ӫy�	��7c'��"�fw��F�)8+� 2��V�����~_�����}>�!����y_�ن/kn�ˈ笖8���7�u�GGZ��b�a�XI\�h�'gf'��CI�ȏ5Y��33]�q�{Xo��3�Q�ϖZ�v{#4���.�ob���k�k-:}w��6t�t^&QcN�ڝ� ؛�Qn�T(�x�'~N*t��1q㾡�tn�T�L:�rvX�>�gu���7@AV�ϩ��A�G+��v�7�೴Ơ�7�c�yޓ�N`U�}#��<�YE���*EC7��"����~f���u�܈xx��Ő����CnoRm��Pl��K�;��R�aÙ��є����݇	Ք�V7�����`�Y�������hT���[�,����c���KmqF�� *w��7O��_
��$NL��n�2�3)��:¢�����yP�"���� ������3���d��=�Ct��"o�Ĳ�l�![nH�.��B��aMO˟�;�@��w��uL�ӹn�a�׽�}�czTAt�t��?n�GV-��%1��� �]e,N�1���zۺu��ϟgJ�Ks����J��U�����	2��X�	`��8n��ӱ�W67	�dn>a:N��ٹF+u��2��+zR��dLZ�NNe�ץק���kָ����f�`��k��|���}��x0L�7k��"ږʕ���g�y6C)��	�5%���`�Vl��7�N��`)j|�����aƊ9Uv6	�a�[d���G
�:���q�ꎊ�J�L�ɻ(n�GE˜�>㔞�+8�x����̒����t8*
��ܪu�.��,#OT����:���kN!������N��FI1����n^NF�خS.c�a�6�r�{���sE>t�0��ݜ�{oJ��Hnݲn�4M�,�B�\q��ѝ!U�1B�Gjv��3f�6����ß�#|���=vB1��o0*E��d��2�c��JPk.�
d	�yDnh!P9���.%�p f��j�0P7�U�Ϗ-�&�VFu�U��4�5�|��>�O�u܂�7jh-f��;:�Ӥq��2��V(B�;	�Z��ٜt#�-<�O"z,�,�$9F^��o!����#�ҟn>��$��_H�/]ΰkX4�w{;GlBF���+��c�5[ũ�P������A'm 0w��Ąs����4|���h�c#[�`�����pD#� Xa��Rp�n�X��
�����R_�d��h��}ƀ�s{�E=D��Շ�4l��CRKRS/����\���!��[2s^
��+��d������?l淟!�����Ey�p�qK۸�ذ��-ѱ�����R��,k:��v,P>���;�G5x �*�{["��uۚ[�8�]QWp��@}��1=!9����LG75��k�n@�L-\��p�8	��|�	�c4�m]�U`ږ��h6�5v��-b*��v��c���X��T�ڍl��u�٤��8�6�c:���Z�kn��X�*&f-�㦨�,E��Ů��.�i"
vŉ�l�
�C�5TQq���D�F�Mccc3D���ΝWlU=��E��N�5���֣g���#��n��ke�ƪ$���b�c���5m��%�Z�X�w=	�K�cZ�BU[��Ӷ�Z����Q;���h��IDSֈ��؊ ��1cm��Qv�E���h�1��:�bQ���PEl�0F�"-�N�A����v�ы�*�b��F�V�5]�j��6�OZ*��j-�qQ2SAAOZ("H����c�d�mT�]c����g[(� �5ݢh�f���#�F#��zh����h*��#m0]�j�����МwqS����`���4T�GX�j#�AA=�X*��"�"�("+������`��TTPƌ�[9)�f��]���F�N���>�zo*n	.��+�c�^�_�b��Ebo%�o����]�Đӄ!�dW�v�Y�^+�۱��� ��A4�E����wמ�n�o]���~�'�UOK8��)��,��b��bU~�0�����'�'V=��Z������.���o���\";��M��)W)j�O��Q�)���j��`�u����痢���5�nYw�M�re��YE���ϡA�'��F��?�R5�q�u��:��k�v"�s�`�� P��Ǯ��>j�No���k$����m��wcX���R����{�S�j�<����dEjk�!��us|2��xS����j�zi�v�����1�%�����x���f{S��������=y,���$��d'��R�K�i>����2'duD9���]R�4�`a�#\*��.z\��vMu���>��WMf�ҋ�/��3{��.Zd;뙹�hD����;N�W#��	H�)��^�=���p�q�Q�6���>�R)�޾2a�R�.��k9�*6v�i�]��Ǽu��T%Y�;IC~�xD �橅�UJq+�h�+���r��<�/P��Qa��4'�[>{�L�5{|Օ�|��!�Ƴ�O�o�(��ec��~#�d�@8/�Ex��]%|�A�y��,R�p�2��p����Y�
LZ9��4����6������]��-�:A�.�O���vQ<)�.�+3�s�k/r�9C<HT�Y���24��A��u}e��		��.���%��=��_���f�)�*�$�*;��྾�_G�o����=���<���`��N7F�5,��bu���@�R�D�oTz"̊�u��m�GA읾��>��`�,��g�P�!�c�'N'q�Ғ�hB�N)E	��1Z#���l�>�>W��t��(.�XE���X��	f�2wk�݆����ra��`�:6��k�ر�8�����]eڑ��HLG�+���	�9����1�&��FU�`�^��lin�<ߘ8�z��,�͊k�|}��5F��w	?xK�8���Ѳ���S%�R۷{�׍��a�@WFP�R�u�ת)��r�>-ZԾ�z�����ص�N�L�G��m�픧��|������z��o�e
�S�%�Y1>P캼�{*�TK3+���R��"���}4���S8�����ƛ5���*�ye_]x�a[�/�e�r+X-��t�nB5Q��܎g���Eٸ]��zMs���F�'�O�7����`I݄F�L�Ӗq����{6���Y[/C]�4����K�Թ���4_��~�]0�����'�lZ��H�^��nۿ�.�`��%�N�N��g{*(q`�5��n�򃭘�3#�D~j��>��K���P��/��pW��y�j��]�>�g+�������g�
`\H<�����}:��ە5F�#�ws�Q��n����|����׻ϱ����&j����0��9�v*�ֲ����ˎ�=�?ef܌ϡ�7��$��k�b��-1O�Z�QY�R�{�uLu�+�]��s7ju�9y�ˋ��iY+_�(�P���J�\'�&㚤3ѝ��OxZF�ʻ49����k��q�5����]8E}ݱ�z�;D�TW����&K�`��������o	�1�1]��{�1�͉j��hQ<�S�;ө�Z��.���#G݆�a�D�S��eޛ"T��P���3DZM�n`����cy����LwQoP$ⱹ�>=Z�g��7m�x/:�����YLy,q;E���A��`�5�A��>5�Q'��'�I�6��4�F��N��6����������1���_�'ڍ2�oʂ��;�pG�EAX��=.�|��+�� ;�s�����[ڶ�T��_��<~��dT��+���{����&&�y+�\,�3P+**��؛�0�1(s�:T[N��N��;��<D�Sl}�m���5����ޑ{з�l�33n��U&:z���yQ���j��:e�IB��T��6�P3�Y��l�C���~��%2Wj�yZ Gmٕ��M��a�x�V����A�S(�Xe�q�%���������������Y�7@N�t^M�ݵݏB>f�G��q��F�}��Uw�"���H3:����+8ʾ�r�-�{\���fm�R�p�Rg��=����}�}��`� y�x3��Y��ɴ���uo�PjKP�	�}S4���nj�Bm�R1��WB�����E�U�q�q��ޮ��mp��Th�s���*o��1q��3.z�>W��,���I�M�F�4c<`�{�����o�5����F��W�����C����`5��QAu��Hթ��x�Z��|�$�gl�~ZUc��
��x���+83n�c��ȵ���*��m);��c���Y�H;��^s���S�3�$�
�ŷʹ���C��|i�T2�R�G��mH�� �א���ig�S�`]�^*V�5ʀa�V1�輼nOQ\4{[N�`]w�%j�	P���k��{�	�D����	ts��ԃ�LW,SlT�Y��N���9k�א�, �>�l݁�|D�F��t�և�<�_6#r��*9��m���]��{�'����
����M���֐#w���;��~��a���W �{��N��x)����I�~�dt� ����`(�/�O�1^�1��|�k�R��e����N���Na	Bj8��<K鰼�ǜZ��x:������q���bcZ:ҥS��)�+�"�����7+m庋q5���-s�
�M�i�2ei�]���[��Nq�����:���;cJ\Ӏ)�N쳫� E�X3 d[˨������ $|H��<�=��x3x3fSc��w�kc��p3�13�����"LקMKC�P!�\��m�`���!��f��S c~J��38ȯ�_��t�V���L�mf��7r��ي7�� �#ͣy)�bs��~�R�[S�󩜪7�&Qhd$��T���C���dv�i��;N�e��D�⦣�ob���I͇����1�Q\%�k�KĔo�+139�-�%���q�����I�h��W)fǫnԈ)H�n�Jt�N������}��?p��6�bLO9O�,}� S�#$_tO՚�&&�]�2�P�U":r�ԭ�����5�~=����M���Z�5v�+�zE�8"����ʺ�p�Ƀ��[)�kA:�Z�(�����|��#�3D�aVǭ�~o�HƦ�����T�����I�C�,W�H��&�����|���-���=�N��Vl;*���[��R�6\�����]n%g�vB9"�N�P�=Ѫ�8�ҥs�*-99���f'������۸.��ĹП�k���
xD�c����xK�䲌gt鯖�EBi/��P%��a�t.�����s-e��;/��������2��7r��\�i��g0��炋r���mC�s�@V�ō����W2���N������d���|'kga���̵Z�N�(��V�fTX��!P�����H'�t]�U��{��"�_��x�j�i(�A�i{��1	ꛫ��?ec��h�p�^=K�C���O��yΎ�źrj+fvV-薹��ϴ��|��}Р�m�Qۏ1�,bHFB�@��be�����P>�{�Q��{������vN��X ev�וc��=�[u�	]c�������V��b�Uy(᷇��}">�uRrX���ux�崕�����������=��6]�
�6>�J���[�a�ڏa]UwԌWSN�[���%ƥ�Ϟ���Y3�Ɣd[+�gҪ��q���8��I�Ll�-:�̚��,�ܤMk�`ֲE��k=!��2�zA���w���\�Q�Ƌ�x<\{���8��LsP9Ҳ���L.!~u�D�znc�6�^����~/���g"�U��Lpy����P݋��zY=���P�J>�b#��!ã�������xaEu�RmY��7s���r͎�!�=�,��Mt����h�)U�)��^�ж+C�?*7֪pTAedt!{�UK�?�`�|`��7_���s���YP���(w�Qv�MH^Sܩњ�>1g��6������_��>ٶ2FM�����7^8��ǧ����ꏱ�]߰?��B�D����N�I�@�v�β��:�v��u�������ȸpܭ�))�+�����YC��K�����Y(���B��V3?��{�`��0�ݬ�qe�@ed�ϼ(E�ȹ�a!'^�t ��j)>�K(V߳��I���P2Z����Kš��]}zf�1j���3�Hx�f��E�&5���5�s�Z�R~�YB���qP��m^��;���OoeR��p�y�����1�L���,�E��-B:M��es�Q�ݰ��<OK��WMZ���s�.̡�$�q�@yRB*a�{ЭH���O�G�P/��iT�}|�|��˝6��K�7��>�^)��g�S�R9c`���75��x�1���S�.uO֢�R�����
��fg�%�t7�k
�R���)��F����B?�+s�Svr~����R���J����J�m|��%���Wʌ8�6����𿻫gǻ����Vk�X�a!d�Z�<}��Y��˪�h�z������-^0�̿�gd�R�moT'�O1�zGY��w]^9�y̷����u�;�<L���lg�H&纤D?j��\���G<��V��[<����KЌP���ک30%��l߻��E��A��`���>""/Ʋ�$��=8g^��
�7�u;�/�~'�Ƿjۭ�qr1-�%)� ��#.c]����p�W��33V��W ���=�Ks��ƹT]��7Z��r�b8�5���d�.P]ڨ��N�Zr~⏛�IxV���{xhK*N5NJVs��v�z��S�Mn�)c��,�#�/�(R����R���O4��-�=RZ�Зc^��T ��k����z��G���V]��w^��mC�y{E��Mu�����B���a1�S�u��q�^[-����S����Ÿ�̭Z�u�H��:��C����rX�[�}9���$�9�_�?D���*>�V��VΫw���UT!Z���(ME���>2���v�k�N��A�8G�3u�6�P3�Y�+�z��x��)��z;ngV_�|S��2i��Sa�'$^���y�8��m������"!��f踶 �o\��j����Q��(�hd�S�oG�蟴��F�gA噽:�HʚsR��[�����{��{k�fX�ŵ�-��S�=ڄ�ц�Q�cA��6)O�"avyz.N�6t���rX!�gYn%Tȹ��]QDh�wpāV�S��������Ǳ沱ӕ����S�YԆ+ݻB�3�̽���,
�Mڔ�b���ɜ�Ƣ���8�b,y��НŬʩ�p�т�@-���"�ҮNƢ��pK@ގ��B7�W�,c�a��v�n��?�d]y���J�v�v��NB��`�� ߪx�� Z��j���6#|�s����)P�7�p��U�m?ؓ=�'j�7q�;��� a/m�}��;q�=�r�����:]��3N��pYK"�8�U�4�u�����?�|�dG��ɲ����z��~�^DH�*�=����H�x�D��4ۿ]��U^/�7�����$Ϙ�o�ل���>ʘ������ٽ}���ֹ'��'=ޒ���[랳���1z*��"��df0��j�Qy�*y��>l�M0�����Ǟ�:\�(L�!]yڏL�`%�]���|��z�q֦N+ճ���Q����M���ל���0]Π�	���>g�[<���.'��?f�-i���[pS���b�-=ڇO�J͈%�u���>�����4�ħ��C(!!�V���Dy�oX�d��h��1'*�Q��g�9,�T��}��5�����H����f�(n�SAf���1(�L�MI�W�֭VZ^<5�.����y@�vN_�}��U-Cw�;E%(6�v�OX�2��/35}�m�X�zˢ��K�q��HLG�� ˧��%��I�w��1�G��f��L��7��}�ʽ^��{p��R��R�j����,MbM43W���A���p���]� �y<��R�}�)�*<��?E}I�Gd���lм��/]�_3�;�R�~����eq6i27���ܺ���<��7��v��K�5�m4������0�����s���H�;�iE�*mA��|��f��)\���&��|3��_�fy�옎��Ǽ�^=�rg��u̟wz<fo��f)��%F���~��y8̎�:N�G.��������y��/vA~xV�;���}����%�BJ���?5��]�{^N�|�(����{UZ�`I����)iy��R�p
Ό"~�R��%Q��g���V�*�˗e�f�I������%�G�n���o�)����>z�/H��߼�ɂ���2��E���ws�m^�vn���kb�m�g���p�o�eF��Bu�X�5�ز����0�}�Θ1�\M�uI�6Y�uʝ��F�S�F,GF��r�遉 |E�]�0�b�!G-�rD��ꥧ��4ѹ��O}n�2��]/yP[�[{�_�EBU�I#y�~˛!r�W;q���)�3�N}p��Ü~��|]W>��J��lyl�B{W�E-��l���d�d����ZY���y�-��PΙ�\�K��+���F�XD2��,����,����Z���(�^��R�{���&��ǒ'{R0z8�8�r=�Gr��� ���cN�L�||������}>�O�����a�~����ϳ�[�+���y���
Y�3�b�-�1��5N+廊w�O��j��Z6+ɟ ��36�'����n��ߎ.����71Z��KD\![|�X�Xn�����n���ݐӴ�uD�dA��E���3�Դ�WbD�/��d��	����NF��o��.�u��K��0�b��,؜y�<���>��t�������a��|���'����X����Ǫ{��[ɪb�L����p4�	vh���We���=�}�[\.N�uW^��"2ht1;J�7��b�^�+�u�����cyr�#�]p��fMʳ����-s,���P;�D�6�\��af��!V�6��9��4�9�,�R�i����7�����>���ʤ��{���,`��g��P ��sȹɼ�
$|{��Z E���V��%��9/U�×�@�3{x�(-��gx�R�o�K����zs�4�)�[�W�R�m��{藜���	�R~�m�y��s^�C�L��y<8F� �O=�uPxg���>m��H	�ܓ��'3Q�$:&��v]���WQ� �WϨrw�s��r �ӛ��7��a�(�,���^3B��G��x�	xx�5���P��H����u�5���Ԝ��k�����Pn���ږr7]��� ��Q:��!]D-���9Ai@7p���e��T�g�b嫮W��b�lZW#m��D3�NF5	��ئs��ӓ7w\z>{ �9=*�Ol�[:�/_�L�
n���gK��).>'b�y�'ˍL׹%�`�K����6�*0���!��.��0_M�m�k�ɛ0u��-�-1���74�dzV���3O�����r)���|G6��s��M�7���e��������a����*H�;�b�k�b�sp���$}�qy�����u�w@֨#�D�8��u��ف	�@2�xZ0Mbz5����=�-��r��ҦU�������f��h=��v\���0r�]l��7u.tM�ug�Һo����	�Ç��;q�;y��r:��d���U��6��=±���@���` �Ck��R0�V��|���Ʃ})ɗ���*�z���3w��(*�R#L��w�����kf�<Vx��}��l�X�VeJmA��n��ybP'�"�xL��$�+Uʋ%��ڲ��#�I 'U�� ��7��`�WN�B1y���1ۛ5{�-*R��l�3��9B�j��Ձ8�:���S�n>v�ge��F)�1z3Ǹ^"5�����;�L91oP�7�0�邵�c$�J�ä���/e5���8��������{Et�8)6�`n�(fл+&�MdZ><�������ݾOٶG0��,;juu�kX�ķ�WT�@uoK^�'���|y^p�>�ԖG15�@-�ޝ��[tD���S�(h�d��@#��	�Eժ_�A�����P��ڠ������v���٦�2t:"(���v�]��Ӣ�(��U���� ��i��th)���F��b;�j ""���N�m��J��]�(��SkT4��D]&�����h��4Nڪ�)�������4t�kX�H�6�T1SLu�N��`���&��b*h)��DAL�����1Mv�A���j(:tPEIDm����������؊�cUA֪&B��h�"" �i"*���*���kOll�h���cEPDҕA1EQ7[�����{:�*5����h��)�(�d� ����-$�DQT�ԔWcwM-%1�h4�4�*튩�jb!����tݓ\Hb[��b"Z(�d����Aݻ��!���RQU�6�ެ%7SEG��WH�.ٻ�:4�l�R���]�a�Z�����^��8��)�G�v��0�F��N��#2��L��sV�CS�[��{��j�{��P��`���H�׶9�Z+��5�>
(Lkׇ<��*ؿ
0-����=�ѽ�$~����y�_p�r>F�du�ͮ�J-�����L���|�����1P�`8�� 8ts����u�C�t�X��=1ᜍ܉��G����=�I򟳃�`�Vs��:<ڢa�^@{2.���7&L?L�ԥ�����,��٢������S'B�<�j �zNt5>贖s�����j_S�Jf*���؋d�U�#��S�B�F���o>�Sl(j��B�e^�3e���ʱ�5Kje�@�Jmm�_FQ}�8���.��_R�	L����Eq�`f>=��G/`���S��rT9���-��߼�e֕�����}�m���gŚ�m^����MQk�Ž:Z!,�l�1s�f:��3�l^=z�܏T�׮a#�L�"������lh7\d3Dj��z&��֑�v���a�����z"99�'�n�8��f��rg2b�?6R��� 5ǱH���)�Ʊ�;�1b�L��(t��*�u��f���;3����w�(}k�����'�
�D��t��#��i>�� ���	���\jPͤ1���{^Ga�M��ea�9u������Hɓb{x�qu��ht��� |��q�鸧.�V��3�kr�S@J�1�9YS����t��SQ�:Б̭�F|��G2t��OI�v��
P��)z��ew^��k�Q�R��Yc�7�c,��U�|hÊ-W0���K�z�	�Y��Z+�6q�� ̦�:Kt�P=��,�O�M��$D%�br��_��^m
��R����}>���,H�]��O�:��u�rk��Z ��0��$�>�ȇ��E2�Gm����cp%�"b���������g?���gu���) }�ɬ�
� 0�k&�O1�u*�T%���k�y�	K��Z\Vev��v���kdB;8�>ԉ�l��h�'�A�>�����I[D��r������w*,]� ��`g3�&�O���:�]���o�?��3.�=5Х�a6��u�ה��҇��W�|���F��R�@k��r�ي�؟���5�K�yyw_��9d�7�L���{'��V)�G���Z�Ât����W���"��7"n�VC�Mƞ�5�Y �v�6���W�����@����K�ƆQ54s��F�4G"�oB��)x4
}Z*�����]���'ZEW��D>J�2d��'���UO߃���H��A�ۋ/zj�
���'/�a?�qZνos{f�3��ak���ť������S�s3�u�!`J���qeZ��,�<r�=&����C���k��6o[�� ��Y:�Խ��w���-�L�v�ɓ����v�p4�{�9IȄ��X��,�F���ߤ޹�������w߿F�%M�c~!�������g�PdPY�n��؊ar����9r�^��a}�e�T�9�Sm�k+QQ�0$U���+/�P��z+o����T�L?A��K�F�wظ�fd�?<��T��X*�7v"����y��[y.'_np�*!6t֎���xy�K�v-~�8�6����E�S�ؼ��:�ڒ���.���Fo�p�g+;St���~4��������1��dۃ���c/u�{��~\�Vw�t�zX�vM8��&tD��Ι�q|ň+|�Ȅ���m묪m����y+��=�9v�f7Ref�2[
N!r��6���� 5�GǞj��F.2!A�+м*��6�N�ieY��[x�s���Aeyډ���4���8u!�?,�yv��HmW�MEcߝ.��s��*��yC���Ybr�͏�ʑ��ȍ��3fZg�<�l��z���9?Rk��٣Y���5��H���\%k|3�d�|mc�K�
�'V% � ���z!��۠����ѧ>H�H�[!�u��R� �d+�yƝݓ"�7;��"�ι���-���:p�����z���/�'h:a���7��.j�y<�����%���^�R��DIF����q��\�b�XC@��#W�:P��;�$���E�	��ץ����!}�nZ7�3�-�ݽ�َ3��#��Eqs{7����TUO�b�u�;�<߷��ņx�t<I��x�X�o�����}���spL����I��;�9�˱�]&Τ��s�9�tod�R�����}!��¶(����>� MG���m���q
��Y<��譝|�7����2}�%%�^�ɦ�մ�$b�m�a��U�^��
����PѶ�Ե;�y������ �:��y�$����&�'*�m-�k�U[/-^��)���V+|OwU��Y�y>��R9#3�9�HU�1+��x����_#Bۓ�5W�j����/����۱���e����o9J���}k�YфN>�.,Ī<�TZ~9᪅���U�mb���U�ym�r�B�z>����q/���ҫ�F��~���m�mf�85�3�j]�S�;�e��A�Kht+�����!��'ئ���<j}��z���R�T�m�;�����[6�K�e�a���AGlq�[�|��A����@hO�ǒ�r�ae^���}�a東y^�׮�n��*c�3RN&�gL�S�/�̪����]f���¶�@ZG%i��c�+6�&t���<�u��@���k��%��W��5�qJz�Wcs\e4�{K�'oHE��o+�45�OW*�ڕ����a"�D�ty1���d�J�Q(
�)q�+�Ȧ�`��q����'c���1�D�~���R�l��&�-�n�k�/:��=s�O~%Ra��y�=zU�j𿮞����|�����֩�x���3�q>���'���է�rc��v�`��N7<��@{�I�ǩڻ��)�#n�k틾�]�D,C!��Ȼ���%�C�sY��45P�'��c�w�у�+����n�����ȭ[��C�#%퐘>G�F�b����lc��k���N;���%�#b��K{��)΂hި�I|�%�(?*
�ľ~"�:9�v�ގ�8���\K@^�*�U�_��'�BfOC��x\@�����ߓ�j��oέ찣f�e8I�EC�3�&���.��j\*�-��eIB�)�l/Uk�ϹM��O�C��G��0B��N��.��F0�`v�s{:�Ծ�]�Q��=��A�K�/)�+�'yV������O��uM��'�kk~�h��.��+)}s��V�^���&��|{�^#�;.�/�ZE�q��7��u�I.���^{\�% cŜ�ı�,97{-����}�Y�6x�o�\�'� �U��Ck4��y��h�UL=M����=J�I���sS�gOkP��#�V]��2�$U)+.�V�r��ʽ�N�'�0��f��ɯ>듽B8��
����4^C���E��M��C�][�b�<t���N�:�Xl�۟FJ�t�⃛�x��t����X�^=Y�6�;[^��qL��
���mA	θ��R�i�P�mG����̇r�/~�f�ZE7k�%>���rg2b���ށ��֡��޴�U�����3���Xk�Z�o����L$��ܟ����~�m��k����!�2�sU�aTA�75B�B�~˝��^7�㚦�b��_B�чr�s�E9�a8���Z��\$���ʋ��؇�֊���X9ʦ#_��L�2������<�K�����j;�m!A��"�����ݛv�G��2֮�A��<$� ��؛^�z��?gQoi8�dA�F�~��b�i��ϻT>�xULd���E�Ɓ[?#�|��ax�MD���6��u����Mm���L͌V�^&5���4[蝘�v[�7��(�R'.��ޯ/gV��o�>Y�]��28�Q��\z+/)�7�d�u�¤n�D�uOP�]^GX��>�_P��׷�~c&Ft6{?'Y��k���yp����Vm��������q���C�\%�mJI���9|xb�xj�@e׏/0\ܛM3���ڥr��K2M�5	so���7���a�,�ւhM��J��-�����ŕp�5lG>�~���o�+��[�űYI-���x
�U�=[HH*m�O�M�'��~�����P�I�cD�ͺ�����"��&%�ۡj�Nn�4�^�cA(A���$M���Ѹ��N�d�A�7��7z5cAv�������+���(<>���n����g)��c䵞W��d��5�2u�mʞ>�
��$]q��dذ���D<S�oe��M{zx���3.#�8lu�^l�h}x8�C�K'��4˯c{������_���ϩZv�����3S����3Uze�:꾷�]3�]	ׁ�0by�wL�[�U2.sڦۨZ��y۶'궺\�d���S��|&f��y5<�4(���_՞�{cqW�c�XE|fa�M�m����Ի�t6���RT�}3����n�>M `:}����!�E�9�E>:�O�`.�n�w�Bj5��|&6���#qe9e*��P���t6�az��z�_M�~��ۮC����`��l�ab�Q{L�۶��1m+�Lv(�:>3��֔1bZ� DBm�2۸��7�9gre�e*�jE��=����*ݔY4V%p#{�/Nh����7:�2'���7I��M��^t��:�z`\�V/[��bm���>i>/�b7�����G�-=���,�('Ɍf�
9����ƞ3&@JN�f����Z�t� ���C;)a;�i�Rop�g%��S��׌c�#�cN�4t�p�F�k�Gɏ��y�@�����fY��#bf���]ʅ��Q�բV�yg=H�D�Ll��Go��兾g4��\��5
O���������00��n՜9��_�j:}Rgdq��O��4�{�啧�W
�������2/�n�60㝭E�������� υU��ܤ��w������Ǡّ
���h�k����8�6�Ȁ�q��>�e�Hx����&�׬�{wv�`sj�2U��\xfy,��]xf��Q�H�ޤ��2}��lì��&w�ѓ��Dk�`�:GD�M�/�O%!����ō�/�,f��S;�;Ǽ�vmg<qfj1��m�M��˚%�`j�
�X�A�VeV,w�M��2�3�mZ�b�&1y�v���0�oHx�R9����v�X|0����[A,�����\���K��[���`��Q��v�oUg.����O;��<	6����Ɍ��ީ�Pw%����8B�g+�4�3<�hi�˴/UY��|���� �[�^�MzC�|*"ojt���ڒi�b��d���X��G���*7V�9iͺ��b*;[��PW@Zʳll�	+?3~�����s��BM�|���Ԟ���IQ�`�r���%ܖ��䞪�?�{�-������wf!oiG����6�d0�4KHz~�/��#:��݋=�4��)����e�e��p�4���o24&�[���\ؒ�f��ʪ��~�h@�H�9�a�zi�s֌� N
�<:d�s7w�`�ƪ�ΌI����~P��r��_o����D��+U���R��1z��@��T;���+1�OO�ֶ�Mrf0#���M.2m���߳}F8;u41��`����;��,��WAgds2ɭ�K#՝c{{�� ����w�`�m��F +2,��U��'7�y� !���5�f�=��9��y~����:̗��z��2>Q3�dU��+d;Nv>����|z+1!�y�5��H��pޞV�zL�K��b��U�P��K³���ݵ����e��}�m9<-w4Ehv���ًQ�^�e
I5^�R��u�իӨI���e%:�=�ي����/��{�.�S��;j�۸��>=X�=CXa8�&Q������yg�46��x�&��Vmbw#��f%C��W�-�ź�I�B�y*v�.�jmL��(s�mkL!�g���t������s>�W}x�.���#'J��Ռ��T��[b��i7�?;�f�~Dw�����j8�=P*'gJ[^�A<ғ�	9[�_�8zCߙ�^���m�0����.�U���Ao���YCp��PV��1��"{w:qu�H$���
[�k��m�	�d=j����Y۰�WI��̍%�a�y"V�@�[��cȼcB�aM� ��e1R���q�O�雎���������г%t�G6������g���G`8��r�<��Jh3��t��W�ߎ��{|� M"�>z����w'��B<:1���l�Q���ӳ�����C���͎�j�Ev�����J�sݱ��Y�`���7�o�YP?�@4>�C����H���gR{�\���>�g�����|�~�����yz��"��8u4L*����^5�e+��o;��a��
<��[�1�N��W����'3W2V�s��V] �5�6Q��Gs��T�4�(�CrVJ�\�n���-�>\�z,�ж��<g/�5M˦���1�o!Û��iX��6���\�r��aJ�����ɚ	~�+O�uo��W&z�+j�&����]���f�j���u��]b^L{{ې�9�U��y-m=6��\�hK���(cF�Z�LXf׃�r�l�r��
�УY�'N|5�y�. �%�Z��3�ݕ��Z�߸�i�X1]��Yjv�W�ۭ"/�Hqh��PR�������ԈZXUhV�D�<a�ΖT��nT� ����Y��[{�j1�*�p������i����Y������L�=�oyf<G-E2c��d��j�X���D�ݲv�؍W2�ǰG�N�̀���2^;]ڞK�����<��Xp��:U���v�t��I�]���sw&P=�f�O-�5�R�lU����-�̬[y����o9l�{;h����.��WN���c����X�*�.�]4͌�I�n��@T�`H�IwYn�3h�s�@wV�F�2�W)>��©>�J�E:�U��=��2 �3�Ǜ[y�?{�=RJ�2ܼ�,dRĩ�*U*��bIo%��D���q�=�5�ό�_��e�s��9�ݗ��A,i���%>�[y�n
�V����w��Ė�#�fZ�+s[�SUs��2и][��(�yU�5��?����c�O#���b筯sc�pZ?w�� HAN+a�����%Y��@��H�Z��w��GR�{�8�:�Z}�G�Tf��7��������Έ-}�b�{����Hߖ�&�p������vT�'[(��U馻��W[�gY�p���q��k�$�L,��!y�6�&�H��2�T�,2*��ׂV�)^��.u��p��pԋ���T��;{�I�btt=��GV3ྼ�a�@��D?¬fe*lW<�Z���W9�U�/N-�u�h�O���L�U�G�-.ӛ������Q:�*�2e���i��'���zv�r���}s���0ɦ)j<��:*������V�A8v�+�\��k�ij�Eb���E"r�Iέ�W�o8�;"7VҸ�q���%�5���������\�-��$)��^�!������cy�:��z8���1��-�����[9aL>
��Ҳ����K�o����

n�\O���ë��G��m� ~=pP��5�j��!���5�1�I�Enŏ��X}��e��zb�����C�EUh4�^;g@����5ޭ�;8N1�ѓ�z��Ʋ�^�ES�[�w�]4;���O	9X˝IWA_d48���M39��wU�S��]��zm|(�4^q��35OVF�r�$���˃�\�.PV��	�#+^{�*/�_p�9T1�{F�}F��c���U=�^v�r�X^�9��E���%�������{	܃��}����I� j���B��)Jh�
�����!��+Q1PSClh���h
�j*�u�$
��l�cZt��lAKL�Q�RБPQ	DAT4�l�%Du�u�C��"����A�S@PSEm�61!Q@P�TC�@�STհS��MƵ�����
����!(�LAlS��ӵ�� �hJӶ	I�ДU%Q0PRi4QAT�F�SKT豢@�-�E5Ui4�AI�W�uUt���*X��F6���hГRRP�Qk5ACKLUD�DV6���Й�H���ET4PSIT:	*�-�Z)&�&"�{b��Ɗ�i�֐���¾��W����э�x�՘rھJ��.�D]��	o�P��lڼX:�E$�QvA�#y���l�7�����̽02P̔���y+ߧ��|[
�[�[����	ZgI�N��D�C��R"��M���T�4�GNH�W���v��bSo����Q��m���ϣO]L�̳�z}�ي��4���0y�?^��!Ƹd^b[zFSO4���e�	2,��l��v�gn���;�R� ��\���2�:�����_���zv��R�D�2{2�׻Ŏ6���X�r��4��kܝ�B�K�l�M���c����*@��t,���ښ���	���R���Wq��5C��d^I��͵�F%C�GToѮ��|���M�z�e7m��5_?:�����}S�5cL�9�a���$����wZyC�7A��=6�� ��Ec�N��J�I���[EfVB{�pU�L�����<;K�A���i�z֥�/E���ht$R�����hݪ �̚��G�z	�.�֮D��Ѿ�Qİc�Z��*Gy.���kx\��K�S�I������u�稬��t4�����Ќ���\��[X�y/����R�-�4u��^�}�.��rL��K����Ju�tK�d���}N�QӮ��l34�k^���ɹJa2��6�]���*VJ�E,�x�X���쳋)&�x�[�z/�c⭵6ߠ���;�wYD.<�M���j��ះ��V'�7�B�b�	������Ř�-�G�4'St��(~�o�i,���I�};�fb�\��T�7�{�����a�}�z����ʁU�9�ʟn:��f���^z҅Ew,�:p)	k�ٺ�C�*�7a$��j|����}�{9��*s����O9�&�=ŭ�o��Ϙ������s�S�7޴���/N��}?��z�uϫ�`g���ޙa�j1�����*�����mH �6o}�FJ�n�=~c|���,تZ��B���C�у���k�u#Y��-(Ӑ�ޑb����=�}�;������F��S��4ђ��\�XN٬L��Ns��1�4��ԌV��3�����zΉ��M���;	��W�<�~��l�d
�%��+8.�۶�7���2o?ք�l������Ke�4�o�7�^���lR����5�d� �Rk�b ����gJ���/����bU��i������1t��y;����p�@)t�l�yY��$4����$�^Y�u���z>�|Ӷgf����L��\	˩2�OMb�:Er	�$�$�w+w�\���o�h��UD�V����ϊ��S� bK(�
�-J�J�+ĭ��[^K�\���z�7��wMWV�M�+��ҹe��΅y�d�2MYU�̱�2��m�Q+�*����xm� 2�Mw�)�W����D�xM�.2�t��x�BW}�2��'|{��b�}Y��)�@�ϯ��p�)��?h��{�w�&�u�i�c+u,�}ׄA���όV��{UH8XTQj0&:���g����K4����)r�7n�G'�[Dɹe��Tc�����k�h�G��O�iټ��eL��&.3�q]�1;K�$v3D�Ĵt�\���<NUt�߳��F}�ק�oMWr+mo:�[�@��n��!�}_A�q/y9B ��n1J�B��C ���x�v�o%��mU�h8Bc>P^�2K��68��%9���)RwQ�N���0��ѭYΤ��<ZjÃ��s�f�-��+4uܛ��:�N�5У{��ӧ�z���^�go�K��1��j����
�0�� 2=";Q���ǺUhu`��_%F? �3n;r����oS���q�y�+p��W# v������]qm/b;�q��g8�9m^:�}��y��ahZ=�Y>���%�׬�4S��~�������p���K��m|��tG*<�/���?�O�~;u���z�N������e����D�*�Kd]Z������C4�J�#��^Ǔ��a1�؇5]OU���7̽	��>��YU���nLH�mz�c�4��Ռ�&!�-:)����lMd"h����9py�w��E<��T����#�34oV�3�:�_�+�dY���L�Ԟ�\��ʹ�G��_�ro?�����e~]-�q���j����+5T�ѷSx˥��ic�ٖC���e+���i�b�=Y�\_�d�8J]�m*U�6�V�31�f��9gu#�Gv�u�����mbzs������y>bDK�^�X���ԃ���f�-����QXmv���ޮ�<|�eOz(N�͊�ݬƝ��s��;Z�Zb(�V,܉i�n/�`0ּ�Z�&�ASW�qWM��PnZ�.����l�w�����~=�e*g�l���H�����J�"/�e�)��� :���t�/��ͻ�o���+y]Av�������	3.Y<���v���ٕ䷦��ɠQ<���Z�'��p1Sٍ̙���k	ڬ�$O8�T$w�<w����u	큸�qI�Y3��l�Lds��dt�渟t�����Z��E�X�����$)��(.�+W��π��v���eY��{J���k�!7������[h��R�J�?Nb�٫�{/��}B�P��C�d�aU�-�^��H�ÁɹK�܈H�����q7������;�]� ڱg7Ϲ�[- �%+S��Q�8�8뽈�hʺ�=m����m׏B�a6+aO�^F��N�:lÎ�C6�;]y]Y2w{*FE�Z�\g̪`����ⶤ
�&�]�u���,�1����I�a�B��7[1/�N��6�N�z��rw}/�/{�ɗ�8n��^��ʸW�#t�-�ˬ;;|�B�F���Ṋ6%�8�ʡf�4�ʻ;H�ۘ ݹ�$��7��m�y�����H�F����Y����ާS�M<lSIH��4経s;��5�1)^m'�y�:�U�KdrhjƵ.���d=�7*�=ɺW61s\�׋�s}�c�N�>���w���7�u(9D�Ү�Ӏb�{Dț	�{��~ʫ�k��W)ֵ��{��}	e�*��5K
̅�J��.��R�Nx�,b�n�3`���z�)����.� U.�	V�3Mb�Z������e��Ï\E��^�QS���S�Y>�Q��<��ܴ�3o0��vi}�g�2���"5 3�JK:�����.�fl��D-����}�o��}*�nAx�ټ�]y�����?fO�G��͹e��y�9A�x�*e���q�XT�Ï���sNE�k��?����Z-���d>�e��^��
�����QN]�¨	����|�p7��&��#=�����og)����9��3�	a���>ISW����n�X1�)�����[�H�{-|Ȣ2��L|�g���D\EN����/���
���![:@�<M��0�$��ok���Hh1�f#���n`:�u�L&$y�FVk���f��R�ōӔ��{���^�L��A�7��V�K�D,M2��y>���r�b�������״s�'�gW�&�b5�/�`�Y�G��d��Y�{\0�yH�&�R�1�Q�'�������7���M�Z��rH�7ъ�AY�Rt���6/X�ƲxX��SN˹߷_���[\�*�j��������b]������+������Q �uX��7�H����er�/:WV�B���ȝ9<��_����9�K�}}�E*�WjF#=B���
C$��S,�n�KY��1ӽ�3��y�T�������,a5:U�^�UZ���r�VOj�8ƻ�2���i���{M^<��<�W�4�<�f� �
�ݩmfN�[э&F]:Zl^f�f�^'2���5]���4�b14\qb��$߈���&� �7��{6�p��j���mr��;�!��k�� �p�=����+K���9�k��<sZ�r��\�1�~T҃;�T�/)���e{Ko���#0��E=*�jN��e��ڠB��@�H/|D�p����Ҧ���6�%�1k��oc\ݨ��+>M��y����5��{_�x>v1��j׃����D×e���w5m��OfP�����
}'3B=y��F�B�����~�݌�L�Ml�ص��h��*Gt�7�4�8��Q���K9���ȿÎ���a��t��	n{z�v���%��$T�!Ӆm-rv:���[uA��osM�t�@��{#���e�ۙ��8��-n��Gv޳���Bk��뚍�Ɏ��R}��%�8b�Dv�@d��d�Z�&��:�寳i�b�/�#�dq���1��ͼ�b`���%O��8�p�-���p����[^ꖁ���2�s�9�l2��wY��6Ғ��=�Q��V'�VPs)���[���T��Si��S�sC�s��97T�`��B������
9�ϼ��$���	P�5K��c�8kF�Lm��̾>�	���+���ʑU�X�&���"FN�6�J4V=7iQ�*�*�yZn�q��3�]����!��E0vͭ�%��ql�D"\��q��آ�F�k��n�қ���wA<��P�)2|� ��T͜��J�B."9M�Y�L��V%f��P�g������XC�����D�u��Y0s�H
��{�l�=���^��!���7��d9��Ow\Y��>�S�#m8O+lĝj"򧻭N�;�Kl5T���%�:� ^���^Ѷ�3u���P��Y ���Y�Sx˧�wic��W=Қ���ϳxe<#�2_vz��w8����Տ�E�������1�7��{�cG|���ue��j�=m�nH���5��]ݞK�Q�~7s�����v�z�I��k���j�˵�% �\�������.�#��>�+�{)`�q��Qgb�a-�ս� �t���z'�b�˷mͽO	}e��}�;nk��S�6���^0[���u�{cۈ�m�AMݐ�T��;ϝw�}��9�<����ֱ���1�&�}CK�ˑ����i�����	Uĭ��E�iAc1�{:���_���G�T�3u�Q9%�k��P�����쨰CG35�G|�zs���o��P���L��};2$��?lCB�6�fϽ��l��������"ρ���^t��f^DXW:��N��I�K�=���ف�y��ĺ�oK��&
e�M˘����yi��'˚�9���b�18�U�G�N��7�;m �{�A����G[i���)�U:�!�����z��D5�=�"ڱd�gs���7�3r�}�փ�-\h�bMҾ�j�wS�!�;m맰����(�/��vz�|��S��^�%4Zq�{���=������3��T�3�>�N�hVMS��_*�WO9k�}�c���P���C�;@�N�l�|��L
���ӎ�(f۴A��:f"o�V�.JX����v�ކ�Q��pܩ��U �3R�yy�u�k�@���D��xw ��I�4�@%b�����WtdFCN��\�Nn2��[�R�������GA�Җ�F����M{�Njb�kbT���,_���7o:�UO��bZ�[�anԺ|�U�K���Ky���|��)�;j�jO��U!j��!���4?�Z�9��;�2<����{���O�����{G�����x�ǰ�17r��@C�%�0��׍#�Û�a�K�I�T\`��h'V �`����y<�|C�*��
e5��V���x�����Ev��R���p��g���PmJ�<�l�����V�x� z���f{<�@v*���N��b��>�dP��R�0K�{}����5RW�ի�0!I+�,u&=�K�}��3��w�-{,�q� �R�kYQ<&�� ���t&�޺G�H΃���MX�
$��\��F��ؠ
c�N`�;�V��m�vs�Ew��8�F�;����=ő����
�P0{�v�
�c#�{\�,W�xu��k�.؃�����g��Y7��2=~�ay�W��&@�Mؔ�%[kn��)է5�}��<�0�칣�L���>��u��
�	rZiN�]�-���Ƭ����tѬ�J�x�V�ނc��:�w/i�$���5��F��
��D��}��]���,���[fo-G��жIX�;��1��{zo�	=�{t��p�OiU�j�����8e((>G��TP��@8��f_U��/��\�(r"��}�#�ۆ�w; �լa8k��cYA*�;��F�8��wo�q�udt����୫���s,N��)������w)�7e��a��<�8�j~@�������	��cV-|K�M�A���h�ہ5��o��[��^|�7i7��.�v��hq|qK�y&ܢ�V �6+-]�5�=3��G��k��٢ӛ���)ů���ҝ�1�7���m�<Vsľn�|�q�f��y �G8�k�0��E׹2H=��Gri�|����t*q���b<?jՇ����ӣ�IS�ZB�,���^�4��&ij�g����e��Պ�
���3?��:�{$��-���|�5�L�y�廰�ֆB�r��4e�ev
�+uY;B�g��-��Ԭ����c-�]Ŭ��W�(5���Dtꭡ�L��R��u,��8�t8!����]R��r��,o��3���npM�����ॆ��uJ���P��eg"=M�����GS�o7t[]��D�U*�[(�yjs�Ѯ������.	z��B�d��|���1=�\ֽ�u�����Y�
K1�����N��8�:�˜��M�PN�I���V��cZ�;�o�'�A�,T�����rk7��]
(�.�;����V	-
������c�$}D?���f��Q�MI�]l�-U�6��ֳx�����Y��ƟU�I����QW��NQ6m�[�8�>�]�jx��.��w�P~��𛃂�O�Ar���	�W�|y�\s�ӑ�	���Z���+�^�c�a���(�ⵢ=�U��S6�ugwZӖ����?�.�	b"O�m�֥�u�}z���M�7RD]@��[�8��!��f��S��m����k�uv��:���Y��&Ax�
� �hTasr�����`��&�o����q|��[��ǝ�EIATQEm��***&��� ��b���
X��>�݊��*ӈ"#Z*�ҝvɬGv$�Y����!�DAMhuր��P�PE--%WGHq6ՠ�bb�i��&�F��M:�13�TUQT:ŻD�ACAӪ*������讒��N����N�)��v�Ei4%4���S�hh-��kIN�4Хt=)��t������z�:ZR�!T44��EuM4�����A��-!�E4�Al�ZZth6��vN��'������� 4�ݓ��
��z���1%&�CvSKE	��QbtP:����|4q+l�����W�
}p�����^ yX�1u��gs�$�b)��2ܾ�[W����SU�²�ew j�5�s����~�3+���.L���1oIėbF�zr:z��e�m�8l
�4;\�jf�8rޢ��fz���^�W ���fO�@f6�XlC�]G!�e\e�Jl���k34��ٚ��֔�r��Xt�[K\�c�:���/�
C=���{'�w������1���~�ꁵk�\�uߴ��^����k؈��wc'FF���A�`�����~~�����f���S�o�|����<���Y�nk���z�n�|E³טdb��G<��y��߿pw��y���ğ�:�h���F���8}�0QU�$���~�6�7�v�R��Y?M)qj߾��}�h�U)	��F�b�������6��
�l���~3���ΜF=��OZSBD��Jݣ�:���oD�,�/r�{a�^�>]i�������p�~���.#h'��*eʝ�yGM���;���`1fs�ԫ������ @�{ˤFy$��s���=�bl��/zn�<K�>�Kӯ���-�Ӯ��W��Ռ����Vx,����蜾3���J�"�a�wOg�PEZ����c�RXU�%�?y�7�h����s�'tY��=�0�:ڔg:0�Xq�S�����߸��?�JkR�j�
��o��̑pt�gFL�L�5�
f��<��}T��9�j����� ]����,�rI^8T�ӈ�X���NQ���3Umy�*..�����k�HW	��ȸ�`�L�أn��r�����M��I�~�W ݭ�W�wg2<��[o$�eq�v[���&�y�VD{v���$���6���ה#�!P��,�duuf���Dk��jF�Lh*}q�)h��=Ҹ���]��8����s]	��ѧ���`1�ǐ���\n�S�ļ���.�[����@�4�����#6��5��3[�#��3:���T;�[ky�Td�����x����#�I�ϻ�q��u�����>lm�.����M�^���Yl�U{u���;H'�R�|�3�Ɵ�w�Ìq���)���S�/�����Φz�AB�쓙V�G�Н������1��{���$�|�9to���B�i�E΍��f�S�=W�1���%$��YÕ�xr��ɝ\@l�;�\;�pI�k�3�y�c�4��4��9Rd�5�-�]��Ξ�+F�/�=��t+39+OMEQ�&g���ú�:��pC0n����`8�r�"Ex��ڸ8�H��"����.����[����q��-@��eP�Ci2�v�nE�z4M��6K�YS}�gY�g�r��ƌ�-��)����*�����M�9��T��q1��`5�{JDMu����<zp���O��;��FV=�ѐ�g(�����Xܔ�CZ��KY�����ZKfu������<ݦ�k,�6�8�yT��W�,w����U]~�a��@"a�6u�?e6��3���q���e��-qjR��|U�P����]>k�������}5���pUC�	�V%���O8���
Gd.��)�V�F�此蛝�{r*�*��]}z���Dپnrj�$e�"�c��G:���y�
^�6ᮍ���1�z�K����-?��4n�D�(�������c�W��S�On`�^%�-�/1#�9-R���T�a��@���]Ra=7���Vi1,5(i!�Kn�`�ݔFT`�}Y���xy8����l�%$5�/6�9��P�F�4�r�Z[�X���ҷ�I���k��<�H�n���E���r��z�����ƞ�O�ʅzh9�I�n�9G��k�3=���%Xu�+m�Gk0��za��-�d��;�$�ltU8SI�݇=Do�{�<�x�}�ue�cy��N���>�o4[��OI�L�b��ʊn}<\�ݘ���Ҿ�\�4D�n��x�>��Ww���{�k~����o_b#�w���1��s������59�d>̶mvBFL��-�m6��eՙ�l��_O����Y�/w�W+'�,��a��h�q��k�|��6u��������_K)9�;t�e���'�D�Q��~;��
ayb����q[2)�p�5.�,��޲�5U��Z���<�-�ji���[�~ePʿ]R���zf��8qɛ��Fۧ��eZ�8����j��Zۈ�SNd
���Lځ̄Фo�&ޗ�Y/1�|� ^�r�1۠sH�yض�!ӕ3��/Nܚ��Xʫ�xT����47C���9�*���r^�4�Ŷ�NE�&�ޅ��gL�	��b�o6Uʶ(�j�*sE=�d����rQI���=�K��t�d�E]�lX��Oq,�[܀�����%��k��5}���JT��\a��(w �R��I���3j��s�by�/<����H�-��۵��p)a���]Җ�R���͗�y�-����pt��$fD��ֈ�a��r[|,
�g].��<��j�8�MyW��=��o�y�{�9o�
����~
��,,q>�=x��aφ�OyI��ޑ}}��OW��b���%�Bs-����e��n(LAQRkm��SP�����e#��=z�\�2�T�O%�Dppۑ�Y���>.mU��J����j��;�q��v����3��4u�
�]�/Ε�5֦�����ƴE�g����؅�PEw��@�c��(����]�_9��
i&1>c&��Co#�+�w��d��gg>#�-��45"�f�V����W�z��U��?��9[��oY|�c�OmS���anǺc�a�vc׫H�V=S�L�1v�R��G�m���p"�_f&f�]Al`{�$�ț�歌��[%�s�L��
f�\olvP]���f��v�)\���ŭ����%�[�\�\}���Zr��h�Os�8�[Z��'7z�,��<�\�\��8�yz�ѷ��s]#�C���k���P�+��[s6`�3f���xn�ߨv29�4H� �R^�H�lR���(e��SZ�{�#����8�J=������M)`���S�~	�2�j��C��m�[�9�n�=����e���M���Z)�kx��P�b�]E�bg����nnmS��j�]�Kn�O��2���N��R�ĕ��U�[�.m��A�ن�����uKl�OF�ۓ}N��LzC]���Zސ:z�"Upy6,�0d���i�����a��J���X�V�A�4� AM�WCj�{��y��������.��y�#�G������� ;�!� )��.���JO�F�X��R}�m�Ǉ$���a,�+�+�֢{�2�f{3v/��]��8��;�Z_s'e���\Y����{��b�6��l���5��p�s2���K�߰����~��dH���T��|�9Ҽ0H��Ǹzah��=U��h*�kb٭nе^ꊓȪ�M���^� ���.�5���w9ݙ3��5�'WC]M��̻�+�
��s�)"���;�$@�ӍA|G�Gm�dM�TIj-1����~׶�H��wT�6�}h�_i1A��
J���Sϥ�p�k|�C��GKl��?|/�HC=bsf􈂍O>���Y(ִf�*��ˋ4էkk�mW�(����M��km��X�������F�JI��΋�˵���7#N��'U�ֹ�D)��O>��ky�����6��3B�J2w��ק�)��5�����r��-��1��Wv���v�OU�}��Ƌ�Q�� -�]c-�:�T��Z@&��q<���zά��OyW�s ٧�n�$���� ڑ|�=ݗ��H�)��X��,��s��Q[�9/�7ޅU�V�27 ���a�Y^�<��?4����$�&<�]�ʫ���tT��d��e1��#>��w_��&|#����($#r:�.�ۻ�o��D�R}����;�6ׄ�<"�\�u��o�ϓ��剏�"���;�U�Ǜm$|���u"���2�Rz܈�I;�A�J:_�h]����j������b�Gr���-[nm��ؓB_y��j�\��/��Z��Up�H��$����yX�Tn�n�.sm�q���&���2�&�T��~��WU��*�8�|/t��t��w���T�s�纪����:�ː���]�JU�pU�J��9J�tk>�p��øm�3�blr��$qآ��Hґ���g�l�DE�n�TkϢ�6�ڌ|��Sq���θ�z8.��򑆚;���(���!�_oo�<�����u�M����͹R���Ljޡ�b�4�L��R_]xQ|f���b��Y��ٽ�w-�G��*��n���p^?2����v��kj��yhۊnK�W���%b�s����F֦�3���k�u͢I�^w���g���xb0����C�bҋW
B`�����5��=8�"���M�W�d�ڮ�-t��H��f���;�=��{O5��x3�N室�3}<�$=bn�~���͙�o5�{ql�~����2�R��y�mGV�^l���.$�8���az�,���O'-�lˏ���k	��c������L��<W'��
=�{cz�;���j�����yp5d_Y��Ip��/��֓1ŋ�.���`^��mv�����]��K�O@��[�7�����-~���Xh��>�wS}{��P�c���!(o�!t<90�ba���<��m���,@�I�r�\����"R"l�L��$H��ވN�YX噉�I�Z�Cg܅B�v�.�ϓ�z����	&&\+w�2�=��c�B�_���Пy-�Qӆ��w�R�{�fΧ���n3j�4v�e��,z������=в�܂�)Aʂmm��T��TÎ��D������]WN���U^eW.�\��^{��`t%�
����^�<��5nA��ݛ�/x�ݪ�_ϒ/L�a�Z�9-��U˱���s�e��f�N��qݎ���D�S���z�{�r�] �3���_q��~�i\k߯�Y���.B�{;<�6�����K����ɘ�3y��a(�"�f�Т1�zrq��T:À7YTs	W��4����lH����
__R���t:;GJa��Y�/�'N7�>U�W�u��I���z���K*�/��1\�{�v����;�c����Ȥ�1= ZΗ����J�cxh�Qۗ)i�9S6C�k����͆N��Y�*NY
�v�v�q���>�8���g�����=�=ئ}��C�u%n��9p�����ѡ�8P̢�D�4�N&�->��3�W�vw��t$����WQ/���p%�;Y̶���>�kh�c�MCG3�����*8������n2k��})-CUݥ;�ڣ����1{�3�}�`���v�v�<�u�Y���5�ۯY|�oXn�i���E��[�;��� �;U��߹�d!����P'n�:�5��1#�U)�ԍ��!�9����⯰�Mt=�5���,�Ϣn���3%�n�d���ςV��:�4�5��KwU]���#���m
�ֶ]��_Map��(��
C%(��Fgww!��`mݦ��KU������쌵t�i�TLIe�F�8���eB�2/��4��=q�x�P�k�
mMwa�G��L�Qk{���=ޏW������}�>^7�x�|Ă"�.kSd�Nk���SQ_����T�+�ctꜸYMΩZ�!u����vb���C/-�ٲ������'�W��ks2���ڸ6��.HJ͟,H^���f�щ �rWDMuv1��a;N0���u�Z;q1�.7��Ld�0t�3�ev���r�W�����h��%�I����Y8��l��7����S32};�]H�æ��5��p/��P��5����t�����|�=��9�ˤ��!
5���Y��<]���:���,��yn����	��b� x���|X}�Xњ�Z_�g?������]S$k����\�� 3Yȸ��N%�ю��|��j�'.z5���X/i��
U���H�7��; ��v�X�X���A	�f�	~�B�7�@�q�#���\o�笐��̊!Ay��zZ��2��k�H[y���_<�u1�>�C)�����N=]�>It���/0�׻'e�[�\)�U�ݴk��t�)�T��Y���m|���y9�xy�b�0�.�w�`umY5����o���ﻱԳ�bz�yd'�R9]CY��l���s0�����nG����J��y�&��C&Yq>ޜ�bj7L�m�q�j�t���<��q.�f�]8U���a��<T���:;��ݾ/d؟�v�s�=�Y�y�f�@�q�"5�s�xoz�ls��!f����De�����d2�x���F�rYZ~ݷ�3��'̝Q���"6�����4#ґWG�Z>�����JxT�)���m�@�y3�兲�][��o^�e�]b�Xb�q����MK���8���d�!�PHz�w3�����r�s	�;::|s'S�s��+������ޥ�-��K��aO�;Ȳ|37�_P�n���ٳf��<��'-좻Hb7�b�z��''=������A��W�����&��9�gaP�wN�3�ŏV_}�(�Ui+���2RZhG��[�6Qo���+9��U*��^Q�@o�7���oN�����cQ=���3p�y�OלZ���<���ܗ��,,~�QT�xgc�zV�pV-ФM��9[��;���c����۾ϋ/��5
Yf���FS�mmJ�Ӝ/�;IuR�;7&C�-�ex�����*v'�ס܏�5����Ԓ����s�|{(�ym�$ўX`����K��r�#�`�L[�5y�s�:����vUa����|�(õ�gv�6���/7�1TA뇼}ۈ1;`x�/��"��0n�OK[��Ɇ�к;���H�f�3���v�?/��=�x�e�t�L��EYm=�7g3���\:ϓ�D�ZqK�/N�P�O'��k��q��9�VL����`bGs�>�;t��cHB
v���ef�����Ҝ�j�p2����)�nqˮR�J#XS���i��*�W]���8�Dؒ����KuV,���.��'%� ه|z�=[���}�C�4jm�IZ�A�:�X�5�A�����"x�*$J�WA�֪����i����wd�����S��Z
)
�����҅%t6�iAѶѤ�H�R�!��ִb"��:3kPS0�L��[d(*���� �CK�
+l�C��C�ch-��z�I�����6�!T�������UڃEU'F���
v0T@h)�zh맚������M3E]���V*��3-�6�-PbJ")
#a)h1+@�3qEE5�CHWn��t��W]JJJ

��IA�4D�g��t�&��Ј%��?���I���.�w����ŝ�Q��fhh�!��vz�ڱWc�/$�J��T��l��r��ӻ9�J�H�.�9�0�b�}��5�������q'hX�G��>��U�����n�f�n~q�A��1�s^�n�{']�<=x�}�L�0�,$���j�I�[ʞ�dkf;i4��E&k�lx헔o1��<���l��.��J�y[��D�����vă��jJ���Iǽ�9�T��C���S}M�9s�<��?n������il;�F�����Xk�6��y.��lX8tC�uƟtm�U|K���<&i�����a(�Zz��\ޅ�clɸ��J4��>�LAF�<�nf�Bޥ��͊1"wp��j��9�Gv�q���M�;���͡�b��QZ�`t����i�����A���9�WB�W�+�cS�3N�{�2��,уe��Σo��o6��!�>�Zuv��v�廰���%�9��
�;a��77)���v��cBE�z%@ޡH��1�l���y�t���C�צ�W�Ot�y3|l5��I�� �I3�';�u�w�/_a��h[. � ��h��.(v���;��Xi<�Fs���,x��a�RY��b34Sg�ț
�ޕ�8I#�v��[D .TS�/���+�k��ۜ&��}\j.�yq7��������뵧�B�17ʀ������<��u�Ɨs���	�`�{;/zȐ@͡�_�jmK��fʘ�븭����n��LF�My��y��\��#hr��V�U<e�[S�Rtۈ;b�<��D��n��Ц�z�bݶ��dj7F����;Ǻ[`5T7.�V`��-�5�
yƣ� ]�N��jIW�Jڳ`d�+��wm�d����6�2v�ի��F_�i��\바���}J�S�јjw�ືg��y�k��M{�+g��V�iؑ�tgܧ��ˇ�t\����$����f����8�W�����p�_�vLp]>{P(�e��TOw ڄ5�l�{2{b�qy;D�/u����G�d����;��V�9x{���׬�at1���cxr|7���\]wO��}�f�|q�m��ȝ{���>^r�78&d�p��,���R�D�g�o�B/�h��y{=���Z{5�m�ҷK�}�L���C�>��F��u�Xԅ��Si�l��1��x�
%����g�Y�^q>��³��q�߭)�����j┰�Q9����qV��q^��N	f��3������������l��~�yz})vq��$�B�s<wVXH�im"�_�hmFę����˨-G12m�1dD��^��(��!1�9;� �̷�3�B�˕��$t�z��ǌ��#S�vܘ����Շ���p��+���-��2��FYd>��ژmy���f@�����/�V���=yB�2�SPs��;�w)׻����]�ϋ����B�`��������ze�YО�,��d� ͤԷ��Y=߯j~!s�׬<@��R�3vr�!sdm��y�뎧�Õ��x�����Bmm;i�WOm{j�)���`�d
`�ֿH���个�̒�[ B�}Q]�D�	��ߟ�ߖ��%yG� `O���?�<��%� �i��4J�q���g-�).K�:�3>j��5��2Q콓َ�Cv<�PU�}Ms�R�!�8�t��=B�KO��\�|�.�0a�e{;�K�b������<΋:C������Ѹ�����8��&P�N�6w�򗚍g[�ގ��}����1sW�<�(��ǻ�Gfj#>А䲻%�Ux)�a4r=����p�z���<N)�r�D�6"k�B~��{����o��z��n�����`}�-T#����9=4���t+(�\����-���ޥ�C�}=7c2��ͩ�������[�vJs��M)�OWT�Uv]�w�7.4�{�.���s!��C=��L�즺���[dV���z�6����.|
�>O�W���o]��f��۸��l�yP�v=ހ_z�����0�LGoW�7mE���#��TWr��ړŶ��E^n�Ɋ���L�q���e�qwԳ�;���J���г�������E�ث	��t����l?`�j�~�P��: T�5�0L����\��\��9#���\�c�h��c�K����k��˒k���;����ڍ�sG�=.h���{��)�t`+ٶӀG]�;z���^��[��{��H�=���~�� i��3�~��^ʆ{��O��t�1;���h��Ң��RK6�b��J�f]��Y��&U�h�Q@CGR�v��^�y�Zۂ6�g{�6��?���L�=0m��r�ᗦѶe@���;�!x�N����X���:��hdz9/��o�"p�����=����Z\.F�AV����?�[VMA�� �Ђv�:2ߎ����CR���"&�л촧���$1-5���t������������׼BbrJ��a$���}5"7�w��ŬG^M��ʲ1�kZ�����r.++ma�"ջ��#-w�Ct4��}˃�jɜ�j��8mR/#��X^�'l��*s�ܯ� e�(�0�f��jj�����f��#j:4J��#	��C`�@1�v�M�u��T��+ȓ�O9�N�nz�:��%��d�\����!���K�.�NS�ݰ�D����-�!�p6�3�3��F��ݱ��4�o�H��h��#�Wb�<�T�"���_���EA0b�dW=��E�ɹnΑ�aq�.6�)��N\�$�Zw��6>z22�~�o��~QhSd�{]�6��Kqd�Op�A����J�L	$��;М�6��YI��~|�����;J��YgOg6���Y�#�{�|�s�+y�����.��hNr}�1��Jp�b�J̾Ϋ7&S�"�7hoP����{����ir�-�S���׹cGp�[+;V�R�Hi����u"����+�������.J۳�s(�{�[�e���G�VX��(Z��1��4� w�Ì�'-�U��S�lO\1��۰��M"g�t�&��t�ݧ(A�%�9�9QL(�Gb:z�K^A�����v^#�F��b	��LʢzkbFt�|�{5�]\e a�K뵗�
���������n���9o�M�z��y!z&�=���[�|��=�"&��h�p���s!��'���/�����={H�T�Ռ@�O�i���[+u�{~�^t�4�1O�m��m����xg �@�rI��Ê�b�x�m��\�(�mܡM9g4Y��6� ��G`-���gI��mzԥ@Z��Uܕ�����m�h�_4,ϝ�S�٭zZ�K$B4�2����M?A����)x�pye7`��<췯sz�����E:)��l�����X	�;�Uc��a���(.��rX��9K�j�s����HfR��Ic{RV��o*Ʈ����@�wZP^fq��g9;c� +�+�$XN�]�Qb�?þw�}��R���	]kP�.�[��D���*��*����
l�+f�q[�Z��c˅,��W��MR�VG\r>��ifz����w��Ỉ��C�G�r]bFE��g�L�-�*�f�S�v{�l�C��	�m����u:.��8�s��ս�๧ř�7rx[�\r���\i~��B��n�K����Ի��7<�ς-�Ӝ�M4VUI�9���t�}dJ�xM�)<*�3����F<���N3jݭ���5���{K>Mm�@ִ�6WLFl��R��u�8��湤&Nwk���h��zj��-���I��'}�+^�Xݴk�r�c�_(����N[Uj[�͡+|�^�G��7z�λ#����VdX��z���E����9�=����c���,�.�)Z��Y���!�x�ȋ*��ɺU�x(���u�P����ZB�O�FqC���N�a���Ժ�B�_H����'B��n*Ù*��=�au�όA�O!/S���t<^��Z��L�i���9�6�aN�4�N]�[ikĒ#h�����-^��b�Kt��J�_er�:(��`�$J�z��a���b�X���Ǿ#��ي�=����gYs�XT���V�N�H���5"(b�%�B�:�Q����=}�Ew]z����$f$��Cg����^�N�e�ٻ�-
�n���*o����`�i��%9�[��@�!9(�}o&��r�*T��!�{��˟d��{{�Eʹ��x`�u�����!�wX���98ߨ��Y�^�g�4n��w�(v�c�cy/�� $���}]�K�n�5�Y���IxN�>ᚎ�ǲ󣴁frA9��U{2oOy�����Q[|�̖��oE�O��3��1Ă��[�T{�"���;����H��3FJ"���pƲ���G��"(Th�w@��ǉDr����j�-�2J�u=�w�=��L�ޘ�8���e�Z7\�y��Ǥnr��	\�>i�|�*�s�-����3T���[�0�j�w������u�YP��n�d8��<*�W��?Mɉ}'7H�ic �Ο>�n�s�fgR�3�7��;��ۮe*��a�"I��sVM�)�]Ԅ���h5�~��1���߼�,b:oY�!O>�{�a�frU}g#�
���氭��k���<�Z�
9��-E:*��1n�+gQ��������b�}�W1�W���꾝�=��8+1�{oGm)l��v�&o�;R��~]��79��=T�����������ޟ8(ǳ�,;eR}��UUu�/w�r������c�]��Mc�gg�h9���pw>"���)(�,�_���<��Uf]�����c|�=r�}�!��y��\�J�ja�(^�ȹ���j�_wu`���Ӎ��rI"� U $�:�����������T{k�7�{�bo��\��@�/ n�$��!T)�N����v:������JUS,���U�DM�ԛ�J:kx���,�^f�j��k�d��������^�	���~��-zT鋉�j�*q�v�g\����"��UjV�y+��VL�����dd5�ʆ�i��Ӿ�n��cb60I�j~����ك9��e'l�� �ʢ��U��cS3��nd�A�U�i�o�ɬ�� ���Xӕؙ���M����ܳe{�="Aq��f��t|+�lre�=\a�����3p�M���zVC��)���Jm9�ԛ[4��2������mv�R�IK����5�8M4�α�}`�͏xTJ��5P�xA�'T�fXA9�>eT�N���$��Fr���x���3���C���Yu檺W�x��䑲�wm,v�*�eLgL��vڵx�YQ+���!��F��El��gb�j��[���ʜ~�E���ô=/,Z�����W�7)��k�>����jU#j�S��jm8w���X����ɫ�9:g����Ц��f�a�[���g���߱�]�rb���߄]���U{Lq[��D�˯i�:�۝��<�3��K�l���7qS�Oe��*��\��Z���(\�0gx��{���9ZV�n���*c�CY���B�#G�����(�޽�є��ۘ��ܖj۠]EX��týXg"����Q��	U
�hϻ��W��g˵wlP��%�2����j�\w;il���؉�TqweϽ�n�n�󍦝��cu3�e����#���`z�i����5�3���������?��d�~ ( ������������U]������>�oaDp0�2�2���� C 
�Hʳ*� L�0��*Ⱦ��AL2 2�2�0�0�0�>��>��� ���>�p� �T ì �{� 0� v�@;  a�=�� e `@d@d`@e@d@e d}2���@!�@!� !� !�@!� !�@!� !�@!� aedDa`ee c�Up� � 2 2�2��� ʪ�( C C
0�0, C� ��ʰ�0���0ʰ2,2�2�2�0,0,0��� �2�0� C*�
�*�(������{ߏ� �P&QU�?��o�~_o��� �����S�_���������`����_G����}O������߷��@_���O���EE��@X��7��� �~���}��C�� ���p~��_\�����>�?�?�O�@o�����o�� ����4 R�  � L�� � B ( I
� �J���ʪ�  C
���$�.%U`� !�U� �� %I@D�U�! UXHPB �UV%Pqߨb��/�����*�- )@Ѕ�x������(>���@����}� ����������;�O�������ov?�����D U���O�ǿ$��@_�D U��?�x�+���ǽ�U }��������_0�7����=���p��� *�z���Q �J���������_�~��������������� ���������_��1�`�O߃��������$��=�@_d��3?���?g���?d��~�QW�L>���(�+����~��g��P�~i���
�2��$hKX��������>�����~���JTE!%R��(���RU*���T�@��TER*�*��U*"D��E%)!QR�B�Q$*R�Z���( R�@*)%*_CU�4�H�D��$D��"�RE*H�*(B	P������IJ��R���j�lJ��(AE T
�YU�P���(������T�T$ �R�E	*)* �UR�U@�����AR��R� ���ش�m�aDR��mcj�5�J��0m�hkj�Tց[m��I�fm���[RKfff�ښ3[�
*�AR�тJ�h�U�  D:    ��� 
(P�Ba�� �
(;�à�]�Ym[j�ZiM5��m�ZL�ԩ�6���3J��V�mJS4f��f[5�AQ
QH��K`�.   #p�����Қ��Z�i�Y��m�P ،SR�
�[#L�m6٣ hV��6���U�Em4ڥU��-��Z)A%P �j����  � 1Lj��j�cͩY*�bYD*�h2�U[lU�EaR��#V��+mj�R�Q��T%�2p   ��d��UhZeaJ�Q"�J@f��(X�f�Vڢh�	UU��$�Z�0
F���U	DT*)HU8   �*��d�Ѷd٭P`�*���ՔU�R��+a��4JmX�a��U�k-�VUR�(�R$*(��K�  � P�`i
SV����I��
�ҫf�URk	A
R�  �� �  UIB�(D�R*�  G  	�m 4 Z� ��`  X�� 6� cK  �` 1�P -�  U@@ (�I�)P*�  G@ 6٦ �1�  SeX  �H � P
c  S  �` �*�� �U ���E�*I� g  �0 ̬  R�� Z+ A�X  ���  � $ ئ  �@ � 
   "��JT�  FL�0  E=�	)I*4��@ �D���"2O)��146MO5!�JU%       �~M)��4�@  @  �I�R�Fjd`�	�4h� 	��D���bZdhqA��@b�F���Nww����N[��d��!	:����=B�4P��@ȍPUD�Ah�̀P����������?Z�!��T �Q8 E���DHF� U!�+�".=�:Z�X�9q�ۿ@z��쿑������_��w��Q���u���?�O袵R����HP�w�K2�T�-��L�Ͳ�%F�n�T�cY):�^�R�1cϳ-��qe���dZǊ�T&,cH�ɦ^����l:9����ĪR5n*f���SERj�d��V�-Z9F�LD
�en0�J�e�غl��Ц��*��u�PL���;�Pse��IT��e�H�]$NޙD�Z�k%DR#l�BW%��n���ʳU�Y�*P��۽E�Gq�L�r�p�d��!��c�`�1��/)�tj$�,�]���Pf-˧Q�V��)��A���d�W�sL9����H`C`�W��8� �Q 6R�D�/H:�#hIR���<&u�st�-�k0�r�T�[6f�Kc��i�����,��k�HK�����&%1u{.�֕�QX�#� ���s(qa��J�7M��é��u�AHɷ�b��`y4n�ۺ�mi�雖n2wuw(�{n��b�,�N�
���Z���b*tOh�ںZ��v���eչ��٧Ak��5/Z��U*4Ј�X��ڼ�C��h#YV���#��F��,Ӂ)y�l�L�
-�Gr�6n�%����A��j
��D�!.&�f3���d�[Jd�PF�n����:�D%6m� 6��Qk]hŴ�)��`^���W)�rnFӣ(a�w�l�YZ����(i�`Fn��vH[-j�R�A��zeL8Q�cs)���j�;�6�q�u�p�T�*��'x��&���!V2�]�A��Ip�������f�T0���a�� �Jt��[��3j������l&`Ac1���_���&Z؋wO��e,{nk�2��:A��-�����Yy$���*fb�ʊ�I[tB��ZKv����V��S26�@EMc;T�Y�ƫPn��1��-Ye=�,u��*���CT �w��6�Q�K,�'�
�!����j���.�4���L�d:�i]M�ǉ���� �B��n�V)AF��[�i�&[�qd����0�+\�6�1,��z�����Ԡ\�6���62ʶCGB̻:o��70KQ�i!Y Ǆ�Z�� ��NS��;2hM�hd�{`�y�m�̨�h0��L�X�s�ē�+�d�9�S��8-'�W�YI�Yd�x¹�Fu7h��8���K�Ӗ@wX���� �ͺ�wIݠ�,��ne���N�d��-Q��F��ɣf�`f�+F�����hc �i�����^U�b�<[�5�N��!L�FE����h�aSF���>ɒއ�9�0i���e�uv�bU'µQe*�74�mbwy�b�+8��m��9��1�;WiӰ�Л�/��QD�6R�Նf�pkЪ��SJ4��u�t���3U=���u���e�qc����G�%�e��b�:l���Б��jRɖ�¥[���H��Y�Fm9HR�]Ƕ(�jn�eb7�������b��"��4��ж����
�Y�6��e��`��q-Vs*<�˨l܉h��ܻ֙Cn��6�Jf���v!�OR� ��%'N����=�qހ�C17����e��-f֭� ����N���яT�@��Z�L�;@T�V~��,��	,���u�0�ƫf^#H"���BnŅ��x"v�!�B�
�:�Ô�����j�n��n)�[șn��<�nB��C
��Qu��E{V�4�wt"��q�Л!y	�s��	�+�f� +jƘ�H�A�z�Hq|�ͼ�Zn�1n�ob���5���`�F�r���|��^��Z7j�eL����he%dP��f�iV*��N�N[oQ�m��b�1Cs�M�OK�[{�;5�XͳYLGK(���yf�n�2�5�#A�c�V�ڻ�h���[P�!�6e�*᠙m�e��%%�	�%gZ����ECY���1cz_�/mk�A�.Y`h��r䲱�-*i�1^���א��w�Am�v��P{r[ҩ�X��6��I[�0Mh�	�\��9`i�Ә��zF�B�Vq��Ƕ�b��P���"ڏ7E�t(YT�Cub�O6;.���Z QVûR���\(��rAS%���xt8 5��l�xʢ�,`V'�K�L���<�U%�vQ��՟]3�M�1Q����j{���r�2�l�E�A$��J�CL
 \d���(3)fa�jȫ	MȲS�ne�Tj�9n�FP��ƴ,b�efE��⺲�e�~Ϣ�3r�]`�ݜ5����De��ɩyT`���;�8D�rnPt�ٹnPS���|�P9KEG�0�k5�6�m`/I���P��k&dfn�j"c�O镉�f}d=�n�rP� �)Gy,|m�X�3h2Av#�����拠�Z�8b�W�����j���zY"XY������W5����i��.D�Iݗ�bh�z�)b�@~�:40۹kcw�J�ubD�n�F�i�4?�ןX�L[B����Kpy����_
6�+akm�yg&�f`8&K�McCl�d�d��t��f�e4�^��ej�u!�{�*��Si��o�6�De��R�)[3t=�cYV,F`Ƥ8 &j�6�Y�����Qh���njv�r���n�m:r�GkpY3eM/1)si��ܑ�B���wXԌ��f$��Z1bK.�1M�KjV^؆!+"%�5��v�0�Sy���<�ѭa�t����f엲�L���w��ki����bb�؋uxZ�)�]���+ z��7"sb����PncN�1����i[��YhJ�����b����
�w�R���`�h`��A#��e�u�oQ��v����R�Z��v���m�W�+\`�4�-"ƝgnD�9x0#rB�����n��1f��mIt>X���IN�!�Z
R�m�nѴ6��E�[A]�Р��*#u%��ӣWt�W�x	�G);�z:�ۥ�]_]���9>�0�b�u"̽a��ה7n�7n�*fmH��n��tqef�/Z�so	�)�Dmc�n�Ļ��`�[�KՉO��&c˳��V%��m�w� ������5TC33]at��y�K��Yk#7���mjxk�ce�#W/l�XړkN"5�9O3&
�����SԔ��]�(]�&��ءn�%,5�(vX�)PL��wT[�
�0(,�����sQ�2h;��޴6��t�7yzb5��	M`�bNa��P^,��
�h����.�x���T"�{Wy�ķh�I�����v3��c���)4�%Q2=�,���P�M9u�����K�BlJ��f:L�i�N��ٌ��_K*�G�H#ջE�љn���K*%-D��
P����,k��f�R��Yܓ����8�[B�T�oN^I��į	^۬ z���C��u 7)�YX�����ƙ+,�WO���fL:"@|��h�W��CM�n���I��H�-Z	�1+��S�S
���еv���!ʓiKFI*`6.��7bf��%��u�x�8����o(�ʸ�{�	R'�}sm��K"�i �R��X�䰰����z�ç%7x����Zf,�0jm��7Sqj��	�t%f9����Eu��@�ni�p��-Wu�su�
L�!��>�c�E�fS3�,�Y+md�bГ��Pv+u	C@�t��Z��%�-���ݨ�Qim��نܬ��G]��-��e�c	3,�I^1E�ŕ&��:���E�RL7�Hn�anX�Nl���ؖ��H�*C��MkX�[c&nů.��o$J�<�F���-R��t�2���&�T�j�/l=��dF��P�t�2��a�����iJ,Z2���c�U��&c'?m\";��bKU���<�46�T�(-
�(r`�F۱���R�nQ�6X�X�,�y��M�9�b͠��{�2�S��㤷\p�v�*���	��;t�FL���� �b��[�H�34թ&ɡ�<ߖ	RQ��8R��Ke��Gt�me�҈��pv��^H���41S%�&�.�iʘ5�	$k���XP��% ��:�+�n8�zr�lVU�)�2(�W�߶�S�kT2jlP��,,�X�uus2�e)J=����PaF�uF��鋫(��+i
��`�(��P[vO$ځmԭ,��/j���k��i"���mG�5śꗗ�ˏc�i��E���P{m�9���'��,�d<��1�p6۠�{��ohLE;o,8aE��ۊ�Ħ)4Ӭg�ŵe�J�H��T6��{m �Q8Jx�k�atjD)5���-Ra�鰈��� �R�}����Mb�YnmV�l���и.ؔ�	v6[��M��m-u�LN�V��e�z@�"�;,O+�B�dv�;[B��%��E�E�XN�u��������CojޛSN�;(Ja�{��+�f�˫Tq4Z��E��l�p3N��V��R���fn�T����V���^Z���H7Sa)�VA�#�q�ΰX���S[��a8���Z,��-lVCM�$V��̦�H�6� 1Qz�����C	���.�^'��y�{.F�;rk�n��^�X����𐙤%�8�U��t�C��H0R�VUc���u�e;ͨR�p9��L�Yk�}t��Nh�l"�-�*�xcIIF�R�iȶTV����4mmp��];g�ԯ>M�l*ʺ	1Ee����ZRV�a�>��/I����fU�W#Z��>�a%�� �÷`n�U�ؕ�*՜u���
hkZVe�t v�&X���-_&�ktZ�Em[Ucd�m�+���;�xt-2�8��"�6Ukh^]�$襹�%��,�bO?�fø��=��T��nT��,G"�N��]�ǁD�"ұu6��Z�m�V�a+G�O
��ǲ�^Bn*ִ
x�(�i��KVJ�y��cF�wh+	fjem�_l�j5���je��mmJUp�7Z���QP�k4dv$����F�eѱR��˩-�U����o sn�[E^���t��B�X�Ow2���(��g9��e�Cn��6-")�Bڎ�ɺ��ѷ�i8v�bƎ�2��p1�а�Uު�v�m���"d�ݻ��9��6�"J��I\36;2��̭���k)<fFE�ui�4a�]n֢���Y&��-�r�R�gBI��p�õ�*k���� ��I�a'M&�9(�e��B������A�/.��M*@0a�&Th�#t�һqt��̛z���$9R�Ŭ'McZ�n�znJ+��Y6E���6iSZ��E��7j�C�[J%�ah��r�z�[d� �j�f��3Yz����i7X	!�\�c1�$ɥ�G�-�Vd*S�j��]iխU�HbaX�e[�)$M�z3BR�2�M��衵m��)V<t��0Ҋ�n|�&�ab���Y7�k*@C���0�?ekP�䡯.��\T˃&B�+�Kf��w��݂Ź�㉜݇C����]D�Z;#�Kj��@нQ�A��l^�0���HG&1bV��A��F��z�<cm�["���n&t]iY�J�4*`Z�{��E+2�
IH�m�;�؎���j��U�W�e��շvˣ�eAr��u{�N&�n���[Nkn�ܡ����:�Ԍ��8������H�*8�ǳM�MD�kk`	,�,^�B�ѫv)��:h�����`8Ў���2ı��MZ�5�� ���R�P˦�{]�╵�!����l�E�r�ke���T˕y�,�/+I+K6 ���L�-7��3�@2�����II�ӧp�k��"��i�;1ee
՘ފWX7�y%d�j
��&\����Z��j'��i[v�
":�����F��ę�]c)25PSH(bY�,��U/s[[gV]i���Y���3E�tF"�Y��BA���n:��4"�5�òҫl�"���6���*�D�#���X)��E��M5X�L�B����fP���mƬ�-�#�,h�����&RH�wm+�E  M���
4�L_Ite��q'��p��j�;
�ZTo.T3	!^��+QI���9I�V !�ܼ+쨾�2`��vJb��5x��~&�h��pa3�C�RXN�)���"���V��-���)0�Y�4oj=7N*�A6�<ݫ/��*��c�t4벲�nmF\MӸ�껋t9"yrĤ#q��Ň2�n�6 �G]5H�a#��&�ܺEk)�t�S.�t'1T���y�M����t��rf^ 1f�,
-CR�ͤq`�h�`�#)���n%��[W�̼Ȧ���be�9j�YV�
���t�9a��ӢQ�U�c�6�˥��	ñՍ�yf4��]���j�����EQ�YZb�u�j��z�V٨�!��]�xҳVMhZp�j�U^��F�7y4�Fj۷n��n�j�U!z�"(+݃�XUk��X5�����l���ϋ����L��Z,��x�n4��Úv���u�&
)���+pmmD�2���n;�5%�(o���q�S-Y��Z������߇�:<N��O���GV��(]m
�^~���i?�|Ak2�f�i �	��%�U
�T-]p���|��Vk�|�8��P��wMt�
�զ���ݖ3�S�v���G	B�2O)�)J�0֋Y/]gv�05����Z(��šZk��^��� 5�U)��W�.s�坓y�Wz��m�:����fZ�L��g��tH�l�D��wSn�iG�04F������B'ت�����&:�#��`�s}�3D�Fen�惀�M�Lv��V-5�u��$�g&n��A\�\w:��gL�2���ԁՐu�'!?;�oz�F���#	n�FT1>�3��_ܝ�v���4��9����44ha��u�U�u�Lf��~�7�\d��F�+�kɲkj��f�2i�v��v�M��[C��]mnʺ�ü-�n��q5{i��}��V�U����e��֭ ��F�b*��.ݺۺC[a_)����Ҭ7��z��u�S,�\�GH�����-k�i:4�SOc ˴�Z1:?�Y�Z`�T/r��̚x�+I�zd60���i�Y�JYt��T��o��.�vq�a��b����gtޮ΋����e��,��G5��:��[켴�\��I�Ǆv!��1���z*�*��/qoE�^�ˇ���
i��ޫ(�L,Z�}CE��٬;��[|�8t�%�8s4���ub�*b��*��C�&v=�G:���x�d\J���P�d7��4���ӱ ��J���I�n�T���q]&`jf㷁�y��#�=�l�
F�Z�^<�A��0���Vj	R��*����ð)�r v�.7����%no"�S�u�f�m�+���x˧�u���Zͣd_L�^�&�L����2���ʞ��ԏ�l��D�s�k/��O\�*��u d��B{:W`}�gM�]'�3
�qG	��I����S�v��﨓#*��#!�n��ƻ`�b`��t�;G�:j�ي�
r�/�Q����3���P�ze�Uv*"��TцM{������0Äs���C-��X �ҷ���d�mvM��|�r娋Ky�\fؿ���Tx�wh:ۤ��&ȉQe�V-��ᜭLY)aӬ���+) �3靁^��X�M,z$؏wb}�a�`n&����Ķ2[*�c wJo�+�of�%����n.9}�n���9����th=܊*{��U�e��+R*eϯ`ա��HK��΄�qu���:�̐E֨TZ0��}��5�����V�ۥu�mj�V�s�X�Jun���7��;p:��'a�%KxZH�I���&�t���S�+Yζuuy/] �fd�'R[�s�
��S"of���KD�}*
K)i�9���s;yȴ0�,P
<'+����t��}����7�|��M�Dv�zW(��H��5�fv�=].�Q�{�*[���Wg{:Sw��*]ө<�
:�X��c�K4+����-�)	�.�|��u˙�G�X��ئ�%[������ls
ő���n��k��t��K-t�7*��ơQ��+-�f���b��Au�IX����WX57�	+�T�~������]���)��.��1Π�o1�Qm��JnE��mi�2�v�� �ԍ��:�ͼ�8E�,��'v+�`9x��B:����D:9����x��[�hu	`�P�@h�/��l`�WX�onJ';�_1ڲvؐ	�-�m۩+�T�v�3�U�u���HZ��0E������/d��s����-Q(5KWL����һ'%H1[���p��D
�G�����Le8/��83X"Q5�p-Oa����,MDuǙy��Wx��6�fc���w>'�H���2#q�Wn���l��Qꗳ�K|�qW �c*h*��/Mk+��f�[P��r
��ol`*j��[���D�tN�m%����b��D��*�ޙ��GhX]n�(js5���6����(6��p/�8�[���"��q�E�K$o׹�(�d����//���D����T�V�]YO2��.�eo9[���Ol*�
C�_`�ES��Z���Tن�3]ZM�o��j��P��'��n��:���R90�������כ*����M�[���y�`A��r��(����(�.���t�W[+��fé����k{���ba�ƺw�HP�>w"�{�'Yu�(8X�-K'���Ѿ�6�:ژn^
��kR���v*}/)2�G1J*u�������u|�Obw��<�'F��3_��[�v��v��Io��`�;��>���{�ԡ�j���0͠��9�E�v�ӈ�z�,C��\^��ep�E�J'S�hϧivpw��=��y��շ�n:�����8Q�������V�[΂��l>W�9���h��VJ3�jS��n�������%���h�jΩ*��,�e�vշ-4��r����ܰt@�R����nD �r�˧Z_Ru&)�
��0�W���`O�TP�W�l���0���9�ш�5���0#wK �`�ԖLHU�eH���];�[�N�r���/���	�Mc#F��7o�=^s�;�f�[�݇���g!����J�y����8��L0����s���y[N��4��XźM��p� f���.-����zpb�V�:Z�����M���
꾢�����w�i����a5"�/\Kոb�t�:��e�j��j��i[��U��1uޝCa}�<��8��(�s�B�촲�P�bٖ�b�0�6�r�����˓)�S�x[m��w�"8tږ�odc��լ��,��6�`��C\�U�ڶ�7ׁ'��Ҧd�����b�=ˁڱ��|�%��=���$�gL�)-�+g�q�۴Ei�C��x$�ۥ�����=Cl�sNo�PZiO,�,��j��^^�V¸<���L�
���Cf�Y�zL,Q49U��׶�7����ó3z���Om��s&y(��c�K՞jLg(�(z4`�,�D.�w��RjڣĬѳE_fo7HѢ�ͻO�7u.FX�#�j&:��W�ܹ�J�kb8>)Ii'K���Q���z�T���z��q��w5k��n:�}[j�`��WQi�]�:>�le��h�5���!���4�A]�����]h1�p�M�g�~Ӧ�����ݧ�S���J��<��(��wC�C�\+���P��H�Ǜ�pf>���f�$Y�HxʣV`2�]Zw��E<��]9���j��s��M�◗.G���|.�B�7CM]����|�:)YO�7>��������bzjEe�n�7�s�(]���u��׸�t�1ۃ챶��3	�}�~y��u���������<�j�u����G�l[b�(��wj�,�Տt�]��>�����R�p�H2r�>%*�O<�8��oc�8N4�D�Ac��ͳ7-�}.���+��h�^�<�	��vI8�@�]���E@�+Z��vA�����](���z��v:O7�{ե]��1�Ov���wAS�w�ǜ��-�*�H��v����JĬǴn�v�Ǘ�k`�-��G�Tڽ�>��4a��J�1MM����\�ջ�,�.��bkP�u��/h1ݵ�VΩ��u�W@ؤ8��`�a�9��V��&�5E����m=i�Z8��Lft{�:��v���dU,J�*�]l�Z��5��	�G[4���/Ǒ=<�ψ�u�_I|���]����m��K��^!�e}�K���i��\������z��Σ8���4�(6D�l���NR<M���:�u�-
y���sw���$�o+�A��ŉ}���Jy����i�JZ]v}�d� y��B�];4d�()���)�dT}A�Hѥ:��ЦC�}FMj}�v gn@�#�Q����駖��#�0�ǎj�9}-��9y�f�l�[�9��C�u8�wEw<�R�Gp=��E��8_8�h:Y�����-�����XxR+�C�G/F��(�{��+dۤ���
��v-�/�e���
�,�cq�v�OX���fb��7*��(e��Ԣ@�D���vi䶷+	�+$��4��b�S[ʲn������TUgl�]Y�(c�T�l\-/r�3�z�o WwԒ�16J��5��ݣ�ַ� ��UK1p�L����7��mH�fQ�c���s�Tp+����a��^��G��ǹv3����
:_�Yw���o:q=vI�g��0�Z4k�̛j&�oK;WS�յ��:�u]��/�OO{ �ȇYY��'��)�
7{��6F��_��fa��4�[��� ����4�CS*��b�ky���P���⺺�`-��b�Ɖ =R�I�������s'M�}���^5�����CV�p����L�y�X03͛����:�ĳ��D�$ޭ���<v)�;`2���z�ju���q̮� ���l��W�ë���#_�-e�W��$�K1�W�չ��J���6&^���W��`vm�2Zj��cbU�g_\��>�!01>���5^κ�iP&����E�V�В�8����GS���Ӕ�^��3̚�q�Ǉ	�4NԽr��7]�)�ܹ��o��u9�]�5\�v�_#A܈��Z6/_��ܻ.�&��ۉ�B�,�CCu�LL�+r��_F�y��y���]e��o �&v��cF�ƪ��|4�휹Mj�k��f�֤e<�iu{v��5�Mf�I\���|������N��0m
����HDk��f�V��]��g;ZN��:����6멅Z�.�gqO��t��{��*!�mV1�������V�竴ô+1�:��w���촆�y��ܝ�$aQW]�lچ3^�O��J��V�����ͭ�cjW+r�ܴ[J�+�0Y�Q�0jfb%���*����ږ�"R�	<Xfi���l��wG��Ҭ ��o.^܏����x�a6�;�qR�9�h��)K[�kR}zM�j� c�)���Q�n��Q� IJ@�pn�e���w]�p<�zx�l�rܶ4YR9�-P���
�Q	���*��ݥ��m\al(�he��w/5`��̈�B#������-7�m�K��d������m�#��+T���Ĉw	W�N3�gC�N�^�5m���JÕ}�E�2'`;t����L��k�vm1�Xt��C����*C�-��O�����]���=���"�,BNو��xR�y0�%1Ỵ��UK��q�9�l�ʊ�� r�o���ܾz�N�������-ZY��c� J�����YQ�=�,peo	V�k5�N�j;[#k�Xz��z H�m]h1�GQ�-jʶ�|w��Lp�,k�wte@$�5:7�R0�'��l[�Y7�23bP*5QY�G���S��V!��.�Μ4
|8�M������K�U�ov�	��5� �[T�|9�hK�����.5����:���v�]ȯ����qfb���I�����P���3D��
�O��Jq���z�.�s�st�xFc�������̏F��*������݆͸�gZ׳��Of7{���� 4ɣ6iC��.m�6u�����Ƕ��{�M˘���j=��sE-B�oi�*&�V�Y�����i�f���Wg9�M����A�y���FrD^}۶��ln|�f[ᗹ��A�Sv>K��ԍ������T��bmk۹�IB©�5:���%�>�t�!u3���yj�q�b�/9�*1�bk*�*0�s�s:�%X%<Z����x�기o^�:�H3R���\��z)�r	iG����uɍ�f�5�
�����}1�nѓ�{n�ɱ5�\�A)y#|�ҷh
���7�=���P��"�{*K/�oF�ei�ULu(�w�a���ي��<�m-3o$�um��B��pV�t����;L�C.�$���I�vu`���v��BQ9�� ������TL�<���ydN�ju��7+Gm�n��h�YR�5����|����j��苸�+��ie�`䡮��R���͓imK�+-��o.�C�.��J���.��{���L��I}j�d�����VM�P�m�}�CH'��\�j���\���zg��U�e��\En�;�M��w��N!D�M���a;E=�����r�������C���O{yU�[�kv��`p�d����ϡR6�wJ��ag���os��g(.�w�r����J��GU�Υ��#mb:1q�]/L蓣ٳs�é�H�aW*GWw,�.���q�4�i:�5�E�Vw<T�"�l66���{�uH�M������J���)sZ�N})����O�i6GP�"<v�d����h��^\G�ٮwZU�m.ru�PoTtRk�Eux����/Ewc���n���s#�֫�M�j�-Ҍv}�xE���LjN�B<��(Jnܸդ�2�v��AQt�H��n�!w�'v��)�ja{X��Zpc���-��X�鄍ۇ&˙ԫQ�n��;��^@K����p����g���b����[�z��m�c�`�:�Uw#|�]��SE;Vqn�lò�<��9�Ve�=叄~>��Ư�fIؕ��vܝ9���d�m��s�{���]iL��YW(�ʅ�~����z6�y챧����� ʴ�Ȃ�.�ƈ�Ҙ�� ���'��^[#J�
l���mzFE):���C��s�v�6�,I�4�m�_$�hw��������3�}R��݌�\��yM-�hwM7xd�x*�MTo@��c��\�8��.�����il����i��v�v��
JH
[����9�@*ܘ�c����1�����`�y��K�W��c�,��67��U��ӍE7��tˏwdu����~�%P�Zy�9�n$���n�e�$/Ws�1�\��;��f�����db1I�F����A�R+�&h��P�6U���y�}. �S�����B4�h�����AE���X�QC$���E^}�͏^j���X��Gl�j߅�^�W�)�z�(������X[ �����v�q+�ţ\w�u�ܬ�1+�k!;��gj�����h.������r*6�G�f���7@D �1�\T]�:m�YQ6���fQ�x�7{�:���_fO���J��L!Ie������4&S����}��1|���R�V��F/���Z���\�}�ؕΡ#���+t���p3�p �*��M[h*Ǯ��)أ��p���*���79�����-B��������[H�s!r��dдN��]���+�G`o#����h镒v����2Đ�w������!v�t��č��*���YLγ�rQ���V�|���̝Vj6p����p�W7`�^٣�:�EӨ,�n�Gxgnҕ�!Ā{�։��s�/���[mZ�XcN�k�7�=���6�,�w�'9d�=]��SF.�h��9M���H�n�Xȷ�W"�w%��R̽znT:��ր�V���� ��%p}�5J}6�#]�ܺ��|~E��׍5���}�K�@�{�����h"�������e�߯�s�u}˂e���+�����i��`�&�]��VgZ��.�[�˝��Yݫ9�x�~S�j�k����+�W3:�E�oh���d��:�FI�6�[��oS�Ts���Als�*>��az)�d�� �JWyV��7�OJk{l���� Yˠ�SrCaX�[-̂�Y��6���P��P=T�oDT@��:�����_@$J�:Vl�����K���w�z�+���h]�wb���p�Ļ���0kb��[;�t
�n�h��u���d�T��4��/^�R�^ثZ4�*3C�=�T��#��dL�rÎ�bbz��gm]�:�#�n���˼���!oR�]�Ӂ�ɦ[|�˞,�␺��t� 2�rgq���z�d���P;�)w4�\!���w׽���ˋx��Y2�\Bw6�{p1KŻ���e̌l��;E/�����	2���.��r%�r��Nw[U��.j��>5hV�*2����C�8*hb�Sa�`��+�t'��i���5�uu��cO{����׈�T_u�Q�$�W��[�v`O:c�~�ГV4u�)��Z#�0�e�Y���q�M*,o�KoL��U�3��qZ�nS�iS��ҙ:��c���3���[g�a�]�q�P_;��[�o�Z/p�#�z	8����g���;9��K�ۼkD̢/9�2+@���±IjK�3�X�ˍ��Ӗ�����3�.�7�:�/X�U�wJ�jT��{�l)���ވ����Aĕ�@r]�̗�ſ]Ҭv��\�u	�I���
�� =n7�p�sH��̧�5�.��/v�I�aV��b��tզI��d|kv��\;�*��;"	DeN�:�Oa�(��¾Q�-0�{�G=�Wy�*��vԕ���e�j��ڴ_Nn�̌[��Mw��F�6���Q��WB�H�,)J�R*ʂv�. �ge&\]���5�8��fY��غ��9+߆T�6��r�ul�؞^�4{�zo+j�9���lHc�q��7�%F<+t�i_e�V��4V�nƭ��"eѦ�V4�EZ<H�A�JX�f��ɳ|�9t;N��4��i|ջ��D���Yk@�BY��gV�K�׎��D=���h��|#k��9��m�&������7��2��])�� ��]�<��ٕ�]�s]�)񥗉�ܕ�^R9�n�t����962��c�Ô�oC��1��m��IoeM�ԩ�Ud}c.MwO����\p@+q&�umV`���[�O�z�"h�]���60A2�{]�@v�����^�*B&ֆV���V[�m,�T�27�r�c���ä7/��&%�r!pz���r�PR�\��{Ñ�v+��YG�p�a�*�7����Ӧ7X��n#��i��Z�PW�\�z��\n 6�w%o�~YWKwq��Vѱ���E]e;C!�vIL�P�"oz�Z��+�;3�#s��w���������T��I�����Blݖ�������A�w��aW$������ljU�tS����!r��<E*�j4���^����ݭ�Gk9���7ٛkڽ�w�+z�ԛ�s�/6��	:�us{��F]�����pN����%��WՓZ�f��[���F�rw)�Hf�((��mWfkf�O" �ee�j%���.�����V5��|�6[��BP!�KVV=����[�G%����]��RCv��Ù�	t�d�
�.�n((�E]�ʔ����Ϋ�X�`�]�Ȕsi M��eY[Ǳ�	T2�.`����L��R����=x=g�a��W��B�b�U�q$Y�ʴq�ë�smM�&���O�K����Ҋ�	�^��ݏU�:(-�n4����o7o��,�5����-��0�Tu:�}4�@�u� ��+\]��������auδ�Ef��¸�Õ�H>�E+�8B�&�8^
jv���{�DƵ����`���ڑ�g^͖�<���]ٲp+��+$@;�#��:+5۴�#��|�m�5|��NS:�p����.n�%s�,!��u^�ڀ�S��_\sh��i�(�B�H�(nŪ\Xvt=89���O���;����5�N �Xc��޶CZ�`Z����s
v���x�@h6��{�F˹�:��E�[@uv��B]v�imt9��3�:���h0�C@Vv}��|��w&�ݡ7� m_t衑,c�n�����ufjv�v,�W����Q[p.�`�MmQ�b�����GXf5b���ׄn.��n�9}�4i�[�]�����L�W@�V�)�$�bwS-�ݳ��e�a�|T�R��l"�ͬ/w9*�˅�'Q�U����[�I��/)5��|{+��߹�k�;���<�s���z���}�A�?\�'��Ym].4� :��n�j�bB�Ǡ��Q-U�9�n)�7���Y����@]�Cy`��v��.��u�%z�j��t��Ŋ	�v���o�s��ַfm2�y�b����f�s.h�ZWM_$�����C�9���5	y�΄v\���4���r��up3\o��$f�6�Fm`dpޜ���KQ�\|Ukܬ���z�����\c�eM��{{oF$�,����%j�6j�R VuB�e��z�lz����n3ӧQz��������\ŲJ�a��X�W	���T��s��0���(]�y+tp��,Պ�'P5�n�Zou���і���Yް�����3N���#Y�ޮ:�]L��M0��2�9�wr������踆�cr�6.�!O����R���Hv�j�Wi�[\�]�?:h�XK@�y���4=�t�P��\�0��nT谧��ΰ����6���_N�̋���]���v��`���Ъ�8�S\JָiM`�-Xp�(uXܶ�1j�'��֭�]� �)�2����4����駗�:�hY(�e�D�ц��ā��o��m�]��N�p;CE��cvn�/XDq���Y��'{�볹D�#c�_[�b�ZQ�,�f��#rJ��hƸ�ʝH���r�����v��9�Y��m�r󻮗�jy�M��r�k݄��n��6�C^Sa�ֲm���ڊ�ӏZ7$;4e2%Ct���g:���Z�g��mL����OF����6�e��u���[�S]���wYv-|u�u>0��a��;fj�q������b�b���,n�i�9;o.�2�)1ha�8 �'m����E���&8r�H��w�9����M�FE�b&�������n*�h�����RX��zr�b�_c��.�M��\��%rvR�;,v����Y�����k;ݼ��/�9"�X�7���	��|�[�Ң��r�H(�Vg'�vm(�+:�P#��*g�nG]���k�3���+-_*F�ȳ�t��9\��a���>,Uܺ�����=�]#��G����&�û5b��Ģm7\�鴮���P�o�0YΚ�Y��/>�b�&!HL��*��<����i�OK���⻅�H.Զ���b+'P�Ys�uz\��gO�&�ŇA��0���uk�*��&)o.h�Y��p��`h�*��J����z�����t���>�2^�k�5���s�o+2���$�+g7A���u�1*��������E
mg%���!8�?� ��%*d0;� 6��J&�[������Q�����s�X,�t�]���N�!йd��T��k��b!�4	`�!�pa6h������H۬���pX�w$��s����f���c�CEEj�N��6i�4"�*��ܮ��%��=;��)e�5���dQ�ł�
�ܮ�s�dSR���j{joGO�-�S���h�:��v�H�&���ge��n�/�l쇏Wn#gk:̶v���̾����K{Ovn��7 ���w�>��^�8-�����%���ڮ�zC�b���ªAHA��Z��}y+z����<��$O�I*�s���WM�AF�Ӑ����X|f]�Y��R�^�[L�"cs[b�z]/��Y�)���M[	��������yG]��[]�!��k��iP�Ǐ=4ݕ����i�ջ{�M�x2�60��^̾7����c�ZS�w�>T�n^KMHn�Nq�h�������������g@/v5M�=����B*�P0X|����իD��2�\j:��qU7�.�ol�	�RJ�2ROf�9��]ڼu��ܨ�T7�r.�z�� \Q56j�on�}�����)F.��en�L��2VKw��ﻘ:�Ʀ��U�KNƗS���<D(���}�{rm�k_T��������(*�v,T7�pԩ�{�.y8�4��:��j�����D�dofS����5`a�kh��%�;X���VDy�\%�p	��x+j��Y����2���7��)��Z����̭}t�Sa��˓
��F��E[��m�@+��qФ�������m�y��{X�=T��ohN����2-��s�ZUA��ך��"pK����-Bq(q��ܵ��+���ǹ��ㇺ�De�ms�t��ML��{�s�lWچ扇g>P<�;-3hἺh��0����U,v�C��`Ρ ��1��yWL�L�Ý��7�K���C�8����]�\�W��W-'Wuu42�z�9Vk�Y%��7a]j�o���Ur=��S��B7�h�R�m<� ;2K�9�3GmWk/�Z�1ۥ|]f �0W_p�1åoqI�5��q jj��q�7sr�[��� ����x�".�[<�͍�ct�t8@jZ��v#uS���D���dAQ�6���o0�APR�v_*�ұ5n�u{�|.��I
��5;����G���C;x*��ɊM�[N��(�4�F�q�Y=Ԯ�*�Jk�nӍ屶�]G7$�p8���MBSƱn�'�P���v�l��T�Pյf:���W�hEHf�&M���@��G��/��v	�c�z斫��Q*�+��Z� `n�n�M�5�ռ���b��AA�{g��`S������}��ۚNV���"�@�]�Y�\�(tw=��V@���g^�ι�<�ѕ�b�m��>������g�i焌S���R�Z31��}�Eͮ��ʷ.����o�Vt4��
B��PP�M�� 1�e�����c�L��].o���q�wH����J����*No\�&.��!4����!*t����:v6�VP�\�G�gb�9wwٵ��ۡ��f�8�z��5ʰax�j��c(P�\��;�UX�־��U��,��Ԥ�]#٫,�9�Md�wvL��J���a��.����D��t����Fs��ێ$T޺V��ƚ���3y����<m�0CA���;��;���kz�&�Q�����ڔw�f�㏨jTɴ{�zlH�S���&���u�6skON����E3���m �ķ������"`���*ج�)*��;E��V+L�%�5�r]�ɷv����E�XbېۨD��ۺ1������{��wf.9r�ᤵ��]����PVp_A�@�>\	�W�gS7Wt�iU��E+ڝkw�]��;Y�yB�ч1��ٲ��(�}�V.�f�F���q�gc�@��wu�qR��j��E���ޔ��o/b�8.��u��L���6e��ַ]�IiX�1Mu۶E�EZ�8�7vd�i]�����8w��o��� !"�_�@�Hd���C��0=)��w����]��Ʒ���m
�{B����N�K�=:��K�tsN�LS�n�\����/�(��ڼ��hLg\�%�ocw������:��o�P��}�����V3�w}��ؾ;n��ڨ&�mvJ�i6.�>�.���/ G�@��sF��c!�]>�0�6���Xe;��S�2��׶�]�,39#N5�B��w���}>{�b���"n�ַx͠mu����7��a��4EA�K3+�`�bE���b�wP�t�ۙr^��	�p���u�E�Bgok�^5Y�cY���=�v>���J����V�q�ӕ�Rr��"��4x�O�
�W|�nj����;N�J�X1r|"���g;-�-3�Fko���l.��u�|^R���]��#!�w�8��wd��	l���K��-�9|x-�T��r@��$��d���G���H����Fs75X�.܊#f�9��u�t&`�&ݦ�璴�x��?���hF�[��+t͕ʃ�B��k�h�Mu7&4�kZ�d�߆\���piS��q�/s:�J]�FN����e�n�_�;^<���5O�32��2Fi���o���OvfD��7cU;|��k��p���͐.X���܌$ӴJe�LXxGX���	�ֆ�v�s�1��˶�Ó�����tfS�X��\�r��;�Z�j���>=(
�������.0�&5���%2ְ��L��Q@��F-(T
�"�BT(%J¤Q[Ea�D�Y]�*Quk\@P���j,-��2�
�XVܵ�(2U�UcRV!rʕH���E1��r��1��3��TXfR�)1 �Tc1i%��J�Ĉܤr�"�5�WWI�XER��q"[��,1ƙ`�bT����TJ$�(b.*c*F�
�hcP�Ur��f0�1I[m˙�8�)� Q"ʶ���F1��*(��HeVV[,k+XT&"��-�-*(�dQ�-1H��am��@Y��-LLq��IZ�c�¬����c*,
��*A�TS-�R,o�:?[�߻����ՙ�t2C��S�][k��	1љ��)s��h\3��|�Y|s��w%�+�u=@��פ�-��4�ﾫ�ӷ��U#�����/���_��YF������g!0���,@��M�P�nj����,�+T�`����j䎧9'��.���0O!=���K���y	M�4���}�@$rU}Q�$�5>'r���c�����o�eZ�,�n�(�6�%���xD^H����Z�+�r������`�+~:�E$9>�x�n�L,��8�](%��-��Ϝ>U�^톨צ6����9�b�����p�"�eWW�C�U�ִ\ �J���XV]�^u��U��V������Ѳ�_���a�����x<���'���k��э�^�m�����y�pj�Tn*D�1�wr�����/4E�N��o�������Zh����#��`����Tjv��Xzzn�L�����Q�����ۖ4_��x�Ѱ�'���L���iq��5�e*4�6.V�8s�;�['�a�N[)���`t:j����q� &��K�g4�Q~�-�$_�a��xubm���ќ�U���4�cVk�H�J;{g5�+.�Z�洱c�Fگm�y�������Ow=i�>
�Ё���6�=�}-PEM��lԬ��;�IM��^��V��*\�7�]�SNL��g�{�%������{ftm�7�M��p\@qǴ�'/�ĕ�~�j�VN�̌ f�ec������cWKu��|L0ɭ-9��B&):�#�U�|'��C�%;ygǵ���q�����}ݪ�}�Y6�����,9�wP����5S��{(P�H`r�53�Uʉ7��^m>W��@k��vf>H�wM
+i��%#��9n�J�UCe�9w`⼘�K����Vf�9�X ��ʑ_%IP�`���J�Ù �wNA+
�q�e�(�z^�S�f�}�Q��]b>G@k����֨� �a���O��Gm
�}��U��+������_wLE��P���Qʜ�ŷ?>*M��T�_5,����U�c��U��SC3��V<��X�,t�C	��
�;�䠁.c[T$�Gk����T=w�/mx��z5�7�� >�;~��ąx����\�3[P��,1}3��s d�r��D�*oL-W���f&�h��#��l��6'j}?u��
�ݤ �� .�lz�#v�މ�����{ n�خ�4=�`y��EUz���h[�A�lH介=xY��A|�mm�X9�Il)��_Ko���g\O7������X/e ͬ��;�[���d�U5uO����ةJ����M}���22�]���7Qv�\b6ë+:#�o��vH�y��[+2��.��T�٧TO	��knկtX*��Vr���
�Z�c*�8��ˋH��n�s�����K�
�����+���N�J��ʚ�J����{�߅�޾8�,ώ��}`�\��HM�����FΘ*
�.�r������iM��>�6y#���tPA��G	��6�(u�l���zs>,>5=�q��?d�Wf÷�O)�1�Q]v�K>�z]Sb���,�QuQ��\PQ�,`���'/L]oG�j��<��U�ʔ�G{��A��B��&#]DO�J������+q����8Q��꫘t�_jO8�Uݧ��0V��d���R~#��,�/;j6;�ԯ�4�pJ�-i䮴��5��z'<�t.��
�#P`��LH����a�q�$ld6|����37����<�9���}�xS���Vz��dˉ��j�o�zJ�����H]f4��7(ٿPy�WR�~�w��V� ��eɈԞ\J�rx�Z�+��6@<5>�B�d/$i��]"�M��@[�U�P��Pz����E#��G��{N��P���rq�v�`I��2|q��Q��:�J�;W��ռ��/���3��m�e���C�K����Ie�{;��̸o���ygYZ�D�E�́(e|xP�*9s�e�"v~�no�B�HX25[��إ �-+��G]����9b.�
�u��í�_�t�b�T���A��u .�l^@����H��� Lv�:b��7���d����)�Y]᳒>��;�~3�� �ƞr�!`i��Ol�;�0�³�ׄ~Py�o�ڗ]yp���yR�>�Ҫ�%~�| ��0X�|����&0C/')�";�*+,��o.���K�����1K���)�}��;�d8�Zb��������G�1X����l�S���c�ifW^�`�U�ێ�B ����ȊS�o���v}=p�(�
��ə�I�.�n�꒯q�G���_V���hb�Yޝ��-S�⯫v$5��'V>V�v�؎p:3Ո-N�����:�kx��ڞoC�c��fhO��@y'/{�F�k�Lp*��G$�� Ftsq��Ω�ӹ�7�G����o��ї�2��-����)��[y=�c���j��9绹�AS]��<p��ax!vrĥ�I#��ٽ5S��Qc�`z
�����Vd���_-����;E�5����	눍T8 f��w_m�Ep�/v��*wB�wl��%'5Uj-��2����Q���Ӷ3Ǯ�+�8��H�uh�p����6��t֝At^KU�����l��J��\�@�%ܡ
�)�C����X9�ݬ�h9W����ɢ����8�e�V��4P�x[{\T�čw�q�&;�oOtb�`f)5�O���e�sU�&&(�xn	\c/��(;�oY\>�*,��@B��g�f9)� \ޙ�o9_]āǄCeq˙i�dR��7�݃Fw3L_��[-Q�S���:�T�-n���#\dŀw@d,u"A�7(��o~+E������9�h?AJ�Ǩ�j^���g\�Wu9�DS���7��I}��Ox���tU�Pc�����Q_��g�� �e���-f\}�GSy�����W�������3gb8�f�$�1G%_S
���r�'\o{q��4u����r��ʆ�oc�ca]m�\'!�/6׹n!N�^F�t62'��^r�UO�رNz�
�����r:ܤV��@�E��uψ�-��1�s8��y�50�����_�ǋS�%]�e�.�_V�t�,�8d��u��
�K�^�t�%b
��w���h�Iaۦ <y�fC�c�D�4�8�,����mZ�lW}0Z������yk,he7�n|�N��)<j>}1�b@rϑ�>�b�\�y�2�qU�T��6�"o��Q�|(����&h�+�r��X�W�#��u�ʞ���^qJgG���?����x��sUgof��FɋmL�]��m����Gt���#t�CR��}�x��߉C�ٔ?mq���_'��#���q�S�6���E�L�W��Q���1���B�@�]׷3��;��CI��?�oc���NQs(+��;�-q�7	��q+�qpB�
���t���:֊�����{{�:z����%�egF�IΉ��ϰv�ӹF��/*����9z��4My�a�<�gS�7��|ђP�Uu�Ζ&8;���]Qj�
�wo�.�xj�]���>\D��a�Q���Y�!����]4*
�x@H�t	��]����}a�0�vc�mo-������/a��TCRD�%I(!
���ĩ�9�
e��o{�,j��;�+x��c�A�E�t6���*���~��q�0��k�]O":M��7�tߕ�{U�����*:Rf�y..����z9�>K
g�;��+��/I��q���A��mZE��AӁ;'ۇ��`�$��9\-�å����#��RU��tFK�C�jר7m\S���j�gYܚ��T�-$��"dy���W�H�8TU�Ҩ��j�{��N=�'��Oׇ4�C�&r�71p����ˮ�<g~�&�J�Dh�؆9�gW����M�p�[�^�b�!��N%�kj���~z�Ԃ!#��E�����~�r����ݧ��zk\�3Q ck��2�dS����jX9s�p�r�J(�p���0Mft<�!�M�~+)^��6z�����DĨ�Z�~�>��Iǻ��}�����LH:�@X{�@p~7���v��2Z����c.��Hkt��*ց�<���{ۡ5��1��;��N��nlV�vO��uQ;=�+*�C�~�$�{�ij�f��N��;�NUs�� dSck���k�����a��c8]4�Rˀb��<�.�[��~99��gB�����~�m����_ʄ�埜P.�3��l_+��·��ހ�� ?���d�}=�G	Z��Y^��k�����ř�����Ih�.��RM��������<�܍��LR{p�P�J�Аt��NF-��*d
m�V�l�\�uGh�ނr��v-T�����e�)�,���=@�i�z��P�J�۝�c����.E�窇p�
w%����Q�Ww4G��WJ�r�>&�7��:�t���;�u%�³&�+gt��s�����ɤV��x`��q�k�+���]Ƴ�����ȭ�~^󱊦/���.!�!#P�N
���BẨ��"���R
�/i�5B�#}x�u�F�m�ȑ:q�l�j"�Ws:!��&����s|��֌t�V���jWo�=��瓫&�S�~��������,*s���e�����VK��˟?j�6-9���Q�q�}Xw�s�������܁(eA�?!Q�ղ��P�`=��dHqWík�{�Cx�0n"s�g�B����x!�^ͧ��{R�g��ܯ^� ��Rֽ��B�<e,wg\�F��t�|O�hs;��6^�� ��p�#�8�MGu�I��7�黜,���;Ě��q��]h�%��b5���Eo��;Y�i�~��F�R��H�q+�"�����;��c^u�p�s�œ(1�*')Y,�ׯ����Vغ^���@��[�cλ����ㅅaWv�ӗ��Xb�� ]��*SS����\�YjR�MMdܡ��2���t�e�+Ep�/��y]�v�T�q͸g/:qପň;q��y]�I~!�����Z��޵2ot�Fy.����uc�\p^��m-5<�̾�#F�97e�k�����7X�����*�D��KJ�;��9�yZq�.�Zc>���{����GN0�A�ͼ|�]Y�4K�rb�i0َ��\��if}6�eM��z��o�����*~S�Ӧ���Q�Y�!��u������<��<����}c/���nRș��$5P�Vt����B���9["�rh8yc<�U)�Ӿa�[����鸜sOwcD���P�.�9��7M��"��l^uPE_��L�nf�պR^��P��Cu~��4b�g���N�1��,>1��b@�rP�q�Y�ºM���S;}�tW��s�h�ea��,u}k��PP�x\7��ND>����ݐ���\f�>����)��+4;���Z{��X(Ȏ��sƅV��/r���ʤk.$;2�G�6&@Zm��r�c1|&��f��+�A����/ U-��y|�7��@G[��Ry`W�H��xe�+�����<����u��a����iu�ؠ�M��}�-��=u־��x���S��kU%K���O�/u�y��Yc�n�"��zw�e�:k�=�@<j�mu��ѡ҂��C�z�\8�u�KK5:\��H��-f�L��lN]�Ⱥ��/�7���Z�x�⎭y �����)��ڛno-a�^ͥ����m��r���ԀѸuU�q�H�](�܃(F��A����T,�<�]j� Oy(q��(*��3������t��P�ڜ7`�B�"*���h|3ZY�j�-X�����Dg��5P��޷��S���6�hMr�00P���Gu�{�]h���ƌ6��P�,+.�0+� �U> >ܤ .��dA���ÞZ�a6��G=���eؕ�0��}���*��s�y�6���}��H�qI�u̜�志��}r�Έ�ǽ��F���ꋹ<r�e8�:<��O�CW���>�^M���tc�GgG)෪m��a�,C�_5(h��h��4�8���] hv\�Of��[Nެf�Q����)U��x�7�e#��4W�_Lf����� O��x���'׋�a �*>��Z�;���qth����wM���2��:wO"��J�\i�#L�+�e�.�x�&� _8��$�J�̔!}I։ڿ�	�:�|~������>�O���~^��np60p�q�V�q��Ѷ��ua��J��0�8__a���f�� a/1��n+��4��9ڹ���X������} (��KB���h���*Sv���,��'WS
�=�wE}�+8�1R��їm���f�x�۽���ӂ�f��u{�F���#Zun���m�ͬW�M�/i�B�='��%FZ�8�<挾�z\Z�h�csa�,�J�]{��T�-��u�J���0o,V[<_����'��f��W������P}�cݭ�*�oIt�W
�tD�M��%]�<Vc���5��h��Ӽ���h��oG��cV}�U`ȗ]�ӑ�Y��d�Ȥ-?��գ\Z\J��(�ވĘ���ɱ�i-����bɤb1P仈7�Jco@}�2��\�-*��6eg!�<�u��Ux���ME1;37�K'>�Wj|�|�_tMYǡp]�Q-���촫,�*���xwm��0	Zyem�����AK[��lQu[�i�/VV=�χ'� ���j�Cy�n֙ϋAVYջ��.�Z��D{s�[ƖAUՅ��֢ǲ�A��L�[Ί���9ݘ�(��-E��pP|��I4+V�RT{��\J��Y��ioj�	�jJ��X���j���>�2�%�Ø�VM�+4����2�m*q��B�)RA[닩��]�t�ao+o�h��D�WR��-���v=e�b��v�*�X/��[�(n5�+�o���*BS3az?�'�X���,�EQ�-�W��.+ǉ���n`Fk�ފ5b�3w��w"
ȳ�h��t��Ԟ��p��W,��A,cA�U�Lլ�7qvgNѴOh4��/m]����Nc��+���YN7F�^��\�w;3
{�ge����Qv��
�]���W�6ڧO��Rw4ކ�!�f73��S�J�қy��[+��R�H��OF��YsL��舷w��|N�N��i����Ɣ�Q"q�߱r��k���K~.�yҷ��(WX*ʙF��Z�X�v]�E/��#&������wƳ�]ι�5f�Y	�E>��`u�eR�)dk��S�AU�A��\�h�i7�@c�n�������]g0b���2���QaQ�Ig�&�60��F�&�, :�JR�.���r͍ъ]���&�Z��7���vY��\4�����$�Hv^(S���5��/�n�Pbˍm5p���k(��{�p庲Vg7rK��]Y¶�����=d���''v�m�a��ŗX+�|Bo��ct.,C��������h�7��/WQ�d�S1U�"Q�.��Cq7�c�R�:�e�^���� ����(1��yH��K85\�������t�Vmjp�\o�EͽV͛A�6��Y:�c��	�k�;�{�)�Z�c[[sz��7�met���r5��et
\T���_�:���o��#1U �H�H�*��\��-(�aFU�ڔF�`�ZYm�EF���&fei*Ae)E$\�@r��j[`ԡX�R�*ܥb���嫍r՘�J�eQ��+YD�*�T�J"(�kF)Q+m����,U��RVF1�YT��)��U�(*��*-�X�cEW32�EJ�G)�	�l.Y�X��(�B�R�J"���TQ
�AQ*ḙ�1�)�*�aU[j��(b\�)\B�&Z
)[���L�be�D[J���+j�V�6ʈŊ�YU@A�ar�ikeF+R���*.4d+(�R�UURѤj�-��E�Dm�DTX�Ѭ������U2�#U�
ˍER�ĭj�B��F�6�B��}Ό����?u�0�k�sy3��t�2��.�^a�WE���}P�)�%�s��缙��Y7��ll�W
�׋���W@�)�����o�OR<a�g�5����ATY'��ĝ�{`T=OS��l��$s)�|���;C�*��>C}P�A���=���Yĕ���ʏ���H�U����a�L_�]����{��!�11RylRt�gL��g�3L���Y\v�Y��������EX
OS��^��;`Vo)�&�|��veg�z�C��� �O�V�����^��p�]��s�>�Z�ϧi�$P�����c'F}�&�x�Lx�߮�v�ed�����i4�a��}Ձ�Vo�iԯ*;̋&$����q�V�O�g�NُL�ӽo�|�>�]��y�>��<Cl6�OS����d3�8΃�d�(m ���ğ!XL��t�ۦ�ϲOl����^��IP��2�*K�&3�.��xɞX�c�DBD�zx�|yQ�yy^�ߝy�:f2T�~2�>d��`:;�|���z�>'r�1RW�7�d�S=a��p�Ԛzf�����I��c:��$����u�w��4�{q�3�������>2��ݾ>k��y����|j�l*t����A}C���ͫ;IP>M�k��4ɉ�hz�C��-CS�I���|�4^����/���~v�Y��rM%C�b��>�A�`)*}�{��q���}������7��l�J��ueB�0��&!�+<C�b��^`m �O�gWHv�����Y��LC~P�4��*c�7���XV<���R|�N��M�ۯ�B���'��y�}^�F��Ϲ�`�T��>��zm���.�9���mX6yg�k(x��u�C�q'��SI����û�CiY��v�I�&�t1���b:C��3�R�VT�>=��x��yϼ�s}��=$�J�C}o	�g^�1��t�Z�d���biS~��IZ��+��!��N�VM�1'�W�O���@���i�yM�q���+�>c�>�f���l�螸�ܘ�Y��>�`"O_Y����4���y��4z�L��&2=�Y�8�'hv�!���AT8§>��At���w�Ug�+&�zM!�+�vɝ����;Ir��J��V|��[�k�|���^��kF�.�W����k���yc�
����'�z4�q���Q�6�^&y��*+;��������B�~��]E��_~{[f9⪶�j�C_:T%�b����T�;�Z�nu^8�����V���N�Y% ��B�f�λ��O=��t��8�I�@�㤂�y�=d�T1��ߖLH):��4z�0��q��3hqS�8���d�!�1{�z>C����,�18�09-^0�,�Ę�	~u�=�߼b��}����mu���|M v��L`x�P�v$����bN�Bn\I;g�nw�L'���2q$��܇�z��;gf��Xxɰ���$�'��_���=֯��������|�[��i�!��ydSx�AH��q1�M'{�h�@��޲x�&$�T���K��]��������oG^��& m/)Y>k:d�������!">�O�V�}�r}�9�>$���}�;���m%{/y&���<z��SI=v�I��1 �<~M���S&��z�����S�Lg��'�g�m ������#�F� �k^���
�M� �u�{�9��j�$�>=�"�C�+�xÿy�I1
��.�����O����w�7�p�!�vZ����H+8�R��1\`T��v�N&0�q�ϬE���G��Y8vaI�qsb�zz��T��P혝uC�4�P�����N!��Y��*<}I�y�Tĝ!S��}k�N�m
ʝ{�Ci�'���V���L@�+�l8~��>������ �G�����Rǚ�^|ݓ�c�I��'lǮ�C�=q�N'i�C�k��c�qĩ8�N{��;LCר}�z�HJɰ���m��I�*��>�GǏ��lyy�n��i���Y�����;O���(bL@���H�|�v�^���4�d��t["��+�y�>N�0+>I�k���'_SI�3�/��:f�ĕE'����I�DWdq�7��W��Ub�"�D��|bb}�3�z�'�j��a՚��ă��a�f�Vw݇��>I_��[$�
�hn�.�
��+����&��01���z�l�>P���e؅�1�g�-[��{��}�J���7� �_y��*m�W�1P�1�i���6�Y�g]���H)�Շ��&����XT�i�M�|�'h]�sGN3��}^���d��fdb�V���CU(\�4]I�������A���'�'��4h]�S�~��\��Xj022�f�qj3p�_J�R��)�g4�.�]d�Ѹ��ыEć�,�Vq��@9ݖ�r�'L�-�Ro��><a���R|yߚ��+�Y;�{�P�J��W��d�E������fY<f+̡�8����te����8�wC��6�Y��$��ȡ��� ��DA��|��0rz�՗�og^|Aza���N��mĬ>>���x��T�<¤gi.��['Ht�_S��桉�;IP=J�'Ͱ��4��*q���Y���^��ш��>�"!���	J�;ɮ��^�A�F;d�����8�}��i:�� ҰwM�3i�'�S!�qgbg��CL�z�&�δ!�P����LC�1��Ϭ1T;Iw�P�J��cӾ�{מ���n߳z߹�=��LI����ݬ'���|�uz`c��>dՠx����L���C�G��*AT���v�La�
�ߴ!�La��{��t��f��:�P��H?vo�}���=<��]�λ��q%eCi�1�jɝRTx��5`�z�'I�bi�z�{;��W�
��g�i�a^����CI*o��6��Qed���z���v� |��}B>�x���ó]�){�G�>׾��<�q�P�����&��Ă���WI=��0�Ն+'IRx�Vi �@�3cC��b�Y���go�1�]�!�����RiH/]�经���������˵���\�#9�}
�E��Y�>������S��k��`):B����&&�yI�d�SL����%���I��
�:5C��m ���Pơ��g�;�4�@!��D��G'=%�b=��Q��`��6�U<��O�I��c�8��!�i�R��J�:��M���u悦Հ��=��+%����VV?:N�@�z�R������� }��:�
��{K1��{��&�q��>sl
��z���'��t�Y�wO��=OP���ZI�*'�g�aq�Af��ړhJ���I�1'��Zc+%W�����AA��DXy���oU�Wq�����|N��J���4��QeI�<B�a�W��z���8�|`T4���>zI�z��{�ڊO]���1;�� ���V�����N��z6���b�s������{�]����W�R���p�M�5�
F�6��L��곆V�SIu2;V�G5J�aֵ?]Cb��ѕg{b��>�軫{w�:���Ʒ3vۮ�RC;+çOW.<�w����C��ժ-�Λy��p��N��2�p�Fk�9ι��,��v��X��Y�k���hb���2g(v�̲z�E�泧��M$�
�a�=�S�`)1��X�d�1��S���M<d�i������>��w��{�9�=�s��n;�|ּ�Y��Y~�]�5�H/�դ\C����$q�'��OP�1 ��<aS�:C�Y1�0�giա��C�{�x�dğ!\��Rkv�:�Ϻ�^����%����+�-�X�����2lGކ���J��ף�<�i�d���փ�b�C�*OS��;O5f���z���:�|ʚH,�o�3hx�Ctya���T<O�M$�ozSS�Q&�[5#D]�nv�JN0H����g�����t��2b[��8�=~ޗ���"�5�x���9l�O<E��j��;�EM"����Q�/L`���\�h�j�h���a��'�L�"B�)V�e��g#���w9��5N}��t��KfkJ��3�����Z�<r۸�j���h�f��Z��x��g_A�S3��a�,+1�U\��na�N�{�ʩ�F˩�p#,�H+��;/=�ݮ�5﯂�1�m[�=���𰬺� C�����H���W
��u�1���k�}��c�q��UrZ�X9u�@��j����`��Ό}��6X����.�+u�]�, z��k�˩�X����7�g��uW�|��_6��n��˳�K�G;�	%��}Hp�q���hCo��՜�N�8r�[����:q�M�=�*s��z�򼂹v΂0��}`�&��꾽��I�s�f�&d/w��#6:�f�79٭�*���j�R)���j��o.̫�(,�.�o1�
cr��#������D�(p;m�OT�u�3|�Uﺖ�]�K�cQ���g�n[)��Ɗ����}�|!Yw�&�]&:�z^�/d��55��e�5:ȯ�t!3�6���G��5);��F�3l�ݧ��߶�H4V�)s.��=@
ф�3̭ͤ"b��9�_'�{N�y�!=&������� eue�����|����ҾoY�wϬ��֏In�g:�G�/n�MU�������qp��-�� �c�n|f$D$etТ��%pm׭�'��J�l.k':c�~���;��5�`=�ހ"�eHHΔ8ED(:<>�����gXX�y���8��wH
��&k��X���rre�]�?Z�������u#.�����e̭��1IQ��Ŕ��(ewUɅq	S���~lҩ��T�{2�����Y�NK��ֶ��H�fakʌ
�'B���2\�Cj���y������
u��w�-5��e��q�.�]�@�W%O�����(���P�}���)hܠjHN���b��z�h�����FĦ�y�f�ĕ�tC=��ۣ��}QJޡf�h,SZ=�?���,yc��^cq��[��;lPO�t�\Dޮ�������1�C�e�T�i����U�a�y0��k�ja ^�0Ʊ��po����ɭа�����5ٟ�>���Aeq�>ꢱ^��0�?r���;��Q9��.�@������(�t:bC����lӪ'���+Y�;��Ý��n{�'�l�p�\\qP7��'���ݱn���\?bȑ�4e~�l؋��	<�C���N��/����
�����U+<�u�}�Nv>� M��������:��'����3my�
zN{��xx:�_�&tu�o]ŉ��6~���h�e�2];5����)���Ⱥ�����*�������i
ѹ�n���O��/�W7���⊖U�Ҍ�1�����pA8T�ڐ�j	��S�e*�o�<�4��krW��wޯ-Ry�ov�G�OJ�c"�!����?+yp��x�l��i�G���8�U��Qus+�����׺����Tr5{��:�8܁����嫡p�THV	��(�E�o詐E��M��.�w����œ9^�*sӠP��ǏyLy5@�[�UH�o�HkU��
܁�2
�>��Q�t�;Ϙ5�v����.�xC2P ���.L<��:�u�L�a�-��{��Z�yr�K��_
�$?��i�����}i+����ٸ���p@3�WC�"b)U) D�P��;�M�q6m�y��p��J��G����,B����fcy���[��9����sf���G�5\�lW��G����JQ���M/�k���̺��d�HW�&���Opfoqw��wK�T�܋�p�����w��]%�9u�*�a��<��
��c2,f򮫻q]��-7�,���*�B����6`	hI� u�cnxJM�q�=���׷���\qb���lP8b��0�,����	�;��_@�?p�gk3� ku�:����	��q8�V5���M�ia����D�e����r(���<tV�����,��Xe�+{�V�ز���+,;�Mh�GgE���l<7~C<�n.eWl�U�]��vH5�q��q3�+�jg����x���[@ه�a�Ԕ!��1s5�&�@��]��B ����s5M��	Ωi��csʹr������������Ү�cY�	�9i}��U�է'�X�/8uH�S7���ױe�HZ��AP��]h+{�Y-A�#!�:����ISK�h=T�T&�	1 Xv�`��-R����e\vј5�]ʷ���+g)�t�,d�G:�
���^h�v&��D�C�ܺ����4x�t�v"�:�䓷�}�7]���d�>�{j[[�"�����k�ˉ��͉(%7���bu�+�G"���q���\ۭj��Pl� ����c�)�M|'$_W �*��)L���te��ipO{M�C�zv�H�->�iM��?!�n�G�<��e�A`�[#�c�3͛��ݢ֑�kE
r�F/
Py)�7)�Fql��0+�2��۔l�39��6/���]26	�{F�,j��񢆳������wB�h�� ��'��"D�f"i-&�
>ӓ�T�|��i}L���Oi����U�X�O@���ۭ��]�p6΃֩ �fD��,�1�:M�0�>���C���[u����*:7�<�SQ��2,C��4�]4�j@�jb�I�KH�F��6�H���k��Ut���D�I|u�F��	��L:I<�:Ԁ���#���I)�zp�#���ѝ���IX�L����1�b���q��zL�=��3�]0Y�}p�{w>gjp�K��N���c$Y�J��9	."� � V��nz����h�+�:��v��+:�d��V]ׇi��2�r�=|�֕�7�4�wF�vc[Nu��s�Ƶ5T+�w��y�R���֓t���d�C/*ww+sBJQu�[V{v�W{ﾈfK��潱 V�}��tmp�beEa�w����+��~��B�����Q�/靦S@=1����ò�}��b��n"Lpʜ�B�����³|@�eV[�j��*Ts����s;�N��M�Sbn�m��/�*3����G�����R�s��ς b9N��``�ܡK79�Ԑ���T�	ݲ������c�`0efu��S:<��R��H�-jM
���uf=�͘(���7d�����8�a���${��ٯG�ŁO�:���<zB�
���x�l�������1jc6���7R�G��w�Smd�P�D��X���u/{%��@�ː�I`�"��D�i�>�c��;��N_�%�S&e��ە��Ԓ�!�.dY7A|Mh�_���]f��y`�ͪ��[�z{�P�[Nڌ�l�Z��j�Cy���ˌ��%uR k�GI����h���̞��F��=��Ε���f�h!�ur9	� E��0S4����f�`!���BFc��@-�e��v��Ȃ%.��Y�)�Ks:�=�K�.�����T|�}8�ܽ�J�b��^^�c��A1����@�֦���}��=��k��R��H���M�p��,��n�w���JjJ��C.tζV�7�Q���y<�>������5���uQ��~B~\�Ȝ���A}Zbw���R!����8EA��&��GA-)����������7tq�6K�\���>�,��\�7 wB{`T<�"4�	�h?c3�{UN}=�L�������$z�v�=9�
�\h�]��\�3��J�@u��S�y���޵[�[(���F�cM�l�V9�^�,��<<뺮J�sD(���T�'�g>wݏ5��|c@�^�Y#tٵ����,0��F��f�Z��[ĝ�qwd>27n�Q��j�m]�
,�c~��'�΁���5�m���r<�v��kwӂ�uz��P����\0��G1 ��lF�:'��p�f/���J� Cw����V�)�{|A�*������@w�����}��������F��.̽�G�f�F�:�.��֊z��v}-,�R��q�_f���s�z�i���.?F_7�ݫ]��o����I�|*
�-y@rS|��88��ZX;fbGo�e#��ۧ�|�"�^�.�
��_�S�W����-�����kB��ٚ��V�&T8���l��ܚ+�b`wO�7(���wҢ����]���Ԕww�M�Ժ�����{���*�'�&*��]M�Kb��o8tڙԍ9Q������>Xr��R�"�4)�s�'*��`�7T�q�X��w����S�Α�6�c�Y�-�*�9Sww'��	��a�:@f�37R����X���5Z��|�*zjm�Uf�Y¾骹_=��m�z������
�[�7�Lv�U�h�e����β�k�v�[j��e(7��ښn��%mD���,�ͼ�}��ڦ�
-�i%�;_J����\p��;`ы��ӯ�m}Coe��Z�yt���b��v�tjd,	Z�O��żh�=�8wn��7�4eJ�$��۴�Ǹ�)��+�xu����{����ƥ��pT�i�[����>P�l�oN�Pv��*��~���{�.�i��ms�m2`t��+�*�4�wl&��v�-3��Pf�bs	�;=� �z�.�@M�������^�f�A�>�"�pu�In6:����v����PW���5:1|��Mi�|�]�덅/8�C�wWͧ�B[�Ȯ	쩋6���uw���Wc���	-�ttC�l�0���7�]ҊA�ܸ���OhA�vf�����Z�"u�S(%�;əX�;���jS�3��xh�tl".���[&{Bjө��lݪ+S)˹G05`5VIT�x�L^TЦ��]e��}ԕNp��h!�:��!��MgN�6�#�����&�ǲ�!l�YR�֊[���A�e�m��f�u�)=�k'�I!u7�kIe_�+�+P�����R��	 ٫���c
���(]^t�#�6.��z⸒��k�BT:;Pi�8u�`�r�  E��f!������]���׳
f�L�
�_u4�Zy9T�T�q�����x���Û�㴋m�5���[�p��&4p�.NL'���}��ߛ[Kgq{8h��$�U��t4XOWb�L<�ۛ��;�i��;�ً�� ����SJ�1��/R�ʐ'�Vޡj�9�W4#�J!e�k3q!af҄*S��;����;]ݸN�N�EBj���-�
���b��Zr������kD��]�Y�P��;c���ȯ�R���Y���䫬��u5;R�	�{��&�ZV�`�uL�]̫�ס��5�7��]{�ҡh�����5���u�r��zVF��^!𐴁3�EW`EÝ�
J��D��#m�[3 �ZH�[�Q������R��������ۤ����@�ֻ��*��q_/���:���H���'V;҅)�ܮ|�5g9�R����?��b4oY���b����Ȣ�r�Y�̬�mk*���Ĭ��J6�*12��Q ����AE��h!l**9J&5jUJ	kh��EQ`(�h�e�mal���iZ �������ZUam�J�kcmKJ�mUjбb�b" �Ze�X�6Ղ9J#��h�X� ��ֈ�&6��".2�UEQH�"������m�%mk�PF�-q�8�R�V�dZ�2��K�ۑ[eU�T����#�kE�`����b�0ATE��@�UTE��PmDU1+��2�+*�1J�U++R(��R�ֲ�2QDh��iF��U�m+TT
T�J�h3��Q��TkU��Z�-��҃Z��cR��AEA\�����*dTV*�,ڕ��B�
���"e%L�E�*�QT��
V,c����<�+���;�}�"�ۉ.fgt�:R�5�Z�A�S}φU��*��vQ+X�7I�\6
����Z>|�o������)����;sj�m���B�
�:�����U���0�����~2����.�0�=�h��Ѓo�q�e���w����6ԅS_��~P%)��<���5��;$C�AM�N���{�o6��2������#'uQ�(�t�t`��1��V����5}��y���-��0�_Y�?W�)�Ga95����j��SuQ!\w8j���]��,���V����Q�˘.S1b�7q���I\M��l�1�%��#���Sm�Z-�����ٮL {h�J�o�T�B�ʼ,C�jV���nz��FÙ��h�7`����O�����U[��~�+����z}J?��^&'�]Q"�KӸ
G�@��נ���i�W|��X�+�.��H��4�� yՇk�ƇΨ�}u�evn�y��<����nM��L1��@n�R��� a1'LT�p���B�ݬ��*G�9���yS���T��+��R�l�,�c!*�d_�"��M]��6w��j�Y>+�<U�h��q��kDh��|�x^;���Y���(R�i�֞��T��_�zO@5wu�t�J�QR�u���Sw#/������B����()�y�5-�/8��q��ٯ,]c=ZR��ڃ�zh��Iy���+_P���S���6�nH����W�}���73�$��uԵ�MW
ǯ1�	�ǕY�*O*�404�^����8i��bF9��ٙ���&��8[�[�s�o�:�����s�v��TB�XlJ��=��fVTtoc�Ɨ=�آ^N�,��=�D��ZU�y��D^�m�f��&�ّwzM�drn�;�a���ϛ�C��TQ�@�z$ňڙ��|:�N @�J������G��Z�n�d�pW{�j�|�8n}N���V_�/����OI����Q��Tt�B��g���
���K����D�?tj����c��:yj��ͅ OW�tsء�h����{��H�#�Gx��;MCO�B.�:>C0�C�B*�ldt�VI͕����Qհ�c�$
 W:�vP���(p\tOjv���W3�4Fj&C�31}��^�r�\#)�JK
F���=F��{D0��c��]���޳�����r��wNJ ���븜�H�c��@�x�t<7�1��(9����:���7��B���B��w��6s$��(u��;�g.��(\��7�U���1ֻBGr9Wi�p&��B��L�[���Ӟ����'������K/r�ӷ�dkMr}�x�L�:{�*b<�W+�����ʋ�L�U���UV����wM��sf�hVx�� T�dH�Y���l�:�T�T��kB�/�u��t���VZ�溢��B6�1m�[8[`VʮU ތ��B��^l��f�SY�n)�w����;��I�L�:�+E٬'�b�b"��6v�;O$�����p��mAsnx�߼ϳ<QOD����1Է��E~*�)g�x�H���X�TF7t�uP�؇0�L����vt��ϨX�=Gtӣk���<��;��S�\͞���=�F���iw��V���t�ǋZo�q�5=x�`���n�:��xAaY� W�����'���q�f�rt5%D.�9.�oԽs���bu��e#�}��@��\�B��C�e�)���=�� n�n1������R��]�]l��n�?A�i8 F�Pó#���ҵPzt
=���V�NnW������s0Ug;L�!���p�ʯ{-�;x�C7��՜ze��{ba�� ��+ҭ.?8k8���c��+�r��Nc����Ѫ!Լ�˨lW�͒�fݛZ�N����{ĳ�J�N3����t�]�W�w���{���|4�9qG
���Q�Wm�Tc��\c�Ai9,�gKQ�+�ؤ�P��r�L�?��cn�����;���3'ϩǧ�>�թ��h�M�~���>��(���s[�~��t�Ӳy��&�Hq`�Ncz:߽>��}�	Us���KM���tߦm{�d�\f�_�4G��Ī!7�H8a,k�~�\)���J#uި�G�{���ޮB{N�'���1������vS$E��]r GW�wo��:�Z�+m��ak�{����t�#�J<0E��]RG{�W@G�*]�t�)n��sf��9z���7e����?!˺�vUCf໭�;�S̩�RFt��l����H�\���e@���%�Ù�<��Y���}I�p�fٙ=��Nr��	�u�`�Oo�K���`,�n��B-�c��?b�grC*:h�Uʜ��g�7�a���p�v���3����Y��r��},�Ĉ�U�b¢�I��y�rP��H���Bv�-90����0��l.���I�7'������Y���Mk�v�����tK�]Z���� <�����U(�����o�ϟ �ʬ΁���rzo�L@0Au�m
�L��C.�I��W���`V	/]+G�,Ι���\��b��2���;hR�OV>��O++,��c��T�����}��c�����at�sզ��Aw�L�u����Ɉ��zu�
���_3s6߸5����y�,⹘�Uj%�ۿ����>�R�9�X�=~�����@�@P�Ǝ+���:�!b�u��J�8Aj� έ&Яn�ťz;�ת��Qv�b�xV�p6�;��B��ǐ��ÝuD��c�y+�_�ć���wU;�#(���C��'g����4�}X�����w�q�9c8��K���XY6�����.����g��PV�k��pQW��D���Kϱ�ceY]���X���? ��IoUU�v��7�'�,�d�����5�@p֍u�蟜C1��0
����[xl8�/�
\cxjR�eLf�
����S�)H��BsՁd<���m`�=�k���<�P��8�7q������.eJ* J@���%h����ԛ
���ۉ���A{:�܍�H��?iN��7 F�m�*p'39��Μ�T#���I��側\A�è���!�w�I��&7�:4\���6TmGb{=}��:�;���Ǥ����R���=%�.�����!�u��=Nc��tt1���~��9����5�uv	Sɼ�+�(@�+c����^
whw'Y[]��SI2b�7��5&MV
YA>�9^d�Wtqu����-�Ҧ��ކy�Jgo��;纫O���:>�� K�w}��{�(��;�Ͼ�������'��K�gL�ʘ�P�\J�.�R<Z�./I��A�/ˠ�_�������l��{��h������}�C�S���!��%�+�%��Sns�nvMD�J�mD�6���-��"6_�Z0RVi�&�mP��.� KBN���x5cnxM>���fW���j{��G�Ok��4A�	��r��5L�"��F	j����ØC-����L5⡛��ɫ��H�ӝ��k)Xx{R����m�J���Ox�u^�p��<~U�"a��N>�<ĭvW/�,��P�%�";nX�,���n}��g�"����j.�~~��)����~��6GꀱX�)�~ ]�T�
���p��'g��J�_ -^����v��ˎ�ݸ�V��� 5���[�횮�2��z�F����n��L&k��P��g����sֹ����q����ܭ�ȍse�c�;!���&ݬ1��<7������/���ٝɖZ�=�Y5W{��G2�Og�1��-�c�)�.%gZ�)�"6ԁ< �S�=p4�B�/P�bή��/��y��5��:�`9�l6N��T�%L���2&��UmMu)Їk�Or�w�Os?,:���"��n�78a��4��c����n'�_CʷG�½5��W�؂:�}�)	�7�}��D,L��ʍ�ޝ����ﾈ�>���0�Mƭ ,�DQ`L}[Q5��;KO��L��a�̡�;B�':ũ���ŕ����� CT���I���r�F.0��q�5��F3�*�mq@�z;������"���r���)��*z������/ֺ�=�[n*Q��յ��%C���Vt8k��s�3�^DЈ?J�Lu����0c��Le�����I�v�d�72ߢ�_�g�H����w�+��� U�W$��?j���kR�:8�:�N�mc�����K��=::�*� +��NH�!���"9p�v���-"���3���{�9�h?AJ��{sG�H�uU�B6	-ً�x�,�c�[2�כ;d�X�c���[��W❮fj4�����Q��L[��u� ]���'�����S��0�K68@d��0��Ʈ�?���:�^;u�,��P���@K�r����V��O<���Oi"8Y��7�/J��8k���aJ������ڎ��K[N�a�<N�%%~>|�ǰ-�}*P��bt��/���f�p��Ӕ�� ]<g�3/��]H�㻤S��
[ٵ�m��Փ�����1�6�� ��PdޝK��������o�M|P4�3)c���{3���nvD�Ήo���}�W�U�é�f_�4��f/H�������.��΅A{af�=g�m�+���}�^$n�Rf�� 3�]��q�'��;�]�E=��.��_���d����!��V�H�*���v�s��'�"�GP�nɋ�t�zaƩ��(!ca�Q�ٮe=�n�v�T�S��\O��o]ü�G���#@Ҭ��2��s��M���n��^�K&46�q� 9��y�\9�\X4S��Z:�w�2��.�!%�k6.u�z�tSk��ӈ�.$�s���0�m��Dizd[��7�xsOz�v�[�����i�=.��ZԮ3k�H=�_?�g�g>�jጃ�����D��UH���G�޽��P�����*ۏ�6���R�)�q���"�쑂��d7,�.�C1�U�$Q�k�-�o�+�7�/��7pO�O݋���l�S��H�dXRzH��eR/g�lv.zlX�`����zw`)�ӐJ�\���>�b˛��yD�*���\ٳP�lC��Bgq��a����4N�t�8��-�W��"��ͼ �R�SO⭖��"�.�谈P���J-�ݔ;�~�j}[\2�*	Eې��v:�mJ'����^�Yך��3�����G��Aol��.�{������'�>�����_+�����L���~qU����R�D�2Wh�}�}a?;>��P.�q��>'��Z/Su�*�XVX�;N��nR�����&}\Q�O{�F�o��|c@��e�����{���B���1]���Ȗ�g�=[o[��_ʣ@�)���L�#���絶��ϕ>��9�8��ZmJ�+s��cǒ�V ��e+ߐ|� ��ܫp�]����]�N)�	g���uE���I�:Z#��֊�k�,�,U/�}��f��7f��@������'!�T��S�ښ׺��j#,���p�������*�#�mb_]g+@�b��q�I�ӛ|����\Ӯ��>����]�Ι�+t���� �L0�}s8���j��k8�b����FMw��r�??��O���ꌴ����Z0W��uM�	���ѡ=��EG5]E��r���������t�/�wJ�/�.����Dq�|�4蚬�_(�"��t��E;��U�F�v�\�T�n�k{9�<*Ԭ�ۭ��];Fkl�+oo�g��VrC��k� H��̅�*��3�q��Ji�.���俯]<Z���B綛�R^�~e}�pN����8�K��z���f��� �7٨��%ջ�?��>����JS��{^�&� �0�y��B�-�CA�p�q/N�4�G�wPŞ���H�
�GN�Y�Ψ�NwD.ءz��,oݝ�{]�H�}�:�-�#OD�yj�eē��f��Vgv��Q"��F�AR�ňC���j�Jbn"v�7�h�#7�s��IP[�O.}�h���r���w�WэR��I|k���p}��ѱ��t K{��,H�d�3f[j�]w�R�+́����Q����]������9X��Q�O�,�x���X1������:T��bG ���a�+����MV����>��z�\�aj�{I~+����.4莚��0Wu�B8�ca�@>Fd1��4$����
���Q�ȕ ���J�az��f���G�c&5�2�Ī��jb0538�N��ɷ��Y��_��;�L�Xn$�nlz�NN�̡��1�w#��2D��r�jx�^�]�:A��Z��(ۿ\�վe
ܨ��|�yO����}_�\��k6����:��M��������*쬬��#�ra�$�hk&�Q��w�d;V�(g1WdYV�N��}����z���RM�):G:���ׄ����+�	Z�9��5��1,d�2������&<����}�"K�<�0QK_=��l�9���}�^ʐ�g�ʹ�\��F�=f�
g�ա�nb�L�������x-�]NQ+*	�T��V�dۺk1�p�t��vl13kb.�Ш�i��"h�{w�Y��5a���U����R=F�|��v�.�u<�l�v�JM*�\z5Qc[�iY[AuŘ�a��i6e�72.U�8]um�f��݊aζ�����>�/YE5n�8V��tId?�n�x�n�Z��p�A�����'UHE�u�{�U�.��uv\G�Eo2rũ=�;5�E�O1��X����_'�v��M�t�E�2�K�Z�K�{v/vv���2�Գn�/�|�/�����t���.`=�g�F��4�f+XjV��x�d��..�1^R�2-r��ë3]o 3eV��S���i�T�����<��t��Ӧ��஡�Y���N�7x����goo�R,x�1�P/i�Ą�ٹ�M�kk���S	�T�{���CB�χGe��P*��;���׃`��Gg'%u��.�@jY����N�Z#7�v��܌���e)+�ɚ0sU�@�V�����k����j��t'	��1p��4�틤;G:�9T/Ӓ����w_IS9�FU�m/M:�<b�����]ZE)b'O�GW��Р�K�V4�XXS�)��V�`���V9]�[HL�u^II+�ĺ�}ʁ�FY��
��-���V���1�:5���9��o"�L:�<�2'%֟ݷ�5 �4N�r�	���L�;��ܩ�U��ĪmE��
�e�r�y�&�6��C#�̠�Gz��Ѕ[��Q:�Y�}��E�b,y̺��t"�=;(%Q���&� �Nss�Q��օ^QA ���J�f��?���$�M�ur�f�E�ժ�7-ݪ��c#��VD���I�+y�u�H/;�f
��ћ"2P�j.
�wJ�DQ�|�n�-��ݗ��\�\��ʵDfP�qq�o2�����|��D_ٮ��;��	X�^�Qb��v�����vȴ[*�nvU���b��+�21���$y��x��b�Vك�]�}j�<wufFb��7�1��e�|���ϺWE��%/��6�ӣ{ې�$$g�g�	)5�E��ƶ�K��ze�F���aD�TW1�N,�+�o�:��Z��V����R�q�]��BppH�v��۱R�uIcli�2���g_N0c=J��i�8�J�ATXcX%�QQ%E*��5�eS1�h(TUTF*��**-�Őm��R���f
cQP��"�X�Ԣ��*��#ZE���C-��\�)��,�-b��X�YA�3*�-�e�aDEr��
�U�V�9h���X��e��`��`�s
���b�&R�D[V��DDB�2�ʨ��Q@E�2,�ZR���\J����Z+F�1*T������elJѩTTQ�+UV$QQe�L�X�Uj`�QLV��`���Z�TĪ�б\CEQiJ�Zm�J،���k1�-*��"�ED�������EƳ2�6��LLn����������&#�je)Z���1��1��U\q��
����B��"�nw�Fo)�ڐ�=(�(��{}{9�[|�싕
37��}|��Z�W�r#Mn�;��O�o=o9�֌�e�[���}_UW�U����H;�v�
�����_]+�ؼ4�v]#½�W��vx\d�1Q�@���\��s��26��BW���|���<�\R�p���(����ňڙ��|:�W�=�jf�H�eݼ\�������1�Ζ���p܊t��ʲ���������(%2#�ƎVsVkj��S��$.53��s��;��!��c��*U��Ν�#I�����Gr�5��-;�)8�(s!��"b���v����>�]6sO�n�{(G)�a�A�*WN�۵AkŽ��%X-��� CH�R$���NPh��:��O'i�/��Ǳ�^e=�����^L�
����Q�:(d<�?$zH�Y�e�� :z���R�R����ø�i�qS�>������p �"sϕ"bh�xL�f���ħ->o{f�[�FXOg�a>�P9d�Su�52��,�0�� u����]vv�j�����L��T�J��a�D�3L7�L�-�֕@��� }~hPÏ=H{�j}m�+�'v�Z^f9���7r⎭��['���x9[y� rR�{�\�E�L�6-Z2�V�n)�;�_�]?v��er�=EN-���ĝ�<����#��L���/�}V�*����<�3�U�|��w�㏳q����^�˔*K��Z�8,�8;'I�38��ﾪ���C���Zp�E��������l��/K�|c_L�I:�/��f�M�ǲ�����:�=�O)��?�J%�A�#!�/�"��p�<=�$��U֓Y��w��z��P��P�ʔlh�6�i�F�CWg�V�W���YP��S�8�=��^'�ݻ��v�n!Ǽ�11r��,57��1�m[����/�p�p>Z�@����U6�O�� �T����c&uψw�]���;��e����Ŝ��&]��MD�#��ٱ����:�};j�7�1n5��2�����r���`�-^Ipe��Y�n�Ŋ��GC�U�E��jˁ�ؙ1u��3���Ȗ#t�R��v�͊ش];z�^����D�K̠2��,%�,ƣ�]V+`�Xi�l�\��-�]n�NtR��9����1a�wβ�U�� 9H�4�sH�����\�*����r5�hv���R�3J�P6W{=�[��n��5+&����"8i:�2�i�U���X����y�!�3U Nnb�v�uKƥ�|zk��KFu��N���J̎�䢲�tۊL{��=��m��[��}��Aܕ�r>��0�P�o�B�TGd�7Zv�#g�e��J�3l�ܗhx�I.Ys������������۝�̺��V����Ϸ
Ü� ��;y�O	�G����2D��(��^Ļk(=�Ƙa��T>����*"S��7+�[�#C4��嚅 5w��Tf�K(��tEqt��D���Z;{?1<��&�T6n:^_��u"]��fTs
{��^�V=|���"�!��
`���N3� �wN��ܝ|�L1���rf�n�9I�ɸ����-�*���Wd�YU�6Z�WSȅ��U5w�X<-��t ���!�����jҝ�7g��=��]@/r�: ��7[��X���ں7�5��l��4�|wK�=�Ktc�7���`ژ����
�tC@Nḓ�v�~tn� �+6�t��\Kx)Zw�`�r/T�f�~@�����dtyP��:b�u���GL�v�Ƕ"�f*R������
�W���1!�R�&�ܿ:�ܫ����:bA� ,�V��K�=Ƚ���&��6;L�kE��^�\���T�w��f�0)�fmw?�{��kv��NV
U4 oՔ�*Iz���{5-�]�e@.�*�#힐�+ �k`��P���]/��Z�G��η��������݋�����iΔÁ�t���A����Ep�J^Bj-��62{8N�h�ռ�z">���{��M�/{�:_��X�E�!��:<�vzZY�� D��~��V��@)�d|���nEZ"��RL���L>4��/.�f�@rSu�QW��Wά�מ�wQ�U�Gejjun�ۄ��Ȧ��S}���A�lnJ���Z�-ez�s�=��ݗ2�(�qT|٪�b�jt��(��"^�/�\Nkvi����byC���}�<M�ㅺ����aK*���������ܲQ�Y�Ϩ��W_.o1wErB��T(�ꅒr6�.���*��*E�z����{*�@j��tv��Niw���R��2����y�,�~��1W�ʲ���A�s��ב�Y�����|��/	\�)N��q���C6�C���M�Y�k��يbV��Z� � *]�]J���[�/�U�ӆ��%)w�/w��}���f���.
*K*��@��`��{<��Ssh�y�GX��}�uԮbd�rh�t�U�m��N�ү�|uuj���!S�uJ�=����W���W	�U 6i`���c���:F3®P�zu����`['kq���v�V�cGµ:Է����؝T�g菾�����{v�^�zm�W�'�Yuچ� ����o3��Qչ�^�>�>�������b�c(��z�\B�.���N�D������dS)=���W�e�{��?~���:��s����m3}�s����*[����+��'i����a�|��bڥԽ�uK�xOk��n�nzx�������*�d�o��p��/gu^!�ҩ�{�r�Ry�R����N�)����&�r���fn޺�<�A�z��8���O������&�T�s?y�ѭ��Uw��@���SOݬ��Q�3��,�:��m!8�}��/ze��v��d��y��>�7'��y�t��gP�%
�ޜ}�O��qj��va��P��@���޵�tuj|p*P����Gv�o�����4c��v#��;�r�[��	�z��V�oq�;���e ����BR� � 8��X2���B�n��;�;4���Ǵ�2殭T�X�)�d��q֎.Y����r�6U�8tr��s/pv1QʽO��Na#����\ �ݡGxx�n��k����Q�j�F�\G��U��UU��.y8���g���������	HJWL�}v;yQ�+�D��1n.�$��;��}��hOE��R��sj�U���K<�uIUŔ�$Ro#y|rn��,r���[��Zy
�a��H���Ͷ���4��jm�����Ky������]�&�j7Q�joySK�p9����cf>ـݝ�A�����Xm[�W=�UDrf�����/&S�q��;v[�X��4DŴw��=&i����|�ؤ=k/]%G�
�D��F��FGb���6�|$�,��5�NҖ�T��"@�Z$�D�;�M�ɸk�v�ʊ���M���j?�PO��(	��~�Ӓc���{�9sꚽ]�n�h����x�W`��۪==i�㈨���)�{.�6����1꽴�W$�S�ڞS~^A�='k��50WO��^��^?]�^�n4s�t�.V�W�L���ڤ
�*�Ɋ�-�����(��r��}��C����=�jum�BnԚ�wKb��l��7W[WɅ�ў�۸F�r$`���C����N��d��'�u�u6�ޘ��[��U_}U�2^���Z.B�މ]?\��6��oToUe����U-���cv	H�kRH���C^�z[߳�Uk�m�j#�Y�)`H&;[l��\���So�oV����C�07�Ρ�V��^�~<'�@N�5:G�]8�)n�[�[�JՋt��GF��ݢ��\�&7q�����mv=ަ�c�J��[�FJtݎ��"L�Rw�ۭ�n�O�ҍ癞��}~�Q�^.��QO��Z�e�ŧ.S&%L�"�9[Ö���7�n�veF'1˸����ގ���;� �enyֹ_Q����0�D��y�O3B����s|���5B5b���r�fiq����`���훾Oo�J�htev��֌/���Y{:�q�M������y��JP��c6����ޭ�i�Q�Dw
{��;�iiE��آ��C]��wR^��+�5vbO�GE�el�"-�7 k.ڃ�M����$ȝ�h��5AR�+kJ�G��<�5�h<��;�<�v�%�RWQ���}�GЩ��ە��>�seZ�w�?7Ы�r��l���ۨ=�9�9b����2h�����ĢMݭǫA�ǽ-�.��z2a;�VkP�=�6�0O8u���;i��f�'����dG�S�Gk�*��ټ���p�ǫe	w
�tq�^)�}�z���S��}Y��GR�>��7�<���3�11�ս�K~絓�.�n�+�HG�ņ5gx�=kV�u��"^��x�������oD6����_�I�˽�syo�����8�y�1m<m=�M�D)�ɸLm�ЯN��+3P�t��5A��j_WS���;�V�Ҽ��o��(N]�,�z�ٿ��y�R�J��&����Ok��Q�o�?Bv��^r��3ݘ�+�;n BR6�F�
|�\b�\3�O�ێ�3��b��t2���jI�wi��j���[:#�bj�zz��E���Z�uu�1@�M�36ĵ]�5�R�/-m�	�M{��ol�^��},�U�{Ί�*���^���Vp�s����:����[ܣ�"O�2�H�n�h���͝�(���V���}�}Z�+wSy|��)�5jWJD$��{T;]�bs�b�o_I��*�d�+n�[.3oGZ��ٕs�Ivюu��V���U3��������mP��w� ��a��9;0����
يa�%��ZI��]o8띜��b�n��'G�ơ���=�i������3#��gx �����������0��k�&�e�j\)�H��ܘ�ty�+�z�VO	��(󢽔�XĻ������h�&L�o�ތM`"��`o����$���?"!������X�w��z���n�z¾��T�Sy�WCz2�j�֡�PWeAʧ���+c�rq.`���L.�2��d8ם	�X՝�_N��-3��>[Eb��j�]M:ͷ#��R���-k�{U�$k�����I�1~>�7qrA��7�l�{�V��2�n����t"KN�e<70M�R�+��\���k������߻��u�
���.;�4����˾sF+�ĕ�3+o1g},�v'I�TEC�u����pu��Jf���u������Y��菢"���r�W���	��&�=˪��z5���������� JS
��V$�9�})o�;������d�HN'��t��}�'�G7��⻪�׉d���
L�u*����Z�׽=�ǣ���x�X��֦�s�3���еB�
7�$����1����{:#�=�_�x�He�����\�I\�U�JBS��ϭ��grZ����s=s��ܹ��q:���o�\z1ܛ����sL�2@���Ó�3v[�.���Ὑp��]�kv��O!S�3�C�,��sv/1�9J/qsۺpat�H���N�B���[iW���N�����qW"��E���/�W˓=�lt�<3��j���*�93Zke<Xs.�̄���imE댞�h��������I�G�1r��.����B�kz��h��un�
����7�����Y�]�:�=�����/�b�<�!��ӝ[��^NX��]������n��F��;ח*wR��&9��pi��0���Gg&��tQ��h��ܚ�aWʭ)ʦ�V�b��MzX�5���[�����ۃAҩgS�\��ʍ�r�ƶ�Ѻs*p
%��U�$W����_<��V��T'L�Y���3k�w	\���"�g���p���1-���\y�<�!�ӈ"�\�t��b�V�٠J<� �~�fb��U�-�V�H��Џ��s�Xj�n��B��e�A�>9{�5��w	jBd�Ʈ9,��VqMTsD���r��Gz_�hGPż��.Y;y_-�Q#��7��ݩz�r��G���yӺa���(9K�5Ӝ��:���-�k��x���V�Y�.���p��]b��P�n������_8��]얻�9!ŵ�׍���N��t�l-��Ἦu4���so飫x(�j�8Rb�iC���@�4����#C�d0;*�7oi�W%�X���{z���A�pr�4�:�ާN�9.��r��jk�u;1����5��ꮺ�e�e�%An�����r�NKqmvo*�)<y�deWrzc8_T�~�m��m�W������,Į��T�D�/�{e�)8��fߎw�l��J���maAcf��ӑ��Y��x֣�r��MaeK_B��<�u]H ��B��z6���Zڟf�[�9܂��`ӕ�%�v�6d}��D���}�V��C�� k�Y1*�h�t���G���ۇI���ҟs8�%e���z��N;{���<
��z�U�fp<�Ԕ��qr���eާ}]�D����c��F=.+jF���T
���u�)�h��f�P�H�U`C�+���[�؆��PV���	��+h�u1*Ӧa}m�tq�T�rɩ�;��y2{��攑�3]q�Y��49�R��v�����mt�C]A_%q0^u��ѽɉ�0l&��ۤ!W,�9�pU�7bpR^qwm��R�t�JױZ�йhx�K�����S�P���nb�m���-��㌦�QcS��u�|���fbd3�c���}a̋镒]�[K���L}/�����Vນ���J�q�W�&�}���U�Zt�V�
u�mujS~)ws�%C(�4���,ݏ��I:�ǐ��z���s���{oU��t�+j[�j�!s+6�a�6�Luܥ4�e%�F�kk_C8Q�ܘJM���O,��RR�cְسOQ['`��0�,�S��gr�T�P�WwH��u�z�>Z�Yf�.�p���atv��T�t˧n�6���q�n��̩4c��Z�[/2�a�7�wv����ގ�=��u�\�)8�}��&�p��מy�m
��c;���%-\pD2�[\�Q�E�V�IYeJ�s�U�e����jf�J��,YZF1m,-s1**�DDE�X���E+ePU�Xԫm�̬T��Y��F"�L�b�X��V�e��VcQX��DX�Z�E�UDX��QF��%q1���L��&%؃1+��V��m�-A�+�qUb ����s2��U�,e�֪)B�j-YR��(���R�ĦZ�r4QL��RR�QF��[mh�V���TUTF�\q0�c��V�*X��DR�ܥL���"���Ֆ�c-�D�k����,�j�-R�h�Z�(��Z���5����KAƸ�YEb%�k�Lq��i��aJZ�m)j��2�Z�Z��&Q�31fV�\�aU
���nS11-R�JҔ)a�,�Z�[lmB��W&Q.\1*��V��̸Z8�UU-)����6�DkD��V���p(�iH* H����Vg(���r�L׼6*���m��2�v�>B_�S�iw;5�����j��\�('���I�39�>����}�����>������{�#V����>M=�c�b6D
�zV�6D��c������Y�z2�zͿ�8b�v�9�{H�(Z�Ԥy޺���j��]Y�߻�vk�ϓ����iK7�p����?y����/h����K��k���Q��g���I�6t�ۯe���������1��Q�V�{I���b[�Fe"%uCo=�͞3���-Fz;�jK���:�����SN=a�a��j��-^V/O
�F��U'ɾ-��ζ�.��='u�J�ދ�����٪UD�ud4����9v�����%;�{C�f���@��?|��§}6�5O5⎺��1v\b������id'v����S�g�F���x�a�q/*j���M!�I���:�]4��AO�����	�{�ƒ��Rz�+�o<��矵�vn��L�L�e/�|�j�J7'٥3rn��p/����\�e�컼����0j�$�>|���A�$�������l�
�wY=o<�#E���f;�76��v�r�J���Q舏�����6�^t���o�f~���_n�P���-n�
j�+�8�f@\$��6�u]aF%����3��Oc��'�a\�7�M��N���n�n\]f�j5�y*��EnT[Ql��5Fw��}5���.?&9y��Q�8�:��}җ�*��c���Ɩ��v`��cF�i�OU�
�Ի�M�0{k�F�9u�6D��A��J���M
h�1gt��ɛ=Esڧ�aq�7�鹞�]��^ԾΆsi:�ӭ�A#'�f{3�^?U�	�:ӇOy���Y�G�9Gf�Z8r��s��۽��/��D=\���#�?h\HQ�fQ]K����.�3u�{�g��A%��3��}�͟��f�z1}�.��Z�/�+��7�W�ͤ��w�騜�9ήO��TZKw"�m|�eC���;?��<�T���k"6%�>�%]ג�4n��FX���2�s�zea�;��QK��d�K�j�C/
y�e
�'�uӮ�A����l��nN�X�`�է��%�xe,��Z���'��"�hƸ���5�.*c)M�r��b�U]�u�����9J����,��=���cV�OS{P�b�y�p7>+t���6DK2v��;��Ê�1KU\�r�^�����oz
�Q�V9�a��S����N�^T)VOVJd��~�7^�?����n-׷��qb\tj7�7�ū)�P�P!)?�/����.��>��/GX�ұ�K}L�2��:��KYUƕ'�W�|�iP�v���
�v�������p��d�<��5��GتtwS�e���cNbbZ�y!�uy���,>�M���:ᰝ�T'�~�r�9viZ��ISɅ�f[�T��Ȣ&�ˌKv�V�+#��a�{�n5�4Ɗ/{-�W^�J�w�%��y��[�����~so>�n�i��S/>��8m(�J:s�{;bv�F�v�=�^ʥ���S���ܲ���$uh��=N�}�,�"���rh�4SP�RD7�]�wٷ�nw��Y���V%h�Bη<�a[��f��cv_)ͨL��wU-L����	td=
����M�m�V�ܣ(��O��5��Kz�\GK�Q��9���ޮ��h�s��6NsFN��}�W�Y���}�\����K. ��^��:��������$�w"�^��x��o��#E�Q{j��V�j�v�w����{���PL�ݜ���pۉX�y^�����q
��;���k!�&�����4�9N8�Iub�U�r�wRU�7�k�� �ܡz��7S^ߍ�|qW��y�]��m��D͊w3^~�k|�����ou�Sx��̀�yS��Ye&�;�du
��8X�t��'��I����Ѡwe>7�鵾(����궏F��TOA��8�=CD����ŕ|��s���ݑٜ�M>8(J~�P���P5�`^=۫�٬���S/����cǛ�&��Ʃv�#�v>-��,���Mepy:zk	X�u�f�&�5*y����G�����!��rn�{��671�aq;9
;*g�z�k���2�UYy�`f���n*C�em*}EZƮ�����H's9>�<�W �=L������C���z�U�\�	��$�3�C�����\����4���Ұ`��*�Ã)s��ؑ�x4Mɮ�}}�>��f����M�D��\���e��9wF�np��&.����^Qk2}N��}����b)�k�^�3�,+�e�7��4�A�d�_W���s�w�<�>�xKЎdY[�3�����|s�4uΡ��P[ U���	ڴ��������^�WmPו����x.V%|6WS���5����"-xĖ�:�9U�S���#>�v�hF��
ei;旋���W6l��-�5�Ƥ��(�m������Yf�ff����,�Z3���v�U�n��y�%��^^k��G�~�Qٮ�>]�mT�kk�a�J����|_����~��ܪ�>�<�T����,����W&ќ�:�@��7�b����t>>A�7�8����9�gʏS�O0�;��F#7c{�wx���U�\�z;��t:[�Ρ��YSs��ƀ�]�q��R��p�2]x�)����䫵8D2�[�ͬ���y J\ҵx.�6�n+E����|�u�gmis=�2�1���9�T����"V:�w�:�څ�tln�.幅���׸B�.�ΖC���	���.��K�����p��&yj�G���}�#h���4�L�u�ʗܔy��1dy�gw�&��=�Ŏ�?/Tl���q�`�F�LʷO�'��;
#(!��>܆�K�)�*5����)=�m'�fs\u��w�f5��U�a�Ĺd^�p�I?[P�;��J���'�P��z2�4sQ��0��S�}]0�ԋ�~�;�?n�.�����k����X�yǦ�x?j̱~�/e��(�G.ڃ���/���5|D��q^��6]�)�p��ݙp���sqԞJ�x�%fű;djz�Uv0~ga�����E�J����P���GCLu@{����F�v��2��7r�.3h�y��Wq�ɸ�\}����xs[�<�Į�Utss7R��^��w�x�V�o���ĸx-Gx���7xA�W���Lv̿5/l��n�$�Д+zY�<�@`z+�ʵ�Z:�w�CWIo}"F��d֫�9�RW 7��H����sv�֌�o+zJ�`�t���w���TI`���� ������R�N�ꏆ�@��=ԭ��9��w�~�#Kw�v�wa�^t:-��w���4�Gy��w�O��y�2�hG>[U�mf*z�MDw��Ƿ���W�y*�Sίz��I����l~��ʼI��7�ɍ��Ci^{ry��+�U���],��c]7�S���s״zr�{��b;�V�m����lO��Y�Z{-s��\;:��Tgr5�{Ѫ�����b?w�zh8����]��YJ{�`�u	=Z�mQ����Ɯ��^�����x��d�ڷ�B�LeG6���uC��A#�J�]__l��փJ�v`�;Q��`���CU�9Z�Չ�����07pS���OԸ*���"{]L�;���ky+�	t.yw*���ʸ����?�C��K�*���v���`)>�o��;^�z:�Lb�yf'�h�r�1�k��{�m�5zk
mV,��Qe:��7Q��1sa���r��a����*������l��d V,�@X�\|o�^N4�&p�O�S�9�s�<:�Q5b��\��j��Q� �gҺ�H�(w���0�{�Z�U"{�B�L�������t�ƞjpnn��aޯ�����lTB琮�A��]�qZ�͜�C�9�S��u��-d�rݱGu�Q�Ӹ��=��7	�=�s��&�(v�v���w�ϯ:����j5d�_\�0���/��v����tm�#��=缦ݛ"a�m����T^b�{�,m=�!���$$.s[��Zq�n���w���_ǎ��?���ſ.�x_ˌ�l��b�3�5Ku/O}^���;ϻ��}m_B�*���;��Hٓ��˷�tݫi�ާ�]�ug�z��ū=��>0.!T�6=3���[;�q�k/�\#�,��(�z������Q#���^�./2I�d��sn�{^�8�eR�쬂���4�s��5�0zW���̩�۝�˭�Kv\s� ��z'����Q�d�HN5m���J�G�u�uh-yM�=8��n�4����C����X*زn��gD1�L�4F4ۙCe��)��ΗsҚ��ɮ�����f��m�{�=΄�n�tY9K\s��R��ۼ��}n�o1�\y�緔�Uɜ������ĊK��[9ܿDG�K�&����No���of-��Qѕ����j�Ҽ�s��<�1�ɋn*>7�+�[����3������<p*�BR67��& wh��E�;��*��%�{����t֚�����(N���ʸ�%Ʒ1@��g,�K���/��]�Ԯ�6o���m\3z�FQ�jx�x�N�*��y�3�*��r�3�S�b{]�]�p�]е����¸ޕ�q�l��(�8On�s���[��e�W1�˯�j��U�� ��K^��K!�F���J������8��}�[��0%s+w[�Zk/L��ZԴ$�l��]�kg���M���E��k1k��m�T�>�8�������=�xi�o�hF�O_�^1�~��D�M��x�3n'zۿ��E�wF��+Pۇ.�ƺ���F�.��>�ݽ��`�}�}��U�;�V<�6[�����V��O��&tJ���{H�P�]\��ݍӏi�2�G��3W�ܪ�+D�A�ޝ�S�0�͓u����w��c�V�2���aU�����:�븪��ۯA�u�U��c�5��k��.v\��˚��܃w���ǯ]�."��*�To���gF:�K)����}r_VP���NL~�|Ϫe㾳�`�A�o�\���:�^%�*�z��xj
�����
�sc�_{�o�����I�:[�����쏘a���Q���ם�����6��ue�CP�� ��s]J��v���Ewq�MEtÈ�ݨ����`N���Q	1�k@��_tt�
Ն:�GK8��_.h�m��Ȉ6�>j�M'�ͥoBݸz2S��0X�G�k������Ѧ!����Rc^�5��W$�{���!��WVQ4A瘹fr�l�T��G�=�#����j�eN�qmy����y�o��9�1��7k�a�R�W.�0�D�3���y����o �%ٰ]��wOoԫ4�Sݴ��=�"z2q�=z���-`ܻG����y����JR��%�'@�F�Eu╋��jt��b�4��ɣ�&�}�+��2�怣2�*e�wKK�u�U ����Ȉ�GY���+Voukm�]�/�l�ܐd�z*��UǆU������gz���ڸ6��p��)Ȯ�M������t�^�wq>uw�Ӛ*%Vz���5���5ۊ"�e���0n�&JY�J������Q���t�fXU�h��7�KÛ�0M>��`�ײM9�S.+Gg�i��8��N��S��l4;�j)3,'j�-8��ܵ��;�e�C�]X6ä˜�Г���
�%9V��<���ą��� �P_�꼶n���w��yԚ�� �Xq���V-��X��6X��&2� �o3�ۓ��盓��D�-C�����c���b�-�M����2_��c"�TZf�*a�bܶ�b�+��
݌Q��VM8	on���33[mu�������Fजu�m5�t�r�������lԽa���5V�ѵ/[݀.ݛ �!�u-6�P�N�^����qc+
�Оn�)Pet����Ą�2�_f!3,Su8b�
}�m��k��9���釡��qV��Yu���.��Y��Q\�rU�u�+�#gS�%B�5�M�U�j]5ť�c����Zb��`ұrf*u��N7.�]�3���=ٴ�����Q��Ћ��!�*� 0=��.'�z�9aE�΁u\�m��N"gN��W�����ˏV�����a0�YX�wH��u�����k�j��c�P���P��X��o�[��� ��TJ������XY���͗�a5��eu�jaE���';���n��d�"�a[��b3���-S}�rf;������&c���x����o�9[�cH���2�dj�������J�1�և\'9���G��n�9���7����,s�4��-2
��b�s����*�'r�|�t3��������yxAaZ!�q�I�/m��ڬ
�\���1+��+ѵ-we��z���K�M9�'�rI�qS;Q���z1�6�*�
��W�|l �\եr�R�w��Fd��4��7�w�VZ�K��+/m�M�'�`â���.ĘP�;:�e������WG�uqG(:��9|���sP�m�F�C�_!��O��Pm�(ԭ��L]]��\�k`ˎK�.�"�f�m�nS��l�Ż��]k��Pw]ӓ�x$ՌUz� ���)y�=���%���X��;�
�W]ƥua�:�X�"�I����G��h̽� x�܁��ǭw����T����YӦ���˵m-�ܚ�I7M��w�Go7��o>pڽ����V*/
-t��r6։k*+��-�A�h�.e��
�l[q̫�p�90�V�B�m�+X��iV�K�mimJU�#R���e�2��k�j����9��m���liEm�(�mQ�ն��rԩYm���q�E��J[Z( ��Yi`�E���[k[EiL�\�
�h�6��am-+*Pj��TQL��8�&4˃�Ve�AS31�ʮ��ʕU*�V[ZR�h���S.#T�"+�F*��ɋ�-�[V6�"��֪�.e�[Z�#Z#-X���-�0p���eZ6�Ym�(U)V��mY�
�������������K����U�e��"��0b!�D�L��Z���X�T.\ƣR�b����ت�s&LUC��bQUk,TT+�Z5-���PU�T+EF�P�mV��F�S�#V��T��k*�c���HT����S[�U��̓Vu>���624j���!�u۽�#�spw++�F��u����]�)�7�����j�S��w���$����<��O&��-�4�����(<�5�w��������/����K�N��Q�{�O�1���b��qOq���n&�\���׮֜�s�Nc����][j:�s�<E��Ǻ��mV�%rk=�Q��]��{_j�q�Kit��f������[��Mw.���-�%ô:-��v}���Ԭ����[���_3}I��w5~����)KU~߂�s�Qng�Qlp=Gw�d�m��P�&3u�8��u��'�\P��[�m+�<�y��*�(���:b����T'{�m�)����o�J�y�M��!��8�X�~��mH<�1OQ	�~k&����8�nT���xvq��ؾ�3M=2j:|�AƵ{�9 �>u�M8����Ŏ�5^q�����n{�h��f��.�̋�#$�̸:��x3Sf^�R�L�zA�*��܀{�ݺ�82����U��jQ�*��Q��`��hٿ3y��:e�g��} �:���T�0�wj}d*��n�WҁMBnŜ��)V��׹��W���k_�����y"ݎ]w_�:�('�q��\OtMj��i�q���3�1�z�{qZ�x�z�YӽSGwөS�[j�=�F���	���=[Β���U��ތ�wI;r��	L
�Ϻey�y�3�8�z3���w=�tY�>n���\��B�lc��WH񘄻�s�1yt�].�smӵEwl�!�V.ˁ�u�nw�0�_@w����=�]����30�rK���3{-�����nM}��أ{��Iѧ��.�N���'"�����7|�-��mc��VOu��\_wd�2C_:���w�j�̛���S�#[Cg�<���a�2�jv��:���n�_�#[=���p�W������N�o~�����)컨�Q�/=������9Rz�ꋇ�$��w;��kGEk��{Ix��Z�r��JVw�"�o�a�97�m�c�n#p�8�܋�Lden㉑tA@uN�gwr��2���(�W�'������@g_v��[38�v�@�81�ԫl:�9�9_�:�b���X��{��f��'��pK�r�X�7�x�C/6AC�.�$����>Z�f�=��I�E����P�>�6�;�=ǱK_Gfo��M��v�o�[c����m�l��<�K��bk��(�rN��5��r��z�U����9�\�����c���1=�*}�|��k��wQ����r���9%�}�HU	�=/>C��C�C�]����\x��l�_{�]�o�4q���|��B`t���+%M����mv�`oy��sӇ��ĊkC��c��doTI}�AA�[7��nT��o���B�i�������Z���r�<r�B\�`�t�b�����jc{5�)��r�����騃��7�7�����@�K1��j��X�s��wave��u@Z�:��%��T��7)��c�c�E�5�F����9�`�ܬO2do2�3Co:���e�l�W�g���;9P=J;jZ:l��+,�KV�:��d�|��W��)Z�l4�.��ۻz��e+ɩ�� kC;�vRb�`���6�	;�����N[L�V��C3�>�#�v�6��n߆ou��d+��L訃���4��b��V.��3y��@ًđ�H-Ys�ܷ}ޯC��/*{���ו��]�h�_wM�kX<{x��R�]%�'�6���ϼ���Э�/Z7w֕ɧ��K�}n"��c-D��7�ˊ���N����)�5�Q�v1�C�t��]o��+V��gh���X��/k]Y��1[���(�^��Uc���׏���ZUؿG�fm�����3~>z�?�&�u�����]=ʒ��V�{�E�ӽ6�L>!o����nD�4mըޗu��Q�k;7����܌�ok����w4ԙC��Ρ��I�������U���UiZr�봹r�O�U�j����q�tuj�a=�}x�7��L?��D�j��!������#g������L�g�i��1��'Tm�^�u��`e��r�$���y��e���3�m,�1�>dyb�@����y��YJm5GxnSWH%n^s�����!���M�c���g�&N����Wyw��W�*=�RfQ���]D��*��������諭���no���"��"��l.k/Lu���"ҿ�sǌ�ޡ�0�2Ӯy{r��S��ԛX�~�틦V�j�zMMG�����ת3��ʽ�])��ʱDwLv̎n�������e�:��Wq���[ץ��,�+��0���<bRr����"���.������$�n��ߓ�w�w�ۛ���~V�
���4����޻+�Q���/9|zs6�{��Ni�����?|�4�s�#�9�s*�c�}�n-���QoL����b}�V.��Q�Y�Pa]׬\v��a�~]����#[C��������Ϸ\��_.��|R*a����ܹ��{�ސ��o;�D�\�C�Z�_v���y�jV�D�/�ύ��ꏽ�KWx����Ԥps���Gߏ����w��C~}W�~�R<Q�΁�͔5>ǐ59N���4K��<
��9��]y����Y�7�C��>/6��z��\� �竺�}��s��t���ܻt�i���<�El[��k,��ǳ}�s8�Go�����%������pvN�7��w�m#�)^�ENQ�a�5oa�����d���mi�n��D�����{mĒ�Y}X�LF)����˹)����^!��m�P��{xWo����i9�GE������2ߖM�<�se�/��Sݕ-��+xӚ:�l,�1�5ɴq�׳�;��K�Q/�T^�=��i��x�|�P�KƲQ�{�~�]Q�-=g��/��㕈L��ކB�s����=��Ć���LP�#|����}OԽF�Q�YVsðʵ}�������޵�%�)��eW��	Ot���p!]Ne���g��9�.�PV�n�u�cC�2�T�ܻoSy;"7!Ö��=�'9X����⾶N�Ο�y��UMC���RxX.cx�e��˥om�*�SWm����5�����*���C�i_}�xVa�%�*�3��eJQ����]��]��,�us�p���H���#��Gjq�@g}�'��/9��R��I!cT̩W�e�nT]וr�r�L�S
�`htl['�o^�e�M�x�qG].�����4��5d��&;����m��p�܂�6����:��_W�'�e��z�9dz-\OϘ��[y����;�b��]	�w�X���9���>�%|��$.���buU�+�1��M�&�/BϽ�1o��S�=>��;����+]������+�m�էT껭�֠�'���Q�-�5\� ��Ds��M��G������y�,�k��݂z�3�U/R��]YVT�՚�oi�W *�e'������{�{8�[��E���.7R�t�\J�����P8Eɫ�:�Lҷo���m	�^͢����i*w:�=�5u����'�/�[�=���lջ�|:�ؽ6�sIնL�ݑ�nV ����[/��ݘ�}��Rs�J�����J�A��R��O}]�	�"�XVG�ZY���mOzx��b�vbk8�n��W�����ǃ#7]��p��N�1)N��,:�ce���y�('��
<b�n+�����AbF�Goyu��R陙�M_DyT�jv�������@�{غ��.�:پ�#W��2{ud���:X�����j�4c��.�65yw���.�N&D�ԫo�k���M+��c�؇)W�ەvU��^5��c�ل���`'��vi��5���OFW7F���f���]���5�@��#����� .̽)���YZ���s�&3f�/V�={�yP��ٵ9�0bV�F'�a^ॕv��n���ͻ��)Z��K�:���u<5?Y=F�W�j�޺�ʥ}k��{��T��M�79y}Ő��x��ۏ��f��˚�����s1��<c���B�->�����l��@�����"����P^�����;̘�����9j&7�����\8�	����;]l%޴�l����C����V-�y{~k�*#յ]�;��c��O5��z���9�}�רw*K~}�;r�������Q��q�cR�s���
t�,��S%�WnPZ�����:�#k��0m'���-�}hǼ�j���x��O0<g.$C��n*y�zzuf���"�Wx��0���gv�5����Yֹ�X{[�ʹ�_J髱I�CSgr�{"7�IF��H|a��q_m���q��~��Ua�]�.�q�a�!01Ṏi����}�������ڙԧ�0a�6����s��)�띭�<��o�w�w����}ʄ��X��Q�������uD�j���KԺl�yn;��[Q��޷��9�����)��s�wa'dlk�������]4����W�зo�V��Q��o���^���]������m���`j�k��b��ī�[��u�kFuT����o�w�N�JeKP#�
�#ʞ����^ ��jn&�s��gt������y�)!˲�3:.r~�5g,��~��QjJ��������rj��牖j�TΊ��V*���֠#�@uǜ��G��;����4*����<�7���%��oh��]��B��/$|%c�Y������3Sʺ��z�]>�3�5��>��f��;y�:2��u]J��u��V.�}i��z�0�&�k[���'��9�V�5pT��c:��M,�b��͗��e�mE���X��Wi;;��P���_7�õw.g-z���y�Ja��j�k�}�@}�?w�[�Ì��ϭ�!�Bz��5��8���*)��Ux��h8�z�T=��ʬ��81�ai�.7;L5u��_��`�To���_8���1�'�ղ�����j���W>fg�r��+;Q�=�to���S=�a �L����ȥk�/u=��\u�9�ŎFԆ��Oi_Ig�Ӓ; ��������;���7Y�
�n�}�VE�9�Тe�q9Kta���o���o�Yk����D8�N_%��}�ޕD��i*��5��tO=���4U&�X�>�&�^�o�U}�<�I-p��^A3W�R[�5��f�yN5V��uW){rP�$��}k�wh�-���8�9u9�WO�r�1娄��R�-1����(�:��9$�}N��c�`o;��c��R�5���u����-�X5���:T��j��k{Z̾����|�m�l�j�pN��2���<j�5�6�cR�soiO�G�f��m[��mU��-��7�5��9=�Q�m�T��]�p��g���:�T��sy��h��Y��*F)V�<]nsߖՂ|>�e
;ӻ��K\ga�ݛ��7F��2i���z�-=G$�Fk�������Ǣb�ڀ5)^��Pmܢ�:࡝M�ײ����\xh�`�W��VkI	|���ɼK�����J3{�u���:^�������n��l�iY�ԡÚ9l'�	vccR�4>�����x;�me�CH/�l���Y�9�k�
�I�o(���|!X���vg�3���MƉ�r��V�7�"�VR�0z@����,9��ꄬ�_Uؽ��a{��&oh0Z1�/���6z�/~p���S��.ī,�r(:NuH��g{X:+;����Uh�b�+.��ŵ4�CvA9^��7�er�ݼ�&Y	��5%��R��/zT�Q���WWBu�m_gq�jN�l�u7F�YNBi�M�낽O���-0�SğclX�3��%�
�PK����A����RMvK������ �A-�>���t��:=N���&��L�ʽ��a���KҧRk3��mU�6�a��EM�oV�*��!�['q���4�c%�����.�hP*�k��T��}��n�$�C�|���bNZ{�f��J�E�B%�N}2q���*��l��K��U�XA����;)d��vj�Q�V)Aݗ�c,���J��C���k#�u�w����ԉ�e�V�ۼ��w�!,�E3�ݖ�"�ġ*�_&IH������Oorˎ�vf�����+�� ��N�z��G'��=v/�$MΜv-v��Ŷl�lN�V]�U3�Ǽ31�I�>���i? ��[�{-Ҹ�p�[���+'[�I$b�렩�Y�u����|h2�
���ͼ������R�n/�7z���t�g_[Y�W��8���KX�S�o31t� ���{/Fs��MN�U|y1WGV���0�WL�������-�/#R�c��G�v�w+v�;���Vh�D��ee���,�^q����:t���.��׃z
����@�M�k0�ȺH�iT˝�ݞB�y®�q�o�m����y�p��-�B��nx�ծ�y��	��q���rSr�g��Y�40P��.%�b=�ƕ�9��i�Jܮ�}��� �+z���/[}��Os�%m��kR}X^��[��S�2CfV������xmL[|8Qj]�ccw�Խ�k��Ngu5�J�
�2H��vfhh������J�<9��5h�;��0��8۠�%vv,t�O�2�^�li�+��=��6�٦)�}E��AoV���t�˾*A$��os��k��'epS���vd|�����9L�QF2�Y�Q�6,`�)�\1��A��"+1��m�F[*ZTQml��k[�����s*֪�e���T�"���,�ҳQ[eA�TQk1��1��2�b#�e�"�`������%a��
+��TV�q*ɉX,U�jY��#b���f0Z�"WX��D��-X����%a���b�8�b�&5�+F.R�H"�J�UJ�fe�Bɖ�*�V,�nR��1A\�"�2ֶ[,D@�ҕ�%d���TY�`1"��F*T̅q
 (\�(�(�\J�jɖ��$�و(,����DF!KDD�Q��aFE"�"ȱAAd*EY�eT��
LKQ2э��(�m+mUDAV�k��<����k�;�W���]A���S_`��#��r��[&՜���:�sXQ-�L��x�{ �bn���J��&*�r啛�s��Y�w��	�Sq�[ђ�'�W�|�^7{�;d��/i(�1�/��cs��Z۬��Q�r�r����gL3�;KSsz
J3.����@�=�/�usϘ橨�\��0ܙw��ʴ]��eq��k���b�%nN'��n��r���C��;�C�=mR]qz�&�a�����ؕ�y���s_j���U�X}���<�����C��.Q�'��S;B5y<�]�E{�9y��<��])��I�۝�HY`�ݘJ�%�ђ�Ҿ8n��K,��La�&�&&r�n�y�<�ãX؟��oSi��P�d���_+��Cq)]jm幪��O����أ��-^��S���;]Ѿ�&o}�F��lm�T��ǯ�����z]e�M<u�(�Q�r�q!P��>ʜ�h��!S'�x�������V����k�
�{�����Yo����Ƨqu��7;��צg=��E��q\;)��(�d��R����z�F�J���s7���
~�՛>���kQu��s,Ʌ�c�$�Y}�Ǩ&L�4E�E�m>���~��f�1�U~�By�H^�.bɷ�Q��Y�w��ͫZ�>;؟Ͻ��o	�p���ҡ3���u
�^�C���A*j@���y�7�,}�!�&��Ӳ��*�kT-P; �k�Qg�6�V�c�qS�r�{���qk��,ˆ�����6(���E#�-uF�%���c�}먾��~�ҽq��VBt��<�rg6�55-�r���ua�צ\�Ac�\.u���f�����e��㽙:����v� \F*��t����w����}5}�#ʛ��<&�v���>���	���0�);ە9�0bV�F'�on�h�|�L��6󳥶�z7_w��O]���G`;r�xk���g_�7�uK6�[�t�f�W�%�fZ�ZԵ\Y
�}�n ��R����[�.���n��*��Jԡ�x2<���JU�Θ8c�Y�ݻF�L1�i��@�*��I��սY�ӪU���H�:����n�WPu�{zs�{��-�Px��5qb�tz����'����w��crM�1����;{������^V>�IoT��5i�?r��ɜ]��ăV��{�7��]�}�]�E,�嫽a���nڕ�X����a���g-䬸�Amz[ʾ�h'�B�+��}B��,�c&-_K�k�x��^�9㰸_h�­�U?T�U��Όm�ƻ'Xmj��ݻ��r`�;�S-��M�S�l�g���=5�Qp���*/5+���]�m%8��j�ު�֥Z�Kv��Z���R`�n�.ū�/4���s��Q�ي8��koYm��-�|z���7&�l����)T�w n*%?�Z=:�c\�G=���Ɯ��MF��E��y�96�V�zI�$���=��~�ˡ#���"�M'�ͥpf��1{F�+*�(���Ʊ��7p;P�遑�_D�V�5���z��:�������n���s�N��%�q5�+H�l4z�
����E�vë�\��T��=	O�^į�޼�Fب�LL�X��I:����vP����[Xw��}.�hW���FUZ�se(���	G�F�=��S�\���n�W�fq�9�o{�l�ǝڙa���q�相�T�r�\�#�c�c���ep�p&�uZ�9ʭq�f�5kw��OD<�4����Fh7{��Y��z6���e�,��y��O����2��.x�����eU1c�̼�K���imZv��i��+*3�$�4�����i��̇Z7B59���}����[Cy�c�����Rh�=�s�Hr?R��)���z,�����=����^z��ϗ�as��6oh���Μ���݃�Q�]�O�5�]�G�[SW7��s"�Ct�:q� ��Jȏw���ڇUw+[R���Z��!gum9��/Fc����nf/�f�����[��;�Ӎ�sV�����)C���%n�f�E.��3=X���g:��7Q����n�-�O1�T�ROY�w�#�W,�<���8�XB{/4hM��JP��/�AS/��I����Nz�vj�7��:��1��mZ�Т��B�uG�]Ҳ3{���vX�K]��
˚���*�^�WM��p��_Q��u��y�������K�靑Z�Γ� ��<m���.���Ҙgq~~�t�|�8���-����.��/���m~�,�>�~�r�Ô�vT60�3�	5��H�{�P�:Y�O�FF3�{���t(�z\ɚGi
��]�=���z��J���x���g�[9L��%���n��-�9Ǣ�>�p2�8��\c�\'�O���W�c�I۞P#�S[~�;�J<���|��y����:]�N�w�w�8K����;fdS�刖��6�=�Q�6�Ogղ�s�?^���9�o>v_S��r����Tvf;ަ���qo�ܩ����+rj16�U�oÓ�������x��I�g=��;Жq0�4� ��[_E�M<8y{2W]i˼}㸇�=�g6���@�P��S-
"ڍ�=�_�W��gTf�,�b��Ɂ�	��+po�m�o�B�W��W5ѽg��<z����js�f�]m9�u��OgQ�٥����-;���c�=x�J�K���%�C�h���������i7��\Bץq1�Zb��̭�2�sL�����r"�N�����U%ݵ7{z`���Ob�X3.��,�׬�NY�4=��yؚvuE��67-D����iΨ�|2b݅�W�}BW#<����=OC^3,^g3ؗQ������oo{�^>��RX�G�WG'8�N#��'G���r���/n(�Q�r��ą'dL��G��[�5k��R���&���neU��Ƚ�B������wW-� ���弚Ե>/q��g��BEW�y�����M�P�9{ha�T��k17)?����WTa�v�]�O�hq�O��=B`t�A��R0����T;�Lz�s]\�i�_qj��f.c;�m�@ﱘ�{�m��M�$��G(��`���w���ֽ�w/SO�����AzgP�yyV�U�L�]|!(J�f>����n�=�j7�!�	�:f+�9�+�-�G�����I��2�TmD��:t�8>�,������]݋���]��<4#}'/����;%���=��X8���u�pԸ$䦕����z�������`�e�Hk�|�s뼮Ogw�y'�r��kd��Y7�["�hɅtf�z�.��J�Y�]�p�������ЛԺ�9���93\��ϫ{.�e|*{}c��E�P��)n>�U�ö�k
P')���&�X=�rk(�k�6�]v]�r�"�ax�V��=��p�D�C� ��v�eL�)���f���D[f~ŀ�'1�J�]%��3~��Нw����!��1r���f�{I���P�^j�9�����ګ�"� �^B|��{��B�5�H0�r�irϑ��<�6�c���;�2C^��;=/k���%�U��*����-�'���j��ځOo=�¤����>:�?{��#�߽�o��[��VO=���vk�ue���M~PJqe���5W�3u��Bķ%fjx��q��R|�W�mqG{�J*��:N��nm��^]˖ז�JǢXQC=襠a�9e��c���ꢲ�n@ɪ�G���b?]g5���٘1M�ewn&��t�'�2w^�u�p̢i	���FM�h�+��pg4!�f�oS���o\ə�'_Lħs:/=Y�+d�s�.v��e-�m��-��T������P��K}������d�UIC�qT��ȁ�g�WU���c��`�A�;o�Q�����EW�/X�D���
�qD�4O޹���\M���0�V�� �\N{=��^'���+��}��)���hp�W��଩
��)�29�-e,��bG�=�k�������vo\Mϝ�sޔ9�p8;�n�~�IvO�

����ӆ�͊��|�V�Ǵ�t�nUq/��9ӜJ9��z7'Ùr@�_��������ߑ��ܕ��=�Mx�T�;��Tr�ǟ�W�e/L�M�\��b��}��__�ym�#�<�ф��G��Q׶}V�M'��wɏt/u+�,d?M
�yP���/Wf[�=��/.��{ޠ��ˀ*=�R����C���0�=]&�NMDm1�_%f��WDp�~��^S;�0gl7j��N�}��\y��s����x�̡�pf�}y��6���8�&wÓ�"b�,H���5W� ��ͻQ`w<��K.�X��c�Xc��r�;&����	��Wv�n<�Hub)m	Ύ������1p����[mI}�2�Us��˚5ӏoS�i���2goZ��G;��K2�<F��;��6�ט�=%NM�7���l�g�7��˵?"w��~ʶ=��k#���q�J9s,-7�챙釳���dTׯC�g/I�\�og���qC�3v��[�ȸnu%�t��뉸��Δ��K��|_O�K�g	�q-%C�3Ц�����B��3Ө�5k��gI�qw���Y��B���>�O���eD�̰��:2g|n7� �Fj���S������;��J���걄X�?dKӻ�?ϙ�)	��j�������L�8Lr�*�_9XU`� ��ĭ��ț���*u��n�:�=�8{1VB"<3'\���:�x��n��X�-M��;;������W��Zӌ��߯Å�+�b���g�@��t���PI\������#��;o��u��Xc8�{�q�}M���{�D{�C���ɖS�������\{�5�;/�O�x�H���w#e�����~��x�V����}v�/��G�^�%w�{c��5����=�DoeI���*y���c�ա7.��/�����xj�Ú��as )��"�G�����i9�U����W��r��ɱtiЈʏ!6f*�����=l��[��]U�f �R}�[���cz(�hK�2c烤Z��n�}Z%��t%M�FA��t�^%�EÇVq��@�^�ƌWE�O�.�/�CZ�\���0=���ţ�10�r�����8Oˁ(z��^G�!ם����O�yV�q�HC�u]��z6���́ކ���צ�\)l���>7�c")�m��{�ŀ����_���w����Z9�:�!�`��(
���Q7>��c�&zrLփ���j�۽�ݞ��q��ب������H�5U��r��d��2���f�~�޷����:S�q8����!Q��38����x�T�b��t����p�����/I�~��;��3?6�
�Ԃ��8'}�|�;V{#���p=8�}��p}Y;�X�S�@������1�����v�j.�҇g��� g���e�5<��sVT0#����NW��9�k���/���^��V'0�Ixv}UN�W�x� c|�nJ�y�^�Z��͏U������O�u1ݱ�_�0to����(�ŝ�������^L���c�wѧ/�����p�#+���{K��O�WW�0tB�+�X�E���D��#;�Ʀ�ѯ8�F�UV� ���Բ�Z7]cZ��WfH��ͶsRwuN�&'sD:c9Z��|�2 �Z��W��z�-ʽ��:!�b�&�M�$%�ӫ�w�e�N!k�oJ�	�v�B��4N�v��j�3\�7:�q�܋(kd��s��-/%��}�TW)JKK&L#�j���5V�NkĘn�T�o:�W�h��:��Y�\���͘�`�	����Ґ\n·,f�M�(V^c�AS3L�7@������JҘ�t�ǼgP��J�5�܋�%�V������Q�܇{dÚ��0���ݥr�2-�Ήc5Zš��a� |�._W�������.���$=%�:8��Yњ�Sљkw��-S����#�����A�e�X���R�b?"��o����������v�c��U���,[��}�������5��1�"��"	�&jQ)���9��PS����� f�P���s�XB	aߜ����/w��O�aU��ñ�[��-�84�j���Q;����{H�S�B��tVWo3�Q�(g,�sHx�n��X��t@:�Lp=l�IV���t��#���~
�a� ��fp�>��A��7ji�)#�8>�W���w�v�C�u�������1��Y�K�6��S.T�1��M\ZV
��׬�t�h�+x-����IR��#���&��$�ZQ�C�r�ot��Tݭ�@`�t���w	�S����G�ݼW�����`��r�˧Y!��)�m�q�&P�S�C�8�[\U�����Ե�&�J7f��0���7�R�5�]�)�@��A3��B)�f��T0m+tN��_��� ��`��O���g`{ 㬌��ȬW��Φ:n%���u*�&5�n��@o�l��cv���[F�H2��`���5Hh����ں}vt��(�lg��H`�[i*��ް&^�E�kRR���9��b�9:Noj�(^EY���c��6r��M�ʹP�H"B1��	ncGlD�W��4�p�}6�h�t�Ur�t[�/;F�ݮQ�C�.x/i��񨥛�q
-�쌲|X;�"��=�FT�l������PUv�.�#��Y5�A�4)[����;9G��{]p�$X�+���{YV̼�-�����`g
Qx;s�P��ް�VeZG_:��%!B4Xqk&�oN�
�q[�u:=A���/:r�@�})���kB�j.�ο�:��z��fS�;Z��{�o����;���Q�tzB������smƨT꓁�6�V��M�3M0��O:�.CK\�.��9>z�������P��+�����쫭=��P�|Ά�v��H����P:�Ƭ��깿F��J�{�4H��U��<�h�� B�U{]�<������5����A`�"��AE���11��Db�T`�X(,*m��(�Qb�U+�R�Eb2�������T�$�X�*�H����iTbő-��B��[lF�
H�iEPcX��FTR��B��b2,UFVJ��[DU�"�A`V�[QQ�ԩU��Ԫ�HV��R��,X
�A`��,��*,UR5��
��b(�����"2("*2�Q ,��)PUm(�� �%�TD�X��b� ֠��A�JȪE&2�J���-��1	�

��c-�FEf0�Ĩ���Q*dRVVT��R�e�ńX�R"�ٚ�]��yu��㎠��cv�}y��(�x�>a�X�0�7Y/��a.�Mv�����G>X��f�=N�wrk����'�Y7��P�uL^uQf�T­*���x�vߨ�x�\>%�d�{�Ѣ�ԝ�Y˒��y�G�_�:ʞ
�����g���V�~/I����{v����iY��u���cѰ_�A���JG�����_/Z����O3�mߞ8�N��W3[k��x����G����� �h�n�ңz��Z>��j:��w�����X`m�7�7���^�>��H�0z�d(�n� ^-�}^�G2��?���\ô��e%��>���_�v ܠU�?[ ;�����t��n"`����Dc��)L�&��n�ۮ;��^�>ґ�9�5�j=�*��Ǒ�u��~��y>�$��s>���p��/ڣ����V��RGz.}�Ek��,e%f��u鹌��)q&=,��vR���J�*��O�᜖�D�>��뛨����2X���:�m1䦃�\_�ʁ��F���/�P�wQ�-o'C=�*DWp���ǵ�4��E�?�~��3Z>�����'F�?Ƒ���с�+���̨��m�mE�s!D����n's2��5ʭ��ƕ��+�%t�à�d��`^)��ސ�ȅ�:k��W%��t��������=+sy�*���,wm��:�gp��R�Y9���e�FwZ!.v��^繂mW��٩�m�����_���X1|7��|��e=�ە� z�`\x�n=�*5�\���V�Y'N���t�{[p�>:���/�b��\��3��(S̱���_���Gw��+ت'�}�<U����꯽)[�8�Փ�b��䞊�M3돲gT�����7�T�ˁ��"Sg��Y�_�T>�ˬ��\��LY��n���U{��}.p]R�x�Y8�FL�WJ�-��}�z��m����K�9.Q���.ı�_���0�	GQ����������ۭ����O�����D��k���ʟW�<�Er;�;���\�C��Np�!�u4O޹�bi�D��W�܈چ��m%��o�q�fk�yW�6��~�U&s}�v}�#C�z�ɖT ��x�AR��-�*L���ԏoj�{Eo��	��9
���H��Ge{�tT{/ף>�˓��}
��I�=>��mw�K�㒑̀x-9��*�Wr���<o�EC��.��r-̹ {2���Ն<���Y�1��5 _OLV)�*����o���3gw(������9������>�0@Z�8D�t;�jG��k[ڀ�q��zk��ٺ�.���|�%w����/�A���G-�z�+o5�
:��Ҩ$'p��2�q7=T�Ė�pߢbc΢�1J{�FJӹ �5ܽlx�]LǸ��}�]h9��T(�Fv�/�fVw�Uנ��t�����v��\ex����h�>�%�JjK���u�Y�Oz��Fn��-�3�ѵ8��ˀ+�?
@�ϸ���C���0�=]&��>���ѵmǙ˅�d���#ˏ�n*��ې'��ǡ:ɲ.!d�8J��L�d�f׸���U׀ a�ܽ�7K�dϾ��P�e�d5U>#�0p�?e�42f���J9s,-'K��_�g6��V�-��Q'���ZofX�L��|�,�d{"<�Q9J}�߱\M�G#�wH�pz�L��ovO����J�2�2kJ��X�7���`r�p9�g!:�7�\I�c������� fGl�fny}^�1�a�I����+������޹]�����Kd����=��Pbw��佫�_�kۜ9l�0�0JF�K�zf��:�,�oLO���+:�����kR�*EϚsi��3����}~���Yhh�~�H- ��K	M�5	���q<�^�?J�7ws�ΘX�U��{b�b�/x�x�T6��t�paثs���{
�a�<e�^�5��z��nlܶ5u<�1���e?V�\�nq�oL�=�U��P��ƥr�O^򖦫�ţ�e��bCMw{�.�ݰ�z9�J)$�c5��Ż�����dBR��w�g�"�lx\K�l^|��=9U�;�qE�^�Q�B��̩���O���ѓ���M����=���9����K�}~��+jYx���^U�3�麚���kW�[誑?�"|X�8��aT[W�o��m�k��}Ǵײ����Y�^�e��%k������D^j�t�V.W�fς�jЛ�]�G�����w���Sg�FǢ��v=��+��̉)M�����L/W�H��}^ӄ��� ���#ᮃ@�O�����ͽV<����>��W�<���7n4S����KG�&@|j/�bi�m�v�3�VM��U�x7|�V�bB���^6_�r3`����%�>�f�q�D+ŪC���[^;��ϔq�I���q����{Z�͛���q�Tz�ʒ|ϊ���^�{�zB�7��IO�g�օq��Οi2v#K�Kwv�U>���N���Q�gjp��x4vS�uv��_�����x���x{6p~�����gr���N����Π���-�ǹ���
�ý/��N�o�I�K�6��H�c���|J��A�*�mv�P�����ث����u�h�C�۰���m���UL��[-_?��]p���ב�뷍>���	0�F��O�\����P���^�>�ݳ�<��=%��f�FW��f�i�r��m�K���5�~_���I��[�n~ˮ~d	�돧��k�Z.!`��r^,��xk+j�z���5�}��do��z���:��G�u�n�W�hp��B�$��,a鐇��7�7�Y"���$��wky�˟}�X,�s���~�q�%OŮ����?k��%FH�e��\��	ǜ���x���U��ɟ)�ɞ񸍥ViT�����#���7�\ns�,�w�]�{�Y$���:3�x
g�.@�\U &*{�U��IC�����VJ�3�Њ¡�������y���{����d�z&�
��z��.�A���H#����^�F�
�߯����;c�_m�~O�5٘�[z�<�N���Dm}�~��=5@!��{�R�W�a�Z>͘j��"�#?M�Y�Հհ�-V����8�3�9H��<=�]���Q�yMF��_W��=y��fl�d۹����sG��	��?%q7���ep+�@�=�r*�S�/�,.7��c��2��=jm���F&.ov��YMPC���{��*{���^��5`\������Y��P���]�#*�[C�=Q�N��K*9����E5���)0�fr�MyG����@m
0��.��v�Q�^���f��*qu����T�b��m�T�Q��������wN|O��ܼj=~�����}%���w�@L;�I��qޑ{����B��{��9�c�ꈹZdT}������*3b�M�\{·��:��צ=7��E�B_�mv��'۲�����뛨j�+t������3��Ǒ�X֨��&��.g+��]E���^��'v	�&�t�=��~Zد���24}wc�s�;�����N�y����������!�����bE�s�Z.9��2�۝�xo��T;�6�N��ZLǬT�6�Γ�*}��@
�.׀1���\j5�\����Y:sc�3��vX�"��i��Go���8����g��o�>\�s��]��7�G�_�+ت'�}�<U�7����M��yC�51x)Nw�O����5�ד:�5����z��m>�g��=ơ����`���y����;�u�����8K�|lت`Y�62gY�ɞ
���Y��l����^G�����*N�ף>���;�Hrs��N�܏���0�	G��7T��ȁC���1���M>,(��|���v�t�q����wU�>w�9����R��x�����uPv<��v��f��1r������FhS��� \�J�X�G��]�0�$�	NZ|{/&���;�L֐3.�;��%��r����x��p�z�W��6�9��g�8ٝ��5�#�'H^F�;-vO�[������<�G��އ!��<x�1��"o
�z�{�c&�_��嫻�H��q��H�z'ù��ޯS�TYw ���ߨ�Sx1�,.�[�����>���F�y����K��}��_��:*=����UzKρ��#�9TNNK���]�^k��)���~9���F���Ȝt��n<W����.�ۗ#=�G����4n���[������s��=�ta��;�\�h{>�R�La�R���_W�o<c�'��\vsΟ=����MGe9(��O���n���x��j��ƹ����UrX��o%@����e��m�GOP����� �?
`�ϸ驇��V�q���Q���E{�dL�/77%{q����5��̳�{΀��5C���+�I�2�h4����Ӡ���]m.��{�����[&j6��)�׆�N�CS���Z�8k��r�XZd��LOp1�F���+�����o��Z����zM����=�N�Ĥ}ƾ�g\O�Q¢"ez(��g
}����>�[9������d��w<���k�KvV�'��wnE�A!b�
�2;د��(C*�*|r'��J�tFu9w��;��Tƍ��{>�j��=՛ӖF�V���
/GK�*J��'����Y��̱�*�q�V�&��*t�L�g�˹�����9>����&xm��!�5��X�;�o�綘��@��kJ����k�^m����ˋ�^����񋇂wM��)�/rkK3�:�������)���G fs!�+�}�{�n�uǞ��w������,�ڇ�_b�b�gY���[q��5p]��|��|�?C<���/W�틟9��w��(+��=5Xjnj޸w�ft�~�>̽57���s~|V��Gν�8����Ke-�_�/��
v�=�9U�;��]����Prξ�n'����g�}4�?+�g��ٸ}�-����ĿW�W2��
a{)�4}xENtc����,�k�U"bK�o�,y���Qm_	O�ٍ�t�>�t�����z�aC}Wb�F`ڴ)u��-��RXB�wmM�6���òx�=|jd�;<=3K��,�?���~ۯ�n_�$k�6�4\9f�_��*���^��LLS���9�X�Ke���>�+g�w{8���G��+�@w�܉n�n�h�̀����T���x�#��l*D�F����.��E��\��ƿ89�x�>R�F�{�5Kn��\�7����|`���x��+W8���,�j�d�=�k��6B��Vl˾G�]mJ��l&dv\ݚ�N���
����o�>�񿏕�d9� +~���� 뉌7����p�l��^���":fu��>"����Q��]�/M%f��5�7�:�㪨���$���W�����n�>���>��7>fօy;�5,i��/ƾK2�UU�Rt�:����f55�݉�]~�?������ӳ�~�����Zo\�w)��r�dxg�s�T^��\*�'.յ�]㦶愥�pǻ�{IGL;�qb�6kN�{r�������~���Y��ܕ���Ѯ���cF�+p�Ix|�a���ڇg��������g������K��K����[%i�wz��R;��B�2J:Kzd!��f��1�5�y�����������wq��^�������㸕�w��w�(��%C��h�1;�{M�bk��$�U0&Ҹ��d�s�<�����Y�~����ߧ�n"V+�x7�C���%�TW�ۺ��Y��H���2��yg�G��q�z��#>gFo�Wq���~���z1��v�Z��Y+���-���`�n��#P�Q���ļ��AMU����"�s�Q@\+��nVբ����y�92�k�ش*c���$76�v��+��.U��L:�mG'm�E ᰲ��[��
�-���>|�-��a��:w���.5�q�,�c�th�����$�x��8�e���hH���ڡ&�8����K2���,�p���y/ޯ\!����� ���R�zU�����i��f�zc�%{3�wzyf�	�R+��@��u����[���� y�� 6i)�eV:�K����K�7��f9�	��Ҹ�T�z�B���`ߕNe��������S^�;3��{ױ�6���KӸ
gt�//�s��6Ϥ�Y@+~��&�Oв�uǑ͜���֪�Rp��.;q7Lv9!���"�\�f�cuP�|��s���:he>�#ψ�^�Ζ���w���&�K'�nO�����������Z�A��i�RUrX�N}P�Px������j�Ӟ�v�	���r�Q�{�\v�v�z�L<����O>�o������w����7� �w�V �3>!��P��0PX��rt���gnv���T7Q���a�ױL�Zo���T�3�+Ǧ�m�)nz����G�UN;ڐ����N�p�K����}�oM���?��Ŷ*駔�br�[�ґ.��+��kz�Q�Ť��m_�9zw�%�1��l��ü7R�Q�r�+.�@����ǭ��.V�M��#�=e^d�x�{�@�5�����Պ���m��cႎ����ga������:)K��H��:�8𯺙&M�����Ʒ��x�z���+�:�V,��:cS7(���O@���'.�T8�<4�ޝ�.�%H��o4�
���6����dH�d�x�e;z9=9��$wwu�t��[h[�f�u����Q)	��*Տ9EZ �]�v���P�].��j�c��5˜r�۴��Un��.�Xq�E=�9O���7�Q�5��#��C%�<iv�]'u ��I�n<׭U��ƈږ]W7Gl�4T�jrE����J���;6�+�L��s��]�5'T����p��Zڶ�,���)|1v��3��)ٻV�9�,r���k�v-��6qJ)�b��8���&	��`��qV�C��u!�=�z>Fr�i>8z70b+�lE��,o���q��O<��f.�u��/���s��nmmv�����������詼��샞J�wIFq�]B�&rT����2�X�	�a��t��"�rj�1��'�Q$�nsg�h�u�����>IwT���,�νg�%�r�z:S8[�k˧b�*�K��t�R��<��.`��[[D�Ǻy���#*MJ�Ӡ��%���ۮ�?eN*����H:t�rjY:��}��X�'�rYT9������腠wB�R�)]ܠ��+=��"��XY:v;��Ip2��$�����Xi<��p-���|V�� V���j��܈(/�]�VC|��k,���[g��s)�1�f�������L�9���y��4k/��骨�Jv��*b�!�\���΋��,T3'����0(Tܢ������+;@�`ՑVF���y.��`ݡY�����Z����lnYRL����x��J���M�X��ys�4臘haޚ��x�dZ!�d�b��(=
��Z \�����X�I�d���N�u��� r���Yn�u�U$7;��E�8%@k�N`1�E��]��{��Ѭ��,�ٸ0J�<�e1�R�0�sj.X��^`b��6�-��\-"7�:�'�^��D���$�فC[s�q����k���\������_0uJ�\���b��m��yBj��P���MՠJ���Y��-���#���F�OA����]�Z�3L�{�{z�"9�9����n"9����]�q��j����y2�̝&8P��,�d�J���(���S+F��������n��t�|�չqm�[���}k����Zλ�;UH��dPQVD@PSv�>5�$P&5YiaYR"�$�,����Jŋ`�*�c%��VH�Ĭ+++DU�PDĕ��h��a���&&$PDb�em�T�ńX�Ȱ�*DeHc��"�
* �0U@Uh

�!X
�If"ˍDdU�V��
E�Q����$AI��"G-b"�V(�"���-aX��UEE��Tq��Z�m++%�,�j�Q"[*ZB�EUW*I�ADY��a���b�R�R��
�*��X��1cZE%f3�-k �ŕ*c,IXE��Z�31�eLJ��������T�\�J� Y�$U ��"���Z����}��g�1���6�]�9O.b�播*���������,�X�F誜ln�\���#Q;C�m�*G<����q<�.�U�To�|�tzx�>��d�ϫ�K��7�j���S���1��Ϻ�k���]���}�2��zpqL*�ɭ/	�Lc#��������n�g���9|.��u�~�Y� �%)`�K�w��,�a�{��~V������ig��Dv�sa^�l��,��;�3ƹ�ԗs�=瞹�~����*>1���>eM�T���D�쪎hVlkś#�ڼ�G���GJW�#\J����7���c�w��:�8���P��7H�c�=$�S�}�Ok=�V���V{����6n7�,.�Q;�����,�nh����r��ў>�qç���pЉ�}ΐ7<��چ�E��$�RG�#����	�Q�t.=�Iw�4���Q񛬷�K<"  ��G�*|�`,-9�/Ƣ�W}Mg�t��Q~'��y�w#g��Nb��z���H����g���L/U�&b������V����r���R�LV��G���ٗW:qyN��oL�jpq�nD��ID�����}s�c���7�k���>��gǁ�o��љEP��B{�v����|b\<����ܺO����*ވrP�)�JnF^�E�H5v�)���*�+��%M��f���E�z@��ط88z�'0[�-�C�"N����Ҡ�R��"θpM�s.�h�3��(a�O��ٹ��u���꓈T�=��Q�2���0+�\�	���`z�U�~�'�qD�C�����iZ��6�Ǔ�"�4�]���QU�V��vi�������@y32<�$/1'�\���^>�<e~t�����^Q���{N��Ͼڇ�P�e�53>!G������{6s�-���ّ�wx�Ɨ{�cl�螔2�ևq���zX�L�NK�_v�\{�d�):k}�q3����xE�M@��cX�)�>��}��}(i�b���d�V��#}7�,�� S��:�w3Cި��%�=�]���ŝq7��_���dU1�gK�;�z�w��o���H�yi�v���ؖ�{��o:|{nt*~����(�X)�𞺨~.���ig���/��*D,�Z����o�s��F�߸�{�^G���e��o�~�O�ɣἥ'^74���6:�f�<g9(��C�N��j�3p���Ωw�;������.R��9E���	Qys���
��2�k=��2���|�V��U�x������\{!Sg7��9����^����j�\H��U�b�I�9��n���nTWX�z����"��Ew�w:���0�9Jg���<�뮶v��S �AyR=ut�ț�L^�-WC��s���*�dإYE�2R,өu��)���O4�5Qy��+���U�zQ� $}���qU"J���ޖ<��a�j�;��>��DG�&���kI37�Uz�xᮭ�^�Ҥ�0a*�J�A+�aϋ��>
��B]�8a�q�@������Xxyv�.s�t���ۙK���@-��&��O��p����rv���EL��I�zF��Z��:�7�(p�7�<�m���@�R�ۙ�	��a���*�s7���qH�d	���/���_�:�>sX W�����QD�χo8��q��v(�����}�V�d֗��o��P���m/ea���@o�3��.������C5�jG���oqگI6�xs7r¿�kC��w�ke�35X�Ww���Ƿ�t�dmM�����6|��g%^������&^������x~��wO�2tV��u��`o+�G����{e
Η}>w��Ib�@�K��/�4%צ�+jz�k�ǵ�~[�Zcm���S��\��/���y�@�eg�V���\;��:5�
��$;>���mb�o{�5��^�M�E���w���y���B �u�k�����\�oQ?�r��*M4��%ׇ�w�.<��������L���|�o��J=�����ƍ�]I(�\L�x�5J����ݬ��۝]}��o{�wO�6J?�����}v#s��2jNq]��
����8{6PY�Pۈ�cI���wd����@�s�(��.��N��aa3q���y���Ǻ}�b/���{]��-����Nƹ������v�s�x�\U /�Q팙Nc	�{�VF��||=�_����lT#謸}��W�%��o��V<U���N�늦�O"+�	�����h{!�:$�|g�ޘ
cӊw �J�}�w��o�y�!�Y��K�G�WR&	H�7�^�m0��K}!��a^�t^�����=��V�C��[�Oi�~�\xa[�xnj ��R�z�� n��Y[�U��~�*����ZFE��$s����/�D`ｖ>5<栐=
�u,�n=Ε����z��3�a���D���x��W�?g =��Z*�S�=W�乣�陝�cs���2Ϣ`���1J{N��wO��.���gǋ�����VP	�wz�LM?F�G'3Wg�s�{�>6f���:��C��V��wǲc*!+2��_�TnQz�������]:��cu)��Xtz��b��/�����^��]����s4��3>v~u����n��O3�go)���\��}J�	�/�*�#O{n��y��W>NLԏ,�3���aĬ�<����Oy���f���4�����_���V����g"b�'9�'.ݶ��x�?�g?����9RMG����>��z���j�K���{�s��F���~���}�L��<��TU�Dc�^��r�� ���>ǵߍ-lW�{�޸�M�����bc��[�vt��߃S3�����3�ƻ5=�s=����y#b�0���˝ld�Q�Հ~��~�`�<&Ϯ�k�׀d:�['�k{�E�z+E��:v^8׽�ٜ��r�p�>�R�^V�,>U=�i��s�˽^%G�u��◵\L�/<�K��v+����>��ܒ;I�{j������k�\�"ާl{֙H�����=G�����Uʣ���v+�g*(ՔJF�Ӏ��0&.{ŋ���p��i]��ba�_	��=�=֣��=�^G��^�q/��{�g�F��5'ȩ��`O�<�g�N|rz=� 偕���-�q7�z�P�O?^����u1��HM
�B�!�����0���u�>�٨Y����6O��+va��ߺ��ϩ���ǲ#�Dh~�W��,��Cr,%�F=�f6ck:�M�",΋+K���č�hY�HI����q���
ʣ`3��Ը���[���6;2����j��$�yE�ý]!駧R��]��񙵓[�32X��Nv��|�4�NP�ԣ#���ղ����%�U��ʢ��%� wL�=�Τ�h�sj5m+���~��Ǧug�,w���ǜ8>s]csu�nM��q8{�ϑ���4�m+���}~�Ϗ�8�t����[�{�>�O]�x����G��S�蘘^��D�9��a΀X���CܒӾ����K�ncޟm�3���ǝ�w>�Đ��u�+���5[F�χvs��v�Ⱥ�F|�2��{F�r�K�׊��C�.M�����x^���W�Zخ�k���6�,>�:�~��|]gS9P�)����@yds����yD;'M����=��U��O�v2*d��<�����������}��}��;���j�|G�`�~��m�Ñ����I�K���v�S�(��gB�q��\c�ó��ic�3q�����^�g���ϥ`t8����[˷�>{�tߊ'���Pۉ�c/�Ү2|+M둾����\����|C�kb�Pκt[�w�����d֪'���V��/�ESQ5��'|z5������DLHSc�@���"���Q�J������stu�Q�5Q�k7�w�L�Ƽ�7�~R3>ͭ7�w:˷:g0���k��D�u9���s_fu*=s0�Ӟ�F�+C�����X���#��%�@�ӂ��v�kf(p�Q���*��9��߹��->2������hw{jQ��R7^��T?�WLUF�^Y���n���&;�4���o����:����n����i�(�Ia)�8G#ʻ̽������@z"�\;�h�ڨ^7
�\<����s�-��߰��c�OQg��s�>$_S�������=7������ygU��E{������o�����O�6���V�<�;z�����E@�0��d�T�&�,y���aU�|%?SfSb��U����[|�;ˠ�l�T�/)�>��Q`@l�ӥD��r�s6|��#�8�h���Z:��}T�c#�Qs{d�V�.$W���,��10�_]"bb�W�������j�_����%��=�§�H�dO�_�e V?^���q#m׍�E��2�]�9.����3��t�ߜQ�}{�To�����1�5�%�~n��� z�R *�{,
��,�y����(�y>��Z�����6��#���;}��x<:���5�7�<�C�����z��>�70r���hj�"��P-��gs���_g����Z�ʉ���WOI��wSn�I=��*s)Н;���v,��D������i�x���K��`�����7��X%��v8ݕ���B�N����5�����z�Z���պ�Wa�{,�h,-=7>
�6�;����e�35��RY��U^�w�<©xS�������㽕Q>��8k���/ND�3�g��d�_�:+M����07n1�Zu��M_,^����p���� cTt�hN|����'���Ó�2�ŋ�6kM�y�����ہ��=^K�	q�@yuk [��M�j�Jj����kE�,�nK��P�ܼ�;�~�^_�=��I�o�=^�q��5�;�q��6�ut�sÒ��2;�i�Q�	ƙ�ԝ�"}b��9c�X�S�:*����lxs.#����~�iyO�Wl]F�Pߵ燳<�iЀ=�c�^r�m`^�v��0ze��}�q�)�^L�;*h,
^��>�H�r#��zx*c9S�uz��'q\nD/u�V�
=�z�<����F�*Pw�z��=��+��:��$��K�[�i#�%za�(�(*O�H�H�R<O��y�~��=7'8��T�|��so��~�3�J���#:!����9+ơ�!��t7U*1�|j�\�{܉Wv�"~ʅ��Ϧ����n�/;�J#�h�Bή��9v�e]W�N�z�r��Dmbu�W:=�se����Ѽ�gheu�h9�
7~V�A�TZ2�K�b�K��o���W�p��{|�ٿ� ӷە�r�`���P��Vo(9?��_��"\y�RG�ïRG=����н�����v�2��_cÝ�Tk=Z�����[��}g~�|3/�Ǘz�{�}~�Ϗ���נ�ʑu/��ಫ�~��|�׶H������DM9�;� �ӑ�=��Q��yUx��-�I��X&b�'iI�{�^[ʼ�����.J Ǵ⛦:��C���EF�������9���z��6�Wq����va���<�#�8=p�T�Q�>%iȓ�z��������Q�t��ޏW�F��sݤB�wޑ~�ʹ:.9+�ddy�=5�C�\�#=��J]�	�V�w�0<�����^�;�|�|P3� ��~������6��.Ďxg�9<p��.9 �xO{����X|�T+ͪ�q��=7��q���<e����̄����'�9ߩ����?���y����M-Z�ꢷ^�g׉ �3y�%a�s~N�����F%��N^'��ӕ�����m�Y$n��s`�\?e��ҭ,��g��)�����O���_���ڨ��0�H`,�1n�p�_/l�8�M�#]��]�V�i=��hi�#��n�5�S�k���
r{C'��J��7ǁ*�$R�v7�e����:&��E�O��S�f0���_�S־񋟱>�˽+�Zu��wڔ]��ݜ�]8��oS*��x����#*9ůӆ���������w�u�	Hܹ�u/u�>��_ZZ;��ն%*oG����b��6x{����{���q��g�F��5|���*�SȀ�=)�Nge��d疕�;s^��GK����D�=��������:�g�%ѯ��;��POn�x��Y�_ny��$z���7[>�چ�n?,�o�����C�a�'�z�ldڔ}ro��g��7�_b�:��N�M�FD�N�������F�uD���>���#�����|/�ɧV��dZ�gWr�]�t�\ >0Xu�UB���9����}��m�Q=
��Y�|��Z-m�uG뜽��ؿ�d��T~�"b�U9 _�0��t�������>��`1w�z�\��{�A��Y�Mw�>�=����V�0�)zg=S��TN����M�h���>���LM5[F�c�_K��󛽜]U���].�o�Cn5ՒſMxڗ�Ҽp/���K�i툛�]ԧ�_�T��em�y�zt�c����u��Vi��g��R���x[�4Ey�<s~�4_�U��RAO�Uc��9h$�����s���up�s�7��p��M��YT�ڭvp�$Y���|އӻ~��v�Gk`�;:ܢ�Ʉ� ^�Ԙ�H�c)>\z��:�1��eۼ�V���$Kg�?L;KvS�öTb�+�᫯������h4^�fhut��͚O�E�T�hs{#s^�'�5a>���R�5Fo:&�c�a!J����yˢk_-ٻ�tGu�5�T!�/oe�1fw��	J�]C!�f�uz���+&���S|���K���b}�n�ˎVg5��!�O`'���PȖ�S�-�voR��9M8�Ge�J�|E�J�m���\hrF�y.H�γ��!�*�������er�o1�s  S_E��Y"��o���Hi�����I���rQ�䬜���[��8��c���U[W��p�;�J��Н��p�v[�s�0vZ̥�]@b�T�6�շ֦op����Sat2��1��U/UA\����t���+e����yl�	Y=��[y�;-��׶�t�c�e<V
0k{v��<�!W���I˯�ghِ���n��Wڸ5#.�� �B(OGR��퇛�J��IMy����V�WՋ���pU���;X�C�n��w�h܅�b�i
X\ts}¹�c�����PO9 +��[ȫ4n�۫���>�K���yb6���64�ɼ+g}�^��{�W��`�/S��B�N���m��{�Z�[K��2q���`�׼�C|��,�2�ȆCc�ꊃʹ�ǎcwy�9-�����w���ruJ7YB@8r�+��:�h���sz�S�����멽� &܁�+}�h��LCv����5Qc,�np�{�f3Yd���S�&��9�:�v��W5�n�bO���^��]��ً5�*�c`%j�fU����A��T���iRUK�P��m�\�Ż�Q�?#��w_a���+�Za\�~�AtB�̼��k��t:����jJn��st���;�j����#c3��K�
^�vv�(��"���o�'�5<�[���B�4��;Ӱ��[x� ڛ�5�S�%�Y�X�Œ�ۓ�R;��@��!Z�=����ӹ��*��ɝ�v%R��+�7M�3{�{�Tf��.�幑�n�T���pؼ��.��o�-$�g6���WN8��ϴ�w(d=h[�LI� �i)���l��/��ΰ�T�/���~��M��m!l�[�^[��>���J(�4tm�ԓ�%n��5���#�]�'l}ϱ�-v!W��������$*j��H��a���+hhW��tͅJ��gCQ����RN�<n��M���+�a�F�H�D6���Awqh]b���g8�=�\J�(l���0�[lq��y��v`�AE;��s���Ͷ7I��v���n���,�*���������m�(�(r�UaZ�T�1.P�R-HQ�SQ�Ud�Vڵ���UU��ij��Ĩ
�1R@���E�J�"�9Ak���
�H*�̰��IP���TUR,QQ�)��I*(�+*
E+**Ŋ0�LI�ER
��Q�(�R(�b�D`�5!P�*ȡ��,F
T�,@�"5���h9IQE�Qm �8�22���R�IR
���E�V,J�L`Un\X���1DUƵ�eAdZ��s%E1�U�m$��Ȫ,���e�
*��$1��CV.%d������
�D*.5Qa���U���@W�G�FEs0w^���H�^F���S�S0)����Y�p�8_l�c���	��n�D�c�e��!�j}�ge�Ϻ~���T0ߠ4��z�i�/����~5�ǻ��T��ٌF���dJ��;�Kw���s��}�����[��,{I��{����+����e���q����D���J.B���ڋ�}��:}ٷ�Qè��踟Jr�֏�5�+?^�j����z�Q����[�W��.U��>�z�<���ʝ0�`��q%��Ȫc+����=0��!����޴� ��n���^$=r��uî����\�`�z$�'�*���2�9��S�՚���<�|��gUA��ңq����u�{b߬��~�c�G����7ގ>qQ]�\.��=o9(X�J�0����ǯ���6���}p�i��Ke-�_�/���{Z�v����U�u�������<�v�b)��W<���h.7��x�M���;}���iumo�T�;|�\}>�����i����[R&
���zX�;�,*�j�J�t��y����ϧ���]���Ӭ��'O��C�E��� CnT��%x�9�������LU�Z dN�T�Õч&TfPβ�]�աIӺ��c�5�;��US�U�'��M5������9Kz�̧��ra�pnɅ乎��T`��7ێl9X�K���{�e�/�nTʅԊ�
ۜ�Ռ��F���v��1���Yw��*I7������J'�C=�|&�+^,o��E�ǶHn���0)�5
�h��L/U�&=�����+�:����^�9����#��W�A�R?V ׷r$[���Z={ޮ���ή���`,>�&&��h��S=�a�K�|=�*�>t��6 T��~�z� ������nY�}<;aPxl��ds�x��>�����_�к�k�6n=�@yS���<�+��ӭo)q��9RM{������ܰ�6�;�ͯ	��cL�F�<��à�¹��=�R�u<K�;1{�t�[w�gp�����$��q��� ��)c�a�,e�����Ma5]�׀y,YdG����Q�X�M�{s�9��zKGnv���{�Ŷ�Rxwu��Y���
�&}ސ5�Gm�)mg�	�'�j�u��-	��5��X't�Ix|����*ɷ$��	���~�Fѹɍ�g������Ѝ�:퓐�y�u��{/��4���s^ɸ����5�[��w�8h�T��
�]ÿ�g}7��K��ߣ���}��=�/��]{��0g�f��c�iKl���U��`�3/iN1��伺�%�0�xcj���+cxCՋ]Y�z�8�}���f�ٍ|N�6Q����_V��trJ��5Ǫ;cn�(����bb!k#��SA��E�����a+��)ӎ;}o�>="[���,� ��������ɞf�iU���w�3�gQw�����%v������KD�1{��,���%�z@�L�2"*yg�G������t�*�&iGyR<��|��tf�U�_����y�b;E��� r� ��&�=`�0è��<u��+}޴����{Θ�O�<�$b�_�Ϗ3Q�Z4K�}?�̺�7��=���'�FS�|O2�6���v��p�ԑ�{���dh��[��W���V�U��WR�����r��� y��4���%���&�$�Ȝ�ҿQ�<
O�z }�0R����^jF�+�w> {�Ċ���7�U�"i�i���r	xk��G��W��P�	�e�3��1�|���m������@k���7��>;M�Fz�vV��|6zs̢r�mT��ݽOWEyy[�����Bznc��9tM��^��*�n������'ä���<=��ݙ��R��>���ԟ�����r'g����ʐG��HZp������b�R�rg�.��p�;ݠ��=de�t���Қc��!���D��z(=�]Y�c��0]�S��X�{�mk����k�+&n�X)�1f\��5�+s����;j�F�t������
C�-��jV�n��k��5�Y�B��M>�O5^ O+��d5U>"ו����]���������=�y������=\�/n;0��مy3��_�M�� R�vg��\:�FD�v�ޘ��5냓��m+��;'�ze����ˌ��X|�p03��yׇb�x��Nq}9l:�&?�G��.�TC�-�g�(%W,;���(z��o&w��'=&E�Q�_�e�mc �Y�{]��ѻM��L�w�yu�o�8JF��8L�2�X�ɝfU{^S>��-��Cg7UΫw�3�[v}�4�xl{��;�~�x���\m�{�<al�ҥ}T�sO)�e��u������z�2�9_��8�V��%q����/-1N�q��:����/?d�Z?���5���MC[�d�a^/sj5���}M��ފ�Kz�h�~�_������d
�s6�=�����@#�h�zn����p7�h�va���q7�i�zB<ϮA��tN\ ��?,�A��_�]�%���_,:���g���Ni�Q�q���:���Ҥ�B�J+�j(�ἰ����'���{��Ւ��즲�K2�.��G)-3yPݴ�"^'b�Mt�Ho@�/���*��LO;:�w:L�;�A{OW\\F��V���nö����6v�%��n��S���G[���qI�.�.l3����g8�r<�S�ٷZ*�S���똘^��D���ta��;���Ճ�1ΟguH�Þ�Ls�L�M���"k��(����ۛ�}q��az0�O^��//�:���Pr}�}�P��z�\��O�~9·�q�������)q3�;^���˂�O� 7�w�ݞ��Dm=0��I�/O���EBœl73>+�@��!�P�F̐}=Å/
�W�}��Ǎ�O��ٸ�ݨy��:�*6���w^UO��uA�v3��.2�,���{y*�n���O��2��t�{���&x�=�7�,
�ݾ��^�v:��'����7�yi�}�G��^�8u�O����a�+���7�o�")�'�ޒ��{@���-P;
�{dyq�4��AG��y�o�/�U1��Mia*���}���3�3���<�l�Q�y��T����$Z�V�]��A[�Z��E��%"C�xH��}o��fn眵��>�2���&w��L�-2��b�=/�w����~��Yhh��4���uzۡVn/ݞT.��"�c�^ȳ����E&��V�w ����@_���8'*<���̽X�f0�G40�Or�<�[5ڲ.���jImQ�x.Z���:�Pfv�qb��4R���ZN�����`�Eǐ-���Ӂ�˫\-+�>�Jf�5���Je�mT/�+k"�:��NG�e�{�Â�	�;�ѭ����{���=~�HΖ��t���7p*.yy4�<��=�#�l�����b��b�nT��vyB^y����%����_@ 6jH��T�'ŏ3����Uv���y��O�^o�#����0��~��|6\���h��5t(���bK�]��;ɹ�����#��a��Z\��
=�\���#_��$m�f�`-����D�Q�����{�ez'�LU�� od�')���m�_��y�N|jN�I�%��C�>'�G]ŧ���,ߦ@hձ11K�h�~;�&�/�yU��:ə��x߄y��%*�^g�:����I(nA�m�Ӳp<>��3��R6�SDTRך>���{ʼq�����N���˙c���a_ٵ�����*4z�<�L�_��W�<��l9;����F�UJ��֨�~۸�C;S����¾��v�v�?\f֏\FN��>b�Z�������*X�gJ%YՕ.�|5�K�n�w�u
N�R�}��4��f��|Y��:-�+�f��6t�cZ�6�;��ޑr�h�|��Dwӧ_
���ݢ��X�#�,�R`��Q]oW6x�L%�6m����S�����������ݗ�,x�<������)~Zo��q�5Sב���ǵ���?7ޮ�ܷiL�=�Zw�]�l
[X�	�.'!����Б����g����<�+k�x����L��^�+�4�e�����q�����r�������U윺�E�3�=����]�`��t�=;�Qcت��L���>	��wq����9���烶&}�����G�s�r�^���گ�[%Q�$���@��0/�P��L�7���(��U{�A�� ��^q�^�V��q��Q�<U�Qg���OH�`LT�"����-��L�gzo���6{���>G�z=]�x�Iw�~SA���Ӳ+����b�m��E��\r]���l�}�Y[��V�|$/y��!+�g�����Ǉ|V�nD��S!��9ޞ��Q��乑��tb�:����ɇ���̌�^��}�(�0k�WCu�'�������;}���}���Ā�Z22���Z;�&�&�ė��}����*����ٓ1�b���ƻ�����C�[�����l�Y�+�����Ѧ�� ��}}��ڎ.8x�6���]@��-:���\*��,�����Ά>�������J��ݺ��R�W5N���@2��կ~��J�$�ǃ�b��ْ���ye(
���1%� w��r-L�#T�.7�TZ�&���Ȁ_���%�����{~?x�]����|��g��ӚfO�j@U�{�`TC���A��6&鎸�Q��ZdV��l�|�{��Ww=�o5b=�����嚇|���_���9���g*I�9�+N}|�\M�5y[��r ^�u7�U,Ǯ�vc�ܺ����k���L:���6�}���t��zh���'����ꤕJ��#'Mk��!�Y��za�m>7ޞk� �W��Ϛ��~�#wߑ7�jy�v��V~��H�NZ��~��h��1�g� ~^�_�'�ÿ~%GN� Z�v�9��Md7^�_�=As��W���ߘY����:v��������ۅ��G�4�7�G9��]��7��q"��x�������I��{���Ψ��{����F�s���߲kK�w��Br+�F�S�˺�^�/p~�)Z!�6{���i�k�����}e��s���0,��~���_�V�M*����,�Y�l�
���Y�|Ό���yؿW�ܼW���>0�be�>EK���Kא3���B*8�Tk7{,�Y�Hej��oe��l��k󣯝{������o$��%]�,��H}a�9r;��t����F	��(�1,^��5p���č���xwی+t���,�}b����ٶ�T���5��b��we�F�֌�E�I��Qq�»��m��8|.���7�1��Ņ�K��ϗz)����_��-Np���cξ�:<�ۻ��t����:;�j��ax�Ʌ��o�q�}M��D�ݑ�4L��2&���������^B�����t�A)�{����j�l�%Q���ZEz�u_'JF)��{_>^vϵ�\/�~�'�Z�@h�(*j�T>G3�XZsK�8�U�ޮ��ɣ��R�v^�'�8�"<o�EC��/�u#m�9  �ޘ�^��dLS��ѱ/�Ʃ!�~�Z��/���;�Zݠ��s>T�3��\C��MC���M�h���>��?R��~p6�)����W�޹|{c*!*�,'�·�q�������4�d�����a�ZK)'��9麇�[�=y��5��}W��*2ƴ���#�@�5C�g�����;'�T�d���:�>#�D�%�h?̘o6����&j6���w^LψĽ�B$��p�j�{�ܻ�x��.�-(s#��_�a��x\��ǝTV�M/Ǥ�l�}���t珢�eJ���"8��/w��>�����~�WqR� :�q�vլI�[{nvl�W��Է�!��\��bO�U��S7|��U�\�m�Ҹ�s�<ո7@$u�NIѾ�rw���6��L�rʕo�=+�<�N�����kh���6\�%�:}[1>]G�}>�6�v�̙л'´����t�1p;;gi�b�)���}��W��x;���\k�9�^6Ix|�X��>�E��+o�'�%�%���@�q��ol�HO]>=�n�q~�C}��a}�%"����ޚ�A��4��rMz�5��W^�:��7���/_��o���_���U������e�(�X&�7}Ϫϴ- ��$�%75
�T=��Ac�^*^�'�״��g�,Нǳ����T�z�J�~�h�̀P:�TQ`L}M�
��E^M����<��R�m�>� �;��gA9�t���[���(� 4z@�qU"`�\M�X�;��:�M`�9Ӯ��C����n�m�Ͼ�B�g=�t�)�;�>�I`@l�څJ��^��=�ي�]觋5�>�9��K��,%��hM§kŇ�}#�Uz�L�t1���c\�	^�*�q-�N:�&)�xv ���@�sʻ��g�.��� �y�?�ُ�G��?��§�)Z����a !	1��?�|;�\� D\���E�"e�jY{��
k���]�F�5�z2 ���#$��[���[�P�"�!XU@�@i[�.�����̬�!�6�R D^�#H�(����_e��&a��y>sK��¤P�Ҳ�T��{�Hay����#�pJŊz�8[�d�"�I��s�J��c� ��x���� �����bV�Y����N���p{��ğ-)��@���=Z�H'�@�S����Dvx��-šw����d;`l��{	� Y��P��І�w��;�s�q�u�G���r }���" ����Tr���K�X @�E��n~Ӡ�@����d9�S��{d���;�ɯ0�T��Dtn�'�~i���y]Q��!���k��3��+���y�����;�w��dӨ!�@݌���.�����O�q��j+'���4u,�. �:�W"��"ɹl���1V�h�2�=}���rv=D1����~��Lql�B ��&��qT��D�Q�D}���}���LJ��5P<�L�fX|K��D[�͔��!����B>f#�0A`��#c�p�����jԑzLL�z�:��^�w4��L�-b��$>E D\�g���]��E��`}6=� �	�|4~f�ƀ|MF���rP�^�Ҳ����n8�N}onq	���jS�C ���H ��sw[i�7 �w��*���C�B �+�`�c�>�i�e�3�yx�M���ûө/d����$��%H ���8�-p6�]��� 2!��;�<=^�9jŵ�:�"��]a�	�<j]1 ��$�fN��jz �C��u^w�X*,��X^��l	 "/���C����<��:�����C��R�].=27mf.��B��,]5�D�|I�=�s���ܑN$`f�@