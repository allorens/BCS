BZh91AY&SY�����_�`q���'� ����bI�                   �U(EW���$Q*�)IE%R�")@EJ�I"�$�H �d*JP��TTT�T6b�U�CMZ��6�*T��:�*�PRQQJ@��B��(P�)EJ�"�@PJ�! �"�J�)P� �����k�7)"I` mU*)JX ���D` -)UR� �A@*U���UU
 ��I@)%JE �DR�9�  ��A�   � O��H �Pw��{�>ѣY���c
�hQ���� :�e�M�X�e�۝4�ʺ���@�����iKb�Vi �"����D��}|�Jـ��_sP����f�v7cm�:wggR��Q�*�
������+J}<����f���秸u���y��ς��G����΀z��UUB)h�Q$��䤒 �{�<����#M�^q��]%�qp�Ck���+ր��޶!��E'i��^� 5�<p5@�s�C� �8:U��p�^���^E	"��ʒ"T[�䤊 >��V�h���Ź� ���ׯP(�4O8�vk��y�Q@�+�z� �CS�w�J�{Z��z[mh��;u��P�]�w��]h����*$�T��$�� `� s���P5���ypz@p��W�m�h��h�){���l��z;v�} tSO9y�P��z�/P��u^�s�PoSp@z3ƆD�*H��aN�����)( ��|zӴ�p w�͞ �q�h]�h�:
�� �� r�� 껊 ��R%P�yb)Q_>RR@�=�=�| m�� h�� �̻� �t� l]� �� ����� W�p i�
��EH�n�J�R���)H  �=�A�,]۰�` ˸ ::����m�� 5��;	�@��G@*�M
�
lҪ��I��R��� C�}�W}� �� 90� �v8 'p �� ���@=��O a�� �%H�${�DI	o�RJ@{� �V P6����P  `�  ñ���� ;P �ox 4C`>*�� � P@*� �  ��d�)P�?T�b �4�&FO�bJUOU      �� ���0�4щ�CMF!�5=�AMU(4�4     I��	U �4 �  ���������4�i�L�i���H�O�����?������k�������&��0Y����Z��zĝ�D��%���x{��{��P  �J�"*~� AW�Ux�'�������H�����>T��(���u$�M� (
�����������DP�������!lm��0
`�1�c8��.1q��\i��.0bc���.0q��L`11��L`��0q��`��0db�8�1��bc���%38��0`����.11Ɔ11��bc �&11��L`c�CLLbc8��8��0q��Lal`����01��L`���6�b����&1b��1��a8�1��Lb�8����L`�1q��Lb�8����-11��\b��1`[`����01��L`�8����1q��`c���&0q��)�11�lbc���&01��L`c���L`c���&11��L`c����h)�lc�bc0q��Lc����&11��L`�8���8��&11��`�8��6�`�8�1��1q��q�`��&0q��`����b����0q��C�0q��\b����.0c�.1q��1Lb��1�b�q���)�#�!�\`� ��\`�1�Lb����.1)�1�8�1�l\`��.0�L`����.1q��8��.0q�c �.0f1c1q��C���6��-1q�c�.1q��\al`�8��0q�c���1��\`����1q��e�1�S��1��\`�11��b�����.1q��`�1��aLL`Ŷ0`���1��8Ŷ0`���C�bc1�LL`�0q��bc���c6��0q��L`�hq�Lbc���&1q��q�`�����Lb��11��L`�8��0q���&11�l\bc8��F&0q��Lbc8��.1c`��.11��`�F8��&11��b�8��11���Lb����&11��L`�@��%�q��`�����b����0`��%�q�3�Ķ0q��11��Lb���.0q��Lb�8����b����1q��cbc���11��\bc���1q��bc���1q�L�!�[`����.0q�N4�Ŷ1q��`�4�bc�8��.11���0m��b���1q�c��b�
b����.0q��\c�0q�n40q��\db�8�1�c���0
bc��1������.11�����1�0bc���1-�Ŧ0q��bc���c11��\b�8c��1q��\bc)��L`��11��\bF��&0q��`�8��&11��01��Lb����&0���L`����.01�21q��Lbc���1q��\al`���#`8��bc8��0q��-�1i��8��.0c1��L`�8��.11���Lbc���0`�#8��11��`�1���11��\bcc��0q��`c���01��q�`�8��01��bc��c���&0q�0q�01���bc��0q��\c���.0q��bc���&0-�Ħ&0q��\`�8�8���.0q��bc�����\e1q�c �!����!�\`�c0q��b�1��\b[1�L`�1��\d`�1`���Ŷ�0b��0`8�1�[�LW�0L`��F�\`��.0b�8��1����1�c11��1q��8�1�c�c�0Lb� ��b�@c �.0a8��.1`�1�c#1`�1�c �	��0b�1�8�1��\`�1�c�c1q�c���.0`�1����.0q��8�`���0b�&0`��c �.1q����1�c-����\`���e1`��.0`��1ƀ�S0q��0m��Kf0
`��1q��\`��hi��\b� �0q�c�c ��G�0L`�1q�c��\b�1�c�`����C1b��-�cL`�cBب��Fc\`��Pq�.0U�*��G ����1�Lb+�q��1E�����\b��q�01��b�Tq�0U���G�� \b�� q�0�	�)�1T�"8���Lb c\b�E1��1�
�38��11��L`c���01��bc�����&11��0q��L`�8����&11��bc���&11��cb�8��&11��bc �1�b� �0q�����&1#`����.0q��\bc��!L\b����.0b�1�����b��#�S�B1`8�q�c�$`c�.1q�c���.1q��a��8��1`���0q��-��Z`���1���0q�c30b�0q��\`�1�����1�c�)�`���\bc-��b��1q��0b�#���.0`��.1q�O����^X���D=�^�Q���ytU�[�j����O�d��A�B� <b�梃v��M3��l�2�,�J�w�܊��3ז1�aef��rlj���!݇E,Ms鋴q[A�a+���������H����b@�]>�&
{�!���ke��@誓�S�E��P��J�nVsZU a����QI��U�7�����0^S:A�w3zG|U���8&���s���)ɍ�TCf����%\�MyOq��E��ɶU�7g�lWe���N�L����L�Q���A۔ch�t�A�jh��*x���fI�2�S��F��l9���%��Fc�z����1��b��UI룐�f�'�S��εC�C�/J���.�&� ];$�cBI�h՝�MK�f^�r��X�����]C�Р��z@�#qQ�o����\�R�����*V�tol�[���Z�F�����TOr��N��^�z��0*��9q@˻�8D���Tm���p֒j�3aу�o��W�E�E�s����F��M��:j�Li��=p�۩��s.��BRa�i�n��;m*Tҭ얍<ݩ��#����b�c&Kk��[{l:�oi+S
x۠��u9��+-b��ː�ڣ.�M*+���2��7-6}�,�&;�(�kSc;�k�a}�xÎ؍�;!�"��4�ѡ\\�9��c��"���5w�.�QCt��6�kn�0e(F�&��J&cK��-�*��7u��\�V�r�4"V�PI<5�+�ˆ(�X6��B�3r� R�<�2U�f�)n�Ү	��C��Ƞ06+[n:���Oc��*��MK��M�U/Pɸ�igUy�����%�Ժ:h�Z0iT�ҥ��W�����A2`;�[��GY�QVl����3�4Q܆�:[Vf��m�1���AԤ7`:^�ܲކ�ĵ��Ҙ���gb��4f���(]J���x�-�N=�iW!m+&�wIEɼ��VFS�F�vM8r�0�r�ke��ޛ�(74�J|�ܙ2i���j���l)	�yk֧o-��%�r�v�oKa�2��p��&�KYw����/�P���j���thOL�YG�c?Y�l��=����4�iۥ�F���5�X��͹�x��y*����m$��Q���D����[�j��ͱ��򔙄c��,v(J���VWh}xE�K{�M���Jb��Q�kȹ���p��j%Paj�o�Y��ɺs��βy��k\��[b����Z0(���.,��^=mQEɱ�٪�ml�tx�}Ʒ�2*W��F���ER��Y��7
��8VĤV�Ni����ݥ�,�g%�������$���h�T+F��P�+D�"sJ�F=�HqQu���n򝢳�@�"ܮ�-IyY���[:�mV1m�kdD�xk��n��$�����Uً�Z���2]�ī%M��zZ2���2M�ifYz �y��OK���0N��.�.n�Df�2���7j$XF�<{ �{%�<,��Z
�ȥ�c���Uu�WDzK��Z�~w�q�K��H5�0����U�CGHB���U�n����X�.���vW;7�$-9�ʼ������ș�W �ƺ=�B-I�c�In�,���d��E�9a&bF� ��K�w*��ȳ���1��t��HF��F���En��C��UmK�tN���ZK����#[9��55b�2266���y4�6�����8���� 5d��{Kj�֕�;#ܙ�2Cm�;�/[#F�V�!P�b�W7+�ٻ�ZM�W��������c)�(M;�n���ZK����h�lK�$Z��/Kޓ?m�*��L�c1B�lR2
�o'���ʩ�*�E���7�%껽�w��^��e]u%�6�e�$��{m#�5[q��l�(�K,֧B��x���^eк�=�k7�ץ1A)"�6�$9Kh�$;�A�ݡI=��í*%�(]�����C�]��VJ��q��q��FXUx�ʻ���ʗ��+t£���:c�Q��+2��{�a"�Ȗu�x�ͬ$�x��]�Nm;�G3$U�Sa�5���m����;��������;��X7f�D.��uTP���R�P/�-����	\�l��f�.�q��4]��Uk]�w�5��Jضj53�����^�;��M-��w�Ҕ8I�gX�N�0�x���RL�,��{�U�s�La7�E�v|Z���H��}Lm+C.d)����ՌIX0*VQ��u=�a3!Z+Zŏ�ζ�	�a�j�6VWq�ׇ&a��I7e
��s/%�Xp��*mndo!��Xs��͈����d9�W�v^�.Hw�eՉ�`��hg��q��e1��m	x��yuU�jp�WDY2�b�r��ֺRj	�Fh�8C4ۨ9�*�į�uB��g^�0N�-�
M�H��&�JA�6��b$L�bC`��!9�Xt�.�.�o;�ݗH��&\;5����W�����0͂7��y��(;*�<s͆��f�9$��<J�3��7��CYR�ɷ��Y�x��c�c��լѲ�9H�n�
�("6i�we��ډ�3*A�T->	sy�܋g�S��h�ޝ�*=���.<ޗ��#�3 �RU-�lJ-ÿ@�u�;ҫ;,�92���kɢ$�G���h�bOt�x^�m����	c�)ƶ¼�&y�0����=,h�*F��Us�%u+���%q�I���˭��ʪ�q9VJ� u����o�=R�3Z��NW����6�q���k<�Lb<c�ɪ+V<ܺ	�1�Ԑ�����,�KTV��x����<oq �WQ��_ْ�S��Fr�Nc�ou���qB�g5��
��c��1��h:��b=4e3�*]]$z je�"�xe*1JD���'5G��S'�[�{�H�i�M�<ZY����$e=*�L�XkJ�g-ӈ��Փ�y����m��1� ���{�����д����,���F;���E/34��Z��\��mnRw0�Q�T�E���K��H��x�`<5��k��V�=@�l�g�X@(�Ь!�cb�a��œދӐ�f�͖ܽ1:�{C��#�zA��S�6ҹ 8�)���4�|��c���uJ�vo��PJ��������껌�0p,*t��7f��x���/$YR'�4aM���.�"��o��/�_i�[��n���ɍ�tys"�)^GB�:�n�[wJ�ɦ�l��e�3�BZ�u/�Q>�O��c3X��,M�wt��{Z+5��t���s��\��a�tr�s�YU<s]]R������!�	���}O�ѭ0G[v�J�}]�w%�sjS���)�-�0�u+4H��en71f;�t��	1�uV/Or���u��_]���sV7�&=�ƵZ�j��*����+1�����f�!K1�c�<�����s�!vġ��n����:7I`�FfR�j��n�A�U%,L�{����$r3��K6�qL�S�m��[��>.1��Y��1q�[8n��m-�+�U�z������8��{t�n�}*�����9�;����%�[�R�IL}�K;O��V�}t�!2�ܩ�s��꼶�,��[�*5�DN�ּn�*���o7�\�k����3XrL���Xû�(�r��б{�p�or���tE�qϮa�ʆ���yٹʛ�1�.G.��	����Y�#�"�vN�����l�+�[�J�PiZ�`�sn��S�.��I�)�ז�^hNVn&-H�`�[j%4LZ{OK��׺��o.�/M��|Dn�]�`L����p\٩�fK:���o<31f��֜cNd�6���x'u�w��ob�ͫ���Q'j��߮
wk��6��AZ%���9��Z��s���Λ�@���,�4#62�e� ʏ-s�.��C�{�y����!��-8a�ޝ��`��\�Lt���V���u6k�J��DK���wmr�yF�xV�&�L��*�Xh�%�gٷ,���'��LMm��򂲨bY��/�����=�nk���nFh�q��һy�Z1�w	�,�Mt�T�X� �ik~Hhu�S�b�;K�7u�q-�i82����-�6���rE,��f���"�cKMޱ��Fhʺ�o���n�)����-�UK�v���Q��H��i��6#�q�ʨ�1%KH~*�oA�	QD���N�cx���
�������Uqh͛�j�[W�S������T�Fɖ]Ln���]�Ul�z�l8/��#�u���J�ѝ�+�[�L=Ĳ�v�Uk��ka��7(���V�3��ӈ ��f� 1��S��:Cr��I\#$�%��[�0���}��!��>��{���e̋U�M[m�=[���,cβDb+�� � r��s ��Yq6vy�<{j���r���������M&����8�V�75X� �D�L�;ZxĬ@p�f��5}��u�ud⛒����n��F7h�W�&lI��81�9��Wv�:��*v�飵�^�B�ʊt��&�3�#��	�fbx�]:���d_M��V;$�\�w�)Q�=���<��X�I4l%J���ۮ>��y�	��J���M��3I|K]K�����ݯ5(�!v�W\"�E����V>�OF\es�B@])�̼�}ծH�K��A��6�JԨݹ����S��s�=S'k�8��P[;��-��-1��맻��ax�l�{�U��K�X2"�˃b�34�o2�v�|q��wj���Drީ��Z���ք�غ�E����跲s��WS�nv��Gw�i�h񬀛�������+:PH��m��VZ��s6�KMlx��WkiI(�8�.�sr���q�Y5#�d���X��	f?�*��5���CŤ��d�N���:vͲ�&�y��F�ǌ=]mqh��G[�c�0Լ[wOR[a�Xy>]ɵ��T�6',8�V,�	�ai[�E�!Nܤ��۱��AN��0�p���jKEj����C�"��^!gvfV�����b�nU9G2��J�L�Xb]���ae{\�qc��$	��L�n������b6LӔ"/��e��ʇA�p�`_���O��kO��^`t�'K%�xS;�Q�n�gY<p��ht�'���r�2ܮ���x�Q�*Eh�%�G4�Ĳ���=�q�>��a�2���(�Bj��<�7KFq(��+��>�d��SV5��皚ɲsFB�r��Q�w��i,��#�� ��75B��w����did�:M�[ӹ4�<Ȳ��)�'�lֈG3���7b=AP�-�L�x�P�Bnb���_�g,�9�ng�Ι����t�N���h���|2��s�s�� O���y�6e7�'S{9C��)xm9�����v'紧)�ڳTŉ(�*���d���	d��n��M"�D�$� ���m;�faV__=捙p�g4�-��@
  xK�I�p{7�ٰ�"w!�p�������`w���vy~��^p��|M�Ǘ�c�&�'Y,���Yt$6*5݆9�9MGj�8�����Rw&�o�!\I"��l�N���|\9g8�Fq�:oOBa6u�%�v��l�p�Z7áZ������r�<N�ʶ��&x�b�xΑ�8��u-��'M�������x�/����9O;�v�B6̄C�\9���r���Q����]�Zƒ]���2*堞OWiv�¨[2���Y-��i�V�JɒM�*��l���I<ϴ�1���sHD��ck/Fg.3�r�f'�l������Ӝ-�0�l�]�;ў9�a�_¬�
�;�6�v�r�9 CZ�)��Y�a#i�9@iL&e#t-����F?B�_$Os�<m��U�-���q-�mcL|��*T��xz3��6N�x�i^.Ct�^F2���y���"�8�Qw%������i�p]q�`�6��6e7�O�$�iնU	���-Ba0�T9��B�S�;�iΑ�r��_ո��Z�'k5<Ui4E;v��͓gi'����'���fզQ��U�[|�]�,�-NKWړF#���*n
l"p2���@Ox- �J0p�vZt=��pΏgY:Wd�Xp��Z�&��r�^�0�!��v�پO)�4�yӘg4vd&�;�%�E�,�G�+s�B��9�㳇p� �91����v�yRv��4��Z�N*��]�f�)J�i��ᗂT�Id�n'k��i(	j�f����Y���	$�Q�:�q�� �A����6�@8��6�TH�b�Uk�6�k��mgt�e��v'���G�|�6�MZY-c�R��>(�Br�eÉײ�D��C�I6�9���Y�K/┇.G.>ݳ�ff��g��xE�ӖS�
Ű�(���s
%���gE�G��S����7̱�E��M&�i� ���Q�I���5��ĘK"��yM)�ڤ��7��b@�GT�V:� P=�y�[����8�gb���	�.�'t�5X%+�i(�(�e�%�%J}+�ڎ��p����iT3��R��*�7��zc=��o'Y�'��	�rfP�=���&����]��QY�골]['Y�/��.��K;	�um���#սg��9���fC�&-<T1���^�M����I��&���T��~<	�aS�����l!�&�C�����M�{���x=�чN�y�w��}�iН/Fj���n���6$7K�@M� ���[�u>���: ���� �a0�Щ����M�����Æ�4� �2�4�#I%��ou�E�Y�7����9�����L�S)�#l�;f#ݱ<��xv;���Mv����Á����7Ͳn�9 
z�gi�+�P�2�\b/
�w���q���M6v��J˸Z!�g,��w������x���ߠ�������?�{�k���I$�I$�I$�I$��W�n�t�NĒI:A$�I$I$�,I$���$�l��ML�I�I4I0I$�%�$���$�N�I'KH$�I:X�I'	rOrM��;1�yئ�S�M�Ĝ̼�-�wj�})�Fl�/�>=I�د�y���ve�4�1ٚ�Zb��s�ͼ���x������=�R�O�"��=T���j�;��}w��0�ꁘ7<L={��Y�����軫n��Κ�:S*�olb��>e�R<sK�C�0��^u�C����LMv.�m�#q}[��Z
��f\��g�sg�u��t�v%�M�*��m��S;���[�d��J��+��k��x���᱔v��G����-�D�r��
ۑ��:���A�/oo��-�Ce��K3�Tܶ`��$R���f�������D��u�m�\�QV�^�ݾ��2�P��)e��b�f����g^B�5���J��[�IX:�e����X��t�e� �ov^���Q�K�ܻ�"r��S�q���e��ouXSgIq�N�>dH�`�+S�����`�;N��*e�/���5v�l�G(M�.�g]Wct�Wrr
�]o)D�M}N�ݼ�^��fQo;',��#;�e�ۿ�+�ZϮe���KeL���Y�|�k��� ��������q�O�i����O�<�LB� ]���Ƕ
�X�A+l�Q��}ہù1�Ĺ���L)�9�m�9�ʛ��Nx�ҍ��J�*�s��H�c,�wn�3����S���D��$��hڀ!D���-��N!�J�6���)7.t�Z�)����LlE���k�߯��/ݡ�����
Y��뽻;.Oy'��g2��MGVٺ9�E.�05�}b��̴�>U!����t�崔�V�������{�����2������PB�Wn���p�:���W^�����E�J�m>�!6�꿥�QZ��$���t�u�Uң�&�n�(���0�aU�Ww�)��mq�fm՘n�Ṋ�^��K-UR1�.�V86?���d�6�t�X���yz-�m�w]�hv\��;|{O3�W5�8�t]K��V`�nH�GM��d62A,ͭj������)qu�"��|�PYY�^�{395}U�z:���s8rm���U5�P�q��p��1|�-��`�ɝ.d����w�h9.�<�5�Y�s�r�mǍ�۫�1V�ìJ;�7Un�����}U�5~��emv�-�=Gw���Ȝ��ڬ$��V�u�ӎ�kY�����j���1u���v��=D�ѣ���m�dU����)O��+,�y�Ƥɕ��|����S�[Q��]LuJ��j��n��#�Zj:�u�M���';��Y��l����]ׁ7��bpG&������ހ�W�0Z=�;z	C������G��hgk�ӄn���k|x��og�6��-����ʙ�lc6u�Y�%��DD5`�;5Ճ�+��1��<�]q����j�\Êu��)b�ȟf5�8��dE���;�8��v�j��ՙ3�K�:��q!��9,׼Fz��Vq����/����Z��N�OR��L��%H�ׯ���k�"۝N�,�&�G��f������\Ϲ��w�$��b]�s����1j�l�2m�z�`���w����X�àa�W�_)٬�4gpދ���\�]�x�P�6�.Sl�祥SVKߵ�
�PD�c��8�Gq���.9Q(�R��;�;���e�]���_=�ܒ���w�����C~�=�Ss��`<���[9�
���h��(dm5U(�C5]��j���7�H���(�>v�ZQ���N*�|5��/�[�h��ޏz>�f1jU���1y2�-�soM�(�j�Z�Չ�.��A�\����!y�,cm�ӮC]}��:��p���F�.`C��N��gf�T9C��]m�RT�q��"���|�#�WR�N����W�������C��Zٱ:�]�{z�(o��0��ӓ4#�e��2�����|ž�]>6�p��wұ���fX�	5�� �Rk�(�#��c8�2��<7.�q����otR���ɛσم	}3�=Ǖ0?�/0�vj�c��T�[j�+V��)�Pہu���D��rݥ� �Vi]�7I⳧	�'��!�.q]���5�f��l�$e�Wn���β��w��%�yo���#�]4��W;y)Tf��k���-�V�k9
B��*����#�}U���H;�W�Ρ�tY}�i����auۏ�cmc<L7	�aw�|3��i.l�8UI��Ρ�6뢕�;HtG�{U��S+I=�Du!Iw*�c�I�m�ow.j�f`߄=ʐv	.���F��L��D3��)��ޠT$������tt$j�e��
�����d��;�ה���Z���|�WS;V/�ٝ;ӂ˭mѼ[�Y|�]EhU�$�i*ѝ���(\�(N]ʎo��=��zbs6�wd�}ۉ.ot���.=�J�����pj4.#�:^�v�7n�z�u�iUT�;�b>�j�io[����G����о��("������
��0TZ=
��w�Z®�R��B��o8��/��V�u���2�D;���u1X�S�=����.;���"Q�w�vf[���6���x�h����I�9��¹,�:�,sH���yRn��`MW1�Y��-[����=-`�B�����Z���F3V�NL��e�(w=�E�Y�-3�\P\�z �X]��*�s�6�)��h����<�����Z���7�U�Qe���\��U��k%S��e�^�n�æX�X����9\l�N�e���Ot��ҲWA�7L�'����K�K�}�Wnޚ�jt��O\��+�;ts��yƄ��� �zf�7�,N���+w�	t&��ǒ�L��ۀ�:+��<W�a�R�w�}'7:��͊s��Yw/:owwqwQ��3��)��������*���Cg��N�㇛�w���	N��G��9�fa�h�Ҿ�vz,2Iǅ��N<z-Vd⺶�ݩ���w�p\h�|r�yu�I4�u��g�-D�#ْV�ۢ),�D�f1�h�c�Z��t^�F�$7@��U��ںv_-\Z�wFJV۩�xKQtٗ�m��0��G�l�o'A�w�%9��펮8gfӮ\;Ů��'K\����Ю��YH����p\y�W��]a|��0-|�i#�:ֹ�;�e�x�M֠]���05m���p��t!������U���_{�i]�![=�h��h�6�ޔC:8ݷ�z^q�v��S=Z*���R�p��-c���U�N��Q���Ԙs
Ǌ��+�s�s>�]��O5Al<��I�ܖ٦�����!��7�R�$�K�ػ��[8G���+���9]�;�]��7�x����{&r9G�\�YR��*e�{`���e���2�+v=�/:��EOK�1G:�����N�J�g�k��s��Ydep�#�і��.�Y�bu\����W�o ��;��a�r�CÊ�y��;ܾ��&��{I����ijs ���������R��6�* �(n��䆬T�ǹۊһ��I�5A��U[1f�m.�i�&�]E�S�0m�\��9�lCLG�Ij����^�y!�s�����o�0�����C�xFl<h:����.�����v�O{�����ע�#HM��u<�b���R%+I*�RRt���i�;/��ovK3������g�W�F���t�3�S����S'��=Lq��6�PV2rT�7��6���8�A]B.)B+}���Ծ��ڱ�J;c:rn��������ڋm�޺���bT��I�sռ�Wa%:Ҧb�(ND�vH>5j)P� ��]9���Q{M�[�:]ƛ��b��儓e�_wFOX��
m��P���^�������񧀠���GVLS���.�ɘ>�$t^�q����o&�i�uݷnEw��v���7�u]�/���[��ߓ�R�ܬZ�Wö9���2p���X;3�k[�J9HfT}��)w,�cw��6���]�V���N���R �*�:;�E��n�*Tq�a"{��l�Ň����a�gNG��n3ku[��tū�s1C;Flj=9�}V���=�����Ŋ��fS��d���O9�]!,vV��z��l͵e��N����utmu�9x6d)�L����2��6{���i۝8ՈL����]��]��6�n��u�[���C�����Ee�_L[�i��
��]>�nQ�]\ȴ�^S�o���R�5�s�u�O[U���0��������S���5v��caY]����w ��J�C_PПe��6�`y�f�E����7+u�ك�r�;������#�����[A1�t������-�gq[�E���ҩ7��Z���5VԚ�Vʜ��J�w����n3��������ݹ�j�7
n�����[aE���Цm6�#ʜZ�CPT�o���ղo(��nT1nn��D�̆��ڈ�5+')���q7d娗A�c^nP����8��
�f�
C}�o4���,./+��}[�G�4.���PŚ�.�M�\�憯����d��Ums(�o+��a��X�sgt�7�r�ֲ�j��'^v���W�ͳ�X��2SV�7�#�WwV2�Q�f�6��ĬR�7�`�70��k�9)q�����g=c�kZ���)�q�,�[��##��oh�-m�OgLxy�79�n�ud'^7f�um
b�pV�
�+uV�%���]V,r�Nm t)v$����8o�yIfk��4�h��g�~̫f4W�)�Ĉ�=���;`�@֋�;˭�|�s[�MtW�bT�#��n�ӡ��d�V��68U�EO�7��N�^�/�b�wg1�.BS��V:��
�\��mZ����ʻ��K��j5�yP���q]�P��<�Qy#Y�Z�}�8ؾ���M��ff�ó����->�nvJ#�/WTx�7:koS]̺����E]��f��{�Y|��}Zs}��wrgX�����wi��W�MMU����$�I&���\����.�/� ��)YW�ћըl�����iC��u����=��^7;$���%yoS��C�%�(:���G���ǎ���o�����Ҿ�0��T������6��?_����������+q{��b�r*+;lv*d9+t��� p�P�A�JN�DByݠ�C�}�z�+��!�ꨑ��w�,R�Y@�*�7��3r�2�$<���m҇�`��.���}`C]`��;{��ہ�	����z���/�ȠyT����wG��u	�B����Z����\��8u�t�F�[�pWy.d�����w=��w/�_�#�,0�W�}
ܹ)����+�(��'@���o~���限����0���N�m$T̹f�ٻO 5�W�)�B#�v�� L��x �2 �ǃE�����|�����>��}���z�H�,��,����;��� T�.N��e��A��q���ҁ��	q��	�!]��T{�\�yG7+�p?�AO���>("(�~�?g߳�O��9��()�ȟ��?�?P���?}�7��n��w�j~�λ���2bJ�t*�l���st�����=��q�zjż�fћ�q��0��6����:�h����3�`fIř/�3	�/r�KcT�� ���]I���[d>�Q,�v+v�ْ��t�:��:�VT<���Un	�]Ԭ�W��8��9��;�*��;g\�yݫ��˙#o&X�K����k�ty+���:'�t<�
�&hǪ�t�l�b�'X�3��$^ຄəb��M�j���îEu�v$��Ӣ5+3���$��^���M�u��`�jR���w"3�|�����U������'[CU��:��Jġ�qӾ��S׫Kȡ���z�pI��	q�=����W�*E��Ѫ�����sn)�Ɍk$E�RZ2���{-VɎ�b��
�$���D��eaȻ0�����Ұ�:ڮ�_oB;��ACZKꯏN�]���e�o� s
����A7��W%Z�������$-�3�L��s�;��:�e����.��� �7Yy�����.޾��N�r�V����q(�nN�V����gfv$�ӼAP��^=�H�%\�VD͸�g����z���w������뮺뮾��]u�]u�_]c��뮺뮺:�:뮺�뮱�]u�]u���]u�]{u�[u�]m�]u�^�u�]q�]uק]u��u�]u��]i�]u�]|tu�]u�]u�]c��뮺�룮�뮺믮��[u�^�u��^�u��뮺믮��뮺믎�Ӯ��:뮺�뮺뎺뮽:뮺㮺�N��뮺�뮺㮺Ӯ�뮺��u�]u�]}tu�]{u�_u��u�[m��u�]u��u�]u��]u�]u��X뮺뮺��:뮺�n��n�뮺�?�������_i�j�,Ám�oxvn��9t�qm��}T4am$Q�ٮ�_}R�oVk�^;�"Ʒ����|s�}t'ʪ�s�W�VL��3���]������#K��CM�
������#��=pU)k_@S���S&w��Z�Vt�D�o#�X.�Y��v��Fn�����d�ۡCBF��{@�U��/Z�ob�us/z8�G��f�[���V@���H2�z=To�y�T�cT���t��ƹ�҈%���7;1�o�H�z�:+�/��B�n��E���'N�n�ؼ�DWx���:���U��� Iwc�y���m���5F�-k��hf���֌�]V���튡���q�*u�y�8N�F�'�V��B��6+�=��yM�����c����&���(瓸^��5Ŝܘ�
��(&��庥Nׅͧ���i�O�@���.%[-T/�y۫i�fgt6��0�!C2�GFdF��/]�7�A9g.Q�qtW��&��_ph"K	��>�ǧ���]u��]u�]u�]u��뮺믮��뮺뮺뮺ۮ�뮽�뮶뮺�n��]u�]u�X뮺�N��:뮺�n��n�뮺�뮺㮺�:뮺�뮺ۮ�뮽�뮶뮺�n��N�뮺�㣮�뮺�뮶뮺ۮ�뮽��u�]u֝}tu�]|u׷]u�]u�]u��]m�]u�]{u�[u�Zu�]u��_[u�]u�]u�^�u�[u�]u׷]c��뮺뮱�]u��q�\u�]u�]|u֝u�]u�]u��]u�]u�]u�]u�]u��]u�]u�]��Wu�W��ݞm����鸄��[��+������Q�/v�ὸ��H�]�z��Տ�!��M|$��a��#B��*�e�~�k�lR�h}l(���֙]�9�|׸'M��G��M	�2d7w��t�m!L�{{��n�g������xO,��LY� �N��S��KyA�i9Jm�$��1n�*J�ʦ��+�Nks%�x����ɏ��urC*���Ŷ4�,���l��n�^C�i�ie[<��dZD���țŒT�HL�;~���y�)�7[V�����Ǿ�KWW��K�u�ۚ�m*'n�M�o��'ܑ���[�\��I�l���%��\6���t25�r�y*���,�R��|���0�X��v�n�W5Xjauή�v�t���Fō �|�ٍuk�m�U�t��u�e�4��W���-�wV�;%/w)��A�x�ĳi�v� k_)�uoU&��u9c��+v�Qn�)�*��$)�ʏoY�,�����UB9HMW�j�������fTi_-��v������~^���]u��]u�]u�]u��]u�]u�]{u�]m�]u�^�u�]u׷]u�]u�]u��]m�]i�]u�]|tu�]u�]|u֝u�]u�]}u�n��n�믎�Ӯ�뮺�뮶뮺�N��:뮺�Ӯ�뎺뮸뮺�Ӯ��]u�]u�X뮺�N��:뮶뮺�n��]u�]u�]c��뮺뮺:뮺�:��:�뭺뮺믌u�]u�]|u֝u�]u��]u�]u�]u�]u���]u��m��Zu�]u�]u�]c��뮺�뮺�n�뮺��u�]u�]}u�:뮺뮹������+�<��F���d�AM2�ݗح�%Ml��4�q�ͫ{�z�t����lH>����=;���
��K�I�W37����T���an���j4�
ޚ��D����xg7�j��
B�<l�!Ї�}��"uX���s�WEz�D���/�jttk�%wV,��f%&������z�*Sq�����X�M�ںsIWVh5o%BM�Xoz���qo'u��9\f1G���m�a�y'^�r�wC��!��.�ފ�=C�Awt�ףsL��\�q�h*c�����,�.c��oz���$���ac�,�҆��ɪ�Ŝ�E��l>��oc�wHO��1�	��f8)�bt���5hZ��k��Ag�_\f�u�Űv�5����W ˞�87v{�U��l�Rm�m���6#6�j�}�L��O^�;�r=Ԣ�������թ݄t�-�/��/8��7i;m��»�%�
��n��U�����B�Um+fLK:�*o���R3+����f5Jv��o�\m�T毻w�3��A�;_tW�3�֖�t�����o)
UgLje�v;+��t�g�{�}eu6u�z���㏮��N�뮺�뮺㮺뮺�뮶뮺뮽�뭺뮺뮺룮�뮺믮��]u�u�]zu�:뮺뮾�:뮺뮺룮�뮺뮺:뮺뮺��u�]u�^�}u��뮺믎�Ӯ�뮺�뮶뮴뮺뮾::뮺뮾:�N�뮺�ۮ�ۮ��n�뮺��u�]u�]}u�:뮺뮺�u�]q�]uקG]u�]{u�[tu�]u�]|u֝u�]q�]uק]c���m�뮎�뮺뮺뮺뎺뮽:뮺�Ӯ�뎺뭺뮺�ۮ��:뮺�	��\߻�q��ZCH�V�vNqs�e:��Է����L���U�q����-]�)��(�+j#j��N�H�ź�15�Çz�p��<�ď��x��u�B�P��eHS{w�H}[�7x;��\$�n�w��B�r����kSv�r��%w*�|���s�
ZqcĈkgf:Ժ�[��蛨b��i�b+���V�����F�ǁ�2��}[짬�ݍ�B�3nu�퓒���Y~���M��]�{]٢���Mr��Ud�)�*7����zFP}�y5sk��Z���H�(�/8�5¶�m_�l2u��yN{%�<#��܊��y���vma�l�<�G���El��b�D9R"���T(ڹ}��`��J� ��;�����;�R�}ú�c8�ä�Sxm�Ж9���X�����4ڽ��fQ�̅�������:�gU�R�!;�R���8�m�:�6-vv��t�E�m	2�Q�W2�.&����J��e����<P�}mi� �Ci��Bv�ojF��gc@v��3M���)���>���$��&�B�z�f����w"��F�Co$vBΛqȵ�bb��Li�ۥ�/{���^�R �Z'ڔ�00],��G�(�k(L��?{���^���'�zE�3���&e���JFh��u�?\=� {)��z��{*�8���x����v,ePW���Ò'^���Q�wo���P��M�ueg`�UJC�����B���ZS�ټ��}�@�ց�L�=����Dv��bx����׏�F�n%�L���r4Ueۢ������{���*�bM�M
���hX,N�h��.��UX�m�����C���V����+Z�G�<�8V��A�rOS�n���*�L��#T�/=Pf�[M;5�t0m��qL0�Ҩ��
=W�.�H����	���\���ŵ���{�+8G���W��&��!��vd�����/��xneZh��an�pO��s=3(p7XV��;Y,%�й޼�x˅-�0z�*X*߇��+�������4�#��#���������]E��, 
��I�U���L��=�L쑼��v�is"���<�eη�{������fUýI���wtZ�*��f�0W֣��V�D�;1�c�=�/+��z�]���M��]���E*��b�L 5�:`'��s����@ה�,��G
�ѰB���ҵ��ި��N� ��ek��'h,Yv���M��2�r�� q�ro.��Wn�ˠ=�]�}��;7~g�
˝lJ
g���urT1�����ļA�fv�f1�x��*��9�wWpY�/I�vF�"Q�r��]<(#F�[�Αp�n\a��.�Ɓu�*I��C�!���o�C�ԣ��V;��}#39��O�#{�ֽ���Rv�ɢ�)�z�n3CX��V*Mr�����:�mL]n��=����K  �8֮�M�
G���1-4i4�ڷ�u��v��O�>'ev���q�xxBNHKU�y�
�ER�9Ørp�ʅ�>\θ^t�@E���+ �Qmn˅3��J3�u�GP�hkӎ��T�U���N�`��j�߽�Ѱ����G�\9�q�kPod�۱�6�\}��"� /�*\.NU�WW��x:Bwc�Z�z�#W��䧛�U�'��u
�v����+�ʓv��t�麏)fK�����iϾ�荳��m���^ڮ+3�<���*�=��Y&��U���HWe@k2T�>O(4�k_r��Rq{3�ZFD)ңґnf��7)�G��w5��6�ϡͼ�F���qd��m��r�p�����c-$����ZI���c��Lt����r��3-����+�!���"��ym�T�!k�D]�b�{�k�c��݋�0R����SBg9�A�)��&�klɰ���p-F�u{���.s��w`��wj�K+vRp[v勲;���Kg:���)[#H�tK���]�)˴���Ѫvy���H��[R�t3I��HE9�o%�r��U G�,��5�j�lb��$*)�eMOh0ot<��u͋�Y*({�u�u<��ڄ�yUn�	V$�T9�X%�\[+�;��v�{PGW���WZd�b��͋�/d����9o$�ep�,��%͝�JUsԘ�r��JÖ�����oah�Y�N^�!�Y�����	����\�����|gYN�j��J���ͦ\Ǯֲ��R��
#�\�E��!Z����S`ƅ��}\����cJ�M�O;��lGW;%�WQ�TOm��ԳJ��CKz� vpN��1��U���[�K9ä��Z]�82�P~kC�c���r�VMW=����Ug�I$�R܎�)����P�Z�q[J��]fY"pG�֚���sۉ��}|��E�ZB�8�I�B˙|,,ٷ�9ҽڢ�-�G����+����&R�x�S\��^M�s��b�6Z8kg�����Qѯn�<��jD���:Vfѱ��������x�=�&Ɔ*�%J��;\޾\^+KӄD��Κ�V5F�ǭ��[�T�,�l�uVTk�d=u�ܳ��	EKX
l#����ң�/��0�k�)����YN����84���խ��ZWf	�*�o�?x�Ű:hƄ��T9�[}V��u7Rr�w']�)RX�V3�U{w��i"��Sy���g��;mW1d�J"�!1&�n7m��:މW�ʧ��n'�Ŝ�0�\p�i�}���:4���U"���O�+�����_F(=52��u�N���Ӈ�ڸ@����X��k;�u�w+�(&B
(��¨�}�6�i�X�Үl]d��q(����dc�]��9��A�X��u��7��L����V�,�R�J:w�� �$<�O*��� ��~�Oz�M�=�/�����X�D�M����'3�:��qC*d�㵎wT���io�*�l�rE��:9�4*��Tx�\��I6\���Ae����ԺS�Ttr&'v�������ZVu3kQN�X.M�e�Nϥr]PL�t&�df1B��h���ͬT���ѽX3r��n	���ۘ�p�>��U�2^6�\(�k����=<�>���]+��lZw8��M���9D��ڢѥ,1�V��ݥ�b�eO4ʮ4���h��PЯ�Y)�G)�y���Nr�c{(��`���<8��ͺ���z���2ͣo8!*m�u����{�˓�h�T��.*li����6���ܵstk��Ie%ݝ3�j�j��*C����ƶ�ls�Bh��ǫHK�z�/^
�7�=9�dL2,]4����G^�]e�r%Ϩk)fo)����Ңf$n�i�nB���jƞX(���9�Y���U�L�fv޼ޜ��L`�-D� �0��;:����%��K�;P��8��Sa��dk��3�n��r`t�Ѧ��q��KT��$�;��N��;�Y�H�߆M�|��~ڢ *�����������?��r�������A'�T�~����v�e-�������5&<V�"v 2�2$n*�Cc��[���U��A����f��P��ʫ#p�Ȫ��	"��EU�����N�eԐAUeC�钩�	Qcm���R����
A���E�a��e�
�XVލ�g%ka�Wo-�ŕ���$E��]�B�oQD��Is@8�hM�G�\�Z��he����֜n66�VD
D2�j�b��:�Kz�+���z�vL��z�F(��s �k	�Lh�T��dLT !�d��B+*�j���P#*��0�HYF&�m����m<��d��Ĭ���V�l���6vJ��'�U�! u�-�R��Y1��mv���@Y3���O2�nL�O�\�������N�-����MTF�dэIX��h��bhi�I$L%��%,���Q�&Qd�`���c����eA�Uć����C��E#j*�q�)P�̳��p�P�.��B���=W�	2I�3�V�y}W&]�f�m�]�b��]6/�qgft=���\d��&�0@l*Eum.U�\Z�-ܾV��5��/�R6	�����S� �������קk��#7ws��j���`�r4���Β�zk��f�0�n¸����d٭�����D��	m+���;ep�5��<�L*�ۏ����ƪ�d��4���)<���Xv�ݤAJ�p;���ZL@q���˱����������yRX6IB��AAݹ&+�A
����x$��tfӃU9�Iޕ"�)u�)#Y]�D5�I�H�\�nB��p��n��RE�<pPT���8m.��O�&g[��ǲ�S%����u'u������<�p�I���nrY��Nڄ.X/q�Q>��^������5� ;l���V�bL���ETZ�7v�%���;�k[�QN�9��VZ�8A/�P%u�U蓓!�u����q?[[��ª�����3�yܬ�L�k#xuH��z{�3xҮ���*�d+[���6���:���+�Go(c�W��M�l+i�cu٩S��	�&Z�k-��-�"e�@r��n��G�2(��D(��el�&�*+(

�(�\��@Ԏ��"��	��[��iFf�j��\�_Y�ƈ4奩��#N��mK!X�
˧u�$i�Ȫ��nX��i������TǨ7T)+��j6A�VH�R&KX@���Td��	,�Ye��2�-+e���Q�;K����I�+��*�����]���d�¶�����m�_qb�����5�ۚ
����9$�ъ�(Id$�eգtC��J�*PZ��H$�
6[ko�a��	"wV�'�����E�J��6&���U��AW۔��ءI+e���7l�C�A�"qX;`1W5bl����%QKT��D�n��CT42�
�,rId�"B)I]C��ziס�G��fX+��)A��Ȅ�jWP;kn��(W-�+�ަZ� D��LPv���2����G!-T.��j��]n�H�R(dz�uB������`��m�q��EP�tJ�n4��B�;eӎ:�wD������=9$l$��Pժڝr���DQ��ٗ PX��r��q�Œ�P������|�N�k��sq�d򓃡���ˎ&�26��Jӌ"�#�st�o��~#I�Yk�F��d�(V6"H�r�ɤЫU��j�x���dQ��u���B�؞�M�Ҕ$��"��=KD�危�hQʭ�դvK"n�n�0�$����R��,b�j�ƀDN+j�U���(��q6�1[+����(����R)F���6'F9-r#B��ME)[R�R��!$M��V�A&�Q��[r��UYP₊�F(W,�% Yuh�rټ��dm�RTԅ�R�$n�G+m����kI��C��� �(��\����"�I�BI���v�t���_]u��뮺믮��뮸�8��{'�((��q�B\*%Dj%�I8����~g��󸲥JeD��э��n:뮺��u�]u�]}tu�]u�q�^��x��4$�LU!&R�Q��Nן89�ޘ�L�wn�oO�����:�u�]u�_]u�]q�q׷�ƟaP	簶2
��<ɥ�/���DtW76N�x���8;�G����aud��ʮ��N=:뮼|u�:뮺뮾�:뮺�8��¨O�u8.��"�;���n�Q]���x�D��Fs�.c���<���/L���O.�켆9�u�@e��8��m����\��\����p�屑;���5��QԻ�c�S�J�0J�"Mw`�GCs�9��m�I�����4D��~��<�:����l�iSI�vNN��dGV9�Z�{���S 
SD획�
���H�,n����I"8�^v�:{���7=���N�
pc��[�k��,Ft(d�o;�����S�y:�v�^�. �x�O~�_��ҔyT�FIyciZ��6�E�$�*j7�ZLOI[�r�t�-�	^w�xdE�8^�w����)G�b��s߯6�:�z^5H1���a�Bx�Vk��MOp�n%�V����Oi�~^z�����Q��r�ޮG�y/��u�r�y���T�w*C.N����q�ܬ�S

�п��������x����m�2(��uRJ�q��MJU,$R"���E��@�Ue��k���B�DT�ҩT���	a#UJ��A�IQ�"�=�?�9�u��2��6/� ��������Eo_Q�'.�O���o��s���[�cQ�����Ԏ(*�:�LR���N��֣q�E(��J�쳗2�$�N�]i�i`�7�r�ז�(����h�f5J�`�
�X䴠V�X��<ԒA�KJ�Ua%���;Gjp�R�X�u��u�:�,nH��FՎ�IP:���XK�F��8�)[*�;l���J������c�Z%�{פ���N�_k��n�$�]�A��*JĻ5�b�v�^��V���0�[�N3�p�;47+re6�S���qf:���*����|�n*]&x�޵f��O����э5������}Kk��q�LW�'��{�{x|���L�qt��7�ut`�55��x֠$�r��s-:b�M�ڬ�$�M�)�ϟ�@��fz)ĸ�3�C�*���sEY�XuN�V'eܵA����u��|��}�q$�e)���0��F�*1�6�fNMꔥ����om �)���@��e4�	�E�x�C��42��Kی@��Q�>�Y$���U��Xa��'hR�<���&OO
��'�o�~�3>�ڼ����U�U׶�P�GG�k`���}ݿ/w84�mS0c�����Rwή�(��Y�{��s����]v�H�|��Lܼ�bg'3��y^�x'��|r��z>��Fo�,b���967tT4-i�;�R��ð�{��� ��of��_���<��"��>q&���fV������GoΌ�j�'�N/y:�h#�5�+�ʫKݥ�������t��[�':�M�'��fu���'�e��c��->7�~ ���h���:Xa�Pj���x���0�{>��
p%�m�Vq>���*ww׶|*'�Y�B����TlD�0&�X�|��$��e}��)!R	!�0����x�u��*Yop/Q����������?p��œi���;.5����/�^�����2�����jG����X��p�@��)Fh͊�n�����C�7��(����Y�r��`��.�f��$&,���3�1�j��+0�xvg�ڻ���j��B��v�O/-�;�t�����>���T����O���=9哙�)�U��.�N}~k����|���$��Ei����晽%*AY�n�[:4�*�K&[vrŋ�:�V�����k(״�x�>�hfd��[>kg�on4a�S[�"P�mE,�WZے�������]�p۸�N�߫�?Cx(�߸J�j]���� 
����q�Y���R�ױ]�-uz�U~��������[|9b� � �T����RZ��e��� �����V�wv>v�ȉ��ʪ�UL�4��6<'��7��b�fB�
���[Z��v���"RfS�zQ[7%>H
�	����.J̖��o{utR�7��]�m3�+#�$�s�C�d=�>��6z��Kr��H�ﰯ�`�;`������
3`EU�Ndҷ��tۍ�֌�y����ު�#
�'�쑀���|�<{(����lkijDo�r�^����ߛ&A�c����-� �f�36����:���ts�hH~�U����/ۯ��详�G��k�I�bP��V ��!扰����=�ct��6��7*i�������R�yIPK�U��be���=;T[B�r%���7�^�z���wu��6-��R6����K_��&�R�u5ǰ��2��7�޽�<o<�:�+J�6���2�\k�TU-*;�{�P'�w�:f�� �����x(ν�����<�;�=���;�'�K����{���*c1�b���:vp��\O�,
�͝�v���{
�������îF�xM����S���U:͛��I�9��֔�;Y>G�oxM�:/lkp�WoFb&!��fh�Q��S�W�f=r�׹ f�QR�*e����
�j>��w�N��E�Y㬗�4��:��Sx�m� �XLø)��ii/��f��Am�[a�)��^�M�u�:���"�����ZiI��j����{<��P>��dNϩC��2 �ʻTKmWmT�U7�H;ΪO������"�@���mv'��fß["�5�ʛ����$�{��@��M�N��2���@�y��0�aTqW����D��%B��[�;�d�e��o��P�d�xv�j��$��h��*�J+Q���L�ܟfz���y��X�g�,=f�P3�qԑ��s��[��(#��>w�Jsz�k�DZyq��ʰc*+�b��^F��|XA'RW*��]��w�P�vv9!��vE|˦/8��و}����սUn�]��d��������"�=Nl�*Ϫ�����Pڦ2.Á���,���J^�~�Ǖ��L�g������-U�'7��(��.��IⰝ$!��Ꝫ��Ʈ�ͤ�#��?y��A3Ù@\�C���+��x���> Q�h�	`zӪ����T�)�9�V_�<�p�4]{�?�N}���5o-�B"}��*���ݕ���捁u}��\'s�-)78��Թ�j���E���$d�t��7�nS�C85�	;C��8j�,����"���S�	��0��ԣ���ׯ<++�̚�.��+_��l+��[�s&��"��y����@5��]��]d}�}tK��^��}'�}��(9k���EHrQ&�V
�oV��S*a��Z'Y�����M2�4���#s�s��oP��1�zK�L)���Rz�Ạ��f����Oz	���6�Q�V�$,��OB�mR�JŅn,�h���p���l���
}&����meܫ�<����ӷ��v�Q�s��z�=���J�}Co�A۲��&m���q i��C�G�G֐G���#ʗ�!�7_���@]��|q��b�	��z�s��w��	���e�Q�|&����{C@�<||�y����$ʓ^�^�Tp�+$��g
g��*N�W�s̝j�c�ح�)R��Q����([Y�:��z�%�*={>4,�h�3U�V��V��%Y2����W�;�#�5[��1	�դ�s��1S�鏔w����»�l����7@���#/6V
2�(a�-rZ+e��1�Tj�J����srv��΍-A���"#̮dR0���4�����k��������gCl-�<*/��6�B�S�Ij��Ϳ�[�8>�;nu ʜ��^k9|�/�^��	$�zzR>�;�K�.�˭S�����x5�m���ʟ�;:Q4�EDPS�".Q��A�T���C�fɑ�W�a=���J�'76�{(õ���-X]�
U]�1���|�k�u�*�{�cA���Z���^�f��;�.�Z�a�M�Vd�Χwµ�O��Wk~���M�E4=E  �_r�zK��m��=�V�d�NU��r{#]\]הD�Q<;��]K}KG�����o~�u�Fk�1#1B�޹}�lG��τ��L�������AU���(�a�cŧ�q�6��  �ܬ�Z��(�G��������բO�͌�t5�ID�\��±�g
����;�R7A�`Cw7hY2h�YN5]��{r��q6��+p&wZ����Dˠ�_�y2����>����� �h�ҵf%��N]�r�Qp�,�!׈�&Ѯy���S�ߔ�>���0�����H������E���$��)NY����*̨�R��EȒf��N]�tǢ�L�P�A�"���}~�;��a�qn�a99�{�(��-�^o"���+r-AN�]eÜ�R�Z�:l.��mx����N�R�2[&�W�o5���^j��E�Рnʰ/զ1��ɜ�/�<��us\��F�/��7h�d8����w�8Ճ�6��^��Ț���?uX7�SZ�ȡ[���wX�}U�Ͼ�@��_��]V������M9��!V�T8<���N�tA8�v�h�5^.Yr1ق�7�Ar،��*tC�`F1�f�~o���k���b��+z���-��~�6���n#�qk��.�R��ޔ�8"�ro�4���'�K�zR�ߺ�W�|��(�~���Iu�ߎ�ozY�zO,���9'�������j�z�4�a�$f(�d��>��}
��}�
Fs�U�~1T�NSQ$%��u�b�<i�fN�ܳl��ў�kV�-W��ub; �M�����9owl������+�p��ge,eP���했fv����ZЉ� cui��T�k)e�vu�[�;�FjEm�hf��,��* 1|��b��'l	���/)�J&}y᳨5SǱ�ct�Ÿ[�L��)�k���9E�e:m�}Cej2r&Hiq����9u�����bZ
pS�ݻ�֯gS��d݇j�qA��v�d��#ۢ�N���}�������<������G�e+_����U����{�}��oc"��7��LX�t��P���������u9�m�\H=��Q���`��w$��y�^Okv��R�^���겏U� <�ĳc]��p1��B��6�=�Qy;��>8�D�l^p�r���6�Q�����w+���0]�s(�M�)U_{�����wda5�J��M�Co�<��.��U�}W��J/����ՋO�<�Ŧ��4�����[�<����x�S��&��٩huR"�
�k����s'b=[�7[Z�!�nC6o� ;QgJ>@�B�����#�|~��Ͻ�9������u�����s&�zʼ�3EU̓���&�C�C]d�*(T������U����jĬ�����>���:�������^��|��\�9�ΐ�#v��H1�sE׬4���D���@r���$��� ���#<�Zf�����N�ñE���Un۬������<�<�����A	�e6�u*�`Mz�^9`�8���oj�X�=��UPVj6���mS0I��R+�ޢ'�J=�wM�ِ]R���`ʲbP� ��
�0�\Z�7v3���X[Y�&:���:�l�S�5�9�ˈ�,�Vh]J=W. �Wؒ��ՠ�b�WLg�����+��d�2ӷ��wf���V�S��x�||�����g7�ϰm\�k������g��||��ǝD��xo}b4��Z�X��'�O������6� �4�{���*��R�f�w��C��n�u!q�o���Q��Pl�Ԉ�u���w���ȉk�Ѳ�Հ�^�Z�su�V�~�^�Ѿi�&}�Z�N��voeLb�ف;���g�~��	�Sa�E��|�|�wE;�"%Iw����~�ޮ�_�Y�S��S��o�|�y"d,֭��~���{�E-��0�at����p9˘����S�#"��I�����J�:pš��Hl��*4%{��l��Y�M�;����­���E�.=C��򱾊"��ݯ`��M��<�»����6�3���&�Hh����0s�21�x>�����#�4��5�&����3��u}�L��DsNXZ�@��LZ�7�`;[�D�,�칻]83�	r�Yّ������	��)�a%��T[dV*��B�U�q���^:z��Hsv�����v��YV2�ḍ�S�Cf'Bo9R�&p�Dw���Ы9(��T�fU6��Ӂ�뽆��<Pq�m!�S;��eps%���h�{F��/��%���gXg�Z#>�(R�A�;����Lt���H�[R��M;�7O�H�U[k3���B���$�h�Gn�O��W�T̆q/����Q��R�����0�Ūo�2$8�J={��{�ͽ:\deR�g��t5��2��N`�����;t�U��k.�f�1"]�A�e���7U�t��n�e�*5Zi��Q軩v���J&1�+�Djܽ�\SI�ܼ�pL���V��ͭ��t���]p^�vml*��޻:�sc���Zk5�N��]�_w+��-�0���ӳ��W���f�ǝV0u�I���GW�d{�� �}�v���Xi�֘޻���wo.N�hlfuH��^��ul�����F�JI�
�,x���n=�����=b�H��KN�FN�Q�2�:>y�^�j�v:��MĤC��X��^zNѶΠ���[���np8����������!�|�2.�X4D����	�,SD7Aʀ�>��=ƍ�����.u%y�X�M�a,��B��a�)�M���S/,�z�WVN"b���/C��ӽ֩6�nQ�6�5�q-�sFw%UZ.�q�4��Gz��� Ҝ�=ʢyZ��~ޮKZ�����
i�v��4���uv����X�;�9��V����gK!g`<�\��+&�xz��4��v�ξ�y|�t���0�{��#]�49�T5���� ���\��K�%Y��o�Wz�s�!Y
�Q�P�ۂ�C;]ƥ)T��R�>ڡ��w�7�t��V��peʆ��@��Z
$d���(r�뵡d:p=�*5�#�w�Z�-�`�O������)�+(��Wׄ��f�2Q�콧ѻ�=[K�C6:����k��Gn�O�<;u�Y/�'Rӧ1.]�hRA�}yW����Eu�(��Tj-��^�w�ml��x
���*V�U�;���
]E���YpJ�#Rp�Idv-LȲ�5�$��R�I�<�3�euQ�S��y��n�h�y1��n8N���f8�Z��Ԭz�_wej�ս�lIJ�[ʚ�1�޼ͽ�1��>_Ɵ�=4�I�B3O�v��w�	!�P^|)�������H6�4	I���P�"m��2�C���mǧ]x����Ǎ<u�]u��G]u��m�^1�]��"m6�2I�q�غ�4لzm�S7�r�2M�d?%�l7ksm�=������Ǐx���]u���]u��m׃߄<'*�c
��$��L~yN�ܨ���"�Ȼ�W��X�U�(��ֵ�v�����x��Ǐ4��Ǐ:��뮺�m��o��=��|�����v�!#Zz�Z�j�G4�̒5�%�cۊ*TdIB�U\�q�_^<{u׏x��Ǐ><u�[m��x��>"��/ع�S�e9���+��K��(�DՑ*��$�PQ.�~�r<�@褉kQL"�[�Zp��uH��P���?k�`R*IU&#��'NH}�:/��;�U
��
���/ZWL��q��K���)�t�CE�[C�\�EЂ*��b�wJ��q��Я�y����} =px+��H��XHY��$"�~�x��D�|�9?wv��.��%����T�-�4(h���e����o7;�R��3 �.���m̾� s:��1��{�����w��w�]�oL��44�(g���/z���H =ED]��UU_���V���&�qM������f���&�T+�
��CY�j{��6���
�O��� ��%�����vLܮܑ���b��+?Wx��D�Xܮ;e�-�|�^���׽�3���t|(�r�}�$k���Z�w�,���>O{�nY�o��9������x&]}v�j��:��(�7���������_�,ʮ�(z�w��Q�`+̍���tO���xdt7��Vv/��Uo���g�a��0J�1��u��^8�>���e�)�<���8�hq����fo �7���$�$�T�� ��v����tqS`y�'�|�uư��y�e*��� Z��}/N��P��1�C�{9�����~E?"_��~C�(:g��Su������Y��[�T{�ڻ����nD��l���b�ݴIkR��u�����.y�7S�xt�Q�8����i�rLdW.�{Q�.f�NWfu�y���{���U�-���ZϷ<�W������=.�'�w�l�2מ| �y��;��[e�nr��ʨ�'��� ;����E0���b�����!yð�p/]���?k�>�~�>V���^
�r"q+�F�-��(����iE*;�/�N�^�v�-��{kr�[�-�+V�C�O� T��<�9�Uݷ��ڧ]�+y[��e�U�w�uu7W8-�c�u����%�V��Nx��(cLQ��3�3f��K��Ϝkm��y�&w��w���z3�����I0�W�C��Rm�������;�����Y�nO�Ű���(cB��R��	���G���_o٤[v�3� �(�Y�[2���.�!M�}���׫ۿ&�ם�����4{\6�K�J-*9�#������M�E���~J���69�y�����!�������&���A����U_�_���ԓ��@C�NPl����*�{=�bSO��de'��ޟt�w�4%���/3���\��5][=���{�����7���<�[���Ϗ~/�O�S����7��Ӓ�5U��<:����_� ��������q�״�?+���y�]�[3}<���o�V@��V�SC<@�����KvCg����W���y��mm�}�4O�0;6)��>ǆ����qH?��J��{`�3}=2�ݽ�-�^n������N}�����`u�]4�@=���n�==�ط��jR�^���j��j��e7�i}���<���BA�ߩ?.����k'����\���="�����J�9�<�slQp���M�W}k�ޗ[/f��p��ܲ,E���n��ǚ�9Z�s=�Hy����[��S�1�C`�/ ��@�#馽�ԉ�������+�����d��x�o�n�A]IS���XT����ZI�w~�/���:�Y������i�1�'���b�_�[�e�lmH~�VK��/u�{�i컷�+�ݧq��˲ܑ�b;�ɤ�������o�W�Vo���U2�LӘo��#C�F.U���P,�ˏ�<�@����W�aOs�YW�ԧ�^*ͭ(/�;�=���n�d�o9��ʟ@��7��wMs�6��[���� x3z�����%��
2>O��oGU۹�vI�up���s�6!_=�U�2�:ƻ}��%�C�	�IiV�V��6g��< �1m�b����>�SK�E\��]���i�N��!,ps��!�L�/���g;�����q|�J%�Ew�������wW�P_�p��w��q�Ǎ{����9��h�W�&�� �������	�>`7�Y%8���,&�ؤ�[�B{mi��1�19d&��n�r#���\��c��^lnon?��x����)�[�gG��x��c�������R���i!y0	����`~h>'D>y߲�M\�E;	��OLkv�u����Uw#�.
��g�iO��T@d����C�}z޼�����X�����wҘ\���%��u����x [X
�l3�ϠpDx)0)�c˸�@��*��m�d6���8��ء�>B{���ź=J˳����n���L�����C1��l�o�!۪�Zw˴h����
??F��5E@��y纲V���ރ�J��a�q'����ˡӞ����Evӭܘ�#O7x�D��<}�(cM4��&���=�pd�ܯ�����P�^�@]��V}�C<�!s0��>����Rm>;��
��Kx�iz �{5趼�@��p!�c���H8��uy����������2��DC�cTB��=��,)͊w"��*^��!x����PN;���/���|}�W�0z�b���^c���+� [����,I���M���֕���~6�OӸ2|�D	peTx��Ig`���3w0�g.�7r+��7��~�U�50fC\	lN%�b<�:}�Ml��m�RJaڪw�/y�{�ֲ���0s�\��O�q�������%� ]��g�_~8�X�sY�y��a���ڻ��Y*��S/��y1Ww���|Á��@M�cZ��� Su.���1~��9q}_�B��a�a?&\�י���� k�q��Q������Z�-���\o��[�k��6�5ѧk]��n�c-f���c�p{�>lel���%��+��{�m�mj	F��E�q@tO��a-��1����s�w�{���yt���\���5�p���Tt���cj�q�jp1�����[��������?����N�-�Yh�5�Q���:�����ْ�KǙ$������v�L��E�d�Y ��66u��Ó0���AW2dYկ�wG9kj��W8%|��Z7���{�[S�_�_;�^����?��1�hֳ�~���l������U{T�-I��2,�Y([efY�����s���-��= �dޑ��b6�d����սz���s�q�y��/ w~_�Y�[��;����0$ =�_�4#��@�GCq;��ڙ��ʜ�'�����<Ǽ���k�v�nǐ=�e�����{�e_*B�~�� ��-I�Sm����C�̬uYZ�{ə�������l�`+ق4Mz<_������w�����d�v�.�f�{�{�{�_�RJ��!����}f��{u��5��������耛Ļg���{u��� s/-�[��y7���0˜H�~?x�����cQ��pa:�Y�%�3�z⯴�mq�~�\����ܢWe�0&W!�y	�G:ُC@� SO_��C�oE����tr�V����n��b��Z��슍Un=u!��T7ݹ�W���o����A`�����;םX{�=�M�x�fy���&��^�	�XW��k��*�Ԍ]>F�kw6�=+�_�Ç��;V�=�}������=N?�m�c�L���Ԝ��f�5��[�z�G�G.��h�{�_R��#t��3l3{������|�6����1Cc�޾2�(�}nV��7?Gmz��*��ا��^GY��hKy�A#���Tz�� L��K�d;��;(�*�`���G��~�_�l����%u�Ƕ��hi����g��	�����{ɲ\\:a�8 �zh�k�34&��M���O��˺y���W�yld?\�j���u��^)�כ��0���,�
���/��
����.�=!�N�MI��\@���{9��5��Ȕ)�NUU���5i�ީd�r�S���0�/9�5<��,�W�n�^y�/����ɚ�����)�-��sH��ha �k�4Sx@����|3���kqM�}=�����p�������n��X�S�y&��xq��zs_�԰�8ƶ����}΢<=�ڴ��XL���Ї������Ul.
��t���5�ln��&�!^v����Zr�+7���W��R�g���Nv�|��������O58�����~�[����$�F7v�!�w�v^��7���&�"m�R鵤vNҁ�q���a�����S�8�ɀ-n/t��sGx��"<�����g�-����P��[}����<:�}5���D��vd�K���K�++)�<5?�#n��,}���kUqnu�g���=�+n$]�x"{����?=D���ܭ����|��n�z/a�ը���1���2�]2Ӱ��8xzTB�T�u�
���>�Ҍ8�=fո��[�Vm`������9�(EǇ�V>����ybWiucv��a����`�>~>C���4��	�W�����k3޹������lbtԛ۰-}}ć�ܑ�eɛD5����u��ƺ�{�a���-u��։�@�vkK"�t��R&�PUU�N�6�'��r�����pƪ�ux6>�W����
k͐@�E��t�ȸ��<�Cq~��}ah��kJ�>7�l����Z����ѽ�#:�t�<�!폛��Y SSsKg��w�sh{����[h):]��w��� ;_�R��J����>������Fe�P]��a�y^�U��Y�l�	>��_0�+�hJ��My���p�gV��KV$�5N"b&����%�%�"r�@�3����qL�n�O�[�5:�ʆ��ۣ�����;W���̛ПW��޾^�5��	q�|��+k�����Ö�O���v��1Y�s7�c4����	OZpr���z(�:�e���lz{�Z�=#�|�]N��$$P�b��y�����M��v�{\	�:/b��t��ʱ= ����ޘ��qμ�[�E��q=SR�(<�^�����g�q2����஽s͍"�k��Ps��^���u;	�ކ}���v�p[�1]��Į3k�\�a��Cף���~��f�k������fh��iV0�������(������-��cm���q����[�g�ltqJ7i�c*r�Ҷ�<j=��Z(p�w��)�{���
��ȹ��^&'Xwq��-�9�J���׺d�zq��}+�ZT'�5(���N���g���Oa/�0��44�
<�7���Q)�n�`.�?�k�W9��f6�9��hΎ�_u��
�<wFqB索'6�!�{��j�G�� ǻ�g�	A�<̰���RѶ2l�iw���a#�0����v��s�>*�ER���>��cZ���5�s�99��z��#�|�t�������(�f��z�2�Ǯ�j{3N����&v�!�K�&�K�aB��EC�/�A���v�-���-����:������B2���~Ρ���$
��� /���^��f~#�Ri���K=��t�@y�q>��E�0�f���[?3�ڟ0Ǘ�� N���ν"H������꯸�`���S���*P�_r���g���p��>���ݖ{ĦX��Y�������﷩|�>7��=;��W�I�����[W��x�s���~�i���:��Z��5u|��վ����ex"�o����[}w��0�9�5dG�)3�n�3M�4��1ƫԸ3<�j��xd��I��u�6�:�7zO�q����Z'��İ%Bޜ�ڟ!���oo���U��n�~���Z�˲����{$��.������y��W�_9�+2�S�̕��{>��?;�n�}l/����ܞ�����Nh�CB$�r�u�}�9��wr9*�ow�[G�G��� �:�nw���rO���CaCF��l
�1���u����}���s��2�31���C�`y��)����;ʹ7��aNc�n+�2b޽����g[rK���[+'�<�S//8�K� ��g@�r�^��~o.���i�� �*��+tPw�f���6"^*��YY���y57��]Sæ���9-���Zd<;��=�}j�Qᵉ��<3sd؍�q۷X�JɁn;r�l80� ��=� ��:`${͍���'np�-�����3��>5I�oB��ˮ+��fiUUO�ګ��v0�����}�a�B���<�9}�,�O~��HI��Y_���|���{�ټÀ��ϵ����Oa_zD�����{a��sx����:iُ�x��O��G�A�À�^�L�`[{��N��� ���}l1���~a�?W���+���臶��v��7ץ���oޗb�l�r_y��
BIH�� ��������s;W����=��l`��.�&�k��n�=��kg６P���Hދts�[<0�e�0�t��G"2*�q@x�iǖ}�aИ4�n�L�hoSr̟=J��L3���v�e�B��f����<x��Щ�҃+l=���t��\dk�Z2���'\��ۍ/S���^X��T�iME�\��:�vml��ܓ��b�c�gr��Z�X��wdOw4�$C�<���� 䯡��>�M��˒��ڲ[�E�bB��B2BC|�o���|�ޟ�A)���WɎ�q�\����_��z��su\���ğ@�zZԜ���*���+����TSxw0{&��s��\/������{��^��'�,�P�ڌa���N�D�@����I����Ck��vE�9�~T�0�c���7��=ZR�#�@������7w5J��s"�3s� <�^?�����4c�^q#��>tAc�w��-�~N����>��w�j�h��n��ypX�&k�8�p1��b�!��>���[-�:��=Ҹ�����33H��K�0H�1\m����C�7�_)Qc�����y>j��k��p��3H�t�/ln(1�j�ag�e�+��Yt�#�zkh2O3P���~o��%������xW���ɓ��
��3��Ɔ/=#�[�֔��'��<�b�����L�3tP'�U��`�E0�l1,�&�Pb�lT3s:j�;[�ˀ��� ��&搔k�c�bJ���&�cQ/�.��ߎ��,�۝�h�Ȟǵ���	�1>�*�,����y��\�?�K��6)Ϡk ��>�}�C� ��}�e�����J�����$�V���.��u�X2�G�-�}�i�齂��Ϫ���6"�,�^k��l��Ⱥ�7�_��4�,�p'��u�uk�'B��3�|���.=eS��eK�u�	^�����DmM"�;j��^��a�})����/kz�͕~Ɉ�E���]�(�"q�\��/ABf-\��St7:�rn���q��N���8�j���cu8��bs;,;���h�]H�-���}�!%B��Sy9�7��T��{Ӿ��M�(�J�)Y����E��ـ���Ft�݂ۦ&��w��p��uU�tF�.���A}#��IAt�����l�.�C���(�d˂;��Z�O���`R�Vf��۝*�`٦yՉK6������ҭX��sg��3y̱2��R4���fumˊ�g]�E�ii�3F��\��F�;�������w�Ɣ�WRb�6�лtm[�D|&q���A�GK[��@�`5gN�˷y�(�I�u����ζ�N�P�����1�R�&1�/� n:�|૥gi�
�"�<�ՔF��#:M^U���V��ؤUU�ZR�4��L�V����酈!H��Ƴ��ub�.t/	��fUC��R���)u�2U�8+��,�ꩂ�����dGCm)UTE�%U�6g���W/��sd���:� ���NۤY�>��PS����7z�eI�%f�%�&�	/�6f`��]��udO�-��h�;z�r�H�1�WNL���Xߎv�$�����ѐ��\F��J���%qʈC��$�Xy���e�e��x #+�*^H�Od��-?��.�����VVXN]��h�k,pJ��V�]eśfWP#V'����R\��1˥��
�L�X��"��/�e��S��v���)��ͩ.K��s��Æ�_4�*��|���V�M��}x򫙼�qq�dy�e��w�Kd�m���J�&�N��c�ad�tub�˛-�h�RZ�Z�Ґ��+�~�/F���?Z�j�'pw���bA��Jœ��5�U£.e��l�Z���4���	65:�}�r)�2z	c�)ol^̲��k�(p���1��u�+Q�� �:�U���ݬtE��N�]�5�hb�E>�`��K����a��f���%��Mt��3�jG����/1K��-�\m��wLgG��\����{tv����`�����$|_���/��mpV-̲��@��u�������g<�
l����;��z�zK���](��
B�IT�M6�ۯ�u��]u�^<x���ǃǏm��u���<fUޔ]����ds�v��ǑDy$��Yj�_�"o���z�oϏ�zu�]m�]u�Ǐ��<m�۷����]򙂘�aVc&B�QE�Yj�����^m��:�OOn=���^�u�[u�]u׷��<m��x���gt�<�/�:��JS@���ޭ>y�:]M�\�J*��ܬ4Bwl:cN8㮺����]u�]u�]{u�<x���m�����4r��j�N��BARN�Q(\MH#ChQ2}�n�w�&v'"�֜��H�(hJˬ�.��~�p��+��ʪ{���fA��+�{��J�,DS�*N��TE:�+��Z+�{����.(YÑr�Q"��Ĳ�Y�����(�D+��kǮ��(��d$����4���2Η��R�C��s ��(��Q�����@��$Y��/G<�l�4�ZX����*s	���r)a��3�d��m��|��s̕"�R��H�O�}m�Xi	�5��Ik�� �d�!#��卫����I.��8㪍�����Piƣ�v�`�"���,Эn�["#�+-�(;#�B�ed��Ss�{�羷z\{xsE��m�Hw��YL�����J��<n����F�'>�ţ�����oDRm�Y�-�)��r6+$��YT��ƅ��r[$��e�����Bt�����]�h��U$)U���l�+��Ek���u@��!-U�QM1��V
"Pv�8� R"TW����W�TQ`������OE��9-hSBamW
�(�U]T�&M�B&�M�R�B���r�L���:�%�i��d ���kd@���j�AIC7����9��C�`��uF�L���:~V���˻�c�/\�8^C�r�Ȓʚ�ΏF44�K@\�^tȳ&/k2��h�G'�]���Ua��;[����vz�Eu�a�[z�ܟu�l��5���u�sz�|WE�o>�$��xʾ�_�ʞ�%I�y���߹�ͺ��L&#$.�	V�Ux�"۪��Q\��`��M�A�:נ?<3��b&V �sz}N�k�D��B�M�SR{������l@���o1���K~F�Ÿ�]�~��cK:��x�:>V���+;��W�t��i��a57uy������K
��}��3Z�F0ƶ�4nd�n��|�|#X@w��&ͦ.��vy+�$�����=�M��d��_Aa#z��������ش;�@�nS]�1�r��ز�w9�ϓ��i��,�H~��5�����v�2r��(��J�Qϧ}�f>{�I=�y/?��7�s��oc
��魀MMm��@`)��<^}�5A�s����RQ�\��-E=<�ԻSDKPs[o�Ǩ���6qk_��+�����S�j� [�uf�[����ٝV��=�#����)�-�1��{�m��C�W���:_��������Z��1�/�Sο6������뒬t�m�;f�b �R��,U�W��Ӻ�^u(���@%f�TM$ �^����zfV!����u���1�c=��f�6������1�hj�8��YT�gc]
�m��8�=����6 Slm�n)"6�m[���Lm�������Y�}�}�z��s���E�o�9��>Lߌ�{�f<0�����!��}40Xu;GS�^�u�(�pQ�|��6k�v������}W�u�xK��H�E���ޛ��T���$���܇y�g��S-��spV\�xSr��\�{J L��
�v�;�{yK9�:�e.dT_oj�<��}E�V���D�~���:7;��R+u���K-����zB�7�Z���5���'�<�E�G�~p<0f�p9�|���(���@������4z��W����8�4���i��_}�u�p���� koy�_��t�ϛ��y������q������(�}����؉���\��3�<E`��c/��:V��������޽�eK��*�X}*��ۨf\�\v�?gFguln�ř����Z:j�\�}���ݿ&m�n;ӄ�����tڂ�M��m��=�p$E�G�\@���HB&Q�E<{^��]��ޖ���@f�h(�^�����G��v��Ϲz@R�Ox�Q�=^�u��,c�I�����ō���=���&~,������}��u�	��������+)�4&͊V�R���T�ݧ�cOa�{�ޟU ��}�@mUmyA�B��Ǐp�P�	����#��8�34�y\:�+[ftz%>�q�K�ݘ)v���V���fZ8A�	���i�6�M���m��H�d	I dA��$T	,���3��>�=fg{w�t&����&W�i���������.���U���Ҽ��
����T�.�O�g/Q�=��S�ýw��1��L��l��:�`0s�w\�}x�!��5�*
��
�g�ͬ����HR~0Sw�@]�>�Y�����Rq,��qɮ3�2�Pյ �|��=�{[��G�]�`ө���70���fq�^�� cD<�{^���ɻ��Yn�v =b�;��<gPhx�x��[�l�Q�`3��m�Kj���8������\/,,������|�UUq�������28!n/�F0�|���P4{���5ozx��Ȧ� ��S��2h���C(������ñh`:�@o49�moD��d��ԁ��l�'9��46��kѭۆ��Q�5�9f��8����Pd��<k��������zڃ�SףK����_G�5����FNkOC:��8�p��Z��B���ړ��@�~�����F��k�a�{��Ј^�޿L�KP�6���J��ۊNi�#���a�߫K��Ah�=���Wk�rF0�gP��)�p���S�N��_r���|m���p�m@Gi�!~��p�E:�.�G�ݍ7�Ͱ�0���P@�K��j��vj��� �u˾J}(k{J�k��-����䛨6rZ�i�[�}F����u�T�y�״ftU~*����b�6��Qi�6ڋM����"� 2 TK"�.��>���^X�6K=��#��k6����s�Lnx 1�}<(�J�x!0|��"�٪��;��x���w�{�t_�<�՟`��˩�df/g���>��X���<ӻ�/v&��(�<�X41,�������aAW9j���}��0s�E��n�$���Ԁ���۾��=�k��y5�z��w�����-κ��������y>qRW���X��}v�&�gGuEF���ߦ�"�7+s�jqQoH��c 4�q}��p��y�=oM�hW364k��3۝8��9�6m�)�b\ �b�@�~xTd[�<����DTzj]��L[��۪�ǀ��Q-��X	�'�8*<;�Y2D��S�.�ù퀖�x��p�Ç@�O�w�ͯ&��=�y��:�E��AX��U@~����_�/��=+W���yq�l�uN�i��a\�y����@�ㆵ�@|ED8S��>_:{����f�u���kj��'6w�UoV��c��8���ǜ0��O���� ��ò�y�g��z8	�WA��;i�-�<�ZX�p�V���g1�4ۍs�(�(b��sU_d����oK�O��Wm�w{�N���$���m�A�,��nS�P��_��mF\�>��Vi�2�����dwq�q�G�v����D7�9��w��[ߵ}uߗ*���zc�h�Dm�6؋M���Jm���Y ��U$@	���ξ�'��צwէX��IK,OJ�c���3xr��Ὕ]�q`�o�ï�`Ө���P�V"������w�8m�ܮ������JG@��v�*~A��ޫ�O+��h�8��8k��??���r��^��1m��]�Jֽk�٬���p���֍���g1�͋�<5lK\O�e��0����Cz��C�����Mj��28z`5(����sh	W�u�3�&w}kgo���`��Gl\���=��js��MF�?��|��RǨL~����x88�u������<���k�xV"���EN����S�;�ư�����=���c٪Euy�Xa�����zLw�X�=	$c'��j4��_]7�rr����y���%�.���f����sO��L;7���W�[�:��֖�2.2b�Y����WS{���n���^��368���7ܹ��������9>��ky�黍�x�
)`�K��>v��4�2i�AP�D�%锌�
w�ޑ��X	1��!鯝98XĞ��o]�p���i���f��]��Y1���ax��P�����1`����-�^7FHN�Dg�E�Q�:y��Ӹ�&����zk=�˟�G
�� ��3�ϫ_�鄓<?_����(YF� һ�J���~���/93��V�>�n�Jk7%H�Wr!�AΜ���X�We��)��_�����o;�K{�vSᩖmՊt���5߸i=o�u�`K1��2	�@�r�C},��-�yG��ѻ�4�����6ةM���K��Lm�R�cm��$FD@� $���*�tWH�<�q���|��Kܽ0�C�r�ߏ���gA�׆x�Ѧ{:y�?���_z�7�}�\���8����A=AK�?�>ߵ��7�p'2�j�+D��y��[��t�=��f�ʕN�������6U�b ,�촑3��"�~���������[v�h>�ݖ�駎����P,��ݐxB��𻍼k����z���*6������������u1}��ȅy1���#��a��������Q�M�e�H�`b��;�{k�E�%���k%q̳��
,<��#�Ϭ�hKli�|6�3e����ڼ��i��Mf�n�:�@z堦�ihg�L/XU�}��ɀH����ҘS ��#Q��:�t���x��§�A�N^���FWn����`�A|v+��8����e��8�]/�vΰ�Om��^	F��Cq�KJ=���y�� <���{��nbʘW�z4�<��0d���y��O��S��������U���,?��^�o��Pk=�P!u ����!���;7]Ao�F�ƛ���q�Ҷ��A$�i�9g�����N�f�>��P�oU���Ȩ1�%g,qeJ}�E�N��k���	'b�ٶ�S�$������S�\�sӽ}���'�	�l~l@���j7�-�6؉M����H*�RH��w�w�y����k�U*W�N�R��8�(��AQ�'�A�y�φ���`;�9����c%���_��j��n��L$c��̹0�J7�!G�/37�	am�8((��V/��w-\�`2���0�l*,	�<7��̵�&@�f<��w�}~0u��纑$>��Z\�&�f!��������� Ah'=_�3=��o���4y����嵝'�k͖	����������zcX	g����8?7�=T�{2��7��s�߭���K����uЄ���P�]�ڮ<v*����X���Q7�x��]y��*6xQ����񫈆-L�����8�S��"�Fn�3�p�#�#͌���<J��>���3^�ᦜ3 ��M#�K[��;+S���O��ֶ��x @�I�G��LD.oO�W���{g���	��K���%�c{+��z�,׆���U���_Th��Q��W���?�����M��C��aa�;��u���݊��[ȡ��j<�
�w��7�C�����34�~o ��T!�_��{��T�.�����O|��͉�ԅ$([�š܅ba�c��Ǻ����;��ӧ,�ڍY�K2������J�5b��\�RBJވ�J�9/
{�3��Jٛ��ne��7x�l���O�]w�^�}�Y]{�_��ͱ��B⥴��
m���B�cm��c��u%�\pI���S��;�3kS �hR�o���09�{U]q���/��7%�^��d���<S�^�N�'�E��u�#Kn}�ƍoO�����^v�<'�;]h�c8l�/p�m!ݦ^$CĿ��?zcrr.@�&��7��Ӎ�oss��[:A/c�竣���;eŁmu�04�_1�?�"}>9՟
�@���>7p��4�l[���Op[�yyga���������>&�/�����7�����rK�m"o`:Wq=v9f���y0n� Nע�K=)��0���[Q���m�c35zډ��ߛ|��0%���h�_j�.�(p��w!^����p5����Az/~黨�x6�M��0	=�� ��l��|�������f��0�k�m���z2�}��s)���2|+�*c���{L�w���.qp/� ��PoN�3?�=�	�c�v�榱���0�� ]{aK��se�MLTfE��Ġ<�lW>~� ���0MXc�^�',3ߑ4-�08��s�c+�)��o!_U�+�A�ssn�a�����HK�p��a�z�M0�y�2�4g$z�K�/k��:�+���^>ۼ��o)û�'�];��7���}���7���� ��Lm�R�cm�\D-�6ح�i��pFEDU ��w����I\������6T���T�un�'m9�z%k�`&�w}
DeS����/�[����x�F�W�i$���>�_�Ξ��XE��<��U� 7��< 	�WhRԵ_(\i�[��`��M����<7�l_�d��9�m�`c����b�,`��վPu������_�n���gn�zwP#��]	�Jh�M�"��-����ٮ����E�#e��k���t���J�V���������ϭ��N��$��x)�������!o�i�7���.��3Çh�M���P�]A*-�[^���[��>9m���e���P����&�P�\�f�Ô�q~`3�틚�N�&���9��ѱͬ���ent�g����!�s��R�#%�eG?� ��y9��-��myO����n͡(���\� ���趆��mmC�[�Od�(��Z=Om���&=�2/h�^�\�Ed�Յs�N2��y�� N���2�s{���eK%N�y��
��lKҊ�_r� �:�U�J��X|0�������G��\N�D��˝=�Z��0CߵD���2k���ԡ��h�D�7F�\w?��>�`�"]uS]B�Z
sf�YǂW�5�t�1�����pm�Vhci]�{n�A���]U[n{��"U�� Q��"��]�?q���}�h���Vaw�eeI�o<�|v�|�S�E2oWQ�Eo	Ƒ��.�N�*8n��g}_�ࡐ_�cm�4�mD)�6ڂSlm�. � ! ���V]<�Q`��Q���/������^�rF����ʻ��=��NO��@|~Cf�;d�N���&r���#Ė;�݁��C�e��/`��S����N��cqiqM-z���kYy/�mF��Nt޹���&���^4s���-�_�8~����;���H���jd���K35P���ƀ]k�O����o��|�
F�T`�1�XZ�^O+3�#���d�|&��ϨLn���Y�T�@N54�}���Kg��l���[�gx�'���8�T>Q�g��:��\��g��@���g���k��7[Ǖ�;�yiw8���ҍ͵�.���|/�o볬��(0���L���W3ۗ���-�<nsMt�,|L ��mB����l�	צ�ŷ��h���D8�q�+��2��^)~_܏���o���{?6���n(Ȯp+˒�A�Qv`.�^<����%�6k0�
ݕٹ��U1ot8��<ۏ%�8�T[{=�-����ϧ=��o�a�ץQ=��LD4f�hP������v�cs�@6�2@�8���'!�pP�n��+�<�
œ�ʕ��a1EG)�w����z]��s�"m�;�1�l�O�g[��9q�g�v"���u�oeW&��=x����fn�bwN��s��l�����#���0I�OV�w2�� ���]I����+ks��bna{�y�}�r��z��;�j	�YZiU��%H���e)L�DpS�7�'�7�q���ڧLG�˝�0�:��NE��	IE���r��+��� C3dwF�#:�=i���-�,ۙ�����"\��8�����b�u��#�g!X�<7���g/'"����:�Z�l����/�K�q�R����AP�'m ���}I�Q�Ԇ���8��2N�̭�A�[3�R�y[�Ά�KnƦ�Y��ep�8�r*1;��En�8��Զ�ʗׇ���k1J���2�U�J��6z�Wq��ǻ��@�/Z|�p����tfQ9��;U[w�L������aP\�ȡ����9�y�r�J#8�#\iwu\n�S[X@�3��zeR�v��˛����* ���(�${T&mP��d*}Rl89[OT��ϰ$/r�%���fAv!6u��o�i
x*�MfVmL����P�ڦYb�ܮ�JM{,73a�	$ܛ[so�n��qR^�����mZĆ=�RR�C��3z+��vd{����}ܓ���Ю�Ōa]��.�q�rG3�9��\�xM�0�<�nF�L�{����7�nN����i�ۿ�����B{�=��Ef�}����ј��S;��]���Yˎ�T�}2��O�.�=c+5B��"��9X�z���Ov�]���u��eZ���h){�+!��
���0�֓m�ʝ���I}�ê�^k��eɵ��o�n\�Ov��ĵ}�^޾
�'���"`�6�#�7����|*r�=ɣ�N�qv��92��W�做b�'t�:��N����f�M9�ɡ��>ӯ�!XV`�e�2�5���L3�o�鯏	���h֬;A۶������7w`1z�M�V�\�V��P>īIyJZ2�r���Z��[.gJ�����˚�*჆+�p��P��p(nƤ�����ɗ�Vr�S27��*�J.Md6��AI�`�e�sJ"i�7|2̱:�S{�J���V�t6���z�7ީ{Q�x��ȚP�VM����A6���������ݛ&J]��Z�9ط�d�S�z}��?F쪮S;��
���0��r��9K9D��2�����Zp��b����ǧ^>�㮺�n�뮺��u׏�q��O~|���UU�x4S�O����U<�%S����R3"y�n޷���׏u�]m�]u�^�u�����y��o��|�;�a�P��QWNl����U�^%�"� �(��Y�	Bk{qק_^:㮺�:뮺��u�^=8��o[��W|�1J"(��%Q�}xW'��"�Aﵳ"��-CZ���n����}�7���mu�]q�]uק]c����q㏿��%EEUrJVE�*�+D�dUfG'ZuEeb	��{�w.I��g�� �Uʢ9D�Р�S�\.�a�I:�"1@�Q��,+�TW
���;(/��bTPE�Rn�TA\�PPP^��TE�\T��n��͙!!bPG#�p��EE�*�̧D��42KR���6N��Tz������"*��q9TU�9{��y�
,�� X��*�X�Ų%o�)N,��ۇs���7.�D�;��͕t��-�b��"���S0��(7燼�^o}�E
m�����mF�#m1����" �<�Ϲߛ���ª�n���O��|��x�K���z��9�-���@_�}���u;xA�/�#����*��x��p���Cލp�C���몶^���7���U�����p0������~��;�T0���kkJ@a�, k+�4~�?����������}�����}�m/�'��:ޭ#7�~@�u=��k�W�T�p�Ϭ������72�3P�ʚ��T�{͑��V����9���`�վp(3x�����t��,ZD�:�z��?�+��D� �M���aD	�D�(;��� �����%����]��}���_ɀL���۹��p��mƼb��=<� �����Ê�}��[�:���ȃ������8?�����.7=�.�������wg���f��a|�{-2<�dV�<��r��u�h*h{��E�����y�x��c�]�j�#�ѥf[���4��U����l趄�;c�[����t�+u�o	�aԢ����������5c�g�C�\�_�7���T,,��:�~Y�����[�`=��E6�b"����:�k��&��Ǹ16�@�~�vfU����}��J�]u���)��ua���s���9�3���w_���<�w�vWY���G����M�7��i�� 2M6�b,m��A@����s�7�m?%���e�9�+��{���՘�����0�g� {j�����-yy=�n''��j?cy7S�Ћfn.����X&�]>]���}j`�=��u�Jx��9�4�W����h �k�����3,��k�|�ɡ�-�j}=�K��`sxX
m�Lfc63ZWy܋_EO���<#���o@��M��`h9����xP�:�b�����ֺ`Fv֚���o_	�a7��N�=ئB
G��B"�ɹ�
����Q��6�v�wb�)ⷎJG��׶�7�E_�^տ+����22�~�7��O��l>�\����t�:DunU�w	Z#��>n��z�ɹ�@��P�.��=��x��7��L�=��ݓ3�5X/��3	��KI�-�'��1?0���,�+��@ߔcxn�Æ�1�5ř؋뮳��N��w�~�/�^��y����O��9�6=v1����t5����2왻c�nrG��K����C<��d�Q+��]L���oS���p�<MusJ����^�2�f?,��X�Er�ĄSHkj����2	�n��~�!_W�
�Rn}��q��1;���J +���9u�U�wS��KS�]��N�s�� �8ƅ׀ݱ��Z!��cR��X����� �o����6�M�l@)��m�%4�M��*qA	ï�G�_S��~l���V"���%��sq02�m�5��s;%��S]f":��pS��6m⃱w�b(g\n)219��%�m�nvo�y��Ǉd��q��QE�>F�/��$/�������X~��C�M���.E�s��v�ճ�M�o2�ޭd�׾��}�?/��b��"�-���7;������6Tј鈧y�N����v��#�5����|��pL/���2��kK ���
�Es�6F�{�mi1�<[��̑8��%��5x[{b��p1�I�k��޻�ݯ��ZZ�s���g����N��1�=��[�~^��Xo�w|����<4b���h�JjhK���Yܨ�A�@<#��	��~�Olc��-�̛AcM��v��m<�1���;y�J1�ƻ�2uU�Ö_1��Rw٨5���'���	|�5�9�����Λ�;1h�뭋�J���+�ֶ�ۑ;�p�y����f{��C�h��M@�2�1F	x����e�!�3;�g����,$W.��jr�_�H3�{j�~C�Ā�@RM��S���[��e�w�zv;ˢ�E�n`5���29�s@��ח�`�DKj��h���=���p���m���(���=վE�=kJ̐�䌮�v���F*1/`�� =�'t����
�j��{�Xvp�J��EH�s{�P�B;�4'w�5���Op]*�w��k*���ƛUcm�ڭ�i���M6�b�$BAD�^{�s����~�r��k��l���-��Ҕn�y�3�&w|kg`C�ˆ��
���{��la�.=�TG����EO�ϔ[ޜ�B�ό�y�r=�4�j8��տC�~�qKy��*�Z,��v�f�Y��!��>'���g�������M�4��m��r=#�(^,�	M���1���y�a���D&/�f�Ʀ�'y���y��9uۯ�m���k ����i��L��A������z��[�ׇ��,��(�g�36���f���r� ��;�;/U���/`<^ת�(Z@P����ʃ;(j����2�|��|�D�'�F��=k-y�Zu~Ϩp�)�D�\����[)�ְ��������Mͧ�ú3��	��m��7�OM	�8�����&jPb\-���xsy�r+UCr�j�Λ�����?�P���4���=�����3SM s�SN>��y�v<o�Q;�w���ZN⦾�'�����,$������M܃�*���Ⰵ�+����U�wl��]Dn����0��w:eV��#��Z�%����1y��+��)$�=��.�v7�/tC��]��U�[��M-aY<PWNp|9T]�:y��[�[�u��w����޶�o���D��i�F6�M��@)��l@#m�؈�W�zs���EC��@wq��=�ә�Q��sW���:U�QqYW�_W��~*y�O�+��1K�33o'���|5��fbî}��\�_��]�-�[=��LQ�oHkj��]>�6Â#��4�,&������.1���[�J=��ll�λ�����|*��|&���Ф濱r"z�����S��J��O���ݮo�`sN���7�r��!�:��qR+js4��������ۏGC��-�� '-�+��x`{C��x|+�v.:߹�(,ӱj:��*�]$�v^w�f<��/B����?A�ێU�^ޝa�iI/��= ����N��R=�i����?��,r�X��U����@���Ʀ7L��� �ݦ�|�;([{ܫ$�:�^8)� _[���_�
��֦v0h5@��Z  �>E�P��ʻ����1�����g����P�l��I�h,���RRy�#��`*}�~gl.�Em
ǋ;��3�X#�����M��Z&��{����@�eߚ<9_+��~��X)������߁�>�ta�ci�m2�hu�;B�N��YV�WeMY���:���s�w-����|GzX������VA|��K���oh���V�e��]�Ѝ��m���[+~�;�gh�4]���/���Qח����m6*F�i�B6�M��]�w�����گӅ;;+�->V| �g��
'�T|��:&~��M�ـ��M3�va~�5Qxx���\���sSH&��S{4���m4�l��٤�]��n���Dv���Y����5.�ݪ�����m�w��4x�̥�VM�ץ?#�P̿~'tiD��c�Q�\�L�Won�����9���}��-��{_��L�iwW���'��Ɵ`P�D?�3��+�v]��ďc�|�� �4N@��j��H�cк�5��6�D�����E6�5E�$�lf��fY%o���������6]�1��!ny�.5;x&��Wd]�k�l���+8s-�!�t�[�h36r�^j����q�`^X��sοx�M	�49^\� c��(��������uO9Suٛ�;Y>�w�1ʭvY�;��U^�Ϻ|��U�o�g����%�ҧP�)�������v��%��z9������� 3����â|�D?�a�9���'�7W�w��i����f��=S�\��\���xmz���_�V~"�wPs=��`'��nA�S�o��]F9�u>�"[�[]!�Nt{yJ�]6����YT�(N�^1W�����/���}��,�?�p��=}���%+\C\Qͮ̄���Y�3R���c��%C6K9�[��������~4��ah�V�m��Q��i�F6�M��pBC��-��%�&;d\u޸��||�/&%5��������@:����l�oc<�1�F�Qt�Е�^��zP\[��7�5��0R7L�`���O��a�B>�t�o=[�wwW�w=�^a)��fG��>����z���j5�%u�x�z"�l����s��[1�:�����*����?��8���X󎓽��49h�2p;��^�M�~�����y�4n��\
�rs����޶2�w4����} _���� p����,uQ?�煀��l
���r�F�`�ݳS�j��-�ݭڝ���1�+�)��ǟ����Bo���Iu3_	�/�*%��S�z��FO�w���TY���#o{x�[�+�g�N�hN"�1I�-��2q��` M�bm��a�:.o]_i({��"$\kx@�0�6�ۯ���[�؉(�����2k����tf�"�7��	�7��K�c/��< ((�������N��Na߳h��oǄ��S��C9�.�y�AwQ�q�����]�U2/�gӏz{��\����ȸ���j#S�*q�#�m��JX����X��Ru���޸ �u�g႙�����Y�Z7����q��|�0��8!?n0̐�H�WUU�r��vr� �oX�jM�ʳ���;�a��7�.���3)��o��*PD���,X1���د^�v{��l�������S-����N��m�G}������ٵח}i��~4���M6�`m��D#m��\E�Q�{3Nj���w�l��c�V��y����8�xO�u�a�h��`9�����e��me�gc
ް��<t��+M��y�
L�X���^�l�T����@�Vj�n��0��E��:�M�l��h���{�zW=�}d��\Og�7�0Zy�{5w�����m}�k魟�j���8���z��OP`�*x�P�>�j�L��a1��}�`sZos��:yW�XZ1�B���]���\���:�zcx0oi�m�}�V����m���攣u�3�@O��W-��{an��������~ �~��Z1T/��2 ��S@dw8�p3�*�>h;�٬�(~�{Y^�ג�b��{�ɫ���$?�]����ōG�}�R,?���ZE�|�*��Y���U��F����걵��`8����i��ϔ���;�?����^Pﹴ�v#���	���l��|`�Y�"� ~���4_�?Ef-��}p�,1��q�m�G��ۆO1�3�w�����	�o��E1��n��ǿ@Dq�n��b$(���d�l�o�1Tb�X����dܟg�QiS㺮�ʕ x���L�jz��1� ������'l�ˊ�.�GE���[�R��]ȺK�����z:�Eg��F$��I��W�쾼����;�����=:�m�Ji��Q���`$m��R⤊H�� ����,[ݽ�n�MU4LMok|"kuJ��<�j���;��?!���r�(g�@�f�G~������X�9��x4+����g�"L��+��o���n���]050�Y/M�[#h�ݚ��%�2���˽v�R���W�.^�T8F�Z=@ts[N>�e{�a�vf�U�����ؖ\_ѣU�\:���aU��;0�O^����|nl�V� �Gf���QEG�4p�]������U�0����{�	�>���f	��--�l<.șlx���ӡ�;�h�-��ۺ�*�Ph��qV#gO��<�����c��5��ث]�fn�M,ޢQ�vK��%�Xi����q�n(Ȯu�H!�Qzw�xl�S�Ӟ��b�o�Ts;?0us�@N��kG<���~�� �<e)�B��`�W�<�+�ֱ�m��^I���AM�7�$��S?�Q��Sý08?���oz%��4w@�B��H�3�jQ���6��:d��:U5�R�8"���[|��c �;��18��?T�7�W����k��|�_�yՠ�X�֤ࡺ���� ��2�h��n�݀�]c� �;�i$|��	'�e�a���Ji�4V�*�s[����+����:��u09��}J�j��R��_3]��H����=��M���i��M6�iqB�m�G����uگb��#�����Jw<���z�ኽ@D�4�&�(_�R���Ʒ+�s� ��+�w�	gE�_�;�!9��z��G�{U�{S�
����ǼT�o�7�=���d����b@������O��(������������^Ey����)���$(z�#qgn�8?�Y��߾w�㔍R��z��ؐ�T���bt@9�Ce���Y�5��n{��8�{w��������F���Ϭ7�[�z��E�U�&}�,����i)��X���7�l��<���/~��ṕ���o³�����8SG6!C�#�י�&Sٜ�����4��gxP�{dp���O���8�c���X+����sŊ�{�5O�!�!g8����O�X�`�f݊a��lǢ���gA��mc�4��	��Ф	Ν�[���n�=7��8r�V���e���w��R�\�_�� ��t^8f����e���uR7��~�l����F<�����Gz?��y�{�rX����z�����xxx �Z�c#j���̭���\�f�Hf�QJJ�B�R�z!�N�,.C���Φ�n�Ѧ{l��;�.}ca��q��X�����jZ�r�D���V�q�!�)%ջ<���wHR�]��wMY�V��L�u�k���J�iu��E�<o�N���9��ݴ��j�fnk�]Y�R���Z��w�yN��X=�t��x�'q��j]���w'#Ɯ�M���&K��c�CH��=8ŽwK>M-����U�8�<ڭ�5(N�;��{�"̣(K��fwCp�0r�fu>BV� 0�����:´+���Њ����3c�O��e��;�����H7�^� \����R�*y�r�nW�w�z�������pJU� �J�5�e�p�R�����1xƞ9��J������e»S�Og���W�!\�"��=��|���&����l`n�&��,Hv��8j>�����]�ki�6����ku�t98�W��T���ݭ1���n��<��V���X���螖�.�A����j�+�cso343 AW#�7 ��̫ͭ�Kv�^�Nٸ����(s��Hͼ.�:̓���Zu�傘��^N8v�
$r���f�8��|]�[vK��oҰ��<j��҃(�\B�T}���a����:�����	$]�I?t�o�o.�h�.�5G�
���0�3L�Y�8����9լ@hݸ� k֤ޜ��w_w$��;&o;���$�Mi��+�t����;��i���'%�^`�����;C�W���S��{7�Jɂ��z,�]�0�|��1���}3&���nݱ+���Z��zxU�΀��݋�����l�8��)?��{O*7�"�����&����r��,8��&==O���u��0Kp��Y�v��8 ��R�=���:�h_:ۊ�U�[Mھ�领�ü�eb	���;$��&p{�HZx�Ҫ�X�32���m�����6^u���.�I���5uY���b</s��(�^ۃ{�4CN�Z%�ͳ3�o;#��ƮA/je�۝wtu+˂�x7��hcW�����maY)\z�WNw69�2wl��
��T�����fWB���`��P.]�v�}�%�i��7���+h�=�fL�|�D/��K~�c �=Tes(Lv�HfvPX��Ʋ�i��!�U;Uu`�eB�of�<$�¯�򎚮S�����C2�D���]�&sณd�)�&�]�4�OpI���l��A�4B�!�T��=z�N|~����ة��TS�Q�'u��~{�VHBwV]J��Oi���׷_]m�]u�u�]zu�Zu���q���|w�\�J�Ŝ�;��;�#�Hhhr�/��<"��F�I�CtQ��oN������u�]q�]uק]u�]q�ӏ��y�|�ʈ9VI�$���� .L�21��>��+�mR�#*���*PT�X�n������]u�\u�]u��]i�\q�<o\�9q�(�!���ޜ2hN6#_�vQ���q�H�;.�5�m�����]m�]u�u�]zu�Zu�x�||��5?�N�
�����?�����jU�r�+���ʢ*�$9���Uⲹ|N�)O��XP�_Y�f)i��VJ��� �6TQ*
*�L�UPD�/\Nʯ�.TRaI�_L(�zxw	Idr�H�R"�������"䐁ӡ2*��͙"���`)?VUL����B��Q�KR����s�G_�z�aPh�2.�L"�gJ�
���>�W�IS�T��7�Uڥ��ⶶZ�v��PI"�EL�VT�VJ�+���A�MF���Il�E%N�#�B�H�nr����cr�t�"�4i�l�����J�]�S��^c֍��زKZ�3��)��R��o:J�e!����L�9Xx�n&�}��R	�̚�]�`�B"֛�+�F��u@��h��Y^��`�m�E+$B�2�KTem�db�i�Se�UX�^��R]Wiu`�Ւ&��C�E��Z�*mT�89M@�SU�DTJ��u��aTuG��(����P�d�N0dj�����Q4ӎiEwx���RF�ib4���Q�]z�4۱0��7VUh���C��M�ط��i��m6�q$��i������箎�mJ&&xL��&)�c^6f�'r�����P�4�����M��m]�3#��j���j[�J�k^^vH�a��[��oO�����rԘ>���g�	�V@�>��2l��I�9N��>|<�^3Ay�og4mWR�Q����`J�l��r��/B��U�����o5���`g�Ԗ�|����/�%WNfd�s���/-]���6�����^[�?�92bna�0��7^^��Ei�[֜q���{O|嫺�G;��O~ji݀����!�s`)]�oF�m���A�L)G!A6����5��B?/��^|�ϣ���o�K�s�[��yw�p��a����)�&������E�P��31��,1?6l�0~N��̪�M�[���B��%����E���r�A�]��\��;�7����n}�>s��C@݌c�Sr�%�r����`UO]�%�����<�{��b�	J���N/�~̅����2�?��[fl�{�c{�6w,�(�XdNQ˸*�p���'�������{_}W��G���L	�y�����2}7��>��u����-B"��i�M�^{$�4��]���OS�iv�c'�bӮ��cZD:nm;[,�ۚ�2�m��w.��w�/:�u�;k������K��"������WKvTO�V�����u�#ת�^D�;�3Y���\h�+U����;���gA|��u��Uf��>v��UH6��p]��ː%�
�<<?x�`���mK�M6�`X�
i��PK�2#�~y{�}�Ro�e~s�u�BVߘiqg��ߒ_��Ӷ��k�{��'��t�on�/�=�s��z%�X$������y���@&�a�נ^=o$��B���+h�r��!��[�oh�:������{W@� �[��J�a���p�q���Gv����x�N�7��5�mwWmP�?���54�9[�8�6���\c 컗\�UGv#xcб�m'�.&>2jgk��x(�	���0��K�Q΄�AH�ֺ�{Z�WSS�tLy�57T�֜�T�����@f�h`���H�r:p^'Ԧa�(ԟ������Wx���MK��UP����Ժ�zQ� ==Ǟ2-��mƻ:��wl�Rq#<Dph�^mw�0Zm�&�y��ldsH�#w���i���3�fugUҝ�i���U��Ml�`��z��[�E�Э���F@-�8�u��q�v.t^���+�>[�w��vp!��ckty�	�~��ح�j�\���Ȟt�?m��	��l}l�5� �5�
�U���\]Mɣ��1�:��jb�R�k�-M��YR�+���P�$=zP@�<i��g�WV�M�Yٵǣ�W6��$���w��\��ެ
�2�\�b�"��DC�x�����{�SM���m��#m�ڀ\ �3*��DQ��gv�����V�ͻ�$�~�#����b��?�?O����QagF�.����uc������静�z���zm��"�3��]⪅}K���8�	<7yޫߩ���d��v}�qv�h��ǆ�u�e ��^�ɤ'��.��8�5�\��l7�w�%��w�w�^����:z�\�D:P0c�w��~/������z��"X����k�C{��}�5��"�����Ԟd>��s��G�{�P�/;�i�~��r��&��	�j.�=�����y��.#���d�'}��9�L�9a�(2��稛x���\�Y��g����z���ڲm|+���P�k �v����>}�k&��!����qr���us0k�_.͠	>��5����)*1W��󉇟J�inj��P�M]M1Yܤ�`�;_�SH���ȥ�+��iK����f���0L MSC�zz_�b����k�����[[x��g�"�! gy��G��֣�r��#�Թ�dT�	�����'�7ͅ�DjEɌ��w缴��eXʐ��<�@]~�W�U�����4��z0��eC�V��(
��@���$��Y�8�"� �[H8φ�� 	����HEa����8J�#��\��lq�i��qL|9B�R���ڶ��u�W]o~�s;꪿?�i�cm����mn4�M��P3���w�=�|�{N��_���ǚ�T�p[y�2"�#ظ�`�6-�Zy�f��r����}���\���ؓ����ƾ�x��O��}p�77R�}�SP!>���)�,��¸��j�`�f���=~��Aҋ���!��>=�S�|tb�P�Ѕ��kX(Y=�$󂣎=Y�.�
q�3�ju�N����j'>��w��_]&���ܽe��b����QX�%���\\�k���A*��d�d��:�<�e��ƅ�7�¶=x�v��P�=�'��Q���:�~S��t�W?|^�ז��C� �9EctS���%�Z�dK���E��>�MӳszmՇ	���0[���!O��� Άf�_�{-�1̺��"����1Y��n��#�C�[ʘf)홪F��0:�ѻ�=`;�����Ui]d�FF��q��c���r�0~��y�a�����[$N򆧮�����<� _s����y��[�l3hPǺxcC ���8�B(�y�?s焽[�P��>�<�m�/����p���%v�v�T�.�R	7UnUXSc�撤 �p�S��0d|(�[C��������T�'��W�/�Pn/������rv��H>�k*f�C��g3�s|��;�˞w'�~A$X��M� ��[��ַkv�ݻ[�����ؖ^�[��6���<caK��8�k����l-I=�Fɕwū��9���F��;e�W�.vM)ܪ�{����&���L�E*��Y����~��?.64��c*���+�ˢ���4\r}u�,9���&+�=��"�yA����F>���3^^b�Nĳ���NX��&��oq�\�k��(ײG�AoˮH��͡��h��Ww�׸��F�~�¡��fI���f�:7���-��Z}���vTϓE=��p��q����	�.�K�It�wߖ�ٳ��(W�}��,ؽ(����H��
��˷A��� r��=3.r�_E�&�iVǖ�&�)��{��cPT>��q����x܇���oJu��:2~:p�v��?�׿�����c�M�^���-�;�mji:=!�#*`&��w[�O���,+{�7�S��l�'����-~U���<�l��K`&;�8^k��s�����2��FS���h��8;�=C��{g0x֖��ǟs��wF�]}����ʸ���H�#��둲�< f���V�������3t��굢��ZG�o��>q���>S�3�uXh藭f+����ٮt%+�5S2�u4��]CZ��j݈�y�y��ߥ���FK�^U�H\�~> �	>>�UR�g/�����l��5���������y7`ni��H�eo�V�M7�%Nª�� =��/X��mX�m6�m��D.ɫq9�K����`�1��~i���??6(]<ٿ�7���{��C>�}��:�)QҪwOa�`8�<�u�W��5�8"(y��;'ɿC��fTr|�{IQ�S|zξ%��W��١���%^^��e!�[˺XP���:h�4y?s�3a�_3�����{���� �;�z����4'!�{��E4^7��#� CG�I>vɿ�Eآ��qos4�y�D��}u�"FBa��9�vMD�i�so#\4����Ȥ����o�$q��q�(@^.�!̹=D�߾�Oՠ���5zh�{si���D�c�;��[�1����ZゑN���⃔�ڌ`�c	�;�ۂD�j{Ɔn�0�z����X��@�z���F��H�=�0T��44��c�Mƶ6�rָ����٘���pÙ��Y�q�.��AO�n;���}�_K�Y��汽>���wڋV܎X虇W�R���]6��K�ys�n]���f}���~>1�����m%�{����_�l�j/���mh_��Cb�i����'k��mg�G����}u{����F�:��		�X���i�+���3��6�u`��Q�Ϊ�U|���gD♙�%���:��/N��v��w�l��C�צ� ���b�1���)��m���Ϲ���y��\�x�`���~��0��]WfK�W�Ƞ9t��םvx��n��ơ�г0���c�`ա���v���[-�����7Xσ{�p�����
���[˺Fj3�aA�&�Ý%��@���sV���̓�L�dl#��T�Rj蓄0I� ���%�t��w���A��7����zF�A��lVI��Gs��j-�V8���4H�";�������{+�мM!���A���~1h���%�Z�=r�gv9�<MLwgi=l;��/�9M��z��
����C�_�΃Ip�(Bb��x�?1���(�pU؞�R'���c�;#&�S�����S�%�kP.�4�=�7���ܤ�Q��#:��a�$_zj��~��z�8�b�cg��q��������e@tr��_���:�>�^��4;8��5��y���=MA稯C6p}#c�u��Y�΀CN�f�;�9����zΪ��O[�4�s����5�ဉ� |/�ii�j:�~LJ�����(�dh酓�o�C��D�������A�ĲJ�d[|�kꊱ���%���d�6X�!��1G��0�f淇\�m���U��%D46&.o	n��+2S��w`v�b��r��b"`�{x>�^�[䳁�Bۊ���]u�O��Ǧ�B�4�M�m�����bH�D��6�߾��7z��'�f��� �}f��t�LA�( >���F�6��͵�;�Q�b��˜�9����Az�?-��un ź��P&�y
�B�g/�m򟡘~�~��t��wpw��?��ijd��~��g}\�Pn_��f.��0M�ɚ鍍Yw{}��W��\N8"C����4{�~pϼ���J��`A�a%韉���L]�-+��ٺI@;{Cb~輳~h���u�k��<�rn�O�9�W,��M'g����U�������XG�y�7�m�M���~�_���~0X�>b*�Ev����D�k�2�0!�7����"�S�<z=)�NoF|�
��jq߮�QW���2�iba�r��Muc��P��.��tz��X熟6�>>�3��o����;��l�]՘�s3�o��;�U�a4}�	W�Xw���ZړӼk�g�=XtBDJ2#VX���&���ܼO���/ϵo�b��د>�|g�������T�h�<\�Rq,Z�db�G�O��ATF��)-k�q��b]�Z�T�$T:�WZs����*7�J����� }��U��U>��o�Ƿ�=�0��d�.�.�cw3����\h��R(S�*���L�a%�;m�I=���������M�m��cm��p*�Nwru�E��r��_�;(ח��R�υ�s��@uΒs��+�.M�&o�u���t5��ɟE�rTk3�-��=�_)�������'ƫm}�6���m2���N{B���D�������0M�'���J�P�砢=f��tC��<R~�t�Wpm���{dE�D���p̱��-��h�ϯ�'���F���$h{m5������C��M��������~�a~6�Co�f����jz>xT��k.��')�w/N�4�[�q=�v��|��z����1�}�18v��s��oM���KK�3�����[n��n\�Գ�Ïب���?o��^����R��V]��x��%c�؇O{}�8珦{e�\B����`��"b�^���w�����-������n&����n�wp�ch���.%�k�Z��9"ۄ�' jz%e
F3��Y7]͙{��Ҵ�xn��A�i�8��pId$W����Ё���8�^�M�f�ڽ�����'���hg|��\'���^�����u�G���^�Lh�4O�=���	y��"�'��d7Y���f�V�ߴ�2���}PA�a'.c��藲�ʯ�ڌ���F@�'�����Ӵ�����^}Y|��}ا%c']��7n�鼗��aw<�$�ީ�3^���(����|�xQ���#���S:�fNhR����x�[B�(���j��W�}7��ӵ�m�����-���I�~�!���M���m#m��F�G��6�;
��M�>�����~�6b���(V�;�gצ��`��q�:���kf���;�xKp��(��qX���I}m	@������!��DǷ;�&�{ɼ<U��*�v	s�[����w�w3lG�'pD�w�uBc��q1N�~n��K��By|�V��'f�.����ӌ.���͞h�<2��<�B�L�n�%��{��@m���N5햩�qF^��۟���H/?o��s�<g��BG˔�.�o�g.��^�OE�D���C<�B��*-�zƾ,��8k���S(�����}�0���@`�Y�s��6#�ϗq~c�|����|ƺ+�9\S�gx���>�\��h�6�3��l����F�"(2o�`��<��i��3;Z"V&���W�����d7E���˟}�^���ҏω�>�sڛ�/�BKP�/��[��=�ƌ�n��M"i��'�*M��}\��k��F�frH��xn��VS�yדs����=vy��t��[K��[蟾�0�Š���G�wP^�=�`ǈ������5��պ���o�l6�X̮|��D���i=y�!w9-��`�l���L�F�EQ&��]W�ٰ�D[��6lYu�B�Y�;�*�8��S����&!�Q�J��	����HQ�حvEb��{j�ګ�9�/��s�֍��[�n�h2�W��TU8�:�/��y��"�X ��Ƹ]˔j��d��=��S �e@�:�.A%`�Z�TuG�ӝݣ���70\���˓:2J�N����4��Ub���a��,�����E�T32��`L�.��ku��%m�U+��О�d�$-^��b*��,��۾vl�%qÚ��uԃg6��
����[�pW�u�e�A2��bf�,y�9�qC��)T��֋��F�ư�Ճb�]��۹0���lE�-�.��Z-�����e �<�!�7��]�ƀ����b�r��8���&\!3�P�]�����n��A]�TA�\��e����-uN�s�����A��mv3����x-���~��"��Y�X��e?��]ŉ�anɣyP׺�:��UC ���՛Brs�M;%.WG�)]ݏ;����u�/�*��Z~����h���+ʟS��U�D���A���lע�n	�:��>?ED�[���,L��F��)Q�Q�PC���5���ñ�xz�y���k�����j0�댺�S7�� &(pI�_f�]��W���i�(EEI�;��צ�[�e){ȧ��:��^��y�=v9�E^PL�^���וKH�Y"FZLJ�B�X:�VߦnC�����5�t��f�$�&�+d�s������z���&���˱S;4�a��ʎ+�}��%��k�<�9�l�
����moJyha�V���6��ei�0�ܙ�s2������e>4�y[l�;ۂ�ke�q=�V�A��J���3M��4CxfY\���!���os����t7n��a9[�y�0i&B�}�|f�l�k�M	�:o6���D�z��QWx��E혻�uU�JUVob�]�r�t�d��E�XE����<��1u�c4����a�� �����K�����������uwq�:�^[�'>:j�rf��3N����7yy�w��8��P�;�جhei���lMV�[��M�Eξ��좻��/�V�*���kG,��^�նUv�h*�]|���euݵʏ����^�-�޼�С">�$7;M���ˁxр����&;d*���5�z���IZD=�#Ξ)rќ��!�s���{o��*�)Y]wq3�t}�U�mC���=�ʧ=��ɽ�X�Y�K8�k���ou�iټ�۵���"i �M��&�s�YkEz+'�O�\���WS��	$.cm6������[u�]uק]u�u֝u�8����?U>�C���2��|y�UɑQEAU�nݹ��^�x�n�뮺�뮺㮺�n��x�߄ y(�R���*M`EWĮ[LM�$"jK�.D��Gv\McN:�ۯ�i�]u�^�u�\u�]m�q�{�2�+�hDETW�۴LT.jT?&�G���v��o�����N�뮺�뮺㮺�n��7��ς�ď�EFeI7�c����c$���~�w2�DJ�
I(�_T�N�*4�T;�s�}WD�r��_���TWw��QO���w8��e^��Lª佶ܪE$�*-Y����(�D��$�?{�m��2L���DX��Q��f�#�H>G��* �|�X��a�DG(��L%-���1&� A�_��V�{ߝ���{n$�IORN�ױK��u>�X8!�l��yC7����7�I�;�8����?:�M�)��n6�M���m.Lm�)WIo�O�����z�A�;ӏG=325ù��UC
�}��Fd^ׇ��ݾw
�3�5�S�>{���Þ��f,%�#^�����s��	8nPi�Оh����9~���ͭ7g��Ğ��w�j؏��'��D'�|�ԋ�9Q�Ңkl�+���o�� c��Ct��t��w�T���d?Q<��`�,�m\��=����������}H�J��S��z����3r�ԘK �@�.���)�hzZ�����y����! �B�\�E��-9>��ծ}]`c#qsL�PyR�a�oP��H�f.{�oxy��
�Fs>C@����&��=^=�'F=L6���Qӆ���Ǧ�\����Qn��쥞�q��b�:n5^�����Pҧ�|��/�ؿ}���/HW�>���e�~�Z'ooH������Y|NƁ�:��#�~�j`���T��٬O�~�i�]h�3)�	���)ɿ�>��v'/�auXˠ��&N���	�>��F^Y����P'�ί2	�A�� �@h0l���[�*yt;l���s�3����ɓhr�l����%o��4�gM�Y��'i����#��M���n6�M�()��$R���{����~����qO�	$����oM���/�ݢK��z{�m�f�@�D�8�$�">��v��O+9��m��<r�cW�n�.���s��*�"g|]"�:w��ѓ^|���}�����ԯ=]�L�G�~QoL�Ԓ�kSз����l�C���~�e�722�\J4|����9ݯ�Cy~���Se(�`��r�V-�HwK��s�N��c�F؇�|����G�5Z���]IJ�v�\�~��_zY��u���6��y��y���D�p�[�-J�ףT��3�o33��!ފ�gۑr�יgx��#{ϊXy��ދԤ�R��؍�ob��X&�uA��67}�Ѽ*=} P��V��ZDKz��sgtyAFxl���-�D�%*rR&�ljc绞�cX8��l �E��{;����w�9;�i������~r��utvف��ݠ�����5��gs�������e���bM���q+`QlcP[���uĎ���$��Y��J�7|o���6�7n˃9����S�Ϋok����Ϛ|i�6�M��i����d�J��ޗ�nu�w:&W~/��K�u�}�6��u���KV����܂�X�凂7{F6�w��d]���7��1t���m9"�L<�߷�3�o8���jq�?�!��(7v(x ]Rwl���Z���R����%`�z��vԝcL�C7������0����nw#^�Mj1�5jigm0���J���� 2���c�+T�<�@l=SW�����6ou�Y���E��̄d��3i��j�^m�g*f�O�f�?�#�c_�	�8;sD�οd�j��z�99�����k��r���o@����g�[/n�E
q<�Ʋl�K�Z�$ΣxE����F�b������y㞕Nz���W�^�t)��r�Ķ����t�Ux��|+�r����R�컝�m�X�LU��w�z������5~�]�<^_O����-����|�_���ޞg{j#U�졽������5F�K����G咵f�Fӊ��et�*d����+�J@(`���u�N-ۂZ>kY ��3qm,�(�ՋV!7Z� dx0r�oeH�WM:9h�`���q��Y6�G).�NEf�s#{�����󪮏N��W{r�����1���6�MF4�j���y���}ٽ=׮��xs��˴����ĸ9��� �����swd��;������'�^�l�GE
��H�ܟ�*�Y��>T�Q���/w^3{zn�kX�`�!���{�ˀ�2�ŗ8���U��^��վ�h�t�}��o%]�0%��ӕ��쨫���F���ח�H{���,����nSn܆��9h���q'���Ɗ �m�R�W�FY6�h����
/�zl�dkr��I���)��gP��F���W�w���k��¤�{��bن�Ao2aFٺ��}�!��#�S�嵭���k��%^ݠ��l�>,��������S��^���90�:DGC����;�3������L�ea��S3�5V��e�o� ]}a�_+�y��&����o��@�q�ߵN�9�e-r~2'0���5>_L�1<)�y�:�b��Au�="}���pHZ�%eq]N�ٮ��԰n�%�ԫGvp�Yl�C�/C�+"�R0w^�
E٨3#�Ӛۛի|ʾD�(p�2^�^T]Cj�lo^	W�K�*ç�w�r2n�
G��?m���m4�lm���=�ϯ�Ϟ36^&#���P>f����:~R7ٞ�છA�VKs���q��dܳ�SK��u<z��ϣF�96����.Yu�{�Vڋ`��概󜒰BL0Vǟ�Ǧ�W���&"ѝ� m�񼛑'Z�n��Moo`�w�����N�IVK���z�j� OOX��mk�NţYy���9M�U_���{��$~�}<�X���qg�Z��g���M*��-+���h���ED�N��8wz�B���e�!���"s��[{/:�:.<�b�gz|��TK2w@׋<KS�R9�{�p���{`�Y�4���}<���>�����\�g2�T�7�O�o�Hg5=�`�[Gy8̱�Z"^�Cmy�Z%�f"}��V}�w�;^<Pi���|z�6y˛̚�5�5]�Ks��po�s���ö���=�ףx ��fx����CA���v>	70��n��	����a��|�5�!�ן6,Ş�È�x]
��
!��n�W6�񷯵-9�V�wu����W��ה�������:ܗ�oU�g[��ߕ�g�4����i����ı]B��m��~�����C0yLF�����螽m�͎T(wp=��9&��m->���J�՜[=!C_���sa�5�+�B����uUr�g�?B���va������e�[�JL��~�J��r�r�-̍�9��1��wޮ�9���>�ɑ���^-��o��JQ}��t�D��� '��ur@�u���no��	� $`'��i"v�Nvv���xZOÑW:W��ػ�^�^*��L�������::�\��!�8�p�L��5�N4gz�@a{��ޫ�z�����L�B�ѵ�RJ��S��]9�DB�O-5uB�c��5�c^�m�V��ݳ��@�MU콡��H���sUA>���U�'n'W��xLZ�{na��k��;�p���ٜ~�>YYB&'�ķn��ʮ�- >n�@ˁ��].ǅ����+9��O�������)q&��lˑq�J��0<�g�����I���!uwX�r�@��9#ȉ�'ni\f����G`��wԴ�CM4���m5%�^�s���M���1E~1R�A��q�❽\�l�i��q��\�}T��:��ht4�t�xr��%�YݫkhJRIn8�?�J��3�r�{�o��T�V��@�������OQJ6[��@�/�.*<�`D�5j���*O�S��bݟ����6����u�ͳ��s{���+s �-�8����[��sW����F=�ܤV��4���mmx{��3#�ߝ��=��;�ZmA��0:.��o:J��x��ip�/��賉�����Q�,1�K�=]�X:UW�^w����r������;=�J[�7H�}��k����3�J�*N�Y��X="�E�
�m�3����7�T�84�3[m�s�7ۙ�s}��=�v�\sZ�]�72U@�0��m�/9��k������b��O���&�_f�Xɔ����l/oh�f����x�{���/Ř1^3�@�O6����
8U�Rw�j"��=^1�;���-�bm�}:�X��Sm�\5j��;�m������R�ST�����iםU10F���m�;O_U�Ȫ\A�ۭ}�U��u���or��Ώ��i�ƚi���
�q1��7gv7��i�s���,=3���Å���N�<}��%�.Nw^�8����ګ��V4w.g�����C������{���!����O�ҭ��x!߃V%⮞`��Jեbݝ�5Qp�!�z��-��Y�E^��;���r�"��cc�M��8��(L��>�<������4M�ř�=�������:�J��w������(�}�
��i�q�'u9u<�ު�n�QݪC���\G��,7�+닷�r9�X��&�Cȱ�Cx���	u�Iز��V�WD��<r��v�����_�>o߶����~Q"v5��u�߉'��xݚ�^�޼K;��/7�= ���Bz�e����+�?,��s������;�G�կ�\���t�l�]�����Oc� dOM�x���\A�}@���z��Q9�yg���g%�;y�ڌ?&-!�nс���([B���c���w�tP������\�&D�2qm��X�e�W�I�y�w��T���tXn�HB�8��v��t͹Ұ�ѦC���I)׎V�u{;��~c�CM44�CM4�K�=��ϱu��0W����a����,v�}��4���	=�YN/6S���kk58����P��WN�p���O�s�6h�vmi�wp^�\��L��"���7�O��{� H]���қ�TG���x�>'��I�sd_W�wf4���3Y�1c��;�\`:"���ZYٟ��SύQ�ܡ�4���$���z��ޗ�pN���䅳칛Ύ�+I�藏Z:065OE��`��l�I*#��X3:k�ʗ��&����#[�[�U�f�jS���Þ"A-e���K�3;��ګ��d�i��ty�ƟL��]��` ܐ��!��$��;eLR�o(1p�z�����i`T� �z��W�%>�����V���G^
���+"��5ڎa
��`�t,B�LO���vuWP�Zވ�i��'���G«m<�|vUKy�壔�2�ejl�i�kq*��YR(���<�q���(�̆��r��}d��K��C���fi��jN�2��;���K-6�uTPg	|+;3�uޯ//~F�ii���i��#�w���s�o~��{���}9�6��(��n�Ǯ�>@F`��L\L��K�F�T.�!����,f�ڥ�һ�� �¯r����xڝ4�vg��� �Eh�����k���I{�~�MǸ���[v��þ4�35�=_[3�f��Gh�@��c�W��L#!�׍��m�C��NTzmGH��Ժr-]�4�Kvzth�W^�vz��y�\����٢�l��	h8���3�6G�=�~�� \r��yOin�bRY���j��v������ۓ!��]�����=1>�7�7��b%�G&c��iJH��4��QJo�߰
H�̩�v56O�FfLn~��Z��f�/��{z�l�۔V}97�[�IF���옿=�׺��tv6��_���n��l[�(�1�>��շ�/2E�V3���5�l���Q���d9@剼�P���t���q��R�&۩���u�T�ʜV��}�|,��4�d&�{y �Z� �4�p~�^�m\5���1Θ����x<aeU>��6�����~诟"q�kP��]c6���Y8��Ͷd��['�7r��: y�{Q���9NÔW:=P�77��:�6���2���\��o�$݊�\�ne�S��f�=���J�6��,@\wn-����>��]��܆�U�gx*b\�OM꛽���'���u�X3g�=��x8��gXP��Z���o��jG�C�n��.�.�ω��*�,�zl��0�x*�7o]�����#-�j��E��ta=ܙ�m_L��黵�)�E�Ŕ9!�!|�O�٢�9��V�/����6r���s.&⮨ݞ!ud�ԷR�d��g62�u�2w�I�ժx�S���hӃ&hX�0�m���r��[Q���^��r����ۮuU�}U�s�����8��z7�3w$�H�M��H]K+F�6z��۠��
�����<��#T��Ig�r��M���W��%{v���,{�����YZڭ��<-e�v:���E��ِ�B�t��XE�sj�����\��v��ɚ����c=j\�TndA"+�<Hb�s�����Ξ���B$#����މ��_wwv�W&g=��b2��W{��=Grﺐ��δ*;-ԝ��;m��{�t���TXs7�N��+WǨ�|��CӫV�c���0.��.�/Df>�1}����.��v�Ζ+�h'/�M�+nͻU�ը!�Z���nM3Y��K�#wre�����T3�\īig����![9���K'q�1�ӼQ�s�q�t}.��ɴDj�B%���z�g%Kw����e��|��������+�Y��Z����5�f��]4/������w�<�YsUk�t=̨��T���PR��ց�7Y���m�)�Phv������=��_u�ʅ
]�[�i�j�Q�%d�P��q��e�����ˈn 2o���
Ӿ
�1����)��(���w�c���hSekK���^��wCd�3�E�%]�n� �������a��5*�r�=����ɂ�q�	d˄�7�%��}����4��eP�of.�l�=tֽ��+5)p]�u��qg*���	��rXxujF�{���9�D�*ZbrNV�,�Q!��(�'6��6����㮴뮺�N��:뮶�8�8���6�*�B��Ig~����蓠���GUQ����q��Ǐ���뮺뮽�뭺뮶�8�Ǎ>��C�%~����l�U:�**�I����QA���L�浻~u�_:Ӯ�뮺�뮶뮺ۻ���v�������"*LV�d����I�ԃ��Ǻ���e�HB�P�v�M������X뮺뮽�뭺뮺�8�ǌ{>l�Ȅi��[˹*g�l+M���pЕ���U��e�6r�UD_(��g����XO\YE]��zd�W,��8<w��V=t��̪�AT\x���D��!��a��d]D+6_Q�)�ĕby���^�eA:$Tw���Xs���Ǖ�B����,�y@�M"�e�2����'��9/>�z����Gj��T����N���1(�P�brD�j-m;\+UU H�����uV�%U��D��P� �)��B#&��叅���航�,3��}&c��/�q�����ݜj070u:�:�[Z-!}���X�2�+�%�0Q)�SWF������T��1�"��""vH�b�$�T�"������ª�����[��)�70f0��J#��%hj7"�"���GlN�#wA"j6�6��«d�I��48�d��U��R5]Ӆ��z�F	������:ȇ��&�L�X����T:KTHvXi�HX�B��4���j9-����Zi���i����\���o��-���.7�-l�gq9��g
�҂�Ȗ�M`���Ӭ@��Oz���C�IO��7J������T�g��3^�D�C00(d���x���|��y\3���dz�/N���^�7�.oѸ  ^��|�EX�����_&}��K�y�n�G��b�-���@�����n'�sk2��]�oT���/C�̓�od5QQ.@����>t;���QGoOm�ut8�b؅}��h�@'�����Z.�TK��z�F�(ݾcv�Ga�c��Ҷ1��ĳ{���@K�C��=NU֕���_�j�����͔���}]m��;[ȷ�Uq�:2G��2T���t�tb[Ư`��Rg=���o�;Gh�3̺�=��b�9�XU
��)ԫI�-l�\�4e�;H��`���B3!a���Nm�ԗ���R=7^��V"�3�>�#7s׷ ��@Ύݖ��2z`��W�.b��kչ�Z�d�.����:��M�|�Q�UO8����M�xSz�ǁl=��U0�L�f��1 �3v9�}��ևsw����r\��\][}Ԥ������D��x��m���i�����=�s�7���!���`����v)����M�����V`n��d�E��,�c͞��_�z'��oi���͋��}̔e�%#�N�e��r"!�"�w�m������G� {�pːR=@�����|����±�F�7�ۺ:h�]�����mO����ɘr����d�5d���7oG��q�ff����ϯd�ǰl��}���|4��+�x��uy��B� �ݫTgo"��h���־��֮Y�j/�PT���
��)����6�'�<�oWxg�1裬��� �ltV#��l�n�h��G_��+�����%����0Xnѭ��i�s��-_W$�3��y��|.�/������D֨r7x�)Ӑl�r0���W~�XGvFMD[����dz��ެ���S�|&ޭ�޷�c+(�7M�h�f��)d)�e	�w6��V��^�G{J�E`�Ok��L��w��,�gM��{=�i�]3#�-�q�t��b��[�n؇x仼���˭뻽��?}hi���hi���U�s��th�xhw���d�^��©O��wl�M3��H`��Q��1�8�a�M��.7�;��{$BƍN<zy�;�u���o�A¡�z�s�;������8p)w�@�6�Vwi�2@�+�H��a�h��x�Շ�^�b|Fן� ��Y�e#��+c6�t6�*I����k0�k]�ٝ��s�%�="����4��~m-�U�=�Ŧ��^�g���Sf{���z��0��ѷ�x�g���.�2�;�N�yGc�]}�g� ɭ��������837��f0o-@ψ\_,V��/Ʒ�'I���YL��36�+�=ݐ8���5e{_e��������Z��.����ig��٥{����]�{W�����N�C���39���By��O�t��9iF�P	6��a������_7�~�Aծ`Р[�B�軒��t{�hc�n�����r&#���d)a[�l�2e �z�J�us�%������+���wJ�w���j�cU��G�g�g�y:�~�&u���V���j���j1���i�$i���z����J�����Ʀ[=���u�|�*���L��##:�Cpק��]u�yf����r��CX�"N�30nS����H�ы��c��%�]ٳ�6)u�纆Eq�S��f��s�|���a�}��׹�}��\���jZ�xz�к�KA����w�U��9���ϯ���\]j�yⱃS�sO2�l���&N�j�@���6��lGh�-�/�ܕ2���n�&��j`��вs,�C��׾�a��S ��>Է�t���Tj��
f�ɋ:���U�Jxz�y����4�<�rLC��g��Ǡ �<kͳ� ���v���-���M��HU����Xّ��ٽ;3������N�t�7	�ŒQ�>TF�6Q��6=oO��FߤB�ff��a��SQɾ5�h�>m��D߱�b�>��� l��g��:;y���گ����Uh�:�k�^��,r�7c��U�y���΍n�ç�OX��gWLUcecT�y�|�䴀0��UރӘ�L��Mgqw w�v7����v���9��﯎S��6'��^�u�{�߶��Q��4��M5���w]��r���m�I^h��s�fNI�Z�ܱ[
P�t|��#*|6�)�@���3�t��r�&T�)�h���$;d��M@}��U����#*���5�/ט;�;�؀�6{1e�B��["%33cO��`7�W�f�A��i��%�:k.b���$����Gz�zڱ�Uݙ�8��K-�禮�8����8k��ڌ���Vq]���}e�8�k"n�*�D�5d<����E��_�������.�W���^����+� ���g�����[lkc�f�O�l�v:8)�`�j�#��8�i<o�N{�c'�_��T^�j��kK��R��u.zhf�p��6duD���W��Fg�K����ו������ξ����g"��،5OL%�z�`�;`?4?o���" QS�ko,ť���T�=D���x�)�zT?(E�	��P2�\�.�-v�byUΓAd���{vz{,�a���Bn�#��w�j��}SC5U����/i��Ri�^�q��>��E��~D�l����q�5�x�T��ޮ7[:H�;����_��=Yd���E�wg�9�q�����_[CM44�CM4�L�y���������|�~��d�{��š������"#^��|�����峦^e=>:}\�-m����S�����>3藗�|x�7��Dih��f�or�������#uG�l�����T������W����uggwy�a^��n  sż��Z(��)a�\�{0�<�#"��h�� �n��sȤQo0��#������X��^��j������nܤ��a��(����9y�׺�C���9]ކ��b��=;�H���/m�U�Ue�o4�KӇf��������t���H��}���O˭�;[����5�;��z���O�E˳Q\-1����6)��gl�F���2*�{_t+ ���lY#��u�t%�"\;;�J�rͤu�AJlO�<�xw,���A��ʝ�0�{ܖ���;�-ݨ�F��Ype�uSKj^t�7 .}e��<F�u\YZf�ŷ�^�=-4�.e
����9��7�՛]����@⳧������ƪ��,�U�Gcw�|v.Á�E�h��W�CM44�MF4���s�w�ｕ%hxV�f&���(ߡ��I/s��*ÞP�%B�0�97��޿N���F8��?�Bf�՞����vf�͒���_oee"�+��u�7�,oe�
qA(�IH�����S��`�f���b�0�7�sU�Z�n*i�
s�nC����f�yn����´��g�i�q1 ��L��.[�M'��*�pk˕�T0N�tI�"�w����{�m���W\������V��3:2��.�*h��3~1}��܏L{ iJ}��"X �JJ����n�&B���'���y����4OB;�c��0�b*����(�>ٯvg�N!��)l��w{�8�C3���� %���*�}��w&�3U];qm�s���2Ӷ�STV*[�@B˔��ԩ����[���=��m{�g��}���dl���x����i�
�sxn���g����QG\>ä[�ܶ�	�]�|����Z�ۢ[i+Mh����U���*Q[{�������,�}'^찬0vk�D�إ\-��)�O�]��{��ו��{�V_��H�m4��K�T~�m|w�7�_�s�:�P�s3r2�j|#̵$.'q��
F��Ko]�m�}���w4s���o������IQc?D䟫�(TV	߾3x�UKz=r+z�� ff�q�L��;/L��8��0��Q�I�q�;є]�7HiYϙ��a��x6���^ި���L3�Hi�뭝�dvE�7pwV����d^r�>z�f��}��_���qy���a����^�ȷ�cbB���k@�$�8=O�5��6��°o���f�L4F�o��F�z����:���G�+M3��U����rG4��f͡Q��ӻp<x��}����
��{f:���$_/tE�0�윙�㞞}�I�d������8n*`ȣ>�c��7��7�e+����ztg��ǔ\z�%쾎�����t@O��D@Α�p���R#L�T��6�WY�.}�#B�S��o�wK:�]�n�w}~}+O��Tv����]m;�:�#��� ��4{�U���ě�zμ���*	�u�:�RԾV�S0��}��4hZ4hZ4h��b<�|���9ǔS;��Ɛ}[ؙ�ɠ��3'vڡD.�;�r[����sw��"�]]��[C��G�0S���y}�N�Q�@Z��+d���~�hff\��uQ�弯V�#u���(�/kJ�&��^��ʯ ��1��8�Q9A�"���ׅj�9)M���Lz�7{u��5�|�=O����T��������\a.�l�;���6�wt���������[;)�U�s��k"�%��zvJ����Y�<����7�of�T0��[3�ʏ`O���j�Ϟ!����M�:��6�����!&�����[@{2v2��Y6t�xǚ�]cw;��X2���7�d�݂��g٪�ptCcuŷe���ޡ��Y>�~�L���F�yX���̴���sd��[I��x`�՚p�0�^\��𽧄������Y;�t���Z�r�qYѝ�3C��N@Á�fI�Pa�Dh���|�Aיy�Z�4�Ɖ�8��rX�=����M���û�ʚ�u�z�a��W�rd2r΃��&��>{P��}��5�
��f���\�0���#�b2u"^\�͓3�|oXm��{�	���,��h���CM44�@SM>_}u�w���6�~��*kd���i���F�33'x��F�OT�MvQ�F��U쇹�D�z�������R��<�H�X�ǊN�������;����A(}�}�l,���-���#z	a��gj��t��w�����U�]��9�W]Wܷ�3��uLG�*�3�5ݏ=F 7z&�b��(���.T�p��������H^ˏt��̰�&9u�B*�Va8��rE��'�g���h��w���+��^�a�մ��Uf_R�YD]AE4U27�	�N�n�����l�vony4��6	�40P��1�c/VQ{h36?�B�|��,���t��#7H�imX�O��ϬױvRF�;0���wp����Cߵ+� Evת�t���g+�N��ـ��;F�D�V_����<x��Ϙ�T#�w�g����a��W�Ƚ��>�B�Pg�_u���R�u�ʜ��H���K�Rg�ڹ{K�.�]�n�񍷺�lMik5� �[�H�3/Z �<xp���35`te�9næ"¯D=y�E]tx�Un�+��I dRqJʩW�i��(,�]�l���Ys��B��㢱�k=l�S�v�h&L9k;��J�b�ґ,�G���ٴ�/�,#�u��_��]
���i%s.��\��[��-ܮfNg2����8��Νؕ Ij�^�`�ȴ���U)�Yڶ���t�.6�j\���#���T�'>��nݣ:�}O�hН�k
��x�3NV��-������7m���3�=�8�)�3h]f�J��j�S�
V&�3�g=��p̘�N��]�:�ի��+%m�ls�Y#V�n�?W`x1+瘪ÌF��Y�k32��C{%;�6+�o+f�]w�'�j�r���*|j�Žα�\(�)]m��/N1hu:z`�����<Wy}\7�n��e 儑��
Y�a �vݳ��Q��L��%X�� زS�����ruGKm�ΔY�Е��W�:XF a�uMN��F�2!w;5�9X0�5�1��@(�] Qd�p�G��>�Y�`��.����$����E�d5u���,��i�u�+���Wgs�{*��_�ekwl���XY�2y������MUdDe�	�D��"4V���!��qm
�'ݳ��yϥ�_q�N�V��&U��k�ӱ�i�{�Q�:���}��J�q��\\��&��ln]��]�t᱓7�����v����K��0��]4xM$p��g5Cms�Y�x��3v]�sk(�v'sU+���w��X0�6:�eww���r����XM�.`�)�0��܈��T�ۤ�Q+�ۛO�����e�8�J�o8oDQ�l��,�����o�@HB�GOi����z��EJ��MR����lb5X�s��Q��g���V`�\C��]�G_
����|R��Q{��c�鄽�=���:I�m`�6��Kȳ1��ĺ���o:ݰ"�8�L(c#�*��p�F�3�)o*���� �.\&�Y��ʶ��\:�$�\�E����#�{]&վŇl�i.w�;FA���af:#�`����]Bgi�MhX��絹i����#��v��vި�6�\���u�Sk�m��ǻ���I��dq-C"��vv��9��t��uB�<���:r��*.O�Qk�.��n�<}}}u��뮺�ۮ�ۮ��8�<xǿ'�S�L�T>ޞ"'�����Jej���Ps"��������<u��:뮺�n��n�뮸�8�����B�)�L`D��@��b�U��r��T�=<i�<x����:뮺뮾:�N�뮸�8�ǳ�ڪ�P�=��f�+**��U����I]	'OM6�����ǎ��뮺믎�Ӯ��8�:���9^ޟ�~v��'�*�_�UA���H�p����p���� ��P�r��܂$�y7$&QW(���Q(Ό�PD}�t�3QVRF-����m��(��B��!LI��ΕSHB�8UY'#������zw�K�� �i�APDp��H׏8E)>��A[�)Ɔx�����i�]1o)�'�AM���K����:��'��#��]��Q?{=^C���yyy?��=����&��rÈw�y�`�M899>5��,���������w�hÃ�F���xk���É�je��wn��=4}a��ը�w�6�mxȕ�VF"y"�e��װ�M���L>w���xBK�Ґ�ʫ��S�]ެ�l�G3t[��*��9W�|��g��4���#��Ԙ����<�˻n���G@��15*�x����/L��� �î�#;�
�O	�z�B���w*� תh�P��3�*�y��lm��y��+��:�^����V6ǩ�{�b���>M@\yML��ܷ�;Յe^�'9�eV�Ӫ^k��Wa�ɬRHc:��rwM�gf��፡��w��Fਜ਼�����e@4��lh�D��E��Y��R�'�ί�/}��96�R]*�����L������L�������":����!��5v�2*̮��<M�F���>M�}d�O��=��՛N���>�"	�]��Ӛ�%��:������~t�YaN={�/8�Z��]�u�]���Y�[��%|��CM44�HSM/�]�Q�q��x��fG�����
;��yL[��n�ݹ��ƹbw�+
D���ou�8�!���ڢk�f�)3�N���ɻ3'�W��0%��k���OA(p 5���� �|Ty���:o��-����6i,�(R���`ĭ��6ڽ���g�;[��z驦�F{ޙ���$����+����{����3�()�������y��Qra�nMn��x�o?t�%C:i��Wvs��魁�3Z/)�ƺ>W>��X��5�Mz�*�$ �å�dT����W��3��<Mv	�s�����1~�]Va�n�2�.������:���ݶ*�W��Лz���J8�9<�(�Մf�����V��0<�\;34
�>����ɥ��	��a>���k}cr�g~V�����(~_=+��$���'���n��J�xM\�fS`���/R{�ש ιY�e�l4r�yZ*u��`��b�՟/�9�^�	_T�bS����4[�۸XS���w<f�Q_KWQnl�֓y�(���M-4��M4�~}�l�}�9٨,�ޭ�h��Rh���ܩ�zN��eP��}�jվ�F����@L�:�<�>�����o�#E��U��V�!ٞ'���,�Q�X$�����m��0Qc������;��7Iv�O����fyu@�G�lѓ��f����+�:+
ӊ�"U��!�ײ��M����{�^J�s�f�=Y1\Ҥ:N��-��w��#�k.���Q���z��r]�J���C
���#.yQ�K 9��y���Gi}�.y������ċ��6"D^)z�:;���`��'�ŒS��\w�ґ��ƀF�|�o�\���aکh��f�&/�ś�H��B�<��g�����k�f=�pmk�֌;=�H���<en�.��g4��m`@�Δӛ5�x�fffa��b���`��k�7�C��)�U�6X�C[vXw�Z��]�Q>`��{��X�O��O6+|�7��g�J�%x5~�^�,��z��[Z9�����Wη"�o�ܺ�z̵u:���k�iq�ؾ��)y�����QDa	>
�q�&mZm�7u���Of�X����"`#A]����u�[Z�<͗�����X����{<����<�8����ݼ̹%l����|��k��Û�r]]��m��]`��m��M��Th���$#����l!��_WP�Ɉ�C���2o�,�l����'U�C��.x�W,��zιE�昜W\vM���v�eet]3�*7��K�`ϧ �}�`ny�n�U�U���#����|��^�U����;� =:��C�P�,!X�pk�bǍ�~b�S�o{Xxz����$i�R�fϞ�z�(.7=Ր*3s�X�h�T�w��s6��xvz3�*m�P9����" ���a`�Y�c\=�a}��*�����AS�\�k��曇�ܻA��	��6�ڪ�nIL.}��Ғ�sʙƆ�n=��I�����9vLgn�qy��Z��ƫݏ^���H篗uhm���~��+�_x���k	������<xؤ��E[�Ս�֬�#�����yY�a���f�U���t�3R�Mvv��h'�u�Uk�kj>�R���s�k�衯��42���FI�^*�5�͔�R�K�����>�4�KM44�I�^���O�fb^0�F�dR�M�33N���4H��.�F����l�~717B!R��QhV�S\��l�W���[�ټ��2��Δ#��*�;Q�nXI������Ⱦ鑹��)=ϧ��~Q�Y����L�Q+��G۲�mכ����j�M��,@��-W֛c��6�[�����G6z�����}fO�up5�#9�\*�\���t����]�ʙ����ߣ���w>�8׶%yj�vxq�]�[�M�9^�>f�)�$�0G������M�e�5��ݵ�I�&��
�*E�w��?�����l��c��sE�?�.��s���[B�`������ߊ���xhG\�g���0�ǋ>G�7�E�yVf�ޚ��Dn��	{n$�{ hN�\���r�����?k�E�xu�굸i��i�B�pO;�΍��X�U�sFm���AӉڐ��*t����i/�����@��ߧ�.��3v�N8��/�ֶ-��uz ��3�vƲդ��W�e�N�c���Y:���ֆ�i�#m�4�Jw\��v���=:�����uK�g)�W�0�lt+��G�E�dg$oa�P�o0�"z��8��m�@��C����щ��c�j��ݾ�"C6Øq����Ϋ�z���`0l9��U�+j�@�:5ms���Ck3��$��#��f1�{XM�lwO�}���G��%�y�o��x/���e�A�Z�[֠�T=������v�:e�y�L��O�y9f�|���wî7�R,C�,��*�G��?��v��0+yX�c|1e���̝"X��fgݥW����#�܌ �A��{�ʌ�{.u�ܛ݅m7�6�
)O��o+�
[��o���syDb�٦���b5D&����˞)Ux��e(��y�(|A����'�X��{�#.+d˫�=~��'v�H�_A�򽓹~�ͪ���Qo-�ݡe�v�nn]���ъIp˰z���]�lk�٠�{� �	#D"C��s;"}IUr���޾�{�=v�ԮT���r�>J��;Y��ݐ�O=zֺw�k�y�Z.Ƌ���ֆ�hi���i
�:�6��(��Vٍ���1�=�p+�]ٽ3Ҷ��t׻�g�V9}.�Xa�ag��1s8�"�/ru��I����>Q�
��,#��Һ�%�38N�̌��ޖ*S��l���d������v�y�=tb�<#�1�r�g�xwͫա�<;Ъ������9��%2=o5�ެ�	OKMf�޹���0�f2��F_�Í�#���Ȩ�{�h�r�����j��"\DE��/Y���!�Bff���I{�o]O����,����r��UQ���l0�>���ff��[�b@���d�ۊ�ro�ʌو��Ȭ�HZǬ?��?(�1Hoz6���&���s��q�4'7d�8���S���} (���~��@��w�W��|�T޺���fp�[�����.��Tѹuz�,*Wt�'�ٽ5)�,ϳ�8zy	`�T��� �(���Y��p nO���~�x���Շ�;�	�՗���@����k�.:͑�ֹ��!qZw��xl����&���y�d��
�P�U���j\��V���3�W�`<Ni�c��io2�w79�T1Ig_,;ˡϟ\hi���iJi��y��;�����y�L�7�����W�gy��,�����X6Þ"vt�����3f�'�d��Lz���.n�����c_ygLf�q+&���;;g��,��;�N}�o�vzn�Jm_.�{�g�U�c�I�j� U�|{��fK&'�Z�mG�Xg*;��R\6��{�ʺ=�[ֆ�㾮>��g���@Ηq)�3�u}YZ�{q�������WA4������(�L$�j��ƭ����~�;�[�p���^F���x���}4��0.�Oy��+��333�D���+z�B~���G��jL��(O�mSag�˧UΣ�skT�ޫ�'�kxc6^��#J/�}Xs�W54�w�Z���I@`�E�V����fr������t1� )AU�];����zn��E3��q;=��5Z�w+t۵L���kL�ةгd|�Osk �V[F/���LU<����g	��]�\Rɼ̙$'p���k��Fw8��B�+���X�C5y|����eT�O������//!���<����>�O��j�$�Y��u����=�l�مPJ��z�e��CCVSL-Yq5k�/Vmez��Q�1/޺�q����ƻ��x�y5I�g{4м�=��7���V�}��M�㙂�wm�O?{ƞ�� +�ksN��{��2�N�2ʽ� 좒����R��i0�|r������o;r�8����t@I���ߟӎk��_t��ɿSM6�OD���ޘҳQ�d�����ʼ���j�8{�GJ[����Y:�Ѭ�M7p1<��Pں`�m��樮}��e}�s��Q��or�͆wm�׌�is0C� �;�Gv�͏�׺��Z�b�K���x�5��u�� ��l�33uEm�g�+�=DG��.t�w���\t�ڵApy�C^����1���A�8[�&��EU�P���o5~�l+}B��cvr��T4C���k�"k�T����(YewԪ��w�Z�U��nr2���዁�Qӹ^t)۽�8>���ڥ�<��A݉!��8e���w]Vy����/���KM44�CM4����u�6�|���ף�r/����� >���U���u�+7�Aoc���X�gڿtO��@��}O X
�ض=��^o����4�_��n��^�n�N��1v�:��iK
�����!Iza�LMI�a'��SYfy.���9����:&��Y�OCoڂ�5�eC��P�:��ƽk����*����:O;d��o�=K�<��)���l��DCzs���Pֹ�	��sBH%Jګ5��b�`<Y {&�;�������N�_Xv��)��K����{�W��O,���c-��v#�p�F�R�{��"�޳0�4P�;巓�|zz= ��2p�A�yH�&��g�+y��=�E	�z��#�e7��rt���'���-/h*���#��zϸ+j��ݞ���|�ޡ��vUq��)���R��説�29�e�[��-���*�1�	��ع>�p��CuT�S�	��O:#H+t�w�z�rHM�)��������.�9�H�Z'�u�gC,�Zy\�$tU�:'n#;G0�R���&���+������,M˼���2Y�Ig{or3:��rqv6�ɫOe���k�m�̊�N{�üT%��@�I�e�|y��o�թZ�ֹۨ���K�u���A;��5��!|��"�����������Sf[�3�*b��Х������yF�Waݛ�tz��È�-P��;�b�`X�mx��S<��z^�<��tL�Wz,_MU����'��n������êZ=�P����y8��o��;���`�a�ݷ��L�/]�'���QGy�l#p�J��px�ei�Q�1�V<77�'�WU|�EN�6/��v��uO�_#$WҹW<x:�o׹jw2�w2z���sR)j�w.Z�ic�<^=�W������)!��u��������W)O3� ��
Sr�-
���:��k�N.�PoS��];.C�b��F�QDՊH�Y�������(f�Wag�+�.� ۣ,�1Q�$�_<5-�ٹ�'bu>#�wւ��2(��Z�v^�=V�B�P�H�Sm���1�X&\�Wf�L�����t+�)�6��H�ݏ��0������Z��tw�M��>��������\���]�@S]ӵH;���Y]���M��;�h��4r�:�p���T���w�y��(�ع�Մ����j �M�h�}�,0�7�溛���ûݣ.k��֎�W�����jY����=��9n��r��mh��}l�*�۵Pv��w:q\���z�
�p��Jn���NX��,�(p�z�]`'mB�R��o[���Ip9�s+&���د���2R+�Q��o���۰��e�w��7qYKm�89Sv��i�� U|�����`��p���][���r6�sMie�tiu<ƨ*@�lT8c/V�!u�'!u��m�����sw��l@ؔ��X\��F�l
��R���m���f(6�)�u:A@��֦�חj���`�K�S�[����f���F�.i�/�l���^q�(��}p�|q�j�a�l<��o�����1V:v]pt�_!o�o�i�VU�&����0ۉ��r���'7a�s]ۼ�M�Ν604�:���|�v�ޞOn���UqL�@�EU���+Y72Sn嶂1ky��`$�A�UG�!p�>�?0��@g*���I'��<q�u���G]u�]u��]i�]u�q�x��d]�}���yp�8B��T�E�x�2�ƞ�x���ǎ��뮺믎�Ӯ��8�:�w�y)Ȣ(�Q�+A�9��.wS]R��M�:믮�tu�]u�]|u֝u�]q�qק�;�BH}�*��W���ˑc)��=WmǏ<u㣮�뮺믮��]u�q����d�B����*����D�V\�]��p�C�G�u ���3����~���J�N�2�ЕfM'��***�_l9ۥSĲ��<��F~����K����)�T����8ETEE�9�D�Zw�^��tYw�H�dN�Qp���U�+��xCzM�ڽ����Z�����#R!
��u+r��ɠ�;[�f�m��bqى�@�U*�V�ej�D*��
�б��twT�rO3��>=/4�,P)�L��z�Si�3��ډ�p���us}R���1�t��t�s%���aַ��=���W͇Z)�I4�`I�H�V��z�R�t�cD��6�R�XӒ'c�I������5),��,X�!��,T���ӡD܄UV媤5^�Edn����T]M@J�":W�]4�(1��[�R�*SV"����+l�"�\S+"�q:T)S����!a+��R+mphV&�M5jr&ڑ�]�������Q#ӪGeQXA~���F�/yyy///+#�X����h},U�!�ԙ�w<6�:w��A�Sv-�°tw��쇐w`r�����c����Т����SMڛ�軿�����ކ�b�u�]pln"}�کX轍�w�7t�{�5m���5a�\}�]��^电n3�{@>,�����g��λ��38��ޝ=��a�=�f������ٿQ��NR��ڻq
v�(=%���U�w��>˴}+_�<��m�U�ݍ2��[I��2�ޚq)ܡ=M\��l�=l+L-,ի�*�����m	@zL���J�
�W=׭p��d]&�,�vMN�-=���=���� sF�wM�]I��:EJ��їݹ��t����m����s~x���`W4��n"M�sV�ܑZ��3ޡbWB�m@t�����I
[b$]��3y����y���D�5��{��gWW^�h�H�ʳ��6DH�n��w�l�mx[tI#��SG��Zޫ�@+��8�;�'۠AL���6DfT��6���}qN�7^+��]�$akڟ�VU��f[�ܣ!]ոF2�Xzv�Ң�W�fC�Ió3Ws{n�HC����a辏D��u:P�Y���5���]��뮻�y��l�>�����b��esu�8��4���x�����{���z�|�&�:���U�˺H�ݲ���W�c�[!�ΪDSg3<x
��[����ʫ��5۲{sr1)�|����hi�]�:�Zə�)�=���`�@[�r2<T\{����9��z��Doz{+FHU?�2��a�H{"!����YzMz��Q8�yt�v/�K�����^mn3K����D(̍ԉ�^���W�1L�_Q�>\[�Ĝ�>yN�Ϭq��芈��<g.<Tw���!���>�osC�.��=[�#7�n�M=�*������kt��-�W���oVG[⌾HEw}S7r��R�=s��rv� ��	�{c��[�N�q%w=�f��v��k����;3o�W�p��+��ۖ����M�(7V������llL�� ֦���ʘ���7Y���<}�����&H]�h,�ٜ$k�^i׬i�N�>��X�bD~�,�@���g#���K92�������CT v���N�Y���/�.Գ���Q_S�/��{M�U|�Ō��@�̞u��UU3�gv򍰀� ���`�>%��`l���ռO�;��Q���{V�t)�f&���'����F�ʚ�����ڈ���B�!�G��ۚ�ES��$a����#���K�������9VU�t�x�P�`z�/~�smӎ�5NHR6���>��m���q���C;��;Ҷ�\�/'���'�fh�C��ʆm��12���˺��Ӓ+��g������2�f�o�썀�Ǣ���M���4��wpp!r��>�i#�������nb��g�f�i�~�u�t֔g��!J�gs�D�X�{|�[-t��gD�Tt�ɇ����3��7y�G���������r{������B��eQ]9G��6=>�P���733%�*�
/�g���˷b�7���	��)�}"u`٧��[��6�����דٷ6�����}{}�˖3���h�$jP��J����:��ʬ�>8���2%ҁ�������;�-ʾ��Ҳ�p�"��.�t�M�gQ(�Z�W[��.��F�UMWyy����7��o0���mZ+L�{�K����l2��oG�}��z��Z4癎ĭ�s��zs��R��� �_�1�mC���-h�9�Ѵ�:Ք�q�PeF���yN�W�u����V��ŷͥ��E��Ut��Μ�$y�X�<�}��[��Y&���G�Eu����%d�����ux�L��j�\�r36	q�m+�̍�{�e�^��r�晆]1玥Q>����g.��q��>>�w�$L�R���5�Iw؆��}i�77��!��p��>��Nx ��2mn�k�g�N�|��d]���;�����&+nS��g���B������S�<���9#^��'��{v���l��C�����Gc��nn���5�d"=D�j�U�[w@D��G���VӬ���ё<��e��CR��/L��?�ג�U����d�⒏�w*
�g��̚�2�A�"G/�jK��2u�]��=�9Z+_u*q��чz�}�T�=��o��x���D��0��T���M��y�+��� ����J��I��%4�s�w����~o#v�-�,<�ly�k#,���]��0�P��S|������8{�ްRw�ގͮ�`ۛ"����@Q���ٶ�֦��P]���-��4���Uܬ�ʖ���-l��]�(��ܻN;��UF	'��ﻣ.*�ԍg
�*w����um�Ouy[�<"t��W]����P�՚�|	�,���H�~�a����b��q����T��7��sxy�ι(ӶUUHlx�ia:��%\�*Vu%������;w�=�er�
��T�;��y̜�%���.���SL{�%��Wػ����k��}������F�-V�Gmb�C�Lɜ]��M�d�gg`��5�8���:L��NJ�)���qV�1αta[��W)��܌�O-��I�_[��5L��iT�Vn����5���1y����ϳ��vR�'�p���@mR�����J��*�=�c��=# 5�[ bf��3j����`�l:�ؓU�=�Ԭ�h��xf;Ϙ�8�P�siؕu���v�x�EShJ�Нr/V���s��w��
x����<t��Gb�)���)m-�}O�N�H�8���D_k�4(9;y�2�T�r+��Je�]d�w|��u{�7��T|�0c���L�Y%b[>�V{۠�� ���@�7;�#���n�J4�X����D�Im�ͯH�熦���#W��߱>K��g.giۺQ����$�Ȑ�u�WQ��'yU�|�)�^%����n�n�0���kkrw
pj�_���T��3V�3sP�I�M�w�E�c�tS�u=RsUq�FT0��CB��v�?7_]]��mT�ΗP�ʘX��/z�2v�}�oL��꟔�m5����˻?uʣrI��vj,���ʍ��@]�U���N�H6�)���ۋ��z�x4��]�&�8@ ��1���k�m�WQG�7�ݽ�o��0oph��죳������EN�ǞՏٺ���eͦ�36�K��RQ-5W�ƀ"��O����Q9"�'���Kt	��Pѣ��d6a�_��;K�	�������&�+�hn�U�;ߣ�_q�K�����_Z�������>�#���� �B���3�%��g'i6�
��u���Dr��*%ٛV�ڵnNw��3��ﾯ�<��']�D����ŌP�7޷��³t��" �w�q�c��a��D-��3��7|�	��)��n6�k	�݅�}Oc|�{V�;��9����o]^.��)��wX�+�ݣ������,[^`��;�_<��݈���3�њ\kf���}=��XMAH�X/�X��O^g��z���^�Ә�w}j��|,\�^o_��HĒX�ZM�9�tK��ü����օ��a;�]�u-Aٙ���	Ѿ�Q�wA�7��du_��84c�+��x��S���V������Z�m����u�Y��͍���*�C��/ù��Pn���k��ݺ��$ŕ�N�C�üL����V����+*���p���c�}˞�޹[툺٤��"��m*�=!�+Խ���@� �gRo��c��4/|i?ܸ���Γ��F���q|�w�N��HP/g�e5F�wN�^o�\�3Z^�"�ap�b�x��-��p^�n���Ѐ���Vl���p������wu������w��w�l���1�1�!^��p�Fk�+�jk�_ *\��w�ÑM��}�n����\pY=�vI"*uto��!��2�u㪼L�Z���׻�-.�f}�|hߟ龞���+��u��=y�0��)|mr�6^ueGaD�-4d3��L�G8Dd:qĪ�>�8rk�&�M@���Q�>:��8Sp�V�k�a|o�m�t�m��W=]\Ѓx �=���{��Z���|��{��Y��4�7֘��w.3�%����:V�!����So\����d�4�NH���y��H��gȈ�\�����އq;��d=���0�u�d �nn$`Q�PM��܌]�$p6H]A�ԁ�*E�[������c$���v�.$��O�"�'�Նf�����3���O���m=��>�`��n(ެ���gA�g}N����>#����*[y��o{)nZ`/��V�����d�#�f����֚�MM{č$�K���;�vR�<��&��*�du����+���V=pa�Њ����iۢ�M���|���X��A��������}�EVɣ^�)
k!9���;�ْ��2�}:>�"�5�kN�{Z�V;�N���eZ�U4]�u}�򛂪��'����Ҷ��QH�\������)��8���h�)�Vr��޺Y�U�@�0XeD���`&���T��h�xnw��7d���P��fv�F�i�#v��Y�]G���:�q�:�tڢ��1A� ]q�N�3A�P�걺�mU�M:C�k)RCw�.��z�3Y�8�f�8���B�ߟuku�s8fj��(�ojΟY/
*5S<{\�ew�x�F.P�`M3��+���i@�{gSerbZ&H�zŹ�4����kz���n�H�2�X��Fz9z:kiޖE��S���2�]�8�l���L��v�p"=o���K=1u���'u�#	��M�2g9#l��}���hd�zw[a������;��ܞ�&���[�6��'�װ_w+�Я�)N�� u��ڕ �?1G1�UӖ�������ѓ5-�	e��+Cu��[��fj4����0m��r��:r���o���uc�xw�Jh��5�кC�S��fa�h2J������x����7��te���7�ߘs���t�(�����Jl2.Y���l��z��`���5f��~��|��9�������//e��q��qqP�j�.��2rFF{$o3��f���c��#f+e��eGVl��ao�V�Vs�W�o!t�"3l�0�hH�g��9�?Q���sf�(雹�ނV׻ϜUzFgD��$m���.[`u�
�HC����7"�.�n��z+�v�yez<����WY����t�#U�Jf�rg��֧`Cw�J���Y�P��7�����F�-�{
�M�<���תּ�g^Aly������ {ˊ���b�{�Fݬ�'s=]Ю=Q/��x}B 5�{����*�P]�s�f�{x__���*w@^��[]�̪�r���s���� ~V|Л�ޡR�4{kFt�@R�D�y.��e [�[o'mά�oi�	���P��'�����^s���m��f��M�^y`�'vq:��������ž�EYX��2�ؘ�(P<��fY:�XC �.�Dg��i��o��*ݓG-O��Y��(�\���c�r�㙷F�';i����R���&�RX;��1m��l�SfB���r�h=Y��	}�	�NM��*�{����L��&\	_1|����U\����M��n#�4]�{�ru}�E�ݬ�j�A�æ����5�'����޾���-�жr��sc�]\���p��)�*G������OD1�,�Wf=��#���1U�%e�7.��vV�}*�e�QX��V%t�jЗW��{D&����׵<ͺ�z#4^@s�]�v�������K�{��5����+�K�&��y��-�F��[���XUj6�`�����0>��P���5"�S��q�X��>\��a�qi{��T�3�=���#��c�i���C²Vt�b��LɊ�;ݱ��Cw��t���i���m�%n�y(�u��1����a�6�-q���n�ln��Y��P�(zU�d��1���C��H��U��;c*_��@���Z�:��bE�нU�+b���6�l�k� Bt	���ILz���/ʭ*�CI���sMܳ�����9]��ۡ�헋Y��z˴,�ꈒs;w�u H���;'' ��R�U�y
�=���Ω�3���ۧ���Ëw�^d,ry�'��^�S=^�px��"L���ʒ����gjy�����g��d���ʾJ7,N��ѭY6�؜��v�����9ڮ���rꝜ��q�=���.Ez�]ʈ��G�����D��<�0v���aj��+_U��������ы����pK��.��M�k�rG�d�g�Vj@��o����tG.���o]��������^,�bQ��Z���;f��uUCa�[�Ԭ�;�7��L\P�1���2�����=�	��Z
I}�Vf^T�.��Zu������Lw�d�y�R����IE7��9�+�fVQ1M�D�S��Ա\o0^�CP+E���j#w��m�t�Š��]Q�|��u�Ō<3�5L]
줈;6��	��͎sݾw3 ��q�ok��wX5�{�#��Gq�,Uכ�D�t��]��}�]�Z&��7l�kkq�i5��i�7N�:�~Gޝ��_8��\��(EȲIr�]ܟ�ۏ:�u�]u�]}u��뮸�8��rHFB+�!"�{��G��s�p���$�'cM�>:��Ǐ]u�]u�_]c���8�:�x{ARA�eU]KΝ��H����I=Rz�����n�o{����ǃ��뮺믮��]u�q�z��T��P5G.�F��ف]��q���4����1�8��㯮�x:뮺뮺룮��8�:�� �<����#��&��Yt�>�]g ���p#��e7������Ǌ�J��/�
u*!��e�JI+��2zO|W/ݎ� ��w8��Т�BQ>V�[��q'�;��D:q�dr��+��>8��hY=z����!�]ѕ���%�ʞ��$�0�x��a��P�j�s˾�>�����+�H�ۗ�U�Y�Q^��/�#��V��c��:��V_v]o%ȸJ����v^H���F���.h��x�3��+���(���,`�"�y��|�}�=�eʕur�>
7qwH�w=ۍ��Ci~f�~�(�W�,�f�V��MwMo�.�xz�6�O�=(і�x�%�F���}x}W�yل�>��t��"1�w�ӏ^Y��ݹ����>�E�5F��㋲D�M����5 <v���䗍��f��7�w*�58|Fa��=�-��6Ǹ� ��r��޴�:<���[��st�{�H�YYQ'ƃ�8��a�a����q]��D�2r��6kQ�@�w��G26/uVO��Ƿ���F¬��
�-�-.�+mf��f*Ù���w��8��)��aja�=Ox�kA�ܼC��q>�(�5Q����L3̏��t$�.p'�����"��"�j��d>���3xǮ ��ݾ���z&"#٢���6�v2B�7�Ir��߅T$-�I�4��p�J�e�'�PҤ��8��"�����a� �\ս��m͹v�q���j]��M�8`���]`̶p�f�YݚZ���L���������< �9�����g R�A�!�)[�)5 I��bM��،��w]�z�Y�֊�����'��b<�([ġʼ��j �P�d��Bی����Ć�:�Ͱ�߰D�O����x�h��-a
�EP��.�kx35��#{ݭx3�f㰪J� ܙ��U�y���,1	`�p���|��0a��&=��T=r��e�)�)�����}����⦏Kq�{�����ϬM#�ޫ%I�Z���r�pǻ�ܼϸM����M_���Sx��@w�d���T�{�3����܉�J����'Og�]�KXk���q��t�J��,8ˎ  �f��j����$��Ƽ3��_�4�!�8��m\���GNCΨ���9a��%2Vv���Kw}K�ʮ�i���zL�a�N4�ܵ��n[����j�./�2�f�x��7h=V��3I�b�$a@�t�\��YD/����'��q�+�-e5f{���N�c�7�4�l�6��l�B���.s���{�������y�U�k�1#�:ۧ����V EZ�o]x���@���NhF��:���C���Qƺ"��2��1ԅoG�WN��s�p������c�����W>=ջ��GY��u'@�`�B��ۥw`�X/3H��-R3�}|j]@���>��2�wU<�H�/ֆ��g@�����By~�pK\�\���LQ�XN��B���G�A㯫�>{Ş�o�{�?R�T?+�����.���r'8��wr;|6���?�O�4�.W���F�\N�ty#�*Y�̚�6z+xnO����l0�x4�'.���y*f#Ӈ�N���_����7�(��X]����g���XO��R�w�\f�dDV���Ug��w&��zeE�>��j���p���Ǟ���[\]�/�����zwfq�Y՞�����ó�UnN�2�U��)��r���Ee�����2�n2�ݦ*,>L�H0�ƶ!�ʥFǴm��4�-o>ц
��U�e����tl��\^��jܙ��rv�8�)��l.��YRq}�Κ7yi��\�7caٯ.Q���!�9Z�z�[�����y��o7���˴����ڼ��J_S��>��GW��0�b#L?S�+bwNQ���n,��⩌ԕ�L����68U����#F	�5NT�̭��0�Qe����<L�?W J�tٞ����������m�gw�g8�E�l�7�}�H�C��{$���3]�!-ܥ�R���i�_8��g4�`}/�L;��7�N��M�O��{�O�Sql�PV��]�rP������ĂB��d���%��r�X����:lk�i��=��g�+��$���v^[�(��32b"��[uѶs��%0��;��'�I�Wޗ�ppn�5tHu-ٸ�x�N߲b�Q=k�A>�\6�7��|=��&l����P���`!���,H����|�}8��5F3��a&�fy����g���~�K�R쿑�}�p�ómHb�请������f��s�2�����ҝ����p�_�f��[I��}+=m�F��c�O=Y�4��^j�]�.c1:`Ea�JQ�λڞI��w3�˕'�H�0#����\}fn]�É���	�N���Q,�fj��z3��U�Rn�9i�xQ&k0�/Q��2=z�����ܙ�3Tո=6Gv���vb��sP�O�Ŋ^������@g��Mu�Z�ݹ�OrF=����ݏy��#�U^���귏`g���ϧ�~~ߕ�Ȯ5�˗V$v��h�326���%�h�IK���ӯ��~��@/��K�LS���vD��gq�N��OD���֞^��u�zR�-v�ς�$2���ʼ�@�N\����[~�T�x��n�t�恰��;0�<E�đ-��ٜ��e�������"'�{׊:�c��me�Om�|�o�)�0���z���53W�5X[��C��+|�b���(��`����Y8���ѫ����eT6�X��'�%9��:���m���Z�+��\5�6e���kss'.�U��'�v��4e���{X��^���t�L����5���A���k�jP���v��a{��NSE��+�6���L�̟�����?�_��������<�yli�w_�[��8i�����m����|x��}�އzy@��[�Ġ�,�3!F�-�
0"���Ͻ���l���*�k������80ec |�0#��fB���e�YO5e��=%��Q������߇�/+���7��f��;E�-!�U*�Z�Ǚ�r�g�aЅ�<�b2$C34��K��Ʀ�z#$��c�㺆C�(�b�oS�CP2�(U%����5�H&*��&���\T�ж�����1�A���RG��Po�wY
V9��"A�[b���I9�b3Jmu�^!6�.�W�jK���L��M?���z��_O�bQ������5^�6�z�)���6W9�\(��8���H�u�o[�� |��N��ϼ~�Vߚy�zBFϯ����v���>1R_E���NZ[7I5x��+&��Ωf���'�3����,���n�"���*������<���F�X�V��%�%It����Բ�o�]n�b'�혙�ي�S�V���y}|�1�cK�W~��\����=�GFfHv�:�h��ZgwS*Ĭ�4;7�U�=)f���I�s{�U"�[���B�'��۩���1���EԵS�׸S��E�*kپ�hg<-�e9n�����cϵ	�����SO^�"#Μq+b�{\��׊�޴���\ސ��3�~�u���S��MM�"+l�u�"ъ
� �����rԫg�� }�q�5��(��\3!�Q�賕�f�û��P{����0�b�t�d�6vY�'�E�66��n�T���<�5�a`j���o��|��tN-Q���-�U���g��"�Cw6S0F�/f<�
�`��7���P�����V�譛9�ƪ�i�_)�7��/iﶅqڄP����+���E�ܖp�2�!�_a��l{��7ӥ�zCܫ���耹�Z�<r��s3�2�/�m��l����e��M��fm&i�0w�@�%۶d'爋S���ur��F���\�[Ǯ���+��/&�̭� Xg-�p�_��������݂fGKKj����sx�M��=Eus������;p�,롽RB��NovUM�[|r�K�j�x?�y��a�&l�Z���=�N��}U�nCü���μ�^�h�}q�sǊ�;���2�_���*$�a��&E��<�V`�[{����g��N^�i�;DK7�3ٓ��A��T��n=]�w~����\؋q9E��e�]�W#q��V���e4W��r��u/�J���3.�.:�5�yL���T�����9OŁ��z`�'^�LkB���Y���@f�{8���r+�|Mdϴ�o�*lRɘ��Zy�����?t
�L
)lvv��.mg��kl�k"Q~���:`B{�^Bj����������'���>�&&a���#t[��@PrG��c�Ds[�����9V�,��8�pz5VQ+No]���<�>����f2⌦���"FG6��zx�W$�[��5}��n��'4�1KY�&y���tG�c~��[mV����+-K=%��-�s���i6�CS���?�b���� QD�Aa}�0����uM�=�:]���Pv�o���G$uq�Lk�%T�.av��6������k0#1��9~�|�xos�3d�]�)������=�b8��o,��]��ml�[f�~oo.�勇O�Ӣ�7v0��q"៎��i�.o��}�괫(��Dn�^���{��ؐpl(��'Ϟ�I�� �^4i��`���Z�Z%v��y�O��g�(m�t�i��Q٣��l�;�4D��;#G!����Uʠ�}U(0i����ug�KR5H"e�>V��{��1�)i�w���-��c��P�뺮�U`O�Nn�ީ���Й�ҽ��hVk�hl�Iۧ���*�P����[<�MVtZ<�0:||����פ�
�n��`ݓ��õ�k����E=���!\*�~�<�x���v�:{��o%��˘�t��*���(�W$��TY�^���)��8z<Kmt��t�z�&��k'�o�	���ys/"��y�q�Eۮ��n���&�nv���lk��5-�O�(yV:��d:;3�튤��z���J�IW�s�v:�{#�oJ�b���8�MJu�����y]���U�~?1�cc��w�}���|'s��6�;�''uc�������P'C�N��Em^�	oW4��cS�!o��eC����zz�z������rR�����9;g��h.ϗ>{��/�ܙq���]�U�^����a��=��7}O���PK|ˣIɼm�}�m��c}�h-�*�=4��L8���$�e[N@�@a����8��3J�F�b�����k�����>�%I\ZPd.�G��.�y���f���`��f߻�zſ��3v����f�������Ju#"�n2Y����v���EG �,0�k�U��*��/}䢯���ݹ}��g�ڂ��ժ�"jf��G�γI8�߅��7�3�X�2H�/6c;D�rszp���^���~����r(��_� �
���H /��TA?�QO�Ƞ��G���(`��ϫcN.S8�9r�6�dL��� Ü�r�lG#�;`�L��e����X� ��221F18 �lk�6�\�BH�220T# �1��3�e����\�G;` �0�A 0 1T��C`)�`L�� 9L�6ddb��$@$b	���r�&\�d�d� 1D�D��HȄT#"�d˗;l e�dr.E�E## �R!#H��0����E#"D�� H��D!#HA#� 1��!�#"D��BHD# �0P�H�X"1 ��P !H@ 1D��K�i��BP�C��!� �@H 1��B 0��D 0P��B H 0�� 1@��p��B 1D��B HA 1P��BD��BA 1D��B H 1P�� �P0��H 1��BA 1����BA 1�� H 1��B��B HD 1P��B 1������@3�d0!�0� 0����HD 0�� H 1D��B��D 1��HD 0��B�UD�0)�D `UD�0R �AHE @T�0 R �`��
- �� mD �@ A �1T �P@  @@�l ��0`�@�cbH0�0D�� E  �!HH� �B��  2!1D�0P�1�1�1P�0P��
��!1T� �D �!��R �B �D�1�� �n�� ɔ2�6�e0 �`�FT`D`��2v�C(d��0j*B�,*�`�@b�D"FFA�!�FF ��"���@��w?_���� � H��
F'��+���o������������G��?����(�����J�������w�'��QD@U�A������ _�� "���?���@��I��?����z�������C����鴃_�O������_�����I��A�Q`!D����"��"! �V � �B�@��@X�EB""�H�@"	 "A 	 �@ �@�$P !  ���A�$H�@����(DH�B ��$A��EH�F
�b!"��B�B(��� !�$�$"��$�$ 	 �(�$R
�$"! ��9�C ����`��� j*�H��F()�B �
$��"!�HB
�$b	�@@Ó ���6q�@� H1@�c��1@���"��� @*A+� H��� H�E	�DB �B*�@�@B ��2���?��?��Ο� �
H�$����$�@�����~� s��P�t�y�DZ�A��F������H~�3���G���:?�?D]��O��̞@W�QW����O������(���oЈ
��@)?������z��PP�Γ�p��`��������P�����
��?q���@{�<;=�����~��t?P��?'����x5��t���C�?�(��� ΃?q���K��(��J��?�����s�8��<���
�'a$ܔ��a�7�,?�����o�h���� Z������?� �?r�b��L���F3�	�� � ���fO� Ĉ�|��6�b�� [X5��0l0��Z�6�65&�����-*kZ�m�%�m��a�j؉5�Zl�36Tf-3i�eJm��fTѨE���+Zh*l���ekZ1�ͱ���[l֚ȨR�4�m��ke�Fc6��SY��FLm��D�6h�����V��Z׻��kkk�T�5fȃm��A+m�f�i��Z6R��mX���Sifdڭ�!chUU-�eZ�5[c-�����1
�l�Sj��L�5�Ŧ��Qv0i��Vx   ��w�-N����]�۬��3��텗rܶU�gf�����:꺭�X���sv����C.���Q��wj7[*u�m���ǻ��T�ur������j���5mVJ��f��#٫YZ��  ����"G�:;��x�xz>�
>}�k��[��Ms�a]L^��{�w!��շnۜk��u[n�v��Sewu-�wj�����m*�ݹ�Z�����۫���V�w-��eTj�m���m���MT�eV�o�  �<Z{q]vh�u�Fmh�;����k��4((����J]�uѲ]��[j��m���E �s������i+[Y��MRiRQU����   �xPP�i{�{��u[b�3]t֎vλr��4��nv��wj�ٵ�Qc���UGS�:�k���-�m�8�5Z����ڲ�ұ���K&Vf���  �z���U����v���3B�w\�*��ٻ���Ut�]�Q@�k�-�5�v�����N۪���e�fJ�MĐт�T�m2M
��  �	��BV�=�Y@����my�@=�w{dڶ�m��z�(��ד�-���神��KM$y׸�魵wnֻѹK�*���Q�"�=�M�Lɬڴj���"ٵ�|  w|�W������Nz	N��O=��ש$���{�@4.��z)QG��˞JQR�W�ҝV�s	�/=�(R�w�n��l������QT)���iVI���ՙX��m�Y�  �|U
}hV�j�퍳ݩK��]維�E�x�RR�Mv{Wr��S���y{�շZv5��/{���N�9׬V�6i�^��[e���m��E쭳U��5kV��NK�i�M�f��   6w�{j�
���sҵ��F�yOz=m��zn�����l��u�6ҥ{��މR��3��ԥt*�^�פ��ݩ����Om���^�y��֠=�ɭ�U6��m�EUSkZ)�V�  ���!T�	㸻(��Uޑܧf�^�Xyn��J������zW�ӇUUQ�{�;�AAt׼=v���U����<��aE��x�s���� �{A�R�� 4�S�4�)*P)��	J� @T��%*�� hh"��Dƪ�@  �)IUH@5?/���o���ɟΑ�������qa?�\�d\�3���bPS
@z(��>�>������~���cm�m�0`��퍶1��xm�1��M��1�@6�c����>|B����@b[Q���x����L�]X�[Z��N�ւ�S)tKX��1SgLb��Z�.��U�=��0Y���n��D� � �m+�u��o%e[�n<J�[�JM8��4�E@^5Ha\u�;�w)|��j)�����	.h�1���T�	�sv! D�$S�L�í݀��:��n�V��r�)�Qڲ���Ʀ3v�����Ȇ��`"&L�Xj��^�v�nH�!�8e&c-�*Ԗ7.�$�,� ����ۛ��ݐl���eMN漇k~��D!�`�
�0=��Pdv%��nM.�T��R��+��0^*e���q�-Ы��2��Ւ
�[�E#���'LѸn�]P�&Rړ�aze�ʎl;n7gM�&:��U�^�d-S2��;��:��m�\%Q��،����#-�0^k#X�ѩkF���Ol�aB�.��O,^�9B��HF)[��2�u�Ό�n&%�^b-�hӅZ��ir�s�;�2�b���^��c.���Q��f�I����@T|�u3���K6^�ʗB�J7�A�m�$ID��	kC��/�]�G.D�|���mտ��l�f�$�Ƿ��*#x�a�f�*ŉ��r`@��B�Ӛ����Q�ɥ��ʕ�SPQad��l�ړ	�cR�A+*�d�y.����(5X���eB�d�t����"�S
����7X�hI��u�{WN�z� 
��km�Om��p��U���beF�K�;&H�ZL9q�����t.FN��SK�v�(���.����n�]
y�Hfc��v�ԙ�uPe���u�\�xj�]hqJڋ@�oM'm��)��S,%�%�v��5b�A��в�8씢�A����J�"spL�q:)e�pls��*#>����i��C��R���߻C�6�L����A��Y1���5c��hPE��%A�:�6����v�Vە�mdu����nl�(�*�@@�:PPP�i���۬0,��ܔq'��;V�3N��k6V"Ėt�Xz�,�)&���iT@��J��y�;�Z�sܧ�d�?;��dhU�$74!�)(�+��j(��)�vs2 6,J]�vmdEm�Yq��k�J��U�&��שU��Cj޹�f`�Ssٿl߳PJ���چSZ��,Ӧ��͘M8��R�W�����K3p�/r��:��$���0���nĭz����t�!	l�� ��YB�칧kQ���Tc͓x\S��ȹ�n�y3-%v�<��f<�p[ı���M����ڔ��XLS�c����M��z�+!�D�"��a�ړ]޵k[��̉B�X�1�h�b�'��nd����ڀSb�sf�dm�̤�,x+"�����"�Tۂ���!Ӷ�4Vݱee�e�r��y�6�lݭ�y��<���l�Y�'1��Pa�F�ɺ��Mn#u0X���*�d�:��[����p�i�4[o�p���wL��.��cf��K�yͭ�p� -�������da��`�/��9���B�F�\���0�C��A�m13X�(��U2���S��q�9i*� �c�nU����
d _�-�&;����Xf�"�K"��/lX��Oe�ҧ����B�1�cJ,�yv���ne=����t�-)h�b��Ŷ�DTt͊�,N�5n��5�u�̽��i&p8��T���~�j��u�P�ǳ�m��^�2��d�a�
���5�ceph��)+Vh�e֤�]�N,-ګ���R;;-���M�y6��yM�0B%��'��"�X \r1%a�:
h����غ�M5Z��W.��C)�%eMѶ��15JJj	��=Q�3(FMd-,���xq�uQ�E�J˂V�W* ԩ[hj�9��5.�^�%6E��74�0����>����Udn�\�F�ͫ��N��\"�k+1��B[nV��7CH��tS��+�^�a͋G�7�)LL�u��ei��`��^�k�%	r�/�$���d[�Y2�y�U��-Ԥ	ŵy@ۭ�x\h�˫m^�Ō���ef��v)5�-�pS������h��57n^n���&��ź���e�����;�yZذ�AF�ͦf���[y�%I%aM1e1n�*m��6h�J�T��ZdjU����4�sR�5ޚݦ���J�D�GYL���'z���#[(X0��VT����/�S2�Q��
tR5��.����"-WnT�4ζ�h��`�0K���5 6���vC��;H��]=ȒY���Cpa�h��2��n�M�Z�kZ�QR�(Z�Ҁ�w.��+"�.�i���!0���IY#a�u�ɠ*J�8S9�
`�v�30�V���t�E���[{qk�h�+���{�۶����#ݫP���V�ӭ�C6��I �;nMn2c+:#X�*�}���KHё�X��r��2a^��XۇK�r��s!NT���:�����!�OB�2�6��� *Î�ˉؕ��i��+&���4k��U&Ps���ZM\j��q�r�m��&Aۙx1aN��jDfMK�7!.9%7 ҵ���#���`��#c�4�4� Z[�"�j�D�˦���W�Ц�e�&
B=�
A��WIR�7;[������Ƣ[D+tl��`x��dͬѤ#��^LVКu�;([�K�Y�5XEZ�[��KM0Ѝ\nnQ)�fRM��;��
u���s&��Z�[	�U����u�i5��V\�t��r�)k�`����5�@�n���e�^���2ۃ[��Ӂ��(^�X�"�Pj�+.������I�r���`P@G��Y�'�$�cj� g��"j�ۃU))n*y��hV�n��J���uD�^<��Œ�yB�XU9nFTwzE]�;�Y&���[����^���M��&���sSf��T���m��)�q���d5��"��H��K�@��+HFg�@V��m��U����<1a�8���_'������p�r��
�G����!��S+E�P��S�`&kf ��*�u�Ʋ=��������h��J���j���uR֑��qi���y'�u�J���U�[�4�
Kƕ����������l�\��b�Qe��i[�W�)X�Jvk^�e^SmEj^@*oss(�To���mbm��U�Py!��Bڍ̘��P�Ԯ��ˤܑd@�A�v�b��,���%P��q^�qM���%+P2ճ�@ӽ�s�P���L�x�Ҁ�;��#����a[�k��7S+.���n�f������"�����sh�9M r�B��H���$ɮRЩ�z�iL�R�0�Y�9h2N�i -¦ˬ��S2�.��/+I�bVѩV�S�S&�c&Ee	Y��Orى�֠b�5�r��-�r�WT5�%�B�ߑ1���Hx�a�>{��'���9b�)HhI֋�n���8t.vN�z��+NAZ�2R;�cʗ�����L`�i����h�� � b��j�rd �0ۭ��l"[��Y�6r�nĒ�vm��3ql�ĥ9 ӳT��U���j��K'D6P*iu�M��4`ݺZk	��`)�@n:�Vm�r2btT̃/MlN�u�tv��ɢ�<��Wd�f�f϶৻PZ��c�sL��.�bQ��H�PnJ����ML3�T��W�h��J��]KH�f�GH�yY.��&�"�I�zJS�J�!Y��#�����mf�:޳B�(:�?ٛ	ܶ 5n��ۘEǉ⧄��Vd�Xk%IBi1�2I�.�5fU��h�1�Ց��Բ���P�����q��&�Q��G�Y۷2��<nC��eb�rR�q�QZ +�0^]��n�����EA�Ԉ�F*x����c��D"�֙@PU��9� �lT��pM����GB�T�w:L:��,6^�7&ET���JӤ葈h7�t)�0�v�C]�ʘ��[v$YZ
�c�Ɛ����,�s��v��N��(:t1�g-��$�a�-�Z�9&�:Gٛ���Sf��b,�̠ �N$	P8[s���4��̀��9�",��dv��W��yJ�z3	����9�CyK#ʗ�
x�[��Ш��^�{v�؀��*ѡ�K�z>h͙�fe�10��\�ڗ��"n��Ct�Ȥƌ��b�b�`ك.�F/Qsool�N�P̔6�K�pMnr
���«���B��6ٌe�����2�I��0Z;��!O��9)�}eG����uv�
R�˸�X��fIel��W2�, ��pU��N�IyB�
[�t�"�pV��U�Ù�#+v�W4}(!BG&XvŔ�H�)�����L�jYwV&ۼ�]�Pt����#H�@jՕ6�rh��e�X���FP�-<Ե^U�Ea�Դ���*}&; f��n��R�L=�f���U��*�(7�nE(X�KV6�ݫ�K!�m��ݼ�M"�f��#0n�m(,P:B�k�	Zf�r�`Kf��6�Cs.E�QN���5�D�cڀ�
�૔!n8�ԭ�)�e�o@y@,�YQ��9,��뵖򐕪�X�[�f��IТS�n&�T*�87+�JJn���sT��а�M��Zmjb������-���{P�ȱHƈ�(��,ojG�׏�}V�6vg$��j�LeDk��R��b�L�]͡$����(���q�m�-��A`�"���7Y�ZI��J�u$������]��ݛ����RyuљK&;�u6��"[�jn����b��P䶀�K0���/M?�u��-�1y
�l�On j��H\��*�z���2Y[F�2�ʹG��5Xuu	��q�n��ay�\@���.�:I�G$�m��)j8���@�1˥O�2�R�R��0:� Q��ׅ4]i"]L�P�k���j�`-;�f���I�,L���萪k3Y� ��Y��;j�ZL����s%�t��Xⶋ��ia�C��� �V�h^����-����ݽ�7f��hp74�$j]�a�^�B䙑A	��Ye8vTWGljܦˢ�43q*�!ɻW����#�-�5�j���o�!T�M��t�sJI/(4�n�j��V����@��"�Uv�x.$��9��ˠР�,���W��Mbe;v4a��YV&�N�Yu�m������)���J��4��kn�i8Zݍ����H���(8�U3]�x��5�&�4o-L�E���h�d��T�ڤ�3w0�����̺�U�f�p�@(�;��N�`ѥ�%��b��:qiu4ZI����Ҕ�T�Ѧ�-�Yh]�X.�DYs,��n�E������U:<���Zz��z��n��8H&aj��lX�ƍO x�W&E�^�ve����F1���)�hv��p	����ۅEp͟C)�kP���a,R�����Y��Sj�`2�x����G�L��[yR���xJ�N��sG�/�h_��p��*�y�f ��Db��{�FƢ����B)Y+d���-c&9�@�m�4] &���J\�&���ht��oRƌz�蘬	J�2wj�[W���D���7��np�e�Y��cڵO2��G���0�5��6ֳ6U30�X�l���Qm	�0m��hf�R�@cʷS.#%֕jl!8�E��X���1�����ɢ��)����h`��b�w���*��c�Uީ�f;�e\�m�M�񛽉'����v3L�i��R�����10w�JŢSX��Q9��M�$[˭���{��[V.�;�7u�m�2lHnSQ�ED(Ǵ��sZ��m��w4[���mY"[�ՠͽ�>���cB���*�	��4ЭT����GQe�`��c"�`�RCdn�Մ%��@=�Ǭ͘ԚڙJH	{���ô@^�jf�"@��Ø�h�oj;Wg���اW.�d6�V���Me�Ch�i�P�0ncY�8顎���z6I�͕	*H�t@Dدr�a9��9m���^n|�m�R	��\����y��0�s2�L��p�=��(�᧍ܸ�?
���-�[���
zؑ���t!l�Kͩ�Yzu;vбZ⻫yZ�`[v �M�)QA��j�0��H�-����:`��ސv�.Sś4I�"�Vi��v'�������y�k�ܷ,�%Z �"�o%�VLR�LJ��!U5%`iSp:+#*V]n�g+-hdi6f۴�S�a�����!M��3�VV��%�[�/G#���`ܛ�#�7��Q�m����+�j����q��NT�j�2�Y�XFk�~q\Ϧ2�T���hV�܊]&)Q�P�%�-iT��u�Ė��l44k�y&�0�v*Sp,b�'�c*
��fг���H���YvM;����R�@������K���a�&c9�Z���n��X��ۋI������IX����j�a�[vAn�6�b�h�h��3TM�D����B���A{E�$N���V
5�&�9��ɖ��OBF��Av��++^����+A�Ah-+"��IG�i��\�ֆi�tP�!������^��
YI�VrX�n�2*D��ID-MQ���md�I��PW@ ���cf�"���t��c����ǭ�}�d�Y�7��Q�D�ӵ��àc���V�`��N�S��d8Ѻ�E�F���4Z����2�����ߎ�l��-�(Ej%n�aIV��,VRa�M���R�(զnѰҴQV�U���Кn����Y��:ƽ`����WO)c��8�g/m
�5B*��j�j�N�ŷwh��һ�i�Β��3*�E$y�jn�`s��n>;Gp��դ�4۝Y(�ْ��};u��}�aI�	�eeN��e삣�ճ��F؏���-ߔ�KY�k�,Q��2+�K����(r�6�����k55��������������gT;i��;LL��Y�G��
:�s�yn#3��";�{E�(Y�'wC\��/�'��v=(�+�{xZ�+5�i��3y��f��d�q��y��ޭ=�s�uSu#3@�<��6�������oFP!�9N�<�����e;��e �*[*h��Z��Mc<U�k;&T��Vm��
�vR��(�o7r���\��@��#��_	�6Y����^�7n���@l��,�}Y�,��ۥ(8eq�u�����i{%o�8(�.�p���ri�m���-���@:�7�K��֋e�R��chq��yL:��:<.���Ч2�[ڀ�}Ď�I{S�,�-6q�7�9����Є�#V�<4(���bOcՙ;C��U۔�e�U�5P��l��� ީ�QR��¢(��l���}�r@��4D�|sWvf�m-�����O&I ��|C��S�.���7�Q��cݛ묛�|���_A�9���jJtt�,�����޴���I�6	EZ�����d�*�v7�`�39r�\�G@�+:=x�5�r��q�dq�(��4_J`�೶�@�k�wb��M�R��U����r2�e��X�WY���E͕Ғ�*�!1ßl�IP(�=�X��:7|+b��`-	��,a�;Q>���V
�v0RX�9n��Mvk�v���T�ӄ۳��;��Wh��zT�c�t����b�ě�o_j���,?��_BNN7)i7����efP�o��32�6�J�o27W%L���]�R]��yڈ��x�V��=��Rg�R�y'p#��R��ݻs�A�:��W+�G9	u��$��4�GJ�*���vD��h2-�ʻ/T57R!�Wg-v�����lv�a�� ���@��;2D�DO���h]q�;��;���z��#�����"�62ɗjW-#�*���v*T/*{��6�_ilV��¹Ra薡�ұ`j��|0qU�ҏT	䌊�+�I���)[Sb?9S�iuy)�jK�+��J����j�l�5ևw�}I^F�G9 ����=6e��+�Q�8(���x�(�F�O{d����hZ�e�Z+���ܻ���Ԙ@+�T��-���־���ӜH���:�G�,�;�hO"�B��h��H��T�w�2�Aw(�<�(�[��Go:�͡$�qU`/��"�u���T�;��z.d������M�{KD�׎Pk���x6����v8l�4�9z�G� c�0���ݤP��������Beg.���l�9��#����P��[�����:���ڏ���o��l�ȹ|�xDdc��4hn�Eֻ�f�����|�U��gV'i���bL�C��v��1QY�$y���mu�U�gu,�8��u�]:.�rmAv��X�.r�},,��+�#�������69�u1�
�xz�BQ�Հξ�|�_W����"�j���U��]�E�WI%iR��.�V��w�9��ilԾ�K�f���λp��̹��&b���H0�k�E��qT�u��c�5��1����(1���3��/y�0I�s-���-�R���;�Jj�E�7S�e)ъŽ���gK���mtT�QI���������EG�"C�u����9��1;(Q����@�B\ȸ����|uN�9d�/�i}�w��g%iڕ����7P�[V	KU�i���x�AhJc�I�)�9��-��dls�����cO5O���W�u���4;��6b���3-�����x��w�e�v�m�ƥ-%J�M�]}I�Uن���l�y���]�3Z�ŝ�� n�r΀c�V�L�EL������2��U}3u�}+=Խ&oݑN����p7��8�����܇�z����� �z`Q*x�6es�6�F���f���"V*mWm."�k7
r�����Rtpd�R���������`�.��2ݩ���Bp��D��T���w3�o	]v\,L�}��F�H��w;�nk�#�ʹg>���-�N�Ҥ�dYD�i�x��0�1C}�2����j��.�.w7������;�E-��QmU����V��^-4��]��v�����.���rr���3P�Q�."�RYP����*���=�'i���K�.�z��4�8���ڗ@��^Ws��y���X��U㇗\��zty���!.���־�
M�SjCǬ��iNO4t��v3�e99��X
���(�G��R��k3��o�+������4V�%���y,�z�*}�~�c��;���7���U�T]t��ZWPC&���*�3�M�b�0d\$��;/c�ʙ�^�QK��Z�BÛ�9�)\�d�H��sB�q��!��F��.�j_S��6u"ɦ�q=7�.3��� �cVR�]�RV)B�]��q�/R��{�S�Պ����&�� ���E���4h�mN�����	�H3y��X;s �S�Poմ�szR�v�dr�7� �nݾ���8٫��g n�8�	�FtL�7�4���Kv]�>���˥N��+���c��c�[�e����y��X�����5��lh���<�թg�\o������t�BMJ�]��R��@G\F�Ku���q\��҉4r�=|�>���y�֥�q�yT4)Nh�F���B�Y����;��g]K�N�K�n��
���w����t�6��I���9j�f>�g�t喨��0n�@�����3T��w#��lZ�h�/H���fm�Vs�:b:�N��ȥ\K:u�(u����:�S������d緔�F�!'P֫��ݛ�+�MK.�NmXֲ�XO�4��%S|���A�e�p���)�K|,B�G����ك,r=�)�ue�v_?�JL|s�'��]�YͽoX�\ l�#��󆁜U��z�\�>���8N��c/���9�"O����EW��a�J�m��޷c�א���\+�˝/�q�@ӭ��z?n۔G)�S轲ܺ�L��WWm�]8������% �ov	۱����v�wq���'EJ��WǍ>�\�����Е��x5_Y��;{V�=TM�Aހ���QG:�iS�7�r߽�o�T����eݷ�(��� ���Me��M�Gz✩�c:A]����ާ�ս$�ﰜ�JT�%�)�������7��h�IPීn\zV���e������l��w���������3&��x�;���g�ڡ�js�JP�HWQy�A�>�)�h*��׫�W����< �2���jq�3�Ǫ+}��P�Bo73,r��ҕ��}��%�}`�s��G�n1;C̀n���s.�;ڻ���wps��ܬDǦ�f� +3�d�+�3(;���������+�Cnphl�v������� �{[+����Isn�VKZ)]rrM�#0��MF���@t��S����-�0P�z����m�P�6�)��Y+�r7��B��t��yj��\'��ƎK9��\��[7�'�PJ�k0�a��i!��C���z2����5{����O����;+ψM�!*fݮ5I���9�J9�O!Ivܾ�Sq86�B���Ʉ��lh����qh��Vgv�'s��mS�)E[M��!����Ⱥ�0�4�k-�5��J�*��]xy�嬭�?�������V�UΩ��]V#`T�N�XJP�2�Ő��8c��!�� V�V�R]��;a��JE�u��
6���,}��ӝ"�]�I��vY}>��Q��N^�;�nZ����(X�������O��_m��ނ�(0�N~���S�Ʊ9���IY���6;�	9ytҫ���Y�r���1�(V��-8(�Fc�g�z=R*喭�'
�V}d�fQs�j[����ն�;E��M�܍+:�N+�Cq��{f)D9�TNi��ʔ��sE���݉e�����IkhX��E�Z�i�ٕ��Rt�³�X�cyg37���O��K�r��ᦻ�P>/��u3�f�CqH"��]�Ȼ����X�=����`p!#�]�� m�9R^ě1���w7W�j�.��iV��P=;��Il]�]Y��OF;�X�Ҡ��P�	���ų����/oV�mnK����G<x�=��o �#�7�r�"�Xv)v�5��a;Wu��o4����h��j{js=㧵�ٲ�DDȟm>7k�p� k�r���#��I/ep�\�V�f���\6�ǞS���[
����^+��c2o*V�d��k*5�e�M"� R����9�D�L��L7Sf�նث���m�RY��3r�Y��I�G�el���e(��v�+�\�� �}�.]9��ĄI�Ĳ#kP6�V#�N<��ٗ��.;�� S�里S�0m:�1q�R�B[ڔ�"�Gr�a��^�R���9�4��V�c���8�M����Y�Ŗ�����%�R����nr[�l�ܬm��Ot#q46�ɋDs��]�۲��1\p���{M�6$��֜��.�%M9I9{��g=]��O�[r	4�k+���Jh{t���j���y]�����OD`�y����'%�q�l��E�y��G��],����a<J3VD�)��-���#s��VQ�<<E�e��5��9M��vM��6�� ����W���9*_
P�9�ۯ<�~���<�ӑ��� [��mqGf15^�h8A[V��F�
J`��anuE��f:8�ʷ�v7��*
���\jҙ���}�ѽ��`�9�W2�.Nc\�(�Z����'��ZOge�5N��ӹ��rD��:n�(�{K�L%J�.�2�r!wճ�79nV�\�k�oe��/�]nkCV]q����ڶ�����ӁUo-�d����Φ
�)�u�ݧ�o�����.d���QI�Ì��,����FW<���l��dN�Z�Բ6�_��@Mm�=P[�B+��tT�r#�R����ۼpg�R�=z.w��������Q6̅v!"T+6�V<�Yi�X{�����mJ@��Rqe�]YG[nu|�q;pk��)K��F0����9z�Z6b�`��ĕ�>}�iIg{Q�\�J�G1�޵�ܬ��wP�&�3,�Va�b�I�&3������۲�_p�,��:�|�K�[j%��6��y-.q_%��[�����IO^wv��nԫ�q�N���dg)vL�#��D ��%3��ox�Q�S�.�� %���}F��o#%���������m�a�,dB����A�;f�6sXw��̤��`Z�-3B�sQ*�l���Lw��	�V����;�Z0�,Ҹ-�5i�]�U�h˫!n����z�]Y-�-����N�������M�g�l���*uЅ��jm59h�O�n�c5iැea�]j�l��fb�})���N�⫣�駹�����-Q������|�g���LvF���YL�T*wu_oKH���)�Q����G/�׻N��=��X95'I�p4�K�.Y��p����Z^8�i�t'�P�w	X)�u:�l�뫆E��d��l�"�86��BQw��w6��S{��wV��;V�7-�鮧Qu߱&j�
Ӡ;w�u.j>�Ԑ��̛N��"�v�VS����y
,Mm�V[U�8pq����<�w�x���s�lW����X�V;��s��ķEӼeo �|���Of���nn�a�
X�Bc�ˌ�ұ�/v���C��y!/���FU��fǓ��B��)��X��\�9]kt���]s�ŦX��l�j!9��)�\M-��ۘ%�프��d����ݒ��:�����k��N�wV��%�m�
$�K����B1dg8�nv��+��򜾜�H�!kn��3�Okޙ���R���	5���n�Q���0]:p�]@�;�����r�{[5��aNŎڢ顉�3�f���&"���Q���zi�F�u��Q�b3�����/K�����QN����g>3N��ܝ��
�w�Ҁ�M�s/)��ۇ27�]��U��`v<llk� Ƙ��#���ٓn�v�"�)���`�Y� �D��&��R�{-��><V��	�mM�b���J��7��Ig{��ޗ�j�����j$�!ϦVѲ�١:���5���̴�r�uZ���#s����w-�W�w��j2��L����wF�KY�iZ��q���n��T�,���T�>��ѹf�����m$�*�vĹ�:5S1tԅ�"[G&�L��u��t��JweL�����d�x�xd��b�M]+���X�͎�60�Ͷ�,F^MؠO:f徽��j�����^�]�d*>�
��ۍNA���D.<���:�� ��c��uqUk��T�ւV��4G��>\s�J�YJ�JZ.n+l׹ c���+m�#˭��]��Bv��_�֥G�`�`�l N���V�c��K�뤰����4*l�E �j��&U�ǵ|���]����%�z��f�80�L�A5μ�6^eT���ll);��eP���V�u�:O�u����{p�x�ao'r-��]Lsq>���aJ,{�͕�']z�΋�yR��m�=����W�d\�o��@N��w�AB�B��Cu��n7��.���3��l���E]�^���u��˖�=�Z9�}����
�'�Iñ�ݹ]8�=��˶�wPZڵ��L��ECp�3aw�*� {�u'�9�Z��7��bPooN��S��ݵ�'t|�S�"�
�,qG��a���g�&�����ILd9O��o�ST���C(f�LudG�c��}So�m���߿������l�?۱��6�޿�������œ�qS]��>E⫛�noz�@�RV�ЪC�۫k��1㝱����0[������-�N��n�G
� �� ��r,Yd�:�����c�6�n��r�/�3DU��J;2�j-фA�6��P�@'��|�! "�7�"�1��ĿMAkt����g[4��.b�j�}X���\��J$�ɖ�c �.>u���y,͡�w_W;�g$̭�ޔ�Ex�tYikn�F�eQ#^��L���H�Wr�ope����5/8�g��zt�6�@��js����fHʓVѷ,��΍
�/�t�R�K[wz�Q�+�5pc��fM\j�^&lm�N�wb^i�I�Z��+�ku'���\$5Y�e>�1ٛ�P"Ns�sV����y�p介@�4�E<D���\Tԁ�Z� v�=��E1��و\��V@,2V��]'soF��:EW�+i�R�t멪u�+
�f������u꬜�
n�!��oNX��e�|!�]���̕�0c�q�8��|����{N��L�����=iwТNU����-5���I�n(�#
��5����O�v�9(�=���Wo"� :����1k��;���ܼ�]]�����;�˱������ t�%s(!����V��CXy�{Gv�u�F��P�E<�n:�䗵��̿�|7%``mm�����N�zL��f\�Wf-�����)��;��N��B��r��W;pM�)���!�8�o;`f:��eYۮ��r��AR� �v���.�dC�3c�2�]�+��`�g�V�#�����[��smd�F��y^8�v� �E�L{Ab��H2���w0��?q�c�k��S��h��8r��F[�sN�n�{йzC�qdxU��[�M�!	��68�]�x;��;�V�I>�g�f� �Wn����
��R	��g@��XL�f]H�u�꛵r4��{
�߸�]��C:V�滨fC6�V�e��3"r�aY��TSʶއ�ַn�p�8�����х�ʨ1����ݬ/��b�7ˑ�Xݠ,�䓋>TY��L�b���B���`P{�[�""1v����]�9�7)./�d��\��C�ۜ���D(��f���H�dugOot3eѷ"���Wu��S7����X��OW,�Xő5�(�wY+{��Ĳl��N�c{Aa�YS3�&��R8GR�y,���o� ���t�E�д�Y�X6")\�D���D���DGP�Nu�W|��X���9����C.���UYFFL�H`��Lۦp^����c�x:7cH-�.�e���CgA�J(���q�6ŧWt�`����-t��=� f[�sG"˔s��k��b�*i�Db<���]^Kx+i��Ϟ��T�������t7�ӷ�#D͠�}�7���9V���%u�Δ�޺�WnΜ���r�=7l��é�]���:��y=�ӫ���v&�uӚ�7ݫ8)/�7��u���a�,0zfM[v�����J���	r��� ���t_J�oc�K)h��{�P\+�Y8�q�,I��8s5|W�l��3B�(�u�Mڋ.�A�2�_�v��n��;�@m1»���wpɤ�h^�O;D8ۣ��쁠�Qz�ŒD�]X%��/��*������G+���G8����D$�r¨ʫ��Ė�>B�rp�'�v�Gq���,�=��8���R�՚�Y��!X�P��u���j�WJ/�]HDs��+��f��v�9T܎n5�.�g_uB�`yM�
9�)�/�#����a�/�=�f�®p�T��𛹼�������u�Ġǆ��r+�w�Ǜ��\5ҥ��1*O6q���z▅��� ֥VƂ��=smt�Cg2)k�&����^i�x�WV�F�tv�[2��p=7�[1풻��u:��Vҙ��LhV>f�8Q�1��0i��f�1���{�T{ts��o�w��N����ۖ�(Do�c��[�zӽ Wp�n��O^�FQn��Y�GлvI�OS�K;^_s��<�E���C����`�M��9)���p�[G;�[�f`rt��k\�)V۾�yD��묾�:�T�V��.���̒7���쏝����]�.��6c��\��]�
���E2���*D���F/����a)}���yoN�W�K��N��g�})�v��VY�F2�B�Υ�8��6DK�R�r��nn�wE_B���[%���70�@�Y�	�2�od�/*wY��2esѺ˚Ⱦ׫��5r0a�cy�T6����2w^rÊ��w����?fG�r�%8H���2�C�8gޗS�́��q��:���؈�;	����;�pvf�^��&)�q��/f'��N��7Z��acޣ&�O�m̮`��y���0�hI#�u.�A�^�j4&����:u��V\��!�ygFm7,u�\'�����0�Q�aoj��[I+p�fg`�����?
�U)�����xnW,i�z��>f��V��[F佴�'��9b��M,�r����7Uj��e�
@k��Nנ��k������W��
�sF+��u��-Ңj��1��qA��ko�rW89[��f�t��`�յ����9Ca�;!�*��w��x�Q��Ȧ��ɓz��u�[Aiy�
9mwt��R��|X{�6��0�ۘΗy�5\�9���L�{��ط�����X#����37�"���|Ĝ73�`ފ�)�V�lу�Ï2Ͳ�<�H&�9a([O#�SA��l�1�%��Jݚ;dCv�OLS���E6�]ӎ�q�v�\�I����Ƒ%��3:����z�o�it�,�/)X[6�SMn���m�Ҟ�M�Q*u]+��5�0�� ���"��]���}l�˒�"��d��p)�o>�5%\�sT�8�f�ǎ��I�l'j7��wr�M����Q$�d1�O8��4R�F�n�DM����j�wU��mq'Z6r\�[�����<��8oQ��u�M�Ң6��M��f'֝�;$��� ��xv�un:v^����;�e3���Xj0� �=7�xx�n�n��.����twu6a l�y�ݝ7]�k�LT�C��2U�s`ҭ,Kf�|��vl���m�``s�P@��8ݡ3�5����m1÷{G\*�,u0y���x�C�K�ɵ�w(��ֺr/^�M�(�i��ˠ,XKa�]�}	jx��%���ܮLwu`��+V�.�M�f�6���BE�V3d��F�܌��g-�F��*V�0/�a�S]�e��yQK+�,NX������k��d�D嗸�lu�B�YV�,O	�W&�Ì��]�ߙ\2�c�2&��������}�<��ʡ�5�K�q���ݭ���x;5��f��\-!9�nn껩>�U�L�ҳ��n�-�]�ԑ����7��G��nEzjf8��rT�}��:�}��u*_WA��Y�X������F�	L�Ú��c����:�����j&��D!�����;d��ܧs]��h�l��ԄU�@��7A�^-�D�J�4����-���K�VPZ"2�WN� o�^T��u�R0f��y�D`n�vܲ��ˣ�'H�k
"�u��HΧ�[Kn��ޘxc�)%�	]��T�l@X�[ՅB�C����]�mvK���K���f��g_p19��탘�<�ݓ7y<U:#Vr��OtE�H=u����[���5[YX�y��h�B����ؓ��,�e�'��g_0	j9u��`ݧuH2g'�HNDmݻ�Y��c�1��d��޻��0e[�At�۽���k�Z�oa:J,��FwD����D�q䫰&;�5U
�/���s5����)vkZ��]iJ�%��:|�pF�;{IS#(q|�=-�P�c�65��7�uAZ2w�8)v��q��wa;���r5at;�o����1G
Ŋ�D�oM��]m�n��,�lE�����nd"qm2��2�ec��{Hn�r����E.�1v�[�5�*�{�*^��p���W9�����ﳍ��k��fm�4y�&�K�rE����#�۸��*)�"̓)JsB�L��n�y�Sţ�\kX8���B��s��s�sU][7n�1����4��T��&R�D���/39�OqpoFNT�<*"������Ωۻư��'�G[�G���X
)��f��\���h���z����RIJ���[�zn�O�᝛��a����KclƋ,��*�����j����IS꿰�,��L6�]9j�k��!$K�,��th3�b��M�(�`�0�ι���M�����w�(�ꥆ �彮��굤q��}��Ĺ�L��o�q�@�Ǖѷ;��Z�]*�Y5ڰ����+T�cYN�ٔ�G-�m*�SLe��׏�[�����ǂ6�����:K����#PWVaޑ� �\���f6v68e-n���K�C�ae:[71k[�hK�i�Tp7J�7m�I��{�f�/���3�A@�V�ܬ�Z�$�bL�#�qn�����e2�����ث��������Ou	�]�,hr�[���ɬw״a�5�U�\�����J��{�ur&}sy���d�2eK/k*�7F#��@���EAg���j2p�bh��ۮ�S|�H@�!�y�.˅��8'N[V� �Dɯ�E�R���m8��d��I7����h�$좏�/7�w����"�:U��o�ɒf�����#@��Pԧajk��yڳՉ-N��F�h���^jlA��1���6�7.57i�*�T�1ܒ$T�z�k�E�+ls���S ����贿v�Q��Kv�$ЋY��ѹ�WcW�uGDj�.��܋����j�5k{����_)%���)��:�2��J��#�q�x7m�Jů�W�/�؃��U�଴�N�G҇[|��Ӳ�_ml����Kx�A�l �E2B�]�vi��w���vH,���Nՠ���@tc�낥�J������Ҕ�8�7NRJ[f��G9PJ�]u:قԾ��_
�W9ֆ�r6�K��� Vs�h�g���9CuJ�CL�)���}-�<4���8�4�k��	�Y}���T,�#��L�h[]u�����;�)n�Ѳ�sjn9㾬��G;j�iR��s8��Q
��ÜW���MS��7�T�K��'5۶0-�Ko5�I���HB�����кM*��T��ھ����/�vLm��f"�36A+�����TСT�LIn[�.1��tW	�T��>�P93����&�o��Q�J�̓^����ά��wÅf䈡����+Z�β��Qu<{*�=#:D��
�"G:�G��u�s1n����̐$�b�N������m������]�6F����nR��b4 �)ڮ��_5V�Tɼ����j���:��n��-j2s.����*{l�T�!��0v�W4��m(4+��$�M���Έ%�r(:��;��(֕m�F���)�S���v�kFg#Y��������N��O�%���9�uGS3�b��zFW	{P�8�=E����uԅַ��k(��۶Y�!�^:�6�u^b�oL(��i��K��J�,U��d��[@���1�eN\sv����v��,���S������d�ݳn�ӻ��;�,��T�r�*��K�{u�t-(X8���s�	/�n��lk��� 	�Q�x���Y�I����!}�mon���łQ	t07-NNL�ZHλipd�:<���V�'�ٜ�%Hz]9D�ܛuu�
!WgZ1�[ʺ�R�ԩ����7�f�Y�"#�]_6��E�{;�
����wU�5�:�z��yu7/8T��Eҙ�\	��RFv^=��~Yh�r���!&�CpU�*C�)�r�,n�77�N��zt�ۈ���]����y!���Y��jN��q��bk\Z���Y����6�)��5�������S4H���<λAR���f��1�C�+w�tJ���[R���vq́]yW9��?pB�Ι�C��ǖ���@�QPqȓm�i]�y7o}�%���<��Ԅ���&)A[����H�Rj5KM>��wP,�ĺ�W��W^�Ux{c�k�V㡉�[769Th�N7�vA��M�����m�	�l�U�O%����J>�7
#']�A#��l�9�Ee�wG�
:ɯ/�r.*��E؃��ʍ�MY&�uc�7Z�z���_9+���22̜��u�T:P��T�lf}0��-�e6r�4��hptv��E��d�*�b�j4��o9e�3#_��{�P�T�������e�t�t:[΀�0�m�����Ǣ@/y��'FmԬ���c�N��v�i���fݡr��V�d��B=@�C�e�v	��� ���T��@eX��'H�,��z-��[X'����-�pL��`�2^T:�=z�Zwr�2����8�%�6`YRR;}�`J���*��|�@�nu�6���
	����Q0�%t���e�ҕ�oi�����A�$Ł�q�*��Ҁ�L�Ƹm��s���)��g��a[����%��ݭu�r�Z�r��+*v`�K%�8����X�"�G��vEE�wl9V[��(��0n��!��}�-
���7Nf�,����$����:+u��J�����4�B���h���y���k�eq�AlV��Z6/�3أ���C²�F��+w*S�u:X ͪ�;#J�jjq��Ӫ_3v�����b�>�#�ֺ����]�v�G��,l�R����ʚt���6DI�T/jW���Æ��h �����^QD]O�5����g&��9T������B)`[N� ��q���U�w0��Hb����]6k�&������>���~��đ<7�t瘳��T��,�b]5ܮU���ER��YzEu.�;�R�6_P����Nl�>'䚎��B뻸�c��:*;Ƥ�ml)Q�ꆗ'�2���;f���#��Ńz�SR�K������Y��i�Q-h]�`�H��}˗R�v+@����7��N��o*�Lc v4&����Zur�y�F�i�.E�Lݼ�I�K�)�lV�IS�P^аwX+ek��dU|��׶����%���l���F.�hr�����b�ި#۳�cf�|�G���d����z6�Iz�m�| K`��֓�;��
(8e�fu��Ѩ*:���_�!�iY*�	h�K(ӫ����<�����wf�5=�IV���b7���s���'�o6�����﯇HgC��)C+��'�)l��i��T;�F[�����ͅ��)X*�]�l�U����#����PY������P�(鵖��^�z8��o:yd�d*��Z7����(]��Y)�Uݮ��ֻ��iW��@�?h�*ׯoIy�Q{|�etH<Y|̾fT�f�R�k��[��o��h�4:�����t��P�_I�e�CI�񦻺�=*H<��Jబ9]Sz-�eE��/O�l����[t�7n��J���	�:��p���e1׺Yӵw�:�F%e[���pljۊ�Z�+x�ݿ6^���(�����b�|8��?�=5��Z�IZ9�aa�N��O/�s#NU�bl���:��F����Y���H��a�t1�K0��"PT�wC����2��e���*F��%K2u�<4↻�(�ET��M#s§ER+Zr�]�'qYI��Y&���:���ꪝ�*,%B>y(�Ú!GK4¬�r,#ȖWJ�j�y��V��%�'��M�D+�D�|Nx���VUG�wЧq!�B"%	i��$L^t�楁BZb���E�H�-��tWwT�$�Y��U���B�L3Y���w�P�3�A��J�7��x�dt+�vG�!�����4���DK+ff��]9aP֙���fD�d箎n��S��JA��Rs��ή{rG<�q*�""�����֙�RD$SH��2�����e(�Lɠ(�Q$�M �}�{��L'���f�BJ�}��j��O�f�Rl�OAO>�mJ�`A�7�e7�>���
5[�f���l�[1���*�c�nd�>���-3�%��=��Ҋ�Kt�ѭ�E�,։}b����e@�z<��9Ӌ�v���f�Ux�
�]�^>0�=���eBٕVw��pS!]~w��uM�S���{�+��05������_P�bb����v�7�Y9�u�Ȱ�K�=R߻o��Gk������p�~�o��[��\�t�s��ܥ��u�u��׶4�����x<��S�g��>�$ܝԃ����> ��5�u�
������[���3��k'"7I�
�x����������wR���AE�z�c�1e�Ȑ�1�	���o�V���o��v���-�9s�����.��/� =�p��jAtXȊ�HD�s;s��àJ��V���og�֝�O^eI߾[s<�}S�_��|�uH��b��_�l�����ָOY����0�؈��=^�^��c�5J�s�R X��_�Q����A� �kyaJœq�ڏ���h���^Ua��Lk�{��C���^F��1�`�� ��B»����!���Bab�N~��rݹi�^WM���R3p�kKs9�u�^�j��yN9��fP���=��],���ryt�'�`l��ɸ��P�ӧt�%2��QpO�W�ݣ�]�C%��ʸ�Nd�#�v�O�z���Y��3�yl��E�ŏ�������tq��h����^��� &�Vy���Ο���l������5�F��uL�t�_�*�������Rc�*������L��t�K�_L��go��j<��v0U��|:^?�3�A?j��F�td�nH�Yp��ڱ���;��O�w�u�*C�q�>�d�t�B��l)��^N]qW�z�+�k����Ǔ�����7�A�x@y���*�E
���W�����!<U���-�W�ܹ��|��	d&��N�y�K�3*�_{��"ꖡ�@Q�(>ykS�S�O�w>9�{�l�Y]8�)҇�%N$�s���X"f���X���A��	���N&�
�������!���v�]O{9����*�9޺P���l����|f]>���9>�K$W��T��*���`��o����hu�>͵RO��9t`d蚩nX����/g}m�ݍ�n�uU�B�q�����G�K�5�O��Bk@�X�됙5<d7q� z٫�0-���j5Yti(��ƙ�'b�^��Iw[�Zc*V|&�:!7�M�x�iw�ﺮ����F�hU�-��HoA+e9��H��'������VmoT�l�M|���KR�"���4�Y��H�"
�Ζc�V�;��W�y��)zz�ͧt��(N��xyo];��隯iu��e�r�� ������=ڀ
dz�^�����;�������#��K�n�4rj�����}8�B��f޹�;w � ��_.D�r�Ca^[���To��sB��d�b@U�ǰDz	y��z�'��$�u�~�VK6��>`�L�eQ��ʎB�lMd5�z��l2�+�2���k;��N�;D��T�4����w[��Յ��_
v#�Mݮ�c�-o6q��zD���rϋ����?']A�E���-��^�T/FT.�	���؂������.��x_����� .���#�t.�^���_ѯ
�S�5�r�u��rǻ���Yc�3-�{#yS���+~
h.��{��J�a�ةa���lO3�
��.��vD'ָ  �)�V�/����X>J������a��;B�Ⅷ��R���w�	Kcf."��y�&������1���W����5��A��=0� �L����]��sC�$��1N<oV˺��x�S���|%�y��
R,{Ȩ��|�t���깫!de&�{��,}���Ȼ�K����:���BP����&�*�nC� ���7�v�f^<�����7p�����9|���xI��+/%�����c"�Ą4	�̽�k�*�?��п�`������q_A�� ���Pܱ��<���cN��%]	�q U�Lg�
���½+<.yX�����}�s�"f�Y{�˦	H�}�Rϳ�I9�P.��]yr�嚂�����k�J�=�z�z��S� �=x��=^��=�:�\���dC��`٭25�gpT����.����J�#1Tk"�fz\�	�9��\�u�-��7]؝�C��P�-�zP�ta��q�]�N�p��g�q��o?<��C�j�@�V�so28��#�L��1���zX��-C��*����@*�3��Z�yr6=�K�i���5���yKŴ;�{��r�������JêI<.�[q!ᮧ��r��/i�EK����:�K��[��3�u���.%�[t�!U��8�uVSI/�)�����a	���T�l�j���ߧ�c���Wzg�O���*Ώ
�������A��V���	�7}���G؅�R����<��ҍ ag���}�97`"�)�1�r�����m#4�`�O�(���K�KN��F�Tg}ݧ8^�����~�N���o�-�� iP۸�W}J<�=�Q��nmJ�7���SI�㲳�v� 4��R��%ݵR]���uB�!pc����Z��E>�4��+k�P��������Mos�N=Gޫ�W�4�lR�N�1��ut�룏Ͱ��#�*��@Wzd���w 蝀�Vz����3O��D믆Ď`��!�w�����&cy�\:��a�]�8N��n��_!y�O$F���`p�'A�p��dp�<~�t@\�C��8�"l�"��,��q�����B�0�׎d����^���/�������>ad�>������j�0ꮊ����4�s�֯��:IX�B)�;��.��P^GG���/_f6%<Z�6�+6�oUL�s3�n�w>}`�1`|��`�5�{:�^mn{��~^���sC���pcş;�#YUs��]to��/#�:�b�{cH��m��G�7[j�r쁼s=E���\E:�76��k�9
�g��vX|)�ｶ�����	�b��`ԥ�n�{��9�Fn�DAPQL�������٘/���Ԯ5����z��1��/&��on����-��Lu�"�[���c�Fq����ʗ���0�{��n����߹ש�I��͙�k�t��n�5���x��o!�V���B`��L����7)����t���̍���u�����,�kz�����\�b��		�ow��ѓ��5�����A�xR�`A.@zb�^�6yO���u�g�TW.ov����bV2��_��͡����, ��έg���
%MFU971d8��/Z��*����.1Tl��֥0�C�Գ��Y��R�a�Մܺ��Ȣ�m��ڻRH���xj��w
��!Χ�
\Y/4V��+&�uJg�f�z�A�%��N)Vˊ��ꡡ�>�:b�#_Y#c��#k��n��<���1a�i(M��0���_�.|a��\�W+�(V �������UWx�s��2��O p��ٕ�y欿`A��_����6U���`5�r�r6�SQ͙Υ|�54�����5v�I�:Ψ��V���QR�᪉�����D$��L
������v��+7ٝ�Sz�9�A��|< �߃<������~ͪۥ%0�%�ɍ(F�|�嵭%��3�h�� ��@g\^A��C���G�Q1!�00��5S��{�& �m�o�9��hR<;��+2����vo�s�O�e/W�F�r^�0��1�q
Ӿ�Ii�L����~]�;�������;�Զ�P59;4��<x1B��+wT��\|i�{��T7����Nn���꾫Wի@R]�uv���,�����l-��y��^u|��>���-�u�f��h�ܝhWR���+C�=Y ����M|)��> ��V8O)u���"�|����:�;qr]�sv��u �-�ܣc3e�f��$V��*C^ƫ0���X�x:�WOY;��s�v1��s6�64<]ڹ��E��蒥�vBK{^9C�[g�)T�x�k��/�`�Zנ����=��w)]���z©��A[^�[^m;��{Ł��$ �g*��nc
�Uz�����2�Sޭ�{{�ąSq�߅x>6<&w���g\GD��g�:�PG�w���S�.����*E�{��f�^x��u��k�t	�U=�s��
�U��n���<V$!׹�D�I+TK����=�T'|רo�+rz�J␇΋���kb�C�S���n��W������L{���N��|֕�pO�*��%���^��~��O��|`�!�Q���W�_>�����.�G��a�[���P�s"�ip�����Y����u�/7-v���zz�����ƺ����r��o �T����}���\��/S.�Bp�W`bLz�:�R� �-L�6�����7�{���s(L�WC!s�P�y���U��P;&mN�ޙ\��+i��oQ4������I��M<����s�Wm��g� ���x�|�� �D��t,5�)����y��j�� ;�y�|�-ӓ(�����Iّ�<��Z�J��=�Ā�;�y�O9��-���ۗ��9��s�]d
��y�&��\�x���|���t��ZI�~�)�5%�al�a���o �S�����Xl\Fm	W����0"58�q�i�0&�2�D\��gV�׻�mDN$Ew����H����k�_����!�q�I�r��ʥ�L�&�Y�iWqKo3���M�[��}K,t�U��8�.�
����(�M7a������߻{����s�������!�mU[U��;��VIuf��.�t4o]1�y5_N:^t��[V 
��^�h��\_���k��|�(S��+��c�x����c4F2)�1|��-@��b }��wHz���ĸVv+�^U!c�0g�!�wu�+`�6�ډE5O{�$�y,����ӫ�`�}�Yƃ����^,xfϽ����0_^t>�.�%&Q�����|�P}T�cqek=�]���2����g��:�w��:��	�*�P
��!k5��s��ð�j��n���9R/�Z��;�z"����]����8r�s�ξ�F��v�ej��n�8.M�oy�'S�u��soUT)�aB�e.C�n�xu:��x�kWN;�U�ƴW�kso��a�#�-�"���cZeWE@W]r�񿼯�Қ]���ć��s;��:�މڐIy7�ZP��.�׹�뿟��Y���T�=�	����Ɯ���v�7���g�&.�/9:���d���\+>�n�2V�����¡<��Z�/
���:N�)����ot�2����fR��E�ɸ.�O�	���	܆�{���i�F�<w|>�o�҄�3�k��������*Ȥ�{#��i�/x��3�n�1�PBB��+f��@�?~���� :9������j������]�� A�.y�+�����]q�}�{�7����Kɝ7�}l�{!`pd�!&�
�\=m�hO��	��G�n�ߡ����%ha~�* ��_���������9�o���4(�F6��g��p�ͻy(L��[��am{{3�h��~��!�P� u�����ĵ������bX��8�x�M�g9~">�ȹ��[*�]o0G6���������2%8`ǀ7F葐�����^����D��i�ZXg#�X���3eH�C���WS��*���͐���|eZsa�	3U��)ĥ>��+AɻY�pT�i��W�+$3�2�]�E|`��ݙB�Z2��$��lE� +/}v'�FyS'��v|w*�_���;��7�8�$��fp�SRӚ}M~������S�z5��#��]@Ƕ$���+K����#u���z�F��=z6Z�?].P�me�����^x����{\%η�o�A>2�&d^�͏g��$⨉\kaA�O���D~��o:�?Բ��L�_QiR'8�������m��F	}p�/�����p���XW=��| �Y��8�4�u��N�=湟s�4_���OrV=ew�����C9�N��PBC~Y��DR�*��v`�M׮��/�'��[J��w\�DoT9	[�ë�r{�[�=�,F��5�����T�9c�ֶ�d���y��]�;0�d�3逇\�b�.��O����^�=>�V��nĉe1�E�-%�8B�T�)��VS�V�a�Yg}ܤ��������9�wI(�n�Վ�Cn��Ԁ�����`� *6�����[,{����w�u|>��~L������JM9�1)G��N��B��|iS	�"��7{�����"�,wR}Ӭr�Ks$�
U�
'��V����8N*��MO�{�#LǇ
�m�M���`uي�<oq4�5�7:�sת�6XԷ��I�G�-Ͱ&�@�ֱ��>�)��z�q-��w����;DO.�k�p;# *˜��Wص�(�l�;���Ӫ��'d�986��p"�3p���q�۩��<�q���2�樊 fS�/Ivu��R�߽g�����K�b޼Q43�C���O�.�o�,mN2棵��[� �7��	�iɀ�[����*tW�*Vԇ(*1�{�iVL&�SP���M
oE	�nǅ���AwX-7 ����IJ��/����޴ot�ژ�

�2�m�Ӹ�0�H�W�M���("�P.@�����A�H�'wo^�cZ��t���0�.^�|z.����������q�N�ܬ��Fd���=��jt/7.)Zۢ4p�{��1�r�:�ga˖�gQf���%�;���L��s]ԧ�m�'��j�u�$��
fw�*u�3%rIuu���1�����Zՠ��/�\;�.L!u��]]=� F>����y�PTyC�E:ч�w^Z�f�K������R��[[y��A�>���z��ĸ��&���[�G���0��ר�8�K]�H擹W�l�%��!��|ŕ3w�S@]'Crơ�%��������Y(�:{U�n�h�ȁ�ӑ�yL=8)�,�ۻ��d��.�&�.�u��z�l�z��E�	Y\��t�^,��nRk,R�b�����.=�Y!*�,M�W��\�$.�ٳ�3y�t��{�C��=ڛ@R�(�����G�!��{F�����fm��b��W-^�b8�L��#�"�B�>��E��$���h-��O!v�>�V����rƮJ)x�.��F�ķЏIL�워�`�Icd���u�y8T8�f� �,*n޹���g+wך7_�M`��5��$��ڇ��;�ct��7�3��v��'L	@v��q��Q*���ON�i_M���<����\7P�m�n����?k��-��&�k��u)VːG���y���;�X!��X��=P�4"��n�;�-�L��rVŀ����]r�ݱ�(�J�z�I|9�5�7r��U�rR��������G�0�ά�]�L٧9*�O
Pf�� �C*T�����[�3�[�ܴeY�M \�+?��;A@��a�}�7�Dt1O9����݄�P�[7���:|уgɡһ�ƴ��3�AVd�n𧴆+��D��q��24��c���J䈼ZK���j�E��q����;�;KOT	��яr����_*w�a3�h�rN'!�����6գ	��J����Z�z�F�>��y���C��
�/Es"z̤��ww�8����lR
4	��Ы�����čE�-�+���曻�^d&Ri�2�#.U���Z�W6��)YJjt�d���,�e;�z&D�,��J��OG�病!�����v9��0Βr<��m%����F��Yy�p��J]4tD�4��If��̥3i�O7*�F&��30�aU���9][��.K��ssX���U9;�������*9��(�I�r(�Tb�y楚 dYU�4�J�u����gNQK]R3.b�P���p�N*��&(�g2wqª�Q��E+
Ts  �a��A�9fDFЂ�sK$32���܉�50��	�DY��H���q�!0�)-�$]:�\��$� ��spB���*Wu̪̣$��\r�J'w<�UV�2�BI4��*�̺�G9s�(��8U�J��#�-e��͢Tr�(�	,�&V��(U@ h�Ĺ˱�oz%mt����v�T��WR}�u��S��S���}Y�*˅�S�E�*Y�4WQ�8�WaJ��p�^a)�}���]}Ws����]�N�O
����ǈ�'�97������o�~�z@�v�����ݷ�	$=t~���i7zM��;~���'�$���{�r~���12b��t���z=�{y����<}�~'*o�;���	�v��Gߟ}�����7����~�zO������I���@�7ߐs�����`��=���I�?S��=���*b#�f~S	Nf�0j�"���l2�~����q!��}��ߜe�Cێv�������[�oa���N��u?�}�$ߨI;������18����'���>&�˷�һ|�����_hQ,F��@F"+�0ԏ�ۿ1��ORݬ�q�~�#G�DX����>���{�'&q��M�N����>F��';�O�v�SӉĞ߯�� $��[���ՂM;Ͽ;�������g�E�}D��/Ա$��JLH*�O��@P��>��'�1���7�{}&�B�o�ݷ�>�����O����=��ǧx��_�}�(��9wϖ���t����A��;xC}4>�?}""�#����^C�y��%�`��H��"�b�E�DA�>��s�N{O�#����~�I��o�����9P����������#��/��m��O�������6�[O$+��T�U�_,4���Wz�Ss���,�[q">�g�vL@��(DE������=;���&��?�9%w���x�8�C���=G�������;���~���ސ>$�ף�מ8�����m����>�Ç����g�^�S{�9O�B��XB"9�>���]������+����~'�~&�߿~pz�c���!����}���aw!��������aWz�?�7�oX������?%�N'~z�������e����k�w�J]~���1���L��$��w��S_��~|��=8��=�	�}��x��i�������~F%v��~��o�sɿP�o߾��������8}�PW��}�����)���9�����a���k�^� }�G�P���>�;ݲ����r$������|��	���zM�	S봟������;�������=��zO�ow�k����<��9S�����ߨO����6}Q�����+Enq��+���t|����XZ�7~=�U���6t�qY����a�Lc�m�8��R���bG��!�P���O�S�9˃iM՝[ �3L���ˮb� �.��|�ˠ����u�ӧ#�X�LO�'/{����Q�j;l�X�����|��N=;������<L/��=�y[O�������M��~��=&�|��lr�?����ӽ�������= }In��<쿮=��_~��`�隘�?ELO��μ:�=�պTg�꟠;N��7�;c���ޏ}���]���q�G�e7��7��v���<������������i���>yݷ�?������ˊ�R��n�ۧ��E��B�M���I��!�=��y�7!����:� |I�����x{~;r�I�z�x��'�/���w�o��=8���n>'~\aw�i��{��ğy+n�	�ԥW�e������B>��<��};��bq���ϼ������_������;�ro���PP���}�&�ˤ���������Bw��?m�����x����^F�O��"��r���{�u��=�%,�D�?N>����$�v��~�}������~~��ǉ�'�=|�zK�bq��Aߖ��O?�~q�j���>�;�.l��G��=&7��������H��o'���13Z��=ۛ��@~$�i���oI��C��7���9��u��e�������;����}��߈$�i�}��z��I�O���������~p.<I7����;o��� ��P[�=�u©go3S��rapL�q����a��X;�Ǵ���߿�x�]�G��ޝ�Ǵ���;���I�!'��8?c}C������1���'}��'�� zK�Ͼ�ޞ~���B�-���}�������_�}��v=8�N���{��0������������[շ&��&�����F'��w�]�ra}o�8���~8�}NC�F�?S�������Oߵ��t���� u�p٧�"���DDH�;��x��-��|���nBw�N��o�!z;���8����|I>�~��I�u��O뷟�x��S|B}�[x�y��_�|q�m��<M���>��1{n��8R�\�.~3��������0�?Y�����������|������ rN���}���=$��$��ɼ\~��?=X�I��;�U���>��_1��UW��o��K<�� C���I�q�f�Z�	�cf���E��Tƀ�"����q�)��p��	�j�&�{Y�w��r�4R'�
�N3�g�JeM��U��&� �������}���)�(�SS4*:G<�ܢt��G"������\u$m��j8�S���>H�ޮ��e���G���݂?bf����(C���׵bI�{��X��ױ��3X �p�쥹.�~bo����}��p:�F�w5�\:%����Bw��y�q)יx2��.�J�{ЂV�}�}��L`��4z��\�v���[�U��[=��?*���2��Ɨ����ݒ1=Q�����X6�q�Ǯ��]�_��V���6�����-�v��IA���zz��"�t\��1]=�pG⯋�b��<v���΀��<?�Wo!�a�'�oX��C��Ҷsd�[��]{=�i�4o/��+����W�
�&�qV�]��|��!{�����QC�����yfr"WmS .�UB�9ƣ�������͎*r=6����.4ja񫛌�lVB7Y	�s��>y��,���W�S7E)�ų�bn�>�����^`��
`���y7�)�6P�w�>�;���~�F@�WԆ���V�0���J����p@xo:�58��oEa�t���j�y�2��X.���K�|ll�n��X��Ac^����Z�f�}wZ�,�XEe��ψ����Ƹ��͓b� "�'�K��n�Xz9J��WR�;�ܜ��j�5����*<� tѝ�n�=�x K��k4AW�)�}�����-�*󹙢��_Єq
Z���l�I��iȎ��p�����>�6��e�� ��4=�m�~PA����FHw��]�)T��Wwu�8Uo"�J�w�� �CMv���,�<~���A�Xng�0��V��j�k��#d�v&6f�N��p[�8P�](5h:�h�v��@��!{�G~�`f�绱���&�����C�^WW�f��s�t��LK�:9	_���hI�=z�1~h�K�=�5�P�]�Q^��Q����g$/�"������xHft�%�6��%D�s}ޫ�}�ͽȺD>�E������/�T1�96��͹�J��A�]EJ��Q��jn���a]�S����>Ϗ���O_��E]k���>���=���۩��F��ܵ6��/o7z �x�X{�tFd��ƶ���>^<<�8<4�8��n��s��̚���u���_vj��Pc�ndZ`��:���Jj�_g������o	��=��u��K��q�L�ϫ�!��^��|��ʓ�l��@���:��dP���[7Ϲb�41�SP{���\�jwm��6�>"��CMٚ��×��#{�����,�h�{w�E��X���5u;��ɱ�RvRY�b��;��3���2,���b���[�D��زv�ξY��0�q��*��A��!�7V�R��e;u��Q>��R�P��|z�kUC�%nS���oԷ:rw�i���}wyx�'�C��ޣ�V��B
h��7B��u�vg.�g�xf����x�>څ@x���Z�D��]ͥ7 �{�� �~Դ"ሞ�H��<�ܮ�b�ZW�tBT�?`����%����-ک���k�3�C�s7k ��]Z[Ɲ���w�wZ�\�nk�����3��z�@#&��͚8�
΢�4Y�,�^�Gc��p^�cő�ٵ=*q����vƘ�Cg@���ԗv�,�U*n��h/����{GO@w*r�u�h��~��ݠ�Cոy�*�]j�����"�x`
���Y伕e"�v�������x\�R�y��̊����hn�pr��_M$*�x�9���~�� ��0=ɏ#�^A�,�
M�k��ʊ:0D�	.$џ������E��!u��0Е:�	��qíit���O>ѽв�f�U�vF�
��`���<i�����lpg�:�� �7���6���K�y|�7�E�2��������Y�0���b�\��2m����`�Q�/s];Ɨ%{�gS̆�klΡIDin|V0���ճ�VlC�ἦ�\�g ę����3�����Nm��K%rT�jr�K
�K�3�*Fl��.=���l��;���T�Nz�1=Ѥ]d�ۯ�k��f�-WD0�:���roro(�ћ*_���*�|�R��������u�K2Uy]43�謭���`ns��B�W:�3lr\�D�='����:<'�y/a���3�.
���	�����Lf���K�+N\uc�_>������D�D��AtP���W��6<&N󂮽�q�g�L�,z:8���Gv)���=Se視fKh�ʧ����ל��{�x�k³yT�s��JDZ�q	���pO�>����:���(S'z_!��+]Vy�*��\k������u0+m�����fy�΅������6� �J��J�8'֕At��ޔ�ゐ^�X����1SԨw����f��W28j��� ,w���>�W��D�U�t�a=u��y�O kj��1�Ӥ�C}ylh��gb"x�4�yX�μT>N�  �l��Q��o���h�^�ȧcsT�|�t��m����[����'fF2����J�����j��������s>���٣�$���Uۧ���3uo�?_�h}���j�AR�i��wn��4U�S��CF��or̲�Ή����a���d�c��uu�U3�H�
xr�r��D�&X�S���nu�3�"��s�2í�9����7��"#���5������� c5�9�ek�\�d��}k�'|����^�^o+ӷч�mt���x����.zY����_	��@�]���m	V��i>�ƺ���{N�>�ހl{����o��ͣ^��E�^���.l��$!=���.�5�)����[�hkC9A<�Vvk��޶�����h��g�W�%�TKYn��=�%X�N�)
+�>���m���JI�k;ZFЩ�0�+�2_Н\�qu��������P�}j�������)��g�]`���լ{��`W�߃��Bw��y^�B��p��&Y(������U��^����`0��^f�`<����/L�]OC���˔j3�o���yT��*����Rp8g�sdcӯ�i[8-�x�xX��_��V���7��W�q�Ñ�����esYg���[#�10�:��r)
+!���g:V����G}��y��P-O��u���\q�g��?n>f�����~W�Kӕ|������
W�|v����+�mN�H�4�X�5��S��V��H����*�C!��F�kB�݃�l�R�{�"���8�*@��T}E��]���Β����gyP�4�o{U��u�h�*TS/"�:��kw��m��h�0���#�MgE����n\��o� ��w��R�3������UA��f�b���}�>��*g`=L�ի�$��"���s�$+��,��9*)�|��+@X��ҙ����]ܯm.�Mnno�tz��CuVVq��-^M�]B�#~]Ba�����{�CՔ��e"�'�ރ{}F�E��f��*��Ne��q~��E �;��l7Pf�z�(�w,K�6��)�1Wb�=�,z��:n�Ԁ��@��B���!�f!n;���K�����Rî�A�b<������uk"�>�Vj�K�B���=
��;�G���K4��+b�;���p|�X����a퉍w���zߑ:Q=�|���QV�p:1�����O�z{=f��"����^D�u�:�^ePU�����ĵ�������[Y�y�w+yr�M�=������XcU�y�]�`y�> A��w;�ܑ7��>:���	�f��R�h���>�z���A/�#şc5�4�\�>G�^mR�Bro/���z8��sꜺ���٫��!��L[�cF���=��v����P����nJ�,C��o9j} w�M�u̷Xvw�m����)J�3w+-���w��@�Zl��q#�]���ε$Lѳ,��:7]	y1����YAQ��G�=e	\���oFɟ}��P�0Qq���k0�x�\��z�/]prR~��vXP`�M�ny��p8_jD^p�{��Bïv]�+��Ʒ
Um]�[<Vt
���3��� 
:�K�O5���w���V����8w�v�F���8a9�+�%yu�e�ۨ�z��A�}���ם�oN��ש�vkYpZ������^��|�]�����٩�㜾�w���� �l��ztu4{�Vؽ���*�j5T9��Lk��s�Ks��{ר���p$��1zS��v�Ƿz�4O��:�Hp�4o�
:v�zع�!S�:�98��s��po�w\ �tf�t͉��s}�dV��A�y.�Ù��	�ia5<�>��]e��r�>�<5���K�!A�����˞��b�����W�a�|\�@o?���]X �N���pU��-�d涤^O$��2���Gdky ���U��u����'��w-��x4׬g�%���E�<r�=��cS�R�َ��F[�|�l1t��4'��ӉR�P��!�v����nԴ&/2����e��&
���\��/j�_,�
�-d����[�JBvJ��S��+a�$Tz��u�P���0�u���x�sgf�"��:�{ḋ2�����yn	�� e���X�ݮ�Ȭ����X�i���p��;��}�D}Ö��Z�ފ�ɨ-�\�l?����zq�:�y�k���Ev�F�{�a��?B�{�_�K�Q;�Z
����E��x\�`o��׀
@X��J?jz��]R):���=T{01K�(ۯo�;دu".ۇ�B�q�_0-*q%�P��w�e�[�Fqx7�=��y��O39�!Ws�=��b��d0_��x�*]���z�����8.�]�e���n��J�_���v�yV0��qZ�<$W`�1D�{u��T썽�.A֟[=�)�]p����ce�kog;�u���b�/3�ϻۻ[�섖��r�
����PKW�m������n�t�� �̽�P�nK�c�|#_VI�d��n�0O$Y��],��]��6����P��K����Xz�t$O�7��¼.���+�����г��hw�e�>{�s�Nީ�l�b�Z[�ыU. Ab�'Vs�����=���V�[�S.3S:h�x��[ZFp�B	���so���T'z��
�ʪ>�t���T�L����#��tȺ��% �u<���U��̷q�\�Eu�.4�!J-�wn�v�A��k��S�P/\sA|�+z$�7!�_ �bL�����[��ۘZ�Q�7;�*tU�r����G���8��Dm��W��<��Y8HÃ��0wWIE`��_�u�O"�7��X�Քv=�o���:�9Ͳ�,�Lx���v��7RF����4-`T!�>�B�)u�3��%R7Y�q��|��{�X����/E��Z&��S9:��S5��yh�G�'� Պ��x��\z�}G'a<��ݧ��k�G%�buWY�vqV�2���땆l�'R����ǌ��,
��=Y@q����}�s_=G�Ԯ�%]G\;�,a��˱��y��B���Q�k���]�boV��MM��ANŹ&�u���P��R�
�\�6�P���:���<�#��.f٩��Y�w�v�li�X1��K-�
��.�S���gdx6��}P�]ҁ�a;�4��������%��rt�\�'��&�)�����-��X����@��X������hS���]���V�i��2m&I�f��]�v'\6���#ٓt
iW9�	3w:QCD2?����|���ì�k�t�0i(y!��K	�Š�
陜�o�!w�k�0���ѹ��X���CkOe�{��Mʟ���x��n� +=��9꒓�����sSy�u��,����K���̓k;rZ���!r'WmU5s�m�7�^P��V(�`˄l�kt'?&�:䫷*��	��t1��LE����ph!F+$Լ'zV0���B��w �������:h�!�$��Nu���EY�}���|�\i\{ZZ��E�W\@8����ۺ9���R�%�ڹ÷&K'(�a� [9uJ��8T�Wnct�dx;��cE�r�<��:9�ni�힮�7z�M�.E:��\��i8��
\���׼�-ڥSk���x��m�'U2�������a� Ԯ��-�K�ݲ��ju��T�U&Vd8:��{K��W09ֽ�hK�o�/�S+fhG�a�\����DQn]���[�wi������	�N���94�ٓ�S\�����z�gM��)=mՒ��I��{YM޼��X��\
Ltoq�q�K�.�U�{h�hɌ$��o6(�ʰ]�
���V��`��s�}M��uӬiAB1h��Rc�  ��鱛�!���o����͔8l턓��V¨PL����=Y�>xj��U ĭ��S��8��E��3Cssn����~��>psfp��9�tS�^����b+C�&���|�{[;�>Ҳ�+wk�s��/	}�jp�&�aJuWN�ڶe�e<A�*}42�)�씸Z���zp)v��bk��ñ�yն�Ā\��t#I�^�j�T^����]<���u;��fMӂ���v�+u�Վ��ô�#!t�����n��MnP(��}n�r���֩�*8n��������A%��$*��DUe�(����,��6+8�bE�J�ES�B�X��jTj���YlH�u�PШ���3(�#j�T�LR):W4�T�P�E��\��1*,Qa��C��3�-Bi�!�*�������*�!,�T��R
,�Y]X�*U���1hW#B�T.2�͖(vDJX�9,��J��������H�d�	��B,ʹ�3YAV����QB�J�H�G*J�4-0�X�QrL�I�&�RB��*�&�r��E��$1,<�4HEb-D�H��$,��9A\�$���ЮDbEB+�U#&UUQ�ՠa�&b�I��D��jd�fPWDH!)"ŉ�3T�
�%,���"��1:�E�Hꈣ*�Z�E$a�aRt��S�ʍL".h�¤������e�2�N����D)F�Ě4��a]Jȟu��G�.a�2�^��_~�o�`
'q�f��84+��J���"�r�J�ʚ���.����<��4J�������ygW軟^F���|�|sϠ��m��j�TV��_#c�ñ��&S2%����j�f�����{q��*��#e^/�_ΔQLj̜��i��Ȯ��F�Iu��\W]iO���x��\�����]QњW7�C�t�w	�y;�uz��c���t�F;=����?g�~oɞC���G*�Y�ˌm�i���?��S�Я�����r��O����<{Һ�֣鸲�%X�M���*P����Wb�/�DF�;��[|k����|��fz�we�5z�;�a]��J�b�3!�joో��/� �r��������׉�|EE��Jk�s%#8B�d\CN�+l��j�؀�_d@^��{9����'�rkBo��>��㬋ͮ7ޡ�����[~�%���w_}������8��L����HnN8��)d��KC���7��<������^�~����� ;M(x'!'�_L�t*p�X^�F�(�w��w��h��T����UJZ��/!�[�'d�}{��V�Kk��(�����L�ۣ0G�@�&���[\�A�p�̷���; 0�ru�W�se����jx���諭��7Y�Q�pg��NEn���ۍp1�Ҳv�������V�.M	"6�ܴ9�u�T�Ù+�A����5/��:�>�E����%saI�����1�oJ���Ti���X9^Oj�u�1J��:�ש�CC��Fn�N��/>�w4:�}�����U�2�vC�2��U��������ro�+Rr�����[B�a�lZM<uϲ!V]���ʿ�(�
�����r�;���������Ȱ�z�B���i��<O�W�eK�=z�-�Y{\r{�B�l77��{���:��mqߗN��ӭ�y�w�r1�h.s��ƾCri�������Q����.'���ڸ�&�3�=�Yw�/T)��l�<���7���!����՚��V1q-�!ǻR$�W�[��[ʕ�c�Gf�ؿ�[���U�r��q���E���^��SN[B���h���*�Y��&�gV����@=���:��������[��]i�V3]�ô�ɔ�;ܭ~'�j�b�^�!��܎�y��^���²_r.�+NP�K#;Ws:h�tne`��ք�+�[=��f� K���96�J�w�}�DG�<qC���Kn{��P��Yk��lRx���R�!����MXP�\S�=/�7�>w�T����Wٜ�_'�Jا�q_5�OT�q��[0e�~xgmb^��2SԊ�9W6�Q;EV����6WPXV_t�կ�%��&m�쇧�g�������=����ض5�2�r�͹��5�d���������3�I�K���N򨳯O@ u���
�+׉?wC-����}�~�6��zew>=�[�N��|��T��t>җ_�����x�l5�~�=���K���#��3��=W&�{[Kz6��u�⋋�d*��a{���5�nyq�d��Ym���&='�z��C:��덥��bLZM6)3+
KGb���d��6���`�N!V+��=}�K�E��w� ak�����J.��Ud��7.�{QWt�&������ς��z���gϺH�^8�l��RP0ִ�7�85������C<��..���=Y ����ʒ�,���fs��܂�	&�s=gJP<�8�uWVV��77nR��t0���~�ﾏ��]�)IK]rݻ_��w�˸�J(��"�ۊ�>̝�a�wG�0&L{{��/���9�x\Fq�������q��V�EK1Q8���Wٞ�^M����}z��7�V=����؜�W�K��.ʎ����L����nO4��
\�Y�E8�'����JHkwn��W�W-gѢ:*+3������0v�v/����n��wʸk��KبN�XT����Z��ŵtr�[�F�,��*������-��w�pq�ĭ����U��e�j�dk�i-�U��c�Ⱦ ��5�C��N�U�^ʎ��D.9B\^�qB�z;�--Ү1X�Em�;	X\��Qy ��R�p�:s�e�?8�,�D坞��s�ޯk�/�V����s���h�H���^V��q�U�ʒ^����e��c�ډ�3N�>g�'���wOW�[@(��'{ޥy�؂Tӫ/pv�[KoO9��{'\B�N�v[uj�w��K���k���aō����_
۹�dɧF
���qt�V�P4���:쓶x�YF��կn����th�c�K�	q��%���Ҍ ���஁��D��G�DG��C/���}�;z`F"�89���}{��l��$PU�$�s�݆z��p�p��]t���Fh���rM
y���<0��;u)n:m],����[�R���
�}�7�E���rn��U�-�[ԜXVYp�t�8��V����L��V+b���3�T���2���u.�y�1��8nO"k�C���:O�y��M��ʔTV�P[qA� ͂]�H�5�iq�\q��oQ���9cyl���_r�J(�����:���U�n+y�#�:��C	ȋ�w]u�����j1�ۇv���q}�"��{h�3}�������}s��jA�O#�ٮ&�)37X7�u�X�xվ��C�ӗ�V�B�i����`��DP�Eĵٲ�k&�2�r��蝥�i��92�������ܟ��G�K:�vC�/�@�j�ӯ�eR�4 7Fh�Q&����pz9��ь@��&�a�b�]Z
͜*v��|�%����"*o����o��3���g6�T�ړw�WX�ᇿ�����;�eG[���!d����F� �c�J���G{h���-�<��#]�u�:"BeҝZ�f�;����������<��jNƟ�/b��61p:���;(�����XÍ���"���������dE9ޑi8/���a�cB�}�Qrs.n���X��q����s1��ۦ��Ϝ;��b�8�p�m�\e�>�)���>��vʎ���}n)��S��L�գ/7����5�����˓���prs�w�(,��j�ׇ�{��Ay�A�y'����3�E�ʑ1Uh��ez��;[�2��i�ʄ;��+Bs�T�f�������P�-^�p�NwB�/z(�����Z;"l��:ݿ��T4v�(}k��wp�*�2��YkW��L;/E��Y
���e2�w<S)[R�7��D��"Y��r�)j�-��#z1$5&�|�q�ϧl>u��u�겶��3fk��Ҝ��C:��-e�W��B֠�&����8%O�RC��u=����hB��0�JYz��q[0��n$}�o�G�U��̎���8Vmr8g7QXp��}t��T��ѽN��=B]�pJ�[y�Q������pȱmw�sf��������gGN�/)x;0	�������!�}�}_U��z��>�v}��_T��ۡ����]F����׏�[�j��4*�A;���9{���{�m���N�FQ�t~�<3��g�(�����(+x��M�p�����2\Gj�ۦĳ��uJ1_D�"壐���p�]y)3n�D�����ĳ���0����9���^�=�_B�VW���K�W@��֤���Gl��6;�����x���~Ty��C��ޝ���?pN���;��wo3���*��PJr98���^�iW�xa�T
�	<��'z>�����	�ئ��V��V��VT1$�M�η��`Ʈ�I�5ɉ'G%;�^Ov��v������ի!��p��۹�q��>��7��f�!��ޚ�� ��+��/����{�K�ٲ�>:�Ϭ�R�����{[����;��#�Hd��W�&����H{�}�����%�Zq��\�otM���D"�|8q؃>>�u���{����L^�6��	��R��u��VrQu�}]g.f����h��ŉt�tWS�`8,N���4��9&�+L뷶�X�|onI��79����Źّ٭]�	Q�/}���}�5a��Tǣu����p9�ϛ�{a��gt�d�3�WݯzD�����N�o���{+eC�o�|��9rB�iMTC׀�͞y��ϸ�����x}'T����
	]i���\��I��:��`-����z��wT�����d�=U���Ѣ��K�ά������>��8�{���ڝ���O��Z�ns�6]�ڙw
�QnP[t;�L�FgS�~Yz�s���{Y��X�ҍ��ۆ�6U�/�[��1�N%tD�W��*��	�^�c��G�z���s�q���]R���]����GTJ1CqSùƸcˆo�9�χb�ԙK7��r������aݺ�%o�\�:{u�%C�.���\��*���om�:Fz^�/�r��jv��x�ʍ@�ɶ���7��y����|(j�LƙU4��z�p�?
��U��v*qoe�]%mӴ.�^]�{;��3+:oZsÞ��q:RU��N
��M���9�Ǔ���P��&*��|��^Z�#N�� �㎕�#�T7�L�e�s�݆�e���s彛|B3�kn�h��ŞA�Q��*o��Y��~�ټN�����"ʾ9v��,G�Sq_7�,uK�����aߧi�/gѐ����瞍n��e8uOwC`�7N/�^��}���}����R�p�덒�bl�$��ŭ#j�F<.��[1���>�*�>�o�㻬P$S�];��M�n;���kh��{}�ϙ�\���s" n�=0ѽLB�����]Wt��n'U�N���[���x�'L�����w{rψ�Fc�3�}i�����Eȥ�TFj*/��<�UoO���=5q&��n�Es[|^�����������*;b�.����b,b��<Hp�>��V�c�V_1�ͽ��L��X�!�{�C8(�tw^ ���c.9i�p֮�\�n�hoR}��5�sȂ6Sje!о �Ϣ�֫2(Ÿ9�R��K�o�H�qc��z�%����9cfrQ��+t��Y�b��H�������-����8!Z�G*mn%���B��˭�5=��ܡ����q�J�B_m�>Dg=�G���4��a�k/�N�}��N�]?���*4���� ẜ������D����Z��uq�������F��ތ]�n�.X��n+��B�}��IE���Kq�g�K[t
Y|�+�J}����x��I�K�fajغ31t�V=�*wP�T5_��p��{�F7�}���$��=`�������������vr�G�)�I�/���(����k�Fl��5�q��Nݲ�C��Z�6�5&�0<�\V�^,���{J7�7޼:e)�zN�e^�o�Z&���ި��v�����a�S�w0���1�C�F6.\�K:�}M��u���~�jz��{��r�J��	��\�z��\����V�U�ڍ�W��хC�V��_���;/��[�Yx�Hq�w��]�Wn�R����jՐ��+>�|b��ř/�P�b˗�72�)�?V�qh�	cp�{;�7W��q�ߺ�̩�Q�5��:�~�=��ly������d�q�W�jZ����_`﨏���]�~������[���4�����utr��]o蘗�zH��mU��;mh4�q�Ԧ�r9�ouS�	a*�D++��qP4=W�%�ܠ��J��<�ɝ��a=ã0y�0�w;4x"���͋��ηkƹd�Dyv�3�z���+�MS؜��,����|�2F����ˀԖ���gM�����IB�	����X��G���'�)����t�5�tژ:l�aԤT�;��/��ϲV���]���;Q��ne�8�Q�7�Cc`�Ӌ��\$F�治_mvo�+"X�&R�PJ��9f
����ގjז�-ʗ����@�ǲ�ή�m���R�{��"���n�7���k㫎�ma� �,9�*�}�5V>Y8�&�4��:Y�
��Ĩ�1��L��[�l��frzW���g2x���χG�����p#��oVk��O��p3�(T�&�v��gJt,�7,Ŧ$��۷�Y;`���%i���X�e��eꔭ� ^��yXP�u��9�PZ�dN����;���Y�n� aCL�ز�V�vˣ��%.ģB�]o&lۨ9[��U�\գ5���n���ÊUr�4���G#�-,[���4�=��&��Yq�;l�����h���n�&n܍�p~��&�9}��՚�'����X���N,wWN^i���do��0��ÃEд=[#i�m�Y���3f��覉��*��;�WQ�+8qsd��D.�u�K��*�І��:S6T� ���Ʋ�^��a��[���B�[�f��+��'�n�G�����;x��We��4�;܅f+�w3�B�e�M�[�
쒩�)̀�.�K����E�k4��'�N�W���h*�a���KQT@-+ OQ}C��o���CFdqp�8��{X\E]�*�쏞ފ��'ΕqU�^�,�b7+�����bW��+16�87;������4'˲��<>X��:J�{�n]�Q�B7���nXfн���saP
V[�e^�5�)�r=�y�6S�9WIp�Q���q8�n�o���|���%,��r��O�w(gc̫w�ñ���aWl\��ԻA��IW�G_�5�怦�pkdf�C��[մ4�� �е�q���ŭF�@��|ܨ+�;2�k@mO�����B�u8%�)�]���ACWFpn�r1`�I�Wî�-�������pqw9�ڶ���;��۽�pd�5c�Y�L�e��3Q����ڵ�����a>\�� ��+��
8�K�5�J�����35]�X��;uε��\Ñ[�HP��mژ���s\�i���f�W��zW���{+b��Ö�)�5�YN��&�s����l-o9��Ti���H��%m1�-�c@�k�q�v�����w9�9M�M��!$�]�2�7Z7CF\c�-���c���M[���������?����"�2�QZ������Y��TA'"NG9XZ�J����H�4�tR��J1$�-Yaԯqۂ\���YX��DbU"��IÒ	���\��iG2.�� ��Q�J�KE�":��Y���E&�)J�E
��(��ȭ�&�R�,�U��6�F$Z&�$id�̥)-dEe	�)&iЫDDDM��(��$ҳ���Eks�I6��2�Y\�H��3�i$��,D��(�$$�:e!l�]VUR�E��&fdTEQ�R�dRl�Et�$"�%RYDZf�E�ʵh��*I-��Qr##˥��YDDZ�;�YȢ�Pջ�T+J�f�bhIEA�$�TW���.WV�H��(�UH�e�8jz�gT�HH����-j`����u4�ȫ�e֤Z��QTig+4ʏ0��r�"T���TR�#-2rU� ��X����ˠ�6�gv͔k�0h�V*��S1���g69t����L�5���)S;*ݨ�6� U�dΌ6������ﮒ٭庩�=�7���i�g[+Gd,�G!��J�����VU�����q���ًpL�P���[Ӽ�e�e\*�p�-���S�a�kV�k�f�����U�+D��B�H\$��\�>U��Whx�L��<�\ƃ��a��+�B�q�=h��-ui �Z�)����&/k�.�v�{���rq�[�v�EAM�N�������]F����w��}��������V�-;�j�O��3�t�O��)g�n�܃����� �)x���#�n!��ݪ�n��b���������h�M��T�컝}�=�e-�d�[[��%7�n���J�j嬈�Q/��w+]^.��dޛˌ>��]S��q�n�pnZ���x�����+�7��;�ֶ�C�3Kp��N�_���{�V�vШ%9�'䭊��qn砬v�8���sU��@�o_�{�K��P��St�s875Sٶ�m�3p��F��3���G&RT�*��팼
/惗�}�챻���2rf�=�{��zPLyݼ���C�ؙ�G]G9*TΤ����# ��S;f.����a��}�}��!ۗ�
쳈_ }>�/z+�TW��e�W�w�El�**��.g���.5��{��]�{]���n)k8^�mZ��ȓuO�4���t��oc-T�yS۩z0��3�OZ̍vu�
;B;u����Kԗ^�#vm�/!�:�g�{����5��>MI�W9��2_���vl���հ�	��T\Z���j�}�h�Nv߂T��h�m�t/4�׽=V����qF^�����$)�MW�^�!pEt�Oqe�z��ޯܪ���](]���#b�I���>��\ogi^�f�;zI~��>|��O�r�{���o����u��iH�R8��}y�-�s2���S.�(��
܊D�3��"ވ�Q�[�E����f��<_K�c��n�3��F/�0�bY���ݴ]��1{�v/EP�ǲ�ѫ�V��d��9�)�n����Ae��+�HPbv�[�J�%v6=y���/��Nẉ�[�ƽ����ާ��|[,�<�7/��zKòY�EP��"�m��cr<�5ӗ܅=qK��oW	�=���?/G��DGҭ.!�/��}}�]���wN���o�wj��7�]��j�[QdS����T�G�<o�wL���Z�ٸm�n���!ژ�J�%�������gQ�8+!�2.%�͔wY��S�WK�ܛP>��\0�=սz�x�ag�v����CWm�'_F�U�(�� �����j��7l�J�b���Ts������uK�VWe��j�ދ����YfD�-vNsXL�R3��͎8֤c3���p�m�����k�Ӛ�`S4�����/T�$��qW�kp�!j����q�>������q��v���'�;q����s���|�Ow2 n�W �Ž*����1=N羃��-/V{y���=�]��6��ʢ}ٷ���맜9��}~�A��s�����(}j���AeE�I���8n݈�x��VFٛӘ�����Y:��޻4�܌�\�b�Ԥ��em]a��Vh�y!�}nc [�|2�����ʯ
��"{������:<.���[�]j9��\��]�j��ሺ��m�J�O�Y�}�@�ޱ)��:��}a���Ɂ�Vw��>��V��UGN�Ư}����Ws��!V�mu�J\m{^u~��Z&�?,)�_M�p��o>�V�j����)�*�p�=}�WT�����;�l�O{���|���Ze;MK�}�*�S*�R� �ARp�*Oi���q��Q4��[0���\��6�wO���ϗ}:1w<�{Mj�]������m����C�#J|w�]:���-e���F[���o��CrkO�<��F+��b��F�)����Z��8�ۙ��i�]��|�e�UJ��U*����0GT�*"!�1���d�p	:�4[!a��T���se��ً���<�F��+ƵiF�'T��G��TI&��8K����Ǵ>fWBȕ�Q	ۛ�,b�T����J#aٙ�80��n�m3�=�����'���dd�󐓍jF(��b��b¹}�k�fC��"��<N�G:��~\�߶�]z�˯���$�Sۘ'q��16�c�c	=�+v��{`5��;�����~k]��C�G\��8�I�AZ�ulC�Dk��h��cc�:mcwt����37�&0�l�r�YKP����#溜���7w~�=ۮ�W��j՗[aP�'�:ۈ}9y�6�]V^�~�ޣ���1<��ӭ�^�]N�ӝ�ǵ?V�h�s�c���Dks�0���qkw�S�6ցkd��^��qOgn5@�et����!"f+S��k��f�u��<��K���u�C�Ϗz�V�,��y�w8[\N�Z��k���l8��oO5�����{S����Uu���#b�=ܡ���H�K�6��u��(�W.Y�*��y�l���L�U�
u�s�L����Z��k�J�qC:��	�h}�7B�i���ʰޮ��[�;rSY�*�u��`�O�J:K͡�uK�X�zIZ�9�f��WU�V̗'���1��8<���y���p���n�7�ּmv�9r��v��X��M���2r�q����6^/�vWED��s���mGE���n�th�R���	�N}��
,��T:]�i}Ϸ��������K����(�B��Ş����w�*�'�b̭v����,��Ȝ�u���R���0�)B����qr�Der��7�5�������Q�o��+FH��7}A~�����(r2�D�����܆��z��wj���q��uDJ1S���у�)<<s�K��aݿ�e8{�~M�_έՅR��k>�$t9��i�3O���)`���6^��g����9�	��m��`�ဖ\'\}s�'_e�b��+�S�yƧ�����0-��2u���sKjrF��|=�"� ��Kh���oi�9����$co����j򻹃��4��M<�_�R�k%{���=�ޮ���g�+���{�X|ъ̋ղm��k�3�<_xk�{u/F�5bg�~U��yG��q��^�3�ɴ9��X{L��7܋�}N�<���!�+�5U�q;��-NR�/c�Es��q�/z6#w���X�x��c^H�T�m��v#
N�d��.ا�7�:t:���T;�)����:r�����V}�c����E^�1� �=�$�.��x��99������wY�4?���=�o?B��gF^��~�[��JUx�����7�f�s�Ne��Q� K��L����u-'���ֱ�W�
݊[4�:b���ά�N�N薂�O0��.ܡ�΁ UG�}�}�ET��j�`��}��u�X&�(Em>��1&i��Ww'J��yE���������oBϞ)�j�Y+��/o:��u=~9舐=��$��r#oxqM=Ps3��ͩ�j�Q�ۄI�fe�|�/:�S�����o���f�N�7m��G�_r��(������p�J7E��	�k�ԟr��B��K9}9s�޺����j#��_{�����גLV�����@���˭��-�<���|.y��G�d���`��Ͱmݺ���U�Eʲ���N\�ϴGTD�1r�^l��LGeg�k�oQjE�@��Z,4��̱m��0eo���W�鸾]������|:��2n��v��f���@��y����^�: ����*v�ҷ1XY�;i�\^���q��YpŤ��
����U�@�+�T~��x��,�v8=;��?T��S�RV�բ��DCwtbL�y"�uKR�ut�ACܾ�da�uy����G�\̆��8J���֋'<.��k+����5��-�{ffL)ER�*'7�����ŐR��j)t����)�Y'��ꈏ���V����r��m[��o�1SS�|�.�}�T5�9\TN���XaՌ:�D��n"���f6���������ǝ�̷�_;�i�o��b�X���9Ռؾ��6s��z�7�R�쀨��^|�3�T�]�{F�I,���{�w��G��n���Ϸ�R�e��r�w$U �ݻL�S�t-E�g��'�����k��W#ϗWm��@�ė
l�����s\�ӥ�|����7��ot<S)Z�=}<n��!|�>��w2ֶ��N�޺ƐZ�)�k�xFʿ�S*�T������Y���b6��{���O`�\�����Xa{F"�@X�D��ʅ�h�Z���)Q���>�e�}y{۔D�,��f�}��Z�?p��Gj����=v5���i��}��.�v#P�:5jxT���ʾ�n^�ܥ��;}kw,TSp���J�pP_��e�]����f���������o	[�����u����s�ʒt��� �,�=���ˣ˼ٓ�z�D�.��{FV��M4��*���1'T��fN�R*��F�V����$M��vЂ��t�%�U}_}��nv%5k8�����7��T�+Z���R���m_�g�o�z���u��Q���+F_l�ƹ�M���[���.T��b:��#\f��a����29�u$��l���Tw#+!����̫cGT���������Ge�������Fv֬\@ز��I�yV��1�`�X�O��%}fKyE����v��Y��ի.��
�/�)�ѣP�kXv�b�����u�vݭ���jy_r�'3��]R�%�;ʢ����[�Vr�4.��5��m�H��"V>�F��^g�/�{�K?En������c+���㠪Uz�Q]g�ul�;=~��:k��������7�x�Hp��T{�:J.��w^�\��݂l.\�L=�5��\zڷ���{~·_8;����f%1}'e#�tqx�~��P�S��ӗ���e[/Gc�2��t�C��������v�6�6���{v;]i��,���ڀ�;3j�ʽ���vy���kj+�^��h�'.��n�7T$x�.��g���F��J�2<��vi�լ7��q�%��"�m0�KŴ�ni�i����Ĥʗu����˸����>��y�5��p�<���]�C�P1$i�Qj��>ә�]+�.�BH_��.�{�~o�R�9����U>U<��F$��A��.1R7AM��r���έ��L����WC�J����"O,��fQ�4^z)+rv���&��Ӫ���t��K����+�F3��b��N����k<�[B�l���$�|���T�;�36��p��\7R��d�lJ1N�6��9��.OG�7��[>��n�v-�!�%��M�[�u@U)����@�W�Ib���ެ�W�_C�;�ʓƣ��X��ylW��v�),�nMf�M�0��=�����n�E<;a7�N�;ެ� ���8�ڧ���^.����ן�^�j�%ev7)w������~#����!���V����*��1&ڭ������Md���c�v�)o���}UC�{�h��^G��ۏ[�ʆ���1����;�J�{vr�_f��ؼ1y�c�"�1CP�i�klwQ���i��xbA Qނ��@��ϟ}Նsa��bû��U�h�51� �^R�hWZP��=�!���v�w���[4AZJf�Wx�%�o:����Y��E�������m����Yנ�Z��quN��ޗ�ų��u�N�%��!��;1�桠(��s.IW|�D6k&M�}Z��q�]���RJv�.��0f+�	,���݀2*�~�-��r��|r]�&��FFm���M��ytqE��݌��V���%L�jK��!fe��fGa�J^I�w���.t�{9sB�/��&�oN�zfs��4��X�4h����t0�{�S���� �r[d�t�<��-�KP��n�k'|!��p���+�}��&H%f[U���Μ�CJ-T�(�Q��w[k[�w���8��pu0u�/������*Ze��(-�!����K{�*�eKU�\u�u+0��˦���Z5X��z��me�6�ِ�u�5,�3{]�1TO1;�L�ݗ���{9S�yʹ�$T��Rr2����8+H�]�&>kt;[�w{V��'Zо���sل(�=�H�w�ҩ�]\e������gWܪ�u�!O_4Z��<bkw� *��J!V$+P�����A�V���9�*��ӳ� )�y%�3R	塽�W�jGts��[c�w<���f�z	&k�M2Ă�l�c�V{*#�ePunÌ]�a���\hV��(�q�d� ������+еsh�BR@�o���7�>T���kΚ�����L�X��Ϭ�g%�2�'/��u����[X(:p�N��Up����4���A�t�*^�՘{�<{�6���ϙ1:H������v��U�$]�1�a[u�@
�%×�34�8�!Ҍvz ����s쇴��r���>&0�ڮ��ͤ&I�M���sz����
�-���kY�q�J%�
y)�$xi7F�f�uiͬ�lre̹qށ9ʓ���_-�.��,��*�$%�����򒜪U��*ww�[��Fn�gu*Ԍ�3{��9��h����J�\HWg;�zFDw��P�!6(aq�,���{�=�T�u�ظ���l"�^�K'�:�^Q��v�u%H�}��$z�h�ܴ�(.*��+1l�O�ʝ��;�3��6�"�Y|���Ð���>����w����\/dyf��ˆ���k�ɢ)��P��	�2����2�
a���9�aΒS�M�ق0MM�ԋ�U�30>��¥Z������L��U�\)�XE
�G�3��F�������ZQ�������I�����ܝ�!9ݝ�il��<�v9+����kK��s�G���K[m�\����u�k����#}N�\1��{Ћ�ʇP���r����_�����~�{����H��Ch��m)LĈ���5�좣:Ej��S3!Ѝ��40�R��Ő�2U�`����p��X�b�" �XX�\�"�r����b%��aERW.QZ�(�	��hg,����G�"�YTJ'*�2��Q1bò$�PW2���"p��Dr�
U#D��hIЊ ��\�(I�� �I*�wiD�r�ZHr����dZ	U�k.�3 �E%h�۲+�NE�ېk��ZHs6�r\C["�w�X�ye	UW&'(�T��ar�Ay�@��d�B@�f�E�"�B�f)A;�ʨ�bak.�㜣ٲ�+Yl����1P��D�E4Ԧ�I9�'t�$\�3GSւ�jҳ9d@s���)@�evY�(��h~ �E!D/�g'��~���m�&��q���ۃ��)��IC��4��%w��P?�]d�щa��'[GJ��*`]-�q�D}��ikV-i[�F��\B�tr�|�s!����34:����)[��i�j[fy��Q���̷����B{����?y��ߛFW���>�3z��a��}=F��^������^Cx�kYׯv���ݞec=��yVG����֟���AJ��إ�5GV�Yqp9r�V���Heg��M�7�L��ngLꨶ�/����TB�z�f�M�ߗw�j/]7c�6�Fwk�w����]o6�'}3��X��ھ!@=9��_�P��T���X�3t����v{Cz�8�g�y�)�2��D�������j�-f��)${j�u�Q�㫥��Ӷݶg%��,�Ǫ�rz�P=��4�y�_v��4���jS���w��ۻU7R��uN�c�p�Ou����=������z�)�|i�䟛`�=�d�#�u�����r}m����K�.U��iu<��X�ɩs��ɮ��9�����D�"K��	��kp���o:�f����8.;�ܗu���к���9ܠ�0��LԖ��ӍA+wA��F1Wh��1�y�`x������֋�3�W�}_Tk88���zk��!��5�v�F�C��eI캭>�ݧ��=���H=����Hຎ�^��8��:�o�ܡ�"v����0u�6��%�^՞��t���pÂ��[��W�c:��F��r�yI�)�dQOKE3�o�hTY�B�p^B��v)���}�Qyв�ށn�A��WC}��N"�x�{_mZ������B�1[!:7�2��� ��򲳶�S����8���kRC�9;�K�=�Rz��ǋ�y�0ZX�>=k<����M�ױ�o����\9E�߱��T�Y�n��8-�M�/��/g9c��o�wND6gu��:��*Z���N��ՉCG�1���5{�k�e�ޝ���+Gb͕��v�b���pyy�6gFͣU��8i���-�0�.+�,Um��޶ގ�x�U������qL�3�d.�䘜�f��u;m���\�>Sl����}gb{�;���QK� 2�˵j��$�tkj��p�[L��N�w;�$uP���]��\s�nNÊ˸D<�C�שL��R����^ ��)��}ۉq� �Y� ����n��M����,�!z#ﾈ���Kq�������@�-i����������
b��z���y/�¸p�{�E�=�ŎW�u��e�}���cb��m:�m���㏋���Ҋ ���[P���W�3��{D��Q�~i�#��ɝ���M�3g�_5�N�jW:_Z�W9��:���>wQ��f�"����3׷ˆ��N *�m|���:1wNJ��qm�B=��[Sώ��̬C\�&�\:�V1c�Wc�/��9�w4�!��@�^0���}������'�� ༉[�����'���C�=�-_�3W8Ynu��ovݼ�׊�в���o{�*]g�V"�x2�]�Y^��g�龫�ٽK!��<蕚�9%���T��~S���]��9P?h�}w�����7oE��O��c���nR�%��+�y�̕��ޙ���_�!R`�0z��Xt�͹�Ky��s��<�|���و����*x,PA띎#�K�fw�p���4�C-��&���t_NF�����A� D����0V�<�*=��Wn�	u�����r������Nz�������}�}Awt���5��5Gп�����"\x�UW�O��c��ۋ�Ԭ��%�<��գR��Yܜ�EjD-(޶wq�Ѻ]Z5\$9En��fT��
��}G�����{΅&���r��ܼ��^�3ϴE���!�X���r�}Ĭ7~l�oP���(��qժE��\�!U�;̫����n3�#�u,���<���p�HY�3��r�|cTII���O_M��1�'-��囖�Z��b�W	u,9Ѣ���������"��D�J�iݚװj�]˯4e������<�6U������g	Bt�Gw��xU��¶��YT��ћw��ߟN��ӷ�yF˼_r��该��9��i�jR�ֻQ�r]�뉸���L��=`ۻUp�K��|������q�LI
��<�?����<r��"�=�0�ظum#������d�͇�o���vdv("��֫*(��۲�\�!
L�{#�sdb��.�:d�%R8@��U�p32:죧�Z�sj��u��� �M�پѯ���%�U�8���C��`��tٗ%l���kT���Ty&3�{�l�Ic�7k:��C�k�-Z�/�>��������.N�":;�DF�rURx���u�xy�YL��8���Z۞Vo%�h�%r�=/���ŵ[��*o�b��ڔ^r*Г��O�8�t�z��뗽>;c��Yc�GK��Nŉ�Ԡ��>�K����{��8�q�l�د�� ���}ݻq���T�z�w�CT�T��f
W����3�U8��%��@5�X=��^�8gno`�;y�;��]����6��f��~���4󽺕{���������$c�l�+i�eh�:�}�����Z۷�W�L�9Kt!p���n�={���P�p�*7iC��Q�ŗ˖T�Ϩ��kҌV�n�/�ں	����Y�l�ȅ[�B͊��(]a�F(�v���c�Jk7�$7���V�j��~�<�π�O�
�E�K��N��]OE�GS��ܽ��kL]��8�6z4F��Q���Z�3��VAW3Fozw�g_(z�r�.�V�֜ɻ����l؛��ڱġAa�eY���0�p�t�Q]��+M6z��q�(��f�F5)κP��»:�lvR�F�`�</}�}�T�\.m%�B�M���Xg!4�����6�]�QD�o��)b>b���{��G�l9�\�U�w�_kK��{l�8n��#e\b����_u���w���h�_8U$�����}v���ɜw�q��Y
����,�&�����zpͳ�>������LG"~��'�-kf&���·n�F+��_&e�UJ�J���|�4GB�1q-��l���lZ�}��U�b�:vu���T����i��{	ӭ����+��__��T]���[8�Oq�$��'�-�M
e9J\k�[��V��:��@��M�Nc������ds���"��;Q�6ʆ.p^![>��k |ǵ}�+�ŗ Kշ;z�o�ٍnt�+j#j��]m�\F+`�to�q���>�+>�X�v��A��V=�0���{;ju�mq�w8/>f�p�����i�hK�>`���'Y��a��p�Z�����L���V���v/.��u)%tb�iq�Yހ�2�sv���Ϥ}G�9�A����\��ʆ��k��w�ȩe��J8k�y���k���¢���ԭ���U�7=�(w�"#��t��Z/�}��za�T� M_Օ��';�-��|<�>Lb��wدJ����^~1��O+�u�y��G��ϊ::��)�ƭk˦���c~�e��	��\s��ٳϴN�}%x���tƦk�ƫ}s#mL~��V�x��[K���:u[}��z�z;)�p�k�6d�k}m�EN��}D)�]{٢L���r�����@y��JX9���[)�%�h���p�Ep/r(=��}c�͵O�Ӱy�ϳ�J�2jH��lc�%<��n�&F˸��;�J(����[q�	�U�;�U��D�r��v��k��NS��;n����q��X#�l�s���t���Kr�d`(_t������a�w�fm��wn��U��Y1д��Mi���E�+�R���m���#x�����r��0��_�S����t˦�z\ޥ7o�+�w��V&* 
��E�3eH;w�c������G�} �]~��ͻ�7�7��h���L)�.)>꽸�fl�|Ra�9��J�ӷ:��v� �샆�]WR^�A%�����;�x��v��vҸ��t�QY"�gu���^�>��>��_3�������u���etB���9��Qy��5.�Q��N�����z?Pw�� fU��v��v��쌃e9���
Տf�(�Nؔ�G>�)���}cu��ΎIk��΋误<����Q��*��k�}o'�ܶP^�X����a+�s�Ng��.�A.�yE}��skg���<�T�A��d����t?�o��y�D��������n�Ϋ�^��&t�\�U0�Y��#�o��Z�C�7��O+�u{�F��k����O�t|�
������3o�+iy�~}X'kƱ�j�2�v,�F]=J�M;��h��/nI���8t�2�g��z���gN\s�����w���ޭ6��.HR���g��u��X&��J9_�_ڠbH$Ӵ�aș�p��E�ԥS=ZT������}�ǩ���|O�,γ�J�zV�<�R��x�`��d[| 
�.���!�G�n��)kL�ۧ~�YGz^a��
M��i
Y��k��y�Iˬڏ!:i�R�#�	�n;zi�u,������J�fu����I�&��y5L���L���2�8��=� n��$ޡO:�U�E�r����>�X������Y��qM=A�yF�.�}<z��>��[�zkW�)�:Z<�v��n����Ӯ����v�|Fϗ}:#>�X2��]˓��+�NJ8��*��'8�s5��Jgq&f����v��,���p�Q13a͂�t���qQ8ȹ�r��������ob�պJ�W�I��6�goaLC;��״�����U�Ws2�㖈ݓ/�m=慌'[YX!��˾�QsED���n��US×��Ç/[�۞��W^������W��n+汋r�>��=��Er>�^��j׸�qM��}Z�W�\1p��7ζ�ب}�5r�gn�q�h�'�/wK���zz���x�<P����������lƘ绘��L� >���3�{zz�^z�����{��5���W�y�z��۩�����{��pS�N�9K�u2.���G�F�c`+ވ�h�|W$�D��� %�W�����~����{cȳF��Y�&�Y��MU�7<4%ӻ>�f�A�7���~ic�5\�	���v���a��ȞR�^�/� Ыrj=ў�x@ʅ�����;�J�N<���&�Í������*Ö���/^N�2�Wi���gugz	2���<�.R�����S���o�EƮWPɋ�E�S��Ͻݪ=~�W�vO]�~Y��>U�lR܊��v��[�wk�+�LQ�$�էګz߽:��:�>��+���rVM� �Ŧ��Z�RH�v�޼i�-a��4����6Sje�lt���TuOG^��R������.�]u�K��K7�>������5��0l>��7�u������c'�����C�~��3�u�s�V�Q�7u�A��v��	�b��R5�k�2�sϖo6�����*�&�W���ܓ}Ŝ���y.Xy~���+�@�Eķכ*���/T�z�VF�%�����9�+����:�
���T��/��ѫ���@���xE2�����%gVlɌQ�@�v�^R��L����C限��' K����1^���f>�:G�e��l�fV�C7�r?b��us�m=c�v��Qަ8��ܱ.*������sf��`Ql��]E:�ּZ�\7"l�V2V���^f���yQ���j�b)r�Vhb9R�W�'�:�h[���H��L��0��Gj�J<.h}���5B�@��+t6R��n���쫑��N���j�U��u�l�­�\�੬�L�m�3je/������G�Ԇ�۬=J���d���XTvve�¥�z���&�n^�@Ouok�����bqʽx���i�� N5,������X�L�d+��R�em�:iܥ�ӦQ�Y�n�[��ø�����e���F��l^���wQ�D�{n�N�G3��\���+2F�XњmU��SV�ڽ��s�u�(���tSW��l!G����Kŗk]��j�B�o��7�.��י���Wx5����J+�[Al�d��܆8�ʼ�1�c��:�b��Gxܹ�höI�t���A��Kv+z㹕#�x����ܛ9�����h//3a}���,>�a�ک�Jl�.�]��'A��ou���;6��k��+z��3u��v��0)�Gg&oR蓑h7*ݝ34gP嫲Xp�E��k�\���aս'Hg���s#�v>g&��3��Ȧ����HTk!!�靮�7{skbS������ȁ6��l�+%[wםS]@�6����[N��u���5NV��:��-�ޜ�iق��l�9f���,�|�V���L�V���V�L|�~5|�"qs�/*��ݙ���̂���r}8>툪��]�-�;���D�^v<,�t=�gwW$s*��Y�q/�w��{�6V��(��Vd�R��VvWNU�	v�w�t�����q�2�9r�E�P�6�wiV�]���TD�jí4)mnswa�9*٣���)��X�|_iŹzF�ņ'E��H/8ӹ�SH���l�=����X�Mjܟe��Q��� ����s3Mi�WH���t��\��E�lE����Qj�ax(��k��(���B�y?b���nQv^U��5��R�<M�j��r		�,���4���E|D�za�WGfb6!��@�ݘ0�B��R�_��N�o.��X�̏�gѫ�b����^F�)�r�XڀJ�0gS%��}xknk��
��_%�P�s*�e�	��*�.�(�]%��t.nl��bJ�.�F{�܈i���v�Z�mV�N�=6�����T����ZN�34R�D�y6K;C×u�;�JXI�d�J�(�O+]t��3h�&�	ݕ��{��8N�-�XR�t�wVFz�V�3y�q\�ff8)�{��*3��
mU�U������:Q�n��v@�d��AE( ˽���K�P/���/�Q�=�"���MT�Rl�Rӆ��P�*)!L-H���JTsS�l*)ft-"�H�YBh�Q�Nj\���M4�س$�wu���;����*��1�)H�s&\�u��V�J�A(�
���5�;��N�ܒ���AK$���u�E.�$���5MVvRI�SbqUfP�"F�9^��e�ۇ".zУ�RB̭!
f���fE*�9���a��"��¼�	H�VR��$�k��:J��XPR��\���jB�����9)y�d��%%�H���G��ng������u�'*�&r2��Br��Dj��d��i$f��vN��*�s	�,��S�(t�.H��(�/5�T�0���G-up:�jM}:Ktn���4H�Ď��W�d��_R�7K��uCA�0��u%�5&u+�"a~�#�cu�����v��VB�[��W�c�_�(뀢��m҆h.G�_s���p��k��
*P���
ۈ};�X=L,�[��d�Ւ��P��w(�y�}�Nv|�w)?W�vx>�Ի�GA�����(-ju��R��OBV���3<[{K��;ʢθ=�Rz��x>A��w�c����W�N��#~�&G^Cxf)I�k�%��~��YXu���̽�e5�~�;�^	�S��>��wK{9�<�
���ۊP��cs��gӱ�=���=�PW�gZ�w�T�<�y&T{��A����B��aT)S�;a�tyr��G�����*R�q3���j�t�\����~��R����r���Q@�W:����дy����k��y�#Fך�����k����U������А��nft�f�ٺ&ٲ��S$�s�;��de�zST��y7�{��$�g���J��"���U{Sn:M`R*����M˂A������ȡ��i�˽	��L �*f�Gǂm��u8=�Cݻ���pv�)��Tu�e��eqai�9S�]���坮}��w^���Pvi}���w�W�'Vn��Ɏ��T���}����M"iqR;����a.���P����O��Οlp���̧K�]9���I�EHA�eT�ꅪ��U�ʙQW/�x-uշ�ܻ=�7���C�;�����FG�k�}x��k����R�{ڱR�Y'W?G�9W(V����q[�7ދ��"Q�����%���c��P=2x�!�H��(_�dkh6��8���ڬۭ�;=b\�,�M�v]���v7�T|?{#�s��*�����Dv��s1׫�}�]^��0fڐ����TT�w�#���ԅ����X�uG�QΝ�O<؁K}��5��f8�~����O�&g ~��3u֣�|�xo��Ȭ�����	˜E_�+�x��{�ݥN½�8|���#ʀ'�kt/�2=c �E�o.cK�N��ή�zn;�U������/�+]!�h�=^�!�Ig�N,v�v��4l�9^����ތ=�͎ִ�נ��#7��k�M�]I�~���̒��/���ļ�G���mh�����ދ/�R�� �3>��9�*���n��m�s^�=�m�d��9Pl5�{��.�6 ���Ϳ:\�v�v�G����o�4������iU��Φ��A���l�ALF���<�G��l�9����M���qo]D����BŐiVi�WVe��lo(��ʚa�C�z6�>lj�;zb��\���aH�>=ܗe�F�����!�w�HX���������y�!�������߼�gܨ���Ͻ��!0-Vu�c�fn�lb^4��07��	
��^Y�F�] =���G�9ӌ�|�v��J����U�Oj�N�ky���K7}���r�k�``Ǫ�AرZ�K�Lq�����f��M��qt|4V8��*o�=W��>��A��=���t��hy{m���2c�<��uZ�2�֘��Oʌ��*kƞB���|�}��T�T�x���~y�-_��<r�Q���qp0=�1]~�R6
�d��w|�(!��mE�ո{I���n�f��,��H�)L�![�]�,����3��Y9��Ɩ��9�������N�U�	�%���%��ul��.{}�X�t�4"� �ܼ3@�쨴	�~^�O,e�9��k�^G)��E��q���7ة�q-#�X��7鑥�B���5�3~;=���k�W���
Y���uʫ}�2�`4�¼}u��O+s1S��d���_L������bc��_���]�(61j�8(<6�~=�^յ��1a����g�����]ו�{�y^���� 7�Jq�w�}�o�Kc�oRarΝ=u���L˧}�0v��^�z�.��p�m���wܮ���A���5n=��-��loe���/(vd\jΰ�}�P��
GZ���?C�|L�����/ �z�����N�,�����?|�}��G����:¯��~�WPt�P�=�$H>���Ƈ�	�����>��>��pf����?q��^�i��c��Pb�%���T��b�(�qDsݼ�yu�c5���A���;�3�7|&����%i����2���E��r��w?�����y63��Z���hFR�Q����t^W�}>{�n��tp���r�7
����żLTl�q����qٍ���2�8���.4�1���ohrt@2\z쑑�~�v�p��qڇ�9��`%����Wg�^J%�*�^�=��kC�ҥ��5���״:w��u[:c���۪�QLKU�tA�8��k{��nd���M�l��s��T�=�t�il�3�]� �t�Qe�����Ag�l�|dy�N���6�ژ2���ko"��W�������B=����l�%˸6b�s����^a���z�l�3�jg|d���T7�B٠�ϭ��P�/���g����d�&�b���K�|z�9��٩�/���עf���HQ��ș���F�[�wnp�����72�����oQ��z��� ��SN���dS��:�b����q����e�o+�L�e����+�����Z:���Z�C�r�t���G��Du���4���G��LO�������@#s�iL��7U,uB��8�0��>���Bw����Az��dS��W��������֤i���304v����Y�M�|�q|x��o3�r��x�]i�/����H��ҦUO$O�K�؏L��v��3}�Pj�IСxz�d����;���K�[S����Y/	�3�O\�9L�戮rju";m�Ch9�"�ѧ�9�n���r�=�3�m�K�n�E�?`cze��q�zh�C�NMN�Cެy���B�
v.��k�A�5b�vvʨ��<�Ն+�Ĥ*�A��t�1����Q����wq���5V̧���R�$~�;�S;)k���}ە���ߓ��~c�]Vy��j���Sm��>6k�o9b>Ź��|�7#3�;5T��W)_-ۯ�Y�3�L7�.=~�}���j�&4gK���K���/Au]7ޏvl�}����P���3j/n�Ȱ�\L���/1{�9>+PFw��ۋ�1���}�y�s,{5�Xʇ��8-�G��,[<��>��[=���T燛��P��1Z/�4C�6n��rw����j��4�����ma���ᆳ��O�ܪOnݽjxp��ᶱd��
��(G���}y�G�"u����Q�:�����:/[y$��6�	O����֪��Cx��y��>KE@��������;}�[��ZI��
f�� _ܯ���O����N�&|V�p�� 5��2`�Isn�]l���ڪY��;h��^�ơd�v�=(=�u@��O��ޛ�SA��L7֧
2}૯����+��>Q���*��2�?\��7����]F����=��%�x���n#δ�]#�;)�ͺ�C�.C��`��M�s�;��dg�U�LX
_AW�����m�Jb{$gl�}��TȤ\^�c/�wL<��@鯚�3p� ��� �fT7��Lf�Q"�9��^�����;��8����V'O�/4�ʶõ�� �0o�{�6ݑ�]ǇC�r]��B+ԯ�G��t�&���N4�(zy#ơ�H�Hzc����~�{����i�^�	�sN��ך��K�x�tϙ5�7Q��\Xb�C������5A>V�E������4irׇ��ddxz|������X�Tx�jWS���y�5Z���]פ�d�ӑ2�(ǊB���'2��'�nqu]�w�o�_{ ׷���x�͎�������.�')������\Y�L.�2�6�+*��U��N' �-��i�7y�V�V91�gV.�*nWEO%Y|Nu�|E��-�a��ʲ�.�W�g7ɧ���vZS�a��u��=�חurB蕃7˩}]�XS�]�fpo�W'��M�{꬧Y#ʷꪹ�OV�?Xdz�ȿ�.�y�ڟu��x~.l-��N�=<~�j���@�t���f����	���]#�G���-�Ba�}��Y���5�]I�IS���\�)�(����~�[�������'������J������;	l��P���>]�O��D隍}����F�f��s|��`���X���Nus����Ŋ���Nbݯ>#�w�/B�P�r�g�����~�倅�N���6l�����kxB��*6�t>���R;Dv��	�yF��u����V�o�.^���T_q�B+��q5���-�e1��s�w�T��m��0}V�Ŋ�3�%1�A��������ү*�K��������˃᾵~��/��Vh{}�� �S�1ÞA۪�Q�w�L[�>QYN�����q����5'n�
/e�"��r�r�T<��W���<j/�z���0d�9ˆ�uD*#�[)o-�̨�1u{K�+���;��P#���d��fxG�#��ᑮ*e5q&�
�!�;]/�JF#��W/=�$Dn�5�6����í��
�����% ��Zu����NIa�|L؟/?~��d�`���?n+ON��w+�z�d���>�z��5t����d�\�˖�-��Ʉ�����20_Tﾈ��xEs������萘����VD��dmd���]}9�~���x��}�\=v�.�B��7�+�[Y���v�B�^l��,�4#؀Pn{�c�-�m�xW�<���9��p˭������E��n��@>T�D��OqD�;Y��b��t��@������LԘk�Wzǽ^�����?��X��s�`�����TN�{f�!���{1$�U�hdof�G��,���*68����K�JJ�y<ɓ��=���(z�������[?�St<�;#�=N�/c]c}��T�����o.r����_�5�t�5��Ƈ�	��}h������uQK��<��V�WA:[��7���O�ˈ�c�<�/���C�j�k�3߲���knn�X:�紝��'���q��зMw8�(��>=~zln��m��ξn�WxŞ˞œʗ,Ƥ�ȝ�����y���C��[J=�;�� �>���w�:�%~�Ѥ|ʯnr��>�z=�����G����p���XN���j��U�/%�H����įYo��zR�)bɩ�R7c:$�G��J̐�;Z�{q��C���A���d��nM�s�mh;���;�s�j������%C�2L2��Mn��R��m��v�@�ū��ɱU�!l)+��Vs���Ot򽉀E����/��"y��W��K���ED�Ѽn9Rc��u�?5rp__�����2�\)�هIH�65>g��β�]ޓ��/q5�߅NC~��mR���+�j��<o�|�=�hu51�|y�\��\�:�m`����#w�2o���E3^�QP��=���#ˁ���,�ƧL�K٠l��?�%����i\����dd]R���/%1��&ϝ�8�V<;>�Z�E}���r1�t�(��R�"�}nDt�G@E� Y�>�3���UK;>�=/���qLgT�ui����w�۸i�h��h�4��6�s|@��F�J��v'i�VHR�g۔e��/����1�����GI�����-�Rz=��P|?�Tʆ�+j��E��/D���;�>��1�W��W^��P׼�F��ǉ�Ohk�s���\��ĵ����M����]��E><�z$?����\\�*=�G-�RaFg:<o�\q��D}iɞ��fx��6�e�������Ex#���W�笪��Q�1Q�HQY�9�����5ǣϾ�y��?	ҋ\��P��Q̥��g���CW�����ĳX^7��X> �6WV_XX*�>U�5�(���s;s����|�ɔ����XwM�whW'�5��K{�r:ǝ�T</Tp�#R�>�j`��u)vMF
kI�3�Ԇ�[�H�l;��U}P5�}W�������ZE�����
>1f=���~8�p�fϯg��b���U�5�{�8�6j_ْ�TCquP�zf_vg�v��q�n��Ba��Qx_�727 ����#۾|[� 3M�I���<�Q���w�I�[H�㓁MLّ̛.ܙ����bc=�wr��I��w�\�;�<=��Xʈx����|}q2ű��B|�Uf�)�\�f{3s�O����>?(>s�0:'z���I�g��X��{t���.��z�i��>�b=}t��w��b���H�U,"*|�����_{"�SN�;��y1z�'��_,�q�]�دf蝷:^\�N�9Q|i�u�jf��B�z��hڏ5ADE�._w���������o�(:�B�/<7����ִ;�ǆG�L ��W&㫞A��Ⱥ�Jcc*����'ѽ�/GP�<Z�W>�{��gF��#_S��n9��#]���jx�:�ǏY�t�.�i���y7s��E��价�=�7�p�&�=�vE�:UǮ!��,��H����b�ﾎ�g�����&����^J@�~����9Z�<�����|�u����R�:�D6�Y�����uH�F&�xէ}{�اr�-�;�&{����2�301sU<oJ�m-v�-���c�F�e�,W,��xwf�NRL;֜�����йn�-��;��L�(�iP��٨v���S/ud��o�����k���^[8>���N{�|�ea"�f�ǫ&�5�a��@�[�uԝzs��m���Ft��wC�y��Q��N�,iJ�:�b�\�_u /��� �s#�������5�&D�S�j���F�yjP��趧�[�u�D�hNO�M�N�ﺢ�������z�h�*d�j	�q������X�)Ӿۛ݁TU��+5e��}��0��/'WX���;xr�A�]9�.AJCjoL�)���k8vm�Aܖ��o'u�R�M���$�ˋ�=��-TKm|�`�d5��%���ی.Ov�$�7���h�k{�C��8��V�C�-� x��n�+��J=��K�aaYY�f)�0+'s�Z'����w�Y���i���u�
��d�ީ�e���.1n~�f���+Z ���)���<�N.�!ע��9?�M�*<�
����nQ��M��\+�83�Tۅp���ZfF2���ݘ�-��I��`����[Ϧ��qnQ�%:ڕ���q�[].�r��D5��q]����|-ɺ��0Q���G��%�e(l�o�:r(��ӻk�o��^$2^a�>ڹO�JM'�i���މ��]mVY���%�ڐ��:�h9�(�V�6vHm5�����I���@��rm1�pJ�%�sD��kswLec	`̏`�a���(���׸���g��Qb��ܣ(�P����c��'e6 N�_7+��w_:�#	v8�ٛ�2��]�ʝꑈÖ��g)�3@h�ԗ{�Y��d��lwh6+dׯSPQ�ɐ'N;��ݚ)=�u����L�;/%F��nS�
\p�Ҹ2�,����\�6��ٔj��+Aǐ|�L��0M�� ���+�J�wʷ)��F��uJ�E�I���
��&̰�q湼�8)a�Js���;��S6��x3哚��b���4fS &k�<��Xsda�C��2G-������#"�8�[�B�sx1�k�C6��ss��QP�k,It�>�	�����RZ��T��6���Idڱ�w=�u�_-<�T���q4�O+0l����'�^����N�1�#�4Nm�Rnv���ف>$��fwW����Dq������ q��I�y��_�tM� �}�.�\N���ܤޜka�7Jg7�-Q�c�J��x���X����q�p��{r���I�y8Ց�����I�MvE��r�ɸR�z__ ݵzoݘomj��i����F�@�3��0��S#T	��N�;/�����B��7x�DUI��(��V�uJ)E(�H�1iũ���«�dSBH�$S����dB�%t�.�VR��U-fe�r*9C�HF%J,��q!�i˅��х�$D�8[P�bē�:�C�"u
���! ��ad�ʣX�f(D�	�$�2ҘZ�jʦҝbIʋ��:g(�Ms��9HJK�("=���ʤ��)���(]c��PQE�hP\�#�DeHh�wp�\u*�W2KR��$'�`D\)Ȧ)*<x���.��ܕ�̵�d���'V���OWs�D�\*̓W<�U$]����R��!���2���"�z."��C�UM=ńL��Jr=�N��)�P�G�wU�M~����B�QY�2�o�6�F���LrtM�[�ح6f�zP�t��y=�{����3���;W1n��1	����&��z�s�O�(;ʊ����VF���_p�{^�ۯp>���{*�B�y#ƢD��P�>��Lk�f����	���6�� gj���k
���x�6����=��u
0uހ�֯�͍�=
����#9�F��^����E��.x�]J^����L���,UT��(�r�v��$���]�"x�~�7���ZEU�2�O��ܕ$�/�%�X-x��Z��{���\vV�n�=_=���ϧ��{73s���H�dz�D�ݩ��:�b_g��|��~ļo���_4��Hz��f����	���������ǜ����&��N&y�g ����A��Y¼Doz(��]�mo��˞������P������ڎ�O���BS�~�OEI�>�#�'��vC��L�K���W����4]}�^�;z?���[�{��}N}�JB�g�B�5��?_��A�3Z�M��:�TN���\�y���dF�Kɭbx�%�����v��mlz�	귑v�|n���]G��O0�o�K��>w�����L�(C���jx������ݛtk�ӷ���c~�ֻ�\��3V?\t
~�K���|�oM��\K�����]�d���޹�/������|�i�t( *wj�s(w��\9^�àƯ%��wIlɤ�Q�����ݡr�8IZb���ʅj�������W�߻����ʕ��`3�wZ�z����T��Ɓ�ﱎ�������G-N�����{�i����Z��skF�c��=p�9 7T�Lp�v.�UG���1�ڸi���$-]�$Z���L,�*�u��O2�;a��{����=�p�!�j����[�����4o�tN�λ3;z��R���z�η�)��k#&ϼ�p?5@�g��}P�S0�0�d�Yc�Lؿy�W�f�\`J�8����5 ����.����[���+�:$�W�/7]��o�w�̸O�9G[��Y@h����3@��Q��=��'}����Q"_[>���߸�!����]|��Nג=5��_4��#b&������T>�L-N_GTK���d���Q��f��8� ��0j'���;2{e��C�G�K�š0�q��^���JA��~}є^�Lb�%%}�;�ɨ�hw���C�h��Xrjv�gH22������f�>X�-P�g�_�}}�f�x��7�Q�)0���95����Hz� ({jd��-�U��phfՓ�P=�Qi�kw1�Yi��i*8;9�{jH;V@>�ǿ1�^���`D�ά�t��Wg~i����#�䭾�i����~����n�S��0�/Yw,^m�c��1Œ9'Kź�s�1�ۜ/�\���z�9Ӻ�G`����;+yE�������H�9~�����&����W�F��]R�u���	1xnt+��:%x�+�ok��w�������e��sM�(��>����y�n������κ����>�H�e^�����qw�d�g��6W�;�
���H�a�35����%2��ԋܚ�þ{d9���m���}����z�'/ya82�^�fyB��^4�@zo��0��s\+䭈��w\���I���L:�����r�=��AN�M��;�'>�rk��s��X넩myr�r5����FiŨ˙�Q��3mR���ҽ����<o�k�!Ƴ;S���������\l56�RS��⌍�󨠢���j;�˜��}P��W���)��G���R����7�5� ~��nf�sw�dg�T�{r�S�����xuRՂ���R\�u��e�.VT<%�� gt9Q�x�{��L��7U,uD-pJ�:�Wަ��u�Ob������w�����q���#�%�y������թQ�P�癚����ɽܥ��n�6��B�su��#����0t���7�ϴ[+�HNڧ�y~�U��S��A҄_{���@���^��\'N�f%�E��z\�{/}<��G)Ĕ�e5��!~�O�����kftzءI;�)W_d����ZtgR����fp��J�+�Kw�=F����O��>�^�u#����D�}H���õEZZ�K}�Z���Ǝ4���EzF���	���]��e�<n:g̞�6��e�@�+�-Z毬���簽�ݣ7�G;xH7Ӗi�r�Q�#�����3�7�.;�У�@����aϮE;���ʗë3�S����d�(�V*}�������<Ն+q)
"��s5�,h9�69���վݵ}��(	���]ֈ{pL������B=������yR�X�x�Ş�۫�w���5]ٻ9LY�بd�޹C+\]E=���|�l٧9��60L{�+#�~�1_��a�߯�qy�x����@c/&XY�<�Q���v�d�����:Tt����ix��;���y��q/�/��a:\C9b�n�����y���Lf�.�~8-�eN�H���1&�#,ʟt�́}���GB�f�x	�ʂ��0*'z���T��{�]�_��<#��������g�\�O�����!V��}f��R��W>X^D�}���Y��iֻ��yx�{��T���C>tshu w%p�3WJH�4q���,ʝ��ʅ���O:�=y;dY����I����U����}��h��~#�j�<�ga�k��6cy,��Λ+Mmޚ7z���V�&���B��M�Na����SFnU�:����n�q�YeB�_K���s#�[�������㫍c#�~�4 b�L��n����}˄��Z�u���܃�Qr���מ(7}-DW���xd{��\8���y~�L���)�K�����c�����\���Dj��������˗u���g��}|��MO ��T�i��W���{��R5��p�=��e�ɸ����=��x$���>���z� 79������_���ɣnB���R�O�6j+"G.��FK�+�1�{���t�&���NT:�e
�H�î� A���k���M�^��W��� �B��k��v�ȎQ�`���X�7�?z�bj�3�2�C�Jyo^8O�r�$��;xH7��H_M�aUS�.�؈��jB�ְ�Qy������*�J�3u'�?�j<}}pORrb����$ދ��h5�2��:�.�}���#Φ�������{�ù/��4��_"ދP5�3Q=4ٸ��1�������z����N+~P�6s�wS�.<�FW�/��I�r�s�<�M�z�&C����qw����_��g� � ��^I���12u�7�����<9���^įp41�)�f�:;l���=��V���B�).Q�:��ϗ}m��]�(��f�gs/�<��B:��ud���l5����>�h�G�ԩ��p�I�YdS��^�Z�"��A�����x{�A�!����#�#;�E�j�7ޏ~˞�~�������=#ާ+�R�(�(�H�;�틢GNZ�ύzf��vC��L�K��U~��Y��;��4��'���#����l����
��1i�W+ƾ],���倅�:�W�:��_���
�_�۵Y�x��t����>��� �h�Tn��yF��g�� nG���&��U��#/M?V���h��Y���w��8�v9Ͻ�9R�=��d;�c>�[�;+PȰ�S�o��@����]�����ۗ!8�@LE�f��᾵o����S��vh?e9 7T�L�q�w���V?��E���QU����
c�A���k��NC.�õ��{�z��o
2ϯ�z���n�\:Z����flk�2ӑ� �Q�uIz�#Jy�2l��I�uoj�!��a�C�[4���7�N�;��6�G��3�0{�s���s6�|�.����}'[�p���9�>˹��zvi8�/�u^�U��G�E���B=�n{��e}hq^x��/4*�z��Wݚl$/&�)ur;\b�֪���]��ג}IrW��ԆI�;l1��&{�M�ޓLc�/�d#�ב޳�J��ܸx�˅M$GMnWUv�J+2,졝ڧS�t�u�h@H{ݕ�
��Ӈ���چ�(Z�x��3���,��(�S���m`�k&q�"�/^^l�{f�%�����p�L�����B���u7[O�D�~≀��]f��Ѹ�7m�W��|���x0]��s�`��s1�H�͹�_�)ՙ���<yR������=u�2}e��/��IQ�<ɓ[���r�d�/��ÓQ�%���ö�5�7�h��(vouo�/���`��p;��и�ׯ~mQ�	��,kR/�������w���s���G�ӱ�> ���t0]S��.�P᱒�Qx�t��_M38����%z�� 6�wu�X�=���'6v<��_���/t��,ӯ�.?��ۜT���4���[�U���5)]��%�����
�;yU��T��[%���PҾ�ܨU
���=: q�<��}sN�e��<�/��Ǚ��<;����4;~N���V�1귑yn�q���Ǔ�R�����>Է�$����S;λ�r��Lk��I���9Y��
w�i��u[:1�T ���������\�t-��of)d��Q+��{�	�\̊�湛��p{��4ܿ㫈^�:*ЃBm~�����Og0�+��o��c�Q���卽�,_�;]��5(�Dq�p�c���H,*Ԕ����O8�8�nm��볜���Hg�јm�n�ot[��tke�$J-�8m�Q���$Ȳ�)��������c��ow7xZdj�&l�QɽV~ ���x=t�_�����5A�]�
���2n5��Y�y9s��>�yk�^�Y)���[��{+vyn{0C3��нL�V�o�sv.��@)^��S�����(����k���ݛ�h���暇�|���7��r������Q
gGa��c����x�]v��ĥ��}�*��yؒ�E�Dz��WP�E�_HznH�;��35;n<1^ϫ������C,������[2�>s���6�FW��S*�y"xS�E���5�O���YoϔeKW+�EW����G5Yf��߸d)����'�́﹪e
�Iɻ��g�R�ZY�Q/7��3��*�Ɲ��Q��. �	h�P��~������w7��'���{L���VŐ/�nK���L��<��]�����q)
��s3<>�|Dc��n�{�vq�
ߍB����멒�Z!��L���N/x�#�/.1p�^T��z'�^���	[R��go��|qq؆���T��s�=�ѹ�yY��1�)W�7Vl�R�����vPt^��{�Q�Ƣ��y�z�V��΅�	��SWR�d�B� q�m�ܤ�JծUУ�"��r}�Z��ύ(D���ĳ ф��;7y�D��N�+��U��Lz���P����\e*����g��ȫAـI4q��#���Ge
jv@Ul�nEj�I*yC��}<�~I��x{��7��V3���|�L��̝9�N,�	��nW�� �"��#� �=u��ϐ���6�9�=�.�~8-�eN�pI�xi7g�o��+�÷7�u���;f�X}�}�gys;ʓ�D?f�Kg;��[�D��5�i���ԇ���^���
�.h�@�n����|�������ȪTӫ��j���^E�_2��>3�|��?x�!��`��5���~�'֔��� ;��8v~V-L�+U>Gл������������U��kC���S <��É��y�=���Ӳ�޵.4���*/���.5���ɽ�l��Ixn<�1�����������5<ÝPT틚��S�{�������h<7��S�W�pz����<����=N�q���t��e.�mo�R��;�65��6`@�dĸ{&��n�[Y�*y?��΢r��S(��U=�S�K�{�UqE�lH��T@=�B���`>;�_���`�[/(�m��I8���4�-�T�уδ㒯� ����	�a����g!�/ T3:��G�s]�hn6�V�M`1���Ziv`YJ��å��t��c��3۩]�5�r�Uݽ܅�/*b��.���ә�j0/�F��>V��ж�+h�]��rfH��;Nw,��P*u
�\��Q��ā�>/T����.����j#�3䇦���f�`?b3���#J���+�yo�A�����)��������$ދ�}�J/|e�:�-qމK�m����k�/�%��s�*���՜�3_wS�d[�j��nf���j�=�5��B��VDo���e���-�'XmϼW�T�sfl�t���_4̇�9V4fyY�SG���oR���x��eD�Fe�	��n�����y�
��oz/��}w���=�g�f}����;��������P�BW z�C���::k�@�i��o�!�n�����=��l:����r���W��\�
�^��L���Nl�����w�@�5�.U�Y4�X;_yp�
1�T��*yu�����r��/.��{^��[+����3����3��$dz��]�)��r7�M����~��덁�3��yY\�\͐�U����|G����*V�{m�x�)�4�uG��f���e�o�59>��ZZ��1+���N}�U���?Cw�~�V��Y�9�f��S�uJf���Ըq�X�u;��,�<�[N��\�iu����|�S`V#x@��&��_^v�r@�6]�=iv�;ڼך�Ө0aNtT�vvS�ξ�٘��w<9���G0u��t��]掎�۔Ӱ�t2����s�_c��5:K��h�4�U�j�)g�;�0��L]]2�Dfs:
���wܲ�Y��X��tR� �u�PR<�]6Y	������51�VM�dq���"��9�3�#;i�K�EƷ8m���ޥ N��{:QE�r�5`Ru��+e1[A�/S8��V�V�os\�o�P�倘��%��{�btnv�_A�!�ָ2.� W&��������ŕJ-8�M�1���]�yOOs%⭦�]�e�< �\^t�tԊ�=Km�����]ǴZ���p�֝9�A2��硺Zf�A�ǻ�gv���]��S3O|��b�>n������٠g�;]�61�d�9Xy�W�Ԅ������@>�&֭$:"�hV�J��u�2��X;+��ЫdX�]X�O����XǗW[�nVЕ�b@�c?r�S��5.~�âYe2����>�#��%b�0|x��9�h�c�{�]�v��j#&9�c�7�Ȇ�{��`��7˥[��S6lPޛ�k�ͦ�U��o��N�Yi��PJ�ϯ�wJ�����^`�#�ڊb�m��m��tX)�\�9�n]	��#}!�֌���DJw�c���&M����n�۔Z��1�뛐 ²hJ�̾�QT�ЅQ\�-F���A�b`��ޜ��k.��u��X�gk��E�Kh}-<BP��F�Wcy��p7�W_�t��]LC���v�SŶtx�Cpu�{N���f�E؏1WT��\u��-G��HrT�*��#��'ʎ:H���㇫�� |�s��͇�:��]Xa	t�y7�`�m�<�t 5Ь�5dŜ]��C�n)�w�@�����/%�]�e��o����>�P���g%,�� ����`ǃ'�ғZ���b�u�Z��ݎc���4a��D�S��9�b��Sjɻ���+nM�'/1"�nV�y��H����f
#�� 4"�K5g4hå��c�h~]C2��&E�n�Ͷ�;f4q*�G�R�Y��l4��s3h��W���GM�wy#�S�w�@�̹jP�������J��sq�O"F��" ��`�S�i��P(b��1�4���C�M3(k&��UbbQgI(W�Л&=6*4�1;���;2��h�/m����
�A�˝�yx^�c�JwQ���d��֔�yɚ���{�Ҥ/#݉�ī�癒t�h��b a[Ȼ��=lp.��W��$��N�7��|�)�Lo;��xX
�-��:��6l�������\Z�4��#�cp����.�c��VQ�6l�����+��+���A.e���%ٓ^q��m�L������4�?�y����{�?�~?�ϖ�QP��9q�]�p�M+�97*.�ͤ�ʪ�j�'KN��K(�Be9�!���r��P�A��āi�Vr�q"u�
m��U,��TUI�Is-d��/:B+$�RI���I\t���iS
�s9�D%�β��؋�㬸�QAGyj��w$�\ZdT��' ��NIʻ�*��p�\:���9V	�U�ˇr9��Ȝ�ZTzӹ��\�Ԋ�br��S��"���<��t��®S�Lym燝'�*�Js8�*�a4��!dXd2P�®w[K�8\���p�eS��RG������yr��$|dy��׎����<xg�s��O<��t5#A\��"�(��HN����t-\���q��j�bkr�ޓ{�:�nҏ�YA��HJ���k8�wk�\c��x���v��q�ΌE�Q�WL��)@[��ިϮ������y�(���"���Y���T<�-_q�|���q�~ϬZ�5L�{�Ћ ��l�Da���>�LR��r�ض���y��Z�G���m� �l�۔��{�n�F;�����7��h
 � ��Q�Bc�\����_N|���� #/�/9d���n�]6K�:���j��Y����Y@hG� ,��,v\��7�(��ٙN�,������{B�:ug`�Y9ͬ��p�L��>�%���Ҿ��u7��SQu�;i#�%���^�L5��+w���x0]��G;�O+s1S��d����v�U;�;�ʭ��7�ߩ}I}"�sB�O��>���y�'>�hw��_=F�_>V���Tmg��)�݀q,����}B�Tp�=	��U��T��Ra}�	ɮ�pW��{{R0ws\}�Yu��-� 8�2V;Dn�>��6'����c�<�/���C�U��9�;���9���+I��=��Nl�]P��m���9��ߎ���>���������_�c�9��sFM�u݈rfƺﲷ���.�:Y��!H�:�����wg�{�pk�{Wd<�ʙ�LBem&�T�Yx����hW]�W�;�nR����ٕ����Sv�k��B�2��yy�nH{sf��44�I���K��Z�̠�+#=���ߖf���(5����s��.�,ɜ�C����r�T+Kơd�_�$��hP;Jn3Q��ݞ ��3�EN�<�u/�6+O���Un�귑c����:v��_i����
C�~�z�:�09�EN�ǥK��\6�:���;�<t����*����9b��q�E��
f�b��횏�׹@��fG���m�N|�C�(xC���ޏN��{y��7F��B���A�*�}�?2����_w�ё��_wTM}�N\��PƇ4D��.����|�L<%��nx�������Z^��.�U;c�_�ɀ�ݮ�I�*���K���h�5a���Z��P�:�q|�� ok�|^ ��~��/��<��oVdw��ˎ��ybР���}܈�5o�i.ͤ\��7��-Hҏb�x��t���V��^�(��訜����2����T�y����k��H��ҦUO$O
}H�����Vz-]�8�cZ�Q3o&&�j���5���U^�ߝQ�g�fm��ŌC]�U{�^��>�יi�Iw��W�6�]'3Ǘ�޹]Dg�S�wM0�{en�piچn�p.�0�:�V�]��Y�%{�z��H���d���6��A$���@mc�eNd�/�{<tsw�o@�^u]N;��Ud���n�{���uyP�";�Ҧ���ƀ�<��䬉�)����Df��#�o����tx�L��{ر�&�/>{o;j����B���l��$= � �V:���ʬ^Ϟ������rZ�/��Mc\/nbiuvzr�˫�yl3P�j1ǔԦK�l(`w8��Qa���s����]h=�Byg�$mz����Qx�fj�Ps�|�����UC���}倮W_-ۯ��r�Ư�q/UϜm��̽�u��l�
�Ţ�ٗ��3��&�<�Q���w�d����H�/eJ����SĔ����'R�P��||[�@��
'l�4���=�����Ķ&U�ܨ�r����~��ŉ�>䈵�V�Q
m
��χ��+�0*'z���I�e�n�����{�u�;���OFo�:nω�fl_��\P��ա��XY�|� ����}��p��rs�ѽ.��Xy.�z���Y=��z�y�����z��Q|Y��yLޚ��������L۟��67��V�p:��X&��q{�U��kC�rx�t��ҡ��W<��)����0����S�S����w��ȥ�O%M��ק�0#�Ѻ�AK�}�w�t�Qg,���=u���Y�O^�*ˣ�qik��;�soچ�;3lѝX0JQ����:)�mF(��^���.��(`�w�Fd<є��=��nr����?��y;���I/t���r��&�]6��C�4�&2��u���=Q|����|�o<�e�3�D�ŭ�ah�X���2���j������l���G��ǘ6=�w*�j�t
���y�a�)�@jLN�QF$'Ց2}쵝�27�5������dG��֌c}o�:8��=�Ѓ���X�@}Qe��!D�,@�+4ؗp}}=9
��/�K��)�3��,^
�	殽\��Y'=x�/"�_�dN�Gm�(��HSs�R>��؈�Q��Ƅkm��M�W��'�'=R�Q����1��ΝA��ӓQ;(���R�G��t���^�<��ނ<0W��>�����fる����*J��\�&���(z��T�Ng��@����C��I��F�W.��Ǭ��#�Y��}��/9 ���@�t���f����O�3��#ilw��+���?���G�����Ϯ� ������y�
��ދ�7��~�[��s��ANQ���ڒ�)tR�����>��>�9���}tH�ȋ�s5��9
��	zρ����}���\�N���bV�VJ��y尫bl��wC���C���<�678XG:��/8����H��d���{�w뭬����Ѩ��81uc�Z��V����'����79���gKhh�:��KhJe�DL��rU���&��15P6ʥK���ĻR!�����꽲^����;��N�x.��x�6���?�Z�4���Z(�ݙ�.F{=譾=K�'ǫ�d��v�x4w��C'릢\g���H|����?St�u���2���fs��3_�b�-[A�;��������[� c#�u�xS����=��d����#ƞ�\���� )\]��k��d7~�᾵o���f�V>^������*��;��{�b���yd�r��� ��v��dEڵ᱂�e�Ǹ��ܥ�����|Z����y��Vґw�7������Au�p
0�� �Q�T����:W+��<\5@��7�%y6�v�ւU��Sn�yU��a�<j/�@޳:���s��V;�/���೦K�>���Pw�i���+����Cv-�j�D�u]P��E���TY@h����4��+G=j�t��\�[�C��O��;��Y<���;�Q<�鯟M�ߦF��jwW�g�}�b�ܳ�jT�dW�F��ws�w�ְ�+����+�(�t��럒��r�1�ڟ��l~��y"�N	y���%����}.w.����%+�Un�,���yo����ɰ�+y'ǳ72�x{�A�sb�ZH�|Zsbգ��sE K�]���"�Է13R�V�U�D��&d|/T�mjb�ot\��vpʴЧO��f�Ҕ/l�O�*�Tpo�<A�f>�%%DfO2d�9�`r�d�3Å&5g�}Qu�nVc��=$�g��C!��byͅ����J:��&gBrk��pH���S!I���!k7�v�����C�S'����{w��x����$ǆ����z~����8��q��1s.;&��kQ>9��z�[�S%C�d.���5�4��ˏ��&VZ������^�L3ڒ����F̌��w���l�<�Q�޸���2g3��A��z*�Y��f��������ݬ��&�ۭ'��?^bѤ��:�y���<(�����4;S����d�L0���G�̺�7ݰ=n��a�G =5��5}�@O��:�o�I�g5��\�9�b���V�>�����Uſ	��TS�lׇ"�']?
��K��җٙOܹ�Zݻ�s�$�RY�6<}L��׮ć��e�cd��ڜ�l`�K"<�(+�ꉅ=ޒ�pj��n5+��x����]p̺���a�x0��2�W14��4�w�V�w���˃��z�0e�~b������C{v�@�z���T7�k[�g]�.%���j��׭��dk(�&�X��A��I0���ֱ�����W��y�qvsuȉr�c�;@;��{��l�j+%C��<ֹ�r��}���|a����Zu�����&�7��qy�4瞢�W�փ�P�����6�u1)�T8��M����o�7��M�i�t~��T����v;����t�l�[�G��W��s�_Hzk�R4���%�T,��Om_����w�``�9u>�Y�I�/�9��i�R1�L��$�Y~��O�aqf�=�lfb�� :��KϵR��ܶ�^u#�O�;�L����#��A�<��x���f�:���Z^�R�#���P�����Df�?��	w�Ћ��~����u9�=�g�f=�~���(�(|�wZrj"u"�(`�C�>��j�x{�h0x="X��%ލ��|)�}~Cfk�����D��06]L���n	�0;���G�^%�dk�n{FNǻ�А�<�`��J��C��J}9�PʍquOW�e>�vi�eCq��q�<�����>�܎�1�q ���!eb᤻;�@�-�L-��c+�~���.�D�r��Y��$.��ψ��
��
���|k�m⎨�@S�6y̱�׵c'�Ӗ�zvګ�~����5.)���>�����}�+x�L�lucz�gb�Õe�H� �j'��wrB����L�F0���x󓡇�聨��Y������8u ����񹵙Zu�F��w#�^�Y�J�w�c'����)��8�GG���C\��ep��N�x+St6���|� �3Q� _���"Bv��Vt�P�zj��ܽ�磭�V0Tv3���=�[�2s­����Z�X몉��ꧮ���M��/-af��o\]�+�myV���yXP�����C}��^GJ��_9N�-Lޚ�t��������N:gFgv��$'��+Ƙ���/Z;K�jև�����=_t��
#':��5[�!�>�!6u>]޲(�G�*�� ꠭�q��b�/��c.]���=] ��}��̴59�X�߫�`p�:?�b�~���Z����?���=��x$�{/j��7�o
�>�5�풋�!�S e�5��15 �d՚�ֳ�F@f�F�^���ˣ�c��zv��x�AU����3�ϩ]����|�jg�(�K��;/瞍�m�]��P�[���Ν�f��=>�u�!�u
��9'fH�ϙ@hP^�
&簤}���9;���B�`�Ӑ��=Im�J�G#t�Z�{�`y�Q`w;w���$�^��&R�G�H��P�j(T�kTz]V� ��O��:�6ħ����̽1^�w"t�
GA8�f�L.- �+z����v�;�/�T:�C'IC����J���g��m+�L�y�6�1DHw1��!�{���i�-͛��PPN�`�Hcj_HC�NU;��e��}Չ��ܾ�:��Lzˏe�7�Y�����`aweT=�����}=4��U~����VsD�^���B��Z��B9����=�<�Gc��Y���_4�jE��f�{�Αu�>
��6�2����ף�������u�.��^�~�S;�|��M�ػ�1.�[�;{��[��l����P�؏����_������ӟ_��pә��}�r!S9k��lA�y�:=��q�NS�/�9���c˵A�Q;�����X���?/���D�鉖�~��y9~{��!�<�eۜ^��r�u���gi{D���FG��Ӻq�2
�f)�]��G�g��7�K��^���8��-]��9*�=�+�|���k��O�7Ǿ�쵛��ۨК�h�Cv�7�k��zP�;��îy���M�n�/�ǭ[�f�qNw���t�1���̚%��T��wnf��A�1T�i���H<>���M���]ׇk���J133�C��r��W-�e���FK5oQ�<���j�zb�L45�Z�ɳ�<\*���*7�M�3`����㻸�b@WYȜ�/|&�[L ��;*_��A��J!��"[7�]����{�� �U\�λ�Ų\�v-Ž��b)��/r�N�r��R�@;��/x�*��>���omP��kx\�0>��!�ш�r\N����F.dm�ax!��ފ�^���_��f��@ޯ�V���7:�������|ě�_8�S+`�P�S��Ȕ�s����|�m�>-.P��E���U��� \��<�ҿ@�W�Y���1O0��g��T���s+�ா�U���fpx���X����H��>�%�L�'^��c�$���^_g)�!�.{�h�~G������&�������z�*�*s�e;�w��} ��P�7�ΓJ}�Y��}��bH���&MF�@c���E��xǱ��s��y�$�'N�I�2����\��/B�Gn��$�K�S��j���2�n��N��~�ݜy �~�=P� rʪ�'�@�=��R �[���^�Dnǂ��&���F-�m�o}�s�؆����3�Ρa�v�z!�)��Z"v���a�//a���}�.�eF@06�}d�T�j|o�ӑԬ�ϒ�ޭ�*A����c+��qw�d�g�r��QӹQw^��w�vW�.�8�W3�Dz,"�- [�cI�������<;�+��#��zN�uU7 ��c��Jv'����p4�)mq+�c�u�T7$�@���8m������qV:�L�.��`���
�p�7Z�e��uz����Bu�:��ݼ�f�2��9cZȦ�shɱ\��]��r�,c1�r����Z�JJ��1��3�r,U�o1��,���ʗô�9;c�ҺIR��t��A���V����6�􍚹Y����5-94f�X��tvm�%�U�3%�dMGj��(���Mއ�����hln�<k�R`��V�G�
����;�P��N�[���tt�K��z��ȓz�A����8�+�{�7%��Q�Hϸ�j#�D�k̴�cc�Eն���CR�o�d���*Wv�yB��F���P�f�.(g�ڴ
�mj�0ڌ�g�q�N
Y`���S(v��n���i�)cr�r��xLw���U[�^�|�{V��%� 7}���)�;��<�/��S��V��Y�k5�����A�W`9��T�z+�����Y�Y�U+W�ݼ�*���-7W&�$�e�s�nl�.H�7�����ݘ�F8"W/�Y���/k�ȁ�4�,���JyO���,Y(������lt,Y��������t4�:k�>�maȦ��F��S�C��s���/�&����GJ��m@l�V{6��)���fF�MM�y���ĳ|5�	%��e4�9������it-M���-J5y����~�X�;���]5I>��lK��D�Q�b���+l��l��U�X����������}2_R������R�Rި1�1R���TB�u��kmP��;��;�X�����p��kByH��O\���}/xq�}(uku�V;/,���Gz�E�kyD�����-b�ofN��P�7����G��C�we<�1��e�ϭ�����<�u�����Y�]�'>Y�w�^�F��>r�V��*���(VQwJ�j>���m�&=9NY>�N��|w���Ϋ������FJDm\œ쫆�F�)h�5�o��ᆻ���f&ܤ��74�oz�_N+Wv�Ks��%;���q�@oa��hjW7,��+%�]B�Qs��X�Q�i�ēdX���\9�I�e�=�1QB�*ޜ%�Q�@�5�s4#i������=]�5vN\�8�4;|��YN���;z\�Ȯ���o{wX������܃.=�WWQ;��.Ty�/s��J�������Lm��{ *c.�#�P�z�%�������m�Μ�� ������&3@���Z�ul~�,4--��u�}1o����Y��c��R�"�ŋt4��{Ϩ��9n���%Ds:E+z��g��ST�Ɛ��}r��lp��l��l�g%�ȍ��y�9�J�\�[�fi[�`]�W:�G6�@�l>�Ta�2Jy�h���-�_��q׷�0O%�V��غ�c�^�&��B�K�`��b}���������AH�:��*0�ή����RD
R��
L�C��R"�(��㠜�뻹+)��ݷ�]�	<�����]�����/�nI�ʻ�u���^C;�Y't�+���Oy$���Gu;���cĕ]�9G��O�8����Y\�Ar��$�$*���g����Ô5�� �֓�]�Cď!��UX�X�y.�E<a���Ą���M��G wVb��H��e�z�3�>!�<�D˗.RH|qfg(��D�ΝVY�l�=)���kW^>9�e��"��NI�dTC�p�����Q�;��*s�������ʫ��<��**�� ����N\;��D�z�T2��<���<�dA�g��V{��Iu�p����N�H��'-
��V�ʪ.k�XU������7t���^�`k��"��^\y���ȉ"��az��qϝǋ�nT["պ���*�9�]�s���#��Ѓ֜Q�Ue�]YE��Rj܂�U���|O"bJ-
$�Uy,���n����<�\S�p�˕ۢ<��!�WtK�)y�M���*�L�-��/L�D���r(�8��%vn�c����sX�sh�=s8ή�Q<�$9ov�������n�:����^9ʱ}�1��U��x���rq�2*up�7�*L{=��ޜ�~ٴA�ʟ=�I+����}�lx/%�'ſ	�,�V���\/��ʄ��?|dWs\�����h����5>�Z��o��y��E1��bCb�Y�V����S�%/zn(���P��@�vpSL���r��x�>���6�Wl?<�v�����l1���%�J�0�cЦ{�IѮ;ہD�����>����ɿ����sT<���|i�u��\D�f6��;�4�r/)e+��vf��E������v|<s���}ȏ3Qo��uU�72\�t���NE�ʹ��{�1�\�|.^��C�Qu>P��5�=��g�`�6�F5)�x��G.����3�X�_f��f�:�����v�����LM��F��w߸ =�0�Q��U(��m�O�o޼{T�@ە�--�S��ĩQ��R5�h�O��P��U}�=��&��k>����L��ώ&P���ԅ�
 '֜��H��=�X>�vi�����whݙ��/R�J�ۺ2�vw���j���2%��������bC|�֌��8��a����o;'t���&��9�g��k��7k������k[��S�ۂ��Ԡ���F��RV�)W8Z�3��&�̾�1���z�h�e����̇X�s=Ł�ơx�8����O���&P��պ;j�SW|�����o4z��5:3��O�+ƾ�hq��T��2=���*��L����3�Z��4
�kK���J/�R����_��S��?�}nqUx��k@c6�&�<��ՊV+�.�h��L��R�)�=7�}��;�sg�떽dϏ�d��=m��s���^g�����z�+���狉tqeurK-�%���7�Îd��gV�&��zH{5��7�Pq�q������dp�9Q�wX�z�yh�u���?C�l����r�ߡ��X2W�?/���<z�&>�Χ�%]c�{���n����L�;�"�/�'[�;��yXP��{�)��L �\k����v��5LM�#��#܋L�����!�G�PQܸMw�����>7�V��xm�3�z�㫇��K��,W�O�ous����)��U��7�R�
����6��C�4�_������)�>��Ŗ%g��| M}\� �ﮍ��
��fR�J�vS�\5@�do�	;���k��{��LQ���Zp�n��ԧ7�cWj�z]���s'u�di��S���~:�Dn3� �p\�Los�]�4�y�@zA�4�G��=�T��S�3����[/H��zZ��wP��ڔ�X��D�(�|#�x�Z��{\��a:��/Z�n��v6ϋ��z� 5@�Pz�&�욋5>�E�����"_������Vs����ɬ���U\P���<i�H��P=�B��X&�|v��":�dJ�s��D�?w��A�A���GHf�9��zD5N�2��u";m���z�(���+��l?#̛���/��i/U��ؗ6K���p1^��kf��}�2)�z�D�^��K^&�:i���T's}�K����T�Y~v�Wے��t�g;����@�C�E��Nd��P�tL�֮!�d�p9ߒLwer�~���>����GV4�j/9 ��_4ʎt��t��1������e�>xפ�Q������X�ع=dٱ���(�2�b�,�S�)�fd�=�F�S{���=�վ=_�֑���	�_�^������P����d�q�S������0��?ef�j�×��_G������z=Wm�HX�����|W^{�� ��}4�u�3��ݖ@~�`��ͨ��~sq�l<��y��g���6���F�?z��[�#��Fc�:-yN;x8ˀ��!G�����~v ��\Z���棄z���8n��&e�K��.�c�8��m��fc��Y�rng͉�M6�";��E��X�ц����.^�.T���9��:��u�LK\���wSO��G�V�R��ݫ]��ol��?���]G�s��WxVZ��uW>�y{��}��ʕ��`f��A�������RHH�:n��q�Z=��حC"LgƫҲ���tئ���G�[�f�qO��B{�{�	<�vk��'_�����$�}�p
0�d��Uw�Ln
A����������ϗX�~��j#r�8��g}� ���FG��BCQ�3����Y�˪I�oN�C�иX]E���/���W���Ty�Y 罙���lxf����R��A��f��>�|�;4������.\���!��2�t�7~�3����U�
��E�����Y@h_��Ub3��A߱n5��٢�6R��s݋Dl��{����<����� ꃯ1`y�x�^[D�ݝ���M�m�
n^�����Lr����Z�z�8��+�(�t���'"zc�F��<;���Н�fN�u���46������PѪ���O�P��s=���RQ�k�i���f^��' ;�h���"y���S���?|�w�q�����}�����&��#�3;L֋��x��פ� r}C}���]y�%�.�MjRv��8�A���x�va��ۆѩ-�Q|
;76��*(���6\�Z�Nv�`����\�"
��0t5c�9�����u�Ǹn��A�<�@�������H���{[y��9P�K윀r��!�Ƈ�	��m�������H�4��=��8�b���)��������'ި��ƃ����fr��P�ֿz�_�qL���DN�+0øQ�$�}(�Z���?;�j�u9�������6<�-�ׁ������A��y69�w#G��Uw�\K<�P:6@���{���k�_"���& �x����"��up�7�xw��Xז�N�:�DP��C�#O�A�g���
��^YKƑ�O�@�� 1�d{�\7��ǳqfBR�W�쬕�;9�����>���F|{�`��o�e4��[��p���.�k]�
�~��+�Օ#��g-itݽ��,}��4ܿ�;�A��W/#�[w뭵9u��pT�ba9-�z���z�w��O�'�j}�Y����v�:��Z�0�\�8��%�J��>�x��}�>����5Km�I{����8P~�]�=ڋ9Qփ�MӨx.O���z�ʎ��4#��%���u{۹I���FE�t�a��Vf�;�a�#�������i/$=s���S�]�-��z��^�I��pW]3��Z���6�u�R\ƻ�ѕ������9�݂*���yW�jc��9�'*����m-��Ѓw���~B%��޺��d�ܢ x��1��;�xs���.�Lu�$��x�uJ�wV+��~ &���/��\.[3@��5S���0�=������>���Ê��z}�fNGyW21�Ƨ��f��N
�"�|H��D��옚�[ٯ��c�{�᯶e�<{��'%� ��n�䪾�ٗ8M1��(|���O$���J�K[����SRh�Df���<��f��̬Uo2l�k!KY>��z�%��߇(�/��D�95:�o�e��>������eG���Nw���/3˙	界�2=Y�t�wK�q�^5����S%D>�C���&��K3C�����%���c�`��z�&l�[��r�k�Ƈ��T��2=���*��L�V�{ns�j��1��1���*o!lY�EK h�~F���U�2�����am��}�m n���H�������~���T3+͞.���wO��|L.��	�z��#L�*'Z�>�-�~
��rG=�Q�[���w�mX��^��m�*p硤E�uhU�����G�?k�Un(B��=��ۚ���M�����O/�x���*s�s9Ho�h��+���_�X��o�x�*��x3A��L%n��s��B�᷽�cFc�y+Yv�[M�ι7z�鑶v��t:�S�=�R�HTd;�$����nv���N6GE���Y��]m�*��Iz/C$q�
f\B�+�l`�f�e��s\wݗ�)S:�8m���D8v�����}ݿ����Uw�{(����[�'�L^�
#���Cc�L ��Ʊ�z��g櫚���{�ܸ�轩��ԩX]��t��1�cَ|������(1��0�}��^�FEId�����ё>�O�b,R"�R�;*��*�n#}M���ϕ�{b����W��Gt\Mm<����6o;E�&�4 nk槀_`�2M23�����R�U��z����^����"���4���Ԕ�:;v�Y�*����ƾ��z� 5�@7�b�B}Y�'��Y�!=���Q�(狵�{/ϝa}��M[u)�S(W��4�$�e��2����{#w�F'���p����y��m�R��ƶz}��݁�=>d�7Q��:�Q=)�;2GnD2����Н���Bo��ޮ���]�f��Ǳ���H[�a=|e����xt�	�NI�$�5�qQ>��Q��籴���};��v������nJ���������q�E��uctx�ν�s��!���O����`ϖ~I1��\���?3^=�<�GW����@95� rm�cx��	���S>3N��$VN�(i󻣺pd�楄��oAl�� �X�����4үJ�W3�����y��ݜ���R�oe1nHt���ذ��s��A�G{;�����B��7lwK�&L��%���K�R�seǿ�붷�W���&��8�>�������<�hT��<����Vd�]2_�Dˇ�+�C0���"�0����䫲<�{�v�ֿ�s��g�gc��H��k��:�}�Ht/�'$^�MX"�r0Wo�>�ˬ�3�r���(��g5��<����~Y'3�TQ�n�5����g��u��]��Q�Ks� �38hȟr�9�+gԼ2|z��Iq�gi��|OeÕ������2�6.���t*��'	�K�D,�ד j�� &1�xVE�h=�wy>#�/v9�w�T��������)��i�tKQޠ�!�Uo Ԍ@Ň� zWDs5�����_���gj7�������m��wN��7}C�m���2c�<�@b�?]��UO�+��x��DT�)��~�qU��O۵,�|^`���D�r��_��z*�iw|�c��Fb���Z�V��G{KF}>��݋��<�|��:�a�"�E�H�r��=���g�g��=�e������J��F���X�Tk�;��jۨ8i�uB�nQf����E����|���΁qs5Nt��-*�K���vB�����6�ntr�d��ϋ�G 6���Y�0Yi�t��1=��7�vP9�~ �����m�,��H32zt�2V�t݊�]>�����Qʣ"�vZy���C��J�w���Wo.�ؾ/�N���y�]�l�V�]���k�G����~<�_X��n]�|�pdl��{��\��+��*�H����aE��ucTNk�� �B�ꐦ�P�g�v{���s��	���W�����3�ڼ��=9籛^]`�+ī��gܳ�X��:M)�)g0���:;��
�j��j�p&5��a�|���SSxѢw+I�%��SuT<��X��]Tv��꺷�8��T�����џ�b�����#��=X��=�2_T�� ����
N���R�i���ͥ��[�3Y�����݈.�.�WY�ǒ��S}���p�ޫndg�);_2����%^u_=�h���#�\+���A�*o�7��>T�ɭ�����Pkf�������qw�fL�n�A��yU�w+�x�G�8w��Z^4��;Q���1[3�EN�f�^��y���D<]P�=�&(����Iu':����R������f���E���U:�Y�!���킟��n�g���Z�̝�磯yp��+��Q8|�Ԙ��o�g�r���=����B���i��U�{Doe���v`vS��7;������X��R|8U��N��� :��1�}q��]�?]�ȱ��T�cJ���%��J�;7����9X�v�E��D�ɔ�8�I�rb�1�X�� ���Y�O�Y�6��M��O�5cBy݄H��s9�������~�j��f��7/�x۾D���c��2��I��� ���Cbm��E����hJ�� �����r�.9�C˂�釓��z��S�1¹�=���9T��Lv,�v{o��L�츥C����ADy��8�Տ�R������߸dk��N�8�k�Tc���W�z2'Ý���f�L��7U,u-^:^ϻ�f��"=Pꫂ�ꎪx�k�RJ��u)�Y�osM;*\f����Hҏb�y����iɬ�[3�_9��|/�&P�xI��j�����L:��S�����^��7�?���@s�I�K=����ܯ U��E�:]��[r�}��n��{yRv���uG���5�G5L�ze���Dv�2�m|)��.��O�30ki�'/�}~w�����v�"_�)0�<w�����Т�}iɯ�R!�F}��V&f����<j�����l�>�8<�ج1Q���X�s5�,wj�c�(��S%�Ib�1z��'(L����Bt(S���H�e�����¾�+Ưf��Ps�q���QY��=RLh�Q���^�+�c)�
���(�g*�+Cv��Г�u[�'���g�Z�R$�,�;�ջϜ��<�n+���3�t\:�!�ެ�r��Ύ�=v�r���JNVs��FvC�4I���$�a9�^�3*j�չP�X�V���u�����M�F��&Q��X��}��N���a��F��#g��ų7����3u�GY��%! �+�x8;�[����]�QE�j7:=�*�Z`����l�ǳ8����u��1[pF�ֺES������W���p�u&6N�d���zf�6��VR��-�ͤͼ鯥Ǐ	��a%�񔍺Ki��e[�-gR��3�;vB\�˥`40�P��p�K7h=������R��v#�ל�֮�ww(���ZЈ	��C�:M��U�ᰥ�M�n��w:î��j+���ɀ�\5u�hy�7hB�VVn��K��#AoW;y:|~8+&V+�����҈�k"�uk�ʺ��*o���4h�w���z���8��u���$=�a��l��ϱYl�U�*���X(�n���4� #]��ƒ�8T��q���Yg5��oN5 ��D�@�iluuֈ-k��N&�L�vF��w>���M�\@�(�#\����Ɉ;}��jd���0��w�+�ʧ4NNf�=��a4�i�j�V��h9Q71H/4��B*vr�u��Tn5(Y�)��xU�X��4�\�ڥ����ʹ�9߷�yc�EQri[/�E^�{�'fu<[r�P���g;���b�90�9\�A5��8|9���u��8[�bU�Pх�e�mP�np�Q�1p��0��jY�R"�5i�έu���2�A+YQ!�(Ү�F�,Պ�7�ء;���i��ӻl�������3�
��kw5�o�����Gjg^�F��\��׏DW�8�*���N�z�U��[|�`X(Ju�V ��4���K��,��(JD9�*ĹV��GP�{L:�J���9l:�5j�}�n���Z�wP�_D��%�[n��@p݀���W%�E��уAt���+w@��3��K�Q(�7�Lbm*�91	�K:#܇�i!;��B彠��cۇN�Ô#�j���4�˩�	D����LlU�*l�}P��Ϡ�U+	ҏ K;e��Yl�2��:�E���fS��t�>ԅc����ma�ݮmdSR��s",����f��c ��-ݣ���jt/��g�},1���iZ��JȎ��H�� )�\��Y����[���|k��;;YZ·*!j���Ļ�<�}qԋR��ܶ����^�� �-�u6�6��\U��8�[�����@(q�Ev�9�ܧ�f�\��=��'�F���a��N���je�,}R`���K� p�}�]�gE����q�I�뾮,��Tg��̮�p�q	0�[���.2E7eԋ,u3����ͷ��g���d�,��Y� �R)��w
ri痧]wS���4�4��C֑E<aDI�D������̫Bw\C��պ�����N�ۙs��+��Dn�ub�棺���X��8I��]�����ۢ9�M�"r$(��V����,)�2e�U�2��kp�3�ݠT�8��z�� ��.#��w;�y��k^wns\���R�SL��<OȊ�U9�̝h���.��+:���.+��I$�9�H����STJ�NVHQ��z4�I�<�PYZ�Bs��'%�yo��Th���yw�I�Q��C����Y�HRaN�{�� ��s��#�\�-Gw;.\s�8G9J�VUE$-.[�8y%ȣ�rR�I&d��9�0�	��L� �Y%Nn���	*�f�.G*C*ČTsȻ�(&(���rvʾ��O������[ܷ����P�fwq�؛ˣE��em�W����z�c9%���:�h�ߛ�f.�dh�NTRV��ݓ�BKaX>?�ȫ���aV̟��W�.�/ƷZ��$��E�9!(�W����F�Kw=�~�3���x�;Ӌ�ia�̛>���Gh9����IF�NW�K��z=޻S��f�S���*p�D[:��bx�����f�Sɇ��uߵ_����'��O�S���~����\� 5��'<*عȳV��z�my��i�W?j�e"��$o�W)�AY5���Yj�u��'�G�XP�{�t���� <�W�U���5n�F�gc���)��P�@�Q�#Fך�F�nk>f�Ǘ���VWK��6��N�� ��>�{��1{۱NI<�:Tt
��lW��=)���R��*�w������>W��NivI��k�[��9��-������������O|v��]>v��i�q��4���{<ߍ3e?�]�J��g��}i�6b���15 �d՚��qV�)�csF����h�˜��K�k�n��}��B��<i�H�,�6a�k��sDzK���޵���ٹ�p57�*��e��"^.�yc�K�Or����ǜ� %�����UG�-t��0����,3ioM��.\ޠ�������m<}�r�2�(�ʘ0Q��/�\���7IvFn��GA��i�ַ@�;mFZ�?.��:�ܗz��|����}<*6{(�m����zD5N�2��'R#����Zzf�л�a���K�._����;Q�D0��n��{~�,󛍙0���Os�:0ُd$�}��U�'Ө����oE�;�J/�e��u�Ty��[�����L�Ld\]g�wF������E8�^L�D��wf�Lo���!C�����_��ׯ~n��ɺ���J��~9J�v��]��6j����
Z,��Ł�͋�)��_x�*<�GHl ��]�[HM�n�=3�b==�l{��6�߲�#߬�l�ߟ4�_��O:�:�}�Ht/�'#�o��bqV���J�&|O�:r:��	zχ�S>��ڱ��ڡ�o�$�yʃk��(o�̍�{$K�5�^{�r���[>�yhm`!cΨ:��o\�y���c)�{i��@}Q�i]_�".��]R$���c����YP���_-�;},�������h=wy>#�/v9��z'�.��}�gm�ז�'MCS|k�+�=h��\J`��]��Dk��cw�~����
�u��K����@�s���C�m�c�J��p�k�l�ⰅB� <�!YE�����E�oP
�V]��X&Pc�����M9O��p_lt�-n`��}�v�|�~�s�|;�����.��	8��a��[n�!u������z ���Xݜ6���ns�±��=n�OWܗ �vA߮�UEW�1�)�}y)z�̼5>��t�ʣ�V�y���S�z����5���}}���W ���hw�)U%��}�u���7��>󔣲}�q��E����I��Z�G�7� z��<��=H�+���@Dp`�JV܆��oU��͜j����\��in,��z��O	�n�ᯡ�uB�nQf��D��Õ�*=q��I��k)A��O�&�Pn^��t<���*<�`��yc<��s�m`�;��*�5+���O�W��٥;*\f���zdiP^�
&��@>�}~��䯷Z�{��`��o'�@ØŇ婬��L���HȊ�ꪀ��U���Q�Q@o�n��MC�n�{�U0�۳3&��J3ׯ_#]��2\vb6�^D=F�O��$�ΐP�<��X��G�M��"���|t��;�䍧�]Ќ�Ez�7^��t/э�mL���n	�ww��h{=��QKr�+�緖�Y�>��P�]^9ީuK]g�v���|2<�͝��7TT<�Dt�r"`	Z��EE(�>��X�S㽿�|
�u}�[�Z��cM<�=���Oc����**u����q��Gɦ��y�����~WÞݚdU��O`�	*�Xt�;��g `�\(����G���d:6�p(��ڔ�9����PQW�ӧ�P�/zu_����i_H�>���u��}���c�A��y62���q|��J.3�$ϥ�D�ދ�:���<�vE���=�� {�x��ٜ�*"up�<�_�fB��]�n��P�WrY~R}���C�����]�)��Q�x�B=����܀�s��wK�>����/%վ�Z]�����:7�~G��%��e.�3{1K�5Fk�w�˰d(�iG��e���O�["�>�v�6#ז�Ⱥ��}�x�cc���Ҭv<l{�6�SJ��b��k��OWjI{�W�T�aY7�o"���z���?qj�ø��x�7<Iu�J���l�Q�3NhT5w�����S=�Jg륒��.t��C���^�Ԃ=��ǔp6���G�Mt���n%��l���@(M���R�oٕ�yj���~�O�ؓ�t'm^�A��O��;�j�I����{����H����W�{.y�����VZ��T�{�����KƀX6����J��Vy�z�o��cR��D�D�ԋ����s7�14{7�c�`R�T|b�N�@�*�ϻR�t��h�� '���QT)2C���U��g
^�fӢTx>�1�`��_��O��;7�s�߽�b��V���]W.e��fT�����4IR���6�F��������e=�ܒ4�p��k�݃��-.*����d#��(��7ܭ�:N��/�3�O\��j�B��rk�Ԉ�bP�g��}�|k���@@�3jY��7RI������N�@�?�(�/��D�ӓQ��#�:�t�u'ݾͥ���KŞ5G���Xb��JB��A��t�1���Q�<�/�]L�P�o�ogVFOeㅌ���2�'�k�_�e�����*\1���hx�����j��E�\��Һ�r�'���6.)ǟ�צek�vj:s*�/x�#�'Ƽy�勅F̿�u�1��-ʜ�3��<�6�3�|m�W�T<�z�.�,���_!�yk������3�PUY�(�z24����%���������:�X�o�j�T<^��m�*p�"��|���t��ܦԽ��j>���O39��d�*=�4���u���&=���*s�s9Hl=�[�'#­��ld��P��u.\Z��ڞύ\�}q2b5��+-[N��O���(FG�㔆�i���������h�x;�B�-u~�;uZ�!2��n�J>��ݹ�f�Ǒ�c��kCU�h��+�~�Q8��#��W��P{<ǯfT[��Ƥc����U�����\`���sKΝ����Ջe�;-[]��w)�7��E)���f�rC�W]ʑ�y�� 8e#���+�bC�9Cz��QS��dW $��4�����4G��X�p����G��� LT8��� �dP�ŀ��U��S`�ϭ��	Yr�N���6�`�
���P��w�O�+�:}�(���s2�z��19��4�ȋ����U���?~6�-{oӘ����j�#|�I��^0�#dxc�<�HC�@P똚���]<E�
�����ⵙ��E�r��F�׸�n��:�e
�H�D������a�q��Z��W]9����*��^��ȍ(�Q����m����=��u
��_�dR��]ІV�7�g���w� �6ԅ�ܼ*�*}��$��5!F�Xߘ�L����3p��������bNӺ�=�oٱT�%��|��2�
/����T�Y�;\7�Y�����`a{n0����uezo�;j����]@O��+^Vܱ$��5fTϡ���и���Uh���99��4��o�p���=3�Gf S�C���z�&B}h��'O�-Y�A�4l��cX�GԸ���K�z�Q"3{�}ᯮ�6�=�.{߫|2{���9u�������SRƾ�i��Wu�Eo^W�e=@J�>���$�``o����bY�s���LfK�q>����\{±�.��DWvy���齸q��﯋|!�-�����K��.䙦^>�L�୕�d���0�a�r�S���t�@-o��/��.�T�w�u�udmt�� L�F�d)ϕx��/gxy
�=/��X�o�$�30i����z}39-�����Xk�Ӡ�G�1|���dNR�}K�'ǩDy��g����zbU@�Cr�m{�Al�C��FD*��yf�MB�鹿7=�	Μfk嫴���P~��>AO����;���k7}��m���� 1��[�;���*\Jc��zVs5��y~aһ8����][�(�}֭x3�x��A���� �S��.�T]V����Zc~�H1�p�&�pzk[���+�د�p:���2*�K9sꇗ�c�(�c5�z����#$j=H�@އ5������>�k�`�K>���e���~j���,�s����t��2��S=o����O\8��s��I���zؙ�L���dmd�2-u����-��;��Pp��B���,�et��F1�F
�&��v.��|(e���������J�ó-�*<�`��X�z�&��X�+�%���W������7ة�r�=Y��j���u7[O�d�/�>�&9}�'%F�XDԳ�u뚉����~R���T�K8*q��3dEZ�R�K���E�Zr1�k��ms���u��yƭ\�;S̧3^*�*��%��I�![[�Kǣv\
޽J�^�f�Yk }Е�T�p��1gM�]�71c[�+/����'Z����J,E*�;ˏ#&\��П��L��}U��O+s1Q��d���_L��s�B�|x�zs�DxLk�බl�m�r\G\�&�|����=F�Q��$���C*Nx�O9��z:ἎDF_��kWZ)o���ˎ=UBr�t.��"��> =��6��@>��1�� ��9B��:,1�w#�ÚѼ����<�+%������/����|r{ٳ�Fꄼ�3x%*�
����	�︿q��q�7T��2�?��_����۩㛇��[7&�,�^@^�^�]���A'��G{�>���󫁡��~�ix�#̝�. M�Li9�gӫ���J�9?��p��������O�|p���XN�i{Ɯ��U�x��N}��:y�&�.};wTYz���/5}�}�G�mO��w��<a���w��S��6N�D��V��O������k�S��~��s&���fEw5��5K��GJ������wȃ�f�{�>���Ԋ
��k��͍�I=/�f�;H�*/#'[w��^�G�b�P�oa�3ė&��[�1<�������	}&�"�L�u��CM}�}� s&~��V�R��W�ӯ>�׳���v���wG���L���#�|4��L�dބ`kP��9��"f<qb�w��r i�jK���q�ui��R�ќ��d��+a���\�/XY���rP�Ɲ6{t����@8�<υ���S:5�*ơl����>��Yʶ����4=
����&�v��6����"t�G@Q/h
�ddE�)|63+��-Y���	nğ>sҠ�yjS7���x�p��S䏓�y ;�"8�b��/~)�<=�ưy����2��_E�Y>�gGf��^�7B��n�eC�L��y"xWϩ��@�옝��옚���A���~QQm����q��x[�xO�2z��׀\�2�}<��Q:��J�@s�B�T9>!#��9R83�m�J���������t��9���ӓS��e��g�:���F���΍v(��ڷƨ�~��Xb�q)
+93Q�,|M��mD��}��L=��]�{�yET<V��%1��k��3�~ܭ~8��]V��ީb���'�մ���q�n_Y�q���q�}�s�8�e���;5Uq�ȥY�����f���@#~�(h�V,f���v�*}ۓ���.1��m�U��~����$Ϗ��#L�N,
�ZXid0��UϪ�u�ۯ5j���h��_��V!-бSc��K����~��h�H:a�;���M�f֎���o�nE/�� lx���b=���7�˚ՓP�u8��M(���o[6N�|��o&�4���&�v��	�A:��[Wa��)�� ��&���?�0X�S�y�s,{*�/x���8s��"�:�*�6����~�Պy}����.NS�3��G+�"r)<~O/�x���*r#��Rh����ɋ��w�Ւ�c73(��Z�s�5lg��>��.��&j5��+-[N��{�ΰ���㔆V���(<�l���'�� ?z�5�U~�;��jn�SύԩX}y:�9�f�Ǒ��\����3VJ
OP�=���G�ᐽL ��W'�;�6)����,/U\��S`��eD��K�._w/*~�t_�Sq.냸�3�z�� 7���aΨ5��5Ξf�G?B�,�`�Wg�NŤ��j=s�i��=��tG�Ү=3>��葧�贀�;�TP�h���~2�8�|�{{kЍuk0���o�^m�>i&P��}���"NɜAMBu{���_g'<d9z�&i܋�!��_��ǧ̚��=�j�B��LLDu[��>��1�3h��B���փ�����P{%	RuК��d�9�Ю6g��G�}�}}���6��������cm�m�lcm�66����v6���� m���4�lc�lm�����6�����lcm��������|��ch���~lcm��lcm�66����66����v6����lm����v6����cm�m��b��L��r�"�\L� � ���fO� Ē��R�*)E"*J�*�!Q(RT*B��%DD*��	
%%P)$�	PIJT��"�(�T")$D"����J�T�*DD��T��D%QR*��Q"J�Jf��hd*%)RAU"R�U)Mm��	JUAP� �!J�DU	%EQE"���II%$H���"*(T�IQQ$IU D�@�R�!R�H�D#mR�  -N�
6����k`a j�4�-��54�Z�j�ʱB�T���Xj�km@�fkF�!�DR�!U"��G   ��P6�iS@Ը�� ����QEQEt8袀���t�tQ@PP��QEQEQ���EQEQC�]�P
(�F����Cl4�UHB�*V�$� �U�  c���桵-[i���1KM�сT)XkP�[ ؙ�
ѭM��iZ ���V�kTjX�MU�S $�QD��)J
S�   8��4#d�mm����j�i����0�ZP�Z��Zi[!�dj�҄  
�MJ�4X�����jP���d��(J��R�*JHS�   l\�UZ�m��XڴUB��U��`i�5F@[���X֚��h�J���-����Y[��@qUU ���JUD �   ��B�m*f�m��K����J �F��C�h�M[
i�����!��a��CLb��)@ZLiM*��Ҕ-�T�T�TCF�m�iO   w:�N�����S 4U���-`��PR���Me�hkM��*�h��M��[bK5���`�B�@Q,A�SZ*�EBDB�
IBE�  !΀��ƶ 
��6��Mi��D5j��h)Y�i�U��-��MZqV4	55+H��+L�`�H5��UEE�R�R  ��  3um�T��iTƉ�l ��+j�SJh�
���kb�
�PͳJڥowu�H�Ҳ45�LP6�ƪ�ka$I*�J�BD�UB^  ��[	3H����2JUQh`P�T!� �H�Zek5Z(TұZQ��&@��54��<�ʒ�j��S�0��� 2 6G���  O��P  ���d�M0  	4�deT  jP�bc���́��Cd$�MT�9V/@HIp��+sw�D��+���{��{������x�$�$ �	!I��IOԄ��$BB!!�Ns<�g���w��֡�Q�/��m�S�mXڳO#ݚ��ԃә����,K�al<(8�/o.�x�f���*]�Uo���LI:&
���5*�
Ѕ��5��85&Sv���͏wD�4%Ht퍣���h5(M��p"eY�nA��U��7��6�<W�*ū*�ѻ�dxr��� CaFÿ�Se,�2�Y��l\9b�v��J��jM��g�s2�u�x�X�x6�*#��l�P<S��Vk.�vV���՝a�M]�K3EZA�F�رH �v���w�0,�7X�U�Ŏ����bb4�nG���#��Eb,- ˹�v��;e��V� Ь9/I#(Ѱ*�Kk.E���m\&�߬�ˠ��,G(9e�Sa���3%�r��n���GC�
Ŷ���/s\ϯ)�bV�_B�EЋT�&�*�3!Z\�,�����T�'��wa���!gj#�vX*�T�^�ɂ� h�n�X�lF\B� ��2|��e<[��hbtD��yZ�����O㗙m^Sh��~X	%XW�.�$��wEd>*���	�*R�]�� Jܦ��W�2Ί�r���/6 ��6�R�[�����]ټ,8+V%��K��ʴ�Q��R#u}$��W{j��t0�+Z��A�W��ݺ+K��H"��h�u�
z���Q�Vh�1�=������� m��b�
w���'s7��\��,��P�F��㆐�u�v�GO�6���������݄�	%Q:�a��K%��%֪F̨��-eY���]���j���2��oU&�в�al��J���9��B	O4�CYkE+hh���ܶptD|����t�q�H�6����}t��*��Z#t��	�Tmm4]+ƤMV�u�������F�%lu�n��8+Ra�O/h�H�uux�RI!��S[�B%KQ)!�F�� ��7me!������\��m;�7Ym	��E�|S�̶��hA�7Ec��#R;j�R�?�t�W�/#%T�Kw,+I��Kn�*��k��-:�*+q��k�CS �QU����ո��[Vβ��`�ӛ��l9�U4�LN���ҍZ�	fl�(�F�ɵ�W�+ve���������z��ۗ��Hi�DH�Zi�a��*G�@t����d�Y���Mw@A��;a�`�dV[Lb���o~4�t,U�	�����a�Y:�5uX]�(U�
Ȩ�yb��e���(�!�5v�̈Q�4нG�T�&(%Ճ�AD�WXWu{,L�����<���w��HR�m�Kt
N�mv0j�$.��3n)R�����/+uT,�2`�ee
{�%j�CJik�0�� m<�0��$�`�Z�;M���޴0��vhKø��7%,H;�i�ɡ�t�Y��
@i���K+f� 6��,�2��EKu\��Ư.�v�j=vo�r��5<�l��kk°ƕ�w ���0��@��#Ef�
J��q[;jj鑼)�) /5R#!�]��X]�)��ZƷ>�����BݒM�^�I��yY�� F�Iř�^�6�ee�(���=#�yp��ZeFY�w��;�[�L$�$�M��8t��j�6
�.��GK�ڐ��[K`6��,F�u�oVa��UmX���D��-�����sl��"�n� �`I��5���!TǢSf=�؇̂�K�I��n롲��e^ZWwr9(H0�(�8��H�Z%�tK^ւ ��V��ݷPN�/U�t�E��7f�&���	6���E�%�362ĕ&n�j�e���<��l�m�l�J��w(��EX�r]�͡-9�v�4(��B�À�3EjY��yOi���c����3n�I�en�j����;X��yWVS-h1L`�ɫ����a���hV���κi̛��ݩ�ʢh�ފхޱ���A
�qɑ]�����B%�h�Y}�@��&��1�f�w2�[I:�Q`8�2�օs bv2�F1Ql�ai������^D��9):B����ӵ�b��`p�7L���wy���,�e<��B�SO@7pȚ�T�M�,�ǸlV�{t���Ĵk�Z!�kj�v�ڍ��0���4�Q�t�H�m�(47)Qy�X�U�[ֆ�dee��n��j"��˧6Q�FQ9n�X�7p(q�yw@C�\ҁ͠�DoI��_j��EVe�S
Ԫf���C�D�)�ܨ��O6����Yi͉���-�mm���#Z��#R��������cv�9�L�Ț߆8�2���~7��0 t`�Xv�|ɚrD�5��YK1��b��f�ӻL��pC�)O��Sn�6fQ�35\YISkM�܃i1����5flm�dU�i�K&c9�Wz�^V�"��MF�8&����Y��!\�Y�&�B�`yN�J��h�)P3��J��j�x�����5�Gx�W)��J�T�� �1Ng*U����v�-:V�A7�U�wo[t�ǏM3W�f���STxy�W��A����6VR��1nrh�� �� d�����Җ1�{�+)8C��q��v�7x��U;ǈ"��gS��2%��mI�Yd��ߒJhڼ�ׅ���]��l��Q膅�,^:�V�#]�����O�=��q��5��Ʊ�5�*�F��4�k,*��b�Y� �ͭ��j�#��-��qHau/2]��i�{�U^]I[��9���J�c�H[#��4N*_Z��Oe����6�sXk	ڏj��ͨ�1��MJ�M�M����6�iY���fTla����[dk�:�Kv[�,;���j��X��� ��-��q�<�)��7�E��D�� � ��B'���:m�utNT�53"8��hfV\�h�ǉ� R�41�f�X��m�1����2X���a]ܫuiV���ǆ��c�I'JD�K��1`�2%Ҳ�f��Lf�LVQ��bce*�`�X�oZ�ʳ�´�2��X�U�F��cl�UfY`	3uV�Wq|���А��2��Z��Q���P�"��3oT��
ww#��P]Y��dPy�#�r1Gr��#h��k����l�1�vЭ�`�EJ���[um�?c�zoi�&7ifj�t6	Ju�G�A���!����Z�xX���� 7��*|�@Х���&�۵$��hݴl|��=T����N3��q]˦u��m�
tU��
�EXZct.=m�&��E��d�n���9E�Ňh�6B�[Qmf^'�$u���1ne���m��Y(7��`�P�<@�Y�.�I��h9X�M�-DЙ��.��%k�i]������I������@0blٶ�-V�ʭ����i��D{u!Rm$Lƴ�n[�w*MK1jq]���t^���5ȅ+"�Y����<F6v�'n���*c�7c6�%�d�Aknݹ`ҭ����r�<�w�lܡ�3fn�kPx�D\
�9h�¶LZ�%�tNT���T�^W{we�Q�3*�Ad'60f�5r4�h:���F�j�C��i��2c;&�U�sv62��wz�Kr,L}��ɩl�K2�.�K� E�1I��lW4VҖ�SU��/JջU�t&*;u���"�e�������`�Ve�١"�UǸH׬���65"o,�x��@��Y�Y��)3v�/�N<�ݨ�[�襹!���ΈEhx�A%�"˼d��/#�6� FT4ع�EHM$Э��'�n�y�U��j����m�!�eڧ�v���Ap�X�j��WB�P��^�J87Sp�'(NF���\5b[j[�P�Ά1��\w6�4mF1�/���L*U���ѓE�;x2���51��On�n�,#�(`���j\R�;[u�ݱh��.S�%�
a�!�j��]���0Q2	o)��Z��*�(ک٥٠/;P]M���T,) f9���-*5�r,f�d��k.�nP7,m  
u�E��.���Y�Lt����1QШ���@/�^`@a�ņ�V��F��z�u��`;y���n޵*ق���0f,o+Ubʴ�Q�F}*�U�T��KU^,��i�]�rT�A�=�q!�u���Dಬ���j'�X�Q
T���V�,���� 'B���iU��p�w!N�h�xHT�2����J2��V���aI\@;��$�<kP�A[Z�f&JY������V���@�f��P�x̔F��aǿ^������� 1V�ݖ�ES�qo^�nVZnPXժqe�ݺ�d݃r���e��]˂��h�Ğ��Xy��sK �MJ���sJ"f�聂�N�NB�����Wn&.P���WWgP��Ĉ=m��5n=�(�٪�uPTi�����Ϭˇ~A���B�&�&�j�f72A�ڣ�k7EƖ꿓U�]r�iʹrR�	OQX�'�փp^ڔ�F���XV��`�⹦-��bk�)n��V0h;ϰ(�X������k(�E���cZ�W+TX�uJ��@��:�K(b�C0�m��4�Zu�.3G+j5e�BJ�3��w0c�IA�k4`Opk1҉�Y[�6��KР1�,�����`�M՛x�*�5������Qm?�^Vކ�P��2��&-Ԓˣ��̥P	�qN=��a����f���$9-�X�F���&fb�sue�"ǡ���D�������P���Z�g���l-k0��b�aWN��1��a�u��6����cjZ5�I�A��3H�9t��f;�4_L�A�X	�]H����[*66�'j�^���0�͂�ZB�A����AȚlvf> Z4�L�Y��HC5z���)伙�P�tN�<�qڣP��&���]�bN�4%��@i�6��a�2�����
+F�u��gE͗�i���3Z�&)\��^�7��
�W4%��B�\��=*H�s��[u��[�J��=�MD��
t�˽I��n��N��W��l2J�Xдk����["����R���45�/f'���� �VĶ�V�YGd��E�� �(���� �����`;�--��ȫS�rk7j���P�
���B�#2����.*ڻMɣa{�k�b�2�%f��� ��@�_J�VV]�ՙ2� �:ưLЅ�z��J ��͋�i-(��a�Y�-�B�b�y�͑8v�5�4~��p�N޳4#�͖�lC�X��9�$Ĳ�ij���������]��u�mTT���9�<�XXoC�V�R�m�Bi-j�[�CPˁ��V�6��E1���ŬY��s e�Y�!��F��[%�Tۑ3ou��Ѫ��[�,j2k�Z�Ukj�����hzLV�Bm���В8Ĺr�j	�eCZ�2�iWt�6�d�sc��V��IY;n����e��E� �]�	�ݙ����
{E�s)E[d/PCX�(SU��(H�Oq��:�tA�L6�*�2�/�[u�����$���{�;�����X�т�߯X�x�e&�&�V��7�1�4���ū�ڎ��l����,�7��w��ںW�n���+QXv�{37(Ma�@nR�S��x�ԣM�X�:-��ܷ�6� ڣ�=:ԙ��,Б�:u�)QM�x9v���&m2�V"���Y#�����Ȍ{�k.�7� ��)+PP��"��2�=��ӸV C�+��{3J�O�Ϥt��f&E<xf\ߤ��"�X�&��B�ʍ�hV=�rl��v���k(���D��ǧa������au���/I�q��/���j�sśa�V�������z��p������l��؍֠�X̺m�r�6q:��f�%�Z��	�.�û7b�y�K���]�a�XT�2�5T�4f��2�˥p*n�+7)Q릮���tN�S�V2� D�����){�hM�ͫ��dЦ�h�r�[�:قn�SBQL�V�Pp�Im��FelE���߅3��ͽ�-@�e�I��>�p��[t�㲂�{Bk������F����Q�ժvX��F���aQ/��݁�4mص[4���$� ���J�2<
�w��T�X�MR��kA�Z�Q8�]1C剌 $�4n-�9�^��<X�2	fd�K5�AEl����$�6��BU��� t�G��k-���VA-p[cFްj-�cn�'5��Or�-�
 K*�0�i`�u)�ۣQYS�%�ә�Q)Q�+U#��\n�'F�հ�.M�$n�Wyb�4��I�o@�oJ9�q'Wz��۫-m9����#2[��jj�n��k�r��:dk��p+Fh�u�;��J�$��x�J/���Q\���a���,�ޕ�̺�t3n*E^�����Ѵ�b:Ѥ�c5��]<�`t�w4�a]*��.��3��<�L$�Xiʽ���b��,
9q9$�&�:~��%3�cSa4Rr��E�qa4�.�X�q֋Z��na!E6�K�@�I��l�F�ڗ,�]M�a����#�#���U]�%�ӻsMh��+��
Q�L=��7J�͛�<�Dnͷ��v!M{ �/^��ܨ�MctJ�w��t�=xN���X��,����5�F�����<�kv�(fVZwV�5iS)n�n��$����mB�IT݉��VF��&�Om��352Gt��w��3T�U%�/XhE�v^P�m	��rj�5[U�l|*��ow-:�ST�It@Ӎ8�&�u���mݪ�,�q(����ƣHGj�I�C�u�E�je�T��b��P�h�rS*�a9x�h9D��N��s �g��+���/�����2�&1۷�±W;"�)�N��Z�6&�m�؄��63=�YKٵk5c��N;q��yM+ɂ+��ݮsB�F;e���2� �:�v\����B����=$wJ�wU��sR_�5�����}V!!� �S���¯�
�0r��K���D�p5�7�Hha��	K�w��ܾ��V[Z�D�7Yd�hYS(I��U����w}!���#�Ҭ���wV�]��8tZ��͢+W<������ab��=i*�J��7��f
Z���lm�z,V�ڏ��և��Ӡ�kx���F��{CM#W �".�bU�$CSs4�Gr���X6�XC�^��:��[�Z;)�A��E�n���q`Vr��������������v�oV|���o�}��1}��ӊVc����0���G]w�,R��w:v�����vV}��7O�Br�r�C����XEbtU-ǁ.X��(,Dݬ��y3hH_Ԫ�Sk�Ú�R�'6��]�x`�ެ���P�t���܅��h0Y����YS��l}u9,��X�Z7��De�>��Ф՜f�������\X�O~�rd��E ��z�5����csr���� �|���@�;��N	�[���\z���Rč���e#����2��s.�1ڢ�L(l݉��e�;� �z%Zۍ��ܵC���g�<^>ӵ�(PwF�/"�e��uaD4���L.l���-o)Y����-�8L��m�� ���{S��]Jij
�Zy!�Zr.�(��^��"SJ����0U�ݞ�e\����j���ϫ!�+-#���v��q���䤫�^��$�-��s��ա���]-��8����[�L�U��YW|xɫ��8��������#�JPT3[�+x���6�>���J���t:U����m���m65kNLΗ.Z�RvN{֊/�����]k4�Tx�+��޾]�lU�cv5�k�,����x�˒9Hh�`�c��XYp�ͧg��a
��=���v+7u�����,�.t��L��C"��=���tf;���������TՁ�ݔWV��dH�ّ����,u7���Q(�\�0)C��]*|�N�]q�:��L�찄�{���֢�_Ҙ����㲆ElSM�$z+`T�#q��T~�1+�ȼ��]%V*�5�}Wk{��04��5�A0`qa�Ȼ���D���ٝ�4#4�Oý�U��EWm�.6��H�=����c�p�L�I��3���I�k�����aާ*�e����������tvJ�N����6��
Y}�{�ykW�fn��gY3j�R�i5Y�n��	QGv��5٥�p��Wn���k)����F�K��;�;2J��]K�-X��^O��RV�kCCxq X.�/]�,<xj������>��,�]�禣̮�]ӻ�9�:���i�ς��]r�R��i�B�s��$ʽ��+1��Lef�M�[�P��U���+�kT��8��Քy�kVSї
�}�d��[@_X4F��0L��xi�{�y5�(��q�9��BD�g�Ԁ��+�Ne���.�tѴ	�e �`�l4���Il��'3�d�5Si���y ���� ���E��^g%��$ݠ��"�n��#�����~1����Դ��:\��3��=��Ȝ%�8���#(p��ly�*&�T�dWv�����618�l4����|{�i���g�ۻ����Y�S/OMu��/��r���ъ�� _TFη�(O�k�����z�Š0��hT��K%JH�h��-�o+�d�M�c��a탨�r�w2n�%^{�ox��X�F�=���.��'Č�l�h-�k~sKb��mE��ͺ���śV���Y�QwXƶ���V�4\�����f�X�vs�r���+��l���3H�k��t�G�y����2�,�o���|�젥�׿\5�v���̓�_��=1�8t<�񿵔4�O�_l��c)�[����*m�kb?��*V��Gt^ujƑ{�;!ݦ��aH�
�A�a��p��;�-���9�Q2WG2���ss�+������B��}���֌t4�/���ƻ�5JC����J�-����y�+�[\;K��s�0u-�NvK�yܓ��r����2-��_ug=��<a_Nü5�A��OKUc��}�����6��@G��|u����CK�K�FR^�m��ݔxe&�N��oVҮ�JX�T�onq&NR�����k����*��1�WRB>*��vp5�_d]H(��E�P>�;�fQ�����w#I1�`����-Qe�����P�\ܗ�0^Ik���u���u�h]4�ܩ�[˸hYݝrvM�`֞T�ӁM/3K�����7��h���כ��%�qM���j��! Qd����r�y�q�weh,��AʽV�%
�m�^V62ޡ����W8SI�N�<�Ϋ�����k�t���ٷm�y;+xu�ю��l���m��h����e�"�����	
V۰S�Ԓ�\j15	���}]��Y}��o@��Ya��]���;�wz|������y��O�C���G8�'s�vQf�AC\��^[] �a�ev��]:���!37�j�k��wV��[�y�K���gS3���sQ"efQ���V�8U����V�z�f�[�Z���\���/,PIYvf`�X�Q���f
�"��&�ˮ��tjdu�*st9P$w+�����^8hܽ|��AW'W��G%Ț�	�6�6N�N�u��E��N��<��mA�/nt(ؙc��x@;b�}-Z[���}S�u��v�i��*y\��jV�Kf�z�U��}�V�˵�q�/��Ta�l�=����+w ����z;jn��oP�S4�WK�9�����=�Vp��5]�=�ճ���v�M��뫋�i��gP9	�k�IG@bM2XW��(vwit��
JYaخ���=��3XY���<��b�
�.r���`|�bCi�gm覴��=X�%�Í�[v��ԄkS��zx��CuSsl%�|�5���@�����t�)��Yg�]�%I��F>k�ZEe�0��.�����o�ۊ�]����[O2�j۹S:�h��)�Y��A�u�GP�{Z믫;{����2J��iI1��VX�}NT֜��b����]����y�]�_X&�W�5�쓐��R�F�n��N���ɢv�9ٷ����m��3��4yK`�؝{�U��V�����K��ѭ{zp4�v�mCH �[罫罇��G�y�{�͐�I<�ڎ�B�D�z���q�v/A>�nk�_%�,�N�� -J����D���t�������۩��u!Y*I�i]m��T֙B������K	ѽ4R��9t�Y�u�Ӄ�#]�n�o¸���A$��ȱB���_�����o+½W�/5uq���&(�ٽ_\9;W&%_o$.Mv|):yWX�T�T��8)�Ln�F�N��mۈ��R����v��\!�b���nP\�$�j�c�����%���L*�ֺ�LYas�ջڃ
�-�7V�;7)�i�Vi*�o��!xiᱚ�ɳ9W��w��7�ХC�,��`�u�XMj\�
��-+ȓ��oH�NW��=HḲ��7
��$�������[������g�o�v�j�mA'm`,����Q�{�%T:<�(aWnk4�j���*d�ʍ�:���	׫4Y��[���Tb�S�E��}z�#j��m�՝k��-��9�EQ�D����W���m���r�GA7E�J��s��բ��
���<��#�s嚻�)NwodZZ�R�^	p�gV+� F�t.�/\�u����v�VNJ����"ͽ�§�}J�T�nXWRqb�KM�rgU��%��]YQZMN����y����r������Vi7�ব���B&_S�|.�)�% VA2A�n@��I�[�����4+�s!nw�f�4>���=�ӕqs�Ӛ׬lГ���P��6��<4ì��R�:ź�/`����?���.��ٱ�$.mp!�s�Q��gűzΰ`���e������v��dF\�P�M�S�T�]*q�R�᎖H24��۹�u�����f�>�]�}}�Ae�Ɏ���pgP:݋c��Ƹ�A=��;U�6�aF�z� -+���h���A�i��r���NI�:�'����V2��JT�Oj�:#(&�M��Dr�-����"�+X�9�x:a��{@���@�o)5c%�4D�Q�u�M�܋f(�o}an����ӧ��ֹ�+Fne�ǧ�'��hof+|��[ǎ4�1�p���Qϊ��ٗ����K�Wm.m�n��ho����U�]Ƃ�W5�v3������3o�[�4��8vҬ�A�v��h�w�;	��eZ�'j�G�5t�\����G�Qv:j2�fMUҦNK���>�*���b[y���\ �S�ֈ�`#à�i8��V7{���\�#�['eЮ��*R��1�|I��)b}lD�2f�9V�<��TR���Ɗ
�m��K���39	��aeº���v[��&/�pEӫӦ	�ڭ2��+���j��о��.��Gܞ���S�Tۺ��-�l!�p� s�r��|�K�4����&�M�������?��k�����R5zwI�N�EO�`�,�C;r���i��	���(Խ%Ұ����}��e�D�����bb>J��\�œwk�75Û�i��u�X������9o�1���vTֳ��p@���1�4�;����D)�x�V�8W%cT��m���)�O��=�m)40+C��ݚ�m_N�5��.F�V>�[�`VA�2����V)��� �rR�}�P�oc����l���j3_��/��9���J����m⡽��q@��9Ej��gM+�h���Dg)��Ƶ]��C��Já�(/^{��h[O`�e�v�,���D�ٔ]��^�\a�ͪ�\����S�*]HfS���ɥ=F{�B���KN��$����t�X�#�Ĭq���Y��@��kT2 (^�=��.�d�Dj�d�� mY��Y�\�t�$G6�bu6F ��	oL��&*��u��WM���̑l�V��"q��,�<|ŹY��Uɜ��p��&T���!�a��u5��1�F��e���HU���i��2�ت:]�g�oun�}Ifj���I�ݦ���PW��ő�D�ܤs��"�6+�"т�+�EK�=�=Ҏ�p��dy��)�v+m�J�9�-�����6__K�9�m��]�*WR�}X�5���sQ̬��ĕ+��2�Nu0��r*�F��o�J�EǏ3)��Vp]����`,o�`M�[�G��[G�����~��[�C����G�vP=2�8��[tȲ�n����� ��f�w�	���]�Qg,[\U/�^N�m|�т]x��d�a� [U��,}�S���ic+{x�k�K�7�c�+k��h��F�����Z�n^�@��Q���Փݡ23ʡ�B�zh[�ҷ�h�5�;C�"�h��Ln�rmڒ�(�ik۱�M�R{3w5G��7�ڠ�+i�˒�����-N��#[)c������;/*���]|i0�j�wwծ�����92�����7��d46�c�jK�6���V�1��'j�[}��u*Te���f۬A�*t�eDi�=W���u��\��i���8;c]�p"-� <t�n�4����={F����O$o�:�Ɛ�`�ΊΧ�f츲�w)����ڢlc���vd���e�Uj;������U��W�\�0p�_�t*�p�a�|�S;�o�R��\��W%ҏne,5�f�婫]�D
��W\�=�*9J%\��u�/�tv(U��לG={n��R�I ʅZ̀�{v7���0�:o+��>��:n?�nk�Lg��{�tu�����E��$��ˌ��ۡ�ŌY�f��m%N�gmv�Y��.u��w衼��c�����G/U��ʶ�x3��`���]�9l-�άu%�����]�Ns������@֑��V��8{����BWE�@���6��%X�lC����_n�2�/��MNj�\鎨��M�|0v��T;k��ԡ'WfI,�CknX����q-���1�E��ğ]M�"�<�(��,���rX���Sf� ��Ļ���a�lL���C�ob,eҾ67~NAJc	����5r3���k�3�0Eo��HaN�����>�;N���m�լs[A�w��%/�-�aъvt�@v�o\قrU.ޜ���\�����	R�e=�̾b����ڂ^��g��zMT/F,�4��A���p��pg�g�խG�:�;Q�u-;�"���f�Θ�4ٻYL�:3x��.�a���C`�*mٻ�$uU�
�V�#�'Pvv�&�|����{j�n�t���^�:s8��XU�-�Lo�N�[�9_,�LQ��0o+2�b��,Ve��pZ:Fg+&P6M�l����o:5�G04b��4z�LO�9����p"��S�5uK]��X\�����a��-3�f��7~�]J��ۖ����id��׼p.q$Ѯ�|{�q걋������O3.U�	�Y3����KU>u�:7W�v��RA\����zc��|����3�0�Y@w7��q〧��������|�]��9�K�k��1s���[�J6����$V*An,[ki.(ݤRW-�[��p�k�v����7>���=��TW�`�[��x/'4�umF�rMQ�iW6���F��W!�M$�@�W���z=���	!I��{6}����{[���u�:����9�xI���t��B���BաO�=��§e��j�$��8�=WM[0�vU��K���w]��%��/-T�q���9;2��e�۹�ʣŞUd8�[��Pr�K��ܻ(d�ER�n����W(��^a��n��^�Yi(��G��b1������(cV�]]���,ԇnW:�#%�b�����[%�!��'ƢZ��n\C2�߲�dm�ۑ�lj��w��(%]�U���9��=m�K�4��s�n>���^SU;���s���(��/��4�]����qշ-��}��mS�p�Պ�VA��T`ݍ���o�W�����{K�a�gê���Tec�<$u6�,�7UH���y���ǲ���`�XFe4%�1,'D��8��wR��+��f�\�(�.ehF��5�]��
a�x��Ә�hCp�Pt{��X��h�b¤��\k�vx���t��'yN��VȰ,j�)w��s�5�wWƭ���+Y�)h����&z�����K;U�L��3��;���dS{L�h:p��΃����N� /{�Ȝ����S�@?2/w+7[ӴZ|+�K���ͬ���ǻ2+��M���eStƪ�3��X��+i#�Y��v�/[C�O#Qv�GJ#�ur+���ǯ�e�}$��	9��*�.a�f��y�ҏ+����#��ՠ��oo{07��e�GY*(�vVV���s��/�l/����[i�8�x��ds��c�y���]U��8rs��t�N'RbJwk:�B�ǖ�q�qM蓮x�XVH���d�մ4���;���WOw\����n%n�֮�
N��Wnuwc��O�ܠy̾tu�C%��msÃ��`��{j�X����78�Or��ȵ�l��9Gթ�+z�>�����n����9�t7�٤'a�zƝ͗	���M]������H���:$j�.�����)�a*G�����*�P��k����!j�P��W��rm�7W�Sx�����'�j=]뙯�}y����$���l�Q�Z�iup�/�tӼ�`V�,�>\P9���|��1�ďee챈�c>�띢k=o��@t�j��\`��
�3{^}�b���qB3�({z`�.��&^b�	U�(����f��V[:R����:�2��j}��8��	�����,$��z�-5R�f�^lX`慑�݈�K�_J2�}F��q�%����FF����6
&��iytu�.Jht�+<(J}w�WS���E*|�qg-����c�H�zk_X'Y#^�7T�s\tT
[�w�]Ć�c��[yR�>@��TmU䲞A� �;Ɋ	��Q�N��v�y�M;��t�w>����z�aũ̴��0p���䦵��SZ�̇Z�,Sd`�pb2�T:3��q�ܳ��:�]+�n�i��<҂L�7'Zb�:VS��o6�������V�ɏ��rO-Tb7����hEǰ�l�A�oD7%m��.+��M�AVE7��\x�(�g;][���n< ���Ja������|���g>b��Rg��9JcJ��TV�� p�՟Y�s��v���M��#]ZY1bM<����w��B�/#�:���MwYz�`����9N���;�^[]'�x��i�Yhv�
��h*S�)��\X(�r�|�T�[-�%-��k�]m-�3]�]+CY[�����>��`z�3N�ܺ!����ʓ��5Y�Д��VV�t�e�RB�����VB�Qݖs1��Kk�HI�@6ٻ�/��^���=r콩�m�(Zjc��x�l�wTz�B{zC�&�LZ�d[q�.�F�<�\��q�ܜ���f����\�z�9!.���Q��&�4���/��O(c2��.�'��g@��ް`�6��y�u�PU����v�H������.�t�,8�1W�N7�5}.��\VW@C�h���I=(/UK�����[�Dq-�6��Q�xV�nv�n��V�&�2�ܨ���EN�6b��w�T��9�(Z��',�y�`mLN��B0��;��B)]�0�ƪ���M�O���F�\w�Yx̎vk�*)�X���5�mi�+b��j�z�#�,���z
��`��O�}
ql{f� {m,B���s9`�e�-�����ܳFaru(��w�{z.����"��ݡ:������ ��+]�9 o��Y�\��I]�%]�	�`�^�V�3^CK,T��Nq�JۥF�qӊ�ӹ.�3}�a��(�8FlQ�Z���6�&L����E"ky+����8,��O^��
���W8������0��݋*;�n"0���L"O�W�����z>�G)�Dݒ�����Q��Ċ.�6��R5өY��Ԕ;q)���ܔkf��G/��2�;��v�ܤТDu ��v��VK��6�U�j=�6�Vh�I��hˆ�k�9��,��o��\���=vb�ER�.���n�\aY�ԩ�>|�aNDF\.��BjFz�N�̙���E��޺Ƒ�{չ.�]�V)^kz�mhݬ��Ʊ��7x�f�V�]7Ri&�ܨ���B�U�]��bK�O�sD�쏲�C��y�br�&Pv�ҳ[��t2�@�e�b��ƾ=u�ϴ!�����-�>vy7 �r7:�w_.��ӭ�V�A���f�yYO�����:+�K*Wd�t���;iSeY�����D䦃x��}ɪʳ�b��Di}�n9L4�Ō����]o�j��d�Wat/RǢ��+�nm��SA�y.��)��G���r�
Wg��.^T:WK.\CWf��}{,>��p$�<�&���m�ye�x�S�"���C�\�Q`,��-�l�WS� ��|/el���ܻ�B�kr̜&b�RKS�K!S�_s]r�ys'�a�V��i���XQ��*hd�o5���rz�Ʉ�Y�������^٩K6���;:R���c�u�*��[�<�؝���y��7�W@��Xr�ك�ѧ��	n�{��Ʃ�c�a�
$L���pn�w���3�������=@�:� Z`�tN�Ou9���a�A�p���Q�r�x�Qq
���k���}6�36��{*��S�X�Q������uh���m���mO��֜���Ʈ��yg��ŗV��Y�GW�����\���#^r�����1�2� ��w�-v��/Żt�l��|4��)ǧZ�Av���O�����f4\�9�li��� %�|n�m�q8j}�h�c/V�
��w6����N��cw,�ͥp�����1�fW]��T0���L\"��XB��v�.b:��޳OMB�C9�;�d����6U��͂X�Ǯ��'�C��N�*&b�9tz�o7��F��;c�LusEu�'�]�tST�S5��tɽ�X���.WXJ�IsӾ�Q��Ȱe�X��U���qp�ݣ,�oqC�{j�n�iX�b	��9��٢�9���wrԗ#�s^��HP�'h���M���Ud�=ח �<J���d�E�oY����\��	�m��/0�o���	k&t�յj�#5=j0O�U;{��f�tL�"G�k���&��:T;��H���ۜ/0�AR���a��:b�J��:M2��/��T���%�m]������T����~��9���iuL����e�\���pԩ*e����ޥ�����g6�"�Kt��)�wL���Y��ڤ���XHS[&v���X)�S4����!�ȏ�M�s���"^�Yt'����K3m��*�V˨���1݁�U���r�%�7,ց��Z�6�CPf��nu�S]]mis�N�*��Ӌ�ʰ	�<c`���(=��(n'-�ۛY�.�n�zv��!��[� V;��v-�7��I��١���j�j89�6������,�[�5vVe;�i�A�9����7*�� ��1�cH^�Y������]���.��v`�B�*�ۚU(��kmʇ� B/�+�Wt��Bh��`݅��5�U����̹�� �So����Z�t
�����:w��8��ew��.}���vӼ�ނ��S9�K�n[��MЉPw�Jd��3���ݣX*N(e��������)��V@�s��DPf�c�̻s/+�$�*Qб^k����LN�w%�w���l��c��,�B���p��q1�^j���1*v�N,�����౮ZX����7/�=���/(=<N�Ve�PCp��
��9`�5��<�q�\0v�M�W����sF�뜲%M�M'�ʆ�W�����X¨gc�u.pj=�$em�J��5�7c�n�}������v���7J��o��WXq������ֳe��3b�u�WgqΫ�v�ߎEY(��|k���+=�e��{)�d�_=�\�0KI�K�&u[��+����qSc1�1()ʺ�#V�'�����y�\RU�HM��t7�ӿ�f
�v����6�=ʾ�4���β0p��J�Xi��-]v�Cu�g��o��j�lX�x`��L���5� �w�6�o���o�
�}�1��m:@u�&��wn.����5�e�/T�P�V���N�lٔ9������
�� �+�Ce	u����M^��&�|��R�2#N��<`�HL��P
8��W�ѼZ櫁�v����&�ur�`ҝʰč^�h�~�-�eg-Ӛ�U@wt�ɂe���X�o�
�6B����`�V���ZFֲ�v��ɰP��-6.ۏ�b����1-��h����[��H�]�&��N68�7}|K��F��l%,�'\{�ld�/mލ.�u��qe�j��(`;�:�XgU���;]M]��i�,�5I�U��:u���x��h�%i�baOv���h�R��^L�t���U��Tw��䰰"%��Ug:�gk;:�{u^��TZ�$=ӯ�xt��o�3C����y|�P�
+�\28Q\,��M�/v�\�ɧF�;8��`d�u&F��ݳPel��F��X��ina��v{�j��c���]1TJ30�M �9,�T&c��ՔC��]n�.�|EY=��N�˟�.M���Q�ȮD�U�ݠT�m��.:ùX]��M�'%c��P}��#���E[Yq�N�������N����Y��sv�T���*������yv�R�Lmyiw./�i��B�7��R�Xe�&*��f)ژ���p�ե'HFu���wY�-ӈ!���]Ʊu�!jƘX̙�W����B3P����5�)�T���(��	]9G����-����I�*�T�����̣�&4�9e\�Jn�
u}V(dh�D�J��n�W֢%�u+II�X�2ljޔ�

��oUp���K~+�9�C����'��-#}i!�����t��]ܵZ����۴��a��I��3d��yP�ae�� 	,ի-�o)��ݨ)7����ؠS�GMɭ���0�*���K�do�G(�sskI�9-@��r�����yK�� �g1��� ����Z��ժYԐ.�cX������t�y�������$o@Yz�ڝΑ��UҴ�Ԅ<嘻p�٧+��H;+r��t�u��W�Z�zr�7mKe�]Oc���&u#�`����]���w��Oz����hw]��Z�Jp�W��Jt��n�Z��ſ��K(���t6o,QIuZ���8�ͧ�{��[���r�w��%n䌼��ʾ�k��o$�핚����^����`���bP��*�����GR㽃���*�)H�nŞ���oU�Σs�XXޙ�P`��#��F�-\Fİ-��T�h�Z*�A�.�ϻw+������)|B7ԩC�Z��63u�}}"���ë�z�pS�Ə"�W]��q�y���c��
��Ѩ�5e������9�yJ$r�c��g^*BJ�u��x4�t	�,�	p��݆�6U����:8"��u�ܴ��1��n�B�H��+pг3�J������T�*pU b�jR�[�V����c]�@7��/��m�j ŝ�)"_V7�6�\�c�'�����*6:�uhՆ���K ��΅��	5<P��N��Ǖś���8����d�Y)=�J��Gһ)���L]��6�J��蝐^�����/r�Li�Ei{X�Mj�i�$*\��VXe�B�|T�z���*�M�78-�dB(�5��AwP�kk�ɖp���S��a�4u���뫱�Pc/�^W_���v�I�1h*,:%��jX&��ܬNoR�ݽ��D��'FHdW�n9����ټ��ki�p[���K�֏�@v�,cF�f�4)����#�-3Ω6S٧����0m�4���>�>t9fNSEM�ܯkq1L��G�i�γ�+d+�x���b�/��+(m^`T����}�<1R*�<���S�a�Ǻ�s�5ҩNЛU�d�+6�"��+qs��ے)����'��N��&��ѣG���b�Ǧiqe�"h�����ZInqi������7(Sb��qq��gK�Җf��.�Wڴws{r-�cqdU�1���'�d�#��I����fJ6�^6)��ZJ�v�w�*�+]��s���4���V�v��ޢ��n�}ż���rxi-{q�%;8�y}Cn�XM�괫����5��eKu��e�۷�xA6�Ζ�0�F֊�u���g_m!�kL�/�g��[��2���:�ؠ��ѵ \�H��;'[%�HGc.�r��P9Wn�+W,�N��nQ�LG}�K���Vs'{�7��#XҢ��1v.���_u�G��{��{��AE��J'�d�-�3:Cmv"����h.�8$�`��\��â�U��ȱV�v�j�n�{\�\8w�W��vh��N�u�U��μM;��c��ς���Mf���y�d��yP������{h�kwT�uq��)���u�敡�}��;�Kw��t�b���-�ﵡ���%ϧ[�P�2�س��x#R��P�U��,�:��R�M��f�U]�\�ٹi`���P�+A���
⠅u�%�ά:�u0�W�QL`:W}�1&;�Y��4J�4j�&��v�E�V���WY\��ހB4��W�m�Y�l �K��+����R�Vwk�������f�c[�P���>�5��H�+{���1�S5����tC���Y��Y���\�앺�����H�ְfTƲZ���[�h
uz:�1SQ�.���x�]�w���\9��:��7��\M�{�ń�1�n��i����P�v:�S��ύu��k
S:�VٓN(�,�BE�ʈa�{Ծ�5��C�!᳌��"P!�������"�i�ﮎ�7]����͵�\jb�'N���>5les��hf��]j�l�W��A}��ǆ�T��:�!e�z3i!��2�U�(ҕ�5ە��u}�E�+-�CYĉ��+|և��x�6�ӝZ�:ev�̶�]�}��n����6.�=c�0�E|>@ (
�QDTV(|�"���,�*�
"��5PQJ؂��V�@�H�cRQTU(��� �H�A�Qj(��	R�kmJ�F���Pm��)n0d��j�QDqj���
���
ť�Q\Zb�QJ�jV5�c(ی02���0ap��V��1T+\`�)Z�,*ږ�1��������
ѢRЪ�[e�����KI��Um*��[K��
(ڸ�C[#bՋ�aqX��5J)iU���U*�E\�b��EIZ����R�B�l���-�(6թU�Z���F�����3e8lDb��l����Z+
���)l�me�[m�0��TQ-
���-ZV��ʢ����(����1���le�*
�4���G�2Q�K(�����"��HJ�� H�Ֆ�A;9�j�І����*��]�0˦�l��0��*���v�j��Q��Uib��z��VaAnp+:a���Dw2gu|K�غ���|�σ/�N��O�Y�]g��o��1K�z��
i����{*��*�������|��<�5h�5����A[���姌�~�0c�=�e��V�Y��n��>���%�UB�x��q7F�x�VZ�����<z\T�l�K˜T�lZ�f1=���y�:���PkOU�9�g8�t� u����)}�Vo�WiK�K��uYC�6z�V�@�9J�T6�`�Lcu3m`�|F�#��U�V5W�Yq�Y{��ܐq�˹m���0r�՚;�`\-����BX2j���22��t���8Z�]<�r�/_�Xs����?QK����]׼��U��z�Lgu��֭p������L�ѥx��''����ⳗ3Z�	�{��wm��n7�,�_o�aH'��v��~�{k���k��^&*#9O�J�ݷ�ruw�ީ���˔��K�a`��l�夙f�־�Te�Gw9��n�i��7)ӲsE��5�ce�[=�A�X\�+��vcp��B��3��v��l0C��mܫ����I՘��u�p[n�f�*�]
΍i�6����[H���]��9��3���fi�C��y���e�+����kQ�P����4-�,W϶�:f�̕�8�ۄ��«HJ7�î�ivJR�>Ъ�������9�� ���
-o�� ��<ۍq��=�m�.�A+*\���e*��S�nk�sZ ������Mf��Ozێ]z�:����QQ�-��1�=�,�]𘳙��9=+�v�py]@]����R�9�{��*sue���ϹEΞP�}~��FhW�k��ה^�W����sr������<�Tmn���i�]{"�BXbip�S/�nV[+�Lby�]�@�m�*cEv"�5{i�K��W%�
a�t�8l%�)u��_�<1}:φ����f]\�d&�ouN°Dqt��Ü����c<=��X�`%��u��f߹�q�q��
�C%��p�wGG\��ڄ�{�]�ԥ�P!0����S˕
���n#��r���������`�rY�(.ו���2�U���M#�-_O{��aX��\�Ot��Q�d6u.���%k�;�V���+� 3Ւ�s��4V���f�M싷'^�7;y^��x���!��`����E�UDZ�5���q\��h^����[q&%�H�r�����69`
��:�V�Tlf=qW��Y�E��������sX�V˞��/�rʺ.9�3P�f�#7nQϫV�m�G��~��u��C`�g��=:���W�{<c>���S����r犋���g-٘t;=;J˴㞲q�}���㷻p��:�:P��n�pea��*'V��B�&�8�S���c��f8Ui	Fۍ��2����uB�֢�	zTS{�o������+z�<�k�u�*/ ��4���������
+�V�T�/�Ŧ���V����^����:i� ��fn��w�v�=8T{�[pc�k������5Y�en����3��������K�Z�~N1��14��2ֈW<��E8!�Q�tY��v2��g&�Qק/W�Y�V�OfU�g�'��c�V�VjX�J�U�Fm�So �9q��Խz0Х�t.�cwY%q3xC�.��>�o��I�[�@��k�0D�����v��5�Xj_&dgrf�$�o7M r����ɀ��^��:�2�S����p�B�ǂ'Ԙ�J��)���"��lP�|Y��j-{����<�[��oh����	��8T�웉X#i<�UO{w'�yQGG>೰�;�I j1%��*�B�2#[+7-�%_��*	UI����I�Oqyu����N��bgz�bA�W����Ӟ��3J*�;gS�{Ctv?2�)K7=�wWiKv�x��j{Ի���"w�"Fo�������4�v���mL�5ˤ�������\	�)�J��6��G\8�J��p����Yb皌چFv��T����o�r[H�"5Qyo�c�� p+�]�;���r^mOI�<c>�߻#z��~���§
:T���Vo&�[��8k�yw�z5�۞)ס����5�wEH꾕����J�$\����1Q��9J�)嶞�C��p����O'�����k(�i�Íf��ĮV'�kH�
K������y�v��S�e��<΁9������^2�֏,]Im�M��yp��t\��غ��av&/4+�'$	T2�µ�$�kf�W<G�B�fHM�Ȼ4�q%�ٸIYo�'m`^~�l�2���Φ*/�����uڇxq���OcR3����r�&f�}�|}�9��7=Ep��k.1)�x�P;��@Ëz��s��f���~��	�B���=�K�j�}���F#�җ����)�Y�l�m��2�����z���혟6����Ɋ�S�8m�kx�g��s ��k�ͷpZ��U+S��{���yFRC�-`Ĭ�l�&xk���U�7\B���(5{pU�zs�U�ĥUTmG+!�*��[�VS��ɦ�vn���M���b�d��w��W��i�ou���`�����ۼ�~�m�Wt��۝1E֪;�<1N�o��5�=;�o�J�)-��	�B~Lg*��
�uG^�=_g<���R�������uiS���`=o"��x+�n�n!���FG�l�������|��ym'�-ݵFrGuV$�ms3�Î�zɓX<���C:���@�F����BqƯU�+��_ojov�q�ݬȊ��)��j �{�R�.�\zJT78�1�W &�s���w�!7sy��W�F��J�S��(VuE�:)Ó��y2�������<� �_1P�=�O���V.s�Fmy���ðWs�w+���WƳ�G�J�m}��>ߢ�71��C}�����2ߕf�E�&}����O�O{��/*w����KɊ�QQx�Vr��7������+��!@��܍�UϬ�ʳ1�;fi�oW���sq:�e�b�9r+4����bZ^�o�Q\�Unc�ʆ흸��ԅpU���H_9�(��i���H����/r�<��gyU��i���O%�>R�|�BR��7�~|������^c�71KG���F�ΨN�B6���9}��5m+�A�^
e��ӽ��M�8�������;�6Vй{��헙��ke�'��k�mC�v��u��ҵ9�{�m�ԥ��MJ-�a�Nl������u�}��5�W���W1��D�W8��p{�Qަj�!v�.��j;9��Mr��cY��� ǘx����>�7�	�r�o4�EDm�0d��!O;s'_5�ήE.Ltô/�t�kj"�;<P�S6�9r�JhF8r(�����7�w�9�ֶq�����i��
yݰj��Y��SƖ.6�ۛ�I�Lpٕ�%^E����&1<ۂ�@���gQ�p�sW�[΂�@O�1¢e�IW�Y��>����K�n��vV�D�[���qг)Q��y��.� �l���J��`�����{��U���0s�Ew��-�;
Ż��5P;;֤��V�5ʹ�]W�Uޚ� ��ӗ��u��2���N*�k��v3�G׮�n��ź�G^_�\�eu��o��G>��׼���=��+�h��{1y���ԋ���i�ͦFnܫ���x�VZ�s}��1�kNX���w>r8���#k�{�1�(3�9�0k=�uC޾=$8C�6Lh�����ܕ���mV�NOzr��ލx��]�o�`|�d��4%�(Wtڬ�ǝֈ��ڇ�i��S�W����ȇov���#H��q���΀���խ�2x��������TrV�G�}�����Uώ�H��G�/6�}�)ݜF��x����=�	ҹ�Fn�r�Qf����g7؀J��8�"з�g7�����9��]��;J��o�[ka����O��*R��hm���$����i�=�����䅥��Tq[����kZ�έ�'[u� �<;��h\y��u{�:N%f���x�i��Jkqr|�k�\cn�\=� nC9�7��*�ؘ�~���T̊�6d��o��^����/�p������w����t���z�y혟RC��kl�Ɋ�կ(.���P���:�ǽ�5�.��v��J�rS���;)�+��,��*�{��9ZI���s`�)��c�.��s�U��oh���n���c�L�ɪ�+��4�5b�ѻ�-��x]F��J�qI-�*�B�2��'g>\߽�ݸ��3|}��s�Y��;��-a3����P�w���3;$,�딶��L�s�v-_�u
Z�ȗ�U���*�-2g�߱�IQ��;�[�s���ϐ�TBc&�MCX3�mLu�l�T�*w�uR��\�H.�pҍ6�W�i�n�d��M��O�wP��w8ĺS�+`����A��[���8X_L�U��1�����ݐ�+�Zp�t�o$�5�79bU�G���R4��J�V�q��W[S�s�!�����l'C7'�fpH�+rJ��\�N)7��<�g��ס��sV�}Ԟׅ��g�[�T	��:�2�R��*����>��j��ڞ�~�1�(3��1���&��׽Ml����8j�U���{��W��y��^-�U<�������ȋ�q��Y�[7��s�6��M��Ԣ�1z׹J��)��i�dC��vM�����`�[��)��n�[��'ek��vJ�p}:���E�>媣�웦���6"l:�Ѹ$g�q['�W9����o���{+�vJQk=�o�N�cbth�*g�η�R��W���z�:���2�t�l'��ծ��ep�o��e�ݴ��w�Qh��z��k)�O7��5�s�1��
+�[padL��F��9�t�.��7Y����N�'�٪�jsr����T��RC���Z+������m�p��E�s1�1\�neD�B���-W%)�Q��n�]�ak�њD>����Z�p���Ջ��D�\��C�<Mڻ@����E*Q�c�f���0u�)���մii��G�2ڃx�)o=����ኞ�"���|�K����eᮘ�K��G]s(

k2�Jv���hԈX��OP���gE�L[
k�N,�p]�D	S�Ӈ����[v�eMg^u34қ�eT*@O�!�m{qJ]j;�<1N�o��{rm/4ӫu�Rs\,l$�HeÎc�x��þ�D�'��~)ymə��]a Ǯ{�<e���) �4/����c�6�H�©(١��߷���[����eU�	�t��T5�CB�VOBX2i���=FW��iWzK�����c�z����>{�i/e?Q�k����~�r��	Ӵ�d�����i�쏴�lg�~�����D���QW�EFr��7Z����=˶��3�J�n���c�r{�t0f�6���B���J�Z��vvy�y���2Vcu�;�S�J�	����r��n�ۈ{T��pbu1W���t��M�̽�F��i�^e<���Z�#H�p�z<�V��q~�8ׂӲ�s_ml����H
��� ː@1M���@�b# ��*Kj�npMu�wx����$U6�P@�&,�y��Uky�E�},n/E7���=|�����Mkef�<5V�ϝ�@� B�NXf��^2/�w5ܷe`(Pd�@�ǈ-$<r9b�f�Ð�$�H��2mg:�uw�m^vҦƊT;T�;��fP"��ϸQh��;7�X�ti�j�FPڕwm���]�0N�c�b++��L򗗷�An6��$y�)V�s2	6��C��
ƩJ��9�ٷoX��W�a-�z�k|x�C�Y��P���_e�t� Ku����Y%��
n��}�l�&3j�|�λ_[���R��7Z[X#,;��-�"��Iˣo.w-����@�a5-�՚���g+Os"r�7t^F� �s�H��i̡':��ݭ�6� ;v��q7}�nP]H�]��P�N�a��}��.r�>�]I\�k/1��*f�X �`��2�[˷x���̐r�Ũr�珚�xIR�G ����umj��K�5�(W[M���c�.d3ky����Vj�2N��������B���Nݷ�J���R�=�pP.$�o;A��h���PM�����.��e���l�]���1�{+m
�X���WK��b�ءV{f���A�I���H�<5����K9���]�q��ܥ���S��D�Az�
me�vMvm�5g�IR!d��%rㆎ�l�}�)�80��p[{۹�A���w�3��j�q� ���S�{��@[��3�8�f�Y�Fm�K,m�fe��I�4�H��<���?f��ZW4e:Ky��ŵ��姏���1J%4��o���^e(E��W��T��z��R�Z��>=i��q��1�^��<������
Y�Z� �Wn��P	�H����ڮ��y�5)%y��hֻS�n�.�.Y]�oU�C��cLɍq�e��d��T�r����9Ig=l�/��r�E&�l����^�.��G��>ᙝ`�om�qY
��2[b�%�i�ԙ��s#/�|��C-���7��W��3qԮ�`�=�4�\8[����s���]!\]�f��|��;�6L�w��eΩx9y9���*xu�%�b�H���|y��K�ъ[#��fYF�ͧ|�`u�c-q��u�,W
˟���ӂ�rBU6����%�2��Y8uz��/.+v�Y}F���G�y���7�1&��c��0�V�j��mj�dgv���
[C\�`�n�aۘ���_�ΝN|�����Q,k�#��� \-$�%�pt�[�j��3��w��d��!b�L9r�.���� ��ܝ�Q�hT� ��@���L Y��<5T1�;���b�@-;H	���̰��{�z��j�/+�v&m�dd��B�6^��c���&pX�y�]7ܕ�%`���d�K����*Z7�Q�Z�FҬQQ���Qk%kekPDKJ��⢖�-��1lm�-�ڣmUkb�m�m[R%�pV��Xŵ���Ҷ��Z�Lc-�j%)mA�[mlf��e"��R�QQam�Q�Ř�mDf�.j��Z5(�4r�\T���ĵ�-�e(�0R���f�iUj�Z��P�ҕ�\Z�V1#AFQ(��X��m�m-*V�E+h)mKR�mT�,mj6%�iLS�m���l��1������(���e��P��e+Kmr�0�eiiQ-�m�r��mj�iiR��[m���("�R�ʥ-QZR���4*�*)j��J��Ҭm��(��U�kj��V���e�EV�h��c+h��\��D��aXҵ��D�K*��֊g
6�(�*�6��[[V�-��@�
�S,wP�@�R���f�n6�u�>����k�u���r�v�F�Ρ��JɏHS�L;�]Y H�o����7'sՉ!��1�|OOz)�q[׊m����#h��)vn)�+|��ڇ:�v	���L����Ewf�۝��S�~�6�x�]H��=*���}���m�7q���].��������s�d��C�xm9�c"Pl�|���c���h����,��"��>�үq�Y���aЬ��S�i�z�ĽV�G'fRc�zevMĬ��p���`�wl�-�uX�K��ï�	و����9�
@o��S/�n%d�g]e>�I�VrX���Qs:++Jqٵ��A�o�z���Q�uӗ�&�s�n>^ey7�9경�jZR������˩Ew��!��;
ųo&�U=|6�0�\���ys�>�J��"��Q���c�m��Q�G$�Ǵ��gM]K��:V�6����V�_������Ϩѽ��7>��k%�JZ��� ��4s8�^Hٱ�9���3(�+=GE�E�]����M�j��փt��=N��KX���ш�\HkTu�_"to>wN<��;��"����G�=z����U���F�n��G9,KBU��1�"r��gWG3�VgPm��;sL�5��ݸ�sYJ*/=ը����š]��o}��Xc�NKÎ�WE��rN�����d4��)��옣#�z��Ի7Tj��?w9jojUy��U^>l������M߸�s_a�;Q\�o�����8��EE�B��-\��|��!�ݵV��pX��vp�t.��q�~]�S��ܗ�)\���}S���=U�o^(y�֭"��p�/)���6�T�֕��[ss��O�5��JkqTr|����C���uv�oqf�%i�q��Z�XQQ�-�������.wq�^N^�<r� �U���4����)���1��訆Z�
�+���y�9��r^݇����DNs8�YZ�v%>���;���J��0�S��;�5ٕ3����t�5�[��Z��K{^.�����p�/=:��[ĥ�A��q渚�#�{5(�:^bϦ�ܠ�yWgG�nö�㫘�,��Y��AX�ޛg>I���ۛڣC�RKq��o�;7���qT�%C��5�Hk�O���f�j�cS5��;���h�хw]����#�ċ{�1�uA2�vt��a�?Ϩ���O\�L�M�m3��I�<�ĕ�&����:����6���e	��s�e&�Y��0�z���}���� �)�f��t������~��+	پ�ԕ���5�pO�>I��l�Lꇎ�N!�a^�=��Hm3d���S	�߰i��)!�����x&���p�{ӝ�,%g��vB����O'�5~�d��N|�+'ψ��	�$��l͐�����8��VCi��W���a�����{�;�{��\����=�����N �:w��I�'�Xh�pB��&N���$�d��d��N��`�M>�9l+�:L2`x�O)���<5a�6�q�:^�=�u�}��k��_^i���:��T�9�OR|��s�i'Y6���y�=d���y��&Y={��wI2��"�O��
���i�C�3�z������n�}׻޽�|q���|��'~�q���I�>a��a�x�{�N$�+!�sx�I�O_Rl>� ��}�g�����'�L�7dXi���;��s�o=���y��C�|�'sHq��y��u�z�m2u���'�8�?S��I�x{�N�w�	����'Y>}I��"#�{�B�k������RO��wd��p�������ͻ�I�'�v}�H���!��14���	� ��ϸ�q�j��d�T�n�|ì3�8�I8���`�'wa5���'Rz���{����7�t�wL������4G�|�+���ßk0�a	�;�$P��$���q�I�=Ml4��c>�I�V�|���J�2d�S�l���w�|}��5�7�s�3����d�v���@�&�Y5��N�=C��w�d'RsfL!6���8�Rz���|�ә��e�|��$����$�'3�s�{���ޓ��x��R`n�c;7p:��,g
��r�P�ݤR�����;����y:��^���J׌�1��FQ�E��h�hNT8���G����D_���O��BK��`�%NRb7f�Y��8.��6Y��ܗz�n�]L�lr��Q�r��ԖvM��8��~��DD`���	�N�:��&���6�ɯ{�)��<9�d'Y_0u2q��c8�>Jԓ�4��ɖI���s�[�lN�Jϒ�z_�z�������N�CF� q�M���d�)Ԟ�!2���'��=��6���;�&P��:�d�~� �N2z#>�o�}����g)镳{�#ѣ�Dp0�m:b��Nj�y-2|�O�4b���g�m���&9OXq:��}�=C�i'{��8���Y�(Lx���ժz~�7R��6�gf�=G���$��i��M�>P�����,=d��� u'��=1`q��=�l����=a��)��8��9��N��>8���Y�:��5�@��D}���0�$�y�|�������u'̛r�6�M!ְ�a�(|��d3���m��u!�=|���[;�L��_}�C�j��D��=� y3�Y/��RN0�癒�I3߱ԕ����8'Y>d�ˣ6�L�T<v�q���u%}d2j��L0ߞ�f������ed��"�E��>?I�&�X;�T:ɴxw�!Rm�!��'���4^k2T�'|>���}�ù�:��M���Bq��x�]����}�'b���+m������т0Hw��C�a�C;��,��7�2u���b�Rm��*M�g��OL�w�ĕ�$�͒�o������o���b�?*�[(����z0z#Dt�=g�N��T6�i��k�$��PY%MoX>d�T'����N����T�d�cԓ(9���	�m�ITJf�w��m���<���{�B�:�N٩�C�&|����<Շ�<d���I�:�}��RM3!��q��P�ݚI�M���>dCޚ���Z��#��Zj��H����/�a5��&�6f=e0�R��[�z��Mg�y`��tA~꺴��m<y:ed:��û���Y�.�����W_j1��M;[�{c�>�w��J�ڹ����y�! h��ݝ����S��fE���d����#�8�眞�����ӑ_���e�W�����L���$Rm����bi�����M���<d�'��m�q��	�N!�:�d�3^�Y:�	�}�ߍ����v1�3~��p�����{�|�z��]��I������&S��,=O��x�i�	�� �L��N �y�&�q'YSɺ�a���#��MO�BI�p���!�������l&�;���d��'|�ui6�9�I��{��Y�'�jw�a�x����I�<���I����'R�.��|���ܴ�x��oY���������'fr�}I8���18���Mo� u&�Y5��N�=a�y��q!˜�&���q"�C�O�]��N!�cyt�������D�w�;�}�^��b�x��z���R|�����d��S��N0�}�N$�����@�M��h����m��wY��C�cY3�D�_}j�B�,�Q�V�r������>N��M��xf���$��8��T���'̝�2d��o�'<�0u'��&����q>d��q{Ѣ!U�ٜ�+,
_o�r��Y�*
\�HVO�Xt���I�5��q&�>X|�a8�1C��:d<�8��'����@��v��q����C�Dz��ESA���>UܗI����A�&�;��
I�2k�d�	��1>B�z�����$�OY��I8�i�,>jI�d��ԝv�x�`|�O�T�!�}}�Gs�1������p���L�w<��8�!2�g�!��d�<�,��=9��L1By�u�d�+'�9�I�&�Mf�q�i�VjI�x��=�<�>��6���w�h�z$���LY6�ix�,'P=��C��,�=ćP��Ɏ��XN���2T�&C�c�+'�Y1�'Y>d�i������)�{`9�d��d�VG�R���U��[�#�h-I��<���w�e��;̨�]\����mv=d7Lo^Kb��o%��h4��]i�w�7��O+�w�d���T�w�u�APF����v��M�X��k��ۺ���7w;�ju��meݤ{�������(�����!��8��'z��CH{�~��'Rs��C��Ag��ćXz��8�I:�e�%J�u��Vy�2~ɬG�`}��X����3��l�d�4��3��<v�|����ġ��Hz�	�ݓ�%q��<I����b2m+s*M��{���{���8pjD�z��o��hn���zm��1%I�Hs8�`|�N�Y�:��g�<z�q��VCl��W��S�0��i�IS�`�'X�>�0�{� �G_���ٺ!�&�f�!�)mW���'~��,��%t�u��ĊM>�<�0��M;ML�d4�<������6�8����hu�g��	�<��߽��p�w���[��J�s�4�l�Jçy��z������&<��y'�L�ydRi����0�����f��!���g�8���j��">�_�4�d}Sl}{Һ��l���L6�yN�)&����z�Ĭ�7N2u�n�s�l�d����	=@����8I2�C�Ċ3��<Hm�����!�}�4M�ߴ�k}���k��P�'�(ݓ�>d�Vy��C3�q�I4���`�'_XM�@�O�Rw�'XI��y��m����0��	�5�q""��D<�?F��P���럫wTU��g&��:f��RL���'�yR|Ì�J�&�O�u�g=�N0�ӌ�t�z�>@�O_�l;�I�Dp�p�yQcރ�]�}_JaU]���6�}�M����E��O�G3�)'��C��~Xq��X�'�8�Ĭ�Ր�'����8���`�O_�M�bRm�'���z�vqs�u����u�o�ߥ�0<a����O�\�:�$�O��C��&��RN0�0���I�Xq���'Y>t�wd8=�=c�Ǽ�{;#����!Sp�}�-��N]x(m���"��J�-w��ƣ��۶@�|�|��7\6���r���f��r�[($����Kٽ�/�����r���Y����U�$���T��v�q��i[�����6��Vd���Hr�Sj��qtF8����3�z�)��?E��#����O�����^�Ra�y��!8�y�bu
��)<�c8�=M��>I�ϔ>fRO���O�- |������8�Gr�k���)���A������ē�<�q=a��.��@�3L���d4�C��2a	��bq
���w�8��k�q&�>X}l��޻�`	��V[W��%�!�X���LF�>I��kXa�}v����y��M0�u3�@�3L��w�RN!��T&��:��|��ɜ�0��D�=�ԁϜ��f5�.�G��p��G���d�3>P�J��ݝ`q&�P�Ł��z'P�`}�m3ĝAgs���^� ��0���$��#���/�h�����p4�gf��<G���}Y�8��&ܦO�4�Xn�N��I]�6�C�{@�Cl=>�P�`o��*I�y�`'��p6�@��C㛹/�[�&��=�!������9�q%d�y��$��h͐�i�T<v�qXm�z�ίC����S	���)"�<��	�>��k�c��/�A{�ŝ9�HVd��5��IԚ%�%ՒwG�VO� w�@�M;OL��=L�(x�	Ğ��O�j�!�"G�D}����Mf,�]ӽ��~􈀒T��pu�h)wi:��V;��6ə�u�ē,��%Ւu���)4���s�`|�N�A�!����#��#������+��@nK�p�L�M����C�:{O�RJ����:��xs��I�OR���`Y=d�k?2L�xs��K�I��������g�G�4D!�E�߶>��ޮ�/�!�Cl�i��	Ğ�m���T�H|�3��e�i�Ow�Ĝed<�7���d��&��p�$�}�g���ث�W�1I����`�S�i�*�*n���e����7V�})\V�vub����&��P���+��V����J!dac�zY����"q���iV�K�ȬP��*b�V:�����ь�=���8Q�/�r' ��9��.�N�Ϋ����ĳ�R[�MFcof�Ɵ>Ze��E�����i!�8�&�Hu��d�}��,�@�d�L'�8���0�<g'���'}����d�'��r}�"#�{�+����G�pT�u���g^rl�wY'\!=C��>L�9l�!�f���
I�hu��(���':�<݄��Xg�q2�q��3{�i�z�_и*������b��=�$۶N�u�>`z��G��	����a	�=;�$P��$����2�8����i$�}�8���5a�N2q*^z������w$��ں��BA�$��֜dެ'w�(I��M{�:���]�Y	ԇ.q&�C�RC)=gqp�>Ci�6L�O�YG�����f�AȚyY�`��h��O=}g��8�|���d�}�I��^��}d׽�����s��N�Ʋu2q���q2|�����[���Ȋ��v7�N9��b$��Xz������:��Hh�!�!��m���'�����	��{�!��'��RC�|w�fL �2��A� zUɳ�����rn���y�ϝi>d�:`�OXm��P�2�u<Ň��Ր���'�4��F,0:�O������=a��)���|���d��y��?lnvED�;'o3ϖ�y�0�����
��T��8�8��Q��&��(|�I�����M��yl�Ri�����!Bu�S��b,Dz�ڎ���|H��w4�U�V.�t'�x��� �O��}�fL%I2y�8������q'̚r����T:��3<��J��8��=a�I���z0Dp�
��b�+�5Ծ)n�g����L�t�؝L!�'�,�hN��'�;�b�u���J�$�~�RVO�`h�8'Y>d�ˣ6�Lɪ;a8��j�RW�C�������߻w�] ��m�9�=@���w��Ƞ;�s_^ƾ}-�-�sMl{��3�놠v����x�O���YEG9z5��^=5�t{eD6�ҳ���C(��V�rD*�`6���t���wS��b�����=�����^��;����}��d<C	���$:��2q��9�T:ɴxw�!Rm�'{��2N�Լ�d�RN�\IY>Ձ�s�u��}M����}���S��|��_G߮u��q�}�ކ_�O�|��4�27~d=C���Y%L�Y:���,+��*��!Rm�'{��0�d��׼F�{�g��x�{��#nb�U�1/g����>�9�o��v�6�Ι�`i3�6�!>I����x��i&��i8��*{�`���P��IԛeC��`�I�L��Y�$�<�ݚ��p�^��|˽�����v{�H���-�`m����4�L�M��'�<ՇS�<d���M��=gX��3A��q��P��&�u��i=�{�u���7ۖ-n�o�{E�"��c��>y_��DE���$��	���1"�o��<d6���zf��Ci�)�x��O&��C��A|7B|��g�:�d�f���g�2�����eFo%G��${�AL�	=d��;�b�������$��;��'�L��7���9�M2C�a4f��Y&3���Ad�VM��N��.��O�&��ߐ�گ�=�=���S,'Xy�`����M�2u��l��'P=I��5�M�<�u��0���H��2�����I�<9CH,�߶QQ��(T�ܿD�Q�������WM�u'u�<�	�N0��8��q���$�������&��u��^g�Bq!�1�C��hh;�H�P�B>�aљ�O�]��\���!�z�B�1I:�yC��J�ɪO�q����vC��a��u�!Ϟ{����o��׹��uB�������%Zӛ%CEwY/=�+�Ůy~Ħ+5TJ{��r��%简���5�m��J��M�nAc$�f��z������\�ɨf�|��Ҡ�6�� ז�����;h���x�bc��fi�]�l횊�V�7��HD�U�y; �di��5(�B'AՁ�ܹ�^�9g�b���`-�oV��\�w��UU�+��bb��J�L$���م�](>��]�x��f��^�!;�.NU;t�۾z�Ľwi�t"ip�^�)m�Y5�LV���\l�/�+�v�f�¨ )��+UNĦ����Rxb}I�2�$���=P�H�K��o���\����ځ+y�qޖ���u�����aI��<�[PN�|�5�V���u�V����5�ׇR��A�T6����qX�t��|Ϋz8�Ʒ�=�!�^�){W01u��R_�gw�E�.չoyt�.n�z	��l|��<��;��ZzkT��98���!0�w\����g�!R�4�J�٨k;
/j<��ˉW1Y]Qo)F[(F�<�"j�mh�m̜DF?sz)�-��C��[�e���-6;Wڷ����%��8��/���	�9�nbM��Aby��'}�������i~�<�B'��p���r�m�XW�e�Jh�E�6�l��;��
ٰr�yv��M��f־��s�ŝ;�ecox�љ}]-���]�#�ŝN�%57��l�퉝�����*�) �0��l'S�Ӳ[8�̛��&��u�+w��6iGe�ݝ�w+`r%�t��$���D|8 �@_+���(�7v�E�L�89(Gڵ��OA]7��V҃/n֍�ZjG����)�6t]t�=kv�Tmq9o�k8�]#\�-Xk�ѮZ�Ħ
x	{7A�p&���'�ˠ�e�㹏Qt)K��\�	���j����`��YO;��]G�: �Ѭ�]�K���e�T��^Z
�M�F�U�s���;���>����%iL�8�&�}%R����W~Y���Hޫ����s�� b�z�9��xFd��RV��+P�Y�%<�ze��ԱM����u7Z�(bc	�W؎L��9}�`�ڴ�=�K����U=��O2U�}��.9c�
�;(.��q��-0��L۶Qj�mX����z�eH����Z2�,�ZvAI�
�{�fm>��%��j�a�/�/��H���a俴���f��z��;�j���֝l��ٗ�8�z�p��QK��p�t���S*��v���z�jY��Bħt�si�[��nY����L���EEY�}x塔��&�NJ�;�X���ē
ȧ��݈�G�>��䵪�\)��d�Z��[���v,[%����]v�1�j�²�y�5��*ѼM�`�PwP3rZ:tw��ejv������%X����}�J���;�2�E>9���YF���@)��* ��#��$�����y 5��,�PZ�6��b<I�ۼ~6"�Y���d���1�å��.Cq�7v륻<�X���7�y������r����-:s:��v]�fWVS^En�z�ZK�%�4>�V�-�V�A1x��,.�{�2l�26���4(�Qw'��u�u�i��
=�N�9�b�
`�Xc1처��eERvu�w�ً�J��gPu��ءbT�d����w5-��a��r�5����e<��>vM��J�X̴(�4�]����e֥J뮡��]�WRw7�@�.�F���r��w�4�s�V�E�\�WvY��3��h6.�z��:���m�:n-<�ܙ�oosE��l:�*����5F���F�-$�ۤ�7}J���<0��3>#�]��:��Ƒ���m1�k�wL�;��h֗m&��fP����V$)�{#�L@���q�r�H����Cj啈��`P�2�e�t�i�|�^n����R���7>vf�z�]���[}}��͜�����5֙���C�M�>�+;[���4���s�m�y��vl�{5�)��(�M�,GSe�9V&c_Gn?.�<����\6/�X���_�9;��r�������ή��vGg@���ke�����j���)���Q�+ij�)iJ5j%��KPk-�ETJ�U�ь�Z�(�����(Ҭ�KF"��m�lJ��+)lU`�VX�����m`�(�b����Ԩ������+ib
TK#T�2֢��-���kF�)Q��ֵ�V��
���-Th�k1j(4VVP�b��ƴb�Ս
ԭ��l**"ƉQ�KYeh�Yh�������-�آ��kl����ֶ��Ԣ4�5(�klmXT��JeA[e���bTX�eTe�cF�X�[h��V��Z�hR�V�-�IKV��K#q��-ij�֭lQŢ�	Q����*%��F%��,[j6��b�\VZ*""�mQR�
Ԩ[J�+Z4DEAF�iU+UJ�TD-(��AF�*Q�DEFR����mK�EVEV*X��QQETTdkUDV0QR���Q��Lb��Z"�J�ʊ+kl����+RѲ��j�1cS*���ZՕ��X�[eaZ����Mh}F�g1���x;G@���[p�S��z>(��Uv̱�s���(s�}+��,�����u�˽�]x�o׮�M������GO�����Α��`
����r���jv���0���ˋ�(�>�ӷSxmz.���9���;�15���&g"� Mt�@��R�7(D�rڅ����^��a���&�>F4�Ҟb�.o���B)�oFB>�=~U5s�Y�Z�Mb��a�)�q[\P�2����L��4��,��xjsVa��F�%����U�G<N��m0Í�gZ"]������4�7�q<�ds�5�yLX=#V�F+�2Hó�N����8�����=�t���L\S����Vq��-�T����/Ć��<�Bo/��7#6��(<�!�i�Ny���sf�ȨW�l���Nw�k�|-溶�8}���s�X�׮`1S���͛�(f�u�R�K,C�uE
��W��We��ǇwI0�_
Dߪ�!��Lm{'IB��8�Ib��xuXA f�9n��r�Z�i�3\�n4[�T!��.B��{M�pw1�K�E*��$���=��VQ����y�5j�κ,�Kֹ�Y<��"��:�z<{�^�L}�/Ȣ�]b���k_{#p�.'�(���b�;Y��뫠�mfE�ܗM�otЫpl[G���S�uxG��\^��H�i͙[�F%� �r5�E(J%Nlӕ����o�������>�΢�]�IP?y�;�s�3a͊YR,ÿq�ا���Քφ��'���{2VR�mZh�}<�P��%���1˭@����{�=��/��X��9����3��.�4��X���oI�zw�n�����:"cTL�L�Ju�'Ӣ��:�Z硍�,(���W��^�;u����j�\d�F	�"�7) an:�=��w��Zus�j%%�+T=��[kc:���q��)M�U5��'�x��4��:��Ρ釪^��:�����ج-�}S��u6V��Ü|��(�����:Pf����R�]'q�����Uyz� ���n���yLwg��]`�OY� ֶW4�JR�����C�QjVFsSǏ;r�C7�d`~MS]-9�}�q�˫�9ͻ����ט:٭̺�EMC�y��>��Fb��|^��[�b�c����D\k�����ؿ)�rb2�F�����AV���%=����{�S�ǢU�i�S�'�.�f�+�T�Mf9\���s~��}ۼ�t$qz��a۩O:<i��9�e�@u�;qb�}>-M�tr�m
`&���ޓ�bi�8_:�;*��Z���y]��;���v�^*�՗wgl'�������7]��s<������V諢gok�ԷKN]s��錒�f0"��諭����'{Y6J���p쉉cj.U~��+�OYܙAנ�B��<�ȧJȾ|���V�U��51�r�0"i!\M���,f���E�g״e����%_������8�I���Ύ\�?��
�@��泠�pE7[e�|���X�;�Z頍���έ���T��Xq�Xc�]�YV(��|+lϛ^�[<1�̕�g:���{w�ӻ���׫<��N�5}�k~�+�����+(��"�m�zc�����&'�<�^SV�!.����c��9�5%�&�:i���
ɲƋ�edt��y���[�N����X"�o�	W����u��9k�~�~v{�0F#�P�q�W���דyL%�~��p�>B�AX���gC�{Vf·Q΀�Q�ݑ�7M^�V����g5�J�**�GF�mBsME8n���f3d�Ȭ�P=��茞x�"�˫qzғ�Í8��X�U83
���5h�S��ɱ��쉉��P�[�u>d)�z�N�ۖ�3�W�;������'�u:�#K*�)�;�,m6*��p����"�����}³'6�+36�4]�4�t"�l"��R��hJ�y6��ݝx-�q�UcV���"����,*�M���B_;w°s�����ܝ߾������i�(���Vv?D���5T��6]=9�Pc�!��Uw���;���#b�� c)xE�rV-}J�=�.< vx4��k��U�Sӑ�%�㌱�n�!^ST����:3y{ux���*xLC�L����Ur�#�gc

����Y!oL].�󘾞��ˡ�E�=����-�~x���f8��L�{$�u.�.Q8ʺ.�u�X�;��[C��.ϝ8��3O����� o\j�0"��!@�R9�10����.V�y,x�S�8sS�Os/43��X&�
�u��A`&݊�u3-�10��c����W�����4dgR�*-hj��ن*V��R��aC��B�$	�'G��So�Z3�\.-�3\V��]��R�t�֞zr%�g\
�+ܦ������`:�NDd�&��oj�V;���Ԧ��E"`��ŌuT����C���nH��Pܽ%�T<#%텧��������I��ȕ����2�0��R�X�b�Wة���*���|pYn�[:�'5FuT\E�ti۫Vi��U�cVN3X�&�J+,:{�s��	j�9�y6���Aλs�.D1�,=0��S:9u��4�5%]4y��6˭���#���.�Bm�E�g��_^Q�|�GXtP :ee�Y�ˁ}n~�磌�s
l�_s�DW��\(W&�>DJ�q����L`�'+�~+��1�<�q��KX�A<��n�p8�,n��+*(?5�n"/��G^b-����E@��D�]�p�事s�}5��v��ÁbVm"n�1�F��	/*EsT7����1V�Z,���Q��?5��y�U�G!�{&-s1y㈢ib�;�����|c��YC��בX�������J*�K�����!�x*�SQ����Bg��s�z���`=����Z�S���Ѣ4>q.͹�H�z� Mt�@�R�:P�Y1�<�q�S�1��k��)hHٚ�ϼu�˖�i.��r�3������u�m�r�.�xx�l:�Ђ�����Nk:fj�4�V��s�9�՘aF��#�ȅ�jf;=*���R��]����*e��xˋDa��b�9�F�5��=��G]� �Q�PB���8��~�N�,L9��y� z{/K�w�Ñ�X�ަ.�W�炲���6�*`U�EpHai���"�+r�+bp�v�����q��z߱:{Mwoy��xu��ƫZWVb�ʏ]6�u]��G#2�T:�i��8s�8��U���	���X�mv�:�ͫ��U�͂��Y̺�R�t׊��rݼ�F.sW�.��u�2�0��I߾�����#��1�">��1�9\�(vl�IA��c��<��:ͧ�P�^فѰi��ձۗ���^�e�ĥ�E@r��&à�͛��m�P�ƫ�Yb$���.pv����n�����$�[B�7T���3rt�*�8�Ib����Q���d�����C�j9Q�!���1qX��Zr$�z�XB�%��DR6&JY�h�W;�u2�xg����P���\5DmG�ؠ��R,��O\�Kzv"�u��5�kz�0�S:�M��7����|I��3���m�#�܌xAP{�J����n��^�U�/�t�[:*�-ڄ���r�f�1���S<|��~����C��`Ce�)R�����
�m[��"9"[;���2�jü���ao�ȋܔ��[����r��goW7=���e����=�lV}��Q��k��J�^�%P�P��P���̲�[��P����-�/8�m��j���w�\ܝ�~`��`D�=�(3~�A�\$�B���Ȗ
�:�]�.����1]06�pިo%93Z�Ѝ+q�����L��.W������q��ۣ�2r�\�';�,H�9�7j��2Zh�8��"O�o5IR�K��-�g�=�&K�J�st]�H-Y�&,��������V�D>	���.�j^P��uw6�n;��=p�j���LLE��3�*��w�5��L�.6�a��s�\F��fߛ�5��w��Ûw#r9��@�(m'�I��
�+�^�ZRn&w���V��[�b�c��q<4E��֞[�8�C�9����4/�m\��m�i$ص��%[3�}j�p�N��]*|��y��sz�}Î3�u2B�龼����S�T�.�쉉cl�/}3�,QS�t��U-O"��8���ٲ�K�z��[��,��t�����HW~u-Ș�6�%��z�^ٔ/z'!�#��39
�v��8qM(���"� �\�oy�#�m���-5ı^�'Nkb��i�sO�Q������¿
�+y�� ��TK����Q���U,v��C"��=�9��Ք�ʔ�3�㧊�F6fv5϶:e@Ȅ���m�!��ⲉ.��a�nD�Z���sٚ�4qR����+���1z�g\9�Uz��mI�����p��ʞ=em�����rm��eܽ�==��+��W��C�Y\w@2�+6����|O���5N�F�u7�n��8%�:f<�gW6[.P|����O���j�͝y8�)v�GD�E�+��	 �P�œG��&��y���6jk'4:-3-��U�U}TJ,.���/����������Ko�v�\b��P}�H\�ɸ����Js䧵Xh�x�*��:hA�/��+��[:�8:��X<��.��g5��h��xK�an�q��D8���t�BSï�,��x�U�C5Pf�'������W��w}g�y�s�LM�YM4E���I�����x��j��¯y��\i�=��}����U�1�I��g�e��I��L�靊���O��UHir�����ǖǵMU���܎�>���ٚ�����1���s�S��[W�`�y@LWJ U�	���L*�ON�,f��XѶ��s�M��vӺ݇�*�T�Y�w�N�Մ��7 %-1Vl �[ۅpH[��%�JrU������8�)��1�v�U��a��_L�{$�qR�r�����g_iZ�GG�/{nˀ�<ϻ�3K��p9��k�7�ݘ��
GL�t���=%�Ye��AU��	˩]�Ψ�dy��b��+"�r9�X	�b���@B�L,7�T�e�Y��,��v)�{a�E�Ao��8��C5#E�`��m۷[ͻ*��L�ͥ��	�i����rMp���	�&(�A�v���v��}ĥV��te�k�O�<1�p������d5���FVA�/U1�c�[˘�k�����TG��7�v�`�������+ݳ���Ҧ��u�H_��@�N�3=tp4���k<��1��t��yOD=X[�Y��LW)�e�S�zn]�1p|t �'�KAr�	Z�g��yrl�|�>�Z-�X���\qS���}��6»p.�# Sr���kIZﱮ�iJ�[�&����IB܉Xn K<6���R�]�]�|���> ,��Q�|��v����u��!`��rFW�e\<(ᆀ*ːx^L�a����X���!�zݞ�u��,�Ountא|���p-%�"5���kF�<���R��ז��\��ޠ�\����˝����c�@�&72n�1�"F�ڴ �/"{��S�$Fn� ���QG���u=�vƸ{v�`���F�����Q4�S�|����}:�e���Yˮ�խ�_�r�3�R��)�E�N� �<G)�����	���N��;���óv�-ꬥ��#�;G��q�9k���)l�(F�ڎ0gy��~�F����*R���̧jou��N�3������U:�[ɜ)Nr7��Ӿ;�F�n���r��L⨒��V�U�����wh�[�	��[�L@���vm*a,u��B��m� �Z�G�}ڻ���+\���p�C��*Q�i![�����U���U6��~��^I���r����N��3�֪j碫 p�RɯF)a���^�`��Ӏ�[��wW���c�R�������cY�0��]��P��2#�5�v���v^$Mc���q�y���27^�W�����9�q<�g���Ƽ�.d�*8�_���kn� ]��kr��ߎ�"ы�ӵ�l��ì��������&��k��neL
�oG���E$�l֟wuŮ���=0tEp0�Ƭ�%͜�(:�޶.��ɡ,�QN�c��ڝ��6�3-s�̓�c#I��ᖩxd4#���P���)3a�=�1����TNQ��yθ�ČX+�yӭ��p�Sx.'~oφ;o��:J a�S�]��3keԄ
�6�wP�q=]�;"W*�sb�O�@zz󐕃�&�z��/}i�u'z���)��Q��X�}X�
ʀ�/֨��9�A���x�웇R�ޝ�,w�������԰���=�O�Wě�4g���ఱ��#EC컡l���t�q�W>��@|Iy���œ�Q��Z�/�%v�t��_|Ȑ��@Z��P�3�x��A�sGӭ�Q�S�� �Y`���V��m��٪���+���x�lsku�Y*���]�D�ޛ[#�ƮJ�c��7������bv�јi�&���v�Ŋ}�1|�	}�1��f��fj�]���t*��j>���/H�v�$*<������}%�G��l�+�I뭒E����B�k�S;Ѝ}]�6>Y���>Z�y�w`�[���M�����W�Lj�9����.��^c�k�NЋ&^i"�X��mnJΥĸ[���t����j�WDy��O������M�T�5�ⷰK������;%�%\H忦e�ò���]Ƃkp=Ó��@�<�9�8���Nn��ǐluf�L뵍\��]�����՜"ۺ.�e�좴����5�ls{|���p㄄ݎWJ�vڤ0��7R6��YַHd���x�Jep��ٻ����RJk"(2Z���J����^_+����ev8��,�EWJ���cx��ܰ�ץ��t��%m]ep��xD/��l�k���Zv�RT��c,Wq�����%k����*lWgoP��wR���ΉK9�Ѧy8�[�}��9�ޣX:���Ы$���G��ͨB�-�]9ki��+vu�����AHt�(3��q�Z�f�Y���^ٽ���n�\�q+Yy�-$�O�Y�M�����N�M!d�@���mp��%�D�ʴK��DQ���5��#'�q(�3�J�}��.�6!d̽����7�{��Qo���ys�k��/X��/:�M�K�^�96N��� ��@ʸ{�T�=v�r�4r�Ȑw݀q�NT�ԁ��>ݷŎ��]r��Y�->:#�����㥵�]PN{ը�PK����:�h���𻺾V£յ/PUܒg+t�܆�hW���hb�7��[�"Q(�_[��Ϻ=�j��dJ�#�gS���+�M�t�vuyp�2�%�����yb΁�1W,��%�pR�C^`$�N�I[o���1rhb)�;\:�����U�k#l�s.͑p��7Oz��e4���)�2��\��)�N��\C��h�e�_inə�$.��V
P�)Ԛ������o� 7���u^R\O�U��-l�X*}jn.���^�Wk���G���P���id݋#&R���1-l�`��;N�4�錼E��Η�uh;۰��J+�1�{��c7x\u���n5L�q���DpGϲ�v��&�M!o�$w�����Ę��l��x�C�?z�ޓ����x,��z��e�fΚ�	��,�Yf��X[C&�h�0�W��3�	��6y�@�t	Ge\�Q�,���Ts��S�W`�r�CJ�;4j��Œ:�M�֍��+a=�R����wm�ն���	�z�S�m­�.�i�2WJ�� �]m����:�+����v��u}��z�h�ʈ��#Ymh��F�*V`2Ь�R!mV* ��DEJ�`����1URT��VU��*�1Q��ѣ+-���ű�b���"��D��V*�Ub�`�)E"���XT���DE��QjT��!im���(��
��0�*(�F����F!Z�UX,�ڪT�U�T��Х�0EQ���mPmR���VQ�"��%�mZ�A��EV��Rڌ��R�h��a�"�(�`�U+
��[%AEVE�
"��T�UPF5�V�J5EdD1h"�*�V�E�
Ȉ�
�(����@D��iid�*�R(���F�**1JʠԨ�#i-��Ŋ*���mQ�*,*T�"�#*6���A���@����S�Q�P(*�,�Em�"1PUJ���� �������KF�Ѷ�e�*�Ţ�kDe�J�KmAAE����X�"ԲШ��m�U��U%�JŭV�m��",�(�1��1HV�6���`,L0�����kc�Yxv��-=�d.vXj��G>Y�H�w[�j.���ځnԝ��Wf��t��ĳ$�w��#D���'Dqi�2.������T���V����E���p�2wn\Ӣ5��{j�7�Ju�&�������r�9����S��n��?t�c/�A^��k��Lv}k�%Z�Ϋ�
����k��[���9��	�ٞ8�8}�<pOn=E�e�0X�*��o��a@��l���A�'T2vGN��'Ӝ���\�5ĘZa��wN���ݞM��~�`�g�\9���:�5t1�z�Ғ�<h��m�.�hD]��� �:5E�R�0\6���yLwc��Н�Q�pky\+)JT|y�*���ך�q�
/�t�.0�Y�a�����.������e;�b�۹��EM%j�^@���C�u��dC��Lr*̈́�����,r7�q<4E�\N�'��B�甶یR���T��r�(|W�$�2|��Ғ���[�V+�'�p�K�4���s;�x�'c�U���bb�Oܮ�BR�P-K�8�c(�,�A=grePsL!{Tq��=��]�ȧ�NC9y�A���&�Դ{=1,m\�X�����m�\b"��>s�",��	��1Ӟ��P��JA�/_I\�qB�+K4T��j*��9{�&�V��V^�Yd��M�v8���Sw��}}�L�v&aϭg\*�_tb�T�m�b�:��F��u�n����L��R�O��*CG�s.<���G�#�Kl-k���{�	C�@Z��J|�H�@4W2_�y�6�N;���.��B�7-�m�|�~�����>�h�xXؒ�Do3Vވ�vU�"���n�X��`����μ���=n���W�J�k�S�*ē�/��o�ZRYظn��P԰�%�ɳ� '��[٬kmaAaܩ�w���vfTk��1��������NW�.��c��F������o��|0��*����\�~%^c���9��+r�K�˝���}+���`���}������,WP�s�+��[:4�龥O��1W>��+�-�o�^DH'�E�ڍӍ��x�$\>�7NW��j��W�R|>N��(�*����S��U��B���x6T�d�����u�t�'����n)�Rɱ�3+Z��T;��*��/$�;�P*,�<n"}�ϹU!{.��e;r[�TJ�^��˚����֣ɳ�2���$QA��0o�(	��`
��	xy��ZaWONF��7�2ƍbF�Fs�J�<�u9�h�ju!z�s-g�8�
��ٮ�er�4�"D�͢�F� �<�Ɇ�EMɆ#�ZrQ��K�@e���ɸ�ͥk���;]󱳪Q���Y����H*=��X��V+����et���(��gw��� �j^h؄|DŮ���W�_V�g�-5wP�Ц������,�SLt܀���!�*�2����u�D��T�n������g�)�Ws�gE
f*ƥ�v�\25�xE�Ļ��W-p�񩱔j��>PZnH��4�08�u�3�^a���WL�w"bam]u*�)\�g�!��}S��:�`�KZ=O�[��̂�L[�@Z� !�:η0��0��p�P��-u-6T���e��0�J�Xk)Sg��C��@����X��mo���z�a��u0|l���s�f�Kzr%�g_�S�aYq�N�鸗qL_�v�e�5V��M�X̄�Ua#�m��J|���,m�Igf1�=X޸
������lr4��evx�5�ǟq�f�LA�ﳉ5��O	\��0/�7 VxX�>�l���	��Wf��#���D؝ TBrFW�ʸy�(ᇈ�X\����?�U��W�;��\5[i���sͨ
�-K�D��V�I�5DD����mhۇ�HΛs$,�,E�UC�-�v]i�X����������3u�}�}�_��n��W�Q*���6�*�Τ�9uĘ�S��E���YB�g��͌���B���ݩK�be�[��g�ƶ�w8jgBw�˖�N�΂�邇Zz �������&	�v[3v�*�;�Y֬�;�W��}�VD�g����'����ie(6����T�[�ƞ�Q�EC��"��܊jFt��Ī>�ُr�n�<el�!oK�2�n�!�dţZ�,�(�����*�tt@wӢNaA��u���$�o���:X̬%z��x�O+y�]5��&�GC v
���e�v��@Й�""zDj_&8����g�]��ܺvi�&d�^մ;�ك�>�8��,�hhɉ�����S*�MJɎJsKƜ�+>�8�������uؔ��'/��r�뻊'�T�=a�EH�
c��R��f���9�y5f�6��2�t�B�q����F'�nO_T���v��/�g���a�������9���{���F�� 2Q�PCoe�=����.[�z_Tt� ��u�T����8�����>�7��=�'Q�yF7�:DM�t��U�{%<��pH��n&5�aэy4J��J�ϭ�g��	f6��Lv=*593	��ڝu􊊌im�;�Loφ>�P�k	��^(��C�&]r��{��[�ԩlh�K- X)	B3��gE$�k���u��I�^R�V�M,���@�^h����YB�|�~"5:�t�Iү2�˥}����S��m۶'e�5��Qv-9��A�uw&΄�&���g��:�wB�`�\�G�򾯫ﾫ��fy���\W)�z��LLswD��_1H��o�;o��'��U_+G½p4T��sr�os
��]
hh���a�S"�*�����R�RZ;S,`Q��� �{�i7=�f�l��"9Bf�+�I�e��HK�/�Q�	aR,þ2{&�KzI|�����E����\Ӳ����xwnoاĜp`�g;p.�ƛ�j��O��"Ö��&2�m���]rbNmu�pw���h����X��U��wO�(�x�ݏ� ��Ӣ�c:y�cY����7u�G-���UW��7���n�c�����gޙ{��1qT5�*K��=�^�t�Q2���$��~�{0m󠮝xV�3����
�6[#JP����b��<M	���p�Gi����t�C��݉�G4��ظ��U(Q�g�P����ٛ�e�Ů�Gla}\9tX��u-�OOlC�c�!�dhN٨ރ�uO]sN�R��� ��y�<��9[\;OQg�F�a>�s�^��f�Lc)��Y��|rߴ)Y�K29N��F�R6�x�I��P���,{�� ���f������!��u~�M	���6QP�b��ĤV:�J�����j�'}�.��1ܮ{]ۙwͶi<��J���nʺR5Ŋ��2`��9�kQpM��_UUWډ}�:�r^����,m�ȅ^�|xG2���z�����<0Gk��ՉD�o��ɰ�9�fb�9�!FB2�G#�2��R�
�c��AS�'�.�͸W�T�M
/2��	deV�^��5�.���x��
nY*Lq��l\�.�&xE��Q݉�ȊO�G
��뉦-�:�&0O.ۊt�KCڃ&)!\Méh�Dı���|՘qa^�ى���:�n���?��E`�(-vr��|�H�@4W2er��ߪ�q�ʨZiڴ��q���U*R�����<_��F���*P��jÌ,1�� �AV(��X����վg����,a7�;{�,�+8L�쭙��>�T�ZRYؿ7Dh�u,�~(o�ݝ�C<��`�F�	q����]>���S��ԓ��*+��^���x �+C�|tƽ7��H��#�l�=����s�s�\"�oÄ��p_� o'��*ـ�{y�z���������u�\7�tа�f��
ł8;�5l���WT�h"��W@��?^�c3H��5qWpmZ�1͚ǰ�l*��F�Nޕu�bY0.�^�ݙw�.��>aӷ��)k7�q{hޕf���Vi�//[�N��Ws\V���:��aa���㤶��|E�sWa�Ƥ�4��i\WmAӝ�
M���9fd�v�W/�=�\�r�v��Bt
���{��<���x�$>�5�n�����e\t9+f�X8��N���̀�$\VO^�tp\qa�Q1��F�O'C��QK�hr���l��!)�vu4�򮫴L�Ș�SE�E���#1ʩ��t��(1۞��Ƕ�]ਜ਼\�=V20����)k���5�͆nP;(	�� ��<�3Qi�Q�SӮ��v��[�1����7��
p���3.M��p��re��Ee ��H،S[ۄ1���=�3zU�oS���&�a�q=�9�&5\K��&*����Cn��B��'B/\)���K:po
��}�H�fE��a��o�Fx8�u�3����X��e#�k�]E9����S��n{9 ��,�V����m!q�[.y�ŻZ� 
�a���bo:pT��wS���^�0p��co�a؂��,`�v�1R���-�
dR�g	4D��LL�l�b&���܇��n�Z?`�4:��Zq`��տ/*��T�r�V\dS�zb�^�x��O����ۗL;qJ�.�.!����'A�#����t��Ap긍勱C��e��{Q��:�_4��.=�g��%&n������
m^�vp��7�7�I;��-Q�Kv�r�wwvt��^M�|S�ʹ5	��8�o�����D{�G2���n�����tI�č%.X)m%��Qbƺ��qS�X���|7��]���Q����ov*��Ϙ�DL��+Mʻ��<Q%��"V�r��J�vxAv|��W;����""o�3��� \)��BbX��2�����Q���ɖ,t]�!�1�;�m��#Om���ܝ���0�Ξ�F�t�8�mQ0����Z6��#:o�d���lM(�k���M9s�x]�n��'�rc��ږD����m;w�%����앸�L�M�4�o"�3���.6d��r�^�O���ieٔUÀ���lqx��at�a���w]}alZ&wNEn+�a/�(qB��V��KJi�jt0a�ܦ�/S���j:�Nr��kIFw�j,j7�������1C�`Yh�)�H�EN@�WKd�-��tT�$�[.���w�G�p���+ۊ��j�)؁a��W��_��7�!�uRfo��
�,�l��%e�,΅
ԓC�aӘЅGJ�ᚢ^��s�9�p׃�S����¶}�v����J?cʇ���V���ݏ@��]J��+�=�`V����]i���$y�<�v�쥜�����V�O]�KwS��y}}ו��,n��A��fk�IN<���ty6�ꇥewvL��0W�e��ZH����Һ)�h9W��Hf�g�~�D{�蓙}���R���v���R���a��1�\k��{����k�b�d�
�QUѶ��mu��b
�&4���/F�b�������&���k��jڕk� �����n�Q��1m@�}0P��adדPJ�$ �m0��ɠu�\_�����s��F���l�o"��C�^��M�:��Ꭺ*��lX����xݎO%�gT��]��1��/�a���,�Z|��ϻ�4�o��g����t߆:���V`a]�5�Pki�bF��$��·8<'pNȕ\��:�HWz �����k�u�~s���n6�S�ۗ�����;�RD_9�ÓC�����\CTF�BCT�0�8�옭Ywb��^��'�&:�z���2p�s.n1ω3�&s�`,,i����.�U�(�
O���޻��#�0�Yh:�v(����p�'v���:"u���T��.Y���=�c5�J1r�a�~Ƒc:sc��g�yU^���xL���k�'֬s�$*{-F�;��%d�`�e�+�:��՗ea�l{���L�s����]�,Un��fr/u_��u
pU��Lz��=NY�.,�u}8�yB�QS�_sJF��tfί���4�E��m$���.G]<%���Tt��l�!�Z��k�F�3�>���=:�dk|�p9(�����nR7�ӂU{q�,J쥂��1J�����l��iu�̺�Yљ�-�'ڡ�_��i�-1~z��N���݉�G�Ҭu��o+a��P�f���yc���˳]�/�w.�(3��E�A�t��ڧ��S��#Bv�F��:��NB|�n�Q<��E�sq>�(��*2�b�>�.�Zr5��6۶5�W,�5��}c)�Ŧw^�О���8�H�۩�S+����q�#Qoi��q�у�:����1����aX�W\��2�93,m�*��&c��<�s�S�p�_�A�ξ�)m�a���jh8f9����wf7,��K�:�R��U3薊��[Q�oa�����:��ma��A#�a����VS�Y8�@�P�����HWp�Z=�1,mD\O���R�:u�S�y� ��0�����^%�»90�>R� �(t Er���T�;Y�q���m ���^����0�c���p�����@��k5a�Aa�.��$\{���j��}\���m}mh#�֮3�s4�� �f9��N7���Q9I�ô>�����]ť�B��::9<Y%��=e�ZǇ}���N`�a��!<1����6+v�Nɔ�Ym*[MA���P�Y!�p�+�+�}���"���e�M�%��N�u��M�����u�4�� ��+�>�=W��#�������Ҋ�=�|H�R�sS����ѩ5Z�}�@,�k��c/�%ۅ�@M0��� �+�ukZ��K�3 1�j����Q��ϒN:����5�ml���^��q��Y.�LIom�����(gSzFI����ֵSmT����v�T���fjN�Ԥ�*�OJ��t}�tU��S��16�ھlm��n���VQ�ϵ,W�5WFc�C7�Zko��"�ҥ�h�2��|o�CL�Z�E,�\�$�n�]*+ [��j�nb�-�v�fsS�.����D���EM��Ǝw�z[��z�yT��g��;¯�VA�pJ���[��4,��pn�zd7���f[��c��S�S`\�ެΛ*i��S�7�v�_EyF��7\-�|�ή�$�֪�l�[ǲZKNe��[�	]��7ӡb�{�"�1�M�;Q`Ŵ����BE%|��m����tGpڇ���no.Zn�2�=_DmT�Г�**�Vѹu�׏Ol������vkW8��/��j�G��%W,-:�ݬG�,A�R΢3ju�עt���b�Ӛ�eղ iK�X=yr�:�.��a�������nwS.�.�.n���Lt'��=���)�ε��x�5�K���$`f��9��pH����}}N�@r�J������<ܾ�>�+�z9�f�̡��&����z'�ݾ�������V��u�W��45�}ΰ<�o7K��#����-|���Y��D��ƍ�Q� ˝�NZ[Ϻ#�r$��Br�"�NNZgQ�4^;�+)ԛ2���oP�wLY�tص���]�I�٭l#v�q��h�Z�*T�M��Ґ;���[��2Q���G�#�\jg[�WѷAM��I�Z���Y݃����Y@���t� in�PI�J��uG���%����JV��.yn�vb��L�w0fU�9O$�$ba�����A�/�E[���ؙûyf�v�"��p�݄Vp�;��u�c��� ��F�Y�f,U�妵h�
�5#�B��:�o+�̽.����J$W9���:��{Û1���-�-��(h.��)�\$��ݫ������3�h�)�f0�=�5��ڬ3��wd��N��I�����+I`C�v��(�ԫ����V�s:��q�]'0�V���f���p�KepT����Z��v6n�n�[L�iCy5	�������W
����1m�7;s�1Ƭb���ӑ���O�ӛ�����T3��R�_9�Q೻L�m�s��w�N��*�U"�
�����P�-Pbf� ��ⶋ@j�Q[E�,m��Z,-�����b�"+TB��AQ��X�AX"V����TB"*1EFV�(��FH����F$S����(��Q�����im�"�m��b�J���VV�%VTYmX+m-
,PET�ŋ0�*��AAnET�
)TQDc��h"�IF6�B�QAQZ��QAK��U�j*�T`��cl���"6�
�D[VĶ��X��,FDjJ
"�[Eb1���*�R�G�,��+ZQ���"-jʘ�kqJň�eh��b"��[ci,TDQbV�
�UDDQ�F��XUX��QUcQV*���AA�1%\P�EDb*�JҤQER�P��IQf-+%�#�b��V6�cYVb�U�*�e�V,�A���c��1J[QX�*"��YV�UUQU��QbT[�VTQX�QEV+UPTE�T�EU��QE�*"Am��C�T>����[W����H�Ky��x�;�Y� c���/f�9tv�1�z�kb�y��8ҾwDr�9��I#1�}��}��f�����&�����Ʈ���J��^:��V$�Vy}�uR�iIgb�#G��Ñ\�1n	�ݞj�tM��p^Q%\3$E��,vȊ\2<u�k3ʦyjK=F��s�P�,0�d�]�x�$��Ɖi��^o.�X�&ϥiDe��/�������yi��X%�Y�o1_)�qR�� �t�P�R�s�ԝ5��)�������k�D��~��ь��^jݎDE�-,�m�:�Å:{�����"��F���sÌ��Yg��k}�2U�)<�V�B[���K{�oc�����*��K�R���G���x���S�0�'���F◤</^S��Y#]������3=Y����q>�g�R.���Pw�>��w�w�Dxsx����ݫ#���F��ƃs���<�+� e�	���¨�黷�
�v]�����Fc��/��Ѯ��5JN�7�,�u4�g���/q!�|��Ϭ���Y#��P��X���9�!����q/zs�Lj.��a�_L�{$�~�tP,�x�NnY�t�U������T��yj��4�}7��=픍��.�����6��JA�Rڗ�j�y�MZ���"�zr<N�UӜ��.�>s0e�{ɕ�Y�:=�I�}I�g*K�$x�nɎ�kB��}�Vu+�G%�#`Wh��K�z=���z�ˋDmϽ��������呐]7�@޸ט`Ey�!@��H�D���Q������A�v{�R�fDm1�͔6"��b���̂�[� ]�� w����.������w'�e44�������r�vci�6%m,5����dRs8�-�'��1��kPf,6�U�xZ�x:�Qi��f��StU1^�0��yw���]Uc����m��k��^�]P�A`UW��D��~�eD\���e����ͳ45���^��ne@m��+��7.���YD����tc��
P�<*�����!��� }��}̹2��3���Pa)#+��\<(ᇐ�����J�,X��MF)9/{�]5�Th}Ӗn��k�*�����5DD����p֍�y�gJy��r6�n=Ա�V	�s�B2����*62c�@p,N�M��c�y�h���3~0���86��B^�lg���]������6�H���Qc/j�âVLZ5��0b(�����1z�me4^n��g�W��d<
=��F�����^�݈�� �z��B��t�8������,�W`����n�X0��`L�B	�l��:e�n�J�2�Ye�G�fh@�kL;E��0�`^�I��+��I��.�'[)V*�U�zT�7������Ѝ�}|�V�ԧއ�L�<��s��fK���:�^�5P1M%��\�P�$k�:��4{N<uñ^^��lp�bz��NRFr*r��[ \b��o\��2��Qq��m.pͣ�!�j��3)�Ƶ/zX��ꫴ!F�/C>�=j��nz� p����i���n�b�\_N��\���0�Ƅ*#�m�ȍQ/5_��ᾴ�\��/R�[�f�
�mssf礓nv�e���ӻ^9��5{{����L_���o\O#�΀�oZ�^&*7y��C�;�5�y� p�T3Å�0�&8��=�/��f����壡���>�.�1�ם��)Rv{�L�E�!���B2�L!�r	C�g"JoS��kt�u�'U;s�|�4%T_�ȨW��DZtB&�>t�xc�*�XM�C��r�ww5=5ָZoK���pG#�\�r�:��N�w�"i��|Loφ;o�,�(,v�7���UY�Ê�P(�����4Ą��!�L�Ax�����Դz�����v���+s\M�9�@٠,/h"�TX�R�d�G�q
��{ԡVi�n��]����w�;��J��ֹY73/n��*R+X�Bhp[��;F8��N���f�S���V�ۃ�Q�v[�����l�S�$�f.�Ftw�������NN���}�RRL�u�[��0~zc�/�+	;|<�m"�j��hH`"(Å�e�ll����oT��*�$�Y��E���0nT�9�&cL�v�XXX���1���t͝�3ܺ�U,٫J��8#��!������g�zZ̋�/
Y����ܲ��m��Vl�Q�RgN�������Q�����:j�b3MyțӖ�s-`|D��c�eG�ήd�o���P�|��0�n��r��o��^�z��lW�Z��[���ҽ�OR�즷�sj�k}<7T2���>�I��,�'ywOX�r��Æ���%�w���&�s�9����*U׽u(�,#qH:�.���0\6���yLwd;̍�3q��7��VL
o�U��Qu�@�<�MCj_�����ȣyH1P�S��Ӯ�9�cY46b���u�O'�;�F�ixп}��'�2P��L��W�9���m�ބX�L�r�4LFaJ���]�.Q0P����WH58�C��2�G&e���*������X+�:��%��9�)
v����4+�3��՞u��R� D��ܑ:���}k.�ʾU��C6;�)��̄�g�9�]�=�\��ƧQce b�BV��2���7]SG6)�LU���z���P,���&s��wɚW͙Q����#)X7a��rh��OI����{V��h!�c~�M)��f9\޸�uc�0)�d�
]1��r��xE�N	ˤ�z;�ۗ�����Ni�*)jy�N�d�9FL8I	�\��W�bX۱����u�8�J�P���%�i��׶eہ,1P��τ��D�ЁI�=GM������pS�<�v�9�W"�f3�c�DZ���΍ 1CvJ��Xq��:������i��s��=:dz��J�a��GY�#��[�k��Wʱ%�뱋hmI����l����>'ͱ������� ���v�'�iDT��m�����L�ҭfyT���RN�=J�	Mg4z�vS�0�8����S'��lA�M�M(�����U�'oÄ��	�nٻ��Q!��S����'q	�VW "���q�:jg\U������4ӑ80�>A�j+�HEm��J��G��4^K
�΀�]���j7N7<;���sME/7Czl�J�g�M��e�ޘ].iLVU8#8���qrl(��&��S�
�F����GQ=g%���(4a���׵���h:�J�L®E\'S�]�8<����T��<��ܡz�_+�
w&r��XzJp��(��<7�)Ӊ�����u�!��V�Qq'ı�R�u��BjL��&|����7"U�0�YBFd��V�ܾ#�}�z��Fꧮ�n騬R���陸1�]0�TY�Y��#1ʩ.^e;q^nk�5W4�\�ʾ�����c����6�@�Pŀ2���<�x-0�gdw_Kj�*�V�S*�Iť�'��ȆXѶ��
ST��n��&P�Y@*����aas��X�vf�#%���>�����e�՞so�Vt^���%\OP��w�Ep�My�)���B'3H.Ԁ��TK���~�AT^V�%>W
�˦�\��z��2�(�)�g�eR�[!�E���ܞ��
�t��R��r�f��ͤ%j�)E:�p0�H��Z$�a�Ʀ�-f�sέ�@"���
ˋ�0�/�鸂��X���`��f�Kf�E:k��E���;�������������Ю<uŧ��٪ו^�L#��s�����ڻ�C��1��8��ϗJ~�k|H�w���R�p�����qU���g�JL��#��`��_�
�
�|û�	��)�zK��{[$�J�Y���q��Ë���\L�.��f	�{�q��ͮ��ff��g�D�ԧ��o�s��3�s���������L�y�kiP�fk�傤���]��v��Xo8L�7�I¦����!6�wv��Y9gah���H��r��S�ó�u@��v*w�y/�=�q��o�`eNٱ�9Rf�e>يd
�������=�YG<�"Vt%֋��Q96wq�/gA�Ƴ\=R��(p�)��e��	\p=&ڢ"a����Z6���sp�[i�9�Զ.v{�/ɬ޺[E��k�)h輘�j�b}���kv���F�}B�u�i"uS�9t$>x�EZt7���#7U��nd��*�
�uj��n���r���-�K:_(��/�ή��}1���Pf�4̖)�E����<�tKNj{j���D,�c��q��3�]�ѽ
��1C�`ձ=f��)#9꜁5�����S�o`u^�[�;Rv�:!���O&:5�|�|,1�|R�]��v�>�!������'ćW��{$�8�Xp�Q5�Xf�)��hC��ѝ���,sɫ0�)�m@�W./��.z��Yء�p�";I��U�B.x�E��i�+��LZs��\O#��t��H��5eY�gw�r��`�(��2�`�LvDK������b�3_�~ע�^�� �R;�m'����ekQ����:;��y�)6�9WVIK�pEݑ�/�_��^��&0v�d��,ݑ�׸�@4�,�w��f�6���Ũ����a����E�b�F�&��S�w��ca��� �@D��,��+h��z#�oo��4�p��Y��5�m�D_�-70P��
�Ƽ����(<*����dL�Z�q�q����C)�u���*��TӼ��c~|0�𼊀��b6��v�n[9Z�qh�[����c�G�ƫ�)�E�Tu�yrL_1(��S�6����c=z��gӁ�˧jy�E�<=��z��k���k��p*|��?�6+�= t������Gk91<�o�ؓӏ����c�xH��[m&�u����TFלؠ�Q�*>���9�����K�90K��_^���.#��3�N�(�3��r��.�Kswu[KB6��Q<�������x�u���k�cg=V���&
���;����8���a�����C�j�=i���I��^(7"*P�٠���BM#�� �~:z[���D����;1V�i�F�����'e,���)�|,�^tQ��jV.zOp�Ǒx'��s�xc�Ϸ�c��r/��T��+u�.�}�vS^gM3D��Y��BA�c4d�����v�uF�Ӳ�d���ĕ��:�u�)ݥ�w���xMc��)~���? )��v��+(!�o���Z���Q<�m.X�]��WNo��ˮ����٨�����K�4�c���#�!
�y�ټ3J㕭�#ѵ��Z�ΕZ^��b�D�3�n6�u
]/���0_���#���\���*w�NY��2{%�����]A�jY�4�J�JT���Y5g�F�a>�s�\F��f�h�y�(��W=�N���ނx]��+��M���Θ�pL�6�dG�̬84�X�^/9�or�S[z�,��dW	����'Zyl#n�8�FXh�e��>lt�J�g��э�+{xwc����cSe"�v��.W)��oT�q>�uF7,�Ժc���׮U��12�Ozw5�����헓,*��a	Z��u:哑�Uj���q7���+�y���)ĸ���s��[���K�S�l���(V�a���R�
؉W`p�
�6j(־/��&�,��ҁuS�q�7[��|����u�X0B| ��k��3A�x��_����iGsa�j�pMX<}!��gͮ�]3��2WJ�^:�_�bI����P�҆�v[�Cw���kP�(�?'Dh�
�X���.�J"�~>g�y��+���V疤���{2;U��^���ZX�`Rx��w+�ɵ�,WU����^��u!G{iaA�>ޝ�V�4��6#좀W�#���I�$0���휄�VT]pJ��wz��)E�Y�^�I?V��NZݵPv�5>�o1DC��E�ef+[���R���GWV�-2�xLt��2BrY��;�n���w.3eS#UlEe0���-�F�!siV>@nN�`p��5�� �� W��zD�����Q�C`(��Ȝ0����:�wz��_���x�QB�mX�3�:G}@`����ݨ�9��x�$\>�7��}����v�;�	���a�yD�>T�p#Q^��:]d��LF�֍�D��@��Ů�g�,����Y����7��V3R�wJ��]A�7��R�x��m.^5ΰã0Nwbc��֢�!z����۫���܎}!
� nP],Qg�@�dle#ov&����D$c�"�t渖7�`΅uT)�Rpcp���SLvz��Ur�#�LR�'�<P�ғQ�\qaխ�VH[��Q/zy��J]�*�"T��H�̽�e@t%�qHzBFÝ�&��X��E�hB��p9l�r�Ƽ�*b	��Y���\2m��n�]�~��ݫ���˕��\�ّ�Ǧ�i�Z���u��`Dk�A���+"�rWJ����T!��MʖA����zV2j�Y�di��#�;IUI�Pͳn���{w��G���7�[����WUٽ���qz{w�{ooY��8B�����J�-����i
�]�'Iy�9��t�s����'g����͇��ۨ�^YK��bXNT6�j8Y��j	��Au�6)[
����L���h��i#��
�ƕE%�IwHY���vuNz�|�^�)*n�9I^)c)�dl��А+���� \"܉�Z�dnl&��|f2d'#o�Wҋ7��h��Q�:'ڏ�3����%�u�\h5��$e�g��L�]��̈́�l��#p*;M����9nS���31����f�J��e�\�[��/��l�x�#r?:�p�{HO.� ��H����G1��T3{V���F��M��U!��MX=^`��HNG}�V����ud
������uTSN��5(^�3���
��ym��)7O����f���Z�le3�l(��nʲK\V�8S�es*�,��w?�M؊
�4ڭc�3�+j}���A���:γh��Ԭ\��:�rJי���m�+�^���Y���R2��R%ළD76��5�ъ0%�W}�r�:U���{s�V�|���N�wX��;c�(r��8��]̩z՞��� �8}�tO����t溇��[R��zv���*m��-��]ʃ�&'��,��v��".��*c�]�4V�K9��6*JU�h�Tr�t�k�˼ ����Y%�H2%�71��qݦ*H���u*m�S�7GX���]hv�0N�4I��ع^�O5Fqѽr��<&�۲뺈�2ƨ����N�����ȸ/h�c(�������C5.»�dVP�sh%��Y��e9*e�:���a+�˲֗�D�Q!S��v]�\p�;6����M�Ӵ[̵�m���J�+��yb\��d^k����ֻ���|0]���P�[6�qoд+I*��C!T�7��5	�jQLc-�h�}��.�n�*��AYҸ�n��R��!X6�Χ�ϕ����e_Q{��%��mj��tTj:�9����t�.�t�л[;A-����oEi*���btһ�/��b��s�k���A��0���ַ�Tَ��9U�gJ՜�ᓖ�1��aguvV�\�&�r��τw���7�X����{B��*��-cu�Ľ��x+�,�K+�JpA��m!o�~kf�W:r~����_v���އ�� Mu͹77w��m�P��:�,5 ۩V_&������)Y�u��$-H�a�ܶi�5�M��=� Q�X[�DWsx"��l�nvR������`;f����}�衍%m�h���G���h=[�{�I&�zk�AN��	G��vA��h71Wvƺ� ��s~b��=k�k�Lp}��ϖ�����ݴ���k���
!�|]������EE�0DEb)Z(���Z����Qb���UJ�"�Ң
"ŉ�PF[᪪*�QS��*
�Ab���J1��me��,�(��ԫE���iQш�EJ0�,Em**
*Ԫ*�1EJ�ª�DQcL%A��Db*��E��UՌX����b�
��
1��F$V �c#RQED`��Q����`�Z�+Z�KZ�����H����Z�m�DUb�b����UV+UU�����UEV(��V
�
1R*��U��"���1F�F� �b��EDA`��PEE,Q�b�m���ZZ�"�`�\YPDE��
 �k(��F*��V�"� ��"*"�A�(�*T�5*����UX�����"�J�m���.-�+EU�*�-�e�}�����j�e]_m���e|�ټ�.��ﬡ+;�|�V�\~�>��p4�Ipuו��V<�Ȕ�����s�������ٽ<�6��X.���+����i���/���}�X�Q�T�����V_nk��z�m�f�.7���"���>�:L��­+����ŧ�[KʯM,od�XfN������W�³є���qLYwD��̑�̹��2�Q���坘�L3���e��8n5�z\3�]�wn�$F@l�;�ww�$�q
D�7Y�uHGE.�If��r��ޥ�ޝ��x;Ո�X�
يD
�p� H�m��5e0�+����^���{{x|/<�E\/����l�N�vԑ	��m����^K�_�%!~;m�t�~˿/GK+¦̓��V�T�U~,z�
�qS%nKj���'5Զ͵{F$Pu[����e�A��1��y"3u]3�o�z�����Z���y���/0�v����1>r8Q.���w�:�\}:-�֒�[xxŚV���'�%r���<�֊򮦺��F�N�p��e�&����3�q��W���#�lOY�9]��a����<*A9�eR����ѹ��-�����j�V����Df����p�)q��\z�<Y�6wd�o)�P���x
gtU^�^�
�)'M����;���]>��S��9DٽؘiJp�p�r�Xhc�&�7��<uz�d��_UB��������c�ɿl��aoOf3Z��w�����NS��x���v�G9&� 'sw�q<�����V@b�d�)a���aҘЅGJ���^��G9c�MY�8��q�v�,J����i@�xF�)�M�]Tu�Uq5�R�ݖQ}�ŧ1�޸�G������q9��i�ܽiUv��g��u��CE^a:�2�td��=���+�Ñ�X���c�Y�º]��}i�v�Eұ��pxs\N�z�
��/ď�>TxRzp��WD��Ĳ:����.���9�h�"1��h_���ɡ��:ͧ�P�!�����Oz���1,mE� �����9���hsh���7%��
��)�W.z����*9;�&6��D�S�6��Kșݎ�97�����Z�'G�c���1{�����*�Wk��U�:��v��o�<�����ͱk�]JG�"�����l�jpL�e ��@�*BB^�ԑ�r*Bl��W���w�T4!��x�������h�͢Y��8~^π�P*zz�(�^qJ|+�L��_4I�W�K/Hz�^�+&p��s��N�[�x׻��v��OP�0ʺY�6)�F=���i�M��`�Dn�jA���we��#�}�q4�v�@4"�������Q�;&݈/vdʘ����.�E�`�q=tr�`Y���9	%w��uwn����.�
?y;#EB컠����qDm�C�ɞ��k2/P�:!�`QPec���6�N�Pq*�\y9�x�N��}�t-v��W�1����9t�u1��(�*\T9�Oz^wPܐ�a:p:�u��1p�]���#h���M�؝L�����r�)Bֻ��h�&�.��l�E��:��Ρ鋇��t�<���Ǝ���t6�1<��r��ӌ�pM^��o�2�JV�P.3�o�H:�.�\ō��==�����d#U���Tzo�����#+l���i�
�R�3��p�2�
O��\�2�;G��=��U�w#0�vӾ�C��/�m܍�tţ�%�TȎ%p99��Du��zct��s�T���E���\Oq�pu�yl\)�rb2�G&e��2��u���q���,)���-w�/�s�p�>SC!��sq�'ݎ��l�z�.�옖6�=�(�,�F��D$mq�tEK��(:��0�R��*\�L�U箍
}�i:'e�e���o��v%T�u�ҫ���6P�W@W�̽��1@��w��U�ƍ^��7�G��U��=��ыq��C͋t���W�~����]^�l��u�����Рl49�oGK�]���ӕp�m��煗���kv1=����t�\:�q�?���l�����C��g���еM��T�ګ�89椬��u�3�3��.�˞�`�n�@�}�^ci1,Z'NƹѢ�b��@�Cy����M�;)�ѿv�⟻����1�F���xe��xc��J�V�u;�Ig���|p-�G"�JйY��X�$ڀۓ�b��4PwR��YD�q�H��X�;%�ʅѓ��7e����B��n*�ܜ�jfyA��T(	Ig	����]�J5�;��<�S��Ƨ���VM�2��媮qL�1�䶬^t�5��3��^k)�-��g\SyGP/c�k�}���Z宪�H�09<.�e�h(������ݑov�t�{�.�ʲ���C���������2���g)@�W�R|>T�>~=N#'����G�8�ɧ�����&���寋��U�Ὦ֣qOdr�g����0�u�E��G}���=� v��A����q'��XC�[�5V1�w#�HF�s������WK U���˱���:�巃��H��4$x��F��%*4���+!�Z �'#�=k��|_�sPz�J����i�n��oD�'�t-��Gӝ����4�t��%YK����k��{���f��s�Mf�\W[�J1*��q�=I~���Tq�j�{���ч^�U=:ౚS,hۅuW��)81�uac��:n@N�BTù�5��j��[D�F�s��� ��;Kޞpc;��z�W�'ڗq��V�Ġ���t����뫦G?T�.%K&��~�AU�hBS�p�8�u�3�ݘA�M�CW_gv*s�v��n���2@�VW����.V��̍�=Y���T�8���v��2l��V1VBi�{����] �oB�s���5��*�.hUΧS�B�����f�#pT+Os��v-�B�5qN��n%v
):<M�U!&�B6�B��;:yҸ��sy��I�%����/��V�F�uM˔�!�d�7č%�ߞ�S�[�ō���S��Zmm;�p��k��e��:8f�v�6H�����q.����Ib��r<%��9�o���l�L��!��?B5��f+�ҁ���% ))#)����Q�\�s�E����_���Ռ.�M��͎´�f�v���6�莣Hۇ�D���r�p�]A�5�y]��J�+Ԯ`3n�����|��m��nc����I���c.�'��\e4��n�$��G���xΛ.oFӃ��v���Xx��J�-s���游h�ś$�2Y �3��W*��S�Y�-/��3w�i���5t����ۅ��ΖI
��u�HX���f-����� �=�u'��g�Vc�#��l{N�2���+��j�H��W�>�7��1h��&��Gl�6�Les�X���VƎGIW҆�k:�C���kIN����y[�*�O��a�~ٸ�<z�M��, �ǃh�^F�o�	�����.v�V�˧f��Bb��w�8Ȫ��vr��Y%���@�[%l��ap)�Íj�)�a��t�j��0:�����gE3�|�﫚uq)CD������p�?hñ��-w��JtG^TO������� �M���2�u�̈�7諪�r����,=ͦ��a3� �{b�<j�2�q���)z�Y(��(!fp���1�� @�<�~�[�&�y�I����/��!<�DO)��^��F�^Q�m�DtZn&
>��0�k��[��V�*�.-"�����!o[Ny��ȧ1�m<��p�n`U�D"n��`���^ߞ�^|]�v�:���.�.�b�Y�缻2�����ڠ��ނ>�ꂔ�����[��/�xhİpZ=(7����(���p�N���j��{R��J�Kk�����m�-�;��-�xh��\ɭ�5����w�D��_G�뜬�\�(l ~�N��4;��IC6�:��j�c�NX�.���˒b�|�"X��F/b�2�[�7�kxu8�Ѹt��;�$��f�Ml��0�5͊��կ��D83�VEٳ{ �k�Y��n�]�Z^2�c�x��9X������T�xBw#r�(�6�ge�׽���P1�UB���v�#�׉���,�E/��J��T]YX
��$���b�n�P8�7�{nF%xث���a�\Qx��3׮��N���q����Sj�ʗ��(��0C�q0f��)gI耴�}�lO�q�.yU^������yo$��#m;��J����xJ!��L�~ܤ����w�S=�B7�C잓AdQ(B��;�d8t9gn���|�uHe_U��3e2.6Pi̋�s�zbު}ӯ'����K?0��ˤ�c��	�����n9�w6�+�n&.�J�J����,qs6T��]V���8g�/Zs.���s\�cvqu����U³�R�����C�xʷ���{_���>O�+r���ˢ��d�`Ě{�y��ʁ�%M-	�w�5�+$��(�+Zڷ�9E�N_��I�+iVPw�2���]�_	�ˢ���_u^��-Ɔ#�Vb��6�������N�'m�x��� ��x^^��0��A���h}�������Ι��&V�8�fߓ�5��yL[�w#w�����ᑤ+Z]���=���u�8��^�aţ����S���\Oq�''t�)�rb2�G&e��UAV�v���m:��u�sPN��'^NALEf�)R�M�+����uc�0,���c��LKg�mn%=2�cH֥Q�P�OYܙA��o�jy��Ny���A�PI���I*6�k�vm�D�S��o�Q,_ð\���P��,1TЭ�*B�9�eF\�Cz�و=�d
O��Sk�q�Su�\c�Z��Yу`�,m��	��r8����t�B����T���b�c¶��[Z�\�]-x�w�X��ٖ�.�����-h.Isë�ê���v-�#Eu,rI{�H�1�rJU�{&��׌Z۝���16\����zfs����l�ԝ5����XN~�$nT'חm�UҶ�	yJ�u"�tE�p��1~�ڱx�A��@�@Ʋ���8{ϳ�*έ��Ge��3&����C��6�\"��"�V�,��	���ł.Nݣ�Z�h���A=���eu#r+5˯�j�t\�.�]����_)�w�����v��.���>άș�K��8'��9�8x�0\�ꌗ��S�-�{w%�I��`M��{�꫼�R{y�`r?{dKB�e*�Յ:{����ݑp�j7KgF��'vX�1_d
���T�e]THՈ�~�1����W�U'��T�(U��8�OQ���,2y���+����N�Q[(F�;��"9�p�����9O��5-�j�=U� �>;K�������~�Y�Ľ�
]v��(1ۏ-�m�U�o��}A�)o(	��� q�l(�C�q��~=�,����+�)xq�c4�Xѷ��fT��:��Φ��q��{/Yos�焽+��y+��qPV�� l��(��9�&5E��3� �M�٬9y��JZ�X�z�=�E`�Ms<%/.%ߗ
�k��^V�/ԟ,���r鸍r��g-�#����_-��D=8!@�t�GLW�G�𔼺�>\6��ʝ��gO"��یXg��N�Ƥ�[��q�X��\,S�����*�.��\�k��(ga�07�ƻ����T]���4�yl-r�0z��=`��y�&6�U�p���u��N,��ݱӔD����zk �֐�Ύ��E� v޻tcO���%_ISݥ��5�g��R^=oo�Ն�f�o!��H5�Ya;ԪBq ����{S��Aų\fa�A�X�1XT��ϰ�juj�Xγy�d.��u�;�3���U%5k��Z%ޟ�f1D�����p�!�d�T7č%�碔�K���A06Q��s�-QFF�q��LW�Nʞgw��a�D\n^��wp��$��*�h�`v��]���$�xc�|)T.���3�g
J .�( �"۹�aJ0ߧ蹾�����x�?2%���ym�Xr*�����b�n7@l#��/+��޻�/;)0�%�RD8�nⅥ�n@R3��B�ؚb2�n��%F�Lc0�Pp�F��{}4+0-�Q��D���q�Q�C��F�nmȧ�^��$Fn�g��T�<,`��C^4�]1l>�Z�:���({��H����S�^Ύ�t[�&VH�C���9�2��t�������{3�da������SQ���1�3�]�ѯ���[&�ӳβs7w4��#������,2�S�&�S \b�ɸ�B'ܶ�_Of3��>S����1)�SF�E�y�����+F�):��j�Ud�'qK�e0��cB�T�5���al��L�\:T�Ѱ�W�I�}��6�w��D&���[�������U�E�!��z��Ν�̣dމS�i�E �ʙ�������7z�X�����Tt��9�j¡���j��v�^�Zʰ��ug���x�M��y�O��aޏ�[$Rv
����Գ�uh�� (���V,.Wf;7���Py��Gl�a�i�Pٽɭ�o���Ԇץ[�,j��{�+[F���r�<�T��)Vs�ZJx@{.ɢ����K��(�\���>{L��}�m�;��Ƿ�J��D
�kt��pT7-2�(#u�5ѵ�˱D�>{D�T��������د�V9ׂ,��w]X>6	u�q�e�B.c�2s.�v�f��Ĕ�2vA��řts�F�n�
��J��n��W�J���S3H�����Sk+���Rq�n��1f�d��RTĘs:�o7v��]� �}��b�r��;���h����*`ܫf��;un'+ޥul�
te]]�~������������+����+C�
`��n�^t�*�.�T��;d3/���I�z'�����r��_#F�l❘-p��Rᴢ�j�j���:4iaWo*,;K�goi��8���(�:�Vf���+�M/7��ļ��G�X��;B�WB���>�u|v��BJFD B�wA��Gq��&3u,0�R��i�)�1m��s��(�}���f'�m�����)��J���0a�帳6����NV��f���F�=���5�/�n���
7�0����jg�քywf�Ԑ���+ދ_.g^e�f��3j�gK�,�����p;�T1`�H �-��M�ս��ɨ��.�m5�� (�9 �S�;�둢da�V���V��h�����ՙ܋gi�Tq�c� \�Q�տĸ�5�1�f�����&owS�YCyh�����:�%�9S\��x�)$���TlLIdG�Ƿ�w.FC�k����g��:닆m����;��0�Y��0���O��O���l�}�%u⠄�h�Q��qf5�2�L�u��zI��"9\:s� ��e�͙)[g�S�����s0�������M)�
����)_gl�M\+�`yyx��>@�\�l5��!�S;h���F���-�����YK��]���eܚ��PJЍu�V�Q��46��܏U�!�#;��us�6k;I�Z�8ꬕ/�4�\����`M�j�IY3�U�ݍ;��������˙��ǅE�@�m_X���yz��`�u}]6�f 3��b[�V��Ɓo�3�E�,��mȜR����O���y�c(���X�2��S4WW>��Ŵ��D�^������&D�������N�C�(�p�l���-�n������u�r�xc����N�4�Tܾ}خ�ظFq��V���][ݙw�](��µ�+�QAF"*����(*�%�������A����	AL4PX+F1�Zؠ�E���#J�EQ�Ƞ�
�AKh�B��X���X����ʭKic�U�b*���QU\b�cZ-j1��*� �*8e%U���EŪT��b���UG��Z�"�TjQUm��I��U�ac�b��DDT\Z8kR�EG� ��*�X�h�V*
"("��k
�J���QDe�Ub
 ���cD�(���b+Ŗ*�QUPX�)��"�*��X�1X�ab�[EQm�Q��*���%�G��b(��F(�V*F--1La���QAkQV1�Dh�B���(�֫�UF5+QF*���TVb�c  	>0��yZ�S����S�ܥo�JśP�A����7ZA��\��XQwZ����WR���v庼tT�e��9;�����ϭjY���(�e3X?Mr�3��³Ċ�<�u�s�j1Ksi�/�X�̮��5V����r�L�qq	��=�΀�o^S%
��Z�����0��/��;d�]yK��l�so���@�SO��M���渝F�^Q�m�D �&^��Ы\y���*k�|���0���t�M�se���ϲ�E�28���^��+���d����s�O�0MJ'0�g}%�s|�5\��^^�>t�gz�&����[�g����Q7y�z��[k��oV0=zEZ���F�/�1��n���ʸ`�.&�"����u��k�p~.���M
Zr�Z:���o�}x��9XI���kY�
���Nn�n��u��!b��:#k�P1�(�ק�Q�R��xvjC�6��b�wnn1ω2V���x{ANU�M�s���~��`\��7欍��wB���X��J0����l�S=+�5��h�̇�UV�����̝>�YC)�> �v?���ފ��G��5^ʤǅ�Uؽ7ry4s��Q��v?x�,�1S�ܶ�n�����u����NLN��	��Y-��h쫷x�������[.�C��>��v���L��vԷ�,S�Ok��bu����E'�VG�bSy޾E�ݝ�w/���)�߾���z=6�Uy��'Eq��S�u��H[��OBr��o����CD�֩�U�Ln��m�fp0���uLeE�XP.3e�/�(:�N�e�:��/�U>�vtn���1��խ��U���#8�.�{M�\3��Δ��.K��u^426m<��!]�N�yHwgי-<f��@�R��������lr(�Rej94��@�j�MfV�d4|8��.5��6�cY�yL\9�r79����D��K�u�c�4纆�c�_^�!h���_ͭ�:c��k��.5���O-��w!�#,4r&e�U(���\�ܹ�m����1��Y��R�N@�f�-�*|��ʥ{\O��ـ�d���X�N��nj��\/�4l_��}>KE@�-�/�y�op�Z�EdE:哌���VF �t�ڞ|
��d�F�M�a>ֻ��*^��|E��ϫv�{�!b��m�s�Y 
I��-/��c�=�@4O�Y�S�G�����k"��`�H�=�F��s��U���ɨ�B�\�ˉ]��UӢ:9S&�0�)g �S��\���p��Z�m��Z�|�bO+t�����AΑ�5F���v���6���_n��53�F]L����f۔�j�:M��\M��51NP��V���JӆEM�-���c7\��]��|���ѐXc���*�L��d��S!��ۅq��M՜�*Cbro4U�{��Aƣ�.f_�O�@UJD����!��VQ%�q�"�u�؊�6�-�ҧY��������'��b�z��f��`�p1),�6ԝ5��VM���pऌxkv�왻؛��}y�U�/��%�8%_���7��N�����N}�qU�Ix����*M����F3!�Ǉ�_���V,O��Q�gD�*
;gC��@`�v�d_��F鹥��:-�BVܵ�ҽ�dS���H�}�n*��c5@a����m�	B�ǩ���|���U��vZ�h�G=�%�|����j����=��gN{�S�X�IY����"�ftoePEs�G��aU��Ӫb��ia7C�c�p�����vy�l\9�@����;�p��]_<n��3�r�#P�U�*�����a��c��5JN�p��\�* -{l��7
����fm�}Z�Q)�*1L,7PU��\A!oLb��g��Ƣ�X���7��6+�m,�`����=�2��2�r�0h���N�|��g���ߪ��#��9"��Z�̏��P<���l�G�Z}��5��0\���g��j�b1()�84�GWm,�8�:P�����A
T���:��H�!#�9f�\IArv4�F�v�D�j]�mᑯ3�/J&������^V�%>W�{f}':�5�n�o*�؛�DR(B�^锎�LL-��(lK���\�ٞ�c��HK֍&VT��]J��Sw��m
qN�� ��2��@�DVr/�¾��|\��ec��S��B�K)Wc���*�F��
�VjT�l7Y�;����co�Z2�p�<sM��zG�$�kZ ��7/�p-s��3�U1Q�aYq�����qLYwD���MU:���v�*/�����h\9���,���v\�qcz»b�ܑ������<(��|��%�uY�ǒ�3�k-��}������g�P�>��b)��gf);�@���۹�*h�;��7W�f�㟠<�� �=�BP�Ȫ��E\�p���S�P#/�`j���b��ss�\�HTK�tDJ�ۊ�d�X�/T�$G^_��U��p�f���Ɍe���w%*��9���su�ߡ��\�����[�r)��+قܘ��z��d���%V�%�W�%R�[����>�-�ٖ��O�m���{)ۛt�f��5���1���y��Ia���Ħ�����_K�}�[���n�wۣK[{�Ɣ}r�g	8wFlV���[�DMӛ2zdeq���]Ӄ�������G�Ce8rw2s�)�re�q��C����z*c��+עMX'�V���li�<��Er.��ʮ�o;z{$�"�jk��:��u��/S����iv�F��lp�y�`p��t;�|o��Vl��{�T�	����[&���Lrڅ|e=�֗�W�����N�F��z^	�zS{���^�S��|~�vW4��n�hs��^�,3yL:S����á�N	7�p�RLB�w��竽�sʫ4���r�g�K�l��
�2�n���r����6�b@�;$F��t���Y����a�0��q<�dG:Q�yL\�DTA�}g�B���TY�r�G��7��GM����,^��/gDJ��Þ���F���ۢ��CI��8��q0#K4kadv�	:%��ɢPy��%P����<�he9��m�T+}�0-9!zw'pY�y�~��Sɣ}J�qPjt�y�rP͸���X�S� {+*H����s��̞oE���O�R&QC3b�����P���)�,C��4�Gp�DuM@M���e�=3�1A������Jp�y=<�[=�=K�}�alM@��WpM{2ʠH+1�rY�$k6��g>>����s�E��Hv�y4�r�]�`֍d�(V]�Y`�����шQ6�)rW4;���ne[[�)��\�%�61w>.�n�9.��O����K���:����k�u�7��/�DR���L�֮�6�[��7����㷺� l&؝�/����,�a߸��u.��u��7�Y��9�A8/�N�Û��֬����2�Ii����֠B���VF��컡l��㌛:�#�'h����Aծܴ͋��O�`��=23��tDƨ�3j�6��<N�EC�렢���eRb��m�k1�����S�<�a�tOT��X>�V9��G�������;�]�W��Q��1˺��.�;�����R�\���o��e�.6Pi̋�uL=R�e�Zz�݃7nw4.������ӿ}p����r�ϴ������Δ���.Ki�:�������t��M������w�.!<fㆁ�(��^R�!�|K�w���-����(N>G=���vF](7.�����f�Lc.�Pp���܎tţ�%���Uy�}��oC��͠\|^�ѫ{L\"�#q�'�������b��,>5����jv��Z��a�y.)8������:�<�q��{+�I{H��tt�/�[��p��O��Üx=�37��Uc��>�0^��9�w�C;gћ�W+c'$x���\�iyɓ�����'jQ��FhR˼�+w�VG1}G��YC0��I�a%��3�×=���w�vb��y9SYP�U=頄s�[�_k��Hh: �F+��~~׎�=���K�\ϧԖ���[��4�KSȬ�\�Ps�M�]�RWv�]}B1�0"Rĩ/�艉cj.Q>�j�0�}2Q\&@�<��e�Y�uP��w��i�{(S�S�.�U�. ; R{��)�o)��.���p�y`�p�luw�v�T89���Q��� ��W�݀�T$�e��7�c������j��辗�<��w��58�t̿oO��U8䤳�ܑ�C����ѿ_������y��J4q�{�Z�T�N�WƝ�ē�4oUu�%&�R��q���k܇������V�C�8�V����5����ڱq�tR��@�k)�9I�U囱�n�}�寯SN���,A�/���U�����U���o�*;[�=��WY�ܮSYY�zW(�QV_����Ď}�qV��f3����]B�_�S����^��@-�{"�z[�Y��<�Y̿
�?p�a{�<���Z��ںk��`��䥯f�71Rc�W:$�Ⲉ���ݢ�r��<�矆���]u�!�]kj[�^��v���5[{k.-WI1ն�}�V����d�=V� ���+r��z���oJ��N��,��r��fu���u�ҞN�kQ��{C��loL���bb�a@�2�јW�
7�Y��U���E���/e�Ӑ�v�<�=�
��_��r;PF�7(;L;C�r�MU浲�J���R�84{3^L.
^�q,o�Xѷ
��5JN�����Swדy�Z�}�?���9�^�C�0��AtE��W��1x�^���Ơme�ea��|�^v�?=Du��e@:����P͊�E�(��r�e�%^��Ѕ�'�#/x9緞�7m(�jZr��՘DT2�(JG7�j먠YVC(m��=D��`ީ�S���CM`�]\)�:�s ��h
��� �3-��_	�^�������CW����b���F��gF
�`��f�Kfǫ���=`�����R\*#�kd_ge�l#k]T��CED�t�����If/�©��S
ˌ�P�ܻ�b�]�&�x��˸���F�����bSJw���+Ph`ڋ�vb�N˛����v�d�����]���7���Oʬv�`�v
@`�p��uwh�^�č��/*F�W�������g6T��z����tu>+��/h�~J�غ��vЎ>���$7���rr�FVv��׼��6y �nkF����wh>�aۜ�>xԓxv�`A��i��-�ӈf�q��׽ln2L� �̪N�ip������w�Xx4���n��t�*�V��-����DSO*�g�,�f�u\B�>@𖗄R*��Z�`��3�@"c#)`k�햠p%p��M�DD����~kF�<
Ft�9�nDM1{T��ePzt���73nq7xtf���+6���ݦ8�C�Ѣ�N�ݗ�+��j�y"3u[>f�kD8���Ư�uש
�	�v���},n�:�\@wӢ�Lq2�G.��Хǻy���Ν�#��S��D�)��8-�5q���Bg��s�U]`ǔ����*�i]KU��#C�q.���$g"� O����1Kd��>�
��{1��S�6��\��n���Mt�Ί2���p�ٽ�}�z�
��nUd�'}�Xf�)�P�4!�A����Tl2�V��t��L�_�Jޜ�9c�i�^�N3�֥¶y!]�S���\���R��}n��-<\�;:�Q����"����9�F���=��F�^S(��(!~0c�T���DT[;��H7��G���|0"���k�%·)�7`c|u��E+�<�9^�x�8§D�Ew�6¨��rW��A�ږ�[<�΁��<{�\k,�,�ڗ������\ts/�Tot��b$�f3c��{$�:Q8�.�f��;��VLI z{/H�Yq�X���b_O�n�,9�q:��^Q�m�D �4�Ӻlg^���/f0�p�LmzrɢP��Ȓ��-�b��ɡ�Nc��7�P�ϲ�
��7U:]KxM��wD����F?��9|�a�����y(yןܫ���;��6_:�e񞅩���5
5�yrLTE�)q�ٖ3rt�,P�8�}�F�/�1����q������P�ʈna�J���VE>b�ƽ�]�7����/���%mo�}�M�Q9��ii��8\���I�zE�Dm9�A��R,þ2{&�K�s2�nQ,���]Mj 6�����K�nos%�9�&c:&�r���ƛ�Ќ��#��X�Ҍ9>���f��BC.&�fF�;Oe���c�>�y;�(f�:�`϶ղm)�x�N����B�m5O|��a:��vU�4���r>��r�u1��k�%����������Z8�)2���*w��-��c�,J�R�N�`��7��M�
�l�F�s"�L,1��啷x���_G��tn����]�6:�_s�J=�G��rJ�`[%fe�x��ؿ� ��Ȳ��>��Xѣ�����j�n�Hf�c�Z��%ҵ�9']��m��v(f��!4[�>"��N�3l�ؕ.��X�2�jEMe�)��:8�Wî�ǵ�z��7��s��]�v�\Jɣ-�������9�b�2Q��)u����$���+y[��O.��O5�Y,�Ca30�֭vs�Q5����� ��`�t+9A�R;�u�������J��2��E�5iԾ�4���2�2^�M�bҭmԬx������V{�o�_G�8�Q�]\�C(���`�ע�ãw7���l�cb���Q)�,y*'	p �_gLG������P`���/��W�Z/�ŰqiU-�r��&����y#�k&����%��1oY!ت�[�ɫ�b;d̧*a�`��f����[k	����k��'���p?��Hl���R�)��i�x8��w�hՐ�#Q:<U'&�J�M��Uݲ����aU��nP
��hc�2dc��:��v���]D��������|^��פJ�����]���Q�O.�V���S��|��ʒ���ԋ2qB����5��(v�3�SE��]S����r�"[�)��8q/3�,�0H!�;�ܹ:���f�ݧt�nu%��1�ց�#u�{V�5�l�Vo'�V�cDQ��)����)N<Xꡭ����Nfm��*W��;�/1j���#7����)J=u,=�&ʾƳE����2tv���Aa����i��A���j���L��ΰY�@o;fP=��뺹My:P�QҦ�+�7�nr|�`��R�r���un[��/gW.����2E2`t�,���-lһ}M�!vmp"�/��}O;8r����Ӓn�Vvq�@�S��ă�<C���ܷ������~TNm+Y�_;yJ�@bKqќ_-�7��H��q''!W:�*pL�B�MrΑ�����A���'�N�ܪ�e��%*V�O�K�o��ŘF)a��)�ϝM|�W�fY��Y�p>b��;st��{f�ZD�ݬ�gVQ�mLmM���i��u�[=���D�K�)�8MY:%1�s��Y�˻ճv�:��>��)�w��C\ѕ�;��.)qLo��}�#2ܪ�G;8�1��]u,����4�uZS��ƋG1�8��9יU��'�ڌOy+�'&�fh՚iH�)�u�..=�؂�]�\L�Z�i��������4t].����K���z������Zu�X�s:��Nvͷ�����{'��[K�T+&��a��;�h1�t�-p���5�kr裉�)�NY	OD���f�g^5I�{��9{�@�OWd����:�''�l��^����;
�2�������.p++j��u�-`�k��W��c��y�����ԃ��/��sP�9rH��.t�B��Kw&�ou.����EEDT��Q��(�,p�QU�)�TX�EZЭDI�Q�e\1�IY�QV1"(�����-�H��U��b�* ���kq�Ը�*��m��X+bƵb1LRTPUAI�b.�����*
�
�L!����QX��,Q�b����KmDm��
��b+����PX*���bR*-J�AY��AQ�X����kPUF�b����%J�qe�D�����ղ�R�*�E(�$EQF���e�DDc�V(�B�QX�������Xb�\Z2�����ҌTZ�ZV�(�1�QU0�b�-�j��*���1+EQG)l�Ŋ��Da�V[AD�q�j��1p��-U�ƥ��*��"�+b*F
�
*(c�{��g��N{��ޛ0ڃ�u�v	�\t�]fmd�����v�vriB<��}ts�«!�`wȜ�����i��,�y��%Ƚ�Y�`�f��Ç�ž�s��3�o�H7П[�T��s�m��p&O
]F�j���yLw]z]�	�z�em�Z|��
�JR�C8�E[��j.'T��/ڙ�6\m0�C}LZ�KN�>�n��\;�b�����r�qBd��٦���pZ�z��F'�ܭ���"�L�P#�Xn#
F��1p��Ƹ�"��pu���6�C��
@'s���n������ѷ�A_�c��G�ϐJ�nҧ�hg��W7�'�
��	�!]{lwU�ݬ��T
]1�1,m\�,�@#�s��(:9���Z�EEt<z��qr��c}&���d�pC�{P`D�)!\M���dLKe��N�.}{fP����H�2q���#p�$xw�@�|��I\�D��@�Oy�"��mT-8�cbԝ&R���*:S��H'��8,(��o#VdAa��D���b��2�v�T��S�E��W����{���#�c���<�򬙚�s��P%����Աqeׄ���gf�v�g�.=��j�4x�m���D�hH��l��`6B��ݛ}a�+GD�b���&w���Uj��h� �)6�6��$p]�6:V��[��7��:�Um�h����P����I���7(��v�L�]�\xh���1]{�ojI��%��R��{��Ny��m������7�E�:fk���p*���8[��������a�
��[m���/�vX�J�^S�����W�y��-�����n�Q��(&����<�����[{gM��f�A�c"J#$�ȷ�aFl�|�u�ϗM���Ʀ�Q��D%���<:�,��}�n)���ٌٸ�C�YT�X�eAg�l�5ZHf������k�R��c�'�*b7֍Ӊ�pk����9K&���Ed�1+n�.��n�tȾ�ب�{�'܎�*�4�xy��wL{:]�n�Hއ��������T^uw&��[`��t��	ч���/���a���Q�
�{&�gd�X�F�T�9ëM1���Yh�����{p�;5T�����o��C��j��>{�c��ʳ¡L�%@�R;�e�T�(Q;�P���Є����BzN<�֜�虥��8�o\��q�0�a�P6#�R:`���]u*���C�P�ZU=�L�ą_Z����]OF{e����	��X�����q^<�m�՚7z�M0������fu�`�q����U�U�yY�v�� Y��)�a��o6�{��v���NR�b�e��`N�u �&��o��K^��B-�[�����I�j�r�ɽ��ܜ����E�s�O]�R瑵�, ���4�� �f[f&��0�Щ��UF%�2�gVr�m�OMig'�<�0Wl�����{�)KEt���|*Ѭ�nٜ���妝`�֊���Gf��X[ӑ.c:�U1�¢㢝C�q�)�����L��������P�<�l���|)JKE�ŏC�e_,^R��gXWl\7$F@l�#(�\w��uܳy�`O]mtD������o>o�*�]��v|��S�\
�T��E�Lz�����3��!`��9#+�U��(ᆀ*�:�nU1��w0�^NY�=3�*پ�ޫ���Ԡ��ـF���p=%�"7�on(5�*@R3�y":��?
������{������ש�tHT�=r��S]���[�����hA�^D���j�H��W�G/0.���c����2zջ�Qe��H�À�]������_��W��(��ۯ9e_Ч)�2X�SL��Q����5q��1�3�]�ѽC�f@���6�3|�|�AJ�}��䯫�`��F�������\ݰ�қ<Ҧ]��]z�C�N��S\��OE��2��a��IE'G��}�4�j�0���U�+RN��'�_&��ବ�����QO�u���H�Ω�<���ɑ��ȱN��yk�n���;���\`��e-�W+}�]SWAU>����oe�[P����+:+��g_��d���n[g�.�=��v���G����ꬁ��d�F)a��S(����;m�sd4c�R��f���9�^�N�|���R�[+�
�2�n����$!��֧����yA�xX�z��b�/��L�"��y�t��厀Y(��(!~0c�X��i��N�2���H��-��v��)��#\�^��b_O�n�,9�'Q�ה`W��(�V��ԳLvW
;����&�L:��kġٲBf������Yn�ap�#е}�R�ۚR��e�J��Da>�����ۘQ�pdlܔ3n�hƪ����E�"��}Ԍ�\ntC3Y�4���)�>�����'���G$�0�o[=�3���T�t�wB�GNǫ�'�NU�.lWz ��|Ӟ���Vz��[,nl�
r���ZQT�՚��F��bgf²�$�5�#i͊E{�Od۩aoN�9��<Ǜ�v�ݏK�+�*9kn$��՝�f bqs����ƣ�E�r�z�`�أ�:������Y��vsč]�yEYm�{kKۆf'5����w��g9�!(���f�_>��͒�>�ep�[v��-"4��ٸ����Fw=Ys6�͓�I��f{�?"��8����s��ఱ��"��z"v�f�ߜa��g�*�"��j�D�zd!o�z��'v�#
���v?r
�Uz(v�Rd�x�:+�U��n��i��\B�9�s�(c���k�%Z��$SȻ�����<L���%�Y~3�1�p��x���Ǩ��b����R^��
�f�d\l��<�P̾4�Qo4��IQ�L-1�On�!�~��U,�0c��.=�~`��j�f�P3���0;��w�Nm'��TtkR�p�T`��==�)��w�.�em�Z|��
��*�Bk��{��[��]��:h�Z,��{(8R�i�k��kt�2��)��w#r#�1h�=�R���b�v��]WƇ:��L���q�#V��A�Ek��5���	��qUV�����>笼�kN�ԅ�W�i/��>�*�hq�E��rw��|��f9\�[gu�5�n���.�N��&+���فIJ%@�.���LKV������aˤ�y��\	�M5�5uk�̖�h��f��FǸ�j�R�W�{�����	���B�;%����.���YN$��N
 ��0Z�+1��S��,xe@˕7�kx��6ԍ]�X�y��]wMgpXV<�N��ט��r���	���w%-L�Df��k=�Z�1�N�L즹gE�
�������q6�Z=���\�X����qϯT�,bxIy�x1���BȽu�\4:��q��%s�u�)S�gAH��x�vU~���f�jv��T�� Ԥl��4�B���0��W�݀��b��X��2X�6B��H�����yj�.v��꥞5{#ff�\�kê�����p��L�����.��KYH3,k��n���DPxxu����c�L��k3ʥg�����G9S��Ig	h�0U,�x��qq��9��{��0���t&��(��9���\�Æ�c�U��^s ��| ���w*۴g��<�
�V�rt�.θ�ol�t:��~AX�)ѫgD�&:��pg&�b�l��D���7�E�ݨ�7�-��)��N{�f�@�W�'����U��=��M�|:x��_q
�����C�G�a�^x����Ѻs��pk��{C��y��ޙUҙz �37�T������S
E�g��3�����ON2������*��p�;�م�Ȏ����R�}�"s����:M��y�{�38�=�)
���4o˴�s�N%�t4���Cr6�m�\���q��p�e7�77�*u�����(^>�b��B1(W>�W�2[��G:�]�][��k)~��K��P�K�������6���9�D3��U�+��z| �<������T��F��7�2÷=�
����نwi��1�7���!c��;"��Ur�"��aa�aAT[ۄ [��1<�b�L�ȫ�\�bUܴ�cU�]�)L�%@�R;�&P��K��ĹDױ��(+��^�7���kz
A�&�F@p9tߵ���ȍ�,WPV��pѮ��=g����k-<������;u�۽)E���ʸz�e�-V�e:�s !0��V����Am���L�������~����dy�YR�vcGl��[KdR��u�H\��I��zx����ا��3�[��i���U
�jhu��N��{5]/(θ�T�r�V\e:���.☒([|�f�s/k����$���MEWW���F���vb�칾,o_��a�EJ�~��(��_d���9	��dq��F3���.S��Q,�58WgS�X�u����E��׹����pM $ ��P�U����y�Xoͅ�����r��+��i�Q�1����4s�S���ݭ�ն�Y�Ku��p���k�{r�g(t�<�[�����n�&,Z�����R��rg#ʃ�[�������6�*�K�,d�Ϟ�'R��'��Md2���G��ve�6�W\�z�K�����joJӽ"�ֻ����{WP!}�ް/Ў��TDK�ۊ֍�x��2B�2�^8�������,<[n�](�<����*d�q��X��Tɸ[��u��	yo�g/O�m̆��|}���72��Zh����C/j��a�*2bѯF�����z*c��ή�2�c�l��r����eƺ����biM2���<q��3�4&{I���z�g��2��`�
��!C�`�[�o�r�3�S�+�d�-�q��O,uĄϫ7��G��z�e��z�]j�&����ꫴ O���h�U5r"� p�Z�Mb�	���\,��z�5B6����pB����Q/zy�5���0�4�!�2�u��M�U�G�wF'�j����=����K/Q=U��v]c����t��f�}KFJ���Y��@@�'L���_H�t���OKꎂ9�!�D�6n	\^�,T^�1t��Dߛ����クσ��I���SYC�d���5�a��s��P���IA����Y��4s��M�4k���e,�;0ip\+5:�V̿6�W:�{kһ�A¹IY��+X!��/2�4�����SP�݀v�c�m��r~,�����\����:���KpdE���Ú(��� D@�]�[̍œz+�J���3m�%�+�[��͙��3�{�ͤ�����*�s#������� )8M�<ٹ(fØs�A���LE��՗;X���T�Py�p��T���DM9������t߆;XO(Y��S�X�g\]�ٚ���z��p��#�Bi�p�����_��*1+]KG�=TƊ��c{$��4oO$��Z��Ez�˂O귣Qt6Pw�"T5Dk4$1�*E�w�Od�:���W��J���x�7��`1¼�/��#�M�0o]8�Pº����.�[8#�S��Oe�oJ�G����g�zd��28^޻�q;�,g���mS%#��W�R����ٯaZ��˰�[~�sg�ʪ����5���Y����c�H���Hs�"ys���y�ؑK��򉕷��r��F��}��h\-��͌���:��x��&.��.�[q���!9<����1p�S<�y��j����[����Տڠ�'���h���pU�;c��ˢ��K��pڧ������#Bv�F�߹s�){ՏG2�2����3�ˏtR����CP#UӨ������r��ۗ�`�cB��F[���km���-�(`�ܬKcZwf�ǟ0��Y�&��pN�ж�Ω�OG] O��.��sU}2[�fB�J�5wC����l�,���һa��J���c�G�)+ПS
]-:���Cn�6�F�m�2�>:�Nfc��<*�.0ICTȎ���ׄs+����99�q<4E����1�Pr �ky,�
�V�e��snB��e��Ḏ��6:RU��<�֮�p�N�WJ|���F]�Q�N_N��W�Y�Q��E�ۗ��}���
nY*�t�dı�T�O��8�Pl]&�8�R��8���)5�.y\�3�=�0"���KG�3b����.2wi \�΄ln��*'gz��6����P8�𓜀h��
���΃]��7]�n(�ݪ�3���(h(8��(�4�,m��B�y���uK��*���I�5VA���}�t���R�GFײ�㰣���1�3Q�}���J�RYظn���X��%L"K�I��۝�|���W�0]ڂ\A�η��q�X߲��̞���1���H�l��s�%���yu��9��HY�����m�g��FY���&����ɡh�=��*"�Yg"χ�þ�o��1*��0���VL�V]�Ji0�u%O��u���+�O�����;x�(�=�jl�_rc.x�#�k�ƦBǮ��u�ʁ}�N���פ}�&K��+�l���5�a�>�{�Y��b+;\�4���\������r���������s�J�b�77y�]oeN�!T�H�]Ιe�X��f����;�8�ͬjb����T�}zNp�\�W���]5ș�%�,���RkU��a.8:l��s�K3xB�����SV����e L�
OP.��͉�q-��<ũ'\9iᚣ���&;�]m���`�E-��F�b���Ⱥò�8&L�_R����E��FN�@y�Y�7B��(4o�Ҵ�ELT.]v�*�R�H���KFvvo��y�B�v�N(�q���~�VG�����T�ǻ���.�}ҎưWe��S��xæ�%j�]���[������inb��΁�r�r��ۭ����v�v�^kc��p�T������F�?]N�+#�^���j���S"�Q�Q�B�mMJq�tH���rp=��F��4�4�²>�@A�Yl��:���h���d��q^�u}�J� rm�۵W���M�Ӽో]��G�^���(�:��d�oJr���Ńn���WD��f>Ļ��=�u/�s�w��b�8�[ݝ+*��ż��8���ݹQ��5�;��K�˾A
�P��s��mn>���F�ŸLoe�S9Ct;T�t��c����s�)/OV�}(��ۘԒ�qG�him���X���y�a��kz����\3YV@6u((pwݜ��b�"�MM�Ċ�. R���e4���ni��7[�ɼF��g/6�n����;�^�@C�=8�#Һ��:�Z;�p���Te{Y���Vc�͘,洋74���Fw�=��\�L�eg.�ˇ �e���E݉v�n�ǭV\.�Z�SF�v*�t���փfwT&^��
�P4�|5R���RY����B���J!��e^��4�\=z+��iZ�b��q�6s�1�$�r6�e���vtߴ���u>B0���
5q�V��X�
�j�3��I�>�|��q�xW1|�'���u����N#�69[��pN��('3L��:��|GvY]>ݻ�-H�X�-�.g�ŷf_;q6��h�szP'WMN�cf�j�*������ly��)�o,��kk����zæw��,��Z���p(thΔ��Kn�.�Y��>�����+zF��Uv�+v��j@H�C#5�y��ܧ��:�j}@Ix[���H	ѕVr��a8
��T͸v֞J����Y��i��gâlV�+C�xc�J�Jw��$�'����{k%?��=�&e�{ݝ%��k�A�B��:u�I��W�ZVݧz��軶�"j�*���--��-�*��kUKLb����(�k�,V1����J*#R��"�����*
 �1Ub���T�DTU1eqhT�DPTH�Q0�Q�h�0�*�*
 ��� �-h*�Em�c�J��#�U�`��	EX�h�Z�J��EkX�++L6V�UV�&-F�Q+%ڊ�X�AbEQDV8K��*�J8�UPűU�,P(��m�)
�QDE("��b��b�mkEV
�EQ�j"��ib�E���"��
"��0ֲQ�(��X���V�Qʠ"*�"֌b�ep�A���,��,Q"!Z�F1�*��
����eH���)���H�U3�#�E[��U�
+L��sq�X���[UF
��~<ǅten	����۝8������N�I.7���{Wp�E���6簵��.�޶­���8�*k���Q��u��w����Cy]�盓���:⟭�,`��אV,O��ƭ�����um�v.3*(�J^�`���@���g��6���\�,���5���0�^(���`h��x�T�ﯟ�Zw� 1	<GK����x���S�0�{\.!�F�!�S���k�sO�n^%�u]��flå0�X�Y�r3����ONG�A�܈yl{T�XN�����g+�e-Y�rvF�t���bP],c�@�a�j�
����5ı�eיv�E׎?f�tXz�`�ro�ظ��Յ��i���Yh����(*���\�u�!�ϕ�jl���s
�c�͗�q1��,"a��e#�e�䡾��D�9B3�*�����E��\Z3"�m0��|��-��@޸טDT2�(�)ɉ��u�P-���֣���;̕��g�ip+�Cγi�R�lVS�G !��h]$�f[2#j7 1S���2�����Q}KM��3�����+ia��*l���| ���t=�� K��^ܸ��}qY�H���f]�otr�oVI������؟m�@5Vb[�Ӏ��l��_ܕ���s�B�e����]�xn�)L�lNJh�wB.Ƀ9�w���Wf?�G�o3����c�0�Zl�w߽��a��z��I<�Ķ9!��7t�}�&��?V��ӵ�Q���G!ٯiA�If/�U1\��N�����������5��tI�Ď&�碔��[��ca��Y�_,^Z</tt�/_��Wbf��I��ͯ��sȉ��?�i��wq��IbԉXn��j�T�*���(]�㈭Z�s�ޘHqe�v��Y<�LU�*�	I�޷+��k��|��-.6kB��;<h�V�ev�/@m��apZgO@#7�.!I���{[QC!�p��HΛ�!f���R��z�:Q�:.�c�۶/e�ɌF
jY<�i�9�F����E-͹��tq㇝x[������^�H�{U��nd���
�uj����F���mr���r�.���ۄ�c'�^�=-r�ʜ��&jP��9��3%��4�GC ta૔�e�v��fÙ�q��n�5���d9s�E`�]��\��5t�x����oe(|�o.���u䱉�	�9�2�f3Z��b��
���6���3��
��nz� p��,�����������ܵE�;��0�k��:����|٭�P���7�( y��y�`=��y2�N��7/dqc#���k�]a煤W^AѩV!�*�O'6���2��.7eN�@��49D:�YJ�/�K���i��t���,X�q�W\�����;�KW���6�Y�ߜƄ8���%�O2Ƴ4aSh�2�u��L&��E��Z�ԥ�d���Qg'I�PX��b�����9���G����� 2Q�q��V:z�sX�����f`���^�]��\^�,^��/gDJn�,9�'Q����]E� )Oz��W�v���h�/Ą��(Ep0�Ƽ��P��!з���<�h�a�r/��J�R<i��j6�O"��칁i���t��ı�`�:NA���$�����U�x;m���p�L5s�Yb8���N�I�����r�V�1����V`a�|Ql2�d�Ϊl7����Pd1}�i�ja��T!*��|Ĭ=u-��0uWs�.c�.�Ty�2���iI1}8&j#)�&:���HK�/�QP��"�=�'�bCwU�T\]���g�xRc�3�Rd�>��&�ω3�Q0s�84�5dh��wC^�HX6���5�j��j���1�8���x�G��E������
7���p��<M+0^-iE�[b6j�q�]o]��!ep��������^���]=��Mf�w�i2�+6��q��n�U�$�/U�[7��+$X���Maݝ��sv=�x�*����A��[	Ys�Y�£[�ד�wK���Ep���u�)�!|�N��+�1�<�O-��A�<wB�m5~s�k�D�Ϛ�nc��Z���j�?$*vu�������К�G����_ql����*���%We,�����s\
�6[!\��Li��e7%��z�6�h�	�Naa�z��N����Ǝ�`�f��Ç�o���WASZ��o@%��*uy���}3�p�\������,qs�xu��c�<�24\Bx��dw7�I���hlFw�VN٧��װ�č≨�<�7H1I�1j]-9�'ٷ�˫�3-uv�E���K��M��3B_-O�	B��]���=ƞJc���ZteU)�U�p���:��V/��mT�
���cn�6:RU�ӣ�}j�p���5�n���=]��Ӝ��jh!�\F��uDc�0*�J�~R�Ș�6�Us< ��;!��S���+/�c8(��פc:�1/S���:哞g*��M$+��R�옖6����%��ٗ��;uwژ�m�pr}n���%+�j����s��Y��:Sk�����AT0�n�ci�0���T��7A�˯��mv\���[>0V����Bln�P�nG8rDos��mm4�J�*.��Y|�r�8�F�9��c���l�%)|f���Z�Gg
����Π=ys��ڶ"@3��b����(��]x;����d�l�WF7��Y�����p��,%�Jp�o3VdAa��w`1eX�#i:ꫳ\Ӎ��
�f腆d�쩑�e����O{��γ���J�%��n���S��R���d��wD�O�S�����l���I��}k3ʥg���g��&��n���ir��Ȝ-���C��>�QfW0��)W���ݫ�A�:s��I�J*WQ �t�^O)h8ԝ/��+[�:h\4�P�'�.�m����9�՘6)��9P+��!�Lf�nxu���Yg�G�>�ۘlI�^siU���.�mv�|rǛʮ�b1���
�]d�<T�n+����mj7U�t��M'ٽ={��0/jV;�Pս�P*�"�Ϲ�T��˧�A����cۙ].�¤i�X�v<�E�ī'�8O���>����9Hy@W ȳ� n0�4�UU=<�(��avd�#1�f��a�ST����Յ���쬠E�D�F�(��j�䚙A{ih��q_	A��]1�[��cb�ۖ���#�)���w����A�����M��L*�n��ZMX����En� �OH���U��aK��W0NW-k.�]׫���_R,��]�1>`�Z�V�z����Q�+�$�,��r�"��C���gIC����	t��8��9�&59���OP��qۤWG������y�h2f�ͬ���Qh����w���O��.��r���#Yb
锎�0���V����j6�i�s�>2��8v��ۍ�=5�HJ�LR�\� C�Y�+ֺ�j)`�R4@
&��ׯ����Gp�f�N����(gō�ن*V��YJ�81�E!����"���H˥�k0�m&fP���ɶ*�;;P{Ӕ���Po������nA���s��JQ6��ʯ���6���)���498���z)� ܋�:�X��i����5�P�����p8�0�7DF@����J��:�&������e���r���*��;G:Ƃ�G.����q���	-�����8a�"%a�^k���߆�V�	.Y�k˽K
����,�*��	I�����Q"���8��c��6�ت�D�8ϩ�b���EE��3P1���p��\����@��g:��u�v܍����4���[�h�O3�8@�D���V2Q��r��S�R�hֺB�G=;��ɵ΄VþL�_E�e�)uF�91k��Yy\��܈<�i	H�s��nJ�sM���)�r-ή:�٫!6kq�4:a0\��cr�Vtc3HW�N^���l�U4m]Jtr��n�4k�z���,Nk�N���qqX3�����٪�ʀ/Z�}��W�5�U=O����?����(���0� q�XZO�!*I�6uqph�����o�^�f�жQ�V����/q^��&�)�څM�O��N�t3h�i�:Fyd�y�O��<39���N3׏���*��\&�B��W;����v��G�.2�u
cBҫ�(.�y�c�MY��j25JǻT�F.�Q[�nf���M���n�)*d�aAe� �E��-9�F�����@(w����IN/(]�c��y� p�Da8�0���$��������.8j����U>��K�Z:�j��Z�n�{�14WFBJ�"�-7�(Eq���hq<�����\�Ioi����ӱ|����49�f�ȨO��"�ז��ʗ�:����p�ĵ�w�Y�@4�u��X]E�
���U1�\�P�J���눚��q)k|-�k�u� �8�=�'7㕠��������U/E7R��zz�<�zm�Ln�|.Y�������4q�os�毢��6�kE�x2;Qx���z��!LuM��Hgf�/x�#��Psa�}�s�^!7��>��GS�Xc[lr�5V{���k[ݑ��v�u4��s���[�&���#aL!�*��Ržb�MIh����|Sz�c�Յe`����V�$E��f�:QP����6(1pT�m���l�H{ʗ�j��s�s��1���,��B^��s�L≃>�v�XA�4Ց��T�F�FE,O�];�5iPp����#i7
̾���ܦ���]YC��'��Ii������<}-(��l�����Z6_�T���.Է�X�f}�QYՆ��H���k���e`0���nR7��{��h\%���g}T�Y��Gk�n�so;3\3��kӡ8n�g9�#��Sݝ��û<��K5W[�-�5ط�*��+Ͻ�܂�V[W���P/�X�Q���RP�GK��m�c��1���#E���t��7�u�`���*.�H���a�u,k(��<�7�Lr�B�SӮ�9�cFn�8�^���wޘT�t�p�)�ȎTţ�&J'�%p<#�Xn0�j-�������I��}��wu�������u�5̓.���\�nz�vp��G����L�n�jyTL~��[77Zs�;��G��6���ы|f$Z뽤��Fcu�X�XZn�ն�n:���lZ�1��3�q�l[Hh�fh�ܾ;-��*< �	��W	�p�(��2��2�˙��jy��Ak/y�g%�ę	4�c�*iLdC1˧\w{ـ�d�'E�*\-����S�cj<;x66��!f[)E�&�?`��U��"��r��g�|����´�%#�11�5b9�We
��jEoPH�����נ�ZXa@Z��\R�-MP6���'�����IЪ�x�U���g8��U:��8���l�c�4Y,X�(V�0���K��ût)��:��AV�J��Ј��8?L�ʜ�6�/n:���N/�l�^H<��tm��[�{Rj�P����y�o� ��������t��R��F-&rd�9ґ�Ӎ�˕�N�T?67b۩膬[�:����J���I�UM�Cu^c���%!DߪuX�^M�bv�U�1=�*�ږ��$zك)�8���mx�=��8�&um2�Qjz�,Ƕ��{]�[�f�Fm�*��sV�jF�f3�u��!�5�1׽W�'S�[SC�Gf񖌭���rm�S�+�lt�;yۥՅ{�P\�61�p)�ȝd�ہ.M'�-%�8�vu���G�3��ƠZ�Hx9}��=��6�fu�s�-Z�E�
�nd|��K�9��=���o�~*z�s�ͥ�=܅{���Lͬ0�b�oij��eƸn���7#�u����r�S1���m>�u��M�2po�����MU������0=�V{�opw�[��,k��œ;)�]���]$�i�m�{�
�R/��z�:��)X��)��j�����8UL�Zh�D���ء�޼�����J�=�(���3C���Tȗd�ݩ�;;!�k�K��r{��r���άv�
8.�3m+�v�wI�]P1�.���U�ڮ��Vj����7�w�y&�n��u���y-�V�O�vه���]��o�/�k����̢���]�E�zu>U��*1�,>�ÅL���=L)��Y��&hj��m��S/��r��.���P��p�Z�*�[�&1���9+�O��Ӭ����J�9���^�qlcs����Yǩ�i�I�]������Mq�ӹ:�v��w�z��R�{}�:��l�O�CA��·v���>Ꚗ���y��҇ȟ�35�Wms4(�%*����k���v�̢m�L�5�
��;[˴���ٵ��1��TS�}��7� *�j�g��4:�h/shHU�\����bt.�X+�,�;fU�b���7�})n1.)���֑����#g�x=nJԯ��+��(Dg���}��+~;x�7%uժ+m� Ȳ�SA/�C�	*`�����}2����s;����kMݬ�C�<R�����U�AH jrW��4J/��8�i�����s�g�N4�5L�:��WM����{n��ʾ�1^���壒�}C'K�ל�_���ץ�}���/]:ˣ[��+y�t�. ì�����w2t/s�]��Iq��#�Wj��N%���.K5���0I��|X�o�7W	�8�
R�h*j�ygT&ޫ\��N�U�����fPf�)Q˓+�u<cۥr���s%��^1l�8�ڔ�;�M��:�kgpG>�n,{���*I%O��2����bm��@;��[dL������\���_Ұw�w1�
��vL�g����έ�(�>?8^��7S���ܝ�=���f�%ŃP܇O[d^V^R"|m'�1և�[�iX���$��1����5��[�o�]a�y���=᧧@��u����o+0�^q�3�:�w�	�©�.1��Nf�t��j���g3d s��+��M+ J���v����M\���j��͏�(�֫���Y��D/��'�%���b#sw/s�g]�ؘ�v�B8H���l�O�Z��w�P_*՛2�S�t�&����ؤB�]ص��q/�T.]���뽧�o;Pܣ����\x�\�Y�q$�����(�u�	e�f�=���#E�5u�\�ՠ�6>���B�w�V���U��c���,��v?����k^���6g0�r��}�!t�q���s���{qV�*Y�K����X���۾�}*&���K�]�pJ�Y|\�y~�xE�ҥ1�R������)v���y��T*mi�;N�8{���N�<[��j�`�1�Z�T����\f���ϭ���0�H<�X#%ԑ�F�*�(Zr㣒���o�ԥ���Ұ�\�r�W=�aW,(���h�&sZ�Z˘6��'6�i��\�	�����h���v�)6����b�trvl7b^�4�s�]���)z�gW&6&�s�X]��M�ଐ�6(q�8��+����,�\�[�hw+�[�ׯerm��FXC���uۮ$���Zb��]�R��<�]ף_Sǉ��[����xrq�k��sU(U-�]��{H̲q>���ݜirֱιm�Ib�עwBڏ���d���Rՠ�n)����s��_R�`��0b*��UeJ1DB"�,UEV"���E�8ZU�(���AES4�J�,�"��
�E�(��*iUA*��Ҩ�Qj���""��W�(� �l*���Q��r�b��U�j*�JŅaUX��E[h��KJ��b,DQ`�je�m@UDQdF*�TAf�1m�EX��YEL�%e��ET���Z*��UQ�,��b1QA���̥��F"*�($jW4�,b�36�"�b()QTPU�fR�a�,��bFEQf[D�����X��EEqK�X��mEF,�%�EX��Q3j��(��
[UJ�Q�Dc�����Je()��bت	P�� �(uy|�nu��w�!�"��.w_=B�Vof�gQ���눭W���S�ۂ4<���<�/t���Ի���f�J]
~�L;���Ǜ��������ۈ��ټ�t����z���;O�&o�ͧ��)!����V-��P�:�B�}YۛH���6��U��pFsqQ���42a햨S�YE�����v�R��69`
�ˉ���R��Ǯ.6��=��UM3�e뉡\�%:x�.�ս`���눼�Kb�m|�mG����k��E(�$��y�L�՝���{8�|�x�,����gg����A��ҵN\�E�e�<�O���S�ȇy����;p�:�@LTD�P'��U�9�s�bǋYԚ��w��:S�o����}�����z��]��Z��^��Q�E�����9y����3��?��z��|����4�K�]]q�:�_7��\;�W8闷r����/�b)���c��_�g$]̩\�T��v;Y��	{��ir_hn�AKT���-n���ڙ5a^��f�Ez*^*�J�X\{5��b�7i7}��0�rܢ}��7�(s̮�'���ycM�ҍ%˵[L���>����O.J��R�ɡP�t�g6��ݻ��9�]��mT�Ћ`������ �~½�Tv(�}����,�]����q�(�Hto�kD+��>�wP^�N{�^F��:ɑ��r�gp���}�q-��y
�혟R�We�YL,���6���H:��vU����ܵ]���UF׷��4:K!kg�U��e���t��R�.��(�[��vuF�ڈ�xJ����T��1���SaWm�諒m�ޤ𧸼���9�g�����}N�����2b�us�.�%R�<����o̅U=ٹ�}U�t�-2g��ROy9���:z8�[4%�s������"&�Y�5ziKt��]W�D�r��Ls��nP~o;E��{;9�dך��U�.�k��k)wn��j�M{Vw+�T�j��r!��u��4�%��
`�"����#N��]a]6���F�"����ï ��o�u�oI:���Y�Z�t]yl� i�D���[఍}ԥv�:�M �j�l��'J�6F�D�ρ�n�2��rٝ��p�]�=��u�R{ܕ2�T݄4��P�2���{����=�OE�ɓ��%(�x�@����jrp�O��.�3�-��5�񥑽<3O^jV�Z}�:Uiqqpg�������=������O2��V'���L����y�;k�?W�k�]�z�״|SX�K������HM'[�����55ԍ3�Ү�9��7�K��Wi/E<����Uf�8�k��V���ڋ��'S+�OԦ�����ZČ��Q稾�\�ؼݫ�k��;�O�h����%���uƸΨ�b&aEDAШr���=�Z}+ڈ���]:�<��f��j}٪�jsq/z�ͩ��b}K���gs���ϱ�v̜L�� �1K��W,���U���#������o+9���3M>�����ak(���o�0�w�T���۟umn�Q��Z���U��j5�:.�Wdߥd�gT[7a�'��F#�������#Y=^v8��YF�]灙��W��qn��#�;5=����Q�ݡܕ�u�'Uh*�*˦�ݎP`-�UL�y�i�=���9�W�4Ɩ���Չö���́4uw%�pԦ[|��xKY���XF��g!�C�IXIjÄ�yU;
�u�#���Я*�T^c�ZO�MRܭ��*�9�l�ed����Ra�H^7u^jŻ�ֈ꼕s�W *Y[�C��j�srv�U����|�z�of���En�:�&p3-�q�g[�Nt����e:�S�W����Z��\�����~,o4�fx��OѭM��p��,r�Tg��G\�{����w��پmMUqink�oy*�)r���h���ި�o4܃�Ev&*3����bo;����q��W\o�!��E�/�1�^Ҷ��kk�=���m~��bB�3��W8�^Ncd4�{��o6�{���#H���3�~��ٮc#*��\�V<�͎�JMc�����f�P�n5�7M	G�qK���8vE.��n��JV�w��k.1)��S��[q˯\gc��l(�O������7g��:��VVw���]�Tn�%T����b�`�5 ��Ȓ�^cLle��p�>���xn��#C�.��q#%X����j��r���w.�r����v�5<v��py��z@W��w|%觼fky؜B�gdC���W3���f3&+f`-��ui��U+Y�oz�V&vt<ZP�xa�X$��|�v�_X�Rۃ&+��V��YG���u�\���S�{4��KxZ��¨oM&8W��Tz�?_<��y>.��9I�C����Q��Wё-�Au�/���/m�K�^���Е��y�=o��QVu��
o�;�ImT�P�c�����Vd�]Z��I5x�����n��&m��ͮ���K^
Ż�qz�Y�C�=ؑuJ�S|�j�J�=n*�^\�'��rǢ����r�Wh� �Y����t7Gc�qn���˚3k�-�(��z�����K������煾�9��w�f�R�pj/)�����VTծ���no��Q&;!5�GPo�#]��Wx���\���J�<��{��H�{B�M�D+h��yaT�����pC�,��1`Sm�7E���k���w�/8
#�!���,L^�b��d�޼�2m�˨�څ�E���=]�,C2h4J]�^d"���U;����+2�W��G/����|�R�K82�G�gj����W�߻�v�ܶ��}��9�盾:�:yB�j2ı�;�Qok79�"�gj-r��Н/zy����i���z��#T��,r��ud��3g�d�:�<꧟mA�OS�mb^un�S�n��֎�=�,�Y�vKԗ"VlM�W��1o��}��W'���ltkG���_s��bb��PU�tg���;}<M(0��7��p{�z��lu��uJyj��/(Ĵ�E2ֈW<���.��
mK~tHV.��-�.��8u�K�����B��bb�h�r�+ȦaG�6\�{N�r ܪ{}n⇋����ܯ����E�l뗵���LdL�m��ׯ�����C'���k�ar���v]c�8x�f�(;v�nr{�\�w����ϱ9ޥ	q��������-�U _D�jj/�ڛ���a������.ӑ�ľ}��zdM]gV�W�W)r��Y�����N����<|4K�r�9����ۊ	�B����X��$Y����Gn|�e<�yaSsv�B�Z��S��n�BQ�Ž9"�ś=�	��ӵ60����L��R�7%l�VU�ȴ������Qk���}oN�]���%�_Hp����ӯu�����k��EN��]�Rvʠ�I�{�f�s��)�D���h�k{']�-?u^x�G�����+��j���L�U������H+����6����K����H�߼�ni��/�c�=ob�3Tǹ�׵6�<�W��澮#�Vٺ�;��Mc�F��q���M��J*���>ޞ�-�i�g�����p���ڱ>���U#ت�:�!Ql�gW����i���p���ف<��Fa]�'�NiTG�Ү�s+MvE.�^�$�����5���9����߹5�����N�:3L��@D<%�T�z{	5�1ߗQ�'��s��S޸o�^�Ψ�b'Ͱ����~	�z�����e��T=�M!!���ڝ��6�h�.t�V����=���������r�N�R�FH�Y��9r��>��N�(Q�-^��o��0�L�c��GX�;щV�P�r�;���n-
�]����:Y�}�g8�XН�w�ۨ3D�'�4_Z�������9��U�9���vژ�B&�0d��2�tƌ�KZu�������泲���s��-W7)Uvm>y�����y��m�gq�OP��r�]r]ףּ����{BV�\�����rk��⟻��5V���oh�nJ���6nßbz�/'��X��j5n"����q%C���W�����p��#H��������ns�]�^p����Q�{K�(�r�j7���+	��wTՋ|VׅR0�2;�\�bw?W8�^��W�36�_ʡ�z.0��i�kk�E�p}.�����i�ۺ�/���.}Y[V�EEۜqs��D,Ƕ��{]�U�7��]���'��ݍ�2�\b�G7n%d���T^5�k��Hr��^6�0aa�rz�̠3}]�o��1��*sx��N�ؘ�[�SdUN�!�Yu�f�{l�J�l;W�K�<�R���f�̺��6*U횩Z�x hf��ٛ�K�4�R�8B�[o�?'���s]"N�{�q��W0��QUۄ+cNw6w�J�U���&G2[�5)p���������!��`�ۈhc:�lW	$�q%o%ۍ�ݵW��ő����W\D�w�O3zb�,���Ks�M���N����mft�8F��n'j�e�Ʒ�@�d�A\6�x�A���Ӷ��(ⷱC��y���F�Q~�5z��n��J�:��S�Ŵ�q)�S�������;E����WF�Y��Y��T3B���f_=����{S�蕬�7�|�������ΚZA��˷��^��?r�K��qkD+Ȯ
b����<�q��E�u�ؾv�ީr��9\uD7�)1�bevYY4V��by��i+��']��\�َ\��o�j@p��2�$��Ό<�\v���mM���Q���3���a�K�[]����V�:�[/�j����Ŗ���
��x�fT^;XNz�9��]�e$2|�ӄ���V�{z$�NYu��#/3 n��w���m^�Z��lk��8�e^�s`�ǫK��#���y��9��#zǧa͚j�w/:�G|]v��Y8%�tL=�MҾ��ٱ|��te.N�@xFK�����:��j�*�ovq�5L����U)�G���QƧ�ITE�U�7ؠ��c�p��ت�r4|�����3H�N6a��/j���M��r����1��U��gj�6�.7-3wu����A�{������{�[�y���Nڧ;iɾ����#=呹����+r|+�e�ݯ'}����id&&��J�=�e��We���ڮ�q�婺�M��=O�!�es�n�����B���~�2�o�y�R�(��a������Ʈ�α>{���ګ�(���o�.��{Z�������q-���y�+�"�;�mjWg0���X����'�q���9���ꂸM�c�����{z�j�@e����z�)iŮt��W���=�ǰ�����t�S~�ܥ�]Ņ�u�r�=����n���YF&!vĢ�,�d���V��=������	!I�$	!I�HIJBH@�~ IO؄��$�$$�	'���$��$�	'�!$ I?�	!I��$�!$ I?<@�$��$�	'�BH@�~IOԄ��$��IO�	!I��IM��$���d�MgJ4�Zf�A@��̟\�+���|�TT@�ک
�)(�
�S-*�l�H�E*�ED�(ֶi*�P!T*�T�����ƨUH�`HZڴ�m�����f��6M�[V���̂�Q�kYZ��ԔYm4@l���SZ�v��kT�-���۬��f���l,��bkk)���ٳt���Yb2J�*���i�m�#j�m�I[4թ ,��kKm�cE�h���6�6�M��6���%�Ĳղ���f�5��V���^��P�V�Y�   ۏ:4�Z��Gjڠv�E�k�-�ۍ+TiuQf�F�v�j�)JU�f�m�+m�ˮU.�;�k��k(�[q�M���Ur���Rh�-f���-��  �4�dlʷ�:������S Ъ�wfn][����@��VP[m4�Ύ� ��Z�Z��;�U�7[�^��
(P��Р�{Q��e��՛U2�V���   {
(P�
 ��w�xP�B�
(hmE�B�
(P�^��
(P�B����
(P�@P�K��B�
��ݱ�]n�᡺�[i�K�5Jf����Q�D�ղ)�JZ��e�   =�+l�Os��B��p2�m6��&)֛j��pt)�*�q�:�:�tp]ݪuևX��ӭ���02�U.t⋰�2F�f�K5mJխ�S6�  ����Jn��)�U�5ݴ F����Z릮����:��X�s�s�n�QBGk�a�
�mv�Z;��骔��`k�٪Ͳ�kZ��M����  {��@����PV��q]i���E�\�(u���ݴЭ�.ҎR�qZ�5em6N��U�ƁM7���WVыVV��e�]Xl�X���  ,( �����뎠T���X�n�d�� 4�ڢ�n�wZ��(V�w���n�����R���jja�j�Z�  �� ҷ��(	Ik��:�n'$
�ջe�v�
P
뻶�l�T�iT�B�( Gv�U
��4�5Y�Zm�U$�Y�  ��0ͪ=�ի��
����R�9��(�2]:8�4�8փ����ˠ�r�v��ӵ`�]ږjʡ&��i�khś,m�   a�J�'�S�p�hi��XnҖ�w';N�B��0
�����V���s����)vɮ���#G��@�9M��٦�S��)H  )���@  2mI� �  "��	J�� �5S����*�~J`  i"&ʩ@ ٪S*s
�F�ÂDR���&k�*+��$t�vJ9�.l�JnE\uA:Ԉc���I���I	!I��HHt���$��	!I�IF ���������l��'���1�L�<p$j���Y)A�3�A�t��M���ږ�Lt�j�{���
��
#6L�����hQ��ζ��ѥxq�x���.֓�e��&	򚊨^�Qf�6��j���"a�)���A6�!��B^a��XM��:�*�J�]�|��X�~�˙AK+Z�5{zf�2P�i��q}�%�4��+��HȾ8vK[&�[UB�7yb�Mh�L���Ztu}�E����cv�=�v�/H�N��,���+n�&��a���z���jJQڣKS�Vd�3\d#w��u�P�_n:�0��*1�U����uw��5ɽx-��� �J��Ԛ��:�J^��6*R�6� %��t��4�km�X����&��ѩBޤ��W3	'sK�����z�x��N���H�Zj��@�S0�6��G��F�Z�e���#5;0]�[�ͳ#Ja�I7��ڒݲq��e&���+5h:Ǻ�nC����C(
{�$�ۈ �X�\B�W>����ϯ��WC�y�]��VI�S�����G�QT�Na��J�8�̬�K�,i�M�(�׻c��k̈́�t�w ��N�1m�nY�E����[�jZ���%:4�-�N����1������JD�֛�ሄ�Y�k�ɠ�}�� �R�C�w��d1���V��9�k1격��P�,Fc�I�^�jH�n��t`���a�d�0�݀��6Si�xTˌ���	fv���u��z�O��bHb��.wB��
��e"�� ���"BQ��7���іD9���P�X���)$�>�8��jݛ4S2g\�¢m���#������F檎ᳩ�J�ax��8F�E��R�S��2�V��"��bI9@(v��N���Z��R��!L�h���@3�ŻCqZ�����Cu"9.��5�5�@e=�Ed.�˛�A�dV^�_ۭnB*��NĚ��+:��
���9<੭U�<��e���GA�g����9���$̉U�b֨��)�̽�8`b��>e�f=jL43>s-%�����j1(Q�)7I�B�Y���6��K� Ƭ
m*T]i���Z�Զ�'�ֳS&'Y��Jv��!@F�8�h�I��B������<���j5Z�TMU�h�7�̠���Z�.��jm^hcHh���ӸI�W�f�C1�6x޻���u�>���T4�in^1Mf��vvKnܰ+`-6���1��7�2�m2J�e^�M��
��Tmi���n��� R]=�ꠔ��٬?�mb[N]b�g2�x�p�j�&i���y��b�	A�6Y�V���%���&EA�޽�h�׎�i]Y�7V�=U�s*�nij�iH�!�V�Xn��1d�oT�/s/d�m$����n�!�(���&4/mm,Nё�\G5����J q�j���m�N��{���˶f�m�wn��A(��-n1�3���2�������Vrh��x����
6t�#����<���9Dj�]<zv<T--"d���\8/h�r�;�6�c�3t:W[1n�@,`SA�GO��1��DةL=:�Z�I�P��������^(�'h�����a	���n9�Uh �:�0Gu1�c��_DL�%]ʽ!<9h'�Ax�4Fm#ov͔^�1��f�X����ݎ+%=���	FB�n:�fや�U�u`fVn�J�t����)�k8.,���q�����54^%u��k6�RMfƃ���Bv1��ޜ����(K�9i�'1�e��v(��,�I�q�n m�o(��\�0ӻ� �{��ٛd7�����)��;�DS��<cPj��[2S���l��]�($��-�ʖj�
�4�D�<��	�!$��0�g�vum:�/���77�XX��X=71�ā�	�q�dÅéM��eX�n;6�b)��)Z�[�9f��˱��Q�s)-���4^m2����(`�U.V	w�C�"�Sǚ���4f̫N�Zފw�Py�f'��Iy��i���S��ʹ�%vvԗ�:��E�$ʼ�ZF$�˗�@��9��P�[v��.�њ�u��&��{��*=�ui�\�	Ӑ�H�l�55c���[�j��z�]��`�JU�]X��X�k[nX;h.3���D5 t5�ͳ*9�ʸX RsL#����i���l٥!4l�Y@�Y�.��ѣ3h̼d��sj	5C�dՈ�Q�,m)J-�`��X��dM����d��нT�0}P-��PL�t�YZ�&f���)ko2�,�-:�C(��fc�SC+���ou�ڒ�lt�5,�؍6�ᎩKj����f���&�R�$yn�殂t �4�h��$3P��)0�`�:�JF,��̕�T�T��l�!�J�*k-Q�����Bc�Ct<1�ia���v\�̛��j�H��V���6 �����&���.�)i�u��nɖ���S4�(�J��� Z���Y�5�c4d���EO�ܭ��t�\D^��+.#kr�[�
����Ne���$�)���yHmgر�j^ZPM�Xj���4�ڀ�Yב���ߝidS;�c,f�2Q�̖6��(�.�����)ˤ��jw�㙰+c
f�CrMu�]�[cn���Y�FE�SX�LfM��N�!=�d� :8��z����lǘ���37r�nʩ��n���2E��o2f�۬k.����Υf��O.�{�*;t��K���n�U�[��0��ӻ�nȤ*���i��"Gh鶥<{�N��Ŧ�Xxh�y���Ʋ���ۥ�VJ�&�d� d�-�Bh���ֲ��"#�h��e�8��n�U�2���,���L�Qe�ķm-Й{`k�&RORi�W3TYT`ǂ��o*���E�rf0��2�s.��/l����lf��A���s,eÚ5$z�@Wn��A8`���o���/Yc����Z��n�ą��Zq1���/M:�$�c�RM�K챊%�f�A�tݘ�u���P5�.|0M��x"5z��������6]Ǫ\Z��G[FU����:Y��Gu&�	�L9x�,���
�ә7-���k!�0�j��d9N�	�f\!Ql��d��R=��P���g���
��vByf��]��X�u�@�a�M͚�NQ�ZpTDe�֔M�� ���J,[.P�����+�Y�sj�ϚP�p+m��q��ap)�E����坱ū�:�A,U�)���Ĉm�wXa�t���+�*Ӌ*��ۀ�H�f��ed�u��aA��Im��Ŗ+V�
�Z�j���/��bkI��2��"�7��b�Q=�TYr�n�R�J��Z�e�`�+HCsv�X�-Twm@�8D���b0��km�B��SF��XF�)�N��I�@������6S)��w(����H�����\�D��6�^�C!��Ʌ��2+�V p���-�-7�3�j���F�6ln�#��+��XW�2���D�G2�"m��E��T�X&$�5��36��;�?�[��㉏�L���@Lģ,��9>o`��r�N=�� 4�����񕗲ڍ3�1A�f!A��mA�a�j��Vv�����Ď<�,��	2�H530�+0=
����
�i����;�����]�r�ͳ�*P:pm�,CG~��K$vT#wEz��7�����'�{}�� ����d��	����#�7T����e�P�݁�f5a�12٩PU�Z�)�5���w�JF��bցdZ�N���@8���o��^���XS�4R�]n;á���gko)��E1�ݷP����t!n��̓{F��P=�-LvC�HYE�e2Żɱ�/FػY����6��M��7��AK���ܘ7�\��do���*�����1*��J	6^#X���A��!֮SSD��Pn��)Š��-H��ѩy�˭eLov�R%z+����V�݆6�|3ņo3F�@�FLh��:�SA�]8��P�N_;sl�o6�B��0�,7����D�\��M��77N@���ݹd��]�q�ON!/`Y�)0 �E���I::��"�M�ܑZ��U�����.*�Q{u���eA�$w��eJ٪��1���u�:�
���<�ݽ�;�!cc�(�]��1H�1M��b��WZ34���r��[Fv�\�t�!�eB��C;���a�j̟a ��f˘����I��*+lϘ!��Ҕ�e��u�*�R�52U��[C�XB�wu��q�*��fJ743\;t.-�![/x*^��@��fշUtZg64[z���Y7�K�GE��Cpm���g� hb۹7Jù#T�B@��`�5kՆ�OE�nP;O�*C��uG�yl�m0%��x)���Xwha38�D��;�t,5&+CEayH���D�Y.��+F�e��)�bq'F�fQ#�8УA��0�6��.堄���v�w\���{Y)ڱ�U�+)}�*�WB���R���%6*�R�V�v3/fV|&m�G�j���ln��7Y{�����ɗ(�VI��_,�4,� ��Ί@�8�[t)��+۔bMId ���V8J�N|&��5����J� ڷ�!�T�SN֑nM��60���)�mh�:���4�u��)Q�!��YT���2��+]��Vٸu�̀`ًd�t����t	��CBYM�8֒S�C&�hXWrl����$�X��Ł��ٳ������E%�*7V�l��s��b�&����r���m�x�$\$�W�I�!�����X�-�Hާ{[:ą��#?V��CjB�kh���+F6����l��,$�.�Ը�� ٬���$^�8sj[�°9{ZQ�˭r���
�QŴ�hL��e�cZV�-�;ɚ�ۤ�څ�^Z�X�ٵ����U1<���ܖ��6�&�*{�^�|K#;�c:�շWz�/d�X�E+�7uJ�j(�#����{&�[���i��Rk����7}d�{�6mm���0�!r;ci�v���R���9e?����`3&S�h���X���hiGn�KAv.��rUأ���!���N��0]��hEu'+}�t!��t�u�-�r��ȴc�ʈ�B{D�����"&��r�@��.�����X<q~��w��&`zA#L\Ƃ�gRz�^��=�SU���7W/�W�m=5�sa��>���m�Ӕ��* ��[�[�5ܴ�xo*k�@4h�r��Ykq,��`8/ �iASr�)��|f0lh�]��,ˤ���Z70K{���feܛ�m�i�����?e�%���YePJ7ZT��i᷀�q�7���X�aZ�{���u{GsQ���H9����ФUl'Ru��z���ۋ^�[]�.a`�Be w)�:�ZF��Ycihnm��$�nkٟ�)��J,�1�̩*c������+1_ת�)�U�;dw-K�L#���E�yV
`�,��H�ʺ�卢PN����F�<�T�L[� �b�QʀD�kNd�*eb�Z���S/&��a�&����A�����BkToCT���vtR����	�!����PW��K��Y	�	����hTh����ڡ*����XNf<"Tt�_$��6�߈�boPᲀ�9��	� �pc��
L֞��\q� ��Ο8�Cyp'y,d4<��	]� ��V#m�ojD%�h;��=�؅�%�(��L��A@Pjkt�-���(iu�P�y�e��:/�蕳k�P՗�����lT���VC4��X����� Y��M�Z�6�1jh�����C�/vb��j�$`*�l�n���e��wFXҵfu��Շ��(�J����؎�D��L0m�ڪ�4wZ[��7��m��f+�%�h��Z�b�����/[\U�3E%�(n^f5������*�}�RV�̓",�X72>L�[�S�R�eޜ��#(�y"[#����b���q�C�W��dm<'"xB�P�H��HWw��sW�.�ձ[r�.�!�#I�"'vtj�X�U�+b���r]�/,jzp ��
�Q�4��n"�(vn���M
t���V+ON�֝Kʖ��Vv*��z�M%f�1����`�x�%���3�f�pM�,�.�b���Բ*Ņ*D1�ý闅I�xj��-�pMVqy�7Z�mÙ ����׊��k8ħV4����F/S��F�����72�toaj(a�h���e��k6a�8�d�IV�á+ ։r�\�-圻ɐK�T�!,'��B�ݬ���*[�CXm"��"d�و�T��+��.���/4��{�1f���jX�F�؁���=���@�ՅK*+u��ۢ����2aX�8U"���:ի���r��*I>�f�ՈmB4mn�T5m�t:���#N�a0�'f����@�˩W�ij��.<sQE,"ԕ�A�ڭ9bXP�A%G{*��1*TF�m/{��d�%�
�e�b3ڠ^)�DB:vQ���0�H�W��V�ܡN�h�f9h��q���\z[�Ɯ��T�W5�Պ�Ͳ�N��j�q��JN6�%�F�Z3)��*]�5��C��;-n�*E* Ƅ0QĚ�.��VŲ�mk���Þq�x>!%9�#���W���f����j� dC4��[XJ�LV60譭�k4?��y�(�'ܚ�h�lf�V�7��Nl��cI�9��p6hr�::��Uz����R���n�P� ��m��
J�w.��,�x�2�wk�+p��m���v��0Gyn%�i�����i����X��t7��6)�\�M��ٛ�
�4@���1�()k��n�%e)���n�X�_; C�R{�Q՗�u[��E���c��/q�ɻ��r�)����垵��N�Y�E���&��cK�ˠ�{�m��+�r�ޫ"�w�E[4����T��.{ɿV��>H�����f���i���l�d�#$����Sp��Ҟ���8X�R�V�O�}�
̥�mF1��S����.��X��⓷h��	�U��s�V9bל��Ʃ��g��A�ZK.����Y�V�,�FI}ώ�U�&��*C\��F���@֜2�U��.æ5����-^��׷�Ez6ͬ�2�U9;j�Vt��W�|#��v�s�����Z0A�!��6�0�-V0L����!2�ڦ��n༫`�I>O/�8zQ_uZ�w�X��Ź����N����Z7�ݥ�jj�$�J�r���7{�k�@��v#�3�h{��85-d�#��5u�-�#�ӣ��w�G'Ju:�Z���w9c���r���7�(��4t�KY���S�ȍ���׹�H[��([WZ�>n��Y �)s�z��+t�WaX��U ��|�H���8�d^]e��
r�Aǵ�H��w���o��#�݃#��^�"T��5�f����̚�2���~q^czu�G�����\�����DFfhq�;|&M����ώ�ZR��uh�T���ݤq2s+�� n�ކ^��˻q�3ʄ�:=2����ɯC��vvi�te��U��j�i�iFO�����҃�6�9o�\zs�w1\���\�{��pĽGS_���/�e�����1����H���E%�|K���1�yod�C������Z�7F��5�fЎ�� lZ�����p�kWM�㝬�6���+�0�ݠ�zvu�\{��9}����k�r�5AE�Õ���t��&��KC���s�;	�՞K��0�.l�%9���2ڜ��>��AS��n�xi�$��PX�09��۔���خ=��M$��ǵz�V>�z���[���H��i������N╍�%Z5���2vN��ged=�$&���VB�wAۺ�qPۆ\��G5͐VrT�P,�.�����^17XEQ��.LZS���ep����7��S�����|Iwno	��>n�R��D�D��E��Y|C�;r�VG�No����L"��=0�HXk3	�|f<�V��5ǃy�!F�#��kԏ[�r�M�X��eif�-�a������%�'7o�v���S&d��
+W�t"\@5`�M��0�V��m��N����&7*����.d���c{�#�/\��a�>�ܵ�v1a�`�����$� +@�;]Ƭ�Μ���=\s/�����>�ʼ7.��66ف��9�sXr�z�k�E�e��Y��a8��[Ff�ZH�n��Wpmѽ�k�Y\_���XB-���]l��<��W(�Xʂt噉h��:���;h�����m�|���)��b�� �{���	�����sB����tEmt����/�5�^�jF�G6�F��mtM�'��>������7q�볂�{���+�&�5�����ْU��wy�K�ɛy����o/n�c�����&j9;u7����Ě�$N�7ԓ� ��ԏP�����x�5�h�+0ݏ#��=,98{�%���3Ʒ�Q׸�:���ͰG���d�R�;;�S=��	%�A=(��ݘ��ɧ�"�fw#ȵ'8�Q�j�:(��ɛ�i~���r��#�.��pdvYiU�Lf�z�h��bwϥ�ʝE��ug�����M���2̽z�uZ��{�L|7�jgJ(�P�8�`�����D�h�
�30n�����=\�9	]�'�|/KO�vJ��w���W�]�[�r�l+��`j��<�@����-�n�q9�,���S'�J�s3�Lp'z�pp��3M�K�y�����qT��*8�7��
���0o��9j`���{�ً�q=�ջ�M�=�u-���!x��>l��h��n��m)Kf]��2U�F�62=��>"F�ju��{eE�r\�Nu݈�D�d���^�Ƭ�\5�ƯBzj��(����;�&2Nj�t�G�$�ze�r^L p�ti�up�6S�e����v��k�E�kl�Y8�S+�I�q��N�Z\���#o#����;�x[��71�x�wުV��;��%O�t&c�V2&�r�3|�Y+:[�r�{:�e�m�1Y�����Y�l-#�quƧ3�}1Ա��Y%Wa�+0�n��7�S�}���)S�f�^��H�6 OnV��.�K��m�x���v��U�&q*E���%�(Gf�;V_3u�Qz���+)���fc݋��UI�8�]��Ӳ��Fe��0B�2P`VZ7�5á���1��_)3��:��}��HblS�p;���;�%�EpulP<{�N�bx5ab>Wn�^yb��c�s�����Y�=y)��{��7.�,��{�}���*k=x�MH�&'��Q`��7y�0[i������f\�A��5���u,e��o��ISo0N���a����p�ʗ�Bz�w]l����]��A���)��U�,��ڪkY�)`�7c�Ƅ�ko��� ��ǳ�K'MTe��ڎ�JB��]s��Ӯ�о]	�(:d�l�oz<=׶\�IQ�&C\�N��.X=�L2�v�O!Ţ��G�R�n_3�ݗ��ܬ�
�MطS�k9�R�2V'�a��+Q� ��_FU5��(�Y��qf�������j
����X��ш�`�Ϣ���nd��Դ�V.u��E85�W:���ݝ40KLx���V�#�2���3|M��U^��$��2z�y	��:y���,��b����Q�'��7z��l�ڑ��|A�W��+L���c��쭬�ɻ��X<L�<|z/��n v���|; b�
�;Y��yض����}r��Țz�pYt+��%�����MG��O/�7A�}sKs�"Z6B���=��+!��"�un<�2P� k���fO�"�h嚇EnE�%i`u�Kr]$�S��B�W/��>G����Y��fa�%_mGr*�=�%��{a�.�m^䐇O5
ӉN#�|� �����*A�'_b��lY(��E\��y۷4Ƈv�ϒ��Ng�^�k�C�qx�TՍ`^�r�>3z�٦��"T8��#.9�:�� ���;G+�鹍�p�@s=��i9��^w[�3�}3����E!����O�-�XI���Pw��`Z��;ji���O(B�ۚ��W�ΫK����t\ˮQχ�ܙ&{r��g�.�y���4Ry�ws
n��0�X{��{I��͝U}L�\�{��BAW�=#OW_�pogI��;�z��g��������� r�<��4^�I�kD�P�t���r�0��+6k5�4}g��PH|\ݘ���垠�yowV9A��/���gs�s�h�����us$[0Z.�l�J���a������>D����*0��F�ȏ��_t�4�]��8D*�r�ZG�WI�.�J��0j�:���
Y�����y�Bh�K��fuR��9* ��O���Dw}�Ĳ���	�Ve[�Ue�OJ��xr����.]�rWv%ئ��θ��;t��qj]N�X�D�'�����J�}p�'���w)������/D�^�ϝ�Jx-<q�-��C%�&��V�[����j�2��O����J�%����g�	�.�D����[��3}L�����5�.��C�hi(޽�~�3�ּ��������w�*J�y��eCO��$5�=��[��sCb���ڰ2��D�4����էʧ��X˚�se��u4��H�=�-��ޝJ3�^�կT�ue𘓕y�N]�K�:.����)�O�O�U��	}���X��WS��M��8�WQ荁���s7)y��<Z�Y��wA���\I�{������O^�������ru����p��&O@��ꆨ��JZ�����0͋����d�F�$��o��YL�N��O��N����zIVxw^�V���Y]h-Yd�˝7e�������
�`G\w�r�+���h������uϺ+P���ZFs�#M�o���Z�jOg`w�{����i>�W�����$�{y����}z��lE��z�f�5}��X�㙷Q z���!|.:	;qv&���b�����/T�6�g�ݦF+O����U`͡�{>�'��,�����`i�Er��K�Z���P��;&���ѧ���p+Yo�Q�.��ܩ�	񳽏2������)�2�,��Ё��(n�s�w���x0
X�H��rD2�{&�X�K�4a9�e;�0�1ƻ������S�a5Z�r�WQqw��Ѕ�[0f��V����p�	(�7ł�w��R$����Uq(^-]V�p3���4�B.�ٵ�#܆�Xu{R���ٍh�p�a��]l���6~�v���R���!y9�.�[��Aї���ܤ�yl,�Z5��j�n��Z�Ĺq]��p��Te�M��zv�VfW�FA��X=Ee����2�y�)t���k@�b>�Ӏ9z�2]�*4OV�PɫY2�Yt(-zW���3�.��Է}�|n����"�ޓ:�N����x��Ĕ;��U> �m����W����Ah��a��:�E+ֲ�D��J�L�\��%t�xW�����M�}6�LX��˛�]x}H>����2bp6��aK,�,�p��̼��=��ɓGV#�>������Eogf�Z�s�3�n,	�Y"��M<FM�z��x6�я�%��.Tį6u���l/�e�FŔn<鶙p|捾���gD�����&B�Ņ���cz`���췳�'�X8��-%w�soZݺ,�|�|q���#�g1 ץR�*���Rj��ö�M���ѡ^{��`��;��ܱ�&��R˫D)�^2�УL��WɎ��I�OMY6:*۩@k[Je��Ëu���6�
�6�q��p3�> ��:��~bv��y�����#��7��;������n�H�7�;�[�
��;4.:#΋*黃�6cK*΃!�z6�E����p�0����X`��앧�٪H��ͮ�r	����A�[�c/��P�N���t�V 7�aJ�2ؠ�o��]�_^S�ȴ�[���g+SU"�Ȝ�<h����<.Z�����o�o�Z�/k�v�����{ ��-�)��&�[��]�C������A��d`g���5���4�&��_Kv͗@=�+;H�z� �9i��gy������vW����ް��솃UzĽ5t�ْ�U�l�g''���j�`<T����i�y>���o�[+Į
�>^F���.�w'���;@��q����f������+�q�R�o��'N��ޚu�
�CH䕏�Tt�2C.C�d�9\YL�\s+p��^��st0�KK��a_\���Z��n'��W.M�^gp5t���b�f�i����i�Tu|2���w5N�d�Q��z�����;3��)�*p`�u�M��1&�PةY&nל-0��* �}��;qXP��Qr�8��nYT�Ch�ӬU%bT�hcl<Of��8��pv�F$�y}Hq�Gr�w'K������f.3J�z�U�,�F�F����,��L59۹���p�����t�>��v�DV�z�&���^�A�7��a�՗��ˮ����*�m�q�c:uam���1A�u�6��v�WC�� �(Dei�#�3���Q5�Ԕ��-N�[��#͹��MPH�~�n��x�֣��@�[S���_d�s�kY|�p�r��j�6mn�g�կV���$�[��byCw�
����=}����	� hf�l��B��F�
ΫlOH���
�˶���?<�S�R��&_����L�R���ѭ0��#��o��X�I�ol�{v�Yp
�eʔ����%�b���\ϑ���yy7���X¬�8�֗X�]nb�&���z#�I��L�z�S�})�Sb�k&�.�L�O��GogV��sz�>�Y��U��2:�i�e(0y\^^t�{�R��
�Y��3�P�N|����;`Τ)6�P�$��l�G�Lq���IH��.��s�oh��F���z\����x�X�~�ڍk��ri���������u��#�/����b��W�F����$k�jƕV��k=���K��8w��q�����:y��ٓ!���2���b���(�W:ӡ˨�O���H�ؾ�PͰWRꙀ�^��`�&���>����ϻ��f�����ͻs�=��2nt�[|�;/+%ٝ�>���M*�}��er��J�)��D֚w�l�F�Ɛm*���*c{Hn99��f֮�ՠ~w�Nf�5���av�F�9Hs�i���y�t�,G��yK�1�R��d���:T�.��J�*�H����xN�I3Tl�ntőq�v�<u.��z��v�j��5�L��I�Y]wM�
ZO,�l�i/O7t:��m]�Z/�k���킌��E�c�`�vW*����+ip�@N��Yn���Ǻ�=�۷4�����	b*�u7ٗ�x�/�E�=>��/+׭���?y�����}��!!�HIOĻu�?OȚ�E��ڤ�nN�Dٛ�:����wgj��	R��V�l�ޮ�;*�6�:�@�p葌X��v0�%��²�r,�b�t��R4)��{-�߶7y���	+��.�����C��V���'���ElM,�6��oQ�a���dw;�gFu��7
#�v�k��0Ґ�D�"�)7[���6T�-��LCr8��Uxd `�}PN[WһTL�K��MSv�iJ&�����yKՆ��HȦ^�la1\��<�[;V�Zh�b��$���ٶ/b^�K>y����h*��N�=���/:�Y���9���+e��N���
������^�i�$s��_�s����F̫�毦k�$,B���3�Q�2����P�Q�ZP"A�1�oA�X�	A���ܜ6Yy�����

AͺM���L0��|�  �'G�Cg4 ���u��O\��vꃢR.AMv�֏y�so�ow�x:F�9��o�eo��9ӻ�j7���'e��]i��E�����m���/����E���U��2�ހ�<���0�[1;�P
Spd&Y�PXmm�D��������+En���fr�U8���{g;��� �����OM�45�If������]l���ձ�)�C���@���D�<q��&�����Vd��8j(�Ϲp�<���ԘZܣ����y�]Jj���u��]�E�jfqwi��S�u��|�oJ����ȼ��>ֺ^���.�fV�c&T�d��M��5'm`��议�X��U_k���gX��c��d����r�mFU�qs����
$�p�˵C(�����Q�J�ƞ����,SQ�,�ڝ��f1Z6�F�p���_�NMꂴ;p1��u��/�;��P�Ry|n���/{n�{Z{�I���ohN�������f);��rN�cvWs�i|m��4�!��=���i����H�qnM���3Zn�j�ӄ&�n����k3��̛8�̷e��m'����J[�j�K[ڙ�s^�D����x^^�l��z�D�������Zj��\(��{a�;6��=kj۬�K;^>�g��;�QZكd����b�[�jJ9�ݙ�_�U�՝�寵�	�;���9��j�{` _v�IF�K��U�L��	j>�ذ����[�v�X5n��)]$��+5:�XW�ך�oqgT�B� ��$��V��b��瘼�~r� ���ʴGi޹fQ"gwwG.��(��B��[�͸-��S��a�/�u����i�(�f�s�#Ѥ�-\d
Ȭ�?*�L�Q�Y�2K���]Y����+~&��Oh'9�u�\�}ˣTb�}�u�_f�yuՑX�tC>=\+{�oo���`n�.7g�`�=<F�2��"��r1R�6y��J2�U9�m�v^-�zJh��=]L�7����Ӽ��7�)�N���@�,�)B�l-u��hD7*��|{�+�r�n�0�f�g��W|������[ID:?P���<�nJ{5l��a��v�nV��72;�%i�`�4�v�pm'$�O4�h�;�QE�3h��+"Q��V�
�2�{3��Y��\���%�]"�X��n����1�`*��p%���b��MJ5��ㄬwK�NAB�U�R��tx�d�4��q���O�l�S�,(nZ���E�m�I�-�s��s/;R�{<r˘,�?���V_!�-"Y�Ҹ4���+�4ʀ�P�+�H��`>뽥���m��6WЎM;�>����*�����>��cu7�U�Ke$B�A�v�rzx�[PRLa��I�q��2�����W��C1_u���=�%4o����� ��u���YCGK�/t�I�ڵ7V��#�_r�m����g��'��:!>ds<�{�^�Y���v䧭l�e�v\�)�㯮S�Au�m��ٶ�K�>�{f�wŕ�nm	]Zu>u�
��(خ�Bj�W�AS=X����<O9W[v2���+��-w�
���$+r����S-����5<u3G�}��η�Y�Q�«e���x	%���vy�;D5$8PW۳'^
�>��웳&�r�}��-/��:�v���[:�$6������'�mb1]5��p�;O�<�[���3%EՀ�ۺT�[�j_m7Ii@�#9�e��k�d#��g�����z�X�v�*_:�<M�������wieHZ:��A ��2���L �2u���]v-�
H�JΉVb���Q�WJ�n���em S�Y.Jی���n�n���'�:���H�3k���g�����]�ʌ�֠�`]*jzӻ�ܘ7m!�
������\+Mu��p��z�q��L��G�Xk崭��p�/�o54�{��t99;7ǏX�[�h=5u�4\mcv�f�=R<F��=u��NvW9�3P�t.�c�P�=㻔4@�F�N١�ŝėXql4��;��p��{���F�a{�-^��i&4�3�@��N��Mb��2[�`�W������1�v�������&_tYټb�+M��z�O��DS�PV��O�+��4�RՉ�2�G8=.����w
}�2�<ڗQ�M�ި�nZ٦٪�z�{{n�w�:�̇�4�U�G�]^ܫ7bS��y�u��9��Mo8�YG@�xB���K�d�p�c��X�v���Sm��8�D��m�/+`�Y�_M�J}�X��1aQޚ���`�B9d6��F��/u���w/v����b��M�c���@3U��6*;��u�T0c�<2�I�˷ß�[���U-H-۫@�B�cU0gK�{�fP��C9��}���f���xOc8Y(:}i8���HeŐ�Վ�o]K�����:��#��*pS�!6[�u�7�٥��B4�R�������Q�w
J8�"	�����B;��5K������]-��u�/GO5r�*q��j���{����v�y�]�'}���x���앋X&<!9��/x�h�t�S�Aգ�����
�u�B����O�R�iʙ��m�+�HM�QW�r�5 >D�״$�底��(�2ͭd�p��ҡ����B-N�U՘5'%��r�����;,��Y/�6��zV�b�}d��x��\�C!�	�����N=�N���2@w$�"���b�3����"�YۂL�hT�*�׬W8h��6��):}czԷ���yiƪ�qJ�3��ڡ�`��s�mt�w���ޮ""���M�?vU�ɑ���aAH��S��3R��8:Μ�͊{2P&u�e���*A}���Պ�"Z���EJ����M�7淚��	6�.%�v���c��n���Q��J�y-��F���w��Y�t���qۄW
H�h�]BR	��}�/c)g	�I�;�+�sW6{ .�ةr�Ν2�P]i�Nn�wN�ŤV��N�\�\�V�����U,��ݎ���Q�Ṛ�hǷ�Q�[�|�W���[��3jV��^���n���/���;�O�c�Eωפ.�h ����qo��1�>��-8��Ys�m���O:Jz��.4�t��ԅc�R�����p͖�33�-�� �Cz��-�;��L;v��?�{(ޘ@�1pvׇ�J�i|�͏:����Sʼȸ�t���~4��0�8��f&7�:�]|!7�)��A����u'��j\�+R�Ch��`��N��[���b˼�5��;tu��-����_+"��Kc���@��J�/���w7��oj�V�ע�{����l�ݬxq�F��x&i/�#ٰdre��/����]ݑu���F�Y�ڛ�i]d�W��\�WNՆQA����5�qX��X�!�-��`ွ�������4��-�m�*�n,�e�� �u01�r�e�2��`�-��`�Λ�<���#w�r)��,Yw��>L��� 8�Ƃl��T{�$>��ׄ'���Vs�ʫ�5R�o{+oҋlF�K9������E��g�6����B��˂7ZYn�`�KN��<�L�Vs�D�U�\
��B#h��[$�˛z�u9:�ۡ}����ռ��R�26��ٓP����?�<�c��t`!t?$h�0+^be5�Yן�����]�z'��%�����@�����wUxbȝ��a�i�y����w��e���3�.�Q#wU�����*X�+���k�� ���|�H&0k���PX�Ō��Y�~*r۸��f�h�,l/���}5k���z�&;ɒ��.���TT�9�(vY5ܯ���{��mP�Id��7�y)%���ِ�"��v�nҶm#	/��W��ZzGN&u��=��:�53dP��.���m�ż�3qa�X[[.|����v�7эAVj�1��U�Y�{�;lfZ������&q�hK�y�r-��Ƈ�;�oh�;�����6��Of0�22����E3�J�������H
�ޮ-���T!�zF���� |>�R�v�8�\lW;�r���c�����X�R��)��9�^������{�]Q����K��1���L���l�N�uNֹ��<i;�)�)�̭&���Q��E>�ts�|�Fo��VN��y�4X}� ;����zە�Pr[�+_{�ˎe/٘<;��NCf�w��a�I��md�|&��L<4�8���n�Ł�B��t3��ţ N\HW���>�Q��e�	H�xtp���о�mI�2�;t���ފ�8��
�f�f?���=��M}��L�Wu�1�YX��a�C%�t١Ď���;�]��M]��>G!L864)�vq��������>!��X�����V�ü3�!u��{��9.��O�!0;�iP���}͸#�;�����]�Oh���x4��Y<��`��a��u�H��@s�{�5R���A�u�A�_g �г�n�[�h�;�l�o3B:裄��֫��L�ˡzV�'9�5�JUϨ����]J�vu�k8T��1����ٷ���I��I���N�[jLu���P���#{1
f��/�W�6��ˀtסo�fk���Y�R��� ���d\�'��m>Q��c��н鑈�XT!uz&m� �B�1�c�%Jj�s)��R�,k��=���0��kϣq��(�՗"��$Voo���K�=�3�gأQ�r���_��-�}9I¢4�ZG��-���*M�Xx�L)�s��K�����ک�X��@�z���N�f��H2GYw��jeH�l�yI�9#�N﹌v�j����#n�ks��p�v�Z�Se�i�ۢ�a�á(��T��p�t��pr>̓�.F-lI�3t�u���*�<�F)srN�X%�_R�*�iN޲TY}Xl�����s��l����ׇ�����݃����u��uVS粷Mfr&&c�u���P=<Xt��{�gg-ki	��&��Z[b�ʊ���D=�D���q)iW,�iZ�(���>�ŉ�|�ۧ�_��|,=����T�w$2�ra�u���Wj�gD�Yuc�v�.*��Ў�Uc��nL��+���Me��얌6!`�-`S5ԣO�+���ib�������ZwUr��h �p�/a�_��wΧ�#5����-B��
�>��U˓o�����f�g�gUj�P�tm�ٗ�u\�K���� 9k�+��V��լ3�w[��.���Z�M���l�S�{ZȰ��ʚ�-=y�GX:�ٲ�oZ����b�d�+{L��rX��b�y���l�K�\{b�
����3��<�XR�	����p6;�pܠ���2xfa�-&'�|��b���v��(P�k�y�� ���D�U��4ޖ�>%�ح\սOL��,���Ĺ^�a�Xn��>rL��������Er!|FRٻ��kyrTZ���IjC�@�g"-t|L齯t�:��*p:���w�=V���y֗��j�\���i����M�QTI��nSwsQ�3���ބ�9z�1�.)p41>�u����]w��r��J��V%�|o��FO��j�q^�N�scBވ�jt�wVVm�@]Zv����_��T��.Ϋj�Y�$�''vE=��rH�׈k��ً��T���smjq��񵸅mf9�WN1�3�W>�XK6�25��J	�ΰ��hk�*R���WT{\��y���g'cL�T�4���H�����G5�0�#��e�$i�C�k�,�nt�����]4�iU^=�}�I>9�m��Â�zl�.g�4��*S���H@P=彈�чL_ws6�Q��a�2Umu�V�t����ٛ0�;��=��L>�:��(:���~�6�\���Օ+i��;���#���Rv�2�ۘ�e��i���qy)�#d��bh2M��9(�Z]l#�=��n�~,.�o\�W�_S<��ܓ�!�/������9@��M���gs�:NC�]��g�7��,�i���Gb��J�����b�-�M@�� �>�n6�1�r~wP�Po��'��]Z0�l�
zmX�BJ�(���R���Q /t徭�L���F;kY=��<2,�ګX'���ă[��7���h2^\��C�)T�u�b�,d�өe�3I免�P�]�eox�ڨ;�n�q$���v�1��:]�^�t53�{�vr5<[��T�^��l��Zj�b<���̚A!�d�L�H�����Tի�����ڊ��崏tGh>2�Γ�0ÚH�\���������`�t�R4�j�{eh�d�ד	D��R5�F��ǒ� zy�E��j��,S{ K<�2���,����Z\�v�O�����+�M�5[$�M�i�㺸X}�n^�6RɈ�{a٘O_*�|Z��A:�wV�{v�킃����C��pQ�k�����5��Z]*�nQ��[�
�M�[Į����複m�6��<����yV��J|J#����0���'�d����-+χR4��E���W^>e���j���K���X��`�3s������g�Խ[�	�-�$�:�21��󯶾͢�><YLy�s#���~���s!�2e<��bI�R�PB��`%��tw;R�C:V�;��{��v]�aov�x;��t$�麢���i$0��b�*H�>M�z�W�9���ۏ�� m_l#�����&`d�e�˽�O;$��kxu'��uBy��`��7�2U��3��p_f<ƫ�n�
��}��-�Щ�f�h���VޛYgjkR�&��9�H8'���M�[�'+�����ae:YZv�朣n�(s.]f9|62D�̩��mb��Q1���7w�m�ɗ'Z:L�W�y�S��X�ޕУo&\#��:�X�U쬤,���䝡E�\CY�{���2��g(x�bD���vB�f�W����d�3�eҧ�\��,�a�+'.�ſ9�o�<�˯� �B@��}��F$JE�*���lKJ�ܴUm��m�,[mU��X�-mmc�+eJ���Q֖��A�h[E�-�Qh�Z��Kkij�ne�aDK[B�)Zխ�����lU+PU���h�j��m��*V��F֫ѪR�X�����X����ZʈQ�ҬT�m�)E@��JDaF��"�*4F��f0̵E�6�k*V�YR���R�Zֈ���j�DTR��1m�B����+��1B�-�jUE�V�ձ,E*--Y*�bR�6�D��(6��Z��J����cQ����%KER�lT�F��m�R�Kl��D��"��ѥ�E��&Zմ�(���1 ��eD��P�Fm(�2ն���Q��R��R��Р�%�������m�ѥ��"��B�EmiJ�FҌ�*+(ĵb2�ڵclU��l��R�-B�R���ƭm�(,cmT��m�-�ZхVTb��*�#e�`��|/�r���c��ow�>��U��S�g���ޒ�5���%�i���v��}�nJE�^���� ��6~�*?�k/�O�,M�f�c(d!�©|�R���ۨ�^�[�V�N�Dn1k�ğj�y9kr�q�F�^�O���ߥW��p\iF��{
�i��˷�<�C�fv�����>v����セ% �r���!'�S��r,M�~=!S�����a�m]V����5lHҤO]���d��q�R�FE6y�|�i�6Ȳ�/�7�C�%fz�{9tB��K�	":̖m`��τqn�s��7YPlE|z	E�����I��Jj���d��کzc����\,}��^����bp�j��]�=��SX�^�����;� ǾIT������A�6zS��:�ui��>��>�J������z��U��#���q+��x`(؞K�.��bU�>
����¤ܾ��TY��*5���l����ҧx:���>K�O~kO]*�����cOk��IHR�����ӗM�Um���;ӄ5��yW�&�5YA�Uk��s DFǼldzxo��a2rS����b���Q�������l��y��Z�'��x�/o&�/.p��,3�D~��5�d^��к7��jpQg���`�6y���z��+�tؑ��|�Q=W.�n�ԓ�DN��T��S�+^�F�iqu �:rb�8՞��f�YY�s�ī�Nha��DOx[�3M������=q�WM#�v��Z�]�T`'�ҁ�C�퀉T��
N;p7u�{<��e]�8��W�7O�y�ym�C�May[W�9P��"�t:�=�O�����~7���Gy��|��H�ۛ�F%{~�鏦VC���JKE��<2�����=9>5��u}�+�t�k�̗�\fM�#��l���*,�iD���6q�(�R��'��^�J�t��������X�ܽAy�;Bz5D�z��s,�������&k�Qˀ����������63����[�w�4�*����UdGX�]Ě��WJs�噡�!e@�
�W�[��4^v�����M�
2
����(dR�Q�E)�/G*��uY0�2dhWH�fIdWtD��Foi�Q������,�2j'ٓ����a���ԍ��O7|p7u��{#�2x*�W'u�ͭ�I�F^�0K�4�o�YZu�̛�t��:�J��zk#��]f��N�����ƠK*���s�@��_v�f��9ݺ,톎^*� ��Z;;�-b�n��ҁN���e.0P�r�:p�+ܓ��(%�A��7%���f�W���{0��k�� �[�^XP^����zx�7���z��;�Y�������9��i5Ȃf:� �5�I{��eqyk���@/y4��{r�j��9��"a�T���p�A�1��t.��(D	ط�"}v�Mxi@�]����%�vᬚ,t�k�f����1������3�F��G��j/]냃�x^�r�-��_�2X22,WuaV�.$�� ����;�}G�HQ�aw���s��Y����C=�>�!�2��H�%׹_޾��V?e��Z/Q�}9��>Х�����v4��vE���.����=���|��������{����O/sՏ>�<fG~:���4�������S��#KB�V	� ;kWY���'^1o���`�ߝ���+���=1N#�*��΃YZ!ZNC�v �3�I�{=}+=�za����>tv�����D9;7�Q���^�S�*�U׀؞�&�^�*3*뉍�xa#�OA�<rrF�p;ڦ���N PnQ���^�J���]A��J:����C��+̤�+JuqZ]�5��*t�w�  J�W�����U���p~2 ���s�����w�w����y�I`��������O������Wf.�ɡןW���sW�{";@Jښe»Z�2r���Jk�>�܂�ϴ�j�}S�����H��\���qeƾ
��"4�'Y0�	2��f|{1+�]M���x!Π��P�Ixr�W�*�ʀ����ҍ��]؎I��T2��S��\i����*��S�y�X}��޺���H�amz��%�vxL� �#��{����ǭJ��K�U�����(.�Ks�l'���"�k%�P6)*�i3^� �[�U�7f׼j�}������^�mێLs�O�&y@v� ssb�T2��u=��^�����y�J��� Ժ-3�n�s�GtP:eC�R�:����@�PNsO��7j�if�koi�뼟N�rg]lrT�u�L1�}�����n,h�(��L5��pM�'Y�"%�N�s��mF�6����^��J�j|7!�w�����p��PQ��>�����9]}Qm�o�[}�W��bU���q��V	�UZv��H�2����>��(8�S���Nr�-Ju]�ѹt��٥p�t�Ĕ�2o�V�!�J]o���A?y�mu~{�e���OD(H�e'�F�4!�9#I����޺X3UzY3�1���>�)��`�+A,oH(��d�y�+j3J��\y���]Ȟ����NX��Y�tfܜ:n�&�v,#�������*%dq����i�f�u;�S
-�ge�$O�n�SuG�aG&�s�)�f���?e烫�kY�U�U��:�d��T��Kڸ�X:J��`�R�o�d<�8U��F+�tr��p��{&ѫ�ۍ��h�-�w���t���2%�*=��z�S��3Nr��0Ʒ\a��Q��#3�bn�g]�:�̩r5�՟��q�)�MFtZ�~��:�j sr)�y�VVh݉���!&_GЮ��_��穨|3�p.�{ ЙD	�t�V��6��A(���J���d�.�ދ�)�˗{��d����0g�;��F/eW�"Q�n�����r��g�`N[�Ri�l���;�/5�B��Qy9s�G��5��9&��zB/���1���ױ|3�J�*8�.5�#J�t�hn�f}�$�UJ2)�A�:1GT�]ÒN{������6Nz�S�0�#�}�(��u���3bV��TE���G�E_'��CM�Y��u���H�T&�i�PѲ�d���Zj���q@o��KA;�A�>g���M��zg0Mθ�7[�������<�産�7��At)�w�T�jم��J��9�/jv�A��ܢ����R�+e ���oe%�-ͤ7gi��L,���6�s�N��U4��?�v�mR�V��[���{��7��4�,z�Up�b�_��Ҝ���i������#��5�[1�/f���՞��`�	4���u�@������K�|��no�6;��Vu*T�Z�F{�Y�f���s�ҧ�DX�%^�x��H��H��n�z�s-ƣ+��L��Q'�(�p�)�Jp��34U�Is����������,�HO�e�c;u][�{Js�L!�Ta~ʜP���͆KUV[	�:sϤlD۝3�lVjKK���d��������{!�ש
��č��p�).(lJR��S�Ɩ�p��������:��8�ݰ�^fƴ<��tL��{��Ȯ���`�}^u����V�>�c�Q&;;E������÷Ȉ���FM�W�H��W��ʔ���ip���Zzr����ב����Ǭ�է.�~T�H�(�����U��@����J�&��\\�U���"u�lC3'{+ի��c��,����V:�R�Ɂ�@�$b�}���J\�1`o��ok��{:���cKm��8�Mht���]��rr�Qy^ܤ%�ۢ�����4&љ3�.I)�A���ួ���pW\/�����-�ԿH�A��Q�.̹�]L�BRl�/���"��\m��x��]f٦�M�륊�]�x�aCw�T�'�>�Ǳ}��i�kD�S��
�Ӫ�#�zwh,Ut�!�3��r���y\�4���./?mΫ)��S�Z*��;
})�{�<~��nџq�aS�����l�"q�K{z�3Jx�8X�W�MD���w��6Y���F�T�w�wZ��Ym�}+s{��ut�2���F�^��ߠ��FM�t�+`�Q^�C}������lo��G��t=k��=��2���IVk�  �x�����w	�%��k�x�F�'�D;��	7=/�����tR�ŵ0pLP�]�b����n2��S&���-�]b��	��{ ;�)��M:IR��3M�h4SE�����S�N�Eזߨ5:Z�R%:�y&JSdaB꓊6d�d��;�
P!ĝy������;״�*���]�1O{����ype�d��=�>���1��K����yu;O=tVϊK�(����W�M��͋G�E������7=�\%�Un�W��҂��4�BO�t�͚]�Ћ�7�ʑ�AQ�\4�Meu�+&����'Z���YM���@��sjo&\�����2��(��{��1r�b�W�,�w:dĨ|�y����
�|s,�"GԂ�U�sÒD�4������X�(����Yt�gy�D{|�u<����iy�}����4B�]�S��S�Sz�e`����W=w�׶����s�����*��N�b�����F8�p^T+�/κ��9遇�+Bq3^�p������2�9�\gTy�n�Y�:���D9;<���?���B�9�����i��է��$���"�OCq��P���*q��m�9u���7�OXZ.']�fk��.DU_�VZ:%9��ԫ��R�=�G�P�ߵ�!�>Z浌E�d���HGV�q���p���tP���=:Q�s�������GYw��F:��3����^���8J�?�U�"Y�P'aT΂&2Q����t��R�o6�d*q�N���bl�����KȠe)�u3^� �[ڠr$\#F�-�WD�k���U��L�4}��%�u��5S)�v� P��E�E��-�ji�V�������ѯM�N-Q�1�^ȧF� J}$�oSY��	� �Ι��ZYF�:����W�U޴��+�є���i�֔��S6��&Ɨ���ש�Q��.4����Z�d~FW��noq��$��g�e��u�i�y˗d��--֤�@��
���/X��w4�l��C���eq��(�S&	X��v�,����}��O����W�<u�o�3(�� w�L)99`���q*]5&p�>/����'g"�Y�Y�>Ka�S�;Y�ƛ�9f\1�0QGeϣ���V�^���o�7�'ۙ�!G�L�N�S�m�V�̔p��n�gMHȢ���TXR�[�in��/�Y�����r�K�պ�G)u���O�z%��0��jgչXf{�p��'��]���x@�����~����Q�3�T^5��2��9o|g�V��ve�j���5�np�2x��,J�"��á�]0�ԌP�k��;#
Դ���������{$�C�
�8�Xh_IQ��%C�����N�4��8�B�c�7h��PH��|q��Y�5%u
���#2Fߺ�ϨDq�Yp
C��ޙǦ���ω���>*%`�o���n"�-���=���0��Y�=��U'�C�Ϟe����λ�׳򱶪6Vu�L}�����g� �)��X�0tgz}<̰]�U��hQ�pm���W� �χ���A3��6��E�3e�%hC�p)��v��×n���q9��yEDM����V*FT�H����An��荱^����A���q�Uf��IksX�dKTit�%B��������{0_���}�x�;������n�
=9��*�7$�,=��*c��P�C��E��]%�¿l�p+�% �cC�%�$���`�t/j�W��]5���PG&0���i�K�TΠ�^̋��}J��F*#�T��s���aI�(m�b�����	"h̖m��28��:���ڃqE�c�x�c�����Ԯ�N������T��ʄׯi�h���}:g}=LP8�`[N�{{2][޻���&X�4����%W#�^<|��d��C`����\]lkL.S���j�e�*9��c�D@�
�11���'���bS��o�-��c�$�kN�:8��`���5���Ҝ�:C�l6h\���e�[0�4�{"��ڢ��Ӫ��y���lq���(�n
s�/.���ʼ�4��F����:I�
��oHf]�m��\��)��e�a���E�P43e�+�.�sC��lD׭֙�ج<R�b�bmOe���xa��K��^�lV:�VP�P8k��*���
S�Ɩ�p�UT
���[�+x���_ͮ�='rD'9�t1V�x�/�ۗ��]W�j�2慄>����Ȏ�Չ�gt��Ө�\�F���\�#����$����� ��-b.��wJ"�����c�qY��fv%�����K��������!�ۤ)�Aye��AZ䝃ϙ���|.����3�D x�Nm֣m��ĥ:e����U�9�V��Z�$��M���)��T��F'�+����
���^��&�60X�q<=\n���)+i�e�g<�,w�[�P4Z[��s�t\�
�k�TLx�q�n��ϊ|"��'n�.��F�7��0�/ ^�����o�`u�����O*���I��h�=O���liT�e{�vK�,�.+��#�G˳vh %�����G����ilQ�u!���;^���2�O�=P!]3zQ��ܥ���\������_����Y�$L��ޢ�{�8�K�F��M��f��m�S����q���Xqc:6Y��U�3Qb�d�|li��E�svo�hF�4jvɒ5��s�8�`D]-�p�n�t�P�������]B�9[�Y���G�c�ξ��ᲿYʼį@q�8ۂ����SY���vT9E�WϨ]8��z(,v��nL����w"Kq\tv�D�g��x=��LT?d�k6��%���e�߶���0Z����*�ySE�}|xJy�5�/�bݦ�a�KI��3L{������B�1a&Л$u�3�n��+�#߀���uj$��eqf��lX�Sk`��(��3��E�t����Ru(�Y3+Q�7%gu-��b"=��O�P����	74��V�}�6��3��=`2g��H���CVht<ӏu��9J��(vs���ÆU�	󽡲��5�]�i���εq�6i�9��f�-Ǯb�kd�i����Y�����h������^�4�7�a9gG��Ye�����Y��r���ST`7��n�E��P	�]���I����̪��8xS��P[EA�I�75m�����zґ��Z�N�4;�IҤF�ӽ�
8��9Z��&�f��r�id�^j7��H���KG�+hF�`�|S��b0r}�+��6u�R$��7-X�մwjf�����l�̐ث���NYZ����Kt�J����Lac���P#Ľ'����jN'��o.��M�*9�_
��ȋ ۝�*cA����ט'e#�-{G�����<�%d��D���WX�u"�p��X�cV����T�.�+��Ν&�3��'0�>��T����%��Gˍ5��Ž�/�;�B��._��L��Ze���ɚ�D2�1BNº��"EZ��\��u˘0Bz�bv�/�n��R��3Լb:5���;�6�n���/wb<�^���AFqOuj��U���_O�Ʈ�V9Ft�W`]KR�����)�@�v���L���}emQ�Tm,�X1}�.-���Kh�R1JR��TTUb1ml�`����ŢV,cmZ�mUkUkPb�-,VR���5�������[Fآ���R�[Dej	R�j�*�֥��,�6�$Q�E-��e���A�)lIZ���eb�%KV���
2�Ub(6۔+�kZ�Q�ZTD�Ҋ
�VĴK`�IX������F*�-E��DIT�,YmH�j�UEQFF�֊T�[E(Ѵ(�ZQ��"��E[iU*��k6�R5(%T-kiU��R�Q����J�f&E��+m�V5�b�TE-R��[H��R�U��ejTZ�j1����%�ʨTQ�*���b��5�\��F�Vҋm��!R���iQ��TB�E���"�[X��E-�*�)V�D"��(�*�ҵ(�h)l�E��%��
�##��!�����;�	�M
�w����ם� ЩҔͫc�k�����h\�mk�g�eF]K�鰞G�d׵ ��3�a	P�[ް平�T��RB�;��.�ۥW�2Q����i#�
oP�~
�Gm�� ʀ�RJ�۝��Wt�":�w�K����=��;�:/Ҵ_��K���ei����w��N�W�<�K�\Ep�MXx�ޑa�쀑���U��(�R��ܩ�h[�1����ON���}�Eu)[��~�`}���;���Z�s,���(D��I��U�T�����&�Q:�'+�rd!�c�豑j7U8[S��5VDu�wib��8!�3[>��skQ�\5&.��@�	�V��n��F��q�2�H�3��s��g��g�|_Z�-b�g=��{ۻ�<z�����٪�����<�h�dà�L)��C2/�1g����JPuV��P,oH�#�3�H�k�0��.�Q�~�t�ҧ�	u#-e�y���\��Z�Q���:�3��.���� ���Q��$�f��  T=��i�cV�V[���ŝg=}�y�襱���~PL�*TcS�̺r�q"�[�B #��eWY��������{咭�lAa��r�H0+R�:�+f�R�̬F�pY�8i�|�u��=m��"��i��ws`�o<�=�$��B�2�ٽx���^�5�n�#^Ʉ����gt|'�p�'\#Zz�� �Y�o�7�M�%ѵi��2��غ��ӷ��āY[��E�%��d�7@ah��k1y�\� h����̉{��2�ц���Ⴛ�nˇ[��|t+hk�U�Xz�B�*�P�4W�+)�Wk�Z�/1�+~�c
�l���Wo놺���$�^W�k˩�ltaUӡ�t�\ϧg�;�ә[���s�Oɒ{V����OzWF�C��puq�}2�x��N���D�ٻ�E_j�V�/�V��u�
a�j����;>�+n�\/$t��k%nͳ�M�lQ�+U���s��R�"��LPp�-���\B���x�T�-<mX�����sQ�{���+e�8׵O�&핎�l<�A㓳~�(�<�>�B���[M'+QJ�<}S]*2,�/k�JK��Ũ�SGqK��N,)U���[��RB��~�������~�4��q�ؠ/��2�qQN5��}�����Ѯ�c�,Ol�"�3���t�����ăMfa6�hB�|5`�2y�7O�v^񻝖�BF`0�f�XsC���O*�u>���4cQ�cN����Mw{�"�T�7̂	�j�*�a]uۦ������-tށ�O_u�&�]�d�Q�M����D��VΘ�yq�&R�rC��!�x���x�3+�f��4�[p'r$S�lyۗGԙ+s�h�S����"Y��gA!Y{׆���9ָ�;���cp��.8�Y^��X)d���*�i3^�hI�Ǖ@�YFNj��stB��+���L��\���1�L��76*5\�"�
F����9zO rsc�U�����s�'nLC��&�r+�FTo���^�&gz�*���	�b@��:f�����֊�Yy�o�s�@J�i�3�]^���\)\�q��P =�`���WT����g��K���<yf`��;����=:v�b����zhd���pŎꂊ֨-2ĭ��������:;V���> ����"��`���c�|0K~����ǖfq���*sq�eU����t�j\b�ܪ��պ�7K��7�3M��W�O1[���Ki�jcp�U�|��.��mW�a���u��T��B}��C#�.�o1�[RM��}[K������b�K�dO��P=y?ⷥ�)R�mL����;1�ϩ��p6�_	��h��K�9�`Wk&��A^��t-c�>�Dp5�o�ګ���;��%E��Xh_&��,bT�j�dZP4:'�KB{"���Ί���4��^F�Oq�}7"7Ֆ��[�#y������U�*�����{U�垺2F�#�L�V'W٘KW��;;�S��Y[4�j���کCºθV	�=�RT;��Ӡ�9\qB�ce!��J���Kg����?n�ҍ�j�:8>C�|+C��+ӳϝ_N̨Q�z���s���#��T�{������3�����E�	�U��烕>����E0+��~��z��G�֘~(�O���J���������g�~.�0�t0����tO��o;o0�N�U���S�Q�tr�a_�C��Q'.b��(��$�
g����D�"z��+��
6H�
�Ʋ�Q��i\�.�=���ȿqG�a��ԣ�7';�R�4�N��2�"!W��Zs�Y�v�'���K�:=�������2 �{�x잎gy�F�>�� 8=ɓ",���1�|����b�զ�z�>�|�`��F&�7�Y������'	�]l�4���	�p�T���Lɯ_Z�W���BL�>�g����Ʀ)�Tr,D ��$�{�׃�Q�=7��';��K�y�I\�=F�z߬�^#�d��p:��k
;o'"�,#��YH�� �t���T���k��|�]r��:�>W�Q#�Ӝ�/�ύ����1w_��Sz9ۋA��y��I붰Dm�C2�RU�r�t�M��{�E� p���83Äy�x�.�k�l�a���-�B��	�"�(�>��[1A���E�<�N��"����j�]����dFlc٢��m�pl�H����WkU�GWI<D���T�=��|��)��Q�K�u�h]KW�@�l�]�w��,�xj�[S��<��Q�:ån��>���О��"T�/��6+�X<:���p���hS�Ɩ�˸]��6�=[�v^g=�>����G�y�(��\{M �v�(��"�%a����u������:��жC9z.J�]��PR'�ugE���2e>G�A�R��nP�z�w�W�nQY�XY�N��쀭D��l)�ޔe()�8ʜ$��-DdS��L�EzLixĄz�ϟEj�=b�=X�N9�v`"8�^��	��WS�I��GG��X��ȭ}v$R���fq��V=�_wj�������MR��9fSX�NfXx�^Kw��V��C]�eY�/*lr�OK��0R�nǟ��<~����VSz�=Ǘy���r���y]�Ѹ��fUݿ��x�p�޽*v��Eۓd��;q�7D=/�c��1=�i���=5���9� �<���:Eb��ۦQ�s,�����C��j���ӲwU�����r���4�-w.�����+.�$����A�#*Q��Q�Y���Bd�N�v\�cF�"���u#FY)&��Y�4�X!>�}����\���AHf	Re���ⲑ�B��<J�]2�t�R��ݕ�]mI�ra����!�N��i5�DP:���@X&I�%��qʢ��K�qp�����9�q�	���nm�3#� �,\[S�st.�,W^��nQF*u.yY���l��;j�׎�p0�n2�J�K���3M�Z13��s��w�;��f_j�q#s�W���N(�2P3�b��
��K�5�(A����Y�v�SSZ�Ok��^`�� ��b� ���K�o�Q��Axu4Q.����![FNf���lt���|ja���_�ş�x&��[Ϛ��Ox�YCj��oW��o�'��*��L�P���H��ob{�q
�N�U��TŹM�c�YX0��[e-�$�`�Z���:��2@RN�达� ����R�"���pJ�vE�]Vt���`B�IGv״T���*��#8ᕱ}</�e&��U�3�M��ݒH���UBwSq/�9Mڰ�MWes/����ã��Pւ�kP��m�FdV�w��f�P��%W8n��>��UC�מ�������z:0ͨp�C����M�:o7f�����9���7Q�bY�?^����<ߓv��:���D��MN޼T>�.i���rj��2���u����	��`�%Cq�ص��h�T�p�8�9u�p"T��/��1��v�F��~�� :�xdP��S��TZ�VS/�u�օ�r�pz��g�L�RL�*��ل�ޑFz�t�ІH(�Xv�W.���=:Q��\�|rL�����;�N[��Ĭ�}<C�5]���4h'>�ޑ,�(��4b2Q��T��}s<Y�W�zl^m�J�v��«���.���u�C���(�A)��,2v1� �]F>�X��1C��j;8��8l�!N8��3��UC�t�n�\����
�
��H���H&8[����ӫ��Օ�Dp�k�4.E8���}�����Lu繉8�L��B"������a<Ňr��ev:�
^�D��DMeSqz"J 8���vai\�#N�Č���\]�[Tz�	�D��$5'a����|*t�{1X�~�u��
�,�R�Q/z���"YR������9.�-YW���*a��o^��y�@�g��w������(}k�l�cӾ&�̤ewY��!3�8�<���}:n��RH���݊g���Ŏ�x�"(�H�_lDh��)Z�cv���A�2r�I���w
�{�x+ũl_�"�1Xu}��YO�{�Y��'��"<6��*�$:ݟ���Dݽh5w[2�VD)-�G�tQA�taK��fn��T%׶��C*�[�n��ǩ���kpmn2�d�ev6�A݄��9�\8a������F���g�ζ���];��Q�λ����qU���`�,�2Q.+zX"�*F#N6��>�ck��n�y��x��!WH��/h�z�]�p���%Ǩb����Bݧa�r��ƷN]��P�>�ܝ]�!塴�1w��5��F��ڮ���������������Ϧ�&�	�'9*�O��̮��Q�B��2�Exϓ�P�3
�{ ЙD
���T�R��������?q��S��ϷE������h�=����fx
x�0���o0+P�of_0���[1�����4�b�N�-6���,�D�I˘zD#���!���5��1�������i�D�ojX�5_{�i\�.}*����g��O�T�!���}7���C����+��s�~�k`��z*�iUh�|.�h���iVP��<$�;�}���HѵRv2�^�� ��x�ɘv�}o)5t����_����2V�v��!����;՜���t'B����H�Ը�]]A}��UO�]b���kS�.)uy$di�j7#��θ�H��,۩�-�,C��T�4֗����u��}PXG���(߃W���Iؑ|�M��̽�x� �O��{�\�}��#�Ń�mE��"ɖ��	����P�,�����8P=���ee�z��](-%��C	�*'��3b��`�,�}	4ߺ�x0Q�<��]I���mb��{�;��A��Ua��Nxٓ��-�B�7Ht6`L���>�
ي���-6�o	����C�l�D��#L�y^��q��(ۖ��u�R��ɫ�5��Ȇ����'�����P���r:2Cr��c*(q��԰E�P4l�]���	�:p�6"e^�i�R�Y^���=^œ���xaݭ9˼�,�<�M�AgC�~[��W�*�t��=
'������oT�T�3�_��5p6.��t���vT�m�1�d�����b�S�Mo�:���%�	�"O��?��,<Y9��޿\��}����Agx��h:�E �ϳ�C��=N!�=���X��x�$>��B����&�Y�k���h����m���'髦0�z��|=�@�8�P繣�{����9�o�~ƶj���)P�f�ւ�v�,�[�^�Ov�cb	�k�W��|�^���g���:�(0�ɉ�ܞ�ˏ~�P_�C:p꼒���V�]=�"���Ns�q�E��Zd�ٽ��kcp�$�&�fw;�����0V�ea�{������{�w�9�����	G�S����$��'S�+�!Xm�2���C�R8���_~J�'�̊|���r�~�bc?N��H}l3�T�qRT��i��T�G��O�8�|���^4��:l}���ɦ[g}�I�0�<���,���I���E:�����$�
�%�\�B��>=�M�2z�Ձ�u�gY+��YE<f ��a�y��I�޾�f��U���Kr�ގ�
$�R��w�5����x��XjVkd6�C�b���,8�gW���RW��Nd�@QC���}q|��s+:��kWg=����޷R���ׯ˰�E]�ӫA���߇���T���UR
~@��w�Y�ă�<;�o�,����V� �lS�
�C�M0�1S�c9�?Y+m8�7Cim'Sg��l��$� ��]2wp]W(˝iJ�Z��0�9�!�ه�6������
��l9ܻ��Y�J��0PQ0*q7�M$�o,���Mr��<a��O��R
y��?:IԨ��§���'����"��<v~����[qhL��9��s�M3�IRw�b,�2��C��
N�Y1����l8¡�QA�O-�eA@QM�kˤ�I�*o�']v��zC�Q�{�'��l�$Y>���9�'~�Y+�M�6}�AO�Mg�Vm ���ua�P?}�;��YY�3þh"�ƥu��aS�CfP�Xz�g�WI
MU����M�\�Ȭ��,�3���L����Oy�ӷ��o��4�2y��}t°��';�<�Y*i���6��S�Y��mćy�W�i1�}ܓ��x�k��!PH>�ݳr���>n{��HG�O����1�7`g�JŚ��:�iZM����g�i�N�����P�����Ri�aP�4s�N�k�I7�6�����x�1&�1�s�'x|�}\����b��µ��9��a��>�#�O�s)5�O�|�O�Qf2T�'�0��ΡR�5M0�l1!�ɤ�⤬׶�'YS��Ͼ��OP��O!�c�:Ɍ4¨I_/�.=����{}�������'}�bs�'�8b�	�>�9-�8sN>	����++����wys=:�:񊬼=��u7���=�n\�I����E<�]�O�R�}�=1�Tr�������{�����3���q�.�F.Pb��m�MMޱ-�U+��I]we�nL$:H�2P49@Dau�2U��[�BɛR����k�������tc�e�����;t�z[���dQkV7�T�.� X91V�Y��d�ch!��RYJ���4�x���þo��ɔ{��`Ǳ%��!�Wv�<�c���N���,LkN!���-�-�	u��Rg�-�.�N|�yE[o��C�3{�Z�S��.�V�=��**����=y��x/����8�^M"�kC]�8=�;�İ�ѻ<2�y�,j�H\�'xD&��v�yC��R1���TD({�r��u� z�YOn嘁�Ŏm:�N�R�Df��iV�m��G�yQ۹W��\�u���܊Y����f='r�[��j�6����H��ܮ��L�n�V>��ßC \թ��r��2f�w�{�I�H�1�Pӏ,ෳ���ׯ^=�{c����{}ke�A�D�q1�l��Y�Qt�:��j�Vrg�b娖��f<>M{�|1��D/p1��"��	۾C��T�$��m�Ђ�{|�맦��/�u� �}�aj&-̶T3MЧ.��n���Vlѩ�c��Ȕ� F��flA�gr@tEH�X��n��Y�;;����=�O]����"�b��p<r��;�����ا��Ye��e����n޳J���>o�ch��^�_k�.��q��ݫ�T���i��0D�Nu��]�G�G={p�+(���@��P8�d�~#�,�Ǧk�9�{Sj��:e.�1��oN���E[�&��4��H�;�oL<���)�|4�lއ'��Fl�3�������Cxh��z�Q��<4VQ�`J�4�Vӹ�W_��&{�����W���@���w�0��!��-�Y���D&Z͇�������\�>�mm��d��$�Q�ͦ-v��s���;ouPrq#0�]�^<�{�e��ɹ*8+ol�K�>6����u@[���Z�m�9ʸ�:�P<�Ա,ܮ�[��*1�����EPvǤ����Mۢn�G���c+u3BfZ��ԔW�ۇ��պR%�/_N�|��g8"8'J@�8-�GJ�Whgl�+/y�L�uk[%]x��V5Mxs����9�w�]�E��&��eq,��ݗ�(d���:�
�ܗ���Xt)ī����;���^˵;FE�{�EBq�-�WZ�a�e�Y���g;m]�Iڦ��RW�����-U� ^��9�'6���1ݮY�Ƹ�&�]�OX��phRww��B{P6�SO&P��}���Wuo�o�0����{�w�_-[b�Q�Ŗ�"PYkJ����mm�[T��R�`��A����e�X���mQZ��c(�QV�j֭�2�g��mmDVЫ"�[QR��QX�iZ5���V�"X��mT��6�(+l�U��aiQ��� ��eb�����kFѶ�kQڪ���Rڈ-V���1�4���JZ6խQDcZ1F�Qe�����-Xe,QT`�Z�`���E�J�(�[h��R��DV�ZTR�5R�lU��F1�)�m�4Ec���U� ��EPUQRV�R��TE"V�-TE�JV�D�QJ�P�YX�V1F5��%�
V�X�lQ�*���-���\�@EQ��V2"�[-��r�-bڥ��ZTZ�1V��b�p�TZ��J!EQ��\J���1DUDAf\���TV���V��4�+DU�J+2�(��R�-�0��TKJ*%�eE�U`Ŋ#-�X�Q+TJ�J�"-c��Q��,AR�eш�

%h�1��ʭJֈ�"����%h�ek���pmv�Yԟd<a37Q:_(��qҳt�qf���_w%�V^A��Q�+����7�Z�5s���.�UDyl������ D�wr)Ѭ�� �b=��?~�mE+}���
���XVO��!S�wy>a��OS����g̕��s�w�H)��0�VT�ힲwVT*E[�egS~��Q�>�.�sIGE���~@�|?{�m�a�z��1�ل|���f��������0�{�jzɈ
)���1ӤC��0���Osy'��L?0��&�;�6Ag*x{�&�R
z�e����D�gj"}��0�l��$2>FP;�g��x�Φx;�e �_��P�x��*)=��O~f!��=��
A��X�9�
x�im';�CL���xwxiaS��<7v��+�g��r�گ'��Tv� i���{���X�!��f�PQz�����Rm��}�C�o�B��\�P�=C�P=��i�I�i*>��O�1�l�`�B��7���}�0:���;�a�+�6 Da$z�*,�2����a4��VM�̚�u�|����N �C�M��4���f�w���
���w�i�O�v�����|d�{�?}̓L�%q�_�}��~���ʺ�CRWW�5 ��H�=�Ԃz������ya�Y欟j����ߝ���S|�%gbu������Xq�"��x�I���,���L@^��$�� by���u�_s��|�=�[��}�>d�{��fB��
�CG߲_��8���w�UT��o,�>Ag�0�j�9HW�oϰ�C�H.���h~B��vLM��1��N�m �d��^_�k�����{���i����>G�����|@��ud�<�p4�����r٤�B��?gr�(�T��p�?n�g��rAAE��yE8�Ri�jO̼�+<�Owt�!̤������?e�|�����^���O\I�]R��'zs�z�H<�������s�j���ڰ�n�Y1�;��
M$��,��̘É�՚I��3�jq��(����{�;��רW[Tn�o!ym�`��3$2 �ᤐ��'��SL>a_�<N��4C�%z���C�(��'{��'�ʁ�{��H{�T+��27`cY]���(��9�J�+?0�����sv+�c��3�/���等a�7}�t`��0�����Zα��50��"��E�.����wv� �GmFa�v�����:yOj�&�{G�Զ]<R��غ{(���彗����{�ӛ@.޾���_c�}C��8��h�R��N�=F� ��\v��x{���cO�7�8¤7hl3�&�'1�TP�%q��w��Vu�y�<���0��oZ�w��u��{��i*�A���:����q�<�z�����$�ϻ�� Y��u���sw��tS��@���g�?&!�
��
����=��8�����Ym:��������Qa�*w�o���VM�ɾ�@�8��"D��Ɉ>��!cJ���]U���� ���n�I���t��.쟙{HW�Z���Rz�2�����?8�g��H��M��`�B�_Y4�a��b�m���� �O��4�h�e���o���r���H��&���f���c��B���5?w%՘�P��kEd��u��Z����O�v��݆�~a_̛=�yH,��_=�I����&	8��#��08��8W��W}�^T[c�' x{�+;?}�He�8�w�g���r;J��14��;̞$l1��(���Zjw�
M?�L��s�ɤP���=a���O�V~d��sD)����k����FUW�P{{<�퟽�a�3�14���t���@��q���d~�+�xs��u<Hn�y}���S��y�H)�f'~��!������X�i�1�Z�OwI�>ۏx�)��v�f���E� $,1�N��������Q@�=g��u'r���̘����s��6� T������=e�@���l=a�Ri���2��1�5�0SH���m��Dʌy�*I�.�)�aW�&ρ>�X<�P6����biܠi+??�����&���I�RT�!��N2�:ɉ���0�N��jÚ����5�
u�����tN!������pz�ev��|R���W���>��pS̤~a���Y<�)�u� lI겠�~�<�?������`ny��+:� (���q�Vq�'Y��H;��}���u�Hs�������i��PM�O�y�u�_��d�w��i?$�?3���N!Y�>�;��8¾]`�}�y9��x���ٔ1>@��6gr��
�|�Y��C�C��&3l>LC��ރw%������YB���-�E!���5�����Z�g ���=9�>�Ƒ;��p��p�Wi�	����h�,�Z���cG��1gp��J�tU�0�d����q�4�|���iv�i�k&�@��
cG��< ����Ī�|{�$3�.�C��bA�?�w!�,�:�y�d>�'�Vk�9l�AaX~9���P1'P��]°��P+\�T>I�Zɉ��%AH���@�|�X����˭~>��Mw�1jqU�����=�>��� I�����כ�q'|>̇P�>M�܇ό��w&�@�1��C��ͤ>�J���U&���O�IRu��2m��[g�L	<��Ϳ�{�a�����{�Agl�3�[����qh�����z��j~�Ԭ'���6�h>�'�&+C�`#�H�`�=�}��S)�I��V|7;����p^2��1!��Z�Z�����^`|���솑gXT�i�P�%z�d�g�C���x�5dR~B���P�}������x��Z�
�G�ޒ(��IPN_E�>�X�)��F^�O��M ���Qv�{`l���PY�bC��j���<LC_~�i ��n�&���C��X��1<@�):�f�Nya���L�}�N���> Fd.~X>��k��(�����
p
g}��m�7�����Vu����9�����
��2!��'�^���M0�?e&��`st��$����N�R
~?8�x�C��&Z�w�j
���a����s����� Y:�z�T� �r�����"�����2z�l��y��:¤�r���d��ֲM'��8�C��$�
��l������W~}�x��Y��e?�����梬���!�IO��Y��Ld�,ĨI�M���9���uP�C��ɜ��Vz�2xr�`xԬ�>�1C��y��h��+�2������H(zG��v6^O�P�ﾷԻ�T�����B����<��B�������N�Y��J�d��>�1*N&���L��Aݓ�s&ޠ����{�T�Ͱ�bn_�RT��gyE�C�id��Y�t����5��FR*7�Ώz����0Hyi<B��y���Aa��N�?'���ayE���x�Hu'r��9ܓl��PS�PǬ
�d��si<Cܲi�t��0���e9���0�LV	��~�n��]�ƥJz���v,�a�B�W^K�=�c�����O}��pճ:��/AN�	��뙙��у�Q�h�p����	�B{�]�=�^���u��,P�#���b��)�C1���xJ�a��f��<=��=Z���tV���"�x� ~ڒ�'�QHjg�h�����*b����9�ć���S�IP��d�eN"��g�~CL�e�u�s�z¤�xs�kt���̕כ��}��T_v}Y�B��[���	��d�#��&�|�M!�s"��B���t�&�Z��Y�&?2y�Pĕ=@�N?�3&��Cs:�8�T����q�Vua�����J�3~~����g��.��]Ǫoua�0��	#���_�a�,�³��oT=I]'�|w�P�h�m������d���Cû�0�<d�氞���q���W�T���*zo�:� �C����j�G[����W�ǉd|���}�eA�a�����*)?}��f!�qa�5���JŘ�3Ý�ć֓HW}��M�(�g5��I��I�g|�m��/�,��a�
��;�5�{�ɵXB��1���zO��#�A� (��*|��bM!ܲ~J�R��s)�y��9� ���w��ğ�����ȧ̞��x����~�bc7;�Xm!���5̕4�*J�����K�5C��c������E�H��<d��ٳ��&�u�I�����$��t���d����I�>O���ṳ+�g�ɷ�OS��=�L�%2k(���O�(�Ͽy��|]���mv�d}
-�I>dx�lz*<4�!������YY�f0��4Ԭ�d6�C�b���,8�gWLeRW�ߎd�@QC����}q|�3�Y�O3XB���v��;�Z�ߏ��%���&��4�a�>��HOH���J�a���U �4s���~q �N� ��?&0�V� �l7y���
�Cs��l:�C�ug��&~�V,�q�t6���u߻��Νڷ��V��~}�=� A?oH|m=���a�+�������q�CL79ܻ��Y�J�s��f�4����~���!Xm���O��R
x���J���=�W�*��ġ_vBxA}�2|	D��4�~�m3a�ڇܰ�!����r&��RT��LE��T�(~9��B�c-���a���T��γ�((
)�&o��q��t�N��UG�cn���r,˾�o�~]�5䆠�H�9��z�5�oe<|+]�)�Y����w9h�BȐo`vٚWۚ�ˀfNԍ�MDD��w6	�y�O��z��M��-4dNi]KU��P��Xh�i�]���-@,ы�j���&��rE���hg'���y�P< ���2m9�'���VJ��yM��AO�M�U�H<��^d;�U
���û�?5��C;�`cR���?!�1&��n���8�~�׎]�1W�U�|�	������$�A�;�̘�����Nߐ1&�=�L�'�́�+
�d�u�P++%Lg��j�8�r�&��,�ć�y����Lf��I��<Oqy�o�_dڈ�N��/��J��"�@�	 D@$�f!��{7`g�JŚ<���5i6^`Vo�L@]��a�;�>~��0��)��&�V�G?d+4�g{�AAE��Sϼ3��[�>��q*�$O�#�@������R��p���>C�Hy3Z��'�$��{5d���ny��*A������$7o��i+8�+5=��Y:ʝE6}��z�d�{��!@����#��,�zϽ'���dRl��Ԛ@QJß��L@�=C��z+'٬�������2z�Շ��c>d�̛=�z���l<фⲤl�퓻��Rs��9���|׿���'�T���ȏ������ A08�g�f��'�~C�wa�E�~�Hyhc�����������*M;t��g)�g̞f�O��4��
Ͳo��͐Y�J�������~<�vt�,�l�ܢw�ȒH�$i��	#,���HW�,�3����H,���8�!�
�N}Cl=f!���No �d�]s�����3��LI����,6§��wg�9k����o��9�ox��+0��}�L:¡�>�wv�+8��b

/�u��
�h}���23R�}�sT�!�P?C�a�q'I�����!���f��/��O��L���͞�?]�a�)�?B>��'�}�*��A��%}Փd��>O-&$�
ɾٖβc�z�N �C��׌�@QN����i�
��;��N2~s���dς>t��GTzy}���וU{�㟾3��vLg+�v{�GtR
|�|���eH=�9�������}�ֲ�������4��a��:�>���Ì1����?3�y>��}� H�=�i�1_Mi��Gvj˺�X�cA�Z�2��ę ��l�v3��m_U/��^�C�4uc.4*�c�;S�VN�f��MS'S��x�i�N��{�	��Yox�B#���	�o6nԕ<1�Y�&WfP�]e qѮ�:抲�k�{O�����j�z�d�����G���$ �����&��s2��+1N~�~�,�'����ĕU ��%O�Y�1��!]�����m!��~Sl>M��
�<ݓl8�C�r����vb�ٮ��שu�rz�l|�f=�'��gɌ1!�����=Փ��p4�����y9�6��V���[E��
�9�'�����y5܆�PQ}d�QN T�A�2O̼� �k_Պf&2�_a\�nt�0�+�� vRvyC�'IԾoH)���ܡ�P��>����x��XbO9���x��VNw6��Ɍ������T=/2,��̘É�Y���m ��]�������wGGѰk�i���	��d��� V��bz��9@��i��+�'��zy�ϙ+�ٮ�=�AO���ؓ�e@�=�]�=���,j�Ʋ��*@QI|o�?x���q+�?{;�Y;�����
���������&����
�ݡ��	���Ld�ERWO7=��Y�M�p����0��oZ�w��u��bi%UH?w�i<Af�g�9��I�pL��Ĺ����������b�{5�
m!�@�>�L�Ɉ~B���������a�6�udߚȳi��ߵ�N�Y�Y1�,+
�ퟧ�IP�4�?}�}��Xq��������M�%�KG�aS|3��2M �����Ci�
�����~e�!_5����'�s,��&3�O�$��p�)1�A�ٶ�*A���i��!���������ӿl\���k��>ݯ�H �O�|5M��(ߗ*=>�l�"~Rv�z�zv�\i��ߴ{�r�%�#�gd��P�x�B��;.}A���5mXȯ:�2e蝘sM9�9�T[�ZԪ���uQ�R:X��c�t����Xq|�KJQㆲ$�jE�W���!Q��+}\@���bh5��ݶ����.���<��Z���^h,Z�G�Q7ꆬ��{l���єmI�8���H���ݫp-�3�E��	��SY��WW<����.r�f�նVǜ@{"\·�7��Շ�r���r�5k�|O\��xx{����)���X#K�?<�[^��}�檮u���r���|�W�!W��m����W.TR��b�P�@lQ�+&���>�ܔK�ޖJ���yud���x�'LZ����;o�L[ԌW��������]]+l�`s����!������ ��e]�T��]����W�z�΍�c���1A�Q�#�B�����4#��AW��Tw�{�"���˗�3b���*ε:�t-Î�2�Ex�0����<
����� gq^��v�$\8�5��O���j�Qşwc�h'.�yEq�^\D�[��;M�׈�f�e�x����a���V�+���k�ws�k��
�C�! �	˘���f���cK���˩ː�O�1
�q�j�ߏHF��q�\4�ip����^̇	I}C���ԹVWWLq��Գ!p��ب��lL���:���$OUv�'���Y���oI�}��<6��|N(��*��s��6"�>�B�Q�5{z^ԝ���4/i�PѲ#i:s��O`��ay=���Fd��y��=�Ƌv��x�UvkgB�v�:=��N*sh����Ή�l�c`��je��˚��[�T}!�U�Q}�G0�&F�J:Os��kV.��`��%�WQj;���G�|�o�M���`���Ю��x =�:�"���9�T�T�@��P9�bp�j��vcK53#.ś�c�d�T<��6:w���S��܅1��l8H�D�1H���� V�i��S�
6'��^�jcvy��ނ�mVͺf��f��6d�A*Gd�`%Lt_�fELQ�}6����\b���uj�70�9,��0ᛷ^��N7 ٢�چ��N��]!���3l�1H��ܿoW�Mk3�7W�¦����ax���:=�A�h1̦�k�W��1!u����P��z���Ua)����S���ZU�Ai�jR6)W�$me��).&�@jm�qۮ��]Q;׬h�i���]8�in��y����1	�Tx'�9�]3��P���=���O��=2z�K*m?e:��Ohq���Qj;�L�֝��)�������3��]����}t���fz3��q�=Y5Ѷ q��+	ˬ#��	��\k�^sV+���M�̣�w3����k���Ѝ+�|�5G�N ����e���T�7w�ջ�:,N�[#8���fD5�����ƔHϚhά�P.�N�<[�Y�ي
�)��!R�so'
ו�RAlnя�%��kTn�����M�x\��K���1`~�)doq�|,c�N"�Q�.���/���W�|VM��Ɉ����^#ho�]�U"v.`Q3\��*��\#jǽ|��U��Z�nW��$��;[����=y��>^	���RT������T������q�2�;��t^��ừJ���:�B�e�SQ�����E�27���4K5�����\$�����n���I�S�bz��Hc�06c'��9���,��!�&UF���v �;�7[�J�����d�[L��Sc`�Q�i��(+)�|�i5Ȃf:�=0.�H� ��P��dyO۷f��>4ӊ�u��L�6���ʀAC�	�B��J�=���>�"v��s���4�����J�惡��Ղ=�p�հK^Z�Y=���hm�M$e���uZ=�`M�׺���wM��e�!�2�Q�d�p�X��r��G4�5ծS��3�e�>��o�.$�Y�����߶���Ɣ���$4fݿ��]@e��2��S�ARy�B��E�w_����67��	y4ctr=CY����"���E��?<�;
y�n��h=�x���[l>��P�B�֪j�o��΅�����cw�㺟��;&��$[a(�Gr�"&V��r�r�^��Y���ϴ#�ut�b�qK����SP7�rb�7]]�:�,9�f%O���`�����̼����4���%�uu�`\�b�O���p"�LW�����s|��w0��R.�RT�J�:X���l�qqwK���
��J�u��3{6q��z��r�m؁�7���e`sy���U]g�u�^�b����R�"��DM���"�ѥ���>�)F�e
̋�ugAɁ�َ9�jK������ݲ���f���;�5m�I5���(��c:Y�X+�^S�*U׀؞�&�n�4��n0lZ�CT��1O�a���۴�5{�J؀��Y��S��葠����|�Ȫ�\�j�G��;x����/H��������8p���:�/�ϵNDi���LX	ȣ.�QL�xC$d,;D�����u+n���]ǡ���Q��]��̑��R�Z�c|�U��A��f��)�^5B2����Jm��q�q��1C��=jr㋡//�m��h,��U��2�J�>�'�
#ɮ���-}�Y�[t,��C������l3��O���0�HE[5�s��:t�j|�M:��>ȴ*t��x�6+>DYO<��	Q�!�Qg�[��L�=,���J4�=vy��Q-��-�۷KvoN�ܥ���+>m_QH޺�� �X��,�\@X�]]����@S�<�[(F��1����3��XȻyբ��j��]�ŦDAKt�/t�Vjo�M^R�F#�v�K<~pP���I�t$fe��5�'j軣uo&�у.���o@�μ���F�4��:gm5����~��=PP�e�����k֢��}�����5��<�u�x�rބ��s�5�m�M����]��:�\��[��B�b�g�4<��-��0��^�]j�g8��
�['vq�L"��Y����P��ɩ���N������(|�I��[g������U�s��yDn+�����S�p�E��_.�]��U���z+/���3y���^ɬ�A���L64
�O%��
Qz!���N#��	Q��6�(.��]+�|�zt��M}K�2��z ���6U�}V�2tQ�X��ˢ�YV���||dC�Nӽ���9����-�y��i�oe���j�CMF����n�s �AF���}sX�{�aB�6�X=d����pfJSj-��ז�������V�^�yd�s�k�u���6�S���e��	��8D�	c/d���lq��F�f�q�=b��6f���2*!�z$�H�t��fGou�d[ >��D�Gyܑ��"��>8ݐ��`|J>㔻�V�{�WZ;����9��zuu�n�s�h��d�d�J�3��\�rՇYǧ(�u�@\�,l��'q
o#y[K��.�c����7��[X�@wi��t-*�b�jK��p�[�n�(�k�ΐ�ۢI|b[���E���Uυ1[��d�6�J�`�.�i��C��x#ߞ��<���������sr�Y�㠼`K&1S4U�����.�$�O�b��9'�c��˭JC˨xn]ݲN�v��v��y�1�]ac�ha�ݒ�^�\0(t�]��:i��[� ��Ax4�;�Cz�S����m��u�*�B�1���ݮ�1i�
��1�;�d�lV$���/y�A7,���]�����	`�7j�0:���6�3��#�r�&�4m�Χiûf霻�_Mtg���������Q���[�3�ݚ�pAw�D鉕KZ��FJw� ��2����n{es�`Yn�4�����<�j���`s�-}ǹHNg1�Oa�ֽɡ����A=u�KΝ�0��r�5}˒�p%�����.#]�u�I��<���Rލ�Qx�w3K�c �t�}k#%���4��s�@�{gt����J�ֈ KgQ"֝��S�=���{jPw99��v�w׽�w�0civf��%z\<=�,r�\�u��[�C�-=]6���!W������+6�zSYc��=�5u��m��X�,e��9�>@=�Ĕ�߼����{�����ւ��2�b�A�h�h"V���Kj�D�Dcl�ZFJ���+Z+��V�b���b�J��B�e���"*T*��1Kj�F
�[Jb�"0QE�h"¶��"��"(**"�VV��b�("��R*"���լ���(���
�QF�,���DD�mZZ ��b����cJ�TjՍ�Ė�D��U���(" �TUV�#��D�X��ʈ*(T�"�2�"*�ŭX��1EX�Ԫ
��Fڢ(��DUШ5��PDPb�

Ŭ���+R�X���`��b+��F�(ԋ(�*1AE*�#ET`�EDb�J�DX)Rڈ�+aV("�(��*(�JŶ� �[
F�e�2*�1ilJ%���[F(�H���Z�U���
��* �6�DQQ�k*TUcmm
*�b���*0_��0מ~۞s���C�Jk�Dx-V��ַ/n'Q��-�sx��幰���8���v
�W1�g�L�l�t����}_}U_rE�M�ۧ�luA?����t��TkK6��|q�����+�x�'V߼d��̠H[}7�5rׯ>��d�N��$�#�0CPv�&v�a�N���cMu���V���9R��Y�w!9�邏�>��;W�Ռ�>&�1��i�7r��1b�%����2�:Ӧ���c�t��(8�S����,;(?r�K�m[��&�����=��pzQ�ڮ9YU�3Z��Kll��b�ͪ�� l8�����
f�L�V^M�'&��W+9P�(���V�k6�y4U�O���ג�q���#U�]f`=;J��n����Ta`.U��F�c��!�ז���m�p�r?Z���t�F��Z�e6�%��5�[N�5�9\qF�L�1�ݣ炑F̎�
�8>Q:%
���n��~N'�����������Jǥn+Q�7B�[��2��!:�ؖg�W�
�3m��7�t�PP�`��M~�Z~�sG_΂Q����}b'.�yEq�Aq쾃*r�K��<g���F[9׭S�p'k���o��9�:F���(�U�n�!+K n�a�:K�(����EM�;�iZ^e���ܦ��N��K\-8�݃��z�� )���oz�;<Lk�y-.��sbU �Ӣ/�hj��]юkR��|i 6c���G�]�|<�ek/��V*AQs���%Ζt\���4�b�N��Aw�C�J#����V��p2w�=�b�!B󄞁A��9NE`=!���u��J*��K���6���s1���ڶ���2:���uJ2)�AױQؘ7;g�k��$J��d�o���uf��=s�~���4�uV��T(���	�0{)��M�Jb���ʇ���A�3R���v��Gh������Qҁ�x�s��5l�0F�rfF\,�Ö���2қun{Tb�v��5[�V6]���HBzAq>�b��!:9D���i{iW���o�hx�0���M�lU{ݺÊ��l�s~��G�:	]��V%LtXlȩ��3 뀺M���%��u���sӤ[�$a�7n�W2�n�(ۖ��N�����B^UȊ�kx������aߥ֗�:�x�T�asQE��s��kٲ�n�fĝ}1��������Y�;�����,�V�lM��u2+�z:�A���B�%��%��o�_mjH�4Qs����w�����:v����7hJ
�fѩ2���mu���׷�ww ��1�������>)�`n�Y�J"���d��9WT�lb�f���wK<4���9}éWA@&&[eM�
)���;��%�r�`e롭#%++��UU_{f�Z�%�=����W�*	@Q��n�L�>��7m�u�ʚ˝�%�U%+��::-�G����!L�W�"���|}�Z�
g�����A�U�
D�B�Q}$��h[�l`�p�*�4����������8Ҋ������z����S2�n �����3���;)�԰,�ZN�B�+���V��*�|�5G�Bq���KWfz%խ���#$���Q�5���z�W]mM"B���B�NF��D�Kqf�W��x{�e�v���T6v�o^�ݽ5	����P���->^	�b��u�Xk�����[*�e�x=�؉z�j�����p=%���V�S.�U�=~�U��&k�ົ�����U�����lT�� mN�:��[��t�4��S&#[�)T�/�da�@)�2��-z�G�y3$����IT1�r�7�Q���I.c}�4���b���`7�֓Q~�T@�֐l��J&ς��]��l=�A3䓆��䀁��]կC�@>��8&g� ��b��j^���}Ì���)���'�����W��G<c��t�����5ٞ�	5׆�_D�WU%s�f̂^��ۚ����y#�t�l��_W=�Q��Ǉ�N�X���
i=�Rւe�L�"e���)�𴊾6a� )�\<�h��_������J]V�EABc�n*bxW^��n0
�"Eک!�P3"Kq~ܚ*��%�Sxo�Rvz��u�����m7r���h�!]W���ϊ[�_��.o�鸣fJ�s�Zp���v7�{*-�c�7�
P!D�4P�4U�>|*נ��c����इ�j�ר��\ϼ�^�oTe���=W<(����5๹f��V(���.�����	�p�/�}:X��̡8��AB��.��f��"����Ww�^����'�*�*�x�n�$φj�Sc��^��J�&��r����X'����Uʭ`zeV�|l�)͌�(�&�D�lᾛ��ޗ��J��&
��ծ�ٕ^z���X�#�(.7���hj�4�2�'��][��߫K�4��'<1q��F�X�w.�{��}��������mϰR����J<��۬�Xɒ��>vWZ�{2�]��.9Ɇ����+�P@J�د_W����Z�;[sY�]�D��K�iz�"4���&-9eڊf*%Xv�V�[�ق27u`!�'��#Ӷ���Fޛ�6����tPn�b�e�y��jH�b{Y���|�<��l.�ϸ���~d��Z�.��V]���o$W��<c8��Ǣ�8��	5KsH���͂3�#f���quf���N�\�)�7s�t�V���ŗ���>�=��xz-���8����;Jy����خR�V5��ŀ�U��z�"Y=94ZɳS�����p���D������`�p�8�)W]K��Xn�K%�P4�j���q��I�F<��0?�XC�T!�|Q��>����{�ƪe�:�򶃃ӫo��ե�H٪�TuC24J�q]Dq��Л�*0`�iE�An&ͷ:i=�1��
c���&/e�pMsO:f�Qx<"O%�B��U�|U<uo��B����\��S�!X�@
7��%''#C�l:��A�gD���=�L0�>xz_|���e{e�FOa�۞���y�邏�>��Qؚj�Ɔ�^�X�cղ��F��}��fTo�H�{2��c)��4}9Pq�0�	K�#�IƤ\B흮�W;)�%n1��w��te?Q�L�K-�7�
��=�(������UY�oj�<`�`b���d%4n�d����ً8�}���]�}�
Y1uq%nD�E9@��\?�W�R�)� ��GF��� ��X�>�g�ڔ��:�D���ɬ����7��zv��7&�Z��	Re�Y�c�&�����N�s��'v���gLͼ��4u8����&R��qbk+M��Qݚڝ2���o'"fs��v��?xxxyb��8��צ��2F����/>�b����Rj=�k��m�B�:���ޗ�b&﷕��h��r��=�����3�r��0���1@<�6dvHV����4v��1��.��u��Tnr$C��|6)�X��*�DnE8���
+�Sg��^hp﮽��&Guy�䧐���ΐ'�r�{�}Z^z��u��%��>���qOW3�{]=:��[xR.(�;�b,��'�Y�h\iF�{�:��Ν�Zl+��9�;��k�{�{�D��%�R�%���Ng�ȿM�g�#@eN�.�P4��FDH�~.����t���vܷ��ѫ^�>�R���b�����F���Ϩ8�d
\F\"�ؙ�w<�ͳ���G�������*z(�⠔m����o*U���`h�fJ��j�1G��6C8LCZ:��zz� 's��5l�4&�k�fF\%Z�+yا݅�R�\e�t����b�e�
`������b��	���&3��@�����������V�c��ws�_H�t�D胷W���r�-u������X��ff�Į�גA5�ws��M��{1Y���K�_��ƛ͔xC9���^.����� ?��D�鋆*�.�g�t/6NKL�h�fz�G'I���К3�j�݂�����x�6�)(��o2��d]�a�b�F�f��h��	R;%ث	SZV��[�).�B��};�vc�Αk�8g�j�W2�nl�@�ۖ�8EY���Έ\����[��[�����l�뺂�jE9��"#^�c]B���R_�gol��@ϲ���6���M��xW(�g�􍈗��5�X{��L��tl5)�XJQ�d��չ����w�TV�d�T�AN;q��3��|tb����2 Ǟ}=�^��Xu��d�q�f�*~�͑]c����1F(��x��N�ɠ�*��(�A��({�Sװv{;+����������y���ہƔbJ�r�ndA%��e�_�-�ܗ�B�8T�8�fP"��ĩ�k�덡J����%��w�.^�ެE�e�1�p���{=r�e���#V�!W�5��R���0(��n,Ҁ�S���
��k:�I������d�Xͥ�Gq&��WJK�g#� ��l~�\6/ҤU��� !Xݍ��^���M2#0jGF��]��]�0��cn!*�7%�ӵ6y�vM�=!w��fzy@�m!�9ٕՇ@���.�(�z(l�jjw�S�5��j-	�u)gQ�Wi��Do��G�޳5U������d<��sj�����3e�L��
9#�u+��_}U�`��{�s�f32v~���B���|F����3FE+�f�4K42 Ҩ	�����w��tk�\S3���z�E{cv���'��8�ւ��
0J
�"�E�q��'�Nٵ��Y�'�T4��A���+h��+gE`��HH��n���Ⱦ%�!٪�V���T@�&Rvkm ,*��T�5c%�+��nl8&yH�1H�����Q��[#�H�b�po���#BC�l��ک!�P,�n8ɢ���������э�I0��왮���u����S�R�8*і\<*��qF�li7���Y����p���ehR%Ěy�����`��;s����K�F��Fؾ�&��Y��{�x��l�e��E�3��$�^r�3Au9xsƦO��>���#hl��b��A�{<-b87:��g�u�Cj��o���4T3P��}c���Y�����5�H�1R��t��KdB��b�6`I��ކ=`�~�{�U\�`zu��Br�.����&{җ��y�q3��=c�CF�E,>��8߬N�S�7�D�{ö�����ov�mD��bB �����8���5|��
96�|�V��\�:���
z�4/�v���p��"�����Z��%_!Ey#�BG1S�s��7�By.���W���|�i���=M��G�6TE(��*���:L*���jK����hj�=��JbD,�W�Ư̈̀�է*�~UOa`�<rvoܥx'ݪ}��AW^Nu�PT7�(���U�Bڅ+L^�czh�Υ�iÇ90�����(s�H�^��WV��/djR#3t;���8+�nފAq��:г�����#��L/N/��2AFG��RQW{��6�+�����D����Bq��O]��/�P�r�B�wy0�M���[��M�QB;a��E�9r��X%��20�EM�nƝ��q�ׄ��u��`&�\�8%��z��o��uv�E�A49���XC�ۡe}�x��.v��>ӢvU���3�wM"�u�G
~94@�sb�B�fE(R4���2`�H�t��t|�:7;��5v�t_�����1�Lχup.�pM�H>�L���x<	X�������!|9e.�������j�G��,]Rq`h�<(@zX2l$��XpM�$k3HjN�6&v��B�x_�e�o���}����pյL.��]鬵QJ�"�^̕���;�,R��c��z��hL����R�R&�Z����k�)װ�+Wp��_t��G;�e.��qͮ�8�-�.��3�}|-0G��]�[��o=�H߇���
޽`�&V񟱻s�};쐁�2)��eϛ�9ZՌ��L�wn/#tD��)�����ci�hlRC���5&m���`�/ܧK���dI�Ɉ]���x�T�z�wL�~�(+�"*"N���A�n��T�vǶ[�w��h���o�����ф<z�͝sӂ������_c�ӫƵ�f|�1�������p]Yxn�ݻ�]ۻت'U�;8}J���!di�ڮ�O�Qb�mxr�q�s�0vB���f'*��z�g$�An����p�y�IP�j�n�N�4�q���m�1^x)D�|����4Vظ�\��N��(q�6d1�3Z:���tu��R���@��t-Ň=Xe`Q^2���X���oi��Zo�L��=�-p��2&x� WO�ӥp����|�%G��@c�i9w�{�%vj��CLGnZ0o�0;��*�9�(�5q�!�.4�w:w��
計B�m��DZS3�Ѭ��ݱ}��dH49s�F�	=�q7NEo�HG&0�F���<5��wP-ٳsǭSL��z�T[��\n#���w^\�wg7��������WM{-�S��KS�P:{����ꇺ�pYWI�:�k�tq��N@���ЍZ�A��{�Q��m>�v7+���ˏݡ�� �u&��������K��o�w6�`�=ՙn����SsZ��̒����kV��4h��{ei�}h�[�;�)ٮ�p-%;T��%F���5��ۗ�b�IX�5n��ĸ�״8 ��_h�xB/a��ظ��(�U:�pp���Uoo������`Hh���q�g)�e7V^;(�K�2�������]�U'��)l�ti��5ݪPW�J�_co�"B��Qg����Ǳ�F���e�nU9�x�)���X�u�醟 ��ٵ�EPTl�Z�s֜����N�q�9��X�fZ!�H�o��8�ꨖU��HG][\7����*@����/q���W����U,憄�ֆ��`~Y�g�pL��/�ݔ�|��P�yj��q	�/7$�����bg��-�w�$7�]_T{K8(j���mY��ʣ��{J�ܲĄ�Ȏ��T@Z���̮�CZ�=gba���#�)�=��d�W��|q}�6ߴ=�"vNd�;a�F~ZR~]H�5�09\t��ߖb��-LU�n1���0��h�/jI	��fź~��c(X�dsGh���z��Z��%����w�9NS�������j�٫AgF�ƪ63�rs-��ύ�R�wRQ�N�����^�� ��N�s熩�kwR��/W�*^���L�Ocm����]>��m�I�m�g���t[�5���%��:��-�A;z������r�t�T3�̛t����
)�\���G�X��s��Yw� ����ګ�(BF/�A����hV�Y�A��-6 ����U�ש;�=�o�G�Q�=䈥5�^��#s8)�n�!Y"�8�	��.��I�5b�̆���1��d��L�`ʯ��g��ݎ��XxjN�zv�ё�
3��Y[="���uLQ�z���*]��V�]`�����F�f���l���no�p�{�kfòfҽ\�mɵ��v/`���5C��Sc�B@~䴿xO<��vd��n�]/��
�[>�)�4S�f�;z
*v��6�q'Ot�:��Z
�G���L߇T�eo�z�r���:O}�oi���*��'�%7��w�^j��ءW�z�x��������+NJ�S��"�vFQ��l*,r����}[Mtrs�m|�=�ep�tY�	;^ZA�N�R�f�յ�l����i�G��/H�)��Q�^�eU���G�kv�+ �����!%Zƽ��G|�n=�P.']�:5�c�Wl��{Dʎ��bn`C��v�cE�ׂ�0& =�4��n���d�z.`��o�&�N��v���ъ(�Em"�DQ%J��
���QAUb�E��UF#EUX�+,Dm(�h+mQ�VTcѴA�����RX ��(	P[Ң�Z�(�F �#")[+B�[eQc��,DKeZ�b ��UKBԱ��� ��� ���1cT��kDUTX�QAX�������cDj�b,Q�b������l��+A�UV5i,-�Edb ���������U#�[DQFҲ�ZYX�TPQE�UAkQ�����
"V����
+X��m�UR� ��T�F
#YiPADU���b""YQU����UEd�QTEQb��0QQ�F,TX�b���*
��������X)YX��DcmA`֪(֣X�+b�D�h�������
,EEEX�� Z��_Wo�n´3��[�v��Iz�-�5�WJܡ1xf��b�EsNeu���+�3�ݝ&#&Aw�� xwf%
o�hY�Ӫ����g��O�*�d6$=���lL����.uP7�E��i��ǉ��K6��^��8d��9�ڃqE�L)%�B�O������L2VG�<�1o�}<�4l�k�a;�V��=LP)Ń\��3^jـ`�,ֆ;<YS:���]
��])�~���Lz��|h{�]�'���#p��(�&9��Y��}ۚ���ē[wJ�{�Q�=m�aT�Xo�5{4��'��J�B����d9�|���K��,t?w1@�>�����
�t�Ņ'?�>���Py�H�7�29
�jIJ2�ٙ!���VۖPs������uZ��H��4��r��[�70�
U �"q�ْy��C��Y�(�/�Q.»��'40���6"h;x�z���[�bT�Ѱ�F�t�hh�RgS}���"�6���.(lJ��5F:u��3����!]�6غ�RjU��+]3�2A'}C%�>w�W
�QS�g?��q�������#:��p�t��:qzb.6{�����~��T����k�
�qd��ݧƞǂu��{>�[d�q���A�'���̞�j͋ݐz�׹���溈/��:y1��zb��|�|%^ٯ�#^�Yx
��n��g�l7.A�ӹ�Ăj��йX��x���'%*��2D�F��Q:'�U����ui��F�>7���zE@���WdѲL��!塴-B|��[h��R�"���>�8�$i[}�Sǹ�P'�=�b�\���H߫ߝ�s>3�qa.���ypr�����2��\�Ӊ戇C�Eh����.7�>Y�q�"�$�X��NC�f�ς���l~�\6.R��]���&�g_U��}�o
�ay�\i��U�=z�b�3FE ���L�,�Jgb*s4I�1�k[���b%B4��j��dP�݀�mEO7|p7u���dW��`�;[�С�ڻ�9q|��*�ҍT.ބK��>�;Jo����D�9�
�N����f7Ӣ���=9|��N��8���K�h:�);5��@XC�?*�i�v|�a ��� *�fKiy\Y��nVn��%R�������E�o��E�z)�M+3�ٱSv�HfT[�a��*���Fޔ��b�M��J��Y3M�k���f ��^�{�
[�_��.��V<��D�/~�+�uD�ƻ��>1��AlPb#E
��P�ֽ����b<���M22��F��N?{��+�Lލ뮊�'�j�@���Z�KGc��q��;����W�+~C_B]m3�.�|��Րi}�$̮�)�I��ݺ���5�GH������AJR���"�������e(�J�� �S�^�2���\ͱ�^�c�s��=��{��Seۯez�p#1JMK�W�h.�y�Ȭ�.� ��nt���c|���JJ;Sӛ]�Y�5B��G�p�(�hj*�;�2s��?��z,�ƽ��ݺ���:�3�^�`�FƢ����-��1���0:V*�V�=�&�\φ���z�����r��}�&�(`.��H�=����D��]Vtj�:�h�G��غ�h��A�zcmެm�K�|iz�����-�I�s��8��x+�J}��^U׀���5n�!M[�Hv��:UgYEGl>�p+ڦ���N Sr������2O�-=aX�P@T�p�}����8�cy����d?c�"�Α��V:gT�F��d�p$���T2AF�Q0�򲷃�w�T��)�r�ʀ������m�(���������\�UY��#3*Q�@�M��nD>@�n�Y�:	�U3���ϫ��#^���O�9q�ץ�����бP�DU?0�^�J��� o�+��QAs�܌�'D=�A6=@��V�EGؠ�qVq\�⳥�03\����z"*���,�0�r���Ӿ����K��{A�|�2TW�����#�mZ�9���j�|kk�CV7���w&=�=�ͼ��5kn��l����U�gذ��Ǖ@�H�F�FKqg�eP�%��9/��#��Y��;��jϷze:�$�7X*C26P�i���"	��Z�f�`ڍ�lU,D%2vs�]93����_WQ3>ޤ
�`;�hsH�Lړ:Y���s �bI��O�g�bv���C��ʦ�A���Ƿ��&�I�ذ��H�f���3rzVeEpZ7njS��|�QŸ�z��eq��"�1c���@��7�v&��X�u�U�����S%~'����m�Ӵ3)�7�ݎ��2Pp�7�w6�����+z�>����w}ǜ��iBa�O�j�d>�=kwM�&E7\o�*P;{-�5� '�WT��PK!�7�~�wx������ӈ�#ؼ�P��鋨�
ɢ�dO���x��,�n��|3�sz�W��\�L���i�ڮ�O�4*!ʍǫ�z�cx����$����$��~w�\;�[���h9��5L�1���x%{�Gd� ;�s���l޾�̾�C��[���7�볇y]Ã�H^��n�T��gt�ˑ80H0^CsSb��]���^��#�'�JK~I��g�^�;-X���;��4%,V�N��EH�b�W�zfW�=��kf.��8˴�j:�u�;��8w����ls��1��~&ĦlW���ј^���|�D��p�̮U�E���ꮤ�8J��Z��!�x,<�K�r�?��qO������}�����g���d*iͽ�ݓ����Ec���'���T��
�(?����C^�ҍ`�H����y��2|�|�أ����Ԃ�9��B+��+�g�ȹ�B���Lan�ؔ����0���ċ4�=�� �}3?4�|����_i��*9�L�=�
5��ZO��+��":�%�x.�2#�p�s679PP�,�|�`�M^ޗU�Қ�U�ηP�ݘ�5Boe`���3�V��=LW�q`�18L�;fAg����uS�|��v;��cԒ�#����βV/CO	!	���1H؄��J4=��wj�%�t
���$�{���lO[X_NP9��9���V�}��+�5Z��cw��wv���ݦ:,&dT�x�>����8�)@�g�v��s-��٢���$��������X�Y���u�b���e{v�k�)˛����^��rXp{t�Y��Z�Z#��;�pr��$��$k^>���r�3X�nv^l!��}H'M�-B�ٸ-�qn���̠��h��E�p����Y��L�0���<(�.TX����U�ri�eU�/� �*�@Ft<�ȓV�����@�#��>�x�w�ˈL�]>�����q�m��d�
����çH؉���+͊��΢�E1Ǯve�fX��=����Ԡ��\H��@ٿ���6%)@�)�u����-������8x�o�5�J�΄9�1<f����{s�T#F�=�E0�C�WWf�{B���}1v.��v˭���
h��q\|=AU����>kb���X��8��J�?��Y�8�Nۢ�7zW*nLSJ�]�؉�0����6®6�(�8�8%NB�q� i]�>���f�e�J�Z���i��g: ���ϒ��C�FXF��w���%�1S=~�ޤ�y�R�︧�ri���z���9�;><=
��|���x'���L��K���).�-E�R�Z:d,�\��J5E"WUa|�\{��dŨf��WH�fIg�FS��ݞܑ���YO�&�Fd������Exln�wR6�9�������d?�Q=��5b��Lj��N�"D��v���*���X��G����CS�Aj��_��wږ�@�&T�s�s�U�ꈄ��z9\e�k�33����-;:V�0�]��t�+�]�<�:u
�L��m�Ȟ�nDp����82�u�
�X�L�!���b�>��u�s�"ne#��4�{��0��.+)�4/3����K�C�i#�����Β��'�.���ե��7�i5�DP:� ���iax��.3�@>�ɹ�Tܡ�ݺD��@m��ᨃbcy�aѮ"�'"�I�*���i@{ˍ��Ȅ�������b���5�E��V�k�e���	���{��In�hݛ���Y9j����kz�[(N��1��ފ6d�g��(wV~R%ė�$A����8�Q�t�H�K:��x�KN#�n�了z�e{(\���H�%׹_����/x��I׭�i�&!�b�g����3��G�]��k<�˿�����p��U��J0�AGW{a2-N]u��'v�QR����y>��u��fob�H��3�J܉�V�� Wg��0%s�h�R�����`��;-�[�Vz��{��:N׍p��Ka��=peF�s�m��~�	4b�<�R�S���^>��X�>u杲�Ωl<�A㓳c����)�*��c��(j�D�n����7��%S�%t��vD�%���'�7�tQi'���Q�/G^�\�W+�In�@c��.g &���n��Vk�s>H�==�D�QF��D6�g���w������[޾s�O�S�I6�<fn�۪)�.bɴ?�U'+�u��������]�p+T���N Sr���.�a�A�OPZ%�tVM�}����
��sۛ8ѭ�V�B������_�h_g+'��;FWySӋ�-��s�����u���B�$X�D�R��o�N�o�n�F\wC6*�W)d+�w�z��nU������ɽč��B�%�vL�"Dd���+������G%�)���5˵0�z�v�켑`���(�%PM�zVo��*��ãk�5V3�����sp�琄s�x�L����n�TZ�fEJ���4�&�k�;x�Zu�=�����C#M8�}*�&w�����&��'�3v�֖lL���}�R��ru�g>�����W/*��"J 8�������	�F�GN�f�m��|��i���2�v:co��7���C$ g"�1�0Q|�}Gbh��1��=���(�)������ �2�#�k�o;���~�����V���������L]�c���큝���}y�u�E�ơ��Z(���ڒB'Vy�mq|oV�Sc�m����A�h�wRZ"���[\HJϽa>7��D�j+���7zSA6w�G�ѮT�Z˙dh3�qtƬS����Hr�"qc��}UTQ-��Z��ӊ1�XvPn���ڷY><)�L��9XW�Ȧ덁�(�l��T�x?[.(�k}M�@��V�{�ҙ�k	[Ծ��U׍k6���c�Y^�і��9k5=/j�xy:J��`�
�#aL���j�a`}H�E�����{ s�0}�y��n�1�ԑ�f�EDs�z�J�c����B݄�2�'���24�7H���FF-{���ې�b�g���"nF�M�G�q��]cgԱR����Þ�2�RSQ�<��ִ�sڽ�וnx��D��4&Q}]<h~�ZV\ێ����G�ܡ��0�!@�{���%e���^����'�؞ܪ�t�4z�J5p��g����#�xwc�#��7!{5�����Q
p��BO@�3��_���HGu�9nž�cP���+����X��O�]���ّgQ�yT�"�b�����F������q�������G���+�Y��d�o.�2#�p�ê�lsu��>�H���{�(T��lm��Vi�Ef��mJ�p�wD �v&����d��Tjx3q^��D �^u��}�.���k6�����;cpx�$x�����r5�U�M�Ȓ�i��Z�r�u+ua'�X�yZ��C6�+�Q����un�Ҍ �D���� �q8�ٹ՝�gfG�ʄн�}Z6B8LC{զ������X<�Y26���Dd��7����������CԍA�����jź�|uSgJr�zx@�����\����&k7<���0)���S �2M.�U��
6'���)9ؗ��9���i��V_�%�0�k���sw�8<[�������P�l���閅b/�傧Z�$��Ľ㞷��n����W'��������"����p����_�hh��fb|��Q�ڢ���vK��Ta~ʜVG�,�j����ç�4V���a��3���TnҼO��귰Fh����F�"��C��*��5��v4�wZg�>����.w�Tմ��\''˱hGG�x'���E3��U���r��6���e�-v�u��x��Ve:��Zky7�\d��W�H��X����~2�.�m��h\b���zQ�8�`.A�uY)��"�����������®6%@����N�z�U���VHbp�]C�̼�7V
Ƶ6X�)��"�+,���E�g!��wyt��yxZ>�pd�EI�sWu�f��{Odrq)��t�YͺZ�p�¹ن�zh�
��K����3_
�2D�wG�Tꎭ7�T�������0�w%�YЕ��Vr��iƅzfLTU���o��`�A[h��r��	�o��U.]����}�����xF(>�M�ry��m8d�\ljx�Ƀs�r���wj,d��Jg:��%^�q�m<NP�� �/��t�S�b-vv�h�}��0�ǶH޵�Dq�Td��q1T3�ޅXݛ�؇m4��r]Y���Ed��Jl�2"��Bv@~�����%o�s�!-��0��,�'��,k_Sh�C�{ܷ̳';�p9�N+K�3j��/6�n�ԁ	Ν,�p�qSM}��]J�F7��ڙH��K+vk��K�/�ی�ѷ��U�s��Ԅ��K鏦I|IK�.�XԘۺS���s5���c1�s7q�Y��v�gv>囋h�� ����c�R��WY
gz7I�k-��]�ԩ��R�\cc��ȥ��|�q�N�Y��:j��s����W���U�\���Xp˵z��䲘<
��2S��s��92�)7�܊���R�"x��0-��=ʷ��%~ͯѽd���z%���~6b͈�Fw���:�V��R���ǜE'���S�.u� S�*�߷ ���Qe�dZNd��9�5a�U��la��C]�	�r*[<(��ؼ2yY�����a�3/�ͽ�˂+N���ȨHF�-�]�-��3m��5���h�-��h����I��R�ҧ��̸���RJ?b"u9C�l�Ade�δ3�v��W�N�6�ei�朽��g2]�&��ծd�����r�򔕨��͡����9�;	m�l��{�����<�I�1��"����%��d8�ܦ'f�n�ц��-5jzF�c�g\�S�.J"uLe��v)��� ��Jq��-��]�-������C���BI+3%��TDe-P��;��n:�`{��9������/6Ƌ���w1I�v�{wq%k�C"�$5x�����x�c��x�`=|�sr�y2)!�=r��E�6kE��H����K���т�^�10wE�� wn���p�C�U�v1��u`�mL�p�r��]�g�!�����V���f��ڽ�{}V�!eJ�g�=�>c�V]��H�����d��)�+4�42�]ܐ�]&���n�e�!�cS�޻x<K�Z��غ�kN�V]��k�,��I��{%u"E��z`)�˰W3`k�Q�'ٰ�(i�A��r�\N�W*��'�VvE#$�̻�	�"g��j��*��r�W��o���Suh���O�n��Ij����N�Ϯ�>>���eDx�FP�2��+.uǡ�S�\=�`�>�e����~D��B�E�"�E�X1b1X�E�*(��#m�1�U1AET�k%V�0al�(�ZX��,AQb�((��,TF1V�,EF�A+QDb�cAX�Ȣ�$b�l(��b������DEV�T&e���E�6"(�A1UĮRԮR�Aq,V�F*�Tb�(��"F �*��E�U(���� ������(�����1(��[B�(�#���U"*�EU��8� ��QP��F1�b�%nZȈň#1H�V��Ƣ���H�"�-�E��`����Tb�f	E`�(���\��*�b+QjV*�Te�("F"�aV0�bȇ���|>�N��;hE�WU#7N=YAY�l�z�kz�-]r����@�;��[4芔ۙ���#�O5n��|N�lo�������
{t �B�������!8��1�b�s,���(D�������H��_n�Z��+wE..�F%�����^�S�QuPX��Ip��ςY06Թ��V�6��D��U���24�6)F��\i��X_)��k�ɋP�஑�%(�8��r����}9&y�ꄍ)�D�c n�ê5�G˪&|F��}�ۃj+���n�A�tb�Z��y^.�y]]#���L�g�k�0�X��d��lp��66	u�4��Xs�{'R�˧��`����&�ùL�\TL�@Y�p�n=Y��d����W[NFI8Dt5����$����L�H
�P��".��yS�0�S��Vg��b�I�'&���w2a�M��'��v���$�7&��V�k�e��y�51Z����B����ti�D��r.i��<��)���e]RqDA@����)@�u�f���`�4��i+7��(F�Mʝ��:u�W��Bf9@�K�W�iu;͆Ed	8'q�۹S��d�;�(T{9�,�۰nj�U/�k�ƪ2h=0�2���.l5�{T*��H��A�F1Q�u�ˈ-www���^P�
����*�8h�VŢ��5r\n�GHޓ+]Ԣ��p4���m�k��3Cg�Hg(�����5܏)a�t��v�G������Ȭ��T-��ʐ2����:PQ������EV���]��1�ӈ���0���EmWJ���0ϼ�1n7����]���4����ʃ� {jF�Osg[�t����1�sc�.�!���D|(E�� 6��۔���~���9'o77��k�+/p��ג��=�n�Ned4"���x'ݡO���X.�YLٻ3�-^F�8軒^*���OCq��P�4v���@n���q�J��gAh��qyV��.T���:X7%�	t(��=���K}�#M�70�nEuw�)׸r)��`���v�P�����Ul���&OW(ˎ�f�@݊���ck��uV16�����v�:a�:�BӯA��f��]�Z����	���g�ɓްɍf�2�A��lM����`r����y�U�Lץa���P9.�B2[�S��jN(�Ճwt˧��q>�]B��5@L��.h�^�`��r̊P�k�SN
�DY�T�J�>��uz��Ki;`U��b��Ҷ���z��S�2��e�P"^B�"n�]�o�-���\-�d��]E��l/���q�|����'RM���Z�i�vO���b�^�:�I�vŝ�M�*Kq����N�X��-�`��gF�5��X�ZQn�َ�ȧ��8 ��I��`�!��1 G9f�J�������Yk(��'�:��]�����*��uց�Mƃ�L4���~pM�:���R��&���V�Ez���RX�a�Ӵ3�7���Y!9�邏�߷��.]ǙM�o�'ۙ��٥���L���;0��{U�k2��~�n�gMNEX�u��I]�
j�����]���A�5tb�(P�r�O����'�t�`^�"��7�(��J�vCK/��]\N�'���v�Οz�=j���V�/�<A�Z�g]�;ذ:�}�^Sf�l�um��8���\P���J��2F����'ԌW����Rj=���g��i:U�3�BM
�����_IQ�PT>�[���9��4)��:۴cl[�o'v2�O�:9�]B���Wj�V�Ή�)�
Щ�s�0�;6}J�������3�V��RyV���cir3�g��**�,��D��4&Q�8��J��6�|�%�}2��P֫��S,� ��:����%Ҳ���!���f���MK���TzR��'qX^[����5� rb�*����Rn��޾�V��8�8�b)������cc�y���]��Ϋq�	%�;)YC�E�
42k��bw"*9��"^vo�~���X��~������h*:t�q(�4.4�W�.;lS�4��A%!��v�عe�Zl+��R�DH4���zD�C��(9�'"�ۡi!g,�ܷ�r���HZJ�����)�F�
����dX8⏔�2�Dt#�3o��gTLm�f��䱷�!ҟU��a$C��ͼ^��-�7��n��؊,�J������u��Q�p�v[�|�eߘ�y�yP��Ϩh��A�n�V���`��
q`��jR��bi�;��a	�e�ɡPt�`�t�����]�x!�6t����'��dl��`�N�����b���Y�,��w�4(2	6�����~�������=�Y��}Wv&x9���Q��6	S���a�c��fEL�m
ي���-g�a�7j��p3�.Y��r�Clʸ׳E���'ZE.���ʼ�5a�Ȇ���#��2�H���¸E{W�B{�mJ�{��a�]O+!{6Q-UYz��ç�XJ~���ԠѾt+j+��벂t
�@��+M�1j=f6c1�n�z��񙓕���up�n]�k�6�c�[cx;�/cKs�C�#'i�|��U� ����S8�Q��S��CK�����q�u8m�6Gi�9l�/���}F��W����c��|l�1KLYudȃg*#�č��pױIq@lJR���-T�U9����h�6�	g�Dx'�|�E3�����r��6���	��zN�L}kȓ��y�6���t¸p�=~N�ɧ�W��R�=~�����ipp��l�8�z/X�3�+�1=\��*ᄚ��ӽ!��r�M�\l	FP"��Y4�y��{�p���`
+�Jߩ���5<x�{�:�S�e���q�HT��_�R'bL<�W�UFa��Fw��B	cgE��P����^��Y��E�I������3�����%�i��Xn��t�9]��<;�*�e��\`��)X���r�q�����E�3^�+�۬wP��az����U�ZAč�f���(667`;#j*y��q�#W+{�6��A�Z�@��dTqf	�F���#� \
�FMz��7�:�߶	u
�Ψ�}���a�ڑd?G!CF��<��5܈&a�D��$���S������~�"Eî�^�uj<P�H�k��
kU�O�]fU�9r����1ԻRN7���������A1_�	ՙ����W:�mw8b������>�4����Ӣ�K��u��w�p<SFFԖ�٧-�}�� ��^I�Nt���n7y�[V�jI���PL�*T`j`���n�>%Ь�Շبb���OS��S�S}�lJ�7%��t
[�ܚ(_�Ir�&i����f`�4+�cf�ML�o�������n%���D(�~2P8C,wM���q%���>=E�5��Jy=v���)X�5y'"K���S'��̯e�@����4h�_*�:���17T� UdB�?w��g������9��g��x&��v�����p�h^d��4��|���{j�=��b+�Yz�T��0�\��KZ���R̮j���6a� 1x�����ك:��M�1�f�*Sǌc���R�Ic�;�#�ʅvE�고��y��\"�F�9�Ϊ6�qx��+,H�>u�J�ned4"���)F)�u)��糆�^��3yʓ��P/ӳ�н�M).��Ũ�h�T�7(ی�[0�D�Ld�L�cg{6Ο8��+d9H�tod#rc#�mR���K�(o؝dûE�9��*o{9�!�qFU�i�y2f��٠/{%iU)��u�^Ն��Cz`����v�m-��4�\����[.4�(�z��;�Բ۲(�Quz�9:LX2�Y/Z�o��Důp]�J.�A�'U���,<�*���]H�R%��V�b�E3���*ĺ(@Fd���τ�TrL�����{����ȧv�S���zs��3n�c�M�z���	�U3����}E�#^����]���|N	�����b㊯J��[t0%�P6�T�A�^�hI�Ǖ@�H��[<�Vt�=��!V����>�*�Q.�tq��n��9��Qa\�"�
F�������ǡ<���rv��J��Ȯ�Q��u�L�KA:�t��u�.&����/]��X�Iܾ9L�Uz�/p�v߼r�4�ަ�����ݨ��.�Be�G�4���^z{�B�W"�n!��;�7�c]��vW��VWU����2��w�_{��I�I/��+WKg~�^c
s�U���/���^j�O]7����������7�*��F�;q
��ã!�.ڗtF���
���*�p�I�F��c���e�Y�|κ��r�J�p�n1A,oH
����\�O �gD�^@؉�'۬ȳ��ꌨ�gBw�^
�S<0�Yb���5b4���d���q#� �N���~6{���-<Vyy��!]Ň�Ҥ���:�&��o����z~��x�W�}�w�B����]�4��8������\Zr^̘��{oN�T�h�{I���J-I{"}[ܟ�q���#jd<�8ڮ�XR1Qb�m�I�r1T6{���h��C�G����Vuq�L>�A:��7��Glw(e轈sI!1+��Bwq3uyH�v�*mM���|�57�睍�<>����ˌ�[��;#��8�a:���`�bEwH��|�z��+b�6�Y��ñS�ܙ�]�QOu@b��MԻ�3�^R���B�
��jYϤlUۘٮWxy�s{�]���M��+:�;�b�q!�
m{S�7�Q��DV�n�P� ����p��WZ�B���d,s#B�CaԪQ�^�"�ɡ�6jug�1�:l��Fc�u�"9�~.lsw"mLڼ���-1=����q��g��Z�k�h�U���<«�ӕvx�0��#A�k��Ѭ}쥝O�3Q�'�[Jk:D/\�lJwP]���V�ۿv5���K�vm �^��Ԓ��y@�9q�KpE���:}�dWP֧�ka{�h>T!����.џs�g�(f�oDZ��{ϭ�ms�`�٣�.�W��Iҙ��ö�B �3�6��n0�{������Õ���`�����d̆�����yv��Ҝ�EBc����/	c�⥷�>���Lm�ć��Cc!�ڋ�۬�����-$I��7����VҦ�+zK�6�j�Ve�vC�ѧ�n�Q�4����̺�.kU����:
���澬��rsR�LD�^�����r��Њ�F�����\l�he{y�-
��(ǚ�F*�R�"���)�!X���e9�ʎ���i�Wj{'nM�o7���>�
~vW��9v�=a>����huX+����4�펮��2�491q��u�J�K����˚��|/j����9�tE��R��<�5̰����.�m>�]թ��}j�p�<ui
Bg�Ȼ�4Q�u�ݹ����3Z��|@^���]�_�|�J����o��m��찲U�=WB��ګ�\�]���>)&2Q�=��qc�]���)kēkSOM�R�јry��3h�����zZ��6����+ތ��YfA�!I��W�-m�V�2\�����_k@]XA����K�]DޡȨP�|��#\0��ڨ��wep�r,j��F�}�NF��-�'�U_M�t���Q<-{Q�V'Qz��1��N�[9(8���n�]�\ήM�S�k��?f�
X�EzS!AV^�w"�
����F�Cs^M�>��o38��ԑq��Gpt
v9��*p$B�������qhte�x�D�a֮v�t��u���@�a�`�	EV���r��*�ת��1�3J�ΐ���mD�Ӛ-�۔8<�b%&�Y��Lf���l�*�{�v�>�����̛��r��J2�ִ.�4m<�V��כ$�6W�M6M\�IS=��bL� w�
^��:�>�����5��I7��꘷��/4W#{�Qc���gHw*��K������<�j�cc5��MQ�E
��/x�]�ҫ�j�z�ȏQ�����(ar�)~�T���3[�2�kv�5fGiu]�ʖ&�]�(��Q���l��P#��tЮ��߂6�v����˧������S��YM�Q�&Ć�c[p��JX�cKl����OJ�?T<`�wh�[�]q�6w2HnVp����e����T���_7g�����>�W��4�.^d�x��v����l��i(��5��F�Ԉ 9l��W=�g:�u*��N`�*�m51�E �o�Ó��2��Cs]�s#\���Ai��'j�T�4O]��kE�T�p��j�� z{ч�ѻ�~�gx�<���9(�iojn_9G��vJ�;tݼ��^�9� .�R�-zc����|N���H��Nf�@F1q������F�yf�Q*�Hv�)��m�1�˂�;��w]�x���`�QK=L�C$IoqC�z�x(7h�q�3ۮ�.jˇ���������{���T��F�멤����ʯ���՜ٽe�QCˎν�5ֳ�֗��S/%���@1�	:�c3�|3���J$j�Rq[ �>&�ГHY�ޗ��qym�u-ɲ��aϑt}���S�Ԑ�][�v�ٚE��1�PΑL83.,J�ݲ��q덧� �I�w;��������c�r�e䐢(Q�R�G���A���e��R�h��s��9��@�����Q0��piG�o�29��.�6�!!���$m�w�q��,K��(�f�[Wp:���r�-R���LL�
���W5�6�Q],6�m��[��j^�O'm><�1��,�zP\��jav؛��!J�М�)��#\�@��o�c��3��^\���lp�:P
�Z����}��n�6��]
FƱ3�A �[U`ͧ��ד8t~�}���mw�Q=ꞷsp�q����|c�eK����g\\H1��衱���+o�Pdt˖n�"2`ŷ���#��� ��^��٢ay���X;+������EmW3��"g�ڍ�	^�-�j�Q��պW�x����=s�w!��c��^��fWT^�8Yw�3�R�(dd�j/FVg���.g��� 9�ryf��������/C!��KwlnĩBy��x��A$�h��J�y�u�7;;WN�33�Ԁ��T����^��u�:h"�*29���{ݩ֢L�Z��%�=���E�S��7}�]�b�In_b���]�.�5;����m���&Zɓ
亹�q�K�HV��C�ka)��e��CPk�mJsS}�Җ����7v�9�g��q�Go��\�h��=���	�ӏfsu��^�l�3+�e��)�J|����^�n��m�Ds�j��8Sc:`�,�B����I����{�p7t��Eq�2�z�u���>�~��5/p-��*wpi��]k�n��ʁ�!O�����O�u0o%	��#v���tŋH:N�f�-� �$6"���#�'[��s9˃x� �Tc�l�Z?�#�$�I�ADb�|��2V�r���Q"��`*0��1DG)+A�,QEF*����IYH((�SX�[h�%�(�"��J2b+1
+"�-d�Ո����J��T�`�ADDAD����-���"*"�Ua�KlYY�
*�B�E�������Fe+hfQ�؊�*"�*-�V*�h6X2[QPQ[k-)����U�2���X(�cQE[b��EX����q��AQE-���e�EF2*��1�ZX�eEc�(8�Eƪ"�c[Z�1���)��PJ�DU+D`��Pk@TE����3UW�E��Xʍ3
�5
��V,U���Ue�J�V[P����*	����ɳ�d�p���c��{i�|Ol�5�D:���&j��'K��
`s��N���+/���ÆPqH[�f��.�>�|��L*��OÏ�]�ɩ���^��A�Ql
��̨���*��Od�ɧ'��=�:�|�]���m�r�ێ���$d;��Y�"��q��L�5���P�H��w�ժ�=�m[e�6�:<;�B�KQ�Ў�W�K���l�>�5�A�GT>?zIՇ_Su1�Ս]�=ǫ!^�te��n�~V��^�*eڪ���oDcɧ��̀�h���[1�+�,f�w�U��L�	���>��U.}��z�મ�����ȅ�'fy_@�[ju��0���X+�HR�6���r.-賁�NS����Ncd岱����.�fc�a��	�N�A8�b�v���Vi��Y�XǤd
�YN�*���7�o0��b��1-q�U��k�w�R�����'uDN��̛n$VҚ%��H��y���]=��?o5Oo�K;צ�ivs��u�؂�̙ЙEdA���u�j�V�|�a�53��Z�'���犲�ʾ�S]y�rn�Y�Ҷ���,��=^��w-��u��rV@�u����}��faH#=:��j�g����� /z�;+0��RK�a�b�V+=�{���Ϟ��met�J-�PqX���ٵ��7�=ۓgJ���4V_FF�;��wf�e\��/.���/Ơ�sy䷊:�}ֵt���&��!𽡨�O��:un�t�Qg���2\���S7��U ��S�p�������Y��X~���&>a�[��}�=�ԡ$V�X9�I��AϳXT��F<��Ь=�l�1 ����{���k���M�Ub;��H>�A:�M6��v)��f�ۅn0S̈�����S׼k�eCπT2�飫�[�A�vn�vo�,$y��VjӅ0;���Vq��u�g��=���b@�����|����5T)�������/k5'���}q@&�Z<w��8:�eB�7l�G#u��kQN�]=*�BL�};��[�9a�N�@X�Ey7�>��S1=�V��ǰ��#�Nw���u���^���I���=e�����{OjR�ă�r�d�1�k����rf��}��A� ui��3&�òf��u�w܊yjvn��� �'+6I(s)S�s�t�bdN;;vJY�陷t�c���޻g��]���d�k�B���d%��p������v��c��:
��^{8��Ϊ/]`�Y�_
ّ۰�P���,��]�����zzC��[B�H��'Ս֍����=)o�����	�˧�İmX��,D�n�Ɍ��Nd�m��Қ�:fF�&�c�1�d�I�q��!�Q���b����d̀��Q��s'�kȻY�b�����;Ed�\�[s�漓M�|�60Cݵ�q��2����]Y-$
��-�U�=������X�t���{4��h��l�f9��kPq�D���۫�5�.�М�V�C��B�GVy"�x&��2u{�~���P_uL\*9������*j%�w`�k���w?@TD�y�?W��"�37��VTt-����AI�4�S�S[#�\�$��ͬ0��q��ԃC ii3-��(�U쮑Do���m�'�Q�n��p��ݱ#G�9E��`,q�u�虢u_'V���H��Ly�:�#xeskk�ޔ��[��&��g-��;�dXtU���v��R=�29��,���.�.��9:��_�T;XR;����n�3�����ws�&�Z���;���ک�m/9X�넎��\Q�O`\�u�H��r�|8�P���k���5wV�z�>�a�x�Kڮw\�u�֭ �jE�F�-�:Ċ��]-VV7k�ua���r��>5��R��uZs�k	�y���!�ʅ2{U���nҜ{��!����C}��,C�[W����Eu(��skڪ4��qPz�{7[�Ld�6 ���₸�u�r�W;�yc����{q�.�E���κ��cpի�6e�GjУX�� ��	�N�k2�zFB�!�t�69�l�lGl�?b�8���	���	�捈�n�I��u�{D����>c�/��2{�<U>|�d�^۔+���"Rc)�u;����sS��څ`S����a���08�|�05sn�0��/7�ղ�X�D�ٕ�7���-:9 <Wa��.
��4�h���敽;���[��g��;�ݛ|�qZc[63L��Ɲ���ӛ�f�ݴ	���N��.��P�N�� Ӻ�X�Vd=w<�)v��K~'�nhd�9M��Z�\홝3�_�e^�LXO����l�ԕoҦ/kg�[�|��hz��h�f�?��	Qw9Q�??�T�7�f�VD��-��fc������7םD]���{�Oyg�rr{� ��G����B�r���E��=� vo@h��b�goP����rv�;x78=�t�%�1����.�j
Gf�4��)%sA�g]��e��1ժ�&ڿ9X�8썾H��;��y	�]Bv�X͍��bi� ��[�8�3�V�y��ţy�޿ z�3�u�Gs���öR�D�Cb�|k�u��zD7m�1�oM���'0�C3���з��eB��j�t�F��aV6*]b�����-������%�X�Y�T�M��z׵\h��Tf�ZorE��W��z��F�`�je=��{	�S�~��ZH� �	��b�~�<�Hy�O1l܅v��i�v�'�%6���{:�|�dq��ξ:0���P�r�T�.ғ��e��h�$p�����5Z�p����CXn�􊭚�u��S�R��=ݧu�a[���@,y"��@l<���;�����w�ߣw�O�l�?*��K�]v̈�ݗ6+��4��3�������rf"�]���.��sw�FEj���C�C7\"=��	���wc��Qu�+y������i8C/��N�d���̟[q[*s�-�(g"m��W����|lEW{��H�L�C]Dn��Neڼ�NrYو���;�T�
ʹ�/(?o!l��7�bZ���=�v�	ݛ��:s	�v��j[��Uk%�r�^].i�dMU{�U���(��M���h�����+�u��l�)㫔3��SO9k����M[ؐ9�Sx��\�s�'y��F1�'k*��흖�����R�6�k�l�MN��e%g6[�X^`���YNz�X��WH>ш'�^��v�3�D�CC�X'�y݌������3=7;+9����	��������S1JEN�q�j�)
p&N��Â���Wd�_w	�+x��
�˚��u4�n��D!9Xc��C�VSg���'6�-f�r�-'y���\�-u�� <t��|«��8[�Z&�w��7�ή�t-�mC�#�X
�b�`��#���M��V�ݩs��	����M[���eE��x
�~����
�ٹ[��N5ӧ`
/y?����uo��}qI��c�8���!���.�i�KG�a{<;��q��<y�륮w[U� r�Չ�W�*�@&���yrc�Z���`���T�f��^�ݥ:�Э��Y:���X�5��ݸB37 U��}�^�[�o��+1˜����Kf+��V�Ev��^*em=��^�P�:��u������`��0��� s�,����0f�lPR9�#�<��J�}=�>RLI1��{0��sR��čy�E1u捈�̙���K�c?$����V�}^�W�Nًct��n���vK���h�H�������s���C����4��#����i��Aer�;3��٘#5�q9<=u~�ֵ�tn�!Gxһ�N����E���J��.�p7o�s��+�l�j٭1�sK�ﱡu�+�u�}�YZd]�RY�Xo�֧jQyTc�9��ҟ}7a�dt�jȦʫaۨ0�n�u�5���Ͼ;�f���xr�@.�4�of��#�i=ʻՈ��t�V,��+I�\=R��J�:�8	���n!�^��8�����oH^��Q"u͉�Uq�M��9�C����z��y*�ſ)ۅz��������h���_{`@��x|q����9'kKyx�-�l^��J�P���.�.�я�g���ar�ִ:��ءP^�ӸVj�&c(��:ű��_b��6չX��d+
8�auxB<�T�Y�d�3����ܜNա^�/�>�z�I^��P�֭��v��拳�{a8�mr��i	���ގ]�sw+W
�n�t��bu5�܊�kib�ٽΝggyg��5��B� ��O]��+�c��rZ�.X6=����'��^�0�r�H��D�C�kڨF��8��Ճ��˩�)W�cɫ|�ə��7��z����Y�M�ɠ$�����=���*�ܤF�]�˻�gٶH������n��_�EG���#a�0=�r�:q���&��{s���-uZO��k��b�f�ޒ�\]@�^P��û�]���N�ƗwvPr\9zt&�\q��+�}˯��
X�EJdJ���n;�V(��+hJ/�"��o�l�29�r�v��0���n��a`�R�ވ���ޤ'l[��kةP!�Do0�ŴhFn������
*��\o�^�}���Z���G��n��(P���!&-+�Ȭ
�|�آUh��ct���΄F�8��W�幠2P��ء݋g(a�S�luZ����/1��J�>_�����'�Qޤ��\�S۳�H����=�^�����g��F�ޢ߯p�ڞ�4�)��ǙS�
�B�k����^*�?W>~qrj���s��h����Z톭Ԕ<�w��b��<,��\)�C�c
s]+V��pk�X{��]F]��Y��1^�i���6�gW�:i���Auj��i+����Hr�^(ɥ3~n(z�'��4�Y&f���+BPo&�J!���
�&��	q
۹(G�W�,��>�}�S�0Ǽ���2��-����M�P����<\�w|>:�*,_���yŰ�Y�yx��X30�E���n��˄{ۏ#�Y[B��U�%Bd����-M�[��f�R8:��B:�>�A7ciu{U0�����1�Ȇ�z~z|fgԳ�ηd-<�Gǂ���P�bk����V*��wPo��^���{
J��^j*����C�����D>P��ǵ�I�&�z=�S<����w���/t���)b�q/Hs�^�B�FSdM��n�EvE�l�Vu��ʜhB����`��$W�(��sꨗ]��9�"��jug�mȸ��֌+��홎mߋ����/쎬�Ζ�:s1��Ņ#����=YK����"7�HD�f�|R�9�����Ko���"W3P��c)p�ɶ�kiM���!=�Rˊ�{��abݠ^s#��Ph؉��e��DF�8��]��t�#
�z	܊�}��)╡��;�ղ��-Q�3�b\������B��*���������ӐZb�J�Q�̭�&h�7(���陬^�����*#��O���ٖi�71��C-LT����.�i=Vې�n¥�#��!�AeYX9�n��0wP��L�ZM�Ң�%= ��UK���� F���*C��\�U���WE�ob.�׺��Qnq��M�yl�΃y{�WY;�~Mh�7���[�|��s��U�Щ�j�Z\�(Df�Hh�-��I�B�ʆ�>�d�o�靝�wGm���E���A	�qZ+/��KK��ٻM�@�t�e�΍�[բ����F`��X����(Ǖ�B�6��̻�fٲ��T�ۘ�m�M�r�]-�4��P����� �`�O1^�[����+�Udv�Ȳ\�v��r��: �/
@tj�4���/���T�d�O(9�e��XGd�m��W�	�q��U�1��3k�;zyt{΁V�Ә�M(m*l�x�v5c��*��v�Ïv��<�Z��(%��	\��xR�u���ɑǨ�t��=l:��v��=��"�/Q�����V;u�s��u���%�;����Ĩ��r��!�%u�
Q�����s��6�<�085��eU��	��1q���Jl1]�4�*$V�3Q�ZLj�?>f�mv�oY��7YǱ���N��5)uM�}��%��/^����*uC��֊OX�yŔZ|B7�"����眷e.ʱ�v��:VL��s�<�T���"����G>���m>��f�s"��ݰ�0��>W8PX�Ϋ&N��j�5*�ٍ|#x��ط�k\ѽt��7yA�z�Ӗ�Kl�}�)��|-u��k��f@OM����Gcu��Q>f=o��� #t�hu�u�D��S�Q:!�J���N�וޭp���I�F4٩ ���������ы�L���m^��*g9�E;�:o����LI�2�n����e�oBoA��=1i*E�r4ts!]u��- ꃕ����׺*:LW8��Cݎ��wk���r�e\�;�mm�ٌ��DJ̥d�3i�����;b�iS �f4��{�-+�X�t��v<L��ڻ�k-b;���ZT��B��8�ԥ E��k�:a���mv���#�JR��0@>��ᛡt�)k���8ܱ��J�zy��Z�)څ��W������o\�]6��c�<Ϯv�uu}\�+���"7�̽\i7(�|�n���VZu���V
���Ӧ���VMbKY�{�R z���e��Y�؇^R��d*�Ҽ�O�N��0��ndȲ4��;J��v�B���[�Hv�������$}��=*NW�L���������{م0���rN���dqp����*�	�wVΗ��K�街�	X;�J���Π�i�V��JY%&��S�.PǕ���~�٨]6��nM�$Rk
\��|��b�DA�E#iEUF�Ekb�e�AEX,KAJ1eT�dEPE��2��ҕ��`�A�3(�ؠ���k%�Ȍ�6� ���b1UU*m���X
�mQE5B�D��Q*�(ŭ�����J���m����1����Ҁ�Am����jU��Z��b�ePE2�%b�R�kb�[lE��P����T+`�m�U�[DEr�PU0aUX�F5-�kе�A�1*��E�,�Z�EX��*#T1���YH��V��&9X-j"��eQ�����*��KJ�#�`8�Lh�[A���}���3U(Vr�L���z�g:�N=��S촲�G�;z;�Ӻ�4�.�B�r�E�;���]3�v]h�b4�b�;g����cFS��].i�dM>�{jc�82����0kn��]�.n]K�����r�W��9�%4��j�&{��0"��ݗ�W��t\�Ob�E��4:���5�ART�k��
��:�K��**�[���j3�b��
��#�P�٤V ��o$�,�Ն�%��E�7�������3�au#�Z��@GX�}H.u+	��z�����)���=�U��Pm[�����a:�J{z�s�}w�ʩ(zѦ������-�{���Z�=��57R�(�#�c�̱{1�ʇy:383ԬK��>� �9��ƃs�����m
�{(M���P�ūaCFT��=����W��P=�'�[����o���Fj��'kP���0����@&M����_��υeiPz�`�T3;�۽7T�ӗ���V��h�����3  ��TG�te>m?;�o�9�6��r�ペ�a{Vd�:M�o���ٹF&ۈ���L�]->�x�$1�j��E@�ҭkgM�0�yi�1�:؛/9�K�f��wt��1�����n�8��i���Ԡ�]�8�����EN��4+q焌�Qu�֍��MN1��뵖X��)z�������,D�n�:��fj<��-��f6��w�8���;
j�h�K��D)o0���F�H�e��};n"uj�17@�if-����-���r��B�>���h�K�d�Wk7�w�9}�E�q�n	̻w�\�C!	�lP��K��y��O�r���a�a���R5�wn�2E7��31#���UՋ��1�p�H�0�����p��T�ޠ�y�ͪΐ��V���)uxz���q�I�f�_�pS�O�b����u��g��ϓ3t�@��a����=�]ݜ�Y���O`�$1r=��5]��]v�Cۧ�݉B|�]b�Nc�����h�ƻ�S��jܬvvG.:�fe9ț�{�vx[3�U�:
�|��Z
�Z=�;�z����;݊�ޢDr�+@�.]]���7��*�hn �b�ԋ����N�%Za6�5�z�˨���7��Ws8��m�N�V�,����)|�r��� y���+F�+S0��~��'v�!�XO�ڶ}����Z���<ز:�"���Ytjdu�k�\��e!�khOhء��ݮ�XU�#��lj�(�ڞ���z�n'�è��ρ�T6���5.��.�������Ҿr���U�9��B��s���l�O2�:�J��T3�C5Y���v-�,	�>�O���Ac��s*�kێC�c����su����8�Ŏ����K�;fDsTS�C��48kֲ�����P�wz����F@�q>��X�`-���¢���,b�W=j���j^���q���=���qw4�M:S���a	���!и�H�q�ٜ̱[�hva�cx���#wzs&��sY(H�lm�idcS�K0α���g��s\�lM{�fG�y�ؐ�2�,�'[�/^��f���ayNf�7h{���ůq�����0]'����n�Ÿ���ϋ��M���´*0{z�}^RKygs,�F�3��3���Dk��לN\|�ݶj�u�.�fU�?y��#yS��ڱD�ؒ����8�{��LeG)Y�I�O��nr�ʿ�݊��yok"h5fCb����H��7*��{�	\���d�e[*��Om'��\��5]��T�(w�&��]�29ϩ�L�o�BH���Q�\��pS�֨*Iw���V�7�]X-��v�
�!J���̯t��q������|9��N�m���:ioMR��S��Q-���s2�.�#�)�#�H��H'^���z����]tcT�J�|Me�Ӆ?-w��W9��g��v�3�m	7�G4��׈(�7N����/i�o9��S�~���ШQ�պ<�[��[���\u�q�D�d��[��n��@by劤&��+����V��񾥳;�õ4o]�qJ�]C1:��ұZ�B���b�r4*P3:��0i��+�����`�)x���4���+=�"9�~.lF�T�(¹���Z�h��1�Cs�um����b
��©�۷�.��	t��̞spc�S=��#�kٚ��^T��n��	��L��"�bt�f�}���HW������J]��v���\�'0gVX�p�o����h�أod��6jו���m{�^[H;��>Aʬ�t#*c�tȓ�e,�5�˧�ĳj�p��2!t"'-g�2E��-�Oe�w����a�.��H~л�Xi��ѱɋhk������N�ȂGf����#CCl��r�)��Ü�ؠ����Ĺݶ��:�-gi}�s��i���N�u��I�厗K�yY������M���CEGB3E���95�K�М��[����,�I��1�!)u�5L�3=^6rV`�Z�K������� ��:��Ի��l�&�w;5/���X�]���4ς�zЛ��e�b��)Ո'�����o-�D���K���1b�(펰؊�
�M���
������KڰMeU��
^_Y�\�C:�{�mcg�(�-�>(���N�=���ȮqԬ_F�*��+鷽�5q����'ݲ��f6zIF�������ڛ7^)G��6�F_�Ŀ>�(�}���=-���g�������y��3�o���+c)�T�b2I�4\����:��!$��-����{�R߱�Y������U�[�F������=��W�wk��c렛�v������,f��0e���vW5�t�@f�]BEju맪���ya�����ک{l�����Z��U�ڦ���HV�j���Cc��Õ�ޣ.*�yͤ�[s�Zڵ٪�WR�L����Tn*�^͋j�c���g�b�G�@T��??kþ��9�������)*Z�]b��o�4��IGx�o+)GjZDv�	��<�	��B5��B"r�	���CsSY���+�[�f�Nk:��S���aP)��ѱ�fd45�m4o�,�x�v�:����V�2}v���\�CnP�pp;O�c1�X����.���%��y�n��̐.�P�o
-�ب.�+�-	�P��~$��8#��L�Rf���gY��v�3'��U�C1�gyN��Xln;���(]���p�n�WT4!�s*aٔ�3�\{\�ێ&��O��$�I�=!��޷:���K����KSb��b,77{��1p��7��1���v���v�9�Ƶڂ|5B��t�<�+s��p��d��Ҋ�y�sy5!y���+ޠ����хz����g��1����+vOvP��u�<��Y��*w�s���nU,Z����`M�O��N�x�͏Q�jW�'�T	�����}�.�#��WY�{\m0���1UHq��p�}X�j��\ܬv�+���jt#.�/oa㧫����Ò�]�UÚ�m>�5l�����Z�u�<�J�um����VV1�}�����!3�R�g�=�b�{ǤZ�f/{��=�u���Ӆ��Q^ʥYn'��:��y��*c�^��n�ИM_V�����6�5��"�Ɂ>�&C�^�Q�1��U��0u�[ZWvp�['��n�W������`�<�BW�eK^�t��f����ە�P��,KSX��������sv%K�#�2�ғX�M[������{��R�г�tm/�7�+4�n���#�³�:2���T��-��A{7҆����v2�J56��]�q�s7%�}�%HgVn�u��B�2.��!`�gή��q�0$�{��l��v�t�X$/����n����ܺ�W`�1U�HȮQ5����`-��=\��C���8�Mk�l6 ���+=Y}T6N������j0S�5�ޔ89�Zf~����#�o����lf��LsC]F6��R$o�픷��\�����u^X~�B�SM�ؚY���a��=�<q�����~�ƽ��<q���|�
�,tK���Țj���ƈ�QY�28Bȅ���8�8Qp�<t.P�oFoW
�\\�@�y�N���j��(]s��9Kսax��{C�SjW�?uyRT�kkc�z'i-UNZӪ{��S?6&wz�xj��@�^l��-��HȺfy��N��]�؅Xv�H��H)��_����N�{}��D���4%�=4����5nË+���3ȳ�hS�B��w>��3���H]WJ�R����F������\��j�n�4۔��U��VTt��� �7��R�6&��c�nc���/����i��T��`��u�������E�x���8��t4���t�a��s�{{ �`ĳ#nH�S��Y�=�3Ɂ۹��P�u���C�.��ڃ7כ��aC����]-w��n�[���؞B�257Hwc�����h&ק����ޣ��� ��c|7v�ֲ���Y@,y!҉��f[]�I�/r�M��n���J�1ˡ�3��ۭ[��gEl�f^�T����A�5d�S�"R�n<�Zf��U`���#n�,�r�5�@�<����1�w�W1b$4��Ɍ���>��a�r�� ��@��iJ�~BЯy�&.�F�O��2��^n���b�䘍sWO�ʓ�b��]5��)�]�O�˖�dkTe�2��+��y"4�����[Q�n��r*���-m���%����:�&��o�ٍ1�V�}�)�tS�J�mcL�Z;�P΢����xp>;����^��?�6CnܓӾ"�()ܔ��$�)��1g���z8��a��e[�h̾�!��SPΦ!�ETN��}���T|�w%���%JP�3\L���W��T�A�w.ZW4���}��t��6^�B1a���reG��MɜA�m�o��wPk�p��쫜�B�dSBE���8U��5�08l�|��^����7<��4�J�PC�9
8�uzs^ +��ݗ�t�&.S��:��Z�F<Xv�[a�F��MC��_v�f�>�;����;H^�2^�ΥC�mc���(�>l)U��Mʞ�3�s1��C�$V9?�����]կ�Տ��y.�Q����昊v�g�B��]����t$V�y�����p.���v��yS*�9c�ɽΗ���B��#U<2��|w:�tۺݥb�>YU\��YB�5���ݽ;��k"�:��F&]�j"tn*��l[[z�D�P���b�zv��M͎n�)p��!����E��6b/)j�1��b�9���}od���ņ�v��N�s����B�"r���&��ĳ<O[�!�_<�ɶqjR��Y��E��A[�e4���5Ś��H�G^fn�8l}X �k�&�U9�O%�6�;gd��øV��Ç}M2��|��t��nd����c���{Ӡ�8�#2{ҟ.�)�Kz�hy��TY}�g�������Ր�T]�Sa�E����U�qt�8��J��1ʺ���|�'8<�ȌZ�b�Ƿi��n��]գ31ф���81Ӳ/�
g ���t��]1|v�Hv�141qv�P꼧ێ�%�[�j�#c��+ŉP����}�uz���ywJTʅ���{����,T�eѭ�P7])�Z�<g{e�U?Ѿ�6�X^����q3�o�b#n���׉T�a�L�̟b�.����.���z�H�3���éVsP�eî$r����\Y��9�VzK�B�eu��Cv�X|k#;� nj],�b���ә�	x����q�ۇ���t
�3"��lܾHZ�|�\�XE��\����7J��ڽ)��Ypй�"o��h뀁�m��E�'#:�n]]H�5�u�K��,l��*���>�f�ND�%��-�ΚG)}4B9��2��W.�R�9�{*�+|�O�1�w���&bGS#W)8���my�������������������@�b\���M8��
����ϫl�}˓5+�zc������˦������ś����;\V�-f�Z����b�%l��/m��+7������2g)��o!�_t���N���K�Ѻ/r�]sf9Y���U��	��q��8ts��Q�\�Y<˖��ih˕��qԶyd��-�tz�������Gô)o�p���IE��]��,ޮB#��pٻ���B��ʒ9�r��Ԏ��k�4�������_�^U�=��՗Ԧ9�`�vM�C�=����(������Y�֗;zw7u�˫��W�6�7��@�5V�����v{��X�R�a�!OQ���jE�����V#��i��\�y�u����=��6Ė#�#����֏�a�]j���ƍj��r�:�ecZ;Z�A�R1]Aaֻ8�L�v�n�ŷ��m�����I�N(nM�i^��zF�F%38N�����dW�t
�S�+��mi}&�Y�bf�lә\� U�yjcb̺��,�
��2K�C�J�X.��h�����qe"8��QZ��Jp��5O��)���-����;Eͣۼ�V�c���O�^��Ķ�in���
>��H;�¥\���f�����*�Z�Ա�9Sv�}�۽��q���8�MK��=����n���*�\�|���$�z�-����p �s�쥠��z�O��(9:�G�Ķ���~{M�7�Vԥ��μ�Ywwb2�U��"<(��'�Ē"�kEF*�*F��k�S����EQU��Z�ъ��Dj�"ڴk�E�[c
(��TXփ�\Ej��Q�f-��8e�j6��[m���Z"�2�fR-�D+R�Rŭ�T��V�Ql��ڥ��Q��Z5���*ƶ�B�qE��1\�R��E\����m��"���ѭb*�Z6�����m�Qh�1E*U��b[PKekYR����8YQ��qJ33¨����U����J�R��L�\2�U��1*�j���ʦ"�����-U��ZEDL�r�-+����TfU��˙l�����8��R�,m
����Fe00XR�TV���b�L�����J4UUQ����qU�Z�Z�����?}�~?o�*_<�[��'0�f֣�{U���1�ͮt�Ίt#�ܾ�g�|�p2G��:���r4\��>{�>z���JBw��'Օ�X�h/��¢������
�p)�3I�k��U8����>�٥*nѷ(P{�Ĥ�zi[�Kq����Ī<�����gthy��R�'�;�
Y�wޥN.ɾM�ZrE{��=��ٗ��&���|ϵ���۱��o+�(eh!��]���p�x�D�,c1�j��Y���&����3Q��5�v��f��E<s��U��٬ܤ����R�<�n�9�
��fn��G �[����E���u�<<s���\�=�ds#]��=��]8k��Z��=�ܕN(��l[�4���5�5S��jÕ�����=x��W�T)�'�Qcك:��t��P���+�5~�}CV�gLڈ�L�q����d'W6�b:�C��x�ZT�3�PS�+ЬO����οU6�ٮH��L�&t2�]VG��!�y�����&��.�;��3��o�����r�0sO�׷�h]Y�w�:vzĢ���i07��_T���޻eU%OOo[2�w��pjVF�r5wa���u]Ja� ������S�I�l�յ��9���S#�]6Lޕ'�v�����ި�j�X-�?,a۠/�3W�J��o3�O��|�|���6�N-��sq�&���	��Z��S�j�|��1o�9G/�E��_h?��ۻU��y����r7ҽ̪+��f�KxVf������՞����Y�+�*�.��3��W7�n�w��oMs9'9����uQaW6�Ue��}YJ�ʬ�p���r(D+N�����[���uV��^
���:���qw4�O�Қ�n���jͳgg/0w35�A�ݠ^s=�2�Ѹ�d�������ǂs'�w"�s��խk	�9╣��}�|�\�oF��j��^����x'u9g�,�-R.���!Jz�W���]��>�;)��ާ����"����t�'/�a�s5�h\��1<�����˓]�Ty�:#no�s��b�I{�bA�R��W�۝����NL�Tyw���CT7��=��j��b��u�.��>"wNޗS���ܶ�w+������[%m�h���I�5tw#�ږRl C�+s�퍊��W'�����ӣunJ�&>r�ʶ�Oن����*��d�hmg#5��Un��p,��T�_*fztu�h��V����O~�Ql
�d\eoW�2���ʬ�LZ�L��է1�+��܍i󰺂�ʔ�
���4�|)�<�}u��51�J�������W���m[��ʮ�3���T�W�Xۼ�3
�h2vn�F��X��۪Z�o���P�n�ߔ���Pn^�u�v��v^�+=X���9��7���.��*���:&�����ʎfT�^�s]+٦��R^���~y��׼��b��H�Ԓ|�+���=�px-{p�����%P�.�fM����U{��}v��O�&�{��p2R�ǒ2<+L6�`r��f��p�n���maB)YH�����0��1b'�30�������{�X����7��v�s�%9i�㵚��ˤt>��s��}��8�')��ۊǰܺ@"ѯa����%nf�50$�Ie�Z�P�\�znbia���Z�^��$ƃ��	:�X]�
5�9��mJW�9s	���ЈD�U�`�{���M���N+�:6�C�OAჂ����&.�6#�1a���F[����}�g��0z������42VKc;����I^��C��6�WLc��佽�9�w^�Oll�e7^厼�\���Ꮼ�^�����⥇}�e�#Q�y�6'&���hМ�M=(ۘ���Ѷ�Ko)���Ƞs}G�o����U����q�hH����Qk�s��vc��v��
c�p�b��W��'|h5^��4�=1Mi��Ԇh��kzJ��#���eχ$��k�v�[a���:F�_�V��m��u��w� ����vL9��~�-�.�X�Pmc��<t6�h�M�ٜMO�D�21�s�*:�w|޷��P��C_Ǩc�Mܹ��&�ZՑ�q�Z�t6�v�/3�#�p��t#�H�W�����﬐ug�E�5����r�"�^τ�B��]��և*�o�j�Iyg���G��M��-r%���p�97ޗ���-�yW�궱�bX�#�g���<�',PDw>g2��O��{v�#���ʷ1:zNsJ�d3GM0ov���a_x�j��|��/:d@�+��l�»u�g��y]>�<0�Q����J�;���y��,�%׵����Y�ԅ*3ɗ6���
�R�DMָ%�g��.�؟c�b�f9:nlW���J�_����l���;N5��ѹ�<��ڱ�y�|�*�ٰ��v��9�@�b��b9�|[�����
w��k\�Z�k)�9[��;�aQL]y�b&`L\	��qs�QȖ'8=Y�˞�n��ϖ��Ohr��۔+���
�*�Ղg6y^���5�4w�C�;��Q0�u�~�����!	�lTّ��%c���2���f%�:\�f�My�2��tK�۰#2E7��RýF�%��-1�2���ʽ:��
��Mz�<�=�R�����Ƕ�AG'�sW�Ϝ���a�L[�����f��*|��o�w���+ &f�ۃ�Y���S�|���T�����<�Ĉ5���XE����vU����ϥ�j��/�f����z["��1]j:��m�b]CQ��w�F�����M^��x�����,
�Z�.R���+�0�4X}���BZ�}4��ڦ��s�E�s���}N@�[��{UC���Od�L\����ߤ^e�)�
��n_'89JEm��}3b���W\[[�-�ڷ+n^����Iȉm��<�6��/�H.(�H)�"�7�D��,z>s�����a���S���-8SX�(y�Q�iX<<��Z'�lP�^��X�][=K�>mά3i�P�U��q�HXuT>^�"U���4v�`U̸q�R~��Bs�X�rƵ�ƅ�G5��skڅ�v�gd��9�ß}q)�
��aߴI6�g��
�_������l��I�Z��qʊS���b��U�װd������sn˛;�Q��]u츊���n_<''`��n<𑕮,VR��no�jb���b=���էn�+�?w<�PRu�K'2ۉ�Sp݋�Q|�P��עť�}�|od!F�K�dj�Vf�����=�9W=XTXp�[�Q!>�;�TL����N��lp�6��U�G)�59�r	�w�T�ປ���}LͰg9{���|n���Z9��Kl8h��hAЫ�|)pf��l8(J���9:�v���[^�K{�Xi��4lD�&Z�Dn㋼k
r��5�OwM�\��)ʖ6��b�	�SB�qKa�7�bk�Y��z63�wm�V��z�چ�8ۈS�J틞{ce	�A�,t�^S�ȝj��>�5�q�T(�Sm���o&9�:Q�b-u�dN��3��*�سWVD�/Ԛ�Z���7�������`��͸��NJ���hub5��T��qVIY�]77�<7J�lt�k�B��g���r���z�)�}�:/ݷ��0&��؉}o�*c�T��X��:�h˰�eCθW���C+�-���!�R�:��״�T�cG�ͫv���!2�z�=��&����EM\��=mLga@v��c�T���ujg�}qA�P�(��2�%�Qm��t�M�\���дWk���w[���:���=|�_ç���{O�[�W`#gk�N�({mWG[�"���j��:��U�G �.���j.^;B����M34��� ���O]���_ٌyXwW	���t����Y�8��%�E�6��l�*��H$�{~�&�c=zSҮ��5jF�̹p�$��ub-犺z_�����4�h68�~��|k#hr%t�����x9�[v��5T��R�>l;^�P+Eb��ظ]��5;֤T�Ux#B��tw���o$R�D ���y�Z���m���Xgz��;)�;y��ݳ1�*)ء�X�2��:%\�Wog�\�a\f�w�-�1}*X�N��BGy�^)��6"G2f@hk����Fgem��������V�2n�U�S����;�[s��د4j!W��2�#��!���y按�N�����-��e	M��:]/{]�#���_�\�G{����C}*ڧ�̊+I�����V^uxJK˛e��YAn<�
n��7�f绯bm�hn�?m2��c��:��U�����(u�;���T�B�ÇwZ�^�X���A0جq�u���@���rㅼ�"hZK��R�.��u0�i��t-)-V�NK�����נ6���H}��s�	DI��i���Tw����X&-��ql�ʆ�m��Z0S��Ǿ�b>��1��	�y<��������\r�pȐ7��:	\�@<A�9E�/%��W� ͐��8�bǨ���{����.��{��t�n�~��:��{e}<-�^�Q�!��2-���I����^ȳ�vK���lEs�[��F�71�B[�87��C|)��{_v������֝�Y�f�DUQ��m���/s���y�M�D.P�O���t�L�i�%�w�xMzT}�I>vl���تU��c�VF.s�(E*�|2�����	r�<��T���YV�M��c���2:z�#����f+rQ��p�7�u�q�1-0�`�P:Y��~�Q^�n���wZ��F�`��H�BF�i��TYJs�B`%�2j�R68GS��%�W@�&9�'6�n���&��s�=0����̓%�%
�Q���q>.U��f� O�5Uk���)�o:����M˪�h�(Le��NxWQv-�Q����t<uVP�����V�=I#=�Ӑ^�����j��r�������9"���T�<U�#K�����i
�q�QJ�Qr	�7Ԧy�k���:�L��y��7��2r9��Ǵ�YN�G7;��>z]����Wsm����amjT��	��1�l3IZ�B���G]�f��:�}T��V���/JD7$��b��n˨xU��~�bP7<�B�\MjN:2��0�{ՅZ�*$��� ����;���I�]]�X�pRC��|싔{7�>��^��#*�`�d�U�w˩�l2+ N��׼ş�x&����˹n߲]�^�Ҿ=��}N3�/��ɀ.���F�Y��(r�|Fx>�؞�^�%X���f��ڳ[��������/e7���VS�`t�W+X��^��.��yi����x������2e�-j�}Uf�V=t����P"��hs�����@�5�S曦TTF��F��[��C�n�.T[�<rvo�J0�O�a��^
����&��)IP�fŨ��LU_O^�oIuZ�ޣ�*q�NQ����<�<bB���uP��(пQ�ݔW�X��H�{�|$����
!�&zj��9����&-9e�*����Xv�W.�ξ��6z_/��n��� #aE�,�\�t2��W)d-uW1�j�4-:��C1�]CSh�Vr���|'n�=���3��8a��`�'�$J}9�*o�G=��{w4n%�s#��h]��X����zJ�֭,Q]-Õ����ҤMIW�c-IR&��J�
�鵵�#7zn��"4)D7SZ�k�H6���@V���<��k��C-P��/3{�k�U�Z1�j�kt���Zfز�����|�]�/ٛ`Ȋg�����b���x!�S��{ЮP�ۗt�L�(9j�^�s6��B��e��)?{"���9t��X'f���9M�$��D|:֙���Z��!���ҌժʐpJU�!��kF��+~�����]S���a�9�,(s�^��"�y!�����;4(nkuǦm�Nfv�O;{��ԫ���*�܁�J���v�������/���.�u)����a,z�؆�lJ�\��\�U=�]�{�d��8մE+���m#fH�ƫ�����K�w�}(�A�.��A<�_47x7r�g%^-��r���
:s+�K��xkf.c�XN��榲�r�i�{������.�/K�����ү�Y���mw)�	QjO2q�]C�ӷY6_f�s��;�&;ʵIO%_S�-AN��S��ud�����"���2��6��ٴW.��ѓP(��!#xH�w�e���<b�H�gV�\-��d�ytɻ�������=x��\fp齿�Af�Muc�৭[��@�av���M!bj<�3*5�����ف�ۼ}_ٸT�l�Vrz����{X^=c/�p�նM���=�xs�=�&��s�5���6Ch��H������ğ<�����N�����]���94veͤ��.�<N)>��Ҭ0���dKŚX)���7Y��c����s��ţ�N�{%�ǳ^��0{����X���������v_A���i�)Ν8ٮ�F����6#3��, �_uu��N�
�FV�A_mwn�i�r�C"�M��ni�t�ݴ�L��eCkT�+�j�a����\�9h�в3�=�A��ݶ�0��֊Te�K\'�`���8�v�O^���Gz���FH\Mmǅ�*F�c��3g0C�g0`��:KGs�8���K��������:��Z�J�S�ڲ��t�G������!8x�)���--d�@��r��sb��&^�,��X��ϔ�˺�:���r)�C����%P���+L��b�tj���}���m+�ܧ�X����h���Y��5����%�u�'-4���ȫB|$�)9�V ��:�0���J�2�;�6�=@���B���X5o�N�{Ϯ��r�I��v_p|_�H�ڎ��MǴO<Ӂ�>]=�=� �#�V�9i�����W~7i� �}�|D�2��z�;+��f���w ���tW	�r^����O���3:��򸟪q-V\�T��\�H�<�;|R��Z]٫�:V}P�  �	Q֢��Vʲآ�F(T�ܬjnd�YVڬi�0�fmh��j�`і�h�F�Ѱ�ƩUm���af*8iU+lQ�2�cC-lm�X�Tk�ԣ+iU�j�����ij�h���J��V�*#F��kU��(֊1�DEeK[*VĢQjA�UFµRҲ���*�K����Y+akR�Ykm*�J)l���#��*+mUQ�%���Z�m�QFѫZյ��QU#)J("�j��
�E(6�Qm)Yie��B�Z�U�im���R[j�ne����cT��F6նŪ��`�![KTh�EQ�li[iim�ڥjYJ�De,�l�kJҍQb(�U������5�J6��E�Yh��V���D�UF�D+Tke���V�s\�k[UXŲ��3jQ�J�iF*6���iZڢ���R�(�Rԭ����*Z6[�������ARB��ޏ�Cc<(}�x��
)_d����$�,ڒ�)d�5�ox�2���re�V�WY�޿���h�O�����[N�X	�_	��>�����x���q�З���`4�^E�8�5OD�oT'�'r&��H��2��|�n�
'!��}�U{(�P留W�[�ʲ@4�mr|��ե�H5V
��fF��ey��Z"�y�I�T���>��|Cw�p�M�8���2���kh�gShV��U��w\���>I�8�av��"��"se��F�X�{�q:%�R�r8(1 (��0d��N��$�#�0D��;����=�ӽ��h)ڼ�]������Uצ�Cr)��PQ}�o��MXj�E^&L��N�f��ͺ���C)%�4Y�~�gs%;�ݎΚ>��(8�_x%.���{h5"�_o<�6�-�j���=�{O�lS%,���_���P���@y���&2.
��}� ����.~��{[�٣=����mk40�:b�3²h�1�(���q^ޖ�¹�|{{�ҫsV�qFf{�=�WY�}����:f������=C�;!Y�8-Iq����r�ب��C*T�GÈ�
�ô��ڰ	�}����|-?-���5�"Pim+�DY���b[9�gR�҃���Fv_=�v�Ϯ#�r;\�b��@���G#7�E��25�:�gL��)��1�f[��ŜwN�^�r�ؼ�y㣃^�.B�+�Tz-����n�4�+�(�24�[v�<�<��
º��#��Ğ�9�i:��1̠砑���J8Ӆ��lc�:ۡntٕ�+�S�P͉fx�d�t�x!%T-�S���&t� VK4���.mFߚ��_C>����w��t�]J����8�K�K��B��y�0N�Uq;q,�4.4�^�+�p�\������j���2M�x�ro{H�X�1Ai�T���:6��H5WmX���5��U���Sm��Ռ2yε��Kn[��`�>��Q�M��*#�TeAȽ�M�,�@���+�&���B�iI`u<Y]ᮩ�?F�P�ê�o��mA�E} B�Q��oK�9�:��6np��߮����./d�>c�f��f�զ�����x�{��&h5l�504�S2Γ��*����V2%^���Պ��p+`����\o1(�'G"�QLs���T�b��C2��he4�X��F	wT��I�ľ��½�l1�ޘ*�˱V�!�)c+ewY�v����$d��J�<�:Yx�c�x�3��׻�ݪ�hJ�=�Dd�n\���X�k��w��W�Ƭ��W��N ���A�v����ܜ�����ɹG�������Sg1�:�T*�=@K5��m�t��Q���%�x�A�� �Z�M��W��Y��WS��D|.��fS�_��S��AaI��Q/x��c�<��"Wy�i�j�mP�1���~�)"p�����AV�E_ǲD0��3�ɟb����{1-cM��S|��'k��&���>SC���O,ޥ{PiW�N�R��\�X7�"5��Jڸ</d����T�5F:u��3����>WF�M�.��I�A�^��'|���G����z����Шq(}�BՀ����`S<Du��H["-��b7�-3���g}�GQ>�'���5�i��kC���X�~�#��9�O�K=���Ώ�\�v����F�@�L��aE�����������x��D������V��s���}0ű{�K��
�Z1zB�خX�H�����f���ȵ����]*��0�r��������Q㊸�K])�Y���R��la�p��=txU�#T�;ȡ��,��o�Otr�q�WX�«�k�k���Y�!y]#4��Y��4��5O*�YX9Ԉ6�y�Z�*5�o�2wE)l��;��%�5[`�Lzܝ�xX{�Tkx��\W��[�����Y���!ƻ�X�W��#Y�,�6��|��1oV�,����]���y38($�}��ٓ��8�om"�G�|��{��}|LA��Q�o�zQn)�������g�h�Dԍ��n��S���F�3�Ti6�5�e��Ʀ)=g_/�m�}�D)�&�x��O�K���4��b�	̓���&�jUB���d��1�S1���(L.�$���$w�����\+�&[��f}ʀJ��eh��٭.���+O�QH�*y��=ɥ�x�3b���t<YC�3-1սv�xg\�����-ڒa�;&hwPZ0��m"�S�I-ӂ���/�xUĽ裑�Y�B9j��莓�#��tX��­H�^h�t5^/���}G�My�Wc����1P�q��/WKՒ����u0D�K�W�k˩�lk�xiz��B��<G.�f����*��$����\S�f���F�T��8��((�F�]��ob{<��Dz:�j�T̹�>qc�o=��~�����Bӟ7��O���@v�*�UkӯV��^����郤��G��Ǉx�^�\��\+]s��ey�(Z5c�Э��wl�G��ۖ;�:隘��`n(β�I���MFf?+�wq;�h��M
m�t��kF�33ۙ����Ȋ��r��G�~;b]����<��iye�7{*'3p6��l�79��]ҭ��W}�\dQ�?�+����L�aZ�c���w"1��S�yVS�{A㓳`r�b��^�G*��lON@[�R���������&���t�1{�颯�Ԣ�p��L4A����r�
��ȯL#`l��ed4�&��k��[1�VO�)ƼT8ꌈ�i��s�&S*���a�%��&��1+���2^=�Kư$-h�+'=�uP��f\������b֪�BӯAR�9HL)iÆ̩�'�M�?L� �q�#�#>�=JW�8�����`%��T�:j��ڗ;���uL�3^�hI��*�7P�a�^�C���<Ϧ�38��=>W�Λ�p���t��@�rh���)��5����54૪DYO<�:"�Vf�n\�S�*�+n���e��3Ϩ���\��\ā9�7j�m��5���7�{~�l���;�3ͫ�[�����"Xʤ�ƈ� �oSMy'Ga�h�k35a�����:���KbsdT����z������y�^�$ d�pŁ�PQ�����Qؚj�ƀ�����|ku6ﯺiO
!�rHQ]�q����}�f�N	P۫ڒV��Y�,M?�4�%l���x=�%5�y�c�"$��s׷�)'c�r��LB�����p�Of��S����F�l>gsn�v�v�vyk���H��{���3���[fe�ه�or�N׳)�9)�݉>�(8�r�.җ{q�齉,g���(Fʱ�.�n�P�}wV�Q�L��X#�����,��V��{.�9�\+�7���:���8��͝sӂ��,���:��>~�?�kY�c��O�����g�����p�ǵ/98f�}-ꫧ�e���r�xڮ�XR1Qb�mr�q�󞡀�#�8�n�����"Br�B����-Y��w�T;���;Ӝ�8�B�c���F	EGd�a]Y�r�G	!�b��t8�2"4�h�j3��.�Kю�@�n��q�fW(��3�E	�)t�'���Z�R��XcGFg3{8��h��~j�Qc��uc�[�Q/�L�ML��r5��J؎�F�g����(r����J6z�J5p¸uø�c�{�2���4����myǙ��,���\��J4!'�8�&�)ȭ�#YS���4��f�:�UYp�u�,�gV�5�!�qG�a^u|�i�7L�*b�׎x��b<�ynu�bHb7D�5�p�.�9���Y [[�b�0�f��GyS��ui�{���ʯ��&;we}
ͫ^>��q�j�;%�z,{��eO��;�Q̔�}ג��8�[�d�3�lJ*�=�bɷ �,@��HⱣ�E^���\x���meצDqN.f������,��%�+�T���M�-/muT7��TmBX�Z}CF�f��w�5^����8�kØ�&h����kվ�y�aq�)���>�P�k�1��U�I�^ك�{���\N���tr,E���n������+'Mo��)ֆ
6'���*���~���X����|���G>��N,�*�q��n�I3z�q�S7�%�;��}3�l�:�"�xH��n�z�̷�f���;OD�F.����Wa�=���B�z��u���;%׺����n�!�H�,{�Íu
�}��n�U��QX�#�������(�����sC��j�%O,+ާcg���0��5�]�VC�������d
���а�Qq^���5B�v4盺�=���\��9��֝��:�]�d*܇Jͻ���Q���i�\!��Bի�}J�v.ݗYw���1z����cd�!��!��g�ѐ߶82�Z/�����3^o)����t_��#K�s��n"J�!]�������{GY3]��x2�I�4��z�W�,�z$�:*��������ԕ���
�"h��m�V��G�h̗��ٚ�n���,��)��n� ����ì��ۤX�Yz�/�w��;U���P���|@S*\Y�$̈�1]�OԳk��U��@�
g�r�	�u�� q}O~�0>�r�7�Vc�����U�%���/ಾ�8�~;0-@�$b􄙞t��0ϑ�z��,�5��f{���ۓK-�`c���.7��^r5VDu�E�I�����9fv< ��l�xdlڡ`p���.�mh���!i<�{��`E9�/��1��&fL�
��&h�G�*��pEE�)��]��z�<=��A�j��dV��06c=<�����m�2+�C0L����(�8�<�QJ��y�Q���ɠ/3~�Jo���H��~)�����ݼ���H���ހϪ�* ��6�vk�  C�?'i�rס��)�:'��Y�}�=w��h�=�U?|"�f�.�{��R	b��v-�z��]��^,ҁ�p�o���]D���wg�ܶ+t�c���Q3��i�51CY�5M
�3=Ѥf�Xu�4 ̤=|{f$�J��z��WY�����;�
�)�M<�B�U��L��z$�u���1��V,fvsx�b���{=�87ʲI��=@�]=Ϯ7���Wn[}I	W�c���JY+��
�df�Ƥ�h��Q+:���!L��l����~a�ǰ^�=�gTv��{��M�M\�=�Z�07]����ˑ�i���5����.ڕȳ.�{*�p#+ h�D���חS���8�&�U����{M���]�O&5x�\1�e�������ڪ�Uk�Ł��]�厴�M�OO
�UĽO9�d�d��ίY{0]#��do�H����|Vk�G�|^�r�{1C���|���}v�c�VFtwE��LS���P�Ȱ�΃�
�\O��.6V.�Z/$�]����VL�+�}���yW�{!?D9;7�Q�{�Dp!PU׀ߧ�	�n�R�nی؅�yA�E�gaEGt>�p(SGo8��#N9˭�y�����]AP�xd�UOz�0Y�ݓ5�l�i����db��Jt�*)Ƽ
��9��:ɋNEvU0��85ɑ�bz��ίf���Nr���dtig=��`���ء��+�VzKG���+���i�§�e,꼅����,^,�:	��gA#%�W��G���ǭM/�����K5�;�4����u�@�3edP7\�	�&k�hI�Ǟ�"}p���i�UV��>?|-Oy5��l?NTR�����x���E�&q����m{��s�G��9��(��<߳e��LT��� �
�ܨ/ƭU���kc�y-A[[:�tv��f��f���c9��-k��b�}�nm�Ӄ�d�V�{�%�*�$�t��3㢕f�*��EJ��*��v'�Y��L�nh���i�s��T�u=�+�M8(�
�*[QS� Ш+-^\�����m|w���/���ޔ
:�pkH�L݅F��~�����2���|��㱹aw��q���3辑�K�U7�$�P�oSM$��2M0k3HI�d�����T���;�o.2c?f;oק  s���(��s��}Gbjڱ�pNF��+֌�7����r��j�A���P��!���"O��A�r�-(u�3���.��ǜ��iBa�O����C�L���9S>�-Ξ�Bk�-�+��A�3�Y�3�5��o�;�]���VS��տc�<X�F2�C�����˨m̾~E�UE�d���%c��D�k'A�J�Q�a��t��ԌW����Rj=�s�2���YةY@��|�����Y6{/#�gIp�]v��h9��7�L�1��0�O+�Gd���'#���c^��X�
U�
�{\�M�^/�r�k2��F���m�ߜ�HIO���$��IO���$�BH@�2B����$��!$ I?�	!I��$�	'��IO�!$ I?�	!I�	!Id$�	'����$��$�	'�BH@�BB����$��	!I��B��	!I���e5�m�P>kU� ?�s2}p$��<z���$H���
�H%"�)D�)T�R��R�DJ)
O�[3l%M
U*OF�$U!H�QR��P).�����R���E$����Z�*EZe��*H����"m�������UBJ�(��$[-�H�E	7�J�D���YTR�%hT��$DRQ*R��f�*�(*�	QU@IH�E*J�QJ*�R��.̄��U�  Uw�m��gv�2�REuvYC�v��d�N����V�7
�P�m��:�k�r.�Yuݶ�q�p*�JenI�v�� c��U[mN���Eҍ$��#�  �׃�ݸ>ާ��v�v�r7[IZ�wa��0W]n��U�]ڪ�r���K��]UM.t�*�vʫ�]-۲�vkLJv�ʚa]�u�*��lI �Ҿ    3wږ7w �9.��MZ9�����ms�NW.���N��u��ٺ��\hi]K����(���zދ�QEQѢ���J  
-��(
 �(��!��+Z��OF���   ���:4QE����(
QE�����ky-�ݺ:����kf���[�p
��6ܨ٢V�b�����iZ[��U!]4UH(��)=�_    f�2��� �gUC�v��J(��uVk��A�юTu�4�P�8a�t	q��(��>��B�)T�����   �憟.�`BB���
1�WB�t�e٠u��q��C��]d(:����[���n�Ν���澱p��v���n҉R))@I	"D���  .齮�kU����N����Uֻ�v魻�5�h5�j�Vu�]n�t���Em�s��a�vۻ��lf������9Nٷ;v��g.��S�����T���X��R�+� g���M�]7i�ϱ�Uz�;g�ws�w��m���m�5�uɥi���t��WW'rP�e�\r\�;v����gjkN�Ď�WuKe)��R �JRJ��  ����V틶㩻�n�J�W����+L���r�u�;m�QN��mݫvWN�vf�]��c�:f�$V;�r��[uKtխ�n��m�J�R���Bx  c��S�N�%�ƻ:�[i�5v�wWAt3�E�k[�nJ���[�q��:U�8Us��j���r�%��ө��S.�qm�.mR�w�"l��%*  S�0���   ����z�%P6�  E?�M2  �~M�U( 24 $�I3Jj�2���z������4;�ʞ]y�^j.�e��y��l��~��|ׯ���H@�xo�_���$�HB!!�(B��p$�	'�!$ I��HH}����������5�?�z�=�w0��1�[�S"��v��5`�`��$U�v�;˖��+$PU��ҕ�>�SRzWh��2�:��+3+I�-˥�ɬ!�v�OuS�x�Q����c�L��m�Ah�MGUlr��@(�'� ����������e�6R��!�P&��+	m��fƣ.�+/J�guBu���,wue2�9i؉f�[%�r����c��[�nl���R��Rd%�1Ս�Kx����؍�r����U��Z��Ů�aҬ�#b�=��{{�(j��h"6�����#�:��"�N$2�մ��hƉ�P�o�T�t��*K�l�I;�Z���m�v*Q��7J�)�&]�!��Y�^����'5
�,[�͝�E]��r�� Ճ���m��-|��e�6�GUB�L�	��C�,�b*�3%����cv��I�$�f	���u�(�2m��:
dj����(���8��-w�]�GL����t(�X��
�i�.��Cm*�{z.�9nhoS���[/�JT�)nw(L���8DM$��e��S���m��V�M[S1�01�u@/0ƪiق���>�yE&�AB��N�w�R!l	�vd�����x��Q\�����*�eY{�����m�[1�e�cA;��y��hat\(����)���7"���+�Cen�9U����7.ӕ��,q���D���hm)�+4*��W+0���B�t-:�)�u��j�֤�����k26i��j�1��C�� *1�P�Ym�EF.���#���Ц�/R�1��G)Sx۔&)f����[A�$3*]��nZ*���7��P��aCU�#DЬ8p��k �.�7�k[��+L^�� ��6`ܩy��u���إ����S�Z���7v�-y��������_���`��ז�j��(���~{6e���#n�h2��&��E��ո��X��ࡴ&L*��۴iU6nb �vr�$��U'�R�f��h�͈�r�>w�<�{2�^�N���ԡǬ�i������J<�r�B����Uo*%�j�9M�J��D�v�"���#/�Z3�̠�̹�U�A��{D
���պk���Q����,��p�I�/EM���) YX�D�)"*�+a�����j�[wqç ��4�ۍЎ�ey���"�*��՜;;N��T���P���P�.�Ym���P���z�����񄔉�-��3h��I���}�+�EՈ�3m f'Ө����v&�Kqk�����Y@�Y���PV��4�=�ܣ������0&CZ���S`Ge�Q[��%m]�	Rm��`˛cq�K�2�،	��-��Q3��$Z�ckY�����Va�#�u��b駵*Q����[	щ�,sh;���M���<U��l������J�@Z�õ5�5	��MD�3��Ԟ֨����ٺ�Cwoܙ5*Pz�$��Â�	V��Y���f�,��Ѱ���vq�g.mf����v��JƊئ�q����G�܃7v�Mn���Af�G��;n8�!��
��Ф�I�S�a�.f(�!�M�-�Z7� (SZ���� �͚�.	�R8��m�V6+��ص�ej���1�,��Ŗ5�re�	&&�D[�R`��9���*�%*5�S���DUk6v�&m�*e�N)en�����cQ�aJق����&�0v����p�W �1na�4�{VH�V�R����3"U͕�7vIJHiC�)nn�6�H�e¢z���"Bh�Zu$� (]�:[Z�[�n��i�h+h�C�nj��e7R7V�+2ʅ<k@$8�	�!�u��� ͭ�OV)�V M�5�Ŷ��b�^�=Ph��,p^^XB�KVnS4%p�R,[,k/K�ji�f�T�و�Ӵ�0QR��i7�U��clq5���%L�slK�k	ܩ�֍b�AK(8�lf�Dd�[I��I<T�۸�쇣K5 +5�uw��I㫐
V��oP�%��)�����(�t6�JM;&ӔS�
�
#
��q^��Ȕ�Z�	����{�U��KQ������� ���T�3>	UvA�v4ID[w�L���6�K�fCln={F46S��pU�n&��,��[k.���
���[�L���b5Ӊ������;j��R%�V%�E;/2�*���䫧�H4"���X���WA��lfZ�w����!v�=5w�V!-R���U�6"lml:�ϭmc5n]
%ᗂ��{���?EPffl�ɔ��M��;QU�I�����ʵ���OX5�u]��Jy�0��EZ�[kJ+&���	7R6f��_ٵ���V��emU����e���C��U��і���л�mc-P��f�r��4�j���Iߤ�I�z�e�#��M���6�2X�[$p(d���雼��N�خ�Xr�c�4�i�?b�@J*�F+6��jQ��ǭY7�]4X-[e$`B�fBV9��(�Q�K�A}�X�*�ܦ��-��^�i���b����v��X���"ʃ\���w�{�Ln'�1H*U�f�J�l�X�jlK�h�K�.A�(�ks)d���j�}YE|jg.�
�A`Zv��ݝ�9�5 ���n��:�����i�R��N�!ջZBX�OQ����S7#�r�\'4�5�eu��U���/tD,��9u(�`��j"�Y�n�M�m�j�Y��l� h,� �R��j\�6̬��] ��b��J`��6���nR
��\WQAVe�KAfѵs�M�wG/���EU�����Pb ��ѫ�j����q�EK�d+4���{/B���n��f�	�����Gi\�V���e������*���*4j!�Ѱ8vÅ�r*u��%�Y�Ǒ-.�N�/jZ�����J��V����{ERP;���t	�F������d������2�$뱪��{n�۰�D�7[�d�d�vǬ8n6�<ݷ����|�a�A:������	Ϣ2�ݧ���.Q�X�c�ӫM�w�Wg5w�����1f^�,�*R�s1��֣v>�Oߕ�.]�-��ʏ\�m뺈�4nH�
�p�/�����l���WGem�e��"��+6��,�-���3#�v���Y;Z�oP:�t5C��]��15S"G /B)�$�!�x��c�#Le��eY�p����FJ��)P�eսnkЌ��]��!!Z��F�4��1ip+5t�6�ee�J��̄Ē`��#�X����ذ�u2�;�LU�nR�����%=�ʤ~����8�ܔ��GAT�f��Ԧt�nj5y��c�Q�5�.��W��e�	Y�6m�ZB@̐Rw[lQU�*���:I�T����5օP��bv�p�Ge�5�؎�W��"���0�*@�	�*�ʘ���2�v��-ܢ������b�[9)���GB�� ����i�){�ܧ@n�
����9M�a�V�J��V��ܶu����kXD'6[��f%Gh+	 ���nU�E9fαY5��r�)6�,]Dq�L`��=��,nb�( b�m��eK��G3&]��4^�r��5���S�n˃Av��J Z[V��t�b�8�jch$B�c���޼8I��RT/d�9�m�v��i��Ry>J ��pZ��e��[��vk0�[y��r���M����Ǌ�*�L`N�q��P�SR���^�f�ז�E:#2�P��\�'fD�wf�,i-�)��x��1 h�ݚ��q�5�a����'7	��ů1E����Fh-Oh-���X��
B2N3-5�˽�E"�D���*o�Ԡ�8΢-X�H�#�a�/`F,w5���(-�l�g3��%wv�B�9�r0�,U�:��E��q��-�����<02.T��VP۵C�TK�BT��[��z/���˝QhQ�\Xj�V�RlZ��X��i�U/튕n%r��T�T&�N�jD�����/�ZG ���c��c<k���k5�;!S/�ER1GS�ʹ����cJ�հ��n6mc�W��Ÿ��2�����i��6��b[P@�;��̥���im&�q��^��JSB
ٓv�<�\��1�ݺF3@�jI�|��\�-!Xh�:�˽�	�˕q�Sp�3.f�ۼ5dk �8���F�%�a\McY��z�r�H=��]kF�P�I*͵�m����ò�R�܍�nnB��Ç``J�Q�r�^��1̺��,,���J�l�xK*��Ȫ��1�Gcߕ
��,̧��m��y1�	�U��T����geIY!��C@���2�j��<����"Z�^�d�ِ�m"���n[ �%ZJ�eEӼ�X���6��;y���-�u.�MjQ��V�+�~WG~%��t��DIf�{z�W�)�ǋR1��hT�Շ6�Is"`kSwW#�G L
ͬ�V\��E�h:r��A��*&�ɽ�r�[�f�����x�
F�J�O/H��"������e��l̥���DY[u(�x�QVle-˖���SsL����P|��G����!����if�V�c�ډ�ݚ�w
�L޽ �+^�cB:Sz�.�� p����
Vm�V����S+��l�mn�����V��<$���+\�J��܌3a��V�9R��
�"6�A�v���KY��ef�6G)3o1d�"��>R�JN��1ɺ��G5v��ۊ�ZZ����+R{�,��t8v�as^���Ы*��E\���Bk.��VԼn�n��ܘBȪ���.�n�T���U���V��j�,^X5>��8��[��WI� B��1hך0�Ӹ��b�j�?m
J�-tf��t҃a���Sn�"�|-f*P�3p�dҦ���ֱ	z� j
�&?��b�zaƃڬ�� չw4 ���Hi٢��]��5K�(��+
��M6�Y�v����r�mA�{y��VodʷI�Ԭҥ��W�^�(U��Z~Ll⻎U2���ܗ@�&[�U��R.���XfRe,��I���a��(���Ԑ�P�Y�sDc�2 ��Z[�@⣴LN3�N�sC4��m �Ee7X"V�x�����Y��MW��.=�׋F$�Uu���nmZAVۂ^��F�7W��͌LE�!j�G2=����Kj[�w(�X�7(
���Z%3 ��p�G�i�.k��Z5
T�R�R�6���AV�jLT�.1eY:��{��w��U�F�BT2��YY���D�:蔮�(@�4%�v�j��jkCQl�0�WV��/2��ϳ�b����  oqH��I��maX���kMJQe5���[x�i�qֈ�-Y��=�S�3_�j�9��	�f˫;W�и�Lw�7mD��U�*�H"yy!����mKu���HX��t���-��v���֛W�`��QSf1cM�c�Q�ZfJ�PA2�F"CYB�<� 
�7C�2Z�Q�5�eĝ]kg�P%t�Ό�7e�%@�F�U6�xd���J��fZͮ2�Ƿ�h�E���Y$EN�U���fiJ:z���t���'��R�ʭ�V5*۽�E�H�XU��v���!J��-� vua��+'Q��0(��̨���u�Ō1��"��Q��qL�-%�Ij%�y��"d�n�Z'�5IPN��Uj��A@L ��(Ҙ��6^�2J�&��yT�S�bJԨ��V;�MZ�+ȷ2-�N��᡺�cv��BTZP.]V KQAZ��CMm��0r�0���U�P�sn�l{Y����g@�E�(�4�\�+L�.I)��;(�[����)0R�l:6\lꩺ]	���4�&+��K&غT����wD�)�ކ�̒�km�X��J�v�hlS$/v͛�f
�aY3(`��]��o2�&Ve��=�5]�8��~Y/hTr���m�g4&�ѐ���2#��^3{�:TB���^c[r����7B����v�+ �ԍ�Zb
mm�e@)�ҘV�Q��%H[�L;�;coq`4��5t=?+dHE�*�f9n�6˴�how3�zHa䡩XZm��Mm�$P�
9m��?;4�2ݔȠq'��.�3es������:[��h7&n�[�VٕX�ܼ�#��NksS�F���0k72���;J�^`zӎU�I)-�+	84ލ��f�*n�4%�m�R��3>�O���ۅb;LSӛ[5m\��*�w�m2��cN����6�̙�#�2���3Ujv�+JV޲��L��5�N5�ط�u���8R�1֌xd���/\�-V�veL�4�B��-��M
������:�h� �j\��E`b�gq
a�}Ҵ"-��ev�'"P���c��ۺ"'E5��
��R]�*2�5�j�+׮�����$�U�-91�TB7aw�{�U����m��Qf�E��4UA�
=#4"�}���L�/SȑI���[�IO���V)�x��2b�Jr�c8�J�˚eɶ�x�J��`��N��x�LiRS�Za�"e�.�[aMT�6��;��)�2��wn�Y5��<%��n�9��[�H�긅Q��;�B�"ua]�1��L�e�dTǤV�W+6�K����iUط��4#mu�U�U*��1����&٦Y�����d?���V��5*���x�7R����zؔ�V��I��J�q-�uzq�*��Yy��H\�Ʋ�F�I����ݺ}n�yV���}ù*N�B칔���r���b���2�T�@�0s��c3��K��aJ.<-`4��q$�.�}�O��CuIi�Xw/ )u��8�4��������1�9e��m�
�GA�Rb�
ՏD�)+x� ���'1���1��ԧ����]MڝDltuuZBb�pr�K��IX�K��t��_�׋���z���kҳ:��Y:�o�Ѹޒ�ˮ��b���z�+�rg������A�y1w�:hѶ����M.K*�}Ӧ^ɕ�iE�.5���b�[8JWWj������C��Ǟ�	8*�*�M�7p�\�݈Ƈ�mÕi
Ԥ�vc�y3kg͸h��c(�pV�ɹs~v_x�)Tٔa~��jYX\M�1�ٔ[��T|�\4�սb��Mt��J�����K���.	��a=�0����@�lu��do׽�4��"������3;���zYh�+�ʛ�}[u&u���W�+�b���E[Z�>���,=��!�T��A:KuW^'1ڔ��ؚv?F�ɳ}�F9!MT&�R�����j� �&J�����}��s����4��>��A��К�Gİ����k��J�����L�u��m���2�&�T�n���b�f;�`wy"�;��p(�7�v�D	����<i�尶�����Y�rd�-��ej��U֜���g|��ẜh1h��4Us�B-뭲�z�W�����}%`.&��+LЂA���u�|�l�U�֙�ȭ�tkH�6���ฏT��[�3t�+g>=\��úvD��:�9+{Y8̣s��&뵐%�$ ��B�p,��u�e!���;��F��� [�m�)��o&%��]r��:ʜ������+��u�:��	�%7/��:�=hqת�>����2�{�í�w�pX_Y�����ӆrL
�(�5�[`�q�ڰ*���j�Fu�#h�>�	�p�T��n̙��<�{A:'��u�I�%���s�����ݬ(�\��{�b:AW����0<�0��#l����=Y��՜�B��uֺ�.�:hiҚ�l�g!
�Z���	ڵ��t��wV���W�y���m��u���bǝT'Q,��Ꮱv8���p�رM�r��;n5�nR�/>��(֣��u��PN�g�gh|-���޳�07]c���%�oY�`)s�]m4���K�-�ͬ׼�u���S���W��m@��: �mq���*�-�C��Y3b�AY��s�4��r�9�p���Ƅ�>��Z�}±�Ŗ��������ʶ�5��"��m�ҸSQ�n�.Q�4e'��
 ��볗(��M�i�)ֶ���Ц��T�9]�fu^
���%���/�Κ�b�P���eI}y���}�����r7�b���x�C�e���ʟ"�Zb��a�8�mIk6�)ZAʽ�vα��So:��Y\�ᗂ��1�k����z�Ӭ�[B���yă�%����kMUv��5uBU�ue�`�6�ȅ�[M��Z]�0�ҵ�3��uW�/6�����G�Ed1��W5)Z�=3���ǳC�N�ڕ�j��\���n�y���e��J7�[t�F�ҍ�7���wN�uh �!.߆
�t0o^R�WyRR�9�-���ݹlg�uk��md|�
����7j%���^S�F��_s�0��|� 5V ��	�U�dI��.���\��+/{?�hA��u�8�(��-��\{5ASw�rĳG{b�!x�6�B�#x�^�\�Zؑ�6pU���ܣ�P��)��(k7�Mv�|��.r�ko����E�/������ۡ9@em�i��M��p1�>���J5�C8�m��e�H�ɨN���ܶ`�}L0��v�GCT��콬EN�����.�)|@8�/��۾D����m�YwB��:m�����]t��A-z�_'&#+���-����ʾj콨�S��W9W�t����-M>α78|��͍<���B�Y<�v�ܢ�]7BI�M��׸�F�|5B�z�iN�vt#�,'#.����a�2BnPr������ރXĭW��Cn� D���uw(zU�=�m3+#4��8qfƇ�2����r���8�T%Wg0wd��q���+������5n���u��U&���ђQ�x��{.�f��7e �"_��dM�ܬ\&֋�� ������]�U�:��"��&�$�Vs:��叇۪��;}AAc��.h�k�r)�"�.��S���)'EV��K��+��H�;`b��ao:�3������9ua�v������0=���y���s�n�%���]LI�)MT�"��jZ7sZ�@��d݉W�����V����dGz2�#�ӆa����n|�8�Hm�̑аb�D��{ �����mi�;�����&�g����Xy����L=M,u��p�V6A�.I�����U�ѧ��e�������]���#{\�<V �ed�����Z�}΁�Z�]��4 O1*u�jv�ֱq�NtRnq����W��;Yn'j1�t�x�ڕch�Щ[�5�=k�o(���:�N�t�1�a(�[�P7�3.�Z�H-
�̗���+��,U&D�S�C7��s�р������ۛ�%+�U����_R�W]�>�ղCm=�IV�Ĵgy㹠-[�.���ޥ�Y�汌�r�ڇ���Y˂����U�×%�b����5WA��e�W@ {k��j��,�C���*۬eI�
sS��K�Z!���>�A
��[�f��C:�=p��Zn8]("�Q�ëz�.8�4i���9�m%7/��Kx���αt���ػ/;n�H���@:��nĽ�{_:+bu�Ua��E��/�ȩ{��Fu�ZP�pW3�8�����sM��ȗfA�]�|1u�O+&�8�i����J�e%�*a��9mU뒊�;��M�j��c���0N���WVM��,�	vKq�5��-�ӎ�5�}Z�u�Y62X�wE%��ʷ�Q�on��3.�K��u�`��	����U��/7Q�I7�ft��4j�s�G�t��cS��<q�#�����[����.�*��ÿ]-!ĳ%���"��r���cv��=�h�[�Ωu/��e_V���$:yv�]���ts��7����/���8bѥ;�#���MЅ��۹|6�Wb�x;k;8ԥv���V��nֆ���y�V]V�C/���������=X9�U�]�*c����#��ӲcaI�"i^�ٜ(p��¼�|:SXY���<��;���gy3Ԉ�k]�ʽXo��R�#-�"�ջ��4�w�J��.���{70vC�w\x�z��Օi0�c0�Z��B���s�����; #���)�V%q]���L䩉qך�ӖF�	�Z�\@��T7E�vS����ժ�� ��,�&�_5�֛�*���l���_��Nq=}�3{'Eqj6�kbkyW/�ҭ�j��S����m�\��=�`	��BI�#{]���PJ��j��PN?u���B�3n�KzA��c"�C*c�`��Y���>�2��*�_XX�b��xl��5�u��e�;z	D�~̾�j��W%÷��5���v%�tՑ�[������ɸY.NCi��2�]
G�-w�f���-��Z�F3X����rQNŏWd���:��$�,�J#�����#._]\�Zmx�����3kTG�\�o�W:IeP����!ʁ(q������������M�s'm�w�z���XP��v��zy<6j�M�)�T�-��0uC����gN�%w$>�fЫ�im,ۇ�;�\�Qݎwr�0��8��b��T�F�-��!�Ǜ�-uB;���/S��f�h!}K3J��������wp�,��5�gj�m��t.hs-T�o�r�l�Ĭw��+�m��z�T gSr���sVf⩸��Qr�d���͗{�Ievgv^D�s��Ӵ�3if�^�r���4I�eG;:�#wStS�܎�dG���:�����ŧ&hP��c��cYs��2�Y��� ����_·UI]��O��	}�gnȌݵ-��U��"hU��'kYE e(#z�,��i]��{�+�V�.�4xX�*�3Ը}X]uwgW>���5k{T���Ip+���Ό�u��b�.�YS�5F܎�d�W	f�eP�P�A��3��v-�)'χvT�Ը�Or�ݰo���Ӷ�k��u-S��Z�Տ2`TEt�v�<�
��d�C&˨5>zej��gT!�L�ʭg-��~�`\{v�w��Z�����B���i����ĺ1�8�l��B<���5oorz/+��9���ӫ6C�q��V��TU�*��5��<��]]�4�g#�1K��54g_d�)���;K,�DN�����4,/����y:_=��L)�oI늝<B�ؐ[͂��5:wƬ�J���7�^�燬���]qZ7��3u�k&c	��k5#oWj{B�^39hi|�η���oC9�B�S��Tpe��`�m��9�EQ�x
<�菰X�k�,7Z')h�w�on52�d��o�PY�Ö],%�b��kOKJ������
򡣕ع;��$y�t$�j#��mI��8U�ܡ�b�*[��[�V�y�h�����k�%�|R���R�7F����V��Ǉ"O�7t���y��o-���V��F�g��ݓN30�L�W��0�=���V��/\�oxK`O*y�v��S	!U�V9͜�x�]��!m�{����4 GX�̨_�6�*̮�#rۛԝ�}̝��;��{f�|�Q��I�_5Y�һ�M[j��+u׉)O{�G`�[Y�n��8V�C����I�`Ҭׇ�dh��P�b����[0>����&�᷵ù
K\�������������xq+2����Y��Jn����,�m�������v�w��c����dĻpu[`7�����35V�%���X�RO�����2�0oNFPz&����W����u�����o�$�y���]��p^0�ْ�f;�{KN����WkE!3��-kޔ��g���l;�/l5#j�v���X���6�t�M{/qeZ]>�q�-��uur{�Q��Y��ݡ2M��f��ݝ|N.��@4%����SZݝ�^i�ʴ��5�GI-�Jogkj�xE�W������{S'(�r��j<ʘ�<�U�{D���,̡�8b�Gy��Z%�-�pܠ�3v�Z�[-mY���R�Yϛ1�m>��}�4Q�*PT(U�ss:�]�Lo �mG���'ʖ�s�q�s0R�Y�8��Csf��?p���ngv�Ri��]a1���uv.�qQ5ka�΃ua!����b\[�p�y�M��1V���mÎ��*U����.Tb�rZ1wl!V�ƶ�鋲��od�(,a�C^�e�M�Y&U��W���r�
�� ��v2��k�ems����*��[��}i�w\�"��/�Y4EX��&��n���ݮǝ�/i�J��G&ҩV�H�8a�Vpg:��i�mvAyJ���1u�>ϲL֘�ǫU;���}��R&����I"��d���d]p�DQ�N
��W!�{Q�S+�vU�%f�S�ӫ��Z�s��v����D�I�^�X� $͍M`f_d;Գ�� v���zZf���$h2Q�S�K"vZ�j��#f��o��˺"���9ձKy�����NBg�p��ۨ������`9�d�xk��;�����B�E�ŏF'|���9˴ �Y�&�=s��Ԑ�;vI�\�ʍ��n��V��󂰫�K۽C�5�r����u/_���Q��yē�N'4ͦޔ����x��ѭ��!�)_�t�;yM��8�YϢϥ�E�o$��Vt�C���V��W��b�^vԴ�r�1�R�d`咱��� ���l1����t�s����,v<TGn��D���J:���Hcǚ�VR�����4+o�d�BJ��̣x�"4]�=0:.%tB&ԙH��޴����<z��f�Z�{�hIfM�z^�E`iWl\�ފ�]�:'f6dcM]��&|p�y9�j��r^
�Sa)�܅�IU��{�d}�np�u�u��\r�nT���	]�E�!�S=��WS��*.`����=�û���c��F+7��Y%,����w3�fK�6���vs�lѕ����SGb�C��[�eq>�U���d,���S8xʉpoHI��Γh�w��T<�4��ޡei�軴�uc�9z��W)J�w�S7�.�Ҷ�ذX9�s��o��@ַ
G��܃�Va�+�e:y��kU�&�\�۟A�uiw��m�[���j�`��t��8`a���}&-��Pǆ��s�Sbin�����*6��ҹ���{������=M=ٽ�;������C�.�}NX���j���N����g6�gaٌ"��P�;Z��͝�I�C�U#��Bu�j�����z!�,Xs���TН%��k;qb�z��f�k����)�4u4�ެwWzeryYZӝ�V	̻oa�3Y�㋚�ۓ���b�rc8k51Y2
g�q�-��*��|�q� .������T��^�{���������LJ�Uv�}���1��:�һKW!�{M�EW4��[�D1��@�{��͍�d£�,�LA^��o�,�I�)�kpbt�i�+9ڹ\�Nr.q �-C0bޖ�^�e�W���&\K�#�`���u �%o���egH�.%�.J�YX���enq=gvr���AFB��*0���/y$�^K�$�I$�I.I%2�"V�%[�RM>�boN�S�	�z�vc;�g����BC��$ I;������������'~�͗5~��1}������ e50}Y����K����)�]ǁ����Zc�p������N]�1����KvLu����k}m�p������k$M�݉�%�T��QPԝW����5��eeK'r�s3��b��������p��א�g�+U-�p��m�1'I*�kF��V�x�����ph�	�3E���rru�%�7�ى�9[l�5i;J����6`�h䣱�Y�8"w]R�K��J�V��V���b�ίx S_F黦�*%cP���h�ڏ�YnI�G�S�=[���9Ca7ܒBvWr���) �bQ�ЊWS�R1fc��\�lX᧦���N�㌻=��n��\y`�|:��I��Z9����mS�����k�	��Ke�5�K��/�A�lI�:;����y"�_*��� �訥�C��s��ԙ`Հ�����Y=:s˹C��F4�3+���!%�G>�t�t4��,��4� ��ְ�<��sL��$�U-<���������%�n�I�����c.��N������>��b�.�B�#Uah�h���i����v���Y��Xa��<7@��������o�f����������p]��ji�.j����,���S�f項�j��ۙj�׭�JqP���ͤS854�ɿn�2�d��LΤ�I�ګ����̨v��w�HK��pըV�r�uZ�6C��F�����7���{�a�	����.e� ��-&��譔�W�ֶ���z�,�sM�*4��ʱyMEx��ᷯXoT��;V	��XJ�H�3#�YXazi<���H���,�Z�"F=h���������FI���㽘���y� .'OsD�U˩�Tx��H20���F|ʎ�C;WSW2����ugE��j'�f���F�ȢU�U���(4�l�}ԓ7.F��4�!ee8�}���f	,�@���w���e�@���i[�)U��7�V%SAO RY+Q#}�2ئ1��W5�lХ�n�;3RՋ�p������;]�Y��5����ţ{�b1�-��-�2��q�E��3�^�Vl��M�%և�cl�n�$]�&Q0����c]���`�ef�,V-qJZ,��\W�Zg;���]�+x�aL�Z��Da�Λ ��%�ymr܌٧N�ٴ���Uk�6�����f���^��H'l���;�"0��s/$ѿ��b����՛o ��
��EwP㊋�@x�6�-�3\Qsu�Q���4+�XE+\�`��'1y7��?,ZA��\u.��h�4)�En[ty[��r�v��dZ�����-ر�'q+��-� �`���ͼ/q#ڍ�$�V�uy���K��,�(��hkϠ�Vj�<��|�����UpN�B��ն7���c�K&+�s�k.�Z�e8ml@u��� �yf�U�YB���E�_��Ƴ�*1�q�.�9b���F@;���M,�Z��kv�Π�O�q�N��7l�'�:]=�����Ar��q��l�ˮ�˼X�
���@�/tL�Yܧ��WE!$��e:u�k����O��,�j��<�뽈^bI��Ae��u��P#�±�3	��gi��¤�c�)�6�bv4����W�c�+�G�`��u<�8W�n�|���\4[Z�M*�2�i3V.o�T'�m�o�F�25��d���� T�:ĨU��]u�t�*�Rؤxr�I�M$5l{�j�*�̭��_;��C��H
rxy]���rR*�ӕ)�R�)��	E(w v������&���V]�&�k'q���-�Ժ���᫷n�o���7�Qq{��1X�)��j�Gp�W�#P�V̠(&�uj���X�B��b���F#sZx�A���%I�˓�!�U����M�Rg�2o��H�������*S۴se��"�VZ�s�
��&���;�Ik�X+HY��ca�GusHu��c+��,H�ض$7$;zVw$V_:������0_&\�v�)a;T��]v\���l;�UbXz�a�m��ew.r��:yc�y.��ܴ�C
�9�j�9m�U�Zj��x��nV��j��<d�7��=]wbݻ2�yPs�XYO��h&c�j[��B��{,�۱3R���S�u�\��hm����:VI�ZD��ɦ�S�q.���֪]�lVP���ک4>M�F�����[lQ�٩���Kr�+wt�eh#�����<����U����aA0��V��cS�x4=&_'��(TZ��]�e�m�mb5d4��f�q�ζ���F�0��CQ�t�Fj�Ĳ�n�]�4kl5-��	˃*Րp�:����2�JٹI�:�",w��P5s�o���<�p�k�V*S��	IW��y��5lƨ����r�fT=Ocݩx����uݨ�����
��3.��W�O�8���6�xO���:TC�z�Ɋ�&�YH�쎴x�8�D3,S䲦�yx���=;�Vvv��[�9���Gd�Zuf�Cz�X���)7�!��{�<��oQ��M����(K5���(e)��8�5v���&>V�6t(�W2ӳ�98h!������������1H�b^w]�y���e
�,e���e�*KX*άqoe�.t��R�;Z�A��_fPJ��k���E�2�гH�;6��0��.e.�S�C�t7�r�֟.�Uۨ��l��^�}�;�wv%-�H/��{��T�SP�ec��d��_S2���]�ʖ�k'<Ҳ�˖I��(�ge;��OY�R�Xc�Q꺻�qM�f�և���nX���v,ʻ��,qpw����06+5�Ґ�8�v0��ڂ���v&�m���޾�kX��w��<D�ׁL��|�õa	CG����.#�eqV@A�gwG�M.�i�Y}��v��Q���Q:��m�J�H++A���cP�oW� �{�;h+ݰmuo^�ʹ�KD��a)U�}��S4���+E��U��Z��Km��J�2�)���y,�4�����/+��g=V�?E���vl����^d�
[y]����r�v��9(��s�gpqИY[Cg��c�o�0 n�4*L;ۤ�o3�v�l9]{�%���DN��զ�YQ��r� �A��ה�z.����h^ڝtPt����4��<�*��@Nl��/3zZ�:�.���4��5]�鎆Z�o[��4qaTl��]�[t�ܘ������[��9j=�yr��CPn(���4h��G0n��vƝ���%*}�Q8h�K��RU���n'm��+��T�kŊ�C�:��o~�w�L��h!�*��|�Rɕ���y��:�v.�Z���A��Ft���\�W֮YW}yU��r����a��/o�3�_ �κv�`�˙��)"(Z�ׄ���R�v9S�Ɗ�BO����=��dE�!݊��"��Oumsrر4ۉ��7��x�Պu�o_*b�.fM�[���ۏ1<|䲏s���֥���>㻋-�μ��=@!���xy�]8���zq+�V����
.�Rn�yu���;Ug��-��u3���ȫp��-��V �%�6u|�Wa����cM��!�A�Z��L5�*� �k�!Pg-z5�
�/�]��V#���w�x�U�����E����teJ��Q��*�wQ��=6�ѐrI��5u����<�\*R��;�|�\���Ó�S{@vR����ٳ�
�w����l��0�4�BbۃD�,�-���o&������v�e�g2�2�B�!] �-�ֳ#�*S���0z
}u�/8c�On�Om`�EC�Sf].�][ל)��e����Z�:���T���0:������^.}�2�/����p_^�g�N��[d$Xv3��x����k�lJD��&��@{�Z�A���C5�9AutJ�bѻx���5��:̀! ��WV�qcfao���v�8o�Z���d܉��:�8�)kNc�fY�y��;h�-dHh��N�׶�D�䊎�eh��w;E]��]���-��gY��aĄ���]'u�J�{+l`ȃJF��+��lb��Q��m0�z�}�؞�Ű��$�^�(��>�����"�(7����,�޽�r���Eg�nE�Uݝ4�D�SS�.����z)f��6�N���C��o�[J�Wc��B��ed[���ݯ��������]y����5i��]n*�P��tۧ�,M�N��Qm�3�$�P;i���'#�B�|s9����HBg&etw�Nr�M�4z�FU;�cu�P�S+��TG���\�	�@� �%P����1�!��i]�}w`7�o�L��Z}��u`	Vh��,^M;������d==3��=��hJ�Vi# Wu,��O��0ՉB�jwH�+ߤ��z�V���&�VV%��,��y��z�b�@����n<��_F �cp᭖\//1Y5�(�-�3��9�tm��V�$��M$��q�"�UB��̩�q��-��iKl[�n.Α�����"ɲ����o+�s���������ʭt���P6~g���|�[�}��u�k-sz�a��7Q��C�L�4MK��ڿ�G;�S�27n�S��a��T2�Q�b�}��=H`�;AP�|u.%WWX7{���V�<��u��Y���sqp��а[��n��e�[T6�E]7��x!ӗ3�sP���eu�X��s떳��u���Y�z�]*��B;{(�>�/�3�����7�nl���L���J� �L߁]a�#�)��(i�n��H��v2��#q�P'�[us��$s�5g^��5�OXTn�	a��(Y�n1)VWMj���;>�vq�Z®}�2-U��ي�e1�a��	i�K�0�ە�a\�.�uy��m�t�T��F�)ր�]gZ[t�0�66�>��k�7N�N�֝��-`	�w} ��ە+��n��hq�B;��ˬ�6�4�N3h`֮|(hW5����(�(#&Q)��9���oh]cƘ5��y����[J��xz���!6��Y�ݦ���A#j�zL���םa��|����_t�yƦ���p�qqŉb�2�N����(V��7nT����Oh^U�ɥr��Rp8F��]��]M�Z���]�i��t3�S�oA\&X�r¹G�u��k���@]z�N�V6���%����J�M<z)Y�ȴT\�0��J�Uk���>�|^�V����	�޽ʼ	��$q1oZU��OWmF�>�2}}ʐ������@��ff٘Ud�.�����g
���NXB%N��L�Y��G;���5�	Ĝs�����G�%��ka�-�x��mhW1Ic(�K��5f�S{����Aoer��+O��s���@Wf�������	�N��6�{]y�I�@��џ:溍�^���oP�`��Ig5(���3{m�n����Ƴ���y^=�O�}-e��#}��u�wwak�����@)�ձα���M����:�l�f��]2�#L��WM��6]u'Vgh���^	P���e�m�WJق�r�l���}�2q��4(Q�so�h��)�y�V�`���p&�dU���7x�]$�\s��8p��bYt;��ٹ�m�]N�}����F)�@<�K���Y�u���U���C��3��v�ƅj�]�n��s�ʲ��tQ̼�=����Y���hЕ*�Uwe<e��&}h@¥��\�3�Ⴔd?m��乄v'�8���F}ܣ�mV���p���Y�࠰s{]����zyu�cH4�
!s�4��F��[d)� ��P�G;�� ^���[��C�k;sn�SJ.� �J:�)7��^um�J�Ł#��n����G�C�&2�:��ze�}ǆ�+]Ӧ#�R��m�m�,93��]��B1D��nW��4��q T��}r�C׌J�;V9t�s��<k�w��b���.��)�
r��n;��)ԝFh�s�1Jt�k�]�Y�w]^v+�S���pA�V�c\ى�i\��������pR��x�S2]l�4^)xGT�l�/���ೖᒑͲ^4��͛�[�֋hI����ރ${f��"�T����1���?w�p���z]�b�rp�F�ᇑ��ݢX�]�差f�[����ԡMs7p�X��o뾝"�`�1��o�M[����������� fsh}d*݅P��h��Vބn�kkz�Q�Ԧy�� �kn��S��(�o�Tf�n`��N#�1��=Z���ͥ�7�nS"�r��Ԕ�>���z�՜����+u�D�;���ɻ+j�!1C�ܴثu���/X�_K�%@WrVn	�O(|�$r�i�z�������P)e�<9����U��,u�Bۃ3qW*A�aA<z��t��ql-ӫGe	$y��EpkM.r��&(�W$���a����wn����[��6�=&�f}z��q5��ӽ�*r���&�gr�$S����Y�
��t���̧W�HL��"��#,���7�b�n�.����:F�Y�6Q�i;N�w`�͚�"��l� ��E�m��*^jd&z|m%��8YWm��v��B�wr������]�[q�ީ\;5��5t�t�w]$:@�K:�u�-��(��sfu�zp���<���qTr��&���@��QoM��h��]غ酨��ɣ�;i�,�B���x�T ݺ)wj������T�A�� :�W#��l)>�I��k�kq�5���YԚ����ۂ�y��s��8?�~����.�� ���-�m�A^^:膅��ر��Q�oc{D��(�F�OD{ޏD{����U���=�YˇCmfU�;��n��Ԋ�>)����Z������r�8���Xn��.�[O%�ߓΣ�F�Ȗ\"���ߛ�R�e�Ҁ�DY����u�9)�����hwr词�]r���N'jeJ5�!��|%��q�X���K�ȁ�7g�uݰ��j,�U��J��X��(j�su��U,����s�`�`]��9m �ړ5��F���ΡB;x��)W�v�3������u��{G)�+V0���\+2Sm	���a\I�kH�� Ჳ`8�@x���=��O-�u>�3�܇�7����)�0��6�nӫR�;E1@�w�-	Bs���P���W\�:�;��GH���EN$�5��.�m�W� ��fb��9Q]q�ҕG�r+Z[�"ǵ���ҹ�����۴��\Wk:h�X�1��]ٺ�w�\�!�e� W=�}�w��]�2__�Ԭ�����lu�)�vvւ�C�UnYo�dɷS��R�+�Z�I�2��Z�Fp�:�&]ۭVU� 5q�i4�9��r�n��CFb���*-�"�b� ����sB^sw*���b��-�!�ӂ۫V�6;�=ۮS_TV�/�����g\� �&e��'���3��(���#]��"�E�P�s�#�N�Y+��1�gwu��!���9p�;��g1��V!W��o�8s�]k�B,gNR7;��Yٻ�V��w*I�� EB�[mj�iZ�ckcj[[h�.1G-D�q��(�ֲ��dSL12�m�)K*T-�E�M�5��,E˖��Ƶe�h(҉[6�m(�*��T(��5��V�QYV�X�T����2����b��d��ڍ�s�5E��2�X�����TYr�T2��l��V!iKlQL�ZJ�҈�TQEA�lX�
ʕ�K`�Z%l�*UJՈԣ��ƮQ�Z�U�Ke�l�FҸ�#JV��[JثR�Z�mJ	E��V%���Lcl�mJ)e-��ڔ��խU���(ڔ-r�bU�-���JR�kmJ6�j�"�U�-��ѥ����-D[V���V�neLm-F�kYE��KeDh�V�[q3
դq)����,X�2�[E�Z�h���iJ�F���hҪUX֕��5�(�b�X�m�\��T'�D�4 �G�W�c����a�n,�{hجv�@]^t��~*m��uY���9�^$kQ�Z��ѵ���xI�]M�v#��}�+�O���f��A5*�?}wt�}��g|�a\g���,
*�ڶ����;j�q�3��OwuȨ��Z��\��F��e)�Z/U�(���3�Ö�#�Un$v�C׉, �Q�λ�qw��`�ٷ]J^0c���`h�l�Jt�V��=3�pT]�;I~���Z
�Z2���}<Ctx����xmw�X�4���X�/�9A��tN�9K/�r�*
bs���FQ�~�4�������+8�N��qew��/WB�Df�L�~���4sf��>W�A���Z�I��=�j��m����Z���^>r�~���ǡ��q���w�f��R��&ajt&[7<����}:�批��t�ݘ�[j��~3�6O=�4Ľ������n���1�v�G��T<��'����SU���QK�q�*��>�Þ�.��3F���J+/�	�)K"V������~���{�7�Q�����M���eg�w[�����樾�
\`=�T�:��a���۹;mh[͂��Z�+R�z�V_;��7e^�c�D�N^A����F�����8WL9�gT�Xo~�N�y�l2d���n+��z�V*������D�S9�h'#�M��g(�U�+��TF�=�$���c�2���-Mx�oi�S��N�W�MUv��.��ἥ:�;���L�sB��
c�.4d�/��S���)�NN�30�s#����oQ��0�-��^�Qm-���^��I?����`�GԪ��W2cǢz���UMV:Q;7{�n���Ƥ����z�P]>ܝ��6��NCUĚ�\j�V��C`�4ٖ�:���s���
�W;:��1��I�r����HS�7�NS�=��A����j�$��3�B {��w	�Կf\���z�>=�*�|��b�+0�����Cذ�+��4vs��@�t�7�@n���Mt�
M	�ׅL�*����<ER��S�5mS��d ����I6(��/6/z����7�7�`wDɴ�3�9	���I��5�Gg� ��z���ٷ'�.��r���@��muY+��f��EK}�*j1��������F^ͭ�"~���p]�����Z�ఞ�j�P�Gκ�9�(����*�z쩨-U�d��L'M}S$����cV���J��fn_
A�����Ό���:��2�\x���F�FM���*�d��W��w�*�{E�v�#��ֵ{�I����+�u�c4uˋ.��qW6�x�vwhTR�S++9ň�wT�w���eƻ)�y5*�����Z����-7�l��,�h�!<n��T�0n|�S�]�"��wKm���v�k�V2���[{�Zb�{b�WK��谒�s �DXc��9���	G/ݹ��}��x`�:7:�b'c,kLCI1�����!�VQY�##���S�������*H�;P�!b��+�^Q;�����E�wHsu
��8�����{�U�RԭY�V4��Hh�3�1�Y�,t��`)�����5���\#�N�m_>}���#G�X�Cy_5��@��!��S����S��VZ`tn�*�lKnґ�q��R�ǦQp���-+��>0,K�df�*;=q.F߉v#&�<	͛�r�=ݽ����X���~ �O�ԟ�C^P�:U��'<5I��Du�;=~�pv�"^]6x�kv>�$�o�1�j;�<�X�-����n"S�ʹc@���d�^m�F��s/w_"*�\�*پ�`s+l�:�}B���+���0a����mHQ�}�هvI%p/�˯'�M*�n��u�VfZ��2p�&k�#X�% �ʪ��<��r"�+3��!����������Goj�C*6a���K�)�tr9��guk�J&F�%�$��J��o�O��ĥ�'�f�k���NR��u��n�v����քU�p�A��e>����i���J���_4�Ĺh��\�Rǚ��r�Dҝq�}�q+o�"�������������\h5~��l��ђ��P�mg�.j	Q͸i��a�M�l0ʔ�ch'e�)��U3����7P�,)�����:��h�x�[��̑�.����'ԥ�G}#$s����Jf4B���V�i4��:�[�	kK���.���w~�-�����[�a=�ᐸ��p&[P)�1�\�nE-�K�^�?r0��+��^�0��b��LU�L
U�lF'�E�Zz6T;l���Vw�qr.h�	ȗ��p�n���D��ȁ����!�RwjL��m��+�i�{�7K�����!���B����W=l����_Nd��X|Əb�ո�x[9a;�7K��Hd�p�H���Um�tx�%#�ܫ�ƍi����8��F�
���le'�Ct��v�v�+��{�
���k��2��G���٨��gl���L��֊�=Km��z���2av�Fhq2�@Wo�E�lu��,�0t�Fp*��=��+a�����"⬚z���yn̩6�G=���m���D�f����M�b�)G��-޻��w�+9a�5ۇ*�}�B�4S'g��>��S��xLǒ�M��-b
Gէ	E�6�OP����U��p�Kp_=}�G��{Y�ؑ�\��8�EҥZ�gs��٭ӆ
��˴�c[�,u
�6��)�P%����E��P+vwS�NM־�o3��vu�3�4e#�7J��U���1�Z��6��j<��x������4�R�Hق��'7I�,p��տ51-����ʜ��=U�x[�Sy{;�2Gc)������26U���xo'��v��Ll�+�+�M{�a�u�=Ԍ/������E)7��ns�c�ÈD�spɩs�����4林K}ʢ������h~a�Y��Ís�_6���%��}��ks�r���,r����j��˅'��mt;@��6��{1,#��hT�H"V�Y�򸻈0p6�:zS�tמ�`h�� D�l�^!G�=�wI��.'���dK��O�$OJ��=�i\ni�*�!�8��!t]Yt�p�����û����Aј���qQǘ~��e4���˵�(g��o�x/�,z2���wVv�aW��:&�T<n"��\�
OX7��sV�׎��q�gU*p�#���[����K�y=�lf�h_q�t�����W�l�U��p�W�^L	}ŐW�Ž�:P|j���+��1����S��7Ⱦ�F"�=����vd�]����f�Ȝ5��0���^�xv&���|��`���I5|�d��H����:z�h��}6!)w��+���@���h�t'l�>^{�V�ܖ�� s��N~�}�v�{�s9:�v���y0yʆ�F�,z���j���+K�o�d̼�Z��8{�t�Va�YĎh�y��1LJ+K���1-JY�������˘8�5;9�2��Ļ����L����Xu�o����r�Ttt�R��Ğ�*.vtD�n��z��w>{�@{�V�҃�3p�d�଩�e���Uk�~�ޛ(���+7��q�#�$��[���������sė
`���^6����敽c�=v�l���\*a�F�n�b��z���'
��}s<�VI�5\I�k=$�pd��Q���>Q7Rg��o�,��\��eF�Dp/E�Qs�>%�(��5�}[��wA��sTH���JI�m�.j���s�^WZ���IuO�h"j
���V9W����.zx�?R�W0�qz�r��l��4;���U�Ɵ(��)rҭ��"���W��7��k������Q�{�NT�E�+�b�׮��ꔴ�Qt��V�ó�ZN�d��2�X%�!�+��#����1�9�S����CqB𗒊�k���G�=�q[k(X��4�f��uv�I�D�x�V�M�6�\A�S�Q=y����p�o���U�nX|4\�1��Ɍ����H#ý��\������n�ӟ8�E��6������I��5����t7t����q���W1�f�e #��=��S5�g���yFTױ���Z)���Χ�����N�䶉	��-��3�jr��+�
bU@u
&���V�a1��*K�*�vFU���J�e[Ivf��<�Ř���s�����5�K�#$��FP��P�1gb�<0�p�^����@Z׾�?�z`�^�2��º]şE���a�d�4Ct�5����Qᅹ=͖���;U�_��b'|�,k1$Ʒ�bJ���r(�4$3��cw7���;\�UwB������-�
�Y�:3���3����+R�a=�1 ��=Ӛ���|�r|��[� i��Q��1S�B��"5�.�1c�׉ṉ��9x�I/v�K�b���d��.��0ta,H����y��5�PT���8"��M5]
��+E�`q3{o�Ӣ��J&S~$���,�'PV��R�:<5=XV����R��T;O��s+�^]�38��A��p�����XI��rn^E�(p�]���H���]�FF��.��G2��__����������	/�����;�m<����n�9��{ʱ�fs�gU���.塚=.�ޜ�����?�����	n��~][^z���#�6[���ܻ�x?=;]`$}���Ly�5�	9:<!X���
�<�GC=զҨlt���9��\v���*p�=1�L<�h���1hyc�����3~hƁSyՕ��1(��A��|d���H��p�g W�̘�1��F68��乹}o�FH�S�W��9|Ԝo9�R7�.�����Ur������=c\&�W�'�ط���}y����,�I��Fn�[-�=;hޤ>�3�����<�e鍏� 2��-�+���罻ii&`hS��5s�g�Jm���Y�o��9�R�.Uq�;�g���y;8Ӱ�o>G�W&��������R��aV�Ԍ��Ar� �*g=:a	��W��!��s��r�vv4j�ҏNE��^)\]�m�����+���W�=�ወ��e��ټU쵐�QH�i0��o�+��E�kL����4��,fT�����۸��Y���A�3�R]���=認(?.3��P�^���[�t>۠�y�����=��P�{���
�}n�#�"�㣐z���3�\&��BR���pp(Q��t��n���j�X(]��u�g^���q${�#X���tsj���굲�y��)��u�",b=մ:h��.X�ֈ��%\d��<���w+����ܴwz�}Բ4�k�k��<Ί��Vvo!}VEIV�����W=l������m�]��A_��zO���#�=���{��
ϧަQ����[1Վt��WG���ҜK=�S��bGE�o[z��X��*�UDTD� :���=�8o�����+�Q��MS;fOX����fq_7�fyfU��x0��[�ƨ���ʑ�=�֣r�E������*ə�kh㕞�N���<+N���v��u�ve�
�6�
Ky�����f6ݍ��w{�Jĭ&��g�=��jo��`������se�cʏ��9!#�X�������KL���0m��N�&L��.�e�n�3�_7��#�rgkv��44KK#z�S��^���K����}�q���&�����=0%`<7�.%��Q6A�TJ6�]��kz�/��X�K�(.sa7y7�;��u����K��%(92y;t�2Չ�)��Jx��$`v+Fk1;�U�E�a�>{��SE�^ynD���%��r�[�?�E�Qgr�KNpL+�ghk��7� ]���b���淩u#o�TS2�y�z��y����SA��S�
���5ۙ���KA�WQ�e֩t#ܹ1���}:pv����GO��f4�Ut]10�[�=	����4���b�D��((�U7Ҥ�����S��/!�4�B���5Z�r5k����U��Ul��Y�6r(x.��D��
zjm�Q���91��\JF%y�ד��m�ѓ5NPb��j1��tH��sVUf3�׺�oӨ9��@̺��c�|� ������jL�C�ӓ�z٘��e@�.y����X³;)���*o^�*zo�0[׼���W�+��ӌ=���2��.��U�G��D�V����7�Ԯ�o{6�8/ڰ�9l�/���=E�^1����JZYf��`��o"�VTˡ %��O]�"3�m��k�oR���Wvп���Vj&P�a3��	�`Ô���t6Z��4���f�ڴ,z�[�K<�c�8�瞏JխQ}(�r��o���i����)�~H8y�l�8"_��O^���+�"A���a�ծ��o�aP�Ϸ�����)y�:���]��ղ�)����L�heҕ�x�|j���R�r%��]�����{</���h�uv�+��o'�Ge�iU����M��)%���7�W�Rr�ؽ��:gk)F��n:6��mC�EB؂����,�,Պ�wv��G��ؑ�Hu��A�g1LR��7����o*��\7h`�{r�ē��X#���U|B�TO1Y��ʻ�d;���[�8�ޓ&!}w-���NL���;��B�j��z��]_ �k��o�{���fwP�b�gv'�QeFo,�)�J��)\��n�y(��i� ��;X��5���n�;2��*ӫߢ3��W3Q��M]&�9�.��7]8p@L����׷Y�,uv6��Anvݚ�N���}5�׫u��Y��.&ec�{9���j��o4�^�����Z��s�=���U(�7F������ۚږJ�wFr� ���p�����[m�Ae;�*ub6�$�4�U�w5���\���A!\rU������(*����mVd�XU���\B���KĖai��w�	#�v�*f6���d�^�h�����o$0vۮ�X��̎�ρDFW���Lsn��c����Eӣ��f�����{���*:��֫%�%�JT��aTJ;�a��P��4�Lh9�=��P��7i츗4��K뇸bui��;g9�`BTn>\�b�/�0�E%k5�P�s��G��&]>*��ݺ�¥%�bziS�]��#�gn�WWו���F�h�\���њ��@]���L�]խZNo�ھ(nH�vQ������0nQ�����H�}l�e������[C������M�\\�W������/V:YCP�+��7Ms6��)x�E=��(#"�o-�aP�HDlU�<���<�b�/*L���7�g=Q��L$7�y�W�|���M��:���R:8訥��:Ju@0���t���д3X�=D�89���������6=A�;}��]fĠ�8��B����O�S��li�\&l`��95RJ]ϑ�7sGk�-R�Y}ÍŁ��:��ǣ�u��VLOH\�j]�cYܝn��sUHk��d�9��Bc�JܥYk5(N�j�곘/�e�㽊Pݥ)(_u�V�;
�5�1�X܇c�+���}�n>'j�˫2V�F�����c�䱝L�&!sVL�W3�����~�Sb�*97W3���/Kو#��̫�r�(n��'�������[�7U=�B��Ҍ�nky�}��w(v�qd�dkmG�Mˀ[�����b��ʼd�)8�-5K]l��&H�*$��O����i볊�|���w(��Rxn������z�P���+�yV}����vh�v��c���X�l�X��ǩ�/��<�j�=Q�ڙc�����Ρ�9��f���R�d�4v�Z�ς�C�\ӮIY�+�(�ݖsZ�ى[��$�n=�9W`� ��y�Ys�:�u�<���n:�j�\�w
���jky`����"䆌���\��� ���R�)B�'�\FX�-mam*�b����E�T��*���TQ�Yj�mbʲ��jZU+mm�҃ʍch�DF��V�F���F%����+\eTšlk-��Z*X�F�iV���G3�Fѥ-���Z4��kF�[R��j�JѶ�ж�YU
���*�%���\V�E�m�j�KE�4��Km��AQ�*�,����ڔ��kVV��UF1��ţ�m�b1j��4JʩR��(Ԡ�V-cr�"3,���h��Z��Am*֍ih�ը������5�iZV�`��F�Z�V4���UbV։F�-j�Ail�-(%��TiecJҔA���V�U-�e�jѥ�Qe*Z#j2�* ���Q�j-��ikm�*�m��X�iAH�-T�b*ڲ�Q��1Q�����b�����+Uj-�n�XV��NB8I�A�N8Wa��黻�6ێ,H�WyPM� i�.%���)8���D��v�S8��f5��7�%��'CG�˷��,�d��oM`�}ULE���`$0��������[5	�KD�7�.��=�+��y�P�z/�EN��}T�cꋚ�[����f㚢F\D�JJ�2m�o�����a�Gf'�F}+D���P�3Ѕ˞|�籘Z6r�ir��p�ü[�\�Y�Vnv4��t>T��ծTޔ��*OWw)\���.T�kO�� �,b�s�-B��`���g��v�Zq��,wD�zХ����C^�@��3�{_n��|��+�����Sk�j�,�g�8�=�������)�X�Y�-��y(3^����Xgun��٠^���=)��{mKR0�)�U�(�����{ihȠl&+�M�s�<qZ��v��U�%�us|!1�vV��ՙ�|)�0��ff��2�\K��� s<��n�6sR[C+���GrH�.��N!��@�}p��].��TO醉�AF\ܷ�vx�؟���<<���Fv�V@��:�bI�g��,E\B}��ٳkJ�l��zR��1��g��L�����ST�:�NF3�F�;���S��V��5b���)G;�ff��LܽE�R�+7����\r����L=L6���(e:zٻ�oo�q:1i]��a�����73zK����9č^�l���/����J�To�r�_���/�Z#pEt��)ќ}-���}�lz����=��߹���(nJ�Nc�4n���fR(wQ��}��+��Ŏˈ�@A��$���N]i�ݠ�u�+�s}�M*�k�׹�a{���W�@���6�8'��:MWC�Z�>�l�U��;��^��$Bi�Q��5
�̂���D>0,M{M�k�d��x���
�a-%�|jr�s�W��=x������C`	�ꀣ�P�z�&�G�+���,�UK�o�ޚ/5mf<ݕ���s�\�hE�րe箐y],r�X�-��X�&�)��f^8v�Y��C�K��ɂ��FN\K��n�l��p~��La���j1�J�r%���0��rs���(��(��gN������������VfZ��w
bf�F���J����#�iuj]W\��ٜ�C��\���ޤ�!��G,<ᇄ�j��,���;mM�|�#3�y��ܗvHS-#��r����12��c�%)��NO�#�L� !vm<��Ɇ����s�Ŭ��r=dɓ��v�)im�c*�h��l_h��*Sof�a{8?�&/'�y]�!u��S�Ւ����^�$H}jO�M��+-�w��*tYyyC�飣��U��Z:ց$�w���B+����\;��Y׊U�+/�oy.�����!�3�z3�\߱�����y>�/<­C"��^�5π��`+��~ZDǛ���&T��U>���+�t��I[gg#x��z`l'�|2�1������V��,���ʄd�c�1�&%�cG���6�Kº�fy:��#�N0����|�D<WM̞r��1O�fp�A��Ə��	Ȗ�\"�&}�s�[��{�}�Á�MU���xB�	S�����vS�w�f�4�_�����f�o��W=l�-3U���s���I�����Oq�֫pNhpr�r���a��7R�ߺ�IH�f�\�W�8�����7;��Tx�=Wm�`�(��{b�v*+c��SM���ѩ�:r��:n��v��wf�ʋpN��-�l�ӄLʪX|�;|�,{}�Ś�R�t��!<��t�ȵ��^l*���d��|2�׭ٜ��6��,1�)Y��+TX�G>��(�_�m#�xt#s�����5������c�C�G%-�/��3$�gCЫ�Qڑp���u�v�o�`�����E�Aϱ�*�΅N��{3T�*Ɍ�%J/�0���:��m�=���q�3�Ӷ���bVWWo9i�:Sjޚ�4�=�RXFus���p�=C!�.�i��+^�M�o��J������T����|1�g�yR����g�ZK+=��b�z��7���V���h�������9��G�3���,�X'G�'�loJ�Oeq�ʰ�q	���]�|�@ޜQ\�Lu�oqG.X��n�0t���Cz��w��9=����x/��v��v^9'�gs�d�8Z���Y���A�o;*�R�QrطW^w��Jh��[�"����O9����[)RZp]θ�g�&aN�2���<o���I6E=)��=��2�TL��b���bRp`$P�:s1Ø��e� y"D�@S�SVҺj���f�>='4z�����7є�hW
b�NP�~�f%+��O`M���7M(<'̱����7��#�k��GV�8�ű��ۓ"t��NLLL\��r��OX7��sV ³;���]L�0վmf�J�g��Ut�B�0ń�lBR�I�t W:�2���F�z�1��[΅�g�����=jOG�=���nu`:g���R�����yʂU/7~7��fPH��y6u/n��de�瑗���+qi��t��R�w�M��9�,�_��R�:���?�xݜ�xzL��Y{|���{Ss��}���<���\���*W�;�zK��3�r�.af�l�+e���9b]@i�-�����fVΔ��5*�'�D뭚V41��A=�kTĵXK���1,)K"Y�=+�9���=���1��C���c��rf�lzi���˩Q�ҁJ���b�5��UgI�d��:��"\y�B4L�����q�&����#���x��ޞ�D+H�ɋ���=~��qS0���|��&k˘˃mV�j�*xçT0���J��k��5<:�����Ԗ-��_�\&fu�:3�G�Y,t�zk��qi��ZC�`�6jkv��[�U�˽)�v��}���k�L]J��U��	�Y�՘�g�A�g�s�\��s
�Js�z`+:Idc�.bxd�����u�_���\��ή{��f8u;�'W-�䣜�cF�Cy��O��?=����m�����vyRz��J�jb���6�Ջ-�J�XSS��f2\*(^���n-8�ytL�����D���ƀ��T[ŕo�/y����)?0���ʅ.� 8��
&�w+�,c������C��.��7ƽ6�w�+��vo�Z�[R��3���z�0]���\��˫�b� ��-O.�}�%�o��gk��I��.�����oy�8s�u�d*JӺ�����+�׵�)��a�����J��s,��ufkM�u��a󓻒�J�]3�0�a˞�g���Rt�Į��N���5�Ǽ����w�Q��d.A�ܸeP�������CC.0���0�W)4֥,dd�<՞%H��}�ٳ3�ڮ`]��iδ��@�z��`�W�K0x��ŚÓ��z�ݏ �'n״�ߏ����Ol<��fj,��M�����Oƞ�by�KT����yY��_=Ɩԗ+g��A^��s���/�44xZ�Qύb�*�KD��{>�t��Z���v�1����q΅F&�"��ˍ_�:R`4�¹��"Zσ:�}o��t.p�J���o�^��Պ�"�,)�]P%�k�ˉ�s�tQL���=9iZ��b�
�/!���V3ꠡ�u��/����� ��K�+E�x�0:<5=E-=�zLɚz�Ɩ��ܹ=�/f>YN����%������'�P��BM}:<!\��0zN��^��{��.y�T�
�]JK7�Eek�ʽ�X��p���U��S���y��v� �+�	%������v�`RQ���.���X���}՟>���:����z�n� �_[�0���%;�!_FOp6`6g^��Ʊ�s{G^��]2n7�V��	ֻ���<�J�����k��跊��6�}]+A������wa|T({�j�%��A\{�G�i�g W���La���j1�ĭgV�Ϊ�nJ��or��Bdʧ��2o�Νˏ��cs 1�B�?uߖ;�g�ks&#
be�ꊢd��Y�mY���.	�����
W������HF�@u���b.%#���k`�Ǵ�Kv���*��c.`W)\#W<��P�ch'e��M�(�(�,�ڛ��<�>�u�5Y\�U��,+��a�TF4*�R��­A�!(.\���2-U��:<�-^�J�#�fcl��rfP��J�Vy{�<�jIZsz�\���ɀ�E��O^/S~���dWJ��⫀_^�%P��Y���cֻee���\'�;/[9o;ӫ&�9��߭�\��ʾ���(�/���P�^�'"X[����B���:�g���\҃�̍/��.؂q:r��Rf�LE�qE�̀�N�([WSdl�ϡ�ܝ�N	;�;Ӷ��xK8x��Z��p�L�����r�y�Eܴ��/vֲǔ��$֏Gh佻��A-v��'�b�J��O�o=a���F�J7�]ژݗڀֱk�l����gV�-���ľ �L3�oh[M�Wz�09��ɾ5��T�|b�H������Cp=���/�뼹�M�V�ꚳ�~0!(]�I��ě�8aEZ=+�Z��E�o�UlT��{���V+;R����'����:�捘{���ТY0�{P"mk��C۾�<)��u�_��f�TA��3ATtpZp�lyhʇ^�f_T^��(�B�:�v��q��J���<"^r��ͮ�$TJ����N陵њ2�¶�������CvwP">B�$�N��j�SH�Q��#&��`�p��l�F����
�̻ՍLKlk�(L��c���z��\������b�>�p�ќ�N�������;����U�jW���W�����3���=эʼ~[[b1�	��y�D�s~DԹ��\��[:��p,g�S��Mqs[����Z���~Ok�VЮP���'w��>��r�N���Y���>�r$,9ǵ'm�=`����X(x\~lW��
#�������T:�R�g����헴W^o���\��q�E���E *S~[�=4��M����ÞT������@�[������XT�@�۷u�->���+P���2��\V����1��a�2yꈘf`j7q:z7���;�rF(*97_�l�o;�A����3���u,,NxgU��LL[��q������891��d����z=��d��n����%��<E�8�+� �֣0z�$l.�5`uVa�g�i=m�v�U8z��+�]�Iv��s����6�;rf�k\o�C@��Q�9Ar2sn�ğ�o(p�y3Fwl�5hc�c��>V.��Z�s�}J���N��G�X��IЙl߆<�M�t���éw5�z��Ձ�nz��L`m4���!�6'��7�c�r�]�=7�)�ͯ<|c?fxk#	�C�gb�N,�+�3�v�N{C�4X
'���=e�ڵ8�Z��-���M��q�TeM�$I:��93b�=6��p���Ԩ�J*��b��9Ȯsٓ.x�/>�	���@��2�v��ϊ�~`5au�`y��n4�)����5���$��vK�ffEL��D�C�2��5ZI���)��`B�<Ҹm+nofz�*fw�s�Ա%�A��Ӟ��Fg]ã>[��o+$�5\I�6x�`FN����;�"�^�y�!�zim;�@C�}�'ʽ����>���9�.�=ъ��e��}�<�9	t�j)�D!��dv�v�(^���j��97��7bf�Vt�W ̌�~��G�蕷����LW{�n��i�^ZeobٸR�C�ҺT�X������:�v��n38�C�MPN�;���.�M���pTj-f�)��U�m�+᧥W��Dv������V���NM��qT��`Q&V�Ρ�
�;ϝ��\�ujjL���z)�R������v�sї��|T���[�
�V�����<F��S�������>���.y�4�^Ip>�3���N8�E��%�tE��&�s>�rܼ�xJx�{����%�z�yQ�吃�Ss��c�5]��1�Ow��Sȱ��&I[�{�O�Nw'Ⱥ���ܵ�*j��A��1l�ڜjN��B����(�G3�=�84�Mz�n�}��ۅ�`~�.kŪ��h��`�X;Vf�/�!od��L�]x��WKIeIŭje�z��`;�`�2�mQ%���Y�y�к�xƟ�1]].�܁�F�F/](�ޮ���ټ$�)�h�p�G�3ߌ��N0��XI�p�cXt�p|���"�ي��y�-g+GIWq�
5�Fz�:���#%���p�/b��B����~w��登	��1��t�qf.]�k���P�w��k2!V[���R(��s���&'�g���M���8��;�P��x:���ngsк�[Y@nK淭kE�N�ѩ;���đi�����+���\�_��#�w��.���D��Y�tnK�}}TXwȤ9�Zx+	ٌ�xYׯ���r�;�����?/��6�% �4�8���]�%<�Gn�8�]w�TeC�b�ݛcH�m�y|���B���$P����� ���]���֪�,��h����јD����z��~UI�y�t�:m�V�"W�L=�N+w�Y����I$����ʺ���wV�y��d��iK�����-�[��,] �q����;��F��2b��9��XS,���R�(!�zL���`wr�,sI�6�:�Y�t./훺v�sJ� ٬5
�:�E\XeP	���fC��f^_VP*��<�_�ڣJ�H��T��U��K�Ǹr'K��e�å����e��q��6���Ο ��nL��p`��z��9�T1�*���ӥd��w��l�x̷���6�Z�a*�kNPĢ��Ժ�����n���\Tufg��FqI�b�j7o�;��:�G|�r�F�+���&�v�Y�+�D'��8_�Vv.�o��[A��Z��*x�Q�.����Ifk
�N'-jܡQI�&)q��	��gF��f����l�u��8a��_cܳA���Gx:t�5*�pp�0�\kn����g�v����۠�%�۶���vV��J�ʮ�Jpp|"��EC���e�kǪ(��a��갸�n�+#�4�]�A)n�)��B�Fm�Zk`r�ۊ.m���)7�a�Q�Ҳy��#4�$N�oVA#��/��z3Rø�KɈ���ޫ�*�,���Sq��m� ���ع�ђ��Z�"{�м쩩AD�"�澭v�7�2�ФjV	��_�����p���{�s5��趕�n���o��X�1��էij���i>�U�b�����oT]�RP]��9�F}qR̳����S#o9�u�)-ϭ�髒7�����8�:P�h�gB֬��܈�黏����2�G%�\Na�\�J�S+`Lv��P,#YWEѷҖ'�R$-���5���������t۹��̻A��K�:1�ȕ�]�]Ӂ9�'i��S��z���PN�i�e��bi��m�2\�'�������}Ou���V��|2�R����W\��Ag^�zb�Ydi��Џ�Wt�B��8eL��L�eL��ÖJ���.��dR�����g��K����>�;5��_��^c9�����@� #g�Q;�v��zE��ۥ�݄^7ݫ��4r˂V��8����\V��!b)�`j�ЧO�U�y���d�ewp��X�nH3�N��dm�:~r�WE'7�\��Էm�xH��/]�E�#���5e�[��|��7�~�K��PUj4F6ԥk-����Tcj���k�R�Qmcl�-mVT��V�*Ҷ�%���VX�h++k��7�q�)jTcjR�--��eF��)Q��%b�-�V�Qj-Ub��Ѷ�
�Ȣ*-�T�j4��DB�T�+[m�Z�+VҔ��[Q��b������m�iVVQVV�U�ԣR�V5mDE(�[kQk[EX�[EJ����$F��Z���֍FҢ�[b5Z�Qj��b��EE�UB��X�JV�h�����DP-*������Z���m���D���(�(ֈ�6Ҥ*�-Q-Z!hUX �,b�b��F�5���EE[[V�QDDAR*,����lE�5*6�@��V�TEUb*��"�PV	e*U�m�B�j�Ԣ+���*���-Qm�E��AcU[e�b���+��QATQaXرJ�����(�hX�*�R�*� �T�ml���bdDPPE�TAJ5Z��1Eb(��UTeV��,�UUUc�"��R�TZ6"�5*��EU�kbҖ#QT��m��x��oo�թ:f�c`��%]+���p��[���wc՛!��9�yN7�ٌS/F�T[��v��wo�g���G�71��N���$?�4EGq@=P�ua�63���c�uf���Cpi�]ga�$-���^��0W�:՚�#�7I����ǜ$��,�:��g�����^�뺈�d��K2�k��30w�V:Ȗu��p����u�C��>�ǝCLz�&����j��W��۞�5���;RH}d���N��pvQs�m�s�+��EĖ1��Y�9�F�-���<�u-��R�s��J��Y�h+�9��	�ߕ���UyN� }�@��[�oe�{�qs|�i'�<Y���=ݜw�.<C9��:��K��ȫ3-^әjog{��6 �V�O�-��D���B%��U��؅*"�}�����n�u���b5��P0Y�䒍OX8Ĝ~�����u3Q���Q��H�C�t��Lm��*���$����C<�����{f)֚�Mc�`�Q�\�c-�q��
�}J^D0�P�jN�Q�F��g�����x�d@I���ʸA��U�Ҿ��՞b���IX|7��k
�_4�'���i��މC�C�R���u��t�-&l��Mv0�Mf�x�� �sHk�g��tᖜ�±}�b/g:���������˭d���v�b��<�-ɢ�T���=D��wH���P����L�_�t3t��43�mN^����ص��{ވ����ܦG>�;G܈��pf[�aL�N��cG���(gz�˨+�6lrw��s��r�^q���(��z`R���	�:��QK�cG̡9��p����ؠ�{���U����=���ۊ���-��);�&l�LE�qE� �a��j�n�z&�r���č�d4W%P��<c��m�k�?S(�čׄ�Q�5>֘]�x��[V�ʞ۞ai>qw�O}[��8��EP�e����D� ׉5��U����V�\�;6Ჭ�]�7�'�I5;rұ�U�hXw[6��ZDcu�Z|�����,�:��Z�eN[{�]S��.�ɞ��_o[��Q�0W7�o�E�2��5�2���=��K���m��+�;o-{(V g��~�՜_a$o�����1���x���¶������,�O�gr��Ow��.9��m(�Ǒ�}�ي��<I?�=�(��Ɇ�x��+dsW��� ��]����L�������b���;N�_��Y7�wdv�1�Mk=$��L�G>2�MLU�+�]����_l�%'���b��^���Tm�@�v7�ᚯG���r� 7ۓ��K�h�)u�Y?h�s�޽����3�bDf��&n��ʶ'˴�Gl�X�s!�:jâKC� �r�Fе�n�8�t�c�O%����W���؟�=�{ܭ>�
����t��߶�D��I�u��T��MK�M�;U������nR13S��uR��R�-tmW�0���r�Q`��=]A�A>O�����3}�j���9�=���Xy��p ��k��
�+ADn��ߞs�P��w!CP�)��..�����xM��8sKH��p�@
�����eY�/��#n�y���]�{{NOkT���=*�=..��,N8�+�Q޵��z�$o������u�Yɪ�܏�3z{�5�R�vl�X��-���h���7�h�� ��0�5'�d�n�,�����r�-�wl���*�΢VM@Ҵ=�^��o�|�˝�gd��>&��{��.���>�ÀT}:�4M�n2��9 ;q!1Yr6�}�:����� ��n�:d�A%��1��{%��7_<��{s�١y�@0~��m6F(����4�Z ڞ��esv9�U��<'��1����"�<Ŝr�<�zj�P��:��(:����lr:���X@���]]v�dN�[�&z47}����C����+.k�bb�����η᛻:fe)˹�k�q�Ž���hv�ŋ�LZ�Ы��A�hw�y�<�Ӈ�U��`
<g�W��讨Q;ko���f�%o�����D=V�>�U�r1 d�O�] R�gDJ,�h�{�
b�Ն�k�����:�rA�XƇX�k�T����n9�2w�\��_��j��*z�O�PPÛ����1���{å��%Rؚ��}<�����tg��:�<�Z��Ww�^gb����m�$���6��tr���ߏ�H�{P��Z/�Eΰ��<�ͣg�Plq8oۙ�����'�74�/RFx{��g%5�CK���+�и�Z��(k�.\���qH��l��h��ܮR�3�g<�kHY-WN�K/��O�a�qZ�� ��Ҁ��*A��u$&��b}q�Q�K��Z�r�"��w<�pG^I0}�g`1��Ԫ���̷q�f	�W��B*��x=ԗv`"gwJ�0���Tvy)u
TN�څ8�I��c���1���#��s���4�Gw}�RX
�V� �[)xua�Jb��S�I��)�TB��}��E�9��;�2�^���7�Z��E�R59��e`��ՙ�K�H_�����r��.:/�HB1��Y)�;ۣ׫~����/��z!���j,ަ��uj��b���_����KI�ߪ�-�Y�jлv	�����K�ّ=�	bP�if��6�!�ON�\��r;�t����X� Ɓ�ڧzz@��T<{�UW�i%%*�����z"!7�nF�s31xl�ɉO�&�:ui2�[V`󯗺`�W�A���T钕8��[����9�rs�:6=P+�4{%�h�,�Q`�ش��+�U�'}Z�6�G=1��!�w�����g�u�C<��^U~B	XEf4��4y�n�{x� ~���˷��<�O��D���˹�yjU�#��ߤ9��y���A`�ˍX�JL�<M�l�!1]�[S����!��c�x:�MA�vs%u@�5�u9q7�u���Q�/��6����6�G:�?�I3��"oEك�K�S��l2�(k����u�������@�Q�:�;%M��Î����9���6���==~�
�@�f2v���;c֑����1�P���	)���gr��%v�Pq�-���}Y$���$CW����XИ=d���,{\`�b��Y:�n��Sn;�����������&�;����{_Q��*����M�/pڄ�CLј9�b���ǟ�+��z?[����+6gX��g��K�v���j��dބ��~�}s�K~�q6��Y�G���:3n�(!{���?4�o&M�	��{9w�k�����[^^�1���BF�=���Nr�:J�T���r�w.�n���<�q�R��I�I��� Vf�HY��[�����]hs�C%غ.��aE�d	��T��
�^q�z=��{�ϗ8o^$�\��y	���G�H����؅5���u�O��6���,�QMv���輯�s���h5o�ݿN&fm�0)\B5s�b.��	���<򜁝*;�+��O+X�mML9��0�m&�AX(Tbusx�`�F4+��)x­BR�CAkG��3r�����pCl�-	<�>�U�O�֠�\�ع��Edim���.br�G`��-����u	����]�����e��*�
��"�/�̠C�(<{]`7Kuи�H[bs��է����2��o��N���A��X����9����iZzP9P�N�����8�F�ߏ�|��C�z]�ѿ�S�y1U�J��ç���=�X��N���!wx�;���_�s�>��d��>�l�9�i�'P���hu����!�l�u�A�y�d�I�{�I�u$�s?jE']2"�Q�T�A�y���3�vg�ߧ�g]���|�����C��~�����2��8��k�	�:�P�{dXN3��ɦbCP�a�IY�<��8Ȳd���2N��w�ԙ�/8�{�_�~>����}�Ͼ��d�O�`w�d4��:�3��!����]��m����P���'�^d�����{N��I�x}O�4�d5>��La��C�M�ֽ�����������}p��\��T�ԁ6w�.RW��HB�R�pI�[�:ܭ�@7�A�uzP�?��`�����ۼ��Wqs[����;ޝl�|.	��F��6{��;wJ�vqt��5�],�ht�b��k�v�#��u	�r5�����"}����_��<'����x���3g7�z��0?$1�]��si!�y�P�������g��g���	����4�N3��&?�Oo�~��w�{�w�>��}�{��i�d�;7@�3S�ߒE\�tL!1�wy'�11����!��m�l̇���=d�����I��+=OXN0��=��o��ٽ��ƚս_x�O��3�}1��9N�)=x��P1���~�o��>O�LO�y�|������Ci�^dXJ���z��>@�k��g<���6mw×Mkz�c����'�f<'�1���zȰ��~d�CiY=�$ٻ�d��O��I���w��'����C�������hm�`y�rm��b��1��H����M_�C�)��g�b6}����M��',=�N?0�&���>�$�w8É�O�5��!�?�w������w��>d>a��k���&���zw^o�3�i�f2~G��$���ya��$Ǻ�̞<H~Շ��&ݳ�i u���7�$Xj~��>z����a��'��ćY�=���{�;���t�e�O��X_Dz�ޏ���B�t��1>��0��4^f�'�O׹=d���sL���ڡ�"���������������'L���w�>���ڿg}�{��1���N���N��v�$6�nw�+̕�$��rT��.��N2)��!��I�~�p4��hLe ~�DZ
 �ܹ�W}�薖���g?}��矺m���)�N���l��:���܇̆��;w���0�������I��E�I�㹝�N$SP�d>x�T<�d=I�hO?~��i��o��{�}{����g�a�x�O,!�.ް� y�>g�!�z���g�M���N2La�w�I�6��s�V�W�~�H�,�x���%@�lþs{��޿�S"\�ӣUe�q���KRFV]�tI@Q�)�Ooo׮�;���ڎ[���2�2���vyq{�c9c���1�{�j��{7���j��(��:c]��.���K)�����Պ=�S\Wk�+�g_�au5KK�wb�Z	_��S�?�舺m�m�Vl��vH��^d6�����UHxé�?P<Hu�|�6����O��=d���t�Xzɯ9��&0��I����g�}�0��P'�k�5���J��6��>��O�������~��a�o!��̇�,q6��~�P�����!�д:��%g�yl�u&�����}�}깅�?�>��3r����|&����z�w���,�Ձ�oXM c'yO׸�m���m��sYXq=d?k�H~C��YC�q�힤�1��p��}>�t�Qa��|�A�$�gg�g}��8Ȥ��{�'�<�u�=x�T�9���N���z�iu8��d��'��:��&XzΡ�!�k�	��>��f��}��yϬ�ءm?���Z���1!�a�J�N��6Ȳo��0��>��l�|�$�']09�i!�:�O�̐�C�{V|����P�b�'��b��8}-�=��w勬���O�L;>����m�'1����H�u1�XdRW|�(���I��&3��$��&04o��é�m��� �<uc�6��_2�S��D�~��w!���I�+??$�0��L�����}By>��Oyd�9@��g;����{�~N0����I�`Ϣ+w��C������QĶ9�v��5��1�#�!�!�;��x�X�l<d������"�~�S�I�<�1���'���I�l����a�l9����Lz6>C{w譡�8ګ���KE/�i��c;;���|�0<�o�1������6�3�wP���|��j��?2Why��"�~���%I���O�I6و�1쟦<���~=�/xc���9�f����&�a�v}���C�7���	�Փ�=f2m8^�������I�k��̞<H~5a�E���x{d8ȡ�6�$RyO>�{���o�����k7������R�>��l�k.|)�3zGϴ��y�u�(n(�ei�h�Ů��ogO�<(�e)s��7|OG]�.c���xKT�t�c�Ƌ��e��U �9Y.��at�u��<8"�F��K�(2K�I��`�o�򪾯����[�o������d��	��vXq:���$�����{�!<��ju�����+%M^g̓���{��u��?k�2~x��5a�E����y��o~]N���|�r�K~�ELD\�}=�G�3�Xq:�c�Xq8ɾk�Chq��3�	�C�o'�'��'|�q�d��eO��}阸b:aϽ�Ϸ/�e��O����{�{��i�N�՚`x��Xi!P:����u���8ÏLw?X3�u���p6��:����OY���a���i7��VJ����h�߾�>����oy���2)�w��턨y{��'}��T1ěz���Ć�h�a��Ol�:�!=OǶ�q��x~�ta1��;�I�8�~�;���gs�{��ֽ�wߍ����a�%t���E"��}�?h�l�h��봑C������~���8�!������a�C��ϙ�:�~O��X~d�ܿ^��ZνoB�����g���=s�>�'��Y1����T�'{g���*�R���ԑC���u=B~�R0�|��E��?{N�=`o�ݞ���י��㹾��o�͡�'�;-����M皛a:��;��u$�s3�E� y��<`T�ퟥ�T���:�a4�ɚ�zÏ�Oƪ��C�p����������w���7�rE	�~z}N2u��q�����}l�u���c$�'{�'�%xsY'�N���ް�@Ĝx��p��������	��������ϻ��vo�����4���	�י!������V���=d�1����u���l$Y?M���u�ϻ����xo�OY>��Tb.c�g���'�n�W��>���������}��C�N�����!:��?SL��8�M�Ԛf2��dY:�M�:�d����$��w���L�k}�*&�
��~c����ZOwG~�j	Ce�w���}Jup'8f�z;�Њb�m
�+��o��7G��k$�j��W}���V�2oV�;�̓PZ�K]�����苮��{˾�35�>�d_�u�	��g)O,�*�~�Dz"=����y��|�L*c��x�é�6�����]�͡=I���~I�|�0�a����i�0�CϬĝOP�Yԋ'I��&�I�~���w��s���sKo~��X���L�Gѩףf6},�sy'�1����C�m=���>O�Y�'�|���a�%g��l'u�����$�ed��	�3��zr�������<>��w�{�����r�����I�?sx��|��|�c?�I�>f$>�6�b��̆����;C�M3�Ʃ:��%v�P�H��������x�ޮirޯ��lǽ����1��5���d�i<Hu��ӻ�?0<�ޡ�|�|���$�6�0<��m�������i�d��j$�`y���g�����}�{�7��xȲc�;���"����H���8��l'����N2s)4��S��8�~�0:�P���Y=g�bM���ԓ��{���{�|��{ϸ�ן]v3l'��o!�����V$Y:�{Hi��5���)5��a��	�ou�2y9�'���~�u!�'�;�N��OėZ����{��ϳ���?{��q�{��`~aY*t�f�O�=g��=d���]�i��ć�Y�9��R��?&ޡ4��q��&<�`u�g<��Cl��<�������2��3�U�>HoG+[a}�)�Ɉ���D�����<;܁���|��$�E�/�'OɟXbN?��Y�2o�@�Chze�m���i�N2�/~���U6����I}@,�]�z ό�9�t�y0���ϵ'��	��aXz���<�̑dY8��;��H���wd�=�d=d�CP4É���x����tn������x�}t�]��LT�Ч�E����B~N0>g��s�;��I�<;��'��	��~ԊLN�y��"�d�����+i����E������D��6r�@��Q��D���}�?,����9_;�:�<��'���4ƞ�	��'������,a��8u)��<�*fi�V��
��Blv��һ�X%.
�[Òݣ�}�=�Od�i/���wu�!�֝*��_v���R���n���n�w(Q�O��{9�ywn]0y��Y���J��90<A�Z���k%��`��u�]�]��V`�Ha�m���Ƅ���9�j9�.�@M��M�APYx&N�ٕg�ۢ^�Mr��J4�a@�X����q!��*�w��l�r����C�wʹ<��f���.],�g�=���C�S%F&j���Ĺ�����ϓ��S�!n�h��2�jϋ�#�F�̠{�Vl���5�©U�ǂ��7����a��X�՞ D��Y��7S7��ʅ�&]��Z��T��u
{*&�N�&������tm��bY�o��w�_&�l��Kn���TY�Q��\j��)��G	��h���nX�cݥƷx]������Č᷐h�X��⓶�J���:3bhwd�ܹ���f�v�������f���o�Sذ=ݻ�Z
Z&Ɔ.�l
ha�j�8���*0�v�X�g3��F�M=����2�H�dy�Y@�ۓse>;�S�}��b����jNO���/7��J��}��e���YDVCVb�W'!óe�'su�y��ॲ��[�����8E��f�z���9��|ۥ<�F xx�{���ᖌ�4��@8��Qj��&;�w]��X|E����-}����ُ�C�oyc�o*F�@=6�ݛT����.�Ό ���	ï�EQ;$����YZ�������a�ȭ�����+�3�d�R���8�GGwEA�^��P8Y|�g��M�� S)&�I�f�k����s�0���˵�a�H�L��vm2��wWX̴�n��[ۣiɹ`[K�@��Ĺ+2�i�۶q3�9��c�6�3���5JUc��ϳ!��:gl� ��b7u6S��$-!	h�ޡ��a#��2�m�N��l�`�!m�f��U<{�Vk5��s�a�ᕓ z�[�f�W$f�u3)eٽ���
�b(��u�N
|�A-!���to�U����,g���/m�Eɕb�]HxH�j��,�[�s�!���Sb�}f��
��\;\��֚�f=엾�b�.Mn]b"���ظ��W0��<���3-�o@T��q��Y*3+v���#k���Zk9���I��V�d��3���ܭ�%�*	,��Փ5[��XO7��"�,D.Ri��5N�w��b�f�-E1nj���ۆ�R;:[l˧���V3G�)�鲹6�:�I�ws:�sFу�L�W��ztm�{���̭��dSJ����}k��X�;j�"����m�����!��+n�Xc���V!�����:ق�4�L7FY�9�6�Ρ��fV��� �����TC�Z#���7�Ŵ��pѹ�_�}c�E"Ul+O�AQ�[j�V,F���b�#���+j�b�Rգ�[
�%eZR���F1EU��`��E���Z�#
�()m�Q�VT����+E[h�Q��Q�A�Ebb"�`�TE��"�TDPm�ň�V()R�ZԈ�AH(�ʪ�"+QEDUR�e�@�F��(�A�X,��j"���J�F(���Jfb�J�`�QFҰkV(�jE�҂°Pkj(�)lbV��m)mj#"ʕX"#Z�U��P��E�h�UQd����"�KR�PTkJЩX)X�J�E�PQcl�Z��+DPT�k�������B��AE�6¢"���jQQD�Z�jPbƢ����EH�Ĭ����F�P��AUm���QXQ�
�B�Z[j,QE�j"�2Q�j5�҂�ږ���*hUB�+X�DE-��`Q�2���m����J�V*�(�J��J (�m-�/߼���\��7���ǹ7{�������iR���p�P�.7�S4nt�as4�r��j=qᱦ�7�X��W����@�5�������
Cz�����Cl�y5N��4[>g�'Y�=��u��MM��M�����u'�Y'��R,��ý�x�Y;�~/�	P6��w��U0��o5%�z�T�z�<���tƲ���<gY�~�,��q��=d�0<�:��Jϐ��0�&��5���<�u�=N���3��Ru����4�m��ѫ��w�z���;1���d4��;d�m����'����z�!�?{dXN3��ɦbC_�8é+:����"ɓwX�:�����o��������߾]�L�d�߹�zɽX���0�m���!�����N���?C�:�P��$=g�Ǵ�>d�g��|ɦc!���E'S{���ڀຣ�n�b�_G���=3�}��g������D�l�|��I�L`k}����v���!����{�2�y���g�N����a8��=f3I'��}���E��6����u�}}윟G��B>dY:��i���|�E]�tL!1��I�L`h�p?$1�ͱ��!�|^��O�z���'~d��w���N{�LW��%����ޮ�����|�Hv}f��'P�VN��'���"�ש<9@�2f�?w�O�&��C������d�0��������.>���xJ߻'�s��S�I���^t=d� c'�<IY�;��"�!��~d�Cɺc'ܤ�� u���9�& u�ɾ��B~Hx~����C�Ѿ�>��EC����XI��R*�ۮŎ3�:]�m�d����z��>@�j��E'l�	ċS��%I���I�)'����N�~氞$:�:r!��z=���������}(|�7���0��'���ɴyx�=a�>��3i&>�̞<H~5a�"ɷl�!�a�o�H��I��&=��s�s}�}�\[agNU��G;컭����;սe��<{��SMu�WS���}��6�^<І�f�[��u�}���Y��utiaJ,�@Pv�A@JMB�_i�v��+\�z�$��f�v�cyI�,���|�nK�*��:mwK������#ޏz!v�~��}�{�?�x��8���9��d9�`u��x��;�l+%N�m�~a��{���I�g(c'�Ć!�E'!�!P>a���l'��>����u�=�翲3���8;�m-qS�3>����>�GLu��C�&��79�Ԇ�;���Jϒy��0�+4]�P�dS��C猓��k�d�'�1�Nr�ߏ�w��W-��*ĭǢ�".}<0��똈�Xm:�z��l��:���2gP�sz'��	��°���i<���,�N'�IĊ{~�|�y�^oZ������U��洶�ފ��؈��C�b"���>C���C�k/�� x{O��:�z��i��z���wS��^��i�Bs��?2W�?w$YN<w��^��=�����Ú����}�1�>�}�ދ<܇�:��~5T��8�0��@�!�u�j�Bz�է�q��uY�C�=dל�Sl�y����$��߼�<�[���;���ߍg�bq���$��N;O/�	P6����i��܇�:�2�Q`xÉ�~�P��������Za����<�C�:���kV�ݖ�x�����x"}�>��Y�L��V�1�{�op%@�5/�u6�i��Xq?2��H~C��YC��Th��{��z
�CXm��T�q����?~��0��Y�������IԞ��Ԟ�a*s,�$��& c�ӗ2CI��ܝv�i��XzΡ���uf#�>s�F__�iE�wn|�-�y�L�$�;;N�i������%q&�vYL���0�S�wRg�H�o�'�:��5�Ć0�md1!���&}��{7��E�9GU��*W�����'�k�	��~Lg������&�P�O��E���8��"���p�@���ԙ��c<;�����Ѿ�+��/��u�,��?*�v).�2r)�E�'�k/sz�6[$�1k[��$����n�0�;V������S��/��'].�%�^�QV�ځ弞���uN,�t�T%�ٮ��b͡j��*I�M��׽��4�RyX��t�n�1rT��&l�Em�Я,j7���{�}����y��=Bq���C�'��N0����$���i�x�q���c'_P�}gR,����(��L����@�{����Le����z<5u��}���;o~gd�L`t=�d1g����#ʡ�O��T�a������	�E�����q7Ld��	���D}1��{���"*b!ϡL_kήv�[|�eg�4��ڕ���c��BW�����>�6d��!�'��hLf3�P�6�3���xϐ?j��?2Whx{d8ȡ��8��T���d���Y�f������Z����_�����x�'~��C�6��rĆ�wz�g�O���d�!�1���^�������I���|��ć�Xx�d�m�{d8ȡ|����ߟ����}���o~��J�H���6��l&>�:ÉĞsY'���?}��C�O��P���{�@�
�SE�|�?0�=���	�>5̆�?<Hw;��>��f𿽹�w����^�,�Շg�C6��}�H���:É�7`u���sX2C��s;��I�߷ϵ��|��϶|�p�0���K����Q�0��3g��h��b���^�I�wv+�ӓ��K�͘�o{�ۘ�>͐�w��n�+�7����{��a^�#I��=�5,?l����s<�'�u��NJ����K};�. �-��B���]I4H�R���ݭGT�vw�Պ9��0)0�;��C ͙pb�׮1/=�&�T��� �T�B����3pB�����tgT�^���Z����pq� �.��/����>�k�������զ4Q���D6};gN�&�3��st���mwv�Q�%U��:-xp�V��EN�-�x��>j`�=�p�
V��[��^^\\�����E�jW:o�n�z�Y��9W;
U�V��Fd�����SU���@�l5{w��|��qyϳ:�v�]A�g�6� �u�U�]��vo<��5�y[5�.1K>� �rr����,ҩ���J��zg����������]fA;(�l�Yȫ��z���oW��̖�c���ŧ��,��Cג��.��XÞs4���z�=���I�t`:{������Y��`���j%�^ߠ���bg�(�SBSݯk�_of⾰m�x�@�[���E��5���0<����ᮖ��v��n��7�9,0���p�^��v�󮈷ۻ���~�\)�I��3Z�����d^�F(|���Ғ�F�ߓj�����B��Q��UW��)f�
�:^\m_��wTF}|��cy�H�+�p|�Ĕ��(��y���~�Fr;�g�uBt�.��f�W	�r���:�2�Ӟ������������o7U��R��i'�͞�9�E�sÃ�ͧfT���t�8m�K��U��%Vm+����R��wk5� r�&�ȱ�na���JS� fF�C��,�ވ�{ބ�sa6;�Y�ߡڙ2����Yq�VM%q8���z�B��\�]r�zź<���w��Y=i�����ˠ��U
ĝj��]Y�*$A�e�/K˶XkXՄU�֝E�������^��Pg_{q^�� NMT�v���oN%[lR�����VU��{a=��ߒ�s���F�Qș��ynOP��6sS[@�+���xbuc�vyW
�N����!:�W�o���{�MZ��̣������ɬ0�҇y����R�4��os}��w���t2��#���TM�5�+Ʊ;�BvA���D��@�,u�n�,��8�#"��#^�C���f�yPk_���$9J��kv�2��R��q�.�%k`<G���=��5�P\|��i!�Ʋޅ�O[�kZY�������E��LP����J�KK�35�2�,{����m��Ix����]ô�M���DK[�>�wjӨMfߵ�8�V*w������MB�AN�ŉ�iڀS��P�Ïvs㮻����7�_8�7��AC��fpM nJ�gd��k���j8d��V���B��']�E�����#��G�����v��H������pyZ� ��Y���zr�w�f�����=<����Ƿ�z�<�Bު��8<i����E���-����٭�y��B�X%�j����������ɍz��N�{"�dU��WZʼ�̢�XKync�[�\��~�xT���jM�g�ά<��V}n1�n�]*�k\54i���ɧ���L�]jw�(ڸ5	T`���V�E�4۞[�.ܑ�#����B;�K�S�!�2b'���ú+�;�jA�R�RZ	�3���E���S�[�nz�>����5 й�ӵ"4��֯��;/f�����"��Uq�]Y���i�A�rsr�݈�5��W�Գ��{.rmħ�Q;�,�-���J�/%U<�{`�yG�f[��׃�ҤMt�k��U��;�H͞���6�>�W�~�=��ӝN�q���a�&�m����;��/R����<*���.M���تcG���7�ܻdy`�[�oIH9�Wq7��L��U���%&]@p��X��օm��ZT�d�l�ܯKX�
5`��&�=V��R����O���]��`���DBZ�,�X}׫�:ݖ)��e"BW�s�i�_�nӼ�X��ٵ�rx_a�KZ������^����l[��m��$5rץ�41���$Q�fEe����OS�ժ�H1��<�Gj�����4D��L\�S�K����۵1v�c��U�Ta��^j���㞱b��n����g�ju�(��S�X�o�Sz��UTk�U0U�co���#4˄Ny<K������#ތ��{~�Y�Z���K⇏�դ3�>Ū�~�Q�gV}����n�otTF��%w ���w=^�ֶVb��:xt3��.���9R����4���]�n�n�~�ۗ,�J����eTv�V�e[r��J���X��yyzڶ�g:S0��"Yx񳩕L���]r�vy��=��(1i!�.Gy)}�����nf��;�v��#t�\����DY�]0����p!gk]�Y����6����m�+6Zӡ��g6��#ɞ�or�a��:�>��=�S鞡�$�9�c@.����qoN�]|&�z{F��2�k�����a�5w ��v���3.� L։��=�@8�*��=���])ݤr�>���Af�-�i�Iz�y>N��ZUݸp��z�K���}۠s��K�������F�P麽�E>Ea�q!x�7ި�_!�|�Z��uo�W����ۊ��Z����w�������}&Ǿ�������o�&'<�`3f!^��bSْ�^�W��ͺJ�����.�g�s�*��azJ2q��\�ͺ��r�9��H�fb������b����`��ډL�.���|��^�$%�^�� V�7�����	OӯM@��5�.1�9�brr��ïk3���]�}�Gk���4��A��;�6��4��ͮ`g�C�UXZI�幘�W\��fp�q�X��z�	���и���7��*�p��c��e8�}Եq�q@���b�ؕd���fk0e����J�{q��L����c�rz�n������ʄa	����� 3={�'�}F�h�����.�B*V�JSk��}����Um�7m�][�)��z�(:�j��l��F����o8��q���X/���a���E	�2�UX�X���P���J���4���=��֞6֭��*�E�A
�׹=�~k4Tk�.�WhX���,�OWl~�.�ŋ~.��U�]G�:{�|����.�^�}�PY�@82{�6x7~Oܠ����'1�ލx��H�	�Qm=��˗���L�M7��l-��n\��eVj;��Y��֓�$ Y*�bi��y�[��׭s�;ݮG	��Z��U����w��*�f$I=ӁU�9�`r�����ny�2��%Ӻ���X$�ڮ���=�5�,�l��;|���7���Fku�{%=��-��Q��x5�:�ۊ�if7Z��q��_{�zǾ�w<�������C�������\���'�Zn5kS���C�݂
ݺ�P^�X�"]�<%2�(7��v�s�Wv�u\��v�ud��c=Y�Y�u�}+��hN���{���w���N�����h��GH/I�*�d���f:��,ڔ���B�m��氶k���-��=��/{р��M�퇫-.������X��x�\B��V	kE�}Ym���M�ۏ��*]L�K�|u\u���Mu誝
��?G��{w��؞��a_~�qƣ�C=�6��Ŕk�d!� ŧ-O�:�;Vu�b��x�z��L����q!��;Q-�λ�5�/��gR1}/����Ռ�0}�؍}����-N�
�`���z殧R-oL�[ם��SįC�]X�T{\0���|Ň�{���/6{mV�q��V_tݓ�{��;X���P���L���� a[���E�ZA8�&�\r��7���q�NZ�q���>��K��2��뱶�F�fn�jj9�R7����F��%�
�Y[pjb���oϜ����w�XDy���i��IS��[��t(k.�Q�����5�^7�wy՝}{s�X���ħ'�����L�]j�,��m	E��
m��Hr:�\�U����ꪶ���#����M6u��h������Q���-{h{���k�]���o�������e#ώ��г��;��.P��zc��+]Ǵ)����+]��r�M��Y�/�|�����ݙ�Iq���jP���3c���I��ᤌZ`ڄ�Y��%����e����3���6�+b��mմf�z��X}}�GiOkI��5ٯ�v���h���-�+e,�u�rmˡW6���$5gnA+(I[�:�9�d-��N��]�
�VvgM.C������Q��DP�厔A��P��O�M��b��찝�m���h	�/9��Y�Nce��w#솴>=�=C8��j�q�LNdp�,[��*gx�t�X�{q]��h�PyJ�(���2ָ��g~�،�Y����0*)�z�+3;�3k���O�뺲�]$�E�9�8@�/t��"]h��
澝�3�"�۹r�J\����0��@U�vQ�u�!�8f�4�r]t�w�
]W����Ft&����B�"��v�nMl�j��㫍Ip)J�ṥc@ �M��uf�S��Ge�$�%c��z�̙ZR�h�թ7R�;7+Me�(7��n�W�'%}�M,]7Z�i���M�>�V���w�΂���S-�Jʋ�4)*�0U���X�
0�Y���X�]��e�E<�U�����m��=pU�\��N�M|��|����;�Ֆ���������ɛ]���&z�$	�u㴣�0�Y��ĩ���2��ɻ���F�	���q�{��lԍZ�5R!�;԰�K�I����3��ᦎ<9�C�љ������OPW�:�i��z�힃��B��!U�@�O�љY����A�j���W�2S��S{�nr��7-�5�E�0����b,k[0�9٪⋵�6�����*�s��,� ��foh\CKwd��;\2��G�k����Gsx��,��l�=�뇯��8�%�e���kvD;��#L�}gT�Y���^�K�Tl�r ���β�u,�{�C��82�It�4Q�hu
��Aґ���ͱ7��t���妙Mm���s�ȶ��&�MPkJQuv,v�9ۥ��]�_����.w�5��fܪW���/�ߙ4;�S#�^� �|Nj#�"�;��9�=����|,S�_fa�A6^�L�9ˬv�qB^[`_�����ӵ�zl���,�p�e��G:ɝE��6�֥F��פ�ڬ���fY�Yqj�` e������}�v�Z��r������C�
�.Ы������۫�\��c��K��N`����n�8��5r�&��8;y_K�*�g.�ب��C�Fd  �N^��vN����Mkɖhn�m!F��d�=��f�Y�s/ZA��\�V��{����Y:6�ɽ�ur�멡���ƹ)C.>;Xo�[R��c3�K8&���n�
pS��h�l���v��g�������WF�
�v�-���-m��iUP��mb����Db�Dj���QKk+!TAA��PKm���c)Dkci+J�Q� �-J�K�`����X#�V�Œ��m��B�-�����
ыQ�Ъ�`�E�"([*�j6�1�"�E�PTb�,J�P�DVډQP��*��6�JbU(�
�Z���DAKJ,���U�Z1m�"[b�kT+Q��Z"1
�mFe���0UA�f4R�j��mkV4XUVV"�*��#��*�)�KaF���֪�B�5
�l�����XTZ�f8�Z�)J*�,R��DQ-�j��*�F*�TUTE"��)h���-,PD��J�DV��[�0�����Q���U��DPD�b*"T��UX1˙k**�\�6�(���k-��elUUX�EUFD��L*2"��cl���J�,A�eP*�h�U����"cjҋ�kQb�-��Y[(,F+h���R�E�R����Q���UZ�����EQc���F��}�^pN�)��̓�}շr��s����y���UҎs
ܗ�o��{+/�J�ze�jI��Kӕy��
�Y�W�3��z=��q�Mi�oj�В��"�U���S�������s�ג���Z��fh*U^vG%G�͇��^����*�W�jyq���4(=��}����E�n��������G�.xħ��W�)m]7G�άy��m��]\@�saj���i
��_���n����N���)S�u*�U��z�[n+6r�sι���qr��l�*N�3n��f�!(s�4�ׁŗnӨ�Q5����P-�`��ڈ��6Ź^�m� 5�Է�(2`�t���C��Ů[�j隽�Ǯ�t�����	>Z�Ez9�4���EV�>u+v`�ug6Eb�;�3m�U��6�5��P�q<�s�,jvmi��UO3y�Z����nFmOGd�5q��*�<���<<SYk�j� 3V��ۼ��	��\��~Oj�H�U�6�R>}�Pr�uq�~,9�-�[Jq����FCkE�ʺ{�g+��2�f�o�<EHsvx���{(����!B�h����m6��G����]����Yz�^eG�lĆQS4+۝�HQ�Ȝ��u0eܳ@El�_C�"�X:�]n`[�{ވ�=V�>�)��_F���뺹۪��u=������c�,�x\���vb��G$�oP�q���x�9��|��rS����x09dس�ۚ���v�4�i-�C�puk�*�i涔E��qҙ>���U�ں�Ec&N�ɸo*�f�3����s�`f/�I
�z�W>�{�i���\v�z֦܎ޡs.w�*^�R�&��P��U���|�'�Z��v�h7O���q�%�S+�5��9;�.�d�@]U���{:k.��-m�ܻ@N3�	�+{9.��*�}-�T�,���t����MS<�j�%��y�c�裃�8�v��t�a���襱���mL��cP(���H����<>�X�=.�*�,S�B�&̷ޜ�s�	b�r%>m���/K�;�f):��#�ד������sp���;-9k{6q)������"2s.p([��"�۞�t)��J�Sո�7ct�cM�@�ͬ��a
v`����P�|��1� mb���ѷ���m���-̙��g�j(ν{ooV�p��8�qQIα�1TQ�(^��8N�t�C�FWJ���)�+ꪪ��[֡�������jo��Ǖ�X���1�A���r��a��*fk;��.%�h؃}�O��u��Y������u~}>�2$謹f���={�*�{�ٌr�0w��ӕ����t�:��fƳ�6��a����V+[�ϯ�U�s�"��AS�b�i\io3X0e��^��G��5z�I[p�=I^�u�py^ұ� ��|�`ֳEDk�.h9���Uͺm,715/�b�ì��Tb�k]p�ҭ�v��ۻ�t"hN(b;!��h�&?wi�a.�����mt��gQ~n�$����Qz��ɾzo�^Kp�.�5��~�Kr�%���-5��,�(>���sJ/�_`]Qp����\Z�3I8Нy4���3ޕ֮t��ͫ&����/�\t�y7��<�]۴֐C���!�M�_w�NOT6�]��N�:V\[�pEL�L\<c��@ȷ��B��s�mÅ"�o�~������'�橅�c%�,
��V�+����T78��;VI�*�ka�}�M��b+^\�
���@Ɔ�E{�Z���y�-��Y�)ɴI\���� ���n��7�'j�%��*�����ϓ�����R����3SV�L'���r]zג�׵�YN�v�?X�p�U�5y���9O�S۪F�N�wڲ��B��ޖs������:�����y[��)���D�Yf)mE�*�y��K�G�@N�wf��()�&���n��?Fu�p�|\�jl۠�1c=�4K9��((o��W �K.�;]d��7�+B� %��u�o�⼈5��BvG�d��m���P0�S���qr���!.�+�J}T�XV�'m�����/n����Fj�{����]d����g���BO���P� y�}7%���lb�fu�y�ʾ[	x*�[���j9^�E�����X��:��2���Su,+}��p�O�ї�Tݷc����1[��`�q]6Dt�	���ޢ�.�@q���y9�+n���(���j�v�+����=.$2�I�𹵉X��2�~G����`��s�S�j0Y����:w�Q8*�X��'-#�h�9��wu��uEc�}�����wA�z�1�R��\{U,0����W���vl*=ҫvu�Ж�R�@T��0v�{��=9���-�{s�DDz5�7���[r�����B�U�����+�em�����*�;~|����іwһ�=}�rw���ۺ��u��%�ˉg�x��wlafi��vʶ:��s�z�O���;���i [�p}I����L��֮Yy~(ک�������U�>Ɩ\X��s����w������6�c���Y���Mz�ca�L녕gw��pk��v�w#I�V�|x5KW1�рqYz��[�u���\�z�r��V���łJ{��a�>�)��=�3��!�X���J��$���V��@���{uX���c��<&x�Q+����]��h'�z���Z(>�p��U	�7Q7<}4��ׂ
ދ�[�O�B�F�Mq��;˕nr��D�;���fݡp�"BW.z)��qa86:'0��F�{���E-]d�8��c1��'kҠv�鳎n�j8����g���+���(w"\gucN-�I�V���d�;P��i=�!�j6H� ���]�e��y���r`��H��
+e�ȯ�y^�-��I�"�t���}ͮ�m-ݸw5����޺t\t!�<w��T����9�e-+X����?��舷�[���t���kʃX��k�� �r8�B��U<��Ö�)V�n��{����A�q�6�uZʌ6�Yʈ�'~�#�=�X�ٻ99K3��^X����	\�ډq�(�^�}��hyQ�1G-��&8�2���w�eA�pa��.jU�R��c���y������$'�h�$T��F8���?>���{����l��]�#\
�X��&�q�.]�Y���u��V����>u��n���^�gn�-��0S�/����s�s
/_�E���b��*�i�ƶ��{��L�FU��X�U�|�K6hV�l�hK}��_(1��*�;��|CO�e�sP����M�Ĥ��Mڙ��2wV)lI\P�i�E��^��A�߫ܪ�Ӿ\ܮn=ަ9q����G�ePk۪s�;�.�wU�.����+��mA0^պ(.],���v�&���7��GVm͈��aډM̹�*�3�
���}-�n^���Z��)�ǝ��Iu��_esO������V!���$�����-Au�Y��t���/GEl�\p��I5|�}����CG=cV��9���t'Ԯ�K�[�T/��};��k���R���鴫m�[Q-;�E�ӸO`:��$`��/�7^!��g�:/ٞ���ӵ��(9��Jɔw�;>2�w�C�\ٖ�`���
��6]�֨^ OC�)��e�Gc=���}+�Ԍ[�ȱ�-�ỉEmwl�+�E/	����b�r�31��>��\���3�y����N�کC����Tr�k�� �7�8�Jͪ�dGq�B	X���� �H]�V�qQ�$v6߯���'��U�ʕ��^;sS�)���bW�vxd�W��
�K�	R�j\e�c�� �i�͎�ۢDӷ�#�DpyQ��1�n�9=�p�h�|�Fv��=��*�n��Ȭ@��V�W=Q��u5W��;}o��[�ݴ/:�R �Gh�̽�!Tc��Z��2<ɀ��-��S]C�2>޾n��{sy���F��<&�*�U-j,�NRT�\����г��N;8��ur�I�n����I�΃���ls����9)Z�F�Q^�+�����������ة�n�VAFjܸ�x�����_(:����4��&-Zc��`ޑ��WڜiLHOU�܆:��h��,��E��
��޺���6����O�5p��M=���̙P񷜇���բ)ґ@,3���+ɛ�n�K�$c��b��T�'lvu�>��m̾	A��wJȕ{��������F}�޴��괎uQ�,�ME�����l�^K�P����a�k�㗲W{u[���T��^�N�eZhW���O 8�q�����\ܳ��{-����+o��V�ߎ�߫<�����k��$���;��P<�,��&�wXY�4\\�7s��&�^ߌS��c1�<��N$8wE�yy����8�C5�z��5Ą���&����'~�L�;㮛I��7+e�g��b��c���(䥁��� lH;^��n�s������]t�ƫ�뵇cee��7����d޳�)� ��d�S��Ǘ]��V�t��[l�ʷ�sӴ�4��#R�jf�s��t��oF�cK�g;�U�p�Y�M�&헻��|�a�v�&�R�mݟ��:��A��W���T{�������OWѫV���qڄ��2*�;�A�l��Zj/ems�,�v�1�mu�Z��A.98/��O�-��Z�jew�b尖ga�%����w�W���C+|�)��#A�n�%���*��f�
��Q�����5�%d�y[~.�1E<]5W��T=v
�*8̥�v�S:��w^�ۻ��
���_p�}^�-l�Xg���n��V�e8��`���վ[���lq��4o� ��6�[�<���	��owk±%��j���Ir4���	����L�]j嗛0f����k�_d�������.���������nv��3e�g����\廤�V�/l ����>��Qm,�f�oy�1ػ`j�3#�}}�%�M�O?.�*��o�m�F������u>�4� �?_�xr�}s��R��$�5����9�0�F�Ӕ�u�E�SE�M�F�j�0��ʺ��c��V(U�z�2Ǳw"�7˩�=�oV�۹���<���v��.��F�9� 70b��k�]c<��������!Pf�(����n�oy
��W�J%(�۟�ވԻvjq������事~Jn{"%����՗���o"�]��H�W^䧰T����p�R��~B�$������łk!�ma�F��Y�=�)Tz�6�2'�ަ�{\3H���%���Y�9��2�{���z<����d5J�%�~V�T�y��P�v8��^��iyê��]��s��x�*1ac;�y�TF�����M�c"`ù#\����Zڐ��C�R�f�:�ʠ�|~�����kT0a8�ݻ��y##*W[]�8�t����� ����$f�K�ʈ
��5<\hy�(+�`�]���gS��
q�*�Wzf+�*5.��{`T��g��Ձ&�dz�}�ӜП�-���̮Z����Ez5�R��Ay[c
ƃڼ\��p�=ڊ;>�\Ӿ٣���x����>���������)qT�:F�I[��4~�"���XQs0�(*#�¿����,�4+������]���2�-i�t3�y��s��xУU�,S���c�t���\�Ge�x��i���HR�ۛ�[/&>W(����7�a]
F,e4x�ۖ;-0ci�f�#F�9��U�A�
&;XS@=�N�68�Z�F˧m7�6��tˈ_p�5�'������PÌS�z(v���`\f��S��F��Q����[�[,*k�<�8+*Z�&���\hL�h��Ou�*C�t�k��)�$?�J���b�l�cw�(�i�w���a�{ֻ�.��sƫ��A-GO�t֦�������z��Y�ה���,��)���qX哎�˙�y����$�mP�I��fT�;/(N,�l˫T��\K�p���r��ld%'9��0a��3qQXXcl�557��k�*m仾���M4�vim�%��p�n��g!Ď����V��Q�+B��b]�J!ۖp�LѦQ�Ӝ)�X���|��d�y��u�\Z��S�ړ��u���@��`D��'��̐
�������ֺ��A9���T�bR�:���is��o�	�6����Er���[K:ƻm��	�_Wo��ڮ\2(�	�5OmA>�u��	�k/uL�z�k����i@�j;��D6��sF5YhV`X�'*ٝ�m�sRS����aٺ�%��Y�s
��E���n��n�X&�@;�^�N	Һ�S˽�[R�������J�zJPN�n���Y���2TT�(���P�ƺ�ңn�b���xf�44hĔ��:�E�[�v-��^�G�jZ;͢u�a��;t�;�%i
��.H��nLR۾Q>�6�ۀeI�k�$u���t�%�5@Q>Jm�7��ͪ���M�0'l�d۫Y;��h]S���77�*��h�����1�'e+�X�G�6�������\�
�
�wRupY[zq�s#8FI�2�ة�SVZ7c��;�'���cj˚��g3��w�s�݈��+���3CT5�n}0��Y1G{O.�سf��oPÉ�t���Z$���;��]�ݙI�����v#�����
�wH�L㯁`�$DM�:52�`�V����nù4�<[�z��d�z4c�T�k7�f�b1�upN���c'f|�]�O�zi''p^d������mݍ�T8>S���EW:�ֶ7�5 �/A��J�����k�I쭗Q!�k���M���r���4c�G{���\��N	u��K�8�Wd�6�Ɔb�y�"s�N�4�%P��*:�J��jX�{W�}h���W�[�tn�T�.����'��"���-j��O5ab�9t
ӻ�.z�lλ���j2�� 6��f���I���Ѫ�=fE}u��:���.�5�ꬮ���o/ �҃=�rʊnd�i`k�s�j��"ԭJ��V*-h�����Ա2�ֶ�m+-�QQAT*�(��B��UEUDb��PUU��b��U�*�*��A�-��Yl
ŶU���eiX*"+D�����%���**0b��UKcKh-E�6�m�ml*Q��h�F�R�A\�e��Օ�V�m-*�hQ�jE�*��m*���,E��U+aXQTE��*ڌ�E�b*��J-kQc[lX���Ī�B�PAE�TQUeB�����*V1T+
�+h��Z��H�F,�F(��`�[��X��k@DDEUJ�Xր�UX�%l
т
,b[++*���UA+X��EYF+Q���֍�`�Q#Em,Uh�J�V�Fժ��B�"-Kf[U�Y��"�Jʖ�e�4Qb*�*�UDIhX�
�1�����iX�EF��Q�2�(��b�֪����Qb�*�%4�	5��
�9K�^��
�=V_g]�-Q�ݷe�qI1�ѩ��Է:��{G[Ve��-�pWP]�i��I�\Y�f�z3Pȟ�Dy��o���B����R�P��_(Ռj��]����-���1��=^+�w���ؙ��no�2�6�ơ*���A���sJ���4���;E.����s��u^��&������a��M%qC��:��� ��Ed֕NV��.K@O�ɻ�;��]3�5��P�딋�F��y\��%�j��N�%ٚm�י��->�R�{9.�o�P���o��;�3�����c�ݔ���[S�}At��]���?=LuG=0)�a<v�&���2oOfޥ���.�-��F1�Տ�"]��\�3mM@V�n�)�y�������m�Nׯd��P~��z�̊�a�}+���v��Wl[s'z����W��� 5�D��CTŗ�r�a��fL�Uh�,�b����3�bT?kc+�ٜ�����Aږ�lk��WVm'Q���z�amηN�ӭ_j�hoN�Ӄ�Zٹ[:�u��=_-0��"�Z�Y�
��ҫɮm�z�W}+�L�Ve�gcO���L��;#�ٝ�A^��q�fZ��O ړw���@���!mR������&���
���e_�����o+V0}��Dv�+X��y ���fÎ���oZg�ލ<K�n�qN�įF��Tk�
,�NC�.`#���y���x�y�UE'�S{���!����Z��Ƹp�>;S��5�L����|�t+�ɰH绀Xw|U�b��z놪��v��;q-� �Ogcp��%�]�j��c�Xw�C�P"/�k�\J����ӎ8k�n>}�Q���[um=�t��U}�W�.���ͩ�����b�m	~���k5����K!��H�+��4�nfR�N���ZM%;�&ҧ��5W�Y�ڪ�m1m�O��;:����6�\�;�����{�giׯh��E=%d�X���N�����l�^Hr3I�3ET�@�to:)�ng��pE-��+�"u;�v���Шk����ίL'1� mǀE�r�V뗢��x9����t]v�-��G��Y��/�b���Uupݛ!�m��!�T"�<�!�[@Cu�8Su)b�ܻ�u�<-=z���B)!�Az�3>��X�E\��L"U�L�%���p������]���Y�{��pێ{�U}�ޥg��pgvb��y�L�w�;��5|��q�wz�s�#���9R�הjKQ~�jl���̛��{{ȕv�˥��+��M*�oP�g�	o��W���Ozzd�m
�z�If*U	�A��=R�v��2*#�3Qć��a�ˬ7�L\�m�6�$�0���ܱ�cݥ�E��}��}�X��
���^��KE�w�Ԋ�(�Ȼc6��>�KX��p��"��'�#�c��\�F��%�VH���y������o#����F��Q!=��p�zq�\�]6�U-3ɤ�E��c�:�d�ו�]�Tb�z�8j�M=&�{J5^�Z���S�M�����w'����K�[����:�R&���rޡr�{] Ӵi��7u9n�B�Ю%�˖xW��OM�}4�l+�&2H�9�Y��h�B�*��ѩ���<�A��4uL��Y���*��o�^��6L���M��m��+�OW-fo�u��N�S����q2�;K�F�w���/F�Qd=e�����rʰ^Z	���W��N�H<�����M��y{��C>���)c�IT#M�G�	�����t�]�y��
ҽ]���k6��}|��B�r�w����nw6:�:�z�F�'����欑�b6b�^�M#=�k��m,�f�V���3Z�6���!�S�:�m���T事^J�PguMN�ˈ"��Uq��S��=Є#T���iT������T�������W�N�wע���-ɲ���꽲���Z��{���	�U 'N���9���s�KN@z��Pi`��ޣ��y�T7�[�s�)�oSr�=B� Ke�+�z�O�짜��9�`��I�b��c^N��a�8�Ѷor9f:ֶ�읾���[����m;�Ǫ�t�NFs��Hܭ���T�����8Y�l�p�g.�a��@�n�u�S�g��ίX�$�v{�:J�Kw�R��<��g+k�O�1k�
�Ј�3�8�fq!��:�g���i�CP���U'o�Wf�=�h'�t�Ϊ�lT���zyח�Un����g���v��=O�`dꮻ�٣9��0��@[~�[���r�U#ef}�Bi��Z�젢~����b�� 1�5q#6B��m�}�Y��.��J�9�.t���A�����I��NԲj]�f�`�ۂ�s6��y��V�ւ5}�jJ�^�~��B��J�Z���o0c�*�+�zu�{���u�<�%�Ռ��]"�ν[�����[廊�BZB��/fC"�sH�͚��<P�/i٨}X�_(1�X��z�����
�Q�D�}��%��f�:���v��BU���֒���:�,�{����I�N�����nf/n+������5>�=%���C;sZA5�Q�w�b�ӓ��ʠ�o�������}�,�vz���<�I��%]n*�F���VU��>+��r]E�$o�'

 ��D�V�_s���j��1Ol���:��;�tdqt����a�>Z1��)7j���݃ܺ�M*r3���c샞pp��6F.�T��6������9oP�.��A�����I4gU�����U='-�d�*u����	��8��9eg;��'9�]���#�cv�v.��ŗ�EL���"�V͚]�,�W�D3�c���i�_D�Vw�1c�����.�Gy�19-��*�1Ƀ=��t��v�5ڝ}r�>�W�~9�.���jtj��g+]���x�) .��OjuF�n���~���Nܷx�\�^�z�\��.��5�ȧm�q�����6��J��I�1�'�Q����-��Ji�}�<�Dv�>Z��F��b9�}�6�<�oH�J`D�^t$v�i�;U,��WT�ps�S�F�@b��7YQ����H�.���S�)s�r��uTpY^��CU��G'�"f���fc��n�1u�C�@]z_h�++l��������;}���0XV�5�h��ܤ�=�Ļ�k�ˉg���)��<��̓3rlש��O���6��R�<�����V���:�
�)nCn���ʒ���f��.���	��hO+$�b�ʵo2s�1����2���Б� c���a��V[k���Ff}�i�n�3��*Yp�C�+m5g�z��ӗR���EZVF�mn��%u�f�V)��T��ŧ�ZR��X��0���J�v��Ȏ�Unn�u����6�}�w\���>�Ҥk�K��es�nd��W:VYf�Z[��n;Q��%����o]W��-��O���;9���6�\��f�۔\����~P�,�c�F�l��v`�I����[�0��-���F�k��]��L�C�lny>���YpE-��f�N�}���ABg�q�ܷ ����O.�qƬ��-y*<b[�N��1Kj�AxgV>�<�n�͎�m[�ږ��S���/��!py:���R�^ي}^�ųnВL�;���[�5ħ.�Z>�A�g�׸���%�E�3j��x)	�GO{�C�7ʸQ8��ڎ�y�2*9�5ć� ��]s�_�y�.}ٺf��w�V��3���ѭ�����ذ1������gݛ�s��/l��Aڗ�1ڿR�iTd�{���ރx�J�J��\8i�֚��	�u�6���G74��Y^nU<g�2������hI>�W��ϫ4�X�s�C���3)b�g0�l�e1�5���xC<2^M�Ue��2�m��t���P��Oh�O�x�]�7�Q`��v6oiB�K3�����q�-���� ;�:�VmD����o13Q��b�k�M�@`dH����׫eA�i����J�zIF��:�f��`e��D�[ڄݜ�lg�{η���fuT9z7�Nb��=՟I]ʍ��$e�T��F�磶*��0�Sԩ�r�+ˉ~�� ƺ�/�A͡R�oɻɷ���W��,����,�\mKG��,s���1��n��1�9�0����Ѕ���)"��{��Jh���+�8�Lj7�E�(㜻��`�E���,J^nq�q�1�Po�>��wƚF�Q���)��J���������1)6#e�q�O:�=ʣ�x�R�Eў��b1S^�R��Kq�vQ���uC��3r�q�m�Ĥ�
�BUκ�9�(����Y��ֆ�\x��#z�ǤN��	|��Zc�c�����3S�~��)��$x�7��`�;[�V��-{ӭ!4��s�x�s�/Թ�˘X3��j���AN�o�\̄+�ɓ%�q�(}�$��7ٹ�%��G�O*�w��W��w�M�Ph�l�]Kk��R�=��e��Y��,8�Z��%S\+;�����/KδM����&#�}ċΥk�NvR�r���";�e<�m!��緗9S�K�&�j��$� �V"��o����%��|:�nO�;i[�g�¹�c;61�U�����N�O"%`tX򢏽��V]�XD�Y���P�@�<�:\������)c(��^�E���u��]�1/�)�Acmt�Z^�n��;��5�h�
#����F�f�����py���Q`��r���nA���9$�Swֈ�"�y���|��P/u��6�.����t7�P�<�crcͺ]�2?�N�j�Եq�x���s5���O�Ltxjz�Ui�0y�J�fƯD׃�+.��kX�X���`K�Q�ĩ@3^P��U��禩1��\�2��m�X�8]��\����#^ }K>�k�C�%�b���]\ߥ��n1�k�dڧh��N��s
1�Ě3W���VM��g �*glߴ=F/�Z�K����|�2n1����%n5����vuyNؐB��β�Iv�14�[�Z� =5�/�=ǧ7��>J�������8VߩΑT|v��54���Yo��7�2�?�!�7�}:��VeGe��dwm'"B�e��v�!�J5���n���7}G�w���}W85�CCh�T,e���
�/��&��u�n�7�� �ls���ǎQy�:�L\n�2�L����77>i���굃z��޳�dU֗Q��ѥ}�m��,�X66��#�}ϓ��o5�gW��6.!�]6�!�y�9S��_S5�4
�U�y,f*�U�wu5ك�Z�7�͊�}J^y�X'�+b����y�b�`��]J/�1�X2�����j�ˋ;PS�����M�iS�TO����hQ�̥`Ի.�6ZX�`��?{�"�7����a��1�n]�7���fB7&)����]�Y��*��PD��L�|��o�;�GBj%���A3�_g���j�s����w��Wj=I4��������[;���6� �h޷�8m������0,s6<yX9���+���`�e[�e�}}Ҹr��C�)�rߨ�A҅��2rMX�F�z��&i&���/923�����PJ�M}�����"������aE�MNܷ��O=0$Z7���y�N��뭣���|�'�)0D�2_�:�l(p�(t�Fp(j���m���G_�C
�Mڰ�,�{��6�E'�(�B�2��|��J}�H1�f�yT�:�U���X�Pܚv��1h�W'*6��'��5����"Uxfb�.��U,O�애�J��E�5fL���y�q��w�*Z�y�������N�a̶	�u��}ڳ��@mf�r�:�e��&'��*\!�DX�M^g>��������O+��iv���ti�F[f�b���C᤼V��=]rX�bçfؘ�h��r|9���I}R�1�̄�����ʸ��.�����0��bj�e�9�%�h������s����{o<{nn����d��F�<�Q�.���r���eS*`�|�4�kL}����� �Xi]G�YO_4�5_|��È=�oCҋmκ+��v�p=�4n����E�.�W�[U݈�un�>��U����ϑ7,��;J%uof	(ʳ�D��v֩q���z��7�-����U�ʣ7q���:�|�ua�P���mY�Wo�JWl���eq&�]Jy��1���0��;7�-ej�5u�i��y��y�eWn�94e�|5F��e��[�^T�}5��PN�V�)�N[��`��y�w�XU��=��C����A�]��R@�.WӉ"�Ҷ-�`�ۇyor�m�VĔ�\pY}t�ǌp�w��Ŷu!��§�ֺ#{��+6�f]IW�d:J�\f�;���̬J^���ќ�hR�7f�ۮ"�a���:��M���U���7'R��s���J���u�g��j�̸�*=>�d��c�{p(��wƶU��n*w�RӘ��Q�<�Xǈ�l�9M�����ɝ�
�܊�B���M7�b�f�%R��>y��ζ�:�u��k�ה����F��S	lj�7]�ƶ�t�L�6o.l���cCh�2iH]G� 7ŋ&��Y���eGmA7K���&��ə1�u���j|�=��H����^��r��'	�^�m"�}�h�c�űњE��`�0侏E�9>���\�	T䝇&仴2�P7������3e<�${J�+���Oӛg�K��*ڢzpԖ͝\��e��b̀:����ܣ}D�����κ��'D���m��w3�,V���Po�q=�zC6�C�1.��V����w���;��,��EB��)��+>Ә�yP.�eu���Y����`'�8�n����cm�8�׼���rav�f0�hN�wH�thy�x�+U���'u2�+�7)�nM��ƝQ���́�Y8�ƕ�p��B�ұŗ�����ω�F��� ��r�wS�L]�~w;��Q�	3M�6�ִ��'n]�r���{��J���ɾ�v�꺸[M���758��
��m3�fc\���}�C���y����R�|�8�9�=��8��c�Zvl{�}���V�+TD�j�,��ϡ"pI���.t3�s���5���;%Bl�z��B���[ί�k��)rZ�\'.CzH�C��C�Ld��D����Ye�ˏ�,��߷��R�5*�j|�h����E�Ģ+",ʢ�1*#��
��0Ɗ�b��Zث-*"�J���m+��h��*�,E*QPZ�Tr�E�X�(�Ub�Ȳ�W3AH�ˆ.fLQ���嫍*X0DUA-(��4��A�n5�!Kj�imEJ�J�V�)b2ثAURҵ��n&
(��Tb�e��J��#Pm���ʕTEQT�KeX���5ke�aKb6�cZ4A�[*[(�%-��*1jQP��V�b)R�R�R�J�m*�KB����G-bel*�+iJ�X
ZPbĭQ�����kj��jUE�QX��)AUE���QA��Q������E5w���s��؝G���S�Q�g_j�X�����d�S��eFrS�.�gޔ�6��*wF���l�>E��[��}��ބ�;N!��D�t�ĳ:2n<Q��K��R������P��V=)�F��҆��8�z���s��;Y ��'�΍j�̻Ձ��b�-<tA"}�t�����n��8�4�V��<�z<9�ݱ��v�"�f|�q��=���َ��������_i2�mu��g,V;l8D�sl��:��V�/N���y`	x��*�������u�:�.�ZKI��uTMF:r+�\������MS�y�ȑT;]���C���j|#1=�y�G7ؙb:D���&��QY�$`��|T���bu,K��*$��7\'^N�]5JwI]2�!��@��~�}��U`x�e��ޱ��Ҭ�0zkB��}��Ågc�nĦ�A�f%;�u*x�̺9o��4��c���]:��i�7���U]�J3ǣ��������B&.Qް��Ʌ'�=��L�r�����V8X��6�}('��z�
vT�鄢w��i�(���>�Gr�R7vGӫ&�W�ͽ^�TC×�.���0ڰ�3�ᚶ��u�����]{F�c���g��9sڱ*X�YY,7U}��t����e�3xr�f����2Bp�tak�X2�d;g������F]a�2;��jKf�Ӛ�o���wmM��t 6��br��2ʙt.IJ��:-���欸������Dn�p���T�ë8��7b�XL,{��w�Ѱ���:�C��[�O��7�ZL�:^��Փ~�8��;-q�k�0ځ�������)L��ɥ���@���������?a����)�T�a�
u���L�Q�#,U��8�Gچ�^��z��$���v0O�����/#*���x	�)��c�U�	�u=\vf�Tg����Ood��'�Z�X�����}	����V�]��h�ձ�j�i.[�2�\p.X�T9z7�s]�{�E���۴�˖�I�1�7�7�r/�Ε�v�ᢧ"\�5c}���Щs�	�ɸzah�Ug],��\f�ȕ;wQڳ2�{�9���KU������z����0��5RF��~�禣ɪs���RD�ůW��s��" ������nڸ���n ;�cB�;�N�s��{�mW5�y�6���r�Om�{�អ�����p3�=��6*��4�6��P�"�_a�C�i�|���i�����y�c��y�بnu;�͛\�����:u��x�˳6���:D�79t.M_��.�t��|�����ɤoSZ�v=�CmH��� Ɠfw��kl+�����H�DO:�=ʣ:�v%$��h�|��<��o�=Y�WՃ`nw5�HLt�l1�J{�I��b��gκ�9�(���;�*���q��rGL7\ic۴���9���F���O�_���fj|��֥,dd�<�VGTK}q7�V�K@$���u�vީԺ�:֬1�^v�s�>��M��.��h\̄*�2�a��t�I��嚟6X�z�vH�^���!v�_�=��H���[�1:�<�`��ѺC*�+:��=w��xF���Gv y���u�Q���`3H=��U���s:\H���6����N���i�_.�G5v��%sM����0EzX�oÃ�4F��:5P"1�Wp2�=�{mOS/��NV��VG]I��
a��
Ӆ�0��u�M�]˃ȓ�Ze�Ǖ��k�~�32�*fFG's4���O����[�K��u��Lu�LoҔ�KZ�OXz�ں�`K�Q��\�"Y�(I��<!\禩?�RK���NX�s馽�M�t��ݪCy,]��_=�u*Ru���A��rԚE^��n+���0��C�9�{+���%���2�SA���B�9n�"t�ֻ7�2�=��P�s9p��.V�����E�a�o��TyKʔ�;�%k7�VR���p.�
���R����pNM�Ȏ(��6����a��x1llB�H\-us�`3�ٍ��k�u�6�r	f�P[�>�XxWNoظV�b1�ĭg=.n_[瑓��cWh�1V��=!�{����Zt��}�ng����[�hl��/�o4Vx�i�=Y ��)�7�����Nƣ5R��hC���`��}�_#*1��O<����0��S>(�unvt�ݴ��0�:�!�Azz�6�v\�ҩO�wQ��S5�4����C�}ٚ�;ԮM�f������B}J[�r^ȹ�� S9��j)�s"os/^,���h(�y�=���t��L>��x�EZ}pS�>#@�p&R�RAގw����oޫL;[��2�����=.�X!�����ゎ�7�X��Gs�U�йO��9[��`��Vp\�(MD����	�m��=C8X[�{jǭ$7Ua�KI��8�<Ί����è�IV��u����Z�~�ߣ�3c���ɪ����fv�4�v5��}�k��J���f�������h\<��"�x8���
�����8H7��W{V���%ڮg�V6��[˺V�o����	��f�RXՒkn���{V�����ik))E�tʷeĕ���v�q[�n�W˔�S���t�Xc�Q��؆��U�V9�5�V*φO0��]�:��+-)V�e�4n��rT�WX����Q�{�����i�`�Kc��S��_Ʃ�sv��/ϩ)�N\�x��nW�Ὢ �M�U,�TR]�d�펱
(�:&_p������Wcj�B�����sȺ�9�ݗ��1�W�?'A����D���\h"�k|XĬ�$1��m��jlO�(ʫ|<�$"c&�<f���p]Tif�&�Ui�i����<g��u���Kvs�E��څ0��c/��������8>��=��̎w�����,UC�βowdv�)�%�yh���#��9L�َ�����J��*x����oX/x��r�Ѧa����KӺ%��^X�Ӗo��b�P�
ڎ��]%�SƖ�#�Z*3]D�b�#���*��puҚ/E�αc��U�!|If��n�I^�����t�#���w��z�XʞT�R�����8QBӲH�/�yǏ]F�J�'f�}���Hบ�k�vpX��[�8t[�n׏�A�\=%۠�P{�]�#X&5�o�XO�����D���ҁ^lΏ�˔�M	�Hl��ǰm,�jw
������_v�M�,>�
b9���?=��c���Z�ʙ7�ow٬�I�ӓ5�u�"U���UGJ��8Ҩ��zU�CO��q�����ےa���k�0��8�W���j1��q%�����(8O�c���Lg�巚��es):���]�D'��3pF��&`1q}�t�'0F�Y��g۔�ޭzq�����y��i��0V����7'ܯ������H�3	3����]Q[�>/�[]B�k���r��䫦IV�O���Lķ~4=>j��X<r�]�G��z]GZ�q�"e��V����b2�2s-Rf����jED({���|wDİ����k��t�]`]3ϛ�q8���W�������V~Ӌ�N>2�W5E�B%\�4;|�K�a�]Ћ��/WW�z��Vha��fƇm����a�ծ�머[���3����O�v�^��yϵ졐��O"f�C.���Mz����N��pb�yP��	�!L�wVk�[�{Й��#��v��'�<��SOod�5ZI��zIF����*������{hī����>�#�1�~�>U��tU��]�z�,�'2T��qR���F�8(5|U���ũyH�ن��'���o9+[7���%�k�9�WA�VE�\-0u�K5˺�h������O,�2��	�\��$�}���)Z&�xM���m�s��r�*���;�棉S�&K�O�.k���Cct���Ǥ��pEN�廰�㑄k�o
��O�h���
n!
�����=0�l�+���n��<�D���w.���ꡩ�S����k�UD�Z��(�����n��S�]���z;{8_^LR�@
���Ş�m�ss���
�|j�s࡯w�+��A�aL���=�7����h��l��+�&z1�o�����xR(wdhhu|���ɞ�gUz�r����f�J��s��_��9I��J�c���}aY�~ՍU�x}n�����*1=�2b�y2�LT�Mq�;E�_0��69�9�k�b�({E��bߡz�^��`�L^���V�t&m�`�ty�kk�LY�b`_��R�lW��"��]>f��ڗ�d�w�OȈӺ�R��N��	;�,h6FK�?���<�f����u��y�MwtjP�TQ�C�Y@��C̍b.�����gր|��e��`J�����q�.��&��ә	x�\Tr�&FUE�^�ȭ�ɭ?q�c� @w��m^m���۠+����A���*�!m�����5�/�XS����y�2����\���ף��ޮ�;sJ�����z�c|��a���ԯ�\-rF�-·:�u,�>�[���j�(_G#Z�u��"	`C����׬�Ŏ����#��[A̤�fL�~��^��*��DR�ز����u~uf����t����ú������/�,�T�Mv��$Bp�T�r3(��ddrw3O���r9�Ih����Wm4f'q�՛琾�q� .���WN�ϒ3�����BL��xB�ղH��@�I��Ͳ�5)5�)��e��׎%����\�=U�B����y�9�6���]u)¥em&\�X�VDf�2r�]t���&�g���;B��1�}��1~�V���7/�Wp����nE<��'r��(��(����b�v�=����i���d�@{e[�+��%�Cb2YT���΃���{��{��X�!ME��#���f�h��p;��F�5�0�s�cw`���vHS-q�^E�W�r��9��&8Rg����e�)畳�u��2s�qF�֖�b�h~�jk��@�F&)>�/!�[6�NH�Hw��S+��ُ�H͐�ex�ڜI[�Ja�£�{���J&5&¥a4Z�*��f�z���ڍ���%c�%�N�b�T�+��XJ�����_X�
�9G&%����<�Ti���G[q��έ�'e4`7������:�����SMw]ݜ3FꟐ�i�}/��ob��Nά1tM��TA���h��ଧ�u�G��ߧ2`]00.�|IF͑���6�t���9�*�����A��>8�(<{]`���f#ri��;Y
S:�w�U�o�v�:pu�6�1�t�0P��XS\"����د�Վ-o�������|�Hǻ��Jmΐ۾��.�a���n(�ؠS�
�f�FJ�qP<�D]L�m�����jM�)kU�'%��rė*��.i��sh�tx�%#>�|j�{�h� rտ�*�;�Wt���툡���kUH�.�o�^\ C�'�Ib/��S�aE�j��d��hZ�`M~��D��[Gُ��?i�zA���F�i�2��C�̗펱P�Eu��{qb1I^J<r��XʛpW7�dyhʇ^�e�Bb�-�l�LD�`��w��܉�ֽc�Y+{�m#Z��k��<�r�ܺR�6��J.r4<dҮ�D�bK��ڻ����@���ɿD��Pn���Dx�:eެ��1��j�j�3գ=>-��H윙y��T��q�y�X:�c��שX�F%�b�s#��s���h���tDm�)�
�p�ە�W#���pCX�f��c0��w����Cu�gsE���y��C�ET�]`�ʸwˆ4��V��{�����	y��-���L�.���ѹǈ�D�ޮ�@~�Oj��$UP�)���	��Z������z����u}ٱ˖$���sD��u�J�DԹ܅%���p���y����؍%��=${�ga����W(C9?�?'�w�/ةȮ.R���ヮ��&���r%#؁�y����C�}���g`*���SdRG�=����
H��-
O�Kr#��b��v���JNC�� :�1gT�e���Txhaߒ�܍<�S/9$&vrT���w��1s���,v�j+� �֣0z����}e��ڥ���9������b�'�k:���[�ӓ"p��	�1r�>��arjOX6�xn�g۽��˫��n�&�E�U��eWM^����uȂ�ۜ�bffg�0�������;������t�n��z����e4^��!�[��\��^WDƺII���W|��\ۡx�1�']hr�+�U)Ş� �QꇼO�C;�bZ����ߩ�rfkB�ͼ�y]Qӿ���"�F*gegΥ�3����w<#>cp�=��/�x�U�dӎʒ���w%ݛ(���j�Ls1��M�+�i>�Mm�K:���jt�ն�h0���Y0��)rE��.�A�il)ӫo6���n��w\k2��B��OY	��JQ�r�IVj/�ђif��{��N�I΀�ܮ��o�;�F�m�ݨ�u&�y�0#�$]�<ďJ�9<<�7��
ʮ�E!�`*f�c0�,�F;�G�廂
��oM'h�퇏`��po>����E�"��O]i
]۶v���(]�1lx�1B(*�1����Pw[�����n\y�srԒ��<�m'�~�{Ք�U���JN�}���=��T��%՛�[5��|�� 濲��m1�lE�M�ˤ5s��V�E�zd:�T׏&��rL���Aal�	�Z�fn[�`::�Y�a��е��v(��Q�yh�[]�^�5a$9ueij�|�W|,���%2���:I��g_p�æ�*\AxșPl�U��_B�:Z1@�3sHD1P6Y0\hsR]]�mv69h�M�R�vI@Ix�mpB�Χ³ug/��γ�4�q�̕*h�Cb|�KtQu|��8��Ӷ\�5ޚ�%B�Am�q��+Dw
%Spt��u��e����\󰒖I��ZcQ$�֥�Q���o7�!3x�ӑ�F�[qx�繀�biZ {���;�2kU�8����$���gV��@u�L�3U��*	ܻ�{9�x:���kh��]/,��X�笩ķK����C�m�N�_ujV�����>���#��/��]�!��&Vq���\�H��.���^�T��Y�����o|����´6�ۈuih ��c�7U�1]����!�x�6x�58P�j$VJE��Y��.kDAz0��>���@ݣ9���k5�s>r�+*:1$6@����=ɝ|�$F�ݒb7�h���z*��=Se��{}�ݫ���[��VvY�9�\~�B�q�w�_s>��h�x���ui�kMw.�.��V�����F�.��k�]����5��7�B4ҹ�[ق�e��]�涪wݹ�s�s���u�Ób�U8N�<�mʺr��c7���Lw�p���Soa:4���v��mTQr�\�ڙ�_m��o+�،���WBh��n�t88r�=�/�
S�l�b�J�ӓ�T*
.���u(����<�}�Q��%�9����,wv�:Բ��SF+��V/��󴷞�}r�;<�F�PU������]�K�����ur[�pM�`�K�!�/Q�ףSz�ʌ��}�)�]$����,W3�9��'���pdDr�5)�-T�͢b�8�5pً5Y�yǊ�rٸ�ɩ�wçn��S����FΐY\h�Y
�v�Տ�M]v�����$�}.py�N�X�fv�wH�(|)U+UV(�,f�b����Ԣ)EPej��R�֊)���A�mF�EDm["PZX������*VU�X���kUX��Dq�eZZ"��#QR,U+S̸���#"����X�ETm+PDTb����2��T�Y�E%"�KE��*Xւ���h��9j
�(孵�F��J*),U*PTUURѴDiiiU.�QPE�b����bF"��S�kaR�Kj" �q�%pLXR؊�)U�TTr�bU���A[eQ�*�KZ�(�E�KiR�#Z��_�<������w�:�ON�:�N��A3Zq2�(,U���;�}ί�9��vRw��e�ͷb�H��󦎹Z�����{;�H�_�1�FJ;��܅��5�Y���}2h��+�d�Vt�b�e[�M<��r��z,4%j�B�ލm�W�orG:���?n�_j�j�� �ٮ7p��S��L�|a�q2���>�{UO�!es<:LY�G�V��D1X�2�:��bޡ{/�x8��*��4��ND5ZI�:IG��1�*6H$
��L%[{U�v���sX��P��P�Y��>϶�/�S�{����Hɷw32`N�&њ�gIqF2��Q��^��LJ� �]j!<�߭��x�5��;�%�t֬��uv�q,h߆��ҥ>yq[f�szD�Z��7�ܼw�}��;����:{7���u�q&�Mχ�%.nq�q݈��wƟӹ�[`W ;V�9��ڝ/y����))U1�#%�%y$�F<	���9O
J�����g��$^����K�4�K\S�Xv���{mNG���,	tP�guT��Z^��y����tp<$��k
�#v@��lsk�rg�\�Z�y�=Ӻi��h���ds|md�	�Qw�ﷺ�s�[P��5h����A;l��=|�SEYc.멍t�XR�U�%�%5r7�q�AP���I�6�:������j�p�c���Ӡ[�o�[��~��7j�/+O�X�F�j|�zԥ���+����U����iK����w�v��:׾d	�S���`a�L]a�\ْ$���DkO^���k�WVgz�u� ��h����ձiϘW�$�1��C	KOz�*�W���u���>��ׯ9	Ձו���2X8��n�j$�X.�Z�έ:���3�r�U8̂��X�8�uֺa�Q���@�U����ғ��ζn���g��
r����5��\[y�Z�XF�@����#	�e�Ҳ:��Vjx{~)�ٸ:\�B=�I�zu,]f�h85hv���l�ez�%`�K&r	��s���d��@'g��._Lڢ2��.xWzwr��RT�Y�E+�kN׍~CX�J"�Qrj!3:ٹ��}[$���]iף'7��v�ZH��EJ�pwdQs�n�1��jHX#d��Z�HR�W.��0W�Υ(����Z)`�}CRc{��+�W��QZ^�	�����N��%k6:��U᝽y����&��s�F��ܻW֕./�XS.��1]��M���I�r�f��*�v���Χg��L�/GT���)�����Y�Ek��~7���S���vf�Cw]Y}��V�ż�\�\(�;Gwi��9���v�����>�k���W	r�_��U��+%oK�2�̵{Nd�
bg�Z��s��hݷ}ia�����dԽ�؅5�i�Gl;�*W�;�(C�B�R��c��:MK�jOd��S����6`�d�P����+F�y�])�Ad<� B*n}��r�'j���oM�M��,TF'W7����B��R�Z�y�;!\.@�v�v�u���T��t}����D��z�JiM�k���$�9��B��'����U�m�]��{<�K��|�-Jl
���fyX0�U^� ��Y���%TPy��X'�{ү����g�	�!~��`q���&
_N��+i!�G�
�/��A3�8���Od�����-j�\;��#�*�Rf�Śb�%�f�o=�G��3��#��e:?{ET��&7ɷ.���n�&jq�-
rFܕ.��H�4�T9B��;�jJG7*����/7�F��RTS�ð�N+�G�B��m�L�f�I�؜6e%����h�l/��P��t5,��m�z��w�ʽ:�<yԺ��yK�Z$��u�Ǳ�m�/6m䴖�����^V��c �v;�ն��e���UZ��YӪ���s\p.�CC-����%�P����29�dg���ݼq��&2�_
VG:��Z8����L�:��:rԨV v�F���7�ë/�ɇ^[TS��Ȁ����{c�F�JA_�Lr��� S{�AD����
�v�
��lyZ�2���:�bl�O��FF�o�5g�M��N���<"\Fr��ͭƑt:���c �o
��������U'��
-�dE�ݾ�m�?o���.8F�,����j���Mk�2e�(��Ɇ���� �:��s=���Irޮ::\"y�d�te��βq���ꭋ���W��'�\Xlm���y�s��{�:��`0���.��9R�5.ww��:���u��N�Nl`o.�6��Z���0xxĭ���0X�>��z��X��X��T�_u\
�4�OwJGoPY �P_�<-y!\3���S�Dj���0$�"�u)zz��<�uk�fb�������
�@L�����l稡�2���tmtxha�wJ�>�WX��oV��͠.]�J/D)UmGL-���{���]:�sV:�0ѣ�J���oe`
l8s䅣����mr��`CM#ca×92L�*Ƶ��K��\S1�E���[H���S�%v`c�8$ݶ�е�C8��m�hd���m޻�)��F��Q�v�+_SƳ��'���T!!�U�n)�d����֎;Ǣ��;����ڡ�[��z\4o�Z�B���A���m{�Y�7�1����n�}:�gi�\�Qu�^��h{��W�f�rxX0�\�́�!d����݈���M-��(�]%�=Bf�7�6]i�5�R�����Lr����Y��Lkm޽������c��=���[_n��`�WMY:���U�L扖}�P$�x�D�0a�Up�$��Zܸx��B�Jg�km�?����y��,���QǨ�f$����G5�n��繛���
%�b�RjΈ�.Y
����1U���]g����'Չ���r�<wMg%��/�ZffEL������_��j��!eO_�<:mAC0�ʇ��iS�Bjɫq�����h8ںsqĽ���dO�+w2���;�Nf�d���@R��b�S���pC�饵�i\��W��⽋G:�b�9�}�LT��[OA�n����|e�	�ª�&�Y�*�#��*rn(�P����`Q'Ҵ@:�P�c\��|�%OB6�n9�����b�������*����J�Ntfgׇ�a&[\�����ݎ��ɐK�ǵ�����.<âZ\{�T{izX�K��h从3��#�3~m�}a'F��+�0^Ws�!9o�f$����z��lJ����D�9_.P��K�(�/�����J�w"Z|T~{�d
�x��Ҁ��*Y���*w4lY��!����U/z��U�m)r���ӟG^I3�c;n-8o"�����-w�2d[\Su��vg�k�^�eIp!�4�������6�O:�=ʣ�qTn[�9����s!l�v����W�^�ܿ,1SV�0pj@sҘ�g��皓�+�
bU@u
/~�y�^֮ʗ�e>�z22=��|2.˚-U��D42���x��0�:��㩙�V�ܭ��WUfm�Z���1�Uݺ���2�R����&�8����b�mA�<��ޗ�MF$\}Yux'�N��+�p"{`8��fj,[�a_��;�Ʋ�!��ӑ�O˞�V��V����F��G��&Q��Ə0�"�X�k
��Yv�i���=�7�S���8�&_�1r�bna�B��1�V[�p��(�ߕζlR,��`K�A9ǚ��*Z����l��P�2��0������:�&j{�L3�T��>�ة�����g��_^
-5��~��ݲf��� �"��:{��m���h��T=P��q׺��U�^M�������շn�;q<AY'�)��G�G7����_e��|��Ļ�}z2��W,�f�[Ae�,��S�t�Z��ˍ򚞳,�W|Ӯ�&{�c#+5BT��~4aؿI��U^�ffW�Vt�\�
�bs�T�<5=S>��^�gLs�����C�j^hY����F/hq(�C����>��& ��G^`{ZęC��$��$�~2����[��P�[�Eek�ʽ���a`(U��\�e޵%�;���Ү��=�\Jct��F4
�}FN_�Wp7�u�|���O��ˮ'Q�pS�{,]i��{Սu]Z/�����qs�ƻ����ǈ{9��*�
��򦉞ʄ���O�ʋ���<�q��I=�0]���b��h,�UW/�bմ�#�;�܆b���7 ~��\�qJ�9���h��~L�����1��:Q7!j�����t��Lm�鹉3z��*լq9�|�.j,��[3W����
�_U��2�7|�O���ppԝ��FudH��k�\�.T&�pV�$D<^���-�_J���<���%a�z�水�7���Q`�GJ��k��O>�;C�F���2��0�L���>���(���X2���]}P�7lw��v-�����a��1.�H��U��XA쬂����[���5x�53^�FͰ_Pc{3f��y[WKk2�]*��$c90��C-���ʶV��>ѺS����y��żw��x��i5��z�:�^���>o�$;o"��]&���H���&<���zh���M�d�4|��ϖ�X����G=LD�Tݷ�w?N~�Fv\�l-���Rg`�LE�qE�̀�zv�!P-���#e����:]j���\��{�����2^�c$n�J�H�F#b'F:�Ι�z�L����=�(��6I�ٴ�|��ڿ�֘E�Jm���)��&�bp�2��X���{݀]���$Em߷��;Z��<c/��\p��EYx/L5���K#�L|4Z�~/�|۾�J�ӲQ���Dz�U�)fƇm���=KF	K9ߎ�Ys�MK��o��D[���fm=\B��/�=[(V g��p�������"���s�ǇlGVj��
��_�c[���gL���c�G���5�+����(j��P`�O��i'W��A��b�ι0����|+5��Ky,�2���7���c�N�_�ܬk�#���8�ȱ,;�u�'�6�J����Ǿ�j�4��]Bj#��-���5.ww�p׵����	n/��U(�܍��2
�]���θj�7j�h[ �A���8�
D)��J�z��M3����3��;�jK���^\%%� �R�P��뽛��x���p���@��XE
�"��\�0-���+���w�OJy�7�7�u�d1�߂�Ο��C�1�������}X�C"��w^w��L(h�ѽ`*��v%6�t_I�
)�<��Q�+�Dx�����`�<b��^��a�H� e��2��%�;u���7�S�a�-"���@�N��i��{��қCYᡂ�;���ӻ�vZ(7��e
���-3�/���t��N5稃�Z�@��葵��I�T�VcaŁ!*4{q-V��TvnY�W0�s}�P���ɛ#ht�rbX�&%.���=�5`}���a|�/���l�A��}n��k��8��xXO��"�v�="��*N��dl��+r�+Q叽�����������u`h������C���D�9P��Ȍ�]Y]�9V����t�ơ�_vٍ��W�ui�CS=�e�ʁ&0<�D�t\�Ќҹ�y���cYA
�c��§��X��A(�S�7[��|�>���]J�K��Y�}�m�<��P)A��׻�	��Z��)o��3�T@�n�g!�V����K�M���z/�Zg��mn����К�љ�i]���t.K"F{Z˿�w�ҿxG��_�-��)ws[����Ƒהڪ9���䶘��������{�j����ؾE���1� �����:�y��}��׼�ҵP�QhDab��[��wP�r�j�Y��Ԓ�T��'U��L�A�[��2tYb���T���<aӡAC$�-v"Fm�8�/5�n��D���ML}��U5tD���z�=1ᦎV��J=��R����������p��p�2�f��`e�(�zadp+G�Eӛ�ٴ���U�crwٰ:]���7�L���i���)MU���\����O�h�}���P�2�sëI�g!��t�S⸢�ܮR���ѳ��#�C��e��|R��|7��x��xB�`�X4�|��W��JG��'Qp�ܽ�T�ME�Ncg<�-1}�2K&�ufe��3	/of�"k�>���K�02㻩ɸ�4����!,x�������&z1�Ow��Sȯ���D�l�s��r�-I`*�[��*q3��@�����ܮ�ԝ`�1*]�-��~���J��t�/^�>=ԴvT�j�va�}vV�MQ��Rd�z�
q`(Z#r�bi�9�� 
�8,;�(A�;� N�*�b��I�g~�-_��V 9��~�����`.P��t�C��y�U�$S���V��v��_uf/�)��ÈWu����v�N�)���_5�>�%Ǳ�vlhr��٪�Z�2H�%��f�b�����&�5�c��5�`DN�4s���-��o:>��.�V��7S�d��=��+�YT(�c3� �{`�9���[sL\\���e+�V�5�r<��R�P^V�7{Y�)��}��+5ם�Huwn��F����n�� T6qd�M�F�6�rhR�7)gN���k(0pq&.�wū�f�*�nm%�$1�\����2�^lyk �J5�kW^�2:W������� ��(�ͧ�.�n�t���Cݨ���Z]��>5�Y��E�V�v�ꛤ�K t⋧�Q{��h�p����PBY�Y�:�\����	i��B�L�)-0ֳ0���q"����/������`�}8��C� ѭ��Ź�#7��Ǫ�Zt1r5o|h�,Dz��}-YX�yn����;�)���*Ӏʽ�� �f���J;p�f���pT�gc��c_K�0*�h�������p��Kz�^�t)������ޮ���% 0Z��Yt{��lrh:ͼOx��t�0dC��᪛0��H�ۭ��[Ǌ�1��)K-��곊�J�e������κ]��)t��Gwy[EV1E�s1R�h���.�hH3;�$-�f
���wo�W��ؗI>��.��c�w\���:T͘��3�W�]�Ү`��m��J�%-��`gY�˩� ����T�>gB�Aq�%Fw�.���gw�:t�vB��1�3O�V3;�]f*�܁F�:3y�d�Ӧl���n�p�R셑�dhI�����9�7��:��Ū��SWx+4W;h!Y�1X�T�TpeD�PAcE�ELV�{���d����pG�n��� ?L����z%��bB��uvd���t�f�rﷷ�{�D�mǽ��_C#�z�n w��Wt}��9���h��P�l�F�Htǫ�1X�O��Z����suV���뷆���c���3�f��w���9ۭ��3"�X!ku����5+�r�g z���N�I�醃��v;�y�����uO�J̦b}yY��k����L��wL�G}��n�N�j%��ʸ��<�HQ�1@Y���+]�R�sJ���t�p�s����;O���l}:�P��g'��d.�����╮q��藎�cw���"�y�M��,��86�W}f��+��8����'!y(9�vm�������[�U��M����^����F�򶴞���h��U�N�\�V�����>J��D��DJ44_jr�X�n�����*����+�-�C�d����`Vm�z��z��k3+r=}q��!��@r���΁��P9������o�9�Q�����.�Sۂ`��X�TV�R����Ec����i481A�h��jRҶj����4:C*i�ȣt�K��kb�*�*l˦�EEDR�Ah�h��2�*��*��k&d������+t�Z#[Z���*����*9hj�*e�K�b�-(��X,��AX#b,V ��E-\��
)XTD��"(�Ĵ*Ċ�Q-�J�lE�DV�L��Pr�X��q�A"��V1Y�Ut[Q��TE]P����`��eb*�"�SbDDe�2%���cTL�-�t�T��*���\KD�L�32���5�L�$Xfa��T2�T��Ib�MQIY�w�Sޥ��:�9z�ٛ�
��ǹib��Kkiw�E�B:��3���/2=9�M��ā׃�бKs3RԐ�˺����d̄-@�o�ƈ�ϵ��N|¿u^"w�e�!N���]�����x�������8�{e��ʔ�!��:�(��<-B(�aXځh;�3��n����Wd�T`�TJ�sLK�J{X<��V<�ғx��ζlR���HU�L� ��9��u�3���
kۦ��E�iO��0���=��y՚����8�e�G���q��Q����c�]nnT"�Z}���L��	*��Y,N��=5`�Dy��>Z{��ҹ(p��S,;��m��ha�-h�lz�3�>"���5�����(��1zs;B�]�[{	^�H��l��uVb�w�ZǸ�b�5E�D�����4���b���[N�nZ���F4|L��wA�[7�=L�
����6]�5�/c5Ů��í�s�tr�>%�13{��=ݜ|t�6�_�o��О
��ߺ6"�ʆ#���ߩ��%j�\q�&j8F�QJAb��}��<X=;h�� Ϲ�j9co�,{ V�s�TD�ݫ}]a.-�Z�f�S�9�h>��Ӧ�1OE��u�x�{{m`����<��3��#Q��&s�M�;f�+>���x�Is���R�&o=�t/닔��v#�J=a�]+�^�[�U�\�(\�y{" �d�s���5�\�<�����8�l����V�ƶac=,d�B`uC�Z5s�dB.��	����9��8ysC�z�nt���+�1j�����e���X(V'W7�e�py�����U�U<j� LsQt�h}�bRg�G?��?�>�U�J8Z�қ�p��wJ�Kl��F�sNt0�s���Ku8�Bo����AEy%�$j�����J��8o۝;!Ш��h�|�[�5Z���f��\6`?*۶#�Ž"%�>ND�[����~���&��[-�{}��~��/ oǋ
G�^ҡ�wjL�f���n(�pٰȝ�M�L�4P��]J�=���;��֧�/���N5�jaJ¶�x��e_�6!�UԺ7F��f��'��^ j�F{Xs��Շu���h�n���D�����\�D�	����9ս��y
����K ݞJ��:���&{[����e&O�}�{nl'=�g��{�iDz�9�#�@Eo4���Lez�:+|�.ѕ��ٖ:�b�{��]F���X�'�Fw�����J���4?7^�*����r�pv���)[�����Ms�=+�k���r�ls��x���ؘ��ɵܡ;ݩ��O*�G;�A��;Kf��A.S٣\�.36����|Bn�C�)�W3%-\b�'�c�D�\��3o���v<��W�~~�+o_�����cFSx�]����c�oPY=-)��u(�Ǒ�h=�ڭ$׵�3Q*r`F��Р4�ce��o�l,}�4.�L�a|�9�������>u�x�vGo���N��A��O[���w�ۼÚ��B��=W�V��w=�J�z�o�Lø=%἞�Ǵ�nl�9yoȧs3��6�l�>'F�%�e>t����+5���<�*��Eq��$��ĳ��5i�܏����;���/�yO�{��]��ϟ6+�M�*����]�aI!��Ƥj{1�B9q��]��kdj:x�M�5H�4_�<I������t��_wF���v2r��O�{��ڋ��vfɜ����ni������Lt�ɲ^�f%+��W��0&�;i�y1]ؠ�ġrX�P#��05�pO�q�k8������3�p���*٘��*q}}7�,��)ӚE������aV�7�ii����U�+C݃rO�_Y��N��H�3v�0����U���FF�tnc�m�ק��YGu]*�h�
��Q�{�ܠ���C����z�n�[^Ң���3/��2�<�=P���J��ln�a<���-,�� OhN�;ʻ�zR�<�3k�Ie)�A����$z��1�r�t�㼥<鏻ts{�2�@R:�������D�=]�i�m$�K0��L��e����k�
�n��o�u�Vr�mc'�	/����n>--�P��Ұ�&c�ئ%�և�lӗY;ْ=���0�1���J��Վmц�(�����Xx;������|�oT�ܣ��Ú�Z�h�2�1)C��lL&=��P7��)z�Q���g�2j�ջ�ytz��m�����,^��.m<\o�ޛ�z�+�,�spZ8I�"�5~����8k��=��3��=����f|F��ho����SE�33���>V�e���u��MH�+��OoW���;ϧR�v/�+_x5�X+ؘ�	����sEx�V��r9F��O�U'�wA��际osH��{�*��g#^4���
Z k8�p(kV�ї�q���ҥ��sP�*i�w�x�-*������`�Z����k��)�(������w[/m��Y(�|Zf�ѹ{�ʕ<�pG^I?����1����T�3��@��}�R8�H���˚:-�޼�C]��j���e�T�)F�@�ޅ���z�c��e�[�Ty��%[��M)Һy'`>����i��A��±�}�=�h��)Y�r�ev�}�قw-ש �n���j���R�K�3�R�ǹ�)�{�grݸq�P���j�����Tvy)u
TN�1,�x� 6綺��$�O�;틚��'{>�6���mA���u~TÜ����9s��!�]+�`�)�D;�m�-6w�Ty�,vu�����ea1�eMx�W7��e`�MY��������wu'*bG�����iz�I���'�v+��v�f:^�ٸ\���v �u��U5��,OBҽx*Wz��<���b�d�q�+�ϵ^������=0�v�~~4��,�����[���,�^J���Af��b������<��"��{���=�0�O���
U�5��0f�:_�9�=�1$U��yq��Ν)3�A�-\�f	^{����� ��̦-�Y��c����N��}Q*`z�5�a^�r��ҵѵF�q}�f8L�;�["�qR��MZo���:ՃV����&7�L�T$��K&r	��7�v��}�7|�ފ�+׮���)`�C��a>f���vܨW K���Q�E�`��w�5{"�G��f!�{����.�K��J<����{��.���p����vH����e���t�p�,c��ͨ:�4OPw��0_G��mi���8�h����}��R�%T*�u�R�w����wrz��׬�Z=���퓚�쏱 {w��2�]�����G`������8�6n�0p�B�p+D9��2;.��>�T�uP������oҘ�Z�n��'.UwYٮ� �4���ٱ�o��U�9��z�d��u��K�p�ft�b��ݽ>���1����c|�]>�8��yU�ng>�a���M��,�bf��kJAd*����؅5�i�Sۈ
�}$�_�<��h>��S��Y�b�U_)�V����s҉�2T!8��+�j��"�K��PY�E^aFF�Z8����
�敔�:���C.��@ɠ��
�N�ol��'7���U����Y�:��29F=S�0O���'�s��\$��u��)�W�TAJ��#Kl��$�R�5Ww{�����q��-��ޅ�h_���nʮP��"P��Y�|rE�d�Ls��Ǐ�in李����2�U�����C�Q^J �acG���K[��.��m5�.�y*�Q��*y�' j�al�8�R�:Y�"Ѹ���l�_[�#��khf4�g}ϖ,�^}S{>�%V�8��X�8^�U�uK�]�M��N�����/�쌆R�v͛����-�rq�+��oXO:���]s�{%h7�Ώ���tլ2�u,o��N����[ʺ��ѹyfQ���xs�D��_3�N������%��C�M��j�������ǩ�a��C��l�Z�v*yD�������`<o$�P�7Z�5�lʦ��,�}v�'��F�k�&�7�x�z��
�z�|�b[aH�.3�ڞ���A&2{�m���Q��2���I����W~�J�N���ɓ<9Ț>�U��aDW�-ѝ��go�����A�X�o���&��\�u�+7������"�C��P� h&"K�j��I��~:�y��<�¸�m5og.�L��㴔>�+�q�].oȘɨ�g����\� �L�q�2n���b�/u7�#��sdG/���%zP�n6�Ɍ+���O0��������ڬ���*���3εa8�g1��ݒ�}��+T]^!?���Xj��X�I�]Bk��/ȗ.n5.w!7y0*Bcű�w셤e�WN�"���vA�K�NY������ܴbq?���cs�����.	�Uĕ�Wۺ���^N4*si�|/�ӑ!KU��A�9>|خ���R����Tί��b�Q�g9��U�`yM6q���9Cr�c�8�.���#R$m'�8�;��tH������vuM���z/�[�]7�D�=���b���<|�X9a6�݆�1k#�pJ���s])��+���xkW�AR���d��X���۶��0\q|���R�������Xҝ9���d��=�Ԕ�)r[���KN%]SsS�f���q�ޕx����4{N5����c���[�B]:��w~��v2���iA�U2�ژ��q��������3�w��(��9"ffbd�癓�����^Qwu�fs���׎�с\��Q���Z��0���>�w�-G��K�M��#�9�}�ae#����>�X&���1�0��)ie�hz(����_t��9b]�R�����̠���25�'��),�UY�WX@�to���q
�{:��S�t@B���@�,�_�oj��F(��eNL�u�~�:��,�h��{ۚ���������Tj���K(v�0���u��2����U3�0j��m�!{5�S6�k�	x*��Օ8�4�<���ffẼ�D�>c.�U���r0��X��_������a�,�4��bDƻ~7�UMW҉�b:?*��%��oM|��Le,�L���
�����mB5L��Z�;�dv`���l^ft�W��	�+5E�˻P6;�8��VI0�k�q�쥗�F�� %u��aV��w��U��պf'4��4��-��0_	^��G�ξ�,;I�c���ک��̊�v�ƺ��Y܊��D���'��'ڣ*6l�`e�(�oj�B�[E�cU9D�[�P�zj�<��B��N�AȄ���j�q-R�Da���'�J����C��F�U5�j]�B�q��O[�y7��ѳ�
�������r%�@ߢ�u�9Vfc�
����&��˩�K�-둱,Gc0ji�F��GS�5�j�pG^%�}�ga�ŧ��T^^����>����=�=�K	�1�kb%�qR�bF��J]B�:��K��<�3�C5��{y�~���z�\��<�DT��teMc1S^�R�������=���@�5����U�>@.L�'�㫠�gJ0n>�l�{��E��jva�j0���<��J빮�Ӽ�r����A��I�30��L��&Yخ�d	ڥY����'�W�@j����Y$�|W�bӃ�ݗ��V�+���#`>�t
!�����=����Wڝ�{8Υ�n�r-��Zcz剂�<�`���V"e,�G�xRl�$� �V��/1[�-[����fOX#�gH(Τ�iǻ��B�n��;�0fE�0#nVR������.��^0Ձ�ݯ-NX�������>�Ԙ�)�9�5Vk���.�@%�3`{�:�$9*k6�9�n\�P�����C�%�k���t�k2Q=���E�w��i�IOb<�-еF�o"LT��U�ZV_j��:}���wnѽ�`�&&8fey(x�t���TǪ;(�edu	B��yӗȟ>����*�׬H�ڄ*C�X�>��{�&Sp��ћ����+#��2����W��^ެ�����8F0B.v]�4c��w������zm YFC;��^1ę����s�T�Ɏ�u�Zz�0V���8ޗ0c�.naٗۗ�9K�^���}ck8�,c�
c��Lf+��V���W>�J���M7��z�P�r'��hw�t�)(�ϵ+ڙ�)����W�V a�:�Lld�vq�Ӥw�&�J�۰VD���{+Wr/���KK�fgU�9��)�����q)���_)�s��6}-�CͿ/nΠ�6��ȥ�4V�6���3X�P����U.k؝L�F2�)w���ATӕ�{~���UW`�C�)��(s��RzU)���b���bM�E��{��a�Ta�C+盵�C��YHpʙ&Ф�+���(4�Qͩn�@����o0����U��l\�q��܂Σ��[��E��.ːm�Z�$vΑ�����b�4Q�dݕ]�f�&�2v�OZSS9&R����t�f��U2�K+}�N&�)�,���3�o{�&������4��(��qg���޵��wx�3�J����7f%�cچ���m��3�Jr�ڎC3���Ӻ��YX#.)z�]�c]�*Q�8��̝mU�}�� �W��%�i�ϱ	�Z��n�TT�{�e����o|_X㣷@��rW:���T����Yݗ�cKv�8���L�c\�j��x�m�1WU�.�a�&n��X\�ҷ^*���@[�B�=o��8:��8`��ɺ�5ˌ��h�Mh��]E�o*�	��/��Mg�����¤�rx�X:NF��ʓ�t껫��cAG���+���m�0��ryj�:9�:כ�\*�b�e����CP��r���K;��I��v�r��v���Y]�T$��% R^;��P�{fn:��A����X���iT���K8�e_�D�S^1Mks77��pC9�98C�.E�PJ�0-�_H�ƃ�	����Y���S#��z�@�c*�]i�W�L�+WZ���� �w� ��չ�R�'%�v.�	Ӭ8.I/�n��#��>��{ {U��� [}y�K��;��6�qSh���㼠��-;r��5�2�f%��˯}'e�^���x�[Q�,
���yNd�ݕ/kt2�hWE.t������f���mc�r�^r+*�Ū��N�/���;��iC�)Lڏ��푳���u�����/�rjWA��pV��q-���6]`=�g.���Ώ	�|����e���_5"F'w���S���\
�7p��2�`±N�l��[ZS�M^Bz�ن�r�M�YZ^41����{�W�^W:�Lj��5��,#�F�c�o�����&����&u��7Ӧwuįq�۱#���8yt�$���"{�9��P�׭o\x.e_Q��B�f��33���-��X�wu���V<�cR�b�80>47�#����٬b����4�yygC�]��ysr���(T�(准�Tھ��}�{�{9�0��;����Xn��A�թ�Y�y�!؁U�s������0�����
�9�I�:��3�q�\�yp���X�p��ͭ33#(5]}k!OeqL�����hs�SԒ͝���Q��������W@�'1Q�ɅM%�qB(��nor���_��EM�A��'�_v<�=��s2��E��tx��ht�،��.��u�9�o3�������^13��|����Y�2�	�甥��܈j�B�<X����)��{b1yV �|վ��#���6J�c��p.o@r�4+ԴsT��'�ݝ��8&:卨2V^��f�9����w}��" �Fҿ0�
�,1*���PX���QCEӂ��*����c�U]%u��AE�V
�7)�������"�-EQ4q�ƫt�ի�XŎ�0uh�����VVV�3,(�t㦳V�փP��U-��㬕��D5ji�nf&�`�E�.2�Ak`�s����Ukh[je��BX�dX��m(�-
�(��c˙dS)AH�("�4�-(ĭE[�9L�Tc�F%bʋ(�Ym��,H�Z6Ԉ��Kj��R�V��%��U����e�P+D�ue�1ێ9\�Arʩ��-�-�[K��T��+Q�j�r����1ml��V�*T�)F�jZ[`*���XZ�q1kj-�Km-��B��i`V��2�i\�LB�-l�\�b�j�b�˗2�U�KB�5����bW�-�����J?_fcqovq��ai�z��,.Ӭ�u���+;�L��%]=豦��-e�w�N�������֝�/z���F�P�m�spY=|�b��±>�r� �*g"t�%a��&���pwmn��>�4Y�N~��8��\˘��������.#@c	��0�L�|&�t�`�Hmu�Tܱ<�����鴨lخ��~;��Eਸ਼z`R��`zh���%d��?��7�=*�'nnn�ޞ֪��(&f���U}Z�؉r��Rf�Y�!
�PlPRpɷ���Nb���5kE(?#O�[���8|�Xf����E9��Ε�]�骀5Y��+�E����jJ��W8��Y:�ߪ�˘Ș[#h�]�|�. t��	>�0�n�ٮ�9�7��﷟ܟթ��v�$�@ڸ�'�����d��XI�+-�Ll�=�Ӈ����ʉD9���~Z�蘅�Ft�Fv�����J�UżT;38�:�A�nw5���ԧ���
"��0e1���_a$C��.�v�
��d<���C�!s,-��F�t�@E�z5��n2��qr��/�_��2㩦NԜ�����wk69V[�ͺ��O��:�L��4��ʂ�Xӭ�I��z� �b���3�j^V��n�j��q��3@���w����:���I�B��9d#S.��꼳,<�K�qɍ�=�"gw!�q�t��Z���Nާ���63'g;��D�WrԈ�@�L�.�VaS=��s~D�[����βq�ۍ�v:P���v�.�/U����,8R����'��j��zǁ�u#�l^���rLxdu��q15����y�ɪ��s����׃=^�t�8X�C��K�.?*�j��u{΅���2���j�#O�k��!Ə����4^���܉��;��P���\"hw)T(���R����oXm��X�^�粰��y�x�i�/@�4o�(	�3�ǘ�Ƞe�UY���Kkk�쵭-���Q�k�,����]�V11���"��������q�s7�e*��㗲WX#�u�
%�e�v�%��r�g���3qm�NLK�4x�6�_J9�֐w �Z��zz��1P,��;?E�'�����9&���T�N�8����K�݇�h�η��P�#jv�yJ>�X�7=W�i����if^r񴣙������P~�Zvl��c<�Tˡ {�h� �|]�o����Ҵ�V�=���!ǎp�ź��z�0�j�=����5�oG��_T�����TEw)ˑ�T/��彉W5{�sh��k�����iw�U��������X폺���I]s�3�G/M�lP܂�(��w����{Vo:�k.�ݑ�9/'g3P��w�w�)�{�v�w8�U�蘗�%c��_6��	Gs�*rv~��v���|%y��7=�)k�:������Q�K���L&�]j�B呪���Ȑj}G)�AC����Q�� ߫y��l�<�:�On�5<f`"�A�O"f�1�ڭ$����|OT�b�V��o3��)�Et��pc%�敽c�=v�luT�}(����g�Y��S�G�Kk�(%y�0{���bI�-	r�Vz��	CЛ?u	=��p+G�WBT�bn�uc����w��N��o�t�u��5D��j����qE�O
��LJ��15$�^ޏont~�yjr��,Y��N��"Ň��i%���`�z�u�9Vfc��<�\���z_�Y3���N�0`Bl�O�H�*^qsҢڧ1��� B��.��~�gq�R�.�~�?���W�y�^��Y�}{Fb琙����4�*;<���1�f6T;(�����\u�n���G+��_�j����	-��2��9�@�A�=)�g���Y,���W��[f8��������8�gw�6��% �Ӹ�����z����5��O�gi�fK�t���� �tq��p)y=lT�=]�tpي3;"*kU�Ġ�h���[����@vT4C���_=Ԡ��i^�2�*}`'y)�N���˺���N��̩Wy�POm-@�Ld]�5��\ވhf��'Y�F�e���syGj��D�'��+�22IaY�h:��v��YBf��.��{%�&�_r;=ۻ�l{��a�=x�A]븡�J��
&A��ϋ>�X2�-8
��=:��w�'&`%�z�ݺJ�dۍW�F��^���X�*SȆ}+���FK��G��EMW�q�u�����K���|���'|ƽ��+R�*C��EX��B�!�N�T� �ްkO��|U!��s��#[e�,z���'I��D������g,�R�������y
��_���}�"���$.'��k��C\��6��@y>~ ��,e�γǳ����~�0,J�eV��S�R����jQ�g9LO��^(����p�[,�z��C�k�r��������HߢH�,�V� �<��ޙ�z�C���G�w�/D\�1�P��MĦ7A��5&6s�X=]ʸ8��/XΛ͑�lY<gc���a^���yT%���LcD�ױ���.�.�Xҩ��[�nf����:]�:-�H�*j����+�mY(Mo}�̞����k��}�N�VBgX��b����[�.� ��C���ޏ�Aq���TI��v �K�wU�IJ�<������'�=3�6W��q+Y�sr����d�5�K�v���h�[�`���s�{�t�y܅O���|��Y^���lO��B��}��
j�}�ˌ�$Ͷe��׸���6Ő=�"�8��J�3Q+��K��'S5˘��W�� �n�����V��8�iX�q�p�S�(s�b�\������\=�����y��+�'�؄��&�؝��h�A�9S��ACRvB�.\�x�S5:k���Q��=��7�I��h>+��fi1|7��~�.b��@�'�|2�1x�̷`>��|&�O�� �v�ʂ�f����N����U�[�X. rw��l���*۶!=�XX���ְ_b�\�uA`'�I�2�����������ؠ�y��[�{AP�;�&l�LE�qE
����=�P�]��7޵M.��#s͔p�\��u�8V����9#n$�t�H�6�1�]�'y���LM��:_��OQ���nU��Wd��qVv\�D��]���g���K��_I��� ��T� ��2��́����,ȴ�׀$�f7o��<w�b4�Þ�ޱצ�Jo8+ǔxh�li���|'�v�}W�f?B�և�)L��Q�7��Xr9�D��K����٧�C=uj2h�F�ef���Us���)-$l��rՙ�˱8�gR%�db/�����5a�gl=c���Ц����u���Ƀ�f�O�r�b�����L���E�펵�E����1�z���s�~��8�z��]Ԟ��į�Kګ�q��k�ȨB�4/�q��"�K����mP�^���{��w"��
����_m=ޗ7���bm�@�5�#&�{�G	2��w#Z�8�Og��ї�L��L��Fz��6�����9@s[~N�_|�&nxNI�oI}Ӷ�gd4��Hڎp�Q���������D�]Bk��-��1N���y�v�-�;��w���G�W��<0\oB\�q�N��ue���y�Q^q��7��ξ�����_)�h��]6������ ׵A��<��\%&�r��z��N-�j6�R�3N;U����q��lG��B��4�zJ�I�}&�=]�p�Î�L���zw��7A�礉R���D[J�sO&n0F˦6��-`�|e_!C�D�U���r�쳞X+zxf��3�im��D�Iy���8}�ָ���C�X,1���׷JW�۴W����z���p,O���KW��TZ�b��;y>�OH�ד:��������#���8zp������w̬X3횁��ѪTkP�#f��`�Y9��]ݹ;ӯ\� ����SJ	_2Ɔ�\g���+�}yg�-D�&՝G_9*OT���v�x��W��=�j�³:�;?G\�׵M��5�w2�|�en*x�����/Ǖڜ�bfD'Be�8���ߺú��V4M�U�L�0�����8���-�ذq&1��T��-���l3G��<���zK;O�Y�A��7�!<��kgn�e���^mg��\�%�蘆%q/UY�{�mц�4u�*rg۔���0�{}�One;�1�g-�����Q}(�r��ݾL'�Z��)h�Fw���9�g_+|��S�b�;��^S��5�M�oM��HU���w�X�X�orY�[z�1+��Iq�.CۑY;7��G�V��=�oǒ�������1�wToi��T��)����j���t��'��*6a��|�E��W
�=�aTwm���-��]z[��*iD��*ii�#���H�-R�Da�E�.�P��a�"�Q����n�+���tc��R�M"ۖ�ZW�
�JeZɚ]-��Rf�=Xn�+���O^��pi|��X�PF�saN�V�y���	�5/e�-�N�����.X4����/2����"`��CqRݰf`���6*wWf�Mf�98wwNsA=��/E�Va�t�62P��8=z��Ȗ��rY�	g�9yTb+��*��N��x���k�;3z�'<!k0x$�*6f���<�e/$�k��)`�o����mw[�m�%4��zcB��9�)3#Ш��� �ߧV�ĎN#2o�-$�v�`�1�,>wX6�DU���ʚ�b����a��9�LF��[^�����A(�}�V��	��\(s>u�Δ`�}��P��g�R�8&��4Q@���4���XC֗h2Py�ٛ������330�+<M'X6v��X�7��f�����/r�v+�T�Y��)pً���z�튺�w���w%������ce��Ƚ�2F�s̾J���ə��X��*bl�����Jyϥ`u4Q��Əz�M�����w+sd�vޥ�EkV�_�ܢw�{ҵ.���{�P��� �V�Xl,��׭U�������b����
�����Ĥ!੩�YyL5�h����5���Έ��u��{u�^���IP��'m��O��E&֪������h`�XbR,����P��vQ������J���w�S8���YP��� ��[N�M�ȁ
��:��u�~{��~�B�KȜNܤ_>fq���y�G�����GT���՜�P�-�Sj'�Gy�59����6���6|+�U������TEj3,�6���"�A	��o^-�%L�|���3Į6A�nK�;< �کha�-h�l{F<���9�i.���&�>%�J�������Y0/��Rd�T������[���P�Z�yVžr�{cW-IXهv��p/G�ƠP4��M�ct�hƁ^��d�# �����Ӹ�[�vNS+�1��2p�ˮ'Q��V������y8ֲ�W	r輵B�kO���1�;E��HA/��4&_(�s89��W�X��_alB�혦b 4͕�ԧ��~̱�[ԃ>�3��~��TX>���X�FK�P���޻�T���W�]Z��C��7r�|U9�a1�y�9�>*|1r�����p��q��`�<˩�=t�u�}۴��h�>L7�KP­A�!(.\�x�S1���f:��fFT��J�M��ON%Wӎ ڸ�������*-�@���B�4/=�Up���}�:�4ہ��wm�*+-AQg#ET�8�x����������S�U���x�ր���.�ņ���ӶE�h���
(��Y��h:�i�ɫO>��_NbqXʵ��VM�q6T�쏧�F9}�Dx�X����f�	�NԻ�Qꝡ���mD�B�w=����^�2p��;��̄^
�z`#�LF��E��2A����t���93;��~ڻG�7Q,5��n�g<ۇ[�{J��	ݩ3e�b���_�9���1e��`%��
𶮦���5��s'���Ԭ+l׌^�榵����3��_zv�\���n�qhsY�0���(:�Jq,�)N,.�riB���5�2��T^�>x���J���v*+}ҟSf���������*�i����*Cٻ��sPt�9+[�����U)�/�LC�ɢǶ:�nP�D��g6\��N�h��-�=9J�Z�g�^U�x\�R�Q�
"����^���*7;])|��~�Q�K�C5�,��8/�#�6�����t��D�MF�8͠e��#&�{����}�Q"�oQCY����ɚ�90��ёA��L�����O��wR�u}b���̂��^�>YÄ���}S�4�V��`!��E��̡��m7�W�߷��	!I��$�	'��B���$�	%�$ I?�	!I�IO���$����$��	!H��	!I��B���$��$ I,	!I�!$ I?�	!I�HIO�BH@��B����$��	!I�	!I���e5�*�a�7��!�?���}���� '��@$I(�TH *T ��(*@ D ��)I����Q@��TJ��
'ݝUD$�"�UJ���J��*� P)ER�ER���)R�(��)QT�)I)H�B@ i�H��@�QT��BH
E%$�j�*R%UQ*(�)B��IE"Qm�$��R R�*U
R�Ϊ��(  �UJUq�4�a�MCRTfISf��Hc b�H֡I��5)T#*0�b�I*T��E)A)W  � �S�Z�E,���Z��Ief�2k5 �-�EJ��4i�V# )46�E�d��UR���%$�n  J-��`jc
+X�UI)�*�j��A��U! � 
����6ֵf��U�آ��B$UJIm�� dJ��e3m� �m�m�P�3��Q (QB�P�+�
�
9�p� �B�g.�P�(9nP�(
;8�B�R��Kl P� 	�*�R�W �v���FY��j���eR�m-�� R���Mah���U*���6�YKU4�V��5�m�l-��TF �UP�(*UV� �*4Pl�SYZ�X Y�F��6
hkj2ڪ���@��Ԗ�ҡ��+Ya�Zh�6��%V)miTYRQ!J��R �kN  -��j��jj�")&�jҊha���Z��LV�Z�UA�[#5FVڭ�j5���@*��j�T��h*��P6b�UJ��   �ph�3im�+B����m�l�QZUS1m�ʖ+5lV�VV6ŵ��A��H�MFj5mj���j)Q��UDQ�  ;�%BUae(4�̢���L jIZ���@�j�Ed2��i[E`P�ՕF!��֕�*��BE"���  ;%
uf!l�5X�J�����
��V���j
�E�j�`�b�S`w� �!
O@2�$��� &�� ����@       "�O)��dOSe2� ��  PE?�% F	� C�Lb0� �A�2i��SѢ�z��=4$�HT�#j`�#L��F a����Ӿݽ�Κw����5�I�1XkJ1V����a����19( ":�K���dh���=g��n����`
#e>!UA++���J���d�A���#
��F" ":Di X"�E* "9���=�c����ϖ�
��\�B��k��Lp�ʇ��G�.�
h�x����Z^���9b�͵:����b���Y[��/]$j�
�6�B��(mjNTA�h� �H�U݊W�0�ؖ3�mÁ�"���3M���H����J�e�K���욳)���cp�U{�T빖���]vo�ӰA[xz�o)�Z-b9���m`��;��egc����C
��,˶�Bm���%����%n0t��X^̥��%f�S�1��Q�{2m���ǚ7Q�݆���2*7%�t*b�cp[*��۔U�,P�7vcx](&�3jx�t�2���6�1GkVV���vbX���\`m<�Z�ʹ�N�]���(�Y$0S�*íW ̷(l�e�J����N�";ζ�/^v�/�}C�*����C�c�ٚV���!�e*th�g:�w����jS���XB)kkZVٙx4�ʲ�P7x�r��.T�ӻ�sf�o��CD��2���V-L�I�X僫]�r\����0�8�]�&�"E)˭�ywz�[���%����7PAH��ݺ��oso@�G4�1��6�(\��ɍ�eF��z��V�M,���R���УK!���W��eZ��YGr�pȣt��3(;wi���+4N��v����SA���J��CM�Z1[�����p�6�&��M7Mܹ�f��C\�Yd�'M���%Ž�а1րi%�ҮK��gp����j/���;�ܬ7��z��%f�x�V��݅��ht�q�gl�I[J��X·\w(�U����.�	״�r�5[��;(�n�lkN�&��YyWY�
��=s�'�A���m�Xq%WV�*��3-�l7j��Shm��^�V�e:7�\-	i�W�X�wt٫��rҴ�7y���v͊(�f��Z�$.g^$�6M�Ic4vҼ��S�g:��΂8N���c�c�YU��0�͵�ko,��Z	�
&�)�.Ց�QȨ����[�צ��ǹ�}�,` �+�Q��c{V+tJom]D%�i*$RT	��e�u����0
=T��,#{�;k	ɬ�t�tt�l����H���*�&�NVa���KIb�[���`Ф\Ȗ�Hn��Z����4�TN;�*$���߈t��mv��ns4��X�Q�����9�f�+uN�P�M�zl�ݫ�d1Q���^��#4L�$���wm������cb�Ms�&�����̲q��P�Vc�L,��t�cl�����/`�6�!���Y���˦���R�ũ�َ�&��W[b�˫ɪ�5EM���[Ǡ�#ִ�X臇i���Z��Y�t	�ؚ�7�ET�
-�y`���,�	x^���	�\g�"�@5嘑�O�j �f�)nTN}����iE-���VD܏Un�!Mb�0�7O(sǤ��f*����(���Zv��(m��1-zJJW���,����S{���0��3k��z-���;Z6��p���$<����5s)Ѻ]L����k'4�h��ltz�+�tZ�w��f�,�U� �Ef��B�ōݽÉHԉA�&ZE���v�����4�Yauǎ�3���9����uͺ���b[���r�&VqS`cz�8�Z���R�6U���N�{��F��ZlԖTm^+�t�:*I&V�#�*�+/M��*a�wlʴ�Y� ��k�t�O��r���b��73V��F�Zjܧ7��Ś�j�����]��/�f�mT�f#/p}:�]HV60^dɎ�X�DIu����m�]`44�Ҳ�S��-����aU����!Ó%�݀��Vei�/]�Ң�Ŭ���,�vT�EѰ� ��Ԗ�� ���꘴4U �I4ajY5���;�lm�ƻ�-���±�P�(˽?�aS7�n��:�
�)m�H�\�D|0�c�jӦ�)��MQ� �Χ[�f�������������(��jY-:��JŸu�wp`[����&S��yhdͿ�t�z�c��Lm��;�y�`�4%��V&�F�t{c.�児�Eں��v0Pլڭ/k
j�����i8���Xi^�XȬ-�U����C���v����.��{n!e���WD���E��h����a�_9k�Ij��԰nQ�Pm�6��PIH;�)��z#�Q��+��.�D`��gXYx�d�B������,zЎ�����l�-	+tƴpX�&�((�'W��EbLZƕ����d6N71f�IPכF�kX'@"�E����.�772�n�`6��A:��Uť������w[�W[�+�͍��\+��-ޙ((]᛻"Ԗ�W�)����e:u�m���/5ut��ۖ� VR�۫ۘ7p�J�c �S���U`i4�¦eЀ��m|����QQ��F�F^}��P�d��>�q,ٙ�gQt���t�fv�����tڽ�m���4��M (>�kmM�vn0�+����UqiW����G�Eaf��ջ��e_ʞ��b�%ԓ�7(�[1�CfҪ��6�d��&��Y�xp�%(��+T��,;�6�U]�[x����̙�Y�.����lێ��Ch�`�23Yo*��B��&�8ܰlϯ-Yg.�d�(�^�c"�v<Yt��ÖhޣGd;���+�ԧ��D�ٺ���+p��QRi�/&dz*� iX SG6���e3�QE�(U��u��!x�T��ֲn�6�YwQ�:���Tr��0h�WB-XiwW���1JVVi5h�����ḭ�Vւ ����/M�в-�|5�eL��l����jk?gӂ/)�l��ث�rѨJ�Y�-������=��Fhx"�r�-[�<�ƫ:�1r�R#۰�W��6����Ot��6sW��9�'��|�cU�$��֪�ps�M���n�r�������%*f���dj�%,]x^鱑� �Ӕ����4ja+8�tl]���gN4Ly��XW�tҥm]���cP�Iwk	E�7jʧ,�� �W��y�簚	���B�Dɢ�7]����F`/-��� �yn�W��Cɲ6�-���ܽ��E8p�Zi�^���,��������Q�;�/(�{�F�]��*�v)��.���m6W4�Y��qԨt`͎ӕ��-����-�c���N�]ٵ�4c�a��W��ɶ,Qm�w�{}Y�g��X��t�q�Y�J@��WK1�hC�P���,=f�{�77����=�&��Z�
���"�����tƄ���b�2���9�f%��I���2���ReL\Q�v�I�i�f�0�U5�c�� U^��V]��-u��r\A�*�e-�à�^�0)SզGu���GN���ʿ�ƶ���L��j��,5��3�ɺ쬵w[@n;Ư
k�5�th����[K0��t=�[���Xd2�%�0��j8�ܛ[n�R��ܗkndő@f�2p1�1TZ,k~Ż�$@��H�۲v��@����9g �9|V����N�<�eӍ�[km�CF��� ��L�/!hٶ�݃2#��98b���3v� A�X�.4@�h(]�O���l"y�3�g�U_��m9.Kt�Yl�2򁗔l
Ċ�z*�#�Gk&�7N���i��QR��m��/h�rk��Tl˴���֐Wbo�i)��κ�,��Ǹ�M�IDk����%�^M�ZA�z54���(�	o�r���iv�-��zS搾x�SV52.�ݭh���H�j��<Vi�@8j��f+5��i�0F`T��M�K�P�,�a��*nj{d*Ȗl���ܶ:˲F��o�����v]�2�^���L�FPm�Yv���H�l[�v@[Yg�q)�2u��)7x�*ZH|�6v�V�&;�Z�;n�e$;F�:=V�a�"��x�/s)ݥ6��Q��k1�z+;+7Z�(F2]8����ej9�ͧ�
��%BH�lnn�ͬ�P6�U��#S�,��2	/-J�Xqݖ�h��-&�DL�zIYP8+*��,n ��j�D��J�F�m�9��)��=؃�;*=��ʭ�2�,�U��F]'�]��z�Y���p�L�ۼ�$ႎ�`��좕��e�ڶE�d��B-H�u1���PͺYV1��1H�3�|q��k���A��R�a����tCܽq٦U;wk�K#����.�.��9IW&�Mݥէ9n��ES7u��S�bB�ӻ���KR��i���@6�ҫ�NDXy������h՛oQ��5��,����h�l�㹶Y���+���GQ�oY&�Qy��`��U�w��R�f��la
``��ʻ�5�n6�[��.	�Y�>u�3!��ŏ]z BM ѻ �	��A�%����]fS�n��Vw[�V���1[�v��z�M��S�Y@fR����gv������Nܼ#.��9J�YE����<��e&��a���Un�,Kxi�5�n�N����6s$Jd(�Ӡ2��F
t��B�TX`��#b��Wug*ލ��,3)��n�X٢���֦�hj��z)c�@�����h�e�[��'n���{^O{[�M�j9]��l��Vf�C3c:����mJ��٬X*�u΀-���W�[���M����P���z2�4)]	[Yg��C=�Y{�4�	!"�Ǎ��p�6=d���ƅ���I��b�	���I�5�e�lnǸ���߉n�U��ۭ��h��Z3����ٱ\�ʹ�f`!:&�\��.V�8B���@����olX��0M,Wj5��y�Ս�"��Zf�匉"�ɋv��of��.�?D&���E�7fȆ^��$��B�����17]T�%�1�=j�A�6���L���Ք�OV�|os�ZЧ�b�g�E������d]�x��*���&c� �x�5Lf��q �7�b��nS'Ju��k��́�ބ�W:7}�wot��`�Ve��"f��H��ؐ��YL֦n�A��aKQQ����g5
����&��@�^�xP	�x�Z�m˨s%�1����!1z㗂���ܼ�nՠ�I��bԵ�ZY�����H Vٻz�urS�{�f��U��t3#��-�4�|Wݘ] ��j˼<P�&�gQ�)�Qd7�ɕ�B�[m�7*m�t��p�j;:��n-�kr��P��U��x��si�C~)Mٱ�7Ebx��wKSXBز0�e�$��XR�7��^ݍO~�P�<�W�TĮ��\_G�*ٵ�q�i��Z1���F�͟#���؍�f��'�Swo�@�yB�n`��1��,�ë)E�1�B�r��bޙ@n�t�3Q�I�ͦjZ ��WI3NIJ�DW��J��_���2�P�Ń�Y7^7�0P�b7�v���3Zݚ5f�zWs����"��J�������Vm4DqI��qD��xj��`��f��\�[���t6�9QZC@)i�O,5�/�.�y�e�v��	���d9�U�6𱺫$q�4P�T��lƒ�X��V"oN���v�9x�ɉ� �L	wf�UGW���-��V1�+�ʰ��+�{�|p���A���9V�̓V�鄱s@	3�؎�{������e]Iq�_�A�&���n��:f*�1c��,m²�JԐ�,��y`U�h\L�{1O��j��V��c�O�Ӳ��.�3���,<������Cee֩���ر��$�uen	I�Պ &�m(p���IY2�v/vŕ��B����i�{�0���m]:�V4�Ƶ,�����́щ8���.��ld#hf��V���4�&�T!��*/i��mY��$�{�mP���q�.2�%*Ƚy��ԥ$�e��2;c��e$Ŗ(�n�� �H�&���oXɪB���a��c˶��u}���|:�c��<�� �4����������r�4�%g(����`sX��n�u��<ɯ&h�]9��#?x�Pϟ��:N:��Q��X�o.[�8�.E�m���bRP�r)*�i1�
c�)NF)M�V���"9���A�]���8��Ml:�+;q5}x��&j�ɤ�%b_fj�W�T��^��V�/�^e�͇��˷k��J��\��R�N9lḙ��s���ѫ�ս�)=Fd��<N%E���-c�cj-;�TJ(_L�\��mvp�\�E���]�԰�h���Lȫ��ɴO( W�g=yѪ�%&f��xպ�&�����՛5���V��ڊbnQ�(���(GeXbj\�Φt���[/*|/ŏ/q�X�42�.��6]'����(�g���4r�N����)��%D�}J��B+{���}�8_$��}b�̙y���^_rw������S5Nb�&���TC�M�<v[ݾ'�z�K��*S�ɥ���ٸ0�lP|z�^`%0>kc�O`���{إ�p�*�(��ڣ�#8�9���sʆ��r}ڝg.��m�Yt���{3^����@9!1<]�KO3OW\u|8r��f�mY|Ȕb80��)^��"�ޮ��ێm�}2��Q)d�3X�&]�`q^�/U�9���{�s����9��Z���`�S&ǘ�V���6��%��Y\c���e��9yϢ�޾��VZǲ�j��fU��)6[�I�����S\�ݏy^�V�:l5��
���/�@ZoG#X�&�]�b��U�t��[����*2��d��tzKޫWm*8�V�.�]��&�F7��<��:���'Wvё\�e�Yd\�^'�6�d�'{b��Lɑb(��\F�f�Y���8m�j���<����Z�Gv-�u{�92���p�k%���B̹�+�t�Q}�)l,��R�JnBK<�0b�h�+�<��hqW7��K��F��#����z��0����\K��X��v%q���&�[e� ��q�+/^*)oҺ�F�� ÷Ɂ�	Q����U�6���ְ�V�ka͋���̤��B��n&Z�eWmNי�����>#	@���;Y�MU�$�ة�%Ga�F��j�q��^U*B���V
{u�T{,mH�a�����nX����Y��lo(SL]�\W|��&�n�m��7��wQ7x�)f�{���סjm�T��	魟mWY0�W��(n�km�Ʊ�Y�#��=
ɺ�m�Β:t�E`�aF�]��삨�iyEt���J�!�cA���q�}�o�N@�5��.��E82���Zs��`��8�G8����4�mE��xE�!U���E��1���uq`;hWTE�+��ʽ�n�m�77��m�<��:A/]���`��J>��������j�&�%#gC��󬽤��:o ����S�+rY��k.�V;4ܠ9����HX�{������*�.Qw�vhޤ�-���:�8���{O:C�A�jK����K�2r��x70:Hr�jKgqb��A�)/�b�ƵTH�B�M�Wp����]���<W�(�@y�;w�,U���u�X�s"M�����d��:żK��S
�eE{��w�o��%%�H�o� n�-�
^��g�����qWR�r�^�{d�D�<);��\7�;��޴�v1Ѯ�&���zWB�����fq.e�uǒB��]ҪR�qV>���G�7~�����f��N�3Y4)����E`�]W�r�W/
AV�`]�u;�LoaN;���Е�B��!Y����ci�����3�7�Vlu7M�Pq�U�O�o2+f��DK��奜�'M7E�飆�VP��XFkq;n�70�8�����5o�"�ή����;@��X�̱���є�eaŷܭ������l�J�u����L:D�6H*-��-�����2�����_e�%��1�]�?B��88��of73�Qu��ϋ������ǹ���d˟t�*S}�e��.��b��7�'Ӯ^|��x��&˝R�m�1�ä���!��:�kT��p-y�i���⍻\݄�J�����u�SK���R��/���hޮ6������EW�n���9�z��a�w�R���P!��+�0
�j3��ɮ��KF\w:/][|Z��V����K:v��^�%Ѥ�`⼸�gȝ}B޾��k�ݫ�lL\��S��ҊS,�t��Gy:��.��lc�n���k�*��H���e&���	1�,r�;W:�ʅa�6�%4�9un�惔�%g<wiRݽ��ݝ��6ݜS�j�Am�S��f��-����&�mE��/�'�w�ɺVdʾ�� g9f�ޮ�6o�2n���k�V�e���a�o�}�9ɵ�fTYc��ߠ�k��H�^�SU
��ۏ>�]��NX�������{V�����v@���Y-��R�`�D������v���S��@^Z�]ˡ|+J�]��c����E����=��n�:�� pr��p;��M���T��X��L�:>�ԕ�ZJ�p�,��!5l�����V���1�r�n���ku�����-�\w:^�
.@�{�����0�RS5)�ܖ�D��v��˖.\}�yݷ�-��NY���y�93���h���]q�bt����'��U�a��C���j^n��f��g;i�{q�(f�oD>ka�S��rwsIL�8:wph�9�v���GZj���C���&A�̡H��%M��bH���{�wk����KS��8\����`9\O�P�q�p�R9�&����r�)]Mn|y�u�q8�!ִ�o�f�RJ��d���[u�Tl�vcƢ�a��W[�i����Qj�9a'f%E�q{rE�Xhʾzs��Ld�x�i�8/8�L��*�^B�!r��w�]ֻ/��`36�\`�.������I.7P��#���N���e�����<Ȋ���<B���jm戔%*AH��mK.T�*06�(�Qt��o>器�4�?8{���̫�S�v�f����n�c��P;��Q����^w��=�-Rh ��5E5��3�:���M�+B:>�V��,k��렺�W�ʝ�����%z���n�E��P�����X�ͺ�m���6�L�a͘���jJ�ؕj�F���1�X�C�B����;#sfrYx�a�I�4���dG7 HRU�v`ii->����b���h�C��{	6��	�Y+1u�^���$'�D�����g_c{H�5�x��9%'�G_b�����J<*_0���p��bzP)�3{L+>�u'�M[�[��A1d�RmoM]7����N�|��@�o�mԬ����xM�1Q��}�/�YN0g#q�ȷ�q���&<p^T��\�ۤt)��T��n��e�s�eb�/+����Ok8op�D�5�C���o6�[w��<"TcU.�+���ݗ�	4r��\;��q���H��c-�+@��h�Zٌ_v�rHB
^u���38V�5u�`u�E*�*'��׽�.��IJ]���v��խ�����虡G�4�&�����}�࡝�k�c1�m�v�P�����,� ����S \�6��xn[�k���.R�'D��CW9�� �ї�j�n��ʰ�].���JoT�7T��ӖXKϺ�
��\��w�����n�.�*-(�� ��b�Ι�@U:1��,�����w��e�,�4��γBZ-����yu��`�CYs��(����ΧZE"Vs�=���-��(�2,x�Y�X�z�H���������IWf5�uf�{��v�u����r���kQ�aQ*���8x6K]�����;���H�I��.�I�Y1m���ۙ�j����Y��kpJ�т��Q�U�i�%��ЃR�s�/1����H99��|֧d��[��r�.�)l�5�<Ԯ�372M�gj�n`�6wT�|�sP�B6k����z��C �1p�L��ش����:mUʴ�]c��3v�Mj�<�̲NYk�R�X3Pg����l9�H="���2��[���@�jV��\W�١��U�tۧ���^����\t��w��q�9�Z%�8kE$[{��\R9\x`u�I�K�ݸ��,t;�<]�R�̺3L}xwT�llp�F���ʖe�R�l��r��L�ju�"�Fڥ�Cx�U�RVn�\W�:� ���-��>�x��w�eKj	���=s�F�޸2�	�V.�[+)s'*ٜ�&;�K�-��wR4�6�|+�S���9��n�Ƣ�e&n�KK�Vv<;[1L
�l�w��/�v!�!d�;�ٹ�&^��Ie����%N�j���+;��Q!ΦQ;���c��3�W|�.H̤X�m��-���� �
ވ��դ_��G6�d8�
ʑmm�#ee^8��7N�oS�qTF!�ɤ�gU��1�2�U5S�%kx6d��v�'�@'��޽������ ��Tn.|�y�eĻ����ݵHE-K�v�u���2&���i�l.��e����[���;c�l+0���cVR�,�8/)δ$�Y�W/[��'���S)o���MW�ꗁ�A�')Z7mS�J�[V�AQ-��.�L��1U��X�Z�aG�&�)�qq�&�Ü���V�9'94�ڣ��[�WVs��c�3q.�ͨ��}�k�R�X����TM�S��9q��c{ �l!���d���"/��^�W�V�uv�k{q��+�T��$�*����o�'}���5G����r_n*�S���u8pC�`�~+����=�=�N3�tq�8m�#qNF �*5��N�v���s����t�[{��$:i:��є�Rh�10,��
�g&��x�&���r�#c�걯i�ˑ�N���+H:�y^c��2�,�l����C��<;mu�-͗�Y�vNU�GR�)��pV󵴧)QV67;UO����m04����	�͋���w�L����ıL��t�7UC�e�A����#]�w`����ȝ�� D�b�d�;���>4�5tS��,}�"����(�r9�i�{J:R�·�0�a�Z���Y����1�շ�{`�bS�u(��y|��!�*q+8U�������*�a0C�kE�Ty՗�.�:�b0V�o 8�c�|��{����c�sPq��A*�����Kx�Tź�"�Y�����ȱ����r�!�/H1}kH����tU;vq�$�n��h��`��k�s���H�n>T��3]�|��9)T�� R�I>h�k)>Ŏ���6�p��%��1E�]�MI��J�aɁ�q�C�-��3#��\[�Z֖����Z0���d�{�*���[��%�\^���`]^-п��#�{[�~vbܻos�,�8^<�C����e��Lɷ#�!\��7"�1�u�.ʨ��#���#r@lZ3LoFas;I����A;!����j@N�b��#bv�`�1b����ԝ�yP�������x�M���,��o'!
K�t+F�EI�f>.���4�2�&S4�)W��Z1�n �q0�E��yiy����mY�֦�wv��\8�P�H�GYy��w-��D�˭�\�%�.s�BT�������A╒�95&-t�۾ᔋ�����&6�Y�����{v���䫗�C�+v����`��t0ofլf#�Ł��$ήM�׈^�^�K۔P�s-�Cy�H��-S
�+r2�4ÿ���%7"��kȵ�:�4Ҙq��5����SLW��3���`k80J���Sf�D��q*���[��+�)���d���A�>��$,��5�!��6�b���h��B�[
i��`oW'Q���>�²�."&�5�b�ev��%Kl^2
�枛�O����9ըR�W7�����4W+u;�!�H��lޭ�AP�]]K�{�ݐ#���[3��ijڗE��s�vК���ץ���8��L�RJ�<�y�
��۸�빕�.�֭u�h��#��;�ݛ�����+�^gr�/���/�;�ݏ��@PG���[]2����k"`�zCqdG��5z�p�է(�q���nH�	�'v����AG��5��B�u��#�iwjY{3m�μ��ް:�v7�u���0�h[��#K�^�s4;��v� �reʃ/���쥑3O�L�ɿu��!�z�eΨ��3XW+��]�q�7ZwY�����E|WS�D�Knɹ*�X75�B�%�a}u;{b[}�" G���f��z���N�*�����DP�7(H��o�]���ϲta� �:0�u�D��ɸ���I�ŅӁ�M�u��\|���ǅ,�u�+�ܢN#|@o�-���OYx��d8�������Y�kA��2D���Y�kA��.mfw.-!��d����M�t���	k6��įe;�B�f�{�N��Y��s��|L�Nn�/���)fJ,�+�oN���,|Z�	�v���!��h�Im��.���U�XU�ՉW�n�]�9� A�p�SΒ@��0�U�Ve�Q�@�����+4�r���V�,+r2ЫY�z��v�.�\��P�Fge���$RJ�G;�g;1tSyqA3����̏��%�XΊ�Ș�!���H���7��:�gU�1WoZ��:�R�����AWV�4��U�+݂�jid���A)G�+B�����L˺��C-*�m�t��6�F��F��"^����Ü��T4�j�b�kl���W3��6J��X�����v����:r���)ذ�]Ðb`9�+�s��Jv��/[����p�s�l�2K���@I�8_^��J�����{�ϥ��9�AWVfl
^Ek$���hb��WY'WnG��� .���r�k����v��]t��p��BM��]1iE/q���P��7Sj�^�1&�r��V;ω��l�:�-G,E�����	��+?L��0�3�_�B�Y�b�jeƞ��ͬn��E���v�ʶq����o�'j�.*fY���P���U�ź�{SU�6# �Ne�\�u6�J�^$j�L�Kx��{r�k�P/q!�j <�!�ܥ�Z�[ �'Ud�7��n$�twV�er�bN�c0��j�%)�\�����K��-P�޳���u����f����V��v9R��d�E2��^C�*��v��u�r��b�p���(��iU��"df���fkw��1{���'%[�|���#G��{Z��wd���B��2Uϰ`����H�wY�WX�q]e1ɻ�b����sp]w!1"qI���?=����;V2�=Ӭ? �V�!�V�J���W7��73��L����o�JU��v�n�=	��y|��
]� ��țk2Vm=yd1�"�eӽ�//�i��岊חVc��8��l�N���eg��wQ�B��T�,�K��]��.����sPs/�x֡��fV�yO��8�q�>Y��Fkd+�#[�IK@���r��;�����yc�:��
�t�3� U�<�F�3���gQ�h�N�t�d�A���m"��-ϙ�<�h������Y)f'{�f�L#�y!7�s��������M�	�y7�f��;q�Nq����k5%Z��b�+e4�J�P�.D� �׼<AfQYi��ɭ�[��[`�hW0m���r/KX�[hV��C8��"�+�z��*�_r<����Y:Q5�
�jR)Lע�VɪB�o.W��z�C@WJZ�u�����&N���ei#��Z��V��i�Z'u�\f�+�:�mm4�4������w�(�m��-|�!���?���N��z,�W����e��bCM���:}r�3��/��Vp�#x��w�LY�Q-
�Gmʸ�=X*�0�:�٠����Z=0vIË��']�'4�`��qξ�X,����ټ��3�q�0��_X��� ����.n�˺� �d��t�/�k3b�f�N�Y��u�P�b��\yu�>f���\7@�=�o��J��e����wW&��z�s��l�J*��m��RqP������5��Y�����lZ��V�S�G��*&�*Z��j���N��:���4�Q343;����ͱ�	j�[z���"МB 
����K�C!���\s�V:�PR�em�oD��ϝΚ�RͰ�U��0>Z�[]ק�A�]:��16���j�u�z��x�ڥ\/S�H.���k�uK�ڞn宇I������{�!�a(s���(�T/�h�yl;��)%��3�qe�������'
6���(Q�����f䏒����\����x��Lт��l+Tc�!�3�4TU{�m#��"�1 �P�-��{dε5��D��f]@Z��Q�� ��m��R�:�*�b![� x��HO>�䳄�7��9�X�447���fX�v�M�k�	r*z)le�����j�E��r�hv��xB}���8V�:�d2>uc.%x�n`U>hսxasNЙ2Ҿf]JW�Yg2��7\cP����D��s��yb����ZlA�ʋ�Q�ku���9��d�tj�ܲ#�J-��k���ӣg�r��	 �y�w+79:S7;c���ӽ��)aX�>C:XI�UJ9��:���˰�+@e�++���^ۻ���voBFZ>�d�y�:Q�M��Z{81JM�#��!�.�V�d�� ��J>��Y|Y����b;׏Y�ˊ�oW2z����R�EP�;�^��m
�\z�rm��Z�,_6ep�	|Ș��3V�Wol�&PՈ�`��q9�|ֽ�q�N�B�9e��w�k��ۻ��:��;� ՝�]�/:]�J��i+HLX���f6��gUŋ�`ÛA����;ԋ[>��^�˫9<�
v�'�+�+[��7�)�rLN��)�u�gpu�4��X����xE��gu�����Uˬ������u��Jg5��4>��WMIv$*�vv�������s%T����{9֪�t�M�Frx^;��ևԷZ�u�1��1�d��;�-%,��VS�J�Z�o.ih����P�J6v��u��CZy���3��Y6�ci@�k6����5qYXZ����U�R�>ró;�j��z1ދ��^�˩+"ԩ��hb�v�[vn.m��3l4:��ǻʳaE+�*��䧆��-Z���]p�R�nT;���X�Ӊfn�r��hG!��s�ge��H�Sӽ�M�c��W7M@l^.<�8VK�Y�$���][�/�^�Urܨ�[��
3���Z�����A3}rV��gbϗ��z��G���Dݤ����w�x�P�n��W�
Ҧ���;�J�@���Ӭ� �;��#Z�.�i��G9�˚�v�`G�_7��]+B���Iwo�|���C]�ZrcKnRj�ʻL^�f���(k�{ϲ�m�mm�$d��ṉ���Q�-N�̪�Dj���GM�]Y�Ҽց��1�0o�ic�>6*l܀:�=�OR_B��׻P�4�3���c3oH�`�u
��A�x���OyU�{9���l+�'6]���v^��>T�F���������յ�˕%$���v�L	�;�����A#���7r-l�t7&�Qof�)Q��t��i:���Z3��cb�.P��H2 ŪT���Y�\��h�Yt3��aD�m^�k�}��m[�;��o��B���R\�q���ܵ��K�����"㩷.����
c,y�Y�A��]�ٌZ���t�Qrб�Kc��ŕ�h���HF�$k)�)⭊�Ls�����:f�g,4H]��d�p5K�{ot�5[U=�82��N���;�
��2��3�QR�r��j��L�nm)�j!2�2�̲��b����E1�< �n�v�luX�Uω}�e�)ZĘ4�n��c��u�7�x�U��8���u���R�%5Ӗ8).͔�����鉶f�\��Y�G�q�p�ߒ�ɨ��*e�����&����+�-ɹ���M	��jԥ�QV������@"�����V��-$kRh��u�ї��u+�
̜2�	��e���ks;l=@���w���|h�jh�٩u���zf������w�^��)M��Rr��W�<��oK��4�3;�y��	wuuw�@�q$�U�Ki@U�+3b�Ȍz�Y���S��w��
�R�o>�^`R��NN�(�������c.��w`^
�fH�Pr��2֋�a�[ʃ�e���k¹e"��Y ��`�jܗ��ЭWoA��MI8�7W���Y���P�8	jL�aڰ�l�[PH��WMФYu���ƞ9>��຦>r�m���q�`��t-����6��K��Ⱥɕ�d��K9�{U�?�05_1xƌ@�V ��oU]�Ee=�]CY;��N���m�0�5]�n^t�Wz�NG��:�������-q=�>={���bvjbT���h�;��X����|�\�h��<D�Xt�`wvuf	��RBJ�i4��׃%]�-ONn��R�j|�]��*��.%�!XˢX�[*�eN-
��,�����W��3W��b�&^��<9z-a�L����K�:Y�A�Y�E�B<�'
������]j�%�cyBQ�w|^F��Ds"ְ�]����v*.b��.�h�w�Y�,�HI&�o+��M�f�Y&W0wo��Ӝ�%;0��:\�6�iI$0�����U�1^�'��Uu�
׈R��$��3`��w>�ab�\��C�u
��2P�Uh�E]l����aK������m�&��;k���W��ک"ĩ��&nZ�a8��8k�R��8�T�h`B�
T��ʰXc���J��N��M��޾��Hޚ9�6���p�Z�%>��;�j]/m�`
��OOX���6J����U�m��lǃ�:�Ւ#c�ᬕ�� ��\N�n�dIRiw.�Un��"Wh
�ܲ5(̬uyc�cA9�n�K��2ƙ�>�rG3��N�9r%ڵ�TU/sau8KB���*�:��v�]!y�tP.�v*�	%(��W���YI$�r7��Ի�r7��1��Z���F��7E��w����#s5����.�����E����5yN�Y)�����7\�  ��\T�i{�,Gb��5�a=%��;�Qz�bxyu�ȉ8�oul��:�Y*��P�Ȳĸ�X���XF&�se�Q����[�	��2�Ղ�ƮԩԍY|iR�);)VE;��/�։װ f[X�������9[W�����������BZI��H��a�ї@�Q\�� kHY��\r²��{4��yiX��evK�f��y�)�ZƹҜ�� �����D�;�GjVS粹ز�8��IHS��&VU�T��,�҈7�4�۴麰_)�����.gf�o%��K#�����1S9�&�_j����3��qL�֠;v�ύ;�ձ](C�s%+��nT�`�_՚��v��퉫)M�
��>P;��U똕%�@7���&-��7��2뭽�JXF���nSHU��q�V�_��)����v�H5����F�.Z�*]r�]���T:{p�/#3��a:�p�-2��fZ��8����5|�p��k�j�q�z��Ӽ3f�c��w���R�#�V1j�ĉS:�39���B��B�����wK*Β����N�t��k���K�˛�.�A�Ze�\c5>�|*]^i}�u�{��pV��@�H�\�l�x@҃ieK���F�3�l]fɆ���8��˞b��J��
�]�C�I䨱w�KˏQ�}��
f˥T���3���}R�&0K�-����i�X�n!�řtYNS� *���Hb��sc:��PK��WL"�L`-N�_�Zܺ<�D�ֳ��כ�JC��e�d@ӻ4k�;\�UZxĬ���/�]-���R�Ի�nr+��T��I�o5��V�U�u���%W�l���;���F�9*�7�#Ϩ:�\�w>b,�u�9��RobgUN��<'�$�!T��h�)y�{\{���?/~��ch�̵�=�/��W���>�
�c�q�2�#�C��]uհ�C�nv�a��|
�4�I�Ȩ�eh:]֛�Z��ĨW,��P�|����2���������Y8���z��]v�4v�z�-�Т�h���j]u�ʏF�)/F���[7Spfn�n�T�q[38<`ǚ��	�ܮ	�e˹HV��mL� ����,_m�cjrz�pշb��6U�qvY��e=ޙ`$)|-�r΢�u����Z��a�-gv1L,��or�������xIZy�a�eu8����01�izM�y��tL����;\� r�����&�]���=�0v��]�	�2�G�\��f�8-fe�jJ^���?^|� �&b<W�˄�0�m�`�!��Zj�>DMB�h�,V��^��4�!�hQQw�S�D.3i�g��Ŝ���X�q[D;0�������A���E@.N�T��Q�]�y�l.�|��+#"����J��\hv�U_2]cJ�r�ٸ�9I��s���i뎌��HÝ������z8Q9�2��:��SPG%��ms�/l'm������d9m;�k^Q������������Ob/���V)�*�+S�Tb�DQV`(�X��(�T��h��ƪQAT��X��E
�LiZ�)mET��X�M!QTVQb�۬��"6��kY��RQR(�*��(��TD���l*�EF�ŌQ2�*�Q�*�KZ��q+H�Z�X*��0Q��+"1\j"*�`ł*(2�D`��j�Ɗj���QQF)Db�Db�X�U��)`����U`�X���iA�
"������mPb�S�r����Z1DĠ���EUE"�"���Ƣ*����PA1���*"*"��*�PZ�b��`��UAAJ�2��YZ�PL�"�b�Ķ�+�
��E�lDF�*>>�O������*�L�ű}��e�GH2c;�n����{i���N����N�����y���͋�_-���/�����哰����!)d4����:<�"���^F�|E��;��>ކj�B�s}��d:��U�o��UN��[�Z��� �ygʫ�7��E8�"[��K\O�d����y��n�O����6J�u<࠭�0������f��y3�ӕ�>�6�g���@B�"]OTh-@�{z�*y�S���ڭ]"ӽ�ْ{��+��I���ul�-{�C�}�#��"�KI׭l���z�;T���P�-ZU�R��t�-��=��ˆ<��?qK8�����c���ͦ�G������Ӟ�]쀥^b�4�]{b���9{�0�o���Փ�N�f��ض��d@ֺ�/�.T��u��÷�����_~��d�v��e����.�[�Y{�(ȹJ�Mg�G,p�ʺ](u���|�U�ɨ�-�[��e�)Ek$"؋������u'�li�w�`�"�}�W�M�)���8^z8X�e��ndw\�j��t)4=I��ȑӲ�-Cܕޫ8�(�`b\�a7kR���1nЎ�FZ<�:�:�n}tGV|
�HU3�֌���Z�ʐ-�D��϶W� ��:N�����S�Jw�ߟ�0�g2��^��8Ԝ�{Ī�2��G�(PgC3F=6��իy�蓕����S�g6�EfUx�k�l�����Zp����,J��پM�;�l��+���O��M�󬕯A�mZobѭ����2�����+��fm�oɸ;�uj��\>�xF�wz��~�ӝ��'���\���gx���F�B��^��"���D�&ל{'�\}��uB���V���c��w�7ȝ����y^�󭬞k�cՊ[�ה-fs	%rg5���zyU8wjd�������cY{+
̱{*��#�	N�"�G{�jC^Lw+��[ ��FY~r�e�Q|�X��i2*y\�u�=x8���=D��Y+��bs���]l�a���'��PN�;�[��4G�2���c���L����F8߆��g�S�ō�����%��ͷ�9�����b��*��.R�5��R�-%X����p��#{�a��n&�-�������uݵ8�6('�mϩ"'�U����9���ej�q�X}-~-۰!܍NGgUzQP��M[���r����չ������U���<�hM���s�T�k�AG:Ԕő�ۋ��
~�[l��րu.>u[ֻ���NtJ���y>�����l츽q˴�	�r���Q7T���ű1�6u7x�\ar�f>y�Xr*@�eP���6:���o�i����ډL���
��!���։aGr����]%�ohsT�
PԶ�1j�����g�L���g(%Э���s@F��ʲt�����5�B ٸŝ���W��Yy����:��a����m<B[7:E&D�A݈�Z�;�ţ3�=�b���pMJ��t��K9ܣNu�%NYk��9�+��)�����r��]V�ئ7�H��{w�;2�]�l���+X��!c�ޝ�|a˛w8rKP�'��ǣ{�A+��/<t���j�V�y倓����6c1�v������\v���[�!V�~����T5<���)c�p�-t��4���E�uO^e@��h���j�Yw�wn��	H�R�ڶ/[�o;is���!�&xn	o(k�1׏��<Wbs"6���(��ֹ�m���y>ԓp��U�*�9bv\�KYs�y3�݌n�T[N�MP�t�FH�Ghs�W]��r[]��l���K���g0G9�n3��{ɍ\����jif��!TXv�8�G��SG0O4͌N��ȗb�T�
ݣ �g��o�2�;�=/����.��K��wյ'Ѽ�9T뢯�>n�n��.�P>֦���{���m�>Ruܼ���T�д���U�g�jJ�/�֠:'J�bJ:�Aq�E��&^e䅌3�TP��4����Η��,���~�9k!��EDoI��{�u2��seckDGI�Y�~���Հ�{Ύ�YNWr��9�)�� �����\�u%�2��q=t�����ɭ<��i���t��eP�̌bKt6�����7Aq6�4s\B�|ו�^�v�<�aݴ1ָ� l���o(�ʖ*�ǯ*ʣ�3�B ��.�Ә�[��tC���C���̧|�T������֣��x�c���x�3~u3U�ݖh���-�2�q��/��o�j�}���\�.l�����Q�Ш��[�)�7T�iᓷ��z&\P.���U���Y�Ǆ���N�;���[��M5�WZu�씛���җH�JW2]�e�SU��!6����G;U��d�'\Z�vv��O����t����b��f��m����Ŕs��S���������;j��n�c�ƍٺhQt�Y�o�@+�W�k+�i2G��U�$3.B���¶�^�k>����5��o��ld^�r������G3���|0��W;��o:��'�
�ze�����އX>�y����Rq�3��>\'��A�&?���yqij5�;��C�3�ȍk�����o��F'{��QI��IpU�vX�ڱ�B�^��1��Ӭ�,��*��ʁ��;�1��a �|��X4J�f](�B:�>ԣr�����F�2~ϩ}W��͜��W�U�k"3��ķ��Fd���2(���}]����Y�v�x>�-�� pU�3�މ��:�i)(�l�>'g�U8�m��̪����!i�sfmV.}�*�;��>q!�r���Mb8C�n����W�zŠ�l�|V��F�D�4��H,�.��mAb�j��Y�i�!t�d8��}-^�mh�V� :Yj�8-B{񊀬�ڝ9���WÇIK$��8���*�ǚI��d�DOw3qwe*����Y%��̒l�:�'��S#7�ͯ�����
�����Ƕ�b��ƅ���3�K�M�{=�57�;(�ӛ:J�gj/1�-M�:#���nueK�֩iQ���d�V���d��O8���Ѧɢ��Yc|�*�v�zzW���߃��O+D��UE����5x�ڇ��AB-)�ɢ��#/YuNEv"w_+�.�S���q6j�:�+R��M�5�����ŞӇ�׃�<�.c���{��8n���.s�mi7nqu�����n\+;�G_<�c�U�����<�Q�F��W7��s/6�j{�c�C�X�w&�5��
cR�b�e���^���E5�体�+�T������"�����4��X�B�����]�-Y�w#uر�%��:v�P8p��r�kL{��mxY���8�;��8�R|U�\��Z����ؼQ]Fw=��&���0a=De�%fqt�Z<ͫ�u�z��<7�$]�jZvCîiҝ|�ðb�G$�t6��=X<�̼���h�v^'�{���y�^��ލTk�yޭ��Ev��5aM �C���-��u6x�������q���@aC��ER�z����䬛��wzKy�yս�fJ+C
^��Gr���h^Ӄ֣`�E�b�<u1SY�s������Ə�'A�9g��C_�(�NzV����^�'�DfS��t-,3B�FbJ��!��9����UK7Z�Q5�$�%�%��嗳�L�	� 6)����y�F_�ަ-��I:۵��&9���`j�5S7��v�@m8��}L��۳<��v��ϔ�֑��L̨��#�H�\�!�0䫛6�o$.53��Oz���m`\���X:R�v��=6���;v�kb��*�\����%r_o1���7��,�.+���
�ڏ	��ZՖ��Ԥ��;$PW�M�յ��f��l����+^J�R%s zU3K���d��¦\Ǘ��̋R��E'R�q�M���NrA�`c��cO�T�y�o5�y}6�p�I������8^//C[��U���j]��Ȭ�Bq�O6($�K�k����i�etu�g��2U���㵔#��z'螽�e
���n��D�LN}j��kW��	/��/2U������+Wp.�Q\��WFsJ�W��V�0�������=�zvy2ɮ�xZ����}�E���J��B`${�󘎟Bq�� �v�)�w��^̶�¥zT~��"E�N�As�
 Q�qAq=t!uΉ7O[ծͭ�|��9U�Ve^�lw�[�����BF�6j��bĢo�v�΂{�ˠ輮�Sʡhcמ��%b�j,�M�j-'�'��Ay�թ�)Ì�ԃw�8�珷����I0[1��˫�'�V\��\��tJx��9h�I�Xkw�[���I��9�'e�Ń�Ջj�3��.�*) 	�
���VMp&��@�͚��D3Vlұ:�>e{&�;2��R1�r�R��;�}o��Cy&�xi�ۆn����y��y��D���72�+_h>�������Ybm.:c��k�m���<��vm�I�u�=H��7QK4%
{��9s�oSwf���O���z��'+zyj���U+�{Ië5��v��!.q"�Q�m��m;���=�AǤɻ�Y�R����-v׸7B	ȑ�U_l�x��pŮ���g%w���\Z�H�ؘ�}Ζ��!'�
���?wQYŜ�����b��a�'<��(��.\��GX-�!g��+�vV�ݑ'-�.�{\�s�M�I�v�&:m3 +"5��\��J�W����),n�u��6��V�ϳ��>t=��I�>��q���������ش575�N���f��Z!v�.���GB���>?oTG��|?��?���+����0���[|�)�8�]al=|�LSwP����Lݡ]+;�1f�.��bC���9t�%���O%��ú��0vi��R�F����"�9�����k*�'w9��N��+Rs�����L3���u"Mcn�;o�������*�Z�Q�q|w;L'�ԑ�c��-��4�n���S�Ѵ:�͊���p�J�w����sR�Xj�eu�WZ�o/�I����Z�r*$}>����%�Ge��qi�	��]N�%ݗ��f �+�RH�64K^^V]��^���nԣF��2�%X��3�\�c��ZZ̽짬cW�ύֱ�;�D�c[N�ۓ2�@���NRw����W(d���4\�V¾�\X�<�=�]OTmg9b���RJc��C8'ť�+�S��y��>�B(�R�8��K���V��kko��ðꧽٵ����.t,��6 �䱣�L�&K�P� �='.�w M5O����Y7���ꊬe]w4����g!��`��VO��1��8�.����u��9�!${{��a���lM�����Ϭ��)k�^t4o��݊s��ܺ�����J���S.�s[�!&ﳏt��V+�%��mis��u5r�u�B_7{(�4�[���<��p)�f����V[�lZ}���u�4��ٚ1a�方6-䕊������c��57sEn���ʡD*�ԇ��ή�Yt9���f�l�'2v)��b|���:v�X�^U�n��s�]T�S.�[G&�nlr��!K�w78��U���M�r��=;�M�a��l]�p�Iu1l����|�a��\�
�H' ^�	���Ħ�b��X���}CK��	��5�6�b�`v6�1�������������R�|���Ze���C��4z#x� }�I�L�֕���8��/�i��|S�fϛy�I��p���(-f��Ρ�g)f�a�ޚ����]x�o�孫'�nb����f��V�2F��Ui��ޔ��2'�1p��ܫfU�0� LZ�bC)r]jLB;%�V���9�J�8��j�)�`F+Wz���Ay�q�.D��ٌR�*�Zf���B�kz�p�d�'�5���LQ鸏��8�=�9Xf�G��g���1��̘ࡴ��/b{'0w�]�_�9�z�y3�&�0��JHY�@6S��p{Ko��>t;!��9S�sjrIVr{�V��Ol�m'3��+7-��
��D��.l�MA� �=�u�JfN�R�\U�����0=\��9;2�>&����̊�Ub*�-EE�������YE�TU�"�A����iQ�����F*�UE�E�aib�X��԰H*0�TPm���kb*��Ŋ�XY�U��AQ�#*4���`�"(��+Q���
�EQ��U`�#V�Qcʌ���DBТ�V� ��YQcmkQm��(���*��EF[Qb2#�+E����R��J��&PZ�Z�ʍ�mQU��RڡV�� ��m-�1�#"���UZ֭-�*%eX�[Q��m�(ڢK+*%B�)b��mm�-�J���֍* ��Q��U���Q��,DQe(�PR�"YFK�
#�~���%�����D���/��9�:Fe��[�n����I<ȵdi��e�eL?7�3�|�d�����ƽ]��������6�G;�4]}q��+�oq�Y�Ne\T+�={�Օ_��ꔾ˙�Cѵu7nӈ����Rb��ɏe�����1"ؘ1��=K��Q�+����#;�̪����$SWۍ��/�-q�<�P8��8՛�pn|�bb������I�����r� ���<���ܯ�:|޼{�#7{��E����n������1�iΝ<WC�=�����gy�l6���?FU���S�TgVFZKC�ԓ����b��Dt��HsEV(ƴ��	6�g~k+S�<���3���2yI1���8�)��#�/9L���}s+�F<�����ih�`�֬چ�T�x�^KT�t3��qȾ
��˝������KꌒL]ӵ�9�>�l_�����b��ǣ2�c��pl4q.�k����[�U��c�I�^V�ܣ�.P>��L�r~ �~b7�35����Q�V4�:�E��u|�T��x/��W�Si:�u�򞧪gD-�(.��9Sb��ϴ��X��u�z/��r���t������t8�n=v��/����9M���2���K�k9]�$s��E�޹�ku�
��������}l��W*���ROe��Э��bsvk�F�_<w
��%k��9�nZ�yhN��bhȘb�4���T5�k;��_�U����U�5*�i��FM뼇kഝ�#ڰ��{�oy��f���L�.yXz� �*�%�R2��wo�e����cwR}��nw��-��az��m/PX�m!#B���9A�{N]�Űx���D�� 8��:��o�����&�8>de<�TA���o=z�#�̗&�%fU��f$�b��-��br�2ON��<�x9�/ة�*�./�H�t��*�珄u�ۯa��d��g���� <4����:�k�jnB���#��rߛ<g]f4qИ�U�L����J/]�@`�F+r�'���ץHshE���H/3�����x��l���g�U�M�37Ky��3w	>���>>�����P���L����X�v(+txLa���P�YV�����@�j��Q�3!G��ʎ���3l]J�n��ek����{������X:ReI��1j�֍��xթ�A�R��O�T�ͯ%���t�	7d����䶻���Z$��׻�3٥@|g�'�7�#���������<*��=HaJ��u[������ӝY�Q]\4�K\W&����4U�:WS�t"�%_��H��L�BEl���ܪ��q�V:�T8I�n<�ڰzvy2͡e���RI�b�7�㒱K�1� yjVk����01���A�V�}��X����[
�<�����-ܧ�@Ip]�bS�3t
h�ǋ[�ˡY���޲7W��ܾ�С���8�׃��]fNg�YKc�ָ[Q]��[{�����P�O\�ۗ�-��B(%�n"iI@�B�A#ʷ�l�R�����j��Gh�sc�}�������(��?�}���F]��fU[g�o���
<����ј���*�n8�:��>�w�]��*���v�}�/
R���^�A��6�Ys�x����˕�&3��[/_�N�[9���6�9�����8{�C���w����yk�Y
�]�Rpͮ���7���Th4�uu���ʉ���)��Ry��e����4�7�o��\�["*g�p�է����;|�}'��8�V=U5���	�ȼi֕޹}�����Q"':j1��] Zw��&�6�q���z"�E2wA�m��	4GY�̥���}�3i�=1x��r�y$�#r�St�BP��J���ဩ��^E^3h��c�!�2|�E^W� ,pʚ��U���ē;��鱦����R�ݼ�Bb�mekd�>��:y�pL�/1)_���=�d���=L���>���Y��G�u��;z,.ZmV:w*�}+8���)_EףNؓ��%�]r�iW��(�1���jTu�ڬ��)w�?GC�b�+�hѹ��n����v]wH�J��&:�)Y�pe�^d�Q������Sѽ�>	>n�����gN|�{)1"�#�V��$Ӝ1/�6t�s�[*�Vr@ǎ����Y�@(�Q�P��*�Z�uu������?%"zOʯ�?M���_H*ztr6M�m-��BfHn
�ٻ9�g�D�����0�G=���!�MeB�R?C���	a��v2��q;*S�f���2�۞��>�n��q�v�����P����X���"�8C�]�x߉Ts��{a@�OPŵ~� ��_7�<{�t^��Zs�ɺ����L	߃ɵ��y6�a�s�E��^c����5��#F����@v�mG��)H���\n�h���Ë�m�36���2�W�8��*.��]eZ&{U��M�k:�z���6�V�x���]嵒�-l�̜�[Qc�s�˰�P���X�ܭ�ӡ�M�`���Q\���ϯ��������`��'����'��
-zit��9=�$���m��{�A%�ƃ��Ή�^z_�ȇ9u�ۙ���z�b�ͥ�:/ �U2��] #u�6I(7|���%�Ӭn۷�ג�*��ݡ�*���Q�ۦ�a0�V�mwe�sK0���T�k�	y�k������³�dv묆v�����R��91����7٪/��b�}mई�w"�.�Y�VUuS\9���`1�w.�[�-ޕY�o��&����gl��Z�8��
��j��Q��ӛ�Bh܋��+�h�:匈���W&�:f��Y׍Qb6,�0W	��a�De+�5eY۲�bwQ����^�����z�}:A�%i;jc�t5�|;�V	5�w��@P%tL�3�4���/�+�������|VW���糄�otՐ���>�x��	k9����)���ٵ[P��!D,	\PWX�:Ƿ����ڈ��.��p����7wy�֬���ޞ� r�S\˸q���P���Υ:� �e͎��̷�<��^2��f�S���X�uK��5���HhWܢRG(4/o�@ѥAǻ��ig�qo:����"b�T`�-�<��)W��Y�8r�X�5T��"��ß��<���to�&�먙&��V..5i�9��;8z��ht�����=�^C�g���CC�%l�v��,�s�_%�r�����vS�P����z0��7Ųc���m0/Z��}����=�R�Q�3>QÏm��P��mI(t�ĕ���jַ}OL�}K�~��uj� gW�K��j���k�#5'�O�W<�Ky���s��N�v�K�ǻ�\�>�r^0z0�����:�[8�<��J,�g�!`� 7�j����ަ���lQ���u*����c�3҆v��Ӆ.ok2�5�b��Y��U�ݻ�I��������зP����|z�T�[���a����ks�V�=K��xiu(�໤9><�-��ܓ����v-2HuQ��뮚S�C�C
��2Uռ��<�q�ŌN���ي�F�M�o��L���Wk��2�rb�z_W֠
����k|]vbF䄝+����t=�c-\��N{.������u4����x4Lk-�d����+�S��=�zz�g�r�,:�U��y�t et�R�U�炀�F"��+�4r���z��	�b/.���R�Y�i��#%��C�zy\8������A-�`qW,@�_X��h[Ѯ5�d�8m�{�r�{W/�<G;����2"�^=�fwY�w�%�zK�%�3��^ޡ�=���{�������q�6���9���L�P�Q�N�O�*o�����}�V�a�o+64��NWR����W��g!p�i�M푛�֨�ޢ�S�h����X���&6b٠���#S�1ɂR~��+�Ǧ���9k�7)������ĥ]K��7��[���YR��:��:�v��X(N����4̴&�;ɦr��n��d����M�s��r��ޑ�Tm#�;\���Yzg�Њ�� 	͚�T�U��֝���Re���s��EI���=-s��иIR'��_n�x���
�H/�]FG,Ǒm�5����Oc��XJU섟*{��]��y�Ů�g�wW_p<�v�S[�^��\�jTpmY	+�W4�D�eC�n{9.�w��ۍ�6}��	�W�i�VDk\pV������5)�V�f���+��vuT>uRbS!t�
��x��<���Dq�޳�a���*��eҎt#�m�P�g�kj�RU=�,}?"zn�yV~�-�F/�eq-���Y�HteTk�u�ת˸��y�@R�j��oO�|y���T�>�]�x1I��໣�U;ga4�5v�lO���ŽO���8+�:�Fs[�����ڻY\��5Ԃ�}Y�c�����n,��si����v�}���%`V3�u�@�2]tڗY�4�bgpqv��)rҎm�o\�q��hC	�#qu�/��o����^���p�A	�v�ssZ0�%U��X��ƫ�Q)#������$id�[�4����T��s���v���DE)������pE�����[�9�!�1y�<�f�1U_j�NwT3<����vVm��>q͸7Gu���w���o!��AzAΒy����̛��w�1o�ZI��'G��\�Fv����T�/g�QT��S+T*LĻ��+�ŝa��jGFtg2�� ��H���\,�o���lS���"�q�u��mr�Ƽ��*�C=^8{�8�P�95:�N��LF%��`��,n��Vj�y�5�'>��M˅~{����y�;���\Z�Lv�z2=��i�eE��G�<���K��w���o*����4B�54Z��O�,&�#C����<��+-a=|���ؐ���#:C�ig$���!�C�R+���E��6�	ǎ��Z�M��hO�r�A�I����^K�i���Y�C|��ZĹM��-�^q��\�p��u������7�� �i�8uɵ��أ�V�w{q|��]�W���p*�fk5|:�1p6Q�9��8c�0�!�B�ޞ�Nڅ-zn�����|᭗.Zr�����_x�Vi���i�i�lZ���x2�Ԉ����Fǩ˫^���*��o��@�o5�6�R���9w:ۮ�̶;�O^�y(u�%+Zɉ?
2*�B\ݍ�x���1[W+��B�l:��[�v��ԯ��βd��m:�h�ec�0�N��<������{jRNf&t���X�²����|�5:��q�L�U����1Z��:�at����ٛϩt���X�R�l�;�ga�v���Q>����n'eV�^Ʊ�z%,��"\��5��paՃ��e�)�TO�/�e�e��Yzr���f��(H�4�,[�C�2T{�φ����X�t�&A.e��;�w�p^u<φ��G�Er�\xQ�R6�7H�A^��Q�۝к2��G�Nǚ���Σ�*��ň����+���{Ӎ�b��]�������V�qʆ�FN�G>��f�V���X�ڲK9z�C3C5Ze:5�S��Au��1Q�ʺ�)r��X$�r�5�����JŴ���ò[Z�RK-��;:r��M�i̭Ua�*�wp����!����mB��v�Le�L���:�;��ڐi� �  7عO���|5>c1���V�wJ�%��_��Z�b�4f�<}0!M}�m��gi[��nò�d^-G5��Y5̰��͗���ռL����Z)70d��p�f�����N�ha���j�_l�ތи3�CS��lm	&> /����1r����F֖���7����8[�yL�"![��X�ǵ������p�1]M7�6���H�pv�p$ħ�Ps�n+a����[K@��grn�S�\�V+7B֠\���M�9�YiQX�I�}�&8�bG+G:��2�lN�o���&Ny[C�����_�Gc����Y��I�wq��Ø!����.R
�D�56��ߎr�tk�����=�P��B*{�y�z���u#;F��5�/�09�5���S�3����՚Mq�:���0��8�Qب��)e���-�"�vN���Ў������c���I��O�l�(����[%J�jR,-,�TPDPQQe���ER*����،UcPX��(�"���UA,���TDE�"� T*,U�+,QF�ň2��V��E��"���R,�ȱTQV(�!iU��#QE`�
�PU"����(o(cr�V�(�QAAX�2���U��Qb����)\�Y+D��((,e1��"1E�bV���Q�)Q�ģ&%FҠ�""�V(�[�p��O���ݪ��zQ� �R�L�,�,ӣ݇�u�LnG#g�j˽��<��ld�X��9�e�~N��p����Ұ�gG������T!����2�q�sP��o#�5���tǟ����.�_,w
�B�z��Qή,���k��#7�z���%1>��a�De+��� �;7e���9�6���v��ȍ~P{�5ʵ+*+��2:��;m�?Y\e����H(�ܢ'��%:�pP�q�q=jTp���]��{�M{Q��y_�)g�岕Nn�Ie���{��_��b��=�LC>u��]��ǒ7�t�^W�N�Vqq�k���$�<�A]��~�vv���� 0s<���s�"�6c3p��{���*!�̄�}����ن*��>�ۿuQ��O�tBXy�ie=喓�����-n���|��:ʽ�1Z���)����}�`��������	���1MU��:����ۚ�v�k��k�����8c��[�h�
�Ӭ[`Y��kp9�9ʹ���s�3�N/y���n�q�[y�I9NQ�
Z���r8�,�JM�m���^�}���F ���2b�WOpj��F4�D$�]-�����q7Fx��p��ߠ�����B4?,V�Oٜ;���3ò�P�J�7cV�皖�^׏!�N�Ȭ������;_���֫�Jz$��x���bsY���̨���E�i���nZq����U�4�EmQ¥^d�o(�e�=�Xe�}���&��:=��8���]�5�^d��9��@7FY;-����tڛ`E@��F��~��^�������e�u+#sjf��t��u��$�}����}�cYn��OW��8��XUq��#�9x�/�L������b���i�ڥ@t#��(�$�!����)73}'����lg��nN���>�#%��Aѡɳ�V�ۛwYs)/+f�x�����]˵۸RY���E��kb;��Ϯ����]b|��9���e�H(���qѢ)�(r[��f��2�r=W�vW��1��m�p�mWoL�k	+ o^m���=.�>���T����n�X��H��v�\M����7���pC}h0�Qn��m���î�&�V##����87��}�B^?���'Of^����F�@�Mj��&�j����o�t��<a������uz�dU�OS��fՄ�G^#�����U�ʞp�n񛛡���Y׃{�9]x=Y�>x2ܙ���m���*��Ҫ� �e�9�q6���ӽّ1�F��j�y1�r����}��8J�.�W}�)�oN���utkC��w��bw ~�rm0'�J��+��ǱҮo���KL?	����ފ�����G_�kX�'��T�#~�B��-J���w<��|���Lv�fB� k��gb�}CE�O!Bƭ�	k�uV��Z�8�������t{rTUw�:�Rs)I|�pv�v��f�_�Џ��ё����;���Q�.���fst�l��l���� x�|���R�K���:�)�saŹ
"�%g�����[�ۉG��Y;5��ޕY��gU|�ϒcu����}h2�zf���@yvy,�V��0�~R�D�̴y�O&�ۜ�^ֈ���H���������V~����\��K4z�ڪ�����d�ж!��ZN�+�f)k4n����8!�����J�5��h�����OK�{����wz7}w���S���P�^%b�X�j-$r�Úɧ��r9ȸe�r��'�uvŻ�z�[��Y�^{���;�bP��[p^>Rz>6�3�K�o\���k{Z����bIE�f:B��-��cMA��}�*��-.h���J=��� �I1uv�^V�S�C��w	�yex����g���&�ͼ��O4JS��,�ް�4�Ȍ7��w�Z���G��
ܚ��og�Y'l�Z�L cV�r�SØ-�<w��ܸ������������Ȧ�q�]-�`�ϥ���HE���V��LVJC���`O�I:S�E���}j~�Hk����%}�d�j|:3�/�T�D.�T��Ά�UWq��yR��03T�y�����^HR���W���W+˰=A��	�L~�s�'7�F=*C�W��V�m˅t��Ĺ�[]�
ɚ�{�ƴ�2������y�V�)�ژJ�r�l6�	�O���Tp����ռ���W#[�vu&#n�瘾n�ZUh�(MdËBjU�:WS��~�ݚF��c�
����>�_<�ǒ��_:���H)�n;fW�2���Ղ�ꛆz`d[�ټ\vfV��c��Iǔt�Ai;X�u��&���tkG�oJ�W���b$c���pB8(��V.'��iZ�����{t�����ԕB���3e϶�Ьw(=!Ի��E���px���M�/��915^�p���X�
���N�1����z�k]ۚ��f��Vű�x��%�yw�N�߱�m�w.��jW�3��yDZj,�\2��I���*��m崵��s�|-R��Nv��
s4��h��\�C`35�;�L�{,of��b�A]��Dw�	�ՠ�zL�6�z�������iL�گc�w��އ�s����36��t��]��T*���`XlO����ʉ������U1����k�u�.v�ax���aލ�h�g��~�����~ƽ6��_�c.�G��Fd�]�Q߇���G�{����g�����!��WZܽzs��;�~���A�$�#9�cH�S���Z��������]�FjC�Ԑ��(Je!�'�M�#M:Y��]�BX��I����{��Y�k�����P��4�T��-A���+*����Dz�K��/���>���L\�<F1�R���U��h�G�����~Sa�e�=���s�I��A%WQ�P��Q#�B�1����Y�Z;دG�L����J^JuYy�OϹ�f@fv
X��i��|E�f�2������KJ
u�;�yݽ��F0�u��:޷M�i��WHkM8���J�����0�R�?t2�. Q��J5�Ebq��-��,�ݼ��l�	�����d���}��f��ߔ"'D�����>fL�uQ:ni��������یm�V=���^+rϲ�����b)��ʱ�����q�͍��딻e%�G�����";"Ĺ���>�1��ڸe��8x����1��sH���V�z:�.I��D��F/�Px��H��U��B�D���18�<%�ΣI*5�4�a�"j	aԁ.(s�żP}��u޶���`�tE�6�E�9�e��S�,j�*ْ.����l"E-���Z�/Ԕ�Y�����HO)����������J�O�٥Z_)�8���7^?�pwyQjF�9�.=�{��}���va� Ԡ�%�
C��`�GEj�[֧��z�q���B��Ǔ���W�)��9�fE
I[+�M�b�5��U-±)�P����G�@��ͼ+�`0Ҿ�\����)!��4O,��c/_��L$	����]��#�Kmp ^����c6��V��Z�8ɜ�q�!G�٘ ���tzZY��KP�(�]��Y���ݵ-Qq%���m<�'~UW�W�ƣc|���Ӈ��n�F��%.�}��BQ:Ynx�\P�-D�.K�iiXF{-E�Y���}V}ACq�gf+j����'��O5U<�z�@G��NC4�=0gEԳA�W$X,���(�Rd�rj�.&16�W.c����.#���Pe׻k�:�ĩdAN	�A^W0N_�<��\7��Wf�0l�e^VT:�;�,���1������9�.}:�v�Q��r�ԥO	�%�D>�J���x��!]M���_�r�M#�#̫���1�ء�vo@�L[�
AJ��sr/򥨱3�b�ȼ�s���͹�3���9��X�sX���.p��58���O
1���7>d*Z�����H�{��X�wo-I�X �!��$��U����.@Q����g��Ј��GI^Y(v(�Mu�2�4�s���;��.�6YQ&�)A�����`��j��/,$���\�iJ��ٽ����g�u"_����~�}�(v)H;�4�w��we�yE���ǩ#nWpƍ7�G]ۢ_{�����N���ͽ���ދ�I�85w����ɉ��r��C���{�q�OJw��h�\�I�ɢ3�`W�8��{?����I�N1�tW���D��ZMcx!�o�<�*"����v݌��t�1ѥg��`�Ąߨ�b�չ�<�L=��Jn60o��'��*�?9�g�p�>n��x\<K��e�T�,�\��L��V�>�?b.{6���(��!���BW�]zE�Q&��3�䘎�ꂴgv�&w�N�2�c�E�Y�����=9�$X�0�2*!l���[9LE���rqQ,tS���*���3co���e�5殑�[_Y�ì0����"�_�fC>7�L]߆xsߎC略uLB�@mx�Ȣ�s���-a���쮾s�S��{M��o��P$���E�my	��"Ĺ���=o�Vё��/�zԂI�r���A"6�������Qf��7��[�4��W�ܷ���Q�5@'Iƕ�(,qDҩk���1�&�p���D��c�/�/	��5�z�]0m^Bh�~�wv�Sݻ]ڱ�t��_�$����9T5��14iL��%|�9y�t��[���f�d�N=��ɺ�u-{'K
��j�nP.3�8jXu�B�\��������鞞���*MF)���T;>Fa:&���;s=s�.��"�A��z��Ry��(���uΔX"K=)DlF���''�G]�=]sn�*����n�9$����*Ί$�5�o���T�m!.��٠Kb�^^\őf�"Ĕ�'���F�b�װ���,m�ص��VwI�xb�t�l�j�	�·�U0�Ah��Ep���é�dy����؛���Ny}ӓʹ��vyj�6q��􇒶d_=���;����+.^�
�̩V�E������<͎:�|!��O<�Jp��Ċ���a����>��e�]ѿr��A��*^�Τ�������yB,�z�ߛU�V�&3�ŝ��^�Wn��%�lJw�x����_h~�:�Y��g�~����߮\&
7�u�/���)I ,�Y g>�P��z)\cx;[�.�X����g���}k_r�wc�d��\4u���W+H��ݙ��z�?�2����{���j�0	}8���l�F�*x� \�1=���j�������52�H�p�;H.��q9����0���M��ٰ������*���a�U�{�$)���Y��U�'�����A�wA�;���ʵ�:&���S��8l���P6^Y�;Q��'�-bu;�S�*��)���x����mΗE����kh���f��t8Qׄ�H��s.T�fMV��\�թ:��;w��DG<3���Y��.�%�J"NVl�A�k+��0�ƳAY�=�3��a~�*0�Lί>:VX���W�	SL�+͠�V�ރ��8s[�9!��v��Q�ΰ��s:R»7�c�6�֐��q�3�EK�r睒kSS����Cfd�B٘��aܮ�w6�4LSrF�������A�����S�cJȔ���޹�G.��j�����<Y�/9X�Rcw�V)c%+����uH5�+:>��oe�p��?�h�W��L�����p:J��:��������!$fC:&:Er�s)��X5Ů<Kr�Z���<��rȲ����q��â`��K���9���
�x-�Ÿ����x�$��	�q,ôJ�v�5�g=�zv�O"ZU}&GЩ��2
��>�wl�>��������YT{z�ˆ���o���Ͱ�W�׃x�u�h���l��X��q�ᑘ�"cq��h�P��ׂ.T�|9��n� �"�ግ;M\�pRSp�}^kh,�:�q��2B%�Z˾#�&��Ky\%io��ޭ�a��xb�4b�wv_3�i���w(��zG�Ǧ>��VY�MӦ��j����I�W�����Y:�\�d�ȅ��u]pč��T��o~-ͫd��]\�fP��;�;��X�w]����q3�L�bR�]�"�Y7��f��S��l��o]*�:��v��������uQZl��1-xv,xCuM�t�v_^����h�o�6�����##���;"�m2;��jt�i"�XҴ����L�x���`�[ۆ%t8a���\r�3^XH"�@�d�M9�!u�&��1�L��_J]ò��;��,e$��Gw����.���To\vʊ���Yd\�
o�<Zz:�{^�º�G��+mb=��.�XgZ� $�jK����K11sa�I}�V���9RD0s���6m�ъ%^�~�;���3B��톼ςR��L͖c✎���hEaľ��XVc����,�ȡ�ѥV���.ud�n�����1ꬩZ"�[AKAU[�b�IR$Q����Ȉ�*�E�����E��J�"�"&26�J"� �Ad1�X�2�d1dUX�AVe�q*�(��X",TUE��P*���!U��(**�QeE
ª�S-�E���m+Y�Z��f�9J�E�AW.R����8�V
�+��cJATm�ETb�,��(�Ke(�cEX�T1�DV
�b�UV#R�I�2 �I���B�y�'e�gS1�&ʺ���Yˊnl'�Y�]���k�kص�p��HԄ̗&V�xPޔ��
^  <7���4�AU#��t �����P'I7>3���B=5:Ut��i���Ⱦj@Ų�F���5̢��#Y"BOh���4�t�f��E������^�<�H7X��i��D��]��f�+���g��e@X/)�S�v`)n7�Oe��q�He��0J�b��/�>.�hK���:�� N֐��u=�u)�:��5�/b��g�u���'�)rrK,�;�rz�vN<|5o�lA�n=}�"�,���'����R'a×aO��t�&��φ�՗�˺/@�޴E@��>X�Jܳ��qF�N��9��yWL�3I�j.����<\����Y`1����dϻG���+nYӇ����wF�Y� �}����#���\��{���*�����#n}��_.yS�3��������2�+%[��$'$Ϻ�	U�Q&�s!����`��3�(�PK�N�3�Ru�os���;.-������%^D�� �i�l�ECtwt⢗-.���������|�Q?]$.�Zǃ"�kM !�E�͇���k�ٹ��f���΢.��zb����*Q}o�B0�.���� xx���rV��Sj<�fH��'=��]x������4:Ù鲼�o�����t�X�z�m�e��;�G��ɂ���8<���ٵe�F�5�9.�*�8��PT<b�|݉�Z���`�GEj��Y,�_N��q�M��Lt�Us�䶜Ɯ�fER��r��ؘ�L��}5
��B�8�0��Z]3�Qd�
�Y��=�:TJ��%.�au(B�&�6
-�/nc��t��4�s�i�S�⎗Y,�>�>�Ǖ��P�"B�Ւ��n�Ω+u�9��C��6@�7���)�s��ĄY��l5J� �ʆ�}���Vv���Z�&�f�~���O��DPE�ϲ.u�ʖD	�<S�:֕��gb(<��7��J "8����Ys�hl��&=z��t�@��΍�l����v��%>Ó�S�`:�ZH
��K+�lWkP7ѥ�J9C��	�C�p����=fF`K�-v �K7�������L�m(5�gy�W.V�_��[��Y��y�N�
k�#���R�3���F����5f�|�r��[��|$y�S�zw%L�T6,��@�9gc��%Y�Ek�z������xen�����n�=���	W*�:�De��i%�Q�N �S������N�b���t�	�ꉍ�Z)׈U�$6��5}���{�D��F��׸��9�{�Ŝ�C�v∌�I�e*g�'|��G��S
1pDk�(��]����^�=���W�G��ãxT3:��C�%���l�K4�2��"��VYk	�����tMA�{E�\��e�*�a�P�}1U� `�Ǆ�އ�1��[�=�!�����9�I�sgt	Wpjrh��������1"��*|�XbbI��16���3��<Ȕ��������8}�:h�yd���7O_����$�ްyI�R�{�T=M������mAK�`i��VƵ�O��I�+����aP�z�i��PY��q�����=g-�!�?y	'��(���?> bmP�|�~������'��R

GÛ���=����d�'����H.ٴ=3h��R�՘�IY++-�9���]w�y�o��I��ى9ް4�Y>N8��J�����!�m�:<�l�0���f�m
��>ʧ*ISG���=�`T�Xbͳ'-� A�"�o���s��>I�K���Ag2����
ԝr� ��R|���$�'�=wC��t�P���"���1']��%A�~�2q���T����'I6�A�q��d�|�U���}��?�=y���n���yŎ�3�ӁGt�e��n�˴*ۻ,�Y��u�m��./t���㾃���|�N�\F��?�Z��@�-e�'��Y�Y��R�o�FH����z��M	����Q�e]�p��FcM�R�W�����h�����#�|��q��&G�>��A�hJ�XWhbi��>J��W�N=���7�S���C��k������bC�C���<�m�� _���~�Q�[�}i>@G��T��:zM�L1'�s���;�)1��P���DR&�3"��W��K�&Ь���OP1���' qY���i�D|h���}sי7�6�~J���yI��=�#��fӯ)�v��P:�� T�����2��6�C��* �{�y4��J��γI;B���:m�Ì*w�冒m
�ġ&g~�w�uy�fo���o�<�HORo�0�t���!�>@ղm���4}��CG���L`(}��N��k�I�N���&�a���ݒJO��k������Fi~d�*2�d�+'I��%N�bO����٦t�P����1��Y6�~ÈJ�YϹ��t�d���Z�i$��;��u��AH/~u���,����;T}[�Qd"<	���V���b�]�ćv�'���ư8�a�VM������&3�1'�f�!��!�����F}��)��� ��G����w��OOo�L���GW.����u��M!Y�%��!�J��k���)'�����6�ĩ�
��=�*Axϧ�`q;`q��d��+��t4��@�߯%��i�M��z�o;*>�A�:IY9;�
�&!Y�M��1���*u�{����{a��Ch{�4��<q�{<���1S�l��@����Xr��{LC�����z{�7y��o�oy`v�14�H)�=�Ϟ�c����b���o�19�J��P�z�D�L��k��O����<;�I�Vt�S��m&�Vx�8���<	�����Ó-�u��\~�?'�*�&�����ÖLCĕ�����A@ѿ0Ӵ��M$�_5�Ob�-"����>�����Z�4��+&�S��&�'��eiS���/U��t?b�aRVR�?�okT[��˖���ء�ت���o�����>�S�K��ʱt�ኞG�e�N]NN�ۘ�v��f,�;*Lb��r���Þ���[�L��o$Iˤ����y�U_B��{�ۻ���hm ��:f!�+��oX
E"�������݇I=B�l:�5�B��J�_0�O\� ����I��Βw�`i<@ �q�	��H�$x_o��onf}���rbN���b
J��Y�=a����M!R
h��l�i+!�>B��g��1�l�8��o~�t��+;9�6ä�
�ϙ`� �q�G�wW��2���5��:�����c�y�@S�
΋�=C:�*N��b��,���H(,8׮X|�$�w�ޘq�d�{f (���t���J��L�%d��>Tt���/w�ZW�
�|�dQz�d�Y�%-�bJϜf}�I��r�3I�J����*q��{�1�W�t��״���O�c���&�56�yI�S��7~�jb��Ů�u�:�G�D𽑨t��Y;9�8􂘅d�s cSl�Ne��Aa��u
�IP+�)�S̓�i$�>MY�B��k����m/^_=s}_8y����7��3��{� ��Y����!ߴ��@�4w�N�����3�i4��S�>�4��ҡךȳI6�|�'I*!�fI�V/� ��Ǽ�� A����O��+W��>�F�Y=ea�p�)��I���0�|�Y��1X|�CR(q�<�S�`)�
���6�z�*��&��M�'y�J� �����]$�����Hb��6����7�p��g��~C�I�
(t�:�4��P8�{�������Z2���La���N2�y�Hq%IY��8�PR,�}�q�&�*T>�$����W�T�Mu�Qy��:~R��H��}�I맴���XL{I���N��������q �:����`m�=C� �����2,j|�0΍a8��7�q���+fq�0�}N��V<��� <H��u"���T<I[�gh$�
�N�����B���gi1�VSˈ)�'>�*m���i�Ad���Lw��AAC�S�}�Y���y�^��7>o/Te���%���!~������[Gkp4B��AI�<M+&�H��g����w��]��ez[4��G�Y9�jW=�7#��5	�:��[�N�f��+��p�9�V�5��X�`�7{��h)�  < �/������}x)���m�$�VN��&�1���K���R|�g���H�m��g�']�1&�Ӻi��*q�C�6�Hz�N:N��i"�P��Ε������~C��&��K�h���}$	�G��1
�̡�r�N�
5|Î$�lćSkF2c�>|C�[�4���m�`q��1�Jɶ_��<f���&3��6��8��g>���^�Q�3��޹��g�|p=C��%N^���%AH�NRv�'�*q&$�T��oIa�{Ν�c㤂���*E�;}M!����b��ǳ��QH)^��1��S����O����9�}��rM���!Xp��f���6��i�N!R�a�T��$ӈ)�{C:eCht{M?;@ĚB�o�6��R����4���Q퉐 �H�#�w�v�Ψ���k�ݽ��R
bN��:zH(uil��L��H((m=�Y&�R
w���J�a�
ɶV.��1��Rz�w�q�E��Vo�q���P$�d$�v�߫��j{#��8�Q��4��<��$�x��gZ�PR(k<��:V�a�՚f�����ACԟe5<�i�AAu��I�c'S�M�Ï�f�a@Qgo\��z��x��뷩(?Y�������|Ȳ�J��ߜæLeO����oY�l��g:ԝ!�J��k'�L풠�頻������I�6��a�R@G��QG�gM ~��.u�#Z��\�v�AH�$��4�<�bm�a�/�LR&���ިm4�0=o����
t�g[����6����x�@�T�0�T������0G�����Ssz�ѿ�n�����n�1'��U��^R�ݛI�m'���ĕ"�������AN w�։�c�:߸�f��i�g5������S7���+*A�fa�:IP����y޽��<���}�f��l�]�;���I��i�jE���_P�'�P1�M�Xz§��C�*0��OL
��M�q�f+O�����ɳ�ɤ���y�뿎fo�Q ��'~����=������4'T�)�rcGD�i��{α�Ƈ	u3�V}����y<(���Ĵ����P��=p�ܮ�f�u��4f��x�W�)�VI�{fnS۝K����9i�L^�3���ͫV����BB�7�׻���=�?+R
~)�4ԛx�aٖ�2m�|O'�� �(��t����ua��)*M�f2zʟ&��TRm
��W��&!ĕn�fޙ�J���y�m�_46�k�$��� �����|L�@'�T�}纓״��<��{d��N�,���N�S��)��t}Cצ)����T=N!�����ALB��8�0+S��=z�]�>:�<�߯�}~5����5�°�V�3��AH��N2��]�4��6�ݚg�����J�$��T�TAH�l״S�I8ã���}fH�=�A���ǜ3{[Oz>�'�6��!�i��'��
��&ӦJʁѼ�N0�bJ�u>� i��Vu�k]���'w��1��"ɴ﫦���P1��������M!��4�k�쏦�ev�w�.,��ÇW��V�u�L�8�nýXi ��4_ro�� ��a�I��1��ɉ�O�a��t�I�[օ�cm|�NҠ�^��|�[����}��｜g��eM&����'��N�]3�J�W��i��8�Pz��c%eN0�11����sI�Lq �A���4�'�n�oV��Q��]BH�$2 ��F鯪u6/�8o��	�lR95dިv�Cwl�Xj
bk�i���
�^^��$��VaP���i�Z��7q"�YS�)��q�!�� ��>�(��g���D��}ݰ�u?"�Vt�׼�PR)�<�z�=��<��I<gN u�1 �g�q408Ԃ�Z�ҲVT�!SL6�IS~�I�l���;IX�3}�9�����k������xi�H�����:a�*y�&��LB��Ng���J�ƻ�x����,�*g��`ui�eghg)�hH(x����Z�#�I �`�"ϤKP��n�9�]�e�!�v���;v��
NM���C�bG���4�t��氞3�OS�����&!Y=5�M3�J��w:�I�x�8�S�)�OYS�u=��@G�����\��dbJw~<nG����[��;,�L�3u[�k]��&�m`|�XV�pN��Y�)n�#�+w2��#�e]�²�_\�t�Y�3�-+ٱ�Q!P�<
���Z�):�V�N���C�G�ut��:�
�^r�.�����7��CT��砍>�"��+�'�N���R.��)��v�Sě�<���)�v�'�c7��x���PS��Z�;e`w5��|��bM�_�a��{��Ӌ�Z�/;�s����|� �>�H�z�������1;���6�waX(m%g�}O{��7��6���S���IR|Μa��Ă���!�>L�O�w�C6�u:��CiY++;d���p�XH,�N8��J���l>CƤP��f�q�O>��4�hV!�U8�P�J��Xx��L
���2C�a$z�>��g��S�w��ZϼHD�ghg5�� ����:���I��� ��R|���$�'�=���4�P���>�ĝwgΐ8����2q���T�ô�$���}�ֽ�����3�:f3*���&�c=q��w�ցH�m�:��@bT
�F]����>J��W�N=�߸CR/ɣ�>�i6�}P�)=q� p$�����&"^�c�r�K��^����4�d��'�Y�I�4�|�� ���Nw��`|�>�a�&�3"��W��Rm
ϙ/�����J�'F�z�� �$�v��}K1j?#�f��?kP4��c��LH.��u�8��8���AB�d�����4�a�b��T*Ad�z�S�.�Vڸ��+8Ԋyl6�Ì*w��m�<ߚ�_s�l�<��>I��Iû4� T>I����8����j�E3l�C����eg����|�*Aw�I��+Y龲M ���:�׺��'��� I�Ѿ߲7Ty�p|9&�B�a�p>��%A坙bɶVN�P��*t�m
�{a�i�2T8�7a��f�g�j� �Y6˩�����Vt}̜C��'�0��S�D��}�յ����{��g>��"�k{�<}O
m��&������Hwhbm�O/L��ƫ�+&�P��:LgbN;f$C��!�����Y�H��Xmݯ�;��P��U����`fz�1	ڴv�X4;�٣��x��Tݕ�Xa3&:݄�`��ⱂ胓���e��:z�e,Gj��0V����v�fn��i2T=�N�����ڊ��&gj��WF�P����� Jms��o��A� I�Ǐ�Lz�� V|���!�IY٭{�x�� ���P�퇉�H�Sh&3u偉�4y����AACiO�J�#����I�1Pp�wz���?}����AC����V/�+'>�q&!Y�Rs3$�V����\��;I�+���
���uM!�{`^��Ċg��N��bm���P��xA ;�N۷_|>r�yS���$�,
�`(,:jO]�I4������08�PP���'2�\@�*��L�ed��y4�'i1'�y;�I�Vt�S�鴚IY���돹F�^T���O݇�
 <O��끤��@���4��|�;��b$��*m�Ă���ߘi�O]&����P:�'�1C���R��S[�A���. ����eg=����uַ~����z���|�:f�c{~CI�ӣ�4��Vo^kH��Y�P�Ci+�l�$�
Ͱ����
��+��$��R:���E1����� I@G����^M}O㗯�D$�)�}��;N�j$�(m+'Yf$������HTtw�6���Ŕ~<��Kj`�ܪB!�8��M,�A�}�e.Ua�:Xt�iu�����+�OcO�uWq���v:��o-r��z��=<G.�|�a��i;����b��+�okk�]��<�4�_Sd��m������<_�K�Yق�Xr�P��L���Ά[�!4�f&iE3<��h-v�Õ�!�y͍�d_U
J[�G#�#C$HT�&�$�63Y�0{j�M厸�R����|��-�Ɩj�g&O���76�mv\��	Lr%��Q���2u-���qZ�@x�:�^m�Q#Y4�����֏G-���81hz��ӝR���Ybwj?84+���Ї���� 78ާT�r8~#����
�e8މ��d���\��:c�j�5�T��:Z���ʠ'��{�s"QT6C,�8z���f2z5C>�n����fg1��i�u����B,NnM�MFN{!��H���=�EbqB\��n�T�A����5�wOO	�K�D	s(�"s-��V��75��4�2=�dNÇ-%<�}U=	_ws��>�	3d�1Lex�d�zg*���41N�M{'�]t�]���p���� ;�x\�0# �dϺ��;��Q�������w�ȵY���,(ù�ze_���J��D�J2}��Ц`�8�i�W�
sf#]K�$㱴ȑ�I�(lQ[�N�U�yS�53�9C��%�n4;��Jq{bNU
<sj<��fH��N�BΛ<i�pB-�e��[|�;��a�ݩ>�`�r�c�o�*�V|>�0���,��}d}��f��ި�R]c<k&��kf�{ʏU��·%�.�C�t:[H�
^ǁ�.�b�2�x�l��"�l�{/�?^�ʠz0Z&p���U��"5����]��S�\���AX�hE�wh�)E٭��Zeݮ�s�-ÓcF��QV���k/k��x�����s���X��rX��tV��e�)�%��)�֎@�f7�)o�YXkif.�@h��������8e4��j�UhR����+�^bȏ k ��Q�̭��s&]�ms0fU�t��v�.�	��]�] �Rί3V;%���n:k=�x��0�O����;�&PՔ�^��t����m�na�'�IV%�� �����Y82���6T�J�����A�f�ըdv�+��mG�� YyҠ�8wHe�٤8�]����d��v[�42�������<�K�X�5t_=���q�ǉ�����Ș
��V���:|*�x��or[��b�Hܬ��!�Y�Z�K��w� <�4�@Z-j��yNQ�vy9Z6�_]b��In�j�SZ$��ӭ�� &y�_gv���H-����]wM�5S�(aO^m7���E��"�I��1�l���
����xk�&Q���\��H-������)�ʴ��sM��Ѷ ѽs���'V���(����傧!��n.2��:xft������Ԋ8�s�o���f3kfH7�-t������o%\���ݞ��ܝ�ȥf�Va����Kq^�.-���!0wn��Q[��Hȇ+k���GD��:���Ms���*����Ǒ�H�6»:��!&���B�%��"��p=�4ԝݵ�#[�+=F\xGTA�S_֜��஛5�\W۰����F쌊���-�i�5nu`��tq�Y�}Q̍��3���H`<ٽ.�j3xq/t�>c#�&��Dk��Ź�

�:��m���8o��SQ��[Ch0O�]��\��ʙ�Jpk��1�ѣ�So���\Yv�:%ۛjӺY�"�pgT�<�E�J�|T�{ϛ�t�N/���V{>��Ӎ)�p$����@�s5��ީ�������M�a3�V=�(e��"��͝yt,H�֯�(���f�yg{#y1���>}\Ae�h�#��U��K8��D�p<M���j],rY�o�Lw�*k�9���s��6��J��e)J^�%r|Y��
}�]�ԃ��bvJ�T�X!P����o���EV�����Q�9��.�xk�ز��8Z�I;��,կ�uc�eZ�^�8)�qm���o5��s�?QSY������)b	[TY��q*ċ���ZԊ2� �R[�IX)*Dj-aX�
�H��AB`�e@��b��ł��)�*��TF�Y"������Y�$̤0AT�Q��RV,(�`Q�(�"�m+Y��X�)����*� "�*�DPS+26�� ��"�� �Y�1�Qq�YRe�e���s2B��T�!Y1*�j�Hc& �PP�`TUE`.[��11Tj��ge��{�[fR�͹gu�>�Z�B�T*�s}�o�rge���I�+c9��9@��sof��UUUU�/y�߾R8&f�#o����Q�v"ZபЭ� �/��t�-Gz=�����w�[,dyb�Q|��-�1�BfE
I�]�E���Z���dʓw}��ij�q�bԼ����!'aډ
 P[0��r�����y4PWu
��=J���X�d:�gj��8ގ.���>�>�Ǖ�vaB��UTˬwzu��e~�SY����EDI������7����e8���B,Ⱥ�j�[�k�b��.0D�G�ڞ����VD��,ݰ����>י�u�����1g��\�(�n-�Y���V��&��At���Y�x��:�e��l��ǯC�뮣�}�
�ϛ�K�(Z�=�>�=�p�OLaqQ#�*l�E�t��;��7d�;�}.��O���(�u3���Zhg0)�"6��}�R�*|��Y�_P�Yy��C�'�g.G�(���{�,�0����*d��+ˌ�\����c�{9e]��Np^�J7n�ȹI����z�pg`e۠Uw%�
,lt�v/�%�u5�ۙl�ˌ�#�S)#r�٬��"4wN��	�։�q��Lj3�J�7\t�5)�;�ds�:�S�!s��Ƃ��u2eM]����x :��m&k# q����sj,�DFC$�gJ'���x���Q��F���t�K�"��g�0Y��_�o����ߋ#J$�إ`#�[0���}��&��dS�E��dXrփR��p�}>�V��j���κR����jE���l�P�G��YH[�Ю�����t�:X��M+>�i�rX�����u�.�P:S��(�c,)��hΨ�YH��h����_��9��V�b�����na��G��8{�rf�r����Y�$�1v��[Oy��D�X4�"�z(\�����dn)g;#�ܼx_e֌׀��Ǩ�k8�Δ��1��K�_P�����g���V�����ll��]��5�����H��(��
g&u��#^/���5�}��W�i]S��'��6�-���������f�,p~�~G���B��h|�^�%�G��"�N�����sev2;�q⭦հ��ފT<���oQf��i�lN˻	e���w�����e���Ir���T�taج튄�EF�E<��uV�j�B��δ��
fm񚬋�@R[[�呵{`�]LJIgB��{���ub��s�MϾ���\􍈥�c�m@$��-E�#�j�!��<(��b56�c�7�}� ৾3�2�)�n`5�;A+dW�8�_5Z�\�e@gyf���;�gP$����P�7;&��4]�)��|�NI�su=�y�[���X��[��?|��Ue�ֳ	�����â!�P�(��u,mQ�P���Vz()�������c�;���T^9��DDN@y.���L)/K�GUJ}��!2(��i�ZhDh|�$^��(:}�H�!Z��/ٕ��N��F$�\qib��@��DߒW{���,hm�ʋ��e��$<f�v��'�,*-��d�,�=R�X
0�zG�d���jv����+��4W�I�E��GK3�/���<32QK<�L߽���Y�[\�y�_��>�ƒ�I���~_�<���f�hR����-���}��{�c���<w<BN��'���H�ȍ����q̬�b�ۛ[޵1�Tn.8��-w��7:6�Vד�7�#R��VJìɫ���H䙎�u�v��:�ÃN�(��+r:L�DGTvV!*��j]X�xx ����{�&��ha_���t��V(iB3�h\ϑ|�,R����D<�bO<�;��g���b}�qy��!����ݯ�&���tY��{#;7`�3;nu�̷�ի����س>\��t �;0R�r�W�4�z<+:Ym��F%��d�_s
��F]N�����/���dM�P���2���{d�6.oT±�9ϔp�F�(�~�3a��';�*<��3>�J��̭e�)\�����k�w�*g�)l\G�(D�u�f����R�PR�蠡�J��̔�.���zb���d�\�O�fN�dX�g�u���@��*.k�GG�o�ި��
K��	�p���<n'2�/j�ȳj����)*V�B���QMn���Q��d�L�):��0E�\xhic��p�0xo��^�k���M�~�^���Ϳ��D��7�%�Ĩ���
=Y�{М�e �2$3ow� 9'[��[����٦��|��u�T�M�z��hV�ܺ��"�Km`�2�pѓU	�	R��nl�&D\a,���i�]���1��uGg	H�f#�iMY{��=1�]�Z����囕�Ї����+85����;oJ1Cg�b^L��u��Tgs�j��S�Jg��X�%�}ݦ��ڂ�����n8ݹo�&ލ��������$��B֖��7�uG�̦�F�f3���;�B	��C�4-O��"�(��L�+�[���!�a�.G��hw��a�X�^/���٥U���8��m�o��=�4�S0A��e�7yQZ+u���e
����U������ۛ��$[7�7����\��9m)�8fE
I[+�M�Q&��+wsq�Ξyt�Q�	G8�j^l�q�I�z�jQ&x<�����)���M��]Q,���ۆB:9��X(�y�>�>�Ǒ=�Uk��jn��y��gN@j�u�@�|Oi���RމOʙ��OM�E���M�S����P���ҹ"�eC"IEf�¦�M��VW�B.����θ��mk��.Зæ��\t��k�;8�+4�q�7u��l�bڕ�4�w���Y]a(��YCb]������ttL�K!�ዋ���!���r�����3��BR�0
=���0�\re�\��U��V�[�Ӄ5�D�'��A�JI3�t��C=y7P�,���&=}Lt��2�8�V��qC���W�5)�s�K�\kĀ�ׯD��X�a�])��f���p�Y��n��m䳔������N�a�#9�N��f}����[%o_�Z�qH?T�n�to<�\pS��e�"�$��L�)A-D������vOK
�[n��{��}�������q���tX�DNJ$ϲ�3}��|M�82�Y����A�3gס����P�o��C�:Y6&v)A�33�afa���j���΄&�*�>�USYPs.�Y-h:R�*���@���*���UV�c�����`�7p��:+���U��D�p��]!bc�6|ȷ	��o���
5Q�,��íM�R��e�H}�FuE��D_��Y����s�Ws�8pJ���s����3�P��M���J*�\�m��(������ƽ��}W�[�X�����)X'�1�+*ڵ;I���I�߽�[G/�.���=5���֍�w��)9G�7�0����Vv�ҫ�h�����'>������n�C��E]���3� ��Z�j����\�dTo�B�Cp��ȬR�s�s� 2�5@�R�y���N�Uj�ȍ��J���UD��g�H]ohW�l_C!�|T�v�l�Jy&:ɲ�\| <H��GN�?p�� /��a��^�C�WT��E�=z<�w����R��Yne�.=�nD�r"��ͬ���Cwl��j�	�U�^~�ĤC��Վٵ �s��"	W"O3�1]q�\j�E�e�w�l2�)�o����J�8�iT�7��k����w�mW�;��\1B�2yxW��b�y�Ǡy�}/���N���K�n%��e�J�;j��/sp=9&��:H�DIFGLÇjCeب槡��u/��U�	���h�k�NI>A�(8Q'n��l��+Q��n�Zȴ}d�L�Q!�Z<+���8�4;���]�׈�NL�B?n����ҵ��kZ�ޱՑ�{ۚ	N�������X���J[.f½P�
�kU	�syV�}M^��U�ds{5'K�1G��T���M܋bTF`{��u��J/3X	��Ș��w�aK���W����ڭraS�:��UU���7��A>�������ܱ�a�w�ɶ~ç;qQ��x��99cכ(�#�������Z�J�o��5<j��l�T7��.c:��="�6*g:/�CfM�O�fJ)b�*���cؑ�-!��\��Eȯѝ{C{<s��G�@��s����cjH�{<Y����2MH34��m6��J��@;��}�b�V(iBS9��K���u���~�d=H���N%��V{���x�`)���y���ikq�Φ �.��t7oU�G�;.\�'+����e�4x.t���U��(��������Vث�X�]N�l#��N�]/zE��oa�>��	Cs(����˻Zyv�먧���ē"v8��C.�f�4+%�9މQ��^f���k�3x�qET�kƅ����v���;�8G�qy��#LB�c��OE�!]/-V�]���{Tv�6��2�F�j��+A2��Bˡ_��8�g��C��5J݋��$g<�T5��PZ��$_*z���4�Z�3�����s:�SY�X��B���c7R#�B��eR���{\�je�U|�T��x�����ɿI�ɲ���G�s\�.��РFK\*++1�� a����Q42��Y�b'2їӅ/
�����C��DV��wb���Req����;aϑ�`��TM�`�4#Ʀv���;�E�oׄd�d�l�{��s��+�}���^�O�q\�U�<o�v͉S�:Y���o��8�eb5:���N\_��1^�d��3�۔OA)@;���ʠ�Bbs���\2[��w`�^�C�UZ!âNTé��/
��@-j�/. ������}�p_|��"�~d�W@��?��Qf���'9}α!Q�Q:Q
ee�S!-jcR���b�����s��*���*��X�����&0�|�ݾ �+��o��}�GZa�/�|�޹=�-34[��0��{t�6���[�K���&Y��/iD�^���>�r�M��ΛP����#�Ҙҙ4���O�l��=��zN��1��o)�WN���顙ӓ>3&�O	�������|+J73�r����$���G\A�Cr��q¥DV��������g$��3 �jk�+�	[�Ĵ4j�y�$;k���^;q�I������t;i�wG�'����)�p�<dZ��8��!'aډ
 Rل�9*�<�[���I�y�g_�gQ ��ll"\��,�k��z,���K8�h�������c�c��8|FT���u�[c����U���^��j';��(,��'ڭ��p�U<kUu��,�ȒQY� ��>|�mK��[���Z��g�2�[Z�d�1;<DjI��ҒL�*�+��e�g�+����q���RR�caOq�K�����L.sb\�RtM( ����(���i�Ŋ��Y������a�Q�s�]����h�#�Dt28b�F�Aۅ�R�9�Q������w��׊���Z�Y�b
ྜ�%k���E
L�)A.T��eYy((��<��{ݹ4�9�#�O%��5���H�#rQ&r�3}�RH�e=��U�b�����RW�r�Fž3��*���#7,u@���,�a]��Cz2g���^�f�h2F�W�C��� �Y���	yI��Kyt�tb�\k{�u�PhGI���N����n'�n�kN�Էc��O�|og���h��/=~�(�b�5���a6�E+N���m�c���qk@�B"]�=�nM�]G{����*,��Z�����koV)'
�q�ںG4'KF��š�Ⱥ�̝��dM޽�{���[ ɍ �IO��&�u��D����sd�M1���sq)��i�X̑n��*s��D�z�U�o�T���`^�B}��(�9э��*oq]]�� ��Z�?h�x�h�s4��D�+�:hC��j��{$ɠx�3l$�ܖ ��U���B����f�(^K�x����u��HA�;.�դ6賚*�j�N1��]��p* ��q�1�Z�-W]���Y�K2
ˢ���y,,�uwJ�j�-��4쟢l+��V�6�se�����6�"�o���S4�5�`�ӓ� ��7�C����{7 )���|�p"���ܥi��B���Cz��w�����n�R�%�'yD�Wu��x f�z��դf]r�33l|�\] �\�'7,|5��ٮ̴�$�յK����B��Kt'v����9Nm+Wz��sJ���IՊ&.oQML��&�D�q{��h�2�쬲7^� �!U��2�����+�wvd76l�۵�2��+7����&�3$"U�]h�q�����M�E%0��k/�6�jq�KH5�5��,�Uw�H���g��1�c�sЕ�����Ab�(a7)�����B����7���<j�v�Rf�q:]����֒/s0y�EA�����dPbV�x��эJ��ݚ�׀vԻ����ٛۚufYQu��i�q�LE�7�iǂ���X��ؒ:���C\!��M=�������t�p@�WM�#U�IT���&�ʷ����V���n����и�͠h�*ƛ9E}9Ey��r�ɺ�]�Y��\e�3��ǧ �{֎U(i���2f��['`�V�M�C�2��N*;%���֏-�K{s;MJ9mW"	��s&=���7�^��K�)'׬h�]]Y�1�=�U��\���l���c9S�V�,&E��	1�.]�g��ڋ���yk<�ST�r�]�o7l���Օ�
��f�J!����l�FIsf�?6;E�[8tؼ��S�ֲ���ثwjfF�o�|�@>�<��T���"ij�%̠�3(T����b��̡��P+!Y�
LAf$HV,%J�E�\�bE&8�eB�RbJ�H&Y�0�)QI1��HQ)"�H�
c"Ŷ�I�,�RAk
��J�ą�B�&2J�eH�1-��B�P�f8�1��q�"�ő`c%Jѕ&Zcj̨�m�,R�La��r�6���ciU��Y�@Ī��Į[* ��(��++��`�SV���d
J� (�T�
��{��5�{��۠��l�-���+	�#�<se6v��$D���+鼺�gwe,QN�*�:������n$�ʮ���\�2�
��̊u�E���,?�kA�n
�ϰӇ@���oq�/4j���E�YyF�M�
dlEYRB6�a�]!�&;��t��������lM�����ٓu����S�
<��X��{��\���cj�؞x�8��LDmB.������E(��QD"��l�JCR�:�9��r��u�h9��� �&�F�P����g�t2-C7��;�
�e���}�&ҩ�����b�e�5�8J�]#!U[�Y!0뼶��@1O=~��Dl�����8�j��z�Lts1�t�IQ'J:ܡ���&m��+D�S�U����o?T��Q��C"�4�S�Xc�d\��@s�_���=Σj�M�o-ÜQǒ�{���r/��lE�c�m@$�p�A!lk�U!�M>�]]�)�HI�*l�(,ޘF�e�AN��b`5 �N�J���7-�7֜���#��#Ք1��םV�Ĉ���\��i������Wb8)u��w�D���|F[�v��|Q�W� �A�y��vSY���d��),y�.�Yk+i�N���j9y��¯���y6����Zs'��H�9{]
{>��o<�k��i�ܮG�Y�4!U9p�
��g��=4]��#ȿnD�4!R��i\���U��b\��Lm�/sp-�ȁf�;�Y�D�z"3��e�t735f${P81���GUW`$cҼ0��%����2�k
��Y��;�B�y8Y�&�T8����3�3�ؗ���ιոH��Z$'�8���?KЩ b㉕T��pM�c�P�I\l[�/�E>XЕ�!R�_�S���7�5ǽ�,����5�0`�?_�k�dsɜ�R\z�ʃW<���^آ���+TǄi_���]��g껵ú��o�Y�-�f�|1'�I�ѕ�r�r�`�G�{'��(�f�ƅN5����D�=�:EC�yiٽ'��+�Wۤ��4������ʹ�n�7���{���Ι��V���:��֟�c�r�̆|���/��dׄ(�I�M��̮���}\�oԮ*Yh�2���
F�	�#\��lP+j���E'���":zk�����5嶳U�ݸ7K�B�C%�'�7���m�=�2��	{��j��tsnf_�,��7�(?{���$å�l�j�|=鱐��h�s��B
��(��P��$�蛹Z�Yz�ܜ^îYO�3�V��!��"�d4���r:B<��2{�j��!�c}:���-oQ,DIOF�l���F�Y,��*<��y�9�Xc�.{��gZ��Y�:���':+�[�O����U��ōd��2R`mi�N�%鹽�6�,��.����ir�,ܛ�����(���dQ%lU��5mu��^�p(��G��I��|*���QWs����_�C��g�>V��2F���N���u�b�N��ǎ�����V��WȊ���:��.1�r��*&��I�#��J���/�����"|��W%��_��ډ;f._C�=��op8lh�,U�\7���^c~<���_*�O*�gqd�<��>j"�ճ���d����qƜ	9�RN=�F�d�v(�c��餍�>����k�9V���l}����nˇ!4l���
��CE��ƀN����zn��v�Xn�fK���ꃎҾd�Y���prb����P�/��s}u����k��g�c4�n�sAO���Y8�Pn�$�{��[W����GvQf�
��9���E9W��]C���&�w��9b��(,:�����Q�_cC�|�*7��ۘG���cW���{��K-����b�Vŀ�=�}��j�ND�U�,)�D��93�dV�u��t�t��u�]�����.w�ۏ,��]^�[JcN&dQ�*�]�e'o*�i��!,��(� VϦ�a�r�+���/6qǲRv�ʀWr�O$}�f�-����ދ\��~�����d+�;��d#\�z,���K9��T'��9�P��VǓ:��K*���L�7H��kQRމM�f ��`�n�Ƚ�YT�t�ԲԪ��Y�2$�Vl�/��u��Y
�	
 �{ʠe�uU|��=dߜd�'������J	:��u�eB�֎�t����FI�dD�z���S��äu@���aǰ$�C�'T�����	�V����L���f�E��]�<�YfZs4���W���*7Qg�������|����7&�He���D-�n�;�Q�{��;ul�P�f-�ֵ52Xw��s��vK�d���XU����͏�>�m8��	b\��o�����m9�P�߅M�qY��ߺY��M#a�yҙ�w2:|uQ"�,��Z����eȏ�����fhn��ʥ�B
�U?+	?����1���\�L��W����Nʍ�)�r���l�5�>Y��񃇅�� /�����D�Q�P϶x�ٶ���&�|K��t�Ј��w咩Ѽ�[qU��������S�X�.�;>P��d�A~U�Á����ȼ�DA����Kp	/`<̌S5����Qo'�ІI��E�����6#�̐���;r������k|�w�<�9I�=M-<%Y��ɓT.Qp�����C��=�h�S�W�&v�Iں+�P;�|�Z�|!8*U��3ø�b��k��m䪵#����\�EM���S#����1DH�ފ29��dW�C7��k�Tvb���A8i����u$`���q==�*:��������Ô�o��e����F/n���M���0��w����҅��--d@��]?r��,:▶2�VY⻅�5�i���o3������k��*�˒�.�`�v�GC]x1�h7;����㮻��yƇTS�F��,ϗ:F�8��rcN�T�{
�����w�9�'{&�pt�צrE�n@n0��)f��DHIӘXc�nq�r��A��p٪������Z��(��E�޿T�8����(��;jA#�5Ki�J#m�9�+D�7z����(���D�{�����dJ�N�V�Ό�Fa�JקV9��%L<mVy+�6hB�j�J?3V���L�
eC��U�%Ҥ��Ge]�RѤEUtz�V�P���V낡T������>���K+���c$l���z:Ev1�r|4D���d��ٞ.�I�V�"�L��v�˕hp�Uv���� �QJ!���Jdq�����M��pt���]��X/�4��Y7�H׬�����U[��
��*������=ޭ��I�L@q���hK���^O�|~�: X��gx���Cs]���e�ԅ���}�=h��j������aZ�q�� ��)�P>e�涺o����\1�E00����06�İc\�h�Z��д��=�rNQ����L�vf��l�\/��u�yl@5X�&��9Y�{�V1���+��=�)�k�=�5E���3��4�E�~3��\�3/����rw�M�f�qS�ƶ��wN��C�w�S�Tt�%\��~��\f�ol�1HG��m�*���O�Z��pX��l����#g֨aoJ�C�>U�o�%���	U!����0�/��5��[���~q���,����|�]w�:H�����J f\.���k�Y�IE�Qgi�~���B��-ř�#`t�h-�)E�T1���1��씹[��Ib*|$8E;8�Բ��P5�C��Ks(بATZ�f�k�w$Z�+�veݠ2�^���p�E\q�NY���D��t�&fN�H�Fw3��n�H�Qt�Jp�1#��~�(�����X�3�?�������[,M,=/+Iq�b��g]#���1O�2˳��e]~��ם`��eNgijWi��h���r5/m������J����g|�h�������V�u'���q��IW�֑8v�������$[�F������c��UaY�������Ωr��ES������O\��qE��f��X�G)H�]�H���5Ze�w|��SI���'�{�8�{͗���>�d!;aD�Q�_���&�)S�x��סD1��DS {���MOv��b��)���/�}�I>��<x���$.�I�qI����30�Z�_���ҵPQ����'�>c~h�/PĂ��^{V�Ʀ;���o��Q�^�����5�B0�G�(׮�~�dt�&�\��p�;7*}�9ə�M��C�Ti�ZW����P�tCF3[{�~����OLd��c���v�~��,9�ƻ��_�#�i�����6�#k�t���t�WW=[���v���<��r����WY���E�{]0Z������1�/��Z��	�T���D:��DayM�%6�ˡ_d��5֦8�̊�B����~�x/�,قR;	7����\q]�������*F��t�f�e�ծU�Qߖ�u͹U���P���lk���(�\��ӛx��Q�w=Pywd�7b�2�3M�n�)Bb
w��$���GK(I�8)՚�:wĕ����u�䗻^��׸��
�?K�6��d�x�j��5v�!�y��]�� f_=i(�#s!�.�o���W&�| ����{����]�>|x}�Z:w��ڽ�
������h"'՛H���j�ӕ����z�!E���2��_]3a�w$XH鸒x��J���b=�P0�Rn�^v�c�k䂬Bƚ��d\�C�:DY��3��s�}G��WWQԏkSOY��%q��.��e��rc�:�:�P!CS:%ϥ'B���	��W+���gk�����G��Əゝ"���/�����S�>>t�z�e�E:$q"ғإ�U�'�CI=�%�e%�V�ʥ��D�}���j�)2ȯ(�.�:�Wǩ�	v�F_��I��c�m���Dlkӗ^S�n7�"27��Ni�p�ofg.��4D
��5G�3�}�s�L����ʡiW]5Q�Ub^zQ�DM�NВ ��lr
��B0d$�?rd�dh�\� �W��F�j��U�mk�8��P#Q�%��B$�@G��3�*Y��	{�hV�*�oJ�����Y�Xx҈M�Y�g.�����ۖ.��}Cj-�(��7NEմ5+{�eU�R���Z�s˝���*\�t\���;rC:�|xȰ�����%-Hs��6�e7{u���i9�CqX��I�d?�}U���������,�̜<6�ܭ ���,w)�R���Rǲ(��IB�J���M�<�>��,Z���Q�|=f�(4�24��B:��qx�"҃Wq)��m���@��;C��|+�X�݊�X�N7��db��2�R�ko/��n՟N�kP�9��+���ꁪ�:�H���@���u�.���*�<!7�8y�:ŏs�����w(c�:�E��Q�<�J��+�� (�� ��[�[�x#J�8}ζ����(([���^Ȣ$$��,<�P��d�Iomq��֐S�`�)�x��e��{���Rr6"���n٫R	�CtD�`�ٸ�5�ѻ ��%�M�E4���l�u:���B,�y�A����%Tт��MR8�S���Ɋ�*�xVJ?3hx�y��7��Y}
��{-7E����&@����n����؎IT}�뵨M/��+��c5��yzuĪ�����{M�F�`ԅ�G��c���ų���0���Pbˀj�x�8�Շ��Crv_^Tk�*ŗ�w.�D�w��g��W-v�/�G�;�v�XVu_��a��wu-`Φ���mC���35��`��Κ�($�ʜ�%!�n	�֖��7�a���Rtf�sj&&�`�'FWb�������L$=��.9\u���H�h��]�r�ڏs�B��V�nq�gEE���r��Mgc�����ͼ�M����9.�e]�N�T��X�iP���,E�N�'e�eР�_R����90��=�1���Z�D����6���7!�x�ΐ��Й�ՑC�5��M1vL�sgA�E:�{�hv�L2��_!k�L���G&�o-�M�{8U��E+�rؒ�:��k���m�oŰ��^�cOk!]��w\R`��9t)�*���)Z�1�Ta�����7:�`�an�#����JL/N�JK�[�`yvE�;�fk�l�Z���2�u��ݡ�Ɋ�Z���ko�KF�n�����WH=��;`�#ݛ�  ��zh$\�nt�t�}u'�t�+�x���/����J�i(�{���	,���k���g�
D.�S=a��]ƒ�	�((��D#	�K1��+����jLyg�����H2:�@�N���Rq��:7Hi��E]��ڊ�H;oy�V�2�+!0�� �ݒ��T���i�.,3�9���^݊]u%�ʋB��v��K�[b��]�/%:�x[�,���e��V�;�oxe�ӇNY(���A���bn��f�k�,��;�y&�]�P��ۇ���ڨm9jl���n	|��H�;:��L2�f��Jq��QX�#F�9���l{&I�\��CN�R+���wVv0p�4|�U�M���;&�O��n#s*�V�d�5����;*���-4*U:��k�vҶ�z_=�S�W5S���;@�J�t��=z6�����.�:{�Y��-���8�E�M
����_�w������4Z�+Ό�Q�����^��wB:X�hf��R]EW��e�IEa)����e��g����).�[Y��G��w2`���v�r�7d�Yg)�%�W�}.%u��qӼ�sCq���1Y�6�����;c:�f��D��Rc�?+A�6:�;��u��.<Rॲ .��\. �I՗�-C@�C
�cs�}���#�Z+����3��.���c�gu[�%���2��������t��P1\���\��e3&8��3)++�S+d�Qs)%�HbR"���T��̲�eI1�ŕ��@Q@1��n8ԅk���X��"��T��Į8ԅeABWRbEQar�0LJ�Lr!�)�����Z�0��2�Y�LLC1�b��̳2��QP\kr��\@m2��Lds.0̰Rc*
��1�d1��",UI��"���TL�倉�Z� c���� ,�A1�11��+�� )-,3%�bVVE+��r�.�e�Aeb�+b�)mf%f0YR��1 �1�n�iJ�#n$�e(ȸ�����
J�[���}ɰL�s��V�ˁ��v��f��Q
�<_��w��?����z�^qe.XzQ��ܴ�m��,�ϕ���yW�����T���}���N��U��?�]ñ���W�ŁI��
����t�T���w���)ޚ�.��,.<�+gC��ݥ	ܽ�7��ɑ�L���Ы�X�2�F��U�r�7��N,�Ŀ��{������-�f*�b�;qp�e�|�Ɛ�v�K��Y�6������jz� {ۛ�x�&�D��Ui�k"ժb��0�(��,��u!-�R�1�D\���Q7����giT�.��p�4A�oE�x*��]cB���ƃ�ũ��2�q�kc��3ٳgt�l���?p�>U*,�|}8V��]g&��Qw�C�M�k�#:��iGqd�g�[�,Apmd{���)��f8�ɴK�e��Қu尺+���n;"���'-tGa#��2��f�~��y��v*�x� C�(��vj^B���E������^��Mbz�uY���I�6�n-b�;��}@�R�I]ϯz`)�	Q �Ju�gSZ����ݻ3\�9�	�t+\`�֫�ѧ;̡���e=B�V;�+�3&��޺�*Pֿu�����d��e�����/]�1S�;�������i�\����㊴:6�����y��-�d���4)�8��LC�d���#��{�'dǲc�^���
���i�O��a<���D��y���|^4�w��T[��w��^��8�����
�<�lDx>��>��.����<1����ʽ�.�JP����y�>G�h�m��e�0t��@C̴r�V�(
�:bm91�5faM���
_�y�҈�V/���i����p�`��}"n��-��g+�vj�X8aES�Cg�FϗDD2�Iq>S>�uD=�g��P�o�;;&�I�>V�U������(������c~:��*�@s9�1h�]`�;�ϊmI�aӧ"�v$9�=v����WMm��ȑԨ�����k%>��^p��W�Wx?�^�B�ƳU�Db1��k�Ӛ��"x�Of�+/w��Þ�*�q][�<i���;1�rړ��ӽ&(�c'���]֥��,_����E	/a�al��+�.�n�+9��51���.���<<*Wb6}Zh�7)���t%&�m�[��[L��)�ޒ�������2F�dr�2*�qyZ�%�e�֪�H4�xr5b�"Y��p��1*pJ�A�۷�{�N����{�	�A�]y<�ȃ޵0uE��G��	��4ky��I2�Ȓ��=� 䋔�߃�.�P����5Ԧ4��{�(�1��$�^�]���˶`�� :���>��;h��}/zp�N���I�Q�8�$P��Č�~�P�\)�[>*d�8�s(�E���W�],&��0�ܳ=�!�cs�Zv��Y�}�rc���'�����"O�B�y�h"�Z᧸¬�@����.�G�:�B,Ⱦ�fۧrE��t��#C��0:$��h���"��)���r�y[C�S����.t�(�ŖP�* �}���k�yDoN�A�j�P�8^�3��Nzc׮C��:�T�jf{t+�@q�T�kr*v��;���2�z�a�tP7J����L��FK:�1K��|��D�95�`��"��w��=���`�_�?(�ڡ������6F�P�;|?i�������a�y��a��ǜ��6�xM����o�5��"�a��w��U�Ve�5	��[��q,��2g^,-����-E�-�Xy�M���}yZ�>A�KP���M[tV�y71���.�̺��D�b�Z�Db��%�:d���O^e�I�e6�\��[���w�`>Ƀ��°�9u�96�@(����5�r��t����7�.�e�
�F`��w�ك�CϪ�ڝ�]�*�����z:!7��X�X<B,�ا�hq����̊~�����s����������:������C�DMB&��3����.^�����,�~;�J���4��On�wL���8ϙ6|4dyHɓUsę �IM�R���EikI�P���Rm�Y����`��nփ����9��_ݢZ���ߒ���6���M޽��Am�e�@.�CnE��A�<݊�X�3K&�g�xpk���f�W� �;ޙoQ���F��F8Ѧ��]�DR�Z���:�p��x	Tn��;��ǅ�;�Aۑ����6E�\��
aYم	�l�v2E���#-�>q�)�er�6=�[AWK��ls�q�̑�:s<c�B�z�=]]U�����:U�|�3���W%�	6���9U����E~`�n��I�P����
�vi,�&@���ޖ�}n�u������3����z;v��&c�Hm*��t��BH�.ne$/jԼ1j��큽�$�Gx�*Hh��wHD��ҳe��_�c
NF�"�\ݲ]`uDU<צ��!�i�gCW/`�C���%]M�E4�TO��x{�}��t��r��tN�<%������x≠H�@9��p�5�*W��²��<x^�D;���۽دQ���~��s BN���ԓBz�W1�`X��aLT@�p�%�x��}��=�mwS����D�:9���2Q=S��W'�D��N��k1q�j�g�phb�j"㋠6��� ��24B+�A��L�7�U�H��Ū������~��X.wb��܏���L�8��Jh]�i{sQ	�����Z�:#�ɜ"���B.s#�ʌ�C�j���ƸX���-���y-�F`Il��G�Ր
�P�]_kv�V��k��eU����-�/��ɤ�֧�NF��yXv���6u�H�iQ��X���3D/��.�UP�m��i^Ad7/�i��/��0`iA���'/q��N%��n��1ymq��+k|������o=����ŵ��
Z�*>Vt���7r��M�[�8�&]�8\��;v�ŧ���M;hA��ت�';�g���QE�R0$6���졥�"�!��ͬ)9S�į�k��4cb��kN�e�팵����҆��M7#��Բ,8�3���:Dql����.p����1������x�^qL���EL��m߫atYE�R�dI�������CE.���K�"֠�E�HLL�$��u\�;P�Cޑ)
^G���|��Xx�%��I.S<"R�g#�"rO(�T�¡Oo l���5Nq�f�<'K�x�^�N"r�D�{>e�U'���Qb4ϕ��E]<�Q�j�EWJ�%w���=��!�-�tq��2TVC>�sκG�x�#���)���da�	�Yb?^^��>�3eT0"�pp��ȣ�yƁ.F�蝸d�ly����ܩ��w��>�5�UF�.r���8��D�
��qR�y��5I5�T����^�D�37<�z�������;nYܨ�7㈫?{q}��J!�jK�S>�ʝ�ѲbDȷ��yZ�
Ӝ2�m��aK�X�*ՂWAU:f��I>�I
�E֤�s.�	`V���|xM���V]ub���o�q�nfٲ&�YR���qok��+��CI}`�\�Fs#�޼�+��:���VZ��&�� �A�{���\�n�Ȳ"�Z�fxm"ve�qD�>�g��uӶ����	�q�S&%e(R,�J��+���F�Y�>����>�³�ZSQ9�� �2��&� n�<�J�F�w���`����h�Z+ؔ���P�V���]�+Z��������>N���]XS����玶c�L�\��FLQ�oa��uv�s�-��^�3;�uƁ�c�a1�n���q{(^�,���p�z)�r�j�;��y�^�^���n�9 \��Ï.�P��v׳<;���o�#��� ܦ�+ojf;�i��
&��s�tkB������׎[���9�ut0��B���W�Gu{DݻV�*p��z����ۛ�v�V���P�s�m3�Mg��QɎ���M��[�b1��KE��?W���*�Zn�F�p뀋.��n�����e����-�Sα+ą�d��D:ݧ�u{�^���w�.`�N�%��u1R���)DI�`��o1z��W:�m75�N��SU&P��1mN�ѻ{f�(i���l�b��t��a�w�%�a�Ԅ�׻Z�m��5Hh�q�M���\��H���v��Zߦ�es��:DY��2́JTA�Ι�jR����T�Ie�6_��'����qu^2��\��GT
�-Lܹ���Q�=Wr{㕎��DǕKȷ3��͌#A�W��g^�P�4F�|�GCu�E�Y�:c� ��5&Gd��<h}2є�I^_�K> �@]������Ǝ��Z��d��K�*��$�1s�T��B59u�b��ŀQ�"
�u��Y�����Z(���(�\�!@�H�tw���.���[@��&�����GE�悱�6G�7�Ȁ6W1P�O��ȧ�@L����s��"�9�y���ɍɢ�*7
�K;@Gc�"�5���КhlF���؎�xM����K�
��J���,��Q,>>�HYQhܧ��R�%����(3�����o"���N\��<;�s��KE:��3�oc�WK�-�L�.eoW[(�f��@j,��b�������457{:�?h^�/)Cz�ۤF�M'������(Aq#D�=�|�p�|KEh���9�+��b]2���i��<�y�gnZs1MT���z����ۄF�P3g�Ϥ�S�Fi��_J�]�U�`YW�����K�p��dW�8�ߝqu\"�UI	��i;
{kuI/زUSr����a���r3�����F�P�,���fW:F�8S
��(VH����c���3�	qSD��)9����
�K���p���YD���'��B�;�O�CKk��,�9HD�3�K�H�ޯl�8	�؍
i�j�Qׅ��nG���sF���"	
U�*b�#W�hc�j���
����s�~ޖ���CK����8�iT�5�;A�a���\��#�6�z�C��Ǚ�*y��[��G�U�L�w2$���I��\_`]�C��L$_4�s�9B|��1D��gM$@�0���AE�r`��3e����-�<[Q`�0#���Y�Qj*�Qy�v��g�*;��t
��B#E��{�[���h��h Yƶ�Z�^f�Ac@�Wk�u*$nkw%�4ڽ���jxl��J��m�j+���9�Y[:*�����Ewt�5e�ӛ�.���9ΐ�t�F�����2��0��p2�֤A�6V����=����]a�FU2�gGȥ7����9�m-n�D�l02"�PRg��9�9���[9W�a�����}X�@���r6���o�I�Fߢ�zGd��^�9���A���^W�|j�u�e��&o�Zw���R�Ѧξ�jD(�,U��h�xދ�����E��ӻ�9�
�.���1P�O�l8�l�ĝ)�����D��Yj��
~ۦM;�~��Y<7���K��j�uz��<E�*E�x�崦59��:l
�n�Wm��"W����@/�XЩ�cқw���諄^@g�5'L�����]-��R�Ђ�L��PQI*<7a�W�k7<Dc�eJB��щ|^r�OJd4)4�tԴ$h�\�� ��~�E,�;����5z◭\1�-�����6T�Oar�1��!e]<��D^����紣��4;
��84#>͕Q-j����1`��K�V2���Ɯ�YL�}��r�n���&@Z�N��WYzS!+g�ŇTN��t�`k ̱gw��V
��Z�T�]J%�5����99�*�:��9fnۧ�)�D`1�\{��;v�
��k�:mah�e�r��s/*Q��eQԫ��ص�\�����5r�Z����xi括�PRF�v���<����+�1�F)XޭIǬ��\�{��n۾�]�����O�dt�R�@�\�*
J���Y���6jуngZɂ��4G�g��xa{ؑ�˖G`,��s��{ݢNc(QqT�
t�Y��j]]׋��{5��c�8Ɖc*�h�s�����5�.Gx�	7��l�)]�ɫF���3���t�u o�%\�f��K��f�Т7G����n�^��{/u�-LE҅
���B�F.�
�p��U�V�]$���{�^t(�k�Y�v�]���xhn`#�~�w��}:�k6�}n�+lԀe�����r��C���h5��V�f�I�D��$�o�cٷ��}Y���R��99Ic"�w�ܩsmv�
��#7T��F�5wj�l9Ej�ڷ�eZ�:��s���/R"��{�.��Hv�㋙y��oj]-���Y�t�cbf�Jw93���UÄM��v�inX苳6�[4N@���jY�Y�F�ν���Ovx�E���x	� ��rB��}Z5Q7[(�ܽ���_tR��TC�X~�ՁT�C�3V&�7w�LI�9�p���#��RG&s6�F���sH�mQΥ].>�����Ƹ��rW?�w�x��9�a�T���|0n֌��
Ή
R��&XX1��J�� �6a���WA�����[�Jmrk�8��X�h�,g�kAru��q \Js��WKS��3����4����X�*�J�nԒVD�0x��E�$U���cSk0YU��krˠ�GfI�b[�ӡ�9�@a�g��ě���ڛo�@�k �7&^�F�r��`?[W��_kY7'�{/syQ�Ue�=��mv뱷nc:눹�V
��p���fk���j��8�s��Ty���ʕ��.�5Ԝe��G��+J�GIL�u��6ε���Ɖ�b�c��pW=��2��,p�rSº�w2%�H��'z�؋{K�.-Ckg�*�:O�$����u�&�m"A�:V�d��2]���>��TڷE������R���Ɯ��V��hYo-�7�����:vjؾ�ح�I(�}RrJHp�w�� ����b�.Z�bT̲W�
�3,�C.`�R���������&$W,ƙejb*��r�J�"��Q��Lek%(��J�D��dr�J�,J�c�D�1�drܶ�LJ����A.f(����-E�AbV�[�
�-l�+b"�nZ��+�1"�1B��G��ی�[aR-
UE��ʘ�1*�(�1b�+�S*���*
��"���,m&"��\T�(�ڗ.&*.!��U�m�ZՂ�V���6��d��EA`�2���mX��Q&5�(���1��R�-���B�h�`�-��P\F�Z+amcnR�q�c"���cDCQ(�qAeaYU�1J�jW�Ř�(�0�1*V�#i�����ƥk(�J4faTZ�QIQjr¸�1O]{�k����s��5�r��T��7#t����{Vzŝ���:U
ޥi�5z�}iu�1��d腹��57*bVU���u��9*Y=Q�\�3����:�vo��F{8��\)(}��C��Y�'g�T�I;&�� O�di��yT�j#n�/��mC˜��>�6�!Vˊ��AgO��D�v2��\��یm�jǾgF��?��8}�E`���ى���>���1��e�a������<�`���q~�,��Ҍ\
"*)Ũfe��L�S>���Ruw���dZT��y V���R��x�5�'����C��c�{}&=��u��N�v���&�w O�#��I�U��k5P;��h�kJK���n�A���K� ����$�إ_���A���;1��ԝY��zӁ�t�$���s�)���������z�����{�	�A�]ey=7�E�x�Yx���G��{ܶ���1Xí��\�L���&�R��.�Qh\����y��;e��Ԫm��KFaD]�2L�_��t_���^"��}|�����1�	 �U-�1(��:��؅F�΄j�p��X��Od��*�S��e
�ؤ�@�P*�s�wÝ�N�@�6�Е���qo$r/=lj��f�S2�d|�[�w�|��O�Ч~#)�����%w��H/BQ窐���ߘ�`�0�\t�P���������G��]Xq��[Z��Ұ���n/Ŗq쳚�Y�t3��`8�*ĵd�`�����5��c{�&�@g�m;�ҩ�p4�:�	�"��ӹ"�t�P�4y�cM/��?wW�ހg�{�(Ǟ�Pe�ϔ\��� �P�P�Y�R�p��]�2,-�D�S�	.��>fϣ�WWP�\�{fYyӓ����t��	R��ːN��
cb��J��P�𪐈�@�#�^���(^�`���+���#K>t#*�(L��;����of."��$0����򈌪~�y���}qf>�G�ox��F��W����.��!���2z��D��#�uT��Ɛ�eO�VV8�F�1���7z�0�ADD���ԫ�����$PP{qT(��`�Z�����7m90��@8j�3q�C���Y��eA�C��y@��Z�ЧC�b* �9�q�N�*�6�d���]�g�{;�4P��]�/&�p@�cGmM\wR�xo,Ѭ��x���^m�P���Xv�&��h��%�&��z�r�.bU�B�
U���P�OITA�&���{#+��h���c�^�Em+�!¯�x}g��� �.^��m8��c�s/��D���)� ��=�'r�_|�:���`��h��,�5qĜ8RS��v�����E�<��V��t+4�,x*||�:6�	f�(4�;�C�,.�����?��B��N-C+>����`Po��DmE���<݊ēFi����J��,b�}���w!,k�Ed#z���@�ҕ;.�{�T���kM��O4	�^$�s�8��!~�b���J�w�K#�dY�ΑC"r^�����*���� ���f�4N����um��)}A�/l����E�׏��\�3��8n���-9Awh�/3�H�ޯl�8����8nq>K+h̝��|hZ�0G(j8D�ybJ�T�dQkZ=�<|�����=�F����L�WW����V��*��B�Ds��s�>� �g�k��XdWi�u���GwK9�X�F���v������[z�N�`�k�W�L���=6�ĵ�1�Q��+9\�R>����J��7V+�Z�\�08�x�J���8�h*�ƃ���gLb���,��~�\��R��Ψz�-rh�s w2$���I�=L�TKܰ��Wǩ��D��K�hr���]�#��F���t"d�Q��;v�<D#��Y��ȯ�
2T�y_�q�~?h�6�.{UH�Y��
�6��B3-]hE����>�/ss�4�"�&�~��l؞��Ys�o����,�8��>F'�B�z_5&dC��!H����|�І�܋�!��a��� .��!k=ݖ��';[<��sg8�<�;�(j�hC�n��B����e���\�6�.iĮ�u��x��Xz���6{J���G��PU���	^I�������g��#�᪣Qb�b��$]gPf�J,�p�ٳ�	:S`���wozϰܮ�m����a��hp*�����5E�#���s%���[0/31�ɔ�.虜׽�EK�zxK��`^�u^n0��Gs�^[fų`�wCW:�h0*ήͅ+���vk^�����ˎ�k;h��Ӳ�#ڒm�X��;o���Ct�2�r݋g=�̧$<��#��7�~�L�æjg
������,����kL�u9��»�r�IR7
D���r�+��L�S�#a�W�vj^B�t�S�݅�V��qm(52(�Ϫ�[+�K��Dpv�s�l��։G����V�:��r�n7u|:�ZrAޘ����3-R�=��Q{"|�&�SR�Z��y�4�^>�z"m��=A���:�3�ʙ*+!�HW0L�z�s�N�=�.v���[Zʘԧ��-�diy�Q����|�8�Nɡp�	4gv�����7�o�Q~�ܴr�V�,��١��q��&B����R$�S֬ZӞ��qｾ洽��j3���?�Q�r�eE`��刧�/��ܫR%���GWM�̅iV�zs�!�Ϥ�v"NC�
�pp�V�
t��2�33[H�����a�� ��+�B�u��x���Pݥ
E�������Y����z_��T1[׼4�z_6miא5�f�*��^]RloV�6�b���6�%̜�!{J��]��wZ
���_SMϲ6ز��r���S�5����]wmY[�8�{X-���ZO�@��4���p��䌬����J�D�@���Q&����O&s���뒶�Ӂ�|r�҂`>�[���i��@y�/��`,/�%x�Ol��ړ��x��.��WwL���ԋ*6��IC�\3N�_a��XLB@������5Xf�k�_es�I�J�EP��d�]�#�%�鹕VE����� ��IJ<�5��óӻխ�i��u9�<�"�\Y+���1����b�tw~!K1=DY��/%oK>��*��9�*��=��G����Y���9�����qVj�O�E�<m=�v��>�t3�Lts1�C�$9�	4�H�M��F#Ũ�3h2&�ip4�:��f����Ԑ���(<��n�h�f���4_�z��4�؈�m{("�g�g+�X�:DY�Yт;��#�':�����-$z�߇΅��8�:�yAp�꿑�N���:�P�-L��!��If��s��w'b��v�`=��T0'�v`���u_�r���c��4#a뽳yX�gX��$��q�Y|�����գy�S��}�F�����.�p�rc#�U`B_&uqg������{}�9١��w�:.��	u�B�L���Ne�Fla&(��}(�Ȕr��h��m;�g#�5%���k�\m��TS�Eyy��K��I^������`��Xa/�\� ː���ͽ�v^�pXwG� ��d��D��#nyT����N]yj��ι:^ѿGD���HvOC�∌���*g�Pw�I��E��`�(�3�h9V�����Œ��{���FT8;�
�xR�/�x�qUZx���A�+��1�mn�z�:(��2/��3�x�L�R�x}-xc��>b��ڃ�[-"�R�os`���s�8����k���Ь��)v�g��vZAà�0ﶎ`fbɻ1����_����G��S+�}φ&{���eq�x(4�;��#格��D5���1Ed=�+�\����Cn�
�]V��I��$��F�mr�ܦo�{F�o,�w27��e�,�(֩��5�5�:�H���������7��w<a�I�:�f+�ɜ�-a�(��U���{��>~�I��UyJ�Dؙ�(mb�*n�p�x�f��}m�Sq�kk1��4�W/)[�z<�'kU>�B�v���[m̥��yP��|[̚f���M�;r��)�ڮ�hS{AZ������ �� �S
��!���:�E5��f el0�����{�i���K<EmS	�W�Z�SS^�N�7��Ҷ��"VOL&y���(�r� �ў:^f�.����q�q�*�=�,wkw�)+�b����q@��i�@�].R�«�tx/PNf�D�ݨ7+ME�Lb�,L"T2v��`���`r5���{j��h�J���f�]��[�զX�E?��8�g-��$��I5=L�T���P3T���oh�3Q\vD�i�4�#\ÇjG3Q� N)���;�0.}2�^KA�%rT�\���gC(���<o�AGH=:dh"��)oDt��{�*N�\�h���xE����Y�f�@dNB'&Yy�PHP�ˁUsV���\�z��#w�.3�"��1�t��vu�g*�>���/6��yP��@���ۡ�Zg���s �j���S�Nu�)T/g-�nu�;�b�U���D��ѿ[�i�����fa�f�xw1%܍p\�
û}b�S.��S��!6r`(�+0��}��U�����jv��T�w�Ww�ݔM9��q�p�����Q�{�zrE^�8���gE�6�]<�M��pH+c*NPs᧏.�=����5�H�R!E3de�@��uK��n���S7
�т���*H��AЋ<�3#�k��"lg��旻��P; �S��X��qʫK���_�z�Ϗ}�R,Ҏ �:z�b����҅Y܎{���0#��]���`��V:Pmߴ���E��6�U�MXqys���+r�v��=B
؂�8���
|4��dq��K�W�̈��{nm���4��4�C���U�Ks(���(д��w� #Z,����7j^I����ۼbC3cWNtX	�(��Ϝ��3!�W'���{dO�+��D�aE�ގj79�j�'�~�E��D�:�K;6�J�,���dk�yFc� �7}�x���̀[����գ��#��\@W��5�"��8�RtN�5�V�h7\ݟ\�|ޫ�;�H�J�_Qq��+U.���(J�Z;s�|>�w��+�E��zq��hc����yj ���Fi��p��i`X_u��%�k7zf���	�E�'���3���@l.�$T��Lע�S2���'���Qq����Ɖ���.*]�"K!��b2!�Ɨi��M�l����G�y,3�r�dV���Vb�ʱ}Ƃ�r����g?8A�tk�-�ٟeU�y$�'�
������/���^	`�_f�lA���ns*��%�U�PQ�ː<� Vc�ʥ0�H�����c!�N�ە3��
�@���`m2$u*%�lUKrռP}��]�k5]>��k�M����{O���#��5��cSƀ�g�9�N�P�<[�7��`�n���h,�y��v5����Bx���%��*ZcVg�f;��P+��ɛL��iu��jWYc��A�
.x�:v=Is��3\J��DZ����s�Kl�u5�-3U>̊(�{^�u��:�6�.l�)�5|����������X�K	��ay1Jޜq�s��tH聖:�saʠM]^*d��!˙�wV���3�wf��Y|󄻢�J��R�s 8I��b�(ӡb�a�`�qZ��j+��u��x��;`�BݍY+(��/�	���(�*�9�T����h��;]أ����7��������$l+�y@�u=���)�W8U�,�t�"3#s�v�"���Al ��V��NoE�%�v9V�L�E�������ʸ��
U����H��<n�!�-_��؁C�9�Ah�ͳH�ّ�Ϧ�v�T��n��;ֻ������>�v�X��B|���F���b�)N
v�t�Y��BS, K'�WM�a�ݷ���t�	�z���{kp��-�CN@W�|��;\s��#NHGG��ݨ+^��:���:�4%Ҧ�<�P�l�Y�em�U?�p]'v���ݔ��pz"��M�<&���L
��^�[�r�ٱvS�{�^�2��o/�����ے'�&���,�]04�1l��Ί�3'.�@
+��6^C���R��^�w�e@���s{�Re��Aq���<3��+a�t��}0�̢R#�6�^>Ù�y$�_r�sM�h��yʒ^5z���-�l��KE2��p#�e�Vv�.��kj���}�a���Õ,VJ���a:Ύ�఺�_k��Sz�a@^=��&��n�y�/w1�P�`��:[�U�#�u��G���uw�I��0d�̢�m��K(q�Q�V(� du}l��yt�5+�8��ʊ U�v�m�H�b�ѰAΒ���:�9�Y0
�$����Q�y������m��ȇ�����Ve�f���js�G�	(�;����j�и�,Dh����T�w�bѲ�W�]�V��6��g�V[*�ղ^IZ�+�h�z�ܧ�L+���:N���L�6�[�R�>���H�Onf�08dw�@CSI(�,V�	�2`�سvuaE\¬��M�Y�,&	4)�j�U\�vTO3&�+�����f4�W!tqՕCvUˉ���ck���9�z�q�+��qr;OyW;n̓,w>�����٠ܟ�*q�����5�����|R3��U��~�>Ӽ�|�}o*�(�hC�|�_\�.�Q-����o8�;N���^�JA0}$�@Z��&>FD�N�Y��%��ncO"Tss9�z��|$�
59`{u:�v�N��K{acJ��oSuؘ��K��\�V@r��x�д�m�.���-69YV�E��|{uw+��P�Qt
��Z�"ڜ��y5��{Şss�|�����ד��`xΟ�%X&4�E�Ak�+X�ֲ�Df2��TD-�\�-1\AKl��D�6�\��C�T��j��%2��T�˔��m��k*P��bEJ�3,
%k e�Xe�)��e%IR�֘щh�m�5b�1*Uq�(�6�ec2��
��W�1�d�(��a���Ղ �K�Ġ²cZ�0��UV*����+ƱTr�[m�a��nc�Sq�d�E��L�+cU2�XфR�(�
��r�#m�kR�)��b��6�*ª(T��q��H��-��e�I����娉Xe��G,���(
�7VTPU�	\��+R�\Ŗ���0Xe�c[�I��\B�cږ�AF�-��+�%ImX��VKj"e0r&"���1�\. �
������(�����p��L�-�Z� K,gei|� <]y��;���FX�T�'�S�ܕ�vÄ1N�v�"��%����ee�ēt�*��oX�4I�ub�w�'OP�Gӽ9�`�g�9�U����_�l�a��;�c�|���Rڙ�$��(�q�`���H�9k�0��"���t�H�V֝�oJ�ɎKk��0M5m�f��}۹A]��6���
!���Y:��&{��L�P�<$�b��A��#�8} m]]Gg�p��e�8&=s����:�b��s]��Kn`�R}�/+T{�_� -k���<0^�E�����p��s_.w��p���$����\+��*�tH��?��6߀��^
b�Z�F���ڋ՝6TvF)��NMC4�dR��L���I�.3�j�����`)w�#�n���Vu/c�]c�,���r�t|����Qaq�=�S��k$��?ga�^�!���J��SUp�{�8P5��_��C��������:v��q���;��C���j�����-hg���Q�
T��Z��t t�^�ܣ�N�{��'_W��Z�lbҪVfӯJ��=�~GfvV��4Wyl������ӯTwR��x�r��H��I��
�\+��g�����"z��z����ԓ��+��P��i�c���&�`ڇ�<Tje��}/Ηb�'7�Ь��l ��y��fϒɓB��m��O^�q����o��x��g�|���RǪ�"���iG��6�g�x������,�sDQ��B;�a��{�B-oP鑅��l�U�(}]FK�;�V6��t�*b�\@Ů�(֩dVB7�x�7�\
n]*��ul�$pa���B=�x����9ͬ7�.�!���oh+��Y�(�\���u�d��6��J��1���G[���n:h�<[x���mF<�("���z����{��bl�qDO�*S�%���$Aݯ��m"����U��;}k��^�KQۨ^��p�Vݳj$��Z��$%yBJ�Se�4�ver�}�=��o�)�=Ƙ)B�S�,��Y9�[0k��X�����קԕ�F���?c��O!�� T>r�vz�$�G\uC�P� I�:��.z�S�b$9�w�tȅ�9��T#��i�87�W�]�a�����hW'-��E�硲a �;��kCF������jȻos�KfЇ��"��w�Jf�
��޸�A	��uu�lkK2�fʕpw*f��s��\���\����SqnD�H�D��0���2Q��6�E�MMDsr�.{�n����p����uMe��l�8Q&�u�NQM6s�^�yo+)	fi�<k�dq����lONd&r�Vk�U���Kv�F�r�4�s�mid
�=�T{u�n��0�Ah�厝Q����^��0��Z��cX{�����E.�>`LQ&]NNl�G(���+�T�p���\�Ch`b:bz�IC��?j��������<��S�Ѧ���"�H��l���{-y�ƣb �~�o�Y�/k�'�jH��"�g�dvmaIʘ�';�y�TSY�3}��kh#=
� �LP�.w��L��;:UƇFr�Yݔwͩ��y��r�o]{}5`O�.h��Z�:% *�	�J�O{�燴ʟZ���<͜�߅�e�+��d�L{PV����PW3Ē�¶�~8��ioW����3��u<��.��VmZb�"���ؤt/��4����}))O�� ����,%RhYW���:����%9�����{
͜Gi�:�Wt�%j���sr����l���Jj����tq>�$���y4��r4wmƥ!�qY�����s(�0Q��!PO���U�����tU^�i:��w��dqp��8�ӞQ;{s�d5J��娽�>��dYӽ}y���1��	���%�[��e�#�qBT���������&g��=�.���ž�ɮ�\y��,�y�7��Y��B��Y��"���.F�S;��+���K�om�7*xM"]� 8���f[9O�j\�l���8����!W�\T���j��j2��K���#���� �D��.`a�3�C������g�+��|��}��k%]ѣ��MpI�\s��L�#����3�����<*m%��V�
0�q+Vʯ?b���w�EpK��
��=(�$��1�*��9����F�Y�Y=��@v���(F��.ǫµr��[ڷ����;��jo����f�{� �x8膌f�|k����]���&v)@J,��܁���HU90���c��u�.Lũ^\���Y���\'*�Nr{R��Ŋ��#d�Et�ʎ^6ͮ�q��5.ܩMk�2���c�3��hCVL�D΁^��
X�����9�:���h]gp���&0�ԙ�)IѴ�"���-C=�X�$!����P�Wӿb_*�Z7���<�t�z)<���u�'M�Oh�S��r��n���).pR��eu�]���[�Ff8]��:�lz�8y�?�׻g#�<!��=����Q!Lf��T�$.7���2�+�����AW�$t@��͇*�5��5�s���j���_�5�v2Y�gӽ9�8�o%�}4|�C>�>t��0Ql�����B�ۺ�/���ǎ�DM䢅9k�0뀋;}t�vԓ�sܲ���ewI�"�IF�=�U��RO�te_l�E�8R�H�3f*]�q:g�6�V�:mŞ4��r�}^8}j��;.p�����rZ�"Z|�S�lD�~��s7= �	:�8�duJ��l�ƑL\_��x�nlS������V�a�bh��}��zC+AN��<k韔DmPs��f'34�[�	-
����h��O����/6���H0�����o	�����e��$Ƒ\r�֞T��J6v��X��� S����ҷ�;}�[��ݣ2r���r�bD�-��!Y"�i�ܣ�P�S��PH"��¬�/��3�Re�@(D���4�ɰ�}����l���r�eD6�pw�is;w�ʺ�x�9!��,�*yI"����|G���w��DX�,�,��G�N��])���x{��X�+�%bC��ر��o����.�T�	��,��Z�pT�|)3�C�Uk��J��t"��N٪�Ɯ�l����^E>�Iױ���Ь%�Q��>�ߝT�H���y��ߟ���[�<\�B�U�{���n���I�[4c0��J���Q}N 
�oy���oey�;^�kv���mxe���Z�^���M�O+A{^~�����~k�@�Q�F�i�:�E�ϴ*�Ј�YZ��{�k��'���6\Y$]�Av��4�ARwaҿG�2����/����e߄�E��k�702pmpΨ�����d˹���+U
�-4�p[o/L3�
�Ŗ�'��]]��CoJ���.�'�E�#Z����Y���BJ=]�����L=MK��v�^N�������v��b�\re�\�fP��/|QϹ�zy°u*�@R��1�G��'�)ޠ��1і�9����8�f�O�T�t>mP&�T�rwս��[�N�nN�l��Ȧ#6V5S�U	�Ll�&g��	�\ξ��|=qo��%���sqI�ս~+ܮl4���bc�w䘞ny�C��V�*�~\�z��Ց�f�Ϻ�8���ms'�nJJ�<\�#+L�W[��}��jh��W1��iҸ���j�힨�(m�kO;��1"��H9ǫ�q=t��G��.釰��׆WY�:L���������n�	aG�+�Յ���Pz�9����<�}�j�NfkQ+
���'G�J���*�C.x����Z���v�W����b{�{�rp�j�]|��ǱJ��	�c63�O�WY�][��-�G��
l3��묅����\��smu�o$p����le����Ҡ����u�W�޶������ݾ��N�\]��+���
heB�X�2ۛ�ǜ1��vK<wr�z0��qYd��N[�_e�,��}�����O9�~�W#�ӏi�H�pAɳ=�5��9�(�}*�j��Y���;k���&ś�>Y�����1g}ZL�����g��]�zsf�ڋ���R7��6bS)j7,U��}��tj��.p�B� ��XO��q{�R\�����׼����r�����Yҕd)	�*�e�������9�<1.~8��͏M�P�'p�Q�[D(6P���r�L�;�U���c&���|'��M��B{����P�(��Y�����7�5O(T��J���N��\��t���S�}�gZ�o����&�=;>e�{r���,{�W�L����5��L���n-z��v�meZ�V\�Ȍ�%�F�j�]�c��왇 ts<���:��{�2���}��mp�zōyi�{ts4�s���*v�v�9+{�s���t���G_r������ED��[\o�3��Q���7�fvm�u��#�nN���d�6�3Ȟ�8Q�uZN�z�3�����D�:��w�;�����b2S�0pP��.Gv\�3#�ˡ�Ж��'��8]����v�P�(H�B}� �P�7���WZ�RU���-�����޻#�7�����:>Z]*Y��;د��z�����O���E�J��Aɸ;��5zc[.�I2��B����|Jșڋ�oKSj������
�[g�x9a�Ã����>���=�<���zZ�P��zC��5�5\���&*6[}Y�(by��O���Ό�̪�-�;��D�� �πs�9������V�gdz��oZ�V�v���Z�e��k�������c���Ǖ�M��P����2�n�����g���ٺ=W���z�[똍`��f�Ah��e`���)n�ދF�ں?�֧���o�ƽ���*�p�{���O���n?\}ӬuD��a7p��X1g#������.4*+��-�7�8se��1��)��w�uZy\)�9�P/���19����:����[pf�a��M�H��6�ၵw=uou�U^�!D��L�����w���=K$�T�
b3���
Y���f���q�{^$�Fi�4U0���y������~ɴ�f�i��O�"Z�=��^�l�����T���&�C�v����F��{�E4g�s�s;�m 0�!�oPp��Se�M.�ou;*$���Cc������jF�w������Ƅ]C+7��k�gB.%C�G(4/Y��b���g�+���>rg��>!i2���镔����ls����q7r����)�L��e���pS&_1����g��C�6���x������	�f����^tUDU���j�v�ll�CD�d�_|�!k�\�]���ᠾGD��Z�Z�\�ܜ�<�&xPw�mE �M�� IUCkx��[.�n4��eP�/�vPJ�>-�i��R�n���U^��(�a �Ox�>=����B�V����q�S�{Wc�S�8,��\/*i�*�{�1�튽Ȭaqs�t���AF�44�8ͪ��v�p��1}��x�hp���q��Q\�w'���ݣ�lm*��\ue;T�eҒ���k&^�b-��8���օ��1�/:M�"����[vD��3�o�R5x�<����-��V��ˑ��%�n�k�]��t��s�����Ev]#I��޽�>m���R��7����]�n��Yo�a ᫾�ڥ���o0e-�!�v�غ���Z��Q��ޜ7杋�XM*�\�8RVV�]�+��*e`������	r:�� ����,6�7�*�oS�q.8���e�6�� $s�Vo(��&�{�����,��Q��,��q_e �ڻ.����u�w�5^�B�+�Cꓺ�|RU<�yv����!%m�e`Y(:]�x�e�gX%��,�iY=W�v�c��7TO7.Cճ�f؜�!
�uKm�������������pŽU���C!f粊a���C�<���a�J{�腼�>�5oPĎ����)�{����{���aS<|Q�-���;�GI�B�R�]g*t땥8��e����QB���X��4�V<K�>
�˨ra���b��Co����Uoy�����^g�S�.����Vy�]��V��8*��S�T���E��G��t�����ne�>y�9�A\�o&��+
u.%t��I�B�;��j�%����2acq��f�)f>����[y5K�KL����G}oF�6-N��\��[z���0�Y	��19����1��
�e�J{;W�C�=5���N}eerµ��⺅蝍$���wuu��K��un,A\�V�J&�jw�Q�N:�%L��-�lfͅrt�o5G�0^9�i���f-�]ut��d�5�a4�nR�{�q$�A�[� L4.r&��U��pٕ��&�]��
4�4�.�o٬�ĴV�C��=PUwИp�y��QL���>rA����I���)�xğ2Τw�V����/��/���̺T�̓9�'[S tkNv��=0��*ĴC\.��)ٷ�$�TX�k)���y���4R�`���2:r��D�\>�ߵu.��Z�ĵ�1rEL,)���1�l`(�ĴL)�A2�X��2ؠ�A��Lq%dU1�F�Zزb�"���d�$,��
ԅaUX""��`���m+cP�+Tb�ET��*�\�q�*��ʕ#
4@���F*$QH���U���(�
(�E�b�TA��TQjJ�1��(1X��Rc�1PVVEXJ���Q�K�m+Qb�-�b�TX��K\VC"�Sł��+b��VH�Q���R�2���e��"�fQEA��XTDX�1��`�QEX�X��1Ub��� �`�b�����",E����	�ȫQ2Ղ\lAUA`�b�X�.Z�*�*�(���DD (DAb�*�V,��"�E�Qt9Vv�I44�^ð�,�I��ig�%3n%��U�k�v�Q�����ϸ��^;rI��d��1p��ȸ�[�c�ya'+{�-�:.�k�J}t�/�u�㌬'f�ztmy�o�x霶?5�"We+�hN'z�Uj/��8q�:����ۡ�\��by�r���+z��Ltsv���gJL��4���ዦ�l��<�2�s�v5��w=y7ԓp�J���'�,%M{o������Ej-����)g�{����O6)&�e9�*9��
W�+��v�nO\�Y���J�9��u9�B2�ԙ�nB�3���SO:+�c�r�8�\�9#͸�����py�OU����B��m&�;l
a��!�����������j�Sy�o�\��*lNqۥ/�Dm(9V����"m9T��Z�����}w�5Ѕ�p�9t�*�jjx�ׅ+������=k0e(r�94&��׆܈��\dn!}�K�c,k���#�k�&�4gn�k5�o��J�wΦ�[��㹑�w5�
7�I�1&�gM�GK��(\1��q=j:��ѷj�fUL�]]�,�l\��7o�J�$DN���i]��[�(=u�;>7��鞑9.��gI^.���R���'�q���N�����7��I:%@�w~�_{�C����=g�Gj/1�܇e��{�Ɍ����O�=�o�A��#z(���nUCT�������q�D����u��q�ꇔ��<�s���{�ûsV��0����-xǕ������	ShFv�V�h3z�-��C�~u=+����[m&�(���8J�p��V��O�v�{K�w�j`^*x�sޯb׎�N��7
�:R����Xcj�y��En�Ng�~5)�<���y���r��J���"�JoTSܞz��ҏ���յb`U����tO�!y����ua�ZKۣW�(��=�Ց�K+Q)�enl��nCS��Z�Jת^�����z,*��VQ�G��߳ۘ����Y��!ݨ7�b���v�d�RE���r���uG�	�e`��Bد&;d���k�qn'�4����<�ux��u�J����tB��gV��+L'�Խ��[�!9��hJdl^���>Ȼi�j������ry�Ba8Vn�֊�/���8j�5
�n_�WP�ڠ!e��U�W.u�s�|�h��b�0�۞���R�+��$g�1BҊ�r&� Ү�I�j#���B
�+�vYJv�XI���-�Q�u�f���'v�j�Y+�Q�/�հҸ(8�4��z�8�21"k q�"7��o��s���qu�#�\b���M��D��<�o��%����O>��=v΂�쓎�OL{��V����y>����u#KveDu+�B���e�3{1.��=���J�ֺ���91�2�c�fA��ԡE��ʸ��vfE�T,�
/�����vfupΫ���Ysu׏�{�^Q��:��sz��@��I���G\���L"� ��5�yq�IʁK�ݵ�����=�<����|}ov	.>������Wkh�i5tJe��B�����'�md������eK�t!M�-�ORS�w�E(���e$��1���R�~>��鲯^k{�y���r���gu[�|'�OP���b�����}=TJ�N�E�c����u��Nd��ϸS�~56�y�i�T�J9�SNa��E5��K��B�"y�Vl|��V���s܇�cK��g"|ٞ�=�%��X�!�!����p$t����7fN�D��H��o!永"��;�s�T�r�G2�Ďn:����!�nNt��{OS6r��Y�Y���R19�*zt�(���.v�Mk+2����m���{��B#.�
�t1lF;�n����zv�]p^�M��Nbe�S׶�9[b�� Yr���!��[ }y�o�N�J#^m$�ݫG��4���՜tfv��+�M���0#��}P��k0���q���Ӆe٢V��Fs�!�w�YZ��Z.V��Rs�jc�1څ�IP������rz�z��T&yR�,�)�FX��Ӣ~;�3Y[�8����B����ANĈ���s>�-�콃�.j�0o�z�K�3O¬@s��9��ߟ�+�9\vh�,�f�C��������o���3�7:P&I��>�|�>	�Q�iݽ��;�TO[{:�δ���o���=�D����{-�ܹ���l����1��T�DuF��Z<��T�3R�����l�ؓnT����O��:z;�{Y������p�����̨��#_�/AkǅzI�z	�jҠ��g�H�m��wn&mkm y���X����e���gR����I���%V������eo��۝=FLҽ^�r͊I�)ȥ*9��
�c�%݀�ѡ�OP#˦gŨ��*���DQ�7�������饎q.�o�T9uý��sR�l������\��B1:U��흦S�-ζ�"���Xrd˦�S:�
�ջQ�䥄E�ԩ�I����_��>G��NuT&gɍI�V�v�=���qN�A&��u�r��.��N7�f���}/D�:�t����b/;o��U<"�ځ>r��e����Y��'�&5��{�p�*��q>\ml�`�#ۯ)}B#vu`<a���WBWOd^/`	�
�lݣ��\o1��a3�"�q=t��=gj�Ve3YVTe��mX!��Һ�]+>u$��7}ޥ�߽���X�C���B��{aݪ�G�K�J%b؜x�Ï&�^�<ҕ=9u��W��W��Z�Cb���P��os����Oo���t<S2C��L�>>aǲ��;ޜ��-j��<x�cEN{kC�m.��A��$��9�U�����p�})�দ�ͫʾ~�h���;`�~Wl`�$٨1ڢ��B9!�C��u(�o��>~ܺ\N��[�;%mo�
��n�#\�Y6�9 �xp�ޔi=5Q
�WܒK���$Ի��V�Y&��<O,�� ��#��X���)}�������8�S��[�gF	ͺ������]�å��=}6����O�n��T-)3�{F�̞�R�T�K���1rv�E,U�{ص�;}<�q��H�EK9ӗ�[�V뷩,��'����f��d�tތOE�]�3.�!v�u9��w�{+���yʼ�sN�>W<�e`���m$@�=^Y�>�;�9���߅v�VDj|yי*����
�6w��a����f�%S�n%�=�G���)2'�d��^䫫98��ZP�yu���4�ZÒ��9!#=N9�t�N��*WP��+*�«��UK�94��r����e��-���:N�+Iڠ�3L�����[s׈���T�}P2[�B8$N�*#�Ee���D��;7Y�	�$T���v�ֵ�,YU<sB�����n���'���$r���N�\�;\ta𜊯����ܬp�K����A���r�&�]jc�6�P7G$�,��}2���\���2�9m��}����������R�YKeb�s�:��M���=Z���͕.���.=�?csj�����Ss�Zs�Ϧ7�C,���z,�!�gx����&��oD����p�-�<͵��S����f/0�Z��%�i���j���\K-u9U	�L^��/��|��r;7(5�:�P�S
���r��f�Vc�n!.~�BEj�*:C�՜���}�OFtW�Gd�˜����Q�r-v׫��m�\���|�wxS���m���-�y=6R�W�L7)�H�֘������Uu�sӏ�czT*j��I����9��k����:�r��#���*/����_yRV�pn��]���.���"G6�1�w=b�� �W`�h)/�A��"T�Rٽ���9h^�1�Y*f�K;b�'����f�Ċ���jb�Rs��R'D�`�c3t��MR�-�߳Vۘ�sJpܚ�ox����+%r92]Z�v�5Xe�w+�-��i=bT�4��_L�|eT����BPX�	9[�#�u8�v]~�*b�N�R�4\�Ō���T�r��ԔĎn:�luv��ס�{�D�Fұ)�gf��>���=�	ǔu�Ds�'I6�=Jʉ�Uе�cUDe�ʼu�b'���8!�ݜ�"V�W��k��pv��\O])=e�7+���Z{5	�� ��o2�D�=P�����BXO��%���^�{qמ��wɩ����ԩ���OP��MG��b�A\^Ѕ���f.M��Z*n�Q��s��~�@�'C2�� ��	�o�H�/onN]�_erɝ=\ڤ�7���I����54I�n��;��EM�`v�Q}����Bw��y�Z�ڬ���B�q3A>�r�����͔r�1r�a�Թ�Z��g{\���_h�붣'xi�]ᗛ)u¯22-d^�\��9KCp]��������/rh5��*�p��S6�2�)���nM��u�v(1e��}�ͽ�6��t�NSwڌ��
���=�4v�=��Q�sY�ܵAK�'6��Z�mS�y׷s\Z��:R�
A��@�3�wp�,]4���9�KMK���ͯ5����o�|�p��R�'�H4��ML�T�|�Z��iZqV�q��=x��5���U�(�׻Z3��|]�Ow�zi^�<�q�Μ2��&u�Q׼*�Mk��V9��K���e���}��E��r���JG}q������n���:Ș�#6N�#;��9]�҇g���L-@{�gO�/��v���k�d{@-�U�񆷽Ѐ��W��=�S�2Cc31;��W�>�.Gv��y{B��
��Nm��	�!��p�&Q�YJ�nҼ֮����?1�G����Z��j���HH��G�⠪����aPG{�e��-��mb��Ѣ؟O�r��[]J5��Ʊ���!��[��wG]�.�-mA��(���RI�J�]�}S<q�����~��\2�U�c�cx�a���1�5߫c;o�!�e̓~��о�*�?`���͸s�}�^�EPG�vTU~��FD���o���)�A��p�Cf��g��v|�f��!G?5PG_�e~�.��~�{�D�jCF?���f���͢���j���<�������8_��J� �<JUf��@���7=�sg���UnCf^I�E��
�-Z�7reӆ��\�zTA�S0J�s���ޣ���F���		g��=<�谿��[��Z=��ӵ�7�҂�#��Z&��}i�?P��? �FW�qħQ�)��xqTR��պ�v��ܒyWkj�̍�s��#����Ϙ���f���W�'�!呄"� Dl���AT�>�ތ:�=�<e4�V���p�{]�L
q0��<l� �����HFn6$_Q�4 Dc84"�G[���Scd��J�0��l6\� ��U'�B�/��\Tذz:�V��'X��#R�>�)	�S.��4��K򁠺`kɀb�U�H��Q���+D�8��iZ��:E�����ZUh1��0�!�)��6Ae�0ӥ��#�İ�4�q%B�6������>g����%�Uv���^��~��}@mO�����Q�]���õ���#�t�u���n��SXx��8��C�ܐ���<WOI����»$TU�#�,�0-�Ve�Z�D�����sN$�����ˌ-.�ij{��N$G�!��۔۠���ܑN$2�N]�