BZh91AY&SY�$���߀@p���"� ����bJ�@         (    }| QJ�ͭ*B�$I
AAD%M�)3���`��4+cF��DU�(h��()L�hP��P
֩�l�_`B��H�"�U*�PTD�PJ����!$��ER�
)EP*ET�@p A@ ,��D� 0"��]�q�R��*	0ےID	��U
*J(���HH�UDQT(�RIE��EP �G�RQ@ �/|�TE���3;�ˢҖ
��_^=$*�԰
҉��EUhf�� ��@v�sT;`�8UJIE��">})J 7{��J����}�UJ�IEw���<��QJ��=�J�P�ty���*��7�5�PO9Y��R�x>��*UT�T�=� �˯�y�O|���(P����U��Pj��HV<�RT w����jR��y�J(T�z�����UTU)G�;�UB��ҫ���/�¥I<���ﱡ�U���V��47�7����������t(_m�m����z���)�Q*�$��*��|)C�խy��o��B�V�9��� )��}�>�J^����>�_<��ϡ�������Uyþ�D�B��q@ER�ϻ�R������m*4�ATiB�J��I 
�P}�$ �!�(
>�s��-5*����U*���R�B��E�wYT�Z���T�F���lY
�Ww�������\޻�U�2��u����ik\�P@"�
�Ek�ԩ@z��m��u�U:�Xw:���T����	Pw�.�*�@�Wv�`�wfˀ��ntX���uW�z �%J�N&*@�Ba>J)@ �<> ��w
�V���� �l���s.��N�@�a� 7$�cusv�Yv�T��� WYP�w�JT����>� 4�؎: ��0�Ўw�u�@ n�� �s  Օ� 9;��('(:�U1�����|���r>+���r3�4	рӠ9� S7l�  ���� ���@t����� �^��
�*����ѨT��I) ��@=LP�h� �F���M�  ����ٷ �t�`:P��]����        �   a��d�*L�� 20� D����Fa1�`Mj�� ��P ��h 2@L!R�Q�     ��J�  ��L 7�SjC�)a4S�MO�=z�=L&���??O�~��~����O_�V~��[F�`�5{ƻ;�;��9���I$����@��$A>�$�?s�r�I$�L�?��?��g�??�( *��UW��� *�l��[��������c����cLXŘ��b�.*�bɋ�b�,��b�K��œ1S1d�J�������������,Ŏ�1c1S1c1dŌY*☩�b�,b����b�Lu��LX�LXœ1S1X��b�*b�,����������qf,�)��ŌX�J�����������������&-XŌX�LXœ1S1R�*b�)���������f,b�1dŌTŌTŌTŌZ�Xœ1S1S1SLY1d��T�S1S1S1c1SVbɋ�������T�LT��ɋ*b�*b�,����qqS��Y1c1S1c1S�������������:T�LY'�LXŌX�LXŜV,t���������S��XŌTŌS1S*�,bɋ�������U1dŌY1LY1S1c1SqX���,����������b�/K&,b�ŌT�LXŌ������Y:TŌT�LTœ1S1S1gLX�S1S1S1dŌY1c1dŘ�U�1S1S1dœ1d�t�X�N,���&*b�,����b�Ҧ*b�,��,��������*qf,��LT�LSLX�LT�LZ��&,b�,b�,b�,bʬX�LXœ1SLX�LT�qS8���b�,���&*qqS�LT�LT�LTœ1SLt�1d�N,�����b�+LT�:��b�ELT�b�,���&,���LT�LY1SLTœ1d�LY*�Ɋ���&,b�cLX�LYœ:T�LT�LY1cLTŘ���&*b�,b�*b�,���:Y���LY1S1dŌTŌXŒ��LXŌXŌT�LT�J���������������T�N�1LXœ�LX�N.,t��b�*b�����Œ��b��b�-XŒb���T�LS1c1S8�:S1c1LTŌWb�J��,b�,b�,b�,b�LX�1c1LTŌTȱ�&,b�,bɋ������f*b�1c1c1c��TŎ*b�*b�*b�*b�:XŌTŌXœ�LV,������&)������U����,b�,b��U1S�LTŎ,���������'K����LTŌX�LX�LXŘ��b�*b�,b�,bɋ1d�&)�&,b�*b�,��bʩ������������,���'�LS1LXŝ*b�*qd���1S�b����LRb��:Y�"1I�PŒF,Hŉ�T���1d&*CBb�t���H�IT��ŉ�C$b��Db�1d��Db�I�!&,��HbȌY!� �DdY�Œ�#!��Db�!�CE��<aG0��
>0�Œ�#Hb�1Db�ń�$�!��!�C�#$b�1I���b�1aQ��Y���$b�1Bb�Œ�TI�$b�1RF(LT&(LX��$�T��HŒ&*IT1H��LX��!1d&*	�"1bI�HŒF(�
�&,�1b&,�ň��"b�LT��1Bb�1b&*"b�"b�:Q�1dI1d�1Q��X&*#I�:Q&,'Hb�LXF,H�Hb�1Q�#I��RI�ňb�1DbȌRF*I������&,t�,b�*b�*b�*b�,��,���Y1c1S1S1d��,b�,b�,b�,b�)�VLSI���LTŒb�,�I�'K1LS�$�1LX�1c�ɋ�ŌXŌT�1S1Sb�V1c1c1c�LS+F,b�*b���b�,b�����b�:XŌT�1SŌT�LZ������������b�*qLY1LTŌTŌX�LT�N��N,b�)������t�1c���������LTŌY��b�,b�)�������:�X�S1c1c1c8�Q��)�&)������1d�������b�,b�,�qc1c1S�VO�'U��|������2��W<7$��߶��Ri�yUv��Mܹ�6��� �fG��2�	Hl�m����^��W.@�8l�*����Pقˎ�GiwO&àk�U9�_�\sr�`�;�bF�!���1�QC4�jț���1��f�ƕ�M�3U�A�y�n�C5��Rj��W{��	o;KX�{V�j-��:�9��5�D{r�e�V\�D�;�c��ʏ0շ_P2�*�����Iyi7�Y�(#��0`�9CN�~D�v�Ux.�ͥX�v�3m�3$�&mڙ���JXV�x��T��Clb�Fhj�n$[�][����BX���I�>���4ʴ�V�aR�m\�'J���f��\�R	��Dd7#�Ksq�K�K*(r/JX�9�'�j���P��֡wrhVY	ML���OnSh��.�ٺ�s3e�Sn�ʅ�	шn��|f�kci��2I%ne��!�\V?n����c��b^�B\��,�e����-(VhX]GKC�Km���U�#/7E��ML�ǖ��H~����R��p�ma/1B�^چ$$�*�^��)u��u�&��v-����[W*%{PT�n��\'�Y���@������^���OX&�d��������j��/n��0�,Z*�(� QL�������0�.9�I&�+��U�{�L+�C�Es���۩���ͫn�,�^��cDʄ�)�fݕk%�U⹳�Cэ�N'��1nZ!��f��|�Y�7�T�ԥNM�W�Qm�%vD���1�X��M�am�t%Vx�Iz��h�p��Lcot�í&E�ŉ�Z�噁�j#]�b��6Xf�+2�
CWsYݡ�lHm��ՃI�7�1j̓ڒ�E�T�*����omS�zt�����NQy���gN�Xhڎn[����QAQ5j]`�үa��t�V�ۂݕ4e��̭�Yzֱh�r�rJk6��4�rPU�5�L`x�X5L �r��7��)�j�v9%�33\��6��j�&� V�%��7*��de�(���k�th�MGPS4��n�������	�[7��up��B�����QU�P�aY
��jO="��WO�tT���.��lX�PTW#��1�f�%�P��Z����U@a����p�_^�U��[������4ȃj
e<�J�5���EMm�Ʀ�l��k3�e�Y�#w�*�R�wws��+D�!���Ʌ���֧��rrx*�0XL����.����*{�K�e�8�^�j�(�9��܍��?+�Ea���b�4�I�UinR-k�N]�Fm`Y�#UP@�Kq�ͨ]Uճ�q'Ln���s.h�-,5�a��,Goc5�CCA�A�p�խG�1iq	E�{0��d���X r`h�@F�(cڕ��0�m�#��M�(��;HJ���u�-zQ�
EEa�b���b�Ɇ�\�ʒU�{:�
����ڹb`�-��k)�Yk)�e�N�cj�`O5V�n��j�6@+#b��N�ABe�{�n��#)6��`���lY��8#5�2l�j��ZS4B�G�1�ݐc���`�9��;�j��9&�ľ��ÎB�����Vǵ����Uu �U�M�2T)/JoM����CS1�����Ц�f��:E:�]e�4d�|GoT&�v	��J�^X��gI7�N��m���Of��r
	���׶nR��n&캎\�ۼ�W�h������蓟sHa*�-kT���ǴMKN%WR�Լ���u�6�=c(lzKyku=�:QON֌��"�f�	M'j���VȨ�xg]�-��tUj�1���UH�ЛJ�(,�p0��5�$ۼS*�?O1��B� �;��� t/I9�ޕZ%�k�ji��[���ބ��b�D�Լ4��)�Riߜ%fdX7UN�Lɕ�4r��ze��ĚP��H��f�Σ	�b8�/�Q	e�n�*���{"&U�[u{������43��7qڤ��wSAo!��fL�,K��ʙB���GCqe��#uD��7�<t\�4�N��ie�+.lw)��Yd�Uj���
2I�Xs@7n���[f�1*�"Z\zk��ne�m0�k9�C�2�44:���{��)��͂�E��fe����[��s�X�Htb�6<�>m��ƘeujV�Ma��������M�mm��F�%�c����k0�ɛU���(HhL�YO� �"U�Gr�`�2�WB�Kة��7�����t"�3��K�
R]l2��fGn�[�t�"b���A�**�uN�V�v���3.�SO�Pou2qM2�֑���V��ݺ��a®طkP@�fM��z�j�e�:��T��.��P�7�m�s{�n5�&�L�x�(�R���)�݂�&�*�;��V���+�PVԏs�[��v7��vmR��I2C7�c��{͛m���i�8O$9�f<���1�e����7���w����ki_���{,����,��P�ڵ���ybڽ̡$�4ǚܴ��jY��XP��q��h<"�a�Y��~qV���ӊ��tS��[C0Ô*��x���r�w��v����/a<ĝY����n�����m,ٳP��ˢr�Ňp�Н#�n��mH�M��7�������`5�jRvk$�LY�p4�{�Y��w
d��0J��0�ZǸ,<��0j,����������9c"�PM�&��5D�Z7q�gw�/�i���h�lau1�E�ъ�:��$�U�5��XR�"��Ʉ�	��n3i�k�(t/o$�0R5('��$��\�k@۷2�-�޼��k0kĚUX��M��Y"��E�[����0ʨ@i�U�y�32�[�af�hةJ�2g1�-��ag�kl�e[��Lriչ�K*ln���W�T�$L�x&�%݇�"���e�W���ij�S2C��0�IS��J��朥��Eypl��a��YV�/(��

U/*�b���B�n8&˅�>�G��^��rXc������9�ťR�����+u���Τ�$PՊ�-M�j�@�
)wS̷LřpMI����N��F�c"���l��E,����1ɯ	��E�,<Ę� F�E �ʧe=�8����ܼ��jT�i*�:77V]�i�Nd����.��-^��b�.�R�1�E�w6f*l�>N���`F��N��F2��ae8��+e[w�5+�6�ȥ�Փ��i�[D�ǁQ�/Q�(��:̋�ۢU;�U*��H��x"�b�ՠڴ�c�)wm��̍�T��2)^Yٔ�׮����I�cЋ�6�/�Y��V� 6n��&Ey��ٱQ�v�OAk1<˺ZN���e;{-T��rͥ��-Jt����V�a
�&@�KL�T�Y�W���MC��a�Ws(�b;�K8E��5��%���b)�{z#�*���n�V��N,�KE^�.��.�T�qn���!77��+"Z��7��ŲfD��,:��L4E��k�5���b��;QVۧ`�����c:U`�����Q���C<@z�5F��I����C�)d�K
�m����*��"�iu4H#�c��6V�q�8����ш�2�VͣAL�׭]̶
�~����2+v��gn�-�(fKn�����j50'X�U���r�,u��J�v��b�;
��:�,���J��Аn���/�@z�Pb�t�%��nf��6��'rn�q�Y�o)&"ȰPb����:dx��m˼�Xq�V��	�Ò�aaN5a�sv�6-fM��4bR���,
:�731�M��� ���.����:��������U��"(��{�P{PӷY-��	VPU&@��\���sP6�eg����`B�R��F�v�G(�V���rD�ާB�MR����E��+v��oSR�Ҙ٤��n��b�زdY�D�&[����a�m�Xa`?@��	d�nc;YY�C�V�j�(Z������k���S�@�LM�a�Wta����5�e�D)x/b�%��˨�ш" ��1L�W��I�r����M^�-82�9
I�Xd�`�]�m�B��Y7w"n��.��Vv]��̰ud1��t�V$�Ƚ�����Ù�����2�m(s6�hI���m:H-�GnJ�ݓ(MY�Z���G{��d�}Ѫ�������j�ud��L�ͻ�1d���f�ٛ����Ҡ��nM!�xsm�*$��nS6�ɆnM&�����W�5�HvS�k94��)�w@�Y1#N8U��m��`��b��.�F��?^6�+�/�i��׳X{�j��v�����Z����Þ5)���m�B��%�,eR	j�.C����fL�J�i5ga��m��L�6�~���[nLv2�R����ʲ1�n �9�e�(�h�.V7y�G�[H�o���ڢ�.���7���1����70�p��m���ۭT���SZ����b&��*���V����E��f��V��~��`��CmD�mv���΋+��V:�&��<p%�yz�,���ͣwGT���v�*zr�C$�[r�!�]En���cQ,�eUJq�ٵ���5�.�4���.Y'�[Q�BT&����,e�֚%����ՙ
`�~il�s��h_��,��{�TT��������ls\��i�[*B�rq���אx�����A�a[�*jI�[&S]i�R2]�,��w#���)gj�ose��o�{x����c9���z�ZF�����GqAwy���enՉ6�,as5���1�Qt�[�%�#��XV!Q5�u�[W���x��9���E��XAH��)�W���D��ħ���f�%�ak%芑�CybO&��a�U�1�b�$�nm�i2��`;L:�9Vѹ�̩�;Ym,Z�70�X�:3r��Y�����2���G���7`����m8T��B*�}�D�:��X9Yw��WX�k�S�����GZ�K]YyJ�WIU�iǩ��)i�2��*�*	YS�KT7�(��,�!�!)L��^����7W/�v"=#t4cz/0C!���(��d�Q��[u����u����׶-����k9k�%5�V������3N�LI&��������f�zjsj=x��z�s2ۓ2���5=������� ����h�*R��$.�,�b#�k�2�V��1���ˌ�ŦڍHYܠ�*�<�
�	F��s4z�R��C`߶ɔ@�z�6f���wS1-�í�(M���l7
:Z�Z�
Ӵ�ۧ�R&�\�7�[ʴ̉6@���ƍ%\R�ܱZ�G�J��y�J�t6���`��V(�l-�1ɽB��,Y�[KQ�r����fۑҧNk�r�A'Q8��2J��0$H�:h�toVR�t4�i�{��Q�W5�f�l����n�ÈѪF�dح����x��1�Z�W�q��9�p�c[i&!n-�[�Xg�s,�����ѴERI���1��Pnպ��c�T�ӫ�������˧�ݡ�2P�}�r�E�~}�[��) yo�*�R�K��䆚����w."	�鞦�\�-�<R2 N�2ym��Jh'�`g��X��ض���R�α��gj�rQ�km4�A���WNFf��6i��;��d����U�y9��=t�ш&okJ��*�H�Ĉ�(g37N>E�����h4֪�S����A�"��H �r��LG�M)֛Z���IF�ĝ�(N�w57Ƣ@�	n�UU�Zm6Z�������&~p]��+��N�n�T	��L��jzdDт���2�kZ	m�Ŗ��A�ppf_;���h-/�%��u隷D��W��=���6O�ݩ�Le�BȻY��lS��:���`���G%"6����K�cQ RRku����� *KS.!U�u`V�e�·t�\t��>o��*@bI,48]]Dun!F��멠R�r�)]�NP�7I���j���igQ�ƙ
�e	lc�*��,E��c3[7t�����hY$�J�Q�Z�*�����F��w�c�%b`�׻i=��D�Vӹ!�R�6�AU�l�F��8j����õ�-�j�I4�+'t�h{�
ɤ���>[0��fP+�����V��Ne��4)�j�[Z�4A]Q(c�K8�MJ��-�h�k��;���xz�P�o%�v�Af�d�B��u�,�ĚI����[�K�z.�5���W0�*��ז�{ӧ�jaE*��]b�[�7�#JLC��J\��֕�q.�N��!�N%];p��p�w{4�-��EE@�Dd����/����ƛ�(�G*��B�˚���L�y����b���Toh�69�Z���e�X�.n�-[��X"G�J-�)dQ2��Y���l��I�k�Y�!N4,�Sj��-:zV�Kr�B�5�G+2RA�ō��B�äH�M4�$�\�!ڗ)�ՎA̻Ք;% �J�!�!HG�Xz��'r6��8�@��2�B��M����!5�*�r+�P�Vy�� ��|��J�*(��_)I�H���D������$͎����M�j�1���"�A�w�.�ٷ�'+h��Uj��&R,24�܀���(�W-���5;�ԱAn��bYa��c)�E�e�5��HY��@���VbX�/��t�J#-nιچ�-�qY�ᴍ,�A1���q��b]TGR�
5k��P#�ҕ��!�B��7�2������H(����^�̢�Iĩ���k���{�f�;n�@���-�r�٦V�@���Cy���em��k�.Al��5��z�ّtG����㵥h���i$��S"�8+�,�t;�����V��������Xt/_�~7�@�?D�)�������R�2n<�"�����7y��o�f���m6��]0s��6o��T�_0Y��=�a�\��mu�X�6���ov� ںC�rf��E�V�u��N�����S�޶v����������3�Ty79������7��	��ַeF"�ٰ��C��ag>U����Bv�,n*�e-}5�>�ҳr뀦ƍ��FNVwzJ�o>z9���!�	���N�w9m�p��WY/�t�zw�M����]����� ����VL���Ը,nss����z�6����ē-��7���7�J���Ne̜����v���O.*[j�5!��;U�t�)�����'����f���U��e꾰�t^���F2�RC�OS��^A-��ל�㋆J��1(�B���:�Z-)�K���Bb�V�$�ՠئ��Q0m�ʝ�;��Z��S	����U�-�QL�dC�_v�m�Z�z�0v3��3���N�$�!mԷ�ɩ(7�Q�u��6-^���>46w���f����y+��!�=}���6�Y��FW'y��tU�;��:��g��<W7����Js�Q�i�UUq���S��v�$�-����s�dtF��B�Q@�do3]�7���,uL�J_LP�x�Ls;�=�8�G��U�Z�AL��v79����l�iQ_}�����)�H���8Q��6����y�wn��}x:�.�˪��Z��wN��	�b����9���sǅ`�֘���3���5�����S�"�*{����AQf�!�^<cs���E�5���9A����,ct�WV���S��}¥��ͼf<�w�>I�XJ}�s>˔���F @���K\m�k��E-pL��X��4����W��-��Nvj�4ҕ+}ӅmgC�X��t��OGI]~s���$=�������C�u�S����}�W=�>�<2�@\�8,�v�>�S��X��s�1v�E��X���76�Zi��P^�U��jaGs��(E��%�@���#a�ݝ�n��񾡵��c$�����t�C��m��G���6VZ�'']����3s@sN.�SX���q���3V���ד"�iU9'�1L���{X�U���M�:k�y���*�615;��C�b�����q�3�U�E�T�=ܶnT�jNT��\���<��o�YܣÍ��9�I���n�@����:˅r����2�p�vtG�����LN!-���G���9��I��2q�����fww���F���f�Үkk�
��4j�}��=�I�H���N�|�r[6�:�\�J���z��KYӶ̊�F�T]�t��;��uc,Q�h*wN�{8����:��q�$�s�����ؘO��c�o��io�.:'�1Z;��=��I*+o��g�*����QY��_���Q�g'�[HHo%��r�q�����ђز�<4��[��8gf���P	�Е�5�%q�R����ȣ�!J*�RD����]9{�s���=�/U���*���Il������w[z0�8�Rc��[�u�\�6����P�u�
'ƽ����:��[����莲�D���]�z�b������B�N�¸#�I��:�Wݐ���}���
W�9�!nkzo�/e^tTk5���H�m�ϐ̬I�k��S��J���s���C�˵[yצ�Z��7��M�U2�����v�mM��t��(f*�'wE�m.U�g#|#��r��WU�F��t�K���
��ɾW��ĠO+��,�+����s�M���(4H"p���3�3P����-����+��V4�έ��.��͜�nZ;|Nr��{����H�ܚ^��jWx^��6��m��/v����8#E��K�_l��l�P�/7�nC�gm�.b�Nۿ����,mrҷ]��i�8���ɢ�1���{q�U+��z��b��;�H!�AeKUGt���p�.�t�v�B"�b���m�ɠ�3�U��H��൵$C2s�s�__6/3v��7�{��Vw�<5�ڑ��z�H���ə�v�T���u�<�Kf����9��w���	*V3�暛9F�����U)��^ݍ�t�����#�Ms@���)ƚ�Wy[��H9=�u��]#%gs+6H�rsT)>�;1ޱL�۵�-�x����ҼrJs����v�z�٤�ל7`o�vb��=�ūUH#x	��az��q1U{�X�o���t,P�Z�Ն�\��C␠�A�n�t�y�wGA��;�V�' k
#�K���X�壱t'�1{X6�/����^:�E������SV/�.�Ц2<W�3�s2���Ǘ���+�z�2�{���vv]n]�R;޵x�pL�֫�2�N�K��љF�wnWCn����d�{[�;VX�pn�_��M�Z�ZM0�l�d��;"��u��,oU�J�-\D�U��E.\�i�9WY��˅���X�����05�UY�U6!K4Tv�<�At���g5��+;ƄW����OY]{�Kۻ��$�}|��/<�.����y��7d�6ľ�(^�Lɠ���{&����nc�t�9���Qw�go2������F��dQD^���c���ض�WD����z�th3�l�m��s��Z�$�A�,�9�a*����ckV
���dQ�� c��PIS�+�7�5�J�{|��u�1v䓎��׀�U�/�e��,`��JL�V�O�\w|$��
z̽��2��p�9C�oRq��.�gp8��^�AG;�"6�C���i�q�-Ѻ�I�}�EvS��g���=6f�Tl�;�.î�w63o������豝�����<�4M�l��o��{N�o�x.g)p����`��9jɋXv��ʲN�*�e�Y�kw^�n��/'�O6��{yI���b��.3 w������<�n���_�؆\EB���nNdU�������ԃ䳥�������Ua�TE��+N�8\�M�Ryk{E�<�9a�1�JۗW}�n�������Z�˴Gд�2��.���YӟS�.���������4��-Ѻ�۝}.�Q�&�z	�U��_-nr�~�z�I�Y�->a[���۪�M�U�_Sa%��wr�{���d�={N�0zn�����(0�9<3�s��)Q+'XΉ>7�J,fJ��|Pf��Q���#\�5X�%����r��U�_�JX�hY{�]��#�%j`�N	L���So*�vF�e��t�Xٗ��ԫ��[�]n�)}QƠ������:��鼝-Q�vލn�b:Քբ;�4�IGU��;sjI'pq�'�p�	Wf���}"J�Q�Ԅ�4��b�(��]��d"���f�r�����{�A'�v��Wk�+�-Ӷ��^��1��|�	6Pp��/cѹ�[ϻ���9�FN���xaW���;Du�/RC��Tdݔ�b��W��lN�2�>(F1���2���d����tڄͶ�`oDx��Ɲg(���(�9s��ebD�۵��]�uj�#@�N�P��0^Gn]��]��M�[����{�_k5�W���L���y���������7u�v�a��3:��!;�W�cR��ɘ��$�*_f����5&"���}S���A��]��w�݆�o�h��f���o��9����uh�(�X ˛*����&����ᯯUP%H�A{p�x8�٭���T5���Z��ki�;���N�-�|N��ـ��}X
�}��3��ڞamUu��K�s[ԗe��j��灓ӥ������=إ�-�wn ��ƫ=wof�O72�����M�ĵ�����loB�eΡ��q��^���G{0!2��ݮ��糪^;xZ3�-�������P��ٮ��+n�$�1�+�6��*���-��M�iS���*�r�Q��0Tz:�:���;ֳO 2�(餋ז��;�+\��0��ֳk�� ����o��\০f��a��Q��_��.u��Ӄźr\ꛝ�n��ؾO2�V��y�Dߛ�z�B�:<Y���im��96>�����֯���A����ʥ����Ao����׽�oq��o]��V�z�L�O�7t���Zo�δ䥫{7mVp���M���/ŷ��:��*���Y��H#���w���(Y�[���[�L���e^w��c�>o�od����S� zAͻ�A�s[`Qh�Vk',˾d��6h�ܫmp`�K��t��(�{�^����IEy\ �ݚ���e�氾�ڹ�z粏v�gv<�^����0뮐��{[)7+�+���J;S�U�Q0��~�A�.�X*�)����<�Q\�.�z�Y�d�"MyZ�e�*�w=��Y�d��]w7���2>��@nk��D�3��۝�L)lhp�&�m�s� K-�|��
;\�� [Na�n���%�w=�j�$����W2�z�=� ��������Zt����[u�z��s�n͗���s��Yn�hϔ�:a �a"�n�x-9���!$m�$Թ�z4ؒ���yR��۴3�9*ySm
T.`;9�
i�m��J�r^�ۉǜv������T���2,3z�anitF%R���{\��{�^r9;u2�f�;��Խ�B�9� ��rl���s}NhlR{�1�j�X��nn۔��U7��Q��7�-���z�.�wչ��rUr���`�uݱէ8%�22�c@�E�ҽ�*�>��;Z��d�Ҕ�s3{��.��U}�oVK0�\�8he^�42�y�]�q�#�s�z�+M-�^����қ�_����&���+�{fL��T��Ö&�b��8���!�j��yL��޲�V���4+��������6�Ã2.2m�ප	���R�s��+"��$��'��gk{�e�`envݱ3T}�فu�������2� ����Fsp��ޝB�xWISJ!`noo\�_8(�}Zެy}fU��ˢ파ՓD�8�a�\��$=�i}�<�iMwN�W@�Him��ΓfuÚ���-Q��]�#t�1��p�:�9�s3R��l&&ܟ+�!�#_����3Q�|��S�n>�7�����ò�X��������[],h��7d�BŜt+~�2-����y����{C��m�a�71�ι���=�V��������50Up��&�	k�ӱ�':-�z���g��Q/yh�|ҙvw�M>��B������A��Y�ԇ.ݚuqFtqlL��.a�p�/���y�owS�����yi�_+�Ҭbw-��t���N�Y�����
�l�w��� Mt�x�`Y�c�v�^L]ϲ��Oc�z���6���X��l�+�շ�p�`�ͥ۾�\�=f�#�$hc���5�y�N�֒�;�v��ˈrW��=��0�֌��F�t�V�+���qW��N��^��90ﳍ�y\������\��r��8_[C*�os�jK�������o��$�9�N�NI,k	$��$�I$�I��I$ޝ$�I$�I$�I%�&h��v����sr3hZN$d�a"b	�2�(�
�N�0e�	A�R�X�A��D�B�h��	���1݌(6d�+]F�槨���m�w���)��5��/PSt2&7-�A5/Tk��r�ޥ`�)��(�nLƐ�0��M�M�yvnw^$o5���00�`����C��KL0�&̑�fPd2������=l��W��ej�n7�z�-����j8I ��;������	S=��Ǚ-$�@�)�$%��7#XN��"�N�4c�2�jI�� ��6l�w00(BM0�b2�mÆS0�R5"L�%��B�"IZ��[f�[	;!���2�V��.�.&�%H�4D���4D�8jȲ	���%>�b8Q)��,�%�#A�h8Q���R���͛Ӱ�m��8I�ڈNڌҖ���mq��rք!�!)���Ii�"aGB&6;vl��WH�Q
2����j�FR@��2�B	�h*IDj�!0\�ŗe �f�i�T��D5h8I�m�Y�����I+X�0@Km��@�-k4(i�fH	,�]��S�"I�,F\m�{�ܾ�\f���!T�P�M�؁Vq9y��Z�:�Lo&�a		q���O+m�:����\a �1!@�if�\�� "[i,��$�ca�8��f�H��e��%�&���9�r�/���j�fH�3
(2Pq�C��8o�؍��d%xW7�a,��bSe^��w2�ih!�@��
 3q(ۻD���HM�M@5�ټ��Hw)��5�$�30�p0l4〔:�]�SPl�f �
5��������X�A�0`�0�%y�J�Y��A	M�:��"b��h,1�e"Җ���8����jFP2RM2�β��	�?���$I"'�V_�����O"�G�R~��~y�՝~�����_�{�����8�Bi|���o<�<���"�ZG]�WΔ0�(iTu%r@�U;"�ݝ�ݳks
�Ճ�����s���K7���6�g+ }���qz��l��fu�J���_F@"�w�V�Or��x��g*��n�QQн�G�U��]��k��,��>wr��U��KT�>��>IY��p,3e�D>"����}���\���eN��oqS����Qg�E[�c&`��\-�L�t�a9����oQ��i�u:�:,YP�e���#����9eVߪ�K�BEc�ι��SVى�[�9�W��K�U��s����=������QR�*}@W`��ȴ@{�cʃ�l�X����楠��T�&�V�����a��T%!x��ك��R��6��/8�v�CR�>�����h��緶w�i[.d�\��v	�y���rͫfqR\��yY�.�]��!�#a��b�f�'n�8�q��`�[���yǯy�\"�դ
���g,3� ��4s�S�b���Y�o>lكGe!��͛�!<�n���2��;�ݑ�Ad�KK�q�֮�#U�r��|����������o�Q�kZֵ�lkZֵ�k[ֵ�kZ�Ƶ�kZ־5Zֵ�k^��MkZֵ�|j��kZֵ��kZֵ�|j��kZֵ�ֵ�kZ�ƫZֵ�ڭk\kZֵ�Zֱ�k\kZֵ�k���kZ�֫Z�8�kcZֵ�kZ�ֵ�kZֵ�ֵ�kZ�ֵ�Zֵ�{kU�kZֵ�V��kZ�ƵZֵ�k}=��w�WV���g-RC�S��2[x��Bвn�0�s����qPW՗�m��&&����s�{ScT�<2�JW�qf�̱X�
�����6��N�"�V�˒��maͼ��!�sY-���т-q�к���N��C�*��SkjmL�fjI��4�q�YBGUU��u��Ӓr�W_R�%>��ɋN�ۦ`�8���  굆˚Ġ9�)e�"�UsUJ�8H��\�=>HFm5/5�� ����`�w� ΛV���;Q�L^A�;�s�����S�i٭΅6�4u�ʻ�C���1�fʂ�MJ��V&�"�.��L�Uv�x1`=Ʈ�K�nv�T�`D��T�S��i���*�Z�g�ena
v1F�nRTe1�$��O�S̍�Wv4�>�4N��\'	�﯁'$qw]�%SD�=M�̶;g+��1#�X�(H�\�b����V�֤7yإY������i��ʾ<�ú��s�\��&;K��k���h�݃� s�UM�o(�]\��$\U�ø��Ͷ�P�^�3u�J�,�2_\��󎆚��9-P�[.J;C_u�!/M�� (���Juu�uu�����v��Zֵ�Mk]5�kZ׶���ֵ�j���ֵ�|k_ֵ�kZ�Ƶ�kZֵ�V��kZ�ƵZֵ�k_ֵ�kZ�Ƶ�kZֵ��kZֵ��V��kZ׶��Zֵ�zkc\kZֱ�kZ�k\k�ֵZֵ�k_ֺkZֵ�mkZ�5�k]��kXֵ�vֵ�5�kZ�ֵ�cZֵ�Zֵ�kZ�mkd�n����9��wݍ#̪�-����`�͙�OWd�q�p��=�k��MfY���*�̛k��?��(�}nL��KWCf�|�uX��6��jC���oS��Ԧ���#���7a3ݸ��*ZcA�κ�8�1Μ��f#*�G�)d����K�,{tU
"��3�w^��1uU�-�>�J�j��f�ub�j��TL���+���Kw��_z���漭�6��N���J�1�X7B�+�^�)qՄD�&ʃ4j)U���+Y�iU*���LbRY�H����)$�c)�=��v��������ɸ'ī8r76�s�\�گC��:��q����sa���}.�V�s0ᡄ�K$B6q�t��B�N�Ӯ��7��2��]ئ{t�'j��n�,�,�wa�l�ۉݪ}�����&L��R�Hk��.�n��oMyB0-5��
Zj_5��wz��wD'b�X��t7�Pf�٫u�d]*2l�
��sx�W��L���zr�ޔ�jJ�L�Puढ़����hL�u*^\��پW�G6�{����NT����mo�f�Ac6M����fc]����s�}�vc�1�k\kZֵ�Zֱ�kZƵ�k���kֵ��ֵ�kZֻkZ�kZֽ��{q�q�k^�ֵƵ�k^�ֵƵ�k^�ֵƵ�k^�ֵƵ�k^�ֺkZֵ�m�kZֵ�kcZֵ�k_�kZֵ�k�kZ�1�۷mcZֵ�kZ�mkZֻkZ�5�kZֽ���ֵ�k^��MkZֵ�k�kZֵ�mk���o�����{�~�w��ۍ����4����l����;�)�|d4/��k����f�xαl�c��K��3����u�)�m�]׼%�ef����-�0�xz��E��7�Z���X�8ݫ��7��e�����Xj���>�k��t�m�\Fa<�ʟSO����n�b��%��r�ԗJ:Ae9W�la]��9us��HJU�\Ί�:X�@��s�u�F�#�sMˬ?d6x�
[%'[��R8�=��TW��.�2�)�@�7n=ʗ/mVx`�L�q�����cZ�̲�AIfq���
��jDp�Nwc�W��B��s�Wcm��W��Ū@���cz��B�^;|N�O+���yQ��ɢ��oK�[;Ϩ_��MӚo# 	��)�+�ZzY{����5'���&��/{�u{y��$���k���`��ʎ����$CU�R�=ޱ����5񣮘��މ���x��;�m,�,�%�n7��S�Qb�m��>����LP�Xi�����]s4t��le��Fk��r��QĹi����ɭ������q����٩s��ˠ3���uD]-�S�u��VN�<A��c��L��ӧV4mvUR��z��G���@�f�)tdǾ�i����Y�������+Zֵ�k�Z�kZֵ�tֵ�kZ�ֺkZֵ�Mk\kZֵ�Zֱ�kZ�mkZƵ�kZ�ֵƵ�k]��k��kZצ��5�kZצ��5�kXֵ�vֵ�Zֵ�{kU�kZֵ�kZֵ�lkZֱ�c㶺kZֵ�{k]5�kZֵ�ֵ�kZֶ5�kZֵ��kZֵ�kcZֵ�kZ�ֵ�kZ�ƫZ�w�]e�3p��^;܎7�2���ܚ���B���0Ї�ACxW��M�*�������,f�-�0�WV�e
�*Vc=K�֟����aq��M�'�V�<��J�&���̧��q�:��E���=q)�n����m�p�V>i�Q����,���ZT��+�fd�N�T;��,P��>U6R�)�J�.�ru�>M�^ G��\c�q��{�T�Ễt���|3 ޛY�cl��������m	J�����8��0 ���;}͇��&�^N�F�h]���z��c[Y�{��I߽^��
���n'sU4��3ښ�o>�>-b#�Ȭb5��a���>�6�4yh"WQF���N����E�;9Բ	�{܀��՜�ie�Ud[atl�t9�I�TJ����w�^�eu�$�Y�YH:C+ӵ^k<j+��*q����ͺ�:kʵ����ܞ�2��ڕ6������
WC6�~�����:�!��i][�;��u*��^>�=�i����Ҩ0� ��_&V���ôñ�K�H��<����|�&��#�+$d��@�Nb$>���|6Է_GW�Z9��v"	v�DZ�*�k�¯������5UT+htŗe.'ٹ�1�Y9ӂ��Qf�/m6�6X'n��]cWw�*���
�k_B����n��zi�(v�7B׶����bO*�2�&�x�k�꛷�c<`(���v�udX�8�ї�k�s�؝��&���U��fY����Q ����Uy53E����K>P-5��]i5ӌ� �ٶ/�A(�uIǱ��mq�w�̧ONL�k)t���΋ �Jy6���"E���sg-�-m^�}ԡ�n�A9׫ܓ���ɵUU(�Ya����5�5���)W�p�-�.d��x[� 6��1��v�!��j��l�
��Ɍ�0�݋�����]��zl�{"*��0�����IX���=�%�;��*���2>��\+L�~����T���1��DoO{�]U4o~)��(;ܦ���KssC����bʯs��boSe�{ޥ�܎W@���tX��G_e]���q�t�Q�K��jC��IX�W�ݬ���ԓg%ֆ�n�l�DSGq�v� ��[Pm�s*�u^'��՗OgZ��pn�!m�2��`M�6,�u{^�e�J=��
h�_D.>][}���eA���W�6m�>g�7�F���V�и�]|�z�ۇ.g#˥&ME��C�8�a$���k�Y�ا��wרJ��.{�a�k';^�)���n�6�����wS�5쳑QOx��,���q�HZ)[��J�)J8[?U����5�� O����v���v@Q��,�.���׽=�R�y� k��%�LC�Z�]����8+�ފ<?0N���7Y��G,�������Ax˔Ֆ�#DCu��!��&w�R⣝��/�ft��Lmi]��U�JN��f���uZT����uFⶌ�]c�[<w�f�M[��T��Yxf��홣u-���Vܩ�鎣�c;X��"mQ��ͼ`b�ҹy�"�7���t�̎EW*"�q�LeT]��{܇;͜��ޙ��8{��T�N�J��b2��crⲶ��$q!9R#h��Q]�V-K*�Â��X2�L��V�fM~��me�"�m�wy^��|�-�/N�rL����+-Nޒ��[`^��cyI]r�j�v�qL
�ueN����,�AI�J��=�E��/�t[��ˊ��o� fիw�r�R�Z�Au���1�^� I���i}8�f��{/7-I����;��,���y�j�2�TC����a�2�ڰ�{$m��q
���س]���̄�:S��!�)9ٻP���	���۳I�!��+r���*�_i}��{ �x��y��pl��G-$�b�� ˥:tk1�`�^������i�w�"V˱ٱ�X�1H�Ʃ�F��GL��7z�P���ʾz:.$d���LU��˱C.�]p|iR����-�K����훛��r�/��煝33���1v�������n��M��P�UC����}�L�����nJ��j u�K1����՛�L�޼۱�����W5�*�@�ݕ������m+ӖT����%�KЎ�wo�f�ۮ>�e�:����,��n���.�FG#��"p�Q��Wm��͆�����Ruϓ�y
�uq��x�oy����h��D,3���n��e;�e�ء��1w5�z��2�0��5��n�АT�R�(�Ӂm�W�V;�Ti��v��1��P�Χ�:@��vsj��oq��6_M�/!�n�܀��Rk�-���Yӄ&�n;�k/5���nl�S+N���ܾ)-�JxvJ�i"H��a|1��
��Ѽ��"����o*��g��r�.�E]�U�3r���Pf����O��"-��z��5LM����%���;U����ƨ3���]R���@@�2n�l�W��AwbWP�Wv�*��[���1X*l޺��lm���>rY놝LB�;z��@�FJ�۝2`�*��F���L÷�ג��������ȮT��
M�&r��n���i��|{V
-MĮ�Z����B@��wwc���X�ɫ��v�ZPVs/�9ohr��	���	�DR�UC_^1/�ZjB/��t��b����b�Ā����v�[t�U^��9��^�����ٶ�Ӕ9� �z�zD4B6W���P�컧�i�6�c� ����쪶j�����T$��c4�,�s��L��i==sN[X�o`���ր�=1�ڗ�1�JG4vI��аm"hY�+��Ю�+I9��պ��;�L�b��.��T-�����#�v�1uS
��R���a0P��I�'.*�[�s.u9��.�Y�	0n��R5.����N9\-��	�	}�_^:�25�v�8��2%F�\�[nY���[���S^wQ��ӝ��,j'P�'U�n�$�n�j�SS��&]��޳fP�k���a��*`,�.��ו4K�F�ܻ6��sA�ϋ/��٩��0�4�4;h.���Gll�q�T}�0'�J͋�����"י*�72�:"�ѣ�r05��zЊ�֬N뤌[ȯU�b�:5�Ջ)�
C��Jo`�)����eu���zrӰ˦�eYPQTjn�]�VNe
���1��ʀ-Ys��Zf��[f�w]YIi����ṽL����=P�gxX(��p�14z�����Z�ԙ���#�6����b�k��O����-6/�L}��/���M��k�^�;o� N]"g'T�M�T������뫖r�ƄMм��6��N_6M+4��U��ō�%6�I9��V��D����-�̒�ۭ��� O��y��E�|.��\f2�_��ӭ�L�I��L�Y���H'�m�QN��GZ�X���;We\PgWP����D���%��V�\F�`θ��&��;���`�竞�U�s	wXT�I���I�k(2�����F�ف�յ&���n���pC��I�ڜw__SB����y�ُCŴyg[A�j��IUv�N"sׄd�(S��v*�6>`�R۫���uCOtfB:���wP����:�V�lQj�Sx�l�9^�6�.s
�i�^e�$ �`ۙ����Р�?d����������������տ�뗟�?^�ru���� �!Eb�Qj6�A,P�n�!��Ii��i�J��I�P�S�8�""a+�$.$�H��NKD��-/��S��J��4ε_�?$�?glwBe_s!�F�1��c�Z��,\�qG��P4�SJ����txQ���ܲPC2�YF����Vs=v���=垈�1�	SzȞ�g��FN,�2�f�R�v}u|U��P��CU5��]	�r�7����P�)����С�R�÷�����I����iF��ڊ�z!ךR��y���"�ڲ%1��XG�p�5�8�i�9��.��������AI�6
��b�wy5B:g+SB�V��[���Ψw,�#�^�k#V�0�k�<,�qǼh���:U��	JI2}��^�v��}pGd���q{P��[xq-{O��x�uob�ݮ1(m0۳��'f�Qˑ��ʷG���Z�MM�0�*Kݰ�Gv�]�)�I]�d-��n�X]{�+�l|{��ļ��Y�Q�.}�Ώ)@���vJ6i�O�e��N=jT�wh�b��,fX��΢bH%�o�ep@լ�᫝�V���m�{����s�-q��2���!����a��*�Pu�\�9��.�S�����zqk�A>����%�@�on��p��h��� څ�Y�ȱD�l[Z�H��&���w)�L((2�A�I:�'�lK1#R�G�KTn>u�9p��K��TD�05�DT�h����I6�H�-��HQ��)��5��xT��FYa�lYJ$�D$SA�)�&�2�Kp(� ؔ`�B�(�V�%�5���?q��Z�zs:�'Vu-��N������ֶ5�kZ�۷nݵ��l�j�-��1IT�JI��h�3�r�ԫd�m��q]1�kZֶ5�kZ�۷nݵ�|�-[���<�kQ1AUL{ٺ�4�b���lDTRD�{)�8Ǧ��kcZֵ�ݻv��Z���_����Ry�k���UD�Q{Cd�=����o��o)�`�Ԕk&ƭ�7qzs�x����ƶ5�kZ�۷nݵ�x�騌�����v��}��DE�4��#�6��l5^�Tl��䫎�?vE�<1vlm�j�b 5�u�cY7d�T��B��RQF�۪��@֋`��T���c�Ѣ���uJ�*����F�8!v�T)EEZ �hS[X��d�[d/\c�o^n[Eh�Y
(-.k-��ѣ���6KX�lj�j���qgF��F� �6ն�H��m����QMO�^���:(	�
�d��+��**/rt���Ilj�h���5��
J*"���c��5{�Ji((�|�AML��QBS�0 H�o�6�r웅Z�Jd���V�y�3;y����H�ݳ�45��=�1���ݪ�wmd0N"Ӛ��vӽ{�to�LPpxURJ��8�4XrH�p&
	���Yn�F��h�t�͔�N��v���Jt�׭�� <6�y�a�ܴ�/UDةE}��Tt޹~�탻�+��_0-|���[S�v�H��������nw�����)�P8ը�&؉�{�*���x߈�Ǻ�̂RĔ%Iz2���Hvt��ʽ2���GuT�4��]�ϧ޽bޡ�h���+c��
K������=A�؍p1������X��{���S�v՘��Z��\ڵ;��eO��`Y��Ǆ�PX*��Dp�]�_s��f�:\li����	��$��QOV����CR"Cw%I���{z�/%�u�Bo������^��n�^�2�YsCF�>C�j�;���u�UI"UR�P3G�}����}:j ��=��IRD�ҧ���n�� ��vq�Qn�5�#@��0�Q�5�pV�xc�Ź��;�J��nW�۪��KY����}%!�7~���֛f�j���D+rl�l^���9X�A\��>r����uS�钔<RY�_���Ё�|0E�fΫ�ny�S����۪
묱�䮭�L��2K%Vп/
�
��e��|�c~�fJפ�z�(h���z����&� ���"f�u^�G4��6qZr�u�B��5����9Һu��׼��
���*b �pu��w���+Ѯ&�+ْН��Y������S�ͭ�VҤm��I�@\ƾZ�Ѩ�г#+&|�f�B��[���Ƥ�S'��@4�[�7�����}���4ʒw�7��7�J|��7�T��k[-0(;�ž����d
dDF^����h�e�������,�>s���h�t�b����k�R�\+>g�
�H��[6��m�r�F�ɓT�FV^Q*��'ڃ�^�b%M�f��e�KX��Nh	�6}���ù|������Qj�N\/6�{w�Δ�S�m˫�L(J��^��j���#d����օIZ�C/ВH�HZ�{��V-���+Z��jح�����T(:̪sm7u�U��v�� �AgeuɁ�VpW{JM�2�ͭ�ACWA�L�C�V�G^�.hɷ��[t�}k�օ�+ֳv]���흈����]𵓷��ot��u��U4h D윲wt��h~:���Z�2��`,/�rS��5EН�{��;1L_8$l;�}|�K=3K(	�>�'�KqP�3Yd��2s�gu�eV��Q�DÇd��D��N\����!f��я1���$�n��#u�U@N�U���3c���!���� E���cgb�aM�ڻ����2��>�|�>�<5�w�}��ٓ�l�v�)�WL+�=Ϯ=�#+Zh�D�5��4���l���Y>'N�AV�aK�;���{�������{@��E�qRswC��Hn�>s
+���q"BJ�i��!���a��֊'.c^FY3�<����W��LTx��������Q=6�xD����wS�罭	����1��T����_tuu�fHz���c�a��R3ݹ�c��+m����Q]MgMݩNco�V��R�u��,��[��+���A9S��7{˕���=��z����Ԫ���.�+e��<�+0�3{�9k��훢H�;��mK�o��1WIyr�a���<te���U��y��`<�o�tN�5�o�E�ۅ$�i;q�s#z�A�zM��`��v�4���3V�����<��4<g&N�#�LcȫgCs�jDX�M�`�;ۍ��I]��X4/�Y���4�d��4�EJ���*�cӀ�[`W%����5�-[ykL3��"+ׂjk� ����5h�Ig���-��V������pt�@�u���]9�}�P��ja�V6eat�m������ʸnr�|S��f��B�h�G���iVf�&e�����sS�uWzE�=��s�#tAO������aOI�m��
S�R|7�&���(�J+w��SJ�� �l6z�o!�7�v%\�˫�B���+�y�lS��F'�S�I ���ٌlϴ�dy�!�<�nf���� ���JT�`��4Ld��tڿ(���}��������y�'Oct�G��ٺ^�Ǽ%�yL��2�iα�>��4.yWk�.�_=Cu�.l%��@ۄtKPȳ*�l���-N��J�ZKd�4]6JIj�R'��1�4�Y9s��o�v�Թ�#ӕ|��3%���,r��{��<�퇞�o�]��n��]Ltg7�2x�^Y�Ӥ�e���4�$6���,>NW&g�*����vw�s���|�z��n�㢙H�(��!h��������{�੯5ei���t�����gV�'�(D�6X�B�h��V�
X�ih�0Ɯ0Yi˛+iF1A˽��M|k��ui�v<5P�8�z���׬�����WkA`P�[�^���:2�����ǥ�C��D$}��22定e�QZNa9;�Qu_1�(I�h Ϧ���ws*��{&[��f��YV��J�㗯<�BV��w�4�н��-��&�r�ʂ����w]*}�4�2P1M~�o�F��ۊ����O�j���ʌ񗘒�٩�@<{*��Ķ@����Nh��y{��Y��.T��?|8�� �w,��(��G�&�����IHm^���F�@�^���>Ν���s���MV�וG٘��5(:Kl����bh�(9CM}ZO���)��?�,X�����SR-7���|v�WF�D�˒Sm��T����K�̻�O2e��y�9��vGlaζ�ż��ܡ��a<��>/�A��7*l�����N���e���8�B������h������]�x�޼��=<<<<*��URN-]ܙ��r�R���d�[EG�4��P�!�%��qQŪF��0��c�fgu^�&��Q)nʽ0�.׍�jsf�8m��K 0N��w��;�{�[�b%L�wc�޲�vø'7&���ڔo�׵�d\!�aauBvL��kD�'Y�֭�m�Ң�Ӈg`m��a|5��%�Ŷ`��\l�زٶ�޸�������]
���&VD}�����7�Ƌ�!	��`������/�wՊrM2	[~���~���>ؘ���M�?�}�v��¦Ԇ���KVX�AϭeE\�ؘOf�N��bPO��i�YN����er����Oؼ�yNa����9��Ig��n�$�3=�:c)� V�N��W�əb��w��\נM�T�T���ѱ��:f��K���{3ۛ�ߏ���s��2���-�5a�|�p�~�k6X<�d]��5���Z0�C�e1N�>�-���%����� �\��Oa�2��>��v��TU�t+z�J�����y�[��VN�=�&�t8�F�"�����s��	� N�۹�M:������h^&pڨ�%�5����$�h�D]�倆�J8<��o�e���4�^baB���W��V��2+N�J����я��q)IU>����X*d#�N�FL6�s���`
�����QT�,�/W��M�f��|Q��;��u��AI��Cy>���[魭G4�Z}X_IQޡ����}�����^�ќ-�F�]�������<�o���N%m���a�FmH����eg�����@v_��EA��S��{�zˈ�&k\�ue�r�9�&nC� ^�l�o���� ���De�Q�7f֒���#�XW�t�N� �G�*2FF u�3��5���1�M�	�yB(���^����vI���:  ��=|e�]�����[��m�'u������E��N��nnj�"@W��Vy��W����EvVe�̒�S�3-|m�-qY�|��7w�t�|6�ro���4v��r��_R�O��٥��sQ����{u~�
��������� C$%���*D[�$�dl��6��*QrӱN���j��tW��:�����s��U�o�5/c�r,�����i�3����]  �HS}��̺�rfӻQCC
(��	�R%�]�4�Ҕ�d*�6�v�q��k;d��4�fv�rna��t��(�5��Vj���q\"v���ļV�Ae`��m�&v^�"R�3�R(q(L��4w=F�j�N�W��r|�jS��!�k��^��`��k�B/���`���.�<w�P>%-z��K+H&[B�Fn�*_b=��G�a&�}x*qӥ�<٨�l�N�E�ș$�R&����A��Z��]��a��-��52����-�Y��Fb,�[ak1�j�c����d�<�B=t�b	��YU���:����3��O�/�Kۤ�y��O͵�1���׆�
��Gt��%�:��x�a����6�WX䫈�.�T�5��ֹ��׌��v��Eʺ5�{���{�:�^�l����{�}�܋�3λ����iZ�]Sy���N�2�t����)���A�`*̀Ƒf�hѣDF�Rv�gI�U��TeQ��*�`��g�͛qi$��O	�-��`1�t�mn��-U;�M�Vj�U���/6kV�n7T�M���! U�Q�_g�{)]�/���g�'f��>� :2#n �*_�$���ɴ5�[�'C�ENB�F���K�I���gݠ�󌻢ih�k�I�a� N�Fb��C�o�qj'\��>��Mpν��Q��fF�0�Ӳb����igQba{Lx�6�,^�q���M0�D�9��Nd9��=��u�n�f�NZ����`#�}�b�g�0n�%���H�J�*-�)	e1���%{���O}1�(;��A��gӴP�9�E��4k����x�CD������'"i�})��{5U��r��f���� ۿ'�e��v�>U;����=�������r�K����^H�~�'}^�k�M�%�LD�i�{��cj�&�Ut�k��7��w�f��WF+���Rf���pm�<%%X=^b�������^@�����A�9r�\�P��u@�ݔ�e�s�&g�{,J����+d����J�Nm����m:��K��:�j�4@4h
�9�}��𩧉�S�e�&MV���$�q1ӈ)�F"���'׈��Q�yw�t��+6�PC�������y����ޕM�v&o/Q������K[k@���B��5�y]�u�ux�KݿlW�^���:Fߥ,� � Kv�AZ�:���:����/�(� Q�$�҉+S��8�2�t�͍��)CZa/x��v5b��ձ ��Ko+�k=Y�����-�]��<ψ p�OO��P"}�lW�U�{f!��S䒩z[v*ާ�p�bV�����<v������j�&��S�[Z�j�J�lj&�jY�����v@�>�;{{6<�4C+��ێ*	�ɬ}�آq�ZA�-��<!�0�6��� �h����w�]�
���u>��u����6��o�%J:�e���nd�w�T��כU�7\c!�ݺy߮L-]Q,��+i��;P�Ȭ���Wt��f��F�2�\% �`���N9��ƅ��1V�r���]�}�q�ͮ+3"L>&�eln��&\��bF��������A��뎜�2�=��ڴ�n�z����Vɾ�yٖʭޓ]��ƞ�B�Yx��<9���U���7�ǭ�L7��6���"떩:�f�w,X����T]�t�to���u��I��md�^�g�����g�J�"�Ɨ,�c����X^�}�����:x�ON��C$+,opPqT�J}�^ӹsxVЈ����v��{)��S�/��\n���MgS��E��\;�����i��@vy�'n�\�qOj��v°ww+Ƕ
��J�x�*��v�����2�^�'�%Z��5���lJvhM-[��	�^�׻�kڄs�>��GkRJ�qX�M�ܛed��-�m�3������xv;��cUL�E��l�j��V��ۮ`��n��o]�*�nұ���5u���Vz�&�Y�gP����s��oZ�uh�����E�^�Ïy�w�3���,p�*�l�n�Qܡ��ȧ\l��#/����^TS{fv�mTȟ�Dr*�����n����^��sBS>��ȥ=�R.n-A�uW����A��춟2��6�L�W���\�i�Ht�U�Y�/�K�o�6Ϗ8���
yۮe4��;5ۻы���*��_2�xC�v��kK8�zb�DI+��A#'UbfeV���j>T+8��pvU���\�;OI�mf���t�z�7���{I����=:;�o2�}�1᮫�T�5�X�gV�Q\����|�wL��s(í��|����`J��y��n`��T�I��R����Ѯ5d�d�h��_[��oC���f�Z���	Tkd��꼣�k#��R�_{�-�ڊ�R�J�o\�uU�J�B�we�V�*�w#��ʔ�&�쩽z��ᔣ����n�q���8����0�m��շ]���G�N��9Z��i��Ցgd*X�W��GL��i�d2r��<ss3]�Z��v1�1���8��;��.xY�񪲽\%Ze	�`�B�j�x��U�̭G����7���)���ɫf�.R��0��v�����}����i̾�޹�N.�:��˻���"�3�-�\�,��5��4.��
�<
	I@QA�:����֊h��j��(�L������~�ֵ�cƵ�q��ԲȨ`�h����0���J`��j��<�G�9�����~�5��x�v�1�kZ�Ֆ�m��m~d�GT�QQISUF�i
*"&�s������|x�+Ǐ;cƵ�jl���%����:?n�
(�h���h;y�{�*Jd�Mzk^�׍x�^<x���>�_���'|���|�!@S����$A�T�ɪ���H�

����&��H�(�9B$M4E�1$KU4O�t�,EP~�GE��*+�8�r[���F�(U�4j��5U�F��E�;j���Z
)�ii�M17gT����(�(*�����#���{�XҤ�������1;�2Q���L�RJ8,:��/w��y����<�y��0�)}���-�+�F��DҥL�t��u C0>ei������/�~zw���z���t@Y��FnP�O��/��y�r����&����e{������hl�^�ݞ��B�GՏ
,��^��a���hy���G$a:jB�o��O2}��-�<��{�����}jƆ��}a�`�C|��h*ua��a�3כ �dS�p)�pzY¹�+:�+sw��{�u��,�@5�O��H4!����5'^�ʬb�|��b�U5�k,��=��J&NÖ�d^�m`�ާ��}�H��1ю�a+���A2/���o���<��d��;:��t��J���k`8s��=��鯎׽�����Ś�.b�dYԋ�����p|����N�	y/��5Y�P�j`m�o2Ql[�_<�_�.�LPC�����xaȸ~Q��X�k(��G7s�����kw��[�0�  �O�:jx�Q|�Rp�T�,U�4/�e7�b�byL�4�jmuK�ލ��}>����r���������$�y����sج�I����g��z��:�χ5��z=�,�9�xxT�7��M�ߐ]�^ô�n�y���E�Y-�Z�k� 4���Uo}�}����-��e�+͈	�,�+���k}��
�î[��T��h�C+{�U̴��z,f>���uV,Ø�ci.��Z���Ҿ��0w<ݗLK�o��W7���r����[&�l"������5�8��ǜ�������-UU{��������8��/����ώ����X= 2 ��K� :{��'�?Q���S9�Fj�:��{��xi/e�`J}l�����!5WPC�[�b�,���n�B!��4��D�#Z���-H�N&��6Bg}^�B��?k$k�X8Α��
*���}��z�؏�����5��jt��Ѩ���9�<<,�Q����ٟJ���!><p����<3;y�q��X�s*|�:k�'i�۲%���g7��o�� a^�vQx5��)�j��x���@�yJ�s��z���)C31��t��E<�jUh!��謃���"	���*���c�����ί z����䀓�'��To ��v���_��UOP�J�P���է:��@?o >��>b�J���0\#">��VJ��a6��މN��+���;�����Z�Ӂ��.��C�U!�^HlQ�,�.�����Q xk#���Y�<�A��{�7���[@NZ�}Y�r<%��J�����$\��`38���w>\Ʊ
s#s6��{������Ӆ�k�@C�a�濏o=ۡ~�=w�|��ަ�őp�m,�:�Z�NeQ�1
k��9F���Sԍ=��S=S��]��Te�7�Pl4,��w0_���B~NWd�e�h
�vƏS41�0%F@�j�g���6���$
'G�]aǓ�h>k��>�T�W�k���؜��v��>�;��N�/��g�e�=���B��у�*�^A$i�Q�,�Q�cn��ː������s�<O<� ���
E	y�{����o��@ r �$04?x?�76��#}���tZo�[��bS��\�ë�{�q�3yخ��T����Y;�Kx <��8a��=k�dӨx~�c@]�S���|=��o~�b1Ʊo�9�cn�\:��uܹ�����l�G�vP�G���R6+���J
5����� !�X;sy
�-QN��n�|Q�v�E��� 0�=j ��r���1��{�(����1@�����IW������t�UP��}�z1`8��B�����
ض��5 r��w@��FG�J���,	�!���[2�ѽw9����%��S�K���,r���OY���@-��:�560�;��Æ9*��S5J������=����p�����H�2����	�y����I�]7��s�%��kh��~S}yI*���*`����3�!���x�Ɖ�J��=� ���hr�f��Q�;�0ݛO�a�øf�y�رgzp�E*�P8B>��� |VR�}�����x�)i�<���׌̦�wқ�^�DQ��/{wn����1>��ކ`7^��|����Y��k�\@,T�_W>`]5~ZE�W0��g��3tt������ܣ�/�j`ڻ�o�����6V�4>z�:<��e���k~�:-I�87�y�6k�fvd�N����bݚ:�q�/*��8��%�"}���=���tbRw�6u���ý2��v9�^s�'�_g�q��8��8䜲-Ib*$�%������;�����5������� ���R�f��)��}�8^k�Jt"�>|F�s[�n=���v����X�/M��͘�-��p!�[�#U���#B��^��pQ��y��q�|��^����mr��{�C&�+�B<�~Y�b {���y̹�k�[�u��͏_��B�ŉԴ�0s��
�5�^�}X�s��:>ƕ		R�������O��DW����9݇�Jp+t��&��0���Y���x{��G��@a���XQc��$�N����!�C�*y��#���o����o���j-NoD�=� �}�(�v�0o'��
4�^.,+�	kp!�����˖#ty��ņ��d�b�������z��N��^��i�W�~p����X}~����/�����A1�`x�8��K!�3J6��Vw��Pn7"�9���M�no
F�X�)��]��d;�a�Ftv��y���ý0�o#f{V�b��c��J4Ԫhi�>�}�<��ug�k�-(9�ˡ2�q��y=�|�[NCj[�۹x��*� ��:�4{03 ���Q"7���x��L)����
8�˕��MwG����8��ۻ.��j����l�\&���˹yץ��:ܺ�6yGL{HR�-Y(�,[~4`��3��XV�L�] �"�� 
�vE
��#2�����g��k��3&o�h��\�����Ջ3��{$��Z�@��\�g�ђ!�U��ӷ8�#�8�',���*%���Id������ל��__>z�C�]H@��m~l'��C�:��\=ʎ�n��m&M�s��Z;�[]��h��< �r�)���w?��m��>.7�� ��O/�Q"w��@C�{��������<K���SE��o.��ׯ$ނݼ�]xh��Xp��9������0�Z�zo���/]ŷ�3�*�=��|c����_0x�� ��J��h��Mv��烖*����s	1xEc�L��o��86ϨS �ij���|��i������+�f���}���T@�~d�Ղ�MT͵��m��E��9�ʻ��v>ǎ��C��쥠D��V"�W������'jz��P�8\S��m�[Ǭ�����z�L@3>@B���a��P���|C8#���k��ތmh�@:o�_��̿	���
��w{ѯL5�#�^H�v*����eb���1+в�E��~̯և��g���p��Il��Q�0�=h>��n��!���s���R0�c5X��O償%F�p{�=M��w©�K��6�ʖn����TV�q��.�G��^P(�d��/H��]B�Ϙ��c�zMr���$QL�oG�o�T��IO����2�l8+�������8�����=kY��
�=�(~��L���Kv�!�7�S�ͱ��α	߬���}��r{�Ay�g8:-���;��a��[�b�}�0�ur5�F>����3{̾���B�~�SN�:u]��t�L��ҠD�H��xc��K����=����5˦\h�����3��0����j��@s/c���%l{<�/�K��Z`��DwKa�\���PF���C�S�g  lE�v[���S��˨� �dWU���bo
fzf����D;)�:���=}}����J*0�S�*���%mȎ�K�������ƪ���@g���W�ߩ������|�}�'���#v�-��d��|��#�_�vG����,�Ë��@�@#����+k��-��*��� �Wt�ݫ�`��{8a�Xˤ����4��(��ZG%�_�=����쿱��^^a�˛�U��oe�S�U�9�j�S�����y]�)�w�q�T�����z4��e����C�euVۤN����M���E��5�3Y�p�u:ސ>\�R�a�� ���M�g0���8`�8�>~��LSߥ�d��<3.����s4�'�0��TZBp&q�S��,�������;q��C<`�gd�S�sbcÛ��Cc�ҟ	v$�a��c�>��k�n��=��m 	�l�</LVW�a���i�P�ÍT=�����^5��s��1��ν�Ca��o��3-�&�t'n+,���d�RX�G�R�ő��vS
�e����XU.���N�d��Y@�¤GGye{)f��u�a�L�aG�P��gl�u�����^gH��ռQ=f���=i�_Al�$�H�(%DĚn\
 �L c���.G���@ ���`S �O<�t<���<��t-h
&��E
6�^�����z�v"c��)Jș��l���+�ђZn�φbf������f��,!��6���`����nA�x�yq����#��n8xɻ�\Ml�ٙ����}���++��i��_Ƅ����u��` {�r�Y����.��&}x�8u0��}���y�?0կ�>��+��n��t���.b���`2W5?De��Xk�p��/á�@v���
 ���������ZO�L޺�LhZ-��j�0���[c9�����Z��.�w���QR��Y�y���X���]G�  ���c  <~mנ��`j���[�5C*Ȑ�ݼN��ՏR��6m�$�[�7�C����� |��-V�C��ǽ�1파�M��Y�=I�fq����}b�^ua|h�K� �G9n���[��j`Hמ`:W3��֤W�z�l��<]��>7��yc�F��e���^���� x�a+>aǣ���h�!�">Ya�>�Ϲ�M�MZ�D5�)���܉��>����$���c�m�c��2�ǪH�C�����=ƫm|�qbLO'w�w��0<�[��Нd��3q���X+�[���|p�õܦ5�^>��.��Rڹ�&�9�=�Ͱ��~��d?�mm��#r�L�!ܒa+{D��i�5�&�/;�w����,Ct]�8��5��Y������c �#�:o���#��Gq�oR���Q�>��8ɶ_�����',�+�8�XI\q�(3�<(p�4"P������6��9��y�W�?��9��<{�J�|?]GCO�rV��{�;}ϕЛɭ��Q�7��5a�Z�(pG"��=��½�0k�a���}p��=O�Ix�@4<y[�A�\3��S��%�(�Қ��n��eL��5H{�<n�y�yX.�F��x����̡�$�}�@�~���%�ƪ*�[�Ľ��_D〓�v>�(> A�C�B�Y�����8��E�cP��Ҷ�j��r���.9�@K50�iNe���s�䁔0w�K�D����`/A�%����Ȍy=][���W�
����+�d6r׼�����}�R�-����x�uy�'�4õ���9��1�٨�#D���Pb���U�k�ѝ�,���5`�<�mT})+%��"�J����~D��>��v�T�o�p)��|xpd!�S��M׽��U�BsXLm���pzڦn�:^���I�k��]a�F�՚������<2��C���^���cy�s׀�Jݖ��=i�ͪ���.{����1A��hx�ߠ��]9����Zp!��ﾧɴ�7���U§ۧn���l3v��>bܨ:^�[
ov#���z!2D����{&����m pJ�i,���X�$R����j�:֞(��w;5Frɭ�m���yw{b����/�ښ���u���ȞX�_gӒ$���8�$��y���z�
�%�"Y$��-��|�>y����ϩ<e��y;��bX�����7wt��>� uU��zFSy��,M��'�{�7M��2on�A�xm:/�m��n������X� ���#��O7���Æ��n+��q]B�u�i����!�=ȅ�g�yi<@g�-o�`;�+���@(�t�]0	q��-��fև=ד}Z[���ނ����8Ƌ" ֑	��X7��3�x]�=F^��5���ށ�]+.���&/Z��f�����>�G��ޯ�\}򴻪��>v�QF�R
�i��v��� yd^�^��U�� �ی:��j�>��؀�-�"�?] �z62�,�� K�$OA�[@]#��~dR:~Ê����&�nG8}e�g��x���K#>u�m�,龺��}K9��%�6y�������m;��mۋ�kkM8.�e9�U����	o�5��z���&���v�o�nM�*�ڞ�s�M,��40�v��i᱀]p����Pw
�y�k���A�@�k�R�;;)0gî��w�|CZm��c�p*ΌM�����<Փ6
�0"�$�z` �U�ƒ�j��U�Hz��uJ��hj���*�f�b�G镳��w�F���K�����H�f� �����Q=�����n�ۇ�[Ʀ�tsH,u)g���9]oH'J��o�gs�;��z�v�������it��k���-��%y��J'�x9�� ��J�E�B�� e���=���S�͞o�d]�E���*�t�~- p�0��5c<��>�OL��!�ֱkK	1�=�ޔ���Z�a���[��� ��;����"��41R�w�]��]_�#�Z�d��|o���^咼zQ$1N�=��� !�_<s�Jq�+��cз���'�vl�������H�"���z����o�?���1�ё�<�F�����M7d� �(f?�p����i�jԌ��_63�u�5��;�|��	��& ����\
k.����%Յ�)�wK���Mp�jA+D'wLۧ3����zS�z#Ϝ1�!�8@���#�lE��%�qP��ӛɭ� �`O?�R��z5��srN��(az`���bzw� �}s�q|&<��w��g8t��ff�,�nOŶ���]��/:w[;��������5�jy�|��U��<��@Q*&D/�i|@|h��ݯ@I�%�m�Z�۶|��@y \��a��ʣ��7�qw7���k�;̏������д�)i,���l�R���l�����/���M6v{�R�:k�򽒘��z����ă����0:hB (
��_}����3ңk��_B���$J諳��5�����of�潾+�w��X�8��Z̶�d|�}�}��i�Y ]Dqhk�*���xjth;uW:�PW*m���q�e���w\:�UWy\�h[.�v"�����@i�GX�]�+���>�
p9EV�gS��o�dY�����M��[=]���1��8p:Smf�ծ�(��ݻ��+`P���H�Y;"�Wי�8���{�����*`-S�u��ڎ%x���Q�\�/]	��sW[X���o�1,���a��K�����[5�w�u�b��0x�j�q�9�%]i)QOo+4���MԍX}4!�ҵ���c�����N�4b�\�� ���:!mS�5���N�����{��56ܕ�Q91��촴۾� �C�<���z���nu���\��k�;�ma��e��W�Kա�e£�CTc*��hC�B��v�]�	@��rgjye-)��*v����۩Zq����Qޱ�[spgt��y//�5�:fJ�[ֺ�e�L���v��S�ds :F� �9�^=gx���ȩ!�����닙�O&���z��'1Y�h�Bnb3��h������Z���fX�Ȁ�� q��Ѿ�8[%���a��n7�+va�l�\@�c),�!)�p��d�md%�$�&FȂ-C
	�(u�L*�!lHca!�`�/nJ8�P�G
,��̭���k݄4^"D1@hv'6rccB6)�6�
�y�g2Q��|d?����Y�q&TĞ���s���ߗ<&f�j���M��oV.�n*n��WT�yGz�ht���Ǵw5�s9�5op��C���typ���K�3����3c��3x�n�Fޚ�D'���l[�\1�nV\��l��oEϋ�2�e��<���5Z�%�[!���Ŗ�A��M(jF����DҮ��8*�+d��r��-�\��8k.�w��I劈��f��;S\���.��,��x���s���/��wV�j�k�q-.�4�=�B)t)pޅ�o���a�q�����{}Oq�/����wV��Mo>��(_UG7�-�t�]JH�p��f�U�;lՓʊ+�٘hfЊ���={H��P�w��.ܙg����YVU�A^ikk`�^�ʝQ�w9%Z{�v��⚙[�.�@·�N;���gG��Ӫ���:ýc&��]MFv�[x���Ұ�\��qVL�Ֆ�z�V��&�.Nv]�J�Z�˱c*���Ke����S,��&�L�3���q�]���g�*7ր��LkgH��w�;���V�O�'9O'�~�o<isܹ�:�gm�篸;������Eh-�	�%ݤ��i�X(�4κ�w�'�ґ��EJM�IE2��vR�A�m8I%"wv�Y�P�9	H� �d �,m��x����l�O�Ў7
��(Pf[	Ě�2�H$�m�-�,��,�w!!{2�B��"���DK4��-T�b���؊�%�����z.�??"��4�%5HSQV�QC3�����-Ke�J���׏mk�O<x��1�<x���lud�Km')��
h��"`"i-��q�kZ׶�Z׏=;v�>�_���Ȣ���N+�4JP�U1˨�P{����VYgӧ�־5�k������v��ǽ��vN�%�/�yjHK��J��JPPEK��u�Zֵ�k������v������h��c�iiMU%�&�2EUTRm���h�C�����]4����{PQu��֋m�l&��64��i��,�v���)�[4�>Fbd�#���_�t�A���im�N$�-z�ˣl�I�4�	��jƵZ[m�h4���xA������F�����EN��?OX�]&n�#M�
g�p1}����2˕�o(-�\qS�<}9���w�&,����Ά�r#�u2���)����+:[�m9r�- ̀(�*�A�3�<ՏMo1��z�	�?�
�	
�y9�P���I�:P���Kd�đl�H�I�-��7��������h�G����H�@}��"쥹�����Ъ�Q����@/yNoO�}}�#p�ˌ���s���Z��v�w�8g��1��:��>Zk>Cw��.��p�g���%�w�<�����5�V��Ǉ֬Th1��c���L���G���>����t2��'8�W����vÅ֮��N;57�j�O�gC�ш����W �?�ib��ɏ�Hæ�~��Y��y�=�ƾ��UCL�W�g������%���3{<ŵ��.��t	��k������7��ξ�lH~S���h"��p%�'��k"|C�q��RRsdeJ�vfhx�\
o;E�����nxZ��R�V��=��}�LF�\�k	�M VA#n��J=L3ꃎ&�)����1"5�^wo����������_=�	�[�F>��Y�_��%��ȔB�M�M�ܮ�U�Q��񐷴�7�5�p����}�|h-aO�gƙ��1�y�(tH���8���>4�~Q�����]�v��?e~��)u?vd����VF���c�M8��j{�`k�eO�����Uӏ��~�^]�/y�D�7%�������m��QkV�엩�X�`GT�p޻7ä3nP��y��eOuu���;���]£a���T���w�_=�P���E�W�#����#ٙ'��{ޱU��$�8�I�q8�9bI%�IbE�["H���<����0�=�����bܸ�|�_��X�]yմ��4&!�����@������`s���n��{-F�e�Łe���wf�I�%���@e�ڜ���fu*�`�4��<<[����[�b���r��O�m�d<��&��I���5�x��s�����'�w7;���Q暖].VZ�����J����qN��NEG���ϖQ��&�Ժ�Xg��CY�}&���<����x`�����L#�@z��ϒ�ۭB�Ws�o&2y�y5��]w3C�;� v19�z�F>�w�e�=6~�]yE+΀��6<#��\ԋ7\��m�#Uv�����3ҫ�Y9�R�M�<>�.�t����Ͼ��{�zo倁���Xc�Ap/a7���`K�w<���ݴwO����˖Ͱ�1<�L3 ��(C�ޘ��(��3���|"���@s���ͳWsRŉy`��� ��)����nW�'��^A�f���ż57���i��{����ZyO�	��������5-�՘}��Պ�����T�}�6�
�7i���|��,��a�V�������h]ޞ7��]X\�o�4c�̡;�>�z��������� �dw��S[��H�f03�Q؄�GeoS��r�h;,������W�t�moj�O�l��_g^�sw>s�s�ﾾnK�!><}�刖�'�w
�<��<򂼰��H[:�����}y�|G=u��O���=#���!��K�`��콫g��[V�E���+�wJ���SVt����@]d��s�8G�6�aؾ��
�������X}�b�oC�,��M�2�<�\�L�'^����1�m <t���s�Ǉ�06:�u��l�-�9�^E��m�(k[Xkc��<�x|�����[�`e���������G��>W[=�ӫWee�1a�B3�����c��`6Kmx
d#��#$T9� �yͶı� z%E�@��;��<�%F���s�������/�T�{up��od��`�>�Cv���@��/F�|>>��A4��=�8z����^�a-����$��W�g���0d�H��QtdU�#R����ד�!6�ӭ�ւ���ffg�Й7�毝��-��:�f��:`p���l!�iDC;��;�ר�9иt4�x�=#�F{�k�L���q��ƻ%n�9� =6�sg�G�;�d�K���:5�?�/5|�t�`ń"I�ïD�"��ޟ�}�i���u�/7
�^J�Z�p�'�{q�UR2�-�6vt` ���gm~g��R�7����VMH�ʸr�_��w�i8m�{Ҏ:�g��:�T�C�!��m�iM��<ثU�w�w>�_Z��a��҈A:�჌���2{���r,�
�=�7�_E��%�M��t��v����2 4(
5���^�
�y��
�y�P��E�iiPJ<<��f����{Q�=\� �6�o�>6���(�Ǭ��Lp܁!�-���`/5��ɉ|���ø��.m6>?uz#���[��©��pl�hz����3�y��b�DE�=�}��e�8��QA�)"���9o������ ��D�y>F�Mn��HQ��Pކ>5+�2r��b�����#,�$�8�	�����#��@�5��{�-f�/pl�.vPs��Y.�����v��䩆�nj�����c��d�W���q0�L�VV����a�����K�mf��w9���V�NS������ڲz� �*�������`a�������1�
�0/|0�]������_�Iɫ��I;G��lag`{�&��(0��"y�{�x~uf  �-{�PjD��Q����|ܸ;ݥ�����ٵ��`d�<����@^����ᔄo��.Rn���+�����^ǎw��3��VЛL�����C��2D����C��.��5�c姼�]'�CK�]"�]��5����+��o�q���ƽ}u�8=(z��I�#J�AGNy��N�����>����jig��WV�t�*�W�A�C�>{ h�J��CG�*\�*���$�﫡M�`�,m��Ew�ݭM��
���L��b8]&*��j3j�ޘ)�m�Q�����Dwf�9ݤx5�״��ޝr��5��k�Aawc	v��&D!u���u:�s���,�pT7G.�0����1"b.TJQ�4�����n�v󣋿��A'��zA(�Py��y���B $�ZT �Q�

���տ{��}nh|fjs;!`��%�
|�<���dmxD Cd���]��v�0X�m��1Vҭol�&�&5��5I�(��y�I����#�=�f�_}.��_��l"�i����yzߋؕ�y���u�+W�ކ�]�"E9�BoNO�su?s�sώ��w���?�iDVm{�B]���	�������xX����ˢLX��������ya��W�#Ъ�e�-�@�`ҩ��.�eۤ��Ϟ�!	;�s��xK��gº�5�k>7'Б�Uç�#�[l��7��]e�d���!	��DЁ@t>� ƴ���G�`�#$\w8�����a�ʣ�f;�+;s��s�R�j���Æ/T*�JY�͋�0^��z|�`:����8"�-�ɀ�^k��s��z��>'f�䡛�t>��ev�%�B:1]q8���j�y��Jx�F�����MV*�G5�37�	�4y�������'���4������X�(�����}��ͳ�W�7>��!�+����4d�"aʺ���C~��@�}J��I ՛8�F'�m	�y��S�{��C��{o��V�mŵ*����o���8"Y}���}��,`�R�Xz參�a��,ʻy�:1!�4o:�}/*�DH���Vb��7�h�׃�OD[k*�/�t�ֳ��Ȼ }����]]����y����I'ǧ�Ȓ8�<��@4��<*�JI-$�iK�~o�Y�g�Ԍ�u6\��ۏw�aSp;�)��n��^�6�7Oq�l�%3�+SuY-l-��ʮ��V�����Q�}�G��}Ch4�������a����z���&�9�j.��q���oL��Ó��b����9oWB�p}�l>jam����~в:�,Ȟ�C��;�}����qs윸G5Y��p@��/y�����쎱���m�dJ���ǀ�Ƕ̞!{��ܭ����J|]�[;�<0��8(Ƒ ?6���U!��U�Yҕg�keՓ�>����b������|��=�rԁO�Te~{Ո1����}{��|E��:�"�~��&����ɸC�)�"@7�%͹b\�=��*��$søh�B��	ٻ����a��K�䆲��<�e�{D�P��N|���,)a�Qn���4�t��˄f������]<0���+�O����O~����T���%<y����{hA��Uq�����]��Z�K�7��[s��YE�}m������r���'���G�Tӕ�����(m�	hNص�R��{�ѹ�Cly���1Og�]�̿4*�3�߆�ܔ��#bƫ��;s9�R�Q(�]�+��F�°=�5����r�uU��v��'���^�|�&�3���$�,�*[!+g$��8'*"Wp�<��(��H�@��о�)�]�x����4^�@��%@ǝ�u������&�A�D�O�'[�o{YB�vP�*W�<�37�}s��n��a��>�w�a�e�IG���Οq����H4��]s=���k�IĎp��_bFb�=N��l$.a˃�uV�5���ѯ��{��UG�p�g��_��U|<>bv�4��6c3��a��j��ʌ��}��o��4=���V�C�O����ﻝ*liB��8^���/�L�X�K+�2��O� ��ܗ��`J�'�1�A�2�/��(v0ҚV�eC���@}��݋a�9s��e|�� ��F��x�ϼ6U����l�Ei�����{ڤ���W��-���X���1�W�Nť<>xg���Ƥ��wC�Q���nEmż�p�My݊.�wIa�]=�.�{0���e~N+J�^|���Ex�(���Kx[)z逗�E�[���>�ؖ/�F-�������p�l��|�Sc:�Sn�=<��O�F�������q��zה�½��X�_����D����-�d����x�+�<@����u`';�50�ff��%�!b�{0t\�J\)	��������]+O$K��9��sz�m`��S�N�W��!��ϻ�]��ս�K�d�w��g;�O�k����P�j��'��ʧ<��'S�<���� %�!H��|�=�v�=�_���M�:<��|A<���9����98�Q��(�r�W��8��j����]z_8I��栜K. �v����`p���y��A�l��_Ouy����zz�)�fk�ﷷ��Zg��"�Km�����cޱ�]T�����'�0���#)�A�]X$gx��'�s��wt��Vp-�̺.y�����Γ�?S���ض#`0gF+�!)���Uە�����k�t;o�����03��j[�ݝ���3�W��ۍ�{I\`�+,�>d�7��t�x
b �l�d�&�|%�XG������J�|��U��	��lFKA�Xb��m�+ H�&�мG���`p�|i3�������D����>��p5G�{ÖW��/���|KD��r�JX�2�|g�ܵ�7sЗ�zW��<�09=ԝ�������`�e�@�����4LP��
c�ڵu�%��y^}�*����=��x����<�u���7oEg�&Id�b����А2)�0B�Ъ��q�>Q�(8�D>���'���;�\y��M_�}4s�x�T�^�˚ϐok�(��Ve����]/I|}P�8�f�H����k1���$m��
���E'{yl��ݚ�����
JP�jx��¨MӴu�Na�A�E�3��m�",�w�/���ʐ�RD��&2��"��-N���z�:��e��Y��숯����<�ȧ<��'D��������ċP\�߬�߯>}{��oԏ:�ϴ�L;g�>�����AZ��t
S�)�z��[�z���w;͌@έ;�ޠ�+�DK5x�H'}�M�7zF�"���5'0���4�`�P��A��fDl;ּm��5�:[=	�߽"�&�P.0�U�x6�{k�LK��%��Kr/�r���&�c�VU����mgʁ�Xmb�k~t���1�t](-i����
::�H�L5�8��}����k��V�T�I�>����Ű�ã��G�M�	��=��t����ة���7۝��u��s�9�O��jy5��a��s<󧴩X��|pu��RݹcO��>�����;ձ-�3dL���'/�u?s��㸄���!��_7���5\�1C/�^��r�#�r�E�?��Bz�0%��N�w9�'�'��u�y�y]H��
}<`�	�#�&T��}�o�-I��a�jD�$�W�~k�1z���#�ܞ�HϩD��/-�ǥ�mwj�<�����d�遭>���G��y��I7���.ypҹD5�Ϯ~�?}����+�9����dl�&��u�w�Y=ה1`-���b�3I.�E󏪒Ă� �Aj��"TL�Q�$�$�G�Q� A�_Q��k��t��Fćyx�_��͔�k�_sBc��$�e��U��8�.	����o���6A?�U"�r�S�Q4(Jy�����y�C�y�$�I$�--[	����߯6yϮ��������3�`�,�4>�MA��5��&�9!�ʬ�15jN��+~������9�]}�$�̐�������ͣmA�)�e�|)���;������f_/3dޢ�^�ǪVzD��NyƆ�z��~Zj*�3R
/Pu��_z_��8��aϑm�����@�5�8�rq�A�����HƄ��ҩ��D�nv�tӭw�:`s��S�l%���:f�;V8A�܈e@$kY�Nn�n��f��z{)�T�C���oV<�������d�#[o��f��[�t7�_�c!��A�����r��$�9�����6=ܚo��V��<Ɵ��u1����qM����#1���m��t�gW&�~~�-��IPk�p��]�1�S�ȶ�C
��������n��d�r_*��Z��o�7�W�G�`�p[�`��{�(����%���Ք�1��i�5�$t�R�x�&Έ5�p1ӷX�LZz&�f���Ϛ۰�&������@��B��k�I�t���{�MM,�ώ���jVkq�ܬl��F� #sfP��gy��ت�Ih��}yl���ѐ����M�v,^Y���]��v$VOM2��0m�<7�KN�'����Ζ���Jm ��w���B���|�6�V�;7k�e�s���&>��B���{�|��(3����Fȴ;8��(;����-�p�Ց�޽���^�EF��ЫvH{ٷ�\�Ⱚ�3��֌��/�*�W����I9�z��{9���o0�����%N��v��y��5�f���Cv����#e�c������ʤV��/Mj�خ���[��R�%��PqX���+��t���ٯe"�eyyߞ?��Z���՝�����rm����)J�m��,%��bd.>���XX~<��c�'w_[�ѝ� =NP���]yV�'w��}v%�T�j;qr��,���r���X�k��I���A�ˊ�!�զ�U�X�����Ir�7G�ގ�P@z�����<��P�sHӐ�jrD�iz&WB;��1]��n3�k
�:����˪72`��
��wU�N/��-�+ ��-��J�N�=�͝�wYu]�/��Z����r��	s�j0�hVH#w:�����h��g��#��V晵mZ=ί���S�-�Z�G�%���0)�mm��6�e�Qh�lt#���T!��5�vQZ��]��c����P�����\V�,�c�����\tȊ%ơ]F`8*��mH�`g/��-��g�1�:uض%��4ƙ8�,v�`.�ے��ib�N����zo��&��uV�l�Z�Y-��w��	Fw�)G,T����6�ݳB2�#X���,�����n��a�]�A)�Cy}�^^󵕛%5�mp�i��CT�+\/b7C�1X�{��Ѹ�fM�4Mү�Z��H���N�D�][��u�hG�����	�W�5��U�'QW�I;7����/u%ؿ�7�v�^Tۗ���sqN��_�����m��뷎ԅ�58K���WURh/_4�����P��7*�ԩ{3�<R���n��4v�*N����d��ʆrY���(R�ϧ�m�N�S޸�!�JAD��Z�N�g�]�{��
�7�Vr�u��j�Ǔz$ï��U]J���vuV�:��Z]��>�7�K+:sю���V�r���7{�rˠߞ��^>�Q�(��v�((�Q�$�_}#��e�\t�۶�5��Z�Mk]�zv��Ǐ��Ovu�]v�b����8��顨�]N�ԲZ����t���־5�k����=;v��Ǎ�bUyd�_���.3I@�m��`�y���Zֽ5�tֵ�ǧnݼx��X�F�G�v�x�|�����KV���c�kZֽ5�k�k��ONݼx���|�|�|�M�S�tuT�tt��!��I�렮�%k]:���l����4;�H0�癡�饤݃T�Ov+_���ytt��%����Hi:Z(��]�"t-m�^��t�l�)���Ƃ�I�&߼���KB�SKU�6(:�Ꞹ�i�C����@b@�"����S,,��y���c��GSF㥃���3���م�x՚�����x�����*��-.����u��U�t�,�}���	\q�'q��%q�$D����Il���}s}}o��>�jt�����)IX?�O'�A;��# �8�9Q��zY�q�S�Q׎�m¢sk�247��u(r��S�i|^y��mXoM��U��
Xd�Ue�����z�,�gu%��8s��zt���X�"T��.G���>���;��:d]�u�U�{x��u��O���2���ε؁ �`���y��C�-�}�����=�~B	�z{�v[U�"�;�3�vgY�t���w�v؞~N#	P+�A�	�z	�2���������O�A���ϫ;w��ó�-���<�u��2�����=���P�y1��r��_��]Ry��z0��Y���q]��$pQR5�r���!_@�w�=�2�s���3�7_�$����N��u�w���6�a�W_�@Ե՚�ܨ�^87�a�#X1g+U�3=��Q���\<�@��Ra{�@�e�k,'qS�;�[Y���11�7b�ϊ��T��{�j
`��n�.��������%�����$���4D4�&.y�)��q��7��7+�ޚ��[}qAr�0��T�]x�S�p��\<7�T�}�D�=B�u޵�*�f���/w���l���gWG��uU�t���y}Z���|&�KI�.��n���dm�C�瀒��rD�q�T�ȕ�H�q�"�ҥR P�*d�}g�{�y����;
�����Ю{�N>�[�Xe�p{Ҍ�����!^�g��Jj�Z}¯��ph���������Ú���B�"��5ퟞ���Wߧ�:E�T}��u,�P�?R2�!�k����p�Dy'��bX���ܥ3y�| ͗��l�O�v�+z�N�oT/�!�/���h�qCѨ�1��G*��\�V�]��m���d��V�Z�1�e,����]��噃k۽4�G�"L@M�a��+o������'#2P�]ȮՖ���c���tǇk�u�'�3�����#�B~��q�����a��<x�M��-'v8o}����M��n���O�Z��׷ <tk���D��>�
�yi�3�)��+�W���2%��c���>��Q��B������+�u��+��$�2����y�k�w����6�׌�HǣR������g".ބ�n�l����#�"0/F��<�c��f�p�ZG'�g�ۡ²My�t�mvb�RW~�?-�ٛ�XAY�;�lrݷ�'L��G(W� "y��O\�	��T]� cx��vS�̇ut�˧uM���2��J�>w�h�M읻�ܘ��7�z��ö�윻wD7!��+7���x57;JUY��{&���,�ºQ�:�(C-r��д&F��C��I����� ��I&��:�\q�"+�8I�r�(Q@!H����������~�sٹ��%��i��x|r�E�4��.�B�PO�>���i���:�d#ڜ�I�
M���hڵ��`�,�3w��on)ʺ�����0���V�x��f�Vd�a<H�m��M�X��c��Oi�mp�Q���C��a�X��S���k�cČ�ZE��\����E�h����99�l��>4��d�fv��S�!�[7������cMjz~�g��N���2�Z;�VM+��y��?����>�f�y>\Ez�RZ�dO:J-���;�x���+�e,��<�Nf�2nv.�z� ay쀟�׎Cv$�)���5u
�y��釾Y|L�����ol�da��Ԋ����a��8�T�.5����^��Iuך�8���:�&o�{�[{U{m66-�'"��ǨY_�Q����XG��S�s��v���C�=Wo��}Û�M=o���D�Ut��~�ż�q=�Ԙ����y��p���B_Ͱ�5�lS���+v�/�媢��O��~�,S߭)�u����6��<@w6�,
1^�<�L8bf&���>�Έ�9Z�p�؍:�T}\_)Ҵ�u}�k���"��i��Yu9���{�k�ъ1����zg^�Zغ@�>�!��=A [�^v��{������/C�0Q����$x��n��U�ǸV�WPV���M�k{�~������%��8�8��%r�0)�(Q5D�j.�<������?sЕ�VdM:oc �n����6;��IV+(�������h~��y�'�}��3��{�0�'��C�9����rz��,ɓ�V\�T��u�8��x��'�_Q����d������ù�~��hrbz}����ʰ�¸�Q{�W{�lk��Bbh`ѡ��W����P���llc^��_g���y�o:o;n���,+�7���R[|��i0�Q�D�G
�Oҋ���~�և7u3��"i��/��v���:~
�8��׉�f�yE �3D&-,�<�(ZLx �\8���G,��~���D�}���!���ʟ�=7c��_�4�B ����V=�=�*߀d�զ���b}�j�ՙt��?;�oeF�ڑ�/C��{��U��))O����4���"�����i�]#���4�{�'VFns�W����%���,���o��2w����څ�Pip+��l�褧s����Ϩ��?}��̉���~B�&�r��>V|`���J�B��P���<��N�_^٤�?gDk/�;�a0p&���5��;�r��QQ��v$�`O7�����v���+�Ha���C�q���lL�QTz,G��U�>Q PywB���s�tJ|��z������ߤ�ݫ�I/����R�+�q��9�Y� 	��_]]oR:��P�z���J��9�8��+�8�8䜰��Z-������<�}w�����{������4�-��k�� �|i�;�/�1�J�짼C�w{��-��-�=�[p�`����4������o8̜�D�/�zkD% <}�<��O�0���_�PnO���Ր �Ll!�2��/�%h�~����{�U�m�6+���s�~}����~/����G8>3���s�Aئ��ǵ<��f���ȥ�62l۝��g���m%�(/E_����������M���Q�ax.9��A�,r������$�U̝�I�jp��w�bwǷq���>09��L3�p�~�]������̵;�z�f1���&�mr��7է�WP� �����J�a�~=��7O�����=��Ox{[��^�m���xˎ�<_}����P��.Xo���9Y�@�_~O�P0����7�����*��ާ;�r�j�s>����s�P'_���`o����{^��Р?��|��+��$�����>��&��;1/���]	��v$�a�k�J-<��+���֐�y;��ڍ��{7c��+N,�X5���L(�ώn�'�\��Y��)��ȭ}x0.X�pg���w�p�v��1ƴwzS��pЛ�7����e����ՙ�k6H���nG�d�B����2�s����|�:���}�UOO��8�H�8q���d�[$K$����>����w��]}���x�F������np��ɡ�-��#n����4���n�R�V�3�@�ӻ׺Ge�~��x�;U�ft	��/�'`��,^�V�b�j��3/_�iN�H<n����U�ӗ�G-�����c֠�`_}�B<���ƙfϞ��c�;�[�o�
�}M�?N�ڂ�f���*�t:~o�!���3`�0�����+)��`]s���ocY�e�7�|�vdm*�s�(��(�z�o�{g�;�C3�cLW �����N��¦Gml��S[P����ms޸G��Oz�cٚ�l�+X���qWv%-���pq��>T�/�[ ����(��m�i�=����V7wT��d:�ŏ]9Ǎ��=2���'����n�5��F���
EE��s�~aA�]9�9
���_�'sM=�k����б�W�d����2 �W�<8鯃�����\�q!�J�d�,�W�K���^�����������W���W�h�YR�Lm�n`�"-��?uh�"7�q��/�ّo��b4��T�xJ�B=�$�+c"�*��������w����ޟo[�z��<��Y+��!)2W*�T)R�`�%1ѡ�z_��<ӌ\��%�TzaͶ'u�[��]T��Vu��v���WҸ>�.�E6�0�T���^�!TC��h�� �1�Tl�r��s�U���D�� s�;�y瓉�4H$D5jKܝ��={�d3M0GH�	�E�3~�8���Y�~��	:8}!�Bzw����y������Z�u�۽���&a����L�#'�n��r;�'�{y��
0	B��l�����q"_I�ܹĒvn6c�;s�vf�{��eQ�^^},���wO�^�sܵ�nO��VHtE.͠s&J�7!��VzC�w�0��X��u6��偬�߶�|ȣ�ۡ¹���4�Ym�fg��ޭQ=�a��\���M-�^#+�{��L�dZ}��P-�,�z��g=/�K��7�7��=^�1����)ՠӘ�^�K 8< CB���t��R�o���:i�wfѾ'����i�v�a'�F����Sߵ;T^&R����l�?1�ۻ��p�1�UqȭF{)�1�ך}��Su�l/,!	89}挣;�{^��ܤC�=��M�ց��;W-�ט�
t�a�F�J��7S�\�U(��r|�5������"SגS�(#��1Kn����A4��i�fntW��@�an��V��ӭ��Y�A���^�n��g��a6nꯦ<V�]�!+��Y󪦀�`�{0 ֽ���W�.���Us�BӺF�m
G.orVcN�9�եvu�oW�e�	9��,�;������8؁�cB�q]'kW:��!��9�ż6�f`{�y��Y_��t��b��0�ӦU�7y߽������M����Җ�(<�ד���C�c�T�&�!�{�_3'�&<��)�Y��.q�ƧDovsko�l�Ǭ���,=��cH��!��<��af�;�_L�V�D�Yۮ;�;'���LRc)���0ut}�ߛ��I�;!�7V��")9�
�M����;�'�٩V��>q�����U��nO`+��=�s�y�OjyKf�H&zN0���t�}Z�������:�qn	�0�~c�رF%�"Yُ�`֋/���[���X�s㸄�8郰���Y�qSs����g�zz9�0��&�������p��/]�>��=~#xPE|[�����ЙM&�$�M�U�f��`�)����S4<'/����L��ݟA~����3D���1���֋Q����3:ҟm�
�q���߈/���v#���Q���7b�\�j��ͮ�5쀻��6]����������X#K*h}(��W��(�k��}��8�fz�����6u�������LIza�4�(f��P�}�s�)_���֭�˽u��zl��zZv%��L*���o��R��T���wÆٶ�)�ŉ�q[�׭�/��z[�W�ZY��F�Wm[#cOM�-��O�r�����!gw�<��_R�����Ovkɴ�E��u��"4�5����d�N��99'rr�q8�G�����r�v����D�X�O�^�J�od3���ew�x��t��ߕ��<�t��M��q�H�pf�0i`h}#���N�1����HM_7�_��7�#T����ɕRr����'�~�1�yxĬ`���}���d�	`L�Κ�����n:��l������^���>�A�s�6��yYV�>_Q��Zt�ZUg��$O)ٔ��N�J��7��7 ��Jm&�t)L%����Q��y�����C�H�ϑO\��f쩍3�ַ��G��nlXx�.�r��,Z�����UP���e�k2�Ǝ�8މ���x�9�n�k��+���8v!�K�����`���s�m�h�7���|�ڤ6�k�Fc�������p�����4�7O�����ƛ�<�����&�`s,/Vd=�_	����9�y���0uS�>�5��D�����\u���>��>���y	0y[���_6aV��^L7	G�kR�~��=���HM�}ֱ@��{�0b�\^S�J�f�S���),!y�)��?��w�<������؆;�V2_N�*��������N�'r#օ!n���ӹb݇3�Q�D3���|k�����^�U��ͼ[�N�o�6�i�n��|���pYJ>���y'��=zqR��̏hU��rNY\q��9$�9q$�fo3�N��������j2�U��a+�V�V�@��p�\B���@���cMnT�P�i՛|8�q�c������y��IeṈ@`�'�3��-s~�}5D]D�}�Ӗ��<<C`���;2�)�i��#KlJ}J��_-��C��@m��1�R2]y]V�)�{��Ax/x<����w�ۇԾ���{�m������z&�]'�<sk{o��2G�����Z�Z�h�_�P5>XB����E� �@nAޮ�>�c�;�v�r�by�$<��N������{%|>}�w�{j�^�fb����S�Z�ݗ�W�ӳ���l�XU{��H��t��1qފ/L���a�z�i �%�]���ϲ�g/TO*<+A����o��ڂ�_;!�)v�B��64�	�p5��-���Ž�xQ~N��@�p{�N��qA3вj�̞�,�S��ȷ��E�S�X��v��e��!�μϽ�w��2�f�uH��pM�����,���Ϸb���L9��]�ɼu^ , P(��gޙ�\�'��0c��1~:G1�R�\܃5K��+U�qf+,^�C�H4�S�E���r���M���7b����ؠn�Š�[� .e��hQ��ټj��F�^6�1¶�ye52�2Mldl+��=F��N������6��X�Ȗ�֭�+&�i�v���E��۾�v汗&uv�Yw�L1�kK!R[���l�U�]K.��qP�瀾��3��,[��<��1�/�=x{���G�E������4�>��j]N|�amhnv�}F�9�V�u}�m� �<9"�G��������A����q���B<ҹT�V��˅�ђ=�Iە+rG.���DK�"'즢q��_j�w�|O]d�Z-�H���2��2�ҝՒ[Q�x�Y������X\��_klͭ�]##���5d(��rZg �����6��-�������n��m�Vw+�s�;����o.�b�9	u�^��C�Y(��-�VT��O��ꤦ��O`��AI���W�VW��m��ݺM�+�ս�,�6��]�*�ו�1{'S�nŃϯ�WU��b裼Y�ޮ'��e�⹝�F�a-�3:����(��Z�Z�0��]��V�5��P�;Ԥ��6i��&=�"Q�uE*����Xn���(Zǎ��U|#
����A���NF&��[ɗ�fd�':��G3+�G����ȌV�m��yאU`�L<�߂���՝ۺ�����\uͫ��Q�\��/*db'9^'H�5����������6�SH��E��X+V��.�G����_>l�ز�q�����Ի����㖆īn�s��
�m�g����)9�ͧX�,)�$�p������h|E
���<��j�sz�uu�w�����eB <x<�n��*=u����d���e����|��,��V w�kf��u[ �b#x4\a��&��[z�3����4m�7�P����!%��|u�VU6�b��Y��ܝy�*��qK��YR��gq]�UȎ�u��xE֚ݨmьp*��X�2nn�N]b�5W^�Xj�	��C:�	�Ѭ��r�u���awn�t���L��c�/����nl�xs��ŭc��Zj;�-ޙ����cү�Of�+q;@���`)6Ã�'�����0��C���Wn������3G=��'�[7U�V�׬�Y]�P�y.�šG�];ۉ�|�Y��_MUrPy�`�i��?��k�_�#%�g�>�o�!a�wCo�}U�L�S��%��r�P�b�|�ּ��4mc�����m��r�wS����i��xw/�G���nw�	9IZ��ˠ+�F�L��q��)f7lӬ:a��͗E3+�%�:�*���h��7�L�m�\�E�V�w��/�s���xM��Pu�u!��C�gu3�.	���3)�j��������ҽdZv{�O�����]X\�hml��	у��i9��]k����s�/��}��no1�n���d�Bg:�ks{�˾RVq
Г#ר�ipݳ[G������Xu������8��ޭ��{���TH*X�A��L�a#��*�.�$2$�50R%C��)$�q:�Ÿ�F�`�j@�*�� �%B�H��HF
�:�7,�tʹM�"`�I�	�pD���1�m�&S�)@bz[A�w"29!�d ��f0����ƚ#�*9�BA���	#'�@�0�f��7Zľ�C�4m�`�=��m��:�U�w]��cc��Ƶ�k\k]�����x��S�l����h�_`ѡt�(��H��ެ��ugJ�cZֵ�Zָֻv��۷�>y<-�՗����NA�h(M��	��):���Ut�k�Z�mkZ�Z�}?_o�����~+���RET��%��8��j%�����d�WOƵ�k���k��ǧ�o<l��y�r�哒�Υ�� ��C�"m��l���M��7̆����R�ݡ�b�(t&�����T`(H����&��ih4��E���ҧK���������]51�յ�LC���l�j�K�TP�k��ժZ���(�PP�Ƈ�qt�ci)5�T퐭i�.�#��\.��M@S	C��$�K�t�/}����8�f�}g�0���yM�D#ė܂J����ꄅ�C��C��2�qq�v����ύ��HX,�"�C�(��!��Y�$�j�2�z�t�Ӫt���Ӧ�Gr�=�>����K�x�M8S#�\_�\I�
�_.����(�8���NF�1�Z��~�l�o��r֓���� � o��>��B��o�p��;4 ֍zCV�w�y/�M��OzyxatVg֣������A�+0��g��eЃH|s�a��~�}�lz�����U��^n�O]��r����^w�1��ǜKG�c!��(c@�#Y\��uSWMV�&���Θ���zdU�4ꗠ�R��K�8-��� ��dD�i��ϗ1{u�#�G{CBs�bX�zdKt�I�8���t3�'�{�UR2����6X��t�\�]e�iō��*Q�����>t }>P�[<ՙ��|�`��s�	O�^�P{�S��^�<��E��#���l�^�����������|/ݞ�ѐ�.9>P/�3)j�6w�O�s�ޥ����z�2��D�t޷.�R_����s������M'�]7M8��GF'�|n5X��z����}è�v�]�A!�,�_{-�3@p��S�ŗ_zh�L�}��E��a#?)wy�?��CsNNxȊ�vn��θ��5�m�I�܆N����V�u���7&_�l�~��5�ۺǝ�+�K��G�oa
��t���jdr]'Jι��W�f�����ɛۈ�+'�ӯԨ*T�R�J� Ƞo;7�uO]xo|�,Q�:�܂�&w���e$��q_�z�&g*�V	�e�3�>�~ua�-�٭�9����.=ѓ�4z ��[�@�D��A�LT�y���{X  ��9�k׭�e�� ��}ץ�tӇ�p-0G���x�<u ��>�<#�.97�`��3	�W�Ч��_�j�tQO׳}��>�+1չ�	>��08FFǺ���JǹJ]M@t�� YϽD���'���o
t�_&\j�U( ��c�թ�]lҁ��c�p����?��)�
�e��9ј�3Eba|�-��.R�^���<��x3�Eê=?����C'�{N���vi��J4�M��#��Ȍ����G|1��c����|t�2+�wR`�/IF���So��/l+�G�.^7�ʅ�Ʀ��_��j�z����nY'I뜷���5�T�L$���hx�*���(n�����0Ĭ���뇖3�J%[����������tYo?6;���hIY����}�/�;]4�A�ի��.{�(F����_L���8X`�B�f���^��,o����ߛ�ʯ���J�!����\Lװ�c5|�䝺:��{�})�!�F��s;̯l�Z�.������<�u][�����ٛ�-�3�tw-(6��Is��J]�;�s�,ck�� *�N�*T��nk�K��|�� �Ż�^wA."�y:G��(ӎvO�g戢F��*VԿr7��b�.9����3��:�?�m���D��~<�P~q�|�.���xgA!�n�"��������g��c�M;���4ZQ�1�LS|`�`���e�/��[��#�o�g�%�?��>1N��@

͚������Q�)��ݧ�wQ>9���"�
����We
O��h��1C�[�Ys�o;�Un'��*ǃ0b�'�j�9���?mёc��
�OC4x�5OE��3}9ݵ��x�	��y[�Z #�h;�范���|�b`���L3��B^��%{�j|wE�-�*�/'��o�a��7��utį�`>���b�.�1�ld�����Ammy<k&&zOhn ��<|Ce"�Ε�bdv׬w���8"y���	�[sN��8�3�|��5�۹�6�އlU|�W\�&W��ơ/�6���c�A����{m�}�Y���R���~�L��Ey������Jx��}�J {�{�^>L"W5�~뚨��A��X2�@孻�a*�$�|y��ПH�=<���Z�w{����d�wrvt���7`��tV,��W-�3�V�TgmS�>��/����v��휔���ef�ɻ㱳�u��}�珏�����D��l�_Z���c�������^�:�M����=c����g���#�Ջu���|a�����sv���/��G<o��7,_�S��7rZ��>�]�mNOS�C�e�0���'�i�|����8�&��$r�\Kx � <����T��I�s�$H�]e�"���Np���I�P��X������za�3���{va�[H�
":;~c�:�/mN���,e�9ћ�����K+Ԙwi���E��4��gO�A��YH�=_�o�wLMS�Ó<L����Z���υ��A\=����I�uAa(��Q{c&1��yڅe4,<^6cQ���#z[��s�fܛ�a� _t���/�i�(�
�ZW�`&��Z�39��4٨��˃ϟ����ɤ�q}�2}� �NZ���͉/^&����V��:��j��9���V1e}\w­�6��G&�dΫG��o���6aOr��j��9��{�������z����i�X�	�X�>\�ʚ���7�UP݅�e�ͻ!I�\�����7�Ջ�Y�|��bGq[�ψ�41���n�r����F��5죗�]�7Eʭ���dxI�/,�Q�ud#��%D�"�0�CHn4XeYO-݂k2�	ܥE���Z�K�Y�{�U�WM�K^-](�������3$v!��Ǫ�Wf'ܡ��5j��Q�7T�L:L��bB3B� �RL���R�J�*T�R���6=���|Y�+�Jj6� {���|�׻pxs�M���mx�ut��X\D��>1�f�"7�.ms��g������B� ��*;��2���+��vt4w�A[�PO��T�^x�%���7G���+�oQ[�����bqe`|"8��l�3��sv�~=y6	�^����Y���/}L�e�WҢ�b�߽���|}��c�M%9��v{�|��|��^�"�obK�ҘsP��| Nv�vn*r���ʬzn��+�6�T�!�ϖ4>9Wt���(�0|j��,r�t�M���Fe��s��	m|E����d�.����ߍ��qr�u�H�A/��S�S�;wK���ׇ ��������K�v
��g�-u�;���g�n�!���#�A�JTrf�J��ͧ��W��9�I�ѬS��{��N��!q�����Ǝs�����1��Tey���ۻ�qthU*�#�B���
���}�to{�^Eadkt�uW���pX������"��"B�P������})��Q
��/����LȖS�{�$�����=S����P�������߬���ʹw�)�u���yad�A�n`7ǱT�V,��V]��Ա�����o����v��~��mK�Q���}���G�hFxX"��
{,����guev�#��yѦ��/���*�*T��N��N���La�Itd���p�����fft'vj~m�f�y��L��N7��9�Q��u�z��=&}��#5���'s�/���C��ΠL��o�\�5�m���i 2�3\�G;�'��]��\殺�g�����J[�emwC=�#c
m1�GxA^�mD��(�r&w<7��ӥ�@���l*�z��)�����z �H*k��V�X&;k���z<��Յ}�����gkx�[�k�Ƅ���LAz��'�O����3}��H����N�/+�5��!&��Ұ��#�v�	q{P�����t��!�i�l�&�[T��g�fCtsRm��VG�0�h��W��:��,�au�� �u-T�	h������ L�IZ�ħ����ۮ���엻ٻ�1_��i���d9�XxaW�!�4�祰.��-�l�wtӉ�[|bMI�e���3������M�w��+˂�&�P|ï'�b?��/`Q\��1��f�ĳz_�ok�}l�lO�`��wK�Kq]��l�z��E���Gt�/��wf󧶮D旤�q������@�u{�`��Z{]۪��]>�(�gQ�"�T����1�C\R
�$��i�b1�`3k5�;r�d������,hc�!c�b!��,���w֧H��'��u��on���>��IN�^�J�*T�~N�����}Ӈ�6�e��O�7\d���v/�ҐȮ���Q��l0�m�U��`�����m�����F�w�D�#�G=s������E�����z|6��0��L�*�_vA�4&��	�k�(`鹽M�TL��)�0�D-�m=Q��
&�p}&��v�;כ�<��b�∯ܨb"}\|x��6/��g]d��ݕ�Xor�����oY�=,���cJ���N��5g<=�j�̐s���"
�.�r�����G����WN��TJ�I�{�r�1}q���`��1�u�<��2�^|_i��m�>g��Cx4
̚a�x���'�:+di�Τ�y�Ld0��f�ئ��䨴��wĒ�|p���ZPű�L����r"SeI��:hj"yʧ�xvy�"Ӕd�co҄�������+�!���:��t�秨�������-߇�cJk���/�]*������|�0pb�fov�;��`�	����eo���MI逜�k9H�;�#`L��Z���O�B�C��]LX\2";9�i��=A�3��֫q�Ķ���_�M!.aΓeq׊��5�ܨl�W��K��������G�������A�ڦj��� #���]<j��C�_k��ԝdS<9:�wF�k69Օ�#u��Z���]�|��f׿����s�8�q�8�9b��������|���s���=I쪡ȵ|��a^P���1����VhXx�ݼ��|N��-p;FNwn>ur>r�3��[�%[O��#�������A�q]������t�7��{w��F���ˢd���K�;'��N�����*��N�Kh��9>��{lg����D7A0�����x\Lrxὢ*E�~mק؞ub�8WM�1����FͰoI�o[׬��]� 8�U��*[��� ���aC@����[<���ߛ`�	\��T�Sk#�����u����M�DJ�*�E�C�-�����-�c5�^y�&)��-��s~�g�zҧ��<;���8�ɣ�ݗ��K�%��a���<6�窾bs�&K4�����v���ż���j�E�_�2C�T]Dy���� �>����Ccy�8���П��)c-�q���Zp+[\(�qT9u�G���θ���H��~�aᆅ(������V&���x⁝]05��2(�x�pN�s��	=�t��̶#��`�8aPcK(㱱k`��t�iM�r�Z�1k���efR�ڡ� UA�2�sNG���X�t7O{z�=���Tg��	��xhUXCh����Y� ��(+c+kY�Z�Ŝ�S�P���Rsz�S����6����,�:����G8�z0�G��^�7��@d�Ɍ ����P�Ze���'g��o�8��q8�E��y��9�;�s��w��PM��+�����,�b���M��~#��~��r��+��-���ҌАmft9�ы��8E*]�`���.�{��#'�S�҉������!w� ��@Y>��ĳ��!�+﹛��\�}V�:Ѳ�R�ӝ���8�@���.��>�+a �,VQ�I����DM�W*�����q�q~]C^*�<�	����y�>��m�WoL�F$F��<xݢy7y9/5�Ͻ>|��.�׌�WI�e�I��=�w��<�Ģ�0F��8Zs�: 5_�F!��P�̭���]�-͜a71P��3�7�J����R�7�pEų���^��wR���c���ho;0f��%Bj��>���$ވ̊�Qj�Ȯc�������!	�yiM�𯐒�\c݃җ�[�(,K8
�s�/�ݿJa�Z-��DFc�q���`�:sv`0rA��c`���p;����¾P�ir�^~O&4
�H��Q��;���\�#�s���c<��ߡ��A�>�z�~� �B�ۯ�s�&^a��Gμ�<�¹���ٮ��E��U1z.P�ǜ½O��V)稿4�uX=oɕ���po>7yf|��Z8�[��ۺ;{J(FA���dK���dS$� ��Mc�S�CE�U�vs
o`��7���g�*����zM��aj��&�s Ӄ3�!Ø�8�DDH��Ν:lN��N�S��Ͻ���z��s���F�J`۟��n�ګ��P��58}vji:'�&��D+lqޅB���M��M|vD�zm�oT�P��9eΙ.3�t��)A�R��|G#69�t��պ�H�Y+����1�_)>krz�8
����%�3��m֟��)��?b�<��T�������8x�Hu��a� _�3��;��:�A=<���z�^�ҏD��x�v����k����(�b�A_�������T#�d�x�t�3�\�"���e�����^�������7���G'�!���h�Yjo��?T���ޮ��h��u����0w��m�����2�a��4��W������|�U|�^\�%|�95���Z	����uކ=~����f|P ��4چ����
|&�t���Uq��h�9cUs�=�c���y����/r�a;�0��H�2���
b��N�z��z��ub�Mş�G4��0(U�	D�Z�$T��_i���|]晠%�d�I�D{˛��%�brZ^:�uf=ǲ��yMEVu-�-�q���w�cN�^���9F��^��n*.;�<��#��ɋ�wvKOv��P�;�ۋsr[���d�q܅3�R�=��u/������(��7G��j*(��.�ܤA|I�^ަ�rH�z�7�u�jK�1�z��|8��{��>zPOe��������U
��}�fD�*[i��v�:��Gb�1����%��b�H0�0�|����6�=)�hE�:��n�{�x1Wy�8��%���Xk�@C�;�Ո]-�hk�n,㪊*_3a;l֩0�5��6=w$�['V�2'B>R�K��+p�#�Ee�P�L��\�(Kn層^)�a��"��h�J#���6�&�lG6"L�x����:g���b�Dv2�s�<��X3B}�3M^s��ؒ��X�)�I�܅u�f��f,�f�%�����ͷR[u���+�Kq�i=�ϗ1���+&�[��m��!bR�C��o����{E��m��V�)��7��N>����R�״�j�ޮ¡a�-��Ϣ�V���YM�Ə;�~x��U�|��"���[q�����p���.��$*�[/mLފ��ʙ[]-q�:l�\�����U%(�/�R�8Ԯ��W۸!��e��#��[���I(o � $&(]�ά��0��/��Zj�n<ah��Xy_���	�m�B?���w/�'g$�*��vZ�I>;x�ɘ/F��tooM��æ�X'8n��, �U�W^�ģu۰��]˸� ͽ��6��]��K7��T2�e���zv�4��䑅�Ψ)z[�c(�t�|��*S�.���N��\۹��R��6;���ǺP���Ū<n��:��}˦޸�R]���Y��]��(���vsh���]`�NuYkF��{�̍�b".�.l u�.=%,�ܝc4�7�e��vy�N�#]a����:ήug�ôo+G#�.��z[��B��m����q;���9�׮���_�����a4�WXyct�d�l7�]���ı�fX��a��"7;`ڎ>7�Bo��~��u�G���%�w�$��箮Jq���0�T�W�N�Yn�o�=u=��V�{��e�ۯ��|��ƷMێ��7��Qq��^۾����Kk��nΐ�-�8S������F�Ld�ڽRԕ�2C�jG�uoI	MZ�t�%��.}]PikeՄ�ECuc|����D�].�a�����n�i5y�D;��Z�����Ue�w�9� g��p�*��HS�������V�톴��4��V�ؠ������zk^;kZֱ�ݻx���Ǐ<�_��)�Ѩ t�1���UՓ��]<x�mkZƵ�k�۷�N�<x��Kdym�յK��F�& ӥ/�zB�*��5�Zֱ�kZƻv�������~|��AAE�IH��E'mIA��h47�u%qǍvֵ�kZֱ�ݻx��~�_����Ί����|�����^6MI���Tv�R�V����6��H�V�dѢ��lz�����kZ6�j�Ť�l��uTI2Ľ<T�a����׹�֩Jh`�ӭ��8�IF��n����nv�V���L�`ՠ�ւ�1����~GTuI���'4MZ�h�ִRmNm��Q��������Z�F���V=T*��ZNq2(m�m�Ν1H��WfؒZ�;S��E7�9�Gns�;j��I�ͺ9\�3��`=w*�2f�?�>��:t���:T�S��k�����w����k�y�I�ax6�|��<���6&+�!"��喐m�bb�!%���G*�����M<s�;��1@&�d�h�:'�`�}xQ��l���m�pήA�PX��IMc�u�xM2{n`��;^\+��I���?����������Syַ=<ז��\���$����H�U��a��}~�F$VA�X׹a<��`�>Lsg����ݝ�T�I@��q�h���G��b׈���!>�@�P�s	���w������	��ќ���i����"ZZL�w���v@�����|�f�d��諦�)vl �'�Jo�W0��ڞ����/���8���(�.����PϚ-�G��`�X׹1-�}0��~�w' g?S�ܳ�#5|��{�>z�8�5�>'�0h]�v����D-?��{t^�����0���F��5}��eaӕ�JZ㽼eo�^vJu�r��<HMD$k���.uA}V�+�.�}ѣ���s8�I�2��O&%f�\��1���o%�}T�u����d8���}Ȏbݣ%(����>�D�rg�T1RF&���D�!�ՑGwK�uge.t:�^��3Jj�z�Dxۑ.\���6��)�ުd֛>�CfKO���P}�z�S��Ɖ�y�%�Z���gnR�f��L�}�f�m�v�R�St�ҥJ��N� �E�v�v�K��v��k3-��+���%�" vRT���Y2i�� �1��ס�>�㥜(gd)�y�:�p����{1U�a��|��|_�W�sXٛ�����DG�L �wu�7�i���*񆗆�H|1����_:ݿO��τHݔ��@��U�N�J���2�
�l�^��h�f��D�"�y�K�l��Wx����^1��y�1ܧ���n��jL�Å���3�%>�a�P��[Ү�I74yWB�ꩳ}Ǆ@���ɾL{q^5d�w�T�U�[���30�z��^�Ǐ�}��Z>}����x�k�n��Jq�9��c����;�p�k�,n�Əc���}�,m��M  ��<ckڇ<7�֣�X3�p���>쉹�8mI����]��C%���Tu�חz�S���y�����CGXra��N������5��sм�zp�H��'I�`$B�C�hj���[`�`1�\��p�8 �Z��9�y1��|{��������>p�Mx�Cc�p�|�&��0y��<��xS�����᛫"��G��o^��P��+�QD-/�j�Y�?sѩ{{g���w=+]�Y��ȥdn���EY>����5@�6vTn1�ꓭ����n�Ko�ҥhoÝ�eX9��
u�V���_u�A�c��K���ǜ8	ԉ�(�&�MHl�,�i�JjF��d�VW�T�R���G���L1�U5�&����{=�?'�zǏ�����y�А<L��K�W�A�P鳌T�=�s�̙��c�J,8|/�Au���!2\����xa��zw�>��k;�ѝ]�s*��=T{m�쎷��p��D =��#�=[�&��gK�VA/�,;=�Z���r����G7L��Çʀ�a �9��+�<q>:�{�{�'����ٌ���������z�Y��{���{��^RY�rH��D~#���8������/y	~�-��_�q���'I�C@c^����0���,�ˌ���"r���!����]�?D{+�kB�L�l*Q�܄��X���>�q]�lh?uXO,"����?M��ɚ����}�DyP2ߒ��;�$��{H�<�`���e�]�|���yz��\�Y-E���l��i�i �=}P�b��Q*�ʝ X�A�ߝmZ�_}K�c[\P��D� �FR�90�˞ǹq"�SAP,f��;�X�]�~��Ƌ�KƝ2�����[�"-{�ݲ/H�ޕNV�1�vN�<i64"�ł��F���"�)�=�pS�'SϺV�WY�k��o���X�>-w-˥�<�)�a՚����@��G��Vb�vXx�w	]�7�=��ھ�i8�8�I�u�չ�⺛=���F�xaS�l��s�<�|*����O�%��E�+�qi�����xg�^�i�[x@v�-���Z. #]>�{k!��v�4�D%�vX�.u�	ҙTv0-�p'�ro5휿+�����t>,O��yc�&ʕb�P�˟���Ke�_h�7��xm�䢛�=�_�=VFWv�ny^ X���7�M-��p������������M�� ?8��Ϲ�:aH�JO�
߮yP4,t��0��ãэ�D�h�8T�F4p��Bn��5$��0��I���H]�P���h;�&�MV�цv2#D��>��7��D	¡%�@���Q`�`���˨�W�Q��ҳ�Ns�+����M�[�@���Az7+_�ݙu֓{^�]z� O_M�?Y
��"�/���-�Bc���ϐXX��椠��}Z�V�s�����=���q酰`ێ8��+�B]����[ߨ�2�"=�3s�+,����Ň��b�Cu�q,��nF����R�8?'v�����~}�.��v���%���ճ����ӯ^���$�+�WV�v�i1�+�(m-b�����lC>x�y����)�0�[2�L�F��	m�jH�A$Wcx�n>���^t}�L�ʅN��j�ڗΖh.�N�w�����B��u�v�W���=츁�F��R�J��t� �Ra�S���~��Q����g��7EzA�׳�t�v�G	.1��#A�G^w���}��^/_��8}x�k���l^IV���z��=8f��1�?,{�'
QW۪dp��2-�C�/�z�Y/����Z�$��8C5KW�n='9wo{������?i�,�@�L�+��@���2��ނ��g<쏭np�O��lG��yR[d���wam���qE�TnS�h�K�,/yGi��lu���J��*d��Qݵ�Q2d�x��:�F�g���\����^ZI�/�@��}�V���<��$vU��^�޼v"�s˱��:40�q�q�3L�R�N
�o���{��<����,:�{~��̽���n�ҩ�`�ь��w��q,.��?wD��r�kg-ꁀ�T?Q�5HYy�%]U8��R8e�����!�S�/6&��.��2+��D�oQ���\�8<^U^QT���:�Ą&=��>1��r�n[�y�|���^G3XF�,$��VV��vf��7��i��ql5�q9VW�ݫ��b��4Q1��]Tr8��Ao!@�>y�)��Q���z�W�}�s֪�Yè5/zI��D����}y۰J�i�vΩ�Uv`\�
��%v�^�J�*T�R�_��9�]�4ȣO�~@�a:�ϡ��� yp,�Cژ��g �0ܯغm��Rʝ��آ�&��^�Ӹ���5��{�'�q������� �/X�+��ֈ���Y�A��ܑ�4(P�*i��y��\�3Uae{�u���`7^p����jeI���F���M��T�sy�p�{@IM(��d������;^�^�!�!!5���!��b2n�?WH'�r(��WvI|�J���W�ͪ2Bq��͍�0��B��L��E��y:�|=�yR)qF7C�����yq=���3ۇy^i�MOp��3�?��s�-��ā��u���>n�Oeix��;}�܄H�ɠ���F@�
S��?*�{*�]+�6�������X� N�za��W�蠥�`����ps��������W�J��ya3L�]_z/׽ƣsT�͞�͏ո5�?~!*3�Z��CR�u>P�w�:0�nX���sYF.y֫R�-�MCU4�w#�r���S
+���cui|�F��h�z����4
acV�_U��*��uuf�\�Idt�����pD7���G{�^6f����!�/����ج�v^s��h�6��H4j�l$K����!h�L!BAM(����Z}�^�J�~t��t��f����Z�V�5��ԜB�F�&P_i������~�y��c�p�ڽJĥ{��{����ʗ�g4NVr0��
�|�)ʩBj=���G O�WR���K��Kp�0���jf��*�|��V
�h����:���=�Q��]��$��E-��O{HQ.4և`��5��X��u�G��X�\3��
��r���stc3Sot��l�l�8�G������P~ʉ�g����w�:�W��=G�k��O��Z���,l�6���3�O3� �U���i��^�w�UH�`Vt���Y�;��B���4�#ɽ�o��RZM�������0ͽ�އ���.>�ܑ3��O峄Ļ��e�e�i�-Y��}5��Jh��u��ڿ?��ho�[��o��l�y���9ɋ��e�j��q\U�wٲ4h���f�O�jధ��|=��n�_Ml�#�ziI7o���=��ъ���:ݺg_;�{2׳0�&�]�;pCխH�E$����G��e�⇫�Y7}N��'T�U$�4˻�iQ�}���1��Z<y��:�Ij�lv��eJ�J�*n�:T�Sg7�Ϸ�eﳻ�>���o���#�|c��|�*/v*���|j���5�O��G��sxoO��<���!�����A�;��Jj>*�n,��9��U=V�V�n�RUd���"�
g�g�W�%0v�+)��LN�&T��)��Y�;u̹d�4n��w}ye�k�d������v���x�v7�>���[�0������ݞ��+��N��ݹ0�՜݃%�K��� �Y_#P{]~ab����Ky��~*�\������f�|���_W�s��?=���>r���W>�8�G8��9�w>� iI�,���{�\t�ƣ��K�9�7OӠ0p����A�.��}�8z�ґjL �PҊ��=Z=�ܫ�wgO����	���uY�f�H���'�D�H�,9T]v��� �O��Ӓ��}��f^�����{�_h�We����k���;+��hs�Lus81��7m�G� ��Y6�,�{�V��E9՝��-�a�6�`�v�pN���{�k��U+}&M��ckw���J2��ӌ�����ʕ*T�St���|�w����f�w�?���+�7E{�	o��{c8�%n״4ؗxM��'+�ܾ��=���Oiw��Dt=�;��-���#��s�j����7+i�����^q\pY�>�Ɵ.�FPtƦ80ܜ7��ۥ=C�;et�[�G��(f�� #��9"1��~�N�͝�ڈA��:��߷��|�t'p����n���ޫ<���U�Ÿhj��l[���fW�Ђ��=k�aVP�>��=����j��MLC*�C��{�ȵ�F�L'�����f���nY�g��O]�%{c{�ո����A)��|�ܫ��?�*{"oD����=����������{;���&Y^�_�±ʃ�5��_j�*�3��fɪ�1x����Q��aђ6�I'9�Q+�ӡ�����OU��OK[؎8��k�"Y�6�ѡgN��hPHrj���=��V����a��������Zc�+��U�}0��ݤ=Y��(�H�ީ�O;H�ܝ�UuY9I�{�Qa�h<:��*�ݒL�����C6o�oAx���ev�%�<}��8�9'rs������3�}G���4�n#��}&C<7�v{�&|�[zt�<�v����Ooڳ��x�;��F�G���秺��]�:*6-�)�ݲ�^�{S2͊0�D���ЋM�bD��������yz���+�4�x����,]�vu�15��Ǯ�X�2�s
���I�^Fx�b�/0=�H��D�{���|nzH�H\�#a�@�5�PC�kX�`�j��Z��8Ә{��F��8-ڟvq��|���]��������썵��2������=�U��?��K�����ҫͪ�r��,��zE�2owY�$@����$������o �����љ��)"Shp�b2�~���3\�w�un��mu���j������Cz5�j,��a�Pa��~��{^��6.yn9�	Apⅳr3����l �kA��b��'�M�I�r����!��ˊ*�n1"JȜ,�yG��ص��)�/WSdfj�/��ˬ���:uX��彷�K�N\}|�ob:Ҏ���'���m���޴:Jd:�� 7��#&���vͿ�#`�GC���*�f>ɣ)�"�#XT�v��HCC���27^wc�\��V
t���%���L�*���4j�P��;� �v�ݴ�	��j͏~Ƕ�X� ���>2�+JX�w�z�p{E1n��ԥ������s�w����L��u��q����ݢ�G2�XA�oJ�Ǣ�۸~�0]�V��>Ւ�w�᝸P�A�1}��.Dz�&>n��1}�W+*,:ɪ�֜�Bi.c����ih�7�Y��+�h^�{*4����;Ʋ�8���+��&�3�f���O=��(�Pe&�{Y���u�q,�f����ۅ\�Z�O��9[M�}Y���Tt����G�=Ӂ����MdI
ݑ�oFm�i}uC��7b��B���X��m���҃���R�i�J���%��d�Z+`$��}���ݼ���0�ЅkjK�z�	/]�:&T�5� e5�V�M_`�����j��H�X����p!3�W�u5t����3*�a֘4\+�cq	��)]BЃ�"�xE�������-4gJƶ>g��S�m�DP�)�����vb/F�񓌛�$�Zĥ�C+mW'���gmV�B)�m�A6�,�$v
�X���bN��[��S��|�z�'���ygL�#��p�1y�v�4�L�L�Ӊ�rq��v�z+eҼޝ�M�so�$�⬎��]�N�5�ũx;�;Mm#EL\��wWm���s��s��C+�a�+M�uE��%GhvE�i��%�4#�]�Nen�P�J�uՍ�X8���m���_Q'3 ���:�o\�պ�U�Z�b�W�Q�Nw,j�T��K�L�1ͺ�\���Pp��gyC�0�"�̡ת���a"�X���a������eFy᛬<#\��VR���@D���}��v9��êV9�����Cl5�����zU��1�0�����ȃ���Q��9Rb�E��u���V�E[p{H�Z�q-�SX���H9�7���2b������dU�n!λݥςahZ�*��o-�4�}*_s�g>Ĳ���p�;Y�x��G	���n��d�]��rC(U7���BU��A��z�r˷gmvV,�8��r���{2��S3j���Y^����xHCz@Ѧ	Y���`�h"��ݎw.�ݼMg����vf��ݽ��r��X�M�R��E�h�A4�rջI,*L��e҆��'-٨��!m1��BX�q2&;��I7h�TQ�"K$�m�f]�bm��
(P�!)#��*H()@I`����@]I� j3V܂/�{	Hi�(�B�i��@��2�(�E|��}Q�K[:e)W��;#�b�������iP�
�F"	
M*�l뮢�g]:t�����cZֵ�ݻv��zx���I�]Kg/V[ie� �j""���l�m%:t~΃�U[i��f�x��^�ֵָ�k�nݻx�����?>��F�N�%�ݵ�P��i�N�����٠��L�~�������uƵ�k]�v��ǧ�7�j���ESMD�D����|��&�*�]��(�ѥ���ն���Mk\kZֵ۷nݾ�߯����4��f�b�Ӧ���b���:
h
B(���!��j�-�b���AZtPh-�Ѣ�RS���;G���UF�(��6��^����E�c��y& ���Κ���"�&b��cg4Q5S0Vآ(ђ��5OY�F
)bJ"����UDkF�O��D�1L�1{��MQZ�X�,DE��i�"���EL��MTFƊ��"(�����e�י����>j�z��mᝮ�uҴ�u\�f��ճI]`�Y��"��w�;�Tz���n��=��ޭGA���鴑	@����,���������*T�T���ӧyu�WzW��o��U��`�ë5_��,�z�2�? 4gO�^Q���4 P�4�]���m����y�4c�/�e�{)�9�8y�Zf�{�LM?�wDnMu[�����;��gI�zEf���!-��w�"|a�X�C�=��Lb䌩��wۧ0�W:�����'P��p���9����깚�d����I���z�(��R6��w�/K�Y����]��T$ߊ�s24O5��uM͵�f|*�w5:T�@�C� ���L0V8��qE)ݯJV�t�5tG/�Ei�ٹ�^|�2��`��p�b�$@��)ϯ�^�=�,&��6-��L���gRebCgo�T�q��\�Ct�6������t���!�
2��w'��+JM�������9D����c0k���B9�Ga ��C�����Y��/��l�绛��{�oB���L����\-O���x�
�����4U��xe�-���|�r���X���z�kї}G;�N�-��q���W]�>�+	�=�����88Z�9��F�����cYշt�X��ww3AS:��X{��:]����Sc�[�����=�:����*T�������q�+�Mr;�7�>��s>�;��Rw�|��oD{�sV F�,�o/d����+q[s%�p�៥�+�[���ws��"k��=l��Ģ��@Y�V�ں^������yW�u�7ΐ���w�A��	^�x��I�U۹�S},�2��0�K�Aނ�~m���Z��񭁙��?H��c+nf��گwgT:��7�>��C��-�f�ÀpAP�7�gC�뿴�V��d%h�>��9� �YA�CZ��+�]���'��k�~'3�l����-XM��$J�T�����z�=��s�gKy	 �ڣ�4��&w/��wK�դi��`5��i���.=���E��2��q�tΣa�����H�r��e��Q�x�	q@�>�uG�z� �F����H� �~����g+�ü�������sr���_)��β���3��Q9��Ӷ`��]GH47�H�o�=M�?A�O3�0����yt�3e����~�[3��1�4�[.f
;U�Wv�ކU��3B�_h��vb��uv���}�== �Jv�z�bi�sk+�*T���ӥJ�67���~�}D7�����o}�=�W��b@�q �sY^�@3�I�-���>�#7˛ϻ����'<Opu����g
�c���#��M��H�F����8��'`Vs�j��3�S]���2e�C�c���<z׈�m�/��W=���@�O�{\v��~�,~2B��7Ҝ����w�D�������ܯ>�_�7�t��v��ۼc|s�E��cس�(��d�Տ�f���ϖ�o�
w�r"6� s%u���1s�{�zd�Y���O&��{7��CK���{h_K�t�zW��g���b[��J�U)k+����>C���/{,hVg�7
�p&�1B��V��|��9>'`0d3۷H�E:yY���~�៩Tj���6��\�uT�HPb���+$�v=c0α��3{��L�i����'�Q��H_��&Ħnx�9�_x֣9rLYюV�-f��i�p��)'v�;i�;%[�EE�q+�#!��PᲷxծew.B�k���}�A4���j6f����o����������*T����<�~��f#+\�4j�P���<�=�\��Q���8�b���td'��I#��!EI��뎡�����}\�ze��Nr���R���Z��:x��A�U�����݋;1튍��x��F���n�e��g�E���d0���Ӊ�uv,�*���z��17�d�$���e{�/9^m�`ݓ��3��74#�$���9�z��;r|Nx����U(�ώۿ����ʡ\���fZ��ȹ�)�8g�E�q4�nt�wr��\mǺ���i���M��J_a�.x�#ޟB9�Fƿq�a����z���
5�/o�sM��
����FZ=>˞ol��9z'��[�*����p�k�tl��`/>ó�A�|F�~�cC8������}�dԵAm�]�>�%�'�;�=�#W���Z�5�H�Q��8�-45�O*N����9�"��32������&s�b���r*��A�;��+k��":�RU�9D����Z�4iB�%�f˩BZO-<��&X�*0���ڋ�v>y�{���;��� =�7��G�RA�l̺�e���ʚ�	6�t"�LR[���ʦ`H����@��J�*T�R�J����d���=���n�+8ƻVbdˊЀ������/>������z}=��=���o+È�<�UWU��F_�#o�o
�:*7\G&hI�]�}S�',�oI)����'so�7�@0���";��rU����&�@l�b/��.��I�����q��כ�s��9��'�g�.OP�,9l9���S��=����t��٬��5w��Fˇ�v�H����ux>�`�|�|K�Y}Om'�7V�U�6�k2�� �4��R1�� ��'�Erʫ���b�'f�dow���mQ�c;[�/փ��Y�9��%[�>��bcέd�"8�fm[`��˞
�ҋ���E��{�wac��ٍCR8Ipy4�J�TDK;qqM�ݷޱ�F��)�����z�	u}�9�x�Eh�+۳��>���㦩��C::*."'}~�[��<�Yˌ�0�˚�
ޭegq@G�K0�6�Lq��}�jm��/w�=6$�c�'E��J��y�pM_�ᴫޅwl����Lp7��u9�s�Y7��|#7\�f�&28��m����[R��s��˻�%J5�T�R�J�*U��Χ߾���y��٧��L`�E��r#��!��~f��DV��+4�x�����F{�!���P�q�m���խm��i����Yg�	����j�ݪ5�oe0ら�����f�yq��V#�z=G�MwWq+S�����iPޫ�2j]oj0ԘNwk6��K�EϥV�Z!e``��c��4��Q�������ؽ�:�^x.�G�w)����� nwrD�����߷���Aل���@�=��������l�m�c�g>�*�l�0=������U'z}}�s�֙Q�ۜ�1a͛5~�S���A�pLc-qm����������Kf��o�(��-��jI}�n�gM>3 ��9Wp�c.�T�v9דgL�w��i��w�^(88&<1��lkp��͞�s߆ޛ��z�
�nL�D8�ub9��ivlG(�v��9ͫ���9�XxG��î6�[5:B��h(ZF�)���V~
F:�n�sE���v/�������� ���si�;�zv��-�+_E�
�ä�I�ww^����{�t�ҥJ�*T����>�� ����_o �����)X�uc:e������۬{:���sǫeLQ⛢���0f@ �j��r����r^�ZDd���EX��X���G���������)�n�W~�ggz���<�:��n"/�]r��N���-�*O,���$�mR�][��a�W\G����AK�k7Gwk�lg$�fLgfgh�w�P�WR w!� 	�욽��g�Gr���-�����Z�J+�ԍ�ǖ�}����ނ��ûό�{��tpyM���cnеnxxF����{؇���DH��[q;q�*����Z�z�7vm�"y⁇ȹ����=ES�#ޭ`�����g�t
��e���v���E��(�a�w����~-�lU�K�߆rO~��+����rxóG
�<���6�P�[�U��[�{i��u|ou���~�#�FW�X�\�2�K^k@��}�9�%��Ƈp��8^��G�c����_ct���O/���]��+��jը~6�w�i���^o�*!��q��[�;w�*��S�X�w��eUI����_�=M��-�
"pXf���?������=�MbMѽط<�Z+uJ��F�U�]��U�#KС'̷�n����iu��(��N�Iv��:�23�W˧�ůˢF�o��_;��9���G0��|��1~��p_%6��:L���[Y�z�� ��t����ٔ#�d'��땻���I�� ���Cs4�ҫt��#�e�6�w�K��v{ ��U��:ޯD�-���;$,6� �h��]:|��7}��O�006 !Ϗw�_�Ϧ^zR��|H��N�3zv�S6�+d䈬�~�k2^2���w���R�>m�e$��.��7U��4������G#�W��Sí8vz�C���+�#LL�bTV�=��yWFqݛ�1'M��'"�j�}��[�W9-�۽�؉^�9�L�+k�V�z_!*=ܻ�z�z:�luD3b�&♀��x۠b����Ξ�fl$�=옌i��6o��9>�)���>ѧC��B���K'stՕ�Y�A���J�����4��`�%}/.��%��
V"�X.]�+�d�ֳ��wv��z!�v�+���9�Z��c[�)cd��)lF�P3n�h�AAI��ffA�8e�JP�������T�R�J�*T��&����v�~��/��Ci��.6�K-w����a?�mt'��Mo7v�l<nc��Q��5a�;�p�{����d]�m�Ю
�vg�@�@�ؽ��#s��$���#yGgIްˣ��O��O���W��|���XV�^y�Ɣr}3��0�Nwi�&Gjx�v|���p� �u����l�M�ތyQ_�s�1uyyf�J��dF��3�y��1�[;:�!���y>��̈��������s���(�nx��X��l����y�(꬘�>a^мK-f�Z�n=%EO0�k욲��nS��bB};���M���X��:<V�e0������zh�7�_�	�/
�N^����"[D��._t����8��ݤp8/h<.�=B*�u��Ǭ�p�U�T���^����I�O��L�2�p�!�]^��v�-0��&������Q��zx�Q�_D���zk�@O�d�{5.�3Tf�Q����GYs�I�
o������ �MѡD��� W��s�m�Wr�$ch��^�"�,흺��ۦ���z���ݮ�Ǖ�NcqS����+��@u�T�R�J�*T��w��ϽΑ���ܟU:[�+j�$%�+)H�o~���22��<�Sǹ�<�P� �؅�I����f}!�D�$�c� �<�AvɫW������4S��|�_=W�6�'^^�3o���i����Z*��D��Wl���:���Ҏ^B}5`8oTI�=v�yӰ���oD��6B� O�%M��5���2�ܥ�/FԒ�2+���=rѺZ��m�Ԍ�rY������kp��{�s�	����k&aaa=�K#�5H;=~�q��yZ��1��(�]��v��ۼŪ�r������U����A�(����t�ׅ�������3q0�(<wV˳݆z��^�����b;�j�\fF�ԳW0�����l_C�s��{7������|���O{���]��9��{�q��� f2�e���i�^�S�`=�YO�ʤB]s9�'v��[�2E��e�Ѕ��5V�sPuv�|K���%�V/,��N̏����������z�՘�9/����R���؝�|�uo'ϰ�����M��>�cUY�MJ-����\��'��"V�m�7��5Ց^'V&4�>g���'�)vS�{XmJ
��&%J��U�dY�L����s��(���A�LJŋ���*!3��P����ݭ��ON�ɡ��z���w8h��>$�X�
��9��ք��v#YX�ޗ�,��
1sw���E;PRË6�)m�Q�:�a�U�C�����j��)N�&�7�<FmH�\壸�49n���M� ��B�j]�y�g'���8�f���Z�A�s浩���R�%���s�pÑ���=�/@�r��rWw�`�A�C{�,��9s2��&VuZۥ� c���� ��#��]6�����"hD�9Z�{���ԯx-�=\�ei�zGom(i^�M�+�y�G1WW9tL9�F/FP��eo �s+�&�����6T[֕�����]v�{�L�:�m���N�x����ĺ�-R�
���nC4���vg�r^Y�RD��ڬ�LW��r�s���v�oxfb*��U�{��q�����b�E��L�(N"�w/O����?5���FR�D��t�`%*`��d�[���K�����*�
�z��ۏ)�_P-�E��&�]��e�iq��>n�Ê*��'bŻ[Z�q���no=��Ki�PE�r���o�I�8m�+j���;ײ�67�-ʻ,��X�[m�<;:�wi����j��E��ζՍ�1V��^��3a��,��r�qX����&�Wwǔ�;xu�L�ʻ�\����+��@�˳q�]�i��e��c����ڣ��ī��[�L �r��7�uL����t�u�k�+띧�]��Q�%N�چ����|�4O�Y�k�v3]fo\��"I����*�&�����C �qgo&':�+3���<�|OT�p!�y�bӸ�q��S�k��){çj鹔�����F,�����%�qf���u*�7�����V����ދ��Y�c���a��MB�S�o[�:�
pUˊ�I���$t����ުU������O�D�WMzozԆp���P�PǦϋ��3`s�P�B�n�s���6M��&�+�r�ly:�_&�W���x��=êu�T\��;+�����k���w5�}�9K1s���ûdFa8I$6��T�����W�2z�]lI$�:mlCU�tTU4QI������o�����y�kZ�nݻv��Ǐ<���R(�)����LSEm����փ��X'<�~�_���ֵ�v�۷n�<x�,������Ū�QS�N��<��N:�5t:�3�|~�_����Zֵ�ݻv��Ǐ<�V(ѪX����wSE$J�|못��Z��Xǎޚ�ֺkZֵ۷nݻx����|�yg-�����QQPth���PT�SU�*	���"��>㨊��d�

b ����}Z�
����n�y�|�r��ǛQ��3�i"*"�$��K��M�
*<����(�"b?6"$���b
g��y�m�w%%�CMI2v˅-5TET_��
��d��[����":��5GZ�L�PS0QCQ$QQTRMQ�I��4H�i HF��73���^�y�����P����خ��%ɘ��!�o7�jmK��i������	���go�����WԩR�J�:um���:��V�_�~��h�����p�L�6}B��n����^g\Ff��2չ�F�Gy�S�:�(+���ans��Va�9t���F{�j�̦�� m���ɉ��f�mi��X&,�V͔���Į{�;l]KHgu������S�c�I�^��[����%Ĳ���~a?�UxȄUz��M݉E�ۋ:�0��^݁���\����Y�%
�x0�Cz���40�7H�|��3��s9*wZ��bL�+�Ƽ���Co�U�lriy�J��f7'k���ɫ��)����՞��������u PopUs`2/Kvb�F�'ި�El��mG����r����b��{o �|Ǭ���ʱ6:s�}�w��
/*4x���<���v|�����Iu���n��β])~Ɏ�ֹ�/M��͋ʂi��Xx���T��^]*yx����i�6��+7�"��<���f;�xJ�����]�v;�gb��P���{��aO7�W��h�l�tt�Y�s�y�Ck��ӧJ�*T�����Y��[=�@�ߨ��ӻ@w�*㣷�P0gqֽ�Е�yuzkaQ�wg�)�O��6��y�HLY�!��9�3����a�������$�T6/��H9�T}����-}����]p����� ��S�e�,����9a;����v;b�>:��1o��7�$��<�4v\k���7
zU���q�g%3]@?�����<�m��@ep����j
�u�ꡏ���Z:��<���he�a�_uzd%�g=chlxlz���`�m��^��fݢy���9�n+��>�m�/t�Aa^ӧ	�oi����܌Ӭu�0d���.�h�wt��Ԛ�FI����Q7-w��֌H�p���U�>���N��L߼v�M��ڞ����|M�rR�{;�-������S�
����G?�ﺄ��vL���5��z��A��*�Mn��)�V�Th��I͵c`�,��U���R nm8��SD��ճ]��nil�G!�ʺ��
h�	��s�r���I���WQ}Us�w_P���DJЩ��g���n���J;��'��1�oL�z���)��eHgZ���A�p��N�Ww.�(��*]*�*T�R�J�*��a���~��q����"�B\���M�9_������RU�|5��L�d��.(ro0�jkME�3݈���u�]
�@ި;`��u�Ko��cC�WR�|jݛ��3��}*������z��K�� r>�R_���z��[�ue���J$�i�P��v�a���C&�^UWu͇�r�t�ǻ���(;��Z���Tb|��mә�@��.�r#7�ջ�3��uLK����o7�<��v���4�y��^�|n���PFs ޸Ƃ�kgy����� ��r�[.�	n. 0hom#\��5Tx��l�$y����L�>�@�_���R����;��P�O	�������ɕ�n�jO;���������D�cc	������J`�1����Q�{U���]Vl7V5�WDFHh�K;��K�`�aڦ3��߹�X��T&�Nף���C�2Q�(#���V�l���D���l��l�t?c�]��E�ѝ�F?��m�\����_+O�ge�d�.�M�yZs������.�L(&r4lN�x���I��n��=���[�Î�>�?�������?��u9\�t�w«����W��[-�����]٭pMN�	I��3t�Ļ�����7Xnl��w�6��4s�~�Q����{����{ŵ��l�ԗ�#��)<��;o��u�1��C���M������m��7u�P�z�|� N��jɬzv��?��xx����L�vjjj���z�}�w�����ùX�oM�PjH�T�oM���O��?]$U>2!_�(=T��_����Lb�{����jQݻZ�p�_��'NR�1E"�+얻|q���0{�%��}f��Th�:Ք$qP�3�L�%F�J/v@�G
����3uy��\�N@r:ÿ��ro��\��Aԗ(I�O�ٴ�XG�e�췯s�CU���Y�^�^������{�@ޟ���3�$�!�{����R�3��K-i��Y1���5�wss\Ԝ�Z��e���yV�+��)���z���C���)
D�	А�`�+)@�LA~�����׹��i�qie�{���A]����8-�;��Ρ]����w�W�Ӝ�|��*�v�J�*�:t�R��}~�}���K�g�'v:yH;]��Wv�������^�o7۵h�{y��CTy9x��O��?���-���^J����������*�-+���!)��*a�ul�>zg�w.'�ٕ��\�g���ՅR���-#�����1�,�l�sa��� Aη�|'�n��.��4Ld	�s��y�Ϥ�R�-6���p�o�7h��P���zs�tC�P��]�g,ٵˁ��ωR1�N���@�o��t9,���d�ݵG<�1XN�٤ j�^���7�P�n�?�<
��1xC��졊�Č�}GQșFJ����X1��>a��(�g��ٌv�'��TU=��/Ś���,R�Rj��):���G���!��	�2ԘW&�^��g���)�!���8L�p虿w%J��Q1��γXX.-�v�˘+k�z� ���Wln�l_h��T7Xj(Z|0-���f����~�a 2�A")�}��Op�(t����W��"�i�J�U)�[�}�,��f;�@��;��!:1^-ެ2d�	~�U��*T�R�J�7�YI(��8>�=���=ylc�f�A�,���c��E�ڃ۱|��/�O2s�M.p��[�T!UY���%��n�%ųU^n
��⓾��bn�m��&�k�wz`�!���^��q|6 ܎�G�t��쫑��5�p:Z�t1ݰ�fM�9�dw)FDk�p��H�2�0��7�z{�G��a�˝5�(����0#e��9���(�����"��1�)����{�i�7�>5w�a�p��8p�ͽ.�x�Q�n�;�4o=V��mQ�k���ǟ|htJ���=�@a�F��;4.rm
�!��O�6i��'u��:Y�����%�5%���3�3��`\��i�<�/�y��&�Sz�=�H��)�]Nf{�A��0O�zѵtwF�Y�[�F�K����.�suf=� �]�'�j�XcK3�:��?;���"�{P��֝񙒯tžg�k�D7c���-_��y�<�m�Bi��T�vsw��5���K���Q(��`���� �
TR��X��7�"t�����枛0]��uh�{��p�c=�ӒG���
1��3��[��wV}�@�6j�T J��I��I�Bf�m&��"$]�e#Y^�J�*T�R�_�����O��c�#H&]�� 
�h�jE�\
W\��fkǲ��~�f���c�sw<��g�Zd��Y�����h���ц
�ѣv3jW���>�4tT2��U{��,J���{�[���B}�cϧ�<�+tQ�7���ڤ�hf�y׭oN��"�%ky�6����ozd!���]A�r���0���p��y�DFu�	h8j̲��p�3��j<)�7Ҹ�]FuN^tչ�� 獟J���r)zj S;�H4��C[K��⡁���|1�~a�����073�Ў2�I�SИ�ѷ�Tʫ�R�`���}�6�3?T�9EO�S�-��}�����T:=L�[�="V�N�8���$��&ߪ����v/�ps���{�!9�u��̇>nOT�8�X�Ŏn��ηU�S�H�oak^������ѤU�̓
g�.� ,�p&6�S�g%-(ӨV�h!�/8!C���A�5���z�ɉ�X��d��z������Å*+���ƃ���Y�����o���c�PfoL׹ۼ��iX���齮�8�U�.����{vY�O��x���?��G����'T�����6��'݄д�{+��z��Z��������m�w��d�^潄��Q����L��*M���ܔ�����9�+a��ȫ�;�5�g{��9^���z�^���u,'�u8Z:��crxw��ņ����Ӳ�jK����i�컞l�*�F�*J���ᆄ���훁x�7p��O�=t���ʟ�X0���;��%tWvG`����yY:Nm�u=�/�۳�ǖǔ�
;O�=�3�n��k�yP���-_sVu��T%���p]�0(�!d)��#����g�������ЇU�j�df�̇��+�T�O���}�	ɡ���po�$�_)����v�⵴���i|��>�{��r�V,ޔ$�Ee+y}���Wq����Q_X��#�Pp ��L��~��_���C7'x7�G����ľN�8�Y;*��:ei��u&"�s���uX{}������JD-�	�jpc�n�1:��w-���3����Xu�=�h�gv$k���_bWw0J��}���ڝyCl��s�{��U���g��x��� �R�J������{y˹�K�se]d5#�����-C��*�����}���1=^�mQ3�Oj7s�4�&����t���Be9��ƎWx�d�z�[�3�
���EK'xw�>�-c}�ؕ�zh[�,4TR��QK���  mz���<�3�ܔ�֊�W�l:���L�;^���J;�G�?�a� @=G�b��p9��6��j��ݫg��i���{{ږ�4����_$6��B0���9M2v��.&1�5�lI=�Ii�o�>����������
�{$_&��'���ಕ��2�g.΋�ơf�[����q����q�9��`�v��f���/�n�!*��w��_^S�������b`�a���S�n$h�sd�� =0J�*����׳�5��%��G�A�����b)-G��m]O��셬Χz����&��z�
EvX7.D��^�Ҩz��Ӝ���$���S��@�I<Q �� �^?t ��m�ӛq�޾�Ź�*-��r�����3f�c��ܮ>TS�,�Ի"4�kw���_��{�N�*T�R�=��{�{~��~Sƻ��I�1�nˠ���^W^IΌ�T���x$t�������B������ ��j���2���[����>�h}����s�I�K�����
( 	�C���=�����3���E˺"jMiE�ۊ�H��X���k�O�~��OE�)1[�����`!�����A���~��C��Q�Vj6����[�ގ�wo,Ⱥ�9�m3�l��>��f��6��55�x�ۭCl`�f���䍨����G2}SN�VH��9����H�Hi5��]��?��Lᛆἡd�K �W��:3ιݚ'�n���[��f�v7�_���t7�ZDID��ئfdO_J�K���3N��+����W'Xx�s��T�Ȑ��ٝ���+�_�wGvR(��vO9 x��ۅS�H�R��ͳc�?������(��N�(��5Dж������҇K﹤���@W�е��u�9Uй��l���`j�
�H��JX�v�a���ܑ�:���ͽ��Nڡ�3R=�T�,lU>�-���%����e)[WҡB���{>8���!b��Z��JM��٫���$��c{`��vbG4�O>��z��c��� �Vow'�K�y�nS<9ֹ��(��ʄ�D�]Q���GUݵ�&'�Qx�.�O7����gl�Z� ��x��.��E�v��#v��WBH(����V*ت���	���ESۑ����y�t�;�m��e�+{5�0�-�b#lgx�/ˬ�Ƌ�e-����b�Ⱥ�y�˖%�Q+W�t�oA��v4wd�����nF{8�\�Ǳ�i�I}5�6�cX�:p��SQ����[��bgi�d��fc�ЛH�PøQu�0*���F�)ׂ^�C4��J�+� _�;4�l�t�t��N��^c�͚|��(\*�����!�PWh�Cg���n�Z�ò�����(�_�i��68J��O���X��\ak�;/���R��8<D�����d},��-�Z!ZJF����ET�8SH9�\*�����/����[������Ot�޾��ڔ����T�l�wQX�f
�"�s5֙8��,���H ���h)m�U�3�
J���4�G��#�q�K3-C&<qEO���Q!P�L�5b��L@�K��Q��;�:m��B�,+��������$�O���n�D���lq\P�I�I

� ����mq(J�u�,NZT��v�����:W)�����SVy�t����8�M
 V]��� ��w�����1��,��4L�D��녽ڗH��]�U�{�w��"B��Y�ڔf�ۥ[�U�Vge�5jwF2����V�a��*�#H$Ig�Oe��Ff�Ô��x�ɋr���}���5�'��9yv�+wjYJSs��@�)3�^�b�+e򬵃m�ܢ�m��U�4��6%Q&�,)Q��u�J�r)*K5׼�X�Oo�BY�S$�u��1���Y��4i�Ip�	�W�{���S��Z��*X7v2��I�ܑn4�6�-aV+#[�TɄ6�EY�k��{b�Cm�<aHzו�@�|X���j$×Α��]eS;���q�-تq�Ę�w�>���Pt�:�w�OU����d���n�MWqS�Z���m�ۜc"��[ҹ�s���P��k���%��+�q�ɹ�<pZ��{����ƕ�x�޼e���8��h�CM��U���Mb\y��bDb��y�VN�p�ja���9�L|{L׳��;�%k�ΫO�www�j�	'h�w��h�e��,7}���H���$h6ᓊ��!���m@��	T���`DE �
	�I�fE�
E@�a�bf ٩
DTT�qBSN	"���b�����I&�\@���:"$P",�[bSV,2�Q7/�v�l6'���9��#J �H �]�;M}ڂ���
j�*�e�,��d�%q�v�׷�5�kZ�۷nݵ�x�KV�-��V>؟��(��T4=�E��j������MQm���<x�V��k]�v�����~�_�����"� ����4oyǘ�'�=8�*�*��U9Υ��eWx�����U�kZ�nݻv�<x��|�qzN��/DDPQ~�QEQtj��6ŷ������l�US9��������kZֵ۷nݻkǏ7�-��UES35k��ז"m�UQ40D��S��33����4�][T�E4�D�7�OmAV�=^s�����tГ4QTDG���Z�DKM5y�E���=:����)����D}���hh���z�]6��ATD�4�t�=#�H'N�6�gU�]�j����T3S��H�b��+�wX�������ETK{��.�k�[_�^n<�:�0i�!7 p����ꐎ�C:�r����M����6��#y�Z���]Ns�W����A�;$��e.��#*�%@�PTPEh�)$#�������;Y_R�J�*T�R�B��������!$`.��Ꮏ�ʽ�Ď���\�Wrb�0d��,��9�CK;F�E��;��!%� �tJ[��W���5�=s��8�0��c��6zc��<C��x5d�5�v���z��L܌�����Lj�R.{N���D�s��
@�Iw�mљ7��ޯ^k�*��2V��p�y�ͯ��2T�*�`Dsu������VҸ�'�Í�������0u��Ub�`̺i�es�ΰ'�Xm��A������5����єn�;������2	��������z=��9���\�]b�-A���iY%m�¼���CA���w��m�Ԡ����h�������57?v�VFe���.��;�Sz#:J���^ғL�e�/��Z;��v�������S�ݢ�ʘ� �S\)�T�����5��D����:,��OH�"��J�mk�k���+M�qgz���q�����f�w�z���W4�n��\
[���X�m�䄭|��͍3E�%�\��-���.�&�jvu�������y���xU
�]����L��.�hWB�[q�}��[��ǌ(�z!#��ٌIV�^�e\��p����2�=��S塪����}���?#��k�����y\g˻���m���q �=k���D�#���%I�'K�r����*c��kzT�#��p���^��~QP`�#����� M��-�Y�"���P+���xͨ�M��_$���d0���2��Q�]��+h��F�H�|�/��Y�{������[>�Mˎ�V������> ���,��߻�>0�<cgCU�X&8�d��Ƴ:{ʺC�ݙl���+sc%U3�y��Lp����u�S���w<9e��d^L\���1;ױ� �o=�	�T�`�SG
,w��o\�(Euhͷw�׺���f�㨧��J,��T*06��Gߨ����ot���Y�������T�a���K����U�,��Ɠ;��)pU� ��z�!Һ��E�>�C�9������g>Հo�f=����G_.�o&��;[�,��zPP�wEm��۵ooZȯO��7���xI���o\6����|��.���܂�D�r���z�N
�d^�dD����:���! �e,+,l�<RoKMZ���>��G�,�V4�ɞw�=��6��/v�J�/ b(F��a����H���I��+4=s�5;vEC�nb6I���7��z�	`=T��G��D�wTVo�x��a-��g���H?%I�U���*���p��t��XYЧ�ɘ���6�#*{X-g,S��� @;��`���EW����k�F,o]yۤ�:���������Z{��������')�9=>�n6��J�2fW-IN��[&;�9��	5�ݣ��ͳ��Ͷَ�� ���l����-��)�`L#�A�(����1��k��)qN᷺�:�X�[��
�RI������2gW\���;3�k���O���5p������zc�JE���j�n��ʭ�;������V�}or��{�v�Sh���4��,sN�Nx�ԝ��A[�놣]��6��%�fsSBʮ��/�Π\�w$�w����-���߾�่�-��0��bN���^oa��~,�n7b�Nd�/�s5�,'Nvc�v�xPO�}@n[������wl-�u)��w�]��[X�Zo��ov#�0�	
UE����<�V��&{�}�[S�L3���Г��>��m�#t�,�����������[� �d�3�챯�Yy-�Y��;%�}՗��"Dr9�F�7$��3�s��`{�3��y-���v���`
��vȱu-7gw��o�%���xř؋��!c˙́��qF<�=*��_�3�y�[����5zw'����������Xڏ��}|��bKn�p�.���:�K:@��_;�:��,^I�C�5���hX����(�;,��m��ĳWj�����t�^IL��^�un}U�m�&7gC��ݬǚF��ye���K�j����u,Zm	*��g�gBK�5;e�w�����Ѐ�AUD�  "(�)�(����\5
I#:�/J�(���)���]G)±�rnt�]���2�3�N�گ�dy2����ΰ���ٽNZ&��l���IH"NDԒWl��aeרѣF���X�����~c�!	��w��z�֪���܄�G��O*��ō�ݙ{e.����K�J[8�� a�ʧ4]0��{�@��������e�,8�[�����Q��P�u#XP��Gcy`�����µ粴��z2MZc9>��׉�i��+�����;,'Y�p:n�a����|�):�kr��+IŢO;Vz6��������7����dy۩��+"I�SG*��ܯ3�N�8�蔷e_@Rϖ��͸w��k���mf�����N�lDt=�H��!"zhu_����ק���HƎx�ݾ9���	F��oLez�Y�����5�+=T/��e�v��ol�6�#�����C0iʺ��w�0��ֽl���r���W�1������;�Т��opZ���!�[������hB�z�kK�|/VHy��3M��Ri���`��H;��Z�m�<tj5�G�yV�D#ּz\�+|Fa0��7�-.�����(lz������23x�w;b�-��v���8WWe.=f7b�����%)��Oi���>��v��33��w����y��;Ŝ&���R��ă�Sx���bދvpC��o��/]�u���;�����*�oeeL%D�O�~@��J��O�U����fm��g	"#�J�V`��J�: L������y��V ��P�;�}�.D�{y��~��TX��>��	��j�t��x�^��$�TS�W�_d�R=xnTĹ!����gfP�{|�R���Ԍ����19�><y��*�s��%l�ώ��޵�U��O��G�s�|w�C<$Vf�2��Un��ŶƝ�� L<��w�g���@b��ϵt�>�D�q���N�|*�T�ʽ��;�6�\�V��i�zBG�{�̵ن���{�E�3kVdOI�����!a���1\���Awv�;=>#x�LUm'�$���D�d0S�۔���"��������V��ʐ�ų��k�-ы/���AA������o��x�*y:���ϣɶ4-���e�� ���Y7{;����Yj�4�¢j���.���rc�����m�n���[�)���p��!s��b�h���@���o7����m��U$���y����q����Ǫ̬&!�����w��H���QǾ��ce��|�s�#l0��J9�w*�\���[�i�7Xl������鯼��G ����R��Z���d��S�B�s_��Ց�`̉�!9,+���ݚ�@Z�X`-���zza-��E2��_��|����)ik�����!��Ÿ�ێotr@H�E3��mCBgy�^N����FtH���<v4Q�����?�F;�7Cy!�@��U�nn��-[�y\�IM�r�!��:/��İ�dTr9`V)�oJ�����t��Xfs�&�W����צ���B�`��R��ʀ���M��"�&�lg�3�C[�@�w��-iF�TK����'�2�eJ�pҫ�}K{��b�����ɝꡦ��/B���<�Ȥ��w�i�M!����ؤ��_V:����~`�S$�[���� a�9Vd�<[E�6�q�M::�ʱ��c�[N]�ᬾ�w� �IYҾ_5.�SL�zbQ�T���md��R7�A�=����|�;�8��W �\����쏰;)r�F�4i���f�.=զj��3�{�����й?�T�T�];M>���^ߤ�&�VdέΣ#-�6 nzD���
}p��׃f���t�b�}�퓕�73���#r�����i4e�'���m�a���Ñ�<��R�H�]>FsM���n�l�)l���(�j՚hΡY{!�;K�9��#)ó2�P�W(��k[���>Q��ڤNI���-O���8�6�
~��w]"��m��E�!�m�d۾ZA2���\ݎI��^��0�o簳vC�̏�����z��C�ɽ<d�=5�����r�H��N�k^Vܶ0`�<��4���şe��9�A��O��bsރ=u���(�Q&=���F�0dzӬii�;yʛ��x�����j`r���FF��H$M�%F�-sSLs�4��F)��D�;@�	gT��|�_��SW�N����k���Z�ɻϳ{���mv��)4���ʫ��,^�;	)m)Q�H���WT�c7�����[�I�k�6����i!yK��a�a��vӘ �SA
	Pػv�X�G���Fu��c\�Gg[b�1���b�������b:��N�9	�m�vM�J��i�����m*��*�p�[2�$Qs��UVJ��S��9}��yη�ަ�V�`LH�+��/^�/i�6З�Q�]�蚓{Ǭ�������)m����,���f���+-H��[޽UbA0�p�~�-s���6l�U��l֯֏E�	�'�7k����f��l�6YЦ=�<�zv��[��`.����S��1��ka?��2�a�un�fa�O6Л~ڽ��3������'r	���;:zSKP�ׅ���J��K��M�����[�v�djx�/U&[4l�g�餓'������ˢC0ff`�8T�ͣ,���3�]2�u�&8��xq����U1>���vA6Bj�~��|S�e_���ॢ��b�"��1ۙB� �E����$��(A�����XU�����d�35z�����`Cy �b"�f8nF�vQa�� �������ؐn=�4���_BK�4��O��}��O��|��Ө�,m�3 ȻT
���=�S���U�v��)"^8���*��M�5�0!n��Nr#$.������u��f�a�E;(@�rC������t��l�h+�]����D����L4�sZ�}|����u�&��t�W����&+Dp��y��oB�[�C4z��z�b2S
�
�;��'���a7�0A-��$�eM�f�1�'͸���qدc@�*_�1�{�.�i*-C*q�Vf�,��k��z��9�{ ��hYO��uߞ�u�%��!��i�ةs]���a�.����h/<�����j;�k���dк��Z���D7�9����@�Q8�C3�"�@�g�kY�R]�z�+U�H�����)��nmFjf6���N!���8dt�_�H��_�b���tHgvw�Jj�/�bw��~u7Y�z
ď��n�k�uɑ,�1���v��B�P�i��m���#O�ۇ�ƺ��b�Z.c�ݪ��wxa�䷛GNP�������F��؉��Պ�D��{�DƁ�U8T�^��O�L�pN9�Lo�H�<�����[_s\�ȸ�,��4Y�o,��5[��&�0,�<�-����j�ݜKH��S���}��{�M�W���4�/I��d%Pj�20�q+���j<k��J�;z�*��֕��B�ΈL�*��6(m�l5t�%gm�rq��;93�n�;rKY4�V`֏]%��vj� �a����/��V�N�rd���B�vf�xk��#Uխsb�(�Ð�ѭ�!s���;��6��C��1���7�I܆��]5�T���sd����Fy���(<�"���VI��9�+Z���R�Pv��X|���E�&�J�:&^�è��f�,��Û�h���x]�#S�mfb׹C�e>أj`���}�eY�)����w���o���{�E����Q�c4�����0gAZȶԥ����5y.��q�z��{.�`�*G���m�w�»�i2P��8H�u�ڹ@����4d�k���o�jj�g�9�ۚ�݈yQ0mY�ţd���ï�H���=�|�ix��֠�cT������@(�xE�4Qb$�
�U
���l���o]1z2��s9D�Q7��H�;�������]_k����euFoCX�j�	NYS�6�U��=��y��%��oO'XҪ4��c��)۰�`�,�{��~�`���ӻ�-���H����j�b��P�c�<EЬ�w���O������Lakp���y�曾�-��Hn&�C����$1��ZY|��z6xP��]�[��2� �Hjb���V�P�4-��Vh$�SX}.垇\w(��}��j�M�/'
={ך<�����q��:z���k����G38u����X�SJ�=�w4�;�"�\��r��@U�D�Hy�z�-���jdcE݅یv�K�a����4A��������mpJ�r{�>�ʋg2"Tk$��m��05lӬ9s4�֡�6�@�.��9��w)�m
�\~Zzw	(�./�>�ݹuADF�}�	�[���l\9�զ+��6(ت��%Qgg3����Wo)��|�q
m��;9(^t��Uf�����;b��sLXօ&,�.�7�E ���J�FE���ќF�u�H�8�ܫ�e�y@B�Q�ԗ5w�蹉ŦG�R�=ب�tΫ�s�C��F�Rb����Qx']ޔ��X��������l��r[tu�2�Mϛ#.U���XׄgG
.�P���e�����b�<�Z���9�-;ܦ'��	��i]����1����1P��r���}署����.+�[K3$;n�	�Z9cFn4u�B��O7ES�=&Z����oY液�'�s�kGT��C%�H	������������=�é�̓���GE���43�KՁ�R�"jٗe�閫��b�2������fޝ|%΅h]eL���BR�n=k�/s��X|����w���P�u�ouvQf�]Q)�����6�d�)�.�����R�4޶T"�@��zk���
~�WZ
�k�����UT�kAC�N�H��ϧ�Ǎx��Zֵ�v�۷n��������qRLW�h&�8�,V�Hb�D?ˠ>ڣ�(��KV��J��Rt�o����65�kZ�۷nݵ���'�ߗ�l��,��T�q�(�a��h���T�-Q��؈��Q����*��S�q�}>�O���kZֻv�۷o���~�~�ϸ+����t_���MMT�"����d��Gd�T�I�,��Ԗ�+ݾ�O����kZ�nݻv�}<|�x�I�u]^����O��A�b��((���UE%���/^�8��cDEv���]&�����q9/v��͒��+͵�j)i���Q1�15�]Em�A�D�P�x�65TLEQ�C�EKGZ�ml�MS/l�!E�f*���{Ϟ��*(4�0k]W]�:�.�$Ku݂(�J֛�h�N`�?6`��b(���Lǘ���\�S�6(� ��(� ���h�	-@�ͽ;M;l*(:���e9�c�s1�;��-��ʖ|>l��"���jf򜳯8����{�]��}O�UUU7>o7}��Y���dx�1�QJx���O�n���ꈇg���y��f{b2�u�XH@�{��k��&�7������ҧŎ�x}�^���:윬;��o4_��suO����	W�ݱ�_$��̮BX1춗�\��N�X������tȮ�o{���	iկ��̋@lvw�b�Fv����A"G������S���Z�5 D.�[5�pm�k��~����pi19��H�f�mW0V��6zly��9�����7_fӺ��ɇ:�ox�z��b�:vo��������PF�XE3髼h�Ô��zZT]�of�
|��{R+B�06�fh����b��ŧz����mz{vp[İ� l�׉
�'r��|����ŏZ�cV�ESS �7�6`<"�IV�5�ӽBt���D�V���'�ӕK�o^����FA��W��^c��H6p�bt�d0�vfGq'��kU��D:��&�;��d���/sB�eܩ��w���\�6%<뾴]����v�b�ݽ`��E�&^ ��������������E��A��`̣�\�&)��<��+7�40�y����67y��߬ N��6z�6��d3������:�8��`kx�"�^$�;��xP�D����[��_���>z����q�}L96y�!�Y�11�;Xv�n���tD��Kg�	R&2�����l78���W݆�ٖ����4�{�u�.=�BUA��|H6;��=�u��7�ȈT���ε;�'�<gH�%����x�=ܑ�R�&�2�,F�i���{��p���!�8��wms;4��6;6j�d+m�ۥ�8�Oo�\����;K��d>&�>�\��x`�}S:�+	�5y�s�a�;^(�S����T���b�`����u�\�s=\)����[%S(���Gv�/`�?��gY��2�5��S�WS8��`};��u7���]�Y�F9�-��%��Y:����pms~�����!�wZ�i��.��f l�V�/ގ-����rU��](�Nn�`�nkh,�瓚Ck�w_f��OS��Ɨrm�[��Ic �{[i$ �-�i��ؼ0�D��B�r�F��5ݖ���Y��P�!�&"}��:;s�Y*�����&�:��{Kz�|F7w�kEcUݔY����>��87˧�qq���6|��J<�V��-m�y�w����OTy�s����yk>�|�ػ�rR�p��$vf$�-�M#�%
�gӬ�v���x�T"�H��\
������z�I�Γ���x׻�yo�ּ��k!�(�p��hy�]*���Mq�nj���/�71���RF�YJ}�O!y��1�;}��!�b�����ƣۥ]"�D�	���	vy|��:����玸���s��'|K�l�J�(q��*�L2�a$�eTE��}Μ���iR0M6�)�.(�j��?�L���=��;�y6���3(�֍�x�e�'Vn�P�e\�1��@�\�C�l�Bw��}�t��7td	�}��bL&�܌s��a�-��rw��8;ܰ1^���(rU:c��ÕҮ-�Y�t6�O\�-�G�`-{Q�s���O	��{�㫫kD�ŕ!�z�n�(uC�N�y���F�4EZ�yޕ>��;�z�gx���~�*��m��g
������q3%�{d�=8��/y�u�8,�1��O��ɻ2&ڐ8s�
���ݮ^�S�7�������^��gFH&�yq=�Zǹ�a$Zvk�{�>�~��T����.W�S=K�8I�Nz~k��������ވ<��
�y�����$�w��@ =�{�{̃�����4M�v�;�d����d�LA��Z������3�o,��2��׍{�Z$��o~����k�o��8�@7��?���
FFko��-�l@�z��zj�Pj�Y+�Rݢ��L�����y�B�>��`47Vϫ�T2vqa�U�P���<��H��l,�BG��^ʦ0��TH��<��FJ{S��Y���X�k'����]y�y�1���9=;Qt������ZhKs�4�T�"YO���hG0Y�����wQ�]k����e\9�[YT�;��B#�?/W��Š_�@�gKS0�N��K�6X�Pb{�2��r��7}uɡk�ޜz����Jx]w2AS�K�}������ª�
�(�L���p�MyS�隧	^zEb�ǜ^�{:Ѕ3�~�Na���*��+©�)g9�@�����r�=7#�tT3�2yn�y��N�#ĥ��^K)�CW��ԊZ|��ud�A��۶v��h�Dp1nJ&z]LXf�U=��ঢ়T�-1�+1U�oq*Nm�^��p�B8D�ǿ%�u��}������E賴W��������q���=�F�E���zQ�!���w�S�X:�*j�iRֈ�b���*��;�iL�g�����"�i��:�Z�\����.� u�h���Nׯ�'��&�v�p"Zf����]i9b��p k��mg}k�H�]��p^�':T\a�w�ٕ�N^��Ө�&iW@U����=ٳ���|�wN�g�a��3H2v{0߱���Ίײ���o���3f,k+K��.GxN��
m��izg�Vt�nz���ږکZ�L���2�-��n��nm�UE�kt��U�]+g>u����w�]�_ƍl��C١a$��������^�$���6׵6��KH��/���^���v ����G���|�g\��t��?�Xa�&����I��|����>4�4��'�o/�76����n�32�>dS�jq4%���gU�#���ך�ZQ����Ж�p%�S̷wqm�iS�9�E�s���p��}�2{|��VQUP�E-'	�
:�u��p2
^�>1}'ў����Gta|#�?l���Y��, �lP��vf��u�)��g�t;���lJ�~��Wj'��ԯ=SW����in��1�ޕG�ʺ�=ܮt��W�@jy|y-�;����2�ॲ��*E�T�2L��2{y]�����t�J���5��K
�ճ�	R��O�%@S�r�{�[�=��N����c޶���"'&9ǧ��n�6�`� XW(#�=O3ߵ#eS�C��䵣+ff7:S���{B9aXSuU���,K'�R��PqYe;�,�A5)��ߜ}ټ��e���'-Q��[��_2o7&�()�{ݔ�I�����e�ޜV��\�W�����!�� ��I�\2(��h�hѢ��'w��w����4��m)���3�3�S�s¹u:4�S�ެ��y���V��Z�mi|���}C��y�.�;�kIfX����l�Ϲ8�;�u.%j~އ!����G�3TV�ʹ�՜�U ���]�Ϳ\�W�;�@W�e��l�t6��J�Pز���ۥ��F&�Ƨ=�������޾J�Mv{��Ƴ�o�<In��7*a���Qō���� ���=��r��d��5��׵M���jQ�y�37
�`8s8�`�O�p�xW�X�*�n΅�勬��b���j�ޗ�n�������R��R,Y�j�tƪ��L�w켵���v�D�ѩR�Qg΁��**���0h�#1��X	��(�w�o0�m#��a+���Ӌ}��	Ud�y|�g7K��&g��֨�gv��X�`�M\����*it��������5g��̔��xx�i��C�L�t��n�]F�V�L�wRq�l�)�o�iE�! ���t&����8T�z�_I����}�o�w�f _�����y��*iV$�%z�K�D�����2�$�^R�b���2��Y��62#=��2�=ԕC����k�aJJ��Q��� u-���s�S�GU����~�^nV�w�A�;�+��$����z�T_��?�N]O���aobB�Wq�9�'v����G"�ٺ�pu'j̩%�4u�@q�3y_��1�}��Ty���o6i��}7n�7�p���+ў%��jI �������3�?֫/��̟w'y�p�A8��i$%?Ok`��E�ް�ϧ�>�W'[k�9��w"����zD��Ƽ4�Tʪ�5���5��ڷt+�Φ�~�vy���۲�g�V�̽Ѝ;�;�{'w�}���i��YڛI�q�osI��P|��vg�����{#��N;�U����!_#��-~;(|t���:�n�gE�d��-lfڮ���OkJ��i��R4V�tx�� �;��8�gDw�����t�����n5Nv�����f���g,2���[�]]�'y��(�Y�<�p@w����y��׻Y�NV+9��w��u��{dO�Fk8��g#9s�-./?�h����eU�}gyw����l���8L{s�0d3��`��pa�)��k�q���!m���u۫ڵ!M!���z�.�J�]����JdRC/�"�	y6�����{�q^G�|���P�bp:��"��S�Sn/s���xbq�LjI���f;�XbN�ޮ�2R��/N� ���s\���Gjh)�3��흲�xc������Y4}�5xN����hU2��J�&N�{D��G ��4��\8Tz��&�otC�NvWV����l��V:v��G�S���ޫ^-O~�gเU�r/-�C17��ai���"������!wuP�ׁ������{�L�]�B��礵�W,���2/���r(NWV�`Qk͛�����FB6{���x\E��.�r�u��]*�d���d	���{9S�J{,?l/[*�Ws�io�E���Sg6����2\��M���hbV,6��b��D�$b3 �%U�4Q	&�$�#I0`IÂU	� �y���j�5���Y3\�Mu�Ǯ��b�%���3�evCbN�.��,p{������<�M��W��P�O�>����:�̓iEMq�O��G�˙�4�ڡ^��F_d�a���Dk7�C�l�Dg�B�c��ba���-�|p$���@ԙ�o��W�o�^��	��=�z�����]0��"���d�a�x�ݯNQ�}�!�ý_�t��e{m���v�zv��gwɎh�}ӺL����l��<�&��@�k$ml�m̻,L���؞���T����ٰ` 
0�~��HF0�J�H�Z��Iv�%�D�#7+we��>uB�C���`E�{�`��p#$��;�$�_;9�U�7�F��Tl2��۾�]>y��c�g�DJf&Y������d��Ol�o����Uǃo�(��)���
�<�ې�*=���<o�>o)�$�O�EM4힑����=s�^�������u�?$�_�$�I�?��B(��j���q�� A�}�>z�:d&$%�T�&I�I		�HT��f��
` ��f��E��� fFB$$eRP	
e@���T� ��i�DI��d�&!���f@`eP���a���abB	�E!��i�P	
ed�dR�e�!�I��T	�i�a� aVhi�b@&��BU`���Y�!Bi����D��XD�� `D����H`�aE a `RB��(`RE dRA eB eR eB P��D��D��H��Hh`RQ D��HD��H��HD��H�� m
��H��HP��H��O~�������@�$(@�$@�$(@ʄ(@2�"2!�2! �0	�2� �>l�@Ȅ�@���@Ȅ�@�$�@Ȅ(�2	*2	(�0	(�0�(�2� (@Ȅ@¾2G8A��`Q��`dXF��``XE�`��`dA��`dF�`dX��`dX��`eE�XDd�*�@ʀ0(��@ 2"(�wp
�@ 0( � @� 2�
*�@�  �PQ ��@ `P `D eA;��������H@��H�"0	 �0	
0! �``R aw �!L�@�$@"@�$"HS �HB&��P��Hh`bB dR!��H��$ �D���?�����S��
DT&�H[e������~^���I���_�������y?���>���d�|�����������__��"I$�9?����b$BC��	$�,�O��Os�Ԋ�~������$��~ȒI�����~����%:�������'����rI���d�~7�o�DFT !R% X��H$�$A�$RP�P�HV$YD��	P�HT�IA�	X����Q�ID�	a` %BX���� �H	D��%A%D�$ID�� �)D���HBIT $�J!�H�H`R�J �
!�
J@F�E(P�D)T�I
��@�TJ!P�i���`dB�J$�	 d %B	FT�9?��^������O� �E�I	-�$��"I-��/�6I�������'�'VO?��&H�I�i�&�/�I$�ԟ˩>߯?�~��L��v�~�&��~�'����H$��b~�9�'�$�>�I������$D$:�I�G=	]$�=�,����'R�G���$��d�rK'�$��ޓ�G'u�{�ɒN��I$���?����$��'��I�����O����L�'�'�$����~�|��t$�@��������I ~O��=OҤ�-O��|����I/R|O۩?��?���$�O�$����I v�������ޝ$��L�~>윓�}�>�|>�	%�c���>�X����u�?�}~���$�'�O�1AY&SYZ�P�TـpP��3'� bC޾x���wJN�]h��E[������n�+T�PWL�4�wi��U*�Ŷ� ���V�ER�IQ��H�V���gm��:���B5�Yl-��]�k��Vvjwn�i�-*�ͭ%��m���f6�*V��J�R���j�Ki2��nk[f�hUl��]��i�ڝ�ѕ���p����:.Y��}d�ݷmU6Q�e�l�ƫMj͡E����cY۸��[f�dV����ʥ�l����iFֶi�Z�,936M��ij�J[C�Uv�Q�u��   w^�_|�{uۜZ�8�0݋k��n�v-�������r���5�:��z�J���s�Wm�T�8�\{�=�\�:�۷��޴J��w,��v�z�֩�l��-l�T́L�  k�}
(P�CCC��Ox��
��
/�xP�D��｡�r��Pݤ�s�uAJs]Z��R�ؗ�ݝR���{��h=)F��ڮ[���t=<�V<�r՚u۵Xֶ�il�W��)�ڬ2kn�  �}��a��+.��v��w��l��תO{����{w{s�g������՞��j�������Wl��p:�w-�S�ևn�����rl��cNC��j��'� ��م� �v���V�ܪ�z�Q�{=鵳����u;�V��1Fc��l[V܇'FW;.�f�ӵ�j����l�(��j�fŢ�s�ZU� �}U*(���*�6·N�*pN�wh�̦���ww3s�ᵚ*�Zʱ�(f.�vn�D�*��qÉRT��v�ٶ���V%�e��m��  <|�[G�������I���MUUP��V�P�  �Ӡ�3��ݎ�ܵ��
b�Z �t�)6�j��3Ui�,UZ��   �x=R�n�:�>�8  ��נ;�C@$-��  ݓ�A#@c� Pl�P khw` ,�ͷ����յ��5�P����   k� <�Օ�  ��p�	� iT)\� @;�k�A@�6��%@UΦ�R�upwQ  `ؠ)Et�jٯ�Yڵ���ڵ[Z��E�   >��4 )'ܻ8@]� *�wC�T 	�wU;S@:� (]��:	
wЦ�9��t$I��Y�t]e-����m6��5[j*ɵ�   ;� h]��T }� =4�r�4 u�p4��8ӣ���
�(gm(H ���h4��8  � �~@e)Q@F�OhaJJ�=@4 �{%*(  S�!��*   ��%U6�  $�TTڀ O���~?:�~w���~!����v���z�^5I��G#�P��@���u�~��>�>�����>__����m��m���������1�������6��� �_��?��n�?⿛�;2�-�ך&��:r�lE�6���f޺U-8�M=dTusteɶ/4+$�Y�S�l-�f8�Ώ�ҵ�zc�ZNB6l�1� Ǻ ��l��e�yR�BTJ�k[&�K-��kݠm	{��O ��'U�����3ˁ�ǈ�۬
 j�Z6S �v��;�Y�o)G�*X��K�ݹ	0�f�݋SU/-S$�vZ�'�b@�h3�b��s�I�UҺ�9r��;�xv�M�-����[T+@(3�,RnhM!��K5:*���C�H2�'*֡D蔓�3��/,'+�%͹����
�S#�LФ�T۫�̤�1�N�6抂�v5n�&V4څ�����`��6d��JH؞���b��E���� �{��I�{�AB��5[X���۲f�y�V��0�h� �t�ю��b���+J�3�[d�ܚ�����P5���e��]nc�IH��r1�U��i��iG��73�g2�%�V�Ŏؗ	x�0�Q��čZ6��u���i/o6��V ��ꈴ�V�q�[��nJ�Z�H����;�܎�*���ի�)U�,�	�C�Y뾦u���VV6]�%��b�D�*�r=�2F.�2�)�u׳M�2◲��M�������+���^���.E�:��a=�݋���22�Ң��+�Ŕ희r�ͭ����im�����9W�dP;z;���E$�&�S4,���,־�i��Z�����1��ޭZ�Rm�VO�#��[�l�jh�z�������7u��a:ݲc@�tk1S���S+o4Ah���V�$ �ih�F,1Lr���#��Q���2H�{L�R�z+j�j��5���i�'/wD4�KT�����0�D��Ws2ܵGj5��ƍwR�۩�f2'L��-!L����h6�e� e��Sk]�Q(MX��h���NI�lf�"�K�u����!dA�D��5�Z�w6*������MGo�8,�mlMF�X���=t]Zݘ�-^b͸�������b%j��IdyM��f��z�ojh�aR�6,[�z.]Ձ� ��s`��[�{E�e�-Ltd�fb����BI�m�K�+_2E��q3�g��X��U���&i�p�:kh��m+�A<U�� �1��q�D1Q.�J��ޜ�%�:�sD�h^�KC٤��a���WVM"j=��ȡ�3FXI{gK�Y��F�0�l�� +xE�{g��MlKV8#M$l]�ݍ�̧u4�!�9K	K&�l㰯3*kAov���$vLז]��T,�KOY�AAM�5Yx�M�n�~�n�+��M�V�w��Hkr�9{�:�2�ȳG�N˕0��e��:����ad��^L6vT��l���Y���-���r���r��Jz7^��-�$��r���K9V��K66��t�[�Df�H�:��f<�9��[������6��S�2��x�sjK`)��X�d��7b��وhӷ�,���-/�t�7e:FhW
�M��h�Ak�7�n=�R��GZ���(�Q�G�BR�^[�fcj���R�^ն&f�X���cL�N~"�$L�6nn*q&����%�uk+��3(�"�K1c*���ߴ��ň�+s4���J��ZVh(�V�9iej�zw�H�5���4�i]��iX�Xp�Cqެ̨�+hX�$PQX
�re=�+߁k��s5�e&*"+/ �q d6�ڼBa� ����Q�xY5��3~uv2��3)�
B�=�mA�'A�U���tPP8��V��cL��8^]G��ܨu8
��%wR�,�Ʈ�`�u|�x~n���E�Y���٧mŻ���pmV��f������bi�b�M���.��7WN�GLd�B���Y2�ó�A���X�*��D��M墜�E���J����+o���P!A���J.Q�OUn�N"�9�X��B��F�;j�7�Ɠ�c��^�+
�Z��7C"��JaCKu|qY��e�y�Ԇ�j��Eӂ-��XsE�%E%['��el��dZ���l7���лj��ܢ�	��(f8��Sj2�+b	Y��#UK��G˫��B�Ɋ���.����@�f�;`����0�O+k�#B������LN�R�H���������y�GI�S�cF��j��6��b��J�
R��y4TW�bG7��33r�^�
*�e�w���N!z\yr�X�
Ɠ%�۸E]��*�ܽ�b:M7`O�V��u�օ����lU��a��BJuy�f�K�lHP�3Z��u�ړ���v����
�2-P����a�ϡ�������&G��:%���ں��k�2��f�̩��T4��s5�6�^P���3!KO�s1x���tdƪ�ʄ�'"�tP��U���fژ����t���Jֻo��倛]Oxe%�u�Ѐ6Ke�47b������z�6�ҍ�n�d��{�jh߲l�<����o��B�ܽVu�.�Z�fЙ��zś$��� �%Oh���fVI��&�tp/�(��6�/S5��l�����Zі�n���b��/%�qA
wyN��Q�/���H&��f˶C�oZ��V��h����[X#��²Шa�bFjz�#�J�Sct-$�^$n�j�"��Ҙ�	u�"�Y&��IҚ��w.Ŷ�r�AjD/�Yc �&�|қ�iL���X0[̖� �kuL&i�Jb��t�Blf���Z��FVKU�S%���-��@]���t���EiԨ��nYOi!CpQjحZ58𥕰���=[�s!J�����\P��se�p�6M��R��,���ZmhN��mھ�o���// oFt �D�Fj��7f��2n�r�mk 5)mY��w�h�Ug��l�Aiz6GK-!���ь�`���0�܎�x��e�ח!J�Y���Y���'�ȡ�V���I&��4[r��*�]���j�5m9��L=�[�\օ��rh^T��`�;yLmҢ^8ٽpǄ؋^�O�X��ɻz���1���JT��Os)�њ /^]�Z�+
�3⚕�rI��L�w!���6EYv�������*���A�1-t^�i)�I,�CC�J��^�F����l"�)EiԒq$f�.TE�����2e�F�7hm���n����w@�5*�ǋ*ܡ�1�54��l�0542�7��� �V	�,0��v���3f�hǀGmm_�aLxҥ���cvh:Z&n���`�i��J��M�,��w���-��(��!v�!�T�TU�bPX���4f:I��Ȭ^j4?�B��-�������F�NJ�#���������3a��;%3���K�@�/N\Tņ��;l��x]�n*vn tQ�ͭ�Y�ע�7,��a�S�J��	Xy�"�U���⒰.ei�v��;K8m!T�N���]j6�2��GfJ�E�r�Q�5j��)�T�'�C�K7H�m���e��N`:����R���p�����Ɋ�M�X*��m`<�r�ґ_=���j�h�&n����.˕��ojkn1Je�[���sSU^i&��o���VPӮ� �:��c��CB���w�e�ņVAY�j��iJ-��):�2@'f���2 ���4EJ��f0�'�f��w0e�/2 h\�C����R�m:�wr]<��&���oK,<<
�*�u����"Sֹ��V���LlV+x�"C+iCB4���xCڅ�Aҽ[3E�DZ�m�(�
m����7X�+Sd�-�$p7
6���3%h �"w&�h�@��ojׅ�х<�(�Pi1O���'I���4,/tę�-٣��ӰVXoE��n��Rk`��!�˽��yP�0^�긷v�����������F�*���u�D�[�bR��j UֻL��h�v�xqk��#�F�hc���2��2�Q�F�.�C@�̥Y[��J�v���6*��"qV^[0�C해+,͊�����n=��TA��`�/[��HAV�3a���������{l��(,E�R}hle�{��n&�ܴ��c���֌m&MbWV���iVM��B�F q<��w/e�F���7L�&��@@�S�Yn�X��42�P+������B�]�M�D����ؖ�j��0����RX K�V�1H�M��j]B�5GV�pv�fQ�6:P��`�7QI�Z�*n�@�� �f�j�<Q��j��Z��[�j�Mm]��c�u40Hʇp�0��;�b��m\F�*��ؿ�Ŭ4��K�p�	�̧)P��P�V���.�ędh��i��jCv�J9��U��{�^ͽ�RQMq:!cA୺��Î�2��Xݗb�J0�{��4�x�9H��;���T�jT���VÑ���像F
�+n��;dU�B=�r[�ܦ0l���f\��o/ukl E�6��VՌs�P+M:8N�D���OkcC8���A���Me��**�1�D�FeI�q��� ����n|�*vcuh/�BVi���=�W���Ӣ�wQ�<�L��4dgpDR��y�e��Bhmb��R� t�,��If^���%����z�x �S��g@;��POf�3��D�g�F1f9V��?:Dl�{6Rnh������2���+�:uXDd�މgMnޕ��QT��D�G���U��F�YN�!��+fP�K�,���y�k�W�V0�x��ЕML%j��I��r�F��6��c���2F�`!��d�wJ���V)��@�3n�.�Ò�#b�k���)`GX �!mHoF;�y�^n�f�̺����Q��tV�Ɔ<�x�Æ��J�����/j� ���L@j�yd�`3n	���X�ҽ��d[D�PFjAY��-������������u�q@�b�d2� wO1�4r�d�)�*�vp������k)�!���
V71Q��7P�����e�D.^�#�-�X�i��F��b{�ɶb'N�5�jm˰]�:�;��A��b�I�#��9��3*�e�`�������c��єv!)��p^�dF�������r�[�ڂ�j�n-�4�/@ ��B ���6	��E1�Y�J̽i��WY4e��eju4ff�r�#W��4^�@��bƥԧ�w	G%hdFΨd�f�E֘!!����6���6�Թxh��^�z�4�%�*$Sg._��ј&� #u5��O6�a� U6�m�-�ws0�;8N�nM���i[���r��V$�\�E����O\E�r�'VaՁ�Ǻ!�B�:X�9I48vBnE�wsm+.�ɄZ���a�n;2��Nj�2��x�U�慮����W���8fPbփ��*̋`�M��TI\N:�F�*��Y�Ѳ5�Cr�0��y��u
�Y!��H����J��
3�u)c�mA���Z$
�Xַm��'��m�Z��BD��ʻh۫�c�5��.V/6��Y���2�(�m�L��W`���W�і[5q2��.�JS�*�l�)�D������NQ���`�L����6��F3#�TMA9dLQ3.U��w�P����MO���z�F�b�M���[�i^��r�:ݴ@d��yX��.K�Av�Ɇ*�//>�ۣ��}� hs��`��ml%�V�41�	B�� r��v�Ӎ^���;B���S.�b(S�嫽%�.��W���ـ�hăt(�(AӷĐ֯K�̲�Q��e"'�(f�L�Ycv�^�=HҺXu3Z��I«i��w��O����+��y�)�I�g8�.�w֨2���Ksu"N�a���#f˼"��%6t7N�?���E�	���03��܄�[�HHh�sҊň̺0��:�:&�*��~gZ��>&��)ޜX�çh�E�I���	�n���*،�\ �'�M��t��[(v����������SZ?R�7ze٭���l	��Jb�E���L�Ff�;��%�1U�5��kc_mMYL�ƴ�*'�if���cV%�e<aK��BY{wJ]�7�3��O ���.�P�q(���ua+*�q�j�z�փX�n�P�2�6&�À�\r�A�²kh��jJy�nG��p^�Π̊*�A��d� ]���Xp��.�q�8���tF��;7Q�Mk�P��6-aP��H2E�uym��`^��C#7�#͠~qV��)D(�[����S������$�C�4R��v�I�T�r���&�6�ʍ��atEmAR�n\�:�5E��y#B��lX��\����e+��nfm������@�^�Tm���/��m:���wSeV��RN �X�lAє����:D��hnґjF�YR67դ�w�&�R\h��\�*���'��U���qs+/�۔)m 5Lu�-i]D�3i����*9+a��JH�b��z����).H��$�ìJ���ݣʯ�f8�Ȃ���⚲D�]�8��ч0�,�����:�'�e@k�P�4�,P;�H��[���-�U��q=ڻ�#IAx����R�z�M�.�̌m������Y#yD%�TE7��le_J�5&�%���+	k,��4��C��:��.�P�Y��1	Y�;��J°��a����K-h��w�&]��T��L���Kk���ٲTE�r�Ҩ���t��R��Fv�'2�����с)�0q��y���!�s5Xb�]��#7GU���J���9XX�Э�b�Lb�#�-�]�F���x�6"�i��z����Rbx��@�oq�s���i�f��V�ʼ����7���m��8�Z�_�[�r�JT}Z�j4{�2��9�C�3*�u)�tj��+%��P�$6��$�n��9W�!{e��-��N����hn��*v�R��T�\y)H@����^T{��c[�-6����E�4./� r�I�6D��R_o-(��)�mi�-���U�tp�yuat�1��K�Be��ZnV#�a��-�S>�J7Lu5�u�&���y��t��}���w��u��5L��E��6fht�tb{�$M��|R��t�u�Õ�F+k�q8��TI�uh5��0cvK�j���Z�l��Q<*�7ʻ�u��t=�f�]�)��hs����*Ա����8���;C �W��7����U�xZGw�KM] �n�2��/K�N�[��R��;	�h�J��7{�����J�K���m$�Y����ڬ��
�����%֟�v(��
_Ym�Ɲ�[/�2��o�җ�r:;pq[��n�:�i��\?=mή��mog<M�� K�w��T۫�=��q�i��\��\�ԽI�qS�e�3A���.\����s/�|�#�"��Dv�AR0�Ū�ǵ���'�ܝl
�&�Gn.3�7RСUw��>�n��?J9'J<�l��v�i]�ޛ���S�e'���6e���+&e�I�<�[{\��mGA�֎\e��#u��������	8����v�]܏-�i%Sn��6��B��a��>�u�~�b�+�$6���^�&:��,	�#����i\���oAf\���w�lp�[j���v*���Z/�zxg=�SY�'1wO0\ޓ���MS,ʽ9˄L_#/2�)��"��zg
�3��ytWB�^>��c9FN��4��WP�'20h��>Q��WYi�1,*K ��s�W�8�S�ɚ� �`�+�~m$���P��ٳcC;i�yS��h�+�]O��yHgY��J��M1�sK��#�8�64�cI�T5E�k8� ��t�Cx7��9 ��Z���m�������lc�Z�T�a�m:�
ɶ��ab�;�8�2,݄����JN���hY�f���`	�;w�5�()�Yz������Zֶ%�z��-(I���V�"��w�Y�����M����o���
��ǅ��\���]q(�w9��&�ni�i��O�+t�:e��z��ϛ0�ʛ�����.�n:ht�r�4n�v��%�;{�)�E�F��!#��\�o��=��Ѡr�$��
�r:���͘��=�Lu�J��k����a�\wL�-��(�]L�K��ې3(u�y��8wi�.��su;	�	�6��D��b�������hn�_b�JS��PG��)�f0��]밫��9(3���6�R*��:lT��gH�N���Z�L<+����6�}0CY�R�&�Ykb�Y�A�4x�I.�:�av)���� �Y�XFܭ��rM��u�jȎ<A���.���҆��!�r�W�|m�jL��s������,��a��gZ��M\�����ۏ�V�3\R��ds�}���*3�-j���q��g�~���Y��h;G�n{v^�Lg�m��땦���YoU��%]�	���P��:`�K�/�vP
�]{Yh_g��D�y��%��v�Ȗ7@�ͥW�ZyWK�Q_H5�2w=k����)����[�ҍ���&�!r�_X�9��Q.��B��^V�MCc�D�@�A��P����v�h{�	��d�Y�+��y�\�zr���|��"��u�;S8Ρq�,�Y���}��C���I� v��4ϋ��D��5}�3�<��%�}��&��Qr�!m��j9Z�� �:���'(d�+���	�w ���wh���n�bxH"�I2��*�[��˸k!r'���x:Z�EֽX�5g���A;�Ѥ�y���/���޹�}���m��2gǷ��0^�є�Ա�%4Xo���Uz$ћ]	���F2[0a�˻��H�h���Cl���8�1�����E�D;t�+:sB/�9������%�9�{uћ�:��-m�!S�4�t�����}@�p��Ңʺ;�y[�e:�P�1}}��w��Y��ҭ��ĸƩ%Wݮ�,䎴�pU�6)���1Jkh�����Z�w�n��֪w�46ū����'9ձ2Y&����E�K^:��0G����|��"���#�@��9w�Q��f��C���NmI[cEʎ�p�Ǌ���az8bܩ��|_:�!�Cُu�z�Fe��n�OF>yPW*a��:;����A{H�$^Tn���>e�$&�ַ��% .��:
V�	�����0<T̠7\J�
��_f d8�U(�*��Ԫk��@]ޜ�8,��2pR�'�>��tɿG����*�x�j�c1�Q_5挹��Q˗�搫'^Փ]����]9ΰ�1�YF���	�n��΁l5[]+-19|4�V�%-�R��7�]���m�N�}�m��c%g���҅Y�� �{���Em����G���_j�6���fvE��-��R���XF�F�F�E�9�7��\̛��M�ڡ׵+rl��{u���7<v���3JƐю�c�Ԭ|^���[�����M*|�C���&�Ү��n�:��aS�KO�ѭ���,�z�]�(dͺĂֺ���A̚���t�B͌RwGSs5�j�y���*}|~tu���kgEv◨�����f�]���5���7Z�u^�D�+�Ƴ�>���gNë
	�kFG���[�s�[|Z��!`�N�]�oC2��BD�J�pc�д�E͠�롒Ԩ�Q�`���.��y�k�	v�差 ������[�P�0v��$���k�@H�A�a�3y������k�M��W��畨<nݙ��ݺ��KO�5%��r�h��M���=�z@�[e�GP굗O�J���}��+e���wO�Hi�Bs\�U%�3��]`�IeN�UIv1ҫa�z��h!�y��k�2����Ӝ&����5�7���.�~�F�	���܍��6]�l)���Қ����CZ��ؤk�֠�G;��E�90��Q������NR+%Ú0ct�����(]�rxC��[�
oeVZ�ͼ���������r��2�Z#io[\(�\��C]bU����c�I�׺����C�q��MӰZ�]9�7|�N��Ĝ������*}���G%%Q��L��]�B�s[��h��wf:o6Y�TޝB{�aF�ѵ�B�nm	���څ�Bܨ�	�AR��!�Y���/M��R���幖���(�I���'j�w6�ەm���U���M/��md�Kް�:*�좙"��1xT��%��u;'n�l��n�+H��<�p��E��5e���L�N���Q� Z���4/�:\�����i���ɍ�7��Ͳ�sx�.|�/d�.Z������6��M��g;��Q�����͊�0�Ce�0�<�>O���y�����}i�௬'ej�]v1^�Z�p:t��n���'�]ŉ��8��M��DXxx�M_m�Vn�n�ͫG%�q�B�9RV����W��1Ij<y�؛K|K��8Z�[�]��u.�L��Lv����m����bN��G�X 6Ѹ�^�Q�6�ca�Z��	��prĞ�*\)�IV��No6��t����a�tͻ�ħۤ�[�$�/*N�=,QN:U��|5f�&$3��+&�U+n�a�Ev8�5��uhڵNԜ�t��ۄ�x�H��tc���wDq��6iR�٪���:o��]��JZ8�!pݻ�8�m�e�d�V<G���f"0;J�˾q�Oo���4J�����S��&�K�SJuvs�mp�E�۶b�u!��v��7ܣ��e�ͼ�4��u���K�0�ۏ�Xk���������,
�1+��*,�5��ͦ�?p��L�����
�ms����tv�}��̾ܥ@6�έRk����VZ�}��-�;v���G3^�[;b��4���P�.�}�û�y���T��\!(�eK�\G[R�gE�v��'�-Y��zR��s��i����#p���\Yt����
�*M�o%M[��UM�����Y�7�����W�^�BjL�s�"��Hh(1Wth�k�|u�Z;U5�.i����䣧,��f�*��ү[�}��tR�N�Iѫ�
��`y�_;2��T��)�Ԝ�v���W��+��T���P,�{	�:̋�5QUݚ�=l�J|6�'65vm\ڏy|p�/���7}inܢ�<�?&y�ޅ��+cz�T�o\�Z�˛�P��sL��n��Z��F��úb�yɁEe���nTb�j"\�sV9��� W}����r�aX�	;˩Ҍ6�sǝ���tPˍ�U�Yu��+�)�ت�'C9�y�{�0'M���R�xI��WK�jۺ�=�%D��쳡eu=�H�%v�1y�<ͷ��=�30��]G�Ԗ�)�4F���U�S9W�1�$ݭc�L\�����f��������?*�^�W�9g!�9��4��<��V��X�6��4�Ê��%�ۮo����ż�����:�j�Wj�s�.�ʾ�Q�%1C>�p���fZYmtmNe��8'E�q��=�s������0��-�]��5���X�bn��"�O��Up�T��M�
�<}X������wXp�Ʈi�f5}NS6�i-�>�ej��k#���k3�XX�ඇQ�u��7��(�ݞ����k�\����r�ui��il��sE۴�v��5�S2�����S�{N�AZ۰�b��]�%�VS�h�*mc%8��V���]�Y���Z�n�f|��7	��m���ƴ��9WJ�u�#�K�#f�SF�x;;I�F�s�&]��Pj_fG��;���ˎ�1��Y��I��7��B�䤀���lŶ�L��R������Y�ټ7�S]Js]f�:v�#�[u�}�A��Ңg5�^}j5eWj�ē���K���j�/�M��Es
�c����K���xq|!�H��s���%@�G�rf3[��a�D a������N�M�9��!���[�����Pm��r�W6��PK6��`o1��NK3
n�$n�_d�nt㸋3:<%PJ�WM	%s����ڜm9uwD$[��A���Ѯ�R�j�>{g�f<qR*��L��^�}��l"�W3���U���m<� ��}�h�P�/vqh�7�����κ��,�(��c<J1����̫���@×.��պ�
7A-�k����?;!���ޓA��-#x��WwvV�.���$$���1�lnO��gRQ"�����x"o��SʌR��`��HtV����9��y\�t�+ �`�o��w	,t�̜��>ţ6��Ϝ�@��f�
��
����4u\?m�]J^�ܹ��E�D��o4i�]%Ⱥ���lv�E��Jw �>���\�0�c����"� �c;{�>z���Zu���^m��
���ӽt_��#�&2����K�٢ZJ&naY�	K*�S�AL�ViF�1֮`츳*r�u�P�YR]��%�)�y�1.)��V��M�С�8m��C1��w%��g:�v6=ٻ�qH/+hM���ᭃJ�M��>�ݔ�Cf�&��2#��0o�4�*m�#4#���o��,f	)w=��:�HH�%�-�g>�aMr�KA܂��ŭ#`��3�os�����X%n]G&2�\�^	Zc2U�囎��fh�f����q��1
ǒR�%s��}�l�|ĠZ,,Ff�$�&<s*��q�
#�������#|�5V�W}����`HM{��Vwra+�:��i�)�d��,
�����v��v�KS[&��e8�3hו).(��B5�{�1�k�S��Z��:-Rvↈ���.��L1#�#�fp��������1飱�N=�����6�::��ܥ�2�knK5X������x�aU�3�Wј�2x]�x�hQ�W8f��V��D7��]w1ki����e�(fe����=��퇖�p�.p6l��݉l��
�64q>��;F�cV�O��s�	���jʷ���|j2���o#��.���:ڼ�Dr�#�r`���S�t�����S��C]�9�L;��N5u�녱)d��kV[���wZ�0L*�wJr��ˌ��ڧ��<�1Ԣ4�+)�rm�oԷ�i�bY�x�R��^�^b��������_�c�3C�3���vQ�YFd���NAݜ��g� ����i`��&�w�n��u������frZ����:,I�ɣk!Z�Nf��n�6�vԺo+��BU�Rֳa�G��ɢ�5�]Y�jP���3��IW���9R&�r)Y��5՚J�\6���V���F����	�̂�r*X7���S��O\�{'d)�ᠶ����o�Cgd�E�K��SP���} {�m��5�}�ۚ�c�NԒb o#2pu����u:ln����a(E�;O�FWu����	`�]`f\��=�����sy���Ԛ3Zn��<�̹�z�.K�׫7p���o�:eﳒf��)��-�0����fV�[GQ+�[�9f%Z��e��;v�7����'X�=�i�;���;5ѐ��&�� �k�u�*��lŃB�}�!Կ,��{�B�}�ؕw�I6�� ��c���Bq珦��/��2/�7Ԫ^�N�ί���<N��lY(
Ѝ$��j�S��Z��k���*+Y�f�P
���jk�ۊI�f��x�]9�=N��w]��	N«�i�SN\���m9�;�rR=��#�(����U}�W�U_R@�c�`��6�|�����'x�}<x�������h����2۵�d���DD��(��VӤ�~�W�����N����	�N ˱G�:4��4)A�f����˷�:t����Q���oZ�m�U���EHo���7�N� ���tق�m42G����DW_��gʏ�����K�r��L<a��-XD�t�ʒ��G���t��IwW��}E�x�s�B�R�b����[y�ɀ=�}�����h�n�G�ѳ -땰~�Ix�[��E�U��G"��n�����tһi�-kK�s�]��3T��r���Ѩ��kz�w�7���u8�)b2�B�y�Aΰ��V���{���A��A{���vM��[K7���X6�;g�T�`�ڥ�G�Vk�b�ayVZu$ ���u�PfT��E+�F�2��"��qt� wر�ò�!��i�`Q�-�`���N�㧔������pty�K�ԄwB��h�8(G����T�8Yuwt2ut�v+z� ��t�`���,=�4K�F�����;���Y�K� �gb���J��.�1]P�&N��uG�i�4V�Ha�s9��v@oH����Es��d%{t�}�g����B�{0�[�GN��Qz�H;�ZIn^���쇨ɒ�
zQ{��]��f_&�sۿ�7�:9g�����;l7��
��B�	��Z���t/��f@�*w�9��f;T.� bh��*�W��x��P����ĳg�J��k��vM0��V����o]���5�"���º���*�纴ܗF�n0�8*K�R��)�M��*�l�b��dyښL\�}rZ����wp�ʶ��t�3ho��zeN�r�����8i��wyK�����"�L�t�VU�J��E`E���}������C� b�xF��wL�겲-9��bԫm]Y��COe2x!f|�`�z�i��̨$|j:�'lq[�d�h�oΟ^�ua�xk�- sksB��S�}PR�2�(+vӤm�ɵV�THΥ�Z�����T�,_)Srl4S�s��ަ+�2���;M�`HWp,5z��cy��Tf��;�Mk�X�Ղ�
I5n��f��[�fK��}�)�����!ʓX�!f��3Vbl���JW�gL$��Bc{���-��E:�4�حry��s�/�%l��]����.*މ���.���f���/�w�y�&a#������42�6Y/9fs٨˾�iҹ܋64Sy.��W[	4�s�v��"$QŜ�*o7֫6�'Q�d��F�r��#���0J3X�fu�������)ݩιպ k4��i���R!$D��|�0$+�V$A�0�G9Vʲ��>�^[C�yڀ>Ūf���'ny!}���wB��=��&����K)���K���r�!�l��o�w.��]Z�ηC��.P��.�7^���A(:"�%�R慳ܡ�bdےƜ�4F˗�8�ئ����wM�0YB�u�θԦ{%�{�xU����d����S�=Z7YR��v�So��9c��-V2�N�k;9��z��Q��Ռ��46���I=4k���Up���)cfRu��6�Lq��'a��n�UZ<�,�Ŝ��!�E�9�����:[�̇}�P�@^���r�!�m��A]G),�b[.:�ҦL��8�(�fv���R櫾��� �=$^,�Ɇ�tqA!�/3��lh�Ż6�ږ3�d��BQUkh�U//lڛ���m�7��:��v"�v���s�f��Ș�6�j��B�Q��}�u����Ҭj�n��ąp\r�ݣa�	j8dGg-�n@.�6vQ�Y-ueq����Go�vaHͽ�m���Y�Z{d���h
��luY��(��靽�ݱ�X^7q��jŧZT`P�֌;VQ#w]���`�r�U�#���
�Ç���t��Ԡ�iJ��� ^�t.n��A1�gvPb�j���QT�nn��Wy1PR�r:�6�M�0,4��ZKTų%ӡ�2���|.�U�;;�oS9�`t]�{Su[�i�9֘ �ic��Bj������#iK}�u�Ł�ȡlU��sŭ�\� ����Գ���H�N�k�^k����wl�id�l��g�4�@m��e��]��y$����P�M̤+	�����-n�2��Ǩ��%n,��{��̜3&=�`�-�-M�{o5;C=��"�J���y'�P6.�vv͘�U�ohk�✮D;LX�T����Z��#j	��W>�Zb�H���{�e95��؋����fK�f��ɼa��B��S��6+�^=���ŒΠ�p���t��r���L�}l>�R�Som��yl�R�t��Zz> 	9�[�o�ӮB�zT��/���HI��]�1K����;˯	�)ёWlXc*1lʗ��@kf���v�#sR��QKU��3Z�!��jK�u���z{k���{T�7.�j�43��%'�;,Ϧ��]�0��Q�9e�b�{AB�����hq������pj�,��f�굼kL@�;��P/�hm٭q���c�5���(:Y�n �R���m�ܨH֘�K(��n'��4M���E�Gϝk�� fd�:�:�|,��\˭�U����v�+�g>ёי��}���uN=V������+t�J����2M���1�'u�I�a��5D���L`�����L��z��DH�6n+c)�70�Ǐ�\;V)��kg:�2�a��ڿ���<(�b�U`:8o�x�U���]��Sz1�ӏ&M�n�U�;�����ݶ���wa��wC��2�E��`։PT}��y�#C/��0� ����0��4u4���SI��O-V�ξN}�ۇ ����{}��[��)V#� s+]Y23��r��v�P�\����J��,T��J��5��B�޳Z���Cv�͋��ر\����G�`�7B��������<�ht����_�S��0��1����p@����Vԫ�.KD�M��WYSn�#�i���>;���׷��&
�]=�ًV���n3����Ud��6ؒD�[[l�0V�	�㾶E�3�U�+h�WNgFc��\
�#KyJk�Ƅ�����-9q��V�Z���#�3sKxâ���(��7� ���aY���326��b����[1�/yrY��(>qj��;!�#�L*����+�R�X;;yP�m��զ��{�Ìa��h]���\ڣ՗��84:�W,�{�E֞��fWN��	����p.�E��S% ���;����R��L��[������5���a��ooWTY��w"��GS\��%@�j;�����,��Y��fuc䃾���J/��tX��:��p
�C֑��64��C�)&==%��9e	��fgc�#��VO �`����p����� �9̡Q�=Ƕ�or[���8��6s���s�N�]*-.�aO���.յx�C���g#n���=������N� �`}���4�Y�ON�Q�ьy�� ʱs���5_���g�9.NJ=��e�fZ�C�ڻ�{W)��4�L��k������e�u�y��jx�=S#�of�5d�|N�57v�#����,���ڊ�X��Ձh�L	��`�'\z���h�,���L*jA�TQ[�-k�n���T��s��T)L=۳j��g���u�����R��NV��n�GI��#ٲe`t�Q@�[j�pl}b��:�髵cNȷ0��CyO��Q�G��#J�����Q�J��"�5,�];nP�i���ɣ&���S��+8�U	��눎"f3��>I�1��)ۈ�1�c���.j�\����5O�k�ֻ�-q
�L�j�����n\������>&�;'�'U�9�͎f��KfșӢ�{p��HN��;,�*�=�n�M��W�,Ǌ`�W};�p��J��/9��f4y�}N��y�8wn�Md����.�W(����-i�˔xY����3���p�A�8��(٤"]����Q��@�h�{�cpݞ��w�*9qhهA��il7�Ch2�V�P�zL�鎸�J�X Ԃ�
쐝�î�ܸrj�v����I��m�vJl�@��s�n�ӳ��{���(��[A+��.�;;�Ư��p�q�s��ٿd6U��9��+0�����#�`�i6k�)%A��q��e��[��k�B���w%՛rеط���z�j�{zQ�,�<]d"u���T�l:��9y�2ё����.�ou��gi�7zp%�a}��V%��L�����)|�w!v�^2��;�Ĕ'K%e�pL]��N�{�b��o�PB`,J"�f�j�X�s�k�ȧ�������`ڻ��<�v�l����~r�����k��ʟ\�j��ؑ9�x	�xM-�ɬI�0]�f�Kʺ:e[(k,9�f+�F�VM6���edn���*Z�@	��b�Yϭ�t�����_S�˻8�l�2\�S�aT2��w��ѳU��9s���M�K:��9�`O�T��TFfYb�E���Vi��ӽ�
�	�*ɝ�͑��ï�]�v�@uoe���2e:���T��Dr��� �5r��.��Y�KR>��y�=�͢!�᷶�Y�ݘ��+�J��5��=M�n�a�cE��!Ҹ�h����Iu��of���-�JcW�U��Yg������*�a�(���:͙(��blɗ���ai���6$�J�e�3��8lwbn��6N��s�W�r���M[���x(�Q��V��&�����+�ҹ��B�tZ� ���wq�W���֯x�wx%�mEL>|�|{�l���hG1�t�[5��	�v�3�(�r�ۀ��#R����K+P��4�(PK:��]7��Y���}v[QY�
U���m 6+r|�e�>ҫa������k�ܫ�N�U+�M�s��XCIʕz|��T2+<]D�A%p�,��fQ�S!����w�n�Y��Q
�V"D�FHB#��ul2s����'Y�Ot����SP���E�n-��9K�o|.��c�%.�uY���t&���K�)��Zz��m����8gE{�卽�`Y��V��I�O��Z��$�m���M]:����X�-�.�h�Ç�6Ƨi���+�����x5�[����	�_oE�p.�ƛ��A�� ۂR�@�7�J�ިśW]eaR^�d��iu��Ƌ��ћKN�h��b��޻�@V%�Qd@t���'�rﭭ�y�3)�an�*EM}��-�.d�ގ62Z��ݤ�ʽm�s���U�3{o�)�mp�U��rl�n��̸�t�C�E�]A�����[��VÔ*�n�X����]�{iY����uP�d�>�<����P6�h���1ɫ6l�b.~�˩JEnh�b�Uᠧe�h��]��ۭ4���	z�_0�#ͭ��m�l�p���+�T ңu��Ca�L�2�1Dk��a�
�>�gZ��l��������z)J�ٰ�6�#�D����WS�{s�cVE}�Ji�1�'@�lp�31`nn����mK�Y�v�G�΢Z�u�j�Z��;m`f�9�$�Vuj�qYz�`����Z"�qE� N;W:�ꓶ��8�b�.2y"���R��L��K9\��,�P:r'dq�n�&�\P�C������|�Z&ӟ-��Ԕ���r���Ue��z@%��&"Cɽ)��1n���i�hԺ���o��M5^�ڀױ��-�(�mqT�3���cbv<����*T�3�a�b������K�w�����eszܬ�a�Xi]��)4�}���K�>c��U�cjY����۱��I�F��!��W����`r<6�{4`w̹n�h.�q(�U����=��^U��Ž*P�;�$�K�Ǜ�ƾD��,w=6Yb����_X# ���: �����Gs3���Nոې&��m�ݹJ���f�C^>&#��]��p9Q�GwK��v8[�@�5��TnY̽K���AiѴ[z�`Y�r����Wk��1�gA:a��:��Y�+e
�f�h��_NCKs�V�Vte�B��3`L�۱�]E(9������t.;=}����8#ǵDP�>J���k!�;���+;�'Q�Ym�Io�g*k�t��w7)r�(=���ٳV����e��? ��=B!}M��Y�t�GyqU ���!T����8�c4t�sL&d��%n�F�BEM�T���`�-�+y6���v� z�r�Zj��䫆3.��R��m�$�X�C�mp݉Ҭ6#����U�l�%�4�49����.g>J�J�e�P*�sru��Z�nR���2���v�<	��T���Y��ݥ��������3VK֤�h�lm�:��]��U�1�����m"��]�5��su��hr������d�/gP8�p��A�9��Nĥ@�Kf<��r�X֗�onËh��n�]uni\Z��f���䔳k��A�� ݝ(���?�}��,�:F\��Z���MZ-:�鯷�%-|lo[���s���@�v%X�s�H��h�J��v����r)�D�l�M1(I�s��")T�f?�&��E��,Ƈ`�ˁ���U���Y�f��$�%��oG:p���ۧ����r�z�����yΗ7z;(��e&{]�`�n�Du�tDs ��+�O#�^�K��'D�T i.Rej��>3(P:��-�n� �}F����%ZՑtu9 ~Ǝ�cA�����
EƙNV��:�MB�c��1����6mU��y[7y�X
�i&e���V���w\#/�+WJ<�yRV�<��A��)�WIS�n�٠H���]mQ﯈+��4��_�꯫������JfU{b��|�b��T��MԵ��
�J�,�w��VL�q��7�Bj䄃��tdEC6�ǚ�:n<�f9G0�\(��:ao�J���81Tۗ�	�����J��R������K������E���r�|ܬ�["�պ�;�]@����7P;�N/�S46nJJ�pM��iP��j�;�}�N�v�U`ۋa2j�t�B�qQ�1�*�*���\��e�胦e���.�9�����/xXn�V�&]s!P��	ۖ+�_m�o)BM!N��dFi��#Oim�YB��ն�e�veN�4T��vk��ܙ�H�a��N:��oaP�=B�ђ_A�U�-k�(ӵ*Bv�p�@n��Ws)���n��U>;[O^��x�;^���éR�zcK����[R�v�5��D=Bë}��g��/nnu	e9A�b�r,\�V�V��o��x��4��\�:Ɇ���,LO�{��S�U�^^p]
a4M�0��i�������"8�uŏe��L�Z��zL޽Yg�x5���z8v.{w��e�U~��4s���qqqʕ�)�
��[����t6�<ʺ��hmH���Q�]��8Jӧ���3Ou�eKE������o��:ʋ_:Bz�9H�h6�<j��ֳR��W[�K�[%��}�ԕ�*� `Qf�[Ѣ����)M[=%L��l�ⰷ]�e]6C�^s��f��ߞ?����=���Ns�ueEEE�%!X,�s9�\�@��Ҿ�9T��<��J�r�����=b�x<
x�UEʈ"=+�܇9�_	�*"�%utrwJ�L�Օ�xNs��G��9QQ�*T
��V�Z�I
5&�Tn�EN�^�EW*�VeW.a�UP^tr1 �,,٩�L9<uè[#��ndR���:uS��H�+G>�iE����V��_�J��R(�^rˑs2'2"������IUQDp�D�J+��EPd���VIp�2"�7�Y$��=n5XiK(��DvzҨ���r����B$R�3*+VA�I*�f�DQU$,�����<ܓ�"�����)�!T�U&QfFBA)β��*Մ��A* ��D��AQ2.�S���
!D�PUQ��r��s�"���!�	g=��@� ,w�+r�D֞���f�6�sdg��.c�\�೷���k�)�&+X`�`�Ĉ�6\��ۏ�ªr�㹼NT��;t�۫�J�߾�ԥm3"#@�����p��AK:�<�d:�,[u�����^%����$�׉��A�'FZ��C�WS�{]����1@)D=���f��l��k��<�.2��E��&� F�7T2�]7�+mW�^��x~��-�{ �98)��%.W�M����xṯ�z�5��i��N�\V��N��ق3a��/\�b��0e�72�����V��%��B�g���b�U`���k9�Kc��CEp��������H�<�����O=���@xWq��O����W�Ao�e�Q��7?=�Ϲ�hQ$l�wu.ta�}�}�ZЮ�=C���Pu����R덦 �D�:̪Tل74�woMJ@hp��ey���e�y��~2.���q����U��DW�}�{q����x����C� �]�Z�SMyz>?v�:r�j?.�&�2:�iQ%�E�R����)�j�/�����w��L�豢�m\1B��^@��(�S �'��<	j�sM�VlC�W�]z��n˶uP@թ�M"�t���ʕ���VX[/^!L�����t1�x<�Z� �=)D+sd�����;���n�z1�l[�8�)�{u(�xoQ�ޥi뮀�)d��躝e����ڥQ�]z�o6S|gc�Ԯ��o.9�#�!�^��Puh�͛.�ijN�g8���1�nT�kD�˭nC�!�i�F�jM�����0�ry�#nl!j�_��8�ϛ��{<��uiq�as21�5��o���af�>��F�ˠ��U�1V�����o����Y�ƴa:A$y����f�g������G�)�QA��9Qq�D#ڐ�Qt:�/�
��uR:�;���l2n���'�m���@��Z"ٌS�`ڪ�S&L.7O�!m1WR���+K�:�$�;��ig(�~pӨ"�KdɸM�؜c��b�|�����N�՟���s�3�O�&g���r7���[�^��݂�xPܸyԌ�t4�Φ���Z�Un�ecN��d`���E)�b����V��}����-�`�qZo�y�o����uֵ�o��r�+���8}��
ƍn���刪.�Z����Ń����s�t��s���kn���k�����r+��yi�ƭ����TY�n��e�U������F뀁����!.կz�����.QR�ʍ͹f�Yr��7W�tح��A�۔�S��}�{}'��Qy�k��E֢����-A��=�Y�a�yV�[-d[/��V9n����LtK"���Jtl̵#�S��&ŧ�Z:^��w7q9SS�d@�N��T�c_����
w#/<L�*��\p��W�*��J��(�C�}2��;{�3+ E�C��!���^\%q£���"-mJ�0���v{���ʾ0g������h3nt��fB�'I�.���qu�\)x�?s@��b�i	S��}wp�]e����${x�`�j�UGg~���;Pڸ}�Z��7!�������z��-S7$Ӄ:�8�S0�L�y�ՎEQb�@�0��go�s�=f���6Й�{��5��^�<\���UJ�g˸�K�h��G�9u���\w��5�5á��{�r�U ��-��2��bk����� +��VT
�l�f���nW�އ7����we�s)jUB�q9���s���n�s�����K����<H��=�-��j���i��-�[��s�\�M��0�[E�!��q�����f�˪�8B�	�������E7����ܨ��*0�5�$:=���}ܝ�q��k�F�"��8@������*i���l�E��IZ�j�؊��!����͡TU,B�X����pР����r��33��i��ݿ+��s���p�������Z���
��{KmBS�,��fm��Ŷ"�Np�ii+S�Z7�Z�ҥ�R��]-��Z�gk
{2ͪ���e�U��TKh��5P�g��+�|Pe�������.�lr�-u�@��2\%�BYz�����C̔,w�h�Q���\g:�U��rþ����V� !���jhEs����;�W�,hc1W}�wN��Qb놄l������ݫ�%bBE���C�����z���z�8b��fNuZwP��'�k��;ՠ<X����^�St�i
6��꘎�4��]q�n �Փn�լ�<-�//ܶOS��A@��j�s:��y��e�PU��2D�/7}�/\�7���s�Z]�=cY�����P�2#"T�z�&��W N)�~�RӞاX�3Ʒߔ�fS;�rF�ZK�>������^M/Co�α!���a����_��|���.��W#itkG�P��q;uǰ%�yP�>iq_ ޡ̮�����'��}��ު~�4���	�D��z���C�OS���w��l�}�XpN��@	��0
~t<;��T=��Ƭ�u��6�'�^������s/�x���buKt.�x��l��p���:I��e��B��*J�"�X��.�0+LR�����^o��C	p���^v��
W2�v�?'W.��#8����-_!kl�֐q9O��ko:t-��T���(�%м�n:��稦˧����ea���aq�}$GS�r2�բ�9�"!�l@.ӫ�j����㷶�wN��5i����nj/��J�1�@9���71�+玢u�S47�UE�ā
�pm�1��z;K&�S���+�5�:̃�a	߁C���1��Z��c&�w�W����wtP��b�v�lM�)I�cm	�@�h�$fO�<�GP�?T$�x̰9��c*���"&/p;��F���V�Kp~u���F�>�(� ���"�̨B'��W%Ba���LK�ݩ�Y��3e��df�Ac}C�s_/k�(����R+�R�J�z{$8�AT�_�GQ祩]�Y��^�J@r^ �nd^k����a1¡ͯ_V��T�I9�,��o��ݴ����5�u�wL=1q�ⵜ�T��DmD�����cY�o�9�9��Rpѽr1F���r�69Ծ?T��9q�����\��^�g#\�)s�i�3g�-��'��>�ש�
���Wy�т[��g���}��b��F��{{\��m{��f��W�L�]�Q�Bn��uȏ�J�QL�<�x񮣉���t:�� �y�ۃm��F�#�����̰�N��6�XTF��}I��:8�z�q���,n�f+G�}9D9�9	�ӆM�pr�W)s�:J��py��u�{�-���rX�������Ϭ��9��A<!Tƾ� 9u��
Y��Ns�h��\�<v�~�{�x�d5�з:��8�V0j{_tc[t:��%��F��W�C��Ȭ�c�tF�W���n�nE����_H�xծ���]����3WT��"zҀ!��]SHAL�^g�]J�j�o�=���9������.s,�,h�6�W_%�>����y�C�`��4=�p�_>��i,��_���/ꙎF��ʡR`�k]�Z'(��~ʈN��v7*Y�e��|����KV^.ޠ��fx	0?<���cb��B�R����xn7]��=w�:�gN��~�]��/�LT4���������L��8do�_ry�|�S��z�_���V9(q.:�.bȫ�Ȑ�s�!�$u0�)���e@���/5�e{����.$��҅J�B%ƥ\�f�0E��v��U���L. }��u/�ёq��b��fI��h��^}�����ɓp��9�8�����h:9Q�^5t41&�y��6��|y�ߵA`v2��@b�^�H��~�j�7�o�B͡"��ѵ��ޗ\��`nYR���l��=Sdc*�5�	�剗f������nNg���ý��]�*��K�����q2;"9�
u�0�u�����Jc��+���q1�6�1��-7�B�ډ�w:3>�5ܸn9��#���'j�uOO=	9�Ί��yJ�D��
�BɚdwS�\�	�;p��i=��do�o�}���'~�����`��5�w�:�|<V�\���/\�f`]�X�z'��#FeN���-�f]=��|����%�^�mY��Z�O6�p ߵ�8)����)7��vt�����@71�8�'���s��g�V��1`V���HXyQ}�u�U�8y���j��J���ڵ��=pY�LC�J��F%[G�E��F-L��������β�y�{ޯ/S��\�q] 1Q�8ub��J���ʗu����B%��j���"�;go��L����X%��Rr��P��ΩLE[��;Pڸ}�V�����ovl�Es�UMT��%��`9���a
����"��#p�X�CBZ1od���8v���U��+G�^�L�5�7CT�UJ�0.�uM.��6�i�Y}�����#�]QJ���tޠ�r�s$��U��tR�ʂ��.G��U|[	1�E�P]YΗ�Зx�-I��st�m��K�}���խaj�~��8K�@$9ԇ��L+$�s8L�R��D�l���O���'0�ф(j�V:M=�W�.�g��֤=�$f����_BuR��� !C�
ʁS3��T�7���Al�}�R[�F��Ժ�qL膎9��m�r:��X�C�iq����<	辷��U�OBk�9%/B���:��1��?H��fS�&�+����f�s0F}�A�t9]Vo��jW�k��$W���+�-��B��jLWrvYd�cBb�6@��5Yqv���k��JK���� ȉ�[Q�����a����ouT��s4ܰݎ���!���8ޙ�XF�����U�!W���K:�ʎ�:�٫��(�'��O���:�'B3j�ک��8��#�%�4"��Wύ��C�����2��u-T�p�.b����'�Ftgw�/yP��ꘞϽ����e�/PW�#���
ⲫH�;=����Ϯ���:��
��-��ݘ��q8K8���S��4bƼ��Wr�Yk��S��ݽ����#v\F��N����`Ȗ!��w�W/b�c��x,������G[�{����s�fT�y�">猗��z��U�\옹����6���uZՍ*^$�)��Q��J�)9�u��V�"q��@�ug�����{��"{���>TN"���kU"���^���5�e��i�9M)�Q��Y�3�	��X�x]<LS\�u��K��r�?�r�{�i�O��攊O�����~�u�*�1�."����
*>M/B��]d�nh(��j���zz$Ĵ���!C���u_Ϯ��6�)�|��oP�ew������Td���i�C��)q�v�_����E�:�'���߼����	;�Z�X+O��|{���jP��s���IH�/�AY�{�0������ˇuh���D���Gq w>e��Y�k�SIa܀����l�6�V��6^���4C�19���b�sg��0ySȊk6{3�m���
`�EKuM�
G�{���Z��@#5�n����*OJ֐+a�V���\���Tϸ"t����˃��!
����$�q{�(陵��l��N�ht�2+ [χ�-y���G���uG��o�3^��uz�}���;�M*|��Vil��W��K�f���\a�1ΡɥS�}#M�[[��D=���w:��;[r�>3
{]�+�t,w��ܛ�U:�3�$�d'm*ҔT��T��k��Ah�еs,ܪ�3&r��m��貢��b�eCR�m�Ld��׷��:��d&�ZXo�1H)�'��6:�G�6k�2��"y��lͣ�W*{�(�@�ttXi�_guޜ�t�q��#j�z�i�,a1�0���Y�ΰ�Œ߲9sۅ��|��V��ه�;N3�e	���H�N��d���q�Øψcޑ;ڻT����|�-�d�'�}p�Ī�^�g#\�)o;��5�����ڳn�\�������T9G3�uXf�5�[�O��0\K���^�/8j�d�>��W��~� �l�؜��JݜԺ��1����a0W?�l(W=6��J��wp��c؅h��������ڂo�\���.�`ֶ���T5}j���ɴh�W�C���p$���s�P��0�|W�t��f]��,T�&S����f�.w��z+�x��9�D��M5��^�Dh$IHק_�[�C�85���-w��:�]!������^|6pJ6�T���f��V�X��x�&�p�j��.�c���-T�.�ijN�g8����]y	Y� R��+3��r+����� &
>0 4�3�@<�T[�Z������܆븑G��(����.�5v�rS����h�<��TU��f�k+RZ� ���j��WTά���
��X5.G]���}�	h�3i�p�\�h�ʱ��k1t2e2�k�5ٰ��\N%��"���8��D�٠l��cb.wh�.�6"S��7������J�wfɮ����}r�+p�˒Bn����<$��kb�s��ڥ���)7�/�=�piT��q���+�7���
u�3;��\��BE����.d�g~N�{�N�"؅F�;�(�=c/ffSh�5�ckh"P��.��OnP�^[��I35,���[�b��w)�)u�J�Gm,��F^I��ڗ+w��,*k�Z;�f�-��rV�0��A��.�.Ӌ`ᖟ�sl�Ri��gc��`l��6h���`�6�:�2�������Gr�2,�R&�;o#oR�e����6��b�
."$ꖱI	,�[�3G���;�}��:�)��b�!��n�
��pw#���mwP�t��t��'#r�b-���nH��4(���X@�y�M�L�mN]|���:��V#�@̗wMT�#6���(p�Qv��"<V��v�*\ĨR�q��d5�{UE}��m�vu�H���Ge{O��;����&����&4��{��h����y %��X�<�q�����T�vn��*�I)
1�4Eƺmk�+b+��v��	�#�Z��V�Z^
Ky��ޖ9Rwa��K���剭��.�i�U�;jZs����I*!���A�}�1����3�ڲ]�P�:v�4�g�?l�5/���-<Gs�j��������Eq-�e�S@U��ƶ9�UK��0�r�O���Է][�]FX��J��hu���\(���G�ב��R *�'7�P��3[[�ڿʚ�B��㡎�sl�N֬�S*��L8������	S�kj�=����_pG�D�B��.��y}'wP��j�%�؉��8w#=L���P3�_�oa��X�*�mvYn�#�>�;�	�)�0�f�Y����W��x� ��2΅Q�yQK�6/kEtX���)S��:bQY�t|Q��T(ɛ�5�@�4Ѯ�#��"!�`X`�oe�'�e�cj�=�aĮaR�z5[F�KJa[�������G�4�:�-]���J�!x���=���!�L'i�ᯰ�\%�-X�S�䍴�,o&a�*�̈�d+Z�fM����:�����I�I�B3���1r-���h�'"�2�L��d]u�,�W��_
�e�N�6{�N ���f��,R��N��F�2�<	��R͘n=%;'%�R8�6�K�s��nb�2���pi� �V�Ǎ�vE'.�[Eӵ�ӭ�X�<v	�&��!U�t�Cw�3�0�I:�($��wjn�CoL[&+"���w�����e6(T4]�����Y:M�z��҈�Aׯ��J�¶|��D񵮗:�$�7[|x���8��Kws�ϗ���>��B���	ZQ�zaG�]8y�DWgB#Z<<�N.T<\�Dr8UDFHr.Fg�S6P��-H�Ad@��T�+��"sx�ʸ���S���"�QAV�����E�
��j��@#�(����*�9	lK�UHeE\(��"��+Z��w-�q$"9gJ�T4+��Wu
�'A"*�32O8�DDE���ZdUEU�*��D��"9N�
���J�TAfw;�����m+��C��B)@�$���h�&��q!(��I�TD�\��[���bQA&Dr+�)!�")P�����i$�X����*�Re�j�(0���N�y���L�ZD��gfaTj)BI��
��P����"ٜ��j�"�k��u���2Tè�Z5"���=z��Y�r��}��B�o:����\V,6�K:et^o�~�����{��������<����yw��U>|�ȡ'�97����[.�����< I;|t�����I!�����O�i7y90��n޼K�i�I����0|��/ͧ�U�=�Nl�PԬ�����v����o��M���v�￿x1��ݪ����o���]�=w����~�����<*2o�`��X:�|y�;��<�xI7��þ���ɼ�M� ���^�7�Q�3��0�I(���?~�����9۝�}�'�|v�ߓ~��w�k����7�$��}�����1;��}���{M���L>��;r�}��[��\���_S�<���و���:�d3��Pǭ�������{w!�)��僝��s��|�I�0���?��܄���ﱿ!�χn~}��~O.'|>�w��HN��W͂M;���yC�k�������p}���}0>��6����
w���_w�?On��ӷ�����۹\�o�}|����޽�xw���8�y��<�}q���\yw����=���e?'!���ۿ[.�ϴ�>~���'o��������" �"3��PME��ѥ���E �9�C���zC�a���=��]�� |HO�oo;Ӵ�����nߓ�_�97�'۷���bw�k�Ϟ|�������~~��|$�ϯ��&�1����O�O�W�9湡�@G�O?��q�?�z@�������]���'����IɅ]��Ϸ����<'&_����|(>��n�[����N��y�������q|��o��q�}"q/�=���ؽ����p��!H��x��.һw�w����O���='�<��F����|Cù�|�w����n��:?�'�®��&���������M��(Rp/�H`o(+��ע���/���!���>��i���e��w�z߿x�ݼ���{�?v>;˽�N={���y����WoG߼xM��&�B�����<��7�Γ��<&}w���O.<��9�k1��J�5�Z��Kq�Mm�=����?����l�w��� I;~>|��yw��܁>�}�)�!*~v������}G�z>������;y�������^w�k߯� �O/�o�ʞ���&��/.�W��()���O?~/5ƛX6�:4��M��g0E����W�\kjw�kԍ�o(���P׆�1i�/)h���ӬZɝ�Ά/{4�3D�r7H��*�Kf+ڲ1�{{$�^����loR#\8���_E�M@��M"���y�w3��h���Ȯ����I�*�Ig�E3A!�~�1T~��B>��O��[Oĝ��ۜ�7�>��)��x>x��w'���'���m�<��~q��?�?�=���z��}���8�~�f ��
��� G���M��U�%߿��{��������s�����.?�.��y��o���ǎ��7��7���������������7����0����x�\�}�#�o:�����Z/f���P_��Ǥ���p{BM�	'ϼocxC���z�x@����G�� }I<'&��q�!�|M_����yw�i�}N����~t�nӿ}�1>?|��#�e��/�n2=v��HI��M�?}����ɽ����~O)�ߗ�i�Ǉ}NM���H
(|O��L?-�I믯��P$��u�;þ���oG��xM�	��׬y�yH�@F#��k�)_�z}V���.������8�߻{O)����8��< rO�o�����r�?u�	}�N��a���6��������j���>u`\�}��0ї<��ԅU0u��>�)2���ʗ=�����;�|q������<�<�>�7�㏈s�޷{�L���}?x��yw�k����	;�>�]�>�o	��÷=�1>w��zv�~~��~�G�}� }@#�>�:_�O�T�o:�{�����#��gۏ������~+;��y=�pI�0��~���ߜ}Np}߼w���~BO_�p=���'?S���y@�IĞw�ݼ��� y`Ϧ"�}BG�|�Y���*E�s����>���ې��׫��Ǉyv��ǝq�v�����[}K巷s�����]���C����N������ü'&�Ϝ}q�=8�~NC���������~�@���B@_<J�	�oE��/9����|&�	$���cۼ��nq�<��SxBw�=�7�$������v���;��c�xO���w��(R};{=���aM�	���獽'��ރ�}�$����]>���y�1�����^�<;۵[O����	���'ߝ��S��{�N��㝼������;�}q�/|M�90�'�n}��8�lw�$��?�z?��ԝ��:���A_Y��U�\�@�3ȷn�:�vD�cU�Uo��~*�*����5(�]H�K���[$�x�0��u[2a�,�Շ��'�o%>��p_}��L��U��:H�!ڸd��p�������2��QcGD�7N#Y�z��]��`�.��������//�k5Q��|���@���DX�6���]���]������}�v��+������U��s�Ǆ�����w�q�܇�rz��'��﯇{w�~q�9�åq�	7�/�|�Ϗ��ڌ�nyo%��gh�}�}�"DzϷo(�8��xğn܁����(I��`��x7�<��5����[yw�i��������Ν�ǭ��P$��۹|��x��7;��y����q��]�����53Y��w�g��(��P���H�"�h��Nq������9]�P��?��[{<|��yw��7 I{|vߝ���ۓ����yM�	S�{7��ǔސ�<��1�ە�ݯ��i�<;{y����}>ub�����wd��DAF����@�M��O�ӷ��q�����o���xC�F�~v�oߎ�I0��w��S}���|���?8�[�HG�����?`�#�">��_zO�fG��k���P��|E��x����De����~�y@�����Gx��n@��g�cG�U�>��?1YY�C���/g�~��KNV�{Fc��:�6/kob��U�}<O
U[ݍh�>4/����1𶗡�ϐ�L�c7�Q��zz�Y��f?R�Q����>���	��,K���_���C���V)���dTp/�Ze���w�ѽ��:�p�(ł�'���߼���Uݹ�'���ˉ����:��n�.P�# �H�����=��)��I��܌�wV�Ȁ�D���	W"*�G:4�[�����X@���P G#�@��j��w
��,L>�=�Y~�4fy��sC�EJ��͎y[�Z���t�)����vz��2�J���We_d�r��DrLS*���)ѹ��y���1~�/=ֲ>.b�z���L��=�_�7n-,�u��'�N]#����F�]�;�q��g�1�n:��n 7��}aݛ]\=4l��h�#�:�"�UCӃ�?w;���e�c"s��O�o%%��9>����}^�����F�f�6�����'AL4�ˇ�k#����ו֚�VP��v���TwQ:���Q�Jt�Ԧ�Ѿ��/�Qj�k(W����Rs��Qĝ��iW(�urn0��ܰ4�Fhm�\a�<��'��t��w�V����G�ݢ/����>�}Y�C�t}�0d�w��NF���,P�P��]6�a߆筷~`����ĩ�8O|�Y�w����x,M|�tװS��,��'�j$m'Q��\;�:�'��%�f5`Vh����/��#� ��z��Ok������|��Vx�鹪��ݣسT�N&��(P�Vf��0F�P��(U\��,���A:�d�J���R]��jy���u�zL�'������]#B,����(��D�,@�s� ���mU���ʞ����]��\��](�;��ݯ�=���ˈ|A���5�w)K|���Ҕg�[�[�W+j�\�֨�Jq�u�ȱI�J�����0l��b;��Gr���f���.��ֺBA�Wuϫ�5� �m�;��o(6�ĥ҆��A-t�j;72����]M�7�u]�4�QI�J��Mї�Hܔ���yY�E�1���������觔PS�l@�����`�bL�:��[9;�b�Y�� r��Y�C�L��=`t�F��@I��S#�W�P�~V�w�s�e���|ڸb�L�/ l��]^LmF��_c�{���ح G������zr��Ҩ���)A��Z�#�ԝ*�q�+��v�@]�e�bVE�잠$~�i��A�� �;<��<�[4ߕ.���xlr�F�Q��xL�}*%PZK���x�
�?Ss�Y&W@�0V���vdE��S6(�*��7�-Υv-b��3F'[u�\:ǐ�psʈ��D#ڐ�C�A��ꬪ�]SN�e���$���L=s���p/�h�1	ݰmUc������ڻ_��$��;���?5�v��zkX��7����L�)�Z���*:~�'�Óc�T#��@[�j�}5f�����>�v���
�5\�7͑Nq��*����:�5x5^���0�W�ΖE�@��6(�U��I�V�
�7r��O\Q'}n�W�T����I?�=}x�h�g����!�>W�{�v�ed��k��/��[E���)�YY����IoG�6	�c�
�M�����hW����E ����k .;77S'Wc��tJ�)d��Wː����QYr����-#l�]����6r�G���I�:׀(�w���i���.o�1�}��H+�#^Я�X����L!|�M$�8��ޗ�ʒ�*x�'��{���o��N�~Ł'��Ց�-�k;�`~��QHѹ>��X���y��$ ��sX'�c���cn�鎧������Rb��{0��=�r��F�����r��2��[߄��M�y��*��,:1x�G�1*�<2-mJ1�+׏`�
1���5p���<2I]1(���1���Lt�Y�P���ߢ�_�3�y ���:Msz���"�>��h]b0P��GӗYB�>ڬ�`�����Buj��I��E%:�]�ow�p6�ll��i��Br��e@��iWI('��؜n�׆
����x>%{V���B�1J �������χmJ60Dr�1�$��(�H�T��هw��>�����|��]Qϩ�1pVR���Cق1�NBuR��[������|!ڹ��p>��bx\C�%�:;��g��+��w��絰j�b��;X�n�uú�P�$�+�Ե;t����A��+�(����L����IW��+(EV�uԗ�~ v_id�����i�ذQ7{X(z�/���6�{r㋜�x�=��#���U�)�:�p�}ܕ�n̫@V���7x�wW;��q��"��Zb��,)!����|���">�"#;#9sn�+�#��`�nP��_��0��h�c�	��%c5�T'X�Io_d���aC�T����Ş�(FkCa�BD!�b�f��p̘}��g�F��ֺ�k`Vgoi9݄ue8��=]����,)Vv*����	Ю�g�޼�H���^ ��]*\K�{�]@tˌ�@l������k>�~����tP��(X�N�L�i2!�R�����T�z먥A���;-���2��}93=8����;�%�Jʺ׫"�nOއ�p��!��3Y[\!��r0��T��C�P�\w΀8b��㻅B!OF<���t���I��0�� #ԅP���P���D�3m�1���3f0�ј�U7c/�n�r��TW�_ܕ�� �g��.%���N@��z��)<3s��1�����b���%�^,/����kՇ,����d.G�ю��U j��~��XH���r-v�T��˔�u��b���kn�婂A���˅��
�u� ӆ��]��L��@�;���J��!�4���^n+�XJf,>��S�� ���,s�btr��%�YOi����u�o%���`���Tt+���#̴������ٗ�V�aE.�u���MͱW�ct�l��)Jy
��=[3���꯾�����xӂ�#�o3P��-�:����z�Oir�w�4��c��:�>�Bv���特�uә���(�C�qs,ECSz�
�U��tOe�U�]���)�)���(�#5��5�GU^�޶q$�pDhZ_�e��E��BQ�:���C�":���i��
�*��]�3o���x�z��4��H{P*�G��G-����w
��c>6^���4T<uK}�;��
.��P���i>�$U0
� �bvC��}��Z���B*6�KY�ڷ�k 8O�=��W�N깧�n�m��('A'����Pu�D ����:\P�����+Vi�%\K`�5�"0	�:��땿3uQ������G��3^��r�"p.�
�;ڭO9J��Q"+�����A�;�健�#448�#�C�_*���h7k��f�3�u��]��ci�b�{������yGr�^� ��~�a #uC/]7pX�c�FNX�bڷXK&׽�����,��������	�K{~��5���}�/�p��s/v�L��Vi�d�6�ͨH�}Hu`�i�׺Ⱥ�Քt������ga�Razǹ3\��]��BeX�>��iڼ�TbDif1���o�}�GZ�n奬��ӑh:7���ӈ�Ij�k�G��y(��ۥ3�:�|���e����ǅ@��qR]����_W�F�I\�KY8f�LW�S l��N3�ĩ�r�%���UX>���Z�,|���;�N/>g}Vc��{���pw��*�5u4u�ʁ�>�jU��FԺ�ɻ�i�A��\��=�Z�&V@q.�8�~y��gֺ�d����zT���ٗ~o�� �l�7":�67 h�}��e�*l��uc��u��{���ǈ8��P:�"�3K2w�ۍY�m�>\��"�dF����ת���T��&ӂ�#�l��s��9�Ew�엄���y�C�"/+��[��p�N�o�"���n*�k���Rˣ�4CM��-L�/3ȑV8�o���U1g߲y�C�`
���U�ҩ��Z�0[Z�#�IҪ_^�S0:�h�c���P0�/��G\ʖmh�9��c O39 �1_[�Z������0�����:nΜ��?��q/]D��J~~@�u���'K](��k�ızlƻ�N���0�jJ6 �־�1N�3F'[u�[�y!���$q���Һ��X�0yB���~�,�z��j�z���w^�^?d��TK����m�L@�W�YR��^J�J+�ϯ� 65�.6������G������֓�M̾c�;$F;n��b)(�䝸�8U��ok�I�&e��z��w���ӳ�
�z�y>�T�����N?������_'e�n��ӕ������U�Pɯ�u�������1�L'v���V:���Ʌ�GZ����h��R��1j�U�[�Y���_��_�l�C�x�n��`Oex��	��b�	��w��t�H���ښ:)��?9���)j�+UΫ7͑N���x��f�烮��{��bC#��*ע�B�^��;p>�A�Â�)N3Xʌ����u>����SR���!6�Tl� Co*X]=ըw��q��?=|�ՂEsF��U��E���a" $��F���yy5��W꫘p������6�!����&ս��36��\ᘾTY�%��6	�v���[�o9�'��}���`tt�ͷ���s��q�+h��S�U��$zakM+PxA�[�{�z����V��1ư�E ;��#~�LC�x�Gjr�����ƾѕ;&��p���s���rX2�Pe��*�|���c��UzP,ȨI�em<��m�h ��v��ޡv�pK��˹��`�\Q�������U�3�_���(��M#r�ڬ�p����l�ɽ��"��ɫ+�V���$����"5�>,hg�A���}�]�yw���DQmv�gB!{�r&�j�^w;7[b���@� �N����l���!n�F�}0����+k']b�f+±�S79mʁl���tP��bw�bU�-Yk��Bj����~�c���tvi������q��qs����&�G��N�ȼכU�J��ճ^���!�>;�&��j�J�ҋ��}�2�x��x$���n��7��{�J�H<8�G�����4|����u�C�F�PX.^M(�2�r,۫7ê��*$�K��W�iTvݮЧ+��s��QW&3j���9u뉀�R�]�[˓	f��VS4j���H�QW��v��\�fQv�IbG�vsqZ6)�T���E^m5{5��=Lt:���jTU�������F�;C��!m�]r�u^)��������Ю��ކ;�vh�²�Gh���/��0娥ZM�E����{�q��k�W$.�K-�	�&�!ʸB�X��|2��i�j�֛6�=�.�K�h�*oabL��s�1�W��j	�U')��*���z
j��Cɹu��%�ݚ f�� 5J�w/ �!O.�=����A��� �;�m��ִ��C�������#<�k�i�`^���͠���Wϭ#G�`A��y��h��[n*Nn�6s,-�q�i�Z�ʛS;j�k :eSwG��(�����*V�qp�;,��ߝ&��\qI�ڶ�LȮ�o�͵ G l�;���d��q1�v~��&�Dx
�wW(wc)�qu�y�����H���W&�Rg-����ns��1	o��\ݽ�RU٥�����N�/iյY����WZ�%\��b� e��V�kuϿ���x��z�G�v�F�A�@鼻��ŝ�\�����D"̹����b-,0������,����٬/90E�u�@+j�L�kn�c�!�}����ױV�q�1�C,/�]@e�Kx L�H7��v�B�7}��KO����B�X���Q�.�GU%��\n�È�Sbԗ@ɹ%R!��D]^�ߠ�h���q�"yay��bP�+,�h�]�o��ܱ�@���׶:��ek��W9���2�`Hr�sa��x3��;o,���t�"Yq��]���XVnAS}����}�x�`n�5v�(���k�g;.�g���:ɑ��Y�l��3��Wr�ԣu�R�D��6����!�WNo</��b�,�H�K/+<��M��scT�ɦ�ײ��O���IX};�n�+a����ԸřȨFfiY�	���`!�}�b�kcu��"�.ա����/H�K�Xqۧ����W���i�d�l��y
ó���nІ��/z�1��(f�B�)jQL1��l��-1%4�I0���U�r��jFZ �Ԣ�T�kR�H�D#�Q&J&�Z��r�$�E����,�f\�D*�����M���$Q�UG*"�'��p��,�QTˑI�ZW*/K���TˁQ�j�TS�"�e\��\�(��"
�sԐ���
#��9QE®\��US(,�%Bu"(��r"�BU�;=����I���"�s�A�\�(���*$�����

"*"�\�TTUˆaQÕ9�bp�DT��Gtw(,�*dW����$��$U�+�3�9p�֮�\�*��B��B�z,��T�p��9�2�*�?A?H E�92@��Xbǖ��Wox _ډ�[���R��3
��H�b���3q��������]�;�@,���LE��W�}UU���j��@�ƿ|�n;�
�G돴��*�$�* ����4�����n�㡊[�p���T�3=��P��1<�[�,�1��ߓ�p�mJ60Dr�1�&
����P��ҟJj/�z�HB誔R������Do{0FS�M'UT�V� !_�,�ݼ��Ir���Dg��.1�E�~y�l@נ�Ŧ�n�o;�5
bIAU��bn��=G7��۩�̖H`=?I-�X�Y�aR]ms1����2V3Z�d�$�#	��ݯt
+,{������	�a�1"�!�b��j3d�G�Ԙ��N�.���x��V�ؤ/���l�U�
�v�h����\�dl)�h.�0�^�Dp��_0��e�o��*�{ʗ+5}!�΁�4���F~�O�T
��Y�Qe�@���};9�B�uÒ4k�������:+;��^s�̆$9�lȉ���k�f:�� ��7�,Gz{�!��3�~�#�������_U��=�@�:1�1=���^�{.�^�����b�ɻU�ꃩIKuX�R:D�J�����v$���7d���u�<��o�7���&h����^����bo �*on+�c���B��sl�"e�Z8��%���]Fn��Z��n���]�=`}��rB��6�L�x�q���Y�+���˘7|��B��}_W��h����H��8:�*���y����{P�'�� �l�uLGf���Q�k�Y�i�s�t�1m
X*_�5��9�N���,7\ϵ�\K?�9�<�3�ݺn_'�6朗��0V��.i��Z68`���b�P�]<LS��p22�ڝW{����@P��{�Q���<~(�t�u��b���kn��Z�"��=(I/�Ґ!d���6����0��U�^����j�^uW���5U��ڗ[��X�*�>iu���;��+jb�^V��-~��^3�gG#�2�-SCb��c_I
{��d������*�S S&�'����k��%��8�X�~5�E3�s�_Ƒ�7���C�":�x�F\;�EvLf:�\�mi����5sR$C�8����ځ@�3��Q���+H��/ND71��;�R��?r�]�{�����m�Ǘ6Y�ā
���A�0��(p����| ��Ǆ8�y*ʿd�"��cg��޳��3��M��Qm�U��i�限�@d�%
,?>�U�|} c��8��9����^����-�«�N���>[����W�����Һ�KL���i�H�w{@Q[��>2��Wo tE�f���8sV{V�y*���B�2%8�%v�-�x�>
��#W�XPN�ω�Q���������̨R�IF�<���'<K`�5H`8M�~|����4}F�Ѡb� �y�,t�(a���I\���RڗXWo�>��aH�0����.0��uMB��}�UH�T�O!t������e�@Öz��&:�H*TUy�b�609�q�7o~3,���gI�:i[ي7K$q�M1�V�L�5~�G����t�Z��r*������9�o�Osir�5
̺��[�c�
��Ua�N�Q��TT0���3��|`��f{]u�%���9]��k�1�����I����7/�*���G2��_�f�4*�b|�Q��֓�����>������4yذ�]AĪ�f���Ns��z�]#�f0��]|ohu4u���%o�,� �\2s���/[� ���*�g"�6ad��mG�i�]���6`�$�j4u�a��:��,O�����`���]z���%���@LF4�0���Z�K��p��ҡ��̷��[����o��&`g�z�B
t�	��Q��Ɍ���n�׮.�u�x$�K�|s>�!�Q]�g|��mK�*�YNQ1�m�5n�Wٻ��=��[%k��z-����,�=PA�ܨ�^��%#��J]���.�$�K��xR�M%3��г�5O�ל%of��GW*Axe��x�R��L�-�>Y���jU��8A۫)H�.]�}�}�G�f ����O����o媤_�H��jiLI1��Q�����ֻH�
��f5+�#��}�xӈ=�쨎uC��,��D����`�w�����௭�y���t�ܭ�7}��ު���ics�븛z�'���?T70��`5d��zcA�}��@�a;F�����k���C�� c�up�S���C1�	m� ���(2$!\�h�!i-]�$λSv������<�{N�	���	�Q�PɨI���hԻ?Wy�X|��41��[�~J;�f��M!v��_s �\j��T�qtT'���ڂ+�S&M��x�hc�%���:P���a����@�۱��m���{�Zu`U���Y�l�s��sͥ{�Ng�P��MX�}m�sF� b���hzeZ<�L8�5���2��h���TsoY�ܖ.�<�G%@l�6��7�6�g������>ڹv#^Я�X�����O���r�<�=�VB(���<�y1GK�?b�9���37��W����J��x�W�{��#�b	B����2��ɢ/�Ѕ���XYW9�3ٜWu����p1q.mT�މȘ�$K��,gձ�|�z�W���Lզ�j�iN��뱙9	X�f�m���E��j.u�u��i��K���P�39�:i֐鹦�$5��݈:�fIv��D��n�����f�r��(�='x�q0�"���P���C�o)���VǕ�bҝ���o��>{�(�w�ds#��SbuKO}��ꂀ��ǔ�T�1a�c7!��#&�:7��#�gU��s�g��sZ��X2�������xGY�2s��v��UE�����]ݴ�����"Y�j�ρ�"um����`�j�yUz��LemB�cPP⥞��R� �{�l-�zuy�5r�����\�������\l
lq�۷�Xc9��D��)���Eɯ/tn��E¹C�0�������N���R��E�F��j7s*㺕��ܵ�s�8��s�T���ۑ��x�S�SP��P�G$��"��
R4��qsn�+�p1Čl�Ko)q{��k!��M���x��݊���:'�Շ��D�oX����<�ׁ͇wcԋ���q��V����#X]ږ�{�߹ݺ���,0t
���#���7%&�G��\7�h�f��ңf���HW�{�*,&��(H�S���`o{���=�'����uJٛN��B?f��>�c�5Ś�ݥ��(���g,����V�
���>��{��́�M#ﲘ�S{^3��՚uK��G`K���`k����Bf��DD}��wHPﹻ�:�~ң]��-������/��@[�Jy5���e��G�ѢN��i�Q�-�P�C�mƻFr��ȟ��-P}�i���ԇ���5�>Z���Ybwi=��nj��9�6�l��U�	��p@��tn�/7��y{<�f��{*�)�x���5��垿޽�zٷ7,v��l^�T�n�*B��W�e�&���g��2�yM�.�en�QPf��JSj�l݅�%�^_�8?:��3��3s|���j���/����y��Y�F:o��mٕ��������X��'P�;a�s��J�Ny��`�gN��O� �Ѧ� &�r���YԚ�뤈Tk��R_K��Zv��r:��M�k��0Oc���Z}pVr�8|�!Q詺02�vl#7|�{�$s3\��>[�T�]|���!�{_<�^7cp�⣹m^΁0{k���r�V�:���ܐ�Z+k�֬Rr�6�Pf?�잹dk����[
��Qg����Ϙ�
���b��n��׽��5W,��v��t\�z.qZRWY�v����ǺJ�L���ݑ�8٭m�:�Fd�s�$&��U��\�,u�	$&3_���G�2��[oV���0*�<��-�K��ֻ���99y�Fxɮ�D_N�z���\
뤟�8�Y7��[�E�t�w\#��v=�!1=m]���m�T�Z�?�R�*B�!����'V���/01[G���冯B��R��E�w�3�6��=K�$�x�����2�Ϲ�5{�%v��������j|��օ�{�;ٯ0y�P%b�<�E�W����t��̜w�}��}��j�0jq��ô�F���j&��|��K�j��:F	=W˕�Q���Ю_L���ޯ
��m79�0�J�D�t�ms�"�����:��g�d6w���6ky��Mz��;]]}��:~�e\AF���u��:�7'"������>~�:���W:���fsy$�د�mE��R�=��y6���g#g3�Lq�)��� �CP�z� jڼ�%{�	T����Q.��G)���G�ڡHb��s,nY��5͋f�Sړ������T/%vR��mٵ�I0�uvVU�W
������̀�)v=��nvC�Ɋ��z�6k]��U+�u�EHJ7*5��������9
�$�kf��']A�����&���E��EXpR.}��=�گFܧ 4狧�Pn?��Y��Ϳ��Q�l��D%7��*�pn�οzB�,ծ�����FS0A�Zj��Fr�Nt��b�D�Υ*I'�#Ό�.q��T��U�jg�Z<�<v͠��g8��v��k�m�K8�Pz�?�}'��Ur�I����NE
Q_U+v�+g58�c:�����/~X#��D��f�-����N�=�M�<r��E�i\�8�r�ڈuJi�`��GB���,?�=��R�譄+�޷��Ty�3�y��ҙ*��h9N[��^�nvℷ5+��2)i\���ݬ�$�;��a�#��10DȺ�ꚧ�O:��0lL�f��W�����9��̪Mi�LMƵq�l��S��$S����,՝=nw{��Q_��ݿo�X�P&o5�!n�P}5�ՄJN���H�Ӛ�p^2�����H�pQ����6p�ﷹ0
"��ژ:Ѯn�T��FgD���;�!4]4����lǬ���9b�.��z�+7������J���i�����+�����Q4_\��<sh�FN��h^��hf�K�s{��ʎ7�s���>�`�;/�n��Y;Y�/��8�a�����;����8Jwo�ġ���3���w�z����v�3k;�ͦt��%���n��z��Q��<��?/r�x.��[U=�9��t���+tob;~���w~�:��u}�޼�Ӫ/�;}��1�κ�O<����s�8z�qÚ�ʀyTM�Wҡ�F(����.
i��������Lt�y�<��W��js+�{���d���є�xƙJ���$gTJ�[-�%j�*�Yy��ke���
����ё�^�t̂�S�>����%��:�և���Vr���U�!�Ǡ��UR�S(.}��]�.��ow�Z�3��Ԟ_��އ��T'M��[���@2Ь��-}T	��P6���k��Q�Z���;��hA��
\�� ��lr�x%H�ʕ�8Bh=Gm��HNlQ+���z���b�s��I�I�Y�3�u�vU�u(�t����̞��^��6�����q�M'ȹg_s�O��cB?��������ƒÿj��Z۪j�.��}���x�WΩM'%��SY۹}KUQ����o1vm�f�"~�C��Rޗ���k>gpWͳ�^�A	�2'x��������D[ޢ��#�Zg��\����xv��E�t!�����ig:�c^2p��F�S�K5�%u���-sR�&��кk5�K��s�'���r6��/�k��\k�r'����ճė��s
w"�f7sS��T����Vn�WՏ{��v8sPۍw�S�?s�Z��V��q���K������E�Ē�K0ʸ�u���(��k�e>�z&ݎ�[�UXٽ�I��M�p#jʱ{���/*;�k���߽Xb�޷3�*z�}���T0��ٵr*�z~�9}E���/���R�R����ʬ����F̨�_�_W�o�zwo���s6s"Tz:ΣW�:��{����`1�OP�'�b�{�� ��GSܰ8+j#���ǐ[lF5���Z����Υ}�`R�F�uLݲ�J���Y�Q�;Y,�[�̠�T���ٸ]a���Q:�TWK���G]����59���:y��O�>[����vod+����$,%Z�e1;e]�6gv�(�}�U,��i�U�<��k]>ǎ�]u	6�_wS�9yފv��v��r�8��F���fzD&S��;VV�99��;�]���G���4{gJ��0�d:����\nM7S��摴5��K0�����*�nҲw/���v��E��s����;���Q�F�f}��"�u��˒��%�owI�0�:�RA�j�l�7��M���c��ةAyz'r[a]�`�i�5$�[���%Kta��#���_ q
�|h
X��*5Gu&��u)�����2�J�޺6���i����L��ЖX2Z��Sq�4�����Lt�=����̣�;QP��g^�6Y�]�v �Zd4ӫ�v����⣡g:s����h�[Zz	���;k�nH͚��Op�I*JT��:?�!��h�}VD�w9v H<�G����J��gTe����pJ�a�_��Kon}�ggT,�h-��HbF�s
��Hu,J8cM�{��
�-ۼ"���C��/$Xؽ'.��Gw������Uw�:���$�7�k�;Ն��� F��u�4{���o�{���]N�i�ƭ�Z�vK�J��Oo/�#A��i�"�J�Ca�0���1e6���/܂�k��4�#Ӯ�G�B�����N���u�2	�Ѿ����ޔ&ծv7�� �T`�y��M�\�2ŬH�Ж��!p� ���j1.�ݔ ���lڨ٩�u�b�a뱸�T�:�nA���6*D�Gkz�sp]�]%��J�k�0W�����kܮĳ�J���x��N�Q�ώ"ˆ�	�{���ݐc;ʐ��Y��'X�p�.ȉʘ[U5N��`��ڳS�u����%�b���$/'[�oGv�4�Wy��mFMb�X{+Mz����ȕ�p��hY�6��ۘM`
P�X�Ε�r�k���k�r��Di˹���4L�)�z��C�,�L�8͵�a���:�0�^��K�IQ!J��U|�����9��8�f��&%ѐ;�W,�M�*���(S�ݰ���|�n�tcpw�O5Ce y��zH��^���"�����VK��ڗȶ���p\{��pI�P2�QK�����8:�<Y%_$%<J����Q�0�wZ��L&lǬ�Kg&�
n;m���6�i��pv$&�	����Z�wU����q�O�rr}�M��Ӎp�BK��u=���4�n��J�%B���GJJ�N%�[�K�w&V5�t��i:c�y��e�c�
Ίf�r�)���s�村��e�}��{���hH�)��ȇ��u
/CA\����E�6QG��y�S�O2.Au��AR�r�M(֜(�"*��2�*k<���s��� �9Qp�r9���
�U78�W*��B*��(�DQ(�m'';��0�J�I�W4Î�r�$&s���(.�F��"�ki�U�):Qr9p�J"+�QTQTU7$�]�"(���IӜ�9��9�p���@�U2��1������] �:E6���r� N'eU%�N�jP\�U�ĩ�`EY�QD�̢>'�X@ B"n��9˝��X�J}��|Rh����A�[���l�Y��
�Ue�a�wn^)hpո�[҆)j�a�O�������S���S�*T~�/�����C}��OJ�ܢ��V7ʋ:�=]����E��d�d�6�ey���g�τ/g���l���וaʺ۵'�b�[��+�G)���X;�OGb)ͽO�Z|��8&�Y�l�̺7�obAް�<��p�'�%:�J�tyW�U�-e�|(y�o��[��"72�c$"I�O�Q��I���� ����U\�p9��s~���?y�r哄BJ��$���Y^����0���ʢq"~����[����FD��&zmC���������v�S�*B��!��G�ծo���0�8�p-;IBǩ(�=�y�����*{m�)�<I]�6��-��i��/wta˧�c4)��j|��]���1�m�GL���]�uZ-t���,Ŭ��ud�زc���Q|�-��Ќ�Dk��E,�� 5l�f�o\&rm==«|��ub�ih�Z�o:�)�ON�M�f�1^��Yj��R5.���d�b4�|h�\+�ɇN,��#9�,��l]K�}�'jm�Dm��ʧD�����s�\yhݜ1�x+p�Y��N]Q͵K�}U_}�O�kўɟ���c_b$x�Q�lҽ��^��U��,3Ob�q��{�n�Ǯ�z�6��֗��d�d6K�9�[�,���.Ȱ/^
�	��i�M���9������q��X��ޟ���_�Q���Ͻo��x�};�^S��-{�0�����<}��Y�O8_z	3��f��,�.��s{WY�y(����j7e�V�I6������^V�u�bΞy5��_[�T�p�ct�(=˙��4�uy�)�}:w�A������D��s�5e�7��Jsh�=2�S0A�'���OJ��Kz��r7���K'}��A��r2?�zu�3�g���z*x��f�l��]c���:���S���Z��UQ�p*�h��npGsn����;�]ȹ���j��gS�9I�w��.�����N��)���1����ɟ�Gw�t�˔�Իr�&��W����K��o 0zS�,��3:%�nƈ�l��P�/�݁�w��k��W�r��{Tq�Ҭ�xBw��	�+ɬ��XT͚�������31+.+Wr�A,�}����[�PI=I��v�:Wu������v��)��:����j��3�r���m�ޅñ8m}�f;���S�k�G5�gpT6�*۝��	O}6'ʷ9���/��]A��g����9�
~��k�C8øG#��5�쬝�7=Ǵ�G�]�ԗ���mg�ͣQ���5�~nz�uˆ�9Ax��+u��G��a������;�j���^+�|{��r�]�ҥ�x�;۬�&G8o�!$�>~ô�F��í��������S�Nx/$���\6d�~�
��i�u7�����?x����v������W����YF2߲D7E��ï ���]�v��z�\�<8_���|��������r��������tzuE�J�p�����V�q����e�m�yDl��Ø�+2#F�T>��Q��������H(�S��}W��!��+��%k��ym쓱��g��j�as+���͊	q���gZ��^�g��9�a�}�鬦�7~��H��z��o /�$��b���а���b��$4�oqu.y����+lS�rU�ܦb"�MY�ˠ�ǯ�.��D}����r���{�F6����$�ս�Tdy�2�eX�3�|��VV?c��w�����>���zS��J�^������j{����Z�75���78�6�=��OB�]ps���e�s�T��g��'���.Ț�+��y'��k�;9��9̒2������H�^ޫ�U�e�}ᜈKv*��K��GnCc:�3���������;�o�j;Ȑ���}�)���OV�ߨ�c�*`�C����̓ʆ�����y���5莪鯏H�����~��|^Ϋ���s)���ݒ�Ɍ��;ʇ%s�Pǧ86.2!;r���q#���;|�.��gx����W���4֤�䖥
�%���q���lT\5l�L��w -����}2D�>�jJ�vyBV�5����m{ޥ�Fq��v�Շ�.5O(K��0^4M� �׷c
�N�>ˈV
�Y���r�/8�z����u1P�u>�dZ!��n���Y����+wf�(q�.S ǔq;������oe�*��q�[3u��%���b�Jy���mn���+,n��];���F��b��UUW�QtS\���HA�����KČ�ۭ���3Qn�ۆ�y��*_=ܸ�:�v�Ot:@U��/`��&��9�i�q��]�9g��Sf/��eZ�Mq����}����Urr,�w��S�U?g*rS�umP�K��+B�&��
-���g���81�{c��f���Qf/�W�N�嚗���"^�U٧��sXF��	��䝗O5�����VR�� s4x�gt��������j�z��E��&&�ȗo���Ml��$B�C��]F��}�{�$$�}�=����n2�soT�2������<�a�ݍ����7ݩo%��	��0-���}%��Z�c/������=ڂͻ�I-�91������p;
��ξ=�H�Oj�R�ؖ5���21�j�ñ��W@t �k��UM\��,ʌq�Ϸ���jݹ���&��Z����0`�݋�K��.�u��H2�y�%L��ulf2��x�W��WY'�׎��//!g��WETܥ�pK�����\=Xv�G1�c����_T�E�̀���֛�����fC>2�� �Shַy6�)D]��8:�Yկ�_}�Uy��I���P�ކs^������;N��AR1p�?�`��6�[=��Ef@J��A�Թ
ǌ)�k����3�Sob��͙�� �]-4sE{n�p~����]�e,ʸ���Lok4���!�иϓ�*!M���;#3�щl����S�}�$���w&���W����I�Lۍ�����[�0��n���b�W�G�V�7]��9"���T�a]3�=�����v�C��Pݚ��xuJ;������ޔ��b$C}�������׮{B��֥㑪/�����q��`�����b����H�$OV�Ncm딯wDÌW�z{�ƣ\��u�����ݸ..`g'b��e�����x���Q�_ҝ͢뢻^2�p����ɚ~gO���	ZL⼝�W]��������D��P��m�_w.f���Y.�m�]���TH��Eg$<����}w30��r�7PR�%w^�Qr@Tk�6�p�"
sh�T�LoF�T��ہM�s�*��*�ԩۥ3�JF�/,�S�����񩝔LK�ɗ[�e�7Hv`h�.��Sl��)c�;b��!՝� �9��7�rQ�\�$�ﾈ�֠�W�[��3;��C�] �/�Tr�/�F}؊4�^o;����)�t��geY}��ڨ��s���E����Nڦg:�13UƼ�.��=�n6�7���C��OQ���K8����U'���Ӝ�:t�[��������s�z�M�@�.��G�Y��w��U�I�X��j��h����E<gi�)��:X!��{,���M��v��v��8�~٠��^?v��/[P�௛{m��E�y^�_'�g�챪p���q��B�{M[�a9�
b;��I�v�0�
u�sc.?m��̈_� ��K�p��!U⨽�<�i��gɭS6\�^����]��͝@��ظϵ�ĵ~O4y�Zۈ�9��Z�˕��+G�d�|��ZP�no��5��k�T��K��3,�N�9�l^�К3"\�	�3�yrJ�8g��^;���_�7]0V"t�/!�����ۤ�=P��LyA��'��#-�V�2��Z�9lL{R�g%r�A{qZ��*M����J�$���}��s�A��QK�\74����N>���ﵧ�$�z��SG>9�i����պgm�ڎw�q�Aʀ�v�}�P(g(�l�ܲ�_�/��'�ecs:�J����(�Ɲ��â���.�M��8Vp��%��z[�2���^��J��V;���hة���;�K[B�Yu� ����ÛY�w��e4e7���_�L�s�;�]�;x������˲�7p6�I}R�v����f{w�u(�.H��d�|�}����ˈ�-V/J���)u�x��Nz�"�/Q^�ή�W�����{��NP�!��59�qۆY��gci��^TI|���*O.m�^q����$�$x�yY^L�!�yu�f�W��p�qfz)�����z�?��O�aE[���@��Γ��9�A�!eeZ�V�߸�מo�+э�b��y��9�+�s�BR7}��PǓ+i�+p��L��O����O:Cͬ��̖(P�:���D�P#qcW�v:���T��%��Es��Sn�ͼ�91�K9�5��ڷ�BC8v;{�G]:����l��#�=H�]��b�b�$�������=�_g&.�\=�>giU)�������H�w��o�ۗ�*��}�]8�B�F�>+��gL\'NG_L��w -sR�$�0D�v]�7����%Y�q�l��h�Gra�2�]��D�b�9�K��N�k{h��4���ۓ�gؑ�>9G���̯f׽��q�>��y+��u�e)7�7��s`G���҇(�ͪoڸ�W�~^�	)�;��nG�I���X��� ���W'�������9����o�^�f��ي��݋��s��-:�������^��Q�?@�F�dOxf(�z��y4�����ix���%@y{���f��{c�z����1W�XvG5%.�\�mnlTR��n�\i�O5��ƴ�]s����j�3X����'��6�9=���m|ec�잞�����uw��]��aEx�k��aK-v��&j�跎&h��S�:�j,;z�t[Zvw�����*������5gU*�vtɷ����z,�LD&IA��&Ї:2��G��2��<��k���,���6�3-�������hQ(�u�����\� �v�Ͽ�����(��<Te��߫������`����y�zy���^XB�t�5b#+F�R��)��!���_*����C�QNڋ���,ڊ:��������p7i�������}|(5�N��ns�}3��!���~X�����*rs��2����,�G\�o3�n$��ш�P�r6������3�r9�r��uNj
�����q�A7���&�^��avT��s>�}֋���)��Qm�B�sQ2Wp��{��*�eOR�J��g��\[s����I>���鉇��s���{�{�D���T$f�9^�a��U;1���|�=�n5��Wd�5�»�;=K���5�t��f�>�[��N�B�a�y��(ν����U�JE��UY���TL�k���5�=P���sKro�U]us'6ry�ڳ}ie��4��.��J�ĭ��V6rUk�$�@���l�y���Z� Yn�r�yW��ҙF��4k�w(�ܸ�u�J섍�n��k��KlfXF����e׬A�ob�5���F�ˍCq�n��w�1��d˨6BΤ �:֧����]��.�G3Ʊ	َ���II}��Y��j9�%u�DB�w�j�+�8�u���X�ѩ���8��h�qp�lZ�(�WJ&�[;�mk�cJ���	�Z���ɢ��k�wu�ej���i�kU�V�ISL��3�wR{y����O��Ѵ%�,�(1�ЄZ��Yؖ�*��ͼ���k ";��CAM����a�o��t�$�ə�*�}$tM�tqW�ڡ���+��yXهTs�PV�f^"������
�u7
j�:��d�A��g�G]��������N{�^Q�xj%�t6�]9n�М���\ő��`�{�"�y�}��7Xnt�F���sn���s��
=.����]�_l���"u��-Kl��p�� -ڋ8��`����"�l̳Hր�^�����n�E��xv�2>�����p�0c�6�L3��^����B3p�R0�𔢷�P��m��_oD*�U�7�h丫���w�I�3*�v����v����U&���1!r��k6�a��h�;� ��M�z6)�6��X��w���0
��u��P�����7�i	�7-��JMo�-m+�>�%g����������kՕ��5C�SSl��+��x����Z��%Wf%�+i�G*m��j�[f�!@�7�i�u����i¤uu��u݇s�=��)̾ʔj� 诈\�ho�,�:��6�峘�x"X���#C�>�j��v�+!T��uD��+m+��T	f�ǎ�����K2rL�|�pbWTyw�m]7��Cc��{I�.���gT��#2%܆`�����0Z�zːR�ne�x�P���0������C�Q�[H�0�m��T�YJ���1��K��8�i�����;s�M��]z���{�2�^&��p'z�q�GZS�J��X3���1M�]�^�a��bZ�X5;s��T�I���1ڣ�n��AA�e��m���y��y��� \���W��Q����n��#6���Y{u2���;���'��ɷ�����shH�!��Q8�Rcyct�
�蓻sq;w�sf����N9�dw|ӓw��[�|��ۿZ���	]�b��va��خ�Jf�*q�`Ve֫�UGE�W�";R�M-��@Rۨ�c�Ҹ���W�5ݪ�֩rNL��L�u�41��bZ�G�k#F5}��Y�)c���l��r|�Gti�HO^��\p����޻�u^�<8��| �.U�u8�!5o0��,��8���/�%�m�p"9-�F��#��Ę��V�l-���SUY��
��e�+�k
�2#]��\���	%��AϮ1U��P�?�$�J��aTQvPR��)D(9DjEFB_���.]�t ���"��E@rH��9T�����S��
�Qa�uAR��;SUPUU�dt��8A�$ʹvGeʪ�I��QȨ�8QdS/!	�'&P˔I�b���r��˲�v'0�DQ\r�r��l�N�I�t��N�@PQ.Rg.pH���<�m8S
����I@d�����YQ�p���S��2�#�0�A��5B� �T��D�0�N�Ge\��D��N�r��/^<�|�>x����K��	�Ɲ�s��Q�ڎ��9�b}��A���]��}f�W��8aW
�98�����V\=]���U_��78��逺8��Ļ�/w��������T����tL9�JT3o���{�/o:���\'�Ê���r��]�:��<�\=\�ʆ���=vx�og��_mα����0uꋃ��ݽ�}��z,j�&;o��-��nW���xBtU�M�Wҡ�c��P~�\��i��w�zi���y5�\�^�v;�RY:�Ar����{��7挡L�+��� ��f��B凷��y����R��B����fy���j�^u���IA��{�ꕡ�|�{q
q���U|��U���0YG7tF��*��T��s�HR��>��}�E�6�:o����t=�`�w�|��}$!}�.�n�+��Gn7�*3��S_7!��ޱ�Z��V��]�B.؄CȘ�	m^=����o>gpWͽ��$�djwt��.z��x���#g$�� =���tu�L�NG˭4K�3���rev�O�!�j��c�6�I�ͽ��E��zt33��1�o@��h�4��,I��(A���6c�d����Cc�ㆯ�\�o6��>�ﾈ���.y�N��&�����C�0ynM�����Y�<��Vy�xV�/U��o��<�2��ȟ�ZS9�%t���D�ɯ�d�
]�w���g+]>h,Viϸ��k�r'\\LCV�Dt�}p6�ܼ��v������w���SJ�{嚶�z9�e�9����e��u��UFd��Z�둖�)�$~Ē�}G7�M��3V靶�k������YhwRΕ��I"�:׾�f�t{��3ʎ)�L��r��c�t�.��-P���2;voi��Z�~�M����&?Zte���)]O!�L��F�gE��vF�z�-^���8��K�x����W�z���V��R^;�us���W�{=��k\EJ��W����V7���u[Ճ�rT}��w��2	�בP�D�+ԋmI��j����!{S�g���#�r��S�x�-�)���S.޳Ɗ����!��{�t��E�Es�w��f�oj���A�4�=�7&KZ�)E06��+�)kwe��EYLP��.oNW��ݖ�aC*��w���*�X�jDљo�T#�nH�Wv@�i	iJ�5�
:��CJy�/�Ȕ�����������޷��9?f��C{Fn|�ͽjOl��zp*��O%5�U>|�4�We��'�S!sڮJS�h5��=��qʏ���X������sƚ�&�^�N�A�<��"9l�IR�ۍ��6kJ��k�
B���]�|�+ѼN�#��S��Ge!����w�Ω盒���YfC�m��7���1��)6v��9��*�E��`-3��l>Gg�6ٮ��\���'����|�\"�6-���LBv栩g�+��;?�t� @�+s^�9���_Ѽ�3C����w&�.5�q���t�/eA�f�!�c:p�:8l���Ta����I�5ء�}��p��|�d.Wr�w2k�~�$�rǼzӥ�V"D>+�Q͛M�Q~�	U��~���^V9�v����D�����꫓�����|a�T4�OS�֦��g5�1&�
�1�ķśH����n�a�b�b��g-��
��4�4�d����lT�~�ރ�1����j�H6��L�T���Vgx�\�^�b�	�P*���=olkٜj&�e��̫���A�ˮ_i;p��虀��w:�[A�>���'�)M�7b�t����7H�����"�39�Xg��:�ҡ�lp��Y��QO>Qk�&%]�<��^�y��OˈS�I�=N��Qfq�����ӳ������(��3�C<�����7�Q�l��*1�C�B�i�v!ZOL�$p��dǲ�uFK��;3q)����VuBkg�s����w���]��	��ܗ����_a��9�b)�����ʚyU�7d?s���uy����q�.1�E�)T���*Z�k-b�}�� k�6C�ɬg�B����ecwp������H-�-��|�<�/oM~�k�ƫi�>��9�7��+��X#��dL�V��!Y�t�7�9�Cy�I���o���s^��9�:�\�!s��uWLe��A�<d�[�1es�U��#�� �4�1Q���6�˛���Q�����e��P�߂B��N���!��s%��:�J{o���&<ʯw��	����oA������[R�ռZ4Xǐ�ؖ���HQ������N�Қ⌬������`r��-5�䞂Wqx1�|6[7�d�.�W8��*���$����񰼤^�� ���Ԥ�����*�ok4���q���ۊ�uU:<����x������#%�Z�n'K���vg�ލ�s����)7�o��sK�l����ΩG���⇵�x���H��9�Y94��M���9-f�t�Y�N>o�no��V�ʯ��=�Ѻ�w0�}*�����ܷk֚�y�z��9�ja��S�N<1�9�S��q�M�h�#P�Qo�A"�'g~.�5�!�O����y��L��w}<�W]���^"V0�m�gE��eI��k�#�X���?Aת.,vݽ����8�\�{���E���|��Oyd���U����������~Y==?gmj\p7㺕�vU�,�͜Xطx�V�jTr��F�T�o:��5��k��	���k�i���ꇽ���!WǠ��_D��D�{���Y��K��3O�L���7��7�x.��TnUv���T +��G����
��\#'�%D\y�orlY�����{�`�ζ��`З�*���sj=����C�V�x�0E��Us�����<[��o[]���������"�fU����Gߪ��$�L�-�/��۟"�y�E~[�{�˦cwl���B�=���s�wi���\ٽG�\��"/9��\��{k]�>�8�'M��-`�Ynrh�=��'v�\?�b�ʥ-�KT��-�tCy���w�r��������Cx+|+H���_��^n_/I^ߵ!
�s}�'vH;3�Eq8���g�¡��s��Nc����X3��op�.d�V;��C�s��r�
��J�'d-s_N����ř����=�ȭNH\�c���5���n1�9	���V�}�T���̘;S��>�S�[k��Ю�)�^S��tk���͸ڈ�9_k����`�s�ߪ���>�]���kp��]��\�f#&�#u��pʋtζs~�V+�X���]�/:FB�,o��u��V���{����b2w�y���9ga�ی9��i�����#�x���Sx�n�-���Y���uH��=szؾ���lmo�c.�.�����3��c]�L���>�s��*'��P�dC9���t�D܎��]Z���wx�:t2i\��O[-WGc���\�	C�+��婸���+N1��u�{���}��{{��y�|Udp��o>Zj��Y����ϩzK@���=C�z
Z�QD�_?|�o��U<����e�J����Q��ά�E��!\t>��ǩ���p�݁�5�t�r����ۊX{���z`��3`<ǣ����sKV��xܽ��LbM>�w��!{U=o���CQW�Ck91�L���4�fk�7���U�����b)�׍���~�sl�� ���2��[1���l�D�U%s�[����h5�C�y�$��1܃W��t�x���aU�#��/��n�wT�*]Ic�+w%�Qk'yw��ƈ��mݭ�G�vU:�<-`�]8�Y��c{*ݣ6g*�c�um#)�UC?��i���v��9��*���t,#V��t����7�%��	x��˻�_p�1M�Jv抖�;]^yz/S�{+f!��*J�t�le���_t�8�����P�t�v�O�u1s
�#!���Qۭ݂��T�5*���7}�]�-�	=����L�����ëf]��U����9��q�bYǖ����J��暛�����}Ǫ�_r��r��R�%��O8�[��	ͣ�U�(�ks��q��G"[���ӛ����}�Ua��|�����<���ȵ����I�n_͸�h�Q��`�����r�\a�Y��{�����U9�y�yc������ ��sݼ_<�پ�G�J�?F@{~�Y0q���~G!K(�Vx��ج����K�O'tj��,������dw�f?��f*��Ƨ�R_b�q�,1i�r��wD��yG����;���k�緅;���첢<.�蜿P�d�����j�ܫ:-h���Qpy6��7�o�u������!��7MHT|�U�6��J�ۏ�E�r�n%4�DK�j�Mӆv��c+:��O�33���C����z�����E9�����Sx f���`�|4���W�3����ϟ\q�~�s��<�<�hOZ�n\4f�V`���L�e�i;Y�W*/��P=z������2xI�1��g��jΙao�j���J")Ib�.��/n̕��`&���˝�^99u2%��Κt���n�4ۭW���_g͍n�oz���&�����DÏns�@\F�"bxe����55�����b��I�Ѥ��F��I�ۂ��TB��t_����n���YfW��֗��k/����uC�s�t����,�u��[Ԍ���Pc��gӤ�X�Z���g�Ƿo�7�����C�3�Rs��ٌ"����W�c��6��f�)�}֎�3�Wͽ��6�0�<�����E��#e�4	�'5��钖��w�dwk5�O���^������j�C���7������KҫI�C{<Gy�S��f�>���ES���,oXsjw[�z�o���({]�4#h�UN�}�a��Nk��Q�/�ʪ҆[p3~��W�����Iy�"Ru��͑�tE�m�曩n)����2���i;�^69W��Jq�no�kb�O7��V>ډ�Q��oU|zV�k�����7���Tb�+�$�{,�Yׄ�`�qa�z�6�51��7\:n+z�va��@���7s� ��o�G���#��뵸��SU�{u$㵶)7�j	�m��Rng��}t!;[*�Y����5b��Z���2J!��j��~+
��Z�h=g�7�l&�\r��~�憎o'#�8Vp��J�/�o��h�5�Q�Ti卺y�=��&w�g;B��y AN#w��m��P*����{Qj6~΃�s�(�뚄C�E�r�E^=Qj+"g�8��S~>�l�4k�
o�<��2�yH�;�����,�m9WWQLp��d���W��l��h�Px��Dw*v����'ι7�B��8�L��K�nn�����T2�W>!�|/���l-f��79�s1�y����\��{8��+�߼X;S��u�&k:�/BJ�1_�D�˭�PT>�ʸ�㋽�	���q��{��1U.�h��������z����3���j�}�p����h浹�u7�B��0�+;*� W�қSP�J�tZ��q�{�{�A�!���-ͥ���-��zT٣a�М3�&.2�
�Ι+�N�Z�'xJ��G���ٝ5-�wY|J|ܗ�f���>ں8p�<!ɋ�m�g�yY+&�C���㑿I����ܫ�>F�I5Fp�}l�1X�Ը���-Q��P���
��{G�Cf��';줗�C�νZI��"NM����#�m��]{�6�SiPE^+	�Ղ	�>@��e!H�]+V�[]�'̻�u%�S*D�(Դ���Q4��"�:��u��y���;^7�Z�tQ���s��aи��k4ˑ��mhH�\�'�i��GǗu�H��S�T��ՙM�]=��H:��g>ڱ��@�Ŏ���:�����C9XZ��5_5�Ӿ��&,�Q��Cl�bF�������V�Ũ�0�x-��'�'%�:�_<U2&9㗛���F���ʶD���;L�U��{�ڲ;��CӔi��ph�a]���G$E���k�L�m�h�J��W��L����{:�5ts����&���+����,�Y�����9ZK�3�te�#��1&�)ŧ�E�ug��o��>��1�L�z"e)sO!uF����4Q�m�So��0���̥b�\6��4+���rd5��J�t��w�3!᚞6N^\v�2�Tw��%��h�]-v�N��Y�:֊K���u�/�D��Ԭ�b�۹��g$i9M���Wd�7����sY�Ԗ�w;4��.�r�C��XJlK�:�W�pEKd���X��+Uaj���D�,�]Y��m��ݝ�;ݬ{���ej���8�qR��v�e�)`��wWl]"��|&� K2��B��"����Wt[�+�T�sV<�U�����u>��&f��t�"n��*ݵw��%i�Ʀ,�FT�]i��*^.<"ǻu���V���-U��*��Пn��!�%�8��K_w�ͷXGU���u�	awTo�t�^��`���ྑW��#J����@�Ä����`�3��Z�ӽ����Ȕ59U������1V���/��pg����Qm^Y�������$f�r�n=���A:_^U��s�FZu�V5j��DV�i�(3-��EH\�r��R}��o5��k��2�V&�:r������gH���<�u�{��Z�O�j�r��z�!�Uq�%��d@�O-ʷ|i;��t;��6.h��ۄ>���-}v�"QZ͡��-�v`�;�A=���u0ai�����-�ݽ��&�cYt�N΅b�ʜ�֣c���r�n�t�9�^e��V�FV�⌷�*�i�T�o�SW�q+�̝ ��D֎Lp&wm
Z�����/Lr��	fw:������EN<��sf�oLY&-)o3�P)Y.J��0Ի�x��zR��a>�j�
�=v�(��=Z��ze���D��\�����Z���u/�]����ۜ�Z�6J����\-ݎX��moXM��W�ڭ?|� �%{�\�D�P]��+����QE�'wn�"�Ô'�5�TBY�2[4�yD�)$��Ң�)�dN�[C�Ҫ/$����NR�[���'aI$� );B�Y˕@�D�����܌B�e��F�h$�C���H(+XG.�V��ΙP]$""���rL���4CP��U��
�PPjM!R�KP��t��Ά�B]0Y	��C)uu����J����uls3�vDzۓ
��s����xd$\������#�PX�R�r�G"<�E�6P^K8� �t&�C.��0L���U��HD�4Ԍ�v\��+�Q$e\�R�"���N(a���Z'\�$�΅��D�4##
)�$��/��?��3jܝBU�m�s�q����.�%M��1��6cq��\�`��r�́HwWd}#C�^m��R�_��}]�X��H�!��Nw&*q��G!�Qpճ]!�@ڹ����vkV�eS�ܼo�P]�wrk,ڥY��}|����mG9����}�W6�1��ͣ�%�&��	�.�n��5���g8f��3���2<p)����'�����\�ꁘ�&ܕb���N�A�yo=s��0��u^�������<U�p�[�P�i���f����P*,�}�0�/8��3�/rW�؋��|���8q������U:��J��5֧��s�ǹ�P������0��l7��bU����M[�8"�𢗫��#r�N'a<=֣��	4�"]���Ψ���J�:�zw%̘݋Rލmf����/*$�+����9؊r��Ci��Y�^G�%���N�׸��<Em0�:FJ����W)Z�[A�znH37�R�:��������Pb��\�b��`���74�Õ�Ҷ�84Y�4ij�ݟR�Q�}'$:���c�RMzmzf��V�>vc.`��nJ�\srN�M����S�6/����Ҏ�Xh�IxlwW�Z'j2�۫�O3qCd\������P�������ꓽW�j��͖7>�S��DzF��uMWʗN�^Ť�-�M�QNƚ�N9��x�T:�I�u�,ʠ��Ș�og�kY�ڒG��_���cO@W��a�qêsPT�_sP�!av3j�K<}�ܥ�Q�g��z�U%<����;��b�Ȕ��E���J��}�z�T,����s�U�^?�Zɨ�o'��7��L6c�Șn���a�ٴ"�W>�TԦ�d�,��U^,�#�=���O�f�Q��njq����4�K��|��:���-���Ve*���w2�V:��<�<�O��w�t��3ݻ���ꦥ��õK�wk̀���:&/��������$q�gZ��y����T�Kr�X坸���zY����fOƽ��rЍqx�9��x�==C�I���7��{��/�#]�=�7p����9P�)����j��DY.���}h�����`LA�����YI)vVms<FA�k�͡λ�ŭX�,�����ܦ�6�z��	1�{��r��e��f�g�Kع&�Sl�Wr�B���$2�M��n�we�\Z��r�]g��K��$�t�1i�ޛ��Lg�Zk���G��Lʉ�;R��^��<��7o{9�V5����÷�|�U�m�n'���OXsk;�J�>������==g��Q��=!㎗c)���QIg��AsF��;��Jsh�=�(3D��1N��~γ�~^�4Z|K�!{TcBg����?��t��/NBv��Ƿ�i�ݼO�w���O�<�އ��{pV7pj�b��
�w^��s3� /��$��B�'T�u'�cZ��Χ�r�N���]|�G*��wh�/��wM�7��Xvצ�[n��]֎>܆�ED<gi�)��=c���a[��f.̡lB?�!�4;&�t���\#��C;����֨����k"�gT�fV稄|�����zh�ܘN�.���i'�nU�0v�n�w9o�,��tc�����hR�s_t�]p'ak���ը��͟<��^k�d�k����~;��F_o]</"�ҥ�ΐ�Y����I�iV�Z=yu��p<=��X1���.��d]AoWN�����;ܼf�E�}|�r�K&�;�l�"��^|qN��������[y2^ѭTZ�=��K�sF%&� �p�=��v)7��r&#\\Ls�5�M�6��2����RŽg(jP�����o���[T{��_8f�p7�����o�n�m��=�Cl��O�#�V$�&r�o�����\9�t��s����^��nQ��X..Є�)��O��:=�l����PzV��z�5�;x�[�'�ONWgzyE��c�ɠ�	]�d�������6���Qpyca��sܑ�u�u�]�qak�w�3�.�����8w��8��ۉ�鑓j�pn�o��P�JϷ���g�au찦�1*;2u���
v��P�D�/P�X�jOO3��;��OE��Ar�:��a�
I��g����r���½��7)�'��<o�59���I�ک�����Su�MbLrJ�v\?�'�%:�+��r��'��=i�N[`c�L����K�H���|��w$���B�ը�NH^<'�尳v��i�\��/��uNy�M��54&�H�oUK�nv�{	��](Zxd��Uoi���Jl�6�Ё<��Q� �F�Vط�R��3\�aǚT/�t�f7%��pc��'`�]?[��F��qf7O]T�����,�XWXa�o3�V�jW9�|3���D<�T�j�Hox�����Qz9���^%�`���=�������C�r�+9�k`��0���Ck�gnj	r�E7ϕ��;gV�D�v栩g�+�N��7:�<�]`V*�v�n�U/9�h{�'>�L;eƻ�G"b[52_([t���υ�ؘM�-��a��̸�Y8�1���;|��mƻ���\d�j�6)>�Ɣ��X�t��}V��"D>*�C�6o��QnQn������F�Ӗ�U^V�on��{�h�����f��;�'_s���m>���t�)=��jSF�����=W�K}�xc�狼�o��\�z���Y�}l�Khk�9X�^>��4���ת���zzy��۳<�S�f:�`�f�����Y�h�~�5��kĵu��^ �#�A���f'���� �fM���#���յ0�s�֨������Vp�6��2r1a	�͚�nӸ���zM�,�V�����Z�ӺJL�v�_ٮ*��1�{vT�	�d��rh�9,19�������W5v��*��w]^\%���V{���LSuZ7'��\�Yjܩ��v��˙)��%��+:�5��#W�����3sW�|�Z�=�Ox�^�\��T�F� 'mHA^��-f_�/u1��c��j�u>I�7'w����S|�������r�� b�yF[73��ȹ��w��-N_�HE_�*��R!��C]HvO��=rKy$r��(	��x�d_����n"2�86{޵��՚dg�p���Yz�;���n�`��w�2O�m@�y�'��ȋ�ç�ӽn)%�$<�Ͼ�N_Щ�F2�_�����&�����]ߍ�K;��<����Z�)vk;x��K�g���Z�d@,*͢^�N|���w�����:���q.k�wۓ��ًfh�7#�w���nO�fxHI�V�չcսD1˽R9�R'��o�7��j-����Ϙ.'y��Mz�*�QRfJDI��}[F��ڸڇ��}���Urn"��4=伈�R��E���bZf��h��pZh����ι4�=�S1��"D�7+Y`��5{!2�dR��c�X�p[�B�����
��U��ҧ/��d㹵�r���U�36��K07>����	Cc#oUU�p��m�2���~����wB�k5��ݛ��y+o���X��������n'Yꛉs`�H�C�][�C��=��٩��P73���[�^x�Y���k�'�g�@�z�m��i��(���>�����*ѷR��9W=O�N�5���o������u]Fީ��z'|^���{�ꑽ�Vx�_�77����P6t3ߣd��r��س���!��Et�wJquǅ�J��>����Mx�������ma�|�2:/�Ǿ+~���9wI1z�AH��VMi��K^׀���{���O}9���)��Z2��\{��66{/4�腓���=8G�<�0:�y҉pi�W^ *�t�$�x�S�3�EH7�jL�u6�U�.�p="��=�~���AS�$���h��Q�#!�L�>��@]o��YVC�!f���@�xͩ��>��D��5��.�(I)��b*�qS)LL�S%�t<|W�g��L�-�/��=�RN�{�Χ����=�q�s��t�^��Z�2������y���%�mR������z�=�L�9�A>�v��Fy�����'J����~��GdϏ=�w��C���Ą�r������0�}�nd\�c��"�?3�nW\�vP�w�vЦ	�
ٷ!��o�c5�5v�������M�LevY�y37�g��[�#@�jj,���fS����c��'H�B���>k�Qs���f����0˔��
�>zWV�����2㲙���M�Κ�2�߽�\M�{}q<o�n��K{��[�����ig����:����.���U�Kk��!
�yZv������3���t�J���{�~����w��N��rH�7	���9����EJ��k��Dä��%B�w+�zH�ܜJ��d��0wD��_�k@~��;��TŪ��� �CڿZt�����{�T�P�>��n^�]��_(��}~��|��&M�ޠ;���O��;�c�w�s��=��Ea���4����Lߎ���~��.=)��7��Kz��޻��b�W�߽>�z׮��w�i��FM}�Q��R*;׏~�{Ƽ��7����ꖎ�gY�>�j�1%^쌮���"����ʯߝ-���=.��M{��E�Y�,ɿ3��N鎺�H�zt�~�?��ڜ��,�>L|�N���w�Z�;��ve��V�G���ˡ~N�OpsΝڇu�Zn��*��`	��W�S<�"��5�h�i�q�6	�=�qEϐ�}�yO��^W��}��{!��<;�9�`ʨw[U��F��k����挘����-�,���+/����.�8�����c�GO1������N
����9�����ku�'MP���=� �����,��Է�⃭��Ʃ�ťkj���iޚBX�]��L�� ӮՃ�6�"�2dg��;�:�Ȕ\�9^�܏��hZ�N�
H��FxD6브�L?꘼oo��먡�ojYdؼ�3���3�0w}�6�
�h6�sϖ�G�7��4�^��?-w>2-�S�[��q�׍52
�
���ǽ*���^��I���Ꜥ.*��9��	\o�,T-e߅g���_��=�淍z�����f��o�ooI�؉�'�q�$���L���ua3q߯G�>g\{���Ƕ��)$�6Ցd��}�s�b����Y2��ɀ�� =�,�[72��]�*�K��B���v���;��D۽��@2:ϣ��#n��UǽT}/I9 qE�@�/�l�7*Ճ����7o=�2��U�G���;���}��.��~m��u�[^s�����&��O�¤I�A�A���%��9��~�����3�O�Dzg|K��oƃ�u^�p��CX&�{NƖ#|�3*bFG3�+_%�>H��9�5q��j7��W.��	?Y��>��L�l{�l����;#}�.��[��ο.͢\��@�/�oFW���e��M��J�E�������O��c7��8��3�fWelZ�j�B�hY2�6�TFy���U�s���
&`�X��$���,z��+�z���/��V�-�a+���h�/����j�݈�p��N��"���>�h' ݹW�3���c�AL)��duݺm]����l3
�����;|iJb<q������ùiA�1���2n��WLZ^�㚽C⾠���=���ǈ�Y_)�����>��ё�^���򭙕N��wj��
�����ߩk�Y�W���Ɍ��}���_*J����%@s9�	��^�����d/PN��>��A���&t�Q^'J�3�D�_�����U��u��ە5ȁ��[�{�^	o�޼�ɝ�Sǉb�l����)�-�u��K��y3����Ҁ��������03�N߉�O�o{ִ���R4�IK7��('a��c�f�������qNC*�hy^��&15�ϩן�lW��Z�?VN�;��~�~~�y���rHףI|������Wƾ2���|�Ӑ�ڐ���X����t����v6���n��:������~�$�a@ώ*�te�u3���Po]X�Z�6�yb1x�)V�V4��K���ߵS��`��.��9���������d_�ub�Q�C��L���ͽ����h^�~��"��Z;�'J����mǮ��8'Ǟ���H{P3﷾�S zk�f��*�gYkrgv�{L�넵2����F��Wh�P\R�-�c��Lh<�ؖ�r���D��@w2�^U��vrԕ��}��Md�NJ4�;Z!ʚ�oӲ7\�MA� -Lv_P���"��[��zP�3ls3AOv�mL����3�j���8�u]f�2']Ń�b�'B8A�,����jϯ�
m>�e�[[�˞5�b�L˼�DKD�ck����� {+D���3^��r���]���It�[�S=�p�m�{��9�-C����Kt2du���.��t�w)w#GZ����l���=\�����1E+�dmdN�
�]R����M�x��d���u:�t�]�r�eNv
dne���r�n����n��#�QF:�xf�)����J�oƦ.!3��d��S]9/o��م�w�]:�ѝ�L	��QZȱR�	n����9��R�<Et�Z09�;=0^�#joBzcC��hF[�[/��عf�\c��֫���z���ݓ�����84���Z�yJ�9��@GZ�[������v�e����J ȡՖ����$�kN%�]��P9��/���#� �*�&����܆j��P"r�Z��낯�%���ql�_N�؁"Óxjǒ����z��ۦ��­�h�������E7e�1T��S�9S�ZN�&�ɵ�Qk`���p��ăp�W�d�!u V�Q�K�+�U����2�����J�n�w�iͰ�c&.᛼��o��G6�&���XUǂ4��b�
�|���7%@���k�蒖=08��a�B��'"ɼ)�ۡIfm,�	�F�Co1*���@X}�q�	��Ҋ�҅v:�y�.d³MM�7l��|�'������"E*9�ĞP��lm����;����uE�P�r�Ql^`7�[��]�e���%�
�ڏ-�S�7,|�����N�� w�HL]!o�TFĒ���,�zasw#�&��Rh��R˩&M`W���F�(Vj�ndz2�iX*�\/�vJhZ��U�n>-s쳆2��|����[v�n�)�~_K����D��4��_*���鵰k�����6G�093�50�p�okr��t���6e���a<��kzl���;��C�l��Рr�1"��̾�!�:$�m\�L�s����(U���4�!H:��"���ث`�������i���\��#��[������˫V.N7�i&峔�����Pr�	�6��U8���˺����]m(������A�#���aE�f�MJ��㮍�Ց�ڽ�ɿ��6���gH�6V��sC>6%�XaS���X��z]	K���ɿ��w����xf��Ou!��k��F�cڵPײ��A�ۭ5ψ�Qݬ�B̐J��u1�Ҷw"w��(�Mvh�X���.f��ȫ�]ќ�ڒ��ͱ�����AY�I�v� 0�.�
"�5�3�-��d�Z�w��֚���`��%n��ŏE�Ni�}y%w� $pI$�V]S�:"�(8h�W��P'Su�B��"���� �P�.���IK*���酅-%���QE�HBy#�Y�P���ˑ"�16Q�aJʵ-�P�������wvyTXr�X%�NzY���:*��(5rB��DȢ��#S��ͪ"R�Ui��s�tS"�-<��'D'ITũa��QEP�����&PI�P^E��+(�銞{��P(�(��Z'�yQ�蒃�:	�DAY�g=�L�')j�9y�+�HKA4�dYI!�"s��I�)�¢E9I��J����"����K�4EJ,�-S*�`�*�qD�P��:�Kd
HQ̒�� ���j�QW.	%Q�(�-A03��LSiDVA��:��$\ҥL���.ӹ8:Ң�	���U�.dr@���r%T,��J�m:I�ӡ�)E�Ed�������.κ=�#���o��)�*Q	M�c\���$nގ��*:y����u5����V,�M�y+���&)�x��V6��i=��{�x���H;��;�J�}�������йuE��� y�S��c]��L�G����ҿ��w�EDN���`,*͢B^��>V|s�;�o�{���g�+c�pL�V_��i�1e�>���'`@@���=��ח�ζ2<.�ȸ��H�dxπ�^����� Hݹ�F�a�˗F&�1�����=�t_���<;��)�JjHǾ��*�]��ܵ��=����`q�}�47�P5y��]R�~���c�q�=��p{�o yط=^�f�����W�w|r5��o>��g�43j|ƛ���+�����_R�����pa�T�s|��^wVG�3�W�S^���9����߮�\~�Y��'/�Q�}r�U7�=ʼ��W�/}S�x\E)�v��`N{�*^\^����ޚ�K{ׁ�f���>��S×�K��Y��'{�P2��ٜ;�z|
��9�FO{�@�T�Ӟ���)���Ѭ�=Cdb��>c���^9��vK�>��6eT;�ʤo�r�π��@$�x����/�i�Ox�3Б����n����W>O��@l�Qv�޳���v%�X9�~Żt�[�y�G�ѡ��`V�:��i\9b[��k��f�ε2�i�שm��Ǆ{� lV,vA'Q-��������LM��-�J�<����r�����R�O��o�w�Gg�����]N\�ʉ6�=0�(ϑ��&{��S�-қ�wX#�{��nFxru:f��^�Ȧ���K�B�֫�����D���+9W�=ʧے-��j�+�c�Mor�^L�̳�άt>�O��������39���bYY� �e�������vǻJ����1u3�����џy����Rt��j�����vL��=���^��A���7�׏��x�A��� TJfnL���s��;}�\MǷ��ca��:/V�U�tzo���>�l�ؐ��������-�����yZ���ƨ����m�펼���yz�u�"��T��^���`����ڣ��1K5��UL�^m8�J�MTa��w(V�ל�Dst�����>LցO�~�uY�S3-OC����7����-�����OEֲ�@I�˓o�zh�X���9�ܔ��2T?z��dC5�9�C����v�ǰEa��~�W�k�cK]��6l�>��9��{K���;��ܘ�N+�}��{�롽�@��ero��[w��\0?S2mX���'{[��y8�[�*#����j��O�-�-��I���gP�n<)����˅�[4�<ʇ{ּ����P�:^���(J7y7S��vVh����� �� �U,�mVVt�8�K�z9J5��=gz4&V��v����R�fdnE0w���\���^���,gmU�-*�dd.�T�zo�{=��x0=}>7{�;/޻5��u���=˨��g*%\	�1���=Nt��c¶����N��9W��z5�;�8�'�ݔ�y���}�8:��r�g���{���;�����qEx�m0�{��}�f����MU�4��%�#ު���W�[��쭣��t����7UC�ڭ2#N������f�w˻3}�����P�&As��\��3r!��.#[���[ږ^D��<���(��[f{}Q��滔y71﫤?MƚE\k���s�"���O�lW���9�_��^>�:�\�a�r�� ����5��]�C|����R��%��Yu�J=�|z��q�ȇ5�Î���J�pS�l�~�.����ﳧ�O��& E�����S(/eՄ˧���b|�g���}�h[ٿx6�&��Th�>J��`�f�{&w�P&���[7�L���JVތ�S�y��Yb��Oz��2�����}23�wlUǽT}7d���I���K�P|g���(EC�y���.��P>�n�q���: K��Us�Ӭ�?��X�#�M��QE������:fSg� ���\-��]`�'e�=:��S��0��zB�ԗ�w����Yl�a-i�hZcD�;	���#Z���9U�׆nK+��r�Jsp����y(�q^�׭x��>g}=Z����G\z��j�UIaz�|���&�pQ�����"R��e,����^x�f���W�d��e�������hlD��I�UR��{>YUԯ��r�J�F�d�4.�>�W>��!�ܺ�L$�G��g�;��F�G�G^�3�'{�;�$8��:�Cg��zm�_���W���`�J�E�'C�7�O��k&;ӂ�
ڗ��/�H�v�}퍨	�9�T�,�
Y���{��3�?L��C�v�.���p�~TQ�^0�O���l�3zq�hu�F�]�V�ʱ��Q��P����7s@senݙ��/m�E�c��JN@�����{}V5��(��z�81���*r��D�\���j}�0����֫3�z��>g�3�al��dU�����؎��gF��T��uDd{��5�L�>���%�+�g���GEפ%7��LF>�'�\��/O��7�=�Zb�Ϯ��ꜟYh�.��rQ�Kx�d�Fpg�Qb�f���!�l���8��D�S�?J��`��d���E����v:U��[SϾ�nw�ӡ3B��|p�Ècv��T�Ȓ���3�kN"c�z��/np�eIz�d����	E}qS�3���墵9��ʽ��P�\�΃�r��r�v�3�ݗW1���\u*�Ε;{S��ҍ�*���c	7(V����^9n\���Z5eS�L�� 'q�!����~4�>�S��1�4=[ٽH���DR�	�Pk��Y~.Ih�(qT;�2ٸ���\��zt�m�^����9;�H�߬}�Fyk�!�_=T�g�>�������9RP1T�����;�E<+5E��!�g�]��V�i��Z;Rt��o�F�޺�^N��zE��@Z�4�V�����k|��K���t��>}9�c���Fίi^��&�����]ߍ�uE�RM�������mf>ۡ�3=�i�q>�s5�
�h�Iz�C"�Y��L��]J��>1�X��(5����?�b~F깶�ݔ*?F�G���x|�2�]�pߩ�;%�O��&��oڹmԏp�f�@j���W~�j���5<+������{P��F�)�{�^�A�_r�]~j�,5��~T��~�������c���Ϛ�5a}�(�c����6ϴ�͈݁�=�;�»S���E+�����).��ڽ@zM�{�������a��(ߧ+��1RZW�S�B���ԁ[`ƛ�͔B���U�>�.q�m��K� �-F��=��z�V�j�J��d�x�_f��u,yt��L��?6r����tĠ����Έzl��SY3��fG��m�*��\�+;����yiN���h��N��,ɳ�K���P����e�nl��~�,9	����S^���9�	�ߪF��7�c�􃓟bR}4^�r��=˷�2;��u8��S�����T1���A���ޚ�K�V8K�R�ϧ+�m�ߜ�M���A����J#&:��|.��zm�|]k�<�!ҟOe�����9�1^dÅ��S�}��zF�O�U�[ڤT[���zc0�P�謪F��r��׀
��@vi>(�hJ������S��g�^��{^�;>��b�Ϯ�ȷNIf��4g��F|��Qp#EЧ�U�����՛ѯG{��1����n�>�����K�B�Z���/�Ē�&PC��msBze��<�|�~~s�����̣�}��>�O����>=�:�js[��ӂY����_?e�ړ-=�R(�����K=�{������%�M
���熌�Ͻm"p����ۇ��8�]j�S�f╚EX۩��O��8H���>�A�^3����c�5hdC��������mʟe�"]���/g9��`_�h��w�p���zL4$$��*K�6-�������}c��T��m/���Re��ƠAYx��Ab�w�I�wka;{���Π��.gU�b�í��v��K����&�T�G�pï-��yd��풻55	Ĥ�&��V��9B���pJ
ש�84�)�~��Z*Ү�����ۗ}[��p��P>�6��TUMw-��)P\����D#<4��-�]>I.^��Z?x�8��4��u�	���o�$n[QQ�W�\�Q��~�?_IOҁ����h���\���6S^�D�����:Ԭ����&'����Q�qzkxLz���rn��d����C5�Wz�_/VQ����Sx"���,6gٳ��}���=7/N��u��g�kj��z�L\bq^�q�O��^�qޡ�{��"��ߏ��ݪ4��R̟}�*'`��ji�o�~2������Y��>j�g��*{��f�k�ż�R<̗7�A²��z�2v��r�U��0�ӝoi�
���.%S���rBz��U�~����P3۝.��f��8);ˡ�B$��W������T=wn� ��k���Z�[�w#;�=껈�ULo�{�^Eo���^�+h�D7]'�zg0�U�j�����y�W��嶐�@�>���T��x��u��r}u����P��,��L��\D�0����EZΞ���g�^��S^������w>2-�S�S��(.�~�Ƽv[�뙏(�ͺš�m��*�Z"�][[N�F�U��KݤP��!GH�U��9JL�Rkfw<���3���۾6��)X�B����}�^\H�>鱮;��8�f	�����<goui����5˸�|�8b(�����Y�.MsmU����K��f͝3�� x7�|~M|и����	_��Yu�K�Gǽ�Q�vmm��h��xz�v��{p�zeJ7	˒}fP"��L�n�P^Ϯ�&m���������׭�3���f�3� 3ƽ�p�6�~��|;jY��`'fa@�/h
>���S(>9���8�u��w��5�|�<]T9y�zv�Ƿޢ5�o�F�z�ث�z��n�9���/j��.�#��#t���{і�|�c�w��֩�G���;���}�T������ê�,/TϜ�@G=�5��?b��vJz��z'�<�X�G�DèK���9�"|s�;�^DxցO՞4.]W��^J/���
�c�i�;z��?!��ǘ�x���v���=����9uܘ�I�Ϗ���f�c}��)]�tb̭_w8� }U����m��Dds��9����lo���Wr/�鐴tӚ��K��%�^�{Z�h�f��CCj'�d���R<�����V���vX�����/��n�2`�j��[�5��Ϲ�&�37�����ޚkѷ~��2W�� T���B��c�����a?k��E��D묦��у.V؋F�-�u~�����9
Y:�ʙ�9�'���:l*�edj27��m_:`сqt�jk*�9�P��\�r�5Nc�a�&�og�R�ͭG��Mvc�&	�=?i��G�UMuEr�ʉ`<[lI���೰�웱'�~9���o�\?e�^�>��|vt?0�J=����k}��s�P����"t�iP'�]Q눕5̀�Ӟ>��ގ��}�h���j�|2/N���k��C�~��q9GEӐ�ޟ8����s0:%;~9>������i���y������{�"���-G�+o�W��O�Ӑ��#ˣ]���D�:�����8A�'>�.�/UZ���N�=���b�7�H�rK�3�T��ϑ���	�Ԅ�Ǯ8�H�W]���@�v���醲+�Ǒȗ����Y~.Ih�(qT;��-�'�3����EoIz�r�*��5�^oׂ�IjwQ��=T�g��d�����1T��J�t������\�{Q�p�j��Wa�s�-��N�q�����ղ� ztO��y^��B�ʪeC���v�x��T
�u9�����N[�i�;��>��%G��ު�	�]ѤŵՏDϪ�#�����	����/L��{Ơ1�3h�e/Zc�+>9���iC�ǧ+c=K*�1VTJ��;B/�:�����j�o�ee��e��J7�%8�Ջ�������p��̆�h�G% ��(�3hc,5H�{fK��۾�,`0t�C��j�+,amgl����2�a�8�j�8���JJj&^�	�jZ]+�.�g;��ť`F@�ʱ\UʚRmUT������t�n'/��G���>�'��q:��}"�Zid��2w�e����=���n��F�MI�"O�����㕻P�����`a�k�W(��y��M�c�x��޿�����ѷ��?"�Ȼ?�φ���V`���MXE�����%z��A�������i?w0T��='=� �}�]��P�w�[&Q��i��������qw����g�t����i:n#O�j#j���׸��D�W�����oD~�Y�����}k�U{��Գo���!zΎ��g���9�����\1J��#���r;�^)*�ʧ�&�����ƚ�������ۜ+�d���@ʁ:��Zn)��U�0'�u����s���&/�q�k��ώ(���>np>S�/*�q�}t�[����7M�Uⲩ�� y_�^ *���j��jg�f��]��ͺ\g)Sg�k׃Gg�[��Ae�rK7&����|F�+����ߵ�Z���%��V��e���TST�/)֫����1$��@8�y�RÜ�N];W1��}��(�\�@v[lLzE�
��f�%e���6�I�����j\�ɽ!oc,VnQlVc,����(����G�!���]+�ܴ
�����o_]��y��N��:�9�#���P�OS��rR1��Tr�
`��y�]v"otN�r�����aT�;���VE5vSjph��m�w��Pk���m�
K��Z��ղ�dcKR�)�;�mN3kMdŗ!�.�W)�������u�SI��߳�K雀����!ت=E�����{g�\�8{bJg3��!D��R^WR�=C%�T�j�y��&$�X��`5�noȝ�/
[��R�ZXh�V+�4�P[�i�XZA��_��E�Օ�&�&��J�WN�WZ�CgP
�驲.�>�R�a8b�:��۪<&��q��-ڧR�F��*�\GP7���:�>́�<Ԗ�"ʬ��p}s�ݽڷ�U�}����^A��K��֫�������a;B�ZD��U�e���T�w��o(u_^ᬗl��ۥu�b�t����qw9�dK��}[�P��z_fb;�,����P�*5&�Źg��f*U��Vm)�Pf����@g�V���Z�"4���N�d	i�V�Jkl�����<n�$Ҿ�r�j4�σ�1]�nF��5�n)ZA���t��z�$�n���ٱ1�s���q�X�Y���!�hWz�mR\{)3o��V\3�k�[�ۙ��j��� �U���*[�+���#��,� �����������\Ej+��8�Q�X$��K'^Z�s��FY˘�^C�J���.�Zh����j�u�m�(�T�vݾF�TdfdHi-Kz�5uV{s��yՂ�i(*�}{���!���"=��@�kņ��1N��/lí�x�G녮6N�X���ָ�f�a���gM�"U9�9l
��b�G�%Vӻ�9�/��/��<�lZ���ے����'�ͥM�,���j�U�N� �5u�Y�yNsJ\��\��J� w�:{���Ǭ��s���I!�Q۫�f�nL����3)���������:�j�En��>���wg��|r�tR��;������*eG�d�r��ȉ�(gd�9b��[��u=*���}�
�����6�[3sO/�����k)�[�2��0MC-f%7k���̏'c�u�2yӅ�	p��%�ZN�6�]�:���I#�o����s�GJ�uNT�v�nwiyZ��:�+�̨�e�1���z��ز/�NU�`�W)��Z��g��Јմq\�u���Ь*����5���r÷ȥ{\�7[���V9,ݬzr�^Yr�JV��3���Wyk捓���N��{�ry�7u{ڄ���:��ơ�x������t ����K�;���e�nQ��\5����Y��r�b��ڛ�Σ�lr��x����{��;%A���=ha!@S3T�B9r��(�AE��Eʹ2�5*�sX�,�h΄dedf	�BHBbKJ��j�Y��kB����ZiY
IE�H�"���9&rYSNVd�"�h�̒�6I�'1Y4�I*#�Ց�5���Zl��А���d\�rr����i-�%�#ÒF	UPUT,�3:e\�\���
-�b���%@U�Q�*(�ŤEP��p���H��)�r��TQFV	tR�r��Ps�1$S5�QS�ꊒE!���T�-�D *"3$���4�E�U]�B�D+��p���UK:BsY��d�r�""�6�EU��+T)AZD��B��E*NkNʲ���Y&t���sK4�
�AY�YX���"5(�B�t*(�V��6Qp�����q6T$��*p�D�Qi�∝Q&fZ"��z����=�nl P��g,�NRL(�ӊb�^ņ�l!�#�&>��i���Xf��n�gb�x�{�v��JWM�N_$�f~�$�L~�t�Ϭ�.�}��o�S�������;�v9������ޏmኹ����f��H5�3�L����T�^��a;v��Fy�����'J������L���V_^{��y�[�Ġ$c<��@^�(	� q^3��z��V.5hc�������]��fϢ]��_:�Ҫ�E{ޚ>7�=��Ā��{@T��l[yD!����xCq�(3[�U��*�K�{ӵ�>���ޝ�=Y�s3.uznO��B3�R*%K��!7���+ƃK���MF�Lz��nM��@�<kG��C5�?]x�U���UU-NA4;.�;n�`������+���wNѽ>�Q�1���]ɴ���7ޠ;�,g�a�x>g���F���d�_s��";�ӿ+r�t/�Xa�v�׳�rb�8�I�z} �����=c=n��0�[����~��d�Q�Z�t���������1F�Xb�J���#�2�|�M��"�]<v�m(���w��^�r�o�@��Ty՜�^t��������i�
���ld����Ή�}��8{q�3��ﴘk%�ل.$��'�)�ov�a��,��q]܂�B�]�tL�D	���F���30r#.�-S�:7���}W!�c��`�\��?H����|�\���c����m!˫��8�Z�v=�k�X�-��9��\�mRV%y���s�4==9�����nP���;��ݘss8v��)��¼�^����Y�����D��Dd*��ȏ{+ȭ��z.7�[G����{�[��ʨs�؝O2��*���vu(K��w��Q�	��*�t�%�^#"]x?�]Fn7؅Ʒ]E��Բ�(�o.ۇ[;��{5u��	�6I}1,�Ҵ׊�05k��ߥ���\y8�c��s�"2�rꔪ]Q�>��H>���P
,g�*��>Nz"̄��2�½����9�v��U��]�}*���8�/ʟ��(2�����2ٸ�����fݿ^�q^��5UF&��[�v4��_�z�=~�Bt��������{&wa@�/h�ْPzz��u����_�=ܺ+н
���>s����#8����m��ث������9����ځ��|o7o
�������}���9�0��^��9���v==Z��z�u���j��T�-z�|�&�z׻#��#ss��ҿ�ꉩ�������h�iuy���'+�5�T?Vx��K�����~��������-�7m��^�]�tȃ��I���V�v�4��e�gcZ9ԫ�ar�bҧ۪RY&`zV_��Y�[ۜ���g9g�E��l��л�^G�� b��B��[zE\��R�ǀ��@�P��n�7�qNg:G��1��T��E+F(�y�hN���|��ǰ��^��؈������}g�%�	���	X�}�s��8��Z��
K)I�UR<�M���m�}��e���`�J�E:O6�'޺wD�o�y]YL)�DoK��Q8w�!��{,ɯ���yd	�1뮭�t^�vGS&f��S���}{��\ђ�{��_�n��禇�g����\/F�]�V�ʱ��Q���P�'�h��Yω�����m����&�Ͼ��B�U{NB^�;�#}U�+7׃�!�/h��p�}>����^�}K�$���㶚�Y^���U�Gx�8�uC�3��q�����3�ܾ�^
���b��꾬�D���斥E!`�t��QP6PwS�t\S��:�>�5=��`gҝ���׆�����3��՞h�f3wj���vKy�`�>�l�7NC+L�.�w Oؚ�D�'��	ҽ��;"�v�:|�N��`k�Q�~}t�E�rK)2�����2�	�Ԅ��i���w��)�mA[q�����\�c�c�"�ly�Pk��e��%�0�LU��g�����Po�!����#N]���/*F�nF��t�ټ�ж.���C{�a�"��O�=&��ݔ�)K�T���ͣȾi޸	)��|���Y�Z(oM/1�� �ъLY\�^��HT�>z�!�VP�Q�]�F��-΋�Kw�[a3蹖<�Վ��Z�ϟQ��T�exz4�����(��r��ˎ$�n81������QA�kN7=����{}R3��V�χ�D���V�������b��Y�D�G��T��&��o=8<��Fͯil������{վ�y�t�wѫ�z��L(�4=9Tt�܄�݉H/L��u�5�¨͢|����Sq�V��ұ�6�t_g��>���@�X�(������Cݟ�}��������D0w�^���7Z��ai�
՚^��^t��}�>���h�g�����mTԟ#��P3���=��:|ճ����z���#������k��q�UɼN�߽~�����T���?��<���Vܲ�V>�swꉊ���6��_�5o)M�v��KӳS#{�|s�N����#=� �ǽt6��4��VɔU���#{���)��KP�����R�u/Iӡx���;����2�}N|s����L���ؘ������ԗ�Y����A�QCܤ��TB�:=�9����;l�3�P�Ī{�s���L�6�xSq�t�^��l9gT�Y3*�T���|���p�>������K����0/�Q�t�֐��&C�#1Y�+��;���[6�T��U�:y�E@dh`�]�ٌ�a�M@K�ƫ2;���Y0��Z��o+�j�_`�N���Zǃ�g%_�@_���͹Ï��{� ��e	�X����S��X�	b+|��]�7Q�]��)�+�=>��r��N�*�q�}t�[���"�7M�U��ʤn)�M�16�{ٓy�׻�͏h��Z���E:�>{^�;<�ظ�>�>�NId�G>3�'�$��oޘ�w��B\�G6Ϣ��L�(.�@L-u,��7P�L�,qy\��t�^�$���e�':���C�����	�g���t��*L�Y�]��ׂ�}�G=�|{�u���ׯ��5I9�J�ț>��H>�2��(�[sS)zr,�Nݼ�ў}�h�yIҴW�lK�녠�V{�*���'#zj}BmO��� 'fP � T��7�)��M�:5hWyB�N�Ͳ$�*�F�Vt��нK������>�u��M��v$$��*>=/���-��^���}�Uܬ�7�B��(�Cϼ���;]���	���\ǫ=�V�\�/M��9�d��A^��: ���o����Ѿ�9^�0�k4L:���&�� }�8<�3Z|���]y)�u�#�;���q��[���7�㷛� Q��8볪�*q5T�Iqz�6����4
ٹ��r;��	cU��f��)��zk��BÏ�PK���SS��d�]b�'UD�;���Yv^<���Y)WhLL4���qd��N�A"N�c#^�h��2�y+Ա�����U��;F�KӾ�.��iK�2m��{!��+��#75�Ļ�h����We����꺞+>Xk�iє���wZ���^��h����#u_|��`�uu��^#�~�.krv!��4�I�5	�G����Ӣ��qc2f�
�vG��<Ct��0=*�"i%D^x*�D%6���D�^����d��J��a�VW��s����ǁb8>/���9kw��Ό���.�������(|�uo��ז��w�#&�.��w�eV���-�U{�v�%��z��R��S���)�3�޹|{м�Eﲶ�g�7]'�g��J�+�:��t�q��W5�/��uZdzG�O�*�@J^��3�u��r}u��b��Q@�V<.���O�ُ{K[�ߧ���<�L�1S������S�#a�S�[^ˏ/w?1~ߥ�Hٻ��9�=x}�=ƙ�n���E���T��U>Nh�}���_-e߅e'Kz���l�*���
@�F�u��sZ�<�vT�p�.I��@H8�S-���A{.�&[B�]��^��֨w�0F�6�nR,�����Q|݃�=a�3i����FM9:�"�ף�ΉF:��:�1��*B��$�Y����k�,��S�Z�Q���kws9|\;ohuc����R�Bl5�:�`�A��K_I�G�t�*&]��Wj�n:����?�~�{�'�W��Bt�?_�=�;jY��`&(^�}-��;��>���/[[ _p�?Uڨ�?�A��_�f��F��~Hg}�b�=��zH	ʉ!4jz{���'˯��>�}���`0��ٹP�W�#��w���OV�~��G_��Ư�URX�&���"�-�e�۩��O���uD��>�O�d�k4L:����'ȟ���� �0=1G}�nmq��	�������,o��sm��j��|X���]�j���Dy��v�w{�~;jbK�h������)�o����@�Bc#�Q�w>Gy���E
�鷣��]���[���YR��0R���޻�۾t�Y���GL�X��V��P+��%z�G�	�1���7���JD*�V�}�����C���\F�W�#W�x��z�zzr=����m�ߕl̫���0���Vq����y��;��4}�D�<�mux_Ҫ��/H��}U�+7׃��/h�B� t�d�(E�g,ѝ���63������xޛg�:tz纡��gY����ު�Kb}x~+ʾ���^��K���rJ��/�J�k���l�>����n�	נ���O�U�/s���/�lb�93u��9���k�# N���;�oE�6cQ��M��MjΣ�Q�P�
l����r��Y���o`�]�sS�w%��1��f���g��ӣP̯6F:�z��t]?!�+���}pj{���Ȕ���я��Ľ�w�]�)�>�}�i�oj�Q�d��գn�|.+&����e\l���P͛�<���f����R�S�_S����i��}����bߟ]#�[��3�T��L�d��&r`=�]��g�VwG�h�w��j2�iG���ȯ[G%� ��f���rK��0qT8�Z]Ϯ�}���A=�cy+yG{Y�TΎg>���V;��Z���C�p�S��`��-���e�p6�n:�E��V%��=����~7FY~9w(7N����>�):U�}r6�ul���������Nk�+7@C�!���^���S���N�1�w��v=�@t}u���X�4�gZ���X�&�
���t��'�?��P��|n��(�Q���vķ	~����y�5+�:�t�:gQ6�뎁~���\��IS3!����F��{q;�x}��;����'����i$�|E��ԏ'�D�#�|{!����}�n����y��ajG��2{�<���CФ�H,�}}f���g��gV�xyX\J�z��:˕���W����\�6�c�v�|=YQ�&Gƣዮ�J�V�����Wm��P)�������fZg3�!x��$��RГ�)�&�-X� ̋5�����S ov
}֑3�7�`�̹s�Q�\Z��� �ʄ~L��qMI�������_����߻ѷ�z��7^j����������[Ͻ��ן!>����Q���;50�7�w�S�=%�@u����O�����N�L���gҶ��O�*����A�O�����t�����]���rCYU��s��,��:[�Gvj�fu���W��b83��'.=TB�:��xK8N(�`Lg�ዕOr���VEL�����7؏���Rߣ�x��ٷ8q�zOvA�@�:�fp�9�*��&����Q��}��:�����v@ȕO}9���)��Z/|���s�_a�F鿌��92�h���^/gz��y,Ć��}���H���2���8�^�����]�[�$�q&��&;*+=ag��)ZIf'�g���	�'Ö�V��fẄ�r��K�B���.�x����h��_{<���G�$��@L�G�*g�be�g�̢�z�s�T��9�>=~��/Aj��b'�d���|=��q�(�j��e02P4����e/NE�	���xh�>��g+��G��7��I�3f,��{&�R��`׳��ٵZ�؎CHy�L��i�WD��51(�gi�R��~�8�]�L��nkVhef�`©�]��1�C�#�z�9��c7yf2 ��[��PU���=ݍ/�����魦$.n�٣�`_gpKv��f�;�� >0���g���ڟz$��~�����3��z�1ԩyX�`FŜ}�}>Kz�j��N��v�R�o�o�'���qW�M�׵z��>�1z�E}-����ǭ$=��=�j��s��>��M��z��g�*��T�������$#�ZFe@�z�����s��u_zG�Kӵ�&<�h0�.�Ioҁ���}�ցO�~�ߪcP�m>O7�+�Ù�|ﶤ�s$	��b�������	�\��M�R�L���@w��k@��t����t�<^<���U�?Լ��QOբ��;���;��]ɋ�N+�}p���F��Ǧ�Z[�Z����s���{E�}������4�~[��gF�Xc�G��JB���/��z���'�����}����z���m��l�9�9Q*�7>⢜�:.���c1�귽�>����G�E��נ�NO�O�(�~�p���3���dT4wj��p���:�׽/�r����ȗ{H1�����Ǔ�ULo�{�^El/+�o���7+���+�b�W��޼�H���b�]��KHA����K�R����\���X�ͳ�m�^M�x+(��}��o
c���-� �@��*Д�+Eo9����(&�yf�꠶D�2����gV�7)��RNZ�<G���̡X��'���@����Wp\t���J� ����5���3{�[h�'{θ����z[�ξ!�i%`�t�}d	�jQ�U ��A�ې�ثTI��;���\	_�],a�ܭ��nN��^�6JV7�I�"��#��6FT�'��Ef�17v&�����I�Q�Y�}N��;3pηPJM�\�S#���q��]F�|��dG1A�_YB�V�t�W0��h1�03����Q�[E1>z� 
��b�\	K��*�/�I)&�t���\�Vv�҂n.5s:e�g�w]��Wrڋo%Zu`9x�	!�S��}'��;,�\`9��*#��S�4fgs
�D�mK�ss�sYY�qyZj�b�oC���5V�J��Z*Ў���4�kHi�19�hL��Io'|�d��Q���գn�F,HTz`��9�K2���m;�[��֛B��?[�;����H�o;��@N�\/�1K�rq<��ߢm����3y��GB��E���a�����V��-B����r��\Q�pEۋM-�����Ա�>���7���mtUnCN�a�B��;J��o74���C̻��g!w/{@Bm�^��o���V��36�V��P�Y�i8�R�@�R��w��yw�:��wl�Rt5(iY �}�Z��h��!�\�
���w�,!���K�Wˏ����U�P2M�{�Esy���s�	�8cv�,Xr�Zͽ?^�a��6`୨���lܵ�):�b�٤w]:0�6��X��yV��3_�smݱ&�����ݮ���6�r������+*�G��L�G��!T���G�
��]滱ƞN�i5cA���b���m�� �Fw����`WP}W{�N�qB��O7*�&J\m� E������=��o���fNn-��Z���x#��f�Cv����b��<�!z�޹v��,��'��j�V�[��
U����Ǩl�vfھ��GF�
˳;R�@�S�	E��y�u�.�gU��9���X���1H�����{�ϴ��YW>[n���J�d�����i�v y[1H�Q�էa��f�/�l���}�����╵G�1��b7�'[��֎Z�1_EL�!������.oH��*Qur��`�C�Za��t��ėـ�6	�6��S�!���E��v7n�A�,���[r �P+^�Zz�����J9oI�S��������]���WZ:ɽ۔{���dUr3��:嵔�0��n�_i�D���6N�.�]*ɼ�$��yR��!�^��gg3�M�*��X�(k*��a]��|���/E٫��:�&�I[���[F�'�hh9{ʢ���N.vu����*�ֲ9A�H�T���vf�EG9\�*"Il���T�L��/CJ=@��8DNg2B:E"�q�PEEtDe�]:j��E��J�qD�T" H͔*%r��2�N���������y�.TU�#�s�B���T�䞡y�V��EEDuY�¥�Tr�"�R�)$*��vEj5m(�U%*Z@\�U�\��3�+$�c���Au�hG%.E�0�C%�%t���!�b�YA�J\����"��\��D�V҂��D˗$�U*Uʂ���mR
*5duB���9�@�ՔFK**"�H�+ԹQ�)%�C�g6�Ȉ��\��2�PJ,�* �p"
�bK���BԪ�QG+EZ˕U�6'**":)Q��E���:r��A.Y��eQ��U�E+Xi.��Ri!Q�#�Df�����4��M��*4H� ���{�oF��5���<�aL���}�+f�6£RJ��S����F��M�
_��vjR�,�R�p�f�f�q]"�mQo����"�ʟ�EmV�G�O�*�]0��x��^�"}u����g�՗5q�;C�p��}��X����K��RX1���_�ܪߤ57k�k����ȸo��U_bh�/�-{�ϻ)�>��=Zͧ/�xל�-A�
E�*P��s�d%{������[�VvD׫�Q�	�h�s��?:�k3�a1�RͿK�}pe �,]L�n>����hy^�����wG�j=MV}�|�g���\{i	��^���R��`&�0^�
f�[�N�\3s{4�ϒA=G�EL���]�z�T�8d)��=�?Q����T��]�{�G�p�H	�{~]���:�7ַ�v��i��T
>���ܨv�֑d�3㳀�����R�;�MZ߽�/WF�H������ �}Q52�O�d�j#4L4����s>D��wĶ�Qp.���z�_z�xݏ8��7��6��`LF<�Ņ��^����؈���5��R��O_|�]qw��掯>��p;��� /<�I��UT�,B9���s�5q���u��?v��-x�������١�/{ה��R@��7��t��W.d�^{����``�+bj�k�x}�oQ]أXdd�ajԌЃ[RN#�w]_m7�wzI���s̼V��͹"�x�X�.��g��R��-���F����A3�+��z�	K%c�ȩ�)~�����_E!���z|{>�����2`j�Y�^yDyd	�1눮��]��Q8#|5K�]������/Ы�����֜�H�}����zhu��m��yV�ʸ��x���_��w-�n;�W�i����7��5]L\D��iK����UxJ����z�$�/-Lي��Ww���;�m�G��3Pvt)ɝ;��'Map'<�Fy�9W�|r=��¦\y�}W�b^U���|ѱ�=�5^%���5�"/j�������ܯKc\ޮf�ܙH��{jgJ����{����7��֘�=�ED[���A�h�Q�ɤn)�e_�4<��ؽ[�y�~��#= zk�'"�7�S��P]j1oϮ�ȋr�fbѨ2����|��j�i�Ι���{|�~G� ���Hc��j��Ɵ�Y�<��ly�yH<�;E���\���([�����~H�c��^Tςf�A��x-���q����Lq�W��NIy�7�B��Ww��&�����oO�S�<c�0�g��(���Pw��ӑ�x�v<��^�T���~�W���j W�mp��R�ܼ̃:�S��9g!JU��)ϻ�A�{˂��dYOٯ�I��Dن�U�׉��G}�+2��`)�c�*��y��RZgnְ�Y9I��@�=9rك�}@���9��pu��Q��Z�jZ�:�5d�.j3u�{��$r8��>��B>��=�/LM�)��zpyˤ�';��/�쾯`��,R{�iP�O�����û�h\�����<���<26y�x�¬�!φ�q]d�sO%z^	i8J�W�c��,��L��q�/��g�(�>��*���|$�}R*$�ɯx3��E���eR��-�C�+��#ýΤw���>���*0z�p[��Q�U5'��Ƨ���������j���j�yQ��r���Q��9*�7�'^}��|�����z6�WнY��q�#˾�}�;�M�t�p���6����>�izvja��޻㚼�����������67 ���e��}�k��	+ݵ�e��SOJ��R��7Z{㩪�q_i��Rߏ ���9Y�x�tn�NӀ�	�G�t;�o��􃓗���t=���x\S�'oe�9�`Σ��V ��u�sԷ�^�j>�Mx��޼_�6���;��НE����t����)������y��6=`{��` ��p;�U���{ӃܧayV��ڤU��}0��t�ʼ�*��m�"��vZ�����b]�Ff���h��I�=�8K2K�����l�3)�z�⨮u��n��*5���M�εW��k�@���a1t��PWv��I�;��徠f=�Rc9���9��Q���-�ീ�)]swq$"�#nS���!w=�6�V�'+�z�y�9�X���������T��,�t/��oٯn{�j�����_e���-r�u,�s	�j�Y�����c�ES���U)�h��z���.P�u릗r��M���,�.�z�[�T��9�>=�9U���"�]g�긽C~�W'���/������$d�j�s�L��Ϭ�N����,s�&/Q��*�֙���*�ڮ'n!���=�;j|n�;��Az@�=+�l��=��1��ݻKk��ˢ��*��!����q>�TN��۸��zh��&�^�s&eB��}���s�`C~����H(s��>���ޝ�Y슿��T�^5'��`ed��%9�^Ԛ�J�4�z�T���k L{�4{	u�K~��x֏�f�
~��1v�J&�+=��K�8��S33�>�ht{����r���o�ï�uܛ����7ޠ;��_�)����QU��ѳ�a@W"��ܫ�j���gæ�D��:�X�^��ۯl��j��_h�̮<��/E��c�@`䯠}ލĒ@���H������K����K�mu�jK0���3P�7���]��_l��`���KQ����H�,�̄��YǬ�Y���2���u�-�QNV�ᙽ$��a�A�>�{j�JO:�e-޵��b�J�ʆ���\������ o��2���c��(G��Ӣ�?-�̋�]��<������"��g�h���vC�#�Y򿊙_}t��o~�FQۯ�:J��w�eyQ�:|��g��/ӳ[����H���������������c��lo���/��ɇ�CVA!�<����4�ߋ��G��?�f�Z�'|��3�>����B�c|s���+ay^��a��:_�wM�]�~QJ��/?,
��$z ʨw[U�⋁�n4�
��t�%�^#%׃�>��ʫ�1:��=�1Op\�3gP�~�g�*��x���(=t�򘸧!��>+�]@����G_���R��+b^v��P%>ge]B��8���|k�/Τfl*Qb�RU>Nr̄��,V/eg�Nu���W(=�衼���}Gǯ�w�sZ�<��R���.I����8�S-�"�~:ǳ/�3Y�"�%��)������T�X;�O����Gǯ�m!:o�~�\z;&Y�{&vf�Fz~T��F���i,;�<T���σ�Taj���
�h����}���z�ث�ު>�xU�-D˼^���g~5����h4 m詂I���w�Q6�R�M��j��b��ǲ�!]0�[���YZ�@T�ԩȷ���l�\�j�/,�M��w;1E�+F����{��M>͌���V�/�d�9<Y!������6��+ݙ�3�k�G����������sO���s;��匿A���r'n}��W̵�gy�4{j�d��<쿱����/yq r�='T�z/��~��Dä���9�"|z����/=c�v	��|����D�<k@�u�йu^�*������	ea��6_�}�C�nG5y��$l����^IVg�L{����zg�;��5�Q�y�zM����	��oFE9����CZ<�.kڗ)���~�X8\rWr.1z��n=���f��y��fMG�QPz�y%9;��6n�N�g^�7��>27N��=�t��^���<e�ǧ�#ޚ�Q[U�2�z���5�';�j��O�ڇu���zN�'e��>��@w�F���VG����'�^=/&����x�}�j���r���TQ��·u�Zax�;\	��w�� g�=�� ����w���y������1{��W�o&tg��Sǲ!��eu9GD�<���1�A�������>��Ѽ���3 ����'�^��Z��H��;%���Ѷ��u�H�9��۶'�>�a�}�X"�<T�o.�Yy\^���CsOi�yu���[�u�[�;
�2��}z.t�������+�!�$p=������
ʸ�a������+��t�cX���qV7��pl<�|Rޑ�J����K%����mu�i���˓�X�}����z�ydZ�?=�EE�rK�1h�����V{�ٟwwG�pK�Gy�譐�6� �]X����u1垻c����y�h�p�.It=�J~�3~���sK5vz2��Tl��v*e��2����[�-N�����LvO��=���?v�{�죏�MT�d߳���MĔ�1T��qFQ~9w(;�۵�>n{ţ�yI�ϩ��@1l�]�}%\_P� ��w�`��>7D�]��
Cځ��'`�s�ǻ�N�1g9{T�����oe�*JΜ^L��q7�������h2Y�^��L�Ȩ�u�5��Fp�U���'*��wG�ڒ���w�1ϕ���������P����N�y?����  �_+���K�}��-���v��=���!��]�m��>���������A��]������Z���:�ro���+W�R��������v��zk}���Uro�>�x>L���F����q�V-�t�4��t���_~֬)�(�c��n���>�q��ں�oz�jt��g�@����ˉw��Le���߼�<=w(�O���|9[i<+-aA��q�R�4r��׶�5�<R��2�07�4Y�mN7�I[C�W��=ٵw��s �}9�#�ubB� �x]�������<�k�5�����<��:�V�.��}�$~៞��w�j+��������>z6�i:tw�Uk������XS 9�p?N�s�7a�>J���߮�_�՞83��A���TB�:��ttS�'oe��+���p!��oo�YΌ�G�2��!'}��3�ܾ�^/�k{��Ά0����OO�_l����7}喐�p=�^�#"y��D�{��zp{����}t�E��/���ӏ��~`Qy�ѣ�7��M����?��R3�]����@$�x�E:�>{^�;<�ظ�|��*΁�r/�}t�{���G�$����=P��2Ѻ.f�g�_��	��������j�W�3m��r�w��E�����/-�K���@F)��T�S^����޼�3�臽=�C����)����u x�~k�g�k|}���p�T���(	(�71u2��,�ME]8������9O'�ԩt���D?r�#��'J��j�����@�񿞉;�(	���x�-�Lt+��}Cܖ��V_�Ձ��MZ�}hv�Ը�����q�qW��񸇲`y�@����E��{��+U"��� VjA���ڀ��>��D����O5�j��eE<3�ȾT�{��j�������2,Z�S֜�����\k�Wk7�_ɩQT�9k���V,�=�=dg�WY:[@s�ʱv0,�^�&Jc7z@��L ��������D2���yd!\���;]���	��W��:^$���?�ֶ�U׭���sY���>$2;�Ae���0�j��Iu�M��@�<kG��3Z�d�x/�~�u�@�����`�X�sU�%�(K���;k�v��zw���ڤm)~&L׫��1����Xﷷ2Fx
�xց\�a�`�Uu>+ t�,���?V����������M�.�m��:Z�ײLz�&���ֽlmϘ��c(��}�B8>��M:/��ߌJ�P������3�{7�3�ѻ5Jێ�]�����~3���q\W�*��{�����bsL<�b�o�w{��坋������V�vx!ѵ��r�ރ�r�w�?T�1�?V��K��q���FJ��`���7���"�l�}B�c�t�(r%tF׀�{����dt*�7�>�{+ȭ��z=E��"��rc}�����g�G{��//W%-P�\�JHu_�UA�;����22]Belz��������J�Wy�g�Ʒ]E���%��3��Tϔ��9M��`b������t8�k۶��u�Y9�6�jHyd���K�[��)mp�Y�J��u`{�fŎ����41�D��S�5�u�;AXY�I�;!M���]�uv�._=����>T0z�J�)-��q�&��gP���>$g`
7����l�}(���T�[����Q�~�Ƽr��Aw����e/�T��T�{2���c������2�y���z��
�u���Ǹ9�a���-�\��2��q=��ʎ��MO]W�r��/k>��tsȺ�����^���{#�Gǽ������ǣ�e���	�^�����2sw���p= 4�;S,>9s	J���V�G��~�7����H���v�+�T��������W�C�g5�V�Ȉ�!���Wå��˘jz�8�w���OV����-��j�>ƙ��`_��գW
���	�O�8H
`>�����|*��Dä����=�Uuy~��t�e޹��d��L�'�5�?M���N��\����&�T=�BYXkv_�HNs�����)���\�ԣ�Ӫ���Y��>��w��������#�$>�A1S�^Teچ�2�>>����[[��z:X�ެ�%w"�z��}��7���7�6�/]9yDy]�G�'w&�ܱ��}N�M�Ei]�^6jXĽW�:�#�gɏ��U�ɉ�V:r�}�8�H���uu��iY��M�Z�i�����ǣ�2��6,�"x�`Nٗ|�ja.��W)�������q#pZ�l��u,u��V�MY�aMͱCo�C��p�(��x+M�7n��KtL:j]u#b�z�T��ㆥ��F⮝GjhAG$Y�}��/i+�;���NM�����l�6h�pa[��ۤ�u�̇�&�����vCd�� f˺ugW(�c��`"���@]d��y��j��㈲�`���Q�{�f��ڃ�W�=7�L��k�&�h3MgI�-9���{i���vS�(�l�z� kE�*�Zo�<OH�k�-��,L���#��կ;Uu��VX���F9T�(�G�*��E,Ǯ�e���ƻØ��i��x��B��:]����H�@�k��C:'.L�΢�,��4��v8uG�dq*ΖN�e�/�!Μ��F(;�{f�E���l"�=K�I��c�W���k%���$l����l��2C�g����q=z3�p����\q�l������g��l��ۆ�2�J����A@��i��dn�%q{BŖ���[��p)=���C��Pa�f�k���0��.��[�T]\��7-�z蝥[1�y�e�Щ�s}�㋴x3ͦ�����[���X�&q�vYe�5�R�,�T�sa�:,�ۙ:�>;��銻Z� ���.��]���C�55�v�ī;w��#C;z�F����-]�j� Kt.�دFf�$C(Ya)�py����Du�v�w(1T�dW�ݕ�`�72��c=�@������ ��;�ˠ�8�������KA�=��9�DCjq�Z��� ��2���vN1j=�*�W�S�.q���34E3/v��>����*�P{ݼ����5���Қ���OM��v�6s�>�}�m3S'wy��ٹ�6��y�n\�e-�\*��Nά��8_H��:����\[���Zeu&���u��d�ŷO�Un���\�����k"�\��K�0#�g5b���]��v�%�}z+���3B�w�*��s|��Vu��rq[��&�\�`���0��Ӿ�6⦑VkoqS��J٤*�-uCe����3x�s�.�Dj-�e��/��o�����90�4�ꥯt�z0��u)v�Q��i���kiM�yi�;Ql�F�N5��v��3�ko�S�ʺ�� ��*7h@�-��O:�fWz������X����)un��:�b�q	9:_8�ܻ{;_V��'e7���ɚ2��A:��ה���h�M�Y{9����pNع3M`�LhuX�k�t����)۔�N�a��d��|nS�!��v��g9�2Z=OeB5Xn���ԅ���w&d����8�u�F����Į�*A��z��)��<5x��ƺZ�̗6��qMN����$L�s��hؖ��P.e�k�|�X��)P;��4a}y,W6�#�c�;� ~4(hR�O�(���;�Dʉ��Y9$�L��wi9EQTTUR!�Z$�9Ty�*�"�Ȃ�,�U\��j��:�TQDy%QȺMa9�Iʠ]�
��W+�y%�S�
*�Z��qR��A.ȏR���,#�\���E_��DR�j�kC
(�EW2@�4��r���'�n�Drŵ$-I0���Q��YHQG#2�T�I�r��9&���*��#��d��"� �*�ʊ�
�&��Xs-x�9E�9��EEEQ2
!̍x�E3U�+��P�J�UTP��"f&p��B���xy�hB��*:$*8s�!W(��tՑT!��4��*x��jL(*�"u�*��R�UAJ	Qq#̪��:Aj�I*�^뚜�I)R�!9N��VQI�ʂ1.$T�ZBJY�
�rt[-x��Gu���3�
��kJNY��Ids�<t��,E2"�_�ù=���?�{������u�ǨE'�ָ�J�=�����+Ju���.@�-�Hڼ/�N�b�}�\1��i]Q�ޣ�CɺFC��D���_�����Z�Qv�2�w�e��}�%��w�>�
~��m�Rͥ�v�W�������9��N���#0vt9ɞ2�´��{*k�RrGl��J�9���qA���a.�X���{�x�:�2�(99'F�9SzXv>�#���;���>���)��>�c7���1{��H��-�N�Q�&���=��=7}t�5%�Q�0��C�q��	�M{"eϟ���a�S�c�Ϯ��r��EVW���᝵��7m%���y� '�B��U�����c��L{����ϸ�{�f=���2����݋�j�d��f	����ї�$�&z.eq��}%��}D>6�Sbe:3Ҧ]�E�Њr���~��U�R]�����ȁ�����d_�]�ݻZ[;��ߧ�ĽZ����H��)@t�\�Fy�_�ϠztO��d�����yzb`'��Fzpx�Kj�2!ֳ��|��U�F=��z��a�WG������ƅĺ����<� H
�"���]�]�]1��"�Ǖw{������.�N�����mֈ�O6�@�9�j����6�D��.�l[;R2I*��O!a�,���H��PD�U;8y��;6�+��{�m.��3s�͇.�\|�K��z�"Q뗶��1s%���YV����Y�4��w-��z��7�C���>V|r�K~&���C�:{�y?��m���*���^�QDw�sf�|��#�Vdչ�UoQW.�ȶ�H�dxπ�c7G���6���K�n(e�Y�{q_��Դ���7V2����]�����MYޯ>�x>P��Ӷ¹j������0��dQ��ׯ9��j��Xb��ӏt�2����izk�w��:���%ĽU%8so.\���7� � s�����CM�CU�e�ç���Z6��zN�Ҽj6����E&���.�%k�O�0�D�>�}U�=�~���ߍ��A������CgC���ǅӝ'Zq���'=�x��^�Pח
��c���r�z��n�z�!q�ͺÐ�='�z`^��E��f�H�X���̝�����ܣ|���P/ent���2U=������)؅�Z/���i���r�ޟT+�X�lw�֮��a�u�*��S��� k�r�g�)י�د^�����kSQ��S��]תx��������'��M�L{"����&t�Ѯ�����fẄ�}�o�#�� �Mf^p�����g2�7*[r�Pcm�gn	C2n�uf���0Q���C��S�CdVk���>�[Ѭ��hƘ�o�dY7ڏ`<�܈Łr�hj��lYx��"ͷ���g^���[����b�6K9,�dq
9C7���]*B�ʳ�Y��w���t�W��%��@F)�$�1�^����޼sǒ�P&��uI���>�%��q��s[��8%��z�AwP%P����e/J�Z_���,�X�/b�X��~�4b�z�;�'J����~��d@��@N̠$�/�#�6�E�E���X��RH/j3�|}q��1n��2��z�{}q<n=v�+�2|^ʞ�ި�tz�O�W�����ҿ��}@>��[yD!���r{��<g��{ޮ��g�)S�q��+0�56e���,|���g+Fq qjB~\���ƾ�����oԁ�x֏��m�_�3����N��ɶ�`��j�����:��� �U_�~����x^���uˮ��4�H�U�K���z5g7sgɓ'Ѽ��}�Z}ޡ�R�`���v�ǳ��ê^SN��z��co��$���H�b��z��>������7�7�O��^�ޑ��e5��TyG(>榝���)�d�Nߨ�y��zc�}�o�Pk��p��L���1�W�+���Ζ��f���e��:]��/�w)/<
iݶ�����r��3�?����=�#/x:��}�@�Q[���و&�`9}XSڕ�-$��Pȥ	��iG#�f��O�أ�IK�u��7Ky�L�ɖڊ�N�rB�-8�jW��ãVr&��w�i�lzo�'|����������S�cC6��^���Īw��o��w����|lo?f�����S��I�\�g�';��4wj�Ui�>d��`	��W�S<��S��ey�F���<9v`����T�z����q'�f�+�z�=oM�Qp<�ƗTk�'�K�BĤx����H�׽�����]�f��݈\ku�Pϭ�K/"V��2�\TϔĲ��^*��\���5�mb��֠.��@�'s�E�N��߫�q�]j/��~u ���T���J�0O˽�m�Y�ڒ+�9��\j��P��~��������Q��,���'���;��I��wp�^gFvy�sۧ��g�n*g�<��	�OՃ�#���Q����HN����ǲmK%X�.]y�:'�ތ�r�����>0.�f:�m L��2��s
�R��m4{a���>�L��U�ԩ��Ϧ���^ w�+���鵲@^�����G�:
���CS�H�3�|�����H�D����ԁ^@�<�r:��[5q���/]O����ꉩ��|+>��٢a�鉶xJ_O
vjSr.�����"�Ivy�J�P�]�a�C�D��"̦fbݡ�*+�tD�;�&L�aݾ��}K�z�ҧ�}^t�`�r����OR��k`���7�5s�5(LJkT,H�B�vgk�f^lj1�1�����,�\�w�\��bk����)J�^h�L�O�G�wĿ	�5��ƅ˪���UT����{Ƅ���ľ^�[����ݯyU��>��IϪ���O�|s�>��bc#}�8@������UR<�Ȍ�c��!1�E^u��]�Y���Et���᛾��܋�N��}��7ɛ���2`mw���moN���%�ko��ٶg����]�w�un���ﺘ�Q�tť�9��P��=V==9�M<�TMdn[�~Q�[�,�?W}5�K������\VW��zN�F�S�����/��>m�k���6_�_P�S�x%����� ������*���t�p7=��wq����{�w��=<��z�����s����x=��gF���<{>uDe�����r����V�s��Y��6=`{=��u�02"W���O��7�=�Zb�7Ϯ��rKk��ѷ �>��Ĳ�w��ݐe���k��w�>���ϯf�W��	�M{"eϟ��W��Au���ڤT[�$��f�]9�����,���Z}�V���g�o� 'mHA\o��B�i��D{��,��G"^Rk�]r����U4f-X�ճ��T��q ⬼���R(�Ne����wW��š��W���T���Pv�d�+Sڱ%���Er�]����m�:����3�N*���)�A�z��>���:E�gf��$�b赐U���s+��2dӆ ��l�����H�/c���G���Y�I���N*� �v�|9�\��;�p�KS���|k>�'��o��t_O�o�_�m�X:vK��@Nn$�& b�5�ٿ����j�Ӯ����{?O�%k���>�S>^��\{}r7�4ˏ��8�O��@���&}/��z�OS���f��>����]��^���z��b=�\O�����\�gW���b@S�#O8�(Υ��ԯ�q}������!�^�gʏ��L{�����I���\�7��]i�2���^�z�+�=qԊ��d�V��r�\�oԉ�����Ɓ_?g�	�zU�5fr��{�Y:��_y��kM�# �V3�}�mC�Q��b����'^o޿��"�V�h\MX1rsh�SݣgW��p�|�6�Ru���M��=6=uպo�/G���ս���n�l��k\H/Z��r7�'�ٟ���߽���>cM�}�Q�|n|@�����hۊ���ҼW�.O�.q�J[���#:2}����w�o��'������g���A���$-�����ǅ��@��96-�\&�7{Ǵ辳�-ָ���j��ҸRw^L�o-�Yk���;>,�\�c������Ћr	Mj�B��l%���#�ٲn&8铻1u-Z܂��F�I�C��5w�-��AKkD+"�Y����2f'z�]�&�sa;zܘ%�KL+�����H�=��/.�/_x�zk�-�^/}�u�>~���=0-g���s��ۙ��k�z���sZo���+g�o�������O}9���)؅�Z.#}���?�W��q��{�GQ��y`O�u�0�������{^ -r|����������^ڽ`;t��dZww��z7�����t�n$�5�r���&_�3�]+]K30kO{&{��ї�2�i!D8��]H,�{h^�]%����]��1L<����.�ԙϬ�.:�n����/�roz�ۂ}bw�������\{��ݎk|}�:pK/T�-@L@�@���<�&��Z�N-������6���ё�޶��IҮ=��v߮�c��3���H	�@<�egY��EGzw�yM%�� x�����=����æ�s��;}�\O����v�*�������=���:痢��b����}�O���o(�7�~V�9=���<4��{��;�}�0��]�����Mz+��Z���h�ㄎ#萿˗�ן��|sA�ot����\�MJB_�a`eRiW��j`�6��ɵ/mA�!�{aRe{����'���E|����ѻ�Պ���Y���N�u��Z6���#0cՂL���'Aw��P.�ko"�l2Յ�YKM��ZM�8Զ���j[���؋�(]��%��e�f�&�e�>C�߫��S�~��|�rI{�%�ǣ�;k�:�֟i��a�+���t\^Uj���V�"�Y�)>��H�7ޠ;��h�F/VQ�Uu>*8�ߥ�iџS�h�'��\�׆�ږzw7G�}�uz�ܘ���I����_}lm��1�S�e���_v��V1�{��^<[��ޟ6P�t���ck�ګ�U���ޡꛌ�ߌ�}�\W�������2tΡ�=��Ո��֡7��	za�KG�΃�LxW�]L_ҩރ����ȟ&>Qf��G�j�7�-o��~�F��盛8��������[������� '��W��J��FB�c|v���wj��+���u���^��5�mϛ��ò?Un�T�ح��!��=\Q����c��]��3�{�D���R����f�7؅Ʒ]E��Բ�V��2�]L�L_��58�a���ة�����y�t�����(��~�ⶽ�X]j/���?�ͅP��{���u�kC��M�DUN��"̄�5�X����½�|u}�;�v|]j0�vԳ?K�}�X,��g{h�@�ï'�ٳ�]��;�p�bVV�bu:��ƈ����L��n�nv���J$����y��)�{ȭ��>Co�Z�Xj�b�m���_'��N��f��oW8��W�7Hs��i̚��ׄ!Ʒ)"��aE�K�����GW�|{���+����@/�E���e�싫	����^���{�'�W���6�~���6c��7��9�qkti����Γ���(}�A��n�P|j�-�K��Y-P�Do��)sO��ҮT�s��������_�;ȁ����/�vA�ܨv�֑�G��[>�m��TogTKNΟk+���޹��uU%��z�|�	H}Q$���] ���7����ڮ�[�(��G��3��|��ϣ�;�^}�ZC�g��]W�ڪ�`���s�VO��3�W������5��Q�$z��]ɋ�����}���FǽG��W��*���2/yB�]����	�2Nnw�t�7�����g�/M���\B�C�>����V��!��9��c��ŨiIeK2}r��'�º��7��ݑ�Ɗںb�/U�ϵz���z�zzM����j����T=���6�Ӝ���<Fd�VW��QzN��+��k���7����sܧ�7���w�Z>J��[걾��I��� t�Da��"����^'MƗ���"a��V�sD�p鿽aA`�#mLˬ�|�؇sѬpCF��"gr���]�+{��F퍱��u.�:��OQ<b��=�����-��A���șN�=�6��{@�WC���Z4�Jw�5����' ˾J�YH�è���T�#�bw��Ҿ�R�S{vt��Y>���pA���~?|��N�^��W�h��5��dc��������Y��FN?W%��喐���>T��}�"S������i��>�G-��lzpg�>�>vhM�N����pz��7^�ʽ�W� �׮'��y�V�z�y8�tC��{��؟zI~��ԟ7��r>�%��1|hϫ��|��9;ڐ����b�k4�k#�Lyz��q��ǌ{��\�+}��`�G�ͧ.I`-L9���3�\��|���KS��L��Yt`�OxA��1����5ԇg���=��d����	��b�1��2��Ȼ�8������+M�x|�:����\{}r6�ul��ztO��w�L��=�/LN�P��t�d����ZHy�Dw���N�1�w��}��J����z�w~4.]Qf����b@[Qe�oÕ[W�{K��J2=<�Y��Q�D:Kւ�Q�zg|M�޸���=qW.k�c�ބ���^���yG�]�A�n�.�����U�Y����2�>|������w���Ǖ�flcm������lcm�\������m��61��L����81�������6�����m�����61��L����lcm`��6ތ�����cco����m��61��L����pcco��{���m��b��L���!Z��� � ���fO� Ăw�|�U-�mmV�-m�lն��J�ƶ�l�kj[w9.f�n�nó6�+l����]9[j��e�F��m�6�M�`ŭSk,�5h�ۻ����S�y���N�2e;�ݮ�Ws��.wrܢ�]�ҕ��kuݬkm�V�gY�jW1�ή���r�۲��5�=u�n왷f�\�������[��٦^wv��ݹ�S%�j���ݴ�;m;��֛[�u�ն��gm�]���v�ɳnZ��ۻug���m]�Wd�Z�i�3���M���*�vw]nw5�l���;�q�n7�;�n���EWx  uT�q�}j׼ު��=稨�=��ۺ����W��^��s�V���ׯ=:�خ�U�=�p�^����;v];fݦ��k���;l�ګ���  ��T���a�
+�����+�  ��}Ͼ(�Ѣ�(���^�E� �.�}�(�Ehѣ}^�����(��(���۟|
@ 
������E^|��\6��_v�5u���[n�V�eZ�{�  }�*��Z�b�UF�wqv�Gvn�:�Z']s��:���ۚP��������
�/s��]�3������8 �:��*ټg6Nݴ��۱ӚgMo� 7>��E5%N�^�a�U�;ѣ��4k�y�^¨&z�YQ/n�wi�[UJ��Ǟ���4�����5j�VS��x4��ӭovn��A��zO)ZcMO]���k�q]6���| �}�Jj�c�Q����w��6� 69n�l��/]ӭ/n��O]���Tsn����S/@�9ס�j��{{��A�Z����{{�g�����ۗm���V뚑4;H�w� ���t�Aj=��=.�^��Mν�����w���lomڽ����m�Mu��g�n��E�7�ݶ�� ����[jJ����5��gz�����2��okn����*�k��@����o6� �|
t:}k5��C@�q^w��m7mܸ�C�m���uS�j��ݼ�Wj�Z(Nu8H�3J���yPoo7zY��h����ԺӬ�\�m&f��m��v�wuj7v� ��� �/{�z��ZƔ���޴���u<W��=h47�gy��v�(sf�����TN����V�m��g�5,��{���h�Ҍ�wf�u�n����ݺvj�,�c��  -�㮻i;c]nw����Vڛ��΀���k]����@���]v�Joy��*hv�7tҕ��Um�R��n��a�����z�����@��=u�w\�َ룺��;wb����   =��iD�ʔ�u�҂e�v���� �oI�]I�U[��
�5��PU��G
�M�Wt*�u۶�t�U:��'�S�2�)P  E=�	)J@  M�T�M1  S�A*T   5S�I�R�@  �M�R` b/������?�2�iw���)���m�>��<�����խy����$Wz�$WJ"�4W� ����D��" (��������k���w���c�+4��e�����N$�� (cEE��z7IB�#Vwk���)���v1%����	]�M[�뫳;W��7f�F.
���� � �w��򦩀b��F`̱�M�Bp���(n'U��L[7C��0�H���e��x�Ն���sp,'X���SR#�l���%626�GK[������}��j�YZ����_LQ&�q@�ݰ���W*�%!X�, �{Z��jIZ��#q�SGa�ҟ�{<35�X���d:��ap��y.B-9<����f��.hA�pՂ2��L�;ک�Z�����Qc#"����t��#�<[�����v��-'��j\�����s;�@s
��6hH�qiYB%qaú�^�5�q��<hQCgȩ�J.F�@q�%<�4�-K��eMڑX%��.V�J�3�	�Xr+ˎ�tn!�S=&A��:g��6Zcic{���s�u����/F�P'z/	#7 Y0Mq8"Xm�c��OREM>��䬭�0�|�ؒ��w�Q� �"�j�����\�2��̳.��XN�<h�,u;�<N��>�����-KY-]+���&�">H���!�Ԡ6i�5�^풥	n������1
�e�b���-Q[X�4���KQ�[�[4-D�*�(��ZΚ��kF�,�0
.�;�"81�6���V=.nk�*|����,��b�l��D]�K!�ѕzhE��޹���n��-�0K��y>q	Y"2��cm��@��z�v�>
�4<i��7EXWI����:����MZ�2Rz����S�;X�{J���_��p�*l^;r���e���B�f�g\4C��E55�Y,�{���R�a��JnJO/lR[%h�UEQ��)�,��l1�6�Y;Yww����iX�U�`܂�&lT�+q�L,-vVn�'H���e��(l�~'n�e�%�!�]m��#���˻rKT(T���z&ʁZ.f���mu����N��mT����� T�Q��cP&��A҉mm�:
����7v(�Of1 5*�̊&�����`p�Z�[N�hKЙ�x���@���xn�$��|<6B��y@��FE��̻��Qb�TIJ��d1VƆ��B�T?[JQ�n;*!��TDbF^ܒ�v �Ź�rj�)ϕ'�3IQ(�� �%�f�pE�E�X�����d�^;�5���:�Ң�������wDR��gd� ӀC���nA���c_Tti��@�t�JO�dfB��:��Ӊ�=KIQ��῁�N~��*�&(1�Ԩאg�qje
nM*�B��WLV'52��X��x^�W)��Dk%�۰���An�R`��y�soqz¢�5��L��м!Cv�Q/Y{e�FȐ������]'*7bP�dL�N !N�E1�Z��[FM
���p���,�����XΠ�V&҄����rb;��3Q���(�~���ņ{����]�t��̣؈"Р��ۦ�\��1KSc{g ͳQ���tV�wW�hM�r��������v�بm�R9�j��Zw��q� �pl�	�H~�cso��͘�ګ���F��@��C��]  ��v]�]-�ܒ����ݦ7�<f#!'3nݍg�;0�cuT�����`�n
Y��;��Mݡ+vc���1:�[!P+m�jF��=���N�&J3'��$F��h
�ˏXn�ݟ#J�m�d-���ML��Y�Y�y�i�$݈Hn��V�[Ī�֢��bQU�Y�-^46�ش]�5a���}�n �WY.%H�H\C
]!l:��B>���Vn��3&��U�7��]c0w�CL�{R�����|6��{7�S�h�7�DK"�Zg�����-뻄0f,��/�n��<Jr�Y�,<!̨��2�_�KQ�G��ȶR��n
�īQ�f�fm�BBݓR��6��i��&Ի�a��j��"Ɗ4H�Y�5 -�t��T4!VR�⹓^"�vn��X��V�P���%��5b�(]�NQ��hn˘�'p4�ʽrm�KF�2�e��0�P�$��QZ�P�%,R�	ɡ	u"�}��?m-3&������4����X�ӗdtZ�6����Hۘ&�+d	��+R��; �1�1G%��Ve]Q�B����&�0O,�F]>��>��A��ـ�y���Z���,�|XS��U��p[F��U<��S�[D�{!��ʂ���*ܩ/�Ŋ�{tD��qюnJF��Z¥vJyAf�1����N��t�c������ܪ�qÕ���Ւ)|s�t,AR�ë̲$-�tb��q!��hW$N�)R�6�f齢��t���FUDjj��+]�����b˖Y��"^�����Z�ҧ��ݎ\T_a�*��k1�d��Rʧ:��JX64eI�Xkj��:����M���zB�)�hAڭUtq�6rc#hc�����A*x�kJ�cI����d��Z�"e[Pb�Y��k5eՊ�a��I��,E,)���C)��T�6�ӌ-Ot�lL�sr��D�U��$�:�qR�p��Xb���áe�VGK�Ҫ-.m��^n�����)�7,Yͫ/@�D�
YhnGt�y�X�aa�u�]�.R��E���Yj�5*�J����d�ӦnJ������`��i�6��x���g�{th�B�%6���k�m��+Ń*��jF����5&%z��S����)9f;�e=K�B�6����F=>8���mOZȆOH�;M��Ě&:^�p��� �e)�u%�nh��ЭJ�O
�*��6Ցێ�clT6��!L�Y���D	W�Z[w��
t�k�z[N��Ӳj��+q� �]Ök�Ŕ�()/�!��N�C���	y��n��y�'D�}Ö'R��fPxЪ8���Ԩi%����So�Q���I����������V(%e���7�\�W2 <��&a�F�j��ZU!�����Ne�t�ʅ�՚�>�"�;��(��Z���k�bv.�`�ǖ�U�N��MnK�Pn<R:F-����K�.0�͛l+V�D��{E݉��U4���uS�2s6���]%ǋc�Xj|��nk��/��X)	rJe���fV���a~���	�15�Gh̠�X�bdc{r�ɲ�ܔ��EB��^R��*����+�T����hE�-h���0=J�iJYEd�neYӑm�[B��PDZ�h�U�y�;�8��	��y��u��ǔr�i¡�{��c[�h-��)Jtb]�O���Ք4ARե�6����$�^��f��2���%����|V�*�\�ӮVk��C�k)�+p�����@#r	yx��I"�QpG#F��Z��9E�؄ݭ)��sB�r�lAB�Ɇf�l���vZ��6G�kIb+q�z+1���$�n!aDФ�t�A����.]!j#Py%�YW��#Azw!��V�xwL�H҄-��X�P9�2���-��(�Uh���M�����&)�F�5�Pyb�ګ���l�謏+�qҦ�a�Wn�bք�PV�K���T���&Dt���m�&�z��nR���E[)��6�Xv�tڍ�H������ٔ1k�u��Wu��`�$��ctt@6P�*yuxp�"b�<H.F_��طِnV���S�0��˚@"d׋^�E��������^�O&(�$ 3Rݬ�X�P�w�hͦE Ӭa&�Qj&�	H ���Y�M�O1朢�NS-
&���jù7v�b�:K*]���,��ܸ�:b�B)GFV�qQ��Y�*ht�)�u4en�Z�cL�
 �X�PX��Օd�r�����Z0�A�0��8^x_H.�ۂ=X}�w� ��Q��*ʞWw=��U�J�V�t��bfk'	l�u&R8�\�36�=�:]2&��v�C��nQ8��P�F�)Yon��!��
4�ӎ����h��ً)na���`�ն��>��%�fIJ�]�b4�V�b�k
7�G���,�t&n�⦵ΰ��;F�W�+�ْS��]M�D�����"�L�B�0E�1&��2U�4���2�B�a�Sd��ϐI��Vwx������0v-��L�ùJ-;rA��
��*D\X�7�{@�P���wdFC�M��e�GأA�Du/z=6Q�h�332IhI��z�*�FS�#�ʶ���CX�u��^��		���b��b��P���n�a�l�j'EL��wճ����s�pX{n�T/t��I6���7�u��0S�VZm`vt[\�p�*�Y�tb;�l`I4�QKC/�r�bpZ��n[2���@)�2؞�h֛D�7�qjY�݈k���wW�2�i��۶��b"�T��,SD9z��$Tf�K�یl�B������EF��Rѻ�TS�	�y@��:*�]E���=[k�e]�RLa�07�]n�a��$5n,��Z6�"�u>���M�y�G�Of�K`y��+�n�n���C�c����=�4���*b:��$Vj��@%��R 7�U�E��je[V�uLn-�4��*��`K ����勫�Xc�tQ�����t�[Y-)�v�%�C%E�nٽ�̀V4$�D|O���mOJ�a��u3
ʬ�D�#���0g��=>>.m7��w71ib�Re�4�]XBĵ(�y�%X��&��.�݂�Ů��M�֊�e<�[r���i-1)g֚0�cKͼ�d���7���[Rʶ�&�Y�눵��p-5�����"\[Mf���5�¥b%4�ۛS^k7��'f�!�%m�g�r�7�A��+V�&ئ�)�`�C-��Җ�I�LL`x5��ݔ�
�	x�����������*M�����n�ysU���K���C��r��ߦ*��vm�/Iil�9rG.l&��t.dR�Q%�����ˈhA���!��aV�Ƙ�t�V����^#sIW�B�ԓ���FW`��G�����Q���%7���7D�,�Go��h�kE;sڴ��P���=;w��k��af={�n:�� 00ݝmmec���*���T��lc]�����M>�f!v�W��0үF��p�&��U��*J�����V鲦�r�lk)�]�K&(r�ܲ�v Mp�u<�p�QY&I}��!j���Y5bKI����䡷��\��z�S�?��)U�a横��de���K�_i��.��c��=�+V��u8�5)hMiZ��VmJ¢!�LB�Ef�⒰>��ˤ�(v�~�b�m�EB��{��E��7B�ff�7(K�f��HD��#��g6�I��M4���1�m�4��"v(�t�/S�Fع��ѫ1�l$mfYv6�*֕T�yJ�#m�1M�$�hxE�aiz��q�f1�ck^k�t&`��{�Q�bYi��*]@
��3ؖl�;5�������ܧ�,���Z�-���FZ}j�W�
|o�;��L�<ֈ[�����u���sa�yE4J)E�D�eLiU�WsYi�RZ0�"�0�)�8���0����˴�i�v�hȚL�T�"AQ뉊�����)�I��U���(ek���	���Y�[2����A�����Ŧ���
� W%���7���K)�n<��h�1��3PY�Xϥ�B��6
�'�� ���J�rk�ކR���j^�Bf�&���`Tާ� �s�j��{w��[,�صd�
YY�"�^�SQ�b���4��X��@�ǰ�zf}�l�5%�V:#n�!suXh$hM�>�v�Rl���7nf�jT�	���٫�RD�c��ɞ�i�o��B��&�+�c��S�廡\[�:���nX.�8N��>�N�7*�GpQ&��B�MW����&ҫ�w�	"3,
ı��j�g3қb�.��l^��Ұn+3j�;0^��,s0�q�b�6�jK�������b�+TU�E^��O6�~��
�k�eð�=0iaۅ�W��L�s�^�YQ�s�^������H��!7I�\[}Zo������V��Xz&j��m!(k�Z2GDC�T�[gA^�(�wф�JR����03��l�F�
�(�I�뉵�J�'�Y��ӏ$M�g"�z�;��v�E2(�!V�Kh�2`P<�`GtTY+	�^�`�/r�O���������nh�L�-����n�g([�cmQ�@`0���7�\H���㕷[���@/i��P�_Kn�VnR	K����� zMj�;Q�Tumbw�l�f\�ܩ�*���e�Q�ǻ�CwM��lU
U�����v�D�ّ �8�m�G��o,kE��J]n�	Q��h�e۳�ݜ���y[r幩:�nwPP�U��B��@�J����)Ә�~n���0���9ow�J���c�l5���Jl/kkӲ�ڡ�����'n͊�q�e���>m��[���~S7�t��OGqMYb�vi�wU�{��`X]��"�̪�n�J<B��A�L��Ѻ��yi����Щ����p��0p=;q`��#�=�&�h�!M��pFJm�Je����2񌧛0*��:��L"�MҰ�<����*��8v����3)���m�X+En#��u0�=�ӆ�]�pK���ﳺ��ۻ�B�X���R�J$N����R�^Vg��[�{�_
p�̵���z=��o��e�-�
��X���7���|�6y��
A��k����:x���Vy�J�������p|f��p�PzV9�w��pcq��Ξ��|ۓn�T0�$CNx���W�aZ/|x��L�ە�紾�|2j7H
W7���i���d�އ�O�5g���L�~�v�:�p��뛙�(Ȧ��ٯ�ݰj��&��:��{�D{�)�+!��#9f8x��%�7�|���a�Q��Nܥ���V:i�"r���5t���j(��HL����G��Uo�����t�O4q��N�R�f�Q%��Q3���N��4�c-m��|�EJ��F�!�"�m�$���wR�E�SwVMĹ����Bn����VѦ�KY�!C:4�X7pj���C��c	�%,)���z�-�D {�,ĥ'4���9��H�Zs����kK#j���l^{o7� Θ�0��{vp���᳷h���;��ãN�=C8h�Vush�;�!�0¬� ����ǲ��Qv��+ֲ��
c:ݍ�S��JW9ڦ�mY�1�h����3.e@°L@6�:�$�2�I��7=N�I�>�t.������-p�LAe�=ϙ��*(���fd�����i�N���o���-^�Bl�]/C�Tqe����R�dw��i��՛aB���M�v4��vw�w}]e뻠�`��b����isp��r�m�WY���E��N����{{aa�ɖ�����kx] ݛ�p�,�<��*k�aݥi;����py(���,B�p{;F°'l�6ӭ\v�e�L[����%�
:@R���Y��m�Sr�=:o����k���1+�O�Z���{�͇��#�5��^�gi78����i<��j�qO6��U���5Ly��;��v.�A}J�Ɩ�;�q|���Y{�) �L���'>ˎ�";~�}fF�����G��B�&�!����N�Ln�oC��`�L�ɣc���k��1ן6΃q��݇!��	�n�0��no�T%�\d��'8y��a�Rf�}y<²�3	�l��hyqg %����r�����zIX�ػ�G�n�q^�x)�6�JG`��}���W�a4=��	XW�b�PV�U_Ɏ�s���j���˦���S�����B���<$~��|�ы=H%b�w���6�@ozg�	a�)�o
Oj�G��l*خ�&����m�%��{�B����<�����1�#_
�T't������\/�m�����"�2;�Z� �N86듃�6�?>]�u �0\�`�[��<����fK��I���''I)�	y�;HQ��P����^�"=�p��Z�[0�4ќ�9����K�%��x�w@�vR��c�n-G.һj'���r�{&1����`�
�Am��ݥ �u����c�<(�KB^�}��є�H��%�s#7�"��nt%���_�ԭ�C����acy�j��$v4ޤ�6O$��>���+1���Y#�oZ�@��Z]��O%ww�����aÔ���G�7�qq=�v�Y,���+=�X�J��B��P����v�k}����"L'E7���X��ᝓ���Y=ґ�&�<7U^��	�q�W�7�<c}��ޑ-��[/�����{�R���FҹO^R�ePgYo�[2L���7�.�\���G���Uk�bh����6��o�E���<3e��j=1�a=�N?���fz�f���S�77�i8�OT>�TBxM�P�_��;��wx�����r���o�zb�K�:�^ۆt�����b��ɧm�r�R�c��m����S��Rd.��u��>q3g�����,wL��뷒�T7�5\X��ҥ�2u��Z�����K�H���Ti�]�{/�q�g�7��E�=6U̗�|�Q���kk�D����Э�n\�O�g-�W�2�f��2�;p(�#rlX�����}�á�Kg�D��4iX�3y�T���1C�We;�(��ZtQ���ù�,C��Ua��M���BE�{�4/�.k���Q��1o��g9�����FHt���J�`̞��p�f���Uά,f�7(]!�)�\��m\,h�[�k2�7��TR�;�i��]V2�a���Go{wKx~���V�Ԇ�,��f�[�w(�a-|Q���1`��̽�{|O�L�.�ޡ�Ţ>��)l4,M�o3E�J��&�v�$�N���h\���$'��
�����n83˯�&��2/M܋���ۖWl񏸂�d#WZ_���l`[�L���_�w*��u����\V���ʅ��{�~yA�ކ�e'�l����E�e��)�۬H��G�a�l'�%���c;� 6�oE��Q�غZ/�M��ݳ/9MWN��1yo��G��^���-�|wSr͠N�:d�?3x�t�N:�c6�m▆�tX2�r�/��G�;F�qk7�":���t��.��wP�׏SA>9�7y
�2Sߧ=޳\ف��~~m�"R�nruoW��&)佲�9iE�7ah�M8$s�l�_e	���0:��H��9�3I<���{�z*1��N��v��q����ҁJV��f�Q��*��#S�s"[|p�5�b��l�k�:L>&=���!<�o���_?\�^/B��u2C
v���ׅ7��\��4r#Bj��ٱl��{F)�ʯAԹ�PK+�[��=�b��PJ�wr�Ě��= 2�۔�x�yd;kgqn[|8�Bp��-��m��*}�y�tn.쫆��%CX�y..��r�B�ק���1v�ѭ�`(#u�#�СF�����XfCi���u�mP�����d�I���(֬s�1}8N������O�Q���Sw�������h����f��_��*P��Yf���|��Z9s� C�{���:��,�kq�w���7�%��gz�^[ӿR��Z�����(Sk#T>=J�+�+��Eo8�ʽF��kDZ/0��8s�]�"y2d$���n*P�!���@J.���Cx�^%���}�zG\q]b�4�Ibe����	��XNH���^�.1���v���;Ö��\���C�D�o���Z�N�+�=>�G`��|(w1V�M�I\�v���>#58׶x��,�&hs%��ѭ��6�L��G@��ܳ�y'mH������Z(�_Y��;�B�G9W[�Ât���j�M#�� u���#y�H��ܶ%����}���ջ.�Dvǀ��$�e<hz��֘�m�@Ƨ)���Tt��ͷ���,@&�/�]M>V7���cHxe�5y��̩Wd�Q��p�����Q�wC��a%�__B����{}�m��W�p8����_{��ؽ0F{݊��k[
y7r��doh
�����P5���Iݍ��H�����fv�gn��;P�/B�c&�>b&ޖ%�� l-�g��u��M�\�^mSZ�u�[��V,G˨g��;.D�1������!������*��^u�}�M�K��.��}K�47�wD5����Aw^�(�N�+e��A׊ΎFS��7t�Uu�cP2vα���[ܧ׷-dg[�T������1�`E�s��v8-4�Er�l�,j`쮨��f�Zs�FI�Sm�]���ws��)#�G�*�Y�`� ˲�6�������Iq꼳��q�R(܅���#� Po���o�eA���+��-��OQwB�f�@B4Ӻ�[I�z�Y���!Ǩ���ġڧ�<�9I�kmn��7��Q�1.�}���eԻ=;�p[��r�}�������LLj�nMč�y;���L�|��	��~y�h�9��ɏl�,��bE��hA?Aݮ�wy��<UoGXOl�du�n�Ccږx�9R�����"ȯh�A(ƍ��f���]3��s&s�֞�]a;��WG#���K�Aڤ�� �iv�J|%Em�AP)��*�q���oz�L�e���{'��̟D���cu�p�5f�U���Q7S�����ǗW@�5�W�F�-6�6�ǖӘ�����g�����T�5.�m�)��tS�8�Z.$<C}b��/:�x��k=�
�����s�9��-ZU	��f��	��(	�c�|��A�Pܬ�׈z��j8�چ�d�8wX�U��l��QiJ�[�dꝻy��;��=�._j���xy�)�ccJY��̚^��q�p:ͩ�+�mo%"��e�G'^L����M��yD�Þ]Ĭ�]i��H&��ti��y��H���:7���t�k��/����/+x��{WJ�Ss��{;O��׮�f�Z�%�v(}{�|�R���'5,�ɣb���S�h�����\��0��.o�83/&=ǧ�Bc�(╷��SLU�un�1p�ӄ�E������U����n��.�Z�Y�w�{�;��r�,�v$�p��3ٌH�x�*A�6{R�`�h�����Z���E�Yc�i�(�,���~)����'s�	&�����=O���[/L��pm{��<v���@�ز����*���y�]�z2EJ�׼[k3hl����c�ʼ�U_]	P!�HM�p�R��n=u���7կ%k:������m�����륧N
V��3����1��� ���a/���4&s��T�ap�����gS����+kYW���r�>� =iޑ��YGD�չ��94n)��=����/�O��ޘ��Ƿ(������w�My��諍��<xiX���ß����t"���q��o�^d�+nD�:#'2`��3Ie�Ȥ���^oA�{�o0"�q{J���n':�^Q��tX�_+��*n�J����W^;�:c�}��d��@��@Zʙ91�=��3����+^Ʀ^���]NKkI��m�{�y �-�ʑ�G�/�w�t��g?�WW��;� ,�p����.�J���Us�r� 'kP_;�Q��z�A��@r��N]`ˇr-��e��[m�'I���#ߍ~�-j�\ܦU�_+��6E��%��'
z	�.b)sJ�ł�є�K��������f_	@�#-i�q�wh7�!�c�`mJ͌�D����{�)xb��⛗]�q�R���jJ�*]f�M�N��{u3���:��t�"N'���<�-��/E6��gfb<!8؎��k�=K��6r�(j�MY�$�)�^��цl�+�<��۷��ZqF*n�����	��\y*�̮���ӇiW����l��6nM����%!�k��Щ�_j��w3{��VR<���h5��2�:��h�N�};p��b�_e MCL�&ˈ�����-�3���:�6�C�n�[��j���u�ӣD��q�p��I��Я����+<��Ÿ�}*Y��Q 'Ԑ`Kw��/��r)�(ut�+�Q#�FmZ�.�Cxg&y��*M�u��\	���Z�	;��I��X�#R���z�%����8]ZY��0y������������@��l�X<�
y�8׼	9Z 1�</�;�
�RDw��WTW�;z�$��{�����k	�ɥ��At�����fe]�=�^Oh�d�|S�-ir�Tq*�VrZ�m�h8w:�%��TM*[�6{3N����z�+QM�(|�͑P��-r�.Y��ʺ�+�йw��z�A�Dq�B���v�>��\��')帎���:���!W�^��rާ�g-��1��|]��6���Y5�f�m�Jb7zˀ� �>V񄗓ʢU��L$�R�M:�+�0o޻�µb�E�BS�*��2=��})x(^��m��}���p:ɕ\�{�A�H�h*�W6��L���I������)-K� *��|���i#�t�2w��L�����Щ_sԻМD�PØ@�I��z$͚.n�6`\�V\�#ơ!�O�5>��%G#8N%:���}$]ט� �!b�ʂ���Mm��d��t�6Ed��d�}�QQÐ&8���.�i�9Qwq�PD.�՛0��b�$���A;�Y���B:�ocb�d;���nY*kZ7���<�����*���oK�Yc�����l�ν;N�`�������&���Qv�h���o��u����b��[�!�c��	��:�ټ����O�t���X�򓮂�Û>��v[O'jH��v1
��/�/6tw�����h�+rq�ՎU�s6#cs�)љ��M�Rm�G�/�{������&��i+u�x;c�r�
+Uŏys�t������Dn&��0�p4o����b�y�3��_uN�.���<��T� ���Fq�ջ������R�t��|�:���Ǒ�Wk���s�wPmof�Wӂ|m"�c��=�l� 9��W� 3���}��� ���%�3O.@�<�fEcjevRڝ��b9H�'Xv����[���9�7d���y���q��36.Q�Uǧ=���Q��k���Y��x�-I�J���a:Iԕ�ڽ�r���1��{�'c2l��:.�m�񓶼.W�}�fB;�&�l<(�W{u��5��9A.�$�X/J{f.<q1k6��X���l�4y����j�NAV��o�ӝ���[�o�0�k���ljQ���6�#G42�*kV����3r����������V��&���>h���!�7��,�4h;,�Ӝ�Sz��lg���-��J�u�3:f��>\��lZj�uYP>7���A��~�5��{����|> }���� >���}��<"����ݿ�����<�1e�����-����d'��o����J�YޫdV�w	��ʏ4�-�tye���en��Z��t��9۷��[�������1��2��1ͨ�f��^x^��Ko���x-@I��uc<o^I���<V�uX��ImKNk�7���`�Vsy�0^7�q)��3������vo�����/+��Gƃo�2Su�+q�-��p�}}���;�h<�R���S���Xtu�ӸŏTX��Ч���鵆���	�:ѹ[g��*E������������V�-]��.��F=aL�=b��AF��U)�.��s�̋ֵfֲri�F�`1��R���=�nS�^NR@��i���g=�ݝ���)7l3����L]7a8El/��:˭�i�ڗo'C�<6cY��C藐�8%��q��q��Gդuk�U�K�SbE\#N�NK��o߸�A�N�ܠ���!��G�˱��`��m�<�O_G��<\q�� �PW�i�I1Q���^<��\�1��Y�9}s(;%�QoK���Z�+�I�G0vz�p�E��ƻ�B��<
w��׶ٌa�ހ�����K�Z�޴����/F#���Tc�2�S
�Hn�;$����wr���vf%��e��sg ���,ugW�x�y�Jt�z���Ԭ{8]�*�m	ׅQ+=[�Z�5V�p�	��z�&�Zq�\E���`���Šx�P��S�<Ke��A�W� ��g7�G�=nH	=�ǣ>��Q憱y�VC�|��M���h�s ��Q�e���G�>�hȉ�4H�3W=�V��U�����V� C��]귝�Ҧ�t��tP;X�i�w�ǫ�/�Rs���:�ϕ�5�M���k����]5L��	Z�V�{kQ��VR�63�<�@��2����+gq�����Ni�m����zV�P㎅ʅ�E�r�N��^h�&k+:E��z������c�n��YX���޺�{J�T�eN��,�e�q��ɂ�w��Mu� D��
����z�^*]��6(M��R�HVp�F���]=z�+���n�=G�ԅҋ*A4oѨM�ٜDM�J�z�Sկ^�v�Q�i�q�=&�Ez�@�oM~L��:ٷ�[ �w7�����Eu�`���cCHЛ��}�R�Jo;�u5b�TgFֳ-�(;y:��������$_)�@DrAF5<�ޕ0\�=���ez'}+o,�1�V�Nm�!�f�W+J���A3�ώ'�3+J�RD���w#�h1��1�4P�:L���5v����}]ov���h
��÷��i��U�;}��V�zB�L�$&q��f�}q��Em}i��wy��jI���V_�^��x��#�e�Y<�O���<���I,���X�2��.
Xw���{e��˥p���#�t�1���m�o�囆�C�Y���Ӗb-�Cڛ���K�8`�d�ۋ*;�a��ǝ�ZR6�U�hf ���Y�NPs��+��4fmd`ҾT��q<!ૻ�e
�;[o�9S5,,5�o�����[��D�yU��[�<jl��S�ti��anǹ^Z�����PwYu�D�)y�#��~����ȱd���Sϝ���h���mXͺ�#fv�w(� �f��4��w����/�B�2VL<��G�g����&$��0TEV�)�M(e�d����*�r&�!7�ݫ[����.�9�M��3������ �aI�/��잾����xˋAp�@��nթ��0N
�S5\Nֈ����e���ƣ�,��I�Y�n[-���Yq^|+SAհ�E6�����nYaܴh��υ�6���@� 0{�o������cA���TsQa��Uud.�U���۰��i�f��peTp�� �e�V�-/�=&t�n���v�
_;����VZx���#��՝v��[�̬x]�Cf ����I]ս<;N�w��l���/�V-Z��G|��V���<�<����נ�}sdQ�����N3�a�q����9Y9�s�u���G냡�{9U�7|n�K�m��1�k�Fgڵ����3����K.7)�w���g�Ӻ%9��?6����l��{��s�8�Y*��Px����1�� y_+�)m�Kٜz,�:C��*[:�u[����'b��Ore�0�<���+��D]�WS��)��U��������ڷ�\o��t�+�u7ǚTJ�;��*�����:L�;�c#��]�0r���2�hm��Q�����w9Aa��bS��7s��w�#\ﺔ�$i	{SQ�s/o��@ĥ �+R[;Sk��s��p&�U�ql���ݝ�g��~P�����3�ܹ������{Q�ue�G��3���s���>wt�}E�{ٸ��:Dj��jo�]־�bU{!w$q��-�����tqf�tyNV.��N����]k��"��V�p�OD��k|��f�n<k���c֧�Y��Ff�e�㓨5rT���\�P��k'<y�2�y�������M��'V]*�m���t{"݉_k��L����T�W��{=����&Գ'.Y�7��b�r�U�WI��F��A��S
p|�������J��4vT�5C�lL���ӭ�y����!o lw`�m5zo.@lׯ�w�qtзtéI�����ʭ"��h,&��������� ���r*7'<�/Ç
�z�cp..dծ��)���"��R�8*u�з;|�����*�����#����NQ��Sw��ó�Cw�CP�^gq]��,��	�Y�Jҧ���M��`�/:��xª���Q=�C��;���..�t6�?X삐O-��t�w�	7���8����ȩ�f�؎�.��83i"�6��쾭��.�Z�l�ZA,jN[4����ՙj�i?��Ѐ��N��n�AK�ѹ�b�����z����᭍n���������%u�432�]]�1�\�R���+�x?4���P�ȏ��4j�q\���b�#�[v�,�M�f����a˱[�o�7i2q.�n��Q��$�F��=��l����RQ|��-��J�[��+8�a�FK������v)AEt��]wf���Z�n�Jt�<75h��t�S��⑨͇�����j_1iG�3;���' m���蛲�m��t������3I�%E�86��sB�Z��'"��7��eխZ��!b������6�lf����͢��v�v��)3�Ǩ%q���u;3�7ۙl�k� ��z�<��+%Z�O=��yǻ+��7�����M�B��
;�cP�Vn
�vz�7;�0e��l�t�7������Z{�k1l��3}sp��H�M�쾽�T�A0�[�uS�P�J�j��'���ҝB�_�z-�ѥZa��p��1P��{�^+�/��i��Y�V+��%��q��6�E|��9��g`̣��-c�A˷��\��:z.�����6ɕ���<���ҙ�IKLݲ�p�Znnʫ��J��n�Y��(ǈU�3QŊ�PW��W��M�Ie�?%��'���Y�IM���V�;�C�՚��i�pp]��u�z+�#��\������L�N䫑w���.1ga+���w���U���F�:Tќ�"���r���`]ܓ���`l�G+�}H�������.p���������E�PL^S�.�o�Wu�ݥ�mF�g��A`�';eg#4Y[I��kC�kU�-�*��}|���rOM�=}*{��'���4%�b�ܰt ^vY��.&����ګ�l*�I���#�F�����Zh�ځ��3�i5z�k4�]�+�ܒΥҫ�g�}���fK����^�*�ʨ�T�ݚ;;/4;+�=�}%K��,�|�����"]���oQr�y���|��Ѫ�}�n̫��LV����D�]�Qѡ�ht�o�A�0V�&VXq����NX��K�J��̠�9`4s:�e��WioQ�lΩ���ko��^󺆴�:��0t�"��2��ǧ��Z7� ���h�5����E�)u��ZݥÎ�\Ըv�"�4�w�Θ��P����zٜz�s��tD���$`�q��0l�8��y�1'Q�TK�ڒ<^����s�P��~�����W
*�z�w���/1��n+%g�oܐ�o[�pJ�n[��C���7��������ހ�u^V�`u���+��޹}����F�[F	M���j��k�e��R�u}|B�?h����){���9�[=%�]"m{r�7y��k �r�d L�s%n�(�d��q^*DD^�4��}kLBecMP�2��<^g��A���f��;v˒�G���e�q0G�۴�e��c�$��FYY��GH��}w����-=�fb�o���s%��G�1.��<s����f`>�)l���M�n�����}v\{&���%1-m<z+.L*��Ar{��ݘ��F7^Lŝ�8�3�Ix���y�ֈ��;t�)��O���6�7&1��ɥ�����`���s���f�r��XPu����∻nw<�Šƛ�/��`Q���$��V{Z��5}�\A3�V�ή^u����IU&�o�1��'��Ռ	FM@��Z�Ttoe�Ԭ�r�̥�Q`�S�4�&Vw
��+LY��]���2E�(�f�cI�e��qD�T��N�
.��א����3���������!�co��OU�A�.�9p0����{0˸���1�^Z�'���.�#pX:������uŪYc,]m����K��2�6`�/��%j���	>�*洞ؗ��J_)�s�[�{�_|	A>Y��ݡ[X���8]b�u��P�e)����ɚŽY�8?m�zo���>�WAwa���!��Ss��yS�r�D�D�
ں'$*u��z�0Gh�\�i5O=�����B�|f(ͫ�D;��7�6�R��;��ӄ����d�a�b��"�[�t����b�z�;��v����ɻ�Z.�ɞ=>,j}�>�S����y&�d��.E��H��ŷS���Zq]֍w�M_S���D�5�q�L��������g]�U`֧q����!Ў� C��4><�u�Eڽ���R�o���/>݈�)7�l�O^���w�өg�9x�hۼ���ȸ�j i�[���ef��ށ���-��-A��W�|��{��� v�W��M��<<OQ�G�.]q�%�hĻʥ��L�s١��lҼ�������r�v�oa�s��)��=7h�lc��:<5vz-�zq���Պ>|��R0��je�Q��>�����b}5��;��9�����:��}9�rF���ջF+BpOP����=+V�85:�UC\��6Uc��o,�J'�Y�)�e�Gb���X�pmG�C֞�1�9�)C\����{F�y[� 9'2�ȓͧ)�μ(H����R���-t�Y���NM�wk4�2�o-�ӝHۗ�?wo
��e����`�Z�mt4���K��>�C�:�T�|\Gkj�.�AN��]s^�g(�<��|{����n��Т
Z�8kB �[�Q�٢�ږ���
��9�ڼ�@	������5PJar�Ú����cƴ�z�J͝	�Gf�d���sY��ޭ��V��1ș�q�>����k����i��l����2�ׂ;W"����1v*��o�E�+c��[�l	ȟز����"���bN\���K�����8XzF�/�4�]�-1��;zҔ��8����F��	�p㺄�um�+�g)ͬ��1(��̾\g�vL.��]�����gp��u۽0(X=�b<����N�Iz�Y�DX{3^�Ⱦ�qS HecQ�ӛ�V%f0U&�����X�:�Kd��K��yb|.�gT�,~G�.Y6��*wiN�kv3�!��|�E��k|F���'�#���uFSy�&4Ik���)�u9ji�9Ad�o�54��YwD��1G�ѹM����FZ˺U�<�Ma�zø���I|J-��F��� V���þ�`q�E�]�kU�%��v��!�Gƍ�H�Ї;�mP��&_&nN��B׹{p�mG����U������i�
붍DŽd�|�A �/T��ἐE^�y1��5]A��"v��2��u.�7"6�L�}��>�We[}'0������ԧ4>�Q������ �@Ş���mĤ�<�q���.����a�T{��3Z�k�f�dvM�jס֑t�N�wP�p<b��-�Ⱦ14.�:n}i��d�v�b�:R�h��Z�o4��Tmvc�E���=��Ml�����D�!�����tu�phYz�������]Z.���&�v:	p��-�Fy.�=��e�!V��΃���d����,��hLXܳ�8�m�^�t廭�C塪��b�p]oV�Og��s�!�m��k�N0���u��e����S�6���4%�����M	p��d ��u4Fk��nՓ���<�w��Z�t���hn�m�␣����t:t7�W�#̃�����D;�����}��š)�}8��x6\|�E����'��ק%�MmK��j�үcC:� ��x�h�2Q��g�-]�mm��i�Zo����N���K����ai�v�N��M��g�.lY�i���zz�Lon&�eRG%'�w����:��u��_�AQ{ߺ7�������#�AS��uwloWd$3m�幃��sF�>�fU�bP����x��%�%aO����r>'V}�z<��r�|y�J�-��;<��ޕjef�7�]5��0>��Vdr��L�[�a�]kf�v�d˩s�� \�7��ɨ"Ӿ��]Y^�J��,']�{�����_���,���;}p7��Ooj(ޮ����[�E�����]�J��P�g`�7�d���*U�-wb!�ȥsgJB�?wc>͏x�U�=WK#� w=��8��B���log[�G'_1[��e�&�J]��Ӷ�!��-Cɐ�go�-�fw��Mc�GZ�Yb���m�~����j�a=���x)��_FK����w׆4��5�nN>v4M���g'�ox,�st+��:2L�BI5����cY�9�_���~񣆩�a�&;.�y#�]�[�P� 빆�W>��Gr�:�g�o�ޙ�bA��y�+to8&���:�ǎ#� �K�q2O?ae�ܙ.!�a��Y(D��W�\F*��oxBVY��sT�×n�s/�w=�L��n̙�"��&2�nX��#L�*Q綯���z�����Fݑ<�Y���i^��!�ˆ<�ZBy�Rx�;����S���VJ�^`~}���1^���"ڸjL��Y7ٴ���{8�u�!o�v��\�r�{�s�u��� T �|����1 ���b�*�������&�"���*� ���2K$�� ����������j��

�*�̪�(����*&���3*�L��&�0�2���*
e��������3*�)�̪"�k0ȉ�H�����$����
� �(�b��j*�	�',)��*�,j�����f����!�����������)�h*���&�3&H**�� �������b���"(��"���*��((��*�(�(���J*�i�,̙��Ji�a�j*���*�*�")��"bj�d"�b"����"���%�*�"�"b&����X���(�����J�C8wX�v��/�lw:�D�-i�K�9�I��Yӗ�R��n>��*���AB�+&�w)�0���[�MD�����<y���|a��;�o�c'��B�|%���۵&�TW���A�p��t��~���jf��d����%m���9K�A���%�w�ؽ�pҳ՜ʸ��b�߻�_�T�s��9�]B�y��}T��{H�x_�.���莮�*��y�dV�-��d��6�F�	y���c[�ă��\�X�`<;,'�����w�y�\Ͻ	Y��pSwg�m��7G�I�8c��'������]tҳ�j��GW�ʱzTxh�E}~�]XO��e�\��q�ll�^x���ٞ�Ner����-a�-Og� ��{:��eWO_�{�7�&�g�>����U��("\����..���n��H;��u;��t����y%������}�̑�-Ų���V����k�s��S�~�&6+ͰM��ͱ�@��}ge5s���i��c�,���XٌC�=����&@�hw��x�F�8�h�i�lx֧���(��N�W�j�z`$�0��.1����{,6�n7(�8�o�3RU�*�Am&�v�"���,��������,���iOg��X��Y�W�%���k��sf�ʎt4]nwV�tIF�ӄ�>>�G����2��,�-g%��W��:?S����þ��KH��h�I۽7����s��w�q���)`��ϳ�s�+�������=��������4��������$�������n�D}x}^���ؕ�d���9�gf��r��l��3����ʹ,�g��	� }�?unj�u�|b�������ʽ��3pu?v6��_�.;+���g�8�m�n�=V���жxKc���yG��-*\���(~�f��=�r����o6S(V�s�� �!W��n|}���U�ᓬ��w�ux=;q�9���U@�7��L��5��R��̡=�{�&�O��>Ľ�;�_��>�N�P��U�t��p=6:T�u`{����o�����v*��F -�ٵ4���>�iE��ާ��ԫ���! ,-e�nљ��*��9��g�͸�dYnH�7�騄1f�sֳI�b7��~U�����[{�6e䌳ܥ���=�X�~�c)�&�����^ pҡ�p�O��˷��N�/��y0��t��6$Ǧu�^e��[�S��S�ˠ;�ƭ>�Y���O(�Ǟ�c�<�X�Ho&6�ɵQ��c��O~�xdX�y���o<���~�3ю�:ꗘ�B�-�t5�	�0r�f�_U�g?kM���S򙇭͟�7���Q]��8Y?m'� ����\�r�5s�}#�����~���[��Zgl/�\2u�����}�����3��ϫ�S^s�����'����k{��I�״|Q��ڪ�e�eJ�Y�0}�'�ͼ�89��g�q�rӟ�ז�.�WZ��c�u�Kz�ڜkO`�u���u7�8y�<{7,�=G�'?ug����o!���޴:P��`)�m�[�W�r�t��>ʥX�f�#�-k��2��E}|���b���ry�t=�'ں偭l��w���Ի1<l����0̕��qr���7/#���y�b۩d��o��g�DUիr<�-��%��'�I����Ks�Wo�-ܫ}�=%��(�Q���ϒ7��e��0���ӫNv�yN��]��1��3d�z�3���ܫny
��.7��~�g��,�d�5�(�ȵ�����{S󆧶I|2\ە�Xk��E��S�WOy^����Q�;z�ֵ��;��~Q�N�d�eTfќ#ِz���ۇ�y_<��dy��4��^d�y"��p[�鿺Iu/�E
�ՠt&7{��	��[7�J�9��Җ�y[����z����/3��9��|�)��WbӋ�=�Y{��~�:����=����禲uֿIb?u��,�b-$��5�&�`u�1��[�&�f�jέ���Æ�{�wrow��k^�������G;|{o�3� ٽU���~4= b̰�=&�
�o��2�:�O9{J{&v�K��~���U���g��1�a5�U�fml�|=���wF��������ܜ�Moz��p��<].=R}�������=pz=�d/R�}Z�#�5dM���44D9e��T�K.��6{�iU4!}S����g�s;��Gxw���bZ�C)<��qpj��v�ҚݨA)��ɭ���&�.5��t�E�����SL�j���-P�+�gZ��:3�J���N��˾������TB�5�sf�����L�x#�)�י���Un�ȱ˓;A}�d=�ŋ���������7A�m;���+��~�{ks�G�of�#�:e.f5���XC���:����Q�"�Tr�zz�bV�e�����]�s��v�bm�V��e�����e=��$�xz�v�Z�6�<��=����'>�/�vx\�0;��(_C��}����I�֮׽�#>���g�ֱO&~��,Ԓ�`�6�R÷1�\�s����_V��&W?n�7�ͬ�
���K��=S9����()����vk��n���l��w�\>�N�j���rǔ�%Wl��w
�n'�E{(O%ܾ��Ж�\'���\��,�������;�=���8dqf��_p��>5�Ϸz���}X����3٤Lt;e�jy��f����C�,>�fjT�F5sEս�:�-���d}�p﹣V� ��odՏk��o2!�һJ�g���٠�Pʷr�4ap��8-�d�6��g� ��v�J����3���h�F�g���v��r��z�%����4�Ϸ5>�r_!ګ���^�^gHl9�N���9_�~^��m�=��2�W����5���z���C���et��t��y���۳:�����C���Dޜ�
�z�LY=��=E{�쩝���7&������W:�W�|�WJ���:��ո<6���kc����59���UV�쇛����~��%���ڥ�~u�ප����p��l��3qЎ���z��ͩ;:�#�g�d�|��s����e���z�\�q|w��{�^8��]~�=���93��6�ޜ_�(}-Ms����/�a.}Z<�Cgf`U���������6E�6ү@�����̝��m�BHX�o�S��j��8;���7������y9�yI{'��L�<�����ۓgl���{��i������}�.f��~����$�[w�ͩ(B�s~W��l�7������Xn�o��ʀ�Z��YJ�щB�� Yu~g�Ŗ�*FB;�-t��s1hO���J�Ki�y]��2e �85-óe��_>I�z������j���.��t�k��.�?$PWT]��άe�-�v�έpz���>��z�U��C=���SÓ�k��i��]�*[Ӵx^=��'k}�x@��,Fi�x��'���췴�+�Y��~wWɸ�IN�7�TE��	2�6��xvXOs�+�����O�+6����uv����0z��t�\N��,��;��g�dg�	�RN�f����nP�9���O�s�D���u��/$��{�A��b���q���������eL�/��1��=c�<T��̕��BqL4�7N�{��"��Y���l�Oj�����:��{�NuS=���e��z]MB�����޻k�^�-���=�V1��Ş5l*��y�-8���U}۾^�`���;Ȥ�o�ɻ]���d�Xϴ'�'g]�!gvM��y��L�wo·S���駽�$�]����2x�i|<�r(�+sl�U|(�ݣ�����'���r��߲��aH��X)�� ��I;�y�7�p\D��7���oi��/li�23Z.�p�|���}�̖.�$����cKP������u��˘É-���^f0�,Fa[!��g�xz������y��`sz|&�����a�P漼�)b�5;*1N�Z 3u`�/��.���m��������ڔ�F�Vy�ێ����p�S����B���_�s�O�N��o|�}oysn��F&._;���}��=n��c_���x�O�a�|]��vo㗓��⬷�<�щ��d�I������r]�V:��;"�i���=�]��zE�^�&u��x��wa��s����Ϛ��$����+f��6E��S�^�U��g��u��^�7՝Ç�jze�1���*�;Cs�UF�#4fG�����{ػ^��ϓ���ue��{���%�uA�����\��_����]Ix��nr=���(���v�K|iy�}W�ީP(72�N�y�T�����6����&�D�=��;v�Ү�S��0���z��W�(���(�}���ӞV�����vr�[j�.3yg� @T�hm-r�<h&wr(�O��~������j�����U~�1�Kn�]+�o�f�s���B������hv>��}	�1��F|cۑw�}�W-�;�hu�k<���v{���c��^M<�C����̳��Z��v�{�Y�=��%��!y��y�r��6oUc<�a�SM+>�~��{1z�J��3���u;�{&͓��Mܧ��纵��;5qKi�=��Q���a��5�͌X�l���K����M��rv�4�S'W��l�Æ������^���A�ߒ�uP�sgF7MΘ�໩W�w*���}㞾ꀓX��;^S#,������T�/����y�VE�T��s)�w��yu �`�9��:��;5����C�_WZ��[^���;��5�@qs�}_\�V�v^9�	ڝמ�ʭ�[}�*{֫��n/�+��]0�ðn����R\��%��ʝ\�Wo��=r�� ����t4{�D� �S;�Gz_��O�&o'�ڛrKУ�t=D٫�g��ݛJ�r�K���%9u���ʒ�4�b��ٳ��<\-jJ���;�'�-���@`r�/���^�富�[���=��L��t6�x�ۍh�"P�/�Hĺ�_���2��兙��^�	u�O!ښSަ�c��vw,����?_=}��|}^~S�s*d�h��������^�M{uFe�$�u�3W���S���P������;dHdF��m��z`�sh���I�3�d�ò�}��r��������;��:x�{-�w�ut9��=8:��u�M��Ͱ_g���
�
e������C�|Oe.�3�{�x�qK���u{�=��5G1de���P���d�Q�V�=�����Ho&M����X��;�B�+���֕��/}W���r�^򧫩�����iuxI�6G�,�fL#ö�ܿo��Tm�ET�c��z�c�Vѝ��S��u�MOh��Z�$�e���}��S'nS�[~u�����Ke�L!Z���(��������OYd�⣆��^w��rl�S��e�>N�O?}R��B��I~]�-ޱ�V���A>Uڟ��X�m#N�u��n���ⱄn��u�f��~5��	���[f��Rf������l��t,������=]��qS�)M���mj}�S��%!F��X;ě�q�����6kS����ג�-��ݧ/e@[���130����qTw��l��ĽAKG14�pywi��/KW�SxM��wTDf�0;*�N�$��E�c��
ivj�ޚ�c���{Gq�k"92n���܍�N�?A�n�s;eĮ��M�*B^�*a)���~#e�W�; ��8�lc���촖���p���PX���ؠ���<��z��Q�#l뷼u܇Ԉ}�r��0��� ���d����2�ՍX�}���v'pWp�:0iǵ��suw�G��<ImU(��t,a��-+}�`�^NglɜSX���Ҹ<ܾ{�]��׶���^j���vU҈iR:/��!�kŵγ=��_
 �>fV$��e�N�-�u�����u���6P�gZ���2�	��2��=Uف�1(��Kς>o���L<W0�%eX��淣Ξˇ��5������=�ڎ�y��0����S���v��o]�`�+��+�a�p7��8�
��1�2:o���K���3��if�d�x�.n&�w'�.r���������94�N��RN��r�v��h���f7a�^����&�Ga�t�"�pki�M��:�Hycִ׼�Էݰ�o��T��s(�؉mw�u����e�� ��c�*
�*F�ZS��Lr�7�q�!���΄����ڊ�wƽ��9Жp	��N��\�]D���=?u@�(d�����]��tX��]��n�6b�+<����*�e+Yto�q��U鸯h��]�iAԖ���o�bL{��$Gūڷ��'c��3��XXm�l�ny��c���v��7n��v-zj\`���¼ಕEFu�ZsyuX��Ƿ��Bx��i �����n�P��V��w\��e�U���Y0� ܦVgL���@�������tu�2e��6v�cMm�r?DC�'N��w��I�P�5.s�~�N�.{:�A�Hȍ�wե�K�J�ugQ�0�����fٵËoS˂�Ա`��4����`�J,	�K%�{z�	��y���9�L{eXc���;��B��=�xV�����_X��&��=l^Kk"5�K�.�`ڳ�s�s:����l���ӓ�(l��ܞb��8U��5C��ZvC�jƪ#ה2����\������\��NN������ �N�^r43&�-��d3�ޗ=Am\<�ּ]���%�(��YV[�a�݊�YQ.�	*����;ܗ��t�,�f�h�iHm��}�~�LI^��{�z��6q�W�����`W[v67Ig2����߯���z��y��(P�P�
�C�QMD�Q-5M1UQ%3QT3�%R��UE0�5E$DDITA53LAHUQEEM1ST���E34%�RR�RU�HU%PčP�5TU%MCM%)DQS2�RTM�ALZ�	�����(���"��i32*\��*�������r���)j"*h�"3������ �"
R��`�b�"������,��������
��((*��**j�b
��!��
�Js2�Zfi*��&���("
���	�fi*���(�%�J�,�',�d��|kοy�}kZ�^y�C��]_�^B�:�϶>�jy!�x���Uko��`��9�������t�w]�uB�`�!}0��"�'I��>��g���j�s�l�s��Rˋ�j�"��P_����ڋ�+�Y'��X�����^�����sz��y��uʹ0��{[��K��
%er���v��~KEIW�-l��n���9��K������yu��Yۤ���zwb{�>�{e�kKo�Y�g)]��}��v;ՙ�y�`���W��[�c�V��k�ȸ�O�V)�|2|}�?zk�2�s�v���|��[�9[ށx9=�#4�ȷ9Nں}@e���6eО�y�b�v���5ro�.�;��-��Xpz�˙�X�&�̪��ѷ�+�/{o'{P��^�{��O��aV��OA��.�ÓA+�n�	��잦/˟5ez�E���%�T�����p��ǧg�?~���_5&v���Y��Y��I�_�G8���έ�et�%=�_P��K�̕Yre��sч��	��d�=eұ���;;���B�À�&3�md|k�h�F����2V���
�c���vi������R��L��\n���,g�D,�I��r��jS�����_�x��ku�g֩�ڼ���I���8��}��_��w��ܓ����S6����֞ޔ6�ݨu/��R��U���'��\���VAp��ҳ{�������\�[-:�jS�}Ԣ�a���v�ޏ�z�V��=�%�2d���둳�r[�^�i<z=.�d��v�	�ʦ4q�!�x`ΐ�t���99��i�k���O��X���|�m�v�rg.������,����}1��M��s�M3ݓ��]��U���ޯK����_�tQw�O�}=�ͼޭw7�eVg%�^���c�+\����N5��3�hN͙���5����_9n�t��2��_�T�U�m�/�ܞ=~vE_Cľ�:U�w���Q�jS���=�ނūp��}7������U�s�d\m>�X�͗�:�k��[�g���~����&fw���J��\�Vͣ�l��#�5��S�W�?E�N�V�K������V�m�]�P&��	�����2�%8��\�p��75�S��%K�ۚ�P[f����e� 
�:���|u��2r/��(��� `��9�L�ط�q� ��GB|��3�T���..�fbkg꯫�S��{�%g��Y~�gnb��Ӭ5P_1�-����+|��|�Gsbʝ��F�ڏ�꿩��~u|s�/u��z�q+7�rwj���Ϋ}s.i�sG#�`)���S˨�2�O�	Nb�A��t��'�&�M��9 ��nm_O/L���ˋ����u�ԘJ@k;1L�隱��· �p��9�2cӁ�n���}���'oC��/Q��49������T��_W����sy��hY�SBo��e�I�٨�/�)x���?A]��A�:���ܯ��i�<����7/%������~���ξ��!��~�Y�>���_|��~x�e{�����}�u��k����߭��^�#�;���AԼ���� �K����G�7'G�h�w+�����K�؏�?h众w�}9旒��y���d?��y�.�����u���5����ps�Z��Of��G�2:;��/_�9/ �=<��˸����NI�a�����}����>���w��~��������o3޿y���:�䇰�k�4��gzO�R�'�sX����۬ԯ�9���)���7'$:�O�ܻ����7.����r�W�s|��_��כ�]{޵�}}�>��׿�����#ß�����|��]�~�s�y�y	�z�n2]�Iۘ&���۬ԯ�n;�9J�v�p�9!���份�������_�f���{���ۈ�qb^|30�a{'��"�B�OwPVl��n�隝Ǫ�hG��5m!n���0�������1�>�����r�	���z����ݵd��."�k\^5�:�[]�8��ݬ��A%0�'wj�=�>��U�$r^���}�D�����#Խ�oG!�܏����>�q�s��~����r��4nK���	�>���ъ�&磼��_��3��e~�~����y���	 ��/אx��}!�:{ޏ��:��}���=Ǜ��ǒ�<��C���?w��
��2_������~�1˒g��כK�ʟ����3����`{d�㣼M��qN�����>�!�A�9��p?@x�I��_��=��~���|�w|��K�(����wXXί߿`[&6���m����x� �>��vh�~������u�'�r�S�q�!��'��i�{����9���_ ���4�qoU������!οg�=n�~ ���HO���d/G�5�uӒ����/�WoX��?G^`{d��w!��OOq܇�j9'g�hB�v�Z:��4�3��%��]�ݣo��	���H/�)��z�~��oΎ�y'�ם.�!zs\�R��C!�K����rGO����N�0=�.Ju�nSج�����n*�o�����o���V��c쎣���ܼ����4����sBP�/O9�Gr���z���</���y�w���>^ǏX�9�:@����K��U�Aۛ���q�����+��h������>�G%��{��w��<>愡�/O?y�܏R��=�u{+����>\~�B d}��쪩������߯+������!�q��'�!��C��]�]�`�A�:~��)\��>ѹy�9��w��9�C�}����u�}��c�:~Y��{@8/+?~��w��涴=^�Ry!����X&�tu��Լ���}�����/pnM���ܯ��ߴr^F@��|��������~���Ǯ�y�{�]��'Öo�Cl���x�����:6,�׉!=%���1�<{��{�6��������T*�9	�u���@6V{6>��9��z��/c����|;�����J��O.��WȔ�0�����9�XcW(5L�ĵ�M�4(��������>��}�
u�z�N�w���~�wm��ԏQߜ��>ې��{��cS�u��w�y�K�){��9/ �`~�p}�wJ�;7��K��yy�_*�~��V�ܽl�����������6_a����t/����֠O���~������9=�n
WG_��pR���NG��?C�<�߼�F+߿n���r��<F��~������<w������Ӟiy�?�:ߝ�{߽��x��~�����R���j�J����d��{��Ϻ�y������_~������#�O%�O���л��oO!�쏜�i����;旒��y�=�BvoZ�K�=��R�@���FR~��@�w��q��ۻY�<�]{s�7���q:�%{�%�!�0w%��n]ɾ���P��������}��~9��%=����<�u!;����pRo΍��3v�{�9���߾|}�\C�7/��a����b}J��X���J������)�w'G{���]Kپ�r��=���Mǒ��t���n�s^�˼�k���f�{����A@�ϴ������n��p��GR}���������07/��~��`���o���.���z?A��w��<�?g��s[��}��߇�߹����n^y�z
W�}����}��;�%�2^�`��}�����t��������O��{)�a��x���|!� ;�r�����v�x9祣��>�۴\>������{��;���K�}w�R��|�K��~�G$ԿFK٬p�/�a���=<��;���>�/e7�����9o���\��o˳�����������}���>�ox���)�x���^k�t�!�޻�u��k�j_�`2^O����~C��~���n
o��~�����ܾ�kf;j����9K4&6�|�f�_N���f��xz�����C�.ص�\�r>��w�����藁e����oSԜX#z�4��br�X���wl�<W�[���:��n62��y7��&����s��� �}��)�-����|��|?C��:<�B{&�Ru�����y���<���1(7/�S�`�>C�sΞ�y���K��]������I���Q�̩���{oC�M~����>��u������awo�����S���FI��������<��P���IA�FI��4%���y�܏S��~��^���I�4���U��gW߾�_��^�.C��bnC�|���rGGx{�ܝ�bOR��3�>��t{��AJ�t������N�~ʥW��п�����.�y*��ݯ��������^��~iuy#�q���>ߤ(9!�=�G�X&�<�����^C�|��K�/p^�䞛�C� ���@;����Y{��g�~+I�<~FJs�I����󘇲�������z��y��u�~�z\���a��	�ƣ���nG��=���~_}��� �K?n`VA��ٗsw��~��{;�=��<�G���<>�K��O9�%俯a�x������B���=�~���;<ޗ �?Hv�r��"Ư� >������_�h�7�<?lz�o�nw���]�쿣'��?C�3�7=H�OO���y{#��kp���=s����[��}��|���u'��L}�K�o��U�n@h���{\���3yǹ ����P�:��}/#$;<��NK�����A����Wr~�Z7//d|9��C���K�#�>6����/��gٗ_����d)�7��|��M�Կ��a�_�n{z����Ox�������份��qM˸:7�~�y'�oG!����~�>��u�u�lu�zN�g��a�_�kw\��&��{��Oe9��nu���p}/���?C��:�����n_�$=<�ܿK��<�C���/������#�����ĪO�\+��/��|�s��]}�`���	�5����E��R��V8y���!����V�ޱ����1�&�s���~�ʲn��C<?;��k2�6i��t)�w#�q��>@s<�LY��?ө{� bn�F)�^��<���W�m<���N�Ͼ��{�砓��Gв>��f������i)_������
�|Ӹ5�P���|�%~�q�xOR;����~���spG�|@��q���Ac��f�tc���������rP��������u��=K�����������]���d�FK���|�%~���x�f+��O�s�����:��<��~��#⟤<����ZCr�۽��?@y���#�~�����yr�λ�(_���=�u��k��_�%����x�U����,��Vߦh��~}�QI�b��������!�}�A��By'����?Hx�Op�>�@�����΂��=�ם�/�Ɯ��������t�/��D���d}G，����_e��;��_�ט���~`r�@����=�S�;7���ݻ�K�(O��A�>�O��A�����~ ��#�u�����.��¯��;��rG�}�\����X;���Q��)�#���aw~b{�������;�O$䎣��w}��#�^����C\�6噜��~���2?�Ҕ������ܯ!�z�ט�<�K��y٬M�}���X��<���;��{��=��������pO�����m�w��v�~U��(\�?�h�^ABvo�|�r����`���������R�sޗ^⼼޴9����C��y�	�O'�4�?}��!9���|ոկ��/�'�}���_ �'G�Ѹ)g�ߴ�NJw�4���&��y/��?s޾�Խ����P�GsC��~��3����8��r��R��;W��)�o��3�:���GR�/g��>��Wo�/�rN����ܯ��{��C��N�9�r�_����4����<����S����n��n����LO�U���h�:E�v���e�%��:���O����=K
�̀�U�x�qN��o�����K���5<# ����.J:�����o*Xpv-�P/��
9X"Bf��v8k��H�*��7�SSV���N�����>�|��x�o�"��D#O�� 0��e����9#����R�������#�����Ѹ�W���y/=�vs��K�w~����C�}���7����߻���g���f��=Hq����{-�Ծ��c������P�z��伂��O�ܻ��$I�7��l����x:��~���e�9���u[�����;��uW�n^���^�b��������7�:Mƥܟ��5�~���9d��9�bn
G��p�rC��O�ܻ���1M˹>�]�k^��}�o�������y��o��{nW����9�H�s����}/��K��n|��!;w�&�%����n��9d��n=�9J�w�M�����1��_�cP���x;�x�������r�����h��#Խ�z9��|?sT��n7/�����iu&�=�h���);3�K�a+����o������5u�����nkg���;���k�~��0?K�wy���=�G��K����=����ǒ�s���w?u�����n��)5߷9�u���^~����9�_g ��|�h�I��w����G]�~��❙��~����u�7!�;�4}n�w��9K��G��H�=�پy�R��^w�����y�g���Ne߿��{��=�\�!�9n�����f�Gr����咻����^�u�;��>ߤ���!�`��<����iy������{�����4gy����޻��u����R���;��2߼�!�?NK��_���������l��N��9{)��0��(���� ~#���Z��+{U<���uύ�W��'�����_�S�`<��s���W�oz��d/G�k��]��y�K������w!�ty������a˒�繛�}~�N�#���������+���^"U�r3�8�qN"pݖ�!s�]tE�Nk뻥�Ŵk'=Ԧ��3M����V1�i���)Vut]��`�	�a�LD�wwX:j�2nt}�U�b!�V��*-��FGm������o�}�� ���J��z����ǿ����?��MA�ԟ���~��'��ܼ���7�%��=�sBP�/A�y�ܯ$�z���<�����!ްw/��{=`;��k:�>��x~��Z*~����l� }�}��yK�8�����<�AJ�x}��K�)��A�;���}�	C�^��Ύ�z���{���W�f�!�� Uk�������~�_��,����־O�<�����!���:��W~`�A�:������ϴn^F@��i���ro�_e�~�}�=��:�����ﺵ��w_lu~��=����
M�y��u	�=a��/$�>}����߸/�n���Gr�ϟ~��y�1�K�=��5��~>�5��e�ð{�|��R�e�_K��O{��u#�voK��nC�ǹO �5=�`r��w�AԻ���1}���
������Zw��>�����o}��y��}��￷]W��w#�ߴr]˿�>��H~��?�o���}�C�����-'��_�ޱܯ�����������
_!������~����g}���������`��gx{H��y�����F��?����iy�?���B�!���A���{�~�����R���`� ��UΜ�[�~��3_����������?]p<�������NGr��rs����^I���w{#�?ZCp�}.���`�o�{�<��`nr��~ p�,�����IfJ�c���uy�é_ �:��:���XK���0~����=�7.��~h��G�{y�<��r?�bC��_�}��O`?z�����<`��w��,���u�A�AI�1��_c�XjG�?F��5+��r_��(7/�y�qM˹:;޿_B�^�ގC�����|?G��?�}���W7/���`����<�d88����꧰�f���AE)�yg.:�_���朤t`������	�er�6��XU>a���pפYq^�2
'�<� ��7�9��Q�;��Ӯk���i�6�
dZ�ks����}ػ��W�U}_Vm�����z�׿�jWs�;���PP=�O �w%�~���F�;����:�����ܧ�`n_�����hD ���3��?}���>:�ž��O�~�Qp����z�GR��4��8���C�(�������{5�n��{ш�^G]�}d.磼O��t��$C���?>����_���6�Ol˂}!����7#���C��_�wx�@����]�� ��=�u#��h䚗��{u�n���;:�a��"Ǘ��G�� g���N��g?~��ݒ������~v��_������
�94��5h싳T�Ot���l�by�>��������q�����`j���z,8=Re�k����+	<�v-~�z�G����S�]���OB|3T7d�]�}P���lݖ���7݇��:׫��� �w,;=�S���fT��4=҂����G���l����+�}�Poo�Z�2�x���u'��Q�㚷�~O:��.[�ڌR5�x�7ɖ���Y槯j��6����t��fδ��Jܾ՝��x����Gy�Jgާ=�޺�8�^�$��=���m��U^3�+���"�I{�����bK��ƣ-����9��������Ս�\�Y�4M
	|��N(\ �:���qƏV\�N�x3�ރ����Z���cJ��:��]�&w�RWK.�P�5��JQ�;�"a9`1J�ml����jR�u_Ì�d�&t�nm��"����F�+'�A�h��p`�Ӌ ���U��Xb�y�~bS�eG�F��	f"z��O���Vr��q��雞�4ţ���ZhҤ�f�뽧��+�
ɃqѫaN�D���a=�cN��t�zm�<�T�:�.�����,JN���:��Hc/Q���vﳠ<��hzp�����G�#}��QN+���z��n����_�8do��F�*��|+��v��-��@U\���C�l��^y���Q�e��,�"�3;��$k��Z���!�q�	YtW7��P���D����l�g^��C})��X�b�9[�N�X;�R�.Մ���^�ś�F�
L�X����/��oC�(����ꯢ����H1jSr�Sي�μR�V�sĸQ#�[FAW���ә���Nb�o��W���v+��*Գ۽��l;�{RX��z�.�xz��t��2����E�+'n!Nvw��6o�@����Q�������ٮ�u7Y�/L�j#K�L-4��wr�� ������O��gޕt�5F��7��e������V�d{u��RԦ�5y��됣�&��C!�L�w�w4;3�pW�;WKV��5�P�PN�+3��>V^�P�qދ;���q�(�Ѿ�V[�[��WVoF�bQ3m���Ɲ�O0M �ΫyW��,ŝò�7s�Q���5�Y/��҃R[�e���w����	(�~41��ay���b9�|s_V��P���AP�E��wm<IB&VU�nwxܹ�ޣG���Po!�l֥Ul��$B��. o��p�XB
���u�'+��Z���ܗЂ�e�S������3XǗ�5����U<�ް�����ԗ]�%8��U@}���i��D�;ʳwk0b�ߞ���9Y�����`���Ex�i��?=��Y%=�]	̀�{sg%��u|ĕr����4
�[z�AG�՜�������	����V�1�!�\:�C�Θ���@��b�|��d���/���!��ٯ
��>:t�����w�1 ;��NЍB3a��6�놻�ضY��'��=�R��V�]\�5�0wNl,��e��u�z�#?=W|u�/
�����nk���[ԛ�psz��.��� ��P.�)�Z�n���+Ŵf�Ss��k ^ĮOd��]gϫ�eM��QhK�'��3�;�z�?��Nv�Lb5�5�Z���L��.2�Q@�a8�)��kcy�*j���NE�Z?H�MR#�nu���x���_?7����@"�
(���&����J"���#	��+# �j�22R ���b��H��s1(�)���)h)��������	�)k ��r(rrj����H����)2d�����2�����L�B��"�����))���B�\��
�2
��)��,�h&�
c3"������&�B�H�
�0L�J���j�,�J����(l�%��H�(h(0��L *��ri�ʳ1(r2��� ���r2L�ʃ0�22�3,�	� �(����'"��@�\��+	Jk*(20����h�2G*s10 )
bJZ
���0s0hs1��*��20$�*�JZZJ)i�/��>���*��3�+s�<���x|,*�K���'z�Ks|�E�qTƀ��5�u�;f��a]gܷ5噟`	M�)��Ti�2�����@u;y�O`�Nړ����d�}�C��{�w&9��l�Y�0^�+c63�7�t���ܟ��;�������7G��vʔ����XoW�ux�9�A�o�gG�n�ɳs����6��v��Yw%0I�9���a�R�m1`������]i���7�7�r�[����ϒ���2�������䃛��uOZ�\,����:������ᝎ�-{�1];_Ac������n���}w'�X�*�%�x!�l�+}�ϣ�Kof���:��o�ſ\���<�����l�����s�Wd\E��v�O&���>[���Vs�.l����&~��pٹ$�.m�+�|=��cw����k�z����6�R{�hc�pj��c�;֫�x����X�q<�����6Ȯ��G}.{/�?9��x�W�3�w䇫uV�[�\(7uK��`�nr�+���/6-��b�8��i��:iÇ��rI�Rr�u�'kmw�B�e�� dy�v@e��熟j�{
6�p4�>Wk����1��_R���%���.����4�FEx�]�'V^������  t��ɓ��'0{�i��z?J���6:=����:�o˭���n�up����r�+4��C��~:A�76�t����Ͱ��wѬSKޅ�u>�Ls{�V�؟R�S�{T|y�x��Įi�ڞ��Z�<��w'��{"�����^b�b�%k������s��=�_z����h���w�Ni[�����aؿz���r����W9ɹ���^�UD�L��^{2^oA����c5J�;�������gu��qN��#��ߢ�N���A�:��o��ݽ�.N��������W��X�:�>ϯ�jS�W����_�����y�~�sL���^T���/���;+�--�uw0��W�jN=lߪD�^�W�s��6��LF�i����4�����ۺ�{PK��{�������z;{�C��x�>��ͤ ��9�DP[7���44�/�j[����yQ{��
DM�̶��2���w����*���=z�-���er����Z�]��T߿B�qym{�,���0��b��@��P����Y�ye�k��tΣ��d۰@���U�8�O�u�����f��}���y]�]��>�{ևu�+�{=e�nu9rs��gg���,��O�+Y̧����;���x�}�=��зk+�V��L���}��]A�1۶��A���᪵��U������v/��u3ᝉ��2�-q�G"�c�KkJy>�+GI�
e�m�v5;j��՗��"��n��d~[��φ�R�����n��Iu�ph���=l�S�^����;I(�~�C�=}�-���]W�'�/�1���mM˫<�;��<�mLu�"]����({Uj���s�h�)�c�Ę�����^]��T�������uO��/U��3ݩ�Rwݴ�����!v�.�.�����W�'�ߡk~���/8�
�/Tt/����<�V+�\gO�ڣ�e�u'��~�<�I���E5K�l�V��}��E���t��je��7�y^�])�Gw.�Q+��L%�(�����q�ڽ���6�=�ǯ��U�%���d+����7�>;]��Շ�`yg#'Dq�s�A.b��<��!�v1N��"�kz�I�P�'L�4E�aY�w
}����<8�6�|>|��ܽ��{]e��������8�~�k��w�PL����Q�s,�i	��o:Cc���	���96eOKi��o]�j;���!׫So�v��vD�����Ɔt~�|ɵG9�������dҠ��nd�u��`>k~��zp����`}/b���o[	>SkF��}J��7S��Я���c�o�[ʞ��]���]��(H����k�S��j�m�x�Ğoq��o��]w�l�֍iȈT�d{�yN��b��[����I{yq�T'��G��=���{8'��T�&��d_�����=^�y��O݁���
�nM2��j��?xE;Mw��嫭ˢ�K����)��u�gk�~K�N��Aa��83�	2�����;�U޷S'e��7>:=����r���&�BP�aP�p=+#���JcٛP�c�]gV
ߞ>�=�C�ǵ����N��q���Y�u��J3���݋�pw��� �]���������:E��i��Cc�x����y���Ć���Ｑ���s����1ckv�͔0>4���o��3���5�������;ݥ�u��\˩�ro܎�;=����sw�xQ;g����|%�Wp���o	�2�jr7�I�_�F��j�q�<����B��Vc���y���Xש�K~]�Y��O��^�3~^O3ju�XPY��H�]fx��<�}��7�)R��J0�1\���C�M���s�cg���ۗ���\�%tcٷɥ�gف}S`�����:�v�ɜ$�����S��f�f��w_��ӽ���j~��c;z�����$J�R%��ȡ���*shzq��\���~�QYL$�]^ͣnz���݋��j�:[b���񱎚^j�T2OX�	�q�ߖqǗ�vשy+|�`y�	Ʀ��t����ڶ������v�������i�NS��QzW��ڿ4p���,��Cyd���҉e��d�2���x�A.�R��`D༞��쭜���(z������NyGθE���o�yh妃'�����c�K�r���rg��2.�E\P+|�ܭ��r��{��MhO�N/h伤�e.��-nE�%�v����%m����$�#��8e'>�����Q�uݙ+|�=z_j�C|^�J�J�Ձ��]\�ݡ��N)�X�Zҗ^��	��L�h����ꯇ��K=#��L��4�W�g��ԙ��Wk�P��*b�~9�]Qh�NVVb=�׫�gs�X��xط��u�P&Z�|Y����P�x5�yC-p8&T!k��]����U�k'���`�W�V������5ژxK40��שF�<ʨ��=��������v�R�Z�L÷N�s�X���r5�H�^���o�f�8=��_�t�I�L�93��E��m��F.�ʌj���)�Yс��<%W$a�O�������ćܸ^�k4t�v�T�q�kz�����CR��±�Ȱ����㳽�g�T�ǆ���*k=.��N�w��p����3!��J�W������y�Y���
�����]��̹<�WD,�5?v�;<��Z��^!�-�}�φ׌���Ω
9�j�OV��{�"��asۆ��n=U��Yb}~�0l�*��U�m8��g;��ޝbj
_�����^יr7D��S��g���4ϖ����f1�s`c�|�@ަZ���L�rsZ�5���Ǯ�7�أ���u���a�X�	�3Gx�ej2#O��5�;�Vv�.U���N�i��6�`�L��_
�T��覬����m�jH�sQ�l�\$+m~����e�� ��'Wl�Wp�OEMe�[H.��.
����u���i���'���  ���];�s�5��c���]�.���C��C�*��e*E�LP��H��K�\�>7��n�[：��ON�p��^�}��;ֽ�*Z��ymU3+Ѓ��!BV6�ɲ�a�i_y��>M�~}�C��{qdlw	��kwE�̮jC��Ys6�y���p�gʎ�x��Hu�Z�ȅз��X���a�8�\�YeW`^����k���o��\	i�o�)�yM)c+���o�홒���Ξ�?]�USd]�{���#Xo���pv�@��k��O��)����7�Υ�b�7z��qt8��V�a���P=ǌC~G�éݓ�1(vK�+)N[yv/iL�JZ�����f�&�{�z�LAn.�	z�sg�:�va�u�hّ傔=�Yi�����{Q�΋�����W'W�Cj���+�@p9E�Q>:˨q׮���H�Yr^��k����i������Ꭴ�^�k2/�"J��:7�v .+k�oJ<�w�,��s:�Ź�Q\킲����$%��h�\x��qw:��R�ռlu ��x�~�u��:J�䡧�e�[��g\�̋K��F��\e$��F�]�5ڔL�&_-yV� ��܆�I(O[�Z�{��F��:6>W&��7��������s=LB�^Y�U#�E��=A����>�M��Y+~���$ItՉ[���_Gy�ݝa=Q�kgdXX�:��t|�h��_
�}�>�LuJ�c��b�+שbm����޼3Ϡ>7��ln�}%i�������������a�W�l��ElMf
f��?Q�שn�׼<�W��Fԯyh���}���Rw\�u+ �٬�c��fzl�y��p:w�T���
�π�w5{��{��ۂ�g�Uw>;q�x�Ń%���g'�P��ϥ�|�'ظ�V'3����)8�:Бx�r�4��A0k�k֋3�{��W
���J골�^��eઍ#~t�y2�?N���C6
����x���:�gq}L�Ѯ
�CM�R�|���t�Qv(�Fg��c�/��U�s�������io�ϼ2:eN�Q��(qB6����/�3���G�	�h�:���`�Ykg�M���?A�&Qɛ2�lᘉ���D�G�c�X=K���M�t�>�鴦N[�ABt�R����;�[�Ki������z�
�*�S>�|2œl�+�O�yaB��t̸FF��|�Y:6y�ѫ����9C\�Rl�>��#.j�	;�}���0�=OF���+����@�Q��+�Yt.fw���:f��S�����<�s�	W��"��䩋s�1�8��$�\�Ժ��h�ت�����m�����������vW��c_��0i�^�r��W�o���	��.VudUb�W�-�D�tإ���Ŏu�*u|�$�=�]�p9D��qM��/}د���^���G�^�J�x�Zs�v�&]�]�� ��@��7��9G=�{����7� 1!�I��O��x/{�P��,��3���5tb�S��h�K}�M���W���Q���0E��Y�v����,�=[��;;�o��y��[E�]yL�caՇ���:�Z�Cڡ����K�`���ݵ�ܴ �ב�+y��	��*��>�r/WF&Ko���=W��	���Z���������X����o�x<���1Zw��ޣO{?t�t���Qlpf���*� Y�ڹ:��.j�0ȻU�Zv��t�^}��<�4� ��9m�"]+�C�a�s�y��H���S"��{���9�2�V��m�m������Z�&�I!�G;��V�0��H'��r�$����xhX��H���#K�d��v��d2�!)�m�iUW�d�x&���ٲ#�cn���8���X�yL���ht8G�sB�0��MM���5�t)����Uu���l?���������p��r�&��_�C��L�F���`��-�T6e�����W�P��ۆt[��g��{7��/��~Χ��3�-�!��S]F��e`M�`�I��	�T��N�-����=W�;������/�[,؞�pL���H+�~,�l	���Y\�0� �-�']ҋ������r�!߾���ػo�';��g\"�K�زM7�5�lc��U�n<�$�t�9�E��;��+J Cg��{6�u�;�>��&WOP��2�,�,q���(�۾�i>�j���]KJgo>����/������R���fC�C-p,ţLt��꽰���p}�VRtG+�W��6Em,)���{}Y��uh�^�3�B��{�ϷN�%�ub���'�j%�}K�!ϝb6&Ay?`���޿^���S�u���yv/�O���F�N�(n��۹�Q�����?�Y;�0��,B`�K�X&{�^��>u}�ם2��~�=�'�����r{�3��CR��Ao�d"�ά =�[=f�zWa��U�XN��ZT�8mfR��}֯jf�hqv
9�m�x\�iweg:���qmb�n����*�<kOD���ά�YR>EJ����r�:%9܁i
��9�>
o\	�ƴ�>�
�L�}�|U�W��1�m>x&��:W��a����%�K�v=��{w9^�GY���x��3�O�*��΍]�kj����V��l�ܽ٩/@�v9�.��~��6Y��l����x�)ӈ��3�J��V�k	��{���;�a�MC�����׸]�z]ǚ�e(��8q��/���T�o�ؙ�F�� �g[���H"߹�Yx�jgI^Fe� @��e*���Ðڰ�s�P���,�B\K6
jV0�ܺ��v\�4�ӡ��Sp��PS�eѴ���F�h�||�믶Me�7�BEɮ&��=�tP.�
&PN��͡u�$���;�ի&��N��u�-������wR629�neV���ͺ�d^$�m�kn����B�j@�Qs��ݩg1�[��e2�Aes���e�n�@�Nʼv�YE�<���&I���!�m��:F�=�Ԕs�Tu���˲6�hXE%-#.�F�寸��kcw[Z�>c//C�-m�&7ׇ��>�bv��ehh�fP�x�#F�X�@�~�U�6M��4X�sl�\�X��<��XF,��f��?���UyM�����<��ܨ��5<��#E�w��Nl��
��1�2v'�9d�٩��d/z����1��ټa���2��啌GJ�xw�!�S�A�n͘x�ݰ��M��q�6W�]����H�����X��i�r�z/�+� �-��GF�&����lƠ�<,
*���k���s(S�8}Z�a��;7�UѧE�e	d^���T:1ʌt���L�x��sNwZ��pqZ�`��uFz�ѽ�F�Y���B�/�c�ӧ]4R���ex5P��	Ys�V��`�e
��m~�ߍ{����Eh,"���H�瘸���fn���K�%���U�)U[� n��և7H�9��mvOC�顸��->|`���fUgj�γ�dlb�7V"����k�&�/e�ŕy%ϼp�=N��%S�����sq��9�r�������@-�0����j��X��Pﯡ|��j<�IƃU� nٽ�*�դ�;�%��C��&9�k�ˑ�.��\��}Y�r��!ϒV��sg���=#���
Cڳ�X/x��1��*��c���5JU�����ZF��,�b��ǜW�8�X�ګ����3��Tn]M;�������gV9b��a]m޾��U�/��g�Ⱥ��>h�����y���%qCEe�(�:�ݓc���5��>�{⽳��sG�#�s].�5��Z`n�m�L�}mX喻�j,����8�U�qzl�q��@@8;<W��՞�W�8��۰w��f�>�$��G!)J§!(�i[12�r
2()�,�����)2JR�@(��%ʖ����E�*�C,!
���ɥrB����
�
G!�2!)S,�2Q�2,��2(
rC%�k"���� �C%A�$r)�hh���ZP�2L�l�S!r\��r� 2r����(JR���	ɤb,��,�*	(ZrJ2������i0�$�B�r�h������rJ��%hr�JB�B�2R'?}��tu��5ֽ�=��q;��ZU��c�)�J�/�Lnd"�egt����
t-WW8��չ�G1c�}���p�>����35�u�d	#M��֙�m�3�Ԡ/W���@���:��x@=fշ�]KtP���g�����_����xq���զDsk�_K�=�됡��L|���5����SH�O���`��œFܪ\i�f���H�3��>�Ӊf�2ù�PKm�;����n�2=�4�8^]�=�[}Z'����ӂ/uV��;t,'C��T���ho�yme_K��u����z�W�<޷��%���7����>��&�kT�B��0ҖbB�N����8|��b�z��s��sO�8�����k�\ۇ>�-DA���"!��pm�{��X���H�Np>�WD��ɴ�������`�+�#`C�Of.<Xsn��`�e����9�g�E�򣣧$;���ǖ���>�Ko.����P��<���*�f\�DL�]�8��D���j%��N��)�`e31q}G�×����-��gF:�p��X��{�	fgL�x���ٶ"��jWK�{
�/쨔63�M쯳n��� dg�p
�^y��3���G���wdקs�Զ���s�͞}�!������pǝ��.�����&5*v�82����:��^�zm��zp��RĤ6��_t�ìvf��-\��wF�	����uV_��{t�\CQ]�z��H4���� >��l����"����뇎5�`�L�
y�Æb$P�\V
[k3*0�^�뭿�1�C�������� �b�j|����]�^�����T��u�ѰdC���=�^&��a`�m|��.�A}����� �b6��B-�� ��9D��u|z��y�*�0b�_t{�x].�μ�U���.�����ޕ��IW�
۱�����j{-��<������?7ط�y���g�	3���W����?<�e��a+Ρ$Lͪw~��ɳAk�]�*7�o3���M��;g�nV�!���XA,�FR�`ݫ<0mx̓��[k���J����^�l�B��9���i��
��>_���[��������X��&[��o��������µ�eC�.�/|z(o��p�z���^s��~��x�ս�%c	��%VMy{��S�Ik�>�ĻI�^�U�p��k��fɢ�*\�#P�p���x}�^Y�$*����6�ԏ�\����A�|��u5���u���/Pzy���ƙּdZ}$�*�{���y��N3�v^�>��y/ ���I��3lSX���;�b�qekUy~�7R���'�.e#S+��֚���8���)T]��7/��d]g��g!��̛�%k�	���/U�
F�2֛̃�M�����QY���>>���>���h,l��c���i9f֦2"�z?:�}Č���u�Vx;Ӽ!�=����]����O�*��}8�ׂ�!���]��J��}u-2�gG�23 �2�Z�~����.�*u����fu���^���Ϳ\�\P�	:o(P���\TS<�޽S.y=���>b�]��O�I�(�͙K�o�S�q���Y6t�I�C=�B� ��o^�^S�
�͝FY�M,h[�gή9%6$��s�1�8�p�i}��i<ܥW-��<�'����
�}D3��ثZ�W��3eyܱ��f2*>P���L�X�̫�.��=�d�+�i|\Q���C|f ��<�Q�>R����� r���n���=�N���f}�3�×�����yh�xU���>g��|�7~t�:��Y����\���ǉ>�L�
�M�(�X�ׂ<��FJ�N�3���>7� �j�N����s�9Y�y̹�V�Vp�eh(��&�԰Gh�������t��	B��p�{�9���ag�S�����zb����j�]I�$tD��V���#q��[���4���-I��M��vw�f���7|O�nŌ�N�M�w���,R��XdkaV����Z��(������<Oe��9V��NI�˻3U���Μ��  ;��m��}n)���C9hp:wyx��`��Ǿ��;��Õ[�sV2��������ޮ��ݯ;X�l!�A���=������=�_��A�l&�̖��}�w�֔~��^�gN�b�sʭ����Z���Ύ��ƹS�d]��N9�W����.�=v������g��m�&ų��{�:�;�4���ڜ�u=c�_F�/)��U���W�dA��o�d5�X���R��탧9D�5L�9*!��n��>m]n�Om�<p);�T�T�=�K�F	�lI��H�k�R�n���"�/B���e��=Rc��޿^�v�ｔ�g�
柇K%��n+�����P�;�b��J��	�N���jZ�X+g�Ğ��ᮡ���Q���k�;�5ǵ�q�W�.������Rf˶smyO��u`����#fW���.3~\�q�2�z�j���{��QΥ���OS7����}�tZX*S:�=��K�u�+ھ�'��I��\��V0&������)����3���4N�$���8�S�9��>�}�K�9�(�*�.�a��"ZC:��?>�p��3�L������b[���V�����v͡Y���4X���V�vYH�f�EF2�[~|��<������x����I�v�����`�}=t��6Em,�2������h���KLC��[.���nS↚��\C`]��L÷��!��<ٔ�i�>o���^����kL�Z�����*'��4"�a�OWDO�J�fuK�*]�ϩ�kh���;��++][3=�/_�����h��,+�Ȱ��:a:l	޺6f!�1u
�Nr���O@���f�Z�>>�T�2����P!�`�7����'�e^pܘ ��l������Ƈ���B~URˣ�xr�kB��,�Dsk�X.��{�B���Jc��VM���J����qʴ�>�Yb}|���B�������2���vvj�K���N�Y����(����ߧ�n���uW����q�J`����Xu��}ұ�ʳ�[=u.s�XÁη��d�_T�}�zVC�Y4C�*]2��*����c̍炰3�P��E��|�P�r�ɦ��r��N��8%KQx�9jb߻�2�w�]nαgV��/n!#�2vF���&I��L�f��՜/��T��铲9Q��/^*�y�aT  7ge�޵/�A`�(J���ړ�g�q���v�*6���r���wc��Y};��f�n�H�b�n��)Wt�+�W�|\��)\׬;�~��W�ҜW�������쳅��`�+�ޔ)��/u��a^�������e��<;G��Nlt�����[�V>Ҷ��C���s7`GC�����u;�t^>���Dw���K���3�&f��e��E@�<��o��{l
���Kq�K�.�:�jɭ_M�'��F;x���ٶ"��#�n|�h���9��=xϻ��<s�����W���e��"���.y�<8z)l�ZG�M��K�Dv�Tyޞ���p�;�5c]i�L�f�yoъ�� t!۩�!ϝb�lȫl�F���s���gm�v�z�ֽ�5�z�xz��c҆�U����@u�-p��y��<�f��޹i���䃫 
0���e�n��P�I.���`7b�g�e�}�d71×���b�pq�둉Zl>�H����pj(x��W��\�P>٨�;U3�jѷc2yK�=�ŭ'�I{/t� �i��;9�+!��F, �,��Y��Y[��=��dh��1��"o��En��v�ݫ���S���Ҧ
t��*���������7y�,�%✖���N�5�)�������C���%��������fsڴb�}�/_SX�Z#°� g����
*W|�R}��zS�a���{�x���}��+�����a�j�o�.���K�i���c��\~����]��~)<]t�ͨ���������.}�w4D���uT��lL̓}t��ڭ���M�~�}���	���C�;^fw���}�6���Y����
��b_y����R�����ϫ�<0*�1ӧ��or	�]�.�<On�=X�=3�ts��z� u��g�|q�A��sW��L�YOZ�,Oo7��w�Ӝ\8<�U�Z���mjc"+G��ι��$;�]fY�ϯ�u�)[�Y'jn�{xO�oh{�~ڀ6hkϪb���|]���*��.��r�3cҙ�n_�kYsgy��y���+����NT��su;�G���!�`�KNX�C{+iq=~�g
��t��07|�N����9�(�͙x	��`
y/qQ7_M� +��N���ֺ�a��s]��"ř�y�5bu�ή9%7%L[�Ɍ�ub�
znz���{}�cs�IB|��Z.�h����3�ӳ��|�X��`ӂJ���U�����1���L-f�y�C�vΠ>��}JK�|QٸC���H��J	�_a�ڲ�JƧ�«E�����z���79M��,�����Έ%:C��|�wg!�f����QfeI��J�SŤ�@M�������~ާOk߇�����2vK�=���]%z�G����U3�����E�/��Pء�]�B�U��s���S�z��+(���X|?L��׮��p&)�g�+����x����*�C�k,���6���c}�}��P-=6:
d�(�\���0׷�!u�K˅��b
�#���[~y���[��jǋ���P��
>�,tX^��Gh���,������/ug�z�8����}[E^�}�Yu���j���������Y����0��u����&v��X�q��B�����ý��v�M^�W������8+�ժ�|M.��v��V;��{���en�}�ξ+���V"�O3�D1`.�Ε�H�z��M�qw��k�5p2�ͼ�mv��2䎈%��W�Zv��D���m��R瀿��
��xԫ��>���}$^lV'���#�4n���L��u�^���|*�R�_�H��F��ޙ���IǾ$�]��>��j^.�=`9cL%ζ\�S]z:�aFڮ���$2E+��D��Ya�=ny��t}���������fMK3N_NYy�bg�}ŧ��+��x��a�u
�;~�i��Y�s6I�k٨=���z��c�3�C�����1}v�OFa��8=kfqTk�ЋRܣ�LΌ��Χ��ar�؄v�sL����1P4��s�����읏��D,�f�_�}�7<%�A\��D������+�2�{fyy��.W*�.�秫!�Y� �������n,�.���5�7�NyF_WծX�Y&���7x��
�t�f��tE�cU΁�k��bP�X(&)SЫ�Ƴ֝Y-LkG����=�����-�+�+Fxp}Z�g�OxXx:nP/Ҩ���3�*��@�KR���sr��4y}3��k�R��+sշmm�&e�T"�`�}=t��4��3�������˲�Z@��W�p�M�(e�-��2�U�1]Ȗa�ʢ!������z�ə��$gy�b=��>�w��̼|c���PJ�2EG>�f8)�ΔN�ҰهR�'�*�ty�;.d��)����O1��ܼΌrt�yn��	��b���ugL'M�޺3e�]~���[!�W�CM�h�C5V:�x�Q���������f�'�b�s��|�z.K�ڞJ���(�G��ˑbǲ�"���B|���G��嵡^�Ŝ�Ȏ�c������ʼC]zJ8�Q�ӷ�_=\��q�|�A�V��ԏ�:[��q��L� i��OR^��@q�N/;!�.���W���O9�u�m����+�<��Oi�J�u5s��ś��T��iN��|�ӝ�l�U�׮tHC��ٓO{��p��P�;��S�ڡ�V:����'��|�!P���11�%U���I�I�v�X���>�ͯR�M�,MC�q�o��7rOxiϢ�Ui�#�BӠH`�9s���7M�ǻ��4�6����}�̺w8>�0��η��#��~�����<7)-g]�t�7z<rҙ砾
U��T��%3�:g��pc�T9�r��4�ٹ�ε�sn�LU�N����.�i��gueUC0]QuO��!�V1w+�N�!��1�W�����X��z���V:6gS�,9���Ջ��cP�Y�&e�we��C��:���?pȚ�]��}����-�O'�9�02eNH����n:ip8�3�B���7ߓ3���1��R����"�5��Le��O�ԋ뗲{��%�X���6�1�8�5b�?y|��f�Y��ێ����5Fu�tT�wp�Ƞve?.H��z)l�Z�pZ���OI�к�w��+���M�\lc���֑}������ъ����T��P�.�k��2�?x��\��v٬@t�0�ؙ)����b�/U<��`�(فi�{�AE�E��e���̋���n����X͗��l�Xs0@9��u
��b���57����ɷ��^�����n13]��F���uo&��Oca��PҼ��0$_eݾ*%��(]A`gN���S����q��D8�-���r�C�ƌ�O������ �r�Z7 b�tf�w��o�����@��8����ql�z��9��B'X��~z;�T\:��h=+^YL[Z����[�o՝�j��k�F5>.�����6�&5X2��C��=��&�b?�,�0����1og6�#2��-+^N!�Q��s�*^+Z��;����N�f�}F�U �Ny�x���^z�T��xmU�������}�7|7�Q�{��܋�F�Ji"G*�{�>�Ⱦ�=���lHZGw\�ĉ�
ܗ6縓�)����2�z��9w-�D<�<�[*H��;pձD=�J�3�����D�������S�3�RQ�Lv6�>M�X�.Yr��!���$za(�uò����%��F����C�_�9���P�\���65[�Bu�9�Z;1(h_������U�{Ǌ�&>E����B��cMN����pM���M5q��[V)�7�۾�\�WL
��.��R�6������l���r�e���4i����,�gƹ��Ɛ��/u&&dn�X{�u�c�6-)ɂ��Z�����IJ^>�z�L��a��`'��� G�wy�y���Csp���;�Jin3_�2`y�Q�,yEط�u�5#r�n1�d�F��~WL�6�Z/K��+�.�F�у���*�罶Es�=^dz]��,U鿈�\��ކw�9�:e�Ϻ�fK֮Z�ڵHX}���2�-'-fn����w���!��gIDW���Px�]��^�Ejp�����Ry�Fu�_XYFf��:P�����/���
�]�P�V �q�M.�P����'*�<������T�����9����jo�C���x�B�d}�f��/�E�WX:��TsM�^̬��A
a1 n������Mp�k)C��݊k]��2�\[�b�7\ż@;�f<W�Ԧ�������҆�s:���
��G��[��"A�{m>=B�&�a��r忑%�}$��{)m�Om>; �N�ݓ5e͖D�;5��B;�uwY�=)�.�+5��Wi�(%��:��:�e֠���V���7UX���4�=��9^������
q��>�x�T�#�#4�]�0ɽ�covv���TLZ����*.-�l3��ey2ϳ���}
��}��Tz��v�����{��ڸ���R�){عt���{n �WڡJU�4uڙ��_<`(K�`ڥ�Y�l����%� ��ȏ�� 4���%��9% d��BUU�YJ9	�9d�@Rd���AH�E)B�d�TS��-"d�	��@c%.I��9��S��e�JQB� Rd���B�Y�-%NU�9%UR�d��9d�)��Je����+�d�Td�B�C@9f9dDI��T4�d�@�TY�fa�NYA����S����bё@d.Bd�!��eY(ђ�)��Vbf�d�EIY�!6H�R�R�HeAK@Q}DQ4y%��=�h�V�7�,4��0�2_�g^2rM�O*���xo�����=�
�k��=�pe,>��f�x��>���'Ï�����`��j3X��[*�x�;�I?�W�:�o�p(���t��2����޳2�Ξ�X��֠���=�)��˦�yԙ*d�{e$���7b��#����ֺ�f�Ѵ��<�h��,�^+�g�Q_9p����.����#z���/&�;�/��2T�I[ҽi�'g`����g`�U��x�	3�%n��n��	���w�������^��D0�Ih����������_��fml�h~�Rx<�(f��r���g�'�N$(��Ux#5Az���u���:(^Ip�S�>�skK5�����yԡ��iɽ��q�3�+K�J���W�af-��֨V�g�sW��C���t8�Ҟ��S��3���ǳ3�u�C��,d�o�$���(h4���ٓ}<sIοem��	.���ZTA�jZNٵ���������{��WY�Yr���v�ݑ���uLG^9�@�����x*b�t�iv�"���KL�L�{ܰ�
i>���<��K�8�]���u�����e8�mwN�;���~��c���Wk"oS�᝻т������탆�E:��j�|����R3�/�!�Q9B3l��5�zޫ�U��;p>�i������}����YB����6/"��eLPb!Enua캞�����yr���!��d�=��(E`�Zr��Cd���]�Ľ�x���p��A��3�c��9�~��I���qߞ�Y7�-{����g��{ ��憟dB�������*w���N}%6�1n\���r��J�~��=*���X�v˭K>�dz�������~\f��c_�Y�L���j�I\�_�A���;�����
��O�s�.����G����}���m��s��m �����G�T_��m{�� �}�>�D����nL���D�J�Au�K�FD�S
B��zS�ӻ�t�G��=��ʊ�l�fDM��I�҉�����G�^B2S�¥3�
�b��VOg��K����>}O����v� L���
7�s6_���*nn8:j�:R�T��#I������b�=��Q�w�O�[�%xXF�{�ĳ�O[=���N�zz#�0Xw��L�4��.�a�5��ݬ*�p�yiX��|�fxPĬdwr	z���t*f\W�Â���˶�<�y�MG)���������ltM
}�I��-�L�;�+��f�*N��4�6ӻU'f��L��Jur��p�8��J��J<��k�ⷋ���&*�J�}9B��.���8���ZB^��\{�ƾ�*B���һ!�'�Ү��~�L��4�CqeiV�}R#�զ|x���Z�ݻ������ݾ(��C��w���}���?X�їK���h*ٞ�����)��ONM�9�o�I={DZܱ�*�hNO�N!n[����`w��(���[�U�c�Ι�/O9���<������C$����'��4<ؗ�7�m[>I��Y�by磮�W��:c�4�Yv3+n%�P�pۆ��ܔ7�} �i�����T	=���g��+n^��N׊� ��q��R�%ڧ�� d�s�3��,v/U)}�Y/w=�ނ��m�t�i�07�@�JMpJ�>��|h;l�6�^�n���V�5���aW��Y�a�rQeu{�0��Vl}���c����tZJ&}�UC��P%�Z���Y��7.�!}��ލ��;֍����0�Z�j�	��I���L��]����K,F��V
}��zd�8���v:��W�b�Q,������u�ؿ��,��m�!k�dv����5��^z���x�^rV�i]��D�Go�nӎ���s_l�]J:�X���f1����=��huT�M��������lǳ�w����o�B���-�F�{C��حvK2�Ҷ�ϽN�����M���,*�Xa�7Y5NL�N]`J!3tћ�u��0!��K���D��;�	U��Â��(��XlÀ:��G���	�/�{Z��g�1-Qć�T��;롣ҁ5�b���u`��s�G5��}=���]��h��>?1��lz�x��G>����T���Ya]e'���;|��l�?J"���9�h&Γ��8��؄�=�����G��o���B��.:dE�x�,���٤lz�&�{�efpnۅ��W��傼f��Z���_*T*��SB!-����E�d�sR;�]��<�\�K��ؚ��S����3����Zpy�t�f�d�w��:�MA �����LŃ�e�N�:��8�z��C�����L�p�N���i�y�N��s8�U���>����1�UW�)��.uB\�xM5�n9��N"�wW�%���-��u�U��>�v�`I�ՕT̟4�k�.�X���;��߶1]�G��4d܆�(�ӑ�A���P�3)�Q{ɊL����T;�맫��U��c�|
�J�#p1����9[)�Ko��EW�#s٫�attK�to;��Ⴁ�x�ۼzyJ;���c9�5�E�<��c�7Rĕ�'�}} �E�J[���=^8�[@�ʭ���E#��)�#;~+�̨m�J4�51�׹�c�e�b�f��F﬷����Vة�o�a�0�ʜ�=w@؎�;B\2R���.qh��k�Щ�۹�*O>ނ���w|^}+��Ľ��}�-��f��@_
Ԯ�j��w�m���s���E�@u��3�_gŚ�p��]��PߕD϶�a0�3"�g��{�8��y�^�^�>"^n���\q��F��/��v��}�<1Їn�`�����R��ud�O%݂�yM@�p�.��j:���WƱ%���k�s��j��ɲj)�+{s�l�}>�<I�e�86�tf|z�lw�q��h�>�\�� ��hm-�wt���[O���z��Y�uX�ٖp5⼦rD`g��E\"v�4O�����z&������AU� ��%y�$�L�5�i��͔�{"���u�ϕ���Þ����[�{�*-}����<'����!����=cuy����z����|孕��K�~���w��CM�'V)��'�cL_�OuT����P��%�=�w㺜ՁY��e^�W�iM~��ʏ�������5������OM����������t��疊[��^������5�$�weu��ٶ�@»1>.���_#x˽������kzw,cK���9�:�/j[����7�.���X��b�\��)�ǳ���gtX�8��G�V��hoLK�7�����%���[ٜ}�.j�1�{I'.����ux�{�\�����=X�V�v��^�~��X�d��BM���e`P�i�ԷLŷ��ޓ�}'Q�ǳ�����L�^2-;�[�ͺ����Vw>�\f\�]���6<�?.�{��zӗ�4g>i�޴r����C=M��f����!���`�O��ԫ��u-3�V!7���8���ji�I���~<�^[���DO7Y��=�N̠E�`�I�L/)�-�K+Y��+��|�h�j����)���瓞Q�3fC��3:_�qY7��y�u<�X�o�&�a
���4%��sV)L���|xH�h�y�C���baL�]̉���z.jX������%­+�)��E�㾿)���m>U�M;g֢�^��Ź��*�;ѭ��K�p���傟�Ò��YW���R\v ����f��>�^���m�:|V/�]�s�4TՀT��ʤ�����ʕ�n��eC�
�������k���j����W���*�8E;;����z����f�K7B�J�hɡ/wS;8�1Pm���Β�Bڕ���h�('e�N��v$�WkV�z�g�T�$o%Zj�݁T$�mYs��x���Ar�d㝎f����\|+�6�EOy�7���M�)�lt�}rz�O�^Bx4i�(��U���� Oǯ����{��cձWggǅ�z��W��"��,,�Bnn9�V��AJ����ٻ=�v-=�|5g�v���&��%�Lgޡ��p�{�Ľ2��������//˱�~��gHG�Eym�z����g۵�Cy�p!��j��7�j���
17R^$��K�X%嗇�m��MX%g�j)�9�<!�g���F}k�4pB�M`Du������3���C�Eڼ2K���4�����Z������"?��!SC��ߛ�Q���Jz�*n�ʜ��t�δb�����F|��`��6���l�{�ů�_��ܩ}F������T1g�rX�	s��8��Q�vAw�6j�!�z��|Vr�x���yqI��n�Ϫ_%y�3}�ۆ��g���5�`�i��Y���:��:��޿[���ęZ�,��A2�Rb����)��NwG����_]��?ux������Q��|/�� �%5����*84Lb�l������ZT��BQ�I�O<�k��=���G���5h�2E�t������>�0���-��^��l#!I��Wå)���B��s�:��nȈX�yT:��[��+Mwf�z�'�ù���Z��n}�@��-4pԁd{��A�=V�=�|&�_�do����a6�����<W�q�P��Wbs��{%Q䠩L�
f��l�%��w�p�'9��~�bS*���;�)�=ࡖ�j�`���e$/��V�ʔ���y�4N,?]���WMk��%�}�U���I��:��s���s���n���Fō�[b������j[=�G�DM�կ��s	W��S���P�ic�z�a|��U��f �<��;��۾د|�4��2|v������E��f�*�ܦ�� ϊ��{}W+��[5-o!��J��{��iY,�3}�g^#���C5V=q<Z:֗�ʞ=�5L"����*0r}���g��}���� �� �_�9g�|�����1�)^��隽��5Ƣ*{Ά۪�4T��O�����_���#�=.B�OL�w����~{4m�׎�ˤ
�p잵:�gn?S��{�_��>�\�ͦc�vr:�9�������'�i���U�>�;t*'B^|��ݳ<���[^v<�
}��a�8���3���v����ж��iVG�f�����Dr�+G��0�`q!b�8[B�d% �H�ǘ'�d�gt��&d��i�{k�W o���|��iC��TËj�woZ��R���L���#�x��������T1g�l��b��Rǎ8�j��p��ybM��u蝙�Pk's����V��R�Ni�B�!�g/����k��o��T8����q����~Ә��sr^��WC6���栾��T��UCz�������}�<Z<�V��g��I�4߱zV��i��ψ�k:�̨�s�,aP�Y�U32��x+*Z;'�dm���3�G�l������c˜��0�ʜ�=w@�*$���3�(S3�)c���}}���wr|�di�u{z]�0	\Уs6Oi����	a�M���7�`��i���f�.�}�[�󼺕�)�9��䙟d��/�J��^�����Bߗ�.�3#���g��%�ҳ8=wu�������o��lc���V�<�#�����Y�(��^�g�M
0|�S}�ݹ0�3�+�e�;�{�Z-3���>�C�ߕbI�ڼ+eW�B�іs�׋ˌ;��3K�����˨p^�Ja��c�Cq�rd��k3���yD��X��%U�_h �m��X"7�oVJGo��4ѕ+�s����{������rD���9�[ӡ'Uj��k�H�_�;*�bz���6g�����`>/�[r�w��ti��U��F�ݞ*o�ծs�FFU>�*������n���|_jz�`п���-jYҎ��\�N6�h$d9K���*����8�/��b�Hv����l�<��)�ZU�J�I&[Ҽ#���{�[��򳥃�V�x��	�!U33��S��߱Ct.僶����DNt��OX�N/���Y϶oVp6��=sj�߳v�^�~���Ϫ�"�����DŏWc��/|z(���\#|-ߎ�����p����ڧ�gn�`���:��^:���P�}A�b�Q`�����3�.j�%�{�L��ٖ�� �G�
ۚ>����g�x�=2����	7��Ų�ˢ��w���M��/�S�����'>�aT�C�i߆v9��=f�rc"+G���^�F�}��>�$O��NS�(�A6��yU����*oW�45ੈCiӤ�%���J��S:�w�p����kc����V�%c�L�y2��{�h�'?I����=�ve,��9���v���L��ͯAB�;�v�ʔ��)L��\??�s�8&l�s�L�s�G����c'�����VPVs�PhWKT��l���,>��`��]n�����i�1bQJ��j�KwktFj�3.�)�pc�h���׀��OxЯ�sf����L��S[ln<<��py��2�s�i'�5ft�;k����1�(т#:MR�_Q���=�����X;�l�+_��؍��A�6��m:%����=�<(�-�O��}�T�W5���P�a��٤$�IM��ua}I�\`�0�4�PW�5��@U�q����8��ɂ�Z.�s�<K�S�{5�<�<c鳚&�y��Mp�2��S����~X��ݜ�#+��y3��.���L�q�nG	��1r��j��f�9�"���V�=D[9q�U�r������F�e�����4��qQ�Ou
��ם��ԮJ�J���2��psqV�/�!�s�P��FU���|leۓb�Dd��={�35)Sթ>���Ȥ*�3u��!�}BuY���a��3[� �ydH����\�.
U�]a��+c�w�G��/^�=�qv׮�o�Zτ��cTq�S�@i�'���r [um�V���y��gD��[S���ٌ��g�oSr���/t��֟}��o
{��,� �SeI�]϶ھ[���GI�R�yߩ���{k�<ia�u�}{P��Od^�]WH�:.>i4�d��aa1���D�b�.Թ֧�dϞ�ݫh�RC�Ճi�c's?q�a���s��Ó0-�ZSJ�!ta��e~��8E����1xH#�|2E=ǉ���ќc$�DJ��7_f`��
*'��`v��+a��D��Զ3��8�u	Ҕ�	;�ϒ�^�V� !ݎ0R�B����G�a�g<g��n�q�nP�|T�z���m���7���K��N�L}��M�0�� �;švI��!�n��!z
obHL�1@��v�|^9HY�T�<��͔	fe�s���'ŜqVuL�`���b�Ym���ge�v���<��7;���E�$�8�q�w��ƕ�_\/��u��;��D��}4�{�C����	�зI�)EC��N�f���3����t {����}Ő��4��e��-[V'f�Ⱥ�
�Z�[��oM;�zZ�l�jH�$�2�B�]�|� '5���"������Zy]��|j�鬳��V�sE�vF�C1)uin�{�A-�vچa��}�c#�����Y�q�uX�b���h���5�����CxD�e�Z"8��Y�n��`I�#W|d�(�.�P��a�7[��X���Msq�s�_I�:I�q�O@�a>���j�G�ʲ^�\��0�r�^Q����o���j�6��M"��5|� E	)I���q��}�Wё�� a.���}�}��f��K����Hu7�%�*�hY�vk�+����2����|h�ݛ�eH޽T����N�جW{z��g�۔L�b�a�d}}����w���1
�"�J��k�8A��D4�QH�e����	�T�4�cAe�A���K��AH�#ETPY9NBдP� R�CKY!DH�P��HӒd�FJd�Sf#FA
�bRd�c�	J�6`�aHDa d4VFT��Y"R�99 ��%BDdd%��FTU���9�R�Q&YY����Ӓd�Ő�NHd!Ed�X�Q��e�E%+KKJ�aE"U%	��PPR1+�P����ͣm\9�l��;���?^3;`7�4����=��%�F�=s���S��䭢���]�Wm�!O=�h�o84scW���=��&�!��t^ƃ�뚌L�wή9#��%�Ź����.��%�+��r��QfK�p�;`���洙Ip�EЮ�x:�t����g��5�[߳Z&uJ���ޣv��u1p�brʞJˤ�r�J�:CK��7 ��F-��_�k�N�{��V�|�y��F�rTՂ�f	�t�8���ʕ�n���;�#6�&q�Q�����;��JEP�L��q��p&IߺQ>�=x'���!<ѧ���^]�R�voc��=�E�ܖ�="�Z���U���(ߺL'>az�t�E	��,�l{A㔖c��؆����L4��_f��oœ]e����^Tǁ�s���S:��U9ݶ�ɍ��D1cՖ��#yդ�f꺧��f��|t�1i��f���MM�2�o6��[	éA�-���|p3�N�:�^;\�����e�x��8�L$�ʹ�Ų����kl��콼�s'/�EڮJӼ-�i�g���i{~�z�.�y�G��_1~/�G{����DE�t����RH*��N+\.Q�������C�
yrhacb
��u$������S���ݔV�7���9t�|�L���Vpaݶ�Jڱաa�:���������1�����lt�#���ަ��3�W��t����ܷ��L�Ol=�NmN�9���{�D��y�C���Ѳ��G|4ɱ{}�N��M�O�|�<e�2��	��}��S]xGP���~(«n������º���A�.#֑��v;;��:�o�ۆ��g������p��2?Z��B0�v�KXK=����\����h!ŞHw��}�K�1z(`��(�����`kj����О�5�[�sk�+����U������E���2�8���	q��4u��ѫޠg��ՐR9��zJ�+��a���X�,<�(��]�}R�ܬ?�3�����1��c����@FϽՒ�� ���P�\}2���]+�qN��_)yp�����e��ٞ{K��f���Rʫ�h��^���b��="Q��y�^�!��������ܳӠ��4e��=�\���߽���t���"��r��=G�tJ��}��[�4l�n�����F�Ap�q<�����}j�ܣ�@WV�ߤ��^	Gƽ��Ѭ����Ĩt��pi>��<l	D��S{Ef�3�Ύ/z�"��Eӆ�D�z��-��R/�m�bJ��6f���`�}�zE�n��^��&��g:xEVppb�=��[���֫7����C�#V\��m�����HWS��Z�����s������a9l�m����lU�Jр�lu��Uh�[E���G��
��@3|�9Ф9�e�X5�=M����_*���	��3;[Ր|�ذ�ڦ�μ�^o��-�~f�<��S��ŝF��%��T���us[�5���{����,�Z�2{�ku�8�N�k�^�V,�G�Ͻ��i�a��>���l���	���'�iӛU�=H�������_�s�"F��[C��C�Vˀ纙�6ٖ;����<q�sWh�p��uF}�����e�'g�[b��ίϪ��`�C���� u��i����6\���1����TS�;�f���w@I_y�'gk�6��*Z�|*��I&f�QuO��:'�M��W/�kcY���39|��oü�d�t~~�G�˨��E�T/VUS3���v!�qG��{I{^#�93��gL������.s�>���*rDt��䨓���Vu��Ya.��ӷ��B����I-�\F����f}+�e���-�ό����"��f�.�*�eɷ���L�]���.�[���Ń�8#��dԽ���j�hڀm���-�����a9���\�w|���,�T�$��T�y�K����L���e}�CӼ|o�΂\;w��<�?3["������AZ��0xݵݪ�M�ֹ%�
�M���������h�l_�׻�U���.��C~W�d�q;�aL�����ږ�HO�5z���iX)>[y��|�
�F:Z�eiӝU�x|�\� Tt=�|G4�[�B�)\���xJ�!���m�H�n5)�ot?(���m���"�J��==2�_f�����棫DY:l�P�]%0����GG���]>���cOT���E�ʮo�֦4��� ;�r�Z����'o��#��9��B���Rm��tf77���ڳQ�{->2��6L%_��H�2ޕ�-S��^��Z��,j~�%ZZ�j��A{����k�Gl�-9hzӋ����^0�D����E�^[M�U��sܸ��Kk�w'�޻�������7��B���y�d"�����c�\]����}��Y%B�9�}��F[�-��ћnT�e�\�=��;�����R�ꮠ���+�j��c6�i�ǱN�'L/a�{�&�24e��s�실�;����ՋC�)�c%�B��&�.-�o����+wA�,!1}�0C��͘�����mx��y�t�.G2�s�R��ף�����eS�4.�ۤ�����^]����l���KJTZz����3���t��}����e�%#�o�kXs��8�I��$�N�Xcy����^����"ʆ���
��p�7������\��{.LlEh�r�r>^\X�mWyl��鳷��>�F}�C|��(e�N���9���*oW�f�����������6J�6�K3�2)#�~�:SF���pE�Ļ��W>�Ýc��G����DO7Y;n�N��GdU�x�Q�ƽ��ٞ�WJ��D�+*M;֙Q<Z�{Ϯ�NyF^ˇ�-��������];Z��ج��H���Z:+�4uO-R��y�æN�wx���T�*m���G\�e���xc�p������'�Ur[T��/��d���O�<=��b�;�c[2h�(�s%�=�w��|�`ӝ*b��X������%�9B�%u+��L�><����Q_�>�X��b��Z��������<�TC�H�o�*jʙ�'��z�(pF�����2{���5�4�^�Q�+�^]��Ȃ����C���렦I�҉��V&��^BnG�۳;��kg*B��\L���otW^�tw��J��
7��L'X^�҉ �.�T���d��3��2b">�v��j�"�#�,��[
�\���{w�uƁ}�j�TXa�d�e_A-�V�O�{
y/[�r�Wym�cn}��lBe�f膜r��23�Y�K���9�1]�Q���;�_fE�aƠ������w�k<O�VߪF�/������Y��[�d�YAh�B�-���w���;�GM�x*������|�|�X��<����0��-oV���P�ͨ�i_�C���`j�Jz"��l��>y/�i�g��l�|~�p�	���j�4/8U��ᱎ�#x-em���=:{��z�h�&|13�.^{�s'!�E�O$�=��i��m��N��~�s0�}$i�F�ר7+ډϽ��Y�ȡ����'K��~�=����	�oﲯ���i�'���{F��a}H�ƕ��8��{��c)�73k��|�~������Z��	>�lF�]�/f���^��%�e����a�;���P���0؞}�s�(sS���ib������N�L3mT:�+�������b`�=��A��z�9���m���+T�U�Fv;d^/��٦��u@�2KM��^�"�����U�t���h�~�����,o�S�u��S�q��e=���X�,<�(���Qpȩxn�}���x�u2���<��<���Lyn6��L
B�L<q�w��ݗ��Ӟ���k�縔�����ͳ�7�hS�9��b�*f�:�����wB��	���Lc����m.�nL�.��
�Z����<Ǜ�������>ĩ��u�����P�\	�����G ���x��t�Vu�>�彈q�c���a<�e}~V��j�|j���1W��Lö*]����-4�44�gͰGC��k�7�c��4��pw1�K�E)��Or{�	ŏP}�]��{�IW�devu���=�ĸ�2���k҆�������t�:�'����K�@+�hp���r���zqcI��3�:��0�7;ٖpE�<},����ִ�~_<z=V�7�4��t�=��|=^��AO�̉8�-}|����Y���cO��1�ؠj�:�*�OF��]�=�� �|�׼-�sc�#�=�!C��w-r��/:���u�<��"
�ˌ�����3�����ydT`:=�"9�̷s0��ؚ�	���������#����4�.<����w������а�����l��3�f];���T��;���mJ��5�_Oj3�����|4�鲳ǴUu��J�c�b�j%\�Y�f.j�jn^��Q�E��u�Գ���:�q���rk/�!��a43�m��ky����NњWw��1��������n���	�tua�,�3�0*m�D��x�G���'0�0<6
2�kV��'Y ��Oxa�;%N�()um}��;��	F^(�}�p��^�¶NO~3w�>5��ˇ�;�p�j-�T7�*�����O���x��7�]��<�u�w��A���!��z��A�W�g��eE�'.�
��ʪf`�v[:1
�	�;IFL��k��^�1E�����U�g:��a畓��&�P6�`��Fl>AV��n���k�����;�R���٘%sB��3d��h�o�B��(Uט�w
�[����Ћٮ���O�.��|՘e/�O�S�{e�<pE�^d�pp"�
>*2�ʗ|�gp���Y9-��o[����5�t�_�+N�U�x5�9fM���Z𻁹e���ا�L-ZD]x��#�m�g���+�ּu?�ʱ%Z3�<,#�c��t��nN]���\n�8:Qk�9d�f]C�:��SQ#�p�n5��L��g��Y7�N^ĺ�&����oէ�$��PQ�r�Z�xZ�D�
�0`�����%d^Fn��ɽ~�mlt4��za�*k}+J�s	V��H�2ޕ^];݂����d�;w1%ʳ�_c�Ħ���R��q�s֬�\$z�l���A}+y'���q�����&euE{��K���r���|�rCo:�v,�\w�������d�g�_ ��/�nkH�y����v��#�#}�x�MxmTi�}�k%ҙ�{�U��υ&r�����,g�^2�DO����g����oˆ�>���ŠQ��E�����cݹ�S�#z��Ux���
N��U��:�����lX�]��rE�[��^�`�썟���\����7��/��+�J��z�/����o��_NK�j`��Zl��E����Sɼעfٗ��O3�ٖ{�k��Q2������z�(㾛q����{zߏ�Pj�_Ʀ�x;��8�:Бx�i��Q�=�)rce"�z�?�"J�^��Z�p�b�$;�^�*�uޝ�<Bs�����z3C^T�!��:Leb�R�AWy���2u���U��u&TM,���\zc��GN~"y��;n�X��]�6�b��o���\��@�<G��>^ϨP�y}i�)�`R��x>�~��򌽗mK.�����xh�����F����v�?3�B�A��sV)L��\:Voi�Rrc���t4Np���.�����^g>��[<֓>K�Z?p˞�8���x=1]�z�,3��Ң��]7���רP���hծ����_�5�����$^�.�hƥ�yJ\�'��݁��Y����<��v]�k}w&F2�T�碝d�M��vH:�Cu��`�Cؒ6��Y�*��:�ϫV���d�|	O/N�+46�^<�Ju�%L\<>�br�S���Yt��P��]J�*�S:��.u^�R72v�z^�ϏN�N��:ڕ�����5w��4�R���IC�O�ה���]ߦW�<bc_���gDg��D=2ϗ��d���bO^	������FVx�{�z���/T��δ���Xu"�����G�W����ހ`�Ի,h�����ߗ�n�L� ��kl��ו�Z�h_&�����ɮ���1�2-�>7�ԫ7��8싷Ѭ�'% o��%�\Q�?nY��3��>��>S�+��ajv�亣���ڷ�v=>چ%dwr��8έ9��R��L�ZVʅF;�W�n����.y��9L�'�:��$���+w��>�˙�U���٥A�j�m4��R�f��<4�^���'>�ͦE���S�CӦ�v?��\g����C�Io����2���`�����Cz��ډ?:�,��.Ka���g�N55Տ��MT)r�Ĩ7����Q4����` Ѿ��N�cn�H�;~��3�,����u����/`��BH��Ѫ"�)0t�M���3�5_S�9��e�w���)y�7dn��-��\�!�;`:ᯈsռ��y�{v�+��z���2r/*𺱩�3������t7���:W��ۧ=g�{����Dԕ��t�P�qq�˫�[����9+��)g��~�*�i��\�u�<��a���s�;��]r�=�b8t�(���D�v�m7c�9��pPLx��ut퍰�W�z�K����l[�r<����Yɘ����-6���8�:5�=�����'���]����iv�vt���-�`Uͳ�ŜﴅK��i^�&��
q���ӌ�Y���=���9%�ϯ8+ˮ�f��{��;�cq��SdC� H��j�nL��.mJ>9o��V���N�ݐqֈ�u�*n�7��
�b�q�ebV�ΐZ� �6&r�_^	���>���J5.��kY�G2���1�5���v���Nn�P6�EwV:�����7�"P�տe2����n]���t�ݥ]�:O�LFl5�����哘'����ǌ=$�: }^h����V��ͤ�D"�z�`��&5��v�9�yn���5.;�X�K}+�6�!�M�fn�SD�;�$F�.�Ŧ5Y��[��/?h��w!L�z���a���[�sX��d2h^���ו��4v��Ò�,�9lW_ig������v�0�҅%�2��~d=ݽ.��I)3-b:70r��֊i��m�8�2��m�0Q=�P�B���ˮ�R��B����/�[!=�g#�p8���p�N�:Ԭuܑ��t���,@��&��5ǰ�X���z�S+�;�&o��.�o]��#����w��L�w�R�	5���O�R�Wu}m>c�M�w�9�i�X7Hv��O���Mx8_���q,�%�wBMK2ͯ~��`�$`��(��9^�>�T�w�-˻X��# �����ǔ�Xّ��:���Ng��xH:v������w�L>�}����+"_p�7�r��ƽ4]>���c_L偝���W	Z��,	-sXRRg囵�䮽�Q#�,�od�a�V��[G��'i��ƌ�����kk������+5����,�(`��*8^��Ɣ� x^C���K(U�l�rnV�ΐνyPz��o �}�c]y���@��Su�R�)=/g`Ǿz�pe�Q��]S'�R9���w�̱�3��`��
k~���-����|W��6����~qXa�)zu�ΐ�0�$��0}X�Љ���Ay��O�-;������oI�d��Z\Ooh(Y�=�!<P���c׶��g��*z�6�-��$�V�ʁ⭑�ٵr{\8�.�D��!	*6�B�� �H��n�������/䢖��
)j�

X�3*�"
h
hi��
)
�Z&(�2��
�(�L����"�����)i��
���$� Ƞ(��J����(JP��(%hj(��"�Z*�����(��!)���("G'��h�	��r\������(
bh��"������J

J*��*����
��"$)h0����b2C� ����*(h(
��*� �0�
i(JZ�0ɠ(*����"��h��$�!�h�B��11"	������׺����X��SL�d�gq9�\��/?o���5оd���:e�0n;�I-�0�Bg'��o�oY�����m�9q�{K�f���w⎛M�`�I��H�j�˱�)�%cΡ��.y�Y�Ew�m�({�g���a������d�6�C�&W#eC��C�����}�$�O+�fnd�>�}���z8<�����򌾮"ܭ=��Mq{u@�t�
��Ϩ'�S�.msj;]T~�<�z(�V����9�R]31Nu�&WOP�-u�sE���(�-�
�κ�u�-�Ɗ����P� ��'��-8i�c�x�ü���j�L�t�^�Nݨ��/�W�M�t����;�{G�Rf� |�νJ`��*����U�9�fg��<��_c������ ���u����>�S~�1�O��K���U�䊎|��o�O�Qɗ�fs$.�������6ai+BoǨ��>��'��u�Ig�Pl����
_��mlgn�˞~���;Szks�6Y�Ϸ���#T�(Ò�᷊���͙�&
�GO]��J���Nׁ�B�^��� {ؼ 
�{�?(r�Ϟ�}�I��0�o*�A��E���@�u��e�v�P���\PJ�����grȞ�+�Ŕ<�:�{G�� ]�"�|o#�q���__�aa�ZՃ��h�,�/o�^��3l�`�q�~.�%�>F[V�+��U\���d�u��� �w{��9jen��� ��9�h~#��6G��!A�zgr��sA�W����VG^q�-kb�������k�8-����56�+�f�{jDp�c�vs�GbjeN�s�Ǻɼ魋��C�|ϟ(�ڧb���Ӄ��е(y_� ![-���Lśl��b�����ͣ�UAX��\���{�ۻ�Hr\y��W���~®:���>�C�L!�j%��k)�V]��"�ߢ�����r���i�-�5>+��d;���J��ԡ�-����.��I�U۾�.'ۉT����v=i�Wr���d8���W#`X{��TEʣՕT̾ͺ���vkw�O=2�Ԥԕl4�.�_p�ٷJt~�PX�ו�N�G_�s(TI�KK[(�n�W瞞�o���򥣜\�O��P3�a�v̋�zf��>ܖ�dXlfo��5�'����@��5�'�pP�e��҆�un�R����l���t����E����Ea�{Du��]vO�79�W�uST�梟(t�[��˲|{�9(�����QX�V�Cb��>5��cC��U��|%r�1h=���)���YH!^~�g��5�3�2.;�Z�sme�8�&��6��ʾx�pz�]����:_�M�G��5��>�3la{J�H�'B�t�[6�}vv�dh�ge��d�Ptg�J���&�Z6dC��|7���x����2;���^����7ª�v�!�Wpr�\09d��^�V�>�Pp�e���5�RɵWz3o�V셲�A��ua�l��{`���QkR�:Q�I��9�~K�`�H��h�^~�2Y����4�_��sޫ��x��0�y�$��-�Q�g�1�ee�G.:FK� ���谱�P�/��b�G�?�[>�*�1�1X�DO��t���P���i�z�P�L�p�m����?9����9���euҿ]�p����u���=P�v_{�n��6�)�-��+����_�ub�z3��ұ����S�]A����]��g���m������VL�����^~����<>�K��+���m�-L^\�����{9�Zȼ�>S��j��PKr���{A��sT��'�i�tߝG���rcg��M���y߽ٻo6���/l����H����ɗ�v�	Ά}�)�W���ו1M	�Xe5i�z��p��Dh�<��ѓ�0�x�����/=Z��p�,���<s��m��I=���F�\�&�gN9P[��pZօ���-0�%�		�x*���cv˸�[2ðS�O]{1�i�����̚}����0��[V�ǮP�!3d�B�}�hr
*�(�o�"�t��3�R��]_�
�k�8�8��N~�"y����T+J�����f���fP"�B6|��P��+�3��?#=��!����(�g�Ťݮ|��M�x��;ƴ?U�F�]�Y6t�I����8�v3�j��3�n���Sގ^���H��l��WTž��[9�'�UrI22���Ca�y%J�E���.���-]i��m:t=�,��>��.�L�9`<.�V]%c�(�V*W\���N�]�u�/x��X���ӊ�׫(6φϸ�������Yϗ����m��V��m-�K���ù�¼>��9M�T
��]��� ���Xt?z� �{6�˽xl;Qy�w��T�|�!^U\B�1yp�����U�Եp���`*��(��I���u�݇�^�o�S�% ZO���L���ͺ��B�B|:��7�K~,��4���VR��5�Z�Z�z��f���VG��iOO[<�*66-;��Õ[�sT�|3u]8���Cq<�/ϕt���>�17p;Lob��z��5|Wcʒ���D�*՗=���W��dkr�ڒ�9�"�k��fY���>����t���l��wi^��~9R�A��V�⫔�
�y��0��^��}v	�awOu�sy��sv�ؓj���u��a�]��'R���t��,����&�y��W��=�~~��gV�(u*���&p#��K����v�^�oI������If�pz��M�..��w����P2.��e���.���%Ӳd�o���Y�����;�u�d�zU�����9���������NmN�9֌B�eg�x-w]O~�;��o�9����F�
T6`���ƢX�1A�XX�	s����g,[�%/)z/m�0I��t�O]���ڶ���#Z�T9:�y�3|6����oٖ�{}/��I��<��f>���5ϥ���7Á&W#`�x�qvR�v"o��^,�;ϔg}:���|�}8��.��|_��4�v]c$��ρP�YA;��O�e��X�,�����6i�S�,��m{`S�q��e2��nh��	۔㖋K��_�.!+���Y޸r`�U*\5��P��l1���5���S<{�C-p8&T"��a��ܵ�;��߻�C�+�RB ;��K"g}�pk�XO(Y��h�V�����loQXl�fT��ƥ\����
���EO'�+<ba3�P�6\'��uv��b�~��G�{�y:�9��s�܌����/u�7Ɣm+�CF�������+�i<�0ْ�C�6�o���\��{lސH1ͨ���F�Ek������έo�Z˼�Qr��ϱB<���6���KÄv�%�+jr�U}�"�1���}��0x�8{�v���c�rF�iR<6�[<=?[A���W3F���'5���ՈP{4XV9�l��t�t؝��8g�W����Z:�U�u�Y�V�z޷Q��R��um��#��Ņ`g<���/���?(r�>{�i�U&��;V��ӣ=B�t<
��-������,GvG��u�P�OL�ZyoC���]�c����nw�ҷ�[,z�,�1�M���51�'׋�'6���fxGbjeN����,<瞔K��F��tj����v��e1줮�V�`��Lśl˧s(=��C��}M�.{�)D��l���z�}S0x�+<{EWZ��qLP��֢V1N,Yw�>�%����~�z����y)-���_{�2��\ۇ%KQjPז��fRDpy���g,�d{=������,�_�Ӳ�5�l�H��W�9�Qw�ˣ�z�|%G�w�{�Nt��W>yano$���!��:��i>�]�s�\��d�šGr��פ�0v��ƹW��$L\$5Ĥ�Y�|����|�Գ�vJg��1��&:;4(����P���n���᫬gG�7����-�t�F��c'�W���徵t+�/�d�������溽����P�5^^�S��ao�=C~Դ�s�˿�������i�b��fE�
2�x�d��h�[S)�!�:��Iu-h#۴"��$^��(S3Jպ�+��O���9�h��󮛳uw�K��\�����lCЁJ�y�#�q����j�-V6V�4�/x�4fo�wq�w�f��uڧ�
��%v�L�a�X�2!�Y�({n�����Ñ�ה��zM�����b��������Z�Y:l�P�]%0Y#��~���Gt��¤�(]�d�V�y���1k^f�����ᰑ��2�Y[4���c�����D��k�r�xD��xK��e�`7�a*ǝ�H���zTiyV�:���-�,y����/vtXX��xY�b#�
�}�/S�3� X^�ІU�[��xqW�H:��/cH�ܤ���u���l�;�ީF*�R�:�N������qxW'���������������<�]�q�ɩ4/3�59(h���qȮψ[,Ow�-����%�Y̿u�ɷx�[���sTb�V��9>�2�*yδu�Ä0��A�%;�Ț���I�Z��0\�s�4ˋ�zIۥ^o���P7Xf��Y%B=N��ɹ��Mu���K\��aԮ8_P`�=��Ε��J��gs��ER�+窅I�϶��P���=�}��t�;���mb���^\A��6��G3E�؋3 �G���.��T����}8�:׾2-;�[�ͺ�t���L�k<�n���/��/ȫ�ٕFǝ�ɗ�v�(Nt3�Sޯ}��{�}��ߖ��z�.�0/WR�I�^Eq��ZeD�ș��2�c��GN~mQ'z�
9N�<T�e��Dֺ�v�}�@�(C�|��(s����}R��)L��\ b�S×Z�nc��[6W^��r��s!�L�s�G�������'�{C��(63�j���!^��jf�7�M�tqϺ���;ej�9{=< �r�	�d��y�&R\*ѰC:��'���Η3��p��uruz����P�b,��$����X����Ò��.0��mt�o���_W�Y�S�v�V|z��khz-�CqC���|�4J��Ꙙ%��K�������i���C����R�YҒ�����[����0L$@�y^�Ȥ}S���k�в�锕"�ߔ�(���̝��y}��qql����mt��������V�t��Rĥ�s/���ⷻ.���/x�p�
��h�G��rΘ�}2�~�d���
U��|.σ��AU��O(�~ 8$�J�6����d#޾�Ԩ�*������lׯ�]f/.�M�XuR*�,�}�U��
h�L�)���1{�6t�� �u,��&�ೝ43^�fJ�Ɍ��tY5�PZ:���e�my��L{)u`�G��V�W{|���mxX���A��#V���	��1i�_��T�IY�}s�*v���Z�T#����v=�I�wry��%�x��:�c�ɒ�Z�!UO7L�ݰdV�z� ����U�gL���"�^�/�x[��NVE�ˑ��v����1(Z6q`>��=^�:�,�dP�{��r�6���s�gg��jĞ�+���h۞�i;�9vv�KlR��.�<o�u�:�,����8�ކ��(0�tK���'Ǟi�q���P��a��V�ę��֮��P�glWg�΄�X-��$'����3��vY�(sY��\��K%��n+�L�F�*7�qv���"��1?+�T}]7��Dh&����]��7����ހ�gg��le G��Q����S��G���R�i�{|^c��2=x��i�h��ؽ��\v�:���wgx`��\�wi+�9|����;���Q�;=WjK�����ߊB����}�[~��9@���������	�|E���xl�l����-4p�=s��j��vW����,�?�T"����A��?ޫ�({�^t���\e��C}2�9���۔�Kv�Ró�?T�'�MaI�b���a�=t�a�8z�A�L�3/��k�ɕ�AO�:&�d������&[��Ƿr�!�ʹ("g}�p���&p���:�)�C��\^!{=~^���_��ӤF^�fN��|b6,�[��F��g/�{iX�^e̹��Jմ=���N��@y�h)Q��0=GK'o�XlÁ�,BT:�q<U���D���"�4��x��^e�·�e{��ue'���谳�L'M��̳��<g�n�S7c*d׍��35�;��ӟ_��g���NｰXVsȓ�"Ը�'z���4��1�hZ�B߹=� aoY�s�yE��-�����<��s�qݑ���r3��;��\ӫآ}U�sY�c�[���X���� ��qs��=�"86�����Gbj �8o�gI�j��d&���lv
U���
h�\�𷆲ӵ����A�fP��r�s*�Ϸ����ʭW���N%J��H�E��ԡ�*>G�d�w���Z���!�!*{�1��\Z���wc��.�ۨ��|�b};)yO>P��e�?����W�6���,п��U����v=�����{���t�I��c	�% Ug�[VEp���VF�¤�,�us���R�r�Y���5hs��[�+��l6h[����rS�#zbX��ftЪ����.�y*��[G'j��r�|��)o=�e��k�o��Xl�`���\��JK�� �]6,�d濯7RռÍ,�G8:��z���^R��oWu6�f|0+�斫�8ٻU���<R�E,,�Pf�I�M���:��5mb�T�XDН����E�g�%��J����ƍ����	�'�bD���̾Kz�X�EpA�^/dW[�(�����F�����z�ndZ���W%�ւ��w
iwq�t��Fh�Nл�v2�;B[�*�>�c=�9z�=;����)@3XM��g��VeVa�mH!�I�����c���JR����\�ޘ��+9�߲�y�:��wqhx���)�/l�յeGz�^[�=�/lY,������e;2�vK�Ϯ���B�@�of�F����w�:w�j���؃�FP\mU�0���ug��d�&���KF�6�ܭ	ދ9�T��5`M�����ܸ�<���ih���x5���<�i�����`Vޖo��;K-Z}"�u��W`�l��xf�VM�Ը��l�[,p�(�9S슧P�����H�˷C��]/�7�7k��k�]=����_���.vp�jᕇ�J�x��&�4z��iݨo�
�IeI,�sI��%�w��P&��~�<>��Q	7�~�I
�|�R���V���n��X�*ւ!��m�w�6 ��G���ذ>Ԗs�{�8���g_�v�� Y��u�{�B,HW=O�� mB�CӤw����}��IP-Yڤ��A�>^��"�ü�7}M��[�n�UzuU���7Bˀ�c.�:�fj��w��"$�T��"΢�_�W�^���XK(�(8�
V�3��{)���[�_F���B�,�7A���Q��k�e��xw9�K�x��m�/�4#u �����k���=�P�D�zYk�E��o)��v
�A��e�e���W-�v]:�X��o
��������l}�H���wk��B��5�3��0�tPw�%���������`*�q>6�j�J�Y5��پ�e|�z��-wK������iFqwcg���܆�:=�P�r0��8�'nM����+#�KzTd�-"��@k�338����t�w]���'���e>�U:�1�"��9�/�j���V�{���ɣ�VNu"��Tt�&�z_;įv�;����h#�A�CMR�0PfeTfePP4QA@L4E�A��4�N@aA@T�%L�CC���MPQDDJe�%QAESMQ@QKKA�E RQML�e!M%R����K@PY��f`�KKT2Q�`�E�E4PQEfT�AQRPQSU�4�SfAER�PEDDf9Ya��UAM$AH�P9Y�EHD�T�QFY4�E.I�P�5D���MQS�fMTDE�EST�PY�d4�Af.M-P$�A$A ��fz�x��}=!�7�ѧ�U�(�`GXɝ�F�}k�,��&o+�Qf}�6��+.g$�^����͵/IQ<gU�.�kz��+�s����)�[[��Q��.cV8�l��3�fY~��<�*�����똏{��S��8�jힸ_T�;��+<{EWZ�C�L!��Q ^�,�6�ʪ�s`����MN�<D�P���z�8���d;���	R�[瑱�Y�U3=�L2����}�+���K4�qO,�m[��\��`�:F��{ s�Q*�s��z��z�\�;L̇x�$����ى�]2�!�V��+˜��yX'R#��ݮ�ly�5>۔�(=���s��A37)ڙ�W��ַG]�2W4(�͓�}���y�ꮃ��i�o5����X��a*���R|��є҆�ub��n}�l���q���R��ҷ�Ԩn����5�I�� ��ЁKg��b=�n�K��8�Or�b�ψ��m7:�I=<pf�éq���=PH*��P�l
��Á�+F���F��t\?z��g�w)�)Ӌ�_�l�������Ua�B;����Qk�9d��k*��z�pѵ6���-��
�pk�[��� Ktu n��]X'�4���j�ҽF��|�.{�%e^\^u�t�����+' {�I^Y�Qە�wguY:�O(�r5���<�,)=I�k�:�-,| lZ��:�i�,�Zo��g/��%�r!�����V�\�Y�?R����� +�l�b�-y-(�.�������J!3`�.+:� ���`��������N߇	Wi�ߍ��ހ|� �K�����V:�x��mL}2��O�o%=��e���/��}�^&XՆj���u�;ޙM������2�[M��c�}ϕm����Z{���I抰ȡ��타�D�p���}��<��G��h�=�pݝt������D�g)NU���v��%�OR��]к�k��ۙ8��R����}<N%�mK��0��{!�r�g�6e���\o�L��a<}P���칯<���A�dо�I��2�ˢ�Oh1Χ�Ҹ���l_�|��^�gh�K�����������"���d�Q�w΃��&]�s�'�����V��x�V7�/�2���V<yr=B�r"�tk���ɥ`zS#��e���8�%7ە=����=���?�}�&GS�T{���C`�f��V�Z��yu�|�m���\��s^P�Ԑ^�2� �p;�q�^���0��8r���qI|Y��WG���Jr�����R�H�l�_k�92^���֊���D1�M��w����H���)_�i׽$9ٳ<s8<�� eX�i���؛˷A��%��A#���S���muB�U3ވy�q̶s�G����y��&���VT��/+�p�1��E�ӳ�;��[��%\:p	�2��-��!ÀK�|<! _�<֓).h�}���S�1���Թ<T��������oS�C�Ř4���.,NR�T;+�IwM�������]����R�b���c
Ϗb�hhu�+yC����r��SU�}��~lbdd����s���~���C���c����P�>��e��!�x�����0��4��$$:�0oQ>��x yK��F��/.�߅��p���Y��X�w��*��j==��ܻ����L'>�ԺQ#D��zyz��	B����z�sÌ0�|��7�̾М�ُ��G{�F���X8s]4����^�T>:o��{��7�-oV �;�Uz�1�ۇh痞.��}r�^�����Ac�2+���ﶡ�du���էbJ�J��E˫���D�=Y��~�rX�6�WϽZa&����V3�\���L��G��s�}k�8i�s}1>�[;�ԣb��sha?^��sd�M�>��v�zjr�L[I-�X�z���b���L�r.J�u��Λ��S��ޫP�:��nA����n'}�gZ
d�5��4��߮!��7uI:�n:3l��Is~r,�W��g�̳��i~�R�ة��료�砸�A|�{����t|C���mO��>�{�k�|��Y���ٛ��$��u>�8���20'�X4�����*0]�x��Q+�Ρ�=p�A�\�K�}Juc~o��1tű�>�q���Cҫ
0�m[L�F��]��w�_�{V'���kf�h��}��3Ϯ�IC��6
柺Y,؛���er7�P�C�Yy�e�^�߷�A�V�����?���ӎY��r��-�i�;.���KM�A.�+qe�w����/C5|T���s��x�=��aNu����|&Wb��a���h�yt5S���scW�@��Z<�T�w
��e]�K���=�ԙ�w�L������.sy^���$fVRtDV(u�L����V�Q3��w ��uDU��,s+�,Z.��h<�Y/3k�Ad���>�*��C�K�!���cdV�xR�u��p�~͸s�m#���GnU�,5u�{S���j��sTa��=G���م��	���c\n������%>�w0�Æ�:G{y#�<�m�Sm�u,<��뛊#ϻ��:8�<�{�X٣0h�(��2_oLb�'��(z6�O��;jm3��s̺:;���mQSҬX4�g<�i1��v��(�cG��[�/���B��%�k���|^�<{�BzPIg����2�|�t�t��fY�4r��k���~��/;�Ŷd	#M�9k��Ԡ<5x��,+�yϜ�E�x�-;3�����K��^�y7�Q��wZ�}�����.��ڸ���7϶�e��*o�b�����n��$)�g:O�������łVn=e�|
a�-:o�]MLu	x��&.|� ��3ޛ�۴�;��ld�66Ѓ�-���N웃N�گ�v������8=��EA�X)�o�q��y���^6!���/:�+����T=�3��eg�%Է�*E�Gr�4Aww���ѿ)�/H@z�\0�s�	�z��k�Ϛ���9*Z�|*��^�#˭�ُ޹,��;I�Ut*�蟖}�ڿ��e���l����粢ee��n�n�cmZ�2�i�k]��X*���we�P�B�u���e����)�Nu��y�4&ա/ܽ�9���#�n���L
S;�P�e�;S>��0�����f+�s�ӯ���q䵉�M�����z�v�7p����޶�-�g���I������N�j�-t��[��[���mE�9�n��s�|��V��^/V)ˢe`��e����=��I�u���I)���ֹ5UQ�Q����&O:����\�Uu���p�{o��Y�Qޏk�z�4��>�:�(l� G�o�E���B���҇9o��+��"�;�O#O�;���֍��"��L�e��s��'vL;��.��_/]Pz��CP���;[���Y5���S]q��sYs��Q�҄;b�a0�u�Ѹ��=q�j<��Ⱥ���1z���=�(�����~t6��>�G3U�����'M��P�]%1Н��998�M����ϓ7t��_Z!��͢Y�4��b���$���,U�bnQkR菑�5hK7Nj�5׮V?e�ؖ'�#�S��{r��\,�W��^r�O�;����4ћq��+��mP7��O���bw��+�L8|�X����q���T��c��C�vm��~�����BԼ�����q���?9����9�����U�E�������^��;$�^kDʇn]�^>��Q+�.�������O�}��9~gy]�V0�/����5ie�d�w�O�&ec��+�is�g�j\�虇��{!�r�g�6e��b.�ں+����YO<��6)�rߘ~O�s��R@��ʆ��W1w��=w��5Bh���u9��Y�a�ר�7�Ա�-�����$t(�NY���鯫�n�pC��B�er�Ƃp��Ƃ��҆t�:�6�ξ�4I��U�1�%�"�FgZ�p�-X���x��v���WA��	ƙּ"�N��b�4sh���M��4��ejExo�i���}���*4���2��	��Bu�I�1�*�y8����^t���1m:t�8|��Ҕ�b�4�ҙ�S/ǎ/|�7ӥ�~��}O�S�F���D�u����N̠D0���{(P�ԙ�R����m���y�ҹ�_��(u��>�g깽�p<א��g0)��,S|�Юn�ҭ���r�B��N���8�C}��#��l�8$v8�j�9o���y�|'���洙1�SY���������P�w����z����rƿE�4�1p�br�~�������� ��/"'է�K^Z):�t�������:ڕ�򇱫��6!�Jn�KT�]o��@b���%{DH� �=T��c�7л<%���}/��%�/;��/}oo�uY'؉�{�q&ÔO�	=x yK�ѧ�g=��̠��آ [��;��,���*g�����Z�m��L�
�
,�f���pqmi7ۊ����w/{�F��*�h���s�{a����;�e�K���1_m��g|���Z/Oǳҹ����?%�b~v��]�tr޼�8:z�B�L���ι����&,}������ �az��H���,�M[�{�{������Ҽ��Dt�*K=��&��o���(����U�_)����z�U��n���/�{��{C�@�[���+�w��0��z�X���
�uj��3�mC���=�_���}^#}vw�4�{ۙ7�:��Ԟ�%��~�q����:[���f���:d]�r���4L�Օ��h�.����Ӆ�qpx-���K�0k����Pm2+��i�ȓ�߫��ǯз���'sr�}.s��!��~�#r�』Rv)Pٟ]�x��Q+�b�2V�w9���{C����M������������zx]���ڶ$���F�R�AUP����g���o�jM�Y�$��=�q��U�e_Rѳ9���B� ��
gN*��m���~Ż��q�H��;��|�.�eCd�rg_x��~
���Y��;�n�ԣ�������j]�{k�¡�Y��_'��갓=�W�p�>�Z'��Z�<β�m��zz���$1 m�A�r;��3<���qW=D��c�7A+��=ׇ��A�O��+X<�C)l���Z��
%����Z��K"��'�K�b��*b! ��j=It�K	;۸B.�>�uɴ �կKwv�b�Q�:��Y�9��"�.k�=]�7̎$���R��QP��l?�^)U�3��x��^�������;k���B-X��%�CGz+ig�)�����թ2�U_+G���OG��ؽ�I�Õ\^>�`��p&a�.ȇ u�ر�+z�)F��g}�p�Ӹ`M��m��Mw�ս�h��ܭ5]���5f�O��K'b�F|R�&�ޤY��A��m��k�s�V��{q�y�z��6r�y�IW��,+�Ȱ��:a:geݚ�o�$d��)z��uu���4/}a�O�Zߋ�W�U��~�����{�}|�����ؗ����{wc�]mncX\�.��^����/�U�<��pmx��;�=�될w}Ϗy��gkU�\��n��O��h<��ݛ}i�|
a�-:���iC�e��������D�S�{K�9�,�e��B�����1�d���U,�����+hvR�]B�yu]vDƘg��o�樘�+��R�(yJ\�~Z��=�OJ��jV��\��7�f*�߆�a��m��agZ�<���7�@��ocV�v#�Z㾝$���Z�a�r��9���8dʑ<�� �wt8.����TO/娩��3�zX��v�n��"{���l���A�i�Zǹ��e	^�T\��m��u�$�3c�a]6��u<�g�e��0C~Z����[0����'-���q����v*��b���ޕ�6FJ�qn&ߠ��V��>��˪!�T⬎��g�jߧe�..k`\|j?V+���a���{vq+�q�qq�q����L�Y�U3)���v Z镠�]{����u�����m`�џZ5���D;s(��LR��)�����D�T��a˭o���q���^#Z���r{O�Ӵ�Xsh G��7�`�-�̱�҆�uPȃ���[ҧ���%����W���.2�|�'�	+��xA� R���=���v��q|�*v�����r�U&5֝9�U3���M] �<2P�n�a0�P�x�V�f{O&� ��޿Doì_]KP���� �E���V��G3Uߜ��Y:l�P�(�`��&�]��'d|$K� S�ٞk��I���_��I-�(St -�-jM�����z�u�x�2{2��^Sܩ�Q}y�r���g=긽��s	P|o?
+�.���Y�8em�ʙ�ո�gA%Vhf!N����A�ut�6�֋�oAxk����.fN�__��sz+k@og��=������ �s�71�srR�������N���7i<T�0@�b:��c#ѴȤ��|j^�K�_�M�n���b����!#Bo6�`�U�+�nT�4`�b���#�uqF���j:����\�=��-ճ��{h��L�0�pUW��"B�j'jq�� 4,q��`��6c����zZ�,39��O!y��V����\S� *N���j���^�.vO#������͇��j�s�I+��!�fd����t�ؔȸ��U��u��^�������M�]�ӣ��'Q�h�n_'�6Z7z�pG��_~Ax��9p_o���{8�.%�ڳ���x�J����C����u<�sw�S�< {Ը��Ub���wvi�m�z��[`l�X͍�M�}f�'U�9fKrVJ�>�&ד�T=��U���>�Tn��a�PHy<T�.�b�Ͷ��R�M�\Z�"4_a���k����S�j7�Ë��u&Aw����\�k��>���
oD,�,Ng��sZO��[DD^�M,��]��h'�^)���.�3�$�wJ�8�� ױݘTz�{_8��w�E�G!(��9է�os�٩�W�m+�}���s{a�9���r�;�ħXU�E�]]b.k�[��;t�,���#���7�"�/fm�U����(S׹<���[=�Q�P���b)�q0� tg,�;N�(��nE]��^��8�p$5B�;O/'ë��э{'��g�͇ۯd����ϲR�J��z)���K�!��xx�څ�v�yݒ���'H�@��Kx�"��50�츟��Sq^ە��t]�NܲvM��p�U*�Z�z�2��5�G�6ΐ4c�]es�ONv���gk$"A~�?Q)�`*��;oM�0���/�$�GW���=ׅaf�;f5���%ޮ��f��O��:�#��SDHJ~��![�i�7�
��J�*0��)B�-�.��GR��\��"f-�6W9V`+;�m�oyV��K�vWPڹ|실
��\��v�Q�R���۞�f뤷w����5�&3M����L6�iY5Yn!x4�[�N���[��ӳOGɂ�l��)�2ǉ��۹��ީ`���vFq%��k%0�Ӌ'sӷN��rq�.�S4�LJ�z�F�&ع	�:QO:�Ʋ�o�ۻF��jS��٣�]�+�T��s�
sra���OG��֒�۝��͝�:C�Y!_nC�
��*�i7��&��ٓI��ޕv��W�Ik�����}贌3n���
����v'Z��xs�J-�E8�Ac;5"���'��V�d[���ݱ���v9�;�RYYټP%�i��XU�	�9�=7[;�f�|l�6���7:�wk��_V�UH��TAT��AEJET@QEM45DQ4�Y�LIAHD�R����ML�UFa�Q�-4�4�-$KT�50PQQD�U5MM2IB�PP�1��PQM5E,TD�%-ULER�EERU4��E#I�K5�4AH̕UT4D�SI@�QECM�T5M9dMYQT��QCID�EU4$AKQ	EEJQQT��$BSD��T�%D�4ADT��$AL@R�T�P�I2��DBD�Q@SSS3D@M1U1AMMSL�&A�L�4�T��QQL�]Z�_��=מjΎ���Ӏg�]�����o�>bBQ�߷�x�������X9�^�x/��～�pO/l��o�&_h�H ��n®�7�CZ~�3�m��Əb>8)3�z�k~�Ֆ+�t��C�xۛwAW��5�yɈ�ޞ����i���lެ�Zޣh{kj�!�Ҵ&ÝX�`��lt_��O@~}�]?gî�/|z(�����w㺼�ユr�����t6���'{��L��x��Ҟ�B�E}_sU�s�g�R�^~���G��9ī�SEݺ����ڞ'�X��Z��p/��������.����w5xN4δ��B��+,��ź��;9�0j�V=�>G��˓Z=���_*�3�<9�9���=���u\{}{[��7� zjoW�l�֥���:L	>Z���J\x?�%�~|F��ٚI7>�&�vLN���hB}���W��)^�hl�l���I��s��L�|��z���hO{v���07mD�K���g�{�G~5�9�2��S�6��c:Z$�!�ڜ8\�Ì�w�3��|�����Ϣ�)�w���N}#��%��.���!�*�u��Hm��cN�� ��.�q�-ױy..����$��(�nԄoƺ����v�,s���=�����i��]Fh'6�!�4'���>�WVU�Q��u�[����m��/�+ŋw������p�]�~P�f�T|�S����6Vׄ�؟\Y.�4p�[�̨��)�;9��'��E�+FN
�r�m^�f�x;�5��`�"��p�br�HA~���!��oO]��I_���Ⱦ(԰?�!�o�,���o(�bb�[WpEs𗅼�
����H�����/I+�H���r��^Z1��
�~L���6<�Z`��S�p��[���i���q}2M��}&U���Z���O�*S>ڨpݠ�43:���C��}m�mnlz�y�l\t����I���,/RΖH���ೃ���<�|:�j�Q;���-�̘�{���Ы�g�^�ǐȷ�Ps��L�:�����R���3�u����7�7�(����x������o�'�gu:�Xվ��}��1+����o�lv/gf<G�t>��O�n&=�b�EO#��ыJ��\8�Dwզlyqw�[�������4�Sm�9I�f^�: �K�A��ƿ�4�~�H��B���J�ρc+��I�]���u��ۑ��{$��L��x6r�6��K��ȇ}�߼��^k�|F���l˶�%�Ľͤ'�q9[�����ڝ@^Ÿ-3GlB=���t=R�N0��X��;I�?D��4Z������F�lW�	���ks�\������V��<:��7PTn�͵�������>)�d�I�Xj���lշ���jȭ���®���;�Ekw�x���O[�8Á9�ϧ���*�xQ��M�`�I��	�f�C�-RJ��ku���^S�+zK���������P�`�i��K7��W$��U���}k���{�OV3\Y�!��u �T��ςO��ء��t]�iδ�)����՘ꮻ6Fgf	�s�����3\����B� Y��!��i3����f9�L�����3����L�0�me�֤�&۔9H��T�g�a�o�'�KH������+�7�{Wg�����ō��3-p8T"�S���e$/����3�����ԙ�@�W���7�M���n�Ot�b�]R��vUqx��b�����n]�����ȭ�F5���tpU����z:=a�/ϏjDL��U}�"��Y���=(�0%a�IZ~=G�V��t��Vz^{��[*��u>��3r[�C��g����dXY՝0�6'{#
��[ֻ��=c�ok��V'�8lu��V��������=�,+��YA|g {ؼ !K��=�ֽ�O�wkq���ޟ����}Q��Yq#��y��V��ǁ��)+�����!���)M�b��:�j�,�NvG�F0�E=�Ĭ�n�\���1�.w<B޶���7�%z�"n�f�*���ί¾�^�T�V���e�;��)�3�䶅�e骖||�N#�Y^>�R���7��ݺ\�[�W	���k�m�T��J����W5���N�WZ��y�����-:o�]MLu	�����.�G����<�R���k�-��U���|����tۿ}tSO�z`�f1���5`c���N>s���i�l委m��KP�0��]�z�}�s�pI�
����_�q�f��q�׆�ױ
�;ɥcD�[0�s�	�z�8���d;OT5R������������]\)�Չq�(*��]Q���.C�o/C�o�'�?VKwH2��}�z0���~.>�W,	ˣ�z�LͷvZC�맫�2��{�Hј����kܹ�v�>Wϫ<d�ϧR#�M̠lIQ&	��h�L��v�Uql']�Ku��}Z�gtk��S9ԈQ��'��g��z�p�f�,���&f�4����m{��{�)�ya��u�vJ�}�������+�L޻�&1=�.����m޵�2՘�����ns�;K"�a�p�(�.d4��x��hf[�Q���Պ��OS�.��fq���	�:�QR�TׯS� ����f!Zn��3mL%��(đ�VR��Wh�[ր�����4��0f	���˝3+q�L�*�3���TR�p��=M�K<��:puT>=��/H*��>ڙ�Á�+F�P�n2��^޹���해G�O�q�<o�pu�U���m���"�Wp��-pr��Kk7ܽ	�.:�d�:�/}O�=jW��O�HŎˮ2���>�n��ؒ^�+��b-���M�q�ڵ��}��^���D-{�#u�g�J#,ϗ/��U�/�����4����~�Rm"����~�j��2T�I[ҽ-W��vs�^Vw�����Y�Z�a�Yl�|�}�Y��/�׎�
DO����pzz�a}��p��*�4���]�a)<�#�aǍ����D�z��}��/��/�%�T#�n�wW���5ѭ�:���@����G�z���x�U�������Qg��5B��3�T����e������f�w�7|��r��7u����eh�d�(I��Ų�ˢ�Oh1Χ�< ��N�f_���$�:���N�a���[��&��
U�e�%�Tit�}��Ȼ��W���;�L��h�� ��xp����8�۸M$��O�yRFUǾO�4�y.���Ba���Y�����]\�9��Sd-*39���<���DY���u)��q�-wD�87�T�+(�3�yأ����-1�a�=L���wϺJp6U�cc=O^s�gS����
�&�{���x*b�	Ӥ���娮/n��TM)���{:�^�N��9�=���6}�Ǭd��G������	�t{'fP"�0l$�{
��6�Ќ��Y�:�*t�:��L�=�����\_Y��z0wd,7̀1��Z]�7v{�~Ɔ�ȅ�yƇ^u�X�Ϲ��Ǿ���_\��hɐ��/�u���_���q>��D�W�����_3��c+���foW���`ӂJ��o��Ξ�I|��A��0���_�p��}�t��V�:?I��Ki.�c\^8�����>g�N�Ẉ�����'}��tH�l	*jϪf`��RP���/-�|)T.�.ρ�Lֽ�ruQ�8��1Cy�m�Sࡸ���I��	=x'��א���O�*S>ڨr��w�-x]���t�/����"<�:Um�Q��	ό��.�H�&�����'5K�IO7�������{r��ab6ڮ#/�a����A��=��Q,�\uAP�鱲��+�sQ���м��{=��e���"nv{$��q2�]-�ρ�Q��`���id��қ�2&��Íf�{��)�1�k�Ӵ=��x*ط��-���t[M٬g��{���Qq6.�۸w7Z�d�~7��&ãs�Yi���F�2�n�u�lH��z���sT'�7UӋ����BU��ǨcV�f�چ%c#�{���y	B�ü>�ï4��Z/�2�ߏ�@�|V�{.j�:=Za&Ǘc��)�VvWG���sT���CK�V�iŶ�WC��{료�\��]A=^��H�������|����83�{tE�� ����M����c#C�5�O��X�U���cb�W�:r� ow�wz{���O��O/T2JY���g=���P��xQ��j�8d{j��́��`��|�V��B�
�T8����_��Cby�Y�i�����K77»ý�_��dù��7ش�G��S��)��C�����)��6T62s�8ξ"������z�i{�u_����v����]y��GP�X(&E|/�`!��$�O&�p��8q�������m���t�]^�2��,s���;r��1�E��g�B��@�kR��f{jS�F����[����w�s����X��s�I�Em,T�v�]��=Z�_�
�;�M�	8��[w�4�PZ+j���~u.�T�s�D��Lx�޺I��pS)�����]o;�OU�"���]��/�I\ς܈R����C���d�2
9j�7۽}�k�{w����K-Z���_d�N��!҃361lz:�[�i����!���g}���!��k����[Uqx����s��;r�ȇ�#b�ȭ��(�_��ӽ\�Y�%�i����{iX�ƪ�n8��F�
z��N�Ұم��	;�u+)�[��§��m��#����A��yn��Y�(/���[��v�tj^nC3W����݋�����R��
����L�6^����º��[@���]!9E�Z*����6�Wi�/�vQ͛u��5�W�2�j�q����8��l�f�&1z��u�d���� u^�N�^�=�Yb���-6���MLuKP���Z�;g���.�K垹�^��}��MC&ˏ��ӻ&�� ��Ӛ��1s��9qf���o�rj�q���/���11�̰)����<p8�j��z�}�s�pI��ǝi�"��;�U�/�:������C�-`bia��[0�����^�}��2�G�_��
/S.i�R��ٽ%�3�-.Ip�i
֗h,V���V[V�;,����x|��.�]�^�#t�e�	��*S"�o����k`V߻b��X��	R;/�͙<���+x��V牵�W�U��I<���{4'�Mx���H֧�+���AGx'�rl�%N�]�;w�u�h3(�
ݙ0����]7C�z��A2m7i��ۋ��::D��W�σ�ʈ�Tg��Iq���y�P�@��+He榖�!=+��������y�Um���oV<�u":��P7%D�8�3�&f��jg�\A�˓%�ޫ\^�קV�vh�%�{'!F��o�}�z�,�/�M��/��@������|ˉ�3�����x���;�����s���P��7�w)�uvL"b$@;%��w1�r:�{Z��1ߓGum˰�Xf�����l�:s����n���AVxd�ة�L,�����Ќ|��f�j3S#|�R��j3�]\�]>���kY]�¶qn�-h���y�ߠ��7\Xm�3-xLV�>�5P:2�h�%t�Y��|6RKvP��t�2c�ˏ81��x��R�(�.���%�8�w�u�{r�녜�\Z>/��W2G¾fq:wd*py�+��Ĭ��̺�j8_m�:ٳLm	e�_GGCPz������=��e��.W��0�D���I�秬n�|�i���7T�;��W�U�k֫�+%\ku卭/2I���9L.��+�������W� �N�y��2��ר�D��ڲz��~�<�A�V@[w�����M��r�9�z�TC�K9	�)�*�c�D;�։��K���`k6N�*{�
�[�RivuY��ͥu�3���4��������}��W�Ip�����Nmi'u�!���Ϥ�V[4�\.n�ܮ�+L�������>1}�WԵ�3�sW���{g�7����y[��*On�OcEY�ώ�_<����>����tw*����WAcx%��z�tɳ����L�P���a��Q�=�)rcgȭ��q{���u��[����5�u[z���}���Bs��MM��њԴ!���`��{E*���h�����8����a�����̷��6p����D�u����N̠D0�	/Vm�k�pX���zp��[=�;gD\�f.wX�>UO�b��yK�l�H�oqY=���<7����wo�&!��C�{8З�sV)�w���N	�2��-�ˆ�&���c�+�d�3|3�^H��U�mS#Ԭ��Ca���cS3z���`���y�%��7��"L���@;,NR��?	^V�/O�K�墓K�,m�㊟�����/݆u�� \�+P�b�_=X��sF(3:jLh��oc̠��
�xB�ܯ$�yY7�pKw��8)G]�s	۬�N��C|�{T�y[�;a���%9M8(�VT#�=���c��s^ݧ�Q���s�3>�x�p�񛔷�Od��}��)�U�y�h�:��g��u��<�cFL{���d�M�p��>���1j��wV�-|-3�Zʎ���Z摔�8Lw��-.WF�.[ϕ^��c��Y%�=J��(��f��'�?�Y�^6u's��U�V�/)�?Nͼ�=���B���J��� ���_.1��/�h>@�)u�����Y�+�\6-7���F��Tַ���;��4�},���Dmlm�q&�.5�U>�q�Ox߆֩�'�D&n�{FX{sM����+��1��h��@��GB rO�]&�Y����������}-��:9�7	��X�nubњiȅe�;�-�+�pJI+	��t�lCk�������ܱ���@�з�y��wݸ���yb�r�s�6��x��[��mX����m>r5�݈�5���'-gFF7Y�M�3�2��]7[#ng]*[%>��W}(\���k�HfR�X��[�4���N>�<A��7�"�+gJ�z�;��[xD,��b����sv�|�L� �}����n��+H���ޫe�&��w5��nK�r�/dӞ�p��p�#�F4���2�y�G�\�����O�Ř��"�h�A�pc�>x�A����Q=�|fi�7p�c:��G���I�Ju_�)ffC�x����\���� ��Dv��d���W���Ȅݍu�s99�j;�Y�v���pA%�ܭy��݁�u2q�1��n����¬��%�PS".��_�q��Y�����]#5���U>uov����VyvW��.�\�3p�)��ɽw2� ��{o[�e[dY��������Ã������{�[B+5�Y�xv�o���0{}����p�m�w�׌h���#$d%��bq&�N����W��58U�O����SL�"}�C�W�r��7���3�Ǖe�{��Fn�O���f��ֺ��%� Fh�^˙}�Ffh!<�4���w	v��gY5�ҩ����!��ܺ��)����#��2W]�PZ�5�b�=#�:k�Z�� �,�pt�H=�04l��X�_N�d��%�.�Y4)ZN���1f�ַ6�잔�	�l�C���s��]�F������L,7)�)�vz��c��B}v����ُ+��}�E(��u��>����>�OF�X�r��k�^�X�e�^��R.�$躂��j���+�{oN]֕�'7`߻��^DKEx�q�(e�>���^��	�i�lm,@pPc�p��ټ�8E4�sR���3�k��Y��Ɋ]���A�D��Q,L�UQEAEUTSU5�`5QE0TRLDTEET�T�MSPD�QEddE2QEUQ�T�PAD��UUSLDRESUT�UDST�UIMAETQQ4�P��D�51D��U4QTEfe1�dU���d��TDY��T��bQfaT�aX���$�Fa�Y�DT4SeDVe&fIPUREUd�dUDYdE0FV8SVFQ3IAD�CPRe�IIQD���51SCD�TRE9�U��KPEU55VfD5L�Ye��5DEDSQUVa�LYeEUS5QC�eM4�%4��T�PU-QTU4M0D0EEE��SQSD�S�Uda�S�e�SAEMMNFA@��� �3�a�V)r����V���ӥ���y�q����!\��
���CXG��7��hu��}�\�ep�I3Ƿ��.���7��ܮ�9�J$h7��5`���{�t�9� ���yhƗ
aC�Δ_OW'� |���{��|���"���\m�\	�tt�}	=x'��א�h��ʔ϶Qw�h��Y�m��y�{"����Gz�(��d�k���$I��,��pN�m�"sf��׽����D��T#/�b���0P�W��c��%����/
��
̩7<�	[A�I=���{��-�G�obV���	���t��u1�P�����Շ�0n�bZ�O.�����|���G��v�V�=tՃ<kQ[��3�ei[*\G>�i����ܝ��t�����[��;�r�ɼ�r�:d���̻ۛ5~B];4�=�l��:�`���H߈T��>@5�㺻�v�'9(=L���~��9�=:\�VD;���ظv��,S񔧻i�^�uGnn*{EG1y,��S�\2Ė8É��|'��åC��]�F6��/'�H��x�KԸ��u����0c̮UY��Ρ��a�}vzJ�l�?�K"R'�Wko!󙂐�z7Fi���(�Q�y[��1��yf7=�fd}�d��&|�g"1���uw�s��u"j�㜮�J�D�G��ݝ���B��l�C��#s�-k'���d���i�Xxw�\)�#m�ww��-c����Oa������.a���W{����w�x�^��+Q��g���.�9J�^	>S��*�'<��:�����2��8&�z��YgZ�g�u��%��Ղ�dP�4�6z�$�{k�t�����1ёfn�3ν!�kk�ms�g��g�xXy�����E��W���xl4#��ǕR�)R��e���ʽ��Zw���Z�pL�E�����RB��[K*S;x�=��jS��L����-���(N�VUU��'�A��������_#�3ؗvD8y�+z�oL�p4���߮f�|z�E���.��`{6���E���}r*05f`8)�9�K'b�Fi�s�庽�;���9k���V}J��g��	��Ȫ_�e�*;�~���}q[!|G<Etε��-%���m�}C�ՏO��!����/�u����=�,+��?V���d�����I>��c�݊���b;��U�g����\��q��3���/��[�׵lc�;>�#���P�OL�Z$�k�V�������� ��q=pw�kT��c6���5���g��l��6x`w��<��.͵O�;�9le��N���]\���Տ20��[87*+b��oQ��Yc	�or�m^��n�:��U�2�okYjmj��w+�=����mʳ;,�9E���<tҹ����]��ؚ�M�V����_{�T�P)��]�ϧ<�w��OasUb���*u@}�bͶeӹ��c�w5v�\/�.{�I��ot��W�Aco����V4�V��}Uֻ �C��PP��D�4�zن˝P�rޯ	�>PSA�it��,�׋���خp�lǢW�����/�|���M!Z����A_p���j4�Q5�q�?������{�g�A�W�9�QpN]��h��f[�/*�b�u�Ղe2����0L]ޑ��V`&�������u��yY:�bne"�0x)L�
̼�je�O��\f,
���OyNy�24�Yk]W%sB���=��'����m����%��-kO��GK�v����έJ�[�u�o*g;��x�Pߕ��-�ϝ�|g�"L��/W���=�a.���LV�}[��/X��Ե_�+N��������/ �<2P�Q'+";�ʋOem��N�tN%bd:��[f|���Hpܹ��U�W�X��>�ſPy���
�f�{rv�d��.�)	Ua�o
GHυ�	���Rp�5S��m����8�v�&/V�jy��]y������A'�_<s�q�ƥ<�tަr�lU�N�8�<�uv�������,��˂����O��OD���;�b�v�oO4�4�@:Y:l��� u뤠�H������2�7{vf���>ҥ�;zL=u��#��oAn��PcO�u���2:=��ˢw�fb�NE�Y��W��y;���z@k��ɏLg'��*� �~�R{~EF�ԢBz3�|}�?T�}�beT���_�d��_��K~N�����S7���2���<�D��xɆ=98+��LyV��i^�S��=�����I��oۼ��Wl���9��EE�:�o��V2���ƅ��lb�y�~�_��=�K�06鼱���n�
��dl��K{���'�hz^�}��;�s�_v��A���5o�k��m�X���Of��u;l�]����[.����Z�R�7�E���Wz��G��L���9��=ӎw �)e�ŀ_z���~��//
ZY���m��}�R�����oU��oc���;ˬM�)Ș�YH淇���E�-�B��ugǴ��L���h��r�������w�^u�6q�=���y�.�EIQ {��.*�ٻ�58¶��r.Z��;�ӫKUӝ-b7����M���Y�������#]�ӱR;��;��9�_W���s�p����.WV�'�3���bzM�s��z�Ys��E�W��]Od.�1�;7S���Nϥ���4WW��lm]����ӟJ��l��d\m>�X������<� ��W��ث�W+��~��D1Zr�,���u�so�++��/)��^��X9�ϭꦦ֯�Ե.Խ]�l�b�%�v����p?�m���Ʊc�쿓�R�w�+g�r�vu��߹�̼��9��*�E�Pk���3�L���Y8��¹u>ٝ�n���\�]�@�7v]9�����^���1���l�ڂ����^�/VApg�Y{��k<sV��Yմ����-�G����v��si?{���J�7�ռ���:�i���U�:��TG���4��z����Wr~�8Ni�v���3�9���z��3��7�_zJ��/<���_B'��j��z��W8jw�Otq�ŉ='M�|��것#�b3�lhP��se`6f��גgp����K�͎K��h��1�LD;�/�gQ�x��ס���z$�<��}�מm֘��D�e��{]�;�,O\���h8���<�o�IH�}[��z}�yyw5�6s������ڡ��z�1u��v�E���l���W�r��Nɜ���^}��V�њ�]�h<|_G5nN�Ӳ{+za�5�A^������n��3�\�M3ݟlz�T�7�������G�z�� � _"|M��}-}G���&��m[s�}�su�U��B���ܵ`��u;AϞ���hw�t�u�;.�x����pH�q鍮��Lx_���-{p}�&f�.��m��XC�_o�}}z��rnp�3�7Qn�h�Qog��gg�λ`v&�
������Ԫ�]�ը���m���f�ٰ�n}$���L�s�ȸ�S�[�;{�O�]�w|�
�5�}��w��;�2�{�b�X�6Ĭ��ywKq]l�3=�����	�����\U���U�l��w����Vu�Ѵl+�<5�E~k{b��J-��Yg1�MS������	=�q��}Y�'_ۖ��.�M�>�L����L?n��L�d}��h�|�sTG�w;�ރ�7���a�V�᣺�eLh��*do:��ru�H�sGr
��%=��f�W���H�=��˼�����~�����}�6�Dz˷��y,���Ox
��~�������Ae�_B�q�^<i,�[�f���i���g�fV�^��_��<���~ط�����g�r��RCG6�k��Q+�7&�udӬ߄�z������ɻ��y�ѳ�Uc��F��wޖ7�i���y8���^��,t���3��o��V��}�ɷ)?z}�/��﫚�q�[ ���?js��8���l_dŝ��Е$�f�"e_��kl%��@��p�sf�ʎt���e͔��^\Y��/z�$�t���ɡ�_������\_gG��u�_P�L=����9��G]N���ټ'u��Y~[��Z�/�z\qg���ә�ǺgAX�O��B�����9�;W\�BHX���d�[2�B����Ŝ�u�/h�l@r��
t����4�龈x���S�6XQ}���pܯs��`��k��te�1��Iʵb�|'>��ӆӽ�o`]��f@�\Jp)v:���N�{;
��T�wŗ�ˁo�_({VȪD���,��r�ط�μ��Üԭ�3���&�i�:�
n�/�i����c�u�}_!:�����ɛ��qslI/ח�ubxu���L�����Q��i/��)�����<��uOv�nH+Cֵ�����H�$�x%�k����)�I����>����0�+�آ {`��O�����	��v�pzK�ͣ;�xv�VOen��)x�Ҟ�T�K;������~Ш7 p?�=BL����������鬇����䋤��z~tY���W^?l�cӟF}6�����q�k�͒���:�����e��7>���9�{j\�}����1��������3�����kK֔�.���/yU����b��:ꗙ����N�6�'����r("=Ӈ`�={O����p���{����5o�3�3��C�ޤ����6٭�`G���!9�����]�rp��p�H�%�Y�Z�Y�h*��C@1:9'�����<=�U~Z�;x�� �АǪ�r������_t����d�a�M��M!��s��|ƹ8a&v��\.��a��A��t��w�|��5��c��b)y���k��sd623����u|�?z�z���C~���;���6~�=�p<9�����<�}�^�=��s�ZV�{'���l��<L�`�}�Z�i�=������"R3%^H>��=<�.���vy��z�q��s|�PH�W��O���%�䪖��!�z�C���;
vY}��y�����\�]C�Ƃ�C!�X���ЩR֟A�dU�<K��(_W������r����uΝ}�.N�YK3�[�:��b�vE��}�Ok!t6Z�]��۲����og9$�.��-��+{�%��.m�X#6�l���ޤ���G~�j�(Mi��瘮���M�`j���I6�R�g�b2��{-=�L�f{`�~�4\V�=ڇ���R�����}�����I�3�d߾;.�������K2R.f3g9I�ذ�i@c�+�sn�P}\�KQ���Je|G͟r>�;�u�Ǔ��e�ajr�萺=�k���O����s#�R����z��[�l������$����E�vz[�;��L� (�����1����k��<���VW�$Q����{JW3�M{X5�t��ǧ����_�ż�[�=�þ�{��^�z��~�9�c��S����=�p���qޙ��ϻ^�Ez�(7�c6��=�&�ٽ�_���=���W-��~���}�Y�L+2��p���o�y��v�ٽUc�g4�7���m��(�~���]墳��!�ԩy�yɹ6N�}2n�<��纷�W�'��)�C���&i鎌Ԅ�J���^���by���[�F~�]�������Y��#�>��א���!����t�逹�&��͏]I� ����|-����@��ݿO��/���q�<���a��#uJT�T]k6�;����@��ӳ�a�����{O�~�V�ѸnͲ�s��1���<��4'<�:ˌ�ek��k���D��W�W�PTA\AQ�D��* �� ����D��W��TA_�AQ�
�+�WTA_W������D��* ��AQ�
�+��TA_PTA_�1AY&SY�RTw��_�rY��=�ݰ?���a������� RBTHR*!H�@��*�%)*�B$��TU
�D��"��U*�dġJP�T
QD�*֔�J	�(�J�)AUJ�i�̉IM��PT�l�Ns�JP�����aD�$T�lJ��l�IDJQ(�
A
��U(�l�UDT��);���p  77t�)p$�m �,U*��Tʠ�Z�mPV��ڭ[h�X5R�Dͪ٩E6�dR!�v440��T(JZ4$��  v�
��V�j�i��X6��L���
5- *�љ

�+T��Q� �kVQ)�h� 
�IR	(����]� C@(�P�ή@�(�n�� �QE�� : �[���Rr�[Mj��BV�H�0�QH���
�j�&��ֳBJ)J�$�**� 1��՚k`K)��V�[%E[Z3T
P�me�����i���`m��,Z�U	�Җ�m��R(�CCTB�N � �J���U(�M�����P$-�Vm�j6)� ��
Д*օ	�$ ���"b��T�UQT�+p �P��R�� *��f�*mlf5� �� ��*���ETI�V� �T �,A�` V��F*���U�T
T�VP
�3R�*�*���\  \�QT30hi�X�рV���M�� f�D ZV)Z�f��
��QT��  ;��٦[m Ri�(-K�UM�4M,Р65	k 5� ����)(��@�  p
�h�-`3J*�m�+Kj�Qfh�J�[j�6��B�`Mk6¦-�V�      ��*JJQ�@b0� ��Oh�JR��4	���a�h1S�)�D���@#@h h hS�A*UOj�Md�фd4���ѓ �`A��2`�M$��@���h'����d� ڍ2xS�Ht,tX����,�j2"#l�	%)M�!�B�Y�u�x���/w8�1��̒HkZC�{�a�B��Y�d��j�	 `	$�5�I�cS BBI!�������?���Z��� *,d!Ą�$�aD��$��ChC �5C�
�p�BBIRw����5�>����?ϰ��C��'�&L���a�?7i2}w�~�Oʗ�xh>0�5�������aZ�U��Q^ہ����\ �v3a;�-�W�є��A /1�)6�B࣋T�,�����!*#zʱG(hą�V��͢�!�F-�e���sG�ZX�b��u2�^�B��k��"�Q�Sp
�x�i#7�Պ���e���Z,���p�_+�Cl	(;؉�av
i�0�޽R��+/qQzBm�2;�6&�r���6K��ޤYL��P{#��cGԡ(@��z�ŋYx�L��I)��y0�z�V���ٗ�6IU��EQ(Yu�N][xp
Չ/m-��r�,���VmZ-g� ��&��`�8#.� 
�B@�M�j�^�Q�e��ܼ���ͼ}Ù��$M2Į�6�5#X�WM�Z�Mg�Ԩ [�"�pfY��E0q�Y�v�8�V!f�Fmg�hܳO@R�q�H71P�u��1��IC�J�%�Ҵ�4��*ܒ�[�^��H�`��hy]��.��^��l7�09�gfFH��u/kn�<��ӷNd���fՇ�h�i�)!N�nV�ҡSs/e%0�)�Jl��3��F�J�47 �n��Q�t,+sY��*v�<�ȅ6�{�n��i�a
�3TKבP����n�����b����_��B��u�H3�+��	|U����ⳁn#��]3M
L9�fɤ���7���W�[�.��z�判��\�"�,�J�G吣L^e�aVV*t��I�!��U0�GlP��-[�F㵤�u��U����*PZ�;ڇ�l;���At[����8���B1�!4f��2J����G-e-x�;y-��7�l�ɹ&�eYq9���X�fYV����B��D\,�"�����i҂V�K�&@˴.�"�sQ��W��X�d��+.�X*(�Ɩ�+e:WfQ��?�R��(��"�5픳y�m�K0P�"��.���W�,X[Wooj0�p�m�a�� 5.���n� ���. �Z��a�~�25j�ttCa^	7b�����)�9D�-J��:�f�u�Q�[�X�F�i�Hcnε�����B��K!X\�M�Z�-^�*�m��[��ԓ_K��1��5f˖QA)���pfJq�h�Y�iU�D�S)��%
b^X��:K�p)Ջp�H�Ǎ�.Y�28/)慁��GۅPf
���4)a����څk�s'�[F�ն]�o�u�@eL�&:N��5t�&'[@,�#F,��V�8Qu����(��ͱ�s�#���Fj�V � ��[*<��;�^*�P`D�P:����`�ᥦ[����%���(a�*��T[��؜�ȭ3VX3~X�-��E�����9WOAn�fU�l�q���h!YAiV�܃�T/l��y��uzd4�7	����s�H�.��@�<���:����S-60|���>��X"�6�]ւN�i��?]/�t�y�m�%�z̩�KB��/](��E�EH�TwX�De�om�%\������� 1R�dx�҇�*��"]ZH��y�r��"�d�bXQ�WD�m����6��^::�5*�C55��7d�F���� d�:ʳ��*���iP�l�bz�u&��t�2`��*���ŏ��˥4���P(��ݺ��F���n��a�彽t\Slf�؁�
���VLClb6!�.�$����(���q5���:��,��ͣn9�mޕEkܸ쩑(A�DV��kįT��r�����Ы�F��F`�]1P��P�V�Q$υ&��'p��wr�P�LȲ���sp��I�ճ+.�J��U(�+kdOL����f�V֙���#4������p�(��U��.���%)b��!L�F�/k5� 3M�ڃ]�ج*R�CKC �UW���n�L[Z����=�VԈ2�2��2�:
]�պ3E��Y7����01�@�Ej{�����D��+aۼU�6)+~�)o[B�K�rX��
�$dʺ����aj����)752]M�N}&���5 �ճ��]�� �����K�d�d��o �߶"��:y��+���I.�s�Q����e<��pԎG�5��[���
��bη�@
�[�
��#.��3�b��fR��9��\;{tm�N����ۙJ��A̍�d"�'L\�V֌�Դ�`�Y�e�L�բ*L)�֮e��e���͌X
�Y�\�� �*ޔVR��qR#���slkW��-�EX2��wu�V\��)Ye� �T�!j�(
⩛��	�V�q0c��L6�ܣN�"��*�U�f�D/5m��Iw������ʏ)ƚI�����1���p9B�yA+��o�)h��P�rf뙖 ;@4��.zaF�孧���J�>:ˎ$��Ez�Q�V=˰�J�m&ƛ����fe8��"h�2R��V�(5�駋)L����X��S1ਃ�Y��*[��esT�XE%�n��(��ݒ���[B+��?+*Y�a!BZ)�[[eS"�)��CVޔ�^�(�H|P�1Z���b4�V�j��"�
�X���	Sê�X�	��]͎<�a�B��裂]��cU���%�i[Wv�������&,���Ɓ�]�3/�� �V��cw�-��{���z&�wũF����n�/�ʗ�If��X�%\�9�Ԍ��a��mSs�Ljxn�`IGW�']ö+�h��0%�^�_i����4L�1M�����}��!�3��a�|/^�Ŋ��,*x�z���yn`��M�G�Q��hK��j !�u�!�q�+i]�h�q���ccz
HS�w-z�[��6M���Ƈ�c�zo7QG��a�I�� ���FL9H�=to~���ڻ�+\ѧv�EH�$���VٴN�q� j���2��͘����zdyh&6ުp���i��Y�U��t���1�h���SS&&Ӳ���Pd���PGF06�dJ�B�Evd�0V��R6�=˒fD�(�0U�*��r��Ű��1��Ȅ��c5*l��\�V����8N�3A�R���M��KH��W�*I��������ޘ�6\4�d P���gw.㕁Ѣba%�k��j*C��#�`�J{��֋֖� b �n�E;Ȏ8�Z�PDV���c0�a���t@n�ͼ����*̙tS4�!��i����ˤԦ�AWr�3Xݹm��<B�t���6k^�Hkf�΅=��軖+�We�D�
�f,r�\��g6tп���Jk
�f3e�˸��Y�_ȣMbè]65;Ǩ1wP̒
Ũ})K�AhV��u�&VV�DRu%TZ��bYq]��FZhPUz�5�aZ0��\a����L�Q����A��K�$��h��[�$�n�r΢�GU͕h�ҧe�̤�E�*�B��8n���㔌�V�aZu�a�~�+ED�*;�$����%���3�F!�g��+XUe�e�ܸw$�q�a�lE.¥2�	�œ+Cc7�co�;�	d��3L] -������r�Հ�낍�S0ؚ�{����+i��;�vu���&ӒfT�[SZ�vR�K�5�2RO2��&��`���y����b��f�m,��7)��f��#�2.l`�Cwr5�T��&0�ɹY2|��/�X��M.���Z�j�� �b͸�]l*MwI�wv�e�̀	y�,Q]6��BՏ��/eAt�t�U��K2`XѶ���E����LST=��Q���5�9�OQ�mn3����C,��x�
����Z�v��n�! 1P7c#��^����WN�,Ll��Y���69��ݓt��Gda늳@�SD#q� Ը$9�J��h`ˀӗ4ؠ��2���,x!h������*Kc.��ܼ!0)�.�j�;)eG���1��Z]i`��j҂9/�mD�\���C�tc�h�;_`ux�[JȘ��]�gi��P�E-�7���va�����)B*hf��Lzkahk���
�h��F��V��Q{֛�����řsA��ޢ��@��Sm��e�����St,��%;�r��$���V����v0O������l��n�1�E�7 x�DR�Q�ϣ1!�sk����Sfe�B�c�n���,��^���R��&M�w#�^�J ��bәFl�<x��@���>X�B���������+7�B�l&s�n���{L���,0�+s~e�R�n��x�B� �}�-��"*=s��w����a��Crݬ:~�j�A\�����`�k+l^nkU�⌶�b�����1A��*���yh�D1f��4Kr��$Ls5�P��J������=4���ZiR0��,ť�!�C��й�1��	����S�M^��[�å1nj�޽VF%J�uJ�)��ŋԤ�,jj�9����F�u�@Q�m��q7$gJ��,�$j0"���`݁m��w�d�G*h3#jU�b�c�1\�S�l���ق�ڋv�׈�CY�-5Y���_N�[����_Z�
�4�d�h�V�U�Fq��5/!ץ�先)@�ݓ�'E�a��i@6���뛡0X�������1d*p7�M6�!{b��d:�3"Ҧ��w��̰vA�[j�&F��*�#cwm���5��w4-M�f�
�����[ ��U2��Tc/08�7sQ��N�e�'(�J�:�����t�;
�(�!�X�# �g]7L�n�G�ljr���hG�^��Db��h�j�s[��KU�6T*�ڇU�Ǻ��ܥ�TU�e�V�����D�QZ��1���F�RU�-�9����<���7���w��uJ�t-S�"��[�b�ʶ[���a�2+��!���AVڑ�)n�U�0iV����#��U�70hM�9��o#A���V)%fT�l^^Uf���,l�@Bm���.Jy�k%�C+k3�����$�UNn)�`��bה�㰶�j9���5�*�ڬ�N%��(]
ӄ8�=E��e/���-�Q�T�)J┍蘩����6k�)�7-k.���5[���S�,�-� X0=�W�{bQ`��)RuR�Y6��2�{�G�xV1yyn�r��Z E	Tͨc� ��.��1kk%�r;�0����إ� UcU)�թ�G�tcRk��MP��Z���V�S�*ɨ�2����ܬ�#�� @T�u�e3N¤d$C�0��1�ӓFc�k��+v.�V4�F�#m[�C�L
����(uGo&3aՕF
o{��?j~���3���Y��$fO����fo�'T��R������Cgg�>g�y�\�̘�d%��H�����^����}W��%���N����/��;yH �v)c����o�l�;бu� R������������+%M@���A]��c]���J���'@�o�Ly�@����gr�}Y'B_X�'d
WB�f%�S����r����i�[Ԏ��wCqh�9K#!�ۇ:�Ir7ҳMM{U���H��Ղ7S�!��s���en�o8l9N*j��|k�G;-9E,]��u4p�{�ĺڅ寜{�y��$ �j]T�6�V\=�O]�F({Gu!C9��&_;Ke�ԛ�n���/��N��tg�0�����,��$��>�ܕu�;%�{�F7���k��`7�H;nY��RVZ7h�܀��.���%��3iIט{M��\��J���<Ht˸lԸ�k��`�=�T�{�:c2Y>
�΀q��n����H٬	�:�ti] Z�K<f�|�ٶC���BIwlN*S�1�ƱP�$Z-k��9p�pt�RJ+n.0�sI;�v"
�Ʌ����m+�h��2��}o����e]fsn\Շ��}yv��%>�o�[��8��ZO3)�16����N��Lܾ+l��N�Po^�/��޻�]vÆ��.a�0��"n͋{s��
+��v�]]W�n�9�sr���Z�Fd�����a��̰j�-	XZ�ǻc�- Z������T�"����Z���F���q�-'��=�1T�F-�Vwz��qE�im���b��G�C���Q���W�n�.@��z�YYܕKs*4(,;�K9#�J�^,\[�9y��0`��=�j��^Q=%�/7F�7�[�O>�s2q�LN��sN�.�r�$T�G����b��t=��\A��~@�2�А�F6P���e�\J�ZUy��bV�.{���@��sA�L����֊����C�q���ΣxprK)��/r���2�����4`Dk�"�-�Nl��=�eU#�j���x��a����È��q�������װ�w�v��%p-;� <f]��d淒�D����\\Nv\ŷ��c����4;Xtaya�z�^<�0�9R�I9�#��(5u�
r��NүMZ��1��.�	���گ8k� �J� ��ޗ�7�k����o��UnK�h��c�BǶ��m��s7�+'/�[�]��({;��k��;(V�B�+�cS��:�Cw���:+��wVx��/M�UD�U�����r�v�L��M��4�B�k;.�um�qm�n�owu�jS�����=���>���l�|G6��,��U�ᬭ�L�QƦ1Q�ʧϮM�)`8��9켧���c�Et*�a��'�J���]�ٽ���/[�|���wr�&��jf���cN2E.�t[��Օ��V�S����xt�q(��s6��ܐ��B��7�K��@���a�ڴ��J���5�Y�@�ߊnG!a�e��e�����.Ie��W9�����I���4��N�ۈ@HY�:��Z����;��Q���ثCv`}]��ט'��F��v��Z��`k�^#���DAEJ��7+sk��b��tt�U�0�6�GY���C��RwG0+�o�r�s�ZͰN� ��̰�)h����Y�h�6U��Z���r[oT}!�5w3���R����E��d����TUia�"k�w\M�]��jԗ(J��,ц	}����Ν��qs�#v�����Xw���O`ac_\�8���l������v���V"Cxh��n��p��-I5r��R�%{@��ת�5�A���)5z�U��[�8x/
�O��j�&����O�k��t�)\�0�m`D�}7��|��d��#$u����*�{Y:\��j
�jT���,m�殔(皮w��A���Vk�Ո|��,�v^0����YR/�.(eY��yݲ[��Շ���n_2��yv�[j�АӁ�A��]n��T&���9��j�*bWA�V�)*�P;n�� �$5�3;�ӎ�=�EK�6�mF���x�S[�[v����N�(խXZα3VVb�V��yMK�ӧN:��2��gc�I�(�+&��
�����-��[����|�붰I(};�Fx� `�k����I�.O(ñ��uj��{�Z���rO����IҘ(�J��u��k7�+eN�Zx��0�7y_Z3z����(,SB�DAe��A�/1v�u�f]h�O9>�zPȔ�BPK���Տ�p�Zp����uΩ�v�z|9����1��.���WR�mv�/��S���]E$��'����,kv�oK��[�j���T!^���ٜ_c��٧Wk�o�|)k��=H�[ٚi���6i��.��si��v��.p:�´^�c"�Y�|{�
�YpS&��"�"�3�mG.ڸ��I*ܬ�Ś#�10�*<t�Խ�
�"�Z�p�^���1�N��+.mt�A���M�:`
�ܮ�Q�	�V='�Go�͒���Y��(m@��{^����B�ov}�6;w���^B��y�)1`�q�֚�s9ڨ:��	�-��x,�p��֚6��\o��{��`���w��%]���ܖ�V0�M��fNT9ڇ��/���BWQ�i���;�T�ה�Yt�k���uc�vڅ�����9�um����<�:U����W"�機g����W��G�R��z��b�_NGx�g��:%ulks,��r΂��5��dEց�b/F�6��6�K�y�с��(�\s&Yz�����-��\����� вlp�զ'��[���v��F�*�A���L9v˭���u��1nK�����sk��]�v��l�6�y��<�?nߖV�.��kgs�m9
���w�Û�]��Ck$1ZC��z��w>[N��Φ�T�|�2XQ�}�dJ1��&:Kx.���B�*c��@��\�ŉ��b�?���P��J����)lΰ�+ǚy���$�P��'�u����{���	�@�/��A�cfS��Ah����x3�va�\ut>��a����y��C��KA��l,�`�p*�e�L�Jr�F���V�#��A�Q����]����P���+��XO'aZj`��96�ٸ�#t���Ϩ[1�B�f�+��3�ݵv;,�Fa�Y�\�)
Ό���Fz��Ԯ�5)���u�ߤ��t���b �e^noj�=�:StWS{Fe�n�4�òkP"Z����K��fm��w�v�0��{X�q�N�J�B��d��鎺�.f�f���7N(���5 ����2(��
/�f�f29�a��ݑ�&XV����p�W�Ƕ䫤����s&�ه�����v�Ԕ3�qڜQ=V� �Hkد�oK��4;Ҷx���屘T��XY8�
NY�\i���G�d¤��݁�[.��V����s��][�	��,�]g\7�:M�:�G��]]�ap,�hAN� %7�˽(�#�:�(�t��E=�*�eE�f��j�lb���8
��ldT�Imը�WFL�JR�ĳ����J!�f��� �в�w1!�8����Aܹ��"�wZ�)sM{�eĺ�t�:��u�1|��ۆanv8��VaB����MD����6�����(kW�1A'5't�ܧSR���\HT�]�p����(��.u8F��5xӭ�4E��QUd�%�F�]�	����]���n�]]�N�&3+hlw�<w��힚Sƃ�;��`;�e����[�-N�yf�[A�M�gz�Y
�
;9�i�
�v�!�m#[��;�]�!M˨����Ԋ]su���ެy ��p�:M���2�Q���*�0n��fJ�f�P�u��� ��>Ӏ=�;���W�*�� �x뤻[�6���@���|a��t��M��k:�=+i�YO^�P��-�PL4���b����NR.֮b��c+K2(����.���i.�B6�˾�	{�ܳ��N����ԨX��)a�q=#���r�0i�0���O*r��|͕��Be�V��<& ��^�ԩ�|Mŕ��[�)�p��^������HL�,>X�r1{p��>���J���c�mZ�B�_�v��n�W�K��ұZ�ݡw��SޢMJ��E)ܸ8�凪�[D�Jb�UغНv.�*Vnӳ F�\�䭉�N^���:��S�vO'�8��Ҿvu�]J<���>���.��i�.����b����˺o�s\�CyT�!@9v�O�@��q�k$:V]�}���GK��; �G1�2��*�(Kj*��4����-�7n�mN�
��neEf�����͗��S�f4�E�3�'�BX�-����b�U���L�!����a�x��V�h��S#O1�Y�Y��77D��:�,�ݚ[B��#�8�����g�W&S=��H���+��k��@�Q��w�:���lpU,�y��b�&!�c�X�Q� ]��la��ݖ�[��֋ N�K���>�C���E�E��7	 ���"�q�G�̮:'�����;6�R�3(�\i��q%dޛ)W!�������&�w��ӵ)Z%v
!�[���Ƒ3ym�M��v�/��:����0�M�w�vX�s�R��c8�c�ҥ��z���99��x�E\T����s���Ƿ�W9X�^�Y���a���﫛g�7���^f`�"�tM��X�v�,�M�
�R�R��v�:����y$H��9��ql��L�ѐ��A@�\z�6��H�N��b(��:S�>#LJb��6 �d���(�k8q��%�sO*t��^���-�S�n>���+�� M+ٺ�`�
��`u�A����6�O��}�	]O�ݷ���ዩ�̌�N@{�l�1%n��E�b�C�to�^GP
��/��M���!�N]Z�rZ����f�s3q�U�ݳ���{[5�u�����R��s*y�ij���Sz��g5��T��QX(}�Vm��܏5n�*�[`q�%���ie���B����:\��`�)�t~�^���tm��SW�&���윞�L̾�iV�|q���L��&�Oz:�,�u*<��[dg[����Ѫ��)$�QdFLeFs&A��<�6��cs�V����2��0=#�oK�'Y��]�9�=�Vq*튌8�B�˪[��+�����՗��[��ˌ��S�Y.ú-��v�+ h�q`�J9:Ty���o{q/{��&o9�wr]�pÝ��^�3P�����r��YLW,J��9{��\��@V/(�O̛`�-P��Gs",�Ժ(��B��KMKc�vn>\��u_T��q>�m��I$�I$�I$���Im���I$�I$�I/������f�'����W�=?���$���8�;��I$�ǟ2H�@�ͫY�Hh�HI!������׿f�?>��g{I���V�nGubή5���`�1���z\����z-�M=��t�h�Fd*���Z)}C'#	f���ކw��Q�n�N��%```0�R��H*�)�n,��׫z#`�G��+�v8tI��W\�e��u��L��=Vz�gpŠ�Ln�za��uM+�ހ�����Xxb�ݾ��@P�R��e^�@�l�T��[Ǜ���cz��n����;�&���<�٫�mf3�n;�l�ƍrS��!j�cy�W�
�2˦��5�H7c-��b.eD��3m�D류����=Ԧ�P�&�t�,�ٮ�Åbl��;�˸i}�u�{R�3���!�8r�yZ)I�j�u(l/��vj�E��e�<�8�f��CF�i���%�w�-�u����V����BW
r0�}u�Sw	�m�@���=�:�#�Z㝊h)P�$��#8W'o����bW׻�k V��v�khnoCs�۶���͡�X:�W6m%+r�rr�����Ԗ�76�QlV� �I�K�'I��t���SV�UwW��.��a�qd���Vw�jq�eR�t���pJ�v�3�Y�&>rS%JI:�]��*�U��΁<��3s����4�9�'a�֫+e��H�[ܤ{F괝��Mfs2��Q��n$ͤXvY�zv����<)h6�G�q��K���R�P�r<4�b����f[ͻ]������һ0����Ó'WB�f&�+�������y;��&��5*�]|��q�ջ�8�ٝzR�ε�ȍf�۬��3w�����2��w��x�z��G��/��H!�:�/��� ����ڶ��Ś\�l�k�ew*X9�l������쾭�>���TvX-�*�Y]ݔqu؉�r�>��V:�]nc�HvJ��=��ˬL�6�&�*�zX�ltɗƣ�DF����A�t�,A�I���}�*��5s���$b���i�Z�-�Q�gk.�D���W����Y���B^]B��l�7�+0v��@�(�#�8����Z����[��5�."v�Dkϻ�S�A���}R��D�So�K�:�\)��i�·۴���w_V�nP�7�i�0�J���=�ff�� mеy��&�LJ�е:����cb�3�m��b���X�HGq�rB�0sQ8�(�)��Q��Ћ噜�D�fL;(Q��f�' ��子��;G=,y�u���ѕY[wF����ͬ��-S\W��B��N��r(mv�s��e���Hj�]8�7g���ma�hm�E�R�FR�]`�riUծ��k�J�!0�V�{yFQΉ�LJOEƷ4�F���]��ƋY�9�H�y��ɩ��Ü�\3�����Jլn�:��(з�ak����V����)��������Jܰ�jq.�tu�U�Wn��{�'
"i��k��d�}��I�KR-+.��=��C=�S�E���KW���U�֝Y%Y� �e�	�s;�U��w4(J[�#t��s��B)�i�$��g��w5�7T�>}s"JKkt�ҭ�eeb����AM7���A����'�+s^n���V	� ;Jq����\�����p��J���.��s���^X� �=�D�(ۅD��9CgW#�˸�;�r>�x��y�j��g�]I�&���ume4�\��=���]��ɱ�](T�����
U��H�]Л�>��I}��}�T$g���;�u�i,�79G{��aYJ��o�ĸf��uM�g;Q�a��l���T厓s;���e`�bt��:̵F�� ��v"��j .��t)}`_q�q8�җA�2q��0^>Hu���De�n�֋1��*YD]&�y�� �-I�G�cFd޹�L���`����vy#ө�5k�i�"A�,5,���
���զ9�׫Bm3���w�\s�D��Yǋ9��ee&��9-K|�*F�3�WA[��w$c�cn�y8��.�5C*:�gv�o�)
=�xn�4P `��r�4."�.�rER�Ĕ��}�P�))�n��
����F�vc���ɣ���vf��A

��gu`r�2�\P.{�כ�����T�m$6��FH�Y�V��jɛƍ3���qE�y�F1���h�nq�;w�G����ƀD��Fi��4Q|Ry�ґ#7t0��ٝ�cV\���0���fi3˝��\4�u���+��T�7�Wob�L�+z����v�܁�K�N9|�� �{qGf�j&�@eͫ'�E��<��Y�a���/��*[�BfI\�Ѥ���A`���U��j�]eݰ:��=��AT�vٗ�9�	�`V��bz(�\h͎͓�ݫ����2��GV�2�iks&M��V�͚:�$u4)�;x�/�=r�ੋw�核3�.�sU�Y��q9U�����SJq3b���w6Cޢ/a�&���o^L��Z.��ה,�S�db� ���Ƃ����D !�1Gv.�M�4�w���˅�S��qd(S�\���(��օ@fSi�B:���"�zeГy��������A
�t�^�fp�����,��rc�!+���-�1�Xs ��A�݅z�ħC� _h`�u�+�Y&-Qv^6&��r�Z�qm�'7��p�[4��h�����V�Q@��{���w�N}G�L�p*!�+�\���o�h�#�k��UrH%/(��w]e�M�&�owx�����ʻ�DBD��ywH����0r�Q<�h�Sl�5�b��7�>Ŕ]E�&"ȫ�'RN[�;O�Y�Լ�z��F�n`��.�й�*S�Rp��w�h�a��Kqv�{*"���8�K�S� &��t��a��R��!7PT���FLB����R�U�Ǩ�+6��Z��m���5k�I�Qͬv�cD�a�n���5B.+{8A0��v�nQ����qQѣ+�9�6A�W>�+KE�̧C�+��)
�F
�����&��?���3�E{޸5h�<z��7[x!���Xw�;xtx��[۽����ь$���z���w9��G0��X�5ٕ�]]fW�m�(��6���vB�H��>Tˬ���[�rݬ�J	2r=�H��b�b	�+x��dR�0���j[O�p��.�fq�馠GE�r��Oi�̮+"�@w|���[Jɲ�ōm8&�1�3;C��c�� �1.r�QB�jÀ�a�-�"���s���%�;�Z���)���+XV7F� 넏�t��v�:\�ܘ1�V�F5j'8w|��"�� s�Z���̕��V�n��i�"ЮNMic᣺���0K�9�c,��\����=��&�x�gk��pU��B�1���
����T�Suy����<�<�����QDg3�҅g,m�+�0�Wg0pTNF�v���%��Mmpu�����J%���v�*�Ar�yL:� ΐ{����ј��[�����2��hx����#W�,�4�˽�������
�CDe�Y; ����EnVlO�V�����vm���!��mr�l�R�~�ܕ����4���2#ÔZT;���p��1�+"����U�W���8j����frӴ�:�r�*a����y�\x���*?���ɸ�K^G�P�FX�{���2��okobމ��X����c4�ʽ�'E�Ù�Ɯ�,:8n�d���m��#U�25ɶ����I�PW���\�CS�V�wbJ^�"��U��uŗ�FF�iL4��mb����^Ӿ��Q��F�i惷¯C��@tB!�iX*��ٸ���Q7�.�c=g�gv��>�ai"�S^�g�+��F"�Z�H��b�*�-���R����t�d-3�Z�i���	)ώQ�\���`����s6,坍W-On��ꋵ��^�(��쭜ʹ��i���d��	�^�!�Ս
>��9��e�h+����Ë#-J�-�u�Z�['R�di�U�[E�"��ev�������.�|�*5⫤V���hqk���׳�T(�:^qw�
W�̩�jA_K��Re��˫"��GFoY��M]ګ��B�V3!�eIMLjhf:%��g �a���4�Z�o��?�1oQ2��_	m�#����z�f��k��6���}B�)���M�\YI���{�K�l�:�͕��&��uv3��ʳJ�-l�o'�Vt��g�q5���u��w�f����<�G���Ӄ���|�v<��B�@q�9�;�s��5\��/�d��C�TX1@ȏT��@t{�p2VVue��llU���5��i�9�JG:�x�%�h 6�U�t|I���P"��)Ɲ9t$7�5[��9n�}��&AԮ��2>�N)YC�꽳O,�u�&��z2�c�$�yX+�������1tF�^BU)��*��u�Du���'7�A�`� �؀�OK(�����a���v^��^t+9@`�u�a��fӜ2�� +�ۑN[V3&V���G��+�n�b�mR��R�{te��j���Äp���-�E��:�,N�����w�1*=���j��2���r��g��Y쮩�ءOU���U��%e�@b'�����]8����� �.�\G,Ҝ(e��-�1Ι;w�u-�jr���к�LAtps���]._N/��er�ޣ��Z�B*���.�O-.�e�����%7��m��u(�4+@!��I�?=�\�Z[Z�J����g'�I]��8^G����]k,�|c�ݔ�.LR���u>T�%wm	Lm�9��]��,�+Q� ��F�P@��kz�)é��$QWl���2F̷a��Q��Cz �\]N��&Z�a����/���9�ï*p�֖���_nf;���L7j��6(f�`��AP#��u��ڹO�+UgAyu���N��@����,o��-�i�C�W@m��Wk"=���
*�M�q�ܺ:�r�p�l';9���p��y+X/���5ܩ��/W�*v�,k3�:��7��C�Zϭ1*Q �������r�<@j��nV+�&IV�D4�㒧D��	|�Jf��x2��t�p��42�
�S�"������vlek�%��W:���L�c�y!,�Kz���up�N�82Jb
7[`���R,jtǼ�7ś)�f�v6��.z۬.�<+]�%ۜx�꾝�v7aom�1�T�]�TT��*Vj�e(�R��t�����Ԅe�"j�n��Ɵ�w�5��lM�E�3x�(eLG�O"�чE4��'�b�����7.���9���a3�O���$�A"2�R0yY��G�@��2"�ߨ��9��,�8�c���p�Yw}�N���G$�e���5һ5�y�PE����w��U��6�(�$�J�����M9tע����̱cBK�ݘx<ϻ:�Z�魾��s����.2]�x>I
pu�D�ryhՎ5P�WX{p���C�D��ñA֭��&���7�e�Ę�(��K�Ϛ�P�b�(���8��Ok��5�*�9�:�5aN��jc��9�� Z��K�ڃcБ����kJUd:\NlZ���Vn��ЕCN]�s낷����S闍ҍws=0�U��6q�f��ݪ��Sq��l�L�X�w������\�Ŭ�G9��+����F�t8���յ�
���A�-����u�U��Y$+�/���G)3YMu.,>�S5�}��Γ���F���(ݭ�/���7�s�W>]�td��k�q�������5�2�K��ݬ)��b�ahuy����]�jM��&򥷍��S:ѝ����p���Y�c��/0P�fX���q�XuԷ�2�9ǖ��If��� `(����*�b�1��+Db�������X�"2�D��TQb*�P�,QPEGZъDX�C��%E�֫DX��r2�V*�V�I�������2�`�F%�eJ�*�*��)FE�P��"���(��a�J���dG�V�X���AC�L&�m ������Ȏ0�SX��`�����
e� ���D����UD
�G3 T1Dk`�
����r�hbb���[*T31QEt�cQAH�!EX �V�mf4�d����'���TM["�-WEQTc�����H"�h
(�ĬY1&Z��JV��"����*�+)��.Y�iLh�X6��
�TQ��D���w��U�'�2\����^�m+���8��m��k��ն�8`�+;"����{�]2��~��:Ӂ����C���y���|fyN����q���<��3�l� �?����m*�nw=���C�!59����Ƹk?A��˅���7Åޙ��Iюӹ!ܸ
+͗3��8Dd��Y:d�b×
2�� ə7v�wPc�/��7�%y?�|>�\��S�>CM/�V�պFQzAڝ�>-�f 75r���x�!�KR.���Q]�%��)Bk3IO���P��r"J��P���!K{�	�� ሿ)SV��W}���[\�ulv�v}��u,�.&+(�Ҝ����D9z�s0�WdY���3����9��{K��`�?0�s��8W����U�C4��ƑNY��y:�\-�������_
g _O����no�$p�|,j���'u�{U���W�
=��euʹuvH�|�~���p!�'���O���R
��V��tUׄ��˳h�(]�Ǐ�.��C�)fuӛ�wʥ?!������>�Z�j�ל�����Ս_:�7Wκ��X�L�v3�K�t5�7s��|�8�-���NV�^wD��
����k�����`�}��[���bgV٭xϨ��q]�^ފN]x���r���_���9�������y���O\�u�G{7�BP���ɰ�QW>ؤ���U!Y5�P[�Z���ҏ��/\]��vhz���T��E	O�h�:2��V�/�h\pWK��~�X
�y}�찪��"�":f�aP��7D��k�#�s�{q �U�qN��%]�c��q���`%�B� tA��D9�g�Em����$\�c����r�Z��Ԩ�g�t�Mʊ\iM�ˉ��X�l�@�駍���ɹξ��y
b8��\�2�w]PDi�>�Ksb��R���D8����=�ٗo�S^1�7t����*T�NE�t��R1Kw�����}�n^joG�8����e�7</h�.;���K��[�-���)�W��F�ڏy���=���Vs��z�m�L���G�1�2V�;��ӃmVZ\��MzE�N׳��(�m�����f�Q��[����2�_Q��M�Z�p��P+KWwN9z��� Ӽ~�U���U�����>g��\�B��L ak�♈�� 3�+�aֈ�lW�I�&j�
�H�QY�.r����s:9K�1��C�qq'��ô'b!�ҫ�ØlT�g=ǧ~���9��=�=��� ܇l�����5���B�����GL�����O�,�=W��
�(G
!��4E���4��C-���m��⊏>a4H��a���N5Rx�ƪb��.	U�Gi�Y�;�ޕrßd5��C�I�"�|��2�/������[ɑ�S/�N��n�8[ ��O@�4Y/���*ާ�H!Д�xs�S㞧�EW;6�w�(v}�8��#k�:2���9��k����K�G K��3���?>ǜ�Y���R�q*r􎡇��"�oO3�����u�@��f_�Q,�	�~����ǝ�w>����rp���Bhj�pV���ymǽ�y4	Ղ����봧n���yQ/w%q9+2���v=�Wp�i��Z�b�]|�Ql�sy>�mm�n�u6
�@q�'`p��zk�5��H�/ƴ/��4�'ǅݵ��W�t�vK��v�(!�8<�2$8�#��:ed�0����tܥ��D˶u��I�k�U�G���A��Z��K�UgEW�v�d2���z��TΡ��{��F{�6O9B,R@��"ʢhxޚ^<0}�pH��ꩵ��F\�⢨�Q. )�q:
�9>�3NH�+����^�l�Tlr�Ң�n=0��HX���5�Z�(�VЋV6��b���uW��O��n�77�a�}��Ҙ�H�DT|<�zY��#�@X��xcI�����|nC�4厐�C�r���U]rN�[A��X�q1�.g��U#�b[󬕋��{�D��}�/�9��/�'����T�D*G�2|�� ����$>G��gfUϥ�h�{V-���v��L�D����=t���uo`)c����e� v�Jġ=�b�=g%D��r��"�pu�r�a4B�s"]�����>�+���k�Eb��q�މ����U�O��q=�|�b�`n͹�RaP�>��ɍ��紻K�V�'�g�;�+�ojk�%�G"����:E�e�86(We�O�Ȉ?1���/��Dzt<���:�˥xW�X����&��3X���!U
��.<Dʇ��Gd��>*��Ő�k�Ep����G�o[���7�
EH����D�x�=��K��<��|涾���Ƶd%���V�_��Ks�=���J�Q��ttS�𮹣�pִ�w�"� �|�a?%Aװ�"�(n\��B��#*&��$9`%�R��<�c�۫��4�\5!Em��;T�\�#E��ҥD�}1����-�+�Z���+���D���j��+u�}!��PH�fC�
bn�={���*����>�&�G�|E�9o����xÆ!@iA��] R����0�ym��Lu��q��l�4� 3��m��b��#�d�{����ԓ����ָWרKλ�"�q�C��
<�n�<�f'{wn�W[흯���L��Ŏ�AͮR�0.��ʹ����}�C����g��>^�
��2�Ԩߦ�~M��Kz�꼎��##�uW��!N=��|b��:s��vW�}����z�#���n�&��F��%J���3B6<J�@�
���Z���Ng�5�$���G�6�1�\u�rHQ*T	\jfԅ#`*!�� xxtU���͍���#���c5�P�0u�^����V�AV�\u���{�����g7J5�3�[4=~����!�M�����o~�}�-K�&�k��J�aHz�VD�78���-��!)9 ��0�:乜
:��s�����`%b �^��ɰe	D����5�ք+B�j���������~Д��GL�#�`���~X/�~˽�G�qbs�/�o�]���˞���r��[$'h ��~ڲ)nR��Nu�P#�[��n��Ѕ޲����X�[P�xu,Q�J��nk��+��[p�W{��Ʀ,&�W�u����ȵ���,���EU���;���N�[IH�`�*�&zB~Ru����ǝ+M�����uר�� ��j>͛��QAq�6�
po����+�V
pd[����t=o>Vw
��mO����!j�I��ރ
Dk}	��9�sq��e��A���\
�NE�[#,Enu���s��bU������D���|���g�ʊ�6˯���V
�Z��^p����C��5.!MϢ��5=��zA����=<���\e/qǹپ���`" D�4��34"��^#�숃�"��w���u�گ�U�􍉅��=N��W����h$gb!��u�0�S�2���W�R�_)幈y�̜)�L1��H�NLR�D���ʘC;��Q��;�z8�]F�9��qW��e�
!�#zJ���T7^ț�v�8sw�u\z����Y�f��##E�W��9	H����ˬ[;�,��Z5�3 ��4����!ǹx�o�YD��=2��� ݋�n/E�M���e���|�{�ա�V�+���#c�I����".��qW6�SuEb0�bDnҭ�P��ߘ%Nǜ�J��I�"�}t�!�a����a�W�L���^�g�aFE�=!�y*��Kf�-��%+îW�h��<�9�4m��N���W4��	�>u�!�[_
��o�;�>���uۏMX)(��"�+��O��M/��4�^/銹խ�l<:9 X;�N���H�8V5����f6q�Q��Ĺp:*����Dw(���7.L���Sh ����mx�2:�谩У+%Ŋ���O��E���v��_K�1Ñ�{�[�E�i}cEW�:��!�xq,9��V�w]	��:�:*�#i�htE�	�NqS*&de�y��ɬ��W��U�#<��PU�-;^��Z��<m��uz�ӾB,��G?3f�TS��L7C�4�!Ì�P}-(�A�}K8�c��uSp���q���2�IK`�
;+�,����w�O��|�����6צ�s ���/.|2Ȗ"�O����@�Ѯwu�Ƨ�;�;v)�
��.`'b�tY��:!f�z�T��N���W��5���Mu&�77�a
��b�9|@�w�@���U��^Oy�"��=���t�庰�{��f�.���i���cKI�be^���H3�D;��;"⸐ꊋ��t6���ɨn\ꮠ�<;f+���醖��H3;��H��H�to�����$Cӏ���ro�n�����*����*FE>\�`�nM9�
�mQȣ\�9[�������@u���u�
�ƈ%�ނ��}�cO˰P�/�Z{���,�R~C��n��K���*��F����e�����wS����r6������P���T+$��zUs��B��mD�[��Y�����$Nٜ�3���E|�Y%�}!����
7U��g7��S��3��/�lp[�)���WK�zN�S���;s�ي9+#����Koi�6���V��=eu��d�"��d.�u q9֝Ч�oJ��"�0�D���Z١�ܯ\��ε���]ϝ��YQ*mF��Pi.YôVb���+f��X���W���zb~\k�7FR.:�l��~��&6A��FA��%�+)�ɼ��=�Gav/��|2y?s���
*&�x#"�O&W;�䮍s�c�؈�r����܋�"�EÿQ�gF]=�NU��0�5�0��H��Ǩpg����N��#1��7ҭSr�6;���ڠ>�˥"����#b >�K�9�(�f�cJ��0��c�HJ�T��@'�-P�J�ц���(t�E�n7�aLB�D�e�JA����V6/����W7b7��]��x}�Puqh��Vi��p�ڙ2�W:;CEvj�ZԐD�m���I��5�ЧP�z��:��a��XkAت�znIb{T�w2A�r��]�^����Hؤ�V�O���?v��|��To`����������Wեn�e�u)�,u���м������`���E����WHN�b��,h�ϳ�fV�ڙ�oU�@�m����|0H���4^c�.E:�趮��C���J�Z�[]O*t]�_`�,��.i�48��wme©��|�n_\�,N0ZX#�f�yP-�.�f�h��0���;K��{���o�u�Α=Z-�^���5�
Wyٚ3S�}s.km�6޸B��ޗ�E#K9��Aݡsb�/�q�˩C�Cw�Q�]w>b+����f�sh1���s�CS�;t��;��%\xf4�r�2(�D�j�;�f1�|OGkp�a�MRB$���pa�ʝe��s���v��F��6�|�8�|y�<y>�Qm�t���Q֩��Zŋ �N��;��%�B�ΰ�R<+�3��C�G�]gqs7��ƀܫfKt*V�Ǹnn9J_g11��ht���b)l���'��쩤Ws��s�[��֮����#��/+��][ʢ�x:�<VU���\��:�vjk����mr�a��д�����96���J�Cn�诮�$�Ǫj��yu�J�c��A��-�F��Gx�P9�b���'&k'C�v^.G�5�T��hc���}�J�%Wl|#��yn��no>�)�W�^m=۩q�����¹��X٘�T� �>_��>�-O)-�R�,�}�z��J�dEO.+��u�O�QPHa�r��v��=��I]��i�N>ۭ��X��� k�ֵH�����߆����em�H)+�T���!���|y��+V�i���iඳ��pب��*=-���{E�,�S���͇��4���� ��v�X���ض�l��Et1A����kzh�eW���&��(�s���x]��3k����.�!�Md\�ν��*��� ��}�����M�b�c�����F:Tk:4 uŶ�ee]�;D��e�J��-V�󺳶���L*Ψڽ���P�Pޅ��9�,%�)H�Հ��m{��Lc'"K4��ք��p�Z9�%k{s6�h4������&�1��hr�V-j��7��72��)W��݇�r�QT.V镛n��LX�=���7�f���w6�q�\�ʾ���;�/eB���6�12������dR�)޵{<�VrK7���'0G�xD"*���I������R�� T��i-r���*����\h���+$X�ZZ�����YX��[j�PX��UU1 �H��b���C-r®TX�����6���PF�X�k%Q[i�QDS*��2Q�ʋ+.R孶ѥƱ��-�%�E�e�-�e��`���&%F1QE1*̶1�Ƞ��c1%DdbF�b�EQHķ0�*��e��Ÿ�.$�J�,QciTr�"c�*1DT-��LE���QXcQE�DVb��[-*�*�6�+�TbX�"�V�e���`�K2؃Ub�lb��<��m�:�v�z���{�x�^!�����9Ӧ$�{��eG>����ln���l�q9��Vv���� U����+��v �~��݈�;$`�ʇ�	���	N��{H��b3w�6�%����Ѣ���(����K,�C��V89���X��vM���;yg��T��RԄB��:[�C�3|
'�3p�Q��>��a!?	��r�c���u�6}��#*F�!���:v�jG@[�39�S��u���{u꒧�Î�ϰ�7�B2��\iM�ˉ��K��d��=���ȩ3�,�#���"��ą��j}A��؁0���η��6��[�[�J�_�����lq'���B��e����Ls��B:����w]�kר������R�DD��(��#�ϴ�J�\6��p��n��l;sw�W
E�â)J�R��0J'd���C�
<0��RίS��%��x��w��w�K�] p���q�fZ�q�^#�슙�<s��rf:�;N���e���m#v�N�����(�w��Kt�5el����JyZ")x'�wo=���������)��c[�M�;����sT���R�ٱ�f��52�Z�+`����q�벉�pܓ>� ��}��_T��������Zf*�
=�3=���s�ۥ\(خFap��
��B�+�#�Ѷ}�
�d��j�m�Fz@#������k��U­�_�P`(��
ƨn��������ݽ*�Ia렽���4H��0+�u�x�K�^�w�)�Iֵ��:qs~�~p���������W�@�M��1h�1�qJ\ob�&j뤷�K��kӱ�Jv�R:J��3B{O!]�fLX�2)ZWJ�sѭU�2���ʠ^}5���KX='"uA�����0.y��3lCr!���Y
�0�e��iazy��H�c�4���en��W#Ed��F)&T+��q}��/ƴ({MN+�]��{���y*�\,`)�" GA��93�r:$�^TGC��x��#�7��ذE����_5}{�,d�R��U�\�w|������-wǚQ"*i��!-�AH)~����yU]Us�6{�id�]��!�U�3��uW73�7�������wH9ӬB�\��(��SVK����ӝ?�LpH�#p<&2z�>���Q�C��4���ͷ�i޵�'#6X*:���י�NX��DЯ�'�"�3�Ό�����I���Z5v��L]S���T"\ R-��.$ue������J=�R:�z{��px�H�5Ң���9,F�p���CT�z1a܂ڌ}�Ca��B�3W9���J��j���0� �X����5���vk-I�10�TG���#�q���LV�Pȡi׎Hqp\��Gl���9
\EmGq00ݵ+�����-�j"����L������R>%[󬕋��ifVf��gv�q�S�p�:�����J~�o�`}���^�VD�<{��މܺg���ic�ʣ���q*�iySb�7f���U���^�����F��|kWPp��x~�8a�h�/�[�\@R�YժU�C�:�yHd>����:���*�)#h�E��G��Wo�Ec�g�oX�ڽ��\w�g��S�K e��wN�_�������ܘ��)�s�8�m��kY�0���x:w��\Lf
�  ��i�!�t\��5�vK���!�6(�+U���Zk"�%սU^�����
���pF�N�����υh}ʮ��ǯ����0fu�(%O.��`�Ң�A�g:��BD�������x����!Vr`<�o"����ݿ:�KS�"��C�R�� g`���7A �8*S5����{'o�/�=����
.2�(m)H��
7͗3��3Ä��3"�LQ	�%\���R�
b4���2FEu�)T�\�#m�*%�C��ނ�zeno ��T�3'gĈ����5�����KI��FS6���,��[T2�b2(<!P&��ҏP�Ϯ!�{�H��y�O�U�o=}�*#D0�7U(qäd*�"�TL�2܊وvwG��X�L���=��ey��\��e5~�hS�l<��-��W;� ���Y$�YG�z����У���q�'��ې��]4R4�M^�Y������P��V.�D�v��5����M�=����eem%��.7~���9s{����B�b��sr������SJ���u��;��f��w��%t�2nyDB�ʁ\���*d����J�AOq}�eL�։��g6n�o�	Jo$�@e��� �B*�53c
8G@������V�~�������,f�_SK�S�è?��z���h*�:瀚�F[��5�ҋ|�.D9둆r)�\! �F���5�q�Re�^����Ϧ3m|=Y���7b,N̤px?���*ܣ\���R'׬���i�� 1�hlt̯t�t�=T��E	D��s�C����rUBn�q���0�\�!=.t�"�Ȏ��6
�: ��"��EK����t�}�fV(~��,�a􌁱܎\�l%#���V�
�DU�p�������R?Zz郧��_�_^��#*(.4��q4�iGg0�#��l��s�Ol�@�s0&�i��IR&:�A6���Ks��ןӺc@�+>Κ�#E������r����	߲H����pj�;D�ڎΜKՍ*p/?�.���Y��_�e;[z?0�Ur*i_�4o���7מ�ݏ
�d��f��e�Ibj��]��;��{�����`���]J'�1`�t<<��|*��H�����.�
�:u%͚���8!��8B��!�J:<��@{*�Q�'*]F�/�%f�s̖̈HP��2�R����>�%s�!�B�E�*��rd$����r�u�_K�W� ���ϸ�����3^h�ltNH���.a��ӛ��=WY�f׺%H��nxl�B��!��Đ����٘.�����'\�[YܸC���9�ښ���-�ؘB��4��.LZ�F�1R���grYy��4��z��
�P*�W	=����
������20⤜�r��Z��ג�ҽ��-�ϲ�E�1�F¹�X�d�4��V�h���ۺn�Ԁ���S�g� �x]
hɿ-&;��Y��e]Yv�j��"�#�a�F�.F����[E�Ї��B�&��#����]q�`��"�g}u��2�u^��PT}�����.��5��3-gT������Ʒ}�*�����߹��i�Uƕ�%2����Zo��F�.I�mB.^QR�[���vit��O�ts�� W}�y9�27"Aَ��0�{>W� ���g�����}�ӥ��7���y�x	Oɞ�N�����諯���I��/$4Og{�9���a��� �H�$�W��(�zbTۑ�nWHUt��s;V�[o܅�X�9ښQ#�����|̎�H�N�Y.;�܍��[��ʰT�yW�xP�~���F�mg]%��Ώ���K]�-k6�/�#�]NB�}�C�	�zb!�+��bdC��)�A��-P���H��z�fW3�R�Y���*\J(P�Nnk��+�sJ�*}9!tҗ����4�!Ì�P}2bn'Ԏ^�&�c�ԫ��L����|���M��B���ib���ڽu���gz�,!����^�+t��Ԙ�r�E�|wpri��T H�G_B�.��Q�$g^���K�5�=j�[tX�r�H�{j/���R�֛e����-�Lޭ��9tR��J2�f�ApP�t�R�n�]1hom��;�������� �.33���ã�MψS�4��(�m"0TR���ߝ`~U4�������y�=pal�9Ȍ�]��/��\�}��`}>o�>��V�Ҥ�w�څ̡s��������E�R(�S%p>M�s��*���SРFz��~^���*�|��XkD�r2�~�ik��q?e���E�Q��c���LJ�<�I�?A�r�.Ń���{P(˭y�]݋�֕�VG@���R��py�|+B}ά7P��(�S����E���i�0���6�E%р/�zEH���r>����g������w9X�����fmK�OG�[�tk��M����3q'`eIy�#�b��<�ѻ��|���.*�wM1��z���o��":VS�;f[������T����Շ�}Ʊ��k'/����^@�_g��+�5�r1kM�g�1Տ�8�5�_f�z�)�|R���!+B���Z�a!���J���u\��`���u�]#�S�(�w#f_Z�[��)��x�>�-�v�J�FH���ξ�L� ��a��
v=7A1tйQJ�x�� "X��q��wΛ����b��Y�Q�!hÒ:D.=|��-�P=�ݼ�BƓo_+�" ���+p"<��FB�E�*&e�.[����6,�9��/cN� gH���!�͘sQ��'�_��\l�3��T�"	y���uW��L#Nhl�8�DB�D�}-"*f�lx���º1"Җ4j>�)�>7���s'�0�VYP�A!Đ��$�s5����iY
DۭM�wB*<��3jhgM/P�<:��1�~ch;���(zf%;��_����U;l��!��~5�èV�C������Q��E�L�u��yJVGB�c�����W��U�gMY��}��}�Z+��6��������̎Lu�ȼ��ڱB����@X�����~>�}�2�Eg�<OR�q�[��s��á�W�m��GT�6i@���ݓ�Vj���Ej*7��F���4�!�F!��c�����`x�v?N�1"��X؛7�uFwGs�ִ�/o�Щ��.E;+7��=�z%�eo7��A��G�%��^ӁC��Ȏ���T(H���B,����"�B^����ߔ�f�h�޾����������XR:ؐ���ەS��'�5�s_�M�e�lџ2+�����n~/�V)���x>���ETb�p�a9�׾��Ɲ���T���o)Y;q �N�@���c5a��`�L@QHq=�4�lĂ�Y3�%b�SǙ�
OSGt�9�Ɉ
/�mlu)����>�j��LxlR 0�$Xc�5߸0��CowM`Vm��e�Q{`T�55I���ɮ��i
Æ]�D���U'.�m,���0{�A��1��R������+��A��f�d:�Ä���bc<T�&ҢɶT�(_)R%e������XT8��,���A@QM�a��z�R
k�p{HT:�{׽���9�{���9�Ç�O7���]�y����
v�Dі�I�-��a�B�q�1�����3��@i���{�¤�wC5a�a��]$6���g>by��[���lᒠ(����x{@�NOl�z��o v�
³7��y@�VJ�f��J�<`���6�C�!Xm�Lf��bAf����)����|��p�ƺ������q���,Ă�,��X��)�$�K�f�d��sq��T�����1���w�&�V��c�f$���E���P@���N|�A���;R�ZU?x�+�s�r<R
Cv��v�NR�΍Y19d��Ns �hn�a��bA{�LJ�U%f�6�&�Sh���Ad�<s,�&0�
�"w�W�|+�+�u�� �o{�n܀u]��@���m:�r�i��ŠO�
��W}����͉�0�	nXs���:�����쾰��j�z���H�n�^q���Q��%v����+�4 �(��guQhM�+"T5q�{�gR���Ȧ�z�֫��h�9�����x2�h-N!��ڗ��� n�psV w��u�ѵ����;���⤬���{���)_��%�}�H�R�s�%jQ9��2�*n2�۹��C��w-��et�Cpi�h���;2:���r�ֹ�H���"�Ne���t��n���c�R�J8z�1��SPs-�V�[���GRd��Vv=�XT�ɢ��	yN^���� [�g�3v!;^W#��!����V�L�XE)y��1-ֵ�"��qT�
�rG�8"V<�����i͘�����&���̠[�ݢN�4m�g;z�(�k v���t���N��=��x�kl
7Ý`�7"۫���'�iC�wi��2��B1Մ���p���9�M=W�r��v_�,��v[ґ91�[�����M}c������r�����J�g� �uh���&-q4��ڽ�׭ŏ*i�_�~��g��/�@O'�W��e�ò[�����&���R� U>�@�*���5!�☏N��t��|M��A�2��Sr���]p�*ϥT���.�2����mI39nE�:� sy�4����3Cu�+y�H{o�1D*����u�R�"��N�[����F���N�\��{h�#b�v�]3d��!|���P�Oo�Z�"+i���oq�G�E,�`5��S�ҷٗ���R�Z/ A��b���d���d��%u�/~\'L
+�ݎ��E�r�D_K�@\^��$�]ځH؜�7�1�ڵ��p^fZbI�C���B ]G.vbBW\w�;��t��r9��S�)���� �|/{�`41rƵ�-��v�t��WF�m
-��&��;3l���zؼ`4���M���0���sl>��!��X��b��%�+��O4�k�77h�i�[1�
gss�y�CR���p�-�aa�_p�m�%�B����6+�uϹ}/��/�Z�=��v2�9WQ*t٩"�\�s�U�˱g$�	�������z��m�1�"���AW-q�b(�[l�.%�Q�Z�*�"����b(�T��-��R�Ķ�c1TLJ0Kj+pre\�r��2�q-��AV"�b;�f��D@��	ir����ne�\�c1+1���Pr�+s0E��Ll���(墊�DTQ�PG-UG�6*���+[PQb�b����DG5pFe*�[��E��dR�EPX"X��V��U�UR"��E���h�,]R�,WT-h�#EJ�*UR5�*��
1��E�b(����UKh��\�,Q�( ���i��z��
4+�xA��	q�עV���p6���Vr����`jӒ��I���@�Nu׽{׾�o�	������5י8L@�O;֊�r����Θi铔����%v��>�R
t��M��l�z��P��Ǧ=��f�+�J��., D
A|yg,4�Pߴ���c;�
�^o8g,�E8=�&� b���Mg�'\Y�0�ᓎwƈ,풧;��T�����=��u���;�p�=d��R�HV��͍ �S�d6� (��
���bGy��|�V.���NXp�PߴP�k�&$Ĩ��8������L%H��l�Z�]ٿ .<*<& ���Y��f�_X�Xv�RZq�;�+^2� �x����Ğ�G���M�c���
�H=�k�pR��l��30�|e.i}�1_L *ǻT��J�'��n�I�\{�V�1�hs��AH)�7�M (�����I�dѻ1:@��a�
�ɤ�to̓L풸�^f�i���<�|�w�xq��H)�M�X#&�R��ÅB�+Ʋ���p8@Q`h��x�bAy`\���!����IY�՚g��t��I+�� `U\��a��ϸ���������<|-��=aY�o��x�z��R���<z�dS�M��SV�!Xz�|��
Az�SL;NY��1���`�@0<!O�0Z\���u��bi�${��3�l��!�E��T��w�8H,*=�6�a�
��Lz`Vx��]�s�S�
�ɮ����g�7� ��}{��5
g{�|��7�>c����xbAM�x���c �CG4=Nov��*%g�ý�� (�VT�m��P�-��La�vj�$�fO*�k�����;�z�{�q�*p�Xo�N�/�����l��j��钾'z���);C���ɶTN)����׶0+Y^���C��<��Y�`x��7��Ƽh��i�E?�K{��ji��X�"eb��`��.��4]-�q��!���r�"N�)Q����O��o:�h�L��0<���Dna��r�$�')�^�B�h[P���ث�NyOv�vEJ�z+�����s�?}�&|x��sgl4�P�a4ͲVN%�(r��v�Ω��k=ý�4���'����Xqi���U ��P4�dی�rMn��1���ގ��:�y�q�\�:��ا	���& (��R�혆��ăl��dY��`zԛB�^�1�,+
�ݞ�a�Aa�홺(��:.`m%~�1�b�u}�����֟j��{`��y�
��{��A�!^<����VJ�$�Ĝ��4�ALd��,��\�6�0��1N�1IY곉�(
,�N5��^<�뛛�}ߜ�IR
x��e��La��r �a�4�d�
hߚ�P*z�Y�ݓ��0�a^Y9;�:d�>�7�)4�ud�ɶT�pot��7�����\�8��8�X�R��1E�l��2{嘐ua�u���*AL����L�J�Gvb(r��>0���=}��e�̩�v���z�s����i�3~P�z���k�bp�S�M��偝Rwv�S����Af0�1t{�i �1����i �C��dX���ɩ�1'(Vq힩������w����g�@�����	��!�(�V3���6��`^;��&�]��4��T���R|��p�ܤ��+=I� ��� xD m��k�����|kqx`�X���c}���⁈J��m& (�rq�M&�IR�'��Ͳbw՝��Aa��gl�Gy�� T������g}ql��a��l_}�����8�q�0c��DL ����8k'�E �e�C',�)�r�׳���A`k�sL�����s@��0�ua�V���\xtxLB���+hUT��;�`ĕ��Vo�ERW��w�	��s|����<a^e�'yH,�,�����9���T����T��!]qC�z�$8���2$'��>�b�f�5��e�ޘ��"g.r��L��R����5��~:tV��h/q�A�oa=��[8>�6by/��ئqWӬ3��ݔw�|���z($U%�lWr�H�A^+*���< ���������x8����EC�1g��aǖ��+8�>fN
��u�y@Ăβ��a�Xb$��:5M3�J�^7`by 	�s��_��b��,��Α�#��p�̰8��Af�v��Ă��,6��d����{�-�A@�SέT��Xl�1:E%d�Y����6Ʉ'O7��o���Z�p��t�=��	�R$��;z��x��t�,��u͇��23�I�l�	�1�DG��`�1��� �l��H[H)�:a��P1 ��E�!�0���J�Y/aC�����ՑH,���8�V�i��&�^����M�UCç�u��L�o<��['I�LC�,]$���g��4@�V&!��1 ��j�&�
C��+z�0��恉=B��i�H,1�E7� `xFm�u��g����'�	�� 	f�醐�%|a��Y�J���5�S�
���)��L+�'�T�ʓ�\�	6�H)��m������@�c/��}�~<���^���)��,�RT���2����5�2z�l���ÖaR�f@Y�J�yd����85CI9d����B���'	���>�#3��}xǜ8����ό	����5<�H6��)���P�Aa��t�͡��yf$�1���Έ)�7�a���C���a橤���zb����G7���4y� \�}��q��8zC�Or����9d��J���T�k��$�z�a�z���{�i ����^�
�R���������e]+����x����:N�l�H):B��;�4�Xrs�����1��1��{�,4��Wi��L钤ה1��2z�2< ��4@�
��}���\vo�R<�6b��wd5�9�Q�a��`���B�r3-Xi3��{��t�o�u��o� f)�Y��<t�B���+���x�3�p[1 ��3�>�nr�"lv��Բ�����i�ڛu����&�箻��\�����g�-I���530铧,��s@�1��H(�c=T�N-�l��)+=�Y1��[f���9aP4wLH,ᒺ�{�m����ߞy�q�����&���p�R����8搬6�&����bAJ�ɏ���1%NP(���y4�{�.�U
�S�l��ef��uf"�S�x����o��u�>�}s����w纇l8a�
�O,��i+;g���E
�����~`�q�XB�ɫ�3�N���T1��T�%y�H)�N��O��\Rw֣�����=��zǢ<{�:eH,���� QH)�3I�3���X�����$�
��8>Y8@Qg�Xi;ꁉ9���4��E��WL:aP�%y;�{�\y����<�u���%C}P�_6Ã�4�ݰ�1��NN��Y�m�$�TY:�Y��M��a繄(����l8H,8��v�*_6w�o�9����}8d�*v�J�V2t�l��y'<aRr�H,�'G7H
)�u��I:N2�<M�OL��08�\gl���ܢ��� �
 #�4��.�;��q\㍕��,���V*!�3 t�Vz�3�Xb)<g�i �s�3V����'!�J�8�I�:M����08�g���p�n��<�חz�|�yw��a�:d�(l��&��%La�z�U ���XVN�H>�1�L�1�F�1 �L�
)�c�1��d�Y�v�P�<"���6��˚3��U�-^����c�l�����0���!�i��E���XT1��p�f�*pZE�OSZ��C�d�vg��a��h��S�Iˉ6����xo]�s�wϾs�^ä퓷,٪bA���g�w�	���i�T�'��Y6ʛE�*Ad���o�Nz¡��&$z�A@QM�������e��I-���>�wc�A[n�.Ǝ����{T��k,�ͅ�7�/�N��o�ܜ�������ޕ*웴7�8�Ȥ\�d=� !agM���o]�'�
��� j���L�� .D*��8Ld啕��2{�ݤ���f��Ka�XmP�{L`m����{�E �tg�,*AI�t3V��!ָ�̽���;�}��ACĕݧL�E{��ôd��1��q��{�aXVi�yO++%M����*�񆭘�dۉ|��
�l�c8߹&��{�TKB�y]7��V~�@� D}�L=f$��3�%b�z��i �}�Y��1|9��L*oty���a}��Ri�aP�5�v��Ě=�@Qv���}��y��Ʒ��y���$2�uՆe!Xi6w�G�AHh�2v��t�rjɉ�&�a�9�R4=��ov�U��g������d�*m�HD{�.�dW����d/��ޟT{�<*<Wf�H,�u���4y�N*CG��Ed�d*k�:a��NSs�gL�񓃝�d���&�RVpY7Ň��I����n;��w�w޻�A`p�Vz�� (�9�3�$8�&j���O�P�AB����ᜲT���Ri��!��Lg,�g�'<Y�0�ᓝ�,������V�7�n�g��� d{#���'� o�gt�a�6���
Ae��!�p����(bi=���u߇4o�k&̃�t����q�}i�C#X�;ң�O�ñ�ѱ�)H#�d�K�=�kv�߲^�n�i �C�#\1�*�ϐ��������XU^61��l����r��c�s�������Qڱ�* ���L�u
��*�:*�t��7e���y�����Y7�A�՛!�u�^��Vz,l�ӯyu��1E,i1��{3#avH�u�M̬	�_� 8d
����6���I�'ݴw]av�Aj�/q����1L��=� <9թ|{���g�#�R���V�5~$h�S�Ǝר%O�`���I�k{���CR�E�=;� �W�4!H�8NGW��2%�Ǖ/,4;��|������Y�M�t�m��rL ��F' �=����^������=�Z>��ૌ�p�c6 U{i�����*b#��y��)���43�ha��V�C����墥��8BE�����m='2%��W����.�����>0|G������FWF.볗<���o`�O�R��8�&j�3�4�	�[�&���b��n.cY��9�h@/LlӘ��f+������庰�y����W[�ny����"D��R���*Q�i��cu�FV����d�w�y0X�ҡ��G�MCsc�#Z#=T�S:�-�>陉v�氞ЪIz�<#+�2�B�$�ܣOw\z�u�t�'B����vW�;v!mt(��L��f�&�Ev�Er�i.6F-�wӺ�[�军{z��5x�T�B>��j� �vgVݨ��&1\lV
��xx{�U=|�ɳUx�j#��e�p����Q^�JExE�i=�y�u�����<�B�4�x�ٵ7�
�O��P�=�r���x�K7��8k��|��<������/耫�CO�G@�g�:�R|���H���W,�
�x�|y�&E��j�Յ.��P^��h�XkI��;~>��!�Q��A�V�q������^D2Mq��B�_���B�e�V<�-o,G3Bә��yEC�l��!lױ�*�^Q�[�4"��><'mƗ!	�ڴ�1��|ͅXkF�?A�˅��X��t���@QM�br�Mw(�}D�v���g�VQiSĊ.�,8p�5a�_q��d�~4�:;�����n����0|Ξ��{�c�3$l��dlDӗ*)3����g>�lFH|N���p�B��*&��n�z�3�z��������@�]B��[��E�����i�`v���ʤ8M{��ʵw���Uٴ�
�=/,t�d';!xg Nw�v�\��Q�Ļ�}�]M�Y���w5M��J��w�z��X {���]�؞(���P%��!���,j�
�:B�H��Dł2UB�&s�J�6�cJr6"����aK��9j�l4)Ƕ:�U��/if�Vo���t��ʴ�]a���/�Ί��SA"*f�c�t�R���p~�P/,�ER>�%��d��2ˇ�q��%J�'nw
S��-{��SL)�&f�G3�4R�n��O�{Ɨ������Έ|j�����9ꄪC�
$��F�ev�3�l�)x���Jr5�������G����|��<1�m���c���v	8o���՛yVGQsR����V
r9I$[@NS��¶��(����K,�C������\�ecKw���|,{�Ձ�\5�ШV���^Ӂ^�nEr#�kͅB�o/,�YGsZ�
����"���+kb�nY������˚��JA�Ƞf�qG
��4�5�-��6�`)���d��h���=M��^*��j�S����k'i���W��g�&����ծ�Ӈfǚ:e�(���Ϙ��탑��VdO*o��+yp��|�� 7��;uV.��!Pt��&����S�LL��^_Z��]��r��o�o��"_��`5=�&��"�l�D�M�4��%ȣ=s��DͩA=�V�Bl��V��}�W��/�`x1�'C���_m�>�a3,d����f�*F)��2�,B��P"!�=t�d�,���wu���ۅFz�TR�5s��r69���)n}(@�F*�
Ws�T�rU˅�V<8|�Zeq�=��@�����+�a�����ϑ�Ŷٚ�(���Ο��q����:���>t�r�:���8���_�^�S��%m��9b��Ϯ�nF��nC��4�E�c�rm遬"nL(�����2ͳt��s��E^yM4��';�]��xCG@H�T:%I�� �>�MH�y	�W� ��[a�yhf�A�ɞ��;������bK�D5�t�LF��sSBHL����"6 T������tE"�b�x�b!}N�Q2K��]��0r���wQ#apV����׼w^�:����}�UU@Q|۽��c�D�;�Y;H(��T��t�.�BMʂ�v*��A��*:����і~�Z����O�M=g�O�ܼe֛�M����[L.�f&(E�]s~#+*�e�h|�ϣ
ׂ�e����OV�����*%�5�S�X??�3�i�B��5��g��+�,�M+��S�Y7��=bf6$�(*F �K�>�/�ϰ<�e�34���k�k�cd8��#=hқR$��R GG��>p::���8��j�F��E�"a\�1R�>�e�ђa
j�S�G�:�9=�};��R>��aa��ZQ�&2�^��!��NX��b!
���2�q�F{<r�ޤ-���'��3�o��tJ��EK!g�\ �v�:;������Cv|�`'ԪiV~d�VhJ�MyˊRC{�X��"�eLMD��^���r����l��1g�Ah�ip_tO�Z��)��Q;�٘ptkv��H�	kĬ������0Jh�i���@���P���[*=�\y����D�&op�*LZ��Q�o�ξm�{���0��{K.�I��\p��r���}�j��޳�DJ��(�cq��M�mP#v�ᝰ����h���c�w�(�n��yV�ͩ��4�<Ρm^�΃.�5дsY��A����V�j�em\aK�ݳ/��je��|x��A���_ABm��@:p�u˥�4y��۫�����9�]���X�i7K��F�]m�Ek�F�utG)AY�B-�f__J�
�We<�rf�Hrwf
�o�j���H�==�ǛzMsΐg!�P��vr c�D-i�p'�O���Y/�9���'J�T���.�Z�m۬���y
[uk-�����au��(ő��)�2`�j�ά{9���z:GE����ǈ,=�+戌���V�v��J���7*a��ڹSuo_݁�����Y*�c����(�hc�K�K���b̨*;8�P�Ow3|-1 �lg]�;tV<�P�a�ݞ/Wf�sw7k)���~��3�Oj[��|@�e�@�Ov�ͧ3�oF�U�N�_׿<:�Vr��N�*�کdZE2j٢�Ѫ�6z���ڷn�-���.=N뀛Xо#XX�v�[���o���л�SΖJ�u�|^�uv��l(��;@�5��a��V<�lד�VBop�͵�t��)m�Vh����M�W
6�(,uuͳ:pa��=��܈�J���"��$໎_>�s�7EX<-@�T�s�Vgl��-��Pj������5���gl���Şuu�$�0<P�$m���q\�_n��qؖ�ý�.�1x�
�pfۗ���dX��U%�
ȸfu�qG����N�g�w8Gv �"v`זce�ˬ�/������sX^�]]��2�-�4���oqYv�S%��s^v<�����]�yY\z�m���3����s��D���4F5qޭ�[n�3e�-���v�Q��[JKu}����S�2��n�L��t]���Y�d+bG��n�=tN�;Jud9�=b.<0���`����5QChɭY�UʶRX�$�~#Zc�,��-�*(�V�*"�TQm�������""0D�҉��UW)X� ���"�dE(���l�,b��*PE�6�X#�V�ƌQU�
�Z���i�8�*
��",b�TT�`�ZX����"�1X�E�X��KF��DamAK�XU�i�eJem���*	R�R��Y��X��L�Qb�����������[�V�(��F ���Qq�V1TT��*�1*�O8�����h���R]��������*�cT�x:w�R*s�,L'z���m͔�p�d�m.��&?� <=�Q�O�yY"���E�>��8�%q�2f�qϧ)�m�r����ő}{:�����Ā�b���u��v�)Wj��c�BOnP��׶���#v�g����|C���֚�C����/�S/�F�i��a�j�|b��B߳k�"�R����0��\n�B�J��A��j!p�Y�s�2���!]z�Y���ŊΡB�b2�(o:F��"�)I���k'y�p�̍���~�+�viɉ��'�
e�%߂c�j���<O���;�K�B����~*i�a�%
�=��x�Ȑ#ד��R��x�4��N�v�ʃ�C��Շs�(.��h�VZ��1�ps��V��=��)�� ����q���v|�̇�^�\Z���:�"�N�|EL�L�ל�����4}4���<��O���V�}�i�)�-�=��ƺ�� �r��Tr9}��Up��|}b�bIb�n�b�bȚ�zw2�W��i8W7���+ubo� ���'a��N��Wz��d���֡Z��'�]ہ��f�]�;��b��}��UU{gm�愑L���'!E�P`8��F��u�j��F��^=Ş�� �=�wz(�ώ�}�#M"j��iU��p��FEu�)T�M*5C�<�Z�f���j=*TNy�A����MC �������M\-�RȜ�WZ�j�ɉ���^l�0d8%��B�L9#�k)Ǜoңm�]�J�w{��5[@�#�C�!C�MS���8c�d*�"�-GZK��&q_kRJȘu��*�.�V�@Dq�����sB:<��8���a�G5�sW�cf}���
���xi��pc��Е-N��3��}&��|�cټQp+$Tt?]��%��e��/x��Ɗ�0�A�Ǩf�s���.AGm2}�J�m��&x��] P�K�"�J�qш`����r�+r}D�\�� dK���%�(��<z�b��X��hyuu��v�Y\'�a+��D=G�=/!���M�'������&�)n@���o�����S��ݧ�(�Ngt�n�<6PU��k:'/���`�Uo���x"�ԑ�_s2l�`+�p���T_ꯪ���ĥ;�=W?{'�3��uq�Tga�w]E�hq�Mb8*z*9��Af*7*�|���0�v�V$r��Ew3iP��m�������{&h��
��{k;��z���7�����Q�=�=��>����\��x�=nP��v�y\�(@��t�.�<Oەk�
j��o��%��#+zR�\������Hp0B���5�I`$}�U[+����r��~J{��U��o9��3��a3I2�{O�(��TNt��(t�ܗ#����׺335_%�@�uN:�8��0���L CT�[!ƈ��>'���j�����O��Z�s���h��VK��SE�ذ���*D4
�'˘�[�崵�ʠ9�; ����Y�d�*�F��k`��ܼ��������C���P���@h��(���>g�by�
b	�8Cr��!�7��Ed��\R@yP�֚vt�yݳڶ��5Ӑ�Dr\�Sy0����v�K
Mp:u��MH��R(4 ���U�Uw�+�B^�*	�%pݰ�o=��]d >g���ר#� ��s������a�R��?wu��x���S5�&3�┊�I��bao�E�zEj�"�_��F��p�Y���<��g[�@�vn������bU:���>&����ҹ:F�%I��I]^��b��0w_��T3+�G�i(0Y�=&��K;B��7�V:���F�75A�����e�����~�fw��$�u���H|�2z�.�>��T�O��.�nN�Hv���='��#HNJ��`�����=�����T�h�[*kTZ�z9j]	���=����옱BB�)s������˧a�����}������ ���f��<��}�����bQn�jR�B�참�!��g�7S�ôدWL�<�ʢF�Z��EO��L�tW^gg�W����>��LN�����J�sNy�0݅4 �":JYw ��v���yp��U�=��o7i���B��ϭ�]��o���g�*��Z�Wbe]����S�ҋ��� ]a�W�o�}��]���\JՂVl�4�3uM}�.��DG��u����<<:�^ts�쏽|C�T�EԽ����u�no8� ��E�O�Z�DUH/�=�����pW����0s��&��aM�n2��y�.��\�{C��~m�=�O��Q40��`x����*�a���v�d+r���Ț���ݛ�\M)E)��T�9#dD�CSHK�S~�L7;���'��*�)�6g*:�"�P}-(㎕�Mk>�[@H���8�����:�O�� vO��4�84f��NG�LJԇE��w��^_{ɭܫZ�<!Aɧ,t�(�ܥ�] �*\�SǨg
��y����1��]���)����ʬ����{�)q�]��8� oy�=ٴ���̟9�U�Ȍ�P��-LE��H�D[�;ؕ.5U�]+�Y&ldα>o��@ݛsu��^I��2�UʈsY�@��������E�IΑ���&���٧�L�u(��u��i<��|�B��T����Yk�Ie�6�ֻ����1�>=�����79#�W-���ᯓܮ%Lqɮ�س�m]���������{/H��X xl[�����5n��C�8��@�*��ص0���g
|un�������-��
w���^q��,��5�ۛ]��80�t;#1��-���Q�N6���Uu�C!��2��)�AN�H7C-�����v��y$p�|��ʞ����K��C鱿}Y�⧜���L¤�3i<��x�.qp��: ��ep��
����o�����C]�mS�Hh�E>��.��&@5w���w$D���G��E��|�$%:���ff����NFl��#Q�R�p6(:�J��Sc�ĈdtD�An�VSG���w�;��X�� �KI�.�p����TL9�"b{[ݨxL�i��UiG��0���ت%��j\B�ո���p�2��"�.��ڮ�s��0E+v+�T�و��`�T�hGG������(�K�V�s��p5k�W��1g�0U�(��u4m<�˔�������M��w����f�Y��>���e��or��o5Nǹ2��;�]����Ye��1#�D�{�"�+e�������X�a�N��C����\��pyV���@��>�BHE���w�����j��2�dy_R�SܥPx)9��^�P�������l9��}��ɔA�W.W���
�%\��!��xm_��WI_P6�!�����[�޼�v&=|���^5����*�pwj*ūa���Oʱ���4���F�0FC�0�cɣ�J�8ʌ���/E{�0��j��o�C��e�E_39ѱ��+��HjH�Wq6�
�P�N&;��*�L��yj���x���N���P��-�U��
�ܫZ
иkY]��뮿AQw�x��,s%�˰�VO���A��*ɱ�#�*~x����Et����TK�y����oij�٫;
H��H��@��s@ϑ�*'gcQQ�� B�w1�|�+&�#=��y��kO�S!g�Ι��ɏ<�u�����N䭤*+��K���6-��Р�Ӳ+
�\�v�*̷W��.34j��9�FDyln�;Zw`{���;��������R/�.� (�;{l�q�Vs�9�����{�O,�����􉍁�J��j}s)Oށ0�ED�lTC��I��7'g0Q��{8:Rz(l�!�����E#�-��2�h��P"!�TFu�9ѹ[�/szX>.@̗ ��1x�D#.@�#X�X���9�Ӷ�/^ub�ַ��o��P����@p_�������U4��P�p��������}�jyл�b�GI�&j���C�R({$�s�0��B)h���[�j��s*"T�G�3؈n����t਌���|����mh,�=Y�=�Q�*��eJ��+����DO�,�sR9�;%���l������P�a�5�'�ӧ�q]��u��}�E"����O�[ۛ��V,3�hsyֈ�T�^�ugq�@���������fF��w��*����0of̃�U
��ȶ�Gp|��Ѣ���X�=�}�e%̙���êc�[Gi�9X:ڼ<z��/֢�Ǝݮ.LOu��\��NH���d�
��b�\�n���f)䧗]9�H��Z&��o-��).�^��T����s'`|�鐣�{��̥������|��Y����N��S˼Jޓ�g#(H���`.=V�ԏ��v�Ex�Q-׏�R�Fe�����������p�u�{���ȞHu�d��F9 �B�
���v��$n�@�����t?\��3n\	��	:8d�w���B�C��7�o�i�fg��C��2,mut]K�qb�=��n[����j���q,�>��<����^�#O�V)���������!W�׵�qL�v_]�,�ĺ����ʤ����
f�2��T>�k����=����P6m�I]�X�I��-M�^����x~uD���5�=C�qy7,U�^MbY���
���-�C�S��+�iE����}7Y�{�N�m���'8��4I�*@S�,@<�9��!�>h�шqC�!�ՍW��%�7z��t�x'��������6��u����N{lX������S$O�j�ΉSq���8
�A��g�bZ��p�r���9b��NS��Ʒs&6.Pݛ�_�� J��X��To۽cb�+����c��( D��KSAq4�EuD�fK��M�::� �
y��_H�X���[z��Yc�z.3Z� !Yp:�\�c������y�.�t�9��)�0Y(F^�!�j��X׽�N��=�;X4���B�9��>T�W�ٷ'$¸�h�P���7�'�Ī�\�Y���퐢�͋u��C5w^�!�a�>�=���nM��]�d�P^���ᴅg���dxhϴ���(/�SѢYj�>��g��8�kS����\�7흲����]yC�̸��MzN�O��j]<w�if�!�Єľ�$�z�z3��*�_M����}�}�O9nME�%T]�;�ޜ��^�?{�r��`����hU��r�7{:ֵA��\�^�������tW2�k��� ̌�dp?�ׇ�Xz*�Ϯ��E7W{ ��ϭ��;Ǣ��	�(��6"�7�,�p]��/��3��ǧ)	Y�`�Ⱦ���`�\`�%�K�|h�;X��$���+7 �'�pY�׍>�Do.�l_q��gEH����K����s]]=��_d�w%��q����3S�k��6|��̫Y�S�=S����֮�$�jء�C�R�lu4.�r^e�/�b�p7՝y6�Pp��ȉ�QE���c�r�zC����,�ofv�F��yc1�\�9Sw��䈛iv�iŶ����1�:N����p�-q�^^�͸���*"4���u���Y�H��H��e�����o^�0@-X�;О:�l�����0h�02[J�^�s��#^����5l�3����T`G�el{�Rs��(c�ޤMU��ŧ����ռ.*M8 զ��ɗ,+����uD5��S���־| ��{il�t�����]4�Nb3!2V����]�8�/���Ц.��G�
�굽w�KZ�*�W#ˊ"nc�pZ�6<U	R��Y�coyes/J�H]�TUM�C�@\T�˙���F��M�����kn��{�= �����SX���J+bw�d���ՇZ�<��Pn���g�����!YR���F��z8*�"Lo:�7Z�Sݜ��<U�W�:N�lP��R8�R�3�r�u�.�a������NQ���v��h-;9s��:k�bR�'������Beepp�n�(!�(͇|�ume��<r�:�c�!w���x�']y�ؔ6�,Y��];�����gF�1�p��.`�G�7y�B!u�����;�ð�<��5�U����F��jvp��k��*�gC�]boYo!�B�)y�2�3�䬁7[w��][人����J4����CV��er�x��e��>�W{m�ϡ�x���*��4�:��K`lU�lmWJ=��l*��$�:�CI�A�*f���lBI�ּ�Ȯrk"���!wl ���J�L�����3�Xֹ�}o�	5{}���������g:��	}%�����iU37�[B�""CY�u-�8�[��p���chT����>xƖ��N��1�
�=;%�!1��X���}N휴�vm��s��9�DD`����f��)�^���DE� �6�j���%b���jUF,Fҳ�*�ETD�TP�X��QQ�,DƠ�" Ŋ�+R�F1խe(�Ŋ���11f3N,(.!F
�PU #V,��q)��r帢�Vf+D][�Db$QA@�DY-� ��Q\gY`� �馩U"qJ:�X��"�X�",b�**궃�TTU�Z�E[j"�V���5�`�
���V\(QDEdm
Ŋ%�����&o>��$%�E^X�ԈAj7Ω��w{�U�
����wge;_�Q�]�Ѓ��J�����MB��ݻ�����v4�"1ɏh(����1Ң��MC":j�r�4�2���֯z *��Ŭ��2��X�H�1b�p���T	�$v�V����(t{�)WG�>"���`�,@�R�T�bc�)^aȍ��oe'���d[�Ң`���h��[1��C�5��R�9�GG��S�9�[�{�����Դx!�I�	s�9��U�4��1��Lˠ�yL#�����l��¦��>Kv�,6*lU����%�uϼD=�^����3o��p��%�$>���$-����}3�>�Lښ��W��*�W�n��5���h�>��p,�����:��ӵ���ǮE���)I/J4�M�g_�;B��r���|��ɉZ��_h3[M
��T⦑\[��a�[}��A�s�h��	Nl�����u���=�|���DD�oy�`��2������ټ���N��U�Y�tP������#.�K+���䍛v��;=qk���Wg*���O�������E�f���0��%hF�����i犹��]���a��:�TZ���/&bb�����%��5�l��A�p�u{_�7}��54�k��/$0��3\®�Og!�g�~X.j�]��)���&^}�{���H��a�7�
�(А�N�X�G�T��ea��<�i��̼��UE>>��Ѐ���ƒ8�q5�����s��+֊��QQGc�F�q9"a@�%Bc�9�L�>�A��ب� l,kMT����_jN�ꊍ�:r0�엲(�[��TX�!�� $j�z��}ɷ�N��P�_�N��jʎ����*�F�>�GT2�fm�K;u�$�7g"2_�O��b�J�b@xW�+O������� *�8(V��B�>������Z��3�$�\�}�'dW�j�LH�d�nz%!P;1d[����pa�uTD��]al��ҷ�\�]<����|��Xuɟ,^l��@
}�&-�vN�#�	dys-hV��6����S�>��
�X�&�:R\�kDѬ�'J��*)�s^5�mn��^�S&�U�.�������x�Kr6���۾X���{��ųwy�Q�1C5۩x���⫵�c!Wb ��oU��M�{��9�n;Sf-���P�:c,@0��P�j�)*M�q<�Ǟ��[@����n�.���/�]K3�p^�2�XS�'a)��{�T���0�Te4���띉|���T����YgźC�*é�`l����4`��-w�N�K�e)�����is!Ƿ�;s�5"`8[��a���z�[���0�7��N���;�ea���M�>���*j�Nʈ�}����;��[m�J��i�P�Z)}�镧��H�W�ղ��@�1�<�R�Fl��M�.sї� ;�^�%�9
��Qc�.�j���q;��읛կXrA،��9労>~z#=��3^��Oؾ�~�^�Q�p��^�2z�s��r����H~`�8�+��*��pɪ���/���e���R��!�a�A�c��ʼv�at$6"{:e�j��ba�=t�2���tU�_F��B���o�ZN�BS�o:��������nw���u!+&�r0�{����8�����N�.N���jtAH�F��y}�aD��zP�˃�}�Q�3Ԩg�ܲ��E.���0slmĘ �[��\��\^�3IW����^�y8�R�^��tr�"3��t�^�nb)��>j�Bq£��ɉT�Ǝ�0n�9����<@�j���&��9�9jbјLC������y��6�k�mv;���$(��NX�1
�s⥩����vi�GV�=���dDd1ʑ
�j���u�G�b[��n�>Ϭ�����s@����73�O��C^�*d����fx�ȴO�0St(Y(FXZ����v�o��b�N��o�o���c"�L�叅x�ݛs~�5
�I�P�K��B�]�Wc�Q7��7=�8��6-��_�~i��YǑ��!�{#��ٗ�=����dx�3�r�lV�V �b�:,A�p����ʮ��t2R=�s����(��\˅ j�Z�U��
�	vR�Ҟ=?�^���Śd��֓�Z��]nz�C��o��U��3�QoS�]ҭΔ�ݷ6�0�}]�V�n�u4
���}��O�}��8�߄��Z>�}��ug��W���ps.-`U���;��zj��><�I���(F�'�\x�=�D*�N)�~~+>�*���S:����@"/p~?h���9@���*Ъ��>��Q�6��f�)52^�����W.�l���T!�0L�� �ñN�� G*wK�M�X��0T>�ꭌ��r�V�V�wS����б䆭a\��1��ˋX.�`7"�%���nb��F!Ev���qV�-}�j�)b��4�G��i�0��[@�xÆ!C�X��XlD�})t;>���p�Y���[1�8�rF�z(K0�0�[u�e>�LuUG�W�o�CxR�1��\��)�(��M��"��:b.�	H��̒��%�K�/4*h����S��A�}'?��/x��s�֕�a�V�5�n:�^K�y��|
�|7�y� �4���@C�7�&��Q�|]#\=�b�q̀l"��=�g����9:�vOqu�{*�\ewmsT�u����w�$�������V���L|8�l�|ʁ+S&��v�����?Bg=�aA�L�s��i�'n�U�C�x:�������WGC�1���J�հ�=ՇrIZ����l���q�ό}46|�>��PMk�M��U��j/\z���n���::kG�V��x0��'�u��q_U⧲mP�����]s��36���9��z�5��R�2�BS��wih��7�������:t�i�r��K܃pO)Ȏ�l#��OE�*"���_ua�O���V��#xک�	�x��9�W!@�1�;A;��W�!/��¦'.��]�T�=����ʅ�R.eĽ>�cd*�M������:���B؄|T�"��	]R�ӎ}��[�D!��Q4b�v��K��v�ġMx�?���ߣ���K��%�21̶v5Qb.��W�{Kרu̠*;0v�>qc��Ϯ��]5@fRw�X����b\�s����y�����ţ���)�Wd�1W��Y�֎��;�y;�3[�n�d)������f~у�7���
Ƞ��l��Fp��7��h9 �dq�[��-K�uϟ2b�� ��|��S�*��\>t�zg�ԫ�[1y���k���6u������١�f��,wI�3P�F(C�R+�r+!ڪ�d��ngG)jLp�b�"HG��A�+L�.F���8*R2�dĹw�U�rn{ɭ����,@a#$8b��eɋL�J��-3��f�Zg��ŷ:��ĳ-��%�"��c@���j��I]Qg+K�hQ��a:�t�R��T��X6H�[B��cg5*W����W�_[z�^�~{��Rl��k��59M�3���u�Tw���󜝸�4�.�}��:�T��dgW�v����v���$?W0�qa�lu(]H�U;`�u��ͪ���>*A5�o:X�&DF0p�U��9DuD=��������H�K]m>�y\�y���4����)��!W[�uq��g\kdɖRWk����9_͜��Z_���j_&�)WuG~�=W�G=�S�o�;�Ꝣ�I�p*>w�g�i��%��r�]�%5�-�tږ�H/�#a�_��X�)J��|o���������:�m�o�-�<�wjW�9k��]�W�{{-�WE�,8�`�>�r�3gsB�P>����z�<=m�Q�{i-Ʒ/7�Φ!�	7)�zPG�*��R9S�iѦ�yQ�Z:u��E�c�6kL��^��9Z$e����I��є{���(F� s���^���� ̽�na�~ņMe��T�,�6+���䦠�Q��NGq�y}Ɇj�d�F��\�T������ܦ�u�B�m�<���� �@EWc�r��H�6MmFB��[Mؔ�b���[�'
��F01�r����12�h��d�M�R��KQ��j�s]a8e�Ֆ_*k�̞��f�Uد�}T��;��X"��:��\:sәJ��M�B��7Xż��U�ٙ��,4����#�A��j�
1�n�^��7�ʕ�Zb�I�v����qS�ɾ;\�2��+}+U��k��(�~ޞ&�c����+��)n��h ޾:1(݅�Y��
�ɰe3]�S]C_^�/P��WaW{�FU��i��F�z�+�@�ާߒVYs����T�U�$�|Ӿ/v)�o����l���+z�v�"�wv�qx���)���R�⩷��/j3�@���:W7:Ѯ��&��j�Y����ZV���ul�@���(�3������C��KӢ�Ze�$KeK&��A��1��M�P�ީ�L��Do�KrNS+	{{Ych�����	 %�9�#)_��pl��õ�S�?y*x�����MG9t��c�p�B��x����cc����e�v�T��mr@ΚW����M�ud�#1�\�����,q��L#n�GYuvws�M�Ɵ3����1A���t�C��αӣ���ʩu��,��,D��#����嬦Q�-��@�7��(��k����p�_Dν�B�!�a��G�O����i��m��Q�p�s�IJ%uE��.&s*���3���g��-�z����0���n0��j�qRU�]J��T�0�e��+�������i��A�jU�Ut��訽ܣ�ȱ%�i���v�w���7���V��w:O&���k���:�G�8�s��Sa.�JP�Ȃ#�s�W>���P�w$�[i��[��;{hr�ˠ�P����B�����������,�Ք3��RkN>���$
w�u"c�4n��b��m#�u�)"�R��˛���4���|-Tg6��v�M�����֞d60o'��f�r�F���G+b�wXg��
���at��/�4r�G.��י͹OP��,�Ks�z�.e�|��Ƅv7�X�Z)���=x#}��[WVv��ʞ+�|]7�^�	y��ҽ��B��W���5�t���0u�hEIY���f���T����Ҝf�!��[!V:3x�k�91=����cz�p�Oeb�Mk(v��B͠���M�ީA�
�ꚺ��J�{ב�J����Hr��tŌL�ؐ,.)p�R����ۻ�zV��8�K�5��PخZ��}�N��=�x�{e�XwR�A���"��:��MΏU�ޮ;@ �y�唭���/&@�ձn���@n�r���A ��X��N+|m:~�f�n���%<�A����p'~l�E2�����E�,e��Z֣����(_t����o3���i1]�+�_3rn\�׹���n��bN�y��M�Y�w .��/lGi���hu��|wzc�+�ٛ��
�Z�
����T���۩شȟV��z$+��p:�L0>��̦p$̦VZ:*��#��m�Oz�&Eq�iw"�M��@SCY��u��7�����w j�gn	%d���̗r�V��#��sA��wz�iE���zf��B3�z��즢゙'8�����ϺB/j��Nyܨ�*��!����ѽ2���<
|��!Z�(��(�3�m�5�Ko�y���|;��ۭ��t�J�ю��9F�Oa�v�@ӧ͙9V�,��9GT�R���v)�8�$"�^�q����%�l[��d"�\�@����u���vU���m:O]V�́�V�rɭ��l�|�ݳt���(�X�jWҤ7�Ԇ��'W���b����R��`��!��\U[�ʗ���ջ�/�]�f=I]&5�$���!i΢���%�J���b�H�j�AN6AOn��,���7v�6�EA���K�Ř���j�d�Z��q.y���=@h�,��&���i��wr*Q�
X�)���]H����$����" �LO�3���,�*�TPY*��Ub�J���(���ֱĢ�UC)TU���T,h��X�*�5��l*�"��(**,��Z�E�+T`����E�PQAF,E�����je,DAPQ`T�"��,�Fz�cx��(.!Q�PU"�R��11YRVZR�Z�+��Em�B�R�-,m�E*T���B��T��E���R��̵E`��`ZRڠ(�Ȳ��`�cQ��-�8B��/�l�YYR,�lFW��/'>m뾸֯}u��f�ӶG%��p�rհ���U�Tv�Msx�-Nr�R+��o���4_�>��՛����M��B�򶻕+
z �CGF����ީO�3ZF�S�^'6�[�ԥp\Rp�q�5KS��n�%�U�H��r�챧�[E5���0�p��p�g�����q�l�s�x5�{�P�[x�͸o�bUC{W��/�7�U��/�Tte�y���(�5ü��O���L�{ܮ�X��|;�TS��;7�!≳��F6_��0e�խث����6B�r�9�A��O�յ+�[�mgS{mU^�|_W�X<�ͮ�Y�pD6�@1Yg��DS]����:�K|�,�rBjW[5�'��l�z��t�P�og����R���y��(X�d�$�x)Ʊ��ԅ��l������u�7�X͸[}�Ķ7�&d�GB-��
6�f��\ۯ�QLԥj)��%��g,�#��)�'*J�S{$�z6�F�Vv������u=n�/�c��P9�A��y����Wt�w�wN����[]6�Fۂ7�����6���hns�+�2��م��������y���ڷ��Y��$X|��=�����B��X��n摽�����J)�N߮�n/36�f������a�r�Ӳ������WN��C��n��Q�z�����w]��{��Z�o�c�Զ�TI�| 掗ϖ:6�@E�j\N�M�^�y�Z3�����6��|���[�w��ޟO���Y]�3�=�Gu��N�17��������ߠntІ��V�ي�������M2�-&ST"X!&���8��."��z���D8���<NEd_C�c�S���9N�u���o��}m�T���&|��8C��G�Ǜ=ۦ������Y��
N"��S1�Nk4��,�ڕQ×����xuYܡ�	��
^���X��A��8+���4�;U�}��^уlo)5�&�u�P������s3�X$]Ҷ�Ln��<��W����3��s55�ol�N	�I{����H�;�]/=T���4�9M�몜�z�_>\e��%����iJ�PKx ���G�m�gIO�%��+0�u�J���Z�>7i�����آ~��P{�r���Ezl�{Mr�6�t^P|+Mo��ը$)WE_;��h���9Khomm��[q�%���L2m�b7�R�K�|U�^^�y2q4(w����C�KR��<�lR�}�%�Y����:��;��ҕx�׺߲6_O�0�X�+g*�� 8��9_.��9}f2�Hj��$ּN^7��;ν9�����iem��t��	+�:������)U�#
̤b.�r�U���S3y��j{��#�6�OB�&,3;Ʒ�Wgm��0�o\W�m.S����紻{L�A������&j�wZ�ܶ�Q]��wW9���t�imy���b�R���5m�/Fr���;z�&��N��GH�M�e����R�I�)��}�5�a̞J]�7�Ď��m�M��v�,q��?P��}���k��`���eGU7#I���[�Y��2����X��o{1�ˀ�0�ͅ$$Z8�w�i�n[�B���qӥ��׍��
uD��]S�ґ;��*M��"}�vN�)�V�+oS�J%uA����̦�����ˋ{��u#㒒����eM�`��C��7N���=)�������#j���Pb�~�2+���[�شP\A�k/�5��n��ny�(k�Ş6���)u6¹��S�B�N�kq�V�˔N��Zyr�g���*��7��,�BF`��&��LC�?M�Vp���.�w��F�]*¸ݍr���|�7��ދ9��d��t�Ɣ��,���\4E�3T�:�]kJҗ��oܜp�H�ɚN5W:Es���S��L2w�I���\�T��q�utb�L�Vy��::l[�N�98&êz���ܩ(�CG����<�m�	ښ��Ԧ;#���n���+╹pq�N]K���$~��8F���[E5����W(SU�
ȁ�-�}�%sf^�7�zF�a�-g�eP6�-�W{Vˋ�]�X��LPco�P+�c�#!��o���j�vv��i�b�����r�:)���{f���8��� A�]����ʿ{�Q�]$�f���DQ�3�]4~��O9�3yF��<rc��H�>i� ߕv)�@<�-�@��J��sJ��|��N�#8�:Ykx]�#�p(��3|��>ɷ���љ�q��}C;����;��N�&u0��s�4�x��ݲ�,��\ΐny�oob�}Z�"G6WDH[��*��O3R��8��÷f�3��e69gK���ꍍv�xV>;fc8Cwu�q�YVVcCr�u�#Z͉���5Z�T���t�T�ʰl�ohY���V �̜��XMGoV���
�z�����j���NI5�������}�}9�IĲk�z����'*-����}�qW`rb��j��tk}��i��gF�n,>��������Q4`I��wv {ᦲ�M�D=c�s+�z�#�:vM����<�Ɔ��ۑ�H�FR��=�	Me>Vʫ�*��b�-Q�\O9{�b�s�n�(9)+%%�P�dr�T�-�z�[��G�W�6�^��Q������N�
�фB�+[�Eђ����tLX���6�:+8r-Y6��,�6��Έ����_y�m)r�-g�R%d>უ��;ŗұo��A�b6Wt4̧z�&1�j�l�ۍ�=��&��_��K�]*�F��X�3i��&�i�E&��������wz+�2��D+���5i���֏S���K	7)�p����v"j����]~���U{��cX��A�i�d��K ��m�p�B�1�]�Ɯ�#�z!��H��鉷�7PuU/v	��y&�Z��^��.7��짷���e�;������s��%��i�UD�����q޴�i>��K*O�T�.1vV�$Sq�ݤ��[\��`�3�#5:
�Ut��u�>]j��J�d��C����- º���ͼ������̿����Gb��X�GQ�-^���v��%d����N;�]u�hrK-A�s}R��4tsn�gY�nr�v.oV�5y��x���Oݹ�i����֬;C�Q���}��S������"+�6��^.��J�f���۵>���٭'*�v�x,;��ڪޯM]�ᦖ�T���9�Nu;��M��{�*k^S\վ�9[�6�L�����-+t!��^�Kr>�J��������}�J�ϧ�"/z7�[�~�N�)0;8�Qz�Qѫ`"�1a�ޭ�(tVC���[���by����U�Tۃ��{VNv��z�9R�~��{@��J}���e��X�R�jB�>�)繷˛
hr3\����Ӧvr[!K$�&��q��5աf�ii���m�2�pmX��IPI�D�{\��7�W;����R�(3��	�Q6x�n�h�cd3�,b�Oݓɷ���!<م�Z�o�vfIȄj �h��NY�[���ؘ��_�^���~��2��Z�9�zq��v���Mw�:���	���y��5�F��Ɓ
gA�F�Y\d��Jě���9iql���`�B��-}�\��E2��Eo2�&cowv�������!t -�Bṕ��h�[�3Z�AU�|�6{m�J�J�[s��(��Z�ȹV��k;����bw+z��P�Ɓ��T�Wҧ�fh(���bzS�T��T�{JrpR�M�A���(J���[y�ҽW�rX��7@NVt�\��Pĳg���̒\���<�z��gm��S��#��h'��ϸ��R�)�K�_,�복��{�rڭ��ꑣ��2�TD��Ž�5�I�[Xx���x�em�J��b�ݢ���޵�����V���l�sY�|E��.)8q�2rC�95s/�lv�K���D� ���_`��&eˍ�v��{�zs�{M�.�YWlq������ݗ�x����.8)`͹����i������7�:�2��f�_2nݮ�N�)[)=�yDQ��6I|=�>��fq�,��!e[E=o�an_NZ\��v��J���z��P�D�D�HZ�YU�i��U�f�޴j3� �O���(�H6�\�nKN�����-x�"}:ϡ�@I�E8�6+�;P�B��!e=l���'���p��8�+��:�N+��B��I��W�v���36in[�>�#��.�s��Zf�<.!zG�;H��7��M���r�sI��"��N<w�Wf�%k����/:'�){�gW��Ҵ����eu䰥Nq��j��T�ʚ��m������W&�ۮVm1�#i]WZ���`�	�n�2�N0-�����o!(��L\�������C�`��X�,+�-iY��`]��n0���Z�h��ܬ�[�T�
��u�em%E�j�����#8�Y%��-����"֗q�5���c��䫺�2�`��6
kdQc/�L�{%Y�%t�C)ATd�z�@䷊��Z��λL�����1W>��1�+ׅ��2��ܷF�,R}׋�t��o��5���jV����ԭ�D� �t���*��2 7[KM_w
���z��3;T� 5�M>��V[��1rr����"���y���v�9Y� H��{�ڹ֕nf({E�]P�9�RVda&�U��D��ۤn���i�4�z�J���(qR�;53j��tU�XGF�޷R�_]�bս��pJp<�#"v��3�-���f�
؊n�ŀ� ���sł�|]�N�]��XR���He�ے�sp�(m[U�e�gx}>�1�G4j��������$_6�m\噖�l��u���஝�`	յ���^��m�������9�dU�d�#�X���W���홉>AjI={�,qTT)�6Ծ:��#��evEJ\�8�r�wlB�D�|�����w^�������&A�f֬�`_z��u�!������jn��
s�0�Āy�W�eZ�2Fv,�@�OgZ���*w\�z�Do��a��YܘL޶_�1�0��]����P9��}�cvﶝ�����m�$۴q(����H��(D�o	��9���-h`1��BB���gv��R!Ϯ��b�{�\�����W#�m����KZk^r�����d�7��|�n��fH��n,ݸk`U۠�k�ZΒ�d.n�;u�^ �.��im�J�}��+?�:��3Vq^O���=8m?�7�΍0�M�����l���.��\��n��J\�m�n�}:>�%���E@�w2��dą��Mm#A���-���v��vvU�ش>�&Ρ˂�[�3#��q+���/Z��gebá�z��wTY��;�b{�r���Zt����֌\0G�elɴe.Bz����e��gb��}�C��-�ES��;̖ͮ]89qL�v*s��˒��n�;��]X��=��㢪S�:�꾸��<�.�Iva�z�� D�H#�2/�E2�q��Q\�klZȉP+�T,�*����,�ZȫX����YF��P
�JAHTZ�E�ղ�X�[EZ���V�
�����
 �*�@XVJRԔB��j�X*�bWE%@Z��ūV�6� �1��V*+3
�
,Y�)P�U4�YX��V+j���Y�
�±dR�YV�Z���0�PE%B�P�
XZ�ԊE ��V���Db�cݘ�,++U�q�AH��d������!�P+mP���A����LG)�Z#%mj�*K�X�P�\�J�-�*�,�XJ�AHi*8�m�ל�|�v��_AǺ���K�V�3��tک؎��1a��l����)�"��sK���nj�����ٯ����-���{֜�g��\U�8;��O_p����J�}��4�Z�zKʭ���>��7�r�'.�S݀SF�H�=�\��ٳ�G\|8�>0���{t�0�'BF�D�V+���	Me>[�8�X���Y�b�G}8����}Eb'2T�:�ϣn�K*S�N�-�(Sn?w��M����y�^I��խ��u��|����)6(����l�ڋ�w��ŕϒ�g��C��eS���`��x�PP�K��*6���yE�#DM.�eP�-�L�c�6
S'�V�+�F���޻l�?C�MY��r���{D����6ʸ��e:�^�C�V�WK3ۡP.��4�c�u��C��Gj\_d`�#��z��rЛ��֪�\�yN��nR��V橋5�,��5G�YX9ck�Lc�Pi]:��{m}�;��/��rM,w�7吧TJA��dI����Gp��؞�3n�[v�J���7+�!��D�et��R�����4�u�9b�W��f=\�}^w>�RQRB�1"��9��&W$���5y}�*���*�w��:�.���F��Ԃ;.൫��]l=^��le��v��WK0���g�b!*Y�I��BO��eK7S�\n
A�%�'�ܜ��k�����o9oJ~�ڎ
FL�V�w�7�!��Djꓩھ��|�����%�^��6���O��F�7����ܷ�7k~���ڒ�=lB$E�gz!�[���WI]}�*��,�Q�>k��T�_^m���B�����ҁb0�z$�,T 綰�2ۊ����xfyw��O7�y
�r���Ԇ@���U˙H��4%�c�Y�L�p:�"��n���	���T�uc�i��=�ڎ�>��wj,ld��7���X�&feD��ꕇ�R�m-�[�[,QJMH�F������/���B��Zt�դ�j��Uv)�X��Ɇn�v�b�Hr5D�GÆA%OJ�nˡ�Ws�T��i��N;���B�U7�(�4�*��p�Sé�����c�20��rԴ�55g-\wp'T���i�^q|Z�m�+��p���d���m�r����We5���~��g�{%�-�۝NJQ .��A��E4� �%����t!��U6��YVX�Ɓ��X��:�.#�q�j�7a���xT�N�;	��C(b�^C��f���vq�Vf�yJm�++q�b�@�NV��s�R}�t�cc^
�/i�:�cnE�(���AB���4�2��COA��N������]��Z�r�IZ���^*�<Ϛ��٭޾s;��ۜ7�'/�^Y��AK��99�Jf@_@*��Uҡ'>�Mi\��r�¾�m��Ӿ�*�P^�!��o��+���_ny�3=�w�U9��;��ЧS�b�_����s�Y�u��{X\�-{'o�W<��Z_
Aڌ�<�U��W_s��ݰK�r��EW���W��}��۩��<��ތ�&7�E�Vѭ�eC�&��Ycp��
�9{���ߙCQ���Q"!Gֲ��9ڛ�q��V�|��=<)�%{���:�m ��Y7[z��T�ePZau�Ca&.�O�k�],�p�2Ҟ�{~��0p�	X%�cX���8Ӫ�Tb;�UK�gs�Л{�k�80�����O���!��F�+���p#�2����$��e�\�"�&
��L����_Uĩ��=vDhv�V�.��� ;�dW���C�n(�����K�����k��]��ⷝ�\�0/�]��m����c��l����l�0�3�C�ΑVa�4��{=f��{Dm��8��ʲ򱡅bֽݧY�����B����k�K�L\��7��<3%íJz��Av��1b�/Z�s��GZ��K��Na%g���
o����t��j��S�9���9��(4���\�����*���Û�{FL�3�1M<qj>�����b[�r��H\Zl��;`���Is�V�W���4(�mm�y.�m�p|5�T$h��3Ȋ������ؙ��og��ͣS�-����D���0t[��;ŗԢ���^.p'�X�,K,�^�xo���6����qzD�/"zw4'��1
�*\� r4���'=��=9&���z��|=0gt�z�`3�-���n������x�����:��@t֔�3;���ۥ��d�� K_1�R}ْM�	Ҵ�ǲG��	ҟ�YJ��DM-��4���B**yΪ�5���G}ZH�d|,�B�T>�D��0�h��GYcn��=�-�VD�+hH��4ݠ���N���k��	�ӏR��~��3�	��T�ۭ� ��D����}����6�9����A�Y�De�L�V\l���TeD����Mpa�Q!��b��	\72�
��wlVVN���G���`t�n��ާ7�k����LY9CX�d�ًϷ�o�-���}��S����hG���2S-�n���S�V��5�\�Z�v�*�Xq��]��Rs9��z;�\Y��Xv��=�GK�)׾���<�m����r���lN�w�X�݋���Ad *֝�+w�����ڢ��s��D����j2�E��1/sk��ѽv���a�sg-�J)[��޸-y����)��CNM-U�d~��H?=��E�u
��e5�mZ�[�=6�UU�%.+u=��);�suC�AB�K>��Ug��Т�>��E?d�-o?��q���m���.��^��&,}��;�F����c���2�����6�����n?'5�ܱ��mMN�Ǽ�6紉��o�3ֺ�m-��ur�rv���\�ю�1��r��ZuG7�V�L�v�խ�&(=���p���]��a�sk��4���vc+\񉉼>���,�N�$l�C�Q&��Ұ���1nw;���1�
u�]O�%��tI�sRFYnվNh�1H�VS���@�z㛿.���J��R�5l2P���i2����V���2�C�λ�����ُ:�Q·�F-n"F�ll���_�k�H[�����!m�(%O��Y���.����m��[	6��ɴ��w�����<�rr'3�x}wf�:(tء����ڎ�]���t]Rjۂ�wf��Z���ƅ��T�j#UI���s�z�[Ѭ���Rg
�f�`��+9�iX����}��Xӎ�o
��7^�6�9hY���YW6�G=��?Ss9���E�m��o!ד4�T����{'\N�Ue>m%�N�USzz�%f�a�>�H.��^��ԴZn�%�j�L·�'��m���\�Ƨd�����^?r��� �ьN#)WI�ٕo����h�����3V2q��<�׾=�ϥ)�vP���g����{D]S���� J78m��1s����p���8�!q�\;]q�׭7+-���7Goo������M�^��Y��<]�=������	�]�@�-^�׽�Vz����y�9������=�;K��.ֺ�돠R��u�蝵�i_\�ݚ���w���Ż��\D�m2�6%{��Dp�3�@��΅��e�V���ڞצ\6
Oýk��2���`���;��OV���Ҹ{�]3�pn�C���6��톔+#҈�G׎H�Rm7���ϵ������]�������TĈqwMV]�I���)�C���5،7hE��kofXm���ذ��u�T�+�e�>�vu�(�N��W�&���C�'˪Ԉ\:L�U�d�ug<sS�{�٬�o9f��\�j��c�A��j�lQ��d�*����>�>�r��{
m�{�K<e��XY�\�C��<�U�v�z��}��@ί=�&!�.N�Z�7ۧ�2'Y�:��h�Xy/9���*��M�ҭ��=�)���;c2�i|����̡�+�79爹~g8\�t�
0�O���Bn�U��q	�f졖��kf�{�6�p��}W���9��q�ZF��V���or!����/��CU݃o܊�t�� `�6ȝ�O���g&��ˮ7u����z�Q�j�r��R�>������`P�g�95�=�<#o���6�׷ׯ�z����K���g����K�6��x)6(�6���{������dm �wP�U=0ݩ`�&��* i��.����9Cx��) 	��pd�m�^��Z1Y^��������wI�m�4���z�Y���ڭ�7j����w�ds�����Ф�H��Ne��e=���S�ڊ;Ϲ���맢���Q)���[�72����ϻ*�''li���!�Cg�API*?���$6���G.������p����)+�[V8u�-�j.o�h�����oǽ�7�Tz�V�:$��8��⫲�7��T��AKh)���U[[�D�Uz�b�!)��c�E��zz�n�ZU-=���|���Qv!\QK�¬=��f_	I.�6�ur�k�gD2>5r.l��Ո{��Ȁq�~�Q;� �5ڻ:"��R}�6%l�gu�����,� o2"zH���ٳ���O�{�F����=N^DW\�u�_q�W������w���ښM��|,��y[XA��)�J�Ab��܂�n*d0��	*���x0�i���V����I����=l �&ZUԲ2¶{w)8B�r��Ph��]<$J=���N^�d�à�Uy��x�V3-w@n�s���'��p�3*�B�M�L�t��Ÿv �(]h���7ʶ���;����>U+J�Ǭ�<չ�/$�J�V��S]u�+�6��3/��4Pd���4��e��;x�͈9l�m�e�lA�:.�Wqq��[y�e��+@U��d|6����s.u�X�Q�jY|��wb���:��8�l��m���Hs��c���b���Zh')(Հ���%�Ê�[)��c��_db�	�ܽ*Y�>)�l8�\�N�}��eu�+�N���.2{ʄ�����(4�)�Ҵe6��$�ѐD�x��[O�d`�n+���W�h�8+�1Ac:�tX�`W}R�+\�y��P��xm�V�����v]P��\�D����W�=�xV�"��SuK�ԀK�z���|r-]wu�I���`��i�Ip좍gPin���X����K���z������9gC[$q)[Hɔo��5	o�zxu^]�7�˖�5�쫱�ilV�/Wp��X�,�G,��-��ٔ�u�齤�-]3\��]r���,V�fŖ�"��1�B��u�u����_:�;�q� ������ͥ�੎�h�3��7`[e�ɐ���O���X�ј����k��83�Y�]#�0�%}�9RH�2����U��=�GW+�8/f�;J�qY�D;�@��!�+0v��y�﮼�ι߾H,�*���a�l�eU�(�LLL�E����UA�b����EJ�P4����H9J��bbbc"�*��a����Ъ��0�-�E��(� ���,�E�i!RQR�l��`�Ek�Q��B������Q���,0E�k+n�+Aq�Z*Ա/Wb�VJʬ��b��ZŅi[%�qi�
*ȼ8�IZ�,�X)�YQH�ib�3(*�bUrբ��+F�`�Ud��!Q��Uĕ��J�!�2&��Qq�,U�
�q*���Z[`��P�SI�!Q`v�|t�1���>�"����~Y����G��zsy�\�q�Jё�C�B�뵷���53{#�\b�w��o׷η�
4�{N�w=��2P>�n��S������t�uh�T�''wz�X^�ָ�u�=�4)����6��{(N�d���&(=��	�-4�6�7������ɮ}V�y>���o��䕆��^��y��Į91��>c�#��޵�kӽ���T;s�܈"������{kA��^��Y&�7�����r�-�``ش#��z�cA{t�%��!�r~��-���p�8�CG��d�'U�j��l��O��lˌH��>f�w���>o4M�=;<�}O��b3zTu.�Kin2�ѓP��ݹ���K�����}�45g��Q0�p��Ӫ8�ШK�fb������dF�oV�����rj2����յs܀�IZ�4<(�=Z�u�e�7z���Z�8��m�p<�Z1@o۪�*�Χ��j�$��;��_U@�-��;OR�=�˼�*wb�Ň�愠�]؈��j�k��>���Md�ϻ�w�����	�ZpD��}r�F�3<f�[�\곓�{<ЧX�!����O��r��V�%����i�(Ֆ�e���9�DH[��g��j�a>��nv���k�S����d�E�coS���j��,�v��L1�����gԖU���A����w�t>��Ҥ��-b�q�E<"����m��O6�6��4���̵�s�Xm�g�a)Q�ݩ<�u�e�#��{gi�ŚӃN4��I�֝UR�*r�k����~ٟ[W��ҵ�&~qo���]&ܾ_]���J������8Z��;B*���&��S0�<�:�v����̳j�>|��=�%Ҿ��>:IQX\�ڙ}p�y�|\�ǖ�,���^ν�*�-s,幏zNG���Q�zʸ�+��sM1�������.>�f�� <��9s��ɉ��wq����a�d1��N8�{��)�G��YJj��,�Vg��'�
=��c����l�*��a�m�ar�V�j��w(4������8����6��I��;|_��<��.�cJ�Ap�>��&f>P��)!s�-��r_Ť����WFG���yE���iu&U`��5����;�\S[�1�V>��g1�����ޚFl[n�P>�a0��%�|�-��ܹ;p�������A���ѹvZ�댵��kZu�7$.פ{e��\�9�V����.��z?{�J�ԡ\�[<�)a��և
T�w���&g_�+iV�}�R�$���)R�K���d�'�a�j�M��I�!�������K�d�_�*Zۜ����N˥{㾛����q��\:O�ʠl����f�j�;]�{׍ug�u�\)4����'N�-a�*��2���M��Hݝ������𸥺��ӱ�y���
�M9֨�Y��L�;K�3����������JrW��=�Nhf�?o������U�6^<^���BO�L��uEWJ��dN�ƻ�Q4
�7X�{�`��>7��:!sn!d#�	�dzv^�r.��]ɣwU9sX�÷��U|Sn-����
T*�s/h��s2#���Y\Vm-�]&Ɣ�&�^��j��.,���6j:}��P�S��KeKIR̊]G�o�e]�h�b���ti�\�~��PS�.�IU��=[4��ݔ'T�$;/bQ��Q��5z�����*Y�)V�{���KNɱy]t�̍I�wH�mj��y�;�e椂/���������͆n�?x��0�v"$=MgM��t��DZ]�'�WP�W$�Ѓ#�(��|Զ�7�;x����iX�a;�|�d.�%��y��D�9i-)�͋;�k���,qd��pS�%4W!l��2����n���)�y�Vyd1�M�jr�]Pm-7��cʻ��׉WB�7�j�b�j����Sq��w�{VcD�G�*�ܷ��n۰p�zi�mE������޷����}��={iFmFo�É����y0�8��3���&;'�i�y�a�*�oHۈ#'�����:�X�,�E���]�R��n�to����|�rPΥM|y9��~޲vm,n\�Ё������:1P�M�c�±��Gn>������{;��;]�ξ�6��xb�MHۋn�*(jv���u�t2�����EK����,�ˈ��}�����%jz1�W5������>�nm�2���6�Ԭ�;�ŭ��z��_��ާ,�@
��x�����}������%�E����h=c�F��5��H��iѩ��)�٘���%|������ℴb�$9�&��8��6�7y�^�z�i2��l&N�6/�K��W���ϻu�"n�ԥ��,�C�87�t9!�Z����an�v��W��;��,Ֆ��(�θ�l����q����J��:��,��N��7��cu9�&�e�݅^.�jYQ��"}�uSl�YV^V41%�}��P�t!�%�J}�q��Um!}��t�#D��v󟺳R7�$b�3ۻ�0�܃+%Y|���)]vm_g^�z��C%��;n��}��_*�mnu��++P1s�uJ�5d����XY�6l>���g'
�d��O�d��WS�����O��O{c�f��e�(��i���O�n�~�l|�?�9��5;ߚpiƑ�v+��8��u��: ��� Vte�4<�8�k��滢s/-��7��N�Za���l�>+H��r�Uow�V�t�z#5[�M%�Ү��XE�O"+���Q}��ɱd,옝�����|�V�H��p�"q�Q�>e�Q�#�7y��^]m:|C�6��C<҃��<3���Z����-�f�Jn��X��7�)my�I��+��G�0�AC��]o���#�������jSɇ��ܓ)�1� ܈�s�N:eK�Y��O�0wwlV��h=ۮ�Z���(��j�N�f��{b�X���lnϳ�Y]��U��6��v��۾t�����L��s!��_X&+�#Y-@;=��]	�v�3�On��r쏲VԎ�`�4�r�Ck�:��cxn��>�AUTd��0�<p��jK3M��pa�x\�2i�~�e��5�DwD���9� R��"z�,1���ɮt�>m���\#}�u�T�+�qU����Y՝<�^^j)>�k��%uF��ѲD�������کL�f�O����^W:��Du�!p�U�n�{�9)W=���ǅ���g�>3�Sl����M�|��3޾���,�L��̭�o�Mvz����<����>�Y{����#z����$nt�%��|n��i����K;�G�t��{�l��>�)Ar��̚5�oZNwsO5j��Gmh���2^�|�i����i2��5��v]u��dt�
j��_Y�]�om5�z�}s#"�K͕�-8��ӫ2F���V.�y^�s�c�oIFw�����,�>��{7}kyn�08��xo�W��\ۿ) w�4$�9��l6�1���jk���̴���m��7Y"���Y�k�����MZ��Jv��,�l;�$l�Tp��i�5P�!�m��2�������b6�Sժ^�7Ș�՘�q+�G����9�a�8�Pv�dV�X_$Sv��y"f}8��s�$�Jy��luk��ټ�;��8)�9����'���I��<�}�qn�4{�O�c)�\8M-��J�
`e��]:��n&�s&��b�u���y���)E�����㥺4=�[iA9�L]�7ƹ�GO���[����!�Y8����i#��K�� S*�E�AT�u?Y���Tэ�/@zn�7�zP�����^�O��q?C+t<}��=�f�R`��A�Q�`��sE��K���@(�wu 5��K�$z���q�]ݼ_�Ά�oA�ݵg	��h3x�*�̬����8^���3�ɭ��j�0�ۃ]_u8n1v��'ݏ�Nަ����2x���N��+��ٔց��r*������ԛifR��i�Z��sg��N��N���ԍ��sD��bnK��h�^�(�~Xc���X= ��))���M܃c����񕲹��+"|ٱ(O�{է�N��}�ug	�T��g�u�]N/���uU2�{�j3W1%�CVON�D9�M\��YY�reU<Ջwu��o8cRlP(KA�֨�­�V���Z~�Ƈ.���|�E�҆��xEv˳�N]f�o+�S����i; ��c�ܐ{	t���d}f��s��-Ά*/sE�dbp#3�)Ko��W����_w̄�/�zM!��k��p]^ c% �y(t�t+��pZ&�0f�E"�;�8��M�6}�4tY�SW,�S����5p$���a��Z.�N9�F���e�MH�ԩ������:�Q�38)���9R�6�u 3�(7�V���<��sF��WXc���Z�l��Aq�׋��f�bXZ�|e���0����[��8��#�w.��Yn�'�$;�Wp6a�4�[ݷ҇W{#���b�ЇGN��]Z��McPm�ƒ��w��9H��a�ֺݪ���l��a�y��mZ"�]ǜ�_JƚX��J|�3�ˤ���$˪��d>9u��/2���v �M����&Ȗ'y[Peq*c�7�[O
�+��nf��j��AE>wܩ�~)�Ӑ㡅1z�<M�ƹ(�Q���58��)e5�n+�b��+0����#���f�d��.W5�\\v���l-���`tM��m�M�Ɋ�
���Q��&���]nv��P�_.P;������e��.�]��[�\
{�^�ѳ��	��`��K��ڲ�(�SY�&�[ph�S��N�*@�����E���FZΙ5�"��9�!s;��Zs�a+a/0ɴa6����¢����C�9���P���V�VGS�{����_�r@����a�EZ�떿=���� ��3;��\q#�>N��K5����]r4��]FErp�<�_sj��Gv`WflN��>_n��Xv��/�뷬k� b�/f��@��^,�mf����|7z�)]S�yYo�%����O�����Y0�1�hv�*�p=Y���u܆�ŽdV��D���CRˈck%.�����l�h%�B��s�p���"�ZS&MZ�g���;+��G
c(�t�v��jgK��E��WVF���S����������:�m����7��jD�HՎx�]5������ʯk�9Z���bΣ�%��ecx0G�r�7L�	-i��r��l̝�W_!>"�p?��䒒�r�=�z��nq��y�y�^y�]"�@��egl<f�C*,U��P��jV�����V�6��������A`�T�XRT5JPTX#Z�qSHJ��J��AeAVJ�J�4�@QC"���RkVʂ�j�J�f���Vi���#��5�����a�q��J�h1�����J5�E!R�@�M!�Ddp���*�U��°�mP�&e���R)YP��h�������,�A��F-H*¡��4E�B��8�I-��Q�-��U�UdU�ԩ�JTRZYJ�mVB���HTY+111�ʒ���b5�,2�]Xi0CYa�1�1�`<u��*�5�'iq��UeL��jc}�IF�|��p�m홛��Tu��Y��c- �h�l[�[�����LO�r*��Y�X�!�C�&���ǲ�v91��k��4� ѼdR(Ֆ��(pv���C5T��sV��I�j�.�^!9�}fٻ�I�(Yn�;��(���u���X,��m��m�E�j�Yy�W��cn���k('�|��T��B�T���SSt����lOtӢ�8�J�s�'�����l��yY�=�\�jpL�1�d�,/{/'���-���������GܱkN;��e�W	m��!��0'�й)�^��m�7Z<ͅ������~���T��3P��
�7(֫��5�����U�Ckv�O1ӰZ�gʺcw|J\���{o �H"6皞Q��+]���}Z�He#;r�s�(�E|J�9��&3+c��38��u3���0�D��9�������wFw��)D����]օs;�)f�[t��󢡞�Y�ʉL%����+r'ֽ�3�Ӟ���w>[�~4-!s�-Rw&��׾�2:���u�Q��H�};S\ ���va�������K\���h%ckWE�c�ks�V2F3�lY��{9/�6�o!�F�mJ�^8���d�CxO��T��f����%���8�[q�WhVK�Z�fF��:N�}3��յ9N��n���ދs�J�of^4��T�!�C�\�FM�>�����t�.�jԷusO�YҤ���[�D��p�ʱ����J�H�;Il�圗u5�t:��
T���᳎5��)^^խ�L�3���s�b����5}A^�^�_][�7?E^�|*m�̳��GZ�M��X$��V�ҋ!�yT+�5�{��JJ���X�y��p�5��҃����� ����{�;�9����<���)y�)����e��u"�F���@U���2�Nh_<��Sof�G��/�ϛ��Z��^k�%B��o�聝^{FE}F�����O'~����](z�b���k��$�%uNV>{��xzӷ���F��{؛fw�cT���>�i�U��-�:CYo�㢹�aHY��3ġHaU��l�|A���Z}G������M���1Av�V)R�Ϙ�dM��O$E��+6��kjk��e����?�:�Cn�MC���P�U=%'���7T&Vw.Uq�7W?�B
�؏�9�MWj�r=u���O�W�hdC`��y3ػA.���If�O+��uhW	]�b���%�45��0�1�h{���xJp�5cX�V��!��sѳ
B�%L�ьk���۔Vv�"�v������R�ѽ�\�s����Y���s)D��U�[ə۩�U>��t�X��2���GkHg�m�-WU�ٚEqF��SB�>p���ĳ�E�|�wA��^YST�����.�ڱ��QF�R�g��؊�w���SU0�V�鋳�j��h���f���I�5��TS���#,v��-cvՃ���4�NE;5��Wλ)��6�'����=��6�7���^�����y�������!����4����v�{S)�h|����ǧ�Y�l�3;i���n�ܺ
p��n���j��!�
�o?��~5�,=��nG�җ��svf�n��z.,(�;�2��\�mtO�F݊��u�˃�ol��t5�p���[��������4���!|�Aj�^�ӭI�􉢤�N�nre�̼F��,��[�ݩ\�I[��%<�r�����0<�s��%[Ԅ���B�q���P�SQW��)eFs�W7c�!D	�>#6�dOZ��f�wC�qV�>�i���O+�P�MFzu;ӏi��Fcν\�G*`-u8�Jg�X!&Ġ�]���]�0���ޅG�\BH�Ҡ��|	�%z��/UV��\���,NH�M�Re`��������sT�R/0G��|�u�c�gD�_*r�xYn�����\$�Nو���>���{�ږ6���0��s{�WbUu�sn75.\XJ�d=0�;�D�����SW�^^����>�������l&hg.�6	�R�RD�T��/W����O�O��V���i����ڙ��r�W���`m�#��Q��M��>�ji�\.�}֚�x�B�S���޹)h�wݗ[V��:J�F��Wm�KfWT�9��7{e١��:E3sN���.=�����3��GDb�X�&�|�n��/�9_=��Fo۴��-�8�i��Η;oqhT.Ю�+��H��(���^MZ����wsZ]��\���ʄ�(H/O����kUD|�K��{�4�;���q���!��8��D�5��۬�؀��r�/{��f�5���"�T��nD�^씦P^�=�n#�L���N���Oo��ڹ@��7���ݭȡT�rn̦+I�͵���6�,�dRlQ^[�!�^<��[eY�l��͓˅�e��='��6*S�[NWh꛸3y���7y����'�7�+���C{�1���I��o*p��)��;p�5mNS���tMС�[��u*�͋��e�6�_]h�z�h���{����	�
1ki�Jh�L]�ʗ�@�ByM�1J�c+{��fu���H(t�]6�s�����Ջ{���]ʹs��s�:�w���<j/yjY|�6�DZ�%p[�='r�;�M
�"{��v�1�[ީ�K���\`���Em�u`�E�=ջ�u�SUyN�eb`�7�z�R�q��Y��,n���bЩ����za
v�o5X��gѳ��ut&s6;Es���`�г}�g���z銮�͝��_��>�rgֶZ����<6���挂��u�w.���O�O'�#^��+/τ��#z2�΢)�_%A��b�4o�<�O�����vG��`��@��n�;g�=Mm���;��T��Xm��W6�Y�����n�pRA;���)}5�ͼ���l�|�:��܉�ũ�=3�e�V{�r����/�id�����0���%Z{�Мy�5?R
�=�8�n�;WS��I�/C}�&ދ�7GI+��e ��Q�y�ٵFx_�H�.0+�Vc���N�.���7�f}Jh��W])�[KF_
Ɏ3�Eo��F)�mh����g8�E.�h��u\x�
.)ZU��&&�#E�۔�[j���W���K�C%擯]��x;�,pl&��ax�"u�[���T��Yݼ���T���h�x=c�ka��\Z9W]�ܤ����;h���z�#)�C���%4WfU�l����fu�iT�>A�V�*���n�x��nu1c0��`w��g�_�>�PY8��}���.��Fs^�
�P�
�a��z�T�u��nć�ԴQ7mNIy��*�-�l5���P�/Z�K��o��*��PYb�Gԋ�z�gr��֏�[��5��eG��p����a�#�f�M�Mh̩v%��e�v�;��5������b1�g�*��u�E�S��MX�:i�e���.�c唛���h�ɷηX��t�ޏ}��Ѝ[�(���mM�������γw/�:��vR]@ut��.���r�=�����x8�.-0�6��{H�we�����Cz�M�X�)W�С��4H�7�Vɕ�
�<�-90��sR\���^L�m����: f�e��]vI��|�^em:�
�h[�CPCa�5=:����BY�sV.қ���[�����1�6(%��R�L�*)5��ʡ��xY49���_l�����ż���>���ڬ�M��[���4�\��0�w˒�
��e��u�t�4m�r�Yn�P>����]Ϝ��%��9�-�jϯ��}�r��y[��3%=`y��5�S���kSV�k�ǁ�a36�R�'Zn�T�DO��Ձ"���m�c�L�)r\m�ǽ7����r7~�4s�'�	��e���7wI�(=�y�q.7�!�F��])�+��{yQX��N��	�>�{1�>՝)̼�b�cWҥp\R�eN-��9+TǗ_>�Nb���Z�g�^$��k����+��!x��4���WE�t��\�9�o�>�G�-�;�t 뛼�(�t<p�ʋ@���H��^Mis�˽�oP���V���Au"9T�B���˕a�m��Rf�7S����j{�#�����r�]H��ĺ���^�]�����/��)t��E�u��:1�@���*�t%c̢̻J�&G^�m�(�����ӄ}\dQ��*n>&��C�y9ф�8�U����&���N�C���8-���LȧnS���**ȱ�f���F��E�fW>��^�U��c`��es�ܡkc줶��,�gϊJ�MX�������>A�����HO&u
�pE��]�]��BMl_%�򤷇�c�"��3;Xe�EN�V��K����\5��v�R]��*�l����r�W1Z/�#��f�҉Wd��y������i;ڕ�Cس�Mq��Zj��:l*ͳV���PȖ�61�u�K>ㅮ6��*�t/3����]C@6;$U��ݢ,k�m�����	���������rwYA��D1"��v�����779��	$��������O-WG^�9�jM4����F��T�*��i�����dJ�4�߂�ǧ`�H{����b��ʹ��@<Ep�o��K�W�uҤ�&(CY+��^Uej.5gKhmf��wc|�gF݉:k�MqW0�5��]fV`c�uc��3�b��dΫ̡��ɞ�s�7Y�V���w��՚�)�ƪ��j�hmb�ww�.��7�X�3C��Y�
�j+�/�`��{��%J�g�9y�9�oB��6Y9���>���M��|;;k����^p���K�Q��'wF���/aj&u��E�Ō˗��7"�1C��ocw�e.�|�n)\0QM!͝�"vë�R�G[EL�T��0���:���;7[5k�*ՂT���؜0�Y��R&����F��|�-�	ls-_r�=UxwALo�l�8���+�ۛ�Ԯ��듨hW@V��)�WoN���7ED,�#�����P���v�6��m*o_'n���\ѷ 
oN�樖��ua�}s���c�qZ;w؅q��o���Xݓ{:]r�ڐ�".,|��;�>Bh��NN�&�b���R��$�x8������oVinXOD��e�j�����*f�x"S�������g�Ut�[����C���;2��t8�
�G�R�������pc�����0�=&��˦���)�h�^�O 7
[(�[�W=G��������:7�t�3���Nk7�q�īE��]�uڸ�dy9�o���s:z�b�-���T����"�'I��Tb���$��Y+&2�Z(�Zڕ!�P�E���
�����E�"�R)+1�%�B�J��U���(
���PF
E�X�eJ�
�0PP
��j�*,oY�)U1����WI)R#m"�x���
Z�����Q�F�Z�E+1�k����6�T)�@��Y�֊� [T%d�RU-*��R-�a\J�(T%k�VkXa4���"�m%TR6�kR��\��QDX
VTX

�%J� �@�E�X,��b*�h�)�J+&�������*���J�*$�X�X�f��=�<{�F����+ܺ������'�0��řI�s�jl+�0&{)p�P����˔)�o�Ns��ڥg|mB[��I��A�����w��Y�?j|�L�1�����h�zL��!��D��7ˑ1a�ݔ��;7��4���U�[��j�F^�����J�1Ǻ��"g�4m��fM+��^nk{�ɩ�PR5n�DH]�pGۈɮ���c)��﷑��w������C�M.���+�_�ke�ۥk��;��}X�n��9/Jj��u�֔)\`�E�^L�Z:�>��������>{��v�����|���62KCD:�{ԯU�=�:źlPݧ0�YhV����!I��;��6-���n��*-�}��uy��v���!hm׉������e�t�%�!��nM|�e�as)%��8���sy�";�I�v����L\#/�igN5x6���j�dCĸ�w��	*g�Y��`���h<�q����l���Kvz���E�M%�g8��}�R�Z�)�\pS�������[��$��oz�vٯ&�ˤ�ݫ��2��<�0��#v4��뗇�ȁK����=o�c�;�=b�t�264�kb;�\�h����O&t߰�rz]�z��pP��f�.���w��{}HmZ��:��{G��M�I)����+�
P|�g�l���!�+��v��~�]\�bܼ|��\�Rn�peGb��B�*l��[����a5]3�plZi��dq�T�mV�1m�<��y\��f���{D�Ʊ<�]p4B
D�eNy%�5dcņMe��Q�vZUo��t����4v�6��R��L	�3-2I#��([��8O1/�DF��4%um���CE�Yv�l��2�ud�ޱĊrU�l�793�����wW�nS�eu!yd�S*Nȣ��#�2�R�L]ı�net�J��y0]7�����>����ٞ�cA��ӂs*��7���[^�ڣ0��]���u�)=���s�~��\��K���=�AW��хE齥���O:ы��Z��6S�{iGFԣAm$�iن�/?v��'�a��׹\5M
[آ������u���Ü�xB4+��<���I�gM�U�R>�n��W3\{'���1��+�@�H/we�Gݖ�՛�����U��ا��QвoX��[@����C.�tU��vJia�=O���~EDNq#4���];���Y��uvإ;K\�P�4���!��_O�]�*��to�-��7�:W3�7�v+KCW\��n#�dpҥ���ɋ4h���s�;'�܀�؁pfj�#��C6�p��R�㢱�bK�f&�GL;1�`��G�N1���{osG+��#�E.�N�dKeK$��8|'��
���oNZ�>���ŉ2\
��1g ��J\�����2�R���&D����l��9B�P����>*'�W3ҫ��ʫ�x:�9�j�ٶ��<�=/�L�3\Ȧ��t��^��[U��TL7<6L!�ݻiEXW{ܓ�1��_������؈n�iҬ9��Dg>q�����e�
��Z��!܇);)I�GḾ�F� �����Mu�3�Z��^��t�<!�!��5B�IRiuH�yh�f�U��U־n����7S]`s�U�^�ugq�>���J���@:}�`��Mv�uh�$ܲi	�Qu
�痆�_yZ��֜�מ]�]-���}��ԁ�꾿�T�؀��`�p�\�EO9ܐ3קܘ�]�*�~&�PW�NcPv�ʺ����2��h[3�y��w,�6·�t�� vs���x��w���̈́��X��4�]N���!�:p���3��qE��j��M��=�b���dYk���n\��ؐ��ˮՀ��x����t:���|tH(LWp[��	�\��$P�yMgي���J�l<3�<��F���s�H�$�^������8�c]x�h�~�V�R*�
�p���WGox��4-�cW�;d�f��|�?p�\FE��0�\h�	�G�=n��$��~���E4o�Г�8{�,�W���<*�4O9���lq��]yW��=�
^1+틧��ba��w�~�� �3�(x��Oǅ��[r=�Ze����e�>���v :�Sb�q4
�9>�3H� ��\8*y7��c���9R֧����P$xC��(5�CT�5�u�2\.�� ��f���n�s��{&�N� ��DG�.3 ��,s8���cC<�����v�T�~9!�dӖ,q
�s⥩��T�"=�(yYV�/�����m]�ZP���G���Y�pH�&t2h,���e�:S@�]�驟�e�l蠪ݜ�m圷�Wc5��&XۆD �)�}��l:Rj���V��9c��6��q�Kie��B�0�B��B�*.7)��������֨T	R���91ռ-���SUt��׊���IH�����N%�.Z�q[�Α�zu9�F��[Q"�N�qp�K�|��ri�T�W�P����<s�΂���z�+0��M�!E�9��NDZ���ᆘ���8Uz�w^�ډHi�oi'y�>�ޗ�ӱ�.:(t��^�V�l�t)��1�W�sR�97ЭV�)���"�q;5��^�!t��Q]}5�)Tt�Y��^H���V4�:B��'���т:4��[:1�*�:�S�[����a={��^����=GhSg�`�+�^��j�˅��u�/��6�MVY��a�����̹��|�h5	���IXx�p�V��ln�60���ޟw�aZi��|t�+͊�1��t�zC�OCqo:"f�ؗ�\��D`���( na���p<��w�[ƶ���ݗ�d���|�[�#%�C�����ީ�)���H��Q��x�m���ʹ�u˷+���Í�ǻ#Y���p�gw.�~R╪�"Br�~H�wD8Q�Q�!o��'F,�ӗ}x�£b���{�>70��P'K���5A�p(��!�^�J�w�t�&��;��[�[1�sz��磣�\LWgD��2��;޾u=��G�5��T����|�O�^�<�|���=�[7�ג��,!�z�_ْV�|º0}�UJ�B�nr&8F��������Z�q�r�E{\&�k���@H~߉�4!��J+*�=��7����ُFP���:��<5���:����!�x�H�g MXC�InP�ĻyogX���J�!�����_��|��Zxf��]lb�P|*����ʟ�Z�Х����lU϶5C�%;�z��H�����X�
	ձ�_<ʕ@����LP��QJv:�(�z����D��0� KҠQ���Dx�7��Gp��Z;����MJ�ޱ�^!��ܸyr��npu�ҴBոz��N5���g2�M�t����چ�&�uy�U�w��9�7-�3��Y����M�P���k�^��U��e^�Haqg�Dh�: L�!��lPO��>PG�F|�eoV��T�\~g�������{��JB��7�l�6��~������&4��z�gcX��ڦ��L�['��Q9>�1��5� 뼂���o�h�׮'$L(Ψ"4ڟS%��a�(��C���q�k�ԏ*�����tG8z�_.\��h21��)�#<�8bz/���
�Q��^��1��rO��
�Q�,΋������D�:�2�UV�vi�a����{��@��s�!�Q�=<�zbx��^j� W��y'�7� �jk4�#4��>蜑�5 �j��T���网��ލ܌o�<51��|~����C}��a����?^Yj�U�4�5w�!�E�P�U��P�~q��!V� ���M���2+I=\V`� �/^%zgkC����5�f�P�d7ʮ,�s/h#Sqշǆ�t���Ol?i��G����L�wb��>3�ZSЛz��ɒ[y��p��u[����gY��|�u��ڇ��>�=�iʗI{=V����To��A�U�p}���9鸬[y��tD�G��z�:��*���9g!)ƕ^����	�Qn�z�4o=�����Iو��Qp����p�쵗/`wZ��ot� +����~[�W���Syx�<>��[�(J����g��H��u-0������y4vNF�q�q�؞P}�}�;V"��L��DH�]�X����88���*yd����4r8 �w��s��Z�_�!U٭��̪N9��Ǌ�h��x�sNGA�]"ԕ:�J�Ѓ* GCy빙���o�RF�dϱ�#"A�:(*t(��qu!9��i�M�D�������ڹ�膻�E�i|l��uծf�:\���cqU�3�{�b�T`T=���)�>}O�̢hx��Oǅ��Z�:�x�Uy���Z�u�M�(�UϞg���rs.C7\N�^R�gK�`�W�Ve��\����A=K(�S��IH���ꕑWv�z��j��c4Fs�����֎��Gl���zU#,�tS-�����L����
e��E�׊�9>��9`W@�]-��7�<���'���.p����Gpᾃ�h��$8ӄt�\�uo��7������b�$Z���L!B@s��t�4�#��W����h;n'�Z��'�`���"⹟���r��
�s⥩�����F7k7�N�����r.+,U�*.3)P�q��no� �j��c'91ջ��ޅr��S4��L��H3qJ�W�n���\8�>�|��槮�S�F�/��p�O���>� n͹��
�.O��P��Y�u)[�P���u.{c��I�u�?1]f�kk�e�.�ze��������ڨ^��=�c^b�q�t1|cg�.Z��+NF�����#�d�t)
��^�qV	�s�Z�P�`��];(&~�~�ʷ��c����y��!����Z���$!$�4���$�$���'�$!$��?�`��~���%��93��5��o�����8�עz�%�q?�D4�&���r�$@  pǷ�!`�B��#�B�i���Y��2�*@�8%݇���,��$���E��2?-�Y�?��?���0;� ����������}z�� ��g��t�s�e���0�R����oRu�
����Ǿ��� $$����������y�$�I�� ?$�	C��'p���C��~���ɇ����a�C����O��pa�_����Y�'����F��	!	$;�!�������"$��	���$9��Js���=�8���?�ÃB��ZY�����?$>p�b)���'��Ne1'�x(II ��#��c<ˁ_�� 	��$�>�	_��2y*�;��aC����`q��n�����?����HBI���r"����C��O�O������z	�?3�������O!�}�!�"l�CRO��f��?#�I)������9�|>�2�$!$��,���>�������w���p��S���9�S	�BΤ��/���'?g�t^!����O�|����3�$��?�>��~���~2�C�O�dc����Qg���>C����0D��P=��������!$��A���	!	$?��O� Jz'��ɢ�Y�ק�Jw��vp|�$�ȇ'�$!!$�!�LD$��0~���;'�/RI$$����d�����C�>��N	����D9�Ԕ�P'=��$�g�&0����8���Ƚ���BHx������T��!!	$��'��!�ȓ�?�����������z���>�0~?�>�>��?R!��>��a������9���_���d$!$��~S����?I$���Y$�?�C�?�BO��d�ې������Mx�������w�'�	�ć����\��3�#2	�?-�Hc�P�O�����䟗���C���g�?��/��3��D��5�W���s��II!������ss��y���|oݣ�v'��(� �|~���a��)�����8!�%�!װ�� ��C�!O�d�	�} v���?I�C�<�G?0BI��Y����A�C��i9�qe$�08�?f@��89!��A}���,!�����N����H�

��{�