BZh91AY&SY��G��8߀@q���#� ����bA�}T    w��M�R�l�(c��d
2m���J�MhiD[Z�[m�dU@���[m�4�j���m�V��lƚ�����l��m���,�ֶ�6�d���55�I��Ь�ѣ ��1V�͒Ц�T��ĲԭP��(�`�-�m�A��l��[
,�"�Zh>M٫l��I�a�f*�*j�
�dVU-+[[3jJ��I�M[b�Z��k[6�f­���F)m-e�Vl�5�YL����Yj����Qs�V[KU�ٷ�  �kW��9�V��m�̦UJ��wZ����vwv�)Cu��+U)4�k����uv��f�;�ZQJ��v�E������Vڶjl�K�  w���6��P��m� ݫ�  q�t�hgU` ���  ��  :p hh;��
 ]�Z�m��Z�0�m��6l���x   ^ � <f �3��z Fx� z��x{� �/r�/@��/<� 9�^x  �{�x� u�s�x@7;�I��@��U�²�Z���  ]g�P�{ s���Р�=���  n����{aAF�����t��m�碀 s����:� Ѻu�� ��廧@i�=�^�j�Ҧh�e�3��.   Z�� ]� : h��:�:7v� J�� t�'  �-�� ��k[�:� GvpN���&@;c�w��M�miVQ�a��ڵ#� �� 9t�U�  :��:��J�
 �w- �� hP�� �; h � i�3r���^����j��Ҷ��)Z�A��  ��@ �j] ]�8]�ks@ 9v�  7R�  v�\�r�v�V�Z v�P�tz+hJ���ʚf�� ����aT*��� D��  �u�@�p� ;�� k�tW7N 
A�z�kUl%�M��456��� u�Pk�  m�� us�� �����sn  f;�� v�q�R�X wv�@(w6��Ck#fT-���#� � h��� +������8P�9�q� ;�� 3v�ҀQ��ꪠ�� 7k����     ��R�       ��i�R��   �O��JUS�@      ���R� � h   "�d�RzM#A	� d�#�4z�%)1�I*&����424��4��8�yR��T��s�	�+Z�'�n�����+l%ka��T�p_RԋJu� ��R����� 
���� *��L�S�r>�S����y����@Y��U_���J �����%O� Z�<�|�ޏc �l(maC��J0'�Y�"���<e�2�XS���ȝd8���zʝaN����YS�)�*u�=��Y�#�C��� ��:�=d�/YG�+�Ra�X���
u�z�=d>�YG���Q�(��z�=`�X_l'YS���*~2�YS���'XS����*u�z�=aO�)�@�:aN�'Y���� ��:ȝd:�̩�T�
u�:��aN�'Y����:��:��`N��YS����*u�����:�<`N�'XS���D�"u�:��x�d������D�(u�:�dN�'X��0�`LʝaN�XS����"u�:��d:aN2/X���T�*u�z�=`�/�W� u�x��d�/Y��W�:ʽe^��YD�{e�XC��q�Q���G������AG0�=dEz���A� #�E���Y ��X<a@:� � W� �X��=dU:�*u�T���D�*�2��̀YP��=dz���Q���QG���X <`z���aE}�
>�D_l���"���*��S0�X��=`W���T�"u�:ʞ0�Yz�N�'Y�)��"u�za^�p�=dN�X����u�:�}`z�=`N2YC�	�T� ��:ȝa����:���?���ݸ��S�$6s�J���i�S��g��Y��:��wԈ��v�S�g
xcv�_��F���S@���>Y�k�-�[@&�rz��Wj����K�2G>X7�W�%��Lb^�ǈ�$ݙ��դ���K\����V0(r��8����q���]3j\?h� �ui��S�ded7p')�H Q��e 4��%�e��,�&���*^������6�"F��6� �H��m��T"�m���1�S���x5ޡQf�nK{���)��#t%���\�
��2�:��n�����̄�B�Loۨ�U�e�,�z���e�����
9mn���8@@4ӫ�I�-��J=ǖl���"��j�-���a&a�:t�m�rC�n�����Nԓ�Pb��he�ɉ��e?�I�a=��m��,ٴ�E;L�w,ko�n�Ѩ�f��QlT�ḙ��ȍZn�xÑ^������%jK4bڷ�E�- ��"!ђd��8����]�)@���MM�A6S���	l�b6�˖�9H��6�ѳH̟�Ѻu�V�m�Ә,7��$��Ҫ��8"�]մ�G]E�oVPr!�7"e��;�$�Y��8� 9�mdsOr�K��L|�,�f,-4�n3.!��:%dh��6��IGY���˕�	�ف����jۼ�z�M!fks&8@�ә-J6��ӻ����
�f�Hܘ�b�0P��Zu2��%��5s�6��mG�	u,�z�B�1/�8^�o8lޣ���[�vh�U�w�OI�g:���i�����Z����k(�dD��kWH�ܙc������T")�:k0�,���=� oLƲ���%;�j������b��nP��DMVL{���s��݃w#��w����
l1쨭�HW�H�r�tQU��M�t.�ݳ�hQ5ӾLNy�#�;4�`�� &�ղ6������Vr�c�/6��K"��c��K]�7Z��zi�ڹ�ڲk]jOyX�ҫKկN� ]y�m�<�5e���3H[	J�DR�כ�7RA]�e�ӝ�2�y�Rl���Yg亵L��'E��v�S4ު2V���	�4�x�<�� �],�pQ�l�����.�f��͏-\5�nV2�u)Ø���6e#�]���s4�ְ�Q��S.P�fn��<,| 3WϪ�dP�h��&qX��ݼ��m�ߒw3*7\N"�j��&4��Ѷ��zTנm���T�91�[����j[#���2 �&�a��tRvjB�Xi�	���b�Դ�F��A�� 2�C�Yl-���^ p��C��4��7j����X)�i�Sc�b0��n,�Qܙbՠe��n�����@�<�t:�������O�z:�ҨK5u��{��Ĳ���V�#�%�T�iŴE���+,<Z-`�6����{!-=��7^�Ϸқ�j���@X��s]�c#����8[H�e�6å)h��V��rӚ�smI�C!�n�^�z���S�-����d��֦䫚�/,VA̛���A�ke%�|�1%����l�V�B2�X�1]�hY�0��g�2��r���P�CpU�(Gz�a��m	�/k&�X�[�����$
*i&�z��t��Y�Gi���pPy`���
ǂ�n��'�[� �Hnj���c:�gVU���H��^͢46����^��3�yQL���n^3,֪��F��C�$��^�*�[�/ZA�{�Ym&ﳘ���¯�oiAm]��.Jִқ)�י)�]+į aa��&��A!��PeKy���N-lc�b\n�m����Tk
����`���:>ԛevR`���nr��q2.�V-6y�B|XZ��O�M�@e��ՁM�E���X�j� �̫�̘M����@���֛]Z���sm�r[N�i�,�%���ĩ/m����d���@,i�[�j�nU���A%u���a�Ș��w :^��Jb�<��б�u]���	{,T�Z&-{)�G��_j	��6��%�����M�-/�0Ôr�hK8�!�m�P8�-yM��H���0�k�����He1�lYN�Õykm¯�e������2��6��Jˊ��JO�r�J��w,Zcc6�G�\ܥ����R6��+/	��%,E�r���<�>dϠ�w�;���*�1Zc��{��	���6���6005(G%e�P6�f��[�h�զ��u�GԦ⥬J�S��VY�ḛ��L=2�ԬӆIl�)���dm1.�"�x���2�0��+sr�E���I�0�աP���Z�N4�Q:���L�B��6ej�fܭ�%��{a^����,f��ˢ�
�W������=ю��6S�Z�Ō)Kа�Wx[
�C�U��h��˗'F�2��w�8rـ��%Q��V��ٹ��d�󼯘* ��͑�U�^z���[����v4��ʹ@���}��/F��ݠlL��a���0�v��6�,������G�[``�Q�̼g#�9x�6n�f�y���R�*� ����s[͡�f�S����vYy�Ap �uPʛ�˭�s2�8��v@�Eع�78K�PK��r,WEZ�+���:�!����jmnO(�k���q�j*5���e�Hf]\J�0���n57-�c(��SWW7x��;T�lg*�t�I��!b�#2�ޘ܅�p�Pd:���ͨd ���l(mM�O2�]f��3ifh����F9R�A��N��NI#R���	`H���۫5�2����J��)l+�h�tuт�p!@]3Kv�X�^K501N9����i�n:A�A���^�2� ��r�gko&I�u�x��֞tPE|�f7���vv#J��gs�n���Dʃt8
l[wkN
\m����.m3��ݽ�p6��	�S�n6�{>ǋXӪG���� �l'\���]_u$;p�i��ia:�">y��a�;�v
�R��f�e�˱�������ῲ���ŭ��YyB�*�`�����Dj5	U��O5^�LI�pK�@�f�Ph֑�6��t�c\#p6%<�"�-�I�rdx!Ňr&�Gk-�"A�7�͹�	S[É��o �
zl��6�#l�k�g1��$�X�=�X�Pd��5��i�EF�W ��Y�j�-�-;3f\�ӂ�2��u&�q�*�!��1�t�n�X���9�����i]e�tv[4le)%Ѵ1�Ll�1Y�v��SB
n뫭bъ�^����$���:2VJ3V1����"�֩����H���\��*�{YJT��ZD�3jmS��|���suj��î�	����^MB�`���<p?�x!y�h���y1�$��S�,�!�֍��������
ky���f��BX�](�h{�2|wviE�KmX���(֌��0���m�qU�.�A��٠V���\���Ď�ڵ� (����R��ܬ�l�Zi�a*
��al�BB�0c���˗n�%[�QT.� �RP��B�t�ˢ0S�&��
�c�ڟ�*]��Ӥ
J�f���J��_*E�Moj�9Oa���A�0To%������mM�Mk����z��F-���y�a��� �4��ЃwMn�{�`7X��0��S�W���6������]` yD�8��@�#����׬V֜��d�{ÔJ��6�f�f1-��N�j��ͭ�uW4wBېb����6�t(�m�r�]����P�Xz���X�����dV"�
U�Z�%����f���@җ�HP�PIj��MB�*5���R�K�L˄ �z�xN� �$<̳J�O7c{1'SS�aS�%j�n-vЗ��n��4M\ڃ��gN��#n��t�����y���T!���vb��ЋS-[RR���ݶ�,jS�&��no�Le��@��f�#7o��:pif�s@��U��MH���F�M��.�w&������W-�-�i�����a�clBހ�������Ɍdb*10r��K`ô�j����FMz4��#F��)��ХE���� �R�� G�{KR���E��ql����nźr��Y�����qU�)�8\*:�jT��S�CwGi*�/FR�/��?��BE�R�o���ʱ�r�q�ȸD�^��3T����(#U�1�o&���S�ii#3+u���.��k���5o�.b^��fn��]�tZ)K�	���=T�lsK��t��`��U�uP�^��dVe\Df2�;p r��?=ڃFJB�`x�;L�<��csRpI���ۭó(aa�wY��-�(kE�K+u�����=ɨ��T�JZ�h6��Q8�$�^("B��4c�ӳsU�4��b��N�o�����n�����@̻,�
 �n�B],�N*zou��k4�j�8�9��i����Q�݁GJ����9�yyw.��(�:h���϶$�/6�Abf�*�!�ȑ��H�Db1:��V�]����!����U�؄,)e8ɀ��E����^�x˷x��F�lV�7���+��	����,��k��4��Xo`��U��ÙZ�G$�%ҭ@��.��CUmb��'����g�t9dq�n�����n�D=�h�/B�/2���a�Yt�l:&�h�y�
]��N�g9���;��M20�R�uB��n��+1�̑�#M���� �nI������3��M`76�4��z��@��9r[���l�����]�M�7ii�B�kOۘ��Ǘj��6���O)��F����N��!*ɃFZ��IM��g��l�H�,�n�Çj�4�{z\ʏ-����c��Eģ3H�,�n�vLr�m�w��:�ii�7dm�gh%���+6�CCfȁ���Ӗ)�г"͕q��2����'{���wm�#���q���eL9)��M*P�Un�*I�����N]�GMD�����m���BNP�-���D�BD4��3�T�cs&�O7M^�9�)�W2�ZbӦ��;��fSyw��a]�M�FY�km<���@�k����\�.m*�5:�>�v��Lv�Î� �iZ�b�v��᝜��,X��W&�&&��T'� #��Ja�=��&�D��[4�A���H�f���K,�VP�����j��[�ƉP�iM�A�5���0�F�����Vi*ɹ�4�0^��z�8�n�pJ.�CJ�bĚm&�ݥfC0�j���2jcCC%fѦ(�Ɩک7
��Q43F�ȥhnf�.ZZpu��5���|����jͭ��͛KR��UL��v�Ä	v-�#���ߣT���e5q�� 5�L;��+�1kP�Zz�o�coQ���,�ekKUKߋY0�-��1��JŅLia�W{����hx��P� ��I��+�̌m�
��d�ynjl��r�f�.�ޓF8	a|�n0��(Si6c��k2蜈cTg�
�����q�[�A��-��Xgo]T&�r7w�M�M��u܊1�qR�r�ڙŖ͍z����óK.���uޚĦ�.�kt�ք%��K)���%[�5�x^L��Eŷ�\M`���h����ۏc�dV���5�v�έj��61�[��aG+ ,���n���HC1hBe*�L4}�f�gU���!����׹J�TG���d���c��^��a�[S�{!-��"� �E�vc�kF�r�6f��=�2E�Rؤsl;�Q�R`W�Y��{f���KͳkL�Ʀ�:ך��x&���;fRڶu]f;Ln�ѱ ���b�
�|2�C��h�L�?6E��t.�U�e�V�z��w���1-kt��J�=�<ѣ3K��U��C�O(#kI�hfL�܎M�B��D,�2F���ll�h��i���3~47��Y�p����ۍ���iM[��4�hn�z���x�$X�Ź�nu �h)#����ݣ���n��o+w.gJAV�n2Sܘ4m�ǩe�:�	�{-�!���fMM� ����q��� ���G
���em�oX(�~-��y[��.�y�lzټ �Ww���QH�э�e��7`*}5M��0^ɸ��2�à��Rh�a�d.�D桁;���wY���S	h���U�zd/�0Z�5�g������D�Ҷ�la֎�a�x��Q����`#p���[� f��A�(�J�Ǻ4����R�@�w%t��0J�'�Ի���ERabЪ뫗st&8�n��hl�*�*���T���4d��̵�v�b��=�P�u��@i����L)lp�YF����IE��{�sy�m={E`�sCb֬��C؆:+0�%�\��&�c�\��O�Я*\� ^d�iJ����*����ְ�����Z+[����,ދ�X�(Z�1=���L��n,X1��#�6��&a�V�+l�Y.�h��ݵ*��j	��Q��ݩ{��1���ci�͸�sk�򽷡b�h�HR��T̹v�K��+0��4�E:K�V�wa�L<ڻ���8������A�$
`9Gt��Ҽ14����jK��ϫ�ے�?�Gx��֑;�]Jv̆U�IK��yɓ���+l\�uf�wpIa���:�Za��A�"w|atr��\���+�|X�o�`�����#֝L���;�#��Y���@�hwt�K]A�"�3�c�V��L�0��)�1�#{�钟iu�g\��ww���H-g)��p�m˘���s���b}��ܫaX��Q#�S���)8���L�Go2tw����L��q�Z
�&P]-�!j.	^b����Af��eIОF���_(ü�:�`]�΀޺�H���-"��15�oN�̷��	�z�Z	B'S�Vl����]�c���Bt�D�mK �y�u���a�kwnx�׼�������j�o/��~Ia����]���W���rM�+s�rJ�'&��Rr�^�ѕ*V���$��M�/�vԋ&KR=Ft��ˤj؜��{�靑��3\�����t�u�>���Ρbܵ1����&4���Q��{v�O��8��ꅵ��]�	L@5�3�`+�չ��D�$�L7�N66�g'«^^'��7�x;�]Q�5�b��	l�{�ً��KN�s�T�õ�%��0Ťd�΄p�*�A�AM����y�&<�]�y�S��Π�?�j���^�r�0r��d*�_q������ {mM�ّ��N|i���%���+5��um���]�AN
�1*���'��eH��R��t��}�9a���Ѳ�C�mA��e^�8l�Oa�˒Z��TC�
��&p]�xi��e��!3�����e�[�����Kø3.�����t<�q�ocB�$T��o�ݐ�	����i�f�k��d���j����uǘ#�hznpC����)���l6��k�	rڵ�r�흰⫛�|�w�H������5�Tf-�m^�AD�������l��;���V�*�����c�ZhEl�:�U��N�	�v��#/Eu��=��@��[o��8�ry���9�e�޺s����j�{�K���ӵ%��u9�/�v��)^��t��k	�Д�[�8k�����>{oX��ؽ�2`���>Z�
Qw�/D�a�����7A�f��鳔��Ę\#��Jn��h
����p͹]���r�jė.B^�8��{��/����N�lwV��,�5��5f��&"P���VV#Bw"�Ïs*9 �ʷ�]�m)��AM�
��N���W�18S/5���.�g{5<w�����+�
�t�
gi�5�7�����5ua���͉��V�Q�wcś�r����-������p�ܳ�\' �۽~O��Z����L��&�r�U�0�Y;\��
U!|����]�^ʼۣ�m��O�k�T�c�P3��Z:2��NH��gU�j��J��\�:���2f�s0Ͱ�sZӿeڽ�T:3D�v^�j�33R��H��"2Q�n�2�ʸ3��F��{p����1�S��࠺�k��{�Bk�>PY�z��Wp�Sb����˯ɰ��b�����X�R�"_T��ޚ�B��8.�]gr���=�e�n�a��+����=�����Er-��KۑbS�-��ck@�:m�S�>��,�-���&qkϡSr��Υ;A"����V[J\�Og%��C���z�v7�F��υ���/7�=1'(�u ��E�/^��˸b��j���+�mX�o�
㊋I6��o.�47+��km��� 
�h�s�����`���z�u���e��Y�zgqn!c3���s�jń������vб�3�e�_'�a�l>yF���f���7X�7�M]Շ�P�v5�Fa����p[�<C�<E �1к�={�)�\��TQ��K{9i��{t�NVUɂi��2�0�mvը�i����YX���:�M�!T�k���j�m�����,�!
�&�n_)�g��N����\�7h �'L��T��g�omsVN1���x�Fŵ���e��t�f#�#�f�`-��IK��x����-%y �nts�lӄ*���R+��Xʡ�~ۘ�(��P�[ү�Ac׈�bX���C�m��=P�|�bW9Q<�$����fQ�=���1�ܔ%щ��:�8��^]ſ_G��G�㒂v��ݾ�MP��v-�i%��uV��֔!��.����H�w��6ŔrE,�7Rvt�ǯ����C��χ���2��j/�c+��-�'�/(3�ŀ�QnP����:�46�Cu��% �>�KC�׶�c4ӽN���Ʈ�TE��e�H�d�����4�=D��ޢt��Q8K�B_u��O���3�ꊻ��5����ijˇ�X�:t<�{�mO�6_��E��o��5x{��%\i�se�WZ�w�UqN-n��p�0��Ō�[N�(��մgvVu�n��#�2��d��"��LԺ�C.�Zy�9k�#�K�hh"s"_�·��Y%����;�ü�V|���R����j�}3����[�Ӻ��Vb
���D�&2��"}\���u�cR��}���S����;���A�s1)��*բ�嘴Z��L�E�e�D @�i�¥���\��QN��)]��E���à��J�z�X��g���쇩T�`��M�#�}.��I�ͷ8!9g]!��)�!��K��Lj�o$�w��+kX�ɶMJ�6�+�̽�+vM��!�R��W\�1����/�E�X�>�����E o�l`]��Pͭ=�1뮾���n�;����.|3/u����M󊖀���-��R�E�O�����Se�F@:������"m���J����bUr��Y�dӈ�cME�k�LP�~��p�jʾ��νhd��ұخ�0ӟm�j��L��8s�]��;����PT��7CP���*�}8��MN�]f6:%��b|��:��k-�!>��V�[�[(VW*@��gk�t �r<�b�����]}GRU� b�-;���^(�K�-w���zo�3H�M�.��V-����c�.ݢ������m*�A�D�J\��*�Ӯ�V�ǆ�1;�fя/�/"y�V���`�����7��]�6����l:�7q�A�x��n��]nbAs�+*��e��hb !�����7�1��<�2i���'���N�F�t�jd��3r#j:͛�v�KVõ�/��ƥ�a��
�$'���$�,V�s �K5Na�Q*h�C�w�S.��
iY)��s/C+3m�pf�Eӌ��G7kyu���j�j��$��.�[0Zz�ig4��pf��:&���D���Ӭ:}s ɵ�����H�Z��*I{��rۮG����Ӊn��!��$n���؍�h�B�2����.�e�{��C�E���l��5fV��ܹ®��B|�7��6>U���=��[�I���/����ou��P^�6��38��]�C6����kHy�7O;�S�]rC�'hY�X�x>����:�.��F�z�'c�❥^���;���e���ݻ��7��Yڦ��]��6Q�@Į�`R��l���*@:�N�S=פ'�&`Ǿ	}�7\���k	�
ϳ�T��]�G9Ig|�;պ���T�m�pi}��zB���A�}H��N�nlU(hB�y���}Z���]e:Z�K�i�K�*R�Z�٨�P�ۄ֖[ݔ�k5fCx��1���3�ӭ�XݫL�{l�f�*}�Vu�M��^�V^L3�B%��\=9�3�,�b��X��U0��zd�	S; P�v26��9MM5ܹ���N��R;�t�ZN�8�z-��vg��C(C�@��} ��n�Z�ʋ^��}#T��=W����v�Z�b�{�i��%�6�$��m��|:��+��1v���q�wG_j���/���2)xj�{�!̧�*^�Ph�S6����ɕ�-���Ԇ�걬<�O��K1	�XJ�����m����b\5t5�k����y%���
�s����ѩ9�����a�9=�2mvf��}��gJ]��֯���p�_,�cv$j�����	�Ɣ�Ϲ�R�$K�X�5���]
��:������4�X�燲͈UD��ʙ�̈́t\l:ԩӋf��zVGF��Zr�wf�l�QSemrwz�������g��O��[�nM"S�����D!�4�ݙ�y��>�4�T��BO�0�-�E,,23��^��+ʐyWOpe�H�vڦ(� `��O3���TT
�a�Hl��Gi�(⏷�<�A�/�lJC�:.��B������(�����zt`��Nʉ�nяq>��i�&��>�JF4f!t���h�2\��{6DL<l�&����ʔ�[q|	�r�v�(�L�5���2s��k�KB�(�ga��L�p?�5ݐ��n��-R�Jl�_Vv���V�"֏�$B�H'2va|��u��`���=@qe*�U�;yk�4:�P���;/�s�_cl���ܬ�v]i$8���
�7n���� �YXn�'�w�Lꂴv��Ty%K���4�/�:WE2���1��ȴ�y�Fz�tg�6�9��c�\s���j�F٧��8qs�R��T��5˶�cr��rmIJ��cR��ʯ���۶ޠ��q�%��Rl[�+��[p���so!�s\�g����E�`�uݣy]�ʚn��ȣ/D7��n��GB�-�nhW;W%1\	8�ej�Ka�,tF�ʆ�p�fQ���l��Ű�5������p
��0�|��k/����G!Uu8�i���A�g_'V̱n�$�wu��%:4Nf[Yq�a�ϵ�c�F2TR!���7��%n���N�5.WeK��VXuF���P]���Ӣ>N�CZ1ĩ\���u����]/�t��@�G��<TT�A=N��wG6���SA�lit�yJ粔10���D`\4T�0	����W>YYq��f6g40mh��\�e��I����2�Xd�+}eQ��B�[�m������d�*�\}��^<�
:mp�W�^���6����mEj��[xW�d�#:h��� ����d�jVά��՛���I�+��K�nF+oA_Kq�N��խ�N��+��pU���
s_[6�U�����c�}�f�%���Y���7��^*q%���m*��q�qi���_I��{�u��'4�v�/w�"�^2��i_1Җ=�P������bl��� ��L�&�G�mVDk,e��'�u��bS�v����{n%C�՘�W4�y��tŰ��G�T�������z{L��s�@4���]�p
WRusFo"��oW\b�U�YCo9�����(Q�^Q	� 8�p6���R1v�Ls0�G���aJt)h0��n���.�N��`<�u�.?�|c�K*V��8o��̷������P;�0t�ϲgr����VWB��ҩ�u��f���7���8Cʒ��2��v��T�R���3rwM�;�M=�<�5�`�އ_�T� !mɍ	8YL�;{��iΚ�����Wۢ�Y[�h�Ԭ�FS��Wd�ց�`�&dհ��ڑ�΋$�&�I��L�ylP���_>Q�c��T�5�s���.�
}�,ᥪ���B���j�iF�5x�mgdw��r-���|�,s̝j����8�P�Bc`yC<62ƥ�N;����*a_	f�^u�X	q��Ԑ�M���H,C�����[ж9{�]�8���5�2�#�p��WV	ǵu`KsT!��:7�e.aۣ/����w}��� �05�+8`ގ�m&������'�NN�ݣW��G�N��`r�I�=��
kz�j�{""�iܽ����%x-�����!��DL�s
c�OX��7�s��r�(6�n]*<]���w�8�o�zLc7���z��77^8�qJݷ�h�Ͳ�[�w�)�%|3z�zu�'��P���4?<q[J�^K��[؂�݈�Tr���Q�,�µN��ӳ�Y.���'�u��� ��N`:*
�޾�6A�X����&��۫D늍��ԫ����J��4�V̠OT�x��j��eS�Y��\�����B�W��AL�x�j�� 0L���A�K��˺�W4=�(Ԧ�Qy�R��OMN%��D���*"#n;[!����V4�U��|�]FA�#�*�b����3n�"\�U�k����dM-���?<Vh�뭉*�r�	�5����ժ�{������VX��ɕw�W�iB�dW{�f�*�%�oe5��PF�'[�j�K�!1d��{[�[�%YV�\����7\t����#,ٛ��@����n�iu��{O'P��F�15�M�_W!��w��Y0���(<�����N�¨�yN�fu�\��;C�b;���D1Ej�V�Xokr=f��������ݝyL�^I��tq�����#*7{��'IP{���]1N��+��(5���Кb�J�I��p�t�}���L�FK��9}�=I�Z>�o,��n���׬%��)�0�ޤ�oS�K��9JY�����t� 3��0�ZSNo�g3	����>�����N�Mֲ8eq�?w��/7ۍӽ�!mL��n)�A�e�]4�.�ɽ�m��XM�Z�	���Û$��]m��}�����[蹫�P�3[�c5�XjK������p$JK�Gg��[t7y=����	�[9��r�!� ki���;76�ю%�e�����S���\��2�i:�M�bTHLIKm��yA�����^؁�ip�˔�Q+�.1�9�F����y����.�a�78$���1+*�6\P�B	��}4��0�"*�]ec�*l��.=�2���eKu9��vq7³s9Y����Th���L� �WR�ۨN��.^Ʃ�śyӈ�5e�e읫r��Q��FI��2�PݣljJd�k]^��)��=2:�����F(ʝ�	Ze蚓NV��GjKS�D��S;�����p��Ր�4�@��J4�6��o*���	�F�M,�h�c�RQ������"�"�LA��5	��2)2n�O��3�`���to�d\C�*; �#A�
�P S���H!4���h/��"iN���|��P�H�I����)*m��l�!)��� 4ZJ-���P��*M�6��"t4��D�(�F�4[�FR��k#7P4��WJ��!�����T���&��T�f�As��TD^�fSAPwmcf΋�=�F(��/8�Á��u��\#���|���-����np�,Ԣ��x�����
ˡ�zib�30����꙱l�N��P��/�3D+2ut�V��>}Ӎ�ڀ�:&����[�$�/t�����m8�fԻ����Jg�_Q�·b����BU��r�.�$v�T�(t�J�X8�[�:
�PlP��`�]V9���<��؈���FH�+���V�]��ԣ����(��|�{R��.��i�7S=��	|P�iR��Bj,:��Tt�ٸ�r+n�n��;y-�aeެRP��a*p�Ϊ�prL@���5�mv֣���^	G�ON�qKAOHIN��U�E��<gmnpD�}*�U��y���R��*�\�s��I�|����51_�_^�((�qH��ȧF�,�9��{q0e�ǅ(���짊-J�ܣ��`HY�5o�ʉ���O-ho.����7����o[�P��.�+x��1>����E��s�%^R%�k7m�V���A��V�~���v����+ݮ���Pn��蘷5-���Halr_v�N)fT:1r;�&>�Ӻ��){�0�旷G5��F+<F�c�0h�z�4B&�ӎwWm��N
n��/��.Q�:���5�VZ���Z�ʷG=��єe If���|Z�9�Jwt�GWt�Y�] ��p�����k�r��Xk��7�f�����VU-�{�X�xIAZp�����hU=K�,.�f�2�:�L��NK5��[Zd��F��en�m�MvP�ԇ	�ō��8@������J������Ԭ��Ct�9`���6��zH�Խ)���;����k);	mg_��2�N�U��t8^�n�����iw�xPU���(�!��Y�D�vUq{O��0�	�r����útr��<5czdS��`c��o��|�tUShi|�)��ZW��-Ûb�
����2�{NG�uP�W��=�՚�MZZ%���'1id����B�����o�#)ժt5z���Zy�؎���{>�X��e�3̵;jR��i�'b�6��b��Q�8�D���螻�Q�t�Vqf^�寓�-�4i�{3#A
<%v��J���Ɔ�o����(�"�n�!���<���B�E�j��|���O��ٽ˚�^G�����ZoQ�7��E*]�bI��*\�Kt�<Iۭ�����v2�Q�:��k(ֹ�q,�ץT�}R�ṋ�CZ���-�ķ��47�ue�!T���CX)�`�)�8�a��t@wl�Sݫ�*��wՊ18���(��"^Դk�Lݻ���9��N�)�q\��� ��E>97��)om�*v�7u��T�-�PWr
��SH����]J�[h�ƏB/��=Ʃg�kG}�J
����A޳]��Y�����l�Ӳ����nQ�k�*O���xތi����k�aj+q�ϺᥢA-n��\�v��!�'f^:�����[��۷�f:��O������Oq_�5��+5���c[Zup|�f��Vm�����IlmB�4{V���c9m+$��y��
建�`q�U%G��Ó~jN&7����T44�g��h����̮cV���R���V.��v�b�ܕ�dY��r�J_:9,E�JۧX�5�5��]C�ja;����,l�<�fݏ��E҇��VP���
�W
��97JTUki�4AIGd�;Ǔf�i�t˺z��WS��3�c�d�ˈ,���������AO�A���[R�Ȧ�lV3�S$��Y>�+\��/G���w ���c������6V
w(g!O�t�c�u��X��t��t��[�o�Iv���ɓ3��f-�ʙ�@��g�і���g;�����c��l�eR��yi^�j�����+w3]�_'�|�r�y������K��8-j��.΋�����:j|R����wS�d͒JJ,)�5�.�m�7"�1�02D7M���o�2��uL�+z`W�l�^K.�5mw$ɔ$��R�v������C^9f�e9��D&����Ll�����T$�mt�u;S����5��i!t.&��u�8��LEַo�r��[2�i��*�O�;�t��Rpt�]	n#�:#�e�B,�e���M�23�q][����$��5t��2ö�>�xdݠzVNxt��tEn:]ڨ��'�#u.W`�Si�@
�>�%tg�ͩ�<D,}םkjj[3�:�[�T0G�������>�g�)��y�'_=Y%��̥���Ji�5p���X�S�
=������� ���Sp���Y�!䁴��K��Z�r
.��7tMP+�+k�Y��A^�D
#���C7�ry%F�um�{N�������Iݮ@j�_S���ү"�5H%o7���t��0����yh� �͓��<��/&��,Wg'bRd<��^�:�gv -s�Վ�H����TF�kmm���8�f��f��a���]T�K�瑭,J��,|�Ʒ��cH�:�=��}K��KE��m����+L,9K��Bb9���e*R�J�.�ac]��Xn���c=��]��
�5��,�)��&��%d���瓴��ܡ�י��x����eHs�L��8�]���}ʅ�ݰ��n��p�e���M̭��N�H1؞V�g��i��N��ugSU(����P��P��,'|�O��]�TW����U�nL�q�{�]� �gh�K,
(}YTъ'q�� �~�qV2Gy�n��Uµ�$o��Q�=Oz��1w��o���Z��tu|�̷\5��GF�e�Uո;��wNb���/0����;��K5-ݓ����y�g��<!|B�7h�V=�Xo�3x�.�t�j�ȗJ��'��b�}n�+\>Y�;����Җ71iD���Y��.�e��-�V֎uY�!$k��w¯zͶ�QW)�~t�Yc^��yY��f�Z���4�,��	5��d� +<���v��fC�n���It��>�5MH>yk�r�h�l-��j������Y�b�L�$�F�
e�����E@�lc	v/E��`��<�\źO^JԷ�P�0�Ҵ:T�gk/_>�"鴎t��		SZx�xA��oh�:�J��r�[�h��ł�)��fIZ�f���ŷ����o ���8�+#"f�]C�	�{m�tP�彅W�g�7��\5����܌����A[�S%u$��;���m��w[P��M�Wt���SR}G��[7|��Sp��E�;�t9I�'WST�C)o_|=�c��\u�s{�wQS�c��$�E��T�q����y�4S��uW#M���h�&��)�/��Y�� k�Ƥ�WH�
�Ұ��ը����"�+�TR�M*5�m)k.h=Lx��0-�2�\��l�sp���R�ra�u��$V��Fq�ڝ��� ;G'�P6�P]f�ρ<�X�q�shc͈B����T/^�vi�W%�i�s>���g_aډ�̸��[:<�5��k�)��l�mGܴ�r^nC�W���KML۵]T֚Zz��B<n=�ג��tiL/F�|-f��74<�P�ѣ���ZywKw�ج�ܫ�KX�%ƶ���y����=�U�lI:�Į�7wo8�r���I��	i(AZ_�ڍ�>c�	��K;���Ot��8�V��Q*7�`����'5"���"��b�,+�}��QN�ƅ}2�(�&����7o�i:fqwe� ��T��j�l@T#�����Tn�5)Ō�#E�ԫ��[Н���X����b<4�=��W��|{�����}6�g4%���͕n%�͓r�F�c-��0�Cq�S��
�B������h�X�)�>�s�t+B+�6ufX��;a�MA%>Av��MY��tΘ��N�]8�z�Ȗ|�`����	�۲�7�j�uY�|����Ӊ���K#�Ij�r�=��)͋c�_^�k�k�U���Y�Y�#P�f��P���3�ט4b���Z1\�:���p���o�Ulj���nB�r�igk��gu��+r�q`
}q�!p֊M���L�Y�
��
���Nl�
��E�q#�h�+͡iѹŜ�/:���f\�AS��M�uWf����{\�f=�#ƹ�]�
�ӯr=|������R!uu-1�k`ݫ.�r�'�ܱz7�e�X%�/�����Nк�uͭ��2���ni�Ck)1yWZl���y��U�0�\0�7�̸-Z]Ђ��@��ݰ.����vƑڶsν}�=,�|��������ˡ�;"I�� ����9]*ﻂ��Z%fǠ��t9��&��I�c����.��P�k�ǋB�Ȕg��}���b�&�*A�0ۗT�^"a����2b�nۧX�p�P��k��O�oq�:�x5���
o���y���x�F�g.�]�f�dVh�d&��2[���%T�|�LX
�9��\ZM��B��]��Ƀ�ln�ֶ������]���Ⲵ��Y�K��{;�ӴY��O�e'��Y���������0�{Y@ER�GH}���0嶂@6�k�w�MS��<�OD�)� mv�kU�lq��<7�9�a�OQ{IC!XN�^&�7ĺq[|�0��v"�Z�A�
��b47�.W[�r�Vf�������)f����X (�
G��a�ҴI� �[��_!�����p��@�Y�jpM�!EG�n4��(f����G���Kh�$�B�t���Sr)��\�R�m�1�d�-�i#���L�ڌm6\=}�;��.����}���m� ���]��*I���u�K��-ru}[Z��(��R�fZx��]Ԡ౴�A7�U5xLC>�$Ȓ�2��v*WVk�t�9X֫n�?9��u0-��r�_���P�SCj�/�kn�p9Y���Ӯ6BA�7V�e�k�ǯ�i�Nە�� �yl��4��Ǧ�L����goFg*���E*D�Xw������#�cy��riPnu�9��L	�j����Λ���X�v9�e; V
�ͽ7vC}�� �J��2�(��������w]t�#n��yß�ع:��l�I����
N*�x<	�2��>U;j�����b�Z*3X�z�k��_LR�Ѽ��a��4	�0Գ���۹�{�-�Ȯq�/�n�n:�%.��s�HNRi��/
��8��R��s4�ţWv�g�ˍ_N��˷�O�{����۬`��s3Kƥ0v\?*�2���9�{��͵75����5���]GD�ع��^�9<{�:�Q���3�T(���x�p�i��c�-\�%�J��٢��Y��{b>�٠�Ͱv�a�"�#����j��V�7�R��y)��Gp���!&ܙ#V�,fU�W8���ƙ���\5!~��߳D-�Μ�iX�Z�y��Sϙgݒ��x)ҍKӔh�.��Po+��P;Y]�'��J��+�ۧ"��"D��Lm�7]:�ĵ���,���B��ǽ��*㍢�G��\�35��\jsre���T*c����Aؠݝ�vb�wtw�ǵ�	�R�k]��ŭ�dCՌ���֤���wX%n�z�m���NV�eS}��]����2�j�rd�W���먐eR���;�cT�1_Ks�nq�Ƃ����@.�+u�N:R}i����z~�- �gj�@0�Y\(L�v{f��,�R��|� ,X����rd���b�&
7-Kx��z6��p��S��Y�%���f� _x�]��E�K����4l��v.����v�́�[hf.��	�W���T�LgP�9��7OCx���b�RX3+��@�M�Z''5)��8�t�a�]���©��J�o��B��q�Mf'E��bg	�^ak4�Ck�ml㒞i��R�}oC��ڡA[{�|FV��ױ���ꋄUk�Ky�n3��V��ՒX=��_B��-+� j8WBb�T�%n���J(E kYc��aŋ0�tK���guV�"���"�K�Y ���#�B��@T� K��o�
�/�j��3E�i��,��Ba����X}z�j���R��Z�v�������1t��P9���6�S�z��.�$2��h5���;Ъ�{��T���1Z�}Yk[�K����|��#<�əp���NfB�Q ͹�� ���p�x�.�&�"��^N�[*}[{
i嘞I�?	�˫TRT�=��GخG���yB�m�� �"ݣ�ܭ�F�����9Pjty�:��l��T�I]��n���:k�A(�F�� t^`�DG�d-�#�j��)��'���}w�0@�#Ί���JW�u;.�h��U�!�,�m*�Qܧ�k0k�o�]err�cͶ�s�(9��os5d�[�]E��oA�*�a%X��ڸ�(8K�&�{R%��Pޔ���_uɡ��Ѩ"���}���D�gծ�E���%V67C$t5����*�ᚭ�b�0L��z���7���$���gs�
��B�R�P�C�L��$�L	��WI�fv�~m�Y)��8�)�}V3EX�eL,��	�8�dU��������q�V,��g�� ���,vj�!��\�k�I!\����UıB�R�y�I�g8���Ԙww6�dr��ا*�
��^��wM��IZ��MnW���}]M�ĳ�yZ�S!]'sr��Z,���F�=!��+VRo��c0��U3��Xi˶h�e�1�gf zK���ve��>o877����P�>���Q%��`��,r���L.��
�i|�a�� 2�_»�ڮ͹qJ��a�gպ�]�'9��7��%۸��|�VJY-���/y�k5���D�[rRy�3����U�9V�X�r4 s���?�~oG�sM�G�GG��ulٳf͛88883lї���?����a:Kq�3�Wu15B,6KJS,U���bϷQ��^������� �v��#�7v;��9�&��M�!dU��m�o-\�ձ��)^���83&c���`1���n�^����\���)I����T�h�գm���`'��y����J7�Oಧ�1�����ҭ�{.Z��✥<�QT�5�=�Kz��S��ǖ]	��V5cD`��K�9���Vg[rJ@���+㠇�ݜ��I�5�r�U��W D`:pe�^b�]!�ՙ
�&˦8��_'0�['�Iuv����(�G`=����4��n���x�Woba�2h�)�˲[^����S�d[�kB�QO�m�J��3sV�?�={0�Ӛt��t�.����:�>LQ�{��j�@r̎Ռ�4T�zmPE;�H�����..���ܨP��b�s26]�^���S�4���H�\�V<W�������Yj���2�,݆�dM��n&�4��N9���r]:��O(u�}T�7��+u�]*=�lp��|���J��Y
�D�#:��R4╚*�����9�{Z��r��r����L����U�tWG��L��ϩ�_	�r�����M�닭Dŭ҅ˡI���f��D�F�m̎�j1��@�u�@�n������8���i��0.:0��VPި��Ù[%,���;��S���ObP�i����
@�.�
.�i��'�4A��:A��	(����ƪ��b���)�����)�v�[F�J�����f�1Mݹ�T�4ŵb��*�"v��Im��LUhcm�UZ4E$�5TSQQlh�*֊��5�LT���T�Z(�AEE��$I�h� ��N�誘j�S�d�UT�T�4T�PT�L�DCTZLl����f
(�"bh��&
*�X��b������S��֪)�64�ٙ��cZ�&
a��T�TIDV���&�"�*f���Z"���&��H�("��(����""(�����;i*��(��*���������a�	��$����jh*����M�=<�}�����Y�EV�{Y�&���F���R:���+.��+��ܡ �b���rvl-|/,���vnU�����p���/�jk�e��Z���;~�ҡ�"�ȯ~L��6�����Y���Qnֱ�~���]���-��wG����������,��xSwc=���"�G�A"�ra�_���C�H�O}M��{��;F�[�~ã���&i����E����7�o�ٰI��>�9Zy�mx1��׵��z��HWS����E�º���;�KZ_�N�}���z�y�0~fC+�n�z�u����$�r�n��g��tL��r�}$�ڝ�o�����~�R���u��^���~"?��M�{�iM��� ެ��WOzmTQ=3|��W�{�y6�R�bxH�䏳�?gz�>�ԟ��o�uCOa��{>�r?3=!�^.�N�A���&t1���~�+��Ϡ�q�.\��>?L�����Rb��I�6Vm�D�D�V���X���uh�9�!=/���|��O�8m��yr�~�t��`Wg�Z�[W=Q��uB�*��b�s[�װkL�O3"W74�4�<��˱8pi��ukH�R�e+۝�P�t݋u�+�gAz��ަ�<�}�M�KϺ��W�N��*���w�k�*K�}���2<w��g_z=
�T�5<evS�t9V�}]�8_D��d�ԯ}3�04����tV��(=T���2VT�7U�Qag]Z�(su��b=�zb�<�4���#˔�o��=<g6���P/~H�yz�Iw�Q��<#^��^y�X*��F�����A��«� �D�{$VE�� �n�h��3l�Gl�>��~�#=����j7��v�H��r����A�=$_@c�yt$;g_��2<㽯����}GH����7%?���q{n����t2R�[K2绷�'�&z��T�w����v�$�s�'\�\[���Ou��?�T����@������[>k�3�8T�$`{y�wM�PҞ�ߨ{�n�/��w�7�lkɐv�m���*}�bz�l�����\���E���1��A f��1O�
;�x�������:����ɣ�L�]��i>���<�z�7gW�󦂙κ��w��q�怙]�<�����ܺ�r�i����'!�I�2�H/��g4��z�*\��O�I��z���n��ĕ�ûl�\�*��U����F�����/�W���wQ>�ǺN���ʖ��������}ֲ��p�z�ldeW�{��s�5�M���͕�N5]I�Y7t`��?���`�u���7X�~�7f�8�o�u}�@�L;��{io���z76O��tȼ�y�b���z��kj����Ů�_{kw���,�i����7�Ք���?��;R�2��Eh#j!�M�����`���8q�����2T���M��1aS���x��$���<�UO:�ᄵ�zSt�.�L��J�$�Tf�"f�|�3b���nAn��^�Y�y�[6>�2��%mOS�p!�����yo����z��(q�Zō~mTz"co0��$��ѯ���Z�`W+.��YϝN��ܫ��^��s�lu�J���K�I�5��Hh���e-����/RS{�����V�^]�+�-]��TR�]e���R
U��Ӵ|I>�m�;3}������{�K�|H�
��2�[]�O=�#�1v�N��( %ߏKi�
�����I���x���l��Q�˴n�|�����z���vv���ɼΊ�P�v����g~�9Sh�&׼������&ѫ�x���:����p��:ya{�n���D�:�m ���I�&z��϶K�m����|�Y��Q��zw�Z�5���5��mgs\�C�	�&���A��,�yqo�e�����ʽW���4\=��9)�@�f�n�&��{���ޒz\�GGq�#���0�����W`�y�M��E��}��d>�����_��;�z��½�#��'��~�^���� �����" 썞���7v��w�Ŷ���%�q��6c�U=&�!�.��[\ ��c~�x�6}A���0�}��:����D{�~��'���������b��՚��6?O5S4���&軓î�+N�@�͠L8���U��2v�n����i5�n��VW~$m�
+ڶ����,�ޝ����:� j�����a������f�=O�"6�װK��mmf=��rU�K$��S�K�}��ʇN�㛌������e�6:"�ĺ�������h^���P�$���rt��ᰇ>|Y�-��r�7��.�c���L}AM;6�^L��p�GW=H�̗8<��`cN�UD���db����C��`�L�{y �Ctl_a�x� �8m��U��:��o�r�R4f�k��U괲���9���p�i:2f�N�M��w�xw`�q��(�ا��+���}��S�q��[ͼ�Wz�����7;#�=�a�6\k�j !���VQ�6)̍�X��X0c����c�0t��ꓷ��g'^�lf���n|jz+�}f�9G4E��N�k�����0y�>�V,�%g.�4��nW���ڣ�?{g���;͸UA:��'����puG��^$np�W�����3ޞ���X�w[)��#�����	���
E�cm�@��͂K9��S��.7r�n�o���7�c�L�6��U9ߒYR�({�k%7�=�f��=G�����9�r6�3��<l6ɟ���t�� �m����z�����wuDT��f��;�&<�集K���z_=��㷽�{�f��\�|�ju�=�q3kXغ��{O&S��uv�L�;*�Π���\��v�N8;�Y��vv` 1����D�fT	��lpg�/z��t��U����=�2���9�����N�����}�6����MZ��s\�e]��ܚ����{�Iz�����oM��&��ͣ����[�sʛt�{�<�y*C+I�Y��^�D�����sg��0rw����D�[ZbE1y�WyKs�,�f٩�a��[𭫯<x��t���r���z�}�n���jܻ��v\ʳ�$���Bz��j�T߭Խ�U�2���*R*�}�\���$ڗ<�8%��T�jz�������G]�L�������ʺ`�2�����V��@ff;WgH�yow�l�+$�"��h{�~�StQ��@w=�q���#�������uIt��ɻ<+�E���G�O/��Z2n'ݙ�LtlE��w&�39qS�����fA��ܛ#L�^��z�}��j�����H�Ш�����]v�9��ing�ʟy�4x��Z\���N�s�9{q�66{w�9�י�l!��] $�r�e?_U��>ʱ�0��fr��>�^�᪋��s���ζK�4��W�n�=L7�l2���h�Y�s�{2����%��JS'B}��69�Q{��5��wI�M��=���\��}�T۹����pA�"��0�{�ܝ�3c~��?>����8���O{|p�M�[,b[��H{�.| ���N	�O�m�������=c=�uA����zx����s#[�8Up���b�f��K�����CH���t���`7o����yF��֫����^��Q��(�Ӎ�7�����ᑗ�{��;��:l1�:_A��,�0���ѓ����j�����罯�����4�A^���|��'oM9��V��Х>@Rg���^s~���n�h{�A''���{�w��w��w�������eq�n�/�S��K�^�k|nM���������D�OT��#�j�"�����	A��>5����XOK[�[�uq��4�msߚ����<&�Ԙ�����j��߷���/�%����5�%�y���( �"��8��ww'�5�����f���,�hfa������l]�����N�ډ.�����;U��w�
{0�g�35�d�3�V���Uē�fu�L�8�. f���� Ʃ���N�s�]�:l�ݳ�T��JU�)OP���x�6*�Ơt���*g�A�^g��^��ܜZ�����^:>�����Fu6*����M�[R�}@%��B���^��g�8I�#���u����$�F��T�v�{ޭH���q�<�H��g���8�7��S`��7Lce��9#{���2>�ew��y���m{ȼ�Q��{��E$�6۹柤Poj�~�K}�k�>�w�7�y�9˄j���_M�����r�l�[l��ɦ=�#�Z��{	�׆xA^�H��[p�Z�@��I�x&�$�1�u��ny��D�j��~4���VR���4%{)tS��~$�<O�d��;b��q�l��^���l��r߯�]��*��T%y�d���<��_m��}O�y%5O*;�k���W/v�9ϓ�����S����� D�{6?��5�KqxIZ��WY:0��9��-�I9L��N� `=�����`�?d��u�J��Ss�4W�0�� �N-e�q���e%b�QD⮽W)V��N��84�tR�ف�;8:Xf]���C��6�=!$�=tc�n��֮��ˢ;֣�������`��~�+�~�f�����I���`�-�הc��8麧��'L_�O��ojg�2zo��o�*�TM-f�|�������ტӿQ�"���/uM!�Q����~�\�v>�'�{�v ��m閝ܜ��I7Zi�w�����FH9 nvϻ	��}��x;���|��V?6���b~ɡ���2�νc�C�e^"�ݵ�y�f$�Fᬨ}.���ә�Ђ3]����/w�ws>�����T�W��'=���}nZ��.��ݧ��6������z@%Ң<)�F���svL\L��ul�}�A�~����of@<"����4D��Y'^O�lJ��~R�oZ����b�]b G
m��rhL�Ip"⦳���f�ɯ{�e�g(戩j�$���M����]B]��&�ce����&|(��3�M��9}��y�s�U'�]c�;�Q���(v�L=Z���uP*���j�#_ڴ�v��g��5��2_V�֣H|'+��=�b��P�&z��^V�1�W�t�w�T[e�����~te,;�h�����s��SkL�m����jw]�=Z�pO��/.�q�խJ�<����?\�G�X�K~�ە��>\s��l��Vd>�T�ީW���5dF�e�n�G�%=:f�_���U����,N�Բ�q��1)�*Bv����~{��%�%��r��>��y�Y'0�Rlۤ*�Ez�]����O[ю�2�u�xOq^�-3}�Cx��~�-�{.�V�*0[Ĺ�-����{|�X��&�n��;{j��H)�R�W�����R���Cq�����q���4g}v���U*w^Q=[��&���������؝�9��zgwZ��>ܡ�=���Ѭ���0��.\����I�ma̧����u�����o��'��}Sj���԰����y �m��8�e�,N���-]���`��~���3>���f�1{_�
T~��I�������׬�����������z�������Um�)��������-�Z�:��f�*��$��'e=Z��\������K��+j�;e��"nh�H�ܛ-4�ssEK�-w)szy\͆��I��I�:�f�*Ǌ��ܧ�P-���M�PyFr�wGR�ѵ�R$���j_=���!��<G�j�s�HwE,�9}��C���v�X���up��ɐ���B��gd�A3��e	x�⺳s�R�� Nu�"`�2ȵ+��2�i�;+����y�㭂���4�Mz�^2U�W!���+_0�VJ���@�EV�]�8�nso(��W���� ;��A[0�6�n{8� 97$S^�	��=I��C�ڬ+E�]���uv۷jHh��wC�q�z@��������J��Y�#�y���e�q�`L�Jͅ��^.�e��B���h�ꡮ�3���cN��Uřck$�PUظ�g\o9R��]Z2eN-�l �s{X�Z�XY����'pƘ���	Yt��8��Ú
,=1��;��{�j�ا��#��na�*���ΥÎ]n�Mdej' Ҵ6�e1QtΩ �޷҅��V���TJ��r���è�9�gN�����8��G�v7p
�6ok�mల���u4dD�ΡLvֆm�f�5�Gk�$��4G�e����e��2�(]l������!P��1!�F�	���8�>�ǌ.��fc�eI���c��i�&l��*;c���Ki�ϭ��HX�ʛ  >���6ǌ�q�5n_(�n�#�
[�E�ot0ԋ80A���f'�w3/�3�D{��IH�e�>�.�}�6G���_������2�gwF�8ƞ֑Q���k2���V��0�&�jྮŎ!�f��V�]�h��n_m�-
�L���S���P���J	^�H;U״��lL�Sw����m���L���<��$c;.ت�C S>]le�j�[�[��­!b�l����:�r����h��OM_�rN�x�5�v8S�4�n��$:��V Щ��F�� ����n�c��6z��G��n��S�f'4��F�=��e<Z��{*g@)��n
�X ]�ڔM��e\E;��z�����f�*S���o�e��\h|,�!.'���ҏ����c�aطR�$W����W�G��%V��RŢnC�_eL:&^�N���UJkl����Y��8A�vV�}��G����k^�&vF���U��!�Q�h�s"��w�z�Ѵ�!A�~��l�[cz=cV�8��sV[�t
u���V�=fZ�Nh��WrYт���#ub��8\ifӬZ���0�D�7��g5��ړ��iaR3k+\�I�xM��V�;��^��.Q�ɠ��3�`�����٬Z3'z_n���a)̈��7q��b��#%u!�`m_c�+z��75���;΂_���    �QUUE�j$��g�uM3UQE,��PABUTQEMDDPAD2DUML�TL�Q:��L�KETP�$T1A4EUQAEEA�TIkU��(��6��MUCEUAML�E3UM4Z�3�MT��hqUMƆ����"(��j �Fb*��Q�S1��h*b���
?,�4�"ƈ�[g-O��\�Uh�DɬESͦ&��MDm�Jъ#grt�[�LEW6��5�"эk���QVa��Y�lD�V6���na�rh*y��Z3F���rh�9m�ɠ�E�-ۆj�=`�-f�Tش6��;p�.�[;c�$V�")*-�RѭV6=\�&�<����QQU�b	!��`�ٹ�rZ�mr�7 �s�卶#8�������w���������*��ޗ��i]^2*����k.�j� V�z��HF_���mE�E����ÈV`m�mG��>��^Sg�:�n��Q��ph1�������Dx �P��􍈨~��goj�I�� �7п�G���s��C�rz�T[{�wT ��7p�4U���R��K�{ؤ�K��%��gQ}�Y[Џ1x���?W�Th�B}����,��#��ݵIS6��A�z�F0LE�c�s�	��+�`kȤ�P�Mj���~56�08��a�y��O?���8�+Q^��Rjon�eÇ��F�[inݜ��2����^��|gXW��ǯ[ո^�o����́��DC��A�ڨ��M���O*|�ۓ����A	�xr�d]% S�R��b#��Q.���	�[�u�V=O�O���J�K<S�?-崵S]�>'rO=���>)��ǁF�[\u�3c�zgG���POI��a�����Q�~#>f-�vK1���Ho���Y��$�*Iؼ�+Z��l�Ǟˀ�Q��q�j��O.���L `���!6���ry�9��q�M��b�R�A.W_AU���wYU�$���I��&�ΰ�ar�F����0�lĲ羬�n��\�]�=�?ͭ��`����_]a�����c6��\r�=;J?w5r��)^3�w�!u�%U��V�^�ᓯL���E�o���YSs���;uV��N�m�.8z7J�i��~[6��ǖZ�aSDU[F�P:�-�Mh��Wλ�c
"�>9K�Zlt�mm���{7�1�ĥU�m��_��e���%ݳXF��q`|:�`��"��Ό��>�of���`��wy���}��.��u�\>�����H���e��<�@!���������h������3������o͏{�W��Q?0�ϯ�X��w�^�2�[K�g�=@u�v��?3��X�sJ8���9�sym��|>t��kb{�b�j����|��s7�q~$@=��K�,Z���]�Ɏ�*��矏�K?�,�69�c�R5�Vu瓸hE{�Mj�1i�0a���n�ݏ�"��;�b��B����o�0����C@ێi0�u~κZm�hT��~u@'[�� |�x��þ$O���~�w���|�c�g�E��2��)�~�,=�ҌEݿ��ۯ6�t�T�p-����5����q���!�R�%�3�����T2���p)��'�!'v�yo:��f��OU���k��
�**��:	����q�ڗN3��{k��s������r�l�qm�zԛf����qp�N�nβjɃ�^~�:װLRu`b��U&��qm#z.7���3{2B��U����&�����$xl��+Y^�.�j8�u�5�Ec���.]s�>���c1y-��ܺ�qe=�bT7$$ <���Ni�2!f����6��]V:�V�
�.�G��f�B�e��E<��|����g��ͩ�����9Y��u�^h�qi�:�sK5Yaĳ�D[{��5���O�%ۄ�Inj�D&I��N�$�Z�TS�oM���U5ʡJ�f�C��2�gO�� @B ƟC�;�j�5gC��LS>d��;q�`?8S�iocQ�B-��dr��8^���a���B1��O�&��"<�/�;/���-�,�΋�Uڪ���5l��bҴ����z������`���!�n�yO��ަ�J9���STgI|��Bs�y����6������|�Ƒچ	�DC�p��@����Çߕ�jpx=;=�\:è�u�QX�c�(Y���.�*�xRΞeJ�Xo�֮݇{p�5��fs�c��녢��+X�9mi2:����suf��j%k���+�ʂ^�¨��v�����գ3��,2�M�C��P?�G��B��O�>A�R̶�m��@ߓ�ֽ�a��Z�O��v���Y����V��|�f�'gd;`jz/a�HR%�!0��oו,�:�n�s��)��ٞ�VV��V3�۲���ޖm�*!��ƺ<-���^]�2*����!�>0���d_����V��斝�Ё\�w�m5��=�.^��>=�����Ar�k1ʻ�G'9j�;�/ſ3���9LB|w��򬞒e�c�ޣc���ҽWK݊E�w��YYeEZ��Q�L�qu��t%0�vL��h�s�*́�e�ܩD�[gj2;�����]=g4��5cMCصD�1��S-x��'`3`."�@!0_��Z��d}EE�Cp��[z�]UE��XݯN6C�����P\�5�ӦΘ�uC����"F�v�.a:4e��~������Nd�=�
�֥s�-mCQ����aZ���S�:�㢛�N�2�7hK�櫎�]�yL=��L��5��!�s��3���T�3s��M��LW�����4�=�M1��[:�w;؁^=;ύ4��)흗3��.$�����|��|����o3�E�w;n����=x��)��2�t���9�=k�<'�o��@���Ɣ�ژk�c@!��k�=G	Lb��G&�&��]/*3<��񮓩�Lk�*L+��s�{���5���(f��L8�ԭ2�.���|9�3���B��OU�y�.�_��S"�s�%�0�|`Ӗ�p���L��[`�䥻����6��m���dI8i;������!�?7��7�K�d�8�(T���>�{Y�a�P|A�z�s�h��}nͩ���N0-GNл�*��z�w:�R;��xŊ�L��؀Z�s�6��n<�.��)\�su5e(Z2�)�9����f`���v��7��5�g��Z���|�7�f�3ip�H��M�;[Ă�ᇯ�|F��햱��y�<uT���9Pr妨��u�}��;w[/_Vd%v�U���.�LDkg�{=��p�,k�i�_U&�VK��a��J.��i�F/P��Y��~����.��L�w,��L�P���G�{�R#O�e�7�����Ϻ�#���ػ���kr/�l��rb9��ۖb|`gc>3�0C��<��p"����U���u[���Ln^%��ID�Iy�lZ�X�c#�]�����zwgbf��ɉ�;���t�"no���5�&|�M�v�~���k�����v���R����0j���`����-T�,�sKH����lS��/��CZ}�p�4W���%T�7��p��uϛ����� ūy��3��]k�(p@˥i�z����d;r?�[�m�%,��;(2o%۬�M1�3��gM*a��nC�x�kVz3^��׌�S���P)G�˪_�����_F&f�^�T��\��4��������֔�{Q�o
�1�ޭྲྀ;��_G�K���������VՎP��,���(td�!�'L,��IM ���������]T6MR�^U����gw.�}��1�1�'|�Yp���?���<�����g?e�w*���rtG�j���΅%OZ�����l�23�y'ޏ�	8�}�bˡ�yΤ飢ڢ���ͬ��JS��4���2�^�	�1��&} z�Ec��ws�)�D�4!�KU+������z9��'/2W�fϽ1l3q�!� -~�N�ሔ��H�4Q�����j�p�UV�9�,�Z��d/{��c�S!��f�!���v
����F�|s��h�m�7A��ݬ��ԛ4r:5ٲ�s��s,"�hA�AЄ���7'����0�rt�/I�?�c�2�^]6s�Z��Hp'�BF%����l�Q� d��9�{�%�{�5�Ll{
�ko6s���Φ�9�"�"v�79b�p!� ��LX
���3��b]�=���!��n�vuduP�t����Z9Ke��4�1�]�N{�m^���w�)'��.3�뇰�}�Y�^�ٷ]�h!���_���/�-�K�W̏S\�&/x���R��j�j�Ja�^5������2�z�{(��";�P�U����	6�Զb��YG�*g^B9��C�bzچO�	��Gi'ә���1��[Q~��PMh;��vO6�cw4o�K��-��`s*�ܰ�0�}�#Y+��sϼw�L�v�L��-f�v�7��E��F)9r�m�u�p&�:�D��AÈw���u�S���;�љf����oW�{)����Z9��_R��޹�X��!��sD݃�jE����l��J�-$�Y1fº��N�����kvY�R4�e+�u۪�଩�;�ґ֧�i���
׶˨Y�Cz���e1� m���A.�z&n����t���^��[	���_C�)ǎ��\�s����� �����Ϡ�q[@t�.��0�C���֞��6�hl�w�\E!��["�Us����6�>h�O�b�1v>�)`�(8�,�2W6���=��T;XHƄ�^���@�!'��z����A�ɜ$�>�YϬ�rGu�ȫjނ�Xa��<	eA.�g�c���Qp�<�|!?���50���)�k�h�-"u�ׄėi�ޝbՓ��׃,} ����#B��T�S.����U`��D�T���]�a�lwy⃖���,�{�����v�=����:!2O`�Jp��ZTj~5�ѫ��qu��[��)���<Ч����Yמ3w���F4��'&�R6��7�.��F�&�b��Z��^��7gi�.�-�B�
c"��&A A�/O���n?���i�'� �~�ɽ�gmC�Z��õ���������M��Bsr���MsӇ�~y��Ð����s�SF��~�~ո��dO_Ia=q�����{*����(�C��͸�o���ky���Z]��^ěF[m[T@ִ�V�W:��o�$닰K�,!gO2�WZ�|^�>�sۇ���浬�&T��˄�<�.���8�|�Lp̣�~ɪ6a�;+���]��W�4d�ߦ��-�Ԩ��rV�}T�Gḩw`��>o��=�^�)#'s�]�O�����q*�3v�q���(��ӯ.H7Ij�>gcfc�p귉�m����!���{�iG���`���>4�PX�T�m��B��D�q�_�s��Z���o|�ֺ�,��.�b/��	{��a�e ��3���p؜�Գ ��m��@�~��b��0Q�"&Q�w�ʹ��Y1�_A{�@2%߁p��#m��
a.�:��f����3w
`��.۟kR�u���������2�t>[�tg/<��t>'�y/��A�ۡ�lG���5��T�/�p't�C�*(��N��U�6�ƶ6��m7�Y@��u�o�3V*t�hF��G�'ت�Ƕ��Ɛ3!��/���U�B��ךE�ۦ�z�M�n|%��!�ݯ�s[�L�@9���"S����{��j���K[iP�͏�aT-e
W䨷����Km�'	3EU~/)2~�SC��C�1L�cN	��}#���[��fJ��KsW���2m&d�b������܂ڶ�,뜦~�����u=�a���B�T��i�q%�͕0���`:o�q�^�e��^]���KR�K�����&t���F�c�Z��	�����*`�
�x��38�)�\�S��d�T��^������xNZ�٩劓���nh��֏���W�d�ю=��ط�.�7ݐW�&t�˝h�3�%E���[��R�(��0�*��W��v�u³UI���n�\�ۭ >�
i m���#��� WAy_��}_U x���H���"���z}�2��c K$�tS!*L)�+�P{�����	���Y]�휳��Z�E�s�p,6O�D������]0�jQu�_�R�Q�~��ڝ�\�Mp�Hwi6��j�}
Y{��2i���&��c��У�S��8���,ŧ�I��'�p5��#z��7���թ�P��5̆���kL!ݳ��`X�3�ad�2��w:��/�4��Y[3r�F(�t���D��Ɨ���x�!�G�í~ىm]2Z�/)U�����}zx�	�j�~�����
i�턞��pw��d���b���P����u�S��#O�����N��֔�4W�E��_�E�*�+<u>��}&g��`v������T`��D"�i;�,_+41�l~��ߥ�s 3b�_����C�������JtH�MW���v�Tycf+룬a�A)Ĉ��Ǳ��Vh1�����!�8I�i/��z5�<�-{��q��y�S�ĳ�-- ��}lO]Qx�pwP֝�4���`�e�AyǶ!=4�v�śumO50��U�ڶ�J��YLnm���kv�[�%œd*=�GW�r��p�.�Xv��y6�V0Mƹ\���;xe帎7-����K6Y/3 &i�8ks�|
<�<Rq*m�yIо&����:[k���f�^�< �a�x7�D���X�p��\�=y���p%�c����>���{�U7�ϻm�ĕ3kzv�{�B\M\��{ĵ�Pb�
�a�I�͋O��o
��)�x[P���Eǧ�	U�m�dm�h�[�s=��3o�<��^K���޿r�5Ji=�(�0<�o�ޭ�[� �d��am�:7uߥ�k���V�u�9�9}�d��hC$�5tA	�Ƚ�%4��*Mw����c�߈�*��{�ڵ.�Ox�������1ٲ���OcHC�{���:.������Ɗ4����O�٨�ɗ�(�Ո�+�K�˨��(����jc=��NK�R/����2N��?�E������kQ��V���\�
dr3^�#Ͼ{aD!b���@ܞ����Bn�����?0�s�ī�9P��5 �O��ח'���a>=��.�`�Za��6bYs�VM77��2��B��[�'��s-�`��01��uٓ�x�b]�_�!�;�����'��3�Z�n\�拭n0ƻ8��j|)�AU�}Г�,��z5F�Y��-ݛg�a�/"C�����~�����_�>?�^�{���{}��_��"D�k��-Q�j�����x�l5>| V��Q8%��9��r74�e�(L�������X��v>r_:���1枍@Gs��N)�Mn��}�oL��n+GgDt\�E�=�D�/�|�w/E�-R���tYl�!7�M@pe6-��ݬ0�"Ro{9k%�aPL���eee.�7�dR���
�0��.�1� ���L���F��;v�#�N���D�{	{Ϛ}�8�:�KZ5	.%�K(wb����(Q�U��v4�sZiu������������ਘ*�y	�8��ĥE��5)�����io�%g1jø���{p�M��t3䛊ޭ�G��Z�p�;H�k_�})K�C�����I�P����5�;�N>���dth\׶Y���2Q�\Ɋ��V�}��ܭ�ź�8\i;*��H���)o��t;R�̀��{6n*����/�2�TnZ�����<��U�ʴh�SC�c�[��|�=��Q��ͮ��K�$6�dl-N�����W��]a�#67(R�W%X�"鎔/�H3�]f.w��]�Q
A��{��ջ&�#W���Q�n+D����n�WYԩ��ՠM����d!���|6��WV��h� =:�y���2���O+��
cqS1��ԩSd�߲2:��7�V�8͌kS2�y�@��������.�S^f�ج>"n����`�/���[�Ɛ����;$�щl<���![�w�b-� �Sq���h<��v���Gڱnk�����4���[�/{�&�65*���VO�x��+����fM�{�jru�*=���6��k#�sj-h<5-�]�ͺ�X�P�h3��i���Z&�/���a\�9�=co���!	Zf3W�aO�8.B��+A�Z���22j��۵�[�:cL�����f�;g����r��,�/��fS��=���s�o�nڸ��7]�^9;_$TivwD'[��hCQE�]N8�%�+U��ɺ&��oQl�H�f�Eiو�V쬴za ����oMq�ڙ/6��dxƩ3����*��mLY�N��y�I���MJ��$)2*6Q�.U�CgiC",U���PZꏤć,���A6�ɳ+��άFL�ࢦ��V�e!u����ۘgNNNEv�\mw94�n�<sԈ����S�2�T�ˊ��kP��r%/U,�ז��ed�NkE��D��:��]��q=@�Y��W�H@��P���g
J��jb�s�q�6�mm[���#K��Oo��F�Z���P���n��T"�\n���:�ޛJPP0u�=#����gWr�34Q�ha�;�d��kI;�S�x�M3����F�[V�ۗcg���x�3]�2�Ֆ�Ky�u0��_-���V��V
L��Ⱥ�["Ê]dN˘�����R��@��8��gz���(�MB�.�q��W�-���O�8�((�*���T�]:t"�R �R5	}	��r(e/�������:���U�gzn�ߖѽs�.nG9��1UEF��N�qAU��'2r
)�nfv�j&��c���9��1<�� �f�mb����i,j��6rܝiӣNEV�*��EE�T��9j�*��0j*���"��0�1�LD�k�1�h�"�DUU&���yE6.A�)���
��D�QDVƫ��.c�LTQAC��E�U�LMUU:w0⦊+�f1UT�L�35E����f��q�D�r�MS���5Q�h*(��*j&���6�֌UL�U5DF�rb

�G6M�1E4D�sjh��*���"��X�jI�J�-`�*)&y&� ��4�T\Ƙd��m$�1ETCE�\�QQST�SS%TTT�G6	�v�T�s9���U�����&��fI���"#gRT�Dk3QQUCMMMr1MM0T���D�PSD�C�QPE1ED�c��;���1W�������ϼ+��]�ĳs��t9�MR�ܚ����RB�mj��p� ҧ��^�k�n��t�=U.TY7��=M��w�gF9�r��P?eg}���Ӟ{�-.��!�^������4-Z�L:�ƲokX'�z��W����`OP�no6���0��յ73�{{I�^A����.��mOB��\��Ϗ�;�ھ���;����0�"��1\�d��ʎR��WJ�uG)�ȸ��x!3��D��;05�ݐ���B(d
.��i#��tr'b���k:T�ͬ���É�|�9��l�w���ZD�goC$�C��I���|������O��]|�x��v� �� �9v�Ƥ�g���l�w���#Xc�c$�]ʁ9�?+(�'{�z����$��ɒ�!�Fq��͜eC [:~iw�,�67����T�.�X5R�<N�h]��za^��ߧ"��zO�ga�j���Q��X�5eEÖ��f�f\��O5�$n���A���02lD��ɻ&����k��b4)X�I�0≔��|��K���Ӄ*25��ϒ ��� �w0���r]�Od��ވL���N��Qn�:�z������΋�'5[�-�)���{�� ���`�C)�bo��W�x��6��G�U����c����7�u0]�^W�i+7  ���K�ǧ�Ʒ�e�^7t!jY���Mf�>QJ�P�\f����7Î��]��"�}H��$�U�����޳���ڍ�rR=\cLQ�g]N\m^]�Ύ��� <<���� ��e��مWt�m�?���䉠n�z�޶�7  ��X�!?T�#��Ú�5� �^����or���ǩ�}�R�Փ+��]㛖�^����;�r���*���av�ƭ��U]�����oiR�J��aTrW<�Y�E�Ғ��oM����rݥ��wX'�U��!n3z������>��9���L����Vk(Y�Y�:�,�E�)gO2�S�U��e�Ỗ��U�����8t-�!���LZL�e0ƽ�#�hv��aD���s?_:OMW�5��%�2��/b�ٶr��V��u�P�f!�4����3-��,9�J��Zȼ�k��1C���@�U[�oC�ތp��U�3���:��E����1w�~Ɇd�v��#��mg%��,(���,�v�2�>:��Ϻ���5��0&}��8^]��UW7N5��c��;��of˰W�h<�@$?���D�4��-�o��5cT�n��z��ɱ�f^C�8P{2��z�3��cs ��45�]��i����Ƕ�q��*���br1�A@�_�xsQ�T:1G�K����.薟��=�{��a��pU�n^1��	t��=�j��il}����GGl��yC�e��M��M��f�#�t�cAT[���ڷ���l�2�^H���^�>{���s�^���ϗ�E���C� ����}љ����0���S��C�
X!'�̚OuQ�F­�lk�{Z����P����z�UE�^-�����u[�"cN	����آ�.��KsPǙ�&��r��3�'�wU��ܶ�+6�e
n$Ȟz�(]�^9�A�/�r�Q�̫U�[.�è(�LH�*u�NS��nN��A�Am�1%�ɔ�3��S�]��}�dJ{��v�`��$�]�q��Rκ�epv2��mC:�h;��;�%:�1,���)�JS�\��O	Ϸ��T
���oF3L�B�i��F��z�H�i�_Qw��]0FaH7@ʖ����\�rn�i��5K
�<q(��8t�5�<��D&�	�{
7����Q�]/e�?7y(,n��e��hȓ����Ovέw�C�K��p�����Zc�kuz��ˬַ�k�;Y���*�\��)tڼ��"�f�wD��|�����Jzp���h�aΨr�Q?�OO��P�������U��g���;v�u���O<����{��q<�d�]t[�!�8�� "8��v�L����F+;�4�Ї�����hTф�N�c�A�`�e��c)0��D�6#*�]0wc�����ݧj�*R��\+�5]c��p*��f�V��"�����vv�5X�Y�N�j�D݄dgw�.[����|�Ͼ�}����M���?� ?� � ��c8�J��
�5���[6��3�/Q.+կ`���VvK1�b�;7���1�r�q�[&�Ұ�:u������7d3l�J���C׉��HD[��!��-�Р]�J|�]=jK��0��?0����ŗ=���A���l�t�"I�e�'z�w��ej�
c{Lj��6"���K<�-$d��O[��s_	24{����|�+�d쒝
���L�dj�۱�q���!�Ѐ1%�<�{6��(���K��G���kC몑����n�fYZe�.�\��{6��HcV�&H܇����1��G����,:/1q��yMt_5g%͐էw�0�J��>҄��'�H2k�SI��^�通x.���zaPP6Bضs�*���?Vا+���Xy��VJ�j�D �W���:����d�,�0����L�㺇O?���m��%��Ȼ�P.@���Ba0]� ���])�yF�����O�1�Q���	�%���w.�Z�|���2���?��ki�`6�82��v�2�}%�H�I>9�NU��eTN��]�_�w��\��0`�:~�k�^�	��y����SU��Е����x2�).�L��,7Za�VsRȐ���t뎃aͣ}gw"��1<����o��|������Jh<�tja+Ua�Ik�����2e�����yy-�c�{Jb�<h
Ϯ�3?�U_-�U��P&@�D�< �f o6�%rօ�n��ƫX�_��^��}��
A�9�hL8��5�χ���n�	s1��=�y���O��]{z-?��'������<�-���F�����=�S�fi�u.�*��sް�-�Ě�e?�MZ��a�(�z�g& �v����!��?s����J���E��Φ/T����`K�k��ғ�_��6�a\���6^Ż���ݲ�v"�'�\:��	:���@~�n}�2)��SI�P/�\��N�j��4'���f+Z��:ӑ�ѽ;l�CC�<h�Ŧ[�� ����4���	��
$@:��+��=Y\�n�vMa,�������w�%�dG3�H���l��X���pȋ=�ڐ���0ӯR��b=����ޖ`5�s���O��.�qE���~�sV6/i�ѓI|�w�~}�u���|��&Y�2y�(�A�r2�m�cR|�x5�)�0(F4��Ί�L&fv#��.v� �mי������r��92j	d�մ�@aN�Y���� [:~iw>a�/i)��;;��k�c<47�:��"�bw �<���b�r�dtrā����f�v��(]
��^w�ފ]�3j��Ӕ�R�-�c����Q��F�1X�+ �ϗCH�<�; Fc���������o�ɭ�y��,��M5_�{�{���
B���V��U($]���Ͽ��~����_��M������Ʀ&nG+����PB}k;'�-@c��ߺ`3˰��L�[T�^[��ڵ���������`�DH���q�&'���gY5d���A������*��S�S�oc{sV��@nd�PQp�p����A�k�0����.���Mͽ�'��O'y���}8*��~SO�ȪmU����l'�-�W�q��gd���!��˷~�h�f�5nm��9;	�UԘ��1I�[�I�&A~��f�x`w @AƑB�G���i슗[x׫����,C渆�/�;O�*Jz�L�"� c�|���Msӿ3�knD��wε�E�w���w���2��k�F�i0�9+�Z���^o�IcH�CW� ]��99?~/�R�lx�9�?U

��t�+�<8c�?*�3IuV�f��0�)��ήcX������S�]&F�UfN���5d�\���#��)�`��� Lk�R9��i�j�J�e�W<ES_%��A��g�Dn~W�25	���'[��b0t8G����p؜�ږe��E�1�J5u���.8�4�v?m�R�3�}v �V�k��#f�
|!7�t3�������;�G{��&� ��_mR�������b��8��}(ft���q�o��**`5�RH�+f����yM����D���S��ǎ[IOMp��&��V.5O~�����ER�V%" �ZPF!f__>|���~~���o���f��vh�&����/E�3�2%��D&�o�oy��L8��9s[�� ��⥙HŔX�]��m�$̻H��E���_���\D�[9;t���R�y���^��{aC&�,��",c�i�oúA��T}h�;릳"1�x��G�6�f����wm�C��!�p0&@��$Fd�{Qx�ۯm��Oy�Z�T^�W!
�	�'7�����쳊�#��:�@�ј?T���&
��=%����p�q8�U��9R��=�HZ�7ǥJ������&TAڮ��B�L�8t7�M�T9�k�)�B�9g`��j-�>کnm���E�V��m�{\)lCL�ƭ�����Ӛ��z����v�1{砜Q�逰_m����ằ�+B��>�ˎ�3r��c��RX&�IP�����o	���m�~�SuV���EW'ǉ�˰=��c}���ث��	:�1,��n�cE*L(?Es�w0�CWT�:���*��E+{���p���n��7v4Y}E�GdQt�ѩE��K:a������!���錹\���B�ҩ�EC6�U���yB��p�))` v�ч?R<n�Gh�ý���+�4�m}9ǣz�Y����w[����Q�'^�R�=͗h��zg�����POtV`�!XK���Y�@���kH��ppG�Ͼ��_o�	A�fDRd��))aB��T�5Y�0�C�|�����`P͍0D�p��vp�w�8����Z~n��Ƿ"�sĵ��]�+��lC��d�?k��?�̛���ښ.����t���duB�s�Rƶ:wnw5t�וR�ǣS����zY�@/N���:C�G�:��SM�k�SS�i����l�b�-�)���zW=����W�����L�t��6���N��ʷ0���&/L�f���baInT�z�p>�zfy��K1�Xgc ��mcns�W*sbPt�v���>��d�[��Gd��8�zHz$@:Kϳ�D[��Lc)�^K��y��1��7�mU�#����8��6^��5��h1�����H}�"!�i<�WWP~�w�`�����[�v"���%�=!	-M>C���T�2O^5�h�nݏbvh���ݩ�$5k���`Юuv�*`P	]T�p�z��]��X*�pϡ���/���l;r?O<-$����Wkm���{�~u������l91�,U�RK(>l_>���WH�x��� �����%�8�K_sV�*Tfi�H��8�[��Ť5����}���ǶХWs���x'�>J��ᝌ�u������Jin���[���LK��,I�V޼YԞ���)Y��լF��;4�0���@�A+�WhI��.xjP��v��)�(_�C�"- �"
ҴD��B�J4�(P�̠R ĀR�z9�}�����8n�
�o/D���0��"Sm�L�ɪҚOr��
�1�z���ؽ�x���{�Sks:�j�N�B�,.b��� ��U���'��d_Ji���I��Gc�vLHF�L#�FMv�w�P�.�>����2}�)ٲ��,c@#��tD�I˼'K`Kv�w>��f��vt��i��B2皃�\9���P�m"�m���!�*�.�uI�\�v�:��}���]�
��/"�����9��"FǘE���G��M�1��F��Qzu$��J�Z{r��u�6`�,P���Qi�g�H%�ryA�z���'��G8K�ǘ���H7m[ko���b	��G�W4�~ƹ�l"�GbqC���~�
��}^UL��՗�B���\VR��o��Z��Ћ�>�*T+��,\����)?5��M�*���l�l[�6�0�c��<X�.ok*����o3x�dC���;'%��hv���%0� �k-{����5��_�iS�V��P˨F�k��8���ZD>���e>��ʃ����i���dUTN4m)��/	%K?K�yZ7{�v%}�#ʌ#�?	�����`\t��o�f��h�heeN��P�j�e:]������:�����Y�����|U���mv�	��e3�Y�g>9�[~c��ua�Z7tʬE������6�c�MM�.�>������B�R(�����@ R�(���"���<:tĊؕt����I���c��^ø�xg��9�����X���k%~��м<5̆de��{Z��li�&��x�3%��,�{�m����i�q� D�N����q�Jg+U4M��l��1�f����$�PJm�j�e�}o�i�����P��Z�QN���p�e���h��cB,�ˡUs�67b��a���!MId�ԑ��<oF2�l��/�����ᕧq��+wC�@��^1R�OL".;9mCT�Z��	�8�Z�V3�o'�+f!�UKR��3�:�L=��sW�ƃ�X�N2�'��j�d�2as�� �^�LRuZ1�c"�.n6��&��v��T��I�FϢ�f�ο��\c<�-�Pe��a'i���{%72�2cr����f^ffJ=�i�Q\�J��UE8��l;��o@�DcL:A���U��x��̡���.������}�e�{�Rd��&���D�7p�;�0���F7e�ւ)6sO�0T���~B`X���%�����{*Jz�f�X�2��7|zk�����Ѿ�z�^^����z�z��������������������po�%~�W~�Vc�����D>b̶�շٴ��ҧ�؎̫4�&_3����E�RsvNb-܇�ǣ�;t�^ЊqaYZ��s�0��ǧrх1m���l�����HR��7�Җ ���ʛ�GXν�N�0f9X:��d����cRh���ݨLKN�r?��^y{�Ku��`��Ý����W�ҭ�.�g{
`0^��V�h�IFw�L����{{7sc��l��⹽�R�T����/�S4M�9�+]�u�Gg�+zlX��2s)�:5:;r�qͭ'3nAwrg5�r�<#�e��m0��*A��4]]����n_��v�M]�'kȩK�$N��d�m�����*,.n����Z�# ��ب��ҥ)w��Ւ�������fhةu����8e��g9V���ʤͫ�t�//�y��U+7�'Y��d�5R���F�P����ޔj��X�u�ɷ���9}؈�Q�Җ�O�b&���6Kvt����p�ũ��#�n�'��-�.�����>.��2���r;�j�̈�sLyuE��^��̛�[W�u4۶)���]�qn��GonW:�9C7���ZH��Q������N�Zh]��;��fPQ�4�r\ҫ�^(ӎ�uLU�W�Y�ԍ�uҫ������^��	��Kq�[z�T�՛aC�#q+:]��{QsU�&�,�HO�a؜N_t�fWw��Y	�m�ζ(�X�w	3��YK�'�;�.�������Ć�]��X�-�O��=�S�t��N��?s�����`��N�x���Ǝ'/���Urkс�%�x}��jk��w6
��uX4��i��w�pMRa\�@n�k�S�|��F-��E���v�К���u���ؽF����l�����Jwԅ<������b�1)u펧��z)�M�OnӺ�D.�ni�f���7O� �k�v����Ǳ�/8J��mm�nR�	��M�����q%2�i2�c�-�훯HN��.��vK���g:5��:ž���E\�p�hxx��],��%uŝ��!]��YϦ&�ze�98ͭum�B�wjn���x�&f9Yp˖�Gw�U�a��5��N���gS]rR�FJ{Q��Gvo
Ky���MD�霵{5�4w�tb�Go�Y�M6��%z0���O<&�;�aR��U�Y:�a�����V��ޗ�Gsh�壉陥z%#�t����<�1��Mќ�Vq���2�Z:��|8��&��\���Ex)=�HJ�S��a����r�꾵�YѻK�:b\��Wl���>Me��E!�+2��fm���K�hE�j��`h�Ɩ��Cy�[��[o'���u%��!���nS�&�EV�f�ҩ���C�K-�G���T_<���4�K��w��`�ϕ�Ī�ٽ*S9\j�R;��]5m�gv��S��6CD�7�2b;y�b+�����#}��M]���~��T�%U1DD���C��0DES�514UA4� ���֍�͒����*�����	��tP��[h�]�ICPP��E%�Q��mCUTQTD�5Q33T�QL5ITM1554D�R�DU�T�$ETE������ �"b
*��<ܞU@D�UC�N�ґ6�DIM4Ҕ55�1S��4��-(������fJ(������X���"�(���� ����(�������)h�-1@P�U�SICQK�U!BRQEET��km���h�
��U5KM&ک*�(�����)!I���
48��~�������ߝ�~#=ezm BTz*E��{�u�Z�����x
���Fa|,=��̻����Jovۥ�҆�޿�W�_ϯ��①h@����	!�D�d&UX*Z��s[5��B����!�1�yO��hQ��4�U�����/6��(��3*ڿ3�ii�|����K����8<6�	oCM��7Ψ�tf�Q�bN���,)gO2��ѩْs�~����C:�k�!�ue���ʷqU]r�~���{C�е~Q+\r�$*Ol���zb��/���ӡ�	=���؝nj����#��k�T�潵,�Vj��u�^����Wl�wΫ�6v�2�����#��ʞ�!��;�Vx�@�ʑ/���4Bo��̗R�9A��������ۃ���.~g�F��7��{�g����!��X�ʬZY2�V�AQ���>j�#f�u�BPB9<�ξ0��s�NoS��yC�tC���^D�4�l��w0ה͎�^�i���˥�����E�#2R{��Ƕ�7cFd���H/
�!����;U��u[��l�/5�S�.��u�,���E�IāsE�1��<㊦��JB��/,��l,���z�y�_�(��Z��p��Ɋ�5�MމBSkH&H3a�s� z����_L���~Q_J�M1q)��j�č���C�4�`���M�r�ˡ:�S*�-N�����oicQ��_,�~�鮗^\���)f�����c뺐)�z��oE�5GQ���U��%8�9y�f�D�!K;�<8�T�Էλ(��N��{���J��מ���!�ҀD�P�P�ҒJD�R!HT���ߞ|�K�6��Sk~)��HL��CG(Y�}�o>��v�[HN$��Z��5�,C���Q���{�O��P~"S^��RZY��!%B�F�c���|�:���۟�k<n���Yˡ�����e/~�08s��hOa�N��N�xd� �ƼR�¼�Ͼc۱�f���`�%���D��d$l3d���s�ݝ�"U��}�E�F�X��l��y}q6�a�G��ɷ��؈v@��c>�'fƸ���`&��>ta��(➗�.�;slL�TM�Ӟ�9o��(,kڥ;�&��\>h!y��;kP�5��������u�j�B�IyNn��>����xC��J^����B�r	a���2ONd����\�r�?����D�S�����l2��͖�Uk[
q��=+�ʂ^���>�[���])�W*?l������V�YB:�_�!�^�aٷ ��7�1��+L��:��ǧӯD���f%�3�yې�{E��������!�y���B1<��|Ocj?V�m�_��zHz$@;D�x���
��5(�W���bkT�w$�#Mk)��|*��z5���Yó�/t�R1�}.���Xg;����Q0=+})�."��N<ȶQ�̌��(�z��nK����8�Y��8#�1�ɵ!I�Oh���ꖨ�!ڳ��b���%�"�X�ϩ��QH)R*�!J�H��J�P+H�@z�>���m������_0���|*�;
%�r����DJ�/�����4��0v��$<�|�eE�LM2��}0�Bӵ%�[�@؊�42%����I������?eE��`焝CX¯�������ǒ�ا�ut�R]�Ƚ�O@sͼ4�u�x�塯�&||�;A�8��p�j]���N����JTͶvPej-�mH�����cM<,��`qm%v���2�u1�s�C���ة����yM�(2j������
��Fcս[�y�����b�F�E�)�g�"�\� .#V�"�J�j�N(�yFz�ebR��mx�.}�g�تNв�:ɋU���><�On�$t�bK�e	��p��'�}��[��N/LOA��4�|U�Ɵ�ց�kk���ȸu]x��Д�mLpe>�`���]�ǆ��O�Ǣr���͗��Wn��'K=�"�-�Ú�F�>G�e�[!��Bm���=����S5��loq��u��4�������R	z����j�G8~��l�@F����:�eV�N��/�S�ط�P&��-.�	�^z�Z��:����,�NT�-��q�)�u�Qi��ix����f��t�XU} �[E�i���8��trm�b���ػn!�m� do@���ƕ��f.��f*�e Ai��U�!�������$�P� �F�E�Hd(@#|��Ͻ���9����z{��[1��M1�g泰��(�K��,�ד$-X�������$|���r����GX�;��ݚܝ��P5"�Ђk�R~kL���Z��U,����Vѧ�#�Q���ٺ݃.Xpd���]�:����MV�S-��e������?�KE��h��52L3d��=��?]t�B�"��:
�/ѫ��c��Gk��pb܈�d����e�__+�R�f���y��r����{������x�X�f�S�@鶉YV�3��۹=]]������ڏP�f��0�[I�$�~3���>�L�_���o�k�_����׻��׍j������i����JY��t��@%6�5F]���֞�����uYL��i���i��Li?Xd"���aqm��j<�{v&ڀ�	B���JI�z���Z����to4j�k�G��ԁg�J��X�qh�*Sw ������'���ը�%�8���sP5�|��v^b�|{��C*.P�����"K���v�S��!�>��A��y��}�y8�sj`��ȟ���W��#��b�qhE�s�����N���1�Ihּ�Ao�ɞ�!u�)o_�Zq��5<��I�η-K�|����k7��L-�;7n�)��GVy�t��8�k���i��_+�S����8�U��v�U�ϫ��]]�BС0�ĂJ��~|�ƽ�k�E8�1���&��8���\c<H���Р�5��N�7%ہ̱/���51��w[O��smSk%Ysڈ���T-XUE8���a#�-�W�q��i�:A�:��	��GU�;�ۃ^�v��4�g��LU�H���4��.�B�n*y��^��8�+S2˺�~���[���!9�݂�Ӵ�T��LS"�09�B��:���?Q]�`<�@��7��6 y�]8t�a�ב�w=	yO����F��aG!��j��	Ibhd6rk���~ֆaCS]�����_��.��#>1�&�	���q6��K���������c�VT�.O���;�_�d��p��4U}�~����ni�a1�ͺi�k���꾇��(��k=�'�E8��y�'K�QlЍnj�����38#c�}�9败�E˵���!�
�5�ʵ�k:�i�k^�0�;@����0���d$�}A��Ntal���"�Z#�1TA��gz_W���K�����9E�(���^����HG���U`��¾}e�>����[',̓ ��9t�>Y��M���⾴�2��`Y�_�yю����H�H��8U����%p7�n�^����q�Y"i	��R��͢+�J��t3�Z#^��ˬm#�+�#��Ƒ����ho �2��~ĴfwT�w;����F�Z4d�5ܯ�UW��
@�
P>{���<������s��m�t	�b3_}%��{��Yv�N�=yC�tC�*!0���:-�a5��<U�`y?o=U���;(l�� r�Sz����ت�Ƕ��Ƒ����� �),�a&c�6�M=��EwfH`���+��M]1p�)�,"ä�3"���-�o��b[@�]ٜٛ�0����C��$��͋a�1P�XK3��@�0Z@���6�{���;�=��/�o.j�3��@G!)�(ʗH��Q�a�Nk�M<4�3�>�81m7�J�eKm�;M^��i��:���w+�4�)�nBbS�	I`��$�]���z���D��4�2Z��̤���m�E܆�u�|!�	�v1��}����K��ƼR��y19�[�;��;q�z��J�p�\�:mh	ٯ@�L=	r�*�.�o%��z�S3It��쎻6����h5J��b\˖f���
��8Bn�	�;
60�w�ϯ�؞��8.3u�&�>a8-�L�ދO�eAcCT�~j8������@`鵟��v���|���GBf����^O��w�]�:�z����>U��)�:�� ����B���oR�p��}QwSז�]>|k4Q��X�w6��Fg�^I)Վ�U�6R�� P�H��Y1�*�����r�P����/��lҫQmHw������z��~r���+�-�_�4(�7� 3���B��R��8�вT�zO��W���z s�^܀��l:= �+��̻ m���k�Y��=#SM�̦�\�V��=+�ʂ^��+�i
�Y��-����3b;]?'���\^�Y�� �g�t!��}�ێ��2˼eRc~OO��gӯ@��j�Y��rj�D������{>�P_�* �b����HZ�_ P����m��(�A�� ��P:��Q�<���Ұ���X���[�GX�n�tK�XW��bT�{ڌ�I���2q��|f��/q�c~�Zl��\D5�_F?��a��%�-�9m�=�O���G�l�ζ�m]�-}�!��L�f�*�!B98�#F=w��.�KU].:�_��M�����0f�_C+��]��*���׻&m�x�g���U��	��6->��E[ʰ:E;��zŋC�D��ͦ|�t�͡d����o�BǤ�0F��W�{|E&�=�6J�O�Q�a^=����pf[p�Ʈ�|�e��k�~	�^��	� �*����I�d]#������c"j�},��)�$��=�SM�\��)�Ԭ��1���wN��?l��v��T�
�$h(�Ԯ[Ճz9<�c�Jx�6;~��Y��| ,����ܤx�]R��c(�d�l�ZM��v�Z���z�l�%b�Xoqa���m���2�f�N�^�� 7���-��vU����{��֦~�=�Ǥ�6���۠L&��냯^�t�'I�f�#��1Vz�Uen����2)��4���u�5>Eêq �5��R͵1����v:w�ٍg��
����ֺNF�w�WR.��9H{�E*h��х���찋a#��Bm�6\�Dh��Y���v��Қ��T�O�Bn��LZ~XH%�'�܌�	=�CE�5�M�����>�����xo�s!F8�lķk�VM7X��r�ge�P5�?$w=X�8�;��N"S՜�Q{;�^9h�2Ϙ>�1~8:����:����l�5V��&y?5�2[��j�Ы�6�ꪛXef*l����*S7!ю��]�pna�A���v�E�uCs�v���aşfz6B�����So���N��ݱK�k�QI��`H������73������!����d�C��~=Pps�mf�6S���k����
_��|x�a�x�&�q@������x10���N�J��F��!�"�V9�Ʈ^*�'�װ؛&h�P�,Ť�0�|tE���6�kdK� �|�֣���.oX��z�6���4�z��ٚ�ms�#F/V�Cb@�2+��;ծ�V�h��x�&�m��P�F�+%`����1:���n��eBb�t�4�l�	y �`�18^ɻ�f.w�U�c���)f6�H�y]�_ʯ��ti�<Qtw��T��8�n�z}2�3E�<�EM�^�e��Z��E<}�
0fGN��;wywZ:���ا�U\����V5P�q�\B�M��3��Há��{W^t>�,�PҺ���J��U�����9�
�7n��x���U�B�[��	�e�wUm�kP��U��-�Nͳ���C*.ۆk�
͈��*by�uN�jɅ�p�jO`��2��>k3�z��sg��L,%�]��C�.[�>zD�Y�'n�7���ug[�9���s�;PDη5tBd������J��UE8��.�;"��oD�#�
��mo><J<��A�}�.�5�l�ԩ2�0G������@����O.�FN���58WwB�24F4Ж4s�L9�v@�U�|@�nɂ��6Ⱥ�09�iy3wZ��hO��֯�r�������bm���#���t�Ou�hQ���
9�[���^{��$c5���-�E��['�wvm�{|d0r�17��Ό܊:bN���s����s�'҆�YҶ,5���">�Mz��9�Y��Dd�v�kBޝ���F�¹��Q�m=���ʘ�K~{�1=IvsJ��2ZX���z-Jc�9�ɜ�6�1����&&`�܄��4o��偻n��T}�՜����1aȎ(�<w����*���x��͹8U�)az`�W�]k	�{��%q�Ei�@ר��B��W���j�j��M�q���
�Ξ��� �N�V��r���R���'Z�=��Gs��|�%z�p\;�t�p�����O�y���8'P��m4�o���a?Mk߉�iڢ\]75�P0���d�W�eޗvͲxǙ��άB��sw�syR̋��t�t�Qa@���@�f�z ��i:"��9���"ԑ�/q��Ѽ���)�� ѐ&tF'��%����#��S��Ȳ�^�Hz*��16����������tl{��e�@_Օ�NBe��BO�Qx���َHxe��'�t���ֹԷ�P.�W#E�y���7"���r`���K耥���ߌ��ɲܝ8���s>?nXiۧcۧ#a[K.FB׵��*�P�iQ���.b��lS<!	���jxŃ�U̴Ҹ���ލ�j��m���KsP~"Sm�d&T-�£�.�Nk�=[�M=��}�]-v���	�|W}<%S �N>C�# ��|����������RX&�zT�k��ϛ������_�ׯ���������ϻ��}���7����n��=u��˖Uՙl�Dvݩǲ�+f�<�����9�$�ͺ���#Mp�݊���.�\�9!�����(�M�>�N�m���%{Z�j�Z�*�ۺ$�J�V�:퓍���x�����[W���9�����8�����#=ʋ��o��b��N�����T�7�,{�#{�v�%�/m���X8��+���uk�2�];�ŎB�:Q,��X-9��ʗ���t��-��j�3v(s\0�}ȥ+,%nr�x�ڧi�
�:5Zn�n��<�K
��i�gWg0�s��mp��Rl�Ү�#�RmJ�nr�u��#��q�\�*��ĭ�jA<x^$\���K�P̩�h.DZ��s6�']�8c��܂����w	��.���;م,VG��gv�5��<Yͫ�����9�nf����t���*cD]X
��07R����DB8�2�mi�;�,+�]$r�M:��K�b�9���Eln�]��f|^l��f���v3�ͮڐaD�+%K5%W��Y4��"<�.k�(��;��c�d�1�j4�n�1b[ټ��CGH1ҏj���a#N6�n��Y��˜qn�H2y!ov1�_W"�[0�S�{�cߥo<ʍ���s���&iU����R�{*3`Nl��ͳ���ae��-!Z���L'�*WVە���*@jM�#R�V�
3e7���]��諆$�Z��ЩjI�WC�yJp%}�P�{��}�<c��F%nX�2ZW���;2��+��x�O�X�u����b��G}%Nˬ7A\�;�p�9}�u�I��A) ��j� + [{���I��JT�=~Ű�����iaY|�P�8�,��CfMe�_<h$�4�R��+�,s;�50�2�R�]�_ѵ�"%]u�WX*��+�R���P��i@����r5s�+���M����iW�����<��"ܾ\��[Q��л�Nwe�������54��췵��BO K/��F�ٸ(����_\��V�ta[��EH�k*n�.0�SH�}yKe\��NV�P����k7��*w��9N���d�Z���*�'U��=:ڞ��ݔ�X}1`Ӈ�]Nۥ�3J](��df��g�e5�8Х2��oq:ukU��2��d�/�����j��(�$Hkk��5����@�	����Z�넴/���ar�5nq�V��0�j7%>��m����qR�i�ԩ)����@f�I� ����ȱ̜+Wd�����b��O�spݸ�����feaWDxS��c�?��u㽹 ��R{��v@�3��x��=�`R�-Hb�b���� F>�[��o�����|�x�}R�V(���Rm���m�G9uqTv;���~�s�Jgu�I<��=�/5�]l�g^ �諉�9���y.W]��3��P�@<n�m�ֹw٘�r�f҄�+���ʺ7#��u�F�s�v
��iA	A�Ze0�#I��$���G+Wz������ׯE4R���DAM)�(�
(h���� �4:֠�
(������i��4��F�$ј(���H��!j�
��!����
h1L$B�5MQTP�QEL4PREKKET�R�E QLM0IM%MRQE5TR�l�)j��c%,˶��tQQU1%AM@L�Rе@���ER�4UUS1IIQKCMQU�EQDM2D@DQAT�嚊���*����(��&�*d��媉i��(���������H�xl�	I��E4O6}cSG!�4D�4��E1HSTL�1@R1,IL�U@Q��H��=Hb�g�b(*�C4PR�EPSLLC������ϼ}wϟ�����ӹw4�V�Y)�Zae���Vn�Iٷ����A��G���rR�Q̝�J��]L���T���"��>�����/w=�Qt3����k�!Ŵ��>T�!<�4'ð׷��)<�c�:��0B�#�Y^Iʴg�{W0OqZ����5��B�l>�3=x�`� v4�J��.���0�R�ٌ����=P�.n�I��ӳ��]������0��9�;�g{󇦀��li�����:�Ο�@��xS��� ��?-0�5{R�/A�8�W�P[hj���^�+@ϣ����u]g�s�Ww��ʓ&��m�~���������hfyʣ/V����WC��,��>/N=��!ÅVv�G�ʣu�6�������:��4گ�TZ�Z�[�qc��]�kd��{��\.������{a˹�W8W�o[���r.���@�d�Cv�|�6�̪Ll'����"�կ~&fڬ���u�E��<a�3�+�T&n^1���F�fx���ϡ��'���ݒ����I}�u�`[;S�Xw��R��I����a�[�󡷺�������X�e=�9aC��^�������A�u?�i��p�Z���Pt=B8�v�_E��lEC�xdK:Z���' ����x�-D͙�����ȶΪ����[�I������pպH@�v*�f#��^�h�/s�!gwpF?f+����ʍ��L/�뮋���qu���s�NgPu��1�sEmi�seI1v�1���!X�rv����4-�`���3{EA��o׏{�*���w3E�,��9Iw7�i���o#^Y��#�Y�1'�Zݛ��f.�I��G(gǩr�ۊ�;׷&m�o%L�`�Z�`�.�Fl�z�u�t��ڹ��U�Ǩ�B��0ư�΢���&�������N��l(2j�ʭ>J��G[�EuMo�.���n+�1n�ռ�[�h02F�1����������E���-�x	3%�/�rs�7�_��H�a������%}t`d����Ba0S��#�0��Tj��e(;]m>����Y������u�%:]X�(�kk�����ty��a��@���jc�-��o�@�M��f��fp��0w'a�c]�&�$��'+<�T��j���y�Z-�?���q�n��e֫�B��S{k�y�=�Sq�t��b���k����D��p���n"��Qf^E_pG9�)a�����1,��&���ʹ���/5�R5�=%�^e�㹎�]�zwfg�ڭ-��ݾ��<�����<÷�ǦD����S&m�;�'水ɷ��FV��t"Y�)kc{uw+��ُ���1��^d>=�n��YQ[�f��}V7kf����l3�����V!V�?^��G��d�9bcx�k]y�[QD̙��彻Z�r�U�q��׊�5����A�3��C9
w�:Rx��F��)G�4�˿��W��wn�}-{������r�͆����~/>�mt^�����MW��tu��	��&J��O�5�yk�T�Ӭ�>��j�������63�����Ť}l/Cj>�8=u�V�[Y�C�*�p����
�h%��a��]X|<R��V��B����__��K����k�>��nE����a�]����j�1b\Ã��sͼdY/}�.u~cg���L���Ys�i:���Yz&7�_T�m����0��������b�����M�]� �'�'�����[��G������u	��=K#qg���U\��vm�b���!,�\������ϝ�~���y0�)~VgPmC f0xO@��銀�l�h��|Ǧ ������O��&��훺7���ݍb��T�q�%Ռ�v>6K�9��P.lD�Bby�@�:ɟ�]9�Q�����u�mU��A��ܢ����O����W�����?��r�$��N��v�5�z��-��w�tGF��W.˺]�N����{1�_�J��RS����;"�F7��<�,���Wv-�6q�播�}kT&�Aۢ�M���k{�5]�n$m�U}�S2�*���F�1Qr^��n+�������}\��ceS6���]��VQn���|j(e�j-�ْ
�g^�HG�0�%l�|%Y�zz����l���t��Q�_���o �em�&�C����n]�i�ޖm�R�w��LP�].�`�S�`�
�jP�=��yy1(4>5Ð����'�ĊeyƝ�v�����y�c��88�M2֯dmF�[�ײ����t!�oM�}g�8{hA�ןC���R����hQ�)����,t����TY�y��OVoW�IcH�C_��ywf�p^Ç��!�8�Ƅ@����ά�b��.o��&�h���ݾ��t����I��<ʕN�-T���n5�!��ͭ͂�LTR���l9��1vU؅�NvP�F%k�a?J�T��G0�v��P���:�nƇ�=aM�oȴ]�����>ۚ�n��Ø�R
m���@Y�hh�U�U�/�P>��D����X*�ڵ��^�w#:�� x�nleK1N��Y�I`K�=y�&����̻N����^T��z
�o媿!ߪ�T�hw��@��_D<��d�x����H��O4;dgJ��v.2)[��M���CC.;0�tE�����U�^gh	A��Fd��U�m~݌j _�{W�K�c�Z���Vٕ�y��͔q�����G���j�6|͚D�mΗ�LmgH��ntP���IWJ���#yk�Z�1i�>���!AG0��V�Q��>:�ͷ�V遌Q.}ՠ���H%ȇM�Z���d],aKE �+�_�ռ&�OK���,kn>�-e�c��B��>�M�j鋇U]6� `��M����y� ���"TQ���:w�ysV)U-mG���gaUk(RJN8|ض.b���=�	��M�r1�҅�]��O�F�g`��ǖ�Ks7!	�A2*�j<Ԟ՝�vNk�z��Q�UQP,�ı��W2d��c�/���Hh��,�-]Jca�Jsa)LP��@�)V��Mv
��u���(�>�8���{w��\��^����R���L�M��������d�`Y�uv�gNk@����bˊw0�����3c�`��n�h����s��`���ǉ����.���6�AnM�,hvuC*0i�Pw����������7����(���Ѭry�{�	�MqT*�z9���PX֩N�ԜK�{���=�d��2i�f�9B�D��^FU����WW�4���xOo�?��*�2��%�ں�@,��%��ǆ���흕S:�#lfQak�?�p�\�ښm3�E��$ޝa ���a�T������,_�ƫ��[�r���Y��Y�kx�v����87[��ke��73G֌���U[��o��mF�XwzW��|Z�����x�~�������Р�;�P̮[�.gA5i3C�f��7܃666��j�x���]�$u:�W(W�N@����&�	|�Z�{�3=�l��弄�޹�~�Ey�!ٷ7:m��ʤ���S����u�z�Q�c*�M�y�;��.�k.̖cTY�	`�ȸf�����:�_e�?f@f�����wb9%U��B|F>V�vJ�k��aS~<��X�c=�A���Se��Q����^��.�u�m��R`��Hq��j|_E��lEC�dK<!���-6NA0�M; o_�o��x�׽���7qS4P�X�B��Ñ{6���xiזy.OuTw~
��.Y��v�B�醑O���d��3m�)f�eU�jq�j	��3g�]C���۽��&35;Ƿ|�<�@�t88���ȋ������	Xڊ��%6�2ciM'n�<���<?*��*�u$r?ϒ��5�\OV�� ��"X\�Cέ�Ed��?B	�:i}��r�o�΅-E�Ji��R��q���xgO4�� ��
$�6P�L�4�&��١�͉�r��.g(�9��ݵZ��"y�|Bw�����LJR����y���ty�n��P��Y��������߶�F�`�q��������Ǹ�����{�����n����ص%uM�t�P�\�v՜u([́����OEʄ�=�m�ӂ��7b�f�ޗ�["��:FKh(X�hW�1����;I�V=�f�G_6tNv��]�M��q#��i'��)9X9�R��XsQ����>�,(���$Z�2�Y����}M�����Qs�!������ŧ�\�*GR3LlD�I��E��}��g���0�-0�s��p��eϝW4�y����"�E������gm�S��z�;�Ymv��������� ���0~��P�d�h�άԊcB	�k��I���o�I�H[��鬝-�aƬ��7>�U5@d�C�u�P�C�:��h�?�y������L9��-�]���(Z�pz�0��x�:�.�W�b�A�èC�H�`���tŝ����]�?b����1���MoKܶ�� �$��Nf�P$@;D�px�a��tMN(��_�o���O�ǊR9�I�����~M]��>u�߽S�yÆ��&h�ŴHDYz����5�.���i��cUb{�U��;�C��Q`(���w�O�{>޿�L�`'�'����A���dQ�n�,:�Z*2������s��&ivV�u	U�ʛ��K{d^f���7kF(H8���y���S�[�
��7�vBq4��8ݪN��Z��\�Rj����r��V
�`YN��4&.w_+l��K6�E��ܫ/�UԠ����X�ܭ0����b�;�S4�б+{ {��Ԩ#�����J�����u���{�x�u{��v���l1{|��X�=8�^͜�ت��u���ʱ�/ߋ�fm��<�_a�<�Q, ?M��9��2����C-K���`��d�C����(a�����ܣO�@�{�Ȯ����W0'�0C-r^S��Хr�0���N7C�:��|�-�&�4;r&Y���!�L�v�f�&/�r]���M�]�'�b%:�$�Z�J����$ΰ��m	���2�B��0l�,^E���F4�|!Ĉt�����4����F�*L���Xn�k/c��Pc6�oy��)�t�*9ٍ<0�`���B�0�'�s�8�U�]�vT��`��E�C�ܳm�3��wiƻ]�Ъ��]��	�}�3�ˇ�� �kȇ!���S��uF��I�l����e�*�7��1�2����'�l�,k��C	<;�@��><������D�^���Ҫ��$�cV��R5��=�K<����*�
��̥Tzu�����\a��Р}GG]
:8+�~	xjSi��}Ö5"*F1:�R�V���~��eA/maTs	���r�`�4T+>5�I�}@��o� $��6+�El���ץ����'n�M�ew�f�,ũ��Y�Q,��x8�
p��^��y�����T��Q���NX��뒞�iͤ W�L�WyD���=�� ���kn�])R
F�;W>"�/(sr�k僩���(�[��+�G>�^fH(����6���q��u*�����vh� ������h9	�'%\O��x�g�*D���^ ���o�2��']����9E�bK�x�f�x��s
6n% �`wI�==�x����r�@�~y^]�."�F�)�{f���"�,��3<�Qz�y�a�����B�tL��l�:"�s�<1�63�1�޻NӉ���N;�s��f���'�|v�rn���yE
���f��B����m�WL\:��g�XE�IƇ�V���x�w]�+�|3�t~��ۥWߪ�u��1bozB׳��*���J�Tu����	��T9��gZs��ѵ�8r韫��ke�&5���j͜b�����D��`&DZ4)=�9B�?���6=�V*�'Y\Փ��=r2��k�;@�b�BP*(L���!���O5�%1�1)�P�&tF���}^O5���v���S�V~�Z����5��aM�:A�0O#��=��;�):�-����r��l��M4k	ޅ-Z�1M�J�
~���a=}h��2�"�R�7v4Q���~�]���C�0M�l��cJkTgS%,������4p��/����/��N�{���&����=$[���Z;:�`�5
�Ā�Ζs*q��MJ�ydNrU�ԩk��O]�6H�l
B�|�nTr�����V�5���f�3M=v�cs�5:4c�,��O�`L/�T��<�ʇ����9jw��Q�w֯GLu#�2'q�/��,�-�o*mF������)�~9���J�;�Rq.���C�u�F%Ϫ{�^�����;���u�-��O:��`Z�Ӵ,�&\�Q��m]�X�|^�<��"bJ}������h8@p�ar�c�� ��{ji�t�je�J�aD��t��	��.�.T�a�<!{��>8�OAf��l'ä0g:������l�6c��M��*���i|��NŽ�g��խ�k�N��MGrY��������x!�!�_��2~��!�sK�E��z������:����r�1��`���b��!��úXf����E�lZTC�k�0���a�*;�c��1�v����`���D$j|_j���J#��:�=�dt�g�_����سg��9�w�Rw�����_I`J�r�wo3�ٴ��y������	m�۸����>�2��6]�FFS��}<�7&m�jJ����A�S���7!�?���������>>?���������'����=26X���C�h��q-"���Y�����z�V}�ȭp��8˥K���+�]�X�l�kip0	|4'[��t��^P��Qܺr�fֻv_V��P2K����R����8l`La�U�9��&Wm�cNʎ�Q��Jm�Ճ�N�d�u��a=�nV���IeZ5���;Clu=�UwTX�Z��E���D`��iH��� [`CǹҤ66��p�u��T���i`�4K&�路w�&��1��ˍ�:�1+S��L�ܙ�Ie��Fm��)�p�l�&�-ɐ�}漭���n�j��9e���Z�5ـ/�gj�%�����0���%V��P��:�ޙ�`W8��� ,��R�;`�r�)IE��(Lέ�Fe�9��i[�h%�iNo��s���l`�a��e�.V������t݉�b����a�+�G{=SےW]�Ȱ�U�������闸���%P��&�t���4��wX
`P�Y;b��z�V�s��;3Aye��/>Yc)T',H����\_��,�㙵����y�K�2,k7�I�2ke��\�+U^��[MHּ��6���p�ɘ�@�VHȇ.&~j�C��Q��)vʦα�-Y'_-o4������b����b�l�+�I٪�N�\�%���~k�C)�ԋ���w�:wB��_n�#L��ƽ���vV��r�fѫ�� �`�����&y�kc{�պ�.��,u�m�P]���y��;�ֹ����iT��fX6��'Y�5vr[)�N�pn��=w�KV�|�J���+��e��2��)��]w6c���T�S��lr�L��ɓg](��ҍ����O��ܕy�%�!�F������
�
|�ر$�^-U��Y����9j���2����YfM�8�.�k�8}���T�N��a�;oc��˽�;�:h��ȴ�D�5���k��jp[�P�F˦�ˮ�p�5�)��ehI=�GJz�S�����c6u�(��k����e�Ck7qbx1�͒������lE|���Ӱ�Ԥ�9�ljq��m�&��w�1�ջ[o4B�`a��>����{���N�[&�P�;X�I��U�+�zabq�WU�.�닔����Z���{ -7}�v��	�U���{��ދݠ�;[X��Y:r�N�6�o;�C�� V�����D�%��/v#���_Vi	ٜ¶^L]��v�ק{8{Ex�D�8���
^n��������T�+�n^�J�U�=�{)�\��Ժs��2;��p�SBcNꄢp�z����3)Jo;,gV�j�q��+�k!8M[�6.���`I��,����g��R5�V�g0#(�.�3��<�*��RĴu̼n^ڭF3,�8��x��]�Yq��Z�dZ.�ʂ����9+	4�0:��f�B&��^��B�ɣ��O>�����_U�v8�D��.((\l$��~~�$�E5LE@R�R�T�_rj�iB$���("h����i�)"
()��ւ���[����h(њ��#cJ��.�!B{�17h�&���=sRQT���QER�-,O���E��R��4�UԵRPEKM,HEM5T�SA�C�b*��%S@QKIEE%QLA���� ���N���e(H��"����� �)b*���(&��
JhZ4R"�"��`�R��B�퀉Қh�u���DHS��UAMC��Z4�%LLHD�V�*��uM���	l��A�i�h)(�h�E6���?}�������w�|���iQ�ru3S#Մ�B�Ewմ���$����$�K3��!.����f�IN�6��x�q�[�v�3�^L�
�,����BW�F�+��ū_>��X�+Q^�"f�2�&g�g���|��s]V�_h�Ӽ�Q�aAtf=zޭ�=|w��`�as�Hyղ�S��7��{�~&�\��ܠK�/��tQ�d����
F�a����0���d���^�L�ia�Ŕ�غЖw1�����:N)ծ�Lk�Mmq�<͏P�:<�3[l���\�▯_C�ވz�w�ߩ3r{!�,���v�H�I>1I���"��Xs/#���~Ŝ4cL�v|ָhWڡ��=�G7W�m��<Ԟ��0�n�S����P;���vn>l�F��Y�*���އ�P�x�2E��kH�#�H�>�d_l���k����Z��aˆ�hl�j ����t��B��K���V.���M�� �����F���ѿ����D<o��H�8�V�;�'8�UOL�r�oV���`d�VH�
�xR�Q�^b��I̻�VՄ˩�7��E�uZ���S@�k-{�'���j���z���H�:)h�+�R�<*�����o"Ot=�,��9��5:u+��P�J���h� �����)�=�2�X���1q�%�Nmd��v�Ӕ���m�'a�
�d�&�蟃��BT�T@��ʠ]]�(�uק��:����6;�t�ז<�M@c�0TJ��TX��=>ݮӹL�P�^�l������U�w=�j��������x�$��	��
�Iy����-^/a�G<3���C���]��Vю����	����2���X���	�4]��bĿC�tE�@ֻ��z�Тl@�����j_�N͎fgu��Hd�~�H��ZE�k���tŶӞ�ޟFe�f��yڊ�dWs��z�1J�Q'���^����x��ȧx�(>0���E�U\����cO�BA�uMr
�Y��UP��{{_�-��/g�b�n@�t��zw�X02}�y��zaS7 ��K�0/�빽�Kd�J�C��Z��A=Z�,�%Ռ����=�h\gA@�"K��"�!�т;�un��uv��e�3��C&;����^�LRu`b4)_�RaMK�q�uEê��ƾ��a���J���
[���5�Ɨm�v#�kw�!2O`�Jua%B��Ҩ���Q���Ի�������%l�z�Bu���ro�%ۃH��v��T�`c1C�I~��qv�U��W�z��P���vk��n@�B�#��'�s��%�_v��RS�z|�nٻ��,��!��Z���:uW(�Yu�!6��C��x阦�=��;l]Z,�;$�Z�rM�V)h�Ym��g���ܮ&s�� $Xe5B��NA�0\yy�*v�R:�h�c%;<�n5{�2n��5�3�S`�sYW[�:��J�k$$���gl�H]-�(ZWNN����X׏�1�i���4�O>�~g�8{l�>C�Ľ	yS�R�Frg<�N�����Ũ�5R��U��^m),i�a)�ݚ7#=���>��s�M��K׳�"�l��ΆUڻѬ�d�,qZ*�O����e*��&�|n�\0g�A���j�w�}i��w������3�zb��sm�BՂ��\qn��߄����r]y��j��<އm��!s�ңY����e"�4�r]Pږe���,9��T��{�ӵ�MKs��Z"_M'���z�](G: ��}�"]む�0��o�0̓�;����Qa^&$�E3�K�@TYv2~im�<t��O�l?��!�ұҹU��֊@�_�ʜ���S�
78�緩�?�trǳjtm�^�+��h~.d3t=2�xc�g���(>���Nu��s�]sνX9f����-�īC�_9����r5��t������с�
"�lԽ4�%.�V���ÅsI�1���K[V�κ�\�(%G\=��W-4|>_���g�&~��=|7c�]��1.k�N����v_a؛6c��]�H��Ȑ|���C^�Ǵt�>�
b�`|�!����gj�j�n�X/���Pҳ1�0�c*K)H�#ƴ��1u(4��h�N#G�re��pe���z, u$��Qܭ�{�SkN	��#���2Y3��D&�2*�hR{
�T�;\.��9�!ʍ�v�f�鷭YSd�ʋz�xe���u��GF����|�	�ex��_)殄&�����k� A��*�2�8�Aޡo�v��o	��
n.�|��B~�pGY�s��c��9vq��SO�Q,���LJR�6��{����`�XP��"1��Թ�ޤ�m�:��&­,w���C�k��E'L�E�·l�.��:�.g��N�	(�aW�����c~���z�T�ڹ�k���i�8����)a��'��]/G"��ZPX֩N���w�;`>���[���a��� �tvC3�^�6���X�ښN�Ƨ�;B�W�Q���J���@��k=:˳2P��Ӫ:���<�a��G�8u�յ4�j�uQkd�N0�OJװ��OOg���ˎ�����l�l���6Pض��0n��!^a�]4��6���M��*��C+�z��ng���4��<�7���.j�c��x'Y�,ƶ,3��`38�`<��E��d~<>�<0
/ػ��m8|纠�f���/DU'w��f��SԒ[�f�8X�B��ΚX+�$3�]�`�OiPXb`���4)Ľzt�=K7�
��}�����q���Q�G.f[�W�C{9Q#u��q�F@3���s!q��F^�6���_��>����Ϥw���Ѐv�	��tE�x�t�v3�w��3y�K��g�vQi��=����[_��ݺ4f�d1#v�����$=D$�Ho��=�)Z7�����<�Sͼ嚴�_��6�2t�m��^�����9���i�*��E]+��p�{7��D��59�K�?�����P���m.>�/�+^�w#����߿03ؐcF-�h{]�-1v�� &���nvm�����1��xȧx[Xd]����%o��kԸ�R�~ST�P���6"�gt�Y��{��
�1�ޭ�|w��`�as�Hy�A�]ޢ��cC��X{1�V��\.P�/a#4�ĥI��Gc�P�t�)���'�$�6d]��N�q�~�Q�ک�!��8nA�ވ��9w�讞�[�i5��\�Q���E��� ֗�*�䶭��<-3s>T3j���|/�]��}%�OuI�9�NVsȤ���5�L^=چ�Lz�W8�e�������	�`���!6�w#�S����i�p�S�&-9A@%��C���!?W�������o&�2��F�[}�h�WLA 2�1���1;_z��7�R ����Y[���Q�6��^�W�0�^�.���W'e�%��J�<��2���G��c1�;b$7-MoBm��re���� ��T���.N��-y���g��od���B��ɦ���l�f�'���0��Z�:�i��s]���˂�������^4�1�B��������'ڰK�ժ�У�Z#��O�J�����۶�p���J��4�I�#�U���Jr��M�_���x�K6VŻ�l������ !���C��/Yy;Cʩ����[���ևUؚް����u�e�d��_a����A���û�`�8>��l�x�E���e6��Ks!�e��k��~��Nz��H�v���-�ܱj�a��v��j{�&��|Dk;E�g��~��#X�ݐ��.M��4�reܷ����W�'a���ڰ�鍀�]sͼu^88���:�:�m�oO�ј�ͳM��Iv7�z8ą.�v�1j�#��C I�i�ִ��6�l�w��B1�x=Ų/3Y���6U���w�8�/׬�|L�{6�8�Yx��PH�3׳gc�gO��{�`t����b�g|j-�I�ۻ���{P�@J���L �w�y�b��.�g���@eEÛp�~AH����;r�Q?���qמ�G�N?�g?}Ԇߔ�L��]^��V��>�z17�{e��	J,��9f���.���p0S�QV���&��q�[r�4j��^jY�^��Zݛ�e.�N��t�H�Z��	P+�s�kF��N�b"PA'S�RΝ}�4vI�+��������e�d��8}`˩ũ��i���&�sϯЃ-{� ^#B��T�S.��Ψ��B�2�hz{�r��V�{�%�"���5צv�7%ۄ�Inj�2�S:r�	�FE%QN/q�&2�Ѿ��.f�6*T0���}�BB�i�:AĈrO��ۃN�L4�R���LV�v�j���`}����k��"�;���.͔����B1���S �y�%��k�����V5��c�TUwFf��UOK��$���Z^����;�<;�A��Q>���^S�x��P�\��G�7�МD�aG!s�p�r�ͥ%�v���'�vh������M�ڝܦ��{�7
a�v�Z��^m�{�(Y���,�%���̦�z*�d:83F}��˜�;ޘ<v�ྭ
��)��֑#������"�x8�P/ҹ�%�Ts	;bu�o�D]v�b�l��ٮf����X3@����f[C��jR�l'�{&�b�6�)����{R��Z��n,��N�z�"]��<�!�6߯*Y�u��r�üޛ����C���fb�R��7��F���*{F�Jv]�,�n�"�I�������Q��CT�0:�"��`��'[���󇄒�Ӕ��Gh���9���
�dE��޸�w[��Y
k��R�]��;��%�烓���Ő�hN^��{�^D����F�S����k��wK���Jf|tE���-���^g���24E��!�>0ب�Fsf_Z�0�]R�[����q�K�8伡�A!�4�fN��T:&���f|����%�"m��;Si3��n9�պ�UE��n�����E��E\�+��4���M]1p�)���0:��\��s�	� ~�s\�*���ʖ��JBװveB�W�$���oN0���l]j�����L�o��=��K��ѿժ���	&9�C��i��Kfa���%o��!2�hФ�����M�:ws1@v�k�=[�S[;^�G��/��HvO�l�y��	LI�٧��]�&OK\���������S�P��v#g1�_q�=|w�!Ŵx'H>T�!?c8!�c�gp������ۓ��fy9�2�d�g����)Ra^~��	�e��澴����.u��'��*q�: n�󝦃B�sH��}E�G�"���E�{�)�-5�c��Pw����� ��'sn%d����-3k!"۩����]���I�U,U��E����4�N��q.�O�����QMY�/�d�;��Ǒ����7uJ��R��F�K�a�l���%x�4�sgfg�6��Uy�.@U{e#�n�u���:x)��X�nU���!M��_,V�ɠ��fU�,f�0�5�K(����Ԓ��nWw��c����`��A|>?Z�Ϡ���ښ.�Ű-�Nл%Q��Z��R�Gs��=���h�۷�7��x���Ǎ�qF�Rtz:�����j�uQkeb�aD��v4Zݥ��^f�j��sX���tnHWr͵�l�t��@xG�v�M>ɆmǭΛeP��?�|�]��nu��Y�ңѯF#X�{%����;0����辈y��~�F�O�����n�s�N�[֘ܻ%�/�5;׉�&+�C�α�z%�<���$fsm��iڭ��A˅s|�/z�h1�n�0v��$=x� ��Z�ש4yN�o׵0��?���3/��9o��H�ii���"ا�uE����CZ@��L�W�X]9Aw��験�B�^�^Og<^L����}b5���	�FFS���O>�E6jJ����A���ʫ0�1�+��Ѧ�v�:���t�w��Ŵzâ���*��[/>S�wS�n�pk��M{׮�/��xZSI�WN0��ǯ[ռ��|(8"X\� �{����-�!��M��mȻ����i�Y#�,>;�������iK�k����A�UN�k��^��9"�[(��σ��'n'�6�܀�Q3�X���)�fJ�:���S{���Ć����!����/9We`.��ݤX��-ƛ�\���[kn�����l�����H���nt�^s���+�&��������On���t�DԊsf��g2y��]�͊b�d�Ɛ�d.}�N��D�W��)�x�I���j��\:S+�^����&�J�n�"��ks�6�]�Y����1����]���.�L���)9Y�"��Xp��f�v�ه�3IWd�Q�����E��H�=�&�w#�K�QE�mNKϩG+�Q*��������e�;��Ъ�8���
Fi�������`�ZE	�W��1���g~z'�_�YO0pWdB�}���)D��� �C׸�%���I�wh��v�6y��ٓ�ّ:�2���S1�H��@��g+�zRr��M�����݁��T$��(�G�z�x���u-��+[qS\�L^�ѨlsڤR��u������i/���!۵�3Z�]t���*�tV�aS9����=�d�[}��	5ұ�M�,"��sP�c���1�����W�U�k��p[ߝ_�� VR�B��_��<��O���d���ņD�&h�Q2�[��>G��z������>>>>��������[w����{���I�L��J�+4�qVgmg�G�]a�Qfս��+��p���m 3��*� �*8�f� �T�Nu���ap�������궛X�V	�˶9�m��V�CN��c���)�����$�bsڕB1v=����(�]iC#=��Ⱥ��N�Q�C����A�6�t�Jꑽ7�e����9uf9	&qj6�v#(�d]+��q�eV]l�X�6����DH��/;�lV�C�'y7{.����%ti�p�O���)���bWiQ*;��]�z���ۡdh��	�keKm�Ҧ&��i���G��F��]<ˊ�/�;�6P<Ѓ��չ}&ۚ��7�7���|��f�Ubpk�*K�an��؏5��ʼ˩���ѥl���ݯ7��-d��-�����*�g�uL]�M���k���Pl�p9��i��9����n��Ɲ�P�`��Y:��!Vt��sz-�lHM�#fl���t@݄q�wT�v��h�57��׈+#���.���U�v�r�j1h
XZ&dYv�����b����=�J��)�%ۀJl�>#&u�x�۫&J�Z�{��i���ǔ�XB�SQ}IӬ���8���*h����`�ܽ�ѻ�S�����w���qP������FoR[��{rҞ%cY=O�3���gP����#��ï|V�fr��H�,��ҚX�P핕ؚCx`�;%h����V�]XC���У�����8.�,���r����
}�A�\��z�ȍH�2��D��j,�S�w�8��0ͼ�	a�2���uM�yӅJ���+!PS�g�d����,�F�p����MH/���g�^���/s��j�ӭ��/Pv8Ы�P
������6V�"+1��cɳ�¹��ul����b��-��A��E;˕���z�Q ��y�����=��W��M���F��N�ɝ.E�+^f�!=��,�7�;��)��|����U��w1��N��a4�����AI�
��J���1�]�%�VJf��T���-
�z�SM
1mhmS+N�^Ǽ,�Y�8���Ő#�'j{��Q�/3P�ϟ^
�.J٘EN/�W7A��nt}���Ih�ӟCb��W76��̥���t4�<�gt�nm_&��wɽ����#rj[:�z;+8є�q�g{���s�����μ�����U��Ɠ˓�LV���6e��t��5cح#5���C���	Y��t�`T����&F��;:��)����7Rm�''�Q��M���WfEq�C: �Q�Z�񴻐\�꜒��ʀ��|�b��B�B�����-����1�Dn�wcͰ;��w �l�}u�q�@l�7�=�òD+��Y��6�M�ѻҦt�����A6�Ʉ�_�M�r;�Niھ�0��6��7&å��2�`*��񻻬��z+Y��-�An�%��`*'ѽh��z���^��e4��SN�5E�h"J))���lUh"uB�D����@ţl�&
hHh�!F-4N�j�l�P�!Zq�l.��(��t�&�I�؊,I�����))j��i
R�I��t��ryll��IF��KMEA�&��CH�R:]%)�4#M4�Z��Cl������ZM�����4h�
V�h4Pj�t.�4�TE:WBD4�&�\UHEI@m�д�R��P�4�h4��骥4P�iF�e�)M!��6�ZCC�(�M��֒��A�u��KE%�(��b�ֿ�f������|��|�^�-��	2�Æԗ{����-*��0Z,>Kk�8>V��E�`�Z�+L�j�Y]$7�R��*7��ι]������;9kػ���_�՝�/Ⱦ{��T(�[V�~?����}������mD\8m�_�T���v��*.��Ͷ��Q�T5{�ɋE<n{g��:	�#Z�0o�Sr�}��4jVM�����~S݇R���C��C���RFq��l�*�@�t��zw�\e�$�VS�<3;
p� ���[�'|��X &rGu�ȫj�B}c��zN!�;6Όv>5eEÚ��z�ӕ�ҳ�9�̎��u���1�)�.ӽ:Ũd���2�%�:8�
V%RaMAvN1���ݨ��Q1FME6\��g�ʡ����$AoGB�k�0���;p�����	���Jsa%B��a<>\��ݕ}Ǳơ8�{"��o@L�N5C�H�2��.�6�D6�4�8n��E�˪9ʧ'^z�oB�Pc"����n�z�[�	�!#a�O���|���}�15�����Oq��(N�vZ�p�ZSl��c�B�y^=5�N���!��cHA���΂�8I�˯]nk9���^�L��0�aG!s�p�r��PX��u�
��� nC��p��ޏ7�s�����\hK�T���Ko�	���*���E�x�0pï�v�u�Q�(��mq���ʛ�Ȯf�N��>��X�@a�sw�ɀ�1�[<(�\�lR������k��cEdW��T�U��7��� ��8��o�V�?jI�{�[箤<�T{�{�����_�l
VK�럍e6I�d�7��W2���]��wrꈡ���k0����C9��C@���6O�4�eH����4-_�J�[�k���^���9��I��2a�"k�f�f˃��A�5�8G��!��0�R̶�m�u*7D�n��;��M�'sr���uK&��0��̃"]���4Bax���fI��n�P�[vl�����Z�[�`���v���z�3'D[�@�r�5���αxmV�����K;�l�Cҿ�c_q�`��Yy�� ��TB&a���N��@ex�;�&��Ax��,�MS�ƞ9�らp�vN����{k݌ī��P�Az�W!
�k�7^�M~1��0�aY�&@i�k:��u�9�X|.�%>UF5u�T��jR���Z��%G\<A�a0βe}��>O}��0�y�g�[?�p�9�F)�J��[���D��`&\������CSe��<��/�tvP����z�oMl�~@Ŵ��K��&�!!]��E�%�>oV�hƼǖ��˨��VKy���=(��*n�W��p�K�Sz����\}����.�F5��Z���n�.�Ë��Kަ�Ȩ�󿙪՚�e���_i,I%d��ff����>
��#N1�����Llj�Jq�[�}	3���ݔ�M,��d�r�y�_ݳ���f���U&	�BJ�؍�ǯk�<��|����0��j�,W�D�Yȸ��k,���P^'k��	:�^%�u�7E1�$Ɠ
~��u�5��H0͂�)1��F�s{��LT�XW:���>�"Sz��;Ϻ⋦�E�s�2�������-@V�~��?v��ߑ�ԟkA�R(~�C��2i�uL�>�a�F��wGt�x�Z~kJ�)ߚ:-�&f�Zf�\�����h��ͯ�&��>a�6��B5����u~58��Ӓ(�=.�j;�ШM��1��@�v�٪�:3�H�t���zp��#Xt��9��4ݷ�E���U�6ܹ�Wղ�/r�s�'s��ӡ�	=Ӫ~m�Y��E�u΅�4]z�x��D��`�[R�k�i�\�ϛWf��{%Qeb���{���KGl@w@��yP�ʊ!ōl�;�R����7������t�m~݀ͻ��%��Ǥ� �<t=1l�X�c��;h��3}.�xz�GXR���96��cjs\�&����wA!��MCO���7��q��I�j�$�j��i�-'�qⱷ����r�7��f�ʫ�i����6�ͭWq��*�#RHu�c��3���4#�"�X�L����]07T͙rn��M��5i�7U4>V0�1cѺ8(�2��q/�Ύ�z[��8����	�%h�}@�`E�^����^�g�<���5p�E���$���{8P֝�4��X]'v�(u�o�2���ӵOq4l���PЁr����_�g��s���O=xnL�V���\���&0/�ry�k�����
�a�C����F=[���``qm Xt^|"����U��NHyܹ�w.0k���u�}m�|�D�M����ҚO��o�Fc�M<��|w����0D����#a�����(����dC�Hѐg�C��W��d^����:��5p��|j�u����w���M�4H4&r�	�SU�{3��Q��f���OcHBGd�z�DJt�<b%:�.�Lh�I��:�pˣG�L�L�Gg	����!�ly����w�~P͸&82��v
����4���'+=�"�y��@��ͫ==}˘S r3]������G�A��C��jc�l��<�^Ω��rt�}��5$Rx�e�97ܲ�e�jc ��XF�GR3L$����'��r9č��\�ՓMȽ�@�M���n���s�mZ�'��kz	Gs��q�K�NE3��2Ϙ:����<�ob\����=*Y�jzo#��kESbƊ�Q�r�noZ+��ZO[7[t8ҽV�{��$�HNl;���0��wЫ��j��8�4��RD�����pܻni�`�졶7"��ɼ�u>���儻���s�#6Уx����I0��yֻW�V��hH�9P���;P��;j_L��+�Mc]��I�xRήOX�}USN���1ݚ)�3�X'c�U�3u9��U�"��6�B��>��n��Bը�ë��Yk���U�i�a�;B�J������긠φo6�^����C�&��LS�P����hux��?M0�H�ņ�&/��֬�xܥ>�WQ{z���#ѭ�}:��ЇL�2;�~�eHL��Pm�E;t(����l�6ȧ�qA<���������Î����L�D�ǐq�ۚDL$����mNw����C޴�(-�=l�^��iZ��!�aض5'�E;�����2�[xC�["�6�6�Òh��T�w���6�,�!��!�P�o�FCH��e]����{�<VT<�duU	�N�dN��xC�0���(#�v*ڽ�	>����z��ʒ��r�n*aȹ��Ԡ�cL�|�����7�vC��ɱ\O�<k���&������]�`���=hХ`J��,���&�f�M���V�/P��΀�ޏ2�t=0���Л[�!2.\�彾oA��`��3]�� �4��DU������Nݬ��{/�ONg/i�F���4$��յoٻ{�U�A�MI;��J�
��&t8�WG���ކ��A�	baL$���e��q��]�X���&�M�ᇕ��r�A\��S�P��L s�]�;��Xyd��m;��W��A�{;������ȶoM�Ӎ�m@�AāC)=�*��0gR�U�S�#fd�j��}*�W�@L���]"ds�_;5��́���:��/[wxJ���
͋����B��i�)=�d]ct^z��yG����6�\��������Hꨣu���t�IEИ�ca�"Wa�©d�yj���^҂Ƽ��0����܇�E�Q����x�We����x���/0~i���K�QI̓Y@���)$��(�k58���1Tm��j:�m̙nU�^uL��[��?5��	�vLe�dRAD�qD��{ �%�X�n�U�!��J������lN�sۺ�:�f�69�@}O;0̲����T�|��QNƣ���]S
i׳`N��r�nc�,����d�f~ƈL <F[��*Y�}����e�[,�6����Ge3j�s
�Iv&�>�2��'D[�@�r�.�����o`Ie*2"^Rٯ��A{`�f��wS0�^E�w����z� ��L����=*:}�������ٸ׏�����ØZwK1�[��]>,Z��X�R%��R���L<��xF\�ܐkR����em������]p��Κ��^Slm�u0��h&�`�N�z�tc૮��s��DyM�BVe�)�N�����Id-Ӷ�lb֛=Y�{eM���B�����|�T^=���4�A!��	r�9�[�:g�,�67���n3#r��f ^Y�h�a��qqw4^�T	��-mCR��κ�����[�7.��~��ú����!s T:��L�8��\�È�i�%cj����ll;=iS^��{ڝ|{݋�W����
&~~�N��au��f����	�R�l_;��7�v�R�;ݸ�n�o�2Iy|8��$�^��W�n���Q馁�I�k�:�]�t��Ku�nWn9��2�N�����l�:�?WH��^���y�'jgR.5�C��}���:,oy�_P��3�ב���<o��g׹��3�7]�6EDp�k�[�I����H�; nt�� 6��;�괉iC�T�õ;S\�7�N��I�sl0���~��Xپ��jڠJ1��*-�gm>�m���'0���s���k�o^ϐކ���j�G�띫w�������ׅ�9�Yj &;���ۋ�lbJ"��~��c�t�$Xi��b�͡/�oJ��o�C7�&�����
�����V2��j�`M�1�ƅ= ��g��z�@"1g��z>�KX�_[S���Y�*��s��r�a�U/#{�fz��W�j=�3�S�ȼ����9�Gq���z�+�'̞%Y-kpT�9]�w}χ��Lt��#�6���4s?`�nlL�F�.�M�c�pb?�jm5�5�����ׄ���Qh�}>���0l=;�hɽ����1+��͍�J�F�gk�l3~�8	����?G�o
g��<���yC��=�[�w���R>�ͻ�v��臝�%^���=���H�����d��^��^QG��?�1u�׫�~������V��-yyH�e�s	�k\֜ǀNh�4�]l@͵"�l��7a{��V����.�tl1���7ѐ�!�
����t�v�̸�� �tհ��疍u�Յ�i��j�\T7uM��	��*�2����f|v�u[����r�]3&9��vqf�=�:$��+sq�v�k��w^���4
*���2�/]OA��Z����
�خ�un�)ҩ���n~�y����|he�I��54Y��r-��jȚbЧ���o��^4/���v���S��ǹQ(�n������W#s����st�U0j�R���:�����|�ґ�f�n�ݥ�V+?�ys���5.��Or�����e6����)+�n\lokUWT&Ş�8��OG�=d��6�.<�-���;?[_��Se��8��r��{���o�ɖ��|��+��[��<�oO�et������)"�+��ޒi�����H���,��B��u&��i�6*2�f&+��J�67��L�t):��)
�L׍( ��u���z=5],���~�|�<-Wc����8�3Ӟ��H�\["{���mUW��y�.�Nhe[��#�o�`=�bhl���v|q��U�A���G[6�n�;����q۳�_����9�h.Ψ��I_p��d�������i��x##Qݘ�Fhđ|��Fz��w��	��y�)���i���@���E���ƍIjB$i<$D<�9m���Ά�a
 7��~]j<{�6��׍�pb�-A����5x��o��_-�v�T�%�L=����6�������ŝ����6� ��f���=�k(��*EX�I��m�jV�ߴs�.��i��.�_0#5�e&lϣ=��:��L̝9W5��m�m4��M;o6�v��DI��B�����T���Ee-T롡l"��yUF���� ��p&�T��|yԕ���R��.�}
{�pË�e�U�Ɵ��
�_��ǴB��z��2WHn!a(��Hmu����G������EǞhʹA�A"|'Vn�H���N�!]M*����v���<j��r�OfD�p��+m�}��T������ͨ'�Od��D�ml�S���p��q{w�}�����̧s{��)���L�6ڔ������1�Oy���ƍ��ܬ��"������ u���Ux��F�����>�<��)p/�ɽL�˫�3��C
v����*���׎v�v.T-w(S��,��Q�m{��7!��?^�
�գ�ҥ$շ��W����=gǯ�������������_o������ ܫ8.L)aι��!4�֝�Z��܇k�v�m�C�t��;|KD��X��*(V}��7x!h�%�'(��ϯ�F�������K��jI���6;�^J����v�Wh\$j#��l;ܖ���ݢ:*��Zkn�1`�[��+�]����S�b�UjT�V��b݈o����޷)��!v'H?5^��g�}wsk(� 1oYVV�o�A��-�bN�u�����,��U��q�vQ����h**ԢKx��a�э�,[�N<,��b"0W[�Q���x�x������h�oe�A��啚�U�*��(c�ѕ�H�6�>n�T�V�����'�"��W6Nv�1�L��@���n�V&U�sK;�r��M���N^�xɠ�rM��y�wEn0-u+pJ�R�6�<�pX$��RVƮ����V�����-5�-*�^���f�:��8d�4������ SDm#���oJ=��8U�E�7�3��c�n��]=��!�����mk��[�t�����fKG,�����눛�XxJ��|��Λ5��WHP���������4�^����)��&ܙ����G=��rJ:�n<�	��fw��5k�{�8
�e�E,3h1F�PC���'S���l�
ʾ�#�[4"��\,�fy�)ҢT���Dt�=��L�f^m�:НÙ��mh�����<5Ք�`Vɉ;���Ph��r�.�|x0�9tl7%o3�>�ԉ�V�\�Ί	�Y(\�wVۭ��/�H*�v��YAIZ�_s�㴁�醺.(�^��b�x��!f}�j��h���*�J=�����(�̼���'��qW۝2Q;jT&�2�dCdV��0#pK�B�����o_Y�m���]�hQ������v�������շڵ�wh{ΣU��v@�+����m%�5��$�b��/�(�F����/�;YZ�W@�����%sDb��o֩�jkW��Z^�ܒ���3P̊$EX ���F
J��r��m�o�0sy���ɋrp�7Q�M	����|���`�@LigK�P.�Ma����Ƹ,���+����fی_Ws]Ma��J�kx�&�8�/�0�K4���A��J���k�"�5�ȥٻ��YA,j���%�b�Q&�6i�8�J޼Ɯ�Ӛ�TaAZd�ԙVtt�`d�n�RQ�JPZ�h�z�އ�5a�^�K�cv������3qp�1M1%��x.���j<ې8�N��k�w
ٻ�m=��X鶽^5���r^�$ʒ����#�gq�Z�i�L�`��e��`Q�U���O>�!D�_]�@Ýe�{T�MiYY8�ea�A<z�f�#U2U��������)b�AJ��C��G�h���x"��y��$��w�b����ݎ9&�'�I?|�}�=�w�zޯ��o'��h��lM�H�����h(h)HR��b[gk4k�h]:M ��t��c	DBF�!l�4��K�E����K� ihӠ��l굦��iSK�PP�"Z(ҺT�����)M�Q�`M<��(�h���5I�JR4�i4�ъ�ht4U:JM�	�K�WIc4���)]i6�b4%)�&�AM4T8���B�)4-}�C�1-�.�R҆��1e�R�lh��%!ABn��Ur(�W�};�uV���@wySׇ��S?#7���	Y��l|���kn��(�����N�"����Ց��9y2t��kXM���X,�IpD�����?3O~��S��47��1[�v2��� ㉵c���|����<�9C�d�FϻV�����W�*+'=W<1;2���_�7�Wy9��R@�:Y�LH�#�G���2:�$R�ٳY{�z`.�V�8;�t<U*ɼJ��:���<�	/ �ח��YЫ��������I�ڇ��h�X3a��Ul�W_�ra!�h�DO����;�2yo�����"�X�U�����*��rh<ˉ�1S�H��u�O"�Bڍ�K�긚�58��v4�6�}sO�6YЧ�� �'ر,��������s4u�.�qs�56�W�'$ڹ��3V�6��=	b�$�D���3��gr���H�^��	):JwϷr6�*a���@��#!14�/a�N:y�=�,�*�-����oJH���-��<U?WK]:�7���iC^��J��M�%��j�?J��yI�L��2q5Y{V�)s\Y�o3��4+-q�%��[�;�w �]u� lSc�/X�k)��XU-}��;���4UlgWC��%c�y۸(������)�e��9Jo�ۥ�҆�޿��w������Q��!� �Y�)���@�+�����goVo��n��_3����ێ���ɺ
`A��}[��HS@��t�XZf	ae��Rխ%��{��c*{i��º��qǿ:{���2����_�s9��v��d�F^�q�n�2�A��!�A��8��p�;?�&���d�gM��(�'r�)m$MMyWL�O��#��q�]�~덼m��rxu.�\����[��{V߉��&:OX�:Clo6b24�745�Dup��n�,�F�=ٟ�sq6��(�ڒ��8�ʵ���~�+}�����2�vX��ɜٿl�[�tvYy�$I5���$�5��1X����.�<��O쌆rY����yG�n臛���ʋ]�]��$X˭=� J)+�%�YJ}�Nd�{��R4&zy��뤙m���B�޲�كTpb˦�Z��WT�/sWs�v��@Vg#��^&�X��3]�B�u�Ⱌ�S���|���S��%�M���o,J��b߄4��������{�	B��ٷ+E&�]eu�
��g���ث�th�8����"bە��x[ �A�-��sv�n���iЭ�T�z����D�T��ͥ��e��qa&6�;j���Ȟ�Q���(8uz.2}�B�PSJ:I�Tf\K���J�躻����Fȅu�"F��u�jP&QH��̝������q�[Tn5E������j�T�	S��#�t�t�x&�*��T���e��5}��o6�g�{/��6��u8��ä!�(M�oy�wJI���fr�.�oE^�y�yw�Fc�`A�"����; �w
�3#׏Օq�\��=t�wR�T�[-���=��w7Ct�F��	+t��b��o��u�nQ���3=gb}\��	w.���VA߫4���/�~Z��\�VA����^h�L��Rt9Uܔ�^�4�ƨd����s�M�v�T�ɮ����P�#��p��`�����=�@��������q��~��Y{H�)`[9S�li����N,7�D�@�D^�y��w�7;�SQ�q��ؠ]����A�Ĉ�������j��n9n�Xj	�v�ƖI��&˘f��%XJn4qq�|D���3�]�Ù������7Sr����CV��T����^����!oa��/�)n�w�ޘ���}�:�:�nFI݃"y��H����G3�A�u\��%~�L�i�Kel�ئ׵���χb�P�'��K����1�΂��|�U�E�0��xw'.tFW�WZIP/,���xO�"�h嶹��h�\@sԁY�Mʚ�Ry��M�F"jVeō`�u��Z%.YJu[���hQipw�Ѫ��ў�:5��|�P�f�˪r.t���A�EJ�����r��d4�\�ٜ�W5�f�>���ƃqb;��jѬ���B�%��#��x��>.kA�&o��0��UP=y#��&����u��`��dWv�:3l.�0�e�N�򉤞	)&;�_-HܷR;2E�H\����>�4��j�]q�5��j�ٚ�ώ������D����Ndf:e��xH|�I�f���u�C=�����$^u�����d��p�v��if�"8��$�b��V/
�۔r���H��8��|d�����]ڂ����*(���E����j��1��xn^+�ʥƟ��4�1�eG����1&&ƍacgu:�\��Sl�k�����پ�W��\�Zeq�ڔ������b�Ȟȗ�}��{����@�s��T��zD.�u���*�.��H�]�w�`��<�-ac���\�3�?x)Z�{`�B��'λz��ޔ��>9�U��ʭw(��eN̛mnv�鞞�0�j^��,{-������@��T;M )B���
��"�3wr鉛�����"H�&���hl����Ái�`8݁p��\�-ͳ��v���6�z��n�^)�I�2�FOtl��&�p-+�ﴶ�ʽc�����ɵ�?UlØ26��$�~�Ӧ��C9w���U�]�&�m��l��4밌��xw��E������W#BI/�<+|��BPf�0��$��|�Tz:�l>rgG��dE��l��n��Q��{�����|w�p���{��be�}>觍��z�	5������Ċ����:1{1����]<wH���m~���m�Y�E�1��ޱ}�d�mD�e;㴚T��K�2xӷ������h� ��S��&2��Wm�xGb��t���1�ћ�g5gQ|E���謺|2n�U:.����
P�	�e
*�����	��{�bmN޼����o/�&�,�A�R[��{V#�[�v�v��{U{�6Ͷ��4���)A�;W"��Ϫ����Y7�rC���DU�}���v��$+'��XzR BJ�j�YD��{i�m�6�w����C�*[0c��kA���;Ғ��-���p~�_V,9��6<P*p���w�������z��P:�EqhݞJѤ�z��l`{��������V�׻v�x��Og�vv�σ&�aD/pY�#V�tS@6�9�m�aQ���7��Quișԛ�#=���p�7��+b��sn���S�+\�=�KƬ$�/����H4�q�!� 0އy*����ݫƭխ�ƻ:���H��rY�H��
�s�d^R}���5����\u��z�v�8�R�ܐ7:�x���>��;@�����{����<݉k���0�Ţ�4I�>c����\nwv>�e8��ia�d�y�&<w[JHp8�n�C;/�\���t��]�B�`���U4(q���U����j>��4�u��R$^��D�ƭv�jΙ�יִ����(ƍ-�\j�U���J�p������|@�E˷��5�chw��F�<�f uj@�$n���_��NRc�� g��������3���2�Ch3��*0"ά�ËK�6���^}�H�*�����fQ�%�f�Gu�#;;)�FC8^�z��J�o(�m3PR/���Qu�����yl�����E�eg�)�CX/�'T�l���º��mg�s�ܦ�*/�CG]�D��H�O�mO��:��q@�E�i�"��,�����dS�Ѯ@|Rސ#-��r8��R�'ii�ɹ�&�ܛ�NGm>
��oPx`z�꟰!���R.ϛP(�G�FUFs��l�� ό����7�..b�+}�*�"lB*F�p�غF�G��h�����.����|1j-��^���ipE`t�?)�g�7�x���'/�3;�ه��gn$�׿Q�M.��e�[ւ��X�4�o�ΩF���'�7�7��\��㹍&(mD��Ы�O��`"�?���wo��n�)G�6�5�V�YP���[گ��9���q8�󙩡�1qr�<�:�v,Ma�y
�1���u,\� ������'��6��[VM���v�F�=��m�����p�,����/=���l�@�<T�u5Ovp��z!�F�_)�u��R1^K�v>`�-�W^�.�SFy�î.wFeh���d���t�%��{�)W�d�35?��nT�r�'��>�����4�B0�##��w*0S��j�$��=o��^�R�N\ܙ�o^��-�����a~x���Q�w݋d�<�3�B*�eU�m�Ck�K�}�&ef����6�Hcc��G3�	��u\�H����2V[�ÅWd��j���BЭ&�{��}��|��{��%��=Lq�|���|�cf4]�:6���_+�� j�ҙ���]��7�G=ltc�obߧ�W
1[�3c��;_��D(w�^���̸�H� �hPW� ���-�9c��1�?GI��o�#*���'fgz���� Ȣ�?����,0��Ne�dT�9K���	��)_�N5���T���IH��;�n���R�}��֢��ط%:ڶ]eo�����ކ)�wkY��t��Լ�+��dV+����Qc;����.��[�����Qc�t5]ζ�2����}̮}W�(�j$�1uOc؛<A���Z�Ӵ��+0gj٭������Ot��Y�#���<��^t��� z�s�		#����4��vB���94k,ӓ��;9̸�e��$�e,ܷSـH��I#cBh��LŜ'�v�(�#u�G�_@���rI_���D�l�S��a�8n�{1wN�+z���f�`�5����`m�T/�u�Y�WmJ|��d�fʆ�ے�*e��"�M���,��-2�.����X�	I��=$���+g6�W}a߰�ْwk.�̓�|�<T���EP3{';*�r� �␉�m�홻�/9�pz�O���t�|��f�a�����[�s��(+#7�t�I`S�_{��7��{�];Cdu7F��sf�bظ��Udkbr�x�h����8�ԉ	�p��wF�i�F�!�����=�v+Hѽ����#�jNޕ��N
�uP��rѱ�ؾ&��;_���YZ�b�+�kA�F���X(��{��M�Ȩ�Z���
p*f��+�f�[����H���5ܲQB�6��Wk��vS)��Z��'jt�t�:��7���G�1ٍ�Fۍ��狮�l�3�3mq&8w��� �=�����ɮn߈B�knU���;סym�����c�t�x��y$���e*ۿd�3�+��kt��gf�ψط�M�_|E�������Ľ�Fwޚ�,���Y��%q�v������/�a��t���S1ӗ���;[3�wk�7�/[َ��*X�[^R����d*h#�8u���Jb��вw{f���]�;~�IU�*���z��H��2*��6�c:ۂ�}M1�9T�<�z�����d=�R�_�H����c��"�'��;_��߉߾��8Z�;����u���[{o���$Y���xז����6�mT<;C�Ǌ�W�j_s�9���X�)nOl���n�%~�+g���P��fL!���Ne�֓U>��ͼ�!���)�8�dƭ�}�����}>�O���^���������}��7�����������u4�h����)��)�C��U���S������>σ�ɲ�K̉0��<5Zm�����0͢������l�݅�'���2�(ڹ�hc��k�r8�-�������I*�̌�efwۯ����=j�.=T+�[Y��Z�͛@��e�Jek�ר��ub_k7�;%�,���o+<�j;B�x�"%�6)�S��v��2��Id��-q�Q-��sn���z5�6�lƷ�K�s%E��ٔ��b.�J�za�n�#K��J��m�}$�8�-ո������m���G�R�<����	�	�8��:�l�i�x��z��!��x���Ǯ��O(&�du��p�ۮ�����y�x:��eI۳��B��(m���T�ݼ�[ц�1$��U�����g��x��IX{U)D]���P�S�S��4�N2NQ�V�y9��]����+r��u<:�`&Xd0�1��gט�yy�!kx��G�N�&L@h*k���Z�f�	&0t�t��݀V�|�`�����'
����Ν�n\P��F-ح�0�v��)�Bخ����w(Nj�psu,=٢�,�*�5W]Eoc���p���^���ACҷ���P���M��F�"H�x]e���I�ѵ��a�lqu���mZthƐ��]�};����8�vWsh�*Vs6��t��:��«i�F��N[�rXFs��>�f����
�h )����G[�ee+U�Tw4�Þ�#��9��"_d���u�m#�|�^O���m;O��s����s3����k��jK!��m�)�̚Y�^���a�)���	YAs5�~�2�>�NY�|��J�_aٹl�����J�ŴK���ρ� ��e4\\s��D��[9ʻ�g$~��lis�9��{n��/�R"%W��s.*U�VW,����9�oy�e<�,��|K�=��V!stf
�[TP�-=��ܖ������@6��R��ޑjΧ�L�!�M8dq?N[�`=�,�bOsMv&'}qPȣ<�
��Q�7`�j'�6T�R����P�� �N����V%��`O�@F�P�$\�W��\�b��\e�$9v%bP����{����vo0���Wd��kf [�{ǣ�`T��wV0Y����x#t��,�.þ��Q
�Rt{�v�bt��qѰB� ��˲S���j<�����R�L�D�'3nJ
ڠ�<��q�s���$���c���r�B�^X� ���*�vm3ّ�������V�7Ƈj�/��/�l,���
�I����ύv��t�z:[+�����X��lBb�̫=�r5��+
�0Z�f$�C��BS�z�Ŷ���8ӹQs��ek�>�i�8�u�|K�}Vv��D����i>}��J��h�����
��BT?	C�=W�nz/{���\���

R���B:qCl�	BiM:]&��M!Z�� ��].�.���(���)4.�t%-R$B��4��h)!T���KH�֒�&���T%6�DV�CAN�	�""��(Ӥ(V�ѧH�"��LIN��4��))ii()"o�Z�w'���!R�������д�4�j�1�h�N�44l`4h�m����jآ�@�AJiV)/�<<���wׯ9��}����fӋ�%K���*�&<v����
�xZ�����Y���68ɇLik��0��+z�����;WXuR�A$��n��6sU�y��c��߽��\�f=����C��w)��<��ˊ=]u�H���X���Q���wd] �Ɵ!������S�Oc���OQg�L�En���rr�w%��54?�d\�&v;���F�ܚ��tE��0���d��S�37:V�al����N��ǟ�b���� �=oO>�K�2�z���t�h&��7oZ�%�{�\�R�I\�Ct�vmGd�6ř����w@�L<+5��V���^z��<V_��/tv�t΃�0�{����c�	B !|ܒΛ�Qs0��"�ٽ�Ñ�l�9܍���"�{J}��
=��c�	�e��^�L<J՗�u�4vG���L�����8���d�J�8ӛjn�F�Bf�h���%�6��y΅K�n��W�/�E�.!^��1�W�>'�R����{�ϫ��V�M��v:P�Q��!��
i 2��s��;6�"��.K���j�N�����W�U�u<&i��k7S����{�G%e�����N�u��)��B�1uo�����[[�wZ#���p^�S��8탴���	>��+��5;��܍X>��!]�p����+��D�<��1Ӛ͌�Z^��gl���ʪ:��՟<H��UB*w�{�t�k�g,��py���U��~���:�*���t�K�)�}�H�nCtwBPv*��m}���N��'��q:����f<�A�����t�T���{�L�9�Azގ�����I2����r
�n�ж!�	������������R���C���3"�#���]�A����
�.ۦ��˜ިz��씌�7��:�t�4`�w$�3��USO�7��K[6�pM��������d�!��pVO�{$nT`����7C</u���|�����(��Pv�N�m��{|�C�#Cd-�;k1�݇UF�V�M��"����*�dx��=A��Pְ�:��g�m;(d+D�?8���Gt��X�ur��3�໯�M��⃎��Kn�AaQa�bѽ0^�1H�]-����޻J`HY��WY�B���(�ę�Z��rƑ#���S6愯�CG-�;Rӗ�M7�z����X�Q�7�>���\᳍O{����W PP�3��øi��A�F}��� c8���oL�ךC�GC<���Y63U��xIDF�h��=9�Iyf���3b�5]Dw3X�^�J�5u�X�GU� �]�U9T^�Q�ݣ�U�����5@�z�꙲P���Ievq��������27�����W�{OTTK�Yub;�h�J��˻Fm\�m���E���=|g��Κx�g@��.D$f/��Ίq�X��7��u:�dk��.�$�g��u^�.[��#�hY㰹x�ݶ�l�����H7I�Q1���R娮h��&�K���·�+�Q{�#��ڕB��{�J��mIo>_���J�U[K>t��Ά��{T`�K�7��� ˮ�u��J�.��G� >Vȋ�s~33��^��tU1��Ԯ��]�ÇsM(�h�]�`�����,��0��V�ę�r�S����(sЃQ����9��gf��M�7 �,��.nj JD�,eY`��v��Y홓%+v�;l1hE+z���ƹ�[��l���"�W_���O�������`r�ޭ�(
3fNvU���g���؊��龹9�&!n�g1�,2��A��`WNOj�����U�숮"��ȁ|���`��;ǺQ�v�ͳ���h�C��$�~7����?Xq�T�T�/iYF�u#A?NQ��v�/��!���υ�)��Et�6!�#T<]��K�p[0d�Ę#@$%��=�/��NX4��\�-`^uxMAz߯����9c�K�������#~���7{��r$�;'�
��qʌs�*1���X@�k�0�{W>٩��N�����Ţ��8�~��(����{�^�Ίx��=�$�plL�[ahJTӵ�i�ب:y-��4�L$�9��嫉s{,�S�F�(�"&��1����ۣ��/q����������Uh�Pk<v�EM9�V���
x[$���SКmg���˨i���7�.D���e�-���괘������K�(2�y�S��ɶ���p�ˌcEi������r��Z���t|�Z����zo�y��+vո8)�����*Ҿ�+2�.JI� ���s��cι��t�E&�k�"� ]���L���m��y��)�*n_H��2�w2� �������a����ro'x�h>�g��J�T�" ��	. �%^[<��|mmU�g������5'��r����;����5�
Gc(e������f<h/���x?i�d�������qzŖ�l��Hd�� ���,}[��$�.6���&�Y�z�g]dl?��d�q���&F�$܌X�m�WC�و���[:�j3/#s���ܢ:mV�x�biay't���>�8C_ݕ6j���n��/��ѩ �)HɝU�*C�Y�ܖ�L�yS��>�O��Z�����YU����.$Q�����Υ^0�y��w)��/\�t\4@b�'z�����ɸ&���3쐳p����~���'����ؚY]��&�d��R;E��}vr;�0;�c�4����\v�Y�פ��`w_�|1j���sCЄ%��c.�&&���ቴ��)ӭo���5e񮬬i�훱���Ɵ,��N7�W1Em������}�r��sc_YO�K��xo9P��&�fp�`�/���Ⱥ�D���\�6;�tV2^>������W�MS��u�X�������T�v
:��c!� �WX��z��/4��9]�N���}�u���q|"�yZȵd��!��GdK��)������uy������Oc��H/u�d�J�8ҵ�cȺe�&��B��2H���z��b��o��P2]_-q�x��P\)GH���Ļ��*bj�3gkq]C�4� P��4!E��jՂ�l��
�2�q�;S{C.pm��Ί����ګ��ճ�.��tVn7��;�GL��3�g;32OcK��7���;���@����Q�u��p!ۂ.�s9���6�7gs+��͂Jn\k���O.�{��x�p��+��Qr�E"zc�v�1b�n��Ѷ��&�+�s���T����$�����ص��{9�A0����.Λ��Q��lW$c��]���w!��@�s�3F�����N�����߻�QǸ��ȏ#�{���F�u+ct�A�#L�8�ޙ�P��mB�	�U��g;M��Qhve^��6�\<���^nSu����"C�	�8���JQ`���W.9��u��)!u�
���s�r9��hi��ʮ����@^7�`;�o���fut;�*�rR�t�i���whܳ�T���hλK�u>k�e��@ѻo@p�����4���"Y���S��\L���r����zUQ��v�͐�{���] :���f��'��9��Y��ݽ͐�$�Lt�v��1�ϡx�F�m��C�lJ9�e\����M�^~N~��SW���2T��������A�X��<���1j�l_�l�Gp��	c��6*ɼ�-ydD����1�@� a֎[k�
� �6�x�/=�����J<�d��]P�e�$v��	R�DfG�K5=�U���`>���+�^�g��P�S�&O���"�ڒ�dLWm@f}���t�_kÆ:G*z�Wc�xr,�+�X���mZ&���m�[�\��Y���8X�3��.4v	�Sǯ:%�i��<��PE׏�­R��ϧ������7tg!=��P��)����{J�7��V�*!��8Ѱ�@�̝yB������+as�&�y��:.g$�)j��ǌL��HnGl��+2���ti�
�P��_S��5�8�Iݴl��T,�c��L]	�}9gm�����}��F�c�I&$� �}��޺�"�N�b�ӫ��6k����܅1�G��!}66�J�t�+��z����P���t��ݤ|N�û�S�S�ь�\��e_�{�J��WmH��Pi��Ȫ���u�*�h��9��P��K�]>��Y��/����~���d�M1Ӯ�w{�OWV}��@;Τ(`�q�<�|�C�o^ԕ�F�;<v��:p$\\l��_=wKƚ��Z��&)V��M0�����a�+��dt\l���T�m�89��b�^Ӵk�0�A�[ǺW���i�73���|�_�������/;���;K�� e��=�g���'(��1�~^5��i����O�)�R���j��Uؽ�\h$O� 䄓���u��y�OO7�6G2e���7�~+�J~џ������ˇ7%e|��$��V,7S�4f'��*'zw<�)�fH0x�,�I�Vz]�J�^X�{w]��eghRM��lb�g[B��.Xؿ�i܊1+�)L_f��Hk+F݇����혟e���Mմ9G�OEc��L��	���ҽN�=P����t�к���\��Do��3�.V���o��1Y�=%;/�W]����btK����t��Ӹ�Z,��"F�M"�Ԏ�x��=�%w%�NDЪi�Uá�ow=1]�,8�B���ơ�jni��W
.�<bz�)�o[f���rE	��d�v���8���4����*^��:�����W_��i���\'m@~�ՄW-�t�\O"䙛U0%c"�ݱ���k�Zb��A���[@V��Tu�|szRE�&��z���]�=Y����s�|{yS�2�Ng\R譡<xu����,L��x��K��C8��NkfwWl�\i%|�gi�� 5;���,�պ=Fs�ú�ݓ�l��m� RW)�y&��ޓ~�Kt���v��a]���A�[Y*�m�V����GDU�6���](�yExqoV�6�A��ƿ?�����W)U�o5�/�Օifm<�C�;���o]D �b�M0Ov�qX;�яX�ܩN�Ln�+�s�]�y�ײ�1�����\���!��lǡ��%�r���X˼\&�K�p��)��v@c�,�ȭ����Z�Q&������IS���;��&vgM�S��]�m���*M����ػ����at�l�?~�������כr�z�l-�χ(w)�,�8ѱt!�^^�����y�T�cSh��v#�̌��p�������1F-���/m�٣rAQ�;]���3병�0³Cg���뎾��ބ�w;նq�E���ΒA ������	�~�j:�]��^�wc�\��k潃��^鼣`v���ǉW^B��f0�U0Dߩm�!�2N���^��[��o!bb�����6�&T���\��!=m�	2���4��P��w;���������]���XW;Z���q������t��Ɯ3��S1g�{���/3s2ni���@�r ��j�n�j1`����x�}�7���'����'n�S���@:���X���}����z}�#����{���w�����|�|ޯW������x��<��O��&��ݜ7��r��ؕ��W�*�+����CS&�f�c�"uP�J6]iʱt6��	�����XI��`,9N�}�Q`����d�^�{0�)��b\���F��������Ԓ�2k��=�uvR��N���U`�H�L��rIw7I/�aἡ��Nc�C,q����fھ=����ƅ_-���d2�w+@�}�1������}>		�+�i�R�tbF����(��s]p˝�r�[`�=�Y�s�~In</�c`�2�1����ȰUKU��
���_=��u�=S����<��@\&*b�|�c�r��)lQ�g�4�ad��5#״���!�P����������(Vr��[�[����F\�ϩ�����4�Tw�My&��HW���cVF�YYY�Hᱧ�۵�d���q�q͋r�Ɗ@fT��	�k��Z�^�q������DN��G��>F� �W�[*���>t��Z����H ����J��Q�LBI�2�����&�F����}�Ѐ��l%K�B�H��:�ʁ��a&��
4gmGpQ�Jh%w��FE�.���Quc6����:��������q�j�"�*V�˄;\ODt�-PwKR
*��3Qx��!�h�[�
\h���ף~y�Lzf�U� �e�
�'/%v�+�n��E��6�WtGp�
�����8#���|�ΗOdk��{A�=ڃ2�ƻ#"�ҥpe�1R#�z���3]N�0 '}`m٩la�:'�����\��C$�w����\����`���d��H�r���W4�����5qP�R*�-e<�C3U�J���2��
3DE֊�	�Fd}�Ґ+ ��CǛ�, |.�fYwC���{�����w:�b���ނgց������2�G�vȳ�"՝�;w���䱎��)�
�0�/�r:P=Д$�!����s�n>Y��\�e���t�\|Z�f��J)Dx�Z�Ɗ}�d:wy��UeE�1�u!ߛ�hG�a���+A#�\�]a�;��r{�!��C�n�P��1�����gmI�05kW��s Ӌ;�T)�yz;a��7�ʲ��)�[Wk��Ʀ�-�(uuH���i2W)�Hi��A�kM��J-�Ev���#�@G�3���tq��:W�P'��.1b��n��n-۔lj�V��� EK�U��ɜ��ݬybi���P��9yi�6��+�?w��pG���)��$]��{y@h
�G�]�(�d���W�����;c;Z�뷲�q�qT���u�,+��+�Jf۵���ZݝLv�r�E6�%Y�SB�b�fep>�*�Vp�Zyi�bte�����Y�s�C���$I�g8k�����M�����F�U�����l����]�;�y��+t�Ff��k�PI�e-}��2m���H[�e"����:б�a�%�!E5���l�j��*Ji��ѪJ4�Eh
�F� �ERRV%5E�Z]4%V�"�X�cH�AAEF�A�Z�()4�!�I�l:iӬZ�m�b��X�
(-a�����j�J�-3UHTc&6-�;mU&؈��lU4l��@Q�]��$ш)�H�
h����j�����)
��E4�@�Mgb�������b��*ִ�b"��hi��(�N
K�HPQ�4��.�`���u�H���[Z)��N(������?]�O���C����y%���L7�L�-�Q9Y؟���j��P�6{�E�:v��H��V�wUN������p�ۮ���ۜ��߁x&���R�������@"���9����<
�k������-zJV�m�'�p�3���t��R��~�5o���i�m�֦�m���4�Xe�9�<;e*Ӹ���gS�\����}ֲ���t�#T�6V�MOP�S=kb�#�tWCC]ah��*4�Nٻ�=���k��C��y�0�s7�:��0r���8ͻ������}z٪$�l�l�P�L�!� ���Fz{/X�`�f/*���T��A�u��؇.����N�m�7;n�����X�c]s-T�Dun
��:_�����^�W����`;fz��aN�����~�U��	��*��on�ե�:͜����4��'E�*`�z$\��4��Fc��/-��h�i�^Y>�<$Di�^�OlE�2!���t���!Q��L�ّЋ1Zˋr來�H��0�:M�R��Ղv��Rc�1�l愩 �x�_\{�oQh�ċDv��W��q�0e0��紭Ȟ��r�PvcX��6�q�g^���RB�Jۤ�膚`�7�����i4tΩ��b�g��D
,���������EVP\��]<��1�r���T���8r��n7��Q����S��A*z��=�����="�R�0��3':e�z]�ُ2Go��h+���z�%���sA߆H�9�$s�]ٽҒ�2܂�%��FyTy=4�MH����N�p�ͦ�]�,�*��DZtjH��h4�xSg-N��j��N���ؚ�lC���I�a�fz�m��@ͅ!nI!�w��3]�»��U�5���*_Ku>X�B������4�م��J�i���f��5��{ZR�;����_�d���0�z�|�J~{����
�G�*�6a�Ȉ̝�8�I�u<�K����0�t0[M�wߢ����L?.|���;T3ԧI���>�<��r�U� ��0��̀�o������-��In\E\se�:��A�R�����^�tg2��!�+�X0�e��я�4h`��S{1V��U%1�x"�<�}̰w*�ӕ��8Jb��Yc ç��;f�$1��G��بl��8^����6N��*���-Skmm5�=E���vx#0��"��Ҡ,=�8��^U�ПmXc��W7�5\S����L��'`\r_r�����Q���>�ц�-���Z��[ʍ-��>|�0r������`�mq'}$p2X�rwv�dVm�
���S�³O�����3��5�F��k���*er�g�~Ʃ�¹�X������ùhH�x�ݜ� ,�%�5=�ېdqs�$1/sp�����k��q�4�m�����=�A(؜�
�
?��z���C�����ֽ�;�z�PS�J��.���R.i���j�1o�.����k��If@�P=$m�W����ܒ�hʠ�܀v���5n�<l��]�-�}��&����_-�3 ���IH=�nz�`j͊�]�*�v�32��Ǧ��+�Dd԰J{���;Ғ�?�vF�Bk����eC3���ch��%ʷ��YBmr)��{M��(�h4��
����ڞ)R.����%/oR�A]>ه�r��kX�K����z����&'���Ыm�<��^ڥ\����_�3n�x���s(	�E�<s���K�#V�:�� �8�o\��V�c�L�/������m_�]Т* tV���`�l}�r+s"E�Esp�텑��i�*�	�"��P7{+k���\���"_�4����ʲ�����&�e4[�urD�O�<��0��]��y��V;������=)/
tx�6mwj��Q����wM��L�/�#Z�unAꜜ�/lt]{8;ӳ:�æSwQ�K�&����cD��.c����l�7Vq͗FR|���·q���j������/�]vOe�����-�+u�=c�6��g9���3�H�-����zJ����{����]O!םѳ�/�CW�XCǐ�����Y���5�;o}� h��\��r��n�A �s�
��O���-F퐜����h�;�t]��y��^:��tC��<U�>�Ee-yrz5n3�ʍQ�Ol"fVu��82'GZ�,��+;���hN}%�F��S�rގ쑬���܎"�JgW_��㘆p�H�<xR�O�V��������6��)\�>ܫ��T���B�D���@�WB��Q��Vn���vW��ǭ����|l��=g���;���,Uq�����$6��7�J�K[�f9�[�]ٰ�;��0�v���/@@W�T������q+��Љ`�Ѭcxx�c]3\�{����ݙ7-�c"��< �,G\�<5j�p��!�{'t
�'n6����BAd��e:����j�SV�
b&ǡ9�`���ʖ�i���{�dk�c��N��\QR�=�u>������X�fMx�Ww@�����^�ˈ���.&Ώ6cّ\�Ōt����f��]�,$�7��l{njl�%Mir�lyg>4�������&����t�����h[��t�����Sֶ6�#X
71ʳm;ֶ��7;g��v2���f�`z<��fuWI�^0r�J�oj2v�Vo\�g�9 �ѥ5C'i���F�����y`m��&�O:�l5<`����@��}x;?f�fW�u��
�t���|����KR��;��o���@j�f�b[���'-t/S��S(�']@���|0�D���pE��e�V0#@`+A���Y4� �[�[{��A�,��W�V�c�M�է��6��f�!p~T��{��Ӎ�{��Ϯ�n�}�n�NK�j�\SY3A�����^23�v-�G�l-$�v��ǝ�
�q�z�uD7WX��uBı���\�U��tY�>=;���^�6��]�Dp#�}��g��s�42����:�h�i��#�� ���`�k0�ޡ�� ��c�1�}�7��}��<�7�F"W��۹���՚N#�����s���#��X$���ޮX�A�q�8���O)����o;̹⧝��N�B���Z��JUx��=7Q.dag���`r��;]��p����i�=F��܀}�z��'�� 7��(��FyUx���O4�39��/oWe>u����E푶�Z4�Ɍ#C�.I��������b"j�jw�gx�0)o!nB�m���t��䒰�&���'�:����N�ʍGԫ��34U��X�e�s{�Ч}�)�kޝ���������̿�QŞ�u�X�A���q%Ω�Ԭ}�+Q���N}KV���9u��} �In�ٕ���@�tReǔ�s�ZU��$9��e���s�#P�*
����3o��z�CCx�5*�����0g`W9�fUz�h�뒴�v�V�a��!�=D����8��Cv�Yo�s��1ϣ:�&k:�r��=��K��ԡKҤh���P���g�7_�P���O�D��;���w����}�N�<�b�)�{�o������i����d�f�C��i.LܭU�i'W����=ԭW@hl���&�t�S���ڞ��c��	�H����|����ڑ)�r�Fw9�v��R��.�{a��1ң��� ���ְf02� %��6��2GNSL�[wWԩL�����wb=�+gU�׺��>�,�-���T�������J�:=�P)Lu��#J"I/ ��͈�B�����^�;9��Ep�}���X��D>�ʈ�ɷ׶�â�6�� o�sa��ΩA�n���iA�����U�t���wWF�J4
�	f��em�d☸��;́ؼ�[2�iv��u��JuչB�>�������O���X��n��ub�.i�2��i�pO*ѵX&T��rM\�X9���#�BN\�[̘�[���R"����M����ʓBf:r�Җ�:��V��e˿mWi��ܿ��6?Kة$�$6tc��a|��iŽ��B��IW�U�ߦ���L9]p�����:���j��YȶDb��] �p�H=��Ë=�XD�dѮ��� S;�/�����,�u2��x���BQ��@��/WG�b�EBji ��oK{�f�==��ІK]:�5���D"��<��s��386�YosQ���N�*ѤU��*|������aN��Եk�=���[���[��x����[e4kb{�갑2'�Fcݭ��LU�/5�Vf����0��ǲ!*پ��[T	F&��v5��e�nNN�ڣ�:��`{��0*-��`��!ɵ@�Z�31=On�uBk:�WV�vr�T�'[��{�q�H#���/^X�>��h�i��l������ �+�	tQ�[4؛�>��#��ofO�u_�esy^�Pi�HW���F:i��{�-�)����.�Y�����f��#$�8�ü�2f��Ww	W�8<���������
��双M��s���ś�E�w�4��v�o���?����6�5h�!vgvB�<2f&Ng��������w�����ݒ��1�F*������k���C귫A���οUl^n`ͺN��H�K��謝�~��u׏L��U/
��lv��V'��5�o#7�{w�tC��%Q܋@����1UWݯc��!�w#��͸����a�BHؙ��ǬԐ�@�&���S�L6���#6J/�+2םngeS��z]����00̪�*�����Bɮږ��,�{G��^�1�8�v�1����9�ASB:���Ww{Kf��^u��Ә�8X�*��⑵FUB��z��U���G�@��ɉ�c���_��҅���7`�)�k�I�UqEKl��Zx��*��aA�����\�w���rY-��;��:�ܸ�m�O.=|��o��l3�O��k�h���q�7�Zן��]��%�}Y�C�Ҕ�3o�Ayش8�L4Ȼ�J�'{I��eֹ���?z�~)����V�����m��&Sޗ�p�)�G*A��2P��غ�1T�_JƯ��QN(��y�K_WU��.�_o<��}7���[>R��GWlE�&�⧁4�Xw[Ou�5�S�וUvgN�kר��
R;�rB�#z�϶zz���ka��n�����/��kX4`�'�rv<ia n6G���tc��ꮓFW^l@Ƶ.�FI����x>'��{�hҁ��m�7�0f��n
$���a��3�9`C�R�0��~�G��d�O gc��N�m��a��؁=0P��:"0�͑{�;K��]#�{��z��/�Z��]8���09��S'{�èEٺWw�^�ۇj���(�~�f�l�цw�=���DQ���K<wi���}�����
0_X��S�V��4���"Gq��h��|�I��al<��v��o#d��>�Ǝ[{�~�A���<�}�O77�^���l�&��y�ƻ��p��<k�E>��5�7>�^�����-w�&'�����攑� U��TE�=�q?퐠T��PAA�p�c��>�oH�d%�f &�`Y�	�fE�FB�V`Y�fU�VdY�fQ�B�`Y�fQ�V`Y�fE�BE�F``Y�f�e�f��f�dY�f�FaY�f��dY�f�eY�fA�V`Y	aY�f�FdY�	�fQ� ��fQ�dY�f�V`Y�f��F`eY�fE�Ve�fE�F`Y�	�f�Ve�l+�`Y�w���P��((̫2,��̫2,�3"�3*̨��P0Ȩʪ�aC*�G"�*� !���@�@�D@�E � � � �VJ������ ʪ�  C
�(��0 0 2��ʪå� ª� C
�  ��2��ʪ�*��<����( C*�*�0�0 ȋ2�ȳà��̋2�ʳ(̋2,�3�'��*�0,��"̫0,��*ç̋0,ʳ̋0,�3*̀������{��� �$ʪ% � 5��7_�t�~���o��?jS�#���-#��
�IH?Iw�o��ғ6פ�b �I�����TU{0HP@|<���q��@�ܜ�~)��Hy�@]��X�#�ż�Bˠ+�J�S���L	k�����2d �"Ċ*���(Ѐ�*@�B�
L"��� �B� 2*�$��# B*��B���  B�Ȑ � *�ʪ� B(	�B" �$r"w��w��"(�@�� �
��C�?���[��@tu��r+�PVA�A��'�6�D��'��`}��C�ʔ7���
�&��i�,'�-
��" �j69��I�������5�0 �*�N~T�xMh75�$hK$��JC��@�� �bdu�&Hx�<�@[&F���^g�ٿpvfj���;���n��� PV��<�(�
�@�f��@�M|�F`D��� �g�3���	]�Q h��DZ�$�;`o�����z�h
�+�̀�b�򊊠���A�m�~�$4O��d�Md���x�f�A@��̟\�7�b���U��F��JV�aD�2I
��KiBMd��((��TU!��V�CZJ��ka��(EIUU%Y��RU�=�Eƚ1(ٚ���i�2��[X���Y5���m�fS*�[m����R�aCl�m*Z��;��-V�c1�T�U����
v�j������Z�j4�$4���mQ���F�5��J̴�E&�+k��
Ճm������h�d�ٴ��-���)i-���a�m����'l�5f�Z�  r��4WJ���m4Z�m).��v:��V�NuZ5���Վ�:�Ym�kr�eeSWNVwYU������.���4�K�1vݛ��Vwm��D֋[X٪F*U�<   c�bF��d�
Ɔ���^���$h�1J�E�&��ڶ҅$m���}>=��}�ٛ3�p�źk�V�*����z^��ݴ�ss�3[[gl�mJҔi�S�J���ָ(u�i�V\�QKf4PҘ�L��cVO�  �ީv��Ӥ�gv�Т�nG)�ʎݵ��ƃMu��7v��)m����n}p�jz���Ǯ�҇u��Y��fح
�we�:��wV[lWpV��T�����J���3[V�c2   ��m-Q�5��;��V�E�N��vj�����z���ۨk۵�'-k����m�m]�n��;�(45[�Jѥ�lꪥ4չ���t뻭#YƪY��cC-�π  �޵@����k�V��f��x�X���tUJ�n�e��64�F�v�e�vq[�ttf��k��MWZ��Ҵɳ,m��e6�[h�CmW�  <����[�����nm��Y�ݫn���5`eUT�l���sGV�Q���*ݶ��ӧ]u��V�ӣ��ieU-����d6b��  6<V�q���\s�R���UKn' ;Z��5ەֺ:�;wP4�����.�:�g�EAJ��S��$)J/{��袕"�Sش�Z��hFf6�\�X�  8�ԁ*���מ������ǞT�S���B��P����D% t�%T�eWz���P�Ts���
���z��`�QJ�Sr)J��7��Tٴ[4�j��m��-�   ۽��U))M�W�U
�T����W{�wy��E^����g�P

w{g�
PP��=%@�V뫏L�I]��.�AB�1ǛMj#+mH�l�cmG�  ���%>���AJ=��xzR��{x�
U���*��T��%T��秽ф*H��󞔥N�K���U�w���z�ҥA_"y�%J6�  E? �)IQ��i����%*SF�4h�!��)F  &��T& C@��)fUR  �G�G� O��������Y�����/w�]"��,p��v;�~L�Yf�^�5?�W�}�W������߿����m�km�Z��kk���j�����j�����խ�Z��kk�_��T�y?��D�E{�@m�[5�KY)aB�
�,R���MY�b# 5���p-2�gێ�5Z��-=��1u���X�ebw��k4�pF��r�5�������;I���L�ͬ?n�f�Wu723�&�\��J�
z�!&&�I8�P�J䢳)+�GYز�d7X�'��xi͆
�u��hܲ�V�ojax��P;�YH!�k��0J��悟�	�0�l�p<q��l�,��(V�AÉ�Ķ�ZJ���z�B�KI����k�D�Z��f�r$6��VF��u�]��Wn��F^)K*�u8���ܹK)?�P,bˌ&2Qq˖\��Z�NV'A�y���SsT�r�l*g����G��j�����ُ.ض�طS�j1�J�ܒP�u�f�	/ND�aD�[��ha:��-ҭOT�k!�[���]I�=�a5WJ���'l�7�̭ �uKf�OM%��Q^]�C�����Z¬I76�EM�Ak��L�(�f��س�Oi�!� pa���A`��^��%�	DI�L�s �W�Dd�>�7#�#u��x ֚qR�gS1���Z�X�Lݕa:��TǶ\Y(6�{dB)m`L�9G*�Rr5���/J��2�]���C3t0�`����gK���I!��·+b�(�_4��0��6T}z]70$@CiA�mLOi�Z���^#����#�kE��2<#m�U	���ԭ����WD��cf��&`͉`��V^bl� ��3d2����5�U"�J�T`h�l�ʽX1��*Y�9��up���LSF��ˆ�'a����T���\�ܻ��N�&�n��y�S�Qx�T�_Y{N�4����`%������ݑ0�mL�أtj%�f�)���('W!y��ͺ�*އ�*�9P'.n`�$Y
���n[[,������͚�Kʔ2�(���F�6����T���P1Z��-�Yj�%0��q�"C]�L�^f����1^c�{��c`H�d�B�Ƭ�dTh�[Ŷ�=�-Z�*(j�k&��\U�� @6n�O,��ƝlWf�.Ve�1ɶ����ZQrTua,m(8�GZb���<tM����0�)؛x�K�w���f2���kd (+V�c]��GS
�О��Xv��3j,�[�N^MӪ�id�tf�ky�`�HT[n��;��VR�Ry�c.�^��r<q��� c7Ma1�Ŏܴ,X��",��0��ߥicB� V�l@���wc/[����2�Bf��L��f�D)�f��In���mM!ٕ���l����{�`�tU���VǷL���o5�U�� ��`����GM��N4�.�Ov<�w5#�^a�	G��6�U5*�Q]��C�[��JU�Inκ��JŅP��ҽx��w�9M]5��,�M����3a�֫���D��-�(�aJ�vG-M+��R�L�ZM���[�6��W�+3V*�}��[I��t�d5uuԐo6��k:�'��RIZ`��z)��Me�^MFiM�2���Ԗ	��M<mn8��
�F�U٫�w7m$*R�e��b��űD2��4�h�E�R�0.���Y�C-]��+1����ȭ�V��#`Ϸ��N�:��q��f��	��G���<�L�j��L�(@��%�eSJ���ư���۶�41���N�ё�rch�p��ټ�Y������u��Z;lP��!��,r�D�L�r԰F�* q��LMdl�F^5H��R�3r�i�t��&��N��1q�*�b$�"1�un���\Z��'����ę��ѫs���b���1�c��,���I��1��Z+H	+���1��sE$�"ȼ�r4lF�Q�H
�*[��mT��g!Z��b�T�� ��1��G
�^����6�}f�yv���Ԉ���@��L�r�Q�7N�k5-�5��'���)5[��qk�9
AT�P)�pQqi��n㢆_��Ri:�N��#��/���/�.�iZ�;tiӓS����*���HFT6��H��G5fe�,]^��OHk%Bَ<�P\���6��; UJ����Q`�gR0Z�A��j�%J�\u�Ŭkh��R`�u�ut�n�e��1%�w��ԥ#��̏�R��p��F����̓c����r2�z�\����HN�yW�\V�&?�ݕ�#��i��1^-|���ݥ([�V �[�+�IA�G��W���I[��Am�/[��b����;���*�)7NP��J�К(�m�`�^��2'M�(��T4X;����se������+����o͕u���5�R�sj�z�Q�ەuW7�k(�WR�K��nm���Gk)ʽ�4cőa�23Q\��J2�W2�6A�@�\d�u�.ɭOa����7i�&�܆�6�h����F�!i��7.��%h��ck�G0�
��(5����ѻ��,F�rt4�̬�e�w�f���[i�tұ�`ۦ��9nn#x-�fC�MH�mӽ�-���c*�)Q�-#R��2�4լ6�Z����!��J�36�0sm�\V��Z�G,�tn�6e^��E�XA���z*��*d�`�h!z�|1-U��i���@h�+����-̨D�3si�B��$���iw��Cy�,%�Z��g +PHޅL�w@���j�1�6e���(�dU&����d���E�ne##�QR�y���k(�.�wWn�f�+`���K��&�b�Fj�2�֨ ��Rzz�e'�sFnH��[7����!7���� %ؙ�9�,�-vf��l�(	z,[�y`d4�5�C$����������Pa��Tg1DU��&�Bt�{��\�lg�d	��А��1��a �U3�J���"�+y1a&�]�h�X����gI���/f6�n�fκ˧N�a=�,ÓV�a�*mjՌ�k$S����1�����[n[͗��D鲎M;o4�1�Ğ��6��a�Cs$u�D��b�TuVT��`���(J�]I���ۻG.���f�5�ǸN�\�t|Y��U�$ X���p�c/r��A#%�b��hFVh��,��N�;&���Sˈ��ԣAa�P��e+���B���pn����Hn(�M`����q5����*���YN�T��jc׻f��eK���U'�[�b<8�O���/&��Z�z�+T���JBˑ͚���>ź6��vv@�������dUh�Pi��'V��kmܗ�(뫂k�@�� թVe;P�V��`@�ܧ��V<vj�ٛ�5aF�ӹr��IQn�O7+T�y����cq���sw6fe�p+�u��k+)Kv�ɕ��A�(�'hA_Bv�766�%)*��䕸�nT��Ү��]�8�[O-R��.���.M�%"��
�����	4Q�YE^n�˟:P���4�.$MIw��O/o(U��Rlsa�BG>��f��j��<�5G�0;�oR*Ww���ݐ���ZFKՁ��M,z5[�XRU����8`@�lF��U�"�8m��H3{��H�BIR�%;r2.·��'�[�tw7b�<�.*ѕ{y�be*iR̬�6��43"^�u*,���1z�صI-ժU�܋.���U�ᇹ�Oo>��i����m�M�Pam�@Y+�6��6��n$���ժ���^
�VԳ��e
Mf��5>�ɘ/p�B����zh@7n�ӛZ"�O�#X,H1Qم��i�kҹ�h �ۗI��a�M�wJ�,�@�{/i��D��*hy-��n�8UK��%�Dk��d�wI�,^�2݃I�4��i|��r#%��94�C^�N����;f�qQ0Y���^eR*r�Э)�2f�)�t%mis.����{��R�5��2n�W
�Ց	
M�b�r�-!��"�^�V���`@��	ԫcwn4�^���Z��պ]֓O*����sW��U&^�O�<A�Mi��ޫ	IcV>��Ъ^�Mk1��Ra�oj탕oa�kUH��ܟD�N�o6�Ƭ�Xqa�x]��� e�z�^=�R�W�fmc1CN!
f�w���G�Z4�7�ѥ�&AR�6.�A7J#(�Y.��*��6�wU@���D5e#ef9Wmr��N�K`6�,i�J��N|�cY��Q�+!�z�5�S.
d��i�NeEvM��#`l̸�52^lUs�*�^��l#)It�Q[��;�ȅQ��b���{W�;&�u��o�S�5k�T3���^�5����淑EB�^��$Q�J��^��4�i Qv�']Jw���F�Kl���x�c�Z�Vܭ86�Z��YW �����v�[v����LN�7H6^-H�����@ص�����E���ޭ�Z���-F��n��;j�ŃCb�m�zZۥJ:�v�b��b����L���6�b�8M���{I]�tv��2O���N�)WfU��Q2h��u&^�Z�b�*�-�t�Z%�@��?	���;��&�B�xEԙb�ةX�Cr�b��ڱYA��<�:��u�˒Ε�܈�����ڵKFS4Jͷ�dӳ^�l���E#��U�t3��۩��v)n
z�c'm�L���hh�"M6�KI���`��,k�ahT˙L3M�+t7ԙ��EF(i�t
�fH�C�)�s3L�g$ۼ��E��"l��<��t�&��n��EElm��	.�1=k)�f��36��r�Y����x��u���3y�jKl���i,IE��mc%��ʠ�*q7vJ	ɘ��1M. 3�[05��Zs�3-+�ǃB�DI{>gfe�h��"���$�7f��)�;ݵ�Ru��u"��^Pي��Y�Z����	���M2��\n��(%+@xV��s�Y/ST�	a2�9dJv4En�`8\ؖn�b�ƶ��@Vl���e�
�����d0�^źЭR�DX0ن��;wq�����Cߖlr�i�eB�+1���4.�Ռ����䩵�=�.�5 cc�&���D�UY[�R`�#�F��G�'L�Yݙf��w63��N�۽�&m����(��	����F��4����׆��u���:���7��Jܹq��2d��dt�&on��Z�[���Ij��3ڔ��M��훭�@�Zݖ��rLX�V�6٧O`I�e��#�[�p�q�
��{)U�x���ÄTǵ�KXn�f�����a�o�����9�z�*6�H��1�����h\}�I�o5]{
W5��d5�U�+;��xU��X*'y�x��<�� ��T���V���峅7p�u ���TQ,�R��ҕF�:B�HmlX�0�oX;d��du���Z:H��lM��.˸@�6ce,��/km+׋atH��'���;^�7�7KB�]�K������i�V�1is�Pö���i̼W���a]`�����y�D�n�Ohcur���H�2#��X��!�٥P�i�td��S�۶����m����(��O@T�)�f��ی��ɔVKb���3iMHU�#+E���U w��XT�u��Y�1�.��į+Dց5�e=ag-<�P��ȥ�:��WYt׷����mLV��UژZU�#j���l֮��ѷ���nk3$r���X]�HkvvC<���EbY���MC�b�JI��O��� L��ޙKnr��0%2��\
�Spe�.�o.�h�E����E��4��i�
���//7X�^mJ��ed��I�i�۩GuU��12� �-9b)&���Kj��u[y�Z�m����\���Ӻ6"�z骀\i�>.���^0/ThB#f�[HR�;�x�3{�<�$�j�;5e7�xs7�]nX2P�A\�ne͢�Vݐcj����f�\�R�G20�[�n��c�Q�{w�U��a�(G�i-�W4%��lw�{�������ūk��]�:�� ��*�%�vLkMʂ�Jՙ�f���DvQ���X�d뽒��	Pj�OE���]�[[@�ѭb�L2�j��V�%�t5����.*�J�,�D�m1�m�	k�Z��a������SJ�P���`Tp2*mn����:.�T�����Ѣ�Ioʜ�n;F�p���oX5k�r̂(2���cTw(�n��{2�m؍��6Ґ<d[G��=��M��RصB"dߖ��yY7^���A!L1�� M����0V�H`�%�6�h�V�5�Tk�q �;@+̧H��{���Ӊc@Z@�d���Z�co7/XQ�z�:f���5qen:�˿��<�J4r��ݬRB0T7���)J��� �3�)`�K&7�M�lX�2�6mla�XR�9������[�Α }�bU�qJ?Z��QI���O���g��M]�4�U����И��HwXuۣ��Z[�n9��b�^�F�Iɂܷk�yM=ͼ��J�#��H$���3Vɭ��Vc��]f�*M0&���{.���%�+jY��m�^�՚��v�U�m��boM!�CoEXWD^��.��5uz����ؑJ�[�Ohڛ��D:PF��[pP�eLC�)�[K*ɇR�MЖ��N�����$x��<uSV29��N��R�(�,�vjh�\#cZ�:��1�%X+�-�;D��%��V-pB�j\��x\�D��JU�o�֊��+�L��(ޤ#�]�O2��(�9�g%�w2��j��[�dʄKAa�a��,��(��q�q��0F�:�����5Vg��Ϗǵ>z�����h�v�5WN�J���g^�0b�,���lZut�L�Q��V�7b�[Vle�v��b<��q�(�jJ*�,6�㏲i�ڹM��V��׃O 6�#f�����X~����n���NXm:h�s�`;��-��'� ��zƷ���T/[�:5�S/�Q3s�6K�n�u�"����i.]���2��}1��v$���1��-��T�鮻7�MzxB��sY=��e	�r[R��i��7*Z$H��K5�]�iqӳ�_N��8�v�n��y١���d�)&[s�k�yF�{
��2)h�6���un|�������,���j��M����t�7�J΅>����(r�e��a^r,�Zbɢ�${�H���q�omG&�Dj� `�"ޥO-��K��O�h���^�B�'"�/o~�j�Ye+ɂ�W4�A���CCY�5�!����
�8oB]	��[�յ;����=}M��ֵ�oD���/ҳ��]q9I���;5�Y��$j�+Ϲ�
>.�L�cku����Ix�|��R.l�u{YJ�X�)Qiތ�Rg�Ac�j�.�/�����g-ͨ�\z|L*xd��>�[����d\�M�
��[WX�m�!9ST�Ҵ��i�YG�*m�ָ��gbc�ܙ��ڏffEs��@V�d�ՙY�9�W#�]�x���*��
��� .7�{��B�9A]����Z,J�>�GrQ�Ȧ�����uAڸd�]���Ay�TW���u(��R�Q\����hq�;�� D6��!���CfD��*�;7�D��O���Y[[�6]fVR�OZ��'bw$@!������>��`�{�3Q�/9l�Z���G^t}NʩQң#��v�oJ���!݆� Z�Re������jc���y�8j�� 6{c���FjG%�g_j^R�l����_}��+lpS7�{glw[5��OP�.gn�n�:jlݣ-�ltӭԬ��u�6q�;jn���uy,|����)��4u,'t��X\��řv4�&;�F�[KM��ɰ��W�*�Q��]Jĳs���C8n�|��P��:��*�\eިN;������S!K�֤}�ڱi�3:�[f�*Qm����$ށ5W_O�6�pȔ���3NZAFTuֳ�+6���ε�ѳ��,��b؋l��*��d�o�,ёe(\�,䝃{&L�|Eh���oWNϔ����Wk�h�ί��n��yF�3W �6if�����30L�;��yK�h�k�q�ڔ������}զ@Z��k���z�J��%]�ط�({��ΰ���W�«�ǥKp���#����,aG
�ϰ�����,�$�8<F����f��k�KQ�l!i�ӕԬ��U�@�"��m���C����e��-�й��C�$�z�{<�*i����[w˩n|�h�%��㬭�	i�M�Ⱥ�f�������e�{]�"�92��I��j��4Cݭ#���b*t����m:FZڼ��A7�y�7	��X|���q�W3
�;:I`f�4r16}�Y,Ds���D32��̻ܚ�+Q�p�F`�b��k4bK��]��ev�y�w��R��v:��b���S[�wI*׼�.�η����^��%�#x�4yt�Od�JV�u�ԥ�N�ם��b<Uծt�U�LY���]��֠b��wem�7Ȳ��}>��m������Q��-[|r�Д2�d���ڶ��&eKWG!�����P���Z�c�QH{maa�x�S���w�Y��1��I駓u�L&��c�Z ����gRU����R/��Q알)t#�^�u��JP1���ᇞU��S���RZ�Wי��W�JL]d}]�)��Ntu�U��d��R�eZr=��3��ɠ���Q�δp�;�,�Ф{ �Y��\�qV�M��u�v�gVs��;�g����Q�\�R���f�W�o��o��Y����V4�jT���5���h}wή8�a��d�A��$/�i�s۔sa�����Fg=�.�ZO�Z�Ϋi���wD�.���u:�87�g�R���^�nL��U֙��r�����r����.�N�m���[8�O���-������*�콮�vm�����6WJZ��i?�jP�ʆ��Z�F^#Z-V��CAZ'%u�`#��m��I$�L�m����S��;#�l�v�t*q��s�� �J��9Z,�nTɡ���"�e�zi���wc�6_g=�"����t�^��V������D�&l��O�C��K�S�l��[v�q�֜o��G-�Jt��Ǆ��$�i�*o�" ��ޓD���'�X��.�t}V�B�3���m�v����3���ErZ�d�eL5�W�,�Z�<�٫�寺�mӸ�z��R��2��b��D���[��h��wc���7]I��&X��f,(!�;)�2�œ�)O$ۉ����d�2�ebk,b ���v�.��8D��'\��+�����J��n;������N�ޥ�r]͠"�������}���\{e��q_j����o��;�w]!��M����ݹÅ��I6��(�-�^%Ni[,�����\��J�.�;�h�/�
I�m���J���Od�J�Y�2����:݊s�4�!��.�+l�MEM<�޸�Y�jb/��A��7 ��4�ΥF�kq�X���ws�6�]�jгe��|�儖���4���v'gV�NgqW�~w�Ŝ>Ԝ~��!�5}Gk6T�x�Au�3K=��]�lj�«S�S)oV��U��ɇ_1XsB�O>Gz3*��K��b�#I�M�J=ú�F&���:�,��a����J�*V]6��j��Ne�.�+���ڭ˓%Y�{)V�V�
]��YUssyq��
	�{�#9��I��@�r.DRx�v�MIY�ugU��hͧ�O���V����;,�d�7pw&�!P��P�Z�Y���P�m�����H�zf��d\�nB���
��"�Apm�W.	n8�L�|�dָ�cr����G�&�D�gf���f2"˰6�Hh��9w[��g+��ݥ�V}.���o��M�W�gY�hg�XQ�glX6��NXq.��9]^�#��˱"�7�V�*}�Ou�u3>	�����&�	�j�K2��i�m�v�2�T��Hܻ��v�ս)�ȯ�W���Ɇ��5P.�m�"��k%�����p�z�J�`4�F�@�c�lU�K����L��*F²s0�<��3��ұ�YsR�sy]M�DT�jm��+���0�J��%�me�qc7�k���2ki}dZ#���2E�&���������.��)Z�\:L�S6�t��֪��c�촴R�}���8�O���5�,��'v*W�A��9S��!���1��6]�&U�5˰+��b,.W��b�7�ۯ�7�2Z�.]��X{-�!���;�h�Wl��ڹ#}P�9h��m���|M�˺)�o���@�!s���uq��*�:�˄,���Ƭ@K�)�� `��6Q�`(��Ԥ%>�|;s�ظ�b���r������a�z��4�ن�Ϧ*Ȝ��ST�'e�.`=C��)l3�D.�NwS�J� x�Mw�r7�l�q]���$��m�kȋ��k��N�I\χ�(�����F�&�ͯx���^4V��[1�E-���a����nmfy�x�B��k:�R�qޔ�.�Խ�S/�ݗ �k'eguYע�ޓ��+�T�j4K�Іƌ_^Yʶ�q�!�V8�!�u�л�QZ�k�jZ:�E�e΄�����)�D���=ԙٷ�^�@� ����(X�p���ef��hM�1ϻ���D+��9��j�8�����[+&�_a�cz�"�K�<��z)\
�����fQ�Q�bu�q\vTG��g8ހ��b�F��M7v��]����n�Aj���7o�N�T-���Ю!;Y��U2�Vd'.[��#i�F�bN⍝����!A�6�vq����#���x�G7���9hxUͥ��GWZ�m�e>֒N�n��!�q���.�vf챪DޭO�m� ��F���������m�I-K6���������V;ۿ�%3��;������:N����R�^�vIW��y�I|f*���
nS�x���̷6=�
�r7aص`�v��͕o6m�Ol,���oyl�QJ�5���hs���4c�+��{9ޠZ\�7_�\�:��6{�E}�d�;E��D�%5^t7$�h2<l:^%T嚬o:N��!Q<�&�^���0+F{��]���5�Y�rT��P9V��Bq��cz��8f2��� ��w�Q8�;�fm��7p��B���:���'qn++Z�G;zb\�F�Ia��+����u�.R����.�]��E��t��3f!�2P���v �R�GEwV�!�����ԍ��A��B�0��ټ��h.��v�W]q�"q8p�,]�6��k�p �'FC��^q�\��$�7�p�jj>���\�N� r�*]6-R{8J���S�K�:*�!���owa�!wi�E�U-�r��جR[$��EHsBi�fQ]:і�'fJ։�6b��^�nX@� �@x��WZ�纯�l`��T�����a����8�K�Vu!W.�]��+���B�an;��nI����GC�jl���c�V�ľT�J���X��q�ivNz���N<�5�iT�m�}����d���-S�]��[����������玃A:F���J��o��K����R����8��E9�a�N��k���B�S��]�/�6C��d�����xƮ�u����{,Y����3���&��1�Nl�����yi���/:���tGRR�X�ѽ�E�IggIN+�����s���;ϹZ�f-;ux���X����73Z�ڛXS=��Y����2�p�йYP�bŜ��K��H�B¨c�v��T�*�֚���a
��r+w��Ǎ+�V�.͆2pl)j�.m�.�n�i"�0�r�eT�]�1n�J�b3*ޙk���Ucu�mʋ���-u��&���;/�X�:�re����Q+�I^��*�~�o�G��Һ:W��;�޼%*]�Þ�yi��-#��sl;|����Z�/�X�K��H-�J����\�[��{i��Ό����������J�܇�VP�^6��2sX�)���n]�X�n��n�����g�?��GG9�Gh�=�E8|��z֔́Oe$k*��U��J��Jh�I��aU-�ڌVq�n��Ui�x���V�RJM��Z��X�:A�k�ץr˼��z�{Jޔd�y=W[7�5�^�DoV��ӹ_c����6�h�4\4+�gT���busJo	N؝@��)�q��;0ݾT%��ge}�Ao����u�8��t2�"Ľ�]vՀ�grUŚ�������yx��B�i��Eb�]^��z���^q0�&;�u�R58�7�#l"���j�JSBl9n��`���.Ns{H�Ī�ff|�՞�/*�n���7r�q�J���F_|O��f��R����9�����в�f-[��J���V�U��H�4�Fqr�p
.�V"��x��)顺.��O�P���&�v�!�v*ߜ�Z�R�9��f��M�+]�UN��L�m�I8f]�g6��E�����;"�h���ob��L錵������s��St��}���W@"X����Mn��) �k�<!"���cKq�L۬Ò���Ea���h��t�AV&�����j_t��K&�b7҂�^�m�c�[#����vS�dg�ʕ/QȌ�VQ�m�e�؁�ܠ��\+�%�d%rA�Cs1��D���"�G�`��T&]��TdX"�������
���r��ǜ��k���-��R��1>vFvlg���tᴰ#Zt����#ί������K^K��[+]ǳ��9����u�3��������M��ָ��BÛ�z�5���G�������2�b�7M�����wk��Ӹ�u�I���SEm%������t��od��-Vz�9;E����\OM��ٳoJI\��,�y@ûMܿ�lg�[b��}�c���2�FҲ0[ހU��[Xȫ����jf�&��T�����m�cծ#��(�\1q�9�rT�Ή�E%��O2i���!֟u�oŃ�5})G�VZŶ�G�w�ߓe�������e�e�p�Ϋz=��w�\�|��1E|�؏_���iK��^,w����p�b�c�4�_<�f֕OxPV�p�Y���i�WJQ3�\��ǋo�k�X�y�e�����;�a�#v����N"�T��h[7Z���r���-���a�nU��9�f�V��&r�v �@1ŵ6�#YΒ�R'���c۠xTw�P}��2��xV����ӓ�'(N5R���.gYRy���X��#J���͈��)��B�k�g�x�g=�N�Ph%��\�R\&�teQ���
�i��)-T�]�Bŧ�K�f��)��F,4�t˼�o��/Uƞʀd/�eDv�c�<��F�-��jΪ�e*�?�#�2m֊yq��"�]r�!9�dqY{s6[�X�d���1P�}15�͋�?H�{��H(�sbd�fMV.�8q#��Ŵ�m�]dR�%6�;X+�m�Y�%����� �$�T���Ӭ6���ۤ��e�Wh�s�G7'��QQ��,0��a���:t#��s��ȋ�$mcxY�u1����SJiv�M^�G;&-�D���c{(l�R�\�̗�u�����.��y�:��^K�'P����b�]�|�ۊ]�ݮ[���"���>��ےT�Ӡx9B�G�s2�RAXJ����sN[�|n�맨�p�g ��T�+ov)h�R�]��:��q�;�	����S6]B�9}s/�50nP9$R�UW�}UZ����kj����j����������^����ߛ�v��T��nI�jI��+e�����2�@��ۖ���%����WQ�M�[����(����sc�:��9�	R�5y���n�p�&��6Q������Ҟ�Yz��l*�=���2q��[��Fb=����ZX�����903G�9qQ�1�=�niR�NJ��jX#��T���@!{C.�K�h�2��{���۰�C�S0�i�����o�r������f&&��؆b���V�c]ɉV�MWV^�}�چ�Bm
n+
ꬔ�oX�&��b��Sy��ŻdU�*�r�����ptJ��	u�5�����3i�SUF�N�yL�D.u(��П
7V��R�"V�tAA�Д�t���\Օ�6d�-q�lY�WzNEW(̔�tvs2�/ef;���u��
D^,�\֠77B���:���R3}.�he��t];5a��ɖQtŃ� M���Փ�-fH+�^)m�e��GVA�1���o*h��h��.p��:���M�t}#�Bz��z�_�nL�t����nI�wzcz\mgn��":J�4�a��P��d�Ӣ�<2u5yc�=��O�e�aUp�K��Č1Zl��I;�ݯ�m���K��[{I��c݃���	�&�e�Cf�U�a`
˺��e˼��7��9{Xj�e<�p9�l�\������*�V*��&ur�̭�bM�C~�Q|��J��[w�uu�&�(n<q��gf�7����
��4�^k��f��cV�7ƚ飳��J���U�r>�2w.��vV��|fmn�mf�=��w2\�e�3�t���)_aN}VPh�N�ܼ�a����>�-�$�(i����i��:�)6a.��-$����zb`��٘��wR9b�ڼ ]�JU��Ya�uIӷy�i>Y������L.�\�K�K��W�WWz5\��5��#��D-k�<ϓ͍)׶��fH0r�t�Č/�ӊ`���u���\��v�^(�{LH�.��.���2����S��k&���[�I�yW�S��v��[�ᰚ�Mh��J���4�.�o��.��+��1F�i��K�2�\f��T:�w4q�أ��2�mX��Y�Z9 n�-�m	�\��^��8�����_5yLKW��2U1Ϫt�F��F�k�:�٩�Y�SQ�N�s�O�X]@�;%,�v;@;��o'2�ĸ�3h�8p�w�rͦ��c:�Ҩ�vWn�7cie���jX�ZR*޷WQeZ���Xu뗺6�U��;���\�n���p�Cv�6hU����U�.*`3��A ]t:�7[YD����2��w+R�mv�N�P��r]5e�S�D��^�*��_[Tb������~���;K��'zc4�Y�b�-�r���^��N�-t�H�B���fnS`d�zns�r���6����^]7�cu1Z9ܣOUK��Hp���ܾp�9m4������ZeF��#��A檤/6����K�����	,a��k����]�;u�E+��ӓe@]7[��w�N�1��-�X��Ԭ.���	�<��,�.ŉX��n�llh:ݼsRQ��Zڗ�ۙdb��x�I`ԼϒJ�h��{.Y��fI:=��2šP�IQ�k�)M�zq�jT�2b�{u����ح�w۲��r�JҴ�vgX��J�N}x3��t�	��9�`�\k��n�0rp5b�b�2�ws�ң=�vG��ð';(�	x*Vi*�sG躱l(;��KoUMGx�:c���˖HA��_�E"Ĵ��X��R���<v��F4�9�B6��Y�7ԍr�7�J��Z1_Ik��lT��\�$��h��h��D���|N�np�Y�3nL9&��h�@( N���9+2ms��li!�]K�(���*�Hgm]���u8��!\���	������.j\f�'�.QU��L5n���&��N��hN��o��M�b0yj]n��Ks�K�VE���0rg�:l����ݝj}1�`�e��z��fqA�+b9H)�/�tĬ�<}ظ�N�X�r�^:��'@3���mK
J�lh��T�Gr L�e�Q�[Z��Sc��[C5M�ݘр����[�`�9oS׶��7O"��a�	]7+n`�
Z���si����"��tU.m\�������d���S]��9�+���r���B�\l�#YKu�J�[��l�^1�i՚R���
�#B��4�u��V�x�8���ò|����|~V����w3��@�i#Rʔiκ��S����܊�h���mZ׺w���K7T�<'���7Wj0�gZU,��;NJI>,��N���0�mnL�Ѫz�쒹]�k����{[��#��R7Ԋ�k3�j���X���x���s�P�u�$2;y�s7eE���2RO1M�qmvV��Y�����t�]m���e;����$�f"�]�F�R�]"2���2�i�֨�'R��}So��3d�L��l�mLu�'�I7���-���^f)��� K�l7t�TOP%J#��j����:L-ƹ�V3j��<,8�����uwҶQ���T��n�P���љ��u��Ø{���Ѫ����΍����"���]%����u	�˗���wݼ�%3���^9X�v�=�*�ۊ���R趈we�JY���9�*�}]C��L(��A;}�}>/�&ݑ�ѵ9աu,"r41H���̝�MeV�{X�B��?�#[R%]����-XS)sw;u����p��i]u�f0u��ʒ�ۊTe�5�s���S�W�!6~���Iَ�v �.���P��\J2]H�!��K{����O-��>�<ā�]g��̿�Ƀ�)�6�����N̪�n�쵌N�%�X�v���[�yh#�J�`��7[4�j�2c���U�ҡ]��'��d7��^�ߩѫ�����A�-9�pTН��VhMt�[S5j�M��|�kz���q
쎡��ڝ���+%�&ڭ�v�.ٴh�:�1�x�N��:���7�՚Qz�Lۛշ֐غ�}�|��V8�J��7|{Xٓ.5�r$L���ّM�fZR�2�.G@0���sj��u����	��wf�K���ؔ���:4��<��T����ɘ�k�7����e�$���x�#t���Z�:���p�Uݪu4~��.�Ƭ|ŭK����m5Fv��ܽ�&�օe�ͱcvQ���ܡS�m��� �U���
��Z`�؍�u�w��I,�����)];����&�3*`�y��ݪ����ҐE�>�7,�]�����x1����pP�R�M�[���&��O����se�V�9�h�N��N�L�#��N��`��g0�Qs�5w�2��`$�$Yr�6�>�d��E�N�P1���^*�p��*m�g���idqX$���1+ݓ���K���i��ǹ��U8�fs.ne�XXWB%:P��:}Y�\y�M��r�6)ŵ��fLge�qfKF�c�m�M��}���w#���+BĚ�x-r�;�	�z
�oTb�̜v�:��u�ܩ�Crw&f�h
-ܨs�;K����A��5�w��@�;d�y{-��Y]`2Ewf��j��R������k"�$1�%�2s�ؕl��0&<
ٸ�f�kq`P�>�f!�^�.�H&��B�T��1W�4cXtĮ�MOZ�ݠ��v��[|�e��I�7Cd��ߐ}/��ˌ�K]�k�z���G*���Of ����Y�����M�v�v��rUӢ��x1S0��m�n�U�l�Ճ-�5e�x�h]k��V��������N��X�2s� h�lR�U$;Yx��%��:�N�:u��)���F
Բ#K2�"p�uy)��H​Ye�.2�p���ӱ�X������T��%�.�6U!�]��um�I|D1ʻH�D�E���?[��2�9TZ���X�F��ϲ��lM��o�=��7J������ЖÂ���O8u�ڜ�aͬ�?7�f�i�K{�T��(	i�u9RN����=��@����S��%7AY��O]�l���Ӝ�Wp�[��9�9�wo�mҫD��[/E��yJ�ŕȽ���y�5������{�v/�ҳ5�+�o�^S2���1RV�v.��v�n������5j
`��c(�-F�j�gB۝�[ʓ�y7�h�(����Gd|T���]1ͭ�"�-�#f��Y�X�-=HU,�*EV]vd�?cW�f>�a�����r�tQQw	��>�p�{sV�K��x�١5q���pQk�*���z�7��dS�֊V��{��r'P������8�Uz���qΝ�eͻ��U�r�Z\y#�t�ĉ�vmj�Ak�8�FS�� k3�* \�]���|��yG�U��	�.�^�P��M��Z �`7��PnΘ�^��&�6ȍф���+��G5\kŗ65�
}��9rI�Wu{[Au�ck%�\�z�@���75�ۗe�wG2�FYjl`�yNu�+��`st��,�(�B�㱳o�V��.�ך0K���eJ<��^�)P��v��lU�\\6�n�u�:ۨ�!�kp�h���Y�)D̊��'AW��=}�m�4���+XoC�
��f�RI񐡏2���#��7�	�{���i��ʹ�b���mT0��m {_$�R]�ٗLO$��W�~4�tR�����J��EC�eN8Em+���1Z|qhV^��-X���^$t��������F�:��׎�ko�Q6ͽ)�ts9jĦ���q�/�����/zwmK��):�P��O7���i�T�_]���lR��7���y�[7�cq[���%!�ιr��(Z���
fk7LԭH݂m�'BD�ic[�ŽtW�thT"-���NSTQ[�����mv�����0X����GIQ�ȗ&*ĥ<��w�Xz�pTi"U�n'����T�3���.�Ы�m��#����oo�,SPs�Kw-f݅\��;����d��|k��%�ȝF��	�,cA-K�YF��k.����d=]%	�镛a�y�kPW���Y]v�p䦪^)���.̀�svL�Uݒ��ԉ�fDRI2�Ի�]���v���P�/����}g�-Xɷ�Ҷ&�il��zt����Ki�I�R�X�1��gH�G������PF���� ����V��9����R���ػ3�1t0�v�O��IwfvI���:Q�þúD�x��!!��6/�as6�=�&�WX�w�ꢵj��\�gl�λ�K�_)> ��=n��k��R���2V˚�g[PˊX�%���ʨ�[v�k��i;Rfh����іEc����1]�Iyʵ���	���\���1�}��4����Hԡx�co;��:9V�Ș{��r�i����^���\�~�AM�k9k�tS�h��֐ԜwP����0�-�����3q�	8�^+��9"�Rj&��ǽntw��{.�rL�1��[��OE;����oo49׳z�=�@�V��0C��xYW)d�e�;B���Lt�}A�3���q"֕H��ͫ���]J��j�uŭ��Շ�:�`�NR/z��>�lP�a��!2[˴(h�׎�Dp��� zEH�8�GK�C�G��NhRa��U��;6�N+�V�x�^�Uݳ������Z��2^E���Z��bjm�y������K+l3��U�'L��WQ��7��OT�n�d��q{��F�q�!f�T7R.��WXWAeޢד�A��\��<m���c(���#�Hg$����c�j�E_uX��'�N���p��t���J�����ֺ=��/Z�9�]#�������w$�oA�HLK'��4'��e�s���Q��[�UT��,�n%���N�[[#�'��S:�I40J����^DU�J�Z��Fe�SlX*���PP�-�Oa�]�t(1�,�vB6�sZE���o��Q��5�{�Q݅5�G:%͜+J�]s���δ�J=`�AI\"��C.���+@W���Cv�@��E���ƥ�T�!��N�p��4tq6Wإ)��*���YM��yI9�Z-���1��Դ�����/`Sgr��g̮V��c�$�q�8F��3���Q�h�M]���h�Bohe���H l�J6�py�pި]e��>��0�|��}}�!����"�9�����Hޱu�p��8ͥܨ�k�MSTQKA��-�D�."�B�󺊵%��g+�wM4�TL5.�M�4�k�C����f�!օ6�����Ҿ�L���)j���E��AТ��9c�뻮��j��W�x��Q�`b�Uh���96�{L�t���;�pPe�w����(��nX�Q@��2�j�#�qX@��C�����P�C8���wi�.ñ�'ո�*�E������Q�v�oG��o�M*ڍSYyY�/�of��(m�*�h�����vm�v���EI�-ɓ+V�ۨ�TZ����X܃s�xy#�d$���`=�N���ڜ*:j�՛��֐�c���k	_+D-� ́)���8FU�8�Dbj���f̒��9]v,ܺW��Wk;��<�����0�&p�h�&9)��Иju��:�;B�O���n��eԸ����s�)N�T{��9U�:@2M�����n�����h5�t�����\@5�s�5n�jf�{t]m��b�d^��Jus�V47������L�#x�%�Б ��VF��}W��2�9]PC)�*X86Q�
nͬ9�K��x��4�I*�X�;���3*Ōz'B4�/vJ	��a��j�� �ʃ�!S�������Υ�J��o��� 7�j�rb�r��+��:�ke+���%��:��	۾e���ҽ
�TJ�V:0޽���hcC�8�ڐ��g.E0�d�v��YBv�;PguW��Dz=�W���X�,[m���EE�sbob�Z��kj��|H���.�V����ٷ|E�#�b}��^W�qVw�>�tߖv�?���J�إ��
S(�rt�6ج�w������/^I�q�Vmj��U.�mɯ;w�4^���#j^�<����Ȼi�w٦�M���OKRa��M���m��U�D��\�c������}�9Lũ�;
uU�a�_
K��#�/`=ױ�/e`���8GJ�\0��iAI&~h9�X��śp��̧�}�ԕk-���e�Z���I�(���U't֤ͫ�;���us����ƯZ�dTԛ��ާ���;w�u۲��Z+hl�l��퐻�T��)��fR�����6����}F\��eB]�ht�s/0_*�q,K��L�Q�g�w�ML�e❰୕G�n�ݽ���NHg���$�d��C�*��>A�ά��d\��+#��3	��]�ׇF�Z���L79%+��8��n�VV
�'c��O�u=CS�Q�ݵb�,�8��2%����!��PY��[Z��a[�
�L{i�,�҉�	�Mu^����W��v���`h��`�զ�.���6�e�i�{ 4��z�it�u=�8�,oŖ�]c�3�a%��6yz9�e��LJ�iK�h �/gWF&k"�wnmjmaX9����W7YⱽJ]��`��ߞ����7a(C��8�wQ�s���w%���+���C���%�%�ɂlJ�2I��GwM
!.k��c�4��p܌w����I`I42M0��"C�D��nI&��]ܥ3���n�i�#2�;"�Ȁ���$su�sX)��
w\�h�"k��Y�˷v�GwI�0H�:4��L̈����N��1!D�M
S��g8��s�w\(��I��Uƃ�&i0]܁�4���� (�rt!"ŌXLSD�&"BIL� ��݌����Ā(=m�5La�
v�<�3L;*kw��'gV�bL]�u�J�J��lGz�EQ���9��湒�l(�k�i�o�*��E�;:�!a�"����+�F�f*_i�5^wm1YMŵ#� �
��n&�5i_7��7�YO��X����3�_U�G(��{�Ď�+��P��ν�G�hZo@m�3��E��}R{ ��
EU��=�qѮ�3�`��c'�q:J!�삧ӕ��s�J��Y~N����kN+�f�pV�^��b��ZQ1�a#'��	��w��fSIS��o8�84�Ζ^���C�wQ����ПS��ifݢ����q�i�$�[�m��VL��Ce����2\��� &#�ZfFB�����gsԫ٦���n�NΈ��j=��W4^�%M�h
����LNg0}�d�*-O%=���Ic�w�^��|���Z,��~V�]��˫P�����tW?��CZ;������錚{ K�!����2��~N㑂Ա����a1~�'I�.�z:�iq���T8�)t�jӘ�deԚ(K�}k�z9�e��!y�P:'a��:8��(;~6yq�[�<�i}�s���Y#�6�[Dg7���Ȓ�.T���I�:許f�{�t� v�vvf(ǒ���[��n�v\J�Pe*�>�0V��g n:���� �H	C[�B�$�Mh2������j��gc5%1�Nf��NF�H܎�V;٢h�$���3w�j�wb�LR��|��uY�S��9c����;��.�x�����s�.QIe��P�U�j�oo=7��@=0�Ĵ�!�������,ks�O=w�>�9���N{^�<�A�WBL���n����c��S�\��&�-�&/�ņN�A�^`��I[������&Ձ���׌c��ȍ$_�m:3�#��߼1z��2�NY��u5�L\���+Fs}Cπ_�X�"���~@����+�Yt�VN�+^b\��{Tmr]*+jD��혐��2d�m�=���pՒU}q��()�<,s����tPU�ZT�����0Lҁ1��T�zj^\,����|�QnT��ٿ�����"���j*߀j���л�Ɔ����1��ӂyΓ�(;;GS쌍N�Z��{ప�lĥQS��K��t�7�(�o��_E@�멇��8\Fu�^��.�q�n���d^3��7}Q�������4����Bwo�ag���Z��x�����gu�q��'�C"OȘ��G[����K��O�@�y�,�JK#p�X}��������S�S��irw[bq��]s��o��^�J�0����8�:�r���2���rcS��Z3�$�WsBεDZd�^���ą�;sB�R�^t��2��2n��N�B-]����hR�hz�ڳN��0e��aek�����U�7�z�9���mG����!�}�Fk���u��1�n���8)L���Ф����$/]�-<��\v�ҐL>{^�X!��Yq�ee7~��x��ȃ�����p�ZO1v�wgl�Rz+G��{L}�t�����>x���q��Z��(G *�i1r-�0�Y�1����'��D�����u�w�Gz%�.9�4c"I·�]0x�d�+�0��:��z�^K2Rp.O�,�p'�*�n	�ef^��U����7���2���A���o�q�uHT8���RP�J� c 1��;T�|�����������ޱn�ޥ�z{��#��Q��[n�w$�ȳ!@��b���ew��.6��v�S�y݁B�'6�GI��'��ߡ����s����`��"���QJ��U��kG�g������l��8���É̄�_�'fM�1�
�f�aD����jn��R��Ј�X��V�o;��v��&_D�ᾷ�J�k���Q����]�zW���nf˂���:��I��aVYZ��*4�}�"s�Kă�z����Skv�Sf��ۺ�NX�g\�&-~���|���6��<Q��V>��z�T͓i�ek���/I{����MdOmF�Χ���5uW��I�п�s5ܰ	�lz��}B��QO���X�����&V�B�?:��m�½2�[0M�7�U1��fU![w&F�����Ox�q�AG�ʘGm
u���ls7v�\VSF�S1�0g��m�a�لOk�����=r��ś�d��/]�����s]t�p�DfOӁ\VUi�T�|J"89��Y�M[���3QV���u4�dȌg[�����U��̛7�Ip�A/�܍�T4}3/}^O�H7�F�(:���s�2�W�E{��X=Y�/�-��ڡ�G�G�
nk����̈/o���-[���7��~˸+*Ӡ��������T[�HE�r��s��7�Ҡ;5�z\���o�/�������*?L�>��R]��^>����h��W���M`vm�޶�9;��W�˛��\�k�$�}��¨��H��WpY�/O�R��L�w)݀T�Is�dc��!i�=ꑶ���I/i������
�Hf�LЙ�<@7V�¶;�#���o���]��(�Ŋ�m�i��*?���l��<�6����2�m�1����잺f�)P����z*���7��Xݺ�F;0��,�G�ף�`tW �%
Ҿn��(�ޘ�RB9/s�h�h"dB��4�4�Ggvv���Rv���f��\Ύfๆ;NCrDmC�r2��O�T�!�K̅K��7��g˞|����q�t�sx���4���g�;l�D�Z9�3"��Q:�Y��(��t(�&�2��4�WS�9$?IǳB뺡���qx{*�aZ��c%1>�T�$�ө�:������\4dܛ�cu�Oa���
L�\b�7�q��b��>��2^,s@wg;�*4�F��j��~��)���DU��8��lnG��}պgL1��P�v���UtF+֪n�9Ym�*\� `~�<���X�gÏ�N��#��C߳ؑ�W�2�1Œ��ݤ�>a�MĔ#>�Ӟ��'���˸��
�e�t%��������D�+����a�������ȘvcZq\���w^�f��b��Q�k����*M��J�⛸w �='�!�ی�`W�Z�cS�b2"\��������4����xe�����&�f���p5�T��l�1_�!���23�ӿ�3�J��FZS��o����#�]��Hk�k��׸�2c\���*�n=&Q��e���}�DN,%*f�Ѽ��g8Na�v�i����jE��>��R�ϸ9�JpI=MY�=/��^
����v�2�q��2�����N�h*���������J÷K�Z��m�&�R�/�~g�����\�>�R�@wJ�)��,���k�3GX�w�:I�ڻ�+�\ޏ	��ʦ�C.׉:]#<Y\�"�@РV��G3���H����.�U�.�-��fR��NV��ɉ�'Z\���\k��X�yXm�絝��%����>V���e����sڃh��P�Yt �tL�j�Ӌu�c
��U��a����*�g"��X�c�:�+�î3�9�!P�(���n�;��1d�ԙ���@�pd�3I�<��#�9с��W�6X��t����x�Z9\��*�p�."A<����xw�\&WM�hyRźD��1D��\��H�K��h�D�c�y#�;$O�m:3�#�ܯ�TkF�&�{q9}ѭk�X��k�(�&f(z���]q�W7ȧ�Gx�ʏk��:Ϲ�<ڱЇ{�s����eY]�^pڨ�h�&O&���؂�&�*���1�c���5u�ʇ�;B�L�{���
/iD,lC(��TmK,�F�`Y�l��zV�̠���Ә�[�8�)(,�L	��hwWR��'�'�;qH�}�V���:"��	g;���7/�@#�\���A3�e�i�fa����`\�C��c����G�U�=�z�״���Z����̛e@9�������3@9M��T�� ��.W?P����8'��1����;GKێ��q�����U<�b任�;��s3��U�Q�mYSj��GB'1��0º�zk�����Z T^��.�qnu�f&+k�;�cs����g��α�B��;�Uv}��J�`t��1�1+"W���dp���䒰n�TN���VMW]�pU�k�!�i��]��������U�)|��p����<}J;��lO#ȭqn��Y|c6��8L^���H�`�΄��)���s�[m<�A�S���1Yμ�#K�`2��R<⛿u���1�D2�c!i����k�g�i|�����]��1�G��)��;c׮!��0�m\>�8ϑ/����`������v�P���'�,�Ex��q�����o8H�r��ч�����[ݩ�V&��+�=XȮ�G��bх���]A��zM�MO���;��]/z�
�vXVx����v�����'���"N�~���=\w���2�g���<'�G������r�LVa-�`�g�ot�P�R�_<v��js(M��
��dx�ݬN��I�I��}��q9����26^�ΰ���\jբ�<��ۚ�gQ-�9�pB}��ͯ7��&_2 ���x|hɈ
�>J���߻��T�ݛ�{�Q����5�>Z!���+mց�s���W%#�L D�b����O&e����j&�<9�rٸ�<Lc]NOD71���-	��HH��0fc��d@�Ε;���9p����9S$TEi����7�Hv_�'fKf#y��.̓ƥ˖R4ܻ�{��u��M�j�0v�5#��7�B^]w�uT8&C�l�	}$V@z_19��ރs�{[�r�t{v+�x��b�����/,¡�^�R_����ŵT�H`�4�X����8��<4������W�t��SV)C��o��WG��o�`��w���m�b.��o�E�Q'��'��n��ꩃ�=�
��m�iU3g������R���GN̎c��<_L�,j��3̢dF"�y�R�
�5���;�w|����=�w}�7�q|�Is:-�c�ϵ.Xچ"���X9�t������1~�Â��y̯Z>HT��r���A�<���پ���MWi��q���bv�111ļOz�3R]OC_.��M<!�B�@��Õ�*���N:�֭9Jn�]���p�R��N��6uu#�:)ihU�� ���)7Y��.at1T���RV8Ɗ�O<oF���(]L�:�"�4��������nS.�lyүO$��دb)�U�������^�ƴ�Y�+U��*>�JCt�C�T#�n�=q0�g[7]p�5k��e6�~�����+Z%�F�>$�?Sf�V+�U�v���#�y%m�K`a~���R{m�D5������Ɔ�:�$���(	�
a��(����l5��k���ݻjg�K�έ���7�1�q�"5��i�2��8�K����[�0𷛺�U����E��q�[�ò;l�A9���f0S���o��C�<X)���6H}��B׵�$LI�SB�\��
Xw�s��Qu��9j�0�Wy��h�OLk��B�[7%�U_��g�M9E�09*�W���Aߵ���'�ҦK�O�7��=V���!7�^�@?'PDM3	X���vQ���^��ڂ�����5Y*��葓=����ܓ�E��*�������������ug�#��3�O�_}�En49aB؂���E7��T�|+EO�ee6Z�^�~�ʶaQŢ>�s%X���p���sPUx�mZ�,r�+E��ՠ�rYI�jѓ�X�����q��F3Y�L[{�H�u=ד��'X��r1gv��Û��jc�7R���;��}lي9�ԝV��&���%uC4����#���C��2|��3�������<���:1�*�'�Gt�s�׺�<1m8��S����h:qMq��s]�Za^��kU�=�'a�j��(%�5���ONgJ����1�;� ���Cua>��p��׳�}u��y�;�e@�^UC@H���x*N�.����5�O��dd+N���)���W[��Q���/��˶�������)q�X�P�<=�`1v*�K"�8���S�罪{���Ş�>.����M��]Z�N��3ŕ��Hס@�i��aT��B�[�
/(�%	��ON�0��BF��c�r�u�d�	;�(	�F�����3L���8�D�p�hq�LК��o�G9�84B��A6��tq��<��0� n8�zp���s�f��ت���7^5X��봎�'Og׮aYp�3������K9>�Q,�`j"FR�~��	lR�<0s���l����"=�S�ݷ
@)F�E�K�ެ��[�&V��EwY��|kB�K�rf�KC�R��>��c����Օ�Fg�x%�����^i��.�AJ[�R�A���X�d��c�Ң�E����t��oM,�ΰ�*>���kW*�Ә.�4����Jy�@�O�ua�[ǚ�O#n������l9���Q�#�j��n�7Ҳ�H��+��Wo��3�-'Y��7�r��e����oE��(U�vb�N���^��$R��έ̪ZJ��"f��N��뇹��/DܛX�-Cu��m���1��r��V1%یm�I`kop�腘:v�,l��l�{�Vhc��O��'�w����W�7i(.�[�\��x�Qv�܄T��실�L0d��xh[�"��W]�g���ЙB�P�f�QW���no�C��7d��l�˛l	ي�e�d�cgS6J�@����#]�{Z���y��,�͎���E��Hk~["N�E�k�-J�;%�9I��J2�꽘�;�4�W2��ڍ��0��Z��~z�c��W��J��vG)';L<uVȣ�� <@���4�e�t��n�����Pg�l\�Nr��|�.�]`rz���AOpb\��q`����-Z��Nw���3�� �*4���zq4�h!Qh�����x�!=�W�Dv�[��R*gn�u�G���g["��=�5��N��swP��++�e�]>ۘpL�
��U+p�y1�I�;�i�R'��胂�9IcrmnT��f�g2p*�GjN�ǽYV�֗4�8�#�޸��򘫯���a��BS�a��pʻ�$��ĸ����/����������k;�mp�>��U��im�g�g�2D��>oh�b��l��֋)�kPZA�O_�w��� 5�<�l} I�c�>:h匉��n�z֩W�G�Ⱥ;��p�W��I[:/9���ΈW!�f�:	�a:��x�R[�K��t��ʁ�âqP�M��dǑ�rV��k3zR���qUbv�7�pX�uϪ}��9���۹d^��,wDP$�Τ��U��mu�����'�1�C�]��Vt�Mde�q\U��"r��uu�jg:Y�e!�~圉��L��wE���^ۗ�>l_~1�;k�ͮ��wu�V��Ȱ@n8��#A�a��gN+ZP���/$��2�,!��r�a���\1C1Er��{]')K��K����ٸ�z�13lNr�F3��[4�ajgK�e��mۖV�έ9��H��M[�u��!�i-75[���[D�w�<��[S�������P��5ȤX�Fe�pT�(�]�0���
K'\�(9���e���em��r\������WDSf���lܨ�������D�,��C���z��6Y��P�μ$��B5�X�[]`o4'z]ʚl��S�,Rk�J��&2/4�Gsr�7�m_�������뿯�R�LD[_�$�P]ۤ��L7"D�4�Q��31�awp��w.���4f��(H!�Ӻ��*%!1&\�Q��n�#3�e+a2�r�3���i�d�&L��#��F��r����Ȧ�	P���acC@����RQ�`��E�R0��� &K��$A5P%$Č��q��v�Hd�	��%ibE4��sAΜ�1�, J��0��L4����0C����!�J��C���%�$D�˻n��N�&IJY ��3�2H;�D�B��)�������v%.��pk�h̎�U�}��&��P�s�/��/]�0`�ڶ,t���P�l�X��GC:��h.[��C�՚�v�b��S���#Dz �F������#Š�o��\���޷�W�����������ţ�z���m����^")�!x�cڃ���a�{��{�DF�"-���c�����"ˉDğ����n�9�ѭA8%�,{�"@､�ݽN�_�.�%���� �ykt���{��<�}x��k���|���ߝ~���Z���_<�Z����x��{��7�������Š�V��V�0"Y�v�g'�`8^b����y�ٳ�}v/����)�_���#������o��������<�ߊ����W���oJ�+��oJ�<xѧ���ܷ��x��:�k��k���������3��P�+��h�Z/	p�D1�"��}�~y��|W�xߗ�Ͼ���_��t3K��ك��Z�Ɔ�vb�^�/\��W���_ϯ������sow�o�����7���KO��o��s���_˧��Lz�Bʏr�«��bh&��S��~>׾޾�߭����������[��O���h��Qe{D`�@c���׷�Z>~���b+��^7�Ͼm��o;�?��$Y����v/�j�_��`7�ً��P͙���Ax�W[�=31wv�������+���_/�6�_K�oǍ�ۗ���+⽿[x����.��f���l7�?��tϼ�]��F�_�>���u��1�7����j-��n�6~��-n�狕ӻ9'���f=�u���{^��/���o���/<�KA�������Z|���ץ������w�W���w�����y���nm��?~���[�~_<��o�?�o����iUWM�y]5��P�+f~�X���xѾ���齶���y���~��j7�z^ץz[�����W����~������Ѿ+��=ם}o���߮��o�ow�^W��o��x�[�z��U�A�=Aw9�*_}��>[�w}bf�
�޷of̙�Kz�{��]�^�>O�|m��~_>z�{U��_����om�ۚ�?�������o}x��������~^�W�����{�M�����+�_DX�Xb"G�6�UK����}�>��3����_���^j������]��V���/{��|ޛ���Ͻo�������_[w�_�ϾW�Z��o����o������^�zx�����<��zx����ok�N�<��Y98g�����b�Ik��v��LZ�,����L�9�F�g\���l>ʶF��3�ݩ���KA�	�y�B��zI��g�
v��:ݾ�e,Ь�K#�f�銍�:�$���1���n�H���f�樼����{q)�����v��t��6]�q�f��1OM}D}����a��W�������o}������zZ/v�P�/���#�������۝�n����5zo��^/�����~-�ߞv?�W�^������<_ͼJ�׿R��}�I6�Y�M�0x?�ۼG������U������6�����m��޿���[�����[|U{��h�-�����z �C�������Gi!���9��(�?����]���4�0vߊ�z�����x����y�ү���]�����x�]��x�m��k����KO;�o���}_��mʽ.��}���[����j�f�=�oH�M�ӥ�L�u�U��h��N�/�r��v^�,�����x���|^֍�W��^>+ſ�+��o^w����ܽy���m��_��yc}����;zZ7����-�vjv�<Ұ�ړQدsol���w[������;K�?��_��l�>�{[�\�m�����^��\�^����:�7���uz��x��*��׍ͻ��1�墼���ίm�ۼ�~]�C�B���p���_��_:Z�C��_���֍���������{Z+����ս�5�^6ｼ�ur�����>��W�{o�n����[~-��n_�{^��k�B��1L}�ƾ�T�#V>�����C��/�w�x;xc�wD�N���7��g3ܐ�݋������xok�;f�o	�q��+�x���?�W�ţ�����[񾷥x����W-�\�7�|�����^/W��zU���_�;z_���[�t�o1p��;��@���w����{��W�O��W���W��6�^�_�^����n{��5�^v߭�~�v�-����P�0����V�4��ػy��qnk��kǥx��������__�<�{v�=y݂��*���E���������x�_z����Ͻ�ww�^����wv��[�^-=����m�o�no����|^��߯����\��s��������Z-����G�N�!���C�{�y<;C�����c�DT��2,�f��?� o.�~��͹h���ίM�y����zo�Ƽ_�{����h��O:�W�Z/��_V��5�W�~{��^�ur������ivfN��o�oX����]���?�3�j#��o.��7fb�) ߥ[�U��*�� %ܓ���r�����\�L
M|��rXtٹ����^�_=E	�6��Y�+ �T]ܦ��%��U��z�-qT�;4-�6���,�s��5�EGr,�-e,�x��1bs�[O��z�:�7G�/z��3�{��ҹ�Ǟ�����˛�*������+�F�ە��/k�^����W�|^/�h�ε�������:�W���o���o�{o��^6�����k��[���߶�U����gVu|�teQ��іc�"$Gͪ��ާfd���1vOO�ol��Ҵ>v����ߞ���kO;�~|���~����~/So��w�^�����7��y�;{���٨�N����UR��/���I:����ǡ1=����/��^/�:��W���/�{Y�yt�z_���������H-�w�!�����_�A/ｯ_��U�wIO�w���'K3'hv/�[�����Zklb3��U���]�W���"c���/CQo��o]��m�y��\���y'��{�]�٭�z�����L2c��M�U�������ۼ��{��^���׋����y��-��W����~��^gU=����U�;�ewS�[�����^1��W,���^v�*�\ߍ{������}W?=�鷯��F�����^�6���[���^��nU��}��F�͹��>���������-�o���ٵ����h���wsX�E�^�������_�~�������7����^��W-��->u����<�?�{U�s~{��^�����~kߞ{W-�{�ѻNާf�g�l��y;S���o5v�u��ySeV���^gv,������}������ｷ���Ͼ~E���Ǎ{W��k���ݯǦ�o��oݼo�x�k����zZ����W�O��_����o���������⇼we��(s��]nhDszݘ�y���{�#���[��������o�5�}�������o׏Ͽ�_ͽ��\�o���E�~��{m����<nm��}/K���<ǼI��&��=���=�x���5�+��U�k������_������ms~��_�>�����oK����Z�+�^*�x7չ���^_~���ήX�^�ﾶ�U�s������o��[���P���=#�"D�!(�#[�J�S9y|'G5�4?�����[��F��{��=-����|k��TD{!"�ǫ�z����`��D|/�������x�}��^�����|��kO]o��}������^�_�֔��e�86O������.	2�3v�"��;���*1#�oaB6������ۣ�R�Z��.��DEJ����Ed��b�+���j�#��O/VHŃu�P�X#e�zq2	���D2J���d�O/f�w���:�>0sI����3������v��~�p�p�{�=��"$G� ���1���+�z�]y����^��n~{��o����s~��|�ޖ����~}���p�[�������Ãy���)����b�N����O�?���ؿ��<��r���wꬕ?��{����������|W������xޛ��o���ޗ��}����u���h�^���m�zޕ�z�����o�߷����W���o����_��-�Dg���R }TV���C�i���/Ԍ���_�.���C��� {���O��o���z��_^��6�^��^-�ί�^��箵��~���������h��|��k��W�k����z���j�g��0G�3Dx�??�>��=Ǭ�[�5��M��k�6;��]�����]�a`���7 ]��������}��r���xѣr��ž��~��]�E�/����[�}k�B7�c��"8D�x1���vo��eӏ���vd�/�c���7��͎��Շ�����}��Y��^��.�������5���o��<׵r��v��|���o�rߟ�^|��ޗ��-��|]=�<DW����G��(�wL�+���>OQ�?{�� G�}��Lz2�׾�$z$y��"(y�G�$z3VRvjv�;������e��&�C���,�F
�p׫��X6U�y�)�c�k�1��.5q��LuSW ��S�uN��s��Cucz����%A������j��I��o*YB ��3y�Bh͙*@c��ح3#�~�4�y�{�ou�PgL�ӎ�{4�7��SYl�&�o��WS>>�b��L��*-�
��vަ2g(���O%3o�¥������m�2�q'K�g�+��W����+��X��3k�Z.�M�:����n���IQ�+imѕ�,��G]wT��fz�6�=�aU��'SynX+�YN�Q���TARZ���>�}�8E�a�I�����r��z�:�π����s�Kx�Y�L���j].�A�1�V�W*�P<���grP��mM �]�Q�qt�����R1��}�=�t�bJ��7����	�~�n��e��Kh�44&�+|s��2��h�6��\!~&�W�l;�%L��R�m�w�����b(����7e3��U�空�r��]�u�:z�3�t>{3T7q}��JJ�T�5��a�ZH�y��
xE-u�F:j�a������]A���r@�T��%��'���|�n8�`�M�xz��1��&WM�����s4S�=�%��kz��X}L��b�&��ZǞ;������>H׎�W{�;����(���29�����8kMF'0��m��� �p�X
��E8���#�Y����+� y�ө"l�.&���5J�|�_�S"��L���9�3T+�Y&c�ٕ0�GS���瞶N�_+�~UW7m�م�u]Bԝ��k�2k��@;m�ٴ��Ŷ�M�����v��<_�;��B�_�0*�o,&�e��8�[T�##S��H�o+�u�*��D�Z�n]��E��wה�p�%�O-1���1�oC�V�c�]ߥ�=L�����el�"!oVi�ڊ�1W���C�
~㚨'.d� 1�%���.9�g���9����]R�#2)��Q�H�R�A�n,��S�l��P�wj�����ս۳�\Q�)�.`aָ�L���C\�װ�x�c�� ��yW�5�oH��Q�{{�+�R7�{�y�5sɌӛ�����.'v��/��5kIw��V�g#�o|���WJ�˙ q�]�q�&��f㻜s�་Q�ω�-.���SD�ķa���p�v
����n�/P��O2�z�������m���rp]�$ע5���gd�^�ƽ�A��w���L��@���˴�`�+e����<i�B ��V;���܏�>�� @��s��G��ʘ/{����=^\'�2��I;0�
q^�|�s���R��g����I�2���H�;1�Z���)��"�%�3v����#������O#�n����s�Shm�r�W�5(a� S��L��Z�C�E'ά	�e^��ɞ5Y�'���v��Z4�W�Q���#��P�8ҀǉJ�z�y�M�O2��[P�(�������z�t��.tCg!�Vm��^X(�H���]Ʋ�����k�j�WGF'����*���qC��>���U��Z>i��Y����r�_H�Ŧa!�+��QE^��M�F�t�-�Vq�(h=�!u��搾���"��nEۗ:л�������j!�+)tw*oq\�����Q>ku����r � s:"�T��-��<Le5���71��ͲZ`(Sh�WX�p{�	�����t}E*��XųH��i���Zn5:��5&*N̖�F=�����[x�����n��Y��[^V��02Z�u���f�1�h��GBs�=ߠ�=����[�$w8��.��"F%��@	w��o��_ڼLuCt��OΗ�a�
��/�G��i[�����ǩ�fj	F���T�^7A��T�,.��T�M!W����6'��ܩ����6/x�6rT��c�&dGpɄ08�Rѿfڶ2�xM����p���S���ͥp5��+�{��,e`Q�d��m���ZQ=���Ԫ&;�y�SI�Nэg�U��u�lEY�� ף�C�맹k���aҜL����ϝDʣ��]Ӥ���Es��\�vN���=l�	�q�:�Y�#j�8Ӏ��#�+�҅�T�uHEtiuaF������<Y|�
���7��H�d�=;�|�G�p�9�����"d:�C#b��+Ћ���+s�,eQU����G�݁�i�����XЌ?�u=ğf.�(f\�q���Yn1��nt3Ϧ�0}���-%z�G;�8�� �f�d���I���/Cs0�V�O5��	��]j�;�;+z���^N[���*MKz⍎��=舄�^w'w��u���C/�h����a�J։t-]T<I��_Q��k���=~T@��zQU�4=�L��:8dZ>qҩ��C1����=ꑪg�A�^S����`�1���~����8Cg�Ucx�Rj�n��l��;Ny�"6��~sH�)�D�l�:��d��j��1���;귄]��
Fx���yoW�T�Nih�b�nbsr�-�⃜��K�2.�x�UjGK��$O�'�M�r�cr����k����e�����]��v#/u�@ʩi9︿�s�I�
�v�U=FY��t95W+�U�� �����D<�`�����̭�&O�2x��5?E�7DR�x�`��l�:]�Ǫ�5Ͻ/��Yz�r`�隄!�ݾ��*0���4��r�_���=,���Mx���[�3��ڧ�kH;�����Z+�.����NOfqt��Y�c�sEl�Y�#���%�`	RU5z�����ß:���2��<r;�3q�n�jf4��z���V��<�L7w]��[J�
��� Y4�z7Ӿ\�_>Z��e�bq��z�8��˭���\�$�R��g'����������`¤"��ݕb沥<��-v�����r�ԭ
�5*bu-R'�*;��Y��b;��zv��E�y3�M�]?��ذ_|�~��G�>�]�X�l`(��(�ʃ9��W�}gG����U<�J�K���3���s��d�U��(��ʑ��s�u�+��"7\.�{O�v�t���.�g>��9���g��:����
�\��yHs�O���}�p]V�kKg��:7�G.�ҾY��<��loM�٨������j�*��S�����h��m}u�Ո��'	���2@3FUо�u}ɬ'���RXc`+]T.������\Cۆ�\KT�d�h�M:�����#n��z\���������!\��(���	�S���2��*�� V���o�}Y-�=����&	�& t�3p6R>��U��Su�QXპ:\W��:z���e�ڻJ۴�gh�>�:!P�<z �`��~��KB�/cw��M��f;:ڧ2�J�К�Ѯ9Wq/]D�x���*C���IO8�ӊ���ʧ"<R�q(��s{�ޫ@!2b��t��f,2kͺ�.!㸚0Y��|��;$LJ�tL7x��t�9ÑN`��c�{�x����fl������B����S�|�@�͑�i]wn���8w&��w�K}Z�\�2�/(��;�2�ڳݦ͗��9\��D�H��:�j^��z�#ۼ1�s�D;3���Sz��#�!&*�s����"=�5��"�o���;�ѨˎU���p/� ��P����t�}0L�mL�z0@B]�j\-���8��Z*�a#�n7������کjy�&�7@s�f�W�N")Py=5�9�U%Hҭ;~*ଠƉ�o�Ǽ��]+��y�bw|c=�|ɯE�P��ʬS�µ��]wj���E��p�0H���c�xpTW*�b�7egh�b�S����F����)b��T8��:8�?Cu�y��'v�&M7���d5��u�48�7�ր�7�q7�u8��$�Pp�r�^�5sɌӾ����r�.'uѺ�Q�/�����f�����+��8�N$� L,jȿGT�D�"�N�.�Ob�}�j4��0e�]�d�ed��S�����4rj)��S7�Ѹٗ\�&���_o�ߘ�/�f�:��ٹ<4�$qVΏF8���V?A��&�N	���L���R	�����K���Xo��eKu�gY��j�oE�mUF>�:(�ZH;�@���<\�x�)�����p�q���*h����m��&U�K�����!����!������=]E�E��'=�ٙ6�	9�gk��/��qM�0/�"K�Z�GS+A�[-jR��D��.�Q�|v����u���u��:�3����kh`��UG}�:�vi�b͏�)U�ػu�>��EJć-�`Zj_o!�NC�
N�㱎���N��qЕ	c���9rY���V2��.F�;y���KOo��h̳�͐�7�Dr�,H#���N|�nU��1Ӭ�	��r]�N(��j�-��e�s,��';[�ъ]¯����ȓ�����y$p�zDK4Wf�8����p�zdUݼ��ޤF<�1U��&�}B`��{x��<��:��nV��M��n��
�Lɲ��պ�JJ]c
�7��8Z��
�X�K�;1:�&6��{�%�
����Ʈ�6z��ʎ�}K�[�=s';��f;�
�֩�X1d�OAS��h�c؝�,Ьq՞Z���Бl��	,i��/�#K�U�㧝q���q���f�a��V���fn��З�P1%r�=p���Z��u�B���0:�{�d8Tt�)[j�!��K^IG8Z$���������3j��w8N�K�z�=�����/�w_R1���jC
�Ջ��N�o'ƥ2_'J��Ӣ���-�݀�pnM�s�:=%X��ԙ��AB��u�9��f�V�w��(�h4�w�v��:�b���n����`�4j�#6t�+�& ֳ-�����Κ���umsc O�븓�`=�-K��K����b��ƻ�jM�F�)>���Ȩ�
��<(29d�
��&�:�VIsuoP'rk�o$��\�23�����}\w��_8:+��+��ZS�ZבΚOFkMΚ�U�]6!q5K�"�����Kt��Z�\�"b�ɺ�`��=�N϶����D�H�YJ݉��ͣ��F'op[�H򾻸*I�v��y�/��R	BG]
9sel�-�U�?��s,�ν�Z��9k�d��]���RY(��SU�{��jʼ�*�����e#�BWc�_N���ˈU(�.(:vd1S��p��)0ox� �%����+C90��t/7*ƽ�-��� �@W6H������,��N��q��ۨ�p�>r�7���w��([�:�z�]�Z& FtG!���]F�
Sok4�-�u�q��݁�0ZR�<�y�\�cq����Ȩ^,����&vc�z�F�Zm��w+�7�*�;���pt�w�׵�����r�+-�K�i��Z�q���­��47��1�Ǝ���}jk�K:Z5�dw�ˍ����.��5�jcđ�jX��Kd����薮��K���rd`�%>o���M�B0���9�4����ݴ��#i�h�Qk����\x�찬oZ��g ������˖n�������	o*Y]L�n9z�q�'Q�~w�׿�������������%!�S)r�]st$�H� (IA�I .nf�A��RA1� LB���u�3��%��u�)��EE��wX�0�D�;�P��bP��n�q���D��4�y�����v��u���Ei�졮���ʀ��3J!";�s��E��Ǟv��0b2���wp�s�&4�&3W:�w�x����d��p�Ɉs��J�r�S��K��r�	"�S��#�e�.����1�]��0FH�e��:�D�:��W:P0b$de@�M".� d���"x��	��Rd�)%�\D�!�3M ҌP)I%�0 %,�ה)��I��A�If��,��y�k�fd@�@R�(
�&�w��k�FV�%�z��]�>qXYR^��̹�z	6,�c�`�	wGu6yg9�;nl�G��+V���Q`4�A��G�"�Y��&������:]zaY��A��f�*BC;1�o�]AwM�	I�]v(�UT��C�
(p��C^�Gߕ@p�|��h�c��L�' ��V+�Ad^��2�ꖱ�����z��-wq)�p�������ڨ�y�	�$y8@iP��ʗ�H�*]�x��4|�����C!��O��-�^��$r���9X�n���	&272�� {��7�-���)�o��̠�w<w�Y5�^�}e�!�\�%�6M��T��t�[�z�۫R,t�!��g�f5_��
�0Ċ�h���+ju!�Ƥ�D4��+�/���d�ݻ(yU9�S�W/aD�f��*�F;�
�g��(@��o�L�gr���荩���N��2�F�5/Wyx\����c@���c����9��|ow\�`��Wx�s�T�FT����b-9�7Q`騆�(*�Պ_C�����*������rGQ���d����3y���<&��.7����{�.�u���|kV���)<��zv�ƻ���n���E�}Z����=���(�/yC[�j�J��}��^��t�[��jeK��7.��I,a��CrX=�z�AmGenn��)�dޚi>�*�v���mN.�͖��b�cg�0l-2c{����DDxM����w�D�������$�'���y
��,��;�G�����w�n���m��dY�/#�p��V=U%�a8��]�0?����P	@چ"���X9N�=��5گLYą/W����2���O}M�f���Qʡ^�Q�7>уj���!��EՅ�]x@�;��/z�,�m�&�J��^�.���Ed4�5������2g����2${�Ec�����^T�J�W�=�&ˇ�B��w��7::�\�<%����tL������� �'㗈����t^�T9T��!����=���lhm�7�0Y1� �Us��� W�ދ�Z�ًC�E�b��"�W~2�q���9�nH����e��f͝�v%�=�Y��K�����!���B��5w��\2�c�r�lÂsKG<�c��oVD��9�kJc儋�Y��<I����j ��Ȋ�P��,5x{)����3B�]�W��n$؞�:X"��lסJ����r;a*���t��"ݮ�����U^�`�Yq���MWJ�{R�r��\�ޤ��V�G�ٝ�8�km^X�}\�q�G��dOxl6�\;v�z����x�qm6B�j	���_p:�Zs��(��Av\��S[{w�i��[��W�D��,���Ս?J��u�n�tՍ������Kmf�:�A�4d�~mS%�r��DX	���>쬫�8\�u�����'��3[7��B��B*!s�c!�WG 1М�4�G*��<>,��姢"V@�)i�W��>Ь�`�vU��;�R:a�,V*��é���4G��C���*U��a󻴤��}x~"�����mpˮ���Ȏ�L�u��&��4⹕��஭����n��y>�mc]j���8)���5�P��\G�4x�*j��Z�a̺� �e�i8�k2rWvj������{Ɍپ{Ɲc��@6���^��'j���5C6-��&�}�����fݓm��{������'˗��,ci5����2���*a�s�������k��T'�TnH���;����u^n	�J�ʦ�C�J*��O\��S=��Oپ�v�?�Uf�ƠG@L��w���i�-��f.Z�_b~I�PN�8ȷ϶���yGz$����u>5�*X�,'���g��8��E�h���_ ����È� ���Y(�5���S5;r�k��}c�{����̠�=% #����A&_[��[�}�C=�g��?�=�;U{ȼ�ݪ��b���F���b-�R��i�O�#�&�JR���t�^���K�(>�P��e�Tws�:?{ޏDDC�q{ɺ�H�#��8 p�%�0:y��)Z��e)�p[<0s�K��Wv�W7<�y���x����p�a��� H�k��4�r��S�)k�:���QszƉyv���l��9�ӣ']��=w�>�`#1D�N���]F�8=0���br-�r����1Ewb��{�V���b�&��Z�wP`�^���#ݵ�x���I�w�^�����7Eju��j2�C%�<A� p�F,	UJL�t�}Uyj/(ڕ�\��g���b���|&�)��u������J��Ԋ�S̙6��9癪�o\��������K�@��0���
���/��?�L^XT.��I:�0�ϙ4o�Vl	���I�mk/h��q����"�Z��.���C[�	��|<��0xyLf�]�r���}����3wT8��uᪧ�>q\/������2殽���y'e���㖖�]��xo��fl�8��u������9��YWR.��~3Aj�`��]��;-p:*r	$\ά�+�D0~ǵc�G2��*\Ė�8t�Ql�T�vbˌN��R͵�z�A2ﱸ�^�����5�U�S�R����ts��=eVgG��*��Y4cee&����Iuĩ�&���6�G@C�&v����8�ԢsA�f�t&��'1��������w���	9���C Lv5d_T�D�"�N�ws�����y�Hx�.��P���*2��]B��g}�Ѹ��p�,2j9�e�:����c�wJ��e^#�yni��c������H�#�3��/�6+�b��+�.�7����l��uԆ薳*f��7�[eo���ª�tQ�t�u�� |+����9s��]t�Y�~Y�V[�t�PA�ɾ�A��[逎�j��A�f"Dp��=�+��!"Ϊ�ߺ�[�U�i��5��S'*��`��*x`�o)�����892eJ�a��yٺ�/�2b%�Z.�
�7������	�G5�u��\M�w,���[�J�=�#j!�!(��#�}���m�u����]�������ڠ�3�s9Q1�g�{$=Gօ{ǩ�Vp۾�X)�Y\��L�)��v���Z����v�����e�����2�OMu�6��b��d���͚���|���q�� �m)�A0ݍ�bFG���zV�Nd5�/�I�漧���}Y�_cnD/��*hY��{oX<�'�<&:v[�WC��WB����X�ow�:Ro|z��ւn���lWd�N�z�2�-�Z��oY1cT�ӌn��ر=[bkf��7Eȣ����"�����N���G@�(��ؗ]�k&V��J�_}vB��e����foVE��i�&H� �ץ��[�4�����x��/��>�N�GXr��G*��^Ɨ
�r�\m\I^��j�?@l�3^nX׹�Tkʐj6Y=av�	�>�D��7F����/u�x��-H����k�S��fyD:�J�޺A}�������X��8]{\�̽}I���;/V{;Yw\+�3<er�l`!�-O����;��W0E�a��7��ܥ=�F5�%ixygf#�S<�G#fb;�|�i2��Q�g�!�~�AD��m헩m�n������?@������P�bS��bz<���4�N���1�2���(Up�M��ޗY��^��+���j����Q�^��p����𦷘��<��Ln��t}�HU��������s�Mx�W�')�����aYt����}�6T|/�g��,A��ϱ�g�,�C�/sc�[��a��Bۆ��M���끶Y�f`?S��~}֊�:-]�'"��s�3zw"��
7V�"���C1����ީj�ʁ�z�Iu�b5�3мE���F�K�	mudJ�&q��'*l�Ռ���J�+[Pܬ��������S	�k�x�VF�v���n*ci\6WqNue]��^�x�� �Sky5���h���ɓ'1�6�adX�=�f<�������*LMh�.��u�ވ��=�/��O)wX ��K0ƈ���W���Ȥ���g��a���"1��=�xN�ؑq4��{2� qY.��JU�Ce2�`C8�Bޮ�T�斋�u�O3ɟ�;|����U���K9.({�<]s_ui"���q\��
Xwx{�	��(�ܴ��,�kz�����\�� S%w�R�Γ�W#�MOhS:�ty���M�Ǣ�75ҫM�Pv�Cڑ��=G�)d��9�@g��"'�Q; ��ʌܜ���r�qE��&��v�Na��ۄ"�=�2Uto 0���k�LW��i�8�v��C2,�К��_ڏ��G�$v�[fB����Wk��xg��@z���C�������+wۻ�/`�wiOQ�+�6�%�1}Ε�2⺗Ǹ�oiW�)�xb�q\ʷ�tSl��[|汻JAީ7�uF#\i�ʬ<MA\=L�خ#�<K�5p�d0)8�V�uӗ���kt*nL��(�ȯOf���\5�-�v����fp�J�{�O�DM�̃(Ͱ���k�=��K)l�}���5ғ��-c��0�
�o^�&I[K�N[��u0��Va�,:). V�&��%���RL\a{j����{�[؍l���ޣΖ� ][Q�h�9-!�d:��k��b���?UW�W���oR��b���\d*�^O#�DR�r3�l:Me��i�2m�E��E���Է1��5YM(�x"�� ��<�ػmP��E��z��¥כ��b���m�2�$�W݉d��cN��W#x�7^"7�@Рj��\�+O�yp��[��g���A�i��E�bսv<��^��'�% _P�����^���HК�ԭ���!�� h�5>�h�u�6۝9Y%ThpM�v��GA��(	<�����1Uc9�n�j �x`gKh*]�gH�(�����:e��}���P*J5�@�!i#N�5iP��1҇��Qu��["������
�_�͖5��%㨝/�Y�������:Ls�n2�t8��u�(�>���%����u˪ ��I�C �H��3-����Q1��|�du��C���2?72[�|��}sذ�d�^r�1^֍F\r�d��h:`�X��R�gv�5���Oz�y����\h��N�`�0��;�+��}~�6�$Z<ɓЛ�9ҋ�67�/���Wd����c�c�)m�c�UgUѸ`��&�Q}و�M�w��q�������e��Z��{cS����f�y�{d�D�ҽq�̷F�ȺL4��c�4X��v���j�{sq�<*r%�]7�V�G�N�1��$n��/5�Z�;���"+c����xgf'�n^a"��I��8�uGǅ�uML?�~+Uv���v����g�֭�ǕP3�)��U̟i.O@;q�ٿqzg���.�1�Q��W*�b�e7f-�� \m�>��"&A%����t8���^Q��X�������:7���d5�k�z�[N���xv�G��̨�P:�_ /\�����y�����+}��.�.'1Ѻ�e="g��`��W���ew��r��Bf"8 �gu�u��o�0WE{RLb���1��՚})!]���)R���a<7e�U\�;]1��p��&��e������/�f�:���ڸ��LK����Dy�=6ݟOQ&���y��u�M/EV�0M<�?�����]���?cNJ��)sY��m������������FOȃ���!S=\�_en"����Ƕ�����ӊ��R�y����9���6�l��*�1��p
���Ϊ��P^��w(�����RQ^]��ë����<��g�Iö�85
�B�%���P�[ꘆ�Y���Ֆ|�
�\�-c4��Y�^l�!�Zm�\�]MW�ܥxˇx�y��z���(m���:����^�V37u�z��+<���ʾ�X���WXF��=˵s�1��K+\���5 ��Z�5�#'7y�1��R��e๊��������bn�8ۭԉ/N��
�¢1>���q�;���J�c�T��)��yL�����p�We�&�º�4 �?<`�V�p6_��>�5�+ԓ��g6W��Vp۾y�9�v-�n�J��� �+�T"�e@Ŋϭ�e�;�;��&1��'���_�й�}Ջ[�eLY�L� ]o��40�k|��UW�LH��i�ޕ��:��BOznL.�ir;������$̘kuY�p��k�F��֯aD�x����@��?�GXr���ǋ�*�1N��I�SR�ު��&C��nX�6=��A�OT��E�~��5N�'-zd�y�/K���/�wSa�,[ULE��̬u��Xw�b�q���'��f��t�|��	��P�%�$ň��Δ��6ձ�xM5^\n5]Aۏ�s�ݺ���w�8�����ᒈ�e�0�'̪>�<�EZn*g�(�f"c����
��,���'�I��'���߯�H��ɚ��O#�.�ᎂ_F����!谞uu�J���,�o��,pr��!D,c�V�z(w�x�7��:�c[�7�e.B�
�t*�y��5m��U�従��d�S9n��2�EY%��2Z��ٹCaڐ����ro�ە#C��LA����ggv�qv��*9;�ٖC��;��ȕ�}\��	�r�^��'خ�5DV���r*89e(S!NT�Qۥï[�ó����p�r;:�+�#�s����f��qIVb�")���4ʂ��$E2��Ī�P��r���[���s��Z�U�&bF�>�O�I�Z�B�q��GYV���:�E@�N�EMj�����o�h�DJ���P�;gا
������8L��h�:�8V����)Pc9�Ϋ�X�=���1�F���������K���K�y���t�Ԯ�w��:lhn�		Nb乜��s���
�ц4rk2��$�8�v�@Ņ�q9�	��x���ԛ*eȺ��]���p@���yt$�)+J���
���]v�gm�VI]y\�)�t+�]i��WA7�k;�R���	ZB�3���`�X�,|�i\��xfJ��mzYH:�QhVEK��&��2	�QL�󬀐���30t�\am�2���:Nӵf³�,���`}�|(3�����X��]����:�ի��r���.G-����1�T"�{���ao�����q̮
%��9+��i�Pݖ�-��^�R��(�QV݁/#Y��9[�Q���:%���Dw`/kCF�$3l�Oy�<VF0eG�-��$k�-o$�g����Y�Z�suU���L�H�Ńr0�u .u1pZ��(�2Iº
k#
ƸVbw����Bt�t��ri�mY�����o�wg�?�N�b
��������
�
�igq�g5q�,╓Gr�`���(E�cY<�-��wW�WN��ܲ3B���rWf�3�[�eѕ����L
'P���f@UW6����Z�g4��+���sq('�1��Ws*˓�]k�
�Ӿ�E��r�ia!k�����-�6��cYk#rQ�svWYej+I����/���ORg�c�V�Z8cY]���4��]�MGـ����7@�T�و�"U:	�Gz�'hNn;=Å�@�i�Z9l��(�+%�\�r�������N����5�N薃sd���4bB�7'h'�a��I�I5�k�gn�ѩ}/�a��[a�����
���d􍳱Ju���E�k($��q�{����v��
;PQ��gf�Yx����
sP����HD��':�KJ�W��������H����,C-�_%�ܺ1��3%�L���fٲ�43E|^�O�6�^k�T�v;��sŔ�T�T�᪱H�'�CV)w�+9М&^�T��-Qg�Lg( �RVl;v���wY���9�l�j8�����ëCaW�
V;a��NS6�}a�-櫓�X��{Swj��a:Y+��v �6(����bc��J4�7��R4��M�)�$6�u� �Ę
s��ݐTe�k�A&F����\�P�	B/��&ȠM0�rh�2� ���03L��PW;�0^uѢP<�Ja$��3��u�	��D��K�r�H�I1&���!��Fai�JW��@&LI$�ta��E5%$C2�Q%0jMbQ) �+��!b��Ƃ2�FM�.WwL�& Cnr]��h�0jD��웗B0^u�X�ƒܹ��3��dS&r�wnM!l���D$�HY�y�-H^w-ݣ��B�Q��n�-0��$Da(�
k�t�T 
 �h�BN׵���T�ۚ�4"S\8�3���N��zi1��IԤvB�
�����+f�v�̾b0�%���K�_}_W�V{׹;ް������t������1��Ӱ!��ep�@�<-��Mo1ǻ����#z֎��f����j��*�����g���v��KK��Y�+UQ��QQ��u�W�Sɠ�m��}}�ݕsۢ9��e���7~zo�s������fb♛��a�K���b�]���0��*�a��c3��hÿV�������C1���zo�z�m�W�S*x%e�Nz����^���I�V��р ���БW�Ucx�Rj�Ag��0�i�y[&)X�<���c��ZH���8g�C��8�rEĥ^e2�`C8�ޮ���f:d
��[)(&�ԝ�ňpۨ�s,��S%'� l�2y����W���=٤�^�y�[�=N7��1�-�,�"�)��g�R����	T��S:GG��J�c�K����ڢ��b�s��W!��=G�)d��9��PDON�2�#��"gb��aj�ޢ��>�u��-�"�����7��L�0��r�Xp�,Qʕӧ���2Cu��z��SΦ�o��8RƘ��a����^�B୳kM�Pȵ�̤��zWi�B�Ӂm@��&�f�[�2���t5^y.�O;�P�j0�8�����Z�n�8��jY�{������.�2q�qZw��$٬1�,�W��W�UW�c�擮1rM}��96�*�7[/�Gj���*��ow��~���\(}*#SR>{�v�v�vH��!s���jYtk Fׄ�?v�~t��L9"����&���-n_q�KS��vd��p��x�a�H^&�5��>W�Y��{��,%��i$��I[���գ��=�¥_�<v{Ɍپ{ƞ8���@H��u�¼��y�=�7��������H�h��i��;�t�܈\��_{�����|Os�1�V�w�[rcb������}f�ȉe	f�����[1}ȇ|�r��·�h�V���z�r�Z���HX�$�rm�2��C�4(Z��gONi��6aD�Lp�0�8���u2�u�uF��B�6Mh�I��(u�4�ׅ�8�qp4&�R��=�C/��u5wg�����]m�h��"�5�p������ c	@L�fll�}x����7^=n��t�ed�v��N��2L�;�WqmI����)�!
$�o���Pd��@�=�'x8,�>D*�v�*
w�z��(��v�ő��<G֐�ħd���KI���n�%��e��r�{��������Ng���B�Sw�Y�\%dV�;0��3�:[�o��]��-
��Vt���v���c���2���0NI�����W�UW����[�:jpGЖ�1SW�e�nwIp��[;T/��hCl�QD�)M��p6�������]����]AP�WM�����T�-�&.����h��M{�1�H�r����c�Vɿv�T�{eQȮ��^G+����r�d�n��� p�b��$9��z��C�FK���|��؊��x��'���XSU<v��zW���i��+֧�2OK�6�w�Ӡ}LZ�l��{ƴ�t�W�z)P�c����W;��u�Wk���=M�7v.�,����N���;Xa�>D�[� ��w�o��8x@ao	�
�><3�Mz+�s ��ڿv9��m�;"a�m���C�,�^^�x,L۽(B{���`���m�έ���j�����:\g[ U�b�g��y����i��biu����^����3�p���>>��ҵX$��}VD ]>�HvjB_�
�jI�V�[�Z3f��m�VqG=�s�W.�z��xa;d��T��LCF�e�W �ɯs���~c�ދ�a8���VVwF]�5�b�4v.�g���)aa�5,hD��56E�	+�u�c(��6�wZx�W�mVr烔W�pï)V��`:E��8vɯ:^*/��7����-�R�[��@N�Sx�m�}׉C��7m3��O��8]{���y�j�/5��2%6C[��(ຸ�4��΂Z:�^���`�����9`�cnjL�33�e���� ���yw��_��^�U�0�|�:��,B=\�_er��|�"z�QYS5˭^�t�3o��8Ϫ�1Œx�=ā�y��oy�HU�2�JnQV�a�Y�)L���Dc�U��q�R�"�}]�u�������qkzo��� 3���&-B�p����mӸ�e�>:���T=�#i�!-�ttw>���0�V��ۗ����� j�1��bB�ϒ�3���>��!�m۸Sq����o���3��H�r���X(��D�l����4w�j.e�;�;�,���{�(|���C4��h��}ص9Q3rz$FT���)M�D�7t��g��^3ᰴk~N�z�H�v�wy��"rF�2a���6��k�F��K�GOT@���tb�uF�;�4�*F;y1�*uK�t+�xI�f��]w�-'wB�d9��r�%�,?���.�x�Xk�O =��Iy�k�g��n�J���![�ۃ��$�c��N�M5��5K��duڻ���謤�b�mt,k}M�}:���ZV�,m�<��>�!�f�9�3�,�.j��N+�;%`�l��F�f\�e����D81��-p�����G��v�"֚�9��K��~��!�{���xk�Sx�ec��t�s*:��@��T%�����iot۽0	8� �4�9�����.��*So�f-^T.ϡ/ܾ�9��ùԉ'��k��|������膺�hE���ΩD������t���Ʈ�)�J�/��0�9�Pq[3N4���η���`�M�%A/�K��k��YZ�ۜ�J� 	y���ޓ؊�M1^�S��Oϼf5f�'z�h�t����B�҅���]�rc���z����!�}�S>��
-ä"۔�e:��A����� F��Ď|�N��^���L}pڙ�{�ic2$y�Ou؎�e�ў�e���w����A��,��x���$
<�'�o�4��7�;�Gţ�~T{������j#�Ͻ���{G� מj��]d��ER�^� �7P��jKB�b(hH��V7�E&�&�e��~.a��Fa�D��X�q&�7�#H�p��p摔H"���ʿarg�(+�0WP����5vE^��Uۀ-.�M�.�R�YR�a(��*\��?G�aY��v7�$��3-��y��g���]�O��=�]�|���Ǖ�tQ����F���@Wk�N	R�f��J,5|��hNr��\L���oq��哗x:pяfW*L.�i_�'��������2loQ�2v����<�y���6�'m�2��\����T��L]9μ6����	�54���ND�5�o���A�Ֆpl�lע|�TMGRv��s�3{�̷�1�n��wހ�X5Ǵ�?j��Rcd��J�/�<�*�U�tE/��tc�bu�6���^w���{S�Xp���^��2�]p��p�����6���`;��K�#�aq���S�\sH-��2o[~cG��դ�~h����ָ����It�j���=��� 99W$�pom*r�6���$zsZC�i�\o��}�����+���3��$�����a#��l	O3�8�2f����CT���&Z���'/��Vw�ye��N���ҡ=S5Ԯ�ld�}m�n��7��fQW0!.��-�N��^�ҰFjrr7�8��i��ؿKOv���<�=)}��Yu�D�{�����yt����rQ�v������nDSO�s�[Z�N]�r��M���� V<�my������ �K�|�8���Ί|�Mٷ�pA
m��u���+�=,"����r���!��Rb��ي�g�u��v�[��j�\�zȒ�O��2[WEwE��Ƚ�ܣ9:3T����乔�W�u���y���Nۢ�២+@S����}Q:�%�Wio/7���c�3�[�N&�Q;��Vۃx�C�l>U%'q�2Y�RyK�N�� ����`��q�=���ͥB�Oy��^�f�jJ��U�훩��z�Wv��L�L֖V�\7�s�y���PS��񆖁i��V����7x��ͥU��:�k�9i_�<׸��x�l9fQ
c��������c$y=ӭE��9�MM��C�T-ᔓJ����)��^v�ν[{K;9�H��V��:2Ͱ{�h0{Tק�mo&���r�[|�n5մ�:�j	#�U�|��������L�>�o�^}W����������m}��U�k�7'd�]��D\rۃ��ﯢ�mRQL�B)��O9�q�q%c����f��P�UF�7Z�*ь�/f	�(�8�[u��9���Ē���$w^=�u]�TGLa�Fm�Sb��Q��Ϫ\/��͙��yy���~U�; �i�+�za��h��E�p��LR�N[���Zu�qC�t�Ϥ���t����-�OV\��������,6'So��>.���v¯���E}��l�2PϹ5Q{X��KیN5�r7�U*�u�C2���!c�Jo-oG6�Uѵ�^�Ix2�LV4���q�k��lkޯeY��t���M�.���L��N�nr�Jc��TO�� us��"wݼ|׌�;��nfL�57�S�;*�Ş��^�
�1�Q�7��ǧ,�nRkN��3��V��sՇ���
�/��>yV�	���w��$#)[���.�T���}r��z�m����hzq{.}^��D�^}����~ښ�?K�?|��p��Ĺc�mT
��*Ը�R�ĕ�R�Z=W�!Vc��:�������Z����=��ʡ�|�;V�ܹ����&J��f����g�Ψ��ל��ky���;8������Ӊ"є\i0�N��"�Q��Nq1�y���^�u�V�����
�\.����+T-�e�]�t�������ni� ����k�`�d1O!>�+mgWY�����kUc�)��vVV��K�L��+DM��Mj�S�Qʃ�*�}i��;��=|�N:`�x�۶{F\r�ް�y�1hog�`���Ӊ�yq�?���z!j��&*�:;�G��D.�)P@O;�q��A�w�ԉз�fs����n2\-��8ôr%R�lwn`��ϯcXh��u�_K�I�Eo7�zi��N��5�օFF�"b9�[�˵[\R���ls�7ˋ���%�bI��p�����<�vF��o:'k��Ҭ�g��^�z{>�ݖ��o�>՜�/;�U�흦�f����v%�Wu�v�e`Ch��o�ی�i�J����^��'�����ֻ���)�QXO0�q�q�B�n��������'�~¢{u7�6+h�b����͛�m�5s+��/l��͓�V;8�xf:=j���9ʈ����N���x�5)QWs5�v�M6.Z{q+�n�Y�v��A�:o��ʹ��a�)K3����M��p�\6�\K���}�g�)�6k=��ڞ7DSdw���EC�$�ջ6�{��#��@��Ĉ(��=i<P����z���w���H�&��|^�f�	F\�wRשpE\�L̣��Z�ziL9��:�ZH���*�Z)�;#ϔ�o����Y����a�P<����2f��&��Ys�_}�W�ٻ�w��RPo�;�X��#���˪�W�\=i��V�U��6�����#��e��;��rR뮠�R�^)<��m�v'A�	p��{k�:�!Ӊ���#��(��5%x�8�Ǽ��dl�ָ�v���c�A�js\s���(�"[���dC>
zwP��\�T��̨N����6��U	�};���k!��P�:�9�1!*�>��U���2oi�lbǘ�:��՜�6������w�	��T��Ghi	��3zr)Z�U*�妕#����=��������u	����q����tD Rw�E͓s|O^.�-{�`ax�B;��#���'���5=m������c��:뭊:�v��U�$Rݲ��"_T�Ë}���w�$�,NW�	;�v����&Lip����7�\��F��-�@�F��[�$��Wޚ���WYN�Z�����f�j<G���W,vT������)>�o6��j��oR���ʰ�a�jaŹ)���+���5�d�	�[-�e�\�M��ru曮t�s�޴�r�M���sC�m7t�2eȞ�\�늵�Ő,��l@��;�fSW9�K�[ts�ɕ6Y����'/��uw,�˩}�v���b�}VtE���zk��Z�4A��̗L#J�G���&)�rA[Ee�+oo��vY�ra=�^������چ�R�^��j�Z�S�PIǔ���u��&�;1�t�qa�ʋqܢ1/D�u��n�v�4��ϰG���I!w	2�U1�6�Υ�h����;q�����r�*]��$5��4<t��՜�wbT�����W�t ��O�����U6�AM�'���G��ʹTʝk�
\������Hl+���1�5�t�^P���N�����-JWc����vr�X�7ݠ'�u[���ٴ}�,��.Ux���}Y�SN�s*t��kMMe0�&�r��>Mb�0e���hCH9�
�W����X2ŝ�	J��8��MaP�m�I���7)��qf�yNk얦��	:�󂢯�ƬG�[��n���bX׷,<���k)�]E[R�Ef����@�����$k���\�0o5�������I��V��f�q�ɮY�ֲ(`�q�f�ܱ]�%7f:���o
4�;���ѕ�2���]F.����*��m��v��9S����ĥi�'&��u��!IWݗ�
V�a<�f8�������v;[V�X�P8rjZ9�}cBg'{�B�F哜ѬW�w�؞��W�k7,LYOd��x���#�ܬ��gR�-�x�lv�������s���Hۡv�g�y�`h��,gL/R��|(C{n�+��3��Jo�c�W8����_rkI�5@N�j���YSWf�><��*�a�H�ya��ǒ���đușj����(,��$�)������f5C���:�t�s>3^m�`5��'��o^�'�f�jh4%��k���u^ŹG_99N���T�ݠK���o����yS�����{å+j�XA�Ȯ����!���
=������[��Jv
"2���D�ԞjY�F�w'.�x]3);֕�
��O�A|���ov	|�]�KD�Wխ�ç�.�WǧL�Y�eJڳ$��Hmt�"��{��Ǻ�՞A ]#\*�v��
ڣZ���N��|�Ɛ�θ���K��Պޙ�x-��۷ʠ�
HFJ�*�G�s#��S~�۾�� l�^W��4"�)�:�L=]���\���/*�K�b��m��_'��3�F�$�N�۝;�H�9�{������λvI{�;���_m<�OOѪ�(�v���f��]��Du���z���uu�t�M��Tn�^==�[ӕ�FqW.K��'(��Mӱ5]�VhM�2f�my��߾�?�o������Pd�,!�4��IBd�H�Bwd@F]ۻ�� ̃
"+�l+�F&���*r�RH�!��u.�0x�xF;���a%�"��(��#i$�A�$��f�2�JH���+!,2��ā�6�D�h�cO�Med3�scsr	f�I���"�+��U�5F/.](đb�u2C� Sw\$��,lM�K�g:Hѥ4�2�	$�123(�ɨ����,RLJSn;��e�vI5!E9�ۦn:��Ӳ	"La˃C�n�H)E C���2w\�+���s���Y4J+��!F�	�SMF�i)@7��^.�)�����B���d������Z�]���/���7-7��E�
�w3���X��B4f�Xd/vP�߽�ƞ��\�z�yL�[n9��t9}S�&^plw��(�嗔���z��c��:e��5�.��cN��Sc%��~�[�/'�٧��fŴ;����=M�]f�̹S�v`Q��I�)����v���-�����#e�~R��8`�pn��Q==S���-\lV4�穧�����S(=�N�3O6˪�47`�/��c�q[��8k-��D�=��f�wp��f��P�`n���JN⺂���݃&��fj�ܓkR���S)�m�k�9m���PwO�;2�o��9�|�כ���V�jJ��ͣ؋��e��5��fמ3��)Rs�x��n�o_o)�6�����̀��!k�e���{��Öe=u|���o�?fjjl1�EL{�ܯ'_-������M+�vͰ�Ȳ��)�∳���j��"�J��2jTۆW��u:�3��z���Ku9�mY�5j��P���а�M4κ�z��.b	��j��E .KXz&;����5t����_,�\j���5��3
��3S��t�ӣ�Dz7]<E�w'AÁ�;�A���D��������.e���Xѱ�p�}�)�}�'ʘ���"f#��	��b�:���t�<���^�\�k��k{{8$�����]�#7Q��C��*~W�+��YJ�N��׬���[�y��M?G:ʹ�m�'�P3[ʨׇW�T6:���B���s�͠�������F}�����w���q�k���+>��sn�9�\�Y^8�\n1'�#!o8���V��QX��)����Ϋ|�<�m�^k�L�t_iMf`�{��t��v�]�΢nr�Jc�
��HWKM��z�x���`�ȃ�RI󀧺�����|VVx>�6�L���+�Q�ug�'�.�����&�r���/��5�VQ�@gr�dꀗ�P��n[jVT�.p�!Vᬶ�떟Y�miw ]F}�*\ͭ��Y=De���fh��RR$��A�E/�J�N
��zr��;�خ�z�h��X�^�j�rm�3�ܚ�O14���μ�=�p�H|=ʌ]M}|1���oR����[���$��Ӷvf�Z%��Fkn���`��V�L2-��:.]ZFNL�6Շ�3{�.�u�ew�L��{����pկ=jOo�ڡC�#���B8�y���{��;:�a�v$v4�Rޚ�)�<kS�^y�K虬�t*ӛ�-͝� ��|��+�D4'��Btyޅח��_�{ق1��w%��|���x��B��K��hȆ��Ny�LeBM*v4�0,��lK��IA6&��E�p�اl�!u@���A�O���n���/%M�8�+�Z\�麀M8��4������>T����@<��r�p��w��Uf�p�$���֦]'�jL��k��n']�1�l������:�}�M'}̾{9n=ˉĶ�umB��i:��N���yU��iS�����z�l���S�f-��ʞz��⽬m��NV����]y�G�N�n���̲�թ���,>�'+~�:&�����|�����U�H�#M�9Ɔ��O&�Sq��*}�E��M���5�a���M�Ɖ�����v�V�tS9qce:7�����m��+�5��#ŲSv��;��h��7NݍkcHZMնЗ$�o�FVCk�I˕�a+��k���´��~���Ӽ��~cd��]���*���4L6'���U��w��5�C�դ�/���ަ�Z~閐�z�ᵽ�;���s��`�_;��k����f�+^tș)����c��6.Z{q+�m=Y�wi��*�.\�H��<�YIv;<�۩]^�J1���m=/V�{>�۽�5�mJ��40,\��ŕg�-d2��Kyxᬸ��mCi��-9<�4�Z�U�!�ڱ����FQ�y̫2=�x<dE�_8kv���s��0�D�gu��95$vz�g�dC����G�'�U$ޙ�ny�Yl��]�_��5�lw�ͯ|N�Lf��r��0�S���KE�Mf��o��J�IjA����H������k���Y�B!OHJ�������]�����ɝޗ-%�uxey�j���!�a_��R��Gsއ��ɩB:�mk�jTώ
�Af	��y��J
L���0�krs]���Ru�Jl����VCXa>ʴ˼R��F�'�aʂ^��5�Oc]�w�9�*�ck5���a�8�v5N��|��887S{���xT���G��d�+:��S�s?�}Q^?7�γ�~�6�R��mo&�Z->���a�n5�#q���Q��.�t�X�!�A�`�̹�{[�;ڞ���E�􀖷Y����S�3v�!����J�Ћ�m�b��G*�/6�MYϗ��ݭ�B,�y����F䙶�B5n���y٬c_����Q6��ѓ�@o4���֛w]{Ό�&Tj�7�w�U�W�`y_t�3N�(;����!�]Oc����l��63y�I�q��kw
e62^��n�o^�DFU��r�.:r�̒s�a�w�CXo�nr��]q�D�v$ͪM��Εٶ����TWT�s+)ۄ&������ρ�Y��	^�j�cb���"�|�n7�Z�i�;�Ő��~��5��G��Bd�8zk��~�͓E��'B������O��oz���P`>URw�ٲ��Lה~�7B�m�}S�i�n�WYv6�9����b�����Yw�e*}�ͤ��]f�+#V�c�U�x薊h��������@�5�f�!�)!8��>��t���|��pP��1�l2�w�q�3D���C�I�{�;���4������{w��Ev���mƸkm�[P��J�(t�y��s$�����YOu����P����g\��7׼���5�7��*�?�|�U����{���w�S�����k�e��c��C�s\��A�Ү�.Uk۷K3F�~�%>{7���X�!o��W��!�c�f0X�
~�ܾ��C	���?C(�@?*����j'�m\o'Q�ʎ\ɡ[�r޹��V]�iܫ���u5]=���̄ہP�߃�_U���N,z`��{���������y"V>}F�o�5	��~Fn���t�Y^^�{%�ߎ��I��go��fy'��>�I9��ᚶ�kw:��{X��2Is:�.�.&4Z���c��g�q/r�y���N����5/o�k#]�ǕJ���R�^a�;�*0�Y�.�W�����SojJ���&���v�7�:�)��z���p�z�7S��j�$�4�6�_�e"��sc8`m���\�|�:uN�E�%`��)���f�y�1�"�4%�V��p�l�&t�assmΦ���Șzf<�,#W&��3�+���5�f�P�N��������a�]bΚ//�F��7v�9~�f܃1�k�ӟ��4{�`��t^�xkE��X�6S�ꤷ��;2���z��W>++<a�t
g��֥zj>�A�r̓�wn����frd�p����4���6��EW�q��5�T�G�`q��Oί1�%�V�(��u�lT[����D�����v��@hPK׹-�r�og]Wgkg�'���놭D=kͧ�m���;VM����^k���뱀[.�#95�J����Ӕ��{}�=k�C��&�/�ںIW��z��V1Cg�ܦ�	h��fx,�O�C��p>�V�x��LJ���l�:$β�y�;�L	KE\��[��7<6�WtP��)o���z��x��{ʳ��B#�% ��q���8�n�k;�c�xNӄ��{�3M���R�p��q�T�|5�y�S�/GkC�w��1�6%eC\T�}��ؔ)��{�"��P�&�<9v �1�-�3�@GO�S��f�L	[����N��75�k���4aC:�P�LG��Vw���;pڃK�k(7��tV�swh�=�rZ�&�&�r��_���Զ�2��5�����vG!�_`��Il�y�k�'�Xw>=����{W���V+�N��8f��j9�hЗ���,i�&�^�,Ɂ�<�wB�k�3�"^eO-}��{{6�/�8e��2&��1>z����d�V�9h���)�	9U�j��G7�����n;�����ⲤL�m�K����r�g|$GοN�[������	�����}Kjf��Ԯ�lg���mo_��VU���c�>3h&[��o��95N�p�=g�z�����M���ߥvjx�l䱻�8E3�z�-�K5���q��]���9d놮4�V1�Vᬸm>��Ϯ��K�@ʯ,���<Bz����u�u�=�;L���hn�1�YqB���KhCwk5x�����[l�:�A� :J�*��OH{)i�)<N]�37sgFE�y�啯��H�?s퍧���z�4~I�E����K�$���-j��v�G��]x�-�i�G)(�+���/���CB��qve���|Y�m�qg�N�L1K��1�E�W�w�;7�+��WV���]Ӻ��*�R.肳j�qMWs���l8�K��+��C"�������BO���]3���[�֤�7S5���v>�lf�C�r��0�S���)h��G[�BA���>q��!;��Υ��jZW浌���r��"��$C�]ڨV(Nv��j�g �r緖�@M��mk�KBpͰ�ȟ*Ew/��i�>ٮy6��f�=�6�j��]����h����I��7��ml�L�U�ӻ�xH�{�C��{aU��̹�{[�;S�m���{w�uJ�W2cN-�HT�xG1���ˍ{1�����r�{"��:���䃣&�J��8��j�#���s�z�l}Q1W��*[��әʌɣ�.z]�(c�&�/i;�2��q�g���ǚ��\j�S�ĸ�d�qZ�!��]ѵN%Nפ�2�McM�
%��n�u�te337g����{G����k��8�=����>�aeĶ&��!���,nq��}d����g�Dy���V�c>�g%Ϛ��BRm����Ă�S#�1S�q`�Bn,��yQ�\�#����X���8����p�cw��b��J�S
��u9=�S���<V�N�&�+�\>�*&;f�&�i�D��׻�=ֽ��vZZJ^��|�I�G� �K��N�J��Q��ƛ�&c�7��-��ٝ�j�����m��`l��\Ϭ��Bet�2��DФ��׽s��S}e�o����[�(w 4(��ʫ2{͜�����%t�I�r����e|��k����[O9m��T(t��I�id�)Woӧ���jy4�zn���ܷƠ����ע���9NR�AT^M���>oRr�Lu]ޣL��C~��wT-}�ZW���EC�v����f�}�6q�f^�/���|�!��^Z���^[�*!&��o��:g/��\�b���4�D�i=��Pg���CA+\�����{Z8rb�r,�]N��r��[�L��Pv�v�ĪD�8��W=��D0/g|�劼�djC��.S�F�����e_�:�I dݢ-�h+B���rGGu r�Zz!��y�>u�Vd�&1� �%un���`�X��n�G�sԔ�\�-����zQ3/yf1�++�2v��|�T��Ʈ��h�dw�`Kwα���9��}�T=�=������HX�0��6�Kn�L��	N%
�4��c�d�Z�	��Їw����%3��:t��m;��ڎ/_Y�
	�߆$�F߁|�������h���5�z��`s@t9B�r|���D�n���-�p�ҫȉ�qH���-�M��*8dw�lWgXVX�I�5�3U%$>�N�u�tտJ�l���������Qht]GFP7��4K��e@��-\�9�i Er�3&ӑ�t�{-�^��A�i�̼>bj��]�Rλ?h���wL,[ht礑I'*R7�N�I�
VK�RU�,����	��-�Jn�U/�p326�U���8�h�Xf�W���f�w#��7�#w��i���Tv�n��&U��������&chD�+�tEjMS-��\�`���b�7|��T�W����3$]�H6k"X�mt���0%S-6���J�z�p (��2�퀶���I������1�_���w��0��t)�{E��dز̬���h'[) 5���gN��G"]�72*�髒j�؝k�\t�h�o����6�:�����#'65p��e����v�
�k/vie3�׆O9:�j6���T����.�Juo'%��.�����,f��̾��kt�qТ�\�9�xWk�{nE�N��m��8�n�7�[��Nr�a��qJmf�sZ��a���;���V���2�����qR�g�9m�ﰪ�|�r�(��6M�o�wXb���q��Q	�B��U��|��zT1���@�:k&�����$��TKZ]���Y6	P����u�D�49q��ASȊ�޽=�Mm�7+یNs�ҨY3�ge;�+9�K�Q�}n>*#G����X<c  �e^�.ٮ+n����M4�Y�m�4p([�*Wn!G�*tMK��+I�.h|�u,��Z��,��ӦN����U�{o$�͛e%�7�Ѣ�� �����`�.q�ˋ� �:��,�mF��ڙ�u{�v��f��V��5�AO[�x������L؆�𡴫=��T��Y�[�V�6smS�*�3m�D܋r�c6��O��u� w�9G�$�r��5Ğ��U�L��'�[�-9بP�b�ewS� �pb��m��.Gpe�>�����gS]���˲��|�������j�:��w\�J��.K��6����,XD6�J@U���V���n)Է>,��Ah.��)9Hb����v��=�ut�1�8�-��s����f�K��:#u8໛��f�B7E�ZM���u���(\���h�w`�(��A4��oj�R�1��d�"8�Lk ;�u�q���Z�����rd��E�s3	(ƚd5�rhz�4�(
�&x�]۱�Nu,Ɉѓd�$����p�˗!�.��� ��
nnS�tb���;������FGs��ɻ�ɚ��ۻ�	��sn�fIwq�/�w]w:�d�̖2���n����e�̑�%(��b��x�Y�D�AN���K�I����.^7M���v]�D�RH9s^.L�y۴ʍ1I�ha4��㢊�t�F`d��ӗ0�ą��B2�u�X"1a$�H.�F�uβc��.n��3��#0h�"0i!��(�(U
 > ([3���Z��.�F�0w9K-�]Zq@�C�^i�j�*�GfZ�:���.h�|�3��VWoRUk����H���Y=��ƢN��k�7�MQ�Z�&�]�3u�ׄLr0-mP����^��nC1{�1^����@t���z���]X�s��3Qm@��yZ��B�cb���o|nlB�QtCg��N 4�e�O=�����m��Ƶ����m�B=x����w8@��(;��s1{�V��QX��2��|�^�d�VksO��ԝ룕��sF���ʣ6ǜ:{���e>�?>�J�v�H�����r�� g%���?'�J_g��z����oW�x>f�g;8�O=T�����j5��	��)��/�o�:ui������*+�u�B"���f�PW��<�F�r��s�q[ᬿ6�\�����v��@m�U�K�t����m\�8�'yOP[)Q�M�jמ���z)�*y:��ڮ޹R�w�d��>�|1���^��Ӕ�5�F�v�$�V���SyY�cW�m�6�7z�\��홪�+u����*���ѭ�q��@�a2���|*�̹��+�	\[͎�N����P�SF���t��u蹣,�k���܀"�H��a�v-�x�R��;I��Mw[�Bg��,�Ӧɜ{�=Nײ�t��ꌢ$B���'<����r��ݙ�w��]���$�5;���x�Ӕf
{�H`�����y�v�rOA{�ru&��=T$S���pkl]�m�W��(��R��n2&l�'L�5x�΅Y�ug8��/a�f�|��;G"aR�v��A�1SIb�c�z��ok-��Sim^�ڍL����CI�Q��p��ƻ#JQ�ژ{mKs��3��(-�����R�;ؓ�v�3Pہ�z{EG]�@����o/%��L!}^����������S��>��Q���zULҫ�Rrdƛo���D��2�ӄ���$���i�NNw���..I��ꨓ��g�\>��·��UqѢq<���H�Relp_�������8��1��2��w��)���z�ᵽ�:��1�PU�N�F��D�$�S{.�҉�*#�+9-a͠�VXǩ�|@���3E�^�i� ���k�쫵��颩Owo7[I֧�|��7��s��Va��Ǖr��P4o�H��{{�s�d�[K�W/�]�X%M�|{1h.J.d���㴊�4�ͨڏN��\��I�]�Gp��4�Q�ۈ�ٷ��gY�XJ5n=�����s��υ�N���Q%uN�KC��qᬶ��|��i��u�g=];��GQ��3���R�Ȏ��eJR�Kyx�=!g
"M?A��,v���u<���<�;v<[��:���k�ܫ�g.Sjۇ�k�7�R�:{ϧ�A	1�Z�#UE�;0375�ʻ�o6�b.<��Xx�q����9Fb
c��'��u�-�]�[���#{��y�M��~J��k���������;�JWeX@n��N�{	���S\��7��3l+�9{NI�-�gR�R0.4��od�/\�M�ڿo'Q�P�Q��c��c�]N\ֽp��X�ڹ�!����ٿ��?v4�ʥ<����e���}�V՞w܃ص�ׯ"�b�wN�F�}��)�~����s$	����TĶ7�1A���@u��]����c�eخycY)�(��xL�[/��mˌ,Q3o��夹���k+�D�(V���6'[Һ�o�o��ٹ&e�>Qơ�����̋���{��z��/�v{L�d�L!f���U�����Χ'��qγo���N<S���{�B���A�P��j�6��{��)��~~vt%ޫ���Oej��.�q�dk���v!U��C1mU�A0�bS�~���a�ho���XD�w:�EcN��ldD�|��lk�{fi�F羽�:b�a�_��a�H$Ty���V�*�+�k����v�q�Snr���^�j>����˵׳��Wú�U��r玨K��V1�
�΁;��xv��Z��-(����_���/W�l��j3ʁ���*P�k�жz�>�#��Y�w����5�[떟\މq�
(>F�t)]��v�vE���C��b�R1�tj5'��OB�y�l�U�Lw�c�Y1P�3g�oM��;�o>�=BzzҬw�o�Ao�����ͧ��y�Y;f�uVo�Sa
c�J$_�e�mk%�B̫[��Ԕ$i��_\�9�QWe>_&�$�eop�/�= �C�{Fn�����Q3��n�V��������۸{p��
J\\zIE�k��l��4�3)��Ȏ�W$����s��=��rd�A��|)eP�C(&�B��Z�m�J�Ά�D���1$��%mbާ��	m�,���5#A<�j�G��BtȘ��z=��z�n8��V*N�5�'�qo�o!�*!z�S( L^���k59��YG��e�Ɏ3dN7��o�A�օF*Bc�ي{�_�Է�wٙ��Ę�ԢڍO]��ծ`דq���vFG!�-i�6Э��T�Z��y9v�/p�j��ի���N���m�����7��5g3�gy��yz,�!�N�BNU}"�yhۍ��f޵/o؜kZ�nY��m��{��6e����_{�EG�Rt��#���Q1XӸS/ L<��~0n^<M!Բ�r{�yLu�͖�u�*<��ҭ�Ug�5�Օ���𣁃$�{��]�N�+RA�~^{�D��>zR��f�)��CU2㼚���Y�}�J�n%���-Gׄ� �k �R��c�c�]�S�,�;i�7vT�����|��{�=t#��Y�1M��"G}�� h�Jҵ6���)v]����ܣA�S�x޻��2�\�A�[9���Z�6��u�ԅk�����y�75R,�1F���T@��sM�z�}q/�]��휨��yv�K��Y6��W�gg��ۯJ���ثp�[i�i���ה�bʆ�Qk]�[��.44	ոGk��S�T�yq�ˇ�ki�)�n�B��N��3n H��IP|i.�TKzj!�y~��͏8ʦ�ɮ�L��;=Q��.L�`+�+.��2�~���TW� ��c�93�r�s�l�t޹��Kf�2�F����)9_K�y9ؖ<�D�tP^Jlf�]�ޓ~��Z�s6��9�S)Txh|���9[��g(S�\�ݸox^��u���
Wu#�l�w�\*ъ�kۮ�Ò��{�;��5{�Y��S.��Q����k�#q��13^&�n�$=��������w'�ⴝMDZp�o�L	��}��2ғ4�au��v�����O�`�4�ƶ�;�+
v��t�*����
O��V��j񻘱��<����@3'^��:]ّ�kE�{�$�T�Wd�vk��o��[���ռ�B ��V�[Z\q&��uL����M_�m
��m/g��I^,�[�G;���1���@���ǻ��dV�Ѽ�T�5ou�tؓ6�P��7�vbќ¬q��{����H�yaPW[W��Tfi��.��>k#]���(��R���b��=�$�w���z�Y|,f�����iڙM��z��ڬ��1g	�Iu���*����MĶ���%���ؘ��-=�Jٝ鮁�,~;{9Н2��F�I�0��U���U�R Z ͑����<�_[�n��>���Vټ�W�E�����>�o�<�}u��Ķ��s9+�r��i�2���M>�7�B�O PG�'�C���Rع�y�̓���c���~nסgC��Il
=��EcV͂6b��ͩފ�_V��s\!6���g_�>5_W<}��ͨx�T9S�AO����*���Ͻ"?j���
���8Ŕ0ث�+�P�h� �,E�'�I�Kv���XY�)��ym���Y:ڀ��A��E����s홢�7�ɜꄾޤn�Ѿn��aJ4��ws9�
��Fuf��X��jM|�3{2X�f���k-\�^�)�뷕�n<�]�����jZVk�o0T6��Ǌ������z�}6,A��pe�����rS4]B���o�b�ͅ5�ڀz��9�x�]*MC�F|���z���O.��MF�yk8*ɛ��,X�n�/RV����ҷ���� V�����ǲ"��9���<�8f!�ֹ��Q[R%b홤��Mƴ{]�=�a�T��'y�f�/(MF�E����v%X`�_r���'8�8f��ʏk�u�L�[P�ШG�;H$��kK�<�f�W��.��ֹތy>SF�F(۵�w�z�� N�bK��EVw�u7�cO�L�.���i���`�M��j�7xJ�bf�Ck��f�d��k�����E;���r󢰗��6����-K/���{��>+3��	�<����z:G���2�wR^ݭN�s�{[�Q���vE[z邡�������It�2���cM ���y�˂5F���w61���2�VB��v��V�B�w�i္���7�>��-6�S���*q�������k�_>7�'�������/Z��@[�`ܑF��)oR7�gI�������+kOf@��	z%�ا�;G7ms�m�(��\in��W~m��i�Ρ܀У�k��D/yovv/k�̄fB�sbǮx��m(��c�����H��l�0-	���R�Ž!�{�sݳ�&*�-���+1�dr�L��K��p(l�?r�,��T�ΨZ��}��9KC��:�+]��:L�9��|����(����D�xt�rU��f�{��dͰ�6)��B�Z#`t��{�ҝ4o��*�~�C�`����z˅xN�KNR|�D6�;�#q*��(]�]dXg"�K�<s�ĳse�}�q�mF���4�0jq�ѽtE�8la��Z��d��׾VL�����u�֪�V��[�TZp�6�mD7��u':�n�:�pn�฼�����|��l7�H+(`\����j]��G,���d'�}8&vL
���7c�U���k+����FvHV"��[����z������� ur���9�Uzdٲt�Y/c�������M8���r��������DA��@��y����S���pԽ���/%��P����ƈ^��q2�_	�Yok�{g>�Ƙ��]yS�+^����7lz���y�tũ�����Κ�����m!�2nvbp�������jj�L���z�����z�,d�1�h)��I�`��6�w8W?Q�R{����e���6���׶r���Q���C
k��}u�S�ʧ\:�N����E�k.O�"[ڃY���k��͹﹞��9Q���H�ֱ)���c�z���b�*�����Kzf��E�����P0z}0q���Q-���Ê+�yU"\sw�J����?kk��W��B����s7��bΙ����v��{��l��3XZ���cw���r��!Lw����Ω0&W�Z.`����vnu��U�n�C���Σ��42��.��:;�ZūPݎ��f�CB\�Л��oS�3L��o5�7h%�C��_86L���}�T9�����p�^��t�%�ɷ����o&\|kIݩ���~"v���j�tݏF�?~�n���ƶnS�[�`�[�L��v�rX��ak�G����ڕ��ˡzj�!Zȷ�!�{wள��m�Jʠ(&�C0jqRQ*Y2��9J����"�����Un��K1H�,|���)=�9E�iu�NU�@����F'�?��Χ3'�@N"�_s.Q��1㵹���*6�ȇ86�ޔ6Iu���U��t���C�+[�e�Gy��kmom���䨳hb�L�3VD̚)����,ln�J<���b��8�T�!��_f�;f�٢��c�M)�z�s᎜S
׸�-ǃ<R��sz����u�uM��&��ùmE�38��8"ز)�M,n�����c���'Y�\WEAG��1ӛ?�u���{�KJ���B&��ݩ.|x�6q�3UNZu����ԯ�syw���I�ʹh��&����{W(LX�t����Z��Ũ�!1a��\�ۧ���
��hS8f�Fp�M+��E�d�
��tE�(X�y���T��Zr���;���[�U�3]��6ul��fWeI��6�bٖ[ݧ�S�q������u�n���b����p%�
H
ޢ�)R��--��f]s��rH�b䲣�+�\o{�`H�� %���S��YTyJ*��Q����L��Iݫ��ي����2��Zv�2���]���C���5�o0������R0�w,�nF�6Jǻ����*}S�
ʦ�(W�,.�w�ʸf�z=�B5\v�A�3c����U�̚n�#��a�!���M����Wf��\��%��W�@�ja��^Ƨ#�1F�$j������A7؆�R�9vW�fH܋@�q��ԋ�aٺ��G���\����⯌�̣>��=gzP�1�n�Q�p"�������O�[k�;;��qPt�uZ�o�Q2ګ�؅��$�y��5���cѲC�<ɺ�ѱҺ�w��J�b���B�@��+�]>��$^�N���o�dxD
an�V��ݷ��pGp҆�Ѫ�dB*z��ne�б�z����z���آ��t�m�Z�3*�ػ/C�N��h���]�*[����=�Qʹr[cw�p�d�[n�_�&KԦ69��k-����Cs����j���9��-�m)t�/s����tfKO
��V��*��h+�Ð\nȺ���6��	�+�E\�qǯh���.D{�B�Q@iǎ@��F"�$��-S�wuR���|��J}c:���h2�V�剮�巒Y�7ֵ�<u�M�����߿����A����]!(\�"E-:�3+�u8�3]�(�$�&*I����I�l�"�����$(bQ�uw]�;�fD��]b;�qL���9����"�$#ss�S4;�2�N]1��2���2f7g9��ɡ%v�I��B�ݒ�Dh"Q,�
i&��%�h���$��31n�Ta"6#%D�wtABh˻�%Q�.Ww;�\ۦ�IDA�-�X��@U�Ȣ�\�:rL��2i�v�E����w\�.Q�
��w.��]��N�IK�ܒ!���B���ۜ�9�&�>�}�_S�'D�v��U �Z��˭qcY�q쬤�����8N�2��G[�j&?�q�xè��FC]��9ʹ�4�K�O_���I�6��k���v̢�us����g��Iݴ�RWU�8xOf����=�s��Ű�ȕImE�dgaZ&s7��v�����|yAm�j^U������u	���ۍ{�MN�=`�78�w�	�Dn	��V{$3}�K��g_w�1��-m1^~��틨�H����=��/q��ذs��Ң�7r�6�]n���=���=[x�3O(�W9b���r����u@r��l��ޗc�J�5Q{Iڙy~i�X�}�M�F��64��ԁv`������]Q�N%N�����ӿ)��/�y�ڗf���y�����JS^|k��8~�J���.^ؘ�sM���ܮ͝ν�k���v�ZYft�~β�)������z��*���.�d<��h�W^��+C��.U�X9�dt �EЩy6qǂS�q�����<�g�֎H�n�F�S�O�V��� ƍCڪ�b����[��c7-����UC/
޴EZ���Vq�{3E��#I�)2���wc+�4 o"�n9�),�봻�\^{GU�Zo��T_���_T�
�1*YO7�Bɩ��k�]�
�Kau��kͧ��7�P(t� ��޴d�ڿ�{�gVoyz�i�^]�zw��z�א���T�*�y��(?`tyu.a֨��
�gV;�O�9}��g63^3z�L*��q���X_n����q�R�}F�Ϲ����%�^kj_���]����9Xܜ�e5;�R�tP8^���z4Q�us΀����V��YZ3�tQ��S����[N��3
���!k��]����h���4��ˊʼ�����.��q����* �����y�슋�E<2Kj�]ܚ�{9�o���*��kmT�Zh��B3���ta��`�&��MR�7V�䁳��%>W����'[x�3^��כ��f�X��V���m&=�,��T���,����NOq������O���!��j�o�H�ֹ�C_���pC3�"Q���/����ie
�ա�W!����r���r�>��u���ehZ���F�TWk\�[��h��v�]��v]V�`'&fXْ�	wa=f�mΜ�5�$����^T�ѷ��^�h�֜kY��T{0�s���S�/���eg���̘�O+�y���Xӿ)��x��e�Bf�K+f.RzBS�=�mN�:ػ��`=ꛜ���^ؐ�9�8]�����M�ʝ%�R}�p��Fv�; *�s���j'z�z\r֭Jg7nn�qqYs5�����܈��_�vםom�@l�s ��8O�;ssɽ�p���Ľ���V�B�p�}q->��9�ٙ}�5��s��H��u��ܲ�zv��9��놝����m�����"}΢��e��z����_60sok�=��׋O/���|3y�W�k�qWO�����/��e
���Q�H���?N�9�^y^>nul%��Ϟ}�rf'7��e�I�jw����<GN��C�����J��R]+�J2�4��om��O�wx���V��e܍�J��p*U�@�\U�ǥ#�q捚����B�3��3y|��]Or��J���ik��C8�����/Y۳.3��7�:�JM�]m&�:���Ɛ��	޳�+neϥm�%ZN�q'���5�wU%kyI��)�o8zچm��6�3���{� `>��ʡ�����gR\+wGB�xO,i����5̶�5�v�ĪC���/&-�SU�u���r�m�e�Y/�im\o=�jn��Q����I��~F��1V��_e��_̵�I+1B��\���um���Z�m$��ӆjP4^�O';��=���e�ȴ�݅������y�����u�����$r����0
)]���ɓk�co��_N�o���+~�Vv	7��&�4��S[��+s0���;��}�Ҙ��t�Z�j����󿇸"�,/W��N��7y�Şq�1zv%cUŦ�K���ٮ�f_��<��7��E�Mx���{�{Wa��'�ׅ̎GP��sM��?�.SZէ�mq�5��q��׫��/Ɣ�ڒ��T%q]+ب�e����/�S��6����몽܎��rF��
�+)��Ѫ�q���*_�tzVh��.�2j��A�*4�ɔ�K�f���fI�:�i�˻�dU�qf�W�i���Q��N�1%�ܩ��Ȇ�:����+��խ@�`�r�6��RG�>3��*`�4���3{���Oٶq��5��H�ֱ���Z�������H�ЍB���37��a��q�i��o�;�ϼ�ի�wԨ:���C����;%v<r�_8�YRe4���z��9P�*:}��A�
xg�I;�m�Rĕ��]�˴��~��o6�b.<��\����(ϑ	O�G���IiI]̱e�o������u½��ƥ�a浐�`m��9fa6�<xQ0����˰lT��vTS�#uxeC\ղ�;�q���^4�n@&����o1�^�gՇ��9�c������[ɭh��}E�÷�J/Hsy:[�������V�7��1��+aՕ�����#um.z�08���s����oy�lܓ2�(�Pۍv��k�&9��[�/���ů�6X�9�m���S�4�f�N��W�����5a��:-v蠔�^a|����}����V�S�Wj��m��G��;+"�e\���n����~��(��WYʷ��`�~�ʷio{ьY�� h��(;j�7����:55P�;�Y�L��V�흂��G��(�8ܬQ�ʇ#�15����i<��Jv�WT详p�
����*3q�ˏ�]��[T��j��w��Gֹ����t��1��t�#�И��{��yT5��Q78G!w�:"���M����u�q�z��Y�5�c�7���*s��o� �wCw����W�	I��;�����֫�e�ŮMN��w/�I��a��?	�@�:^QΨJ��z��:f�<�t̍�ju���S�t�����oUM����� yT��T]Н���/T���p��iw�x�zި�����P���@l���;i��{t��2���6��}�iNNF���\5��-���ͥ:��^���)�,i��u��ٯ|�M���ס���v>�ʈr��`��LV�Sw���~�Y�K��'��5�{�!�J��{��ɻ�}��z�����	m���w���sٸ�\��U�'�}%mI�:�{�]���Z��3�s_��(+v�Q��K���6�d[����,N${٣��n�q��X�T��z��'�U����*gg5�ͻ���>seި��sp%�u$j9�i`O�lutm�q���]˫����g����S��j�:��!fἏ���]�O(�bT��Z�{�l�B,�x����>�ͤ秳���fwE�8MMgf����q�ѸR��2huɋ��+��E�n碐LGx�7}�O%�5|�4��v�ϵ����;�LV>��)c;�e��×n^���]�iub���m�pʹ1���y����y�7�5�^\�t��գ:l2 R��n�������~�N����c����}������q����-]�|��Ȣ�:٨4%� .�nP�n�q��g��[��V��:�(u_^�3�|�A.+�Md��\�Jz��������M!u��s0�Us��d�k�	t�{s��&�Z"nqj��%�3p�С���q�����y�6FKI@kܓ�!��҉ћ>amh�f��{�a�����3�e�BuAd(nC;�vZ�N�3`���� �f']E�Ĩ��ڝ���8 ڇ��-1��F����t:��R^���i���(�&�pCZ�(��M�9u`P�rd���}�f�ΐ{�;tH���"�	�/� �K���:�-tB�ܱZ�eݚC+s��V'I��Wz��*ɼX��-4a��#\���SRd��Q��f2WGpf>|(�t�_nI5��	�R�ڝ�ubY�B��c~ ��3�1�S�&sֲ�2�ОW�F�r�=��������Z�R�^�yꚮ�t@�
85�<�B�8N��t�gwM2�
Z�r�W)��S�=�<-��B3�^� rvO�M�R��:�K8���0�In���Ҿ/v��o_��V}i�zn3���yV���r
�L6�e�|Z%��{�.isP~�&%��lt�~��|UK��b�&z�2�N�c�j��{�(��	dn-�J-�@�h�a�H����mh$�oWQ3�^kX�ic�-��!6�C\��D�V��0F�
�E;��=�����it�Q�]��Uɷ�D�J�f��c���>7��.�ܶd��ܤ�L���!���r�4�2��=?L�ə���mΌ�k���t��!��d7��H�g�p"��j�Uyu؛��!c���Uo/<�5?�>��au}[��J_��W��q�{D�NE��Z��?V�n�2�~p.�~������N*�Y�U�U��2K�p�P��n�y��p����X�Ƥ`;t�ۥ�������y^�Sy�=�J�~�kn��o�X	6��V޺�	V^�,m��[-����}��f���p�+ه��̫{1��[�S�b�*�{.���z�ld�A�(�Rpsg3�r�:Sc׽�Zv�h͍��݂rQ!3j����!X��9��wP{^_W9'8�p�̼#��{��\h�������]�Ϲ�g��+�Jg���ˈ<���It�n���o:��q�l5��u�3I󚦢>�rS�����T?i�'��^�S���s����{)���u��[�{b��o���N}4~���(d��S?#q\�2�~kE8yL��&J9��B8��Y^"5v���
����m�'D>�-܄3��0N�FL0��nԻm3 ���hO0)<k���ҹVo�#"V(�Y�O����W�P�$�a�)��]4�w=2�
�v�^OZ�H
�")1];b�"�R��O����~�gƗwJj"KCu�+�Lm!%�oo����%R�TKފ�[,eB���RcR"�O��/r�p1ĸ��u�X��W$,�;���};Y�D�ՠ�<��/zxk��=���+�\-�7`JJX�%�$JM0��m��ݝ�o|4+��̈́=��y���2ߊt�`=.�O��[!
�&�%�N�f��p ��3�BU�8�w4��VlK��f���eYa�����l1��
���	���o�u&��h+��T�u1|��df��_G�"ĕ�L���0s��M5�oc�+s^mnF��{6Vdl��'+�eiR!Y�e�r�t͏j�8uM�r4�݋�YK0u��ν���8�2��d�����
��foO:M���yn[2_Z�k!���<��-<���L�u�!-N�ʤ����d8/�Ij=�v*,�9�ݦ�C�r�g~L}pԾ���n�J�Gлb`O�(wF[��|
�¢^q\~qO�$Y�ҍ��cZ�2]���]�p#[�6�X%��n[i�ܦpU�u'����./fs����;���'�_M�j���%s�hQ�rѰ��y	���T��\��͊e�����	d'����Ջ���+/�M����<�·P6t}'$��T�d�`+ߞG�S�����ג�{�|SXg� �V8��Wl�+ �`7�5�,��|uC9�G9�t�rܴ������vF�S���5eP��&���f^��{�^K#_VL���)\����T9�e�tyƨB�V���]@?�ww�3�M|B��M*9��B�t�F�=�P^���C��- ��[�Ac�3M��m�l�1�� .Y2�X+�h�k!���:�,���Q+�I�X
=<�I�<��]F])��#x?T{�2Q���YB�.s
�H��Xܳ��P�u7�!���<b�m��9Pj)�(iw��B�����y!�����ON��*����K]]�ƌ֜а:�qg:�1�p;M�T���h�RJ���&�R��(>��gQ*�{;4<.��,�]���:��b.ruk7]MSc��̏����ާ��"��)�����I�|y�:��a�n�F*�n�G��u���T��WX���W0iz
θ��rJ���{�����m$��]-� ��C[xޞ�yh���m����뼕�r!��Jwi:0��:�	V���{���}��e�.Q,sxݮ�J]b8.���&���[�"��ӡ��쓃�K���ope1������k�VV�9H Z�ٌ����dhC7���Ф�cj��t���Z���.
��o+�s�3�+b���0�|2��u ywt��>�
v����0�);�_lf�d�o�Ʋ�P{��)m�*�m�#ǔ*�&��B�7xQN,�݉��w{J���6x/z�W�}�)}i �\�z�c�/��'���v��Nj1�K������Ta��/��@�tr���MV�&^��)ӷ1�2�:�G{z
���%A�[1�Qgb��l���Y�W��|��JR'v�k,�����-v� +x�e�����^���)WPce8i��
H�3�K���YR����l�&<̮'�A���kf��m���Y{��asEԺ9!V.Y9���R�;(���`�2�[z�[?uq�)��ʙh��w��%dJP���t󤷉lXv�Z}��@mb��ݰ+3(n$���nb}�5:��*J�R��Nu7*�&�Iyʻ~4�A��sR�N<ۧzk!�q>�n$5�����j�eX��� ]�+BZ��Ѿ�����.�u��{���f'f)Z2��{��'�m6P�C뿔6V����>��<�V`s��hm��w�.	yo��Ty�ٔ3ws~ĵ���Y�顿�i���u�lP��&ZΎ���x#5����� d�r.�[�E����j�{q*u�e��V�� �d�%	�ٹ�\bV�F��t�w����b@Z���<2��N�	N&mY�,n+�*��zc���D1Fq�1ˊ��B{՜֛=�UZ�U�/9s��c6�7Cb{��>�Zn�9!'t�[Mݯ�#����c��� �yS��lI�z�N.I�1�!��n�p��~�5f�#�n:�DOq�
��@�>ڶ"�M֥�1�XS�:�^V�4���w��ˀމ�w��;S��7���cM֊��ʚ{@8��%f�����;0r��:��l����aT�(D��Bk�0�|�EڠpYp�Ε]9�jmĴwu��Q�Щ�Ƣᜩ6m.�{�X\�^ �KLK{��"��X���ee�[j�7'��ߑbxv.��]�u�8�wv"��tH:F����Cwr��wӢ\�4��\��X�@�	���D\�АPS��Z�1�[��2.��+��cr88k�(�K��b��H������ruwwNp���P�c�r�͹������)).vd�����.lX�[����p�H(%ݺr��DXɋ��˦���uu�ƺwu�p��w���6���:ls���wut�9�!�����nE"Nt\�c�u��.ݜ�D]�˚��T��7wS3�F�X��W6�v㺅q(��{8�m�W�D�3QU�����\ܬ��
��[�����7.����Vs/�L�aql��l����c��vj��?W)��A��ύ�tK�l����`/U�ex����BҮ�g��O+*�Z��[�.���0)ܳ��Y������BQ�e�B�{zՊ{B�(^�R����.z旓7�ըsDiG�Zy#&���]��C��_9�t+�}����������s�z�VR�9�����0ܥ�	�c�$�H��xO}=G+���lQ��0�}�$.����l���ޭ�&~��dp	8�@bJ1�YR�1Ģv\��9��cOhɆG	$.�Y+:�����	vk�[(�����'w�\"���1���c�y	i�p�h����5`DJ���A�ǄСh����3��-d�fp��C�*��́Q"L3ӎqo�+"E����W�l�x;�����{N��]l_t�*��x��|c"5�Ј�9�ZQP,�NS����s{�3���C�(��Q.�L5~Z�O�t\Ru��6ds����OK�e5_(|G�y�d��'ݷ9�� \ׁ��׍a������a�VW�o�R�A�T��*��̮-� f߻�lT� �*�4��D�:´�*���()�k��?S~��}��eLQj��Gp�^d޷a0���X.�
�0�q`lָsd�:��h8�I3n�D�A}17�DZ��y���y�Q}��V��P�S���<�ҏX7�J��nN��R��Rd�xv�V-Y�ۚ��:x��(-��h��@i��m�0�l�VZ:�ROH�}��T���:�}8ۮ�h\j�#  5�؞� �6��6���OR�\�3����M�>h�%3��ڄ�<�˟ν�����l�6���;�$D��D�(��s5��m�$�}NJz�'x���8FZ�D�S`P�KR�C�S$RP�YmX8=A]�`��9��N��8N�є���IR�4�K.)��<�����G����E�����/�YYTz��s���#Se/Z4 �6� ���3��Y�Һ�	V9y+���갠��;��gr�du����=����Өw�rY��D�x�8[�&�����s�;�a�}���q�)1[����Z2ҮM���H돪���s%� �|H��[+��蔆��\����e�h�L��Of�5�(��	F��K$��@� v�����J׬`,��勣c&� ��x�F�h��})	kZ!�Yv�! �
�97�x��j]Jk7�ӓ�R��ӵ�uV4X�.�H�/,{�4���]i��+PZP>y]{��{6�_�~*�(d���n� {4?�'g	�\�1k��u�&����5>���
���.q�#
�u�^M��(�&+vH6����e�&��,�n�A��&M� C����n�M8e����J7�lv	l����̐һ��%"��_R�v����f��̝����\�'�2��0��%኉koFEk���Gu1�]�c��[A5د>q\s-|Zg�$'�RӮ�%*���W�3a@l3����a\Wպn)K��J��Ǩ�v�C]���r0����
҇@�Z�q�|�\K��Az��U��}A��v4T-C/�\)e�t��1m��8Ҏ�2x���p���OM��
�.��ӝ��T��	"w�yŋ�'�Z��:�gUUf��wm��	\�0�,��k��3u��Ci�.�ͭS�%���6����|ވ{��Ěoq����9<�}�[Ϡ�u����w�g���uG �S4(�2��Z�"�����*t�%P6���j
#�ݐS�889�	Zq~��E��7��q�}Lo�\/4y�H���������6��&�&ܨ:%� @,�5U1~����]AR�Ѕ�	��İ<�Y��3o�t�X�K ?d�SΰS�
��H�J�3 �L9�-�K�`��`�N4g��d�&�)L�X�n�� ���D{fK�l��1v��E�v�RT��*��vh#FC���j쾀H�}��M�}٦�"��j���J���WJ;�Ū�.vؽ��	닎�He�<fsy�D���/�*Jݙ�CNpѺ�/�n`o/;�p/GZ�3�ҬW�\r�@u�Y^�{��a��R ��,�S��n�c>��S��1W��V^��{�Q�e���tSi�ic�/X̌p1�%�1;s<;{CM�M����O����r��1ľC����oD��c_)����%p@U�����AyL��(Zϱ�Ԯ�t��N����l�@r�j�1��[�N���d=��O�̊�[� CE�%Wk���0^�l����A�2|䶩s�<{!Q�-lީc�j�1Ϙ��9����2✃��fG ��kxKS�r�.#�x�C�~ʊ�պsղ�=z,K�����Ⱥ�[��͂��-Y��L�D��E����g*��}� ��+`�������u��*��X���$_e���h��ҰMdܶ�w)�|�����y��3�,^�Z�B.�������s�q���f���t��fBk'��U�ɣP�Q3}��x2�_❎��Ee*p���Y`�X8Y���N��j�Pm{��]L��#�'
1њ�!9�Yzu��J���/|kuڗ���+�i���%���C�@ݸ��H+K-iyݥ��6�,�Fp�%��*G�����s��I�W^��Gt=��e�:�1�h������Z��5���SP��Ge]�N��O�Yyf)��p�i�z���&�ս����;�fP��b�kM���-��<�w���'V���Q7��ɒv8^��)�F���g_}{ppL����T;�����tq���`D^�g����~B���q�Jn{o�c����7\)vT��E�$񨒾5UC��G�q7]��m�Z�
�q�Z�L�V
�3Z.�]2�d��B�O�N>�8�6=�������,�V����]ng]��+Ӫ���W�ӳ��wD����X)�t;��j�}�q�l3>�9��귺O�֪�}���6j�����
5�jДk�e
u��V)��X���/�4�/��l�D���\aع(ה� ���E���p'�WZ�$�XٚT*:���0V>-��|�K̡C�G����0�@�Fв��|Q*��)�6f��<��˦l��N�s i��(�y�,c�D�/� z�����I�������)�u�M ����,�N.׽���$�\*gP��7�~���y�V�`^�uW�3�����+���#�A�\��0�;)Z�m�Yyɇ�_��43w���͠M�=)�OZ4^u\@+\uc�G�Zoum#w�J������ cV�/;[NĔ�d�jNۙY��+�80+:�s��	C;]W�'��X�����`�t�jx���y!�.lҧL�Tc��Gp�͚V	�r�e^K�`Mq��w��K��*$Y�؝�n魲nꑎ��ɤIB�?K���A���k%<����7-�ܦp5_&�D���sٝ.�u�:��*����xd}���Ei�7�U&�����O�t]'\Og���>���N���
GS�����kr��&�$'�6�(�>�6���5���w ���7?i�Z�U�PU�w��j/�gmM_kI0�u�؍��o�F�ڌӿl�ʹ�iK'v���P~U�YU��[Z-�^!͎�lN��_�c���vE�T��˘ǳ�m����B�N�눹��4�f���>�%ǵu�9.+�P�Ɲg\+	L�,��-��/ҥ��/��6~��}6�E�����5!}�E�����k������_zfè(+���LgC�3�����q�J�^d�CkкYnA��ȝ���6j�؁HV2��$�bOO|~��Y�����w)O�X�G=�`�#�gu�m��K���8�;�rQC�J�2��R$Qӻ��t�-	V9}��[��hU�p���G?.M���l]b��':��)���n��q���F�0�3Q�1��UԶG��j������o8���͎�)�z�]r��2��Z�:�s"��b��m`�u̶I�Gw}RU�Z���U�*vST��F���1Z��2r��3�C{_2��*:z�����:�~%��"ʌÁ0[�&�J������8MͶ�1�Y�J�!5�;�+�k^�+��/�F> ���#��q#����f��꘳�!�m�IK_ik�A�Z�:+�]���ݚ��=�{�oBѸ�	(�|F�0�ā��5�v}������ݺ�����&WSqJ�G�hRЖ���l�%�"�+�@.s.��P�E�G,�Ft��4���`KgO��)��=�WF��͎�,���n[2C.� ��zܩXd�gf3���c<������s�&��'�d����kkֺ���u1��ކ$����L}�,���Rɳ$���_	\�w-�����q���ݒ��6�B��-{ջi_U�ګ�&N����EG:J!`�������<n>�j«���� �_;�� �q��W��`K�f��b�O!-Y=�U_i9�G5<�`�k��ܛΖ��ח�`�w������5��}����'x�d�<6��eLA�8
�)��[6��sD7�;8x؄��t���	F~�U�S_瘪"E�6��(,����Yt�����#mT�{��=;g��*��Ҝ�k�o1ҍ���f���;�ZAE;�Ӥ4ܙ�iXԓ��m��x�ef2�uC��n��n�D�l��,�R1a��x:��nZξ�����QӷIA��Pu��t]T�Zk�O;�_Bq���N)�G!�g7���֖\]fk�7�e6����h�eA�>��-Y�2�������9����o��#��<�������b~�i�G�B�u��knI:-�G;�0-�8��^����L��fP�l�Ǩ(���lF���:kLW�,���䧝`1�H�H�J�3 �L;��-�c�o�2mtQ����+��R��L��>�Y,e�t��E���`W��gDs���a����j�o�K�+�)�w�o9�n��E8�Ҹ*k藽�!�J7F�i�~H��Az@�4�u��|�7ݫft�U��Q��#�=DLOθ/���s�����GpgUq�&���Me&"���o~*m��D�ѵH�d���˽h����Ȩ�U��,:��dm���61]�_ꮻjZ����=,��!��'�B�㧡�h<F0����c�
�U�;ާ3��,�Z�|��ͭ��o8=Y\"���]%ЀTΊw�^�-N��YrB�OT!�\�z_V�ta��o��_�n���Ǟ�J�C7!l��yJR�Y����"�j퓉�s�j�痽��3�\��o��G��v0�f溸�p�#YM��8�W�u8������Lj�J]8��tC�����j�Zuݳ�U�qU�1�v&K�����*/Mfl*��W��V�~�r�N��Ւ���\���r��W
�ylV�<�@��3B�NoU�v�����rk+��x3��}]�t�/�����ۅ�ܦpU�tD���7�S~��MY����Cd�VZ2��Eń,��X���TsܳF�`)�!5��ʽ�aXj��Ѩu���9��S|�-A�fvJ��_�͢p�7,O:��o��[Ϡ�|�F�`U��#��_��98.�7�5k���F݂�r�{�Qznj�Ѐ��[����Y5��]��,M�WҫK{��d���t�;��*rQѯx)�dk��82BvAn�!�ZF���F�v^�?������cBdG}>�ȸ�w���Ts�Q��A��nT�i< �j��n �cʲ�ԭɞ�n�iq<GgKvt�u3`P�W�A],�KM4|������W�_C�����WM�� �ħs箆ɂy�ӳ��tK���X+t;ya2Y��e�8�h�M���dVf�t)����p��@�Pg��P5���9鯦-��:����t/q�j����Q�R�[��+�ؘ���=O�!������e�c�ls�@+S�xY&����m�ݙκ���3�i�4�.2�hM���H�ɹ�3&�òZg$ɹژ�{\�ښG'�Y�b
kZ'x�y�.9Ro]"�Ή���r���X�����E��É�����l�0J�j�6����m�Td�}$Y�_9�gO��8,{�ھ�Z��%�j=�L�AZ��Wq6�K�����͡���� �ꌁ-{B�A��:@��$���ִ��͹N�.�wH����@O�Q���JX�~�[ �l�$S�������]�׏N�6	&�@<7�l�nCս��I(�
����N���6�P��+S���V�8�\��4�l}��U�Rg$Vi��ᖥ�0+���rP�C䛞\)��1�Oe��GCө�Bf��5rP����Zt_�__�����߻f庛�L�j�M��Z����ncUQ�܉��/��YG�g�3���J�0��X<�W���I�[�����1Zu�}��s�Y���K�e2fK��^(�-jm��$�c��pڭ��n4Vh=��v�C ]a�Y���%K���SהB��o�F��ڢ^�Sb�ן\������A�xh��M)�&�4�;�}+c�~���V{M| �-���Sre�c���pK�3�I�량Cj"+9��n	��ndH�8��}&:�n�X]rU9c��v��h2����U��'��׭��7��4Θ��&�S�B�ab-���\é�)f��lR|z�`��J�V&j�a+�rȻ�T��;ӗ̕YIj��8�:��n�9��ɪ�J`��sX��<���2��:��q�7�ݮ�D��e�� �
oY
��YᘮRk��h۾w(pՊ锰�:�E.���A;xqG($δ��l	�syֺ����޾+���^*q�H�w �l�V�`&��꼉��A�N���\�.��o-��vL*�ٴM��|�$`HpF���T V�jn��#m�s2K���Tn��3�5F����H�imf������	sy�K���V�s��1Rz�;2������sh0z��B]����Y��Tv���Ȭt�|�ʇ��ռ�k��BrGe��}�8�lإ�>or�!K�r���e�N���ƌΕ2�b\��8�Q} ��*+Yͼ����Wpҟ2ou'���Y��^�t2��)�1�v��t�`0^V�:�O�&ΧεC���=�[�Q���@�H�����#�B��a����okWq^Q �	,��mK�5�մ8c����Eʉ�L��[; ���(�^c]kg���ث�#\�ml�Cʔ����9	f.��/l#4]n��+$���n���@�`�Jw�֬f[k�H�t�m����*�S�[�������Si �ۭ�B<���_�'>��Λ�4;Tۺ��9�ţn�lm�p�5K�e��n�Ό7/\:i��gw�t�@���P]M��+���e�4k�u_m]��W�r�.�p8	�f����u�:�w��+n�S1˱����b�>?Rݙ�pd�J�m��+)^��\h��tΫ*���=��5+���2�C�g@{yJE�����jK;��a�ͻ�w�&��C!��	�s�<��i;PՒ~�5�LHL{\Y'�]
}�e
ב���Gr���u|q��YJ��R`n��V4G1�y-vM���تf�#4Q0�.��c�#͖j��u�zn�"i
�a�*\u��`�-��7s�ˆ����lH��CA+Z%n���G�p&v�=�PD�V{�rot�q�먘]ؗ=��v+�(�^�e�L�^m��1*�j>�b*@�����路��w��t\��*4:[ΰ��r4a�1��8�S3�l�3Qb�K�ڀ�ԧSWkFr��r�b.�8ӒN�I��[��õ�\�ПO����m�;�,!Kc�қ��d�5)�o��
R�m#VV+�NT��[����{�)0��ۢ��J��j�Ջ]a���W�PLI��\xih�ySx�Y�t�᮰U�'&���AŚ�������G�2)�Yե;
o|+ov��pJ�7��FK��Y����K4\Z�T.���Y�t݉���U�U*�2V�[�/���>�>�I�I�S��r�"�d��7s�pI������"0�CFs�E�]�8n��,�˩;�P��[�wn�&���G77�
�r�s�[�N���twtN��&wu�#����n�ĺh��wvu�K�tap�W:�]:�cv���t���(���s����t��WMwt�F��ws��\��.����8˒r�s��������3��Nv�9�r�N�݌Ww�s������戹�S:Zwnd���(.��4t��WL9�����������ι�p�n�]���j�]��\��#�܅��]�g]Н�tnb��Yq�w�nr��Wwg]Ȝ�Q9�u4�c\�\�;k�@�B�`�p�zt������hvK̾u�-YM̓�<\Ui���BEK:�T_>"+6r�y敋�F�(�gdʃInoyu����յLKFθV��Y�BuAe��nCJ�S6�c�L�(�F��������eӄ�k�y��R�J��ѝ8ϯ�K�7�(N&�:b�"���Uv��q��W���.F��LX�2�B8l;�q�,]J���Z�,ߩ��<����4�s��p�.�㪳Qp\0R��],����;%G�J�,	��"��Js�u�Jj��.Rv�{;�3·.6�)�[_2��GO\G�HN��N���B"ʌÁ0[�'���ؠe�%�g�p�ߡU��3�k�|��([Z�J1��~�U15d�@ ��^�ci��#y�%��o�k>#�߫A����{��j6�<5�r��L����F��K$�呤
�O��z��|��L�Oa�X�L �	h=$L�HU�R��Х�n7�j6�j��)�!L��fB��fn�Jf#��T�b4^CF�RϑO�!k���O����}~+�0:)�fa�R]��A�,�!{8�>*d!��
�@���d=�*�A����X'0��'Ǜs��t �M��ߊ���6��'3t;{�5| T�U�:�M;�֖H��
[���Ւ�X	cm*X��c&�v8�.L�A���H����B����:gk�6cTG%�h�;:��h�}s3r�l��B����/�fm�K�H#c�&��%^M�Ғ��F�ĖƆ����Ͼ�D�E;��4��خ����n�svJ7BB��QlOo���eᳲ��Ǆ�ޔ���P�<ˢ
�P��kSN0LG�mXUs"��s�񵔕j�ƍ��hζ�m���4(���5��&���2U}��Σ���u�#^��s�i���q=l��k*v�+q���`�NP�m��*"ā���y�mt���1� 
�k%�ٹ�z���s2߮.r�25E`)�oO:�"��1)��ڂ�[�C�92�V5�������q�k��y�۸�}�y��V`��ה�/CEeA�2?+�,e<X������ty���ę�t*����&��p뱺5?�Ȋ���a������<?�T��L�u��|eV�S�r��~ښ��j^];w���զ+����>Jy�#Z СI@Á����Y��
����p�����۞�`��Y,g�:U��]q������dg:��6J����U�j�4����?I�	��\��_��ƣ���c%)���!�-�"�+P^�I6�̋x~��oR�'꓆�=��*.��]V��;a�Z��qU)7;mi���1ky�粔�]B��R;vX1P7�aC�6�pj
��b������Mł�bˑ��,*uϔ圯�w�t�T���QM�=d�yx3r�(}�+��Q4��3?��A�QA��O�D�u���7C�F�*C����^J���n3�sJj�q�`	����e�x�G!��ϐ��L9�:���N��l���,Z�ͩ%룔�g^E�!CӮ9�@R��C[<t�1�h<FK9-�\��@��=�f]�R�&�.�as@.zL�$��-�/��� �Ίw�L�%��9T��x���U7��̷�]�Ew_	����fq�����9��c{VJt��j���r��W
�y�p\F���)�Ob�4e��`L�SbZ,��{��O�&�UiQ��>�q��D�yt�䀛Z�Uq=O��I�\p�
)�^Ϳ)��c�ه����[�
�W�rh�:�3�VI���gD�b�� &�ɴ'��hN�,�	��=�~�A��c�75S����᱉d��/s9��7 �,p�f��nQ/yM�sCM�A�-��ݿ��~E����u.��>�h����^��ewh�%K�f��\ה���j�S�7�D?���[S���JWa��=��`l�Ju-7�.�Sk}��k	-h�b��-�-8�		�@���o@�|[}Y�Ϳ8�eu�q�Y�:x�}@W:��u�T�J8�y�u+� /]M����*r�w^�������_l�?�X��Ey�lZ-˲��N�,q�*L������M�\B����g�@r�5B����)����L|��C��Zлb��߉:G3"���������K�VhL��5L�g1�:e���(V*�t�,�KMzB}�Q���9�5W3���e�YC�'��@��e>��G�S-��ӳ��0�;�XL؋��+��]j��`"j��n�����56R`k����c��gӨ�������JP��}hh�����'���|� �5*�-DX�ejX�'�v<��5���0.�7�Ft����:�r5�m����/��
ǧM��)�+�O��5Z�8%B���d����&:W��U��Ġ�h�4�>��܎/�}Q��0w�����S i��(�yeJX���8/�er������fr�96i^:����3e���5�ol�%%�S:����3XC�re&����3]U����Ш	t	��f�<s"������'��%�%�0'��PKrP�KZ�	���a��@?s�D��-�3
:�>ti���i�q���������m�U�2�_���,Э���X��]��RŐl��3s�O1+6��R���n#�K�:ފ�]��V�s�m+�qX��97�n�t%i�*gK�v���������f�Ȳ����Is�*3��kj��OOL�ukbv�7+)��8�M��K�DV;ܓ�p
]����_���bQP-�+�:ZCvk=ſ�Sߩ:�{=�L|�w?���1���应Y�w<�J;)�֔>#�آ\lڛyyn��BlpnU����-��D"ŦU�5b�Q�)�{�� *��3�c3��̮sC4��u!q��#.�wo�f�V��n�k���;;$@���aA=�mF�`��
�7'"�F��m����B�N������[�_f�5φ��7!��}�}S:�&~�{P��9}*[�څ�א2���v�[f\L����7��*]5�� Y)�98�-�-1�8�_(��f��8���X3Uo������������[^�Ci�2���A�2��~E���T�9��7MՉ䑑QϾr':��Q7z*]>����u�8d�],����� �^Ѐ ��R$Q�IIXB�(�i����L!4u�r��yM�j�\6����eq�tۧP�g>@Á= `���&N����ݭ0F�m��5薾[,eB�נ���� �ej��Ds��8�b��g݄<μ� ��ދ3#I~���ė�����4�G��z�fmuMN�[G�gt�y#ASܽ�A�R_XmY\{e�S���ґ���O�U�����M;!t�;T�u�h<l�U��ؑi�`�Cf����w��
<NŔ����Z��c�_����H����lt���s��>B�n!�����	dn-�J-��X��'�e��RE�6��L �a�9<�^%�c�c����ִC\��D��+@Bo�Igm��y��%ʘ�ZN��k �6�3Ӭ	mR��x��Ѹ&�c�Kg(.��f�Eʍ��[uf��2n��K2E3����U���E�%�ʠ�Ƕ�ޙ��	��\^�	s9sj�l^ob)��w)�y�r�D�E;��mUo/-�ฆ���n�fsv[yc?nB{�*�mn>b�̌�,|�~��߷g�Ǭ���V�@�5��%+�ym���c���rW!�����k:r��O�Σ묯��%X)�O!>������
]����0�%���zfn�������+�^��θ�rĪ�R�Q'�jD���}���zr�q[�[q�ݦ�:�S��ɘM���9�lMo:��`s�3���):$�t�,p5������g꫹�}�eɂ{�k�
;���y��Y$ع�����ނV��_�)��i;_�TީJ�*�f5�����M}B#Eq��=�{����m��E5A�u�u[z��J)�������xY�X�ҭ��	N�v�����}�2dS���ڦ�>������8��B�z���:���SB}�SaH�a�}�>�'U��ܼ�w���QYs4�_x5L~ϣ�cr>���e}H|��1��*Q��=�a�j�o"��D�v���Y@eo�t
a��r�v�����Zb�],���䧝`�4q��� ޢV8�g#�ٳ=г�[.�e63����0��ze�ЖKQҬj��,���%��#���o^
	"1�E���eKv�}���� -�8�󯁷��:��֍�[,BQ�7��7�DXΈ��U ��w_F�i�QzXc�$iA������끸/���8�|�_8����kbۓx���ċ��M�����B����'�)c��/�G�-�,�����oF����fv1O&l��w���q�+ٹ:����D��kg�t�1��x��r[T�9�;'�4��
���P�j��Zjo�����]<�rْ�˺
��]�L�<C����vyЃ4s�a��Wh�{�5<Ɏ��{�M6d��=�%=2]Z�C�3�S�M¢^q\MH�M
á4��i�ذȁ)�[�	fi�c��LYX����Y7-���g_(wDK+�cjz�Ş6-AX\�	���a-�g�I�3kz~����Lvg�	`y]M��q�J��
�.>�4���=p���+�7�_c&qb�B�1�v�s����Ns��}��or�� �X�&���dշSL��2��X��	B�bf>��9xTS5�KT���e7�Y[W�;3D����6��jQN4C
)�Y�Ϳ)���`�l��KVOK*�0�4���Y0w�v]1�C-�i��a���x%	�hKhB����{6�0j������L�-O�J���w�eMmŏ�
��\��F!��K�Sb���뚃btpr��T9Z9�(ń/W	���XJ��Վ�4b�#\-���C��|�)���!�r�H\jڞ4>%.3ٚ�,E��S[Vi,�E�К:!	��w]M�!�e�H�Ss���>Y]��Y7\)vT���=�run��y���9���@(C��`���q���[��+�]t�Y-5�>�wV�;�Bh���
���@��a� d1:��Kuz	�)�f	h�s�ЬZ��К���:�n�f�f�`�(J��e��k�K�q�5����<�)_�-�25�o�+�	L��W�L1�\��]/�$�ϻ}�-"�J߮'o�a���B�Td�}$dt����[�}�� ����d�v�sk��v�%>=t.�z`�%>[%�J�,pO���&��,�" 7���Cꏪ
��,npQ�H�͇�o�Fox�hf�R�����K��e/T;��gq����|\��f��TӪ��u,.]nIs'�&9��=5U�[k5�8]�֨j�mNM13�j�3jmdGe�+�<]�sb�˵\�-��]��H������}-��>���Y:��(� i�	#n�T1��Q;7/Z�j]!�Fb��آ>�L8�,w#�KF��ג܄�\!�Y��Q	#�3�N�)��E�l��Y6+���5�>�ma�ǘ�D�1Y�-�H��=�9\2�%��0Uc��t�ܫg��'��T*�&J0�N������i�u���y���W�]w\}}S�u�4��b�fH
(2[�D�<�2|�܉�����Q�ѵ��T��E�u��������l���fɃ��yΈ��L�B�jk���#3mM���MA�69��6��a���k��R����f�ƨ�}�&�qn.���v�t���d�P�F�Z���sP^�Ov��F�2��
8Un�b�*���71�VUi����+D�-nȵR���N�_Ny�\y}և�s�g��"�A��BM�c�D{y�n�%��q�Vʀ�ƗW�:d�9L�z�Bf~Y�ϰ�7=�I��Z���1���Q��N�`1��	ZZ[ѝ8�#���-�Ӧ�Z��ȢjD(�\�gK�z��Oʜ��D��Y�Sy�`��k�t�����ڏ���=t9t��r������X�fPzg�	��g0�q�]�j��W ��*�o�2'�)v!�J��ת����Z\��{�6+�[�����oc Ż����w�+��Jr.B�w�סt���F��tL�8�?"�Ԫ_W%����Z����M��)�l���dy뼲�K��a��ñrQ�#�%T`H)1�<[T�ƣK{���6�U�s��ý6���m�ڮ�e�,b��hq���y#�hvu�������
�޽��0���Q@>��Sqj���e�+g_B�Z2Ҍ|Y��/��#��r��&�漼�ٝ�U��*p ��
�&~��-�`:�F�ٯsܧ�:�!�F��V�Y�dL���ﾃ_C����a�<�t9p�C�<�^��ox�y	kZ!�Wl�(�sF�܍���;�uxSD-�,!������!zt���:lg��|h\Ec���c��"]�7����1�.QzL��2CO�� �H�|\奭����dy�d��A�Ƕ��I
����m����֧B��Bu��j�C�wB���,��2uU���.#�PE�kа�#"
yv��`�W��B��1��-�ݔ��Y7)�D,|��=V��`�d�4o�7��/���3t�������3���{q�Q���Ž�]A����Ï 'M�ȑ��YQ���2�3)E���-]�4YJ�X%�9NW]t�R��hp�6��S�T�Ϋ]��
�5EŹ�{7����1�MQj����Q�A�bޓYʌ������nE�X��>˾��wWl��PRKu�I.�U��V���C��6�!Æc[�w�)*����8�W�)�fiC_fWh�zڏ����%��ý#���O7y��˳%�ޔÑdh.9kM�4S�[��wl��[�k�������2���sF��ohI�9ZP�Q�\e���������]\t�w���q6*�Se�iWQQ����ħn��rQ��ک�v,!]�.�Xw��cH^�q�(�k�3L:Ѷ.�q���+s��VP�W���b���t�n��.��[3r�lj��楶r�i�Jޙ32&-^͒V��23�OW"����*e�Zwk��������&�"��ג��cAF�\B�Np�$K�f����n�oa�U�W��=��weJ�ɎP�ŭ�޼�kd�(-�fI+�$�ӥp���"]�����7�O_ mR���[�����gI�I��J�|mmn*f��ZD3�QY�if��b�@1K��C;-���t�o�<եq�Uxf�	���X��������
�4WM�0�2�T�l<]���ҍ���S����5�*�7$5�(Iw�;�ф�RҦ��[n�f�8�{�P�%��8�i�L� (ǻ]��oV^Aٯ^�J#ǚ�����lf���5qSJW:72�Z������Qb��������CS��T姒sA:}K�������FK�n�-n ��[D���Y!&��}�O:�ƪ��-�h]\Q�b����d���{V�X�y��F��R��f;򪼀em%�|�]�`=%�V�K�R&�B%�XK4�m��ҁ������C%e♏,X��hK֎����EX����5^ҫ�Zơp�o���ͧk`%�աZˤ���z��b�L�Mݖƅ�g��<��e�
�l�,>�K�XTzK1�M
��uns;���5X)�ڌ�k���}�)4/fґr��2;w�RZ��-�Ob����G-�g�[����.cY�i�Eෛ��(����GDطzjgP.�ɗI1W֞�A�N��AZ�6�Y����1󒰛�@V�Ǝ�!����ә9�7Zv�)�G��R�m�[���L:��z�x`眮.�F]� 2s�ˡօ�B���A�9���û@Ww7�lICw93C�8A�Q���V�-�W��7F��IM��'Qƍj�AIٕ� �\�<M�xq�!k�1��\z�b�T{��[���SpTU���'׆��մL�x���_\mܘM-Wr�i�������P��B����	�mwk.:�Tؽ��1ՁdWtC��J��D�
�Kl��z 4�cb�-Ѹo2sW[PkӀ��o��W����dʛ��i̹�uc��? h�"�;�u�%t�ú������G9nw:;��$wRN��7]ۻ�4���˧'q]�҆s]�:u����ts�q�gWw.�\�'qsr���\:;�s�.���r��&E7r��.�ws����ww"��s����D������
9��wuw:���5��2&m���(�w[���@G*��ەJ��\��c�2\�Es���)!�M5¹�ۈ`
2F ���v����wk�':N녌60P�������7r�X�I�ܗG��6�n\r]�E�û���\�GJ��&]r�r�v�9w۔���K�w;A����ɠ�)%&r�.٧wD@�;�]9�wX��L˛�sq3F+���t��\v4>$ M�G45Y����2�����޴�s-U���rQC3&�pK[V�����'Q���'%�6����c�&�<v�u5�q�٨���T8g�v�]e4n*e�:sڥ�s���:��I���sS������Oˬy��뫝&���9'@�͂��t<�ʮ2J��p�yo���u4�?��`�����d �d��{�x�Nh��4M���,\�<�rq�E���Zk�O;�k'b��������uQ&�
\.���r-Tf�F*3��M�Yd���� �%���f�V�
�Bd/5��f_���jz��"_i��'-I�s�y(�4���X�ےN�� dy�nC;#+zqي�g&R�^�m�X+�nԻm2	M���s,���G:��h�켑�N�@�Gu��h�ȗV ���WCl��:�=2��C�cPu���@u�U�H�Xe���썷�TU)�����H�ԟ����c�e��V5�+���N�`�!�;�L�щ��Y7��NAt0N�AzH�ĸ���`�X�Fp:_ō��Q|�J�"������b���zr�
(2}:��n�����Q�!�����#V�y���1D]�
�}�fM���؝ݵ�{��z�U�����R�m�S}�m����U�C����� eƚ8lnKK��;3m�Z���J�baQ�H�Jt{`��rխ,W+C��Q��m�sk�������ݗd�J��&�25*��5Fv���֭m�c�f��z���+d!L��'-L��=cA�1�mV�r�fsP�N��=edW_��,�xnY����X����%�wBS:)�p��x�R\F�2�s�ڭG%nc�,2B��*���b�����̆��Ւ��.��5�ўR��*�
�z_�G&�El͜�k*��������U�ql-��tΗ�`��=�}Y7-���gz�C� rmaq�T�X�����Y�R�Y5��#�%�t>���m��>'�wK��u���4	��X�}�e��[�y�`�QA�%�ï����̄�4'BnX��C=�~�h5�`�|�mV{#D��QU=љ��� �.�ܳ����#�'�Q�m2Q/y^lS�}sPlN��An�g+G9�Y�//�/g�̜�7��_jy��<�8�B�Cz���5�h������R��F
��<�50��!?T+�V�3=��\j�+�ݑq�SsЏ:�S:����c�1��^�m.���9�5�"���� �E��my�p����tUkE�W^Y,��'�^9x��^�_���ק7�y��d�%0�}��8V�qK��R��^�Z\��re��&p[WrԊe;�2��$�wX[�Vl��R�Z6r9�,�-Y�+S���'�Ԫv�rﱁ>��{V�!)u����GA�L���bǃ����$[�J�ش��w��?\@6O��,z�X�P�*e��e����7V&����uFdu�!Vk��&��;�?���\>��]�`�����J�͎����~!s-W:�}�{���0����׷�K��ZE��jX���LñrY�P@J��}�HYv�o���D_mg�F�(R~œ�����Z��O=y)��(�U�c�T(c�C5���0
d1_Mo?�ur����I��r����}�F����m��?}H�Ht�%�*��˻���k�f�(��9�����~�tb!.�����2i�e�\V{{e>IF�TΡ;�-� �T���n{�U�Ɏ������n�	��M<1�x�EF��+٧�Nr�eL�L�˼�2`9-�Gd�ì"IY �þ*d"I"�Kp�u�X~�ܸ�X���ަ�̚J!m��1�uS��Bk2�jkK�gU�Ј�9�^%7"p+��Ǟ�v��[��b�c�t�1c�f�V�Vz_��-oB~�VLۧ�])��C�=x�\l�Z�y~�&EX�.�6�V-��7dԻ���Q1x@<8�RA�q'�G.��`�,G�X"͑��R�<����'���Eٽ�v�+d��{nME�\���:V"�H�qT�jVdRƭ\��(M�n�y{͐�-XB�[q�t�lR=�ˣ�v�܀.qW;A���P����]S&�jf�h*-��5�w��Ҟ�!M�6�F�ڌ=X�ő�-sP^�Ů]3���b�V�6WeVro�A�#&p�T�����LK[�/ʥ7&\�=����Wh�]��4�Q�ڒl��^�!@�5�ؕB�م���u�}��~��C�V�C83�ߥ;��V-��M�-z;%�)�\�ǫo-(�2�uN?KA+K��3_(��X�ڪ\>��K�d��(p���lr	�],�����e�$��X�K㔔�w ��,k����3Jl�1H@Mq.g̷�>=6&Q�t��d�Ye3H7K<��4 �2��K>�<�`r��|-W�i#��ff]0�L%X��SoLڮ�[�_�HN��N�ع,��R�c�OE�v���������|.� ��P�3�5�[u�-�wTV��J1�h���`�.���bq]u��^t�V0�w|��䉈�끿��۰F�o��ۆ����x��9">ow�|1^Vo|�����N;�(�@��p|��~�M��}�c4Qģi�]�i��Wr��V�N��},N��9lx�i�}΄8�'�nڬ7����:�k��	�-�{%���7
�7��d����'�����qQGs���K���U%d��@�s����y�����_v�Bn�]w�p!��Z�݆�M�
3e�p^t��ʈȊ��ͼ��B��p:9�?&k �9�HA���30��X=񡵎��r��p�;�T��9���~x~e��}�fHi��R��g�L�!���U3h�1�7e�T�����|!4@Wu��6��9�h�)�O��O�SWz|�!��C�e"��j�x{�p\Ca@l�h}�j���褸�q��zsԥ��o۲�k&�=2腂��:�֦�`J��W|�ܭ��f�W�}2�!���N�3�t���n4V�h'���欞��IT�׸ga�z9�����E�"ar럠IXS�>Aз�$� j�̸�;����e7�}�m�I;�I]# M据]-��/Fؚ&�[Q.X�z�'g�Tyh=��+f�t�>�T���qWs?X�]h��?���W��=-Tf��Q����ş�J̱��`�ݛ�p�Y:��O=�:?W�C��
%���Bp�I�s�%��u�kX!vT�A�zs�|S���u�}K$������ęr�Q�6cv��i�%6��LWXC��2SΰW�}Me<t_C�7}�NK��ӑ��y�7I���G#�+�.g5�ۭ辜�ܮ�7��U�w�cdNG��R��^��D}.�
e�"	\�8��E�WF�^�u��nTB�P���tu�w�*#w�>�e^��2*�����&	�7t�*3ɷ.�Y��V|n��ɕ�q�w��`��%��|��X��]q�e�`��e���Ŝﾬ9D/�_ʫ���� �擄&u�1Ų��������tЎF~��c*g$ծ�03�E��jK���x)��F�C���!�\���g!�h'�+�.��D9X��2u�
�WdM���9,��Nd�P�a���"d���s�12S��g}��k�	Y�w�|>���}��ߚ���[!
dM�:�kg���\q�䶮l	��c�����-���s�~��]7�S�l]%�Ϲl�y���E;����ː{>�0��Q��򿦹���&י�~�"�d]�a!s�̖�ݫ%=%�0%��;�-�S�{/se��QD�����mVd�_1�[R��V���alWպn�_�ԥ�ά�\��|V&o�������]�9��!;�	l��d��帽�ˎ�
4rXV6t;�e|6T�'N�����>m�֝�]���P'���TҰԒh�:�L����	け~Ѕ��%�6t;����c��*���i�n�T��W]��n�x&�rX���n�87�ǩ9�����#7�Yg�jJ�ղ�(ZV�V�G/wh��_V���� kS:l���3�qi�|m��=� �X�p�1D�b�L��څ��/���'hm�
��eN9���	mWC������M��O���F|V}�X��﯑���T�Y;�ÿ�[���:md���}����8m���ei~�k��v���ȯ��{=N��9�.5mOp�)��f��p���x�f�P�L���t|&D.����Ss�*9��)�t����4nvg��ݘ �uyP]KI�f!!a�`�}y�p�����
�z�t���OE��b1��͜Y� �ٖTv�}��
�%#�$��e�>��wS-��-]n"��O��S@�t����v�W���g��t�z��W��2�P@�Q��R�3p:[,}?%U59�?�2�9��,��;!9��B�{zՊ{E�%'O_�����T�;�,҂U� ]w��tNq�U�sa�Ofi�{�����b�|tWG?x+�O��0	ejX�E�fK5�
�ؘ���n�۪�]�>|%�;��g�Ƚ^�]�XF��t߼�S i���w�������B�͍����y���S�p_4K0����Li�5�-�O�p��m�D��\/�g��ǀ?��)Q�K2�"E��{Ɔ*{�����,J�49�
����}a@�e�Iy`�����@_%��ÝY���×AlK��7٥b�\"�j���3u����t���B�&��r9N>*�̧�n;9�Yu�sc�ev .�6�̏�J�R������[�)��0?�^�n�,����>�e��=�}��Y#:xY"�iS�Q����6h��v�I{Z��!��!��=5%����+N��}�������Z��W���(�(�Z�岷���LQ���L�܌u@ȶ���z-�/qoЛ3둨n@Ͼ_wˤ�������Ogu0��f�=.����|���Q.6Z����MA�,�8���1���үf�gP�����~F�S�%΃����~w��u_^�m(�:�D��ő�ݴ��9r��U�yw�Uӭ�v����XT!��e1Q.�_Ĭ�L^Zݑj�7'"�F��oF�6�d����K/��=�5?s�ݹ)�צ�ɓ��>'�@9���0�:�M��~�{P����ΚvG\�����A+dm&�-�4����W:�Ն���OA:���h%iih·ae�C=v�0�sJ�1����\���ls�E��	ቫ�q��3�k��F�ܐx��,m���f퍦�TX:���ؽ������x�4j�s,��S�ױ2�{�Y�K%��+����4k�ؾ۠�$�'l��$�>u�Q�D猡\��z�j����@de�B�~�V�s��V����j�f�"J�j������`���˻fV�����|�^��2��+[�+V�����xVG�@����:�Q�L��3Q��.��I�*�2���.���7�e�]��@vH_9���?]}�p.(��j�\6������\؞����BT򻮏Rğ�g흨/�Ԉ��B�F#��o�עo��b�ֽP�e�Q��E(͙wX(j���5y֣*8�"���GUp�s%M" nk��"b[��KG�؀�5�LgC[d��2
��znˮ��m�`)�L��MŸ�IN;�4��Ih������_҅e*h��E�k$b�����G���w0��?E�˭I�d����W�E;Ǹ� ��0�%��:�{�B��wԞ��+^�����:;�(.��̐˹@#R)�x��u�(����CzH/���ŷ���~��Ep��{�>�_u�Ȋ�O�绩��홷�n�3>�P��S��f�V����i5��v<DNeY]Qe�Z�n�9����B��we><�M�uī�P��SN0�q4��-r��U�1�"��ζj�
�������h�Z'�OX)�O!5�ҟ�*��6z�xK��=Y���)�,�%0�'�j�vMR�S��"�6�-�Z	���y�}�S�EICm��?��
�;�v)���JƼ�q�AJ�4:VNw>SC�D����>�06�{�0˾��rj�&Z�2�5�AZ.*�gea�t��&�_X�[%�JM�h֢�tx9FV�&�r�Ruu]����1,�)1.�[�c��\�Ⓑ/	;��ٸ?�CR�k�mS�&��6�,O=C��\T�GD���yF��&�N]�G4�F.|⸜w�g�)Ķ�����W�;e�g�=�YدKg�=΍�M[��%F�Β�(��x&��t:�(��{P�<�e�L�rP�]mX=�Pto9�uIߩVm_�v�����&��12��+D�d��hݩv�t������@~�d��`7�y�E���2�ވ��z�\�4�]�`���M0���?��Ke*�{Qu�;�]��ST�Wg+w�M������#��d�R �I������ucQ�S�\MM<�ٗ��ݓ��v̻�a0�\7 (^���/s��3NdT �?I�n���,g�j����s	��HMݐ�)���
�WP�)c��!� �^�-�,��xd�2�1�n��=��z�ጂu̳d=�.�O�H���3"m��C[<3t�1��#�zmt�
]�yk��n��.��Tv�Z��P�5����8���x����;.�3{��7����f���mm���m�[o���V�ݭ��m��ڵ���m�km��m�km��խ��նխ����խ���m�[o���V��+m�[n��V�ߕm�km�J�j���+m�[o�V�V������m��ڵ����ڵ��V�V���1AY&SY�'N٠ـ`P��3'� bH��UD%J�"T(�B��P*�"�4��EJI*�I"�R��R�(�k@�P���UH E
RTJQR�J}��*�J������D�M+m�t݆�� �{��%�U�QI Uz2��U�m�T����d�*R�]�v�j�-����2�JE�jD�HEl4�ur�a��#-%&�R����lФ
��k!dkUA$�+�ԉ�6T١�IHQ	U^��n
�B�j_   �M[m�аa�)����W��]��Ԯ�������<�  G0��Y"��Y�p@��iZ1c��풢�J����	���{�  u�UASh�A@�D�[f��0r���X�R��Ѣ�:( � �N��   �� @  ;����F�h��0� 
(�-�Ա�Qk)UP��x  ���=-uUmh���R4-4�UQ�qGKZҍ��2�R��}��@*��8k40-W���+��U
��i�^f��-���  �j�Q�UT@�����j�&�gntm���3TkUCk������ݴ��[���N�J�v�p��-,��QҴ�w���[SP*��6��D���  ���i�>��`.�����_\��:�������î��.Ύ3)�v��;�a��7gUz���k[j���'v�(k2Fm��mz�٪���T�RT���  w�=+v�� �z�o`vچu@.�i��Z�h,��5ڶ��Z����훻�Y��-��cP��)��#�l��kY�2�v���Y��e-�m�6�
�  ����g]-Ia�Jk�������v�>�� ���6�:]`;ד�=�����z�:V�Cj6��CB�[HmGk`Uv��t�Z�m!�E�h����٤�kQ�   �}�m���/��-Tk�]a�nYJ���=ڸ�WgH[mP5Bǧ�Ht���� ]�hm+�v�W�S�
�3
��[V�	scmE-���4�*O�  =�;5�J�1�2�V��ln����Q�N��+*k�+]�`������[���0����C�XUR�%e[�T�i��kJ�$�����W�   m{C"�:u�������2����T`�-i�*te '��̘���N�F�����Xkn��V�ӫ�z�GB�w4: ���T��̪RP Oh�JRP# #S�OM5UP#  E?�Ddb0T���*�h&F@	4�<�UME ��~���������4/�˻v����6؏�W������?o9��g�k[������$��BH@�bB		�H@�rB��@�$�H@$$>��9��_���>α�q�#�ҷ*���T7U��RAK�6&����Q80lK4�4lu����V�n���u&���C��	i�V��j�KK4��+�p@�҅�f撌Ԥ�Ʊ� ����ÎY{�䛻'o)�Ӷi�0����s3p<4d����,+�)݇b��
$�d%�z�f��0?�T�� [IYYO4[Uͭ���'bLXr���I�Cnc1!�^�u�`a�`A����PBe�(��ڻmGR����4�^��UYf��M1��Iu����^n�D00�Jaj࠲c`2��8lA�r9EɊ�ʱj(�43s w�'�}�;�LJV�Uc�����

2 4i|P����54h{�&r�5v�����JE�r�,�2�!��ؒ^뼫���%�ZڣG&�gee���.η��Ah%��)�孶��i,84RƩ���He
��e��Jf&�Gn��;2��6�ʹ-���ǎ�)陯6��HRx�̡��ق�ª�X�������c+`�p��5��)�l���z�ӡ��z��&�`K�HY�M�K
lMe ��!�h��oƭ�t���H4��4��Uu�����i
�B�!k(#A�Nh	of�zjB�U⩦�2ŕ{H�BFſ�V�f�SYi40.�c��w`�[�r��e�o�eT�]�t��4\y���h�H	J�ŧ{�(F���H�Z�����"Zf����݊��Z'@#T�Xe��/4m�.<���r�]��\�M�uR��V����Z0Y3@���*�iat�w/!���Hʰ��V&uB��@Փ,���n�w��Q�`mj�1Г3C77q��S���ڠ \ח*b�7Y���%���T�h,�]2��t�;u��x�T"T[�0�/u� *튇0e�l�f0�d��c6��phVu"��ci
"��77%��(�:1M����� -֛��V����,]-�r�h���6��{JkM܊5J:���
 :�f�I�Q��Ƀh��E�9�]3{�q���V�-e ��`l��O��:���ݭ�*���K_Q?mI�K[E���.ʶ8�8��t����)�nL
�sj,|�|��Y�>��nI�܌�Y{-�7t�;6Z�!�4�Z�h�6�M��u���P��S�cR� �f�� ���Z�(j��c�,��5�u&L{	3L{Y�[t���CvMZ�򶱂q��˓-�lbW�*�k~s�B���Z,�s��VV���Cr$���10en��ൡ F��	�;��

XA5y��p��b6$�����Z^\��q��+eb���SC�E2x���'�ٔ,�0�4����3�Y���wAKm�uo)�.��jV68_��M�I�Czor�܁��Ճfk˥qn�nm������L��.�ꖨ��p�:iR5��^�b�Wt�#��=�7��O�/�tU��2fd��0�b��Z�\��'TK�j�X��Y�R�7I�g /NؙFn�iٸ6��"��(ު�0Z!�9kS�L@!�[Ր6��t��kNB(�!Ʒ7oBAǬo����w�~��p��Jy�Wh��J�on����J���6;+(�Y-����hQpڐ���PSq\�"��Y�Z
n�0�
�L����Jڰ��&@��i������̡�*�	�f���vR��Ɉ�)��=�Jn�� i��fM9w2^�r����v�EB��f�Jr�c����b�BcvS�b�ԫu[:N������&hӛ���;��n
�˒�2]�r95�x���0�ف���r%�h�I����[���S���ĥZ2�dV�3;A-��.�#c�b�V�`L�x�D�w����1Pl8�*;Vl;hZ$m�B�d���kR{Oh�y@MR�j����hq���n���.)�UV�4w7KHY�<�:�xJ�E2��ѵ*}4V�i�F�K�/��i��F��h
owU�
����j�/%My7o��Kph�i+��NЭ�Im-��p�t��zՊQ]҉5�R�M
�V�v�"_Ǝ�rƵWtȼv�c����n�t�4�V٤����(���
�V��2%�����T�zt:v���;�Ad��
P6��wt��1֙#6:Cs1#��W4�Ĵ2�	H�Q�h��B�%[��S��".V��ydX ��Xy�X����(V"�jG3�-�a�)̖��3Q���2Y�[I,�l�(e��5���X*���d�6*���#�������nK��S�V]^���-��z���R�,.��;B�Y�����V���[�ֽ�T�]M�jJ_L@���y�
�F�4rØ�Rm,��t�Ҩ/]�˴'�����١�;OR����PV� ��gl�n��Son%Y�={.�5�m�LqS���+��a+n]�HnS��������z�*�H��9.�vZ{����'(�B��B�������X��GDv�l��E��$}�j�+����Ň4�x����1���k6�K���Y�k&�=�q�iee]�Y6,$72�(5%U�q��0�u���,Z��N]�eH���0���^j�g)팬4�%��5�PG�(�\�,8CF��U�
ų^�`�1�j����x��%��AR�H�ib�©�W�V���F�YATEַ�ZT���#�����Ɂ
֙k0e
�����ł+J��Y�[(��ަ�+	��Z1��4��e	��w�3�5�(�P��l�֖�b5I�2��58�D�"�L���wa
b�XT�b%Ā-Ѥ��@0��j��[__׌�z���Wt��ɵ&R�LrL�Ӌw2��cq%�b�Rp����]	��7`3�.�'�F�sU+���j���#����@L�Âj�i��ܼ{+\��߁�vdW%:x.k�)�Ҝ���MY@��Kl]�J�W�.���:rP��T�I�VEXeJ���uq&��{�&�C�.�@�ȍ�F�h��dCXE��WT�vګz� =���D�!�55����U�	�B�l0��I��u�z�Jw+)��~�,�F7�%��̧���A]�̢k2'nj��6��8�(F�^�������F���<�I��ҭ�7L�e�5���,&in����b�)�)�%���۳w�
�P}#.���l���w �E0!17�P�:3]kY�A�֩%)0f9҅�e��� h�v����6�aR+)h���p͗�f�C�Y��L��K��]�n���ž�r��,HR���k���[��FY�^���4����~r��z�S`�p	 r�YJ���PݰFVՀ��Ys
��b�+��ec�Q�����t���I���r�ǂ��"��a��5���z��RT���̫I��cri�=����b�%��QD�b,�jVQܣV���&ɇeKZ�*��jՑv�ۗ��e��gЭk5{Nӗ���n����������n7D����k#	\T�;�{��)� ��n�Đ���k -�`���A��,r*E Z�%&�L�[t�����T�	��
��OF*�N����������={��FᙐXL�Q��(T eK�Jv���t���J�I2�e-Ë��Hc��J��]7��Sr��Щ��Y{aU�V�Ү?��EзW�@���v�V�	;"���0Ę��U�Ե�SUM���t0�J7kL�{o��47pG(X2�R���18H[Zr&��Af�q_�Tuch˕Z��-D46؞��2�j��R�Z5p��$R�M�'�J�U����wzp�$dM�Z���ʎAwB%�6[{��oV2Y5��7XHWC6�m�#$W*�JJ��a3L��䡔��h,�3 �(�!GM,*7�Dq����ƶ��u���J�i0E���<��M��,�J��N����{P�[h䩔y%�d��5\��n�3]�I�A
�b�jh��<�/!�l����;a�eF�J5��]�	���9=�(.7�d�Y>�[��׺082����iMrV�6��)^ �Żt�� R@����Ϧ�n|j���$�3	6@OA9C5�W�釤P�%�6P'-bN[�a�&���j��ޫ��*��b�6�����,":[z��]ೡIq�R��9�h*�ki�W���f7N��Ϛ���P^l�j�.��A�#+s2�&�����@�Z��Ԙ�Vĝ�u�e�5�s��$[���C��U`%�(i{&�f�ѓ��t3+�i*�
��������:��3h�XlP|.��x �zpf#��4��aDh��l+���r�E�73b:��Z	ЪM�`�r�&K�Sr֢����Md�]�D�6�JygRz�m����+*�Ց��cu*�AZ�"���n��%`�f��cn�m; X�����jA����Ov}v4!��ɬ���b���[��r��,��4bv�4T�&6�Fn���j����v���r

*^�;@d̵�������*i�zNY��f�.��.��8������f=�F-�x�[���W�(fYn0ɰ0f�i���0U�yhk���˺{h
"-8���e�l:u�w6��5�{yWa�-�LTز���Z�xk*�ZN�qE�X]i�[Ys����2���C��6\�Y0�S7Y[�h�����ӵ�Q�yIz���+J�3H.+��wB��N�5u�a��Sy�;�3�`�{���6i��eJ�r u,w��4[	�5c�w$�ص9�7���'�Z�6�&"�wUb�$l���X)e�����c�Lr춱n��ĺr����K
���N��X��lv��L5Y�vZ���4)��4�QZ@��|�fG.Rq؏1��E�ų�K*,T�fT�� ���i�thJ��m��*��*Ҥ��xܺ��Kk7̶�ݸwFU����ˣ�)��4L�o*:��Z���gSġD�C7 �2��F��ʙM��^dݷr��e�Qƚ��1���v<ԡ�eĹ��.ޱ0TyBTZِ":i9Z�k��@ڳ����֕m�b���l;�բ�)�)�����%�t[�9yJ�?]�YvԊi�����v۔(J*;�CUF4�Ս�7
5s4ܒj�5�Y{���[2�
N�1m�iW�;�n��u���YZ��m$3A���Y�Ԓ�J�t[Lb����k^�kr9��ҡ��T�%{0c��U%��u��[��.�;��(���խ�j0õr�׺lT[S�kU��)S6N����
�41�8Z��N�QԲ�8o2ނ�K�tSVM5P����t�{�Cʒ��Kg6���(�!��l��&%�i��e�������vt�肵SL���Z�����*�eC��n^��q��i�aL�zUf�KF-����w����:)��+ԥWR��(`+@j������J�znJʂ���Ĭ�ј7*n�$�)D��V�#L��5��62�8!2�UhĴ�p�3�vYʣ���2��vd�����l2��0<��*2ƻ�ĪjC(�uA.��Ph�G"&d9Q�rSMb%V`A�Æ�ʼT�E��p��HbygR�V����h;�lRj4�s��*a�7�2���eF�u]�{�V��Ļ��l�ȭ+*��t��W,J�B��͠���j��Vț�T�°
N,����o!�Wۙ��U&b��%�˲�ę��n��-��F��DW�*;�K.U��T� b5�HPa��X��X-�K��HȶJՍ2"�wf�ѻ��-gl�nE%
!ѫy��ӎr��f�[�*ݼ-є7v��/zsd��,˧0�>�2)gj\NEq�s
&������7��-{�-d�����Wz>q��QJ���(��
j��",�y�D�C�XUj5�ǯ�sUb�� h0&#t!q���ָ�.dL␜�Y��=eH(��i&�{NM��+Bf�^��]]��o	sv��#玸���_1i�c1�*JJ�=M���ɏK�=n�'v]�EU��7���fT�d�]Lz�n87@8������M�Ah�!�N�H��}��d�R����T&搖VDo.	x�1J[����wY5�I���pc�K܂ܠ�����ڹ�V�%��7�n1'��%;a���5��4��ʔ�����n�̛�ܬ)M4o5��씭�ȭ�1tF�W�2����inҗ2nֿ��(#��k^cD�4�Z31"�K����C��)f�ha�L�X�l3��-A%���KOs1��#	�c������t�EQV,��4i��c0�L[6h�M�c�O0#��@A�2��ٳ�Z��\c2�7��8��e��^`GL�5�+mj��������ܥblm�I4�yM�J��%!�Y{�*�M�cPB.�6�w#�uyvv�a*+I���:K�Q�{3E��e��{�Ʃ���%����ݬ(�HI��f5Sn��b��*4�Ak8�(��|��(2bg�]����`�`ZT$������|�U�Z�#L��Lᨎ���n�4���)�E"oP�Y�Zt;R{��K�76�QKhTK-�M(���Wa�Z�b�
��(��#5��-t�nA{X�b�\������>�F�R�֚8�ud�J9�lV�k9 [۷��ǲkץB_r���­�%R�g��18+^ӫ�ԛ�N�2R�N��,�A� �.�����4ɽ�r������2��r��)k����޻3��!���V��Њ@q���wE�kDF�^�V)<���*s��/hCe[�O;���~y��B^V���t�W�w�-��`�{Km��8��ʹ�m���XW.0u*ۜh�fhJ�{U� [Ƣ:��0���Gm$:�WB>_��P]�;�U�ں�g�9��mn��16��K�t���`!�u3.k���4fF�fµ �B<��Ff�M;
�]�|jf_,z��'wn\F=�A ��˶ ayϫ�4�4)��fbx��WQ��təA��pn�j7K8�<$W�d�yL�Ѧv$�T�sY�;5q����펳�c�]�]�i5����M#�]��V;����.�N��N�|�jഺ<MŒ��p��&���6]p�A�#��mu��P&g3o���X�.=���My9�(�`�Q Qօ��*��7�nMT��(U�Nm����^�U����ы�ؤx�TG.c)���J
M���_��YFm�t�v�qi�VEag�L��>�2��W�g$y�>w�I�t�,W�v:����PǴ먶����nVۚ����V��s��sU��Z�����L�L��Or��uj|�W{(i���l�P���x� r���U�Z/`o�+$�fڧEP�V�/i�U�]��u� ���}��%Nw��F�x��p6��j�~�"�����P�q�c�0�Ձ�[ӥf�Kb��ی*��L�r�w:#.}�v�|����k��ﺛv�ǓnEXQ�s�_��;��{֦��*w�����{�>O��F'}8�c�h�p�+���Wt°�	{9I��=�-\�|%%�%��oa,E�i�+!��N����	�t�@�R���*���\:�δ1s�V,-]��ߪ�/h-�	����u-��o),;2��Sf9�%��>��96l�� �����7ec���x��%a��u��b�s���A�>�����y��Ϙ�ɗQ_\�0�H��K�m��1r9!�WXZ�3�ֵ�����_k���cG���犛�#7�L�S �ޮɒ�>\d��,B��5�6|���%��;8�����a�;Kw�fudhQv���T��#�l01�/(PN�2���Fum�k99��{�Aҗ�wa�Ԝ�a�qAB��n�c:t���:�����]CQZ�[���y�7��9����{�b<�Kp�٦7�̑�"�A��3Xt>q:��bn�C�&�W�I���w]��ulS�:id�6�C3��f�o���O��)Z�K��Vu�����$Ev�KX�٧��Lwi���ǆc�
٢:�(�S���(	��F�:=��Ֆ�=�%ߦ�֔��y�:�p]oL���yl"{v��$��Ӫ��Һ�5��7������=�<{�x��s%���3oS��<�'/�>�
�V�ҚĠ�������Xˁ%(��Ɔ�E�/�!6_F���3ts-�窎 �T�kEu^L=ˣw�AI3�E�Ӛ�f$0�+xUc�[y�Y*��Z��g��ל�%H�U��D����k�	o>�&��Ԣ���e�ުiR�(��1�����Y����ۛj]>�9-��{-.�m=��U��ݑY���P���z0c.�'Wf�6�8r�Η��X����s���;x�{�vAX��F��s����]|��t�P��W����o>f�Y�%|����w\�Fzvw9�
��V�}T ݩv)�ݒqT��9�`N�Ӱ�/2�j�:�W,7Z�G�Hv!�S0c��Z30�N.�u�Ig�K��	��#�Oi��SEm0�XX#�:����t[ �v��p�h�`�A���E�3�6�#7��p���R��n�G�9�@�5��l��	���s��9{�`�IPӉ<�����xm�wږ�l��͗�鰷�՗�
݌K� �2�a�]Y�u%�>���a����A�;�����^�yڭ�7�Lmg��B��6��f�S�����aj� [�v{4j�f�f������+�N����'��os�nx���w��iC����[�4�ti��]��aj���ʇw��^9���A)Vy���KU!4���;e!JV۔�E�T��h7��HP��U�rԧV�z��)$�tA��wX�.\��|;�T�7�Ԛ��f�t�R�NfsD�ݡ��)ՙCa���x!�^��XS��w��>��~܍�L@���!em�v4}�]fҒ�"�Z܀�a(�r̦����9�cK��o����X�t�h��f`��h̠��&/�h��-����5}�DJ���u�*Yr��ck�R\&�k;/EH(Z���u�Ia��&m<��Z����n��[U�{b�{o;x�]*⠫7kr�?v���=2.P]�ŀlj`�{8��odj��r�-�j�i�5V����y}v�����A��,�kv�珪�Y�����W��Bʩ"�s��¶f��_D�5��К�[]��~�N����5Y�k�^K)2f�J�yJ���v�Uos;v��OKy��^˴F6�M�
��#+(M�]�s](�NK��{�.*XiΚ��#�CqM�[=t��:���l./b�5�L(NuyL�<�"���z�"&�'�z��\b�7�<#��A0���c9oVQ�V�9�I�]���1j,C�v�hZrc�n�'#�b��H霘ռ˜n:���Y3����3ᦕ�C�9y�aУ��g�	Z��Be���P݁Ŵ�������M�b&���V*v�C�76�\Q�[�a��Hĉ;9���3�]V�x0�ZV�D�.\�z/����cy(X�m�tf]�Rݕ��>c�2��cN�N���m�Wl�׉V��jB��̅����06qE�K"�s:��; �I[� ��]�0�}�w\J$!�]�����r���o�.��[}X�7���Y��7��՗�UM(,�p��;��Vl$�2�7[���oK�n��+q���P���嫻����Khk����_�^����8�K;h�"�	�.#�OueܠJnR`E��Up�;�c�oe��ww��lO��f�nVn�|��7;����h�2Ãj�U�2��N���ooF�&ؼ�{#X 3/"�X�j�s��pΰ�eѥl����hH���Y:G�*vE1[�k.��fr�ifA$u��g�t�g6�^ST�޳�_�;+��rn,*��\a��I���/�rQ��M�B�8p	y�&{M}!Λ�D��6Q�qR�!=�p͢���z2��� ��ҵ!�K��w�]O�+�n�ۇE�����t4�y�6�c�|��l�.s��,<��~��>O�T��w3�0]�	�p)�$2JX9w�ȍ�,���(j�����C;\���ӈNo�u4�rA�,��e���C�j���y�b�L�����1"հ��o]r�k���[kV���nʑ�z�/�@�R}}
�	{R��Gb�e��*c�n�oe�Q7Y%m̀(t�4��u`Q*r�Z�K�}�K��S����y��=�Yz3A�Z���Z�ٚZ,4�՘��!�=�'���J+;j-���RX^�m�x�}z@W
GA�g2��Y�A�losݩKZ}����g{��{��-;�"�T�.]�ۦyׄ8�f��C��Ԟ����WT������י�l��zs�:m8R���/C{�x)�����9f�..�M�/:L0U��]Y����v���\��**�i���.�N�g)�{����m�ۊ�̧7)l�\-����o(_,���z��<�	�֟���-�r5\���n�{�2���ӏ�xK���`��B�	��ҖY���ewK��A�"U���ۭ�OЯ|���QlN����ь�H�*d+쨩���3M4+��&�`f$#��؀�����,5zGdN��[�S̽�`ڒ�PArz �9�b������DY��Ζ5��ާΤͮ#-�P��y�����f*������ ���,6��"VԩVM��o!Y��v��X�R���8��NY|���2��f���4��Ԁ�s��Ҹԩz��1�B��e)6�Z��C�����鸧a�����^�ⴗ\�f�)����u��;x��դԗ�VcT�q�c�I�7;��1���7Ir�'�ե����H>^�\{Q��z�7��͍]im�����y"�%��;�ג�mcF�����m������>G� ZG:e�m����O_�$��w3�k���p�Y.-��s�Q���^W,z�fV��s�rv�o(V3q�$cM�+�4k�!��[jr;Kr��x"/��1�����^���;Bȷ{��Vn��K0gH:���ą�������#���M�����}ǊO���,���R��$�A7�z�4���Z�Z)�Bu<3���O�3%�b�jBH��������y.��.��]��eL�����I���VCyfJ�����׋�h/P��љ�Dv�x�;&�d�S�,cp.�q86 �(�y�v�U�d�9e�\j��Auր�i��K+�,�1�z�W�O�qs���i���v��\k[d�z��oP�RR��y�"ZD;&n�ת��}����B�o1�7�v���\N:�"4�P�t����՚eۇ���J��ݍ->�4I䳫B�I*�����1+�ƇAPogE�t�m�0�a$���B	��q�bG9.`�D�{�ӏ��)�U�Vu�ޜ�����O��o�IIn��ʓ8L.l�؎�;���/)�,�t�ͺ��	��7A�|���ۆ�5W�R�Wt��[�!�����m�a�[�wY���˔j⫧c�X�V�r�|�sxv�퉾Ė�����Y��D{�+z.��OyN�L�Dv���|��+��!�D��Ҋ��2�3�q����m���e�8�i�S(��� �vP7�o+����vVҼT-���d= 1Yg��٥[I�P�K�oJT�����#ً�J4�D�����Y��8�����*m���Փ�t���}��a��M��&0%��b&k�]^Y����s����_#ρ�|�]�`�Izlwe�ΠAr4̫�uxm��c��bĕ�F��0�^̓�YKn%��b�]sˤ�ma��6��ADo\2V[t�
��2��X�V&yrY���N;W����%�Vfw'guꝎ��be�d�7��TO^�[2��h����8����HOr�p�l�WgQ��t��f��:D���W���<h�I޳.�L"�K��֨��]*]!��y�B|�>�F����D�/:����$�!A��b�D[���p�����ӹi��+Z5�6����P��;���P�<J����J�Vs_P�KM��V�ˆc�y�w����e��js̢ʕ�2��}%"�]�&6h�յX�����u�k�[�ƴ��t�$U�:��MmJP=5K�(�ͼ�+b��KD� ��$�Ќ�K���U��F찿N���<@���yv�0` 㕝����&K~)�v���k�1Ot��6�Ԯ���;7� �o�p��w����U!4dd�]���ꁉRlti�ltbQ�T�;z�]c�w��V����7�4�gFK6)1�R��6�L
�:���y��\����\� ��@�rv{s���Rhׇ��EuK���
i�at4�O�UQ��U�t���f�]���2�d���0}��ګ3u�V��8�������2�U�w��Au�c���`��w�^٣Ͳu23��Sq���֮�J�,�����#zqBA���+�o銚VZ�����{[8�֦���j�Ukfl8���B++�]�Gg2cm��"�vݬ����|*W.��O)(o%._j޷-����Z:�z����1Cf�o�M={[��9��C/�Ε�8��!��p�|��ɷ�n����~�ϮQ�W��tT�:����}@Y( v�\���L�	:��c�ƛ��R���������ՔLC�T�Rp1wN���skeum����1͛�S9��N}����GTނ��ː~�Υ��=�s=|CK�,Ӷ��+�p�q����W��K��E%hxv��F"��V��wM���꽭�ݾ��[D$��RT�)�
�:�NҨ�Y�����it�h�<��j��;�:�n�V_i�H`n�i�:[Ὂ�.�A��E��M�&�f�l�ݛ/�v�X�T�w���=/P��Y��P\0)�|�
�.`;\�^�AU�7u��F��L�Np��|WMz�q�B�`�"6Ei+4�O�6�ܠN�,���ci�X�0����[�s��*�!�<��t�slrf�*D��av͒hy�������k`ƨY�y�F�FW|�W����6��&z���yq��W��gH�����Q��`�[�ǀb�w��`�)#Ʊ�f�}��v�x��A������� ��܍emJK�'���wBM���kw�o<B�4��n4ol�Sr�h��Ox�*����[;]w'�2�A��1 ���F��
�Yw�18�9#����1]+S�'҃�����U�8+߳�܎�������p=|3FC��(^��K2T5� �D�7{N�g`U��CiS���]Ǻ�X7n���O��l�V��6��|����o��-l;6��Wc�A�e�n�,.��o=�|�S�b����w.�k�6��M�:vwЗ�ޘ�(7t6�5�e��Xs�3|{8�e��c��ClM��������6�Ͷ:�o&�RAY XB�%>幷���t�����j�m�*ΎK�3�XェS�?��d}����C6�ڡ�>���w�廭vK�+�u�	�v��v�ͭ�/���V,s��_%�ԧuXNw��}�}U_|H ILaMf�zܜ��:q�����h�$�/qK�f	���v�,�\�9�c�J=����ͱ�xmU���ˎ7��f��31�y�Y=�հ��9�n�P�M�ZzwJ�v	��{��^X�qvFW{ ��df8��+@!���H��ݭÃ�x��$r����C�Fwt��SH�R�[A�ӗsX�\����D�y�9*�W����qSdD�*�Z�S�ܭ:)Z����:�$���ԉz>�5��"!MҸo�v����(j��З������c�W`���|���7]���OS�z�������r�A�V���_��8a5�֍泙/K�&C�B��aWL��:Th��ˮ����s%����PmX����[����f������>��5�YQ�*,���˽<�{�\�i��7�K���v��fG]5gy�����`ܒ &;'2����s�^o|��'��s0�t�cط#��!m�]�#D']ر�Y�쩗EDo(�C^jᨛ��ͩ}�k�om.ҷ�D��$ޚ�Ī�ɨ�-7�Rg�yi�[y�\�9����r��1&�]�Õ� ���1:<��	�zw������m��D)ە�BR��y+���PG�.e���L�tr�,4>�V�D�4�Fe�]&X��E�Su�e���س�!6�tM5ϔG2�fִ������=ݨm���f��eN�c�.A]���ܤ���v�C���N��"��ĺa-��+�TJ�:h�c3b�0�lw��M̵��ܡ�u�γ���Z�ҺQ�gvˤ
MX�Xw��)6�f�G��Յ�{v�J6��'t:�1�7~m)}Gxi�����v� �C��vj��n�Z��h��/s��yP�kK7�h�z��+���J�º�!K��ӧ'u.��=��v�t����Y�ʴ)[M���鎪A���F�o2���up�y��V��kU�{��;�Qc:���sz���S+*6:����-��Dve'JL�'>y#��Ƅx���ȳ}0FfN�n�B�ƅ��6��Z��V��.=+���;�a]k~�Ve-cq6��(I�X�Ç��{� ^ ��w�iPk7e��]υ�(��!�%JB�l*�<������WeԹ��X����\�O6M\�]��գ!�Hb�$,��� �w���y[��sXq��1��`�ժ��˨h�X�NŜ.uDSHc��pv�4��Z�N�����u��n�d�hLⴐla��Y
]�$A!`�>�h���C��ː�&d�_�+�H��IR��uJ�T-`W�m�Jc|�g`����z;��6�0<��Yr��f-�A<��*�o��\�
�-I!꘱���26 ��»f/�{K�)wSY�jtۡ���gq�0SǼ����ܻx�gcz�]�U0�SO<�_%���VHж�NI�6�Dl�-;�TTm�>�üЦʴ�wS���R����V���7�xy�`�}�oL��-j�Q��*����+iڇVf�fG}�!��B)m��m`���4i�Y͛�>Uy{kNV����,}�n�X����^� СL�~�]��$;w~�C������*;��^6-�j��6�r>��ўl�a]t�oz����9�`�"S�쪰��h�ާ����=��J�m�í^MF m��$�piVR�)}�r|&i8J�wrc@y��:%��.��[��a|�9S+���]�"����p���]n<q���/��%Yڎ-�`XZ�	��ͳ�oej�R��}Wcp���Xf�S�5z�n`M
���R&L&�y��-*�"����Ox���},+�j��L��Y��&lx�� �F^s��`��8w��{FR0n���U7��}WY'c#�b/bB�u^�|�T̹�`�dnp�el�{���(��
�;�|� U�̈́��R���6n��(	�^��А�7�;�^!�݅��]�^ē���[��s(�!i,��R�,�C{�Wf��:�Й�4��ؕe9�ou�i.[J�m�uux:���2P"]�w��C���:=K�F�*��e��]�S�#9�F�k�2���m�.������Xʜ�����4�)��/���z���rpҚ.�v#|��U��ə%N**��&/��E��x"��,m?��%�� �X�on���'N�Z�I�3X���,��cerBTT0�rֶ֬�z�t�t���ܭ���D�
�s\��_gt!�{xo��Z��k�,��X�d�㡽����v���ի�nAgY|$�qd��t� �F�������`K��7%���z#nu�ޘ Ɂ*�|1��F��Wٵ�Y1�f�^"+�e@[�����V�cᮻ��@�_�˛�7xf�]3�	2Vnu���pr��sW����%=����R+�F�{Y�u�6i-��p�R�=�uX��h�M����;ih��#]�Q?"��n洆��².�k����(���˨����`9d��\�t���Om�/{{9=�j��4���>[ܺ՝	mu��c��lNU�.��RC�^T��ޔ�С��u��z%t�n�96�ҭΩx��Oqޮ��a�Z�[%5�p"��n�Ɇ'Vmm�)��:����S�����q:۴�8�wn��vr��U��y�o��ήP	jE\���`���]�Vr�\y�/f���P>.!��������n�4��=��$�Co�;��xe���z��d��vҾ���3U;�+UC��ʟgF;m��-��˚F�^����SN��c�^���N��ĵ\��r����S%h���������ܤ���+az���U���t����z��Ӯ��< �vd�7����=8>)��8� �]��9ִ�U:^6*������m��{xb��	:ZI�@*��K\/>�;oJ��,Ez{vR�t0�ܟ'P���MQ���T���S���LW���ns[R`�b����i�7����I��V0y�W�m㽫K/�9��V��|�s�)Q������r��֛=���H��}w���qk/�jYY����Hi|[���,iP�1��ϑkD;���	��7�i��&5[y��f���
�92�$��΀1�p�\��(,���]yLt���R���{Oi�5s���*������b�����q�4���y;&Fu%]�օ_rڷ�������+E
���EϞa�( �m�hu��uLz�3.��#��}�L��h�va|��ƅT�#���v\I`~��o�����m��L}u��%"�Tk�e�
+y]��d�fU��뜝�o+OM�����^Mf��:���r)]�%l��݃Dd~��9q�rfw"6�]�A�_�ң->�T�u����O�#PM�W�a��	ȁ�Xr�+ګ�;1��|�
�l���t��)A��y�Sl�+���f;9-V�Uz�e\�8#ƅ�%�ʱLL�q��u��X'f���+���{���;��	\��m����q����yat��B�d��T�g�t���՗�wB�w�J��F^r5�VYv5B�J�2�������p�*�[Z�^�խ ��^�C�!�=���,+�t.����|t�[��|��)�a���ͩ��o$��aL�H+}�F�خ��3��Sx��1�UQ��S�E4{���h��w8Ӯ���w/����+���[��ꔣ`�#��#75��MA4 �:J�b��r�`q��ή���W�==�,�;'(��A�f�e������f��t4��W^*��9�~�`�C��i{���^Y��PC����tp�4��Yt�u]ӟjrѕ�<N\v��~ξ�s����5XsQZ��^����۹�3f�;�n�k���IN���EZ�oU��.E)�zCu����&���Y4_G��r��ʜ7���׍n(&h��D�z����������*���9+OP���o/m���q�K<��N�x�C_"���$fqқ�[�y��}�l�,��� �/��!G��[�����ܦ��`pnd���|��jhV:]�zՐ�����TU������]a�{���է���Uhvt��o��7�c�jY�(�Sr�ų�3+�d�)�W��m]�5tCC��۔��B����$�³�R�Oz���
�����n��ݹ�˓c��ݤȀ;��ה�;�kjѯiY���ιS�2c�q΍��b�v_+��t�{�	���gs���1 XU�s;-;�m»o`$�n�0JZw�������J���Y*)�璜|��=�G%N�������M�����~�|`=��+�o:NS�F���@i9u�n5�;�ݬm����Q��%��ؚM�����jF�c����ʷ~5��^v�@"�KW���Lo-f框���4�����`r.h� ^]�$���G5�
��r�71A	qU�j�u��N���uE���k��Ek79�%�#V��k՝̵���[�`&�u6U���q�wbc���
ۼ�B%]�������憕��TZ�+8�Ţl�P�GԻx��5�#�i�R��r�(`Iݑ:�駆�|��=kz�KW1�eiC��~�E�	c�s��gn�:��Z��K̾��pN������h�+�np�89��	���Ö�2@�k%u�p����-���4p��K/�XZ7f�iw�b�����O^���)�޶)��(�����!��*�$�7�1��z��2c�V�l-ˏq�]��y]
�{A��	���5���U����vk��A�iԻ�k�d�]5Ճ��(@��	v�n_46���w`��6����u&�.�	9���PT�\�b�ɲ��#;�,�<�j�cs�;J�կ	*�Ru�K��#)6�g<��+�+L��=X6&+A
���K�h��D4��qz7�!Fd�F�Ͳ���7�N[`�,���ܦ�^���M�+C��5m�ژ8��p^�Χה]e\47��e�S��ǔ�q������� 
�KC�5'�t�׆����>53W]޸	�%'5�gJ�Z\�:�}�7��N����7PKw�6�!�Clb�т��f�9���!#�e�d��j�1A�`|��D`vP|T������3E�$k�U�9q�{��9� �.�0vV�U��h��tkF#��ZV.ޥ+|c��J������<*Y����1�Ş�%\ľ6մj�.G��UF�.�sy�{6������Y2M዗7E�v!�멎�N���}��E���X�eP���uy�Q�t��姭�5��Z+�vA[~^؃嵎�`]q�\�+�X�G�1A%M�ꎯsʀ"���u�Ce`v���Y��ۄԳ�ƫQk�os�S��l5��s��Gx�g�V��-���dr�
���r4.��ONP�p�.�*�S����\X����oBcS.�z���V��D-��ӅUB"���d	��A��6�J�}����g<�U���V̥[�4'U�. 
��pX֣�֚��Y�Hk�e`�|�c�y�:��o��T�Y��e���}u3����ʺL=�hW��d�c���VV��� ��������t[�CxӖ�<}��l`�+^9�U���
Q��wxy-�B���3�PI]�z*{�;���5C1WD]%��r̚�z^mJq�MS��I-����]%����u2Y���=��+��V�,�7�f�[fr̅c�v���n��j��;�Z������h��2�{�l���������;�Sr�Z�{q\�C'"�]��Y6�6nM�{��H�*a�}���e���	�Q���/��c��N3�r@͸��ظ���ݷ5=YY$�}����Y_C��Q=6*�-�C�=��m����N��j݌�tr]��O.�R��E�����ʏ]k�ud!�� ��[维5�M��w�F
+�W}�
6iT����}x��Y�o��])Q����݆o^����F���t�U5I�T�[���P�ꖱ���˽hԂ�V�ɋD����q���H���
�]{(E����{p��v�,5��[����T��K�X�*5���;�$#�[k$4�!�Y����1v\��w���#���[\�:C#�%Ȝ�ڻcs �����&^[r�m�g4L�a�,�Ug`r�چV�Z�����	k��Χ���Lc�O�M	�/�;5�����^���ΑŽo����װ�j��r��]!��^��}sq��l�XM#��b�J�<f��
�kdM �;h�ƣ��єTk�ܝ(�Z� �Z��i�
�K!>1,L�+N��W�ne	����u��:����XW�U�"���}:鲭e`��
F�4����UiK�}�wغ���i!�r��37��]�ff�X��jKݱ5��r�C��� ���J�z��b���f�,չz���� nΥk�0�7{�Vv!r�V��r���B�vw��x�S�[�"���)i����V{j��ވ�Q�U���`f�U)�Ry���r�s�1���4�#�t%,���D����-�ǥ����V�%b��D����1����e֧j;J�u�+w�u����`�U�F�;�S2i�H�Y6Yh�DUY��f���/0���]�.��*y�h�ZÛ�­�*v͛\�a�{;U�X��Fy��Q޶+o�z��ڲG���7mK�Q\���6L��co�-���v�s�U�V���yW}�buՍ'(p��2h���F7:qnՑy�0g6iK.��s���Po! ��2�RL�>��P�Y}��*2;X���n�v!V���n�������ٚ����1+)���zo�X^�`�}�ϰ�V3a�G��ED�<����:Q�2��N�����Y�}���>��}�o����'�T;Y䨿}N�o��yz^�#oemd{T���.�Q����<^|��S� w�ϖ?t�������S2A��N�
��h�Lf`X �E�:*s�xI7+_M�V����/Q�0,�z�yB�U��"����D*��k�p�g��Ñ	Y��)t{']ћkl�^Ӯd�ܸ�M|;�ɏ{bfQ����ES߮	�6�K�yul��Fj؂��.u��fok�͍�����h9�ϯ2Qs���bbnZ�T/K9J�xWi�g"C�2��w�6R��s����K�2Qy��ހn�;��x�W]D��,�����E��csmE�ۦ���FU@��d��k�1v���Ӗ0溊�T��n.���n�R6��� ��:���Ю�]�n}hu*����6p��X[:��/��u�j�\u=Y#뷪�]&��X����&���6+6U�K+z=�����å�[�-�j+r�\�^�'Nj�R�g�yJ��a�_0v�ťbm�����G���"Ԯz��&O|5[ղ�ӹ;{	Z�{͡>�S2�q���KoS挡�
\�e7]�;�0S٧K�;���2����J�
�z[�dç��wL3�t:GNW7v�m�$Ŧ��ea����{�x@E�V����#]�0=��ү�%n�ﴘ)�mD�߲3�^���F���S�G^>�ܜ�H�2�iA�P�5�EQ���-
���1�+X+(����PAQ-�QTeD��jJ�b��iE��-��kh�22�QHũj�*����X�1�"�*���h��H����QH���b�UVZ%�%�b��ER�V20PU����Т�b,�QQJ����Qb5�*�,��KR؊-�T����mT���"�Ib��TZ���X"���T��,V��e��bR�Q��J��m�QEE����*"����1*Qb� �X��mEE��j�EEE"T�"��QUEF��Q��m�m�+l,[h��TED�V,UU����ł(����jUH�F�h ��+��mB�Tb	mX������iE��T���E���+��EH��PU���[QX+R���V*R�-(T���AQX�V)Yb""DQ2*��5�xo��}�s����������x�[�ӗU�a�KW�i�؁Hur{Z��K�֌ݽ2tuֳ�.���u���	���}(΍�xh�c��ܥ���t4Į��])V��3AVj 6���f�|$p�얳,�z�jm�Y�S�S˅�Tϸ(e�ʄKO<���f�%�.���'zX�y�m�ٝw�7p�2�m����.��]ёY�«�/�>G��fך����:z�Oj��l���,�-�oۈX{��D��/�,R�y"��+,~J`��ǽx�=~^�Ŀ��k!��	�,�_I=/�;��zX԰k��sJ�d~�l�����{����:u7d����"Ȳ�:�׈�Z`��z�'��f�=W���eg8kio9����d}��"�,n{�4Խ�� ���^��t�����.>q�����\��E����/hϻ/�`��ϼ�2�z9�����׺n0i���K���Y�V�R��OǞ� �<�qya1�%��>��z}Nf����3�Gq�h��xW�x��Ͻ|Qs����V�1�ɞ|]ڂ�Z��P��6̸p�Z϶�2����{iZ��o2��1�O}��"tR�u�r�7-Q�¬0�7�˾û9n��.���؆tm5�
�����۩ʏ�ժ�R54"�	XmN�����Q���ffL��&���Otj���}tx�1<��1��B��2f�[�ⳇXƺ��C�l[��nz��|t/��3��*�S�u*׫��w�b�&�0�s����q���߽m��f�CCہ�3�+q:�G�q�eUq���l��E5xz��3)�|�m�ה��kT�y�x�<�f�a�r�uKW�]H�`�.$3qݖɭ.��׻����O���'�z���<g���[�1z���+�v������]L���ٓ���7�^��\�l/T^'Ϋm�dr�ng�\��nZ����*���6j�U����p��n[�E�昴@�`IL�C��iC�M��%6����b�衾G>�p�{{`�*�Ҧ?zl�TO��!g�B��u��|�xԉ΢�gI���Yp�?)x)����G���f�״�:�*��cc�����[	6]h��l�6���1foL��O�mzv�'���������Y:l	��L>�@T����|�]�K����7���c7ͽ+���T���rX`ؒ��K�(걹w|�K�r'5�KԳ��پ=�*Yh�RbkfTVC�ەv8?ju�p�z�\q�"��⠙�Cڨس�oX6S��V��h6�헝O<|Ϳ_�$��_*0zT`y�έ�~��u�q��?y�n�Mj���9�7���	�ׁ���VpT<	�,���6+�_����p75���v�s�(ݻ��^�	n�ǧ��s��0��P����J�Y��r�.�F�/o�n�n�)��_����F�&ӻ�mqI��f�ხ��N+:|�_��l/v;�-��f���ږ<��7��Q���=*�eK�,2;S܆��3;�w1i�q=C*�;�S���n�=��Wy�bW�aX�ı�JK�R��P��A���Qp�C���b��W�׏���$�l:��9ˮ�dC������[�0�7	G����KG��[�&����xed���x���zT���!0�oWlfƴ)���U�^JE�SZ;��d~�{엎o�E���qFl'�M�e���g=���a�ƻ�L*��+�t��-�O�����H����E��V�T�ozcd����R:皭�O<��,/#�8�j��Gf^�鬃W32��\�^��Ɛ"#%��(P�y}i�v�j�SnqP�$��a�*`0�ch,��>�ߛ�Ǻi��[w�5��6�5�q�o�����Y�t���i5�pX��*VY�&_T�']X���vj'#s(�d���Eƨ֤�L����5��5�C���<��z�������}dq)T��;Q�8��৘�r"ɍ���gc#z����3r��ǉ������ M�9a^dY�(��34Y|o�ʆs}1t}SCն�'���xT6&F�Ri]S#�X!����8�>��*$f��H��5^���r��w��8�kC�&��C����Ȏ�>^Z):K��{�i5��9uw��)=}F�pIf,87��V\P��+�9D�ܣ�<�z�L�<�޼G�0���ܯLUۏ�e۳�.Ɯ�~ʇG-/�tU�s	E��.��|���:�y%g���$mc~��M���R���U���Z|+i'�x*מ�<�J�����<G�� p��E�����l8���.��{jY��k%xd��/ҭ�����Ű�cU<�5�M�7��=��q{��Js������<$&ϵ-�%%�	u<�:�����1��/p�?N��c�K$�j�s��L�����Z1���a�
]�X�2�,�`y���:�c��k��Q��h�,�>ۦbr�N.[�K��m���VLRk�&
��֨�G^l{��&K^�����*�v�#�b�Kҡ����{L��+Z�2��Κ�B��X��P��}��9��O���O;�fNΧ�3GM9��(�C�V�]�=Y}r���^�hq�"8��ݞW%��es�yz��b�2y�z�Q��Co�����q���\K�P��5E+5򹹟Vj���Y��\�.Y�5|���̨��wq���nf�:�P�F)t�I�]�x�8�K�(g��2OX�����o��>���T�����o���޾���R���uK�]V������e3y�r�{�д�[Ͻ�ۚ�׮|;����ΈCx�@떪vl�ڙ�Uǡ\s���z�N��9t��-ܗr�����x�K�Z(nqw��Y)��g�m�x�S��lS���nf�d��%��;!k<it���Ś1R��ɗ�����c��Ӹ'q�U�����L�������O���g�i=�1j��o��־��]�I���dx"�,8�'��G����=��W�wnro���7m״�5�ܪ"�)��">r)+��	0���I�n�W��S��_�JY7:m���I��{����j�#���a��=���>�z-�zs�k�_���q���2���[���nO�@抅ն#�I9O2r�J��Y�<�ꕯ�ov��X����TJ,Al���Z���2�쮈�<�W"�/V�1��4�{V7�J�1na~S#��zS��%+���]cW��(�H�rj��R��{�+�\��(�}���}XT�:�ϗ�����y��&=8��6X�-xz�'茸kv>؝`R��~�;�f���[��U�ܽ�8��s������^��r���H<^Ӎy�׹�QO���i��p�ۗ�r���{�z8�������i���Tܼ�.��l�7\S�/S���[� ��7��s� \~yڙ�Rf^7���:�_��gG�gЖ��P�p��<d�tC�����{gU�z�g'�sһXVtx���v�T�������ߩ!f���loڝ��w�����x$�ޖu������K�6{[�ٻ[�ߣ����=:k���f��q݉�DE��Y��S�=���lW��}|��p__vt���GT��w��}r���u]Xw�^V�k�_?=�~�ĉ�8h'�7r񝓤׀)y���%h�=n�.�hOfU�p�i�z8������v�x\���Ƭ#ɫÉ��۸ZW��J�Z���7oN���r��kUwt:=@��7o���Ojr�2,�%�3��E��戵+�vd�^�\�t�3�{�7��9��I1�	�f�OY�l��h�r<|���`������eA��J�x�
N�����Lx�u޶����J�6�+Jt#o��]�M��>´7=�eK	Z�e���
�޽���K���w�s<��]כ{ڌӕ�ݱ8��'��㿴L.�I�<�QJo2�*X�O���T�{s ވל��[����]N�oE�/Jz�]Z�e����=�ꣽ��bַ���}꼣ޗ��<��'�L�@o1�]�Oc2y:~�þf��yO�}ٷ%oT��7/|�/&M�w7�:��fc�q<֪ƽ��,뿓񫎾�4Ŏ��3�,��c�~��Ls���9�Y�y�8��}s޿���q�az���V��1��י�Z��7�q�ם����o�.�z����=7�g��sΗU�8��x$�iׇ����ƙ�Æ��$s�s�d�z��2�*=�GWAMQ#��{�*+�6B�O��E�T�lvE�{�+YuN��{������v�^6x{C�3�������WJ��՗���Ӝv.��c$˭� Y6���7��Q;t�^�ktSP�u�ŸiXfX�ѵ�Umy��D���z�lY�&s�X�m.��v�{Z�ڕ*_S�ǘ��4�y5�'<�'���tuf�� k�۝�;��)�W�j��z�?}�&��F�w�~�����w��X8�v��<RW�7ط��&��!c0Q�-u��;����ǝ�:�bNy~V�g����߻�.c�v;��JvB�0��s�9������O.uܽZ�6-`�R�vfs����7+n\�c��V�����=������L�fq}�7���^�}���`
\x"��xk�n`�앬�Z{(ԉz6���f,7�ʼ�:���rw�����"�,�nPwN�a.yu{w�r�8s��ޙ���'��$�ʤ~&����M�-����=�o6��?��t_,{=�N;z�T���V���%x����0k�o\�9�Dj�*���:W��1Ӝ�&ߪJkU�ڨV�P���J�r�sz�o��*����2�Y�׽��������;q!�t}{.n`��+ �t%�p�oJ����&��R|l�S;ˮ����Ӳ��n�5�$F呼G�l�pt[�Wr��]��ǔ䲎k ����9۽�}�l$eq�6C5hԸO���#�	j��ݣ����i�ӧRnKٱ/w����;z�񫎇f���,�<��ݝ�f��[��z�Z���|�f�9��~����x�rQx|����cԒ_n>{�D�ٌf����N�8��ǚ�]ƛ�������d?Q���앷s���̆�pl�ܴ�L����/�:�������p��x`{y������u/��A��cf�ĞɦSɳ����2��E�6��z�fW�h�����s����ٿ?9��l�Y���dٗ���}p�� �}bY��:!o(�{~;6gmL�+[VW"thU�Ox.Is3#�vӧ����2��o��腼a��>�:+9������ط���W#P���'y�%���}y��w0:vBY㛴/t�L��>[}�eo3ӯVT��V����Ҿ�t��;�"��%�ϥͱ0K��,>��^��3K�~yx�뮒.=���)���n�/�}ӗN��*�}�����U��˪S�^ZA����X9d�v�lYw�t�֜���Ku�+�cy�G�9��8��f�`p�U�0�ʜfg}�ejj>�q�-���z�u捻�:>���ڱSho�c����Ԓ�O��/��oH��Ru{i��o�_��=��%��ϓ�U�}��z;�f�9�ܻ�ӂ{gv��{τ�t�lz�wO��*u�}���$���G�/��%�懑�9��U�~��;�5�s�a�zs�k�w�a�����n�汳Wv��x.=�}]��_��po�g�Lzq�n�����ߨ�A�r<��5䕕���k���.Wón�pm\ߛ��q�29�O��	f�.��S#�/R��wY�|9m�^N��ulO�e�z��zz#��)Գ-{�m�b|��'ϼ6�(��г��հ��2��nZs�g�ީᷩ�;�4�=�}#�g�|��gh��/S��[.����1!�a]Uu�{k�����v�&�7�m�o�Y�>/��{?(���8f�rk�VB�q�툖>:��(V���lŠp��u�������K:��85TZ����ʹ�K�IZ�nҺܺ_>�Ȕ�k��c�T]O&��c�]���1͹��N/%�	�v����_�lg�S��Oa��!�u�7��[���#�Eiz�v�(ԹH&hif�3�����Z�
��\�2u��7MѨky���Νٺ�ӣ�<��.��'��N��cjLmnRB�0��N���u��Q.NdI?�Gݽ�(�AF5��{k���;�?<'6S����r��S;���Gz��z���y���0�o� /u��w�'�k��f�c���<�oM����}o�y�u�n7�P�Ó�Kd�x�3&;/&X��6�CK0�k�T:TY+�疴\"�{z��O*f
�S�Mc�B����*�*0�a�6���c+���,d�9��X怡ֲ���.��-n�zpz�N�wA`!S
^p��V�eũ���w���llEE���խgzJ[y¯��;�es��3\�i<*��j��tm�bT��X-���]Z��x�ו@�T�O䷡�K;��|�u��`�-_WBh���*A�u�isS�t�XG��:�H��T�h������❳J�Mva����O�z���1z����l�`�>�����N��iSO�NWL�M�O+D<r��7K�k�r�j�Ϛ�5�)��Z,�w�N��rn�{�����M+CE;�j����'��
��{S&O��u�]k��th��rY�u�+%��Y���[�\���:�]o�2���;V���X�1���Ky�O�5�fj�@�=�wh���:�Ϋ����7�x�v��޴gA\���z:�sG�����t�������g���1�^�u����[˚
�M�էh-�*��c�!�2��7�Ou=�����o2���|��|-Ge��v�+��¹>�-IZ뫘�ٺ��W}]\���N�/�߆p�Q����r"iǗ���=�
��'�Ɋ����^rC,�n/��ԡѾu�g%:��ñ��l1m�t6к�x�o�s�TD� �;���Dr�{�V5������tw#+f��z��V��W>�����+H���VځG�q��֕����>w3�)NǕ�*U�܎�Â(�7q=����#�!�ղguj�t���Ӂ�9���c��n���c8�U�[�����,�7�n�9׊��Tw�s��A��,��eԻ�6@i����J��̳n)��h3z�(h�5��A6LoV�B�k(��r�1���mw-Iƃz2�un�/Db�'\�§Eeq�����x�Ժ��;%���lՒL�Z]ˎU��Y�5��g�[�`[��t �lv/�(���ڼ�@%*�i��-�|(��*�7׀k`��2�
�Zw�ķk+V�=�����\��*�V8����W#���z��h���eۯ:�x:[�o�$�I?A ����ը����	Z��AYF���Pm��eP�U�J�+Z���Q[j�UX��R4J���J��V��V
��"[T������`��Q��4����EQ�֢�UTEkTb�*"ְ���QUQ-�%���"J���-���Ղ!l��(�*Q"�m��J�����ڡcb֨�"�m*�"��������c�IR��PQ�PUD�F6�kl����*+)[A�V1��� ڥ6ԕ���1DQE�j,E`�,EAZ�)U�6�����m��� �+Km*� KJ*��R��U,V5���b�[J�ҰUX#b���m��
J"ʅJ����Q0�@b�0�QT+A�eW	S	U��1h�UE�,�
�P���hZ��,���kX.��kZ.9�&=��BLW�����܍i[m�,8��/w�Mi���{[�OCk��0L��j)��sS~���ި>O�=����L��~�������l���%�h�,Q�q���ww���K{�L�#�����J\�m7���xNכ�z�<�t�*QɿV��սz-]���l��k֏��I��T3��"��w{�^>٦�f�S 㔺�<���D��t��0�M����܅�3с�k���c^Ք+��&�aGm�o��;9�6�U5��	A�+�g�|��{[�1���c[S���P�g�*�R��#��z�c}�<496Z�	�z�=�b���j�X^���<�el�C�sFt�X[�z/��t��ÎƉ��
+��}���|5=��ǣ̙��ۛ���q�cӃ��R�a�U<���}�<�w&�<�{h��W-kz��������Ø��Ok	�εux���R���E�W��\h�#�;��yV�������g���U��ڐ跳���m�7�1�~&��I��2�nSK�շ�鐌d���c'�]�۳�-���`.�U}.�3�S��r�n5�^R;�K�wM�n]k����7'b-�G�	r�S���(!Ƌ�g#� &mÝ/�����6�y�=���Ϭvo�⦅��?vb�� ϶��ՙ�1���K�?-sK]��=��H��K3u�v�9����e��uLq�_�]A��gf7~a�d�).a����X�U�_v�v��[8g
5��f(�<���f�N� ~1����%�L.?w���t���� |d��y�̯>�+�}-[�W[.���S�g���y6�G���M��o׋X��k��-g,���E�w�n�;<�+������9�l;����'e���>��WH�ݹs�uᚈ�e�<����;]<<���D7��wv's�SϷ\��v^<��7DX�0����V�o϶]K�Z�<j�q�>���n}�߳�%���v&N�CY��'�nskֆ�]��M��ҢƐ�m�=��C)�+r8+E�&��o�L]wY-��zϣ@��G\�����_���ݒ�{���*?,�y�n�H{����A�]���*{��!�z*R�`��g$�v�Q�^�;#���6�\G-��B�*����q� �tx�swb�4�9F׫,x�]Z����km��﫞��sgz
����t����EL[���Z����i��{�/D��p]6'<�γ3��ݳ3z#_y�h��zww�t�q.�WkG�G��l�[ w]~Ü�lu�+N��yV��4���������yLb���ot�zo>1��8����':����zy�)-��j굧'��f�v=�ꓩ��}������v�{��n?��ߋ�7V�#K��� ���NN_�������[��?W��4�������T�������{�S���϶ܰ����{�=�y�Y�C��L���۝�N���3�F��-6h[l�lg́���9�q���͝M*�k�\����}oNtVpq��uK	l������$��i�M�$a�<����ɷ�G~�2��;;N��������+�u6o��m��I;O��	\�$��ۮ+h�u/��q��`���t��i���M����OP�F��û1�')n�[݌��!ED-SK{R�ﶸΜ4ԛ13�86����N���Wp���*�!���%�Ŋ���d�|@P��IH�hz�e�c�:������;�O��I^���6w���������Yֈ��X�u�C�_S:��XWG�����ԛ�U>�y�s��X�痓$��3��N�[�ϻIs��^�j^��ofM��	N�e�I�c�ϓ���&o�K�ɒ��ӳ��Fyf��S�v�k=rl��=��dݺ�6������� ��|2#���>�:���u��|s|ҏ�'�d���V)��l~|ߵ�rdx"�1�����*7�ޫ~�� {�c����W�ټ��~�m�����̝d?C�`4�&�:���`�̚CF��2L%`>�Ֆ��6�evm~����߃#�~Q���m���P�&Ұ�s� ����s��$�f�\�N�ċ'�`~��L�L��,�d?Mk��4��?gw-��g���f�ǿ��g︁�C��XT<o�<��*~��2q�����I�T5�`��l�~�O2}�bJ�w<�&��<�1a�O�����O�߾?k��}������3��+����m�d�$�;��,�Ato�$�!��py����<�ԨL��&�u&�P��b̛d�ޱ����X��6��~�+|�*��3M����O��p����R��	�u�C�N�>9�fY:�G�&��'�]�	4���w��L�M�_w�:�	�^�y�Rs=��6�����Z}����~�wE�����V��.0��s���6-kL�?��F����%�rs!�b���W��+s�)N�P�-&A;H�x�4��3X;9�9�X�X�Gd�bc%��}��ov�q��1n�A0��vP�5ao5X�+�$�4\=]���嗢g��C������d�����O5'�N�LY�̙L��̓��f��y	��P���L��I�:�����<�&;���$��h~?}�����T�=����=�[�<����4ɶL����$�$��c8��e��n��I�'Y�P�'�O&qgXN0��f�PY&	��2y�3\��I�T��p�<�����������s����^�o	��g��:��:~xl���|�S�q'N��q%a�C�h|���C8�'�N�LS�hy2~��	�|Ȱ�@C�߈G�&ލ�ܿUUx���3��y�;���x�N��*x�ؐ��a����'�h�1<ÏY:���8�|�3�ĝa8�����CE��+'X�O�q���F�B��}�Dy�+{�ܷ�����[�*e�|����:�����>@�'�Cܲ��:{X8�'Y2�ް8�&Y;���8ɐ�q
�6���ĕ&��g��Aa��s^c����߿8�<��?z��ɤ�$�O&Xq0�8�<��L�e��N�{�{�����u��d�&Y4� �ԚI�]�	!~�?z��>�~�?N�9��ǫ��w�>��ݾ%AB~fP��Aa��:��:�$�I��6�I�~�d�A�0�v��?by��'{�=d�0>��O3,�a�����}�����p��ֵ����y�i?2{z�,��~7���1�䕓�Y?b�ĝI�d�a:ɴ��bjI�g�ba^2y���d�}uK�����W����׿��ͥ�H�1t�N�q&P=�`�fY8Ś�p�m�>�d�C���+	�n�aY8����'P<������u�i�bjO2ur��K#�?~�b�}��~�}�~�W��7�a0�0�����Nh�����6���P�ɴw�C�|�����9�%J�vn��d����M�{�(�������R�o�J���#�����t��Jb�%�����3)<}��N�GS�_��s�.��͡�m�Ȏ��W$�!s��KGK��u��M[�~��m��7���;Ww��򕝳�7�ӄ(i��8{�U̬LM�v��o��仮��.O6i��꯾����۽<�w��~2u��=�H/�e�~�<�0�����y��{�~I��}`��O�Y��AI�N��	'Rs6|�}����>'����Ӗ}*�~���cw|�zL��&Xu�l���M?2i�}�bٖN��_2L%aϻ��,���I��}fRq��;�`�G�G�7+�?�����?s:�S���U�\���I>|rȰ��'�3d�~L�Xe�̇�k��M$���@��d�S}�'�y�M��Y%Oƻ�̜J�g��i�Y6�����/{?�_?��:�s�����߀��O���&�>͒�I�N&�XM?$�2b��M�ɓVa���`�e��<��;ĜC,�A����Hy�g{�ɖI�7�g������1�X1�o\�7[����N%d<s�0�&ݤ�l�6�Ú��O����~d�Vo�~egY&���a�a9��	! �����@�~�� �N�s�����e�;[���/M���������t!���C��Y;�����u�̝v���0�w�bJɤڤ�Y?0�1d>g�O&Cu�|�?l:��w�o���k��\��h�\���P���(r�I�N�g����I�31�fXO0�y�̜~a;��0��'L��:�>s1�IY<��9CiY?$�+!�0��ײ�3�������~��}�n��d�C�<~����*d�VMsXu��Y������?{���y���2u�'>qē�2w8��'Y�ĕ��g^��k���}�m�y�o��+'䟙RC�Ob�I<����<��'���u��Xv�a�O:C���B�y�u���O̙w m�&�5ݸ�y�L����߹�_{����o:���|J�?'��Vd?Zu�I��Hm2y*V�:�C�3�I�<��y��Y^�>d�'���oؐP�;�|퓌�I��q�qp~�7�/��_�)n�����/s���V/z���/r�3�]kFn�5��~���%[7]��e�3J=�4�#�wf��{���eEu���9]�����p=����Dz0�΅��q0��pI&�j�F�b��_GX=/���mv������� Yg��e?��!:̲d�
�6�Œ��3�8�I����q'Y<��$�N�P�0�u����'����|��,�91���ݺ���������8����߾�c�Y4ɔ�͓��L���k�fY2wX�$���IPP�g��J�P8ì�N`��@�~��!�d�f<o���w�~޽n�c�߃�'_�m�6�4�L{Y4�q�q�̙a��}�<�d�L��	�?2o��)'P��%J�fn�%d�VO�0�'����{�� +��ȴ���}�_�e��ϫ�Wцg>��&P����d�|��=�)<�;���N0�����6�̝�y�{4�;�������Ϲy�Ƿ�α�sx����}�$��́�Rm��O?�3���z�e����C�����k�bI�T<�'�y�w^�?2u!�X(u'�,��`���L���t��~�3������wZ�8�>I﵂VV��O:@��O m�������:�~ְ~d�'P�s����&�jo��I�T?���IS���:��ƿq�ݵ��{x����{\�8��*9�H,>d�����q<�$��Ogx�d��O&O�d�~L�Y:�~5�3̚aԟ�`i?2y�ݾa>B����>����3��?sY�]{Z��w���
ISӛ��M�Bd�q4���J�S����?g2O2d9�Iua:����&S3d�|����	�S����I��[�����޸�k����7�6É8��o8$�a��`�	�}�<����}fRq�יִ;��N2g���'�3�'�d�'�3'�2�Y�I�*wf��c����_s����}�B��	��`�2��M~� m����8��2c�<�d�3G{��ed5�u�̛~I�=� m��~ĕ���>k'�N��=�cߛ�g���T������H9>P�����d5�µ�Qr�˙�CѡF#��;q�*���]�D;wx�����Ys{�S۩(��Ɯ�]>�^�˴+m�,�.����]
�l�;��NK�B�SO�U#9���W��{���o�$߿s���s���g�!��'��b��O�S�͆زM��N��|k�hu��SSy�'Xy�q�L��a�^by��XM��y���~Փ��O���s�o&��{��ޝ}��sO�Y2��hu���!Y��egN!S������\Y<�!��b
N�u*g]�'Xy��<�y�%�2w�	��.s̾�;�����7���>��I��'���O�'\��	Rm!��%d�!�~I�V�M��&y���k�N��2}�AI�O}CA��B�y��m�y�̿������~�}�>���$�Nc y�'h;�T���3���m�Œ��CV�䬝Aa�����N����N�߬?g�e��B>��~%�����o���Z}��������N�m�=�bB�y����2u�,�=����I��aa:�dϳ�T�l�;�V,&ӈVN��Դ���'�&$���G�m��Z����}Щ��=�؇�;�����O2q���d�	��q�M2e�G��y�d����b��L���'P�w�$�(LMӈVO%d�^]��g��n���}��<���8��OLI�f�C�d�N�ì���=�&]��;�,�a9�y�L����ĞL�q�SS�ć�e&}��:������ss�����k�k�����6�J���>�IRi�%@�O2w�>�a<ɶo�k$�sVA~d���'RO=a��`�2N������ w�O'�M��;�n���~��~���z���o�4���	����T�&�$�8��Ru�l�?O��O�bi�'�:���`���(g��u��y�O{�y$��~�9��׷���c�{��u��R�9�(m�h,�w�	�6ɓ����y�gu�*V��YNj���N�m����d�!���;I�N����g�4�����.l�Y��~��B>8��Ş`'�&�Y[I�B�W@��fӝ��@M	[�io�\�p=p������}	I�$f󏙁�mc���`��u-��ړ��Ϋ�0�`�,�t�/�t�.�*ԯ�B���Ŭ�Jk\�ޖ��K7�w�U���o�s��3��[��&���ԛa0��?2q��N�P�&Ұ�=�
O�?�̓�3�bJ�wvE�ٰ*d����Xe���u�{�v�X�3���}��}�7����~$�O�zw����'����0�aP����,���w�8����`4��6ʆ��Rm��}��I<ə�bJ�w3����'���ۿ{�����~�g|�=����I��=�a�����e��8��;��,�Ato�$�!�}��hd>�2u*^�):��T7;�@��l�ޱ����>�Q���<��v���S��'O�y����'R��t��<b�l'��i�:��i�?2u��bM��O ���C�d;�O&Y&ٯ��̝J�ׯP<~������-w�P���Y��\���|2~d�oa�L}I�R~d�fb�m�d�fbβO��(y'��ͨa��,�9�$�d�Vky�N����'�}�x f}���i�w��6��s��N=a9�q�������$�$���q%d���8ԟ�u�	�a���,�	�?��I�ypd�&MsQ�#�~Dv`��o�mc_���s�{��6���u���y���&����'�5�ĜI:��J�l���Y<èd1d>O̝J��m&�ȡy����iU5.�Mh�}�?}F��IԞeL��HVO0����ē�5;�O0��N�|{�$�;d��q'XN&q�IRm!�Z2�u�E��<������W��ٚ9?���e��^����h~O~��~d�rs���J���p y�ۡ���
����v���I��b��&��b��&g��VI��;�|.��_W�U��ş�M8��=�
�wT2��`q�u=0Y'Rq?fÉ��q�?`:���CE��N�{�{�������d�&���4�.���z���vw�Β�~��:��HL�6�R�-��"����
zҼ��I�7��rk�K7u��+�7�Ef���Ө�Oz�Y����l'�t�N��Y�d&�E��L1�wҖ�T���J�& h�����C��8�dZ�L��\�¡�)��e\P�t�[�7���w�ꯀ'w��=��k?���>�a6����	PP�՝B�y���I�}0RN$�e�-�u�sX2y� ���L�C��̚a:w���M0��oW�o^�=��}�뿿s=�~&��L���k�L�g��,��~�pJ�����J�䬟�@�N��(�u�i�bjI�g�ba^2y��{�&ޡ�����{����������'���'�@����fY8Ś��y�d��$��d�XL��XVN%d�b��d��d?XN�m�_(������_������:�jNo�ԛa�����}�L<�;�d�O�6w؂��M��3�ć��&Ok�I�͒�I57z²q�f,�d�'�S_���f���~_c93}﷾��ސ���&_2i�h}�bA|�,>��$�V��0�	����2��)�؂�Y6�̜�)>I��q?$�I��%Ւu�1����K~q����}�s����}�dˤCM��|�>��'��&��4��>s6̲yo��$�V�� �J���'�u!��I:ɴ�4s� ��L����0<��K����ǽ��\��k^�a:���X��I:�ݑa��N&LXu�i�2��'Y���̚I�gx��2��.�I4��p�py�T�k�<�Ĭ�ύ�0�>���ί��k���?}�#���x��o;ē���kWI6���b�i�&Y����g�:�����k�,�I��$�d����&���uw����[z�~�|�������;�d�VC:�L<ɷi=��M�s���O�$���d�lń��egY'�S�0�	Úq�:����F��cZ����~���y����C��A��Bm'�ɏ`�2�|����;�	���O2q�'s�@���ϵ�+&�4��d���,������,�$�*z���]�8��Uc_�1O��+�A�E����]X�����v�yr���\�O8m���������$R�.������}�����<�.%{)c���f��8'Eou�r���r�<NdY��%vl5���莮���u���:��mhK�9S�0��B�=BT�U��ψ��W.��@un�N�X�0�ڍ.chnǬ`o*�ĳLwצv3I3&�C-[�C�yQ��9Ls1ժ�:Td�(�L��{x�Is�55�|.�+����5���P��\�Yѵ�Π&�"����J�Ė/��:^:�� Q��ǧ8�J�S��"�<�?,g'#ƻ�Zȷn�Kq�%�޻G�8>3�Yw��'*#P�V����������l��y������������p���,��դ�܋.1�,ƪᅝha�u:�M��ͧ������tl�Ξ�ɴ�r�R�*���[kj�=%v����I�߀�K�P;3�i�y7~#��E�&�Eೖ^�Ȝ�L�����C�U*>�^�P���9�2x6�\	������=�1��GdZ+��,��	ƣEfuެ�:��LK�9��&۩��qo[�K:�iq�a�&wEO:�>��;d�&v���z;Kc̻|1��
���0��ZL�'K��k{�Q��:�e����N��+N�)�(�l��i0te�j�3�&��;�C{-����%���V_(I�
S\�]ܷ����w�'2�J�y�w�(&�bս{ɰ��ӮӉ�i�'v;��^R��X�����Ώ�g_r�D+�Yp���-�t]:�1�B��;�mt�Q�W�:�>����ƥ�V�u�D0�70�P�ww%pع��yx%�Ck5�[�.
qmM>�����p�)켤�-Wa��YB	Ձ��o���	ZH�bt������ �C2J���{EU(T��*D�N�㏓�LC-��ؙu߼o�M5,WZ٬�ޞU�z�!�jȎ��]joE��M��Ѕ�r�<��κR��xň� ���,Y��nǃ�{[���E����Q�Ҷԣ˂���ݠ�]��Ž�"� "䱀JKv�q�Q��'_'�o7�ZWmƏT����� �Q�U�j}3:ʤ���;���a2��{���T�/y�Z��,[$�dA�=.�ɒ]�2��Z0��\6��k�]7�Q���J-��8��K���lE�+�;�j����	������ݵ��l���aF*�ׇ��7j"�%&h�8��%c�����BM=կF>�T�B����'���h^�85�k[h���k� v�9�75��`�(5����Y6�
��w��b�Šov������W2jՎæQ��[��ct+�P�%�Q���^��\�x�bUm)��Ɣ�Su��iΫ�x�����r����W��������W	o��:�R�!�n�I���o~�3xc�|/~���s��� �,���Y��q.,��B�Z�������Yb�*�f(T��ʊ��
AV,X�U"�iX�J,V"Q%AA��+Z�\`�J�-�R(���A�,X([VV"�ahPbm��A������*"V��T��QR(� �DEU�eH�eL&���EB�X��h�kQ���Ҭ�1Q�H�IV1���"6ʀ������ƵQQ���TRڂ�`���
��PX,ʋG��EQ���U`#҂ԬA��FH��VҠ�Q�V+jԋQA�0��h��m"$Q1`���)qT
b�U�)Y�Ub��(���QEX��QC�%dX�**6�ID����mF�D@X-jL8qhPŨ��)�E�U�+[Qdb#����{m`�0q��za�	��iWV��]�A������٘;�V�������c0�d�Ү��5|m���`��?���_om�ݓ{�@��ù�C�<�����
O2u+3>�u'�Ɏ��2�y��0y���&��u�6�����:�>o�%d��l�~����<��6z�����^:�|8���)�\2N!�g� ���qP�'��3�`��u+3�����=�=�$��2u�'>=�O�$��'Y_z��߹���k�ɏTd��~��R���C�Y6��ɊC�~d�g�I�:̟�y?2N9��C��J����d��o��wV{v�'�@����~��\7Ϛ9;��5��}�6G�h|�'S���+��:¤�Ť6��<���N$�f~��~I8���C̝��j^�>d�'���߱ �>�i�'�y\���w�ן�����3��	���������ˠ��e��u; �2yK�oo�XO�w��L��㽎�ۜ��L�/ηa��x�_.}` ��-[��.�oz|�V�S�=�LmK�fV9+nL�c遺&Ƴ�+��Vc�^�$�S���[7�f��ۿw9�)q�U�p/M��]<��v��α��I�t�X[:���n_��1툷#�pa��s�_��V�.c����{��ݸ���\o����Is��s�7�N�A��Ɂ�0��\��;�[�6�Nqqû}jޣ���ؠ(=6��ʺ�f�,���r��vd�(=z�v������5�Rʝ�c|EӟoWS�N-�aH��g�������Qy�J��}�YqL�5-��6��p�Z��[j�)g�����־���ﶃ����o>��7Kc<Î�x�v����%x�k}oO{����{�v�����t��s��6�~�;>v�?5�4.�]��6f9�f>�>��m��~q���������`{�e��օz�}Ԗ�_�uud�kǌ�\��f�+��;���`n3���<��~>�\Xnċ��y����g�T"ݡ�y[�l�=��n*h=;�9ީ�����x5:h�<�3�o�X�#�z^oP{n�ٷ�':t��������6���^�[�$���g�'gPuv6ly�=��K3ɻ^O_i����~3��gi���� v;	s���YY�m��Ɲ;'+��T���=<����W�7��������Έ[����I�1	�{]�䦖�ܵ�o���/���*���;v{$��3��A��6*��Y
��KS�o��ۮ�^Z[��8��>�N�#O+�dF�$aiˉ|�m�;@���M���9�w%�Q�*��V�ܴ�{L��E��h��rIՒE^`;h�{z�-k;������PQs��X�Yq�?>��G���m����uO�����>Q�s痒{|p�^�`!�[�]�9�f�d��Ol����Ҭ�V��	C��ɤl�����4}V)�o�v;�crO�oC\2/}U}�wo�!�Tx\8�=y^��ϩ�L�m�R��}��h�L��T�{�N�J��������wz5Z/���nM�2��g�vR{�Q��f������[�L3F^�z�ϵ�k�Er[WX��U�k���Y^��8��6l�f�AVe@q������L�wm��zi�p�8Xs��6�~�fݭ�0�jh]7:�[ٹ�Qn<���s�^�������ߜf�cӀ9��ڝ6���K�t��ރ��Y뿓�����L]g�V�7/W{����t�u��=~-G��ϓ���{٫�=�P�'�B�;1}�p��n �ڻ�5�x:����󬝱�{�s�G������ov�X	�6���y����+ء'xgۮ�;wv��Slz#�z'F�(˽��f�
P&�O��h)*��ܼi���h��L����7eJf`�>@%bK��u�n�p�1���=O.����چ�Ŏ<���t�k�1'��*}6�2��E�����b��\��YW��W?���}�������/Xzm��	Θ��=;ݟU�����v�N��/@�*^��}ջ���f�����1!������3�7���r�XLb�c�����ͿH-ڳ5{v��������Tf��&��8ɝ��Ny8����;3����o��C���*��2l�r5|��W��.<}�G���=0n�+ْ���xg;���u�BYb�3����e�C<��,��+�9F٢�~�B���m�O�u��y�otF��'M��>g�ܺ� �ך-񬘏I�>�����7N��K�*{f�g��;�6����#E���_rƐ����u���EOq�Z-ɷ2��sY�K�7{+���$>}�f{GQ������nE`Il[���3�;����C���W�]۝���#'r}��Ko,G+3=��wm�ވל�q�-��j�VW�)��q!��q*Ul:�8��{�)5�c�I��b~gk�`��/S9+�/wJ�U�QW�P�츓��M̨a���)��.���tW���ے9!�yգ�,��yW�����,=������r`��6��N���0��c[':�Y��w�������H�J�]��JɁ��l�Z�+N�Q+ǖ��F�/m>�X��ʅ� �'����K�qn�ӓߞl��נ,��{/�@vm��޸�`�����lZDM�>�O[s�N��>>m}�rk*���ۣ�︼���3F%3�����LG�����/�q�z8��&}^�)�s�k��買z��\�#����f�E���l�<3���ܴ���#]�����W�����Z^<�q�uM\��Tm8�t��p�86o�Μ��｢��Aw�)d9�s����X��m�������]u6o�I�sɵg0H�-�����s�~����ݝ�Gh/����j���u��ް�y�~��};u)�߫���3|���^8��ô����;��;���闝dJUW��in�UN�xv8%M�'<��d�r����vF�D霚���ս�����Mv��;`K��A-��5�.�g�$:�z�CQ�W�{���Îe�qf�mnPT���mt{�c�P;�G�(v^���tB����b☳�Є�}C���uʐ�yQR܇�y�/H�����K��!�N�g7�z���| �c���2�'�c�w�����
O<)y���K�>��u^�܀KE�w�,)�cV{�9ݾ�pϖd����fX�����`R�ȫ���Z/�&�v�6d�~~ڸ�n�yL�sL�5�}Or�&��;���r8S1��C->T��/yOf�u2�_s��MΛw�N�o���{�ռ�G�\��C����ݹ���ۍ�3���6���Î�{%�O=yn�=1�'��5�{�f����9�66@k�`9�N�k��c����x'��~�.���N�s��w�����y/�����ɏw�9�c�y݌�]\�F�E����&5��_:��m��l�6�XN_�7��v�[��R�ݺ8��[o$���4���u�K��ƭ�6�b�ßm�'.a���hۭ쭣�Op�s^m��o�Xs�����B�[e�y��cp�U�+f�Q�^��}s�$G�d0���[��WyObftͻ�����p`4k�cM�'<̓~pՎ	�F<��5��w8�	�yһ_G�e��$zf]��+�u�=��N�\��A��;��ټj�7r9@<�����ݵX��Ͼ�����Y Rfl�z�}�c6�_;�Y� ��y?%��Aݍ��t��S��i�������ɳ k{�=3nY֎��b��is�h��P�U�m����q�GQ�<����+���f�d���;A�x��d=�lӚ�ꆟ����׋�>��?`/Ͻ�Ӯ{�^L�/ ��<-�j�z�/�j�[�#�9�����Ξ;���<'^����;�͗+n��u�f�˘�zm=1���Cl�65���t������OK����x��o�+�Ay.q����m�0JvN��>Oe]=��l~|����F6�Uz_��筮���e1�8�rm���=ò�{�Q�!�ʿJ��^Q�mSs�6f�9�lX��A�wN�=�ٳ��|8e�̞'��z-���D�b��s������Ø��A����2�"��.�oR�/m�R�Uf�X*�̴�gâ��73o`x�]�-�%!AY}��͍�7�V��8�ޭ}P�b��X�}��리B�|��K��B��<8ި�Y{Ղ$�]��P����LÝl��wf�����Q/7������;k^����m~�W��#����-kz�.�#:_��;����x�����p�k�==�Pp��G���eB�������|�������m��kޓѬS��n6�B�j��Ɲ���'�W%vb�{\3�
��W��ox��׀Q�4���w3J8�����7@ov�XO�lm�U����u�'�Y�x�S|i��8o��Nt�\~�����+;G�;^�IE����d�^�sg�Ra�����<cs��7���r�;r��1n��D߲�~���Q��a)�R���lߟ��N2���y'<ϧ��\�����_.{���q5Q�,�G\�9о�����3��\;��O=��&�M���Ӳn��:�<2���y�����vt� �f�7���^�n?c��,>��s_���i�g]���"��O>�A�nB����%nc��Mmp\O)3�{1_9��o�� ��.�[F��M��2�];;�=��{b��w����y����g�a�����o��u���E��)Wk'V�nX����Ի:i��s��(%��4��`�ם�<=MK�A-�Z��އ���v�����?���W�$�%N�/������~�%�ϥ͖�vJ�x�s��]���j:�U��~�[���=v5�,I��T�>pV�'��utr��'b��[�9�ve���W!�~��b]�툷"�-����y�uz/Kd�'��'�|�����μs��;S��J<�����y��%�:ޔ��;��gu��=U�X��{�~g�ӽ��Z���/p{�Y�d_�nĶ��c]Ӫ�Q󽯻�;5<��捗Ɓ[�~ߎ�B�ޜ�{<�	�\`m�Ǻ9)f��{���u���k���RW���	��6B���<w��s��s醸X�k�6ܿ���n=�s���z���q��uۤ�f��n?k�ɛw�7�6�b���r�r���9��厼����~�����M&���K�z����φ�p��������o���Z7���{^>�����4o)��g���kT�n�trl�C�=����J�ޒ��KM�z%�u���󥱅�"��Ynp�ϻNļ��`�m
;5U�w�(��xhW�L��4)��k�P�%�o(n��"V�#7~���b�ϙ=Y������>�L���mᏇW�1�u;	kQw&�p�'�L�
Z������r�ٞ�=	�u{�K;N��<X��Z\��]]c�?g�^U]�(�}�;K���ݟk;�����x㻘v���b��-a����ԏ9:EK�O�.������\_�]�{�N˗%�	�vA�o|/ivӁ�6��\���]�W.��{ˈ��fVk���d��L�2��G�>�������ğY�s������}�~�s R��w�ª�^̾�����&�� ��N��_�:hn_��@��n>"�J���/�Ǒ����Ǽ�A�7k~��:m�7^9C�C��(���/+ʸ9�s��Ώݨϻ�5�ط�}*�W5�NyW<�Kq�-%X����*��gx�i�vS�k�o\�cӝׯ���8�vz��AzY[�J�ٸ�s�Ğ�qgV!�b�A�PY8��&����7���5�G��hj*Q���q��]MѪ�At���G��okxl[O�+��Z�Y#K��U�$��0
�;ZU����+c	��a+��y��.���6ށ���u�m�n�4T�J��:��A�x�Ūg%�s@7s.!�1���:�Ծ-�Gq-�+e4����o�A�Jtp��F�ڽ�9�\�I�F��v�3&r��z��6�^��W]�w��M&W��`��o�:�}/QY�g\K�:l�@�=ɱ��V�M��SZ���c�6�l*�K�:Z�\��S7���u�n�`�{�L+�[��8�i	��r���P/��Wqz��p|�AVZ�i�in�����m,�q���hY���i��Suo|o {���V�#-���{���YZ�oĤ]����8��6��y��oj�I�Xe�\��:�l�\�؂���Y=k����<��i��2uX����D�Wݽ��6�u�Vb���*��,n�J��*Rת�{Sq�U��t�skd%�Bm ��*e�I��5�b��{Gh��e��}��qE��][جeYֻc]�u�V�mFl�KQIý.��48h�>B�R=0��݇Kt���B7e:o�D'C�BB��Tc�u��8�C�g�K5�6"7���؟Z�I���|&73�rr��jyg2�I�;�<7z�ۍt�h�[ۧ����}8�'����Uد�е��ľ�}���~����Y%�X�WV�0F����u,'����PPnwϧ$&��r��|�/�)��bd��ڜH\&�����^�z����i�WqG�W\�l�/nL-�S�8�: �ŜE���pRړK`y.��6	�k��b��l��C@��c�K��3��1��h� ������n��y�0��3�0>2�$��;oO�0I���v:�+i&����G�E[�|e�B�|�P8m����&ǤqQ��Gl��Ž�8��X�յ{g.V����a��-Ƕ8�-�ΚB�Z����tps�z��>�b갶U�H�oPc{]@�@�'J2ĬZ��C�S��|h�4�N�XfqO,�g3�R�(o$���d�t�ê�y�7�D��2E�l�e.����	r^�4Zѩ:f�Z+%7P���:�����X�S�!�T���-8��e;� ��]D�<1u�]�38����,�%�y"�_=��q��P��\H՘��OR\Et�mn˶h�Z�q
�V�	iQ����8:��}w��5]u}�kL�sl�a���s�v��5r��ި�-X����5��%��>�Z�'��[]��5x1�Y19�X����s�r�@_!�h@U�9�F��}��j�����pVL�Dk^�#��c�3nÔq���J�V��i7����8pk�Ƭ�զ�ᣴ�i�͝�Wd�"�L�O(uolf1����A�EͫX��������* 6EDJՈ��%E*�LR�TQXa�ŕ��0��UUR�EPTT\R� �b*�b�`����#������U\Z�
���X�EQDD\Z��V�(�b*�e�b*�����Z"�p�`U��j�Kj�(�X�����PTH�Kb�Tb�U��AAb������l�1DUFD�X��p�8��ҌX1Q����ũ�L�"����Q�QTEA
���"�PUTUe��E0ш�A`�p�EEU�,�Z��EUJ�f�*�F�b�+E��(�*���+���*���*[UE�)m
�6�Ab����Ub*�"��kUQ������"����[e�1E�
�`�EUQFb����UUqJ(��U�p�FV�� ��5������~�wwt9���3J� �fp�d������,�]�n�ֹΞ����t�YS�;�d����/ݔ��S}�|>�����9=^wW[������[���pm�<�7GǛ_w�څ�=2x��E���K��yw��Sƾ�uٶ�
��3o��/��nskb���}Գ|��a9���>��+Y���]��k�am���k�ۖ��8�-��ᶕ�:&��}��w5���ϖ��i�)�c�p�pl�Vv���άֽ�	ɳ��.r`�����6��ڳ�|c�����]Aޭ|u��T��*�FS�`��4�&�k{�=3lK;_:;@��Gc^��<S���e��	��}�UPT�{M�~s|'3yܿm� }rδ~3�j(�Z�Wd�nv{|lB�_�>�S�uG�/Ͻ��u�=�/&I��L�hv��/��혧L��}������1�qIևJ�s�~s�u���!h!���w3�zn�y�7}�/v��gmֳ�N���о���kq×���p��0�~롹�n6D��"�'n�t��ova�E\�ц�X�!�.\9w��� ݮ�;���y�Sϻ�2�S����tf6��{��U9�x�V��,��9�5��`هz��rcy�����CYX��/]ׄ\�c+0��L5r�Q���,�y��c+j��� $����)������g���*zX��d���-�g<����v#�ǖJ��_�<םσ��N2<����nM����g�9���}�bK��]�*�jO�{��~���GjIl[���z�ӱ�qͫ���
�=;Iw�˛U���ƾ';'������X�s��7���#wc��s����i>�#g���C�ӽ��ܵ��?>^�}�{��u��zI;��A����R�}�o�"z˛H���
ݪ��[��6����3���=�e������w>|���629��~�y��=�N�[.�~5rv���k��Oz�W]ཞ�v�ό�찤�c��={Ra�]�i�^�i��b����Ky�9�g^��Dِ^h��nZs�|\~�N�*�+;I���X[����0���ɟt�O �b�uvHo�Hnx��Ff�I��r�{I�6Ԙ �^��!�It��f8�����-q�O7��r�R��s�+�~YL��Ve{f� Л1�X�Eҥ�ա�_5o2�(��n�o�\S`j��bΨ�2b���	�hϝ˞� 9�Sd�]�Y��*eWP�#�{E��N�M���ձ	���> }���D������Y�G�����é��{��*gk���v�9���0�ѝ��k7S��3Q�ō\#�A$�r�=�>�y���������y�oq���v^	�2"=�y��ү�eC<�x�)�\�J/;�.�q{��i�����3���fs�=�"t�x�{=��kݾNe�5>���׊^v����g��`t�5�<��y�����(���tfz�y�sܩ�{�dy=p/'��{s�o��_y�L��0n��l�M��=bS؋r)+���/���G	��Y�h��xT�ſR6[��C������/�G�.x^.�]�<�I�Evh�P�G7��^p�s��U��a��K���Gʤ�NYW�%v��m���s�y�>�����3��s����ٖoϖz�'���|'ˏϲQ�Z%�em�m�� Kf��E��v!�h߽^�fߚ�7�ͤ�������R�X��P:�-S��h��,_dW�y:�.�6`Z�1e����ū�q��2�n
{��r�kg*�h��N7y�x7t��=���^r�e�V?����3�����q������϶�[r��2�d���_f���N��t0�ɬ��!-�,/��\�{>��գ���;���`ǹ���\��a;ն7v{+E�ڮ��k�y�-�)�B�!�[�ppߛ�ʛ������
ַ��״���m첳��ʯ�mp��T��u%�]�N}�&�u}�ld}��my�o^O��M곴|d�����R���6�6�29'�^���z����^S_i�7��og���Y֎����X	s���1�p�k}s����w�C<�Y��y;/ qܳ�tB�,Q�/}|��>9�5>FVo���w#|�E�g�Nwr㻓:݇�d �0����L��;�/՛��h�Lf_��G�C�\h{Lƥ��ד%�ՙu�;�CA�y�O���g�a-�{�{_o�v;�n���|��ҼVߙR�^�S;�W�7X�H�͵����+{+J����҄�� c���U���n�ӎ��K�~@	��E�Bۼ���i�\h\\���F1�OF�Я2��|�*c��m'��\Ph)��A^ʸ�8�T(��=J�`�:o޷�H��(s�� >ﶆ��9�w7�P�ݻc�:vJ�{�N�83��S�۩�X>�޳�^%�Nn:�_e7�ށ��m����wO���e̣Y�ω(������#Uu��L�s���5�hz@i�Á���ԾÎƏd�y����~wN/�Lt������e�f�����8����_���q�u'�[���i�BS��P���Lk�':��fz���[W5�6��62c���u����,�Qsa�ֻ��~��y[���c~�l��K�9~��/��=��z���=y�{�
^��%c�ཷ�ձ�c��m����^��n{��盅��9ҧ3�:,����,r=���X_m�b�3��t������z��=�����������>1��w�[,��l]g�u���l������|s�y&�A�ف��Ϟ��%�����b�Z$�wG��*n�5w�ݔXb�.nG�v�L�u��~Y�a�K(z������1���v�B�z�d�X9� J��xb�A�>�^�w��ŝ΋.��d��՗z�+'2EP�v�1�w:�s?e���{d;����N���Z�{��n��ϟ�|>6��欗�d��]]c�3~~s}��&o;�3{$g��j��J�Ĩo?'�k��Č�������9�'����������.K�7Ϯ+�sO1ꝺ�n��z}�B�Y�>#���?9��;��u��J�w}�����竣އ�٧�>�h~vB�k<k�Ӫ��}�����Xi+��_J�|�c���:|��j������&	N�_k<h'����2��{�z�>�E;3���'����H%�\��Jȃ�Wl�8*%v]Q��Ƒ���T�T;d����?qS�s�]Y���땤z����k����IX�P�I���(���'�]T7�J���~�L��a��KW��
�G����X죣��Ϲ�azP�u�Ƶ+���V����y�Ü��p�oCْ��E�?vRb��T��c��-���s��Uc���@3b�_?�L���ߤ��I�^�Ps��=��.����&�t�r�N���58�^���F�/�8�;���W���A��w�R��_� �'�xyך�0a�-�,�6u��l����a]�y{Tl��Y�t����X�/����y��|-��]-N�K���l���2�B��(��fu5ԋ3��Γ��Fn7cU��G'��}��o����2׶:Y'{}�)�m��N�,����
��[?W(rݟ����UtY�T����#k�%�v�8y��Y^q/7������E�nc3)�Ţ���g��~�O����@�u��9fN���&�ۗ�P�9W(Q�p��Zk��⿩��}�r�<Fo]�#�a���R�8t$��oW9�ZY~�W�ł���r�v��M�:&B�m(���Lj_4�Flo)�/�{*��i�,��<ޯ`����
'I��Ggȭ��z܉��<��c���(j�W��a�/b{N�Cmu�bm�v.�ݰ $���+����3���Fz����^�oN�~O��v����Y��r�����گ锌�%�Q� $�]�B�K�/�ds־��<�J���T�@����uc�_���qߧ��Y�=l��&C�"M8���Z��g����u<��J�lC�)��ފ^y���*b���xT2�G�}�B������uՁA�D[]����߱�-�z{�E�z`~�+�� r���',�;���n�[�/�nb��o�5��,�J���];���@��+2����ӏ�aL��j�#��w@��*�@�
'��kJ;�5]fR�4��Z��
vf�=,E*6�Y�S��%e˝��Z��j�+���ۃ%a��z��W�_}^��f�ro�U��� gא>�����
�u�oa�/U�L�↮L���z��K���������J���V��m�g�O�����R�:�D�K:�T��Ӟܱ�o�ڬ�<��}N�~��o{IQiz���l�����ͯ�Ѕq�X���Qn��
ڤ������n�y7����Jֻ��@�î�M��c���}�l3����\�*�R�b`�ι�^�=�>T�r������jh<뱦^�b�ۖ=��9�-�~��3W�]��,���}���;�\��Rơ��wǵ�A�m�q`�3�:���Gp�[�log/�t˓_l���������k��>'N�c�k�Ԉ睓	>i����z�x��r�N���Qb�)�3�7�4�j�z�Ei�t���8��<�H�zY?%�M�(%)��{�޻a��=�w��jZ�p���(C�$�R��ܵ�4қ�r@��R�f���]sy�gv|b2�����{]��)�L�zU#ƍq��c] �he�W��[G��<��j����t3\�� ���'�M�(�&,��K���t��u�J�s������&+�ʼ��w�~��P�Gz�w��X���k6V+א�i�K ԥ)a��4���<w�[=���빋6�5����G���}O�>}�g4�;;�_ >�ەݻ['�ݏ~w1���x�=�Hy�bμ�ެ��L�x�D��J#�Y-1����nwa����4b3,.�%��M^�Zִ��'<�/	�e���� ��~�͚���sȑ�z(�3Լ��3@�<78�mި�K�x��v:��vew���)����������S���vZJ�JE�t�uP�z�-���Ň�8����!ϷjLT0.��_�s�:J^7P��`�/猓K��l��G���m���.��tBBO:�O�Oq/p�ӟ5�=��[�k�[D���O���'��g���1"�+3�(S�:�����f<=���1�i��\�+�� (�\�.�O�,_�}�]����4���l�<��V����}gG�G:�'
�-{i�i�,+��Ϣ�ή�O���
hܩ�Vɴ�=d�z����X��h�2����O	���@}�^!�({|�4�J�]�.[~�7���;�2����#Fv;ӧR�/��<l�|�_��[E��'��}�]dx�SM9G(l���q�ݷOJ�䑱]��ؖ���2T`*)u�)��	�WY�N�v��-��-�=�w���¶��i�'n�x��@	M�^;]�8d%ff��H󻕐�m�>`֝O>�l�_��k'��$�
�X��{��U3������yY��Վose�8�>Z2V��}6֫�V�q`��,�/��P�s�K�)W�t���:Ձ�����
߲q7ʯ��i�q�nN�{½h��������9X������ʗ���ԝ7ƭ�>�)����N�(|�<pz
ù�|^
�����Is>�/Җ-�+[|˹�b�C����/�bV<��7ӱl�P�����s阎�vk�����_��Yכn?^�0�P</�$�r$V�M��g�M^�J+{�L^�̐Xf�����C��ɿ/2�����n�5�H��āfh�vf|���>O��kZ���=�<sT11M��Y�ko������V���쓣k� N~���[�̱޶�ɷӟ(�o1��>��mOW�������a���g�R�|p�:���R���z�mġ�gQ/K�z��i[~];�Zޡ̻�z}[Z|"���p��&6It��9�m���$��u�o�50{藏���ř�0Q�\A����P�C�2�À?Fp���5fvݧ������Qp^��ڽ}XC�-Q���8�̻j	Xf]�i�w}2���Uۏ
���UԻr�#uZ:��Q�t���R/�]K�,��Anv�Ζ�@���t`���<��#��[P��n$��u��]��L� �z���Սyx�3l�j�'nY�&{v7�F�- �������W�{K~�ٯ�� �4�)u�7@�cK ��i�/*9(_
�9�Ly�����:$�:Z����,#�͞�6*�{Yx�ESNW^Tю}ڕ�n��r{�X�-<��;0�ՙ�p�ӥ������|<^�� �����tB���1ry�Bs�;tR=��t��ͪ�����x�gݍ����vdy8\�n���U+��9�����G�7zą;�H�j�=�����Z��0�\�� |�e*[\P�f��G�3^�L�F�uH��4*ԧ�����Q}K�Hc����Mf�S���,Fr���ܾ��'%��j �»�*��ʎ�Uc�˛�
��b�UG���
ͽU۶��[�kwu�!E-�6 ��/]�7����ֻ�Lzuq�J@o���K��8�<WD�Y`���H,�C����%�e79T�bP����.����癮�`HmCwVAЄF�H�6�g�e�To�c쾪�F�7m��%ig^� �]����`���m̶�eg.����"h9v�o$waO���3���U��@�m����}��}��ڽ��jW'�}5�-���M6��]lZ�wKܟ�"� 9I.S�M��W�4Mk9�qENoM!���;��'`��fh�I���z9�۽ʩ�/��e��U��$>�7.�u}�>T�Ձ7YU�M��t��%�i3}1��֢1�p�(ts�7a��ė��{OT���X��:���kJ���֭�de�	��ns�)�v�wo�K��r	�� �h��)��.����Ka��zC΢�ku0����Q�xksHx�F�P�2�
{�Eݓe�p�hν��Z��4Q����xO�2��`i�K�Z��|�_U�N�G�yҫU��*�+-j�x©����,ޛ�����ȝu5S6�d����}����r<�]>��r��x��\�aF.�<\��l������hb�sa�ւ�sՈ4�Hm/�����vw���̮�i�>v�4l����A7�pp�e�#�0y,7��E0��[z�8�����d��m%����}����e�I� �p5Zv���-���dt�_$4]P�p:f�;zZ�31=��PI.R/{ЌK6O�X�}�
�t*�!;@���+v�V8�Mf��e���mަ�X��,Å��ԎӾ�Cu�c��&���2�D�1D�}'�R7)�fҖݎ��.�aF���b�1g3:�p�Rp�q���j֦����:kU�J��V��%���W�خ-5qɶ��nkx���s;�4(��,D�A��ڊ*�*1,F"����eT�V8j�*1U����
��*�"�qE���PDX)��Qb��m�UUU""�-d�"�JT�*�AAB�Ab�*�eeb�"��E�1�"�J[(�S��PQqh*�bD�h�Dk*ֶ�a,U�L%-
ZTFԲ�TŬb�����b�1@R(6�DQQqJ�V����&-W�h���kYD��[T"���SEQU�����m���\*�,�`��`�V-AB�b2�QPQH��m+m
�UZ�-���`�5�DEKF�\$���[
F!Z6�Z�[e� �֍����Z��\7�(�`(�ŭaa[n�
T�J&-T J�G�3W�*V��K��g8o5p-��.u
f�֤u�1l�cn1��R�T���R9�)�s�q��s.>r�5�����}�ח�}��m|t0;>����f���}����P�I��O��q�;�-z)��r��7���m����l�)��폅���z=e�lw�(e:�5��P��<RfǮ���` {��6�{�k�<j�U�GʥϓInx�ʩ��z�ǧ��j��q��e�쏝���H��󰫽�QM�k^	�`��m;߱[W�!��*9Y�ݵH�:�Z������r�f)�8<��pzK���x���b%f�JK|d^u�(��b����s�i���w���Lnc3;�����1���*<+a�*��=�%U&��LW��}%�K�ŉ2҃�C�Ѐ�"�]L�ӝ��9sW���{�]�!��t�>��jcv�k{=��1:Z�
�7
������넛tL�d�Q_�NBcR���u�3�p(���E�޺Y''4.����Ps�\kЮ.�Qo�w"Gb6���.u�zLw�O��~u�9�Ó�i�%�aQ5�Z�ilS ���e;L�w.a�[�F�yخ���I7�J�����`a)�s�o.,�3�i��{�����j�p+�6û�|*sh-�؁��B7��oRj�aw��Y�;��ո�gŜ���^}�Zw�k��Wʒέ/o��v�Ԧ�D��=��i���9�X������ >�:ޏ�K������)�ya�~�<s�Pv��q� E�0h%��P��H�q���{4���o:ѣ>}-��{c��#[��d��L�ne\�$�c�����r:w�o�ǧX�!Cb���a��\f��/<��
ŠISze��וg��t]��Ԛ����M䷺��(%D}a5΢�_��}�/O`���2`~]�.#K����%������>]qۘ�L�o��p=�QэD��D���vbÀoK���7�Է����"=�=�{θ7����t|���sm���B�^U/UpϤR�U��Ms�@6��=�W�O7�c�'�����6�I��O��X����x�K���.;XG�BN����CjL{��喜	���(�x�|f'�t����� ��,�[��B�^�ޣѵ��LM��K�����&���y�_3�����K&W�*<o���;
�~��Ϻ:���y9T�f
�u+�P�U@w��A�v:,�`�|�r:�|K$�+��c2�*�x��WJ~�(��!�zx���a�F���s�Vt�/ޮ��%=��$D&��h��݋�Cem%���mU�v�I��sM�(�:��b����	�땷`CM��ڌ.n<������1�V>��<4i"�i��r�Ӌq���UU� ������"����=ӭ*��d�":<�BO�fw����tr��kմ/�i��Ϲ�m3����
�Q_�i��z�ʭ3�vq#��T��՞�q�<g�zM'�n�s�'�2��gz(�:NvL'LZ髃&W���W'38�*�f��ޔ{ڌ��I�5�fo�b2�i�v��*5�)�v�AJ��S�19fg��[���)#�~n����ڼY��0�O7�Yv�epr�x'�2�'n�{H��Q-}�[&��쫭<>���,w(��������5��C���{���;���I�-u�O�g���5�- g�(���cY��צ�r=Q����~!�X���קϹ[+�yl�p+o�� �e{k���t�I5������5�D�,�8�����C}�a=G�9r)o�7e�:��.(F�%���B���Z�/n��+���5������]�{S�#/�P��	V�6২���uD3c���ў@_@�y�H١6V�]�N�ۋr�6��e��<e��r*��)ђ�WCS��|�nbU�^n V:���ݯ+)���Vվբ�q2B�9]�6�*�$!�E)�qoK�2��Sǫ���S��.6Ւ��c:X�r��ۡ,���Ȓ;�:�� ��Iӯ���}U�LFU����V+�\����d�&������`��
z�J'��Di4�tw�7w|�s_���m;՛��k�G%��ϫq�K>���-��:�O�sv?=����K.�����i=��*e�Э���%�������౸<�4����u^��{g��q�x�������oF&�~?m��<�y�sU�kզD_ݖ'=�NU�n9��֝v[����6F�����>ZJ�;��ǒ�ڙF5D)�w�s��P2���=��q��_��Oe�Rf��y;��@��xW�aTV/Z�S%iˮ��;����s��uL���Y��)���NX���Xw �dhtp/6�t�-Y�����+�g]d�F�C���Cl�Z^h�8M�a���8V���Bn}3���L��%"7�Vh{�9���t�q�eU	uTF����>�j��E<�Z��͍���[��T�:��l�s|� ���ݣ_k�_ǋ�~����;���<���k~j8 ���tS9{י�5,�Z ��`�<�GN��r���^|&*l��W�j�Q��{����b^��7�c�+�r�MA+62^��I�&W&VpsU�>�5:.� �x2�r5�'�m��qؚ�Z*�8�+lI�o���m��w�ӗ���Kz�Y��B���/r�=��=����7k�,��h��;�\�'�/hS2�z�S&�#M#���<]\����{�Q��<s���	��&U�G/�j$�E�Ipۑ�*�$䮰�����f"x{���B6�`�j�Z|"���p�	�-G�j��/%��x�;��DWe��ߠ��]�����q{��Z�&
2+�>]��8*(C�2���ܿlB���;�=�!C���p��cs�\�I6�,7|�tym�=��ژL�5�r��yf�{���h�٨
�
A�gZIx��T%���۽}��n��W_x9z�M<��p1��Z��ty^�Co)b�:��п*"��D���Ə�tfu��qcZ���<��ѷ��w�f���zkM�̬����G�h��:U�5��>WӶ����U�ձ���ᶙ��fܸf|�Vt����C|�:�Κб��1Ғ�t���s�g]'�yg����ņ�ޱ��n�89jm�3�;�����z�B<�X�,�"����u��<���Q��c���wUɋ��yu�,�֭V�2�G6Zys��N��k��d�fkN�7�K,���Y���Mn�xx규V���&^�Lr�Z�&ބJ����M��mRf�'l�"��N�|�wTh>v+��S�MP��]�����k��~ɞ|n����ST$���
��5Qw��qX�.�t���"�W��%��yi��b�Ԙt���OV��Uq�(�ʄ��Kew����OO{����7�����#w�?g9Ub�\BvG�A���nǾS�-��>�LR�CMy+��%�z�+���v|7��9�k|'�bY����;A��>������V9*��͡���7�A��!�{��+���>���J��2�i E��0I�Sl�E��x[%o�>FS��ξ�}���/�(�D��قL��	�g0OY0���H4��<ӏY~�F��=��$�0ܰ�5_��lC���`���~���d�1r��[�����1*��\Y��$c��}^p8UppJJ#�kUs�{�r^���3�,>��i�7��+o��Щ^�dN߹��H�w,�?T7��IWJE�`�\EXAyQȟ��1a��.��oL�P����ޙ.��\`}w��tH�l8��]��l�C���r��"�j�sS��R��)vƟ��Z��\�x���]b��o�F-f��S@`�;{w�0β���~z%�Nk��{O��t�h�w6��zw����2�{/fn0_�c{����0��:ڒ�vЙ�J\$�ω}[�t	[3��]v��x�0�-��R���ʞ� ����{�Q^n�_�f4M��2M��|�P���Åi�P�]��ɢ����͏=�4 �������{�ό�Pw�t"|=a3|�_[�^l[��[�|�t��_�W-����!~��s�'ƞ�Mzּ�u/����k��ޮ����r<�����0+7���C���x'��,�U�y*����=�"�n�E����P��?Pgq�z�vg�7��:<��v:�F
�}��Q0w�\�+��]��G<�BM��2���tSk�3{sk5�{�B�^� �f���}Yj+i��/Z��V�����N$z;��=�D��g˓� =�9�k���{�k�Ea�k�`�:b���d���g�J�U���g��=�G��\���֌bzƑG�ܽ�Tk>�H��%�<H0&6�Y`�.�#k��g3?Q"��jU���j�f{�v"(<��gT�W���O�l� {�Aʖ�E30߲v`8L"!���R�2j�֙���.Nr´k£`#㶘�I�s���uo8��n0��e�����Y�54z���*�Vg(����*�	����* 	��er�5>WNw���N�>Fzگ�л����'��Ξ�]Ս�b.���b�֛4���%�a��L�e��"�O%9u�Om��<\���>�fE�uި����T6;)�(����e��6;>�6��K�Z�L�re�uv��W��a������Z�v����t^�ҍv}ѐ��K��Üo�#ʻz.π�#A,�C\��5���%�Zw�W@4t��*s�B}��yh��E�yG�qwzbۇ}w��d�fW�#8:�4N�২�Fx:���Mz*yc7
̞�6�*�d���A[Uex:��tMS�5J��m�X6�,,���� ��XSQ>��΁�z��5xD���\/��z^E�ո�k�5,఼��>��9Z���P��A;dy~��\�AP/��6U�~6���<=�[�6W�n
���+{��9�k�o<��W�G,g�-�L8Ms?m�уΧ�9��9~�2"�����Z�ܝK��O}ݻt�M�F��Ǡg��>XߑA<ڊF5DL�eu�����gf����q��,rq,ܶf
s0�t;�c���ѓ���G��aTH���̦<{v�`��VuvV�P�b#��j).֣�,�FC�'52���I�}׿؃R}h�|i�P}��m�n� IXaR�,�Nٗ��8�i"V��;�ѭ�o�mc�.=W�(j���0삎�����W���]�K��.�P�Bי������}�S��y�r�C��=\��)��l3,S����Ŀ(2lz:(������߀7\�hL/��D���a����T]J����:1Lm����8귐��Л���-�^{+Ӕ�=w2q�fn񰺎��{Ǣ!t�CW*�s�:㬤�0xmyv�C{ۼE7y�l��Oy��+���"ݚn�z�b�+����ٗ ����g�l�����ɝ��,K��p!��Ζ%���<5� W_6h/��Jɖ�f>���θ�����~ڮ�����Z����x�Y�.��͆
ժ�
?^��Z;�w$'k{&����g�x��}q(^��v�b?)�9����p�OY?"HGd���9W'^d{�T�T��^�9_o[�Ө��%�<$��?Ev�8*(C�jݷ�d����Y��M�@;W��_�ј!�ϮS6}�X_�uÛ��%�J�+�N��?yԗ���Y�x|��/qc��:ѳ���*T)�σ��K�[��s�v+(p��5��m5���	��8����/�[�D-)hW�	�ԐHSVo��ӯ;�=U�N�+�Z.4��+�6�� �W�~�{�i��h�͞��7êYl�N'�,���v�c�锣/M1j1��{;������=��n�n�ަ��V�ݣ�J�i��u���~�h6�cZ��Q�{����r�hN�yQ��\���I�7���)x䇣b�Ѿ[܌C�X�0��Ρ$_�e�+�V���X���z$uUY�z����][^�jF���=Ő�"i���?���0'�8<��s�{)�����9n�7y��[�#�l�S����;$az��YuQ֊�����f��k�K���u�,a�/sD��+���A�q�]�~�כ~9�G��'��6�(��$�C�t����;�i}7�.az��v<C��ͅ�Z<zU%��-^@]l^ :���<����j*=\2b�{�^̏]�Ӗ�<���U�NpY*!;!9.9ﾂ�t~lt����Ee���K�e����͍�=�c��g�9�8�ZnY�r�j� ����ވǺ��OE�,���o?rV�`w-��On�N��ռ�����C�I��:���0s'�v_a�/·��ֺ�AB����~w5{�6ǻάx�n?xzd��zz��zɆUV�2��)�\9�@䮫u�|�����uua����dYO]4�Y���V�����Gt����)1��o���VX�B�Dh2������r���)�:;8�\8����ݍ;u���=Z��[��s�Ο�^:yi�8���Ζ�vՎ�������,p��El��S��r����ۧ�-��G��l�I6��3e�7{-I6��w�]v��*�W���Ig2������".����t칯o��*�q�i
�HgvαSbR(+]���4���7��v���ا�&w����AC �|0J���Qm��g1\��h�2��u{�'p�-��).���R4��3u��f��nVj&	�pZPgB��Ka��k���J���@+R# ȡZ��])�Q����YY{ԗoZxw�A,��u���ln��>��Ou�\��m�u��n*	ђ��I�Ss�#����&���]���л��G�q��IHV"�!�{
N�;�2f��H�8S�+I�j��(f:��ũ�}};�=�s��vH��SZޤ+%rw�乮T��b	�Z�DÝ�&�rh�Ǌ�"/Q����������U��u�6�B�5�yG]f[�ty�r�"vˋ�J�[�Qא��-�S/C�R_.(��:��m�ilu6��S�FHI���O���Z�)���=������Wj�K*�]��[g=vų�}t�$Y��G�l9h	Ԙ��9ˡE��Z3cw;�2�s�W��	�"��n�k�O����=�3����t��(�ufl���gQI�`j#l,;��:��}Y:��&�5f��	C�P\y�S��SLܣ�\A&�>ߕ .�ӳl7Pᮕ�%}�˃��'c�ݵF3� )�5�e���~��#��y���������/��{�񥼺����煕7g�[밹�s�����+���|����H�٦�ѼB��������).��Uu��y*��)�XVsm���-nAؕ����*�i�ۣc���|���:��|m��\5�S��p�w�:�XGb�P�N�Ǽ�<�,�����\����I�Vk���'DK�'9��f�Ԛ�Lj�93�b:�l)y\�g��ѧd��t�D�rs�·)X�t�q��1J���Fǃ�;XJ�|��e���TAb�X\+l�x)vl�hd�n���sShoV�5���n���A�Y�@��X��9�P�6Z/G��5�if�����1�3�gF([j��Ҟ�y���Z��d�Ҽ3��d�i����Iw��"*,Ȧ���ޛ�;��J��\7�6i� Ю���G��}�;�������"2��������;4���s�:�b@���r��,شeEO�K.�Ž��� o)�W4�����=�!���f�m��k4�%)���#µ�l�nL����m`�� Lm����-���X��[q�"�Z�50�Z8j��cTJ	�PU��KJ�A��\a�)W���mkja�0�.��E����m�����V��b[Z�%[*"J���ih�1J�6�J��Ҵ*�P��D�-��ն�p\`��QR����l�UTm�Q�`T\4�ڍ)X�EVB��qp�n,���m
���1`*�f�T��4��UX�1L-�VҢ��P�V�U��f0���ň�V0TTmF��h�YXUaP�a�ֱER�-h҈ʅIY+e���iYkAJՖʢDaZ�Z�-�ł��m*�FAm��*U��Z+ �P��j��jڪ��Q
�e��[A�,FP[j�lTD�0�-��e���(�؂�E�-E���[h�3�����K�ھ��7y�iWN�.�w�� �C�[��`�g;l�}d⊬��k0�7�L�P;���B�k6N���w��O=��D�$��3��Ս�6/5�gI�Y�x����*b�V��mS1�p^{�6��l��V].`Do���R�8���r��Z���rd����<s_Q��"Vɺ��w>wQ���]�����ހ#���q�E��D?r~�f,0[iw����©K��w=��J�M����F�9G��yvz���w��5Y+\uT$�3c��{<�=��L��ۡ�qf��+\�Qfr#�ˀ|���:��m�5Ҷ�f�\R�=��@���;Ǝ������0cC�������#�bz�t����ۏ}���D曶7	~C��q����d���d�Z�y�{�|'[�N[K ���������{v���2_v'3�{O
R#gI�/).K�^��Qz��ݎ�9v=���*���ڗ5��s�_�t�q�y�3�7F���f̋i֕`c�k��R#�v!&}C]ep�U�Yӽ�OAN^���&r���Yj/����4Ui��='�qN��^Z�E����Ľ)�Y6u|��Q�wKzz���P������^�w�#=Ɣ��gg�ɳE�-oQs��8�d�|���Ac��תj�NW���;5�kv�ԉ.�P�)���r����j�Vl4��d�*Y�0v�6Q8��G���.�ڻ6B*���H��S����5��kX&T6���-t�W+�ד�3�f8=��sݚ�U��w6q�����o�����4��c�7��Ͻ��7U$f
�����z>�ɞ�px�Dv���`�xΜ,��;�{���N�x9L�W�d��/K�r�r�F��D��?1s�
�Ip,���4+Lz�t�$#~��2?n�Mo�N��w�	�#�)�(��S1�޽4;�����|,�I����f�O�=��3��_�jZ{�Tœ�Z49�-+�ywX�N:�G-�����C�{Q�a/T�q`������P��mʄ\�B[�I
Y�%�2��f���ủ�[��^��"|�yX���>u.M�>G#��f�	�秱�˙=[e�Y�}oOsj�C�`�x	�k��=kH�7�
V<�m�X7󂹁=�j��B��r��y���O�Yr��f������\\Uߜ��6�mk�5,బy�g��$x����^��{&f����C���W�tg����g��M�[Du�)t�j�����T����}'>��L�倸��{�/����r���ձe��;�д��,U6g"�I�>
�l���c�������(q���Q�q��%��t/1l畛��hg1�c�1�
�V1��E��L��w��0���U���m����|�sX=+�q�x�ۨ�j���>ʘ�W���)��Ѵn�1���r��{������b[�d{�kv�嚾�E��(�E��~��G�o3i���ݴ�B���R%���N]��:�08�>�:��
���`0�+�|dg(�׺1t���o=�얶ЊPig�f\9��S-f�f'S�%�gޕ�s����v��;K>o~I0�i�*�˥CH�b���ƌRM�a���9�|�&�o���r36�t}�k>s�=eq�.�p�Q�ʹ��y�:���8'+�m�-�B�ξ�Ϝ�ﯯ�f|�ȱ,��ݣ[ԋ��q Y�sa��V�[��Y��W�,���������Ι��<��}=l�0����C�v���C����B��pF^�QVF�u��[�|�We%p�i��Yܮy㜤Xt�zfq�O]��C�B�j%�Ȅ�A���7�n&⳹IAP���W�@ I��f6�����K���V^���h�����<��9�<
$f�vUx����ʍY&���e����tfN�k^��`{��QJ���gY�.�x-=/���l��R��6��(]�wr�������k��դ�I�:k��̗�ZP��i��t�5�L���֘a�G���O[�6���:T�i��#^~u��l�D�}K
Gb�۱9v�H�Ө���`�rVD5L�
���:��J}���Ȯ6uwr��Ơyvt��E��4_5o˃1A�U��&o�"w�yxQv�����A������֧f�u	Ώ.�,�2���/)�u0�"����H�M��-�����\_��{�l�[�N����X֥�Ҏ���R��S.����9�]q�+��h�}��s�j[{�mi�c�ȏ�P�5�'�BH}��.�8Skƚ�s�^������]P�sz�ͭάU=��cA��ھCmC��`�ݗ�18����ȇ�O��sZ/��R�31�~�U����RV���+�,q�n���0�f'R׎�\OV}����a}Y]��xe���;��=�0<5��U�Um���h\7
�<��L�ӗ&���VV���n��y�Z�ƙ�t�f�o�E��>3䖏G�ؼ sP�ײ����5�q9�OT��.�{��v����]�V��@����T
���>�٫�oS��YH��G}��N���������l���+E�_d
�����l�0oW7�]�H���KP8�Ygto�����=���������xEK�ɽ��1M����h���a�'��N����U�0X	�i9E�=�GO���3pe�]��u��+����m#�A�m#/���g=���a�8չ�p��S��a��㽺/|�e�H7�s��{�jeKP��5yM�G�:����䗇"JL�h:��Y��E��9{3u�M�o��I�N}B�vWt�sQ��|ܫE����d��zz��줊�u�M�}x�l>�'�`�4{�_yO̽ϐ��^�>^k�ϺL���+�xej��=6*�,7�5�,�vn^��F�]t��D*�#Ĵ��W¥���g�ʺm�&�eu���w]7�jx��݋��n}ź�;�g*WK������ґ~X*WW�P_yQ�)eD=C���;ڳV��Q{��_-3��HH��.�8�F�a�>W�˰�w�o���T�>���χL������B8�VOP㇚`oK��\�U�gyp��|ʯ]m�f���	�4��2���ڥ��ôx���jOh�/�kا�>2�����Z:_� Ts,S��IoW��(ǲ:O��BH���� ���)�L�bΥl#��ۘ.�5hŠ�e�ۺ7�l���n�נ=}��
�MI����&pfi���OS��4z�m�Ɇ�{[�u�c���0C��w؄Xkcs�DE��{�2V��7��[ݏ;���r��խw��f&	����J&Mu���#��Q�O���K�Wc�n����7��I���|�`��ӂ�������D�a.��m��7��� uC�����z/�����=2>�ܩ��/�}��3�e�A]+Vl�Ғ��g˖�0�������)����Œ`�֙�T��{�\���[��>�TLg�cQ���8���w��w����׺D*����ԡ"LK�_���<����:
ְ	�`ʾB֚����B�UP�+�u}�*��YC��{G���ds�u������r���p��x-W�*�����h�J�6dBH�.]����K ����	،7��<pL��T��.�qA%{�ۍ����G���ä�|�!���O{l����l:�镜([����+���/F{a�����y��g���6�@�J%�cYA2+s���:m<Ϳ�_��ƹ����o���>�������=S��eLY<(;-\���u��z^��6����+�B��\)���J�z{���	�9e�撕j�8��w���̡���r�@�uH��=��E�^�\1����Cswho	
�)������&�ݙY�����ԧ@����|���X,���ǈ���%}}\<�;'���|V6�r�*�=Rm�h6�L
�p����(e�>*s	����\�|}������)o��l7�o��5��y��懧�Pxt���s�>G0�ʢ!�5�ykrVu�{�=E����)�QT�����J��g�mi�ޘ)_�H��Y`�pS�Em ��K>��xS�wY��7@a%����<����=i��u�$�W���E9�}����&���%����41bϻ�L~�1���/��L9yL����C7:���l,n�}��N��uꓫi���r�/�n��{�+-b5ҏ��R�cҮ> ���Oh�Ow]�u��z<}��0_^��e�̒���q�3��|�야�Ou֬թ\X."�^Z��������<�ދĎS.Ec�j�{S�=�fe9�w�;P�{��VOk���["�)��r{��o�;��>.�J[hZ�"��ٗ�p�ZͰ�N�(K�0�N�gǖJ���<������`<7�c>���O�b�_S1+�Y��F.uC�[�}x}��=�~`�b��U<P���q�zQ�ۣ�3����#�EГ�u���Ex�f��)�ݧ�FZ�*�㚽�D/��()�N�jCv��q+��7;.��mb��jm�8hv	��3���5�6j`�S�z�4Z1�ob:�)�=��3Ah+S��KG�6ۑ��C�B��t�4O�C��<E�Ė�J��c��+>�j������hY7�1�ɝ^]��֩��<^ ��f�XdX�hk�Z���b�\\YA3,we�e�{���M�����U;�<B)�skb���=�<s�z��b�]"J������˩��Řt�4Ow��I3^g���e���Ln�̫;���F��������`8t���w͵B��OvUV�X���U�
9䥕:��_I�gIc_�S3Ǽ�LZ|"��.�=:�^(a�6��;�ΖP=A�(�-(Uҍu��Go�NE�}&
6�dUʼ7y�v���KMo��{ټ�l��r�����+�"�[G�y��pb��ﻬś��%��<#��IG�����{�m�q
ٚh����N�uP��>�V�*81վ~��%����L�ϻ=�6A��ޕ�L��W�
Ė6$�kR�åW���/�9�C�O(�C%�۪E�we��qF�߾���C�;o">C�k�J��p�/�2ޕ��/,���WRQ�u����,Bp[�\u���s����[���ܓ�=�Gu]���۩�����6%�9��k��r���ujҗMЁ�{Րf����J��^�-��,�ʧt�u]�7{�(��TmG�Cm�2S��Q�G�l9���=��bk7;��桯��n��T���/��5������ݗ�0⳧�x�����<w=s}Q�ֵ5�'�l�ힱ�=��3K��ȯ���ؠcrٙN�'j��9�_��ʘ�Նw����Sw��΋w��c`0]�Lt�,gҩ/%���aA�|�Q.#�M�Vy9���3*g�z������������^1�u�:�VP^��Y�I`|bKG��V��%��]g��s����?k�^�>��9	�-��3cZ�m
�uW�y)
��R�/F��W���6����q�;܉�(O,�H�~��r!�Ys�w,�a�֨�$�L��QN#�+5f��xfs�f�����3�}���n���U��������_�X���s/����\����㮛m���>4��`4����(s��֙������:��V4�s���	�s�#���ml�}�?M��>�7���`v&�:D����Pq^�����v���)y���^����l�\gy���:��}&B!㾽�<*e#��&���GR����s��|�������I=im:���\��ܨn�Hm����v{���~gwur�W���lV�ǥ-+f�;|��]���M�c �Knn��j���6N�5B�e$z�FEQ[(��u���]�4��^�[
��t��^�ncU8:��Y����d��}�uu�=]��y����Z3���'�Cbe$�t�_�T�"���Ku���^�r�y�{˧���N%�����+���y��H�\G�yve$��
yf��w�=�ŮU^�}���1"Ua��\=�C>��@���%Zf4M�2M��O�<�(n��;o\�3�\~j���8V�Jt3wב���ׅ�{�N-*���<G��s�申Ĝ~��0]<�J�MZ�pƁ�>�¶�d�Z�y�_3��cP$�XJCz;$�^��N<�];v������yDk���mvd׵�A\�7�[z���K$�j��M5]�|��o�@���qt�>A�RV=\����7[�q�|3��=m�Kfsn��N^	��^� �z�+��SV/Z�*��=�)�Ħ����fl��w��*@vq#��?K�:��]G�Ύ����L��J3�������y�uޠ��')P�>���4�y��o��F_�֭��9�n8�!/�;;��%�aWBԦ�.LzX��n��wzy{g���מm�_ո�p�Y�A�_rp�ڳq�Wm7��.������t�ǃ9��ww�Cn����*�)��`&�PT�l�l�i|�Ӣ��.�B2��k�M��0�|��}a���aj�����>�.3֪p���5IDh�9�u�T�v'	�ɚrP >�7ib2C���1U;��;�[����<+�?Z;���;0�qC��u�Ok~b,�л�A�e�R�IO^�9��"���z�+Ǆ'K��՗8�t�9���k"����lr��W ��n>�R�2��V4�zc��S�5��}�n�ۊz�ix`\U1�E�v�V�,�kGN�=f��oM:��{��&<6�J�if;�I��\�f�i�&XF��bo��;ϰ
Ži�-����F������y`Z�{o;�39S��G��϶�O���ٌd����\6Ԃ�7׃����2�:̝��aQ����⠙��B*���]�OD���,�BWb�u%d��p����y/�:|ٕ�W�L�x��u�j4���(k�"��u��m���D�M���N>�_�8φ��.��X��[uoN�����{6��kw��-��c��ɂ_:\�VV'Q]e3���z=��W+��5�wŢ�ݹ|�j[w����ލ
S{s>�3k�����(��*+*�վ���塺�(3Km짎+�ﮭ�IGs�sڽ�E]h����P6���n_:ڍ�畜�U�z�[�J��k�|y�����P�a�'%�U�&�a�l����-�����E�{G@c���ac5��wi���p��������QC�HY�	I�(u���Yd��6��Z��o�H�ak�W��81�H-��T�h�eM��6�q���I4^Va�9�{�ǐ�v��;�PEJ�A��훰�J4z���:n4J4�,��1�K��&��j�=v���Z�"Z
��&�����[84��QIiǶ�0Wt%�*lPp�3�(�\9,��N���"�̠WW+�ޗS�nR䫷���b
T���F\�k���7�vS2��MwU�詭l>S�v8ַ�F4�ݻ�֩bt�H�x���>/��ǎ����ܛ�\�D�6��d��.�+�Sdzs�d�U�J�E&�[�k7:>��y�
�e�^B��s�f ���J�Y�|��:�$*hw��s��ʹȁ6!S�ʘ��YxK,��ئ��؉�lY]d�R��ض��j�n�F�.���������Sy���X4[�b���1P�O@{��U�Vu&p7�K:1c�z����#hgC��.��W}�iQ��"��Y�m#�]��%H�a'�bR����A�{K�����N�ӭ�+�4#��tz���`��#�n����Nju)m�M��~޹���R���dW�"���l�V+��6�@b�V����b*��%�ka�Uk[F��2���X%�PPZ�ADX���ԣR�UVQ�V�U(�mYTj-h�j��l��QH�+cZ,EUQ�lmZ�("��c-�J�\P�T(�TmmUJ�Timkmb[JѶ�+hڋQ�Vҵ(��[b�F��j[,Jմ��hҢ��#"�2ڥ�B�"UE-KcjT��*҅`ڕ��mUJ��Z�*1"���U��*ֶ�Z�cU�D�Yakb�j4ZT�B�$XE�j�p�1KmJ�RZXT��)J0R�Z"���
U*Q%L"����,*��UJ��X���V)j�2Ҫ
6��Q��D��V��(��b�F�V�-,J��E���-�������TZ��UA0[
[-�V�J6-j�6�-��4j0�miimP�����M��1�6�A�rU6�e:x�wQ�!O9�[���<`2����f�יFq��r�pӛ]7,�.�Q:g	�w��Y��X����v�C���"���^��̑[��]�Ϻ�4�W�3}��F�{�0���v��M�~�n����eNf�r�;,�q�S1��2����(ؽ9���iAg���:��-��<��8��o�xTr�%l3�.��AV�>%�\=�*<)}�C���m�*ydO%ޣ�m>�Oթ֟5L��Y�b���b�3�J��Fh-�G�/c*�X}��*��I����>5>�L��'Z�[Q�.�p�q���g�*,!�Hz�K7�F5^qn�ܫ�7ڍ�SW��|.����B�^Vk�3>��
� gz�i���ac�f"�X�3A\S+ӝ�w�F5O��7
����Gp�=�g�����b�y䊎Ee��o��E��ڟ������t�E����%��|���:�G[����wd"���`w��?y�r��mwt���[�,(;^p�0Ϸ��c�B
���/Я՟{)���C5�����(zٽ����:V�cd7�Ɨ�ȵ.��Kɏ�VZ�k����r��eܭbU�� �٪aR��֝Pv�ƄO�L�X@��t�^sWyOy쮠aii�L�n%��E^���\E�w���sut v���<��m��]X�h�=���n���c��X0j�t1�	�c�Yq�*���.��&�R����jq��W:���7��Z�-L��]��<�2�z9������	�ՃV�q�"�G�&�wW��{��TP�*{��Y`�>��X7-���>���g�����p���^f�~^���콧C�di��<SG�/��Ͻk�f];���rǏn�%$�B����{���E��?"��2�"�1C�����ъ,q]D�ѷ�,������O=uZ`�wB��^����ZG�`���Ih�$�]�WLV�[���ze>�9�uv�Ԟ}��<�`�,2,	f�ۻZ�$X�\\X(&f����%��Ý�on���/��؄O�&�����<:�4����p���8��.qY�X[�}�3��T����Q��L��iL�p�8��;��Ǿj5���w�&WY�B���ˌl��ӯ�����+�ĬRq<�P���ġ�6ZhgIc_�®.���x���{\�{��v�1m�v���`
9�t��uϛ���ƤNu�:Ll9Yj��b��޿eu?}<�j�8�)�@ݴ�e���ʘ���1�so�[|�
��a�-\vZ��Aq�ap�s#ɪ�`����J0�V�B���s{�����'Q4IS �kS�ʷ��)���M�ܷ�*g(�-H#K�Z�l� ]Y�����9�Ǽ�N�Vx4!���f��C�l$p�4���s����㷫��^�rG����IF�V�`�Z��'M�&]��,S�"�|Y��*zFY⎊�����qI��Z�ϓ;jޗI_�\�a�"�������.�|@#��v�����9h�}����&r�\���|�ष�t=����UX��;��P�5̷�{�o,�:�}�7�(ggx\��丠ÀYC}Y6���/��R/޼0u���gN8�������u���������ܼrݚlՙ���f
�5eG�a�`�r���o�w1wjOj/nj{�-tm�3��r��֮���?u8�*�Ľ���d+��`�u�Y|��^��N=~�=�
��n���ơ��2�#��Y��,�K�I����۱X����V�W����]�f�%°zQ��@�2��\���tZ	���=��U�4��4�^�3ρ�w��nߦgx��By`ia�w��	C�ßN5ܰL4&��w~�#;:��!i�E��yӘ�9�Ӽ��o&��%� }�F�skp����K����
c4������ҥ0��*�u���c��|����f܆K1�M�s%�e�G�>�ː�!ס�>��3ekn@xa��y�*�����y#q�B�԰{��I�g]˚���#�(�ek������*�����Y�!�C�f>��۹�#WT�� 5�I�2�w�֙t�yw�mî*#���a;뮻����佫�o������h~�`x9���t�?q}�(8�}����T�&y%>���*��K��9*ooZ�
�ܝ����C�'�Cba�k�&���GR����C�^V��\�%�T���j��}�������5C���kF|���lL��t�_�T�"�s��s�Y�j�v���>�fE��j�ޗI/��탎Q#Aq^��y�z�L��q�t��
���;�.���,V/�V��2�ަtr�1g�z]�Y(�9���x]��d��5�,�x�q��I]�kB���hq���g�Z|+R{G��x������s�F�2X"�cR/L��]��d�+���X�e:�z�o�u�KO�m$ɮ��!I��๡=S7FL���s����y���P����O��G��/ᄹ���d����W*0�v�vC©f�]�%0�"�i�@�wD�m?4no3�E (��������^���h�N��z��\��r���ۻ�[x�E����=ʻroJg�b	�X�ܵ+M���{y;c#��c���y��fgC�t3Gmd��:b��{K�ҝ���]��*L��uJ�;��n=�<`�.͖�%cО8
j*����צz��罧	�H����Kt�ϩ��=�rޯ�����;�VZ���)���^w�|s�o˝�E�y�.-���ԉ0�I�\"�Nv���`^��3�]��4�	�g����7������J������K@��N�e�X������wn�-�g��ۘv��IRyd���-�'(1�����~�v;:�4�j�fo�b0�_=ߜ*׺�we��=i�Seq�&Z<lK4Mf�Öc�?X�Q�-���5>o�gOI��G~=Ӛ� ��L��)��<��L��VӍ{ �hp��O���w2f)�|�W#�s���p�^����~S�,�2�,�����ΑiNg�s]�Vʧ��eF�N��9p}w�_m�]�޲v,�R��EvΘe-�ʄ\�B\��|�����mdˌ�HO��y+��/�.����A�Ȼ�=��Ȭ��UȖ�ȯpw�/���~i�7�����ʅv\�Wn ��In�����lD3G�L\��i�>k��ǽ�p�7M��ذ��G�bs��0�'Sn&N\|2���p7q<���ѥP���7�+_K��@��U��Hu
g �x�ׅv�fG���pl�e�;��4X~�`u�\��[d�ӏ�B�{��D��-��0R��>�o�����{��0o
�I�'ڬ�f�#��i��c5�֘(�^��W���E{����Ui󛺻��J7�c�c"�ά��ojdYz��j����f�>��l��=�N;�v񞾯Z`�Ҵ���*�zt5WEq�K�v�_�y�머+������X���9���+�d�'5}88�	������u������ϯ�2�|=��rV��^D��VQ�4���ݵ�U��r���樅3�J�5e�=�ğ�rى˳��w�~����('�״����Ov�^�}��{����ǔ"z,)B�Ю_O'�X)���1:����8���Gz����9�z�;��^_���Zj�[j`�51�a������+H�R�<�Dѓ�M�>��|��yʇ>�/��N4=��'@�:����������HWV�.ø��]��v��'��QX�}��<�l,��wkU���b���>yhBC��,U~#��<�K���x$��Q����=a2bڑ�O*�^�$���ͻ�ն�ÿ��(����i&^)-����ӊ�:׸���%���kםJ�(VWV:�y�%ss���������qk�{!�Kb��������TݮB�[�jt�=׆�e�/b�\"$J�hn��_<��zs�<�q�j�|(K���9�ۄiŕg�>��>j5�����e����ќ�3���3y�]?S�A�X)6�(S=}�C�e��t�O��*���� {�k�i�uҏ[��S{Z0v^�����H�t����������S�j�;i��}}����uc��^��������{�Y�P�<��
�
�Z<3�G���p��f�k;�A�ß�m��k�)+r�
ę�Qk�|哦��w�^S+PpBuW�Ꮪ%���G�m���ر;1��|���>�T�k+��p7�u��
�Z����p_E=ὧ�]u���i~�� �k�qT�ЪK}g�*n9���x�\�U��$��̷�{�ҷ��-v/-�>���������v�e�uN�4׀�6ԋ�7���8��ϼ��qq���v_���,�=u�ځ����죧�Y�W�̩c�����5LCb�7-��~��l׍m�!���pPP�Y�ngwt��Ç��9�M1=��d�q:��P$��|�@��%�E\��8����vv�={ֲ�{�y��b��&�L�p!;z|�u(��G�s--/B�X�9�Օ����@�nP���.�^-�=��-�������|\OVz;�mJÇg�x;И�Ic>�xa.��R�u��+�I���{�2V��z_�-j��r�Ft픓�9����j�D��hS��̗���M�RD�S��w��g��Ke`�3��\���4=ɛil�'dp&.�q�N�u�;̽����y�r
U�S�/C��#�`�<��g?N�9�C�Âq��a��r�����u�����:�|��D�J��%�4W���g�sW�ۄ{�l�k瞽��{����Y;����C���N���#/�h�	sS
�/�3�;w5x)���cH�����I]�(K��ܧ�ۏ�<��g��������4M}Α&���Р⿷�l3����8����f�y���N����(T_p��9Sdˆ�}<*#�&���du+��w6���Gs�K�������m�>��Y��3�J�a�T<Xr�����o�2�Uґ~\�W�����fw9G�7;m��/RVYb������t��/>]�s�(���Q�a�nY�l��f����xx�c4qT�o}z�1���!V�w�dߧx�������-�e��|8�ٷ1)n}�nn5x5���+e��\	�q��I�G%��˶���Ʋ(�.�Ҧ6�Y{]�(V+��e�,T����J�B��o��t���z�K���I�xBL��v],^�Mׄ��\3NC����@��1�\	�d;Vk7ݴ�ߩ)�.}�Gw�FT��hB��Ƈ��ei𭤶�5Z��./�
>k*����Nl�8}�:A~����Z��f+Z�b`��|�i𭤙5֫^B:�D*n�����tL�c�u[��N�x�[s=n��X[�Tp]�#]���˪��^��uͥ�1�ְ`눃6�tY�9�W_lsД��<��{nq�"��
�&8�+�ˎc�����,V�����ۖ�ޖMv�����N�L��X�\����+Ρ�Yj/eQ��Nn�]�G_�{�T�Բ��vʿ��=�8���c�D9�'�.��gGAZ��vw�b��ͻ�4�+-y	��u(�<.�<l�M+��֌bzƘo�	�������{Kz�N��}c���8.\�G��5���"9�.�`�x�����h*�U��ql�Jw�.��n��ׂ� �^p�/>�h�,�49҄?����4kG3��`�F/I�om{cڗ��%񜊌�[�7�ﶺ�9'+�j:�w2U�"�Wr�:�(bdt~��A�F�w��x���v��'f�}��c��������dLM�u��8v6z�Z�ഡ2�3�oMwyʊ�R��u�B7z�\�}�&�3���z��Z��M���zz�x&`�X�i�wH�D�U3��"�rfo�O�X(�ó��>�m?}R�ֽS/� -��^�192�,�����}n�^���̘���  �o�w�6��jv.��S.���|���*F)��k�6�{*���V���H
�u���`p���� ��]��tf}+/>���d�9���Q�ur�ޞ~Oו��,_�!\tW���-ӌ�n�¶��W���%�?9�X3k+<�G���Ɣ{��e��n�{�9�=�i�aH��������W���<_fw�s�9�^���o}\��,jY��}��'�0p�7��c��
���.b�}��jv'�VාI�͎���{�!{�{��Ҵ�pP��9�,�ҽ ��z���ǂ�ٞ�ݍ�je{K�2��1��O����K���L/�������e���K�7<�2�G1�ђ��l^��NN�!�`�;s4z���~��]��#ʾ��_��VX#ڜK�\d�3�Ga���|�Bzu5����X�X|_ 2]��7s�vX�T�<����w;߃��?Z���"a�>�*��=�h��%9[��K7R�g3�!���l�1tu��h�k̺D���I�X���sÑT���ļN����&Wb���z�l���GV��-�a��򃲊]f�Ǽqs��PI^'��Tf9A+��9�iN�ǏX�JtYA�����E.9]��e��Q���)�E���|��m�.�y�	L���,�Yǘn���-ݜ����Q"ҜwE��X�捥F�ƕ�W��IQ�w��;x�r�Zll��j��T�Æ�њ7��\�4l�`�n��ܫ8y޹z�u�U���h�m��t��ͩ��x�l��o�𼻄2(V�3eh4�NE�Y�W�B2�qu_Z�ս��r>gC�!�i�3l'�y�����}���ut�\ˤ�v�k�a��o6w�f�ե�0��n�umgd�������ȕX���uQ����s8(T!��jH��M���;v�Z�<�T�ۛWcn5�ᩜ��t�j��R�D<��9l�ˁ]<@S�͖�K��d;����2ۭ�Z���v����夫8���B!h�: �O�η35��i��:�Z+�n
,l޶YVG�D�zD�.$�t�I	F��	c�Xf��W���z�魳IW5{��HE��4�lK\4B�Ζ��{7���̫�s���!={��ٷ���DP{$�ȉݤ��'�uʺ�TJ���ߜ��;�`��/�-�n��+x�Kz�����v�\��?/��^������2<`�3T����F��o�4�z������eZ9��6h%0P����ں��ਖ਼�tn�ܺ@�*|�)J�����)�2'Ո�/��f*�l��Mc���ew��)��r��Ev�|8.��j���s�e˘Uoir��t^�wg��vs���_
�K��j�p�pm�_2�ldǬ���(֍���D�)RaUy@�VĽ�.N�΋�qj�ԑV�w�J�[��0&�ۻu�lV�ׯv,*4m��($n��ݔ5�ѦgعR�Ц�]MLU�d&��$��Y\��1t=�ê�к7jf��p
i�y�##ܡ2����-���gb�����c[�q�QP���E-�H�Ǵ����D��u�J��{��y�wW^4%���)�U0K�Q�3C��98m%��:rS\W�1����oΗǷL��W�C5�i��������r��-��	|�*E�;��e���v����H��&��c�L�넢�\?d��>K�fv�[]6 �эQ{}`��v��50;z��y),�x�Gjq�Gh�ծ������SQ{�3��V��ҵFo%�έ�t���Z<��U��R��j�Y��zk'!թ��/�[� �yB�
թ#���{J�i�������x��r�ѷ�}�m� �G�E�e��Ѵ��b�-B�kTX5j �X�Q��Q��TKb���V��jQVTih�X�QYmj�Ѵ*Kl����jEJ*����)*#�EE�T�-d�ERԲ�B��R�R�cU�im�U[m�X�k(,�j%-����R��-�h�V�jR�e������Lc�)Q)[V���QR���qV�h����kiq�8,���Ɩű����VV�����҈�4�L&-+-��Z�	S���KlkJ�R�J�8�\Z#�[YEb�&-X�b�b�1ZRՖ�Ƣ(�Kj#�kb֖�V���YDmFԠ[T���YY0���ŭ����Ѡ��1�FЭYh���*�֪یK�c
(�E��h�1��,���F�ն�b�[j"*ҥ�h�--�.)��cZT�*�0��B�)U*U�D���"/'m\�k�sr���WN����j
<]Ү��oqx��i�$x_�&A��"��'|(
�����v"[o��Ys��3�g�>��eH��8�Ȥ�XOе4+�����S-f�fsu�P�
�_wN���{�kG���]��q��J243�xz%��bƪ5B����ʢ/qML]vt�no��?k�֨�0�:���_4=8���I�DP-�#�:G�e$�z�BX��ܼ�{��=����2��Ϣ���Q\�옼a�`���f�ۻZ��ԋ���3N*�k:<5ӎ��(��T[�=����:`��9��潋�]�'�������m�n��d��-K����&f�rQ��0)�þo4�������rD���"�2�.���{֠ChB4��hS=ި�<&�M%�~S3ǯ=�SԁU&"�ck����I��A/`�\w׸'��l$���Rqu��|�v���/���ә�~��9�d���:wJ�>�Y�w��z�g�	B�TaxR;�dv$Y�u���U���K�ίY�3���pIf,�邒�%Bɘ�q������ѿ��� S�;�5�GF��N���AX)+�W,#�;�v��z�	q�k=�>�g'l6���F����;u���d̩�wz��!����[�.a>��7�D���'7X�������n"yc�R��w[k�q�gpY(���q�٣ا4=�1�MV�dkn��<���[��z�wk��{:t[������^��W|%�f��]%zయ�,0nJƵ.��v��7%���3mX�r���˴�m�(�߂�߬�Ϧ�E�yހ|� ��z>�Nc^�^J���"��^y����mFp8J��#�R��6
z=���nv_�.*>>[��K����E�m�O'6�w���9m6'nTP�n�_J�Qb�5nXdW݆탃�ؠ1n�����3{:�$�y�=V��x�u�9���F�\��a����Um���J�]�ӧ6�b�&���5�j,�C��9��Kz�ju��1��~qz%��F/�Otg���=����7.Y4;2M��%��ъ�1�E�k�zy΋A;"��>5�P�p��׋��i]�N���B�\�/��#�`�<�m#,?N�9�C��8�Դ�4:i�����KOӴO�P��@l|���*��ﮝ�p;�5x6�	?m�qZ�6kV��\A�y�}v����yH�v��5�\��J�o8���?a��}��X��溳�\��^y���pn���O��7|t�=n�f.ً�*�����ʠ�0�=�b��egX���ZD�
v��%�e��:���t��:���s��튏\�� ͒�^6w9��AE�t�\W�f砋����n<�M����]1-=�J˯99#|}� ���a��&��H���B��������>�GڭdoR���u'�ꝃg���A�*�9Sg��9��lL4�t�ҿ��I�l�����ݮ��{�;��=��Z���Y��]�Q���',¡�����#3��{wk���3�٘x��Ե`���XX�>�,��7��V��Ev�q<�V�36뭏v����u{�~HGO�h^�@xK-��u�5�u��,F���h��3N��Sٸ�]_>��{�K���v�ڐ�"��V4<k}��Z|)'��%k�G��`֬�X�۞��o��`���h���,�"���!���wʳ�gZ���&��9�n�>Qt|3���o.�ǢƠ:|�4����e�;x��-�;>��=����!�:��b��H��p�ɫ=~�&OU��^B ��c��s0o�uJ�;��[�i�^�W����h�ݲ�^��w�����<뗢3�^X���"_= J�i������z�.�c<�m#WԸ�-֖���ݭ�7�@�%^V����*���� ݷ7;p�:�tq�X�����nP�;��,��8$��,^��>&�&�Pvb|�k���T�Vs�l t�̵�ъc-h�f��dG��oPf$�"uդB�t��4N�o�ԚeKh4\=\��+琩��h��]dV)z��]|V&��4�G<�H�K�_���Q���y�fW��K�m�Y�tѶ��z��������!kMlԚ(l��4ҿ��C7�N�a�Bh.�Lۇ3׵�y��:N��]�>Re#ҩ>ZjO�#��r�v}��XfQ��έ�߶<�=m�����#��x,�[�\�^	��E�(��!ŧg�ؾT��������٦!_��ɪ�_�!O���yN(�^Y룧�� ���5ΔK���|+���3��5��>��y Ynq�3�Aͧ�\:ׅL�-��^���Y�2�,�.%�Ǹ%��ں��ʝ�"|��t��o�y�@���d�Y�mF��\.�}�k���d�}�eG]��;p��5�J�@Ҭ�ZK�r�����4��5���%a��[��+����{ʼ{�|���]��f��B_
�+��m���s3O�@�*	b��a�;De5���m
[��Q�5e�a�OR����Es���2��9���gD�w֐�c�Ww^�b�9VE���47�~�oa�oW>��g��3�9����BV7��`�O��ih;��K�=��_�EOwj=��nޫ��܋,z����݊�
����}�9Ey̜�ӳ��,�w]��`(��Aer�|�@�pۇ�'�4�3/�vD�d�=����4䱩f�,+��c,�o�0�7��|`�9��󤵆�G��';����	k-q����]�z���"��cpy�i�^^
��/}u}��kO�7���X��}'#]���k��U�¦�m��ȏ]a�%��y�e���|���o�Z��>Y�|�nh�]����K��	��_]ȯ�j��������m���"1yk^�8m�.o�sB�չ:��
���a髋)m�Z�`�Q�~�L��`ޞ����ןq96{G���qCऱ�zu���/���G�ҡ�U��R��]1C�RC�%�%�UX��ʝ�ZS]��&�0�s���C�q��ɘ����m&�<}�9K5�J7�w2�Ǟ�1v�B���p��E5zu(��\��0�Y�Pf��¬sgD7_o:9\ǧ�[N_M����#�8���e�/]�~@��=PæOs����^��.�­��P�̹.��o[�c����z�_bi@LP��L��[Jdۄi����u���j�b�0#Jз<�����Z�$��W�Nf�F�˩�ne�~ҏ\�kw�7f��8ߧ�������$Oe���ՙr*N�'L�'b��t�@�A�H�1�x�&�����.�C9K�̢��8(u]_����EjX|�v� U�<�_HL�ٽ!���Qo[DO:��Q$y���_z�P��-40t�5�Pug�����J{�v}*x��5�8&\;�z�dQ$^�\R..�������X�<zݜ*�����q��8�Q�%dA�T��8*��>ٗf���4#�_;.�fp��M�*���q*ܿY>�o�_���
IP�bL�(���tؙw?R��,�W��9t�z�﬑��˿m��nx��q�P���J��మK�䷥[v���}[����cy�u(�� ��v���Q�;��V���v�4}�P�5�%_��H�L�3oo����N3.���l{���kB�`LY�{Do���x*���*�Q�EM�w`�꺻qv�N���t���}2���:��;ݔt������K��Ȯ�v�ۨ�n{˻�������p���2��Z|\OVz;�mJÆaX6�Bc�XϢ^My���v���o=�!�0Ѐ�m�L�r퓮���]�df�Vn��2���������\�9�.�.е*Rk��&�{N���S�R-5���`���}X^��M���˩�"�]!���]�S��Q�*�≅�5�p�n��/��Xڙ��՗�*���] ��]�r�����J�:N��U�|��ty��SXN��s����-\���5	9Ȗ�ƌS�� r���fƵ��A�u����+�ڠ�������K�AN��WR��܉`�<�m���]eW��k�ݩ�\�ulZ-�s�}��$�b�D5nhrr���^��i�w.j��m�=��ِz�����h���ހ߹{����]�~��ok�E������w�֙�n�c�(�3��;ȹ���M/#��t�U�"���a�*bɕ�����4O4�8Gօm�q>I�w+/v�I���D�O
��)y�(V-r�.�}=��;��H��I�����WJ���'�|E҄i���g�}e���貦L�+��(���	�`P��{6F=-��&\f�^�G1/&EJ�t��SzYk�t����Wl��$h5��g��g�9+��1:��s�ν���ր8:�>��yh����
E.��8=��Ek�J��3�ɂ�����=��>�����קն͚�[K,�?:��爱�m�k׵�Q %����#�NV1��״�Har�[}�O�g�h�՞dk���2zr��J��
�r+:)β��ݸ飯��ol��o��_i�^�s���ig
b��Y�������s�x���4�rw���Qۃd�+�K8=�Kugt�ˣ��0��lo�F�bz�Gh����9�6�u�xd�.�V�ڗ�{5d�>���o|�gq9����[���ܱ�|�M�<崳���r��N�X�-S�1Ε�l&ū�<7U��~VH�}�J��ݙ�"�
s0o��ZY����{nq�$ST�ʰ�+k��/O9u��ޙ<����֓^*}���*Dq֘Icn��)Շ��� �z�t>TE�l�9�d�ΏIĦ���~������8���R%�����m+�y�
�����^s]�u�>�V��eC�+-rJ��>�CeT��i�c�T1Ջn��^�qS[�#��ꝵ8��r|T��R=`K�x�ZjO��"�����MU>C%;y&�Ʌx����� n_5�B/�K��`LN�����0�UZG���ֵʹ�i��Aַed3׾o��
5>H��u�E�5�L�B������e˱ִ?fú@����u�m_g�%�5����k��R�+��6Aͧ���~!�W��,��|s�l�ޠ���;�2�f̋��\�yn�Cn ��[޻�ڷ���zOJ��X�<R@����ǉ�]6��)��X�M\C�F�Ky�^o!a��Nd�ޥ�XؖJ�P摝PH�T[%e��܁��]u�:tG:���(l3Ԝ2�=���-�zf�/��à�}�Hį�����h�w���mF��\/�]��+w�7����V�������V���������4���_˖�8߆�)��oj��!���|����~n�/���<} j�Q8ا����Bp]�����D�^E�גͿjn�c/y�tF�s+��Y`�
z����E4k��E{�\/
^��{Żs2�vwc~�q��y���zX԰k����谳�>�鱹��ayݕ�u��X({:���qi��Z|�}�l{ۘ̾�Z����_�౹��ƖJ�\��ڰ�*gy]�^��T4�&�m��pz�!1}��Mx̺g�9��8/צDT:���ݺk��c�ʆ�������4xx�8r��a���ݡ�Hf܋�U��N%�L�ks������������Q
=3���oشZ�eTH��НW��fTWI�j?D��U.t���z�3�}�eӹ�.����m��t�Q�����=),g��D����`ߍ�� ���Ѽ���t��l>��ί˒�u'�G�Z��s2IamH�0m���(��Wt^E2�� ���M1��(SY���3�7i����H��~��4��t��{}�.�,�&�ۮ�r��K0��]�}]�R�wWsjE�wfDy�Ҝ�ɞK��Y7�9�R��8����8h����x�U]Z��8���3h,��g7��c��HV�o�/�j�J)��1w�͂�"QCvCQ�5N�oi��4��G��fD�fh�v^ ���~�6�(x؞�����(c�ۗ�{�^���N���C��@֦���e�
f^SJX�t�Zm����{q���F�·�y'���;m�8{6�NG�x��!�t!}��J�s]�)���ġ�6Zh\���聽���c����8���T���E�2�L�Y$�5�⮓��>����Uy���V���35o�7��m�$�gI������z�g�Bl˳	��x//����{�6���Bx��m0�^~X��^�d��JD�yxQ�38��9D���.�j�I9�z�Mt��9���V�*01��?{۞,��(XޗIX��%�X֠�o��n'o��$���we�����j��>U.&8)-����ժ�y�s	P|�J��^��6=����Nu�Uy��B:�]�|ڮ\��Dgcѵu|�ayG`��bne���{ұ.ұT�N;]�^�賨�r`y��i�{}�,�Wjb޻�/)�6.w�3�51�ԫ6��`��[37���k�B���m�:���*� �ˍ�r�]�`/mLN�~���K5lVq}�;y@�v��r�ɨ[\��"����nw*OOQ�ڨ��|�;4tw0��V9l�м�e��+ܳ��Z�W
R��*����E<��=y��h��X�<�Wv�a9�������º��V$2�6�&WK���vƻ1���gns��f;d˗�;S^dM���U����#	��<4��;�Wc�8ӯ��X��L>�1��Z�s{V$[L�EU�y�]ϺwGݗ�����Cw�)T���eҲ�蓇P7�K͔o��\����"�^�
1>U9�� Lj(�Z[m��:�M��Iw:zA��!�8�Z��FW�����k�`x�,{i��ˍ��1�\�����tJ:��E�Q,�J���v�vh��Q��a��r��Zo\�>V+�:*U�[$Ò�B�:B��%:ܽ$c[��މ� n�~��#��݊�r�&Gl(���E��訹P�ӹڋaҒ�Xd^!����Թ%^e�O��8��Ǎ�I�N�L���/y!�݆��r��f�tQ�ћH&/{o/����U��H��K�4����k�p����h��׬W����K��u����wj�lm;�<0��a;�r
<1�l_���̫��A��Hj�l��/m`m�����)nu��ȤI�'	uh6d�8�;CU�8I�����oC�<�t��tڵ4R��vf���i� �m��X��+aJ����7�����P�`i9��Q{t���ux)�=q����Qa�;��r5[VVm`\�-9Bh���Ai�8�~ ������(�q{s��⳰�;`�It+.�^��ۺ޾=��G�P'W���P�؆B2�
�Lꫨ��	.�W��Ր�8՛[/T���D�"#�KW��jc�w�|2M2��cs�;��9�|�k���פ�b��%sB����b�{^
����K�w�h���yi���By\��:�r'@���r�<��x-��n�N��N�\�NȨ^�-�S
�ZM���Z���kj�k�W��aU�!�4.��oH������t�m��ƎYz;��mS�X	��R�b-Z^�����^����'i��:�KAr�TOt΍���Z7(	uW,�vN9t�攩r"va:�3�n�)n�G��[�c�q�F��5�h��`Q,�`�4E>F:���Ӵn�f��MD��(蕗ڄv��bUv������w�aB�Ȋx�}���NRjwS羣]��O`�8-�7J��&.����h`��ht�=��sR������Չga;J�ŀ.��{�E�
j����������2Rpo5�}�o;�?O�ƶ��1h*�DF�KamKj�-���[j�%��*�[V"����Q(�RѢ��1�Z$�ER��-I��D����Ab�P����j�+�J��Zҋ-KZ������%Q%TZՈ�[U\S�E
Q�j�B����K-�X�R��-e�+U-,iEF�Z�8ËG	Q�E,aPT�iZ��m�֖"����Z�!me���Պ�,h֭�.���ZZ
[b[
�Z؊�j����8h����m��R�U�,m�YlZ)F%��J����QPF�cZU��kA[E�IR�R�$R�E����QJ�V�VUEQ����R�ň�F֫KZQ�(Q[E
�Q��*���l��h�Pm��b"�*Ub0j4kUKP��Xʉem���m(����ؤ�kUk*V�JUcR�Q�'�B?f�˼qؚ���Y[fp5��v���j�hIU̇;XW�pr�BԎ"�嵣��QפU̧���ŭVQ'GW�~B��zo����G��^�;)��Tք'��	�k=�/h��=�E�7�?s���*-���<މ�o�p�vT�"���l/v;���-��	��%~2R�.��5�^.�{0�:��D���#ܘ�n[3)�ŧ����GP�T�8^�{�Yim((�lk�M�ե��!p|�YPخ�Te��d8�S���t���5�e�G�&��s�&�Y���:�V�_�+�|�32�C��$��:�l�tb��!���q��B3�38C����{2]�zq�@�'���+���)W�\�-�H�������_����%qBЖ�so}7������Y��>Xj��A.I�`%�L��Ϯ��qܹ��)��'�Y�f�v���)勵s�w�Q�6�{������e#��P�`�\�ϨP�e��y_����&�׉{���uS��l��*Ƒrs���z\��O[9��L70�49�$�#��C'��i��m�{�����l6&/Eڧ�I�Y�x��"�~N)ks��8'�Cba�F�ojw�@,�E��*mӃ.�E�aa)G�OV�Z�S:�(6pN1`⪠ܚ ,�!N^y��HXTWCK�����P&E>a���]@���<��Z`�X��k�u$�p�J���pe�ڵV�M��룮��(q�:�5���������Ve{r1b�����Ũ̄��0��*��J�"��9�x>��g�A��*d��"�9�mh�,NO����y�u�>���]�v=W&��n���N�3����:Yk�.�����]�k`�����_������~�H�{���;.Ç ��Cs�-<��tN��Z�h�=�a<����T�o,����y/=�8��Z^�[	�w�O��bvR��·��}���Z|)'����)G��oW*nVo�{��bqiV6\��f'�G��[^�QZ�|��gZ�97:��+��d��9߳SBO<������=5�c�[K�)�����L7��I�{��E̩q�}I��׶�b�=Й�SC`?vd����3�}Nf�^K���_Z���&T87'�3R��H�>���`��-+F;'��߼�$�ۦf
r�@�?/��:� ��}NogT���j��3Ŋ�K���jeK�e0k�Ӊ�y��,��A����3��gl/}�{ޏ]��.��gz�g�����p*����EVz|ߨh�ǉ��|;Ziրb�k"n��T������g�sWޮ�Q9�V�S�1`�d�n�3ܽ�NW��U��ٗC��#Z�Q�۽�,��]h�͓޾a�Wෳb��I�.�.Ųoge�W�cFERr:\^*j���z�g<�S%;MpV��*�=A��̜�>.'�{��3��FX���	��/ ��jZO-.�9E���5�f�N,����7�W��{�v��i��\Ɩ�0�M�ay�b̙[ޯ8i��e��ĳD���Do;=��.�Ɇ�CӮ�� �..����Qk�?&��/��y�^�˗c�o�ƙ�}:��*7ow���q��R�I3�	�[�l<t�~.k¦_� [���=S�E��������z[��Pw�c��5ґi]:���z�l�d�XmF��\-���3�AR&G&�_���g�Ԙ1�B/還�������-r��{����C���ү(�k%�r��zߨ�u�O2��u�O����bDC���Wy"�m�H�X�5i����|��ڬmA%q��+��$TpEe�a�ORϺY;aY�͎VEs���,��<��^���r��L߽��4��A��,jX5�aX��τXYՃ��oj�D��k�Ǟ>���t�{�׍�Ls�~I���Z����X����~��*���ŕ��l2m� ���\�[��w�����bp" ��|և�Nt{�������F(��׫h+��Zzr1)[[�2���ME�����ժ��H��F>���j֠�e݌�;]bR��g_@�m���JEӸ���J�L���e�mN����س6y�!����X�h��WK�ǥ�����~�2#���U�3�8C����V7�͔'�7����]=�Z��U}F52�j���'��^��Y��/��+��>�g�|���
߲q6�wms]��q�ݓ�+�=�G���	T �q�D�OU�g����)��l3/�w9B\�������^_�VZ<��,g�ׯg�]��)�kq���X�� �(K����ъ,�n#s���CӍnL�x�Ն��uz\b_Q��4�\���:��dx�^���m��}��:�W<�&/33ԫ� Gim���mu�=��m��*�ו�HϏ�L��v^v�/)�W}<o��y㛮��D���g���9���P�v��D�H�(����U�~#���t�Zm�֥��=��ww���Z����3�L�k��ChF�p\�ח�<�|�v�����������cg���=�b�衾GˇpOY,�$��qWI��W�7Y�'*XJ
�;��*�{���y$�Ո9�r�^�cA&�mY���a���۶�o��ʂt���W�1^cp�u�I�%Y��vvc�ʬn��I*&�c��W��i:α3f4�eA��>��y�N������{pu)ކ�^�u�:L\W}����<0J�̻0��O��������<9���"�>��šй�ﻬŘ7�
J�B�&c��Y:E�yu�Ny�w����=3}K�gڀ�#�?wy,v|tc>�|�Z࠶K���.�.��З�;�Zx�~�o` {��5�޳\�!�2�1Wµ��J�!��zx\o�݃~�C���=���o���đ�u�*t�3+ҩ�O�0Mg����o�
v�\�r�ܨg��U,�Þsm������H����#�zz������g]��c���ΰ�k�C���!�b]�:w�{��D��j���0S��n��{��j�zi��S�u���Y�������U����O=�g�K�	u8P��h0o:�Qe2WNfC�[���]�da6=��J����wi��v}|�>�%��Ė����/ �qY�F+NBarޮ��H�\v�fn�V�����K$LBvB
��2�����T^�w"G6
�&�3�K�(�/�k$��L����
Ūv��pQį��12]�\�ޫ�*��+;2J�XL3z���#��swwgUZN�}�D%Hm¢��l4j����Nèn5t�4�\ƙ⶞�So���i��9>��v[�4��[ͳ�+�� dc��:�.�u[BE���r�R��Y�w,�L4:¢4�\���h����3���K3�
��aLx|�U������<�#}�O^W�a��<�ȃ��)���"����50P�����I�e�:���V���[�:ו��]�{p늇��$��a����xO[92��YD��H����i�kǴ�X��N�o���V@�������/5ڧ�I�_�R��?�_��Z���	�P���8m.�mNu�o=q�у�K�X�du/���9����Z���X*d����Ϝ�kB����aǀ6O{�wIOG�VK�p"E�Qq�L�ڬ�)ҋV^��H8�k�/��!���7��o:�`ޢF�m��]���i&lpS�E�7~��f�����j�2�j;�i�lܣܵ>�J�ŴM�)�lt�}<���*�A��m&V�
��qF3�	-�,����z��Zq8���plyǈᘞ+�ȫV��`��jW�e��)�_�XԞX_Y�R�·�5-k�GSܣ������==l�mC������F�%�00��L�3���Wgw�pKK+3���W,J�H�	�Ji�]tͫG��퓮����
�MEvk�N�gV�Z�g>�������H{�̢f��aי[���Д�3�j��SC�����Iu�DI6�h��6�.uu�qҘyw0�{3�'3��߲T7��f@}{\D�c��Nf�uE�Os��+��<'+机J���{u[���6�xث
�͖�M�g>\����jDp;�	;I�������#�3\��
�ߵc�Ϲ�"������Z��#�����L�|V&YN$_����E1�m��Ի1�m�{�;Ƽ���y��^�'<��%�Z���PB�������D_B������є��4��)�������Oo�y��L�z��h����M�.y/=��w�zW���.]��oY�ř��v#��x,�+{��2�閏E�᭗i7뺑�\�z�����s�"�x����F���T����Q�,����j&��7�T�\���&��U�h+�|KJ�PL��4��9�Ԩ|ө�����Ѐ^�{ ���rޮ�3M1�+qv&��4�KB�.���K�o�_p�>���Ґ>��<�9:�ȸ�Pj�L#�I�k����S~�qޚ��S�w��_��ٹ��HJ`ӹ;1��W���-S�1�+��@�&Y�εT8W}��C��5b��7ѡ�':f�Ћ��:l�@����	�{QA;&�s����5Fy����h��^�|Ok� �Y���w�P��A��ay;��<rf_IXay[Dゟ#�v�Q��	�,p��E���.��#�����`䞜����G�L�-n��Ϸ�
^w"��+,~K~�d퀬�f�A�zp��LɽY��6sm;՛�������Z�v!�zXԵ�Ac���g����Q�ک�����ݻ�˼|=�������T3�0Qν�&O�Ό�G���;�ެ��x�����=����>;'=Y1�VZ�k��ҿ�+��S��.}�]�������KƷ��s������v�͑��2���ڞJ�X'���}e���1��kTD�q?e8����x)x��_(�oގ߹>K.�\�3�KhZ�v�nE�vO<��=�Gȥ�#��Ξ�	�x�[n?^�}�" �ˀ�������N��brǎzu��]p�Q�����<���-{ס^��9���R�ȱ\(u�C�:1E6ч�.uC���CӍnL�x���RK�(�
�W��OI�oN��`�2,��3��T�Z>�j�J+�}�������y}q��-=�'���V�ʇ�X�8��16q.�C��>�b��؂�$}*����o.�R|H�&n��c�Z�u�(�X��A݋�:'K���=�l�&Nƺ�Z��V*�v��h}i�	%{��kr����P�s;&Tms�J�^[x%���ZE�����f^;��;���'�sjt܃u�D���˒_��=��9>~�ױx��X%K��J�S-�ܦ������Bm#W]���◕�s�sm9���j����>9�+n� Ak5�\�`�L�軹ˮ�����sBr�0�;
�O{i��U��
���(o�Ϧ\;2�dQ$n�\U�x`�/o����k���Ws뱱v�u�:Ll9Yp�?.��Vxg҄;s.�2��ћ�S�
�|}ދ&[d�tԅ���ԧ��1A׺ǌ���H��T!\��kG��|q��W{إ����6�c��+-;�
b�pbo��U߷<^�;j��+�\����0/n��]�y�s�թx7GU�˸q�����C�9�&8*�߬��������Ƃ�v�W(7��1*��Sp݅2�N݊§���er8ww�_
WאOz�#�կ����Y�,��7�P�_xe�t��E�^[M�^�w!����w�|R�=�T �l,���M�E��K�V��x���vg�*9���Ў���w�#n��1���V갵j��JS8E����{�h�s�)w�pE$R�+��ܹ�>�W���7�lZ�%���R��iz�+�f�̮/(����3��ա�n�|H�8.�w:��:�a�=b�j�>��֠��f`�s��z��Gp��Xp���ۏƈ�[��J�x���z�����6��B�a������
d8�S�����ޅW���I̒�����Z͜X���}I���g�%���Ih������7�D�Vyъ�S��=UZ3�n4����ɴ�~��y{�Ƶ��A�P:�/%"\���\^}r���ȑ͂��2LY]�W��j�=nW���H��s��C���
�:X��SoSn�ނ1��ɮS�$��.�	tv������>���>Sn
���}��i����t�/�*�_ވ��H��`�K��Y�;=����N�%��=�4]O��p;�5x)���J��X����d��&W�zɆ��h���7oZ\��=��뼸@by�U�//����v����Լ�+�*b�~I��f�,ԩs��/mܾ����V@�_U�>%�\+Q��_�~Gv����g�υL�5C�˘�H
�^{5;�̵a��>~̤�t�_�
��U�3Z��)�Yk��H�����Y/«Fs����%���b�_DUu�n��k:rb>�2$�bTʘ��R��	Ƈ���
�#�d�a<t�&�HNh]Y�E6qw� �6Vv�v%+�}֐��}|:�J���5^>�ŵ+�^�}�!�[��Xz����$��-2v�DrSopS�*PB���|�^	L�ג��݊�i���N�|b�HĎ޴� lї�;�p���ݶ�k�� v^�ʦ�����p(;u�vT��Ҩ9ڈ}�ºp
�`�ۀ�&�묔�����&!�r(m-ͦ7d��ڹ'�;7iJ�*�w%GLk|(�������N,��� KO44l�3o�Jڏ��'3!�Z���lD�;k �f�\3x����ۖ���6j	��Ϭ�`c�䷪+�Z��ٸx�9��f
8��x�����Fܰ�Y��qQ�#9�}�Y��3CD
�iރ�m���]�G-`�Dqlo�ͭ4); U�[l�;r�3�S�!�㛥�pGF�X�
w2�#�>C�'x�f&�u�D	�AՕ{1��x�7{ԆK�Y����y�ҹ�9|�5��m5P�ă��w)9�s�k_
�[�M�u:½YH��4�s3�F^^����%`�7G�p�wv��q�a[O3h򸞌yu�z�o)Y$�뇛�,�K���|��֞�͖[��*��|�K�ӭ��aN�Lq#�7CG+zr�ˠ\���\nm7x�S�Vn����:�Aqm�2Vt�)�M4i�c gT�T;�e���ܛ���O8.��Ӫ�T��9�9ECjW4��'8�
�O��+�;�Y��K�=�'kw��*ulג��� ���u�9c���NN�m�٭�YZ��4�t�)�f����u�F�w���1����*�j�0����e�jWB9A�c,m��}O~}�Le�ra�_�����^3ֆP�ȹ٩���hc�v������u�E�5�2��8�j�)Җʾ�X6E���N�BvnM���搸^�B1�7��g8�z�Z�%r|������,��ac�xp�K�y��@��,�ߚ:���Z�����Y���n�P��t	Z�BaEuf��eWb����茮Ό�P\�c�X�w/ �<�w�b�(��{�Mu��M��-v�,o]��X�ˢE���AEN^ͥ�����M�s�U$��an�u=apղ��ՋV��ə�I�3�)�k�j�o5%��9b��}\�t��o)S���Vhv��f�^�ۄaҴ�y1Rf�wS��O�QXdS������Sܝ�S� ��;��Uea�����f󉵹���Z2���F�夹��r �b���Aѩ]�ȋ�JvL�N��ֲM����y�[�^�z��[�cd��Gl��$ ��V��EC��mU����V)u��˻h�b���L�:�����CMVF�U�r{i̺x�ꂱi�{��uu5��n��ۻ����[h�)[EQT*����E�eE�Kkh)X�U,�#X��[��,�*1X�mR��Z،�Z�`����D+m��R�h�*TEQDjRڍJڕ�--��V�ҩmX�U(�m��QQ�j� �TeQEj��1e�A�X��TU+X�mmZʋm���-���j�ڭ
�ԥl+R�6��Q�"�Ѷ�F#iV����+T���(�lEFڱF�J��Ek(�eJ4EUVE+,QEF*��B����"�R����F%B�ƕ�eB���ZX�J��*�U����	iT��ѵ��1TQT�jYKJ��5(���ZUeB�E���h�lEX�1��%m%)VT�� ��+-X��D*�R���Q�F�ڨ�UkZ�ڋ(�m�-���Q�����Ұ�������""�Q5�Q-�PPm��������m�Em
�F�V҈�-m��J���1+X��"ETEQ�����Ҋ��1��Kh(���:�'͙���}��n��ix����+�,Lzҽ�^Z��t+�!a5��U�`-m1��Q�F5�i�n�}��x���7ܸ��Wz葠��7]��m�O��o���*�H��f�/q;]/xO\����/T�.���a*�1�o�2M��O��X��zא|�.X����F�ԫ�X-�ly�i�>���׵�S�8��]�Q����D��^�YKV׬��w�b��h�T��,��|β7َ���jL�����!�nX�X�M��ize3�¡�����6(���qk��Zx�JZ�}UڳT:����]�{��� �6�tX?O�����-ȏc�	h�ރ��k���E�⚧	QD�>��b�){e��R#����Nm�3޻]i������͛��йoW��8����e���^�l�/=����ĉ�Ϟ�ޙy=�r<����c�% ��"�s�O�=�w��k �P�VZ�,-4�GRh��9JF#��%D�=�AW/��8�=~SУ.zƘp:��^|jr�2��h񰴯P�>w��N�n,I�ga�f
`�V���cK ����֌.{�9��Y����z24�� qE�ݑ�E�z_�b/�B�g�m������ﴐ߾߽�>�7�T�4&SAW�TU�ɤؗ�L2:�h��8�˯����π>�zѿ_��웫z=Y-��P�����b�έ��J�l��^�Y�1�DFqEb"��K�^w��6C�2��Ө�����G3�as<��ߊ���X����ԃ���W�N���A��.{�"yg����(�}���q���GD�P��|:R�$�kh&Enq���si��íz�_����Us�η���{[����]�qm�f<��>�����t�I5�p���%�Q>�{�۪qX�N� �29�N��0{��;.*��|�Z�s���������:�/.��EÞ��'��t��V���wh3$�2�k�3%a��Um�OQ�0�ʢ!vJÅw�G�SàтC%��ƞ��޿e����/�ݞ�~��7�
W��H��E��
z�J'��<�/���3:����0���B�z5�0j��^��W���Qs�LO�[Ci9�l�����������=�wC�@C�l��:�T��/��.�d3Fu�(�V�z౹��'�u#,]k������A _pV�~eﭐѮߏ��.V=>��10�"}N�x���m{�8DNY�O�D���ݺjce=��FJ�X�]j���J��\E�ɑ�Wr-�m���XV}�3�������9whWQǇ�VҤU\��T]س���u�|ynR )t.��b��z�6�7����1|���η3e���Ћ9fu�t��ᩆ��6��Ҕ���������0�g5��0[��h8y�]�'2��m���������%�=�ĳrى˳��w����j�~t��a��b8�CY���n�
���n�x�Z���e�=k �˧s�%�rma�y|^
�G�����;��ο{C���-�LG�H��O�ԫl�bW����h��fR��8�����˥�9�||ˑ2�a���g˩Dl�Ē�6�����+g�y���~��|D\N"��>�{��>�ו���"�vhk�Z���E�qq`�����v^v�/)�S�q���.��k�M�rŞ^��_�|U�\�pD+�ڸ���h��@mu2�3/)�-��j�.tp�#�Y���I�to��I����9�Q�<}������a�C��B�Y���溏�f��nnEx�~���C�e��}�X��g�y����衾Gˇs��%���$T��\�nT��k
���{�T�T��^]���xۋ�u�:Ll9Yp�?'��|%vm����Ѿ���u_�{v{�i��4� x����ˬ�̓������loL���	36���=��5�J�7���X�&9���Yו�t�R�+"��O{G���e箋N�w4U��t�`��xTH�yP0�9��=��;�pX�m7L�6��5��n�-C[�C�T*�Rr��,Ŷ8��r �f"��"�ݷ�]X�yS��
�H�	��\Q�ڿ}�Y�ϥj�C����]�pv�ь�f�$�q����[��(�����oxpS��4[�q�o|�U�������yT��c���	G^���!����+ޑ���c��6K%h�I]?�&:��^5MhBx/�&	�mK���G��������q&�����o^î��	�gO�v�L��)i��vQӟn�� ��S{N9�U���m��f�Rƫ���태��n[3)�ŧ�՞�o���j�q�k}n�n�[������ �ӂcҒ�}>K����K�WP��Qu2V)��|Kz���FL�z��·�UGX*�&��=),�'G����`^ 9��e�7#��\�����'p��h�ꫝ����ƹ�T0�l�xũ��������vg����ۛÜ����O��M�Lo�{H�Ӽ�xJ��+�g������6��0R�/��<Ƀ���S��=��9@4+�o��C���*~ۺy��X|�x�A��2��wh@�wd�j���C��m��u=��f�Zr���\�8�X�+R�f���-,|/�Ɖ^i�ַ�;W�n;�D��ڷ0`�$M�a�^�ޅ$B�0�tb�PI��1�V�T��f\M�A��R��gr��TZ�8�U,C����+����k���{~��]���]KC�/�C�;w5x6�נJ��I�3}=7������~�Y%l���M�(��s=H�_�v�	���]�z���ʼA��P�'���H>�e\k�ߣ���f>��플�I��#�x��}q~}e�Π�E��LT��>���sٽ�/ӹ�uZ1����ߦRJ�R/�*WV*���>�x�Z�5����V�uV�={��ּw�W�H�\G�˰�)$��S���\}�a��[j�򥄦��>Ngo��2ϋ�7��Z咵3&�pS$�å�yV=+�G�3fJ�K���ϙ�4w�KL�=�׈�U��c_o���˻|5�m��#P�MJ������ghvy.6��f&	̖�ii��&Mu�y�L�/��n�w��4���@�8����nҝ�\��e0rgM��!���9�l��|�>�_k�u�4�jx��.����zi�d��
Riw���9� �Ӧː3�e�A]+V�g,�~+)֕�����G<�$�ՆC6s��S��<EԶ�P��=�Y���h�z�)�LZƀ�Yg�K��I��Yӯ+��r����咢z&-:$�a�j��)���0�l�S.�[=���������٠D��ѻ�hh�1�wSS�I��$���ojm��t"	�W���)�pX��^��S��x-���8���v7e���8�j�z��R��L�*��^"8�����Qt�����X�χ��-9� j?W:
ְL�{e�@�A�:�r�������}�n����U��w�cQ,aC=�F\��0��ڹ���G��v��Y�0f��&^:��Ǟ�*��$Ȗ#�X�v;:�4�W�3|'b0��<s镽�p�y+�RX�O�קM;�}U9=n�/�K��V��O:����o�0��c��:�镾S�"��:�Q���b��ztw[��Mq�篰
�Q҉_�LƲ�dnq��:m?T�u�n]�M8�e9<�����#����XA��!g&Tœ����t�I5��߆���6Q�&zOq�6��s���&�/��ysX)����:a���\���.��^��4��^:��N5�C��8��w6J��5��>����tdVa|"�h�pS�qCؕDCa���m(��OMonɂ��W�OsJ�C�)w��|а�ݞ�[�#7��\<�EGVX6৩`�d���F�𠽥y���ܡ��Gk�*���H�������)�y�i_u�a�+ana�]Yn�|5A)�L�1�vS���/��N8��ZH��#S.����v��L7\�R�%3h���F�;��|@���g���A��Z����o���b���}˖oԅ�O~���Y`�g3%�Q��C7��K5�a_��
�U��k}O�{(������|��s=Y1� �<�A~�x^g�]�z��Q}+H������v3���7�d|�x�{�}�޲��j�ǂ��>+q��X����S
�1�t�aKg���{�{z{��r�f.��:���������74�|�%���@�W/E:��(ub��X�����MI�Vx�R$��2��;���g����'\=���������$mk׹�r��;�K[hE(5t8�̸}��Y��N�(|����Uŧe�g���jߺ_������5�`��S*E�b�X�f%cΌQ`���eΨqԾhz���h�l��w���>s���
�\mm(��WUW�TG_]�Pg"�\'R�d��]޽�w�=������{,Ƴ�a�K46ûZ�u"ŕ�āfn;���v9
Gv�Q/`�y$���8�7����uf����sJ�_>{'6�R�8��F�S/
fk�oA�\A��K�X�Nfe��$�E]��RI�0m@E�*v�����m�;�1lzZKßb:�k�wK!b4Χsod�"�u���ݰv���ځe����b���8��-����HX��PՌ:�\����ǆ���}O��s�g4��,G�Sv��)*���4�˽xw�ߏ5���OL�9��x����Aʉ0��5�Uo��{�va��zu�R��\gz�P�J\��,k�=�O���s������}�P�iZ����p W�-�r.�����7"��W�أ>r� ��0��Vm�ڰ���zEA2L�)^z�60L���
�e#�<Ԫx�?��Pv�>'o;�~�h����
M�M묛Ͱg����%�.��K�r&������?�]�K�F3�t���<�Ex@�F��rop����R����C���J�FϥV�/3ʥ��G�\9JwzW������Zf=����x��0�~w	"ÙoJ�J�Y��>�Z���W�n����=O�?V4��`rj5�3z���Xg|�Vt��q�&���a{��59n�
�yz����{D�����6k�]�2��V2�"��7l#b��[3;����~����
*����������+�i����D�Է �@v�:�Q`�C���2xp�y?o��͌�q��5�_uB��pY��Y���e�Zo�(3n�ګ�	�)�[�+�}#�T�]���Al�9��X�܁Ɵ	-ݥ����]y�{���H��Q}�ׇ}[o/30v%sp%o��Aε5�5.� �"�yk��ٜq� ���:���Ӵ�����i�~a��7jT��i�1%�������������Ŵ�]�uwŊ�{'�nS��A%?-��V��ʈN��(;�(ȗ�PF=�r�1�SU��|r���E�G�wz�Fs'�M�e���g=(sXgںa�֨�4\��ؠ��]zzoz��wͼ��^��r�Z�:��^Sn�l�h<��,>��<�ȃ�-#��@���i~�=����)������ʐ����{f�)���i$��a�*b��������5��s%�{�����8�� ���&�"� ���}��>k���Ǻ/�Uᕨ.^�b���h�[���q�Y�����Cs#C�&���GR������Yk0uz*nF��m7������=>j�x�n��P��xT72�G��=��:1�~VK�;<Yѭ�%&C����mtz�Zw�RS�"�����$xQ���<�ZI�৕����7*z'�����k�o��8��z���ix���tV�d��3&Â�&�Cu�B�YRP�����7��=��mL�8�dn��q��2��u��Tex�ԁ-�v_l.��I�S��ҕ�mC���W���A�D�/��k��y:���pa�[�m��!t1�蹓>������a:<�!e�.NF9k�i�ww|^lӯz�.�Y~vǟ���P�����y8�����8���OR��
��?nR۴d��s�Mi9]~jֻ��Lo�u�z|+i&Mu殴��nX�L�|q��J�]{���SFl|����8��Ξ7�K7�R��W�L�V2T/�w��� ϶�tWG��<2w�y���L�w��v���luG�c�ٞۜyH���ʊ&4)���v��D��aj�ރ�=�_���L�֘���rޯ���t<��_i	�K֦T�+�;�Sn"���y�y����aQ�sBm)��E��~=M�3�t�dP��Wk���A���F��|�9n;�v2������x�����T3|'b2z��{��o�y��ZG��]�������?���bL�a"9������x��^,���F��Y�����K_i�~~��Sݹ����?}�����,�8r�|�!�2����(ؽ9��yF�������x�>���Kz��_4�]c/`Z�h-<Q:;nLi�~�����o�c~�$ I?�BH@��H@�����$�$�	'��$ I?�	!I����$ I?�	!I��B���$�	'�@�$����$�	!I`IM$�	'��$ I?�	!I� IO�H@��B����$�@�$��1AY&SY���� j&_�rYc��=�ݐ?���a��>Gހ  U@Z��Z�@�h�B��` Thm�P4 �Cr �kJ�-�5�i�U�W�.�1l�5�i��X�[��*�FV�f�kUmJ�)j�e)j��%�ݕ�VՌͭkM���mLmM-��1��(���f�Y5j!e���ؖҪ��1�U���2�n����  3��s���n��C�������3c��ۺ�U]i��E֕���gml���uS�c�Fξ�T�K{���kk5l57� ����P�ΧP�Q�m����4��� kuU�v��v9me���S��l���^{:��nT�ލǹ9���y{�u�-Z�-]]��&��x  �{�5�E �=�}���P ��׶�  
���   (���E �(xlQ�٪��ushW�y���V8��:lϭ}�ە��+j������؊ַ� �㾚�=�{ޅʲ�-��٪U���V۵k9���蠵��7Yj�����ڥ\�c�.�w3��v�{��M�5���l�խ� >��:��٪[��w[l`Uw��=j�[���mGn4Б�i��V��nEms�מ�m]g����n;m���Ш-m�&�Ŵ׀ {��jwn[n�;�f�n]p��� 3�r�v��l���t�P��[(;���Q;��S&�4��f(� �(S��l`4�r��w7E]u�&�� ��pwu!j���]��,��fڭ��  �=hwg@�\ kd@wwS��Nwr���v8Gn���˃��w8 8붵[ldU�e3m3x  \�R�X�k����i�mNn�P�+��P��M��iӺ���u�C[Z��f�&�x  �
�ـSm��i@���7p���dn�45;� �m #f��=� � �%IB420@�  �4"��b�P 2h     ��d�UB�4�1� �&L&��~�R�        M hL�56�xDɵ4��i��I��`��h�jf�F�'�m��}}�çmk�o5���Y�f�Z
w��!^�s�·I��GAI�H��?HT	$�4H�B��@�4����;����C���:I$�BA*�$�!�K4!%	!h�����j�Ϸ�>n7H@��&�է�����8�A�sP�A�A���c�����u-mRלZ�z����[�� ˙���%0w7"W��;��4���-�CS)�ܸ�xo���,���[oC� F�@Ghd�	V(j�ް*A�������� H&b+e�h�ղ9!�bq�2�i�D�[Q��K�N��x��
��n1������n��]��k2��V �ʶ͒��,���&J=K��H�
S+.�+�*L+�B;H@���KB6 ��+���1Q��E;�d��]�cͭ't��۽/mcZ0\��v�r���bZ�7tP�4pL�4�T�h��Up��6�>+Y�q��EWX/U�f���A��ѯcF'���#JZe�ݗND�E�۱D�;ս��$8-�(TV��'�#�4��]��E��`XV��)�Xpڷ�g�һ��i"���#�`:5=W#7Yx6�9,�2����7r�o2�%GMM��tD�t68�ɘs���U�5�k!h֚��rd$���n:@�46հ�x�
�l��N:�ٵ,S�A��oVn��L���Q�Ӓ�q�)�m�B�질䔶�XyYPg�m��p��\U�!�-�'^�Y�xT�h1;a'EJ���{�R9�n�j����h`�6=ĭ�"t�pܼv�[�Fl�Ȩ4����u�V�yMyi�㙧�N �d��٣xV���m�;�⧶��e!�������H^*Ź�z�m�[�I;�Ox� �Ѻ�wn�\-M�Q73�$�Mb��+���5k77�1z���T�]�k����<��Y�f��{J��ժ��a]�KJ�GZpae��M�� X��\�U��) �S�f��o(�-UK�Q�S��;��%w�AYw`]fӗK������^1ugpb�����b�h�d�!z�hw4X����JJ�9�h���5�M�n��]3�;�e匑N�H�f@�.Q!-��w�]��׭mro�j꜖��֫Y���M<�@�X>9Y�c�7M��˔�6�mX̀��Y��TcDx�kB�g�V�A0����+��i������F���'M�V���XB�*3-g
Җ#7B�E���e�c+P����c��	� �t��ŷ���ʧ�1�*{:�c���JW���W�m�b���q\p"6���v+�ۨ��	��tYG���=�y�� ؼ4�L�[`+�ł�:W�e��*eu�V���7ʭ�df�,:�>�>�~ț(1ZĎ���jD��-��Q]�k��h�e:�Tp�*�d7���sh���tA�D�O��A5"���{�K,���:��k��+�*�Xӵ���k�!mh]�� 7��$�QЊ{8��XE!�ɀ .�R\Q�;�cQOi�܊
ؘ�#��c��4�l��U�V �T1����
6�4����u�zŋ�)n�����V���IX2<"� FK���"�b˹�� ���%��+�Mb�׋Z��*�U�B�����+4$6����TOr�~�f, �K��(ڽڛ�,3�C6�:i�˿�i��R4��k����Wzq<�Ql;W2�X
2QkEM�YN�H����M�T���F�*�^�~_nб��Ug���k���c.�>��qֵ:9b�̧���$a��,�B�ua9W7~ä��P��Km�U�7�g6P�bS[Jf0�cǮ�KS4��[�l�����2��'�볲��z��qH2�J�]�,��ES4 �K9V]JU�,U#utci� j����lL�Ba��ś�$	��8A7d��v2໰m�o� ��k�6�)������6DB.������(��T;wY�ѫ)�BT{���}��&��;�9�!k mZD��J��J9
��n=�f�e ;$�)}�S�u�]�-j��tF[�1�u6":)�`��d�[�`8�Ж�]lK,lƬ�T��"�+��K>�kq�I2��J��q͡��ܙ������L��n�1�SrF�]�ۭz�_ F^1vjۥPC'�YL���Ԣ�|�Eҏ~u�B�ۙs� ����E�{�as o/l����HM��LE�ے�Fm�d�(��\z�j[��N"e��\Y�c;H̦��p�Kx���
��<�w�]�^dxm��}4�QL ��-�.]��ܚ4ILwY Sa;�Z[�YW�H�-��
�sw�9
zx�X��Ou�j�g�l�4kWo���8-o{u[	���(v$��vM��8���+Y��B%��Y��Я,�"�[$Q�}ُ���,�-m�X��+��/j�Mm�P��k3��L0l���,�6�M��|
��'�`pn�J�t�r�8ì��c~��\dYyF�+�w��kIf�8^Q�ǹQ�pl��L�R��i�
jZ-��HΡ�.�[��%Zt�$��.|�#C,͖��0�\ �c�N���˫pϠoE]�f�(�ҹA �yok��Ј\J��+IYB�+p9�)���:���8�,��:+i�)�3l�p
��1�&qV�"��ufH'L����h�&j(�S�or�,ky,�Ot+*�Z��y��1�;N�j����������Vj�-74h+$E,���S)63��*��v�p�ǤYZ��u�lsk�]=UI�V�\�f��-�E!BKn����#B��P5���������"�fM���Z]-D�op�4�oI�����v�)��	u�o.Rv��t�}y�b�Ӛ2��ڟP�ӻ֣�&�;��i�8���ic2F%3�[Imwr-3h%�Y*�)ƥ�'q	���[�.˹X	� Lk.��Ի��km��>sv���%4U�(<1�;N�N=D�]�O,]�&���#�f�\�K��ݨ���l�wlD�p��|+^�;F��A�H��撢�r�[�Nd4Ju�)�}h���V����Yaڗ�[��V�x�kI\E|��'n�@n}�$$��UjM���vM\2+�Ed�$�b��n=�l--��fӑZ%�V٭�[�ɘ��̓h5�u;����t�0�j�؀\�ٽ'^Y+�z��#��]���\�>a������x㼥IV�
YүlR���9��<����Stʵ��� �@�pl��1aб�q5�c&��c�̈́(����9Y��^��������r��[n�a/�4�+ͱT�ıe�m1�L�xVc�N��H�2�ۼװJ `�;ڱ�e�b�f���8��r�H�+���i:9sv�w�E6f�͇eYUdm"��mXE@<��	��+unR��b7r(��˥��pؘ�j�#t�D�U�G���.�k`��&��-���JN��v]i�N��u`e<�u���v.a�5 �@�HV����YA�m;�pj��׉P��e�f���2`+$�if(�BлG>�1�լX�s4��[Krd���y�0;ɷZ�{��M� n�\�j���Ķ�*�u�f�5�����]�A��c�)=�+�
o��/XE'��#e�� �Q.ռP�!��lӣ��0%y�k�h�Ņ�]�n����Ŧ��pY� ]�4c�@��.���7-��Ԋ�m[��n�!������6����.R�lb����R�)TZ�I��ʰ����ڐK����=�@�5*�:&A�� �JR�*�4�tf��Y�ABa��l�'u
ĩC#ۢ7噍6�8X�r�p�R����̽x2��	�W/)�x���[�K��R�\si;okvt��WV���m*wa�)_W+%u�<:آ����ߍ ���􆴭T�l^ąIiV��6vm��V�hu��k�N��gh�gY�Q)��[��@�в�i��P���a�s.�A�3T��M&K�*96�f�Ӛ,��^޼*�dT�J�#�֛{��k��KB���Su�7E���A���{�.ȥz��;,ӻI�d��D�n�vLZ�IBKs(Z��W{���܆��0��4Jx3�jYF^�#�N��e�n��n�h�Y�,��Xn�:k)�N]�C��:n�d���f���Cou�&�'���A�%֋�=�3)-{Z���o-�q_ϟu_aK\0Ѹ����Ra�{��3/v�:0e굘�V��˽
l�9Q]b�E�G7.{R�/c�Jԗ�ض�6Ad+Z��Hn�n*ɕ���Q��6XUxТ�'3��SM/�x&ʩ�>[�����4�IRJW�����bk(*&ķ����5�ugWX�������r9�N�Ӻ�KX�����&�2���f�5�Eʵ��X-i���(�U�U�C��Z���+& La��&�!]?�fM�
��t�fnTӁ�����Xtad�%���+^Y�!iܭĭ��=�~��M ]��0�3H���/.��[�0�]���p�n�+^-W����;���x�+`��Hy�)�`����w�����Aݍ��b�+5�i"^� ��y�ypg�=���n�Dm��b�Y��~��B�b�I�T���ǹ[�"z��i��$��T�f��5f��6�픞�r[�)��.ի��� P��J�1$�&]�	����(w=v��λc�H��̥������V*�ޛ̩�]\hby�Ԥj����e���e���t8�
Z���-J@���tԤ�Գ#�OM���1���w$�n�zΠ�#g�1��uV��;�R(����;����t���*ĺ�V���2��ЉĦx��0���l�WB�����o��.�fR�͍����/p��/Z���J��{DI.`Gm*�� +;��J��u��ý�K����=�6��8,@��7ŲQ�n�c���\ڗ����n/L�p�8yѝ�㒧�AQ���f��)�Y{@�sDȻ���p�����P��aGy�ɋ2v�Z[X���×Ԕ�ʙ2�p �e't���H����EW�pß�.�G20]�U�G �P�:�S�n��*)w��Ʈ9Q�2#���Rx���\1E۷�3V��w�*�����P�
K�ψ��h&�ƒj�f����9p�f�2e�U�t��ǐ�+��4���*�-�	��»���\��jkB�i��jH��W׆g\Uwݻ����\�	�%��wz0!���݆��u�m�B7A鬚��Q�I�ϟL�`��%v���eL�@�9$��o�#v�������d�p���}�@�IU����i�9�ۭ�"���)�a�U/e���dg7xk
Q�p�Nq*���WgIk��r��ŦPB��vy�M;�=�eܭ��:ݾVã����"s ��mu�t���=�e>zx�P-G%���3\#sV�X���{ԗo���Q�UV�
��*s���/�Yh�F�˳�m��+�A��(�s>�Z9݅�E֋O�Z��Jj�э���P!��ɛ5�c�C���u�4���E8[6J�9.�� �׎���F��A�p�NY��	�B��6�c�q^�iz���l�+\SJ�l�,sD,��}t���!��BTOzR�}[�q���l"������6�Q�/�-����{j�>ν�[�d��Wt�̗�:����P����!��$��;)rUf�;��k9ʎv>��*���{l�w`읷��i!�hrC�]nY�X��A��|��z��w��[�1mӐ��|�m���f�=��K���:SW���A|jwI��d�����E���Uk6��t� ��(��,��1)���%�:��J� �t�\�ֶtS�N=Mot��i�m5cIB�.9�t�1�%B�g[Ҷ�O����y]�_ʺ[�]fd>�^�0�\�$���[oxh3�5&oWfǨ ^�3�}׽��QVl,����)��:ӬT������N
M3�u�(���m�y�Wv��͊<��np�7�&�(v�����K7�w��Փv��=0l�(CӶ>T���a����87qf����0�I^�V�F>�O�X�SUh��V��j�#]�����.�"_`ܩ�J4�i9f� �Be�{*���j[����nq�aC���$�/*�,<}��7����vK6yTY�o�2�E!��Y|��D
g5��^�7Z�PL��Wz�>CV��yDA⫞��fڱ�h*]
�X�ud�ع^����7�:�1Q�Ǌۺ"�U�n*���u��VB�� �:�NpL�5ݻ�_%6."��Z�5B�NV���z���_3��8��iT�3Փn��bwJ;,���.f�|VLC;���=Zu�o���5��(���մ-��XXz��%^Q�_u-S��`���F���d��kR최���'8���2�0�3���P�.�u"�;\�7�8�`��E�a^H�
=�7]F�Zi�X�[f6�=�F��\F�f7Hw����ٝ.o���Z�@�/�]��GN`�����Y�GQ°��Y���@�����=���`�AL��}d�	�g���S�bDi�ɽ�B2j��fԲ	+�s��5P~6]����+�9o3/��h+'J��U>ePw��'qs�W�3+m����p}��qo	{O�.�]m�jW	xa�Zr��+�[��� ��%5�k�b��d*Aފ�� �P��[�y]�"�V{�
�����[���K7]d���Kj���
+�Q�nsx��m�܅���U\������/�;�\�V��Y�� ۺ�x��v��M�i�v����O��4&���U������ۥ%�`��D�=�e�e�������X[9��Ҳ���15e��]h�5_h�1��wo,me7e�q[h�*T�{�ܔ��mI�^��[2Ʈ������]�*�덹��Z��\FkR��U����MNyQ4�l��U����]�5���`���x�N4a�{�b��0�j���oe�\����C�4lt����"�Dn�������K&���J̈p�/8��2����_K�H�ʈP��Yt�ؚ��\�BP��w��k�VP�<�0]qoc#��#k�]�6X�x޴n}ej=ze�;�-�N�v��4ʦ�ԫ�w���J�fJ� ��n�%Vw+�nЁM]�0B���`b�u:s�.���6\ۤ3q��V��v�����[�+���%�d�b!��K��B̡Q3�@�f��I�Ջa�*a���w޾���Bx*\=��{ݭ������t�Ok1F������idX��b�)0V��|s
Y,9���0q\��F��0S����K;F��v�0)g��-JfK6T�2��un=�V�5�2�;��/�o)l�6�򣖔�st,�1�p֍Ef>�6���cu�Yh��=C8R[[C��gv��c�9Q����b�|sv�q ���e�3Ԍ���Ҹf��%l�M����viR��Ȋ��e�0�d��u�ڒ���Z j��0*��Ă����ؓ�wtQ�ŅKpK�΀y�ManL��vΥWE�s�K6�P8�X�l�i����ɺ��1�,��wE�}��sD�@:�ǚ�k��\�(�o�Kox%�F�ČM�R�������M]]�T��=�է%B]��WUڀ�7G� �mP�m�(L�y���{0)@�,oh����^��-�-
sӊ��\Z�S����r�[�s��L�P5+-���� �]](]��8�=�;E�x�J����W97yv�,!����u��,�} +)��Rcb���'��3��Ⱦ�ea�v�H��P�s���=kR�M�rc�d�8o�ot�2[�IM�b �t.��-mЩܝv `�N�nɾǨ���t���A�i"�nglj������;�0ZYdo��k�MQwo���/GmJ3�Qo9�`�.�	�8>Z��ND��a�iW��k_��:q����3l���ɽs\�WL��)Z��iU��=��Qb��䖰�Lkr��O늭�"lZ���зwM`��$�F��M&��o7.pW ��w���Ǒ�xZ�f�"ɣ��Mt{+Q�i��D29��ՔU�dׁ���D&n⾿�.+�I�G�Թto���{.����39� ��34Y�������!���	����mR
�;Vm]Y�kb�$�-b<d��f7C�е���ݱ�Utm����;,o�֝��$)l���<�Pw���͠/K�����eN��9���E+V�М�p7g�c�6�3~��yi񿲹ܫ#�t�F�J�������e>ǛG���Rs�K%ZӍ��?+9.��z��<jCz���>B�hTb����{�x�Qlnj�tJ�ZO��RpxN�#$��p󥜳��۔�lkٲ�y|h�n����&a$;���ɭf>a9gI&�\�:f�r�i�=����ž˭� �_K��fT�����n�r�Y���4���\��%�ә�Ȧw7�ۚ1�[	�x_Z�)Vd���e�Y�r�y��ؘ,پjV�2�%w8���F��M��Z��S!cP���	E�����b���w-C�����/�>ڍ��׋��sW]�D�ET�ۚ�ܫ}S�-�#�c�G2�V��]Ca]�d΅�vrr�E�Y�����ɲV��ݠ�C�n�*��/�Wn�4A@kw�T���j�.Q�M�M���qCSo_n��cz����oD����ԓv4�<��w�Y�Gn�a\).iv���XĞ�J�'z��[��r`��˙<��j���Ln����:��C*TWYp��twWl�0[�KW��]0�5y)�E|Ijq�ʵ!�ƒ*�W,�#H�(E��hǪ��H�ҡ�n��e��|m��)��7E�Oc���t�iٽ���WԷ�;�����d���G����P��
3 \�bB{�il�*ov�^+�zm
���t�YV^����l�R����HX���%QZ!��޻�"������WT0K��!z譙f1��U�:j��y�\�I-{���#aV�:4m�ڙ.�^�Дx�
j%��{@��%�N����mb�+:k���N�������s	�s-�9q��ʜ�U�:��r�G��*���J�mZ���Z3�9��P�\�e���B:D�ƫ�Q�F�S�vvі�d�1�$���w!�1<��k�G���1K��@���Ѻ7��c9�C�ѧ�\���b�_vw#��\9�p�6ͳ�ni ���_cWK2ӗr�����إ��� 1p�j'�su��4�R� �@<�FS���RѴ���%��[�եh޶�r���E��G���9������Ʀ]���u��0��������Tu��V�(	&ޅ�팗�Fdr���38�Ľ�JƼ��j��eI�7P�;*ā�r�:�*�TP��	��I$�I$�I$�I$�I6q��*�������Αu�o��V9�oTى�[�
9��p4���4D.�7i^hJKi��Y�s\i<��<��iv�+�5�X���:K�L��;�C��R�Ye+T�����Β�B���� ��ڇjn�Zz�wHx�eW�f�6]'A�^�2+6��Ք�\�
p�]CM��'7������i��N���+����;>
Y�y9�y�cC�G��0wj�oDؐѭӼ��	��u�L=Go\�T�F��
ON=�MF^��w�ox�B"2�3I�P��![	ZX:I@��K��o��'T��])J=�����K�8̕n�Jh�X�-���9��a-�����^�s��H���)��|���둝N0s0�	8�-��k���hu;�����e�=��nl�w�Pݗw��}7��;� ���J��7��z���~0d!O��f�Qw�@�n��L����f��;���[���7a٧F���*���Z�m:�mWl0����oa-�b��Td=�`ƖՋ��A�[�n����	է��X��R���4��Vp
���M܈����px���q�mX�g���n�t�ՁZ �C厔�&����t���[tB�ل�o!�W-��\j�5�V1�Z��ſ"80�nڨ;z���(�5kT�Euu>]m�G��=��N��y�� ���5��7sl�L�հҳv䥑Z����(꥚W�uI�y��-j��yt륽�[𾩶����V�_5�7#�T�ml_��nVE��" �5�]ܑe����;}�V$�	"�z��3N��@euv��F�k�I\f8��/:�#��ܱ(����	�8f�Y�1�����~�Hu7I�R�f�.��J�X����-���U��i��s����!,gU��Z{���ʵB�\��95����-�I��#1�κ�L�[;�=X��*fG	3T�(F�l:}�M�Ȓ�qv
��,ҙ��؉v*��>�M[yIѷ��O������E��E
G��=�����>I������@LC�'���Uk��{m�Oj�[j���;�ׄ��m]) �J��X�g-r���*-��������ɵx�����M�1�o{��]�H�3���:�h�֋QxaU�N��3���v���=F��4��P����I�0��-:�Ma���ʎM�U�-��}E�<��s!v�b�}��nGq�sV��30�6 B<����aU��X����w�)�9�(bK�4mq��;6)��%ܤ�5�/��'bgD�����1�F	�E�R��n 1Z]w�+~��B�v�Ֆ�A��Kdws�]
Jޓ�w�'���θAJ�>�P��e<�V�9!�3Q�k;������v{�'F�QRܖ�w�I�2��桶6X��<$}��iѦ����H�i��|�̦��XhG}L&U���Ջ7AV������l���߃��Aw�N{XX��Z*��3�'f�ԍaY�ҧ���r�)�ie���JI��K]_(I�5!Ы):���nؙ�s�7Gb|��L���X�#w�!/:��U�լX�3�j�Y"�CHef�١�%�k)��h���b-6�l�rPO��%Jܠ�s;i[�%��X���]�	a�C�db��;EϧWCwT�r�}Z��ݎ S��Gg-�Ѭ]�k��$SmK��
k�kQ�ku��Of�:�P�k�_X��ذ����@Y@v1�*���mړ���XV�w1HgZ/��V��y�ݴ��A,�g�^ιwv�t�KlN������o@*YtV�ɖ���ς�Z�3L�:&�S
����fnΊnK�M�!��;�l���EI����	xEf�-S.W+4�{2�J@������!�W��ji�ㆤ��9SrVS#t�s6���k�t��wK��{:����e֭2��D��Uz鎈��I\����8|ٔ�v�ל�Y-��z�KI��A�8#�+MȨ�H�kv�u��eov�v+��)��UmZӟp\�����b�Բ)�՜,mKRF�Ý5�2:r|�yp��B��lՐ�h�4���V�v���@[�V��+Uv������ɶko0m�0�� m�sZx:�u�w��nU�4�L�*n�<���.cuf���O5AQ��#��#Z.G���T��M]Mw�B��d��f�f�δ�q���Zz:� �yb+ ��}�1Pg'��]"hg�Hg!`�ws�*5�n\Y���C���#�z��L�����pjB8�̠-w��/a%�y�Ӿ�2V����r�AbDG-�VYa�܎rZ�u�ߥԱp�$t�Z�^���fރ˖;�wp�n�yp�D#ӷ�o,����A���>N�� �:��n���oS����|ilX�\��0ލ,o�6G�]DfTF����_:{8�.�nȭ�o7�'���ѳv^���k,[;0X���5�����8}�|S�S3��5���ᷲ:�-4S������Nj�ʸr#�E��������:�ˡ�VQ�y2�mv��d%hWcE����+�) �{�(�1GZ7��-ǹ��m(�B�
�V��&e.�OֳK��3+n٧0]*�xs�W`׵h�ܤ&����S��N�%�ૌ�,R�QRb�ڮ1HE.�<̡����ܓ�h�-B)����/��0����v����G[�n�=Z��Z��/7�n^�<��y�t6�z�i�(hT�u���m(�G����`N���m͸nj�=�m�[y��=�����5��£a����'��(�F7n-(on�-�y�^A�*�8\�4�%���lv�jQ:����J���]5��˭Qq�t,$5�5>|�t�P���L2�ښ��w	LEwX�Y>���RP��rCx���A�}(�Inv�-,(yZ7�<(�u�))�e1.�/I�]B���r�u��֪̹��B�ͼ����K��ggda����A�ctK�UD@�8\	}�x�n���'��[�c�#6�iv:$*µ�(\a���V;SM� >��*��ۨT�k�L��K�{��WW1��i�e�g��SlE��胬�0�֬����O��c��C1�mp��jnᤈ4��S�\]g�=�!��+VS�T�4n�6��K"�9������q�T�n+�\�Q
�,]9+�Nf�@R��D�ǖ�E]\�_%��'��\&���Yg�od\�û�)��u=�H�강ٴjx�	Pvy)^} V�)���v�H���x[�k찷�f&h�9Ƚ�c/r6ά:��0oo�P�UK�Y��t�v��o&�֬�����:��jg#�t�L�F��̛|�b�6��f�oT�m՟���-P�Y5�ct�j�j�c�gX���$CR�R�@�Jr���q'�oH;6�l�+��+�2���xVa�"{A6k�������:��\}v��)����kzg1H=���=����#r�tXW2�Vy��G���jqm5/FQh�0����ƻ*��)�8
}�5p����
�
�܋�|�f�!��@��H0�f��΂��h��k���bI桪�m�+��Y��	;
iK��85�]4�6T�z�60�)Wo�A�敩�6fj��F�I5�|k.���Y��� \^�ޢ�֝N��`/�o����g5PF�J��K��X�p
Gu��V������x�B[ٍS�o6�h�����+�ກ�ME����w�.�oP��,�5:�&$vU��R����c6^��e���h��H�HEzf��(P��q���d���b�!�5|n���A֧�c�1����R�1:��Yr�jλ�g%�O/�l���-nӊ-��p��/�HEB�]��:&��E��Υyk)�5g�i!*F�q�3fǥ�Wʰ�I��B^���nu�1�n��+I�B��?�u\�]�W#��(����ӱ]��RĔG`��:������]��Q���A�v�;m ��ɫ�J�_-�T��Up@5��v@��ǝm�y���g�C��Oy={[p%K����{E,PJv�Sl�S)�tVE�te��%���<	t�7�v
�m
�nE�,Fv%�*��j*I��c	����\i-yV��x'fJV�2h��AԨ��T:��h�����v��DP��y�l��\�V�˟=(7L�Yb4ep��-����A|Z*����p���^�xY��-e�ƨ��F��D#ͫ	λ$�#
�����f�:����u����?d��Ë�� n��f�]eO@������r�	���;���f	��������̲v������[�IwP���\9�(,�$�Z���!x��"��Im��˽y�x�|2A����a�hA�$�K�r�ol��y�q=���-��q�b�c�,���n���?��.��t���ݘ�9q[r��H�m	Em��Fe^�K�����]^��
P��^�cn�Ȝ�ΐ�Y�BT�˛���̸�pY�TIf|���+�neD���z�
�֔j�1w�{��\텘�oK�l=�ʄ�9C:���#�AE�cV�z��B���k��R�.j�/R��Y�w��lT��2m�nTQ]����@f�V�ŕ�T�R�[B,�5�`v���騰ޚ��C�T�$ѧ5�j[LR�����:���d��YΣ�*��\2���DÜ�)b�E�[JpC���
C�D[��r��m��nӢC���x��y+��D�t*e�FN!�Dee��i��X��:�7v*K*�|S�5p�m+�$�0!�J
�y�b�.m�u�q"J�\�b�b�V��ucT�(?���ʰ����Z�9�'����"���SDPD�vm�W*�(�Bf�;n6��	�-.$��ŕ3�r���9��\�gs�Wť���c���"���5j]�:�y�A����m�q8�<�MҝJ�+�Ô��=����9�B�B۳-�g�����)����;���i���T�����^7�r���eg1�,�5|㣰Ww,�V�Q���-��N����!""�� ����{��z?c�ϲ�,Ή�V?T�(܎KG�s6m#7�l�<�am�7�e;���T�Ydc%���ȕ� �GC�-`�~�:6�[��,&�"����M!t��S��s�x��
� ��.�NJʒZ�Y�ء���'F�0A�r��%h�F2���\#�2�5��C��uC�tN-���nS�X;�+;�+N�xܠ����9�oU����p�M��r��A��֎��V����/,;K�f���{}p��lZ;V�����R"觜F�]��L딃�����Tw��:
E�0�A݂�W��WX4�/������jG�\�q@7�Ⳛ��m�о|N�;��EX�J5o'S7��/k]`����4����I18��f%�e����X,*����ɸ��Y!�/qt��֮�@R]:��5��㶍f�BΤ���q���ˣ��vdy�\p)��ei���tI:�0��]�)���ɖ��]�d/SZ�׊x;����>,:���Y�sR���H�i���c&���-�QV�Q����	����2Glau�R��h1EE��Xд��,m*[(ȕm��+KDf�/,��V�UA�aX����ڢ�]��b�,.�:�QL�u
%Kl�ԭ������X�չmlm��ҵ�ڢ��(]M-(���A�Z5�U-�� �L�TA^mXqj1���0����4(�4��,˧�j��fլ��%�
k(�0Ԣ�����R*�%�Q̪����Ԫ���"��5�kXX%Km$bu����ڧ	TQAAEc���j*p�E5����݌�F�KV�j��[�Q5e.r抦�a��6f��N���u����_z�wҭ*���ө�zu��t�uٛ[KqIf�lȴf��M.R���ṩ4���d7��4����RL����op����ݙ=͗umA��$�g�Ƽ=��V8�#�0D97|������ߠ=�!�NK5P�<m1�9��;ɭ��b�����I���#d@R˚v�M5��j�[C�������{LH�o9��r6�ӭ�֞��lH�=c]+�-�<��j��9ҫ݌f�cM�pt;��Y[����bn�! ���I�p�N1x������t�#�k4�vza�X�ub訾=E�Q��}��c]���Y�
wj���q�K�9m��|S[|����Q���>�J�eP��q��?�U�yMx0 =�PSgul���Z�1���ǐK�BZP�кn%��b��c��[&�Ҟq����Ul0�E�L�&3��mQ4�(�١K�D��%U����l�U`���ex���ط�u�<,�ײ�!6����g.�Aek�F�G��b�o��m	����m�O{�f�.��m��X]�0�}ܧ���<�<��פ�E�N8�:�����\_m�pL���pF�|i�k)l��%���M�%�׭bW+���k�������¦+n5��)��:o��9ۅ���JGԃ5'c��h;����R4e0KV5u��m��Ӏ�p[k�^�<�l��E{���Jƺg�D�I0Ts���Z�ե�����r	غį�P�۳�e�MMi���y�q��ڰ0�1�bpޠh� ҥ�Y9G.�A����as���ix�胜H��&���u����:!ڷY�6և�p���ݨq,��*�o�l��Eu��W^ ��Hjt)`��nj�汵��tY8�Z秛��k�y��wSwW�3n�N�>���%�	�J��L1{���zAȖ׈���^�fN�����,-W+�')�܁�M3��#7J�"/��m�meė(в����#7�S5��j�0T]�*�g{��Ճo�*D4����#,�z���Su^��������-���Pf���,��孚�w�p[��"��Inbm�����h����^��;����s�G��QI*�ӽ�K��\���:D!�E�eD�[o�sU��͡�����l奒�F�k�3rsePgh�V�:���r�e����4��krq&�B$]�:��n�[ݚ���y��Q�F�`�����2�� �2��7���+o4����	�����ަ�g=�>#�(�Oy'�g�n�a�˦�4�o�(߻A.fcz���R֩�֕��.�va��q��W��#H/��Sp��Ưu�땞���;���ɞ!�n�[�!KR+�6�ƚ�,Z�8�[b�kG+��mD�D������L��z�f�K70��F����CM�t�����M�ܘt��XKҪ���<��]/WI�X�L���[�n疵���\7ە����m;�2P��*I2{k�T���Oh��@�]�N*����t�E/X�Ʋ	�)飼���+jk�Pq�Vi�3i�����?y;75���l$ˡI<� ��튻�N򍉉�d�4��>W|��� <G�C9����U����\��
�I`WEY�TY4w�u`ȸ����ʛM��]�mN(�B�%P����5�@o`�yn=��E�?uS`��!��x
Ĭ�\i����U�|t�
Ggyb�'Q���9��B���MX��u� �V:ξ�m3|���E��9b�@nA���٧9W(�H7c�TI5���Moc��{�& !�P.T{�����V������*��G~%{r�a�W�/��~><5�S̨)S5"���n�r�ȉCs$J��[Y��o�ný�ԅ`2b��$�9&FE3B'SR�47f-�i}q�XRn�`����w?
c«�YJ��a�L)�'T��V�-'�;�\���!E{W�+�P�Ȩ�5��)�)A�JY��k~��V�������_��pي���b=PaET2��J���xײ��`��}e��׭���7�Tt��Sn�rt�ǝ97-�:}ts&�+��I��ncq��=�fgwZ/L���&��u�傓|{�S���;�Z�^1¥�E�w��E���܎��B�k�WR�v�kk0���7F���!���EfVE�N�_K��M�_p��Jx�{�Yv��ϸ�Ni������导|�v}�><"x�Fѳ���"HOβm8iަJ�h��
�xW���_B�Q�[ۇYvnC�� (��p��>��j��g�_V�� ��,��K�Vm�j?`�x���`�U�Zc`� ���ཊ.�� �t/x�/9}'���WR��N2
�4$�tg�E.�0j�M\��׋Sמ�i}���tU��8e�[J��I�A�\2���h\D'%%�5�n���n<a@BL��2D
!C�F;1c'ę���ι7�$W\z�z:a�^�{8�R,G���N���5<Z?k7.'um��~��Z�/]���n�@Vi�e��&�d
b匭�d߸� i:��q� #��鸺��co[빺.��^= s)@�>���|�u&)Ky�ׂwe����S����/L�	�/�0h��%�xB�r+�jY1��,�S0%�GW���s��p-e�tk�)q�'BE*Quy���&����K U����r�W�6��p��;Mذ�1]�ZE�b��ڿCʸD�gO�H
Nؘ��j3���وnlϫo���Xx�r���}|(mY�R'�C�&�z��~O
ϼf��W:��Ҏ˹~�.�T)��:�Z;�4�җ�8{��K�tNB�\�Ɠ����r�cjGQ:TMo�h$��^ f
��V����^w��e���v��%�����	���+W�}�������vj���͊���t�qwɞ�V�J}���z�p����8u�OW��|>�b�B�<*�_*�֚����pt5O�a�~�+<n��}�>4��"���f7xg�^�.�)���V2in�4Oܯ���R��-w9i��e�/������+�cR�;MmL�ْb�.sw�hܫW�\FLJ95'�A�����uXc�}㇮�"v5ʃckǳ��ս����P��X3�Pp�!�,T��V
��{Ċ�.��R��]U��a���#��ƀ�U�}��\�dH�u*:$��BL����n��ƛ����raE��Sa~�JE��vn@pJ�}W\�� 4���KQzy,�p�
��~οP�7�P�a��R4_y�7�Of�續^y�=�dzȡ��	�}��H�Zs��C��Jf���R~W,�#��O$�����=�t<j���^S
M��K� =��N9X:�H��/$�Ѿ����R�������~U^92!N5B�[�O�����<O�TS�7k�mx�"�W�k��X��4 0�
�d(Փ��E�{�U��T�ppP��� `���Ⱦ*�R�5�	���B�'WO���Q�\3�k%"4��ҼzKϝf��8oi-�5��1��u�tV���=�Thۧ��r?%���Յ�=R]A|����iZY�n�>�!eQ�Ʊ�x^���&�%��<^}jB�WTܞ��H
&;e)
<�9�q��2f�	�'�]z��4�#m��������BU�˔�S��ڊ���N��l��}B懨l	�%MԌ���[��t`�C��	 ���'�M�w�2��:t,-4��@mx���B�����u���3�尟
G�&�ظlכ���:�ⅎ&P���h��٨�z�/{3x�����62�sa��=��=��3�Q��D<~�GR�f�*_�����:��/�ʥZg��΋�Jj��B���VY���~�<�y[����U\*�H�V�����5�����dɞ���/�<��iW�x}8�~QԺi���*�0�{W��_�-Ƿ����<����T��H�O�O��*�v$������pq~�`����:��vEva�֫ �=��L�b[��>����W��k��;XlT��QZy�!�}�_x1�ʣ�-��.׭�л:�o����B�Ho���6��֛��t��F��oh'!@�d���\�Ȧh^��ɷv�����&s�#��H�R��jV�� ��F��l���(b�vwx����Q�Ң K��ߍ��C�&���B`ι׵���(��Ӱ�a�2$���zƺ
,l�Kx�=,@_u*0�Z�5�|>��Q�4WY!wς���O�i鮨h7������M�|$nJ�n}i��%G����̬�N�^˄r�$�;����R$c6)�JT	�C��!���g�*�z��t�j�Ԝ(�)���<Gl�LK*y���h֪���@p��Un�n�sg��>&e
�P_ي�����E@!�P��"�^4לZ�xvy�4�j��X�ԡF���~?n��+�}X�:L�t"֮7_.*Zf�jA��:�s��Ӏ����\�`}�ht��'BjәPX`��73� M�w9[��(!
���Z����>3Z��yrV^�u�,!Jm����W	3�Ɖ����T���J��!��.�Q˸�F��vu�b�ZkGQ�F���χA0%����;X�%�M=��=+�m�0��B�y���,+6�-�����N{0��ï�2ue�����兆��j���Aq�5b�֎]����%*2^�㝫�m`ػ`�����TȫQ��� x�3����VL�:{o��0��aS���w��[��]=ڗ�K,�٤�ٱ�(5	~��Э��9=v��d�y5�oW^�K�v-�*@v,��7rqcv�9Z�]Z�k{�a�G�)��qިo���Y%�
Q���-�m�ٶ��`��������ډ�{}�CA۫��7K�]XV�(V�P��dX�XȜ�ձ%�opr����U����+Ws�X9;��N��i��ɗZ u$wZl�c�a��n~~���;���=��-��n,\�k2C��ŝ�*PN*��l'�W�-�g��w�	��N��e5zf@��l�n�]����H\ٛ��{�u�'9E����e|}t�-�az�VS�l�r��Ҍ�\��P��#Q]��mA�v��\pC�-�c�bx�;>����+R�kg	���ȁ(��3A������|��3�Q���r��c�r����1��IO��F�qXd=�u�p�2��8��8�{D2�3h�j�k �t �6�8��:�x�����������љ<A{�ԕ�J��lR�B��q����MY0`�Y�{ٔ]�o�%'��f���2j�Ah�QU��`�p����q��"ܾ�ttv2�8BQ!W�<���C��.:̔z���ݩ�0��kvn5\T�GN�0ێ��Hr�'utbO.�S7P��Sf�8��P���@�{���F�C�%\������J����3,������u�����q%�������B	���*�9�WS.eb��(��������̢�.��U��TUGZ2�;U�0b��*TU�*��-<�Ԕ�6�fs�0�Q��Z�6,Q(�`��1jWYb+*�`�V+��D͊�� �W4PUR.��TAG[�Q5(�l�\�D���V6�9����U�#,X�8�X�)X"�c�cRQ�PQQ�lYZ��¢���"�1b1�b(*䢈�ADQ5��nf5�jV"�#���Z�H�-�1��Z��xŊ ���`�DED�q�X�ELխKe]ecj��u����kEY����h���-��Q��ET��x��׽��x@����5��RG�.LR��Ҭݤ�c�Y?֦�',):43y�fR�Iv�2��I�O���Q+�1=&7$��r���4)��VM�ګ���f?I�G��b��Cg�!F�P��e��F}!�dѐ�pmï�?<�Q�,�
ɵ�C��G�Z����=B�^
�j��j4幬��$��~} �������%�8�w�mHD@.js�_a��[POK�j�����[8=�_n�cD�C~�Dp����cض7�{ݥ-�!1T��H���
�6\Yv�s䪜"A�9�E�dy����|G���P���E�����N�6����7�n��f�Qܨ��ZS)��'�.�	�p�<pHA���w�	w;�N���{P%����6��B��*g:}:'��)[T6*?<($�֚׹��l߼��^ 5Gݴ��J���dU^�P��\�O2>匚;R��Lu>��^�7���hk��R�R�u�,'mk���s9a�ܷ���^�����6=f�p.ꢚpv�� �tۣ�y���'\�'l����2�ٮ�����XB����v������A��a���\R���B��쓉h�,s:*�.���GV�Ca�^�^����%��y4�P��
z.�K7H������n�ԡU���=�׃m��d��������j*r��S�����Snv��<Z�G]v&�W�q߰�D�W�

G�;R*���5�nT���羈3�[i�o��B��l`p�:�t,W >�O/x��jPT�����=�۷���'�u��T	�#T5����
îr��#��ڞ��Ex!Gj����Sԕ�����Uˎ��M���q�V}���ΐ�ľ�`T��K-3Ś�)����*�0�'A�3�F'WR閻{7�e=�e@Q/(�)�8S>�L���8�r�\P�3)^Z�V�����Y����;zٱ�g�Kz��~�ʽ��`���Vv��R][̶�$ �U�E��#ȣF&�}�¥c|7�{e�n�m�S�wJ���-�)�\j�1r�h�5k_�_W�}yŧ��v��O�"�G	�f��W�(����r�]��6f��YKn�3���j?���� �hAC~�_M>�����GV��������d���%�AO�������AD��f��{-����=�'V��x|��U�XxG�3��/���L��o�
F��F��G삥��}�ЩDU_�%�+�R�{�h�9mw'���ᓰFH�NVaܦ�GU������a�����<�7�*Z^�%�>D+�L����)L�Ȭ��W��tk�� tW��]�Xu����g"���t��uϨ�8.K�.��y��O�ʶ�-�����T>���ڱ�7�j3eL�� (�R���Mz�v����;b|��F��W�z�Mvu��fq��J�W��^���T3FS����5��h�Y��:�p`��18�5uJ�h�\YO7��Q�ƴ�5[+�{}5Ȣ�N�,M����`�S�o0l��d!�`�H�i�7��ո&i����|�N��2�}�U��|p��>�V��k*��
�BVr��^���W���V=�e��ía�U.E�C"T���d!"�p{�U�p���˺�>%��A| 0p�7�^\>T�☪cO���m�Z����y��Fh����Q�Y^���>���֐.�
�*#n|�u#��u��_�nV��`�ch7!@����3EL����/=cW'9CXձfv��H軑��ӎЕ��Ѣ���1�&1����EHs1�cӲ��S)NÊ|o�R�(Fq�$�j���������zM���x��w�K�=�����V'xXX�ռK��P���v��E�d�.���!~j�V/x֊�Tٌ_??MՈ2y�w��J��l>�O%ֺ�¬{���e����߇���ł\�KV�a���Gu�2�d�&�)�
i��m-<�+4dX&ɮ�DZo�R�/�4��[��k�ݬ�sb��JL���o���1ciW�[���2��0ۊ�G���6�wRNMB���X�&ҜR*f�}����Gk�(�����ox�X}��e�P�k���PIi�N�2v�vh�Z鍒{3�M�3!ԫ��E�0d��C������B�����x��F���"�#EHw6]X��"����@�<��o�����R�W�	f
T�W�ʷ(ԅ{dR5�'X�m*�5N���p+������P��J���.�u/��Ih����Y�9,@ا7�AXہp��V"F���@�
��)dc�:������Y^{6�G_��V�p)Q�>����1Y��E�-d	S1���c�ܘ��h��gmg���܀_A.lZ�����e��"�Q3b�PS�
�6\X.ãX��U8���}��fq��}��Zܔkt��t��{Y�.�����ή��Gս=�VO\�M�ïl�!�+�������ۗ���8a�32�,��G0��PG꾔�d&�s;Z3�����j-�zӺ5g�4U`�E���T�>0�����X���=�����CF���4�Mp�<r@ghL]��]��	�=f�&VZ��-O�����LE􋙠�º��PdI�������#I�i&��7���!=L��5ؤ*�.2�%�p^�����Ү����kmgW�W�p^4���Z�N��"� ��X�z�2)��b��֑�8|*���xՊ�,}�P�3�Ǎz�5O6)-(����!0��]m,���v1ߨ\�/(���*�k�;xo�I��#�8U��!��@��y�ʠzj����ۢ�ؒ�9���*�q�͙am�УPѥ@��Q�g����� ��H��C�6􏧞V1���KM�cE_>�V�R��F�S����\�m��0^��\9��-���u���ެ�T�E�5)���}>0X�-�6:��)~��I�5��)�Be8*՝s�i��˔�aik����*o	�G_7Ƥ[|�k����#sا�����z��B����%�3�xJ�W�@�G�J&�t_s{��
���4/���GE���ip�R�����9��i���ԯ3J-v�C�� �U�>��Щ0s��ӿ]J���q^3�E�"��c�\p�}����i�
�.
CB��Ú_h�*�C�v�t���]�δ��0ÓX瘪qH�dр�97�K� =�\���v:O"ӱ��X4���zӿRT�\<�����*w�v�G���xx�E(���s�=�U�T�&!�HB������:$w��$U�i[yJ���t����>�����a�C�2�:&V����#����e�l�f�6�ת�������H��vŸ3{=ݩ�ƴ}�Eh�e��5�γ`u}���P��W���E]{p�08�UCl�Ր����ˁ�GPy{Ѱ�kn�[��V(���k?l�gO���]�ǾZ��/�&�����	\��ۿn!}%2�}p�$��k��P��
}������yk߄s�V*讑S!@����c�_�Y�Z�5���7쾳��0_/1Hֱ�*��,]�\̗�ԙ������1�����.G�i)�(z��u��SW��>uw#�(]a�i	��!Dtڔw�g��-ؙ���B6>7�(�s|��
�V��k��v6h����	)��Ҭ�˃������>�
ΣX�b��@���%��6�>�Т�]HWGD�EP�*�tP�lX٥7��z���)͖�-5&�|@@��@`\eiWx���U_ʍ�"6�ʌ̟�zO�fr{�A9��֚�/N��t�~?�|5��O:*
oJ=79R���5D(~r;g�4˹�h��nG)"A�ސb�7�����
�B�'=��FáN�v%nÀ$)����>��#1�s�F��9��-٭_u��m�+z���W�-F�6�&�D�W��
����j��z���Z�Rv����U��3n�eN���mX]�ϳj�JSZ����=�R-�&���`��Ҥ�����/���Q��-�ǧvRW��OZ�GƘ�� V�UĎ;ƌx�>y�
/f*[4w.ꗣx��m>��`F����p}P=5�Z5i��B��,���5Fvյ��o.�aP���(P=EI�A�Op�P֋�dVe�e�k=�w��q��2졗TP�J	�b��K����B�%�ݟh�k�N�Y�������ƸK0R�L��k2ր;8�����hW�� �Ɠ2�+5ఎ]W��;(���0��kE�臢oˉdY��,���f��]5{�/+��vu����igrP˧so�S4)Q���^O@����$wL���	�z�qyDij��&3�Ӂ]��D���	����傓壤=z,��$5���.7xqٺ�:r�w'(����x�����%}-gy�J�Ӟ֗+W"�{KC���>�m�eܰ���'x�b*�9�����l�K.jW��/�����ޤS�t����!�3n<���#fhp�� D��v���Y��د�}� ���[���B\���UtZ*��^~�����y����ʖ �Tχu�j��A�$$vv]���v�#�>����)��I�_q��vxW�]�@�9��&:"��W4��uC"�w��Ng�����/�����Oϩ��B�i��#�F=G�)A*�\��h����=�^:Q��(ݮ|�șz2�-�M5|�H�vQ�.Ӱ����5-v^7Oޡ�R2y��>\�wڀ� MQ�P<0Z:(���w�'��5�gw����+�<� PՂ8]Ӥ������x��5��+<פ��$��|W�o�^�C�8�{ǾӔ�i͞~�%MG����"�$��遗Ӄs:C�s,ͷ�53�V�w6̓h��K�k2��_(Vj��U�V�n�s�p��T�$�����햖AK�v�WKbi>��*�4�����p��@v7�I"��x�T�O��(�%{�Bh;�;v��#k{e	�=�+�U�$2�R�^�{0����/�Ϊ�4�\w�|�:�h𺻘%���c�T�2�j��Ee�{O��J�L�ވ<56�8mU����'�t<F4�n��*n���.;�zi���7E�}�6�
m�?t�V_hVF���9�R��p�sh7�8��N�����a�3pJ$-�Z[��bÖ��&
�z�٭�[i,��\^�*��Z���ƍ$����`�9b<9
�=[|KT�͸(^VU��*5@�:�X��q�,k���m-g�nq����\����i����xbڴȍ�2�yS��l	�[�p���[�<���uQ����o#�%��v��sMA���w�]v2��[v4�,+݈t���ϣs��B��ܾ��6�P1��������n���a�{���Z�Xa�f�p,�.i>�s7�h(�S�;��Ok�Sv)���ƴ*��N]@:�۵@��n�k�pF�5W2�1�𷉠��D����L�'�!����r��ѿv
ӏL���+b1bm�/ �7��L����ʣ�8v$�ښ��l������eӴ�T����,���=�����ӝYo�a-��!F-��Wq�WtӤ�쥜�����w�&*�9�ڝ|�S n@��Q��Y�w�Y4�W�c��8Vfn�-%����;֝����/`yXͷ�睩[齃Z)%�i��Sx^�n��J{��mwN��n>����#��Q ��R�ͮ#C��=�탁���A�#6�=:8�ՖK�ƠyP�Q��޴`[:��p�&�@%t:��թ���s�u!S2�	�qF�iu��w$W�0�m>K�c7o)��/����E'v[U�ղ���i⢡��6_,:V�R���7[�v�Q�.�b�F�@~~?�\lEg��X��A[elE1��R�~���j%m��N�%J��*��[UcF͢�	\�Ȳ�qh0��b*�`���F,E���٘UG�Vk(�ER��֪�,b�)YN6u�+KR��#�DQJ,�n�X*�Y�;qRا	a�*ƶ(���@�"�pʊ�U�l��YbV���������E**�jR�
���UX*�U5�(���Q��T�TF1XqneT��3y����
�rЬ�R�`�QADE�\Q���-��-�L���T2�Tb
�KJT��[(�-�TPX���6�4֖ �T�F/��V�W]�R����UQD�Ӕ�(�0Ub�եTE��T�%b�Y�QF"�X�#d�o�v��~⠧b�3-s�)��ڇQc����7$0��r�V.iT�S�O�.�s9�o\�I &mk�Y�)L�u�C�!�D<�,������S��V<]AP�z�����.��f�zx��E�j�\emg�����~�V�����������Qp��)`G�:��iD��@�T+�&��H�s>�}��l��7�������׼�ʠU���t,U��T*��^��늇s�I9�x�	��}�<"bp�Y8;�yg̙�h~��R
i�����x�C���OYS�O]�!�q��
���fs<�fv�LT �hͫn.i��S)�ђ"�@֋'����õB���&H,��C����������Xx�!���	Y�՜>��� �Ͼ��Llx	�ܳJ
��7����|�|�zɷ��a��d�yc��2{�
�Ag6Ȱ>k���<g?��) �sNz��(���&d��S�2A��R�tty�^����|��}돳;O�2Az���8g<Y2}C"Æ3<�����wZ(�L*p{@��
��,8@Q~d�QH)���
�I�9a�4�!RrO�J�8nf?}���ب0'��2A`|״+ �C�(z������*AeV�E ���I�
�Ml��0�9��
C}��(��}��~����מq߲~rAa�
�2t�N���W�OɿNq��+�sŇ��H)8��2|ʁ�_i
�*�R+�(d�@8E�Y�6��[i�]/��"�`$�P��@��Śʅ�v+sh��fJL
�վ��[x
��enS�TJ�ǣ��u���'��ٟGdΨirS7_@xA/0���]*.��N�xH=u���L���� &�Q%��@����O�՟0� ��>bp��2fO�j�$�ڐY�'��w��0�85��R=a��p���:�&8p��)����y��}���_;��<��N�
��3��@Qk�zʇ���8H:�αg������!Y϶L��"�§���Ä�ɧVoh�V���_��s�Ӯz���߾��wI�����
��A���Hp��)<B�2Vr��v~�"�XN~�0X)^9�|�����i*Ag���E���&�"v*�3u.?�@
��@= 7�xɘ}|Щ�yfg̕N<ج���YY*r���a�
����8H,��^��t�sE ���&d�=0<���^�}�=�~y=#�c��G�rAH/֟3�2�yI�x²twfH<Xd88�T��"��'����,ȡ�%yI�p�Y�&}nǄǆǄǵ'�k�ܴ��j���#�g��� *��d���L�!P���'	'e����&@^gw$Jʛ�)2A��bϓ����2OP���'�����~���s����~E�l*~^�V���� �0/�vɐ_S��'	'�{���S���Rp�{:�3=I��QL�AI�����Ͼ�ǿ�}�]����������u݆O��d���'���'�T<IRZA�ϙ2w���� ����*��<d���1��p�珸9����w۫4�����	���D@��Oi�Y<�Rư3'��)�
�ǋC$����!�S�a�
ã��H<Xx�3�0��C���f�c�JYL��cި�����}��	����
æ�q`{� ��N4� *�>B���B����<NR
$���p*=��}�w�()�1v.龸��s����l1e��jʜf-��Of���=Ws]2�����vX�6ҬU1���SQ���t�{V�6*�!LФc�*QVqE]ҡ�6�r�8�
Qw�+�s� {���e7����#�0/|��)��1g����Xd��Y���l� ��1�� �Y7�P+��C�����fx�Q���x���X����S��Ǐ��ٔ��>;��X}�>g�H,�'�|���8H(q���X,N|�y@���P�o	 �$���+'�$,�����W~7۞����{��$N��Lya�'�C�$�Ƿ��I�'��̓�u���OYÓ�i&:����>����w�_}����Vr�H|m�,:aS�
�u�%�C�0���!�J��2o���W���Ag�����:g��q�C�H/6�2V�9��������>w��u����� ���b���V|� ��@̬;L�Rd�ɧi�$�|Β�g����@�>B����ya�Aa�8�S�
�z;���^}����~{�\s�=��Y�T�	�85��T�3X ���)��I�
��I���8H,�8��O��9�������Mh&a���}��{������ �=�z�*Ag��%C���V �fa�T凬*Ax���+7�L��~rNg2AO̜s���B��}d�8H,������_���|N^Y9L���d���|�i
��g��	�}�pϙ���T�°�R
A�w�0�`�P�%~OXtsNR
�W����q��k�_x��x��1ᑽ!�C�`pws9d�^;�2ACwa��A�N;�NXx�0<jAfa�'Gt�Xn�!�J��|���߸���>��쿬��<O�0�Rt�gw�� ���'���2A�!��_����?2T��Ϭ
����- �N��pÖP�����������_?U��`X�(��+F�����t��0�n�1c�R�AU��+vT�K����8��c��_t��Wk��5֓�w-̵��
�[�mR�+����{ۙ�����@���rOR�����`�R�^h�a�_}� �psL�%@S��P�%gVL�{��rwC��T>�H,咾�[��y���~u��NOY3���L�R��l^<�+�s�ᬜ�H)^�3�'��qI�&��8H=Ra�R
p�Y�=C0��̊Aa�;9��������믽��7�) ��\C���³��W�ퟐ�E
�L�H/�TY=��B���$>������%@^9�H)1��ׄ�������{����u�~y�"æ~L��*Afa�~•�S�<g|�����=�V,�;g�)�AIP�8�Փ�q����Iơ�tY>s�T���}�������������9d�|{C"����~�$>����<��P���g�<yI�TY9��X5���H=P2f~�V$k�Q�� �������;Y__�@��J�s`d�ݜ����*NO�2Agi?9E=d��G�H)�q5���:N~�N_�:L�������8�S�h
Aa��O�����y�y�=H>Y:fa�Rm�,��!��TRx�C����]a�ö����z����Y8@QC���?���|՟2}��+�������<��=}��!���L�+'��!|��H?S�(0�&a� ����
)O���T>IY��ɽ�V,�=Nhr�R|�ܪ�c����O/��.}�@��,9O*��2A�P�Pᇌ+Ƶ�Y�%E"����ԙ!��>e�8a����
�S�IӒ|�q���~�/�|���������v� �@�7�hw�)��d��RT��E �P��p�R�"ɘv¡�ԙ ��q�(
)�&��Y� xD-g�]2'6zg1�WUv����Jx?s���uI=0S�)Ho/�^M�Y����+Bķ9� �6�����f)�KD�t!�ڧ�:�v6�"TҢ��.[DD����_}��w����:��%h�؇�i�"c0�`�Nz�2�W�Ou<���S�3$,</�0�P���9fCw@��t�
�R~=�����a���=�g>��\�L|$�Q�P�s�',
����2y��<;�0�*C�O++%a�*�Ad�����R�o8!X~g	��vL�c� ��;xw��w/�}�`" d��OYP�%s�d�Y�T�	'W��{d����0��y����)��d�Vg�fI��{ "x	�5y����F�ٛ�=����Æ�B��>�ǊNЩ6Ӥ�9'iQfd�ã���h��X}��H/��<T���TR
�'T8H,��Ǯ�o�^|�ξ��~�;d�8a^��2Af~����7�/	!ͥd�y�*~�Y�����0�ņgL�������)!�;I�*A�g?��0�P�;�~�����������> ��z��
)��2AC�͈�a�Ç��
����� (����
��3�O��O����T�� ��J���w�:�u��~����T�ö��P>�S~�+Y�o� �{Ň���N|�������l����zÄ��tP���&I�Ȱ�O���]Z���[����� xA�� \x|¡�J����������RZ~�+·���*~S3Ԟ9')Q��C0+X��H9#ʠf���yq�Y��?n|"�s�Q��qrAgj��Nl���Rd��϶o���0��^
AM�����x�{���Ad��2t�뼤_�	������xT�t	+p��Y]�{�'���|uc������*A��Ł��
��&H,�s�PX��l*As`n,<a���H(z��ϩ�&@_8�y�o9��;�N���{��'	���ʔZ�����˝�U�ڼW�v�׺z�Fh��H�QfiQ�m	;�L�:���e5���SR� Q"h����fΉ�386tݎ�Xo;����f2Yo�>�`zaǀ��T�̛}���:aY?wc���{�
�Ag6Ȱ=k���<g?��) �sNz��(��,�G��� 8���D[�������o�Y*}���:a���=C�~�ɐ�yC"Æ3,� �;m��Xt§?P3����2��%h�R�P~��L��Ik��?,nǙ�>
�}��u*��"A�s�T$ԱB���{�s� nHfq���W5]y��80�D�+�oY�aGU��Q#%��W����lUe��4b��AO�x@�%��t�^��{�݃�G���J�*A��0K�_�#B�J��`׃��/;�+�<��W���N�+lڌ9�x���	�M��B�.��r��I�ß
_>[��*!i|K���u��;��;�cy'�sU����#����4�+�PQ���-�ɮwuf�ӿ_'<ot�	l(FF���ѱb0(kE{F�}�EY'(�8��6�^k��'����0	�Y���/�K�*z���Q�o�,^ז'���L�{���3��M��q����ǽK���iV�r���;��Q���{�L�Rn�ao�~��}B�X�����#�b���g���ox@B�]-��L�>�p��P�ײe��/�tm�)�{��+Ak�y��G�2�e�~D�!X"eR����C�W<�݆����Q6�BqP0V�Ŋt:dr$B��ɠyf[����/Ƥ�$`�A��iWR
�Xyg���AP�zB�{/DÖj�5�|C#��ܕ!<�Չߌ�<"�#�>p��m�j�x��)9��B�b�Cٸ�9.v�vCr;�DD�&e�vMs���#υe����(��[�~�t�t]���N9*p*ci5W�+�{V��4�O�W���;�����uO|���o��&��z[k,t�\"�T&�!GH�kIs|�������b�*�klc���!=��ͭ49>>�`�*4�a/&>e��=Ӄwx������-�z<�3L���k��_"f�aB,��vG5�-L�.��ӜYq9yr�s������Jyy%}�bzH����a�V=Z8W2E5���t�;���sWJ>�S��3Wc�F����T8Q�����9�3�Tb�;ɬ>7�W��3כ\e��˪?!I�	�b���ב]��O;b~{L߀���?z�~;K��[AU�S�\�,��e`�N.e=�3/D�LR�S*=Bf܆�ut�T�G.+ū6�No��&�;XkI�Y�r��z�4�.�V�^U�ԫ�X�x������V�f�1,���R��\�>gE&j�W�;��'��r�Iΰ$j�M(�����T�q^�%�f�l���l����9��a��65PV͸
fpB��'Q�]�W^�(�xS�δEqD�,ݯL�����c֖���5��:�*�j��.�uk����A���#Ό)�Zjwe��Ƹ֘�����yfGn�(s4�7��ޑIJW+Չu����:�R���v)��vL�$1~$N����kW��
�܈��{KL�I9r碡BD;�Q��vtk��%�dj����(��p���0$)�yˇ
Fq�=Gg2��,MO��(P t�t@�� X��W
�7�J�7o$��(�0��3t��	SaO�Ϣ���#��*�F֛R&���������v��3�L4�0a��-�]�e����7я�?yN缎y*�	����P
� ��0^-��[�d���뀞���ʅSp([V,C�R,d�8��GLE옓��`���q����F����ャx��߯�__Ӌ8�ǜ{�9B"r|���I�;�2�됣T�=T'��ut��#���7T�w����!ۍ��i"���x�v��WH�5{B$q�>;@٠��9<��-���=۝/`ʳr���E��tH���l�xS�7ȍ����'c*���k%�I���D�O!p�,��p�gGsy�1=��S �\�_}�}_�z$�����.H�_�J&<��p�4�-0���D���Ƚ�{_N5֜���u�t,U���B�'Z�H��R3u ���M*d������Q��YGàg�G*s������K�X9V�u/�����q�����t�2�B�f��U�ٍ��ol��q��&m�hV�r��
�|`���y|i+���zQO�dq�a��"�;ʜEDѡ�683>q��k�W��Ng:�rj�;7�P�T� m^:��xH��=O�`��7�i��2\ T��2����C�)ߨ%N/�TH�Dب�yW��i`�1R� A�26�'8#���ƌT�
�*���{}��k(�����ҡ��<򢩪�����}!x~��Ҳ8����v��T�����Jb��l`�Gfȓ&�j�YQ t־#��yyǜ�{��XJ�6+w�`�8�X�d
��v�x5[�2��%iX�tqU����7ӆN/6����;�W�R���£׷(�0�:���=:��`�[,&�^�7j�*�C�b�\-������0�(�&ii%F;�u��d����z���(e����-����U��5)��KY��ǔn�Q��+0#%�#)��\������Nm�{}5�O�l��o"jJo�`�f�S�w|hć����k��Q��@����"�����,�X_CL�A�4�i�7)Rf�97H%kbkXv�SW�B�R̆��&^7�`������ǖ?��	Z"�>)ҏ;tV�Z�]��Xf��aĩE&�����1�Z�]��U�(n�+Ԁ������ހ�mr1�OKbat(/�˝F���(h�#S�ϋH��d�V^�L8GV�b�U��͵7e:%��5>ONJS�U�!2�b����l���ެ��_�~�1e}����B'fJ.�i�H��ҳv���`�/e�ХC:�8��`��S����%b]��]��J���A]�o���Fk�u�6�&�_-H�Rވ��y�;%�r�[;,Vm�omMHHT������+r�W2�fHݡ��nc�\����2�eƶ�5R�`�ظq�D��5X|�^��p�\/N�leܶ��F���&�������KY�G�t����R�=b���&�T��l�v�:�;x���H�	ۉ�P�t���q��֕&�]������vZw�.��H����R�c�27���s���5�A�f$,'6�q��VtY�ЈbD�
�w{g;&,s���s��_V޴xk�;ZGi�\�A�mZ%k��Y��<ܣ	P��W(0�������[�^Ai�`6��%�������Z���Z���Kg{\X3��W
���+�5�`�Q��V�..l 9�y�������qo�gL**b"��QDC���AV���(��Q���Q��Eb�1E�*��+YT`�j�	u,X�L�F*�A2Tb*'QP��DUPDQQ�8Kk���EXV�U�TDX���qJ(�����<P��V,�J�&i�X�,X��X���V����ډŪqlbZX+Ŭb��"TX��kEE[J(�����,V(���s�-ku�b�" ��`�#[X��APEmx�F1X�X��`�b'�1UT���1�,�0b�ګ����]x��FS}�쇷�Q�n9��A}�v�:52"}n޹VzLi��N����gW�܋o����we�/��FT�͌u��	�nۛ����løKp������Gk����*1�"-��u��v���*9>����X�+ܿ�h��6�b�М~R(4Q7�+(z�
7�ڄ��F�^�B���e<��Uzk��?�kE�F�!��Y�W~Y��v��>G����<4��l׆��_s�%�`��5
��6c�j�e�eL��pRÚP�`��>V���`���a^F.2��MoR4ɩ�tMX��:�O�<��O�x���`��poOM����JQ��N��@�XT"H�����T���-���q���>iOf�f��O���n�3beě��Hڈ�renotn��4�'|�����}�_O�H}+��b���NM��z<�7U�OE5Y�(��m]-dX��_:���1DiF7,@��쾒
]gc��z�uȺ�|u�-���l[��{VF.�`e[�vZT�z�w�"��Y��ѽ(fژf���BI'jW8�3�Z&63xw��fbT��)<�a����nB�2�*s�G
W�s�ݸH��ѯV4��GCrGH���N4�ʻ�d���VR�� �HT�6DD)q�������8�\hK�
��)�^�
�:�8И���:f�:^�����Gy��^1{=��=C� ႑c��h�\�#V����q=<�`ٿ5�G8�
�*j�WJ4��&>��Ī.������\�yP���ڤ���R�Gb�~KLQ �7��I��<ﶭ߀�S�}��_]��٭����X��S�]n�����|�S깚H��`�1�S�܊$@�d��9t�k��u�s�>A�XO��C(����x�|��R�N���%@�yu�X+��tD��gqf�Շw5r�tP���Fm\�$LXteۆKH�"+kZ��*ͩ-m���;��#v�N���#Y$�}�)�F���� ������HFd�9MA��������ܻ\�}]�*<���|�^j�K���@Q����b�vtU�A�<[Y�����74�S�P��.�f���\~��_K��6b2�H��A����_R�RP���D��!>���AVK^�y�O?t����%
�5�q�����-?>�Kw��ਵ�^#(��"_��aT�#�@t!&As1뭡NiOF�	c�p�kn)_��Y�<���Р�܈�W
���Z4���.(gt$�p�Im���b�:���w7�|hQ�����oו
��ՙ�l�6\��e�*bz�7EtS�r�X��p�K 7��|oFP�;X@�P��5,E�4R&�O�3�<֚H�Q&KAEG�ڸ����U��5GqA>�L��3aٖ�+��}�	�I����^�+�n$�0�����F���Əm��KO�����e@���ct�.:�@î��4�f1eN�ptG:`C�j)���{��M�qi�nB���U!^���:}ΝƝYC�ᩤ�;�����x���1=�����TDfK��T��s�M��CF̋.�6Y�%m��1�P�z/��_t��<`j�Y�G!^;��+h޺����쀁� �@o����U�F��] �>Q�3V���y=ʌ��&(Pz@�J�L�>�B�L��
���{�[G B׾K�MXU��eyTN
|xf�б\�^V<��g�K����(��R8F_�Y��\*���F��\������o�Z"/�AR�ƅp�IJ.��ɕu�����3���m%=��]B��X���6���+n���+���_Ӕ��39�{��R�۠��Ҕ���I�1:"����2��*{��#��MsPn�-���[�I���gqYaX�y��d��<uyeo��a/u�7[j0a΂�VQ�#r�BJLn��ݬ���٥^v���������W��2�`�n}��2,ٷ.OJ���ǰ�R`@�D��*�\k���ȹL��]R�N��W��_��>2^1.DM�A�S�۾�/sDX�0��L��NE9nL{b�e��.��w��M�i}��׋��!�ʉ�"�џD(�t&��S{.-H�Xh_9��e��~X��s�Fѧ��z܁7�_ir������P�2;i�
<G
��4�MX��X�'�o7{ò��W�8z���x���0`�uT�=Ż�9���V	��P꾳�ou= ��BF�ȣ#�DN���ՇZ|Z�鏻�� ���;B��ھ�k�i^޿`�FgI~���>({O������S��������f�����w8��=�d�G[2upa@��y1�M-��ڣH�-�{-*�c7����YvoQHe�JQ���Bӓm���B��ɗ/4�{rRt��+����R\f�6h�߼=�����6��>C�	���tF�~�8���&|ʥ�<~�&YҲ�d�SpOkcT�jaH���+cb\��T�
�zw���N6�V�޴�u�*��Ĺ���e8
à��8�Gᘀ��(e7�x7`����k�C�ה+߾��*��������������'ٜM�u�ͣ}��~�ds!+N��0OG�I��a�����C�1Xl�k)��az�0�P#"���u���rzGEߧϦ��s�t��:�7��E���SG��QD0����x���\"��N�ϟ�ɚ�M��͸��Щ�=���PQ��Z�Uo��^���i��yau{"���C�
(h��]��r�h��i�^}pב	����O8�7����*�:Q���;���H�=�	��wnMМki���=�����|pzo��m>��[���"sz�h���Uwo����Z_�ډa��lO���3kN��w�Ս3.�G2s��d����Os��7�j��k�������o{������a�_�G��/��:D�=�L�<K0a6�4^Ճ3�����+a��S|�uix?���V�L,Y3}�gx�]�)_�tr ��Wuu�K���W�+������/�cH~���J�{����U-Wb��(-�j��\��N��Z1^q�X�ѝ:>�}��U����������b�8�һ�kv�06@&F�>�E;�uG9pr.��:V�y����}��=�n��N�
���B���tJ��A[6�X�]\��<�M��fp) ?L��
A�n�/'�C+�e��Pc��[5�ډ]�uK.6�X�G	���T��C�S��*u�=y�V�=i���˂
2+�
���E9|0�ȵd�V>b���V@콲�UՎȺ�4���ۗ}[����ZA
���%��'�ݹ�_$c.QS�Kw�X�ʷ%���VV;|y�̩�b�T�_{&�	Iڸ��P�]�M��ܗ�q�F(B�>��xle�df�B!v�g$�5�W@��p/�*@�;Mش���>�>�+��̗�Z[>���_��Z��r"�g���eZ� R���
���f��B�ԫB���������T��\���!7��٦_�+�2�(�G��ܱfꚡ�┋5,�F�:����7��@z�|��F�6�����g�3�V܉joi\s���\�ß:��E	�~��5WJ�#��u�0sa0'�z���g������P�q��%�FkdF��P�!��OK5%FT��qV�����N���?���t~��6r��i�`�Ɖ�3aeW�������W�@��T<.��x:�����l�{�o���"�+�e�:�ҶٌH�-�f���=8v��S.=z���CT���{#`��	�ɻ��6l��&ԣ4J�8t�	:�w(wUG��}���k7�o��������(�z�.}NC��r@�����I��7����)\��b��Lp*R�Я
�IJ����gE	)\3]���4��䰺��.G7F2\�蝊�#�ׄ�Q.L�F�=�U�y�]~��HQ�-H���L	���0#b��	p�P�q�&���ꠍu���V��pS��]���h	�s��6�9�l�������A���_�n��l��^w@Y/�]8So�[Sq"H� ��F�@�$��T���YA�xh��������g���q(��+�̞|��^�߯ ͥh#e�s+��߶ߪeUl����"���YB�?���h�~_30�����<�X;|� p�p;e)�Q�8S�Y�K�=�=ժc;/|u&k*�=�m�Q{2��'�DvDtZa�ڔ��j+R���4k;-��#(w���2j5.�ÆYZݾI���7��wm�J}Ҷ��9�w�Hh� �߀�7r�I�P��Ȳ���2n���T��1�"��#�d��-��V#^�U����곕k�U��xX�EYB�̔�������e�?L*���_>T��wj�^��8��ud���~O�)���2�)��|�|.���t��e/4W@���p"2߽�"}-��v����`��.�Y��5�2��r˓�ܖ��(�b\�~Ҳ�^�=}cZw���.�'��/s�㳨dOK��e(
á�@�3(/��zm�����zw�1�p1�1�23��P94��!���W���N������z7gޭ�}-��5a],� �!���_���{�\܏5.�>��Z��4Y�O%�3�Pl�N�&]����8+���a�-�>�3�,�	ո}��B�?'-Y# ��u�U���C#�ïmfHdJ�p,Pk��䜆�t`-&`$N���GF�fGt2�S9T���;�x;DS:j�?#5�����:�Τ;.��ӻ�a^�-h݂H�WfT��M����Z;������%���0�����v� �<�*[o������gVl%�+����58Y��tZ|�]��)u���{[4b3n��+�P0j��jP�Y.q�z�n݂��F@�`W%�E��5+�����.6����tؾRW1Ϯ� ��6NI��k��k�qʆ�Eӄr�Ä�ה�R��V
�y������c+���y���m9��J%�-�t����{ˌw�t���t&,���nm�	P�m��'�d�ǩ[zQ��w*���Fe,�uEoV�;�$l����I�����x�f�\�MAI.fg�q�3�������nQ�G^>��t�l����$�q佪<��]1w/z^t9V^&�;1WNZa��j�����]W����k/�����O2L�[alH�z�(�ǽ�4��ƢũcG}{Oi��@�*���|R]�1���()���+����Zy˙���\�ma f����M*��4����Z�Yęu�cBB�w˗m]������m
�ts���FzS]�Qf����b�nÎ��λcN�\��Bb�s ܺ�E]k�6,���D��\���?{3���n���d�w+�j�F�cE�:�^>�l=�*TZhS/3�И��(�8-�t=R�`���{�;���e��1_@�LN.}�|E�+����[/D�)RG�Y��5=N�1�]����}����:~�A�[F��֮AM��/5g]v�֎��:AQ�_C��"�wE]���ķ�vR*�^�����XĎ�2�^��ZXM��+W/c�c�x����y����kvv$����j�
�k�z�0F�X{��Þ�;����!�,m���h����1b�J��QPU�kN� �FEF���X��"�*1Ud�(�����UH�*�Db��,Ab"�b2"���E�+B��b�+����8j))P����U
�,��V#+(�)V�)�QEx�Q�*�E�3�J�ȪX��"�"��TkFXUAh¢� ���DTAV(�R��UJ���Ub5�����`��]h�UR�:�;��~w=�v&̝1���lj`�����*ZR�J4d���R��8vĿ��巚�lߊU�{���0) �dUp�>\���tu��^R#wF8,�?��\(Ⱥ�ب����(�*��T)�U��9�q-ABZ7�����d��򣣧�>B2�����{���[�M+BL�T�W��Эi9� hDN�B��)��/�]]���>O�dW�(N����#-�Qy�:�4&- ��Q�k�E�t ��	f�˦s��j��*�X�"��@�{U�q���}{�܇���}W3\$mh��ʏTͩ�ے ^F��E'4*���f٨>��)���T����
���ە؛W�-�G�yO��~���]H�x�!ƕm%���w�{���̨:υ&~��ʴT�+�)�����r.�*��k�z���uգ�@����߮{\'j�(b��[�0twW������R](�B��ߋ_�K��Ԟ�����b�G\�b��sVR�o5i���_��}UG��E�b�߄�Jn�@]l
��̅�ъ�b��HO���͌�݂�Z�y{KưV�TP�MJ�ET��;?#Z~|3��W��E��n�~��������\8ʑ�6'���HD@Ns�>5����Z�
��Gx��^dv?�X�p�(HHѢ����\Oi�ih��Ɨ�Q%�^Q;;\����9��v�p#B���}�;����&�޽��RT�ҁ��GT�sb��iS��0�7�Η}���7ɬa��T���������]a�.Џ�J��^�ۃ�J��ש?i��{G�*Q��c�D׬߼>�2~����.�Qwb-s�{�]�*�zFRJ�����X��>��C�R/�5��������ː���B���~��U\%렭P	]�H�� ']x����|�y�^+�}�Q5(U蘺D�Ւ�p��ł��#�2^vV���o]�\�]�@�\�fN�;7�s_qJ���������t��==�N��4��,N�_��"�p��K�W�ӫZ>Tx�[�޶~���m����Yg3��u�׽/�����i�nI���D Vu�!�b̊S]"3���R�g����o�$���px����/Uh�T��ϼpHj��˟�D���l��Ӳ�"�WX�P:mCe�Ee`x|5�/�yh�P.�]�����<=�����zg�/�76*BW>7;�@D,ȧ�(�s��ˬ�2�ř�(@��3�$O���H�B�w�C�I)'d?)�7�����Xn�b���=�^�#�μ:�����V!�x���DטN�~��-�Q�-H�bw�&Ğ�H����)�j�ݾ���y/�Tj���].�����ax�qH����3od�ت������/�����00�\�4`���r��(El�z6���9� E�b�2NN�-Ԗ<�����"����������#@w^���o;%3��H���)�	�n�|sYyא�.r)ײA�L&�f�0��M�f��gbDPr"xW��cf�D)fFZ���\6ùf�$����'Z�cORT�EK^\M�a��ӛ�A��4�h�^���%��+�77��鷚*����h�����_��j\�e#�=�'r��kJ�mѯK�	��ٜ�T�(@��IHQ�
c%F2��Γ �6ϒ�W��~�%�6�p�ո>�IN7C��q�d��l4J3`TՇ��j���q��UG�(@��^��^^�
�ɹ�yͮ��R2̰D��>*U#����	�Ν�C0��u}�<6��,=�+݆���fj8l��O���H��[�!VM{ �[��$���e>�;����AZ��6��늰k(�F�>����2'k<��W�:;g�d�7\(�}�!.A�iYL��=}y����q�]*������޺M5]7#�ɗ�ev�I������٨B)3���Ц��&gj�-8�*Է"���sֺ,�1�N�d�ȭ�Y}(�����]�Gh��=����ēv����l
v/f�o'Բ�΃S�L�?�Q�;�Ɍ��k7�G�~����b6�*��*�=W���*
���g�����j� F���eMc����?O����r:)�[&=�Q�8�a�U�7m����=U�i�x�!q�ƸtML-J�.�rṁ��OFdD��^ތ�B|��FeH�SP�YF� S�`��}/o����}��Vo!���ceŬ�P����BB��a��o	/j�餞�y�&�/�ǯ�{"��6:�!�F�@�b�T%�y3��w!t����6��\g�g�]���Δh���:��+V�7+�3s~2��T� �w�XWʓ�|�^��d�+Λ=5*�c�@W�ϕd�����2��K�7���)����Z�`�n���w*a�����h�y��5];���Z��k[$�rscV��Z�S�3V�)Ğ�8��
P$iQ]r��/�1����N�{��4���yԃo�B�Z��jd��Y�|*ɾ??��/���ѡ �����`�̂"��o�!Ǫ/������Ln�T���!8έTڞ�l��/z��Mr�۟#f�֪�	�a����(!��7 ���4�Vvu�K�^����tg\�6:���j0�P(������[�vȈc�P�$́R:��WN-�5�0��*�t�.�جy���Gn� ����GP�B@"���O�'�gN���Y����h&��%���Fԁ��pt�D�c�o�T�yʉ����N�rnˆp;��5�ȡ*DDX��ח�s��I�p�$��^᳧��������w[u����v�s�H�dŀf �P�ڙu��[��LUt(���8��X��"`k���%,G)����ˤ����ɺ���V0�{o\~����f]Fq���fz4�-v�
b3�(���n��SeIa1�a&���t�0l��e��Y�c6�.����e6�p��#�nX�ِI�����Y���^�?{�>5 t����v�uO���̎�rg&�\����'��{M2|>)W&�ex��x��w+TC���ȷolջl�-혅��,�>��IV�������ʲR�i���Z��Y���7[qy*�i�3W�7���nR���>hߎ��I��j��v��ńo���nO����8�r/���0:�<x{ugK
�i�Ɠu�F_�T+�~ܗ2H�
��C�I�c�F��<��Z��>z&�n���X_*Ѣ��MT����I׫ޚ�]uv�����0��=R*��ܓ��-*��>*��{O�����^����!�,T㤡Ugi{���u��2�y�s�jX{�o9���9>Lo_E��*�Ѩ��AR��+¶�)AW�vo���r�`b������)*��PN�*�W6L8������lO};�o|�����ػ;��P�|�ȕvKtf�TV��a�hK�F�zcd}?U�q��k�)�y4��u�Ԇ�̡3�&�"v+��s��՝�;����M�P�n-���5��g�pU��i����u c
�`�ż��ӣ�CG�Ot�܍xZ�\��!�|���~۞~F%������kO+D���O���b����a��珮(%�gG��JvG�����>+��xz�Y��*?/��*�>f�Z��#��FRݚ��)��e)�rh1ռȲ���VT���BG7���n�c��
�C�y��n<���ol}-A���Uӷ]�U�˓.����B�	��U�3�[�$�Y�oi�]c0�`c���Uw��s"����g�n7wlu�l���>��.V#�͉.�J��ڠe�������GE�Y��#}�U�UQ�J<64�5��[��z���d:�նK��͠J�9���_`���j�9JoPd�o.��ƞ����s8����Z�96h�Kq�4�O,��3���57D��M�r��ͳb������<%��wG�6+�_�����k�B���/�^�%�\6��≱;}:{�� ��죭i�-\�����O�b���T2k�3у�32�[l�A����]M_/��Zk�p^��X�LP�P��;N"�;�6��y�֊�{4�~c���K�^���qkBͨ�T������S����+<MP�m]+?OGN��/�?.�»ƽQ>�盓/	���<�R"8C�U��Ǫ��ʂ��n{>�������I|Di[����^�4s�)�4��DA�U���2�&��<B�edl�;\�ي��ɛ�۰�m�Xy|k��8�S������)���y�����W�d�QE��7N;BV�� P�DUGH��ً�Pm#�Q��[
"S�*-����%,AR$�P'� �`���x���h0�ל���2�+��V�X���e�±k��[�����3�NE��wx���9mM� bA�d�kn,��q�Tނ�Y���+y%�w��t�2e&k��5�ed׫���ݝ&Op���m٠s�_����#�޿����*����M��$;ݹ5��]d������@b���+e�����\r�}o
M�f=�n�T
Q��߲3�v��i������xCy�҉��ݻ�P��4�`��|,��k�M��ե��S���M9�"HM�B��p��jAT)e*�]]�>���h0s�"x�~��5�(S({lz�x|���P�f�h�{Qr-+�8��eT�)�E�bC&䩰���7�j�	��o��3.�2S7�d1©D�q�'�P>آ�te��GXڵ�s2kC+��{ݥ��S��V/��дjRk/��E��pvLo��6'�KU��{X������1�B��$l�(@�E��6�}����k���uW¦����?\e}����e�Z��|�+2.���Th즥��ơ�i���Y���Qm��Q��Fpl�\H]�������Gi�����p�Fu��o �CI�?.��L��7�h`�\�B���|T���q��[��f��l�Ď��u�BU�YQ���-��4d6Z�����_�V<���_�`<u�H����Z�a@�c�\�������M�ڏDQ�;�L웽s@��6ElÎi!vQ�#nӢ�X�J�TR0ެ�D����yC
;��;`�(jhm�����ł�ź��Pj��8���P���ٱ�ZZ��)�H��,'p��nm>X�jpε��h��`��BI�?XB.�6�\R��
bu�j�^DΣ0����=��"� ��d�ߛ�(0�ԟ*����S++��m�����YfU�ԕ]�UwkB��M��,�:��\-(Dm��V�LE�[r(�დ���{I;D�������9�ׂ��o�5�I�����4���tu�@��WJ�l%q�r#t��]r�Ih�.þC\�;IQ�J��2����
��ђ�VLt�ӱ����zO)�՚f��ƂY=1����fݽ�ݡS��B���$�	���:��� ��'�[�D% .�Sy��̎fc��hۚ���x�-G��\�j��h8LX��O�԰�j�َ�˛�C��^R�JV2�W!��;�Ha[�����N��X�ٹ�� )�ǴX�4^E�Ӵ� �P�.�9�u�R��,�eF��q��Ou�Wy6!�V(�)��ϋT�!G5 �f4�� -%���F�hdm�����K��Ɣ���%��n�i�K�X�J���c�0�O/������׍rk�ܺ0�*#��/8ޚ`��k��f5��0�t�&�!Ւy_0��T�:grW�4X�vY;Y(\�4<�R���;�'i�U�2M]Q#@��/f��7�y�X�����o�y��DW��T��ͪ�2��D�QABڨZ~�QV(�**d�����*��(�-��mQb�*+QA��b#DP`�DkF*����)R�
�+eEڂ�*��֊���Y�LR�"��1b�J%@U+*��*(�Ex�ED�ʬrX�-5�Lk�5�
�u����-�(�����"��sAũ������V�x�AԕDTUu�ʮk5�k�b���F�*��U�EV-F���
.��7<��s��*W�gJ͒b�4b1�cΤjnث��`��lQ�|�7M��̌T{��QI�ǯg��;a�7Gc1Yf`�4\e��E[3�BZ��y�t�����p��S>������<��DA��O��r��2��hl�{�..�Uz:��.Lh�P�]�g�BWn��F(9����N�@#�>�i( �W��m8��E���n��a*b"���-���.}[:|�H
Vځc5ی
���w��+UdD���S�b5�Wb4e�nn�0�&!��0kMb��e��w*�l�դ�yu�����z6�]a�h�4�m/�aP�]#b��|kӲ�N�zu��kС�:*T M>T���GB��9��WE��r�����&v&�Pd���KH�<e�P1�N�E���I�O8��t�������G���oh��*���6���975T���Ck(��Viqu�[+�F�{E�qQn&���	e��.����T5$���Wמ	���u�>y�uy��Sڡ���Nq�Y5F�h��%��q�0�ӿ>s_��d���h|jP<0��]5�U�MU�Px`��J��=*+4�"�w�3O��HT(��3a���ȝ�*:���T�I:x�k*&7<zp=��X��:JVj���H���ҢC0v��t#W��H��4���lw_ǀ1���F�+RR��'�9�y?p���X9���B��zxǀ�U���Rqq%�Y�w��;� \0���o���1*S��!����i47�K��ov�׬��0F����4n�2�t�ˑ�L{�:$ek{�u��c�@�@H�H����y��X��aƹdу�R�w%��m��	�w�ΒpB8l�6`)fi7P��QbI��i�ȪM����
���1<!N�	WJ��x*=���ψ#���7�K���zQ��%���"�ۋ��`}���$cX��X���6OF�ˁ�h��Ƥjwsq�#U���Y�a:�y˴��kG>�d�럪�o���?:�sϽJ[���SD+�(zRI���'jK�7�v��bn� Ejڕ�Q��bﷸ��]z����^�̫mU�r6��*^��8bwRX����Ltą�8'S�g9�e����+n�NUY��V�8�[��(�#j�6��`�}�3���%�ܙ�|J�l��׎Z�Q�ఉ��[ӎv�\��=ܕ�noƧ"�X��6oX�Z:��u�Mu�mG��`��\p�����k�[��]+ܕRb���S6.ܭ�O��\�ѓ�}Kzͭ�ҝ�i��R��ABR���Kr���U�\�m�oww�P��v�x��P�]��Ԍ�J޻u����l;F-D;̃���g���j'���w}:̐4N{XY
��ؚpm[�r�M`��I����Ku��Zs]�i~5�߁/-��B��!�"������8m����J}w��.�v�('��f��DF�Vޗ9z�����wX���ٷ�4��pHv�dL��Sء)�֖��*���];=P�L�J��{ܦ�;Z�n.I`�%�
AؑX^�;��s� �so���q��YJ\���r����ck��7�\U�ډ�n�ujK��o���ɣ<�nk.�ۥX�3=�S{��yz�:��4�.�4�ռ��8^],�.�1�'�\�S�c���k���T%�J�]�{�ֺ�].��|�k�����h̣��ά�h8�G�&����S��	*n㢅N䉕�:i8����[ix1ӯ�ja(���S��N�L��,V7C���w0l��`�42��"�9j�*�	����ԛ��j㕳}դH�ޣ��R�%G[��DJ��q�.VW
t�<�5N#Z��f�t��{�N�Y<Z��Ƣ��bF��H�٥�f���}�`����)��s-K�s�Ѥt�[3O��۬�5y��7/�M�ݩu����J�F��y9��lb��ތI;E�dT�t����,N��$��E��3_=����҅��3���=��z���ͯLf�GsM��9��:H���]�k�-�v�̧����"�溱���hR�	
^��n�ѵ��s�5�ʒ����,�~�ah���'�/�;�K����j�^��%�i7֚	9�as	5�ź��z���V�������������wJm����L�:mt��P���vvJ�Tjl�1�n��;��n�`�(��՜�I�U��z�R�z�H
�C�����R�y{��C�,���M��t��E/�%֯jvTV��߰�#W�9��T�G%b�����F�{�����rew��27s(fд�h�8���0�]E�_#�Ti���R�++&���a���
�]�#�䞼.�E�`g�����_c��溷[���Q�!tP��'I�v"y[<]c=��� gR���(�=Gl>[r�Wn���C|��l֪��%���E[g�"ܧ�(#2��
|���f��W�OC��w�=�W�d�V-�VpXwr���w FYT+%��H��!D�x���l�d~6�7��dT�
��ީ\E�_N���"�]RdD7�-obΥų"�JG4+�B�mm���v/��Nn�ʅ6>��K����Ɲ=�Z�^��'��ݎ.��o7���Y��Ox��z�������>������K���X�x����![LS�Py��ʸn��^o��})c]#���i���� S�W�4�O�g&��b���z%����*�\��I����~{K�a���՜�Ƀz�"=�OjU>���c���]��ѽ#΋�y�$���9x,�׋R���E�zw71������9Nn�c��v%�tr�o�Oo�W8���X�70�w�*��V{V�{̺��%�:rZ���aT����{,�B���r,{�v���gX�oo��)[=�~8Y~m����u>�]����@n��S�WH�S73+��Vu��$d��jg����	L�f�\�Rh��� xL嵅���~HH���o�����c6(e+U�Om�����u��P�����[�'"�{����P=G=Z(<$��O�;+��8.�K�4�:�U�y�j����՜J+�տGC4)�6�4-�����y�ӛ=�=����mokW�d�}�׋���%�wut�M���vٰ������J>A�'j�UnNm���K�q�D���[�o�$Ӂ�H�UA�NU]��+��0r�F����t����$�Q���v!�C�7����x
JӱX��u��u�d]�B��ԗ^!���eRŕ�m�^��6��
���a�=tl��H5���e����&�lf���R2��ٮy�lO�9yվ+y�Jp�/gG��K�k���q�J�s��?r���Zs��v�����Mq�� �o��o,|صݣ�I��u7�yC1U�UV*#'��-�ʙn���(��o�'MW3���;�W����t��#�KBpc,p�4A�4J]4�ښ�!��B3�g�7]r��y�[�k���ݪ�暰o�#;��H�e=G��Ԭ�<c����W5�J��PR����GE���n�u���s)�RJ�mk%�(@��!�D����fΌv+����u�Ŧ��[N���ιt�!�"Y�u����L��i��C)�OPֺ�9id��o�4}"��؝F���7�/je��8�:9 2z�_r/��Xku��.��#[�_EY{�S6䢴�j�|`X��>!BŧB��Grf����%"U4D�dOB�Z��:�"����	�K�Yv�,�{2�@w-Zk�j��sR��� #3II3~�9��Bf|#x�z)kT�=F��,�3l�-��;�l���J�C�1����f�vj˛tq6��3�Pn� h�[���^��g9E�ٙ��Z�S[>�@��у��nT�r���h���=
%�w�����2��૵Qq=�Y!q�[9ϓ�^�V�Ռ����K�"�b�f�:�O����&��c3-��P���n�6	2�/�D��ߍ)O�w3>����N��گW�;SIN��갇�0Q�T�0[��+
�wYiw$��{]V	�7�$��s��Q���Ļ�v+���,>�j��[����e�ܫ7��B�Gzq�d�l����X\�v(>�,�mݭ-4Z��H�Ŧ��j`)c��t�+�v\���adUxN��25HP�P��ZgTܵ�k4�y�S��l����Tth+��\��G�����\�\m�g�4TK]L��v�so]
�ͽ���QP�骚�l��HXȖ|�KSW;Pw�o�[�'v�J.����ZfM�Ј��9=ߚvҀ����;&���w�Y�g�w�,��I�v�G�ivM&���Ws�m�
����S�%LEm �<Մ,�gV��@c���	��_
4a��kLX�GY�����)�����c�wv'K~��	hv�j�k���4YDfH+�q�Tz�$��w`�U�k/�k�7Zݒ��@���]� Z�:�Ζ��j�|ça�'�^�jوe>�]2yC��m:��A��ҮK�%�Pp���*��(�c&��O���,CoiJt^p(�L&�im��R��T���Lԑڦowa1����/45���d��N�Lac��Z	L�U�P�9W7��چ�h!r�8٫�9��#b�D�hZ�X�(F�F2ZW�����JZ�ۀe\�E8�wsZV3H��B�- ��iɏuSvb�*+�Y@0�έ�+*�kbi& Ý��2��%��Wp�v�Cv��������&�P��C��F�*�AĢ[��֍�t�ұ�-vX���}��%�{ �fI��m�z�6J�]X���qN�@�T�f�0m�]�G*Uq��LX��{�iI,oU��L�a6ҹ"���^8�mtP�d�:��ob��� �6�>�V��mú7RFnAw�ݜ���aU�/z���A���sk���c0��IA-}�7H�x6�x$c���}3k�Z�)�p��7hm]�wH��u.t1������+�NQ�zΤ���8^����b�D��Z�軗M��ݒ�	��-�lơĪ�_b*�v�W.��e'�:J�x�_�)me
��-N�m��T\�E5��Mj*"�R�W�U3F"�V�&�
��h�*��V��bķb�
غ�,m[KE�R�٭�*�5Ψ��Eu��*Ԯ���UB�m\Sk��A+U��dN�UX��"%Uex��1f��MeB��5�d6l5�EKm�6qTG\˨�X����J�
�Ɣ ᩑK�F�VѰ��5*�8����T�0�Z���p�TV7�=��{�k��{��ᚘ|r�M%�-�uƢB��al�9�s�P3V��<�~���O���]���<t�[�+��¡��C{(�/-Չ9�;��|֮�bK�� Ց��-ιl�J����U9�!���f�]_*�"���"��X�<�--��x�!�y^��6�/D{ӣ�F���^�ߧ7ۚ��q��k��;\kΞإ�+��W;|��O�7"�6�ף�����'��Bҁn��=��i�Y⩊�R�$Ӏ��h�I��o�	��ws�:��S��!�P�1�8D>�ݩǬ�Z��:Q��޺Z!��p�\�1KM�>.��7׏E�Tr+0Z3j�{��)��YJ�Es�ʗo�\7�wp�<�j�;GJVs�`j��)�O9�xw@I v�q���kNdU�k���SY�VU�,�giݣ|e�6��Y���Nj������"0�}U_X¼��V��������̴�pײ���v�T��-��qb�#�q�GE9�e�{�3R�UF���̆�ӵ�ܚ���5u�<���g�ċ/�y�f�9ƕn����c܁b���u���8��w4v�JOh�����wkG�tv#�v��'S�,ؖ0#BZ�/�z�/,m��wH���Fg{���п:۔'Z�h#��5�b��
��^���L("�t)�6����$�M|�ɼ�u���/�;A,�b;�M	��Ou��8�(�����;���vq��-�P��2��6���;To-����l��H,~��K��e��� }Ƽ0�6k�ۦ�	t�I"5W��ؼؤ��nc���ִ�r�9j�`��)-�vM��%޳z@��R2o-kL��"�&s~�𙫄RO)DϹ�`k�T�}a'A8	)C��D����E>l��AH�dT!*#�t�Ǫ��	0�<v�jZY���E�0F�,���V5�͆�6��H[%t��:��5����h�*�tu�X�i�"��FC����ܦ�:��	�z��rɣ<���$�B�!�w�׼���lRά꾖q7�g��Fc#*�X��ذF5|�[ٹw<��$e:�۝*h�Q82�N9�2{�&��n[��T/�Z�f��vY�.�^�p�E��cP��smui�*��`����k.ڷn��({��k��2�U�ڹh^��o
��}�8�W�;��Iݡ��s�@���(�IbҶ��7j�
F��/�E5�jN��kگ:�sBw+���١���c�)�b��g\�[ZK���j`��T��ϲ�u��V���I,�$n@od��l��w˅��qIWf?s�^~^����,�]n�i�K����s�VUe-��PԺ�g�]#�Q̴ػt��k�\�=W���щ��1��&_X�[�J}���!��'�fcz���kTѷ��C�֧O7���R�����#mU{DcW��rj+��ƅw]�mI�f�E@�#GKހ�=T/[=�z���%p�~k��:R�\�W�`������������5����uҕs�B�u#��@-I�N��st��s�Ԫ�l�j��K��Qf�w�Q��=�]�vڗ�V�	Yrq��,�@7��������A]���w]3dR�\���Z���ORjs�̮Y���p��W3$ ���]P�Gɶ��Y��܏T��^Lx+e�l���l*W'Q�2���6�ڗ��
�Ne�ⶳq���6����,o5��	LnWU���jU)�y��9��C��Y�ۚl�7N��S�4� �T')�z�f�FAȮ�m����I�5��ֶ��Etu�۽Xr]o�:�~��^+���-E�H�RKH z+n4:݊kYlػr����dR�'rU�ш�ͫ�wv�[��ɞ->)u(�����C�ҳ1�©&��j��z�"+{�����;��`�|}�ܗ�V�sl��u�vW&u)��dw�}cG���^�=N_���7%פy�B!��]���f��Zɷ�I�����%t�f4��QkVR;�n�PA#]7[�Į���%�J}*�a˻�rl��'eXCZTU�e��*�3�*�&�7��:��!'I�CA#,)r���'FΩ�������Ϩ������0�AB���� �w.*w7�K�J�) �V��h��ǘ7q=�Y�F��j��N[AH�Ybo-)�[��m�!'զ�f��7���a�.l�Q�M]��5V5�7&wm�e��(�i��Fj��Ne��"�`�7r���ӫ>����#xUHإ\6��	�<˺�$\KOc~�Ϗ��Mk�<�)�A�_T53F�c�H&��E�=k��-���o4��ܛ�Cf��ޒ-iz�3p_2��Ml���Li��c�prd6Aɫ�|�㺻���z����*�9>:4�������\ww���U�mX�d�p�,�ս��m_18�%��ܔ^G�rFSP+ִ�]���o'(���v��J�]����BC��-'��7�v����Ryu��j�$����A	��f��Y�s�O�5����S�_ZW$/w��p\��g(=��Z���{iR�Z����0�6�JR|�bz���.otRr��F��#_Z����I�N��uM.����"�6�9�#�t���τ��s��{d+�F4%��R����SA%�Ҹ�V&:��m�,-'dj����[[m�^��U歪5�:N.���[a�b<5	�k�ΰ1��ώm�i`Y���~��pG���jv>I�w�̕S�d�ޝ�{R�uӴ)_x�k�ԠT4ݽ�T"��7I ;��s"͸N^���R[ޠ뒋�y�ZΜ�#�sU���Ǵ#���b�2��Qۺ�{հ-��D�ܘC>��פ�t���Z>N��8^o�e6���KF�δ����#yu[70����������5����1�)ݷ�4�����bq��>F��xz6�PS�UN;�۝��v�)�콃H��5�[�e�(��$n@oD�Z��V������]��VS=���WܫϚ��Z�#�ۈ��ʑ�u�hN:�o��Ko��{R����UƑ�b��S��x�c��0�	f�*W]$�������th�x��K��TC�|�'BWT��rܬe[��;0�;J����L����xvx�jvZ����G�_U�}�є���e����t	�u6��ֈR�v�e�|�b}D��[�a����6���;;ɦf�ٹ��j��J��T�9G߮���V�Q�4���w�w��^i���αק�L�y�
z��Ќ�pz��:J��huW�2�l2
��cD)F�3�̗�t��Κ��5���v��2����x��~�Y�{���k�5y���R�}�� GQ=�c�WY���mdx�tM��kD���)J�9+)nf�E�01�?B8{�/h�5!홞���#����R��ǭ"��3sᏖK��V
4%R���b�.�w�Ua?ek6]*�mN(�B�%P�����������J�cePKk���􎵼Q�J�n	+W[L�\˝<�	�
�#�OE����$|���?o����U{2ns�J�*�&¾ߢ�V2K��.Ꙕ��s����G�&#�o�N�i�r{Ƶ�6��l���rM�t�EQ��p�q�0��ÞS�˕�3}? ��sݭ�&}�0�ZO@+�6�nb�"�Ќ��d":���GvU%�������7����MI����o�	.���x9�+�:ӭ��H�z�v�-��=�!�fr,�.��oC)����֯��v+\7�4�(h.��+��x�Ţ���֐�X��f����N�ۍu��%א�ؑܢ�bW���l�[�ԏV�t�f�W,�R�>Fm�-Oz��6��۸��M���������/[p�[P�@w36�zݷ�s~S-�r��fcU���̣/�ά��&� F���4�i�{cWJ6�lu4B��Z�Ջ� �4ʃ���kr������S���/{��ƀ�5��:T��E�7&���O�5�����y�� jU����xC�D��SW��Q�t`0�a9z�e�����e�w�l�Yb��h UXX�pt˕�;6�%)��XI*y�1U�D]��������}9�9X-gr���v�\��n#"_Ç>��db��RpO��.F�9���e��^�j�=�ݺ�4M�)��v� t�m�fn��J�]Q0f,N����C3�朢�e�</��i�[i�c{���W(�L�5�B��֡�����YJ �s\���7���]O��˛ucwQ��[ 6���>��ḛ���]v.1Kw�]B:yx�m�U���1du���ĺ�ïc��w�6���+��k8�%'8qZ�m�Ǆ��G
9�ExZ]M,�>y\��x6�'�:�T��W,��Y1��j�\�K���AP�4+ש����Sm�b�Ў��S�Jv���5�`�WbԘnM�#y���7�9�Ή����C�w]���G��� �"��ڹ�rt�6��B7;�l�	�w�L��w�)AM�-mq�[���)CC7g'��U���n�,�� w�/4��b��pՎ�SlQ䵧�_�k/'s�/P�ޑzșA����������W���-�I�tqc��$���$�!GRV���W�v���3�K.Y�v��_��L�'�.�G�>\��/;kh��]��Jؤ�]Y( $Fd�l��v�.ӻ:�`5w:��a;P�)�K~{V�u�p������Ue�'��2iA�g!��f�Ɂ�K���պ�Wu�y�8"��Sގ���W7h�T�Ғ:]�{u�Ȕ�/��	���%�=�`���|Jn��oa����N��H�=�[��_X��$��Y�=���0>�����t���2q�D��bV�Y��4�Dm�\����E�`�}cI�@��\����m�틭��L4vMK\�ٚ�[��3Fl�QMi3�֙2��32��E����۶�j�J��b%�A��-Q��Dֺ�ݵJ�GTm��DW&mqih��ZQmsu���ₘ-��UUKF�F�Qj�Sf�cl��Ю�ڮ�Z�t�h���5�Ce�ҥMh��R�̆�W1��X4hb�@X�5������h�M3F�E3�����7�V�ڡmm.�4�Z�6�%�4Q(�YR���5msJ�FZ�)Z���"Q�����F�k���Ʒj��K�VTMK���"؛�8���kiZ�V���U�j�����U[�b�	��d�mu�\�Z��m-մ�ԩN50�ve�XҴ)���s}P����p#�f���s&�rtg0�#����:=�v-7��`��l��]�wR\�����#ݞ��g��]8��H/���H���e�*�3�"rZ���q@x��QFk+Ki��S~���в���k˳���W<��x��%󉡓�ח���O�	�@wR�%��#�/Z�+]
���!P�#^�C�o�f���w��sA��ȑ����R��3E��7m�N���쟷R�����}��J�;�-{�q��G�����3�䨧]�/O֭�Qά-ͥ'��k��d�Lߘ������]`���*h���On�s(�6����ᬎ�L�'@�j�Ӱz�G+lLv�Pst&v �K՝�^H�l̚�]��������:b�m�s��f���pCw]�-Լ>�i�l>�"�3RˑwmY�|��.5��=���Z�)�-l\��Eb�=��\H�gύ	�N5�C����{{�v�X���
�Cj%pU�d0�![�Me�VO�d�)K;��5��K�Ɏ�:�ܮy:�R;��gN���*��N���8��~�2�L�SuQ�q>E�ܧ"��J}�d��*H��o��Z<�{f��0��8��8�ۯZXF��u�j{���;��Mf�Y���Ge�Imm��"l��{I�wt�>k*l������@������{�bª`�|��ͪ�{���흴��h�#r�7RF1�M�������?N>�������>^�W�Eb�$��jyp"/�V�@����X��!K�����|��[�D@�����yv%/F|�ZϮ��H��d8ّ,�G���5�#�
�����������ؚ�lޗ�iCS3���I[�)��>f�����Km��K����J<J��Bt��4���`伎�I�}P�)%~o�-�T��������sT��'�u��J����-k��mQ�L�H�K��jmx��3Bv|���t5�����tx���%:I��`#GW��HU"Mm�a]�F�\d�ѳ�
g�C ����װ`CĹn�5j�5����륡��C�F�51�E!j7��֟ZcE������ʫ����)徝O6��K��|a��0f3���^ZoPܤ6�a��i4��o���ި�Y9�bq[Yo��^)�ib<l�������!
�ϼ��� ^�HRMil�����,M�Ku��V+q�Z�o	�FI]�C��6������x�ލ�\��@J��PSb�rJ��8���׼��<��q臕Z���dC2�6Y�g��U�SVi�ŇI8�]�jlb��++i�8�Y�e5s+����wV�j&Z''S��"����R<��ת��z�7,��K�Eu�˽>���c��,=��R��H|�ɬ�^�]wf���k��I�9�x�E���oȎ�M,�5=�g�<7�5��ɍ/�&g��o�K�&k8'n���n�a�m�Z^�s�sk��z<C�=�0�����-�.
+S#���\7�2�4��a`���S8"A�2i'�m-rΘf����:e�Ȏ�
Y0P���%D:>4Pg<&נ�����e�[�`9Z�T�����VR
Y��U�J�I��EΔ�&��'!���~n�M����s���Y��*vʳ��9�o�:W��m)`�xE�[��e�n=(���h�;R��7Բ��W���w5��4hwj�u��e%�C�U5ӥ�1шM�4�'G�����QE�nS�����M���\�̲��z���u]�Y[�Nf��[rѯ,�6t>��~[�=貆xB�Y����+9!������{�]5�\[M~4�(m��ɶ���3˻�����"��%�O?fĊ#BQ�����"�7��}\��w��ާn��.��p�4=t�0D��wQ������c.���t���d^�"ڕ��E'C{-{��=��X=� ']��'�	�6Nѱr��S�;|�`��Zݭ�s��tO;JbC�PRu��QۍJq��k	זb#²oU��-���#'&��J+�ߓ�x���}ھ��J�������Y%n�p�:�jR�ѓ�v��v�.�c�>S��y��>DT�&���YnM���3"�Z�}X�d���$j�'@�j��o��4-u��>h�0�1�4s�v4V5��&j�w��Z�@���b]H}٧�{�ЩC��WOx�=M`��xpS�#ڄ�Թ\�3��F�ؽW+��!���߱���)��6��H�]�f�晽Lps��o/)�5������h{�D�o?I۰~tM8A{�����%���+��*Y3�vV�^��b��V�usˑ.��h=՜�(-"-�x �bb׼F�/z�-}�%/<6�YA��[\����b��4,�7%:M5sxI��!I}0m����;G&�OnQ;�6�]*��ڲ�m��#m����Z�}[�4��u;�J���(.�ӎ�{�Q�VͧW}��y]��Mv��h��7(Hn���K���v�ի
fƙ�J�ܨ>h.u�t`��U��z���<١oІP��E.�}�'w�Թ��}�pZj#^����o�ضr
�pN�MJ뤕��G�:�E���δV^��F'�a5S�����Y&��ڜ�gj�<���������֤��=���|����wuZ��I�*� h�{�ni�I��y<�1e;�	�<�(V�sB�/���,�c��D��P�C��}�Ȝgd�[t��"}ivУ{]Q�Co�ۮ���JG����}����W��npB�C�R�+$�<VTCT��"S�J�׹�u$��e�k�I��9�����t�\��v���t��jr
}���o-*r��7�o�
�V8U>;���Ώ�k7������:�ʴ���65q��\u7��5�i�5��s.�[[����Z��M*��	��mQ�U| p]^�F��I�Զ�d�@-����%!o��n���e�u�NꝖ��wxwS�h;���:�֯��[K'']W� �P+˔�����k S����I1����9�ST��rb�C�V>t�Ј�C�#��'��S��'{��yw̾6Y�*ڲ!��vP�����ܖ�/
�s�d@�I\�얡� O���}GR~4��m�A��I<�{!h$v��,�'J��T��N/9^��V����B��Μ�}�0��#�2:�2`Hs͋�Ry\V_U�S�n�]�h��lRE��C}^��/�t����ќ���j��q%z�v�nl/]�r5�4��E'=+�v�Z�����\7�4��p]K�y�L��C�aLN�6��]���Wf�b�g��{�9�ex�����8�V5c]+%��W���x��m�i
1T�s���ɼ�jm�᪶۸�m$���bC�v�c�O��#N5uyQ�����ݭ���*�k��+���%+3�6+�6�he��$��vr��hj�H��*F�3ԍ�|hm��)��2�A��ʴ����#w���s�ZąaC��Vv5K����^č>�M9H8�qZ�����#e�}u�aR�kJg&:W�Χ0��O�v[�c��
%c�����V��x�GY'j�).��"ow�.��/\0���Mʨ��'���\G���I���KnL���#BU:���᧡���yO�-V�R�nΖlA]]����rx>�{2�a�N=���k%о�x�>h'+�c�؂7d��(�(�SWX~g����������Y*ⶔ\�6��͛�=Ba(s�����X}�u-�=�݊1��ڒʈw�} ���@|�X��!�����ܾ�\K��L��		pHv���Oƕ����I{tS[U<RcJ�D��|rC��tj��o!��vcuP�ʰc�4 �Cj'{GZ��|a��S~5n�^ ���Q��b���\ty��l���ƕ�SK�@��uv�$x�#�ZQ�z�+�r�gN@�5V�	kݠj�������S��)�\�J�Xh�Y��]a,MU��:u�'(��=3��K�7{&�;A�`��3o��kl$F[ћ0�vF� O�GqF,j�Z7%ޮ��ݙ&�#F�W��@o[�x�����_^�/-�`��c>u�5/,뫦j|���*T�'9�h�v�i�+Eve4r�� �w�)C'm���0���ɢ�Y��^��}����JR�H�X���8 �d�5���rvi�N喓T�} �Y�s�����B���:2���]���	f�9�V*�6�-]Jn6Ef.al�r��l��WtpQ炸¯��Q�О���5D�Wخ���Uwe[��˙�@�#o)��C&��7��"�.9eq������ur@w9��L��7��1F�t�����H�[�s+d�3+��ݪ�z�L� u�qD���)���VDi��ݺ�.��C��&�\c-d|Mf��]IK2�9f*�-Ո1Kg7;�X��.�3��V-�mi+�yאr<��r�wZ���J:�(c��N���8�,- Tb`QҮ�[�Y˟Jb�3�[�S�&uI�3W,�-�Vyj]�EX�f^�Zp.�5���;J�g� y���1�)[�g^L̬y�7���f�$�"�1�r��.���u�6����9�>5�E0Q��Mj�(�$�J^�k��N�^�t�(3Uv��^N��G5���!pCx��K+��(�,9���6�j��s��n��F�ɜ��;q��Z{�9��Xc�(b�\o��:b����
n��8he�]lE�4*� ��ܱzO>��[ۻ1���\B�Ʈ�uAi�ӪA�~� u�J�f�
�:a�w��h��zr}��N�G:��T���q"��Ƿ���<�ou-ܚ5�لѣ��Yk�'��˄��ws�Sѯ���_&���k���"�q|�A���� ���.�H*@
�H�4�% �v�V�ڷYj]��ZT�[r]��m�\����a(ն֭[�p�����6]��Ue�A�R�l�˚,�V�VV��diV5��m�խl��^.fÓ0�VԶ�%EMvQm#uƱj,h�ʚ�#Rԭ�.��m�+e�+A�ʺ��8Dk)k�dQEp�Z�R�+lf��FjR�lR�Œ����-V�3�S[Kn��֋1��)[��E���*�im�j�Sk�	sxn�*���W:�6*�(�����75Eֶ�&�2gR�,�5�V�j���΍����cl��܍F�[((k8Ӎƫ��.�Z�����v0-�b�sQE�WV�Vf�kk�mD�R��A
C�B��;�r�Fk�x�ۺ� 3M�<����'	���i�4�tPf�֞�L�����ʬ��nk�@�?5�|� j;R�s�_�/EK��L�/d]�4�Y;���ҫN�$����ot��i4^ц3i.�ʪWr��2U�ن���RG�.B�̦�٘6mա�D�ՙ����y��F�)��5�A�*Dak+d[��],���oW�"�<wH�1�k6Y���CC}a3��T�X�����_J�D�x�J��םl�+pJs����h�>iw.|��:P�'*0��oC��y���/����b��Ox���!�r{�3��ER���������.�p�Z�����D���C:>2V�uI���l�QJ�βTLLYo��SA3Օ�jnk��ڊ�\��m$���̷�mE�_#��e�ohu�rĬΰ��JP�\7��ײ�����'	�${oވ�`Mئdt��	]S2#yH���\����[x趲ԛ}i[���!��w4FLԣ�W$�4np�^��k�-�I�*����Lv��J��j3�B�+ѵCn�x3pP���5^���񧷐���7=�Mm,r��<#P�(6.�e����{�.4���U�nUh�n�zʮ�-V�Z�ya(v���r�/f3���]&�dK���
qaEL�(0�7�L���85@��+���`�xV��B��^��#�D�©T�]�'������77�bF���M��M��2�*�{��^z����򀡔�ƾ�ჅNo41w�mm�4lh��x�{ؘ�)�Ȇ�u�w�nɧ����y)!�ٷs:�m����fQ�K�*ȳ��Qj��N<����.�჎���kɖ���Xڌ]��B:a��9ž��E��E�P�$V��e��HΣ8�	�\)��I2�|�1�'`��^��CR��f�X��%e���5q1�ݶqd\��d2:���H���|U�ٕ�.��V'rL���k}Q��^���TS�@u=�Z��s�anl/@&�BX�iff���q�x����_]ֺ��֓�f�睤���c�1�f&�7a�z��y�γ�V_h�(��<�z�)�k�t��2q6訜TK%e�)f��Z�k��=+"���.=��i�3�����PD��q=�����m(��C[ڽ�h��-E7�T֧Q�ܷϳ;�^�G�@�S3�p���iSH��Ԗ����QOqY�,�� ��'�+�UQq�v)c���������^���v�=OF�*N��#:���{�o6{ޗSlKw�Nn�XŴ7�I��-�h��ރ�������cl.�*��U[u�#().�͚4�����Oϵ��U�ˡb1�+nw�_$g*\J��f��;��K���Ÿ�5٭�|;�5���|���9�JP�#�#�s��:��*���!go[�ܞ��x�w_R�1*��s:��!��g��TT3��MĲ����Y5�U���}�}�5}��J�U�ڭ�l����e"GN��f�o����Q�V�-��u�N/;��1NG�WR[Y�y]J�E��|�VT���7�]D�����_e�d3�c�i�c�KE�h�Z�f�\^Bb,��W�E71�
&�&��voG'��=���v��\�x��Gh���,����\�y8�!��f�!�׎��_Zo�Qa:��	��eD�/�HxR�{}c.�
)��{^�;�3����]�J��}��5�������Z0Ƭpr�+�+�0{�/&K}k0�w��[n�^9�"�1�R�y6�������\�c2��e���i��GVWL"��^.S�������8����F\��q��p`�v��C|�܆���n�z�
R�V�ъ�p�ۭi��i�	��-F��d��Q!!�W/e��&��V��Q�n��Ve_B�)�q��V���tGbۼg7.�%Xv��n�mSǐ������o�=%��Os/���g��Kq�U��yGe��m��>4{TwKoJۖ���j���{�<�ϻ��t94l�`�h�mQ�[����b��F��[@�t�Ҿ�O���'�Z��J�T�tHC�B^�%�5�`~Z������ej�^�{W!�B�l�7���k��ȳ;<.��X�͂`�>��J����m�bN&QTS�n��OA��S��	�$2{�th�۫�Z����),��wZ�Ki1��B����%��(
ʚ���vH�(>uY�Z���]A���s��Սt�C�p{F�8�yŊ���"5��E��9�s���&+)�	�|�wh���2����T)]ւ{j�|/-VϊnZF:���N9'9�=ޘ�}fm��T]��/R�a\��|��+9�8jP sI`��@7�d��Z�t���;���]zU��N��f:"���D��BlJ�s�t��}MУ�YT������zX�^�NwYU����G���O�g'�Z�N���ma�U�8.��"�m�OlM�ToԗV���޻�M�o`�E0�ʹ�<�ܘ���OT�q�3�ǷȾ4y\3��Z�g4����<k�衜�'8��e�r�P!Z:	�z�ˬ�
��L>��H�}_��O��SOt�s勚�΅Go�%�\\��e�Йꭦ�;���+G�ԧ2�Z}�V'sdԛ���+D��u��J�:����ֲ��������#�-�I�!ٗ��5k�g��.�o_�wL�L�.�����59Z���l}�x-&l"�e��K�2�)���uv���I��n��3�d`T�;Vd�`2>#17$�~��!m1��u���l񫆤om&�}X�̀�hR�Ȁ���݄6��q3��1���F�T�|�}� s�~���McF�k�S�+�r{umP�ϼ�<�:��L#6�ͻ<��=����R�\�y#P�v�|����橄�������W���Y��P�T�2o�^/�h�a//?M^Uv[��n���km��"!����E0�4�}wJ�a�6p
V
ʫn����9rnf:^ii�x˼��ц'��"�17*�4a
��[�95ո�u�#�g��P���|_��1:I��C��^� X�N�_|j
�㕫y�	�=����4�nu��ܺ����S�L4.ʋ���Ҳ�%r�!а[�	�m.g6�@2�ҽ��`�b��|�S�ϼo�vΤA][�Hܱ/v�����3;��+�z<m
(͍yI�s�e���]���H�e	��F��nSߟv��_�}����"�L�
*�ro*�^s�]�V�HجJ���ӝQ��p��^�����#�2v�B�m��3��]Rg�I/os���=�:N\�����UEN�oYH���C���;0�	0T8|q�о�b=O�M<�'{_�:�	���5���>�G�c�E��5���7�q���t�K�;���d���{�6~�qf�&W��Ux�h��]������t��:7^4-;F��F�U���3�͚���u����{y��w��ِ�vtq�7�n��@��\R>R�sMJ�D8�dɱ�|P^0q�;����;��c�����[����ѕ�[=灂����F}[����0e����M��9;�ɤ��d�	��}���V��4v�k�T�"����[���X�I�ޣǩU���b��=}!���'e	��yv�v�k������Q�r_jg��.O�;k�	�<&�E��:w+�Mt2H��;)u���lA�V��6f^��P�$������{s|�Y�4L�
���s��_)�ݞF�Ofh�-��1M�\mYu,�&�>�mB�ǛY���yɹї�������&�XJܯ`&xt�a�L+Uԓ^�d�kY��b���m��]0�}L��������Eڥ�%�ں@�=[�p�U-�uS�N.�(.�QǸ�mϓͮ"������:�ڡzV��_�g_DƣEp��)��V+�d��o���*�I�*ee?�6���G� n�lM�6&����v�<[��������4�AXK�y��tu��oE�Vl�nTn�<�0E��ց�ֶhJ�4&�ޱQY��n�8���b���9��(�qwZ�no+�0U�ZP��P��$U�oU^�������9u4��Ns�έ��C���mɰs�S6�Ηfa��雺�K�;Q���a��	ArW]O*)D*Ô%ٮ����7�s�7X��5-�t0O���֒�U%>iW��$��L���+�;X��S��&���p��ss��pT)���t��6~�t��6��[�r�[�ܸC�x�Ov�K01=�B8Jo��$8�P��X�A6$qގ�c����g+,�f-��z��3`
�՚�.6�d�TtJ![���|���58���v��e��pI(lB�6C-����XzvZZ�:�QJy����E�ʕ�:W\�iW0uK����vԚWZ�;����J�1�لQ8�:J�WC�0�,w�K�)�B��z���[&m<9��C�*���M]�&L�݆E�oX�%J��+�m��F�p�˺r�VP�����]�{eO�s��r��bom���MHfH5ժ������/u�:�����=�|�G\5�r�x
��tX�G��;�@{��vRad�I�&�ѭ��t
��r��g0�$��Þ틔���,�vuL�]K/Q�Zl�s0�T��wJ�ƹ뗍�*��R�g�.S��E��Ρ![��,f�9�gf˘��!+����5\�s��{ڊ'�Dv�kxIJ՗%6��YH�IoL]d�Ϝ����Y�._kX�bo|�S�:�>���Ӹ�HE��Q ��:�X�k(u�����7+;*1��o:�KX��a��P�B��֩���Զ��+ibᚹ3�p�U[J�j��q�Uڂk\֥Qjے�*�q��E�vюWV���굌\�8��R�W�Tm����L��UZ�m�-�qb��l���m�ѫ���Zqp��E�2kX�J�b����rX�v�R�1A(�l�Q��c�3l\��wW��6"��V+m֢�Q��"�[m.e��R�UJ6եkU���L�9���+�A�c[�X!J�[�p�����[DDE�[��H��KR��X"��rZjMm�!����q���;.u����e�B#�1b
�֪*#ix�b����̠�Ym*g8Db!iEe����֢�"��`��EUR�ɢ��ZܭE�EEMKQ�|�������{��n+�����J�Y%]K��B�n_����w\�j�2��[�%n�Q�.���#��wZ��L&��L�����C�F�t�"��Cj�6��f�)�N�,-��A�D��@Р��#���[����xT$r�v�V�a�uk]��Gl��o-��Vdz�3q]3�Y/*��'�F����(�ʨ���ͼ{5Z�������^�9LVƕ4I��7������a�c�MVIr����hi�u[h����|{7�-ͧ����FŔ��"o_�a��Gq^�
*��ꔽq,2!\�7'E��ź�y>���s�˔����ߙqZ5��7N�,�/2�h��7�;X�^B�0:A::�X���u��X���F�wi+��Vi�����)rv�(2k��]�:����Hҋ���w[�;'+&�2��E����Z��[nC�D�s�L-�D�;k������Tr��v�m5�Y.��c*�8�A��6C#����o6r�k#��x��W��Ծ���5��j�'s`��pK���Wבm��F��Vԥx꧶)kU��uxanP��T�}<�+wk�y^w�} ��rI��<n��θ�¥��rY|��4�43D,�oP�U�:`��M��V�q�?[�s���*�9]M��
*��l�#�����s�z$�09�B
�S��~�YJ!l!1''��Ҧ�NcN�	#P�'t��e�����k����$�s{��V��7(�G�6�=xN�7<��
�zG]��&��S��V�gE��e{CkY��ѐ�LR:�,���JR�s#�z��]bѽjк�[tq7b�
fA�(�O(��~��>47q�ٓw۪�ԋ5�!�/�J;s|�k'�'i��6pBU)��mв2�$a$s������=^!v�;�c�"�&�T`W�S���d�V;;�w_[�=;�bhd�P�b������YoYk�M>��ǒ��s��/�#w^;$�zSy�Or�,"�wRk#��ZI�A9Y�$_K��tV��z��8:ˎf�%YO~}�}��(L��wA��<�}���VK�ք��N��h�gs�5�Mw2�7���<�JS�|�7'hL�.ޫ���i�ug��E�|���%|ԮF�үn�&Q�T�:�Ǜ��+��&�ނ|�J�;4ɔ�a��>D���Բ^.e81)6S��l�D��*�N����_t�ۙcn��3�����7�=µ�0� 0���|���� �kT�=P�y&
��Q<̧�S�Z��l��~4�X�J�*���`��6a�ά}�J�7_so�,STM�HԦ���6�>P=P�!�Y��{yɎ95����Ց��ʭ�H޹����غ-c%���Q�؇�����f]R���)%�n��y�)��0�O)�p�L`��8���F�WL�w]}�ԫ`��č�]r��Q����	�v�Թ�v�y��Y&�X�'�U���TJ��/*p*3��l�Z��q��a4�׻gm.�)�|�w����G�����b�Y�穂�S�n�K�~�Ҫz֓�sN�t�Ҏ0O��Hw����H�l�/�;�e�YRXS�o��������@�-����3m�$��{V�ܾO-+��ԳJ�R1yhwj�f���Yi�ʹt�lΊ}@_tn*2[E3qgͶo��Cs�O��pM�,Z��u�|��_���p8�bw6	�O�[UJ�Pؓ9х�y)�ȎޖecTٷ֕�^��o��3�Y���g1Ad�[�c[���Զ��%da)�����c��H�7hmV�����~�[/M`�M��To
�t��h�,�����V5Ҏ֧�Q%�Y`�/�#V���:F�w7��_���Z�5髰��ԝ:=���R�FLf2�A.�:Tu'��[����d���!���]{���0���-�����k��z2�t9��� 8LI�c"�VF��]ռk�N�e���N�;�-<^�_U�x�X�3Us@�=)Z�,�oQB޾�ڷ�/�st�H��r�؜w�-g#���-����<DwFߖר������Fĺ�_��R!E��vo4�������$��J��o(���-����Kd�$�yR�kqwR�e�V>5�W�D��k ��i�N�9�'�zz�����WΗ���E��-�t{����θ��刦��.���lU5Y���f��7�B��\r���]RV�kZ1;�&���/�Sg�/�߲Q�`�q�On��Z��5m�wqk_�3T�2;�.��f�.�Ǵ���M�i9e_5A8V�F�,�&����:�SB�;���L���y��Et�P6���Ʒ���Z��h
���)��+`�yS�YX��u�Z��uڑM�;��(���in��nH�w]��}��F���!�x�7�����**�չ\�i;T`�u��:�Z��������GD&O��
�S��=qs�JN-&�V��6k��j�����$��'�+�T�c&�s\y�ש����}�����|�����qS���/[lݔ�L	êz�ƫ=�4���]C����r�/-����iu�'@nWU�D�#0�g�e[tE���&��S�l�v��6cA�1���#f�e_6]�nm�������P�W:�,���b�N ��k}sip�8�:Ƅ)�\��kM�lJ��irKrz��+Ĩ>k!]◕h��zĚ�z�����\�Sp�w1C���<㑓��qs����W�ҏ�ĳ5�~��h��������	����pٍv���̵r=�q���e%��ޭ�c7�q�}}bV���K�3�����>���6>�����vs%��J����^.�V�rұ1YM��]��.�xS��.��Г�&kV�jv��]f��w^���ܛ}i4�%ÂC���񫸙Z�f�Kx�Haz���-�ƕ�s�ظ��S�����\� �O����`m���+Ӑ�w&I��ͼ�M&�������{V89>���}O�,���H�o����I��u��y��t��7����syȷ��4#:%q6:bF��f3����!=ν�O�]���{�B���,����^d�����[�Og�q;���Po5E:�Xt]e�7PYd^�t�9W �vw�m�K�0d���y0�ٸ	��.��� K�>)��JБ�h��lR�E�Л�Aܛ��i���ǩI�z���D�4�ev���׆�40��C���[{bF�����8Yt�0:��*8���|�^����_��:
�nr5��?#��9�ۡ�onsMgb~�U6F�Hn��&���,ޜ�]FI�i&��9��G���Z�8!�$3t�9Ě:�6��Ss��[C	m���V#xsCD&Vŋ��MZ'�
���U�N�ɉ&A�)��iRʝ�i'�I�聯��kFٷ�S���}}��-vE@�����#��v+]-��/q��n����3 K�Jހ��V7���ۀ��f�.�D��J.-��'F�<����[�:^�|�S1r�NgF�}]��.����N��yV�O:�gƍr�G@r;w��Ā����̐��/tpΉؗI�_���K-K�V�X9��{j3�H���)���ګA65�t��N���TVP��;5�>o�,�����t��%,R��ڸ��z2&)�O�U��7�3,����{c�T�gz��P5�j�f�|�W�E�^�}�-�|�Ӌ7�Gv�v�Z�*x��e>��X�x)T�WY"�����8�r�I�=�t�{&ob.�M�BY�f�l�P�y�+6�����y �r(�-�C$pn��Zt��/����nsŝ+�|���p܇�5�^�k6B���e\Nxߒ8�.����������S��Z�����!��O�@���$�R B6>�DX=���	����L�ǿ�BJT�a��JG�3
�!Q��X{������J�@i<��E��� @�z��-G��]���KH�}d>�K"��sAHJW�pb�jm����"��(���EU�r��$��-{}Y�Ϲ|,���O !��ư�&?�>�w��!�ì?�
��JH>Z�~Ҏ��T9��;<R B1����?N��j�o�@��`,Je�	U(�_�v� �Ԑo�l�����~���
�� _ߠ� B#��9�4|*yJ��R B=.BP��R"!$u���KԸx���Ccΐ��XV��oq\��^�)G�("���d���ʉ/����x}h���!X7v�&	#�B�Q���$n�ؗ����R_�7���,%����w.k�4�#���V�w%з�w��8�	!������P�_��N�C�?���DD�$�D�v�D���ھPuE}�.���� S'�{��ɂ�b�=��̄�C��U��P�/�;'���� B!BUiT� GZ�T
`ɑAZ�p5�Y ͔%)Z��)!��r�i�����*���CÙ��@h搁O�w�~� ����p/���G۷-�|L�H����)�����j9�HS��A�o2�z��}GOǫq�}�"�!΅8pHQBO�t��Ľe��$�~����X�o;��V�h
��H>��BQ�c���<Pwx_h��`<�/�vYc!Į�v�� @�s9�؎<�"'s�HF �t�ߐ�#ݨ��N��|�
$�z�P��H� B?e^���'�� �#���_f� B;�;E��X)������Z�`i`�V��{�E�� K҈?�gI�X���H�
�,`