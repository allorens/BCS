BZh91AY&SY�Za5�_߀`qg���#� ����bP/�              ����-�Y"�T)c	�"�J���5� Th3V�RRRJE(�UkR�J��ͥUAJR�[
(�
�A����ԁB��@TT�%Qu��dQ -b�
m�h1KT+TQ*�U%@�P�i*kD�m�C������R�+[p �˭FmIn ��&�
p�*C�p �8��M�`C[m)ESX@(���IIRQ�����p:�[4
� Ǣ�  4*��]���T]s��r��ۗ�t�]N2�z�h��r�6}���=�՜wE�M����J���� ��e�6κv Wv�@\�64�	�}Q@ ��J��M�juT%@��ؽ���OF���Ω�4 �˶r�R�J]�}��U��g�Ǧ�Cf-��J�J�{���_mU��Ͼ�*JSώ��f�������4�^$�� ��<��5JQT��<� :U����()U�K�z��J�S�N��4R�R��y�Ԫ��(��9꺬����耪�'<�OPR�){����ޥEN��ޡTQ)K�m����D���I( �ܾ�UR�o<��P�(�����W��H[���P
�׷�� �tkýޯY�E�ͽ�C��R���y�+�W�y�E]�$��I��A굠{�$�]�����
�>>���绞�
W��t�^�� g��U^�Px=��R
�=�{�(P�k�z�B�==�zW������ v�)������**���w��%*�^�)-�M���Vڀ�ϩJ@��|)%:м���⪥=ɕ�T�C���T;gZ��o{OI�J(�M����w;o��ѽ�p� s� ,��  s���#m��)5�%���)H o���V� P;�pN��t��Cw��` �w �� v��� ;�UmD���y�)H �| ��4�� Fu`��`: ]Wn  �` n� M]� �VW@ܪJ�JSh�c(*�<�T� 3��| tō gN�>���+�� + ���F�{�� :���p 軩��������Ţ���	|�)I ��>�� �: u]� �M���:ޖ  �� i}������0 j�p ϐ(E 

$"  @  ��2R�(i�B1 �0L&�40E?C	)TP       ��d�� `�LOM%)P��a0@`A�&h	2��*T  &   р�L�o�(�hh�h�556�j=M=G�zOz'�?O���߬7����l�f�J����{#�wO�,[]�ϖv��C:���|z럀 ���*�
�@S�@!W��~��?����4�_��=T�e@V��$�O?#D@_��'�D�BdN�*"���?��~�&0���b�X�u��Mb�X�:��.�u��bkX��05��bkX����5��`�Y:���5��MbkX���u��H�`kX���&�5��MbkX:�XF:��&�5��bkX:��&�5���`kX���&�5��M`�X:�ČMbkX���u��bkXc`�]bkX���5��##bkX:��.�bkX����u��MbkX���&���8���u��]`kX���5��5�:��&�u��M`�X����X���.�u��bkX��X��bkX����5��`�X����5��bkX:����`����&�5��M`�X:�1��5��MbkX����u�05��&�u��]`�X���15��X��5�kX:�5��`�X:���u��a��u��5��.�5��M`����Lb��&�u��X���X:���5��]f05��.�u��Mb�X����5��X���&�u��Md`�X�5��bkX����1׃�&�5��`� �&�u�k:�5��`�X:��&�u��]f�#X���&�u��`�Y��&�u��bkX���.�5���X:��.�u��b�X:�5��Mb�`�X��c�bcX����u��X����5��MbkX����5�f�u��b�X:��&�u��f�8���5��`�bkX���&��1��5��bkX�X��X���N1��5��5��bkX�0��1��u��M`kX��X���&��5��&�5��M`�X�u�k:���5��M`�X�15��]bkX����u���`�X���&�u��X��5��`�X��ы�M`�X����5���`�X���.�b�5����q��X�`���.0u�kX��`�׀k �	�SX�u�c``� ��X����q��8��.�u�kX���5�k�u��X���.�u���]`� ��u�k]x���`�5��]b�X�b� ��]`��'k�	�CX���.��$`�X:�5��b� �k15��La��]bk15��`� �.�u���b�X����b�ы�`��.�u��Lc��b�5�kX�ǌb��u�k ��g��5�cX�u��c���`��.�u�kX�u�cX�����$b�X����X�1��C�X��5���]d`�5�k��]b�1��0b:�b�G� � �� �(:�@�":�SX#�kX�X � �*:�WX���]`+�Du���Qu�.�� :�WX��CX��u��":�X��]`�@u���
��X<`��Qu�.1�
�5���A�*��SX"k M`�:�SX�k b�Du�&�Q�(� 5���� :�X�kMb��u���T� :�X"kMb)�U5���� �5���kM`��5�&�� ��SX�kM`��Q5�&�D�*��b��`	� u�&�P�(��SX�kMb��u���`�
�X�k `	�Q5�&��(�X�k]`��0�*:�X�kb+�U5��T� ��X��Md`kX:���5��M`�X:�bk�M`�X���	�`���kX:��&�u��bkXq��u��b�X���&�u���b�X����bkX:��5��]`���X:�5�k �5�k �!�]b� �!�b�X<b�X����`� ��#X�b�X���.�u�k�`� �.�u��CX����]`��X�u��CX�u�kX&�`��5��8���q��]b�X����u��]`q��5��`�X:���5��`�kX:���u��bkX���&�#bkX:���5��b�X:��.�x���k���9���Q���w����;��G3����]��a��
�`�V�Liޚ�UO��X��Qѻ
�&c��E��V9Tr��A,�w��R"��Q��(�����M�ׯ�&B��4D��C���Y����E�uqeUnY�
VA�kc0��kX�a��=͡���7E�P1Ǖ�������&����z�S@��d�7TQ��ft̵Cqi�̗�Sl�M�1i�k.�(���KLǒ�7�����-'�U+RA��F��\�۠��O/8��o7�"Pͪ6Y�G(o�ڵ�|�t���woTЛʲ(a��F���u%���
'^���t��շ�D7*��ʧ�j��k�s[�����Ԕ�+�\�ڗ�b�0�4�ª�e���lИq�,R�G�1�]+�<MU�tj�=t	�F�ɸi�c$��D8�*��v&m�B���Q�ukd[�(��]�j)z�V�c ��Yti%��-��UřNħL��om@���ۑA����.���&��0pnk7O䫗1���c^I*�[V(J�n�{oMpG#�:���tA��Р�7���+� ���m���
.�f�xBGZ�Ud�]r�,K��J��JS
�c(+�ٕg	�K]��I:h�cAu$��2�V�����Z��P�B��Q]L�9c]޵Q�ً*�m����x�Yj�\osA�c]c�A&dcF�Q!�vکc�����`�[/$̭,}/Q���Et��Ӫ�ɮa�M0��T����5��Z]Af��HeX��-���0�ugۭ�0�%��.TޑU�nd�	�)�,�
4o4��1T��+)�7hXa+�͍ۣqDj]�Py2*�^�Y�L��z�oz!�6�RYiTr,6�t*�Y��.f�k�n���d�8^�ޖ�%����:j��R`҈���Ln��#i'`Л���^+I�䘷r^*Lb�-'�]a5r�e�j�Sw.D��f�<4I�&�Sͽ��F�Dͬ�KVè����Qc8Un�Wb�̭mScW
lR�=Ӹ�<Ŗ��u
Y�\Uviݼʖ�;jh�a�e*�5'W%eb�ݶŐCc��u��K����UǑn˶7���r'3I%F��
�=�̗Zá4n;�w��h��n�H�J�V�Ѓ���t�܄T��+oiLx%Kx�U33we���ލ�[F�8t����d`U>�T��P�a5�����ᥡ��m+�<7�������Z�*}Xʶ����kCheݥ.�E#GNC�W�$��YiM���$[�jd�lx�W1���mP��K�L�+-A���n��OfJǢ*v���:F�e�����hS���naذ�r�S u��Ը���U9�L�\����R��[�a��NP�)V�ֈ�eLK�k�ia����Y��b�J]�^%P��yl^)Z�ڷLdʖ�6&�ca7�4A�PN�6x,��n�^W40�V仑�gΊn���؇V"�N�KT�6�v��q��l��&���,Ze3�sVd �r�GB�݇��!��=��P4��E�ȸ����~�L��YrG�Taeb�O!"[@�-�����v��ê���Ls.�%#V,�����̬�d;T衙�풫hz��B7�%�+���Z�Ul��i`�`��ɾ��*[��&��͏6�蹈�z�FQM�"��Cp�AV�@��2k��5�e*���$���t�L%[7��rA*ö�֥+�a�:��!vQ�@�ɀu�P�1�
�(=��BDwb�dڱ	Eٻ�F�qXCNv�*��J�X��2˭��˼UR!�.�±R6����Q�L)Ź�쭳�,�.�U�L�9oqmL�Ľ�2�m��h��+�h��h77�QP�L�mJm���]�\�5�YXw��r�S�#�5�w=B鄕����[��Nc
Pڌ��Q��OQV/�+͹yO@�2�:�'-9x�bzb��YWrY�S�mY0�/%�ذ
5�*��{n�;��������5䡙aD���������#߅��kZ �[���F���N'sw@�2R���1곆�]1!ӛ�qi�T��v�����ɮ�e,���P��ʪ�E`B��x��PmG��޻Vou�him@e��1����i��U#rsO�k"���[;�����DY�Y�ƭQ"ݸ.�\�KDt�����r�G;��`�)f��X�vZ�Bn�^�b�P�,��u����*+���k#��U̥v /f,J��K2lqR�
��KËtFF]��ľ�A.�闭e�ج�F����ͭ�`Bt;d�������{���)]�虷V�
��m�յ�e*(�L%F4�D����pY@�˚�&E=x�m;�7�]��ʼ4�:���9z-�R��r�-W�iz�i%�;����ݓyV�T��-�^G�a[��z�f��!�5��Y��Ԫ�t^Jמ���i�#��&��.�\27y$�bT��0L,�T"Z���V��{����t�OfA1�z"��BV�,��x��ͼY�Z�$'���r�onf��q��d��74�z�ő��H�y
O4ۭӯ[B�v�����v��1Sz���A�J��D��j�q&��Qi=��V�Ҏfk	`��%=͗76l��X�ё���tMz�t��[�ppU�ܫm��r��*a���Ƿ��;a2��M����n
5��yL�-|[��^QøS�9�w�oZxC�eґ�Wo��#C)�2hv�`�̼�f;�+,�kx�Â���5f 3%�bˬ�f��b�3t��wA�d�yX���7v)]�hE�^��[�T����F����Qăx�;^��pS]�G�
(qE6k�7��
�`�׋��W#HVJRK��0nT*��r�N�,�������/-*��V�"��ie��^kӳ<�WI�E�(*�L^���۬x���{uC���"<h��d�.�@�d����k���Lx̙-�A^�C5��F$��Ղ�kHm���U�`���H�ic%�Ch�WUl�(�vP(*�ʸ$�r�c���֜��˺pV��y��|�H�\�p�L�-<�/UMO`F�r��p1u��k�.P������x��9`�x��[ʻ�QMiCA����k��Q�qe�k:�Tl��2�
��I5SgƷ]�0а�om��9A���V��gр�x�M�ҐӇ�hZ�޲��c�����|�OUǹ0=������On94��~d�Cd.�k~Z�f1E�"c���n�7�+4P� ��س1ӑ�4Z�`�fD%�1�Z.�fvѡlU�`�V�h֬~�m꺆)�+*2���t�۽{w��OVh�{ԯ\*�s	 FP˲q�	���76jZ��64[ո�7l4�f�S�Ck[�R��FBż�8P��5݁x%ÔF�F;����Z�3��Zp����xd��MIf��˥Y�Fb�m6YK�LAUX���Sa�`��Y��v�-�('c#uz�VX	;N����7J��(�W��m5S<�'0L e����W��c�\`}.�τ�v�w�f�����K.�]إ���Z��Ыǅ%���1b�X//
�a!US��Z�2�U��cKwV5)�.HU���3*(��Cp����թF��sCKw���cslЦI��SW�f���U�f=n֎�w/�qԎ�V㤇��GZI=���n$.+4�smy.�շ�l2�	}5�d���iն]���kK��@�m�ڤQkS��Ek^�fԽ&tn؁��j`�&6���U��i��ڇua�Ubiۍ�M��:��&D*�&����;��\��������`�UV^�RѴ'f�t��Fv��3( �$l�/��2�kxm�C(�Fb{L�q��SpXB�(n[e��R{���O^�˺,!/	���V�W͢�Z��6�$���Oݵh�0�2r"����FQ���20f	�)ֺ-���mb�n��b����Z^ZwE%�F�L��,�\��n���̚��7 GbT�	TiQ�)�ƝG���,��»��#h�6J�K��Y���0���X[2nVҼR-�1Ұ1.�ng�n�#j<\A{S{BH�RF���TR�%e�l%�s�yA^R���+��s#�W����Ҫ1�E�b��[$�8��V�]����ׯmU){Z�-=�7�b�Ĕf��yk2��܎B�Z�5/e�[y��U2��BזE�3n�@�N�Y��p�7L��M	��(\��-D����nk��(Ӱ��j�Hʑ�;M�6Ե��!t�ʨ�GC64�Z��ؗ+��ʓHWa��2�k"�ՓR��h���`�!�.�OSM�$��t��Mܹ���=162��Ơ;%�l�ĆQdx�Cf7ld,H���s*��e�����u���� ��Q��id���.e�j��Z)Z]旬��j+ȭBv����/J2�\Sʢp |���]G��w�**���QR͇��y2��^��,b��G�rHi,��MP�����8tj���ʹ�7+o ���) �Vrt�������T�D�R�ũ2�L/`�w�J�Y��^�[(*v�~.��W��:�f��a�U�+B�؊����y.�f9Z�,-�+U�xp�n5:*!nV�v��f���Ŕ&�2!I�P�tg`����#f��C�f,��#eD��yy3p�6�V�XYۋDZr��r�z�tc^1_7&i��G$���+��+]�Mu��T�m,��2����I�4�-V0��F�%L�	t�4ե�ЖUY����K���\yYPY����.mX�q�a�^M���t�հtYV�[Bݫ(bW�5�e�L�,��=���ǼG!�1�J�#o� �2iTf`�bg`
�LP�9��5���nU���4�ٿ(�3jX�=ʕl�7�)M���)7ɮҪsZɸ��� ^�U:�EGuR`أQ�]'wL�8�N�Ҝ�U[&���*����i�{��PFX!�5!v�b��˭�'
�f���s	'0�
��m鉚�op�R�RE6�Y�����fC~��̬��̙���7P�Z�����j��Nn��&��6P�(�F�i��Z�����֪ͬ�U훵�*�>%�3%ǒ�w���2;�sl,���iT�Z*��u-{%<`���.NI�mK��2��Q�n�wV�v3��p�ITݻ܎����Ǥ�+ڌX�����Lvt������N<��U��b
F�X�@�6�\?],f9W�kܥ3`K.�r�Kj觏^)6�F��*�=ME���4��,f�y.�P���iޒݲ*.j���p�ժ�ڂ��6�u�<ӺX�^ZەOM��*]��y���mSEZ�����L�B8�5��ML��t��!��%V��9��ǫ(]���Umbt#K/�P��H刞彛on^ً%� �r�1�m�6��������i��S��e���D��Y/2�VNK�/r���m���W��.��P��j�B%)$,�;�(�z<N�[yԝ����6�Z.9�g+C�xn�Gh�wz��\r����HF ��j�RX�B��)�	T	�P��٘,��h��Q�TA|I'h]=�M풖CN�]RMh>���$}HѴ	x�-�b���\-�,1(��+��ej��R��"�<�b���T,�Y�����&9�A�P�����ٸ�J��O.��L$J�U�l��i$,UM
��v����H�T�Ī"kn�<��]�]�b�V�U�)u�oD	�����&]F����*�4icF����F�([�).��i�ʂ�Z�%۬�q��I��_�y��9���Y�\%Di�F����Y�.����Tt�f�-:����n�i귊� �S6�gR}:�b����r���:���נ�s�I�s�7R�cp�ui:*�M%��"ϢL�Z��&�
-,�P��Z̖�3�H�����q&0��ܫUid�M���OTI���&�4�jh욣$�֍`�.Y��bw�/��"�N��S�5ڪ$R�vh".TRZ��Yk���2�5�i�Ya�P���"R�#ePITb;�� �Bm*EB����DR�j��4��ҝ3Z�63��Ư/A&��J��j��"b�������j�V�6�+w"ȕ&�"9�r��yt�IV�k���}U��֒	��$4Ko=L�Iul�J�"
D�W\�RH���0����D�Uj{x33\�z�1�5\�Յ2�b`�c�� ��⡇�}ׇ�T"�Q	�4��p5�{�Eva\uH2H�$!|Ͱq�B�o$m:N��ֈ�jЦ��ӢXyD)����S�R�\�c+�5{iR�J$��ֻ/��q�@�܋.\�D�j��UP�Z DZf��#��S���"T����tyT��N*Sn�F��V�>M��'��B�3��V�ŏ'����Q�\�i(w��M-�wb���֖(��ĩ:�*Mޮ7x���2�<nw5����2��{r�#)Kβ�h��:�紖��m�/:�5=X�J��x��¡�iZ�Q#l�Q�yr:P�ֵX���֝�c(���M"\��A̬(�8�W5ܜQ,�q/��V��A���k�4uRU��A�ņ�sUbZ�Q'jR�D�N&I�֩-Jڶ�6�rv��ڬ��$�X�I,\#̮�8w<X9�۹��)��ȭ��}1��7QG��1*_Z���8��:��q�+q$��Ŕ�7�RȎ,�ڻ{N�W��D�X��*�(-��f�Δ��R[�b���Sj����%J�����lأ�����*�60�Wd�b\��^����kJ���v9J;eˉj����ظK�-;Lj�;N�ii$���iMK���\�ݻ�oJT��$�H�/��|a��i�N�����)��+�\�ʁ�2�3�
��>�@u�o*w7Y���2?W����[��`?���/����3��)8��~NI$�I$�M�`��ZX��'��8�j����r��A���n�*�q)�;���FM���x���װ^dE�\�6���"�y�'���mo��D�ނ)ה��T�^>MD��5ݢO���W4:A[L!8�:���I�"���k2�=����]�4�*���ʫ�-�NE|�A�n=��P�e��{{M�ܚ $Ԫc���By�C���lwҎ����U��3;;R�������`�U��(wR��t�['W	Ũ�ms��K�q��
�r�w,�+	��q��>�M�{��O�&�қ᝸LT��Z#0�d|��o8��y(��F�AF���Vz&��-c� ��wf�f��{ ڵ+���1���t��+xw�隣�n���L����.�T�@���W7�X���=�]y�H<��<�0��a�՟A�GV�����c�;;a&��0�:Y�VI��
���IG���{|ie�]���u
����=F�;��̇�:���Sh�,uܸF�j�;�U��g$�ݻ]J:��wΰ\�8�;��2��7�G`klt���F'b٦������`9�D��{��6dp�[Du�ãY����ʜw)*R$���M�G׶�����r�X��R�1��-f�=��\��%��3qң�5��{�q�,���WSy�J�5c�Й�έm]��uŻ�/�`y7��`�����¬α ���ʚIʾ�C�;AsxҺ�P{d�Q}0�w�,�4l��eJ:2vF��hN	�
�����{W��,�����Ƴ_	*�>��p��)k�%��*R�a����ה�V�G\Xn���:9Vlh`����Q�F���.ѣj��hi�����=�ܹ�
-��Apq�v�Z;�#��['�ʰ'j�z�nH���Y]gS#��*�S���-w^f�$�����2��N#�2�G;ywW^�(T1���ݰ��s�(Y�N.{np�rT�#Ox���)GbSY�3�r���;N*�c��nK�ȇUʉ��VU����z�J��Hؖ���V����H���j<�@�FB�㓕���:�|���w��۬�����
�p���1׭$Fh�7^+z8^���V�y���d���8⎹�v�r3����o��OE�W-�E��|���v9�B���$�V�q�W��'Ϻ'�T��v�6ͪ:8o��k7t��mU���Z~}]Ee�0������0q�y��k	��Kk��Ә�MD��u^ms$�4]����!ؘs�kVܵ[��5�D�t����>/w�	u�.��lݒ�;�Q���
6����T��V䠹��=�"G�j"6Hy�:�v0|GCAPemӜ�Ѭ�K��F>4�0��9*qnq�G3S��=��gB�D�x������9��
�4���;q]%�Dt.e�r��;�e#t(�K��G<s�K��,�I�f�����YZE��D�+��d�����$;���ozJ��m	N�ۘaa�+�n��m��zUe.��T�X���nD1Μ��\�2�]t���쎞D�W7�^�>�DC��wG5w��2��֭�6jUU17�Of����0�����T�87��NѼ���s3.�-v�; 9w6;��H^�tU��	(����&��
V�嚌#7��ؓ���ؕ6v�5�;CoG<���Y�S�r"����i��A�뼵�)�4q)Տ�ͭ���W�a��0��:�;3��;���Տd�����x�޼��=/�S�r��
j(��1�7�4�`�Ɩqv�ej;JX�[ګ����#{L?Rzvb�t}�w�dH|�Y�5A�%0pWgI&[�Pq[�kC�9mL7����G��Zlϧ\oe0$��֭��"mp��_tH7�\F�3���&�U�m�"8�!�;�]���C���9��]����D!���C�Բ�s[O,��֓]$]L�_t�b�׷qv%o���׈�j*�!�E_eN����wT�5�#�\4�k}:n���	ȣ�٬�ù�c��+ar%:��aWj��)�����,T� yq�s�d����ݾ������wM�I�o���آȝ�����{k���Q�j͍���b�Vj��[JՋY7��7k�m�Оo�=Vr����p�9��˭:��Q�A��ܵ0h�ޢ���ksz�{8q�����~#���	�H?w��9�.�ִ��[X�<�A��$�R�v��\�'�7�=���&���y�X�W�G�as�����Ȳ�hv�e�E�\,f^:#Q��Y˞ZÌl�U��<�D�m34��%�I�_i�б<�jU��|EX:���wZ"��l�+x��^<�{m��e��V_X�XU>�*�����kr�Y��<�ֆ�s8�m��0���Jd=���� �ݛ͛�Ф�v���O�#7��І�ؾY�u{'F���9D�-�������SXQ��Y
W�ŷ����	*I���K����imv��5ט�Z[Zf7�m�B�WE� J�]̔n�N�'ov��k��j�b۰�Ϊhu% ����-�uVwTZ�8+0� �;��5ԕd��z6d֮	W-���}Ko�A�H7:�#���Ѡ�
��]W[n.e�RC9�3�S8��CWƀ���-5��=�q6��;R�v!�������7`���I�guiwfW!�8�V>�����V8zN|�l5f�7��Zu�:P�-�H���:J��]���V�����S��u�&=�]Z�L=�ވ�.W�����n��QJk6��_�<"�Y]�I�mdͤ�,;�,T�jt�򩗊�Iv�Ć����r�k�i�:�{�Q/T�ļ��jQZ��x/8_QQ��}$2�r�:�{��v�x�衾A*[�.�%Օ�����k���^�W'��-0�����-�33�.����[e�wys�F��Bo9�r;�����,S(Y���YkP9��]�ojtvܣ�&���ȓ{by��ok6�YcP���3�
����W�{��/m
�gvG��,E�S���+[j�q�jSxw�.J����Y{�n��Ql�L�fsT3 �HFe�uD�w�\��*f��-��*�84Pe�r9�T��Q�Uv�C�9ř��WMZ�.��c[��- R��m�*��;i��"p��L�vc���N�EBS4�����
��2�]�bQ۵ln������U�2x�V�UC�4@�7LDr�N頷��^N)n���rv�D)>�5��t�,�����1����9��vl�S�Bk��f���2NM��M� �3��]w,�R�UEu�r����u�J�Ѝ�ֲ��3J�����'vses���E��n�r��C���Bl9Q-����8�^.j+��l�z��K��=���Ewk�(�+o��^���0�*Ĳ��1]=]�],]�g-ᔆJ�+Y���^���	��ۘ/l@�!n��!���iWn�rd��3���k�܋���WEJ���ʖ��&B+	�a�RK
9����<�{Fm܊`݅�Rcok�C�W<敗�M�y,*���1������0e�2�h��l����I���R��ҙ{�,vWE ���4�v�g<�[\RK_u�z�^��ڒ���a��jc(��E���u���h���o���J���hΎugWp��{��@��iiG�7��.Ɔ��+,r��
:�:��b Wt�ُ��GO��W�| �W�/ʢu}�sٓ��%�&�[�\y�ݥ�b:]
k-�;����a�n��u��z�u]�.n��Kw�p���F�]��<:��avf�L��bk�8����AS��p�IJT��,{�*��@�sCvZ� )W?���e�w���9d�;��2������(�RB��U�SSsτY[�Fԉ.t���YeeV��Y�+(���gXR��oI�{�Q�t03J"�͡�.T�K���7m���{R��cQ�`ᴲ��_h�xm����l2q���HѰ�<z��
f*�����ZݼX���������B,���IVс�f���W÷�._dx��v��S�3)<���h�Z8��0ЧHj̶���Q�]�s!;���A`�������#ݶ,�[N�n6S��W�����y',$umZ�������+j���}7Wr���q]�f%�!#'b��uR�}��SXiz����K�������4�ᶪ�P�x%��(�]����r�ݷE`��7ܖ�#�sB\1l�d)͵�1��QN�S|�[f�|�^����
��p�Jd�%�ݫ}*ixi��S瘕��M<�-W{�������E���X[}T��z�<K����ZEc�g*'ϳ^�3&�uvw]�\�����}��-�}����T��Fs�ʓY��U���׫�޵����M�T�>*�Ҟ�H^#TQ��:��`������+v+��7�	�cFv����F!t*��ؚ������׍Q�\���f�Nw��S8�4O6�)��t��-k%1Z]sk��J�p��ށd��X�Cm�{�u�x�ȕ�����V�i��d��������pyPn���R�܎�ݼ��֔y�g�W����Xc�ܴjc@)����^�AS�]yW*���2�zn4lZ���И)���#�<�j�/-��}�e��ڛ7�e����Zf�kF�g,�Cr���\��ة]��fa�Ϋ�ε�wSm��9L�Y���:T�|��W;4��}�ej�T�\�)��F��.ݜ~��lB7m��+3
�S۝s:�[�����J��+���#���9(f&�/��<������Ȟ�+`];w���ĭ6���A[6l�'�MU�U�k�8І�{ѐhgd�s:�෩�4�3Il]�M;���X;�P8Zam�ù���;��f�e�����Bս��`��(�M�Iz��ݶ���:=פ����[/32�m�3��.v�yV;t�Ê2YY�r����N�ޭIR��V���(���N�-��5��M�{�h=��v�*qt�ݮVٛ�t��u����P�]�rL�;C�gn<i���I �����ˁ�L6k�l��nn��XR���{��˪�&P�)�+�r��P��;6�Az8)����[o"�38��S�3�Z��J^��͙Y{�MFrp�U�N���f�uڷy:F��f�WpN�r�x�M��uǸ���ٌÃn1U�D}�/DӹB������oCQ3\��zv�\�|�.hwm�tt��O{�0�2r��:�|��Qf�׶�u^e���$����I-��_��u݌���$a�Q�]�3̔)umA��E�9���æ�\o����]����g3�l�͆�P��%�2�p���z�ݘ�l�{������*��Wlolt�G�:Rf-��z�K�fg���k����c�_T\�d���=�/Ak8��E�m����$ν�����6����!-�{�u%)��ùդ�.���rF^G��ӇRZ����1$�s�<�`�����+�	2^�͋����e�NzgK����ۻ��������%���:J�&ۉFQ�!J�\d@�,[��i�EG^�2��	,Pb�Z��m�!4"��nq��QȈ�1� �PGY\}��VBB�F4�@Cm��DЅ8#m4$D�6Xi"!��8�P��(���ɊG+�-�x�ލ|{�<���r�O�EBK8���a�1o9b��ɨ�P��$���h��Q������E�(G�WlPtyJ �H�l�T�hF�(��-�",�Y��eQT���ׅ�9�r�(�B�5'1�))nP�'� Q�I*P� \%Dv�˰�)��5X��*p@&`�}# L�ҍ(����iF�z� �Il���($]�0�,�O�"�ΰ���%��Dq@K|=�r�1+L�SO�m��.���U�A�!����'�W;��'-k��$�@L��'?XtE��@���%����d@�h�UC ��g��DQ**��Q����������>�^��z�}��ڪF`��e�Q��!���1.�D�L6��J")��n�HҢ��n#V��;�	 �mJE��P���4,�ذ�ܧj�,��uD��@6�IY�$*8m4$D֤x��m��U�`P*d$,�c+��&P�>�ܠ�f5	hEêM�\��8J1Gm���!f�de�as��!b��	ڇ��<\ a��8��J7����q5L�v����edA6A`(�Ɔ1��#
.>H�GTK
����-Cr��-�7'^�w\��G�&*���m�
(8�<d�"�2"Q�@i�y�v�h�F8E
*�1�6�@d0J��F�r* �������A D��O?/��?���O��@�����������/ۿ��Na��̟����y�'9�,��Ǥ1$E䫥˲"���M�D�c��n��7Q�ΰ�d��ѫ�U� ��mb�ޚcT����GX�`Ý���f�oU��i^�g�,x��%(��Y�Z��H�Vnʇ�Ԛgn���1W|1Ψ�����v�bo�&�����v��;p��%����v{3�oX�,�]�ӻ�B­���Ĩ��b�pt�^-�Ž���7\F))�ԍ��ė-�=��s:��q�t���>o�c�� �=�5��S;���T!�Jѯ��8����]��y�/���7�κ(������@n��|+q+CL�mjޮy�V��b�6�pNF�eQ�Y���}j�=L7�"qlH���Z�Ӓ̰S�\��m�x��y�-�I*���k�3�-ӈݜV��&9Q�M2ym�bk/�[+$cR�Kj��}z's�]̣u.�q���Ay�ʽ��ך��!��o�u���!P2k�b��8	B���ˇ��-�������0��2�6�;v��J�K592�{�L�Q*��,��uuB��p�驻ǜ��r^�q'����B�E�5f��2�]�٘X2o;&�����ƽ�Oo�kZֵ�Zֵ�kZѬkZֵ�|kXֵ�kZ�ֵ�Zֵ�~5�kZֵ�|hֵ�kZִkZֵ�kZ�5�kZ־5�xֵ�k_�k^5�kZ��F��kZ��Z�kZצ��u�kƺֵ�z~4kZֵ�~5�ֵƺ�5�ֵ�kZֵ�ֵ�k�kZֽ��q�kZצ��u�kZצ��u�kZֽ��q�kZ�~s�s�ï8r޹����N�/�&���g�'5�jEX۾��Y�gV��w�
����+���tpƱt�1ސrY������Ͱ��V/��U �X
�U,�uct���]ʎ�B�����fEyV�7b�!�}T-�F*�U�9l��Ky���"�.Vg(��qe�:�Cl!�����}o�Xލ�i�l�ܘ���2�o�ՔZ+x)��_Y��WE&��Mk�)qMe8��ݙ�| �}�',�:Sc��0.]�÷2r7č��t�U���2wn�LT�;�lV̩���2��՚�$PP�'�NV���qu���W�x�D پe�[Ԧ-�`��m�^7�ٲü8���4��I���Ox�an����=LnJ]v��vA��L�ך)ju�&��6բ'�>������=X�;n�5�e��_c�S���n՛�jٴ��s�Ua��h3����9��N�g,u��]Ne�7���4�J�\CG�B�8\UX��uQ��v��P��y�&���*�w��-v�b��i��wA�amwr��*�t>�Tx����kA���Ic�1ƚO�G�X����a���w�|���ƿ{c��Zֵ��kZ�Zֵ�mkZ�Zֵ�mkZ�Zֵ�mkZ�Zֵ�Mk�k�k^�׶��kZֵ��k^5�kZ��Zֵֵ�k�Zֵ�MkZ�Zֵ�MkZ�Z׍kZֵ�ѭkZֵ�ּkZֵֺ�zkXֵ�kZֱ�zkZ��뮵�k\kZֵ�kZֽ��q�kZֵ��cZֵ�k_Ƶ�kZ��Z�kZֵ�hֵ�k�sM�o�y�4��|V��w�36���2�w��wjǲmT��/W=��o[�W�-�|b�źs�z��ѹ�0Ύ��ݣlZ3���E�(Q�6�:І�����\N]y}[Gu�]Z�y���7u녙O7R"�a�f��;w�������uMN��ӓF��Cvx�[]�R�P2EM+;x�A0W�2qC�wS�wE]��)k�mA ���Ų�!y�8�7IDs�������^]�7�^=���zNx1a��w��4<f�u�]�hmV�C�d${�\��'3�GcW=B�C��]s3OQ�ăêHٹSQ���k���Im5��L�y����aSk�l�(���	��gb�ӷt����_R���q��A�ԫm-)phe���czK[^z@�i�dUU�aXq�38䫊fTɀ�i��2��㛮wR���x�WI-��뮧RDUf��{WÈ)Φq��n���(��J�yF���X�������#T7�Z��]ծ���}�)���^�.��c�ǎՙ���1����P&dI5�y未�����\�K���T��o�z�����]�->���	����C_()do���|��?�����ֵ�kZצ��u�kZצ��u�kZֽ��q�kZֽ��q�kZצ��u�kZ�Zֵ�kZצ��zzkZצ��k�kZֵ�|kֵ�k�Z�ֵ���k^��5�kZ־4kZֵ�mk\kZ�ֵ�{hֵ�u�_���Zֵ�MkZ�Zֵ�kZѭkZֵ�hֵ�kZִkZֵ�kZ5�kZֵ�k^5�k�4�7�7�7;̸D{mwC�o8J�dʏ1��ZHd�B�b�lw��ԫv�IKλ'�Aԉ���Jf�Κ��J·fvc��}5\π;X���k/��\�����<1��2���D:���h�;�GB�_�*�5�:>+
�}vs^&3���J�S�mE��Vq���|4�2�yA�ޡp�BGH�CG�Y�)$�������w_ΤΥ���]$��n]�uڔ��j⹙>���Ql[*D6{�Rife�@��bb��C�<�ꦎ����]��[A9�ǵ%�*��_b�^�Ŧ!�f����8�B��p���<=�U�O �,���/�����[�e�B��E��;V���x�cJ�{M;�|��!8L��cm�D.(3Z���@az9���O��4q�?��[�&-d����d� Vw"�(��!"bu�`�E9��Ձ�]f�=������28	]6�*��`�x���c9��ĳA:��3|���H������K�=S8gs��Ƌ/gr��}Om���[з�<�M[ڬwH�NM������60��U��7T��y/��)�/a�u8��Ӷ��wҨ �gU!H��B=1��ﾎ�+����o��kZ�k^5�kZֵ�kZֵ�k�Xֵ�kZִkZֵ�kZ5�kZֿ׍kZֵ�Ƶ�Zֵ�k�xֵ�kZִkZֵ�kZ5�kZֵ�kZƵ�{kZ��Z�ֵ�{hֵ�kZ�Ʊ�kZצ��u�cZֽ:뮾5�kZֵ�kF��kZֵ�k\kZֵ�k\kZֵ�kƵ�kZ�kZ�ֵ�{kZֵ�w~h��;����>Ny��޴��j����f�F��r,��NYv���U�r�W�"�5.��/m�-0K�oe'q�r�H�ͽm��R�:��&��,�����L�'L��49:��Tt��çPU��F���c{�E<9�p�ٺ(�6�0�Y�U��:u��9��"4����;s��;vwa����,ˋ7�b���#���ֵnX,�Ucړ{hI��Ԯ$fv��X��{]�p�^UT� �)�� ���/bj�S�T�y��v�J�c��XmuF�mc��3!y�t���/Q��1���|�����h���+��͌����n��=�Ņ
t(����M,��}YWΗ(��	�)�`m`�U��c> �EZ_?{�&�]�V�/۪�b�|�B��8e��mX@���0�恋��G�)�]&j��Х�vv�ʄ�=[�&�ڄ͜����k5|��X�G�bAq���6S���^�,::�;��R�"����8:�Tz� ]6�����d*$�þbtKGw.����gt�:�wj������"�vz,
�x��B8Zi����Q�z���9�;�h��ݧ�w��+.e����f�z��
�qg�B�W�Ĳ�l�kFt�>��e�$��O�Y���Ź�v<8��\5�k,9���zf����Į� Y�����6h��٧�� �!5
}�AvX~�x�3z�&�UԆ��4���Y �DfuU+��:%f!(�z�f��t���a ��!�_p��X<RB���W�7]ݙ���=�Ү��̩�<��+O8��NU廻}�1w����ӆ�g	�Nh��g�
࣭XF�go���o<���bO'^u��*��&��J\E=�;�G1�Vi�#�z�M�ΥC&����g ���/J�s�.�����֝3k�ƛ�5�M��Eᗸ�0�����E
�7^�WJ�1cUUvR��#�Q�z�Zu�(6�mk��ѭ�0���2�4Nq���(rP׋E��b���L�=����+��R�޻���:9cd��opq1�*��!�����8��^ҿ7�\�{��1]|�WD�/���E�{}�� ��c�kO78�Ϋd�XF�d�/��\i�@�\���:r�dL�KU�/�� 3��;����N�ݹUwba�y�Q�xŚ'�b,�fq8�q�)]{Á�7���v�Gs#L��~�ͣ��0���IVu˽������o1���,d�沞#H[�L��E<\i cO%hhx'Ƚ���^�%}�5�"���s�v0k�C�0s��
�nշ۸��n�+n�2n ^A;���6+6�fv�ɨ-�W(�b�є	�;�Ͼ���L7y�*HQ]ʼJ�t"�i���֫��o���������"��]��ü�AnNos5^>����tR)}��Y�:{�+�x0b�Ǽ���
D=�L�/_bc�M���.��E�T���:�x>rs�3B�W�4���	p#+���_LaM�8�׳���47�\��q�Q�x����le4�ԥ-��VJ�Uk��Ho�=�B��i!vPW+{�ݩvK���wʫ5�9>����ى�i�����#E��W�W^�v��UWk|�>�ȷ��t��D c0�v���ܵ���Sh��k��H�;�t��s�A�]�+�*-��cR��@
���|o1�b�9k����j��P}�,�K��,��B������"�-	�#&
�\��f��&]���ʘ�s�|��e���[�fUR�.��:X�k�kXN�q�:ƲE�2�������(s9����[g�[כX�ݨX޽�b��c�%��<9���3=��ﯢ�SJB�u�XD=-D�Ӹ�t^�m3,JE�U���Xo�P��K�4 3p9Wϳ��H��{��h�s�-}|�7ǅx_�ز�US�')C�S���;�Ģުו�㝕�"[����o;�Yr�%�ҬU'�,�+yQ��q�A��w$�9WT-T�R7A�+>
�WB-��|G8��򆊉M�:ǁVM[�Us��ޛ��|޺
���p3��0�]��Db�Y
�A	�ի`Fn<ݝ<���K��}A��B����]���Q�ܾ��Q*��t^��HJ��+m��.&	]H�9`�77��k�Q�v�]a`&���|Ӛ*�T�Hz�J	�Y�,JS+
�v����R�[��lz��]�Aw���;����E�d�E�U�C4҃3���]-BM��� �l�b�ppH䦒)nr�]���UL]0!L6�L-�u�뷦#b�'%#)2�r��'.n>.F�<)Z��*we炅f�n�(f�(w"ݙl��^k�uliZ(mj�ja ��N5��b谌"�]��:�%2%an+�S�w��(���u��]Xڜ�靝m*��U6ʄ�"�	�ce�f���uٚ�b�m>Wo�3V 
Yt:Cx�;���5x�;����By[[��+��ne�"�uM�t4ދ���8r�i$�s]�Z��7]i��Lƴ�J����Mh��P��&���6���\�[�{���Y��ڥ�V�ʄ�/�G���*��1���<z�S��C�K4-= �iqd��X:]��4��11�S��6�l������T�u�'X��è�l���#ՠ��>�j����K�y��%���8.�X-d�P�E^�r��o��3���T�����ڜ���Kę�=�2hR��j�].�B<�F��-��^X�J�\3w�ly�����i��X���,\�sK�FT(�yv�;�#gT����L�q�jfl��I��.l��d��a��n��2lsio=E��]���{�brs��w�0��T�D���i?}TQW2���A�)��*��8t՛���xq�G�ְ�Wz7 �/M.|螻�b��b���}O%�o��}��u=TW;�n���I�w��0��ca*n�A�V��I�5�i��l
y�,O{s�煲od��i_�I��L�kX�y���^x���Y�K�z'T���dGv�/l�Mv��\̮�kuǗ���ov�gi��y�q������-Cªp���>8'gb,#��8
]n���a��F��jdi/�g\�黭�#.�@2ɹ�ve�6֝A�s�lV^e��`��j'$���!q�b�)���^[5}�g����/����5%���`�=�Y��uw��c�����ȗ�/q��0��Fb���Tν˹8j��MJ���%������k"O3XRAo���V��z�w��Ι�n��Po
�zod9Z���Q�<�C��P-aΖ���OfUP3��0�q�oe���#Zi�dmm`])}���V���`Nꝭ�)Q��9����rb��qY�Dwiͬ[��ŷg����ľ�̩s�Řx���'}��1S��\��P��u��;̹��W[�:gK�"(v��%���4Ѫ�� 8��,�2¾4�2+Vj���q]�v�^;o�n=��1w�p��;�z�J���$s�!����0�ބ�1g��Z�i��egq���Yԍ�[E�8eP]�I���,�y?Q�򞨭�/GrC(E��C:�+����Wf�+O'U��A���(S;2ț.ge廤�7;k��I�e2�ǜN�J�W���S����h˳�:�q�yL�#�5`ut2^'���5��aWsz�k�Ff)��D�Iѩ[]�S%m�I[�@iK���
�����Ɨ8㥽&|�-��#"�t0
>$������Y9�������( *�L�����o�����K�+������9���	�Ýp�o!�&�7sPp~�AS!�h��<�9���I?Z��BQ��$�$ģ������.CE�ل�B2F"�ؓ�� �ځ��	#1N�U
�$P��t��J	#�@�`��9:T(�$m� a�M��18���Ah#HN?ؑѩ6���J�2B�h4�Dː2��Ƃl�rk`�@�̮�EQ�ʛ�����fd{ph�\=6.D6wW�8<]C�&F�R1�}Z�Tg+����n��Typ�7S���rݽlQ7uܔ7�-�{j�����n���h���r�1<6c�f}��:��n����W����EQu_I]vūx����먇*�*����O�ʠ��y�x>S��otNK3(�Z0g)w<��gKi���´Q'v:�ށP�b���ܮA��g7[��"��Y�U���v�˳��G9˻�Y��RS��Ne[�Gt� �t�.�9e�ܭ�Gv���ਜf6���(Mb���S���䙑pǑd�j�,�9H+!�)��v�u+gP�U��xv�Qw2� X	-���O�HvҖLC۶'ӊۥ�j��$��-�+$w��KöX;�KBF�6�o��T��F�`j����Qթ��S�I��򾡯ud�?�+f���kI-�Yٟ@ei�)^nΧ��y!"t�֛�Ut��v��Joӥ�ɽ�^r"ﺧ�-����N��]��<���Iz����}��Cj�X$�'Z�0�D�C��:�̡���}&(	NFx�cĢs�ea ��`P�	$!R	��F�L6��� ,#MHA||e��P10�21��PƵ�Q�A��P$� NFЉ�(�J@�N6TjTQ)�UM�ꌢT@�L�AmDb�%��q�NF���A"F��[��	)6���
�p��*�\�9m��eD�	1��:f�C�Q�Ӆ��	B	ģl�"�b%�B�f�P���f0X.�y@�2�T�Cd�H@�|�0�\RbQ8��lH�\p�m
%ц8i$ n&�"��]� ۆ�e�a��d%�L���ȅA	r"�l4G�w������}�u��U>$�<�+��A�rT(�,ɞ��9h�O:r��c�]~>?�Ƶ�kZ׷��������~#�
��"�J����}FT�@�ʊ=��iQ�k�\ȹ\<�H��͗�Z<uֵ�־5�kZֽ�====5�ߟO⪢�k
���t��
��.�Ჽ�'^�Y��\�&�r=_�ηooֵ�|kXֵ�{zzzzzk_����ET��׸.���p�Ru@�s��y���t褄��-"�br|�8'�����h����L,��s�����������cZֵ������}�yq���;�s]�=�c=mL��׽#� �!&=҆�~݀�|�4�y�BT1$�|��B%��A50�TP܀p��T�%��vq��OeېܽP��� D�CB[nxN(22b�a	��q����؊J�jڻ����M��s�c+�ب!��N랚��$�J�DIUP1.E2�فLDZA���)�Qy#�bp3���qK�+8> ��3�G��W�N��ݹ�����{b���v�l��ǜ%���|�鶁ju��u�v�����!lT��������=q�T)P��$��N��x�wQҠ�_G{��v�s����<�+�8�����Pe��"�������^޼�Oz���M�i���=���/��`U�;���ι��l�pr����HRn{���8�\����ݑ����0��NF�A&�DƐ�NW���w�=3����wrS�Z��B-�,5��;Q!��$1�RAn�N�s[����|���晘]���'��CPI���7�|u���ɻ�H�e������ع�8������)}����E��N�wFY$jE�n��i���ܐtϻ�������{�<=�u̫=u��Bz=�|�|UT�v�|@>#����{�BdY{s���n��U�e��Ww'#-��.e,uϩ>`8���!��ѫ��T�^�E]Voˢ^�:��.���vQ����>�(�W��t}�'n榟-Q�4�Ua�dZu��QdX��@b6d4QT��TEa�)A�����\�;�"�W�ˢ�r�r���)B �5Ʃ�0^���ڪ���%E%d�^U/����̛���/C ��	�g�Y���"x��Y��S��Y:y�%֪B�wU��R���ly�8g�ez�a���½��9Szn�[����}�M���Ki"d-O��7!��gw��
�>*OGY�ؓݣ���3�հo%������6�m$Ei���N2�[���Ƌ ��o�,�)�������54837N�a���<.�ʅi\��� 8�L8��ꦽ�i�F���L�)���
�g���VQƕ3�ů�L��1w3�*����f���,\v�8�ީOa��~�!���=5ك����EL����^�;Ś�5��
�������j�����=�.�+��1*�+Z���H�e��³�����{��{*��5���J�V9���s^j�R9��5d:;�)b6mYs寝�O�_�4us��?V�|���!o5�����W��D���b�z��EN��6�;Mc�+����2!�5����~���Bd�9����x�[��>��+�C�� ��<\7���[)�̲��Ӛ�^�5�U,vV2�T$�ek�$Ċ��D53���q�K������J�|B�>�瞠ѹoo�z6o��_�ɽ��B��6N�&��z��F��_���Z��^�uՊ�{����%�Ѽ�5X�tl���go4�P�zV���(E�\��d~\������xйRU���b����$��ڽ�u�d�hJmڕƾ�U,'X#��I�8K�M�S䗉��)l�h6�Z�R�ô�4\�c�Ѷ��Aw�0�[֚�Y����͎K��;�Ė��g���E�_v�'w���=ͣ	ݭK{��;����|ˉ�l�����R;�v9��7+�n�1'y��'B�����;�( x@< q�������f�u�hB�Lk�=�,�kQ���_�l�����l�d�7,��#�^S6�{�s�C+�rccf�@�{#n<T��Ia���]�z��GM}���H�4��Ź�<�_�ͼw���Y6�� �4�"Q�c+Iqz���Ӆ ��Wl�g+<3��ǖ�[=Ey�'��^�1.{=$�*�(^f 3��@]������qנ�2��>��4}�(y��h��F��ޓ�Q��=RW�t��`A�q���\2>�/'@�T�z�t��3��C�B���ّ���!��#k%�t�����+Y�Tx�;���������ܜR�����I�/�;�#P�xk]1;Ee쥧kuTS܍5P�A'�b��zOTO�({��џB롲���N�c3	D��4Efי��F�c����}JFa�nGh��f�Ϛy���b�fm�jc�3 ���9K
����ro�ê�~��a��0���fSo#Њ�\)d7Wx3�����{�xd^[��T�3o���͛n��V�|7OR�� z���/l��o��Z�L�Zyd�e����������������{��^� �s�l[�R��=�SB �-�]�d��ê�S�;�Y 6�Gdנ���z"^%� sڨE�j�"�i�y�z�WU�Y�n���d�?��WI�N�}λ��{��YM�e����EV�b+qF B�@;�S� ^��L!��f�A�T�L�I��T@��,Ri�
��^�m���+�щ�	݊�U��n��č"��rsJ6M\��4�o@�C@�;�}�{,Wλ�\��5FE���0M��vu�z�ngu��I���|�����ͱQ;b��h�gѻ��k�θ���6�%B�ffl�g#n����qx��>��M>[e����Q�-�������؀ږz��Q��g�i�L�����D=�q��+Ҷ0���0%�ԕ)^5�>&0����Ϳ{�ǜ���ч���*�fe�lY���,��(C��1^��z���n�:
����,�Kr�|�ct����}�3�=��˦��$)#M�IIN%q��"���UA	�^3!/o��	��ޭ�;;��d�V���Cʗ5�37.V��	{v��ct_V���e[��7\6�k�)��mbd׈��*!$AIg�����ҧ���� 9�� ����^�ܮt�3��uSh<�k��|�ʈ܍^uV
c�,�tx�� �R�02@���wf�`����Uyq���^/R�좇^�{@�/�z�*��5a�̰��Ԓ�0�`�%��]�F�btB!�ؘ��ɰ�lAa�&���'p�Z��UQrJ�����%8��Duw
�Ohj�5�}O
ݷx�]ٱ�*�V�gG�j �t
�Lzo<sۻP༺y��1�Dc�/)��S��;��5P�h4��w�VT�,@��V�͏��ҳ��M����=y��:��3�R�y���{���U�t� �%��D���4��]�Q6�v
����.��,���R�cX!��4F�u����Ayu��D3��G��]{ګ�ӽ�V7���%�]�+�`�{���*/^>&6��������nh;����G5daHJ�k�=9����{�"�
혼(�|��b�_To=�3n*����]d�Up\w���*��zХ�Rܗ�;a�P�l�����eY��c;-d�Α�0��3\���My6�i��yd'Xj��ɺ�����A�X��_>Ц�cB{
������X��foX�p<� ��1��z�w�]|�o�9^��Y�"�E����k�im$A��>ʇ�lu(��V�.r35fC/��vk�S>+�k��Vmr~��yN�e���cy}�n�(B^�id{ �ߣ�O@�3P��j�裙��}0�Yf4�ڹ�����:��m����T���x�,�S8@�������11O��z���H0Y$���h�X���m�P�1y��7n����6MYB�2�'=����l�ak:�9'✚�Qhٌ;�*BVeR�R�^��B2����t�o
��� ��-���}F��(a)y���DѺ�1��5�Ӿ(����C�I��y7�3Y��F����Pբa�ё ��Їى(��͛�I��L��b��_Gzcp�t�=�#�OfR5J�������O�DN^��'�j%4۝x�;��/4�Y�}6����F��+!��;�M�Í{���oL�Q�YG�N̉_B��p���{I=X0�A}u�?j<:��Q��Ii�*�Y��3��ծ�U"ۥJ�K��`�W��S)j��ณ��� ����zM���Ě�׀�V��۹����AT
P}�w��ab�=�n����Ks�{hו���P��^��W(�5Vi�M3�3��
VH�j�7h\޹mIY�+u8�Ǵ y�5�E��O $�P|�ۧ��W\|�pg�d˹�}ѐ>t3��%I��l�	&�5�����H�1�GkI��2C;�33: �d9XЕ��q�y*�[-���&F��ަw�Z����w��3�^�gF����u,��ܘϟ��������T9��k]��;�'�J��!������;��o=��ʎ�%V��{ӟ�RN�5��VרC�z�=3ߎ�n
2#/%41���VO�'��mI�f��{���Fs$7�=3�8�k[�h%nR��ķ	�E�Q�bf�"�䁯�L��rI�:{_5����*�|"���f��Ϻڈ�P��z��4_Ǻ�x�գ��rg<�k����������^��o��D�ߒ�2^z�oo3�[,)gp��:�������);*�]�x��t/��1�:��o>U�&��~ �����ڭ��t������:�[)ԉ�Ag��w��v��W,��v�kaÇ�����W��3�!i�텣}Kn=��D�g�YWc�V{f��>Jzw�'wr^��v[���#�1O�*�m:nE㠆����NI��Y[gpYв���1߻���PbՏ���o�w]���_�^�Zj����2I��v�TK�o5O��$��o�nj��VF��e^˯v�+�}w>�%�e��E�����̘�sgq+�,3j@��S���Ǟ ������C9��z� >I�^�*�i���}�������G���_���s����N�6�<�s��.��6T&�x�tY�l��FBuwc� j`勾Vnw�g;�K��離�[ޛ6��u�Ȓ����a]g�k�z�煾�T_V�%���;*�d2�V�C�Фnk�6's
�F�Ez��燪Ŗm�+��*�4܂?I�Rk	8�&;y�����Q,'���aU�3P�II/�LEt�+�Y��ʏ��ޛ{P�"���$�
��^3��B�-1/��y��{wy���og9�s���>�IF�m�d��&�U�H*tKjśm�G�����������3�.�
��W�9NS����T6���s�d�u�n?r��¾�YI�ߞ��yS�]�Dk������=����U��[(B�d��n�Ea4�NM���KaB����mb*n=�YL�6\`jJVF�I������ڇ��X� ��(��@��ȸ>gB�^ ���� ��wv(��Nۄ�դ֌�y� -e��ty��xV�H׆nF�D�'�����&=O*�G�Fþ��юz��X`��E�"��mYR��R�V��m<�;��Μv
�޲��2�(�6�Y(\��{3h"J#���VV��ރ��Kd�����e�ᝨ��b�*H�����&�(wa�3kSY�e�B����i)zG�x���J��m K����]�N��W�\����gڨוp8�(��1�rf]�R&�;o�`�_!�W����� �O�I$�`�.w2,�{���Y��:�1gl�:� ���x�6ۼ㋱u����WT��nڮ��z��������|||G�1����nVک�$
g#*Tyр�y�� fA1��)�A���Uk#}j4��۹Lk��v�I�O9�u��S�"��W�[4����[����RIkmk�Z�JP�<�8\�*�����r��gv�!���uxك�;'M��K'�J��L5�Y�,�b�2�'M�+p7�A9�o�Ly���@�X�'�S�7&��k=\3�ӘM�%�͢��<4�����U������T����Y/c��l��vh��%{{UPK���C%��o�0ZdDe�z�LĒD�؞��$ڼ:o3)�W�(��o"�|���nvlS�.[�n׺J;�{�{)���Vc%����C`�r�j?�my�F�nn�%L��Z|��A~��y�01���} �g�gCpg�?��A����osH�"��P&��u3a���|�zV�N��yq�I&�s(�!T��A��p����=:�f�V�o��lM�y��A�Xo�{u��A�\��Ż��͆�r�͹(���[�:�e�t�w7P��sp(��/F]e�"�%�����$�C5�mV�Wȣ�Ԡ��ql�yݨw>���*����_���7�ZC�I]��mu���ԍ]�!�Ck� m�X��Ɋ)��$m叭�9��Px^2�SQ���e-T�W�����qoL���󔳯��#�P�si���ٍwp�lv���r�]$���D�n���h�<5���×�y\���P�{_�کAr7w��!�f�����1�d�QG!Se�^C4и:�H��������U �҉�<;�H�����4��^����j�oD�N�2���e��uC�mT7���c�VjogX)��r�`)Ŵz�k{�5,�e=B�J=�Ҧj��ۂӦӇw$9���5�u¡G�t:��y\�[u�����i�vT"�]���T�~x�_NZ�|^��M<��f�4�@,t�Q@������̝3��ˬ����ո���:�S/g�Ӂe��y��[q�&�"ٺ�H`0�f����J3Q�cv,n{
9Y/S$�FnWh��������VI�⓬:	��F���M$ć e�2efk,��j��0^)N�_��n�!�k*��B�xݎ�ּz�d{��6��r��%�/�Ӷ�*��9P�{�\o;L����9��v��wk��ev�)��۳Ϡ/r�\r�C�ɁQ$�#���S��T"Z�#~#V\�-�jd��P�K:;�E��b��;�+4m�Y��Rّ�v�Q{!�
��ͱ�闍�Ɨ��k�jl=gL�W�ϙ�i���-_bh��k�D�gR�Ot��Jk��՝���ãH����W�֋��ev-�<����[���4!�V�N�M�=�����Rv�e�����Z!kՒ�1�M���WY�!/s��M_vr��U�j��ڻ�nr3����7�N��p�b$8�N,ѵʴ�\���Q)ң����j̼�*�3�.��4�-�}��x=�u-���[N���,gg�e�H���y{�S��M�wJ4�V/TԨ[G�"�X�Tt6n��C�Twsz].l��7��6H��֕ř��.���xj��R//��}�n�r����fm��E�;���5��n����+C9��+���,sF' �bZ�w'�N��w�9M�����C "���\m��]3���K��T��g,�we��c�Ss*>/�*tY�y8OP�Ur��f~kZ��7���_����Ƶ�zu�]kZ��I>K;���{s÷�(��r��={�E�Z�����r4B�G"�P�l^ε�־��>��>������N��k_>�w��*�8Gd��VY)UE#�"��B��L���\s�"��DrU~���kZ������׏���ON����w���R)�(�|�a�
�R�����v�r�~��@�����sB(�N�ݻ[���߯Ƶ�־�������뮾���yy�!R���ew0�7:Y	Uh%*&�QE�Q~ �*iTD*��AU�'�dz\.[*�Z>{�r;?��D��'�+Η"�V����̺��0	��\eEy��.TQRITtR�
)�I"�N�V�"?��ߤEp�&9	DE�H��PȊ(�eډs��+�Ȫ��Pj�-�Q\��]0�(.�WeA(��9����:9U^u�Y��Q�4��"�l"��UGՕQrL�ҹQr"����HG9sP�	��\��t,P���nJ��+ǚr�K�E- ����3M�f�2�rQ��^�㥜���_v�͙�ܖ���훶��������������?��z�^��� =���p��^�>�|2���j�t���$Ղ�?�V��]e9.z^<�A]W��2�����5������З�zO��zlw'�~�xg}	V:<�Z<A� 
���֯�����|���M�!����j���1ǪR��x�#�-��0�)���a�.2.����D�V� W�|.��������RO�A|f�����d}����s�R�m��Y�g���Z�T�Γ�o<��eQ�o���HG��z~�W��;�`f*�㴟�@3p�B�Kx[�E�/��J��u�ػ��0nzgs���ښAq�� K��M7w�S�u�_:�|���QV��EǃzE�T=��\�e
��i�y50M����{G�7'��%9���Su���mpc����?`0=OB���N��$���� `.-���τà�/����0ʐ9=���Xc>����	��wN�sP:z����q�=�O�=xt&��A�`>5�.s��r|��@A_=2�nNy`d��i��<:f�ق�[��Y���< �q�a��,8��r�p`�g���rԀ��(������I��Q�_¾��>������HNu����rS��z�rp�'7ar{.��[[)I�U>�mLZ�qB|�}V���a2��9�A�:����'.�"s�+R&��
o&��-v��5�L�I�3�`W����Ve
6���Y������yyyy�����pY�f
$���	����P�}��H�YD?ҧ� !i�~kO�a����؁��])㗧{� x:a�M	�_�c�y5�3�郋\���
��H��;�[;�;?=�TN�5����t�Ƕm��	ok�0��xw�=�6r��i]���|%p�u���`��%6��D^�>�ꥅw��A���j��B+���~��s������֦8$�4�q��I��[�^Y�����w����G���{��������1��O�^x��� o��5��ҟ	݉/D��t�;0e�O�N���A������?���~/�j�<�5���.^[�M{������X�8�l�]�s��=����������<�� \ ���G��|�Ҝ.�ΰH��I�>��g�� �Ǹ@��p-�75���������͘�^<C��+��$�L��m��gǐ^��ӁO�z��C�3���ƃ�TA�������t�[����7�������m�9oz����U����wV���c���M��l��.*�s�f�U�/������< �ph@{ό~E>Z@�㖰����>�������C=�����KjR1��m�|f�?���p�9��jh��Θu���Y�y�x��<��5�������W0,�OZ�~|�^?����#) HmA|���p��4\��u��T�Mrrf���2�Ӝ��M�\zk�{�Gv;g;���yOC�K!i�p7����d���>��3:	d��$8j4��L��f<�W���5�kZѵ�c����v��5U�)�N®�^d�UYa���3���]4�)@�|�^�>���K4���"�c[s��>�]X\�èGOtz�Z}I�����RVxx{1�xuu�~�5r{�C�������<�	%k�q�	���#�5�u<���W����qv��ҫ���|w�xo	�ـ���Tj�����/�|�w�H��A��YUM��������u�LK�d�<9��S��b[Ŵ;�׏;�W��r<޶�M=	9#��.�eia�{�!3�7�F� [W��#q���������}�D|>M!�u���D���j�*<6*h�U�� a�T��yN�G�ˎ�x���z�~b�lx�7Z�]cxJ{mbҐ ��S
w�ř�����~ x"��>0�����27�º�58'c��Ǻ{l�q����8�XAf.\����-Lr��������(tq\�!w��?]-:{ϖ���#k�ej��xN�s{y`/-L&�Nvi�̱m�w�p��Hm��O݌i���yiΏ�t�0��@v�d��.q������@�zʕ�u�Q��O{�؟5�ݩ�j�߾�0�ރ���$P��=L���D��%-��~@F��ȧw����?D>��*U
�P�D�g�2-?���g7_q m[����r�jR;�D�v�J}�w�\��f�0��k�-x��7�έA`&Һ��|"�����s��$:>=�J��j�ދsT̆;;C�m{sI���>���?�����?�D���=�5����<�?�{�i`��p�����w�� (��ϠǄ�B-87Es�ӝ�y���p
����_�j_;ɇ��WX��׫(!`jT<�q��=7��^Y��2�gf�5��j�]��A��pp58�����ï
��� ׾��!��c<;���~ڏN0�{��l&�+5t��s�R��Ʒ������G�j���u��0�0����	�j�_�&7V��7��Ϋ�w9=��a���[|�6�uLR�Q�����G��ѱ������h�#Y�N��2�;|b�����-�T��h�������l��M=���0�^�^��"�j`sSx�"E+uRE�܎��ݜ��GӇt=�M�<êc[��9�9��C���1zoU���l�i	�X�����N���|P�[�GypŤ7#"���B~oԩ��sxخ0!�w�	��|`w]���|�=v��<��Y���6�#�1�U����=��e�X)>��k�	�z���|��᢮���t��;��p ����wןs�������DAc���z�	�����"�������]��	���}�)Zߛ���u�r
�Ae�&�T��q����&��0tż(��������U�fwm<�i)-�	> �_���:Cj�x�~�}����6�Y��ؾ����V��+d��k�<�×48q��MI�H&����w�P�~^\\\����� ������o��m�ܥ�l	��c�O��� ��O(E}R�>2ül�5��Hq���b\>y�n�ab'���Ϣ�ō������a���HF�>|�@_oDOqK��D�?Co�Ź'������x��~9�zu�r�ht�n�=�9���	��|�t<0p�sM�v?S^�8���Y�(`�K�j��N�l�zZI�Dנ{|��v��`@ڻ��Ouw��Lܳ��kN�Ͼ��|>x�+�'��'x@W2Y�`�_�CK@RT� �
NDT8-�EG.|��v:�j{�	d�� CB�a-�ɔ}��Uh
�1�ۭ�s{0�;�A�yCT3}��cgo:-�a��:Xp4�W�� A���~C�_
������;�|&�4�;���x��^�]5w��^�`���<����N#����|���-��Ç����.?��.ޞɼ�Y�9dj&�+ᴏ��2̣�(�-����n��=�$�5V'�Z �:5� �x/Ղ���ˮ�;su8�x��P3�:��ĲO`�)�;�N�q��I���Mn�9�1���R�o�,yi�q��noV>�Cy�2�t֟vvK�"��0�VtZ�s-ý��.�����[�$�v��<(.ٜ[��flJ]�HuHw���rA�o�:e����Z��3r�u�;X����H�|意n˩��<x��ǁǏ�ǽ����ϯ�A��G��7�W�x_)�9>����M�\k���,]"�+����7E�����)��$�����%��øli] �S��%�3��'b�<���6?�X�������i�	����C��9N����@|����w�����5܆�9�S��i�������ޤ\�T�r�U�C�f8��V���3L9���^\�N<<��~!�<��?hR�	cW�&P��Ȓ�}m�������y𾱤�*��y��g��`�����}ʃh����`|w� �_v����qj��+�ņ���5P�N)��#�w�W��?UK�/��
�xO���3^���U3Gp��������\�ot~>��Q���:�yX�>�p������o��{ޗ����գ�\U�J�l������-������	vNM��6��נn���¼H��)-��,��p�C�&";cw����mA�qxg!��jtA� ï73��kr8eϹ��L�9Y�snYf٨nM�:{�������>��� t¶��D��\൦�_�>�e(o���|�|4�}�ث+y��ٶ��J���ɼ2�]�A��3U�j�������4f�9Kj]�1�������G�r��A��a 6CH5�*�TR5�80���vu��q�B���cp�B���^�����j�[ܴ��֎�WձZ�/3��%����I&�8Ȉ&�%%!���*HԈ������O>�q��<||�Gp�Gpr,R#>���&s��}as=߷k��ʮ��6��L',܄|:�l���|�,�D�Ն�@w�@KS{���:���XA�d���.r����x�jk�3[�M ɵ���S�k���Cu��A�	�k�⭝�
�6�S�]�h�a��m�v�Ul�U��=�ϸ��3�����eÑ��a�I*��A���r�O�<�ح
���+�]z�W{��U�C��;�}@�~�|`���-
0w���k��Ԧ��c6:��k���K���'��b��|�@OC����0>�Ahhu�ɷ_<� Jp�!�݂,i�
�N�����/�෸AoF0�r)����qٞ_|��\]:��>~�7��Ѧ��&:�^�< e�W����Ec����������x�aYQ��>3�0��k�?��_�	ԅ&��w���8{�ȹn��ky6{�)�{LcÚ{S���s��U%G�?
?���d�}��?t����îmW������6�$0	���_\��������H
:,wBe@�Sǟ�4;ϛq�����՘2�:޹�6o,�{�A��q���O9��r�[ɅQ=F<�,WT��t�T�����U��.���-Q����.����������K=���!j��ޗ�xS�<���EI&-^U��ni�v�q��˴��h��7Z4u�)\f��7�E���"��pp�^d/܄~�\1�Lq�#q��`!�$������]|�G�BxN��`1���{}O����P'���_���{�'���� XM�t�n���ݍ:xm����
WH�<�(|)�B�����vMM�M"���KlJv-O�&��#z��N��E�~&�4��i�ܠ=:�+�ρt/���Z폨�� �Ǒ�c�fk2��y�=u�[�a�<��|�����@��������(݂L���O��|Q��P5>@a+~����\�I�����*��a-�� �ǁ����<��D�C��g(c�%��!�Y:e���V����� �*��[^���-���XO���w�|�dS;�S� �f.����l���K��t�)Fa�A�ڄ�,��2A�3�M]涯^���w�u-ri�ٞ ����2�h�ϫ����W�{i��k߃XW�4,_6}�K�#�`E9�����\\���|;�kOD,1SU���x���z�`p8IY^�3�i3Q�;0|�!���s�ƨ����5�xf�OF�{��fmnZ��Tۅ�K����wux]��cֽ��8�8�Ə2�X�}�P�|~�]�_�{ߣCwW+�U�(����q
�Fy-¶ֱ��3�������o{�3H}�_��{j*��=ཉ>�ش]�Wng'�2�B�y�k9��t��=��5p��o��q�|�[����IW-�O�~��&Ac�<�c�8�ݸ�8vW ���*vX���[��\������%�{F ���\ŗ�������i��E5�B����{�ŵ�7z7�*r_<��M��F�7� ^[��.[�ŗ��k��Jmc�0�����������q�fl����7���������X��L�[��Y8�b7�Q@t�������!��$��J *~���oއ�	fO8�Kh��Y W����c�X��`��p���w2�W��8g�<���m���tx[H秿Aw =tk������z`	l�"[�ђ{���l�@u2���;�{U����=�ߺ���+�#��`�����6���_�R� }���W�^��̼'��b�S��P� ���Eρ�x���F>����nf�Nq���8F�5�@@X�� )�����L��U��&ֹ~����;j�% ��*|�r��wB`gtބ78�l0`w�8�~-�yb����WyKt�zCD��<0ˎg+K�'fgW�^�_���3����-�YDq�7%뗨u�%��  ������~�d@Q��>`����ܞ"oT� ��<Sb���|��,^�T�Q ��?U�*�;f]��
�#�/��[�M�y�6�>�'��%h|E|�<� �yt�Mӻ[|.�JW�bV0WV7��9Ǖ����q���͛��}!���x�f��z�-�K�џ�Ac���EH�&@�0�B@�#�8�U�d$$A�Qvv(.�@Qs0f`�[���\k8bva��`
�^m<⤀�>#�,�I��n�8������=Je��]�;�D�i����٭���8��#�����nC�E�ڙ�2)�,������] c�֤>�i���oss삊+�8t���&
�_�҆����� �R0E����xOB�g��v����]@ٛ����f�F�'�0��0�d�q� ��\���WD3
��+^�
Ol��w�"�3�ÝY�{��[��8\u	�o�d&"�p4x'�%�>�]o�.�l_t�S=�$6,�V2k-��ʷ��k�χˋ���f9�Р��7���q���Ona4x���M��}w+�.�3�mno�sU��n:I�x@?	׽C����c����2�s���z�8��]Ӭ{5'��U+�wn9�qFwN�xax.�2�ZGjy�ڵ�0n��g����<%�y}���9R9;`Ш�-zƂM�R[�y'���>�ӣ��g�l�ou8�����x2��b�!��vpm��l��~~�l8r�8��`e�L	`.DMU�%8��@<���W���4[��v��``��B��V�s�C☿�y9����%�w�J�"s���ѹ�t�d������uQ�8:;�9��L��gү��m�ۋ�)�����-�ɮ[W ��E,c�W��,ŏ����y3-�V�� T��F!��!=z�&�����>��K�N�u5�;�F1�E	���-��n��޵7�詪�9R��<a���M���xߵˢ}�׵��@rB"��������"�Уa�$F�ԗ!׉�Օ[v��p3+��脌b���1k�5,Amv.�75ࡋ	B�ːm��[!��4а��c�?��n)�}`ܺ�2�m
�;�WHw���L'�	��w���F��YU󂰭�nP5��!��]�Opm���/.*ш�a�"�I��xU���7f6��o^5�e����C-j���`�(�;��6ơ,PZ�#b�Hޟ�X�7��ݚ3�Ppn�̧%��v����6��լ�W���#��B���h�'6p��Vk�,���k��eઙ���K\��jU��Cy�C\v�>�5��r�z�I�Vr{�]R���CGb�f�}����0S~8^��C�Akz����ü��=Y��S��b2�o�+:v� ���[�������Rz���dM�An��=�0B�֕yo[6��+U�u����P$�E��we|1����4Ӊ�"��Rw`�0�WXY@�T`�� šh!䉇�Iu@ͤ�3��ֱ%�ҬE�yj�w8�f�V��$ܺu8�N�E;�cE+��DC_���S�<ў
7���/�,��g�i�7������(�w��Z�V���Z�1\i�ގ���Ya�G Yw�8a�F�X�yMkW��%��/���T�;X1C�1]�3r?����7�/�����/�v䫚�����n^ѩ[Su�&tާX�CΨgT��ؠ�����@�=�f]J����J��uq&�oMm�v*���)t�ރt�i>����%-Jd�������p���q+��W
}�miЧ������+��)m�}����Y7m�.Z9*�9�y%�)E:��:�n�8�:�N�u� ��YS.��w��������NL#n��k��׽�:W�vȕ�J�>�y��u>�Y�7*���bD����@.a��}lY�urJ�-j�{��ۢj�2��d�#3T��.b˻Cr��dEg�г�<z��i�L���+���ɡ�>�R�Z�]y�he��D��g���s���pmM��(����xV�"^n��Z&k�tf���VC$]�އ��ܺd�M
���0XX�u9)�G�x5tj�� =�]3d�j�;J�6���ݳw�I��P);����5T�����b�P򋢘�#wBJ�F.2��
�) ��H�:�J���B��$h�Ŧi�$�m�����dR�$.'q���=t9}IJ>��;�W{��]'�ދ��o�]�S9E�H;��dO�B����C��ՑD?�
��(��AŁ��$��=8��5���mk^5�������___^�2V�!$PZЩR�P.�BU:�$*(�~P�X��8��$���$yǜ�q��ƾ5�kƵ��ooOOO���!$�2>G��j�
���T�ew�T'������ʡ���NOX��Ǧ�5�{kZ�k������o�������FQ�ߞ���E}q��K�b�2�Dr��(�p�BIs�x���ֵ�mkZ�Z������������HH��Y����X���UY��eDDUJ�(���2�2�#�h�gH

("	�P_��%�C�DAI�z��*�V��N^�L�U��I�,��5~�Î�w
HT+6�����M$ND�&((~�օUs�؁G"~�z�&@YĂ��\��3�#�?)�2�*�ŉI����� ��"�)�������}��S��M�bfq���H"(�B&��ԧ�-�m&�^e�)�)���l�s��X�$/mO���G���tx�dp,��Q�Nc8T��`YW�,��5���e�M0�&m"0�d�Y|q&	nH�e=��n݈�TK�CB�( �F6XjQ�#�4ɐ�'{���#_��Gq@1�q�\X�"��� <	 {�-�װ:�5)݇��mݗ?�O�iZ�e�l^�GM)����!�m2�<H8�D�:��3�Kg���[��/@׌nN�gԽm+�X
Nq�&�w�I�f�)�����|��71��,R�� #G�_�<@��!�����W����� JK(l1s�Z��5�z�Ɲ<�l��OA�#_�O$@	��>$>x�b��>�~��L]z�ׂ�pđS�Տ��ǀ��fֽp��`h�:���� �xf}08������?`���ΣQ{�y~q���Y]��L.� #�P\�zԎ'�� Փ��> XS{\�	���9	�5��~NV��l�s�[2�t����)����$
�A�$U(5��4�ٳ�Ő�ZC���;�n�t���ϲ�9 =��~�oL*��qMc�7�M"��<��eA-�1�9�s�V��zw��O�	ص�zX3p�м���\���TV@��Xp�@��ӷ��<}*�xSLE�*��h�͚��:f㠂�oKe-��qc@}J�c������Os�Wu� !�|��y��0�1xNMr� �l��L�dp���s~\a�a�:�e�'���`V@w:�n�7w�d��N�4�[���*K�w���g!�<G;���=�]�������sz���w�	Ƀ��@��6)�r�"�k/QT�){���Һ<��*���7�������mq�����9T�'`��[i.��;�^8����g�>|����P8���c�8���8〩��	��� � +��R���[S{�Py�_�Ⱦp(wB�����m'2pQ�0��5�`Ž��U�����9��M<���[������5���N��n ������qL}ڞ|5���}�;�z`86���1��P�n�u�s���\�a����i�*�7�K�-��ώ\�=��,�ou;xs;��7��.G���=�Ɩ����6�09���T���)>h�)�%%ԘWa�|�y�@��ь��k{��tu��u#�8Sc����[c`�����*`ct�jEs<k�o�BW?|�|��M�5�۶
�:j�l�Xt�Y�8m�ü/�SVϢ}nY��3!���wfn�*Kx&��=jl�w%O��;{g﷢�TQ	���憼��EǄ�r�Y�(�2d�Pd\3h#`<h�9�<FW�6]�s��)��L�XP��;Ƨ;��}=&�Z��O�B�H0)�<�_ޗ~�{C�sk��]�7�5d���=��)���f��ޜ��|�s�w|x�u����t�^0K�b��������z�8� �n�EW�;8lⷞ��5��y�\��񛍷�� �n�ٮl$�=H��B`�EF�a�4͞����Əe�~O���>��$16Qe���vn�{�G]�HJ@4f�����\��v�+��&�A�!��+d.,_�EA)����)]A�aȪ�f(�W\f����߷Sq��qD1� o������s��+�@{/�\�z�����?��+���Dʂ���҅끞�1�9�
�f��͘h��<�=������0�y��p%�}�$cF��\��ۧrG��� �]�f���S9�8s��؊�	/&�`/v�AJ�0�F���r�������o� �3p���;_�7r''c�%�x��	�(�p��72��v#d�dkC?<�;����}o>��rxM���9�>��Wn���d�ag�4	`9d��Q��#^�xz ͯ?`�����,��=�s	��L���6��u�K{���qN������j	tП��3�tĻ>��ֆQM�ګ��P��*�rS�ͳ�׿ń �|�H��F��rpx�0#|���x�N?����)�tٝ	�Y/�uN�+8P���L!���fv�	(ϙac��OJ+��H霴9��y���2�)52O�V�Ff֙�Imf@yq	�w��Ó�ȟ1j	��n��e��.���$��rpC���|؉�`y'���y'��o,:�)�3QK>���WJ��=Q�<��dvu�
���@N����W�y�8}Ru�e��h1��,fB5�&����{���|0�f���؝*�b5�#��b��ܙ	WN)nR�k(����Ֆ��xy��{�Bw7�]
�`|����_
��x�/�d����Lt��s�[X�v	C�����#����A8�	�8�c��G����ꬪ;������^���6�����ź�'7�n�9b�X$'����fƃ����)R�8�Tp��{i7��/�|��M�ߐ�LW�t89�hx�pZ�^�t8�9�Hl_�mg���sE�d Ql2_�q�Q;��| ]#ޮ�`��g�y��y��O��Z�#����^}���F�k���Cފ���	i�<Z�{�@u�,���b��|�.�v�z�A�M���S��q�	�-��p��Tx!��Hu���Y�p������\V�΢=��.5�-�l���*�w{
����:��	�#��l�{���v�H~���XB�y+C�O��t`�F��Wf�@z���F����� KzA�A�P�yW=�{���o^b�U�c�C�!���o5���b��w.�\�1ow���r����!�������S�w���U��l ^���Xwa�+�Sd��z�K}�{�%�]	��G�����/���|��,�>^�Ot�lowtsSTw,���2��*�검�bL$w����O!�cW�|Aqa���>k�ܟC�LR��pYh�mWX��f��E���#l'�X�����x8�y�F�U�7�����Ņ�`T���J�Q�GE��2_t�H���}oL��!Fba���=��u�u�;��-U�.�)V3M�Z����fN�M=�Ǣ�[�����ע��ܱ܁sڭ�;���^��&Q�9 !!e��$Ȫ6O'��Q#���#��*&F8㈮8ウEX$��88<�++ .)�U��y�wv�U���^��턅Qn[�~�W*>�SL|�zY;c�=�[xp��BG�gCo?����֋e��q@�Ǟ�s��ŵ���K�st��;Sφ��	al�Z@'��K�/�4���s���O.�{3<��1�-�	�Q��r7K���1/�n-^�m�k� �;\o�X�����~����`5�ndIz��H��||�p���+�|�4��_�|�HWs�M�jw���[���R�����a���y�Aס��������t�Z�H�������k����pA#gZ��A�z�cC�������h�!�:���/��ϖ�f\���j�}�a~$@[sn3��!
]��՝5������$φ/��)PH1�)�>�^�-�*�Ǐ�P� ���ֶD3r��Fu���'�o>f�0���5Qzd/��k�#��$a����>�H�Lz��U�m���hU�y���8Y`���������G�<��_��K!M�vW(k��qY�����J���Ԁ�ۖ�~q�oO�����Cd��^���J#��@&{N��l+�@RP!���ߛ7i�wo킒���HlD�Ȑ�gR�$�KE�:O����1]�m%�~Z/���B��W��������Z�b��ѻa���b�(_;�p�ˠ������t��μ���;���(�8A8��c�8(�D��v��Y��z�8�p}O0�޺�
�\U��V0�~c�z�  ԟ��$�ӛpu�y�O�u1�������1��=����g%�
�4�O+?h'��ܥ{���W���XC�8%N�_=Fnb��=4�Y#O�ۋ�����+)��N���U��KCE�����ޣy�7���YzӨZz/�WSy�os����V��#������
���+�\^ң�k��Hh̟{�M�rT�q�<��8d\����~�孡 *��
�$�����T�چ��ͭ�:�6w�iq�ũ33g�w8�R*�	�.K�qt5 �߷��#`k������_�Y�����9�Wٙ�+���y m�8Shmn�9�r�	Us͍T.��fG��;��,�.ý�;���S���+�ӧI�p��ù~w�P�6�ϒ��*A�i��5���H�o�*C���@T��MMS�k�yi�<Z�	n���� x���@t��6|@��1�����E�1���;�C��ZQ��֢��{�r�\a�pf��_�� �@`����Y���p+�yݙ���7�5��#̼S����B�8�d=7U�Tӂ7�q&���b�v�j�N\�a���orSU���38��/J>���Z�����ٚ�(��3�^R�,����x�M���y+�*���p��nh��//v�}�	 H����U��*�$8ァ�8�� o7��#qn�ͣ����7�3̾/�i� �H,��?�QA��b<������!���k�3>슥�Z՟�d�{����3^�fj�VIa��Br]���J�p��kW����K�-�:�K]�7��{W�'�y�L**-���eo���k�w/��;���T8@MCl-��]�q�	�u�ڸKk�=(EZ�Qo/�jZ�V@��T_�W��Foj�zKc +��|�0��Y��s=�$�P�Y�z>�#���(����I���N�v��PQ`|����P����ڱ��g��v�.$��Pa���}�U
�s{�z�˨U|��e���_���9�u����7�p�h�5�yXpi@-�d�w���R�y�k�T-U�2`�������!�H9B��SQ�z���&k�7��=�/�Cr~h��`�)0��l���g����
�p;��Ϗ"���C�j����0!���)��`7x	�Z��P=����x�:�7WwW0�9�,��\O�*y���
��Q�;��zXr�1���@��x��'ք�~a��]`��h	o�܃Pwr�;r�e��t1Q�F��,{���=^4�mױ���E�2�hE�,:Ed�v����3��ƀ
s���J4��]����gI��tY��z�/ee�1iš�p�սܜ-8�F����U��#Σ�}�"�=�3��ǫ��FA�
8ォ�8� 8)Y@%��~y����Ϡz��l�Hw��Ĩ�|�KC\8�����xk���
��t^��=pt��.ֵ#+��Gw���U�Z���!{�azA�g>��J ������-s�!XgQ7�C궈�.��{���c�8�i0�)<�o1�L��r�K�:�&��NC��GIi�mi�s`LKo��NSѹQ�����x�����{Г�=����e�a����˄��k&UmYi���5y��y3k�;3��Ȧ5FH ؘN��F:N�ok����Q��;9=����R�9�p��������ϛ'�2�&����O��A]nV�x�pZOS�8���ó�j���VFrx?�B9R��q��pN�����'{�����d�g��]��7������qq�q���S��X�oLk��əj{2q
���]Z��2������@{�/3{����2����>מ]��P��9�Ϙ�X�˺9�ܑ�ϙ�R����Q���'��d�6���thiz)�j	���;oX�Τ�a��z�����~�vO��MN�q��o�Yj��~=��w����X`���YY{ݾ9�ӫ\����)� �:`�(*�g�0�)��GP�x��&�쳯3_o[/l9���c�������X�5E|7/����V��*tpJ�U�$V��mF�R0a�(5
m�E6
��H*UQ�ps��#�����09X�*8�*8� �G8�!f'ҟm�U���7��	N2P3�9RO_jG.U�WuB��F��q��f'rb�e���S�W��*����4u��]9&�����g	����O^f�"Xt���rz�d>��1�a�Y'��i��~���m�jU���]X�z뭧�q�����9�=���
�a�6��ɉ|�$����8	�v�2F<�_t#{���b� 䉢� ��5�s �W��-�#�>�_ut�yC_l1e�5�fq5Zj
"����Smf��K���m���>��E������v�S���߼L��5�/��p�����_����{��ڞF�������!幐`�{��<poUVnUv��A񎭉l����fA7[�>���ɀ��Q��C��;߮홉���y|H�nO�r�D�����	����'9�^��*��f]��r�T0�hسy؍e苦g��p��i"y�M����Q��5��L�fR+��Xf��r}�D	�PS:۽��K;G�o�3{T%�z�}�d�
�=����T6�k��˃ ���vr��������p�����:��c�s��/�oL���Do<�q[�V�U��8�
��tfus���r��pq|������_����"�D�)���tSə\������^��w��bXxViOd�wV�6�k��l�'�q�	+�|fo�:q���!�{���~� �Qq� c��x{ކ {�\�"���7> �����;NuB�C��59����=��&�u��������.���5'Qà��>��+R���2�H�$1���g�d'�A��o�5�Ν5�S�g�g0�9>�ٯ}�Gy����;>�����oЙ��|���-=jD�A�РKȣm2�+��Uv��Ƀ�&��?��)���z����J���6��m����] ��t8�+oΎ�|���^��TG��޷\��|��X�5V�,�X��B��S�����}�9��AQ6����)�h]|�i���Y� �P����4g;�N�*����k�����^�ۓ{��"q �TBH�/���:D?n��Ci�PR�����5"���>�E@���'%T��j�oz����5ΰbT:����؍�1���`�y"}��{�sB����B�����޸�K��W�̃}�>�b5�h�����wB�b��w�xa�����\(֮��Ib�~D�'+��g~c��>��B>VИ��Z�LSqtz4x�'���ֽ;���z@�ǵ�+�M*�7+��ꅽut^�ALj��e��rQ�ˀ�!������w��Qo=xxklR�`�3�U��tkR��y���P��I�M��]��ҳC�"��ƃ���𶍻�@��3��͵�AAdd�]�	�����w.X�d����9�K��2Ⱦ�)f@ay�[�o�e��Į�SPX��6�'9��]�W_pL��Y�/Hȴ�����X�݃M�{��4\��V��=A�p�r>x�[
��W� � ��g�uG��Po\V�.":�F��*��P�N���
l ��֮F#�_p��U�����]o1�&�Z�7Ns���/��
CM�\x���\����t.d(��C���<����v'f;P�HٶVɳ#�:ӬQs|�`]v�3s*�n3X'+'��<^_T�9�	�@�׮�N��#:k��qW���:p]q��V���&@�X�ۮl:�-��#	�3,j ������=6!�彼�YnizZ>7�Ĺeõw�"�
�C��*I=z�/�F"���'�S���q�oT���u�S뭃(P�����Ɗ"YM�:r冫����|�=*g)ռ��o+Gu!:
3A	����X�tF�{ޥu���-�e���V)�I�KN��7���BDaZ���3jYO��KWڰB��`g�!R��{B�7��l�n>4�ќЗ��4�O�gˋ=��p���1cݩ��r���R�{9m��Tt,S'P�Bl�x����mYx���;1�nNA�!��i�i�>V���1ݷ�OU<:YD���u���v���.�Y�`	҂�u쩷\֩)E�Sf%����x�q��`�J�� ��5Y�Y��TkB{���2_1vF�*p��AqŢ5~H�^w.�]JfgZ^��K(��/���:���p�ˆk�\.�tjȍǸpC���_f�ItU���gi��VTIۡu�dQd��YD�����jn�.�[�d�kY�.�+���Nu/�KwV6�!���Ľ<b�ku^�C/�tj޽�u��������u���&+̖h����;b�.dw�;�r�+��{:᩵�\���%վgn�y�9y�s��]`b�ω jS>:m��lQ��t_�V���Y,묋`��JE�-Sg:�b��Sk0X�a�ƷkA�	�ň�.����[�ӷ����^k+��	��cgu^�듖sao` epg�*]ۙ�jϹ����w	>����K20F�4�U
�ԞS�Iеt�i�wt.peL�����2^$wB��	H��N�2�[E�C��9$���g1���z}}|}zkZ�ק׷������Ɖ&ÒI�9��+D �U��Eȟ���A�qǷ^��|k�Zָֽ>�[�|�7�������T�r�"�(��"��U�&E\����9�$	=c��Zֵ�k\k^�^�ޞ�___,��q'=�S"�2~k((+�f�ц� (��,���ַo����w�k�Zָֽ>���=>���XHQp��Uʪ�*+�ʫ�7_�
�\.s3�S!�)]�?_�9Uʠ�5�Q\���*?��;�(�"#�$vAL�E�ÇL����<6r���EQDI�*�W*
�݉A3�v��Op�"@�6�Dr0�Tg#3��]�^aA�˔_��3D�(�������#��Ȋ �����܉L�9�	��:�6�ta��:uC}o-�5`����m,�S����6�k���x]N�^+C~xo��ޏ � ��*8� 9�Q$	$Q"�@d>_=��w�x��K���g[;�<�hnm�����"3j��8o�i�-47.}�}��ɢ}{�Nú�3fi�!����o'���gk~p/0��@-��K�~�R�co����,(,2[�.��v��K���̮�ű��/���G#I�2qt��?���O�,ȥ^xoj��]R�Ru�_SU�t�;��q�S�t���y��b����h/��xt|��/>"~��/�>��S�{��w9�m����n�R2�}�N��3u��y@��;��P>���G�]�l�_6t�yB�Mf��"O|�fI��k�>qcv(��e��z�#
j3��c˻���yɰK���_�x�Y���yy��q>}�V{��BB�t\Piz��5�X"��.Nٯ�;�Ү�L���7�xyC���r��*��Vlc�E:׆����~�EZ3�桹��5���;�=˥��~���
�Y"|D�וu~X"|\K�T�f}�xlקذ5�����쭵�{Cp�R7�p�3gM�Mms��~Yv>~(��
�Y��}G�A��L����)�cU<*���c�H�rP��\��/U#��������tq<?Y��I��,���� F9�2�U̅��`�}ӪH'���+��3�V9�����ά��1q�\�ww񉾧z��_�qE���≐	�8�@�8��8�*A���7���ޱ������S�#X�XĬU������/j���w�y�7�C]hHO��&��k3������ڽz#[u�?j�@W�q|y��fZ�VW�R��Un^A+�j��������c�B�4Bq+��ꛎWn..j`_��\/�o��c�o?b�����T��Map�^<:a-�{�ۏi���(\b�f>�^��zS�S�<���N�1M�oD��YN�t�^��[|7�9>{��0����{<�|!" s�	�jV2y8�PK�Y�2��T���NM_GAF���n**�O�&]�ް��_6�B�A��E��Ǥt����xd�]�Y9\u�n��F^���J}�Xԫ�cg<�.�
�}#k��e(�Z:�kw�"��q�Z[Ǧ����wL�{��gܸ]����
-�͵��?(���kd�m5?�7���>�3��(��)��X�B��ާߗ�>��z�X��_�P��^��l�jx�̨���T��i{�<3'��3\z�ҽ�\O�� ,�kؖ��F8����|�W4� 6�������dغ����}?|�#�2�E|��:��8�efkt��1[�N���#J�j(ԏ��UDSˎ�xOf���ꕩ�m��޾{"]�)�r�rP_jh�0i)�J�n��΍$s:W����` �g	�\i(�)�f>��ۚrny���~H��qQȱ�1�Q1�Up`�Ȫ{���vx��d�گu���f&B�3h�h��Tc�E�$�݊F�\���ޅ�k�O�Qڄs�~W�Ր�D;P̄g�k1��-K��Tq�-Gm�m�9�>x%����p�4<�K�D�4�M��Kս+�H�	�=S2j�Rw���W	��4���
�$:�^�.���*0Ai�={��4
��2q>��Tu�R/��?}6�����}<�Ŏ�����ZKh>����l���z[a���}L�b��Z+"���"����+�<�ۂZ�z:IN02��)�}���<nd�R����p�3`@8�D�p�los���>�/���	��.�W����n���W'�lH1؍[]E9�^ښ��%�a���2�9 �P�j��Y�ؒ�N'��U��Mg
k�f�Mm~���a�x 0�	
����R:8~����Q�}��#�	�;�����RE"Jh6�RK�� �X�c"��aI�l���O^}�9{�8�=ЁS����U����։�u�y�c�;Y۫xY~
�G�m��=y(��BX� ��%�mf�H&��[ Vc������G�1՛���~♅���J�f����D�drMvM��T-lL�ܺ�y�`��ɮܷxx�O��Q�`�` ����_(����l��j37x���a�?iO�������I� ��M*y�uJ����}�z����8���c�8�8c�8*��H0 �W���i-˳ݻ�!��wƔ�%zi��V�L��б͛���uE��	8�g>d��u�F���EDު��L���^t��G���L	b�	���<�,0y�uϡUH�����:a��Z�)`�g�.9;x7N�0/�S�/��EӒ�|WOvReC;��ۖ��گ_����G������fOt���k��
�+�������6[��h!]:z�$�i�]�;������fs�J��,�J60|���swl�m��˲�p��ƲCzGt�<�2m�P�-c^��ƶ�;Ǹ8��nZ:\��3V�c��:HV&��5�iU��7�K�K"��#М^���}���f-�=>���K�����ʂ���[Rsvvp�B5�y�+��-��ʉd�\=V�3I�d��i�{m���]L�;���v���Z��p��~�t5熹a��f*"���m���a�c�g+�+���#_�b����F�v��8�Gp�r�)U�E��]|�I�V~3���1�56�}=m�9ѳ�3���Q��%��m?y���g�,F�j��iǳ�!�=��)�ol���oē�I'
< � l�<
cc��q��ك�7;����R�q�$�Ū7|���9Y�;��a�������A���w�~yL~�N8���8�,�8�c�8�P����}}�]�Aظ�ۥLy���a~��NN1�����y��ra���.�z������.��[^\��^a��������S�����<�uGOs������G���h�7�H{h��q������p��&�j;��}k4`'P��!� �2�4g���V��Ps]���[�7�v���b����0���f�r��,�:x�U�+ԛ=a�=%�s�q�}ڞC�h#V_{��zG��sQ�wf��+�c�倍-��֘rڔ9s�&j9c����zc_B%������j6p��v��;�,Q!�!>��Ǻ��Gܖө�=��N��2y5M,��Y}O�<��ﲾ#���H5RG�������B���퉼��,~�;��|��݊��=�Cfe�\O\��Wd��;�'��~#~�z`�e{��]^'ᫌ���T/aN�5v�v���[�Sl1�{�|	Nf��q�*]	�=ꂐ��0oP��*���m�9�������Dqa�s˶�'�)�9��������gx�'�G�hp��g��;fvg�4t������S�3f+ٺ��8�B>]s���9���g�]��@9�z���UW�P]�h�&���![bs�Kkq��t��"�)��31��^�'����k
.L���������u z{���Lq�Lq� Lq�0F�úx��9;�� �:�)�E����<R�e�ú��1�fy��}�ST華�.�W�Ӵ;��_��Zk`3g�/��	���G�'%Z�t��Kڙ���	��1�W�x��`�S�;H�ww2�����{9�mt��mA�
�L���g��^�p6\A���ݘ��tЬQ|�	:k��_B>��D��Y��'�1P�#}0�'��xt~_�'�~J����N̑r�@l���$�R���0D8���HM����5�����7�����4l�5��m91mŮ�v��9�Wx�q���gf� �o�D:�εt����>j�٬z������R,�.��Vޜ�37~������$cƺ��m�~��������r,�˻��;h����{�gjL�R�鳒R�y��N89Ɍz���"!0�v��;`)���yO��EҬ3yq)�Fwb�VMg[]f�I͹f`����-�s���&:G6��.@��OK����g>���/�O�ŻwBe\g��W �X�:�	ass�!e��>��	�}�?\)�.���Y�����>����v�F�u�bq�łHn�!��)r���2���y��әH��Nã7,�09K�!K���H�l�bxm�g�p>�Hf�Vr�N��WϺټ��)�,�7p��o��y��u���,pѳ���8�-A	����G����*�!_� �GpA�s� G�������6�=����ȭ��ߞ˝d.��,Z-������C���1 �O���0v��A�����ට�x���Ѭ��*��bl�q��5{�{��O]�d��oѓ�'۪{��=�=ϔ�o�df�0��p�>n���t�sg����'���ȯ�e�\���������z1�%^�XKh�XPu������>@��~>�Q#�@���sJ�"?,�(\��˵��;�Ǳ�����wp���6u��Y�r���0m���H�}�_����V~��$ϵ���2ƿ5l�ѻh��ٮ�C}��G�ǖx��o�:�O��, ��� ����%�ޒ�ll���k�WY�w�'d����090�R�+S�כL�b�>X}0����g���0_.�۵W�eq��>�S�M�2g׾�CH�tG���<�-��s��*��)'�6sS�}j��{��ٻ���q8c@mOދ�L�����c'܃��rPb�f%=��
�c�6qN��r��+(Wd;��O���,,8E������>�}�V�
t@;	���D��n��C	uT&��m۞K��e�eP���8�2��ո���Okt� )�T|;�����&��b��k�J��?U˭s+i�������\�	����KV�k���/FMW}�&�y�T�eK$�v�\ܿ:�ަ}��V=?n"�8	�8�8ォ�DIz�<��������/ط�XkWp��U�X�!�_!X\zD��>���9�xK�h�d��=q�=E���]�<��ܐr�-ߍz=v
�:`;�`@z�XA�D�uR���R4�gV��0X7����\��	��c<��|�W���+�����]���I�8XChF#I3�5|V���<cԺjmb\����7H-ڞ�+�@"&i��ˁl�>w$�&v�x��{�I	���0�;����x[~�r/\��n������1�&w{ۺ�-�����zy\�Uv�E��,��1w�
��͇���g��m��,}d�s�إG�U�vO��5�S�@߼9�]��{��'	�	O�0WO��oH3WH ������D]9/ӂ�g�3����Y�U7[]�y�����E��]� ��Q��W�|�E&E���<~����_=��J�e��闇d�ޢJ�|�+l�a�� v�uo���vĨ}�':�)=��Q�h��
i�1�[���D�{ӓr���W��h�����jSՃu�Z��ȑ��ꢶs%��S�\��Y-���Wܷ?nPZ��R4��Wj�EQ�Bo���~���Fk3�;����Z�w�����_=�T=��ͅ��Ȟo;CgE����H�G+���2c��y�;�]g�9����ｻ���Ȭz1�T�qSq����"�;�|��,�7�LRz�֜�G���q�+�+������'xAXg�����Ӱ-�d��:{[Lpf���Ä&����\�K���\[S$��Y0ޘA�#!�}5h.���\q*:vx��\g���Y��\k1Q�v�}�MXx�3T����C}x{z�
D�p,oL����yӜ6����`�>1rß)�Zz�=��;�s��C���7�A�JNPy�rì?���]��ĨUߥRaL��9��;�O��x�8>��(G�$;��i/EB��Y�����	�c~}��(��±��9�_8Ɇ]��h�3��msx�<H[p�gi�+;q�C��%��i`_��W5�m�[��2+=��*[�|��Vr�y�Fy����ä!��_�w5���<�*��a#����b��9Z���9/-۾��������^B�m8�0�!u'n�OfD�>��Ȁ��TX,��A遯�~��{����*���1�ɀ'�ϕ��*���9�O�_�k/b!��yăƭN$;�21��z��L#�E�q���~\xѭ�����:������M�7zH���Ż�sOA��:�钎妒������W���#�b�H;�2$�AH$�}��^��B�m2���V��՚��?��5��锎�'e�����}�S2���k���4��6fss�e�
		#���8��8	�8� � oz�f�¸�5���e2��Xo�Ξ�	*R��P�i��B>�ǯ�*F7��P�2o��"s�Z�m<�)Ď[+������'ƾ�,'���Q{<���xP�)oߵ^pҤ˗��l3�j�vg�g�xS�-��	��H��}�N��Fo��Z|�ɤ2�����C�����p�ܼ����DV:نk/"��)Ja F����6y�{:�G�a�*�239vI�Ο�˼!�86rE�Dc���鐙��S�M�7W~Õi�n��h�3{��[{��:!�O3ő2���:�(|:놫�� �}�x�)^+jǶ�Z��t�t�m��Y]ʍ��.8�{\cD��{�����ή��ʰ��G�~�3&��\BO��e%�5]q)++xx���Af���W �82��7T3�����3�qmB�Bi�c�u�t�eWv��:�r~�>����!P:�H�DbT+�;�< ���n}oV��o��'FjM�{���-7��� ܜKt��ǣ�5��@�;�Z=Dש���&�;��ߣg1�{�`��ʝ):�*�;&+6�7i������:�N��p�άWJ�e\���o%[�16�5�c����Zq�xU��5�cN&��Ԋ!Bkś�YVM���i�s����棳C�q82,���*M�nnT̡A��4U;g(#N�Q]I�e���Q�}�0�4m6P�y��T/�ֲ<H]�&��&(�#�vhT���b�5��Y���s>F�t\�Zb�cmJ첮�L�yC���T����˦��8�u.g;��CU�9΃�w:ӮO�*�I ��N���\!��_�QV�A��sy���e�g����.]�tkn:�H��\%���۹g�ܻ�������XӴ�s^e�8���\�GPtu�W,֕^���a�o&5؆Ћ��w�%�a��g=�S���K���Ԝ3xv��|i�oL�3���X������DE�?'؇wD�5� Y2��Q�8u�𬴂���(n.��^�B��zlїe�:�V�M��<�*�s�ľėp�1N:љwF��K���+:��hU��$�=��Q*>I�tkZf_�w�,(-l.��9g���Fe9�y6�/%�|�{�n��AG[�^����i���ۇe9���p����kZ�ai�F�-Jt��=3Q�h����fe��J��n��Id>�r� +���J����A`��u:�}�!�{�$+�nP�L'Z\(j���W	v�	hв�l�RGR�Z�kf����EuM{t������呺TC�u��s�&0�-=X٪�<�Z[�V�Q��k�]�bÒ*�;$�Z�:�(gnPR����.���l��h���a&���A�z�bz�Q�Fd�AɌ�K)��N�$WNս����&�F�p�=2�{`�I�ۇ7����i�lv����s����WG����Y��
��7m�F�8� {e��b����+\m��K�q۾����L�*�rۘӖ�w�ɒv_aTf�V�V�[���)�d�lu`��������\��V�8%�Y�[����()�$�v4�!���=\�Zb�mo�*<��*��sg,��
T�d��S-δ�De7�I��zt;;R�3��D�ؔ�s��z��}J�"E=2V�}�]'*S(:2�l�;v�ƈktIc��╹���x�V�y�� �:���0aV����\��/ni	�e�����Z�=��,���֝c�\�{�r�jۼ���mAN���g�+L����jއ#��U�V#�zL��1B�/� ���f��e�2��S)J�%��M<U7%Pԫ���`�!w�a�m�Jk��J�ֳR�	�zqM�puQGe�.�u��f�UR�Vƕ�E��c{6���Su�X����S=���䯞�k�Y�{f�.����˵� ��tSS��+M,��BUY41l��[���A��>��lE���7;���6�%(�`�L�J�1ѐ(�`�D���ĚP'a��p��}�^bꄆ�["�N6d��XE�#p"�"Ld��Q�PU�f� (P6҄F��P�$I4(IFH�aΤC�&QD��	�{��~�y��(� �L��NdQuB�=��\�1bw�r9O�(�H��n߻���7���ֵ�q�zz~�ޞ�___��Ns��h��fs��d�Ȫ)z��;�D�PC���Zݾo���߭k�kZ�Z����������ԑ$AE���Ȼ�l�C|�ʪo0�{�Yst�!�8B<c�k�_�Zֵֽ=>���>���RBB���d뜓!*�������R&���Z{�'OOzk^�ֵֺ�u�OOO�oO���z0䳄���$!$$��G�Qr̮�C��PZ!p�TJ������®Pz�d�D���r�*��������j� ��UD�Ps�G&QաEDW+�đ�7�{��Q;�r*��Μ��DQTO�q�?N��D��T�9܏�"��;���9U�̖U.E+������dܐ�E�*�()��I���
'�������F٠SrN \L���f�$���iv�Ǎ	%�l8	b}��eάw�famem�5R��-n}�Z4�����e(�]s7�&��>H��N�n�Wz��>g��S�u�څ(!�8�\$�`�h�)�
(T�Z�D/��KE���x�8&8�A#�8�8�9���sڅc�߾��A	 ��Q$Ϻc^8�W�Pyer{�xQ�V8�Ty�G'#^�b��-kk���p�o-&Vm�t��ؽqA��9��ǌw�'ײ�7[�u��yO�*�y}���ڄ�k���eƻUZ�J׆��A���!��Z���΂H�����N�N����7����O�q�?x�g`��gr��	�{��9nc���A���~p��v�X)�ު��|aƜ��מ��k\�"�%�e�dkt�M��r;`&�cӼ�`7�"ptS���e=<����Gx�����O�[��7�dl�t�s��^^�w�~�T��x6ŵ����(����ҳ��@7x�'ѥ���qP��Z������ΧxG��x�D�cޮIh�I9>�ٻ�KN�p�z2v3��_���Ӛ�W�ec$�����`�|�/`����v��*ئ�ov�,bF�i�Z���������nq�����$lu4�"�/�������Ň�����LyޣMV%ZkI��8f���[����%�V̰�]�����_��0�~�z�%B.v�WĬ̪���&�l��K@ųy�'�
/�+s�^���rC)�����:|>����M�;�Jq�)������n��e�J�q��
˅���,p�	Y�&�/��7��E���駰\�"�}�~O�� �8��&,8㊘x{�Ҹ�����~>��[��L*s�Tr׵
D_U|�T���(S��
�F��3�uf�W��?E'W;��W�����쑾��	���	�7 ��뀋�W3����җ���3�>k�!� ��jz��L���7+��/0�*�Ά�Q<�(�ֈ�v�E����ȫ�&Μ�q�[ռs׭ٸa�X�_��ò�8����"����?q�I���k�5�ŷ�%P��8��^�ӛa�>���)���8C�k���B�+�t���k��9��8E�G(o^�>��uc����_�WW5���φ���\涩�0�7l$��wEu��d�0UOU����v���b'��6��A�ns���^=���dWW��_����w���ac�G��m5����j�1-�f#��KG}��E�d�'�}=�����zFׂ٦�`@��g�r�fL�����1�ø9h/��;�-x/�-L��EGd�p������;���㥪�c��t�]��/g���_�v�O���y���k:kT��Z�N�E1�3�w݅�8W����ƪ���jb�F�Me�2Z �A�6j3���s��Ⓤ����Z�W9�gW=4oq:7��1'�f��+x��X��!zB�uh\�m�<|�Xk���j>])�w*=�|�qo^�b{z���h��
���Z��D?�~�q�1�b�@}�|�m���2��J�F-�F;t��C�wf���/���P���XlLǥ.ٳ}�%���?���P�^t���h@3�pH��?~\f����*�G��M������aۡ��������6İ�D���B ��=�����D��COEq��W���*���q<��2U��0�i򃺉��}�7ϴ: 4�B��b]���Qޝ�}oa�{F.��b�z�NWZD���cϦ��6_)g�[�|I���I���xpc��Z�@�thU�1UA+v뫗�"g��gP�H�l��'�F�zm��'>ja��b�4n��i޺�ԍm���+fۨ�^F�I���,/�HݨE�s��rY��zl��<^L�d�*��T{h����׸	���t���P�㦶��W3���	��	�s���Ϡ�TL�j�:|���W���Ʊ�G}b�
Ul��-������&���<�����~���Q�� z{����V���N0S�j�۽�1\��H �=�-�-�͛mc���^q�2&�໬i�%&�he��!��~}�}vfܾ9+}�VY� Y[�W����&�/7=Xo�=�������G�	ISB�ޘԮ6�q֦�Z��_l�ã�n,���M��U�m]���ݔ���,��oΤ�O_�ہ�8��9��8�������yV��*�_����H�A�	r���P�s sͰr�2+�{�Hmz�1<Ɍ��6�k�t^0�a�0 �5�}!������lӜ��>w����|�4)��m7-J,��Xu�C0��
]9W_�w+[`�@�Ǉ�x:���Y���?��]s �o�r��ґ�E�P��k#d�{����T[.�ΟT0���bV���,d���⨧��'�1���9j����N��2����E�v���]t�<���I��8[
q�Ϧ�!t��IlA=>:3�:=o����UY=�!���m�6.O����&WX��p�I�\�K��Y'�R�0uf�8Q����p���U��%������!�zy�y�٘,9���Ȓ�(��~zt��L��UK���z�|�5w�Pab%��΅�� Q��،���M��x�޹�D�7�̝�$},9�>���޽����{�SU���s��>���jyY�����_�M�E�n�I��o�,��n�5����}���&~�	��X���_�V��3)C���x�s�����]ʷ[eq��x�����}[����~	����	��]M�bU���U�)��x�RɁX��4VG LU��b
�����!��D�S(���֫��8��9c�l�`��e��dW�r���G���z�U��g�T��@�-��v0JRK��%�-� ���a�9���?n8��H�	�8�G�����<�KqV�"��3{���=ǯ*U�w4���x�s�*D�9��*iO���C�|d\m�j��T���x��7��9��4�.��Y�>ʸ�˞y{}�n�����1(x"6��Y��Z���= ��yYa{1������~�3}E�g�r$��r��,�t8��8�G�+���$�c�ɡQ�)+��ݾz���#v!�Qp�w����nb�s��{�Lx#��Z �zѭ>��N�Aāwu��qڵ���:z����o�j�/�RL�(yw���7Px�CC�0����%�0�[J�i�D�+`/�v�o�þlZ�,���Q�c�p�G�c}�!���^&�6���m\No=�ïjKu�ؗ���#�=+\���.�MÞ���q�9�{��ۭ�h���OS�{ڶ8Y��cy��E��L��C�#�L����h�c,D���6{�Q��Z�]�5�cp���l`��@��Q�T��$wP�&�� �PQn�� k��D)�{�	�d��)�[��0?�?s��y|3�2%���n��?'I��κ�B���w�ۮL�WN�tܪZZ�h|Q8e����w(���`�ۺ$�ً���imyGpr	��q�@�B	U�����V�B�]��;����ʹ���S��ݑMԵ� �R2��s�7¶�l�9�s�ڰ?�z��ۃ�8��c�.8ぁ 뾹�O��a(�`B��;6�5óF0��)���(��e'�_�l�L#wY{u�;�3'��º�O���E�㮠38"�;�(�����`�/��ܷ�]y1��n��y�{֧R�w]�7{X5�r���Ά4��.�I��<�Py��w�Ϗ{O��.� ��H�9W�����h��=�8yBT���A�����'�G�����ױ���!��EҪ'��j����2]�T�z���'��f���]���Y�
��R{������O,�Hò]�{oL����B��Uˋ�ۏ��Fﾛ����`�RYAΙ�s��b�"+�w��7R�]\)��?Y��"_�]��P;|�]�J�|}�@�'r����H��m�'I�{+@aZ��"ڛ�ѯv���C[�b%�ɺgA'�����1�0�;��[NvH��ɺ&k���Z�e8���B��=ŇM��+K�pP��]����ǟ@��mLd��	EEM\vq�-�ޙs�$�7�@7G�����A�r.��h	᭜Gt��#kW7I���^�n�z�p��)WD<�̹�6����'�b�*.�Z�6*��u�*�,����m*���6��I�+q�b�wcr����ܢ���gMĂ��w��׶�ą`��X�LT��ڛ]�����p�sq�q�:�{�u�������y>�ɨ<�}�y=�>��,1�
���8M��;���X%����MTW��K�p�2��{7N>�t! Ϣ81���	�Ǟ��$���ĵ��i��6��3��z�Lf�He�}���7<1��@�� �8m�;+14���{�t�'U�"������b}����w�6��Pe%��(��c�B�cW������}N�Zln�_�t�^5�윮U�*���Q;���\w��=*�p5R2�- �9��r0`�H��l��ߚ�t��`+�P�K*	;�{Oc���U��W�߾~�|מ�;k�`��hA��ZD>7�hXg��T���k}�2@�Ӿ��_e�N( v�TZ|��iOA�43�r��ic��R�*��#P��"K� �"Hlx��H��� R{J����
}+ �g���O�~ 򕷙�_g#d38g��Ђ���MGOC��g����55��M犯��$D�=_^g3���l�Yh�Zw��~���ț����

Ǥ��\2XR�Ә�[䂝�ޡ�1Ac�Cy,��+��?��_���L��;Z�b�swE��i�s�4�i�^e��pִ����0ws�}w;v�{�l5�n'��A#� !��(,T%u�{�Ba�&��X�|��H�xⓇ,��DC��AQo�����샞ǚE�Vù�9O�k��8�8�Ǐa���=�߮�5��3�Rm��6m��Ξ|^��X�\,a}򁪵D+C��\ͺ�pl�f��T��G[my�98�Yw�U����ˎ��u�k�?��2��Q=R`ʉ)�Z7�$��nw���e&�zC��ghjb�@n��5hХ
S	mG$j �\=5��t��7�1�/=�}]�0���}0S͸B@��s�-��}��W��C�:{�]��3y�����Go�9����Ǉ�3&�{qGk{��/����/������?G1`�a����0����M]#_I�����e��~���u�W��#��|kH��C��V�2�{\��&-�\��}�u�yy�t�5��5�L}_l�� u0q�����k��ƾ=��<IA6�s�%fw�*���5l�x��-{PK�t&[�.gwr�m0q��ͭ��П��ڭéJwos��^�@����a�=�N����gO˭R�
��*x��\�̬�������	���Y������	=�K�v�:7ޢɀ�I�iՕ�e)�6��%b��n���Ѿ{:�93o-���z^���t�:M���[O0�E�O��+�#ۡZ��Ө3� G�%�5��t���m詵���)#ܵ�ƹGk_1[ݨLj��6�q�ڭ�o���@�f<�\�ռ�=�]M�-P$�P�Ji�� ���u���q�1��qN�|�>��}ws���v�y�e�7�dw�\W��ϸ�叟�9"OG\GǼ/��6Z����?�*�p|�dh�a�ޠ��2iXi�P1��_R���2|��	e h2�2�0�� ��2��ѽ��[v^'cs�'s3�^\�4�qs�)��^F(��#��o�	�O��,����b7�=<���*���5"��'���5�P�� >���S=����åD��g E�k��}����(k1?w���؅���j��P��pܛ��9�U�n�����R�_c���;H�}�(_�MI�Ƞ��mWn����%�"��M5�>��Q�@�2s�/L�y���~O,��u��^��VWZ�Y��	n���u.W�s�`$�8����A㷻��)eCR5��uHKV��!���fq��ى��˥4y�K�!����}\�7\ *g��ӻ*�W���3Tϒ�R�L��+װ��|���`�7r$��Y���z�U�򂕤�Cؑ��21�u�4MG�? �K:��܌[�^���S~E2�;��/�c-�=��=q8���#��G���t5{�x*֘��&�5o\7ݑ�O&%���Bٲ1�y���J�ղ��3�E����s�����_Pn��V1��9Q���$�b+٣�2b����v�k���`�N�u6����dn.q�6�]���Y�J��i����.���]�fCǳxL���1�q�q�L�}�}}{{���i��0��S^F�1M�8�έx�.�v~.Z��}&O�@��{$�nv��7�e���Bv��
Z�(�Γ�9c���t9c�%���`F��wQN�X��;���Y�����D����0֛JEQ=F^�F�MwP%�pY4��թƨ,6���d]�}pzG�������2�-ϐaCw�s���ǯ�xKL9����a;Wº���$��=C��i�D��uC�A������e�%xz����;kW���i�r$aa����h�r�ס��>˷>Ϯ5�g7���jB�y�޿{oz_$�Y[�u_�bap��>����[��0i��{�P���pl`�_8�7�c8,v��Vdq]���kX7N��1�wKM�%��H��G*j����>x_8�;���뺵7�ݤ��;K7��i����2#r9�w��#þd��fr_���Ui��yH�w���0`.��o�����-;����s�q��Ֆ=�`��А�#ƽﰒ|l$ �/W�E���b�b�	R�t�N���q���J���x��vqոXP9��P;]y`�\Z��6|}��w�����Uvʧ�^���v�����!���˺��:�A�>��]LJJ�H��^��u�ݛuk��3���[��wTw��e6�A%��r)j={]��Rۛ-f!N���eꝎ_1�Q�Ɏ�[L(����ǖʉ�1_N
��⥃�;]ڱ�0��r��9�x8ܖh�V4e��y��%sT�[�k�!^���3�@Z���"k[�����@qC���	R���9�A*��&���b���/�)��b���ސ���1j;ٕ�m�v�9�ڸb��6{U=[���V�2�^��u�I�n7�h)�+dL�&uѱ�mv���s�v��FE�}v���v]�X+ͮwl���]ok�w��O���]�:�:,\U�"�,L�����rW-]���<Ƴ�}�l����,9nT�"�̢)�t���Uy��:��5	Tcw.�*�l����.Z�*�+�3b�Ӳb�yЌ�=�n�{��c��.��R��'q)U��hG�hm���Us<<�p���K�S�*]+|�J�s�ݺ|��Wn�v3����I��:�r�T�#Bj�Z�,�1G=EA_D�
�1�Y;�l�T�>�r�íbl�(���U���mM��*��!lA�Ҭ�@��M{s��+��wn�gw}�1׎�	��-����w�=K͕}J�^�,��ս�Kt�6nX|6��a-箧>�Ɖ�)��zH�g��N�1.��̄���֪
\Y���r�5S(�b�V��v(d�Ѯ�c/����_kf�RT[����A(\H���S�8��|kr	gT�j����9��ν�Z��r��B����+��]õ�e�'.C����*�w��^��&$$�����P��)j/�ugRse��N��5yd�����)ى�Z��d4wH�,ѹ���u��#�H|~�*����4�E�â3������d�b�s�7��>�J����E{�C:�=]���N����|Oq[�M�؉���<,=Q2�G��!Ti�in�.��f��kH�,�A��%�+Z�z�"�u(+�[t�%�l�5��Gf���2�����/vS�3i+��)G��6�7�L�5+c'�����@+gs7�p�'P�$��5�e靷�X��2��}19��ר���=�&:��8n2�!��Y�Y�%����*�ݦ�J�M�ձ���B�9��7�:��Mj�ݱ>����mk�ъ�l��������A��<��)�����\�I�糭��v���o�o��q�kZ�^���^ޟ__�Bs��Y2�s��J�B��s��!��$�E�p篮8��_�o�k�kZ�Z����������$��	U�P^�����FQ�#�H���q�׶���q�kZק����׷����'		,��rB�U9DTJ��K��I''9�I5׎:��׶��5�kZ����������y$XI$$��+��W((�'�eQޡ���*L��b%U�;#����r"��
(�+օD~t*.QҢ��""u"|t��u*;"\�z���`AE\�<�~J��$���"(��;9ʎr�.S
eA��]�aȮ7�eTz�Eʪ.EDW(�9�
*�#��gy!C�	Up��
(Q]��Ar;4H"�����O�����졻�g�\�M�Y[�W^W=��Dt����A�� Π��y����w+�=���Usk6�j��<�=��8�c�8�*������~�����'���b¾����a�����$��[��\�+��o��qQA�n^A��Ʃ��/(�I��_�8½��ُBޭ�ـk��,�½�i�L@I�n�n�ݙX�Y��|�4ŇPaގ��%��9*��Α=�߂H�^ꖏ���'TA�}�)�"�l���F�������7]7',���D���E7��\��O�P�N�S��|Ly�/y�+���M�%��ۯ���y�{��d�	V��3O���/�:j7\J��OnoҘ�0'��ԘI�/A��=�X������3�n&�s�D��W�1��б���J���zs�{��A�m�[�<{�m��i�z�v�)Ny>�,;Ց�F�v�w���� �8��o����0؋���W����9�]ќʈWڭ]q�N�_U>�����]�Xp�,{�w�����x���	���z�)��DYڮy�Y�m��p��vRz�:�Ъ�eln���`ԟXB{� ��I�K�d�2	���[�n�~���<c$��85�3�[i�;9Bsll��<�}���,��^=���8��>��v ��>�ao���L8�����뻻�ފ��ٲ�{�A�ke��#\ys_uӮ߫d�T���Hy^\�*�MX/FrM��8�υM"��ێ:zJ�R�v���z��>�u�����9#�9�8��RF����f����潱��{8^j��n6;�4�ǋ������ʆ��s��w��3�X��{z5jq�vB�7D#�u��!���H��ؒ�L3 �R�`p9iX����L#`��#	Sjc���dդ���K�R�H�M}����c����g2|T_|�H����.>1O�Tioc����t�~�ϝ�����k,Y�imi/�<��{K!���
Ȱ��0��|������̼��̌�z�yR��{C�*��������K>�b��U$�y�,/�|����{`��l��D,}[��{��b�FW������{�K|O˶��۬p̸t��4Jq&MD�{���	�wf��������瑯���vm_�B�bz�g 4W=� Ħ����ŅT�ER�����^�M��t��n�Th��m�mx�([��-�����ѳ��5]�>�e���[�h�:ޏH{>?y��&�]��E����g����p[�2+���9{�n�&Nm�B�l����&D��>ٍx�C���s�NΙ�{�*뻏�J�qF�Վ�1�]���g}�F���ɔ�C�B�-0���g +L�!�\ɪ�EUqmnn�c�#���	�	
��[��X"���p����`c�w�os�9o�8��B_wqP�P5���h��ώ�J�m	�+�0�ˋ��v>�
-8S�K$%*E�?(��\\\o�����ܦ�?@����_�N|s���� n���]�,�k��K�Z�;@���y�����`�����ZU%x��>�~L,
]�}�dOC�������`���;y���px��p1r����s�t&[�.�����v�u���C?!��I����?���v�M+8��i�"��t_��%Ԁa����_G�ߦ��Vt�Q*�	_,:��}����n�I[Ü\��A���;�G1;r<��uGwC.��ۥ��b�t�1������f2��3K�����2��feuRs�VpKlqs)ó@�VjV2];U�֞��&i��|��E��`��XL|��'�H��� ��KD�[)��Ĵ��/k���8�x���m���t!�BqY	���߹A���_�¡�P�f�8�_u}3yu��9�Ǝ��d�L�5�����y{��ɏgD!>0G��GS���>Xh�����_VM���T�m��3����k���G�/��y�]H�@��)򟚶b�񡞬F��!/� b���g-�w��y=���\�n��	�oA���?���ru��l�xH��sm|ֺ�iu�ϭ��e��5�[c�L<n����ª�u��)�;�a0N�t�ۈ+~o��]Լ����N,��o-/���n�}Җ�)���(�ť�ʋ����e������}��јv���F�L���5�d6�oJHo�~�@�����?��	tv���:�Dh�r�\T~�ܾeqw��h���x�/�It��gט�y�g�r�4���8�oV���V�	S���W1n6>��rs�)^�Nh�����/UL?a^��L|~�Q�V�z�M͌��3�\b�𽳧�{y�.x��w��!�X9�&qׇ��I��
r�f��#�7��̢[�(����#n��`�1�.7���]�4L��ڶ.!^�Qӽrw�
�Q����0�N"��;��D3V6�\��;���3��p��`���y�J�7g���p�YH����f!(����w8'�T\�u�K�����.�(����|��b)k��+�ς2����*��%?��l��q[ղ�r9�hwP%�ي���([����Y��߽7���̬0`��Y����_��?@Z��\!������/��
��^�.����ew3OT��b��3˝!�]�����8з�[U��Tt�ƛ�(,��;[�Ĝ=z���>���Ƀ	�m��@��'��c���5�����c���^]��h�/-a+�^xh�����o�f��r׭�k� .��#�ˍ*��F���";�E�c�H�S�7��$��O	$��F�=�,���cն�ojmfW�\��\���1�♽z�y�u�B;���9��Oǻ�眾uxO�˾yi����?x��<_�"*�>��f}�z�V��|���� ,�g��K�a#e+��x��Dψ༧C����.����gK{�_�O̕d�ȹ��;����p$u�f�'����Q-��K����E?V_���`�t�bȀ�t���nV��}��)��י�,��&�M�z��'��$����]t�	��������p�n��9b�!|��y,�ި ��ro��Sr.�X��E-����{�M�Ռ�JT�ml	Qa���>�%K�++��),��J_��L�{��D�Pܥ>�}��T{h�����9���za=� 4\O9�8.|������e��c� �pˢ�F�uI�9�z[�������f�\�B��Mņ�YE�I>}D�HO��>�A1�<Z�t9~�uH���.7��y8�f��U�',q��J~��>��\��#rD�r.���05���{�6��;�w�T��g�m�y8�#�)��~��k�����6Ȯ�����-�R}-���6��vU+΢m����A�C������B|���ɵ���}X�GW����A�Ŭ�$[���-��H2�L�N�/�%�{�/��?\��f��r�?e��w`u]&��,�X@x�v��f�舝&�S�9��2�����g˵Mx8�9(޼,q����{�Fڞٳ������?���������F�	������B��, (�0i
(�PO� �\=���}k}�>�j�JfTj��"oS�ܱn
�'��8>J�}8Q�p>Cxp����l?}�w&���xX����qϒ���M���.#q� ��=K�w�jB��� l��y�� S����kr�T`�������'ϜNK�G�p�U�h�1}�{@�>�'̍-�a[jg8բ��n��8�)� R쑯���J�Hǖ�8�C�q*p4`�,��6����F6��a����r�3|���������ymGuU��^�~���5L�z���{����o��,�a���f`�o���V���;���B�8����:���`:5�Wxy����*���ǲ�Jj��]��IӞ�~�Q�	f�p�r�߱Z: �>�PR�s������/OW������2���9�I6�Iנ��A�dt+�6:�eoT֥~�	,ݮ5)�vt��;G؛�ҹ�`�������I��sJ�콍����l�۞.��'Ia�L�"�U7M�C�^펺n����.$����i2S����|���Tg>3��3/�&Ǖ�B5��o������:�}��#L�
<m6����z������-kZ֍kA��E����)':���Uf"Vm; �ݝ��p����=v��}�H���PI�.n��P��3��/l9=��F�.���}�3�M������\��J��M���ܻ��)&��׮�ۼm�H�Ov=抝����x;�=;{��#y#zo*�����ـ.s���z�{��<�HG.�p��uힵꭖ�sZ�
����7�ڶQ�,1��C���̓kδ��E�=d@,�YVN��j�t�������ot�:1jR��t8܏>�l;�<���^K7�Ij�p��@@�Ӿ�� �:;�_d�0��{n<��݃�U�6����Y����N(� ȸ�|1�����[9�A�ޤ�8���]*�w%�&"�`%˯$.!>C��h_�n�cڛ���֏g,��P��׍�1r����sx�fN/J�*������s?0a�p��^f��oe�۷C\�)���� �6�o�IJ��ⲓ$�����KYm����s�h����F��bc�!��x�dig���hQ�s�ɣ�+;�����1��M��>Z�T�] ���nn�$ǃ��L��{��z=p�����ׇ�ά�g}����pm�x��P���=\{��F�3t�e��1��Ճ�g�}/Į˷���s�-�Zg�� y�V��E�$��U�[�����84��Y���'`�,aP+)/xQ�G����f^�}�}���=�f��!��K*Dˤ�N_�H�i-�'m�VYqg9t�.�y��Mvnj�qM��X���.t�o*�=�@.�����2��ky]
�l��{}���~oHpS^��l����vF�<��hu�`�sM�-�K6(��z&C�NM%��^/tw7���a뭆�^����:�?F�~���I��� 1�;:�q#�.WS�zu_����.w1�	;�e�<]���BJ�m:⻨o0]9��Z�~������uOj�Rg����L�m\�B"��m�foh�*r=�Q<��M k���˵>瑞�A�a���2�m������\倍N��.`! VR5;d� �xsB���;c�Kn��	�{u�?��%{%ݪʐI��b������I���ٙ(����Wu��r���N�h3�o��Su�E�G���������������߽�}x��%��'��c$���9V<f��|�=�>6�$�r]�����E���25�!�X��p+L��"'���L���k�uOG/��FugA�F�wg%)��mEz����N�n0^���)N����!��Q��=�����锶x܃CcO<���p����"�P��2G{������n��>	��_l�T��&��c�hv��{�+֊���]��Wn�5x��O�hX����g	'��ͮO����J��s�[��f���q�6�F�r�[g���{qd�yC<{v���V�"sh�έ:}d�p�J�0�xa!G������S{�(�ރ.�����H��Fb(�kǆc˽���6��T�@g��ÓǪj*B�gfnT.}������;)�ܒQ�X�O����7Ԏ@��
�y��8]��<�N��t9MS�3n�;oh��m��M�	���/���UJG5��l$�O-R�{[��yE6��1��g�� SI9'�F" ��� �s�F����\üSB�<� ��gbW�BoB�q�97c3��o_]ssr�e�t�/w�x^^�:�:�<x��Ǐ��m��U�p)Ύ�N�J�*piX�S'n�Y\M7^��!sW�Ҕ굙�����|�>�G@�m���]����P�ܗ��f<���@�oCk~�9��+��8�a�,0�֞�r"���~>�~�r�3����̳t�6g_>q7�{�z,L�_FG:��'���h��W�2�L���;9���ȫ��z�^Qަ�5ڐ����X:��"�"bUB"��#��߭�^�T�����h�gXe�2���x��B��a�g5���ӦLDD������C�e^��[޾�Rs�/,�����C|����3���u�xx��PL�ɝ���ķ��TMڙ�o���eiO��̘y�ꫲ���A����ꀶs�z�W��kD�����o;.͘�.-��7�F\�[*�8�!��t�3獽z7�lg��g���Вa.86�c
�|rk뷖��4nd���9�� }��I���ԛ�Kޅ�X��n�t��yM]ɹ�9�v]n�Z=ʫ^G��;L��]wO�t�"�V_%n�_�38� ���yw��p�$�ږT�ʹ;K=��}ո����]�r�z���f�zy��:4Y�4Ӻ�<r��U�Pݨu5lWM/�r^�����P�lUz4�e�=D�u��Qav�L�ԓ���]��u�γq���d,�gv��!ä��Y�����:s�]��0��5�b�����\�QN�9�=t.j��p��h�^�0l���1YZ�3U-��Y�+����;r��}_w>a�O8��ΫvF��+���A>�k{*�N]����0��,����wxqQ��N�P��Zt�]]e$��<w�S:�u����b����[v࣬>�-�;�P�����y�ҩi\1!���ȹf��KUi���>������u�t"4��#	�2_⭣M���M�� &ތ�k32�tT�Q�:�b�hVZupj�Dս&�d"��pgQ�G���M5���c��:�=��';:�
��.���T��It�(2�W)�;=6b�Sn�uc}�ʗ�ՙ�:Y��ã��J��dXuu�ÝW�g 7*lұz���b���J�t)����.�d�C�����i.��k�����VR˸�Vv�[o�Z�U�e ��m)��mɓ^\D�k<��Φ1a�$�l`����/T]�˩��j���+�	.�bC��H��X��/�0{�on�7ۓ]Plwg8�q��FxE���D��L��Ty�0��d�a��%r�"����.Ĥ���xt�:hYsz뢚Hdk�������Iۢb	���؎eX�X�Fw�qOhnb�j�!����}z�y(ѣ�B�\׫�u�d{l�!�٦�X�G\������k�u�.��`��ӊ�\��:�e��_3|v�dƪ�WI�v�S�`�#m���|���
v�x41-�c���e�v�I�mŭun�X��[��MX�q�s�0S�@��YPg�w�k�=�ܚn��s�ݒ���*�VEUݜ�w�kv�:���d{��`R��>�{w�:���<���Q�e%��s�=�^����sp����e(�v����\�l���В�.p��Wn�86)�C�'4����b(Ao.�!4,N�ǡ,.���������SG8���s����r��m=�jw`�/c��i�"t����K����gv��3��̙!5��Hxc4���.9�`$J�V�u��(�ॻ��PY8Ы��)�I��R-#;�$��U���o+l^ �=lT4Bp0�A��r% (C��\:ag�BYw
�PfH�4�H��1�� ���B��1�@��Q�B���r�>3e4`i�H��d��P�u���C���T�>]���{~���*��#�r���r�c�l�dE�"(I'�	��+�n�7�oǶ��5�kZ����������|IOԲ?(p���tB�c�;�)̟_׉�������@$M�Oq���Z�k^5�kZ�����������HA��BX�$�$�A��́ܟ�aW*����HA�]q�__Z��Z�kZק�����������xC��:�ǜ'y4�����+J��r(V/$�!�{z}}|~5�ֵ�zzzzzz}}}~y!!��BBIABdȊ"�U@b$?c���WɤOP�z'(�d9�S"���w ���w����C�\�퓞����W#򰯢M�	�8�܂��b�Q��'g�	���;���|�r&���ETO�j�W*�S�ʊ�R!�J�g��z�֑E��E��&Qr�"e3�iAA_R��.\�s���ޤEAC����p�G�{]���D�&!B1B>F�DB(:�#��t��Ol�S�.U�ܬd���)ýe:�k�;��0�:w!�C�֋�kE�����[м�9�)�������8xR��D%Ģd.�㔥�
�q��n0�$��ĉ,��BGUp(�(��'K�������?������=*���wx��v4-:�(��J�D�d�]n�?��_l���[�I~ю�w��_��Ѐ.�Y}ut3c����kl�9��DO�oe���g�g�jE�z�150Qy�f�ؙ�W��� ��]��A-YJF���h|�ڗ�:��jڭ¨e���ַpҕ`� �h�yQ'E��8��\��EC5����{�z���a&���J����Y��Z�i�u�"��(�o�dE��}j ��GL��Y �t��n]�#EO��lx�̩Av�cޫ�Z�r���7�� kew o����Y��L%�d�rם��'\s�lz[���"��b%f��h��1���]�Z����O���e�-n ��qeM�#��˰��S�pwy���3ڼf�B2t��wv���9R���'����m�#V�n���c6�ר���"̒ev���L^����]F"�/��}enm�(DN��f2�*��-Uh�f�Yg`B��6�G�V{�ڻ]��DC-�P�tv�\O��K[F;N�i����Ipw�ɥ��օ�j�i����iMZrѲ����S��7���;�3�y�?�������8t���~��d�G�q�ȵ3;���oD���za�҃��h���M��df�)郝o͆������Z��������Z���ڰ%Ue���ǟ�LPp�=�J�%���� S�i�{������Vu��^fz�=H*K��D���0���(P�n)e�y�d�ǻ��zV��%���[>7�~@�a��+��UsGo;�r�wú������K{�3���yz�kR|� ���!�P�U�Q���g�)��ETM����$O�{Ω��>����3�	T
K}^h��v616p��D�-��	�Uw�T9�io���e*z|9m��u���j�߾�n�e��z������Ջ)��<6^�)\�=�U���[���g5�����'p��W6�A��.�с�}W�%�9䵲ܛ_���`5�����266*O-	H]��!tggN�~�R�����9�g����� �������b��[́��%p��n��52*㳷�v��:*{���<��~���&8�˼:c3�X�g?8����������j�ڽ���/RBϾ׃^ç��gL� 6��m7M5s+����ms�8���w�NF�{��N�}�R�훔��z�h7O�Nq��;��o��β��/u?�_XB��R4�����t&CJ`�ݾ]P���I�1>p4Z��pNO={�W^\u*���=��)�(���]b%�a��f�&�=)XH0�m�֤n�/�W�v�o$=���85uA;s�~��2��37VQ�r�fç��ibGw2�UCHl�}��L�ε3�k����Y�j��q͚�N���Vɝ���Wgy�8-A�iy-�u�����V�qk�'���� 8<��v�Vk?���u�6��6���r��9~�@h�^��Rܑ�~��!�/v.�ޣ8�W��P:�/�9�s�c�i��K��r��sJ��Kg�~>{������Ey$.l'U�+#U�v�؞�������­�1��^�\����c����o�G.�����Ԯ�B�U)2��<ƾ��uh-<���͝������C�.Q��S�1�
@պ7�2:�7���o���k��W�������������^GՓ�Z��@��i�] `�R�<�u[L'�e�3�van��[J�v����$�������~���E�4��!�[d+��%����7۾��S�X��vu��y�J���޿}�ww��@�s?^��~�z�����d����؊�9r�8^�]�o{}��QK���빽bK��Z�ED�yP��:�=Ŷ�r3�e��ʫ�:����\�Ѷ��ǽ]s�g����x���]�����WV�6)x���+Cy�4���l�O�{�;����[ge3g���ꞫҌ����_t�
�@���,�UY���#c���C1'Cf&
���ͭ����F��xrˍ������q�Iw5�P��6j�uAF��1�Ķ߽�����>�>�y��̯���Jw�8��Y[�|@�srB�]�o�䁄��Nі���#���>���ع�%�A�@Ə�sb��~$a���rS\����A�YV�ӗ׈�R]u�X��z�ݧRU^]�� �X�#�]xq�bwum3�y���*K��4fWPɂ�5���[�9r��Y�q�\����U�����[9�a��9����!���Q���Rb��(���$����Y��π\\\\\\\\\�݌Wԁn���VbW���d�,[5���=��#�*�gvQ�ҥv��'i���v��Ta�ɬ;uđ�V��y4Q�/���Y�	A^�y�;Y>�}z�Zb���OMǴg�hه��2xTWvH��$�Ks��*&�/�&��;����0궄j�.y/X;({�o[kj��n;8��Q���ow�w���ذ��� g��ҡ�*׹������s�_Ov�f�&��s��+VV4�����d!j<�ܧ����[:zo�ن`Ǵ�d^��
�Ǡ����X�]ґ��{��aX���ޗǚ���Z����F._�Iz,L����swzg/��8��O�
��v�@&��i{6C0`m�3�H�.6g��3�T�7 ���rk�Uz	W���������;D��ۘ��dFw=W��s�U�m�;	_U��vL��]{_���a��J��F ��YIЏΦ!�`���Ӡ�Z}w�`��+�ƪ��w�3�R��Su�9�=�l��_o�Vs��N
]t/��玤���*�*W�����0�F�.�z�����
%�s�.. 	�v�v��+%����ƶCa�x�Ⱥ
=��9�EY�1�W�rn���d�l��5��y�{���.�fΉ���Z*[γ����>���S*7Z붷V��g��є}*QF3I�j_�����ox��
Kğ��6Vv�=�jg"T<xT\�n]�,�^^��^��5�p�=������	��-����q��/o)ix�L5�����E�A�;����~UD���i��q2���s�bl<�V�^��@k/GG�O�Ha�(ЌΛh�|1��ԗy* \����b���8h2�RE^cm8gl8�ʶA���
\�^a�ty�TI�"�����Ժ�1�E�+h�p�]���M�Y�`{�4@�so�7%����a�t^F^	�;$��,���=Ӻ��@���={�xB{��{c{M���ͪ'Q&�=�����*Y��x�Abq����ᅸ{�)V������!�D�c����@��Φ:W-���p�VM��B�8��u:j�4�����޶�p�:C���#�".t1��uCS��}����U��XW�h>�>�_]�f�7Z9�8&ٚ��$��{�剪��Ow��//////// ���h��P݁���l�&���r��+Ε�j	�M����uy���<{���S�h��s��IP�12��9H�m͒��]q����;���[ ��u���a��3�6�+ã�ʭ��)�4�e
Ɋ7Xv����_Q4ym��Ǫ
�����W��V.<!�[k�b���8K5l<�0fi�q�{����Suq��h�i�p�\�n�fߠ���ŇrBΉ��d�����ܽ�XՃt��<hR���ko���3lع#ϝ��-2M��'N��� Z�݁��wUm4u3x�3zw��9�{����,�?�]t(�k����r[3Z5�c'Ui��{O�х�O���}�`:/w�)[؜�g�{�tv�g4���@��4��\�z��>�ff1�Y�f#:b8(\>��;#��e�g�wE
��R�A��\����W������~q�-�G]0�+(��f=�E�-(G������Q�&N0��I��8�`�Y��;�6��-���dW
FeFz���^�㔣��g����<���^^^^^@u+�=�ț�*��D��UzS��l��i�8\b��;4?kS]��Gz�ӈ��V�<k�D����c�j6Ff��v�L,���v�;�d�V��)� �|�`���\s["��I;��A���W��F�Mx9�Աc�,���;�����5�^����Ǫ4l}[>���!��Ν��s�wW�5i��;��SޟC݇�fl9F^^�"��&*m�V���L�u���9Ʋ���10�mE��X��+�.� ��'G���tqr�id�ٻ��$��Ŗ����A""���e-AI�7>zD]�5���JR�}[���J}��Ǝ��Ro/ORN��0�*%�tp����'��b������ɟw��^f��nq(��B;��>*�s#3�	�7�o�W�5�Ȅ��unz��Ӫ�k�d7��wwr����������k��;���:i�x�˗�j�I�y�]'�p��9^s]��Sf\�վ��۵�}��H%���e4�;���M��j�YE�����rh�`�6b]�+s���'o�њ�6Ά�'A}VqQ�
K���e�g`ط�Z��Y�É�Tj�%'9�8�E��4D�\��d�ϸ�����������SL%�ۓ���^��Bۤ،���z�	��w�غ]�.���x�����Gqg�tHN*�on�V��M�U^q��T�D�a�d9��&��ʌ;����o��om��d��G�=��ڞ7�<)���O����ވ�7}���^=���8w-�i��azy4nϖ���fv�3QX�]�|������s���W��J�d{FR�N�TA�i�d<C��߳=0��B��q��S<���q��iTx��SPv�? V�q!��z�y\K�6��!)[���Ǔ�Q;�+����ޚV��z�o�F^p�&����4��G`�`,�����kѫ��Ȯ���%,-�ɽ�ۃ�Ƅ����D�q����ͱ>�ڏ9���b�=+��z�Ω9n'5�c/"��l��[����ɻ�7�̏e��z����G�꼥)��g v��٭�ei�{���҄8��W"�s���b�m�m����k��Î�$��������
�dj�yۉ;��ܜ\#8�bG��ya�V��=a���7)_��ƍ��S�����sJjw.����{�Rr�_�������������~f�U�ݛ3���dU-ܱXcڥ	7�G�)O��x�gG�JXj�D�Z�T����cșd%�>�5��J�;+bgL�M瞌[�-�m,��j�J�d؆q���.�e���݁��>�<&���θw�5�)nF��{�+.�mz��i�-O,��{|D�� 5�S�Cbp1�3��w��5�������}���}}�j��@�ܳs��ra������٫��F��,�*�.E��I�>��i���������R�2���t�5sWڮ|u����G=P���qq��õl�d	�v� �sI;)�lf�������㞥ҤgdR��?�s�n���{�0مt��]��e���M�3ny��ȱ��R�P+��o"�z;��C,կ)�u���B-vÝok�G�Г�o�7@���K�fm|����k6J�1�w,o��8���s���}\��#�=���s-�����C�h{�u�w���yMd�Wi�g[��@M���=�7^vH(.�ŝ��������h^l����'�ͮ�=�y]�s��#Md���x%e�7�$�f5�<,J���h`<����.�Ťe����X1�����A�p�Q���'*��[Ǭꆥ<���\���Ī�΁\s��{��N�өuH�Q9��m�%{i�����GC�;��P�z��|�Ұ��MB�v�ԏ]�N;/ �*�m\��|�LRmޑ7y<�]�$e��^�<z�ի	\���GV]-��Z���t�d�˒�6��c�Y��R`�e1v���b�]��q�+g/r>Q1i-�)�W��t;�W9���G�VS�E����=fP��[�M��fm(���WpR�er0;�{n�s�Xyy���6m�w`ѥn!�L�Q�ޣ�	[њ�c�iEm7W���ʮzf��(c��ܿ���"���^5�7����]ee#'+�-�kJ�Ν���\(G%���R�U���	���S�m3p���tVx-_j|�ˎeW���`�N����E������]��.�=��!�SY�Wc��b�%ZpB#�[ƞ*X�!9G��r��V];rby��p�yyB��u�Ad �u��O�_^�$�?u�r�co��r>���ҁk����ڧ���g7;�������O���;��R��:�o4d(h�!`��8Q�2�h����Q�)]�t�0��o-�� �dsrn�v�Xx�]�Kݹ�h��c�qd��W��T�6��Yg5-�+ruai�S���N���+%j�譫�D�"����8J�\��nʧ�H�鼝�=-���;�V8�|�ec���ţ�w�F_,�����]���ʕ �L�6�ft�|�;���̀��;Wʆf����5RZXqWbD�X��j���/k��:�b��	:���y�ٔ!pq��oq�.]Wk��RʾN��-�"��R���J�1�$JK���f}�f�A�K1Y�;go�Uj��{t�^���d{�4%���G�/����v��z�@)�`��\�ƹVv�i|qJA]E8^��.�t��;4^	�Z�F�4.�f�+*�<��oDW�]˩]�0_v�w
%H�yq���h�X����QmX�ܵw���}W�o	oF2.�]�� �S�ty���S���*l���X_]8��/�C��a���[i�Z���/Zh�9����gY�u,�*�򰩅2��.>�2"�Z�2��H��o
'���oo�����Ʊ�kZק����������NL�(�����L8QQ�ʟ�8II	a�8���^�_Z�Ʊ�kZק���������$�Y!�ĝ�9ȲB����}{�U����u����|kֵ�zzzzzzk�����'Ȓ#"B�H*��d��s̄�� ��8������cZֵ�OOOOOM}}m�ܐ	$�!�$�	ȼ���w+���-(�e�B��?��E������AD|�U���	�"��I5���"$&r����X#l���gN��J� ��;�������#JvQ���dDܬ�H*Q8kMN�n����L",���-iӔ��Ǔ>���Ni�)�]�$�Q#@Bbp��'9s�˔Ev�}��xh���U�&eu�*�,�~I#G����+�t�_[;xGZȩ�q9�v�ha�x/w��������������(���޸���T�f��{���48CL��N��9��g	�2�f䕦ʗ�4��N�ޟI�``j�1���{�����Xc�'3�P����2*�{�z`f�RN��i��|�:�w%�eT�;��dh�^]Q|fϛ.��g�s�ⁱ�y}w��)�Fpӆw�\��a���8�Z��%��ҧ+��\�7z5I�^F7'y��*�{6�N�Q=�x�o=�Bp�\�0s��q֢sF���D�p��S=ȒkI�������aW-���xB�/v�|��"�����L��1�M&��y�ORK%���Yc��slM�ׄ�w���gܻ�@os{G>�.�Ǻ��g��v��
g�iOқ2�݋
/Mf�r�mҍ�^"���2�}-�
z��wvc�;��f��(�x��&��s��.�]��o�b��׌��w&��v_wU�5��*�ݹ:�ڛYz���n�2�wt��D�$��h�9s�2�G+�dU�;CΎ�}��ge�_#!)\k4�м��_Az�0W�߼��?�����i���wqp�m��z|܊)1��P�3�ی����&*�n����pO� 0h~�oYGhQ�$�oN�55�)�J��U�$`w���f�%t��m������f]B+���m{;}:�v�bؒ^�'�D��B�Ą�e_@R�2��>7�kҨLoy�<�=�[���V�y=Ȯ�0 k��y��u?��[et^`��Bv`xki��7v�y��kǄ[	c.n1�*'|��S�C0�M7��E����_�v4~�^���a�"�|�RR ,��]��ּLL@m���:�R�������]��+�vsECn�>�62��Bs�]��S�꣕��^����+�Ɔr+`>����Kr�K������0ws:��fY��9{���!���lS���_�=����Q�Ubݮ�����	�����U�Y2�#�I�ݼ+��j��+�s}h��j�^�t��M�.���LY���t�N�f��B"�JrD�k�����&�WEܕʙg2d�|;nv	�,>[�gA�6�Eժn��&��z/r����b��PJ�SM�H�[���R��������4�����������1��-�7��}٥uqfj���գ�$D���K� �2cT�<{����-��PT97�v��5x�SU[�r��J�T/;����3�0���4|8�#�O�h��C
�ak���צ��GC��+1Wz�[����"��;75��U�CoZfk	����;+�A˻3�5�@[Q�+}1�����T��Ե(�g��h�0���>�������\
��r/�9�Hd�곪Q/D�ݼ�=(�o����>G7�����ƌ�]R�A���8N�{���{�j�2��.�OW��g���J��sT��ƅU�Gx��9"�@���˻�9ɓ4�߀������Y��lm�v���o0��9lB����W�;���|�}����Ү=*�=���V�Oי܍d���F�'���S�e���ډ�����:oڥaU���f�M�Amn����w���4�Z��m<��o`��]&�����OcZ�=n��὜�Q��7X<uc޹�#��GG��y;��f+�j��9�WwL���7��3�E4��d�[�Y��S�op(^uu��Վ�������������&IÆ
ӵ��U��e�
|jt��'�Q�u{s��b)-���\����塻��	�� ���ͣZ0s��mxF�۽���z�M	�5�ݤ��@�R�o�t.�r>�c!���B�2��^��]�|���n���$tἤ��Y��HԄ{H�@�������Ǜ�y˞Y�6Ef��:p�o1555�G'՝ޔ/�`W���l�u/Dz��f#�S�o����1�窞�b����e+\\;��49z���%�j?��ӯ$BF$����A���7�g���gVp����uyzQ3��Btﺇo� �u6�x�gC79�]���y�E��1�\�F�n]ibx��]��K�%8/�[��ߨ5{�[��0ZsZ<Ma�?i�����Fo�n(����^�>eςW�@�����H�4߁�i���H&��������Ö����OU��{8,W˪�uX�\��ؽ�ڮ�:��J�ǔ�� I�'�@)	�ףUI���MZ�86��N�D�U�|S^��y`Ft�`��q4WIcr'Qޅ˳C˝��߼��������z<�>ZK�o6���>��19��⨚�q@�{y��vB6c���{s17��w�kT2#�j��F=jǧ�v��IJ��&V����S0�n-Y��y:q��V6��-a�Y�X��+���{u2����ob�w��ew�[�-����l�f�v��Br���.P�]BY��a˸��[=g��os���l"X�
)%;����������y�7�CL8އV;bvj���������௼�|I�@#8��[\XH(ha�|�8_�?�5*��ڭU�h�ɥ �*t���\z�n��os�kM<_C�W	�M���S�"�^K8g��ݛ�y�1�QB�6&�n������;��L"��yy�����oO�����y<z��^�a�����/�b2Y�rUV�j5�{�k������8�C���	T9�L��r����*zLv���Z�6D�?��e.�m��9�#�u<�r���ѽ�L	j�N`���>��ə�;��uVi"�� `#�!`�	C�"OE� 'K����X�� @qX�]������yѴ�Cе�8.�k��Gmh�	��St�����!�����������!��zQ��z/�Z�_���L����bR�A��_t�5�؆1j�|w�3�l��G���٨�GH��Gm��z��R(0�\zl9���|�n�9T�4�]�A��*��6Zva�7#����2;n�˓c�\�0h5�4�.�KLR��5;dެ8�]��Nh�9킑~��zz{����|�3OL����v��z)���1nk4s	��E,�5�-"s�#@
�v�M�5����cRv>C'Ͻ�n�	�G��T�|�ם��Y0��}gpG��)�NLn��g��?H���\�֕v"[S�4�:��ܤ��BVl+*7�n�G��򆺶�m0��&17S=Ӗ��R�9��.<�s�DʟHԢ̟˯.�)�N������nڲ^[���[5TMR���,���'���J�W�|��7��r �23%eY���9�X��]^�_J�?/V���K�=Ӆ���m��̸��u��}��Sgd���ܣM#� ��S)%�0}� Y���J\�{�>ŕQP���殩�VS�w���u�w�u|K�[˵K
j`�ȅM�\=ײ\�qXX���&0HrJ-m�@�H�~�}�����������w�S�߲�o=�����.���I���2�e}�p�`��?,�\R��'��27k�r�<�L��Պ7����g����	@x�U��g���4k������P��-���I�XV#�9M՞� ����r�^h�]+A�S����I�'	�x9�_����F��Ǘ���5��Y��Ӗ�a���8fv��:���js"�g�i��	�	�2�i��=��R���/��������Z}��n;s��Dȩ�
|I�A��uH8�E�sc{/z-@X��Nv5y�`ז0�q,<e:1Y|�u(��5�a#p����-�	�:��gYT)nHl��Qq�4Cڍ�y�Q:5ـgg��ˀ;{UuS���:�i@���uJ���;ֶ��Eܴ]S�B�����j�LwU6ʐ�^��,C.�=�=s�
}��<a����p�=]�N��y�8:�����*	kzE�<��+:�L���n�y�Mg��,����H?X#��N��_;�h$`� ���9.��/�f�Sy`y��QS�S9�r��7��z������x����\T_*����$P�����?����hŷGV�����d��A���-/~�h��jG0k̈́���Gb�;�0r���vc+s�=={&����ɡ�|��Z�g�^)����mf�G����/��z|7��/w�|�w��t*�{T�]�X�7.�+�96����C���/��"7�VOK⁻��&zۊ0#��iۘ�gi4�' ��,��ǚW(�wv��y�au漩���LFmΤ37N����W���y�w�F��d-��z4�G;=Ѩ%��o%K���g��n��8m�����0�j��!_�A���İs"េ�������h���ݛ2k�T����Ef�m9Z�[����Bki��M���Ftυ����526�G�RU�of������d�n��.�oٷ믩}�8��J�<�5Dm�*�=3m��3mD�t�;����z�a�CT.t��ta�M
K3�6�-;
�w̿3�'R�35%Ik�Tf�҆U�S���vۤ6����ٓ�8�윀�:1�}t��ֱ	W�!����Z�M��,�aXXz&R�4Xo���uN�h���\\\\\@..!Ɇ˻�uQ��vk��7����g�T9_�D�g��c	���=LТ����w�&�ҍܘڹ�k�f��~��zt�ș��,�i����� �'az���ITP��K].�n�n�]�rhڮM��qmV���/�\���ޤg��)�����0��}��}��3f�wgv����`�����0�v�ڀ��Z���m���]�7x�f�͢���n��Z�p��b8����N6�3�;�TY6�M�9��£�{};3�=�ܬd�,j�'=�ښ���)^�b�����"ON�gf�^�k�k��3=�����Z�.:C��u9�m�P�����j �jH���p�o+_�9�E�0mx���DK=L����F�wM��r}��>��*�\NP$��"�p_�Ac����9��.µ��)��7�&�t[�p3�ewr}Iu�wϸ�mIhVر�N�
�s73$7Y{��\ ���H�>�$��*��2�,"�')}w3�ۨ��&�.ՄG���ȧ8;�����p�[��Wf�S��}�����������z�-[]��j��l��*Oo�x�^���E�`�
�6�9�-0r����CF�򯵑� �{���cF�sߴ[F�'��d-�Sknm��T�4�D"դP$m�����[j�ﾨ���l%��F���4[1�-\I�k	�²�}A��3�/�;� �Fgfu+"2u�g������t�g�Z�g��l��7E�7}O-Ŏ���Ɋ���w�jsv�&ꧼ{�D@ܲj�t�%r��ji��l�����6{����0�4NaR�����M��>�q���ǹ���g�Szޝ����X�&���;�{��\�K0b(ATv�dj�zz|�]֩��MRN��p�7{=�<�Hl�ᗙ4�wk�ܖi�t���ٟ({ˍ�$U�YT�Y�䞎73�k�.�O��'������D&5[Wøi�(~JJ*�nC�+W��e�����{�\:���W��X�}��.i���L��7�Tk�_s]���*���e�cF�;��L��1���ؗ/M�ʼ��G�)�Xy�����I���̼�nX\(��lGY����˨S2,�j�`� #�We.`�=Ҵ��y��V���L�����w t&�VUpBZ�rj�+�a�G�[N�Ou�K�tv�Z�W�XZ�/�'Mc�����F�G�� 
T9RM���C�8�=:,y3M��紳��܄�����S=�n�u>�kI�&�+y�A�b�2;f�f�Ÿ{L�B�WםV�Lc"�`S*vМ��>��R.'Y��3�u5��l�d�g�Qx��>����*�
+��tX��X\�K�w:�38��nm�r=�e�K"�v��
�[�U%����P�|F���uG�o-�AV�7��I �;f�\xT�d�@�Ts�)V+�N��!۩K�ܥ�)s�����a�Y�"�s��ST(�p]^<+v��+��<�6��i0B3���7Cd��tڦ�ml���P����Ǔ�gw0�.ﻒ��-F�&��ǧr`Bos�W[K�N-!J��G�FD7��v��!�Y��:rZ�ۊ�`�	XxrX��*%�@tS�>��F�Ψ;�q�,����%*}J��͒�ԑ���(�b#��E:		�_#1�"ȟ�*2�:[�M"M ��R&�<�ht�:��.�R-��u��e-@��qֵ�,4r�'!�ba��2��"S3w�.�D.�_f�1䃵Yjn��*X#��ɴ�H�X�q��k_ ��^��'@�;�stGq>�l!�q����-Sf�0�5Yj���Q]��)�'=���T�y�q���z�TF��gY��=Ɔq%8�)��U��MV��N��U�����l�Y�e����:8����9�R������]��ʹbT0x�n
�$Ù�}Z�w��ԴzѰ��}:f�I������c^��i5������A,I�K�n%W�&�=����D���Q38���;�[�U�P\&�����ڰ�&]%����ə�٣�\X����ɂ�̴�J$�
�,�N����6�e�ְ�E���ʺ�խ���׳��ݢ������C��rۦ�e"D�����Z�Ӛ�%d�t"�WYȯi3-�̩��g71�ﳘ# ��P�;�e�2�ZU�ۦRٺ�m'�b^N�J�%/_@GX)�Z��Ϟj�����PE���M���{`���虯���٨:0]r �Δ$�8{��a;�f�r�;+���j`�b��B���3�L��&r�I�O�����%�%��d��1��(�G����"�)0�iY$�SjH�E$It�]�͇T�k�'�5�l�$BUTLF��!&�I���H$ K���i��	�E6)BH�'<d���D���M�$z�}����FQE Gh��i˪)�O䓒�|��Ϻ�i�^�Z�5�Zֵ�OOOOOM~�_��c��>�_�� �R��4BՅ��3�u�f��~=����hֵ�k������_���1�'�S8�YE$�B0$xr�!3��"�z��}}}}kZ5�kZ������־�ۜ��3�%�N��s�Rg*��i�sBDI��n�[�o������5kZֽ=====5����!����NM+�.S����}�&����w�[n��fӑ�/Z˷l�wC��q|�|�)3��Q�ϝ�J ]3���|��3=��tqDE�r���-ߌ�·�Ȧ������8�	Qt�X��RT',$�c�r��u��[`�K"��'2�D�!粃Ҩ����$RHd	/���'-�d9�>[����.dj�(_9~��z��$C���j5��򔦈HԌNf�,�%D1�Jx��+g���#��A�����7лEl`��$�O��eؚ6�}3z_K�m˘o^���]��8I5,&�E�S)�q@[e(�e6���f�1qӦ�C$��`�(ѵ@��)��wR���|�Zֵ�kF�??>�����0��mf��O��{�+20�#��57��O�{X�q=��z��%���������ިΓ�f��X�lq�s�Gc=^;��tW��,�l���!2���:=�խ;�+��F�{];����]N�VV�F�/^!�Da��̽���v�v���O�.�u��k�J��׎�Zx�&�>7��=R���$:=� �|���.:�T򵯓>� x<
a=�Y.b�=Y�=�{=�h3�vt.=��;?Yuݾ�n*J������qr�K:	�l�/a��1���g��?�j�W?�D�.e{c��Eǽ�����=̘x�^���z���B��~���A���8��ڜf������R��(�39���]�l� #�&_�z#:OPH��Vc��a���L&M����b��UL�Ja���������\!�izz}]ݻC�5h׆�������7R��v2d^#�[ױ�n�j�������맕��N�+We����¬K����6���N MG�Nu�]�
˛8�$��I�t�� z+�j#�[x���Q�:��ͯ~�7����y��y���3uYo�!U�GU�o���,4UW/s)�;7*�Å]����m����װ]���S����G��j�)���#<�u��{b��.��.n
�{zR�~���a�x�[�{�KA�(��Fչ��:��I[ZC]�{/���l3P�8�����
���"���K��Xe��_'�g��ߛS0� 6�ԧf��9�I9��dW�p�lR�׳����/�)�L��a5��3b�����4�A�[��6�[3;D6w����@^�Gt��V)���{�4���]����ۑ�y�v*P�g�/?�t����{Z)�� ���'~��r�}w�M���3� v�{����0p���s���ɢ�m<�g�֍rNv*Dݙj��p,8H��B�`҆�_Wq<��zOmRh��'o�U�Oa���.8`�!ξ�\�L����|=�s>B�ˢl3�;���0�;v��ɩ��]c)_	W��Ť2e�u�mvm����.�w#�{ˋ�Pᒸ�ȱ��)�뛜�Se�+th�u�*_h��7����y���g+6V�V�yN�W��knw�ؓ�*=��[	s�����yuj�F���<����Rϗ�w��5\�=>��{k�s�����n�Ou���~<f�3�� �t*�q^��҄�%���F6e���L��T����x08�\p]ꤼy�߮p�5�5觘�95D�H�wq!��gw���?�Yh��χg3��Og���К����n�F���v|+[�*���X��n홧�M��8i��ǻ�jͫ��TskOj�a� S�Ǥ�r]^\|�US�Ӵ� �ċu��9�r��4�̾� �`���*c�q��z���ܧ�mn�t�-,�4V���%g�O��l��k�'v:O��nx�`�3˨q�h�e���/�֤��5��W�!����ݔ��ʡ5�:O��<5뺵��;_���3\Ϟ�?2��̴39�J�[��ϖ���b/��Q�Oa����^�UY�Eʑ��j��ŵQu�I1�b����ϩ^N�v��[�u!#z�D������Oywz0���ϔ�G�#�#yU��Gw.foz9�?��
p��C��t>خR:x<AFfq2�$�>����w�h
O�|2��h����kD��{ș��p��'����@_C.��"=�<��myw�gwue�Kc+kc��xא OG�����Gw*�f��o���t��W�	p6N����m�铛�}Y�o`Ő�^�����R&��ȁ���%����j�b|<<dv�S��\O��ǇԸ����㿽�B��o�q)s�F�O��sV�֎���͈>A`^湡#=�&�%ݚ���ٞ��l��7�g��[՝���8�6��@��#3��f�?E]d��Q7�g��w	��X�'i�זf�K�p����]��xc������QΞ����r霽�x�RW���r*iԊ5}�ߺ�����hd��T�M�r�}�iԬ�}�q�h�ѳFi���6��`�/LKXB�X2�������@��j�T]����G=�X�יEF"F�лt��Í��u3�,q��Չn�ަ��z�7:"{��sr�]�{�Jz%��p�6&�p�
IQ�`����M�����wç��;9�9��ꣵ�xBwoQ����8&/wj�f`��:r\��gU�� r;�=���Mw������꽳�n�Ͳ���\g!8����Pfd��*���wݱbn�����+6���6�W�ld0n�~���
v�+�|@����������vfT"}Z|wx2�,� n��Cs9^��pwb.<��y�Wr���G�0f��vԬNXn����-���_2|Kku�bڮHOF�>mUviͯN�u�~�\	6�$%���6��Df�v�
�q��^6���#����1��9��-ޞO�3s���g-��\�A���oY��y^q��[�l�Z���ƾXJ�	oK�¥w��4�3�{���N�|7B�s8�6`>q�q�W�'_$l;�磆�W=f�����v{Vz$3�w�xX;}~x�O��ۂ�J�Y4a��n���"�X���).���T��5�[�+��;9��N�jҷ3��n���0F��j�9�D�H I@�� s]̺L�-ƹ<�����nMŭ2I	��>���lTuɥ�\0���%�q�S�^�^>����y���J�'�v]��(����pu�1p�4+a�v!n��xy�wf��64��L&�'1q���r�r]�r<�c`�=��\�y�+�������$��3��x��%RDf0�X&�F4I�촵�A�#u�h��:}��wǹTY���0�mk�z�Ύ�׋�;�_��y�T����:�
�*Ug؅}Fgr�?T�g��;�K
��^�3+n�z�&��\�z�{�Y�ro�Ǟ+gX6�r�v���8�q����-�$�ReeK�����]��CE���;Z�mn���W<^�����}�L���w�aoV��o|�K�B�y�6�����O���wn��c�tv�g������+�ҭP����-�p
�� I��=�۽�����}a�wf��&/^��U�{Hɘ��4xl#f��|;��t��^��h�Bo_-,�\�ڵj� �"��wFNv�;=�H�7�N��qu!ws]Ɋl�w)dXOv]Wu"�qF�K�]��D��j��#=���=��Vj��ia�����y�~���b;�[u�@��}�{�8���&�n����|�����9�Y����㱝�~���3J��gs�r;�={�a=]�h���6333�^f�����w���2ʩgï^^5�)���^%jG�^���MC|^���j�,��<@��~�]���t���[�`��w�Mw�:g���nso��0e�.#�Vm���tѕ���2;{��v^W{�seo��������N��Fy���@/\#/r~R#���P��2����ES��ʵzPvN�����G3{Q��f��U->�N�#}�p�N��"��O��*��k��v.�g"kؙ?�EAu�W�~����_b��9D�޾J�M�i�j��sջ{ڪD-^Þ�Q)���m��<M3�	��GU��O�?N^/��U��Q���7f)�s\Σ�n>��l[G�Q�E��m5�H�P�܎t7���nᆖg ^�V���I�Kbuv�4�H��JΤ-�����z2>�㙒V�S���n5r�f���zv�)<?x����|@N���In�s����n��.mJZ�i�ܜ�v�im��*�X�wy���g�%��]v�_�`�0{�����ӻQ'�PP)4�"!���T��� DCC���vf���bs������o��=q;=�j�ʴ_Sct��5�fR8kom���C���]ّ��3V�w��4���9�����&��W�׉�}���l�5{a���i��
���k�R��>���K%-;�,��=��U�;{ �[B��|*{�>ߵ|��6����c
�N�;�|�=��H�Wu-�E�D33z�v���)���c���6�C��*�'��^�/������9^#^���dW�)�Ho��FF�i�$L���CDoK��a,��`�B��q��`�\�fCX���F�46�yu�/D������J�_���2��Do�W��W_}2�S�V��6+�v�c*$���	�yh�n�{yAZ����k���%<��ɑhލ��MNH��{4 1(R����u�0��J���Ѕ�אn��WG������r՚�p�.^nu�Pv\��QM�v'U�(��:r�$͔��P�тBZ!!$8C-�h��(q�9��x������V
J=[F��Ot�E[�.jW-$m�[�6�'�r!�U���3>ا٭gA��+��:zbjM�Xƽ
f��z4�&�ׄ���@�!C^�o_��.'��z�t#�DέSS]~�$�4N�܋���sFlq9M��nX�6p����A��5�g������nפ�"'7��z����z�܊�r�۷	'�s�t�Y�^e�/R��D�[��W����dVG3�玀�b�eY7}D�,2���t�z��G=s�W���� F>�=�UWv�TMeR���j�ө���Y쑓������R��15I�dQ9�U՛����9�b���/�[	�G����w�Xr�>��++;Y��0� �B�2�/~�ɮ��$�u%��0wcϲ��X�B=b�8e�f��xdL^u�q��x����#: �4����g�-�5_@R��s�����e\ڂ��]�I��3y̕:��p���-��1�J���˵���:�0��ݴk���g݆��B�̓|h�MW��!J�T�qv��ڇG-Go�C]�!�×T��9����`s��{�/+��,O.k��^r�9�?BF1�b����/_/�/��?>���1�ߩ�����D���36��eMc�	�f�#�&���.��f��;��/1��o������=�I��fz��d�\k3�.'U~�A@�b3�!�9|�P:�ͳ��vإ��*�tS�6��|�2t��De���,N�1������s��U�o���:��su@�o^Wwr����
�Eϥ�pwB���ӂb+�w&�8��<���&5��2�ԩ�ꔳ���{����;RO~3��Fw��]��w�Ȫq��q�/Ai�4��uuuZѼ�n\��6����":�����њ�;���ҁ�e��a�JV̘L�n�ѳY�,��=S/^���nO�N_�e���@�{ �����]>���Gh�IoV]��㸭�ɦ|�a��g�h����
����m�D̿���V�g�[ͭ��;���/�����
.Ըt C��:Mї�$����T�x���]n���|���J�v��3*Լ�Ah��ܤ���mH��y~���9���j�<IF
mD��w�B��4�Y��!�`��R=�o�f���������;�z�=޵�:�v��h
ֵ�c;q�6�����%���F|0Di�/oܲa;�oc����!	��铃���yZ
�n&�c+��G;���Զ�;委�Im�j0��e#4�u�mZշ�C��'i:���Pt�y�Q|��=:����U��`�O���,}�kTa�->۠���V�0st�Ie뾔��`d��J��.�fD�(���>Ӝ��D���3�`,��T�k%��ܒ����U��ŧ�S�8+�#�n�A��D�X���r�{W[�R������X����f��c�0V<a�'�Z~'z��1�*��}�N���3�RA�� %ѫ�(�㧥�q�Μ}�q]�<�RSBb=n��\`սh؊�J��̰e�*��}B+2r��*��D��2�P�6�N���/���um�U&�J]�=��<,,�x��g���z@6��I4߭w� �;5^۽�f`8���D"K�I�S�1GT;i�m*q�4!���>
��xV�+�DIi��F$6^hLt��e3]ˡ����vEw\v����j�=˜ƥ9N�]0㧅R&q �38u�-�,f��Μp��yXcA\��eΰ=�X�3��~�og�ǻ����Ȼ�^H�;�'�m��49:v+ǉ!�d�:M���Wd�Rš��T��Kե!�$�}JXI<�:�mR��C��O�o����W��Em�JõɁ�͝�+���C��P�گ�<w�޾�����R�}��.3���K5�+����8�eQ����1\�׊�J��ZA&u����վu�諍$������S���ۭ����v��m�+��bu�ڷ3���V��K��p����hx�*��풰j�}�b���s$��ӕJ[um%��6�R<�*��gmژ'sV
Q��6��M�.�իi����`� @�P��6��j���{��l�M=����]��:�'Q�ƷGM�n�R���5Z33�%m�-��D�s�rk�)����0���"����Ԏ�A��`�`^7�彷�}<��X焸3�̀G�'��d�.�R�u:sX�z��a�Yͦ0�RX5�)^.3-i�v]ٔ�B���PO��mL��vHo��Q�/��95v��p*���i�2�����Sܾܾ-rɱ�!{�s����/��j�keu^����
��)�5��`!�o*q���3�)%�H*���u�f��f��m^U��w~��8W
ػn�.�c��:齜�GgwF��9����h���>���O�$W��+rHJ$�m纩G��*�:TTq�"t�g8On����񯯭hֵ�k��|�7��~���~v��R���-C4�gy.�Z*����>��UB' ��c?��[���������֍kZֽ=====5��>O���H��SW��F�]�TS����X�Ws9MҾ�����_____Z5�kZ������ֿ<<�PJ��J�N{�;���w���,����j"�cwJ;�H���a�8l#	���]z~>�����Zֵ�OOOOOMk�󇜎Q�Hz��(��A�
I5d�}�v/��$�.U��z;�s�2�����U��!^V���V�����W�nl�Q��r�Ô��ܗ�r����O��J,��9Z������� R�?#���S�9����	�<.��/VQ�MUYp���8��
�Y��9AS��F��E
�}���Յ�.Uz
�YBW?�3���L��+�|$���FeU:4=�G��AW~�U�T\�9\�b���$�D�H$�uJ�� ������OI�S�n&��g�M�˩�{��Q	>�V5Q�܇No�/Y�<z��>�7����y��>%'cq-��#7⻧���>�ܿi���)=�dB�r�U�U��\w�-��E�O�I�64�^�����dndm��1�L�p�h��X���9���NY�DC;�`��{U�ot{�VM�����0��"d��o���߸Z-����β��]'�gl�P�'E%Ԙ��=x�L��}��lZ�E�|�󍩛�����-��ΈW{MQ7�ј!K?!?F�t�&k��M�}��~/>���C����gE%�F2%�ZjMڔO�w	�+��>S�v��Cok��#��;ԅ:�Jb�g;7{�\qˏ]��i2�Oa:Z�B�;��Є�F:ޣYڰ�f�j8Sb�WF���t$���vϱ;!�o�%�@��gR����9D���\����,��=�CG�%��+�|�S��F�X���3�w���Qr:ZU7N���و%�X��D��O��'�T�kD�G�F+�r�����5IT/���{j�|ѓ3��c훺�>��Qřt��� 5��7a��Kr��m�Z�W&�k���s߼|||@o7��y�$�ZuYoW�)���WC̳DCK8`�l�x��
�>��æ�\_.�"�6(敦���爑{u#z�6�C�����t]O\��'����w�v`���L��^f� �RH��@S��`s�l��m �������"�)��+�4�=��0�V�Y����h��]�W�j��(v�-/UMx����;�<�3Ml��$@��[�˥�UO��m������2NFL�N�o^��"�`�ONx	�'tv�b=^�~��U��oDF�Ol�7�{�~�:�βC����c�0s;g�f`��g��X�+o�V���6��k:�V���̰�������Y����j�8ދ9��5���}{D�Dϖ��׽�m�2Ͷ#Zደ^�ux�:�-֚�a�����9�kߵ��RG��Af�w^��^��|�X��o���O9���r}5ۅře[��4އ��{�?+Pv>��ݽ�w0�
�4����7~�}/���Cs\�W��~!�u(���e���� ֺ�
���J���Q���o��B��f�fY�_:�o��s.�����Y��J��#����]�A��	0Ra%�r'8�y��o7�^��z�jS�W�M�ͣ��e9�2���	�c^���O@��{��$���ӭ�����y���kM:����;uN"ݞq��6�8�wTʼ�-��ԝ����N���WjB�u�5�-���=����8�Fwf�B�qC�=7���z�.T!Q��x��<!/��mB/���f:��c-;U�t�7��d0c��=�I��L�!߅�`��*��^S�=7��3|N,�\c���yz�]��@��$q��ȃ7ƣ7��a���mBe.��a���k���F�7�>����v��e��*�4�w�D�B����n�y�9�ʱ���/��g���yyx�%t��\I��������c��hY nBU�Ǹ;54�Tt��޻��ն�s"YD���O�<���"uߘ#�f&�x~���rg��`�Zdw�5�ސnt���S��k�T�X��G=�n��,p'J����;���pf�j���ҍ�X�w�0L�O�z������P��m��wn'�)h
��:9^ŷZ��ܳ�L�'Y��)���}%b��c}�D������ƒI��Q�����[q���8��v�b���&�=q[֓�k��w&�M�^�p��yȉ��Hv���}��5z��wf�z�(�=u�I4������b�Qwf��UH�ͳ���,��D286<��nZ��8o�%-�j~���ѝi�-�z�o*�f�-����H\����>�Gmʁ��^��=4:�j�FI&��a-;W3��yoxӃ��l-����+�9�\���I�K�>|����fv�����5�oz�6t��68Ϡu�S��}�f�Y<��;Fɫ�.��L���	�3��aވ�¯�tn��م�3+�ۚ�{��7Y+�<�]�V H��W~_%���C�z8���o��Lnei�A+�ԙ��c������j�5�ʜ�}����C���5��5ODe)�w�B6'^��KV�;��ĸ�b�/�z]�s�̾y��Ȇ�;���";y�fH�wK��ٍ�	 |�U��z���{��E�ר�5�ܚ�ֻ�9�+��o0W���T{�p�ۻ��v2Х&�A���8y�V(� 7�y�o7��e:F�z�D4UW�E��Ӿ�3hG�Vs�YV!���\?4�+�GN���?�ԃ-C��`������q�=[�I���$L���I3��^��7~����p�X�с��S��qh)\�rI�C�m����<#Tv�U<Kp[Ω�8��ՁM�F��UG�i���w��.i&[!u���	�����t�
�F3�>9=��4�S`P��4C�#\�U#ҍ�k�ʛ*�l�[D��w3�E�?/2���o��U��Ҍ��d�\��]%�u����ƯI�Ke%�5��5�vC+� �ݏvF���`O^��=��!�ej��QӨ���������?��+�ϢLw��QY��3s����c�����&iW*�o��_��z���O�K���AŞ�{{j��,9VX���:�����k6�Y}���#� ��gH��D���a��\8Da�G������_n���M���]�d��U���v��3��O�u:��u�-�e�(n���gM력v��G*}��y�o7����[�qj�����^>���
\�`�Q�9O���3���5�b"b�򯸞��	@��6V;I�V�F�2{�GL8s���L4̘U�o{�B!f4�	�� UV�C�yU>l�U�w|��8/ǚ���f�Kn=21��d������3����h�X,
���>x����C��{1�9	D�Զ��/Gm��
��AB����i��.��Y׳��,5{]}�iZ�]3�-8p�4^ِz� ���z�o!�A�ձ�d`>%�\ղ�u[O)e����%
X"W)$�IۏTK���Iݙڬ 1�(�YO��ǽ͹�UV��1�"�Ȉ�S����A@s37={�gz�~o�����%��7���u��yy��ÆRN%�.@t�IU����&��]M�ވ����r����o,c0q[1�'�1�u�M�z��׻���؀a�����K-�l��t����!޽Q����ۆ���j�$��d���S����.�G�=M@[1""N2ȆN�t��v�LJ���4��S���}I�Y<��EJ�-JC�Hu;5+�B9v��Hރ�k��{f���R����M����{����q��r�����9����߮�gIxH�{�/I�s�0�x
D��!It�^A��@��}��[?I�m����P��{zg���]�eا�Kv�#Z��7��S{g����M�s8gS�\?l%�;���Ѽ����n��=K������S���l��aO�ڛ�63�7���J}�d�_}�eH�@O�ҿ����މ۲�b��?�q�ȸ�ɮ�u��<��n������=q�pY���}�UI��� �;�+6��]��lk�ż��{Q�
���
��uh���)���5�mh�����KM���b ���s����ـ��P���Á�ۺE���z���.�fo��g�����'�L<u*��U�8���o#����G+�XVl���bqa�r��H�hsK����$Q�wt<����Y[9��tŰ���Z���i��ja��b��P�|C���#���`�-�ӅRP�Vv��F���7=2^��r���|uװh�{*�ry����w��v:�T�Tw���A�o\6��Wp���vr7J@MK[���`q{jNfsr�m�ɲ�_k�ڷN�CsWE��>�< p�w�Z�h<I.�be�]sFl Iʷ��n�����%�n�w�WC�3@v`u��_)��#/Q�0�-���o���Ȟ��Vt�0�ʊu#�mG\z[�@G��x���yo:G�/^'(TM�bV����ͯO����8+�?E�Bv(F�,l�����Nl���F�+RW�)	g`̞�Af?q��h>�����:9׽�׾ʭӽs�Q�>1G�U3��tfY3�!��O-�3�0j�v�^���z�W���f.����f�Z�s��ZR丮�����x�{����Qt�in®F�G!��~W�U�s���++���F�W�sB
iR���X�x���^�g�wg��Θ>������@H��ܮ�fn�a���J�̥
W��7=���>�>a��� ��~����=��x�֌h�Bq�c?�~�$y+nZ�����Ob"|�XWp�;��7>�k4�[`xc={y�<]�ߓ!y�� �D�G4X�X=vL��<���ׁ��v
͈cA2W^�뜳.d���ua}x��Y�)�"f�;�������o0 u,�&W������NN�ddf���6����=}~�܊���mus�d�Ϸ���a�Oϓ#v<��f��׌�T�.�;��h��N�������mm�$��"g�-�z;u�d���w��p7� v ���೫�y���{cL�A�˥披�/#-���)�H�DU4���1����ȴR�X��`���/�'��G�7w��J���df�WX�m��.�Lҵ����"2NKfC*�XK�\��}V���\S�Ri��xMf͚�[F���_�7����xmO;�k:�=�=\�	J�{�k�f��Kb`wg��T!�o]ߨi�ț�~�V<uNl;�h��^��ky-����4wo!?0�����M���b��4��d���x/0�>Jɣ��X�wX�}�ie��m������a����O�{���fsy�a���� ��'dD7��f����9�S�r/��nHw}*� ݪs�J��v  ��"wA�U��dC!*X��V�L:WdӸ
��8��ݸ�5wkN�1gV�]��T1k��m%nX���Hم�ˢؘEp]�c�u��!6��w�y�o7�y���t�G?yk�6݂|����0��2�?�4�p���&:qĦ�b�Y$��[O��zH�j~�d���Pfϱ�^��a�⤉}y
�!I'$F���͈�n��Hϳ� =>ggmq��>7v�uζ��M���a���r(���?a==:��ߩ�z�5��qn���ieF�5�8n���>mE5����>�֕�Q�&�۷���K���)��>-��j��F�u����
]��X�1�#X���Խa�f&�Z���ca�������'��X��<F���19��Ҧ	��
%�KI�T�T{!����x(��\�ZQ���Yr�a{�$�+���+Q�Ѕ�]��/�#3�!j��)53�=���7�y�9ln���@fÚ���z`-����>�u�o
�%�U$�����o�����G� �
���P���?�DC��*����U �� P8;��{A���s���p;@3�.A�8v�L�CBF���`�
����b��	��A�
D"��d*����,BF*��FA��BF(�d��c�@d`1��b����dd W.v�9���r8�� ��B ��F`���0`����(1��@b�� �A��d���BF"	��$ �"@`��$(��`�A��BF ���$b��$B1�$"�
D$`� b	�$ ��"0�@`��� �d!�@Ɍ!�����$ ��F1@b	�� ��@D$b��$ �
@b!La����&0��0�H 1D��RH `1D��R��t�RQ 1�� H 0P��B HD 0@��Rd�!���C02D 0D�� H 1��B  1@��BD 1��HD 0�1�� 1P�� H 0�� �BP 0P��B 0@��D 0P�� H 0@��W� `�"�`"���#�0���������F0�@b� �@b��@`� �@b�
�n`(�@b�*�@b( @`�  @b�
�@`�`�l �q�6�g(������@b	�$(��$
�FD 	�$*�)�`C&0�v�h��`L�q��� 1��B!#H��T"0D��r2!H��H�0cH2#"�0�E"1��0D�W��[l88�r�a3�� 86r�r�m�#�ɰv@,��9�Cl�L0�� ��u���;���
"+*$b����_?���y�p����Ρ������������0�/�L��?��{�w���?x� ��O������Az�"( ���?�D t:~������B�( *��������щ�A��'�����	�������$���* �� $ ��P����B
E @"@ D
A$E", " �!HH	H����D�� H�H @B ," �B+ H#H0�AB) H�$!HT"�(@D Q!"0�BH�� �0� H1��	�BE�	BA$$T#	B@I H�EU$@�@EREA��**)�(�"��!"(D(P0��.0#��
`�&0���GCg&����D 	 �b� ��$"X�E�$F ��A�Ab!��E�$P��D������p?����)�����(H ��3�@��~����B@�� �h�����@^��~�ϣ��~��S|�t��`o�!���:?B}� 
�?$?�??�?B|� �Р ����D����"�����@_ �q?O�'�����G�C����s���9�N0 Y���?������T X~eO�g ���;<��7�?Po�? ��>�'��h�<�$T i��p���� _�]��~g�v'}?4���8'�p?�����;�I���Ҡ ��v@�~?�8����~_ `���~�%�A��8oZ("����M������i���
�2�ͭ��x�������9�>�(���|T}��Z[J���Tfm��;\�N�خ�˶�颣�u�t�b�Q�Sv��T���gu��;��j�������v�3X�f����mj�f�k][wZ�-����hwwn�]��7s��U-4�ì5�6^�sݺ,F4mb�Y5YC6�j���.8I�Ҏ��*�gji�������s�)�j��[lV�|��ں��Jt8���u
�v���Jգ]�R��m�����s�s�+Z�� �6w�i��cQk����B����7s�뚖��ٳ��fRhkgm�������� �  gw���흧f��k����T�m�5���zn�ݹY�u�{޻o%��u��T��׽��j����T��㴣[����m��v�{ݩ+�v�lܜ��W�=C��W�ݳ]��nU�x�czt]hl�m�]uv6��  w8�
(}
:i}�z^�D�(P��(�=�"E��������W�)�������{ۮ�n�gm�wzv[^��v��Z�n�׷w������m����Yz����r����׵�t�n���dm�䔻���j+5|   ��ݽ��m���뽽N��i�w-�ݮ�^��U���nj���J
�W:�N�ڽs�[���1w�G{������s�V�m���h4��wu��h��ƹ���  ���3���mlݻrw[p^��W�����*���{c�F�[�j��n���ŷ\;P���Z5M��{k��F�w�
m��
�۷Z�kfԖ��|   ��}'�A��t��]R�L�ѣj�K���F����8V�kl�X�u�9k��wu���]k�ٽ�wZ=k�I��u���µ���[VY)�Iw;�   u��b���gil�ug��M�:���5��7Ev��amz;�T;`�3�  <ݶ您�ܮ�hj��W� ;:�[[[l��{g0�lj٩|   wu�� Q3�:H��0 �{��
Z�.� �X Qaw("�מ׀�@'rn:4 	����*�={Z�3m��W���Պ��  >O��W�� �ήC@;u7Ҁ�� �T�Ӱ��A֔�ٸ )*Z�p�@��� iN��e6�P��j)l���Ƶ�   -�΀�Jf�[� X4 �e�iJ�����  .�{�  �\� ��pt Y˹JC��g:�n� 7�]�Iʨ٥d�Ղ�J�;�  ��Ͻ�Ani�h R��{�)B�=�(W{��� 8�(((zoS�� ;n��ʲ��{r����� D�%*H� h�"�ф��Bb 44Odɤ�T� *�4��@  T��MJU@ e*	�� h f��G������_ۂ�����n,�g9jEm���L�V��,�AͨA��%���Y����￾|���c�{� �����6����m��c�; ffo{ͧ���v�~>i��_�ͦ07^�Lꛀ�@���)�.����Pm�V��2@-ᱬ[ӑ�Y�o	���*oiR��.��I��r����
]d)�*�U����o��m��r�B�3��ц�4����lլ�K7�!R96lW�v�Qr�8�`���F�|[1E�C�@[�R�s��k�Dͽ9�wsi@.l{��K&�uj���bj�t����.k�wL�R��n�6IR��h�v�zF�
;�J�?m^�3 b�oq<DJ:v��jX(�B��=�eF�
Y��։�9HԽ�I)nڲ�a� 0�WI]^��neenb���@E(���T�Wt�_d����I���S��Ɗy u�XE��e�Nj�j;If��W�S3n���A�U����Cm�HB�
�wv�vn��^8Dl�%�H�U��-�^;zBD�J<��bK	��C��{eP�,���嵒�"F�V�N��UK�����1�f �Li~fٕ��-�g\	T0�P�l|3CP��v�S��E�l6([���Ecְ����̚t�K�!tF76]�Y!�[9ۈ�c4i��^n���b�2�����״[2��ԕ���ݣ���T��"�VU�V�T�ܺ9�+O�)Ru��7tV�B\��6�:J+n�*2^Ԑ���.F�ۥ["�&Yd��E�-[�X5�fɇQ��U�f	L]����;1�B�Shв�ɪ�br��^�u6FS�<uT�%���n�l˥w��^� ����Yz^4�Na;j3�j�^^�T�^b�kspeѽw-c��b��M'r��[����"��m܊�4ˬi]�ݔB�n��k��2�LQFh* ڨJ:�YmլS7k"HཇnS:�m��%��ef�I�%s!��:HoB�10�:�j΅3h ��2�r�Z�����{�Ǭc�1Ò��N�RB/Y��U��75�X`�6Ѽ�(P����o,2Ċ����CZ�P�A�k-@hH-�E���Us&�Ȍ�ف6v�U�l �٩�w�Vɭxh%wt,�G�q���e�jYl�f��T�K����Mڸe=�*�JD���GB�Cy��ɶ	h�h�]�� ������/��k M�N�e���(cu�o�ϖ�#��5b�b�	���;g�r���;E: �{iШ/�ņc��Q�0��W��W��-Z��t�k�Q"�)�dَ7q���p��.���°Vn�ǎ\Ԍ� ��8�R���pS�v*aH�y�kz�в�\�L1V��Pdk&���{6�Y{V*i�[��q��xՈYC�Rji_٘�ܶ�T�*�i"���&"���R�����!��	���ۗ2n����t��1�R7� N#�+ه_�T)�L�(�o.�,�RwkjB�!���b�-���v�"q�4�2����u)�׈��4b����ˉ,�VJ�^�P�l���m�#%)R���Љ���v!�E� ��N�&R�0�[������S�������wm�6�H
���H����-Ņ9g
�f��E#k9P{[b����8�4ay���M�n^RLh5�3X��-�L�{�عD��"�H��p�`-I��杋tҰoJ�,��Z@�ۥ����쳺�O%R��i���MK2�f���om!��o&֊��SW�8� J:�N�L���2��m=�k��];r�4ֻy�!4d��M<�S"k���4m��"ñJ��H�-{
&�GGj�2֯m�c#�$t��Bk,�X�q3I���J���f��6f RŘx�Bɽ˥�k��]�I^f2�g�-������[C-�@5vb��u�ڱCr��A�h%R����dB���SU�*G�m;3�}��l����YOn�r���VAim<ԡ��W,�T��raKⅲE��)�eU��#P��E���$�%�m%F��-��KcR�iv�Μi��#N�YG0:�P�e�uXh���PUƋ�X4F޻��v���n����^
��d�&T�'M<�Z��{uf��7�4�x9l:)3xe���aa�6�A��kjXͤje-��<E�5�I.���6Mc�u0�ք.�Xt��Cn�����Ϟ 啦��Q��d��M4�Y��*i���U;R��yWb�N�d�p��/ (�i֭�īr6jXԲ������P*�kߦ/��
��V�L�+[h4�U��چ�$�űS�,Z��l��TuP������]l;��N[�F��2��T#%��Wp��f�՛��/t��"�A�� 
P�W �Su�����=&���'�X���@8����H�/E'7(�	��#HI���|+v�2u��=��o-)EV���Ͳ����Bd��#M^-��Yu�c���&��`��n�zYe��a��]K���uvԧ��f;d�vn����f�m�W.�R�3����gK1�9�{�n�0�V��:E\�&��t��tUjʴ͔�RJʂ�n�J�[.��Ncrť5�����˺5gn����6橴��X����! �Q
oqӸ�be?���6�Y�-�[@�NS�U@g�,�{R�֪�1ۻ���ˢ�]�H���tq�W�n�ER�4ۗ�qkQ-�*�$��jQ��fmfƢ��yR�RGm�Y�K�&����^�w^��u�B�EL�/K�KN�CY���|sS�]3u����8R��l�H��x2�t��޻�������W[�^�iH3*��F�n�V-�~R[Sn��^�])��N���+1��\�{N"��[���D�v;�v~tbv�H� ԩ���N����eM�N��ۦ��t�n���P4e�u�L�l�2�t�/\�3b�GH�0S6c�n�5-Z¤E�2_��b�v�[�>n�MnͧE�s��h�U�����z[OdPlem[z�5nMa��t�ck\R�V��qP�,ڂٵ1�Z��z�[[�����Z֍��Z��x�5�R˱MM�30CI�MZ׏$z��-����x���
'\�B�an�`@�8N������CW2ûQ<��f�A��e]Ez�yn�kbɷe��3m!J�4p�q2�a�xfc/i�):
*t%��h-�]��S�YW�7h;մ�@�h�u���Vmm��L��[�@VP�m�sA�j���7�T�}m���5��J��*f��hΚ�`TV�N�f�V��p��.���ǚPV0�m`p���v�꣙.��VS
�b�F��^��Q��kP�Z�۠�qL����l��C�ѻ�#[z>ƪ�+j��U��pa��E���ޮi*�-%����V5T�j�	(-��zػ ZYWn"�Y.�ei������h��jTMB~�Z���g�͙x1'x�+�F�7oQ�Dh�M�q+�y�[�z4�˭nmK���>�Vba`5t�J��n�)��Z��X�,2�|t�H�l�p�.�Ke	��z�v�wN�c)���l��He�4������n�����Ҩ���ۛ/d*nn�۽o�# �٤�D�Qb^R��:�����^]flg[�b*2��z�� �z�@���[�%NdEࡐ,�	J�=��彷��r��$ҵ�[q<ċ���ot6���L#ޙ�Z��I4An��)������ӳ�v��l�%�L�:L˥�ܢ�Tɣv�j�ݒ�H븕�ި��r�	yM��)�+�n�7���e�K�e�/K�zHJ���ڳ�,O��&ɤ^
ʼ�
����)�ډ�sf�N�BR,SC
��s���կ�_L�����ԅn�'�c�\��$f��@!r�ov�X���t䩚5�Y{�e
�f���Ԏ���ܭ�Π!�֘6hAe�gb�1լ�H�8�s.�i���I�Ӧ�Z��Y�vBb�1�n#)i���ݏT�WX�"S�m��,�T�ƪ���~[N�0P.�wwI
�Tbl����^cQ nGF�c��DíTqJq�[I	4�ȵ6��HSj^)2t�X�IR�@\S��hCl9��@�y)R��� �7e����(�Ճ5�r�ėV ַ�		,U�nS�ӢHL�ٗ����ξ���mZI,�h�	<Y���i�Ű4]Lb��-M�ܳYbF�K�6�mf�|:GJT�n�NSѝ���-��\E1#N�n��	��Q�V.���f-z�]K�a��)z遑IH��`dRid��M`����j�!@@]���֓ݦ����{��H��Ě:��mkGq6�����W,�H⽥ύ��#z賴����iyx��-V�s^��r�c��������c�4��A���Q��� ���5(�[i�I��=�7V�sxim[��g>���l/m3�����`i�q#�n�g;��p-6�֞@4��e˻an1�5VP8si�F�(��e���s\zi����0XfSM�*�Õ�f��րs�S+�T��9�5(��!m[�8� ��eOڰ�4�˱z���pU��xK��:�����qSN��hr��٬��l��x��QG�fO��ڥaM�(�R��X�ᠬ�f��
�ܫ��r��:�#�@ؑ���-סHQ&Tn����R�)P#�m%S+fXԦ�M�.�`�)1�%B
��ؠ��P�wYN��IE�Ud#b��n�D��zAL�[���ӧp�M��W%�x�2,Ä�Qj�K׺�,�JeJ���A���1Q�$I5wK+v��6�3	�>4��#5�e{j*�@��������`;��-�`��V�Xx��i�u����v��&�u5��,܈n\2�6ޭ�W�M�t)=��{�)b�aXݺܫ"�#5:6�M��\�n��ei�T��\B�vP{��eX�J
�Q�*Ҩ�h��WI��N�&��a���[� %����5{�(�[�i�4�&��M�:�K/�{W��f�c5�Z8�%�/kL�AC%U��	N;Z��I��
�
Ȭ(Fi�KA������aJd�P��g2����� w3*h4���V�,V0P��2�6�ZԽe�Y�)�v۬��#z��q8ۚ�J�3� ۔��3V���Ͷ�Z�ìg]�{�F��LV���!j�v'����V�i�2�4:
klqn4լ/mYƱ�:���.���Y)lgRe�$F-0\Vժ�G^^�I���wq�BXeK3mU�ڔ\T�m�l�0�0طK.@��`��8�i�*3��A'�j{����� �me�^V͵��aT�,P�U)��l�Z�T��$�ł�&+Ѻn��kt�8�)+��V��R�#�ܺ��((�n�N�	p��7�[X�	��41���KM�u���62�w7v��뀸0A	�v�l�Ѭz]F�g���4�7���q����-��Ȋ�pYj�!�;����n�+i�ނ�ZՖ�d���5E@�(HT4��'*�E��n���Ֆ��GUf�t촨e��n��:4lm��ѭ6wb��K;���!�ww*mD�F�^=�Bɯ]�-�x��k�WNň�a�mJ�q�Q_^�Jn�g^5al�#gB;kH,E����u����Ȕ�z䗹�-�He�Zޠ�Ue��&ѵ�VUr�t��l�f4-�m��sb
ܺ�pZ\�I5B�+c�BRs7Fǭj�
��$�9���.��^Pٔ�
�Bf�ƪg-�.�T8pFv�F���/1�g�@�%��Ѻ8u�Q�E[,c/e$.�Ԃ�Mel�Cr�T�1vq9B�̠�ZI�	��K�SUel�LL�;��" �b�+$GV �,JC����.���'u`m�Y�u��#F�ؤ(�Ͱ�Cu�Ἰr�-1S�e|l���:�m��[�yM�[@�t墅�U�1�� %�9��9L�̩F�����A��e[�+l6j]��+,Z�[W,���a���2�Tp��IT�Zj�(*Ք[�<�,Mz�=�P�&U��:���v�M�g�D�Y.�c7�Fl
Ӹ
G	6�=a�$�*��1���/V�Bf=@�q��mۄ�J��&�T��ۺkoLݭUv����CJ���1XZ�sd��M�y4ݦ�D�Z2Ep��6r���v��'N�ZoN6�vs�fL�"�	U��["\�uwA�&�%m;�� z�80iJ�b8ܳ�ve�BZP'42�Ϟ]:�E�$<�{�wc�hEI+���Щ$��5d�*7I�����R�(���XMb�6�*�cu�u ֕u+���·#��×���E�W�^����,O#wE虃5�����Q�m�@<�96�?0��=�!�ѓb�����鹙M���62M;�%��9[���Y�Lzb$�d��֚ke�q�`��j&�)
��M�n����
�� &����� "�A,���H�m���ZE�/D��qV����|y��,A���r�ֺ/�:�@�� �Q@k3j�&�S�+�9�ش�m�Xu�p�n��Yd3����n���-�ڷU��,��Y������Zk	[[M|j��fQ�n�*N�{���|���F$m"����Ɵ��X�����oٸ)��`q��E�U/]�͈�*�խb��MY�ڊ��]cCb� խ6��,���؅^�a��J�����hQ(ѤZ�&ȡN��e}i�'joi8��&��q֐4�y/hn�5��L܀��B�b��f7oe]��|6�l���j�R��Vqws����Yu�S�� � ͽ�)�R�;y����=q�3�[a�E��*3%3�����;UsV�h	>����d�i�dlmL�tӘr�95 �A�;[���j�n�ckS�o
����R��m뗁��o*>;�:wT;�8g����6M�V��A�-���$�98�c��V+]�n k��d�x��y�����gL��ѷ7���S����J�N�zNʰ���s��z�!w�\��K)s*߹���
���+0Ol��i�����&:���Ô�X)���΃o�z�l����#��m��ky����q��H�"E�������թ�d����p�$z�Y����z�ӗ��a�⣮_c��"��OM.�]j �vJ�3c��5{D��6�غ	�t��ڼ��\��i��d6i�Z�Q�z�!+K�bȻ��<R���1M5���'f�ߎ�D���c�uۂǫ��K���r�Q��0���gH�1��{��*�^�/��@���0�Ͱ���m��}8�b��GG��a�Z��e
WXMp�A9*�����oZY9�=$�5����H[Lknr��f)�z�]�m�S��,w��5g���:9����1�u�d�ޜ�䫖�����	�i��:����v�WN�6@S�c�vudu�csv���Z���]�i�fp���r���40N�� v9���#!��-E*\��)n�����Q��I��8�A�?��2�����ZN�yn�Ȏ|0�r	�L�6��J᧥�R�d�
���
a�K��EVŽws7���0!����NvL3�9�\BԮ�80���n2p�T�0R=����:�74�{}W���I^_�fx�T$[�O���(�V;!bή]�v����K�I^Ƅ<�r�p���v*�ђrS&f�qu-�5�ZάqL�x�]֍�,�{OC5�E��Yԩ�{5t�tO�U�1�-V)j	�����·iq�/-�7C}�ϖSɻf��l�2p�;p0F�;(��ȁ�tJCu9����A����lC�e�۲���	[I���e ɓ(1�2�Hgs�Fb���
�
�$�Nb��Z:P�U�!��U�_-Kfd�dX+���Z���z@tq�nS�ⴸv��#�ѥn!�Ne]�(��K�6�����F��17�Y�<\(r�wm¬pWI�����6��U��Z���,�V�����y�:R��il3�ؽ�N����)�(u��\�c�i������-#]����aCEYsx���V�`�u����V"���/�n��Ko;���	�P�8�L3)��-ˬӤ�p�me=Odt�E��h`�r�Ƭ)��n��S�c]�ˆ}�3����^�g
W�9�:΅"Ӯ����&�#��q�xG2�=��0<��'F�v���S�ˊ��v�z��}|�#V�f!���U��=ܛAȮV����h{�P�Y��֯)�"��Mf���n���V��CsN>A٨�=Յ�tK�:��ު;-��M�W:������uI�xR��*E�j�}�")���n� S�/�)OfX������U�.�6���d�\�n�*[{ǁ�+��$ܤ���4����YݨwW>mLw�۵ZOj�|��u��pΓ����x�5-� Q��M��)�w�E\�$���yy��'��N��N�s�QQe^T�}S"'&�t�ࡵ�d�ڦWU�ꙮ�5x��{}�p�tz]Xս"p�:��pQ�@�]���ѱol����kW ����6JL�}�j�wsfti�����Z��{��/��$�qy�h.N� ����z��N�˻v�0U3'�m�}��'l���Qb�@�N�)$�o� YwI�0�F<<���7-�p���ǧ�^A,ͦ���mmi9��n�ٖ���[@�up0[wb�%k=�nV�M���Rp5��uxy���k�_�8R�����s搢��2�h���G�8(k�;a�J���0]�՝��z(����z��❎"	�MK�{��c�Nݜ��xA/��ݔζ���Y:l]I��g�ХwU���dd��aP��5%Ձ�Y�с�� i��$�{3;�̾�����è4���q��(�'_Iӷo#��gh�Y��G�U�ą�5�e�E�n��@�{ҕ���������s!9
׆�4-�Yf��<$���:ʫ�?&�ձqΫ�R�v�*2�ث�w��s/ak�)Ζ�5M���<��Vc��;u�@�TƆ{J�ZU!7p��'8H�5	�*�`v945Y����ԫ(v�)f��u���C��۹��v e����%1LRj�^>�=/N.�뗚�&�|mv�<Kѽ�6��r���K�]���>��.��^����p3֚��I3r��^�}���*�۫KVi�ʵ��5��>ZOb�թ ���G��XK�#c��sn wɣ�m�w7�]��ص�9ŵ�}��I��=�7��#���}A;��(���fb���	T��
�5֍�$�,��Q2�O�0:5׻Q�F����E.��Ra�t`㱜[}�+�"�U5��HMT�V�W�Ge��]��-.�3��(m���a<�$�Z޵i�҇�m��%��yL=��z�Wj踅(MnO��H�����v�
f�i��;h��6�j����Zur]��Ӄ�)����#l>`���L��ٳ8��K��c�(A����S����2���Z�s�,��3��},�}�)�D��soq':���a�M=+�,�X%��Y�0�*f��O���xɌ+.p��u����0_\�E���j���g�9���u�+�W
U���&�>����!'�0�g�Mn�3��O*��������(�'�t�|��[�V�Cչ#8ʺ�v7w���t���x��<h辍!�+Uݢ�{�4q�]���7t�`wI���r�Ӛ�ci]�M�ާ¸!Ԇ���؉A�Y�e�;0_mq��^:c�C��Q�4����;��7z�P!V�e+=\c�QV�Z�U���>�\��F�2����"�Mn�7�j["�y��.����w���Nӽ�*���06���@��wǯ;P��ܾ�t��d�K[���*q���}*Kkn�j����o�{r�Z8t�9��ڨ+�AJq��[h���4�s/�J����)Z�s��[� #tٳ݀-�X�����ǣ?����O���A`��}��[2��w0��� ��ֺ��W�J� �+^nι�i|�{H�|y"#�w��t�6u��e����a�_;��rï:ٚ���30m��(��௜�s�jÌ�IHe`�Q7u�Զp����87���Y��W5(�N>��;޶�߷Wom�Nj�.�.�X5�̮�W]�>�؎՗�o��T��oU˱��\ �h�|�n���(Ԧ�Lqr�$�����8l�iu��⯤�.�V9�7��s��@t5�b׼��[�;[���q�O��C��Wjٔ[g�+9q�:�f��Z=Յ^T;�yc�ڍέb��#��J[��yn��A�y��Q뙶��n1��LF�ն��;=1Φ���=�z�,;��୕�Sx�z���/��\OP��kE�M�P��n�]��ǳ�6Y.��u�3�uCX_kۄ�\���wo瓭k���a��y��
�I���$i:�8�F��������N��f�N��:uLAm�@�}��Y����R�!g���e:�����I�=o�Ôۧ�y�Up�31���J{�J��W��Bf�{�f�{�5�̻.��)v�������s���}փ:N�zx�NW�f^�o�5jYD�#lN��~{l�ne��RAv��g�'P3�!M�S�.���jp��
t�Wn�Ht�8��4�uFx��Jt�evTyO-Y���djҠE���ohє�!#f�Ǥ.|��'f�,��=�탎�c�/!�m�̚#�VJf�ػ�c_m�˼
��t]s t}�إI�7Yu�_,���\�m僭h��4u]J�� ���el�.�]^���j�"3'�v�G�i���3��ۖH�y���V�	��T5]�P�[�O����wO�V�K7lc[m�v��r�8h;�Y���:�+�K���9$��w�HG�>n�Aynt�+%\)K��IM���'*ێ��a.�Kyg��8n<u�9�EYѹ�-��b�n�W��f�։P4������ЃW*ض��;�b��}�{��o�[�lS�++3�x\�L|��TKg��E%T4�����h��膜Dg*ϐ�,&��:�wC�*��ؐ�z�a�p����Q�j�5	_-;:�g	��'V���g:nrg*�̉W*g`Z���5n��P��Q�इ?@P!��m�UyCC����<����г*�N�-Tgv���5Y�ʶz��m�)-+-+F�:���k��[�'36��1Ekj��8ФY�j�'�^���N��, �nf��w5Z H�z����7P�.vn7W���U��̣�K�Y��)t-��y��֖��/#�o,3q��V�����$�鋬}�CȥXާy��㔠6�u���}U�Ž��V���b�.��Ly�̢U(2��U����c�w���BjڛE���lk��x���&�i��NchO{3ӯ|<p��t$�>�N�f�6i��0�ވ)�=�5֧]I��z��6�a�c��N�RvPT�#v5��tGm�O�kZ�W����}ǥ��z@ʾxQ[X&Q��Y"��E�RS�����)��Ԟ�{{Pkۢ\W�<w�Z�V���
=�ٻ����C.���q:���,���^`R�6#��tSwR�ݥ�leΩ��wJ�!�I�\h�X;d�F��s$͘�a�apfF�o9�>)��Is�H�P	��	
��Jy]�b��<x��^<[ӧ=Tr�T�Wb�[C�Ht��4���
���\�W]��˩ܴP�91K2R)w���B��y��΂�mJ���K��bN�&���G�y���X޳�µ��� "�M:=l��Vm�r+��+s3`�9Up�z m�4 i��h�Yƞ
������w�ո����^D�P�J��n��.��8���3����"���f4M�b�s^iĳ�
�3H��P�h��5���X��̮p��8�N��N`N�}��t�G�l8�i�;�eN��eP9Ք�I�o;Y����J$�	X	j�
m������P"�v0wT��9Ү܋{u	OX���,�M�|�7:��r7\� �ʒ�ndV�9:]��W%&�Cs#E�3��J@�n
��$]�y�q��Y-�c��z1���0����k���cb�KV�|��FiB3����-��V�H`�5Ke��}x&p�Y���=Ԭ����E��M���k��\ġ@�!5��F�ѭcH�HF#H��͗�}��1"!�$� ���A��T�L�񍬳����OE��YG�m�g,u�\ލ]� u�8��#f���51�4X}����O�ܺr��Emr�c}u�`
�7�����yF5�ɨ�n���[j��j�~��<b�
��@m2r\q���
[���rߝ]%lT#;
O��%N�mJ�Fҏ{fu����pC�ǣgQ���=C��=s�$��$��y�`�
���p���'32�+k��/�t6�n��Ҩ�c:�5�q��&��ն/E)w8�o��JƱJ���<���,*��2j>X�q쎡ǆ����/m����������N�L�ڜ�m�	��eXwў�ܵ�K94V�꛵�C:�4x9�ȵ�����\*�nvcJ�
ˣ�P�I�k�(qq R��]�;�݉8��¹��:��S�6�񓳮�(����ECN���ۏ����]h�<K�;��"m�7y�h�Ӓ?4�
���x��@Mm��|G�ݕ�&�|��G0��%s�w����o�3��.�{(QUт �T]x�%ҏ�.�!eWd�o���Q�.i��l[x�.�H�s U�v�v���OF)���W�3g!P��j�pz�4E<c{�1�c2b{l�eQ��n}ۖ��]��\g��j環�twx[�ܐ�Y�xN����﹫�BZ�C��i�����wjÎ�lo���LpGDKw�V2�b[��V�;u�yqͪ��׊�iܼ^�8
r�ݹ�)CV���9��q�J�H����� �E�8,�;���2�����k�t.#M��c��B5��5��r��"oɓ��
�v��$�֐5��Ah5�k��h�ei�Y�>v���jq�c��x)���HF��_y.�����θ�j�n��]�o_�gn���-v*V�"��w�UL�I��L�z��E� �3m�Y�]og.*t<8��*r�_.�B�o�>��0{���p�md{d��\��8��MBU6���������KxU^�Ĵ�@.R[C9���y����A����R��|7�}N�y�\�\!�\Sk)"/�t�Ӕ�8e�{uّ���u�t2��/���qQ=�>�3+8��vݽީ�I��k�Z�y��`�]%�=��Q�Fs��uq��m)Zw��k�<��;y�|���cd�����]y��7Zޠ:6�i���*���f���VЛFu��c�L#���1|L`i�me�݌r��,��4�5ӝ�	���g2�������&��;N���sl��>p�C�e9-ݧ�ᆋ�̮�^�;sQR�A�(��;6x3�����[��,L%@7�Q8���Z��%z��[CH���Iݍ��L�̡Û뙁�+k	�`�l�tYh�<�Y�t�f��X�a�[\��foWt;+{��N�i��� �yd��o"�l�\�]���ʔ�g��L���n��NY�+Rgd�k��b��=Y�z�ukr�7�θ�2� Msy���ӗ��m[5��KW�L(Nc�a��n�4�̈́�U�HY�]Z]��$}WK��A�jP�М�9��v�t���K�j��r"J�*Wr��.��}�pM�d��o�v��:��a��s��ù���������>>}��` 0��m��661��ޯ���]�ώ<u����ϋ�h �ei�<�n�o׏��]��A��H^�� gL�ub��7ϴs���2�� �����f�&�S��vCN��a���JWg���$�U�.��s:��n����"�}�o���������Q%��C�OUŕ��<��>,#[�^�����Rk=j�C���U�(��)�v�9Wc���7��l���s���]Ղn��3�I����,1ؤ �;�"ٳ�A��8�]�%Z�3A��͎>�=�Y#Lڡ5Z����SER	�l�S%��\���n�5��T�`�ǉ���7#�	A���u"�yW�jTr��+�xf����o6SGec��ca�I,�ŭ��q;�ge)&G��r�,F��M�;v�H��Ju�1u�}�5�M�BR�xw�Q��$�x$�����8�5y`בf��FU7�s?���z�t�vt�U�.���%��0D�Hݩ\5Qt83Yb��*����{ӵ�z�Ҿ�}%EX^&�u���(�xxp��b�c��^Y��+a�ޥ�Xkc���31^S�[jSD�ۥ��;SJj����T;����c�f���S��P@e��ɸ���B��
�W�Jw�I�&oX �na׳i�M�j�e�;1%�4z��$\��vPNV�; �K�����.��n]�]����ݸ7�&y��5�8�-+_ًZ���"�,З�$:ݝֹ*c �yL�S=�V�i�m�m�H�3t�f��BV"Ԓ�Ѫ� �6M��̃^��a�`�kr�t�k���n�؄4�fj���,�q��)�:bw3�u탓KW9�Ś{T��X�!��
�*]m۵	�_,N��x��	i���)_AV������CF���aw��w�\���Йt�}�p�[˹ C����.�;a�EP�vY��a���՝�P�z�TK��29���YN��j��JQ��-Kz�:��py���.�Ya�	&o[M`A[�{�̋j�ޜ�]/�N�������"����X�jV_6�
�����I�M,.�K)^*�\�p�C��P��"[��1��.���8J[��,�v�Ue5��oZ(��'+��-;��Ϟ�3�D�>��#nJvjƴz M�ڎJ9�����{/��q%�ܓc��
:v�ۂ��r���K���kV�_0@��ƅZ��h �`ea�6Ġ*
_�\�����bo���2��O���9����m��L��Ju�d9v�>���ump�M|�jg;�)�V+� �.eu���N��u�зB��${�k �C�,��l议�w���К���[��k.��\×� �u��F�y#a�	W�v�(�/Y��l[��U�䪂����㛂Vƃ�/4M���8�R�4��.�U��2䣂�|��Io��,���h|���OuU�#.��'��9��v.�`�s�@�ح�D� u]X�4S�&=�"���eX8x��2�\�d�N�V�Ėꔬ�K��<ɵf9M�;j8��#2����y-�YK���#*!ٝ���zWq��hq�h����q�������0�s�$�]�[����̔݊�2�;V���Vx�{���J��iG�γ�k�A��y�M8�k����>Fb&���ۉ��-��z�*���-��K@]�A��شm�0�����ݭ��)�T8�+����(�������WZl�7��]��kW�{^9O��ʖ���]�hs�I�`��s1�[�8q�h�!�Y��ۃ
-=I�E7����
t�'sM3ۛ�-�m�Ƕ;gz����Z/�u�9�P�ɪY7C�.�[JPqՍY�G�k��Zp�$��;�F��.�gZm�9�-��t��W���໫������ȼkN�=�T[Y ӳ1-_D]�5Sw#eK�x7���R��	�^�-��Q���Mn���֭���uӦ<��1�����2X4dG,@�h/���i�u�[��\��[�Hg.�vS��VF"�1���JC�,��F�t1��8k?���R��}�Y�v�1ݽ�ЕtV�Y/iYۡl�5݋wc�+���teA��C�)���1���5{�m����%a�ʋ�]�:���vX/�z�]q���]iu%�՝q�2�t,
�uo��h@�;"D���<.ɬ����l_�(ۮ��x�ʀƸp�'�Q�Ҷi$�eZv��w�Ѡ�Vin�w�e��q jS.��u���k�jQ��u�m��.��J�0*'r�=�Y*V�o\Ǫwve�a�vM��v���I�u˻��u̍|���%��8m�]����Tp<��6:P�z���Ok��\[dp.ua�9)��i�8n�H�eI�R�޷�B����,�A�M��{i�a����]�w�̱[�<����^�g���·��=��6Lf1{xa[,�{���b�K-�XJc0�k5]QWqCX4|N��F�i�]�g�R�o;{��W�pL=�#:*�a�(��:���6
{)��)��Π:�D#qe�1��iGg��N�3ӂ�r�|��]u��GE�*��ܴt�Jz)��OB���4n_j��*��r��=�Ҙh�O��7EP�=���EU����X��n�W�GU�Vi�d�#��G�tW��]Zg�qo�S�9�
Xsw�j�oK1��ȥ�I��P$]j�8��]UQ*�k�%G*�c2�E$��%[��>F��!�Az��<s0
y-0��qͻ������K�D�ҵR�y�d�z���;�q�*pd3.ٖ_��Xl��"���\;K4���Y}�tA�Vv��*�j�z�k�3����鐵�{����`Zoh-��{ٍQY�_:����n�h���%^�P���ThWm)N+r>ڙd�م���ր�ӽ�l�=�&a�*�м��rȻ¨+��1\k=�+���D��f�}RC�W\�80��1/�4�B��)�J�opU���{u�W���8�O����\o���,�:�$\t���go��Ս�ݼ���L/�R����J`�!w��<�)@ݶ�=�W��
q�֤�1!�|$�v.��N���O,��^͝60�f��v>3hN�i�]G0�m�LnFi
��44�P;{}�ߛ[]�z����I�Q�·����]qn7-� �a�i�ث�*:_�\}N-��0P��H�&u�4�����]4���P�l@�Q��T�gy��N��h�z�K��'��#���If���";�IK��o.��0���]��g�ek��w�;����b���p���du�co��B����bJ5cQ�%��y�K����3vgg,7��gG�Z��Rf�0tKl��ۙ��E�˃b�p�9ϝef*[��j�7)]
�@|tvIK+�ŝ�F��^���]`�Vk���EDX�@ld�S�ٻP����]�-�D܉ݽ�q����˔��e'��A����=�3,�;/��G��f��8�8^�Դ�$*�=�d*�[ԢK�$zͮ�!ڦB+�d��'��V-Ǣa}�m'b��8mVC���,:,�p�.E�r��-�)u�����wIu�]A��w������o�_$��u0me�#�`Si9[�1e�e�_� �;et"�X�L����KJ�E`W��P9�ۼ�W$�<ΐ)��V�.��>N���g�6�g��v��ֲ�^E�vnda1��<=kQq�� ��;���P����S��Sz�ٮ�� ��Wc�&i��G�[�ݚ*���z����M�ϛ��Ƌ+)�|%��/Vts��E@Gv�����q��rT�t����ݺ���0Xӽ��fF֮�@��2
i�M�p+ƺ��Ĵs�'u�P����&��6
��N�����Y�{%���n=.������F�qM��`�oI`=��y���n�7;fRgj�:NM�Y���Y��op=���wu/[�&n�N�{���I���T>���SrQȺo��g^���]�J��.�1�V��˦Ţ�..�\+�FQ�F4�i��<�"'�B��*ZS	���b�(sQ�����ˡ� k��R��H�w4�qj�}kI�Dh��������y��+O(�P#�;�q��`i��x2���h���L��7�v�a��q�f�d�{���\li�9X��b�����z%ۻֲ&�<E3��g��
}@B{�\1f�J�i���]Z����4qЄ�u�QJn�ڬ��/o!�����F�wz�sW;6i�uґ�S,�Т��Gq�]��]}��n;މX}��Ok��g"�W3E��������Z���|�D3��]u�HՊsH���͕�!���:�[��k%褛��XK;Y��� �X�o3Ww�CO^�oh����{���@��y���G`q��61��dth�q��.N
S���d(�"G�Z��ݹaQ{����>�;nӥ�IȮ���ڄ�*ign��t7� �G�wt㬭�}OOn���KvҖF�Qkx]�X����xh�Tts���>��2�W7�ָ�[�];m��[�4-�[P
�j�]�_r�:B;�+��Ǽ]N|�����a�WP�P�tL[�z���/�I��#:�������B�b���9
�l����@�5��*{P5c��ZT�"5Y�3��� (�Hc�����t4/z��0"���VZ���eq\�MN`�ǭ�5b����:T�V-�7��x����J��ٻo�.�0/^:g��qr�*q�pֆ��Td�W��i>�Ef��K�<�oA<�l|�ټ��w,��K��	�� ��kkN-���h���뽭j��� �r=��Wrn������YiJ
#W�`É�(��!��u�'�
k�R��o��Q�Ka���^S,KU��/��(ne�8U�Ԭ�}ώ6mq󑉘�%ⴰM#��
AP��Nss�	L��͗wƌ���	2���K4w9��q��[a�9>Ѩ݀z0x�N��܍R���3y�%kf�;���Wtދ/��.���ii�"8��;}��Un�*�b#�4����m]�Y7@8a�z���N�p3˷+�gp��f���|h��vI�X�m�XT��!C6��f:��vFs�/��f|k�-We�'����s��.elV�]5���W�f��]l���(�|��C���gPDb�:TM��t�X�j7�I�J�B��0:��;j�U��K;J����BR;���
��=BNqL�h����ȏ7�Y�`��o&3�:{�Z�ޞ���x�+1��*uX�z��6�*�S�Б�+��Rp}����In\����
ӊ=}���ی꾩i�/h�y�V�w9���u��ٴ��a�!-����.K5���t/Y$���!��"�rg�m����Fu�=�c�X��ɮO)���`E��M;/��Ѵ6�X���i'��:���6#���7���ow�bU҉��o�1U�̩̳n®��i���R��=��]0�N.6�F�s��$�YV�p�ۢ��\��� -���ۡLp�-�������D�fs\M�˧�7u]�WEs����9�D(GV���yO9OD�y�"\�;|5h�(�o^�ť���o��e��86�����\��6���X��C��^��ު�D�"�حͬ�|�pV��M���q�,�v�k K2�5v�e�}J�櫆��%�^�GWحk�凹:9������V!�B�*�*�ѻ�U�_)��<��Z̆��h���t��И��y�n�C�k� }��<�>�YY���U�� :���R��B�R[�����jr�[R�Z���1 	�ھG6��ε�X�tk[w7CX�^;�i9wk�J�/{ki�X������=�-��=�\s�tq>}�N�	Y����U�5�E��H��!i������g���ηG�+.:�{�Vn�δH����J���(�5/q'*�Ĵ>���t��E3G1?�����r��e�g�i�'��6��}�Ce3����ۤ S��o,|%I���uQ�rĔ�kG�̂�nӗ�f�#6������l�:B��fT�Ye*�T�m[�͡�A��ОI���Ǧ���6�u�1\�쭼z	�V�UƐmwp<Jޞ�GV]e��ssJ�}j#�ȼA�m)ԯaޜ��4>�T�l��/r���p7`�p����s���N�G�Yur�6NT������˛��^P��o=���hU�"T�z���Z���j�~Ї>���K�:H�qhM�yqgtov�����.��q��1�p\��D�]�毁��2r�u�%��v�9qļi=Rc�pK_�����J�|���;B`��Mm�נ����J\pc6��,���d���f�ج׬�0"'[��ug!��V՗��i�u�j���yɇ[�w",�\�D4QBjv���wz��PWy�)7P;Y�i�>���җ|Ihon$���^Ϋ�Nf2�c���E��uf�@�ߡ����m�Ke�Y� �M��}��\����,��g��#�A���{�a�fZ�Ƴ��c5 SR���/GR��y�)���H���J�h�O�/3�1��lQpY�E]X��أn@�\S�4X��K�yJe��n�rlM�.>���t��1�`��9�n�"oQ�X%<M�h"��:��m����N������\г�]�ۧ���-4��:��w;�Z}��w�wlB�>.�ѶZur�k�T��a��)�2h{��a�}u������7��kf���gRk��fAx]VŶ�EI���n �ͤx�V]uiSj=bh��98;���ӓ���.M�E*ئ�j���X��pR\f����w}��D%Ň�D.�r�ڃ���tn}0>/1��ɥڭ��&z������oy���{�>�b�-�Z�"..�NmЪ3I�4:Kn2���W�]w.���'�gto[�1�U��$�$�6�{��=��ӻ�46�:i)�f��E�s�x/k���4M*�O%8�urv��G��V'�0���tn<� Y��NC�Q��m൲��� ��[F`5ڦh�;��	��u4latZ�]e� ,��
�U�E gs�"E��t.�e�lEMr�(R��uhIZ�]�t�vSX6�pn㕓!��M��cm��lҺ�εZӺ�.r��+y��+�;���es����4Ũ^��)�t�م��A˶s���-�����d=�Dy�՝�����q��ՅWc4ވ�J�<��B�[����:�[�D"�9��\ظV��O���?���_��5���z��6��GA(���"�	�^?�R�u6 �cme![�6z���&|霨E�iu��1��t�VѤkaknPO%���t(�m�6����	u�]�����q�:�S�(ު̭ѷ�6��U�z:���Ja�6,7��.7,[��B�uX;j��I�J6Ki*;� �գ2=��dɋ�޾��^ݥ&x��٦��	��v*eN��[�g/�����[Xy�L�����YQ���V�M����/Y[WOi� @i�C��W]�RfnP{v�_K�+�����T��l5��!���	7BSb��8�]b��g���R�I�J	I�U:��J!WIUdU�!u-	L���m4#H+*�$5*��,,����
��KD�jh�Z�*ŅsZ)�����b��,�����Q�+�
�L8��]2"Q�e�XAUGP�".V%�!���fCe�JH�*MR@֜�J�EfV��b��.�-JȊ��)�ʬ�'B�j�b!%1����GZ�16���Z�V�X�,Ke��heF����\N�"I�Y-�
�PPFU�Jm�Tp�.bauL4C����Bm �ZDd������(Р��K1$�%E,6V��HY�K�ȉ���%ed\��\N�A$ �WD21�o��_<,AK6�h���;��WY|,��ރw8�X霫\��h�P\WI���\ꃮl�_N�Cf<zb|�i��s��������H��?�f�Q�����O�:��������V`�B~˷އE'x�)�!d����D�9j�ڥ� W��M:���Z�z�#�!�a�::śDJ�Wz�ֽ��	�R�SXN��{͌��n�����߇eP���F��`1kl3ڽ�C�z���G'��
����!���-8��T�����<T����� R�v˾r�`���R�����*3��&>�g� ����Y���MQhQ(i�j�r��B$_��w�}ܽ'(�l��9����N*�:gbF���M�����U��A�N�s��y~�œ�]Ի�N-�a��R͞g���="��3=U���s8-���_��9 �Ns�e>~�nJ6�;7W1�7=7no�`e˞��Ϲ�\�`�>^��u\���z���݆�jV����ȃ��qHR��6�������e�����޵��֔P�뭤 �H�Nn�3r��Q.0�:|�Zl�V��� �[>;��F�=��|�x"�� �LP��3��:K/�֘z���f��F�	�{�{[�s���ܫ���Y�U��w�(rO�
�+m����9ƅ���b43LǸa�f�z=�c�(з��'\?.�f�b���o��:���zM��y��4�a:D�(r��#ET�cg4�f$ؓ��&�LCi#�K.�޼�*$g��������mz���ks���˹ח"T�~��jX�kN
wLᓻ�����R�r�d�z��5�ҝ�)h���&=�@����ڝힵ(��H�	�Q����@��Un��o�.8��w��h
�wS���P���Oް��}�;)���r�=���>փ�����>��W��Rmx�1_@�8���(]��b[-Ŭ��:v�{�UI����E94�tc���[i��^�-f��"B*3U�1/^��`�A @M��{<^���`/s��mKgƬh`��?�:����z���;��vx;���7�&���4�@jk1��(L�5L=�4��D*�[�K˳o��l���V�'�\N*ZM�[��c��g"�jl�}s4��۲��
�p�2q�KE���ʷ�E�|��)kQ��s�U2�o�X��V�J���Ǐ���\*V���z��t"��c��Y	2�֢t��r�����y.�aj-��YCJ=乊��yߎ���V��Vf[PcTR���a�+v��z�������tA[�z����M�"-�y1�̡��a4;�-��w�z7Xt�L�TǱZb'%��ݶ:3rZ�9eo�m�Z��U��}M�du� ��u|�q���K��w�7j��ۭV;�$ָ��̇�Oy=ӭwN&��(�����׎-�cI���m�WX��v��-0wrvԍ�`iC=������߫�7�-go]z��Ek�Խ�ݯD�\��~��j�%[K�R�G1��6j�I'�@GL�k�kR���!$�(U>��A��K��"�*�{�mq�ty�t{���o���D/^i�Ģ\;nzԳCm�i<چt1#,�A�#�ϖ�����4���#�>�a� /�a�־�k׆#_U���H�5	��xD52�e(mqb��YmEC%*6�����^�b}ɍ��O?�UJ�t|�����
�m��GN���y�k���ב��
�s�"�7~�&8'����� ��A���*�������i�y��#쫍�{A�Z��E^`L�#��Q�n)�U��W�U�B��ǦZ���"B1��.��oκcy�q���:	�iI�G�u�?�AfQ���E��8�TR��e�1#����5Ǿ�a�j^�Ow'wfT{��i���9�3KF�I޳��f��D���/a�u\���eZ���6�=ohep��G�W�v�Ww)��4���g���Ij��WuyEEz*�7m�Y�;���j����b�<um�� ]��)s�v�	]`�Lp\�3�0�L���G��/��d�7�x7�%n���(;u|q��f��&N�u�����4��|�/�u�O����3�C���'wTDz�KF�l�l���%��Oq���j�G�<����(��(p�f. L�u'����c�d���ðy�3�_����E쉊~�c����Uw��\�ɻ����F��Wy^�޸����![6Ó�G���v1e�}�K�'��2�7�i�Y�]4=Sr���O�\���3B�?�Ƽ<�;RV�e^!^,��̚�т1}���Q	����<j�Ӿ��O~�h��]}NYy.���D��w/b�M���ևe�.��\c�<���h�p%��_���Պ4(lp�]������g������������S�y2�1�u�t���A�T���F�C^��Ti[;�Q�j�j�HÌOz�zf�l�gvR=:!���.�^��>@W?Չ%睇�o^|���M��{��=�@͵�����z��-�	 :�<���C��i�O�[TAv��i錢��W�1&�R���3Ej�H�S]qjm����P�zR<N `����q��x���>�㩐���A��Xq϶��rS�ۦ���e٣�����/�Νx��scm��C(�e�ev
�H����ǫ���4Ր�w���0�r͎�KN���}r������yZz����n�|��RÐG�����A�'1�n�N�r2���K���a(m��0�΋��گ��[�=^8���!���C޵��[P�:W�L�M�'��C�kO�P�4d�!���,�J�Ԕ��3(K�k��Ԁ���5�e.-xaY{�t :�1W�|#8?r�=pA�\��|h@$�̼��4�u+E�|�����������Q['#;��t��i>\=���h�=>%N�����^Q��^�++bʕ�6�}�
�=[�[�L(����G��5��:�K=o�����NԳ)N��Z�6&쓔^�:j�N�׊cl���Sμ�\�EtuX�ոw�'�Xި%Y�(�YQ&6�Z��tܗ�]����,W�!߽vw����P?+~�W��_L�~T��x�f�Oi>������jL�b��z��*�7�+]!�����D���ʀ�����e��Vo���]�Ua�eL󽭖.E?�ZD��������rz�i/84�ʟ�zӏ��0NsT��Y��ݧ��/a���A�N���kB��,ؑ �ɥa�[�Yx��(P��k�Qۛ��<����
vߘi�ރ
�"�(N�ڪU�:+yg�����K��4�U�͌v2�� �AZ{E�Fb-����oN�#���Vs��Q<�5ˋ�8,�C���j���ts��U��[�7������o/�Rz,�Z�j�ϝ�.�>/������rUI�x��%�b��Z+iL��gU�2SA�{|�v�,֎��q'�#|A���v�u	��^����Q���Z�+q5ݲ�c��e�ƏE�Oc��Ӝf��OJJYv~�˗Gw�u������yy��d�so�;
њ|c�a!�ؽ�4�܊Ao�V���C&���k��)��\�{�b3�l2i�dE4�i�%���8��������R��S>\��Һ�Ql�0B=��sT@o�W ��� #x��m(�/^2v�LE�����K4hկA�b��^}�����{���銌.�����G���U���Z� ߽�Gv=�^������.��*�����z��/0� O�$��/;��N[x���V��d�K�Tw)l��/2�G$�6�N:p����<URqL�f��S@�����ϯ�����z<�a�
D��\i���URjx�#���۰�)�R���z?��v<��R�����+��f����a1�b�+�W��_�I�����p��+�гso#��#���E�MCC\�n�k#Y�5|�����[VYXH+9��Y�ntwڱ��V�l6��,wh�;f>��p;�G4��4+T�9j����p����(�X���q�jؚ��gI�zq�wt�����Ҳ1���qs�ࢻ>��������s�aa�De7V=j�V5/=���/������N�˥�o�ɾ��{.���W�3��u�s�5�=�P-�=��.�w��h>�a!\w+�m����["��U���U&zx�ul4���{F�c�{2�@��{�x�����ɞN�w_�VH�.�p ��k�GX�6H'�-,�-����E%r��S�U����{��v׷[�M�?k�k-�FN��o���G�6����J��x'w�vu�2��өWD�kϬ���s�)q.��ɖŮ�U=G�+��������/qW�=@x<5�s� �=���rU׵�֌*�!^Td81�F�י��҄���s\'�B�����.�;l�Գm�e<�t2R4�o�;7���WXo8ӘI����Gr�����=Y�ęe@�r��\J	昜7ơ=�2/�X����L�ލ�(�αF�kڞ��<
T�*�Q�`?�|���4�V��ڨ�G.�J����$5S�W<�nn�"�q�Wk2t�b:��M$��y@]K����d��6j�-S�;iR�GX��J���^?z�C�hB�͗�$�H.wrI��3��ǚҞ���4���^
ܮ}Ѫ͜P��)�j�q�]��-7X��ڱ��fT��y7dǼ���Y��I�
\���o��#���6��9 ?@;^�[�����}�jU�j2�gI3�p�t[x�c�"��&�W�U��/��J��-zV��!��<tpВ�n�6��g��˹ځ���^hU�;(�c�t�- o�N;�6��2����D��ܧ�3��)/gvt\j�6�9}�wJ���ֱ����;���M���bi�-��r<�dWX(Rٮ�Z��tk�,����l�hT�<�����2������{��X�OgH��:m-r�>*� K#rx��՘n��^ۭ|0QG�����'��z��i�&$�<��|��Ҿ����y�V��LU^فW�w+�c�h7N�Z��c�FhB|��U�sӗ=�/Ճ.!H�wd��S)�{��5u�C�7),4���h2�<�qiU���^�M�I�
�fA��Ch؜!�:zCY)��j�ך)Z���0�v�`�VQ���X�={�ݍ��~J3��C�^�~ţ��-!�4�B�K���J�V(Ǎ���R����ރ&!k%XL>n��×)�ל#�����)첻r�\#9�|sJ�ܛ$��^�U6>X�QY��5ݦk��Z뜞cE��e0�R9�ق����"
�]6�(�4eq����w�7X��d���n����ghc1�{���}���Pǲrb
��OP>��;����Y��C��TiiSn�<S��m�h���a�d�M��o�+ب
�8U���6�\�r�~�yU7�W���Q�d��6Oxc��돤�)	�}�	��:����S��9�J*E�]W�EiB0G;q����/sy.�;�5���(��E��B���{>.���	'�#���q��>2I���rJNj%$���c�Nu�Д6�x�d�E�lmV��đ�Σ��Q�9}D��J��د>�4����k:p�G�؜�j1n���$5�8���҆�i���R��%��f`�y87*Z8ZJ�/�%\g�<��(?�s�
��f�U��l���;�U棘���;��ٝ^.f�����?2|�҂ 4јi?.y�������>���V#�����N��[9ڀH������9�#��d����z��3^�:묥�xq=¯K�q��"���V��x`��W���eqLm�V
��yK�����z�:9�h�E�N��kY|�\*��9[��W��x'�C�~�~����h6Ժw���YϧM�]��8��i"�w�L���.�N���:b���i��s6뻠�y� j.=�s�K$L'%�a�D�����!4��YE:Ȥ�[�E��^Rjņ:�t.-�/$����ab�ӝ�>�O�`��Hw��vw ~��g��R�y��գ���������j�9I�N����� `��5�j}-��5^��C|�������=	&�yCH^����R��u*�>����,/��l�٫[L^�Ϳ��uN!m�%9��˻qXHđJ��$�^��A�C;��d>
�¸�+ ���!��N�K���x�B�)��X �YǜG���'m�~����R�>�_�I�!¹0.Q>���
U����^��poz���wNW1v!N�A��)���r}�h�K� +�(�a>��K;} ��E'�/����l�{q�^^ۺPW�/���
5�.So�}NП{*�K��&3|��߆};M�p���+ۯVo���ĩ�,uL �_����#L�ȤX��;�w2���t֊�}A�A{7$������[J��g��\<,{��C��/G�X�d�4i�a����ذ�wՉ���ֺ(}]Ԁ�Y\�� ���!�HljQN^���Q��_����o	o���y����C�P�]���in��0o�����5�UE;G7'B�r�T�W�:F�mu[1�m(�zҝB�)���fm'���xk���9�C������>����X��A m�=��5��t��j��k�#HMTU�z� �'v\w3�++e��V��d"�WM�8�F	L�Ht��Hj��x�<Ӽ.��+ܤ�����:��o�;�N�k�$�<Jz�%@���w.����u�R��u|�91��c��͵�o'j�jjb
t��P�r�h]u�4�׮�^W"xn:hW����+�]Q����.�d,�t�f-��.�[Ηr��}lQ�3H�|b�h��h�92�ރM�2����3[�y"�+m�.���KR�lH�����+&��qAvԮ�ձ�[��T�{\�������,_3�0�ػ��|MZ�f�B�ƈ�B�J��5�����-�Z�c0`�N�2�>�=WC��lYv+)��_-m89b�7�gE�Q�ǒ�yq��&�y�2
3^��]�&��ݓ��=��{����)����l_Z2Pe|7%[�^��A0-��GH�����������[6%����j;��&�Z����ǚ�����癕��4�nI�˭��͵VnWf�ltŶNI�����ƹ���]��wب0�df��&�8�P��OwI�9F�i�o �7�6o�fv�[������s���/�ƵPy�C[�&�9��Wm��]6�v����S��n�0�!}��	{�����"nW���%J1�m����U+�[M2�����[��q�h�\ڕis��ˬˡ:��8��a=׺�޶6�����m�n����Z#�9�eG}�����M���-j/�/sma-=5��\�4o=�M��0�n|Q2�as/�ͩ6�����vF������d�VS��C�ޮ	�yV��gWt馝��J�Fm=�2�*Ʀ���[֍<��A+��ʇ�8N�d�j�啵��W������v�Pk�Z4�"�9w�����z�6�O�|�{`w�J�����	�+��)�V�j�Vc�O:^�:U������u)8np���n��E�$��b�� �]7f�E�eu�U��2%ɀ�zY��M�WA)�k�����ZJ2`����K5Z0�X�����0+rp� �9�t�����es"d����m�{�2�f��BS���suwv3/�jٍ&��ڸggGq�N�2��E�Y���j�[��8�6��e���=�ë9�N�&�>b��v��۫Y� %���6��!��1?�NR�k���ŋ���bb��1���>)��v_BC�`�b��J<�8�ئ8P���T�����'m�A�Q3�����5���|�q[}��M<�;����f�}ݻ ���ԑ�Ma�|�Ά�L��i�=�{��Ϗ��T|aXe�rQ%I*&�)gYdFYّ�(�Y!f�Y�j�B�4(�%�!�
��\م��T��s,%T̠�ЃUf�5
�CD��Ft�����*9p��Y["���:�gUE��si�W)eU���N����ʍ�*W��D*3
霳�A�$�#��d&Eu̚�IJ�¢�
��"f�Q�R`EB��aQTv�F���l�����b�uA�Ȱ�@�S�W"�0ʈ�*�-,M3S+3�i�H�TU0�
�ųkR����Y-�4M[*�sYQ
�NsEVD��9MN�,9r�K%9��F���B,1B�h�Q#��Y���R+-8j�T�e�BL��ȹP��ѡ,���P��D#$�jV�J�TI�_>{�|��x��@���v���w�]�<�oE�3�h`rpΣϫ(f�
���EĩV#��6h�l�:>��9*�4�'n���K/xn�������?T�����
b�PT�}�xEO�ro'��+eӿ?P�G�	'o�������	$<����&�,�~G�o>����Y��i������������D�d��j���~�Y�ds6�S����ݽ�؏;��؟nܝ�~��ɏ.�v�z�x=���aw��w����~����r�L���9�u��ǝ���8��$�C�|O��r&��+�aW~M?O^z�~|��ڛ��}�t�^`�������j[��������<����������'~v�����N��������C�xOI�>_	����ô��~G;��nW�!௩��P���㿯߷������ѳ��r�nj~`��f��;6;5;C�c���s��X��
������yM�N?>w�ѿ!�χn}vߓˉğϰ��o(�!;�|��_V	4����=&�^��������p�ǟ����8��L���$�4���_��C�n�m�ܮ�{w��oH^m�{��奔�q���oI�0��_�?x=8��	Ʌ���(��9w������eӹ�O[��HRv�OG������ I'�?}��-MKg�R������x��"��"�����~G�
r���@��8����w�i<���<>ݿ'*��ro�O�o>����bw�k�|���ߟ��0������m<�o��pxT̛�������|<���F���{�G4�y��3�����= {Ig��˼'���z���raW|q�����~Ǆ���>;r�ԝ���{C��o(Rw�k�?����S}BO:����_��-�Cn)������Wk͎�����ٛ�����Wn����<+����ݽ'����׸��}���s��|��x<�r�̟�?��aWryC�zBM���7�99����N'^=>�t���ͬ&�RO�'fmv��=������}����׻�~��{v���>'	�����yw�iǿ���=�yw+��ϼxM��y7���Ńý���<;�yL.��[�'�]����~����ǞU՚w�ޗ��N>���PLW
�~�w�eӾ�{�@�v�?x�]��� O���yM�	S��<!ɇ�zw߰yW;N�{�yO�o/;���}��<���9S���m�7�'�o�}}�蕥�N�a@��H���h{OS@S��
Ťz�m�+s�����ޠ&|����ҮX��}�q��=�%������ŵ�k\K;�aԹ��/}�
��Z�^���y���vJQ�r��<�P�>#�VҺAً�K��qE�����!_P����ǘ�����<&ט��⶟�;��ۜY7�'���a�現'r~q�|�~�ߓ˾���S���i�0����O�����x��|'�nGf�]Z�x�i0���	�/����s@�<����V�����?�7u��o��o�0�z��lw���1��7���o3�2{�(b����k��5 �m��̇�cP��NG���Z)
�@W�*�ro�$<�����7!���'rĜN=�q����RO	ɹ���{<^������Q�ޝ�|q�;��?�����r�0v��C���ٵ���s��q��3k���^�]�>���;oO?�߸=;�zL.�������þ�&��>'�y�xL?-�I�u������;���;o7���0k��ڡ�N�.�g!���j��Uj�vq9�r+��wk�����1�v�d��xk���~��$�;}N�����	�	��O�;R����O��<����O��:v�i���V���<&7����N��hvf��ʻѭ�:�:�ޭ�� zIޓӎO�߼oi�0����?|C��|v���'�n�����N�G���o(w�~?z�y��xO��������?}�ӷ��ߟ��{:۝?����3�m���O�h�T�'��7&����}O}My��|w!��raw�>�~��;��g��7�$ߐ������7�99�����y@�IĞO��yOo�n@��������f��5Х�cs���k�!ɯ��?jǇyv��ǒ�ǁ��xv�8��%��۹�}�ro���o!����F'}M|��q������?'����{���E���>�o)�|��.e�M-���oC�I��ݏn��m�ǯ{yO)�	��V�������o*�nӽo>������yOGXP>��v�{�ǔ������ޓ׈��A|��n��>�yv�N/l��vq�2��kMjHO3k���+i�������>O߻�<�'ｏo�xO9����x@��>���|M�90���ɼ>�{C�z6;�e���=���N��o܁�C\>���m3�~�&U���p�G��^������S����KN]^�2�]��<���o������j�d��NK�ņ��}�q׎�|����%ɇ6��5:��on�wo���1e�l�y���J����֨Q�Ձ����˸�+4o7���]�J�{�t��n �fwosr�f�`��<Hfk��N��'����������]�w���q�0��;���ێO	��=��{�N���rz:?��O)��_����ؤ?~c� ~�DW�G|��7���K#d�������Ѓz���Bz]������$��v�Gϟ|P�K��z=��o(yC�k��=����Nӿ�����i�v��ޜz��y@��۹o݃��xv`�n����jr�&��w]2F)9�W���c����n��f���mv��i�����vQC�_8�C�a�m���7�?Sr�6ߝ;��nO����yM�	S�{?�v<�����S�������r�f�jv������l.�Rz�Z�0�q�	�D��������'iw|
o��N���'ߘ�����O&��ڭ�����
�_߻�o�ra������w���uo	 ~Iޝ��{���]�����u5R�M�麵��q���?B>F��~����>O������N�������O�Pmzh�3���y?� o��kة���#xz��*l��Q5j�����k8���o����O���9��Ώ�
�*>
�	�8��g̛��+/fn�}����ld�tP1�N)]x�u��������qZTV=�)�W��%"߮�Ǹ [����v�wa��N�Yu����y����1����^y��[Jb���'�5�ƿ�Sv�`R�D�/uV<�M��|F_��]ƽ}�"�g���~�|{?-S��!�(u[|��-�ޡw�ϲh�YN���K<����d�'Ԣ�Q�D��qy�P��IKS2��XI�x=���bg�Ə^r�������x<,MӖX+��Ev5�c��XJƖs�t�ѩ]*�Ν����j� ٍ�v�:�Mm��3�6�{��${��C��kQ��r�N�5n��/Gx�T�vF�c�%ʫ�A|��&�7�׎��F'����8���R��*�Pkyׂ���T��#�����ا.��1:(kb�م9��^��Ӻ�4����d{����&��%Auy��C�`̴��T����q��[w�*sKt�K��F�@O_�Ú�9T�d�-@�G���k��\+���];��Y�F���6��&��8y�%	��"_(&��mR���:د�u^���kgm1�6���E������X�?q��͍������g���^��^	�זQR��/����X�jq&�"noҠν�L,{#"cۡ����-�o���ƣ�����iÞO��i:y�d���{����ﭗq}���(�`5L�����ڣَ�UR{7���9����*p�c7\�-Ii0�阊�o��7n�:!P������������W�A�-��O(:%^��=�������q9S��Ϲ�S��~�ê���������\��P� zn� +ew3D��H��Ztɩ�tșHD(H6��4��l��zm�}5 A�DO�l�`2њ��j%PkRP�im(�ŷ1͍fy��h�u�{L����wi}ˆcUh�69�'����:�븯hnR�9��ݥ� e�*����8v��ۜ�Rg�N@Ȱe$W�L��sT2+b�wJJJiھ�m��ѺZ�36�^��R�j�Dq���-G[�O�W�&s}��I<i�(�\����Ƹ�S�J]	��m�Ӗ�R�k�'��b���(��`��D�c >�(�
��e���:�R�|H�'���>F<�yO{*�э=�G2�}̶A'�Bց>q�CW�!�
i�>2]=�3#�����h^�[E�������mS"���푾����"{�*��CI4�� �²����=3�U��K��je�X����We����J�44A�_��M({��{X��A�S2��<�@Z!f�"5�l�VU�Q�Hkd�c���s׾�ea��@�E�#��Ѵa�76:�W��!��OӖ|o�S���2�	�*u¿!8��ӗ�r�S�36����u�*�orc5�β��xf>~�����|�׀j5`8k�|���ew����X?���y���ܝk2������D!^����C�گO�9�zv�l�DR|~���}V5}<���^Y*D_����Or!CG�[��AV�f����<1�v8H��R���#^��r2醞��V�y�Ҩz�'iԬ`�3͞y�9E��^��1^kYᾦid�ת���Ut+T~O������=<��W�MZmD�	U�t:��e�*��
�g]Ĵ�<fu���x<?k���Rh�빧dL�YFrҺ*{񻧎�UW�zt�%���EB�;����4�:�ZM����Ϯ��_Æ����u�W	g�9���������Y�,T[��V��Q.�Ey�G�J��3=�&W�������k���0F&ߦ��w�+r�'�Xߗ��1*�F_�xyo�����f���j�c��b��6X�Zlh�*�Z:��N��$�ڌ��HV>���۪u�2���:�EwmK��^�k��²!�4�k�ɘ7�ሙʵ��5�3��8BIRP9*��^�C��\J��s������Um��}���x�0�qt�����G��r��_���8�UAl�AiJ��jqZ۩��hf�	�%ğ] TC��SJ�:IA<��2���5b|Tkq�ޫq#�[g)�4C+� ��R�]��^\�<T��Yr�!A"� �c�:��7wr���"K�6,�M��B�z�H|"�d0{���[���� *����	�T��ӳA��ܣrvI�g�u�����3�@��׸_�dۊd�C�*�v���0��-P�w��#�+khۄ�u:���=��W7т70[g^���{�}��<Y�,絟������VVU���qo�����e�n�v�Zlcser#8�I�X� �{ݘ6܌��e�du]#�K(��X�� Q���<���%���}�����W\�t`W�x�TN���/4&2N�"�D6�t �!8�>*m	qZ�k2���bf�#�f2�7� �^`��B*���8L4�x��G:3KF��;�x:�U�t�B��'�%���d�F����=ֹ��͑R�B������bk���z��<�n�C�uU�����f�u�D�.�K�S�6&�g�F��D_�U���CA�`�j�s�ڻ2q�L�+(��m!y)���s�%�5�.��>yj�y1Nz���)M�X#uWJվ`���s*�5�3��N��n���'�9%��ح�.��Bx��|�*鐻��d4ϐ��N_@�K="u�wI���:�^��X��Bmu[��|/�U{��T��^	���G�r�v\#Xs�������T���Vj���+P�L�_���'��Jώ�el X��b��..K*:����c��X��'�,�҅e.C���Ǧ�9���Ѽ�Cu
�WX�[���<F��|�{������n��T�*>M/B��]��!��g��ݘXsl�#��IW:��78���R���;·��إe_͠�3/�������
h|/����؃�~�YAU��`�U1����^�mjw�o��r3RZ}"��^��X�y���
�]����>�Ҥ�+��
�����`�_vv���>�Y���y��crkej�F�EK������>8A��6��>J �oV�&�gp�7EC�etysK��9=s����Q�Ya�s��n��%��W����< ��`oj���^�~��nL%�����\6�c�'%��o�pd�e��|�T=ҩ���cõ�����Jrj^�#�a��R�C��̖yp�K���jQn��ɢG���d���_����v-���0aw�;����m�7]Ԁ�t�P�o:�WT��'�q�g�)Qg5��.�l���[�;	�������sO̘��@�(�*Fa���{5��׼��\��+(�ff�����!;���T�����o��p��z=f���1��p��v&����F���e�tӁ_��|�'|����Ma�T2�m<�a�K�ny�/:��	e���w��h�=���V5\�7�zr�s�� +}���g��y8�����]]/c��Cm�^���{~ɪ�` ��N��ey�*z���o��]��̱J<��y��
���X]�~z�Fһ�hΪ��#W'>vV#oS��՝�����M4 ��p�I�57�[(iQsV��0N�0�m1P�N�(WXg\�E<�v�� �Y�21i�O�����X�2ƹ] ,"�_S�*Kd��]=�	 ��e��}�7����XQl\�� i�P��qwʰ���`6:�i�*�_�w�پ|��o=�9]�ڧ�V�׊~���ϱ\�hL{Ʈ�W�P��n�aVt'>�]���2�f<Mj�B/���e�z��J<�cVE��;RE�����s�ws����g�L:�g/y ��/�͞6��~@*������ƻ?b�z��}�Oݫ.?�� 8*!p�g�F��\�y�?גztu�|+(o�p���T3�p=ʧ=��]��Nq��*����˚[#o#d��ݲL�wL�岽1]��'�<�YUoGT�
Cc�{�H�'r)�U}����0�̂w��.	�f��@�jC��m4�x܏i�%���8��������"5z��u�>~�������>�w9|]��N��3���N�2���:/��;w&�0��Ѫ�Ϋ ��a��+�4i���_�WyQ�w�P�_�j��J��c�my�h��k���9��Q�98�d�l�6=�))�z�V�^�p~�@{��!G�б��:�g���x��W��ic�N���ƃ���c�B�[��d2�h���I��M�4����p�7Xo�Wh"�^4!S�&�*��ܟr�s���y~�180�@��/X떢��F�҇�nS셤��*u)ϧ�k�cQ��\;��؛��3��������+�8�Rx5�=�kոc~ݖ O�S��8���9{w�����0���RV�e�;�΢Py�Iy�L�Iy�La"�,؞=��C�w�F��`Oex��E��������aq��IᏭ`�C�����d����S�\sT��@$�3��4W%���+<2O�o�1�^6(�^�dzg�G�����g�^�x��Z�=t�B��V��l�
�o��]��YR�>�Z��Zm׺n`d>�i
�e��ۊ�.���7�0�N�7�����IkvёN#'T[j�v*�{$���n�ݐ	x�0n��Qva�8M�{�.-zIñ��*]أ�f�n�]�/�x{�<�I���ע�N���ą6Ml��9CC:��޿�r��8�8&�̴M�ϳ�]�n����d��R�ZT��֔�r�事3�͜I�tU�s}��,׫R����OE[��V>ن}��%�����+\�n�eS��~�x��u�Y��h��V ��t�p_�ק,���G�uJ�g��������v�F�@�3�7�fs���Ԧ��gP�X/h���+��:�@���&C8�R깖��v2ܗ[bҙYn��L�U|�4��!B�Q`%��8��\
�ف^��n��=I�n{���g���xZa�u�J��,��.V^{�I�l���{7��	q9@�
��e%�
Wn���7�v������U�mq�ϩ��<&��/�fwx���@T��9�4�(S�WP����Gx��x�k��0n�;G���<T2R�d �0��)�k5�Y�BT;E��$�v�h��+�܆J��Wn��gC|�4D��g �g>DGm��I}J��i�`�Ӷu���YXO�ռU���f������i��7�S%�'Sm���sTN���aL��qipp�Z3s��Wn�i�-g:���)Q�+Q(���H�n���C/	'�X�^�pЖjΎ���e�8�LZ��ZKU����Ŝ�=�l�}�cwEu*!� �L���Pfk��"���2tng�A	��̄ܕկ��Ý]Fd�ʶ���p�7���D�ޖV��(�^��v���vq�R� +����խ�{0
�mj������&
hWS�7����S��ݬt�wV��/���5ڢ�s��oMe�"�U�ȗ6>�|�:oGq1��҉�y�[o����ȳidV�:�����a���,��tZ��]Q�[tƞ���1��,O�7�b��Lr�<�Z�v�Ek9"�@hN�&���ƚmK:/q�T�{�U:��Z��rw�1Vo�9�`5���ih�+r`�Ơ[�\�5��'�\���ͺ�P��؜�wQu�Cj��}��Q.����j��ەЄ����V�L��!/O�=����z6��1�3��G97�;�&�D[\VL�(_�9J�o[�vwU��̷��y�S[�q�D&����co��T縮�Xܛ-6�� dͩiMo+�4M��]��p���sL�I��C̰�|�*��Q���)I� gh�;�[�Ս.T���eY9�D�UEIgXn�y>\1�dBRN���;��
���V �wv��k�<l���pkc�Cf����k���Z�DkU8���k)�6'b�����޽�Ԛ��$Վ�e�@�����fql|�p�iWX�jt��d��ŷ�[����$�M��Q�;|h�)�C������:)�{��]g�yTyy.��"��d�5o�u�	r��L���]bu8��g\ű!����ԛ�j���h����a')��hҊ�NFw,l�ʖ�w]*ʂ��q�syKyVH�%M���Z����f�<��
�H��#flܔ�R�A]ʶ.�sI�9hh)6|�n6=���՞�M�Mν�R�ى��)��kF���s2�˕-@���?��s��&�څ
T�ھ:�.5J�CnZ��;�q��*��ޡnu**���&�)�e��I&h��D!�"�L
Q9DQArSN$��I+�it"�L��Ќ��UQ�+1Z�DDqR�!T�j����F��YĈ ����PY!�*9KB$�Z�	DDI�J��9p�"��P�Tr�+�B���(��M9a&aBE�%j�#K��ht�9AȈT��u$�V-Q2ؙӧ����K"#��ar�*ZmD8E��dd��+��Q�Hf�R����G%%C���D\�+JB���Qi�V�±NF��J��i	u6E+ICJ��Q��.�\���j!�(���t����A�IR�"�Q���!,�I\#:Qa���UaZ�%�S$���N�!�)LK@��(�(�j%XI�¹ʢ*�Y�Q�IfA�*"��rT���E\�YfHQ��ER��֥M 5�TW
�]�]_�<�\����2%:��[�Ծ�����Q��uԎ�8P�	�AKV�k��=j�Q�t�v�w��a��M� �ߛ����ٺ�v������F}E��h^���!��TI{�&�+yCuM*��%�[�8��zT�6r�^�ڍ���K^	�/T6��%R�VϹ���>��J��n��Ǹ�������3й'[�t��V�K���ƥ�9����~�Dc�c�}�ו��@ªP��3`t�lUI�,�E��֍k˟C�!��h�q�-x׽�By�)er�O�8̗��N~�Ka��Ct�@��m��7�d��E��mvOJ"�W���r�3���eu#�#u�G:h���ͺA�D�.�cX�+��YCT�֑�sWHX�����Y:�*�C�~��3�ʩ0*���� :��~f�sdT�P��k��{���y��}��Rla�8�Q��K2�KTهL�؉J�������Y���D	dnC�~x�.��.��'�ʫ/�6�L�yt��#Y���jk�.�S��2퍩�}8��b�����][��P2ײ'I�QGl�
Ck{|C�%;;���:�2�6��}��MT��!ņ�oK��*o�GO痎�W���wO� ��T�Ӕ8��,x��IZ�:���i�s�2�h{���㑛��{�l�Z�<�OU�M�x�.G�&<c;�їW��b�#y���c�U�<�F�.��2 ��nz�o����(�,v�4+ks���{�ٷdI�)O/#�k�4��Yk��X�2���N���/z��N?i�����И�NVj�I�v�V��Gz�dc���4��O��W��U�����U��xV{MG�*x� ����B�p׿o����]�^OX*z��K��/��ta�	���}|(�$鋛��	9*m�pա���:3�b�+��b�t��7O�����F�IC�T�i�U�ꝇ��1.�a�♖Iu����ιg�g�( B<��CYJA9��ܤ��i"�{9e�ޘ�}Bڢ���z8�l[Ճ�*�>���^�G!�ws��s�~��OgN��(X�ꡢit������Y$2}�����SY�U4A�Ӛ�l6U�b��ya5��ε��IHx������ڇ��ND��[�2h���/!`�%��^��
����b/�����Ğ,]y��߽H
�~���o:�V\Я��<e˷�m9ƴ��w��y�E��=��W�y_���sO�ڍ��D7�c���M5AuM敡e�`ոѵ��3���4��.@ŅAF뵽�vGcx9*ԣ��4VQ�}2��/wRY�(ޝ�kT��]��E��7�I��h5h��ش��SKWV�-��;�/������Q���̤ttD�'���[;>f$�ǵ��7;4�2m�u�������{��z1Z�Zbd<?X:<��'�
�E`
���������>�P3ѡ�=D5�x�|=���<X�ꎠ�Y-�~�٨a:p�'|
ȉ|t��C(G��_SVF�G��]�0ke�s��-���&a�.�/9����� V/�͇Y�axyq�b6gX�x��Ӷ0��U���.��h����,z�-�e<T5PL��t�	�`.�粝�}ݴ���=��*�?�b�5��>Ϩ��w��WX�U��y�^��3��Ey��.p���W�i���xP{���v�|�u���{��Z�y��	�1)��h��נ�6�pe�
d��6-�l��#�$[��)D��A���
���dyǵ�{S�����/ �JK���ﺣ��D6�SOo��קֻm������Ѿ+)-�0�On痼F;�zF�D6�G�+گr��B��NPk�e9����^F2L�S
�}�-d�K�yӚ�	/�Ipg:�H����0��^���x�cA������Y㷞EHǮ�h���(�{`�
��=t��s�w�ޭʆ
R�f�#h�#���ae��U�^�
�Ҏ�Uh���S_x�3˫m���#Nqr[�
��q�}���d�c���g�n+���+����3p��\�X�m��x�`�E�UU��_M�ꛀ���:@��Z7�=̂0-@_�}ܪ�U<n�G��.��<�*$��ƚ����'�F&G�Y)d����-�hAw@� �x�q����p�=�<�[Mx�}�$Qͳ�Y�/Z1�%;�R�T������h����({�������ew����<���s���ڻw�ֹ�A��	�JqޙM�ip��ߑ�wDP�	�A��|�'�ݴ���t�b��a���o�۲�	�*u¿!8�ñzw�*�8�3ja�p�Z�r�L���S"j'��wҜ�֙�V�/�f�!ԋ�J7������9��>	�Sj�~���}���,2�Cw�O���=�w������l�DR����9y\�:O�������{��&U��r�������{���V�
�l.7�R��Z�[���ٝ�{��y���vȕ.��C'��X�j��tr"���$W`�1��V�E�����[��uN=�ڮ���܏��'�a�����ɼ��� ���CF�|��(�([�y=<^���j��]�N���
��Μ{���nU��æ��9J=N̲�����<�U�W"h�����_�'.�/��� Tx��'!5��qvkݴ�]�n��I�t�TE��Q���8��|3.�Sά�gɣR�]�	��z���3{�c&���,;X��� �;�����M���ּW���R����ע�������RF*o��e��	QFd�+κ��zP�������x������@OW��1v7rͻVʸ}�rN�|�͏Wf��\M�����U��:�^�:�>(eWw�x����<�D7'���^'=�oV10]�
�!��*�t
��Q�m�NY��y�2Vn��ƒ��(���j�^���d�i��03�z�,1y�P@
�F��ނ�0��&	�DZ�m��hu�-���t��m�ڍ{t\"
�Y>W�劔�(��25��a3o���lH5b�+���1�jY��`�"��OY�V�ϔɉb�)j>� �D�$�/bv�i֔��3����3텻D^#~C-�$2Tʍ!yE��z��lQ�ٳִ�F'�T?�`�qE3���;��HZ�='"^��>���%z�=���zE�����+;]�/�ї��{}�H�rW�D��c�����`Mz@��2�F����k5�bU�:��Ǐ�v�3gOј;�Ǘ� 2rꉑ�a�X�E�"�$QLw�+��6�7b�������;����$����ni���3.«I��J��0@�tc{��諭����Nl\I�H����&Ğ�ئ��T�F��Pj��~����f����=f���;[Zj��	��d%$ث�E�jkF��i�)�cK���w/�dY��!��'��zl�bn=q;;�r��2ԥ��'S\�g��l��v�v���ε`�˓ݓr���oV�dǮ0΅s����k}Ւ˩E�W5c�I��UAm�1��c�o����yO�{y�w�	��^�����ꡮ��#D�q���p��c�W�=G��LT\�e�e�x����́%c��=�n�9�����P{ɪ�E�R�59��Y��T�F��<^�p��̗���çL��^e����Щm{%v�}|2�	�H�Y����b���2r��U��^XB#L��Ƕ�*)a[M��7�x���2���}(z p�G5Y�d��,ޣx4=jh�4�'�Am�/�|��^�v���X���c,	��璴x����h��n�>�+��ڋA�j�Hԑ�d<�sXJ�8�Li��Қ���v~�dZ�Z����S���oA�B��u�\���'�����n��9� �	Ά�8z-�kK�U� ��*/������N�\~�O/�{�fm���4�:�=3��=c�3�SJ��2�N���{�V��KӥUv"ɣ��Dդ���>X�j>�,C��j�C������T�V�j׽���4����׭�iL���#.�����Po�|�o�.�z�ڎOox��ךߩ.k̅��IcJ�P@Qca��3�9��C����d:����sԽ8��T�dq	bV��b�mRy����i��n<���_���IE=��������ZS��I�S-���J�U��7��l��wq�m�<^�ώ>lO��d�&|�J,�2εb�Z��R2rb���ñ)��	<����}w0mҞ,��3̩�~�^��u�T���A�>��� �s��Mz0�D����iu*��ڌ�,^��4�+�ּ߹��*�iXqy��g֪Ⓑ��(z��2����	]&5޿�.`1��j��om晢�W-��CׇRݝ�����k�WeWNX͔�^=��͢��ll:�QȌ��#'u��)����vr:�lс��m���Ү�.P�ˎ�Y��̠��0��IEΣ	|��껜�/�+iec��s�U�L�D�y����A����")�Qx��j���x����Z��!⯙�%�'N;��ܾ&��ޗ�ܞ�٨*����#�X6��)���SV��-�͝w��i�I�H�̍�QQ,Z�U�3����3�M�}al�m��Q[p�4뺐ѧj59۴����_,�m�3(��"L�KӍh��۟Eæ�~oifs�x���[��o�A�ƭ���ﶨJe�Z&`n���&J�#.��**\I��s/u]U�z�̯E�)W�,)�i��~�<6�s+�F�*�<!R�]���B��[���S&%����|����em��%1�%?%��۲r��m�ܽ�L�^%he��KYE(�
0���`�)N�bv�GZS9B��19V�w�%k��!i�yʹx�O3f�m�wi$̦8�T�T&a��i�#ϸ`-��.X�}�=w�N���9�V\�Vr����fJjv����Q�մ�U����UX�YK��S�Y#�ލ(=���v$[J�;��컚�a�Đm.6+�hWi��[��X�-'J�����q�B�b�M���]sՒu,�N�T����g����+�(�evȦ�"���(�͟��f��IYr(�èE��Z�=��}�;���.�U�7b‛)^nWX��BL�A<߻�5����s�/~~�^�����+"[U��ߏ	f5�a�IWp��:nwN���K!J���T��`-�"mZ]��Ӈn[Xcf9�[���ĉ��2�`��6��X���[����;ok��o�;�p�R�C$�&su��Ѱf}�,)b����i�L������w��z�({�>}:ó<6�\%1Qs�L�l�Ŗ�SW�EPR��]ڴ\��;���^-�~y�i��U�u�:�mS>���|<�woE�bF�Ŧ�F�Kh+�(�*fT]̰�_��D���]3 �M�����M���;�M�M�7b�:�d���7�����H����P	���Ѕ�;�M�a�W�_\F�+Eѵnmy^��*Rl�g�}�T/=3z�\�"߱�����<��%L
�񥯐�iLpH+�S�]�;6��}� ਆD��)�:.�ɽǠ�j驏�'����{�ޫ���[���׮��5���Bڨ���Dz#[�ݢ�ս�c�c�v�+yc&�_D�td��m�o�����i�l�L�F��7����/b��v��{�9M2I���"������)��,Y�6a�-RN���H�YH��˶�S/>jϧ*��l-�"�C-�$2$;�r���*H����+e�"���ri�C�v�;|�z+��M��>��7��dn-'�{����	�9J���|���t�P8�Z�YYx剴(֬x��9&Q��354��4�&�L�[AMM�D��R��D��,�BJ��}�=މ��ܞþf�[>dvD֖B|�lT�E�bkhF��i�ן%K�;�*s9H�e]��Mf��+)�6��guNU�d&����FKjk��n5;�EQ����*�����:(R�i�/T3\a�Ю[u6*��Ck��� ��'�c
;Xx��1N�s��a�Դ[U�ֵu��Bc�"yy�vw_���JT�lXդ�A%{l����d��y��Oma�:�.��w�|vx̣׭��?Ccs�f���W�#�KN� Ňq*���hLtnm���t�G���km\��\&���l�3�=sU��>q�й���Y���T��[�� ��Xd�âyW��[��=Z��$:8���K{3�[��n`�+���T;/�Xհ��\Q�(��Ϋ#sw;]������dJ��!�����8��wc�]x����b��]�0�aQ�a�ao�u꾐�p^%Gպi5�~Ϯ��1���]w���0ʵ=P�ʉ�N�!֙Ǭ*�!�ަo����gL.o�5\�Q����n��ǯF5J
��;݊p���pȞb�g�����(����_��4?�q���fj3M6�u��v��6��B̸yV�vje�Zt�q<k5Br5���O��ژӬ���[�%��zՑ�s�t׭˭��ˍ�C��nˬ!n�{�6S۬�i�V�CU6V��U_^���V�A����0%�.g>yx͌���ڏm�Ƙi?�*t�˰�3)�F4�h�N��1l��+�g^�u�VP�E>
�;���Д5.([����C����%>4�>�U�c	pQ�@i�����Q�;;����c�K���OhgsC��)f�W�n�8ͣO#�8;�� S���,J��̢�mr�7�չ\�V2��d�����a��d�����L���r;��ŴewX�`����Q�vl��\��7)�%�����mn"o�=��f4��\Ŷ �#ꓸ���N�͕(=!`=j��J�v%x��8��PM7ۊC[ہ#�.��~��l*�t�iq��or�k:d?���t9��,�r���]�s�7{�y�'��\5}�ҫ�s
w��Y�\���Ւ8%�������9�ĳ�C��) �*�;��hQ�sSZj�`��G��Qݗ�������h�qR�����qT���#�^�M��u��5���z���A��xm+zY�q&�\�Ⱥ`�"���/%�˧��l'N�ym0�6�_�n�%+�sqkZ�.�x��ú�����ii�*�� ���Aϥ�ib�w��'���t���Ql ��=pSp�Y�h�owf'���wM�JY0S�r+�!�n^"�����Mh������,���y:���d�ql:�M�IV���zgQ;��ް���;UE����`����FC6o%�:���2�͕+���/V,��ht!.��Xb���LG��r�7�c����N�֫�-=rK�{�v�7F��Қ�*���;A���Xm�R�Q{g��kFG��!<�����JPl��Z�u�,ʺ?1ná�%+u�^��P��@G��]p��d�oN����&��*�TS/R,*q!9�����Cʇ0'�V�����ӧ��sz����p�[gp�����2I�N�;�Q�]Ax���9@�[7�|�9�,r�u&�ՙ��/w���z[�j��E=�:�ޞ������{p����-FjTX�PE!���4@������Pp�9�"".Q�Ē�9r�!9GC�(�9�i�.raT�]*8Z��@�E�%)9R�+��eH�TD�F`QQDY��,ʹe�6bFT���.TDDDʦU(�TG8Ur�I�(���I�DVT�UkRA!
�&H���V�2*�BH+��\΄&H�)D�R�EA"$�����-�\(�R)E��­j�$%)��\��U�Ȋ��.�r.UE*ih�G(N��*(�h��U��Ra�g%�ER��RU�hu1 ��)$�Y52:�Q�dL��0���!�Юr*�r��,�.E���4�U�K�U���J9fʌ�"-
"�VV�B � �Yp�LΑL�,��I+��QTUr�1� FG#�U�"����D�AIOĀJ(�,sq^'�Fk�ޔP����;���x� ;6������[B���ɳ���R�@�p�`^Y�{<ܮ�V��ّo}_W�_5�����b��#AJ�K+Y����<�[ϬOefQ���s���ܧ�7(,X����b�/W9<7���s���s�]�y�z�!�;�*�F��p8l��^�<����7�ꋇ{y����zY�:�`�$]��ni�P���,��t�xՇ�^hMH�,p����u��VPV��u�sE�daӦ��3�e��z��t��[s�>�u]��U�2&������شb*�s�4/M���=��*�YV���{G����4���o���p������q啡��2�L@3�|��hg6(�s�(ܡ��/mR����[�K��kv���O),ie����l9�v��8�	H�2�͵k9*�a���y�p�bV�� �zk*��04��u�2���ڡ0��p�"o%9F'ц�m\5�3��%�Jq,�lTD\�&��j/]#�P��O'X㆗�v���u���ڑg�,���N�V�e��t��C�d�g��dO��s|�V��YG�S֚�����]^;:�=�v�V.��NӦ�$/���Op��p����gX2�ԩ�m����
�l�u���o{��(�4�N�5��[ �e�V�,�3\I��9MzY
I�˫KnW(�|�f�=NNwө�{����U{��Ϗ;yNy�ʤ>�Viy笯Wa'�l`���sF�y��ώ�w�J�р��e̴�7�V�S�({��/���!��I��cm�ȜTءf�*ٵW�v���6�aE�i�՟z�}|��YgwP��������%K7VV�9��W���J̻�Dm��3:+����<��0�2�e>�_P������s��=�>�ݦC��O�F�o{0ݟPΫ�_@;>��f����� �QXZF⼜�O�*�P�g?r:�d��v��ڥ����9&������Gá�4���^]���&������o��f���L�ھ�s�(и�s�d��;�#��b�u���$�-���ʛ��	�Z���V1R�e'�H����5q��j}�x����h&*3?gk����Qc�0*��x�e'�Xӊ�݃�x�l�[������)�)}RD��ܙso��lS8��%��\�`��:�]�����^��(G� ���B{	�b�v'����w�wR��;n昱s�2���2��������k�������Ɨ�;���T���2��^�ޥ���hd��1%@SG��g(�pہ�SsAEV�Mk&sD19�V�=��i��J��yd�4�E(�@p�VE��-X���:�1�x�g�
ˊ�j�1��K��zN���.f��hU���=,�&i�����{~���Ge�M:��b��[3<f����C���Z��G���ʑY����x�4M�Jx�4�w�.)f�t��Y���߼��k��-q`K=�Qx�����ӭ��S�����>��ve�[��H#ǲvr����d�^�BZ�����WT�p�B��ݙ�S��v�q'�YZ��J����>ŏ�L�f�����gڧ���V���y;j��6����5I��Z^����MÈ?\.�|��c�"r�x��=M5:�YFx�x)�ʴ������v���F�N�(���鏪�'��hw�����Z
Te��g�����M�Z��|})��)n_�3۲F��px�n3�k�y�F�o֮v�}�a`�\���EW&G<|;3�gm�E���F��4:��^VՆ�p��A}��=�X�N�WWb���QO��vf�M����{�Vp��UW���<� $��Xǻ�{L�����ܚcr�j`-�h,vnϬ�we,���x78(�D�W"��jKn-�od���Qw3�;�L�@ݖh��a�Zě�wwWJ$�x�֦�J+�d�VSzi����H������}��^y���hd�Gc~��Qb̝���/�5��W���?[C��};U���V5���ͦt��d򽛖ހVD#�N�y���l�ޫB�L�j,sq�6RgTK��x�X�MA��6�gV�υ	��=���<ف?r����9,��F�v-�M}PV�m��/�gbT@�beѫ�/�τ��5~�E_d���$�=�
:�$��M�'`�ұe�!mU(�1
'�!��-UC����}�r�������ÚA�9gLK���H��؋�YMM�}G���N�1�ړ�7��z�[��}�5p�v�go7dO�K!,�lU�".|ؚ�=���[%��%��@���˘�|��sG%Z�팞~�gS���U�9��� �:�K�-��yA%HҬ�um��P�u8�5�:�e&�e�����HN`�f��Tc\P��'�e���v�ۃ��ˋc;|��Čr�y堲���m���8'� �����_}�U�:ƾ3��Y��י|��5'���d&����f����Rɉ�8K%�`����:��Svե7!�ɞ�\*OS��{<!��٥ƨ��^�'��N��'�Ҿ����(�������>^��1�z��Pz蹜2m��n��~�&w�O9�O��ⱚ�y�g�g*���ŵ�^����P�a@�tz?q�z�>��IN�U��m��V�ҋ��BƊ�.��	-|Ej�û�D�jQ�Z���TQ�hT���(�n�.��Va�r��n5ׄm�s��Q���ݟZ�� �^��_w��/X�}�f�JOV�w�=n�������#���J�XcY�2�]c�M��u�dRKL�O�2Z��O��z׆tL�ҫ�3�L���8��B(��L=�1�m6t���))�i�XSG�d6�sm|�%�NM�����#�ͺ;/�J��n��Ч���˖�b�� I�Kn�H�7�
fB�t�:k*7�6�@2R3�Z ��5�u����/}=������!ZT�Kʢ;n��Y�B=?���ꗪ����grsho1��Y��$�޼]�  ��R�X��O^)��+��y���c�r������o@Vtb(��Ȭ�fB�奸����e2���#�}��l>P��$��d(�c*֫��zL��.��d-<���~W���f!��
՞1V��F�ƍ����5a�v�V���f��	Z蠛m*�ρ�U��h%�K<Ug3����vۡ=W��Q�g)�??.϶LU�8��b.*]�������D�X�5�Q7R�5C|o�3Ҏ��y��M�짾�_)�����bMr�/KQi�U��%�+q��R5��Sw-��ת.$�V�jͭ+vbp*��4�LJlV��j�x�kр��\ʴ�p��+<x���	�Z���2'um{=�lxک<��<�������}�m���r�N/~���kV��bz�Ĵ�e/B�S��q�b��4ڦJ�m���kG#kƭ�2
���Cѐ5�ZF'm�qE����m6笶��3�Q�b{U�ނ��u#��]u�		W`�m�ا}�e�txe�TN��LB3�	N�̆�l�qDbs5.�l�e-�b�'���7�����:x��=�B|�M@�n�I_U�\w��l��]2�л���Y��Y�E
̐M��yR ]e!�ucZ$�����5���f�{�+2�ٔ���Oe'u>��0����f���[m�D��G�����3`L����K�u�ߨ4�Ş�K��|��I��X'?�Q��;�Ph�5�*��a3v,��9)�i&���%]�w'��޼��27܍��<"����V�#��׽�W�劔��,)��/�L��I�"	�������y{�6h&g�5��9����%���hb�1e@T|���*�rE��R��K&\��IiL��0K��nq��zĊo),d%FN����7	�0v�*aj�513n��;h��N\S�V��q	���k�z�N�e�{Q6��^����V̗�+�P���5}�#���i�����~)������)#�7�;�?V�}�������e�*��;[G����|T�wp{�����Ӊ�`�ĖBY$ϓ�.Y�5�3-�!u���m�7c՚�ӱ)D��}yH��y\l��g c�C'v��P��m:��<ˡ�Ϸr��
��iu���L��C��t�* �+.�J
��1�Y.Z;���Q���� ӽ-q�M�c�z暎���)��lI�c7F�+x0v����:cՓ�����������9���7�gvU�d&����d��kр��	w������
��#̰TH�sr�L�+{�J���6���V(B'��L��n��WT�kr^,?N'm�}�m�^U�1���P�z������{��`%'0������<1�Wjg�w��P�ybvU^�L��ϨT���-	�͛'x�D���s�fw��M|����5M9;�r�6���,vn�6�"Bɪ��	�aT���d�2[�B$�-
��7�������f��oiXy�>stQ������q=#z}{1�A�X�����oM3�)u#Zr��w���*�N��l�x542�1i�2d��E��e��Y^��b�*|�C��� 5���hh�3�@�{��}JZ���F|d��^�{��y�:��~�e2R�ݳ��[�	��l���;m9�aA�޵]��ظ=�Q�W��Q�=��w޼�-j�4��*�����(��q �)x?s��'n�3���O`aP����kn�?�(Z�o�2Z���)��yF�N}i�|��ޅ���to��|0t���Vd7�r��������IM�7�٭+�����r�N�v]���W�{̧	m�l*����,�TI�Y������o�s�W�*�oz��1�MOx��������hb�D����j����|s�=̯Gl_�^�����ƃ7���fis�ԝb�-�ij�j�6m<dc��VVD˗:���I�
��V�f��쉭,��I�Qs��U��?!�Bwץuq�X�1���V�3�Rїr��V��T�^�BZ�����s[��FP{h���.��ܬ)B�ϙ���)\�{�Yq�Xl+��ؔ[K[�j�V����S|k'��*�;���Jo�QE���>���Zj哼p�;K�s��%W8�{����ⱟy�~��S����Б��M���2"��)����715xj)�*��[v���rib[b{ܓ��]ҳ���I�N�d��g�X{l� ��¥��G#L�rұ�.�\/�<����k@� ��1�;8=���\V�-l��j���n�t�����k�$�0rN��D���u�S:��%��vB��8�MC�i{g6�ή�D�g]�k��u��PY����t�,�B�i��;W�b4"�l9�ˀv�5����o7�ޓ8Y���FNs��h�	���婆� ��e�hEc��q���X�f��nQ�s���|�{�>������#L��R�G-����8q4r#�-��Ul~��ߪ�S��=�j>�,5�3ּ:&Z�^��>2v��<������6�����K/�^^k۽Ư�{O};EA|�-���~����6�7tp��D��ez�n��/�n:�-D(,b�G��XК[�D����l8��j�t��d5b�s�wu�Zꐴ�+d3Ǿ�|n�"�J��'G��E��J��/*U׎cٸ��+]S �y��]��[���芮s�Ꞓs[k�GM�Ugjk.���S�~~]��w�g���yA=Nq�u�[����@�ӆ6���R�]my�T�F]Ϛ��7��7�q�՝��;9S���:���MV��R����V�e
F�1Lmܴ{�Լ�X�AP�玹%�Q��e4�_bZx�ov��iRO�^�Euv�"�ٱwٵ���t�gL��Ww������0��W���i11�M!�oos�iWMq��r�wj��G+�$*�V�i5���@r�}δ��t� �m�n�)u�0�T���<��i���C5�N}tX
�c@1�eY��Z�cL�Mv�GӐ�}]q����$���xG5;e���K�IQ����������ʥz:��\*� 4'Q���6�^c��������A�2�o�\�!���!���E��l(`c��:
��o�M�Վͧصs�N!XWY�,9j��j],��WS0ʹڡ�&��gPX��m犬4��I��+K�7�>���i����{��;-&Vc�T	��c�� �3�������m%Dc��z�tEf��Wj�ή���Z˽샏C��w�N�f�q�?��T�N����T7��(F�uU2���ݢ����l۽����m�jv�ܽ�ϵ�;.-�;w�ՃX}t;�}�w���#�*8��'y{B�"5 �!&�b�\W��(nf�
nۛ�+)Y1�`}���^��n���M}V
��G�������Nm��9�iUH7��)>�;��ݍoZբ����껜\����b���ʠj��_��/���睯�8I�����X����jWq�\r�"�oD�3��7c|v1r�䔓�o������i6([5��/+5ڒ���6I3mX���1�U}�v���6�NӰ�p�ª�2��5R�U�fD��&�JGgI�����l9���x������ro�������WWSxմe]k�f`d�]�*��t�W��SN�	�lZx�mQm�#֮R����un-;|:��%e0�ǆ
�{8��v�L�ze9�wؤ�X�:Ԯ�j��a�޾B�f��H��2l@�<���bꃃ-b������S�4���6�K�\�9��ù��O��l��e��W�d��x��!�i�"�V��]��Bco/21���ҙ�Bw����*��͝X��;��[���w�38��gtیJ:�
W�=�S�H��}��\�BrY��$�W:��L$n��јj2���*[r��3�)��i���F�v(b�t0�CH=Ak�Zu�\ \�Mdۀl�9��w��JD��cwPk��1�Q�<\�Y6�i�Gp�T��ƻ7[������C�J��je+���(�y}[��	�d�e�(��Z3+h�Z�����_��V%�1�} Ǘ&�����j]�	.�S�(���#��A/����n�L]bN�Pn�S�,u�QN��+��3�hWV�D��j�G[D������c���SD>�x�
��5��E�� +�?Y[˶AW@��I�o#��)��v���`hֳ�y�캒�pg���s�'豞L�����W|���a���j;�۩��h[�O�������""���gPB+Ι	B�TEP��ER�:+9�Pj���*:b�ʒ-�V��
S1Yr���(��aQEI V�E���IQ\�ʤ�L�Dh%t샓#��fQ�VdjiT�ȎFr��"��UgL2�J�Tp궙Ds���I;K��"�D5DD��Rd�AAU�r�ҒQ"���+�P��Vr"��M�W+Ca�	�L� �Ei,�im1�jU��kK2�S�0�eZPÅ(-".UT&QgZq"���
�IȲ.&Av讻#�<�;���D�;��XhETU&��m�Fd�e�.�F��DL�A\�QDI�ETs�Z4ѡ�(�C��R���D\��M�g.��������v�5oޮ��C�0svp�FR�f��y�(���������x�-\�K�_shb!T䣤k+�ѫ��Joy��6�Y��iӓ��0r��lUj��>�D���Hײ�U���?�հU\F:�����;���ĵ�/��߷V*lP�oثe�U�S%��J�劚:�Ya��y�r�^����q��y���D���8�z-��y�mO
�'��7sd���B�}c��,����2���}Rt�g{����NeVM�0��r���2W�BR]ΰ��g��4�6�ꋇ3n%v�6X�\}'�ܐG�0W�̳r*.�Xk=i���]�9ȷ!��ɜ��WtQ�F��/-����K$V9�����5w/�OZ�蘳��9-e�W��_b.#
e)]#��׽W�����ϖi��o���{�4�F-r/+�;��xt��N������8Z�K-Ҵ2Tɉf*@�;Ns0Aow-j����y��N	rr}V�7�1�[!��+hD�#O�I�kCHP�7蟺�8'��zw��Kg�r�0��a��]M�ge���A�H�m/;�.������Fi!�V�9rn�yj��l�������ޝ��{��9° uO9�l���&8�*�o�s�������B\��d���ǘ�]����ћz�Mn�[/��2I�&��y�a�.+�U[��@�+]/�KX��"&7V����;�'��_�����:�J\�eQ�g)�/��}�ү�S2n:����i����#�ĲI�Sm�R�<�r���U{�v�����{	S7]���a�Cl�n�2�'%��ZY�=���V}�@���5m�X;ۊ�uŨl��{XQ��Q�ef�5ĩ��,��L�(A?{��G� V�b�K0���\�ӂX�M�Z�͕dlz�X�!�j�,喢�ڞ��a'k4�|0QX��/h�:ÈO\.��������E�+"��4���O3��ӷ-j�2���:J�t(���zcꏫE���{%����E�/���^[%�Ҹ�UnMx����Դ��X�jgE�啝p�ؔ��T�Ҥ���BIEhR�Xҍ��eE���s��
L�1��-��rTx)-����x��t�B�����'�ǧ!]a& ��טq���ֵ��<�OTT��ș����yL�S�Va���G`]휰f�;���՞b8���`)���S|M����no;��n�R��i�������jcC3�����18tt�k3�AQ���$U�zi��H���Y��<3����=��W��ƫN5[���%]"��3,u��E�	U��i�䲉��w㉆�um��2e�W��z��~�e箈��{19���M�9��2�}�Ch�hg����{jg�
�����5x[�.O0�OSo)!��eD��,��4����8��֕�* %�e��J��;�K�v�i���s�[CJ%�B�a��k���~���(Ո�y�l�H7����>�n���f�ԝA6"���SSCj�6hȧ{17C1d,2��$�J�n�n%�]�W��%�K!,�lE�_�5���r�0B����I;3�z�78�o{>:�����l_T��T��x�2C�
	u��Y�V��t���R��������o��<���S�,�\W�8S�m��˱��v�wnU�Y�J��R9��n��r����5$�6P70n*j\,��{�r�Z1NT��)�g{�Lݡw�}��e:���<���H��eț��������Wu �Y�Q$e�0uhu����W}���q��^a
���a I���ܗG�ӣr���ﾪSݚ&���Wp�{�ym{�%�R��N�r?T���^Q�������� �Q�,}�ܔtٹ6�"�M-Jn)�SQh�ݑy�s�E{����~�L]��Oѩ����0�jJu
�-��r6�Ӿ���oK�ܹ� ;V�s�^<f�l�۶u
h(�m
��zQ�څ�k��v�{��@/~/���="�f��� �^XV�VB1E�Q����奦U�|���K���i��������z���v�՜ԣ��d l\��O����QՔ��Lϖ�Q����Z쉿@ҪgJ	�2�,lPw�ii��9K�p��-{��.T�4��£�:E�W�����	��I����&�
�rmyAݦ���}V�J�Q>1 �#�g�۲�!�-OY������Mh@�0۸�n��V�x���N���QJ$�(�5�O��ؠ�Q5�1-{DSO�Ow3q��^|�3+��#m�]�՜E�ؐc��]g:�c4�$�;.��{��dNn�/�]m֬K�s8V,�_e�A�@W36+�}���R�&v5uݼCof�|e$�mO��V�9�g/o�y��m��s� c���>��e̕V�[7�%k��	�W��}�8o}��=8x���z!�=Z����t���:ˉh*�}f��lݑ5�8$��x�	�w �\��rT��+{�)W��9MԴe����n.$�X�L��>�x����Z��d&�g�J.q5��(R-���3����Lf�W{�z�1��}�潪�h�K�˳�?.ǿv��@'����/���w1�c�u����'��KK��D�VjO??&���x�'�v�>ջ�"��Y�h�ק�;�*.c���
8�������|���OSZ6�_7�μ��nOP�O]���1�9�X�]^�������u
h(�� db-�끺�s����c��R��e��G��N���ux�z�p�%l�r���H!�O{Ѵ"���ypO�r���2�7f!i�lw�����h�BY*P��E.��%jա�v����S�o9Qt��Ly�9[>A�|x����Wz�։��N�[y�{T�ݐ-V�"���)��P.o�'�:X��S��D7X��C��%���U*�H����t//,&ne��S{��0÷xH�,�}ja^��Lq�JEei6P2qܖ����e�ne����}z|��x��Ω���WL��:��`�T�L�aMi�<|ʽth8�0�/O#^��V[�m_y�go�p~���s����2��1߷BXI�?}'�ʺu�[���W�zWg�qn�x�{�q�������kn�qw��,��2��m���QL�E[��� ����*T蒆\ͬӰi�X�漩���g�!���:j�|F�Jy<I�DB2�il^m�1/I��R}�I�u�}�Tg��	^�{�snA��n�Fw���Vf���^����t��&�mQs���^�%W�ǥ%���<T��4��kI��ەk)�n=q9�^z�2JP�e�Ⱦ�2t�`�W�ޜO ����n�r����ق5���'��x�]�W�]�ŤSg:��뼫�>�͆]m^mG���̫i��M���Tuu�"�8�V9gT��'Z�֭��%
�����z��62�̤��"���-j G�F�\�K�|��]�Y�5y��خ6��;5Y�k�ۏI���������:y��t���}̬&��.[}��z�.�Y��4���!���x��t�Q��3��8j�5�/�ܭ+��|$Q�[-e�Nν�<Bsc$����d�2durJ>
U奰ԍ�S�ݦQv�^�5;�"�eq^�{\��$�g��f�m��J(ߚ-�oJ7g]�D�>VmiRKP�È����Q�>�hĥ�nͩ� ��,Y)�kN�X-R�bY+���yW�LC�r��4:V����8Uc"��,u������O�X�Y�ّX����B�}�0��Ln��S(�;��ڏ_9�O�����5u9�n?��S&X�
h�L��7�Ol��-J���L�ƛb�#�r',�nt�C%L� l�#.�؆qE6]�ܵMp��v�.�M�ו�iu���Y+b�Fr^N��:_�%l��m��Y�h�`����	i�5|��r%���u}΄ŋj�5HdY��L���6���B�C��#k&�C:�@e���Zi�ڭ9�d�ټ���:h����f(.� �U땊�����A�xPWѬ�����ܬڡ���D]#�~���_u[���D��	ڎk�x�זD��:kF�wyQ�^3�s)��&?nw����jg̹a��h�Z�-��+R�b.(���]׉hO J>��˩^����}[����U�ߛ��Jux~ZMYD&ڸƐ�ҴP�}W�r�5̶+q��[}�|��Nx���CCG�}�u�c���
���cb%6+A�}�˥E��]��Ve����E^���B�؅y���%�ᐛuR�Jm⭖kUg�V��F��nE���z�(�ܐ'd�;Yb�Mi�QǏXY��JU�[kܲJ⯻I�칾!��U��b�vl~gg�pe�1ٵ��e��N�PQF�d�{��1e}L��+{D���*�;��	�e4kfͅ��l����[�r�2�燗�����+�O]ǫ��Be�(Y��&Pp�r?o��x4X�)3���Gƭ*��47}W-�i����v���CIsP�q�@��լ�ʿ+/	���zr���GۏV�uEɽ9m���cN�b�<����Ɵ(��N&q��'p�s�E���.�+k:����K4�z�����/F��^�#7b�67)j��V�3�,�[L�`��_����g�ݟ9�)F���ع�=�Iz��9I��uk�o���XSGӷ�U�;�����>0���Ԟɤy���oF�k�W����+C%�Ȇ� �>F�`��:(���ȋ�(�JxPϙ�)�E[��[�F%HZyd�4��Q8��aٝr��tל}2�xk������H�J��s����������t��)�6�7�xi=w�fxL�V��ٹ�Y��$a�rDf���5B72�n�9F�/U��*�f�Ԩ�/�2��,�=��F�33�kBݝӦ����4K!��k{^�-~����߫��S~��O�0���ku�!<I���F��fԙ槫���xey(�*��ns�TJ��M|�����)���Ԧ��+z��)a��m�V*�?g���{�+p]��WΖ�)��K��!�s)�:�VehOxs�����������f�^�:,���AaM.�om�t� �kv��Ƨ_��������󘖣�W��V��X��3;q�{J����b���$��r�Y��5�i���Q>��T��~Z�?�}�K�;wI�;j~�ѫ|F����(Q��~}DN^>���L�8)��DeD��t��^9`�No]��-����ԣRz{�>����>{���O!uz6�)��-h�mb^6�a�����WLSj8Z5Ú��9��ɨd��IXZ��|V�eE����3v�=�W^;�M���p��D�/�{9_�fH��l�3��#��F�6��#_'ۚt2��7�x3��2�J�Q���ϕ財-|�+���
�
4wLǦW�&{�iWrZ�0wi��[���C5��ʻ`�*V��������p&��}t�\5����sߊ��	��݀#6�l� ��V�͹jG��^9\H2��4�o6�S9P�nQ�G���U�tvs0�����sL�ZsL��1T�ϖ�KUP��kl�U{@5z���N.���[W����o5f��2��x�]��gqʽ�z�D������}u��8^qQW8�����NvE�pv�%�������nRwS`8�.;VR ,.�<����3�S�5jV�4�cBV"��f3����Z�W1��F9@��+�,� �|"�\���-�%ʷm�-1e�} �5ٚ�Z��7=�fO�]�P�<i	\z*�Z��P�wI�oYh1H�N��o��w�T��w�#q��L�\d��.hgvs6�0B��iص;�V��M1���I�@L�#�$S�\\r]#X`��˙(aOCgZ�E�X�/l/��ⷖ�yv�Ç��S������`=1���&(����p�؄�xɮ�(�S/��y&S
��@+��Y�.�s�l���UsV���	z>�чO]�;������Ю��1���LX��}ƆӢJ���WpJ���gV�lq2�R<��w�r�:d~�ŏU��L�C�c�Y{ܙ](Se�s�E6��e�å��*���nYX;n��`Ql)b��dy
R��L�F��LH1}�7l��Zo�t%3qm+�T��Y��(��aoJ�ރ��k@#�
��,���f_pj�J����sH�X^��g��Ӫ�Qr��;�	.U�:e,�N��Z謼|j��-ۗ�w��N�H>ރ��.*��;v���x,R ��=�k��$*!s��"��ѹ�9�`n	�+�o����@��bs��N<�s�� �>��8��x)�V�/�>��������T�$t �_j�ȸ
�ŷ�$���ZB�Dx^|g_[y�c�]ޔ(�C7Ǯ��]����.�xfݕ"�\���f�ee
��>h��;�[Y]`a|9�].�����h$'p����R�cљ�.5hs����s>��J�����E�I�Ħ_4r���&��+rU�AX5.�����9��	G�=1�ǽek�]`w�٭��V�D��iA퍩ۚ��Č����������SE���&EZ����{N���w�`��`,|�7'��Eu�)O6#�^s�l�wrD����rSY|i��\gp�峗��Y�6�nJL:O�� g'�P�Ǳ�eٗ[�G�
�/�W4���;9��
��d� ܫ#7�����MR�I�2���Wۜ����bg)(�@�h&͈��h�|x�.�:.�dm�-�p�{k"�a惘�ݧY��[19w�����bs&��9g2ML!�{i������=��i`�P��Ewo@�5IJ8&��$���q_:A�MM�{�7���7Y�wK$�ԳF��Uŭ�吸j,���{e��N�,�L�3(��7(��(��T���i�<���K)Z+'7Ӕ��;�d�D�s�t�}o7��V֭^�#P}�,��������W�I���S�hqM��X��]��P���]Gj��@��8r�0�����Ny�hA	+A't���I�˄hH��H�7E�R%9:�Ul88�^��!Ҝ�!�I�ee�V�PT�3*�"'ZEU\�e��\��N�z'�y��"]�=B��ZI�Vd�-T��$���HC�%�<��r"��A�d�drT5�#����+��**+������28Q�s@��\��\�:�Wt�*T��e	�a:������Ľ[)�(�wJ(�=���9���=TN��s�T��r���B*�{��	Μ���q��J9�fNw#�r��ܒ�(\��G9\#�-�K��(�"����Q�t\'E\�*��wZ˲��99��,Õ��E����i�Q�sD
9az$˨�E��'n�NjD�,�Ң���%�G"��'A*
�Ԭ�%�Qr"�V�^�z�����璷[Z0w|O76� G��r�V��-6LMe�!	wìmYiZ:�+w%��TSru���|�\�7�k;�y�faj}�rD��O%&�D[���T����>L�(����m����]Zĉ�
���[&|׊D�idMxڢ�VR�Y,����9�2��3�����]�����7��S5�d'ԥ��!�M�b�p�6u�Y��%i��5��z+�r����ve|�I��݋�N��	�/�)��D��{^�XO���e̫K���ܞ�=B�˓j�/QOZ~���9�BU��P׽��[��X���m��˛Y�[Y���C��w��n��q���X[r����^Z[ԍ����er�_a���:�%�ݤ���^�b���l���S��7�T���(�I�wӓ^�(�}�n��[wo?}a=���+��Sd�O�+h�o|!� �[��JQ���sW�f��m���)��zc�p��2.�,uf�;��Q�ڡ����4|�_v�[l��1�]����WU���o�z:(�1J�׬�s�_y��V�tWj O.�v��N%�|̪��A&�\�.쮮y[�ץ�G)��i�zf��}��*�WJ#�l=H7w��;�ǳ���#�'���9��:KƝs��S�[C�T{��>߽$��;����z<��N�r�+'���XO/>{�ehZ�%PE��L�mcm/��ϛlScʶ�
����Q�I/+�v��I]:HZS*%�b�Ym3����l��r�<Ǔ;�^�Nɚ��V�������O)[AT����9�V�*�����/-9��N��r[NB�f�M�x�ז���N�ب�h�T��㈇ʬ��R6���O�'��s�Y�s]��Z�~~]�@�Ԅ�I�D 8j�t�V��Fb����B2�kϒ�2�Y�ڳ7Q'1E��跔����LO��p�-��/>�Rݧ�bo��������kT�a2޼�z��N� ��N%��L�lT֡�ТW{��v���&L�f��
ܾ��II' m��ҁ��Bg+5'���y�O�/i�U�;o���$��=�O|�{uk5�=�aJ$y>H���c�r�ŗX��q�I������-.�z
�d! fʣlu����D�Ԙ���2Z��lu��(��*����x��El�{����b0\Z���OZR
�zd@�P���*��D�.��"�;s{��(�׸G�:���uC;<~�x��=���&��*ֲ*Ts��=�Ӊ������Y�G���P��U!�)���«�Q��մ����	�0�&��ʋ�x�q�`-���f�����#��ĵꞹ�P��׬�<@�՜��<��8�x��h�>�;k�zs�8�v�d�>n�F��I�h�L�[�����Y"�������:�dkz׆tI����tH^o��ܓ�"�Y��^��U^��Ke�{*�YP��XT}�|5����ݙ ڪ�ZQ5�����Q�>0wK���2[�,��S&$��|�(�+QPZQ�8�<OܽUu�V�Ӵ:��+�{�&"�+C-��,m��n�S���*�5M���
L�>~��BsXo�U��mwz_����a�<&{q�k-��ir穋hJ��*-�l9�g�c�.�Y���ܪnP�=��pU�����-�B��Z5���c�q��"<�Ժ�nR���	�t��&)�!+�[|�6	�5Ko��w���t��z5���obQtr�5p�dD�����զ�\d"�o_s��	��g7�;�BΆ����%n�q��3fB۝[#�ĲI�Qщ���R��u�ϓC��G��^�n�`s�5�'�S9��D֖B|�g�����͊�C#Kk�ߤ��Y��l�z����gw��5ĭЯ/S!4��J2[U]W���Eym{S���z!n{������>�Y�֢��0�xl}�h�(Ci�Vb�9��b�Y����Z%���)�=C=ڟ^�������R�9�ma��a�i��f����)�4�ӷ-j�2��q񟽉mX����C��˨V����pi�V^��XLT]���5t���7��x;��ڠw�#��ut��|�oB�zȒ�sT���&oBĢ��-�od���ʋ��	�q�&����)���u�ur^��+3�AQKd�Ec�ӯ��$]�e�i�)�ء6�)g�&֩�N�'�7�9�3�%]2.�S,u��E�	z��۶�&Z��>����J3ʟoK���g.4�LPF��ڼ�)j�L�۠�
��G���[�)\Cu�����OH��R��1B�O�������q5Ik&��gi�L��f!�F��-y
Z��W�>��*�.�Z�G��C�]Ź�&w�LФ}�8b_s�	B��*����7�2dl��]�Ro�zQ��p���vu��fi��˾�u���e[��̭�<���1�]�������V�lo,�!��TI�Ytk����N���3s	\C���wy����8K�볻H-t���B�
���Xl9�W���/��B�jx���9�5g�I����u'I�Z/LX����J$l:ծ2Y���02r���]�h�2���ԧ7dMid%$ث�E�jlk�!f�9�m�Ofp���?[��Ɩ痛��I�m�9z�JPɃ�8����5��=S��y6���o�y�v��w��>fD��j�-i�{�o*w�zxEO��y2������6g��Ϩ�չ;�ǉ�͹<���\�@�,��ԡf߱TR��F����7���>[���KÞ�e/^ B�v���9@^�܅�`�!��x���0�U�y��>�Cь�J���vO���#�z�b7������]1��n���&�p�����k��R�{i�Q)*<�e�dD]��el٬���(PU�Z}xiv��]k2��{2)rI��OzQ�=xa���IT���m���%
�Q��k �t��~�7��3���=��X{l� ��¥���K�Ԑ[�<��u����Z���|�/�������SOC�U�\�t���%p���o�ԟ�!�|�Y]���ĭ
!��|���kqFf*P�,�f[H���Pڈ.�j�z�-��f.�LR���1�:وܠ�G5�<�q�\�l�W�K��˽�ٖ�!��.�d��ov�����ѽ��r)���c��hM���-�[�7^8+������*�;]��z��s�ٹ�	���!]�s%�]*�j3k�w�vu4muUp��S3r`����ܚ̍�j��;n��Vi%Y��r��r�Z�C���\��(�C��Fp����]7��L�'�n�&s�&�BC'l�K9��Fpu�Ӿ�C��v\M7B~�͐���T=%�@�n����Sc��q�pM�����|�a�7JEB�l&7�rEH\2k%�	ιOZL�
���Dj~���p�]8��P;x���xJw/ef{̢ͱ[N�Íwbf�ED��9��E�����*�P�f��Q�,z�k
��H�q�t�����.;�Ѝn)D�386f���=n�6��b�ĺoۦvr"���u�Y�yu�q��a{�ֽ輻�1����#��]��\�����6���f��L�zo��k�~����!`���&��W�����-�{{|�{z;�K�@�_t���כֿ�!����+���c�{P}uO����������D��q[���ʇTԱ��p����~������O�(��>�}l������q|���Y��w�E<!�_6Bw�;L�WL	��ͽ�N6�[��g^TؿwF���V��n����E&��/Sq8*v9��d�{Q��{U�ߠ�΋n��1����4uE�3�{��'KE�����Mcq�v�vd}92EJ�~5�ws��'�_�O!��Xm32/j.�Y�&��N:���Gh�b[R�ٕ� !P(����U��W�&r�dG9�R�X�L���U_[��+k�5wт9��%�r��7(�yi�����8SDx{2ʦ �ji���Y���H�V��:t�3�z��LpR-�`p��r��
s�6�xC}h�p�Aw�{��ݒ(A
��n�4�l�7LF�B�u*WϏ�:V��``5�i�)�Upn�ܘ������.�]^�[^�B麄_�ԻEF��c�
�]*���Ü[������� 1w�a�8���D�>Y;�RG��.g8p.PK�DgK9�r��]IevA�n�]i2gXI�o:v:����K�#�^EL�ʕ�3 ��������A{��F�̔ƽ9�'�WyD3���t�J4^�gQ}�vt�`��M9ӯ�&�g�ʷ����K��:�����
��
�����p�*�9|��Eи���5�
����L��-�e�8��}��i1L�P��Dه��FM��.�g�������eVK�f����G`���x�Np�w�.���f�a��Ɓ/��g�jW�u�ñ��t�����o�NrL��ro�y�f!  r�}�Bq�[z^Þ���]l�{*�V�tu;�=w�4��ܫ��7�W����pdL6�6i�����?@�wG3���/����差DU�(��uA�]Kt�Χ��F���F<h���	�}�4������M}�6ۺ�tS1�ʷ�m�;7C��=��sh�hT���M�"�F8��O�>��OPeV8�&{z7�?F��_q�m���F7DkR�"z;�o.^�����%��a�,��s8)� �'w��z�3�=3��<������9��Ϸ�K�_x8�h��;~E��*t}�t�`�0�,�ӓ8*Bg�+g<K�fN����^��w3�<��*�^�R��%/Ҽ��������8s@�Zv�R���Z PmC|܁���Be�v��	��2[���!��vcp��H]�\S���W}H=�jRњZ��\��iUb=Ҥ�KZ��@j��<�*��!_n���t�������D?z�\-�:���.q)��dx{�v��&_���_�t����n&��7wu	�	�A���s�8Cי.���T�i
p�]D��P""���$N�y���0�&�`'�`�L��EЇ':Z_<q\�}�8m{�Sv�8C+gܘ�7�o�����
��R;�ϧ���o�'xfqz�LGp���筚���L�uc�q�b��kݒ^0e�Fg���q�̤�2+Vၙ͜��*�;9�ŝ�C��Hl�Z-�������~c(�Ƶ��Dk��ȃ�x��ؔ��L�y]
�;�PȰ�Y���֋ʆY��#���EŹ�p΋�F<�8xd[�n�}��T�	Q>r���r�*WIw��7C/~S�-qL��C7]�O�ꑥ�_r��-�G8[tFp
ۄ㼮���u��̞H�t���u�=�[��̼1=��M�/ޛ��k��ciڨLĮ��ۢ9�zЖƕ���Tt�*+���6�S��(������.зr��Lv	��O���o�M��Cךʗ��w޺����e�4���������\a|�m���\�8l�M�b
V���ҏ�8�k��5*�^��P���5��	�uvoTp��n,=ux��0_e쥰>��lU�]�m�x�;�6'C5����+t��\�o�w��\�AW��0���_Y�we����n��r���eS��*B��m��rjS��Z/�z_�Ve@�n~�#C�����v���l��n3�k�[��������𜝔�}OH� f���'t�x	P�vt�<��]u�/�/zd,21�zng9�,I��H�w7�)X��󊙳g����κ�N|@ƃӜ/��<�q���}}s��ֈOm������zu�ţ���{N��ǋ�[�~k[L&7�Pg���p�GT���N�b��jH�q�$�e޼T�Jmm��<bx��3�@�4�J���ȗ�M����=M�J�]==6�l)�2���q��C�=�a�Tк �CQs�F��w*��a˚Κs�B�%��S��yJ��%�L�fjq���e�9�ܘ�]Ѐ
�Cxe�8Hd�s�$�Yj�~��.}8��.��۽��4����!Ί�a��~����g��
�K�� ���`��B�K�s��c9f�>��$�t��������``4ݝP�M�4���ǎ�MBܲ�g�f�zj�Iv�S�c�R��2��n�� T�@��f��V"��6�L�-��5������ذ�����]�W*��tn�
��ݒ2��.�� %k�K�5�}�f���c�c��l��+�h�B�xH������z�}�F�>����hƅr�Vo�Vo06��>�C��&'E�S���lr���d�n�2�������+
��'�����M+5#��#�6����F^�@v�n[�r������-wJ�˫�\B��5ݛ��Ͱ��{�c�7oAY"(��
ۃ�WH����ˮ�W�����S��u
l^0�^�8� _A2G��ئ@Cm�Eծ��u�,u��a+l-�f�K#��g6��FZ�7��}����YQ��s5�|�wA���;m�݄ɯ�*��nN=�A{E��rs�:twT�$;��*��ϟ+��u
���ccկX��Vj���ru��1 �p����k3��huf�_��z�=�a�'�6k9��4n��. ��W5H�2f谳i!sf�@�-������Xg/~�[�1����ܸ��ֈҚ�ő���'}u(���淗h���,;JuI�Ы	��Z��[����e
}�h��qҬ���#��ʴ�n�u��mR�%�/���n
���\�*�u{xN2v�Hn
5:���@{]�H��K��j��]}��F�cH�S��6Gf�.�5�3�s�@����_��
�<�b2X'6��?�6R1W^BTׯ>��[ֶi����Q�v�v���V�m�s�aA%H��
�;i�)nr��Փ���2��/�~��e#f��;k349���T��iV�U^�k+�>ʕ��N��&�`�_�k��u����-.��3�����V�=��J,R��o\�m�;�e�D^)����l�2��ʔV��i��b�i����ه�ފ7k�O.��'5�U{)`�����F�Ee�T�̋h�32�{7��<�B	bU�wY6�&99��ٖ�t���S���>��^�F����{K�̫��9-�ʚ�,$l�d"�@���)L�CQT�-t�A�[�e�\�����*}Sh]�u�M��&U��x�AA]�kq��8�9R-�N�*���WL��LH�W���p��u`��S�h����ͷM��͔��	Wh�TBz��b[ke���p-g�y�¬	6_����O��0;�S����\}+h!��'��ͅl�if���+G�Ho�.ie�f���uIe����9�Y�"��ԏ"��Rd2�EN�<[Fj����3]:�p����*�%ߨ���&M�݂����wn�u�U��4M:(v8/C灺���2Ǝ����Ӯ��֫+g�41�o7u��Xr#Ң�ⱈ�3*��x6�ڵnq� �J�Z���q�W&�\JC����ر�bJ�a�Uc=���:��Q�N��v�h��� P����J��Z_�C����g"""�J�maQZ�r�UȎQA:,����k��(�8YPQAʭ��#��\ ��DN�s�*��NNq*�r��.EȊ��]0**']�0�5hDEȨ��
��E�UVt*.��c����<��F�B�J�"*���UҨ��[9^��z�M*��s:a�H(H�����Qr�
�(�� �QI��2t:Ep����,�H�TqԺ�Q�e%��TWtw�"�Ny;�EPG�����I�,镹���r�d\�\&��EPUQA܄�"�DQEeK+��T�{��=C����*�eD]�k���p�s�e�㰈�z���"�Qf��A�W
&UAwS"��J��Гd����\��v�2HT�����H��W
�^M�&���(C��q�.�R56�Ω���qn��ܸ�I6=���/²���ڝ^rZ�����eg��}��b�o�p�e��3����њ�U\%�L�!\��>0�[�Ao�.��E֞;���C���'��9�^Hu,OQr��8��}�wKc?Et��D� F�']�e^҂r*aD�ݳ�O���l��~D��ۉߗ��ٲ<�N�C��@��#���l��ŻT��b�X[7H���ͦͰ�n��  "5�Ƽ�-��M!pɯ6K,�	�I������_:��v��=n#�y\�"_7���M��zS�1cb��ӳ�*B��)�,1�N�Q$������_#�Z/�~�M}��7�a�7��UoNp��Zϱ���g0мB�8��y�tz�M���4w�HO�jY!`k<ќ9��y��}�K�w�|-�� \]G��Km�[w͌��^ ��&��	�y���L��V[zs�p�3{z���u�M���n�ݦ������ra��<�&�0���麧��=u��,�>��pa_G{�-�L�{ss�^;�5�E��GP��~c��</�q�-�tKf
e�NL�LҡߎG;��R�J��'���/�>_KD:�v�Lr�����պ�A]���1z0T�kR�����#z�rWiǞM᧑��][�*{�%ڮ�Ԇ_�\+�V;ޗZ�6���ѕ�]�>FR�
K�e�I��!��x���5�+��2�ޝJ�:v��뷃�@fά6� �ڼ9� �Y�C鐌��ϙ�m'��.m�� !P(��ʤGR9B����k��`��NƩ���2j9߸����D-��ι͌�Su�p��.�f_� �k�X-��^�9�u]��اwu>�N�#��U�2ޘ�_lMܩ�o�Np�}�xB�ѐ�8.�'�q�]�l�gD���|M�C�sf�#yD��Z�_>?,�Zq��׻4e2����s��Y^Y���_`F��O��w�^~0;��S3��ׯ��=)F��}%�t��:�4��|Or���W����������B��a�Q���
��]^Y��^Z����`��\O��[;���͉N��M���)���(B�r!�l��Z2m�p��xd��Ǿ�<n�Nf��;ܶS������������͟r�X��Z����}�����b����pv�3UuH�xc<���@��.���N;����=�#H�m�b���u���`��Wy�Ğ���t��{ ��l��TٽU�����M��6�z��z_���ȁ�L=뻮�qU�4ϯY��/�<뱯Tf�6sr��jW���G]���k��k��GMy��_����9W��T�j��9pt��E�;Bh�d�;5���}�-�B�`��3��k�ڱä��x�W������q���7g��}�ٳa30C>��5���?@8-�z3���|�l��OD�m���~�����M:.�+��j{�(�a�'�]�2�����`eM7<EzTc���Oϑ�� ʬqlL��=�����Y�����<�9��1o���˗�Q�fktK�,��ng4��l�����<�_��ެ3o{�Vi��Oz;����X��s�6�T��m�9��e�Bg�;]�f�W����B�{澗tL���p�hꖼ�Kl�bS���#�{�x�uZ������b�sXmY+I�ˆ朇]���b�x��Q���J�s��M��)�)t-é@p�e���p�aЍ�3��8��6�c���ri���� ��O�dp��Tݶ���yJj�/�QWc��ɐ�DӞ�� 7�xgBz��$)� ���M9B��.�~N9쀆Ja�{��nȘ�V�sS����i���Lp�P��W�Cx`�]�|����[5���L��� f�3ww����/���G{��+��<����A��B��C��,ϰ�E3��@�v͕�����w��n�U���^޿�	��z
���r(�tkN���jQ�?��Ѷ����
���݂[��"mL�^��L���Ӈ+6�ӬBe,݉=*��W%CO�NۧsW��]\˭�X��F_Ź���vX��)��0�������HdK�s:H����$Z���tl��|�uMqw��>y��� N��ٷ#
�ۏ����;f�^{�4�kǆD�
���Dg ������fzE4���cL9��Mbi�g�������k�:�B^�&	���������WP�~�g޿!-�,�^ø�Q�i�f�8#�bi�d�%>�~Q�;��M���?j������j��ʗ�����0D�x�&��iͺ9�l�y�.��ܮC񷍠�S��+���O�95)���֍�����7:�u�����j���ɧQ��C��i\g" ׸E�L3%�4��*>ijmO�.�_S��v-'�v�~��X��S'�R�-��y��M>k.��m��N�|�����맍�w��x�:!f��Ʋ�wP�0sp,��cA���Np���-�OJ:�1�l�p���n�pUu.*�k���$��>w��zf��+w����cz�{��p�h�|�n�8��ԑ�c�N�q���PE��3(�U�؜|�q��I*^ȗ�M���#��m*yt,��~5-���}i�^��Eb�Wۦ�0�kק1_
�ts�J]����ө�gB:2��RA�f����TB
k2�b&���+�|��Vݬ�����ʺm���3dY*F�ߴ�+5:��2���+i�	u����]��n�Е����P ��j��c�jI�~�W�=��� xCQ�S�LGR�ܪɇ.i���X��OE �nD�o-�=9'4�t9ޕZ�@���L!M� ��1g�fYSH���P����uwTi)�&�T�u�����W�O���~�>�@Uj]ܨ���̰�?BCuf�V(Ј�=f�wK��x:��{��ണx"8�cz�a��4��?F<p�Zhr4C�:YкI����ѱU�[����h�	lU���
ITf�h��{���zfxK����.���8�"�Wj�nwY�������
�Bm�s7�K�\���C��Fp�-������z�Ǩ���*�
�|�g\��͑ݔ*?F��{q;�x|�d:yӽP��I�f�̌9�5]��f�w'Z�����(���b@�,Lk�[9"p���e�[:�=�1]ݔ�v�Vn^f��Y��e8��w���D�So6U�<�����������7L�O��։�L���;�n�sT��l����U��
�~�M}��6����z�緧 �+����E�t'��0�
��أ��v��$�����u�.�Yi
����cV-��k2Vh|{Z�5��I�5��Y.	���/���	�A�R0�*=D�t�8k��ܝu�46������7L�-CJ��0�-�x���Be."�k�t���@�?K]6���j��$�s�i�@`�`��5-������<Ӽ/��<�m��������.,��y������|I4��<Π�W�-z�W�!;ǚ�i��4Yl,���#�i��[��s�Ȋ� ���:r�|=(s2��7m�Ka�s�4�NC��N��S�c{U��YыP���i 5�fiq��(�H�>rɒ
���tKf
��׮���ߐu���|�8���m�ׁj���<t��f�i3������-����j\�� @<�"6YC�#=!3�5�xb��N'���+��1���}.��p���ȅ�_T,���L��	�� ���e8,۰L��"C��_u��K���o�ruj�S-귥�1�H���i��Sv߂��������iZs��Z[<f:ec�y�1ĳ�;^��T[5
r��R�|~YҴ&��vh��<�]Og)�К��gֻ��Ԁ���~�;�0�<"�6��m��)F��}%�7 �l�.��	�QW͙��sF��i�Q0�z�;?*g�r�K������5��}�>��{ ?`ԥ��Ze�` �F���4�{ё{9}h��ؑ��"��[究��oF,;�w�!J�{�ZȬ;ʝ`sjp�k6��U].;rd��K���e��E$���ٌp5�om�gc(�Y9�O'm�����f�6:�[���+���a�;�NF,C1�=����:��]M8�fr ���!�Z2o��s����q���飛1Q�ˠ���q��[!8�,��R���j�2��GC���
O�]]x?��ܛ<>�#_lsaxc:v�#�wK������������	�Yj�c�wmV��v��rwb�������=O��p�sz�SYM=��9ƞ�{��|�kU��֝�� �=��"���1��oZ��	�}�4���=/��xF5e �Y�վ}�܆����ڄsn�d�*��l��-��02���*Tc�����?��5U�+�E����̒��r�J��՜�w��2��I���tp�;���<oM��b�u�̌�.��!�G[��h���3�8P����p��q��v�z�L��v�ϕKϭݵ;�K^ V � 3��b��C��H�Զt���x=�B�u��Rז�m�HYϕ��"������gv���>�p|�V���s f�s4�tb��P4إ�����J�s��M�!pX'�6��t���h���īsז�;�蟴c9���NyK�.�!��y;j��F�C�����ʰ����YcU��m�H��YyB������ѯ�":
W �3h���;QX]HY��;�ުI�D�	���;�o9�w�:�=u��RH����}��\&��~)Ot��%��ix����y���Gˆ�m{����ƛ:��|�U�7�#��r��йkLWY�|a�	�`V���ce�`�*�Aw�8���$*b��TӔ)R�Ƕ���h����O+�;9���\�kR^0S7uu7[>���P��W�1gu��L:1֋��+;5���f
�n�n�sl�Vv�td�7�ރ���3)�tDt+H�V���]T"��,���v���ʤ���y������y+���TH@^�A{�gSwuC�7T�	�30׹T�Q`;�q����D�6��q��ҽD�sGz!Z��Έ�5��t�;\E�� p�����z��>,]y��*e>n�Z>�}Ӽb3���x��}�B^�����l��Y�`:�ӵP���8_Ds>��	legb �5�v8��=��~}��r�T)��ߞ%�{rm�G`��O�͝6���&��ʗ臎���Z�Q��[MaDOs��ӂ���,�ܮ����~6��ӳ�)�B��{)��&�;�Z]��]�`��ꡙZ2�V-#f�K��E_M?FŷtK�湧�,IN������^��m�i:v��n�x}�t����k���<'f��s/���y�V��G�����}�� r��uG]�������'��)d�Ss�f���]��V�m]�|9���Bw:���K�x�Թ��qK8�"1� 1.�� ���:r�u���ۨ^�������S�t�*�M�>�����.���T;���<�o:��uMȮPX�� �a���r�&�麚��ga��ޑ�
�����*��;��|wL��sM�|}�����D��\W��ҎP���Fc��/�1r1�z��`N��[L����U.��|�n�8�]]����Ő2��p��{ޚ�� �$�m�+����|m�҇�+}t����h�SˡM�=�"�֎�t��Xט����᳚�%�$_�� *�D��)���SJ�r��a˚l�V���T/��1h�[�8���B{T����+�r��&��@B���em"1���bL�IY��;N�,����oLݰ8�[-��E7�O���\�l�W�K��˻Q���+�ix�猑��^����#F!mU���Q�iF�Dg7gT>WT�
��1�5��!K&��==��v���w�fz�ggӰўqݱ^��~�*�j3k�gt�:�6�����Eߚ�\�;1y��Q�4w�hw=^xw,���5N�p���R�OQr��8��m����9.�=i��O�a���b�<��Ԅ}u���*
x<B�0�2}�)n_���cǯPWy�#.�RJ�#���qi1:>�X�3w����X��5.��� 37;��r;Uo�.�J����Y�N���-oqK���lwa�|3�*z�4�Y;e�u(SK�����R�V��s��W<�u�O̞H��P@@��@��O���~���u:}hm݊��~s:.g38�+ ���ٸSc���a�n��T�K�F����`����;k���OzEUo-�ճ�����'��SZ��]���98����e3�1龘���[�~�����XL�F�qۚ���걒9���[&��4���*]�5�K���uK�T��7>XJ�+����q���V�/v�r��*K�Lv��$%�jYQ1=���Fp��Oߏ�_{������-�M_�~��j��.3F˺�3�c�f��5���5��'�2��[ռ7�pͺI�[E<���sנ������_��ʛ��uaY�!<X���4�'�,󀆧��C;.J^^3N/��)��6sMWIQ�b�i�(�=y��ԑj� S>N�M�νo[�o���� ���j�6�M�����;�d�s�q3�E��Hr����Y)�L��� !4
!��+�A� g
_^S']���n���9�AuM�]��B+�K�r��7(�-3���p����n�)�A��KY��
)�)��@�5{S���of��d��u&���`��F�5�6�p�C)�K�\u��/HJT.��L�T��l�"&^m	�98^]��:N��3���l��3qk�n�ݒ�~n�5�c��R+���֩�v�Q�T�4��@8��T�Q�3码�]�o8��_h�.��$z9�!�j�U��N�]l�Y�oj��m<Y�m�d�Qn�@cԑ���¹�
�]�
�y�id���r9��L[��4B/:�1,�-�pQ���Hv���doa�9��]Z���;r)n��/(�(w)u[Zm�[VJ���y��y5���z��W�T\r�Ν�V����ja#Ó�2M|�i��eҼOmiꢯ�o
�Q��%��Q\����W1WN� u��V o�m^��!�%�tց�AwkZ\��ҹ������g?��S��Ύ�6��ru�	ݰT�ApGL�nQyv�s�RԎ�H�/A!�)�.�Ӄ����$��tn�;Krd��[�*��)���L�_Z����ڝ(�9(r�ڐ��X]�a���\��Μx��2�a/3b*�.�/�M�,8{m����͈��_j�ƺJ#zذ���ӛe��]_>Dm�!c+�]JPd�oJ�2|ib����Y
 �)Մr���5������������㝴%iw�l:�V�F�[5���Zvr�+>� �O�����%I.v�;�Jr�y�g��g4Ŗ	��5��V*]�NL(��!b�`2���6�;%7����d;���x��q
�wv��$�j,gJ�R�ޕs��ܘ�i�Es�ݣ|77���#Jv)}S9�͌H�!A���<�R�ۀR�-WfԤB&:A[�A�vJ&dil7i���mq���r�x�Q�H
hk��{�Ӧ�[�ܬ@�g]�Q�/wKc��fƶ�3̍n{3�=n�����Y���Kmsַb�c��Zpã��f:��m!�p+��Ű��:�p��bͩ�ڶ.��]�$I�PkZ�9��X=�?9\K<N�*�"T}s�҈�c`V����Rkc;��:M�vN�0��	��k����p����>M��KC��D��պ��cxJ�q>o%�m8M�l
�m"hL�z��M��J�{��pBdx�8��b��͹G3Eѩ�]:]��1ї���B��o~s�qfb��T����t7o�b�
# Iv�E͊�/��,A�S�{�w7]��$��j�].�l\�/�q�,PdJi�G4
��,�V��\��{�\o%`"��6���.��O7����lc��� Lj�U��i+C��gWac-+�7�P����t$ofP�x[w�j��@��nBYͫ�$����A�>�IV+��	�ԅmn�	�9U1��e�����T���n�wb�
���㻩V���i�,�սZ*��rX��ʭ�(�_n�Kh"�ؙ����:��n�ʲ�A�e�1��v�ԍ���� +E
����*��uT��gGSְ�p��E��Dq�璒Z!���e]�-8\�g*�p��6����r;9��9"�g,�+��땙^�hbE��6�Ҽ���E\T�#�T�p�B(5�Dey9S.U�Ѭ�\�QL�K�Ժ�\(.�X�;����$�WT�\��g�.y��
��N�P'5�tP���8��E�(��֣O0�3�jy�.M\<�ft"�'VY�^*A[��PTvUI*W��k�9Xd:��ć;���ʸ�*�����%���+�@�b9�;��랩B��.��H��R�Tr��$�	D�BSS$�]K2KY�DwP��[8UY4*�rB"<�9A(U�fZD$Q��I�ٙUH��	kw
w\��x���fN����m��]��w�sH��u��.��H�5�T;uQ�\� �}˯H���'~�ޜ����U}scͷ�2�l�x9� L7�;=��� �Kz���G#�3��Sv�9í�1��V#��]\K@�:�'���	ݬk���M1�[5
r��+�Ƕ�H��}��c��=�t�z_c.��D>�k9�r`����z�AwgX��`��pP���ۧ�R��(΢�J�[D�����w�@�e��2��]+֡��W�ɥ�d��ܫ
���a������s7�j�6w;p�N,t.��c���:�M�}m*"!F{�P�������FI���z����n''/R�:�?v��K���8��Ż��qJf�a��F-���E�/�L�h���Q9}�04��nlv�R�v�3��K�]������a���Sqgz��޳�q�[���|t��<�5ӣ)��C���/f��oL�m��z7ts8�=R���֞U;q�Q]���?:��x��F�g]T���M*3�߶�Lӧ�&{m��?�j�	�|b�e��������t�{�2��\���`eSs�T��u����\~#�4>���w?2��V��xEha��� ]�Q�V�Q�{��{��}�RY��;�m1c	��7'^�>�ߦeB�/)"u�Ӟ����؜Rw�q������&���L{���;w�տ��૫U�0��<s�������t��A��.u�4�3,�۴3n���ܼӚb�v8⧵E��K���+ߓ[iW�lEU�6��W�V��+� j�)��5�����$u��W)Ǧ�3������<x�=g\䍶*t}�t�`�YZ��y�C��&e�g�m�ݢt����#��6g3�]��<�O:�q�-yl�m�ģ$,��B	����z������'/I�/���צ �ji�tb��4إ��GzK�p9=t�o�N7V�H�|URѐ������89�o�8�Ne��SK��qQmB�Φ��8��y��7�6�쇡MjݬF4�sQĜW6�xl�VϹ1�� :�xgBz���4�=mSNP�K���ZB��I�_e�B��6�$�`�]]Mͷ�ڇg*�1g�`�]߂GSK���Oѧ�������^w��>m���z�.8�+�>^����O4�Z�^y ;���Q���1xy�˺���gr�3w�zlG3��E5��*c*���9�F�8�����5�30��Z��U��B���*�'y޹祠͎ygZ5��)'k��������o��2���쬻�̿]�gN+�,�W*�רg|�M�m�=�J}-���a��m�:��Y�=o�-^�7w�1�'>���vb�IUv�{��T�3�7�-'�p�SWz�N9���p
§6����������ٙ�+cK��Q��Al�"�k�j�=ke�Ř�n�n9�o���6D��t9O�a{Z��{ :�ӵP��8/tG3�Y�ۜ.\��r)��#�=~�r�x�h���ǹQ�&�!>KgM�={I���ט~@"�xlu���UQ΢:�9�zۅ4���g�r����?���n����R�m���-"�SM�VFI:t��[�Q8;ؔ����ؾ��c͔�\g" �~�8��׍j��o�V�dE�%�w�;��n���4w�$'�;)��fVz�ogL���l��]u�.۔�3�o��n�+y���nz�#b�f���3��� �w�ޞ�m�3ϧ7��Z�/�|�g@H��F�n��oO�ߎ�sr���c���	�-m0�F�j�\L'���	��؝��MQC"�1��B��w����\`	[tN>S�#��"H�P�l�~5����=mBT��rˬ�bE�b�C�LiSo��,���jH�p�	�I�e<�cJ�r��a˞�s�:.�l!�aټ��4j:_���$M��~6�ԟ��Y%վ��� aY�Y����?v�Te7쭶�;P�dk��ک�~u�z���w��j��/�����ʹ��� ���63�����50�-eޓ} ��G��ue���v2n;�Χ׋P���:��Q�DE��B���5�u6��6�K�����B/���Ý1�g7b��R���{�_z^psTA~�v�[�-��b���S��~,�S5�wr��w�k����yW9EV�9��s��)�F���AuM�J�J7�#�4�vuC�{�i�-�b��ѣ�E�
4N��OB�!�C>d�Ϝ���VƳ_E�R�D�B�{n�:vu4ogLcsZ��{n�����2��j���X@r�}������s7�I=E��(�C�a�"��M�WkbS]�lJ�Y���k�bzEA��(  T}�#ۉ�����c#��+Gt�}�����-1���e ��G;�_���y���aL��T�8�a1�,�H�\.y��q�K�?>��e�i�k�ǮK�7#5����w���=�o6S<��銅�[�~Ml�7��	'����D�i�
"���0��z�E�
�~�^��w�0��bN��@]��g��df�Պ��ԳN���{��O��g)����>ɩeD����a��y�<�o�_N�����$W��=f�´�!�POˠ����}l�&/��J�0'z�N6�ޜ@d����MB�@v.أ���f�z����p���;�F�_�����x�^f.���՘i��TT��#��j�v^�ҭ}Ǳ��]�f˳����\�]��"/��}yE�q��^�c.�J�]�����]��i>=� 	�w4cK"�J�b�y��\M�;�F��޳�c���Ђ]��V��:�ŷth��ar�'�M��Q�6Jw���CKHd�����VNi���Oa�f�~��<g��ԑj� [�+0�ʽ�[�o����/Y�;3�s�����w{殗xD��ҧ��=V��|���rڗ6�P
hD���[.�/��<dims�]��V#��C�#�Ȅ�;�QBJX��F酔^���
��8eR��xg�_l��̾�+]��%��#5zg��t �L��ޙoLpR/���M�l��7���g96�nDLT�7L�ĉ���#��zC�^]�ท	(j��z-�S��W=�,�:;��q��ua:څc�h��k�%�sFqڢ_�raL�"�:��C`��pP�k�N�/}׻Qn�3��e�(�v�:vu4h��M5�]*�;?*�<;���1z����}�쨚���M�8J͙Ƌڌ����5�
���zn��i�S3
+ܢ��܌�-��n���%��6o+:�PΚ<�ċ����(	t��N?8�Bq�|��(��ƃ2�c��h�\�|��sOų1aj�q�bⲌ� [f��Jι��J������5������ت������^�.���xܺWkq#�#5�=�%MJ�e�*xneu����涥w��E-�4���o'�L���ٛ��x��Q���\��+h��Xڝ��Q������C�{;��2�˃���:���K߂�6ӵP)���@�]��l�㼶���FX���2o��t����3��`���4[秺q潐�dL2�ު���e4�
g�| {�7�1����|W�O��i��"�n7����i���Tg�l'��Lӧ�g��jrX[�؜��~�ԄT��&�9�EX��ʚtQ�ʷ�;1)�\�g��ʚnx���+%?8��dv�[tN����I�~�&�ŷ)[�{�/�c8S�.��{�nS�n�tK3%�M����rm��EU⬾��Q��K �A��٠�|�}�=���X���8����F	�7�_�=���^�n_�/��&�y�6!i���L��;�'��p��p0�}���bS��T�s&��V6z���3�(P��'ޘ�a��T:1��g�S!�PP�f��n<��%&�茇6V�;lsn��$Z�!�q.m�A	�/�1�D�ru���� ��g;�\M��k٧I���O�8C�k��/CgܘB��� :�Aw�3�!=LBB .{|�4��z
־ךLa�c{�YV������E`A�K�6Ȼz�5�����xd@��2\pjU����uѤ����c��Τ7D7���蘳{.��B;8�+�Z��49FZ[�ͺ�K;�ЂQ��.���6P�F�b��k�ݴ�[ET]��J]�d��sQ�gp�9S}o�^~��i�$�`]=-��&�kP��W�1gu����
<���rV�U�^bC;�uT2�t��{1������Svt��7URy]�P��@w w���狻�;Cb�q&����E���:�W�-��z��3G!�ѳ�)�����5�k̦fw)�5#�4�d�o����辢@�U	'Jls͸�%�x��I��-Dq��Fp
ۄ㸮�R�]�e�4l�붡9{��_��%��K͑݁1�O�ǰ��^���4�T�WP�����填*�bF�(j�b�g'�z�z����]��nV=����=�t�����[eZ��s]]%�{��o���)u�9�8������,��WQ[��~7獡_�cA�����\��%#�W��W������T���Q87
��}4��藗�V�]���%�aqӺ�ה6,������z��I��#�G 0c���r�f{�=.����3��:���u�H��!�o<��;��b��/^l�p�~>\:�ng>�1�&{�Y��;ףz{��wL��ޚx�5��*h"���h��M-{�z M����y���6���y�F�*]"��[����bgky����JvdD�yɳ,<!�դJ<"����Ovw@f�ˡL���1�o�L������ϐM�s�}�t�?Ȏ�.8D�.湉9z�J����Y�T�?�4m���`.��.F=zT?�	���	�oV��pU.���ܡd?e�=��q<].�GVrڒ-\`	_��q���D �m�~��T���=��'sQ���L\��GI��
:)�O��!�rڒ-\'u^�D��)�#���ۆ�q�GF��|�<�դ�Ov�\ވHO7l��)�@W�3�L!M� �1g�2˯:2S+`{��Ia9]:b1�f���^Z�ޖ�F2��C���}��~���
��K�����w3�i�PXEfY�j��\0l��D!�-����J�J7�#�����SH ��se���|l�z[�l���?J#�	[��i�h�pV�5�[�$�,�6�Fy���+l��N3�6����6gP��,�ޖ>�m�Hu�@E@��.[��p���O_3U���w�Y:�6p��\,X@���mg�龦w^i������`@@=v�{���	�љ@��Y����b5Mˤ���9�z�
lw����EOH�A���1�,�k�c������I���I�w��G�[:�]�Q	]G������o.YH���(ձ��( 8ߊ�ˢ��>�����w�_>YW}�1j�<|���R��[E@iN��zÈiiާw%l6����"[�� &�8��H��W�z�;��fTAC��T����O8�n��}hD�o5�>�銅�E��G� ���n�vt	�D�s��ޞ���F���`���TٽU�ٰ�w���.�k������*b�2�B`���2oӊ��Z~�e����m�i:m��Rʉ��m��w��t�<��U�C�F�i07^����s�t����q����CV�]5����sux�K���e��:�L�؜r��h��q��(^#7�����u�M�n��7o����OSq8*Ts�M���q��=yM
Hѽ{����#F���Q�~hR���S�l3�^�[RE�\`m�%����&H�]3��;��n�3�wu	�y=���}�.���*yY=V���%9l�.m�� !M�>�;>�a��o/�̔ǽ"���VDs��)w�SE2R�l\�)���.��HF�c-n��x)��kL�K�'����1��F�eIB�A
��[ז��"۶�7r��͂���YN�r�0o'���!ߨE�Cy�d��\�%L�OD��Z�_>=�ޤF�Lh�i�ˠ[�O�72�s,��TN:�Q�IU��ͷ.��M�N�f�������q�����ut@R�.~WM{}+�W��n�|<�k/�X˗�����#3\X��k):�_@P��� �)Aƻ�8����j����gi��ڹ3�4��F��ٜ��s��o�Ä��i�;�x7ܘ�i��DAw�p�;��<"�ࡵ}6��6^gw4��j�:7�9�r+;]3����t
�gSF�n�T�K�c�5�v~T��]�C��Z!���y��vL���9V��5�A�囻�B�xr�p�|���]�+��DD(<���,#)�SŢ��5��^�5}�.y�x��N�@ԺK���8��	�y]u�)����Yi��:��M�؅��7�u��9���}�O50���`�g<2�iڨ��@+�]����w�U�dm\	�ʎB�b\GÈ�G����gǰEa�_)�FU?|�晲	ɩeY�U�����r��i�!��n5Q;¸��y0���/��[z���:��G�Mv���o�Cᒵ���4����i��hu^:F�nd�_�/����z�훎�@�z����W�<��Vx퍈�����y�I��L%�=?T������qd�oE��K�������{����aa�!�6��N��]Qj��Xv����VO;���|f�3�=�O�-��{A�Ʊ鳮rF�'��!Vj#����e�O�/zo1�;�*�:oh�]L�Z�Au>E�\rX��7V�8R`��Ĝ`0��/5�ُ0���vMr�����OX�w�̤�y\2�O4���[R��m8C8�:��5�r�4c�|�N��� ��^�G���sӽ@����η�W=2�iQ��x��i�|�ۜpH���θK��z`�;JN�G�m�G+��v���c�ى�(�6$Y}z��-޷[�Lm<���.-p��Fg4(�p],x�N�M�]��c�ul�c5�@�[������?�RX�M�n�Y+��Ħj���-'�3/�Q[Am��ŭ���(��d���CCCQ�΂����u��{�Y<'�k��+�!�B�E�ͣ��^��*�8��%w\�����O��4�u�W����rXX���Ȝ)��I��4�M�G��,\�.+5�̕� �ޝ�V���_n��>�e�n0���P����z����������=����sa����[����+����b缊�+j��.(�:}$O����Z�N9��4�&��nk�M偨:�ٳ�8ө��dV�Б�Yh�o�<�ت؂>\���ݜz�)���f��o����Fb�5n�ߕ�H+��}������U���ʀRZ�{w��ͽ�V��{��ӻv�|{n�(���Q[�(�6p����b�.�����W���*|8^�t�Ӧ������Y�V���	���t�ډ�!5Ĵ78v[{iKO*�D��])d[���ggk��T�ə�]64H�+��<��OЬ��-Ti�^�S[-1�V��C@�����Y�^\op���ت|;�v��hN\K�OM���$Tz^0�j�7-_;���v�y��Y�n�75eo4ƌ���WT;�Y�t���N:G'x��{>٦Q�-��f���˝1J�>��%ry��y������$�a��L�A�v�zh٧R��h"�\�k�b`���]���r�G;{�;�3.Q��p���-}��3C�})h��d=�ͳv�tS���'[��.�w%>�gB�f���T��zg,&5٘��oU)4;[���)���%���L`��ӔJ��Cn�inSh<��-e=���T�	r�m>���������.�\R8��լ�pɫl;o�eg]�M���<dE�:�D�sj��Ԫ/�C[ڏی�.=/6��cF����Fn���@��ӕɅF�Tx�5t[V*��n0�.bQJ��R�������/����9]��Z�ұכ�9��b
"��9����t��+=Δ�0�n���hV�(��>_�]�m;����M�G�,*ʳ��Ul�*Y��x�_m�a��1}�ҁ)�������9�f��L��5|��%
v�s��X��eV����E�+a�m����+����т�ܧ1��,��* .\�#,�աQ�*8V��UЍeU�]���#��*8z���9ar�+�$\�I�C�,ڭ*eZfX3"�\6��r"��g	�Gi�I-�\�V��T��̋�B)3�iK#u�!��WQ��"(��R�J���8�Ҫ��ͺ�QĒ���H�N$b�3���FFG
�)$9I��9�r59AEW*
%��(�(!=�P��,�%=��ʼ�q�䲎��MgK5+T�5g �eW0�*'uډ��4EL���UuUT40���^�K���������u�+������l�%.U�����	D�2����*�٥^�GV�V�W�X�^zJ��Z����W��ꆢ:{�h� ���&��FF�G��"�22X���S�HV�(ue�.��^pe��7�5�59��D��]PO�� �u��G*t�Aԝ�L��dR ��w���mYDԈ����vJ�1ɨe@ٝٿ����mq�{�e��$o�&s>�.����<��:��--���^���y��3'����Wވ���Py�*�~Cܴ/�M�}kⅥҸ&�+1��T��-�Ak���y�{�6sBA`��Hp��)̳�!=4����1�E�rk����ou�-��쳲�*�8L݋��ͪB^�Tݶ��Ϲ0�3wB u.��,������.zg�(���{�5Z�;N�][���X�����f��kݒ^0R��n�}Ʉ*�;9T�+�#�`/e?"O���x�ٛ�|����k�U��d�����7<�C��Θ|��O4˦c��wr�[⌗��r���z*���7DS�~�W�,��Q!z9qL��P�]S\%q�`Ԇ��ȅ�滦ε�w[=��āʇ��iw�s͸�&�ᔱ;\B�7Dg ����a��¦ƻ�k�N���͑/]3*E������4yO�O˴��^����9�U��v��k����;t��M�&�͑Ͻ�m���;�랐@~:�.���e��g�4��[9��:��9�L�D���'�[�N�9����ʅN5^+b��=�}L��U�x�fY���⋫#���� W(>���f^8�gvH�TIՐ��hk��Lw_e+�ޫZ��c����X�P��B��x�#�DU�z�Z�a��9%��B�x��ӕv����-\Y9���xh��0�iK�E{�9�zЦ��͒�,ܮ�����h7T�� ��kM�O�U[���c����ĩ�z�WD���n���r��."4���h�S�T:a�N%uiF����I�M#��!-�����`'��8,�x7�V�^]u�.�c���ZעMON��U,�̄'�#E�`�9@`�	���,��;�A���3ϦU��ֶ�!T5nh��j[�OC�ȫ�N{ `�S!�Y1r1�ҡ��`N�ki���j�_UČ꼃��Ei�=Q(sFԧ��Tp5g-�"�� ���pG9�ND�R��5�/��Z̎<jq��,�oNn��&��ߛ��m�*R�Y=6�m��!�,� �� NH�0�)�#��3�����d����V�jy��'�0���SO'����c�?h,вK�}Ʉ)�� �,��{e��6�K�F1��ӎ���F�sqdsLF�! KӦ[��-��B�	�u�:����@hkOB����x�m#�{'�xv��|:;�4�!p���꼩Q���B�o�BݿG�_,�YF��%u�G/�B��Y��꿇�ˣ���ͧAl��YNk>�(]2f%���c0��<�������@g�H�	w���[ze�o@?e(皚�$]'��Y�ꛬ���T�i���# ����w{W:�\:��hJ�����	�6bx].�����#9�#����p��d��8���L�
د_E�S)THk���'��1�z�H.�g+��bTѴ�U\%�DBɡߕ<;�g8��u�s7�b&:�!�&�f�8�J���T���������t�^i������g���~>�;mI붽/ݦ�&�5WSΘo�w��.�[7�}�d)��uu0�Su�)�ā�<sz�l�<����I��� ��M���OZL�
k*y�W����rqy��L�Ǧ�`�k�f�����q�]����8̎
)��vs:��o�,�7��_��w���;��1Sa�ND�DU��&�LX�t\�ѯ�L��4��0V�[&��y���m��w�0�8��#�][P���ڢ���*��n�o�o~�@_L�2���5��'u��Olyu������x����t�lY�4��;z'��ޫr��ו6;���Qg�!=3M��J�pP�*�K�Zm��u7v!]Y&:���Ҝ<��[=��΋�t[����q�9mI�0�!�Ã�`T�>+�^��<	YCm�'1M���ܖ�]�ڷ�� ]�#5;���ܭH���/���}�[�ٲsb}�i�5����]]Z��_�/x=f��7��tC�q<�7���/]�N�j���n+wɔ�wt�:�*�H�{[k�u���Uƾao3�J�%'N����!ߺ����qC������<�,i���崟9d˕P@.��������k#9i㣘B�0�P��P���4͊]��B))b�-�NnQ~31XU�<���E��&����F^�H�f˞pS4Aw��-�1�SL��-������2ޘ�[7l���;�r!Ii��i9��*��1�e�/��{��Ep
�.������z.�9T�_>;�mF
Z�'���8ҷ2֫��X;T�4eyu_ƾ�Z��z�뢸@�H���lࡩ���9�H̄1R���D�o����E�3���t����L�iK�c�x�z�b��z���{�e��7=y�ӽ6#��^�]O�.YFN����7wN��M��ה��!��\oFW~�{՚���r��Ƒ���x��I���Iq��o�8�8�+����>��Ew@~�o[VOI澘�|�fya2�,�e<���)����6���H\~�]�_�	|���S�n��8g��y�K�y�)�R+�jB�K�B����^ʧ�ck�kƜ�N
�z�?Vh���mi�J�07��r�E�QeLX�{%��:��)�����D7���r�wG׃�'��V�,�Q1(�z8��QU�]�� Ze�{�%㕊�ӥ��D��*�ut��P���!�J�H4e�qW�� �q�ԨeJ���h�+�!AV��Қ�9 �o��5��~���X�����O����c(�����[]�^�Fp�m��5�����TmWQ̈$�ӓ����J�kĥ�"��+�m�u4�וo|vbW��O��M���tN&)�{7qFFݛ�[�@�q�ҝ>F�|f�*�œ=���3�>o�^\��)�7m��XX��Յftn *�ji�ܝ$��l�2�H��d�w�k�z�3�=�O�;�;�5�Y�9#p��˳]L����s�g0P���iɜ���[�}-�]��<aO:�q�-y�S�3�T�P�Y�\_S�ޝ��}y!mos��T����C����)g8�8C�ǧ\��3����;����y�]7����x�R'�������L��!�9@Js���w�fv��4f9����מn�6��Sv��!���L!M�� ��8���$;I�K�n��
�ø��t����ľ����X����n�6�$�`����~}Ʉ)�C��L!�>J��:�'���j2*�x��w�P����D�c�d��ߌd��]!��f����O4˦c�ڣuH`tZ����q7&J�G-:��=C"v]��D��Xt�دl���*�_K�㐾I���ea6z�وU�v���ҽpݙ���K�](0!��c�V�$�R�%�lR�ܝr�Z���K]ʶ�tɒ޺�Oe�AW<!��Q<�	�z�K&H��]�G���gm�3�X*�#=D�Q�������44�/|����ܯy�:1���6т�޶}�H�z:D���9T�]��)bv��fQ@�(oWCL�%�ꯛ
�� �8�-�7�^���h3!�a��7��J��k!p�f�uۏ�'O�Q��5��ZalG�;�����%��˥�;����3!���mYso�ң�H�y��wS�;s3w�[�oM�z�j���T�DWts���ӂ��%�y]D	nW!��3��n��ܕl��&+[*�sx��#�;o�%���5)���z_�_D�FF�D����j�oN���_p:��I�b�mn�����C�)n�������{'e=A��OK��Ι烝4�ZS:x!7L+���9HE@qb��21�.#3��L���YT�A��Npݹ�Ľ�w޶�0ύ��}��rt�ڪ�}}s��[#Fڙm��ɋ��^��1ӾZ�a����D�]�6��ٽ�&*;03�4.�@t�=�t�Y�jHT,�E��G=ND�:g7^��d͸�I��ӳƅ��D:�8k��2��p^�1��|H[8iY�����W�;W0yY篾]�.<}�N��F����7�P� ����r��}�PL2�@f����m1Ӂ�ث��m 5#I��f��l1���{��fHg������<����Qˠ���aNԹmI�p�
�CQ���ǒ��D*�k�<�ń��P������b�y�BW	����ԟ��Y%վ��� Q�gi^N[GAg���<���;%��D1	�u�U[���d:а�|1�\�z�u�����ok(�N�49@��wu�� �Ǟ̰�P��H�j�.��,�{��^��ғSn��a
�J��[U*�fqq=�18ou��!S4C��Y,��OCE3��*�-���Q!���6́���~�Y��2x��Pt��3�]2��C�~G��,�Ѫw��8Ni�� �T�6sz�;�Jju���hp�n�����������iLOH�3!Ѷxw׆f�:R̋����|�#��*7k��9��l��t�zfK�����9�z��6;���aJn�EzHDz��s��iVq7�O�t��5�l���r��I��eG8��N�!�[͔�p��0�Ӏ\
�~û��c�6)�X�L7�[�G�?h4ǘ�zv�i���xT��
��K��s��c��v	�<�[��n�:�N���bP���[�T^��Ly��,-�3���Yfi���v3���
I�+]���@�?��'K��n)3'�:ǧ0��]ki�1"�=O�<
��v�	�1��ӯ�kK�NC������Q�gCN`r��3�\����h���_�c_�L��y����dԲ$G`b.�<� Fs�K'�$Mu]�7P�P��/�|�B��qu��s,��1zf�W��z�Z�1�\rˬ��ٹ<����0�J���D�Ӟެ7�����P�2����x�]<OOdV��7�:x��n�������������S>�����1�<g�9mI�q�-��l�K9��%�iߣ.��̥�ng���L�Ra�f�N�g�ǉRxE��O!�'��o��zl�.io^�~�V�C}�qC�l���%���~U���g���ڇr��L��[Ҍ�;��G(]S;Ζ���P����d�N T���̲�4�S=%	pB�[�n��8)f�,���i�f��)C3MO֍7k�_/��Z0"��X.)��%M1�]
r���cc���*3�g9S���p���``5�i�L�n,��)�4;�B�3����n��:�a�Ȏ�8k74�t,�S��4^�gQ}�wI�)�:�4SuR�����Mj��r���.�z�F�P�u2H��þsV�L��=�3BWCq��-V�;���R�v�xS3���B��:����|GR�{π�����y�eb��S���R�]�,�����Ԕ �*���u�%��>'n-�*
���E!�/��	��E'�ʻ���e��O{�������W�6�\�����Eи���k����]|����^B	�/�e�Y�n�V}��W9��/�>��G�Q��k���*�	e�����^K���n��:��������^e�_�o�߬��U��g� ���|?C����K߂�:���ap$�]�l����a�r�qz�w���:��a�<#k���`�ê^SN�~��wZ���^�wH�ЗV!���eu��-����&�����׏T�V��y��ȁ<�[��οSL��p����O�msE�͝�<���f��l,��*_�*�+�m�SN�=yV��f)��KAV^��;���{*����얜�����t�M���['e=A�X����M��/:-��u����������`wwU�MΉ�=�K�0���cM73��#xY)���g����~�)����{A�Ʊ����ɱ�Q[�;n���+��||؊{1W,K3�<�3������Kι
.�O���TI~�����.'��Fg�y�x;'�No�l%�.�_r����1X'��R�=�qܝ�o��:�Vʢ��{��K2ﷹV޷{0Ĕ��QӟL��;��x��4&V�u��T��\�t�%�o�R����ཡ=�Ik�޴�լ��jۄ�9З�7��Y�0�B��ڂ�u��u5��\�r��I��*��v�����=꺞{�a7����룗B�������6���rz��0S�W�B�<-�ԇ
�E9�8�������3d;�n5��9"I~7�Φ��#��Kv���ʛ�!������ ��8��[^[��eա�2GD��՗Ӣ ���4�yR�ǶnO����q�az��|E	�
Ω���=td~rs�:�����	����F��E��2Q�ˤ>]�0�M�T�o%���[�#m�18�1ef��Q��L;����C0�yg�\"�Z*��1��E�(���ctl��0&񷛲Y�>���m��/�|��M4�30�09A`�:�h���9埈�ǆR��q��Y�Z�8��E��M�ol%`X�Ȍ@+�	�u�\%���h3!Ѷx��gQ�%�TY�zXT����������1(>w�UT�]�8[tG3�'��]Aܞ���fC�x�h����Y.*3w�؞�|5+3S�^	��p͹}&fl�~���Y�����,��WQ�@~8E��OO�{I�ZM�hk�'>����O��0����z_�_D�FF�tK�l��fgF	�Ư�&X��dli�ke;�diYOrՁ˴���zմ��aQW{��-�\j7P�钮T��G���Q�w��K��j��d}WS�FrgE�'�+�rE7M����4bչQ�&Fu�K�O�e������>�ij|) ��WR����K��Y�Fg%�!���Z�]�)��Id�|nC<��}����(3h����	���˪�Ԩ�T���
�%�\T�\	%��1��n�����ec�P�@3WE�T@]�+FD�i&T'M�F�V�d�t�'�4`uWku�Sµ�\���=�L���"=ܗhm�2�lmG����k�^&+��5���/U흯C�$�lٮ�Uq��>5¥G���t�S��39�G����$\�.Kplk�h�#�v����e;�(e+B7L�8�77c�o��5��ڳ,���;�c���t��Qo S�����2�m.�5��7OB��Z����$��f�G&a�<��]�YN,�È.ם��ޑ]��d-i!�9�c�ua��5���4�|��/�jg5l�hU�� ��w��)��·�|��C�u;�-35��,>�U�R��D\S�n����憫^�{�ķ�緗Aվ5���U�{�=�(��,1�q��bstJ�#���j�a8�q��L��ad�\�9>lN����f�����f�ۼB�/�wm����b��S41������\�7]Q�%eݬ1m�9�ki�\ƍhԫR�CE�I�'�#�:$Gu�]]!\Mwn�cH[�|:��o ����gc�F�̨8�u�J�q��u�`x�#oV�u<�V����&�熟gc��v��ꆖ1�-�.Y�:��\J��j�EE,Q��m�\��Vp�]�V�]`:ӛfs�B���h04ݣ;v���0�tn��k]���w$���@v��%��}g �Z�u�*�U��4)�5���ڦx���v��h�#0�8���m4ڭ���=�<�S̻������Q�p��)�����>�It���$k��=���{�X�޽�ά����]�Y�"�Ɨ!��s��N.�w[W����ɟ��ZFmL��s�&��B���	���!��XZ���*�|],;�E�5�����k0'\��}n���� yhv��,�r�{��/7U�dh�ɂ�r����3^cu9��bl�27z�n��2�n��ëh��ލsA��_%6k��ڮ2�Y��^Iɶ���ۼ1�Ev�]�V���S�K�+)��@�6o��lY��V"�<nb��1�ە��m�?������?yd�������8GlQk���ui5�[�N[�P�ɥ��{�rr����V��]mRG�޷���w2�Ks)�I�Z�D���ѝg�Tv��,����Mͽ\NgV%�$��88pV��ɜ��3f�e0X;��n/]�W�M�+(�椚�^����CC��kYͭ��3����>�v�wjx�#|nR��>��9��A�~J릒���7��>ɲ������)� ���Z%֥bXsVf���s못6�Z(���8��zX)G+�ʳ ��H�U2Nb,�)^z���j��3��9\�Kru�I�3��e�А��4̶���T���<��.\�Q��fL��TB���U$�+C��[T'\��{�&��Fa��,�G)
�+:],U��2KEE*�SZ�ZW*5�jEi�*Qr*�]) +$"�b*dX�,2P�K�Brʌ�
F"�JRQ1iQdZg5Af"(�"r$R�&aU\��4ЄCB-���F��Ijq9]ML:��lKB#��ReE�AF�bQ�Ie��8�s�GR0�(Vi\�D*2�)e��)��R���+(�$9ZY�4�D��t+B�u�"���Ir�0[y8=V�#��خh��,V�\�ᚚ�d��o�_XT��k@���R�oA�i^��3�pێN��݃y��ʟ�r�W�,`<''e81`��|�͝3�6+k�N�B�1�An��GC�2۬�z�h��Q���}���}j~I��PU�G^�\��H>W�=�_kw�giWU�lٔ�sU[ϯ��cۖ�Ѷ�YƮ���O�}�����Gx�;V7\�ݙV5-�h�a�� ���4uO>nwQ��͜����+�|�G<`�[�KoU�g�t����ww���<��Vu3�3���r��Bƞ�~6�^\���A �D�p[���o�5:ː��Z&�q~���Nÿud×9�/���m�e?��'��.�>��m>q<Ԫbp���]W�f:@�ɞ�̱�� �(&j�.��U[���i����/� /�\5�Zٹ�|���E�˪�0|�P�t]��n�\}𶪂�R��ҍ��zl槃��X�V�}0��l&��֕C�7T�
ߣ8U��! �m�d��8���L୊��[�po�!5{W;j�j�sl�Wn�B����}��zfxK���ɡߕ3<;�u������6���1"��o��B4���7�Ω���A�>��I���Z:Q�a❸�Z��_*ԺS�gX��Ǐ�"H�b�4�M�r��F�
[�KխxC�u��7f�O�S%��`�`�g8���AV�b`��r�;LM��l�W%��:��W�Y#��cW��q�#D�輌��7���7wQr��8��~n�������M�}M4�'�T���þ�Tw[�i�S{�'6���P���҂�sd?<�ިzK����9�zЦ�u���<��h���%�Us��=�#����a<�n�H��Md���P�I��VT���}hD�M���Q���i�]Y'�
�P���j�yX>�!cҜ{��h��`�ɩeY�U�
�~�M'��w�21�ƥy�V�<�j_)���UoNW�.yվƿA�{ƘX
�xdL2�r��VU��oVv���Cs%�;�:#�4��_k��[�|����C�g��P/ᯬң �O|@v���W��7��ߧ�������om�q�z���g^TؿwF��m�,.^0��Pʦ`�����4P��էk��!�3d�5��,ѽ����egE�E�i���9mI�q�-X����^Fs[\r�F'���a
X�NL�S��6O;��R��<"rSOU�>߾���Y����B��KhA�Oq>o]�< �^�D8�n�F�L�
�Ds��.��a�JX���~/2�פ[l��anX�9���(f��x�Z/�<��8�s���OM�K9N���eb�36���זtg|;.s_�Lb\VZ�4[
�[��qF�l�l�"�n����l8���{�sU�¥u���h
b�b����2r@������T��z���iq]��.q�i����)�
�
�s�"{�k>��+����������,:�Э���f�F#�T6��7k���-��FC�����9(j��z*(Xg�����6�<n��_��9����߹oR#8��i�4e.���~}Ɏi�ܪ�.�����w��9��{��y{�7��s��i�Ϳ:�d�ӯ���t
��h�^�M+�G���9�My[/�����{��X����!V{f������Eи���k����}m3��D�A�S
3�i��LP����l��Z2m�	�xe$�t
o%�\u��'�v��RX�o�L��ݼl�On>��|��y�<���l�������L�	�s�)�����ͻm�E�[`��]�7gVW+5�K������=��6>F�u��ꅍ����O�=�W�ΩH�zWVi,�͜զ�y���U@j����;�3��=R�[��差DU�Y�u��|���[�W$fUWn��^�P�%�f�90���C�G_Ep���q֑����h����/��C^�ܦb�a��mv�Lr��,9>�]�%�֚:e.��\��Q��M^���~8.K��\P9K�L-��/n�/ r/�p�����	��vV�r�[���m� 8���m�8��m�r�DS��n�u�R:��#p��,a���(�d��OF8�l�~y��OPeV8&;:�K��������0P��4ڌ��#yf��9�J��X	��{v�Z�J`�I����3:�ߠ�|�m�s�ă��l�j�3"u�wH�R���$.������B�����M!3��9�b�xbzOagd��6��TȤ�
��yC�Rז�v��%; ������)�|��/t���T:1X'��Y�}7No:�m�2j9����M�J�rz��S�S.��xuy|����s�%�>�`�}�&��y��d�ur�59���n�6��Sv�8C+}Ʉ)�� :�~��t����۩}
��7�xȀ1�橧(W�.�{�'�Cm�dp�n�/)uu7[�L!'p¡�ʄWv4
���1��U�0TwX���ip�9Wj��K�W-~�1t��+��)�u�[�;
߾ך�?v�����ɘ1Mj���D0Y,�p�r�]C$g�����uus:�h��Q�-��lJ����k��)�������� u{U)Iw��<�~��4*�u5Z��Ma�*�d���j��N�Ze��,��aӿ31N'=6��ڈ� �k�oXG�y�R]�O��ru$7-�
�[��#ʉ-�)��5�s'-@��κ7�Lݣ����1�����e��t;t��u��� 9����|�����{����po��(����w��|%�L�H�h3!ѿ<K�!�%�Ҡ��kW<�Vqxۈ ��}j�4�T�=Է-����H���#�O��]m?|�w��d�D}�&)�ic�s�Tm�U��'o9?J��4��>�6��L�>�R�]�����SN
��d��+������HU5;��t�2������e�;9�`Y���"a=��Z0�?M}4���(�.�;}����V"C��\������C�C-���
���	�N�z�3�-��w������&~��b(=nv����������m�C�������ngEH<
f����e�%�;"5�d�:��gH���B��;�9�O���}}s��[#Fڙm��ɋ��^��:���֨l���e��1���\�������p�GT���u��d�J2W�8�L���B��l7UP��q�k��+ls4�:Y�k3��z�6T��Y���l��d��� (�۳���Ig���Fy�����z��"��ܬ����M<��%p��O�%֎hY%�6g�FX���~����yZ������G%6�u:	U�/O<+�^�h�2���i:�xlqS��6]��/+v����+�'��[���˰��SO���P�t'y��J�ٱ[\��7��&%��6��u�yr.�i
��D���I[�"�;���)F7d�c�V~���O�F���n�H��4�s�-� �����lc/�d:�=�J��~�vX�Xɢ�p��	��6�{Z�מ`�G�UC9Ѯ	f�.U�*TpM*ԩ�L)�����h+/���j���t���M ��я)�49
��3��ygz��9R�@����J�ޝ$�*z잢C[tf�h����a��U\%�L�!Ƀ�#A��>҇X��=�`��)�˙�n}�uN�V�g�޼��%˕hp������Y���i���h3!Ѡp��W8��*}�I;����L<�͸��l��}�z��.�[p�w޿!M�뫩��P5�R{�Ԗ\Ͷn�8�4lH�Z���Y�~��u�.��~�4o���wus��ؼ>�/��[ ���V����}�)���o�)�E8��b��c,cHX:F:���Rʳz�@�GI��gǥy���v���wP:��ot��y���Uo[J�������e��KSOȭoo[i[���m!V�9;�Qp7bM;���3���_k��[�� ���d9���P3�`��U<p��g4R۝l�Bo>5E�r���'v�����r=��g���,f��.NMֶ�����s�(C|+��Y��Q���]zz��s1��4��s%��q�ȸ����ê�����gXdV�S���S6W���: ��Z��c]ے��u{"�%#�����5��OMV[bz���D�Ӟޫ/~ͷ�>�Bdϓ���*1O�:����(�U~���)��89	��뇘��l�¾���o�c��Y2DeV�8��2*�q��#�xĶ`q�ݓ�$SOC���w8���RxEʞC�zz���͐y���-����u�O�{j_��P
�DH��U�D:g(nDs�lR�qD!	;WY��u�W�#�-�C�	����m����1���Q�̲�LA0�3�P�B��FK���]zw*���G*z�����n�7�Kv�8u��c�h�p�Awk�y�%�ƺ�NF־�^qܾ�����9�����Ϗ~�H���7a���.���o�1­4;�L ��ڋ7˫��d�Z&r4��OY�ࠡ�	�Sn���/j3���7t�����U*i�] ކ��]�Y%�\�%�C�D��^�X5���9y�Ƌ�(�����7wN��u�n��h���;/��=�31���!�b�-7�\&�ᔓ��+̗>�%2�{���t��媅�w�s�m���^j#�V^3��1[�7|;\�Pyq�#�Y�Q��3�[]�BE�6�4n��i�� ���r�oɑ%�.�rZ��ĵC�)��I�����b�a]�X�p�'�u<[�7KWU�q�c��1Ʋ����;�r�8v �f�i��r���N;ϛ��(��ƃ2�`%�]l��4��)�,�u������,'2�Vfji��ܣP;����/a�E?@ƃR8}�yhQ�1�t�̦��ݯ�]u�.�n�r�͓R��L�j)��$8�S}�/��z�G�Z��U����<� ���n$w�A~iP�m��|�d�?==�ׇ��"�O�n�i�^=yV��f gFy����ڭ26�	%�E0D2����Tc��C�5��t�������eO�.Y[��ugTK9���֨��U�|=.��N�'�Q���믭�zP��Z� UY� b5�4O�/����N�>_;��a)�~(/�5�M�s�6�)��m�9��A�U93��!3��3�lRPs��E����b�f�S���j�Kl�% �W�W�3���^�b8�B�F&��Sw�J۽�*�_5���3!��t�:��O��"�B�<:���2� ���j�R��^�����b7W���1���C�X����U�7��6�ܩ�m��!��>���Ѐj�:�
�����Y���-nWb��G�&Q���6賴v.*���h�3Y�,<��E>�R �G��t�w==�5/+Tͥ�+��t�޽L�DWQ9�܆�	��w�Q
�;���N�k����t��*I%Uʽ1om�nMf�Y��]%��ɺ�)C������`��CM1	ʘ�(k*]X�ܞ9��d�������,4��I�H;�MAQ#0;:�ԡ������n�\=Uڮ|�dF2Q�]!��U�n��p�w4�"���q]�j�^R��jܨ�C��vиF�.�S^\��3�H���Ϻƅɋ��S�u`�tw�6q�wL>o���M2��	�T�Q`;�u��>�+c�m�1�	��8�~�T	N��-ɽ'>��V���s����.x�u�\%�Dt�f�2x��u�\3v;gl��V��VV�X'��"Y�`9�;U������Ͻ~E����a�}��n�sd}���DU��	&�}��k�c�N��4������MT=zʗ�n��}��!M8+y�Y��[�/p9	�~�:b
��ې�[<mU;9��vd'�95)螚�xz_�S_M?Fº�u�&�-���O@�k�"���MU���k�"�|�e�s�*B�0S`?Z��<��{�H�y>�.�3$�29ܡٳ)�߱U��.��m�C�]Qi�VUrb���Xׁ�7��?z�e$�?Z� a�o��֮��4T�|t'*�2����-h���4����Tf��P�#��ٵ��Ҏ������ΚZ�g�cW�M2F����Ҿ��|M�bu( qj��v�.��Fސ90L�r����RUr�	���޽�&���΅Ξ�	Np�wL����>���x֌���0��dc������1�*��4���yh[6p����\�c�{��Pg���p�������8�����B�$}�8��Q����=�� Ve��o�*$�!�:���*gx8�[E�T��Y=6�]E�ڹmIi�2�3��pc�Cf�������%�)/M1�Aܭ�L9sY�Nq\$�v�~7=I��W�1P��O%�h}����o�kP� ��1g{0��By����꼵^�GܶBD�R2)�ҭ�^��~����v�Ges���2�Z�w*)�xg�,%��!^�.�P]wi� ]�u��H��ɳ���r�@��{:��%�B��g�>�HC��?���R��5�܄���V�iwq�ž�J�CZ�����t
��a�3<%�DB�C�*xw1�4��X��^���'��~�r��r��f'��{QƇ�f��mg讖�e1<����%�tT�3�gE�G�;=� <��uH�q;�f�8el�>��}�}���y>x=/�lcco���6��61�����1������lcm������!��������6�����6����m���m��c�}��m�����ѱ��m��c���lcm������v1�������6�����6��1�����PVI��l���Av` �������6���ET%$���fP��V�m����*J�T*�*l6ڈlʥRA"����T����
�JHv��k"RF�)���Ml�Y�-���jc3A���*i"[�-5k�M��m����5�svdL�����;of��m��Z(��&�ls���m�o���#cV��jiVm���-��ڪ�&X�YZ�3DM�6��&�lش�V�ʫF��b�Mj��d b�R�Zm���Z��ff��1��ٟv�[�δ̑�[^�  .���]ZΆ�U\7����q��=�={��V�k�5��j::�d7x�y5E��xs-t��3�f�m�^�6uU�J�����j�UkBk)�fL�|  s��*��u^����w5���u��h��G�_n=h�:P\���4}�
>���(��E(�F��<z(ѣF�(��-�����R��}�|Q@Q�h������B�`����Z��m6ʴ̵X�0�ۇ�   o���j��}n���'�����+;f���֩Uoqǖ�#j�C�z��K�u�A5׫�׽�mW[�{��ښ�h��l�{l�km������zj�v�֭���#Tkj��cV6���  }�j�R�z�秬�k6ޮ{n�=m��۽�X�{j�9n1�w]v�M�{î�[۪���g����כ�S{��`s�p�{Sܽ�z����I��n�]45�m[�,��g*־   }�g��qû�Z^�t�Mt�j��z�m�]wz/y����h�[����Y�����<ࢻk:���m�m���ݽ�.�u���b��y�����.��k������QV�L�6�L�f�ݏ�  6�wo�m���wz���({f�{����m*��=��=5m����a�u�z��������wj�Lh���;�Y��׃Λv�m��\�	�t��<��7�n�����uV�ck���5��'�  �z�͙�f��ڷp���/S��w:ݛ��]zU�7uG�^�UW�*��q����ܹ麽��oj�m�x�=z��wm^������1:0ˢ������[%a���f�kUe(v� ���
޶Y�^���mZ�����w+�����^���u[�����n�쫮[���z�ۗ]{���ӹ����{�u��6���a�����Mnk=N�:ҽm���j��m2+Uj�Z�Gf�m]M�  u���u�uљ'v�Wgm�U���=Glk&�ǩ�CB��5��<��*WOy�u�M���z]��wngN�{M��DtkZ�sչGm�[����{W��J�ٲ�^-���m�gc۝/d+3
.�  �^���ӛ���w^\�յm����;�]��^�ۚz�oV�hku��o\�]�oz�5�vg#����Ǽ5l��l��ށ�]v���죾 j��M�JR   �{FR�� ���x��L� ���~%J�  ��h�JT @)@�*�@ ѓ�S�~������G�~���?��H�>w��)�G߼�|��߿�׺����ED�_
�(��QQ�ED��* �� (�������~{ў�?�����fc�W�RN��	�s`�B�r��4���ZN�:�cx.���d��90ᐴo+p���ֈV��dC~�\ˍ�s���8N$�VeܴWj�y�h����T@��?��)�B#��jb�Z�L'(R<�m��Aҕ�붎�7nʔ7�Dā����h�

9�]�۔ �5��&��U�
H�E����kt�
��b�!RVbwJ�Kͽ�v���DR�T�c/)����׿3��֛s&���!n"���v���Ҩ1�M<h�k,[�e��Y-Wb�f�D���[A��u/F*z�LnJW,�凎��r醦���e���Maǀ�hM�X��Ф�[h��5��{l3c/+Iʶv�^ֱj�2�S�c�t�uctQl��>�O-�M˺�G
٤�*ʻ0b3Fk׭�]5"�Y�'���V���j��ǯo�K26��U��a	H�{�V��l�6nV�wS!���zq��&���E6D�vL�l�t�l�GC��z�ˣ�#z�)�t�pn]�CL.��-�@�g��qb�n���bWLc��I���]m��( S��W[�n�d���Cc�EkvŁjt͈�	��(��`�Q)(�ү�/7Tӵ�`�P�
.�҈Q��2�� ���ȴ��&��o06R:�-p�AĮLR%�2�� bi���YN��B���h�x�ֆ�,٥p�i,�F�,��l�F�ԺY�E\�,��|�J"��ҙ�b���D&�Ƞ3.Sd��i��@�oJ97��ѭۈ�w�8s#�3 T�)��T2;	L�	�E_�x�/31�
���6�n�v0��H�xj:�1��W�������i�d��S+aEa���9�H�r�tyD[KM�(@ �[�p:�n�I�5�xln�2��Չ�Ј:���ˉ��i�e�o�R�n�	�L���DdR��-�* �U�q�mB͊X�cP|n��)�2�*T2��x@HnZ�����۫ݳ5�@�0X�oY�-�	Xq���եY�[�U��x�[mn!*���IͣwIYt��R��0��чTn`8bՈ�=��t�b�K��ȼ�C��hR����)�m�ՙ
W�9��nB�b��Hҷ�o3*Ց
F��з�o#7�8�&��G^3�|���]s��C�u��F�
ƽ2�up�ox�u���;��%#�j���8/Q/^m�� ����Yz�Gv�tbjf��6ճ���롣%�ʉ��[~<3�k}5�x_�?'�d	&�N�N��bV�n�;�B3oY�&T�eؐ�Vkb��(��y1h��B���,R76��kV��VBͱ3�C�,*��c���3sRƎT6�l�,ږ0�@�*݆�����2�Fm�k�$��#vؑ5�JcÄ��4M���6��@�bW��L�� F��Y*P[KF�l,�����ń$��5n�n�]���J�U�hP��1(wfu^%�\c˘茖U]2��@�.�J4�'�������y��6�Ǔ(P�bMW0���򮰀>����^��
�m�	��ҫc��y���Q��H�S�eC��A���ƳZ��7.���in�݄�V	7pT3f�K��9��q)�T���F��%D5���X�t�f�m�Kki3%��7hU����a
�7j�`1M�h*{�)�M���ŠX����nP���ˋK����N���5{j��嬓
�F΋��D�7pH��7�d�M�waL�nH��!U�X����V��.n�@h�h����
�Tڍij���;	*��嬵l`BԴډ�7d��Ŧ*�Xpf�@EˬW��Oo F8H�Dv�kx,�J�Yw�%�.��Mm�-���t�$ʹ�,S�#�uĀ�pD���tK_e�խ��l��Y%�Yv�f�
�2�b�ԗ`�,��J�,�Z--��XE6�R��%{�U�9���S��Kfӽ�:��*��-��-m���X{X"�jZ���X)[�
�q��7op�l��/#h5[e�Zݦ�Rw�l�I �E����2��w
ǡ�YStm3�)�6(�)	m�Na/qd5���Ŭ�X�0�b7*1���k`�����pܢָ���Yx�5 Fǻ���4$Ĳ=1�vm���ME�f�qp�V�]��ڗA]k�
�v�hVՓP��X˺NQ^�[�h�J�E<rK�
�f�ք�Q�����lF�i�S-��b�N^װ��܂JD��^����4�욕��ʛ���vQǴnE���n�{�+P��'Qh��pЈ\`^�B^�� 2��&���;c!)`�iQ)h�D����dX@e�n%nԣ��(�Z����7jooJM֚ �"�D���A��l�i��Am�XQ]m����gt�����o尷Ww�6��R4���֗2�7M𗘦�)���k.�5�"d+��oɍsPj��n�n!H�Bi�W�J�h�W�7TMm,$�l!�M[���!�y�Ǹ���#&;b��ac�q��0��F!��� �V���5��(�N���:�Z�u�r<�bZ^�7m�fU�se��u^Xb��+C�n`͔�nV�XQQ冰"������ �qI+hP�1}��zNKͰv!z�@�pn&u��,�=��=��!��X� aD��#D�ԞF>SE��d��q�g��?d��ς�sb�$�Ď�{�5�eJ��D�E���n��h�/Fd�[y�2 *B0�e��֔��r̬�zpS4q�Uan�R�k6��[���J�-�ߊ��n�̩h��t+�����Y6��l�Q�E'xL ��-�n���7M�6L��M�W�,7ڙX�{��6��M��[�r��q�K�ֵ�B�Ṷ��;m��Qyt�A�u�Tw�t���NZ�� R)�om�R��t>��� ;����q7��enG�Qxc!7�8{��3ۚ�̔�R��-@��"^"�ҶmB��W���	*XT.�U29%=����VژV�6���)=JZr$�0ەk6,�1�Wa��ٔ]��=�
9�S6��V]:�f�6�@�c#NDgn.�8.iN����~J5��J��A�;H�����M���ݒ'{EV+J�����ՙ"1:�u�j+xUݖ`Z��F�W�㛿-�bͬpU���`�V���*yL7,�)�[�z[wd"7s�)ěE�B��h�bW��e8#p˹�O��A5��W��M��ƚ�e�f;�"-V9�Wj��cj֠��n�ٵ�h�Pm��I&�c�sB�rZ.�R;�P�V�d�۩3��0~�����BPޚZ�_|��6��]�,����)괆�`n�n��֩YN�W��fEݥR�9�
[@���
*ܨ��mЀ�.��haoui4/,�2���3	�6�'�QĕCU�.�̼������ވDK5�&��ǆ�A�Sr�-�T�i���!����YǺ�QQ$��v�r�kr�e�su8��p�ǰ�.ĞffXf�r�j80D�Y�l%�A��
'e�;�]a1j(`�9E�+d�1]�u�dh���2X����x5���WY�X�A�u��G����"����j�m�v���A�׀�1�p
y��dt�E$:po�Pnb�`۬d��[���[!�[�2�m���ʣP�2

��C�2d�b��s,lr��$4�;��x0�N��qlW3i�M�cr��
ځŜK%��f�Fi�mYD"�x��hM��R1��Oh���ԩ�e�5IL��X�[ӿa�K6�h;*�]hzuZ%���ON����dc�Р)�̒���4�77b �t3.��D^�Î4�Uy�ʊ�
��mh͉��cD�/��*b��]��k鵬^�$�X���X[�V���I"�P�aq�ɋ�%3������B���+q��hfYt�c9���L��J���r��/n���b�"�C��7��Kk�-���%c"���7(,KX��V�j*0v)�[W� {���ȫ�g4�4f�1�3@Ӟ7�ֹ���������#��3� #�ګ8��%W�2B�b��:�نPe����BK�<iٿ*'�t�ݳeҳ�nj��[�Z�l�x�'t�J���ةG+r�N�����D4ͫD��e	%E�S�� �Q����l��n�WR��/)��oB-.�W�qұi3�f���	*�3n@9����k1f��(^��xD�MW�:�"�
��������h7��0[d'��bB�PM���^n���6$�#u�b8��ڂ0��6�w�Z	�ɩ�3Sdܼ�ilL5ct���j{�yC��/)n`��ڲ*S���U.ȗ��+e.�c����aT-���S&�]�V����ǧ&�r�(!��^(�CjS[�����I�I.�}!S�*ś��X���PS�Zu]h�cT���'��E(C�YKd	#�-+�(M�9��L��ʺ�WӘ��sB,kCO�X��
�Cl�4UZs2�N��̫�7`�	���ciӢz{g"nbP-p)X�*�9h+�1��2�op����Or|��h^���-T���V�v�� ?(�
7Y��ץ�e,�L�XSv�Zy�)�*��v.,�rFݤ'f
mMՌ=IU��Yk,2-��	TU����D�Xmc�t���%�.XE�n�պ%*�V�[�m�[B���zͧn�nl�x)���j�cZvh+� �"v��g�a;�7)���V@�(��[����ۭ7�e���;I���V��O^��Mi���j�(��-��U��T��cUl�h�v�{���i�B��a��UH�Xi�T�M*��r�'jXY�,��P�D��TQ��CD��Sk.�VȆ����cL��n]���!��P�c6����{�f��V���v��E@29�DrYS4�V5�'hh��>7N�� rӒ,��0�j�Jw,V��wH%6�OJ�1�Dq,˦{�x��٭��0��*�7ܣ�<-+����oL�{EAP��kM�Ҝ39b���j���IV�sMVn���d[4B��%�
+t&޽8pddoed�G7S�>otD4ZmӠ���=7�5OC��څhu��\�R5k6@Y7X(�"�l^�a���Q�;9��EN�ij�	�h��)�Sbw&�d�4�Z���pV�a�@���(�u�ڧV貝�nہ�ᗰm*Y���-2��%���J/ke���X0���ˬr�8.[�!T4Z9kL+�a[ubb�Y���93j3yf;���"�`�VދnҔ�<�uy���$����l�[hLY)M��GWF��/�Sb�H����x--ҨԤ��mG�ح'K5p�ج7�����W`��jۡEZ�PVӥ�O�X�%3c�+&S�$j7�c�Gbdجɨ�6�{%�*�(<��
T�q�:�e\I\�yvI��&@�UÂ�r�fZF�b�hi��:q�RGt��t�
���(���m�I�r��6����vӂ�+'݅w�ڲ��헖5���0kW�ڗ�2�M��ݭ:��y���s�lƳ�Nc�}�07���֤קD-���h��q������ ��f��j�d���6+N���H �0�ݍ-V��$�T�׮�	T�j���r�1[�Z��6�;����͘��j�� �ʏX��
�A�tdQ573��֜Ąn4��v�
���a"�f�6��О'o-q�Җ�Acǉ� �i��n>7�����n˙�T�d�t��^��=��hR�/`�P+v��*جTo�[n�����b�@J�!@��]ۄ�ą��"���� �M^]��Y6ށ7	���6���*݈�>X�3*��"��:�y(5h���'d13pZ�e��W��ȥ�U��谅��a�iq��v��`���*:2�sk3��Z�M�w"ӄK�f-j0�إ���@m���aT�o1��಻7ar�h��viJa��dE�J;Y�m=V�)�5x�u]�vZ�]lT��R혮��$���<;��Q��X)۴�R�Q�r��A�^�B"��Qަt^��iL;{m�x��t���T�Z��.�����ra��Hf��޼T]7q���"hɺ�B��q��hd��ct���d�ظՄ�1�x�Z.�b+��p�ܩ���&���j��j�l�R���d^}xp8u�bF%�[�nVĒ�b��;����u�V�קd��3@����G&����5b%��Ul�m0.�SK�Q��ܬ2��� �f��â�J-�by��ɛw�e�z��T.�Y)6�a��B�� "��	B�%!y����nj�Oy�����5v���(��Ǡc�E�A4�rbtnS.�]�ͥ�2kpd�E�E�i7f6�CZ$Q�����,f�Gyn^
� m�v��̙�x��x|7;��!l8�:�r�WJmfn�Ah��`#�\�X� �B����㼓de��X�b4,5b������O��0�,��1(/���Q�ax����[��m��c�C�� D��{,����M'�!P�62�c�I�l��n��"�c���5jAVm̶5����)��Җ�x(�;��ڐQ�y���eZ��aB��֡/0H���̘*]��Q������-J7�6�^jm-$yY���5�m/��v[��8$�"�����fGsĶ�$KԆ�K����9WM��ml��ښ�8�s�iXW"�<�<@=�H�5�s����u��������~u����\8���wK��0L�&ސwv�ZU�a��K6�����1˰�U�x�2k�`���C
2;�d�qe^��� ��ǎ�n�����[X��6���3��ۏ����y�0���];oa���6D�� upG��ug���J��=^^��+Ǜg�]�H85��e�����Z5�Q���Oiwy:t�p^�FKaX������=�l0ć�S����8�	w����t�|�>/�� �T����<�.v#<����S`Z�Ce!חo����E!AVe�3xBj��b��O�[�/V���E���gP���Jf�>z�ܢk{�1�v0�S� ���$���rC���<���fK�t�[|�+�*X[|�F���d��EE4�Z����F�p�ص/%�9�{����� @V�+�����v�=X�Uއ���S�|�Cĥ���W�7J�������x�W���I�c�cj�Y�F�A��&�&v����gn�.Wgesc�ўH8�s�"kT��,�b�{��vW\�ʶA]]���)3���P4�n6����u�{VW}�����nX��%��3�=x.�G�^t!n*\ى�mK̻0��o����v՛̋P�����T��yb���:6U��|��{�)�0��gJ@;���BvHۊ��o �fĺ<.��\ޱ�t����y���6���8�A.��R�jR˽��В�g,��Z��>�4虗�h��X���0�W�������������gf;G1�mLj�-�Ѡ�r����<���e����K��爇��.�F���U�����Uce}�g�y�}�)�s�\�H�~WL�.����,�^��{�R �0�/���Αym�ԍ��!�8Y�.���}����R��7My���9��VVY�q>�{����e�y�
>�8>��$��\��f��,0b�e�~|rRg�3r�����/�f�s̗�t�L�PՈ,Yם2����.}��h}���M�E<1�ݎc`g���p��˻Վ���Y{�P����K����[h��X��]Rv����ʜl�d�Zd|�N������mE����SY)�fZ��
b����RtiWh(�+ڷ�rb)ldB���]�e��[!sz&5[��v��t�a*�i7�e�] I��]`nv8��Ԡ�ǠګG@�?^k��T���Û��W=�v���2 .<��%{5,�o<l�	�+ ���I�����!ѧ���m+C\&�t�nG�)����vM�۔���G�lF��bUt�l�N�Xn���Ղj�̡��ge�hْ�l]�.���fh���W���2�u�A���)����l�#0��Eل_h:E�z���N�/`����R�6<L*�d�Q���VjҒ�ę޻� Ӈܳ��)s@B�<�;��5Z*��e$��ͻ��}4������jɲy�����\vLam���{�c���<��`=����6���
��)����/l�R㋓13�)�.q�-�)ѣG)�W�H��#�ǒ���:��c�պmo:9}�:t�ֻ��ZsP���]ɚ҄�{ɶ�k8E>�d�xg*#�>Z�\wK��<�ћ����K|l���緖�4����\D
�f��k�4C�\`5���I${P��D:=|�q�O5��u}����*֑p,���u���K��9Mɑ�2���#w�mQ}ȱN��Ԩe�pVN:j�s�QV�.b��ֺ:X���IX�Rμ�{�Ҋ�|�;��5K�=�O�n	��0,�J�&����*�w7�<��l�M��R��rﻞ��*���W�.�����ir�b �<;�1��,`^��Y��KT@P�K��m�K�� Q�{�ij��c[��-�� ��b�=z�\{z��Y�����ڔVb�!=^���-�'�tZ��V�t\Mes='/�C�-U� �B���R[��'u�T<f�����[��N�K\/;���!K�l�Ax��C0IJ�#�\C�E�g�}���x1�ԫ�׸�G�l��!���`�̑[�@n��>'r�$�#^#a;��l��t(y����bI�U�=�=f^��+q;&r�)w3W���u�J�C�T'[o�K=8�� g{h#���xrZ�4u��>{�C���@���UU�sg6����+qUs�oc��qú�Jw�f�u�/�h�{�+����g�4��%R����wC����d�9�l�.�/.hIEрF]�Λ4�hO%�W�{x}��>�M�=EU��[i:�6<�8 u�IN�$)�{5?E+�D�۩������]%_�0�U���-��^Shd>/ol������l�� ���3�#�6mXT�b�/9.:u! ћoM�5`�Φo�����Q���}M�J��Y����^��;����X��6 ݢ�Ӳ�vwz����m:[��C�T���ľ�	uk@�}LX��i��"����斏de�y�q�Шnn<��^J!�U����-�ZJ�.�}}�l;�Ƣ��l��e���N��g�k�/g����y�{
�[
D��ى��VLU�U|��H��f�{�D��!Jn��gie���n��<R��G��
�zfIe-���+Z��E)P)�V#��:�2޷Pm>۵՞��!��.�X�Ή�mͩ��P�!���ӕ�RgHg
goq��i�dÌ�)v�唓ܹQPRP��e��$�ŀ�6_O�@�l��\�ʜ�� �q�F<�ՠ͙ͧe�q}jNi:����d�e�Ỷ+C��u��Z3�"t���CBYӪ�VI}W��7�/��J�P��Em�o���y�{���u-�%�҅�ҙ�K�B��-[J�vK82ͱF�]am�rNv�.�r��vT��wH�Z=�+��p�W���k{;՟�oS��q�Y�����y8�H{�]���$[[�:ۨn��T4S�u������_*[�9���D�����?�g\�T6Ս�Z�GCݰ����t���)��^�4l�WI���*�ͱMm�nwe�0,ĔvΦ����8�#��L�q4���Vd,J��#�1D��a�����ef�{������)�7
v�3��NA�ޓՉF�t�	M�o7���J���m>炲��@ݾjY��2j�9@>����o���x� ���+:l�5�HP<E�4�'Fљr2��U+�x6q�O�(�	�n�Yݞ>�Y.�t�Oo)-�0�6_T\Jv�ٮ����-ӵ{&2�֧�3q�_q��D�+*�s�{��]��-G;F�7H8h`I>g��TiLUvjq�e����*u�Z�S�r�*�ԭt,�;�Ť�~��,:��<`(+>�^u���=#�+L����<p�uzS��$���#܋luT;w9p�b����#�ed\3m�Euʛ�KO�/&9񫻁�U��{��^e@��bfm��F.�|m��0:GeK�Wv�;2�!9�۶��"T_��`��=} ��6G�:.(�BaS]G�.��3��`�����7�ᗩ�/xC�w,.����ˎ�4�+�� ��l�3��&���S�R�]t���b�B͛7)dfS�u^�շ�ֶ-�6{4�=��稴y�J��p���Myuo���r�f��u����a�y�vMZza��&��-H�zn�&�#~i�C�k����84����p���k6^.��CCaήCk�L�a�(�P���7)��w-�	⾧��3K�[y|�gZ��^|��U� N��ri�������D��g+qޱ��׶UΤ3���/��F�|����[Ў�S�m��_�C~��=�F���y]�'+ޠ:N�q�Y����i��*������Ql��؄+�<e'��vm��nh�cO�퓹'���������ѷ�C3<��]��N�&~ƹM�Ԗ/v���]�4=�\>Wv�mc��%ۣ�V��ƹ�\��-o�wh�\��-�T�9�I�]��bG��\������µf�Pȱ��@���r�'����:$�>/�t���>��te��������AsY�0��N$-�s���]/8_(�ʹ�3*�^�#m�D%���j�km���.�?�luH$�7�x*Ő�/e�v�1yA����Ș�'�jm����:�0��7��Wˋ�tIҏK�:����=y�K�Քi��\��1%���X�]�����3+�QHP���m��r������NXm���{�9�'d��}i�"FB�}�2�6�$6M~�A���Uy(POCW���R��LI>͠(+��L�´��J�| ��}x;9���~.��[}�.��V�aD�	YF��}2���� ��,�D��(�
ĕ�`0b�{��0�r���ײhʻz����r�c0�ƀST+s_Cӭ��ݵm�V�����z��&��N��������07
-�O:���V��Y���$M��:�g*����Ԟ�r�n�`qS�<B%��u��r�nt�b|y-��X���s��No-ٕ
�:[��Ai��6����o+���z�@-1BY�uGkH7���=��f��vʭ�w�t��2�=W�d�:�o��xT����NjE7�NI����;����יP �I�������0I�u�V��l=\��ܣV���;�7N
�l(�]�n3���z���U��4\��R�%L���.��yҦCv���/-4/y�xR�z��ͱ��% ��J����'Fѻ[��M'�sn΃�J��˽�A��$"�)��b�t�0�P���\��s���E��v����cթ��<�&�t��WT��f�H��)����}�ÞIzz���}Ϝ�󲙫���D��͗h�[�ݖ��{,D�.��pS�9�N�2�=z�_>8�z���K:�RǞ&�Y��ɚa�Ӣ.+�U�����Ugr��S(����aϠ��a���ڂ��֮�L�J��m��*�'��L�ޤ�H�X���uw��X�u5��B ->:��r69u;�-9KP4�,�ǶI:�-���{��L���"�Ƹ�F��ꈷ�-Sہ�����ŊŋA=��z�|_Fu;�7x&'7���gsq���e�CBJA&��7[�ݟT��Ǹu%�O;�zG��k6�.��r�<��N���3.�e�hK#''P0μ�奒�.��hPPc��	!��D��o�u�}���R>ۇ�����8�f�RM���r�̾щf��(V+�u��l-��c�! �ۧjB��.l:F�f9.��G�=�u���ճ�-�ĭ�/����Yz��7�:��	�t5CҲ�ӕ�g�����a4��f�h�iw>��<%&
!��$C�%���	����.^YYHU�L��թ����m\�ݡP�-!����ջv���U�D�9��f��lxW ћ��Ә�(��n�
�T���4���Xs1ˡ٘�]�&�8�[;jF�,�h���>]h5�Xzs쭠A�Ow/:�Q� T��Z��.6�8��7�b��^`��M��:�>�W���L�{@WC�HV�^�q1ϕ:�������Z_٤w-ya�X��*jJ��T �ʊ®U��RJȯ(X(�Q(�}2��
�"�����#�%h�ھ_[�{K��fm�V��Svp�Q���Qr��
�r&�̚YGugY��w9�����/vk3NG�ImY�[zl5���Ϋ�\8�Jޭ��#Zy�a~���0��|5�/J��r��x{:u�PX��%����ٱFh�C�E�YK�P�m���<{=NyNO]KE`\W%g�T���*�e�kUS8"��諆�O�C�1R�k+�X=QZ��e�<�,��a�J��뜗,�(�;���"�YD��6�����1e��<{^�-�;�)�f�lf%Ϻ;<-nS��qQ�,�hI����!����%�<�j�ŜRh�r�mËO<fY�V%�G2��|i�y��.Sh<��.��]��?zH�7.\�}sʞ~|V���`�Ub���M -4���	���ݶ�hn��`��Ϯ���Ã4�Xt4�6Yc��\5*K�3_,__::����{��~,�WְNG!�d>�ֳN>&���}|pj����"�c�Q�'������|h�*���⪊CO��n�`���Y��3㫗>۲�8SH�YhW�G&NP��O�F!%3i�ޔ�T����/��
�5S��V�O1��=�u2��m�ua����7��ڤt���_j�u^���i��9b�}��=�U��D��)XN�\�r�9KD:}�c�}}Ǧ��E���$z��.��F^:n��[ċ[qZ��7twmAj���겳��lٹr4��k�޶�5Ӛ�6���p��f�=l7WqS
��)� @*�����������[:��
c#����|Mp$n�w(9���;,��ݲ)Ӷu��aJ�]��[���L���l�qu�ֺ;����>�R@]si�_hi�I֚���ʞ�q2��-Ľ�c�f����ȡ��F�H��nk}��U�p���D��(�W>�;�Lc㱱�X�Ne��Y*oR�:�9�e3����O��_� 洉ՆL��3.�rg���O1��_�E8���f�^*n�-g*V>ĸ�[\wueJ׵�`�7򫊎%�jۥ��Θ&r��D��5�ND�J=��'.�md?D��ʏT��*�i>�2� �N���:��b]�~�ny��K!�S�Gԝ�W(�A��0�MY�Wpy�J�bj�'������k��~�u׿�~ֿ�@QO�ED��~��ï�v{��+���ˍ>��+���4�|n���*H6TbZ��X�%�#[��:��#���Ճn$�w�-ؽ��6�昉���x?j���z�9S;bf�|�P��s�����w�|�i-���s}/;�����FأX�-]����t#Q��0hU��Y�l���΂��"�p��)LL�Dd�iC]��d3&�T~����F!���Td���Y{�p��r�Da����B���ޚʰLY@���M
�-�7m�ً�"Ն�E�b��.�$��Q��:�����듙����X$렒�uE�>�累7�;#þQ��Sf���|D0�]�}OU�Pb�2��Z�Gn6U+��_b����M$N�O-Ǵ�sAhX�[K2*�ʅͷ����lq{%�x�)]����3�l��PwR�>�Q��!黬��v����Zx����4;�v�wՖ�}ҬٗE�	#��#᲻�RK���a��4�J��Z>8��I�e��A*�:}Z��\/��.��5I�b�����8H�Uyz��سH��]wu�b��87�@�fts����s\T���RW6%��{�L7Ĵ���yq�`W4�q�r�_=�)6[Lm��t;IE�n���)�<0u�E�q��LS֬�z�5݉A�82��%6��qe_&*����f���v�������'P`!�<�!�֎�3�������]����.�m��-�����w�!Ě�
؃��V�a���D��l��"]vk1�w�C�+ɡ��x;h��
С��wibYB��Nzz.Сں��P4��۴���μ5��J���R���Vr4�{Tە_�k�wO�ӭ���6>���n�ʘ:�WR���qI�6�F6HbY�u��*���7�(�|�?c�i|C=De��+V�����߯����#��>��o���r�����$$!��
y�K�ZO.޺v��n�L�����o��|`l�j���b���@|�8��u������X�)�E��xx�ҽg����{.n�`0娰���-��K���=sf�8.{���\���Q�)��GHao3q�S57��b�<�������x��>r�N��J��6�iJL��у�.�K[�ɏ����.X]�eJ�:�EB���R��[��k���.̯q�=ΞG]{�\6-G� R�4���L�Kx�\�Q��-��;3YNw|�+z\�^��q�q�j%n���4�x;: zÒ q��*�b�S2�è��}7I*����`m���K�LXD������=��ۦ��;z-^��F��ѝ�]�<� ����i��R�Ĺ���F	k�0aW����	�e6)>���E/�A��5I����bQC�*���o�c�3֓����&�	��S�����0_����:ZX	��W4��/�GO7��%��o��KB[�Y��Z�&��^d�4��T+,r:�:��VN椀yf�<��r���*��6VN9�*�)�!MVʿ�ҝ[�6T8��PK�m[�a�8f�W�t��+(o�n�R�h�1�8|$�ߕ�m=u�2�nC��XT�e]f�fc�V�-��n��>�gpYI�/V�+
�����LĮ[�3s���L�9NL!6C2���;�	s#�,��6�ߺ�9�}XdN���-�͚w	/�ޘ��rIWImwf���1�C��ȃѕ����{AH�v��W;9VWB�Pn��&� 6�d�c("]�Ց]�rV�����"��CZ3s��mƍL�U�h�������b+,�}�S >�qr�n{C=_�C'W���F.ÓgQ�S�N�v;m�>�������@��.gf[�?(��J�ԭj��V5����d+�Y���7��p�p�{(��O>Q���u<�����G��.��YJ���Ru]c� {%ԛi��:�`��K����t�iTկ�$�f���1���&�s�D��h2��`x�\�*���OU<3*�㽍\,ܠ�l��y�� ��e�f�-�^�K@����:tq��ǀ�8&*dQOҬ��G�4�����;���7���ը�d���xz���f���Dئf�dyC���O��U��)-6+�Кq2��}�49�)��i�E�J��c�=t��c��{XQ�wJ�RH�wjа��g��C��{K(,kxZv�蟍��뒥��^�����7�!��p�[hJ$W
�Ⱦ���{@cZ�R�KӅ[֧&�֘W�{��z?d��Q@(�`K�Y�ch���}�����Ψa���zd]��沝�|ZH��Y|㼬�ef��<�*�C�<#�Q��H!��#��"�杮&��wLp��$�`����M�K�㵰�τ׊�@ �|�흓ݎ�/Z���j����9]`�u��m���3�m��]�t��6�$NK4�b����Q'x���
�,Z���sn�B��֭*���vp�/f��pa4�dc��n,ɧ�'�nv��q�e�򛙙�4e�i�i�,�C�Ќ��.ӽ J�^�^Q�W�{\��-B��@.M�,�����O,��]��FȨ���6�3o�**�7�[IH-��;��Q�`v��|���EMW|s��<��T/�M���4�J���"�4yzG�L�֬7#���v��#PЭ�=���ڔ����ast��IB�4�D�3����[����P�8׏zm^�ҭ�7%;�N���:���<�2��G��W����x���\���x�憪��K-�Q�"ӛ&���!._D ���3���"�1�E���S׹A�Y&���:�y���ZL8��)9��T��?7����:��V.����ܕ��t\����|V�⼢�$�F�>߻L-f%h�ĄB�Et����>63M����ͽ˽�!��>Y��*K��,N���HTCu��-�,���e�t6�S���o@��(�e֑��l�ߟb�$璎���+7�"�jv�����Wt���7�u=$w\�Z��!?r�|��6���,�鴎�����(f�F (q�b�!=V.��Z�s%`�˕�}D�z��t�u��#)�(�J:��.�=��%Ջ����_`smS��5uٖEMK����y{�w�Yd�x`��](lU� �%� DQ+��%�a���d[!�<�c�8Kw�9�n���d����4�G�:����sG2(��sN�Y8kL�˾��u��D�Q�n�Gk�M���&�6	z�*���Y�l:W�U�ꀖ��	����������}���R�-�tƺvй�lӑ�U+�6-�g��h��ɷY����x����Y�Fɵ���l�z�@���9�������5�����`-�.�@}�6H��^Y��]��擣-l<ʀ�ߍ��>��2�� �0��O���(_2)�31�-�!ov���Җ�3� ��o]�QH�Ԕ�댽��/`t-պ�&x��A�K;�"
�Ӊ�/��.9�rp.���[{v�W�
V�dm��0!)��Ō��uL��X���]ˁ��*a\�����ܭ��,��o�f��b[H�:ہWR=��ç{���7\�����Bʝ&)��M힏���J��g�^-Y��;rV�(e��A^TS�v|#��GQtqJ�����N���ݤ���5�Y�2�\��a8X�Dr��)�]�f�̣ͫs��OM-���4�C�\w7v)��rT1�;��Ed��a7G1S���M��uJ�cM�#�f��7� �����Op���s��6�������vNӥ���NP�5�v�|^P��X��Tһ;]�2e)ﯘ-�j"1���u*?�T]K1�\�#��n��"9F���<�4,��%�`�ٛZ�;�����ɤ`�wy`k2�h������0����Y��N�(ҩ�2%��n�h����[�!77X<�緄B�m �XT�ru�o�4a�=vU>�pK:��]|��Or	�O���?'c�h՝y�RǞ$m�D�U���S�+T������,j�Q����]�j�(a�;�m#�5�x�o�O'm���r�.;Wu�RT�A��bNV��X�Ɩ���M<+],ʴE�؛V��5�%�����5�[�Ō�2�����'Y�^	��ݙ��l��kӉIֲK��t>�\�P��#{*]a�>������������\e��r�lԝ]%p��#��l1�k��c�wD�5���k�*KD{{�֡\\igjB�p���8x�������5��{�b�޷q9a[�T��֦����ݳPђ/�"�%�^���N{�]cIU�$�-D��^iɻ9� ��\� ���� �v�ا��s!��;b�����ܹ��o�1ᴤ����HtH��O(��F�i��V��XGC�x�$���]yjԱ»�%O��i*�ZV�Q͍�=�e�ȑw�;fƐ��ض�b����H-Րզ�F�n1��;�/s��ݔ�l����[��e�q�)3�<,Zu�`�p�:e��8����6h�8h�(*�v(�&���Y49�S�E��O�Ywi�[B��+�Qd��"�5·PY�h�W����94u5c�2t�{�Sg��0�i��/��d��}�	�G��Q|�:4�d�7��zs9|�Ȇ�/$��JX�h���{�˝��Iw"��Ę��d�u��y°u�T�Gp����k�[w���R�5�(N��p�|3�n�}�79̡n����g.�b,�e�T�/b�mI�����th(C�V �{s%;1ā�hc���
l	X��v��������5�.���+:G�lj���])���qL#�Yb�oc)oL�0���)c3o����Е�����A�ʂÃoi:�D+��V7���"��։�7�S���;�k�M�YC������h��0mk4!���O�\ju��ǂ{\��qgr�n�HnC�Λq(A���U_�2c�	��+қ�o�#�����m���8���CF�Y� {���I�}&<е0̮Av���#���������\f��2�%ti��EH�"!��ѐ	6xe!�#�.��ӛ ��ڦ*Z�֙�]q�iAh�CX\�e�[�#����q�U�h@s9.Ň:p���=΅9�u)�L(���%�˖ 9�ݴ*�i%��X�F��F�WD
����鶀6��[o���;n�M�9�ӝsr��L�E7p�a�ڸ�{�����n��tph�YP"r읮hi��ms8�f�*
O��G �K��D^���ksҼ��dCi����VX⾒��H�IWH�op�`� �j�<�U�+Lălr��\j^t���gH�d����y&�Ւ�p�*�}�_����u9ۈ�{v�#��cz��{e��3����t��tr�Iǎ�q�j��n&%���@�ɋ�����C�za���it�1X���8P�E`�RG��R��GWG��i ��,������`*\�뜖�e�<4w �>�i�z�nSٶ��� � �Վ^;�u$m�#���������Q-���M�M��L��Y�4( 9v��Φ�	��Y.��Ϲk���o�/�zl�m�9\�k��.�P��uƞ?������i㾸�t�M�<�X�)���ah�ZQ�r�+n��	���ܝ�b����������O���Z�Iֺ� W��Cm
Y���z���vB0�M���tN�[�rg�pT�f3�U�$�]aj��.���g�-�09q%�YI#����m*w�.+/5��}�)�1��j�CS]ڸ1��, >���k8ih%�]�-Z��ʍ�*g)�7<�&=��[�/\��xF� f�R֞���e���{#QĠ�N]��(g3���d�Ma�vp�g�4y/x����??Y��h7�h�WM�k���E�:��y��o
�U�n��sqj�"�zv�3���8Fud�-�7T��:��Ġk/�r�?�'/�p�4äu<a+%PZRuër���޳�b:G��]Ej��o*{�c�S�uS�SM��F�˞�˯k�=�n�]ݰ[�\��G\�ьu=�_h�����Th�a�b;�A����*�M!�U�m���G(�����1��ŉ����/�6�.q��ě�/�Z��H*�A֯�ᦇ'�jӽ��6l+�Tn��r�7<��f�A=�+;��u��C����˰]X����OG
��-��z��0S�7���c{�r�f<?#gi�_b���C���QN���4nc���h�7M�4���5V8�],�l]������\%�f\�d�k�y+=��������a�q!{Ӆ���rŲ�Ϩwғ�N�/	�*�r�%#�N\O��vEu��*��z��
�㙼�qM�����b�z�t��ͯhd�%'۴�)���W*%%8��!���;�U�Kee-���� ��N�j��M�tv7�b��}�y���*�]���_�u�"���ǲ����h?tS7�+z�̘�u��n��.�m;L��>�B����Dc�z_t�j�"q�a�M�@A>2��Ȱ�|�o<C����oR�,%�����i�Q��?2+u'�7]��O
�	C,��6��e��W�c@.܈��i�G-�+y�6����R�M�E�j�G�h�č��ĴW:\q"�+e�~pP�%������w��&'X�{���պ�Ԡv��ڃ�&�rؕ�..=��"�bמ�9f�Ƌ��ί �-�J�&�Vg=�C�r�i�X�;5x{����_�"�
���7���k�]k��p������6n5��D�9�Mu��!uf�����V������LY��ฮ����t$
���Ѣ�|�F��d&h𧽜��GԺoӆ�˴+c�&wk�.�Q�4:ށ�-�BN��GUr���]`��"�� ��
�'J����t��h/���9�8y|4�����>K�����J�t�y�ψ�6�GZ��>یg�۪����f伞��z����ݰ�gr��w"�{��j��J����Ugˮ`U���D�1Q^>b��Y]�T��z��X�6�jo�2�/2�����%cp(|}��ݗ�;T\�Z���j����{��Y��-I�� �n���{�e�c����97tnf&�$��Y)3�G��i�����jf����ӥ�b�������[Hm�2�Қ�A�}Rm)ac4�iZʼ/=���O���t�ZZ׺}�u��]襡q�P��*�+wH��RY�anS̈́-��yy/+��t=�]n��y�m��!�EbS��:(��[�V�56r�i��8�m7۞����UB3��LO����ܷq�G5ޤ��=��$��<���W��}�`�س��e1�$=Ɲ.��n�[}ϧ-���S�J�9��ْ�u�Y @��Ga�p�ɑ��~'�����r�4�N�ߗ���}�s��9����u�y�d�C@�?|H�	k �#$(h�0(r�̚B�ihi3 �r3,2r��*�&��&�̦ "����,�1��+0��i� ���� *�C(�ª�(2ȳr��2��+*31�JJr�3�����&��JC#3�3$��0r����2p�h����1r2)�ʣ,�1����"%���2b�̃*�,��0���3',(rLg!ʲLk�ŧ&`Ȩ�����2� ��� �̬�� �J30���"3*2231*�C+��2r��h�+3#&������,�("�#32,��+2
Ȱ���#'	30Ȣ�+#&3
�̙&�'0Ġ����$��%r����(��������ʊH"�3�²�"̥3��@�4I��hǧ��Wnw+f���a��i��������!�z�8��s��g�� :�m;G�v�.�a��8JG�ӓ�	-q>��}�T'*�ʭ����F�d��Q�E���H*�yݬ6��q8<d��g���n��s�Y�n����[0.��t�̩^u�it-�٪{�u�Ss���s�*�Y��;0��e4K�>�Y��>��'ޫ��Z�f�C�ޑ{�w��{��d��(��lY���W�k�2����.|�ɻ�.ߥ_�2��i؁8Tc�v'wHm��\�UDy_��YK�F� �~����Q�9Z�x��DuM��F�_I2�%u��l��{������d�����Af�����3Y�7ܳ�/+9,���+gr�ƸO���^��,y/6����K��O�R����ݾ؎�����]�-��o:\�3�Ols��c~�"VQ�8)w��U�3k:�t5�|�M�
�c9��oJ�s�<�p9��F���ڲ�3��Т=�����s!�o�����;�q:��sV,��~��	���w\�`}�T}a�4���y죞O:J�̔=y/����z)����[
'A�ig|8�8�ꆅ) �g#n�䯕���3U�CI��ՆQO��D���FJ㧏�"S�٩��hK���6o�t��Q�X��7}�}��{�/�}�f��b��L���I�+������3���z]�Jcg�_/O������ϧ�b�����\�����T��鲎^�%sed ��`��<�U���Ϥ���]bzЯ���v�I��=��n���Js�_˻,��NX��X��6�L�4;٤-�<�)�~���o���ח�C��L�y�\�`�{�s�佬���Z���w�����~�e�x��[O�B���Y��jg�?_o���>Ac��+}K�v1wzī�X�N���U�O�e�o�����W
�'!�)ky<��w%7}�AH�l�sX�:��������r�=؍Dv	R.�z�T����Q�s��M�:��Z���`<=���^'��W�{i׍���q���G�v˳����q^<`�(��+��W�����*֛Ʋ����Z��P�^����t�5��`!�ߗ����9��em,k�I�-�Odq(N��<P�Eo��;�)��)�J�cѤ�C�)�s��l7�{A�c=�k{��'^eK����v�lH�ٯu�^,N �.3U	�E?'��^��g���d9U�{�yմ���z�~���\ڮ���t���=@�[P��~~/;�z�Ç}f�U�t/i������+;��|�qɬA��њ\��Ed���7&c��mW`{{����s��gCc'2Rö�rւ�)Z�Γ���{��x.M~����X�:v�B�/��>�ݚF��Y��9�⾓�ߨO>?U��1����F�]����u;IȞ�pt���k7������Md�s[��zcS����9�_�2�����R���-�~�t�:��z�ΟS�jq������纬;��\�5��7�5��M�����'z���7E���_m�҅�;
vY}��������҅c;4��Ƃ�=�<���nu/��a>�C�_W�gg�[���h�dsW�W!V�Y)[�\6(����F@M�S��s�#>���3�9�L��yKU��ى\v��-$���.�ou1K�ѕ\�P�R�<��\�p�����t��	����ז�t��*���E�8$k+�xF�r0��J�scG��>��Uo��[�a��<�Zs��U���D��.�a��%�{U��fW�S7�ˏä�=�I�*ı��Л�Sr�W0߈�A��D1��\���ni革����#�迄��U3�^FXF����\�s׎dd[�rD]�3�.�� \���~��t��=���7N�]�ZG�n�����k�:❛�T�q��ۘ6x���d��3�}S}7�=.�6Ҷ;�ݶ���c��xX�	ך)�ۏ�1nJ��.��fK�[��ט��l��3�ѷ/S��U`N�Ǌ���p�����Vw,�6#����sw�=����Ѻ�c�I��ͪ���4I���v�zlUfڔ}ϫ�R�G���.vMs�����5��g9-���ʞ?R�V��X3���ׅ�riü%I��Ό�ݕ��}����ԏ4��L��r�@��V"J�ҝ�:�":���{��\���w�P��_I.נ�=�r�බ�[���o�:Qݠ(c|���w�q�zPPݤ\�/a�wvÐ�N\#�*_H���E,i�	�m�-���C��Zz�*+�I��w��]޿3�k�/W��(:�39�x�7:`.s�3<�e�>Kڝ"r�z<N��]pWj�/��o��
���ю=4���ǚ��U�|����^�1}:N=@M��D�};5u}\g^�_L�n�ɗue�Ǝ��ݗٵb[}~��Mi��"�<<_m�Ҿ�,���n���Ǿ�}Wɞ�ܹ9�N���u�sC��E�x�O���b9�,�j�&��T�)o��k[�ry���r_�T���EÕV���x��z^i�{r�������K�e���+Cs_���؟�S8��N����8��H^��^��Z�4��K\��\u��p�NM��W��N/ށx[?��[�Őp����js۫��[����B)�{=Hm��rh;:k��3�2��ճ���7>��ߧ`�Y�j�%d��fm�j�d�<����^��� �/g�����4T��gS��*����W���W��&W�>;�3�`xr�x$ԥ]6��G���Ͳ �KԱ����X{p.�ߕ��V�l��|h�ε�B�*pŚ��ٽ�h�<�������-V�]fb\����/�Δ�ך/w;���g�p�s��&s>��~0oːY��U�Gl�Օ��9����)�o?V��]=��~��y/6��I��3O�fB���R���>���`W>7�X�t/�͐o?.w��'�c���ɺ�\k�^3G,̊uy�����v������M5���ь��(.v��W�;.U�D��;R�%��otg<�������x�M��U��6lc�Y�6�\y��ɕ��{`�~ʫ��nO����l��/KY�%��W���-m��z�u��/���u\�'�K�}��OW�s�}4�o�ӛc���{r�޷W�����-�g3�j��c^��C��ھ����y;WM�����I'�bv��ŕ��������rĜ��zM�:������2ﲹ���B�'ϴ񰻴�4_~���{:����%�K�'�kIb��	�b����z'J�lo+'���E�ۺ̼񧞞�r)Jt��O�+C�-�r-K�Ce�/��x��j'�k�?r��s�f" ��^Om)�c��1�(�HA�%�!_����m��ҮW�q��}�v���s��<�V9�B���y]�ιz:,��_f�K���8gcw@�˻}2�=ݷ��+���Mb5:�7)s�=y�=���t�x�W�o��7�v�׳|eA}`��$��6�`��_��7+���h�e���n�7Y9�����W٬t������̵c���v���F�ye�fY�簮 �w�2���w�;��pܚ�p��ٞY��ty��+�ǼnH7���x��"���Q�}L^�}v�X�����z�AY�i����9�����}U��o5]Gz�ћ��K��^%L�&k�w'm�{;''5��%�R��޿�ʜ�
��
s�����hگ@�v�:�ɡᗳqϖ����=ӧ<��﫳,t�O���Kޮ�i��[^�
�НO|�Ov��7������7�{�$���O���.��ͤu��7��XW�i2�`�q��+z���ӎ���飅J{��ķ�� v����\��*"u�-s�yK�y���M��s
����[�.���Og��00�ތ{�\�K5��5�+��z���h��p�0к��D�oo��z�El�yY�c綕���Ԧ:���� ����Ƨ9�3xN;��)]�-�h�y=����+>�����:^�F�w1���]��nBK2��қ�^�N�s�'���h��ł�l!ί��
v޿k���u��qU��"�����;l�3	�|!�vE_C��}��J�ߦh�������m�2�{���vol��������u�&�W��/��S�B�����Ykm����&�:{���%hM��U�a�F�C���^{�\�W����1�e�}�m�_���1�vl�.���z.I�R�`k�V��-�����g)ہ8�mX�+�v3vX�M�}���{s�W[�,4:�x׻��دF�u=/ג�U�w�n�϶x���C�AI�~��c��/Ww�/�b��A�/�@�x�Q{~��:��H�#�㝾@ˮ�u� ��5&[X6w*��y�1*���ɛ��)etOGOC9ҹB���T\�+��'��Qᆇ�9^��������d_^ɇ����D7 ��|=qy�z���e$���B��zC�3ګ~��z�5�0;�L�_i�nި�Ǆ� <�5=˽{\�;?{��?5ry��-�W�٪���Vuy�Ӯ}��i	�{���i�[�v��k�ߧF���w�5��v�7��R��jI�G�3o�:�/7����s���'�9���;Ƴ�߻�cP,tŅ�>Cx�����}\hn���X�Q��_�N|j�5�9����{s��:h��?E�� ���Z���c��4sf�6����aÕkwuF�6�*�{��t���1K�ǅ�_m���u������ӽ��~�ꆧ9���z{n��s�Ǜ�ǫ鶝�<,�hs����N�i���;���6��;|��sk~�ޜO����[�s�gP�Ekj�u-�����i���y�.�����T�zη0?�E�e�*/n�BȽ%<;ե���ٲ�����L~������S���Tsη2�;�Hp�����UU��Vh�2�o�$��H8��}�����zv�T��<o�i v��왬}3;Tچ���b�䮊��7˽�P;�n�#����g����=�Տ}��x'uXe��uף{���^��Ax�<�^�&��E�����⸏f�p�]/b�:�ô5�;��o��h��j��5^�/�bn_kj�Ƶ��)ޫ��Z�� 2���Շ���[�wi�Ezt޻��4[�d���,��O�pS������8eK(?X��C~|��������$ǧ��X:jـ�/�ԉ�Y�w��M`J�/L] ��̯����;\2c������^,��k��4y�滌k��yfG��ZΕ[����gOj1�׾Kͪ�I��>��&U������)���:��8k�o5X_S� �7�.w�rkc��&R~𨷾��J��r��2%��1�O�B����������w�i%u��3��l���{rw��onj֗��
�ῳ�3,O0=Y�h�PN_��y��$�__y�	����M��i���Թ�J��7�l_�F��X���l=|�2�sw�@�H���<�$��>̔j�Y���[k+2�ձ������9���T�*�wk7�:὇o*	�bN�s�Q��iޝ��Gܴ�՛ʙ�A)�m8��|AXwY��啙{���Eފ�=}�ަ2�x�nwP��p�5C8Q�<�n�c��G��M���U��-����,��s�%!�]AX�i\�yt��4��;��+J=���B2���{JDj�*ۡ^�ԓ
�!(Q��C3�A �=z�©�r*���DN���-���y��,�'�b%�[�}I�� �먎\9���>�
�*+ήo����c{�/mJxF�w|��ꗊB�ҥ+*JÙ1k��h��v;�Tu��vМ5�2al��dI;q����w����¢�HXs�Un��g[r�1xA�Vy�Wֶ��*�k��P��]*gM�V���H�)�-w�VV��;*��H�J�v�ҥ���N�N�I���
q���C�s6݈^�}��,/�[Y���6��b4Y�@5sK�[�T5�	{�����QIᤜ�{Sm��ڭ���u�[ۇ��;3Q��X	,R���55�#!"����,Y���e�9B�Yß${��5)d��|�s�]i���8[���ȟQhs�[��w��O����Qof���ǡ܍�j�4o+�A��}v��Fh��H՛��'�]؃�%���H.S�.�����Jc�qb�/��l+CWqp܅�oޞ���_rI��r�Õ|�wSёT�[٪/oS)��2ɹ�f�h�(�ٍ2��2%�/w�ڽ��٠���q������E�5=�E��T�~^��e�
� �O���ͻ�fJ���\s��9�O����eX��Y	@v�t�ju�X�n��$��J�3$8����VF����*���e6��^\�۠���;l���n�k5�Cr��}1#��ۼ%Rd������`CS+�qa]��B6ڃ����[����ھV�D�g�ZC(j�&��RPY���ta��]q?IC#��'��/���k"�_Y�81��aڣ��r�#���������R�ܵj�W��,z�/���e�Ӛ�	�<x�����SX�!�=&]Q`;������}3�]U;�L� �[ԥ,�@۫���a�ъ�����	�$4�Sph��ۈ;T��iR;�e=�;�����
�ڸn)] �}�ΑͲ�����GY��ش�(f���yF�������5,]���*��\�Z'w�m���O�8����8U�.�9�SG��⮗w��x��^0�M4���Z�pŸ}]��a�9�����9�N �s��]�s�Y�{� ��:);F�,�[4�1�p}����4��r�R��7�j��N�"%�Ã�Mݚ��v����%.�Xz[��y��釲���B��@�Pj�,�
21s3$����h������2"��23#1�0�r��&3
I�#
�# ��i�(�(���3��,��	�*b)����,� "(����Jr0��*"�#�0ʱL�� �")i�Z�i,���"�32�&�22�"�J"b�s2!�32b'322*"����&��*)��Ť"��"$*	�K�'3
"���rK,L�
��()(�*(���$�1�$(r (���$���&����*0�&��(���3# �0

fZ�0�0r"*d����30ʢrl̜����*���������"�"���2j"�c#�,��
���r�0��bl����3��,������&���j"�*�,&�,��2�&30�(* ��2���si]��W	��S���&Ǹ�;=�Q�/��7o��.��:z���� �Ac�Y:�)ElVt����:�ʿv�7���vN'��s�	Ƿ�N;��,5��/7*�椰N����������gL��纝Os����{p�c5�D�;�Ծ^k;I��|V���@�ڽ�\�����mt�&�(��ي�L&3ӱ��|׼ß	�E\����*����\�gS�nu�O8{���r�R�Hi��A�۱+�\�M�x��[�?VB���kݏ�]
Y�T������[���7�����8�N6���n;ԟn^�0�G7������W��ӹ�佯�91�迤;BL��5�����/ׂ����vA�h��r'7'�L��7z��*�C} ��zo��s-X�cM>���p~���.�}�>��w>��-M4�����&�u��*y7Ix2!\��T����ϐڱ �Y����U�ǃ}L^��ozC�VR��Oԅ��of�Fʕ�M^�6�^�ΗTf+���/P���`�wث�h���p�:�[�j�6��*��p�Z����^XF�S�K�/_i/�ɬ'P� i�`��\�=��4s�W<p�v%�û# ��-+�(�d�ո����*;�7��ucFc3�ֳ��~�yA���l�O~�(n{��gV��S���r���E�	�XӰ|�/�ueoNm}�6k�\�U'X�Jx�����G�O�[)�A�۴���e�r{������ˮ�z��U��G�[���	/k�;�|�)��!�Ʒ�x�3�F^�	'��S�`�t�ٍ҅7�cվ�yI�ہ,vxJ��Ώs[�������7���~��𕝃_��;g#N�m�-�'����(��4������5�p�Com���P_=���p8]M�$g������r�z���]㊺'w�ew�5�ݲ��ە6������5u�vE�4:=��o���s�G����]1}/9'���y��7�o������⡸$�(^æ�nU���!���{�`��ѓ���o�}���`.��%�`&ܫ��3a���9Y2�9Yͱ�n�d[���ЬS��Wku��P��biy�����{\j����]o�I]XD���m�M[�z��6��+��n��,�����,zyzj.�>yJ�6�w��%:�^@�]]�P��J5�z�(�w.R�h>冷uSv0�4�ۤ窲vV�Ϩd�,>�e�9����.����f���>���S�7��_T:#Y�=C/]���N�H��p[����B�m�z�cs�8�\f����S�S���7_����l��Ӌ9�3'���Y��؁�g�} �3���f�xN��O*�}ƒΧ�(�7O�,v�O��/9)ks���g�7n{�|(���v>�d}���҆��􇁘�����:�܏o=���u�}35������p�u/�R�� ��pW�`���;7��G��O����y9)��:7/%�~��7�@~�|��H�!�>�]��w�KA�܇z�y~��:U�(@@��t�����]}�����߱7&�|�R�
_�p�伌��I�3Xn;��}w�����#���ܼ�w�~9��CP��{�ݣ􇎋�S��Q�~�-,�_�w�����8o��w/��Ԏ����NAB���
��MC�w}��NI�ֺ7~�ܞ��r��G��Ի#�?}��9c�\�t����̟}��!�^}�:���y�r;�r~�%?OP�?�ΥA��M�H���p�rC�5��d~qM˹7�9jW��4�Su����9��Uǧ�t>�u�ڑ��]d!�Լ�.�>�s��v!7����pR~�p~����WPn<��ܮ��p�rC���߃�0|�q��x�ۿ	G?,tۗ�Me)�O5h�����[}�����z]�D؈a�޽���sv4��5�)b��Z�]����<�)����cr�����죣'I��Yi�Q�O����5w��Z<�k]�S^\�]s7�Ô�wY3��ʥ	O�}Yt����jG�|9��C�r>��Y!�7�Ӛ�rS�>��M�xs�����
O�9��<:1]I��� dY������%�*�2ߠ����K߸�3�y/��=�܆��߽�H�/�����>G9�jǒ���R:�����(�7Ѹ2]AHϒ B>g�F o��/n�t����N���W�瘚�_b�f%�>ߤ��]!�A�s�������캓�瘎��to�v�����𺫺����{h���*� ���\�_\����xu�~���G�F#�Oo��W�ߘ����Nϱ�!��'����}�m�������_`	�o�� 2>���vՋ:'�v[U���߿k�����w����2�9���u9/�`�]K��Ԏ�?GϸY#�;|��9})��;����kX�>���g����g�<�̟����������/u���J���Z�A�_9ߝ�J�OM��k�d/o5�!�w�!��]K����r�����Grx���9rS��ܧ�uI�sï��sF����~�i���R=��<G�?��Ϩa���!��t���)���!�^�s��%y'���׫�^{k��׸��`�]C��{��Ga���;��y��޳j�\����û?�#��0��4�������tr
W#��ܼ����A�;�����BP�/����=�z���������C������~�����-�g���w�=��9��@�qc�yy�����tr
W#�}ѹy��t���97�}/�����B�����z���>��W5�����ԭ����y�>��|H������q�?A��>��������y'!�5������/�n�z��y+������<�aܿ}��b��/������c�=��S���gHc޷��E�)�}y�[��/r�<v�ᲂ�V�t]A`��vX���"�6�u�D։�so��Tٖ���k̰�����2��s�
s�����4��^d���˸g>�30�<6ծ���1w5K6�w��ڛ�qǕ��?�������wr=ǁϺZ��Sܧ�}O��r���j�������V��u���];�%}�o����#.��v��׈��i��wR������ѡ���t���������Hx~�ݎ��O�ش���G�X�W����pR���9.���P�NG�:��V�y�w'��C�?@�LY�J����t��}����Լ���0ܼ��R��/ 5�׽�ؿHxov��A��)�;��xu�R���xw��)^���n���#�i��}�Zv#BC��_\��������ӑϱM˩;��9j�zf�y�}9�����}M���9�����&�s��O`��!�~��`�(��́Q��-�n�^/��u���o�&Gr��z�ܿFH{!����)�w'{��������:�#�j�C��}9��%>�Q�{��!<���2]�I�x_��^{����y�?s��^��kqA��G��G�;��7���9.�%>3r�^{����ܚ߽~�ܾoΎC�����jMǒ��v�J�w�q�u���_Y���-����:�����	��u}�?|�JP�g�P�;�Q܎�ΰ?K��O3r�o�{��p��s�[��_���O {��F�+��{�~���޹�5��Q�x�v��<�v9��yK��rp�g�Gr�;�VB�{��?_Jy�nC��~��]�&�>�Y��e�޷����y�^w�3ϴ~����p�Gp5����/�ws�pw/�}��R���s��#${<�G$�u/�X�Կw��x�����r��䚇/�/5ݙy��o�{��3��%;�7�?��>�����}�����k��G����&AԾ�O�s�9�|�~v�!�y���5�$�u}��]K�xu#�O^ǻ=��Ϋ�j��{.� ��!�#/�w26�$T�$S��Ǆ:��d��ײ�+�}u�=$�s��K̧���t�Ǩܾt��R�>@n��3^g\�S,���=�J�t.�xn�Vm��d�ݾ�Xu
�b���l��,o���zغS����#ﴁ����)���>���N���rrW^���ABo����)��	��o9�o�����^��FH�K���6o��_�ez�ŕ�������>��~��@j|��w��}��O���'^{Ѹ)\�>���y	���Pn_�$�0Ja�<��G�{q��g��Y��~R�7�չ��x���Z��G�� q:�䆡��=;�y!�w�G$w'���r�s�?A�v}��AJ�v�����O9΃�7/��9���z}�.�ۿÖ�w�+߇��?|�u���W���k��q���?_�(9!�>^���	�Oc��>�%�;�߱Aܻ����}��w�tr
G�5�w�s���ʶ`�_�?wbN�F��]���ReI�_���:CR�_\�^+Ծs����/q�������Od�:�;�䛑��>������A�}uV�^w������6�b�E�~��W_K��Z����oK��O9��ܿ_C��������9��@y���:���<��-�ԇ�c�ё�؛���}߿nl��#��e,�Z���ϿY���(%���d���;���ѹ�Gr~�9//dto�n���Ϝ�y!�^������Ñ܏���S��~���L�xg���[�v����f���H�O�j
�� 二��I�w:��<���ӿخ䵆��쎹�����}�:^H~���{��}��Zp��_�}����'��5?�i~�P�xu�n��a�/�7=A�)]ɹu!��I�w}қ�pk~���+�=7�G!ո_N~�C��u��z�~y���O˙eN;��]}]i�q����&�<�]'!��f	�5/ё�:�q��'�]Y&��d���n]K��=�ܻ��߽~���>��z
]�����Ž}@�ҵ{
�gm���k�>�O=k���~P@�u�"���Z����%��5��7/{*n�*�{�E��O[S����z;��ֵ�ď#�{���|�1 �H�:��j�7��?��[R�y��~+��<l�
�!{ϸ�W�k�*ÞVߡ�V�}�о��7�R�'5�d���}�k�|�N��u�b�R����w���ϝ`r]^�xf�G�t��v�����g�ܦ�}���� ���8y����>wΟ�n9#���Or��>�:��o�� �{|�O �u/�X�ԿF�����&��~�&����_��sݯ�o���!8f;��>ڃ�b��OƷ֮@���Ө9��/�9�<��y�}�>�>�r
��u�r]FK�����W�5�qr����ּ1�>�����]95�����P���a�;��?_��]�!>�^��<��~��|�y>C�
z��=��;�y�·��>�D^��(X[�uݿ͚�~���G��������_��üGR���p<���{��r�������y�t%u徎��&��A�}�����_~��}�{��>=+�=nT���?J�?����rG�7:Z]^�y��?C��x��jC���B�$�c�?�����>{��9#�y�]_}��H�$���6��o�?�x��|(<�q�o�S$�^罞J�C}{���+�K]-.�`<�r����SrGǘ\��>{��G��OO/����Zr��ο����=iG�߸����?K�(N�O��_ђk�%'������W�u�z^��y~��4>ߤ)9!�|���7	�������#�d��L���=��ݿ���>C�
�}���;��G �~�~�p�rS\���w/��=�:�����=�R�K����]���CC��C����8��;�O�e�;�y{?<���ׯx'�{�#�u/�A�yh���ٽtr<��}~�O!�䧞�r�]_��������>�R?�4��>f��� ���FG��	W×c�x6wd�k�<��Q,����X5���b�����}f��9���A�J��o�VW���yT�Z���Zɉ{�I�6�j�/�ykn��`�	Mc ά��fr����{y�W�0���;X7+�|���=�������!y9��5&�{|�Aܼ����ܼ��}��M��Z��y+��o�O%��G�������|Ͼ�~H����y���3����G���!�[�����>���u/���y#�2;��P�=��9/ �<�P�]�G�:��~z�F�һ��u�����}_~�N�.���<᪭�/�r+�}������<�K�C���<��w	�o��qܻ��b���O�gR���y�&�uw�&���g���w�B5}����9Z?i��#Է��Z�~��8yw+�s�F�չ~̀�>ߥ��]H}�}����'���7.��0M���Ǭ�WPn<N�9�}�~�����'g���K�좟VV�5�Z����z�w����5{ѫ�r�o}�V�y��A�Իy��!u=�>��M�xs�����
O�9��<:1]I��<���6y�~����g�����}����d����.� �}�rCpo�?Z��_���?�@��!�7��{��#�5�<�r }c%@G� ���+����j�����|;���?f���u��:1_�������w�'�w�)�f��>ߤ��t��9��F�����jNG�����=�O���v����y����߹�g=߽߆�K[:��h]�� �>��u���I�|:�7��<�G�����咻�$�_J}�;��?_��X��=�Z-�������<��)��|���єj�\�����z��x�����	��C���ר�^��[�!��=`�]K����#���Y#�;�����/��(�����|�����f�����7�3���俤��Ġ�_`����<���뾎�y&�ޗ��_��\�%�؆C�u/�wP;�����~@�#���Ղ��n3�|��U;�o��5��f�~������_X��	{J���&�������l�̵��I�n���g>{l+�����2�F/����J/(ǜ��x���8����&��@V�^f�Fpl}���!˧&^��*����y���e�@^��Z��_���d����gޙ�<~�a���οtjH��G��
C�|�(7/�S�7Й��tw+�>�^��^���-.��?u��u����9*�V5�%�T�}ֻ�d�4@���p7'�亃߳r�9^�Ѹ)\����9/ �<9΃�w��=�:��{���y#Ծk�v�_J��]-�?���Փ�X�C��Y��~�i z�O�O�=�����!��C��^A^>���;�]���������>�O��Ӑsx���/��=�P�@s��9�����=�}s�y��pz���9��Z��x�'$>�Q�z��Q��/$�:b���wx}���ޱ�w+���9/# y�>ù~��o�<l�����*�-z�?۟���C��{֤~���~�uw#�o�Zm�Sܧ�{O��9�|�R�
_���K�+ϰC�;z�N��_g3��V��?f5��g윤������W�
���_��x�ΐ�_���������v:���>�b�~���u��~�� ����K�)|=��;�����~7�~�3ڧ���~�߀��}����F�ے��%�쎷΍��[��9��P��;�݋���a�����~���u�R���y��z�~y�W\���ȭ�o޿��\�_�,�����~�2>�u9��%䝼�G-B�Os}<�w�>��t���Ծ��K��r=N��h�y���w'�d���_c�{��Ӯ~����Yw����g��A�p;��w+���r�2C�pu���Jn]ɿ0��p���:�#�5t���Ծ�]&J}����רy	�>��=��w�������f�y�8����s���<��C��MGr��:�ܺ����˩y�қ�rk~���/r��:9�P>^�!�7���=����Ǣ��~���� :1L9��~[�^��R߰_/0���|��+_d� �ǯ���;���5o�Vk��N��1
UYy�N�v�j��+��Ư�n,�AE�q���@�c��>�m��\�2ޮ���Է�7/�Fq?'����������>�| Ž;�/~��J�>뾇�(���.��0C�~�!u���MGr;��?K��O�ܺ�����7�?~�a}g�dKx���g}�7�����<������?O��k΅�y.��AJ��o�� �{�]<�%�d�u�nC���b;���y��!w>I��o��!�~#�<@��{X4Ͽ~��P�z��4w���w��	�A�7������:O��'w���w�����)^A��}��d��Òd����X�Կw��x�����r������|������?u�\���߾��� ���{�	S^���bH�	V%��3a�55�>�ՙ�3��ty����[1 �>�5}���<�C�&\��fN�4���쬿���)o������%IB�]�ݗ��W׌�H�A�"�nJ}y���~��v��հA�3ל<����ѓN�{\ �K���o��1��fFv����NAg��w�Q�9���O:��G�t�{�]�|$}��xɚ�N�W%ͪ�I�����7�i��@{�ի:��Z�7�X$��-�E�۴Ƿb�~���N��{2L�s�Uv��0|(J�ݖ�~<�b�t�+&��]m������^'�s�H1�	/úU'W%�p9.HK�tiU��Wv20� �ԩ��,��V���0pʽP���u%��J�\ LQ�2��J��Z8`���[������Z�Q��1r���&l�r'vމo��;1P .
�R[Cx��MG�	�Pjf®�p�g�vH�W:�u��db�A���ZY7��͚Z��:��ph�JɆ���	ǚc�"m�&�I�B��b.��3�ci�1:�β��]��=���|�����<^��9�k$���{}i�ț��%K����Jn��9N-]�7;�U�����1;_Gi�"'S��21g�2�Z�J��F�JbLx.�X�Z�M�j�w�]d�0��sL�LaC�s�K7��1���=B�N��H:Ue=F](�\���D�S`�羫)�|����dl��i�tJH^w*�R���Ķ�,�P:�6!�� �Qd��(�-��s&x��]�O����V7X{i}4E4Րo��9n�����N������<��ۚ�*;�ݑ���:Q{-�X��t΍u�-R!k�
ř2�0)o��'h^,̭�OU��f0k6�k��V�NTc4uL�5�}�4�̴�%�����Zv����E�,��uZ=Ҧ@�v.A�L(s,L��ZP�Y��i���t�
t�-o��ͷ=#���u�L�~� ��
�m�R��3,�ڵH�Q.4hl3>��NP���e(�@$��%�q�����G�y��l<���ғ8��k�0���ڻ�z��e��g�آ�}ME��=;aB�� `�.--�a|��}/�p�^>Λ����ԣY�Gn�p�P�.*�U�����i�3YjT�j_^��F�̵at�r��-��qbt��Z��M3 �N�r�?e�Ց�p��".  ,[+�T,�V]/n�-��x(NC61��HŞ�b�C��Ξҗ1ǻV�<�QEӖ-�j���G�M�]�6,ߘ��r����CY�!�o^��6!8;� ���]���:nr �����#G��0�L[ �+�C/E�*�:(��tۤ_v������Л=�#��0����uˡ�A���WU�{�w#�w��X.,����}�釴���0&c�8��ns	�@��<ur�Qz)���9���EI���Z/#ޑ����KAj[ML:�p��oj@0��y��U�����{I��j�)��ٰ�����\�vlY�GN��!H����ߠ���O�.��u���P�ʦV�E�kA�dHG���xu{[�*�7�	�N��ӳ�S���Z�Φ+���o�:=Maz/8~����`K�{ec�wt���+���n���Y�)�x��v�Աk[j �'5N��LB�!V�/��e����W�rfvE>�<����ٱ�Y�v�����q4������!"���Lb���"i�p���j����hi�L��)b�"����hh�)"�2' ��`��a�r��+0�������*e�"!30"b�l�2K#̨f���((�	���(��30�*�(�(��$�������*2r���`�*��"�"JRb� �l�32r��������	������*�H�*2Ȣfr�H���#�����h�l���,I��*�"�12f*"�b��r�*(��20�j`�$���j��h2L&�1ʨ�kʊJ�3&��Jh�r2�h�* �"��j����("� �jh�̳��1�Ș��)l�"j( �ʂfj�����"j0�!���Js0��H j&���#3)*,̘����0�(+32�$�,*����j��)��0�<�S���G}~�Y�@�a_-�y����2f|�� ԡ��ԛ�݊�u ���M�k+���������z��q��w��>�������~Λ�g^�ϳy�y�\���p8�5��g9-�/cַ��k��w5�΁⻟�h_��g9�~�.~c���x��r{�%�𮫒���g�e<�g�����^�Pu|hgG�5��ј�A��ڭ�'�ܧ��Ut��n��s�L2�L��O5r|hc������<x$dKϝ����~�ڛ}����ǨM�(H�3��z/��
v-K�AJ<�y��0q;~f,�8v���W��t��d���9���vE�<K�r��|Lz]�W:W�����ޔ}V�f�yo��vT鞽�.�X�0�����u��P���6�#OO w��˙[-b��?J���c%����A�w�q�V;;;�����m�+EOV^�C�c�NߏT�7���r�O�A�έ΁K���G���/�K�e�ݚ��y"�VU�(]y��ݤ/o[�����d�v����rEI�"aŏw���(Kh�h��v2�<p��d��n���u��*�j[R��+S���u����ug"�����/K��״{�^�ښe=�U�;!g���^���~�[�f���jՙ\���|��� �n5��ތ���;BL���Y��7>�9���)o����c�)iv<�f6��ف��N{����^�Y<xy�U�s�����J�Mk�R�غ@�!ѽ��f��fg3�#n^�v:��1�kJ��Kj���Swٽ;:'�c�k���Ξ�T��h������-YA��ۓgW�'Qr��]UL��f���%_S3\7��z��s��'Nw�sU��\v���\u��r[��ʧ�ht��z�c��~3��l;ϳ��{Q�B�WqsV�ݽ��3z=˓_�^u����>N�.ep��p{�"벙yW:��g��j���:`�����9���6[L�e�m.v*WJ��x�D���wmrw:�6�0n?n��;�79������i8Y��go��o��{��&%������)��^��,Ι��y�M�ߤ����]d����y�Գ�ԧ��Շ��m ���b��ĜwL�r�\2e�Q�`��j�6Mx�m��nY��*Z���.R�Q��R��5�(m�r���_>R&��4`��Q@mt6���z�&�v[���zC�
`$�?G�����Gf{�Z�&����yh>��([�g���z\���=<f���G��߆mG�$@	�x6ÀN�*�<L����u~;A�����;�Y�����w�y��)����,�~=��.�����CU6j�v_ֽ,���̀�M�������j5:���O�/^�_k�fOF��<�r7W�Aލ_;��E��Г.3j�<;,'ٽ��*��2�]�.{oڦ[����%�t��z}�A�K}�M������)�C/���۷IC�f৔/[��LX̕����5����xj��YR����f��κ��e\����+���5���+�\��r�^y�����V�;-�<����P��K����F��U�wɍ��y��s���7���Y���oG����\������1��=� ��|����n�'2��V;O��Q�q�0w�;2⤉EZ�>�����:�,��yzggF4�W�fM�v��D�	��	b��Z�v.��j�@Ⱥ����zL�9]�8m��%����ݨ�×&�Q�������P��#ñV�@sn���+�Z*��pj�}����6�����֟�ou.����q��rw�����X�s����3D^�:{5Gz�C�D�l��$7�G:p.=���{�M���i���b�_��6Pg7�Q��[w�!�����@<���6'�ϧ�&���x�d�q�_v��
��
�xA����kt��N�����V�C<o�gv=�-���s�y;ք�����C�_S���t�x����\��Pg�P�>p�;[ܩ�ot�]N`�v������` �_�i/N�ďnq�>G�ȡ��Ͻ�5�1݀��	߯��i���O���H!����a��S篝��sJ�r����`�$v%X�m	��.��nGʒ=��Hɻ�ȼ�TwΪh�S���nI�]Aa��Hsd˞�����{��)yw����V��X쿗{5t��z�r{a7��H,8����+�<ƿ�߳(n�� ,�+@��O�����ϒ��[�ИLl��l2�M��ϱ^S����˦<��$�{B(�U����ظWM��}��
r��1΀(�0���w^�dW4{/9wQ�s�<i.KTzC�EoP�_T[������U��}��*\7�fs�a�t�sս������^�'<|m|�����'s�e��k}�~07��	W�<��bʹ��3��㚷�i<ꏏY^V_���ͷ�'ӹ�S��~�W���zM�Po���N��/���iƦp���.9t�8�l�X'��f�e����d���s�Uv��n.�c70I�}uL?N�0>T�3d=��;~2g8�{~�;�Ov��%́l��>�	�ς� ��<s�y[1Ďk�ͦE.~���=BqSz����q>�/�~9�����㌗u�b�!��,t�9��M��J�uC;�X�a�ML�}�p{�f*r�d���1�S�[#炦$ai�`�&F���_����թ?���d�н���������a<��g���g>�Cܱ�\ӎ�e�b�lƗ#`�x�A.�RL����n�^H'Tg�T	l]��B���,���]�������M,���_�@�Y��64��.��η֊Uzw�����z����ܱ�o���GN^�f��N�<���p��X���]�W�^X��]Ə��������.��y��q�Nɜ8�*�b��3�d��s��$�+ɽ�z�M��q\mΥ�HuZ�~�������;��������?�CCm�I��V��>�w����l�j)jU����;t�{=�/����d���F8�v�3���x�u����ܔ%��ʄ:+��"Ζ��M�����.�$7�z��q�Z�xK40���q����]�L���K=1Õ� }K����V.u>�*]��V�	�»VR|�x.ف�s��X)�_*'�o��=X�z���ݚ�*3㖠6$�/}:�w+��<If��CmJ�xm�C�ʓ��fna��zݵ�;[�졚������1qk�g�e�m�fb`�m0aee\|n��jҕ�W5罢^z���*P��"��c5�ĸGN-K>1�l9��>��zmg�*���xv�7�*S����]q�n�#�dE���3�6�(d�z�ōM�x����ё��ԙ���՘��4#eȬmY�|1�x:�3�M���>��o-65yź�cS�2<<�ǳ����5N�x)��opZt9_�!W��sz�k=l��]ҽ���S��(�m����/�<����h����T�+����7]ՊҚ[�BjDinfY��E���˸ޙ�!�o?q�c�E��b��m�C�{���J'd`�9\�U�9tv����v�[x1�9M��)���0�w�Ͼ�>�]�z�`��ǖ��t�i�=����.��&\�gҫ�vR��]1C�3��Ƹ��n�*��>�^Pz�f�s�	��q���;�Z.z��*Z��P��US26���V��e��ŏK4EJ��Y�� �ڰ��Y���Ő�bne5�	N�`��+׻ǻ�q�s��\ٙ}慎b�t���=�/_t�;�C�VN�GeA��M���v���9���+Z��	���"��΢�|��EXu�:��W4<r�M�9�z����T�.�[�z��ۼ���{]�|��X)>^TxnT^'��G����J�7^Fml]N�����nF�V#�-�g��	�<lI��b>ӎU7]���\�8fQ:�m��ەל1��٣7j�]�-�Y���>���a�]yZ7!�F˧k���׮h�:��ѽY�+Ӛ��k�ִ=U^�>�B��2�9E�	)/�=u�V]b�Q"ȕ�a�����|�Ct�wj��{q\�%��X��RJ��a^������͔u[��Q����,׆��^>0���m��]�vB�*Ê��\vr���+��>{���C�XNT>7q�4ƨ�
A�w��Tf�j�p���aY�^�x>-��Sky�f�#�;�ޏ% <��t����8[(dj�u����j��
���n�Yb�]7���  W��҃d�|��������pj/v�>�Ze�9�����$\�o�h"��=o�ٔ皮�MW(:f�W�~����8թZx�&~Ԥ]�����+:Wc%,��(���wbN���R=�Ǽ��O>U��b�;.Q�1ӫE^��>#"�pdL
����-�:Es՝�B�Lz��N�Fu����'m�ٝV�6�z�*����W�M0���ϸT���ԅ��y/��W<�w��s�Lj=ɐ������޳�i�NSw����`�ڞr���q�֛�ݓW*o�\[+�3��K�i�/�3�,COh�z�:�y��N�LJ�x�յe����˳�NH�t���{;�'���k��{(�3��'�������^�<d�i0p�/"��N�.�=X�Fje�{��g�Rը�IV'���b�}O+�p�=˞���B7�S��C����pWT՟)L�Et�y�խ2�����לN��~�c�s랙˦o�i'��zl��H��#��(tW�49��{y,xϽ�u���SK�9j%G��d�����y�%D�d���ħ���ӵ��#�#̅ڧ�Hr��� ��crY�K�B��*%�\y^�6S<��p�����ӗx�?
ް�;�s����z�|���H�����A�C|{F��ۯ~ |>��-�y��q���J�y��KC�ܩ�of�8p;�p�		��e%­�ϒ���;�ފ�-���MT�6��:����Vu�����9J֌K�K�pŕIe.��̯97{+����{d���˅"xm�����D�XΧUV\P���0�JX�W��b�ަnu7�oo�Yt�8���E�7�l��S#qC픊���*�	3�g��n3s�.��I8�������M�����&�+�`�L�]æ�z�61e��(t��uN�.���ȫ�^N�w�F�b8֗䳥�K���HM�9)���@x\��*zd����A���\�y/����^�j��r�Zn�N�+J7��߷��R���-����HJc��=������^"���]3�������^���Je�r�ҭ尅෼����D�h�x�+0/T*��&������a&���خw��)s�@�8��rK��u��s��W����N�|��vi��g�_S��R%�������M�8^��=]��>�x�w�6��+ܯXB���!U<ݺR�e�6�E̜�n���exoF���O_3G�Я��eKL�Sv5��eoݻ�cĺԓ��J�zR�]�uϵQ[�,9���n ��O���y����^5��L	%s�:�$�]���UW�_|:�:8��x���~��߾���xug/pԝ�J��������XΨcϝ�73pn��>eǻQנ�~�l�Wv3�q���:����f�8L�$�k~�v;)�%vh�����O��s���z�f���9���8k�z#�Y��VM���lA.f��;*�þB�9Mܿ���s馐�շ�DȻ{�CM�r�\"��v;���y�lc��Q�#b��Vώ<�[#�A�g�/*o�>ʿ��q�}[\_-�ܭ�B�E-h���o�������m���]H�-L\�c�߆��P��l1�׋Q��/2�BZ�2��2?g���LPk�/����X�"ۤ���ʹ��3몇�^.;���ue)��o��Ů�n�}��ș�*y�>�R�q�#b|�ԻS��0�y�>鐥�3�Ę{��w;N�M���=Z`���L�21�@Ǆ��#zCmO�᷉h�Y|�Q]ot�ju0����e�?P���W�>란��\Z�d�y�؄�V=(r���9�Oz%3�gb�g�XD���SL�=;�ޓʝ<:�ܠ2Eʻ��K��*� <�P'[8"�:򜭵��Rp
�����$�j�f��J�����Y�%��w��9��!Y_2n�X&���p@w�٭�^nʳa#����Wޤ➙��G���_A��͐`A��W���\+(i�d����ԉC\�[���b-�e]�I
øٺY-�M��p`�x���w{-��l�S�'�5δ���t.��X*#i��Q|S`ܠ�E�	�֗D��نU��F��{�XU�\�����0v��a�@nW�£�{��$���5u�K��)�j��Q�B���mP��n(u�Fc�Wt]
�_�����	䧕x57"��=c�XE애7�a����+m�&��g0����]R�47/Lv�N��M��61�/x�Eu�v��h7��f�|.���r���Q�-��t�7�B��m��`�Ǜj�[��̣u'�ԋ�9Ӟ��6���IǍ�݈���n�j��_Mpno��B��q=�_^�R�� ��w:>�Kp��z�]��.F&�}��P���A�6�m(N�K��*'J�����(�۴O_��::�J+o��3�`�Ù+\�8�d��
�	�-��pZ�Tx�X�J( �E	bb[��Z\Lk��nQ�*�ul8 ���Gq(DE�����j+����"��g��'`�H��K�D�0���r1r�jU��,�:��Y��\{LPj��%�<)���]�;\���TC�㉆j���oegV�4�-�bCӦ�ou�U�:�._��1��]�w�f��}�t��V]u��

	��[7#h��9ێj��H�\1�w�;yP,S*�>aÈZ��tҕ�q��j��`�;��zÌ��N>钆l�ÜV;p�b�ӡ�"�c���YP���9�r��j������<�z5N�{u�D)�]���2�c���b�˶�R�RE��BU��T�7{�:��\�뻀k�v��s�� yg�`��6���U����w�:=E��������pY�vQ�46����;'c�
�/�h��d�͝�T�C+)��v��:�귝 S�ؚՉN��^� Y�8��QR���Y�w�iQPW���(p"��7Zqf˚�˺s�^ӫ������ j0��V�+���5т��Kz����=|���fYB�6�q�^���}j�g���P3mњ3��/aT(�8k86՛r�&�Z�N�1|�=����G+}��)2��S+����F���_+f����4�����rt/%[�I)�}Q�S\��.�2����K��˼W�����*|)
�|�5�����C�Q��(�J�Rr�t��[�I���aR���8����Oe��O*poh��h�-��qܽ�m�N�&�w��c��������L�^ַw"�"j�aVNaY�ATL3LU2Q�DMIUYPU����AFYe��5Q���DTUD@��eM��IDEae�eU0e�QU4ET�Q�ELe��DDD�FLDS1Ye6c�LU��f`MUYPffd9QD�8TS5c�QY�UEETD3Q54e�Y9TUPTنfc��fc��DU1DEQdQUQTT�QEY�UDQ�f5�e3Ycf`LEPHENI�T�fce�D�FTRL�e�T�EUAaQ�U55L�F&Y1$A5��SD�1�PLQD�AT�FcEeRD1Y�E6XDULdcT�dDTUQ�fXdd�UDLUUE36fFFUXMAEE�UUEnn�������>xf�D~\�����+�"��S�8��]��u�
�3M}Ff��ܛ��֭�n����N���7{����  y��ŒJ�:򿖡�~�������+3�k�D�YKA�2����)�}i����rJ��6o�ڿ =�+yuƅ��GS2#��ݑ���P͎c�2��b܏r�O���br/x{���~{4m�b�����W�VX9���K �3.��j1����*f��'��6��.g7��n}q�g�,ڦ|1t!�>8NT3k�$B�����M�4�:���]}ɝu,i����*����v��i:MW
O/٫}�yϥ���ԏ�IO�s^Y��0�s��9|։�����}���q�1JQax���4ng���������$C����H�jm[��g��ϧ�ȜPM.xV���}�su�؎�S=�x��Hu�Z��"�݂���DC�Q��v�K��՜����[�p	���u�p8�3�)�c)�/+��i�b���3%s@nPw����ncv�~��~ox��]j���KB�SJ��7-u�^'��MX���������j�<o�(�ͽ��ځ�9;΅s��<O��?6�#��<7ʙ��ۏα��­�H�uZ���pe�̫�E(����F�o���ڲgC9�ĩ3��el����x���]{O��e�uc6_����/�o�4��w�c�Z�-x>�+���?| � zq�x\��[=߁�g�|dW��gήɆE9I�ԙʻ��X�k�ݵ�V��W�Zۓǲ3K��>L��j����&a�����h�P�Ԍ=�I���Y��꾆�Qp|ϣ���ig��z��>�E����9E�Z>"]T9՗F.r��^yX����k�$q�^�P����*RK�E��t��tǜ}�,W��)��=y�w�g-+Tό�|mJ��o~��t�2�,>1�O�s�I�����:�<����W�O��靂�9�+9��q�
Va.4G�N^n�����dh�Uv xq�k�j�dT�G�"�s{M�+N�c���ǵ�~�Ie�6�:b�2+�`�v%9y�Wӱo>KDL����Oay�7@�z}�9��>���F���g*�V��OP��q́H8�-�ɤX���K��=���r�XcP��p��+�4��<��r���V!���sK�[��\>F�9�T�p��ϵC_4���j�8�>kL��;��\j)t��� ���m�{�V]��p�ƭh��A��͕ZB�1oX{�ܞX�؄��L�v�Or��>�^'M��a��I��;�o��{�6��	���T��껔�]�q.��ش*|P�Տ�9�u:h8R�eZt�-��7�0mw������%�A�5L�0���=Z)՟gԫ��rü��7��ե��gh���jf�%U��ww�S{��n���S��O�.�ܥ^=�R�9R���S#3i����j�v3$�{�yq߷sM���z4D9���G�ve!�00��U����)yz��1&}ޟ��Q{��{G�v������\��of[9�V����o:Z$��f��EN�O�i�y߰�^�H_;�SԞ�L�S]\>8��▲�7ß;�p�P��k�Y��܌M�J������E��OO�q�g�k3e7rǞ�3��g�&-�.����:��g��xa9��N��oi)�q"�k����XVt����BƭR�����������V/PJ�c�]�Ι�&���&K	��J��L�5����Ƒ\l��nʓ\ܯl�R�u������&}%���=u�M��OV}R��m�:l]y�����P�|q�2<��6����nw��Xy���d���^��GGz�(^�E\#w��LM{�Ȕ���tE,+K\{�n��{��Mb*���Rf�����6�_���kܦ��+w�Ǵ���Ϋ���m9uwvm-�Z�mV�[f��lM���{lDo`
��t�D�8����v��t(��+O]��9vCz*vO\���e+��o�����D��'�l�Z8��GE���z�:��[�n��,۔Ƚ�ɝ�5=�̡Չ1^Fgh�y���n]K�f��|^!�A���f��du����8p�%vw�ΪM�Y©U�8�ς�2���^Ԉ�e3	7��.����.yh�8�����c�A���"=��[�e����7�|�HZ
ևV�V��<�|�ڔ���ӵ�?	�HI�+�b�����]u�����v�*2��y���2�U��^�<Xf�탇�l��=�8Î�c3���GC�>��Zf�$�3�H�k�a��ּK�>m�����+v:J�{G�lMwF����`p�4�;E������@�hTI�
�!�#%��cS�a�5�B�S��J5ر�Cbf���g_�9c�9���yh47Z��d=u�h[�%�Z@���-2���Z����\��B�EE���۾јֳ�$M��8�@���G��\_�^�95��c���Z���?7�݊3Ѓ.�<�:Ϛr�k����x�o����<�y]y]d���ڳCgk����IKƯr�{��q��Y�C^X
�r
J��﮳z��)֕[���LK���'�v��x����ɳ���E��O_-�ܜ:ԲѝX+���~� �^m�U:�:ǚ�i��	V,_=�HN��\Jgׂ���l@�u����t�k�ۊu�}��õq1]�p:�Ī"�N��Klϑ�8�|<\��-�[y^eȓ̬��K���r?iC��z�a��Dc�(��K5��ڈ�KI�v�3�:2?Qk[ȷ�W�G���g(��hf�aX�L����^�>>�H�3A�fנ�X��1�]�82���V����f:v�>k�pX����P���z|��5Q�)��#7���c�����_Ҁ�+
V4��M�Qi�"8�dݑ�7�B�j����xlRw��R�o�O�S��S>;�V|9���B�Q������<�<﹡���V{WVs��ۛ��n����{vG��E�Tφ"�|�+%p3�����7�e' ��}G����puKs�:ߗxd�_o�=�\�+!�Uu��IV�A���=�.��~�J��,���kk�<�P���fx��|�|��s�J��W%��دU��������Ӈ[^5�vv�<��ޙ3���x%i�ڲ����S���T���[x�_(��й����'m�%�􌜐�/��U��dݤ��Y܍-��Č��iTƁu���[׶�uōu�tψ�E��9/�Oz��9���/�
�Lc�����{�߾ |��{]�ǅ;;��/�,UN+�z՞�övY���N5���x���0G�2���A�ݩ�.��׭���z�2�;���؅�]6���SU���EZj��_�����S����9�r��K��M.>N��T�y�8�T�-�.���g*�h���b�Ӌݣ�����b��Y~[�����m�%c�]�B��*%q����w���>ڼ�鞭OE�uC�$U��ϱ�a0�ZI����e'k7v��\�.�,|�;�Į�u���I�>Ě�i����U1I¬��]���V����'����>��VsP�7����T�j�;��֟'~U�']��wpr�^$�|l̺��^��e�X��]Y���B�H�������f{�P�I,�(/uS:�z�|+��v��>��ݮ>�\�h�ùCP/����T��h�v���6<���L۪�;n��5$y�Oy�u�$��yq��)���o�xt~����+��4�Q�yQ�d��=������w����߫hkwz���e�״$`"��F��.�=�OٙW��K��k�U݃�,c�����o����oC�}���,���}I�S�_,�4�[��ҁ���ע����#�g�έ�]�dk�u=_$�v�_W�}_s�;�c�:��˵6��#�݆�t�;폳�ׅ�G%o��1ת�e��B�z���tc�|V�����-;�o#�F���-s��t�'���e��#Ÿ�v���˩fc�F҃xP��4P�Wϕ
{�i��Ƴ�9C�*��n{�:�7�W���z��:�l�:�|��y,��	61ql����k���7^иg����>m4_g\K{G�g��X=�NٺZ���υ�it��˷��d�u��Qߦ޽�c��ͬ��U� |j=��q���1lTOOyfү�.��TL����r���W�$��ӲϦ����'="�`���;2��D>/��:�K�B�Y�-�ue�-�	{�gӮ�I�,���m̶s%iu�w:Z$�!���V����o[��F|ᡶ1����w����9C�Õ1m̶l��i}xha�LQz��	/s��0�RZ*�t+F)��m_ָ�J�rǞ��<p9Vtd�'�pKSj�|�N��o�7��S��jX��w*�+�9A��H� f�aؗ���X�#*�u;{�W�O����Kt���zz��+F���Y�h/M��#��������j���Lv�W2a��}�R��Ԟ���E�z#�có�=O���� ����>1">�F��墓��c,X�Qx�Z�J�}=���_�*�ar@r?��A�?{��D�z�����ۤ������ђ��K�\<%P�>��AfA��l��Su�Sx��AO���&��S$��D��:z�P�X��D�o���x�[��d8O���j-c�"�C�fǓ�
:�Xߢ��/l�E�~vb�u�(��T�M�[����v��z)Nl3*0X�r��@p޾������aÑaGFv?Y�eo��d��!��̽�WQ!�׀��6<��>���ek��f��^Gp�/c��L���#}�1�q����:�L�֝^�U�,^��a&�-=b������R��	��I�w�r��l�����.�3W�o����X��j��C5ԉ`�23�bްj���2��`ܞʬWOP߄�u�{����CXՍ>!�T6U0|o�HVP�+�wl]�*5r�Uwv'�N�OT.��|�v3�N5=տGC�>��l:f�8�#I!���ADԳĤU��i�䤂�Nm�]\�{9���V�~�rg$Vm0�.��J����)�|���󋹠��C�z����݊�Q��ч�N�b_$��Msܛ�t���]�ql\�j丹��J7bb��F����vTz�e�T_��c��� ����,zY�-:Կl�g��6&��bJ��\ӎ�fm��cK��Kx��ͱ�Ȥ�㤂4��:B�N����x�y�77�Y���{�,o�����deH]-�[��?j����0G�M`I��"�ƃ�=6�$=�X+��`u�x���,��]W�H}�S�t���z����`�ǳ�=��r�h���%%��_5�خ��������{ĺ3�꭛�]�˶z}�:��*r�X��t����|���[p��3���Iˍ���*��N�w�7=��^�uz��q�w��BX�DCn����و��ip��9��U�=�V�����]�����J�f8���Pr�a�/>�	�kդlK����Nxm��ƚ��WS�!7�����_� ��p�������^��6�GZ�UF�A��Y:GPV�׹,j6���uD]z\3��j��1�C�\K$�E���5*c�j��z�<��F8�_èb�+t��n�/jfDgՊǟ��Wr�1b���Kh��~_\��k�Y�9�W�YE��6�.cno�=z��cܛ�䅚_>{�����Nj�-���+�V��h�Nr�z�^>;k�����V��&��nǏ��E,Ht�0�r�l����[Mٔgg�-����6��p` �`�m�~� >$��w��ݺ���o���	)�ڰ�w���E����Q`����都�Ǭc��ݍ��қ�9�,F��u�ڸ�͑�g�f�3�����A�7Vxn�xY�Q�����N��y�-z��>�pÝR�u�.��p��ze����<7)-g|^g�Σ����q��CH�S�>K>��\�m�d9�峟O�=�9����Pљ����Yd�5�x�C`��_0k3=~5��u���_�Cجb�W�;,�..k�\~%a�Ow{/��}�o��M����X�~YI�x��Hu��:鵠�����k�@�Zhu�B/[�=M�;�����N�EM��lGM.tϐL�e3,eqm:�^�tǲZ1���4�B�b�/���7�{��`3B�X ���,$��/�KG��>�C
�2n�}�}}S�Y���O���{K�x�^��Ld���xO R{�t0D��<Ԩ�a���S����}��>�����8+�������F*φ&a����V���)��,�����Eߍ�������K��u�Y-wZ�8Y�V��|�[�ۨZ���0>�ݽ�z�ɃV�ڻ둃�H����
^gjJ��t���N�z8;�-�����f���@���씴��[���'���\�pd�%�[��+/�|��kBeW_L�Iy�d�����{If�a돂hZ%�p��n��3�m�]�U�ׂ$�h�T��I�
6*�ecR�f0jwW�{��{��a�����/��}\���H9}�X�s^�_x�|cncd"��hr��<C^���dI�ӛCF�d$�[x$5��g.��8�n��
�,v��W�(eX��:�P|����U3n^��f��H3�s�*1�4�a�Pc����m�P�'&x�ܓ�ތ\=�4sų��gާ/]uЮK	��[��&�ws7UN��v�0v�Ւ@SBk�1=��6�������2��h�!u��Ϋ�4_֗c��#�
���a�3�m6�Y+���|;e�ӱ��V��וS��	wӜ۰9�R��-z̗ʬ�j���9��ysٝ9����{�Q��Ĳ޻C ��S����Un�-�)gu�;M�|X$�ɹ|.�B�]c��ʝU���x��딠���z�ׇI�C�6c��w���~۝֕&�,V������]��w��̱Z�^:v<��t�+�w�K�V�����|Dv����b����}�{��Q�wQ4i>���/�HЍ��v6��'�IPy��F�j��7�簾�U�.���W����دx��mͽ�7˄�+�]�z�W���j��8����b��7�=�1��0�#�pl�,�o㝔��p��X�ڴ.s��v��O�Ю��<�3��`ZH�o5ց��e� q���hY'A���ჩ)9��fc)��p�	���4p�)WP,��U޳[�%�j;}�*TW����q�{wy��r����!�G�[�S���ŤuwJλ2�^#�T�A��=[�!��K�`�e󶶄�Q��^U9y	T�/���aYG\����@#�x�Y�Ôá˥,(���yլ*��u{+�V<�u��>�^��s�n�N�fnɃ�n�d���&[��L%�]n����>a�3�}ԭr"��v�������Vhe_P���������˶��SQ��s���TbB.j�CtwX9FL�=G\�UBq���^�s����Y�j�s��㛳N�Ս+±k�[�˂�,]t�kfQ���̉�ˈ�&��Ez�%��^P������X�8��ti1�{k�c�7/�/�X�<��]p�3���h�lf�Y���ݎx�v��[\�u*�ӈ������G���47�x�r��w@�y�:f�{$�/v������fݦm�tifK�[kS��Y��7�M>�������P�h5�E/)���!��""� �1'0�(*"�r2����"��(��(h�b#$�"��"b(��(&b�� �"�J��b���
�)� ��"�"*�# �f�)�����)�
�����+0��ʪ�������("�3�&"�*�J�&�����(�(�*�"&���������1ʊ(H���32f�)
������b�ʘ����$�� ��*��(��(�γ)��i��:"���
�*����z�Ȫ&�(�*)*����������+
"�bl�(�ȲɈ�"�"&�j"�*b������*��1*
�jbh��+�ʦ"���&*J*��bbJ�h
h�"���rd����*��
j��#����
��j
b
��1	�� ������&���i�@$�~$��'�����[��E��}�f�"NcC;]�\�J���ݮ��~�b���L�
y���.���on�E�V����U}_}BD祓�ЕuM"�m��C�[c�mE*�����Ϊ�׆Ih���}��PN^+���<Y�h�b���P����GG��2S��T8��c�½��*t��2���s^5�+-)�G�L���5�j�P��;v�4K��eY��g�={���j,~�c%G��#�Sҽx����X�W����V�"�I�#)F��OgaMe"�<���Cr�7<'�+���/�e$;���������^���r��´�mi�� ���ڄ��+��W�c��)����,9��a����ׅ��t��폫��R=�P�p�&p��VJ�1+��(U�����*����	ˍa���}r��/3�2zm�tz��a��싦V�lco��#�Χ����Ų������s�V�Ӟt^[�L.5�<�v��
�+��쮽���Z�Ȋ��Oι��$;�]f����9�4{ٝ�#����7z��f����Vt��k��@mD�����ᔼ��:�k��Zy�:>śl	9�u��c��;v����N/J����%�`C����AW݌=���NΤ��B���l�t��z���c��b\N���-[cq�:��Bp��\�ML�XG�����\�4���&�*&s8�����K���}�ʯ�}����3m7�nw7D_�S.o���'=��>������Y����������:*\G��=t�.�bT�V-�yq������9圙�扖�`��q�zl��H��n�S�:�)��y�]�9�퐇�iC`�[�1C�����P��L[{7Áދ���gL�7��B�~��_^�)� I22��D>��ث^[V5q���P�����>r��4)T.��_~^��6.���m�Vz$x�R��I�o�+:z�ʉа1b�`;aUI�v���Ws�8�G�ݷo��:$h6�i����5��K�Q�]f|��d�.��.υ���/�Kqo]��z�M��v~�&Â�&�J'l6�tڬBp�z��μp�uZzW���.�w���3F�dx�[�����0C��^���(l�k,��׸Y�2x��D7�皚D��t���\#o=�!Ҍ��鿻��X����iӱiD���2�S:=�$��Խ�0NV���9�|M^b����z���1�A���������=����������Ä�����x�d!f�k�Z][(VS�W=��x�w<YS=��������.��#)�a�8����|Eb��9@i���W�5��ep��F�%�h��1y�<���8F�Q����W����ՉM�|�0�8�X�;5uުc+�s|�^�> �N����-��\lXw�X��C�1`9ʮ��x�k�Ύ;��I�(U�v)mat�6�f����4:-k��;����,�bFZ瀺�h*z��S����<�S[f�=�a��� ��hk�(I�V��=췺�k���#�J�����L�Y�˓2�.�x�,�t�!peC,Ia�}�7�ri���uҼQ�Ι�|�#kr�k���x��)_t~���a���V2W��0�κ7%��t5��'Z<lG�c�1w���h(����S��V�р�,�3����N�1p�o���	�U�,v)}-�p��o�gv�����f	�h��D�ڝ*<)=
��k=i�5��X�z}�|pA��:{�W�������rμ�Ly�b;;��ec�ZX*S>�U^P%�`+W���UL�`�=�+fN�2T����{~�%��*J�b��I���*W~��q3�=pI;;'���/9���R�J^h3���_1]�s�BX�lW��d:u�e#�q�<6�M��4-��ɝP���sRU�H�Q�v�~*.=��$�ry��`�m���d.�k�⨘��B~���y�G��|��a��3�j߰1�+��j��UwV��k��	�Rՙ��X�ӫٝ�!0��ɻ~3fju���^�־�o|xU�����|�<7L��m�G/������A,�⣟�����>��a�IZ�vt/�����W}�����KQ����,�ER��S8XOe�D�Ӌ���Y�W���i��n��Oe>qqy�_���~?_��fǮ'Y�������ڀ��"�8,nuD�����+���nz��G�a۞ۢ�;�Qx�)X�Ϯ������dG�L�)Ԫ���ډ�j����B��Iz�IOT>Յ��>�}A
�G�3
@���kd�T{�y���z��ݗ�}�˰)�û������zP��#�π�6��E�]@���`�>��W��=�"^�}�J�/;�,W\0�,�u��z\=�<��.U��D�bmߓ�^��^E1B���Z�.Y�� ��'-��5�{�}×�*�OW�د�&�ݏG�s��"Em��᰸wK�o���'��Վ�^/p�ܛz7�D���Ƈ[���	N�^�}I�c�yT;oòyb��W��Գa�,�
���"�P�e�rNq��uy�V��R�/E���%�+Uo�3yl!���]�E�曇\�ea2x���P�%�ϠqN�IԺ�j��L�un���wgT 3����b��5�U�e��8�-�ogr?����56OL��۹��{-��:"�$G�ۺ㦗Zg}�
fX�f_�\F���蚚�u;ɷ��O���W5����x��v��w� "���R�-��w?e�O<I���CpՂ<�g�P��Zl{�����{K�x�2+�Q3��;�&|I{/i
�֞�u��0%����v+�����M_�S"�j���S��U_��{I�^Wɘ�4r��e{ms+NcE1�4e�*�n�������V%V;k竁��:��ѓT�2����3ܶ����xNV��5L:2�h�%:�����Ȓ�=N���TƳ�vot��n��U�u��Q���Q��`����8���U�/���?�m�:��w{%m���Շ����c]�H�2�}:�r��>��Ց����"�g��35c/�<�կ�%��G��+L���0���݆�t�;��}�3T��!~G�mu��y?f|��k+V{��ȽI�
d�	B�����k�6/�0�cӮ��㘺:f͑Le;��J�<-Y�`������w��=�	��}C9b�X]5ǭ��e�T*9R���hc+��A��K�)�@������<-�k~~�{HgV��7�n�}��>���v�(�� �{ي@���s��Ṗ;/l?�����T�0�]ߟ}FK�o��d�|���^�Ξ�i�V2
�0tbf+���^��'Ҧ�j)l�n�aӗ��W��&[���ۖ7���n-L�u<�z| �e�X4��>��W`��j���)!��>���
���p��3 Y2��ZeJ'��NH�Ρؚև���c���=�4����7�tf�ڜP����Cn���ϒ|����˩i�~+0z�/��G��\ٺJ}�P����6p<��lD�u�w��d��XD6|���,�rϩ����k�i���S=��!����93�!�t�Ņ{;���t��o66b���D�Gm�Cܬg�y`R��ߝ\>8��>*bۙlٰ����[������Ù���j��%�_3��c+���\c��3��x3z;)vU�O���f��v�K�p��V�%`�H�Myh��.�5�㊝�����G^�]�ve1rvf���Up0ID��җv#9T�/����J��˶Eb�Lںr7S�x��N�&��j;`�i����.u�kiL0m��'�=hh�y�u��/x�t�+��ᯐW��ZxMܲ�X��I��wU�̣wxˤ�ϡ�e���W����7Fۮ/�-�ؽ��S�)Y�j�[�/��Z[W�����4wR=J�wT�
tw��J�t:���H��|k�uh���L�}(�s*��k�Z�'����3���WF-��^��]s��B3V=g��`�����<O���-�Hc'���?	�vԕ�nr�|�/ҺC/w=��c:�,���1e����8u�D�FX�����n$���6�1rz��c}�g5O����t�𘗨e���T��|M5A�x�
�S��ix��3�݃Xy�=��Y���U��uq���ʷ/��O�J���gG+�l��镱�E��b�܂�?_�l��ML����˂�������9)s�\]AS��8΄o[3��'R�4��<�X'��W3���o\�Lyu����#ë9x3�:M�*�۬Ǿ���07�\w�k=�h!���V6T1`ۆX��Z�l�������.���L�{��s{Db�k�ܚy�q>H�j��ؘ*_%�C7�p�s_e�昜k�z#�YM{7c�yu���v&��`+R�Ag���au!�R�V|��5h��no<�/���5�q���7+������l��z�op�g@��w�|�>t���e��w��g���x���]R�}.Lh��k��5��Cjfz���^��3}C@�v�=�e��T��O�7qMFPP��@i���(Bw�ӛ�^M`wklj��E���Q���k9��.o*p�y��j�@����ϊ�� Y/�!�i1���j��9�6�מ�gw4�k̻<`�S{B��r�4Xy;�@㔋K�W��_ޠOPM,<��/Μ�����s<kΠۭ/p��ϥ	i��r��� 粒�t6�ϪS>�p�[�kP	���)3��I���Rpbj�٪�k��lM�O����b�%W-Fŏ�Co�{fԖ*���ՙ\���۪��7=l��R"��J�rEG>=ja���W�����c�|�]?����y�q����6)����a�.'�G_��Y��&�C"	&=�,'��:�ŭ���>�b�dU��=u"�<���4� v���*�Yk�_������XER~���4����P�j󓸤��k94��ƙ��o���j��?�����4-��9i���ڪt���n�}��.9�tRΖ+�/?��p?pP;~U֬�Hf��_mƪ����g/Qq�l��8�S�k�������h{'o��}��_{�T��@�c���*�Y]Be����W<���n]��'G'�SP����o�uˡ�R��ӹ�z��Z���y�zeѸ�+5��]�u���e���W�+��r�f#ajs=\4�8���T���@	�
�nS}Y^"�z�v��J��=��e֋�m��k��+���,��N��Xږ0��q�c����<�2x](75�ۯ
��kWZ��ٓD*]!PW�j%�������.uC�9o�q_f9ܟ���4�-ߥ�:���Ll>{�D��>9ix<3�F��t�h.�o� i���v�#[��uj�v�8��Z��ơ�8��fT\�"�0��\=6:|�l4�-���EǵT��*@{c�G�_o�\����!�+�Du�=�@ܕ`�ϳ�̿�������*�G��f:6�o�H�3�1{]�3%sB�OI�reu��w��B���|�zr��]���X�M�צNf�b�p?���/�O�>���{�B�.7���4���E���wPq��ۡɹ�/����r�������r8��e���o�]Ƴ�¬��_u��n��=x����&�4���m��ƣ<5�̕�|um�V$�ݫ·Ǯ�>��h�~yY��n�|�k�p�4�i�ު����kG�I��U��+�D��M�~cE���o�b!�L��ثe*�I$��N�ѥ�ws��Ƅ�i��Gw���*ޙh�i���
����V���hm�{��PZ�r��rd����c��Xѐ��k�}�SL��d�^�����r�%��}j�Z
�b\%��+w��Z�[W�Wp�ז���esǾѡ~��%�,�G�×"��6}�2���J�EN߇AѲ5W�bHo�p���n1o��vyo��>{<J�w	"���V	Ԛs�b�G�cl�U�6�{�e��Ʃf�	��1�"�{?mq���,�ޫ?�������d�>�,6�&^�}���q�xZy�e9k՛,��l����<�u��B|F���qk�Zÿr�%`dw��n���V�3���gT�����Ǖ���ڱpOY�[��O���P�A�g�}�s�e���n�ʾ>�������?-��/f<g�eM�.l�>��^]R�V2Y7�w�\[+>��N��^���*o��B��峍3���݆m�4����\f\�^(� �^|��˗Y�:���n�jb��7ϊz�eLu����x:丞�i����z��BˉvS��Y�e�=_-XM��S*����6p<��BO>��>�N̠E�`��RC�a�/<�s~^�(t��-3�T����c����uٟL��sD�g0J�F���@kط<}ŃuNZ'X+0��v�2�osz��[մ�mlFң�GNm�*��w���o� ݔgI�}�K�Ϻ���e��ѕ��9���?	a��{�RnnM�n�'n�b�;L�\�<��]�+���.��B;��	bv�ҟ3����6���>��
��%J*�v��'�����_b�"�݇��w�p�,����T�M7w��Ň��3���mlʛ��6E⳽��1o��_Z�!��M���ʹ�.7[g��� �$|' ��n=	檆����/�=�o+9lt+�m�~��g�Ŭ��������������	�#ۏ��b�]	�񖡊jT��-刪�u�v���{8X�A\�%!�T�X�6M���
�����Y�L�]4J����+����~c^MO&��4D�;�.X��7q{w���k�9�s��OtYE���)QԺ��6��p}������=5u�{�����	�nTe��u����2@�i��Ő��$H�nk��kq�+(��jx�6Kv6�n&b�[X�^I��*�2����4��A:	�)��o�%���:�.>|&z"�Kn��[�K�J��o�3��Rp��/F	YUu̡Y�m�V%��y�,U����w����������R���l�d�L�ꭐ.S�}�f����n8E��y�wg:���]�Y�脾v�qJ���f�_P-X��9� �2_k�U����ɫ��W���<#{ל��a��z��n\��#�#6�Qy�4�zz���+.S��֒��c�$�7�8��5������7-B� גs�^ݐ��n����W'l�yB���|*����J��
�
�Nu��U���\ic��F]8k�w{�N*�'WX� �uwDR����\V�K���X�,2y���g�!�F��7�θ�d���os/��l����N�t�.��8#��>����nnl�
HJ��\w�G��J34�LM4���o�V�ݗU��܉�u��>��w��p�!To�
�I�I�QVVǸ�Ⲷj"7��'�jWh:�=r��Bf�+GI�[����>���b;��LV��;�����뚵��2�oަ��qX8�r�ڛ�b��Jqnjo(�L_i^��mR�5�uR|�wV�h��'6�K{��2�Mb�)�]h��鬏2��fl��Z�Ӑ��<���6�����u7vW��qY���qUEٮ�o�&��m�g��z��BM���w�1�	���s27z;Z�6����|�KE�s��#.5��*}�a��6�-\�0�f.�ҋ4��Ue)��.��J\R�e�C�s�8�s�v�8]N���c��B�>\4�kU����K��c[N"�����mɸ�<}g�͢��.�.
��v�E}�Lw�=Q5�����F�dݢ���aOUl��2�3kWY{x]]��'����5�k�5�yb����V4iȻ;�(^����y~�מh��)��jj�������"�"
&H��
j�FIUDRMS�`D�RCSPIM4Q�TLQ-5DQD�TT�D����u�4��TLI5AQTUu�PU2�A5QU-PDQՙLAUS1UQDSTIfaE%EEQ1T�M1UDTE!T�0A���DT�15ET�eQHEDQ�c0�EATUP�34�4��D�DD�MS�dE�531EDTU$�33d�4U1S�E3WS�SU)0��MU,Q&c��TAPAT�ET�UPE�`e4E$QUM1SQVa��U%MLD�PTd�4AASEEMD��1TME1DPنE%3DT��zV�;/�����Ԛ�Y6I��0Q5���]���G�����Shs��7��32���:���/3��H{8e�]���]��d �h�t���q��j�
S;������*/h;}���<����̩���q�I}~�������gI�p�G�u<s�K�x��޹a�W� 摎����]M��F{ݷ����/
�&��\1eRZD��ז�D�ˢōqx��s��S��J�o�=��A�qp˸�Q#�$��30Fr�({��=YR���]�%�j�Һu#�~S�y=_���� ���Ρqa�L����x&��u�E}Y�=���8pk����{��|���fP��e�a·z�(���0�i~K�=�=���{1�z[�z�����?,k�6��J�ڸF��fpj�Lj���}q(򸴙��2�ҥ�^�]	���甇w����Õ��j�(^�U�X��#��r�������)o�o�xNNk����v����O�oN	�U��]li�(ŀ��?S����w3mUp�Õ�B����o� ����}=5cC�ֳ�Izv�/��\A�g;e�:�˼�;�Ai*�}��k-�<�Ow\+c��N����Ŗ�ML�kj�o�q�;%s�Ƀ{l˅�'c��?�%�#=9o���"�u"Ā	��i�F�����؝[X��y�'�U�_d�P�4/�շaj<vF��z�h�j�+��=�%��sw�h���K��K��=��9��G�<�:�/�8�����'��WNֻo*�RiWS���=�=r�́��W���6�%�0�:�bq��Z#�ze�a�I�)W�;��dJͰIdz��]˱��%�C7i�g�k쳒P��ƹ��q��z����s�����}��¹.Fʇ��C��ԇX�}�|��Eo<�n]o��Vѯ,5��=�W���~�u���/D�:3A��<G�*k�P\E�C�2�.;��c��ض�d��s�+����ܽ�L+�г�\�Ł�};�@���ϪW��������(��ɻ���Y��N�;�\�=��BZ�8.T"��b�sn�Ά�J&vŗ��>rJ�������S�SK��Fjֶ��P��W��*�� �C�vD8�Q�V2�	�X�Ԗ�N�ɏ�4�(�^�Y�u�H�r	o�EG@;j}sGӭ[�\�E:��N/_�ԝ����<F���6ԪG��+g���<,e�Y~T �+�h9��[�Ks�ί,��{|� W�G�t��)a�n�L�?O.m�{ݳX�kݤy�C@<%Y���b�Ɠ����R��t�I����f��jSp�3�Q���)H���^���!e�񏶸Y�2�����w/E`�>��f�b��k�zp���Q��q�~~D��)_��2�~ �;��\r�����>!�v�BL~�z�B騽����no�]D��|�o��>wM_��1�
Vjyt�~��'��
K�l_m��sm���7:f]���]��}^�N�����{j�0���1}]�:�66�}3<���>�VX9���S2�9�w~�c�Q^����>�r{�ӷe�+�d�Ε2<�Ӻ �be�u��y��3zٖ;��=(a��'r��w&�;(3K��g�0{�_���q�u��J�b��G�D��Me3.uC�;��%Զ������w�<�;߳�ޜ��p�)E��T6׾U�RDn}T��#�z�Si}V�jJ�w_�pg����Ϗ�sS��wӍi�nTXK#�*���1%�˒�V�GB�kG}+����z�<���T2����:��]@'R#�{2��%D�&&w�)�~�Ĩu�����u��������V�W��i���w�\УS�f���ņhA��`�*�����\G}l��SG����9���Ņ���IAM&��n�z����'�zNf�Og�3��9�KI�-\x���4�L��\��:�p*5��:ۺ����f;)����$�(/�<x�;�,y4mɽT��e��(n�&�7��̺{�����Ji���|��7���򥣟�q<s��x)_g�u[;��><��^d�s�Lo?9��T/�d�J�?U�ݕL�#�k��ڝ��MV2�Ǻ�N&p�uT:{~/.r� �>	Lv�j�]t�ƍpeI/����`u�ѾP�Ք��jU3�_�s%u�[W�X�uڼ+S��}�������ywm�h3�tb�~DXʡ�ׄ�m�CP�2�5�_��;�^;���\s-���Jwp���K��-jY/'2�j���1r�\�\'	@����kkc��y%zn�>���ʷ'�W��$_�e�+�M_�f�W���MY��q��	��8�e[��ڙ�Xlp#��i��uf �������}��ϺV����(�Q5~rU?Q=��I�WKl�b����V�7Ղ�2(^ݰp������jZ��K�:�:̒��@����ʊ��2���N�9�]`��<�é<��}}A��Z���j��c:�^l��Y�{DF��RE��\��揧��z8.�����-L�yp3����Gl���������~;ܶ��¹&�
���㺻�[�+d�XR@�[
�&�i('�6���Y��2��H���7_�@�
��ݤ3��{�v�v���_X8D#�G9?�S���/EV_���m�}��C�ő����z�8�湏_��c�z��w}���-���ˍd�\_,2&_����G����V�G�fI7�R��;���[x�v�RF>��xb�_d�
��5=ձ�yS�êi0p$�{�t����x,���e��s:"�ĺ�.#si�`=�q��'=���n�w��d�r���5�f���C��n�y��bX�0$��
쮥�S՟)L��ϲ���̿K��-�)mk�5]�M��}��,�Y�`�։6D=����c:�)��<��f���w����̽�Yn����1��
���I.#Ը�.��������'���Y~|�rZu���1�fr�&0\�����Jˤ�Ď��dV��.՜:��u\H��]o��ǔ����]Xjg���|�4�J�Y�L�Zˤ�<y(��~�:�-{A�f��2ȳ\�ú��ޤUא�}�."\	�|J'o�6�Mk�Z���eE���3�y���b��˅��7�aȫ��W�Bʬw��z��0��$�Y"��ݎ�ǵ����7*�d|I������2����e��7�g�]cz{E��/<��8Ȗ�m���W-��ޚ�l`�0�;�xh��ո$g�-|��s��v������s���K��!Iu>=�A˕�8Rf��b��R��-6Ro���Y~��3^�3 /}�p���`g5m�3�_�Oy�J#���[�I��}�x�W���V�_�Z63���Σ�Z���Z����28_�(��vg�����b�d���8x���� ty�^
o¦��n��8�[��u\F��N��"�vq�Nٹ��0L���n��d��]���_�o���\G�h^�����]أ�a�NUc����p9�M{>�ܔ��[���'6��S�C������}]��rn�W��Y�N�Z�)P��h,�&�N��]����%jo���λ+�B2�
ǰ��#�S�:ś�c�VhF�G��TS�KZ�o\0�}vzJ���CB����gV��N��Ӱ\/mS0��#eC��C��ԇ)]����s�z�]H����,���Ɗ�S=���\^';���L���Zh�ԁf���\�g�,	%����������L̕�x�]2���]��,<��q�E��)�`�P��h�7������bkxn�;�XJ�\�+�fqȡ��f�!33��]-�,�B�PP��X<)�u����}<U�]��	�Y�RW��n�������Z�eЫܾS��X����o�X)L�5m"��Y)X[�ImM�A"Ei�Jꨯ�X{�/��]#\�׫q.����u�As4�BR�x\�Eʱa��I�����5Ҷ������sj�N�z�גg�ջ+iL�uz�uqi߹��#��>�wdB+س0��>���g[ʶ���7<��Q�������s}H�kMWmȨ�]��?"Oz®s���^�w���[�v�ᤖk<5�)<U���D��? ��+�@+�hk�K���:aq��>����|�1~D�׈�~w2�f�\Oh�E�M�<v�7)���Ͻ��Ҽ��R�o�N�"=�a[��K�JqjX4͇3}GϞ�k�T��{�xM"C���3}�F�v��P�#�a��vF{]�P����rV���S>q�ڳ�,"ҳ����u��/-Kկ{��}��&8��3/�s0�JP{�긴��$�f�<yu�k5�їKcު���Uq���yH@B�L�LŞ�bu-BzP��;�LY�sm~��g��_W��B�;3��UǙ4CU�*]oՌP��V.i��m�l���{�A�*���C#H�j¼�-W�w�i���d�[���o�����1�ir������Uf�!��U�o'��Ʋs��3�p��/iܱ�9�p����g�<�]��e�S�F����o�k�bۮ���[�>J��9���<�A���Wwa���/�'��N��C��}o�S�?	��|r��xbK��HV��At+|9nԹ�lָ<���d]8�蹬�q���Z{ܨ�Դ`ϊ��$�����cެ��l=ޣw��WFB�'�*{k@"O=�/˜��9�NH�麟(I��)L�>�W�����U$���v�����)]���lȹ�Gn91�9��Bx!�%�Q���㽑�Gz�{V��´ג�R֚�1�䡱5f���d�S�{c���C�.�~\��b�zly�������0E��W:֕�JjwT;S�jrM7)�}�P���S˫^���z���������,Eǎ?���Q��[f#��7>���,�/e<���K�����ud��#��p�J-xIH���̺�m�S �@����h��L��,Bk6���bnwy?S0����BåX���#��B��6}�2�\����]��:���[=n�K��⨼5׊�9��u	!���V:��f�W�?SVRB�PHZT�C��h�#�]Wg�����9���#��卙��ܖ�Q:%�m�S�}��4�Iڬ����W�n?C̞3z8^L�2�u�u�®�J�l{�D�o����o�v�R��g���:}��Y���Cnmv접�ł��ѫg����T�Ve���:�v7a��t�;�V�k�{��)Z��q����F>{^�%�����T/n�9����-a`r�%�����\#�f���ԩ�a����'_���x'��ڭ>J��(P����Z�K�k�`өBRޱK�WS���y�Ou=P�/�.�<�=5ݟO����ϪS*�Y4�BL͆W��|w�y��V����F�Pb�WJ4;��\k&���g�Dˮ�Ŏ�_R昮�;�J��}X�<\ �'��rzK9�é�w�9�#��ڙv��4��C>�5=բ3C�LBuM&{�����Ȳ���ڲR�.���JiX�L�϶�v�&�'�=�ux���W�3F獨�������?Q�Di	/�m
//�3��=X�3ۡ�C���rg�C���w�WL��mlr{�==�(��f���t�I���P��h;ι�Jg{~up�����zG�-��^�8z�ہ�+�ޯg�܇K�l����Z�db7B�b���Zqy;3��Uu��S]2�SԬ� -[4��˚K|��eּٔ��gw�ց���4��=��ͻʟCK��5�.�=�ԟ��i?.�����z�M�b��0�s}����ñ����@���� �4��[.�{�.ˣ�}d����z�N��fʘ�6��K��%y[D��$i.���M.�^�-�4�6�T�sݸ}:ůc��;%�=}�������J�X*f`��RP�Ɋz����˴����^VWI{�v�ޑX�W;���C6d5�B�&��7҉�soެXƲ�,�[^5պXk+h�'��ip��Z=R���>
���(���i\G+w_MJ�?N�$O���G>���~.��g�B��W��]f���
>�U�``��.�z]��t��{�ԧ�]ë����Xμ�9����(��WN/1�P�guMY�F�پs�2��-Ⱥ]H=S��h?h��� g��>
f����[q3�,�c��Z�>��a�w1AQ��>�U��ǉ>,�{V=������sX��qo2�D�V�Pzf.՘����묳o��*�`�ʍ�k�ϽL�o?ώ�GC>��6U�;������w����[���h�t��J�����u���1g�p�(q�����_N9�%\%���1[v�BS}����2˔���}�רx�m�K6��(SXB��-vb�����%p�����8���2���uW9��:<�%;�L��t����q��=D����P5������l����2�g��zv��&��>�� K!�51^��H��"�\�;rB�)�/�|oV�Ř���A�y�l��JG5R��K;�C�ڃ�(!�Nn�`�7�QO��i�\޽T��>W2��n*��b����63E.UV3Ӯ���˚Wn3�W[{�QtK�+�+^��N�q+�u7��s��1�7=e׶��x�#�{��關�t4ݧ��g�7�����qg��{0�{J"c�K���g�-+��)����@�b�!i@�_.�N��+�v�m�R��K�+��沍 3z㏶�	(�,g2�m�zzk��v(TStʣԻòH����qX$����%{ٺG.Bq��+���RN��ViPVЉ{�El�F]�u�7�lD*�G�ieu����Wr��Ad4,tw��&؈ng��j�q�X7v7�x�����HZ��ɻFJ��3V+�S��8���q�o ��5tk5�k�̾���;��G7�ӓpJ3̞�h��5��{SͷŖ���8�מ��.�hnh��{oݦ�{����x�SAt I�n���o^��a�i1ACIMb��΄ZN���E�#M�+x�c��N�[ݫ��#O��#c&&l���fݦN�m������۹����p�y�j9�ݞ ޺���w�Y�ͥ��#�0]��h��E~eɃ� �َ�S����H
���Kהe������ǳ;{8�^�i�?V��&XT�u���]�ٷ�yP���n��%�՛�mؓ3�W��Q��4h�¦\Y˄���8���W�b��v�S�V�O
�R��Z���ͱ�;��z��dGP�i/{�Rd���ᗝཞ�+�O�>'%=����q<�TJ�-h�p뮺�Z�T�wK`�T�ҽ��P�^k�H�U�+�a�7/�P�ۣ��Og�[^RYh\�r����h${�Y�&����6�x0gc���z�2�/�Z+Ua�Q�3���iB�}�BM0p�5��^ 퓤�����E�{���Q.�+;��F��~2J[�BoQ��]�r��!����}B�%%Ϋ"m큜�Kn�n�g,�.[�
ٹ�%�ع҅U�dl��h��D��;�M��e�me��K2d�q#y�B��E禭�-��۞S���$j�w��Z��z������� �����|`W�����X�p<K���P��on��Y�-6��-/�H�ge�U�_�\ҽlz���n]x-��w-�4��c�v�1�a�U`*���(�����a��\=彑5-���cU~����|\w�q]�c��V|EïD�v�_��x���yRGy�G%l����l�ʞ1 �?�$�f�&"��31�,��f(� ʨ�j(���*���'0²0*�	�
�*�"���	�
�(&*��j��Jl��ɡ�*�)�&J��)�Ʃ�$�(ʨ ��h2ʪ�X���"�(��0�
hj��&���*��$&X�((�
*���������
���(���Z
\�*��ʈfH�JrȠ���*����
)��*	���*��X������i�"
"�(��3
"b�"��
Jh(���i)"H���������� ���(�����"��f��$��ȥ�H��"�( ��i��Zi���(h(h�������ڜ���{\3��xKĒ����}�b�n���'��n��7��=w��(�V�a����=��N닝9�&M��M�8�ۇ0ط�W�׽GL�$�5�\��S�Jƺ�{}p�7���/��};3~�L|��C��yK�ӎ�fm�f��o��h!��]HM�=�A���v��-�=�l�u�}��~ygξ"����l�V�|=2�9%&�0��A2/��ޯr����oC|�*����&���\׎\��B΁r�4Xy;�@����ʔϩ'�>�&����s�*��S���-!��^�������P��\�E�WN�W{"&�6wU�2u�s��X�N��v�j�L��@�u���YuqmΡ�\����r�jNޅ<nz��f��V#B}$6���k�>p�cs�o�_{�U�~�Q��P��\ed}i��p7܌�m��W��<��#������/�u�h�}f�l�^� MY�r�s͞�JM{���13���>>�wGL�4� �^�ͪ,�}���S
��E���Ƕ^A]�:ߖ�(c����hS�R��3a��Q�ϝ�W��Lh�(S�ڹ�	Z1k��Y��_�o�ҶE��u܇Z��N�RT[�]8nt�:!�iSDV���i�)Y�ƀ�s����fu6��K�
|�"�e݁���]�x��v���U9��b󥸊i3p��;s�w[���Έ<������xd�%�a�:���B�L�ڑ=S�Y��|㽵gs�ݧ��w������]�2��k9Q��c�̺s0#~^���ϱ܇XR��Gg�}�Tk����i�rΪg	uA��W�T��>ަb�[1:���],iX3�:W3�Oi]����=�}?j4���/aWd��C��LW�j%�4��a��o�2����Ⱥ��9���&����w��ŗ��mT6ׅUq�������(m)d�^�l��[�ūzݤ�Z�j�Og]���'�t�8֞Ϝܨ�:��
��$���{�u��x��<��ǥ��pU�\�e��ݢ�<�ΰ�C�V	Ԉ�̠lIQ&���}wާ��˧.ӳ���)�iqt']��T�J���7�&S���~6VP��.9���l���B�A8�`��~ts���Q��4=�~�|sp�t���M�9eoM�����X�Us��lOy��o~n�K���r8s��'���49M�B��D�S�^�z�乺ŭo�+��	�b+Yⴒk^j��A�z�@k����m������N�������������;�Q���wG�J̣�w���_�/e~��)���8E��Q}W�
.�=ii�u�N������a���fu�Η��j�=~���n�s�Z��(GjFۯi���`y�Q/�}���ؽv�����-Q���]:uL��0Ih�ٙu:ۤ��H��}�r��>���&Y��=mc��2��Á�IV8,+ޱ��yb^�u&7��',�V�Avțs���E�x�އ+9��������a�۵q`�^*��J~�Iev��t�zgX���Zv�q�w�:_4��w���+0�u�
V�8)C�e���Y�׌-��7�O#P�R���2ߗEV{-�;~�'����u�=��9^��Q��N�R�m���T���k&��v�4؄)�윜�e�3z�>�x[R:gF�����V%��\u��֢ ���ͤ�n���>�|����O�ML������=����m����^\�y�v{nVGo�������v��>���Zy�^���`�k��/�_X�}^���1]�p�R�y^�'T�;$�k@�9ȕ{�vObm#�t�,����ABs�<T�WFhy�LB�qP��[�poj��v�~;¼hW1c�li˭����C!�S��-Pƥ$��ofRܡ�̑�s��$��K:G�u�x����H�r�wۼ�tT7��sH�9}tℶ��9ԁU�A�����|8?:����BN])|�	77��q�����^�T>I��+�𺖙�R�W��dnm2�����Nz4DO7N�}���:��{v ^r5�{G`�̠D,��O��(s����T���{t>�~�����^��Ut���//M���c�=U�蒹X#C^':R$��m����y�<�{:�S|ǫ��t�?/Oe����<`|�qS�b���^�g҉�/e�K�UqJ���ڦ�P�w�v�K����mO�C<�e�{���1xT�5p���τ��J���\E2��:������V�\���.�Z����j����|�4T�R��|��(F��Xu��{Sܻw�+���o VxT��>�D/��O�U?A\I�����	������^��n��q�5���g�˅��aȫ���Bʯ�;�Q�5��Fu��粻.��>c�fُ��7�M�H��~}���]�ġ{�p���`gNRc�hlN�Ӣ�n}���L���r��s|4ߝX���A��#W���	���i�^�^��W�3�IG�aUz��Z~3ޟ���cK�h$�3�~�,���O2f5Ȳ �ګpK��2\Uk��=J�5������.�Y���zN�ww랔��pt,h�:� ��W�d��[�u���+ݭ	�3�l���{�U���v��g.�wD+���%p���:�@gA.�{�`ޞ&�(��wr����E��s҇R�{g�7��U5�ٜ;p��L^���ٰY�L�&�-=b���0v�MY�C��Je��e٫���1�5;G��*����W�u� �~*�W@_S��jD��E|���a���d޹�����A��U�u��ف�<�ޮxDY���:N�Pr����D�k�bچt�8Á9����gǡ��yҩ3q���N�̻63l	26�#�X�v;)�%k�c��
�n+	荒����$�v�z{n�f��|'�t�.{ÅrZ�0���z�[HmԽ�NY�Vl��y����^ݾG��n�׽�ՠ_|��z�yS/�-d��8T/��'���Y]T?A���_��C�f�D�{���d�k�.WM�gE��X�v�nR<��	�v�^H�^��qv2�=k�i��WRg{�.f��(K^ʄ\���J��c�����{~��"k�f�>&}ǆ\o�]�'��U���ΡX�ŧ�U��I�*4,��'�v!v:��4�u{Y���g���ޑ�V��;O�S���4R���7���q�I�����s7�*u]{��L����
8:��2�5��(�v]�u��Y,�踽��m��(�>Էz�%��8a�g{����k��ݸ�`�S.�����^зb���..�s�Z�����F5��Y��\;���Zj�w�ED���̇^�h'�U^�f��wz�h3X��p9hc�(𜑆������S<<�L���M��|��J��nO{r穸��	-�����ϖ���s(��a�iރ�o���#��v���'x!�9�gn��ϝ;\��1��q)�94��s�tX|	@cYR2�#��+a�w�}��n/K�h[��3�7�2��u��w!C&KmH���52pZ}�"3=��EIm�vݫ38S?Qõ��Ey�e����z��9�wzX��Q����������[|����/`��q��z��5]�բ� +��87����̿�;�����{5E�]=:3Ѯ{��|,���y?d�_o�=�� �ef���]�R��X�
�D��\-�`9�+5E�w!�Yn���3�hw��ɦ�����\X.;�ҥ��
�m�R\=B�P�뷏<Ρ�Z�O��wtH)��j�"糲�qsNq�>#�Z{ܨ�:�����X�Qtj�Y�?}��MM��WY
R�y7���JJ��Xx;:蚝(򼛂j�4�党������������{����L�z�n�ۻq��e�S���>�(�S����a7(��^�����QT�u�mg;:X(fu%9[�"Uk��Fm����ϛ�����Z��p��L��/f�9��+'R#�{2��x6U/B���ʧ�h擔<yh�򥣜\ω�L:����\Уc랓|s�m�R���5�����z�S�bo�&� ��jH�[�8��5f|��*�>�9�h�iפ�~��z%�9�+����`~�טL0�$h����_-�]����jh�)������i���X�u���
��(a���&�֫F�v������XE�|�[�p&=s��oN�K*���&Gqwpr�^$�p:�xq�졨
�������VV�Ƒ�z�q��R��\��m�� 2���;Ώ-I��G;�lr8���zI��N�,)��ވ����ɟf�r���ڸ�l�y�%X��mw��� ��R༸���̛�qLM1Py̯+9�Zt�&p���*<4:�,��ƹ<����n̚������e�f�Od�g�*�/��^���6��z�2/j�:ؘ��ž�7�p]X���2NN�;�6!�N1�++9���+ѯk\�|��g�ݮZ�����ͣ�=�)5C�OX��JI꩏�1�~ԣ����]c0M==�7T]C��a~2���O�5���mv�w|�v%���5.�����;���F=����6��(L`�`�V�1q��bW�Gp�S�;��u���]`�b�w�X�]OR���]A5!���}�(j8�bR��c��^PWͪ�����疘�/�2d?{)�i���=��7�J�>�Z�b-���qf�;��6M���,�V5)? �:��q�|փ"������s�rdkt�r��{�D>�9B�AJ���&Z�"ƺV�[��$gu}���N4q�2�Yɲ��y�~�:Zha��y.O��R�2��ʉ���L�ͦ[�_=���F)�v E��W����b��o��u�j�A;2��P�	/� �>}i��OV �3ۡ�K��3ځ�]-~@����m�����-�ϥiG����gKD� �{l*ʞX�tf����"�P�6w,�|��gz:�|s��9S�j�L�l��\g��	��I�Q�\2'ޒ*[�-��|��~�Ok�wN�a�|g��1xm��>�^�,�KOD�$�����3nf�$��sn
D��Qb�:��PؽR��g���s�(��ؒ��T�+��yc*�+�B���Z5ΡЮ���
���3�</-������c�f��l��''r�{�:�o7�_z&��U��ǃ���Ta8�����l�3�E�P�����2�`��zr�oX��=��v̄���\eD�>]}�;�2��S�؟r'��u��hƗ
aC���_$W�\4���M�đٷg=O����SW\Z����.I��k^��a<[���yt߅�"�Z�}uG�W����F�^��o��Ok}3I��@��%�6_�Q�lF��X�/|���ft�&<m���٘�^���ٛ�Әm2��7/���C�r��c:�0�{��P��I�	���0a�}�5�\���X0b�p�2������8�V=:��O��w��f�|����e�L�:�f��^��wU���a�*��*�:�a'����s�����|���h�/�m�g�ng��Թ۩7��ZՐ��v��oJ�T���>Ω�θ���s��tt0M�)�tGhWuY�K�<��pOxY�K��#Ҳ/p�IإA̻`�1�J��1`ۆIC�0�����}���WrD��ޫ����'T=7�(�:f�8�#m"<�ܻ�r^�P�<�%��,�n�K,�ކv��<g���昜k�z#�Y��W�\����u!ތ���+2@{���+��z�^�4�#�4�m�=0y�h{�_o����a�7�-%��S=��<��=˵��V҉|*�1��he5R[짢Qոto
"�\�i�=+��_wg!��3�X3�Tނ�\�@ia�z�肎�g��n������l��-��h��f�=3���+��������@���G>*�j��ܸqߛK���[����?	��v�?�g��WS2.kO}r�m;r���Ӯ��Ȩ)���I��y}�
iO�rёR�*ʚ�lWLY���6˙�����\�F��}��Nh�l{׻��F}�I	��^���]÷��f���kiO�!��ŧ�V7ow2��r֝��ñ��zу�q��.�s�Z�����k��p���5"=���XUԡ��zړ��+{ݚ�*0��2���V0�uK���S��q�\e����d9�K<e�{~Pwkz��3PI^1AOs���A�^�-޿"r�_��~5s,�lu��K)���e<��-x���ù�j氊��cs����԰i�s7�|;��{Fu7)uFxm�b@��H�ֶt�_��q���2����HP{=3�zJ�qP�+Z���n��9�>y]I���Y��S"���ws��Q`���H�S2��ú:X�A���D%s�a�oV�,<xpS?]���˜ܦ��D{�"\���Џ��r{�mE�s�c�3:Ih~�7��s�%l��������yХ��L�]��n��XS��=ӟG.m�T+$��>������y�]���G*��.�2x�W�N41}��n1\�wf^s꼘�v�����5e_5�u3AfL��j�	�);5,���q�T���:ij���vQ�R�4�8ͮ�lۣkF%(�N�ƦZ�[�;Nv��/�V���u�v�P*;���A�z q�	߄�WF��*�e��V�K=����9ՅGp�ƺ��k��ZyG/0�^`�Wǎ�r�r.8�Ԕ4���}�m��gl>��6���m��j݀�=B-��́�'����.r�n,-�Q؞��DhM��&��Ol栙�[�ᏱU��r�
�R�B���\�W=Uq��DC��ē���LwY�SGQ�N��λ�N��q�f&p�;�Bso�q��ތ�xkRղn"��:@_b_*Zm[�8K5 l�{XϓV>a�6Ѽ��=�ʂ*@����e�j��.�w*u�X���hظ�x�e����;��9λ�K�q�u)Ҹq������`{�C�}����L%b�[]mrB���a�6WZ�	a����� 
'b�T���!�n)4����N�rd� �q�m�#�l<5��fr��F��X.��'�N�`�:�7e_nا��]�n�e�ۚ�<T��Y�V��r������4�q �;J�:8%m�.N��k��>:�w�%���F�PMuX8u�X�e"���iIU��y���v>��v�
�܌To�܈M�g_$+u�gSh
��o�os6v����m�L���$[��s[9�9Vx�W+�kpp҅��O34�B��5�q�抬��|�	�Ȟ��R�~��]���Nk�fθ9�hJ�!��,֝|��f.U �'<�w{��&:���$�%V�]�M��x���]���c���mqK'Gw��Ժ�r�qֲ[�-�px��&j�H�����\#k"��i��+�h��r��"��.ȼèpZC�~�I��y�n�+�k˽�0�ur�M#�_E���{�
Sz-�4>���:ʐ  ,�F����� �c�&,��`a�+3�=5��A ��I>-uMu�w9�Mv���-̮,���]���
�����E���*3U�:�y��LK� ����R�dH�uk�3"M�¯"�u6�&�!uyʥr�O�LE}Y�Z����\8�KC�2�Jzk����K�nS�L}+�w�F%���*ص��3�y������*|�n@�4>���x�@)�;�v]bN<�U���W@D��u�5z���Y�z����cS)
�X̺V�g8i�`z��6��x����2v.hUI�.�x�����{zU��|�����(�����"$>�!��*��Ɉ����&frL�)�����h�b%��(�����)"��"()
f�`�������\`�i�p��i������))s12��
Jb���)j�

(fH�+$�)h�����������3((�`��R!i���*��ʜ�����,��i*&�J"��ri�1�)
J*�!�2��B�s2�j�%�J�ʒ���rb
Ji� )*����h()
H�h�b"����r����&��2(0�f�+?~�ύr7Ʊ{۰���ݠ�[�m�Liw��]��Y�j�w�!wLI���C�*w�[����v�(���tyᛯ5�;E��~=��_w��g��w���������>ͮ1{�|f�9��;�Ӯ����V��������p�ٞ��M��{«�vR��&6�x	ro.;�=��󭼚FG�zv�/)�e�����-�q���̇�Tڇ�KQ{@�����f2P�mtǖP�w�_W��ǝ�"�SҾ�<X[L=��p5�q�>#'����E�:���Mg<�<��)���{�KH{��w����XN�mi����9��oz�6��t�8ǃ\�y�mGG]>�XOP�yp����.gҒ�P?�-�/n��	[�Q���'�*��͜�e�Nc��5>3B�@�6��R|���p󨸟�՘a��d��^��5p��v�E�r\e�{��˃��f�eʞ|3 w�L8ZI}-qYI���a��>�ފ���;9�Nʗ�c�c��}�P��.�[􂬰a���/*GDP�Ք��]`�����l'�Ƕ))�>j�A���Z��>�GU�r�^�����f]C���(9,���H3a
e(�վ���bP���ʃ������cb���wΤ�W�9g��Mko�v�Bއ}�s^:�Dc��і�U�}�G.nE�؏�e��<�pԹM7���j���;���ӏ���ov�5ԚB[g�26��M��Z�q5w;�����L��r���)%@c�¿��@o�yb^�e�����0��00��&:\���~���e//��^;~%]��>�,;��;��}2��p����R���*��j9��������Ń�W�J,ހ�Z��1՞u�_�b'	uR��!��ftw���Y�}v���6�L��c�O�٪S�����JN�R�m�	B�&'r�����W3��>��ݧ�;x��Pį�N�C���ڑ�;������W�V�%c �����1�޳|+�]st�)���u��qϓ��9C�������g�b���V�Kkr(����مx��&}r�&ǖ��1lH�C�ǝ�-�3��"��v]��pZ�7SY�͚�e.�Y�WR�l��7��ե�����9КS�V{3�=��9Q��냦Y��:��6%TI��'���*��JL��Oe276�v������u���f��֜�=��U�'�1�ϧz���z(C�O���;�����=X�{n�����!f���Ǉ�%|�VИ���B.:��k]���q�>(��˗��7I>����u��SF�����yo�a��r�ry�TY
�9�|�2|���ky{ǈx`�����M�}�8����z�V�:*m"�p*���}�-�T�ҥ'��@9��i�w�v�/�|y��5�~0މ��d�(񿆼6M�KD���{HU�7SB�Y�E��j���X};����P*���c�T뚽�r2�S"aD����`�dm!���������'*|5�y\�V<�~�u(k�i�9S�JW}/�U$�:��y+��E'4�y�>Ҁ��gd��Z]�8vǫ����JӸ���P�J$`2)���X�u�Sw��L�ηg���"xz��u���юS|)T.�	CuC�"�f̆�
������槏����C�L�D�V��֡4�=Y^\/-�E\%�χ���c�bp�B��<mS�1���
=��֗�t�E|�Y��S�3^W�ja�ɯ�}t��k�Y��D�J��_u�8�LA�1�@p޾��L�-o��l9ZQ��������j��f�#K�g3�����6Oy�s��`ϱ2 ��=����x�Q->����ς����h7�$6c/��^�d!<b�/����O�J��t�~�w�_K�S�8���ǻV93��@�b�y�<�[��6vq7�z����4�խ{�e�5c�������j�w������P�LRƴ�=f����l+��&<�ݓ4Z9�����]�up͢�>qV��.���Te�nU��'��<m�&p��WaFs��5�����'u�J�Z��_d�*�T��DN�ԉ`�2+�������ZL��q�>:bh��I��g��{�.n�3�Z���R�(zU0x��Q+]C�3ڍ�K��Ϫ:�/g��0/wc;8��:����(�a�6���#o��Wr�ru�K����ێ�x��s�/ ��͉��̈sNq�i�v�7=��ϊir6T<l �S����x��=��:i�+�z�������P؛�,�ξ"�9|^��[9閁�)q��m�]��a�{1�ʎ
_=:�{W�L�����fE�i��2��2�9�a������S����z�o�L\�dT�5�T3�ر�׊V���Oaܔ%�כ���ȣc������ 
���I���f�]R��໇��$͌@ꡮ��Ρ ������M�6�䧘���`�}C�{+��]��F��i��Q��p�`nz�)�~�+9�C�B���qFq1\o�+5S�:*8e����c�wҰم���;Gr�)q�u�Z�]�毳=��Z����a�b�E<-Q�"�㈞D8x�u������\�e>��O��*�ں�^����|�%
��LK1V*]d�8��a
/N̮����2��W �3�����w-W[z�%pۻ����j�CVNuQ�Q��kU�C�Ÿ�Ӂ��C��4�( WVP_9��f�|�<G��72�53*X�����l�L��f\s����U�U:v�>a࠳s��Z�|y�m��Q��\��x���fuJ�6o�5p:9X
Vjt�v��զ�-x�:�?G���>o�A2����R��"G�X9A�}s_}�|pJ�c�X���SAiӸՌ����H�S2��è{��0�(�&NRk�z+�v�Lc�=�i�>uXtb.�Z��
B��ٵ�-zxW3g:���l��+��
߫&�:��c����=.ܞx��+�u-���Uh���Wtһ���++\����6�}t�)���nl:�����M5�o�z���-D�
�m���^T����~�n�!�WiV˱amw�ge�..k'��2q�=��ʊ��p�}��}�g����ȱ>+���������U�-:鵠�]|{�^�'a��S�$:.�Z�P��Ҡ����2|5�P1����|�fxe;S*�����Z�J��4��rQ�4Ӷ�_�H{�^�X��СGLڕp�.֫>#�y��W�����'�J��ܥ��ʉ�(E*�۟]��:�GlTx�W:?[��r�q���{�=
����'��q6�0��@��h�#�e�4{���[��[�M(���&��	
�d��[�g�[��~T+�yСI���{NJT�y�\O���0���,����|uB�E�8�:���x�2+�y����;�&�E��})q^��=;��o�מ���q���&@�O)��X�*uL������@���>�vL-b�}#�gԡ�]	�l�2�&�~M�>����jk�UM�B;>.��Qk�����f]B�U%=��*����m���Hf=�r�c1�v'��u�IP���B�^K��G���m���^��3����X�h���|���p����.��~X�;��羻����[�����X�{�OX�'��K��u����bĤxG�CmF�o��=Ze�[r�ʨ��i�\�r�\��Y������|�,�8�9^��Q���:�J������ȼ��|���ԴM�]�\ŧ�1&=:���md�z|6gW��Gz��XZYr��v��V���w4�i-����y5���;�t/K�ZcP�hɐ������y����r~D��O92�E{d�W��z��Y�Z�}$*��D΢k�H�Aq�d�+wb�>����i��f@j���W�c�*m��x�\�<�6���"�0�K�=�fm��;媿o-G�z� Ǳ˂��Y;C��g�ܗsy̞�bT��	׊�'k��3k��p�.X��OW ��l��+����y���ƙ�BE�[��<ك��z�>+x�Q�vx9��-�ԫ�˖K��Ti�=Y��a��R3z��r��Bw��y����7���s4<�K�!�T�`��o��\^]KL�)�{)���,�׺���\Ln�{7ݍ"�o�S2r��w;����.zn�#�E`�I��(s��֙ʔ�j�L���*n����cڝ�h�F��67�~�O~���V��`?���#�����e���S�E>���9���;���㛀u\,��詷1??�d8pK�l�3J&�R䪦�f3z��������'o�B�>����\Zqa�oW;�<��<qʘ�*P��^��3M��Jg�$���U����E��r�I�^�5�E㊝_,^R�������9D���V�DY^����֥L�bۤ���g�+����f�23<5�*�l�iA�%D�]���T�{�6��b� �*dD湷�o�z�P�X��>�L瑱�v�=�[� ����nOicp�B��+|����@)ik+,-ÑcQ��<��(Sr�V6F�3�iY�zJۼ�����+����u���/dR�lݥ������tA����]7W�Ԙ�n;�Cz��/�.�����q���ާ5�]�oB��u�YIoN�����`mG��y=Ub���xN��t�E��s���M.��bP��F��4�V���W��V��T�|��(������{o�+�z��g����a��1��yW�Mw.E#w!՛��.�9�9ץ�ʳ��5k_L���D�:��\1��Ü��}�b�����3��0g�3m��X���NO�Y����Ζ�RnLqh�'�ip���՗��^�;/��񘴆pKS+}\ڑ��I�����7�@T~��M������^���O1�圬iψ�N�*��P��/��^$���sh��l�DÛ�EǶ4���}��Q�gӪ�w�l:f�9�L�$�5�\����p�yq���%��ζ�u���{2���6V���n���.��دL��߻o2��+���S��B���3���J����,����^ ��x��\{�=h�jy����~��T��Us�|�Yx�,�/M	 �U���:��f`S�x�]6��+�OG�!]uU�oz��#�lGw�xՏA����|�_�[�*�]q@���V^��3� 15Iq`�܅c�7~9R�p�3K����;�����i.�*�ǳuM�����)�LT��K�.'�;��k�k�P�������@����Q3�(}�e]�%��c׊k\3lw���a�h�v�g���o�<�2������H_��I�����\k{DU���v�T{�'��ĝ���v�-1�Z�BX�ȇj6'COW
Q������s�.#;<[�U���Z"�f������PpS�8v��V0�X��ez��X�]t��FQ8�t����yae���ݺ��	*�b¿t���������jǍ�ܑyN�l/�6[=ö�����;����9�1��ߚ�+�pXW��z%蠟���e!|;W�Чa^f��X�y~��q�>ʤ��=�Sυ���\SV���:�/��dg�����N�����K��={׾�����O�yw\oN	�Ǭ�+��
a�-:o�_���8Ԉ�θ�x�}j7$柺��9���wmy�+ݾ��;�{�T�P)��>�}tCV�`�����W�vl>��O������(=l���P��0��]r���O<�L��:�[k}�*G'�x����<�"�×�v�b�"Cʻ�t�.�{ᢀ��VkM�����Ps;xSzM�.U�g"3���Z�QaL������r�{}%{��;]Y�J�zMqm���e���� Юf��6q��=� ���[��b�j܃�m�f.�t�)[���k돴�i�~R(�2��:mC��_54��{�2ESj�T�����;�Y��3��� ��.�"o�S��GD�f�Շ������Ƹ���a�wW��;���Lv]�.[H�B�~XU3)���@���=�/˜������o,�nܭ�{���|�"���J�0qJg��
fbt�\E�N������1�7����Μ{&����V�<�ɔ�34 �l�A��%�>^����B��ڸox֚��~���z��8��}�����iw2+�y���w�L0�$o��������.����bR��=��9��Na��jz����qø{�9h�U�;*�Xu�Ѹ�����u��Iaᵖl�;�����>�{ͦ��l�ꪷ��.���-xd��7񞺆*Y�.�ew���+C���"o�9P1�!�t{$�]>���b��JIV�
�;r�Z�S7�v�i���N��{�"�6��@e���WٹA��ۅ�ݫ���W�0�>"я���ߍ�ݽC�+�9;�|�X���%kySRԒD؁���H�!ђe;��1wHо�f�]�ҕ�z���jN��lIҕH�f}r��a�*(�殧Yu�)��^�|�V�q:���=�1�j%�P`�8�¨�f��^�\zgJCM��/�o�+KX�|��b\]�s9	�­7�h-�j ��P:t�f�}�t�K����N�-�/�PXP��躓&�Պ�B��og]���oB��F3�^��KiwV])��r[�̝;�u`��^�w=���*�I�pκ^��ΝD�`m�3��Co]�͚�[�1������l�Zoq9���0c��#����l*���p�i��k�u#:]$]���*N#��RC�U����ӿ�K��*{�e�o��.~ �^GLg-Ow���}��x�cE��c�X�����O�W��>���;>O����$� ֫*�f�s��m�	b��+�K.K�I�,�3c����V)龀@3�-��㽶=}0��L��8�j��Z���<�VBx��r�}�ou�Աc�*n�zt�7^y�b)w�Nw�]�6k[r��x�cB��+��R`_VOd�4f;�w�7^�o_M+(��#����+G+-�N����^��!Uq�P!�&��y��g*^���٨�6����훬�}f�#	���t�
[��0֣�
ɱ[u�.�e��j�Ut�]	7[���)�JH,�2�q�B�]�ˢJҀ��Z� ՗.��q[7��ޭE����G?.3v���n���5;W��\�r"�m���_7J�8��������Sj$�ޫ�����wX���	��ͳ��j�z�h��@���t���n�`�/Z <��X��j̵I|��$����v��ٹ������,�sn���8A��}���9��'�PDOq~�Ǣǝx����ɕs���g�x� ��Y�A�(�W��M���p>nsj���<�M|{���ɫ�hs���Y@ʷ�DK=�g�H�g��+�I0X�w7��Y}�g	��b�J#������-<��%^m펵n�.�G&��T�xW�8y�0�4�'���o���'����C�Ý��h6P߬���p���k;�-��8KR�������uc,L��L'U�B�N����D}����
x��moeh{��c���4<+0�ۤ4[�Т���q�秋�{}�a�2��O3e��š��=�hf]�w����_�����������_`T�Z�)��������c6��N�������D�]��n�}��q���)����p�S(oPYc5Ik)�6o n�����w�4�	���|��u�B�i�}�}v�w�{Iz�k�iOE<ةY�N�f�.���cS騙jgu>�������y�_i��?|H �f�({���R� 0��3)�L����i� Ȧ�iZ�3�(�̈\�,̌�����#+1�2&�,�(2(\���$��*��#'%)���%,3"�Ȥ�[1�0�(rr�i��iZB̢������(�s1�3�"����2L�S ���j���
���X�� (())\���"�2h�l1ʲ�
����Z(�����"��(��2G ���$hj���,�r����#*B�̤2P�J��V���0L�����2i"��"�ir�&���3!�Ƞ��&���3%,̚�2E������*�$�2\��hr�ʚ�*����# 
Ƞ-{�x���{�W����{կsBb^��i��z��M`92zWa�֜�@W}�z�*��WW�͡�bx�
��q���q-��n�Sk|�.�6��5���5g��8թXp����&1՞e�C�jx����NN햼$j��q<���JӾ��3j��^׾^���u;8>�ᖖ�Devf���WC�*E��˭��5C�N�C�}x[X��F�rt�hf�5c����u��j1�����S�b�r�bآ_s^�1��琍C��d?{=�%d|t�򆦜�}�����hzb������"_u�HO�1\j�o�^��o�d)dcU���^ķ�s�p�z�C���/
ug��q�.Y.�ʍ#z�=ZY|�n�kj^V^���e����m���Ten^�����|)W�]KL��)������Q �u�T%���(̽����*^s����.C���I������6��;ޭ�&K��^�ȇ�O{g��׽�����	��gҴ��]�'s��M�C=�T����ք/�x��ꝏ�K�Cf;~F&s�������*uL[��L��ρ�vb�Ǝy�Ŕ���h̬�)V�u,34*<f�o����*�Y�%�G�"k
k�4�AXi4;D���2�Ou.�/��@�Ўɭ�a=�ݲ�nۉҋM_
���r	��u�F���$�N�7W��_c�luM��ٌ��.γs����}r4�\� ]cd��^�l�I�Qυh�8:��թ������X}��}�J�Lg�,O'�2A7#��N���ٝ[t��#Ik��N�.��Qx�W��l><T��ݟ��m�M��{Ǘ�ނ�I��ZR��1�.���]���Z]�]�1^�p�o�t��%�Ń6C�v�sǽ����4L�S$�D湷�hk�Z��X��Jg}�p���IE���17'�8e�_c�
65����i~KK$Pٞ�G:y{�]�?�����_Q'g��w3ڥ�yx�i��P1�3�����{����,af�r��c;��3���vöt=�Mx��WN.c~�cuCO�v��h?�ݾ���l�]Ef���O �qƳ�3>ޡԪ�Y����ʰ�ÍTG�k�l\Z�V3C铖M!^暻�K���Y��#%29}G�eű���Hgt��^�c��н�>�� i�]�ZO|�g�=�J��wE[��7��u��3��]�^��)�V�U�ߏg�)�� �	zݝZZ�?��p�v��;��KGZ�N�]�����y-~��I�a;kh�0��)㲺�^����t��Z�� ���֕�X�c������S	����7�Ka�u1l�[�v(�~���ɶixD۸����c�;�9U�X�{�>�ty~������Nv3��O:ߣ�zh�Ҍ7�tͰq&F�C�@>��Iٚusw)��uo�;X
(f����}�dC�s�sOc�Y��W-.G��e��<��E����.Ӥ%��ڱ'�j��P��o<��:�����z�w+fߪ��t�\|#����SEs@��i���_�PL�ƃ�=2�.;��
��<��3땳(Y�z�y6e�h�x%��[=۞�S�7���㖋K �L�(T=y@�W^KM���WRgz����;x��b�������.u��˕�*ņ��$<3���
��4�6'��B�T���>��o�c��}���shC�e\XsxU�yq�wdC�֣b��m�m(�^�Y�pKy�2�P�s�+5�f�"+�u�����(�������	XlÎ�b>=G��+�vӢ���[N>�w����/�ۡᲂJ�X���2��L�`<K6�{�O�ٸʙX����|��\�K˼T;������1ӵ�kH���¿�^D�I^��5�!���k-����9����C��裨��r�:׭�aG��ר�C�xS^K�A��R{��w|ya�RUY;����w}5�WK~�L�Z�m�<�Ι@�i@�_�=w����M�&����.�j�哩b��-9�wt�Wcdq���%�r�H��I��	W��Ν�\��/��u�Z����6�E93Q���n�.�2q˯ΗZ_(�'-N"5ج��mA%w.>Յ��mY���3��������Ԉ��3�Sc|��z0Ǟs秠��雷�3��u{%x�h�n�J�z�	dcT�*��u
:+<��6W�T{EI�\�'`�&yA�fX�s:K\u5s�p�ٞ��&J�>ꮵ�	��^;��L]oI���)��E�n.i��fΨqԷ峍}��2E�\��qiԓ�N�xQ�7J�Ɋ�jr���`U�.���T��#�z�jm[��d8��8��ں�u=F�����T��>�s�{��	Rу
��eU30[�/*�b�t����=�-�s����M�O����]�W���TԈ����$��)� ���(긌7�uؼ�����U~Ï8Ғ�杙[�Q�qɌ��x��f�����%����)�c)�s.����������P)_gc��{~�<s�"�W�%���� R�#�����xg]뺗W�Cl��(��u��P��`N�;{[un丬(E�Z�8��F��qm�΂l���L���kE
�AH�}�=���vݫZ9�[��T��/r�"� ����j�m�;��
{�f��nCMj��ӏ��w<����>��a���&\|�Қ�x�%�i��U��^\���C�K�&�R;��P���6���J����{�G\ڤY�C�d(:��ڄo���J<���KE��<�l/.��ݗ��{u�|�.��2���kG��+�Z��u�D�W��E�:�*[�_���S�3�g�Y4����`I��s洭Pr'ؼ:�7r���Y��Wl���z\��>[u���ĭ�i$@6e�+�M[������ab�xG����ճ�*��K���7=��T��������z����k���F�6��i�}��
.fՋ��:��1��"�#L�MI��s�ѐȟd��p���Ů�k��X���_^Ԏ�ݙ��s=}~�$�P����������V�U�%x�
���Z�Y𯹪�1��SP���&C���ѹ��f���>~��3���w u��z�2�Q;��BN-�ں+����s�̣0���(��<Ǉ�N5�si�7� i�`�a���'�Y�\eJ%�*4���f�X��~2�X^+�~�k�wZ-!�s�rĽ�͆�4Y��ޱ���1��]˞.QG)?lN��ξy�o�9b�.V��^���a^k_��מW��C�c뻽�Oz���y�]+NY}�u���4]b�Is��Z)}��-�h���
�A�3�-yq��.l���ur3o{��5����}BO�ꌡ���!i4�>	>^�)V��y��yq1��,����؏˭����stE��e������y�?�z��	ٔ���0l$�n
9�Wמ��<��]<� |@���bƅ��t>��z������w��I���4?��`:��v������@â{�[�YJ,T����Jgy��K�C�}S�j�{�	^r��VR��@�Ex/˖��~w~�&�-4�de-"VCa�������S�CX�cL�ʘ�+&�en�}w��ׇ��m��w���[t���#�]E��K�:,X�|qV_,^U��k�ّ_�X����g�Z�̷�w�#�T��S3���% ���*W^]�(b�L�#�t��y�����=����X�7�`��.�=8Ûx&��u�M,SԢg7�p��3��&��Ԧ�15nr�o!�{�<��ʬw���K'DZ_����6g�Q���� h�S;�<S�ujub�Җy*�g�9���!�@p������o�堋���0&�se��7}����I�`�z�F����]kA	a��?S��}/*27�q2ḃv���Y���W��ܞʼ��wf[�e�-��{���wN�2rg$�q9�c︻������5j3���7M�ʧMD{xL�WU��,{�����]�9��t����Uz�r�D�f�qx?�7�#����]��cN(��T-��]k�%;k�U�b�\��k���\�<%��y�?�'�%Z����{M,ǁuwV�6$<<=9I�G����|}��.���%ӳT�=�l��8��9���/�)��1�>fi�c��Dwv�I�ӝ�udC��{��]�^�!�wJ��|��E3��s��=�6�����Q�WIM�g��2J,ϓ���jy��Cҫ
0��p.��Wm���Ы�-�Ǧ�^ovAV�����S�J��P�o�l	���}%k'�t�,Ob�z�����/t^��.���KQ���.�R�v-�'�j߽*o<��	�|E�\^!2�b�۷==�o�k|�3>����n�D^'��U���e�|�����2#�>�s�u����*=���;��uA}'����؁���E��)�`�P���K�u����7ԫ���#��WD������;�n/���ʄ_ҬXnm�k*��>&/.�~����C:\¼Ë��t�u��w��
u�H��d�l�J�\�1*K�](n+ɥHҷ.��j$Ƙq�᧮�h��0�~�4~��J�jo᠗Z^w���t����8�"���͟�wt_tL�,d)n��U�v�Ϋ������y-2��{ �*R�A����ӣ���8:�.Ļ�!��X����X)N[y�[���Xx_k��f��u�Ƒ�Xj����ڀ��
~F:G|%a�:��JQ���s�_lN��;�F�JL����;3�j���l����,+�L��3S>^<K>�Y#�����0���:��#|��A/'��u��眿�:v�>k�1�aX��?v��:����Lnw,�>�9!��w�?(r����1��C��f��\j�\S:��Gΰ�����͌�6-~���W���#f��(z7=���ܸ�Vw�����E�>9V.�+�:��h���vhFf�uz�����`uǮ�{�3e���N��W�M��Y����[ܫ�HDɗ�r&�.���^K�z2h �{��ȡ�+L[]k�}C��s��d�_h��9��+4�<��v����r˃����C�LP�^�J�sM`�f���:���q����C�����.��C=)�
��7��kRI�I��S⬎����糲������X̀��.�תG��peeY8��V��1=�`��L��@�[�0:�>�/qͽ^47yI˳-��U�+��)ޒ�׳�U�u焩�Q�팔3lɛ�X�h��A�_d�QY0y��!�Y���x���;X�eN��6�b�WF�c���FNQ;xl���kOc��:���P�,�US3-ݗ��v Z��C.W�^���2�\~>=�#+}L�Oa�U�S�zu&��1���}�)�e;S*��(�Gw�p�{�7G��gmy�U��u�ܮhQ�s��xM��>3Pw��W�̽&}H����:���򍅗��fW�B���|�F��f�o�EW��~2+�x2[9��	�ZIҗק{Ȼ�n[v�����������.r8l9L��P��=뚳�a���鹄�Գ�Uј�l�_-E�#|���]׭C�n�1��DU1�P�χ7���q�L0Έ��3���/s��YꙎ��.�w�ϱn�~�Y�A�a�� �������x��:�:�뱠�tbԲJ>V��8ZU�O��2�\��k��oÄ���s�P��gj����/1�۬*|�|J�5��w�®����8�r���ώ�7X�]�QǺ���u��%��*<5a��N�'��n�k�e���G�{^Җm3��lH���^w��o��3αM��!��R��4��i�E�{��{ҳ�'��%'��:jV���e�j�CbJ_b!{�7Y�YS�� ����	��}�Z,��M�s:s��-̰w�cD�X��y[�h��q̞��)D��{���V�k�"ۿ�kL_�\Zꖰ�$���]<�6���;��+#S��y���vV��z�:԰�+�����kQ`������SS ơ~��e��u�5�>�����.�b}��F6�hze/.��ɡ}P�x��V]�~A�0���6�3��ݗ��>�5�ء��n�3��=�)rcb+G����{���=YRa�4V�n���^b>�⏧��Dߒ3��5=բ3C�U���i0p�ӑ���<��k'�Rb�ޭ[�7If&FM�]���6s瓞���n�NƆ�l��xxWPω�7�'�GW�Ln��.��0]O�ݮ8)��bg��p�A�1gO~���yX#C�����M��;q�z�[�n"LixBU�B[�������W�|��>��5{<2d8IYC�y�b�����=Ϛ���a�(�����1/
�X������Of��,>�=��\�����:ھM���ƸK�ԫ��!�#�1R��K��ōqx�����>��n�g�}��.���U��I�{��sF����u٦&�3r�+)�x�KQ�V-��2��hZ��N\�f;�:���|�k�>�b����l��X�c��4uܱwӪ/�4�Of���o�CbVk�)�8��I�,�+/�lw��7jsO�'���;sI\��d�|�_�'bHT:�%B�X�x�`�O���so!��瑐�g���k:��"z�&H�+�^U�:
�{��ڹ��S&[��]����ٕ�s���8h��#��D��)oE�!���TP���x�CwO6}�H�����iX��Ԇ3���ڌm#�p邲����]�6=�B�NJy�Q�X��܎+4�㓇�ؕ���O��יk���h%�3�dz�^�7Э~7q���>MmJ�xMeE
��*È^7�[.y�O��~�z��x��Fo�������I�4�°Q�ݑ��Vԛ�[z���I[]v��N�����l��h�狞i;l���+<U1�H���7�s+J�2�����ߚ�;�� }�G�<�R�L�n�����}���6�4�4�ĩ�tKm|�݇���5�����9�B�c�\�E§���#G$宥 EMCC�;��'��H
��6���C�;�6�De���ʗe�q�߶���n3� �nA�]ǚݧ�%�:}�7�����M98��c�zxa_Oi����8Gz��_~�w`�e��դ�M��n�>�v�<�\�*�jW��Eꬸ,Ho��{\���u�2��.;���:T�0�[6�v�]'���c����P��`���μ���y9�<��6A���u�p��NXR�zC�W7j�w�ˬ ��u�r19L?iM��.Ԃ�T�-u��2��س���e�z���,�L��W��0%le[���u[�H��T�Yku^���@�<����'d�"}T��I.�@�,�-��E��]5��U]�]˩��u:�!3��\����}�Q��4�%{֦�^����WuqzVO"�xc�p��s�.{v�b�n=-��|����l��b��g3�a���`7��]��M��m-�tr�x�P��,�w���A�&Ûɢ�M�}+iֹ�k����Ԧ��̨����Q;�2�T���zd�y惔ot<�wi�ؙ����܇:`�M�֨�oYvl�����-%1kU{ R��2ݾ��ė����T{,̡]F�iD:;f�zp@x�x�^�w�{�qx���>�թ?=䉝��|�����_xvZ ��uȟ=HśwX��zZ�DLJ#�JE����z�W�t�9�@.y�i�����m����ՓOdjYٱdϔ�K><B:i#t�^�usR�r��v�DN��'a�=���;V�p��f����𩘮�	y6nTFiꐕ{	����Z�eV3��tZ�VB�֞s�]mf�^u��a,٩�v����=Y���Sg�>�lM˻�^s�6�E���2O��G��H ��R��ӑ���44V@d�YDY�UA1aT�SYd.�dAE#E-�26F�Be��C&@dQIf	FTf.f&YCT�ASHRRPfcYPa�eE4��4�Y%9�eҙPfb9RR�!YPٌAHPPde@�9�I��&Nf&fM5B䡒@P��B9%VK�%��e�9Ӑ�B�a��TQI@d�CM5�E	FBeM��B4�AU�KH�!��Pوe��!DBPPdd9DNI�I��%TQ	�P�Ӑ�8*�������Jg]���\2f���N��s��i�hz_N�W�CB5�mo:�^Pf�V�c���i9pt�繒��|Z�z{&��J0�����DH�,IQ�.�F9e�P�p��ꕥ�o�(]���Z
�3��_����,�3iY�8�uh�d��N��ͼp{�W��g s�֛��Ã2Iݛ�I:mMɝ��Zfmn'�������G�%��a旀�d��'��li�E��4�K�Ɖ~˝]!����%��f���χb�\<2�Em@p����+�R�9fY�FUO�K�x�}��u`}�����P��V�𘗨eY�]N�N/��VY�G�/*��(�o�9��܎2��>{,�x(�쩃9e���bǥ�x��8׌$ޮ,)mՅW�aWyd]Z��;QI�ǩ��c}�v��񘴆|0'i��)�����D�	P�����!��)t�q���(O3\�WGBoT{S�C���3�����gt�EV{����/Q-l�o]���f{��(b��P��c:'�u�=�����/�E��J���7u��O=�"�DcW��ؙR�+�P�o޸a����2!�O�]>��e�S��u^�s�� �K)A�B[�K(��wm�fI���5�]�h�YU�M�g=����]*�ԕ
'.P�}��O7�ZsJW�0��,��rc������K5G�{7�4퀩Mp�v��m����|`��n�MW�ԫ*�7����QY�l�����M�k�µ.Dx�G˩R����5o�Csy圙��Z?#,�;7��Z���n�w�5_=h$��¡~YA2(_���%��Y�����{���s�Q�w�k��.�g@�]��z{7�Z-,�L�ʗ�����Ma64��ǛyX��$��3Ƽ��Z^�==�rP��>�B/�*Ň�{)!gCm%;~����Y/��W�E�	��ݶ��bV5���6�=e�ŧ~�*��B���ȇ�Fŉ����{{�ͧ�eG/�V���Os��o�Ci����.�����21הx_�M�o
� ���q�-�&U�h9��=��K�㬵�X�������3e��,+�L�ᚙ�b�)HC���n�Z��m�V6V�a�AC���9~s�f|�ڀ��<࠼7%�H��ؗ�c������JnӋR�e�m�a�j�%�Z���}u�ڨ�ꗾ��;5��߰�Hj~!��2{TG�n�=�n{u?����9f�|��,N�X>BWM���6vGO��摮�\즜w�<Z_�����{���$�������w�5]�`۝*JmcLԧec��󱆪�����N|�t��K`y�CI'>O\z�qas��O)�#Y/�qT��ye�2"��h��������]�՞U��w4�X5��>�us��:4�=L����;�,F��u�ڸ���n>�jͪg�w@J���w����۱̺�3'L:-J��/�Ϸ���̱N�(t.�4��\�u�xpoA��o�wy��yۇ^�q�Kҕ!@�||�J�sM`�f��>R���k�x�u��|���O�]bW뇟�ti��e�������eU30]Q�ⴎ�����a�쳛��W�����/e��M�*��P���q�=�nTX�Z0g�B��US3-ݖ��@��)�vű��k4���)��!�%�|�f�=^5��ڈ�~���Q&)L�(S2��v��؝F}�^���x5ͤF��/hwlȹ�G�zM�ɔ�	��l�A/��K>��z��{�L�Xg��{�m&�q8MY�_L�V����"EX��-���0�p}�@O7E��t������+��Wc�:��ڬd5��5nS,�P�������>���9U�Z9��g��@�>y��V�,������j3�]\�]f-�(:��ڄo�=wV4�F�n�kw�t��v�������Y�(�:I'�xU�������^�� qҕ�����L��+n���V�;xA�)\r3�Z���4r�**�ޯA�����"�\0�&�(�[Q/��z�܅����"L}p@}{7S�=)9��q]k���|�9�<��o�M�:�U�E�����	��'�j�c�Cq�rd�φ׽+wИ��W$�v�ˬSمtǾ�`��ā��3C�j�M[0�
9�>��
��$<�'[��^�Ԛ8�87:�L�|'�mg�ز�6s��/zrl~�����A��z��j=��e�r3��۞k�LuWy��/��l����2x��{��W����;��O���>�6�y7�C���vz�n8�s{{U>����7s��:�����7�r�8/1u�����\~�1��$hq>����0�K���޴gu�J:�bQ9�'+������=�Wt��x��&�w̼t�Z��.����R���Շ�ٲ�QT����z�y=8|���o�q޷1Ki�/��I�Sq���Ym�������{����{]Q�B���������*J�BgG��>��\�-�I��B]���v��;t��W����2�1ǚ�SƬ�{�bFh��0�wG��2��Ʉ�p]n������{$he��]i�a���d�5H:FL���������@^���b[��[{��mR��bt�xS���k����g3~�}�>ٺ殢��BNV�7�ʧ�;�˦��s�f|�r�/Og��	���e���SazZn����h����}Q�{�R{�C��i��U<9=��y5z��Z[�8�'�9�>��[;�ӵ����ەbXk�:&vR{u�p�������{rqɱ��j^��<�^��; 2���z/�'��.�5��ïS���]�!��Y8x__Ju���3����^8�u��x|A�˘Փ�8���7W�[���;�n<Yu\��s>��[�v�,I�φ����^�7��f�ĳ)�SEOO,kޟ1�3�s�S*����L^䡾�lw�77_��8���f䮶���Ձ�}T��x��^�3c����DN��>����98V��)�mo�ړ{��U=�ޚ�l�ɍ�p������)��{\˛{!	i�Gp@�/
��IC|)�1rJ�{M�w��oe(x� q>:���k�ϭH�����������q!�O��S�,W';��FБ=:����Ǖ�.=�ܲ][�q����3��we�zm��9\�gU��k��b]R*������Mv��2t�R<����O��{N}}���!ù��[��W���ڡ7��y�1�����=�rk�^u�z���t�cй��T��e_G76��:���͌n�ntϋ��x���򦨖�uCè��5+s4�z��GC��I��u֟�{�ktw��s�}8�g>X#.֪�=�������wb�j�,�i�`�a�չ��=�3c���nN�Ͻ�����y�|�.���y;S�E[g���!����M��G)����}/	VOvE'�Nf��ǯ~����6i}O��A��n.>����y�39�������\�{zd�����ەaۚ��x�S��?��yk^0l��G�[�iR�;d�ګ�����Ү�b#:&��lk��W�/�O$œgni�_mJ���sL�z�ޑX�p8}ۓê�%�]u�mb�>
�yK�;�d����Z�]Ӣ�N�p'����w�I��lX����/�>��8���{�]�d���:'�z�XF�tQ�x�T�-�n�[YZ��[�q�LdW�{ʣX�ƻ;���㲨��8j҉��Ԧ���0�wRsgsg� �ߪ�}����MOl'5����p���Y�=]�3��^c���n˥��l�o�/�pS��^�y�L^价�y�h��gi���}�����������;U����됬�1z��xN�,傽&��wLu]=���nn�{D}�3�f���z5�7���?L��kۊqsO;:í.W�S��;I}�?������	͹���y��T~��f�20�+���o�W��s����߁}3�:>ϮM~B�h*k�b?k�{��՞�����b��8t�͌r�s����|�{�7�SzOb�;��t����T��/<���\�T���Ώpkfᧈ�*R�[�=��e�ng�.N>���8�Xs����/��	s�+��N;���)��bޓ�j��.f���4�9�	ں���(	!b��������i%ӫfO��vyrI���s���gIᛋ��X����5LO�Uie�[j���W�4_w3ycMݾ]t@w��fC�J��zW��gj�����:��%���If�a�X��+/("Z9K#�+��,��	�W&�@��?��qf�{��N��?L�{ZL��V�f���
"�׮�yǫn9����� ɞΧ����r^�\wn�L��,� ���Oz�ve��i2gt,�}�`T����;�r{�og���h��q�X M-�ڒ_kj��j�'�"=nt�:�h����އ�K ]��{|�v������e�b2��C|������E/���=����O�;&��_gN:�c`ΗK�1l���a>��O
�4�*Sʎ�]���9Y;�L���i�����$��Fwe�*����R{�:M��xX{���_�Y�sꞫ�s�Fzv���6&g7�7_��ӷ(�%=/Ի�`���&�pʎ�1����y��x<�7��x��-��L�x���޺j�6$̧����}U��v`Y�����k�����bz�mG\��[�^Zpm!z�����Z/P�����e��ܕ

(���̖���ר�|�n<�X�)WY{����2��t�r�=��uyg�v���}@���jn�"��*'s�Ϯvn-.K垼��eP@�yAV���6v��&r�-{�;���ќ�����x�;��^p�6I����+�X����3}�[��d��f�	#�v�^:~Нz�^�X�e�t��v�Rڼ�{�M�H���͒�OLjs�<f�q���)m2ł�d>91��h��u���u>�^��:n��y�����ں�+H�y%gr2�<������{�����`��f�_<�S�9}������&��4!��x'ý�Y��<mN�����M�������>�Q��f�lXuM:���^�,������uɤP������C!t/�Vt��<0߶jUr��w^o���~���&ܫ��hN����m]?V^�S2���,Ynx�O��qz�}�����E�$�S@k�xvZ~���2K�s�l��g���7��R�i�+�\�zltRe�kO}�{�ow��޾��)g;+�BƜ�V��AS�Zz.�AW��+��pL	�.���:3bS�Uy٬n�5����R�*u�<ɛ��F9���n���CdB�6��r{�P�,_kȲ�U�C����ƣ��y�W�ں�k�}����.�V�Ay�57�;d��1�R�_7%�f\���1�4���g`�v�q�[W����l�S�����vnSʽ��v�ۛ���;�b�n��"�G�2�	��S��)�'7a�j���������
�B�������2v���KFrt�F�w��͓='z�����Ok�Q�MKk���v�����O�v��	.��po>���zU��{68��'y<�׫%]b�G�'�Uoش�kŵ=�����Hll_'پl����ɯ���.�?\���ȷ���_:n�
s/. �uׄ���C9�cnt��<x��τ��%�=ɣy�i�Z�93����}4
�֟���^ns[r����/+^{e�s{|o�3�M����f��:���;,���cϾR�j<Y���̋�D�IΥ���sw�hM]�[*����>�G_�{�^�ED����+��ED��* �B* ����
��W�DTA_�ED��+�B* ���TA_�
�ED�W�ED��* ����
�uW�(���Ҋ�+��TA_�TA_�����)��MK� ���8(���1$��}UE �$�J��)T�)H)E���%A!ABTU��J���R�*�AUPE"�*�Q	I!@H��(��$T�J�_cUJT*�	
���$�R(�$��jJ�R% $�	"%H	)*��R�4U/`h��"A� D�u���@QT���I*E*�B������(�	� (�I*��U*K�BkJ����   q�zk��lV;NR-����u%�����f�M��U�NJ�S7"i]L���w!I�뻮���F����5�tI�j�iEΤ�EHlaAJR�D'�   ]w�4�]j���)uf��;����[5��ڻ��m۷s��Wj��;\��ӍV��Ϊ�wml�uS��V��ݣ3Q5��ö��C��B��$(�#X�/Y@J*�   ��(P�  ����  P�ۍ�P�B�
3��P�
@ �L(t:44(P�J� 
 � P����Q��׵j���l˶�ݭ�p�uM-ڝ��ۻS����
��I@�� �� =��#�m�.��ip����-����bva�ַ`c��J�]�sm��7c*��v���vWl�ӗj�t�+��nݚ��j����N�
�[j���T�%�n�  ��-m�ws�wV���sZ��Nݳ)����5��]�n��������jݶI��]�]e۳���k�)0wIJ%Z��1�n�٪7R����-���PRQQ�x  ���.ڕm�U�X�F�+���w]����m�㖮���m��[�δ��JS����wj�p�l����qڇW7:��D��T�Q��Mnj�ER�IAي�Z0<  #���^�NuZ�:�v���n��T!�P �`4��u����n�:L���sS٠�� �$%%KX�R�vix  �� �] �A�F  mT� h���펀v
�u� f�vͩӎ�u���c����TJ��J(�锕�  ��@��0(�U���: aӹ��J�@uN8�P �&t� �e���-�\� �,  �4�i� "��F��   Gtz]�v�u 6�N�u3�mR�.��k��gZ�ܹ�vӜ�\ h]�r�Z+[��q����Z��i�]�÷���eIJ� ���$�*   *z14��=@ �JR�  �~$�UR@@ $�DM�J(V,�����B@z��L��$4!�M��!M�k�t��Y��r�D�߯�>���{��P$�	&�! ����	!I�rB��@�$�H@�u�$ I5|����M_���oz_W��=��|ӑ�Y�Z���6l[�H�S!��p��F�v�85j��?L*��v�<YZ��H��F����²�+@���	f�S�͚�s@�u�eF� T�4���+ �+s��[�z񂥙�aZl����l�L�x� ��ǯMG����ZfQsw#���El������X5��Mb�mX���v���!�@E;w��E�ہM��Z���^-�Uk�z�F��**W�D�̴�Y�:"�*�����mh�M���uּ���L+T�Z�X����&�d��i��a\g�W�[�R��ࣰ�)�H!�W��PFs��J�uL�.M�@��SB�ʍ>�F�Vښ2����TZ��,�|X.�݂>��ɇMݠ��N�Fıj��0m#5RՆ��Ă0�� N�^,��+ ��[���e�]�sJM��o�@RJ����Z�BWn�5�@i�dWRܼ܅ky�~[w�^5zl�~:35m��n]�C�5A�^�[X���HU���Q��6�p;;�\��w&<E��D�:��S��yw���V���1�h(��\ųn�n��woE���5��N��~s��(G6nL+��hSmJ�4Ty�2�ô��e%�j�B�3A�u=�&�B�{b���˙��v� �F�i��w�E�Y��df�r�T���,��\Έ��B��R#�
��<t�CI�/ �,�>De�QU�7%��;��F;�uM�[N�F3jjW2�H�{m��`���H�`0ݧ��АB�7�U��ܙV� �^kL��ܛ)
-���y�����ř3C�x#j�H���BI���;�:��І#���IV�Ӵ�sHջ6Jn�a2�S��ls�N�Q��S���Hn�ͼ`��Uw,H���#���P������YY�#����K��ۦ���+(�*д�ݹ�V����՘�K��� i�b9Yk'�	�fKq��t�t��4���B�i,ߴ�f�t�hn�%V��0���$�V��<2n���cm6jtq��jZ���+ZbT��XX�n(:h"U��3���]K��c~/c�T�Y,�rSx�ږ�U�ЂY�P�҇(���!�si<[F�eq8^�!Mu*�ͅ��N޿��aP*�&E^-W��N��c�zSՀ�.��nv�m��Eآk�K5Cmf�#(ig"�%##�t���p��Gr�)���&�����`Ê�m�Ö��.fʒ]0ehb��px�(�$��H'm�]�MZ��;y�bIdOQB�,�[�c5��Q<�`9��J�J�5�$�32�%�0���U�.�̳e��6����Qd��r���1-��u�͖�$Ш9��keGOX�Cp�;j�04@W���n7�R-�L���㭂02�e�/6b�Q��J7�yw�K������]�CV��2FZ����M�[g��7h=ƚ�����̌�Z#�:�p�-��0.:�c���2���%,f���uyn?�.3ab���a5��0H(��@6`[�(c�t�H�ڬFNe�f�q��x��Ub�&/1"A����Ө%�0��N���V��r՛@�6���f���؊����h�^����Ѕ�7f��8C�z�-�v-���V���l7oJ1��)�i"��+6��/kj�s`-K/`�n��{p���ؗ�Tb�	��m�V�d�Eh�6�D�ky��o��@V�ʺ�T����7�V�_�����ۣ��Q���At	WV¾��v�+z�}�e���#w��P�q|�ݐV��*e��#��"��eGt��;�bG,em��b��4lܬrSi\E���²B����آC7!�BN��Ǝ��m�tN��k��V�]hT�;.�&�/N�(Mxq�m�w���V�fm�&�݃d�'j�Ʈ4��7�����a�鉭4� w
���0f17^`Sjjz�+uF�b�.��
�1���5���f�Z!���	��X$
�S�� n� ��f���St�7��&�+Ϡ�Q&���f�"մ��[�Q(ƭ4�`k�z��4�=��l�3\z�F�e:`��-'�٤M�-�D��|4��w�	Zc,��-qY�T�Ʋ��ow)���7bz�(6����ހ�h�cm�W1V4j7>�e/�S�9R�fml��D]i],
�+���'��XN��4�ah�kmmjz��@�mV�f���T�!�ݥ�̶�<\	�Pe0�0��b0��K���RJUqd�]"�E3*7���V��#6nR�1L{a�Z�ݼ�V5�u&e��Tٚ�=���0J�/]*(|J�C%j��]1V�
�EL�X^i���d��q��4�v��*��l�x��Ą�F6�MQU�m��z�ƶm9�)�wor��"9�+kF	K�56��ŗ��Y �ƺt�-����
h��m6-]���ŮXV2%���!�KxG*@�yVL��f��O@�{h�@�K��f��m}�ki��U��f%D��v\��g�C+1S�jJãob
�-죸�]��Mar[潩�kҌ�buLC�dNY,���
q@����P�4��5��X��ɚݢ^7�E����5t	%��I�gZ�OYK(ދ.��RܫgE������U�.��`�OV�[KU l|�<J[� $���k`��k`{�aQ�GOU�1݃#���&�M<��By%��qm�7ׁ�o,ڕl"wJ�n!J�'�Z��b7X�F%�-�+n�b	*��A�Mbر�S̍$��`I&�5Sk3t�6�9WuL�K@f��IPu��b��4��Eӌ�I
A�ױ��+t+m
̂��)Xְ��]�p6����$��d�e�B�k	T�n3�hů^0Lͼ�+���+�N5J��`8��1#0��Owk7���SS^���T�fI��RѶ��-�゚/	.��E�m�sneD�K�%m��lJo�U�Ẕm�q�i����U�dh;n�F9��ծm�P���ePT�݆�X�own�S$H�DX�>�$��
�Sӄ������j[�C�Z���;�9T����-�:I�6S�)
"ҳzr(�`�&��~k*ֺ[��P�r�[O��K�Jɰ��;�e'�k ݣ�wqX��2k"FS5tpd��J�'���K5(}���cM�w#;Wj�h�4��^�����W�ۤ2i9�C˽�R��խ��D�.���\kX�e�Aͦ��z�Bө1��4h��n��(�%�\�f�(+4^� tJ5��R�7��N�
���%4�o%�����5�)��$�*k!�jP� ��/7V��R����!�v��;�5Z���g͂w7FF��j��zF�*SnÀ�n�X���=�P�m-k@̗�)�I�ۼnX���27�W�]C7o,Ī
�	Im�tt�˥����Dh�6��o�l�2\��A�m�)�\W팳+B��f��&�h�&��h�u�6�G�.�У9�VT��;��e�n��n��҅l��ԫ< �*`�N�HU椝�ܻ��cG^�@�9W�I��ARKR��Ndh;����e��!GjjR$a�f�˭�� Su�ܰㆱ��7F�e�"��l��:T���y{���Е����^8�yb�>��,<��pa�j;�Ωٶ@KZ���d�y��Vf:;rM�e=Ǒћ�,��pm�8������-�	Pc��gp�+:K�ǔ�\T��{*�]��-[��z�[����0��ܦ��@�v�,���6�:X^�
r�����L�oa��=ҟѨ�f�q/�&*VUbv�a�V��q��D�7Bb�.͝x�Ь.�`$V6T�z�4�+,sI%Kk���u��JK"Y[G�Z�Ln�bv�w(l�ٱQ�LVm�J��l-olf�{VXa,�kE&���w7-�u�u��Tt�u`��Ҟ�Fݭɏ77&9("C�t�A��T�5�Oq�y�4<ڎe�7�!T��d!�ؤ�8s����TY7�۴���6��魵�T�-vN�d2�e=W.�@�{"
�kQ<��Z)�����JjebA��5dԒ孢��/5�0�%�Ǝ��QQ�t7.J�h��$u��{�c0�vX�α�sj�S��%�E��X(ϑ�*Sܩ�[6V ���]_�IZ�[l�̚�L�
�шk�ƅoJ�0�ā��0H*ɳ���و����RX����9�����R�R���C��	�C����w����qQ&S��(%��絳PL*�Xl Pˉ��t���IgŬ;w�kp�h�N]ǐ���v����w6V�<u�-���פ�0���+7!�Wa�	���%�V�N&Ї���1�d�u�eH`vS��[�eL���nV�)[-k{�n��s)K7�Wd����I ����҆V�0�jZ�VV浗(����th=3Ky�i8�ջ��*&Y�1mn*ۼHeJۍCf�Dr�֤���@m���1���.�J�T�f:B�%�z��̭��K4�W���'(� MYA�݃x��*c�V^��� )K!5N]'b�XTҬ�O4<ॄ�)Q��"x�3�F����\R�Bb��t&
�gĊ����ha�z�1��Vt�:{-�Q�q���Os�a;q�%���sj�⼓/VUD��Q@�y���������cKLa�]ַO,���w.�)VB�bnMm�e̶1T'm��6=�"�[;��M��r:��Mn���˭4�я#�Gda7.T�z�Uclښ]�WQ<ũ��@4\B�A.d�H������`/)똢Z0kb:7{X���,�ݧZc!a,-�36鍻V��wf:{�BW2<��"�a�j�;�@����X�gn
6�V���*CbEM���(97&���YG]���RI��Utn:���ոv��խjV�s@J�@Y�{��^^�ޕh���Viϊ������f��^��Q@%��#ˠ���f*��d�xKFҙZ��X��va��iT��HՈ�b��3E�bC���*3m�2���ʍ"��1�Z�<� 6�k���C2
�
��5�����<L�&�[�UYقͧP�E�s4.�v����(��%��ǀ.��M�őқ[w4�4
gBm��Z��J�����Q�2�ځ�mnf���(�Qʖ7(`�c����<��3�E6�<Ma��l�((�3P)v�׹&]��+�]}w����`3�[���W�{%Z��ҼX՗X���kM2�J�3 ԃ�h����J�:V�M�j�j㹍�����7h:�V�0����[5m��M�ö$�nE�����ȶ0H�ݺ��T	6F��$h�9E[i�7���c/2e4H�����æk�?��#Q;v*,m��˶��a2��ۍc�5"�ܚ��?M���sTR�,�JX�*�ö�<"��N� I�8�V�Z�,�LP4.�%�d�*%7ke��hY���EB��QM;�ݐV7�Q�r\�#5�n���H���]�Q^�Bf�Ͷؔ۵u1���\a����B�-�of�v�xnGb�MLȕ5E�m�����nP9�Ei��1d�!�6/k0*҄ɗ�2��IV#E��v��g5�J�b"������$�@떰�AR��Qǟ( �/j��3,L4������"��m���u��oZ�x4��jYh��a��Xa�L��a�+�u���Hp{6�D[Ve��Y��)���+Rk8���Ƭ$��
�{�P�Ա�r�Rw*S[��+2bCݣa����n�09gh-Ց�-���z�.	oQ���LݥN�hj�����#��2���p"�$�x6H���|˼�M֊i���Į��0�t2��A8u+�ָ/V�?@�@r�oA�si�3v�K�1}���Z�Ν��PTY�@�w4�H,o!��mXo�=��l��^�krYJ��G]�tû�i�e��knۡ�[k"QV���蛠�s��k���x�Qzz���X�M�m<�km�B�l������d�Z)�.KRcGU�ښA�4TVɲ�V
��2�0��&,�̡��9B�Z�QĖmF�2�{x�X�ֈt�ҐVu^P�c!���T�եܛ��t�Ŕ�����Mh���j
�Z�Ӭ0��ۄӎ�d�j��ITC-^]�.��,;�ѫDĪ��J�� �ZR�i�]������jvmeʘ� j��z"����Ej�r�md%o>	��;>?(����<WYd�^���kǄ-���3. D.��חqKW
�چ�A{��F�
�T��p���Sc���t�����dn�uD;/U[8������t-/���x�V3�aӶ�DP�-`U��t/<MJ�����������b����n�Yr��Q�;�˗�6a�e����X�%�jeL
TX�lB��/[���2�t���T��S0±Kq����ܬ]�q���	7P���$��n;��&e��̫(�"�d v��5�Y��)u��͓&c�s )ĘoB�hKælR�J��-�?�埣�)��x�K6E<B��F��#Q�͍��T��Rܱ�B�L���J�n+�jK�q������k�j�L�O#�R[�+�)��S2�&f�J���\�T��IqY�Y��c�m&�;'e5D��Ո;Y��w.��8]3*��m���M=Mˬ�VrTT��Ӷ��z�xv#JU!��U��M�8ތq'��tmP���90��#m����L���@Ў�Yޭ-2��,�vqn��q���u�X��X������N�Ϟ={u�b�ƪ�����;{Z�s��10�|��,\ը���y��8r)	-C�d���U��.f�ٗ�����EW��8�8�Wx��-���r�������r�R$��4>���g���C�ܚM�@u4U��r3f�E�'��r�'�c��M	<����ھ-�>=X�j�|���U��k��n�r�t���x-U��a$X�է����`q�-� �z�FRl��7.���p���=��P4v�WoAݼlg0��w*�xz&q�����Qױ�gˎ���a[���I蜱�{���ktc���L��40�j��5�U����),u�P�M7�΅���MCXx�9����ڳyR��>
�@2j�n�����u:�������P�w�En �Nhv_J=o�'�q�]���aF���zĘ��A�\;Ҭ=���w�D>�GEہ��*Z��d���f�����3�C��ģ5#f�9Ԕ_F�#벳+��Y�X��9mZ�eL-Z���E�x����4�}�����w�>ܽ7|�ښ��7�۠W0/�͛��n�7�q*�^M�B�W��}�VA4� �N�C�4Z�:d`��I������lc�.�A��(S4:��wQ=Iub�9�N�����Q&�z�A��P�j�s�2%���7X�A�f���ub��`��>ò�\ޚrG*�;Ȭ8��j>CV �@�bͮA�F]�ݛ� �d��� '�S-[e�,cӝ�jV�dQ'�O�؏iR=��twj��*.�*�� 38����<�7��-�u;�[�4�#��փM��j���vZ����u]��S�+%,��p����r�{��bXz�z6������5�5�ƍ�]+g��G�*=H\Y���<#�M�ZKso.c
�xf��͊�ޘ1P ��]�;$��[Е^<�_alT��0���d�MM��}.R\f:4��
J ��U�<�n�L�}f���J/�z]6L쿛�ـҺ��Qy�$�0���֪Yg�֓Q���ݼ��~�[eћ\�n)1���[��_�ѹ˧Ä�j�F��0>��
�=�ڵ�MvCt���L<�a	,m6����8��G�;-ʳF��f�6O@��p�ڥ٬��%����;M��qi���5;wc��۬k�����t�'��ʺ,h�<\����5����o1��3�%.�t�)^t��-���Ǵk��z��.u�B�٣RN��ݨ�̧�@�o�����6~�ڈ�v�c�9�)+�+�� 1�%�-/�f�7�c]�}��<.n����o�l.�Ĺf�b���at���7.��X����M�E
�I��b��$��ާ<쾩tً�N�=�˲u:e�=�|x�Bjtbƅ{0�:���k:���4�s��d����=��N��U��}5KUu��q������xwRHУ�2��:��Um�ONt����y����uf���\젦��Oo�9�PXEWj��EVma]�B�Rp�ُ��k��&wl�K�q���Λ����DC�Z�7Q.Uٜ�P�w�~V���/u΄��rL��ϴ^�ل�E�u��g`U[�n�� ��%��I^9��_B�:hU�@��WdK���3�����C�X�ֻ���\����u�y]�{�^7[����4��#�����{�/T��Ad�+��_)dԛ���˃Y��/�k�ᑎ���3e��ME5�Ψ�p<���c��Π��S��6;j��=+��n��3R�X�wѽ�s��}��IΊ2r7RF�yz�19�[��&ۥ0�,(4	�؍��������fC�ʒ�Z�6A�n�5�@[�+[����NNB���]Yj<�
GAj��E&����.����+7*tӹ���,�7��n���dDb��g1+*L[L
n�*	�A�t��3+��봔�v2b�Ż��DI�ʺ�M�	���ޓ�[^�f.3��f�"�ha%�v�yƲ2]5S�9�=t�y�yǋ�k�-?i7s����S]%��!@`ɑGnQW}A���k������TF$�J�ھ��$�f-��ȐT03�4,�l�Ae�|�ш�	��i�`=�ag���Y�ˋ:N���z��`�0|>��J�6�m힣Ƕ"�R�m�����n�Ef�iѡ��M��%&=�h��g"�r���������p����H*��:�cF�ЅE��t�����V]�q�ج�j�"����;�Y����݁k7�,���SOP����EF_c.I�o�����YV��̹w���G��N�����:�H�]ڹ{C����.σ���`�ً떶�)�xc�%.���c�K4V��s�����xG8�ղA����yf�޽K�U��IQ%�2s�����i���V�����lh[�����{��ܩ�+E�oB�#��<��2^.w��1Չ7@��ޭst��N��l�:d1��%7o)#�poqѷ����K)�$wq���6�_1�e�P�Mܰ@e��3]�Z��iKU�Y:����K�ΓW���V�5Y7�m �L�4�	��ݣ0`��|�n�]}u�,��Zq���r<���x�j��n�ݻ��fp.�kr�kYĹ��m+�����' �ff��oU�XKY0}(��t�*��z*!������R���D�U���/w�©*on<���_O����2+�ى�x�ئغ�	t���ΙZ�J�ع�Wqn�5��m�u}��e佝:Y���uB��'�I�m�2��!���2�Av�:�-�1]
aҩ��C�U�Νټ�:0��t���u4^�[��q�Ƹ-��"];Xn�û+i�u	�Lo������dbf^k\�wq�a���*v7�=糺��Rd�0s�KCc��f�=c&o�=ǥ�W.�Z��Pڐ�W���ݎ�B|�!ջ\�߬�G�b*���s�����ݷX�A�c�vq��-0��|��ܢ/4�/�p��z3L0���Cwm��j�[��>j�5^Y1�O�M��l-ܶ_+;r��}�2��
yX�v��>�.ٱ;��EEKoBe�#;SJ6hr���Y�W��F�u����ӏ=z]
��8p��n��A�,V�[-�gSv�FX��ݐ���]��k)f�ɱ���A�흴^�!���z5��B���`�Ԧݷ륽f'�n�w�YJ��:�t�]���4�st�V�n�Ɋ�Yr�2��9tk�:f��k�8�2_��{�u��F��Jv̮ʖ*n=�y��v��xth�b�e�V��U���_��M��y�1OE�oN�<�Q��낯�\ֶ�F�wjƈ�8�ao�q(�Z���@f�t��K鬨��0h���x*�M�dFʰ�^^J�owsE4u�ւ��Y*p�v�u���en�j�Q��"���L���:d�V�h���u�O�N� ��؋ikn���Wܜ�NEzꋞ!����PFi%R���t�@c��� �g�]���ʼ��N�����QǢ=�u�.4$�+(�V���S;�/(H]�8��]���^f���u�X0@�P��;��uVk�RG he�����W�=m��s�G�Q�Ȯi���&����k��s%C.�Y�O6�e�J�;xu�t�j�R��W+���Q7��un�>�R�ne8�ӫmq	���k�S�r�}o&eJ�QZ:�y���Y�z2CX-q"qH��r,b�+W�?�ӳ9Q8;!E�>��\�w]�B#�Jʵ}Q*ݻ��^*�(`�㋧F����(��[է2M�Y�o4Ȗ�L�v�R$�u��2�$⨌�弇��X�������gw0Հ�J���
��8���g\�(��MWg%dP�V�������D��4�.���yN�!���HX�b��}Y�N᫦W:��k+��)\�T�n����JH��*c�3���� &��:��˧��^�f�S8���u0��3�^�u)z�,vQH�v]�p����� �;+v\U�vݫ�Tl�'q9Bě�SOoM�X��F4C�lf�H*X:A���[�7ej����M��kbD�h�P�;-i������2����ɶ�2Y�`��&��^�-��D/#�\���[[���\Znkj�3����T4��v1�֬�hJ�z �����Npȸ��4�w��Ͱ�Xe��ԙ���i}�iK��\���'�!%�{��1���ϕ����`�B�MXz��+ �d�J�I���븙�q�E�WF�G\8r�.����A�����6��X}W�N(	���M�D�*�"3�ui�/nf���R��5�]��p�~��O@�S�y�K�j"�Sf��v�*��\����V�ޗ�:d|�[�՗n���h?�3Y t���l�]aY����,���^��4U�ǉ�vP�je%]�~���_�΃��խB��5��lN��
V��r�ے�n�b��eU�ʇ�)��z�0h���u�;�M��Ϗ.'�|9���N�T�Gy{�h��'���W�sb:���X�U�O �U��	�+!�G�tfk�Ppu�zn���<i�䓒��R���%�cD��Dy���[羶�9.n{fn�]��v^Ӡ8�BZ�$;���ި�j�bVV�M��"5x�@��f�UÈ[��5��,�!P�X�;�-<�㣠�5,���@n�i�oV�{8�M�\��n�]׮=��YDvW]�$�g'�$W�����=��=��m��L%`�9`��w����O���jh���R�G&mأyWƝ0mG��r�Rb��fWף���\�$��:��lsA�.u&٦1i"���2�B�lKx��zU�u����2����/�k6g4x�_�4>���3IAU����Kd��y`��;�96�q�{e�t75�u�s��<n�f���Z�ҡĭ�Y��΅o)DWNS���\�D�)ڛۛ����5ӛ��6l��3���+��=��[Q�]�|�^,�LK�8����.��xp�_pC�v�G��/Rde7�V���.��/"뒆Q���8X����d���o��v���%3���\�ʊ��A��]_ooE"
����J�;��F%��( �o2�m�[;�gU�=�f� v�v���Vd�X9Q{���E�:��[Ü���l�xTȴg%JP��5�SfQ�SF�{���bdK�,D'u�)�x讴��÷/g1ݗ}���o�\����8�s_#<�h�ӄ��ƨ��A�6d�"�ǥ�"�{E]��E�g0Z�mg]�썮���_��,:��7�[t<�){	r���㋗V�*�:�[����yѓ}jI��p:���Sn*�J�������XVlK�������\�	3��9�1��{�m���$��x���:[Y�Rv��\��+�����*�����۾�J̛�i����C��F��Ė���E�,�ܙ}|�� ���vw�k�F�=�K�/�,w`<L��6u�=�,��1:d�'7�]�p�KI�����-pt{���,4�ky� osEfp²���5[oeof_FC�ݮ���k�0u�e�ǀ-�VU�w���)�V�C��؁-<��lq�"+�v�� ���+�r��Kuo\/�VWu�.5}v��:�ְ�ƍVF�u.Si���p�:Kq�5}�-���T�g1ʕ-����;�[]ƬfR��t�b"�֖+N�wH�\�*${h�  r46ݓQ�{}�)�[�lT��p"��ְ�ԙ�w:hDY}�)���gMI)ʾo�;�Р�oP�Q���3jяDo�A9�iL�����ռ7c��on`����i۩M�ݖ����R�p�$
��T�W��	+����ȓogv�* ��C�Fewf7B]��Et��YIj;Ss'��e��LWQ��O`t���&�Q�D�'��@M`	�[�R��<��7��s/+zYu�VZKX�@�])͠�е7]���������V�@ms���r���Yuΰ3���>D�6�˳� ����h��Ve���Eg(�&�).�4����TKV�w�S:'����/��}�N�b���t��tC6l��j�)[��ޤ@p��n*����v���飣��GlTj��
�p� W|ܤ��7]����1�A��pvq;��υ��uY���v��R��%9�2.�2N��-�r��,(^ Sr�ϕi�u�t��!���4ո�G�b���
ޮoQ]Y7��U�8�Т)ҹ���:�'c��1��Y�)`Ep���e�OB��0�w^֨��oy��X뻂dZiz��m��P(]߫�������FM���v)��%%S�7/y>�G��Zf�����K�m0�����(��<�:�鬍��1�2�b�:��\J,�ѡ�0)��Ǧ3
͇zK�Z&Z=�XM�R͒Ź�u�+68pD�^���դ���KE���;�C���$��S�N���>]&��s�ҍ�7 ����E̕��z�<ζ�K��ui�tƕ����Ճ���֮4�[I(�9�R7��h:�*�j�S�p��TB��'^�P\ҫ�o
��\f搩����՚L�v_"�p�J��brބ����K�ŭ�Վ7
�Af��� Zz��7�U��g#:��������·'jT�p�6o�]J�x�H��9Թ������w|imn�+���.��}m>�ᶵi�,t�v'_E5ۮ�w�j��N�܈J�}� b�����^��+	�T�[�V�>Lk������3;9�9�9���/����p�v.��#2WVZ;o���.UѸ�[7�r&���2���f�Z�@�ڂ���}���B		���$�{��>:yX���W���2h/�ܚ4���D�nN������SCk.��=��Z�Zb
�P̑J/a\�1u�hS��*��/�,�6w4*ttΆ�[6���h�0��j]��V(M�eu���j[5�C�����"xlD��*���Lhª��]�s�3̜��S���y�;Eu�Ri:\���X{q2�J�)9+�J�F�$��Qޝ=+�4e�[�-bh��-�{��C*F��n�w9������6�M������_�;*��?�:˨�CF��S�3!��G$c�W[LT��փ|�u��B��/�*Xz�Jl8ˣI� =�hS�<����G��Z;N�$�p���V7SwD�W�,u��Ů螊�e���pm�jJ�9�z�
�����]tI��9� ��M���l�'�iˮ��(i �]�����٭��C�wG�*��x3��#��]`ǲìg�݀�y�&�v֬`/�%:�v��;�3DJ�`�T^�}�*�Z��!�[(�9��^s�� q��k���:��i8�k�j�8���kSu;v����}�h��b�2��Ē�?cD�I����O<��rLw�gt�;�� ���s���h���φ�4���j�.�܃d�2�g��e�Úy�9&���gS���GX0�J��9PqN�-XY�g_i.����L�{Z���p�;�����B<��Zu���ƺ�+���n��l
�Z]vأ/>n%ս�b=�e8U�V:�d��1r�A�B딧�wz��
E�n[f�ZU쐻U�86�۲'*s����Y��W8�����;�'\X���00���}��G;#��{��[BvtE�\b��hŐ��^��F��;
��op�q9[R�і&�z�]���͂�W�cU���gk��P`�V�w���&3���X��vG�7�e�����F�������C��ŨR�����x(Ow_��҃�f[|:Z��N��˶���$��3ۆ^�4�ƚWz��6!���ǜ;Pº���K��A�%s�x�Sw%��0j!�d|_;{�)!zI�7]��(cVܸ�5��$�qU��֫L�3� �k�fv��4���o
�v�Q���։�u�Gg$QW[�틲)f�j��Ž�
���Z��+q�;��f�k�8��"ї;�ʛɉ���N�M[W�oq��g������ҖEӧJ�x%'l+�h���F�+`!��g�Q�|w��6AW��I��o�ŧ��<}c���D��}j�f�8��͆U���|C��sw1�w����/���w.�' 5�%�B>
��J��eM��N��L: X'NiVTP���h/gj�*�4DGkd�=�ٺZ�Ѽ�)�m�����b܊�.u���WJ��77��{=W�f����(@��,� ��.�m�[#9��u;CQ�ݿ�Y�|9i�a�E�	��ܢ��]�ê���4��:?���ͻS��-�@;r�U�`����5&0����u#����]�QLv�F��<�p���Ǽڵ2���MX��J����C]�Pk(�̆�"v˔7���q�٤�F!&�>y��
k}�gͫ�_1����C3�m[��
�N�d�|[wB�1��=4��Z�Ν[�Әj�s�U&k��WY�%������y����"��DvUB�7����PӒ��{oLֲb��/�V���{˄���+�����r�l���f�5�j������Z7J���1����)�y�ZZ��U�@�|�}r����oumn_\�C�<%=��F��&��#��:��ϹX�v�w����M�ŦT`!P�Jf�.��a�J.n�'�������_>+w:�S��3j+�8h՚ �p�Vo���v7y$�޼�@��=��DRU�!KP;�zb���۸�
��@:�oS�2�,�C\FeuX��G�I8�]�'��WVe��k�\�D���z�J��No����z7�/����d��ni��`��.��;�˴�rX�����U���U��f��\����2��&��kxlm0�i����D��9Y���}2��}xT\���j�����*�I������K�6`��\ugxS�lw�8a_h��:N�k#�Cl�RV+}J��;���=������}�Ew��Ѫ��t�ݘ.X��6�w&������e���X#k��4�oul������b���YΫ����A�P�S��fZw�WN_jj�c�K��mYv��8��7Z���y1�};�YǕśV�-,�&G���χf���f%a�CYlvv�@��{V�|~eiU�-PYJ�L��(������Y8J�Ͱ���En��*�QEJ�Xr�=Hn�-}��2[ڒ�ӧ9��OGPi�
z X�P�U&�v�����x��Ic��E�xU��+B������!��+S�f`��ˡ`��y�.��6�+ݬ��x���3�H�k��<V��vl��U��[8	���,�^*U�my�M�s��x�w���r�v�q��C]E�ԥ���U���<sh���"��u`�Lp��T��3
 zeH2b�j+&� ��%�m�Z���+�6�X}�w[�{A!�x�u7x·7χ.�+�p���1פ�U��[�Ǝ�V�o��Al�`m3u�7��ۮ���ʩ�e�;4�^Y�,VeZ�1mY�ժZ�vӽ�� 5V��2]�9�_2��Y���`ޖ���5Eҷ���u1jT��}���PO�����(9����E��&�B��+��՝�j���Y���PnU�d�ݟ8�Yo��闙ue"7�mdgf�W eH;�Ut��$a�ʝo�i�H<���i���pj��s�L��熸n��OI��R�s����:)쓨һ9��m�q+/Xٜ��DӔ���pV�pa��x�j'�*��1V����w� ����(����Me]kJ�u}u$;���H��Wo���	��N}Yz�u�I���-:��a�'�b���+�L}�N�b�j���;����1�Pg��wNKJ����;'7we!(^ҩ�����+pR��cs#�q|:!�CszQ�'U��(��s��3{y I���a�h��K厸��d���������gc�G���tk���¬�����"_>��dc��W3>�ή{G6!��1��װY�(�սc�kq ��h�vdO���x�(x���F��}0��5��A�6� �hr��Zn,[/�v�l��U�(J]�f.�Kw�+�X:��%O���k��y]�����U{)��j�&b��z���{2ڽ��#���I:�`�1Zl8�7��������χc�c�wz����@ޞ�tR�h(-��q��_!�d�3���r|Z=f��A�y���:;9]^�u.����GS�x��s{t���LC�N�we)�����m�0䨭mX��x�8�w�5�w�a�$�uNC��EX���B��ܠ>�v%�bј١ ��]���e���:+����[�,P\��Y��o)�y�8�XƉ)���S�NՎ�b��ɼkԟV��-��jv�jB�,��tI�����qLB p�+g6��wa��n���ȵ�����h ���]�]^�}9˺\-�4�憅z�r��_-2���w%�(Z]��ϳ�^0Fno p/��C�V���C+]t55�Fiɍ<�R����]h)e�UܳK�m��+���E��p{ڹ�\���Y�Ue*R��X2��]��J _�Y��q5\�ͫ�ɗ8]]��ָ�ʏ�a��<���{W%<���ʸ�1j���=<`C�);�1�!�L�Ջn��|;�|�����N�[�����V�i�#$n^-��;fv�#H��=CLԔ�6ԝ ���kK�=9�f��zi�f- sB��-�̜˱��q�О��!;�5E���LfeԢ���-uL����<���w���W�O��ֺ��lnY��=|✲��8��r�J���ԡ��y�-�ݱ�J�v�AX�*ժ�P��qh�S��s�}8<����lP�3s+L6WҨ��ب�� �b�G���ZB��_lJ+�Qq]@�0�A�kK��k�.�vnP��L�#����Y�Eld�@;���5�sbŶ+�w[w�[Z��3rb��Ũ�����ʺَ�Ǭ�d�)+ۉ����k%��uI)b%#�kE%�����X�b�j�*[W����eA�׵�n�b`��k�ఎ�kC[D�5�X9}�.��h��(�;�����V&��eU�t�)+�]o0
9Sl�Y��ibl��a�@nP� ���IImc��u�E�\�m��gJ���T��t­�X��/��<��gU���w-]�2#g�c4]aʼd� tFZ�9���t���7�G����В�ꙙY��浽�y��y3U��m�s�f�ֈ1;�&�cEJ�z���AۗoOf�bS�2�ӑIe��*��s��.��;T��fCx��|����X;�]KY2Y���Y�k�r��[.��P�j<�h��KOr90�]��Z�YX��*ӻ��˷v�+b���F;���R�LV��K���|������n'oDua��vض3���,����nb$\��\�or�ǶJ�~̮��*D�i��%��qاWC9`v/:;���J�`\�6�����Y�m���V
�zt�s+�K�i0��v���ZBK	��4ֳ]�����>�#YaqR��Rn]*wk_*��ޥ�����VL��7/r��v�ɧ�\J-Vŉ����l_q�;.c��`qb�땚����kR�X�m����� n����:������-��P%���Ju7�&�!�E�6�!t�.����[��o%Fm���=*��.H����k��g]#���h���(Y�\��o�s�w(��{��`����9�(p����Qv��y��Ѽѹ�(9��垜i�B�4�.�;%�,�Os�H�m[M	P�Ŵ2QɬS.l�g8�����Z"�A��`��o#Rֶul/�ew-3>l�/���k&�����J��r�W>v#�)6��v�٥��Y��2�y����m���E�"f˰N3�'�v�O��eHx� #3�[�GV�9vv�h�j�$��@Нԗbk"���X G���Agdj��t�}|��=৮��FpS����f�lR	 2
�ٕҬ1u[TH��Keޅ�f��M�1��_˚��@u�^ͼSib'P�O���Do}*���e�fwG�w)�Z��9[f�:Y{��k��K勰ژ �Le���2�0�D�H;x�٧Q��U�nn���1`_3):�����x t��	�Z/��c������AQ��^v�8��>vO'�����B�%�`Ȣ���*�$�-w�;�	�졭�ʺ[������K�j�Wd��]�DwǤ�����4,�z��X���+V��s�k�c�)�zV�Lk�Ȃ�����۝����J��}ٷ�͝83Z �sX�E�[���\�A��H��1�R�]��~�[d��Һ�.[h����NV�Q�GV�7j�4�v��:{�G�:ڱ��,=l&��$�btTW���sa���f�̠z_<u;�I̼V�s�������XV�����t��FX��5�C����m�D�U�C�c �U��s%m�Cm�<{��!�[3'&+�BV�#VkP!>\GMf�I��%;Zet�F�e�0ȩ�s���nJ���M4��v�E�˒w�H)�1��`��6�PB�u,���u�����۷��m��n����y��)�2&��;�h��C�ٝx-z�G��՚b$)	�V��T��!l��fudQʹu��\u�@t��i�lCh�|\�:oE3$ ���_$ ��2�N���;zL<����9;'��)w}���t󶸜fb	J����s����J�wh�|�z��*:����wY�%���ɻJ��_fP�&s�ml�&д��fb-	�i�̭C�ľm�Z+��hY���Uf��.�fD���xj����9��mn��:=�]Ƒ%�<.��\i���n�G��k��	}����Vwd�@1�N�U��՗|�H�;�A�J���$��� ��-d�e��i���Ɲ:����E��x�i�G1qX�[.�Ԁc�����T�:����*5#��	�����E6:��_^�h@uK�M^p\�3pp�n�i:Ub�)��V�<�\�ʓ�V�{X�:��{�ˋ�/����u�0Ly�u��k�y��_+Nl�*�G��Q�[}%��z'wW�3��*} ;hkYy;t��εێ�=[��R�'�m�-��`��J�$�Ow6)��ou�wb��R���3�10��WVDe̠�[Ӿ�����֌�Ɇ�M�����늹�v�o7���X��ܔ�Z#�֥�{)����ǌ|+���%����u>�3��Fs�;R��*x��2�ֲF��s�Sz��錍]��ټu!c�uvA�k*�e�g]��WG�M5HҴ�Z���zr�[�l�n��3+�����Stc3�1��1�p7ǂ�yݓJ&�p�7N}'q.�RJ��g�v����6�u��>�V�;IӹC@wv)�LU1EK������L6�)��}�v����[�B�\"��i�M���|z�ǒ���k"G/2�nv�Xi
хՒ�:$Ă��<�G.ܨ��y�p7Fd���r��n�63ە������N޹���n��mwD��/���1��U�����A[�!�R����pGGT���Y�����xx{��t(Ĺ��^��-0*=����oPWz�uu�ƌ\��E<�՚hg�L��n���,��v�[�͝㋻>�k�x�*�j�x��r;c��GOY��E}[��Nu<��=��(�*bK����ݑ���xՇ`Ks��YĲ]^A�\���E��pQ2̗V�Ew'L��f��{bi�w�d�N�%LZ�����[�EG��哯�y�I��Ҭ;Q7�d�j�
W�r�M�	����p���{�Q/C-dyq4M@_(2y�]Z�FN�J9;��@����cεvȮ�5&NH���y�d���}�����WN�ք��V̅��fX�^U�˦����ϙ&����y�>>2U�Y��x�s>�e�ՂrE�Z]�r��'���Ŕ��*[��;�T�ؠ���)��K��Y�7Y�^<���)�b�� [��,�uO����v�Í3ۖ ]-�����t���K��:�[���.��Q����j٦�K�/(�Ak���/��=�hD���uN�t�Pq��m1�H�ʇqyҢ&�j����^���\���#�5��9��/�\���	}�j��+��N##+6���N�-�=L��|��K7$�T۳\Z��5_��o�ƻ)�l�bY�k&����M�����\���wP��;ա��t��������"�p���˝;�㪶���7J0�Bij�w]۾�㎀4�$> �����1)R��Zұb��UG2����llWk�m�e*�jV��T�-mmj�3,�i�fJZ��ڃTmkE��m*1���i�\J�Z��*�5��ڶTiZ�Qh����"�J�j����cJ�h�-,�U��Dk(�E(�kjX�-����5��
�.)�-T���ZV�+[j�[F֨�Z���e�h�U�ie���kj�mB��Z�,m�F�UV�T���iKk*,JU��j+m�m�[
���F*�[XЭ��Y[kVV��������,j��(�Q*UJ��V�iJƔj���E��%���Q�کR��Z�-�h��֩Xڵ�imeJ�
��#EZ5R��¶��UZ�J���X����E-R�%��KJ�ZR�JZZ��KB�Z-R�*�������QZ�F�iX%�Pm����(Z��)E�Z�Ֆ[#�%+U,DR�-mlaX�ʔKKKb�b��Z,m�D�����Ѵ�%*%F"ն�mQ+V����l����������iJִU�[*6�j[A�^z.�s��~�2��K:����j�m�_���b�_NWL��\�'q����(A8��hZ�2�;��;��w3����5շ"|�5�#�eU�4�(�xD�;չv�	OFǕ�
����Z���k3I����疞qxQ_|�z�6/h)\`�^�ҍ`�J�z6�'�4ݽ�>�dͅ���CV����G��8k�:���;�8,+2(���E(�6e�ы���Nrt$�J9w^;#�w֡��|��B����6u\^�|g���n����]�q w���'���!b�XZj{��Q�<�1x�X*SU�J����Nݎ���m~M�}�ɱ2�����x�cP��4���i�����E�n.,p�y���#S{=�*��ka���&�t��P�d��AE]8S4&�j^l��"�hT��'�|��+�L�a�GA���u^��]��~�e�٤'B��q�J��]�]S���ygw9=Ǣ�f�h�E��scH��,��s�Ǜ�e��p�aU�5c0J�з���!j��PX\�;�(O����;A�_,�	H�/��4��#��D��l�Z��x�<����"[�ݾl/�o�.�Є�}S�2,]���9mq�q��yV�ӡ1��Ok�;�^�7^�MV�侻�Pq�|^S�c�՝W�WN�����v��=Y�/�Mޤ瀘�QQ�wk8g[��w7O6;��O�a�ѼC��z�}�ha�sXĝz�����������=�=�4>���3;��91((`:h\f)����!�9'V��k�OQ��>�'(m�-<�}��[Gةp���lP(2�`�JY}[�'n<|�N)�U�'�����+��������(֌A{j]:8&v��A!9W�jz�T"��j�;�ݴkbq�㾧x��u�@nD�;�1�W��|A%f�����|/�a�
LX�y�a4�0��.�^d��ç9#�	��O�8|��!�;^��B�B"�b�J�x�� �R��֠��_�����XZlotf�w�c���s�}#�W�����Ǽ)֭�W��L�v?��ξu�4b�%���`; �*��;��l���Brb�W�Q0҉���w���=s��m�����l]�:�H��h�>��!ڲ:��'��=,�m�ȑ�wX(]�S�zr�V�[�~�dAD�[��U�5\i��A�eŎ�U�����t-����3����;uv�v[�}E��[���1u`B��ߐ$�!Xye��g5p��U@x��ek�ČCMw�'d��f�c�����i��WC�ڼ��+z�Q�ګ�&���{�Wn�FS	N��f�y��. �}���p�s{,�xQ�c^s#y���<������7K�Z� ����C��dH�v�*��)ഒМӍ݋�巻��6w53
a0���1��s�-����AZA*�Eb����r.#{�����G���;����2�KM���D:{EA���̖���}44j��+Z��b�k�\��2Zi���%+G�$>Dl����,�,U�!��r
��Q���"b�G�A�3_�����N	�z�8�P�z�z��>�t��B��Q»q��ʼ�ȇ�R�
�W6���`�����E_A�4��S)��CMz0.���ʱ�z-NAn��^�{b��g,�d�������&��
ŝ�lU��H��`��
�k`��^ד!���3Z�9���������0���D�#dz���:�m��tlhC<V�=��f*pᝧ=��k.C�F��_�_�j2V��L�FR�UtIlqU��6 �R��݂��a�n��e��z�Z�bv�+�
�/N���
������kR�:S��C� j���h���kv��sƘ�M�}��c�����������^:�μޮv�>�D�[:�>�T>|�mr��|�.�����	-�25�V��7 N��9D�U����NT��MP\�:�Y���fwIC��IB1��L��j ���p�����+;l�͛a'�vWT`�wHyh����(>�[2�ޣ�e�x/|��OB������`PC���/�p�Pj��d��7K�S�?w�]q�%hSElŧ�n'��K��c����/�>p��r�xS$!V��Fb�B¸���;��y5[�]���)�W��L�{�gۼ�P���U�̀�Ui����P1?.(��܈+�����A�#��9/Ie������D�c���ϫ��Wυl^V+#��i��Ei/��m^�ܨԝ�Ӛ��ɦt_M�>�NӸ�|�B�$p����ך�� vX��إ�ɂb+���r7�XޯMG@���7ݦㅮ?I��fE���4C� �~��P�b���o������c�q[�K�;+e|���^��P_�Ն|��Lu��e�2��x�Z�9��;{�Z�'�=rjFAw�NC f�6��x�A�������Q�+2���q�����sP}���Kc�P�]���I7���W�(�z/�iݔ!��C����3xC�Gfg zb1]������.��υ T٘�P�8bx��e�'N�xh���¼:��Þ�G��F6`�V0�/c��n���x�����\��d.p�\x-�Ŋ��hi�ΕLRwv��8.����z!Vf,��G�4:Υq�z7+-�W]�ԍ�򾅭�94��~����Ն+�+J�W�c�&�4Q�W�5B5Hԩ��@�Yqn�,��J����D�R8�Lt��бmKp�w��MOf�R�X<=S���JytP/���Xd��8�D��|�
2����ig�^����ΫO�(xR�Ǐ�9���(�D��b��;/�Ȥq�/M,������q����:!Uh�j�z��T|]t5��{���ͩ��K�C�㹲������و3>^y=��E�}��A���/L|h�S��䇲�H��,���<S�.�mX�9W}����޿�-5hP�>!R8��8k��@4�w�=������^�-�R}i3�=�W���N��:����ܕ�{�P���|��BAZbGA�u��j#.��������<���ױ@-UaCS�����)U`Ύ�z)�C\�.6nf窝����e��3w٩]��0��P����AGl�K|��@L�>��bj(e\�J׳.4g��u%��d�ܩS`۽SR��v��2
[f��g*�������j��wc�T��8�f���wc�����X>���#���u;e���qb �d9(+G��[��g}5i9��N:�}a
v;��.CBw[�T˻�u���f�����{W׽�����})�-��� �l�N}X��?wT@@�D�>MP;�جv��m��\0���{�&���׃0_�XURs�/��9X�Q�0x};^"n��>�����&cv��m��a�28G����"E�]j�x/��󨗼p|%���~�{�/mc�끳`��u�����jj������/�V�a�R&Y���x�����43~�g�w���f];Y�Aύ���z^�Ŝ;5�I��]dI���h���8K�:�[˜v���C�K��$nJ�#����˾g��!�*;�2s�����q�]�����d�0z��<y;���������DR�_A�;q��jb2Kt5΋�N�:�s�ʁ)�<��B�%`4c[A�E�NW�S��煹�$���n���K��E�����BQ#�P�ta+0�u�����VI.5f�iW��8�>��+a\�2v��ۧ�>hqF}}��`=��1J�����1�7b�d�G#����RIv��;�_��r�̮��T�)g�.��݂�x��̿ojQ��RVu�:`c�zٖ���>�����u_Q�P�ik���CA��m���z�����t���tnͺG����ǋ��j�v��۪�ޛq�9اqSP�R��Տ�/�oG�v��&}�酂G���*��p�h�1jtٍ���q+e��"�B� �$�8.vW⯡˭��>������������=�6��9��)�8a�����q?[���b120Z����P�/>��mJ��׷���Z�����ޏ Za	�z:c�X���QPoqc��UauD7��(r�bYN�.�K�˫�;.�`�B얪@�,."����|ߍ�2/�Rs)ܾ�6t\�q��ppm���LDr�3	�6@a�5�4fI�B(E l����������[��w��9i�V��Q��!��]6�M�
DC����#�������"��o�f/�������]O&��dy��[Gw�v����ձ��!:�2�"�u|f��B�Xˍ.���'�7w�҇�^W5[��ma�11����Q�ڙW�?
,V*]�~%��ø�=���}���jH���y�[^I��)=����A��V���g�܁��e�Y�Xf�K��k���<�V"����q����A�H�Q�2��A���Ka�B�K�Ց.����wV�%��l�̊�sr�$]�ѕ�CS�Wwf.F�f�ك���z§���Cpqֱ^� @�UÔ���ħ˵^�e��Á޺�ޘXȻ~�Y\G��U�}��e�����ؾ軽>�߮���y����w�oV�|����D�R��6��m��)ѱ
��\�F.�}ļӵ�w����Zw��:�
�<h�H2V�ɘ��ϒҰ	}� ���:���8���0��]p3E-��5�Lݬ"��qdW��
���;��
������kR�H�L_}C���2�x�g�<���{I�97���h�"������!F�ɞ���o�"C04�+;l\bꂎ�jh��* B����q�W��%B�@�����9�C�`��g��+�����4=�5�]�}����2�3qB�,�!�K�S���R�ʋnZ�WG[��D��i�Fn�LY7��hlk���#Z��@��R%pzE���w�P11��*܊��}~��VL��Ew��Tm�v�Oy2��U!�� -3���P�E z$^/����|��v�f�:�Z�pb�:������2t�^t�x������Np�}��V~Tu�*�}�n��fa������s�H��
m�-�q�v�5]�ŧ%#���ǫ��M��#�H,ڎgp���F {b_vu��c��r͐��l�5����ڴ���i�s��M;Ӻ�L����܍��D+73���#��3Y�Sk�e<c
��Wʯ%�8�2}8Y�Ƚ���������"�o~��#������d
�꼉V���"�lgT>x�X�g(]�6���F��P^�a�\�T��Y��Ev8�Y����vS������8X��H�/���C��
��q�9W9Y�S�=�S�S(���n/z���v:/f����>la`5�$����o���Dz����QN�uձ�)�ZZ��s��`2�"��+�Z�ΚS�����b���FA���6z����D�34�ޒ�l���@��,�N��r��\_��'c9#�+�L�R8�>�Uge�{[Ts��ֵ;�+��<0C��Q4��[�r�X٥=z����p�̕�����L%EU�$���<��Yc:6��8���T��J�
��s�6�X��8�̎�ȷ<���ٕj�of����װ�U�w(�����X���l�>�y�����������c$�7�r;�l���ETz��v*u��<��q1����=M�;_)\||�4-	�����ZG�čͬ`��p�O����d�ª�s�9����j���������;���M��m�F��i߽W��������t�+�moV'��^_
�j��KJ��w�ڮ�gH�UI���M���w�u1�"�������{�{�2��d�����|��;�}�zzH�*��$q+�(s�:��A�}C�#^ާw�:p;�sh��ZA�##T��6
�J:|���ܕ�Y����(H+L�gU��`C;^/x�s��=}�Ĕ���uz�!�V5;��q���V�J�[BF�����Y0�pke�w]q��|J��U���������q�Q�wS�#�>��S��o��IN�|и���#X4:F����� �Z�o�E�=�!"%�8�r�>�R����R�W{�¥"�`&���N���o�
Nv/�x=���X�ѱ�г�n.�\b��vQ�a�L2ҽ�\��N�'��@�?70V5_5dWy�0лD��#\��O6��j.�n1�ι�b/n�����_P[&�ӛ5��1�dpKև��kN\U���G�}�-d����H@>�P��Q��ؿ����}Cfh��ؒ9��
'��[�֎%����ܖ�v�u�rE�� qLe-<���=����bD7��|0�{ݲ�|���v5W㋚p:��Q]:�����\�K##�H��
����'�M�I�+���hX���z�b.Q�2O+�ʼ�6��Ҏ֬���J�Юk.r�Qݖ�����J+�!{�.����wHU>(h�0Z�W�:���4tͭx���$�>�X��9��i�;8wܒKα��M�zQ�`���4]�e�x����U��K1�]u�%:Q9�~�1aѢ��wM	0�j���jM�})��r}t�K����c��c��kY:�9�0�<���ӵp�/�Mo�Rz�/(UЗZ��W;�]�W+/-�����^8`�I��ɾ�]��ݗ�=N��x�(� 	�\��ۃ�������[�c�X���=3�{�j�,s����m�/�S��&ѕs-��
�3k�oue݃T�k�	���"L����3c��uט:����yb��t�9�Զ�n:�|f`q�%�u�X���k\q��Ӻ�3�R��L]n�ˡJ�]�����-A�֥c���K^�q��ukh;�J�5/���iͽ���'��b�t���/�[�����mwF\u%��r��͈f ��dΛM=�z*�M��+pU�ST*vQ��<�ҵ��V�s*�vV�=wb�Ҧ�vM��#g@�xU�L붂c�*�vSU�Y�j!;U�c>���2(�#�h��"��)q��:�=�JAn��f��E���ؚ�yV����D#�M���#]�h;o̢Kw�vܸ��l&^ʓ/��x�nĶ|Uqč�]d�j.R�\l3�d����9���x55�ѻ�/6q�(�A��ɂ��<{
3:>ղh���4!]l�r�h�ǻ�Ȳ�E8�veL���suj�܍�铢��H�Yp�*�9�����W#��G�j�1JǄ����	f}g]��w�VJ
��4����,(��hB,RG7v� 1+h������&�Q��5��u��2(�a��ͳ6G��=f�.��G@�4�H�wn������F�FJ�NV_-����byLT��K��C^��c�uJg^�"<}��E�����h�b�k��w:j�pӝ9���5��eP�U$V�\o��/����9x�8/:v�2Wk���cZ8P�0���a�ۉ!l����r�u���!����0�Tc�l����8_\w�~˜�˹5RD�ȡ\quv`�����?f��XJ��X�A�Vj��T��o�U�>��a9��yΝ3Q���p� ::Y��n��.�#�q�tv��X:ᬹo�Q�U�3(��L�^��P��iҥI��G"W���oP�R�,Z���E9@�W'v�zn��ѩ�h�ە|���R��
�ʳZys�h|���S�9a �2W*e�Sx>&q�\�Ѿ{"���o+������z��N�%�����w���R���֖���*�h�і�ijңUhZ�YF���)m��eE�������ҕ�AFQ�h���DU����Ъ��V��j��kb�[TV�-�UE�ED��[h%�V�B�"6�X��)Rږ�P���֩YQcb�(T�,AYm� ԱQE*�KZ6��Z�5Eb��T��Jĭ-��6�c
��b�m�
���+P��m�Z�`���R�6�ժҔ�6��EjZ%��eJ�ԥZ�P����b�ԥV�R((ҵlUDkR*���E �Z���j-����,(��ԱDB�E-�mJ��%+K-mjTTc-�֣m�iF*#j����"��ءB����aX"�J2��0�D�h���imkeV��e�j��գF�E�"�6�E��FҨ����m��Rҕ�m�V��e�+RшԭZ4�m[j
Q�X�YKmm��F�PZ�X"�i[aEH�ډl���+R�d-YeaEUTD���b%J�ʂZQ(ȣiU�)V�V(6��*�B�mTF#mb�A��=�����az����.�)z�W-�]]���G:�\�Y���R��M[F���׎v{$�F.{�RY�y��cݥ�o3����_1�z��t�D���>�X$R�C�"݄���v�7'Гv��^��JnVJ�P'R=�G�*��z�i�����ypp�x��mD��YY�{�ֹ�ݞ ��z�$��4D6��LjU� ��CJ��_}|�B�eND��;�R�e�)ZP�t[_{�/N������H��C��=�!������*`�b�9���ߡ�Û7�nB�;[����̫t�A��n��n�I^	�[UU���%G{��nl�#�i�W�PՄO�U��`�Ӥ���~�����aU��GZ�eu�ݢ������k�����4ʖ����b122��'��P�%��7~�;רIx-s��ѹ<R�W�e+�8�D��g����U�Ś�ʇA��k� �u�� ՛�'{�w}�O+E�P� ͫӋ�Z� ����U�(,1��S���_��M`�ҹ�s�f*:IZ�є:P��G��H�U8*��V�J�QX�dw�G٠�7kΒ묄Ȃ���/���i���`�����o`�@%���t��t� ��9x3���ʲ0S�������\O�"T=[�']\E��B�U��ё�`њ�P�Ő�S�8��9�͇����qpE�c��)�<d������7��0~��Ɵ�P�3�v�������>ْ���
�%�z�ǋ�N�O�/\�q�K�x��\�����\KD�
�
�՚������u�D']���\��d���g�@�}&l$4_��LǏ=�Xj�����@�t�m�h�ЙW�+�lGOOb�W%���)�x�IL�O��5'յ�/���$��-�@�Aʼ��jg�ݛ���V,�ԁ졳h��^�t�`h��lI�ڑQn�OA�y5�}hS������[�CF��\�����=�㽌�bzT>_;�|��d{��_D8����Y�F0A�8d^��3�i\��ѥv�k����|��%b��GM�|���A_ms�A�o�XöE/\����W�g���z����Jk�
������r���c]$aZ���q�+m?r?:�v]�<�R�3%8���܋�G�X2r[��(<�fT=Ufm���٬qL�\v��C"u�Iؓ0�x��_���(x�|u������ǖ�6k{)�z߻�{/;DGŪ>�J\��.�\��o	y(>&��=��j����d'��Nӑ�����[�L���o+!
,&�>R����f��vŝ��L���C��R��m��3\O�	���#���V� M��'t�i�+M�-�=�t���;��JH�2�qB�Q�E7�p�F�-�"�q��b�V�=�g0��4ջ��9���;�[d`�-SɡT�M|
�	6��U�ˊ.-�<k��"��R�g��@؜~[q
��0�.L= T�V��=�k�+8�)v�Gp�d���Λ�KSsh? �;��/j��=���������QEzi�\\�б�F딆=�ˬ^���W�0��*ٵ�X�=���龥�����c�?{XĄ�Xݽ	�u�~���d�;BDO�g�|��.��;9W}��?!���~�ެ0��4g];sxv���.sٵ��ɢ�-�DlW�
�H�*�9�0�ر�6��z��2C ��s���l�4Y�Z�bfZ���^�Ԓņ���������4�O?a��q��^���P��^��"�"�O��-h�M)���V+�ءq�@ڛsƠ5�e/*�A��6���+���|����t�"8����[��O�D���rd�¨�"s�I�~v{��쫨2��(Ƶ��u5�ނf��*�n��+�:��@���q�3�ܮ���q<�.�����YTgS�۔�%3���!4{MN�S���/��)
k������[a���	��*t5��_1?��n"�����p��zv���R����*�O��*h��F��-��+7r5�
�W�ύ'7vr����\t�4!)��T����B��(�8:mJ��V��ndK�C��g�������g�����C��/ �_��\|��u,_�����\O��e�Q��Oُ�ȿ5�3�؆�?s��a���f������B��?���6����pp�e`�Ab'�|�N�ӯ�/g�8�.������㢮Fs�5#�W�>p�'W���^�9�}S	oo�Nh=��9V�b�B�x��F�W�Q�ȧ���ٽ,d����*Q �6Cݷ��SHԔ�Vڼi]GNd�f��x��S�& R���+�"z����n��w�U�pc���8�2��Az�����^<���cQr�o:N����Q�1R�7q����ɰi�7�:�zg�G2�{-�}�]��Ǝ#X<5��ju~~:�:S�b~4�r�"�֖��������:��F��7 �h	:�'��bo�B�h���v	�E]��c���!Ҽ�^T�DXl��Jt�cX�2�z/\|�U�p�1&r���z��<�\�Y<b�4�t�9{�͜�]�Ӈf:���Μ���MÝ-��L����bVn�1�u�*��6��-�4���t�쌢v����8�T3���w������$�Y޵����7]3	d�����+ڝ{�<-*A������,®��'e�b�;����uX�sh�"��6v}Al�zsf��G&KC�-��A���T�ysg��`jR�	�A��B�K� �Fl��~V�b��0隅��K�(�y�ՖX��r��b�D�o11T������X<:���[�3��܂�:��E�2�;�;׊�ijt�ޖU��Ο�z1	[�E�Q�7S����b�PeB�"����E������izx��@���%Ї޵�G�*�*���
�� �t�܄�]�f�^×���q8X���I��47�I�#�!��{�� ���J��z����Rd̛�W�c�s;���g���)�ػ�ӧ�G �[t�$n.�Z��+ؽA!Z!V�Q��6Ь���bm�>rTGK�^��E)�dڐ��v�Ǘ�N�e9f�xZF�M��đs���@�.�����3��y���P�l��x_˹ԃ�����ŋ�[����}�V�x��6����yI��ۣ}[p��皹��c��q�@Uu3i�h5dFMefߐ<W_+#S�� ;K9,Kc��%�n�;����>-O*J�B(^��]\F7P؉��[��YY�ٮe���f�F��0�iyB2�pʭ�S1x�����T�@k���>�y�4���J����m֠�+ǎ�!u���'��$�>⟫
UX>sP��>�>mT>5^/�?	[G_)�j��fsY���f�8N��
p�<ڰ|'d�_HŮ"����7�f�E���O�Úu��g�����g�,��`�d���(�y?N�i�����i��;^��s��0r�sz+ɽjȂ�jρ�Z�L�^�����c��xI_bS���ME{=ˇ�х��?N��]f���x�S�f�4T�߼pX��`φ�Y��>�G�.�.�h��z��|OK�{�͂����|���;�>�.�0�(E�h���(`���J���R�ul��^Ȣ��I�l�O��F��[[r��*�H�5R�RR�I�ao>�1n.��v����:�{�95�Ϻ �Yذة�|�!=)�t��gj�~3R�4`�۞@���>��Z�s��qb'b���S"E�lC����V���>nG�>go
q>+:it��8|8�{���C=JR�q��d���ݦ$���[��I�����(�ע��������D��u0���,Z{e���|�cA0���c�֞���K�R�wr9���;�*��U�z�_j�է�}UJC�Y�{�T���b�ת
����ƭB��[/=3J�UtIlu��1cXcn.{�B:�b*Q�P�|���h�/N�8�ُO�E5-���A�9��������^#�T@E�����{\�m��HeړD�kcɕ���S6�OV�s��FZ�'��U
�	����֡�T�<|3ҧ��$�fI��^]�]累N��x� u���7�TbA�G�ߩ����ק�)G�=�2�L��4�<י��{6�t�l���u���Z��B-� *�S�@/���,^u[���+&{VԾ^�'k�^ �e��&R�%C�T�3�  4�
�
q$R�-
.���^!�6�|�x�R#�S�t�U�.H.
���ߛ��|�BĎ�58����nT��?��i�ܜ�Zp�+
�N_���[~񕺘ꇇ��.��N�{�\�Yvl�˼���f��O��"'s6�X���vr��Y�I_:�8��l[F�]?�c}�+�4:��j2�S��C#�q�O�Y�N�t;a�.�V��4Q�)�o8{�-���ܯ7)gl��,6N���:�G)��<���,�����;�6S8w-��mΙygg:�M.t�W�Y��pZ����7dܠ؛�/��x{�)[��L^��)�@���ѰՌ��Ϣ��'¤\d�<�Q�u�Vdar��Yk����-�z�����ʮ8)�͞�j��dl����-�#Y�t��ѿ�<r߇�0�|ԫ�}��
�|kDm�8Pox�Z.�,'���oJ��%}�K�u^�:��7E�n<.�}'�ݝ�Ҟ���P�
�=[C'ִ��G�F���	�Z�_�k������\��t�)*�_B�����P|�ZG��8v��(C�7�܎� ��Y��ԡ�#3�Ξ(R�ާǬmS�T(�:B>���F��P��YE��t�Nǋ��L��mZ}���q�Xޡ�^�7ev��Q���0�����z�<ʋ�l�=W=��?(�Ot�y{�3����̎Sp��A�X�!*W4�y*���=
�Ԭ�jW�����S�zk3u�W���65�w]����և�q�Ī��h'.���ج�aV^o8!l�Wa������Cw�1K��%{���.(r�^�T^��Yj�R8K:�j��Q���j(����F�&{96�oۃ����I\�n�a��]�� 9n�B��U:G��Vnr�pMWT���G\�K�r�v��VnL���ݜ�i���#��ոm��6��ͼ��bޫ���܈�Y��{��a�ky�d���UB����r�Lu'7영JNK��+�"T<���)g���WU�Xwr&�����nYs�b�g>�ՙt�L{XN����tڃ-盰rY��8I����m9�r��v'V����g�]���E�h4/˽O��8Y�o�;R P[�wHL�8�n���=$p��U'
s0�<>EW�i��S�B�O%��9ؿ�y����-�}��%����%3��{���l��#�a�v����a8L�������7�T;�|~�{�13����$��jj�L���{�L�СבC��7����E�}�ֈ�)hqFڰ{Pb���P�4o�<;����p�C�6�v燯"��S�j�y�v7⠸*��J>B�׶���:�hi�-T9W���A�a�6�rTQ+J��x��ՎT�ϫbz�߇D�u^���ٔ��P��>�>
�q7��tx�G<�熨X<�y�?q�^�szB�((c�u����|,7��|t�w&�IB-VZV��u:����PO���II]����f+&��l=���U��f�Ng���)x�뻂�sޭ���'K٤\�5�|wu����F���B�d�ڏs�*l͗��}�j���qTr8:S�����"�~��<a��Z��� ��]���a�{܎�
���L��D"t@���!���!��R�=wPVD1۶��H�gk�e"����$p�C�rC����'�q�t�U�>��)W�� ��vl�([���g!�߸�3�)�Fj7��7S��t����0��I�8�7������
���k
���0���M�4�l�1��s!��Ͱ��!�
�C~fa�bN����ɟ���6�|��Ă�����l��Ɉ
-ٜ��Y��$��U&�r~��S��]{EUe���Cm��77���
�0�{�k���6ZE�'���ٺM$�}�MO=ɮR��<�։� ����u*,?{a��'\`�Oq�[�X_/�r��d��9���� �_�j�a�Ag���m6�U%I��d�1?g0�:�d�[u5�O�Xq�C�RcO-�eA@QN�xo��q��7�']���g�����1��'h��"Oo�oW�>�0}�&2t>�M2�W�'2�C�ֈ)�
&���H=�{a��<T*��a��ef!��uE �u��aS�CbV��Y�=5t�PlL��E[�+��rt*��{�>7���:y�N�P1&�=�L�'�́�eaXVi��MϹ�i���Y�w&�R
u��ri>Ag�0��WVf��w�,4�Y��lSH|�`D '}�"2�_Uq7'�o+�(	��z��ǳv{d�Y�<�����
�vɈ�Xc
���}����x��{�a�C���4�Y����6���ɉ���8�� �
��_l��1l��v����G�R�����wI�!�̟�~q'�Qg��bx��yoP���������l���T��>�!�Y:ʝE<��I����u���'���xL@�%�i�+��j��:�S7�<Q9�捌�ɹy�f�}�w��me��U��ve!,�V���8�I7���,75#pX���u�cӖE��j�:��Ul�N]�w;�d����W�����&�� o`h�˧P�i\V�G_j�"�/5s(�dڼt�`Z�Ǉ9�i��2���K�&��GQP�En�	r�Z���m�ճ-��4݈�E���}�۷Y�f�s/�L�UHP8�,n]6�ۍ�9�B��.�خ���qA�X�uw���Z�"`Ӻij�e�����#zQ��N�����*C�鱥۰��Qn����^e�a���6�+��~��,Y��&�����v.��p�Ԡ�av-�m�o��WE���b5�4�^�A��V�Vq��
4.4�D�+
�dN�1�&�����h���v��Ԇ����*E�MQ�u�����^��Me��Y/4T��ej��k�lh�m@�@�ٱ��ȇl�}�C��9R�tͩ��o|�-S�r��F;��F�.��%V��]\�:��w�1���ݘ��WI�ET9�gkXy,�*�.���n#�_?�����%� ��1�9a�T�J��]Y�&JlI��lAN�s~i<���t�Ls-�VT�G��j�r�䢏�>�S�0gVm�6�v�y��8Ǎ���7Ӣ��D��i7E˸b���aG8*�1+Ħ�����iIIf��5B�>8w쵴������lڤ��,�;��k!Aj9�����l)I����j'����$�e���Ŷ�J�;���d�+�m���AQv�n�|Z��B���su�K����޶8��ޜ1�û��!����������u���&X� .�/�K���}�:�E��VE@���H�U��Jײ�0Q�z�k*�;�1V�����4�h�%]i�kmS�vN�c.թe|̗cq:����%}������7y⦶�D�t�f�6���g��Si?�%�2:�����Իt�8���M���*���hX�1E���y�cu�*D�`F�z�@�*��V��T/5A���MIu�]y�޿�Kz�i�Mq-G�Y���Ӿ��撵�W@k-�'8���o�6I;�J�9�h+�L�2VV�\x=�1��9V,�9^�j�^d�]63�ͣ>�����'ғ�⮑����.�#wzn�ԫy)R�O��v&Ilr���]������/�Kn�R�D�QgWu>��z����p���&��wji]r�T�8�4��:���Ԑ����o��`�C��Qn<(���9կRw/�B�#�D4Bq]�zGX�t[�J��m�x���#��o���/Q��o�T��5of<c�
�̿����Y��ev"%��u|S��5��͝�%���]cT/�YP�'M������m��+�x�y8�2�R��{�w@���iVe���{��N���W��pp���'k�jݟ��_k^��޷���J�-,�VT�b��T�[%�j5-�e��4��J��
�-imk*�VQ-hU��YQ�U"%Q�Ae�����!Ye��X�E�%�Z�U%U��e�V��VT�+%F�UTU+bR�Z�H�h�[E��R�P�#U��V�R�(�J��D@�mjQ���Em�X�J�Kj����iU[eJҤ�-��Ub6��Kh�(��Ҡ�B���+P)mR�QKh��Y�DT�YEQVVTQB��+-m��
%jE��
�4������jb%h�$Q�TeZ�J!mFJ"�ڶ�D���V��Z�
�ګ
��B��KB��BƵ��mQU
�V��
�����)mJ�mmDc!R��ءFV�B�UTP�)b��ڍ���Ub��U
Z�Q-�KVXZU"�[EU�)*�#iU���[maVі֢�F"B�Q &��Xt�[��]ack�E)����}S��{�<����vf�]�r���#P����[��f���۝3�4HJ���� �ޚj�<���B�1����M�(�a�w�bI�Ͼފ��*nj��4�d�1���1��W��wX)<@�y�	�eH>��'ua�B���`,5��D���$�nc�pf�;�UL�	�<��L���z�!�����E�{�$+{��S�L@QM��
M;t��b~C��y̓�4��
Ͳny��ϙ*o��4��S�f�מ�έ�<�V�\q�[}�}�T튏gܦ�R�����y�Ă�s��O��E'�{����bO�ӻ�H?Y+�QM��AC���3^Y1'�Sa�<�ɻ����6��"7/��ő�|��{��v�)����	����~f (�d�|w�4q���;��]�+K���'�T�Lg�?8�IQ���'̘�7��x�H?RsTSL>��l��~�/܇���?1U\(��_���"��T�l�0�I�+&��M[8��Xq�H)�>��Y4���f�;����I�ӻɴ�'�;H{3��+�&���2M3�J�כ��o�͙{߻���c�������qYR��a�B��Փk+4���
�sˉ�|��q0.�:�O�>��I���2m�c& .���$��13Y����]s�[���u�}���C�?3�&��L̅a����{�� ���氩*�AO�e�OPY�jk�r��1�<���
�]�Sl>M��
�<�16ì�:���t$Y*s[=�����y�|�7�������9�m1�$���u���1;�"�l*g,<�d�N�Xb��P+0��QI��gz����&��8�Rm���'�^R��l;�O��>��3g������ݽ�L|G�(�p'�l�� tI�;�>�R(y߰<O{�I��04����a��͠(�VT�ޘ)4��T7�e��'���i��R�Z�d�
)�{��������O5������9����d���a�*�'�O�v���4������7p��̕�l�2�AO��hhIⲠ~<��!�XiP����4��e{�(i�0���������3W�����]{�� �X�z���l�a7�:��l��J��a׎��r�H̖���Js/)5( ^ї'-2�q����=��B�r4��s��2�}a���銎BĻ�Q��
����޾�]f)��د7R�����=�.l�z�$��f3>ӿ� o<����|��?Τa��ϳ'�*AC|�����?Z���+��~��Y�M�p���6ì+<L�ZAgX~/p�|����y��OPY��`��i
�y�㎾����~3���}�}�E1��*L�3L>LC�*/�V%a�1�CIVO|�E�N���ۉ:�f�d����(��
��w�T+�;f�E���$��
�������/�n�':�;��޸ D��>:�@��I�x�쟙~�+����t��Y�Փ�O\I��i��ɭ�6�x�H:��ɴ����ﰚ@�VqYye@Qd�}î˟�~���o���e��4��=0<`	�����Q7l�ɭXyc���}�՘�P�3
���
�g�bz�띰�a�
����m ��J�����@1`l��@�Le78tU;P=�7�6�����o]<�>�+;�si�ֻ/�4�!�z¢����i6��14��;̞$l1ꨲ��<���&�1��f"��+��<7f�z�gY7=�|�
��
�Ӯ�޾�5����y�|��Ԃ���hi8���k~���Y�Ns�7�!P��3�u<a�
�п�+6���4�{ˉ6���w�)�H?�w,X�I�1��՘��+7�%��)�?����~���w߿s>�
,=aS��s@m'P�<�yr�a��~���J��w��O�6���9����
������O�y@�;�6��e&�����+?$����)�R
z�����ou̞��5�ٗ<���{��������
���@�c>����4��;�0�@Qd���4�E%I�'��>e�u���ygXi ��XwVq��w�օ>d��� 	����x�)��]�"��Y-Uã��￾���I�0�0��J�Y�N���좐]����'�ʂ��Hs,8�<�$���egP�|¢�Oh�g�1:�'>ʆ��@���d�}�͵	�}�7gy��?o߿~�>���J�?2c9��$�>����x��Vc�G\��W�u���R9�Y&��J��S(b~@��l��a���w����aP��I�����$���<�x�ז�ʊ�V"�F�u�Z���o�t���
�1DS���\ռ��U�p[xV��M�TEr�CJQ:���S�3u�ܷ����Ŧ�뽶{�C�(Z�v����=3���m�H#&�֘��g.w+�N�LV�c�Y�����ա3{)F���5�b�� x{ʏ,�T{W=�ޘ�����LC���m�<N���I�����ɴ�°��oE���8�g���?Q@�>�C�J����4�2T��d�M�&=��T�@r��Go(����� �>�O��Cm��I���s6�YĜq��2B��7��>0]!Y7���h&0�h{�ͤ
�4Oy���Aa���1=E%I�Vi��[gY0�7�B��2����?
Gz/���6=6�P��Ì����z��N<w9�~I�����'�l>d����>I*��9�q!P��1V����������3]�����V|�3�N�XAM3��׸!�����"ΰ��i�z��N�g��!�~I]�|�2J��+:�����>g���l��R��a�J��UC߿j���ͽ�����3���>�/I��LA�?wQvÌ/,q�gɌ<aS�P1��Ɉo�LH)�KܚC��1!��9%b�'bn{@ĝB�}���d<H,6���	����{�O��h��i����	�ٛ����m����Y���:�h~I]0�ްq��jg0�Y?&'+�4���x����i�aܤ���Y�<7�m'P�=:���~�j��Q���8��+~VE���Y���?yA��s��uRT�Ǵ>f&�IXw����2�4ÿQ݇XT������d�ެ���x�q&�i'�T����v��4»�ɴ�Af��戹��w��&�>ξc�鍏{`T{���4��8���ͤ�;��;������v��P�iY���f0�7�Că�<�0Xmu�`�P�%v�a��ACi+�;�ߕ���>ٍ�Ln�f�� 8PǾuzy��
�o��f�9��>�3�J�d��& T�|w�g~a|�{;ܛa�>La�<;��Ag�116_�RT��f��mɤ1���q�n%5�YYt��߷���gޘ�G�G�Rq
��}ԛH,6y����P1'���M0��
�����I^����6�̕&�������l�w�m'�~�&�wO;�l=a�C�~�9�3�����e�dث��s�+
�Y%�]^>�cr|ʁb�+*Y���Y6�i�����nu��L��i���͖6��\�e$;�۸�=Co.����f^�ov��}�,8� ���e�
q�o�d�d�c+�{�7~}��PbL����hdLa�IG�xx�1<+.s�@<H,���R|�����/P���i�6^sPĂ���3���)�y�'YS�����'�1��[gY�����
��;���?>���9;��|�����G~��@���*����m'�T�7��]�HV!�y�k'��+�&?2y�P��&'�I�g��I�!���R
x��Y�1�Oyf�H)�q�޺_<��=]q�%�f,���?���*�|�߇�<E��V{�d�C�J�|����*�y�����?!_�����W�f�=�OP�|�S�+��� ��
���tÌ/(=�^��{����������}�zE�g��O9f�6��t�<�u
�AM��u3�8�0���k�%b�O���p� ��WD�?Y6�����O��1'��L6��E�f��~aP�J�!}ݶrQ]w��2��0�_Q���z`>����u1:���i'�s,�'������w)�hq$|�w�|I�*,�N�E>d���<9���&3���$��Lg�IP���W1�����m��}���1�tz`t�+�X~CL�e�y�'7a�'��ć�go���u����e@�O���y3����a�o��m�������3����YE<��O�(�����)�������{��=��7�Yă�'�
��32�eg�1��E �f�Xi:���ì1|¼��1RW��;�I��&�wo�1'�u�8��kW�s�9�~�X��v�5e�.U ��Ǻ=�R���&��%La��X�����*?8�����L6ϓo]�i �l6_�����7�a�f!���|�g�%bͧy��AI��}�����:�����~����7�& (��p6�i����!�6���06Ì*�p�sm`Vu���E�ɴ��{7I���ɣ�rk��a����
�S��I뤝J�h�_?��?7��{�{Ν���q��>�4�~�m3>�s��t�rM��IRy��Y=eLE�T�B�c-���'�,8¡��&$<�q��A@QN�a�si�
�HT�}����||;u�0
�WQ���Fv�����~1{W�VvBR�`]ϰ�v�ޛxy�b!%tmj=ki27{$�ޱø�{���p�\x{��4��98��\��@ m�@&Fpu�rO���[�@��VHE.ɮ�Y_�����bg��>����?<�HT?��xɴ�N��Y+�N�>;�h��@�o;��f�l<���a�P;�cƲ���"�H)^L�
�������������U�d¶���5�
/LI;{����W��̘�����&�� bM�Ol�>d�;�<3�+
�2w)���i���Y��ɵT��a�{�I�<q��xw��!Xm�Lf��"<�\���
��+.l��������C��LM0�����1�v{d�Y�<Ì6�Rn��Y�Y1vyq��T�h�}����x��zsXE�aP�5;�&�0+4�}�lUP�B���dg��%׬���������CYa�w�,�R��g{��'�T��̟�~q'�Qg��bx��o��!R��o��l1 �%J�*J�~�!�Y:ʝE>�@�@��>�����e�ow)�g����6½;܁���c��iE+��v��R~C�k
��k$*~5g�2x���Xc=d�Y7<��)=@��'� �f��wvT*G�ȏ��C6�l��`Dx����݇��
�Aw����'�~C�wa�E�{�$+N�6��Sd���v����3�&�'�٦�Vm�g�ވ,������������ܻ������ +�����'�u�g����
�l�a��Ă��w�C�������p4�0��CI�wTR�J���)��;�(c5�zj��0��l�u�B*�D^S�?R͙X �i:��{�?0�S���4Ì*�}���g��f�^2u7߼��
��;���:�v��9s�C���
��}�4ϒ|�M%Gý�'̘�7��x���
G�k�3c漎���.�[�D�s�`wW4��*J�VLE����yi1'�+'���5l�'ua�=�]$�֚��Y4���f��>'*N>�y6�d��i[�W�M&G����:6z���5�j��Ǯ=�C����AO�7�`�>VT�۰Ձ�v*�5d�������
��ˉ�|��q}�`g�a���}���
���d���L@lu����5Ig��2���`WXNs�_�4w����uvK���ْ�3 d�7Q��Z��w���:-��*q�[ˍl��]�Q�EefC9�{�L�d�|���|�./�,�}P�Wp�rթ�wV�P��ʹ\ Z�N&���g7a�z�L)���}���U[;얷����`zaG@�:�: 1�xү�̅a�
�CG���Y�M�k
����іE=Ag\a�\�k��a����m�XT���m�ɴ?!Qf�*i�Y�u;��<����z�ߍj�{���<���އ��%N���gSbAw������1;�"�l*g,;l�N�Xb��(�T��)1����nj�H
/̚3�T�I�6_��?2���n�=�S�y�����w�y���*N�3�?8��|��$���wO�T��N���x���bO=��6���7�f�Y+*h�L�I�*�2����>\����
�W���]R��"�~�y��]���J���/�����ڡ��'���0�̛L�7p��̕�l�2�AO��hhIⲠ~<��!�XiP���@�����0P�>aQIo��^�o���������o��Y�OP��t�m��1:O3'�*ACF��i�8Ɍ����+�?~�D�Vu����� ����<ֲ��ΰ{LO�UT���#� \�"<b�λ3>���O����U�ϼ��j�Xy�!Xc�\�M���@�S��!�ɫ��1M�!���&�5�fӌ1��n$���ϳ��L*w�xw�T+��w&�E��~���G痾w����?}�CI+�g�͓\C��M'�&Ӻ�쟙{HW�P��I��jɌ�'�$��R
c&�t�x�H:�2i4ý��?~��%g��{�_tt�O7������o���E��t���u�&�����>fퟙ5�;�B�L��Y��Mw��Y=q:�Y�?!������{�0��2l��6�Y�%vyܓ���Pb+�8����O��<���>��@��D�>��n��,>Vw�ͤZ���L�g�*(w���g�14���ͤ,1wx��¤���I��i�nj�EWoy�6��+:ɛ狻Jw�˝�9�Qw_	��	����?n�Y��O�4�IUP57�O*u�q�9���ԅC��gSl?0�>/�
Ͱ�1!]�����0�bn�
z����,�c�e���?g�Nq�ē��?�-��Z��y% �z��{4��Ϋx戺٣��ۺ}vƙv�[�T&����y�!�ݫP;��O0�C�S���Y�dSn�䒖�S�
����x���#��
η�ss�]������@�7/��L�-R4��ض���}_}�U;r���������?$�
�yd�M� Qa�7��I�
����k�(��~LC�+���ڟ2mE�y��:�'�'���yd����y��z���~�#��Uj�a��<�_�vw�z)�)6�O�Ȼ`��X
����7�Ow@�%g�fH
,���M'IR~Cܲ|���ü����XuC�v7rXH�f�p�T��m��ַ��O��������<2.�2���K��A�����po�y�P	J.��K�͊�,����V#b����*X|x�cP�o�%��5��x٭�u�wm�v^���u�q�+r��t��^+��U�bu\|���|��X�����ݱ�����P��p��V�m"��K�qz�T7>e{��:���t60��ų/��6���qDs�z�J2�]#c\�u���	���և�qJ�]\;_j�)D�(������
n��i".��V�Ƚ�a���Pr�gnJ�!I��kZ�⯗)���0+�"Al��:��uxU���r+$��>�Ow{�J�Ra�}���BZ���^���C���s��U�J�!���������jG�`rd)z"�5ѕyiS��j^��ᛞ3��/��ޘ�,�t/��yM%nC���7jܰ��E֧�1�od�" Юͦ���Eb7[�<��p:�����-�7ze�7mm�ur�,�;��ceHh�K{�����ڜ�׸g���b�xĩ�fη�1җ��$6X����VDS@�:�eʰj��\TYkQ�s�9zzNa��=�S�H+�  R"\��!�QsZ%G�h5q2	h��E�\�ꁕ�˅�n����;�F#]��R�ny)�m�+ؼ��l��#�Zq
��=�-�f�Z/�]K�\��	���7;�h� ^�p���}Al���L�����k՘�n:�ٳ^�S`c�H��hqFڳ"S|����k�x������R:�̬�]nv�֮r�E������/���� �9wT*��P�!����)1gi���Tw�^��u^�ƐԂ�:���bz�ߢ��;=�u؃X%����o�d���b�
�l׳�VBbE)d>"ݧn<C�S�qUt	��v")����+r{<h��A�w!�B���{��1xA^���)�G\XΡ�J�6!��xrcR�s�W�Y7������!�ga>�J �����Z�Տ銻�ӧ�GtL���#�Q�MI����l ���\�`�7�5��,Ȯ���]�|�s�¯)��u֍��ţ�[d\Uh>n���e�(N_=��8p��ھ��FZ��v�K���޷�rnj�W�����7�L�S��e�__\���v��,	�.vU�)OoV�1W�!R��{�x{��ɝ/�PE@�רq+DT�D9��E��Jl�rXr����L�ʴz���P��x�}c9fws����i��	S�#k�W!X`�M=/��M�5`�P�x�8)���=��5n�%�r5#X�/g����z*,P��Hɇ>?g�P�u1�γ^�h�dm��ZV}���}�1�z��.�C$��}#P���
%���Y�o�Uym����x�,�!6/��>�Z|4-�Cq��H��)��mX>�씪@�,."c��1{�Ϛ̬��{��<�s�Pp;���\��epZIqo"ft�%�y?N�i�4�q���j�yOz�rCo�O�x���+�B�})H>��no�M��D:zTV�.z����_���N+> 6G�w��u=��b�3��®%����es��8�b����}���w�t��L~�؀*����L�~�4��-����E��"�!1!Q"N�F�F���-��Ԏ�D�ǈ	�y���\��(�}S����.�OvD�%�rݽ}IX,RtԺ6�Lo5�޶Ʈī)iG�Z�^%����2s�=�`%�.�-C��˳/{dѼ�)#��QV���Jc�o.�:��ֽ���H��Bg0@D�����)_e�}̝y����p�����(�̕����{$�u�Y�ՅQw�{��'�72S�&E��n�r��w���js�\�O���ֺ��^V,�������{��άͻ�v���щ��a^MlZ�'ɭ:}�OJ����g�o=����X�=�^��qm#�;w��=Z���H�(]bv4_T'K�tw�Ey����d���� u��W8Q#��xfa���lZ�� �+���r�@���J�('�r�.G.��t^�X���S��E۾�Kɤ&k�ܮ9ZԴ��|��Hа�)R�7��������+-�s	2�o3�'g���&B��e��%_���|
��89��ھ>���h��m��j������H��t6=g{)�Zu��>��6=��H-DW��8B#n�FU�峊���c�ɏ1�A'�]sP6�Rw���֩��	�� ���A޼��@�ff�u�(�m��7�Rsb=�H������qq.���T�Ms��ͼźӹ��K�����©�ZIV��4y1RPu�+�Z��xj��<$�5�;��K^V�L��/�i�7khIq�'#���L�����u׼�Y�#R�o�]��h�EԛF!m�A����u��
�q���c�#�{ў[�^]���M;@إ,�X��T�
U7����谶�>W]zj�j7�pL�Zg<�Ӟ���S�U����X�v=�pZ=\��%�u���[Ů�A�\�L�2�ǯ>1�{��t�̜�������m�4>Mg��[F�n6q�5��+kG$b3$���ݝ���q�Ou���o��0L�_K ��9aZ�ѻc7��6���Y*�e<���Inu�vk��ұr]�"��a
�3g>�Y�[f��S��֮��˺��oiV�	���y���6���B,&�z�w��:Q��*����Ɩ�ki<@�+�lR���Ԫ���Wl+\�5Ք\2�&��h��:C�*��,d�U�����cn���-�c,��KMN�n�j�jBe�ճ�*�9���x�
k�~z]��ˀ���F���h�(Y෰�fδF�oE;�پuI�v-��a��Q�B�8��;Fn�k{���8�.��ܠ�����D��|a<�-��,��6�U�`�	xgQغ2kCC�Q?|mI���avĵ7G/��obi�ܼ�.f�gF4>���@�3���v�����֋��Т���m�z������m�=y���v�쵎�HZ�x3�5���y��Q�>؁O��.8��u9
V�ӧ��]ޚ3�&�+J�u%�޳;����,�P�v�N���ӆ�3*gW#��}p��ig:�Z9Pz��c|���t�j�g	a5�#����w�ΩwȽ��:��������R��h汶�YN�[��:(#��Ѫ�� �� ;frპt|F�Ђ�=˭�ڏc��i�Yԯf�4�ۧ7����0D�i}���7��5ABޝ�r�Z�r�u՛5��;�|m�\c��6�1��1)R?XE QM]lyF��bpp3|/ys��%�ܚb��\M���5:��i�D�_p4z�ֳjε1���#xя�n)�N(����&;�mn�;"��Q�r�[+~�}qܙZ���
d���6hG��N��l�]�]KY@�ul�ZS��wr�
"�^XwumGG�_Å�����i}wO����F�=}W|���#-���ܥ�Xt-�rs3;Q����� �;܏4�}w���P�'�8to�,��.G�W[Q����>�)��wm@��1�c;c�K�V\� ;"Y=;�OF�o���k��$�+E-�����u�Ƨ����J�NW{�ǰrM!"���y%����I�.��:\nc3��tu�Ғc���-x�v�f�L��S�@�(�Wvq޶^D��D	�U0]FE�]�N����czq�J�[]C�%�����d�K&էMtR���oq[�{��g��{�����µZ�V �U+)hՖ���Ub,V6�{��4�)V�2����%D�,Ym�*Ŭ�Qmm�1�

�1���[d��D��e[FUh����*�+E�!Yh�ڪ��`��J!X�[j�X-�aR��T�,�ʄ�c��)�V�IZ++KAF�ZZR�TJ�PP��Q�J�b�k%V�ed�Ȱ��Q%j��-�����B����Aұ
�QmZ[DTTV,Km�a�*��6�Z�-l�X-J�d���1V�`�`�,�����ԅaR��*�B5mkP�����H,���`-I
�B1Q��@X$�aZŁm�Z�U�3�*(A�+%eU�+	Z�+�Q�ٕ���K�o+pu+a��d\oev�̮2^��s�p�2�p"^����:\�e�����H�J'��ic0֢�wϷ�_ =�ռ1�q.sKDg�D����W��@��� vX��"`�>�,�����Crt���ȶ8���:`OG�6P,ԛG��������<y�5�3�rò���f��58�>��A[%J�m*���6Ռ�Ϣ�;Su"��Y}A*nq����,oF�ҏP9W9I�����rj�fp60���p\fy�<�`���>��g�O�R���	V�Pɋ������"�"��}Z9�Qu��ҡͭ[Η)NI;�^�� �f�ƽ�3�<�Σ�s�������C�����s��ܚ���y+b�"��7��J����^cz���౏@���y0�s1l��p��MC��5Eo$f4~ͱ��Z'&�7����]> U�����0u%����m�����$v=^/%_�c�b.dwȷ7�U�+��Tl�T'Dq�a�Z�0N�u�"1/[Qw~�¢�_ǣ�W���%=G��{�*��#<�l�o�9��S�xD�3�z�d�H������9�W4$�oCV�Y���jl��hU�� ��r�C�^�Ī�+"̶��-+��5Y�A.��u�5a�l-沬��e[�=I�VF�ٔ�< �֭�d�{�m�8,kCb����V&z4ngJ1�<�=�m
�N�����n�㏊6�|D��Y�-����>�6���(!-�����r5��w4�/o�L�f�R��_�X�mY�h�k�1OW�`���u���G~�%\�ٞ��bj�G�|�B��V��Ϋ��G��?�E�e�C�v�.����.�N�9�M��V�X����||�Е�爈�xR<���c�懦��E�q�]���be���os��a���[�+�pr�?P3W��W�s�B�40�]S�+���{��/�
A��K���e��󈭩2�[�AE]8T&s>O��S����B@��jVfǤl~s��Y^���K�iz˃ch�V�l\y)�|���^���qB��q��Og'�n����A���j����Êl���nwф ��nc;��Pk!���$�8x���NMA�6�.���� ��8�WJ��Y�S�EP�4��c�D��z��W��'��LxٓXĝ.���ܝG͊V�QΡU��uG&y#�v�y����6�WW)xk+�N�ti�j� U	:u7Т3���{�m�W��c��.[�gss6������0�ܑ����L��ei�w*�e��n�n�xs[\����fVZxGTd�['t��"7���j^�W$oe;?Ae-EFOo�����={�q'�>>*�!�:α���خ������Ŷ,�]uu�ʃY���3s��;v�)��[�R�C�c;�!�)�8������L|U
�8��S��#yU��f��XpF��^��!�u��S�%DAs�"�rGd�jht�Q�Ic��V���N�͗cj�����M��ח�s�8Kj�t������BѰ����y�]�Ҹy�>,.�3;g���4 �8�s�%���&*|�5�E�׹>��ْ���qB_��^3�![Zz�s�yIl�'�>��籸V/�_26n�G��h��U��K�s44%�����N�+)^�$1@I���a��>��V��c+��� �a��yu}L�~��Z��tR�w��Ν'c���*�.���Ց�6)=���vtE㡑 �P�@=X�Z�Pu��}�vF��8��o ̯k�kN��=���q�;��X3�6�.c�´�a�f.z%=�����)�U�_�d�`�/��ux[�]��\��%�`Hc����C�Wpw��?K��S�K��8%��+���핵w~x��Ԥ%��1���Z[��dłfN��-��!-����b�ݻ�7{�w�7�^���#v��I�( p�ᇹ�i��J��@(vQ��o�SS��� �����ռo�BQ?{������h��|�`Ԯ
���OE2V�3b�I�<vP���;yP]�X'q#�:�N���]��{��Op-�$-�u=���R��X*%�1b*���nc�Z�{3�4�p���:[W	���X{dLQ��9M���{�8f����e�z��Q��re�A�B�muA�]f�>�囮5b�������m���d�dԶ�y���\��N�F1ܬ8��.�t���J
��/(�_@��{5��}��Y��^.�����vw5���H���K�
��ش�!t�6Z�r�p�*��+�y�&G�Qݶ	.V�3YO�Y}����1##|��������+M��fs�L�=�} �=Y���oʦr��Zax�'gE���/ֱ���ΰ|�!W�@DV�Em(�l��4��&
��q��+/�*�f����6�O�}���W�jt�����^�X&o�|�ܑ�	�ֵ���/u��@`����Py���_���[�Q/����ëO�'�3w�T�{)��٫��*tz�6\�w��̋gTn�wmi���B���rV�F�ojI�CU����[��
�W�8�qY�κ�%o'��t�	��V�ח��0�e�O�<A��\ܽ+�y��d<nc���s�PB�휂t��N��b�Oa�@��<<�ND$tS-���߀����l����wM�:�
�]��č�l�#�������$��k,Q���wO��oO�w5��qMZt�06�>�#T�hE�y���D�1�d�ܿwl[H�3�i8����^0��ȼ~��r����P����#L+ ��#�óR�Y��I���W�?j�P�i�lT���`TÚ��E�R�
���d�8�	/�ĿT���rn�x��DМ_��������q{;�u�!@�:u��֔ d�Pj���C�~lQ�,J�:	�"���Ʒ�d144C��(|<�,S�����`l�0�B��ʬ����������Pw4a㏝��bu�����l���hSܯ1F-S���
�OC>�.6,aN�gQ��9ԙ�h�����ܪ7�k�F%��fn������u�o>����0���ػ.g�;|U��ӌ�2�*�p�@׼4�\�Օ�N�ÉA�?���h�k�;N�&�^����X���}v.J�"�U�c
װZ�}��[���à*��s����7����5Ě��KFk�L�Y�1�U;q�{�]kj���ڨ��D�rl.�`�9*kO-<GZ�H⁞�i�z�*�;W�e1�v[גn���W�^�t��-���sibmwSOt��f���W��=��z	La�V�1}YkbZ�`N�ֺ��k���<�o3K��c�W�O{������YV$�����.C�Uϲ�(C�;�7˒Vsv�^
P��P젬1���CHc��ydK�)Ceo>�m���=[�PD?T�\���C�E����_$�� ��w^���z�L�~s;7�u�z~R����G��W��qA)^��=��z�A���+��4�e]�,4`��#�;7��N����'(.�Q�,<hy	���r)<��L4:,=�M����xŪ�M������@���*>|x���h=T�"�:���nr�l~��z��n�Xn��ۙ��ܢj�9�oj���<~|��BAZbGW�`�y{��<���"��TĐ���Hw>��{X��Г��}T��P�J��N��
b�3���Ð��7ʅ7��H�D�˗}|V�E^Ǹl�����m�
e���l�x�bp�(��0����c����B8���p�n���ς���9�� ���$D�!4���dՉQ�}4�SYtUp����Y9м��;a攌�u�wV�R�s��������0S<���C��/�Z9TVF(P�j�#���ŅmFM��&��8�W1� ���I�,ӱ[ӑB�-��z�4���Kظ^��fS!�3��\�D�m]�w�~������nul~����c���XU';꽏��h�V���XJ�{J�/7�H�xn��B!aW\�eGR�!��l�59 ���v������F�/p�1���Hy�&���}�އ/[kӄt��	*�3^��*�t"�WhqFڰ[��,�K�"��*{r�]1�{MV�W��zOK��=B��ZO~�XU	Y�_{��SZ��|���fV����J�&��o0b�a�C�}��Z!�s�����Wg�_������`�F��8�B#8I%��Y9��*O$���6|���T,)K|����ǈs�qN*��<�蓿K@�ǆ%9����߽��U}�����`ь�N�ʥ\��l�=Ң �8Ұ��{�됹d�ڬŗ�4��IưRS�|6�����l�V�'E�j/�ckϤ������3�-���~Ix���=(��̗0Q�R�}��px�o	�r����Vk�㢩ْx�G�6��Y';yl﹌��S���m�n�9�����7
��4E�*����x]ُ�1���!Y�Uk�*�kGZ}��uaaU�'8�}�-�X��5��'G�>���S}��	z�_��<!�Г6��ϙ���W�o�,˰o5$%��] ��(�B�B�7K%��3�N�K9(#�.��;޼މ�y(���6���v���}�}�U�n;:�5�{g�\�ߕ�ô�t�Ʋr��91@���K`�8"=�(���Hl�ل�*�*��)a��{��s�{8Eb�Bu1����=�Jv�b��8��CJ���,�6e���r���c��� :��g�׵�A��{Y3��1�P������;R�zܞ��Y[U7�2u!��T�Z�6l�/��uʽ����I*G��Jr�+)�!W=�:w<�FMn��T��d]��= ��/E`R������5�P�̋v��Lm�ضys�7�����ݎ�(�ϲK�~�D7U1ӂ�2ˇ�[��ܘ��v+[�3�73�L�]����T6��C��R�1a�1D4}��R9BmL�Y\�R�-U���@Dg`ۃ����X� a�77!ߒ�����X"��EXQ��	��T3�ˮ��J;�q���{e0i���Qu ]�y���js�^P>OU�}W�]�u��c��ioe`-�쒐��`~Ĉ�/	�0��5�E�b�kɗ֣睽����en��`�A�\���w��̰7����]A������k�J�CkI�K���=Qr�Q��v�v˫qC$j�rw��>yl��Yk�K:���vw�)G�s�8�#����x��0z��-���qs���7��ޕen�p;,��l���ji&:o)B�g����G:j��\�l��*��!@�;f,L]	Hׇ8V�9r���hu��TrY��?a>����~�>�U1BN�;��*Q%�>�>�o�M����ʀE�p��k�Ʀ���,�~E�IA^����}}Q!_t|}Q�S�H�W�hrD�������y��1��t�r���#{JC����Y��^�(�;3��:����QSܪJ8c'��Î۶5d^K�-�������t`lr��4�l�"A��
�N�+�5��+A���P�Ϣ&���*YB�;`�=���!���ާD0����=��|,+�jӵԅ��r����0E���CM*[L��]�M��{����|)�0�O���C��V�@Y]�D�RIP���7��/���-jQWr1� ��
�(S�>�)�U��D�b�P~A�aC\���K2������Բ}ГN�t�1L�w���N�°�r�J�P��A�W\gc��Ҥޖ�O`��+�p��8	G��W�	6�7�"%���"r8�Ǐ1E^x�Ά�wm�n���ϐҦ���YN�H���wW}]�9�i<U���x�����g^6�t��6��q��SJ�x��gq���8�uS��E�[`,��P��!��|_]�
��\��*g�R�ͻ�uq6:L��"BB���͜+"p� �\R1{�{������o#`��V}G�(!;jܱ�H�8>�� Xn���V2Hg��X�zV��|��u�ݝ���гSB#0�l^�vu�����L�[W��e�e-�q�O-�㛃�.L�w>�e�B�^35�WY���to����� ���"�"5C{��^�ܚ�qxp+�t��h�Z�N����B��z/U�=�O�*>}��&G��t�*�L��e9��XO(K*/ѱ�����M�*�����z����~Ⱥ���c�����W��{O� ��i�������M�䅕�V��N�lsL��Ur���^F�R������c!�YJptڕs����jdu�2=Z��ʾ.J<�Ӟݥ�{��pw����O���1B�G�T��U����=m�	M����|��T�;�}K�AotgJf��t�WE{���X�vL<��ya�^Bb�!�"�]iޚhDr:jtǃ7��-�һ��Ok�
�U�8�-3�겈Z���c�}t�Ȭ!�T!1T��]��2���7��Q�7�6X����������l��zf���B˕�]t�Q.m�n�=�h�d<�.ѷ;9������;}wU/w���ɲr�Jl��%Y	v���Z+�/')�I�tt��~Ξ�h[��b��E��j�{g��=7T缊U4�1�ݨY�#Vn��KE�olm�;,�*n���3��Z�F�h`�Ky�)���N�=�-�M�*����ܖ �R�*9�+����z ��GDl��t_;J��@M��W�;�OE�]���9_W-�6X�E�kz;�2:m�z&��N���]ӝ��M�`�W���K=,����x��3� m�WV+��@�kc.�BEB�X�8�y�`������SwYe�Cp�[I��� ^���#`m�Vf��f1�Q̧ѸZ7�o�՛9 �нwutCS��E�̛��B����
���Y���,H�9�޲�i�Ie���NZ����2��2���	\{���&�V6�i�_f����?+�H=nf��%Y����Aq)��dWvh���;֔i	RXu���%]�s��2Gm���B���^Q�+L�u�ֳ�t8"o/����s��r�1��W}�]��t	"���p�G��~���"�϶7v����]`{����y��.���	O%�*ə#r��Ays"�+C36���y�d�����ͥC��)Pf�"񧘪;�)��r�n�lB�'o ����l׶�6Ԙ
�ڛ��'+���_LE���$�Ww"_pF�vҗY���x�WT�,<ނY�NLc=%^" ��z��K\�ޛ`촜A\���֫��,s�2Mٻ\����!;s>��a=j8*!�`���J®ɗ[7f杨��w��QX���X�D�J��]�ըm1�wt5Z�8�r�N���x5 %
��RfPp�v�D#O���3��T�[��� .�C����u�(�_;[v6.��,b�L�8�!$P5	�HŸI���ȕf�j���V3�ô)1���>�Y�Ju��4d�]ܺ��F���T
������i�iuupi��Y�Vn�2�u�!�,h\.�zR���ײ�oWj���;�h[A�OqCu�OD�)�j���]y��cY.�|0��bKlS��W�7K��vzPd�L1+�u���<A�!Mi�Ţ:���
ۉ�h�&7��ꌨ��_.f/�͓�&bҰ�d:�t�}
d<λ&YgV.��X{i������a{�bo^������t��OgwB�I棽w]�;'U�/E�"�IO��3i��e�+c��YtU=� �#�6Z�v�u��TK���ab:1*�|c�#}��s3�Ql	N���:��ؓ�t1�[[l�]ճ3OFp�n]h|��]]�c1Ԭ�8��Y�y�^+��ŝYgmrMj嶲�9:{�%�[���A@:�����\Q��ꫪ�U�*����,��1R�HT��X�Z�)T
�(�
��(Q��T��lY
ƴ�Zʱ�T�Q��2�%��[*Jы+�a+`V��*B�TEV��`�,"�)++RU-*"�hV
���
�Ue@R(,�72�Ʊ�-�B���D����V�eDaX)
0��F5�����Km���,U�����Ab��KEIQD*T�KZ�EA�����Qb*,*V*�����`���,(�dX��D@[J"*Ƞ��j�ҵ�aZ�B+�.�r���gA��a*�V-J�*��k���ZӢ�ɩ�Iv�G�WV��q�3q���f�G��ڡ+�Ʈ\�U ��� 	��&,��91���k���$�cc�P���|��R
�:��)^���"��h[<v�J̓ċ��9�ϩ�T<�%��/��v�,!lu��Z��ۗ����tbB�O�:�1�v<tmö��xݨ�t�{@3W����.p�QƆW��y�r��v�����L}�6^^�|kX��IQ"\��./�ь��*=R4OV&��do^ӹy�K)���l��U��';�+���,}�H�ױt�6���p�bX�Y^#TIt�桞�"�U�ړ꜀U�(]��uM�����u"9�Fâ�}ᢽ=3��,��&*�W���V�84�:E�n�p���^��]B��-�k�0�p�/v�+��p��������1�fb��%�@H*��	�|ؠ��j��'9��?`��ikθ��ӆm|���鎗�ݧ�*���:��y�;Ϗ�j�1	�Tx.g��Qgf���s�g%3:���}�^("�d�R�|�c�v��^7���%������3J�lv�����lѦ]v���^�����G��� �#�I,vz=�'|���_]��Nħ'�5t��ܛWè�jfw@�Ԅ���P5��c���¿�Z��uK/�n\s7Mm�}��ܷ��t�-#�sM��p7gMo�[�����8��}t:��èR��4c[	NL�ې��V��J����J��˽�8��t<V��i�rI�h!O�e@6���,��Vx��kӽ��La�c�j�'F�q,�8�����{BG}���!{�ڗ��nh{����w��7��A�z(-�AR)�]Si8G�{y��N�w#��3�)�Fj4H�*�:�v�XX�i�t�Τ�����-Άg�r�&�;<�.vV
��i����'*B��>+�L e.H��ǟ}�}yy��E��Ȱ�94m8�;��do��u�Jv�Ŕ(.0�U�^y��	}XP��y��P�q�	d������ms�D�[#E8P�mX=�ʣv��d����Ȋ���z*}C4�Eٮ������|\��z 9DKx���u�;w����WW;y;���'��m`�P�����V*��Y�'4�|iՔ=�n1sz��e�ީ�3w��i�>�	�:�v���Bq~j���WӅlH�#>z�."��O)]���5�6�X:b�\�=�7pa&���d% ��O9�b���f��������`�ԕ��mn/u�n����LnYܕ5��Σ'�wo[��/�����7׉Y ����F�{N�;�Rx]�YOn����d�n{7�J��4Аߺ�F����{��Y�v��g7�ɏފ�"��
���w�B�Q���"b�h�(>�u�cJb���h&�0J#��c�ɉg(�9aAs�}sp��n<_{��E�!Ḓٌ�f��'J�:�9ٝ#�Μ��X���Ov�\[�KVpr�f��S�^P)꾁�}W�\Z��X�-�xD��涽p�,�XlU�ة��a^Ml[u�my7�E�e�\*���fs�u,�G����L�tkش���p�|�혱1t��V���g>�tF�.%��]������U����ݔK�����˕]�t���ZWKܧ� )�"'%Du��A,��\M��tn�;��fd�ʃ�]co؋�7��X�V�/䎔����l�5�����*y�曆�>63����z��>�̗:�7aA�[3�oQ�7���aI�PP�x�|�n�婙=���������M�/�^|3ҷ��Tcu{��\}	Zvm�cۚW�B+��7(a�s����}��Z�{�N�j�?P3�8�����U�#��S��iܛ�p�Y�ˮ��pPU{�Ȥi-���κ�/ʆ��=\��Uƽ�D�iف�Z�;]6sc�:���b�1n걹`#\�N��)���Z<B��5�cU�ķ������A�Q���B�����8���\5�|�Q̝Gu��Z���lO�W��M����0!��O&�YL��0$qz{�u1�ƍ+r/�����>JSq��&�/3����z������=�;�Xi�P�����-����|�bS��ˎ׺L��[e�>��i�A)�!�H똂Q^��\]�a���s�sg[��j�\%�X�f��n�@�=��Op��:Ty��nM����d?���bs8���z�{��x��}��9���|�4�Y�d�#m[���'��/7Gf��b�d��U����Ϸ=�|�:�������<�q�t���z�U�p$�E����t2��g=Y�����L����)�#mW��z��-g��Ex�E�]C&/x��k���k�9�P۳�Á�xh1�Vr7卵e�v�3A�V����߈ƽ��`�����{1n�qs�1�1t��p-�\_�P�Xl	:�����B���i}��4o�kޜ`�}���.fN�-	t�IOϠ�v����S�UCbz�v�Hx
��;( =��b�!/A�'Oڇ��]���ǔn�1P�z]�v��ی�<����E���ܫ@≰�U������t+��qi|�Ǭ��.�j�=�'KF\�]��������9>Ǭ���K��p�Tl���]��h9\��%f�z�b~����nv�}��{�L�1
:m�Z���/OG��T��L�s~u�b�yU�^ZI8���Sx���cKTz�4�HuIx|�������S���pBS}?G���b�(������]�i�_�w���y �\Q�������@.�(����L]�0�S��N��u�/$�C���>��	�9�|xQ�$q*��Ϗux���J��8�ӳ"#�ۗ�A%+B��*���;�N�k�X���*߬�T�N�K���6H� �x�܄j�lS��_)�\�*�]����]�57�}G����Ε�	MW�#�;v;��}�̕{�=ƽ黼�je�CҴ���7�%����|�@@����\�P���^{��3��t��5z��X�0�G\嚸È���C1JC�$p�aE��
��u��������D�Zi�(����i���ֆ�<��.�(���r�?y{����v�l�h�$T����z�i���;��ӱiQ٧����#�`4��X�֪'?�>�Lu�GI1Sz��5�uE����x����y�hrUͲE��*ijE_j�G��4sRκ����r���|��P���uNorZo}ę��뜴x�"�D���s���Hh��a�l�u�;i��o�:�7��R[36|O�O�O���<T#Ӫ�sT������m��LקU�S�ch-H%v����xb�F`�N�'���ٹ��%t+�����{�z�Jc��	�bN[°OS����J�հ��I{�-�;��)�թ�(�!B�"��UU��~D7 ��e`����}����8�|�z']����諵XC̾�����u��H�,�V1�\{��R�z��T�}���Rk������C���]��ь7�Eiq�!�w���[��˝��~�Jwk��0Qk+�;�R��!��JA��Vx_^��>�cO�}�5���Q{�#�����w��g�bGhL��w�ZF����;��ڭ�rE*�P��ܒ�q�����(Œ2&�9瓿"9��V�+�4=�^|�F�U��ϙ�y��a�k��3��=+�٥S�\�u�o��TC��~^ô�l�]U��'&(QQ%�bL-Yw�s�yz`����M9�Y,�§Ξz�i��x�ڄ��2׼uկ
6)Y��0M�e���k�۶o;�[ضlj��f�q2Qݖ%���F��ܫ=�yV���w��1sE��,����=\�ٹZ����>��̽�ĉ�A7,R\��T9S@Z���1��.G�5ٙ���K��r�N����ۚ�"�����J^������g�Mv���f.&#�6�,P�q�@S��A���8OV�����
4(E}�w8;�O���ezn���{+	k ���Uhw�d�fE����.Z�=(�{����o��_`g�$
���1�u��4fI�A�~pV�I<^��{�L�_!(���$�Ɲk�O��o�7Jwex��%��I_ZU8�5SCF�N�y�Մy�Zͺ�Z���ĥ`���ȍ��ʌ���(v�pń�C��R�1a�1D4}1�񎚄6���gR7C��Uh�ռ�u^UGBy��}렄>�P�뛅�%n<C�vw�E�!ḞnӺ��������ݼ�~�gRh��!�ӭ�E�aE�0� �_�OE��/(��B��h�l�6o����c;���]x�V.��S�i	�M�c�=�L_w��E�Hw*�,�=	~��{3*�V$}ɑ1j[��#y��V:6�F�9�
��!�\T��BfMw����J���"<`�_�C�z����6��y�T%��hs�AO+��\J��g�����觥#�Ա��z��և}�m�g�st��ˤ���r�M�N�fe>Ü�����Fu �*^nq�&��pGf��My�
Kn�0��*�A�|�7�5�����z���Ϡ{�A��βtgKFʮ���R��Ӕ��xj�tur;%҃�.[�,���q��_|*�^.��uj�~5���ٵ ��(�z��B�>>��r��$t��;$-A1Wo�����r[ʇ�J�$�)ȱ��@��:���PG:ٞ�z�nC*h�P��3�>��v�pTپ���d�Af��o�k�5G^>�=+ye�t���wM�Y[�2E����d���罓c�vX�Ϝ4r�z�վ?P3��)�N����4�o�۵���>w3n�75�����Z��B,�H�
�+�����T��Ɖ�"������.�U�z���ŒN��צ��!��_N�a��B���������EBu�ز/�vI�<w{�Cr[�zmO��7q���3���My�a��
��m_$�C��y�L��/��颈�F�߇p�)�J�Y�&���"%����yU�W����E�gY�ދnc�C����^4�J<������a�>vG�u��Qъ�w3�]$�����mp3�艆�'�# ��9�£b����Q�*�8g�����ꋤ�����3i�Q����X�ԗ:rל2�"�L�6�7�koM_i��X���S��$�nfۭ�RU�UfʚE�t�ָۭu�'��H�{�0��Te�[��ނ���|�ݜ������t���N��E�퐫��I �0��FC/ﯟ꯾:���ռ�R�
MBR��|0�sꙓ7i>��[=�4�m�71Ju5�w2��s�-�W]�ԍ�o��-h�Mq,���&�~Ī+����i�@��kZ�Rf:W�s�R`�I��d�l����d�ch�J�@�#O����GJs{�L)��\�S3�R�{�C��.#
�4	����xCQ�i�Yٔ�O{z����5���1�>�Sr�fX�cZg�x�:t鞮���{�?9�=��J�-v_L
p'#�Ks��1٥+;{����Qŧ�,���#A�<�F�����]_������?G�Z���z��u3}*/.rz՗�1��p�(�|����2�]\Q�,<h!1w�ÑH�~S-�����͖�Ϸ�Xw;
�j�	|�9��~��Lt�Ph=T�<5>CHn��m,1���u�%	l.�.F�r��𧗑�7�C,���$L���|�H��C.��F��Z�p�����VI
,nK���Aq���V��X��1as8��Q�`���cl�1?���Z�{q��Qͱ�N�K���Y,�S.�1��
vy_k�V��8�� ��D�*v�S\F�-�x�y��-��S�C;�9Wb�m�����1gtn�hv9��� *mY�_�m�����kMYJ�L�{�[VD�F;��_���h�]�I�]���5i�F���1�5��):W�f/8��>+�?S���hw`0�.�]?#QPE�����>�H�r��XĠ�"_V��#k}/��֌(`����&A $pb�"݂}�B����'�)^��WAa�c�qޝ�9�ڝ��k��b�6o�����#�~�S�Z6)��Px)9��^��y$�&�'�/�¼�w�|6��F�V�u��2�5��iN���v�]*��ʕi����{"��Ϯ��,à�P��ޗ��=B��k��u�P����]P�D�AF����x��xR�
w44ʄ# �r�8���D7!�*rOV�7�Ξ��5ԃ�F���3|�`��G�/'~V�C���àJ���c;�.qN),�(���]Fj��.W�P%?r����W�*�+t���ipp�x��S��T��XF0�A�V"�/�*����@nGd�jXԨH:���	���=|MN�]e;�_P��Z�y\�/U�\W$�q^��ӌ��y���'J�{�����כM��YI����&V�X+[�A�)r�Un.�[�V�	Pl�c�r�{e�9b�q-@|����������P�]�3Z
�I\��9mlۥ�i������֞�[�3]�@پF�up�☠Ւ��c&�<�V�";��,���oM*Z���n<��5r�0��3ۋ�eEKIg�+�ڼ�ݛ*�H�>��+i!�D\�;v݀#e�ot��xw��껫e�M
�bH��t7-A�ʽ�b�F����̴ew:O(��V,����)�0_�(Μ�)g:ub���M�B&��u�ÏsG���:��
)ee��VԶ5�`gS��VS�ގ�t)KUf�WW�����cp��i�s�6��-CN6�hv�F��X��R櫹c�@:/��M�E@Jfo}ˬ�د�v/,2��8�BXS_.k�V�B�W0�Kr�7����:K�J�Lš�|�x��tp
�u�.�"]<�Zj[�5\��=�.��q���sk�������X��]�YugM1�3�}|KM�w�nN���Cu�7կF�/�^ZP��w`S( NA�|q6Ԗm �N�J��Wm�Ǔ��]�S�M/f�4����t�����]3u���~�	�;��!i��}�W��!@�\ߎ��]�o>��k{���s^�^\]�KU�t�c�B��6Y@�f@HI/�bS.�ج���*:�j�Uv���DFT����]�T�gV���]���vӦ�W��fkD�Gr�5�bG���'���#np���UpL^a�����v�5צpbɗ���nк����)Yv��{&��G�<�Gx�͵�+I~�6�q��	��	NCuܱ���Tz!L&+�W�Z�Y��|8V��<��ً+_Z�3jZ�����"�Ծ$b��ޞn��V�:e%����i��;�?,�ם�*2�V�9�p'|%e4&c���а�L�Y �:���-��mljNw;�s8�l���eo1U��<:�d����k����݊�gR��etF��WZ���59C��1>U���۪�Ģ���/��}hma�(���<^G^�`�����de��:�;7�v�-�ݼ�l�9`;˹ V]q��fu�~�C%�׽�m��a 27\����W���ü<���4�d�,���S x)����l�}m[��|����sZ��rD�M�kcE���xg}wuhd�YrVUr���'��qd�eH�EnrМ8��s���#��ï��ξ�iNB[ڒ�bR�V�Y4_mٲ�G3YP��V38�8s���V\�+T9b�1عS �f��0�J�F�ec��#]���l����U=��z�;j��	���Z�o,��iF�>2��A��*�A�3��c�'��fg9�����*'�6�
�22s}�[��)�i��(@
�| �m"���0�ڲ*l�E�VV��m[���*�XZQj-�r8��*U�*��nZ
cDjՔQ*T�IR��`�����ƣJU��-�VԊ+h"�j�1Q�YX�[l�-��V��4UA��m,�ڑʑ@XB�P��R�Y*l��R�
����AP��ib��%e­�UPR��X6P��)+*ThVVUb�H�����&8�%AUH�h�m
+*UU
�X�ł��!Z�U��S-Ĩ-aU�$�ʶ�*���QTX��
���b!��X�
���F���D�"�$�����W�{����c;9,�|g:x��d.F����Gh��ǃZ��Zj�F늝��5T��{�<%��=�Ѱv��.��:�yQ��Z�8�?n��l/x.�����P�BCHw�PG�V��ꭈr}J��H��E����R��9�%���
,Y�|�3��!ԙ����ϝ��X�s#�q�K�)�ַ�ě��T�noږ[ <���T뜹�R;:ܟ?k'*lBrb��ρ�hڒ,x)B��������p���S8�޷����8E}�6C�du��{}ݝ�'��k���u�����x�p�D���B�e�UeEA����x����[��oU==�r�g��p���QX4c�4pCn�"���x�ګC��6_�Ⱦb��*�<�G:���`#in��|7ZɈ�J�:�%�Q�G��H�S�b�8+H��/EuLإ'46��S�"W~S�޵9�%r��.�]��T"y긊!��J��_�����NbַV15ޔ�Q��v�g^^��yA���7ڨ�g�cq�%W�
YF,=�&(�����4��w�J&SK>���1pe��؏b���G0�.C.�!.nC������a��E���j}�T6��S6�o����$�puQ:rEBS�뱂�����1}]���7�7��#����`f5u��A�y��Y�c�Z�o�a�!YN�쾼���l����N�;)��b�*���f48�w�e0kft/s�3#��zF����L�2旕}�1'ur�����lQ� V�ܬ5�H݅R�RVmt(Ay^�kEp��4�S5q�v�V)Se@~}W�]�G�]5b�ޥ0ϑ�'�z�����Oy��+ɺ6iKe%����D���{h����o>���ǩP�q�=�X��9R#��/�)����9l��B�^W7F�Ey���<+e�GE�V�T�O��S���؇*�h����w�x�=��TǼw�O�&2_?:.5��kR�GJ`_����w�Q��o;�1�Ц�iD�E)Ut2\�l�s����3a�%��腛-�r�s5꽓��(� 郆2u/��������=+yQ�P�F7W��Y[$�*,�|�����wyc�,zJ��.|����� L\qP^�\��+t<1����,�;�VƱZ��~l�j]��R3C`�d���¨Oˍ
܊���K���v� .2�f#��*.�T�Cj ƥXk¸8U·���VG�1yvN�r=�EGnr�ͼ��3��(�:7d{���{�\�q�݄!;��}��GP3���i�����o;u�����hU
���IG�G������Z�S=�Ӝ�`g���,0�+y���`fnl�;7���u�۾6�e['��ZA�.��.*�U<�AU����T7a��%2�;�sCQ^��\]���M���O-��3$����)\�3��^:C�G�Ks�&��t<�B(?{Xħ� !U�K��O�>���yC�y8�h�63��1u�vr�����������;�h|�\��7t��C����j�m��ظ�,��s�9�£b�����Ǩ�\ 綽ǐ��9Q�+��YpߺB�ݖ2�����}S8*�"�x�TQl�_�ҡ��{ɑ&p!0)���� {��?��.��v9�tћ�dl�r�>|�ۧ���Vm��E��*E��xf�mx�[�z=��%J��F���bN��ʫ�zƃDS��d|.��b3z	:O]�Ϲ��{󹭋S
T�R��"�������|��V�OqIr�u��n�t���X���iKWB��~�Ϳ���"T(Pl���M�V�x�0���.u�EFM���xdÙ�Y5U����9�U�}(����y����eq��l�<���=m�	N,���8Z��v%t{�w5���R��o��޴��S�j�_^�5SZK���*yz����#���Cr��i�}�hMH ��Qf�:kG1�̷.�E��� 4�=}��tY������ӫ��,�h9��B����F������Ч�F��{��IB��S�Q��yب-��4�I�#{���9C��Xg� ��!�a�C�r�^X�{y�yF�M��v���y
�� dQ,���\�f�U�(�F[���Ѝ�kz�m�|�H0ŵ�|n���ˆ�5�6��1*�|�ҥ��ߪ���9Sg,�Z��jZ���T=��h��P�޿}T�˗%��-�v�,a�K��{t�s$��k��ԫ9b����c��1�;��&�����b�#7i����ݻܪ�������'B�|�åu+��#qPo�X66����"%�����b�OVǾw���^�6��Q�J�d��AxO�*���eA���V���4gnf�ŵ��F�q#�L}�>�+ڟ�4<�����Z6)��PxI����i���j;��N��J/:�[�A����x6v}Al��֙��V��P�A�	�C����7�8G(�7��s�Y,G)�>�\ dt!�\LꞳ�=B���$�+���Y��y嶟�L�R9~�Y ʌ(������;���1wv�����U�-'�gX�ZP�=ع2��yW�.j3����2^m�(U��m���������p�z2�q��I桻I���g@�fdⷰd9%�u���eN�
�RڹJ+�֬Z�Pi@��g���N�fP!�Vu4���_�#C�c8��D7 ��cc<ݝ����}(-g�z5_�����V�ڭ2��Ƕ0P�J���<��xC��N�3���.��$�p#��%�pI�(���yw
tlSxd^��b�[��/u���r��u���A/���9VD#<��&5*�ui��-59D���ը�8%KGKp��Q;�_ZQv61���!tWG\�3|��*�T�E�H��!b�8��b������J L�%fw	>��xe��\%6�{��_�:ٕ�:
��F�V:�Fׂ���y����(���X�)�,*O�Y~�] �:� ��Z��v��k�����3��<c6��õ��3{�{J��0�ymS:���}�c�C�1�+�1W��A��3/��R+�����7���.<Q/��=���<z�*������x�]1�n�b�'&��%����X0��
�ͫtvK[P?�\EMU��l�,Ⱦun�W�Ժ\{V��=���v")�϶˽u�ci�_#�4ηo�_�vL['��n�6R�zd]}��F��-����v�.ٕ&���Ů]��ۣڞ:���	�D��O��i!��$V'����)�����)׌����r��g����|�|:�#�f��MC:�c|=wx�XN�
t�u�正0jZ��
`�x��VFڐt%iL�~
Q�ց�wfI���a�\�Zg5nۣ��3�K�+�J����M��}���	�Q���Jn��'�.]W)0&���H�;t)e���4}8\����ZU7s�!�ྣ��{��a��>ː����\�(�i[��^��n���,�j}�J=�]6�h;L�(���&����X���%;f�̔������uK9uۊ�3��U�.�����rkU{`P�W�
��F���5�B�:������5�ޏ
跲�n�(�ix�c睲�F*���*�L��RߢF�èV��x��>��1s=�Ƥ��s���MR�mF�y�cԶ+��V��%l�������J$��>�{�Т:�m[��{�/3��s�7A�������X��C��s>����QG�BN�����+�܏R�1j�4���+}�wT�R��=MHᖏ@��:�
����Xz�ѝ�F�+�V��(n���;n9o�?C����y%ӷ��R�N��e���{�;��T�{�Iym�o"!X�/h0����6���O�=�1V�B`�t&��v���`�˻�uՙ�k�bQ��gu���ޛ�K#�quA͵�����᧲o29 �ƣ黼�U�����ŏ�c'�����P:����鳂�����ʐ({���(��r�����i@O���ٸ�~l�"�����&2�xS��[����
�3�qo���QN�V�āQ˨��N�_��#mT���wR&��WI^��Lyq��y����n�b��19=�B��~�蝥=�\}��=���kpp�Է�|��c��N��%.l������Q���z�>�n�wHL��:� ���./�9D�5iQ=�����/b���8g6N*��:B�YT�ﻅB�*<�ɔ"���6���+��Rŝy�c��vIh��"	ŧ�d��71������Gl�,o�38w��eƑ�-f�#�5Ӄo%׫��a׀���J��X�5M5�ٞ��gͲ5����w���g'��&LhR���~[��&�|��/��}S9QX�m����=�)���2�5�����"�U�b���h�ȿ'���s���dl�B���# �Sny��+m^N����jq�7���A.v���!d^��۫*����U�l�Q�Zj��%;2|� ��]ʶY��wk�s���|g�ͮ�H���0�����������x�S���9[�}���I��0�;�{u*�h�erۜŵ�lU�:�b~j��y�����x�������ٸ�Yqn�vN�6�T��X�����t�wk�nKn��4��Rvߏ/�Xǁ�'.�'������b|���SһҼ<mh�w��Y����j\����9>�����>,m�g�|��
��S��*:=OFr:{�Ҁ�g1.9�u����|lvJ�Y���Sf��P��Uk��Q��Qc�g��?Of��Z��1�kjg�9�Y��=O9��>��'/�iG;�����2��������f ��Y�)e��}E��C���Ӻ:i�y
�>!R8�\��겈Z��'�k��K���Y]�����.�����k�2�r�gdum���4~���B@��J�vv�kVR�r���l���T��cVq�@�ʅۇ��_��\e�}�V���*W��̗B䢯z�����y8'�۱�0�|/�@�.<F����ڃ-瓵t����3w4%I���=ʔ!��� �(�,á�~]�~7W*hz5��x��]�R��5���w����s�X7��e�`-�c9��tw���D�]Xxe���������Y̺u$���m�w6)�z40uc������WC�����&��Q4hr���x��mc�akm�{�]��>�&��3��kF�<2Қ�*W3G�O)M��O�F<��aQӗԸx������>�	�=����,OJ�����bU�>sD�*H�{�/qv s.�U�q�a������I^�����Tt���|C�(ì��h�v�>�!�ߠ�w�юop�1���_P[&�ӛ5���hE��������ky]WHP�Y�=	�A�H@9.�#6TC�o6,t�8nk��.��Zц���^�orguz}>ޣ�iY^Le!�8����Z!�q��*�Z8���T�J�󼳑I�W�;1s�~lYµ?G�������|�ޡ�����tFZ�:��y"������D���$��e�`���F�XdY��Ɓ�bs��G8��|� �u�1W����w�/�Gd�~SC�O��[A%g�����b}��]�X�������74��M
�6��O�Etu�NQ�+o���:��4����������Zى�]�����J�E)��jB��5��g�xs;2��f�|-#t�̸�O����ܹ��VC��DxZ4~	X�ql����:hyR�-�ٗ}�C`g*j�;!r��
@�vW^���٭�v����ї�+I�.�1�;a�]�W;бJ�%�-�[�rɿ,Y�����m:���u⡴�*_L!�N=���u)�[�4(�ޛ���9X)f{��������N�.�U�zE���;��Ļ���>4���OsD社љ�T��.u�9<r$���p}۔|j:o%AyHZ6�6wd;
�땗B����C�gnn��5Xz	����(R�
%��=��!���*��Ϯ8wB�披ۯn�֪��:Y�w���"�S�	�fՃ:;%���"�ơ\k2�^_�>�"���[���$n߻v=�b�yw��_G����bڅOs!��*y��=�Xg��mv�=�;�^M�+"ݦhƵ
�轻����0Ls;ĺ����q~j���[z)��.�/	��:�~�T�����/Z��]z�ED#������dAo�����Y%Nّ0&z.��%�ΤF�َ��[[n��dfe�B�2�sp�E��W:���]������]�����-�W%_M	�a��%��	��(�a�0�����:�Z��N���7���>5-�g{H������Z�;ޥ0�F���7���VV}W2QQ��3o�]p4!�eq�K�����c��ط�/��y�jd<�3�r�ȬY3tn<bݡ��$��g�:�y4���v='n�A�ؤ:�R{��kF��.�Fq�Y�z�G'3�Ρ�8�t������
v�"�����,T�3��,i4�
�$S�ڳ9}7�C]�{��9j�,�g�Z���<b��K�:g���՝843D����WVqgp�G/-��I�2&f��LM��E��p[|w%&� s�Oq�Ud�n�t��{��}������ A9 څ�s�Wnj�iјh٩BmoN�4�A;�u��ω��E%v���¹���z4Ic
��	��hT�i*VHWT���.N�a��e�w����n�	����7b��:[z��Ԇ��yf�Ӓ�U�)l/lV�쏳_+{N��b��o#�*A��r[]���X���s&�ku����R�1����a����R�l�ӟk��r���b��I�r櫛�I��u�[m�Λ̻�T��Y���3/r`�ǋ�#2c�j�����R�r��mЙy��ll�{{�rc�ޗH���c�2�4iݐ��^K㔈�����e��i�܏�+|��Y��9��n3$6��x�3Ov�q��.={�qjxkcv�I�7b�[�ֺO�@Y�f��Opƍ7Ht��}�'W�[p�9ֵJ�6��@��_]��ٴx�:�����ڻ���x0���O��i�nk���hP������^7K�h_m�d�6��朝8�z�[��]:�U��:�er��ք�򘂬����u���ZwK��%�J|Ղ�ܬ��r�f��ui�٘y�H�N���w�3����\��-V�c bbW��m+wF��m��<�n�EZt(�A���n�n���9j��#����t��Ԓ�Kŕ��7\n�tX�� �<�'i�ٴ�Ӻ�j��X���L�����1RZC���q��)�.y�;*�n�a�S��e~��Ӻ�Q̗C�����0��v!O,�Z��h����a�֫�,@=���i�q��80�q3�Zz��h�kI}�>����^�+q�s�E�����</M`�z����Y$Rp��D&���K̎��\WE�j�8SS:Y�r����������G}�P0�4�[�8)�9�Uv�.=�b��M
��\qZ��ҡ��^.�{�$Lޗ1n�����6���"��M�3:Tw=�טo��']�11ա��z����fu0%r1$�� �(��Wi6��7���Ǝ�tK�epbwM���l�]Ge�ᲡpɶNwK|�J-�6�-XVK��Ql�S[��RF��1��ά�4nne�H�-&v�5y;R���_gu�/j4�V�㥓�6�P�u���*2e��i���5gq{��*o^R�Y�gW �I�%�3����ru��+)sq�Y����b�(���Qә�w�����7��yu���"������J�V*(�X��YTA`*�b�H����5��@?$���AUA�
µZ�DVE �Q���E���b��Z��iX�QU`� ���`�`���j�`����E�VTX�ŋ+�X��
Dej9J�±���ȫ,*KmkX�ԣ&[YY��VUE"��jF�UL�1*VB���$R*�q�,%�jV#1���bȱEUR��E���%ERc%�%AV"
ֹaXbV�p��m�DT��R9aQV-����LA�YP*e�ƌ
��d�Z"	�b`�CU����]����/��/uڤ\��n�A$��;���r�T����8޵�-'�m�=8k��jد#�EDc��t�:2wr�V�6�7�5q�u���Q�p;fo��o-���R��6�����Ѱt�n�����E<�!c��bp�f�����+�6\$+e������R�x<����VV�2sp�Ǹ�m���X�|O����H�b�!_v�G/�HoG��E5+��%���L��R�R����E�Z.�$H��C�S���h�Qd�<8��%����%�/�FL�m�����ٔ���OX
K*�$<1��XP���������c�uC�t�5W�ŷ�akj�v+��_*�
�]�č��g����1�����?P3��I����7|�9zofԨҨ��N�_��d`�j�MP����O�2F��7CI�ٻ�By�\ɲ�x��:#f�X�dS#C2�"��]�z!р�gM!.'E yN���ut��Q�j8�cl�)�
F'�n�~A�XP�/}��d�x��С�H똆�}7�r��wr�&�Ɣ���pVS�貕�q��e!��H��������,��� .^-��9L6�3��T�'qe
�0��l:.�yo7��}�I]�M���
�Ս?�2#w�et/1��ˉ��΃w7�w'o���3SW1��1ή]�ge�52Q�2L,3r�ۧ|���^Sp7��Cc��+������|��]�6܈�D�";����1K�g+�ӳT�w�B��G��մ]x�f&Y��[��&6e:���Fڱ��ģ�0<j�B�svf]�>Rxj��ҁ1�	�Z���O!�~J�8)�l�4Yۑ�rj9�2_#m׌�xUՉ�M���/�g�3�=g`��[���Z#oi������]�_��}Z9�Fo�g�쿄�B�e�/�7Tv����:�r�zqK.�;�Mz�U!yJ!��l��,���d�6�jy�D�%��)�Q��̎�lr1s�.�����U��b�<1>Rib��:xC_Gu��{<���a<�cfI�
V;ϏX���E��
�I�SH�|ƕ�t"}-��K�(��N�-'���<x���*����	�:����@�D|_?���d���h���F���Ɓ�`s�G�S�!�]ٗaOF/,CB�8	J2��d��Zi��F�N$�*ݜJ�[N����D=WG֑�Cn1�b�ڹ5[%�M಑A�ݛ�)�(��6rZzj�L'Ӳ:+�zY�_�����=��vÃz���٘Dj�s�pЂ��/�%L��<ce9�5��&���BZY2qt�7���Ͷ!K-vgs�F�,�P�B����Vb�,#9�+O@u��V��#��\����%�'gt�+����g$�fA��g&���{�����#kc�����d���W���X�rB0'�U+����[���aj��O"�������rxI��w��P�>�X�o��H`5&�+�P�@��W꼫nNҫt�]���$����͞CxA�cp���S�LN��CY��[��v�e5[�2m�&���kqyt����P�%��Xo͝��|"ZY9�ۘ�P����*�M{��)�h].�HP9m��V�����h��)��ޗ��"37}eG$�:���a�oC���hP5~E�	����f��.��}��N]�m\<b����ݧ7(�h-#h��J�����Kc��C�'s^)Sj����{Ь���'j�����7��ƞw�{�t�xk�VW��xv�,î�,�W�{�Lr�.k�+r>���9���ݙq�sg�3ʙЗ�=�@��{if��.�;��q�H����}	����|ZЬ���s:;TaOn�Mq�bp�ͫ��4жu{��B�@@Oג���z�ܬpc�n�\��q�X��{g���S���C��f���#�F{$�
�ۏ}6!w���WAdcI9V��{%(���\D�Bq�A��1�t�=��w�z��p]�jq�=�V��
z+��!�ap��V����p�:	�'���d�w��>簈z��*�>��o"�^T)&�T1�ʼ�����R'�ڏ��v�H���W��YQ<���O�qŽϯ��dI���Ҥv���!�>����.�lƌ�sB)�qM��V�b�~����NzP�@��� �8��������=�^��C+�h�-�i���A�J�p�I��c�U��_�8|k����^��Շ؊=��PM-D�y�ɔ5һe�+ڙ�����o+�x�[�]��,�#)�݅J�'���Q
#�fj��eg+�ѱ�
�ڌ��hp�1�O�g��tM�]�i�G�n�ay�j�fc�,d�H$��.�k�U�&[���ǘ΁+Д����00:`�	r�
f�y��(��a�gr�F��V<;�+�^��f�C�w�h�<�]է���\p��|�罈p��lXK}Kf`#h�ݓsX���W4��q@&#W�������]!�
��̇$8�UV��Q���ӹK1iɦ��w�f��u�@��t�Mee꧆ԅ�v��ӈ�<�a��'�{^�[ޅ`���;V�<p	���oE��z�����$�|�ߙm�+���V�S�����w:�؍ͪ��ysǟs'�9ֈ�u��J����,��NU�s�rPWl^��Qa޵�e`o��#Qz�euM��P}Y�ȋ�ݍ+��;��rj�c�U�����ѷ�.j��\����~�9�H��8r�4E���z�ͤtXPjy���k�A���ETS��̵4c򠆅��H�Ք�f�#�!)M�h���l-J�'���9G֑�ۍ�?:^�S;(�=u��ږuy]ZbHܖ�s�9��p�,�����)��.ݑ� :�T!�/f��5�$�&f�M�f�O��S6�( �M�k�ut�uϺ<X��V�����OE��49�9ѝ|7��LU���n�rWuӵtUPHȮ�H��U���Ž�]ӱ���OY�U��f^_[g�H��`ls26��o(d1�ar��g��?/��}��2�8>�B\H��$4�L�N��8�;�ٱ�V���[Fxgr��|2�FH��n�I�ȇ�)���7�f��T�d��\�A��S����e^P�掕De6Gp��1�#;.8�q�m희�\��Ko�JQ3��U45���³�yo���՝]�bX�����oa���{�}4�&>��:�\�[�A-�U���<�
��3{z ]�o]��֢��`�Ao�YAkZl=��-ʯJ/}+E���Jz�j�d��]<�E��y�ojW�^�oc�٣�yS����}KkZ�h��q!�);�r�N���Y]q�!�l�Eߙl�9ٸ�j��v��_]�j;�����y���������"5.;E��}��Zm���b������f�ޜ/+\��f�'�7��oC�z�:u�E �����sUo�UF1��G.=�;{:�Jھhb9�B��|��q��SV�!�rC��vw�Vx�QwΚFu���O����rD�;�XȽ9�v]�Hr卡�Q���
�.+·��J֘r>�^��?{�yU�]8T<դ8��Mm.���t���⥫�焽�z���ސ��9ip�a�R<�ǚ[�Aq�q�d��i~x��	Ĝwp��q{�M���OEb򠆅BU{�)L#�w�M�?wZW��;��[n���z��*�����v�C�r�
/�w�{��u�s���;�_��e�����iԃ�w�����Ua֚3�!�4�
 d�z��}��G����I����t)8vW����%��8�e�����h���+�ऍ���Vv\^иF��^olEY���͌A8}`�T+҆�鬵uyV��J����+S�U��C2���]	����|^�	U{�<�_�Z����.h�шv�3g^�TFW"��:iS}��T��*�����AwV�-,37�z���|{-d�h�:���>�*3dB���ݜ9|���o6�d53�S�s~
��+�Ҭ̿}a���^5�l�}�J�A�J�rW��f�O���9����L�d��mfKX�i���h;H!s;4Q�p���ŵ�Z���{w5\�o�n��˞Y�HP9m�	eykZlL�':�����T��T�J�~ܛȂ����yYT
X@�C1�W�4��+4���w�5��4 ��u�go&�������ݧ7+@���ha� ѽ▸2ꋎSM�š�X�+6-^?�g��Eb��F�x+��(>�I���TF��;�1��5�������S�=`7�N���uV(N�nR3��'1S����3�TS����-�li(��D[k���A�E�S���gj�ٛ��n.���[��u�)3t�^�ˣ�����xy��.9�����s1V	�5,�S!��l	�y�ej����c��z�r��U�|'��e[\��N��V?*{UNuKD�;Q^�t�Z�wP�8!�iLE����i&9'��2�(o�h�qPz�6�9V\��];�Z䵙]+��rr�<fs�u��׵7e���^^8ʧ��G�
�D%es� >�b
V�m�.�j�c�p��q�.����F[�ԯ]�4+��d���N���%w��nH�rWQ���t�E�V��\v��zѭ�=6�R,d)���9�.K�S��i�NJ�����3�L�=��]t��Sh��g�8l�B.�D�Z>#O�H8�(k"k-c�JN;�'Ěr�o9�,^��G��8��)���A�|-�2�u�2� ���ia��t4��!�XVQ<6>wnM�>�c�g&�ʩh�E�.�]��9ew,��a�A����U�ڳ-�����,p]O��ry�;/Ƥ�����3����~�	o^�'ȋ�0���=�gxM���WK�Ug�c[�����f�����S�wJ��oGn���Y5&*��8��PH/�C�sR�xBz��׳����X9��p�ڷ�y�#s��t�%cJ�m��Q�;|�[��e�,��U��E;�C=s�㜙+-���p+~��ZF�W��ˠ�m_�,v�wM�͉���SL�|Y�5�\"b�t"�}�QLt�8�+����*1j��~sQe�0x�A�]V��hP~]
86m�#���{W��]���u���9:�[���{���]5z�B�M6�z��Y��P]++����A���Pj��JgI9k���|��C����:�im�n��+��':Y'�K*����<��&/x6!����;hS��W�q<���T�l���3<����Z��~�8�WM���K���гӝR�";U��8���7�3<J�?�������*ҩۊ��K�h�U��+��xo����ؔ�ͮ|�����*�>���g�r7Ԕ
�c��9���Z��o;���~���c9�)��!.&S�p����nc\u��o��O{9�9	Ct�e��GT�Rс�=���اӄ�g�O�"������| �>M���5��Ro ��Ҩ�)��)���ފDͺ��׫s'Q;6�O�4Z�����Mfwq�^]�.�>�!C�v��Ǖ��/	^��>{K���E�,	��0b+��|����힯��^
~���uo�2t����4ْ�n�5���qٍ���Y�DF�����jK�j/�J�C�V�L�Ls�GS�vR@�C����N�w`\p_e[
-���*���ؿ���\<&H�$~�;D,��gL��B��κY���B��m��&v���[81�wt��*����N�}X�1�iiJWY�x��u�׸���ʷ�9-�I��%��K�^FNƊ�;�KGR�{�k7�*R���K���̓Zկ��n[\��ם�S ��ٱ�f����FJ��$&ee�ÑҦ�ğ,ڳ��*�v#M�B��%��}�SJ�s#l�O+|�m2�u�B�E�݃9�ج��#@2CE�\,��o��5�EW�d�{;|A��|*ٚ��͝��\�/M�x������W�kb�D.�Gb\ 9�8�P妑�o��ױȖv��fhuԹ	N�t�C1�H��Y�1�B�D85
.L��˼
!��4�Iq�<�[����P.���vD:�|���KѼ�o ��x^��6K=%�Z.�� �c��[�U��-E���Wa���N.��V�X��ՍtZjKm}�d��ۗJ�g �(4*�\�֩��ݾ!��gKE�&��mc���i��*�4���m��r�kE�Z�s�K��2��g2��7�j=�ˆ�<�;�{GCD�w�X#9��G�e�G@Jem�-�n��� ��Vkks��c-�.���G���KGy�����M��Ϧ��pε��ט)�6�a 9�]=5�M�� ����o&�S�c,�`��c��M������gZ���4 �v#�S�g1F�6��3*�8l�YF�S�e�!�
�6���92��A���Hk3%��$P	�ζ�k&n�:�gB4c4��-)�ׂkl92>�Aɵպ���uʽ V�Ǣ�#��β��:���Uy�3H���Տ��7�r�:t�'���}g ��[��k��ʺm^,+~ʽ�m�/���m޺�н�
5j�1�
�5�[SE�ϯ2�I
�Np2�E'��}[q.
�s�g(V��Vܜ�f��mfI�Γh�:��5zu��2��pξ5�N]kF�$*gqc����kR�,Z�7z�d� 1���"V�K�ݶ�����;�gPS�ۭNS���p����p�lf�g$mmb]��S^�s����hf飳��X��^�@e�/2��N��В����Ϫ���;;I*P�fj|��z�y����� n�"��{�jݦ��{�r��7M&��u��Ft>��w>�=87�Eo6ZIК�7#dC���g Q�jOi
G�U�*����o;�D�40�O7�vmN�����Se����gR�1h���e��㾤�aӎ�M�R:x ZΨf'�Z����B�z��,��/6���x�t�si�I�]�V�0c�������Kc��z�O�v�G�^oK��)���PE���k�|�����ߓ���,*����QKnR��`�3X`��5��`�L���f	2�ƥqH"�`�AmiFBڵ
���KqS�1"�nP�*!���RE��\C2�D�1-2a�F�Z�4�F�����i\jVB��Ej�ZEne9aYR�[s3 ��VIX�J�*)�b��JV�&2,Y�E�UF�,,TT��!DX�E���i��
��+
�@�QIFTdV��2Ȳ(c!RV)r�
��ثJ�SRR"4`6�ZX˗b�
�P�)YeH�Z�-�maYR�+U���ʬ�1lj��+jX�l*8Պ
�1V��ƱZR�-��
��6������T�\ʘ�
�ԍ�V�[YERP�V��[X�YG-b4j��,�*,�)������i �%�mwgm��]\�VnD]hC,��P��L�i�u�ްi�]Z{�֤��͘t�R��)8aT���:���� �$Q����ws�Z�n��9l;	eykZ^��h�|/_
�o:
�j��:�:x����N���!�sR������٢lTMﰸv���kڧ���f��p����V��׋C��Z.�-�μ��s��Q�讫�I�\�'%05tS�z}�3�`�֮6�k���gϠ���D��;��n�b-����f�+���6���.R:��X�B�h&�����GyD�8���s���Q]|�_�jݹ씣��͉:1��z3:*kap�M�΋����O�;%�J;���z��2�OF/$0$�[��I!�,%m��êz�KϷ���5`�n��{��"�2n9n���1�v
�V�缰������ܤLv��8���~+����9<�[���\v�s�ܐ����h��8����Y�I{}�0F�ߑC��͹�ۯ�t	�oZMf*�G��]��f�GKq)�*�QYf^!ٜ�E�i򥔍��er[Ǽ������i��Ҷ���Өz.�h�t�/�}S�y/�[h��ΰ#{+��e�q�!��w�;����	��:]�����L�3���ծ�+
�d�8t����IW9�3�D���4�D�J���V(3�l��H)Y�9<s�5f����6H���Ƣ��A�	CY��Z���m��i\�]��rOa�λv��\%�������4U憲&��p-�jJ��ص�su����z�Rev-(t���d�5k�|"�ZEQ[��ss[X:X�����"��CA�lXK+�Z�oof�L:ZC�R�_Y9�N�����SNOUe���У���^D/r�قYr�n��V�ĎM7��>cv�
�Dyc8]|'"��Kܷި}�,�����Ţ��l��͎ �l>��sҴ�u	���+LV� A���7ȷM78�b����}���T;�UXs�i���1|��Q7ll��.W�#J�t�ߜ�J�����\�q0����M����֙�/u�����v�s�:t/�r���6J��A����1
����u�e��t��y��%2�T������.��>9�ְǃRN�h���=[�un*�n=����Mb��c�,az4�`9����ׂ{��#f�Tv���as�P���7KU�|B�� jq�x�r�],���k ŗ�̷&l�MA�=�c��S�ץ(<٥���a���(�Wr#nE���v�.�T��L��.(~T����P����p�v�U�3�;D���DV]�o+��f�g$�i����א�DP�U���� �
�>����K+���@�ﭳ��y �N(j22ԇ�r�ݼ0Q����x��_vqѴϻC-�]-���H����/�fޝ�媶���6�,�A�=�@�t}��;�7a1T��-E��_1���k1]�Nmq���L��,k3[j���Nx���6Gv,%��6:3�uM	��5�qA8�<ʹ}�e1iq�nM����u��{���M+*=��oL�����r�[Ｖ��i٢��>��L]��V:o.P�������ZJ껽}��6�����\DR�	�4�n��8:�G\���Yft q�p.����qX��p{}ϸ�┗O-BǪU�w��8�	��W�Y�����d�E�Oԯ`멐��ՉwR[ܬ��@2����vn�Q�ӳ���V�)���I���\�%��������S��U��Q} �[�)/5�9�b�!�sZ��^'�{<��y��+ެ=�4�L�nldF}'�LWR>�Ґ��!�l����]*���FH�6�DU�k����PXeՂ'Z \�A��iq]��V�c�[�e�goq:�xQJj�o��d䧩C��U
4��4ҹM�Ҹ���3z�������n�����Sшr�:��<�h�Z�="�r�_vF�-��6+{�|����U�m�w��c�CB�ί	h٘�f�\�kn����[�r���>���m]1i6�?5�d��W���A��P���9�]/���Y>�8127t�\�K�������P�b�����5ou2F�6����F'�R82�NވubD�H��~�b��p���&L��	u��t�L�}�z��Lu����eok,�1�ծY��}�N.����ӽ4o�j�E��$�tQ<�V�o�w�+$��3nӶ�W<EmPO]j�ʭ���7d��⠥��-x2k����w3���G����]qߨ9��')Xr�{�Sm��}�"�����}�3s�5��>�Z����CzkmX����Ҩ�7j9Y�B{�q��������E��Nh-�)f\��'^3�o��B^q΂�xMk�HPm �>�,-�Mhj��EPz6kӘTu������K7�^s��t�o�HQ�Aߒ�Z�~{{4@j��iV�Y��&r�������|<�������>�� sR�����oc�٬���L��ʝ4�kj�b�����ڷu��7 -8�dh��-�g!���0VE����J�V�.�������>���m��(4��i87�X��،cx�-Xh��h�W;Ċ��X��z�ڊ��P�WUb��_^�njS'6+��y�Qw����1���ջs�*��9JC����^�J�j򼮋r.�%V��#�Ki�a��AR���5����Ai�H�L�s�W/���x�SN���i]���kn�Q�.�<��'�~�f_��0�F���q���qB��z�U��u��q�qfv�"���Mҩ��s����y}�V�: �3˒�nb#��}~��Gv?�[޺>m�j:4b�(���/o���{���p�'�8���f��[��}�=�@z������r�!v��3�(�4�T<^U��>��N�j���U��dK�������Y�Q��;W��
���^�p(66Ԏ�D�z�d�����<�]i���nvw�/�{��)��H"����鬵!�:��7:��6&x�t��Os��)��5P�6!���X��A�JȚ�V^Y-׃�*���l�����̱xr��"�p���^M}���QS@4"�덑���V\ZǢof�휓Ϸ��un�o���)��pgq�鏝	7���θ&/��^�Oy����u�U��xE�{{HP9o�g.~㷖O���oE�H�zy=C޸��m.4'0���[�.��ho�oW�oe��Ԥ}�G^A�������1���B��zX2]b�}��!V����ǁ�/qiV�)�9~[����{�(��>y��ktW�hN�{բi�����\2R�r�Lz�$�r�Zʜ,'�Q�~&�ڛjb4�-݃c9ImM�Ƅ�;`��3�����٣��������~��E��hgc���Kq��n0�[mD,sҬ2�qf�w��z`��w]J{Oz���7�tn���4^��F$��n�l�8�(���E;�T;�bWp�l&k2�]���F��&�J���Yƒ��c��U���°E^(���*^oo<���9�!�M.���{��].G޹<��zȘ�Y�%�1k�=����������(�y����N7a��0Rb:*g�u!�v�Q�����e_�����{V	Ωh�#�e=b6`wS�aedgY�{��Z�W���U�Y�"�2�(���!������%ȋ��9&�n���U�]��}���+����pZy ���R��#-=L��e��V{�_m��tm2;C.��0�{���&�p|0'�cU�:������k��O9+f���t�3�I@j�m��3�M�hD5j����NU$��h�eZ�(X���X�h#;A���Q�氄���Ta��5�odfN�oGe�v�t����h�0�̉壙�K	q��7-�Y8�vV<k��E�5ג2��8]c(�
n�@&�>���Ρ����)[�ĝWܮ�����	��uyv�<YTr�#�
	C�o�/���wa���5�~�I	A�\"������'0]�"�#�Hj(�ə��a���[���1Z`>���zvh��oҭ�S%��>Hf��z�`G�*�D���81��(-	=!�[�L)��U��We2/ˢ���}���J�֩c�rd]1�b�jV����oc��5�/>�EM;��Eh��{�-��v9ھ�t��t�;q&�̶|�nr\�~�G�����MҨ���m�T<���+�k#ڒ����[ɨ��m��q;�ӊ���+X�\�mE;�T8"'lP�@���7cJ�uh����iRp��͖K�=�v��He����|7��W��;>��W]w༫����"��4ױNN�ʭ���&�nd�o���R�.�)�!YZ����b#J�j��=p��i�n+Զ�~��ޘ7�K�/=��^KE��q�(���\�������	��o�"�� %���;v����6T���1j��d��F�F�{G{�}���&��=�!�>m�v���hT':�:<,�Un���[��~��#�`�e���}W[�]HI\�Y�HVv;YaԞ�޿���7�9Ĉ�x1��U�̉y}m���Wd�>ry�z�/�R� ���{��8㫌l��G�R�e<}���D]H���HOj��w���k�$RQ^�5��b��u�x�D`t���o�][��v(���Sn�-!���h2A��:+'E.{��>WE��<��-��+�Г��c2��)�A4&��Z���s�J2�~��������k�zw#gX�.���P�ť�-է�w��W�^W���<�{x�?ٚ�Q�+�ۼ�Olm p��%�൭/M���sO�D�,�ɕ�̝���p����E.7Ha��x�`"�z�4�3��lR���nE��nJ�+F,�cCOu;KHe��K���T�ox�`��K�c�__cq�*P�7ܧ~���|�L�<[^�;0.��ر���0�7tP|��f�[�&>�r���\�N���o)>̜�
�QU�%�܎�M}��	����ᝫv+)s��ۈ6F�\F�u�i��ئ�n=b�֤/��ӏ7]*�����^�7�Y�@����\'sJ���;��L����8�px��q�k���[j��T\s`}W�f�u{1�g��7�F��4��71�Ҹ�tq���n6�S��Nɹ�19$�6]���]r{ηC�e'�=l���(�#_���]�2�=+�A��Ћ]%`}�G��WWeO8�{U����`;�>Oa���=��X���V���U�$4�(c��j���Lv���Ҭ�w2�er���:"��4�i.Ur� �P)���hq�WY����Z;7����/,�v�s�5h�)�H������5��!֩�<������{�7��r=��C���M��-�j,KA�	CY��Z�WK���N�n�g�A,���xl������*n׵9SF���j#�8�F7[|;Q�4w�w�_l܄s`���^���f�hf�tQb>X��S�9�[x����W�A�����!3SH|�mh���5�юL�բ�)�u:�^-��;����J'�0(e6�U�Mά�h��K���t��;{g �t��_�0�ws��4�Ƿ|��z��#��f�䢶�)���m�))����K��n��7��f�{�jLS���.1uԾ�ս{�����&XX�-�tju���������V��(�*�l�gPXlt�	jт%Zq��YP^v����<��74�����_]�u�u6��7�/��Ǖ�	]^4��R�3�c��(oA���
�"����i�#-�ue�+�lr<����%�W��p�a>�N�kU��Ե���૟t�����Ɏ�tYL�Af��l�!���K��\;i"�(^�E�^�Ӫ�s�5��;p�*�eg·��D�V8_vkF���g�F�ꕽ��`�0��^�	SNDon��kc��p��/��E���)�kD���m�՛ٮ�:y��DR8�8������+�m]���>�R�����cy2f�:��ט�sk9)�+�H��;���:�X>��o4�ΩyV�ɶ�̕3Mʎ��:�����4R�q�#���Yכ܋`���7m��z6�Lw}fG[&T�1V[ao1n�'����ã����^m��;n��)���� GY�\�)9N�H8�Q���(1Yۗ��u2ua
�����vQ;ܸ�:��߹mn3���4��PEC����a��:]�k{n��<�b����:�w2��P��ţ��V���o�9���U��U/���C
M0;#�+���B��;S~_`;[m�"D�v�Ɖ�Ϩ]c�:�݂�}v���p��'e��q�g����k�z���;.�@r�J|��V�Ntn�U�K��#9@mj�4ɍK!��/�y.� 툘.,S���>���(#4ޞ�����4�N3]]�)�t \��X\J��)���p�*��,,��Lw�W���.�v�rqM�}���/���.U�9	̐�:n��6�x��m4�÷�<�f��g�5�B�g#�.��h[���� ��]�oM-�I���9Av�.�C����!f��g�k�k��	�i�G
�[z��F��h���<��x3��y���)�%�	&�o䋏�'��XY9+Q�#=y��J��G͍�},�쬓�g[!��7&����,�c��9���x�S"�ʛnl��|�ji��)�S>I�ǜ��Ҫa�%dw�����b���5��Ĉ{)����K'��Wu�ו2�;6."�+x%�J�,-j-�3H����*us�#צB�A�T֤R����㣪�vq�{������b��,�ٸ��O)w^�/��%��Ϗw�J�Y���kD���Q������[EF[`�1\�`��Vc\B�R��iJ2�*�E"
��ʙ���*�*+Y`�������KX�m��E�¤�aq�F���h��DIm�*[*�h�iA-�U��"�I���aQppaQKlX��iZU)e��ҕ�Kmees
�����L0�T��(�h������ԶJ1�j��m����Kn3&6؂�JV
#i[l���e*Ԉ�6����T�
ZV�+ ,R��-[c����f\S+r�+.JT+KKFQ�U��iK[UlR���4SJ�`�j)QJ#F��Y�L`������T--�\Ĩ�[Z�D*V*(�m�bR�e*�D��QĪ1r�*(��L�YRذ*�*�m�#e�m-�&0EP2эJ*ԨQZ����b*�Y�E�s�Q��qȪ̶ڈ�6�Ҷ��RI�按r���6��ǎY'7�F.F��ϰ��h��vs��ˌ�
�i�s�U���1�'@wo#}b�x)�\�f1������*�>N����)�A4���4C�q�K�6��ԺƗ5֤�]�"�� e6B�=�d����Tr^F��_���[6[._�T�ٯNaV*�]�>�olm!G-���bQ�m[�%s�{w)��,7{4Cw����Bs
�VQn��#5�\�0;������T�*�ŧ&�͆��|קt���}s�ڲ*��	/WI4�!%�oCD�*�l�ś���=�DA�p�մ{-��B���G5r��{*�и�I�E�i�ŋ���������z���xх�v��
����m\��[K�t�$�t��s�+��d^��G�o��8�Pj��dhU8�	�(��Z��_.���V��gh�(t�σ�rtJ/W�b��^T��8JQG�6V��j�t�F�x���2ԋvL�+��N�83��.��o����F�	��4�yWr�oq]׬T
���H]=�H����Y�w��j:������ھ����U����2��4zLj�e��袞qީ�d��d�5�n��;�&cŎ��������1J9���p�������n\W��/j�':��Gj�t_nhU�r�X[ġ_k�v� '��k9&�2����CJ��n�5nb:�\N�sk�n"0bgwK���)�Xl�6�H"��R���3E�����-n^��^$�vd�gzh�"4m#��˰�&Zǡ��w�X��_�_�^>�BP�3Y}#3��')Vc(�
n�LU�xc4Y�	�'������n��蹯6"P�f�݊���4*��o���g6��g;a5�����n��U��I��*���gw����]7O�gQț�qg�b	^�`s�_R�oN�>�sA�&�L+��;�Ȼ�0�g`�rۃ�����@��a���q��t� �P�)i�n�Y�Z놾��w^>Y]��N�}�Hf ��5+�E����b9h.1��5��q�Y��)g�_nzp"�wɿ�vM��_!{��.[�=����Ln��V){�v_���� +���Ív�G(>Bt����!���Ԕ�|�{gG( �}רw;3FG�--m۝>��iV<�ʎ�{ya��.3��\N�%33Q����ջ��nt�:�l�ۦ����u����rf[1������������P�3�b5���K��.�|7רI��7f"��"��<�ׄA�����C� Nء:�x���M�;�K�L:���Ȯ�i��7�_n��c�*w�2��Zo��!�M�w���x��I꾳��������Z�ͥ�c�q��ٗ`)qX��Ж�Y�����v���`Oi	-µX;��/�=��������G#Sl��ȱ{-ʾY����;�zg�$B�pcgwJ�����g:�xm��d���o�C����}#m�qP���2��锸�*:*8�U+[��5�;�̷��]�Vi`�I�J��������h+�.$�k;&�f�Υ�9&M�ϡ����h3k٭�%*>���#��wq,�Uz=�����R���N���
v�֞쇣�-_h�[I�e]u�a��1����{���'%X��zOQ��ooE��Ĥ��Ϫ�Άt�ʏ_Y��z8��6�h1�hY���%��2�{��z���H�͕�ʰV�k_N��{:oJ|+��N	�4Z�8�����̹�(�Dos���B�����o4�3��z��R;m�a(oeY���5p�D���ݲ��Zf+)r����zo�ػ�\��(q�A�YAkZl=���#���}ϧ(����P��hM�V+*�|n�Í�5+Eጢe�oDM5*�ֽR��׳Ef�r��|Nչ�[s�ZF �8��;�e�kLٹ�Jo��唹��vkkg�z(;�r��N�q�o$��s>��[�G� �7I��Y	��:�)ힶ�;�P�S$*�ݞ1�����_&�l?n�Z[K�.����jێ�J6������w���as�B��I}O�x����k�s|��{�=ED�ͯ.�{ڧ{�r߯���:��)A�F�*�i��Oa*�L�fv;�Q���-c�ײ�V��bw�,;M��%�;vӊ�Ɛ�\1�Z��NN����?���w�]ֳ�@�j�@5��Ǧ��/W@k�$0�ܠ����R��na��!��v��ڊ`�:쎼�:țn�Ɇ�F�hO�e-�t�%$庩�i�BN(c��j���Dv�0�w�WA�!�#b�we�{V{9�9�u��g&ө�a�h�㊮�GX�k�1�k��/^[�)��;�V�O$RqR��&�ՁA�����S���H>+�`�k����{���D���j,M���5��0/S�Us;R�Wέ��Mx�u����)�:�h3��j*N��q0�
��[��`F?&5�5���*�aʢ2�+��a(u紪����\L��'��.w�r��4�����NaWV��k.[�HQ�lp\�хi�q�lX6��+�cs���N��4sF��w����/ˇ�n9��r�f%ڜ��F9��ބʼ�V��xX�{&��fT���I	�7�i�����sX�pa�Ƚ�"�qf�ru���zC`�"�0�
���i�n;�|�_5A�R���^ .��	�ٴ��zZ�2�Y�m^�W���TV�N��[�I��NF�l_M���ϝ�H)��q��$Y=..��A��'$őVѮ�+���z���R`���>�- �	\9��E�����!�!�6T#WG�/
﹓�����h������ۦ��,X��z�}����nWp��z�]����N�E�W�M^�ˢ��ww�`�T%A1yd��IĄ�	t�h�B9-+�������݊���4�.��uՒ̓����>c�:4b�4uNBR�<����9�R�4a�D�Ⱦ��o1�[��S簋�tm#*×�ʗ�T�W���q'n�������}�sl�j������t�k>Oq_���i���oΐ�Q�vf�VQH�����Z�N"0bgwK���N��8���8��{2wSTr�D�o[$f�HW�6��A�΍�Ghe�m-G�����S�fȬ�ŜIW��R�/ԃ��7��Z��[�
�1�{�6��ޒ��n�ܢ�)�Fa�\��[�[Pg�(k����y^�SE�G)��f�Ú��B���bؤ��ZƐr��T�b��ǩ��bU���?�[�t��O/���%�{������C�`�jȬ�Q(4l{���>�-=}��CX�s���_Ɩ>��؀;�5cz�e����/cr�[
�@�j��kL`Z�0l��56�V�y-J*[��2u{��P��� j��MdN�;��k��Ѳ�Wr�q=w�ܢ�Ҕ[i���_eLv�	�,M&�V�w��=�ap�/glj�Ʊ�n�>�Q�A�I�|V� ��i��b�
��Ɉ�zk�/�U�I�et�{�A�l8�6I�Ha� sRT�Bz��ϯg���<VS�I��Fu&��1|ث�ڷb����-� bL�>V�ٌ
x���u{�d�wj�6����V�PvC��Ղ�F������5nT�%���TV���s���n�7s����H��C�Kv�ج�����;:[���1����t�qɢ�9{.��G`��F*��Q먎�e5��nb>����vH�{C�tCl˵.+�lt��i�;ע���n�	��'";Y��X;��/�=����6����0-�� dER�ga޾�\�T��ΞD��6}�)#�=�m��ܯI\�k)mxS���~�v�FR�J�F�GF^K��j�Q�s;-�Ɏ�N ����[�e���\�S^�f�"��T������_^�X�^�F��ڷ��5ˉ�<�8sRU=b���m���V!�81�7t�+�<<4X]׵x����Q�JT��y�����r'�c�/8�c|0e,\2�*l492��ȋ%�sv1Z~�Vv'i8�5`��Rk��]{κ�~�k��|���c�N�:Wz����\�d���5��U�^���`���ڱV&�.݈�ɺ�~��#�S��hM7�$����>T��W"ѫ��oUΚ�[��b�׮�ʢR�r�]zJ����>96/.�?m�Gz9�umʃ�-���-9�2�Z�Y^Z֚�ۂ�]�f�����W�&���)1z�T��Ss��"��ƜԂ���ǻ���<[��;}�o�^��ߥ�{��SEY�Qyvyc��T��w��n:y��Q}�:o����mt�z+���� p�ڰgZ��'�h@��t��n����^|�P|.D$���ޢ���L��.z�Pa�\��{��m��o]-=��6�tl^��P��yO5����[�7by������w�E��LB`�[����커i1Âr��v{^rٸ#�ڈd����{qWe��_r��=8f�:S��Ϡ�l��ŁOl���W���*����I�Ps����.�}ηC�`��&�ԵlS�ѩ�J6�S�ñ�W�gtT��޻P4Z��R�k�|������k�8��tf�r��,��/����G�y�Q^��^CB���	J(�����n����uiˌn�19hA��[�����l�-����h���Kdv�q��D^�_-�y����0�*�LK����|-3 �J66Ԏ�qTd���X��4��v[�������_N�rG�H4�P�5D�N�i�\�}��T��\�Kv��:6��h��U��dC�5'�� �m�Q[fN%B��єub�#M(�4p�#]�PԢ}˂0�\����yק�Q:�s��-���٬�'0]�6ʬ��.�ń��\��^��V�W�?.��2��NR{������yv�͗�K��t�j/t{��5OibK���&o�wc����9�r �hce��6eg<��f�f����W�fK���+�.���.�����gD�`�w��T��w�έ�������M��[�/�KC'g0��u뵗-��!����[��l�9;�����?>�Z�{{4Z���F�1wJnt��p�M���bD�z�yE`-k5�E�t������3BwK
z�����38��{�^fX2�Z������-�#h��*�l�ś���X{�@+�R�����KK;�`X��_K���J�&��l�\�Ŋ{g���t�;��l*������it;�����QI����tF4�[�1)�ꑎĽ�[�����R����z+ͅ�G��*y
-+����ǭa���v���%�b7��՚y�{.��W�yPCGT�u)A���a�м���k�P{nY�B��	�v�Ds�E�>���r��/j����n�k:!�Zg���w��^�ݥKOqX�M�R6��o��as��oj"B�ґ����*� �CA[���w �Atx黄�EJ`]û:���]��cbI��2rIO��|���������s�9Brќ(U�����QI_N�%���`������ �Tk%�oF&�=-γ\f���[�ƶ�H��if�,e'�܁��+G0�́WՒX׈�F��}�M�ʠ�Yb�떴ⱻ�� ��Ŝh����F�K���:q}�1e�d��)�v�3@�}�;͡+R�8&��QsP��vB�C��{8S܄*;����l�;$�$Q��i53zm��ǩc���'+.�nq���m��u7m-�"�p��;���h���e�V۩m�5v_-�z�6�;�f�\��9O7�P��IІB$[�z���ڒ`��j����?'�r������_acSI����^c���������®u�z7����7P����$��猲��pW�KM/L�pT��+�{�������W���&)�,魁� ��v����.BإY�Q�ڝs]Bd��X\4à��a<��94��%'5�N�O�5�v��A��P;VP+���"[�mݙ�)䭱�{�:&� -]mr��G��<�t/Lj�����Ӕ�KZ��3�<�9bZ-㶻7x�7��ЯK��Ev���x��j��V&b����B�xv�$V(U���u	���J4�ZȖ"&�BW^�}Bv��+8��&a���77q���u����z�b�P+7F)C��%t�Ӝ�b�\5���wue26����5�QgV���UY�8F�}R^��Etψ VK9|(�3+��Obtx��(�ʴu�x�z.�ҤQ`\�j�]:�?Aƴ��Edن`��0��H^�p�{��)��SPr��+��]�+R,^���yW��L�c����L����b��F�b;՜Է%��2P���#EZ.Ja�3�f�)��W<�)Y�i0~ M��wu�����u�mq��ܩ,ͺw q@�A�](v�)v�JW
��oY��Hx���y�r�������RF:�a��F�P;���E���#6�, �0�X�2��_�.AV�}q	��7܅�cw�����}vd=��w���ck�˘�5u��"2�'�ࡩ���9��i�9��V�����.��a\�f��`�
[F���N����ov.� T�=[m�q+ש�%j�h����&4�6����&�]w�ا�N���|���J��V�[/6�Q�G{o튠��#u���.�	D`��n�])C��c2cW���8�]G�Ju:�B�F%�*T	��}�*s2��UӳT�zuخ�������)�����hm���}Pп�j��Bn�j��1|6�s*;�%G�w��w�����,Yۆt_ ��������H��gL뺻��R�Z�*ڵ�DQ3
�1̱s3+��-�T�`�.fe0Ɉ�QQKmVҥehV�2�1��k�r��-��ܹ��&a�lP�3-T�W2""�9J�#\Ƀ2��J�1Z"�-����UA�s00E*�������ccQpF�FW.�*\ɎR���h���\�LrƫHVnFѶ.Q��YU���
�7��bW)`�T�S�Qcm�mjU��q̖�F�EˎE����j$�3-�+2���R�D`�VV�F%Z+.R��Q��0P�Ҕ�Eq�UZ��Q�X�j�[eJ�)ml����m�UT�PmKmiJ%��ƥ\̆YU�*R娉�k��is
���6�.[U�1ƶ�R�k��9jZ�VģV��h���YeeZ�,˘�A��RԪ����*-��ZU-�V�kQ-Qe��e*#mն-���FQKiP��mW.aJ֭�PF	���b��jڍE�%[m��k���L�ls2+m[���բ�,[�fZV���ض��0����`�E[�pY��h_W3)�]�36c-�����b}j`��1�/D �|��Z+*E:�̩Z����뗓��P���Pv�;G�W���e|(qΫ��l��vW{�e{��w����`h����z4Ms�����de��rq�+����w���{˥�=�qb����6�c5��0�מ��WCs`�Uq���C=���J�>�]��[{�P�;Xg��YE�4"P�f�݊���4YU��foK�F[ރ[����aa,(\�8'&ڠ'Nh.pɋ2�~�wl��Uk������D���ߖJ����Դ�zvi��äE�D���ݪ�х�y\�lW:o��Í
9h;I���|riي\7B�;J�ۉ���L@�	Z]���}�Ha�ԭ���"�rƎ���'K�ܯo%1�E;�̓�v��J�\��bL��7��#��p�X�X6�q{��8�p�J������P썒.u�����*F�����ݮG��j٬�)T����]xf���֯i��ِr�He��t��p�����Ū�Hp��sU�}��b�kY/�ͫ���P�g�����ָ��Ό�d�07���gh�䋥\r���S�X���%#v����6��Pe��3]�l����$ڷK�읰9(�;��glC��s-��[tэ�eks٣�O�����'�5n×��th�9#Gn��i�X�'x���o*�uQI�YZ��ߛH���8�WE�e�8[q�Y����dT���a�0�
�9�)�#�0�V�w�����V��hV����:��1Bd���T��}���fL��v�ڎl��V
�%	<Q�c+�����8-�����=�E�����d�]q����X��&9"e<w��	�����k-_�9�:�c�W��i��U]�^��̭��:�h���Rh2>�CQsMaz&��R�w6����D�:�V�f��t�(������P�4&��|�T�"�yq�覬m����/��;��o���!�[�:ian�i���6v��������H��H3$���^W�[iD�������^ �a�ý��N�:��XT�oB|hÄ�Evt=�6xR�S���w2GV��C3������t]��:�����,8c�a�'��w�I���ܚ`pCn��5�T;AK�u��UF��~ll��b�U�˖�}������
��]���.��en�s����w�M�|p|Л¬VU�t����V�q(�g8;Y]OyU�&xެ�}{4^lrq�9%�e".v���]�*�]�������l�Z.�-�9����J�����^�������Iۖ�I�Ӫ�ce	.�M�SM��b���z�ڊ󰺮oaB"1fd��c9�.{�g:�в��Rj��q]��Gջs�)V	̍����]�pf�6���Cx�Ы�q���5�>u_b	Gv�?~�<��?R=Jïjy���賩����Sы�N^���j>��_��j_<̣�:�9�����z��&��˟s�{������;�FJN�vI�O�R��Cε�B��^�es>�����I��i(��m�C�bp�
��B�q����-Qؙ�(v�<�#��T2�|��k�2�WOǃu��W�ѥN�N�S��/2X�e��ݷԂ��{������tX=�G�:�"�N[��o��v��Q�a��Q��M��pJ�op|�e	�5)�E�
�bg�:��۷�u�ˁ�׹��2��eھ$Jx�C�4�A��Rj"��	ˣ��A�����ā��,��ãB���Y5��qpba�V�d�����ep�7�oϳ�s5��'"��J����w������:I\��2��@L�������;Gsp�N�f2i�q�5%�	l�d�3�ٱJ�Nv'���VP����-�)ڎ���A�{�\�`vQpl6��]W�(��m"�u=E��`���@��[���g=*n�>(I�Ե�0C	P�B�G �!���Z>�����Ɣœ��8~��}���a��@q�7^ה0@����s��%Ǔ�7��b��¤g��6���4Ε�d\3��Δ������P�.@��B.��i� �cDw��.G�Oc�Hسvܫq��nf�Cz��Uj4��V�+"v4Z�X��o��s��..'b��+kh�o_^t8Fb�zq]�e׾��&O��� �J�1�Hp��t\��gU��>]��*����vA0'
�HM�I�C*d)��x�Q-��f��A�����ˉ�"Ȩ��-��ix���1Y�r�g�/J���3ׂmӄ��\�y'R�h�gsjEK����nM�ǯ��V5��J�ec�' dg���}J���v��m�jk��)�Պ�64�ύL�7f$��;33��|�Y�~쮉lW�|�� "+M�>��m� ��R�x�<�~[{�4֙�F
�T��?>ؐ���(�ƺ$t�}��Ha5ˁ���F3��o�華��x��w]�d䷞n:ٕ���@���~�C��1e�54ݬ�`�L���`��9p�2s��t�*�*��V+�W�Kf_y��S��]��';���[�ecO+Ӑ���Vj I�P�Q�`�r�utu�ˑ�e3��6F�xV�{���^^�U��y����	^��&<���܈+�s��)rT&���+�-x�e�WF�WU��z�8U¶/ �b�=�F�Hñ�
�#)ũ�u���/�,��Y>��6x��%p0�ѹ����P�px`��ߍ�x_�k�x?�+ZN<jk��X�J���n�����Y�#�o�"h�44Cs8��ǘ����){��I1{�7���l3�������cq�(,oVF�vF|&:���w�����yc�&�]4�Cz��X+��l���F�q�3h6�孺�<=y��Ց��:����m�����ݩ*>7�	Ʀa� }l�l��i�=��,�-�����3Ar\(�2n�WV˂���p�wl�%,�}F=�ow%�*�ꑐU�NB̮����ciǨ���I��[���轚�f�{}Y}�}��~u[7{^
J��t_59��ص����l�X�HF�����>I��q�\^H���Y��y�qr����tҜ�lt�yX�al�D��6z�+ɯP.����������TOo&jJ}ʉ��
=�����H�J}J%	��r���d�}\�s]��vM�ދ�&Fq�Üy��
'�?>�-�C��*��V#b��o{��b��hC��>���r)b�Z��y��*09��pl���mJ�=;����d[�t��<��b1ҠB���w�n��U����O�U�J=^)��.����7a���{��b��N��n卢��QS۾f�\��|Q��}��9��&6p�e@��-g������e%��K��'���^�Ы����[���4U}C�1�4,+2/Cq\���X�r�ҹ�'����k���%{��6~���B���Ď�D����� ۑt@�V1x�f�2P�>��ڦ`W��拸�j�k���oC�ٮ�X� k⣮n�QZiF���2��t}H�p�5�.��N�����Ӭ�eU�dL˲��o�w��r�,��Y�M�z˺��%�·���؃��#щ�IƳ*
��Vw ����fk��U�� Y��O�<%�|��gG`�� �6��uug�����_B^0�e�o�nuߕ�JZc�}�PP{j����%2�x��D��h[��#a����uR�ϩA�Ƣ�ŭ�s�&8�T}j����wL@C@H�rS@�6�2k}*=S7�d��%'�:V�כ�"�dc�`�F��+�"�U�c����BWMÏjU0�{J�,:����Io3<�94{���G����&� #!�ݣ��nw6�!^�BN�P2n
c34X6��(�0�h=�~zsf��G&KC�� ܅S�O��� Y� jy� ��rDd��Y�N6N�7�=/��0鹬bN��[��u��^к�9"�N@K����,;���MX�ȱU
]�>.�d7!�qG��y��(;1s���ūp٬����.�Nn���Pc�P��+������z��^�ސ��I�(�f���o&x�f�w���*��~�smPFT��'+�թ�
�ArF5u��dB�{OrW���G�`���BxQnP�Ss%�Ĵ6uT ��xㅞ6��%�q�d����5�YwW[H�i����'#=�5�:֜��w;B<彪�p�wX��Z#PΪ��d�b�P��{���4�Tnd��㳁��I0���w��hf1)�A��A%f_=c�{}8O�V�J�������U05��t%������W���n����t^��
���<O���8ʳ<k�n�i����.8��9;	+>IVL�t�A��Ж�+F?�>db�枫rP��g*�|�o���mu�W��~�;<���*�W��S;���d�M�NLP TH!��Ƕ�B���j�f���ԡA�U�v!�R,`�DP�q	���].��J��F,�eC�4�A��uA�Ӽ"Sũa��UAp�cš	/�����{P�{ʸS-��+��!W��$����w�jHŨj�����l���[y�<D���]�/ۜx���Njg���v�z<���k��+H���Dψ���k��LȻ�Y�.�Q��2����x�W+�=0�D7�J6}��pQ�CW����G0�Q���xU�ǢU����l��;���z�v��,r9Hk(Ň�D�5^�|Ɨ�4��,��xϏU�u��	�l�q��|���]���s����̔��	b�v�ОoM�,k��Fd�pm0�L�u8�}�H$[��������|&�9��q�=]-[�}Z�i��'ף� ]W������-S7_T/��vЭ|X�ۘU����']��Y����v�,��aA}�P����+�)�y��E�!�ؖ�.|��EM�}Ȍ�ew���N`�,dvy��$tZ�/RU枋R)�������zq(>��p��K���\�Yȶ�^���TZ�z+5�hK��kɐ���W=*k��/�Ϛ��]K��|��ԍ��G��R����+mu�tlhC<V��˺>���i�s�8�y�u1r1�m���%0&c�)R��lqU��6 ��Q�P,Kڼ���Ҫ�$���iFfN�7�
讎�Êǧܮ9Z԰�Ҙ���W2@օ�����97�4���)��}vTܬ�.�����
��̨��3c��q$K��o��m�Z(���Y��O�^��83Ҷ+��^>�c"�Gh�%�/��T���	�2fa������g��<5�����U�@���E0;{��R�w��N�g���!�=���uf�YT#�d��z)�"��M��QqF�H�����)D>�eKo�)�λ�5F��O��pg��Z)�v�[ER�p��dr�������(0�'zpPƔ�g����(��zcGo�1������SLv�FM�
�y�����e���n_:ݜo���.�Z;ج��lab����c�;�����K�u�𪳓��J= N����¨>�"�x�h�u%�&'�%{�0]�{Փy���-�2���+�w��>(`>54���*{�°���j�W�B�@�e���ub7>���
#	�^�����h�\4${��"h�44k=�lz�RZ)�f��<�<B�o��>z�r��^��PXެ0���xLu���Y��A\�}㐬+���t'�Q�:���F�=�M��|0K}N��(�r�����p�P6��*wJ䣗�z`vP�j�K�U��\�d��,���B�[=��n��}k��S��:�D�z�9�,�g������k��v�3��w}����P�@�k�xV�=�O�*8�Ec�P��r�L{�N�tr/}��b��.,:��v9*ڞO��"l)Q1��;B�{\��mG$�(����s�Y�k��(auFˁ{4��E�;�2Tc��dN�*'��T(���B�����I���Z��#����WVP�����+L��M|Md��u8Ϗ+�V����B��`IO��IO�$ I,	!I� �$����$��B��$ I?�H@����$�hB����$��$ I,	!I�H@�hB��@�$����$��$�	'��$ I?�B��$�	'��PVI��k�f|�I����X���y�d������t D ��t�TB�(�70(�T� *�����̲2���"�SM7]ԕE��4�qȢ�[�.]�TZӎε��kE����CSZq��5�[j�͡IlA��$�6�P�FP!�gG.2�B%wgF�[kCA��'�[e[ݭ�$��@�NwR��%*��mH!N	�THQR:4��    i�JP�h� �� 4)႔�T`       挘� ���F	� �"��	J�       �{Ԧ�� �� �  I��F�SdLh��Q<����2����������>�"H@!�?�d���g����$I=R @��~`�$k�������A����H�!&!$ �R̑�H8�T�2E	Ēig�צ��9����~w��� Az�W����4f|Z~���_�A̅"�����������ij&":L�@ݰl�r�u�q{��T�*AXr��0U06i\�3`�77N��R�b:��y��Et90�#tkr����԰i�j�+2T�Vc�ǺM��������c��_,UlU���u�����a���U-%��Wlx�d�-�v�����[x�6��wpa�m�Z1jF��fV�1�ӄK��sWq��P���r��,-����͙��Jҭ��y�$Z�0��i=�h3Lϑ�� fi�h@�l5���3Ż6�=�)h�Y��J(�OPldp�7XU�����L�������9�(�l�%��d�Q�ȭ<�
h</�Q腝�`�Ȫ�eYV^�(�R[�[�n^�LƯ�q���6�f��3�M��q�����|imn+I�{X�j��G�Л�,@���evX��93���a�i������1��������K��Iը�-H��d�����]U���4��(���+�H�ڲ�\��hn27L���.���'X���K\x�զ��i���^��C,#t%�ȱm��.յX�ϐ����{F�X6��ȭ�t���u����^&d���fe�xш� �Ya��NXZT�PlT$�y�\��qE��L��)8',c�7u��x.d�khܥ���5
-�T�V����-xNfۏc�a�ˣkn#�j	��V��n����kH�B���e3[�[yD�Kh��� ���Q�%ٸ�FM�rVP��'/[�;�ˬ*\Y��5E���?[�W*��?���:��'S1S����(m�'S+R8�{uV�XUHu��K4Rj�`��`�b��PZ��h��*�Rx�M���N�ڴ�i���Yw���5�k7K��MV���@3j��Z���ϲ���5�Sm-��!y�e܋o�4�ZԹ!h�Ei���of]�XR�v3vR�-B�����mef�.��J��L�yuh�6�� ��iMEa:mH6Ry�(�\a�4��Ž,nč,`�A��6�M:kq�u>�5[Y��V��r:��+�f���t�^��w�q��{���m�1"�Wb�^7����:-��`uv�j�S�dY��t�3	�	)��NMkVë{��ͽ5,9�p�8��Q�4�v�*�u�^��s��3��@c��t�'��:�G�1�(H�	���m�����j�T�jI$�II$�9.oA�W%�#r��R�y3f�ꙵ� ���P�=��0�"鈸�P��1�ft���)&lnG/�nSgk)�v�e��tmgU��n�YX_c`l7cbۧ�4�p��9�k�+8�����*m0��f&�@������ř;��u�>�^kWH빗�&G�����{u|{��;ifF��e�5���d�r��BZ�:�sDI,����˼����]�D�u9F����2�AB��J���A14;�Υsq�r����'yt�ǅ_f�/�����E�J>P��ܼ�l�u�^hm�Y���Q���d��p>�V�t������Gթ+pb�\`�Ε%lY��]W��sZ��9{�n�<.v�ymݧ�q�z����e�Z'-�ؗA���!0��v�Y�yS�L����	���e���;\�D*���9��LI��p-�$S���bwY��6f�p�\����m՝�oZ����%,����^Q `���0�I����)���*��oi"^3���;ɪ;�.��Wj� uD3m�3z�%C9����]6�oZ�ثY�L*����}�M\㗷ٍ����\�o۪�kF�j�F��_M���[0�����ݵ6�ou��-�yҚg��{ G!��Wp������g�y��f�6��V���2�E���W��1�)�ed���k�ݡڣ�������̺Z�G�1+/@��i�:J��{����]�aQ��	Ƹ[|˔8>ÉX��E(�拄���y�jvp�ܾ�<y�&��n��X������x��<�]J������"�A��9-���C����Zؒ�`C;22�gNe˹�#1��G��V�ӕ��r*�U��;z���'�k	�ȾVc� �n7�B�&��d,P׊V=��±���gY�M������ě{��ְ�0)sq�J+BTrM�*R�ۓ�[�ai�s���р���c�'n<#�#��74G�ܱ�ԚCpU5L��Ex^��Ζ�T�G�^�y@J���;�-�fwI�6�qI��w*��:�����l�XL�Wp�����@��+2���{��^�}�zX�n�J<�3�Ӳ��b r첁~���xwk�����d�ņT'ۍK��߱�>�ы��G��=�;���$�<�Մ�쓇�:. @!�����E���]Vux�ߜV�s�M,a�.�/�l�N!Z�=��h���c��PY�0+��)N�M�0�Պ�B�hhf��X9֕`��'.���ʠ��*�Q ���ͦ�cބ� Q�:�O��:)�E��oI��i32���˳��JZ��?08-�J���OZ{ܸXӹ�O(Ao#ӖWS��vQ+eu3�Y�핃F�˲E��bS�_	z.]�P�x���k�v�i�/�l��I#g@�ٺ|��� ���Ħe���8���۹�1�&�}#�L6h�t{d�j�qS���|�j�XP��XѠ���@ц�a8`�3x�G+?t{�Q�{���{��B�%�"����b�S#k��N>U*��F���A��xdm�����b�u�λ�H�&E�*��h�a�lLL�X�Q�l�ˢ�d۸^�
u'����o�j2%j����ј4m�TU�t���'k-X�8�D�I.V��WP�d�/v�s��9�m�;Q}�gU����T�m�$�q�Z)*$7t��޴w�鋆�)������`��`������]&2@��_3�hN�w��X��"w��O���ӀRec�#R�F0�Ŋ��oZۂ�]�`�s/:��0Ur���o�xŸ�L�����`Nоc����g�RQ�]2��mS�ğ�ie�vm�Za�S)���1Y�c��7@�]������Fq�6ب2�+D�1B�Tc�.L.�u�|�����X�R:�e�O,#	'.�J�h�T��ckX�����ԫ�%���d��<��.���rS��#W�Q�����)�;�k���&�i�U����Tk�Vh3P�w��vG���_U��u�	��)O�M�Ѐ�.L�N曵�YZ�#�(�X�����G_r]w��4�u-��/���*ϝ^L��jUX(�W���7��H K�� �U�f���ePe�Jw��d�k���)�6$�V?����/0ܡ�&ڤ��
k���i<�tfaT��t�q!����;������Wufafj���%��݌ٲ��[]I�F�8����1C�d�{)�̳��B�|�$�U���F�N]�o�%2���j�+�E�pl�q�nά�6gwu�a$��fu���Z.��q4�sxu���h�(D��6Nx�D�������'q�1��M�j!�5�h�[��s�efd�+v����w;�)G���Q���%�O��ڶ��)�Ó	��{�qJ{�G&/ei�Ӕ��]�&c3�^�}%�\�I��u�MQB�)$P�#UR�b" ��X�b�%$X�DE��M]B�E"(�e0��
���Z�J�Dh����n3�#�L�3~������Zr�v�~1 r��(����@ MW���7�κw^�{���z�cT�aƼ�^f�}ŷpA&��B����+�3^Q�^��*#�"�:���p�Z���0��4m�˺�O�~mopL�}�1��:��+�G&���.$����g �X��i��1>;����S���K=�Ҏ<������k����ΐ���^[�Wp�A�侲�lM�۬�	��[ �Y�7)H��2{z���|�
�����.�f� f���6���u�R`�4��x��tA��d��Á�~g,�%�jӻǟ2�Ռ^l�A�����%��cp+���o���)�a6=tQ�Z}�tE�[T)x��&�LyX�~�2�w�c�9��ަ�y-�2*J�
M��]�z�{���t�zy���g���X��e�w\bf������uǄ�5l���{Ʋf8 L��@5����oʺ�ׯ�EC�>�'%wB`o���%Qq���g`n���+kۘa C�*�̵�3p2=�d�Y�6�K2���!
�ZW"��٤�nJ�[���տ)�3���=�$^�1�0���W���o���~U9"q�]���_m��Ԛ�Kc����8a�W!K�P�5���5ּ�Ϳ�8q^K%	��a�=�G7��,'��Y��;(�f���)v�i߾����3����m�<̾�7
��M=W]t���m�/�Gs�f����՝.�����煌��f�Q�O�������07�A�����p�M�@���f@�7�8G[�(i/��}�x߯����t�m����W��Z֧�+KՔl]�7��o��fǜ+�����Q�#9��ݻ�����S0����^�zdy~�wW�q�ҝ�M��
.��vh���Exn��c�ء��M�0�G�=�^^�ο����Զ{�(�8�D˻����L�
�4ݽ�&�z�'o[��L��g�V���c*u�j�MF^c�)�qT�ܡ`ۗ�I�9��h�b�Zh[��"Y31��opv���s�َ�u�#E�!13w+F��ed�fDs}��4&5əK�u�귊,U܎:r��}���������e)a ��Y���zXEu�ai����5��W3rb�k7����m���n2���l:sSrX"�q��9�Ĕ\֭�R����$��$FE$P��
)�HE�$?���g�ʷRT���}$�{4�.���½뺳��f������Ϭ��~�+8�o�����pH}��&���D�Z�j6hz:�����Vd!W�Q��Ws�rb�[���'#��d�=�Sǵ{^��
瑛|c{]^�[x.��׻`Q��~=�z��tC=vz�*�txL��#x�{�_EM:�l�h������,�
q�mXw���9'hP�׎i�p:ӕ=�DQ�^�2lwr��+�
-8�R����;��O���43ӕB��-~�I�q�����|ކ�2�;��M��yiW�;*Y���n����×v~;nd�i��ӳI���&y�Y�2������fܘ�ƿ'�8D�&�oJE��wL�&Y�^����uL��g��8;���y-����
����>ֶ�Jv�$�rn��Υ�3�w��Ҕ��[d"��� y>�~N��#�Zkc���O�����o�؀���5@V[�i�y)�n}=�t+*��*|�����~p7��MܛL��t� ��=������w1��|RS/��Eӛs��*w��]�{sr��K6�����0��.ݽT��W^^��G��叭���+,��zh�<3��@Qb��i�r;���x�o�f���n����;�/x�I�T1ERo~�e�#�,~Q]� 3'c�ۭ��g�3Ӎ�O�ĵ[��_�	�|�>f�Q�OK����W����=^U�Ma�9�ճ��q�xf��;���R}J�Q�-�gJ)�!1���^ќ`}���*��{V�my��S��l�<��Wyr@(�v�zՅt����߶Z�]r��TKĜ��Š�ܮ�W{׾;XS�P��Ϩ�4cH��4�O73�����(���?\y(���	k���}h~����E�
��'�y3���F�s7O4=w�;��C2�*���E���ߖp�v�9_�Y�_�2����mg�߆u�w8E�9�G��E�$f��Ma�u:xWL��Xu1�ԧ�S���E���1����PL|Y����ج�ۓ(K�,D��V��V�8�B'V��0eHJČ�f���k�3�[ﶥ1����D���gF"j���_N7��;k�-w�H�7���@%zX���ۺ9�M䳻��}8�B-��=��Iʹ&�I2�V�����w�E��5��=r�u�뮻�>�`xI"
D@YA`,H�P��E#6{��ϙ2��mD�T�4�~z����jt�ߝ���g��({��0�)
{��U���(���P!1���aXܻ�EX~hٮ���6k|�%��n�~���hʿfl�k� ��%X�-��@���ws�W�p���/��봛jh���m�!H}徛8�j&�!�I�{r�Kؙ� yhpko�;S_Y��5�x�V7�>��+7a��*w��AF�]����#I'M�Ԓ1��ڛʏCS*%M��w|5�!8��M�C:�'/*���u���K�͐�	�H�f�L�1����ġd���t-��`^��+�3��׬���,�r��06#�����Ԃ����U�����~�=�(ڬ�����b.ùBͽ�L�+u�ac�l�+Ƴ�w�Ɖ̪�E
�[$�^Z-@+���#62�S
�ޝ�{���\�\>i�^cb@��<�u�� y*j����L��/�A��MNѦ2�;ӫN_!�>�Yܔ���0���\�޶��P̿wv�ԟ����'u�}ݼ �GY˛K{O���|�mj��JU|�Z���UӞ`�K�h�ǡ��0�+Jd�B�+���X�-���u�v ������OJ̀�!�)�_��2I����j�е�3�l,�+��R��L2C���'S!���`m��!L	��iS%�i$�a���HkU RW:����$�!
@�Kd!�$7��6��I�����!hAHa'y�9��$���ā0��0�'���f��a�I � d��,��T!��@��q��e��e!4�-&Y!Ψ��M C�>.e��i��X��qX0��C0O�2�eaꕷ�����I�5%���3i�����$-����d��$<���8�xBd��M0�!0:@%��\Đ��2C��N�4�Ka��,���.s�[3S���E<�|�TOzps0��H��۹^��VG�o`�K7V�w�*��N�j�W�Y�24�H���\u4c�P�5Z��	Sk7�d�G�� ��n�����{C�M�˦|�t��]~֫'�n��f�呬#��3R1��Z���BF��cA玁�ۼ:�Ө��0��������W3���H��%8�Q����0�~��yy�i<Yǯ�k������W��L[�5�:�$�uN�^�/.m=�$-u;jC!�e���+Gt�OC�K!�����o���V�~�T��E�<�%��7�L	ݫ;%�i��k
����JMM��I,�-S璮2�(M
��]ep���[VZ�n���
�܍q3j�A�vw�
Vn<���\pt�u�u%��t��>������Bh6�*'0��`�;��J���ÇzP4��Ke���y�7�� )5�����ɛ��uu��N�øŁ�
�ۍ̊�B�9O5M\q��J�
��7Q<��dƺWD�ޓ�:�,��"2*��EPPD"�Qb��"��@PX(,��|��gu�_k^ի�_2��S���xO��B�"��~pF���m�����FP�Tg���fq�J7�'(��,��.MhZ��������*��Ŕ��=ȗƝ�^(�S�qs�J�0�&��5���)ۋt�jA�觘��9�)�{��~��.`�2�~���3^{�Sh{�ͭ�X����&�W����:��I�G�݁�_��
�a��m��㟫�I���C�<��ح����o伭���zN���5y�ލ���m��}��	��'���<W<���z��Y�#(�u�X_���nt�r�t%N,�3|���r��Nc�������3����2� 
��\y�oe�������������&g2PV�/s0AF�]B ,�G���^����KE�ԋ����� W��&/�OU��H�=�]'QW�O��[kVԆ�&��.�֢�X�7�b��MgVp�;h_����Â�gN^�n�t�����D���K֫3q�b^ff`;�K���m�w4�W�5���WN���Z��燍��('j��8=}���24�]L�J�Mf4�+��%�{�U��E<Xtn{u�X�(z�������i|}�2�"Ⱥ�|�b>e�@ۛ��񤓲���c`8c5%=���q�x�5z1�d�������k)kg1W��wK�R5�2�r�o��.:�v1jQ�z�^��0`�r^��F�X���kU�x�r�ċ��r=r�B�>�<(�<#�2H���g+�NJ��L臼���J�g�ߋ�{}�ӷ�a#)��]����<IJ�qo�`_/[��G��o2��EL֏N���2(�Z�)�/�݀^r��n���	�®��{���-����w�s�F5˖�e�
61R�Xf)Aך�oV��;U��e)����W,ީ�-O�gr|ý�h]П�|`�YsFW���`��q�Ql�(#[��:e!q�i��ӡ�=S�F�/�3�ܳ�f^�5��N��}�$H�k��v&��W�*>8�@p8l�A�o�%��C���:��̐1Ů_e���ްr���(\��szwn>��Xu��Gh����7�<	�m���8wA���j�ْgo۪,�%Uh�	B6TD���G8Cpl�6�5	��Fl']�ɩ)M׈a�z
O�64(m�~�!]������d�HYw��"��V2/�n��[�:߅�
�6�s.� ���Wf��u��o7ְ9����AUTQ(�1AQ"�Ab�*�1b��Db�UV(���I Abŷ^���~����ս�`��_J�<m����EnҾ��%�;*���Pij�Zm�B����Cѫ%�Wc.��lur�Z��K�+{��\�����%��GU�w���3J���直�b���������02rI^�]�A$լ�z���yeJ�vH9�w�<&��8�$}­�n��������9y�mb5/�9���Z����
�b9ifڅ[��=f-^f�;����7�*�}�n9��WҬ���e��sd؞�o>�{�Y䤿+�ޏ�5�廒#O.���#C����R"
�FTh�j��DL�M%���,x�y�;X��3 ��_��Oj��J�i��B$�ꕤ��1~�=����-����2c|C�;h�3�^J3�RNQ|��wӆ;�t����{`@ ��xuյ����{y����5,�YX�����=��<P���獑�S�%���֊����7�v���B�u����w����1}l��h�i1�u����
�И������y��Q��uj�PJ37R������|�z(�'��_�">R����h',�u@*�P���g�Բ��|{knQ�H����a֯9�!�,�y�oϫ�mz7��Y�v�}��n+0�j�t&U��f`-*����5f�`�o�����,֟��`�+���'0]�[�	2*C�}���ϸ5�8�������{vg��VG�����>�d��I�l���.�{S�b����;�����ۻV�0��z]��Q��I��ۋU����k�g�h.j�%���\��g��x�ҽ����!߰Qa���pQ&�[��e.��wVl%v���W���l��"̽%��Ý��3w�ۃ��1zxf���[<�%HPJg����>�Eag+/oѣ\m�Z(�*@}5Vk� �JU6G�k/3�o��%n��m����IK�ʵ�������()�����To���?;Y�p���u ܡn\!�N�3g$�­hZvzRI��w�UKG)>���(u��>���������j[
?����V�</��[9���g+mIQ۽�9U��os�t�v�L��\�El�efU���<Vb��&z��h��n���o��f������H��V=�K*���r��}E%`G�[֙�]��:� T�ռ�Y�nnmE�*S��9Af��V���*�E�jZ� ��)����n���s&A�2f��(*�7�lմ�B��CV�.Rr	�VdTީ&Wo��Ik�j<�����<ȿ�UWb"��T�U�U�(�UF#��b���E"����"�("�
*���(*�"�`�� �[�)_���^v�-���K�0a�}_::_�N�d�'2|����O��0�:������F��P�r�ߔ�~Z�]k���) �X۫d#Ⳅ\N\1X9�f���z�Q���_�,����?U�@x�
��;�����p2��������)�eP��#b]�����X%W
"�gx���ea��p�tu�ݶk����:+������1r-�9rNF�ʺ�٩�9ݣl!g��VZ�9گ�Kƛ����aw�=��3�,|����S�z�z�4"�C,�%�J��味�ƺ6Ԗb�8��M�L�'�\6tY����ݦ�vq��3��q��s�XHQ
%�����C�W�ѵw7��U��{q��ݐ;��m}+G�4J���`1G&����Ц����켵V��
��,�Hůmn^�;jj���x����Y�'ˋ��ȃì@�q��t�:RǕ*.�^�`����94�xRF�ϊ��Z7��49�+A����w��"�n�-�g�״˓j��E�y�N�����������<��Z7��b�+����`���a�0��9W���.vv_o�U�4��/r^<y4/\��ǞH%U��ւ�4�T����u�Z�R�\;,\��������6�5,�=�(�o2�n�Y�PA̗�-Ⱥsnt|ӈ����c�{E���������x֜U�dӵ-�	WX�w����)������,��ʔ�uz޻~��lح�ѷ3]
,cw��v�Kלc!sI�p�rL��]�]��WK��Z5�t�v�8����DK��ٷD���BֈO3��eX���}a�v���pj��uU����	�sI5��rh�iyL�!�6</�#8�][��/�X���dU�GL��r�F�E�%I6�05��i���{�㚌�Pr�fWO����x�=�f*�f�+7'.���xvPZiL��' �t�I���/�&1^���Z�
�0�-�m�fZ����GVS;u�U�HF�\�F�[�^R+N��T�S�N�=�ʩ]kv������T9x ��6`��oΣa�*\�]Z:�$r8.�|�2��z��)G�הHrҖ)�'B.�E��:7�;׆�c��]W�+Y��N�:KmbiQ`m�MF�m��\��qà��L�N3]�i�|]@�k�-T�Z���"(� �*#TX�UV*Ŋ"EP@Qb�"E#u��Ҫ��K�݁p\Z����՚�x�(��Ui!8�U�g&Gx�C��<����x�w�9��[7Z�s��O�l$1���h�8�{aL,�f�6�{1U֕�=�^��]���d1̸����ph�āw��L�d�޶�����0���+rYḲ̌k�(sӼ�i�v�m����/��L��u;p�JL<�z���6�(�ۆ��u�*u��c'�QV2�n#���0D<;a�AF�9���l�#���w8�����a(� Qyq6�in Yf����h�c���,���N��Q0�ٽلSn�XJA�i�j�N�S(a�J�Ud�۔�i,��z��4�r��DW8�+Į
�Ԭ�W��4�1%�RiI��Uz����E�5��w�<�Q�
I���7u���lX�
�Y 9 q�2��EK��q�^sai)�ro}�I���9ʙm��%���"��PZt���S���:JL �i���{���'���Ic)��Za:B�]�&�;�`��N�7�,�2DH𚼡ՙx�,v.멅��h����&Uڭ�k!��!K�Y�Q�,q 9r�>����Gc�6	��
t�ݚ�S
i�3W�:�n�q6Ŗ�$Ů��IǷ	�HG,gK,�ŖE���,;�b@���wF��k6e�L%6�"�3V��lϘ��!�DX#�����.��'2��C����yo#��rGt.��]��x��۶q��a-���gl�(����JL%竅UKE�o|�m��t�d��i�UԌ 99ݷ�R���-D)��e�����e3)9�z�}�2�r�Aa����0�t[�7�,4�&o��&I2��U�Q)�����\z�p�	y>����i}뫿��/�4t�0�P���-���HZg�KE!uF^4��:�1x�ӍQ[��P�s�K��2嘑���D�p�#3�7�v��gy���\�,ȊB���y��5���v�&QWE�w�,�2�D9i�玖p�;In-R����yݢ/i:��Z.���3���n���ײ�{B�d0�9��t��S����e�����%�v�f�T��e2�Z�=�ݽ���:�B�S2�Mw�oT��!�˩����Lb�Rctc4m�-�o-J8D�a$"�N�=��a��Z��m�fw�f�6��"�����F��k9��O�B�@i xbI�7?�����	��Ag���i�S3X�Ƽ^���!��ˁ�"�ZH��w��c�����IY�0a�I�^h�ki�T��`0�Y�6�:Lu���2[)�]N��U۴��M��
iӺ��z�uS)���"��笙�N��&�!Ĕ�4��%��z+����8�[̛f.��a;p��Z�faC�t���t�E�cz�d7˹�v�k����ZS2�5Q�����v�m-�坳g�OL��1�����}��&Y��f�F3G.�3�e�5u4Zi��,�ᨀ圁���q�ZM�_l&�kD3���upm_s:`�ʕ/�$�������}0��d�˧��B��s��F5�2�j�M橧,��1�B��
���K�"��]�!���b�r�����QF��2���58��)St%�q�6�#����d��X�%o�Qg�x֘	�l{�^����pѨ��oAsW_U·e��`�,@H�\��;�y������ƭ>��Wq#Gh����S�qrb"�Db|:c[�U�3�HH1�B�t#�/o5�{�{锂Ť�1TUE))E���4�X,UDPi�QUE��S*� �*�b0b��
�Q
Ad�.I�9r܉��Z�'����+�-�H]�y�hЇI�M2���֦���#���p-�U�À8���|-%�Y��Cp�[�x���o*f��;Km�kY2��(AgWE�Z���i�q$"����q�jQ<����M$�n�9�Ke3,�-7�N�}^.�$�6;�vs��2�O��a�9�'%��x�
F;>8�|-0���P���ތ��L�(��ۍ�v6�goI�5�[�`��zBݴ�\��,*�:��Us�`K20�;�,�jKH/i����4�X`�pݫ�M�qDAj!����4�*�}bҨ����N��+����!��q-9�2�Hc����ު�fs�,C��;fY��(�2�{�W���P;KKN��s'i�7ʝ�!X��.�hS&^���ɼo�a)6�4�3�uy��vӴ��RuU.�=�e��J��m4���:ΐ�Agl�e��=��5���ƒ��{J�n$��f���ԷlOt,	g,�9��<^�VA޽����g�:�1�o˼}v���,���ף�:I��/=��>��������V-�}ƺ���Q<Xisp��;�=ڔʮ��%N,�����0䈵Vv�[ILۡ��j�ޙY2��oQ�9b��8�<��Zg�(��/7�:�Q"��}W�t��U�r���8��b�֔�D� h�Ex-y�G�/w���������U�aB�x٩\��Ҟ����"y����x��:B�D�}1���۞X�Q�5_���c���~L�]�_��dJ��V��&�y&�CQ����d������I���a�Nɢ�ǆ���%�~�i��Wgu�>�h�9y��Zc�n���D�[���9�S��r�eu��60"d�bl]��3��>μ�W��H�׭�{�'�Ƚ�X��\�]�4ߦ5\|��;�B�'{w݆��^��?N�0��7��\�75��xZ�F�D@��t;�S/�����L�]���7.NY^'�>������^~��q�G�zo�|a���>���	p�Ǘ;���a�~�y�w�(�>�7���f������Q�ǩ�{��]��׳M�|�>v��uwGј��.�7��>,��~y�`Ӹ����>6�q����Sq�J�[�\^�ޕRx��\�*��.�H=^�8�[Bj�� C1k�=Z��l�/���!�hr���)U�@iwc�B�9�8�j�鳩ì�����jZ��Y;f5آ4��f���\��(��ﺭE]� %�u���W��(Ity�|%n	�Ȟ'\�w�5�of+���e��]P+ WF�L\��;�T�����C���;��3�՘�b�f��pA�qS�8l"���Dr�0u��V""���TP�
*"*�A@`�Tb#I@�"
�X��H����EZhDF�ETF*�E�X����Qe4"����
�Ū��EU"SBȃ��$� ��������Y�����
�zv��D�8׷tV;��ufzQ1V��
��x�$�����wV�0��l��J/��zn����r@�e׹��c{���!��](�'+� �uF*9NrrIV�f��s�c�-Z�����jl%:J/ͩ簲O��T�G?vPꝞ|䇝�W�X!䪯�c�r��Gb�0�e3���!���}i|:M�L�nWp�ߍ�ɞ]Z5i��.�+5��q:x���Y�����m幇|��{� Ѹ۩�vھ{��[���NR
�͏���YL����aE�xDf�ӊ`J9#	z�+�Dby(e��fv1�w���X`����U/e]'r�
C��L{���<"�^���Č=�ޭR�A�}�{.�\H��"��ȷ\-o0�1׋6�]���GMԕ׼}1e@%��Jq�~�&��d�ϕ�n�G��h�� �g�|3ls��S�L����j�n�A�;s�:cu��M��}�z��u�]�n<i5cy.��خ���nۥ�[J��F��r惲o�Ϝ���!׻[dhd�!T�w��p�*�g��?/yG���q�1���"i͓RnHϬfpB��It��U����Cat0��^;v��%�haṴ�ɻ�9�69�<"�����%Z���/�݆���+���٢��Z׬BOS�}�v��'Fa�V}�ǰ��Yt�o�*#�KM�b�&8��3�0�i�³~eŁ�7�B�����\]՜?{�mZ*�'���KR�Pf�ZI��=�-Ik�O�>P�5��c�Ô�~����W��*�vZ�jC~\��ő|��_]�!��S��eǂ�{��yZڃ�y��.Z��ۚ2e���bDd-��5�YN9'�ŭ>�{�/���ރ]�D��2)ڷ�r���#�YG�r/��ys`��F�vҕcݙ�\�j��\}��q�=�~��n��Jք#�v󚭻q��r�Ӱ�u[�]���и5]���ku�]��q;7��d�2�e�4~�!|Kb��7���T�fa�Hb��B�۾����r҆;�Q��]�x{Ei�'A���G ћb�"��K��q�c"7%�gYW�FK�y/8��kD0��4$��6�,����؍]
����4��]��s��t+�J�ܧBS1T�{rdB�ZE-pY��S��H^��{�k}o}[�^z�%X*���TUB�b�DU�
�1Tj���(
#�e �D@T`1�ʩPAb���2)����VF��wUW	􊯈~rvt �ܲ��Pԅ��2�����~<A.��ĻK�b�ѹ�]��Q�7]����h@��i�q��&���]G1�)�m:\�yzd�mcY�1�#xSRF�zG�Hd+y�y�ejZL��q�e<��'B�v���p��̮>N�c�&�t	?	̉4�/Qѽ�e����GH�!C4*��]��N��.1���#����+��AA��gn�o+Zm�^��ƥ�)W�������vr�ufh�1l���^�a�#B��r�*�V��k�H��}����'?V��^r�6��ߦMQ#~ƍ�mKTg��T��U졆ܸ���֩Ň'y���Hosލ,g��t}FS	x*��`/˛MJ�(��OvM�_�oRˇN>D�^�2�A��`����T^��;PNT�y�Mt˞�'*��'u�Ki1G�<4�]r��20@���X�Y����5�+j97�ߝ�2��k� dD��a���>���"ޫ��f��H#���VP����S^�M�	P�ʿVz �,f��9z��Y�佫i-��?9���R�7��xt���kMY����
,����+��qه�V@��%�'����q�Da���ۭ}��ޟ^r����L�늼�r�\���H.wBI�g(�}��{6�������{@���j[MrR���$�Ù�63��xd�~�&�slFĿUn8��=���\
��ڭ)�}Υ��	W�3ȓwp"܋�&�G��Dv���+����0��x�Q{zt�Sώ��}#�k��G��|���W�w@�W˕��Q4>�y+�N��L�[�<��t>��v[�wR7$�ꡆ�ғ�&z7�øN��2���F2�-Fܑq�Gik>�).��E��7�j�,1�	j*���Ch1�DZ-<A�|n���)�UE[�P� B�>�$���rT�@x�t�[���*S�E��f1��50�Ͷou	 -���l���$�`*J�����H�A|������3������P_<v�Y�g>���a\���9�oX��Y��.�����ff��I ?�N���/w�~!
@���2t@ ��{aRY�������A����>�,O�����=����o��$
=�Y$����_���|T%�� X��%�����Od����V� ����/R!�?Y>�W��v�`��d2��I�ϑD� A��c�^�;��`5	 ?]`.�*�u�Qegʶ�����l>�$��?��I <����z�|I�=G��)��\>�R,�K�_z~$:=�'�������`Q��Qo�O/x2�$ ��ʏ�yϜ<��R#��E.�c��S��(4I�{�_A�������>��ǟ��#__����g���{؃ϳ�E��<|	�C�?��Ԉ�D	 ����$��߄�����I�h*O]�����,�3
!=`}�I54yڨǰ.X����'�ܐ�1�5&M���M@�����4��u u��rkT}@�UC�ك8�C�X�̒@vX|}�����l$���D��#�>^�=�?C��C���y�Ώ\?��\�B}?G�x�G���_����������C�}��/����C�P� C�|�z}2~d'��a��Ht�q����_П�ק����N�@K�N��HfH؟d�Q�����]{�H\��~�_�������F���A�g���I !�=E�{����A�*�k#'�r���y����"�}ٯW��bIA�� ��d�O���,�~p��Ͽ�o���?� !��|	�0�c�A���4��*N	3���d��������� �.�p�!��V