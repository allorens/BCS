BZh91AY&SY��3�ܙ_�`qc���"� ����b            �                                      �  ��y�뷷=�       @  � � �@                   oҢ�RT*����(��EE�*��������UQ*��� B��U*R((DUQU%�*P�  �D$�H Q$��ܸEݸ	\�3A7w*�Wt*i�P���Q����vꈖ�B��Y�T��Q��   �Ϥ�@ ���Ň�]�z�y5��)ް<{
9 ��=@<m�B��u �N�9��`<�\� �   	/}�U/�ʅ(J
�E	U�$��|t3� ��`=���� �����O�v8� ����!�'�}� {���� z2>�� {��   �U@
�>@zG0� 7<�D� CϏ�:�5� ;�w� 1{�TS�� vï@z��G ;��@  Z��T�	�%@�����>� ��� {�cG{ A� 1��v�� ݇/CA�@���� w���g���P�   �>z��� ��{� <L� $g�(�Ǝ@�������� ����{�@   5���� r�T*���*���R�� .È�D@wX�7`��`�� �h4@1��{��nH]8!�F�8    {�*( |�|���w�+�hvr �2l��{zP�ΨU�Jn� �0���"9i!    _>�� ��*��Q*)U/f}������;�U� ɇU]� $� ҃@�Gv �wH��4jB�A�   y�JP ���G֊�*V���@�#v p�2�#��B��A��   ��h`(T  �"`R�&�i�  M ��RT�       �Ѫ�E�m ��`�	�M��&�S@� �� ��(�6���      �j3J��L)�"l�!��4��b}�w�~5���"��'��#��L�k������(�a?`����A>�QW���O�hE U��O��{�_ݣ���"�*���I$��P^�8S�������_��xF����cR��LK`[ؖ���-�m� F%�m�lK`[�6Ķ\�c�6Ķ�-�lKb[c6Ķ�m�l`��hcؖĶ�-�lKc�6ĦHK`[LK`[�6Ķ�Ķ%�-�lKb[�6�c���-�lK`[ؖ1-�lKb[�Ķ%�-���m�lb[ؖ��%��-�lK`[�Ķ%�-�m4Ķ&�Ķ�m�li���4��%�-�l`[٦�)�lKb[ؖĶ6�[LKb[�6��%�-�����-�l`����-�Ld��l`[ؖ��%��F�m�lKb[����0m�lK`[�6��%�-���m�l`[ؖĶ%��-�l`�ؖĶ%�-�i-�lb�ض��-�1�%�-�l`[ؚe�i�lK`�؅�cb6Ķ%��%�-�la[ؖĶ%�-�lb[�Sb[L`[4��Ķ�-��[����%�-��-�lKm�1-�l`[�Ķ�-�alb[�6���-�lKe1�%�4Ķ�-�lb[�ĶF6���-�l`[���%��-�Lm�l`[����-��lT#K`)lP�"�K`��*�!K`�lm���ER؊\�U-���B1ؠ�K`lTm��l.B
��Rأ \�E-����6�R؈�Kb�lT$�R� � bl m���T�(�![������(��R؊[K��%���[ `rT��$�Qm����
6�R� �rT� 6�Rث������b�l m��AF؊[t�[b)LU-��A�
��؈� [b���A�
6�؊[K`�l@m���GL�4�؊[K`�l-���@ت[Kb���D��[����D�
�!K`)lD��*��ؠ�`�l nB"6�� �m�F؀鈭�Q�6� ���blm�܄#b	l@m�-�A�"��F؈�-��`#lTm��@-���*��-���P4�Fآ[Kb�l@m��T�l@m�.��KblnB 6�F� �0R� �`lU-���Eؠ�[b�����A�(�[`�lTm����؈�b#lm��@V� �Kb$`lm���T�������
6�!m��Q�"6�F�(� b#lm�1�6�� �lm���-��lb��#ؖ���-�lKclc[ؖ���-�lcl�Ilb[ؖĶ�-�l*B[�`[����-�lar$K`[��ؖ��%�-�lKa�Ħ�-�lm�lKb[ؖ����m�lb[ؖ�����ؚb[ؖ���m�1��t���-�lKd`[e�-��%�-�lK`[��b�LKb[ؖ��%�-�`[�Ķ%�-�lKb[4Ķ0-�lb[�6���`i�lK`[�����bSؖ��%�-�lb[c���-�lK`[ؖ�Ķ%�-�lb[ؖĶm���-�la���?3Z��!b �����e��|��5��z� ��HF5c�x1E�ia�z�GmY�����V��u.��ǒe�OmP!9k4�� �sm��9���^U�yoo"���F�ඍ㗦��M�g,��u����.Bt�%
�TiB��ʬ,J\�Y�y�@�ӈ`6@�W�X��cu�����d�ѱ�h+&��S6�R*(;u�Dl`��5bm��d�t�L2��Acq^f̤�é!H� �2��"K6�'tn�B�2�Ġl3��� ��)����[wQ�W�EY��t��+O#�"�\��J!d+.=)���{�lG/�i��3��&�,�Y��1�R%Z�ҕ���z2�֤����E��mE�`�d���tt[��U�䫳�-)
J�WOZl<��V�[�@u+t��/R�4J�"6�J�Q݇!+ʰj[���2����vYۙa2�Hqb���,=ukw6�TB�bY�L�vj�EZ��K�aV��fnz��X���@��/M��IR�'"WY�nTvS��֭�r̈́���l=@�fS�p�Q$(jU)�mY7��yZ��)�38Bh(����f]�svTZ(�3RVӮ�Ƒ����-�JV�յ&�n��jii���j�+d�j-���[�M[�F�R�'w�<nd0n��X�]+�D�wV�sV,��*H,�c�6�n���ʽڸop]'�W��� �+�H���i�S$\��-/1I��h�12}p-B�-CT�8(�9N�^Htm+��=sn-�m�T&�i .����]өkwb4[���y��N���0Ew4�ͅd7.M�5�e-r�8�*�VY��A�v�f)�
��ՙ��vϷo黼��oj&6�kP$�o[��&�5�S�ܡ���]�:ۈ�KaN<�A]��uae ѐсGD��:�,ʋ�d�oU��i��ɦŵ�CjV-:��i�A��^Ǚ.a�˓�񂱢�e]Z�B��r׋�t�t|����B�Q%J�3=����ZÕ����]�9�/�O2�X�+L���6�l��Xջ�"�f�u T8�T����f)�R����5G!��n&��zVn�d'X�/.��̢�^%�N�,�R�)=5�kl�dOsE M�r�擳*k���YJ��ѱ��ML9�b.�=��z���ea[d᥷n�kkcʼ�U++&"t*��K����V"Ʈ�؛���m�ڕ-)t�.�5g7E����q��� 7`9�0Lٷ.�۱=�q[u(nܲsQoEZ�	j��Fn�u�^&�W�L��:��s+/0�Q��-�Uɘ\6����İ�"��B�2f"�[�eG�̋�,�Z����t�QZ�<�DB���D䧏Me��9��~�yHhXEc*��D�F㧵zm�TKխ��K�2Q��v��2�6�U5�ب�n`�b�aghk�.j�7go�Uy�G���iB
���(T#2	x1*��Z�ʹV���m�.�&�h�R��6��7 Uֈ��&d`EX$�Ȱ�m����Ve�����R�5� ɺ�K#W�W���-7f�O!
�v���-f0<o[pTG]�[zo`1(��5�]�I*a��>�"���G�z�L4�maG07l�r�;��ˌ�]�z5�,�h���M����;��H�G%aʱ0bw"�+#�5���B�2M��ܛAenmͧf�@��V����-赯r��i&�Ѕ�/V�fh[� 1 aR���*lz�u5����[z��M:p�Y,�z�Q�jaݖX�U�é�z�[��a4��B
�<�c��V�i�;��f�x-�5���$�е�r����Q
{7f�,Q�]YG�r�T/T)�����р��Ӵ�VT��:y��͠��$�ĝ� �k*�ˡg2
���\Y풰r�����8U�mQ����֬[i��׍�u��i���l&@�y\��u�u��w��X,Q�+r��۲.�aQC ���*�ckl(VX���m��/-7��
ݕ�jTh�hR�
�̷F�:u5-��ڵ�1E�4��'F�lF��@p�ɲ]h!��^{�Ğ�w���K7��E�Cj+���˲���N���l/=U��2����$`P(������d���73M�Q;�k�����N�;G��l���q%$qefZ�[�HY+p�.]�z�N^��ʸ�7Z67��M�B��wk0�&�*V�n�7�]�.���LHU&LB���Q�~��z�� �{��rcU���
:(V��ɲ�R�%+��ݼ�M�DH"c��Y�&��P=��6�6S��$㷕�
˫����&Y�.� �o�M����eJ2��i�֫v�5ӹG������1b؎ʸB������
k.ڣ�V����J#N- ��A3�u�,n��7Z�wbMU,�u�0l�AB]�E�ĨQy�GoAڙ[�
:7\ʖVT�-�5Lѷ�"RJ�Y���r��3L����w�)���d��Bm�)�6A6�/oC!�D�e[��t��Z!�gl���K3.[��ە��SJ��[AKX�ڮ]n�i,Z%��3�(�X�z�b��ݭ�T���yI����=�%���Pn�˂�*ѫѢФ�����i��Ɩ셋z2ƣ�v�oN\������N��^�������;��X.8k��(���ra�yn��_�1��Z��~X�� �(B��32�a������V�7u�N�L�Iݶ�捊Z�v6�A�/n�fe���4��
a�|��)��-NEɻg�Z���(ca-���jq�sd�Έ� [y{(<���D�8����fh���e��]�8��ǖ�q���5�d6&�9��ܭ�,�D6�d~�B��/v��/T$б7ul9~�4��CUwx��u�94�@��KP�HFʹqOl-ٛs,���eP���+p^���U���ooT�!�FFS�݉��^;�
S%�ʻtJ���=�&�&U��4G��^��6��Y�ǎ7[��4�(n�T�iee�����]�"]���J%��2C6R7e�FD,�b��_�Ӆ��hЌ�^j�Ţ��ۚ^̬�G7$4�k(Z��`B��Yxk0�ۺ�r]�[�Gv�T�����Mc"VFf9��@D��={V��݅hDͣ2����* ���Պ�ܣ�,c*	(f��v����X��]��6�A��� ��hsjf�9G��A�l�t�@ۺ�Գ`ڄ��FyM�Vv��ZݣN���f��[�PY�����n�G�Բ��2�Hj�&i�&�P�-7[G#̦�m��ySF�9I.�ʼ��ƻ�ȭ��7NT���^���v���c#.�ËU�rl�)��~ɻv*B/30	JB�
�Pғ9m�A�ͽ���bٷn�e���͆�9
bϡ#��@�n���N����V[�ҵ��x��D��н���ƃ˼yK,�ɋP��F���7�r�F»��R�$ѷAL�����B�ɰSպ^�B��C*"�Z�Kճwv�ݻuN�G�Q{�TÙ�0i�^"Ә�9����PٳZ.�-�)e�5�ܲ��Vuᷢ{(?b�w��ۉ�F.�Ӻt& �3keFN]C�b-B��Trԭ!$��Me<�r�e�M��݆Z��%,P�KK5B��������W����ܵ�-�/\����[r���C�eY8��˘���WotIZ"��;��fK�3"Í;J<�m]���e`��.���S-b�M7B2���T�O��2�U���t�+T	
ܩfk�N��^��%{[���1^�̚�հ7��j�PjLщnݵP�;�[0Y�(�X+kR�������L�H�iǈ�y�Z7Z/^̂�;rjȄJ��Y��H��zs�:B���JU���K�hjƷW��H⣖^�nì�˕���aۤp��ˢ���M�kL�3M��䫙/NQ{`R�w��X��B��c�̬d����7�����ʺ
���S[�KM�`
��u�/mJ��&�P�f�c�LԴ(k��L2���zd�s+=�l7z�Bc���im˸[�諢��x��%�ZQ${���GP�[�v�^&�5!���q!e�{pS�xmU��x�[���A�h�Y��{a����ЭW�5$k"��u0�wһ�[����7{1�wx��Ԛ$%�n�"�c��{���,�o,Gko�f�3m<iU�nXY�vX�ux�^EÁ�ͳ�A�l�k�[�����2փ�J�ᙃh-w�9�J��A��;w�hؗRb2�us^5�fʺ6�!�j-�����v���dwG`@�3/i�R�(�.��Ke���z-;�*�{���Y�Ǳ�h:�H�ٳ�^�Y�5$v��͊��0&=z[�b�Z5���r���j�G-��b��ݼ�-�jx:ejط(��z��m�{���2�3M]n��#q){Kl�1 Cn�m�sF�� �Z���VA�%NA�dܺF��Wt���@����Ԙ��2ݬ��T0^����ݜ՗�淊���� ㆮ+R��u�<ձ]�mё$sh5zrLV,c�2d�&�q�����[��"o7+���c8�n�f] �%�r#��ݹ���B��cN�ͬCq;Bڥ$�&J��O�e���c,5�q+�Cvi{��em���]Kp��dyD�r��� WL^n��[< U��֛�ۣR�jB�5a�[�1,3ɥ���̩k2l�\L�@�I�tָ�wE����*/�!�����pѠ�/v��X����[{-K��8�������2���S��������hA ��S�]��9�I��]����Mz�y	Q�۫�OYk6�o��S0�)`x����D���'��n�R����Z�z����2���iK1;Vp��LZʅ��`��Fa�e\tx͆�K��H�8���a��A_��/)�I	��h�<�v��, �H���{A٫@���T�mc�XHJHl�b�ƃB�;W��ؤ֕і�;�yu-���?,{�a�;�ojlKsnLݼ�3t=����;c#N�_����ܙdڗ�Ջfkڼpc`f�D�Y��i�Ȳ:8�Cpa���q��	-��`[W��` ��c;X�&��n�RK��/+�I����q=�+snQ�t`���"i��/vU�ܭ/"+.�ف���Cr`��5N=[���S�j%���e7i*�;F��V<�h��Bj+�hJ��4�4e���R�n��z�2)P
�ژ)�Ӄ]�!�1ݩP̶c��HKiVee+T�x�Sho��w2e�u0Z5n�[��J�g��B)�ƀҶ�ݦ�"�0�ҭ�l
[�E�����̚�ieHr�F��׷kcr�CZX�,f����#nRy���q���J���B^x`��0=�E�L�q�K;�L<���q�C*��#p
�{!�%�a����0���g3[WY�320�ELx7K�������ن
�m�Lm��8�.���؆m��-k���b Zj�o�,kmh�*(���m^Q뺇-�/eaݱlm^��"n�w���������Z��˓Nh&��f�F��
̖�x��ØƱ��HI6x�.Ͷe����H�3S]e$w(�U�Ç6�
B^Q�s+,�z��^պ�f����4�˼aY`+����Xe�&�E�2�87t�2�������N�VA��gf�r�Q�i՚Ř�ڍS7L1�]㔰��6��e]n	yR��C[`$��̗)�ku�pA�vj��$�����B)?;F�+(֊e�WwWHe6��oX�J��SҴZ�����&�d�z$OqnHl�֞AW"G}�U��vd�w�j�M�[��]��(��[�b�;r��ʵ,��� �Vp+W�[���qU���+inLw�%5���z6Ƭa=(�vZ�ٙ�kNf�$K��2�d9���F��3k7���wtۖK/T����Lژ���>�w�ywh����u�D礒K'I�	�ᅊ��7�����E 2巩���;\���D�<N��8�K&�$�n��$�T�1i6I.���I����Pd�6L��I��9ɼ���М:��L�d��%�쭬�>ga�3L��|I�3��	$ْ�k�dOkށ|�KI�]-E��4~��N���ˠ	(�-���a�l���x�aũ�Q0�c1akr#�(ҶM��	�(gH��Ng4�M��Ʌ�l�l���'�u�^RxG6�FQ��CIu�3	���'�D�0���N��a¶�-+b�0��N��.or�m�7X�e�鎀F�I&�Ӵ.�D��R�g<M���$�N�Z%��i��^JFc��.+zp�;��tݾ创;�o�il�'Id�YJ�umv�u���"��L$��77wa�[��!��"(̾x�q�[x5�؄���q3��-�t��\2���͓|Oo̲�ĒB2�7Ċ���bBMk���C�w�%�i9��8�)H"w7-�b�,�5��{Qβm�1բp��8�7�o�2H����Y8�7N�fVs%^d�c%q�9Z�R������h��P�ow"�y80�I6^[�IH�$Pe&+&��,�諗%bÊ�n��^��8��Tj�8��cs,�I(��ZU�
�/.�V(GD��nLډ�r��s%�h�M����E�N��C�1�p��������+�eř�ڲأ�ɠ+4�mM	���tm#{��9�|�$�j�_}�#��f�;q2x�A�^�fJ��7N����E���1����G~����2��m%��Y�s	D���;��i|V���չd���p�d��HN���I��Z��bK�d�(�v^,%��]n��-����P���8N��ՂM(�̩�쩘B6ɳ��W@#��&(��%(a�3v��$P�2�EEf���vr8�$�l��p��+l�-��Cr��CZm6]k6�:N���p�e�j�%������M�ъb�9ݺaJdL)$�V�%Ib3�{�7�}7�Z�@������ok�(!�@��ddEj��UEX�V�ڢ��Ѷ�Z�-���V+h��E���ض��ѭ�E���b����b6�TkZ+[F�m�c[TV֍E��E�V��kETU��Z�,U�F�ѭ�V���F���ŭ�m�mkh����ձ[V����6�Z�lU��ŵcZ�E�-��j�ձ��F6լV��ֱ�[[lmV6ڍ��ѫh���j��E��mQXŭ�U[�[m�ֱ��Z5���6��_k_�o��H��ϒ�p��y���/ʐԞ�Ӿ���������ȓ�,�����4JRg(��^!N��� y
�I @MfdӰ�Q	!�9fr��Zj>K������7T�<�爗�A�P�0J���<X2�آ<FC�j���+C �=�Gb;���f&Vj��Ō�Ҫ�3��5�X���xΞ�7Y%�/�g��At��PPP�,D�� R@�4�����<���$u��!�P.~S��&S�FRm��#�d�Qci��Me����R���UU��<6*�U�ߐ��#�7$��Q�}�^��y秞ON�����~�'��!;�N��\J#����^�>��K����.�O��)�{ʌ�|��W:�C (��w��Fe8�� �f�F��%/wy�I?F�$<���7����ִT����dG~wF�;����xJ� ~�����`�(����!>��b�����@�*(#���������~����
�����j�M���m���n6	7��w�;G*[YE����!W����)���"���R]ۻ=D����`������#�Gv�ΑV�<!�Y舭�ݼ��Lq�1�Ɏ���t�hi��%:�!ܪ|Bk�c����z�s5���ʘ�o.�����V�`/��ɺ�z�V���G-f���`�]�\���w�����BEh�_�вt��Ƨ=W�Z���*��Gٷ�8�j�2dQ됞 �I�7����#1sjM�e�"�]�哆�kM:�
9�﹍��!�;lvw~�h��g {$;v�]w��a�a�c :P��� ��g^��!K&��}���޵VJ�oJM��	��K&�NO(�����^���3\����u#�ڲv^�b�Aб����+3j�Qm�s���\�������N��lkP����k�r�V��J�t�g2� 
X���WvU�[��vҭ�̯
�f+��<9��Bms�Cj���(J�b����\G��0��w��9>�x:e����>�+D��R�����eW�k�aE㡼Y���*�vQB\C{㤮�a�;ֶ�)U������b5
�W�a����Ѷ%+ǌt��y�3|�rn\ߚ�\�Fݻ||qۧq�}q�8�8�<pq�q�q�q�q�v�8�8ێ8㏎8�N8�8�q�q��____\q�8�q�q�n8ӎ8�8��:q�q�q�q�8�8�q�q�q��q�q�ocN8�8��:q��{�������
a�%w<IEu�/S���������ڻU癥^�zj�n<v�T�V+�N�ɜߠ���zļ�(m�6E�諂�Ʌ�R۝�+s�$Ƶ�Gq�ڋ��֌�;z����3�J����]�a�EӤ�X��mMG��@�ԏ!�{�T ����"���-K�٣~���%��c)�r��L>r��u����S�(�z�v�]u��\����e9���^���أ�M!�S˻[[�����>]�ֺ �Ƕ��k۰޼uu���� �J
,�SnF�k0	��a�8'����s�����ٵ�$BHI	Fy�6vd�˺W���V�.��6������'�XEo8Xܜ3�����n'r�.�4�y/Nα ��ɕ���*4�vF(�N��y��&�}�՝�ӛ]Ya�����aƅN�0n����t��cq�77P�/]m�٫GU��$E�9Z�+�\�u�sul���1�����N�����
������x��,u���Ԕ��d�P�]c�uJ�%��ɔb�`��wF�n׽zp�7y�m]ʩ�❕�c}v�f���գB�Pm�U*�����YCl���:҇�e�Y3��i���oNW%���|��}��l�5=x��O��^<q��m�qӎ8�>��8�8��q�q�q��q�}q�8�8ێ8㏎8�6�;v��O���8��q�q�q��q�qǎ1�q�}q�8�8ێ8㏎8�N8�8�q�q�qۃ�8�8�G����{���9�boWe;��/�&�h��K�oVgL�^w #�wEV�K���G5�\�]v,7�w��=x��5�$��h=���m�]S��C�w3�b���s����c����o;��Oic����IN�N��C8Ç�^�_�c{�LԵ��.�#w���.!�Dԇ�s؊�Ƴ(��x:���Rw��9�8G��Ⱦ��6��$�9ݮ��umջ�u�^IS���-n�f�������U⼊F����1�&�#����Z��p'�����N�)pؗ	�و:�l�<k�F�k|{�\E=�=�߫Fe�⬙(�\�j�^�ە�Q67Z�5Àm)�"�Ϯ��IWڕ����y��{�RU{��!����.MZ
��y{;%�
�γo]�[���^����ގ����s5:Z걻�Χλڰ(��H(J��,^͈꺆g#��	�Υ 5e`ۢ*���µ�ݳ}��{Zd�m�rI��X�OK��ݳ��3�B������)vF�Z/��	�����bwWO�����5�\� �z�	�d���Y�1�d&��㝝��f�f��u�wn�q�z�B�d#On��k�h޲�Ev�[-�%�|��A]����7-ogM�`8h���c�j�����=�<q���N8�8��8��q��q�|q��8�n8��q�8�8�8�q�q�n8ӎ8�8�nݻv�n8㏎8㎜q�q���8�8���q�qǎ1�q�}q�8�8ێ8㏎8�6�8��8ӎ8�8���q�|�g.Vk�=瓞��ܳ��U���%�)�F�yG0^���h�V*%�Uv��	�����H+��_l��	뽫&��ɓ.Â�]6(�!L.w�����Bm�݌>(h���X)=��UL���a+����\�c��������{Vm�8l9�[����6)n��^5r�Y����ɭV*p"��|����r��-�O����5yWB{�~/�v��+j>Q��4A[���.�ͨ��̩���z�r�wR��w��4
�pL�`�ÏR���Zu0c{��櫭h�5���5S*����q���:AyEپ���ͷ��vk�]�A=S �"O��{��$ǆNT�W�n�%H�M��Տ���u"Œ�u���nv�� �D��j�6މ�I��[qWZ�-o�;��WRզ��v.�xv�(�]�C��<1컨<o���;��,�X(�%��U��]Y�z�Sb7��8ۜI��b�þ�b����:���U+�]pӊ)\q��#z	w��#�j3}�]�È흪�Ӑ!������
���/��a�Qk}7��>�(<�7�a��0Ĭ5�J�
�]3�>uZ�eJ�b��8n�N����@�e�K��H%ݩӋ�~�)�#\"�`�7X!,yC��k�ݗ�*��t�UW5�%Con��G�����o|x������q�88�8�8��8�8㏮8�q�q�q��qӎ8�>�8��8�8�8�8�ݻv�۷n>�㎜q�q��q�q�q�q��i�q�v��8�8��q�q�\q�N8�8��8��q��q�|q�t�>\��h�\(uԉ֭'a�WL�h�}�;(�]���pb�
W[��:��X+�{�ɪ�&�s���L�`91q�sf���cjx�nP���\����ܙ����/�)�-he�[)S�hR���UUPr2VL�:ۢ�k4.��1�yנ����nؤ��&
�x��M�I�Q�,��ଦڢ*��klՊ�x?���NS��� �X�ޝ��B7�eT��p���֤�
0�
'1�+,�E�Ȧjt���T:J�Q��7}���\ӌ1/��Bxz�&�� Ԑ^�8��K$c!˺B�QsUE@7h�X(l��G����j�m��׊�KQ��Vt�.�fgc�z���P�[�V�b��c��ʻ��������i֎�]Iu9���8��%Ŏ�_g��S���-ζ�����V�oG��ތ�>��B�΁6/�VKƯ�
Ø
zXCʇHF��WY���^4�"�i�7�!o(�H!3(��a�+c�a��D���/,]X�p������+e�� �f�o/uf��j��Q��,��J�6��:�q��Y�t�V: =�qڊ{�t��kL��Ԣ4�}�9�7�0�%i9�u�Cշ�F��5/���n�w��[�ʖy�ֆ��;0Y��Ÿ�ގ�1*ƞ��B��yUHi*��]XhM�p̣�^Y�\���!^,�#TZ��E+WɌ��q�3��D���|*����i��7Jš�s3M����Q�C.�Ջ�l�#82.�R��6�T1���h����UY�4��r����l�o�ry�C��BҖ���c�M���Bj�d]��K5���;{Q��ԍf��5�����0<�bu-؅l�X>��i�A-�Z��B��{�<P_T�]�V�=�tv`Xޜ�)T
�����F�cՄn�Z��&@�>4,m�0�����9��3�+�s�7�y|�Xʹ2��&U�oM�O®���u�R9��2�q)�ƫ��T���苾�
�hT2���ڼ�\fWK�(�[�Q�t���3w�khslײmZ[�Zf�Z���v3r6���g��A~ۼ�Gh֌ZW��Y��1�Wi�t��U���47^.5x%m�9Wݻ�L�5��</����}D��n]D��];Qջ-�o;�.�o=��/m�6�m�t}��dWDr�:��n\�(mfY�F�*Y���{n��É۝|$,���d��w'*�ۛ�1��T�Ք����T��r��%e�������{�N(��'_w�f֠����i�L|sNu^C�N�]v-����vB�{��1�qËB�=�7v�%�L��<��{�3w���3s�'5����)��b�o��S|�(�I�fP�X�7]`����@粠9�Ź��n��Ƿ�:���zf�5d �պ���5m��T�P��Lԃw�+P�άur���9�҅�h��VGr
�3��3Wc��nk��S[���!7,�������Jv͍ׇ���2��˝�_>:]���Iu�3��k�UN����k7�u�|s;n�5�p^�w��R��=��u�D��̫|�����o,��ֽ3gL��p�����n��߆d���gx<	�C՝�y
o(<2P���ڛ�6��B����%�WH�W.�H�]��r��S�s�{��v�&�͹��Zv�r��vz�g:��ô�dܽ�i�K�"�� �[�	u�r�[�mV.ƪY��u�{���t3ʢw,���Qj"(�ȳBQ��3n1/@�����k��@���J���t��b��G��"9dq�u` ��ެ���v�4�a�a*i�`�7���s�{�L1xaG�;��m+#F�^�"�$t�]ڜ�-fWwJ'L�O����5W=���7q賽���-K`f����^^�f�gr�ם��n���N�B�E	!�1�W��\z���P�w�����X�-s��x�nC�U�ʸ%�.�#%��2�5�r��duϦ�囙������j��wR�j���nZ��fW<V3l�n=VV[yY����P��i���so�CZ7guL���-2���-e�v��+=i7=��=�������s��������e˧y\�!FH�ƇYX�wXζ�6����x�]����+�SQ���L�i�wH%��#�yy[�0vn�=�=;1hyX�Ekw%ZR��}����GiM���jvRy]�a��`T��wQ�Y�A�A�`�
V�n���m�A�s@K:;[�L��:�U�;X���}e*<4�'hڕuh�B��)�7*^<7o�w����:kkuqN�����J<]E;��)V��1m]V�(��ʹ�m�00�6�Ӏwe���R�u�
��G�+�(�\�{B!
�5�}2vG�B葠S�\��3��vK���v�BdWz���ۜ�9��n��Ku�7�#5��'&��.�̚��tq��n�wۖ��Eޓ{���c��옲�_`�w.�Wm��k���T�C�dc�}��zШ���ks��GP�Tn*�|{���ۮ7N�z:�]NU��uds�u��:6�
�Xa�΍)�̭�ܤ����Bzh��T��3oU�MC��r�5ًU����1�o5闹�B� k��G:#G��p��*�x�o��@̫DX��{3�d�;�N����&ZX0qJ�l����� �,x݈ۭO���u݁��0s�����j\ZMN��F��gdU˺Q���зB�h���n��Up�[�Ȭ����)��3z�X@a�:T��k,�R�n˼�wY���V0+4�����=� ۫W7�L:�c��-j�),,b{m�(���a�0� 錮���8�Qn�[F��>]�u�"�N���fJ��Z��y3ps
=�]����vH����kI�%n����x��]gT��Ž���軕�6������a�n{��q�pܩ��v�<��i`���X��S�e�����/����i��go-�ک�i�Ǭ�=]~u�9�pS����yɯMqU�ww�br�J���q��un���⡷��WժM��uْ�+W��mͳ�q�d��}gN��n��p)���t�-���y�`>���N��Z��k��z�՝�u��M�J<33D�P���	{�	n�[D�w��k5�P������v^���h�M�ھ׌�86Xzl�>���m�Kһ���w��q�f7��h;`��㝖�_E���t����[ء�&�eY�n����ǈ��"�ur��|w��{nY��jn퓻YP�)��Ք2�ˀ�W%BD/.��L9.\���Noc�];͜=f��1vMȩ8�}�0���YʖoXٶ4��io|l"��۶sh��p�]��{�u������ѕ�-�˥{��z�ݽ����l��4%t.��3V&=ܛ��٠r�ѡw�֮Vڳ�XuHoNwr�QW|�S�xm��v;k�]��˾��B�v�*�g�����N�Zx>9�o+�n��)���8�S�K�����[X�P����طQ��[HČ�\A��|:���=�A_n��b8�T�˽��a��w�5�v�X�1�_-�[+ouuvՊ����~���'Vwv�9��F�b���v��4ڞz{_e�cif^kb�&G�=|�_���|�kX�D��W���=4�9n:u�N:nl��h�_'q�2���'�z�J	��&�}���ë�����w��|���|r���
��۠=�XTt׬z�p��/v�˙ݭ\9����Q�u�+E@�lDc
j��l��Ṇ0�v]�=w������;G�E��Q0�/��Z�sHT�:}ܰ�f�"ܮO��N|0�6�g�.�R:p�4�V \OS�3de�ocW��h�;���$+��>.�3O��*d�nN�k��-*ޜ���&����e�6�z���g����v��wr�Dޮju_s�͒a��wOb�\�Ժ����i��p�U�)Tڽ��V.Y{j��u݊�u�}JB�=�fA���t/�����3/UtWJZ�DX�.�\'o���F�wwU{�E�9��P��]�c������|?O��_�������~���̿�Q���'��O�V�T,<q�Vh��:��\ك�?��e��.��.�f%�q����ٲ��)��I�f��#�h��f�VCV�0'���	q]����5�*�4����+���4!<3�{<x<�[5G��2�4O�o"kϛM������|�xs���,��I��;כ�	=����0�2]S�4������MG�O-�c��%sW�<]�.qV]m.�Ȫ镡��%آmH:�ԗF�ۛ��E��y;J5�9L���LTI���9f�;m�[��O*�-��mr�m�5d1V��2�nH�L`�(2�ES�f����+1Kk����W�К�hF�5��V�Me&�nb���Z��o��|ŭz�-���e.1,m �r����"�t�鍍5�7h��P٥[-!T�#���5��4���2��l�IkuT��e��m"��W��IC9qqSجc@[-T#Yn(-ID�G6kH�P��-t�48�� � R�f�6�E�$��j�mc^ K�fBf�q�1H����t�tsi��k.5�6������B5�	��h�K�ˬs]3�,Ő��QL����XME��ᦄm�q��:-	���3\�X�h9�s��5�KE^m�����kP�Yl�M���W%�|�7�Cy1��95#C�K����X�u���l�Xl1�¡���%�c�f����mA�{q�,x�u*�M��Rq�J6��ě+Q�iX�$p�Ze;K��e�7U֐��cH���/<��XS�L\�I�%A7M�0����e�1H���(��V�)�pff�k��[)3�s�ip�F�]Ib��8jM��]a�ąB�7�ئ�f	RT��뭮"Y�T��7b1�
W\#-�3�PlmtnҀ@H�� �=����cf�H�@-c��Y]. �e�Q��cf�0�6k�!�t![p]2��FM���k��k�,n��pG7��|k|�^�v�]�.u\�%+Y�l`�v�[P��%�u�V�E��A��)�@�ke����[���nP"�b�б	���Avic�I�V�Q�[�[ΰ���fpq�u"�����K�*B�-J��5m�a,��[0�tt���Yh��7 �� �h�sC�����WT��6���lp�&���M Y��Xunv��S�WYj�Yc��\$1fíu\X�4�"�2��%f7m5���˛�� ���A.i`����hM��kc���	+�+��"��R�"��ΚT[Kn[��43��U�V7���V��.%��
�CL+m������:�A�D�Һc�D���h0K��VU`�����]3I ab=L�Ap���%���,�%]��e�@˘��# �W�֖%�l�rG78�����0�#ImT���7P"E ��:�X��f��
�ٗ�,#l����kd����apJ�9��u���0`.���3C5�[�a�k5.�����Wd�fv�!��` R��vc�JK�[6�8"e�Nl -W7���	l4Aֶ��`�ɂ��@����v��+qT�/M���j�#TL�-r�v�mic\�Xv���ٱ��ilb+3	��%\Ka*���j��i����^	F�L�[5�j&�h��K�41���eҲ���h�ikFɇ7jM�ʌF�R�+q	ss���F�q�ck@�Ii�J"��ٖ].�����R�ĭh�ej�*�b�-�X%s�3�Ko8�;P����� �n��h�@k���P�t�JY�wl����0�.d��c�R���,(�\VX��,.,Sh�.�#�&�l`JJX��F^�:Tf���,Ű����Y����YX��Գl�� ���F�������孻6�1C]��Ҷ�hJ��x��Qη�8khRԲ�v٘%�tr$	�X<-s���l\���⺐����s�.ib�&��V�D��.��1����u�O1g�1ᶫ���m1��0f����0]i��P��I�a)v����1��%�JLW���	^��`��f��,%�`R��.s6Eї.��6�Թ�h�ֺ�6�Cvis	\i�/(p�q�rZEւ���6�6��ؙ���C&ZZ�Di�ʢ���.ͻ]�@MtwKi�L�g���\���tW��L��l�d���hB�A�:����u͆ћF虮MC5���4�d�B�		��ʤw�y|򚍭4T!�g#i\�+�vvUݢF&٭a,&�
�5΃6i4�D�*m�5��m�n!�Xm&�a֘�I`�4;@6fY�f�ۦLÄ�.��6��B�MI��%���n�҆�a�/A4�)4D�<(���,�.[��CG���Ԏ.��3/i��vF��v��M
H�)�2�ж�V��U�kU���u�K-F9��5ҍZ���-��͋PX2k�Z#��2�[3�Մ�mp�s:�i��6	�K��Éf�(J�]	M�i�#��A�W7m@��$1+).�h�a���Ů�, IW75�:L�뮥�`�
�[(&��Ut�l�4�.�b`lh�K�Ke������iiũ��� �A�ŕٴ�a(�Um����[�ͦ�ja4�tA\Ԫ��:q�1��$ɂ�F��TCl�����]45V��c��U�](�l��n�f.��\�&��X�`�`+�t	Z�F0��P��M�W�ˁf���X��-��Iu
UvKV:r�[��F4�mW"^,õٹ�,�f�1Z��\;We�5)�L�P˜`$m��:)�H����*6\:آ�.�q�V��.6�=U��j��u��Ih��٥�L��ˀ��,e��itLM6e���hd��1��K4
�atq5�4kڱZșc�X�@�,)�˕҅S6��sq
]��0es���y�ul�a��\:�VmW����̘�f�r�^�YFB�F�fUY��.��͜���#��M�٨�U��Rͩ��,��+Tu0�,�bC�4�;h��ؖ� e�,�F֝lafaXP�W���-����=���_&���m��a�m,�]K�u&l��/�^IL1�J�Z���Al�ƆiB1a��˭�y�(�]À��(�
��-��i2���$4�Ѻ��]&�G3@��)����
JCDh�J6�A�k�lmd�u�G@�	J\�c��bcn&҈�VM���3ҳ 4&��#5GZ8f�l�kp]�M���,K(�,u!k-�F�+��Lh�i((i�GKs�,�ԳZ��lK�VcM���Y����T t��i[=�n�Ŭ�L$rf�1d�ee��Am��IP�lqm�l��7�H�XV�rc�i f<&�V��P	fKki��6��lX�e�h�2��P��XK/g1�+לf�,ѱ�!)��L%.q�����,l�XFbF���vl-��l��X��)�`-�*"��m`�b�zj�w[B�l�;�IHP�[��1׆7B)tXB�m��2, T�LK�&���4��3��-��fI�\�1Zכl&YLL�Y�UF5�1GlX�̄%X�vaWl���q�ek)D��!���6m�7�M��^+�K-8F�1vZ�b�v��Y�eq1�bFl�u^M�К��/Q5x]Bڝm��`B���f��ɜl�[e)t`��
CJ�Z�gV����u��ԗF6a�a����[|���M�����,��t&4v%��݊��ⵚc�pO13��Bm�G���\�jRm���1�B�{Z@f)*�ܻ��MP���T�z!]mˉb�6֊�F�-f��Bl�V� Ve-�ܔ%WE�\ư���4ڌ2��1e��(�B���	L���3B1�wdͲ�֑�	m��*����]����\�U��[b��T�X�5T���B�"�ٺ �'2�#�ZD3ݪ鑵�H�!�$r�iM�0R�P��YMn2�)��˫	�K�-4��tv�8)���K&��B&Dn��3q�b3�eD"�aM+vv�Zm�T�p��d1a�niIl�19[\G)�B1hL��j=R2�Ҝ�l�bc$��!������f��͸qkj@��3�;; �aj�����J�V�fm8ŋ�)�jC����&���5��i��g(�*Y\��Q���ǭMV�5���\F�Ų��2�X)��R���f� ��n�I��^,a⌤�ġm�rۡbn:�����`�@��֓�*<�bR�r�t�	T�ײf�+���S13�՚�i�U���H���ɲm��2��+q�W4/N�4��U��h��]1�4�Z.0Kkc��g�X���6����u��T�P�+
K��v��F��J���������R�,4�#e!���PF[.,�<�Tg�ź�ū2\\f��I��iS[1{3lJ�u��kĩ�+֚�m�j 5w$�y
yJg�M�n��7M^s�V�79ԡ`�J�z���.c�1��5�����\�c��ۓT@X��k
�Vj�Օ̺锚��2�-P���saY^�+W[�sUca�(j��m�A���.e�60�ZY��S� �i��m��]noJj���p�pZ"��4�(M�(i��TL��k��ז�<�Jxɯj���R4J:�c�Dek.fGl���]ˡ�;F���؋cԃL��ٗ�c5�6i�-��喂��Yc)-���l�l��+������]�-=���<+�c�_'�j��h�6j��C�aZb.4F���.ǍDX�Ɨ�m/X�T���|�L-��˶m��,�Z�,	j�渍���ů��Y�b(k�����U�bn�ea��_(x^�c��]�֡4�lM�v%\SEy�"M�]"rj�e�_y����TL��*]�]�Z8Z8�T�Il�5A�t�e��⺦�
�,,g{  I���j�b�]�!���$���B����<}q��nݻv�۷c���	$�I��AH���%Hh�G�b@$dH�m��ݻv�۷n88oɢ���QX�D�5DT5`�q��v�۷nݻq��H	 B�3h����t��Yo�5�s%˴�I�[r����6�lW9B�]ݶ����3�m����|�z�۷nݻv�������BUU0�lI�"��Z��r�ꋘ���Q��ߍ�׋�U����ZLF��\Ɲ�(�&��.r����Μ�ݮw]ݪRK���Q'9&F��y��'7��K�����v�v0����M�.�.��w\YD���s���˕�MÒ
%s\�Lx�1y�^v��rɯ{��\׭��j�s]�h.�EyM�׊��s����W�k�ޭ��z��W
������`=Ur�����z�娒6�Ѭ%�{�5��sE����5}+�cE�y|��Z6ɣ<�F�{�sFѢ�BZ4W�k����w��<{y��b���[��R�!cJYy
Y����ծ�YgR���#e�"�pBL���P��-\Q�� �:i�͖��d�#��lauu�ڨ9�ݖ,�@�^.��3Q��dA�c��2�ّ�	׃K-�0��y�u���Ѥe[K�f��nS��Z�%8%�̨��ٴ�E�T�3��YQqe�b��f�Y��a�9�Ơ�WD,��JnKو�[lRQ6�-�/��	�F/��R�B]f�0k�,f?\��6�LM��\�-]��0M���SY��!v3,��[�dXG6Xhu��qx4mKaF�+�]m�"cu�ZC�s���.�`�� Wp�ݣ�֋M�LYs4p�������Xkl��Glh����q���c��إJMb72�9&[`�	]�����%�i��AaGDq]L�gh;M(-�K�9Z#���@ËftC[�s�v#5��֛#fh[Ƌ��XR)�0MnJ����ζ�bEm�Yk�]�sIs�V�&غ�%loٍRU�%6B�"M.h$Y5��v���q֒�0!S�Fۥ/m�V[�.�]r��Z��e����X;]%mWf(��eÖ	��f� [a����� �>jÖ.Ѝ����#���b�4�hJ�Z��@.&ͫm�l��aûX���uAn\�.B05b�Z�m��)���0 V�]�!��
c]��S�0��Y@%���/)� mY��XV�j�[!f�L���7R�X��;Z�K�.Ԙy�m��6\�e��İ"!ΊRb�,��2���T�H]u�9�6&§=\�cCf[ƭi	64*�[hF)���+H�Mɩ%Ia�K�M\lTƢl%�MT̵-�H���(@IY�I�:�a��Ѷ��.is������j�G������+0�m��⦹�^�%I�B����ݴ"%����GM�sH��%�Ѻ�`�Pߒs�ӻ�+�k��P��2��d�D�E �*�h@�`S�0���5���kjT`Ң�Ґ�K��
�%iZÙF1�D�XQ�iH�[
F�Z2���c��ʰ���ƣ��YJ�[��������*P�l	c�Ne���m��(U������>	Wr����~x-]��~�Ń@��5��� dnzˣ�֢;aB�X����m��Q�����cyG>\����Vn���м���H+pO�m��(�*�ӝ���SG��S�*d^��MN��"+[a��2�a�w�FK8֭}#�5JaLׁ�q�� ���V�⌸Sw�Zը�33"��j�����O
�jٯ6�o�}���W}\�y���݃w��	�_>Ϫ�ۭ2��O��G��Ͼ���:�<1��ze�R��7�S��Ȁ/v���'��+Ӷ{/o�ٯ�O|�Ϗ-�4�K�����U͉FakvA��ޫ�'NM5Qz:�HnL��$&���^���/w��<Q�O�>�x��.xxa��m�6�|p͹���L�FI%������㷄�`[��lZ�_�j�>ݘ{�n_Y�16.�V5ٴ�ݠ�3R΅u�J����r��~���^�|!��zG�}/���V��[�<iq��ɖϾ�Աi�=�B�I����N.[���lf��a2�|�;��{;�"�hp��\DA������Sw�[[��0ɫV����W�~>��}��Nٟo�u}bF�w��/-�wMfM�cUkTl	��P���~o^}�>��}>�3�L݁Mn%*S5f��]ne9���$!�+��98����c�P���ؘ���D]��z����f�X��31撘;-�{&vt��j��eɉ����w����X��c.�
��uO��&Y!����L)��Uǉ�K�ς���ր/�U�h��DLn+���ZW��983���Y�m�F�MOo����n�4f���钳1P&������R��{g=���o�rT�CMX��|R)|ϧ:���M�����lL=��=M�o��DF��lr/o*��n���7����Y-e+>>������n�}�n�oI��w�*>$�4�n�������{���2 �T	�:�!R&FƷ&v,ն�,Ap/�93 ;t��L������C,�W�Y3�p�f�����y���X �T�]�z�v7H*�;�ؘ}˼�^��{ M�wi��46�6�a33g(�t����P����k�ks��N5[(L���qHv�F=���uV�\\9�#�7���v�l�osNP��}>=����̽�WAn�y��K���5��L{�}w���zw
�{�X�i���v��efal�l�S�z���_�L�y��n�7F>�#4}u�4zݫ�(�ܻ��h�����i�5�=���y���`P/YBƟA!��$�K�� K�gh#��*�]+`�b��&pR]��a}�����~��z�j�Ϟ?��������^@�夬��[k|�hj�`�*��<s)�ш6W���P[��.r��a�����ۥt|2�o��whP�߫&��z!�a���U��ÃS��pS���ܝ�-˼�V�����g͚l՝Z���{����`�Ǯ�_�or�Ĩ�����f��������"!7�	�&P�^hS]z�5)�W�2���u�~�n���}U�����n��>�%;���]�R�
d��XCŊ�����V��vM1m�՘P���[����m��p�N�Ep7B'Rjl����T(P�u^;�.��MO�B�Сvg�$x�PБَ��;7킶���ye�;+l:Y���mmM-б-uHL���9\�T�A�M�6��ʆ"��Y�h��tT����!���d8⃜�v]ƶR�͈J�ŭ&�XћfL������J�0��K-1ƀ�3Yu�E�e���e���&�(7l%v��W��W6���R�\����`D��o��6j�L�y]5s��TwP\��77[ 2Mp�+�)3�
�f�&Cf-��'b L6�bd�͓͊��W�-5���H�:��[�w(�k͟U�����hk��V���kw��2���s��e	��f��b�˟F�n�� �Mv���r3�ss��L_x<$�s�n���e�W��e�2�S�ˈl� xb|45����@D�o�{�r%nU�z����s���+�Z���MJ�a@R5l���ɦM��f/o6�B{���^�����M���������o�L�Q�x_�(��j��Ԥڒ��f�0�l1��l�s���Ĭ^&�S�';sܮ��R�9�_�}w>�����f�O�MM>L�7uM�_��U����×�_.��lWc{30dv'N�2Ѝ
g�'����r�p�-��P��	�s0�@N���"'�^ �@�'1b��	>��}���;�*�Lր��]W=�j��_7C�K���|[o*HZ�/v&}	������۽�5���|�ʦ�6hZ��wu��:� �d����@��+̜�:�n��Q^�|8yY�4�ff&v|���!�*�صB�YWG��fG�_Pml�kcr�v��ߙ���Ͽz��{,ҥ@��L�FT�]�n�L7r-
M�r�X�:%���e�����o}��b�{���΢d�3�:3�d>�׽�ߑ3���^6����O�o�h>�+���F�l������������>�Vy��{�՞���+P�b��Ȗg�K��ZE���,�t㱦.nȶ���z�὿Y���C^$����J:�>T�Do����rꇪ��A�s}��=�݊}���귓��6}��ݏ�3�N]�.�	�eO�slk�z��/[f�f��>"���t��������J�2?�m]�e?��+����D�䚼����l(ki	�&v�`�DB��e��O��ib�Q�K��W��)vCP[Be�B8��<���w�l��NoJ	�36�\+��y��[���g����H��&��-{@��6s���m��?�w��������dS��%�#(R�ٹn�#�L�nN>l�[��͟�]��ڛд�M,�e�{��p�i����4ӱ�A���q;��ݨc�k�]��B����Gnnf=��a�A���3�V�=G��8�>`+�:�Q<�Z��/�+���[wt�伖����ׂؒ�fVo�z�T5�m�X2��H6Sz�W�Gnd�zP�[*y�x�ȷ8%�>U�f��z!��ʍl���3�*X�������4�.5b��#"��M��"�Z9.�5]0�;�p���''��at��c��*�oo��9s�Y�L�^gt�����^`�6�uw�%�_[�O4�g�ߑ|�6N\+��^�V)�^�s����-ZK����_?�Yѝ�������+�K��s��޺��L?6]hk�^��񬤍}��욾���M�/�|(:�5��#}�_3](�y�l������۟a�?/9�ۓ�����>�e45ˇ�3c_��7&V}��>�P��b�K9�LG+!�G�'8G���]ܻ�f�j�j��/�U����,#C����6e�ʹ2g���V:��O�{�₦�mX=�z���C�>�W^-�!2����C[\D�WBX���1�1�i���%4�*�X����͇�\$�,`2�Cf�\�
ݭ��VT�J��v���q�d1������7��4-��n3	��ƍ���ؖU��|i�N.��e�m6�+���A�s���Y�&��L����������32�f�;M�-�MY*�p�U!Q�I�b����X,!ya��]Bh��a�M���6"�U�134��z�	>���7�7�L%�_|���r�������ꭻ��uV���5bv�fd���	}�2�g��R��ow|�u��wU%���<4٠�*݉�5�&�i0�D<1�q�B����H���)�'}��[s����^�?N�W�o=��9:�w��ij���_5�-��3�������/�F�5+l�����n����f��#��nq�]&�}|����W��or{�����m:�ǒ=C<���={�y�~O?)�����n��ƙ�S��4���\�N���Cj�)����L��#՛�Us�����C�{g�1�A�	t�#�ۀM�O�)݇j�<!t.Ckv�;)�y���[H;���o�i-�Bl{�Q���yMj�q����b"���πYw]N�ު��CT��Q��|��]�ҽ��t�]Rf��wK�w:��j���CRF�����Q|	�־޾�r��l���|)q�ϓ%�i]؝�UWvY��Ҙ���n�-S����<�wfß:�ʹ�{I�g͚������c�z�<Z�t��|��^%;����}��en�*�v�iRO��>�������4,#v���h���ɸ�HV]z�Q�k�1�s!�����3�	�f|�RU���݃r++)��{팈|N����2��l�Q�co;�������<�N��Z���m���ksWP�չ��\u�n��U�k�� �  �0`>ޫ����N~��oe�����쾭�G��D̽��|p<�{�ظ�;k<���u�5]Ҭ���NLB]��,�yVn�h^?l�yj�f�Y�>�X[[�]��#9ju��D���w-^�/fqs;Vr�=�յu{-%wl�*�&t���Z��tV%:n�ǉ9(u��t��+9����U�R�8+3d\�M�;���C9ڱ4�aU!}J��ܛ���_
��e��m���ޫ��ނ�(�1W�է�1�{^00c-Vd˷\5Y�#;{&ie���zL��lgJC8IVW9��������٧��+�C���zb���A�C�G�c���@�%9]`^�ʤOMy�w+:�F�vt�s���#Q��݆0�Z�n�Hr�[J�5
%�t$n�6�P4���dH���yQx�S��!���#"�j�h�=��M��O�G�6��n�[��!e�]:���>T��;�����	�[u�L��Ҥ�V����Y�6�ٺ�-����ra��Zr��Ν�,��^�5�.�ھc����X���M���dS�l�x�٪�oܥ۷�Oj�&ӱk��av볭ѝY��Fg*Â�U��B���@��k^f���]y�>JV*P�Ű��ֵ<�.�?*�pd���B��t����;�X�G���`���[ca��SM��
��Y�}g��s�*�Ҕ�8yQ���AS���տJq5��[
�]>zS޳ư%5���Wi�r���sZ�����]F�A`#�Ԑ��d�Mo<�{�~�����F"�
D�H�(�L�E �Qa4��8�۷nݻw�{�|���x����60R@F�l�(��r4`tF�,��H��o^�z��nݻv�����Ek�:��jC�E�%���IQ��2�}m�뷯^<x�۷n�z8��tF�5�K��zܢ��6�t؋��E�j�U��|z��Ǐ<x��ף��pD�	�Tm~���s�V񈤃oZ���d�����[��Dh��b6�m��Ӧ�j5�F�m�FɫƷ5���y5�mr��W�����-^���}7+��QTm��{�y���h����W6(ѫ�U��%rܤddJ�D�O�c�0 ;����sG�G��46��JX��c�Rv ��`�Ɂ�v����>y�gh v��ާŇk�1����uGw���3d.,	�	�,+z,�G<F9�����D�������ApӋ�X��sn�����td�d>� �<�e���>��~�Xz�<GJpX���^��&/�p�%!���q�K�8"�hL])�%�	���5 �&1�38q�t�x|���|����jik��A���r��ݼL�z�3�,�aM�׹�ػ�f�L$c�u7����0�"�8!N��v�� ��vEk��'mjz����3��7�E�M�ʘ�=k�C��J�7=˾�+���|�c�뗢ɶQ洚a�Ƈ[ޭ�gv\��S3y�ǫO�6������������7���X���T��z��Rgp0���nT1a��My ⧶�;���G��9�pv�����5y��E���}-��vp)�WlOQ֭{u{e;�k��=�r=��Kw�Q����o.��&�[R�f|��RRR�S���1�dG�]g�=��Q��։�Rٽ�q7�[��}g��L��{�gnn����u��&�&#%b�����7�)�6W�kf&���.���j��k��f;QM�X���W��y]�^���A����L�Ry9���EW]��EssCwU<�0 ��b�p���0�&UJj���
���uj}�;� ��5��=�Q��
���9��;�(I`z^ص�)�/6ޑ��&6�ٷP�,6ӐES�pES�MR>[S�:�0om��m*�1^�CZ��q���vJu0sT��\������ܪ�4�<�U�0n��؂'���&�g�q�����Fb����4R� �;������;�	�͗AٳSs�RA�F�Q�;�P,ً|���pW�P�Қ� rNٵWQ������91�=(;����R�(9�.2��˅��7�ܮb���3���ַ3����eu��Ñ���2�O��E�©��FF�H��M� �V2�ar�a��,X����țFTNi��Ѐ��V1�X�^B`j�%T̈́�.ˢ5�"7\�VV�RV�)l�B�Ixy"�n��MPԚ+��e�K����t��cYfZ#Z�)M��v�E!o^p���ūc��4a�¸�U
�$�����6,�Ź,-JK���vv�����"��Ie]��0̽��f<\ܛ�+B��#3(�g�/{K�t� U��N����y��O����vX\�Eq�5F�Z&^%����ɚ�J �^.����"� ��8���v$
���ov��C�Mz�Pܘz{֭�ȓ`0�A��_]�^ �j�Z��Sf�F���ܭOh��qB��C=��&����o"�S]x���v��� s\
��U�5� ��k`���ix��^b�eT������n���wr��`0��.�Ξ��qsy���7J�
�v�E
�%ՏR��ei��BP�s�.<<ʣz9�i�a� ���h���4B��A��D8���Χ�{��^p�bS<��_���XA�N!�v���L,��h �v�4e�)Aނ�@���=1~���/53]�C=�����<��E;��4������ϴ��nf��)���ԅ-�q̣)oele�KuՊ�.��l������X1�j\G��L�Z�<�����%~����\�ѥj{J׮)�0�L}B�7t�`nd���&�4o��)J͐�7ûG�όt�P���ɋ14)ſ�v���Q3a�]�SE���b�fR�֝E���o>���T3�;����J�w��J݈���~�Ս�0�x�c��u��)�ev!�*����TK��N�k&t�iZX85K{);�Ө��f  b�L�<Q�c㺀�0�*LѢ�Y0MN�Ư"������g7���ML�a�{L8>.X/8,:���d �f(,'#�j��GN���Aƈh��C˗������������\�g.XSp]I��w6z�X�x[>}f�b�9w�4C��Sl��7D#��C{8x�>�f!ϳ5�O�'D<��۠��ŝo��� �:�4 �^NZ����j+���aS��z��a���#jj���ì(�"]Ý��
��
@f��a�g��~{�&��n:�ޓ� <`���]�q���L����\�?j�׫���5B��͛�bj�eT��&);�&��L��Dc ψ9|���� v��sdr�{����A��p m��Q���4�3��L׋Ł�p��&r���glr�;p�z��e��`����ou�Ų�i�gBW6��gZ����G���vr�3uή��s���@�p���������Ng���T�DJcIM4$�$�P����\�l	�SW�n� �+S�L�T�`MRv�L�&�t8����A�٫W��R-�r�8�y���gkt�a�u'`X\I����F�p5X�H�[�i���&�9Z!��: 85K�P�3��ʸ��zӋ���Α����3��G�Rfq��] ުqv�+���)��GC�r�@�5L0�A�)�@f%/fg@�e��\3$#��}<�����Vb���p�T3�T�r����D�hQ5y�c��V�	�Y��� ���T!fӖ�r©9d�T�1a��buQ	xCO�f�
b�.��`���̎<�j*�B�8�A��V!lX]�L�c�l �9qa�z��瓂�E�����'ǋ@U�՝[�� ��@H��3��9]�]�hG;۩-D!��͛,�8qL��g�[� '@���vF�b)QU��K��t���tN�`��>��d��\��~Fn��j���F��xE����t]-\���+}Q�.���v]A��L�i9�Uq�6�dR�/��@&M�۷N�ؤ�i��j�~5�g�C��֠\��׌����I�����F���\��V��0p���O�4�}������(�&g��a0�wj�mNw��U� n�P2�r�A�]�ˤDB:�imYl��,˒bRi�DB.��	�1a�U'��vrRpY؄@�Nՙ]w��ʮ��3��!��Z���l��aLF�`�gP`�N�U�v� ��.������鲯�aM��
kdi4Zex㘀��f쿻�D<�恎���rY�Bm.�@�W<!���fy��Mj�L7�h��2�D�����ŅyN|����I"Tflp:�OW�u��'|���0pDS��H
�o3��گ/ML-��n�;m�5R�`MRyܽ����WQu��0�(;J`���ow�8�y� �&�dd��0�d=p�	�e�.�
��4#׆}�:����w��]�˄LU�c� ��v �j}, ��ڎ�\:x����s��]���+C���1vЫ�t�Y4Jq�ǖwr�)V1�B��ۗY�����(f��9�:t��Y�e 32������Q��U��� [����e��n !��/�� O��B<�[GJ�X�YEr-+[�S�tܪA����6o9�A�2X��z���v�L��K�S
E��ښ	1.�1����ZQC��m��V����E�-˂h-��J��mj�ҷ�q�),nF[������]���:(rf5шM�6�(R���v�:cQЈ�������S�/��%k3|���V��h]��X99(��ɝ�Bd����������1K���w�)!;�5�l	�sG����9�Sw9z��}�YZn ֐g��n�� rj���r����k�%Nr�X��lH�pA|)NI̓���8vJ���	��s՛����3Z���0� s���vk��~���K a�BD2�`H�N�������U8vj����wDrx4�S=V��|�ڸDׯ4u���LX�;��H�����n�?�`��{e�y,f8v#- �T�n�c��W�o��+��Bk��>J�S��n�CWDbo�40��+�y7��Rq�]Y@
����N,���Em�TǕ�*K/VE��)�����_�6������u]M��9��Lw��p�M' ������a�3yz���dl<1�x0�\'�Pc��]��l�uĠ&��a b��)´��|��")qH��Y���y����c�#�Ǫr�X�) �JژN��S�U �N����DƇ�-��wϚr�z*fկ���k���Ӄ�k�����mA�����3k�y�;\#����k�8>6&����^�< �pXE�"	��@!M4��AH�4� �`� ��n�<��!�=����Wo��Խ7�x&&�;t���\
�=hS3X�9�Nŧ8MOD;�$5��'����6�u]]{/4(�@��Qd<h�G�� ��1����}��9���K��'���R��/u�upz�M�c�1G�Y<2��xrْ¹��h6F�����C�*������ѣ����H��h E;��۬�'jT�f.��3�<A�p*���h��O�Z��(x�`3�F�&{�R5ke�15���R\��t3*����4�	�o+��u+�����Y`�mc�<�ue��wu�������I�bZ�5y	��> �����"͗ ����~*2ŀ���Ey݈��S�����C�zo,it�QR�'HsT�2v3�J!R���at�3H�v�G�m{���n�����?�};�bc+�C�9�u
��l�ý�������7As�k��Ϸr
�suv��ȉv���ѳ��T>���H�H�4�
SM(�i�����H�k��S�m��=����_ �ŝ�vj�8v(R��Rh�b%O[v���P�HsT�X�)����7����Y��G�(8"��{�7�N���L4[©������cކ��G�9
�=��V����n:?�9t�7I؂�]sC��k���}�p��ٰlKcSh��:鲡P�nE����m��ea�A���L�@��Aۙ0Nې ٲ��	*�nu�5��OI��Z��8>�{ 㿵��3�.7.W��S�g��5I؎YG������\�;i��'S�̾���Wu�����Ǆ����g+k&ߒ���A�3D����8'OT����R�*�G�^�ۺ�L�x�N�ݲRu��m�W\��y���	q�O���Z�I|�G�o�ml���1(;4\��N9z�{K���=�����G���Lvo������+FA���@ߒ�����d�8��M���2��kmȩ��'�]��U�9d~�Ǉ���W�x���0`o��dԊ�H!M4dT	I1U	 VAA�{tc�8��|C����dVC��B��A�+`�Ǌ��]o�z��k8x��7R7O��4E�16&���B��d�^�����l۶B��8U&���f�e��!�5X&��[]��G��hC��Ωߛ����E*!��Nwi���j�7��䇕M��P^x�����oS�	�NMJ�\ i�q���Fz���s]8���E�׷��."{��3�`�I�N�ki@U��;�fc���`���/b��A66d7�ඓ�ً�#���X5�'��P)y�2�u����h��&�R`�n��i �8�U 8���0�@1b����Sit��F���I�=T�n�]JxW���X�:#�z[)8��r���
��b�1h�p�ݡO�����B�1���K�����2�pO|�L#�Ѩoz��N�Z�!>מs������\��w��=��O�G��G�㳴�gof����$B�%�{AwK��/�i�B��ܷ}������G�n�d���l+�k\�5��7zA��m�}W�'�xu�yR�
0i�G��+Q���pS����s�g�nS92��.49s��{�d������V�<�+��h�&�����u�.U��v|b��n�}*��&.��ja�(�nLU�}��D��z6n#�򣾺	q�����ͷ}|�VI�Y���i�Y���W�@&�6.5���b��lŇ��G��ZJ�l`g��;姅g�]�́k�k&S'�Ky�t�l�ho`4�Z������k{�]�-��@�E��vX"��;+�]l�\PF��ͫZzs"��G��q�ə�i�܁:Gf��6���3i.���i�4+^o+��K2kU��,��l���6�b%�;Uc��������4�YV��D�zф��:k�o.���,S��h��'��
���N=.����Ćn6+<A�[C���r��Zv����ɼ�����ה���sd�ʞ��G���ݟcy�1�qZ=g'jY���[�yp�R�]u:�R:�ڷC�!�q杔��@Q�����;\���3z�]]�"2"��ѹ/36fF���
�z�J^f��&\[W��z��f��h,�bL�XO'>"i��8$�.�/jP�e�h�Ցi#����OX�#Ac��q�p��p����7�J�D^G�r.)�B��MUA��^�~o���Ӿ%c�LH0�G��I��/��xcv��Rz����$��e��R�LU�F������q*�cm�|~�<x��Ǐ<z�qL�{5M@*�H:�R�m���\�����;���sn8���o^<x��Ǐ^� I9A�o����Z�o���x��j���|q���x��Ǐ=z��j��Q��1X�j4�=����m:q��x��Ǐ<x����N4�ITT� ���M76��\�W��Ψ؊���(���:E�����H����F��v,m�˘��nTs�s�QW����W��񾦟wr�W�tGMc��,Ex��;nh����lV,F�r�c�D��F��*,Z"(�w�y^5�ڲ�X��m��n�V/��b�4\���}wTX�H(��s\���uy�bة�ۮ������^��<.�!���d)+��2�7z����7@�u�A��-�h��̪�l�V���(u�q�����i�������P�W�m�,� �vV��Z̡qQ��s�����+�R��m�rFiZ�`hT��fu�5��l�����vA��ҍf7�M%jUq���&�ev��Ԫ�8�̯n�љ��@��%4[ہm�F��Ei�mufajDfٳF��x��^�2y��ˮm2�����\��2m�6�U�%�I���t#pP�5�lZWb#z�J��K����l�vn��ô[j!x�K�Me�k±t�)f�3vm�)��v�K.�a1Q���a	K6�F�IRh��&���%꭭Ƈk�,R��ך����Qa;k�%��ąq��vu�,�,pB�*f��պ��*�:3)+3v[�Z*�aR�k*JFፕ�7fU�K�vA�ii�C5�S!R�$�,W�k�uƠg2��ck,�1\ԛ.�1D[K*�i�z�f+.���-�,n�҆Q�Z&��뇨�r���tmuc��6A�S���5��en+�%rK�Y��Pl	�Z5B��%��t�oa�mX ݆�JB�jj�ԗd�B�K�:�c
O	��_<n�´�T�iQ�K�Z�=�С4Ux֍!u���=�6܅�iR���M!	�@u��Ԥ�
;W9�L�`�b�iai\��5E�K]��`3+���J0�Uư��&{Y���i��3Y/RДXa�R��f��||KP��ICg�F�Mn���-̗���Eݫ����6��%n���!q�����u����i��(�ÝŘIR��i�&��\�@���κ��XZ¨li�2�a�R�2�QMeX\c�Kb�r.e�U�GW	k*mV�my���Z�b�sqbmۋsE�a���$tuoW�K5Ņ[e�ՈD���b���Ua�s6Ք�%���ӱ�?Ai�R��F�A�hUJ���*	"������W5��ET��,�MF�4�#�`��]q�v�=�3f��@�B�ٵmz�0JC&t����v��44H*	Z�K���h�tk����H����F;T49p�]����u�ZGRֽ{0�z� ��*Ų�3&�%���P�fl%z�A��;%Ӯ �\� ܎�W��d%2�)^��-j�9��;�i$����7T�(Q�7j�˸�iF�lj�%Zܬ��3(�$x�?|I?=�al�f�^T�o��v�u��3/8O��۞|��B�!��E�s6�����	�ߝ��\����3��|j�+DZ��h2�����N���n:<��'5S�zk�fV5R�d���R2]]	X�R]e��~̓�d]��-9�0g]*̞e��	� ���]˱k��s�ms=�W>r��[u��3i� ��N'���w{�.c.�p@�ր�����V b�P�	�A�h9u��)�dw�������֋c�K�s��\o�*f���. ��r��85H
��2���<�:.�s�z��\PQӼ<;�4������f��1L���E�بgJ	r�8I�@��)��:��6Y�ۇk{����7���'��&>A�A>�&����$����Ր�L�&pj��7{0^Zw�=J��ۻeӕt�*���I��GqΫ��<GVe��0b��h�ͮ��5$�t�
헵�Q��מj�d5�I�����*F�R�
$�ƚ�i@� �֤����N�x���^w�ʏ\e�@�Fy7y"�4h�pn�<���fy�8h�� ��9N�#�w�v)�%V����߶���[�,	�Bڙx$�Y�RŮӂ,ۆPoA�56��v��52�F������s]Πo]*��g�v���F�B�K޸��8Rl,iij���I�
�gcT�:�=���ʤ/�u]���yw�_�� � ��%N�T��Q�).�ip�g��bX�2��r�R�vx�Rc�Xh��\٦���Ͼ�M9(9�9N"fv����g3D.7�3y�눹�ϵ�H�|��b�3����j�Lj���A�^ä���sĶ�M�x�+LU�s��OW��;����b`�EQ�X3���xUc9�7��C��B<�%�g��(��� �?�I��xsE��6���붑�� ��قb�]�zCІ��)>�����p#�
�o~U�록פg�m��NT^�=����Q|~4�4�
T@�4+P�@�4 �DPdQ$$ ����>���]C�]�3�	��A�-t�ȪA�U8vU8{c�__m�z2lL, �w@�7؛�c�݄�(�3��p����NG��z�0$'54���A�Bb�qdU.XV�lw5��8���w��T�y<ϼ���NAl��Up�MRyY��A�LNV
�
�Ä!��5im ��V�4e�.2���	Q��=P��MrR�8���]�u�W��(O�I�)�]ޗm:|�@U ���=]d��e�a��(��%�=ۚ��S�Χ\[j`D�!�yH���=�#K`�/T� �8�7�9k�g4a�c��[3��C�<����jr��=��a���{�㘀�Ր��]
��ֲ��էz�B����P����m�Ga{̬�g� �v���k���ہQ7׾�{�֍s���|̇mD<o�s�ɘsO�>��Ė�ڏ����&өb�p�'Z��*��v��F���$~4�4Ј�@@�4	PPIEQY����pA�b.�c ٲ�v��I�1�ǯ����K[-ZC��;��.z+���:�qm��I�R�,|�n��	�>D	��}~�JgW:Ilm��kt���vV7U�2��P%zBO���@��F�ÃF��LUS����׈�+��#Yoa�1gv�v5�"�y��A�z�5>c18 ��,��o-N�����^wS�_`�Ύ���Y�$� �� �
�ƍ}"{�ļd�U�Ø���t��S�Un�B�dt٤;�_Q�17���A��c�VaIp ��L�U��9��� P�W��xT�e�qÝ8@r��T�Ǫׯ�_��T�^?X!��;�K|�Χ''���x-�&;p�F�Bj��My8Q��+��z|Ǽb��q�[���;ff^p�<,{PpXUM���yx�jk�w:X����
�F*�I�46Z�GA
?Rώ������w�&n}]n#[{�:̱X��n�JT� ���6�X����8afl�g.��� -?c@�A#MTH��\ڴݻV��j-��T33>���'~O��O�c�U](hm�UZ��G81C%�i���ʄ�WmB�֙��xjWe4�#�3XTZS\G^	R�,kmr��-e�j��]ءZ�MT��kn�uZ�7%P�ܔ�ۛ�2T���H�
��f�n1h��M�B�T5c�Y�TP�i�q����[��jR�.�`.Yp5e5�e�}� ��վ����]E]���D<���q��@pjVV0��U����Zq)�ic��Ʈ�) V�]�� �6\v�8"�ݍ*!�׳��C����Y�.�����ZS�r�^����6(P���A(U�-��z����3�\� �Ӈ��_\lGA��~e���i� ���{��iG�yԍք�C���� �TXx�����eE��n���ݷ���31{3/8Y�d	�v�� ��p�B�S�"����Maט�h�r*U���b)QW���~��^^P����-�9q(�c�m�n��	�,�F�5H8֦zb�3�%p�w4N��(zwׯ}����̷�s2`���n�����w��a��>���Ϛ\K-��Ci��`�K�m���$03�͹��c�R'i�N솛"�N �'}��;��يr�g�����{�C�䃝+]ÃGK���9N� ��߈����?o��h&�������ζ�r9CS�������_����nsT��u.>�wW5d� y9'(8>�� �� ���2�CpG��B�����{|���ð�ߍ4�"SM(�EcM"5$@@�~6��vό.]����0&�o; ���yyM���Au8b ��cT���q{N��$�[f�wPۇ)S��
�8N��^3a���ʸ����\�x;a�p����;*TDks>bk���[�T��"O�]�1T�m����޼����`�=�8>c��vS�'+�0,���4�Ӹ,ERpERXUON.�W8���8����<����Έ\ � ��Pa�U(5(��d
��A����H�}����%��뵉�°�
6�2��(� 0��f�<e ���M�CM�V�p)�6�n�=\��Z�骞�̷���j�>�W�;��k����B�RpA�9=.{�^�
�����׵�;{�^�'91�����&�;T���{�/�`]�;c!��"�8NR�	ow]U��m��V�,L���Xk{{��37IҮ��v�W+��*ބ��5o�U\�Cġ��QP|8���y0�K�W�������4ҊSM"4�SR-[Tm�m����T�����z��y�Φx�m�r2�R�ƥ9�'-T��3̡{>�l���d6D"19HV�β����Ϝ��1��u3KJ���y�=BȉwbbY:��)ݽ���)� �v M'��ѳ$���58�V�k�쫌��g�9�ZERI�Wn�\�k��V�bh���& $
xx0[�F�ZV��slՄ����̤��4ߞ�'�4	�ˡ<�� 9N��A��'��z�����e�q笊[�k��t��7I��' �S� � �k���\�۸ ���A��|o7�z�.�pv'�#��
����uՊ�G����wy�Xj�=7B��lP�!��a�А��~�םm 	
����R�}�s�,`�^#� ��:b(��� +�9��B<�}�����&A�`9�{b,�Wy���]bs3��	�� �x#9��C�[#�{.�cг��3�����]�pJy�jjڣM�yWK^�@�f䧕�)b+�;w:	�.��W�{WW%k�({ �ƅ����B�hU��Q��"�H(H
�{�_!o��^�z=|�J�H8��V}��5V�.jo���SQ}�F\�6\�1��� ܻ�dM�n����c� d;�8���0�ЩS@�4b$f]��b��a�So'��w�a���%aj��*Oվ���O�8�Y<���dw�#��_�ӡ �l�I+<�`��8pES��j�v0�-��V�ve���N��vv껝�o��33���YU' �g5J�2n�B�y3,�C�М1��wPpAoU!�@=S���
$s�ƽ��ަ��3��y�M曁{Ŝ;�g����N<K���TFӻ8m;A�N�Y���<��2''��n.�N�U��seG��`�2����Z�\K&^����z����H� ����+]���^op�zL��g'\l�q����&sT�-���C�@��=���v�=�YΦl4-5�]��I�t��ك��~��L�j.�}�v�hV@M��9�5Rj���h��� ��B4�ջv�j�Y�uZ�Z�j� %�1,�;8qY�g��K鸐`0�X�.�Rg��e Jj\h�鐦��iA���Օ����64]K[K1:ɛ��eL;���k�˘ ѭ�G��$3�m��%V�0������2bxCru��0�"��˥ ,VGG��44\My��՗V����Y��d�de�4ìk�hT����K�hn8����M�	����ɨ��!: (�]�ӝ�|e�8F}�e��~>�������+lHb77M��&b�Lf72�hR�tn)�g�@w�=�����}�B��j�<�U �r=�����bs�ċ�U�P(��n�R�x�NE�ᦜ��H2ۯ �j}��f�ߌwf<�>��v�v"jYô2�@邽�]�,w �l��t���I����b�N �^�ԓ�;��H�Sw�.N*^���P���rN�j��A�N�!T��K�\Ů�xb��9�@;]�}�5���}���'9�-y?�K�&�Ĭ��e�F�fiӍfU���(�ِ�6�D
D��#r����o�~u���=��p ��4�ªBv�8y��={��z�*�t��pL� 4�c�6ц\E �5���J�a�&z�=�߰ߺ�1	:�9N��5���V�����+26�MO�ݨ�R����@�9���' �v�s!����!\�e�������j1�q����de��1`���־�\���m��ޙSdHUn}kK��)�S���g*ss�M��˛��Q�j��hj ƚ@���F�
X,�Sv��Z6�jŴZ����������u���L\��a�FppO� �n@P��.��g|���' ���D]��0nӖ�(���!���nH0g��<���-NO��Ac��y�L\� �U ����l�ګ����3-4�u�v"9݈�v��̮]'T�VVd���s��B�ם�y�pٺŠ)���Qּxd�n�rN�&7�/TAxǱc)��ܞS�>W37�w�ך�'C���&�p*�ıB��,���?}|�����61�����R�i,v�!V�%�m�v�h��f�slO!�濄��!���{�t!�Wj�T�g����ŕ>�&}8�����`����p��Q� �T�Mxj4b��/!f��G7Ƙ�Z�E�#k�w���<�z�/9�<u�8���_��_<�0� ���D&��@=S�2h��
�<�y�� �⹠v_\�9�ŎכYz ]�-�3���%�͡�ɸ,�r�ͩ�;��go>����oP���WB��c���t#c7)�ɸ���طs	6
�Җ��X�]}�ް�f�<	J��n��=7�3�����ffv��k�7���gfd��h��3X��tu,�'__h�iVz�+7���V
f�FY���ل����,��烬��.�.����Ή�:F����q�ô(e��{�h�4˕`�Z�|z�U
!L=��A�()O3hN��\��jr�do>�pVNЅv�W�k�r�#��#�j������5չ�3���ݗ�dl-��n�vX���w�p]M�fH����=��B�)u*�n��-���xa����m
]hɏr��ּ�.��	r5.+����Qy��+l��n�6ﱆ�9��Z;��ڳ����mmv��f�s1�����59r�1����8�ƭm�����>�Ӡ���#y��կ���A��z��UP1�f:=/�Vۊ�C3n��+���wT�mMj��L
�h�9���՜���ܩ���_�7�,��0$Fm�1��؜'"][�6���]���2�,�:աP�s%���!�{z*򮮺3ot�ݎ6�mq{��o��jγzӆ����ܚM8�!�^�k���륦��lW�e^��W
��<__# &�o��ei˥���u�ʅ����4р݁�e>$Vd��i����t:�u��8=j�"������5��	��Te�$y��n���הk�G�{��@D׵#�P*������F���xD��޼}q��<x��Ǐ^�1��k��J���r4j�j�HjT����	iӎ>���o^<x��ǯ_z�`�)��C�Pu$m���b�2��myۭ}�������x��Ǐ�z��hj6�*����]n[�-��~��"z�m��Ǐ�x��Ǐ�~|W�v�A������-8��\���z��[��1�˕�طwo��+�M�nj��H��U�h.��ɹ�h�UԨ*5!�{��o;��#<�QVy��y֍��A�Tmr�K�F��X�k�8���c_V�r���4��_^q��o�x����_kW��p�g*��*	Q	ڠ$RBC����JShһu\*��v�Zn�n2"� $�g�d�%V_/�w^�W37�z�8 y��V8^�h�R�C�ϖM<�"�!�bpA5J��=��8�>Mk,����.o�Þw�;�V�Z�8"��8$U&wj�aUm�2Uqyl�۝W���=.��/9�sj�#�7�� �19�*N��!�מ�B�Ͼ~~�3�����ILJla�T�f�R�4a%�Z6�W��(%��f����[ yb.Ӟcv��l�ޙ�/]�vpG�0Tw\m촵�m�8\�ōR)���YnӇng�/^�5Ǳ�$�%P4��Gg��)ǹ�e������y�6�h�2���P�zc�B�4p����U&qJ����/�&vj��<}�f�/9�p ����q���Cc���5��~��Z�|33��,�Nn���Λ�����zv3|��8[�x9��S����H2����w &��A�����)K��3sD� �ٵ���l�ҲMܻإ^�̷�|P��߬�O���z�U]K�(���e�*� H+� R��H�@4�B��U� �EK�e��b��I��kY��j�pn�SK*�����sK�l��El���4�7����Bd�-Y�-�ph�r*���D�V}p�:�{�/d:;�ZR:A� ��Өp�V��b]I�͡��-�$���56�M��{�����>���\SPA/b)Q5�|�;�\��y�����f�mB0����*L���=��i��k�RZ7���2�c�K��ng�N����~�âX���j���ij���؅~^�T�j��v5I��y��b�Ń�P���s��U��z{��b�p@�t��@�p�Ѣ���z��r�&&�lz �a��k�<�vv4��q5�|�;�\殳3�
�qӂ8G�J��n�"����k�<�S��A�5N�jL9<;��1>�P�p����/fǽ^��i�!�8Y��4&zTF��2	��~�A>[��eݥ��eݵ�؜R㾶b��4m�C��:D�	�6��-����z�}�d�S��I|�]�n��<�X��s�W�%�M���UE�4-4�4��I �Y�C����'+W~Q���Yn[�.�C�%�'jh�p�k�����;��YT����W��0W`h
q�6h5��ؽ�eڅ%6qf�+���VƷ5l ��5i6����9�06m*�`�������
�V�;%b� ܲ���t�K�[<�Φn��#	L۲��"91p�1.rg`Ha�B�L9��Ձ5�����&��l��Zg���<�g������XĖ��6�C�.+��
��,����R�m?=_�C�۽rjr�K�j����;�=+�б5L��>C�g�8q,��.�tȚ�pX� �Xt�){Τ�<�V�{�g[W�s������:|���Ny��v�%kn�F=H�j�,Ey;1Ln�v")5
HS��ުX7T�JNË�Aέ�W��=�^���� �N ���%�S�;[+� �[}��bo��X��A�P�sʘ�*��Ώ=���u��7m��q� ��n1�@�W�L:���p3��a�[���\]�8 ��pAk�9Ok*-��;���^���{���^gO�1���;!����@"�ܮ��C��.��H�gYH�%D�׬Jmv!����8��a��֌�fp����^�g���{�jA
wi�<"���d��:=�_a�B8^[����{ˤ�"�CT⚙z�E&��'S���#T����W������t����d>������זv��,z�wEq��o6��Q��S�%A���<� ι2dH	�]��<rQy�;��o��7Z曷]
��n�1��ֹZ-�-@ �1�)���<f���>W0>{>��G;���FB���j�./x�1�>��{c R�ƱwL⩐ww�"�7�����^{j���tb5~�́M�H��5T�1JX�cn�&���.Ԃ�וU�=5�����6U�)��:���j���5t*q���7PAA���m���^�<�m�oV� ���edt�đ:Yñl�g�UJ&).�PR��Z�;�[����FO^�<s����d.`Alw�C���W�D�G��
2����{($�;��%�4C�Њ�q-Fd��A��ՙ:N @.䇆^#��}��:�
�©�涅���y*�e�w�e�3G��>�^XNA.�6c������cT����R3kR���5�A�A�h=�No�9G��}��ԛ!7��m	jnp�H��l��1����]۴���9��g�ĺ�]5x�DM�ś�T`�u$]deCSr˚/V`>Hw^Iw�����u��my������u*'e]��Y���
o�0D$i�j,i�i��j  �O|������=���_�AȚA�RERES���"�̤�xb�S�$� Kݻ<�P��~�J�&� �ds���[�x3x�&g�����ԝ��NU �U�v�C)�iz7c���4��ә���=s�y�I� ��h]�rAn�=>�/��-:\K�wz)@J��FE���
hF	i�1m�֫V�6pLSy%��?e�_��"�3�T�&AT�	�>���~�����0ǚ��ӱO�,�=}Z�ψ@ �;`{�b�-EÑ�S�E�v����כ�Ⱥwb�-��WP��]Е^M�@�+��(ԧ�1K�3¼"��S��a7�ij�������A�/IËƼ��N�$עf��r��s�O3�`�s�(m8Z�f�K]��瞈�OS��q����T�k�Uv��)>VH��sL�DŚ�<�,�ʣD�SU9X��Ň*-�hwS駇*r�Q�3��7�G�|����1n{p]nr�d��5�V��b�����~Q��y#񔑦��۷�Z�aX�'�_��}�F���"X�ӂ`�v#̮�8"+�N�3�X0��k$D�ͳ��^���י~�/<`By{}s�k5O*�3�#��~Vo���`��0�\ږ�;hB�hFj�m�-:bPVWJ �
	A tq�@��A�7��h��T��=X}]�����g�wc��=���-�E[�1Z�5�e����"��oI��EC�Q�FX�����k`�����
'3B7�n�r�$o �lߙR/�i���P�p�{s���j�8"���XE�}��]���lzh:t������Ye��s17L�-^M���N�'�Q�@�S��"��X���Ú:Y�e�eN���^�ì����:D��Ǹ��p�F�,)���Z�9R��%1������,w��{�o���U�Ά.o�,n�pD�ƍ ����T�>2W�����
׷�%+���.�#��-AXv���3��F�P���К[v\2��pJPn?��	�p��6}���U;�%:E����ɒ �-4��)$$�d!!�9���wτ����~k�$Lb�u����),��V�DH���ck�F��K�(U�3F�k�4ټ�p,ɶ�m�2�gDБ��a�:�Y5��W�S8-桱V�)4�շq�h	i 	/Mv��5�Gbi�6�du��]4�����fkYQv��M��Y���Q�b�C3f�x�*�� �@��̺�1��9��P-9��>o�~���_g�,��YYX��Y�n�V�q�#�5�5��F;�@~�pS����kx��y!��	�-j�q]���9u����ΙM�S=���cs�W�%��8�k�ҠA5N��q�����0������j��&�z�r�W�Ot{�^�÷ ���pH�NŁN1E�fa�6��!Z�7W�&|���j��	�@f�v\���D��H$DLL�~���S�����%v�q~p�U'�`�T�2r:\�r��
�rg�z-�����A���`���^�&��ep �b����Y��U� �w��݋X��n�qh%n��"�'޼}:'|�NQ�fǽQ��<�Hq� � g\kB)��OT���B|Ҽy��I0;�!"����8ܨ솎1�m\k�U�����/��}y����[H�A���ǚ�<)�O�B��m�gnQ���Sy���*#��MF��Ǐp��A�`j�85h;j�"��5���J5�/n�LR+!M�L��*�]�&4�v�����"��-S����u���}��	��Q}�W��1�({����������IM4�E0�4�DcH���{�����;�٧~��{���w�pT�F����u�+n68�c� �n' �w�r�NI��q>��^���ƯUO��z�=y����|��iÑT�Ʃ���r�,�葯~�Y�NE�H0TS@�vyP����/ӵ�^�/��B�������yY�]��Ͷ��3�U�4]�M8pERcR�ד��wECAy3.d5Y����ӵ�u�Y��b��N�˙�j\[r�y$�������㻈������枨*� AS-�v����hb(����"ʱn���=���~ُ�,����{0$� �5{Yfzz=S}��	0�sf,�Q9�����]�W���j���3�b}p7����D��F1��,&�܏M_W��N�z��c� Š]�rR#=��o���R�9����LR��-v����iVq�F-v�s}�(
�f��TH]i���E[�,�T�����W�ޑv��asۗgEd#@����f�z�P��}
1��ق>�s,@,Qd�c^��S����=�f&�����&v�p*�5T3�K$iӂ*�k6�GD�g ��E2sz�1���z���EO�o��	;� �Q��3�Yh�FK�R�t�x�#7��^r˒s��_�\ly�X��Fl'�ٻ9�=oW��!�2���by��pn�pI5N/;.%��+��#H���N��DD4!�l�n�WQ�QM�h�*͠�����(~�W�����D�c�]���n���ѓ��e�fh���9r��h�g.��$է]�,n�;�Fװ�������j�[���3��<�<�N�Â'5TG�ާ����Q"E���9 �S�3J�!�'�KT��f�5��x�S���������᮹�'m9$k�n�b�.݃�;;��q�#$=d���)Z����j�l���ѓ�B�ʼ��;��&��^ڲ~��e �������OQ��g�L�)3"�ʻ�Q����[u�2RX,bG������6��G���؉�����*4���}'�Bb�֧U'b���H8,j�.+�۟���+�rw�l�ݝ��D�a�y�v(�r�$M;;�j����䘒A���f��
ٸ�X��x����Q�6�f�,f�+�LS����ŷɟ���5I�1�O5�9g�;%���k���[�\9���ݮ���T���j�pEoa޼��xQc�|hk�<|;;w74���*�W A)ÐA�ɪ�u��|���Aϵ?��z���5E�9�A�$�8�nB��h<��l���=8�>���ͱHtOJ�0A�$�@B���cUZ�����W���%F��^�9�/
�_�{� �y���>յ�^�/�r�hv�@���*=���;5���V<b.��4|@pi�Y;*p�W� ��R�k�?gV^�]"��^uJ�	�N��8&��m�9V����0$�,�qA>�2��9Ǘ>E�S�6��y���A'�&�Lm��(�����s�Y��/7(��ʨkE��VD@���{�4�iZ���I^=��3��u��X�޳�CË�֚���#a�l��{��ʴ��7���b�/uq�`�[��W,�a��`�/�eg���Q^��ĕ���Ic�z��&�t���%C+V���\��2��a�2k��v�a+�u9���σ��K�hwN.n����Z�L��Yom��oP�D��.=2�`�������%(n��wvByJ4B�W��n���y�v��j�JZ�R�vw Ǜ�Pa)}9���y����^KO-w�]W����1�g�����$)�}����5:�ݣ�L�6ۊ�����D�;D	����+���t+vn(��C�zN�yT�٭^Σߴ��'�v��'g��V���K�E[�n�w�^nQ��|�/hPf���ȓ�F�U���	����C��D.�䳩"H���躏rn�g�s��TGP�/�w���䳧g@��5�TjKu�9�Z���Ͱ�u.k���A#H�o)3g	�A{`&�t�@4�t����N�y�2�n�+�m�Du��-t�}�YQ��+��a�g
�n�O��1�.[{F����dv�{�'n���O&d�s:�.�V�ז}O�2��_Ulc��O�=�Ao���)|��� ��!������=�����T�����nc>��aٸ�t+�����.��Z]{u�|����%t��:�g�ɏ-�/���_~����J�>y�i�� '�>�5���^��-=tl[���#O>�q����Ǐ<z�Ρ����X��k����Uj���BE#m��8��׏<x�|�7ͿK�*~n��m����*,��m7m6�8�㷯<x��ס�9��zwi+]-�E��X(5H���q�x��׏<x��������ص�mI�U�Q�~�(����1����[Ƀr�Z��Ž��'u���\�\�,x���rܢ�;����:�lcF�o�W�\�sC7++���+z�x�m��睢�����.Vﮪwv'Ko���k/`�h�����>��<Z5�Z5U��Sihعu���4p�X��*��������3P�u�!�s�-���L��M��0s�F]�uN�"1��ٙLS:��$��՟�Yg�\L`��B�͝� ��V�� 9K�]KB07ZF�0�n2XqM\�j*�`:��t{)et�؃�i�.�5��M�mc��X��Ʋ�ٍ*ҵ.f"̻h���u
Y�\�f�V[b�fr�(�E�\ku���Te��P�r�]��a�ֵ��+�dJ1��L�5�v^.���\�ڂ��m�u�\��D�0����3f���j�c�^��5I5ƶ"0	���f�P�.�l�elчMX��U@#�)M4���mR��%6��a�噩3�c�q+M[���8"	.�U�F筱n9ׯ����$�-+��� df�(��&�)r���\%�i�Mm-�����MpP� �)a��i\e�lx8\��6�fiA��ҮٳX�mi��n#�!-qġ��^�4�Z��F=�´k�h¶j��a�\͵�4aU��j�ˠ,5�"[�G:T�4J���$ɠ�-@�d%�F��jDM�ں��YaJ[Ѹ,`��Q����|�'���H���e�G�-�R�۲���[�,�Gb������^��2�[�]�&A�0�SK����Ͷdcf��j0����ДK� j�E%u-�jmun�m4"�*è�X�ػX
v	cu�`6��2����ѥ�;.��6�e%��h��h�j�(5f�l�f�zj8�*��Vk0hW
K��L�b��0���5��4Gk-&,)��Ks�Bc\Z�T��m�#��[BYp�e,�(��f���i��p�i���	B�8bK��1k,e�K���H]��WY��[�L��嶱ai.������&��B�l�&M�k66Ű��A�z�<_5��`�7�4������Y��&\3Ycf%�䌳e�����%p�#�i�b�aPdd�����Ͻ:��.���(Bx(�%����6���0�BlKJ*�R�B��F�(�洗�]��қk�܌K0�	�5W:�b$��uf�� 8l��i��1��QA�+cal�����uF�3U�f���!T+d��q���������2�˭j��L��的�.th�͐ �5ُb�X}Թ�o{������[{BLf�,�W`���:;�k��X�)�d�K��ѥԲ��֡���I�N��1�NI�84h��;������^.e<<�=�S��u���.�T��&�Ò�N����:�3��M��݈f�߇v�! �'���Ț۝��.�R������Z9�����3���Pr*���N`��滀.e؛�2�����ʡ��x�t��ʼ����RpAu�^-T��N����yȳOH9<�؊��U@������ޅ�����-���7�����jx7Qa�����q�8,	�N&�9I�5��bI �O��7~���2����q�@8�p*���MS�����>O���/b�o��� _�e�Dz����Ƹ��3,˱��+-N�( D@�:D1e�S� ����+8"���X�/1��ɼ�R��V�w�t�����)�|�G ��bvj��i��_�~�N��I:o����le�M�D݄����j��f$}c�|E����d�!}Ϩ�d����v����R鎇����{�x]�]������j���aG�>b7�x�Ll�oN�{�����Ëˇ���� 1\հ�7T_�{2��Z�䳲�PA9a3��ta j��er�A�,ʐ��-�:g3�s���L�2[q�uð yQ�E'�HU;��Sֹ�?^a�e �W'��B�.�2�qJ�Z�˼��NX�Jo=A��|1��65��b;I�5I�$��E�1�M�p׈���j���<�����ћ���9�|�p|��'v"��;T�]�k�s��fETriK�.�$�����Xa�I�&L�15�1�(&�)6���� C�͉� �4�c ���c���𻜛�AݮYO��6�1$�Z|KR0��ד>��M�,�c�v)�Z`�7n����Y�A�6�\�r�� `���E�� @��̽�+�j�.�1��]��XŮ�'�Kܺ�H+�{W��2
��")8j�ES��u�������the�&�_Q��y�1+����p�S�yaɵb��=6�˅����z(j��t1�n�dX�w��Y]�����
���o=װ��$<����RS(�LƉ$XHA�1�g�{�t����k^{��s|���A�i��AEC�	h��@*��P��"3_�7N�u7� n��5E�������7²s�_dCO#b� 4��Q�j���[V'�O�T�8 ��CUD@"�C�ڨ��N���rg��hl��V�W�we� ��:��SB$*@n��c�뤁���~�����ff��ei	[)]R:�n����Rͦ�(D�t���@3i����H5JS�k�u�h�N���}��T����<Xg��8v�HxE�b2�;T\���pA$U;���~.�ry����C��P`=��r���um�s�4�&�N&M�bpX���\�����6�N�� ��v`�T���w�R�:!I���ۣd�Z�ʼ�Ų�yd�#�x4 &��	�O����������g��A� :ט��I�ْ��9'y����o���'ΐ��#��޽�� ��tN�x�SY�ٓs�PV+k;eC��e����G�]�!�R�d�f�8��Ej���Z�����:�=�"�a��̐	�L �LSi�&p{�v5H3��w.�#T��5K�|�=�m<��X�;��]�[�ͳ¯���v�6r�X����r	5HzDEY�%��2}gwr�^
B�f�a��΄m���T��n��"�(L���ݤ���}�'�ۀX_8v"�݉�NKefV�n�*�z�8݉��jTd�90,��4��N�T�����'2 nS�f�8��ڍ�y櫆ss��'ح��OP�J�T0f�'��bP� ��؅v�]�A�\=�UN�� �D��F9wʕ�;��p��A��C�8,�X�(�r@vH\
une׎�'&��~p䃶�ش*�"����4K��Ǭ���Ł9iȪ��7r.cYƂw�$�V����v�ߐr]�r*�`��|��Teމ�e�vE��R�S�;�R��sɶ�1�.�8$�v�0�Y8�u���S���5�������w\nNzjY��f��#OL���۸�j�r����������?��^ޙI�Y^�Z*�L���/[߳~_g|�����>_�ʺb� ����$t(*ll����r��-�1
�E��P������U@�� 3j�
n�i��%�
��:��"�lH��i�f�e��ξW�([0ְ�J�X��l`�m�e��&m���x�oܒ�Xi�Yl��.�٦Zh�Z4��l&LUх�lQ쵛�q�iMZ"
JiV�F�	�߯ϱ���5�ϵV�S�D{ע톪���s	Y�.���gV�
kV�J�%���z�6�̮��<������t~{��5I��xO�g"ʜ�ʇ����n��*6��rl��J�
�+���P���)y�塜�&�ss�z�� ��g�7�C���jwD���Ǭ�׎���	�
�<��+�⮽��=᱂��N�l��4��F��T��V`��N��%[�7~s�]�e�"H6`��a�RC���{�,���kl<�r,�k��	�O��|ħ���#p�X�i^wDOQүм�;mNh�K�F��]˂l�pA�p���^�s�b, 99��w�)9�y���A9I��>5I� ���y�n�7zլ�9*�;��u���ogM0�l5[�J��ke4�VoE>�w��!�U�$��h�pA�qY�ս9>3��:��5�*�;g'�UT��9�f�,��Q,|X{�;A��b$s����w���������x�܈��a_��*�Vim�(X�2+��t�雘U�Κ�bi��%��8ovbS�z�K�a����hϮ�C�
]%��[u݅��
�s�1#	R��<�\�!7�h=�2_-)��{{�pÜ��S�[�f�W^~��X���p�N;��.�c]�"��˲	�[�ۦj�z6soΜ��?�6�v;��9@ZC���R�
Ѭ���دƪN5NB(T�*�뻶�O�5WÙM�@LI���.��8'Y;���cT��Ʃ8"��j�C;����_�$ ֚P=��\o�򬌁��y �qÐ9�Y�I7n g���ǜ�NG
B���kM
��XB�.%�fn�*��rJ�YQ����=���X�
c�Z쳳��Z��Mw{kw�p�7��T��w�x���u�����VC���� ݧ"͸^bݻ��/���>ۧ|�"O�Dj�}���s'ޚ��̫����<�U{�5^t�)l�	������S�iQRq@HrP�(P;`��{F������,O�	Kk�ߚ�h��A�|�4��Tu1�˱�J�Eu�t	;C�)[۠��S�d&`y�&5�HD�"L%z�C1��Ř!�,@���>��xGe��ڴ�pzPp n��,l�rA�A�5N��O���� ���4��Q՛����8�ȌΚ\A)9�/J����j�rA �'$�F�,�U ��j� V~����}��]�7T�����&�ʹ�$>.�:����@wd�!�Ū�޹�1�Z X���k���\V!qΠ��6W3���LG�:�jX�ק���kX�;�,��;��A5I��巢�]p�s�B(���w��+ =��p�t�v ���b�S���_F*ձo�4M�;�d@�ޚ��t���%�:iql�ձ;19�1=���m��}Z	�N$2v��	�UDh�zdT����4'��2�D�_e\�ŞuñNS-�Ϗ��I���=ѝ{I����;�MRq3{_���_��pÜc�����shuu�}����{�a}}xn�Q�XR�CT>���t�e�޾ݭWYW�.�J����Q���v��CU։�ʫ��1��}5����74C�T{�	F׃�.D���v����-�r�;&�{;�}����:���U �4�0`�7� �Ll䠄����Xn�U�a�t֒\��Ff��i�L�Q���?�y������8 ��g�w&{�4"&��s*CB�U��]�Q����n��J��*���v}ӯY$���<jv �we���_�����@���I	�@4h�!S��LfaÑX����ːj�9T� �����,yl�tWf.��|�|Ν@qc#I�x�5I�������'1܏C�e�x���d�bI�́ ߐv"�u���5WÙW�R'
�W�<���`D� ��+�����%��rہT��������1zU��]Ϲ�uu<3E����B-�Vϰ!�b�k�W]^�މ��T<�^~'G��K��oJ6�,oh�D���@���e�=Å��kN-bp=�̘�np�5����´��y _<��h��`�bM��*y�����}�ۊ�Z�:-����j����m[6��^ֲ�Ņq�jiL���%�Md4+Ha"4�&B͈&v�`�#�[Qsn�X���g@G`�,���B���3Fch Ĵ�.�2/b�M�IYn�r��al�r�6͊ܖ$p��".��l���j鱁��+0Ըż�Pw�z}x� F�A6���PB6��k?U��5.�
1[�4�:F�.-��A4R�a�q�A���=C�֛Ї1����H,*���3����˧̶޾Nm�>ޓ��Z� ���@�Ʃ3ҧj�q,���ў��%͝<�Eۇu���4#�WÙ_;a�v"uU�J9����t�����q��ux[�ŌQ��U&�]ӈ�z�.N\�G�7w^ќ,�&�A��ÃF�=S�"�Î�M}��3�x�v!5ˈ$�;KC&��;V�Wvr�x/�o��\�Ł9I�Y	���׮��(�i\���,}��ոT�}�B7,���~�<���\8��f^״P�U�g�v���ę����*#s��sp��]��Nf��k)�e����h	�T%%u�k�ي3�d5�8$�TBge4S�L��]�f�#|*��4Y�u{v}��쮜�lZ��*�.7nW�$��r+�&�wfp~��1��T��y��5ػl����ZY��6r+��E��_���̌���!8Z���u�	KWJ�I.%�qM�@,@,@,@�����t^�_�9.q*�2GV��;n�Z���#�y��V��h,}	�e�6���A�eT��>���XU�|3~�������Y�pM�"u���pM!�����t�r��]��d�_����t��+����Wu�p�af��C�U^����3��:\k\9Nh�pER�U����q�;T�5�&]�ʯf��f>f���v��AM.�hR�cT��*��8�y���8t����tB6U���r���)�ս*J��$����� �� �&]�l`y�@l8v4B�UNeEn\��]����3���{�D�=w�kFyÑ�L�2��e�y����i�y�ѢX٧N�;�y�1����̧�,�-���/1p����HׅSH;�K�K��g
�'"��N	)��1Z@��}�r�#s2�cs�8Z+���j���#&�%Qٔ//f\�q�5�����#5,;��X����ǵi�= ��趩I�s�<D��ۻݮ��lV\���O���k^ZyP�6�6n������/2�a���'k��U��y��Jw]��:��:�l�+��Y� �B"t��K/V�btT����3j
��Q��%�Z�vP�z���]��t�=���]�ά|��ۭc��,U훶u�\�(��xǄW�;��ш��6_e]Y����v��.�
�5K�QV�<�Vɷ@�.��nu&{ݛ���;�5�)M@�j����'N�ju�8��^>Ք�u��֥[��e�:��9�XY�ӻ띹V���[��r�q	�jo^n^,/����x�uz�[Z	�Χ�{op佖b��.Ww��=	y�I��fM.��ܢ�BZ�;mJ�-���L�Mzo�
U˽7[;���KήW���53�aqy�>�}��n�֝��y}o��������V)��0^����s�/�:5���E&p���,�v��U|�gZ}R��L��Zl� �z�b���O������'�n�_ۅiA���ڽ&��/`�gק���:��[��Z��d��v�&w$���U�#����z��x���`(�a��9*��wC�ֶmؚH���;�[u	Y��Ɔc�}��M4R\i-F��N�R9al�)�Ŕr��HUkt�(��H�%���ҳk}o�%���yf��(S̥�����U�k��&�;��Vau�w]�!�h}8�V���Xc �j�I�cd���	@���^"lT�+C�;8{�U�]�/�C���ܵ�Ā4	9L�7EdI#��<x�׏=x��Ǐ^�t{�M@�jj��B�"��O[m��x��׏<x��y�55��$�|��"T�-=t��8���o^<x��נH�ؽ�+���\I���n8�<v��Ǐ�z$��sh�>UJ�x��m\+�׊�ol[�wk��������$�҇t���aK��]�\�m�^w�S����w67�Ti$������aW.F��]ߞ[sƹs��ۡ^wLܝ�1nW5rKEuꪤ���1�P��TU{Z��7܌Na�-����C��!��gc�N��T���B������w����2��!.WE�\�O]����8�6C�@����
�}��@�C�mg{�v�#6�E�@�*���7��s�o�s}����g� ��; ���@(B>��� ^{��2y�z�-�a�V1�]vѺ7�ۚFVk
U�~��/�!0�-���w���p�z��X��)�ܭ�A��-�;ژϯv�BջK��;[����})ݐ��2�����[:s��{۱�ǈLy�V��|��{EN�]X���8v�d ErG���#cG�#g�k9I{L�w�8��3*  ��Jw��p���A<��$�����5��s2��0��-4�̖DˇL�po��%�^MC�_�v���u�n����3.3$t�� ��M��,r���>�ܨ�DK�g�#TsнB��t��ei7�.�ť���yu=��a��m��F�+:�;���+�G�y=�H�+D��bF`j�	�V�'Ԝ%	�A���0 "�W�ℏO�?ln��*t��̬�h��'\8z]؉M�B�Ｄ���h�*�2�(��Y�v^��䊩.��ͅ3.v*�XTi�6���_�}��"� �R�30���y�x+�˼�<G��/w��=���L��8�	��R�c8U! D��ty��=+�,�Z�enf�?.��q�����ǩ8!Rgc2�:�����v� ��<K J �2s,PR��2B�!2�L��0��7�.�}W�O�T�5Ջ�_8&���P�R�f*�(s��`��V��ɛ1h4� U'�����\�e�z�< � ��qV}a���l��4�I�['cj�l�H ���}Z!��{��-b%H�����p��ٗ�:wY�!ճ���	��vsT�U~��Xb5V���>�+�>[���Y��oe�wX��:̜-T̽F�6��MY3���x2�-���8U�S���Kq��<f(��"%�;�nbň�?�x}W�GP�A*T���wN�"�@��Xj�F�ƻ��y���Ds�5̰���4�uW[nw7R��x�&x�3�j"6�Mssq��u�;�8���iU�,e���:n]tu7;�v��F��n��\��[m�#�����գ2E�1m�H����x*�	4ܻY�Z9��Lk��U��h�WB&+�vԵ�^�J�g���i��/Hŕ�-��m�
��9�xr������Z�d@�3l��-��kj�Q���G@g�����:�AoK�H(V��u{N�=���Е3�w�)�1 xFc�b 
vv2���3)�'��x���U���N�q}�5��+]�w�ᇁ���&�s$dW=���v+G �Ñ<��S"Y�BHA��p�[����j/v|98��w0��ˌ�;ڸ[ �Zp4���ݦsT�%"���'����bi:B��uoS�������Ӟ��SF;!�b����3)� ̧ �L��UG�Vv�l�/��Cl��^i/o}�y0�#<�DӇ�L��{񓾍&���=����[�B�s��B�92���+ZK+����81�f_�;���E�
�e4�$�����p��ˌ���;v�ξ,vZMS vS�X���9r����v�w��J���g�ގ1e�|��ॹ�*G�����$���f5~Y�'m޽�Q=�+0��a����T��bF`��p|B#i�����p1�KZ��q���8@ֻ"+FT���٩����ji-e8 ��9���z�oY���~x�dy ոp��D1H	�`��#�k(�/!�`�x����S!�ۻ}�x�g�3�ѫ���������������f�%u^����-��a�ChxV=��7���`�zm�9�}^�c��`"3�l���p����)�a{p�S �����T�<� ���:w,m��[u�6ee�Uc��xxr!�7O-~���I��'ו���l��f? �"[��7Mx8�t�J�HD�`�Dˇ�IG5��v���"�D~L�+����C�*s=���zS� ��vvN�.��!V'*��Et�YDf�2�&�( �Cˊ�;� ��Qݑ�'��õ�y�{�n�֠��
��4�.UͱF3TM�+i�Ϋ5�|t]�+�f.���7/�ݻ��+�iu�> �]���5#'�Hq!�O�_�]���o��~o�wr����{��Y* �qU;;Id%������Η^��X��ɵ2c:��,��>��u�j���� ���8��pJ�z �c�)B���wC°CZ�U#��`��q��&�z�L�1�W	�N!�I	�)��bU�����1�M���M8N��9J�QX9wV���0��Gib�[�*�L%K;�y����z$EyÃ�('y�\F���]�u�������zF����#$m �V�v ��ex�NEk����oj^�ص�b��O� ��=�8Y���~m#�BO�)�9^��h����O���9n0�(9.����������{nv�ќ���΍M�zS�H��A��r	�NIa)��*m�'R��A،�IdD�!K���Wq�~sq�y��8"�F1�z��`<v�(�DD�Y&���XS�N�t�#0n�5�y��j�ñJ�*yYF��u�V`�k,��6�)��^y̿u���!P�'!����h��0#0#�t��2v�oup�7�pA4B3++k(��M�{"[B5���3Z������Y����<��d*p�D�"e�q��׹�X�1�O���kp`:vv:E�\4��eE�]rv���ݳA��ﾽ{���g�Bs�"e$E�����9�{-�G{W7�|c��M���9a,yRZ� MR��u5z�uM��6�`�+�=Vz�]ﺽ��=�t�YD�e��K���&�Ag5��a� ��CG��o$�]���D��P����|��q�B]��X#
<�V8r.�8�o��bm��x�����m��E�pd�����#=��w����'b!x�Ϋ�*�����ѷNA��š	�A���Aȓ�2��E�`�~c�}�/s�^�{�<�|i�(�'�8"e݋"���P��y�����4��t)����ʹ+GU��i@�ƕ*y�Y�'�{U��;3"�	�l_Ǚ�̧+S������G��^�.{���Z5,��/�1�Fg��/0�V����UN�-�\���ND��u,l�a�f�\�&��Չ��o&��!Ea��ّ�c��v��-���#]�,���i��=��yZ1Pa��,��+G:RMb�2�fs�l�4K[4X3j`.��8f+��Z�6]D��R�Kh^&�;5I�䦯d-��(�v�.vQG<#H��K��.�k��p�4�f�ݕ�_��{�?<��i^��ٓݬ����(��	qhD��v�A�Z��MIZ��*�V�ś�W���_�Xާ#��� �R��gEw.{2�5��
l�Ng�V
�t�tO�ҁU8pDˇ%��
��̙+4��"�8:B��ܽU�h��س�� ��|���QrMR�,��P��{r�Y�3҉3��.�l=����c��Q�RJpS������Tx���A�`�������i�K9�Ή�O��2�Y�9̧i���vr"��)�y
�8��&ӛ��F��`�(EӇ"eÁ$���%��pELG�u	z���
��[�h��س:1q�&t�Hs2�pZev*S�F/�D�ߞ�.u�Z"���0�I�r��--�Ҷj&�� %� ��Z̵�� ������5HF�{[�N��=�eU�j���]�=���ر�vS*,�9���z=s���=�n!/Ѣ�;:����w��n��c}a�y���=6/?K`�=��x�༥�ה)Ҩ5��� � l��
�Dۘ�bŋ&j�Aԥ��N��[�Sٗ�C[y^pA�p��[֟8)��U�����ػ��҈>����)�Dk؟W�;�ϏQI�w���V�!�b��1|����d��BX�)�2j"�����xgB����Y4Ç]�0��vk�
���	[F9�[����ƀ!�:BʒqL�RpX$�KL���1G`,)���Ot�fu�U=yy��7B� D�3.7���߿�������(
iU�k�%�e�]]���V�*-M(F�)�&�a�7o8$I�t�q�z�;DMf���B/�ř�����f��ʭ�ōՊH ̀�҂��&n�:*u�C�F_��v{�}�)n%�/���(�8PT�"+9� ݷeyb�HNX�r5���&pj�d67=Z�ozgn�=^��b��zc�̰j�mwlYr!x���Wh�|�W�6>�1�NϷ��w���i�	;���Ç�5UmBJO�$c�>��o'޺ǲ�v�2,ko �/d�p �(f\8�@�#pXVsA�p�݀�@4BU�G�{��c�s�?	�4���쪿N9`��ih8#M ��H8 �UE�LE�Qv�r��!�8{���Q�)g#�s��}���`q�V�r/Qb0vzITb��jFx :2��.4r�����M�,�F�)��eT�b����>��?��؝�2Ȑ����2�r3+WZU=w��FWl�Kozi�-1Â0��*����v�U�o{��h��vqLQ�Mz��f�!~����J�-$"��>�w�-w6<g	��$<ˇId!�`m����:��w�TfN��;�d>�$���L�ؙ!2���N]º~���t�@�&s2�N��_.6�z�2sa��e["bn_��~"�Y��W�:��+K�r�����M`��:�ҝ�ߛ�xM�U�*�:c�ە,c.�D���9��7��C=�������]s��C����4��u�C�Ie×c30�J�	>��[Y��
6�ywwby��A�NA�TD���x�^F���NՔy�=B&]{	��4����cI	]))��i�:�2��m�Lr_^�������@=�Id�.s=t��I��=�d>pp�:��%��6(FӇ#e�9-$#2��̦��1��&�@iLQ�N';��OU]w�$����A�#1���'y�]�=�-���pA�J2��.���4�����ƉiA ��[ʷ/x{ȼ�����,���NƀL�<�]~M�T&�%ut)�B����˹���%f�-[����"����ȠEӳ�cd[*�z�L��i�c�ѽ�X��X������6���25�� � �E�L2�#�RuX���]Mx����Y��U�'�]t���U�$OJ壝��yÕ�ڻ�ٜ;��7[%ѩ%3T�V�h����̯��ϊ�LXnaF�ə�O�[�}we�T=��<�i��xh�ľ��شTb�s�B�Q��v�����tgW���	gE��{أKwL�K�{v��3��m�OcY3m[���{���� ��թL���l�,ᜭ�Ū�����;sh˧�+
p�b��n��|#���qi�+�nU�6\�����ڶ�Jb��JcU�k�[�9���*j5:�Q֠4GS�s������c�xwl_-�R�f.	�l��We J��d�����kk���S&V	��G�N:�BS;�j�Lc�le������bn��t��
v^8��:U�7��ۄ�Ç��:v��l�ְp���yeu���UC�/�p�;H�Z�;�,���m<G���t���%+%i�wS�7;8���s/��{B��}5�k-�)rʔ;��t_���MCd�L��눺4�+n)x���9:%$2�w(si��)�gk���\�o`�1H�l�]�+�!ưP���z�J]���]�x4�����W�0�j���j�9�gu���w�!�6�7�;�ٵv��}���m��|zd/4F�T6����([�0ξYڠ�n�oQ,����\�ecK �֭�@�6EBd&[�[3wvC���B���Z�Z�%�ut<]�m��u�z�(�6=Dx���h�>�<�<�|��l��*ˈ.�TmX��[@�n���
T�� �Q��,U��V�%�k�P	�]><}q�Ǐ�O<x���_�Y�`-��hώ,D��
��P!�=m�q�Ǐ�x��ס���UjT�@�*wE0�ք�$z)�.'��&8��# S��q�x��ǯ<x��7���c^+�]9q�@Q�$Cb�����ێ8�Ǐ;z��ǯ^��E�
cE�9�J"7�t�(��p�Ecb�r� ���<v�	�v�%��u��Dd�.b�]�Xۤ�Id�.&#]��ͻ�5�bH�fc��
LE#-����J����N�J4�@�I1a"@�]���F��t&�.Q�\�[�������\�ɾ��^u�nWc��u/�\4ۦ4j41~O�(�,	e3	v����jJ;�n�vתƶXq 	�.��0bq����clH1�nCj����{W�;�aS=�PBf!v�6WE�l�G�/�4�X�j���K	k��i���ja�(:���,lЕ�6*�(V�qa4+N�vĺKERLG��`����5��Z��)y�b��L�M�n%�\V57�|���t�V�.ڣ`��L��j���3e�f��3X&���jJ֒���%u����f���1�l-�ګ�%�V�!9�Yą����b��c�K�bѠ�LK��$!0�u�[���]��T�r�c%)�e�-W)m5�F�e���hG�i��y)�Q��q��`�X�R+ʇiu��;.	���m���l��lݫ(�F#�a��[j9�]afe�)����0�Y����5[yn�����T�e�0�5�jM�LS����CK� XSB�g� M
J�[+CC�P����LM��&��b�Db3Wa\C2�=k�,ZҎ�V� d6\m5��ʊ��<��V�K��4hJ�uukI��f�0dIZC:��L�\��4�h�K��b�J�8
��ktŦ��&�l]R�� i`�ػ+/j,�f��/�	�M����)<|�0�Y��t���M����Ii����\Bi�Uƨ�2ɑ�{GGE��4�j�&l�3n�E*Zـ0ٍ�lrՕ%������V��(
����q��q�#f�a���BL-��gM�%�j���oZqJ�h̒��( �;*�4�\�h&�%9��+e�0�k���M���e�Z��CkV*��u��Y��.�ev�5�\���R�eVlDu��]��kl#lU�a�h[���7�1���$"���0�ˣ���ֻm�Ú�R^�!��e��q�gu`ځv�n�Z��0׎qn(TZRŶk*�ɚ=��b���&j�1 �bŋC$Lo��4�5��� ��P���f�H䘠7[4cL���W��؍r�Z���vXiF9Ku�k@�Gr��Xm�LT�]���u�Dz�qI]����L��kE�5(�`4j��p��&����Δ��Ky+��*R��L��A�.��2ٲ\9���4��Y[.v��ZZ۰��R�َ��V�.�NEefe�f
5�k�;9ژ�M�\��v��w���f�Ł@����&���`��Y�2L'1aB.��VK���^����>�}:bz����c+sܻ6�9�����.biS;��q�Z�é�k"B7�؂�r�B3+�`��\�Hx�r6ex�[�5�uA>䕜��8�(���`�L�m�˱�y�K��b׈ �'vA d�fS�2c*���Z�Y�s� ��L�6�r�29����y����AK�L�q�%׽;+4�Fk��HS@�Sw1���yҋ�^7F ;i��*.�NyE���s!�s$9�/K��Г2�1?[�X̧��!=�z���'���o#�v���߾石��Pns�B�C��ʚip�9���9�\��0�����K���9�N|�i��Xܧ[���<���3�p��.pm���m<'��A�\�r4���R�;���Ej4��	I�'��/F~��)�G��8a��0h�-�~��%w�ufY8}umc#h��vl��M�4r˽�uʌ�B��s˺�.�߼<�bŋ+q�E;;h�=����Z;�z�ם�N�pC��&��]{�ç�g<z�G1�'k�Iv�	��."�ÀD�Ai�aσ�>�tHO;%^?9��W��"� ���&\;��̦d_v����L��F�9i�7���xɪ��־d	�@ny BYq�Vu�aC)�r[̄�pt�	�
���>OE5�:B�W�Z;�\�:1s3��!2�L�ё��U��ki�[���u�3
�u� *��G��
�3�bH;@VO�����A؉ "�Ŏ|��s!=`����v�f�zm_Q�9.꘣���C�=!���M���DZ>^2��{պ�j�U^e�Yvc�r$��׽"�B�8ql�L3�CL��DK�d�a������ ����u�y�i��(�/�,c쿬���w�#��=�c����9��Q���
�3.n���2���3���P����"?_��m���k,�*~����nbŋ,[�!����s~��ҕ�{2�{�1@t����PA3*�W�����j��&�p,;��؎,�\8�5�E>d�˹��Y1�	Qwrwd���sS�v:Ze�RAc$&�2��A�i+��ƸW�#׽��"*�3��Z���X�v�dS��j>y1�0��'���y<���h8]P�#��`Jjh�p��aJ��x�_RXJm| ���٥��=��
�o62�O����=)^W�,t��*����/;���b�B �� ��@8���-4�1��kf;4�C�d(�Z�����*~�(�[n�E��=��)��<��T#��gj�v"�pfP1@�TMd���/�\_��YY���&�35��'!	׎%�P��B�ðݝ�����l���9e���cD!����ʭ���ْ:qq��NX,���9�(R��;e���biܖr_I;1�I��3%�>�sn��%?��-ٻqAT�	��e��[��a�i�[s,C,[��&�N�[ �T�ƥbv ̸v"MU�n/�s �EÍhcURld�;ǖۅ|
,�Zz� �:gc@��F�ױv	6BE"�#�=��g�T�ͷ]&��Ă+��yo0�4\mf(z���w\���NXE�T�L��ٛ��Y���̅�NI�\|��B�#�Y��8E�	���"�@pA[��J��M�X�E�D1b�C'����Ep���g{�'C-.�5����X��;'�x A�@?�K�b$��q��h-$�_|�l�����pY@�� �@I��2���y����=z�FT�S.!��' �2��:f�{�d=Vfg6p����;�=�(����>��%��"J2��3�>j�u����2���_
{�e��7t�8y$;���X�~�ߧٟ	@��λ/U�ڐ�=��x[yf�n���'�dS��GJ��=0b��'y!���K&b;'���}~O���hj|%���e�[L�0�ŋ,X�ݘ��|�(��	_�=�Ǜ	�����&�3�Ulz��kR���fT�
����Ȯ����h�hCr�h�ue�M�-��`u�#iz�i�p;�%�F�r�D�u�TbE���`ȷ6��f4��J�h��"F�XE�<�K��,fpYL�a�%��K0ݗ`
��`4fiq�1K/0,0B�2ْd����2�eIi�̪��)������={�$3���6���
)��S�&�`R�G��-���%�8B:�n3�X�$��;��XC�՘��vLd�(;z��k�����u��<�{����#$�g�p���v&H�I��e5�����-�^��Z�z�o7�#!�39��[@p@�NL2�9jj��+���V�_�c�F�E�S�5!׉%��#8Ȧ��T��o^�\�\%�X�m�x#�l��Z�0����CoˤT��C|�8#9���e�q:��'�r�qi7�!��I|���}������g]�p�Y>&@�'TS�%��Z��9��j��Y���猅Wy��ĞrpA� Dˌ�����<ݶak��t��" ��v�x�jգ]Q�-ͮ)ᜐ�N�@�:B ���b�3���UM��_�7�euj�'�͋���ԛ=	�#i�eSW���]�-ن+ּ$`7��sN_9�pѪJ��V ��ڻ6M�W�@h�O�U��ɷO6�[bN|����5F��ENF71`X�bŋ�b��z���9	VI��9N��*P�)�����;aYHL���5T
�9ʦx{��Q�w�︪n�.������U�W�l�w��Vd{��f�
�c3�;oc7�ߣ���Nkp�,����Ͻo����Z‪�3+w5�ׯ^ڍ�!�}�	U���/�@�R���|����
m���n��"��AC��P�݈)�
Ie��3-�Tm���ZV��\<:
��A9X�5�a̺��SZ��z�n�*��`,��Y~xbZ�oje;L�y���;��s"���θ���ݖ��{.�[ևJ>l@:��l�-�_"����"�CK��u�6�T���`�%:Nbc�nZ�Y�jk΋��F�з��D�w�^��z*k�P"�VR�����,X�bſ��% S��&#�d���v/�=,޳wp�f ��;����T��m��>�9����_��3ݜ2q�6��V���Ԅ�j5UQ-D�GC��0��f6��z��e�{�ˬ�i�g�g��KCǅ�ˍċX�������%\Y�UD�eUi)F�ٗC� ]�/6m�����p:�9=�eyCʫ���-�xε��n+�/�l�������H`i[޿v�$=�u����E{&��kG���
|�l��qS�Y���<$�������ymt�)��C<�8���Ц��~��Q&���3��s�=��Q78������{.s}j[���imkݽp��H����m�?X
��TfA��'x�Y_ky]l�ٿ~���z@k�Wh���c����/o4��?D!Y�b���`��FĖ���{-^[av�4�]�Փ.Besw���T�<�jU��LHB�uq>׵��C,X�b�`t3Zٝj�k5`]鼸{�k���M�g׏f��{j�/ݜBn��i�q&���=n'��6	���eu��Gh�hl�U�l�@u��)��)w_#}w���>���[�St�.c�V����3'6��>8a��T� ��fh�~ݞ�߷GJ�iTnA�g��6���鞽ؾѵ�FI���f�UJe0��c��+fj��\�\o/C��NT�_�vso�d�r�ϛҙ�f��7��n�,i�(L�����e��̜�.�l�={���b2�	��(L�A��s���z+�F�3xM������&G��O8����EZ�$J����썋"�zf���.���������񙦰շ����_I-:���=΍sR;���m-������AM��dŁbŽ;
n�c�P��I��l;���EB(E<��v�u7���b�+��Zjfi�s�����j����bKY� ��mK�[]F\KH͂��B�9�fu��wk��a̺.�f[eo*���R��IoV8nH���I���1t�%l^�Vݑ�e+L�iI���b-���`�h�.��÷2�G�Yh�BPd�7ݑ��K�*�#:�Aw�bv���4�����������R�j�U��-��M#��A��&B��f�]�$��^����4S��C@�Z�=��bv��~�Q+��)�4`8T� �[����v�!4�ʏV�Q�Ͼƭ�}@t��㲎�S�3پ��ܔ�1
"��]�ҺCSFb�`L�gmA�E���
ުܐ���&�s=�Cڄ�3��h���"�g��^d ���\_}ѳQ�s��a(�xʰ�[���I�\&��CKK:��tg���ӪlVF���輣ÔVA���hVi��
�L�����Nu�\tGO~|),ܕ������Ha�׮5���l�5f4.�H<!у�V�y��u+nX��f��8�~����/8�������Mכ%\�2�65��s1��'ԗ\|�����X�3��[�U>��ׯX�Vs0/����uqP��礮���ʝs��ٯF�f�P�O^yh��>�9��2bť�V��'���{�f��s��	�� �UF%fv��2�M;~cځik�w4�`�.�Y���fxX�p�#;ֺm���I2��W:�O�ȵ]}������[ն�wyָzHO���7��۞>�� ��[_! J2��������0T��Y���}�^NOg0�@WH�����Q�m�ߩo{��9�o�m�����<@uE�8�᮫�\��9<��ӘՋ4�M��C�XU[;e߱�պ;��X����=yV���7j�q2�g�dNA*�M�ۘ�ůw�����G3�,{�Ӫg�iȃJ*���w����	l�c��^٩��B�@?~I3�-Z��y[e�{Oh/����r.����.�Iţ&w6ǇQ��M'ݿK��ܧw��̺陈���IԢ옷���TuotwU��K�5��i��t=����r6yYܾ6�%0Q��3_m��5�ͨ����7D�J�T�8��u�׋��_b�����u���g���4-��`��m��=��ݣ��)X}�Wu{R�\�BVӵ��<�ߍi�*�wԯ�dt{j��o��'`�0;�쮱��owLu�3�@��R��:H�,�J�ލ�{���+����6*�*!�;am�H�OTk���.\��,�a@NGÛY���^��,�wR=N1#��V��A>Z(�d-�5v�+mڶ�ܩ�G7z�J��QO-��4���km���g���������B��^�?e��U;S� �j���k��H��|dST�.s��Ұvd��F������y�\�[G�7{�Wf�o!C.,)԰�����.)��k��k�R�Ց�9���-��W+�����^k|6�Y�Ϋ�U�Ԯ�Q7��v)d{�wXk�#N*�m]k�o�]8�/��][b��e��@���}�E�B��tz�U��4�ηkS��i�؃Dz�e�j�h�W�Y��F��v�t1�g���4�98qҤ���C� �ô/}̞s
��]zE.���
���C�^!ǦT�$�H�B��̱&���X��bɢ�
޼��+�1�ݗH��1ݏy�̧̭x��%j��4�Ạ,V<���՚�]v\��/M5P5"b���\� �D��%P�#	Q�2�:}m���x��<x���!� SIR��9cd�ahU$�H��D�N����x���o^<x���	���$$$$��9���!���!$�M=z���x���߽�~��~���|FF(�o��&Bt�t����D�� ���|�7���7�Ǐ<x��Ǐ^� @�$a�P�,��ƻ��!	-��HL�2d7��^�	77]�h	b
P"-|�P��<�di`e	��u�(�d��#!6P�}��Eι�"	A3I�{.��D�y�E�Q���v�d�I�L��BM	"f�li"1 �(��q��
$%�r���2��"�s1�4޻/<�.�ŋ|�1b�p�I����Ǟ߽������y7�L�4 %���Iy���C3�a�{jn_.poBw�5��¥x�s�kj�����^UxU �*e4ϲ��~�t�V3����Ļ���9�s��47�񢝅Tn����z��D"zRP��1V1I��eԗ"9�X�
P��G��;J�Y�ྷΞ{�x�{���߻�iB��e����=y4ñ:�]jL�Si��MU��H& U)���Z-��IT���N�����@�B��L�Y�
7`u����l�hkf=R���6b�g�y����S�y9�Vg��@L�82�d��->Pu�����qP��F�'��-��'���}���x�������Wv��?����Y�g�\�k�N��cm�ޅ�n���6���+b�XJ$��J�yJ\M�D�i|��,[�ɐL� ʾް��[��i��;��L�j7/�J�V}Ӻxy>a�|�S�q�	�KL�\.�<·u��(r�)��I��%�+`�,�հgB;��	Bp��[M�C)	��s�^UϞc�Q|�9~:e�;�m�L�o�Gq��J(L�2�n�k��+ء����Z;����o=~��n;Z�:P{k��e.��ݏT�P�1P<���N�Í#`.�'sZ�7gs���6��]K��2�r=�o���R����*]��HL�U��W>��=e�9f3��/ab����P�@n�ϘL&v��X*_&K��s�`\�{�Z2<6�������gn�P�w6"��f!躘�N�H�ŭ9���-����˲��ЇI�1fݮ'U��M��`���c��_g*�kU	U_ߍ4��MSM{�o��-����q���Qü�r!�*�$&�זiY��F6�[�э.�e6�]0��DQw\[��ƫ�k�!�F�ֆ�4˦�)C$Gm5`�.�M�ssA`����@�l��L�1f��f�m���HK��M��&��M�MG�l���ǚ�<�[��mvZ�%u�:�� ��.��#���o^�'������u�Q	���"{Hj����.����6�!�v��TX�D��!<	C�U��t���t�߿n�9�����w�-t��99�%�-��o4��yL�)�I�yi�Q4��rk���Y9u���
�p{�L����π�!--s�e �U &G��z����d����ᷗ7���Ҙ{P�C�D��P}�L�.T�o0=(�R���爗�nk	���,�0�N՚վaB�R�f|��zf�gk�ˬ���ëB�僘=�b)��X�9C�������"QN�d�����*Ŭav���l� ���vP�������'�^�gi�]z����o&�s�������h�gm���n�.ޟ	��,��>��*!��e��ٟ����z/���*�{j(//i��������f���\{%�y��S���ujn+���2dɐ	�&L�0dDǐ��*׽5�k>��W*�5����	�=��s�վ�R����4��0��*��(; �I{���xehU���h��� ���S(?9���J�:�m8Aږ�����x��w9��|�����+Z%�x�܄�2��WT�y���G3��_LX��Ws����橡��1��������e��U,rD.!҂�$��k��8]��ql�I������>�[�A�:i�3�z��O�"}����s�ޜ��JG^MZ�L&P�$��M����Ef�n�A��{2/*�`0ݼ0���3wt�)Y� �M�����阁 K��V�s��]�P���zt�b�Z �J5,fU��o����N?Y���G�^=K3�w��~��ۊ�5�f��;|5�bŋ,X�n79�7�U���|�Һfbei���Wg�0�Y�L�����>O�upS�����8~ά�U
<ts��D��t��2�	��i��S3�����&��Q��m+͙�uY���3�	���w�>qZ�c�<N2t)3hCK	�`a\;Yf�-V��.vػ ��s)?����?j�M��N}Ӑ����}S�}U�e<�M��'��;e�BC�,���e���ݲ�a��_{r*�v ]p�� ��"ó��yh
�,��/r�zK��l�7U���9�}�FU{kU��M��Vv�7��=(4�i�!����A}��2��1l���ݿ_�%]�a�2����^��Vr���pSk%�[h�K��.X�e��O���_���˂�V.���K��C�`t3���2»�E��ܹy�l٥K��B�e��
��Vy�8c��1�c8땯����{�'��f�ĭ�OùޟLM?� eƇ�3��-�q
���K�K�{�1�/u�w.V۵�檴�܅��GYG8	���E5����iY�6�聪�9(�gI���Z=�Q~˪���b���>-,{��~5p�f��~ʄ�����%��g�|C*�j��^�v]=�d0��&�n��0���uVy��W�x�v�g��>mŚ|�3����}��̫����Fs��f&PM2�@Qڌ��x����A�P�:�e��;����,q��*nAփ���Y�6^gĉ	�&lnK�"�{ҏf�����-��+/5�P�������BT
�%�U���ߗ��_��b�|�����!�E�O�����Է��v�唖�Diن�������� � (nbŋ,ZE�v*��n�Tm�.A��H�4���x�Q�qI��,��U���{��,�p��fЖ۳P�4�F�4�^/l���mP�S��UcRʚ�V���װ����6��4�0��Mr$�B6�cum̱k.F4��:�
����;\��c3uP�gKPlq��U�S1�q!L��!pBm&U�&C0��t\�ߟ~��?>yo����|�޼����T�Y]R#	���h��6]\�����.��8;�@�xN#���,��)�Vg\��y�[��o�]蛃}!�U)�3�a���g՚��ݠ�T���zw��VNp�|��l�*�y4�:M�8Z���������>nq�=���*� ��Q9�3������ޔX��A3�U^��p���wʹi�2��}�����vߜ��_�׫��ΰ�ˏύv\���;��h�]�:Nv��uƱ
�b�C�Ls�V{;;|��M3��Y�x9�ٔ�g��O���X$̴�j�怹�3[�4�-ej"��q3k�I�����g��+o�f+e��j�S�n��0�κ��xv�,��a3-& �$��_��%�^M?�|�
�M���;���>ϯ��|�݊��2�/e�R����|��/;�-�$��s��KB��E\ItInbŋ,Yܐ}<bj�Xf�<�f�;�v���1�f�·���u�� Ce�1UI�j����^xqMu�}��{�ŝ�7�	��I��������f{�{���!�껮�T��yy�$5w\k��kZ?c�5N�f�m��P�|�3uN;;�v{�1�A3�h�|�n|s:��Q�`P}?1c2��.��������&`�ݩV���:ļ�ֆ����}����(	�i���t��mb��}5)dN�=*��j�C�k2Op����9�Φ���EW���]���^{�<�fW#ni�sPU�%���1���R���د��瓿����h�̮�+��ȯ�kw�}z�^u�]t��
�p�4í�,����om����2_۹S�=����y\��m��,X�bҁ'��nlq����c8�TZg٘e;L���Z��m�&�q�+FV�u���,�<¼��r�g���3�!3V"�!�S�ˀ�'�Ϧ9�С�\z{2o��]�k�^i���5^�G��=���/�Cސ�z��=<d�8�a����ke�#`�����8o3D��Yhp����Q��UP�Ɲ�Qq���(˸��P޾0�g����e��Ni.V����7�Mi��ŵ���ŝ|���͵]>�N.����Z�X��L�&P�����nx��A�|̛�M�����=+�fL�j���+۹~���k%�=7½'Ӿآ��Ɗ?~u7s��O�*�����)���f*��y@]������ؼ�wY8R� ]�)q�IE����f�ʶ��S+P�:)Ss,X�b�=���e2�ʙ�cz<=J�a~St���c�x��2n�-�g��n٭�2W���5>���?H?��9�J'ZF��6�`��+��Vkr7I��Kc�H#��]3 L�ʯVgzo�N�[�ƕ��TA��_����Tٯ�%Ӣ�{U���v�'��-���:VM��R���(��h	�3ss����X&��_\᫐����%ZB9*��7�;ﵗ5�k��~�����[>���.�w �چ:�5Q]��6/ח��&Ɨ�lN!����`L�&SL��8<=���-..P�We+����{�{��N�3�y�!�չ���|�I�Ǔ �?�쓮�;U9�y��l{v�Lśt*A5-������nZ�Ջ�o`�z-e������A���a[T�Go���c�\����i�G�,���F�p�/x�U�wpvp���M�ܣz��=�r�neek�I7�o�fѬ�Q�������;�lK�q�!�5h����;�gw+�5N&���*�xYY�t�RۻtA�j���4nC�.���Z0�оk���{r�Ҵ=e^*�f�r�^�Oeo,;NU����;���.�&�t�JK�����G(� ֗
����8�Uݛ�d�WO��ז]J��_mY*�g�]�
zJ���f����1\��8��A�!vۑYՋ��Șn�� �㴄gh��Y� > Q��:ۚ�Z@�9ٴk:�]`nK��ej�s/���s�e�6A�~uy��b�e�IV�L�n�=����P=��,���v�px_. ��ž�kWij��RM�P��t�1J;�Y:PǕ�E*�DtZ֔�X��W :*�;z> ����)P�f��2�f9*;ª>��٫|��-��_'���j��.�c��|�C��)������H��wgl�co���̀�����r�[_D	ϒnz�jJ�ק1o(�Sy%u�8���װ)M��;���A��S��2m5���֊�9��x5
�J�r�U�G�����M��)��&�rШQ����+:sT��� �{Ei>�����dTl9.���ʵJ��wwز�	�u��G����FČ(�5��A�4�Ժ|q��(���S�L�B2H�����v�������=i�X��-�/�s%	Ff?5�摑�_�q� ���!!�����۷n�^�z��-��$$Ē#�܉4��d�h�%�IH�Nʃt����ݻv���7�|�7��&(�ɲ
E���@�!d$����H�=z���ݻv���|߭�|�>(�W��f��%a��.W"I�3P�(�<�^$3#$E	)#|vH�9�d��) �p$c&H��ut��SD�v�fl��v@)�ĐF`����&Ii32$�@d��d&�5�^n�A(�h��j$c��y��\�9B
HU�ɭ�}�=	�w�ylj�<������D��<�Ձfå���4nŵ�܆�V�^f`��hż�fnq�l��0�lܪ¤Dy�,-�ڸ�%a�ʓ;q��4��z�f�	Ř��.���:�cX�$L�I��\��3�2�7C-Ґˀ]�5%Ŭ���tvJ^��V��⁓^�Vf�����֫ �t��U�60R�Ų�	R�Zl��Ih���lL�J	]�i�e;��4c��&u�	T`[]�C���
�X���X
`�g9l�1�H��qA5�t4����B�k06���:jʆcfțh��:�6�V�V���m4��P�֬�潪�`At��67b�&ƃ5����+�-�,n)����K.Rǭ�h�!�iQ����U�cp�˱��d�b-V�!��j�c���#Y)kVԦ�Ih��L31S6[�iyw+�؆`�U�G4!��QA��f���V������g	�H��hXn��3���,-m^If�&�U"�M���F��%Qdto�����lR+JM���UH��k���0Ўq10�̲���t�8�і8�m��j룮�j`xд����U!�����L��{q��dc��V�B��Ձ&�08CF͍.	��Y�f�z�%z��WE+]CAsA�ƭEhV��m�
-R�h���$f�t�̶#�1�1X�Fݎ1��bŦE#[�aU���p�*b��u�j��+cr���R=`6�Xa�$BP�4,����6M1�Mf��虎��
s(b�ne,p:ҷ����9]r���9������4�"sڥav׉���Z�	SQ�>yǚy�2�Z���-��9Օ�Ȑ�Ymt
)q�iP���j��,*[��8lʐ�ڍ��H�X�-�#�n��̎�&���W����I� Ю1u����s�]��\ׂ��Ge���T����P͒���yg�R��!u����b*K(��7)�V����g��"�l��of�h<ـWVj\���~q�q�~G��`�W�Q�gA���JB{��r������l6e�5l0�:g'8K4&�\��k���Җ��]P�<2P� �j�;���b@���䶘vV��LXT��З:�J�c+��E�4)�K��o�Z���FQ��越T�1.x%�k�+��nvm�`rͶTX��k���6ԛ�։˅�U���Y���
�K��u����o!�wk��۞��r��LJٳ�)�`2���ѳI�%9`4���i��D�@7l��L�)���Y*{�*��,n�m��M{u`���e	�U�]],w��l�io\	�_�{�o�]��f�3M���B�`.E{����j�y�+��^�>>��p��O�'7�d��r�h&3�e7�	���0�ٙPޕjb{e��*��Y��W�
�}!q �@�T&�C4�ra628�����:|��bB�co{g��*���3@�y�rM�����w��V�����B�lPÄ�죐�Rf���5-�!M��j��ڗf���ϟ>Co;��R�#��>O>����j7��#�U��N�es�.�4�d�+�%����DI���`���d��g�� w,�Հ-�M�t{�d~޳GW�Ɵ���
<���M������;��eySs,X�b����z���f��JO[y����^[jdi���\tc8�LY��P�Bf,b>;����3����N���ב7�(U���[֛���8�C�Z��[��[]^�o%8�;�?k;U &;�hu�׷��#�s���k ;���q��0�֪۽�1�~�A��M�����Ϸ��.	��צ&{� ��C0C�*TؕѴG)�D�������v�î验�~������J=�>���oٳ�t��{{�,wX�x����6Pi�$	@L���*=n���[�45��ެ��6Gb%�w�;�<��N׎L�mT�cU��5�h+�XeZ'of�%���X�h��!CJ����΃/,]�2��Wv.[��I����.���s��Z�bŋ-�i WS�I��I���[�ر�:�eL�4ƜsNM]]ǣ�u�m���2�3�Wy�u�(O��3@�C��1ܟ8��(�u���{L!2���N*�{=E/{R82��@eex�纯f���ָ
��M3Tn���'����O=��K�xe��0z��[u��u�g0Y����DPQa#��3\�3�S(L�؟Nf��W��ݺx{�6�ȄXc�ˆ�fL�9����s]�$6�2�E�Vfl]p�뼼�&��,�L�݉�Vj���}�g�MT����΅�Nɳg���js:ocƸ]��3/i)7vr,��Si縪�ʢp���z��){��k��~(��/�yU��f�ɬ��\�߹���'�,ǿZd�;[�ٷr���i�N�[S3�9���V�J�g�d�����߽�bŋ,X�7Bi�߽*�ߠ�g��fu쵓�C��s�V�����w���� ��e	���S��2��S�-�폾}�?`�5�`�ĵ�+-�D�]�;l��*B0RQtfE�w�e<�`����ɰ���:/^���/c��Q��ڸz]�Y7f�l�����`v]�.�ͫ�Ř���Gn!�?yN��\��LN���z*j���ng��Ff�z]��y�֓��y� yI�\L�"�:��ODFZ��vEֈȗ���I�T�i��(���<���U���ا}�Ήף��~ǧjq3��	�ʙ@L�T�qϺ�loL=�+�dEM\��ᐘ%�@�2���r�+�S8y�MU�+Z�"1�
>��N[L�۹[����3{�ٵ`����"Ҙ_c6${ƪ^����y�=�"!2m��Br�(�^s,X�b�0w�)Tν&|��^P��Ce\g+�\,ۭ���V�н��-���*������q5���d���%k��5+t�6��fbm�5 G��J ˶��5���ڐXB��̎vY�8�i�.lB���j��`M����7lY@�)�im�2�oP���R$�܇R��������ٮi����YsYJ�
 �v36hy��dmb@��8r�Z*�y���Ϥݐ��nL�6b[ ִ�V*�&]q]k5Ă��(�Lz	*�u0�S(4�eT_n��dME��e�����O�{�m5S��iy�u��ޮ�Y�5˼�q�Y밟�}y��zA{���Uy�S$Tr+bFӎ����(L���yb�/�c���I8)�=��[^؊����oͶ��i��\�K�z�j9P&P����}���Qy͛�j3bS�Ú���2�L����5�"J��J#�v������϶�݈WC;L��l�z*-&�]���LBE˹�!���+s�m��`&�Zl2�m��	=|���>�~�ou�l�W�����t�M��:��OGݠE ;	�2�򻫏s���~}9�B��'0%��u�3E��/^gAU�r�K]!�z�������b�=��7I���-�X�bŋm<�p9≯�lm�9{��e�pv�p:��¡�0Do���n�k���,L��x�ڈ���z:�	ލ��ľ��7b�M2�d��Dni�N;�x��b������^Q�J�GM?�H�x�v\ٲA�e6cn]�5�dʙx�Y�N��'=�r�3�������̼ᒺB(	�}U�%��@��D�w��f
e1]���WYn��	^B%��8%�ߟ>N-�~{�)���*V]{��}�	�{���U>ϝ�U�
!����[h6�N1������׌H�UM�^�b3<��ޡ�P���^��k���g��b�rzd�t��2��a����3��d�GM��]sP����uGPn���QwK��#V��}Q![���(�sQ��cE����ɱ&������Ġ@> �1bŋ F ����[���l��߹��f��" P�)�޽US�V��x��lŴ��eT�M��u0e���[����{£��{�U!�3(bf��>m�A���.^�hܨ[�UWç��l�2�g��ގ/�W�S��Un(!�0��D�+0�T���4���vdI�B"�"�t��PJ{z����5K&��{�U�_�Y�-x��r�{^�͒��m;����85O�q�$My�\e�o&�k�	����_��}ñ�Ζ�ѕ��C��/�sm��5�a2�(LƮǏO����P�p���e���U�����ɺ�y�lջ��G<m�_U��u�k������mW?�]fU͆�xn��y*�va���oە��ow�>o�&��q�7���.�<��f֥u�n��{w�����e҅�B��Փ����-��UG�	�,X�b����kKQ�Ri�NU��ɭ6V�nMe����_��x�����	�!X�h@�7L�!<�3K]H�&EIAJ����g�Q+�B�ڒ���ᴱ���6ˍڨ��]~��*/�j�#ç�VE��z�Ll�{-���a3��U-��7��[�~��΍���ʼۅ���(���p7��y�"9��I&!Oj�Be4��ȝqă��ʼK29l�{-N��L�)j�^���3c%�h�򀙣�;��{U]���	�b��kACa7�f�3��*����J7�Al���6�&������2�5��NZ�ګ@�
O�TINF�ϟLl�~9PJsv�jz�{'#�kp�4�rh��5c6ig��V�{w��ik�Y�^��[m�fJ��g�FD'�i݁! �nbŋ,[���zO��s�8|�)���!�C�.�$�������MՖ���2�.]�i�Ź���K�,Ԋ@���A���V��BHLj��Kb[[M1y]4�b�Ck)� �l���+n�,�L
8$CD�CHuf�v{-��-��9�U`�ʹr:�g$J-��W���Xv�����cd�f�2�Kw�
�n�dXm�mv��7Q�S:�w>���F4=L�5K���v����є�
Ў�]�ͭ��X!9>m�8���U�w>~ښK�l�FZ���M�2T؜O�ot�W&�@��E��o��Y��@�ں.��������nt���){�3W��Km�{�߇�V�y�� ���_h�5/�j��**�*�@�!ҦP�3�{��t�㷡�y����K��l�FZ�nlc��4�˥Ƿ���	��ϘL&i��À��_>�*�qСz&F\ܗ�����p�i��qv�� 1.��	�)�ȉ<�Ʊ:��1KkDF�­�� �Qr��%w�99� �x�2��\�]�cw��\�TnǙ\7%U[�ʧ�A��1�S�띃�w�>�G�ŭ��;����y7�sw�hҗ��,�>y����__�'8���$�+�*.�\)Nb�6o�r%��,X�ld幢��q*2�k��l�{-O7Zmk�Un!�T�b�k֘L�2�M2�(��9>�(ܯȽ|��̾��^cԽ!>g�߫�/cǰ)���|��׾��L4�m�_ul���Y���1��5<�[w��|�����.ޕ�-��Pؗ�;ԣ�����l��e=ph5ra2�L���ۂH���#�
d�yë�̴�l�΄`Rи����*n4O#��{��I<�fa��UZ�'w=��{�����ن,��_�;_ֆҙf5�����a~W/z��i���}=�f���/.�߱� ��Z��CՍۈg��ٮ�h	��(4ˁ�sָ[N���x�qXV?��
��,Txt�nSh�yf�lr�˼�If�#���H�ۣ�k���M\���Nnk��+y<�ޫ�g�w�)k��=�Ϋ�34U��f��ͧ�̫�@j`�δH�xX�y[��s#�ٍ��w����|�jUu�9n
����ٱ֡�(�.o�n���r����1y�d�u����<��T@8
s�x#˃����A=�.�����ĺe,�;~F���G[˿�ӃY�b�U�c��p�;xy,�s/y�XG��g&��1����b���J����V��P�д��fe�r0*܃���4߯.تF:�m�]��[��E��WMR���n�>(Xs�2b��s�����M�{Bi�HTʏ�cƖyo�̻�T{�� ���[��]C���@,�G,�z�gX���i�R�j�6!�4Lv��WϘ#�&qb4"�j	m�enp�Gޤ���(��Ƴ�$�"q��to8��ݤ����2���3΁���Ʒu���ޣ"r�t�oM������,��;f�\ �;K�Ϡ9b�u�*�e-��xA9D;��:��6���濇W�GgPX��ą�.�j�Ý�,����-��%�0R�J���y���\;Ka�:U��K�cXr�t��7"�^�٢�b/�	,�e�e��<ɐ��כ���sh�f��6e�����>�M�j��//��GkG]�X�}��5ٞ6���[������e�l���b����бi,�U��Ғ����%'�]$LQ|s%�������׎ݻv���n=s�$����;^0k!��:X��D�"��O^�}q۷nݻ}z�띠���pl���D��\�Q;�@���t�o�_^�v�۷o�^�z�!g�����(�5�R&�t��0I��>=z��۷nݻ}z����$aI�9~<TF!$��(����D�C�R�%��"���b�X 77Kz����}5�Q_M�����J���}w" ����4gۄ�3{�Qb���\�F���g�W6c42l<q����Qx��
1G-s����U��,�+չ(�Y4�� ��lc�5��EW�����j����{2�����L�&b�$
�w�=�R����u�W�	���h�d��*���s{��;q?��^��۩�Sm�eJ9��֢�2��y�j��N^]��J۪�������F]u`��yP<�!ا�)�gUݘ��L˶�q�)t�)[7jJ(i�k5'�~��o?}e�OT�1�M;^���_s�wْ�͘�P�/S��75�e	�!��E��r��쎤3˥6��R�=쫌���pک�U)��3\"lzZ���%�SL�<��t���<8�X�m׶�T`S�Yx��1�I�R�C�{n7-R�^�
����	���9�[�}����=p�&��]�P�Խ��l��]E�vic����%u�=�\&��ò�ѷ���'��	�i+�w�y���ޭF��y�xW?}�����š�8zT1�A�	T�i����
�S��_���س��}�q�]<�myĤ��3�u��_O]�%m8p�\��!tK"�����Y��eŠ�p�:DC�!�8>xzPv-�U���w߾�f~�;_o}U<��\����(vc��Ů�b/��"n�ܻ
�g�~۽�;7�x�;|�ʨ�����JͶ;�h�l��HL��>m�]P �Y!��_.����=���lg�.��b���(�Y��:�o!�@L�ʘ�����.s3E�	�z��B��o�����&�,%k=T7�3q�w��nz^�U��0�\�ޫ�UY�����{z�����Z<�n��ऑK��^�a=�wEl�S��^�R��{Տ����V3LU�ma*��w�²R�����
���E�x�y�:�
���q�qǳy�~}�~￞�ϐ��a�d��8���BQq6]Z�-1m�X���Ĥ���\,%d�f��bX�#.��t��4\�8f �N�ֻE�g��j�0��u��Sb
tu`nV�5E��-���-[+�Kf�n�f����9iu;�t�
�sR1�A�z��4fV]렉�[����v(cG[�sM�)���z�~��㽿�iEn�ro-�\���pVQ�@�y���o#B�A��ˮ�+�.�D����|.�ZfL�&�'�Ͼ��N\�WV������b��m)f���6i'丟��Hkc�߿}��k.s3[���A������-��n��Be	���b�W5��ͽ�:���+1�õt�"�� ���TC����1y@d�2�U'��?{�}9yY]]���ϗ��WO7�t��FuT
�v�S�ꄼdg�r�)��TM_N��r5�9���4Su��av	�+#m�r=Q9.�r�b
��LWA�v[+�$ͱ��$�3��8�����O�=��~_�M2��q�����x����o4J�?9vRY7�{B��!B�L��+*|x���sg�п�!ݖG�1e,��gF��ISy�&_����G��m��5`8�o�Ȩ�e�p#�R�P��C��ŋ,@,XS��N�^����N^^WWdu��;���ץ�61^�q�.\4��xD��f�x5٣��~���Ss�-�5�9��<��	�&P�CL�����	�kz�[�����dfz��:�F��pˏn-������Ǫ���iH	�ʙ�V�
���q���͘�NffWP���fdu�8�wXL�K�S��%��ra%�uX9Q٘�����A�r�!"��/�p]�k-�Cy�RLj��U�F��P5�9���3�(���fC?����)�uu��Fڪ��V��ł���Ƙ����}��y	���|a�}=nP��x�s�����i�&G?�w�?sb[��&,7Hnf���Q�_�ﮀj6�5���*��ۈ��z ��L�kn�ݾ��sj)�Q���SrL8���ΤM�1bŋ,Z�� �y��ۘ�M�fV�nĀ�S)�P	�K���|��W��1 JaK�[��<��������8okV��*��5���B�i�� Be4��6����v`&�j����rr"�8eL�o��&P�!uu����z΂Agꯏ��6ڈ@v�,L�qJ�Z;RTr-��*C��SZ�&��@�gCF&�e4�g׏ek�Lg��3)�xsmm���!=u\�f�l}�P©L�(@���^>����C�����yuYu��{��;��lW��/��$���[�3%��c/<#�F�� �?Nu[��|7=3õ�癖peL�ܶ����l�����'���t���/2�-˰x�gF/�$@���~iV��vt��Q���=@J�M��EY��z��Ӧj�sU0:Ȟ�T��N���*N�ծw�Xl).�ň�,c��Znj�j�TȬxz���_�B�OZ�]@�^e�^�T�B�4י��Ǻ�bbrP���9@��ݖڻk)W�A&-v�2GL�u�dB񢖆�a���>�>�{��j�p)xOV�n9)��琙�Ml룲�WM��gET��0�@n�����F��=h���I������Y��l��uL�u�N�0^ُIhoS�庄��0��1.NG.�5i$Ͻ�R�Y@�^8�v�b�;Z=ꪮb�����6)P�I��Lϳ�2��)�/��{���ς]���]�yS*e�|��"6J&dcb�O޾V�궽�����C6f �ӈwl�$�[�1��U���{��Pm�h=�K-�vS0nӃ�N��ܚ�e=ie�@��U4����42���f�ʦ�fG%4���i��xxxxxxx�}��=��8����fU��d�eM��cYc����ñrc&F��+ \��UDi����[B�t.b��ზ��43��t �&Z[p0ҹ����Xŀ�cC5�3mT����^i6.�1��tگ06�-�6Pڶ�Q�-e�GKiB�s�(b\�W5M[V������V9r�õڻB]mbѕ������t�;�]�tעGom=������M��&�^�ut.�ؼ	 ��x&H�a[��җ9�qWD�A���wN��R�t���U&�@�%5��A�Q5���N�;;��(�Ŕ�Ϥ��G`�]R���qo]��V��f_�[k]�\H.��0&C���T���&��.R)�`�B|����b
O/^�eV�fW�y�͖pe4��9��C��l��si�Wy泖q>�&��+Ej�s�|��hygV�y{��Y��3-Ťة��n�t>����]�	'n�v�W Tfv�L�ɽ�ecU<r� w����珿V1�S���"����I�-����E��X���3�P���Q��7r(L�]u����̯p����'V�/�jlo$�1I75�]����}����ْ��gު����Y�����*��v&:�(G�)�����Kd+�o�n��-,�6 �(�E��G=�VI��s,X�b��7��Jew��v,�}�Me�[Z�b:��S_d�Ľ�N����l3��y@L�7��n��c��$�ϱw�����[����t��*e44θ��H�i���3�BfY��􎗞�Y�=l[����OBz�g����T��Rl�@�h�s�x�3-[�k7�Q��k/2��s,�i�gr�T���I�τC�&�]���h@e��1pɱ�Gs��)]�o�Ͷ�j�2��*�9�����}�9��g�C���GsЬ�7lm���2�e ��l�lݯ4�M����1������І�3�s�2:��{}6SD;f ��M<�y��o>P�.���r�����̫�Η�C����M;eL�����ߵ�e����!E�<��a��I�����\�ŀ��QJ77ٷ����^esV�Қe1��U��7�W+�L�]�i���U��eA|�9��ח�"�;��<��Lz;�=*�פ2�/������`?����z��C�!�z+�OF;���.d|��������o^{i��Za��A�.�X�6p�!�)�����T�'��S*e^ھΎw��7y��F���&n�v�P�L��J_7+g��[Z��뜽�¡��������Ʉ�뉭�J����M2d����g	���3����ޕ�z܌���6si����fG_h��Ue��}�y��T���p�^�)�Pxy�ܮ�;�x��X���5*^9S�8L�y1^��}1�9:n�D�n�]s�{��{���,�j��W�	5����u�̧��r�9�$-�[�� y���yYlS0=*e	�����b�ھ�J_��d���^�&P�q��.�Rw1<��u�8#S��"���mH�8�J-�[�Wwwd�AP�<"��4�
�� vL�L�I���g���s=�q=U>��ơ�L�3(&SKe���E[�4�����ye�A��O��{�n�|�_p;�?g/e���S0&j��~ݾoG]��%�w2b�0�^٘ecU?�����W�u�)���+�Ó�V�3�S�Y�ׯ�U[���x�:1�pf�娡T�UC<�{��g��w^c��򚹟^�33�G��'�3jL�(�PG����1���H(����
4U( 0=�����ZA"b�jVZҲ�+-�bͪcR���T�ԭK��U�TɩkJ�m,Y���YkMFkiYmL�2ՙ,em++YX�f���,�R�L�f�5i��Vj3[J��1�[MI��c&T��m�����+56�ɩ��dʦkY�ki�ke�Ͷ�,�U�c�fe���dԫ2ՙ����dɌթ��ͭ331�VjL���3,��&�֙���Z��3kJ�ƥU1�m��6��c-jc�m1�kK,�ml���MM�,c6Ԭ�cR������ifYmJʴɩ��em+7�m��Y[+6Ҭ���iYk+-n:�V��n�Օ�iYk+6Ҭ��ʹ�Օ�iY���iY���iY�+*ʲ�Vm�e���J`�*@`��(>ߣ`6 �����b
��Eh��
+���b��(����*�b"�(���
�`���� ����ZҊ�(�*+���b"�����
�`*���R
+���b��(�*+��i�@�E`0QXTV�hB*�`"��(+����ڕ�����f֔�B��HA 1D��VjҲڕ�Ԭեe�����"(FD"	�Ԭ�R�ڕ�����b���P��@b	3V����f�+5iYB@`��'��!�P<�
=�?�EAAX�QAc�p+������������������_���@;���	�ء���;���~����(* ���?w������
/�`� ��8���@! ~��H��?���ޢ�*��~�>���/�H}��6��!��r������t�O��
��A! �VԛT�mL�M5h�Lզ͵3V�6ԩmF�6���V��jikM��٫M��*[R�mKR֛6�٭J�mJ�jZ�Դ���[SeZmKj[6ԫKjVZ�imKjkQ*��(X�E:��mMM�kR�m6����T�SeZUJ�TեKjU��j�J��j���2ړ[L���ZYUJ(� 2ȣ"��,���Z�kj�[j*�JUh��"�B ���J��~��?�E�@E$ �@P�_���>�$���,���_���"�*�?e�~�_�>��l/b?�a����v����}��W��!�S�����"� ����
�i���?��E��?!��*�
�� ��BP_�=�9A������#��h�PY�!��w�?�E U�C� �M�����^�p@A�@���Ҋ ���?��o�"�*��}���Р�?���4~ J'�P1��gA����D���� ��{$�M����@���� h?���~&}/�( ��l
�Z �S�?ӟ<��
C�O�����)��W� d0l�8(���1O�\                                        nr� � �$)@ �PBT) 
 

� H �T
�

*����J�@
Q@@���I��
D�H�U��J�H�R$U(�!R�TEB�U@��*AQ���A	AP"�"��Q| ʒ��QE"UEA% � 3���{��yi[������ۦ������Qޗ����zem���J�w��C�׍�ZUc�BP��z\�J�O{��`h�J��� ���������A@ ��%q�(( ��h(�`咜FR���3Ҫ���DD��ԩ��!^���^��;Q�KM���j�)H"���ﾒ�T �HJ�I*����*�A�^wt�2.��W��w��驣Ǣ$�R�*��Ƚ����(�=�u=h[\��6m�BC�{m5��y��J�m:�((	
 ��_9�N�o��J��9���=��{uz5*��:Ŧ�gWY�g��B�ձ�Ug�ڶט��j���x���p�'��W*�(**�������UIJ�*"*�H�>}J�ۄ��C �' 5V�H��I9iP�-**� ыR�n�`:͊���uP
(�| �������E\�:� d `��*K�8�r��� =� z*UT���  ��AU
�DRT�U�. d� � � ���M���v�� �n� ����l: 3�� ��   �� ��= ���8 $ 8��; � c��\ ��@y 2� (�)%>   >��$�P�A"I$�Q� lψ����b �"p [����� : [�U+ f<���J)J��  ��� �F� .�R�� à݀ H�;� q�J�� -� v���@���$�R4#MhE?	�RT�  ��U��   6J�%E �'�UD�#	�i����QХ$��mA�����j?�?�_ؒI�rCg���>s�2����e�hC���$I9F��B$�]�ն�ׯZڵ��m��U}�$��! BH�HHH����k������[7���C���h:ٙ��how*lJp�,�(�1w�{�������Z�����q�<;9W�B�Ą�q��Fro[�ܝF�O���R�@�KL9y1�]Z5.W� ��˽��5l�.j�ޗ���j�$�2�8a�a�����n�Ұ8`O��ʣC�<Ĉh��4gm�Q��7Wf���@��F������`���G��ߜ��zq��DJÿ5��S�mNi$/x9�n>�����g��v;�=�wx���l3+\u��z��=B_	S��Up���ȑ���3'����;��ra4=�5�!��]�;���3��
饃�&��y�Y7�Fs�b�^ v�2���8�v3�p=�7$�K3��i:M��K�y��-:Wo8��EO5Δ�ۼRf�c�.���	8Q���ڀ,W�����qn^�V��%i�ȣ�^�X��o�b����e�ݽqn3#����/ښj,�h��t,�d�7����ͱ\�N��N�x�Nջ���vtn�P�4����gyf���ߌ��$�a�P�\�v.���);���PDmUK�W���gU�,�J�9r'1��J�\��x2wm�][�mr�N�6�R�A۳U{�QWww�r�7q�E�ׅT��N���r��@�#��lx(�����s�M���f�ӳ_=sL����{&���ۘb��w8d:͓
���*���'�.>�	�.8�� pV����Zn�Ӈj�zUh�C�]��{�gZ�g�7�Y���[o)}�J:@�a��E���ܢm�{�=pr�Z,�V=웒�FF4l� �dב_6{Aj@��ə�����z�cݜ�������)ӈ%H��ۈ��X.�<ݝA��{8f�Sѳ�5= ���G�9c4dw��wYx�.7=�4b��'Uǜ�wAS�Ǫ���b�Q�-����̑���_ۆWP��X'!n�{�8�(�wX���p�����݆
9~�jӵ�;;kL�����[��p�:[t��v�����P}О�v@�Z۴�b�-=n������]��-��	r�[��:�Տx�LÅ^�ģy��K�f$P�F#�1�s"[53�Y�n� �$Xblsu��_d�X��Y����R���%�T�)'$�CV�X'��L*��2�� wZ�����p��Z˹rn�a�Cx��uI�b3R<�vo�]����M_vYAܺ����7��f&�ې��0�1�5��%k�J�˜V�r%�g���p�M�A�x܏��@ۚM�=Ԅ�X��Y�%�b�}۷��&�5Θ���@k����M���`��H";����˺����puⳞZ�����vjY�N�3����t����6�w�*s��;�wCÞ��hT�J�Ý��I��n}�vR6�	� 9���N
1�8�Rb:�6^�A�6��6#��~<�T|�,����cއ7���8����e�>u��y#���9"����D���'�p����}ka��)��˹q|	5u����sO:�v�lt��<:��"\�=��^=8�p��9��Dg���;l�ƚr��ʣ��n�{J�5v�8����=����q�����Z�>��gv��ȣ݁��X�96�K;W<@���׵���18��{�X0�"�.��Ii:ͧ�kP:W3�ט'>p�}�oJ	ٸ�p�h��Y��b�B�K��(kF���Cǅ���0��ލo'�*�\O�n�嬲�6M�ʲg'e�ڵ��hީ��b7;H�e�ZW����t��5��{��q���O�uS�ɩd˝2\A.�M�sUخ�e��wP�M4�����y�)|wN��Rk`�'j��:�㬩�׳���[0�q�0�D�i�C��\�������[;��J ��	�8�ϧk��|�L�x��V�m�g>��'P��1˻���+KlY�p�u��p��mi�Ǫ�N��J�3��=�ۓl�5�È�X�Xlc�qw[�,����ޫ%�7xo�AC������	 ��y[�P�Bn����6ݯw�2l0nYn�f?yp"9����X���6ٱW7���B3o�z�M`Y+����+�h��v�*ӡ�5Vv�uJ{�,�P9���Cx1��9�-�2�C��!�����u�o�\�&�9t).f5���7+�M`6�fQ͜�.�w��;q��x�1��Ht���~;a�Ģ{n���D�k�ۛԉ�A�Pa3ڎ�'��k(�^�le<��b	T@·�:�ה�`�p᱆�!5u�W,ٺ���ъ��1mup�S+{�#�w(!�2��9�q�9����74�c��{E��h͚��H��7S[�C�VbA��81�Mn��m/��bM�9�0\ٹ�B��b��Q����r��"T����h�r�
v�#�2�r�;l�Y���V6q�Ʉ�3�pc���n�5��ad��nP�UK*ы����Пr�p��<��G�R	�r���j9�k%ۛ�ѵ�ku20���h�5�݇�0g ���)�qI���u9�����uN�v( ���gH��t��k}�y����"��yf���t'
6_���0�6B��K�(�m郷�a����#eu��6r=ܸ�s�Hc�(Yf�^� ۛ�W�|�x�Sٺ��Z�is	�{/|�a�%�]3PC��������t�ot�-Jp$��;OU��bU>�iod�<�̊�wg���U�]I��P=��c��Ĵ@��][��{��n\Et,� �&�wk,l	�u�
/Lv��%���+��w9�j���Ex��H�s�\�75��m]p]`���M�k=1�;GG��J��!��� �-+�;�"�;&w>n�ۺ	���pe:�!h�"�����z�(`�/������N�C:1�f��^Z� .��C�j5�^Ƴ�O�K��ؾX�x�h�y1{Vћ��ևN��We��ķ�>��I���:&Aq�v�Br�"� �钒�sA%AD,=�s�~z��Qe���
r�hջpG�Ӹgv7��.p"n���{�A�O��%���S���Pu\i�˗9���㛿t��C�1|�Z����V�u���9���gr���C�=sz��&גH4L����6����'}���V��l:�@�8n��f�.��R&�n���������C���۹{T�{H��-ɩ>p�ۮ����A^ν�N�q�l�+}�G�	��[����[�;a ����[qt�4�%]�J	z;�4)w��Y�T܆�V$y,��y!�qs���]�w_�ݛ\�Ǹ��9e�3�5��;9���/���z�i9̣��^��ɼcV�Fp����6�!�2��S��(�� 0�}��ʦp�Ƭp�~��3���6� ]�ٴ��"�=�!@&c!�������Ȥ�m1q�v��&���|�p�9��+�H��0=�+�0�\�&�q�PVufr�����0B����s�OD"�G�"��%�pN;.�	�*q��c�����h@Tgv�a�v-�f� ���o�-M7����/^ɣ;7�]e�pQ.�] ��%��û��Ó��@X�m���6v^��Rڻ��(����P�g<{U�m�
4H��sR[��������έ2R��0�Q*��;���٫]�i���,-шn4`痉/j� �gNW�J���8��b�\	�Q᧝L�Os�Yh�S���p	��)�S�-�x[m��=�SQ�M�R<yxR�/���V,Н�q�s�m�2"�q����eǻ?=:���� }θ(�@֩�'��f�XH�az���b�S"��N�\}� b�}/h�~�v�����#ud�5�r�(���&]?z��D.ɡo٤����g����x�;c+	b�w��A�({+ ���"�N\3^݋X���9������p� ϽR��8lc��|��#�U�����Wg	�c����tA��{��H���M��,���� Y�����9�v[GR�$�+畬��VM7�7���uL�o3���-ZI=^�SF��akh�ٷ�Z�N�ˎ=I&�L��Y9>�gF�_[]�k]4Q�τ84׊N�f���Z���eg��j�hi]�X8wCǱ*�JS����h3x�E`�ηb������3��ֹ�0�^�Hٌr�!��+s��k� ��b�,,j��E�K�S���t.��u���v
`X1�=�(��T��PǸ��Q�G%g��M��fK$ͺ,	d�u�ٻ��y�m�64f$�2�K�6. �Km��y��u��흋�%�X7e�o^to-KAa�6�n�_h|c"�{�J3S��j汙���w�w6I�,y���(�N+r�Tuj��QY\�K��n��c�Łap��^����#Ar��ϵ�H��<3{z�VB��N�z]N�v*4�^��P᧺P��t�[���cu��-�2���e��)�{w�����"�:	�.����7IA��&C�$qEøݝ�U�����G!�N�Wm�{y��y�M}��fwn�Ʊ��|�{zΉ��1>��|�-�I��@��a�\������q�	����а�F�vc����3n�67P�GM�1�W�b�sW[�K������a}��v:Peۙq��1f�Ut�s� i=��d�5��p���8�x�Yws^���\��ի9pX�l��8��9Ѳwp��J3w��W��s�"jCVQp�0(�a���ccO�t6
0����ѷ�we[�n,A[7�ni�y6zwv �\�۸peg;V�����`���'��(rڵ	�Em�U��:�xMp;�1��s_gU/v����7Z��b��r)��n�2k/�;!)�.�\��u�܆����s��14gw%ɸ�Ϯv��a:�Ǽ6<7�@�4_�g���X����lѶ�]gnR:4��t]�Ú�׍kĭ����9��	��q��Jf�K�_L�P�om=1gr��g8��:I��S��JIhܧ.����a>ѵ��P2�[����o��E�ϷA҂l�ƕ�NQ�Bg��^�DȂь�[6wv�O�'�+!`��2�� �S�r�۷z	Q���=m�Ċ�;�h�����C��ݖ�]�rp8����e琧4܂�wXbkGcm'z������������{מi]��^��!t��jx�sx~������8u�w=�cyؠU��v�v�������:e�F�t�ȯ�;���^�5�bQ�q��T`*�+�Y���jY;���p$��AC3�aqls�{�H�x䱭���of� #�.�z�Ft�庢��+�q�5���؛sI�;�`��Ҳ��muh�������x�VK�NKH�q�7��˻AM�x�ו㣞U`l�D��v� �|	�|��>Tʳ�BH������,�;OwY�a�6Y��61+Nk�~ m�ŕ��t9���.-�|x�B}
|;�5B`hE��q{�(}ؙ�>��&���޻�����0x�;/jNb۰7o<k�_��:�r�����k��{������;x�0VN���t��l�,_K����XA�8T�ٹ��,��ONЩx�� :z�M�c;	91���4g.ޠ�Y���tXk�؞��o\���K�ENt�E�e�[���(oҙ����org�N��B׃mѼ2(����mS�k�D��&w�89r�q���N\���jWU��K�#u��yŦ����&>O��W��i��c�8ɏ��f��(�A�������h77���^�&�zk!��{�-cͻG	���z�4��T����:�7Qi�/ �p!�,��8b���:�_v⣵���X}�B��L[�TR�f���>[��c��.H�ɝ͏�2��
��^����[�ݢ�˱�xk��lU��q,�CB��n&�N��CE�E筊�"�}�uꙭs�E^�WbR!�C�0��8�h���5��̝�S)Kf��t��U.��][3�NXV��B���$(�U���Ih���ҧ���.�vÉ��"ع�)�_	����x]PM����2A�h/.Z�%{P#O�v�S��J�^᳓�ׄ�$S�r=�}Ɯ��k����$���d9:ٸGs��� �][h���p�{�{�:$�Y���ݸ�۸vː�\�vƱ<�=A09��k�^EVWF���Nݴ�����f�< ��e��e���5P�;{�^�v�$�7a�
����ݦ�݋
�㳰�q3)Rf���b���0�{��w����ݳ�K]�H{Cm ����ߢ}NZK�V0b�;g
�M�����w�F�#F�j=�z�i ?|(w[��yv����v;�ϵ�.4��c�v�7�%p�������%Njnf��y�eg�6�����Stn� �TG��Y�\�EN�P�sY��{�?rݧ��e�b0�=r��`�:V"_:�8e�<���z����s_jL�{�cw:]K'j��!�4�t9ŵt�#T�����jKt��B֝\����
�6 SP���Q}�p�f�}�1p�<rF��t�\[����q�
vM�𻃹�8�����5E[�i��
w�pP�<Ͼ���j�[EV�ՋmE�ƫETV�[Z�m[�Qj���kQm[V������1Z�Xգm���kQ�-�+lk[[V-j��5�6��klU�m��ڱ�ƪ-�5�ִkm��E���h��QU��+UF�Vت�5Z*ڊմm�+kڊ�kF�lV���6����U�Zƭ�[V*��6֢��km����+cV�Qj�m���m�+TUk[�j��j�Z�m�k�U�lmVت�[F��TU�UZ��Tm�k���-V��QmlX��Z��_�$�$���B$���g�W�_�����~��)^�ʔ.Z�`DmEۋ1)P��T,Rm�������P���[n'�[{nnm�9{������\$�>f%�Ӝ��t.}Ў�}�ޞڒ���Hi�q�}XT��#0)
�D#�'���]ؽ���g���&��n����C�ͪא���Ҕ��ݩ�4�
6�M}��3���[�	VĦ�)�-ҙr��;����A��{f1��V^z���S�I�>=���w�X���o��
o�~n$+��/�X��xy�l���<v>�5X;�fv5瞁E�CO�q��Ɛ7�f���c=��og���M۰`��1��=�rw5_�'S��G�=/e>59==힨;�����+Zs�(c�e��:x��x��y��<�91�	v���.֊L���/b~�X�~�V�ن�&IF2��UP�b����T��wʙ���B���Ԇ�yu(��$]���<����l��醢�77:�l]Ŧ"Xyz%�C��|�w7�"Ҟm�㻦iҲ��[�����
�cx�n>zx�n�r�F��J~��#.����D�N{���'�-�0桮b�z��>G���ޏ+�7�缡>H5	�&��O��o��r�uQ��x�|�Џ��R��$
}7��ɾO�φ�E�₯�z�A���ܵ�Ӽ�n��F�A�E��2{�9��PѲ>�$����r_n#��?�ʞ�B�'x�͆���k�P��W���9���Y�W.wi�z�쳲I��Aۚ��&e��g��Ԗ�7f!���:��{�{�t��9�Ǐ�IO�wt;� 
v���F˘�V���)�P��`�kt5f�����c�lJ0}�e[�^��Q��l���|���kX+���ý��Z����<�m,�s�����:&�u��Գ��+�ι�Q8i��=�2��ۋl�}%��A�ݻ�}1��� ��9T�xyd.{~�Blʦظ�/vz����#���`��b��8tVS�sQ�zD�է�Q�T���x��~V�@�T3D9v�}��;R9$&x[��	F����ywr��q@�xo�n��ۭ���� �M�j�ww��9ǹ�i;f{��ȍ~�ۊ���V��I��n��y���������h�	��������T9��xO�.�kWM�<G-c;��;�-�AoI�(e�BA�;�,�=���A�Hf��Y���
uÂ�25nB�=1 �86ξ�A�J��Е�w. ����B9�H׌�������y���߳o'܏oKs�.�՞���=ݵ�5�?[�"�$Q��vI��S�pBL]�K9�������q�vb	���"n��x�v��8�#��7i�'�=9c�xx��^1�Kg��{ѼQp��V�37K�_v�c�S��'�yE֎��$�*#r��Wu�Gn�>��J-�n���Ѝ�0P9)���w�^�y
[}�q 0�C�3o{�tI=��z%vaz3-[��~�Y���NΔ��˕�oH���t��z�6u���^��oy��s~��%G��|N(y�k�5~����;"o<ߦ.����7�x�3��������V�gq>ݯ�V�hd�pь^��0�G�Ϟ;�KE�c#)[Ǣ"帽sQ&�<��QI�b�Y#�W�� ��6��#�����"�l��z,�
�f���R��Ƞē',�WvŕR�[ώ>||��(�`�9�������k�ٿQ:7.�k��ݾkd㨬=��{{u��nW�4i�.�J�x=��wj�k/m?t� ����s/#�7:xj�9$^�f�}�{���K��x+���������48��XU��t�N(ÚS��Ʃ��2ax��NSK���c7��Cy�c����>4�=�o��OU�J/}q�e*息�c%�{6oW�o�7+^>��{謾�2�Ӥ���<=�֭-	^�{Π�R5�H�z�����{�S��A�,�i>��</HB\�!�ܳ��3�sx�/3b���~>=��S�c ��5�o��� ����������m����3���G��[�����=�z������fϝP�]���/vе��1���2f�)�ŵb>q��r%��B[[w*,�i��i�\GQ�p�:�Mmg޶l}D:}�o���ʣ�D3��<�̽�uw�-�@�rw>��䐈�˾�>��M�"w�����_u�=���q�6(�q�+a;��M^7�![�ݍ�ϰ�H[�7
�Sq��19;�����G{�x٫�o:481qӜ�ثc{S�ݵ�ږfc������0��h��������Ϻ�4����p��\w��Y01��X�˯�K���޻K�����)3�<Mʒ��f�?ku^��t|�/
BN��Q�����'sa��"�o'�[�b�������3�O�77�,Q(�^(+��vv�r�b��$t�ɍ'���3��2�j��D��6�&��(B����˝��x���^�H9�K��l�=uxxv�P��<�)����Zζ�lV� �.�n�v�8�˕�+f��Y_�k���Pݯ7����g5���]���\�eGްx?G����[�??��-z78��$�U�'�Z��jg�Dm}�=<A�N����I=�ۺ��u�Nk}�1���g��&S�Fn�;}�i��Ϭ�����'��mk�Z3�i>̭p
��1t�Y�w\�i��l�J-e+��h:�zǹTø}�Dg�=�ɼ��X4��.�ѡw{�l^[H��Mc�ɮ�����P�Y'�����]�9Og�y[���lj'�}$w(�"~TpH�`��5���Po���.m'��*�7��O.s#|x�k{l���[��>G���{���B�o�#px��޻x�(s���Ӯ�{�W{���r[R��7���5����Z�sG��{�y�]\��y���ӊ�F��{{V�ս��<�Б|�w�w���+�т�����i'G�*���d����}�a�KnR�L�E��*����:���ɡX�U:�$��w�龫ú���}�<[�f����^mt>��LHP��|��vW�x^#ş/9�ڂд��S��صv��P��͔ii�L�w	
e��g�a�M\�'�&���5�Q�(�6{s��z�j�nS�j~���Ys ��U�mEbJ�xg� �[7+
վ��x����@H��Qwwz%��ۦ�7SXY�p�l���fx�YO���9�u�y^nwX+v���6DËpjLZ��qA;8�fn˛��r���׽��]��k��g���k���������c��==Ca���݃f���Mi;�����k�fq�tn ��~���G��p�	ƹ�/c|p�l��~��3)�E��,N�y�S"s��ӐW�C�C;S�0��E���(�m�UV�}�<\�ŵ��
�?P���&���Tӈs�[�j7���߁�x��0����ޱ����͂�v�¸l-z�݉$���N�؉T�svn�Ͷ�2N�ȷZa�*�*�4�i�3Z��~�%�vE��S˧I����Ѕ����J��I����]��눴g��5n(	�j�P5v:n��u��=ޫ�sc�}�_9��bZdq/)����6@����=�0W*g_=�o�w��Y'u��CK�9]x�d�#������{�|�D�������1IBpS��y��a�7[�t����d�/v<>�u}�g(�3Fx�-�*�����J'��E���y/+�.�ϵ�I�>��ZX����T<d;ŢR�[�Q,ƴvnYQ�Y,�k�|���΁u�2��ɛ���'�����'��b:K;�4���7|�^:��:�N�Qp�k}�8e���!��ӂ�H{�y���0����Q�xnj�v�E:�و��m��Ʈ�4m��^�z#Ɵd�:w���;��7x���mC[�I��Qid}�,U�Xsu�m;����*�k���i�#�������>���훝�p���P���hy��q3��e`bڱ��4P��S�m�1ۨM{�ۨ�?\��v��=��-X1N�47�V��"�U�+�M��<��a'5�YC�z���g�\����g6J�1S�q��݆�e���ɼ痱Zg{��*wi3ݒ�THE�ll��ad�y]ٝ#2+�s�|���Au��+�7��������'���f���~�ڏ����\�G۠��D�"%:�Ѯ01TA_Zx�11�������M'Y�s��n�ޞܾךJQMj>yxޔ���O�"��7sj��=og���!�c�(��
Duy#�����l˞�q�ڧ��v3�����C24��Fw���ad�<ۼv�F��cLޜ��3�/dP8��>���y��*{���LV[{���������=�H�I��m����n��Q���#<L��۫�y�C���>���	
��9����iK]�ћ�H{-�8"�δo(_%�jG����<�;DU�Lۺ����Y�e����d��ה���IMd7O>��&{�|�a�;�
�4��`���.w��ݥ��nv�ڝr���hڮ���8iѸ+9��g?L����V�oy�"�Z��n�nv[�ĩ��wd�L�x�e���M�$�I�9�}P��'���}���mN�>EX��1�r��*�����8�ݰ����/�fyyw�pT�}�e��gG�z��G٬E��g6����o)��%�^���}�S��{��ުq��R[��v�:�,��ٷI� D�	�B 6j̔�S�!:2{R}7�j�����F�E�ӻ�Ȉ��\5�[�'�>oI�C�>�q�mZ�����(F�X��B�qT�v-�c��=�Oz��N��0�E���@ʬ]���Q(����8��#"���¥�D�ٚ)��0i�T���ZRMKl���	膤-͚ut�T��T�	�3FS��Zx�K�qU��R&�58��q	���l���=��{�]�Xr�{VC_�g�(e��>:�F���7�r˸}J��K:�@|����3BZ�w�S�c/6I����f�[�̃���һ�|p{�{d�� �=d�1nP����`�ԣҰ#��I������+s�sɦ��i�_n�ۇ�4f�-T6^��de��Rd깄Iä�X^�慻�����p�Բ5�K��� m�#~>N�V
4f�|�#�5���H�u/a��g����ɒs�{�Cs~]�|��v�������Ǜ��7+�y4O���nW�x����X1�!˫�.u�.[��xc3�2]^�}N���������`~��2]��OO<?z����woj4^Bl�4h�9�`���c� 	9�,�0�	ѽ��?c��$���.׽�	<u��a���Q�/{�x�௅��k>��wU�k��V�֤�go)��X�_'�s{u�¤�"�����qp�w�x�[��o��7�K��I�3�1^���r!#]���ܖ,���+#��}�8\W���^���Ȇ����~�T��NOGi�&bǄz�t����U�(�1vާ��% �_i����sUWjIC13��f��8V�'`�r�NEě�1b��cgl^t��Tz�tO�1O�^�g��l,��ރ7N�/H�vͬiE�{�D�̍�l���)���8x.�XB�g�Ѣ]�{���-�{.M^�r�������.C�)KM�T����TNNDT�6������B�13U��f�S��{,GڽXS-Ji�%s+7������v�U�v���W�,eѫZ�Y(j�-�]��D}�y�-��( N$<L ���
��Iݴ�]Ы'lTcy����&?)鍞��L!:�$a�s��M¸��Y�5�$�Z�{wq^8v���x��ٞ}��T�o��<���=>���ĵ�������r�e�V	�mE3$ۓ�dny�������d� �iHg)t�w����s����^ΰ��w�J����3V����w�=2�s�������������+N\9�
8�H>g��Z(�ѵ�٣�H�Ğ���|{@/�_��lѷC�}��>̹�-�����xLh�ʆ���T�n#�6 ��N�gd3�Q�z�ݫx�w�:�+9՗�Nm�k�nN��9i%oG�7Gn��p�C ]G���?X|�Cw�+Vx��ɝZ܌"�j��B¿�)Kq���4��C���4��vx�4jб��n�����qrм.���x9<�wk���S��$V\��ؕ��J5�u8�7������)�v�x��M����0^/ñ��ӻ�g9�$�&��x ��$��?E�X�[@;�7l�=�R\�JD����!Z�j`��mR7�Y>�C� ��i�yvK~���n�"��\�
m��(y��9M���s p4h���l�n�D�n���	����|�{gq�:ɑ0wWy��=�Y���xo����On�Rg"=DA�7�F��,hyv�N�s�K�4������R�T�yo����{��!	9Y�܋��g������<�<mx3n���R���|2�?Y�����"�!�����lٴ�u��b�B6;~^��*<Qؙ���F���Ԏ�љ2����*ׂ�6l���%��ۧB�/p�OaO��OuOY�^Σf��5��Q�1�6���{Ӡ�^<ꍹ-^��w2�oS>����ggy��{�K7���wҼMP�0�����G�{�z��U�S�X7	Y$����3π[}��ȱX��וJd�w�~9�*ng�����0k*�|p��P���/;:ʄ����r2����Q�j��=ݸoS�=��zÚ0�ua��s�c�
e,�*���]�'U�u�N��G��Fo8���=2�[�c�T���lYQ�7���g\�Ґi|�L^�(܊!�6ç�fA��1(������R���V\����z� �]��o�e��*�xd�6J�D��jה˺�Fe�7������>}���7��ҕvN�3]��C U�)�/���]�l4I[�9rK]P��1alu�V�`N5�%PYnW�h6�Ҙ�T�H��8�
h6b����.kŅ*�:�
���mG�j�ݠ���"�E]�6��eԾ�Ծy62Ჽ��+5W�����.��=�WgE룣B��S6����(&M.�Kk%I�*�e�D�L���;uՂ��P%�\4�̶������#f��m�ֳ,G:�X�*!�Эn���Z�԰�n�#��0�b���D5��Km���6a]t�3I[�L�� ��o1��D&x���LKe.��6�����.��T�#c�pX8�#�����l�m�YR��k�tT��j ��m����,���.��w��R��b��r��h ��D������v�fׄ�-5\f���[����<�nF������.�	T���S:���ŷ��9�+1̱�j�Zmh�lGj6�c]�q��0�6WGj+���M����Nk���=M,�(�Q&���>�oqv��B��E�ZL�(�]cXT�`�;Kg9�rfX�+�˴�5@���n�,5��:�4��Em�R� �X�l�&�������ln+�U5)��[x�3k]�s���k���t���jѨM���.�R3Z4�Z�:Z�0pe��3���ƩLɥyCF�kAV8�4�M�mU3#�rf���-.jq��R�4ƀ�La����m�ͦÞ���#Hq4�F���f�B��E��ԣa�JY��ᤱ��Yl[qH!H�YL2��XU%:�J�����ħ$J�e(�"ͷk��L$qԠCZ�F�G˱��CMWE�X�fζ��bP[�Ĕ��&��Xm������ئ5��� �V����F����#u��d�U�Ŗ��y��a�)H���[a��Xޱ4h2��SD���6�x�`͂Ue6�`a��!(ٶ�����B�U���òMn,�t��0�-�+-�8ne�lk�s��/�K�Y�jk4j���-�"VYV���m�)*���uݦ5�b%uŚ)3�� T��e�H�[-ʤKkUܑ�ˎrLK,��A���K��ƕ�X˰�b�G�ƛ�n�a�0
����'qB�io;[u�� �-Z[h��W�Yf$ʺU6+.k(GR&W��2]�̈́�L�J1�MtfXF��GU���A�B��x��il�Ma,mJM�%t��)T4���cb�A���i��]0���l45#�mls�fl�6ۚr�8��t�.�1�*G�,��טv,k�]-�,j�b�L����X�{5! �L�`�0K�։j�4��bi��T�v�-�X�ms��Cb��4�iaEv�b��Ui��9���nf�k���wm�x���E�͈�9.�m��ju��Z�-a�_#�M��0@6f*h�RZi�h�b�ݚYG��/+B�z_VR��z��5l	s2���l�u�9؁6:�U��r2k-uB�0�vn�F:�k��^K�ծ�5�ub�X�d�T4�4Fۃ���r96Y��m*��4�vn��s��ۜb�Ԙ*�=t��xM�WC�%xapr��8-4
BQ5�d�2bP��	��ɓKPqa#v�MDю�x�&��ĬM��;c9f��+Hش��h9�]2h����)`�3m��
v�U��E��\�S5��6m2�[��T�Efr;�2��[�ڥ6u(�5�: �&�bmu!U�p\@hܶd
�A�SdtiJehFl�[Eڵ�	cX� .�;e�Ò٭6��`Xj��İ�Fyڂ�I]̥�\і��KQ���:dKN3�l[,S���8l���i�`Z�n΄yL�m5��4�!/�UnVhW[bR�JFXH����[�邙�Sd@K[��Tk�%�Ա��kF�er��%�����f�SHE����y-�p'j�t�k(uf��	K��)X6�Vfm6R:&�ĥ�Yk��)�t�ܪ� �;�hlG6i\b�F�Q��IUR�܍K2�V�6�1����Tv�a�kL���J:�q+5��u�l*e�""sr�v�̩1.pT]f�R��u`\7�n���Es-uƉ)L�	{[�M��ԫB�\hf8��Y�m�]�D�]tu$,2�pu�t�n��GL��֮�iZ7F.,����y�[�k�J!nia���W��iy��� 3Mz���Yn&��]�L�!McB�M�ƕ�ge��$t2ŖӭJ�#���%,R�[u�t\�x��I`�RЎoi�J:�F�T���v��G���r׍�c���5iK��l���o�d�e�%y
�5}=Lu=�Z,]��.�5���69P�V�a�\l�Q�+5CQc�J��V�Ie5&��F1�܍e�ɡzd[���R.���ti��Ý���4��f�M�s0���3k�qGK�z��f�E��"��[�B�&���D�s���քV��`&̧e�bƶ!���vץ��ԳVWYG��`�Cij�Lv��mLT���RP&s��J�4���tnWb��t��ei	iX�.�%�]��]�킔�Q�;�y����@VS��Fښ2��pf���n�me�R8!4Dԭ���Ky2�l2iun����Ʒ9��v����FC�c-R�Ģ�f]���LCX�Z��U	5�C8&��-�`L0.,@�\�M+�*��q/7@���Ǭ�
�K����:�ں�8�l8�;�c,�5��R����x,ڱq
�֌1�tv)�,�e[*��3��1��y�y�vr��(K�c�4Y������۔�A+i����Z5uɮ���7P��
����X�ͺ'l��\�|�g�	lj�1��i�R���ƞCy�{@��Yc�s2���@r�k��e�o,�X��f�ҷ`���4��&�	�����]7D �Jin4�i�{,l�KCQ+W�Y���:��7F]PE��F2����(`�V���4"�Y��,t0=��`�.l3m��\<�
��&�l�M�3W
���n�]�԰�B�(��X�1����ۑfƣ�p��c9�㝲�(����[v�[c��(�!s��!I�gst�F����](�͵J�6!cXƖ,��. �*Bb��+nH��PQ�5��-	�e,�#+��4 f���`��Z�hG:������ـ˵�*ֻ$;M(ʧѢ7k���	CB=�����2�`ڱ��&�Y���܊@��A 뫓�l��a��f�kX��j� VZ�%�n��Q�3����:���]֮ee�⥫�s!�c%�IDUZJ�æ�y���VV��f�`r��t!2��P�!GUŚ\X���O)�4u���vR�.��V�u�8�J1�X��X\�:�&�6*��!���n�R�1)��5�K9����͂�s(�膥J�ѡBQ�8K��1��:�m����5��X�� 1�̊�$׃B�k����v�l8�D1�BjD�c4�Vi�If U��^.�h�h�[f��d�W0m^R�MB�m��Į�0ᅵI�a�ƚ��XmrCJ:	5CQfn�����a1FSK�3T��1iV޲�Yj���T��Ҽ.#�&���jF�0^���M�k`�V�e1�K��͢�͊���TfԢ�[Zͱ)j�[�]��d���ڵ�q�a2�\�K�0J���HN,՛�v�Ms.��&��np�p�A(�,��l5f��p%ږ]Zs�v[�+�95��f/�R�A.ًi�-t���]��	u
9��$ڬalXr.�фcl�.3X9mb�$����2ư��4�ó��J �׬m%���)k]���ԶݙLR%Pe�;5��4�8�rY5(4�a3����f������$n�cHJ���pƢt"3L���V6��:����Йn	v��ۀ���n���P)�:5��1-4B��6��Kva��g,e�l.Bg�R[��n��m����b�a��j�H�Gmc�64��TJ���n���r�3ZRģ��0�2CSp�7&W�皧�������K��TGA�0�6�D�ݜ\��*�W	�]�M�9�oBS\��r����B�f؆��c-���Y��5��L�=��CSTyqs���u�K||(�dD��s���4�3��Jv�c�ie�Ck42�I`�uMJ�ঊ�Km]���[�D�ES�R�ґ�Q��km�ЉU5����X�e��c��8ġ-�ll���h���;p�mjaH�K�(�L��̚��jM�vW�H��2�,�;���ː�t&Vdҗa�`k1v�0к.�e1b)�������aL�ik4����,���aE#.ԚZ���5Y���#f%s����Ѻ���X�P�	q��.�5��3�K�K��9��&l���Qڮ&��L��y�&�fM}�VOJu��rJ�f��i������>���IqV%��;�M�j�B�<��X�� Z��� vȋ�t{f�kY^�`�eƳ@�6�F7M��G6�s��4S1��l+�x���[���%6�Yt�T։F-&kj�\GV�h,pe��f���ց�ncf�֍z�r�fR�hh�[��e��Z)��Aʑ�d��n�a�.�Q���c*�X٥Yf/7% x@mrZ1�qJJR�R�	�!��c���kL=��I�E#�jP����0�"#�`�G\�M�[����mf�NX�*�\�@
�R�X�r&hT�hҷ��1�tq�v4՚�ع�;b%�)����m��,Glk-Dk�t���a5��B���CksF��2�i�bJ:B��/8��B9����&	E��$Ѣ�lm�0a���*ɩla[A�s6��Mz�$����(��m�Q�9ib�*WLX��kƣ�
�en��؂`�+Xm�m6fvX�g�76�M٥�BT��b��8���.���E����f��f��P�5��D��5�v�=�4ƍa3�����v�х9��:�4*�鴭�ͽR�,lV�b��F"LQ�VJ4�5F���lV-��b�Q��h�$X�Q����XƍQ�E�F�ՋF�RPUشb�5hƊƬj,[Ib�Z4&�
�ZѬkF��L6(��bѢ���!h��ب�lT���Z6ƪ���J�5mD��kDQ����cc�شUkm�ƌV-EI�5�mU3�[֖h10.�3 ���G.�QM5�	�ʅ�q��)�-�R��~oP�ަ���SrBXBܒ#��f� �+r�mtHc&�� uB�tƣU]3���+1a29����7F�ں��T��`̒�َA4�au��Yme� ^x��v'j�HM�s��j��ЈE���k�\�4�2GlA�ҘY��qH'%�8)st����B��a��kk\�lܲ��Xq��M,�jls����]��h���jZ��+Bձ�l&fI2��	V���֤R���K�a)Bhhˮ����4bB«p,�����KCm�ī�K���eΔ�cl
���i#xK�(KvBS1�jݓ�WJ͋i� $!�\&F�0�[�au��(mf�#J�Pm�c��!H��9ݝh�ݍ�M�&ܗM�+������ڄ5+��Ύ��Ց��r��90K.͛WJJ�ԧ-�,AE�g3@4Ut�K�إ4-���Z�1�R�D��p�4��W��<��.�]�٤�Q��A6����]H�-&ʂS<2�2�R�hj�*�3!e�i,��ؑKĆ��g84lM�VZ�݋2mx`�e�jBl��xk4f���X2�C<�K�=�f:�ĭ�%^�ۻK�H����#D����ŪX72�,�pb����҄�\�mܐ�g��g]-2��-e(�M����2b��a2����U3\���ѦQ,6�2h�Xk��sl�v�Զ(b		0��W�vh��]]I��c�]4m�:f�k,V�U�F�J�(�kM��-���
�er�Qe�:�멸z!c\G��Hyk|�%�Ÿ]�n�r=��a�Ԇf��Z�5�[z�jkmvbb� �D;���U��%��2����ͥ5M�к�5��hV)�҃*��
ܫ�-�Ρ�WE*A�m�T���Y�����S�ekq�),iI]l�Ն��Y�hi������ɪ�:I&�&,�V��S���#S��[V��ekŶ�lB�+`-c
�H5[b%��ŃR�Ł��+,�%m8c-�<M�X�rYmX��U��K�Z^Kz�R����<X�S�[*�ևZ,Z����Ye�(��T��[,�Е@��E�%H���VXEB�Q*0��������� �a��q�ga�M�KX�-�4)v�#)E�*�z��T���\N<K�e\Ḏ�99 �L(�J�Y� ���^럫2D����T+�IQ�B����s&4`6�~ �,�K9�)}�*�9u���@�{`O�q�$��̜ͨgL��ND��Ls\�%"HE����0�3+�^�Gb�y���nV��dC]B�J>��2IU2�lN�S�M�(DI���	H��8$�\z]l��,��A�s_�ns�hץQ��0�\�����a�2A	*�(8*�g�J���`�������QX7���k���~ �q�%9���{�}�����)��P	��&�eö�Hs�;Ke0�i�.[���f��}�X��$ ]"A���R(v���Du���ź�r�8��j�«2Q�"��� ���U@�R���֠�E�o���د�c�*w{䜬h�~�~�/�<M�=7/��
ϸۥ�>4m��p��2K��:SN����9~����9�֎c���1<�ep�� �?��ԖZ:�s''~��obA�d	*R����X�����]N9�U87���j~{ wt�%%?%>!(�E�FB�Kj5'\���'��䔊�M�Du���ź�r�>��D�R�.ou�
󾳐yʱ��Zs��м�'9R�IN�}�3r��\�O�0M���t{�\��lw�W9���"A	D���%C�37���k�%(�8����%�C)R�����A�0�^�f8	G	n,�$),���������(ؓ�����p��uT���#6�](=�w�j�Df�P�{z��Yi�DG3.��Q��p%�C0�b���}��f��,� �ȏ� -��C��Ē��t8��@�����wf�;�G����fL�UM�\��UMf�K�e ��/�w��|Ie�^��p>l��-��t�k�>|�^M;��ʼ�v ^CC��AY�Qv*�cS��v�e�*9��C�V��g��WS��EӡE��Ai�L��lͫ�K�p3jG��F<R�\lX�j���x	�QpfU�e�f\3/��s�~�{d�!����!�^w[���ڍ����z�x���`�1g���K��xz��L����ڎ��ښ8�����)+ʹ�<�qG)�]��[��;E��J�f\̣�{Z�ߒ������`o}A��k�|"�����Q�3F�ʸ�cL��_>���[���㏂5��K�V��x).c�_�x�C�"ڽ�fȖ�Kg��C�Yc8���^�a�e�*���3���E���m��w�x�Q�A3 �]"��}?��ڡ�`��L���@dYX�� nȐ����*���kq��[sG��s����v���&$��#ш\\�r,�a����ϸp����wMVeùWڌ�]= 1��9Þ�7CF��"p7�&�PlF�2����n�y����٣NeX!�	��3+��zZF���q���%����X2�\�u8%��v~���bb3)WJ���C�����gYv�k��,L�m�pa��t�����mCf�_�9￺���Hy����>|ҕNp��u���{OSÙt�-v^nͶ#���G2�1�L��h\�-��V:��_IB�C �s@{dH�U7�hӾ�·G���$��.��狎�|bz��@�JB|���v'�i��H-�Ry�`��z�s��oƄ}�-�J̽#3,�̨r�9�a{uw�֬C�O�Տ�O�'���j���݌����K�[ ���7eKN�362����̾��j�c!V���̩yK���[8��	m�۳����Ar����\R�Փ^�!95�2�b��_EƅYl(��[�ᔕ���W�����V����t����rM;|;�uH4�w�W#�Z��kKvA˞4��T�j����u�薪[��X������ YMe#�HV�0�cDwtXA$;�
:���kGR�)d��C�����]L��hԪ��U�l�;C�cmhT[�)u&A�2k�,�a4�XQ�î��3[(�kK�;'ZA0����p#�1i����x{@�� ͡M�
�e�n�Mm�{�O��[�]����i6uE��Z�!Yp�ڱ��=KI.Ÿ�����Ğ�C�������A�	.��"��K���P�i�����l�P��o@��e�*��˜�(�n��D	�~���!L[�==j���-;Q�A �c�ۮ����3�Lֶe�Нg>��̢�.%f^�-Y4~�ǽ�{;��v9vb����N���/{��9�X̢�33F�2�=�8�$�ŖK��8�#��W��H �F�����X��ӗ�����8~U25��
�7�\�}e�ʩ���̨`�����bc�k(Wâ���7*�g��̎`w]
;�����fF�Z�S�"̱@g�8!Fc`�v��p�A������1���6�KmZ�7��ϖh@�>|�>l	k��Y�m����`i�Y�Ɗ�ӻ��~�c32�s*ZcI���!9'w���:�p�o�7O�ׂ�w��Ezû���Y�����>_���.h˞-`�g�:2�N	��m㠶�F���o��&f'�O�#s*\�^g�;��}�z>��R��-+���]�v���`����2�f2�fhpT�{d����+���k��k�N�g��8�G��eX�Lffnh��>ŧx��<s'#�'����^�n�v�c���-���O'�Q];b���'�Q9�4hs*X�33S2���u��+zx,"��|�tNnY����	� K�7vl��#���ت�}@���1���T(൹�K�n�B�95:�����!�-C!�T�6շ�L����DL����c33G�c�]5�J+y��)YC�ض���Gb3���9W��ff�1̢Ĭ���ν_`;�5���j�NKҸV�[�O|AM)F�5�(�
m��jr��s*X�)�4hs*�bg=ފ��Ob�n�b�����΋�zdu!҈�°��[W����J)ڬF�-#0����`�o�NQR\��b�N�C����3{�[�dfo
� �} ���n�h�7<ݎ����c�o'> �H����B���	�WԢy8Mҕ���YB�]K�Ag�Vo�q�Bfe���Aa�*9�g^g���\��p*�;����ݎ덼�� ��5����?ݡ��w�g�A؏#*�jkYtnQ��Mq]]5�=sH�q
b2�rb��S��t�ˬJ���ѧ2�3��ZIt����+��37�|V78�B9���;=R�����t�f\틼�o��C0~odP���﨩��[����|~dG����Q݊�+�������~IB_;��~�Nf^�&e�#8$�k��w���6�v͛�a������r�����۱������P�D�!�@�����H��a��H=7��;#/z��	vkevPˋ|C$An���>z1q�O���D��ΡfJ��f������#��d�#%/@�6���/ݯ�uL�����9e>��=>9�'��2�ݠ�s2�����5J����:c�ĭ�tc�s���ϫ��R33�4eX�J|^�㼧�o������qv�9�C�A!�v�Ό��g��WL���M�U֔�ǹ�ߟ�?Y������D�֨��w7�ٺ���9q��߷��ez����,���353+�bP���Uu�Y؛U��|R���ÂI.�zn�\�Ef�Aj�T}wflv��6yJ���.��Ոg���Ɍ�C)7v�zf�-��͚POUu��뾳�}�u���xD�#�wF�ʸ��P��T	����� � {�`��jQ�MY�s����x�׳DA�J�#;/�Cg��9�b1Ĩ"ff�eU��5��0���� �#���Ď�Y�����Ɔ=��ʔ9�zFfY]�/�;�qooESˠ���1�ff�[�
�mvz 	lyб�(�ϕ�'_cm�x���Gף�֭�k����S�;?y��1ͳ?j�P)���i��YM���е�iX��h�!��م��u��Z0�P/-��<���2%���*��fz��e6FZ�ͨi�+Z��ps��2KA�0e.����Ψ�(e#kt�:�.*�J�5u�K6�J�]-�4+���5:�s�,�c\�R�
�:�br�B��az��, ���W���$b����G�R���[��-��v�F�IW^v`�Q�.�T�����u-�[[����T�g�����!u�� ��@�@�wv� �}�<����4�'YK#���c[��՗PE�7�+�$N�n�@�� $���J�����s@�����9Tݜ=�'��"�|~׳@�� �9[�j!@�����g\O�����49�,Gy����ٚ�t��s��v�n)�E^�ؠp � n��vD��>!��1�p�lm
ʝ!�	# �F��uӶ;j��G4�'YW��YF�m��
뽔^?!��kx0Js�A��5z:�N�u~���Ur���d�dY��׳D5H��3v�P�W�K�梜�~��H0P8Q	0 b�⨻D6�*WK�ˠ�:���M

]x��>z�Bz% ;]
;���"8p׺�I�Y��+��ޡ\��+�i�괠	��c��nȒ4�[S�&p�n�������5/<���M�/D����˽����W[��v��O]�7�ql;Fn����H4	��N�	DA[�F(vs2�倈-�:�Ъ휎i�R�c��>�u���6�~�b0������c�9�5� �ȞDH?"��]u1����]ѧ��<�^�s���fhәzavV;��U���ܯ�c> �t��ƥ��-�5��
��� �eM&�ϟT��=z�z�E���9��霚}Ց9?��_]�j�*��e6��-� ��A�~݌ ��E���&/��Q>���P�\ʲh�u�j����n��Jʖ��5���V4�+��x��X<>��2��=j2��{�Y<�G��	f�����>��ʨ���C�V�cQ0ַ�Vd�1H2�'�!�CKzt��,��j���{�\g��ֻ}ٝ�3*��yz3,�̪��p'����~u�;w^���F�{�u��I�L�}����C;.�Fx���1� ���˾˥O9�
8fx��]�=��76<����Q���^�RW�3n�V���S8��K��oA6ڻ�r��v^�hE����˕�#�c`�����ќ���X�bVC˻r4�qR�-S�:v��r�oy�v����pd�x6����sWn�ɭ/l|���|9u�!RY�r�4���Z�Κ�kS������M��ihQ1����T�<��S�w3s�wtS%���]&��+���<:���W��^��߽���+�������F�SH)��n�)�Fe��g�@g��,dE�@
��v��3��h%��Vw����5�{x��J�&z��`�*U>K�77�X��.1�vt�O�h�~؃}�a��[얜��^]�Y����\�]ۭf�;.����Ƙ��k���-.X�ND��yw�����[��j���҉�1˹ډ��TL�cA05T���qL��OLI>tȫ,沤�zx��=�
���������R=o�^)}��Mf"�1�-��m�nJŬ�ct�L�<���v��D�����_�����^%o��jf6��n��93[����EU��|i%��ˊ��^�ۊ�%�H=%�=�;�m�i@A��r����g�/+Ÿ�˷=�1ك���V�#!���M���~&��7�������#ݿX�{W���eT�.��/5lk�v�0wc�"�w�b&!�K#�<3��]#�f���Ld�W'�w��wt՝��`b�� ��֍��֋Q���65�RF����,Z5�m6��l�QQ��բ�b��UF�6E�60[%F��
�����(�F�6"�"*-�QF�dűlQ�[h�LcTj5��Z�E��QRh-��Q��#Q�@RH�
��w9�Z渿w�{��~�(@�(���I ��I ��sچ���r�I�) �S)yP) ��,>#���������tk�~���߀֨���!I~��R�)��r�ld���s�i ������z�s�>��V��=H+��I'�!L;�\4ɱ��P3����w��k��ǒ
AH+ʁI �*�vᴂ�`R9E��
H,��O*�(X��
9�jH,69�-#�����[?]p>H)�U 	=G���J���^�$|	�M��i!AT�E����v�RAK@��.f�JH(��_���LH���El͘�pI�3���*h��,��[�eƦl����u�%��X�S�O���
H)?ü�p�&�RA@�~�I���
�X]R@�����'�޼u2���z�� �Qi�@��������>��ϻ�d�T
C�JH,*k3P�AH(�E��
H,�2���.D��Ü��I �s�ZARAS��V4?f����@���)��ˆ��JH|@}���^q���������WT��RR���p�AH(��AH)yP7�g���{�� �C��m ��
@��Zi�)�����%$9�jH,60�r�I�B�
A^T
@�/|�{�qE��(=�u+,��	���i!EP��R
AtWn$��L9�\4ͲRAB��(�Aa�aI�P[
H)(�����_��֯�0��p�&2�
�4�Xi ���r���h�$��d|	�_������;����@���) ��T ���8j���y�5ơ��wXioP���їJ#^����w�x���(�h�xz�����}r4�j[K&����������W�0Ε\{[u�u ��?~��i
H,�2��
@���Ü�ݤ�B�r�H) ����R�0�9p�!���>���>��~�i�o|>���}x��#���a��!`��A��� W�z���H;�*D�Ъ	P����᎔Ϊr �lLk��pۜ)�n���4��I���-? RAe��`R$��§���`9�-&����C)��:g?s߯Z�Ͼy�xR�������{�uu���������������ü��L�2RAB�9�4�Xj0����RP!L9�\4ɶRA@�}���>��}�I�����`X]R��#�K���9�^�gu0��	$���%?��Ĕ�XQ������l)���e`w������B�&�N0) ��X|� �*U���uD) �9P- ��Ss�3`�I
�s�i �ߓ���"�`�7y�빻�h�}F�/|$��4~�
Aa���O�) �Q�Y���R��)��9ˆ���H��) �5�����S㟯�/�
C�JH,+~�P�Aa���������L��
@��=�W����Y\����R���i!U@{�ZA�D) �GNU�-�v��א1 �P)�s�3l��P��$�) �B�����0�9p�&�I��4�XH/�Oo{�����높��}���]W|~���s�~��r�O�$S%?��Ĕ�Xg=p�AH(��"�Y)��H�K:��ʬ5��9��c_���ヸ�'�(��۪NiKL�#C��kF���1jx���oܧ�n��4���������khR+驮9�slt)%�c�j��Q���,���.c� [u�X���)V�����6�7nkY�b��`
B[p���BP�GF�R٤&��Iw{WD��@��9�F��U�&lƼ&�Z4شnY�e֖�9��%dZ���$�SW�TV��܊�����aZ�� (�Ԛ[�b[H�5Ш^�z�9y�����eZ�b�Zv�l?I��[�-�pK��Ћ�m�.��䌤�es���*��tֵI�*�(�i�8�Xw9a����P;��H:��Z�� ��
a�r�n2RAB��H,(c^.�n��޿Q�k�	#�MD��	&��+�~��a��놙22�
{�i �4�A}Uʢ
A���rᴂ�`R9E���FJyUBĔ�X{������[s��u ��3�ZM!I ����_�:�'^��Y�/x>�&�@�6G��T�E���]v��R�
a�r�e{�?w{���>H(��H,:0���,aI%!L;��2l����A�Y����i ���eQ �C9ˆ��kY����}����A_�,�oLsU:�-{�0�9@�>�Y���U@P���XQ�wP�Aa�9�-&�
H,�2�U@P.	I�3����j��X���E�Q
H-��),@��\4��JH(��X~����{��������硤��?) ��)�;�ᤂ�P?s�ۯ��^�g����AH)�T��
A��{��c�9�-4�I��O*�(\II�9�Ci��R9E�kg���������������V�+�|��}�ô����=�- �RAh�����
a�r�m��
�9F��s���3g<[��qO��
��dN�pY��M5���s�4*������ƯT�Z�) ��х$��0�~�i�c) �Q�٤���I�T� ��s��m ���x����W{�g3�y� {�ZAH,�G���z����q�UC�JH,+�桴��`=�-&����C)�T�RAa�r�c���P9�- ���U��t^�خ۪���W�����e�I�tܛ��m�h����w�Io�,�3{�3�|v�s;� ��_j��������� Ss�3c%$��H,5f~����}������4�]U��R���L�e$z�H,4�^U@��z=��)�{����
@�Qi�@��ʌ�����%$s��6�XlaH��Q
H,�O"> ���]�E��^
���R|	 ��۰�� �*�ܢ���$�wH)b0�9p�6�I
C��I��
H/*�)'�r������u���2le$
�Y����i ���uD�Us���yN"_w��7��+����� RAe����Rk��;��u���k�6�XtaH��HRAd�S�
Ĥ�Ü��i!U@s�ZAH)�T ��)�9ˆ����V~�$R
��i �ў�*�{���Y��㹜�$UA�0���X{��d��H(��X�ʨURs��������>/�ߞ�K)�Ÿ�6ԳG@F#v��Y��j�k�5a�
�%"݆=m]��d��6~�
H,����@R
Aa�}p�AH(��R'O*�(~�9��}�Ω�|}�~�)�����v�RC���wU�_Ύ�Qi(�$�P��)��놙��I
�s�i ��RAyT) ��
a�r�M�RA@Mz��;^��ף�$����ʢ
A�T3�����&ǽ�9����n�16W��O�$S%>���bJH,3ݸi �r�Iw߾��o�s�>�O̧*�(��Xk�\4�R��(���R�]�R
Z0�9p�7) �Hs�i ��{?~����gy��:���u�гv�*v�d���ݜoz�/������O����3�|���D�
5z̳���<OG�)Σ0� �PL�u~ ��p���Z�w3��i ���
@j>���#9�,N5���@�U�xr�ݷ~����% A�
�I�@�dnpO�f��b�p=����&�����Nh��\LeG3/H��.&>���>��쯴�&���h���7�<�f��wő5B�݉�K7\�%е�!���f�\h�k�ѢG ��A�#eJ�R���U��XZT�����ߏ�7{�F�>�K�߷B۲;t�����4�K�R$���1q��У�\�r$�|~;�B�;� N�Mf뻊�����";21��xٜ��9���5=�\D�J�f]Ws[ӽ������M���v�a�������2zj3��M��7n�0��{9f�2�q(L�Ѣ������m˺֨��T��r�e������:�g�K��BOOwM|F*B��s~z�៚�t2~���r��8�V@���Օ�*�N�m�D�D]�o�82&�;<-p��E�%kb��E{{�5����w�^|.���$!��<�bs��r��
0�mxť����^y1�n~c{���p����3�_v��Gwg����~Kc�>�OE�m���-�s
µ#�\%�[�Y�Z�Z�.!�\�ˠd�l�67��q-s��>#H��)w^��]F���a�����4�̉:D�n\���2����"8�3541̢��٦�;��w0SsD�J�5��>�\u次'� ��3�H#O��OvdݝwY5=��g��JFff�e\Dq+.��ۣ�еÆ��f'��w¾� �jS���3(�ƒ�N�o���;���W a�~;�B��ק,�}���|�3�C9�_��6�������Me��iŘ0S��mL ��)��v_���Oܙ��s�U�׺����⻥���e�Ւ��a��zc��/��g�+[���Y=)����?~;���y2(W�b��"&{֛��G5֗�|9;3
�T<�V�ϋ�}������+�*�}c3Q�7b9K�����l��k����UQ�"�@��Mt�c�*�֙�,�[]-��
¶m�h�:�����m�u��ViT�+��&0�0���o%��.�"GG^t�BYd %���"R-��v0�e.ĠFM�J �fW9Hٺ�M�3D���(��Q[�gv�k���7j���JE;0��0`�X�uh[	����-er�����~��/��Ը Q�f��sCm���V�6�2�����
�UwZDV�u�_��Bw�\̯�WY3�&8j
�b�7�� j�WD|$�=ܞ`�����8-���n�N�;�k�(�>���Я�u�O�T�,K�m�0 b��݊�3GU��쨐�V��"S7�nh^�"�S���s,ރ6��s�p;�t�v�J���S��#>��3*���5ʰN��=�V��s���F}��Ӟ����MsYVg9�Ơ�fo};<{`9?:J*�F��e��3*���Й�\fp�l��@MȻ�Gr��ʪR�\n8A��}�A#N]�t��[�i�����3ŵsusk���l��	q�R����vA��
[k5n��-0��gG���#�fe��,�|j��;yU�皪����
�j�zzt��񜪎fhәV�cQ;��}����9F�:h����k��:(�jH!��:o;ry��P��N�
�켭�8"^EΈ��3�%䌦�܉4��&.�^���}�Oh��A!�Q�	y�F��o|�=�(��S���;y�/7Y�߻�x鼲�=E�v�.�����Mo���˕u��We0�m��L6�;�! �ޯ�c'H�7v�
+��ު���D �}� �7db�2͠��ٖ�]P��A��F�)�j���[p"�c��eZ.%#�����������"&��m��A^���+xP ���?��<2Շg�|k���?�ظ��!��aA܅���֥�qVZ2��ݪ\7�ZV�4��n���ꮍ'Y�w�ޑ9�,���\��d1�v�1.�G���r��]��]�q��8��h��Bff��P���v�J���ѿH3�4!)�GM���+=k]H����4?gH�4�5��:���_h��VΥDffhәV�Fr�p7��Tw��pcGb��B#�r��\(��ӝr�l6jqigFB�ܧJ��.�˾���:T��9Ȳv��vv��R4#N�nc����|3K薗p�Cowg���P ���͚ �ȟ��gL�<��y�,o�I@�ݡ\����v�����/)��~3�+�f[u���CS�m��"4��|���!8��ɾZ�D���sD�t�#L���
���]�!Đ@���Z��݌�S��h���bm�Xd�x�7j]��j���+�� �(G��ʱ�\i����6�v{�W�.���;;���u�>�P�ܽ#3,�Ƒs2��W���z�!,��#L����|���n8�[W��pkn8�
"  ���}��Sԯ{[����i�Cͪ�A8pYW��Vzbf^%:?;��܊���Vf=Nc���S@���Gۻ?n��J��T���{�یL�yc�졁\i��o�꣹�}�R�@��Hʦ7C��F9��3�FN����6�5� ëd����8�e�oo���!�wOd�fL�Uo��*�=7�E�=7�T��@���{�Љ��lʩ���7dI�n���ٝ�f�}#[�ܳ�3��m�Z�Ln�p # �3:�ؐAi��v��7���jc� ��?XY·&$%�u� ���mD��vi]��,	f%������Ë�A,����Fv��Ņ�Y*�5x�~���y�o3�����\gjTffW۱�F� ��p����A�}��q$�f�'S}GUͬ流P?�Dz�̿��=k��]��X̪{y|�X����e��w�	����� 䗌⹬[��ˏ��`�3��ؒ�i�7v���x��V���ő5�ջ!�����X*�`�= ��?0��_����׳gFz���{�C�V�cBnУ�;�oyտ��;Q-7�a#>����ߦ�>�,FR�̽��W���ɂ	��6PV�sf����e��7ri#��C�=��3I��{����^�WW�T����+�u�b[�Te@���loO�e9}j�t��%�M���͘K4�.ntk�Y���N˝"��T�֖P��#GN؉��l�>'w,�#��W7wy.�u�z��.gV$
�2&N���.�!6�cH��odoX�6�1[��M`�ַ���Y�?;n�{�Ԯ�F���R��=�.\�J�aU����ld��h�F#6��Q35-�J��eH�v۫71�%��!�m�!l?7�3ݴb�{��<Nԯ�1У�����	
���@���{�ڥ㇫�	��|���~׸�����p0���K��nC�5^����z=�=�m��C��{��n�i|$�;�
��O��3{4���>0(�緰H4�1�r�E`X��R�8�y(�7����o��q����G�:fN���ӓ8�ۄ�}ݰ>��[�;�"O�3�7�0�����o1ǧ,�|�{�x���g:�t��w�f!����t�e{�HQq뺉mۙ�DV���,�lJP�	�V#q��/gj�hRm�$���|�s"��[�����k�p/n�n�efo�w�8q/�!t���ܳP2��{8�<��=t��[��s�S��s���Oz��8}V{����=ï�k��@�^ٽ��Bpk����]��y��8'����}���k��9�۝�;ݚ�~9v�{�F�=T�#���)�@��M�o*%C
�>�:2�\�a�s�c��[ᯩ��Ea��ȋ��F��lDmh6LV�1Dj-�؍�Z��lUF�Z4� �5-�QF�Vƨ��F��cm�[ETj�[�Z-���Eڋd�%�Ѷ"�#� )IĀ-"�J��s{(�gF#��X�uv�ґ3ĪئΤ�ae�R,U"���6�&�eG�f��$��Z������3a-�\ب�Qڭ�TX��v����V�����PҰn��0����L3�P��F�t
�cJ��$#���A�׊�r�f�,� ;m*��[�:��h��b���:��+��6�:W.��j�8r�4Κ��#GA��2��fсN;f:˶]�M�mN�2�0�˰��
遶&���!��s�bi���0�,��$��@����EM,
� j���S]�Z`.�M��/7hƹJhb�nz�L�6�Ŵ�:D���m��F���, �L�4�+0i�ւ�cc]@�f���4�AiY�X����m13qnCW���9f���9�nFQƷj���)�ԕ�V3LgRR6D�]���ul�HL�ka�m]1M6��ґ�\�*��^��vA����v�Е���$�3�Tf�B���a�f=A�R�͍�X�J,��*d�Usv��V�\LSؖcf�`hh���;��ݥ�*T�k	�l�s���@��cW���F�1l���A���hX+.%̥0ISD�iTq�(�xF�/9��YF͛��VhL	JY���x]5ķ.4���FKq�iq�����	F���!.�H�b�ծ4�]V�Ye���A�L긡lX1��4k�V��b��j��H�.�ֵf�t���s���VY��C��;T�cB��B3]]��XR���f�'�,�j�e��.����H_�'R�vc������덇U��3Y[�sn�h�f:f%�1٠�6.�l�����M����f�
��dM�ڢ7��6��"En�Y�U(�E%:i]	au�f(��N!��Ņ�DtK.ʹ��M������In���b��-NKV���\�0�ձXkF��a�jL��V�
bV���\e{A�R�)����pަm�uA�V��AD*L2U�kv&�5Va��@��j�n���]���s\���_�N��N�={���}���(Tx2й6��/X�mPv.p��ı�n�p�X؍���1��.���2 ��%��፞I�uM	�gUQH�ֳIL����쐔�m��Kn����yh��ڣy-���M����ada����vє{�����Ո�-ɣ���\D�6� ٌ
GJ�Zk�v k���0&�nR����f�6V&*ib�u�\.���O��������hJհ��$c���cY�&K�%L���č4�V]��}�^�s�[2��fh篲9��W5�q��q�nD]��n�G��E|Z� i�wn�݁ ���^��y[�T8?f�����b��}���K��}B9�^�'޲�3=��Nf��;�������B&fh��U��?{��e��1��"e`�����({`H#ڔ9�zD̲��ϵ�ִ����TF� �;�O�q76�w��t��g2�"�Yq��/:���_eX#�	��3(�"eJ�fYܪ힫�l�K���"~������ĸ��g�B?z�1���5�ߵ�����.�J��m�Un�K�v#�V훰2����hh0zۦ�V(�������s��C�V���8��f����Fu���g'P�p#H�l� i�	���d��1>�s:N��P�gtS�Ս�^v��v���I�?�$�ǘ[����'�����.V�]��o\l[ֺY`ҩ�&F�]���X<�%"��{!vs&�b��s.>��A�Я��S��Q�l�|�ā��} H���٢ݑ�t����q\n�;tbm(]�"�Rl��z?g�j{,�ƙ��i̩c�o睻��g���E�����m�xT��f. ��s�I<��d�c��_T�1)���Y`�Ј�e��>��^�s���.[3[�	Юu�n9��T�ip˸�/��7�Ѩ�U�.%}��﷙��l��xɭ���N(���PлGcFW;�(��Y�뀫s\c"���	<l�������G����0+�bV�Oe��Z�?��D���׽w�Y�}��'ݲ�c33F�̠��?�[Ҝp�.�q��8�	m�xT���&K�{`IA���ͻkL��P[95�,O�#�ܽ"fYi�T���ē��͎�5�w1�+7N���=��<�~�\�%U�0�r��I�`�T���������Euf��ȋ��(m���|>�
��|-#3{[گ�����y���y��_�4&fjh�λZ���ea��TL�����\������W��0} �[�@�\���%'�V�B�~��W�l~8Dy�(3���`�p����:��b�33��az�(:�9�zD̳[��}����j�U
�QR��t�Ä� l��M�`m9���l%�A�R�.�_�Ѵ�Ȉ�r��l���fm
�8��1;���8e�qhՐ����b!���G��f%D��h\�w�՘Y��-}��s@�����3��.A^j��g�'{&� ���[�n�XR�~ѧ���#33F�ʱ���e �C�Ǟ$�N��}�������ʟ�����w��f�:���{ �~!�?ݡ_.�+n4;���8e�q����뉪��́uz�RBZUd�^T�L4�������5ю�hO%����]�b�i�7f�8à��xw}���	 ������\DO4&fkB-9�~�mB���x��nU����|�
�W���D�~��>;�Au[uHЉՒ�J뙟�����ĩ`ǭ�."�Y�2A4�0�uN�е�;�m��tO�c�@ؒ���\����̌��{Fy-��7Η^ֵM��c�}�^цe�̠�̹xv��3�wn��1�;��]��+�(O)ի3��G|@��["���l�uu���Ki9�hЏ9E�G��-Y���ƞ�g�ӹ���y��}�������I���1��̳Ne\NfW;[<5�kկ����z4?z�D��}�P}}7���}�����߸�>�R_ީ����Gܰ�Q���DnȐF�a'lhϷ�{B�gJB����mTq��wb~ �!>�p�<X��@Fp=�r����{7�:���V�h(���9F�Q,!��P`�]Ōj�+�T(�YBq�u���q��CO&��uZ����~�|��(hQ�\��ͮ��/�&�u���:��k3ʍt�i46ueË2^ٕ!���e��+�+��Tk������+��u���MGJ;�<� ���q`Q!���� �4��-��E��v4ҴЉ��iJ�i1�Ԧ6�h���́u���e��e3��cQ�m�������-�=���j�ڝl\l����Qvڎ�ݳ�XU�pO���7��̦�T1̲��L�汚�LME��l��Z�C��Ոފ�5��}E�ڔ�e�G2��v��y���98_#����D.���������D��Zq��34j9�.8�����.Ԭa�<ϯaJ"�Ġ�"��kS���ǜ.>���H�:e�Z֊���n'P�ݽ�s,�1
����G4^�"�6�E�(YKRWlmT}��`��Ne�[V=������k�!@���
�5��+���x!,�*�p�G� ����)b-�X��5O$iF_y}i�
3%�4ZQ�}��!j�4�w�E�T������y�������`�W���f�L��� ��r,Im��-��cL����a.Z�	�9Z�3smŃ䒁�t��5����
]p{��Z�Rࢣ���*���gR��K�,~�׌_��2ڳpZq`ɣ�n�ô}{��Qd�k8a����}�ķe�L��w��M�9,*��kzp���E<ػ��N�)N]�{��x}�  9��o� ��M>Aǻo#
�N�� ?'���<�����׎r5�7��}}���>�&fY�̫EĽ9�yܘj3)��Ml�Wiڟ�����~q�f\̣��/oyMw���؏ܲ�Fۻ"�\壠FrĪ�'�/�_!Gd��"�� {bA� ��X����[W�hu���&~�c���_Io#
�NW��Ƴ�� �r'�4���^o�#�����_����������L��m+[+	L@KG���!l�ګF�Gif]H�]O<B��4hs*�1��w�8�v�]�<���b�&9;�w��`�8��~8;�1�Ոe`������<x� 4�Rw����*�eEG<D
�B�݋��jDLF�H�T(p$��n��&L��k3�����mr��W�������8baZ7�nA�Z��ƻ���n��0��̫�����\E!�O;;�Ц1|>����E��=ْbr�G����������}mxť`�^�3���D2�T(���H�\�}qA��zZ���y��~ �(�SY\ �/����u8�Q���b��k}�wN��Y��W�پ/�嚦�� �0A�
v$����!��F� ��e���\]��ѻaa�!�6�smE�Sl¹s1.]Qr�l�{顏;E�%G3/I�E�%���$.�� �@���芣v63^����5Q&fjfWȸ���e���كJؐA<Dr���T᧧\�o:��.>�����jR2��Č�"A��'�<���C(#�מ������r���9�%���.&8~����X"8�&fY�\��u�����Q�B��/�h�쉥�L7'�<��5���M_M5�j�Y�隭Y�l8�ǫ��nJYԸdŘi�"�S"�l���녞��qtE���9��d˩�/���wwφ� �Nsg�|�1���Ai�|(�2ڱ�L�O�@��{���F��Ȏǭ�sg�������ǜ,�E�?�Vm��K'R@H�)����n�����^*WM
cP�.�9�؛��_���=������Ov�Li�fh׻��o�窶�fĮe�GЦ�i����ȿ� ���(�?!F���<Ӌᑢ�	o�$��#vD���15����< ���D��}Q�NX�5�]��U��p���mxť|0
1��5�<�;{j�Q�:�~�;=*^��L�� ��N2�3/H�Xc5\�5�UW=�?U� ��8����Ю���t\��إ̸���d
�ڽS���[%�7v���Ne1m[���Sս�x���A=��9������xw�B'ܲ�1��k��kެ�Wv�X���*�����c`���/~ བq��t����� ��6$F�� ��l�~�̟{������I;���	�����3j"���S�^	��j�v��5���ԕr�S�u��9ͳ7�Ѧ�����/8��h&�
A9�̅7f���u��F�ؒ҅xR�̐��֗f����ح\���I��%�)*Y��[����	f�8N�#�����m����Kiv^v��G6�H��Jl�s�3G$��\��ed,��W!g��ʲ�	������v��R��2�/������0�c�`���^a�\L��q�����p�����F�2�F8��o٫;����ʞg�����۬��s.q���@ݑ �0 ���#2�հ���c����P��OVoD��㹱K�p�߳��=+ǂ��O^��ܧ(��&��н���s2��e��[su����o��X�Ae#oKߑ�A���X�e��k�-+�3˪���b!��^W۱�N��mT�A��:�8��8W��H?`�_EDF���~��"H� E�˚̲�k��s:w�sW�;gkL�g`�إ̸��	d@!�Ƞwa����u���ƾ�_,M�&����b��SW[*."9�L��(��2m����}�E�ڕ#��5�e��쥮c�u����=_#�5s�k�b�D���ݑ@�ĐN��]���F��t*���n<�%W&_�ۛ�#_�X0uF�yW�F�b�K��m�����Ѝg��3̍�ïĂ����\LUd����Vѧ?��|���-G��D@u{�"��mG;��s���E�̩Nf^QY�z�޹�t6}�	�*=�nh3,�1�����O����r���C�%���=�sb�2���DG�Zg��0��k���(�G�`g�3���wd;{��ܮ.�=-}���] Z[���S�L&4��Gi_
3�mxŦzU:�����/�y��HŇLp��q��p�A��`������-9���?C�v��V����=��T��3j�8���쭆��&-Z���uq�p:�5���0��W�/|����K,����L|~#shWʲ;����[��2����ݽ��
�b�<2��?����Q�nȿ�� q�^U�eJqȐv���;�D�5��� �� ��Ӿ��x٭ަ�j}��z����Lʟ:F|����a�j�EF�?,�TV������(�GycZ���朮��w=��hRԞ^ C����p��������J��q�s&���WV���/��E�'�U��W�ko#&�=�bH�|x�H���ɥ���l0�=�A:2���R�������~��Tx�:��(�z��zBt�]�k�v��ջ�ғ.��d�r�~�8�nh34������5Fҗ���L�7����L��"2��*=����/]E>��nEw7;͙x���=Ϭ��y�4c�W.�n�Ｓ������z0y���7N�@����q׶�\���v��/b�|nY�(�J���VP���L�������$^ն0-8��(7���/�I���+#����4koZSP��/Y��3h�uK�`�愱��Vm��|�g��Ϲ ���;�D<�B���Q}WO<K�j���~ݛʈ"zA�"��ҏw^3ۍ���#���W�AŦ[f�i�(>��u}f�8�&`͂�v�������p����8.��ڋ�*�	���.��d�ybԩڵ�0���*�bkfh+�JG7�[n<ހ�*��������伦�q}f�=�L�u�� ���o��^���{�#��د<��}�g~����^�nj���U�g"�Q�V0����8�A�hc�WzH��ӓ��]��~�Q��������:;��X90x�>�:�{;f�,�-�&�{���O�U�s���=�a<�Yv<)�-�7N!q%��������}��/�wF1TF��[Tm���nm�����Zƣ5�j-Qj5nmͭ��"�#F�V�Z�I�1�Ѷŷ7(�E�-E�j5�Qhح��&�\��W-�(ڃ�mssZ���k���j��jp͉}ǢS����{��	 ��2ڷ�ՈeV����`��! �`�@���؏\�h��K�F��G�C7ߏf�ߴdw�K�Q>�֦S�>)�ඪ��k�԰�ɧ?v�6��|�>:gy1�#����YbcC����{?^��s���8�Z��VSu[uIy�X���Ip�%��pJ��$�Z�BC�A�J�؟��D7x�;r[��)���}C�l��uA�H��-�~ ����oBfQbcL���O��VsVi���?J���ك��h����f��?2 ���W�v$C�e9Q��T4���[��ʔ�e�FfY���[o���Ur�s���w�����=�ޠ��e�4�̳C��l��2aX"�eE�G�kR(�t�׈�7�%;��o�q�a~��?��Ww��#r���V���,�+��DF�Q�5�O5Pba'l�nV�(a����P��W�Q����w�jL���34�\T�o��|/�럫�RX��33.h̰��ky��}O�>5�����Y�{Df��3qd@#1Ƞwa`������~�m��`�1q8sY(�t1�vq Ԏ�M�MaU��*�p�V6�v�e�ْn���!���T}wf�#vD�hDd.+���6�O�:d�jw"�h�}�ӭ��4eX"8�#��c^�fef��U}��H�w��wu0��Fӻ�f��-��F�7vmc�p&�*����ZՖ	Ƣ1ϽzG2�ffh���PN�;ݰ��}Zo9�L�pX���<��JQ�e�g�y?;�j��|Ev>��74F�	z�1�q\2�!�����ՓD�d��O*$Y`�[t���F���玤���`�׻������m;��k�� l}ݚ `�cΝ��Ӻ��y~��f���Rz!s�Vh6��r[{�Uo={�!Ղ���6���m�I-� �L��͞\���ў�:�P�*������� >�}���j���c���n��vʹ�j��hE��Ie����<��ݩ����t��c6�[�L���K+�Na.l��h]n�����X$Hk�fge�#�ⴛJ��Kj5@8��A�RSL5�Ddpͣ��\if�,��+�@ qC\g�
=f�n���[�0ڔt��5ôs�0Ń��P��ܲ�SkJ��e�߿�`ŧ4�W:V�m4�[V�n��H��J��l�ZH�ZW����_����w���`�0����(]���@}����
S3E&�5{�F��?^�
��'R���2�O�}y�����,w�^�/dO�y��B�v�l9_i���ٯ�?n�b�]TY�����E��K";�B�����٢����Eͣ�����
��̽{B��Z9A���L�t�u��}s"6�lo$4~?n�
l;΀�	��
S3%�_5ee4��w:��.=JL̳@�Qb9R�3.�~�u&����3����5s�7R����ۗ���ZcC���j���|��n�Cu��,*Sl+�i������:��+rJ4c���;UKU�e����v":J��=�NeZ.'�ߕT�75��9.�����9�P����ԧ��Ќ3,�Lj��r�_v/�I��Di��l�$���-=M��,v����4N�cQt�=:����[2k/i1c�e�82$N�#�:��Is����@#�~|�U���3;����f8Ad@#qȠw`��|��k|x}�c�TM���C��T�wv~݁�X%^,
��:x��}M:j����}�^�3,1�34i̫O�g;��||����6���Yp}걟%������M��w�K-@�~�p�hy8�ݹ�ܲ�Ɔfe�G2��{��fPӓ�)T*��^tq����S3�"=J���u3*|�}�k������v^����l5`�vr��(��2SSvF9��f�j�-,�fT�7r}��[��?^$���t��ȗu����I�RFF@ʘ����������!���c��0 Fj�-���m�ȓ�:���swJ��:����_s�?~���͈���Ns�߫��Ybc*=��3(�LB�v�fQ-�)�Vrd=E�8���ڱ;�S�<���yd�H3c+�m=��1t��s�gڴ�=����8�1b��m=!����d��:K������6�;��Nqݭ��1 �x� �[B�݋��%&fh���m|���j�TX�r>���#v���&�-]v�z����׳@��Rұ�� F?�
��ĐA���x-&?�un�ܺ;��#���
��˹�㮮�ɮ�O8A�c�wf�2Վl�:l��s�f�e5���1� ��,p7i�E��G���.xB�%�"�m0�D���AMM�~#L��СW(=�bpv�o3Y��xѪm�nQ�w�D|A��)��h��flЎe����gv�`�[���H�X87��W;��o@'�M�e�Fff�4�lޫ�5����jZc3*��FF�
OW��i����5[ޯ�{�^�h`��Z#�C���̢�2���|{Tø�;s���~g���W,v�8;v�����p �8�q�m�cP~��S�"Z~G�(�����Ӯv�j7�lkV��צ�3�訁;N�X�5���X`{���y/,�k��@���﫨��ff�S2�\J͚^žv�>�nD��ǰ�{����q��}ԧ������*ꧩr�ְ�~�I���B�H�b����%�\�M�F&�شR��j�k4�j����@��\̯����M�m:������9�P�;����]��}�6����"fYi��wf�ze���ɫtM08�΄�C��`�ٷ��:����P�wcMؑ6{7����7�P �$6>��������|�ݢ�)�ΑX��g�y�"�]���ZcL��4-+bef�w�����A�Ҽx;�P#��d��q�;ݰ����_w@��Sl�;�o��T}�ޑ笴Ƒ�f^�s$H#LTB�`8l�֋���ˡU���3=׷�n���s�ѡ̫G���'𿚼־���:B_��lhҨlf;u	^+�`�w!�L�Ź�c-��W�����no,��x�l�'z{�ᩤ�#|��$�5!��j(I��`�Dj�v.-��n1xE���9���e�)����^
��@�]��l���;M�4&H�3"
7um��J��JX-��Cb��\Ac��Ճ��x�����bP���E�Jlu-r:���Dڈh]��IW]"�G�.
MW7���h�uZ7�a�Y�ca�2�H�TśFmZ&�W���a�hE�c�~���a�'�1e��#r�Զ0c��[�ձ�et�U�2�0�Ұv-�g��z�t	����d�"rm�L��vw���i�rzNp�gj��81W*Q�-1��33S2�q)/��V��w�Ӱ�k��}'��.������n���g�ޢ�r�9�w�y_{/�>�.'Y@�T�-X�Pp|2������]N�ͯ0�^��.S3A��5*wc�H�2��Mf�}�ѹ�s�?��'�ݑ�|�1���vu�ˁ������u�����~��O����F�ʸ��ImXŧ��3���e&a��y���P�=�:�N��_w@��?l}ݟ�vBξ�z�l�z�A�,~m J(ac\�6�.ű�� ���GF"	�XE9�.�_�՘���B�ܐy�h���(Lxf.�=�����"�b´��rmX$�F��@:D7v��~;�$�uh8f���S�H�8�g�g|s����D�ʡ�N�S�ы ɔ�93C ^R��V�jV��u�����ۣ��ǌ��1�0�x����/.k�7`]�J��h�ݛl�p4�~���~�+��o�r�9�G�ލ9W�Y��NeZ.&_y����e���f��U�Z�"�z�=�$~��>;�4݁$i�-����"#{���"A����
�B��v_DV�pn[��d8<��O9�]��wbA������i�YO��m_��mH~>��{�?2;�=�s�ѻ�m��?u9�A͑ ����O��g?m��[(�f�05�jj�,��s��in�@%��e���"s�ѧ2�ĩ�Z߽��c:j9�:Ff��Wq��Y]5�j�~��G2�LeG3/IGk[�s��ڝ|���i�э�a�Nf;�	� q*�݈\	�u�W# �ͪ{��0}O�0[Si��
�˺W���<��'�_�/�~~�C�{�J)'0�l_�)��M�W�P�w=����o.+-BRZؤ#�����.;b˝W��7���Q����.=��9�3`I`�mX���o��K�Y4fyuz��
2�y��$<��������	 ��޺��/|��=�פO��D̽#�ݑ �#;��aG�"�?:����oqS��ׅ7N�8O �%B�݉ ��/��*?\�?}�mH4���Xq�R��ֺ"gB2�8��j�T3k�-����T�.���w����ݚ�u�Vu�u�ڼb[!�����S�7��y[�s�I�����(�Ă	�0cE8[�p�4iN DPA��O�#'�9�36G�H��ݝ"���~u��A�� ����j��@�7v�N�1զ"��Q�·1�JN�Tp �"��c"����l�P�>�׎ u@+:k�7`e�Ʊ��nm��%�� ���p��Rʫ�='�!umm[8�(E7�X�ܱ�b}�<B��ׁ�ոϫg��)�{���zz8���!f�A�i��g7�}\�3���49�b)�DffkI�guPG�nb'?Z��袾�4d����ߎba�mO�՝e�F�k��v��xS�6R&1�<d�S@��:	�,vt��ѠjWu�kCMD1�K�>C�߹!���i��v�BiB�c�!��J[����$+;*"�B�J$�t� �ݡ@�� 7՚�8�g��)�["~ˣ�뭬��Y|%��	U�@Fl����h���W��rͼ�[:�3,әR�N:��NS�*��Oi�#��?&2�̽DO����g=zu��wܺ�O�"@!7vE�)b��:"9��Q�F�Ã.���\�yU���e�^i�0S�m]�����|�ft���{k;meg
l�=�⫦�#v@���Z����~iy�%��鿢W5{�%��La`��m�v1L1�V�dQ|�}aU0N�w�}2�y�o_c��Q�&������m͂z���&0��]}��QY���k��7'�pK�"���H�E���y4hMBj6z��L[�l̳��{�JASs�zr�>&���/�6��?j��ۻ`ýoE���K�Osj��:=���鄱��+n/���n-��b&��	Q7"]	I����3P�fa�Ww.k����-�a���*����v��?q��Rߞ�H�iΖ�`\;r�rw=�4(���^��壒���A�wc��ps����k��+3"Rb���P��3"l��ȸ�%\^s��wR��	{����{���w/������*�a�P#�3��^��i�љ��Ē��|4�^��ۯ���n�Һn��=Kg{�΢��m&a��0=�t}�S�7j�Vq��CB�T��bBݖ�X���9�� nmƷ�*��&���o��x��{Ţ`z��JI�*�*��wJ6Um	�鑸cgI6D���uY�w6ZAƹٍ,�k�kl7�O��q��Dn�zkm��^���i�qI�o���=�H����]7�0+�[�v�i"4	��ד+g�}RO|9������cj�n��X����7�.IOv^袭���NX�X��`p�@���*�m�%�⫧(�����G�e9ʺBmsr�؇^���h^���GU�tk������87����v���Ԉ�9l]��^SѤ��)(?m3���	8�gb���`@�!H���\�.m\��V+Th�EZ�j�-�6��lZ6��kEU�k��5cj屵&�hɪ��QW-E��ch�t[;�6��r+b�
1ccE���n�k���7s�t�q��e0Tt���,oc��b=�Me�I�)�F�v�
P1���.����t
�Km��9f.�ۀl�&�Bf�h���-�EŊ�dly�� L��m.u�42�(i*0s�r�i��mm�DnB�W7&&%���q��&!�h�#���֔��B�Ժ`���L�%�+frJ67%��L��*m��5�E5Z�Zg;TjPeLDƪVa�8.�W6���s����%�ZK�0F�u��p�Z�k,��ԛ3e�j�����e�FZ\Yx8�t�/1��ܨ�PK�G)Z��W;f�l���-�GkfF�Y�c2�[KYb�`&s�Nі6
@1b&��F2�Wi6x��Y��д���:YeSQɲņ5�@HU��U��B��Ť4Q�3D3���TrLV�h�`�v�pE��LY�g8pg�COQؚ6h���Q$��4Gnw`�5î�X����-#�������fX�͹�lE"��2�KҢqk0l�s��n�T��2ҹ0�%.�-�.��l-��D��)�R�Fi��MI�p�R�*��k�%�F6�k�6�P���m�\i]
�mZj����٩RicGG��"2:l�ػ��kP�H�D6%�]D�s��:�K�c��UεN!����"KoZf�#)1�H�cF�LZ�&	6a��4����ka�4s�kSE����.����YKbEZ�ڤu!$a��\�%��.J�s]fi� U�n��(��ȓJ�sZ�&�1Ls)Ķk
hK+7h+]A�Ե#�j.�!dB�eʔ��4���Ai���:^�T���-��@�GZL���l���X$�8Dm���4�69�)MK\'0;"�Cj4�CpZBilan��0���ƥ�D���$6�`,�6�b�@{k���h�m�
e��`T��n͚� J�Zr�B�C�1��ֳ^k	�m.��������q�X�.���X{e��MX�	�i5 ��F�*h��0�U6.�-�Eї.n+K5�5C���hˈ<�.�#��
�խ%R[D�,��k��k6��m��Џ3KBGgdB�7��o[B��YID���<9�+e���MT��W`�^�.m���8��;Ef�Վ���lT�+n�ɵNsP&�E�%f�f�U�*�fBZ-�L��QK��Zd����T��� ���:jJKh� 
i�����6��F�J<�a�}�>�61?;^-�ׁX0�u�X�bʛ,�ͮ��m6�J��+�(�׿�ĀA�qP�w`!3uk�{�r�1;q�^oP�x\m#�X.o a��'5�#i��'2ڰ��?/z3���{�|�����[1�O�{\��ڼ�S�ٺ;�_u6�w-�Rs�;���/,�����D~�?��˩��mV�ϻ�M�e��w蜴�屻 s9����'.�[�������V���ݛsg����-9m_Zm���Q�k{*:�N�{luF:xٷ;�>�����4M�'��&�=B��.����54y�X�����m�vsQ�!*Sk5rX�*��95����Uꇏo������a+Wwq���&�������������;�ԫ����R=���t����m�{|N�8<�x%�~3&�Ex��7�- *��ܵ�D�~^����ܽ������ywT�99]'2�ð1��yP9��}/�N^b޷�����7wtȓצ��B�O�}]���67`}���u�\)�#�1MN�{���*��xٶ��tkg��݀7vٵ��z1�N��.�ZQm�u+������J���կ�Uξ���ܜ��������]��GԩA�u�G'y9샗�ڷ[�����n��������??1����@_��(0
�&v�h��ٵkts"䅦���4]l-mS�7��^>�O�����vExu�r��d��L<��pu�f4����ほ�?�m���4�b��.�^;�{��Roc�]?b��VABN�K���q�-��[���vi����P�yVd�j�T�O"!#( c+R1V�����X�~��4��k?_W��C�p��\�wt&�u{�~���t�)�y�ɳ��_�����~�q���N�
Y�p/�\������N��]%��wK��|^Ef5b;�Z��ݑ�v�I��܀5��I�_#�j�y�WN(�v>��x�WG�W3$�j��5�0��mK]�\ZE�M�F�0utd�֍*ʚ0��q�\�n��w��=��0e��wOw7��Wt�)@ղ��wd**,M��+ �I�:���1�m�f��M�t���>ų�B����0���*��q�ݍݟ�F]�0洷^uӓ�Tt;������rӖ�w �A]���/h}k'T|7c����Hї�����|��^�1����V�1GB_�N�|��u�t�r��^7��J��-�:�ݹ;�y�zk�������r��Aީn�o�j�O���֛n��a���u�`v2q�O���mNR�@ղ��Hl��쥝�&T�& �:���i���l70�H���䖱��@���vk�1���[��7b�_n�u����;=� �ۅr�v���#v7b��{Gw�!Owع�;�}#E�<�n�wx>���ݽ�����n�m�v@������A_c�c%²�R3���;m��]�}%���݁��ԯ���L���@���)�n��۷T��wA��N�}T秪1�Ğ��喟�9��Z}�s�%���~��Nv���g7�6��f�v�w�}f������eG�㐏˹�Jz�>����P�����y���5R�7Ʒ-���TP�Y��SBE�m~�qZ���z��-��GH�{n�Ͽ}�<��]E�]U�����λ�V���fjfb�%K���T���k.F�U�h34i�#���Qv�f��/1X�ۦ��2��1��Qځ�*�A���M\��ɬq �\�����7\��bM��G-v	U3F�i,`U�.ar����҄@ԍ���H,�J6��1�a�͕!1{v�luX"kҔk��qf�%��D�VP��5pʦ���>�<k�˥m�W�V�X��4��K T� !�R4Ғ�E�P�����������7vB��z�����K2����e��Q���GVw�Zrھ�����]��n�lU�Q�xv���jvz���Vl�6�Y�rx��Ֆ����D=��ٽ�=O��NGrt���=�x�m�my����Xg�_���wdu�����_4�^��} �ʨj`<:���wg�O֜��O����9��~�G�����߀�{�?d~W�y��nNS|%]�$��0��B׵�-#2���]��R4m��mH[��3�<,�2Ӗr��_~�W�{�ܛ�����d8D��]�vGwN��ݐH{��~�s"(?g�v��.D�K ���/�jq���K�AаXSm�[Rz�B�S��h1�q1�ɹ��W����\�euB�qڦ����������u��Cx�5�w������S��R�Uحg�������OlYu�Z�:+�ՍOr1����r����7`;Xн���i���x�����ܦ���֧޶��ߟ4�	�8?_.����6��ھ���������긊��w�F0���S�G�$�o�М���S̛��,�&�Ox��DM\iP)���\3#��0uA���"Q����=ݱ�t����[��{O�Q�ϬI>�˅m�w�q��mݘ�
�c��uNWԣ���z���V���i����f������))u�T}�VZm?[o�������������*�m�w2Ќ��1B�Ե+N�b���91�xH����qB1{<�[���F��4?d�K#,��X/���ץ�߾����yZ~��Vec�7@һ��s3a��;�n���hc���[��T圹��^���+O֜��tL���c�#s�c��^��ղr�t�w��67vw{�a���ٻ�L�
�a�Í��d����QR��j]��#�"�q���{-#���o��|d��{�O{�+�ޞ��9�\�<�+��������i9@]\��݌ݑ��X�q��:����ׇf��gW���|�Hݏ�m9bv���;��n�����!��e��L�ګ�c�I��i���} f����v>�>Ζ�se%=ռ��[���?W8�����]�
�Uo}�x�-[]�Tk�uZ��lջ�O#^PY�o����eTk���Z�kPȡ��/n�=�e�jr%,r�f�N�X�Y
�H��]�����`n�v����P�蚭��>e������_݊WXx�E���|��AI��46��XU�:��+XiF�`�h�	���R㩉b��L��߼�;�ߌ������=���dV��M�[���F���;B��w��әi��Mz�grVÒ�����j�
Ovf���:>T��W�	�YI�}��~����_��#�����sñ/z�_���b�,�O֟��n�u�t��n������vݮ�Yu|�t�����m��*4&������i̶���n��~����4�OgYI����{�: Z�ỻs�"���?���[�);rT����{��K�U#Y��IP?M��P��Tl���X%ީh��5
��Ei
��g��y]D�0#�tR)�����A�[jʱ-nB���hX���%"k,v�3�̓A�e��%�#q����E\�WAM�K�IiK�F�PiF؞S��m�V=eĉLKn6���3l��H�Ylu�@`�]���se��%��л0���P�X�#��a5�(%�U
aά�h������;752:�طhr�pRd<��M�e�v�[�:��4>�����Ɣ�v�jⴥ9�eQ�p�]ۓ]���<W��U-�_�=yg}����݋���v����ݤ�:���6,%/����wgv ݇=��ٔ���蚽�c��guj��Wu|�t��Ϡ �w\����`v�}�g���n�DBe��Qޛ�᭭٬�{���`�ݲ���;�̧c0*�m���҅g;�OV��y'�����Aq1��,s��i�m����B#Ŭ�[���=��Gk��9Kx��� n�sv�p��0_î�,k�4�gcfmRS7:��E��F�s{[��q�A/�_g��N[S���w����6j�f���:�t/�S��Ol�ݿ���٫t.�:_3�d���t6�LMfۘy	˕����^�LU�2s�	���0�f�5��;��,8/��dJ�0���̋�1{]��:ug;���i��|�VKn~{�F�`m�U���w���wgv>�}���.|:��f�OW-ԩ#�{�9k{������n�݇MUfWE��}#���n�dw=���/z�*�e�����mY�E��o�����Ӗ�o�CNg�u�W����9ܮg�a'���{?f�JJy��Ԋ�U6%L�	(����-��3�+���Wp�Q��XVQ(�@{^�T��G�5��)(uy/��F�1��ӗ��KKj�X��=��8�@IO�BJe�̍��nd�c*�p5*�9���|r��5p����$�R�sS;d����*�js�Ԓ����71��W�{�Y��[.gV|6�;#����·dֻ;7dZ#kbZ��'IN䆉���.2��L�����+��I�e�f��Ϋ�يD!���l�
�
��C9�9eDj�8(�O[�^̲�Dd�����x�7�&��W�N��|�"n�zd�5r{�t�w����l���&{W�����8�x��8sܗh�bn���=��{ܺ�֯>G'�nJ�/�������_�Y��u��7Q��J[�f7}��{[��c�z�sq�.�%�G=��^=�dK����mر{9!
iKd-���P�H٤'���n��/>�y�I�V�7�\���:'Y����5JX�O7�����+��٧��V`�-�U���=��%*sty�V��eH����j�j�bwd'�c��s�1�(�C�7n�\"�cڶV}NG�z{��Z��ô���.J�����]�'�x��%gzc{_cѻ�!��?\�3&�\���-�5��x�&t� Yqv	��z��X��\�J�\��e�{X[�Ӳ�a>�
d2�Y��]�ÓHaS����C�\�R1%��ٔ�h,U
mZ.���7��֟	�v��]����(l�6�O�ef�/V��T*04Mμ�PM�Gvk����:uB!%�P����h���x46�򚗥3��/��Kaf-���r�݂OF�$̙���*r�p_5�'�V	=^��q"]I}Vw�Σ������k���s.��S���˖��{ɒ���y/f��h��`�d�|S#UӴaTr�G7Vp�^θ��+gÇkm�ˊ�"��������}��Y]�rst,�d"0�EF��]�����nnX�V��h����ZME&�RllV���Ѵk�lk��ѱwtF-�VH�خ�;�r�(��&�(��,lR[�,�E�hŢ���E���4�0 ��D3��%2���F����"MA`��(�dԖ��BE�شP��R�1�����$��`���30A&�L4���"2�Q���E�\�o�w���|T��u���($��\�/%lt�?����@J:���]��L^j����϶t=���'�9�k�Z�������"LC�<O|P�@xp��\�'a���\t}����Irn��n������a�&�Qss��#L�T����VbR�@�4yJo�""�Cx�K$'$�%7��K�S�V����fE	��"�h�S�	)IHJhu�1Q�2;:Gܘ����^n���ۋ{�>������wD���;Fzf�lwt���[� ���Ŏ��ؾ��H�M����Ώ��	)�(�%?1��Nt�����ھZڟ�IO�g4*��Ob�V��܈��kFb7�l��'����		�{r�p:;����CA�0�Ũl橉�bR�=$B���߲�g��Ģ����ϰ�C�?gC���% �䔤���鸅1.���|sw"sR�����BQ�O�,�]h������v���3�]���L�.JV����"˳^*W�m��Kx������o�?~]�����R=���u4af��mO4$�+���f���~I%a%"��\S��C����v􋇳�%K�S�V+MWm9f����/��`Wt���.��IJJ~K&����w��v�+5%����~	@	)IJQ59�-i�4nU�jS�>IO՝�T�N���ab�]��l�	9P�m�ꄔ���I6�و��p땇.C�{[���۵i�ﲞj�� I}ki]�>��v��W���̧h��Ԟ[#TP�a9ΟN@{A�����ᠯ>3Զ,JUf�>}=�[}���~��nq���s�"�e����! ^"�/l�Ж2��dGMp1�
�45%�ԪB�6����#@�,R��L(��nk��)�t����l�l�A�\ؚ���A�eG� �Pb4�ea����b,ڥ�B�Z�4ͪ��Cc�m�
�vaK�	��T�)v���m*S^k!s��!�F�ձ��
hX�jv1�0i�J`"M2�+m*�T���P���϶]��j��6- Ɔ,F,�ULm�5�k`C��m��,*Yv}���R�������^���jK���Xe�=�u�-�$�($`�D��A�����xw�aut�O.S
���;#��[��V��o�e�j@J>	)ID9����mK��N��UM]�OW}�ӑ�����������X�q0gaN���7�%�{i<�ʻ�I.F��}�Tc�g~����nBP�))�)��1�sz�;�r�Zה�-]�>�5�IO�].�^�-�~{�̰���Q���-�sv���6Q���F���޾y�|�{�ϺO�M��c�T���I��.�p�Ż�z�|g;$�%#��JZD�Q�ߨ���[���K��Tg�'����; ��銄~1�����Ooi��v"�
��4_��n�A���޾�x�"@vdF�	��}��ʹ��d��$�"�{��#T��99�;3h��N ���I+�% ��"b��.ct�3A�wS)oR�������	BJn&]�%�#i���f�IN\��8T�E�I��#^^aڨ��g/������Q�'))	G�$�|��9�˨�z3Om���ȫ�ԗ"�x>��W�IG]�w�f�1�b�MM�	T��mH-tۈYp��å�-��Q�+(��m��D�@ ���]�;\�$��w}S�K%���������3���%���I%`$�}���;ώ���� .S������B��R�[��#5JCy噼&��mHjR��9����g2��"t�W9eGS�D��-},����f�����+����v�> �P��E�7�Kz∝kq�҇ߢ����<��k�t��59r�5s��4i�}��5$�䔥nz1_v����N��9�V�wڬ�`�s�/��нa������9�r�RN��OيBp������%;X�Ku@����ܺ)<���u[W�])�R��J�����2��T�$��������*XQ%��5!nu5�*2[�
�]��t&�P>�s�J~	C{�jT�i��IsQo8}}R�g%��x�ۍސ��� �����a�]���،�mJ����W�Yk���brI�W��3�LNؕ���S�I+�%���t�+�T�*�,U�����J�.ԁ��% $�%"�xü����H�r��vqJ��5s��j��}���v���'&(N�EU��QM�r!*��pۏ�nv�L��z����'�q�r�m*?P�����R.�e��r���tD�m��H�%nTb�t�ϒ��JG�))����	P�Ɋur+�S��͚����\G؜������	P���,ƅ)�vs�TM�n�#�M��C(��W&��1SdIjO�A��� �H�$�$��(�֮<�V֧��Dl(wW�x�`�Cq�J~	)�(���Q����{�����B]}���Sun�v���I1@�*�ي�������I)�ݶ�8�p�T1칮�ۻ�m�ﻣ�N~IHJJ\�QP�1�l]\ml|��	)��(�V�+k�Un���꼑�Yj&�w2�i%�%	)%vX�Ƙ�"� ��ʎ�ی�Y�C��]��$�����]���3*�c�9jj������voo����lz|G�(��E��s�8��4�ϳY���C`����`���iU��i(|K!�gP�e��[rۅ�pt���6%�,�Y�`��]lM�%� .�M�C�O<��f�KpV�\��Mu�i�X�M��n�d]�ɠF]v�h;e�'#!h:i�cr���� SD!H�MB�B�]MDMifBP�c��-��� g�3w\�e5��X���Tn(���T���krf2��)�V�X����Mέ���Y�[|��ҟ�
8)��.�NÛ�%V�V]��Mye��m�7fQ�5y������wH	G�)���Т��7o��[V������NZ�߆�N�%a%8X��#mh�u����3�_�6�<U�}W��?%����<�:��5 $�XZ&^��0��yۺkso��v���f�	)�%?%5z�[Z��jX/rCp ILOflB��9�|�ڵ�w��+b����~�VJ~JJF���DwU<X&e��6����W��!(I-�VRʦD��8�dMQ�[�J�����J�D��q�7YZ[�he��~\j~IHJ>絼V;��̔��v��x���Ÿk�S��%)��{]$�[���4f�w�34� M,w�l��M��{��}�ć_6�B8h~7�i��'�6_r��p&7�y��Ta3��MR��]17٥UOvF�r�{�k�G؜����8"�*���Gֲ~�R�|���F��;��ck�i�����U�rI+II�:�Wkx���s�k���{ؑ�]{��x'N8|�'��M�E�he�ٹ̔�VJBI,ٕ;�ܧ��G����r)�ͮ�}���)	(��p�&��)n*�2�B�^��
�uP칱-�45�4�De�&��S*My��?5$���LDmv��#����=�}�F㋬`U����$�%?%JHߊ�ij���}W�Y:��t��y?%	%��//�V&Þ����\�������WZ�ߤ<��QxT�<MtNI��n��SF�B�kf鲱�1����J��c��j�����mg�dY�g6$�)֔�(��W������19	)J>IL�^-��׸��۵x�����J~yQ�Ӿ7�:�՛�����0É� f�	)J>IH	'#�]c���_f���yu�K8'J8y %$�3��#�>�BE4������"Mu&��:3ZC�Y�^]u���ʻ�UT"�.��Y���|��mju7�{=���ص�`dƊ��������徟�I+�% 9��uu����?}w^��sA�n��³g��CF\B�A�{e�������R��:�
�w�Wb
��*�ig�Gk� %$���J���
&磪N�dh�s� $�E�-r�:6��l�h���>�7r�̕j0ee娿���j�8֜�U/Cb4F��qH��î����Ό�32�A䉋�qȯ�ݑ_�rAv]I�8LB�EU7:�]��8�% $��Ȼob�Q��T0����b��n����gි��J9`�u��f#�R A��Ma,�c�CT�&Am��Y�v)cڏfJ삲���A����R>J���]^N���	��|2�D�e���8��S�Q�J{+����&r����r�s�\�퍪kv]�uw�.��$��0�{����ꐒJ�I\f�q��p:���1W�ۭ|)l��������a�Un�G\�'�-s�5!(:�P}U{;{K8'[�7�q�2��{�U*�T�������S���F^e�3�"���t�W,�v���>��Z�X�����7�ME�1t���8��-h���q�Po`��W�d�m2f�NelޥLj�4H͸�4%��$V�@�*��8���&�P�r�`���0Y��A����lD=ѩ���q�Xʆ��'5!�(�²�ܐȊ2�*��l�j*ao�cv��]T�޺�gگ����?���Zs�ܹ��e���K"��l;l^�+u<�ˎ��C$�(`�L��47�����Q=�;i�L�k]���v�N�d��a�~�(�"���rv&���b�0ܹ�z/��M]:�*W9a�l�E�{}6g#�oͫ�
i(�{7<o�w'�S�"�A�O���e�ʱ'���ث3�P�Y�L��q1���',0���$�OmK�n�c���h{�]��^95��3SpT��wS�(��Z���j�]��oJ)\X�<�Ĺh%�����3�� ����<�{;����G���G�x�s{Y�8^m��os�bBs� ��Y���uЎT��i}�wB��bcQs�璾���mբeN�?h�%�bʙ��lf^U8O$��ڧs����{MS��!�\8;O'<G�+^�+���{u{`�2J��g��A����v/�o�=}��\Ҩ� �h�r�q��](�f�=[��^���bҟ�
���hq�y����y1<�	yogf��n�Bί@��x�:)9_��Xȼe�A�Xʉr֭�wm:�3n�hԔ�ʼ;uX�{��ۙ8�!�NT�8�	�w��Gz�\c��hߍ��z�)c���;��1T\�W
B��)���� (ł��%�ԅ�H�Ʉ����X�(�E���l��(6,�6ɉ
�%�H��X�Ԑh��(�D�%�bfC!��2,%�,D`Hъ �E�JD�f�d�6C@Q��%��dd�6�JD���e6Bj`&RDT�I��I��D@��cL4K4B@`�ę�2�đB4�@)")B��LQ��"��&d)1
&H%2�Db@�D$F13$FIF*J,��2fH$�,��,�d�&(C
8�y�>������Y�K��I�B�խ��͚R\�Yf�c�)-����1����c�4[��L2���5JZ�4tF��K/,l�o�Z��ԓe-����6��-�C�2��n�j���Hut+vفpC&	n,�z����d[�K�6�pî,�X$14�� �y�⃊��e4&&3���U�iPٳJ��]j�`�0���0���4h�gGUض��[���{CRk,��5�N��!�32��p��2�cX�U���p�ef�I)Pa5�u+��	rDf�Fڎ�lX��%,�blJ���^�����lާ�����2��ܔ��r�*m�ţ �bF��
Čԅ-�3p.�*�iq��4�����"��"�֗4�(�1�;Bٮ¥��̗+^-��^̡�,)ԡ�ב�����L�#v��5����Ժ(WY��j�\G ����p5ق��MJ�7b�qv��t�i�r"�I��e�[�mal�;�hS��I��
�0��2�jBm�˔�L �s-�z�6Q���A+RY���be�&[V4��F��R��c(����%���Jb�	6�e��ذ��e���l�Q���;\�.�J�˳��eu��b�K�au�q6�0P��wjL\&y��Ñ�v��k���Z�bS.щ�����F�3���!hA�L�:ݘf4�¶0VV���`69Z+���,�o[Act�ɭ�{g@#1a�e˝lԋW��	�2�X1-�jcįb��X�g\�xH��(��l���A�ζ4HlA�WWI�!f!�&��,f�(ā��Cl�E0،�m7(�[\]n٘�%��X�ͫq�I5�6 mM�&u�c))�8	���`�בz�1�%s��ˌ`�-��j]��@*��iCM��ڱ�J1@�s�l9eG����<S��0	Z�A��x�e���k]3nĪ� (b�˫K�Sd�m&����W�Q�3lƪch�rir,���������$�F�陫%f��3�c�+
���GbV:bʋKXL�z���8�s1.کT�cr���D&JB�1��:����]*L��V]v�͌*�#p�KuVnlݢQ�k�s���ێ+P9،�3��6���B���:����`��b�#���n�*]�ФqڕHB���m�ib��:��U���`��l����n,�ْ�$p��~z��ן�rJ�Rr�ЪӮ���r�k�j%�RN��fO����I$��Y\{���5�r�9�>��}˸E^��R�	���bV�Uq/����\K:��ٽ!%)@	&z���e-y�8�n3"v�l9l������$��������15���R*/�d�Ng���/_	J~��^�]�)4�΀1���|�|����+"ڧsC(l�����y˸��ܫ\���~	BJ~IM��<es�����T��АL�h�%aְ̠�Rl�\]�Q&5oU#�]�������^>|�Nw��$�2��ϯ$L&��Lb��U��s �s�}<����R���q��7��o��#gߑ����i�(��h��n==E��|i�����&Ipz�杧oKQۧN��X�Ԯ0�=}L��B"�r�������*Ӊ�9|T7����]!,��Nz��v�z+q�r3\���JBI)+{Qu�mv�^��R�	��}����J�IHJ>q796z�[�	�������ǝvH�\��Lb���w��+�TJ�͟�I_�)(I��+��G�΍��뉎l�oW�����%%R�5.�$A�U���u�i���6Kj�u�����kJc<��M���=�MHIH	G���.����8'{ �T��F�6�p���O�)J IKSP�ln�Em�̱{'ҧ/��>8bjf[»��>Ƨ�Kr�V�֭���J~�RQ�J@Iq�j���VES1F5��,ѱ���)@��|���ՄrY}�O�4�,�n:肗�r�L��6��P��˵Z�n���Z��9���S�l�ޮK�%��Q�JRY��gWv��\���%i���k"sVc	��}���6ؙ�nn�O�4������A1o#H㻎6���!f�᱋�}����)�K�ZNn����L�&�SRƄ�:��-�6ꗗk�b�4z�A�e�6�laThͯ�ꟃI$��t.{ƣn�ޮ�{��]�_�%!%?%����]Up����������k"sVg"�c��VJoo*�X{��V�꟒S�Q�ILl���E*��]�%�#�L�lf�}bI,JJEl�L��^���J���nBJ~��3�s��v�pm����4e�+��L\�RQ�m�r�Ƙ���P�.Ï��:[�~9#^>,霵.��yZ�Zv��a���❬�BC�_��׬������d�˻� ��J=�"���#�|���,��Y��[������RON�{��ɽ�����$�M�@���[m�4Z@v Y41�k�34e( ѓ� ��u}�kJ�IN��p���iqpؽ�=&�b�:>�r��J>IHIH2�T�s�.s�_��wzEFq��o����7��ur�� �u�5g�EK�ۑ���� $�%!'Uwʳ�pS�����,٭x�S{��(%))	R�:##)����?j��Jw�{L��d���ܱk���	n�Nżג�9r\>]%))	@IT,����9S?Tk;��D��%��}.���� $�w�f���hް�ELTF/얹�K"�ī[�r��2���Rp�]����٪X�d�n^�1I���b�ǩ�/�^�=V	t�k1Zs,���ftkִ�R+&p�kM�i�-�2KqB=�%د [��l�E�M�KDk�Vf�m�C��nb7kl	�4,Q�c����ku�sX�Dif����24�Zih�,*���U�Qnc�X邚kI1�+�Q5�M!,gĤH<���Y���:�͍�Pc%�,3,&[�h݁���2f����f�uq�������l�F:h�M�3j������w�I�R_p^Y�?q��;�gv�����Kvk<n��V>�WUH�ξ�F��uH%)BHn^aT�K����7T�r��o��;���b�ݩ$��ٳ�g4��T[��� %	)	$Ɇ�`�FZ��q���Ν���m�O\����R���of�*4s�1J] %_[����z�n�i��˵%�c:v�Mo\��HJ�)�%!)Q��c��Ο�u�������<�1i��K>K"����}���o�I����	�ttS���0b�f+
�C�!�˙i���l�H���$�߭Y����XUnc��tgD�L6��Z��.{�Te�R�RR7�}����mȠ[�;�V���
^�Nm��,Un��[����c��oM���x�)X*Pec�sX�$9O�X]�z-����XE���UmNF�w�1p�.PݸF��/����|#��������N�ۦ�U�_?)��-ȐCn,������G�_��A�����n'�ŷ6!�x��uϤ^Y��.v5Kn����z�
n�m���r$ۡC�vn��7+Ly�?X�}ꯋn�^w�S��~���<��x��@��"'T�yqr(�=g�<}� ����!�B�n�n�ۗK���"A6��!�!�Eﻧ�\�v��K�:��	^S�|܉ ��}�|ۑ+��ތ�F̙�ER���-nF�n��6k���e�W�b;#Y�6���`T���or<%g����
�� 6����=���cay�~ߨ_�tW�z����  A֨P��k�ro+���"�ɹ�n������_W��{�E���^����FǾ?5�D��P-Ǿ�mD؃���v�{�I�B�-���_|��5��}Q��7o��Hj���a�a,���}ʝB!}���|����ݬm��d�d�:3W���s�<�:�Q�W�MGj;��9ܷ7�ᮤx�z~���WŷB�q$t�u�FU�ꘫk�}�_}��G�$Am��Q��׵+���6���@��[G��������$6�W͹��-ȟ�i�'u^q��c����=��:���еg���r<A/T�@y�n$Am�{e}�6y����1���b��mp&hVmn�tƹ��.�e��(��j��6�ث��������BO�?6�H?7"k:�=�>�{��|6_�eO�b����{�`��m�����WŷB�q �[s_�}+���:p3�=�3�wA|�{��/�ȍiF�o��A]~ ��P��{nh�f+/E��"H�گ�sD܉!�U�mо윥����̋�C�]��pߍǏݪh|�
��A ���6�P=�{[�q�|b ��W��?hnD���=�Ǚ*kw�e����A�OdzuG�n:���s�0�1�E�fD0l��b�Q�x^-ر��7��4u�(	�TgM=HE���������x1�T+DE\X���B�?jt(�H%�?PmЯ�qon��:�c��qw�Í{kjW7���(��	���n�|[s@���[�MT]p�?�lBX$�T�������P1[h8�����	q�Sh̏�w�#=���	��4'�_�n��{-��>Ig'q��#S��L?e�{ݓ����|WD�Am�۪��Dw�Ķ/*-�˾w��ހ��������Ju���G��9�rmϺ��6?�\�_D�)9��!�B�-�� ��U�C�~�5Q��R��^��x~/�$��n�|[s@��r$ۑ"A8:VK�Q9,WH�F�P��n�}�=���G�Vy8k���N���X41C�ɵ�(�A ��u@�[�$6�Qm���en��xYy����8�k�{��J{y�9���9��r$��W����)��ͣ���˛�e��%�s�n(���\+�Lj���;ƺ�ݑ�g�J�ᣲ�����wuJe~�?r�E<���g��)F�u!��m��,X��v��ک�4��霤�7��c1�U�1�5Z��[�ݑ�[T�l�k��|3�<�5��7�8"�)�u�!�2�Y(H$��ב�r!�������J;����LU[(r�c6�J�Zg�8!���^jZ�`*� ���쐷[4�om��$�MJQ�m�A�2ڳ8�)�F�CFݣ�2�p����λ�'ϓ��~�/-�Ie[�g��YL���ι��l�j�-+�bk���}���h��(�H ��x��A���R��+�⑷�Dl��@@�-���:A��7#nh�fhN�`���W�S�Z3�����%�NZ����/:���N͉��J��@�oH�y��ͺ[sD7b�n&�r�ǣN�y��^���@�}�h[�x|۟��xQyꅱ��N��P�����4�Ŵ�z�jW�9^
G�~�$!�_z�ֺ�ѾuzhS� ��@�����w����zf��7*��ѽ������x�xAz��o:[� ��m�;��]T������d��X�~�1�)�[��	@\X.6��,�j����@n���f @ �1��<�H��
-��AnD՟{�/�7�fRyx�g���3q�z�ǋ�9�A�{�|[u�q�ۚ��9���u�l��F�!��1B��ɭ8�z���>��gx�o�V��hl6ꠦ��9
�t�N9Nsة��Jb6�6�˸V�x{� j���ɧ0{ۛP����8�����[s�Z ��!yR$�%"����!�����ͺ��={'�l����Gor�u�կ�|A-��ܝ
-Đ~-��t({��毯��Q�:�
��r+=�
�U���<�\g�o�?*��麙���Gr�_��n0Am��u�p�=��{�Cv{V��n�5���w'"=�ݥv�xR=�~�?G7B�n~���ſ}q�����k>�>�k(����^M ;Z�гQ�+,]�Db�͚�[������C�߹���$۟��B�v��S��6���Q�:��(e��*�Y>#�R(މnh۪���nwϷ���{v~������yg����^��W��Mr$��J�:���w�(Q� ?9�AmТ�I��ޝ�(�<|N���ߍ���̈ɑl15x.]'a���)yy�u�4&�81E<��N��R���Ehl01��W�������{��Ç�E�QP��ϥ�l�t�˹m��<�A�g����������]�l�rOwv�2�����s�<xo��䆢wN^����������C�-Ɋ��({_ý�Gi��4Yp���D��,S	���1��E	�Bj��k��[�Z���t��Y��e�]׭c�S��&��Ö;�7��ې�E����ǚ}��3<
v��{�̌�y�f'L{Sg:���~N{��}پ��׻��Ԝ��of���o��kp<˼�����j#N]�u�	U��UnƱ�A:��f'XwO��Bff�Y�4ˬ�Y��sk�U�A���,}�n�����|ʚ��9G�7�v���{�}�8+��|�g,[��9,?{������>��Ü:w�秧}��S��朳P�تuj�5���wn��:��L�'�`�k�\�����b���s{�(�Lh���d��}1w*��çV���5Ox����wܥP?Y�{�	.�I��p]ev�3�w�g�
�N34�l�����}����Φ����[��b-��*g�L����[�j���E^=��m1pD�ޤYۻ��4v{�$X�U_e�ۜ�7BНФ3kaꧮ�r+f�n�����=;���Ժw���m�ҍ;�ӻ�A��p��1�8������g���'���0�a��Ob��
��{/Y�����<�F�rU�iiE�މv�F?�P1�d�(�a1&F	�R�MQI����1�h#�$0�&HЀ$X������$!��#&a ́I�!�&��2D"�I�&E�B54� �"1��(T�FB�$(�Y�0�H&"�Bed0e ��M�I�$(�L��
3��$Ă�`$�,I�JI� Ɗ*
JM�Ĳ�cRde�L��d��D�2�L	��a4R�A��#&1�b�DPBP�4$ʘIdD��Q�dX�̌�f���I�A�

����" ��^�ϴWy������^�A~�$�B�nk�ȐCnA�tw}��=�v۟��F���6�V��tw8��G�[O���8�h��R&-/nh�Z�A:�hۯ��	 ��Wŷ9�T,�$�;dNnzS���3�n���#��=?PnD�u_6�R���������a�:9�jҭA��kedk
�Wd�n-M.�;J��T�o�����@��������-��[sA���q�ݥk%xl/P�0/�P�Ni(��ۻB�-���m�|ۚ{�>��E����#���?H��.=�2'ǥf���ǈ'sf�#_H��o��fg��DE1��4�� ��$��MТۚ�W�\oD�9d��}y��f7�ӧ��@�g����H6�!�B�-đU�>�Ә@�k�ӄ_�E� 6����p}�͕>k%xl/P%��=�^C<*g�Ʋ�&����T����Ȁڍ����7�S�e������Ƶ#��$��4��pz���}=̤�^�<c#�y�V)g��9�zD�t([s@[� �W�Ώ�6,��|�:l���}�[����x�z�?^�E���n^���>xkߨ�K�⤺0�:k�D�8�\f�G[]L�.&M���f�M�m��;��6���嘄���'��|Aȑ^�:}y3ޓ����.�P�7z��{����/�H#yЯ�n���-��<�|:M���_n��/M<��4��ۛ*|�J��^�/�$Gϝ|۴����|_޲�߳SB>��Bw�\F�W��۠cC���m�ms^*��fb�[������4��q?�s@��}B,H�u�Wsm�@���}Ӡ��Mr^�u�=�9>�R߇:��	�zh�ױ׹���̯|G�O��}B�q?Am�mР[�L��mU�f�a�鯯�/>���ʟ=�~W��@ �΅����mz��zbO��D.�;&*B��.�ȼ��3�U�9�D��X1)I�ۻ�����40{�����+/߰��� [MY=����N��YT��Ԑ�۔�U�v�QYJ��Ӝ�s�#�r�*[k	���5�$I`�WQ�4t23;JX"��qHсX�.��p[�XZ̏e���f���I��IY��5��q��a��`])�km(j5�PHLK{v1�eWm�v�0�@݀	�]��K(�M��V:�*�Ž��c)4j�Xl٥*�[�Rn��ya炝��4�ݥ��ITm���E�JQ�@�[5#�����]����N{�@��"A���n�h�>:��_,��x�x�{��^aw�p���B��A-��mР@-��.f�x%�vto��{����"���.��NH�E������Dy��m���/����'�����
-��~mʫ���,�쫝�꧵��{r����A�
-��-���������g�����;�'���|ۑ]�����ck�X���� �w\�s�2w�
u�pE�H?7�D6�
��Bn�m�@��A8B~��K��]���E���7ޚ����� ��
���m����<xDi��&�L������c�&�팶j�8�
Pз6U�L�|z �y���(� ��p�ϟM{keM�Ǆj�Y������[�_�h~Ȓu@�ۚ��z�򪞞�|2�XN��;*�8�#0e�B�*i��5EA��o���.A��5󭃽�����@ǈ���~D��\u?�5� �5��q��9uW���\���C���yZt����������+��]((@0 M̮р�)�7��� ��|۟�7!T��#�{�}eR�0n�y�W��M���yȐCn��t(��9����U����%��+�ޏ���xg�Ϯ��������5z�+�'�6L����P����G8Cn��nhCr$۽șR+�+����<�(<L��|�����Oի�+��H �ۙ�?z��?��'������e�X��a��^B�ZJ��qu���cV�@3�_�|�<��>�=�s��"kyS���&�Ԕ����C�(�23ݔ�M�܉r��m����[sD[�~G�y|�Q ���\3��]^�ٹ�<s��@�W�	�
�.q'ӑ=�B��cqH��v�=�4!�mЯ�n�ݹLC��`�Y!/n�m��v�ɟX�ص���"Sc�����K|��N��7��.e�F�Tib��yC��V+$�J�{�S��Ʒ��j�
-Ă	m�۪����Q�O��s@ �T(�鯈!���렿7Ԕ���{���鯈>�	�.�E�O��W���[sDۡE��J<��~��љ�ۮ�l�߫^;��R=�^�$΅��_7#*��l}����1(��rd���ف���3���Z��e�LQ��f&W�\�b��������~��~��<_�r+�W��\N�o�S���.��9���_�A��M��-��v/��~[3�yMG�"k�b|����3��R߇uxP?g���D���G�l?�}�(Q?@>�����
-���g�sؽ�JCX��-��{m��^�A�@��=΅�����}C.�a�N1��J�~��"A�@W͹Ы��P1{��j]q�� �v�h���O�k&wr7p��U�L��GQJf'n���y�}&%��w��}]����Y��2 ]gU�|,�f9����A���2��ޢT��g׎,���Ӯ��n$��M�ͽ�An�ۑ@��>���ƈ��!Z؟;}�3��R��9��	�zh�p$۪������龟��y����v��Z�1�n�%��]�@sqvV��IfE�#s*o�������}��H?r�
��	m���~�����y[{~[�k�I�G5"��� � 6�`-��)K�b��h�+�����Wݨ��	`�m�zԺ�����@F�P�[����D������<�t����I���?kr'���|g��r�}��Q5:�����}@�����I����_7G��.ќ����<f�> ��B��͹��3���훺޶��Mo��������3&$dü���٠A}"Hm���nh��I�y���w_���(�\'�6Lf�u�%ώǾ?e�k�K�(�~ �ۘ��7=���+�!4.�����UQ#��o��_/I����Z{$�$H�B�����E� ��>�����FlSe�p^�K}�����h7�=�i���L.�I`iY���0cVb&�ch6h@,�)�f�j�ke	�CK��v�G(���ST)�.�)�YyI�om�G�@�*�q���uVcM	�#FX��Z�m�� �ZTscl�����(E%p�.���o���cդжf��5ؔ�Jg^���\�L��t\�e!l�
GXv�m3\��`Yv��)����g�0�K����~ʖ0�F�m&�cE�W��xvX�fŸ-�m��*�-� U������ie��Fu{�
��� �܉�l)�}��j������|(G��t�+���� �>����Qn$	m��w����Y'+gi����_�k�^�쮏F���5��w�<��A�t(���G�O�.��a}T>nh~nD�u_�EQ��������c4Lf���%ώǈ ��hB^�@�%�4m��5
.|\�e�B��{��|}�M A�7"k�=->�	Iz����dx�4G���U���^��_9u
��A ��6����͡�w�UC#�>�N{Fg�+��;u����w����I��B��4?7"��~�_=��S���ͳXԇ�!j�l-1��*�7Mt� ��p��Tn?e~=�~{���lm�¾!�C�u��Q��{)�(������3ж.h�;�B�t} ��!�B�-�/��A��4��a�U8�{��G;��s�9�h���yN���:�X�~�X�5�������ڻ�f��ʍ��9��������|R]��p�^�^����D���x�ч�8O|v�Y�D�~����t(�~m��f{н���`jcwm���]��H!�Тۚ�H!�B���ު���>���$y���܎K������ֳ�NyDx�Y�A����.��ޝ3Á� ��M۪��Cn�ۗUNk��J�5>�3Ӝ���n���u຤x�zk�A�O���
��#}7h7�������O'�}۰�2���V�.�ؑ��,Y��+[����e�h-3`�V���w��߾��|����I��5�.͎����ߓ�^y��H���>F~�.>�/B<����RSDfs��c5t�[S�rt(rMyvDVD���'s��	���/P��T�#^]Cr���Dcs�p0Cn�|[s�7"����'*��g {|Cv����1�����vq�wv�O)����3}}�z�6~Z2�~�����[Mce.'V��V�N|\���@��D�ۯ��ۡE��To���v��m�
����������z��{�|.���}A`�Y�#���
N~��� ӑ@��n�ۃ��J��q{&=��>T+��r��t'w��;���禁zE�}%�/���s�'�$�Y�T Wǌ�-�(�b��`#�^B�`*���YI�0��k��0�'���A���_�� �#��g�;�*��V���
u?`��s�.�$sꯋn��H �[s�8��W�@��ϽH-9�ב����V���W��}~ ��
�1iϵ��.��_*���MnD�Cn�|ۑ����{��٪�������N��c�A��������H%�?6����sH٧��0}��+�RsD7~�����I��[�>�������}bL��X��$>�?�ݻ<<���~��{+��#�n�/G�~0�7� ����Uyv�㍉-H�IJh�&'+��f����
��ɹ��n��Мzo�Kc���=�8���g9Z{k�^xW��A�P�[sD��
����T��֊�eأ���˥�v9E�%�aRha�Aw�a0�z�;�4A}"A���t+༱�u�]	�^�o/�c����|s��ݲ���މ��[s@��
���y����l��({4��O{ή���W��^���{���D܉!��=��r�mg���*�B�YA=�h��n��H �ۙ�u˸E�|9]�){y���Z�+3��= O��+�ۚ �"A����.E����������@��"@!?U|[t)r���t';�5���|A;��!���QN�N��>�ϧ�ފ�I�B�n]c�譨�sfX��K���G�Ty$��|_��~>]4?7 6�!�A��۽,FL���d�ɣ�ţl��6�����GJ��Ya��$;�|N�yQա���݊^ͧ�7�{��OgM�~=�ob!^8�]�捔�UC�;�#&���]��"Q�&��츖D	̕��
��A�yJ�r,��{6 Y�3}Wa.�f�s�R\-5���Sr
���Wx{�3�V��h���F��=�S�b.�Y0��zS��fż�p��T���m���N8J��[pC�Gr{����=,�#}'�ҭ;�^�ξk!,��6p!%�s>��.����&'rޣ����r�V�����f���R0�{����o��P�t�d��W@������*A�����C�	�㤑
W����+���.h�݆̦lnk�<|9���w}�t^_@4U�"T�t^M��_lf�pM��F���;�\��<���猑�V-3q�D��J䐞Rzl�s�B6���%�%1��=n�#!��BdCF�\a�i�͌_f��C���c���iPi�봠%��[�+�$�]�jb�Ep�Ҵ�P7+����	�!���2�ed�:�T�y�Ɲ)"����z=��{�L�L!	��y��GO{Y=��V�:�;.R�WӶ
�(��־G�����{xH��}�ۋnƱ��=�NfktӋ݃V���w��}��&��w��{N�����<���������{ǷCx/��Z�m�Y��Ck,��7��bI��=3y蘿z�*Mo_��Z���|  `���hR3,�	`�2"�2eTRB&��0�Z"K F��cA���AA��(J$��b1b��X4�HF�D�`(�cd�T�E�R+Re)��1���1b"H�ȅ&�"6L`"4�4i�&�4AF�S6	��"����FR��Qf�A���`�&4%�1�D!�@Q�ĈlQd�	��Q3Pb�hKL#Q01��LKEIm0�bP���4�#j&K(��&���&� ��AEF�`�Ed����Q!J)��61b�(�� �Q`ب�%,V 
#�`����x��m�ձ�,����*X����4 �%lՕЁ �`i�a�bP2L6�[Qe5)�$n)
��R*�(��Z����K �����˳�2&&R]6bg�[���������mQ�&&m-��Y��$ٶ�6V�.b�K��ec��CT(7k�fe5�,�	kjK*�W����	cE�ZZ2уz�k5W@�k��l�f3F0�lWku��W�QWsHf\ie"Wl&�mL��Y�UV,,v	�-�Y�il�Ҁa@�_^��M�tKJVK�3�u
��z�\%�3B���T��@85e� k��U�Ķ$���#�W��c���i$v6B�Mi��ћ0��1�`ĤjV�pm6����a2[*��,1�sH��4Xr]��5�ůPZ%l��CK[MB�(R�eX�P�#�[�B)�X���lE�:ZQ��55X\!�ra�17fЂC^q�ڴ1��9�&U�������h�nlˍ�[�����h0k�֭��l�Ԛ+���4�!����`�LkA�m
��hT��@���2�g]63�T'alX�o`��Cm;v�1�+�kJ�(ٵ�\mH�6U	qPn����̸Z�74�α�d�T�fK��Aa+�K�����Üu"�⬫�Z�nm	���^�44133+�	V���h��	�m�ͩN�1�n�L��US]6V�&�h�F��Gɂ��R�s���6q��Vh&hm���R\�380F�h���f��$��T��:��l���J�^^b�X�K!m�t��Ǯ�2;.��3��|�����(���2�.fie%ˀF7��^�V1�3iU#o0Ѳ������l�Z;Pp�V��%#04�hV�D!6�6n�`�Ӣ�Ő��:�[(�F��hK��,`�\^��Ʌ�l{b����j$�o+naGj�m�56�:1e4[Ec�1u�%�Ԧ��Q!��E;3\��R�m�n��K��!�X���Uι�32���A�n�bm`��ۀ#i���n\��%�khTV���)�K�f0ӰgFe���	���B���I����[�:��Յqx�,��v�f�v��y&یH���Mv �nl��͡����Vj�u��vi�̦!�,\�z��YU,�H�.�r�3
/Y��nv��"ȸ5��*�Ѝ�ה��i�;2��a-�L�� �Cb�"�c�<�?O���$ɣx�0Q�:�B�M��i���Y��Ce4ll�n����_����-ĐKnk��������S���{���F��P7�%B�}4-Ȓu_6�!�;��su2���� �N�����(�����<��|v<?�Oկ�(�Y�r>�y��W6E�P�A��O�6�P-���r37�a���IS��.�F�P���vz�>N~�܉!�_WŷB�q?Gn���F�G�$�[sC��{�Ğޯ��}�$�7a���T�j~�� ���۝܉6��g>�S>���&v��c��fG��5��lG�s�� �~�E��Knz��:�O�l��]��~�G[sE܍����S+ƺ�� q�lR���[v]�7���~ٸ����1��<��ȟ�c�+z���g���|o�\	�y�w��p#���M����nh�N��b�1�d[�b�3;���9:=�LLι�40u�w���޺0����>E	��h����N�PC�Ӿ}vo���ƻp�Ļ�����I���}��Ѿ�x{G�7���7'�� �?P�۝b��ު6��v�j���z���9��$6����"}�>"A�Q�[~���	����jw�؏|~�٢�_7%�4CnG!w+���,�
 ��O˽:Cp'�dyk���)o������sDe��9����K��������~m�Cn�Ⓟ�c����c�v�=����x{G�7���7<(�?G��Wŷ4A��Y�(�z��D�:��-��\E6��[*J�rCp���@�ԁ1t�t	2I�5��P?��_�H!�?6�<�椋���z��lG����sf"-oc��Dޯ�����-��=����y9��Zƀs�h��=`��:���^x^�o�|��9��S�Y�M��zdP<�H ��@�ۡE��Kns���;��Yپ����KIH*��7K�۩�w�~kg�~���+q=��<��'喔vxt�y�p��L��I��^���5����p5����Œ=�����>�P�[s_Cr$��
�IS�Z�y=7�7 ky�mР���t���z�g�#��w:h�rG�Tro�0w�$�t�ۑ��H-�no���j#k`�zD��]��}6"���xx.�@����܉!�?Pm������h=�'��|-~XR1�]*A�4`�@ըW;`�����c�5���m�؇���!?�����WŸ�-������g��&��K�Pj��^���Qk��!��	m�|Fza^�<����PDnt�Mu
�떽 ���O3�c��:h��E�����Ņ��s_��P'��ɺ[sD܎���ULܾꋜ�`�Z�=V"�M����|(�S� ��6���q�K�B�/Q�5�gW�џ�s^�����hO�^��� m�ޭ��϶���ÍoJ���;��^{Hۊ�j[��ŏI^��6p�3*N��{܇v��ٰ��{WE���Vd�ݾ�[���R<[s@�܉��ɚ�-|���|��9��I���<O3���6�hF�P�S�������7��y�@�Y�'%�.��۹6�S7+���m�km�lcGYZ�m�~�>y��,�)�|۝�r:���#ޫ>�y��]��4�^�M��O�&��mР[�?6��r�R�����I'4;��v�{|3żO5x$�x�H{�Qm����1�F�_w�~����ېm�۞�4�T�vrvs�h�1��ƞ_�ǀ ��?V�P��q?~�4Cn����>&v��
!��G�� ��H�sX=�>���3�=_y)�=C��񮍘�y"<�??9��d[s@�܊����\���8��驥��ۑ���M<�ẽ@���${�P�4Cp.';�Ff��=�Y>�Mf9{&��[4��;9��i�q�������Qp���^�/��@f���1�qM��ў�e�#��MUe�A�(���Z���9�*�=nfպTz��4Zk.(YR��g� �5CW��e[����VnD�`B�%n��SY�T��l� (��l��V��]��3`Vi	B�x��h�;j�R��&����b;�Q���贪�%L]�f��F��\�*:T�1�f��Sa(�(GM�d�a�6��vx �[tTff��߹��o�B�.0���]ve�swm*D�-�c�i2�AM�h�\Z[/����a���!�����mЬ�̦�Y��4�n<F+�rպ���f;���#����|A ���-��C��ڡ�Yu��Y����8͚ �"}`ް�z�O��s��.�W�Jh��"Hm��:�-o�;B�Ȓ;�~��
��H-�uW�>z}-,��o�;R��^��s�$G���nw��ȟ�m���]�ʎB�F:�O۪D�5�~�ӡ_g<�a�Ո��[��q��4���"�}/K��2�H �[s@�܊�A��B�m�{��x_{pg�$/K��4z�S�g�v�P?�M|A�$��W�6�Sc���hD��rCl(^FD��-"��X�,I�e��^-�ɸ�4&+�_c� ����zE�A�[s_�{�_�v�e�K�z�1�PhVL=����G_�O���(��A���	m�"��w�60Wz���P�F��;�L��F�Kޢ���#��\�>����2��S���ոys�)�1�F�]7=�Wn�VujH��Ν͝�[�<�c���W�w��	����h��x��=Q *s��~t(���q{����m����D{@�}�AmР[sD�_�V����e�!4]O��6|9�
��h��"Hm�|~m������:줕��ޡEtH������z�;³�-���m��������wb�����ͺ�`[4A��H6�����܉6�lLcs�x`y���~[/���]k1Z��D{�ƟMZ�
 �Im�e�m�O�}sHE�(X˴,rl�.&��e81I�\��Rl��H�Z]�~�������x�y��7"G���O��7<χ5�3;f�_��_��y@�9���܊��A-��6WN[*wޕ� _�H%�M{������>��_��?v@������{�.�/1	H�G����t��H!�B� 6�s������3�썻���4h��Ü�D�"�#��P��#Ç��:��FS��o��η�O�-�#7�ޛ	�HUR�2�OV��d���ju�*t+Y��Qi�h���P��Iۚ!�T�G��vG�{� _��B�<�~��u�;á�����g�=�~>Jh2�Q���wu
���q$ۚ!�?79�+���H>�MZ�o��|}�k�ƿo�>�#��(��!����z����~�?��6��#,Q���P�Ꙥ��Q�K�c8C&WM���&�о0=��������B�_c�"a������D}��5��;u����@��A��m�|� �w�y��O��1[��/H�=b�{�3u>���|9�䦁zD�Cl��Qꂣ*��=�B��D�A<�5��B�n>�nqLk����z�z��1�Gu���)���A�H��nh��O�6ꃊ��o.X ��D�F�P��mЯ�_=�&c��oqxz"=������}^:�Ng���ݺ��4�35a�Ҝ�U��VU�*[oz���{�O�b�p�vx92��=�FD����Jo����Nh��
��	6�P���GE񭉼�,e����su�3���9�|�h���m�|Cn����M��wc�S;4"H��&e.��R�i���M�F�F(CK�f�q����,ױ���7�"�q �[s�w�;��H��;��NC��os�5P��
�����u@�[s_o�Ϲx�c�k�_w�Aƽ��L/!w���:"<%女w�WŸ�y��O�6�5�h�jE� HmР[s_Cr=������酥�ֈ��ς�����n~�ۡE����y�G�}�b��Y>~�@��H ����W�=�YQ����e?P'�A&���4���P�5���m�|ۚ �"Hm�hr`��r.���-���YB�=�k����ݵ���|~{�A�B�q Knl|>�����ث�23�{��Ҋ<:��|��.��g�����񎓏���'���G6�Z�&�8D��7si��Ds1}�t\��X��Y��.�at�]-eD�s�E���%�ئ4�t!��8֪:�K)KDu�Z��3l�0R�qF䉱NLD�V��lf��,\RA4�䌹t���:���s4eظ��5.\ٵЋ{ j�5�J%�*��t l#]E�.�ma��U�,���<�R���LU5���X���@H(�4��ۇL46��ܬ�H��}w��Y���'us��&�5u�5ua�2K.���<��-�`�M���G�^�$'�(�����5�nc�	���a�K���\�R(�Ůe	�9�n�n0Knh�����g����#n ����w����D�F������ ��P�ۚZ������xxL�ޑ���D܉6�-���Y��R�H;�r��ZNm=|f<> �צ�]��n$Knhې����f3�1÷� ��Wڽ:Aȟ��nc{��G�yC��𯼔��yپ.gL��`"���}��pn~ϛt(�	e7|<������w�z���-�z�2���;�#�oB0�lHMo��\�]g·斮����^��URVX��R�VPK�De>O޽{�[���u�~$���������d똜����E��[~9Y�Y����>~�@�D��s@��P �H���Hߕ�2#����o81$p��j0s�{�y�2K�Ï�Q����{��]'9HŅ5��JU��J�SQ!�t�F�QǷX���=�����?
�=�<2��x�>�#��M|A�t�!������=���С�?{ޟ��B�-��[s+��*���z���Q�S�����)xP l	��;�_6�H!�mС���Z���-��~��|�O�jꯏͺ�П�����(O�c��zh��v=��Q��3R��� ��h��W���n�m�x`Ǒ�G�"E��v}�����	φ����yM@��m��ۡ���Q��Q���'詪���
l�͔�5���`�;+4 Y��H�7�:8���� ��4;ޡ_�Aۚ����{3�',�n�=~��
�;�N�����_����nt[�$6�P-��F��`�_��x�ק����*7_��@���m)O�c��/O���q�8F��U�����;�ѡv���tj=�oH��Ϥ���e7㿄��:(��̿��DH:$=BL���=>�kO,��s:tz�����ڑ����8�&��Ӱx���h����!�x����<%�0��Ϻ[���/�9��L�N_=��b��VOH�v��l�1]�7ۇӯC١����<�b�-�]^5P���h;�K���E�\@�t���tҹ�y����uV�QsR!Ai�D���A��y�����ݾ�m�>���A�wW.>;�p�=&3PP:��Ͼ��9�aX(d� �'�Ð�a���wSa۰ˑ�%�E;���q)�v+�wއ�Έ����;x��
[N��z�v��E�9��}��8U4d�@��BM���;q<�xv��9V��!��nbT��7uHAKq_7&9��ȍg��0�7���éps�#p�'��b���������Q��zf�V0dcn�M�N�d��+x��H�z9�����{r�L��b�ں@���K��z0_=5���U�rS��5{���`{=���Z������f�ȧ�����67):r�N�bi��^;�3�+��Up���o=�4��/1�Z|5bP1�4���<�G�V'�p����)��)�y�'n�Yhd�UOG�_ݲ��D����CK4��ju� ���D[�Ë���\G����"�)� D9�ա��J����2��sp+�M�X��������N�3�>�a�r�s ıVN�MM�£G.I�y[��&����7���/�+�%��E�wy�����b=������Z1��ƈC@QFK��m1b1�e�m��&�+6)5Q��APh(؊ �fъ�&����X�4I%�,TccTTi(�jJ��4h���Ɉ�m4l%�6���Ƌh�Ԗ�Q�F�5�`� �[�K![��%j�`�$&EF*�V2E�ё*6Bƣcb��lV�c�5@�$QlTh��&�-�V*0&�cc&�Ti�A�э�E%�6-&�ص	j�c���I �w+i���M�˯���|���H!�U�m���U���C�k����_�H �׼��{3��Yͭ�:�+W�{`O�U`�Eߏ���zh������
��4n�����e��y����mC~����>ڄ��G������B�n'�	m�yh��ө������կ4-[�*��!��d53Ī�¥�2�Pf�ƀJ����������훡	����۟��+�/i��L`�x�x=��#{՛��O��t���+��m���|A�4��cg�<��G�y�{����<<���o���Z���΁?~�����}~1�s�'CR$~�P �鯁�܉4��m�l҉���F\,5~^-'k�ه=[���{�	�zh�����ψ%�4m��v�����}"�:�~n�^�=}\o�w�~��}�/g���������|�na�jnh^��vQ�ӥwD�y����8�zZx���8���b�h���!�s��a_���
���P��I��m����C^V�z�W��_�Z��ͭ�u�(� O��Qm��	�"��Y�-�m�r(�[�h1�n�wn�u(�,�5eѹ�i��Y�*L��w������<���ǂ�!�B�u�1��=>��I��{�/�7~��:A��
+�A����@��H_jF����zP�h}������b��Ŧk��
�<�?.�?ۮ���(��ܯ��U�z0O{���q�ۚW�N�Z�,����jSS9�ƿ
[��~ ��W͹߁7"G�6ꂿ=��N��鬖A�$��|Cn���C��޺�v��ǀ �yz~�����Ѽ����<A��!�B���A6�P�':�R��|��r'��;�f����'�3�x���H!�U��8��g�U�QY��
�+r����L�n;4���{ǵ^�<����:ګ�4nۈ�����O� ��NF"R2�"�L^��SU��u7J&۽kY�K�߳5��q7.l��;E�:�lv�MW��ku���&3HX�Bj��2��)A�j��2JM���a��M"�M*@1�4\�MYn�
�	
�um��Ai��beIe	]eъ�5�R;�`u^ڜ���bj{hp����Z�m�Hi���.��ͫ�ް"�TL��I]a�4�۴Y`���	X�cs4#��L]�"��]]\k~�C��
���\8K��F��i�����Bc�,5�!+�@rXѲ����/�﮳���7 ��y{�~��T�o��~��;�;�	�ǫ���{k��t~nD�۪�������<eOD�-������{���t{�Rݧ��ܽ?W��B�p}ŗ���|��ܔ�!j���	�|۝�����:�}]R���J��H���؞�����WH�u_t(�~#�xO����A{]}�F|A-���.�WfxxT�y7-�,�
�@�6*��+1Dm����w�@G�"A�nh�܉6�ٵ��1��	鮄<���t��<�4!w�Qn$�r߷ԯq���T�����o(J�̳#H�yY�aZF:�usq�j�mm�i^O����O�(�����=gc�z�F&}��د�}W/f�'2F�'���"Ho��?6�W��H%�?zHގ���9�Dxc��,���u��b���Ҙ9��l�?g�N]GM�*��]�A��5X��7&�l9u��a̖Ć�=��Đ~=�5�'ޮ�i���n[�Y���A���Wŷ%�m!HC��/UpB2@Og�_���W�6�e��pA9��ء{5�*�U&���x���)�AޡE��?6ء��V�@Dʾ|�A��Y��^����RlW�gxP k�tN/S�=�6�>��A�U�ޯ�����m�[t(���p9��}�it��]�Wg���r|ۖ�o��@=�'�?P�[sD܍/ޯF�ߨ�F��2f����v*�\J&Y���cθ̺�-���u�P�t��'ߞ�>;���t	���_6�V�h��y��{b�c���B�_�vb�����������Р8��nh��
��GPOJ���n΂
��+zW���3[孊�����ρ�$�߷N�6�L���H�q��A}�r+��H?6�� ^L���mW��3��L�l)[���^�C#�m����Y�UmU`Ն�,T�Z�윜�wS�(��	��t���+��������t��##��K&*������ I��(۟�7 6򅅊��U���������
��t7+A����y�x�����=4�s�9�^��N{�z4�_9�t>-��CnEܘ4��n�B3dO�>����&���؟������I��i�{���W#������؆�P��)]0��tк�G�4gkGP�"������_��(����C��P-Ă	mϿ'�]��T��o���	��峏�K��>�@����W���|A��mРKn~~َ9�����o(W˺EnV�����Sf�[����=?P��p�� ����!%U�|G.�@�� &�P�?Sr0Jkb��ļx�')F^߸Emk���r�P'���^�?۪���Qn$�Bv=���P����� ���yd����SQ[�E���O��v��"�?���m��DEXܻ?����ݛw�߄��������;�讟���ju�@���XY0����� X��P� �j�%��x�٢9�����nk�Ȓe8.�t��p�U�3�w����+i�c��q�h
~�_�A��*�R�1�>����gT�M���:�0�7�V�ҳU�i�Li��l	a�[�(��\���|{��&����<���<��|/\+w�᷷�lO�y��к-�'��7���:�mТ�H �����3Y1���3&� �AwMx�u��X٨��"����� �;�B�nr�ו'�u���H�E�_>s�p0���M�C�=��dO����{��n�Sm�v<?~���
��� ��m�۫a��Y0(��?>���Ș�qM������x7������]�"둱�(�s����|�` �ۚ�~m���O��ݸ��8�SX'���z��;����=^�O� ����,���;��\P��	��8;?���Is��e��巠�����8ux�"�wӼy���7N�����{8��}�Q�#�����{�l��;E���ߞy^Y���B��k�M�SY���I��ڑ4�]�0<LƮ��P�����׊��V��]m���	�!-#u[��#a�l�JMf��ųE���g�bz� �#���,�-�^���Pa���xs�a�$��.d#�9.*W���@�E�J���RViL�S�K��+-)P�i7V2��m˳��l�4aL�@��&���j�
X�4�fm�y�����Ex��&�5٦Rͥ�e�ʶcTn���k�R4�7g��{���}������x�W͹y[�˼<�l���lx����>�̔?s�{�O͹�u�~��a�y4:�|6��n���}ge�v8W�=)�^߅����"Hm����q�w[�Vw���m}j>�
�O͹q �no:�{�	��wAy.�'Vjc|/P?d�r0��A�Cn�
��=/��[Xg��r~C��.�_ۡCso�g�yVU���(����qZv���D��|yD��鯁��n �t(����[|�ÿ�T��a�����ٞ�د��>ޚ�I��mЪ��,��{sgs"
pjf(��ָB��̑�+�mXrh�wb75l4Ҧk(�e�0�#���ou
��	m��t{�%,��7�;�Xx�,�E@��9�?7"Hm�	m��=D~N�������7��A���7SܞˇZ��n�=P��mo��s_J3�N������8�3ѕ���r%��Iɻ�y����~��jt+so�g�yV]�i��q�=�k����Di�~~^X��=�5�4C��}�Cn�ۚ ��D��S@��o�vr�d�ғ5��xP'��@��Bn��ۡ@�E2�;�vo�t�(�� ��_w���5�/�X�zc��^��}@��f��M��C�y�D����Kn~��H!7��s�U��}_U��S��}�z���M>�?v��A?W���s\)O�F+��w���oLl��WJB�CQ�1M��v��Άs[-�r���bf~5������)�|۝ ��Y2�G�۝:�W�D-�(����N�zD�:����n m�X�Kv�۽�ؐA)�����c���	Եxg���}� �=΅|[sH��9��@V��<�h�r$��
��ۡ����}��5I��iEb��Ț���Z���_sh_M�ۛ�{'�;�6����8t�VR���@�1��f�VZJ�Ŵ�}N<A/T�K�_7`-���m��#����L���J�{�D7~<�S�xy_�[��o'��?G��M��*���Z����E��~m��t(�F_�9==�}�
�M}h^����͉�Z�3��xW��}�B�-��A��'>���w"A�Bc�A��I�������-� ��Evn�')�Q�t0�+2h�&�O�g���l��������+�]^��wkSO�G����.; ��~�w�_��B�>蟈%�4Bn��p$��l�F�Tł�M A] ���
#�+���7�<{���zD��������񩑧: ���n�|[� �>-���{�z��9G7n<�Nޥ��~����Qm��	6��j��:�*٧+��rD�����!�CsEg��~]J�^$����?=SDw�J���C�Q�u��Z��i��1^xx�}:+���M�����Fe�`_E����B��uEr�AG=;J�%	"[0I����~B�'�6��A��B�m�z�-N>����a�̒�x��q~g��/Oˠ`!�U�mЮ�R�����O��"D4%�Z閵��6t��\J!�nC\�#�,�7�.�o�^���鯈?o~�E��A)�����<�=�;V���{��x쥂��v��#�_7Ӡ�܀��@�۟�uy�7sӞ�澤<E�����3F�{����ۊ�I���� �jk�����;���^xGFĺs���~u�O��Cn�mΐ~nD�3�i�ܫє&����to��g���y�|A]"Hm����q�l�n�-�� �ۯ�� �[sC���Ͻ3j����b�
�`Iv/|o�֯��`�܉���P?����Cm����ҟz�{��J��z{{j��R]̯�;z�<��r�"<�/�H�ֵ�km󵭫[o���kmխ�[okj����mZ�}+[V��:�խ���mZ�}�[V��-kjē��	G�	D! BI�-mZ�~u��[okj���mZ�~���[okj��׭mZ�xk[V�߳�e5��;�  �}�!�?���}����c�                 @               h w�   �          uC   ���E��
�C�z�� ��=��=4����/1�ʪ/\>�ԑQ^ƫ�O@���  �/�J5��`�>�==@ǔ9�b��w���^v:=45��>�+�FZ ��   �
�)�%��٤���zS^vN�u��:nYpz��Z4�ݜ � 2nܪ��K��k�v7f�m�c��Z�tҚʻ:qN� �  �=Ov9V�E���!ݷ��]�Md��T�b��[oc.�p�}R�{JM���>�z4�[7�A�{�]�� P�>O   ��}CZ( 
ì=z ��g�Pv =FZ>���`���     D����H       "�����b�	�2i�# L@��7���g��       "{R%5 2  @4�S�!2�$�0Fi��i� ��I��dڀOQOz�d�4<!�'�����XO��߮ƟW�AG�j��0z����O�����	�EQ�_�Ա  ��R׼�����o������v��H�@ Td��'8@Q�D�$F�e�<�v�:�O�����i��?� *<{E�c@�i�4?�y�`��`�~��[��g@�`�C_w�-<}�{li�U�>��EN[��N���}�F/CNR*�KP���Y�-Z���c�c�{���Uv`Q�eX�vw���//.]��]�y�5f��=�f�i@�Y+�=��G��fVtQ��c\�7]36�� ��r�ճy��K���p0cf=M�$nku�t�0�g����'.]�p�F雰4�:�һ��֨X�f�i��C�ۺ���
N�4)�"�1���%3���Į53�EwY1�u�yw,a:�X�u���i`\|��0qʖ<t�P����w��� ��](34k=(*�*��C*!�`��q3��cr-Џj�:��a�0�F�<�h�6����[��y���B.Y[׿
�wl'�Ӵ��nC��M�ε���>�9���O��@#\��Hͷ�v����!y��>W۹�q�{���vabǠ���x[>�:�)Nz��!;J�;��r�
`��}�g�=n�b��t�95\��178ߕ�����B��;V��"�V�G'�������(v��G�;ݚ�G^40Ǭ���!�3:a�;{��ۛD��^��h���.���b�I�e��G�V�s�S�Y��@��̭y��^1mݭ.X��) ��;�vp'{/%��G�:��ڵC�9mߵmN�� ��u��ue�y�*�I<�H�7��ե��kf�=�;����-Qy��N� ��m)ѹ��Jj΂r}�L��>o`KH�I��vpJ��+�x��Z��'V)��NBl8��#�d�2�Ջ��jL����opL[�^8��+۴����B=��>�{�
u�ȣw�{��q��rg�hZ28�t)�6����g7���dx ��N`�#��i���[³�M�0�?)Ê����vA�;v]�٬��i�q<w�HMB��rb�b\�$:���M�t�	1�o8^}8=�eL��u1ݯN��،ڨv��4�)�Ep)�W���s�l�V�tZ��C}[hZ�!6{z��u�Bڲ�A�0-jc�|e����j�����]B��ın;���ڌ�U3yreu�t$943fS�9k!�X=�w���ߎ0�5}�7[;��\.]��k��GЩ���m��Y����Q�E���3�VY��;qd��Jg*����i���ӹI̽�w5f�����&�m���;�E\x�+��)x�����L�*��[�c��KJ$��r���1�o�N[�
���
Vn��+ln�i�"�nhG�w���:ã6�9��(2���b��J�H9A��&w,�OsKCzu=E�v�4�,hO+���ܒ�<;���K��#">�J�4;�d��8�LkR������+gU��z���	��X9�*U��کN�[��1c���>h �I�-�+�l�0>;�ja9 �
j�bw�͜b�f��>��0B�@GD,՜�(ֲqE���W������v����GaZ�`���1��unɻ�R�8�ZY���n���u卙g�i\�����s�	س����G)�ȵ�s�˥3H��$z��0��J���W׺G�cc����od�b �h��L)4��E���ЗP�w6bX��wͮ5��i��p��Q!8���p�)�ܜ��7��;*��k�s���^�x���4[�����E��b����\�[�>��:[�]��۰n��v�'��r9�ɸ�k��xT�*y����uܡ��X�)wU��<
�cA�%���g!睭�	������0��b�\[{�.<w�>�sah���-B�l�k�+��f,�d,�oBAn �٣��I#��:�U o[��^��w톌j�{�����������u`F6ovu�k����p��v�lJN»l�>��T��{{p.���)�ˬn��S@r� 	GBs�6�"NE�'��v�`�Ocm|�!Y�3^?���h: ㏶�A�5�p5 �5�j�p�}ܰ�w;t0Ü;U�x�}=㴇���zd���ؑ�g]Z�lgNMs����q<��Fvl�@oF�9.�Q��Hn�ZZ�p�;��+S��U9�h��n�=U��Fճ���$�x��y�`�=W�����6uǔ+�{L*xw�fώX�+un���)y�c��Y���D��渽=�4ŗ{�饗n-��ȱ^�;P��3mO
�q}ϴ���cI�mU�ǳ]=y<�Z�_�ݗ�"�Ynpgc��҂v�
�DL�5�]
�ۮTN-��wu��'p�����ӽ�E�Qd�c+Q�:&�L�����-�sG5Ķyo.��Z�
5��+���� ��f�ҕ�jB휰՝������z��"�$��;�@oK������aL��P�ig=�͚8��\r@$U�a�n"`�Z�-k1��׍[���8;�vۧ��6�Հ䳔�6��A;F�Ȳ�}���'�F�oF�%�4ɓ��$��Bf�͙��5��EnsuEX&�
i�[��wz�P<$u�H<�j�Q�.'�^�jp����vs�]�tAaD-���J.L��>����9��&��d��A=7�,M�����Y�e�΂��F�1J2�d��:s�>��ƌ�s�f@����t^탙ם�C�8�E��Uf��6���(Q;8�y��.-��p\�f�(0�q��4"/���b3+7S̕�sI��R}�VP�[��oCt�8ۛ\VYe&���q�G^q�rk"��`�fA(���ۼ4e�4;wg
�:1V�1�M�uk3�d����t7{�̝�p��_v�� ��ގâC�޻q�Ϸ�.�4�����v#t��%՜5�s�����Dbe�m��cuem�[M�١LM<���80K�E7ZW�s't-�7��6!lI�����b,�V�˲�3�������hĳ`�vR�O`E勁{��3C�Y�.	� �o7Tj�.�3���ʒ�yoA0�Q��c!c��e'a���w��;�{׻���.K~G�8�Ͷ���ƽ7Wd֗t+wL���6��q���'�>��c����/��h��!�����OQ�	�翙鱞:�����C��
%   �@ ҈� �-"
Ҋ�RR�Ң ����J-(� �)H""҂�H-*�R�44��	J�P�H�P�P���-(�
B R�@1(�P�Ъ���
����|zz����Ǒ���Qy��G6Ν�@@ٷZ
��'|�#�	��
����������LǗy���Hb��J�bͪ�/"��y��Sn��������'�����R,�=hB��T�`�[�K���>��B�{�}�y��{�f<���P�{��Q��p��p��lNd�<6L���2)����h�ὭU�����=ޛ���#�������܄���&t	�m��nOo�֧V�j�����wP�aI;�d�d��q=���v��!L���EWp�w��5�A�[Vh�5n�{��@�ׯ��d��\�M�n͙�/vu0gn	������eD\�`{�w�x���7|;����e"g�3���.W:�|�|=����]�x�@��]�0u���|��zu�ձ�wq�"�g�~��s�u��Ɔ���wf��P��|~�D��칺�g��C��E{=Oy��t�I8���õ�S���������E��fj/y�d��LX׹��m�n��='-��4x_Q�M}Мy�{R5���z1A
�xc�{�� i�-z0N�.���Ƭ��
����=޺m1���'^:�!<�����	���Ō����#�}���{�[��f�;�/��;;�����/K�k�}{^����-(1�bxjK�l��A%�7�A{�
[�N����I�1j�}朙�8B�9��7ug7���c����{�LՕ���<
�;r�R�B��G>�v����Q�*�O��i^ٳ=ͱ�/�����^��R��Ǳws ћB٫�m�[�[+yg:mT�j�L�*��7	9"�/[���@�����7f�m��؄���Mq=���ԇo�@M}Mk���u���C���y�<�Xs�����}�q��;^ݣ�W�p�Y�;����=��z�r4P��}�V����x3G3��3�7G��a1-~�� ��|�z"�{�(4�9o�~����nN�J����ڼ|I>���L_2{�Gw���G�wvuͲvn��k�� �gG��~�
�ʏ�%(/jVQ�6�=�p?n�0u��D�G����.Ճ�;|
|�{���"}�[8���n"�w�vr���s���.�
����}m��.�잶ӾXA�!����=̉�˫X4�=����	=k��^ɝtp�u|g׺�=���{ݷ���p;�r<]&F�0N�n���|��� ��rI�����V{V�:����j.d���2.��6sc�Oh ���˽����'�b��.F�d�狼�xq%1�ދ���>�}_æ ��ͯ\>��s���=sІ:!�1�n��ܔ|�n���#;��b�/^���(�u^wܻ��%y�1���v��C�N�~4\�x`c��a�TT�Rgc0a�v_{:=)����}�P'-�r}��(<�g�Dj��<�Z�+�wiU�3�g]���{�+	w<sޘ�9Tx��O%�vL<����s�b;���(<�o�������-����*&�820-zSq��ٜGV:RVN,��,ZS'������{�^ݾ%�3F����2s�-�9jK��Oq�a,��`9�KD�Y��{�Eu�耋�n���)ˤXۇ�M�H`~�س����}�@��\����mmՓƠ�^}C�3)-�^��}�w�	�>�;l~�g$���p��׆�$Z�����J�v4��}����VK�čp��������ˋ���\���>��E�8����s�=���G�	�K77��̄�I�CwϷ�S#lsN��>���O��9�m��M��w�owf�:�^MS���rw�C�ڦa��7�?լ���V���/2x�����o�-�)G��{˴t��F����6hǞE�<7����}^h�{ȴ5C���)`	���}�z���[���D�{P����6\g8�-�&o���;��l05��˿)�&��pAŻ'=��tk�hOL���>#k�6�;��]^��L����7:M]�5�cɕf��u'�|7�=c)Z�u//_Z|�ha�ϥ:��zf�A;Ǜ�|�X�;�z�z-�g�Xo
�S(����75yٛ��_O��s��w�8��� ��/@��XC{�(ޏNo��Y����r��S�Jiy&C�k��I�����"�b�v}������_��=���x5��-��~�>�6!���ᓵY'�������Ε����!����ѷN�ΞX���N>~}�FK�*������ׇ_a�1��}.ub	V}��z���ҕ�����݅�������}����O���2o)�L3�a�2,�9��P�G�<�>?@��L�О՘]�f0�_N������7>ân�>�g�U��wf�6�v�ɹ�YOj[�K_G�����A���B�SB�}���ۍ���>�G�E��ž^�tZ_b�˦f糴t';ޘ;&�߸w�����/One2�^,�|����f�q�|`���Ϟ_�J��˪��\(���w]\|k܆9�s��ݬ������ze�=��I���s���>�N��z/�x�k�i��}����\+�)�=������w�1�� P�(o7iG�d ���|�\��T�*�b��A.��ҳ�G���H�a��٪�C�8}=E�r�90=(���6�=�y���ҼK~�瓉b|�m��'�o���O�^	f{Nt3I���'��)�!'ďj�H�;���\�����s��Wcx�gnf�`�L����/�{�a�[���� -���ks��&T�ש�d�Һ/�c��φ� �pM�Rw3��S3�n�[�Ql�}�=���ǻbZ�5&0��߹=퉙�n.�_���ܘ���۹��r��o���
Ո�0�����xa_8^]K�<�ۧ��=ô���n�Z|r�\^���Y��h��t��~����0C��y�6/0b��zXwe~�U�e|��<$|�9U�1�Ky�f�ٻ��G��Eݙ��ά����;�:��ú��&{�:AϦVצ��<�cԁ�1j�ע���Y	g:���E�XT���GG�g�1���gm:�=9v�T�+�%���snssW!F<8e��e^{�S�λ����Z;�=���e�����N}ټ��-���[��+� UE ��~�9 kT)X��C�G�v��;?>��g������n�W�O���9�:^
�6�Lfɣk�/<�GYŷ�gvա���2=6�r�e�oK�N���[�Q؋��A۱eyqv��T��n�9��u�^;[�"�j���7n�۳�K�^ݦ�"��cp���t#8�����z�
���s��K��-c�}i9�9����q���ڌ�'��i9M�Mf�vL��s�jJy^s�aø�����0k��[WcO[;�mң���3�O:yw�e��s����Nwg���˓d�g^�h�v��W��PM�-�Y6�N��{Ӹ��er<sp�k�n�X;/m؎f��Kʔ�E=M�����v�i��+�4��u����c����8��W�:�]��-{/�U�+Jr�-D��!�	7l��� uy����ݸ}���6���������t`�s"���$"v{q�ksQ�Dl� Cd�V�!F�S�ng�����m�9�r�.��k"�9��dO^��z�]��5!v�	 ��מ�q��5��M�󽛤��!�Nk"��g��6n�����u������O7��&�ࣧY�Y�ܝ�%�����|�1�0�8��10H�Z�+�7k�k�rp�/=���Uq�����_[���r��rg/g�gU���\��q�糌K�xyі��eݞ����;�۴b��u�{N�&�N��A��A\S����I����<	�v�Zۨ��v�lcY)�%�اq�n����wh O<�9�W(Oq݋������cv���7h.�i��9�5�[�AEڒ�����9� =zeNc /fȸ�3�9����a��]�f{u�-�fN1����$5��9�Aq����7X�Ca}�b7I��W>���\����z����*7���l��c>�1����=Ůp���r����$�1u�=���LI��n4gn��8&��������󵫌��C�U�w�/h����x����'K]�&�����J�m�d�WFJώl7nH�s�U�[�Sn��k����/�v�[�Ny��Ǟ\���ۊE��:y݇a�zό�<c�s�[Z�=����y�7]���a	-ֻk6�<��B�4l�c1��':��J)����������6ɍ�r�vm�Sn��.W���qn��[� |W��>�����wQ���@�
�S��|�[v�o� 6��.s��+'jζ>|>m�v�pz�gGAҁ�ӵZ;M�k���a�G`�\�9�L�4$�b:�Nݎ�k{Cܛ��G�\�^�H�8N-[G��J���k;,Q��톈�;��4NN"pu�tZ�5v�gy�݋�K�-�m��8NݸU��\��1���D���ӃnpN���e�b���[�L)�ն7%{4ɋ�&�n�"Y�M/g��rn��v����1�=�w��vd<&�A�:�ۧ;5kt^m�v��^\��iފ��˷_�~l�yN�U�vx�;����������dO�S�`������Z�N}�L�:N셶gOa�nA�gB�#Q��5�^��ό��s��]�\O\�Onű�պ�VN��Lt7����guK[�x�u�'�X·�Ӳ��G�.gk�r{v�:+K�ǲn����<�mV���d�㛅����1S؇ۗ��ڕU��7X��s�ͻv���x�Ⱦ���a홮u�j�i�v8�тcN�B���g�[nl��-s��٭�;�{\ݹ핮 �m��ݱ��;�-=�����h�]�`kkҬ����3���OZ��vKc�������);QE!`�n��պwd��φ�=�'��[�/Gl�آ�u�B��{a=�n�������'eۯZy*IGlr�tY�nlsG�Z6�ە������n32h�v���4�[�i� ���h��n:���Wj��3��w��s�Ob^�7���o�e��nȽ�r[{�����ms�صN�=��W]��w�G^�v}H�W�M�
w\��q[nA8<ӎv�ח���s@����u�F���&�05���z���S����V��|�R���:�Żu�u�����6u݋[�3�d����ZH�Wf�Kih           dܹF拴     MQk%    �@���V�     5MѮ��+;h�&َ��G|���c!�s���U&ӫr�וnF�BI6�Z�Ͳ�5Mخ�v��ᷞ��ݽ���o�^��i�$���F��" �F"��Y�h�JJZJJV�ܟs.l�SI͉��a��(���R�+"
(�.�8� 8�����7�`��ALV��-ZZ�R҉ ȡ	;؜�Ѥ�MR�i��D!@�%&��4��4����pa�
 �X���1&���^,�M%!�'@���S����������Cۗ���m�6�6{:�{u�pj���e�A�l�nxz���H�l�>���:� S�yU2ձ<m�Vɓu�/�����ihˊ�>u���i���&R�_k�>�\���W:`b��^6�k�f��Qų���tGN�B�i�z�f�u�%��лsy�kt]��2-[�<\��8�8���cȞ���l����q�3����3lZ�.���D��vx�v�g���OT0���v�3) ���h�1����enѐ8�v��8�86�t����C�<dK��^0yN�M���|��ה�[=knX�K��o'-�2�-�Fŷ=��c��O�m�.Lżs-rvpg��n�L&ڹ�������y�e�����8Y4S͞�n#1�ָi�[7���%  &�J  �� �n7&j䵍e������7�8rr"��*�v7��@3����ۗ>���<������c&N�8�#�ll�UW���<�&���3���*��v����?�̈́�{���5���fb���������>[�1�	}{�,�&L��P���G{_<q�( �+�J�&`��~����mj��eXW%Z���l����TLX�$A��>؂�x��k�p�ǯ�o����]ў��1�29�D����\�!�����p�:R��_t�f��
B���R�9�L�Ø���8>�/f�f�Ʒq����U D�	,�;��6��D���6^�;}����;�Y$��T��ro[:����bKL�ĒB$�%#(��/dӬ��'�����>}|�����=����	'��]��-6ww[M��BY�Qw7S	"��E�2�@F�ߟ]�Z�ozv���:���R�0x�����W��E��g�1i%
0�QsV�����5���gz�6oH$����6֛���ڔ�w��c���<L(�Y���!H`%����i��{}����d��M�j|�Kjvl����5��
�ij��R�����qOsm�p�mO���W��}}g�
������.�*�Ts�&�Dɔ&�l�Q�wv$�Ǚ=��.WQ6z���n4*���}��|������oQ���q�Ԍ �D�^�µӹۜ��*c�!:h
��,����ֶ"�\%�9�W>A%eOh��3W���ЪP�	�����
��gn7Mܤ��l8�nP�!%ѐ���o�=R������JS:ӊ��"WU^t�*�U�k-��+GI�N�v�̳[�o�v��>ێ%�&/�\<Pr��u�2���'gztv��R��8�p�.�ػ1�X�C����vͶw1�mq�rS�-���c������<�骪���߇��q/f�4,b:G)��@��T�<���x�o;q�zjшA)��/kwLX�ӹۼ黵�:�7d��Yn�sb��o6��!)�!�Wt!-yx��~�z�7�4hJP��a��S�ۜ�ù��y!�f�4ծNz��l:zŭ���h�쉮K�G9���۾~�w)$��s!T�u���ё�#Nu���x;GE��T�����]uk�7��J[5�s	$��ç[���b��̽��ڡ�P򲧻7Z�������	#	M���Ю�V���w�4<���8�D$B���jZu	��$�U��I�#�M��n�Na�����ę��I%��~2&���S�����i[*�s�3��AJ�;9��S��p	˘w]�(�r2v�^��EҞ��յ�"�%����QC"��v\�f\�m��w�I[z]�!� <�9ٺ��z�%0���~���ܼ�I�n8o'a#59�%4��>�v�D�F^Io��>�]6��v��l(ܻ��J��=Y���淝�IR��;��O��7��[r)�i_X������Voj:�^N;GW7��\ȸ.ބ�$��@�g5����!	X]Ӆ��JR�'�<a͓��2A��D|����鏿���g\U��T��1$�
�h�ЈW5�x�o;̺����!�bSn��]�5ۼ֤ZSuA\�L�(F�-��ֶ=r&E$a��#.�w��x��X��RSԧ_���"������`~Ը����8�u�ӱ��ĝ�I��;):�m��:.�>ݰ�h��A��B��� ݣ����σ@w>��Q���n�0l�az792ّq����۫6c ڴ}}~��b�qn�s��V�Dͽ�)O)�k�i���8,$�BJM����汻J�P���YG5������z�$������b{N^�sZ�M3'�h�$��܈��*�v�Y�,%0��e6�sdB	 !J�2�B���'/�%	Om<O���:�֬WN� �����$�DU�]��f@9�tHư��2"�<B���w��e�����ق�쓐�a�XO�����ZE�V�ڬ��SKs��n�u^�d��($�@Ukwg3�Zq�4��_??�7C����lZ�/��+�$V"�	�v6��D�=���!%1����s�t�������L�a��W�^��>��G�>�?a��eW��r��t��r<��d[�����e�;M}���8�a�}s��<}������}�Z�#L�ox����:c�Y�e
l{�ՙrz����/��Nm-r?u�\��9?7�'П�Od�vI�����Fl��skxN�>��M� ���3����W�tӜ��2w�P؂?5�_%'ް��u}k��=�ɘ�p���\Xw�G-�� N�սod;�7KY�v��	����`JR%�\\��;|o{�v�2'#"��K�a��^�)�����D��:�ҽ�����tG�3��1XM�.*��)Ƒ�i-gF��f�SԬ^��3���۞���K�a�M������Jv��%=��F�D&�F�&���L�(�R��	N��К�k��R�WV�������Z{�M��H�b���4�AJ]��SJ*B��(��8�3b+�Ua1\cET5R��1U�`�s�)E-T�4�EUDEk(��%��󈍅XQ��k��Ҕ�]ݿ���CHX���,���<�鮊>���������}����P��:Rͼ*
Q2�@�jڥ:wg��qW������|w��{�չ��X���C�8mVIŃ�2�=��|�ҝK}���轔�.�E�ߏ?��W�©JR�I,FY������_o��m_K����u30����62�Eu��2��o:#8A�@�4]؛���>|Π�������_ߕk��P�[B�c�.>�g��؎�묆X䇩&^CR�ھ9�{��a�Ts�I�wy9�����?mM$g~Wwa$R�����9ђ7����y���Q�W�͈�䧖�s������yTM�	'BY��g���?s�ښI!�# ��\	Ŋ��;�+.LЌB �`�WeT�
W��D�ED�M��n�8���ݦC�g֭y�Ȕdn��g&ۧ��W5��=��t:�h�v��o[��7v�c�q�ұ9�jF��wl&e�2�(
��~~~���P�8���Ol�(�P$�&{Gb0�����f�Tf�?����S��s0�3���o7��O�}9�$���u�t��o����ЄVn ��kW�-#���ƛ�8C0��GW�!�`�y�jo������T��ߣ��3��k���SP�׫C7�1"�����s�����
�r�_�&K���LotVɰ�b�v�Ȩ'�B6�F��!%����~�G�}����?_n~�i��9�]]�{�(Fd�	,���:��*�Z����}���y3S3/�t~��j�����{u�����.��u(BJU�*]�kf��Ił��KK&8� �9����x�����޷BM>��5�_F���a��5y�=���ۘ��>�+�a$��{9ZΆ���N?x._�#~�*n���=Z]��\x�u �o�X罹���h����g8CY0$�9�^�]�����(��\hZ����������?
/p8�9�y�}���̀k�rD���D̀g8B�lmѯY��;�nq�]s�} f@8��"[a �EU��J[��?}�˸�,�,�%�i�ֲ�3D7绻�{�������(���h+M}����~����"s��nu�w�����l!��� ̀g86:�s��H����0���~u���$��\�����QDB� �hJCxH�p��9������;��w�s����3 Ƚ�g8@�@��;5�m;�@�"g|4Ubh�jw����x7
� 8��۠��~��g�욇cc����GP칞��K�3�j�*���"#��G�=�`@�@5�u�>$L��������aN6��㾼v�̃�r�����`1 �@�w;�}���#`���v+l[=$�����hW(�@Ԣ�4�o�s��������F�}���Z �E������ Ӝ�ƨ�H��=g��<w�@��DF��Th�䢉HV�(/=o�l�����g�� ���h�CZ�����}W�kZ���~�@u�{��@3�ȹ�29��Z��m op�1 ���9���ޠ7�{��#���x�v@1 �X9�(�s�0s��u��:���8�{�� �l��"o"b
֥�i ��e��K�ݻu���'�nދ�����le�$[�e�o���ަ����ATJ�����|amի�e�Pr�]�t�^��%
������Ǟ:َh�|�.��=�k�%ڍ����$��������k�f�\j�̬M�6��L`P�?���~��n��nzv�9�t�䇩�wu����{�������wwƀ5�@k��=�������ARa�����1 s�Mdx�ă� �p�$�i�	����_r�5�A�|�s����y��@�@9��Ȗ�Ď`-uێ����������x��"kP�4��"h����=��]��w����-� ���B���2���d4�:H�@8�t�9���ێ����d�;�1Ń=q��dix9�i
��i��!ZԠ��(+�}����w��@��^��:H���#� �q@k^��w��%��	d��7�ݷ��nK�mq�Th�>��MX��s����������(�~��C�dK\"b]���dHX�CH�(�7��f��km��~��r��w�67��׏�&\�zq����[}�
"J�	�G�s��n������d� �l"w#���,h�A��m��s"F�D+Z��V��g�����럻����%�8GBD��	���֡@i���k����@�,�4��d9��\��}����JC�}�Șl���JRP�62U�r�����_�?�=��`�Q�n��I�)L/$���ď�_Y��z�Q.�_�L$��BЂ��ʞnsV�m$��H��6q���ߞ�&ᴁ��g��<`���S��Ϝ�s$ȼ�W	���DD{�y���������J��+�X�v�]wk�Ƕ�D�r��0��6�:U��j�ܥ(��w����>ID�$�a D��LD��$wcT�%ʻ��׮r��F��!)���n�_k�YZ���[2%]ʸ���x��oosU��Ez���䑁)�X����5[70�'"dV�х�TM�3*svcz�f]U�G�� ����@��\w�]pk���k]x�}7���>�)+��/�,"bT�2% A�
RJ
�R)	)RW�D�ȧ>�������yI(J`Ah�]�iW�m��+�J$Z�V�"��O�$��H��ÝV����e@��B�μ�mS�&�U!)�![욜���O;�6<��F�5���7c~�%M�Am�E�).��j����륩y��QN�%�s>:�ӨY����*oM���zT�m�^�)��}�Oi�9ɬ�O��xYɃ�h$�n�\��d�r�2g����g�=��1�C�VW�]|]Q;��9�6k9�����@wc��zw (�[9xm��,e��>9ᶦ�޸.-5tS�z-�!�W�\��S����g=���� �U����i����r:�,�����=a�[�ZSv�q�+oQf���ǃND�x�U��_y;,�v
n?p�òDw��r^��<�%"�l��<�q�����Jk�-��7�m�ې|��#�^�?1TN�B�P� ��,j�*��
*���k�Q�x�ŷzHD�L�g|&)��))���HqU��D^�)ƈ:B(�-
�V�v�i.Ei�@V�V�!"���B��L`�(8�D@DmbZJ��������iJF�&)V��iX��LT�
ĩ�14�F�LCCKM)J�ESM%A<J���X����)
v����Z)i��
&%�/nݿ?�����n���x��|�m�M<!h�n��L�1�X�nȩ�z����F�h�6�h��`r��;<J�n�x}�{�q�fNQ���e���C�i4P����z���mÙ2>wp�R�9��C�[ucC��gm�^^M����у�r��Ki\mӸꝨ��\M�.��Nr�g�������F6j���׳.�n/u�v��^��=��N�C��ù����"�7S������8���=i���p=fmggp��=�w"v#�������qH�W˵v�=,C��Xݏ��l���ۈ�g���񡝶������p���5x�`�2���=���$LT��W\�ر�\s�]�l��:ln\�Rշ0<�"\�A��N��{)l�a{,��	�Z�v��k;.�\k�o8ٮ6:��Ir�&�%�۹3q��� �f� 
�F��,�Y�����������K�����b#�ӤBN�e��v��l�O9�k8��:r������P;z@��@<��W��[ی��fR�E�:�u֎N���8{v�Kc��5UՋ����v[q�&�I6�n�D��eDJI��;0��սßW=��,ϳ�/�F�P�7f�aZ����e4�mU�s�JR��wl�,�׍�V�	$ᬬ�S�[�f�ok.;fSۼ�Em���R�O�7[Z�ZF��yQ���ð�C�e�p��C�$�ބ��o�s��%��6�*>	���F�%s��uVFIک�U	#��mx��`�l�\g� fE�y�F�u��߻㸍u �͈��(��[���\�>J\�V�70D$���]���:�f�$��A.�",���7u۬��9���ۛ����i3�@�a	�F& 	0B0�ɕ&o��+���s��q�t!7i)��"{{{�e�N޻mZ:{�{a���}�鞟��+gs�2��;˜^��B�)T�M��F��W���r��G������<.�����"�I
��p.��
��u���4s�yrU�y$�('jja��[���W(y��P�
J�Ya�)���(ͩk��W����.t���jFfP�X�wy���wNr`��BMk��]���
�A)�(o\e�Bķ��u=�/�c�˭˻���q���˾�l(��7�0d�K82clA�6�x<a5�n��k:믍pMA��۟~�qb�>]��*�8^�
C�W��WK�	�F��~���t��i�k�17)��A)�cI��{{f��k��1K1����4����1��p�wg7YN�D����hԸ���z��;e�z㜥(BI�Q/w���_�f��W��ސ�kf���ݎ�Bu�UJ�����ditj3]Rs�������������.Ic90��b�үF0�z����[�'[�������3+vtp�ޔԨx�!1۔�m\h.�8L�M�:PN�\s5UU٭�����O{[�5����z5D+>��"�]}��c�$\(��I`�X��Yo]�!Zy�j�u]����������$�VH�����fv�u��g>Y�P��Z�u�U|u��M�0������7�䎸�Ga��8���h�G�Ce�گ��ߏ��_KĒA\9�zÌ���j,*$��+np���󦚶b���Z\��G������>��{���v�c"j�*�����̼�ޮ4KJu���ڑ��[����v�铓v�P��*v:�9;ٹ�����Q�����~|����z�8�<��eD�Q���$��-��W�7>�O���Ihu�s���o]�9}�J�o^5��2R�F�|��=gM���w�pv>ӡ+��#;g��Jw��Q���D��DD�Dc�I��_E�PB�exԥ<��v>t؎���݋	J�\N���{Ա��Nk�)��_)b�B� K��6ۇ�k�!>��w�����5=�{��99�E��h�S�d���t�W*m,�3VRG�,�gI�]}�s\PA$nw��&ǡU��u��zP%�� �X�i;;�2�.�N@=F�s��"k�Q檁J�k�_�Ɏ{��~��x�^u�u�<�z�2z�A�!J�	����[I]kա>���w�_�_�.w��ko^vee�!)��i���*窹��o�ذ��m�z�%	9�P1��Ǯ��BHΛ[�F��U����}/\�ݝ����P��E-K��6�<����ZE<T�%�0u��A�p��y�ü㗡���ֵ��UTy�)h��-��ۖ�wm��:�xS�b�k��g��WF.��nl��>K�m\�L-bqo�m�+�
wOl8�5觗��Xs<�F��`-s�ۙ���F������i�ݭ�r��$(�b&J� ��j�I&��<�t�OV�w���Ѕ��x#-=������n;�z�H��r�O�{����@�M�>�I���������J�%)$��&{�U�|��u����)J�Y}ƶ�T�����pi�V�g�TChL��Z�n���6��r�Dc�E	7�l%t�P���+��b�h�N��nQWj�P- =s��{��|w��
��7�5yg�(��t��wWoz_��I$c�q��Va]Umv�>�`�і��,eͩ�I)�"��N��]?1
�%����������k5ƐFe�Ȃ�DJJ��$�j���m�s��9)J�k�s�}}<�Wn��v-)��Þ��Ja-��c�V����f�E�4{{��g��J��_�n.󾬅
�ɧ�!��ə��zzu}��Gn���5�!Ӽ��ǭ�u���1oZ ��eN��:�h L�e�d��`�,g��槛\F-{��.��=�}�ikĕ�_"=�7��Y�f�A�Ɍ-��#����;������B��.���K�s�*Y������t��p�͜z���G����_��#zTg3������m��ӕ��ՙN���+���T��%r������??~�N+�-�L�v~r��6/h2�����*���;�������;O���`����b��FM�fiRKǷt�7\�!���v.ۻc���]j
ZB���\SEP�5M
PTMU�b����bjj��0�mT|��i]��
��"�(�T)DQ��ܛ`�UY��q��{�IT��Ehԅ�DAUMnK%THƎM]�"ɦ�I�74y� ��mq�q�b�%;kiC�[��"Fc�$�d"�h
� �G�ٜ��V� ��\����nUs|qvm\Z��)I��[M7���ϟ�z�o߇�~E�O+ce^���"���Uq��u�u�~��Cv{V���B�8���ŷ���xZ�k����$PI��
E������BR�� �T�&ro��p�]f�S�v~�I��w`<՞�zX6\�!];��w7ɛ	��J-P��
��s>��R��K�q_!;__�ʻ��=j�������c;v^r:�9�n/AB�*L��|��n��ϻ#�G�L!%$]�x⹾o5�cʔ�ۻ�	#	tZS�sU6�<ԗ�G��E���Y���8�S	L%��u���7���I\�jނ^p�!N����w�⤾�x��/�f.Ł�]�G]�u+B�#C@SI%ECCE4AB4�-"�P�CB��HЁJ�4JP�@�!!BR�44�B�S){���~����v�1���l��(�<�]W���ǵ�>Wm[���8Ԧ-����h��<n����o/OI�v���D��ax-�.y��5IɯUU\�߿���t�t�[����J�^�)�����������m��'�fg�������������Ť�U(�#��A.�.h�Ok��������}q����Uͱx�[���JV���Y�ś���X��U����?�m:=Ȅ��r��T d���1JR�Y���3m���f&&dϹ�u���z�s�Ґ��;��#���k����� ��Z�*��R�������J�u�}�n�p�ٓ���y�6	�	$�N�-O�_s�!)Jq �����T^�m�����HzW����չ���\�������������g�����B��LL(R�"���0�S�׭�:��aTe���"tʤv+�W�gy��
�
=rѬ�0�*2���ֺ���2�hQ�g�wM��.b�'F��>���j2�����h�	-�swib���y�)���WV��!#���^o7�����P����^���kq���Ja�#D%+�'�co�i�	"�\����W5���8�in��q:=��� �EN��V�w���pU)L%=��m��Orf��|\��Gy!�I>�u��2�<3���a�5W�x61�8����q腕�%0�V:�+����yQ'^BY����~[��dz<9A�qdt�a$Mx�����\��8���������B	�RJ��f���2�OFf"N(@���T�y��*�n�JS*�<�x�L+%JSB	0�X�U���η��?FT�)�A�Σ/ �{?>x&�),;��琾�|Ĕ�o��E��.�03���g�E0�Aba�<a�e�:�7k�۳��]�p��緳��N��/,AQ�ޞ��i��]��ӎ����cn`1#���U��55�0� ��s�����q�v�l�o���k� �|�%j�S����`�b��!�DѸ��U/k�<�w�Z`eE9ӣV�JT�w{�2�7[�M��+l���L`�!��f��✋�w6�P���B��=z��]�j�V ��z�B"L$�YB��F��כ�>�>�/�������}7�6j2��F�ݛ�Ǡ�Z�L��2U��S��"�,������< �"�ϕ>_^���P�	茢EZ�!Kqi�=6uַ���A%�E��e&�ͷ��m9�<�H�Քls�vo=�B�$�.�\u�0
|��!D�ȃ���$՝�$��ok;�::i�MO�JR��Z���Ύ�3z����)wRS^�F�R��<0K��k͌9w6av%m�+y�Z���)[W��=�Եsm�*�)Jv:�W5�!&�^������"�0�He;�ud��m��eO�A %����)(���
bxu�DtS�]L7��?�����٭�emKљ1	$�N�g�Ky�_k�լ��30�R�rg��^⩛�{�.2�P��2YLV\b�\�m��=�l3�. �~���ȷ�zC#	�WM�~�"�~mpxOW�綣����)��3���;Qy>�v���t�������U<����W���
ݶ2�B�Q����C�&i��s���E�ٺ	L%<�g
պ��s^�}�.�wB]�d�ȗ[���]7d�EК���{6g;��KV�l��3�" ��f+,o_fk�"��3�5<�l*I�xD�����vq`�2����Y|	]ۡ;˵h�Or7�2��ִ�k�h�A�׼�I=�r��5L2��E��Aw���jޜ��6���-nJV%�|={r�sSi��O������1�}��?v�����)�o��I�w=�a�M�����*䗳�Un�ݷ}�eꄸp7�~�����S���޽�j���p;\��r<����+Ny���N�v��y���s�� *3�X�O�M4�nW��4N���}k�����;}|&�HBr~�Ia8V6�k����Px�N����#Js5<GF��2.��x_+��m����n]��t}���-���~d޷�M_چ������i���슋��v
&����"(c�Z����M�����	O����\\��I �$G顷Ir"V�d�e���\��+[�^����۠��s�Q�4|�7!i�j�2Qmc*&GsZ���ur�]�C|�k���it��\̕�Dw	�Yz!��{՞9���٩v��v�c�j�
v�A=���z3�nB8.Ȗ�ڱ�����;7N�.VὩ�`vWQ��t�`.�lu���r�g]�-��{m�	�;�=i.6 ��s�r���>Ccvh�5LwZ��;[���h���pݝ�3�[�k���^=l�u��Ľ����3���&:��2��:��p�R�܎�6vǞ�2�Q���Q7gx�RZ�ݍ�e�K�s�1`7��s��z�V�T�˙M)ڞ��%ϸ:�*��v`9xCL	vф�N�mc�똫�}o\�9r�;cZr`����ܼ�Ϋ�n����vLQ�c�۞��;��IxI�%�4ܽ�;E�v����V��c���x�b�7'��a����o����>u�I�ND��!��u�����[uq��mZ[n;�
�+6�<p����k%l�3�\7v.�7c7��  7i4  (PV�vir+�������o�>\>^��͠sJ�s˞9C\���n�қ�4�"0��*ې���+s�n�Z�H���4�\� ���m��!�=��Z�c�j�P&�s�۶�LL����U!ӜX4�K��߻��~�[�}Φ�r�rK�<G�57QP"ǨGc���;���i�cX�����2J�Dr�#���o�����ε���A1���=�V���鹉&���vVkj)ϵd���C�i�X�!��v���ڄ�m�׻�{X�>F�j8��{�?:���gvܒ�������8��2z~�w��N��8׷�k�:C&��Ւ�I���!L��'�6�͘��ب����|8C�y_c�E9�4DX�6n_���Fh�y)�q]�D�o7��<�O���ę�i�S�b&B�'u߾��u=N�B{��t�|�J�Ʊ��.�^�A�f��5� �c�x�s{_?���ArM��8�E��ּ�vu<��2JL���;�{���5<켸������z�7nV��}��������&���06�v�;bc���-3S]�z҆�uO�5U�gJ]*��Z�13?Gi�������O�1��	w��Vd5y}�>�w��|�}�[��n1�Lk��#����3SK�5�h� \�#>
{�ϯ���������^:�ٶn7.�%�˻�߄\bq�j�N}����޳~!����{��<�R�bb�8'��6r����Aǂ]f��  )���r��d��1-�#�絫�$�[��w�>k��ơ���>۬֝�����#��:���"+����f�����ґ8�y��A�]t(\g��ʷ���X�2O����?k�w\�߽�{�o;����|�l�~�8�͕��F�u��]��n���=o[�>gw�{Gއ����ZA2JĎ2�`�s�ס��P�sy�}�{�m�!�r�3���i0K�v�21�d7��;��ɭ}���Ƽ���q�b^2&%�q����g;�}�a�At�>�a�Ss��C�A����;�/�#qkw��[��DD��!y���V4���#�o'u�'_!�,�n�W��@sG>�=�}?8,�g�/N��y�烬vn79u�6�݁b6�G�e���h6t3�.1��u�)ǧ]��2��YuEk�9�4=q�k�p�mG^�b�6���w~�ګ)t�d��V��ʨU���y����'���\��ϻ���{}�؎�!�f\B�{vr�4h�LO��so5�!����guܧU�����5S��w��y�z�/R6�n�w�9������E�S�����t���ݕvn5`��%��}��y�i��g9�w��i�LGp2�9��}��&#� ��М�'�8��z�ww�����Xո����w�Cz?!~���1���ϡ���w�T�e�O��M<_�����嗎���K�/��g�c�3�:�d�o�� � ���@�6�H�DrƦCn�ng{3��}�6�57��5�}�oms���X�}�s�z�S�h�� n�v�����BO����ʮsKs���MO�" [�O���uτ�;a�zK/:�Z�\�{-���A�&&����w�o����W�Dܕ�j1.���>�ώ��0 �Y��\�`�BC/�t�O��ֱ-1�G����{]��77w&��]�r�U���iL6e=�8����>�{ﱯ�؎�Ƴ �˒��`�C��"m����u�>���9w�X����V6��X�N;u�4�o�u�9��p��!0 )�5k�pPG�6�/0�y��7J�l�zc&$B�1=�����P�G_6&s�y0t�5��$O�d��clM���]z�E�p(z�	N5�z�}�!%1!	g��];�ޘ���
����c1��� ��9�|��������fPb:	���q�l��&4�ۛBb&�y2�F\g1X��8����t���1����uq �B8��~M�u��w�~ٿO|���w[���C}���?��s7I��s�ܛ��ȯ���ݵ���n�w�����}�i'uw�.��q�6��1�kf��L(�=b-�7{Pc�=C�r�<G�z�\B$!�S=[q���{�9��	���cX�.w�/I��ռE�?g����O=C���ѷMbX��q����]-�;ʉ���g;�������/K�{ ��S����I�4�x~9������OU�l��:c�����^�����>�N0�㦌��h]�v^��:��ڎ2�Nݻud '�r�3o^�����r������8���ď^[cl7-���<����[r��� l���箺�+%�nF��3�F������ǝ����9�?|���Ͽ{�<C|���&�&ڙ� !��g1�ȡb#A�z�og9��1�a���v{�Y�˔�/��s�;u�@=C�! !"���_!�e?52q�s�s����L��76i8�5�"��Aƻ�8�Gn��}��9�s�"(AzT�T띞D������Xkۉ�*�_9�<��B*b�����"�xh�"`X�$BB��� ;����:'U������QEBn�;.d�6?z6��p����{���p�y�P� ��^m#�6�1!����J��5��>b"b�$!�"���jG�D]ς���:�s���,|�J�|�����>c<��}��oky=C��!!��2�g��U���zs����Gw}��N$q�X��Ϲ���Y�B���4�kM�B!!�v\X�=�:��+��y��!���h����!!�<#�A7���g�����5����\�!�{}��y������ɇm���'L�!��1gf]f���f�����^G4,euҾW�Z����1���j/�B���f���v��e+yd���@{��b�4�mc�ohEt��a>���}�׀�m<t3���P��sp[�7��97�}�t�u6���/�1�!Oj�����C��r^�4)�O��7��=�j>�Ȼ;Þ79���ra�4�)��8v��ںg�����w���`,��y/5�W��^��A���~�&q]��iCy��w�֋���]@�5�~x�Y��|�,/���}uL8�(Fh���>�O�ě�>���Zv�bytVT��a���po�5^B��E{r�B0Y
��Oֶ~2v�:�n��X��q�!ƭ[I�5*�c��RE�2U"8�<��apjnT�2Q�h[ض�Q�`�C��S *���5R�m%*-e���]�Od3.�턴dP[�L�	��m�RлdbA��-I#̘�kwUԌ�Y- �KV�,���I��"F1��܌������/���{��6o�Av�6�5��5�{��m 툎%�����޳I���^ֲ6c��"d%cX�����U���r������Ȏڛ�q�����z�r������݇�wuF5���Hy����k��پ��}�"�mZy7	X�qlNK�]V�5������}f��yR�߾�N	�q�K��+��=ɼ��{�c^~bm ��&L�t��91#�Lm�)�s�C�-u�K�+�\J@��J�-k7X�����ܰS]���<�k�[�E�"d#��~zC��k��s�����a�J�DkP�1�w���������EX^�Y9�G6_��IdQ�0i�h���J�v��cX{��]�q�cYd5߯�+�=�*�ُ����b!C���B�!�  c
9gt������5+	�����Z�N!��C�4���y����V��<��&5�_�ѐ�w��o�w�by��C�D�z��
e�7��,�̱��vN���螇�+?���6��"�^�q��J{r�v��AN����䓳�xz�OA[����]�Ǔ�����<q8{'�����K�N�i�k���z骪���_����I�\�N��o89�Z�wߟȸ��G�1�Mw��}Þ!g��f�X #Ã?0F8��s�x�jJus��g���>Dz�� �v}�,H�=B
|����v�h�kmF5ִ���bw��#[M��K��=���k�r�w�7[}H�%��!�>��#�bJ�bc��.|� !����������4�y�N�����="#��F��U�ڄ�:�gdt�C�+ƭ�r����k_nn�ɛ����3ތ�_p�I�h�SV�p7����E���^���~��x|�M?1)�3 �(������r��z��Z����1�=b;����$7׷�8��k�Ua�oz%E��X�!5�c���c����߽񶺞5	�㣎�~�?>�
��]��k�^i��˗&f|[Q��&52�|޳;�{�cY��L��n���j�&5�DZ��(zrcWq���pb�B��i5����y ��zNaa�!��レ �?PI�7���/��.��g���������os���������bbD�����;M$���';�޳�w��!���vB�1LLH��8���Ș�z�y�N'�H�s!J�'���~���q〶��td4v��cZv��ch������}�G�}5ry0G�\m1"bG&��l��ϬD��4�_;A�p�!��}�۲#�!bbk���7��5����/�����k_sY=>��H�Ӯ1�K��8޼��#�6e\�'6�}�n���v0�}���o�/�������M�gd�����"z2J�&!�|�u��RgW=��� D ��>�
��g{t�wWf�WJC�����N$q���ﯺ����K33�M���L�qlM�m����g��}�p�y�Du�y������d�K������5�w^C���qkoΐ�llLB&-o���'�<w�*����<F�J���ݗ�c	��:��<�=��S�<TŐ��O,eM�]�$�}�_vV���2f��� )��(�;�~����#�$�"s�׳u��v��Cι��Cv3q��v�8��L�{OL�M��B�������6��.Ɠ�Z6y�d�1�]nL���/h��MUU�������9��.��ѹ�^z��ҽ�����7��g�D�w4�����LI��BĈ#0웟X��^�l���pb�ޡ�Z�֡(m5�[�X���OO�������MJ���D�B_c�}�Ѣ���#�.R��wA�p���SE�j:k.V$�G;v�I�w�Ϲ�3{���B3���B�(HP��"3V��ϖu�_��������xy	g[��D]b!)��!T���~>~�#=�=v����h^>�e:�=�V*/�}�1=�>�ۚY���C�s[k�^�1�V��X�9	|כ�ѫ��apb�B3��x+�UCi�0o�{��[]O'3&Os�<bm ��b�������Mg���"�HC�=CiVJ�%@0$���K$���v����}��#��S�t��a9��Ǩ�L��>B!"s	�����3�����M$q����h��.�#�#���b),���=!o��q�nV֨�G���ɰnD�!�u�_xml���=b-�cYp�=�ki�p�����ϸ{s[0����j$A�O�y<����]F���w� b"j�������~�V���#���cd�2��"2#DB*bb�.icߝ��d�O�&��յi�9xf�9�mq9Nw��f5ֽ�D��Uı�Px�!O��<ꞌ��d�Ǽ��cDH�H8����8k��>kIi�C!;�nMf�:�Ǹye,۶jw,l�O]��k�(ើ����<g��]�9������7��[|�Ď!�n/������P�=7�f'��7��%F?�����˟���L�qr̼c�E�S��1q������}�H�z�G5�y�8��D�Aq����Dh���ʒ��]Pc�=710�RP��X��$!�SE���f����<G�P"�׊Ǭ{B<�L�}߽�^�ԉɗ��t��q�]C!���o�#oI��n�1���<�ѵ��\<��#{O_v� ,��U��#�Z��RVW����YaO5*;
�3�����k������`�!}%n��^ {o.ٽ���l�򧣧���vv����v��,�wkΕ+�N7�H� ݄��֏$m�]과�³����M�����<r�w�F�Wx�a���;��.t������/��7q�t��A{��tY#�N���{=�s����O8�W��q������{wM���ߣ0��$���k=���]ɒ_z�7#��,���y�Ƕ����R�OL��Nc�|��z���ۻ�p�oz\��wERw-~��Ѿ��'�X|0<�>����|�ѳ�����-[���u��ɋ�Q�st��rL>�'�}�j��Ai^�-�E�
�B�w;vZ���Ȉ���H�%6�rKC�EU�DESR.�Q����J�Ъ)�Eii�ik�*&�d"��T��K���H�@�B(鑂��
"����8�TiEE@TEQ� �9wY����iZ�jR�"ҒJDTd6�9||��:8�� ^�.��hQD�G��g���ַ;�w'�^��=k<s�k2�]Y+����[gU�q�m�d��z���)�d���<�y��5[��7��ĝ����=<ku%����;f�p�3�ܙ:����N�VخN�,���[gdx���<�]�����Rk�����B�r�CQ��6�=n.�f�.��h�@wn!���ݣFr�:ݰu%�.�n�xM����Cwk�.z燱�'��ٷj;n�+ӹ�:ݬ��(]��ɸϞ�l����ǲ]N;c�l�|:�b��D���i������:^0q����[5�n�����t�[����k�.Nxm��k�<x��-�i�vWrvmΡ����p�qvU`\���ݞG��b�n2n��nUR��1�q�/<C�QM�74��S���[$�df�W3dˋ� m&� B�M#w����z����s��>uNq�ѳg�=����6�C u!�Z��<�j�ݵu�m��\I�n�N��]����v�w2v�rs�-�z ��B񮚪����o���M�Cq�֗��������z/� �$�ci������;�5�k��E��"i�KCI��N�Z�p�lE�{=����i<�%��ְX�"E!��)�r�E����&�w��Ƚb;��cV����M��:b9"}�'3�[1N|Ĉ��vn$FL�d��<D �[�`h"����5�0 S�0Fg���m��(H���F��z��ҽ���~�}��y����M�cj����zG�!�<�D�(s���m��NR�������ڍ��Z����5on���0c�De������{�����i���/Iu���jd�lDq���ǟo����k�4վG!B*ѡ`�""�O�����'/u�B#CNgׯ�c�G��qkn�w���$BŇ�3�Ea�L\�!�#.�6�c�i�]doa�\����K�׭c�cmcgw�}������KC��S���X����X����'~�w|�{�f�"��i#���I�<j��b>@�BCs3��?*��ryF�_GOf����!toT���]ۆ�tPw���_����a���[KL����{��o#\� ��ٯw]��Þ	]C}��յms�2�c&���}�����s�'�{�����S��C�&&�6��=�>��$Ri��D�S�D�|����Y��mE�W`�C��|�BF�Yq#E�Oks�>k�<n��M�� ��%�I�S
fg�k���&�w���{��y y�&%�=�4q6���r����s�QN`@c�b��Ӈ1��GeR�6=s��/��nL�E��L1��ϵ�x}����J��O��TOo�k���>�J���Ʒ����o��u��>JV\�jع;V��1��U�����}��V&��]�_{�f�&��#p��1��q�z�m���u��}�a�J�Sp3�����ZH�5�[�#�_>�9���s[����Az�6�5���}��e�0#F1y�NSz�1�G�,�m���>h��ag3}�_�Nޫo}�a�J�i�)��<�u�s��ߵ ������7q��QDy�`t�y�{�>����N����ջ8��g�
�s=��<�^1Wn���\Q�d������sm��Nɮ5�{v-��1M=r'nZ��c[��.N�ѷ�����f�ܼM��.��Ęظ�f^1���#�G0�[���F�鼂�,D�"(BC�%j�DR�!���o���H�P�>���v��[C��!�o�7������}���X�C.V5�r�Z�k5��k|�y�a���'��>�q�iKq��H�g:�ngj�dL�{��okV<��[�q�﹭�����;ܞ�D��Z���v��-I�;����v�<��[��]��[�ov+n�����>�&<��hܝ�ޑ�#�td.�(v�#��&z������Xra�2��~�|��?g������~|�6�<��eD�'!+�bX�*V#�r���k�����G�M5���Yp�̟[C�V�}����0C=W�N5q�6g�<�BC<5��@��]n6�0�D��!n���|��Ȝ�ԁ��ۘv%���P�1��4F�g�L[�++q���Ϸow�:Ԯ6�11�B�������s��u���h��ֶ�z�u+P�B<��nt�����:���2�ʱ�t)�/f�a�{v�'����F���o�~���G��#�LH�!��7�|j\�X�S�Zk+9����o[S�}À�5�bb&J�Z�Z1&g2��{�9�W���DƱ5��u�l�c.�@����z�����}�������� �}[���0�yB�D��H��%cM�����L�{yɛ�~���G�h��/ܽgy������q����O��f�����������ߏ����k�c�X�o��u��9�b$D�カa�prp±g�3�yA�����(Q596:�J�����|F��$�jd"a2�Hw��3��?~����	��!�/5�_^s��2�[27�Nډ���w��]����ݫK���6+�`8����C�Aml���5\j�0�^��}��R&��R̄LH8��2�bO�z���x���]��������G���+�����y�˴뱻�s p����U�]�NJ�1�Ʊɲ�8���Ϸ�z�x�=H&�������x��<d�Ӗ���jF۾�vnЎ����{PB��=����i觞"�e���hd��Y�j�ֱ�x�3�Ɯ��k�%��޵�]��9�؍m�7a�c�՝"\��չ�Ӻ���\��=����������2.mp\�tm��،��s���7}�!� �\e�Wo;��VN�����8��2�&'9�ߵ�=�zֶ�vMtB�7+m��	��K�����c�����y"�Y�y/8uB'�C!7���5߻���4��o����8�2�{��1>Lϯ����!��B�O������g%O�<�=g9�cp�v���o~0O�!��Ϸ�w�����提�[�"�	7g�UW�0fBS��^ab��/I��F�H��{��~^��(�k��u5%i'|��s^�����_0M�����	���� �ޞ��]����{�ޕ֡�DƱ,q����bA؈@���]���>b ��w#}~#�&$B��	�H���z�f����]�5�B8�q���L�c�K.A�_7q�ś�:��w��w�}�{X�!LM��{�#D^G�~4<DF���LM}0�[jݱ������h砾H&��~����C,��S!$�!��}�]��oꤶ�ZjR�x5N@�������w/(3������Hv��z�N^���p8g�g��/�����|��eO����t�=9�G�=�2ч��!�cv��;|�>.�8��LA7q;|��ˢ���w,RsX����y����^'�4���HhwPޙ��4u�&�'�����?j�N�7<�s����3~�\Ycs4(﷍��Oq'���~Y�C�ؓ>�F�a;����>���[�(�$�Y����
<���/{б#	!Ԓ��<��-����|�������ׯ��L�C-v;�sP�N��OP�0gSs���9a޼��xG䇛|wQd�9g:�Fv��{Q�ޭ�N4�+[�ATUE>cN�F�`��/��DJij�!KZ� �DZ���PU4RT]C�"L�Diw �n�P�;��`�$C0�UF��)�J���b<��)� SmQN5��J-
J��%DX��"�B���� ����o�y�|u��^"��C�Aƣ�bu�t�R���%s��s^�����/�7��6ki�1�bbGd{���<���{��G=�D�X�=��|�茶��"s�y�����@�J���I���ɈC�������om{_|�0ձ���Ʋ�4�D�ۊ�E�ۼY[��h�4z�B���o�=��P�O��C���*���w!�BnV5�^C/��D�[KM�V'��k)����4y�7�������Z��d0j��!FW���5FC�fAH���vo;�se�/>��w�Ϛ��M�&5�gs�/�3*��w����q��P������y�=�q�	BQ��n��Pjp���C�<�A#���\H��VUs�V"0ya9߾�Y��Y11#�Ʊ7�{�cÑ��k����cG��!S��j��h믚��~`�8�����������$@����TH�� �S>C�A��y����공Տ1�DP�zBϦ'e^���@���2$��_��U_��o�]����������;ܿ��?�=b��F��:E͜���ݫ���ڜ�E�Pt�͹佺�����^ %����U��L�n�㮃ԓ'd�[��SA��6�k,�^r�IW�瞺Ŷ;sj3�an�i�m2�Rw�М���'��3��=�M3��X'R&��Xո�2��Ľj��y�l砾H�H8�n{4��ȑ9%c� �C�E�I���FU�v�@*��c�c_}�{H#�[k>���;���O�n�K-4ԭB8�6#���>��U�:������zW�#[�q�d>{�����u!���w\��i�f���{�mC�1�L5��5������˾�BS�5�8�M�]���8�Q7��Nh�62���9{}w�݋��k4�S���Ͻ�,zva��ϯ�q<���%&{ީ{wi��Zm�X�!o�ks|�s�w�h�^H�k��LNa�^�\`�C�+y�5�}��||�?4��yZlDt�Ď!�c�9�f����,�]ל�0C=b�<�euZS��"}qr�$|���D#���"<`�ecV1�k����h�Y���Zr�&H.5�9o������a����0y���!��½�� ���a���w��`o�3ބ�2�"��ut�+�Gn�Aw�������9�����т(D������q���-����\h����«I)!<�o]�ω�GՆ|�M�̈�Fg�LI	%%A
T�f�X �ܷ���	 ssW+A$��>%)ի���"�Q<�E�	�U�r�a�u�ݼx�b�Ϭ]�v�o[�9��b�b�f��J��ø�����Pq\n�>�~��k�Lgz]{�*����_��Q/h�Z��>}9�x���m�İ�����>#�w^S�t�s�9=�2O1�2��nM
���{�\DX�a�u�U0D"�[���E&K�ԍ������:q�+DY�I �e�*w�x��dx�7��5ɣp�:��9Tt�;_�)�.i���iZ;;;�;�f�37�����.٢�ܗ�u�;a��V�����c�,y���Q����v��`�v�lu�p�[=�K�x0��oX��݌���jΔ��z�ܪ e�x}wu�0e�e��mH�>�^IL$�-�$E� �v���x�Z&�G��$�U(�>$���ws��:�V�fLAܹwU��/��$�
�"��;[�z�8}#"�*E� �<L�;��e�]���`D�O����M��חP&����n�JQJ�iv��V�{�M�>��L�&�OB}�IH�ܳߗx�d�붿u��'�v"$��UC����uK�������-��ٓD�q���{��Ξ"I7���H��`�W=������
v.�FI� ��캈����n���$�q�����]�m���s�]��bA!#"�L������A��4<A �u��赴��s��W�;,�{F�0N��'1{mn4v(j{U)<#*/s0�U�f����p,DDn�����}�(�0��Q��������o�?d�k��)�D�"�yL�G6�n��({�_���}?g��O�#g����<�Q�L"����"(��u�:q�!�>"5:�=����/+{][�3���ȓ5����d�wM��B(�����gg�oo��+E�wO(�����(�_q=3˱?L�!�-TB�27� �>�epd�#ǣ�ٞ�W=�_}�׸�6�}~߻|-nL��f[t��IL� )2���&��ufs�zw���P�2`��9=X*r���yΜ1�7�.͡DX�$���IF�M�Vo:x�'�d�9W{ո�8�:d�,H�I�9[��0+�����P ���ܰ�-��cÞ��({�ݗ��2�溸���Խ{�\4���&��F�.ӽPk{zS��\�w�;|�x�gwyxzU�5�s�8<>#F��y�}׊���ꔞ~����AC��l���G{{�}����羫rj�E��糷��~�uI7JѸ`7[Hg�t̛Ow��8��k�w�����)�7ړ������,z���y�s8L��gX'O�� ���׌��OL�H�>�9�A�
+�����<2p�`�q�v��R��o,���G޻�������;��ܴwqFv�兡�����y�Ɍ{�bþ �\�vV���՜3�^�Q�x�O�B���&�&���$�z��c̽��w��w�5g4����Z�T�J\��� ��R���*
��@U���ͥ֒��h)J\�--"�vO�˂(����e"�*-�ZW!�E�4��UR-#T"�6�Q�rࡶ5J;�ڍZI��*	�����D�Z���"����Vp�!�N(3&��	��J
�E�<�i�(ER��+�E�
S�Qr	�򿗹~�nfHI��خv�T��Ι��鍊�pe۶c��r�׍�6`xǰ7��O6�Y�W�]5mn��j[�ה:`���s���8�+�8
A�ö���ڭt�۵�����ϐ6���1Ӱ�	�:�=v�U'Tz)�4��6u�8�k�`�״q�u���{]�à8���Bn��W���7h.3��n��Z嗨6�f�ų��'cgS��׃:f�Z1���v��1)����+�m�� �x�s�k�z��3�ʮ껪�f`�s��.�NW���9�ݹ��k7D�񞡗�w9K���	Ę0OK�7[$׃��v�cZ�e�	z�!�sq�y1�q�����N��j����.ǳ㹯���;Tb�v�{f�qv�t9γ�;{9`��W��=I۲d�gF�����7lv��X�U�����D���V@ �@   Y�+b������_�s��[��ۓ[<s*Rz�'X��)��w�����t��28�gT�InxcV�g�煛�=���J771-�v�ٰ�/k��u��F�3UU\������dN��F[W`�J�����G����v;�u�J|L�\�M[�i�B�ͬ�x��+3�̒ ��^tע^�{m��FI.��4�-�o]c2�8�0Ag�>�ݬ�x\P�s$��uA���"A$"d���E��<`6[e��Tq��޽����H[y��RAm_h�D�J6�[ӝsc&��	Aq��c���I<i?ވ����ϭ���y��\@�$��	᫄���n�*�	�[X���Fa�z��s��qw1`�d�JM�ٵ����v���ۅ�:s��	�
!2l䒉I J[r#���W�ہ[y"«$ɥ@�������W7y�5�1n���n�Pd�26�w��fx��6r�f�Er��=9xFC��~�{��u�) �it�̏ Oo<ڼnڎ�{����I�Xg�=rj������m�;�B��~��Ԇm��Js�]��bpa#5<I��so�Ӊ����c�s4�jO�P�]��f�e�V�=�8d�5ǳL��[o�L��^�0A�N�_s�!�����1�ӵ��Y�"P�U`/��w��.����g�w�����[�{�h�$������o�_w���Q;����}�L���rny�LQ1$�*kF� �*�y��W@��"�$�R�"���s��!d:��p�M�sc^u�U�_7n�$A�����$�U�s9��"T�A�%���ܳ��]8�$D{c6�Фr���DMnH�RR���I�|I�3�{�w�_�����4jSq��i^��>۷C�c��p�����]�m�[��<��:�
�=&�8�M�z3�@�zc'%�pX��sӞnI�,��ݦ���7~~�?���M� �P�(���#��q��v��R-D;r���j�q�~�s:�fr}���S�bw�]�:��&FQ��DU��,���L�
#� ���[.��:�$�W7�ݿp��4�F�k��߯���"xū�y�R�������w��8�&wS�KΥI
�P�)k�y�p4ȚN]���&��"#��Dp��~�cU&�Nlv�΂ ���E�vv�7o�,����Ї��ެ7O��ᐘj#2p�0k%<2�_�l�^��Q�bp���_.��&zQ��)��jRR�܈�Di��cv�"d�b�$���A̟P��\r�s�~� �Q�]a�U��A=.a�d��j����.
v*�.c��3Yӽ:t�=����'���}E9�YmD`�k6���v�F(��Ɉ�DA�=��`5�ǫ�:�2�r���J��H�*BA	)))!),�3�3�^���佂0�$m��,,���nߴE�3V�A�I�4���i��\�ޙpL�u!C��Ǹ�)����PT���N��{���yjF�bc;T�\+�ɉ��s������2N�ؿF;�{{3�n4G�v�c�AL4V&�m��(�C�PB Ʉ���$���V�w��M&H�wRDM݈7���s�8�Gk'"�`�&G�*ȁ��;q�ǀ�'��=��T��uة�;~������>" ����o9�x�8�3Q!��Q�גM�3�zAX�=� �lC�հS�\�d�I�(�l��\���aPda  $ '4>��Wc�a��t���<�Żt�9���$E�t7nT���ͦ۔whp�D����wǶ������\c.�q���gn��{*��8�u��;)�y^��]����W�uݜ����D5$x�#�W�X#U�[U�珄 fYu軘B	��(zw���oU$���"$�]W{�ݸ�9j�=`��/�>�U��V�{���b[~
������ʗB��`D�$�A��Q�6�0��]PoY����� M�}_��K��x��7eA0PZ3����#1��?C�uu�g�^?i�,P�����<oj�m���$�[��p�
ق:����v���칰L�0Nx��1COf�^�n4{�;��ϫ����Ȟ4��5M��D�����"r�$�]�|���i���	��-�:��9����o�Raي��x�����Ck��ت�Yg���V�S�zC��0�"��٧��ٗ[#v<O'0d�{���r���x��r�����'aX1g��������aT��츇�z�+څݓ����i��`S�;��A���hn�-��;ޘ�����}=��~|��O[���d{��{^����w<}NIz�����h�:���/���YM�n��� ��z;Kw�غ|Js^�5GS�|݈i÷t"_�黍�����9sٮA��Y�8hp/��,�{�G���f�Ry���$`[�ޯ�Щu���xyܣ��/Ur^� ��ڽ8�tv��ܞ�ڧ9���5%�W���rHΜ�晇Ԟ����s��O�����$�����:��͹�N���$�R�TD����J&M�q!E9�� � �PHEHf10�I��m��P��))((6��)R6�!�QPCM	�J8�h]ȥ�V��
�D#T�B�(
��rT\���q'�B�bj�����	m��:��PR4�.�&�x�8SX
F����ZF�Ťi!s>�蟫s�;��I��*H#�*�u�x��7f߆� �'�ˬ��w_��>�ϯ���k�8L��۪Y=() ��JYq"(Dgu]��w����A�]dy[Vsm����wfj͝�N����O�ݺh�:��=�w�p�����XNu��4��%��R$v��Tg@s�Id������׽G��Y�(�%1��;�����Kr�j���n��U��o��A��x���2тO,����i�ܺ��o�i��T�$z�Dqs��Nd;(�{��	7W���xuB�{5�'�ӌ#����d�AwУ��m�n�p�2Ib���frب��W���Gw���e��>{㟄���fY.C0G8e
QE&�����:�h�[=�Q�x�n�2,t���q�]h�rn�z;\p�0oY0ƍfr�۷e�z�.�a��u��MUUp7����/����R������ԘH��4AU*;���<�;uH7�L�%��,;����պ��Nf#�R�%�q��{�ݾ&@<�gmQ�}��	\�Q�$񫘿ڼ[��q�L��׀A�G��!O��d�B@0@�*d d�*i��ŗ�s���L��"]�"5�d��5�I1]Zj�ʂ�݇��F����w�M��;�F������Q���8��Y"
�T�&qԙ��\�����J�$*W{ۍ��9�̒A�����T^ok9�������C���0���	2� B&kX&�v�<�S�)u�,�c�(���k�6�>D���jp`�'f����t�X����-,��p�ZB��eM�NTv�}�v��1=7h��{���}�ϸE �b�P�Y�k�.0�Qh�U�]���^u�:}F\�w����M�Y�E�:��:�B'/rI�4y�k���U&���fT����V.�l�������&�p�\��oV��0DpT"T��7���kڋ^�=����=�oq�z�-�7s���{��WaNȾ԰!��!�.�(���f�e�E ͱ5W\�F$��g�/�����f"�>����֞�^7B�Ւ{�fw����;��<����@�F��~ѣ�	0������7����(���ʸW0w�wm�i�:8�]ɂ<A�쇆+.<�X^�k����dNq�
�r/���A'%�%�d�ɹ�s��Q���H@!	��dz}kK㇎�f�n{��8�G*B�v�����<q$��Q	�σ`�s��\�]��1ն.o]
�'�E˭�p�Y"�Lp� 6Z��w\���.���������k~o�����Oq�u>��H�2��bµg���i��
��&O�ʣۯ���D��r�/(�$�Ǟ�gEU��6f(ADm�ڋ
����i�
���_ɫp�.�8��]��zt<���A
��gw=p��l\\-$�1Y6�Vu'�.�c)�Ë��5p�#}�	\�HX�P���3�w��[�"�P ��s�#�����]	���2kR4�u��]TXB�G�-;�3�'�,�ns/��݅��iJ��1&&P I�*bT�0��a��Y�[��}�StDP�$�6޸��n�Qy��_b6���&M�m[ʴ�gN�Q��ېw]�|�zV0�4#>��e$����M=�k~�&Liy
RD=V�n�/�����G� �l^͑+0�s�ј;��_����Â���{�%u�4Fh��9�������0�TĖb�7#��ݕ���f��8n+	 �9ڢ{0޽篂2L�>�XB,D�8�s�q��L�Oz���9г�^Wq�7��$�d�Ϧۮj�3�{TE__=��e���bI��"BS�R䞑�:�t��w����������-d� �p�d�d�Y�ar���m8�*�\va��&M�c!�:��7Y|"��u,E��G{��|�P�ٙ���Ze���{B�f?�ɏ��z?�� ��P�E_�c *:X=R 
������ G��	�2D�D��a����PJ1���1����l�	�� �
 `� �E��d�t��u�L4[`0����1�p�@�xg]�^XP�2�\w���@ *?�y[��{/N3���~�;C��t��#Geɐ�j!u��R��(�����l.��,�0`vy����;�2�wP���G�����F������Ԉ��]�T�z%&C������x0���?�`~�?L�?���������y����H *<�S��{��C�T�7�Jh*d�ϲ5!7t����2%ȟ���HS鮩�|�6V��OX<Ϝ�ox�~zٰF�+�C�y0 �̘za�:cC1��k�� 
����'�j��Y��aá��x0o!�@ϩ�q�����yv?�jx>� %�M��\�`���}����>��?p&SD߷凑�{���|��c��\��vd�A����3������/�� Ts�,�h��>�y?��T=��CcP����z`�zC
`7�o������������{8� �¾�߀|#���� Q��%����}C�~G����4"?x��>	�q�5�Q�4� G�C���B�� ~v���@5��C��}82�<��}���G`�="
H!����Nɭ�Tp����w����r�NN��BM�ňp��=l&���B!�������+��a ��=�����=�{� TmB�!�!X=���a���?�<z�#����{�MO_�=����4/C���>/^�~i����'���o��5��` G�z���=/@�1�����p�� ����|������� �=���z�}�O����w߿Bo�n�:$~^�5& �/��<��������s�N�?�}�����&���z���[  ����	�d�����hX���'}ۆ�!����O|� �`��=�T�9�v�p2 
���+�t~�h�����G���?Q��DQ�����C��d��������xd3��v�}�i�e<��������{�w�.�p� 1�[