BZh91AY&SY���Na_�py����߰����  `ٞ� o��&�� � ��
�kM���             �g�ڒ�@  w���@����$B��}�)Z5=}���PV���{{�:�!ӭu�6��]9N�{�v,ks�����KYui���'t�M�v��z�S�Z���pv:�����V�A\c=wom�ʯm"�rw��ۻ�4q����j�>����ywh����W�EK����vn�9R���@ �/�0�)}�������[����s}۳���7�hr����W��w-����j�>�ӧE�iG����@
X3�����l�X������ңJ��-lp��u\�`n�Uן^��ϭ)l�l��N��M�Á�z ��U�֝�������n������a{ {׎�7�����ӾޏT{㜕)Tv�              @
�)ђ��	T� oR�R�`z�F ` OD�J0	���m ���S�*�S�� �FM4h  S� IT�4�`� � ��&U'�1L����ڛI��� �hS�hDM�"hЩ�S�F��驐�� � 2O��L�HR��~D�G>ӏ@E:U���EQM�� ��S>�O���Fa��E98E3y������x�?�����}	j)E�QDR�k�V YU}O��
)�(�2��0Bi*�O�S��@h?��K��G���w翩���EDl��?��3�:���H���j���ItN�cK��yQz�/]I}wڑ���m������RQ
f�W��{�%���~��wT�/T[yQ��'��.�T^���U/z�u�����m������RA�E���59-�_:i��N�*��r}�g˰x�N�������e]��;d�]��4i'C�g<=�ޏ^��nyз�XC`�GG�0�fPk�������M�#�h��B�9��[�����c��Z���W`ݕ{�VX�D׎o�b��ݍ���n�^�l��5S��v����UD�s�u=���A;DvOv�6W��Z�{���K}U<���H����$���e�>p��>l����vY��I4i�1|i|m|q|q|<�wC�����E���o��6u��LEp���Dz�=���}�&�ȱ|	�
4h%�<�*m�F���ʞZ��R�����|=������TQ�e=<��8o�Wvrh�>��cÏj-�O\�Z���wO1Mj$S-{Ɩi}5ǻ\�m�Ni\��Ⱦѩ���6�����I6�ԒZ��sϮ�&���ؖ���%���%�^��򫌾ܮ�5���wU��j��8�V䝸�e�/�N�1�-����K�Y���gi^ԙ�u����rD����4)�m'��smWYѿ5O��n����W�q��>÷�7Yh�x����v����s���Ib%V�h��Ix��g��j]����$1x�rO.��G�W�G<N�%�D�_���Vy+��9�Jt��Iʵ�ִ��Z���S^l!�>g���!�m����L��7�9�9�9�t����/$/����I��8{���۪t��H�_ܑ�LKd��-�{��#l�W�=bN�D�ey6ܧ�F1��\n��MI=��M������u���"N�8�����TԹs�-���!�i�P�5K|j�ϹU\��C���5UMR��R��U8:��M=�F1�U�ꅐ��r�x���l���[j�����$��R��W����xŶn'�X��ddj���n��m�Z��2IN.�^��X��c���wT,�UjM�{j���-7Uʯ�����~�I��v���n����\;�+ٸ���K�uB�Um�j���z0T�7��T��Sl���Sʭ�j��;�>� �a�<��&��}Ԇ���d�浦���:3�r�,%���I�K{+pNCn�a#&�V�T�</����Uzb����*U��$v/y"�cgKޏN�l��^���gNH�-��^HkF���#[�:;�w$~}�x�rGiF�rn�^�ܐ�v2rh~פ�GvoݓU�z66:YI'5U'�kR�)�l�d痞^E�_n�"�Z]Z�n���7]%n(�"������Θt�wK�n-�K��k�=f��p���D������&��\�G�x�3w'�Y�dnޙ��vX��&���k�.�"��8X�֙8V͔ɳrN�ޜ� ���:�y�q������Wd�U��MN�
���y$_
���2H�F�E|-7$����U�e�k�NG�Ea�;��#�H�}�I/�ЯAT�S$��H��G�Y#�ɾnM>��"��k�K�?��W��=�rE{�Z�}#�n�}�2r,���RE�$WW#�i�FI��]=�.��r/8�ȲH����+�H���qܑ^�E_H�[��d�Y%�Iͺ�.�#�W#�i�FI��]=�,��d�u&�����!4/7"��/EIi�\���y�rO!I[(�ISF�$Mk�nlO$Mi�7
��Z��u,�,vx�<<v,v]&ű=[���GCz�M���D�����ȶ>)�!m@�d�X��7Iu%��P�&���͞9��wශ�0$����P��'ó�C�N��M����H�P��g&��=�#GN�Wdg����nNm!>��"�r/�ɾ����]7؝�&���z/C���X��b�0����O.g����>[����s�v�F,[RiI�5�=�}�^/�yGyZ�ڵֱoГz_f/��y[�3��#t��u�}[W�W�W�5�]X;������{��ܚ�7&���������5k�z��v�v�|;��'�&�e�Z��_t[��H�th��r�Z�[<��0�����p�&����4f����]'6�#�2�U�c���d���Ͻ��vh�GE��N|���WC=�/8o~]t����[*��1�|�8}�n��"��^_+�ߕ��yw'9��M_<���q%kAT5R<:>쏇L����$�	�I��wN�����{��C9]u�RԖ�<�Қ'�3g�{z\�k��pǛ\ע�Q�}�^i����eԬ��>9��c��8<&�+�}Ϟ}:�ۗ�i9OυvK�XȐ�G��l�	6�y��6R����Fݵ"u+t�w���/.}��Z�^-NO$�裢��?G�
���s��QJ�W�H���v���E�誾� ��x(�Q�i�����ӭg:�8���{���g���u�'�}�k�iU�!���>����LTj��d�X�a�u��dB�*\J5�ؿ�����i�'ڪ$��S9A�e~��5��gzm�34��:��~�P2#�C�]�|�g�6���.1n/�<z� N����>�逛d �E�Fs伴�\�A��3��=Ps�1h4��D?���y�	!E�n�~y�Df�:*���aMU�L����4�֦�X���Ufr��"���w�gwS��"����pe$@��6d�	D!�D����X�������E��ˋ����C��θj���I�`C3^����#-L�E���������@�D��M~�ǧ���RL���
c+N���os��2��g�wΜ�6�<gI\�$��{"Y0��&A���,dE�7��x^(�t���f�Q��4��jy$	���X�޵K�-��^�M��a0V{	�(pT1��"�QQA[��_g�TH밾��K)���`�Igf������HYg����5�Pel�V�(��%X��C(pF��l��D���w�;��ɌJ1�<��6�!y1����.U"'	�B�
��Շ$���꩛�� ӒD��T����Y;9\�][���(�9�N��EAL(&��k�s5�����${�3�{�/WQ���m�vT��z0�{וш�7.^/�4�Ӵ���������&�˙�,��[wszr�LJv�鷊9�?���2�q���[�-�5��C�"��ӻ'��~�x��,v7I4�#Y9�h�.a�.b�̒߾ۋ�=�]�CN
�XWl=�{�R�S�Z�ǝ_xc��v���-����H���$�U:���/vzk�H�����T�/�F��U��{���~!lL��,����r6�5is�a��R�#2��N1�ټx����I�_'ҏsKC0,��o�X��}J���;�Ձ�<Ugw�4�I��l��*�	y$9�f�l1m�>˿�$Z�|��^�[��,R������CY��	�������8������~��s��֟nG%(6�M��f�ڟ�M��N#�����I{�c���J�����-0%�b���q�Hh��j���2�2��On�u��6�QYY�XN����/|�Oaݥґ��g��/kZ�N�m�d��zpE5v�+3���}׭�3:k�m�R�f#3R��[�h�k	���G`��q�a�>8Ot��}}��"��ʙQ�=~�mb0��x!�oL�Cԍ(�Ft�NzO��x�j���J;C��n]�_�m;������}�M�V�h>sW�,���Zh.�8��Z��oIV�L��$��ڞN����2��)�͖#	V�H�%�o�������'s�<\�c-�$/6l����U�%���
�ޠ�Ug���(�'���ȁ.	�i�5j�l�ŗ&�EwE�! �~�k�.�5�����!Q6�i��8��CWA(0���I���lè3���zw���z�/�X��_�-��'�'�O$�+H[n�ř��!Rk�ɋN�h#�C��ǹ��S�~I��,V��?D3�W�>z����/;�U{�f~�]�.�S|䮉 ��j������6���]̞YmF`����u�i2���E"q&���8^�ӈOMѻ'
pS9-���)��V��J��g�#������ށ���Z&L����2�o���f)��	��W�!FIĞʲf8�2cH��d�9�x'Q7�خ�b/
�R{���m��i��E�0���F1"yAǃ(u$�$����Ɯ���S�]6Q�KT��Z�Ӊz{#]@�v7q�uEac���;�!#s��2��c�a{bd�Ȫ72��n}����tw}��֢'���ՊU��0��{�:c-��t��q�ib�Оe�]�����W��iĎ��RJ:�̦t��A�o�����d��eX�\�� �Kh{���)��Æg"q,8'��Z�u��U�����������|��HZ%w�Պ���r:wu�� s�ꆫ��*7Z�vƴ�Υe>��'ԇN��A�7Ӌ�'��,j�0��O��]�$��e�	ɞj�X�ETm[��X�`}y��$ȭ�rw?w���&W����?j��(��= �i�j���h��_���߯r�:���U�CJ��)9�/^��UDt�K�����}�l���t3LP��1ڣM�gAE��\KN(t=�Q7��D�U�0���4̾3�Zǒ���,#&*�w2Qc# �Кe�Uƪ������Z�♛k�&�b��f�� �zĢ�آ�ʡ�p�Ȅȅ�g��;��O�׷v���bBHZ|�t�Q�3캮��C0�@K$��������3�vʜ���,�}�;N���6�Gj�*M#byVD%麊��	x���o\�|eZ:
9�Vve��L���>)��̘`�m�#�(XlIMbO��t�iw��9(�ukUj7Hi��s
�>�.��Yͽ;�5�)Z���SO��j�&������~J�t*R4��T!T&�|��=�C����v�?C=�<��uuηq�s�;����?/�(�4~�'Q����Y�}���޿&G����:�R��蜟h1������2�}>��c椉|\|֜�P����,�,6�mDR]�D��^2
��� BX��TBq�c&BaF�	d�^\c�y�lA��6��er��i�a�M&��ɂE���Mĸ,U�s%�vLQ�*ș-�Đ �H 8��W
�5���$�FTZM��%���fD�jѿXz��M��Qf��姌5�ejG�7�D�������	�R����0BF�M�0���8��ս�\8^VP��B�CłGm�"p��1@�*r	��a��C�da(DI�z�1.1$dƗyP�2���݀��8�j0D���FCl��<zx�c\#\'&T��##�b\���уI6
&0�m4������bChP<�N�	A��	e�B�f���W�AQ��,��Rq��%y��`����AL�!��-�e�՚hB
�D|m���B_LN�w(:�H�
8!�ni�S��:K1�K��!��d���0���!�i�xS��b��(5��_�E	�ۘU!4iQ.8d4߰Y��@��$J2�T��($R" �2(IN�X�G���KF�i�	i �)���	o�b{b�N���L��ZD���NrD	2>���&X(����0FB	�LS 	FL��ʈ�Q��o��
	H6p�e��>ŕ"�AkRrB�
�A.`����bk�'�NV��l����vkF&U@�@�QHdPz��d�Z	`aB<ѵ��xB �7E9q� ��\n6JDIm�Bm�-���=���Fl����C�����Gʄ �!||����π x'��O�䌜?H�w)��~��?������U���K���I���>��~'K,��,���"P����DDDDDADDDD� �����$(DDD�,�:"&�DDN��4"""tD�"""%��B"""xDDЈ���(DDDO�B"""xDJ,�����b"P����d8""lD�"""X�B$ ��x��Ǐ<5PjH�ֈ��
�SD�O��؈�<"'DDDN��8""lDDЈ���(DDDO�DDDD����� ������""""X�DDO�xD��"&�DM���8""lDDD����6""'DD؈��b""pDJ,K(DDЈ�$�����4"%����ADD�"""%־'��S��� (����
GPcR��""'��"hDDDD��B"""'�J8""lDDM����6""'DM���4"""tD�"""%�""""" ����B""'""pDDDD��B"""'�J<"P������DDD舚4"""tA�"&�H"""%��"tD؛: �"""&�DO�J�(P@�N\J�%��$$�2h�<<<<<<>��"""""�����""""%�DDDO�"""'DDЈ���B""'DM����8""hDDD�DDDKDDDDK�����""""" ��""" ������""""X�DDM����DDD舚4"""tA�"&�!e	B"""'����O��!>a�2��#J��b�B�"��- �@$0k1�;� �H�@%
�4��P�H���G"���]@d
ĭnMì�#�r5+N@���/���_�?p���0R��������
ϑ�}�����>�?�.�]��;g*��%G������Ϡ�c�x/G��>������b�~�r+B�x*�=�����ة��m6����^
�=��hW��6xQ��'��ޓI\�*??s��O��о�^�I��{�Uz.|�k��<���N~N$$J��dI��P�D��#D+
MI�M�KD��n)��14Y�Ej�!M9c�[!d��^d�♗f9_j�b���a�$)���5��	�E� H$܍B�l�ĔG$�F3bd�0�@�����#m�\mǪ1�"[jC���0B�d:�*�J6��Fd)�i�,2[aH�0[�؉"��&And�#Wq/2�k4d&K�I.A�-�!��s�-JpX�|�ĎH��
!14�PiPZ�E��CT�!܉��p�'
|����f�/ruQ+5�t+ea�e�H�{��r�ط!�.CL��-�,�P�ˬ��񼄊$!p[KLp�`��I�b�I|n�	��Ƭ�A��0NH�Ap�R��U�!'7m�E�M�RjճY�[��R��HƧ\p�$��v�0��,a�����5��mTF<(C��Θa�""" ���Æ|N�:a�`����"""p��}��:t�a�""" ���Æ ӧN�a��""""���8`}��j�ދ�{//�-��������NM���$�8�crm5�]���L�嘤���x�Y�B��*j�U�.踸��!d��L�d�T%�m� ����R[���ʪ��#Z4N��֭��N�����ԃ�"��uF���.#�%+�*>��֤�i�ޑ�5ؓ��wZ��;�]�YF����I%�����%�h�.Yu-�V�3Z�TG[F�0U[=�ԙ&h�{f]����;]���^7�[0DDDs.k|7�6�7�2�D�Z7�|�˕l�����65��1�Gj�+ޚl�<F��O���]��-��0��pnV�j���t�4��������٣��|��q�A$�57G�aڴެ�=�����{���������o29"cydЈ���(�}9^GU������v����6���0��Wޕ�w���FoRh�7Q� �(��р�{���pQiors����imZ���;�Ih��C��M��Q����	���ɩ/Fftű��_�$���!MW���h�P���ZKG��7��3)���p�O$�0}�q?(A�����v�I�?*��\�[�:�q<ǆ4��;F��H�0��G8ٷ�ݢ���B�%}w{G�wgm譍���6��yJk��*�"�M��!�d-0�52�[5��F�.�$DУ�V����2l��-�A^U[Er\� ��
9]Fp�A���7�1��-�0�fb�ap�� LD�.@Q�&"�|�! qHB)ٕ32btDDDH^\ӂ�!���c��D�ɍ�!2ĸ]�W05D&�cJg�%:	�p�Q{�=E��!�\�/3p��z��e�����s��+O0��p=CFW��u�0�ap����=s�m �~��a��8�� �0������;��(�Cz��$��{�5��ݗoEll|���=Ό"""):{4���|��Ƽ٦�I���;�o�k��=�����Ǧ�{�o���m�o��79ŔP�sH[�X�_�d6Q�h�b��ja�wvږ�B�n���~~FI��r�|横{�I4�o��5�+�ڎ��Od=�ћ<�Ell|��
�,�]��������1���\�qi]��*�3�-����>#�Yx�����߇�h�0�|M��N�|H�kD��ͫ���j!�9qGDڧ1kJ��x�뀉H�(���[�"-*]�H[,e�\'&�.W�4v��`�Ee��p��A�V�\��;���2ފ���,/wj�>�I_J����>p6W�N,��%�7 �"4���;GCZ�;4�:�p�h�fQ�����\��qi�"�2%���Yy���$Fj�_*�9gW8�=���9s��+Hr)ǈ��2�MIz26>K��Q+�p���NF�P����KQ��\���g�{f���l0���F`F�D$�$ko@ݬD�V"Ͱ���A	���P��j��L��%��吷:"""#x�4�f�i�ˢf�%2W��_�j�Q�>�NV�զ�kp�<�&N�����S��$�ή�|h�!���-��z��8[�:�μcD���;FQ3��.ѐiX���H�v�>��z��I$!����{�=����[%�:I
,����7½G7a�w�4]���m�(�te�������O{���w����B�i%v���H��J�G	q�q �8��a���#d���q��g5�6���В��Z;ú ��lg �d�fA��d,��@�`�at��Z| �C�}b�lC�Z>�>DO��VЂ|�ɂa ��aC1�7�,a�p�k�Ǝ�̇$�QA�(/%bPd����,�1��ξ<*f3><����<�3̳�c��4cY2L��C1�0͐c��=�a�x������L c�C!CC��FC!��;�Pϡ��f�ѐ3��%>d�4�ك6�7��
��0f��%�o}�T2~T�R�PS�E+X@ر�2 ��hf3�#d%����ЬLK�
bTOW!���|�l�2�3^H',��u��S�g��F�O*�F�'j�b�I�L��I��زT\E�`�^f[7�ts=պ�s(�@��0��:x�a�`X���b`|:tنa0�0�f��8a�a0��0�,��0�F�@���0�!����	��a�͖x��{p޽��=�3:f66>K�P�	B�!!A��>�
��rN:�)<&ݹ�N;s��C:+����� ���lKmw(��G>�B#Q;>,���]�X�@�"�L!>����++s��WF���|'���P�[D{�p�P��P�G3�������4|�c򧐐���k9��ya�:�e��{��};��0��#���'��>`���Q �h:;�zkF�f��6_xw�w���Щ�B�!�WBJ�p�bz@ ����l��B�CU���|7��/�.���T��5U�1��k�~� �zgYVޤ�)�C����O�$m:�;��;чs.�A�%6�����e���nތ��N�>K�G�R�ڝjP�l.�@Н��#cÊq��;I����w���l�͙���_,��o���1�S�Bs�F��O���!e4�H�ZR>3,�D6[$[)��CH�I�].+�e,��Iwve�c.�%�)n��"��Ww	Cx�	.��W�B�!IXGZX.��֪-Aa��g�!�HtP�m��0�B'�}|�� �r�?e�{&\����Ȯ4��)/18y��q$�'	&d����1�ﲨ������i/O7[�"�6`�"n�����W�n��	
"�z�ZZc�e>F��l�[dRb�P�ȹr�	kd�����"�"%�Mݷ&PC��{�¶&Q�Z�J���ģt;�sr,�l�ST�����û-Ι������NU	���%QB��u�1�OZ>�Tk������7i^&/)9�o2�t���]6Q��AZ��q�,hI����D�K�����}_~���{>J��!�+��ȋRM6J�>�ь�̠��CH%s�2�q!GSokI��m��Wvr�&A�P;�5Z:Iv���]`�p>$wt�����1:�zH+��+�>`�>m;� �^�"eu�Q��Ю���{g���3|����_�EQE�!$B����Xn�P���C�n;o ϔ�v����=|��$Pm-ː�{s���h�#}���O׉���IJ�H4�%�>��(v�&�!K�@>h�2�:>t��Ժ4c��(u���[�>����;�7�uTq�}�i<J�t�tݷİ.�"�sHn��J8�^��k����*t{G�6|fό��e�΢ܰ�F�!B� � ���Z���,/15�J�MМj�!�]��G>��joy����h�A@�<'Z0M%
|�R�|�!-QH��,øO$��Cw,<C�9xB\�R��YL�ҷ�ÚH|a[L�.CNI�A���NSBdz���n�\eYp���P�@�kq(iMAkF�����ٙ�.�坭ݓ��ˑ��Nj��� �j!u��2�P5�
�������(D�)��	�/���j#�'Hxx�&q4Ja� ��D&Afh��!B	��_dG����rS��*U(|�(��'�.]/n<J���z<i�.�&5����B1]����"��p�<b<��ɑ�ʛ:�bо\TF+�	���y��M'���uo��y�Ԗ�#�PLS�!��%Ҹ�ah�⪮�|�h�nͻ?gKΙ�b����C�f��g�!B�4<J��;;[�ʛlZ+���
�\M]gUl���jx��<s��={�M�d��1˳�iX�ᦃ.	�4-4�٥���{��G�K�M�.������^�od�)n������!�*���ZX(\8�@3SL7G{b�p�Nh�}1陖(�/��UVUj��	EQBH��|{�sU�=�_tF�G�N5��<:y�N�Nê����w�T�O��H�#�?x!����9�%-&r&� J�?F	����t��#�᳛GE8�5(������p�¼q�K8��t�i��V�V��'z9��̾���=����~�!B�!�U�}2�#к7���kd��&:�d����reݬJd�m���	�9�xԢ������2Q���Na�i0!R.�D�E����\Rpi������4zQDF��N�T1�>h����i9�a�f�u�r��kH�77���(�M�����Pѕ��0�o߈��vD�'�y�'��c6d̸mc,f3�o��i��ى�L[�Ft��>DChi*	�&}�F@���2���px�� :4cVl���*�X�hƬy0�\�!��(�2硼(��d��3���f3xCo�C1���֛�1�� ���su�����P�&��C�bTOͷ��=$�1���Al2���P�fQ�(�gJ2̣ &P`�a�A�`Ͱ XT�
��xd��O��ʳ D� � -iPP�E�MD������!�hJ�|��C�GW�U�%��X�O"rO�/�����>��X�{'c��gujiF�D�m�Z(�HQ	N�=�$�'u�0�T�▪b��C�� �mB���D��f1��H��rY��9e��2۫.ԉ6�2>?���r��1{��^�� ��2X\��x�
(\AF`0H$�Ba'B��=B*�sS�4$0;)�H8�����9se=:1p���c��YݝK�u��Z+([
lF�d��Z7��<�Re��;v᠖1_�Ģ��,T]
��"�̮�����K�H\Y�Q�Q��IJLn#A<"�B04Z����U�B+Hi0����0&T|nD�f �$��abQ�K�8PX�r�ۍ��	u�	�����$+�`�
g���^�=KS�7��,��e�Zr$�d��G���
�y��m�Np`�f$Fbb"�Jg��-K��۲ȅ%�YZ��q ���ƚ��J��j.4!�h�3	Kw$f9qR�k3+Đ�NYg�W�i�Cy�v��XIa�|=*�5��o{6a!�@M<~:~,�~,L0�0Æ·0�0<"A0�:p�0�0<"A0ç�Æa�P���� ���Hp�ɽ�͙�33��|���rɊXyx��BK,4X0�9�G��X絍�����f!@��k-p�d�	��f���M����ϋ6�dH.��b��1Ӝ �i�G�c]h�Kw�&�EHA���1�jZt��!B�G&�H��̘�%��Ʌ�ۃ�V	z�\%�<I���|u�j��)�N|L(z�
#�`qgeF�r�)D�4���Fwh�F�]�;ݧ�.��!B�<Xb)G�l�پ��SG)'#�сc�cϞ�����(�?&�h��_�̩|z BѥRR4��~�"��"�Y����l�t���fX�俷� Ue0�EAA��[F��0)m	��� t8�����ڮ�p�Bӧ��Ƒ�KL�Q���#�+`f���[��k�%~2��U�T�#c?I�J�Rf���p���Q��բ�j���+�Q(�si$U�Z�j��@×u��3܌=3�"�cL��8����&�L���ݛ����3,�|��2�&��6QE�!	D@�{��fo\D��}n!��4�ܔx��8��e/B�i�4r��(��Z��t�G�L���fYy�]��h5���j��߿k�>L�k<@k,����(�Z@�~�TY!�9Tw�ɥ��j��:��4H��i�yx�j�z���#0{����8�l֍h��o�=�33�Y|������كZ,��!BQ%�euU?IJ�r�8��%W�ӫ��M�8�2%�	�lբ��5��W�\��za�K��q8T��4�	a劂���� o����i�6i]�@��`U��	�+�ĭly�r��y����C�Q��5V��B��oȋ[GQ���kEh�f�gfY�{|;�;��Y�	���JD��G�""ё8�k(k�u4��G"Dp�陈U���H cE���I9f���3	$��@m��l4`:�VB�"�&ay��E�!B�%Y���Sm�F̀�ZaH��д�`�/.҈����<�P��m��JUJqz�m��!�ԓI��s���I�p� ��rUz�����[hY�c�n��� ����3�1�ڍk��_b�;��G2l���x��i��;DW+��O�\��oF�wGj�g�~�LG�aR}8�&QEQE�PkC��>��f��z�l�8@�e�����܁g��D#J�ԗ
gb�� ��:����u�I���~r���]m�;x8�^t�Oc��n�S���氒�5�YZ�DZ����A�u��P�-BlE���`�(� PJ���b4WiF" �\��Y,`ٽ�Q�2�Q<n��Zѣ�.�g��fY�_,�޷3sz�钷��?�!B���W��Dn���jt��H��8����ugHL�q��\C�4����̭ M	�1�˷/5����J�������(��4qmi�A D�sH���� M�77��5����g�+�4��l���rĸ[m67y,�����j���w��z�yB��KդP�i9e���Kp���M��� �J��u��!��8sF����̳0�Y��ޘ�$��k��!B���+Thd�X�PB=��T�M^W��"W�����ɟj�Q`��'	�:z�3#q��C_s~�)4u2��������A gI��5 �am�h!j���fb�]*k�F��j������5Q'���6��y�Dt�zӸ�O���}d��ƔR�B�E�"zx���V�.�7�}Z�B;��I�4{6^,�3��&N�a���r5/!v,�b��0)�TH%R@�Ӎ&'?Q(�b*O]p�q���NUL\qDq&�"�CӀIb4`�! ��q��BqF���ȁ��-;$Dh�!B�%�N����V��vE,�R�@hژD�(\��zKY�[��CP�S[��V�(F+%lP�F��eй��@f[m�+��(��R<��oK�{4��q�"��v�΅!��{ϻ�T���W������V��w�]�h�z��Q�`}�Z���#K�h�gw&������̳0�a�vI]�.En����K>!B�!Êה��mzlN�"V��2�_kZ6�J����M��yh4!i�Ω0�7�6Jz5��_���X���W�K=tr�v���"	.�w7wqd4b���љ�,<ָ�	�=��F{�=�R6������χ	�N瀨=OM��=��J
�H�73�e����m�2��4L�Hd0h3ҏ����j<cȈ<`�(��<`����"���+����a���f0�8a��эpx�� :0�$�Ġ͔�dK�&Q��s���2���o
$3(�h�2Ҍ�@�d�z��B�f���(��@�x��2	�;�`�@��
f�)�3L!���3(њ1��3�A~���g�=�1�d��dL���X=��F�0�KL 5�f�,���fYQ>~ )�)O��E4Ō��d�1�c(��<��=�g�R�Գ�Zp�c9�Ko2f3:A�B��7��/ ^�G�w'3�d�I�p2u	�d��#����W|u��x9'̃%O�q!į�X<s��9�w	���%Ԫ�@�Gy+��ƺ֐�P䁴7 q(�UU�h|�F����{�}�f�#	�5ç�Y��?"""'�H""aӇ0�0J�$8g�8a�a�hDDD�DN�8a�a�hDDD舔"YFC7�7F��̬ᙖf�:��>�ܐ��,��!B�@M���YTۈ��P�8�����k�m��Vq�s�.�ԣTn�U�u�U�f�z]�ċѦr����L�T�́�2��[e�d���m�8��EW���m:D-���H��6�J�m��-%XjWSFګ ��S�$��bi���Q��P���ʩ7F�sg���fa�êVN�F����B�!(��u'n�%݈Y&��D�!�7�#�Z�J�\�,����T���rA��$�F ��8(F"1�W��kh��s�t�0�1fB�!X���wkM���(s~�k��ƴ���z�<+����!��=�ж�<B�xa�᡹�L���*OL�5��9Rof���{|=�f`�~�Y��P+kʰ��`���UC`�q���i4��mX����|�ر���-�
n�x�s�x�\D,1����,�4a��!B�Mَ�f�[)o.�3X���*l�p g��5v��7F�P-j���Oχ�V"T��كl��y�GqB�%!}"z��D�5P+P��H����Et�J҅�P�]PZ�7E���5��ܶ\�m�ʑ5�����|۞���2z{��7h=�C@"�+Rn���{�ft��;���܁���q��L�u.s��L�7��܎�`��R��.q�Ha%����@3P#���Uj�%�шoG��!B���:�6�GQ嵦��o��"&&G����H���iiJ�ooU����#4�7DKYR]�r7l��#%رn����6˖�%�eؗ,mP�����Y`ڤ�b��-Dm��1eܕwuke��7w	jB,��i.1b�kF�ŋ�AJڱ,ee�
��+P#���
5�Z4l�J�kF�h�s2�-�I-�|�O@c�'X�	�ƝF��׹�Z]�P|�a�����0�u��׌���"�e�ȵ.��`XӔB<�7
��%k���7�Z�g�Pz�d�Q���:�%L�N�m�wfqs�32Mp����p�gK�3�Zzh���!BQ9(�'�=&_l�4:F55�B(~N�`oٴ�c�C����j)9�h<m?���	���&4�@��R�ldF����\}�&��P��T��XrI ��f�P	���&n�T��S*�y���a��߷q�Hel�V�J���Je���Q�0����L[Eu�Ö��K��f�{�ft��;��'�v7"���Ʉ8B�!J!����.&I)�X�%��"f�m��s?����� ���Z�G���1�Nv�D�U�i�Q�?�#LGi����m��&��\�7��6�W2��P�C�OVW
|=�ލYU1z��M�ӮN����<��*�Oh�R�k�Sl�,p��(�h�:�g�	�u���lv�䝓g/g��3:fa����:�F�M��n#F�F���[yvd��1��#����|{��c��7F�ښ)U���HebJ�qX!(����GƜ�ŎY���&O�B�!	D�ޝ�a�/0̵	"��
��#����Z�O�c�B/�ߵ,:�q+Tպ�B��l0����^.}D�4h��de1j�'��]'���%߅Dn��!��
(��"��GS��h�#Qh�E����Tȋ��[�$�4��z̘�"3&\�Y3cc�Ț5�3ݸF��ޒQ�eԜ��^���ff�.!dÜ֦b\�:�8B�!J#_}�/����|���ʢ-�r�7�w�%������7���\c"�ܴ5�S*o�h.�t=Ԑ�0�#�M">%bl��o��4Ȉ|M���W׮\�L�b��)�"�J���	��̶�Ϯ$�]j^���=|�;x����r��;��'4'�J�p<���P�qt"��v��Oh��x����/�!�ID��	�B�!(�G���r�}D+�<T[�X��J*��j'h٤v�C]�H�5�9�2�C����*}w�w��e�f*%AH#f%��)�h֑H�ε��)��""H<M��<w�'�$F�T5�Q9괬��/�Ѻ<�k�c.�T����n1�1�4�<,:�E�lr��)~F�W$��g�O���f&fw�Ժ��P%�QEQ��sYN�J�[J��;�Ȩ<�_෎%�b���z�FT�eb�)��ϩ���=�-�w���*޼��jΨZ���uh�iJ�ֽ!Ə.Ck��E�!�OH�0U�
ח
Z��e�gpzLg����"�Y�$0�.|pm�3lZf��<`��<`�";<��a,1�0�ha���X�1��,��1�c t��cV0į�HC(1(�$� ɔY>2|�F�&Q�40�7>��d5���t�f3�:ͼٌ23D-6�f0Δd2x����L�a�(�X@SL�0f�C1��3 $�1�Ό�e��o�!���� �gLѐ1(�	�a��(�o�a3m�� �0d����\:%��S�L?��E9��6{��l��}�:�ڎ�=a��h���Μ����z}$z��}��w�E�q���%��@G��#�ɨ`��H��SiG�$&[�r���S��k\�d�$����4`cMTl'$p��H��H�C* �
�U2K�QP�#��yJ��8�8�U1[��
�jr%1y�Yx&$K��+���1K�"h��ҭ�0�2�-D�RL6TnrW��у4��b����m�L��*�[Hk�����E�� ���[�UP�I���BdfB����Fq�FFqa�7l�`���S��}nr��I�X��r�.�a/;�nx!*b��spf�bi(dҘ�1���AB�m(����QH*�E����d&�Q���d�Ң�
Mp�O0d!�H�S��xYU��L��0��l�v�jWO ٪����Ԓ��AԤ�F��k�6,	s!#�RKc��i����E��J�.j�S6���m�ɬ�-,��rɆ+n.���.bDF@D18���|M�ArG J��sDf2۸�RI ���6db����b�V�5��d.=��R,I�X�p b�d<����?l��Y�L0�a��"P��3�8p�a�hDDD舔"'p��0�0Ј���(DN6aÆa�a��DD���"'��w�;��>�G�}���w��C衊5�
-�F�R�����!��P�6bH(��j1���$����[�yc#���2�`�&e�Y�K,��gB�!	D͸�n�eː�.U��dW$�	7_]���E��k<M�Q�����/$5Q �O����hze(M\#ȸZ��cG�0&�}m��Ц�:�4��Oh�S	�!��Q�i#_B���]�p���f\������H��"F�4E�h�
l����D��	m���Q޳��rw�6{8fe�xg{(N�!B�%ڕ�����;E�tsp�|�u�"]\��*�]�^ZU#�:Y����S&�[K�\��Z�x�A�i�6�q������q�	�Z8�A�+>�e_��!�#��)���FZ)����5��c4�J��2�څ
B�B7(zm�!�C5�Üi��@\"���;�$ܞΛ=�311�.�!�55�!�(��
(��h����0$����d+.v�h�:��=	G+�UJ���v�ׇu2�3� [�;���VAi1
# |F##�QM�4m�P�퐤;�o�%b\g�iE(G��CH�	y'����m��^�����4�q�4B�p򀋼�#��ζ�*WmF�,T��\�_�b!�sl�d��2�ᙖg0���:z���8h�B�!	S[[h�K�����t%LY
i�jW��nSZ���ZŐ܌�ڶX�J���2I[�#�ZT)���GebC~}ݕ[<��a;����8�SNT^�dd��G(�Xh�{+߉_ ��r)ભ��p��]��d=U�G!(�e2w'$�(�=�3����z3��m��:Aⰴ��	4�L-m%�dl��]��o0ZwG2�8o��,c>Ò`��Q�a�<���0�#m�p�R�BEd� �:�LEq�"�ـ�$��DE��i�b˫M���j�nY��>! � ���
h��m��a�!�Rj���D���\`�~ס6R�`�:��=r���N��\�u۷���A(�,�K�Pu�3d`ݱ��!='.4��
��]�l��C@���r�G˂W}�8���W��E!�kZI��Im��~���%�g�A���ʘ��
��+�Y������1?x���a�~��!](��!B���M�Z���E�?��(5�+)=Mo�Pl5p�G�����+/�x�x��m͵r�_h�/R#���"�2��cw(�kg>������6����Q�f\�q�:֤ԓG�zKh�3�E��b4h�� J)6\(����	��x��)�*Y�j�]�5�I�f�'d�Qv{�fY�w;֛�x�0� �B�ȵ���2��,3���3�u��nd�iy��!�ziZ�5tG�/ˁw���~��Q��⍉�]�QiDJN��-c:4	���qsӄ>���1 �7GN����;U[Lj���IQ�p����R�,a�V!e嵒��{�>����T��~��獨�l��XQ�m��	���C��u���:��������ɒg��a�30�]䁲���(��(���.�/����:���D+ȴ�q&֐�OO7����FSM��!�A�5ce�2��.��Wʜhʆ��Ĕx�v���h�4J�	���C����Z�@�v�[7�%����(�-n��7�i��� �0�z��$C{��Qh����5�Xü�j�V�Er9ֈК=%�+�rL�l~�4}��|=���п1��c_���e��� �C3Ni�(8�)d2��8a�3V4,h6��\�%@�.@�쐱��)����r�ff^]��,�!B���g1&܈��	�<x�_�<��20%:�JNU�cf������_�/}�L��ku �5s�|��!�����k=��uh�r�ۃZ��'���~�z��	���*7�Zxǉ��A�iv�@r!���#(���qa�id��� ��eҔ�C��M��jEֹP�=:\��ZE�fQf�J������fa�3,�=��yw>���!��!B�J|yN�[ꊋ;��ys�<���Pl�M+Q�v����4/�c��ʃ�7˜�<yzpA=�<����Z
h�t����t�<L9]E��^�0�j�n~�ye��g�o�ȝ���P�5�p)�� ��m+�!�4]5��1樛���j��?�7�_ݸ_���=K�'5O��������20�;������cc`�����ض�w�m]
���?,�ோlm:�M��zMG�hU|?7�傻�(���N&��М�i+�?TD�������vu��KM�7���ٙ���6�˝>�3ӗ6O&���>����z�}�E��>
3^\��IIN���f,��5v���t=����=_��y~8Q�<=׎���x'
<t�0�0�b""pDJ��p�a�a�8"%�Æ�8p�0�0؈��4"p��f0�0�6`���B'7�T{�=�ٝ3�������HN<B�!BT.�E.8�O��D Q��ZIF��(����0LѩGi�J�ЙD��!�Ùw{̙xc�7���)�`�K�XM�X�j���j�ㅙ/�Y����t&e_ ^�d��w���)Y��,C�;h��Q� mBQ��E���2�w�UE�ѢQ电� H�F����5)\��ީ��A�uJ9�G��Vt�=r\���{f�fa|�y���"E����!B�%T���c%h��=�D�ަ�4w�ک�5�Yb4���E������rL����d��i���]I��GjQ��r��B�iCN�
�5�P��d�H�i�@��\�jWa���nN�Nd8����"V3�q�����]��NI���xfY�^��{����)"[�Db$�m@�"IS�o&pek�Y��$�Zq ���86��ۑHf�>3eŃ	�T2�RZ[�d
r	�x!��!B�i�.Z\7r�a��C�Ȓe�p�o�j�)�H���oj����i�j�\z�ipYh�uRxyqB��
��!s��ܭ'�a2�]W$�V��T�H�y4��$�#��r�T)�<k���^��`��kL�(�iĸ�K��0�B�e����6n���V���V)��ت�nT�'s�=��̳0����!B�!J��럵tt�[��}6q��0���#h�P��@����Zӿ��TO�p��Uu��U�k�H�J�Ж�%2
�"ˍ�-�lVKH�1��ߊ+iӤ�����s����N�Ԝ3�tJ<�ڽ�yT�}K�c%K���#�G��!��0W�FM�s6�Üu;O;�lGc��G�}�Iq8�{6��mG,z�S{ڣ{S�Irr�fl�>����z��e#�����d!B�%Oנô��{G�QQ,�>��R��N�^V��.�s�t�Mbr��=���o�����>U�Ѫ$�o���G�e�*���i��Kb^�kX$wI�C�r�R��A�D��T���7�S�����,���MP��J���"�״R��9�i�0�c#�x.�-����R�js���B�u)�b4+G<�F�s�x�3z3F[��E�0yw�T*�#��!B�!*`J6�9�yv�\���7�!��C�F�E#t���R��;=LHܬ.�@�U�7�{��<�E�NXN�I�|��i��Uh滑a�t���YƊ/�^}|{=J�Y�RRp;�E6��R-��q�v�q��5�5���O[LKV';= �I�;���.�e���z�]��T L\Zu�T��1�l���s3.�Li$��j1�TaH��"e8\�:�w��5��eK%��rU���E�3��Y�nT�c�[e���:aB�!	S5�d���.K�RJ,J�t�G&d��*2���zU���=G�%��E�<��W��X�'y'Q*�c��v���o�Ҩ�G�']��I��⦃
��T�4�\p�5t�#kzE�E"��niwK-(��4�����ԦDQ3�t����<�FcK]F�`���1�b�����R1�Mu�;��"�	��%��{g�]��|{]��x�!B��ѯ�DêUmq_{�C�ԍO��h�h%X4V��A���~�O���Q$�AV��yh҈[�M#a���Jx������QW>��~cV�it�*�!��1�K 	)!�d7Lo��y4X���D�h�F�k��3h��Q�bQf5A�j������P0�h�+�u�Z�87;&I�f�l��,�/]���*K՘f͐�!B��`?"=�Z�ei�6���]g�����̎����8ll���#[����x݈���xNn����2Q����!K��7��yR.)$6�h��=}G�#ħY�G|h���PZ9I腔/�6\�R6��A��t~����\0ww��jk$��6V�ʾ!B�!	R���?~����Iv]J��{C��ٚZYD��Y+Sߗr����,�o�.-��~�J�)Ҡ�mV����J���H����䣣���_��R1����<�H�V�L���E.N��F�#��)����j�R��h}��z��!^l�nqgy���北b]vq9�~~~~~~~~V����b�o����l��[���{��ihU����t.Ίٶ�ө��m7��~UЫ�}��
���[S�N'i��bq)+�%A_�����c�zu��KM�n{�߾c�����7���ɏ�t��q#D�,���mX���l�����F�B+���")���g;����ڤIr�-Hf�Tl�R3V*�5G$-4r�\����-름����"�9��1��Mi��H,>�y	�ɨ:��i`�"I�IJ"�R��gR��R�kfI8�a�jY�L�8�)��he����[NaD��刣�0���$@�B�nD�{�W��7�|�k�K)c�-�
%�Hs&S�m�NH2u�RIX��fr(�$�]B`���7&&!0�gn.�^��A$��8�Eo�M�A��,cM�@���0����R�|��`9d�yP���b��"4�DxvWE�A��asƚam"h��#2^YvA���$D��FL�샐��$%P:��53ܭcmVBA��0@"8G�҆HӡQ�"s8�>�۠���-�2�-���f�B�&Bx�K��I%���?,艆a�DM���8p�a�a�pDD؈���0�a�a�DM���8p�a�a�pDD؈����U����z+�f�����\b��Q��%���HdP�%���aRi�# ���V�U1�0sm1��^9��5�,cf�2�	�8C�!B�%Kޙr��d�.K�B�E ���۹�7�<z��9�×A�<&7��CL��H���iV�Μil�F�!���VӦ:v��Q������D��эg�E�d87�o��P�����Z��|�9�8�\�!Fsy�L��r�zTs��y��9�R�(����l�F������3��&`��Vt�!B����?}~Ѻ5��N��S�q����4��Zw��!v�*!��@1��'��."��tƈG.jfe�̛D�|E��*��]�/ϭ?%�3"�9fI��ˈ��O����Oȸ	�]��E��IeF��5kw؆R���������>�3^�ݗUy����Ä!B�!*X$ֹ��{h�����"�{�k��.B�I�.���$\񱍽rʵ��(�zS�����V�a�n�FѻVn�x2�Ք,��];���<q"uGz�r��¾{�ή�'T5�k��<[G��;����BM���o;N��ƅy8x��r
䛓��=|.�a�\�M�C4a��!B�Ҽ]�n��\�2�½t<=E׃߬��D�5r�,�.F�\-�TX�~��ÕtY���I_����(�+Ў���{J��3�ۗP��$�
\�3��+���F�J�8��>�YᖲQ�R-u)u������b8�EBr��֗jݝ}�pord��ve�{��{�ʟƑ-����!⮓+TET�@'�1(��Xxco+T�DM"W{u�ZA�P�ē��q!xY�	�.�ٯ,�f
)�t�"�L$#Ƞs�Ɣa��D��b�7��+5V�ZY�L�x�B�!J���7,�F��Y��լ�6�mjZ�%6���J�u��{ɱ�$��c�<���S������uQ�:=���wl��ꫝX3�Ҧ�����5�]Z�^�(���F�m������]+�5�+mݖ�ܸHYvH[I�&�U��%�(�Q�~\S;Q��UI�/����~�r��=�����fdٳd!B�%M��D�u%k�UR�9wU��GQȕ��fl�]#hD6�9(��J�F�xԱ�l}D��X�E�_��í���n0�}*bN.f7-��o��;��x]G �-m���'6��k܊E-���߂Qo�W�h�:-�;RT��l��w����/�_j �ᇈB�!J��j2� h[E��OK�DuT,
�y��lj��wH�S
��-�g 	�\())�E��m�T~�TY[���"�6��P�s�jU���w�4�d�K�

ݑ%�k	�Ċ$�*;�w�J<�˗m�9��FEE��1�E��1�dq�v�pF��f$eo�-X�+[�C�Kt�0.$���2\��]�x��Y�L�YW�1��2C/-%�L��r�ڥ�HBEI"	��kdjbfc	,m���s�W)4'!�T��@�d)D�4�Q�D�|!�#f)�
~��x7�.����*��G���������)��������ힾ}/���$�\��(�n{�
*E9-���ӧ,@6�KV��P�V@䡹)
�ds	��W�fq�5���/3ÇB�!J�ڔ~��Q'�6�ںp���%�is��#!6��F��eح�Z�;��I��m:��4��<�����F<��z�����td��~�ioС3��KG)*�ڭ)��J�ډ[���Y�л�b2NK
"Q�Z��%�w�|.�^=��>=E,	KH�m����:�F4QI�P1�J*x�HIM7*Aa���Y�7x��q�T�km��)�	(�䓄�\iK�u�{7�CsW�G�B�!J�Z�,�7%��]�t�+uu�A�DD�V��ґ! J�3�F��Q>�<B�x���`#C5�,�]�����7���"��Fж��#���[<�5���[��[:��ַ��G*!��AHLa&�K������{�ʟ}ɼ��߾��n����t_c�|=��^��\A���*XAA �P��jH2�[hڶ�H�{�t�qO+�l瑴{���^� h�����T����g��Dm�! d�hq�;[�!:Z�/Qa�:�s"t�lWWv�5�EV�����MQN�]�8������^����
}ld�����n����6ffx�L�/�q9�~~~~~~~~V�3C��E�������66666*Pߓݥ���t�]��`�b�6�N&�voI����W��O�����[S�N'i�'�q6���/����]�<�4�j�&������͙�z�1E+���vC���1��c�C���8�|�p��T;�(>C̛��|Ҧ�>Z��W0���UƱL��$/�ָ�͹_ �O�~J�w��l7;���!kZ�
r�/R�0u��n�7�ba���8B˛���
/��naf	���,L0�:"&�DD؜8p�0�0�0舚bp�Æ�0�0�0â"hDDM�Ç0�0�0���B""lNҫ��;���|-�>��!B�!*·��Q5�X���e���##HRI��+KH���\���Q+]��x�0V��e䙌n�m�x&�\4�Z��Q�Qˣ��6��4oo���sT�-�9���-B�cc��+F�)�2lƹ�MBш��h,U��q.���]��xa|��8/��>�l֎4B�!B)���cW�n-uXJj��6�bL����%�p�H�[�ʩ�����R��w�m���F��qwMI�	�O�%��ρ�nk�ۜ��k����M��@��v6�%h罱�h��=��{_U=�!�Y��ģP�>
b�$���dB��&$�%Q��Ļ�Ͱ�l�R�Ǆ�O�N����(#)�x�d�L�,Z�2���fd�ǌ! � ��#k��6��R�E.����4@ǩ�k�ƙ<X��|g�Ǐ�ҢN��^�vzED�p����#Z]�J��6���֩Ң�<ԫF�^BW#`�6������F���w�W�v���5�6�Q��O����7�B�$FKIp����H$:�n��|�'��kEѮn�2��n:/f{:/���ڽ�jWh�r$/F��!B���.��8����K��z�E"WB��i��	=���}dQ��P����6���r�����r�Q��]2�&4J���/Q�6�3p�6�wf�\�7w���\�ӆ�<��6�y����բ�ը��GH]^��2�Uy�����L��!b�#|E�#؉G�R�Ѽ*HW��~�i����/��[0}}�~<��Cf͐�!B��r�G���_##iwvYd�n��&�Ѫ�1���'Ƚ/.��m4���c֥��kd˻�����KLE�>�g�:���z�y�F���h����i��1E+p�R��z��)�<A�ãA���ɣDg��	�{��1����l>����W�I�Q։ӧ�!B� kz�F��v�6e}Е>�GŻq2���d3*��6��K:�ln��퍙�E*{["ш��ԯ5-k�+V��U�H��߃��lo�8�m��@���[_�zE�￀UU_Ǭ���/g������_��-2�Q�U��1 �_����!����q�]M�̵��
�de��Je$#M�*���y�Ŗڐ�tۨ�е��N���!B���["�vngKI�3�����u{F%M6�G���.�����1�G�j�Ӆ��E%"��J��+H�Q�@�W�l6r�6�H��f�����6[
ۇ�g\���;bd�8 �0Ul23�!�k{�;0(G:�ّ.����1�?�jʗ*�4h��(��(�F��F�J�qɹ�����=W�_�ݣ�Y`�}����v�b�\|ȑ�[�>�ܿt���},��;#>dO^d��!.�Z�+A4r��~�u�C�+;�mO�ilG������0�S�g_Oυ��ڸB�(��(��!{��.��m��Ű���`�RT�ܢH�o"�/m�,6��imz=�Z2�e�m�yp�h6�5�D#*R4X�Ȯm��9�\P�|�q��d]Q������&�|So"m�#hԆ)|.+�B�3��(Ѹ�ԗ���Oυ��`�W�I�UQ�fQAB���S
��#�O�s�u�������2_��g��)V��̒^/�!��ǎb�/Y0=�G|7���3H�-�'�Sbd�~$#ˋZ�ii3���CE���S��"�h��b꽰�u$�uUl�f������a��L¢1b�jի��Zc�c�ï|x|66X�66>�{�4��v*�����t.��
��Sig�7��~UЪ����
�~^�b�{���m7��_M��T~~�IS���vhW�>׍&���{38f9ɝ��MNPB�!�2��d�*�c�ڪJ�6r�NP��
�;UÆ6�,D�B�Jh�K@$�b#)�Ab9 p��o����P��]VP�b�����F������S����!Q�\2�t�c�E&%�Kd$����=�b(�=-�3=�7�Ki}�YĨJ�T�d����IKgf8�� r��{�J'�j��`���¡�KJ��!�l|�8!BE,�`n&:�0������щR�%E�	V'�B#|����@�� ��v�R�O`bc�s����a�sK�ȹ\Ҭ����	m�i!�.4�Q����%�ai8EE6�d�2)%�˕)e�92���n�S�	����`��n�r�%U�v.4)'���R�Y �ch��H0A	r$\�xW
���Pф�&\�6����Y��E��H$��#e'�Ə�m�Sm��i�ؚ$�|E�%8X�p.�n*d/K)�p�yL�R3R�,���)�0$M,䌸#��gO�x��?~0�0��B""lN8pؘa�a�a��Jbp�Æ��0�0�<"P����6&a�a�a��DDN0���h��ft���{�������ZXE��[��1��	n��D	%��y'H��l�(,�I�J�-"҉ 0�E��c��H��Z��8i��U��r�B*��}8YB�!	Xq�Cp�-����-^W�:��T%��*�N���L���-�&�.�B9Z�� �E'���ݶ���n#�OH��e!��w�8�'(��}�˘��V.�~�E�ma�҉$�w���,0�{�$՟���t��ئ�������U�t�!1�G^�"W�qyY������wi�r�Hٷ�1i6u5q��~d�����������2��j���p�*L��.�dV��2!+���o ���բ	�EHq��������[�?>�/��u��\(�� �5�H�ࠆ��J�az^A�^�R6���i�&�	V��L�Mm>�)�ߗ���w��.1�c��v�ii�XӨ�a�I�r)^M��E�D#k7�sЍ�F���G���ln�Wt\I��[����:��F�\�r�3��2^�l�_E�)xz_�I^�k{�6B""'��{5�Ws��v�w�g4A(�^}�D?��.*�-(���eKqn$�.�����	[�Wy����i���W_Q*VQ>��C։,��%�Y���J�k���1�@��B�kF�g��P�W֋�׾	�B}�=�ћ�L|-�^��$����d&��� ���#FR1r$�I���7)��Q�p�;1ҍ)E��?*tęf`�n9��%]e�`���˹�`�b���i��\�:ՓL�L��)!X)C�j�Z��;KA|���U�/D�2��!�^G�E�Ô��c��u�QI�A��]=��e9�8�@E�+u��pkteo���&���t^�����إ��{su�GDDD	�)��e��i��3�O�FL���Kh�-f�oV�`b-y���Xr5�pcl~F�N�S�����v��f�"���5srBI�Yb�vJVƋ+����A�P�n����捆Ӑ�9y���׾��3�ѭh��6{��_b����a&�F�"""5�.�_(��QN�n�A�y�'A��sۆ6�3.��=������~���ߊ��tH�+i*R�dhV���k�ׇa�%�^�Ji;�� _`3��RCjcV�Ku2�A����2���Y���ukg����s����4�v�����O��~�?~�tsFl_�?>�/��~m�ȍ˫!�"""5�F� o�w8��'q6�"@QF$D���#��Ҥp4��v���v=k]G4��5U���m��(���?uI�Ңgl4*��&�[��g~�Q-��ZM�\֢�2Oh���_��g=C������c@�a��*��"��"d�h2��0�E�ޔi������-�$�����e��;d �M�&-�ZY"$�yZ��<8B�����]�(�W(h�?e�	Ӛ���nI&�i��Z�%mO���<[^��D/c4�2�@m�\[--+g�Ԣ�jl^�]n�ΫrVS��H1��0L��jP0�SF8�(s�p^�X��Km�GQ��5�*M��3e���gp���1�aH�h�3��-#����{���"C�Sݵ����(i�]F��m�Cދ�m�~�_��z�=5A�^�//��g�	�ɽ\����L�^<�+���f��n�G��w�ٽ��V�y[�!����嚵"$<��������E���gl�Y��zQ�,X�Z�eܗ$�����޳�ᱱF�����F���xZ�v*����4.�xylT�q6�D�7�~X*�U��?,دGcb�q8�M���J�i�*??pI>���/Ot���5�}��}��}��>��x.�}2y��3�t�O�M��K�fm=�u���������6t"=��$�����̋��&L.�����U��ڣ��(�bp�a�a�	bA�8pD�0�0�,H"""p�Ç�a�a�a��DDN8p��0�0�0� ���Ä�]������/K�d$4X���׎p2���k$A��9Xܧi���4�����$�8�'[1Q4zQ��8����Fd>�sZ56A�%D�$�)[F$P_�K�^�@�$���֊����M�6�ŵG,<���7�D.#��Cٗ,c�8�Ґ�>/�������>�/K�b} �`���ר���?~���~������u/!$�-�os�.As2+�I�vę(�r���������ޑ�b-��]��{^�Ѳ�у�D`B)M�6�m���c�,��{�ajq�'w�0�M��2:f�엣/�1�)�K=	��kXjnj�J�QmB#��)V��Q���iU0�"S��-d]�&1Y�vdX�0��0�f,�Z�]9Y�X�v��;��.J�H�a���
(P*@�p�pҤX�]��_B�z���m��]m��agok��xl�ST�;��qZ.��t֊>~�j�H����cS��'}�5�S�t�N�$w)��RIRt"j@v��V������y]����%@���.�G�^�/E�)xq��U��DDF�^a�h?���i����Gx�iAۼ�k��c���Q�s��v)փt�[H�%C�c͗��I��U���]v9e��@غ��S�+�iM-,�,��R���!�U�:�*����."�̥j4F�$�[(�Q��)�:ֹ��բ5�s��2	b���5gWmR.MvMhvg����إ��zIW4I$��������'��C��ճ�M�y�v�m6�;��
p1q�|�09���>er��h\M[.�yL�kul4Æmm��H�B�k������)�R�[E'�
��G*�ۙ�jn:�#Y�d��7�y�=|.�]���I���Qz0DDD~6�����k��-�%���7�62��S���"I&ܳ.�S-dd�J��9P����&�D�f����C-J�7��m8�t�b�7��'�"�K8���a��3�}R��h�+�\��ק��إ����ִM�Zѳ[���BW��Fa�X�b �5j�'TR��BT�L.&����ε�i(#�s�7��q��43B�D�3*I��$-2B�n��>�M[p.�WwN�1ZrEBk��UR1���6��fe{��U#SU�ٷ�0���Dgc|1����Q�^-�?9�pE��0���\�q/*S�,C|���Z/���3]�roF�ݗ|.�_<}]�u�n�dЈ�����2�Ѻ=[�x*���+��؞��ot�\�ni�����G�&�����=�w}c�n̻�5��!�\�Љlַ�"!���ER3�E#���5w�v��#h�QO�Ԝ��2�������x�����ט��YhY�M"#�ڠ�'F�����L�y���t"��8EІn~d���������ߑH�C(�Se�v�˼��u���/.p��c�e_���:JգHҝ������L�N��.�3&�;=��|-��>���oܩ����!D~��)��>���n�~�64O~���en�x�e	Ȍ�Z�1�.�����yW.���x�-W}�m�����*ծ� �6�A�m����,�km�X�G⹥h�m����Ncg[�E�Vb�\"�$ǎ|>�x/���R�(��E%ST��)��������f����qba�lM#�a�b�� ����\g��1�}u��"�$ �;1iD�R2EQ%���i"�*�"�"���FH�$��d�(�����$�("���������B�gX�TIUH�EQ%H�%UT�E$R5$UT�ID��U$AT�4T�TIP4IUTP2EQ%TI�wj*J�$��b����"$�F��$��H�b h�&$�Fh��@�I�&� �$�!Lb&	�&����&$���FbH�db`�	���(��� �f"d�FffHI���2f&��Vbf$��bbHZ&f$��bh��h&�B&��f��f� N-3L�4L-4̍32B�@D̐�L̐�2M+1-31+PL:�0�(&��"`�&Hd������&	%i�ff&YZ	���h&"I�CRII%&RI��RaH��1��RRRIHII%!%!����0IHe?��$��HIH	I%!%%���0�ADOP�8�b�2�J@JK)	)!))$���CRe!��Re&Re!��I'%IH	I% %$��RI�$1He$'D��)!)$��������$�2����))!)������2��C
I)))))2��$��������)!))!)))�)	)2������K)))))))
L��0+2L$�L$���2	2	2#0̄��mc�D,���)30�0�	0,���̤��$���2�0 L� L�B�03$�L,�L2�,�0�!2��,�L$�!#2�!2�+2!2!2,2+23)0� L�L���)2��23+2��̓)02̳,�L�,33�2	2)2�!:�j)��$�̓	032002L$�2,�L�,��L��03!2+0�)�L�!23!2�0,��L���̓)2�!00!23)2�	0�L$�̓�0,,,�L0��)0�03#0�2�)2�!0�L,,��,��!0�2��̡�0���Y��Y�&P�Y�&Va!afefdffd&�!afD�I��I�d&@�	���&`fe&	���Y�a�Y�fFa���	����&Fe�d&`&Ba!`&I�bd&f	���d�I�a&a�I�e!d&I�`&I�efI��!e�&`fI�`&d�	ްSI2��2��2,�B�2L3�L��0L�,��30�$��0�0�2�3$�L�32L��L����32L3,��L$�L�3��B�0̤�L�3030��0$�L��B��30�	2L�3�,�2L���30����&$�ȲHS�0�̄�� L2HP� R��,�I+�L�� aA"�L�L��h�d���f@��Hhi�@�&�I��	��`�&���(hd�fd	&��&��&f!��i����	�
u8���� P�0���jQɡ�hd�(hfhiI���hiHi�fhJ�&)d�j`a��)"��b�d���"�H��� |HJ�?���>1�Q�<���8�	ˊ|������BA�PUj$8�3�G���������ٟ����_�?j��A�/���~���ͬ�}H���qC��x�O�&&��3C5�9���_��;�:_�����q}l��A�oh�(����e"��g�䥟����"�)��>��������B�h� �� �E?z��8���G��o�����>��r�&
}Z_���� ���,�g��#�?/�E;ȏ�?V���"��Ε������I���G�B��L�������&&'�G��p��磴9:���G�4���Oɥ�73�����	���bm����u���B���.@���P�1UbMH��
ĉ��������4���Px�؈��!���6>����g�<��@"�Ĩ�LB(���!3"� #��b�#LJ��1�Z>�������r��9��?�	��\? _D�|i-�$���e�?`������ԆQ����4��4/�l���u0����? :1/�*����� ���?��s�?0~@�X��I��gؿ@/��#��/������W�/�HHBG���0N���&���?g�~��8X�x@~�t&)���E�����"��h��I_�/����'簵�>�A�{�b����Yg����|Cl��|� ��AI>�����D��R�(�(@��?O@~1Ҏ�4)�@ 2�SG�h�>��G9P�N�n?�u:�f�����<l�������DS����+��!�� ����EO�5���A	&ď�����K��?��{�_�)��%D��֏�������P�_P���P?z@��	���?����H�O�>&ޡEO�����D��&+�?b?�Q	����������~A�G� }��G�	��N�ё�>΀:J�H?>�ٰ �D�ޏ�t~r~m_������!����'�6��F���v:���
(�r?���~��\��I�>��ߠ?A��@B>��{��0�:��!t:��2lЈ�
AX����NAԟd	���e?���P4�'Gxo�r<��N�@ ��v�_��~;�� ��������Cl~���$��u������H�
�� 