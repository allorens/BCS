BZh91AY&SY����t߀@qg���#� ����bJ>�>    �                            �       �����%E(J��*9b(U*�P"R�� R*���B�)AB�"� �
�(R�R��)R�J�T	�C�e
U {0i�P %J*�
$P	 %���*UR�$
P օPP)EUQJR� �R�����TE
�@�   �GZ�\���l� 5TҨ���tP)�� յHh ;�G@������	�$�*J��"(T�BO    ��j� 1��]� Pg
�IP��& t�)����JR��\�0��9��B��)�L�� 5�s���tm�K�x���
u�I� hU	*U*��   k�������z= v��+���M��ڟ����J�򷝫�%[V[#ל���)R���ka��SG���56�^��Ob���g�yz�٪G�*�)E
 QR��  "sһf�[Op��z
Z�+�O<�)�[(7�gCmF��s��ҩm���=�z�*�3=G���V��tW���m��or�)[Z��*wJ
U���@b �B�P�  ��]�m�gmM(�*4e�m�`Ņڔֆ�����il��)GqX������֚�H��K9QѦ�7Ct��m�r�H%Q͔P"K�  Yz�+Mm6�\�M� 1�cl[(5q,u :�98Nɱ���]q��[m��L)Ԛ��n�+����m�B�st6��B�uE	)E

)!J)x  ���
��º�ma@�:gh��\U�wV�J��R��nU����8mTۧUTĵ�*sKJ(��%

U�(�UI>  UH�N��R���`Uk_`DqbUUJv]��%%wڃAt�P�"e
]�� Ġ��B�J��Q"�  �zT��]�F�Uj�RJ`l*�TM,*�j-R�Q��p.�jE*�a�QT#UPPUB*��   =�$����;TP*��N��AV���Z�
+2�@E�m"*�5YT(*�B���u*)��    
� j`�J�i��& F�#d�S���SC@ `� ��#$ �50#ژ�4���	�S�"RU5Q� �   L�j��	����"bd�F �&F�T�ߪ�T4 41  @?K�����?��DП�_��Vf	�̑qv��lkgk�k�j�a�[s�w��� =�{�� ���*j@v�
�������&}|:$b�� `>r�����&
 *�}d� �� B�K�TUp���:$�T�`�80F9���&�=
s0	�
dO2~�̡�D��y�<�`O0��S�	��#��y�3"y�<�>eO2'�̩�T�"y�?<�9�<�>`_0���	��
y�<Ȟ`<��)�T�
y�<ʞd2��#�E��B`2��̩�� ��|el'�S̩�)�� ��|��aO0��G̿�� ��9�<ʞdO0��S�����?l��
s"y�<Ȟe2'�̉�P� y�<�f`2�́�Ẃ� �y�<�dO23	�D�y�|eO0����T�|��>a2/�\���|�>e_0���a_0��E�`_2���)�̋�Q���|Ⱦa_�(aI��#�Q�(��|�>e0/�W��|���2/�̫� <��g�|��`_2���2���<����ʨ�0�L���*����(#�PG2*� _2�>d|ʢ���(��D̂��A2�y�Fa |��y�� )�A̠��O2(�a<�*y�� �����O����2(>`|���Q��`0���P_0 �e �ʈy��  y�A� ��|ȿ�U�e_2<���|��e_0��̣�����Ẉ�D<�|d0����
y�?L��*y�|ʞ`2��?�?�����G���a��tȠ�$Kkc���bMn��`FTIY��.���o��j4-·f�����sV��X�-M�W;�p��΃#�9��ά��!w^N�c��r��ɰ4&N�MðhNcz��/��A�ՇR]��8�i�d��gI5W�^�B�Zxmg\�����4p=��W>܉��և!�`/$�� !☃���f�pݝ��s1^�0'�Wڊ�C*���,M�|@��Kނ�vѻ�dι&�L��Q'uDZ����.\�� �HPƢ4�����u��Z�/��y�����NZn����>v!�={��xV�;�4e�v��v�������g7��ҍĴ֍ttw[���DN�.�2)/C0r�w&��,�=���B�5g ��PVk氜--L��	�<��F8KpynM��ā��95gN!�0�Z;-x��E�|��^h`>vmX�$��.vW��*	�u;�4�#P8�xk#� ��^c�.,wv\�E�i�=��(�Z�c�Y����H���+�"�������29C��;�E�f��3{o�B]I@F\�<��W%��f�;���=��2b9�����֗��d����S����ezv�R廛e�����q0�\^9v�޷�M�u�×:b����A�4+o2��w��H����2[��*KF��o`��<��+�6<��[ΐn���R�[k��|Wp͝�#�k�I�����*r�P9��^8{�:�����W�:͝-w(XFgTv������{��Cd���B��h�.s�^�Y����Q�l)�ӡ\�;m���	�X��P�Â3- {6�|�ػ69�~�,���Ey�/q�np�uP�]��guI�G�i�ӥB���`{��[��$���4�)h��788�.]��EH�1wp5����ܫk��t*�u�8���qt�6�m�Ca��2I�B ��L��j�K'<Kr��;.���4�Ϋb�;�V�Nj��yDf�qΆ]��v��*�F�Ζ��z�3,m����ӷ����MEE8��xե.��Q���c�ח>t�{WV��n��=�y9$��q��w�֊\q���Zy���#�wGl����b��}ܬ�tŧ+//-C��E^ۜ�o�y�2��gc\k!tppg����+���eΖN����Ô����6���&�ק�P��kۗwؘ5���ճ��Ͷ�,ˑ��؈Cp� �,Wfqe[��d�V�\�Sd�����Y���X�f^�Ƽ����+8]��ċ�k�:s�2�N;}���3^�oh
�I��'DM�frIj��������������^'32�z
���Ɨq�FiaO%�O��xsn ���i�L�v�*쉇���2�V�l�)p\�HR�8.�.�[�f�f���"���h���F����wsA�����6[�:�y�yݧu�z-���&�.��mʫ���ԸoP5����v����n]�~9o������\��e���r6o�&�1��G�N���ڍ�UּN:*��W��;Tw�l����%�2ۯy�X�N��7%	(��%ǂ�W0v�4q�1^=��g<qgX;�#����]��+�E���=�)���X<��]�gMμۃ7�P�[Eƭq�}�b��bFR��'$S�Ni�^1V.���2+��s���`�Ñ�iN�a��U��� ���X�,�vozA�܃���@t[8g?�1�8o�Jb�)���J�]�)Hr�hh��E"�q���l���}����	�|��X�_i�5G��I���Ix'Y�����Zb��׷y�o,�]
IȎ�;7wE�ܾS��sj���,�WuN������A��*H���;�r��L�ӈ.�H/�7*�&;Jg��`v��3p���n�uι\AI�3����0T�SWH Bg;�R������w�ܭYƱ��Ú�C��"�׫CF�����0��;+]؇RE���]�[�&��7�e졁�]1L�sGtq7Z�'r�+��^w�|��N�a�ͷ�mԔr��K�2�n�Xُ��/M0���ݼ'��դ�����tg Qc�̽:v�nѱ�8m�>��+�-!�;�@t��o���g��z��S�,o��숭��u�=���3j9���N��ҹ�=�z��W�(��Ο�Ƥ&;5r`}4�7pRwgG
7p�a2����>[���p�as�ڲT�F"����7���ǋ@��4.s��V�6��n6�<F��ɽUa��+6��:�Xg^�r���u���0��=zy;x^��ʷ
���9ծE�5��s��9�fWJ���m�A���	�2�r͗�7}{�!�4����ǖ-�	��t�{�|�]ݗb�s�dE�e����
��r���u�-,q��ǡŌ��3�Fy���pK]�4��28;rkr��pv>3b���eI2�O����U4՝��f@u�N�hE����gl����A�v<{��^�K���ϛ8��b��V���<қ��4hv�r��Mw��wD(Wf۬����OE�)e3E��O�4��bף��ݹ�v�#�dZ���ֵ���1�;�����X����ģ�J�ݧ�]61M�՛2M�M�{Yj]&$cSy���q�r�n�'P��#,�(Y����;1�vr�rTfE.��Zq��1g�Ԩ	q�:��I�.�hM�@���o\��(�vD�Ջu��FS����Պ^�%{�c��8�O���i8޼�O��<�=�4�k�,�Cׯ>{׷~cciǁ�ʾn�2qlFIQ�����irχ9(1��Q����Ǳ�f`�]���+Y;C;.���R�+}�a!qk�g��������	�ֽ2]U�K4��o����Km��:��L��9_Ls��5�l���{v	�f�I�;�<1�i]�}.l��6S�4�E�R�n�n^�:,�^j�$�55����������kh�����ݧ�=�,��7R�*���;�q2��lAe���n�`es[�z�-8��j�/������y�0h��R�Ռ��I;NS��0Q��ӓp�$�� ��:P�eǯ �]���(�75,u:b��#��nw7�ZS�4�^�w��W-WV��I7��+l�}���ÁZ����������r��7'mW��rZ2od��Ӊ�0�11�� �l���%����0oW�>bC�����=��u!ex�;�L:s�l�P3Nt��u2��9�7Y����s��cԿe+v�aw�-�3Vm�k���x��l)M���y�_��	ۋ�Xh�by.�6t��N\;���M�tM�P`�.gH���3�";q�Y���V��C{��MƤ�N�;�4V�H�xVp�q��v��A.b��9���3��Ĵ�}6�t�t�۸]#�7zJ���HN�k�3淩eM��.nD F�xקv�������_ŧhҨs�^���2�h4��̿<n��u�9@s]r�?5N�۠�xBRN���Y�q!��4B{��15�{�R�㜳�Z���LJ6�v��ʞcmmM5)n�3l���.���T��^�|��̍������v�,kr��X��u�[����R��i�)\NL;�y��-���d`+�+YÏ\*��������ko�"g�P���|e��	c����[�)��&��������3�����G8�m��s��:�r�0��n�;��'i�cx4��	���r����r���h�=Ñ��x�Հl��W'-��Ǻ�ӝ;$�9Wɇ�>;r���9�^�'LE��sq>|�ڃÓzgc)p�c��'p�##-��䘏#LO\� y�.��]��N�t��հ ��@ᛏrn�o{�j����t��j�!�j��	0N\������25Զ�ηW=f�]�v��Ň�\�r5.����#�_n�����g!�t�����)c�}�w^+�n���*�W�-�@W[P���cj�������d�r�\�0���f����\��uӷ!�8v�|U���c�L��4���tr@�� �i|��������#/.`�_T,�X�|�D&�cjF<�!����v�S����
�uk�a�bͮoU{2lÉ4t4����7;���r�$��=�m�{�`B�����f�V���l�����6�u2� ́����k7�/���]$q�Vb�2�8)�4j��`ǰ0��hwV@o�n�;l����8�	'����vY�P��B�j<�30t���QZM��~��|����dg|��I��nt[��5F�&�ĜtQ{S㶮(k��(��;�^�l��潀c�u+��#"����坎��IԀ�8>t.�T|G��
<�N�a�)\���Z�f�r0A��$��h�VLD'2dgq��Gg�v�3wX�>�Z���r��ޠcL-(���5�2j{4>���@<p���tۇ�b?�X�WH8ټukǐ�ӈ[���`ݖ���ǱU7ot��(S[{spAr
�1��ܤ�7x�{�����6E�0c�n�|��"����Z>��U-�&tP�H�voh�f��]��c�=��=6�����f��Z��{^�q�i����m���S���y>��ފ�вw7c��[t��
m\�2K�D��Q	�i3;�wa:�i�b�md����jŜ ÀtUwxA�n���kuw4�:#S�N�t�(V���;:\��r�c��{u��x�t�
(��t����1$�v!�F��G�'pm}�lư�e	�A�������q����fHUYy�Zqe�髞�Rs����[���~�T)�G{�R�tB2go�r�X0�ً{V]��ҝY�q�0��7p`������Б�B�ݺ
�R��`\qG��V���Uu�n}v9��v�{��bիq/Z��F(q����PR�3��Ŝi�No��4R����zf����;sn�1�lA��r彳�+��rY_KM���!�3�Ƣ����H��G�]�����mxC����"��×{;L�w4��8 M�b��8��nZ�l+&Znխ<{2�-��������z!���vJgd
��';w�P_pՖ���뻬��3^>#�3<��4��ل�\,���Gܱĸ],���FqǢ�w��ڳ���0�
���h��v1!"Op�+!Ơ��i�\=�M�U�Y]V��x����L��S��:z�u��\�cZ˼�;�b=~��F���M}{9���R׼Xo@������Ӝw�Ǉ���h�t4k"zb�ln<S7������eN��o�N�)��qQ��9�k��l���&(��9�P��ç��I�+�n���k��ܰ�͝�훚H��ۃE�4u���.@�r��]�4�C�n�cU��UG�^nV�Y�S}8�V���8���4c���@΂�C`��F4k�����5��2j���ĵ�VP�qv,��VZ2>���9udL���уvn�����-u�<D�z���k~'�O@D�L��W'�r޹�`�5 /]CzjM�t"nԳ�
�C7m�B�\��:�Qi�"�\B�Һ�����75i�N�,
�fņ^#h*��y�0sU$� AF���	|M5��M鄻��Z�v4/f�-'7�:h�i�=�C݇����⽇=��"�s��]V��p�9���H�|w�p�X���4&��\ކ�pg��W�	Qb:�kX�·,�F�r���(�j�t$�G!��8�A�]�Ha�Y�к��3p�.�;yӛϷ4>�J���@��u�!�'nNE�kpK�&A���0\����i-;�f��ԧ�g|�#v�X�9q��M2�{v�b��ӲPM��������w@��f�;[��l����g]ĉɡ����u6�������b6��̃tE���<\N�3'A�`�7V�pc�T�-��_+�M�{!��ӥ|(�.k2l⠳�oD�ۭ+��\sV�* ��Q�軉Q�:�]��8\�s�������!a̫xшf��ݸ�'�
�Y�իn�}&��q�]�t�ע��F���f��s�V0�V;^��բ@�xL��a�Ą���oi�a"�ót���q�s�3t�k��-�"�<�ˊA[q�Mttz2�Ԕ�n���YeŜ�fh��´�q���x������5���j�c�IY����9 B=PX5-���z��ݰN۰���q����^�.MӰgN�=x=<�nw-&�[V���$��Q�Y��>�$�\�Bfv�b���\뎩�;��[��`���1-ݻyu��85��ᣑ�q���\�t��KY;tE�D�wo�Z:��g�3���p�ա��(���}����Mm&��,0>���&����HeU�z\b/'dL	paN1l_>�o��[��+VD���D�T.hm��7��ƸG����*4s�=v��ڪ&�2jT^i�y�yR�
��;|�YZ������ڏ.`^�k/�n��.���7{���SǄ�L,�+6�JQW*��0nc�EK!�EB4�a���ef5�Y�m�6�Q������Lji-S��}Ĩ[�5�i~���µ��.ۻ��x(D#'c|#�x��j��$��ؐ��"�ó�J�Z�N�)�	�,Zg-L�F25L*JyY[������n,\O��� �>*W�\c4�E��]+���x��g}/��驙Z��*R"���c�*�W�"�^�t�4�,�QU�	d(���Kq1��
3.�u9F�e�����S�����w������%��}���6��lQ�����������m��µ��./��\��ChB(��˥9bIq�(�!K�	m�.��RƘS�u�/b��CM:Q����;1xͽ��R��Hϖ������������/���i {<���O1ph�2%=K�p隋Z�5�Z�e�e�=���{�kc�|ק���W�zM�&Xo�R}�:>A���!�x-�k#nΞ7low;s��B	]]%���gtwݑ��MN�b���=��b����Ĉ�-��gkp��J4\;��nE�HĜ9J�R2/a]D�io�Mk��c=.tX�FyN�<�
�'o����3�YS�!rMP���C4E�J��;�۳������{��9�ctu�="���m:��"�L���!�������|��K��`�e�/��.���h ��r��04�mX�]'���}����W7�3���H�F���Gi^��z�8N
��Ny���W*�����&�����.��Dgo�����tr��t��w]��Qp��_Oq����i�-<��6�~�i�x+��ޣ���g�A�/$������#�H	���V�s�
�v~s61�wwmS{��J�t��4�\�FH���2�Tf��~�)`�F��k��88�`��F���~������M+�:;GUks��U���َ��a���W�gz<Yo׺Ӥ,�{�o�����Y3�)r�+�=go��[<ٞ�a1�N,X��v��v���T�N�71n*�l�5�m�c�t[Ԇ�Z$�ˌ�n0�[���N��i��
�LZ�.)�3c!ֱ�3�Gp�k{YY:-��7�c�����6@�.ֵLE ~|�`�S�n�`��,�ڧ��f�li��x$\\q_�O>�<.�-^�6�ڂygy�	�>Y�V��=|1oD�x5E�L�¾Ne����W���g7w�����_Y'���;�D��O����S��E�)����Y��g��3�{�zBz�%�����y�B�8H�~�t}��'���x��uѯM@�����cy�y�M�w5=�f��l"�����*qY5�:6J"�5on��L�����Ǖ�5B[Mmމ��g(�8i(H��c��̅�X����i����7jw�ט���C]HV�� te�h��������)�Om���;�M� ^���J�GûG��g�Z�Uó`���x�҇�[�#�wǦO(��,�Ǵ)CT�r�XJ�&u���Ix3dnj�бrfLn	������"5X��PӦ5�]�4��;�)=��2x<E�sS)P�o&��6��E7ed��nRU�S���z�,QK���yI�܅Zk)���g�5r�DU�jgQIM3bӄ%�',�>�e�r��/u�'���O9�x��s��"UF�~�I�6>������{�5wqeL^Ѿ�ۈ�jQLä�b�n��p�F�2]v=���1tF.ŒO4��P|1	�^�c)�aSީ����Ԁ�Õ>��z��*������h��x	�g�0��n���yx��W�P�ҷ���Oq�=svH;H��f�C�"^�Z��.�{L�jS'���A�5��ɚ��UdW�qm"w:jaɄ���;R{.�<x{6��m�'���O�<�k;u-�Q��,^
��y��y��peZ�r�����F/vVm3&�3��.�<�I��qܛz//rk_OLb��6"S;IY�ws�ͶD���RӅu<v{��������QSXމo>���G{zW�'�4��NQ����> ���E���6U4Ɂ�P]�EӘ���i
�DN!�~b �YL�"Lj��:e�wDWMW����0�cO��Ԭ���E�O�{�]fj��q�s��~�LJ�=E1�8�t����{/0�O���m.Aӏn�{��@Ţ�v�x6���{ҝ�!$�7�>���ky˘���T���� �$qN[�4U���{��y�2�_������t��D�(�wH�ao�a�0;�Ax�g�IX��YR���u��m�Cx␧�$C�˵Z!�1�6�.���A\�/}.�h���Izs�nTp
fi%5d�z�籽V�������K����n	w��ml?oY���=�LիQ��J#B��
�>�ν>|w7����/�//�c��|+����w� [���^�=�ħw
+��ڤ��.��G�@�o�\���hW��& �U�`'_*� ���uP�b��r(�E"��(��u]ゑ�Tv��D�p�֜Y��!cW9*Tfb�]4o�5T��g�|CA��i����-���F�$��l�k6�4�ި����R,�;�I�8�!�9-5x�o	�w_f� ���'�1����t�E#�T�+pBǒ��Ql¨���^	j�&��>�ϼ����>�6�6,�{��xf�}=3�L@6:�/CỼ9��^j����l-�����P��_k��t��"܅�QÆȥ�;/Z��F����uu�2%*�?&�{Ӯy����,�v�A)��tPCw٢z���*�P31�s(ӡ���f7r���PnQ���3��H��`�͚A���A���v���ҧ�N�T74X���x���4^�>'�I��˱{�d=�y���i�&����׍����;��[{�d�
y����_J+��?~�<S�8�dn鳷����~j<���2S`[g_a�����H�����W7OUtlN�
`� �Evrq%oL!{Zy��}��/��-֌�<��y��.��#�-]O���/D��t3y�o�����lA��X��8�1޷�Y.åk�Z7gZ8��1� W�Gy3���xAPW��n�k7?H���q��1����<�s��@"�Э���iW��|����{B�=�!����0���ש�k�8z4�}�.�Kf������z`��{zD����Wᴆ�Y�����r���Y����č���~��1��$ID�+ZY��]�wM�+�*�A7��밬��Y�ŸMc�fi9,r܍�E�g��>"��5�y>�R~;���V�ψ��a,j�LăvVNKTp�``gP�w'@~)�<�Y��^��z7�o�(s���qd��-���L�!��V��Jr�BW��#�����E�]�����̘7�ÁL����y�l�'��Di��и�R96;�a��� !�M�]���Ż۫�َ�lV9%~b�T�SZ���;��ܽu�35omig��ڝ[�Dvx5F�o"�ޞ�:�7��ح�6�$�\�Z�S���~��;��>�]�K�d�u��%dy{Zn� V��f0Z���N�n)��::�˝ң��#��fLyN(W�ML�ξ��m��Y*�����4v���s�Doz��|xɑrh�/r�:�ͷb�^��Or��\ ���2J�tW֣JՌ�����)]��Q��\��1n0"p;��)le��a�ݽ��$��R�|Ul��� �Y�ꅷj��-��\/�8�p��s��ػ6�^b�5u/"KѬ�3�k�9/{��������ml����f)H����1���}��B=�ە`Y*4c�S�tj+E-��,s�z��.-I���t���1�V�����h����&ޚ|�5�{�������׽҆�a��'MRv��E�G��R����bh�z������cg�w�b.����o��Uw2�g���D���-���K$��*���U"6e���sR���Ɉhq涞����|�N3��n�ዋ��T�ny�����Z���Rݪ[N��G�j8�m�W٭Y�+X����A�#Izu�*R+����=��p�|��*S��g����L�>ix�t1V����}�:���AO��j'͏n܀+�%��Iڃq$�X��ac�2��FS*�z;w�祔��Nz��א|�-�0"F��Wb�٦%6=���S!''����^�]�:��oAX�&gM8�W��Sp�D��^��	q�Xǈ���.3��'������.zY�[�˓�Ź�=ո��}�ڮ{���¹����H�nu�/F��p[�����|�솝�s��oR$F�=��Z �q�+vbrj���e�d�9Y�#Ż�.��龎7
]s&����oW�k����=�z�"���^���;Q�f�8��蔇��dy��7ڽ��Kq]����6���l+S�y:)a{{���Hz����؃Vn�Lz��}�/^9M^�	D�ܘ~��q�l���'[#Ss��*�Ȅ�%�&1�V7��4��:ʹ�3aU3���rA-��	��*Fz���D��!��� o���d��Q�×f���<�N>�{�����'�x��$�{}�]��A詒��
кg=*n;���۟�#��f�l�ѝ{��,�0�@�{Y�sI'���e�L9� �ި*R�Ĉ�$';��&�R4ks�x�:U}0]׭{uY`�4.����Y�ķ�)`��4���\~`��m�ͬ�F0��rA�m�oS58�O�#P��FP��[ e�n� �lM1n�²]�vsO2ȝr�⽽1�M�g;
�R���7����SN�(�oB�W'>��V��}Z����_�4*^��Μ?y[����I�x.�MX��{���<�3�
.xk�p�{�ԗ!���Yq��M����-�6���e�j'��^H�;�~Ɇ��o��I>�2&^&���튇�o�/C���٧}�����o�.OW�T1�/M�ܝ'{�:�x�y'!ƽ�yϷnOw�m\�o�[{B:%u*�O���=5C���i�gc�;�.��� a���o��4N�Wv.ٷ�3���������<������%CD�{�ua�S��q��h�νʙ��1]�5}�|Ǐ�m�Ї(9܆µ����a�0)IUC�y��^� +��{+gs��4�n��B!�v�3��;�������=<.w����w{n�sZ��L$r�x��m��m]����=5�<�o`���)���%r��}��y�(����W�.���
=���j�7}�r2����L�ʡ=�!�>�ޘ�g�J7�{�b��l{��2&��$���ɷ�
(8�*q�R1e���E=2�L�^v��Z�%c�������V6�A�f�Zkci�ݐ��u�����6G�M1�;�K��4��ǧ0��N�|��oet���TmĽ�(�hN^�CQ52c�E��+Hd���;�tGީ%wgs��������j�o�����U\����(u��&���j^^��z�\#v�[�,&��۵L���R�+�����N���ꂿ����O`���#��=����D�ն���.\��U�y�����F<��{��9�i��N��: ��+LLQ7.�C��Kؔi_�w.�S��}%�z��̍=S��;G��8O|�/�G_�>�x�=��{�8"ii�z!�Wd=�(-�l��P���	������ ����M�<��Ή��S��F���u�Z�wxF��������A�h��f{%��x����Y:.� �t#v$��wt���
�長t�ySɂ����29[�P��D˱��S����=��i�s�#���qUJ�մ��)(S�\��1�������� �-��1��BM�"����n�y{w=�2]�gB���
����e5
>d�5��Y׹��}�X����殶Rk�U�_!0ب��\�BJk��ykIt�dL��(5/3�n%�+N6�!�%Y�0�����"kIl�b����y%�������M�[�Ǐ^��&^��z"�N�Rm
�ź�l��M���R���vNqq��[.�D�������������@YVvx��Ӯ�w���`��W<g��'�B���=#�I���]xw��1Z��9�ŖN�Yk2� �`I�#�%��C*�6\����o�;X�ߏ<i��3-rEx�|']�9](�u�/�f�����u�5��J���04��.��w��vns{�1>�}��y��E"�f����Mo.���]�V'�����sz1�(��O��9��GB�
����{\��
�)�核��M���3h��PR����6����Q[����j����n�u�Hù�mm`J�n^�e]��-�3�_b��]��ݸs�d�&�R�I슝� ���ǣq`Jw��P�����k��kmJs03���m'p�ڢ&0� Io��w�(ǖsRn�H�)��i]��Y��C�8�����4x��6�ec�܃J�l�X��t��3:�r�r�$�q��b.c-6�k�����z���������^�U�:i������sa���u'aJJ�<-})-m�'����f����d�f��o��������h�Hq4Ӗ�r] C@����C
Q�pD�/92Sm�M���s`�NPw��_+t��ҍ�{���ѻ����jG~���%����#q��kY���8��4f�3V,��ᛵqd��K�p8.ےHS�G�')�{Gtޘ�5ZgZ���$������N�om1�V�i���T;F�*٘�ҁ�����0��S�r�6�5�Kr�f�zi)a�LUh�vr��ɨ�̤�v�f�3��L�0��=r��͋��Fs+Ki���2�m��m��oL���Z��1�k��ml9>y�Q��	�� 2p�b�7�8�<<9�k?Oo�|�t��/���c���s��r��˶턫pa'��� Ʊ���X�����|2�G��/0.8����s�����X:;�w�1]HI|F��K��T�ad����#ĳ���ǌeI3�G(��5��??������2��c)���XIG�bc��C����, �F��R%t�'(�DD]��n骨���5��x'��f�R*�������7��|6矱��x'�����?��Ȑ�ܛ�a������yd!�W	��Ӵh�I��$������e��>�s�b��\t�E��@�3��-T���~�Y����v1���]8M�'�^2���
��N<���Ou^=7��lw�6W;�����$Wx���q]�f�>1�`���z-��]}�,'A����k1V?�K>����)���"a�ۖc_����1�p9��:��3�u�������ف��o�a��+��~��h㹒f�*Zr�9�; i9[���P�S���׽<]#���WVk����n�u��AN�?��,�a�q32fC���ߘ9{�ܽSK ��5��d��&5��|6�rm��ٻ!�;}��z�f�(��.�攤0���7N������l�U��F�o�ԩP���=��=}֢����:l�ƕ�#��4� �&`G�pa�r��z�le�3���2qt�0����sp����jz�Uh��5�r� �Vϡ%�î�y��u;����m�uI�bQ��(N�ġ��L��0��t��sE��99��:�R�T9;��h"I�(F'k*Ŭ�n�6r&	dĤl<5E�!a�6��y����Gf��{�S�v��R>ݗ&�\��yY�_w��U��,�x��#�t�+�3��|�{�} �?�9\�P'*�*|1�x��ۉ`xp ���u�&�J)Y���R��؝���hoQ���f�_������p$�Ӈ\Z7W+.�S�u�Sҋ��:�74�l�eSHk���n�;��X�x�@��ygY�"��2����)`=�C0��ԗ	����.��=��sp|�É���}'o��v�|�_��lV�u���� ���{L��^h�ô9���Ǹ,�'���O���r��������لny��2&񵰫���g+
��;NcO���_#���sV���#�h�uk�\w��e�>��=���T�^���{@<O��Q��z�7-UW��v���1�4H�C���7wݨ�W.�5��sf=]�7�x��,^<����R9��(�r��=����c��I���ѹ5b�p�.3wz���}��	J����ǎT X��	.�.�L�Z���|=�d�ߞ{8&��!]�pgCt�^�&�M�kssȥ�:}�r�be,:R����?C]�*�V�U���=Ql�wH����=�[��x�o\o"��K�kGoo�*�O(��e�q�n,uUS��М7;���	n:�^�T���_��'�t��~�c�^�s:�L.�D�霡]5�e,���]�Ó'�_V��鸷;�x*
T2�
3s|�{�va����ew4�-��{g��E-�/FW�GJ����=��=����\-�F�'S�MgƯ
���~el�!��v�,�{TT�-�[��zlbY�Ҧ��c�=�R��X]Gdy�uں��,��,�15PQ�pV��H��'�p���tOn�L���N���Fg�g��{6zdmg��"�c�Cs. ��M���d	�ɴ�էTj��v�؛7a�ף'w}����d��6�{<��T��s�RG�����Z7R$����a�����+k�Sn�%�xD����������W�8rݱ|���*PB��vT%6F5���Tب�z�}�j3���%�⾢���^W\��8���]o�9$��W���6g���g(T�qkzcIf$�j�;��!Bą;��	��l��ʂ���A��LٵA�O3��4��p����l��;Ƈ�x��GC��<;�MÇOz���7_f������T٩f���^�K{�{#`p��I����G��'��������Aނ��x��{j��n�A�0��7'lD��EW���]����a��������iZB���oOv��T��f�w�j��vt�fQyfp���b21:�dR��$�L�!F2��f�6�����!T8,����u�F���E�Ǟ�����I0�������kr�OO4^�ZU��g�j�� �{�ayo��{tе����<���#w�W"{�'m��W���ћl�{~q��������Qf����aC���R��gۋ�8�r��oz����;�5��R|��{�m��.�G�)`�m%����Vպ��gTY��$30o_�Y�LGjV�G���M��c�P���?]X�0ژ���M��P$����'��ulC"ɓ�Zun��9y>�g�,�^�5����>1k<�yH�=�&�I��8F�pwm��^������X�/�X�����e������.V�A.�7��"�c�vR��ò��h�6I��i�F��~��8�R;B�"̻���p9�IM�=����yf�{�#a"��7%殮�x�R#��VS���$�FU��"�3�dƬ�/'�v��G[&r�9iyp���-D��x'}����Oc�V+�rb�^�����nm�)�F�T�w��wrvf��\M�x�>���M�4�}ʤ�$d��XP@7�`����ћ�n)D�_fd���W�Ɣ�I��;��#��x\���o~�tT�0������=<6g`��2nH��7�=�������>ƈ�n�xy2f�'51z�{�/j�V{<|�����f��A�W{=e�wA��YJ�&A�gHrl�l�+�e�A������ڣ��aL�x�y/z��Ac��4t4(pp_,�+�[������9�hX�o`9�
��}cH��C\ݘ
���zZwwid:L�D����l�p�[�����)��o���W�� �h��J(�{|�{��[e��v�i�8�Z�nЎu�K��������,�ׁ���z^�h<iLU���A	���I�1%�&��Ѫ�H�*v�i+8ٍ��Άl<�� ��F����{ �l�槯	�>f�8]k�.���`ޯ�}O��W�E&��3�U�-�.Ud�lū�z�P
���O�����0�0bP����u�Z�׌��XAs�\��ݣԦj�bzlr z׻ӷ�	i�}ƋGopm�*0l,���wR��5���B����T��t��k��'ŝY(f��1�ua{�1�<�'��z�hT\[��,������m������;�I�#��l����₧�	ԗ���g/<}�X�9��X��u���|�g���u�]��<�m��Lo�eh�SN�Ì)�F�a�3��b�gxe垾�$<�y�w�&�	�Ӟ{�݋�0#,I���X��{p�n���x+��i^ z�w���5=�3�,M0�7D���wk3�' �;�˛.����i� �-F��ͨ+g��o��M�.�}R{�i-?tF�����ד�ʤsuTȏ�g��wƉ����෰tUU9d���7k%�N�%��eU̽��t�m�p�f�-L �guTX�
#`@�iF�j-Y3m�7��?3_zM8��ȯ����;+.���YoV=�Ҳu�60jNp7�:z��/+	�����������q�sK>c�X{�vU�o�'�\�`I�m��Jh�k��26ˍ.�C�f�b��N1��L)w�u��mHG܍�v���sܟ���O/"�x���s�i �jf�&�L��r�"�=y8��}�o�0��Z�`��6�-hp�<��n���������9Tu�V��80�G)'����yq��ZS=�9��yx�ore�y�g��9�hƅ9?75��ғ�3��TK��h����×Æqǧ4tB�ɼ��;��cdld�:��6���3��"��B�ڽ��2fB8��0����|�,?^���������`���2�3\��d��L�	�����^���1�t�l0��V�s.P�|���F	�8z�3yƙЮ�Qq�j3dɮo��N�/� ���ȥ��=����h�F{�toƬ~ӄ.�d�{����~��� t���:}=��O��gu�w#՜
�Sb)��s��6nX�HcO��|5�d��Ai��~9�oNg�P2��N��vy�'�iE�=��G(��tA�M�����j��%;+v����%&c&+V�qn�4�N#wJh�˶��4p�0�^˛�$W��A�8�n���qi����j2{�V�7���x;���T"���#/���o$���V��˯@w�)�~	��D�˩���b��#�ʋg�)�>g<�\N��ԶL�n(�Բ�1�I�pv�UjF)�#+3�r�ඦ��G�+@��~?7��I/���������Jz6Wu�S�ک�go�/���vk���[��_ ��L�&N��!�<�\s��gvS|���	��C~�Ȍ������|Q�>�$F��������a)a�A*�v���rb�R�S�7�WŹ}�)�M�jHG���ƧY����#;���M	�ۗ�J	sٚ�K~ֲ����ܽ��5�g�r�q��?g�}�u2�����P���5-'Q��8�#0�q4�H"�AI��vE[X�9�������94�F���z�������~g�)^�IF�"[��G����e9��(q���������e�kĕ�|ht;��<P�	�q�3ؼ�#����!�JV�z����1|��ǝ����;ux�(]� ģ|��pR���5��[���Ϸ���ԃ9��,/{������G�{�s�Ú�^���;'�^�D='��<�e�9�=\�{=�˥=�]���Q�ċ۝N�ݾ�0�T�q�5�os�ڶ麕���x�ί=�b�|������s�I�f�5� ��+I��;rv5m>	n�����(��x�۲�h2���=�#���C����Uͭ��
)ae�Ma��qx2���Fw���>Q�,0Y"���� �Ҕ���/�{7.�Em@�F#
���`�3]����܋��ǒd��{{�NNt�R��d���9!�=��-��eO����#�'�y�OCX�[�L
nwb�776o��QwM�ۘ��[�NfI��(��� �6���W�w�_V��}Cӌ\�b�Tlj��7���A���d���=I{�hGݖi�>�_����[:��=����������v������+��!���wdA���O�rpy� x�/���1m8w5|zn��K'"�u���\�����@a$	��<"�@)��]	h��TI�aTF�&l$u15�g�X3|v�̯�2{�V�5��c��;����r�Y���`�~�׻L���ɍ������T�3��r�%h�*9��3.�Sڭܧ�hˁ�.��B�a,t���q�Wcֽ��/hr(��#+1��b&Е�4f�'ְ5���ӟ{hR��F{����Kh+Ӱ�&�������*t{��}7f�=琇/UJ�L��17
v�Q�6�'*A�ax�y�v�����ݒ�V��Pq���z���xx��J���w�-�[ X�SS��*:-9�z��st�L;����'S
�^Ԣ`^-uLPxzN�J-: �/t,�/d�NiŔ1����!ԞjӶ�L��P�Ҡug.Γ�*�����;�݌Sm��ZcK�+^}+-<�{	�ޔ��v��j��8oM��-~,�Am�J�c1cۧ�����D�QQ����xrj����0>��7޴�H��e�99� J3��ϱ����8��Qݽ판�oN{�'Lpc��u���0��u��	v�3V�.6#*|�o�����~��������<S��3|��5M\�;��4L2fbu����ۋ��S�CN��q�F���z�OMOE�{W��@��⦱l�=��p��雼��y}�v�Nm�Û�Ҽ�F�x�⋜���V`����{��n<}g�虻��ړ�U��l|�#7_^��܏���IOϘ��6�ˑin�))� ��M$�w~j����{�0q{��X!��ɒ��%Ð���dk�{c	��t���]R��~���w��������5#���
�BfC��x���oC�XV�Nޅ�&{.���w��2
8lR�Gp,7�J���l1&vaJ��U��DF�c'}5�y�Nl/
ɶ�w�����A�g]o�sȭ�r|Wof�m3&�ra���%Qb8�D�e=HzG�Y@�yѷ�;pzj�#�³���`\�Wg�c��=JXx��[����G���l��|��lS�b��q��/�ˋD�\ޘ	[c鞩C�Jr���d�ON챁
��*����/u���{�����&��E=�ܳ�w�9���ށx���4ދ�sG<����Z�S�������,��!������bv�\��4s�LG�K/�{xk���ž��l!��ރ�LY1R�v9/�f- g�;ty��L;q	Cä�$��9��Q4g�S�~�=�3��7d-zX�K/r06�zP��^��/[e������[0Ő���/Il\^U)�Y��q��;OO��}�>��S�����ܝ�����͙�N�=	ܚW5��$T��{�֬ޤ��OIU��6�-����Z��]X���ed2�8�OA7����ٰ�홣ٰ���!H�w����i�#㻇���l��F@:���/�0�w��T����B�D��{U���/a�-kn�p�`E��h;x���tg'hY���}�ݽ�/�t{��q�&��Dǹ��'f�n �V�s������#��XV�f�A��z�n�1C�UF�W{���&��
��f!u����M�jkw6a�{�3-M⼙m ���$k>�)�]�ْ=ƭ[���;TM8�0���l����w��u��Z�����9h�<�k&���<��bEn�Wۤ� v�Wn����ε�n��n�{���f��0ٳf͛�4hѣf��F�s�2<,I
 �)b,&0��&�)* �-8%8�ł!(��x���.|���'�jY�6\�ڳ�U�5B��[���3�&Sj���1��b�5�;u2l8��(Pػ��0ڕ����m�Y�N�����/[�1��]$݌�%c����fo[�M^��_n�� c�+��lY}(Wv���a� 綩�Q����\��g7�mQh�B�!�`�=�l������W�{�	�����9��p�3�-�SL�j��u����^�'Me�0]hVKӑq�e��[��i�۩���N5e8��A�ꢉ��wHoާ�*`؛��ȝ�m.��&��D�Xu�P�7���H�䆃T�{�R]^�Jy�a���xh�����q�U�ˌ���ύ�**�(��H!��sb(w@���5�}�wb[��j��X�n�'����0�9�=	\��ͩr��^<�c&�y�:0V�wEْy{9o�g�r�����)Q�$��YP��	�NP�HR�`�Yݽ�wiN�o'a�a��[����V�̈����9��-�d��*�d`�+�����r�g}<i��G��֭�p����_��]�<��'c��E]:����6M]n{���.i��`J�K���/=��OK�zOyq�kƕsI�yQ�7�tˋ*��+&�5=��|S��z�y�r�\n�0;Ѳ�hݙ��w��!W��{EW�w������q��DFZX X�X�	�XS�q�q3�`��y6FC"LcĆ&NH�a�1��Qc@���Ç���C0���d�����>�w��;��E=mo��I�J���T���Av�b��X�.�4�DE:6���T�IQm��cTt��$�����λ�v��"�j۹�h���MQ�Z���UE�J�����UŊ��mAb�]ݺ�v�X&-b�U3EQ�M���;j]jf�����7vy�N(�E57c�SM��T�m�����4h�"
6��:tέc�j��v���.ڠ��j�X���QET�S;:�f��4j�
���E�j�cY�62S4�m��:"����gI���F�DK44AUA&�AN�ccю�v�l��vu�]�/�݊��8:��h"J��X�g��*��m���X�����1k%Uh���-�gi����v�Zٱ`��q�(�wbZ.�ݮӷ@qֺ��ckh��b-��h���WA�]���њ���UQ��lb��96ƌT�[�"�;fj�ncF������Z7n�����]�tnݶ�6;�8��5����o�1��
1 ��
�5?G�称=h^*��X}��)A�C�N�[Z����ӏg_q�L:瑣=W.�ek�K�(��+DaP9���i�5��f@zx��}�ߦ�5V����S��-�fr
WO~��PX�F'/X9��r����� ���Y�qo���E|�/��h��n1�t"k�^u��l�]�<6�Xs=!܎�����6���8Ԯ3��3y����KG7��{?
��}��Z��;�������2������5-�9O�����rr���]��L�d��AG��d�C��=
��^Mc�I�KE��Y�oͲd��0�� �.A�;he�zʄ��z��7����mNg݇bE��Ot���|a��q��ǷɧSod�
$�����f���v2����	vv�pV�`��w�z�ݳQz�ە�&D�sØV�{�]������6;U�݂+�]:��e�1]��	�[���80ی��_����'~�f~�z:c��\��eh|����N�)9�g+�lLgtб����n�}��qy�Hk��1�~�'���__b03��/6}�ƅ9�8������;���b����Iti}�����C��֙8�ߓ�j�ԋ�WJg�˹�ء���1�N0M��K1ti^D�q0��|c�Ր��9�_R_X��0�ݒ��j�ϕ0������v�kű�U|���C��U��8v���QW�9��ǲ�Mjgdtj��?'..r�f�k)`���fa�tk퉉.�1c�A�g0H%�y�7�Vjk>��џ.s7v#�^՛�*�5�6A���m�ڭ�}LGB�̼�SIc8��4I=m"�d=�(��go>ށ��E����9J)�s9w��:�Gf�γ�u˛Cn�JD�tf�PY|�K6`U}�Ł��9�E��m �<z�I�~��=C�k�
v�/��i��z�6n��p2���%�ͫ4��;�6�4^4��[�ls�9A$�mn5ӝ��C�0��g]�ǘ��8���q�)[�Q/9���k�;dw_Hkl�Wz��bN�T�p��kt{��KX��*��b��e��`�yy�8�5T�x{ �q1Su�A#^fP�8���@ĩ��P�&M�;���{���d���� ����xB�U�3(�)a�"��5�EH�r[Xd��(�f�In`������-�{
z&���ˆC�b]Y�+���������v콙�.��3�Ogrr	+�`��߫�Y�嶆-G��3���{���i�j5Z/���-l�}�1P�=�	]A����~�y�"��Ի�V��c��<a�0{��be�΅��f@ó���t'u�,�s���Vw+�3fq�px��%O��6�;ܱl<�����*�_O���9�#Ǣ��]�5�-�C���cO6�q�}*��[�u:��
��"\ͨu�[)Dզ�$v�����zp�o�J�d:ϛ��:��M����6�_-&9�l���{��y�=
*�P�շ���W����'LV}	5��9*�T]���j	�+7�5s����l���,U�3S��\�$g��p���p��4��Y���4�V}��d,.�M}���#��ʭl���|��?����q���bu�fk�4�ɣ3��tf���h>͵�].(���a�)ӯ�>K7uv�� ��.�8�9
���6Ss�^U5F�jV0c}|�uW�t�ػ�V���9�^+���`V����GT�WҔPGJW5y��樖#r(fjp��`����'��j�柧�54#�|"4`�N���]P<�<�u}��qߡ��9�o�ݙ�Y�٢k�~]����׹M&˫�Ӄݢȋ"��oW��I��;���݊B����dWa���.�ɬy�8h��$Hx��.�Z=�$�n<hJ���ޅ�����6��p%�Ҷ��"��@�q�"�$+�js!��[�|���]e���[��M>ΘZ�%N�LmC�2�!w�-<zgD��j����ѳ��T�$�ɽ8�tw7���GT�A>f9]ry1v5z�h^kN1A��� ��Ib��F�w<��O;"	���ų�pW�q��G&u�ú�0Q��fq�2=g��rok�NP�Q���C$m�|Z�D=��í���z��|FL����&�望�8��ڈ�h5��֣�w=���U��սH�n��wt{�*�F���ٳ�t�����*mjjc��IH��ETgI+��i��T�����fm@"�BF
*���Ҟ��A��FE��c�[G ede�(�@��f]�]�ѹ1�B@��r��1{C,L��s��}�M�R!���]���w��lL�N�Pf�q�'V�2qR�!�un*�N\foD�`��w0�Dd��#A�C�&��]��������qS��8��an���2�&:Bs@�gb��`kEt=�4&j軎P��w��7��RA�\q[���%s��;��Œ!�lw^������2��'ImW����ǰ2�Dr�[��>�S����ہQ/��.�d��Ѯ[e��drt#s�/��Ŏ� 嬉N/�|�v�__1�JxuN�U��ӄ �+p�EWq�P��������dJ������UW�2��\�pB�E��j�_t㐗��������U��H�2{����K���A�`�9�Ӳ	&[kEK��x.<���Muok���D��M��8z�߻����g�],��㩉W1�Ѱ.�r����/m�ɴ�!ez&g�A�T��iV�~TFBdbYs^ب	A��#��ɛ����q��k�>��6�oH�����^+�F���b諴&*��Pob���p�IF�p�ݛ�SMa�w1yC�X$]}(Ín���?k8�$ �F��v�-��'QM����ŰONc�"8o-���9u,똤d����r:4MNlq՚��\�]Jϳ��߆�m<�7~o��pK��%�[ɍP���-]� �ً��q��LqY0�ŧ��]�>mq��lh�Jܹ��T�]�E��M���'�
z؎��W��+9C��ү~b�¾�Ye�ܓ։�税F�r�Ļ�
َwVCߎG,�=�_t��[ϭ	�*�e��[�p�n�׋b]¹��`=��znG����\��f���S�Do�}�.��6��q���M�f6 ���s]���隃t�vS\&79��4c%�C�������@��foN�+���iK� �$����3.z+�����5�S��Fׯ�2(�{�q��{��."�'������Dnmv@s�`g�!t ��:2cw��� �������g�UQ���Qm�����,{��!f�mkٗNY�Ge䛮Y7�S�T�Gg��d��ҟ�v����\w����nҊ����;X,7R.��U���OR�gE�p��*}�48�[GGz�cÏ�}3��s������=|��pV�-����]i�����٢k�/n)��=P\��3r�Nҫ�Yr�t�{�[{����v��e�l��n}}��L������i�V��A~$s�<y�4�I5A��Z��B��q�d�7�7��o^��(6�.�7��59������DJ����6}"Jo,��r8�<�$��ȉ�*'��E�$+��/��yݥp�o9u+̆��nMt��Fq����L��Ư��S�f�š�f�y���n�i�b�:�r�I#��d۹��&��W	_��,��o}M�6�L�@����4�)=͌��s�Z~�ؽ�6~p�&*<���ޛ�l\r��2CD%�Z\l��Ù���hE��K�3���3�9�&�V=�#.1�}�u-�ydw`�K�{��!�g>n�|�	���bk�R��~���ޙ�p�%}��D�5��)�?O{�����۞�Z�GMc5*�އ�c�;٦)�2�t��D���py��d�X�J;����[�<�F���;��ӊ���:C��Ĕ���p�}����<:_ep=�G�ڔ޸��1Tf�E�s:�ζv�OtU��8Wl*�d:n��>y�&�ڍ8��Q�x�-��Q�ܪj��U(��v*�'�o\}��,�h���ǐ��6�X�u��g]�|����ÓB:�TN�=��Z���"n7B{�p�K�0��j��ă�`mWRɨ͘�V#��̈�����V�n󞮬�sI�anF��w19��y�1��l[�	���D��Δt.{"����������`I���d�U�f��h�����9uWQ�ݭ-a�FDu89De���;�m&w��x��ނM6�z��\��+0�����'��]V��\8x@~ �m3[v	��m��`c�gs�O��B�WWC�.9p���S���}�Fj�����a�&︺8�,�R�ck��ӄ��Yi�_W�ό���ٵId�J7����т+n\Y�Mgž�/�,}����f�r���[r�:6�^Y1LL@�Xfd���
�S��Be�6mNɢ��q�LȊm\Vj�$M��4U9�Li7�+>��k�>ef�����R>��$/�K�?L�� �^m��۾�=��25w3���8jy���ˌ�T�A>f9]rp��'fb�V������t����Opuwo���͈�7vBي���ଇg��K/���p��
 uAv�q������K��7�i���lJ/�__Z��떜`y���'u��㩖�s��Xb7�Yϛ����4-��ݾ螝������Y��\3�m���PT�d<���̀A��-�s�ޡ�Fl4xடO����gt@�}����)+�����ns�d'e�Wo7_�f�h�g��p�07�tA�vO&壽�R��s�����]�V�	>ތ\���d+��Y4!�[p3_Ct��XeraC}@`ߢ�aZ9>L�����w38Pںw��npu]�gC�Go.{A�#`;�}d�ɍ��q��=&��X���?g�:��Y�E���	Ɋ�s�p9���R֮���lp�3�P��ٲ�hǙT�=�˚�r��5pnt��idVE�%���*������$�B�po�Q�"�P��5��V2��sOn6jzi�7��|�&wH^��X�C�!��u��s�m 2�3; �8*6�$�R;sj։�__@ϭt\ ����b_A{����E���^�	u�7�Iv�3�E,�D�k�6�	q�Ѯ�E�5�ԳNP��ֺg��o�J���R���@�Ī�eOйq��(�N���	=k�ή��7�ls�|"VwI��L*�c+c���Z��Z��a$9���&�A�_���H7GI����8FN���V��a� �/3ca�LZ���9��ޘcd���|�>����Q#��-3�t-%�G����bJ��Fcj:+D��DL?��9vB�F��U�2\{�̓�,��9�U5è���9d�����M8N`���#4��}Ζ��
*f��L2Y�';����s��cY�bx�D��	�Y~9�����y��8�b����i^;#�^��[����1�#h7F�8#�_o�?L7����z�~�/g����G��������||||��/g;F숱�L����5���?���#�¢H��,i�F���Sk]�Z�E�֜+��=Ӿ��:9�)܂����,���p�_[�*ߺ'ϡC����ȯ�4��n��ܩ���mM4/^8&��#퀵�F�OOAh��`OTݸ����-l(�"������S�4*ǝ}\�#�NTfɕ� �ܩ LMQp6(�����@ًQ�5���6)�D��U�:���-{��f�s����1Wvb�(��5i��aV�f����',���2ii�m��d3Ѕ�eY@8Zao[��X��{T�v5w�_i�ak&�Nw;�ζ�dVT��$[����tܫ
L��a�z���o�� ��lk�qg�B%ѻ+n L�̀���[ ����Ἤb�)�6�Wf�3��y�b���7�9()�DYˋz�,����kn�3!=$o���)�D�ؓ�z!�Ɗa^=fR�e�ݲb�?W������Ζ-2�$��&]\3.���;���K �wf�UY�li�Р���*i��ӎ�A�x�:��`M�	`�t�cY���ݦ��n�����
�	mKta# VR3�=�Wm�hx&8�����c�A�1N�cT����1Z���6u����f�K����ќ��<��=&еBѝuU��u!���*��{�J�%����O;�c��h~^�u�>D�^�{�9�RU	���������锲��v��	�զka�3��-�Ga��4��,\{	�GԬ'@�¼�ތt��[�]��g����懨�F?��t��^[�ӻK�(x}���+���L��1�<.�ΤnF��-��ձS��M<q&[�J�ؓ-�0ۇ�*f���mh��ӗ��T��
W"�2t�oT�b�_�BN��K����ڳ������v{ �,���Nh��s}�[�&g#�f�׾#���d�?n);˸懗{m֨/3)��ȇ��{%۩�����ұ5���Cٹ�twF��Q=��Z]�e�z{9vkk%^_NX&9��p���5�٣|7;�@~/HҮ��8l��4N��} ��=]�5uo�C`�X�Z���T��v�+ؑ1��}�=>v`Ȕ�x���yH��_�9N����N�Ȕ�h�6�.�nٝ�.�h�s�p�ۭ�`n[2�ϻϟG�g���V��Ճ9�R�m�y/]:�Œn�t1������Tr�rܥ
�c˪VU.TÍ]�������߹s�;׹�p:)��Ӹ&�q�1C' s���$p���){�a|w3���f���1�?f?2�M�����٨��ض����#�����5�|{!�]�������17�i��n��d/٭������t�nHnkK���3j,D���8���X���[\���N�Udϵ�.yj��o�;<&X�$J�h�QS�]}�]���$�|~���>8�a9�wc��Z��n��jZ����n�TV��n�966��ڢ�cF�o�1=�UNثF��Y�;8�΍Dl�Wn�j)��튙��cm�X*��N��Gg��UUESZ,��.�=r�TDC���Qm�TUED�����(��:5T��']tULTD�����5T��(��"�6�S%���b�4n�Utc[Akb*�6�h-�TD�ڪ��ET���h�&���w����ђ�+�n�a�b�����mZtEu��"����3�QI�����TIU��<�V����"��)������փ��*�k�QETլ�I]"�j+Nݞ-�m���U4WI�G��ӱ��m]f;9݌_1�$�v`:zz��워�m��IV�C���1�PPtj�-�m������b펌��A�GlPS�*��
�3DLATMAq�8�WZ���4n�#���Qtwtq�Wn���+l�$Z�.�ض�b�:��Ew"��F�&+1�[c��ӈ��tݱɬs..玦rX�n�Gnݮ"�j
{�Q���=~�}���h�Tˢfv�Ν����A$�L�66�4����u��[�);��"����u�+te��w�f��1�t}����W��N��s�F㣜k�̍������Š�˶�-�;P�C"Y��D�B�WQ��wo9T�M�,���}'ζ�48���D���l���0��4p���A@����d���p�(��;|.�����O,�Ds->C�,��.pUO���fm�䥛{�ʭM�,̽m����tH;��rN������o\�w�-�Ò�\zxP�%����q�������ݪ3����BP�`{�Ԇ�\T�CQy&1�ј�w�x/V��q�0D��pH{ճ�b�Rl�a�+fT����Q�5�c�.��d^�3L��J��T�ڳ j��D�I�b���(�'ֲ��8�5�M,��������0}�O���_?��9�Nmt�eC�*Mmq��nfǨu����wr��'��V&O_w>L��t��1�a2��v����F�I��Rr���)-�Ù�����d���,Vsu�g�����X@!�?��&86���W�`�i9	�^�d����% ��Tt�f�ggx7�Nc�^ۑ��,�~������#�W�bY[؞ɦ�����=0��x����c{N$ۏ,-�n۩��=��
PQ�(�8T�͔���CAMՌ�Pq�Oh+r^�_���3t꺩�F�6fP��שnH�C��	f����#:w��̍0��Q��ɫ����e����cL�b�;�a��|'�Չ��Mo�#���N�W��t��/^e��c�.p��Ȏ��-�[���ΠǄ� 7��n���ny�iU����םF��U��{*=/�dՅ$[� ��S�N�eWLB'-]˻Y�3Y��BҾ���߉���0ߋƲ��=>��Q:dym��l��Ʋ
����d��/.���l'���u�k�E��C� K�چO���G����i�pB�	E��c��/a�Ôm����1�F.9W����F3�����l�[�!�ώ��d՗cp��-�������
g���|æ)Vo݃�}{��h���ѷ��u�R}���c�.��4Pݞ.���w��S�D���{u������?��i�?5�-�v��g����|��z����wIl��lz�NwÏۡ�ءMC�Pj�Fq�6-���-�<�R�<���Q�WjO����ٝw6ʶf������������ʢ���|�׆OV�K*	�z �|�a��9.�@v{
����즙δ�ot��xp�'���(���&>�� |k��b4)\�L)�qm�����鎳K�D��4���=�H�,�q3�c����v��u`��/i�^���b���i|����`���W���I�ɥ=�U�;��<�o�֜`�f�}�m�oo&N�_�`e���y<F5�t�^�s;��v�>K�E����y�w{�za�]i[�&� �ø"7Mہ򙯦�b�e���n������6���~!�d���:?a�b2�j22�[t�\{�� Jsa#BՉT��oD�>�Ο'Aȭ[�K�3�7���h4?���v(8�rV��ۃe�K��R��	�)�^�J��/�.%��^!v���h'1e��-2#�� ��5c���ǆ�[hG��U�`;8�A�t�w.-��n��[jx^�yp�w��(�q�ҵG�* B�b��!���z ��"�S֕�����K�C
�0�%s�R˔^�tx��;�H��D���)�Az\|B���Kh�)[Y��y���L��\���"��2q��*�e�ފcD���)>X}>2��@���)�D�LJ�����n�j�p��`���=Bc^�ʹ3�xZ�R��Y~��a(%픿0�z��^�k��3\�e���P�*C�#��?���h!Bi���Գ-ΒÛ�Ԩ	�k\G��qW�̯/q���&�4�o���)2P=GO^�Z�� ���?I���'����~��,�:��v�;�[u9ڝOl��48��k���vCL���<�˳}�"���b��P� ����5��ٹ��{��:!�%��l�MP�T.6^�������z@���ˉxF����[�@/��F��n�:�I��K�6
� ��usw{���sѭ����F�&˲���Z^�s�g]+��j�SPFIqU�u�sH^=��k����4�3"Z�Z�k�P��v�B��ƍå�j�.���eP$=����Έ�\�Oplx3>!��u�<�?n>K4�ݴ�2�V��]���OmxcFd��כ��VHB�5�M�ۦ�zoC,��9$Σ�55�`���{3N�������=��Q�J�UK`^\�.|.�"-]
)H?{zq�X����Օ��T�w4���g�!64��-0�9�F�J�6�[��~"@M��d&T�B��b&7`1��7mz�ɟ���Ɍ�6��1*�<9Q��G���	����H����-�����r�\,����Wӵƹ�2�&t���F�c֬��M+Iƒ��!\����-[��/����ݜɓ���p3��>]�;��xd] �ʂJ�
~�os��O�����.͹�� �vz�v�\f�u���;��Cr4��i;�<�M�F�O�!�L��8떂�\��p��0"�2{�<I�Sݘ�{g��hg��ܽ1��W��س`i��*�*�z�Y��҂ƗJkL�O� Ԯ{xK��\�N�k��E�۠��`����kL!�Cjh��&q�j��.�Te��#��XWC�������15[K��Ƹ^�'#p�Q�u*�Z��}��4�������~Yz�{�M�m^"����F��-�Wf�g뽃��/kP��\���R�a�i�G&sض�q3M�f�iέ�Q�%y^�E�<�'�Fv9�k"'s?L����8���O$���C�'�Z�w� ǃ�;�_J�l����Q��G�Ы����,ph��6±/0�-�ь���$�{]1^b��ɕ�u��q�� ��XO��(h��\2r��lQ��V�uv+l,�\�}�W�><u>��S�עfy�ǲY���� �fq��x��E�X��y.KU�\�K����ފ-oǠ(}���%��Q>���v�Q^�lZ�X�c�S����
��U���W�tw�y�.�rV=�Fk��q�� �wk<��;��zZ8�v��-�8ܵ��_Vo�{���j:#i]��GC:����-��xb������H���4���,:�WA
���oh��;Ll�_3Q�w��;9�=:�
QHc�PP��22��T�y�b)�˒�n��Pd޽��y�[��7�-Ѝ��Oub,/f��h+��/V��m?O�J)�]�`�J����k#��<��]�y���TF���
��3x���{��
�=�B��~S�+K�!{���V6=A�3��q���	��x�����Jz�!8�bY'�Q�er�&���\�Ξ���A�_/���{¥wO*(r�p��Z�\$!m_עn�5��ګI�Sr.����W�n�.�l��g��x�֛ԙ���*���-���غU9�2��ʛ�w٬�<�n7d����8e�ܝr��ᎫWo��%Y�k��3�)F
o&��ŵ,#0wc,�n�ײr�����<VrU{���vk���X��vJ�>���>K��.&��FE6RJ�Y��e[���d�vb$��1Z{;%B>o�C74�)K0^�!���]����3��$�^S��t�T��`!�q�Gqʼk���ۛ�����לs,"�@�C�	��n{ry����a��&�z�1i�����t�m��֌���!4����#4�O@~�0�`|�Z�9����@���#e�kڤO�@���'w�Ӈ���i�㰤{�uI�(o�H��e�c`���4O�w�6dN�?d���IE�[���F�BU��JJ~k��&ޭ\�T�el[�6��7��na$?`��ūn�I����\�����mK'U�е~Q)�Qx�Z��0��q\����������rw�B`�W1'u=i���F5��t؞�چ/�3��;I87��i�x� ��@�7��u=��[�ob+�#r�:K�A!ڙZdxs� �8�f�Y�\��hA1%�I�`�":f&J�C��>��"Kd���i��S�)=��$ǂ	���Ͼ�\��b�
�G�H홱�}�t	d�ӵ`Q���YD+��x��z�@x�I��t�3����z���|��z!�򖱚�����v(��jTo��h���O&C1q�Q"Nn�.kd5)[��`$}��ʨ(����{�Yhr�=�	蓼4�F�q�z���>���
��emk�h��槗�<˷��yzz����Aou�GE7N43���S�Z��6���#R�\�~@E(�l	Q��
�2��E�U\���$��OLK���˪<��ͭd7�HqV�=簖M���k=�N���+�jRb���b;�f���^�r��W��P��c�\r�d�_�~k�A=Z�,�$k���^ʋ�"�f#�\m�3hI:{ɒӣѽ}P��'��x�U̚��g=�A�Z�	�N��J��d� cd�(��^��wg�UY�|AG3ĈM��,�S $�#r]�M���nt�?y�Jsi����}oѺ�jؐ��֧�3�7����#��ن���=*�c�̈́`7��O���~��_J��I��*��:�<f�2*ޑ&�s Y}w�xa;�A�5��g�c�T� ���ܽ�c���l�qs�������ju�Z��d]&09����'��BZV�AQ|�H��yf�J�س�4��Wne,��mg�0�<��Yc&G%s�R˔^�%%�[N�94��W�(��?>��v���xT��#������X�׶���7"��2q��*��Ɗ��֮݇{w�6y���L��E�ɋ��P�l�vٌ���y�T��"������� �;�{�	чU-g��qt����&~�Y��A�7g�N�������y3������Dz�y��y���-��dA{/�5Ӻ�d�d:���Ͽ�}�v x?�o^Β�gQ�[w�ng��f�}�hZ�R���X���֪ s�f�U]>c�I>^o�hd{g�n�F�`���3�Cg��>'4:��mgQa�^:�x��K���K]5�}1�\��LۈwT�� ��^�9�"]぀�."Bo)m� ���3a?z	���(s[e�������\�Z�.Ԍ�z&e�N��5�-��7O.����z<�R#5�C�}o
�bY��M.��ʃTA�}Ս�L����Hr� ��˰��U�463�����_
e����Y��mwK��R{��Ƕ�{k�����U�B��[�:l�.7��wy���\���:�K-X!��q".=mI�_{FUKcW�)���ej�N�Tu÷��d�6�����K~��W�k�a0�~ S:͍~���Lޡ#���♗_��[�����Lɼ�[B����Z�'n��;�zx�x]���ƚxijgk���I�&C�|CS����2� �^\��
rZ�R5�K�~��י@\�@I`�����ػS�->SJ�bX��Ȇ<9O��}��kݕ��O�a�Z�PtD�ju/hӊh�����=O<����x�����������,��� Z��[��aY�Z��{�Sٺ�K��~Z�/i��a��3f�ب�Mm��P����:�)�emX%�К�xHR`5o'6'3�_����b�?��B.~�{��x�S���{(zR�)�y�K"���OwO+]j����@ņ� Y�"�N�[�1S�u�m�.ar���2��"U_Qw�vEL-��,�<�妡��r��@�e�8w*��WFދν���i�YBuL�|g�N��*�*�u�I��%�.���/�ԭr��{yٴ��������Aq��Lx=>�qk�G�Z�P�K���Y�i�ѷ�����o&�h��!� �|]�r:����q@���W�:�����j�OQke~��3� 
C�sjjM<Ak|[÷:�㡝^��q�>7r͵�l��!�8t�C�~����P'�8bᓖ��dw\�s>�W�"�5u.F��%�!b�;�귴��}:�	���j�o�g; �fp4�"�S�e�nO���^��V�7�x��d�n\bd3ئ9����e�zHz$@:b�t=5�~��|:%�l&�q�}O���ѧ=�s	���4�i�1��V4�cn�$?Šj�2Tel
��aA�w��1��ٽλ�F%�� ���	���|�ǳ��5�۸i�(_Ia�Uׂ���z�&�b�dW9���;�&6Q�z)F���Ȗ��J�>��<��]�NjYá�����F�3{��:��'�-
M�\�B1��
-kG���`Y��MøN�h��v�C��]�67���F�޾��`�N��.�7}�pH�������PP�"�D��kH	�ZA��
R��)h
)�����>��������}]o� �M�r��)3���xs��,r�}<��˒�moN)�˩Ҏ�4j��6��įB�}�2(��3O��)��â�"��¥V0I���pv��jd��=0V/u�go啣4������ޭ�|o;G�P3�oNk�p�E��ެ�ʳ����(d���A8�bX^�Fi�%(�}�#mI�TW(�IѢ��_�綯kmo>M���	.��&>�iO�$�׃�Jt�������$�������өU�,*V�-�6�W
!�p f����hL����v
����F�|s��ѭI��ݘ��sG1�]��J5��ծ7���lo ���"�G�"<�:m�	�O��{v9�����.�
�8��[��];��r�u�����^��<�F%� z<�0�`d0Q�0�s���^�zi��:
v���cv�Ss!����_k�S����cr_������2;(���`�����|�[\������Oef��9^�"�k��k��I��i�oJ��T��6-ݛga�x�"_�o����O������?����������^�h�#[p�w�֬a"枱��.q^���;ّi������N��}�� F�F�{/A��^����DS�����Ю���ne��F�R�����}���X!��JV�M�W��+��Av'�kݫ >Ʈ�3x���P��rV�5oM�e�ќ��9�U�hƳS�6}=��$�A)a�X�hA��
�ۣLٓS�t	f���mvQ��:�2�eN�[(F]�&��0X �)�����Fp�O"|s�K��u�׏�MZk=�#ūSה�w��B��o]��� lK. m-��)��mVXZN[w��M^��<|D=W�d��g=�gN�k+���P��@�L/�~���B� �/�b�zN�`�~8�aܩ�^��mx����ӂ����/���Ǡ�?\����=w䍕n���[]����#]�C���^��`}V[�o�y���&7����<�rUڽ��*
̞��»o�uk���Ti�l��>����Mσ
�3���M��M叺�xp�O����~�]��+9�H��B��A�ނ<����;����;�zxc#�Zͭ���yKʛ�'�%�gk�����w��$���n:aJ^�����|�x�{�@t5���rv�{�������SQ�����_e淇Ah������廖�|��w�����7*�I��w0�L�Ybb�+R�Y%P���/ �PK�n�����F-r��R��S�jb�xѩ�F�,Ϩ�i�RN����ƒ�޷��)t?/e���SJ��}�-�z!�˷�Ţ�k��y��:1Z������>%,Qp��4%�|��&�+�j{�f�_�:\l\l�㕷��X,;�%d�)�b,���4�R��S]�ɖwV�	bnܣK��<y�0���S<��C�	���x;��Y�q��t�~c���"��%�7E����B�S?2��AS@G���~�!�Q�*�<[����q�ibyR!�Z��W�6aT̽��D�E�T���#��u<�N$C�!V�v��٥��{��%R�򾛲��;���'U��z�+TJ"n�NT=�xQ�*�Q�$�����3nvl��W����'�K��[�Nƅ��|n`��2��s#^ZP2�$�F0L�t�Ei��m��R���c;����L@�h�/y`����-�%5����1p�<���ڬj�X�I�w��R�7��qn���K'���n�1RU�2���g_7TY�-�ʧ��6]�W,��߯MQ6��� �4�W�P��>$�vW]�>��� �$=�{�=����}ΎF�Ma^Z��M�e��%0&պ���м�ދN��*W!<����L�ܻzH��X�ܑy#I�)Tb����W����z��p�ɕ��<�2b��3e�X��w�6q�W��нD���O����l���K	�-����7��ٜ�����ieÄ�#nd�5��{Vzсp�V�7!�(W��p�:�����w{�|z"	)<8�<?%�4�i�1�e2�����P����DTFkh��vcb,����m��v�A��+�c6��4t��]�D]h�ѣZl[Z)�b��Q�4�T�ι�������m�qUQ��v�O3�-:ؚۚ"�Ė#lX;�D֎�.ƙ��-j�
�w86:zj����.��kE���ت��]�u`�����N�ãml���J�
j���lm�W�w4�lb)�.��mn-A�鵨����m�i�%خ�EDm��j(��4QA]m�-�b�q6�v�;�H���M]gF��mG`�E;F7]E��]�D�m��j�ݱb1�cR�cb�+�2mlETQ��z�|�N�q��UDh�g�5;����]tf���?6��qQ�n��q=$Q�vx٣�k%l���#��wc�cGI���A�PP}�.��n�)�������ID�Qc��]=ti4�PLQQh4��ب*��Y�Z&�(��)�`�誈�t'ĸ��l��LV�)�f>7���5��x��9�������d�y�����s�;���*���E��Q�-H��E�ҟ�K��r�ih������;���k�a�
$��%Ch4���@ҁ
J���~�|@�!J1 3�|���������Y�j�AE@�A��ѵ���g<��I�0�x�Z�XG���j+�����v���j��"��s�Bo�0dzg��9�H�M����ܲ}xȂApl'3L(D�^y�2�ѓ�Z�^	U��tON��嗭�;�G:��H�	��f�%��P����F�+��X~z�hA1%ٽI)�VF$5ujf�C:9���
|�j�O�dK��
z`8}˫�q��緧�Q2]F�{X�6õ;	�ޱ}k�:��3DQ��e���L�H���@����);b w�A",�H{�9=ǯ�'�4�Tv���y{��X��″1j+��Fq���8ʆ@���=;Ǭ��}o&����6���K�����=��M�T���A=z�	eA#@c>�om�*.��kCzyp��R�]N�n���{��x'�Z����v��u�PɅ���2�A1I�#"Q��I���,��*��t�mf�
�e����x#[�f��I�F���+Y���Z��#��x�����`�#��X��=�_T��3[7�����L/C �D9�m˷�^��W���̃\��ګ�FMm�^�66ߗa�}�Xs^��r(
��B��rݳ@���á_Oa����إ[('���B�Ǎ��I<F*>h}tJ��8g�خx?owy���#�j������`;�]8�چ>1��{FV���a��U��-��Ӛ��+G�{���� �7�
 D�
�?;�������������Yƿ���7H��&��p�|o[C	܁!�B|�L7� t��e�Oә6���"Μ�ш[wvK�*Jz�}{ˬ������lN�-+T4 �k�v��J�n�߅fa�W����\�᠀�J4)^L*�J疠\��a),hr�v�L����>8a���M7UD�$��zf�>lmB &'���s�(\1�n(�����<ƭ]�$x��}`!먦�V��!QIY�4�J\?0`��L�`Lk��[�*��(V�1>Ng��t��y��n���&�g#�OY��׻���º��Q{�z�b5��6'90̰��,9�� ��qS���ѻ�����gQ�t4�0��KsQ��� �y��a1��7���ܸ���MEԦ���kMRv��쭧�Iv��$b�z!�]@�(�(�(��Qg�!��A)��KAy�u���į4�3�x���)�y�F\;ب���P���y`��p��O�ϼV�f��=�n���:_n�/�2S�3���_ �O�;�d�+��4�m�m�����C6��	�g�uȬP�S-R3L�H�R(�l�ܩf�]?U���O	y��R ��EZ�_�L����[�۪^�9�
�Ә~�{�^#9Th$[YZ n��`U��B�	�/�7%��gyJsǑr�H�8t+~�ۦN��o�,�W�0�J :`� 
�)D))iT"� 7�����6��I�}���"5�Xt\=���MF5u�T�5�B���Pg���׍?t�(�]����@�a��}YE5f  ���l�����K��[����� o#�鷔CuEI����Ф��um��0욈��S���@��i.'��z`�����Q|��3w"�vei�=Z��{�Pe_���>�T@kR|��Y�#�P9w��RW 4�V#+=�u�
�.j'�b�ZhiO��)�1,����l��*��֡?*�~Xp�j���1mW��(�nѩ��A`K��W�P�i����c�t�JN.����ʖ���4�5T/�K�oj�w=�b	�C��p0��0��7M�F�N��8����"Ӗ������c��Uw��-�NC�Sp��#�9mi�5�f$��&q�jx㋲Up,Rjd](�5���5iiۘ�������|o>�;B�02�C��6���=�k���:�#�O�t�A�q�r��(">ަ���xygb����Uu=>�d�tB� ��k�o�'�>_w��z7��[�
���D%.�Ӱ�}��5�.���I�w��дVK7H^p�--:���!�bξ9wI��z*�ԭ���E��n�{�Z�P�Uz��Q����\���Q �J9)��N(�97P*� '�	���y	��)ZK9���Y�����H���"U�h��@h�%�P"T)��'��Ͽ�a��8_��a����
S�9�M���u虞j�Y�xņv%�5�����R_*�gn+��з��:چO��������W��rC��Ex�zb�:�;��P��Z�}�����ͽ6�J���pXE��~���o�/5gX�Hv�����H}���8�v�E�r�}�3Vo�w�S\ck�F����y5�NnP�-���=��{87��ZG�p�4P��Û�(��A��=T��M��8��.�EdV�.S5�
`Pz`Ǉ>*���C���DL�:��m6_ZkU�3���1��SlRG(=���1��{�S�a
/���/����Wk�\�B��ۼ��g]�j+�"Skz�0�&�Fi=�(�0�ј�oG�Ac�y��czg�,@�ȩu�5�ۻ��"�G�A��C!O0� �P��9�3�Fi��t��2�+��	���6��l��K��tP6LJvl�0��d��<����J~N��:+�S$����#�YK;��+y�Y9�>��b�|"��2&��mo`���{%�)�]�t�I�9�NU�}>)r��Dk���ze�n�"�E�p�U����2�V�4����Q�wk9V҃*���v!��R��y{�����&��;7�e֗wy=6��T�\1��0�Fɫ��I��r:�yO�{����|�X�>�#����˾{��5��b__��> �x{���H��BH%
�(PR�@ � ��Ɵg�q���nn�r�F4p�t�]�����[Ab6���}܎i4c���"ē3��^5C�z�������׮~(2�K�\�GR3L'Ǡ?H	�4��t�D�1�^�{�J��[�4�W(��=�+�"kZ�-�^id�c/As�Rz���3�; "8b��@pT0nW��/l����-�U�"K��@H�NL�V�I���M�Z��U,��֧vm�����B�u���u�D�̡�G��R<��F�:���'�.�#dy<=k���� <� C�����%M*nz�-T��PǑ}�AZ�ǃ���~S��}�2#����s4��H�u�sn1b�}�wB�i����?}�J)��U52�����_ޏ�U��{�f�Z�#�틟���쇈dS����i��O�vz	�yy!~���@��� B\�a��&9�D�N�b�i�{�1����(�B�{���ޙ�uw,�\x�<�^*m��w���Xk��O��@���<�pV~ݝ2��ۺ�"H%r�z7F}�>=zg�w��A�PJ������3gP����s���Ă�:��(���!<�5�(�n�­�&�����4�0��,��.<��iCBm��*u��">�Bt�\��͡z\ˡ	1G��̯<�L��!W�D�O�l��QR*�9���gJ��j�'�t17���|>�}����_{��
?�KH@� 
ĨP*��>��g+��ܽB�?�����½3r5_����PB~k��'�Q�,����(LCR�էz6��'�����Xf����b$������dՓ����e��������"8�S�[+|�XK<� �&�8g~��.�����E�~c������#p���B8��_���k���U��t�N�/��UxZ�)8�{Fڒ��ş������ׁ�ʄx0mrd4f%G�%\N�����mm&Y�Pm�)81'��z�zw�xa>�#a�O��\.7�a̼���	�[k�U;O�*Jz&)�t9�5�g��FH؝R���T@��W��[��K������� �������R!B~��B��¨�<����d^���θDwܚD���s��e�U�Ffg
��嫂
Ϡ��8����#�"�^9.���y�	T�ó���������iQf�*/ݳ��s�B�ԩŠC�ʘ>�4��͹�{�i�M�����pZv1�L�ڋܘl�'4�^��Ӱ���#���[��#B����i���f��Ion�y��;��Ǜ��a-�����)�,۔K)��N۳S(
�{Hެ'-A���TM����EKR3s�Yo���;�[!���O�k�s�ˋjOm�L�o^~ї�a�+�ЉE(����&�:0v���^x
�4g�ܤ罚��E�{����
�ԫ@� R���J�!B#BP�R!�a� �< oN�$4���0��>�k�0�:L�sqeȳ�xȗx�`<�i�����}�
b��j�����W�LR���#.� -�,	x.�L�z�#�
O�kW���b��-�s�*�ω �&�C|�q����
�Ɯgܜ��;2,���Hr� �#.��-�U�����
2��C�ǩ�|��DʍA�[H*��]�˫Th^; @�~�L����r�g�ފ���6p�8��$�uoj�~e똸u@�3�,,1N|��9�v�/�=�U-�^�ɼ=�a�7�'k��a97������9V�Z��|�c�+Q���������~�qx������w%�F�i����󷥈�7a�X�F����Q��=;�C��
TQ��F��#�z	'(T���S�ju`H8��W�2���A��Mn�����%/Wtx�+��J�T�ϱe��E+I�B�89�Dt���ܛXn�t��h	�Bu���U�脝�˜��ʒT�W��:������D^�t�8c��`-ymbvDl3l�!0\��7`�i�z�}�{"�y��7(��7E2Zf������z;sH?M҉��1�ú5�NV��p5�rXw?-��̈́ �y�|Zab�{���j�g]��ow�G�aT��[>�}p���ޞ������袼���~:���/��[�H����Nq�����^.\�r�Y��G�Pu������>�����������ZJB�
Z�)PiUiJ"D
 
�(�)�������&����yo��kǜ=4��c��C��o�O��<��_F��S�
x/H�f}yjk��I���MU���q.;`>�a�2mj8F�lė[&q��Z��~U��K��i�D8ŷ��9��8��g�ꑺ���1�('�����7Pa��S��4ڟ�F(�(N��953O�����K{[��m�	t�{	A/t��4���6׺-������D��Dqp4���)/����^w���d�L�W��VeRc~	���c��ois�Ɓ��dt`3�J���r���N��oU!��<���|�%�[7���m�ym��!� �b�t=1`/�����ɕW��.H�>���ଌ�>��含w��B�da��y?o�巈�hd��3��'����T�6�
�����g�����-0��=��{9�ANBG�f��~Y���_n�9Y��x3h>�3�p޺�z<�U�yir��PS��� �6NlUO���r�P�-�F�g.���Z�ûM3u��ʽjm�j	���/�ښO��)X"��Aw�}�/�?���R��p������3� �_��}9}3G�kz���\<�Q˪!mJA��zys�ݕ���|P+��J6�ѧh��˩�75�aD�Ҹ�f�v^���f�'��6=H����n��X�F�5�G�{{)x��&�<k��=�9��ԕ�o�ugy���F� g��HL �D�HE@��!�A
�
�� � �KB4��|���?�����xUKh�}|>��Ų����0��|�>���O*��a�wjE)������}�3<���������F�̼�K���<��d^�U�OЂqDĲ/i�O���i�߭�ԛaS�Ufa�B�1�ܱ&c9?##p�Gm�<,mǵO�r��r�������׹b��4{Q��!|�K�E��t\�Õ����f�u�6��]��}%�OuI�1Cs���2���u���k���LdWW��a�D����찋a!�"��q+!s�B�%L�fgM��X��|�P��5��y(���2�K�\�G#���a��0Qm��C��J�q���@L]SGO�~�^ĳd��g_�{�<la�-������<�"��D?�c�@oE�,�NF�-^�w^��\�n���ɑL\���ғ�XZd�Յs�5R�w�b�eY�{}��d��l�D_����(�@�#�/r��/yl#�3��H���0�Ϭ��z}]`�W7r��,%��q�С�7W���zʨC�N�r��������mC'��4#���Nf�/����]����s�G��(�J�
 2j
��V�v1�L�J6q��P�f(Z�C���&�N(�ΗoxX�f�y�������yS��s�{g�w��,^�۾x+=���7�w�19y��s �YD7P7h����t��Uw��Y��鵷k��k_Xw�x�xxe�F�D&Q)h&P	�H�(ZQ�f �Nv�+�B��wEk&�n[A{�=���=(��s�>���&����bl�v�w��Q�yq���רB��E}5�� �����t���yH��H����/=)��ޝ>5+|�"\��E]p�ϫ�5�y(��2�FwI�jM�#{ЌR�\���)?ԁ�0��l��'2���D�������LNVKu���՛�X�#�c&b��Pd�[>�6q��l��.�q�Z�5\���d�&ڈ�K!]���(j�IP;�
$���?6A='��c?"�Q��wsj��s�*�T�k��y�G�B�Pq�\�s����MC&=�A���LRti���R���x>vȼ�Oǻ��״�0gK.�j�.и�x��A�k�&v�nK�	����Eٞ�T��c���ԫXy�/��[�D�64-\�R�\���Ы�8ޏH"1� �a�d�,6���-4�Y���g��7�d�}��L���Xn�I���n�z�o-��B1��e$�P��C����������<9u��`�4�#����&m�t�g�-/Ch�ק~g��z=�O�����x�z���w����z�}~�W�����<�+����cr���ޖW�To�'�n�C���c��`�÷��Uf��1�k��8e,AC��p��j�=�L�q(�^�{4A����W=$��bcB�u�H[F�?{���>����b�f��*����	[nTahҥS��IrCM2*ƪ�}���'MK�ֳ���V�y�G�t���u���4�Ű�VL#�]"�]\��l���}*����_
�N����\n���W�#��xV�I^�_P7C-�[���IF�ޤ]����B��p��ژ� ç�sȐM�IEN�(���;8*��vd��������]���}���s��c��K�A�ׇ��{���`n���7'�7��� ԧvh-�g]�hıZ([�b�_n��!|MĚX]kf!�h�؄��ׇ���>�|�q���}Q��w����F�ŸvX�9\S���FfX�:5q�n�Ǡ�nv�^�@��t`W�y����\�o�{�Ϩnp|��|v���vC�[����(�����FP��&�����j��[e	��O_,�q����x"œχ����#%�p��nbx;8s�],�"��.�v{Q�_��vC5�.\06ݸFΠy�p۾t��7Fݗ]��昷�`$ks��ro�ob�D�S��bf
'�J-۞�[��6�9'�X绎!G�KiC�Cj۸���D���#��v�O��L,�<�}��c��;� �s]]-wn�4����^�&�~���QB�@�l��f�йq0��X.���>m%χ�*_��o��f�+�B��=�����Qw��|z��!�5�ˉ��/����<4��o:��[����p�[�� ���{8�0 �Q>�̾l�nj|Sz{� 5��'��Mz������:�� %��8c^6vt9��|���t���b�`�<�חҷ;��#����q�o���j���]�sܖ�g�R��\�1K��V��.'=��շ��We˧ѱ����$ԓȿp�kn�����M�`�/��6*��ZP;f��NV�Kf-�Ƨ�ȑ�{�i��O*�Cr	�����~}�����w-}�r{پ`�	u�������eu\r�0v�{8	�(����{�@k	�F�~���/&C����}e��m����s�9w�i��;I՛[{��&��;�7��Ff�Zi�э%�1~g�:S纅]\+��Qt�;ӯ0yp)&�y��%�{;'ݝ`S�%Ƽ�ݠ�����c��]�h��-(�b7�6|֯xi�N�	7k~��Ҁ��^��}s�3�p�Em�5�V��s:��v�QX�`�;�ϵ�f����@���/s�&{
W��=��K ���G����߯nnn�M<��3����-n��Zb�*���ٱP/q�8�۩[���9]��K|l
���y�����ې�N��C|N��I����º�>�~v��������P�[miN[W�Nfb&~����������}�:�[`�a�0m����}_��`���!j"b��h�c5��%�$C54�15�`�힨���4PAtj��$�cA�DSMSCM��EID0QM��b��u��)�$������A���e4UDQT�AM$AT�TETTT�5Q1Klj�+N�4��WmRUC�bzMT��E5$�MUQTM���Al`���#A��)�ih4bI5����4h�L3UQ@P4DDQ�E��SRQDPSC%Dm��kc�:��&,ZJ&�)&lZ�*֦�ђ��6�E��J(��ؠ��3%��(k韶 -|�^°�uH���s�!������jᲱe���i�z����0n�wR(��}e��k������?�fiT�(Q�F �
fD	��;���aU���0P߀�k��g>��|�Om��avJ疠����RX���;�]�D������������H�)R�1���t� ��:�����X���%QaAgO1��g��\ᦝ����iS�9Aa�(+x��,;�æ�c�:v`sm�B��D��@�ח.��'��j㍙����/|�x�}BG���Ӝ�b�;�#��(zP7�������Ɨ���}[�qKe�z��'�vf�&a���^�{�A�.���t�zs�Ր��-�O��K{�(�����'�/�Ia����@�f:��;a�ƺ���meUX\�����fR����|���;��C���b��{z��̜!��� ��T[ ��˴ވ�O �ީ[7I6�J��y܂�+�Fc��)=�E��X͌i�Hxj�G9U�Fy����a�ZC�}9Ck��,]=w�Vb�0�B�TO��Z[B�`ٞށڮfmX��C*C%����6�hmCMЮFN8Z3bȊ�-z~�%1��!���7�g���.��@�����),R��YK�˗4��3��e���`|Q��kbT9�Xn�r�:��mVZԎ+�]=���s#Nd� �ܮ�nݸZ�����Hn� ��݉�¡ꨤ5���j/`��Y�ut�7��\7�������ϣ�����	�ZT)E()ZB�hR�fT=�0�����'��'T��P�ߏ�%6�R*�
O`J9B���cռ4�К��GX��FtQ2�l���<��!*���ʞj������Rk���"��]�Ֆ�)�ip��qV���[U��}���X2ʜC�L�n��pE�n�$�s�r�tS*IRaO�|���xr�x�����V�Yb�x'��b�R�7OcO�����=�E�ft�tS,��2�!åW��G:����^4�:�2bǙ�Vg��&���i;�S���]�1�ͪ��L%��NNJ4_���\`���ɄG5'��a_��0��ryvG���酩�\��㖵�(z�+=��{+b:�����R7T��ƘR��A	���7�S�Z�����	�Mn�eb�1��*����*�OJ״���{W���m�Ώ�/���
a_Y�f�KUG\k7��.�P�[!ٖ=j�bA�I������3���&g��d�1a��u�\۶9�f�'����T�(3 ��~�Pj9_,�yn�y����w?X���RB��?�ڧjKF8�
�]�v6�-P	��ɛ�"��3�Z��:&�bs��ߟ�7W���LQ�Ѩ��D(vb�N�Wq�J�wj��\9�BH=�����r�a��6��ݭlM쾛��6����O8C!�5����D\�kMe�~��PF�Qa�?��������4j>H!�B��HB�I0!J�*P}�b��V���Nl�Z����(9�5A#���OB�
��8�*�w��q��vq���$9��MЉ,�1-���3w(��Y��}�/�(k��pS�-!����>��{9����B�R�ѷe\��:K�_]�hV��4��B�).�EdW-.S41AN��>�όp�E;�ŋ�`G?Q��]ѫ�O�L��ⱚ3nPeB��ԑ���q����2����Il����ϊ+Jj.�����coj���"Si0���%ԣ8Ë������̚j#��P�����W;� 8�(!4�& :�A2UsP~�����K��f�\�I���I�d)����< Z���Bk�f����Dڨ�#����ꐵ�$�ħAd�By�z��ry=׈SZ;����;'�����| f�t���C%��SDt�ԇI�����K�y����X������)PCXQa�@�������{aH!�9�jc�m��B��6�^V����x�����Q�9SYt8��HY	�^�&.<��2�K�D�����	�?O�-���F������_odH`�L�T�f^����?���Ov:���zu��d0zݾ\�L���ÓW�j����2N6YzIS�q7٢�J�S��i��c]?oz��-I��Ov^U�QF�x��Pw�s?)�sG�vwrY�i�Ð��*p�V���Ē6����G��  3{���{��\�'R�ݥ˅8����=J3L��3��]���K$kz�>��C���M#�vQ���+�X�����R�P>l�P�.��vL�b��5g��'�Z`��W>�U,ة]��ж���]��M�lC�J0��h~a'�C��/C��k�ƅ�u)�}eo��p������>	,��i����.���XZS��
�׍�l�q�Chp����Ǜz��0XD��sW��k�|�$4�M�zQb�?���^���knMό�*�։����t����IMba����q'DYz�o�D�ǐq.9�ˡ�5o]
��'$��G���D�9!�p��g¸�y���M��b���^�e��Z������~���VT/�U�uVf�WeB�#�q^�E�n<�۝Vԝ ⓠ�ܪd��g���]su3���iA[5W�ȸ��]%)xZ_X}�WjH����\(���9c,0�z�	ez�B[$oC�6��Y�^v��
�O-Y�~���m[�Ðb���8����3������� �]���
���6���R}ᶛUUǦ�����}�cH����"k�����n�v�܇K�/}�*��g�]v;�ay���)��`����چ�2IͲ4Y��I�,mnYV���%͋P�Qs5����=�{�$�N�m5�D|����xa� ��  ^,�;�ݩ��*���1�&K	o���t�C���x7�[Ңe��D����mK��c��E8W3��On��\�͏lyӨ���Hеr�'{=Z½O�khT:q�A�i�:A�ZN�m���G��Y7��]��(�j�l6��wJ�˘�LU�H��&��p�J�22��}ð����M�_n�����r��'��Ƽ/�;O�*Jz�f�@���-/!��U�����|�%E��=�����%j�4!�P���yk�"N�4�U��-K.QzJ�}������S9��N�򼈂�'��ݦ��Sn#��Do�6�QE����Τ㋰J��'�WQi���R�W&���d�u#u�8��̛���+��`��L1���r��հ<�m[4M��UtNlJ���e8+��'��PK�)~a��N�T��C��Zd�����������k�Nb�ޛL����a̵?��S�պ.�����<���{�A�.����o|e���`۰Y἞����w�LeK2N�oo����0�bK�x,�\���^���!%yg���^��lG{���3ٹӷ`Յp�J�X�Y�ǲ��\ޘzW�{��j����y3@|��Fz����7Tˍ�H���y����.h���%�F��i�xz��,�[��M�҅��o�A�t�ѡy(���3��&����9T<vvy5do�����i��3���)
bA
Ti �f  $���~�����@���0�_V��287��� ̋/�	�@A��ʟ/z�l���u���ש��{C�p�	V5���Xwqܪeժ5x��}�W!�C���V���D��������y�\m�5��s^�x��Xu���ٝg2�N�O����2��z�M�����s�P�*���F�Tu����	��T9��M�HBkh�,��<��չ�I��Ehܼ��Gϸ����bD&�&Be^�hRxF�V��ׯcռ4��;G��NM؟9�/_�H�K���q� r��M�j~BS^�JK�	{`XMl*F��Ng��9�}��s����1���0/=� ��5��I�1�L'����M2�����;Qc�!�b���K+���g,�å7���$D����cH�^�]�(�`��.�gM�Ęx3i�.o��[]n�1J9f`����N͍b8Bn�����;��N��2�$��;Q{*;���Ւ�5ה�w/WlsZg���Y��o�0��dd��t}??��r�u
����5G$�Zˀ�n)�5�����@����Kj$�ǋn
$���pw�.%�Ix(���{��=���'f�}�h�O_<ئ�{(��j%Рj��oY+F�1�k�/U4w<����V�����%P��f�ƫ�_��Ng>}�ǹz��j�'�읞��܌\�$��?�����D(�i)D�a� ���j�_-�ͽ���:���e���.����
��}sazp�f���Dÿ��w�^�{�:���>��{ji��%��z�a^'�kߒ�\m�s�L�[1L���j%�)F(�t���9�#��)"yq���'-H��VeRca<u>�3�נMz����c�?0���Mu��z�T�p�Ѯ��1���r��Q�����-�y���.���/@ G$�c�Bʻ�w}�.g����a#��bę�b.��������
�EyP�w����B��N�E�Ա�$cvI��7{�_,����HӴ���Oϐ�u��r`��T0��5~�'���fն6\�6�-u7/T��C�^�S4P�%�QWA
�N���sͼ4��,��斐��Ϻ����i�%�Y��ѷ���s�1�kjԕS�A��(2�jm�d���G{zvކy���N�+���jj�G��vz2z%uz"�==BU_��9�,/���`�A�U�4�ģ8��|M������gl���Y��x�$`�ar"!�j�VJ�jЂq@��E�1,�����[d0�5@�kR�qq%� �Zi�%�_Hjria�*�e���K���f���S�8�RKL)&j���`]�1�sbh>���������{/�D9�nd��)�쫑F��˲cqABj���T�;�^}��,9��3����oϿ���}�]�
��")@�H����YY>�����Vdj��Gҩ(�'��׾�L����^�_��&�'��̖�ق2�cR�ӵʋ�d?��$���ƙV������&��d�Zl3�1�#��{w�Ҍ xC�oN����ڭ�����|��E*��,9�����}��l  �z�M�x.��!حV��Or�܁S��{:��2�'Ҽ�A.�>zW��DL�	=�Z-��_��;�%GNv����0��9��ޚnZ\o��aFu<�d�c/I/I.#�i۸�;]�c�9����W6v��E��|잏L���dS��y�S���´}�B�YD�{P퍗�d���5��"wQt-#��$N:/�uCs��^�Ba����_d����w�^�w�,�>�S_d=��j�5{C�<f��~m/^�O��P�Vm��s�6��9��D�^D@�O��L�h��>T�L�J3��~0���W�,,�wo;�oYL�5�I��	c�[���-�B	�.�4�f����E��R~��$� �}?/��(o�Yb�O�Շ��gB7����z�\��6�^ik7���Gb�4�D���[]��,P.�GZ�"Z�:��%��Z��
k�>�On�cz8����<ÝD�t��2�4����v�EӍ�R�J�ˬ)
Ӛ�Z�������>����#�f xJ��������r-��_��m�oO�2�3EwI�j�Sl�W�v�֤��)?g���S;.sg{�r#�%�P|,#�qlS��z{mcat����A�����3��^���d�����z�{k��}LQ\��Rt<�G�]�"b*A9/4�5A	��zN�F�j�*�(ѭKm��r�x&��h��v�״0J9��<�ڇ�gF3���U9/1.D_2U�F����������C�R|�F�+U&ˮ-��.[�k���l�G��dn_�SP��t.��¶qM�ú-�,�Ad��sPoғ�b��t�!K]cm�}#b������^NA`�pN�j��:��!�e!\� �/L�OuL�1����):D�'�g�w�xay���%��,eݵ� F�֑���x�L9�ݐ%��m�)蘦Eַ@�Ary��ax�YS��fz�3&�apJ��  ��<�P�;�~���dIц�
����,�E��j�ê�a���͎�]����oe�G��K�4��@+9����;�#eή~���Ơ~������רO���&U]�+9�^����Lk
 =>��=�g�<\s�#F�Ѓ�3��4[�"cU��wN�����r�Z��6�ъ��"�߲��������R�� 8-ɍI(Z�2���J	�X��ypVe)��"]��dJ�o
�:mT��D~L{��y��3��� .Y�����Z��/r8�zc�*��L���@���ðB�� �c���C��]�xa�g���Ҋ���[���o#���Oҹ�(%�S� m�#U�5�4/�`xcҐ�#J�o�Uk�7)_0e���T�-�%�7x�T�����fv�MKsW�@��3��.�q�Bw��j֭�C�����9C*Y�:�oK�Iܢ&$�P&Y��2�'D[�aLәw�;�a��������i?b8+��3"��z�i�FdYx�� ��<y�m�f;��d�W=�Nk���vU�-�R,��n���@fh�"^A]��eժ4/����B����abz��D����]{M��H��O)q��鮑�Jv�P]�C����fu���<]�E�h�����ܸ=���� ��(A�WB���p�7�\<Ûئt65��N�Bc�V����f������<�InV6�[����l�	�F�'�nE���c՟D�[�;N�df��q;�Z�*��;ς��N$�P������O5�Re��k\��b!%B�ѳ��{�}�o����yyx��>�w������^�W�������ܳϴ$��bAɊ�4��o���M�a͖b��B��Y�D��W{�� ��x�6˺�kQ�4��ל4���0���N���!B�y*N��)�B5�/[ݹ��ciK�ûwy��`�7ݶ\ӱj�0Y���}�fl���s�S�R�'g�Zѷ��-/�"Ѱ&��Y�
�N��@�0L�����:��C�|�^�;�/�#���8gnL�B�NY��ۡ۬��C2�1li����H^hQ�t���q�Գ|�~2�#�k6�R׋���|K�� v�<�#Gnxt1J~�e;�7���m����/^Y�d3ˇ�]����da��Sc�E����]]�xgm��]�<&���m�uQbU�ȴ��M�f� �l��ͫ��J�3����8�٬�Nr�|s���*��,��Yf�KFF V�r�~���$�r1�J틟MF���Ԅl�fO���@X"�#E��s���)��叆�b6��cË;O���H�_
��}�z�\�o_{A{���6{���[}ឝ{сH��y}"~r���>�xy�����'��2K��v�pT��6�=�;Yӗ�z��;�R�M��w�R���̂��P�(hd� %��U����h�f�YG��Ojk�%�!@��I`hދ�k��4+�L�(�/��g8>��{�q֦(=�9^���Xf��v9��
/���	J�ų6���^�>+[ޞ����@�Q��)V�\� ��v�;��oxm�|��||��~�X��1���]�Ƹ�Ɵ=Y�w���:�8����U$q����ȝÓ�bW���t˕��a����q�����l�Mo�\��w8�V��b��X�Y�94�����¢�8��W�jT$���7��uf���"�qD�t�YG�5n���-��|g�Ix:����(���)�g�a����7��7q9����>�'�a��I��P�uv�7Dg�/z^ҧ�K�;=�.˩lf����Έ�Զs
�r5��+i^����w4��mh�C=ރy8�Q֡�}�<�bJw���'���9�ƣ����K�Id�o!��U\R�υ�ߊ�6Z^Pxu�l�~�.E��5��� ���@S^��8x�Q�/{�M"㼏x���X���1��&��t�,�R�,t${��سx̓�3��/4�Z�:6&�(q�U�z����o���Ӿ�k�k���ia(�����Q���ĸ�j�pXWp���3}s�����u ��3�9����o}�4�ᢻ�s�9�뤨�7O�>�Pu�G�I���z�w��8	렚'��������!]��cf#JP�釬���i����ͳX��5n?Iq7�}:a�>ٍ���w?���[z��++&�3@��*P��˖Xz@���z��]��o�
�/�5�;1��,;琿S�{�sl�[/��gh��܌=w|��}e�o���{���ha%�&nV+M�����o���O݈v�MEE��EF��N؉Ѫ4b��"�F�b-����-��݂��-�D���U-��V�b7�=u�l��T`���$�i�q,E!5MU)�E5l���Lov���) ��*�d�h�ԔUPD�Ӥ�⪥։��`� ����STE1RQl�
)�h�@b(�DAl���j#l��hh��g1LPA�SESERQ[&������t`�����%U�h	���
���DEAD�!A1kkUIF؊�(&�������&�4�&�4j�IUU5F�EE4$�SEQDLU%`�&њ(���(����6uI�V��b""(�*����?o�Ͻ߳��M��6�=����۝�)mb��SKe�/^q]�~�C�>�����l_2!��%�ç����Q������Y5ljT�;�p��8�����Ï����v��Pʐ-T�K��x)���|�L�3�0_��L���E���Wvu�հ�q�6u&q�omK"��y���Æ�k&���Ǥ�Aݲ����rR�'�D���Pe�7���]\���c�KMCu��;��`Լ��
��8Bn�����Т"OT�4��C�e'��)��q����זE�洠��.�̛��b1��k���
а�^Ӕڕ�����9Sӌ5�
�`�F^�Gs�Suo�li����8<#^�W�O��y���Je��{�.��Z��>��ML��aD��{�]�.�N����f�z`�d �1UT�gs�պ�':@A�/���!�9i0͸�/zm��T��U�0-�n}�����6�wr�g��mdz3r���S�Q��)���+j-_��چO�3d;od"���zK�8�ɻ�%���)�u��OC^��������1���~XV���bT�{ڌ�K_�U2�z��9f�S��{;9c����ɠ<M;O����EC��g�!����=�N}�=�W,2r奆�f�;�B�&V�-��(3c2�S�o��Jһ�^�9���|Njby�?ܱ�Gn�O�/����Q��F��E�3��{}�=��o��/]d{���~s�'�!�c��}Y:���3þN%e�'��8�3u��7�Mʥ�ը��n�Z> |��` ����NrO���.�}���i��L�^��è�������z��E&c�PS��|�MH�ʣ�I�ϋC�E�\7W�bG����c���W���֦�&H܇�f�z����03�����2kH�7҅���l:!�1����&��̖u�/0�(M6آiMx�i<#���=�O5�`Ȝ��ɭ�ܟM����?R��ja2+@D>��F��\|�]	pK�.x(K��`�&�F���?wu�.n^�4��7��Ϊ+�M%P<���D܈|GFـD��<���t���e]q��Mf�$�'���(��n:uNoˤS*�IRkg�m|��\����BR͵1���$�<^���&lɵ�R%Zg"S�w�>��4�'I��Rr��E*��7���cK�}�?�"=�{i�b���n����׹�݁[J�,J�-I��`$��.K�~A@�u�*GW�3L'Ǡ?l�<c�+3j�3��]�A��4à�H��Z�ݣ9Vߝ��^h,��e�%�3P���QK�='�K$��[��S��ga:��<�v/ƺ�W?�$Ȧ4 ��߽J|]��ߧ�����n޶Ge�Y!��v�۳���MxMuP��H�[��k�U�n͍��cj�2�zp��������E��zp�qn��!�'j�ͦ�=1�-���;dѣ���[n�)�\b�1���
1�&�V���WJe���llc��j�1����}�������NԳmt[�2����#��H~.����C�Cs�
�plb��S �7.�u'�<�>���k��}�G�\�u:�!��2
�������a�).}�Z���ro.���K%3��&��,�o8)�K$@;\[�\���,Z���xg��9���̫��Co�ŵ��(��5!2W�A���pЊ�j�1i|������TR~��!*�c;s�&�w (���n3�LO�'�z�ϯ/�\�ĭu��3,�4W���x6� ��˵��'����(��m4�
2)����{�b^f��ٛXӊ>jas�}�%x�%
:P�bpx�u�=�+�dY��آ�@�):�����7j���M�E[W�A	��Gr���u��g9�$v.�3��F��m�/	E��g�_Z�T\?U�f `\؉.2���S��%�>�M�Ԧjgf��3Ժݱ�1�IE'V1�J��d�;x_\�:��g�[��3Y�
��&�%��W�yN�/.�,�nmЙ'�1)�FE#*�qv#�Od[B���{���٨�q���2�5PpəA-�R��g��ުՔ��δ��U%"�9E^�.�2��1��L�n���۲�9�n�d�Ɍ���һU��h�R5�z�=���љ����L�ˡd��c���j��=�E:.�7�H�Vc�f����;Y��}%�oOQ�{�o��$C��@ۗn7�.�ҥ2�1���n�I�&A~��1)�g��
���0��.���/�~�0��ʯ�;vL�LS.r�c��*Ε����>�d����Fz��5�^+a�����?a����P��ǲD�2�Ox�ygvE:�x���\��}�]�S�����Dri���AY��{�!1�)��uEs�r���Q�9&�f�gn6*������u
�E��]a��R�#U ���x-3�� �b7D�7M�V��Of�g^��%�������_���{J	{e/�4����B*�;��qL�i�ŕ��,ɬm�]�ھ����_�a�n�Ra�GR�StM��2�c�����~^2
�%��r��q}V/\�I�E8u�� <B�62���W�.�'r�
&$�P&Y��g�P�/�w��f��*{{�+b�p-�y��<P&tF�s�XV��29���z�FE��;��%2�n#�[�s���BWR�����D��-p�~�`KzP{.2}���.��3����W����W*�A�����"���;y��
�L\�!7l�Ǌ\���������։8}23� "��;F�1�*`8۸��N�k���Pväz_,=	���94;Gl��>��a������5�~Wk��Gq�V]`���+t��;"a u��<<�vx#v	/�������C7ϡ峞�?�\�(r5�q���1p�E3���������T��u���Ɍ��󗹒Oo�cu�j���d.{ ʭ]
6�p�k�aC&-�<o�1��x=���N�(.Ey-K�?t��/�9�17�R���D��&Be^�hR{�P��PkE\��j�es�����y�7^S��^�L J�FX�>!�ʞj�Jc~c���b$�Z��j�UA�]t�n�V]���,��}*�dI@yo��*`p/"�p�[��ݙ%�y�Ks
B�����$y�w^+kY�E��qOw0^qcP<��o��S��}�`GH��$���{(Ir�X��m�4f<^�O�J����\s�m�[�nvM�AC6�C��0�؝vo_b$����1�(YC�t8�t�x�Z~kJС���Ļ�l�a�6�Ԋ�%�&�νݣ�Y��mHUM'P��&ф��J�.����
���K s_���E>����)��`0/���:�ԸT��0��yä润�z�'���J-�����h�oJ�Mܳly�����-�E�*�ޮ�*�7݁���nު��˔��(��4.3:��T)IC�����uNJ��{���(��q�s���q֑0��"�D����C�s�����c����j��O�gwy��I�����V<8� SCխQ���`T�i�D�������d���-���x��`�4l�D$�ͮ��a��	����o��귴��������"��L-��ٕ̀��f��1a����8D"�w�����d�l�m��K��,��<
/*��fJg�����k����;oQ��o�ơ�!��D��A��,)VK��NF ��2�t�1�ӵ���/�;O��Cׇ�D���|pJ�����`AW�|���o�䄬�֤�v��̼�<�U>��z�4�֝�4�"�����4��p�/f���xi��4L2�g+/�_v=�,F�e�엧ۻ��'�ٛjS�L�>�(2�Z�`�#rsg��=����u]�����+��0%�[E�E�Eǧ�Mc�mEzGq�I�5.�/R*�ItgU��j����@�;�F%<WJ�|<���Â.rXH$?.�c}�����'$�s-���~}�y�jv�Sv:⦙X��5�omY�TW)4�b�?"n���>=#q���P�(������ǭ�}��E��Juk�S*�J�[\vO5>Eî8.�M�K)e����=Q�E6�L��w�g��|ԁ�{��Ðj7g�a�3F���w^݆&k4�{S�EuJ"и��r����Đt	KKX ��@�xV�5�;��dZ�p"�`���G%���F�vi]�� ������z-\�ws�,��(CѲ�ӽ���{;�e�i���5K�ɵ)�O��RO��Rr�7O�*[E�6z�	�/A�<�-�q�0nuU�w�Yk;��F���Ac@L �F䖢�TDy��&�zŧ'H%�J���a��d�kC8K��ys^e��0�`|_���C�H��K.{�4�c9V���E�H֒�r�z	~�����V=e��;�m"H��(��tꏚd�k��s�dS&i�=�)?4>�^5�x��v�Hkaĝ��.�&˯��[���f	��I������>ܑ:�Q{r�l��I��U�A.�,�/��c�
��c�~Hϫ��b�A�}B�d��1����k�J,L��ts�77��LRk~H���I����0�H�v����Z��w��>����u߫z��'룽|5B%���ԍd��� �@���,Ÿ�w�[�wו�u�L밣k/��iz̈B��ã}�����s�ޟFe�f��yڒoM�C��mYۄ�����Ɋ9g��ojƮuo6���)��2�!�-�{���u��ƜP�qB� �����ﲛ�Dd*�2D���gmDK��o��
�{�(�O��p"��N{���K9��Ϟ�w���N�/nK�o��%O�z�y����/j��=�_��	���tڅ������$���@E{�=W��u��\�_ǟz��H�ڡӵ9:�C5Flms�ΐ�>��E��;����?���+�7k�>u�W?�'�!'�S�l"2<TU���P3T��<�Ѵ�;3�~�; �� ��g/��ٕh\g(>��02�Ƣ�c��{)m]��W���ňu�.�?8���'W�Х
S	m]��^�.��3W�}q_/�|�9��Y�|�����j`�i%�	қ���	�{s�ߒ4-_�RN.�t�	�d[BV��@�+V���W�w/��a����0�C\϶�ۃM�{�ۺT�\�b���mi�����r�t��|Vo�s�}�^�~���$O�B)��O��#�{ K*Ɲ������3l���]��/�n}N��uc�qmn��I��ǽ�1pKJ�D��8Z�!�n�/)���F����_i0*��i�3W�+�����:��	G���RD��j� ����|��[
5pXG�z��r�{���e�����>"z�4����/:��L��H%�J^}1J\�ݕ{�{�H�'���cM5/mHL�b4-'�n;���{J	{kU�OX�nj��W���{��:2��i;U��p�:f��6k�g�2��oXW���a��xV=�_�#O���11�;ё�]X�}h����0��Jj������1a`^+�ݑ�Y��9G� �������Q��Ȱ�G4�ƣh!�\n�iS{/r.�z�+"ʇ3{��ܚU�� _ B�/�������S��F�g>�7����3v^�a�|�@�O�Z��a���DԷ1�+~��5f.�����1>@��	04[�q`e-�s��D�,�gX1$j&Y����w������őշ�>ڼ��F()5��/��$�<�ϴF�yO�+f���#2,�G��i�*�d��l�,n�C4> ��n��'[K�<6f�f|1���.$F�W�Zkg*����L���4���φ�i@Z�9��\�9�S�:n�.W�)�0Aa'r)N�JY�**sWfVf��Wn���j62�[�r���L �EuH�Wt�S�D
�-{�j|�¢����n�o=�mL��L��b�nG��Kc"b&BehȔ��G(]����%�4�{E����8;�7W>�R�h[HN$�T�HOex��Q͠?!)���NR�~p�bK>H��2bzQ�ͬ�𬬗�y�v�VZ|�R��(��y0O=� ��5�脀u���#+uN�m��};\��>��)� ��¼��)������e�&��T�^�i������*3yίR�n���`̭�	�5�I�`[�� le(ӰEi}�6m�mŶҬ���{6�)��;.��ќN�	�â�6b3�,5z2�a�"�a�p�HJ�I,ی�Phܭ(0�S����Z��
�&�na�q�ۘ��n7 Rƪi�֞�+��xDa��ӥ��.�حt��U(���ʼ��72��6�M��!7<���%R�/R�͹��y[��n^+�V�;JU��_ŧ���\��P�ܜK��7<G������K^i���ss�q}+ano��a�`Z���vJ�/K#��XWC��8�-(%�^�2��ga]t�押����~���^a��p�+ji�\��N����{	A/t��9�}���܄�Ñb��b�]��y�Q��S�F@ �j
�P8���0͸�/zm��T��x�}|e�6�	�@1�^-���ך�S�g&{`��������a1���/�^K<�~���cgY�Ш�˛�Mh��q��\��x�0�ps	��7�Q�ū�b��a3�A�e��6��8���T��u�G���>�~�L��ɶ��$=qhON�{���:"��D��Aif�Fd��x7ɇ�jv{��h�~�=�9	ٛ�~#w�R8o?$}Y�M�QI���-&�����G���ٕ,�ZZG���uuS��t^t�5(�7a�jm�j	���/�����x�z��>�G����{�ޯW���������m���F�=�c���K��{�9���y��	`���վҷ�zd)Ћ)�.'r]N��]���O8��{�Eaݾ������)��ױ��,�Y.x��ˣ^��8GŨ%膂Tiz���;-�TPi�@V�Ɍ��M��`U���"����{�=y{��#�t�w��%*�.�������ZG���;n{B�v^�?����O�r���zM!r@#�og��Jb��3#�����NE�S^ohZǐ�x��g�U�������l�x&^�s�Hۥ�YW�;��u,#����Bm���a�bG� �#��S�v�ؓ�9'=�q�x��(����͞z�\���xn�����gC���b]ܕ�]x�.P\�$zzb�OP�n�.��*�g����P��~l���$g0�{��އ�[�M�x�X=�c��YR�4r�r�g��y���-�P��^;# ��.9\Q!�M�19Z}g�%0�����ő!��2jK������2uW��t��(1{�t�}y���V�{�ڔr��x��^�14(܃��f��7��a��f%^Q�	�T�"����}����ܿCp�z������h?��*bj�p~�π�`�W<�b6cU�����X�8�"�����9:�1�\�9��^��P��Y9�^�S0��
�$��+���뽸�&vm>��.��2m�$�&`jK!NȥF�������S�g�Z�絍>5�|~���k�f��9|�r��ON|���n�KXF'���:��ケJZ����.��V���b�:#�	����T�*�Z�4�uۅ���Y�E=��(���l�7��w�5�|ؾ����,��n�$�I��趪�ꬬ3��hV=��������P��c|�|� qY�x��$�`���E#�܉�;���/���w��`��}P��g�7��?�g��aU?��5L���QB�� �9ҳF�2�=�⻱/e
���V~�y��s��Rx��촛e\c}�ݝ����״i�9-�9r���0�3͞�}��Q���c���5��c��#�f�}Nxv@�E����a�_�,���{�~���ϴ�f/1$m��:��^�7��1ZL��-+���}�)���ӷ&�ڄ�3�l�^��CڀvS����&4�L	�̞��f��c��q���K,~�������a��c��U�yN�!�4���g�F��j���cb[^����@��{��5���Y�7QK����=��H�\�@gײ-�=�=����%5xy*��v�t��o"�5>�� ���ꐟ_�w��]uV�H�+�!����Rg���V
tsc�gRB��Q:���ʋ�	]b�0�$$�`c.�b�Y�`�i�8ǣ�ܸ�^���Y=�yI���3On��[q�P�^Y�%�9���x�o3r����'���f"��ӈ��b��ӣ4TAUUMU2EL�m�I�d�jfmj 5���5��j����""�"48�N&*����&�&J(��6ƪ�b(���5A��MU51D%��CV�6�4$U�Q:��;b
����AT��QEE�on ��(�j"{b��*
"*��
bb�(� ��*�*�"�����Ҙ���(����`(b���mMU%4Z��TTTE�LQT�:0QT45ES1EI��D�L�P�P�A53@D���PT[b"&�� ���(��b*��"h�ӈ�����J��(?6(����ڂ���TSTˬT�f~f��N�z�(�L���zΪx�����fG/x{����d�6:5!��X�w �6E������R��-=�tW߱}t9bm��Mo���~��ڢ[P���D\zz�S{%~ڊ�q�4��O�P7�[����6�ߛ�F>�"@�wjE)��M+I��.>����ǼV�#FJ���Q�2��[٧�+����+�zTK�3L�)M]�;�=���{w�<2@Q%ٲ��`�����X�puzwon�f�>3]yr�]���p�[X�����vO5>E���� �6M�����*�:��W�C��Z�L�ӆ(,�`�s�;�&��|s���%ph��%쾾G�mZiC�����w�V7Od4#�,/�p|va�9q�yW�����]0�^�,������ي�zu݁�lVvҾ�ڵL��h�a��>��r9���-z���ʵ��;(�߬�6{*��;w��ݻ�[��>ݨ�5���eǆ1�B�PG��}?lȩ�R`K&i�B��T�U?0}]l����~
��y�Z"<3��ܙ:�UL�SD?0���;k���n}�m]#��F�+ִ{/t�����u���5�=����3��$/�l����(}�iLx>>7��|�٣�d�MIUc*�i�>B�̝y��=X}��{�T|�v��$�?>B8g[ͨ���gr)�&��=�t�v��=f����-U�ݓ��{.͘vψ����z�'�N��8�-���4շ�iC,���іN�l�^�&���NV��j��v.l�߁�I��r���
�h�E�|�GQ���us[&y�kف*��ᲈY~[y�g�r�h�Jk�u��ýC6Bאw��f��,Ťq�����xF*��[$(NE���1qy��[��B˕�|J|�W��	1��_&8S���e
��}pHޘ8�5;��>��O]�«p���笮��-m\�sͼ�.��
�����["�Us����8�(��.D�&��r����|�Z��T��7<�&q�Cf�2��l��������>c���K6%��D��1��{������p/�c ��@�I�r�om�Qp��3Z
�"K���Y���j����9�S�/j����\��2װLRux�
V%RaM^]�7w�.]nF���ER��Z�qfݝ����_����i���}})���Й'b��(�T���t���*��.�E�Fn�j�ʸP�h)�� �4âL9�n]�4����{�Rd��&������SEӝӏ�{pF�9Ϟ�����F4Ð����; K*Ɲ�������=5��c��C?�-%�j���=������L���\�_t���2I�E�f�N��.�s�Y�����g�o>���C����h�u-���&5��M�6�^Q|��O� �/,��[�����-��K�v�Ɂ80�"�`SY�ȣ��m�֪��Q�Ј��ϳHޒ���k����%�ʽ�e��pH�/#OD��KJ�*<�T>k��rٍ��|������y�L��t��L?��F��Z�\��iIc\������ݚ7!��66�`��&��ہ7wBg�֚^��ލF��$���X������3ή~�"<��2���W�Xt#��nYs�O�ކ�����>��}/S�!B𨘷[ak�%����hF6�}����7�6"��z�[f��A�B<��:8e�sjY��u�u*7D��o�f�wnK�$h���� ]�4=��P 0�lI���M�-�� ��^��t�w(��]�V�OkVu:�LsіvN�m�^�.ҴE���l���P�<�F~Q�P��"��z�e3��vE�m�D�UUV6�~��Yo
ԂC�Pi�e�A�ʺ&���fq���B,��̔�Ulp,�vj�*J���וf˞ֶg��k� TkH̎Aᯜ�~*�!C��K��ۦ���u�,���X�P5[5U�w�>h5��E���3lΠv���(_��A�z�Уa*:��zq�@�ۮ���������Fu��-b�O��+#ǹOC����,��Ze����7f#�z����~B���5K��]w=���<��۸	���ɏ��v��|�j�2Y2tC(��w�LX��AZ��F.oI��T売���sV嶡��-�c^��Zn�Ъ���t�����,MdE�Q�}���Q?K?�p����!�s��d��U-�[E&�JG2�F�'�nE<k�c��3�����;����et��SI���L�b�r�sw�mψi�O5?!)���Nj��9��x�r���*��C��=�����+���V���4|{���<9F�c�o����/3Ք6�����i����\���y�K"���$�0����]D'���3d�&��.Ct�j�Va��"���͍Ql�.�ț�y�حt��]!��&�.SJ�N���6��� ����M���jY����7��{B��&e!a�J��P�⮗�r-?2NX�ҡ��8��j�)\^�x����5�y�fx�����B�׶��I�xI�`Z��N��¨����z�+���sn�V�!_N�Vy�G6�8u�0>�6(�8s^�����Z�	�-l�BU�(ҵ�	ɭڛ�Mvo���2��9���/c��6h��{?x?B8�����W�6���I�j��!cኙ�W��z���}:���=p�tņv$���`}���~U��-��=��^X=%�h�͑FaM)�}93�<�։��/	4�Ä��=;1MӪ�6���촡V,�a܃��ub�y�� �]��gy>zΐ���B��^��g����U�
�Ml�
e��ޔgY�a�KBF��>��i*y��p���/c~�����-*�V_�v�����|��/^$@;D�y��5�m���Ļ�&���r��E�UVs^wO+�^5�,h9�����L$�Y琅{�Ӵ��-�>W{t�Nl�5WB�Nm��;�q��򜞅Jb=B|��i��	�)H�L��<釽�7��Cz%(-VEr[�r�{�s)���[[�8\Ҩxdyg����'-�������@^��V����a����S��v�6�Jt'3>����8V�7���VbS�R�E�JW�_E���ߛ�I��G�����Wx�_�J�*h��I�a@�f=[ռ��|(8"X[�$>��A�6褫j���d�N�l�V�ϱ�8��Y���ebR��q�fuQ\�U$��$z�8�'2���z��'b�d��^o8��9�F	%s��Jt�ħV�E2�$�5���j�.�ξ��=�y�G]P��5�-!��~f�B	�f�L�˲���]����$��'+t�U�XsQ1���o9�l�[9D���=qِ���G0�G�Ђ�Bc�n�p)��kdڟI�O�H%��O����u�zq�;���x���70i�/w"���EhzzO�=��T�w��_�y;�C��{���yrXI�p] �5?^~b <z����>T&[�LpYv�E<[�����z�+/���z+dI��5�������r�5h�;�57�|M�3_��͘�TV�!�Dz���x�KOb�#6$��ξY�km�ݽ���R��k��c�-��`��X8���ձ��#�l�w=�vOǦD�dS�Q��B�]�
eWW��E����ʛ)���Lz#�����`����'#ആ<�@h�E�Mvd*�N�Xp�Q9{��:�_�K�_[�L:�^5�:7�V�-8�a�#�EKU1:���p��1�Ƿ|���r��۵׶���g*��v�pl'3L( �b����c���?����r��&�-܇���ǆ�ϭ�0O�f�pőJ���Y溝��e�:s䮒m�Kf��ǳv�W��/�i���{��������+�О|H왳�:��[޶�D�<�O��0�j,C/i2�#��kT��)>����y��)S��U23�`�2��4�����N5��~'�p�:b�T �t[9���e{��K�
b�X}�WjHK'qnǔx�+9�k�:��m��� �����FeI�z1���/P�=q���ϳ����YS(��x|&*����aA%v�ݓ/'�����@�ڼ>���{���'����J���8.6�ccb�آ��\�AaN>���F5���g%d�����r�L..�G��D�\4��~���^�LnJ��2cT,�֭��Qqn�Yv0B��ǒM��Pfb&f/'m�[H$�bW��\J��� ��M^Ʌ���2��b���i�ԥJ^qM�;'�T[�!K[Ր�2�OjM�����	�
�]I���]��E��~f��&P��%9HȤ}*��@�Y��w`�2\�J��#�c��&�^��(�v(8�rm÷�ޗn�Je�`&*z�5��P�Ku�^!v�;����|�ZdF�8+4^�~�<5@�,��ӵ�F
'^�����:�-ۜ�-O}{}����c��H��ꔴ�P���;>uX����K�jrDwޚ��~�U��(YD��al��fd��`%9���mC		�ݚ�W�!�cn0u'nt������m�K|�wk�o|�Ĭ^��`Ĝqd
K���U��a r�Xt� ������a�з{5�ީp�����rܺ�p���BՅ��_���{J	{kU�OX�e����57kz[,
T����g(����,�hgQa�x�T
n���#�T��έ��2{p�f��Ig�\��)�W@�I��	���7������z������Ľ;.Ɛ���;��}�*z�3�+��+@;�3'Wҁ���83���������ݗ�{�#h]�F��+L��
��0�	�T��W:C4C@�����Y�vJ���#X*P�܁	 �]��Ԭ�l�r)\�8���i��@��:��Y��A�����g��,^���;�׹2�o��ʞQ[<a�EyG׎R��1@j9Y�Qg�z��<P���W\�|V�s�1��aU�{!�(4r2��e����f`1���,ѻ�7���&��,�O�_+�^��Omxcs ���}s�W!
�#^i��t���垂㥃�wΙ�Ӕ��wk�Z������Ǳ5ԯ*���r����aT-]
6�p�7�8���YX���y���h�?/(�r66r�����[#�0�ͼ �/!2�F�'Nv�e_�)]N�{<X~t[C�<J���fҨ��tc�1�m�_����oO3r��SֵQE���9m�c��}:�ٙ��y�eE�R�`��R+|#[ӓmb�O�׾xԂ֫��X����(x9Ν�I�C��k1��en�����ٜN��K"�<�ʀIRaA� �qQ.��O�� �5��L:�..�M�
A�r2�7�@nZ�D�z�'y�E�fu���g����/HO����r�K3�靵�w�xjf����pX��B�����Q�].q�?7%��P����R����\�m$+����yFq��S¦�v����oI��	VY��qwr�Q�&+Ѻ_���畜���G���M��?Jw�BV��O淧s�o'���:LZ�2�1!㪣�q�S��%��dUK�ĝ�����D^T�Ln�*r6Q��$��^"�8�T6��oY}2����֨B5�f$�2�l_uȣ�Uz���sV�ϵ�r:xY�=��K��� �CB�=�/� ��SM��=E���!*�0��y���OE�����L�a{]=��g�&S���a� ��k	�{��ƅ�'-H�أ݊25౫��'��Z�{:�o�L� ��jx�3+
03�����<h�^E�*=]~�霃���o<@��N'JmyḂm��I~��#�_IP=�D[�u�v3�w�r�	������ͺ[��qp�M�/����h9��X��}���H�D���b�)���˂�OQ%PS9%m�^�����>2��)��Qx�s��᭻�Y�}}%�W��P�%�8�ꓵb��m�ܚ+��om��B�@��j�������ϊ�p��z��ȊmIK6ل�I�&a�R";1���X^�9W����5���3;�[E�E�.==^�N-�%cj+ҡ�=��8U�����Vu���j���ģ4��w�ȟk�S�)�����@��.�\�	~�?�xH�9A)�z�m؇mZ#����g=9;v�/���*"7�d�䰓K����{|z�%��7%I��K�\pU���:_^}u��Ӳ�:�����|Pc޵`������r�]��7�q�1��	�E[Q#,��F�2�)�ۀ�l�1��'BPЁ����N+�K��E�+3L�JUƩ��gL���RP<��v��W��Wi��^�����uٮ���!��C�Jt�ħW��)� ����;2y�>Eã��2���+ܾ��[Ob��#���a)f5�(2���2����4�㘤�`�+��0��$8l����k��Z}�^�Z�Z��||�zF\i�*�t3�jz�1i���'o�8*�=�׽&�o�z�xy�@~�l��X��9�xeoBw�i�r�k�蚪ng�4��;��k��zJ;��c8�1	�;(���-�[��fD��/�"v��Nfג	���OGM�/�L���浦M�XW>�U,�[�ͳ��-!�-�B5VڐWG뙪����oS/��\��еaԦY���;�&�i/��:�;t�0h7���7�UN3��s[O��bv�mK'��q�^;Io�	�i� �b���Z��18�����}�%� ��2����ˍ�D�����jF�W�A��pȍ�s�,Ÿ ���z��>�o������{���w����z�^�>P��	g�v9�Ll\e�v�+�J��?�h��� �!���)0��ay~w-�}�Hn]L����y��ű���n���;n�jS��Gn����.�}i�|~a/N���pjuR�KMZ]�	y�[�g�b��g����uJ��@�{x�pA���m�f��ڷ�xD����f{ ��8=}+��|ڋ$=
��>�eK��yjm��E4*�I!$�� ����Y˱��겱܅s ��<�v��>^9�i�i]&�Z�<�2}����Zx69�F{�w�T�57m�D��|G��W=tbǼ';��nM�yԆF��Y%��m��˸u�̢���ae��u��Q3�yI�5�'8�}hw �c�0n�P��;�{}KN3���Y">;�z�Z��"�-�O[�l\��gtTc����咜r�cy�EJM��j��᫉֒�0���T�p�V�����V� �s�{���9Ǣ��Z��%'\! �a?jIg��B�fa�U<X�²�}�ې�:��A��x/d#"��^�v�`Ks�L-j��:�J�1q�St��"ؠ����q�љJ����^Pe}�޸�Ȓ0e�Lg��a�-�g�Y����^���<�'�o]3Ѱ�v��q��q�C�+T����e�gv{�6��+4P����[Stc&�H��
�1ZS��uk"�u��޼�ϯ�󆸷}�Y�M�;�7*w@��j�L��A�`���j/u����!S�rߐ��0O5��\�f�w;��	�hg�y�=�sW��g$�h�^��Lm#���&&�0����n��w����R�/����~X�Y�N�{��}�H�c��
"N��b?�޽ݻ�";7q�.9݀��gi�8�y;�F���pm�q���d=Ҕi�/&3��t#sU�b�x�9��үӲ�x�:��FAw�_g���ak�
"'&C7��Z���F�vm��ƨ3���ɵ5h�u��aۜ��*��D��p�������糖��,áK6v�瑆rMc��6y��%"�w>W�wԉ�`gfK����Q��h�e�N�b�s�f]N����	��D}�-si������Q�N�V]��J��V������8/��ݱ3w=�O�/��J��^˛k�E��:��8,]���A���)�
dJ�e]жUE�^��ׯc���)zZ��K�p�����M���c�{/���듄^�<�f�7�ю%\����NDs��˱x�[a�*�>��p-�0u/�2*ʞ�;�z:3��K��}�[h��+{IG=}��Y��g�@�O�=z!�%J�SU��fR��ɹ���2r�0�C"�@�FM��ܴ��!�f�hA�vCZ!2`�8[�S[�b�F�V�F<*��~�/����u�T�{�=��	p)8��:n{X�ɸ�~��vny�qʶ����y�V杻�l�g{��w�}�-%�&p��@a�0��b ��y��axsf��j���T�?��AWlU��UATQ����4�2v����Q@D�S������Gˍf�������B���*����J"
��	I����J(*���������b�8��u��J+��TT�Q�(�i�&���Ji�(�ST�Ph�4EIT!c����Q�j��8��ƨ���)���PT��[n�UM��QMF�T]�T�RE@UMlizlc�7X:J'���"j��0AE��SӦ���j����gcMSDE�AQUU�IA5WZ*���l1��&�)����"&�
�hf����
��EE;%�
b�*&
�b��
j����,�����������=|ʮ�!�����7����`Y�LŹW�lH�&RYn^[U��1�iJBfp��8*�xp��{�Ï�Om�XF @ѡ"ަ��RhB@�W�j�;k�%U�k*=�Q�E�Z�~�T`��7���Y�^�����7(V��ٕ4�;���T޹8�����#TR~��)X�xF0���E����ļ�h��k:"j�5m���x�����梮Pd�[>��2�lQ\�T�C�]|,>�Q����7}������&zF���mN�}d0�	��	eA#X�^1���2���\l�P��[!t��هy�5�`��v�j��5N�j�L.zЃ-{&):�dJ���vN6̌��O��!q��#j�D> ��*��~�i��o.��8�:�������zA.�j[5��ˣ-�SיЭ�oVK�Q��$ȶ�]8ތ�gZ��H8v��j�6����Gu*L���{D��fx]��E���f��:绤r[Ӟ?)j�22СÃ����xj���{�p��G���޻����0n�N�
ڌ�5�{ˇ�ӣ�ʾ��튥)iZ�
~��*ȋ��n��l�W<}����ɗ1�"q���z��o,���	I>�w!�L&�/춭B
�?���=~:"�`��V�yz�,���j�:N{����������sS;#���������ޤ��mh����nf�2&%Cʍ�3�n�;��n�
��Y�r(�����#�ދA�u^E�;
7�Fb8���̾���i�#@3�<�Ѫ�n��Zt$ŝ�TA��E�����]ÞU�B���='h^X1']�����<ʬ+�a�6��B���UI��:ڻ]�%���0�����Z��uH���"�xV�y��J	{k
��eκd�2��d-��3��r�zO
TǎAA�+�=(��f[^΢Ú�G\ ������wg\獗�㳊�2����)/�%O��p�H�W��!'��'��?�o)m\�=�����vl�q>�=�.��c�w�^u]��c����iD[�5�և{���y���3����<+��U�w�qcv.�fE����Ԡ@d9v�l�tM�1����	�l��+^�A�Ê����ݾ�̭����2B��U�B�#^i��ۦ�:b��Tԉ�EOT�7\H�RθG0�pr\L]����TcWXʩkj��!s�tWB��%G\<\���Ͼ��toNҦT�C��G64�`�L�q�8�+کnj���l�	��u��V�S�3d{!��Km�Cu���`}Uź	M�bU|1Q�B<�D1�#���������|����"S8+�V�np���4Ν̅�u�Tm�������|�*�;��o��A����%apa=�F�<BaDؒ���Wn���;a���He��*�*W*{pw.1��s�E�>��b�cX���#Xs�B�X�%uW�!;���l�x�[N���6?�ȟ^u{���>��U<��#Z|��V !G�pWc��[iuz���Ҥ��խ�V|8 {+��)�1,���L�%I�vF�~�*Ldu̟vr�c��C�s>�T�5JƑ*�}E�{"���J.�7E2������NZ��m|K}J�31e�������YBm	����У`�(qG���i��(��t(~i�i��#
e�۪���؋���t��#��M�^�#[�mM'W&q�l&�V��F^���s['��l͇�]V��6��nfep�]X��-�<�j��\�������O�_��a�|�g7�5Z�,�ᛛ=��j�^���U䁮�[ ��@Ax-�����'-]�>��q�'�=��6���ߜ�,Z燪������3<Ǯ�z�H0�Á��4_����;}��Σ��k�*���f�v�������/@� �I3~��-�Vk�	v4*%�&� _?d�s����{*�5�6Jq?K޹'�h9ݜ`탺	@� <M;I}��G�ә�<m��W��{B$���IVL��Vrx�EB�����!�}gw?�lD����j�b�V���_]�f<�O���c�4~�w|=�`� �Օw�sX�U�����m�s���
�a��w����6-���m��S��,;F�g��=�{����s����2҆Bi�'���g7�kN�f����UHB%�N�.�Ye׫�V�z�l���C�\_���?�,5_����~2�v��IS3;[*ާhYJF,Vr7E^C�<�<B!��`Z����@�OX�Χ�JO�*\��ߏ�U?�>}G��ʄ&/���*L|�� ^o�O��bܗ��|xW8���Dg�ݩ�4���D��PW02eCf��K�z��N�������J�jЂq@��E�$f�X��U{�ڳ#U��I�^Go��-u���n������h �vm�0�t�4����'z��&I��Jo9��[*IRkk�!�A��0��Њ�����m���kAG��ki����"�)r��gIwMm$��b��E&�~�f��Y�{]K�q�W��؆��z�+&:#���W��A�ˁR6����zU��
S39��xe�3���29�-/#kǦ�Ot���c�<0>k�PE�Q�uT��KH���Y��Y}��1z��y��BoB�纤���in�!�2]�?�߯���^��A�Y_��10FG�����f�BG'��3�8�[@\Ň^���V_^����We|��-�ot�a� Ɔ,Z�{p��mʭ9g+O[j�p�@���X�:_-~�`�}�78�Nl&.����x��Iw
��U�ޣ���OE�����	X�OnE7 ��Ã��{�ٽ���4��HJ�Lj�k��)8��<^�G��A78�"X�A_x,#=ޝj_���mM��5�c�C��箨R��b��S@�e�a�U3�<�a�>��C�sD�C��3P��,��G1i�M���P���q��vRpl'��	y�ף��&�&���g{VS����5��!3��V�c*Bd�oP~s�dh&$�9�n����lb���z�	ۙ{Lu��/P��^߲%��b�=1�ܧ�(N6�(}�}9�E�M�R���ލ���Q��d��r0���TsM���f|;�T�a|�d�����W�^U>���]Ѽ���M���o����W(5y#!�׳l�tgO�.�`��7�z�f⸝>e�wW�����������PS�X�'�j��5����'�/n�N�z��>܇@�n��S���c��|�
Fȡ\LO�yڱM�j�L)�w�2ε�L�ѡJ�*�
k����:�=Q�d��&�x��m׶���E����3w鄝� o�[�mn~�Ƚ�9�Nw���{4�j"��m�bzF�Pdp���h�͉է@1(�b^�H��1#�|ȟ���Nۋni��J��\ʠ�%��=�#�"���=n﵋<����=��#ϙ�<�ҝ�f�����֤����'�C�gH����!o@��wDX.m�-��.0�koA�A�y�'�B���ཟ���E�.��7!���v���ސu=��][�*5�q~�絍k�`*����36OnGy�/Q5)�t�G~k�l�xjx�TG?��.0a�cLbܼNӴ��)옦�.���=�#�LfX�m8S�@�`*$19z*<���Y<��a��]ȫ]�Hr\��	�ʅ#B��¨�ye��{���^���G�9iR7�^����m����=3���	������P,���zs\]�U���U�]k	����-�?e�7���6�T�ץ�q���2:`Ü�Xڑ��g�D�Q��<�{��Bn���/��&�j�ekm8<�_`�j�{wE�
�f�i���FL3,�{\�5�P/�@6��1�p`��y�p�{��u}��r\�J:�+�>�P� �aq<�2ײ=�l�E�ʴe��z����3��>��ԢK�0�q���'D[��Ϲ��7
$�>����]��/?�1��ާa2-�wdwE�ǡ؃�-�^)Ẁ����G�8U�Rǔ.���] sy�(��ƿO55�ec�7�1s^���"�ʜ�s���g���_��������ݫ��>Қ�ӯ%��	��f.��ά�{�\.�_����Q��~�8��q�,�wg�k�'�o �ױw�'�6E��;��M�J��n�h'ی������*?>�~u�=�hNk�nd��?r�_'�Ց�鰴����nc�RJȹ�1��<p��C��|"�h����^Ե�.R=�W��c�f�z�u�؋>e��w�>*��e��-f(*�I,���&Q����%cj����	��4�e
D[uD܍\�x����1�b#�s76�h��r��g3��XD�¹yA��EN��sO���lfIs��y*��ګL�	�xp#'C$/Rٺ��Gnr��n�P"�S�0Q�0����)%���5��v�/cz��D=F*����t���E-���A�ݱ�y𗝁�% n�͉�Ss� <ضO���8���f�#��R�W��/{��d���w��N�7y�2(��SŷҰ09~"
�F�u@�p<@��B�b|f0_Yz��=!u�ҳ�����0^�^�ާzvgUGJ�G��fPL�7f��4F���YwL�1�)D6�:XH�����I�Nq�W�h�����.-F���N����O73���4���e{f��!��h�<�_�8R��j�nJY�H�$��t��É�;0*$͛�
3�uaG6ަ�;'��P����4_�2~���$MM*p8	�y)�}�#��^q��E�vhy-52okf��:�/�LO><��\_[Ϲ���)c��jn����hi^��p���;�rM�}�v#ź3�Î7k!�!�I�~�M��s����*�b���~����%S���#9�^�{����]͆��mQ��#����ؔ�M�s��w�a] ?���m��PI��>��%��s��Y����3��'lk�*d���!v�	�������9>���Ov�e�v�#�%^H�Nm��e}-@���}>��ֳ�5L�n��y�ϗTGL)�$-%���'�4�EAT6N����F�Va��ͽ���\��	�7e����)\#3�r�[�ݝ۞�zb1ca��y�<����+�q�G��Kn�J�n��*�IH��ż�tA�;3�!��=�CcaW�w,�ތ#���.��x�?e�SI��C�w�x��/�fBq"�|�oB�M��&EML ��Z���V2+3n��+$��S���E6=�,l+�՗��~�&A����/���	b�l�����x��}�_s�j�/2~�ʼ�#06ަIy�H��n�(]Z ?M�D��O��-��GGTn�ai�y�O�������=��'~^���^����^�YA��d�~���9���	�G�cr��򺞄�.���m
�L��%+����GwL�����Ĳy.���h �mp͆��EUɛ��:�^nQ�#&Ir�hrn������5�JP�i�z�w=0b�q���d�:f���J#)8H����I�]�/Ֆ�eP3��C�8��3Z�;
귗C\�g>�6��8 �	�Գ�gM���/�����y�]�Z�sM��[����O�N|��A�����~����ȘU��v;��V�n�������A�9q,pI��s>�g@�X���W����£�V*I�A�{8������T�}%�Dq-���]�}���-7���JSe&�GmMݳ[����o��m��Y�b^#
�s��Yt���=[x�Ԟ�3t1�� �Q��`^N������f`L�oN�e��-7�#v w����A��%���5Z)�'����6o�7|<u?pP<���w��j{��m^�~�s��H���HL��B��;}|GO���!.��Z���x�jIΪQ��=g�4�P���W�oC��r[|A�EI��Ɠ���m�f�B��ٳ���i�h!d`�܈֍d�B��(���f�ܑ�/w:�5��.^��:i�i�\��t�m��Z�CiH�+���P�:��岉�xuc�}��wv��DW�ݙE��؂�a�4����N��٬�����>��&��"��ҥ"gʹ��ݮ�j=��gj`����y6�i�j�h�\�G����Ig>��c��G=&���f�u���ӓ�t �	�B[�4k�WU]�ZzK�N�R=ﲢ����������i� T��D�d:[�6d��fAκ�\���*w]CӯJTo6�F��L��`�q��6=}C+�f�]�
�������w����5qjن͛6l٣F�4l�qlݍ�� �Qm����O�cдth��+���RS^���>^+��_{�cv��y��=��c_h��A�)�4�ڻ�g��;�H��$>�';[�|�Eyw��C7jj�����*�HDM^'My�K��C�����p�͂����ش�d�/j�%~�I�)��S��:�oU��׼v�'����G6*�G
��<DD����3d8�[���ܳ���.�����;5z7ឧ�BV�J���^�ý�?Ose�R#|��A ���M�Z��f�w�X���Z|.�l������E��v���lv���9û�������6Vc�C�D]M�ߧ��M�l���Q�=���w�Vi~��@|nV�'�s�B�K{�Z_�?*�<��l��{k�׮�m~�4p>�)��uL)y��/}�Z��W5����uA>��'����܅Wj���0�d�[�Ve��������1��vp=�7S>�:r�F"4i0�[W���y�l�pq���P�)�
�-�p����������!>{n~���Jz	E*�ǉ@�i�f�.oM���3g!ķ&���}3�Y䯼5�Z�ᨸ��\�{%����}��1�\�Y0[�g���&�h#L�<��/�y��B�s}�JV�s;�]�l��]�Ws�V�N�|2�c�钯f]�Z�*�!��>Q)���{z�	7�gV�=ψLȺe\j��rruJ�4U�o��w��_�o=��ġ��
��Gweb٣�6v�|U!�0��4�G���>�u{}w�� Fs�~px���f
�p����1P��ka݉��FӨ��y5�����w������������ǀ�N����)�_�F�����/4�#�����F�Ӟ �b�湿/9�K���\Zk�o޼�tUw���ɸNVl��'��5�f2�q�hP�*�����qL�Ov��P������d�V��~��u}�7،*a�΍7�o�L��v��́f�pN����J��S&�I�A�Ղ Li�����I(m�6�[*���'�2d6�^��,�\�Ӗ�^綀�S�����~�5|�4��mQg���-d�L��vV
V�3�9�i�um����`�a����{�x�w������|K�|�s�u}�J���g�g;�=�����N�/�J�V���i����ةx�-���ɸW�󝛑��y���Qg�}�Y�Z��95�e�0�RΚ�ꖁr�Q�{g�_Ev��Ru��e�m��p�2j4�'0��a޺ge� Ƽ�h}Gދڋ>���ڽ[��%���0�T(��AS��S�w �1#l�$��ua�%Z&���9agi�aD��������3����g���y�����i��5�n�n�ާI|@�e�8�@3�Ař*�ͫ��8�F����X:o"p�w��no��s�����������������G�y�&	���(i(����b���M6�QVɢ#l|�DTM-EI]�3UD��%0L���H�
���h��h
j�B'gh�H]k���Q]:��Z���ibhd��j�(M8&��kI����#lmZ��#F$��Hh�蠶t�S���i����h��i
��
"못�b�*�E:tiѭ�Hi�3��&��EZ�6ƃ��ZkA�tj���)��F�if�F��A�A�EU1SAm��U�ƍQ�
��%���j��iД���S���kj�uc�A@V;t�mKF�-�F��(�l�LU�l�J�h�ZcMhL@�hth�QQT������>��'����bu�W\0�ƷFŃB���|*��i*c4��0m|�Q5�'p`L��r�R����W&Rӄ)��k$���l,K�!�=�S=�/��j=	�q��WYܞ򳼜��CE��s���fq����O��g�d������F>�!�e�F׮c�mE�C�8=N�6~MH��H$H$�Lv	�����g���ܿI�OT%�z���NY"B��!D��c�k����8�)�F!��}�E��˃���^��W��4k����|��z2?IX��Va&gG}�J���W���=�����@�w&�cd
ȩQ]c
	?=\D������Gwuouf��SsNge����s��X����ux#f�0�0�/[����C���9���'��|pOtkT��`] `V����Ȅ�n|ȅ'�u�T$���[>͚��x�W��H�Sy��y��В��}M����*|L�V���z��;L8^���Ҧ$��b�Ņ+q��f;�bbp#���w�i,��v}�aKk��s�'{���x޵PY�d�����P�@Mkn�(��kL�D���,3Bb�QE\6
ܕ�C
�����������zYʎ�O{�U��6�	����fRkk9��q��$�eţvy$e��*�^Y����?fd���w6�`�m��/C34�q�f�A�N�6�'���ֆ�X��j3͋d�ndJ��J��kl0��G����xE����G;<-%x�9xb��Gv�dzz$�&�O�0q��S��6y��^���l���[I�/����Vp	S^T��s��di�q��8����1�3�����<6V@%z�R�alã�c��lGu���!��� �Ψ��R�!�{�fm��a׭5L�X��͙�dqԓ>���>n��cP�/�|6�ve^n�h�u�����<;�f��Y|ĉ� �YG<��U7]�o36�(J[��;RB ,�s�W�N{�57��Q���の��������(���R6)�䵎y'T�GGw�������vt�>Л��d�9l�o-]-�h�Ҳj���D`Pf�9�Ρ"/oB^�?{��˻�0U0ՈlJ�}��vN�q� ����]����kXȒkN 4�T'J����s6�����.S���jN9���yKfp�F��;C]
�\k�{b[��$bX��7����{��� �Q�r��	��(�$q�6��2�j�#]V�8 ��̫��j���h\�jAf�PS�PI�Z{2E�o�б!�Ca^liw~�;�k�a�|$fV��[-�D�)]���U�/������ݾ;�FM'{Am��Ƙ2�~��p�|�[R5/�z�*���yR�CdVbPm�on4�ˁ�NgS�"���e6��l�?:��e�.�׭�
�G7��{1��. r0�᷹�F�YO�`�F&������V-3A*\�̶s�l,��/㞏9P��M=�\��E}{G�#�s{z8�l��2Yؓi���V1f�"G��r�F|�~��a�,��p���̋����ؚ��rS�{�4i@5C${i�L\m�U���A�³���-@#�{D�ξ�U"�W�n�N�����4�}�k4��$jktL��㾇��ʃ�mm'����4��$�t�u�����e��$VBp�9<���������Z��teOjI� ��(Uj6F�m�rm�/T����qv��#Y.�Ol���fϔ��.M@*��(D��Y�C#ށT#|��������_���x����6�Cz+�`*�x�����Et�F�<��V�*�"�v~��3N��94k#������9�צ�p�Ñ%��>L`d3�b0n0��JEE�Zz�/��W�I����ϻyd�2�y�<$D{O4{ܶ��s h�^J9�\�NU��ή��yꠗ�����-":�|GHR�\/eg+w�ū�x���_�7k��suD�h��窕Bf�VLT��m�Xn �Pu#�PZ�[��m5�Ou���^��ffF����ZgC�=bL0�k�GCq�YD�x5��;�G��֌ݾ�m鴻�L��"<�Ե����f�>���~�l �}�֍^�[��l5���s�s���H�rMW�-nS���@$��	��L���f�㻘�j8�&�(�G|�Mҥ#^#ks�t�w�# �g�b��v�n��|��(��;�3SX\��X;n$ܙ�u���mN-qF��`ӱF@ی� -�m)Uݝ��Dg���z��\v�����8�ׯ��"Ο<	�=Gg�/C�i�+��GNw
��Gg�v��x<�NOw����Z��q�z�I�;��i���(s;~�q�o�U|Z=�%Q��Ecu�.��������z���Wv�i���ǂޟ9��hJ0&�d����\��wI��NN�L�0l���Ȳ�&݂O����y����ó�,n����oمg��[�Jr޺\I	HV�,�lٮ�]�]#'�gI����+����j]R�*��/�����[ґ�=#lu7G��4uy���q��W����踻�Ҹ&u&��z'�>���@.x��&zOfA�p,���j����RZ��գ�Gv|�9�}]�!�(������C'1�Tbs�y�\��'���
l'.�	q	7�#�l �fg֧꧜P�n��ʹԻ���GD-���o(����H<��,����\r�ҷvrf������]i�*�S�O�j���=ܚ���Y>Q\}��=@�0Ƃ���l<	������b}~�E��:m������<�n|����8�B�\�ʔ�oVg,F����.ɷx�;wyֈ͘��1S2�&}�h��RZ5YX0��TUe^�M��K�0�����|FyP�{�)�e�p�5L����#M�Q�� Xf6�F^�z��ՓjE�9�d&�A��tg����K|����$�y�������1��eW�+�-���S9�U��p<pF��1�.���2tr8�Q˼�.��zQ<�zU^}��m2�m��̥��i�q�wOM���ρY�������Gt���%Kd�$�~�h�i�x�Owj�ڸx�Q�8\�+v8.�S�����b4�[t���7�C+�7W�����פ-�HSb==Y���y�������W*�z���Z�����Ā�&�)�N�v����,���>����"�WU��^�3��%%���������,���1�ϡ=�Ncɫ�<�W*܉�y��7�zx���94��-�;�uj��s��g�|�t7��W�r��gC��L�tT�q�B����d7Ô)�_�������{�n郀ĈȋqC��淕aU����aE���=�BH�zz�Z�A�b�f����;Z���z$65��r���ɸ��^��v�oz_B�����L�S��ZT��Bw�n�|��������u���@lX�����i��`n��>XR�L�sm�g{�O�[%9��t�3���ujFHY7��}؏W���ò{�W0�tKښ΍S��'�A�k�*0�Y�l�U�����Ĉ�u�W�W���y�oT&{�1��{^�s���u���ث}_^�_����AF�����_ξ�h�5�K��Ee)2�\C[8L���B�7���i�7��X.��x��5i*	i���{{��`�mY�5�M�.ͬ���C�yTf�.c$r!m��Pg����&朋!�Y/n$.~9����eD���W~���Ƭu���D�4��P����h�S�ݼX-��>�^_Qp�N�p�]��#A�����C4���/'��Uhgq�~��3�/�[%�kh�[�z��Y�{
.���Ndr��;o��wq<��'�}��_z`���?���w��4���0��c��ܛ�*�4�2m�E�Į`:�XޝH^{=f^0&?���}�q�V�9��#sn�c
Am�����Yy(y��༚.��"ʋs��e��[��R���M.�}���t��T/��b�NP�Z��eYJ�%�v��'����og�lO�����n_�~�y>�3B��f��0���������g�kbM�f�K�F�h.�؉�5��W�1�C
���eF?D�Q�gfw�9Qbjpw%>W��@҃T2"9�z/i�:���ʆ�c�=�/M*rWP/�)�XȮ��ާb�2�=��ݝ����Xu3��p]/؍,� �!p�Xr졋���+�Kr���!�õ���=!�;h��`NΫ�\�I�6��qi�grY�Eo��5�oYڶ�1���9[ :(�S��}��� ��q��G��Dr�k[ ����5��q�����>Q׵р�&k���Z�����6���P[�7`p	#��⤄���[$3	k���cw^�qI�Q�����檌��=��k���EI�g��GnD�S�^�;�0!�k.mD�큉辮w.�c{��o#�R*�8���pj� @\x6��{LgRۄŘ@�fs��R��[�QM���E���ٴci��8�EԱk�q�w`����s�T�G��e�w����i:`칃=w��?�h~KpRu�0g���o(���z8X�늧Z7 -��X��Gj�U�3�ۇx�W��U̞�x�g@�yA0��{o�7��[a޶4\G�&0�4�7�{�>2���i"��-t�r�O�2$[�����T��׈��љ{��iZ�cv	6ܑV�*R$l�s����M{gn����)�u�qmJ�|Z:�и�Ԥ-/��͕��E���[�t]�|�Pd��t(�9��]b��_%=㋡\��.�m�gzw��8Me��[�fۤC[<��;!�oV̕^�fNu�{�rjʎ�S���[h�_V���U� �,#-����a��t��{`����#k�eUϾ�4��oS����'����z��Sv�ts9���Y�ɭ��t2s��`�\�q���Y�	���9R�������F�y���?���ָ�kٓhҨ�bܵ)�%���ˉ�Sx���0i�����	���y�:Q'e�R��3��%�vg��7����Q���^���}��nI�_f��f���x�pUR��A��
^%�4yN*�ι4fF�m�R�d����z���O=��=Y!)�l�<w���A�&;�.�)T�W鍟>քsN̩��B9�^rُ��x�N]���n=��7>Y�s�q�FP��@�z�7�F��o���/$Y���f���nG�	5�tp�j�Rg��$w>��Kp��!�իg;�,(|�X&`ȭ�;Q�ou�-�U��K����r�SJ�]M������gB�PF����F�S������{���>=��w$�FUz��۹��2*���R2����'M���[q��s�|�q�<봞I�S���e����j~�k�3`F�oo�^u�+\�Ʉc����Ǻ\�TɟJVi��MS�S�Uq��̘/�k�)�-����
�ѻ<�2��t�٩ٰF���P�<���*��t���M��B|�H�[;�&�q>�t�<��^>>^�w�{���w����z�^�W���e�#e��=tƹ�QP# �H�W�L탦�?I��wK������0F�
� f5�c�����K7	UH�͒Y�D3��C����1��6�%R�Mɋ5C��[T��I��1�^�hԷ��f��gw�E(w�>��>��;��i��剉�	.��(���gakj3\�7.��6���wWd�5�4����e�
8�Sg��"�U�� �s[.����M�u���۹�3rzs�1���HSl�� �賻�>��t��=��rb�ay�;�={`L�"��ɏB|�L�f�v3uM�s�v��cө;�"��<��?PwFK�^÷9`=�^Y�y)����8�	��
1[9�\���eXu<��w.ܣ�4��ຨГ�w�C��б��3��٤�-V��՗�����3}-]p}d��{���rj�nm06>��'�����G
�a�o�����=��y.3�����a��H�w;/�k/����Y����p<e�����g�^�V!�n+T����S�k�Oi�z�vv�Yބ��j'v�A"����MŻf.4A#���sX�c�"X.m���e��̡��j��{�[̈́7ƽ��]X<4���7͆@ĔSp�}����}���K�7B�*wH{3���bC�s/mͱ3Q�m���/^
,��l��H$�0��8�t!+�#����L}�N�׷A�e�$vݜܵr%cf
"�yU�*ཌྷ�#�Ʌ�4+����3G�iDiSNv2�W��|:cY�"/ns�=?ý� �O4�(��j_����j:�Byj���C�j�py�U1��V�e<mZT"η�}(�.d�^[OG�ԃ��f,�F� q��4=�od΅�a�9�[uD�i��d\*��7�Si����B�w��id,U���/n���B*Q�kbm�mC�4�
�x(�l�5�b0
���vcfݝ&�ܯ�&k	)x�d3��hJ[YQ&U)��$��܅���N{7^��s�Z�&�]���=���$�{n�]�7!/ʾ�W��.~:v�"����ͳ˰5���-z�@��J���jT!w��Օ�IXf�j�9�3雤����a��φ�|� ��#�K�O��N����~�nq�싂�-ӗ��������or�ؼT�J��1�F6�M�+.rZ��ŧ}�]�O�>9q
�Bf;�����ܗu�Ό�?
:t7�l�
����k��Ї�{�2�r�� w�y !���^]%M�"��˖��3vctf�v�!Q`��ᾪ���rm��9�3��� Կ��ٽ�o~n4�)�
u���1�EӒ�B�(f�P�xZd����E 
2��eS�F+�"�Ȭ{�N�n�㰻��{��,�T����z{���A�y=���98L /S.�LQs�mވz��`�ح/gY��D��2��M
��TL<�M�q@:�ڴH���`�WQQ#?,��$�"ˈ�Ғ'��!+n��u|�Zŏ��������&��S�(�mf���E��b1���5A@S�v�q�ZKv)�4[RQ�*ѐ�Pj�X���`�kTRPQ�֓g�*��S�j�)��o�Qv�*�[�qm����ѡ��N �#Zj��)5��m�,Th-�+Z�kZ*��hj�T��gA���8�Z֗��1
+������ѻ����k4TI�t�`��h4X����M-��ѫcΫM(ӪشIX�F*�C�I����`մ�%QEh�����m�tPi��PiѬ|��t�ت��X؍�l�jf���~I��6hn�D�F�F�����M�6,i���6���⛭%mQlUkX��kA��%JMGq�R�3��[�j���|��j��:*N��˽�ٽ.բ)P�!2�u�e{�{���pz�}cC�go{����)l�<�N��xnO�Έ��i���=ۮ��g�w ��d~gQ(�J��>Fc��<º���7}� ]g��W[�w�݌�\�{���ZH����q�{�h6�|i��3�����)LE3�'��ܮ�$�&�ɐ�ԫ�-��54?L���� o��=ȍ��sw�kUS� ��T�dn^���><�4'�,O�/Y�k"2Mv�RᜎL�3�BM�r�����I~��p�g�������{�R�����8��Ό�xV_[�f���:�w�K�]j��c��\�0����W�>h�`�#b����:������)�����8o/n����ϭ�C�_�BQMY;cb�ϲYŎ�Av%=S�ɰ8~����2�	�a}v|&T�6r���\�I4��6m,�e-0��j`��xݾ��<� ��w3�V��WQ�#S�7˰:�eZ�$�Tf_�ם\)ᨘ,���`�q;�Ns`te�6�����`�l�b0�г�*��p�<���{dV9J�_Φ��o���R��G'9o&en퐭�݀�Le�:��ÁkFɗu	�0��DNmJ&��e-���O��+qjCu�����\۾�GSB��zuM�^�n�Q0�A��|r�a������SY�BWF���
�q8NEl"��,�HmH��c\�ෙ�
�,�c�?oo��nӸ���F!Z���e6��;�ZC,ϱ��7�/SJ{�p�	�}�+;���Cf<{m.���������[�yyKOt<`�\Z�*hK��[9�}۞ϡ�G�pT�1�:�xwqi1�t9��"K�G`�3#�lI��Ƭ$L��Av%�9WM����m���E�S�p��r�R6gUz8ѯ97]�r�ޚ4�`�1�/-�^Jm��y���r$��~opĆ��(�M��}ziPrWP�<���qU����8�v��/C�~[ī�0��.��F��{�d�1��p:�*���Tka��Q�o����L��bz��0i_X�WN���D�{���R�H�Ut����iV��o���{���{:��s��_�cE�nԝ�m���պ�&��l��O�/�FU���Ώ�n��L\�f桕`ʯ��^�#>�E������9?n���z�j}��z�]V��ᛈx�^�Q�U��#�d��F��m^U��j7(<6���ǽ��!e���=�-��1�e��>�c�d�O�K.˕��]��|�F}qVz���>��w�	(�<���wE�b����>���nZ̎���P�tz�#E�#�_�
�'�.�21�7/r�-����J�I�ł�P�y��Ƿ�Q��\�U���ٸ�1������V.�޶;R����gӂa��ڴr���x4w)��z:��^�����j*�̞�x��8@�r.�	髳x��G^�d-��2����R+�rMS�t�ݸ�isP�/��:�372�w���[!��m�"��a0H����r�-,�Z+zݲr�G�ډc�F�h:�7}��U�h뒫ǥq�R�-/��,p�~DƼvpi-}���nciǼ�)A�]~z���<�]�t����(�;g�_䷏�����m�<ħ7|�F�7�z�3WRsn���	^�0�5US4�Zf�+O&��7�����AU���:{Q%�$��8�����<��$�ފ�3�/�<�@������cc!�{VЌ��������k��n6{e���z�̔��t4�x�QS�3MqNOO��vo�,��eE}�͆�]9=�kDtJ�&�csY����m��������V�9����Vq�~�n��q���F��=ڬ���QQ۽����6m�qu#���+�vr)��[�\��%���O s8����զ롃s�k .�k�m� tq�cX*(�r�<k/5f��N��#�YG���M�67��f[n��$��r5��(-��s֞��5��=�4�����Y�=E8��&l�譋n�L���<�6�$,1���B�Z�b�CP&�垑�jf;6u�U�K�������n���̵چ$ң!.��=�6�>Y5���u%]��I-�6��e^�<�yVL@�Aew$�]܃�s�SNg����,��|�i{M.2�䩿N�����ɩ���G�{l����s?��W�u@�k�k�A��0�9|�Dqc�nL���\�X�����<����Wgx�CO�T�{ �<&G�1���lI�Ԅ��������m���9ǇI+܏��~�^��_g�;�k%����Sl�����e���8^=|�|܂�B��U	*�>�ĿC�u>J��s�x\�5u����%p�T�#mx�&i+c	-�z�b��ԇy��L����$�{-f�B�`���Kv����}6�?y@S@�w��7�
G{_��و7N����}!�l0�An'ѫe�ヌW���W�!a�j�uڋ���I"V�Ԍ���
�N�� �E*�8_3��֞:;��w{�<��䳇�dƣ5�T�R��b��7�cE�{o��ّ��OQ��_ս�b]�(*vd1���o�����:�"�a8ݦ�iy��5�i�k׽J�al���<�h��{<�����;!�����x����8���`>ٜ��|/K��#�_����z/�=p_]��ѣ,��	h����k��Gt`G�>h�����5���-\���|-(��`]d�6Y׺ v���,7tr&�zV�q������V�=�O`�����$"f���y����������FYR.�W&F�"H�zh��&�dM�G���u&�K\�8r.^�/�R;�E�ɵ{��q����q�i�Zo�u
��h�0s�����!sO7`�cb��!�hWC�KP�P�<9��s=�YZ��;o(���y�wyqTF��h��;�[%��B�z
�5&����wuv�!�{�eD����HO!��J�9%o��Y��'�w)܆��8��GX�\�q0ݡZ�a��}
��l���B�%"���q�T�B���y��ڵ{�5���.�! F�z�+��j�7d6�U}��ٞ���#l�7nDW�`�]�oL��r5[��g
b*�#q�@ˑ�XD��o� %z�߾z64�s�$�-���N�ߠp��h�[���<Ѷ7yfli�e�������I^��N��6�.b��C��N��|�گss�A��0���hh�r]r 2�Yϒ;eOsu�p-.�X<o�d1f�X�[>�����kb|m#)wv�`���D��D�{�KN2«�n�<"hC��ma�u1=�a��������RL�f�c'd�Tja�%��t�E��3��Y���F	r����Q���ǰ�7���z.t��oWe�z/tښ�x��k�IsB��f��z�	�ݒ$\j��кb� �?Jܘ����P�&?�<gfw��'\��;�U��oE���M��Jқ2�z�_)!�9dǏ��AN�	��^�T:�&��� b�p܅�~�~��+�qlJ�_/�s�}�dy�̅7=�@��z�F�|Oy�Ux"�&:A�2:��Ch摁L?8���w�Wj�D�(�s���y9|5�J��sܣ{�Y��^�\���d�i��
��y(y�;���C�v�������|���z{3<��"��w_[MK���$R��&�j�.�#����U ��F�0�(�Wn��笾�@�����@������=W������2ʛ2��;��f�`ü���'�*%��g+�`;�h�2l3Lqv����4����h�`8L{	{=&��u�t���8@�yA}~�<C�}����iB��*�[�jݨ�;X�6gk�f�����C�JڞmYdam����[���*�qS[qٖ7����v�`������&=�������HM�٭w���'35ML[�,�	dֹ5�,��6���Ci��6��tݘ��5�2��p��F�EK�4�K庞̜̠��uϼƖl��|OpN����p�����H�g��(t-H�m��ډ��@��DP��o�gi��a�&!$Hѕ�#�F�̪�- u�TJ�5%�g�Kc)a!�2����8�ն�k'd0�%�G$?��q���~���zq�o�p�x1!�kV��}�ޏ.�̅�m�F G[Yٹw�__�CV�oM�&󛒵�`����,�SJ�d���`�l����o?��E3cne�4i�̬9�F�S�.�d�j��R�]�oKu�sR��0ۊup�/��f�oe��A�u�7~�(�ԍ'��eϒ;�gݧP�Q,B��#N�o]?H�,F�P��H*E�d{mq&�I1�c�4;��d������+�+^��a�HG��"7��7ve��p��z�lB|�*�)��m���Z������Ʉ����I�ܞ���ܭH�����k׺M�˳Q��Շ�щ�kޑ���~�4���Ǚ�wzgq���<_g\��G�w�l��O��]��~Ħ{l����%���1}�L�<�t{�E�<��7�
��>��@�v��Q���qp\q�,ח����!f�S헫��f�����) s�YN���7�ϻ�#�>\�8����q'�w�'A�7m��隚V�O@��Zݥ�V&���{���w��X#��\�F�ݽH���iiMC}�z��M{& �!^Hυ���ȩ�/+v�������m<�}eN1�Ö7��|�r ��,�ÒzJCɌ���|S�| ��s{��͝����3	@�b#o���I�C�o)��W�\�u�Q�ɺ�]9�gTy�"�8+�eO�4{���vc�͊�]@x,o��HY�#��|ŷ�>A�nV���U;�cEMVDʘ�VEy��Ҩ����#��W@��ӆ0ͳ�XB��o�%��Έ}���(>�ߝ��5�wt���8�f�����5��Ԋ?�-*��B���㣸�����+vvkȊLu�>tw�v�)��lٞ{���^��)�kƴ��H��'2�2N�q0脡��d���H���P��z��fD�͹zڨN� N�3hܤ*�_h'����=�S�%��V��/L��8����f����q=�a�@p��ڭ��Z��k��m �5*o�2-�莾3X�埣2I���"�<��a.�d��8��Ӳ7&��.���`�Q��St3tAs��Ȼ-��b�B��=��~���=#ȶټ��oK��yd���O�װ��ڵ�nS�\�;X��biT��0���Ĕ��w[�=6N�9��wkL���N�DO�4�v	:���'�W������L�]��hF�K��)7�5�Fu.��7x�T��E�%Xب��Ԏ�[�O;]�(�=�CU��*��\�I
�;I��$p��i��֩��7NN����{2]�8��"�̈�&��8����	AM(9��B{����) ӭa��@D��2���}���bݹ�cV�����ځQ��T�Ţ�ҍ}�z��k�l��%�U%����z��U���`Sw	f�pO����{=�^�/p�{���w����z�^�w��!�'Y�k��vQ�[*�QE*�_LѼ�NնRcoT�F;T�Ԅ 孙[�0	�U�%d�f��A�����'�S���*�7�rK��XK�޽�\��Hq��ᦺ�縮��݅/�6 Fe�:�t��/�����b��.�wq�n��1ՕL�����nZ��qe�s��o�xi>!�M{}���f9�j��f�U�,97�ܡ�JU��Z����-5y�^��]干!�_C�V1an�.jמ�9�}[2��wǇ�z�3�L� X�,��}^�;2Ǩ�N�Ӝ��D��(?>���/KS��Jjc��w7��ت�-�xJ_��5oI��/-GHV�^�vW�l�}�/5��$���cߝIy��MF�ȑ[6���׋b,;�j��\�v���ث���|xN�=���3��	'�<Pr���W[����V�W�b{/���h��YYY��vC��v��[�F�h�f���gw�90�׆�>{��v@!�xO1�_��6���j&v��k���s�z�r�(%�{�s��h�Ƈ��U/|���GN�酩��pa�ƪ�聺�l�#���!�>;Ea[���|�S9Ҿ�z���1o�1h���O��q���n+h�{{n0tSAèP�Wr�ͷ �Y�0'�2��j���y��w_
tv���N�p<w�m^Ё����w+~s�P�(�7��ϡPN���Ǒ�\�k��Y�}�����Vj�yP�~���[�m���x�r�[�5OUI�|��g��<ɉ�-�d#�{�z�5�2��^�0fT�pN���Ԯ�����P����L�s�M-MS�F�h�95����/���bf���{Y;�7^'�����u�ƌ�%�zu�Ri�<k܃��X\�����ֺ_��z�g��iO)I���|��_$�N�z@К��k�Ɛͥuj�OA��&	{���tP����')��ll���lȺ!��2i�xX����y�%E�ѧ��:������u����L��یk�20ˊ����UW���W.3+%����3-���}��yׅ%�Ʀ�P047��}!_o�W��׌�x���L�E&_'��s�vb�j����g�K]�㉴����$oa��a60nS�Ig����ᛷr���U��K�v�`6����B$d\UP�&jɥ�<�Q�j��ϵ�p�)��Jm挍S)b@�w2�%��
'�7���=��o�����y�L1�d��[�b~N�r��7N)�&�՟S%;��7k��UT��*�ؤ�SgMTl�yv��q�o�.���䞳�4���"�kG��׵s�{�kYST/p���J�(R��Ml
%aK�*�_���:UH��W	췒�����7�-�X	��]o����
���c�d�S=7���m���e�9A�lt�ʗ�y� �Gٺ��^�g�����������_D�=�E]�ӡ�t[P=�lSwpvԔUQ�E㻙���N�[mkUKl�����kZ�mV5mb�N�풵T���((���Gv�Ht]�h�kl֌DF�h�u�w`�ˣ���hv��ѭ:(4Q�h��࣬u�S��C����^�M#�t4����8����v�DA��8ۮ��h� ��5�mYvú��hZJ"��"�m�A%CGQh���"�l�����4��m�&�ݰ�u���E;��b�I��l4m�ѻSEFƃGU�lf�����λ�7l�A7X�j����M;j���;T�ն
-���4�MD8�m_6;kc5M%F�:��Dl���|��c-Tlf���d��l�$t����[��[:֮�Eu��"-�;�����"*����j('�����cY��j���`����'Ni3t)�p4e���ut�0�R�fJ��� �X���-Nv��������ɷ�-��6�E�g ,�'u���6���޴��������*I*��q�N��"�/]� ��Yu�;�&�;�.�O8^�54��ZM wJJ�r�A�L�yu�f>����ٺ@�w_*�;�4%� ���m�V�ͲT�wo���_�.�5�vXse�U`��	�F`̯}0j5uн�]�e��`?fGZؓi��w
8��3����;Y�r�9u����pF(;�:�;3��q�A����7w/@�%y�m]����İ�(UC$����=�/Nz�	���ʄ�!ݽM���y�~3��B����^�W��"�פ�����K'{�ͬ����U���K���<>w4��E�%�,w�i�Y綽r�W��,�~��Ē�㢌�1�^��n�K�d�5DO�Gtɇ}
 p��L���lf��!�wS���͟w��O%��1GWۤ�T�a��c��F=M��8ґ���L�si݉�Yoand�_h�⬋0� kWӺ�O���g��9n�מ>fs`u>���{+(U�
]���Z�-�쥷{��{pt�Y������7j���?w���x���;岛��Vn��V������8X�B�T�D�� ��Cl��+}��{eE�-�'���7�el�V�zY���UG<Sx���7�4|�oȯ����gL�L˟�G�t��ג8���Ohadб�0�R��׉E��� гx{���uHbB�%��hA�T@�������g@�=[3��F���)0�o��CWW�jH�J�(�rMS���26S-������Q�;c閜\/[ĊP��6ۄ
��t��$U��T�"u�q��]���֛��Ƀ��N�B��WH�6�xҿaMq� ��J���=�XVk	5�GY/��x�
�u!t�^�8� ��������?{^i�J=즗Cw	��[�=���6.g�Dkl0�a�["c��ud��k.n�m��O݈�[������,�R�w|o`t�|�Fo��~s+�>���Bu�[�D�^�[�Nb��QoZѿ��<���[-�<�p�_m��9�)v�w�&��
:m*��⃻���ELmڃ�����4�ia`����e�S�lQ�~Hw��-���gO5���
����o (�ɩ�/,`�]����G7 �T�]O퓄&	�Q�ETӊ��g�oR��T�ՔOu+�U�P�������D)ͮ�Ƃ6ς{��j=>�-�����r�3��u#���_;�;�f��-\�ob��l�gH���pa����>zZ� ����@�"A �<]dh��ֈ孔�|�(�vё�3�_E�
���w��2ٻ2��Y�b/ Rq6e�3��G�&���&߯���@�,��R6j�Y�i�pJ�d.���]:vt�_�=�d�:��ges���澍�������G.�t3�t�h=؇��裥-���<�]m"�ԋ�s��m4UL4�nb�T�<�����ae>�1g*Ɉ�i;��%�eP�o�z�56�3��b�_v�W����	.g �q�7!�5a����R�]^'�ӳ�_3��K|$ ��EO^H���!(�8��3�)&�y�J�9E1�4FS~`�Εs�@쾫õ�d2���}�'��	'W����3���xH��kv��� ���/\v3sّ5$mUS��"��jJW���ʚ���Fl5q�0B��X7��xfb�uf�cE���x�{�+����4'���-��k�
��~��a����5>�#��:�8��-��J'{y�����,I�-:��Rv�W��o�A�nj�E��@`�%����x���+�oyy"H\��������sD��&��n�]p�!�tz�>���9TJ1*�ē�mv���g�OE�*���f۱�}���z�\F���/�F�ܖ�H���ʎ���)�:�Ot���ER}��q���dnM�R.�}χ+}0��L����i0I}mE���{k<�[ȕiʇ=��g�#�$*����kЦ�����T1�x1׋�{&|�vw>�h���Y��wFa�Y�͗|�"(�����q/�2���6���縑 �n�'_�ۂD=wE^Ծ�9klo&7���+Ӝ��tC���U�ȶVR��Ns��8��wr���<2�̻��Ub��D4G'ySڲ����T휋�f�96�k��>�z �G^���+Yl�|��o�ݶ�K�h)ܛ%�R�y:(E�� �c~U�l-��ط�o��9P���#���˶�EΈ&��j�pM\�Z*Í�[���<��[p�eϾC��U�3?Gw����R�v�i*�D��3���'�L���Mn.���k���c�y��|!Y4.c$j!m�Y�K{3�$�5�m�)tǷ̑y^>gA\z�uȃ��V�rD�=UL�6�N�}�&:��Z��#)ьn�S��pu9�*�d����9��K�h>�>c��t�U$��~������x]�5����f�V���n�mA�JoKGt��.%�L�˨�[1���\�kk�pZ�^Ƕb[E���#�ǆ��U_&�{7�|�'ئ3���8��L0�$�Gh�n�\�X���dx����DGl�7���|�}ֶ$H�-��mY�4⫎�=��2�x��k�+|z�q�lΪ�;�ݹ�ߢ�.��a�馹�i��<�M#S�f���<Fp�`#�8�dt�W�̇_oa�����i��װ��C�kh���r|g{�ޣ�pe��:C�,���x�/Fc3�ͦ�[�P�I�n�@���E{2�	��p��&�J1U�ꑦv�{R�(��	}�7���.Y�l�X�-�2�����7�m[�u�l�{�K��(������oޥ����q�z����;��`B3[�:.��i����]V��J@�vN#�_eR �%Ǳ<�x2�{.����_�OX];�+@�`����z�W1�f�d�'���3�Ih:(��˺����e�fmf�SGvs�q�DyQ�dlU�c�0� ��R�O�C��{�΋4��TD�a�9�Y{L}+/�L[Ί	�
0��K��x^]�G2a9����.��o�6�3�F���dj�RW������.���5��yU�\ձ�QUcq��޾����"���T�H�I�TK���!�/�v��R����<<p�ڵy�o�Kr(�dQ�4 ���^=�}Cƭ�U�{�|����@�s����~p���{��Q�0� ��䚠�ksg0�3�3�N����E�uCȸHɂ���}ӻ	b���t��yGJQ��g��B�V�VN��j�����Ai����&���j���Y�~�U�l�J��߀J�q��93k���� 6���k!a�G.�9ٖ��5�0��$3X�hJt�	��%��Nݧ=�5�AL�{�Ǘ�O��C�$`�	}��:n����r����~="gKU:���J=�$lnUd�\V`�Lbv�����w��L//yuW�|z�XX�1YO�d��3Ƀ����幽�/������¹E-��R���L���S7��W�՗��M����Z��QN����|j�@W���y7��������"c���پ\5#^�F��_!��d$tg*L�ʷ�_V׏wR����������0Lv3e�=���������p�=p�w.R4���Ѣ����ac��Y���G×�������,��#!�+��!)���Ę1�nx��<��zM`J�}�1�/���g@��0��ɼ���y�@O8�m�r�dx޽�vu�i��t�8�؝ח�>/�0��<��ؙ����u��ˣ��/%���=q�S���״����=��z�W�;��`4[D��zp�ĝ���`lV�<��B��v���u�o_m#�-5v��=�{B�V��<�0�J*����h����1����{�G}�4��1{}�
��1���V0H�2�e4��ɒ��I>�܂>�7���5�M����N�x�e������wHF�܎]�1��TR�l��74�N/qA��iTb��q0�h����aĨd��B�䑴eP��&v�z�yAaX/�硄�����l��nM���XE��nAI��.�ؽx��4tl�xs`߅����[/6j����[co�`�JYY������~���c���I*���z��n��L�nOv**�d�r˴�ӘcL[i���g��ia�R����ŶS�m+�j7X�����.	"�bK�?L^�@vl�������Q�i!r~F,v��M:�S��1Y`�����a��X��}ݪ�@%W�4���+�8 �I����{w�h�԰>�g3��L����Qҥ���r[^	S����M��o`h�H4���9��?��_t>����#roz�x����M\�٢u��(�T✔���Z�	���nWX�_*ER�����z����s�� ~	^W^�>k�����h�G�w�E���\�i0̼��e���<P�]�"%,�PHH�ҡ�^�0�7J��x��`���%՗RWj6�����KQ��kzX�/P�����1�ȕp�R�=�Hq�z@�x0@����y�_�~Q�,������7�H��Cؚ�U5��{���z)��vc��R�y���;�`�W���N?��A��~�u���+��n)�v�A��3��tq^�=x�.�ފϖ��]y
�"ײ���*�i�\\��|�U7Y�d\Ի���1��TM	���ع�+��e,�I��}�T��U*����궛��l�.�+ɣ�	k�uD�1�7�W�w�V�����!���Z����{�P�'�4�E�
��u����7����^�ٸ��z���䒔k�T!����吪�-`�x59��|���3;k��	�Z�L��epԴ�A~aD�T��n��u�J��9��(�O˺�M�s��e��9)�H��В��ƛd�<��(g��[6Df���k��{�6��R�P��yMg��{��,>�����;�soA� ԕ���C̘�`šT����8�F5������ ᯭ�W��$m���YY���-;8���L�̌�}v��J��}�����(dM�LTd	PL��7;x��U�6��Ro�:��q�\:_���*��D�D��	�z��Fqq���il/P�4��Qź[���������Q�kb�*H�jj,�j��M�v�l�*�3�X���e�ǐ͆�q؍O�{m�"LW�r6�4{]0o[+��?.��a����=f�o@
-S��]G*5�Z�aM�^�k�����u/�7�h��w�B%/���U��e�(���"��k�����o�kx�=CL_0����]9�s�-���[������=����� v#�6��3�u\��J��t���"w\0k���l"b�]=��+�S\��'���T��V���̲��|�8�x6�.R��Qg�sԣ�%=��ל,B���ѡ3WT���>n�œŦ�ݍ��	^��d�C�nL�נИK�H��7,�I۳�?�z�JH� e܊�"���I
܅Q;�DT���#��������(�2,��̫0,��"�+�L0,���(� L�2���ʳ �2�³̣2,ʰ��3"�0,��"̣2,ʳL2���"�0,�3
̫2�2�ʳ̋0,ȳ�0,02�ȳ̣2,ȳ�+2,� (�2,���0,ȳ�L+2,��� L2�ȳ"�+2L2,���*̣20,ʳ"���}�'��	�f� �`Y�fE�VdY�`Y�f� �`Y�f�Vd���0,³(�0,��"�0,�3̋2�ȳ̃0,���(̡2,ȳ�0��3*�0,ȳ0,�3̋2�ʳ"�0,ȳ+0��"�2��3̋2��`s
L#0��3�3"�#0�3�0��3*0��2"ʈ(�L2�� * L2 Ȁ��r�ΕU̠2 � *�0 Ȫ� 2���` 	� & �UY� & �UY�U�UY�U���V` 	�U� eUf  �@f�`Y�`Y�fE�eY�fE�e�{=<�0,���2,�3*�0,��� �0,�f�F`Y����~/�� b  aUb ��K�F�a�������H=�.P����H���J�Ǖ.���xOU���� y�����uQPV�H @~]C�(t'_�?�؇� U�ψc��й!e�/�L��"V`K>!�l��2��� Ȁ!H��"�D !$"!)(K�@�(���(@�0�� �
J�² 
�*ª����*� �� �� ª�*����I��3��A�x�nO0 Q�


 ��%��n�A�6����q҂ *�8�8eB}��c�N�t� ��0AC��CbiA lP�L�7lL! U� *�!����] *����E j$�Ԓ9�Ix�!�0�H=�-I��d��̑p�V9�3Y�=Ԛ ��2,���y0/+�Aϼ���hu��!?���� *خD�>�OP ��
^+�T/���$��H*��I�و3��L6� U�E�a�$�8L�@\�WC$�+�T�3`$ZMTT�{�[i���$���PVI��N��� 9�` ��������{�>�/����#cF�m�FF�����H��l�BJ��Vm(�+ZV�V��Q��HR��5�
hdT�16��Am������m�ɪim��ϸ�ٛV����f�U[m��kJ�H1ZƴئR�lY��v뭃D�Z��g2�Hh�*�ժ�5�m)MPm2��ݝ��Q6�c��AU�M�f�H�-�4EUm5[J)��)f�H�ҕ4�Jm��mmjm�1�+[blѶ�ə)V���,��i$mm����b�mZ�o�  Z��o��[u��=k�S�L=G[u=z�4�k��U�m��s�����<��˹�볷ot6�L�z���޽�Zm��z����]�j�ם��;��Ov���2�f�{�uT�j[M�m��LԳM5|   s��/���bض
��}�(}
(P�4����B���
(y�C��B�ܟ[�oK�3{t�)k��{��N�WC�^�;�U�n�7{*��P�jU�v����*[{�{^+{z�]��z�ۦ�5�j�l��h)-�k4��   ���>�ݽ�=���]]�[i�{ȼ��뛖��{׬�׶n[��^�x{wK��������\��q뗺��n���{��r��ҩ���S�b�ӫm���wo-zoL��^[l�++c���U��X��   �yt�v�.�s;���O�T��\=nҷs�^�����-eU�w��٫۷[�n�]�f���n����3�N��+�.W:� ��EU*�)W5k(kmmM�ȶ��	�  7� �0h�z���
����h>���pgCS��((u��7[
����a�k]���Q@�Np��2�cVͶ�6�F�P�c[[+�   �hV���f�v��(s��4�7�9a��wr���pm��V�:���ܗP ��u�+mAe3+lҘ�x   ���+���]hV��A�9ݮ+�D:l�� ��[��`X����y@ �Ӏ��6��`�-L̦�cf���&�l3F�   ��
 ��{{��4�wҀ�۸��4 ;�ކ���sp ��W  4z�s����i�� n�`�����Kf��l����ݰ�֙��   ;��}P �&�@��G� {s� � sݖ� ��� :Ұ@������V�B�נ�^��[*+mV�J�ڬ�Fd{�  ���@ '�W �ӻ�8= ==t����, :�׷  eX z 7�N ���ǀ= ;{;�  �S�)J�hF�4Њ{F��)P  �L�JR�  )�CIJTM?R0	��M�JU@ eH�2��S�6jo�����e�_��M�w�5��r�ܮ�c�N�<�,��=4[�A1��_����x1������y���l�}��ll��6���6��m�������m��6<������3������?���}��� ��uM�� N^]�ڗ`��Z(6ӫk�*BF���MܤŅvf�en�:v4�r��&�økl`GY�aˣ��Ve[YPh-l֢������������`n�U�Y٧pi���f�M�&Gx�+-�kTSc�E2[ܺy��b�r�-ڀ���4�3���(��zs��� *�\8�� �Md��E���6��d�ô%h\ך�U�WB��g$�IQ�A;i�#nۧz�W� h���zZS�[m r-KcHP"t'�!��ՁK4��0G)��	% ��VUl?$J�Ke���:�� arX�30��4�`�s� A��-&c�Y����	��%J�/��-�sT�Q�%�Kjα��u�p�7��=7K,�,kӴ�/�Xn��vN��@��� 2�z�,�li�����z��� �3F�E��ʡY��X�k%<Ii��{WW��Km�k(�ˇn�T��b>�z�cUO>j�Ź��!-�![���/-���k/Q�f豆�b�����4V1Pk	�+vY�I�HӽlW�1'����"��l�6�t�X�g%��������1eATN�?�״[2��ԕ���Aʓ"p�V�5�w�)X��ڸ*�f��E*N�]�f��HK��&��IEoC̫�:�YCA&����ŒZ��/	j�*���6L:��1�+��i,�6��)<����/Om�R��mv���:-�r7�,�`;z�L1k�
�[1z�6�b�޹�)R��74�t�Y4r� �+͹l��st$��˦�� ��L ��h�r*0�.��v�vP���Z�+NeX����T�P�uR����1�ӄ��l�`�W�L�Kot�Ƥ��F���s4ۓ��Clǵwe'02!�l�^fj�߰�=cY���u��{�Lr���Y���B���cya�$W��f"�tZ�b#Yh�BAk�]�
�d��9��;0!@�H���A;�yRW�V��Xhw4U�Q!�GEU�R�D��lޫ��r
�	v����W��%\)H�� �V�o!°6�"�muo		Y��hz���M`�	�le��M0wj=û��F&��q�1GV��#�v�)��-Wvv�t6�ӡP^;y��f��t`x���CU�l�zt�j�O���$l�-4��Vu��	t,�6���w�<r�`v�l����*�]P��j�
��T��k�e�
b�"�*��M/�e�ڽe�X��c
n�m�4�����Y�V'�1�w�']&�����Hcr�2kV]6�l3[Z��k�b�yzp=b�i�hU�wd����j�'��c�ï��&F�e��ae)�/jB�!�JŴ[�7	Z�hD�pV
��K�0�ԭŚZ�ա�Q˃`i��A2�K&A���T7� ���j�2��u����ݢv�W�^�4��e,�����q�ܥ8�iiZ����ҭ� NV^�#�l;��/c��[3	Uj�����=��\W���΃C.ac�	�Y�D蜽�[�.2����PV���r��kuɱB�!t,���;
�:dX�Z�7Q���q�p轶��U��N��5[��ԪZ��Y��"����g)�0�� &��y6�U����A�xSjemf){�PR/�-V�1�.Q�]+N�4֫X�e�z1�.B�r�g�V��v�q�/>₱]x[
���k7"iR�t����&���gk.��63&���Bk,�X�q3I���J���f��6HU��W.���ư���H�=a�F���J���Y��Ȉf��[E�6�j�Ł0�Q�b���0�@�J��H��C���;oiMV �9��|�c��2��C�|�m��V�=g�o+sR�3M\�1S KEɄ,!/��F �m�Vv��B�Qr���ԃ"������,U�J��A��4<9�l6�,���#j]@2έW�EU�V�Bn�M��Y�Ֆ�ѐ
�n�YlZ�*��a��I�ק��ܠ�]՚���o��U�d����6��q\Q���v�|m�=܀�Yuc�f���� T���2�@W�F��]
�9`e�G��f���>x��V��EM�������*-j�QQ9�
e[T�H��1�]��8b�1�ܼ ��Z�[��٩cR�,R�8&]ؠ�6�s�_�i"�]���`�rHR��Hn�{�֪��y���[l*:�IAZ�`Iy.�g#���`���:RչQ�X���5�ڳx�Ӆ��ȮPCdn �R�!�Q��>��zֻ�;�Z��r]� BXe�֤`�����uF��x.����Se�v�w��I;yiJ*�X.�&m�V�ς%�y�:�;�+L!ei��m���e��p<v�H���!�����^������$�� �ح	e��2P�I��]��:��,F��-�Dք�(!vZ9�4����F�X�4ȳf��2��[]f^i����u��=Ot)w��Q kJ�5Z~9��R���Ш^����	�� C�m�ɑ �]C�F��wo`�R�}�������2[Y��a͆f�,�B�FjĨ,�P:�䛦d���sfB�Xv��g+F�4�j�`G�v�{��d���ń]9��;ȧ0/�n�7>Պ��W��nbq��ݢ�۩%[�ܴ�T�M=h�'3V�٬�2f�#�v)��В-#q�(47r� �N"�n�Z����z�yL5rJ��^�N�m����tڋ_����=)l;�[��c���J��RwX�ǹ*1�)�7Z)�6�6��3�I�զ��-�e�˺�H�%��Ttj�@XѪ�����7Z�r��i|�dk5}���x�L��ݶ�$g�� ���m-oe�06ŉM����*�;���	U�5kOu	��.,e륓
aպΗ��ƞ�۶�*+M�tEⰃM���Rь��nуm�����N�;�T-�h;"�Ow>�0�Y���bb�5��i�$Y�	0�;�E���P�X�%^��BX�m�p�R���c6B����n���7-cٹ�U�{&"wfS�ژ�ْ`x�����H�;�6�D�z��׻aMSl1p�I�[N��@@��ݜ�Ja�����&I��<����Tj�к%૖��0�,��zZ9J�n�^�ۢz�m��%n�0ֽq��M�i�m�̸�M!�#���*�� ���*i �xt�ߓT�<����=��ĉ	1wj�s5]M��o�&	�-[�Bm��ٚ��.ȚeQ��٘�����uf��҇6��%e�Wb@-��٩3N	��r�Ԉl@�1�4#����b�U���x�����$2ȶE,(��b�Qa�nT��a�K^Kj��*�&R�;��PЭP�9�􀐛�G�pr�ed�n5tCF��È�q,ߜ0u�̺�`�ZӶ/D
�^%[xƋ��e+�n�QhT4��ܻõx��B`����STt2f^hȞ�wk�(�� 2�-͗�77@0�+�$���z.������,Ӊ�:�����^]flg[�b*
�JU��k4�l=���PJ�ȯQ���4e`��f�or��n���щ4�u��O��"�9�<�#���7JX;b��ti&�[��K��U��,m;=�i���|rZ��ujQ���J�o�Q� �\� I��͸ݥ��m��Q��D�Y�Ҏ'�J;�+�wp��f�R�YG&��R�C�^���j���zY;��ou*kH�Vcb�7�wq
�yQ�˅���+k00������:�+�a�y�B��y5 �6+1R_Tӵs0�&�
y	��l׻u�i`�	�rT��,�Ӳ�m3OpQb�GXUƆ�V�_Π!��0lЄ,�e�S([�v�8�R9�{4��B�2����aU�vBb�1�n#+��͸�בJ�Z� OKNiG��i���b�~	��N((-�6��Qʌ@���Xk�j ����s#��f��H�[6J�lI�I�Ǐu���7Y�&dr�Vm��IR�@\S��hCl9��@�y)R��� �7e
���d��u{�e@P�u,4$l$�V�L:�YI#x��������v��$�N�iUݻW�F���G;X6h�x�[F�B��@ə�D�1�-�w�E����H
v�Y\�l�Cu#{��mVռǹQ*�4��X�-G`�srKª*�
�K�L�JF�S �"����r�M��F�k~j�!@@]���֓ݦ����{��H��Ě:��mkGq6���y�mR"��f��+�齶D��f*iE4��v�Ũ��f��P�Q[
*׎ܭ��&�:Y� ��
!֢�u���7���l��;�Փu�h�J�YT�d��G븬��rޢ�
a���W:���;��a"�6��j����U� ^ui�Q�ɂ��6V:hM���M2��ۦ��i��[xr�L��m�C;��D���p-v�V�N�PI��ڰ����@����&ѡZ�+��76��t�����A�Ӣ=Z�r6k!u����������۽�NÙe4)ʻIc����U�V��*r�ʘ5�@Dmf�HM�aX�e��f�rI��x�ĹT�JT�IT��lcp��s3eӢ!�KC��A������c��B��e*P]���vo)B��:V�w^�SV���u�^-Z���®KZ�
dY��ta�E
�su Y&���
5)�c1b�&H�j�V�m�fL|i��Fk��9�n:��ܵ��V��!�t�����1��m��B�F� J��5��kMY�ܸe&m�[V�
���"R{Yb�lR��(Ń�(��A�è=�;�#3T��꽰�D�"]��~ׁl��AV�AJu1�%���2�Y��D�ݬ4p�x��7Y˿��6�*�ܭ�פ��0�x��ZYx���ڽ&�7#�,���)���LAT���l�+bŕ�\�&@++"���42]-clZ7si�)�tk�	C���A2!B��SA�����j�����[�Q����U���.�&�kw{�FY���*�&fM+AF�ܥ7�� �4�m���vc:�+״(�vj2�J��b���,e9a�Ӧ��T�ZX$lƷ��X�kp��ŋ4��Kn�C���4��x-0\Vժ�V��\��[�7�Ԙ�R����μڔ\T�m�l�0�0طK.@��`��8�i�*3�yF�"��١��2А��-����ٶ��t�#��a����;�m�kZʚ�$��x���s-إ��7z��n��S�c12F�Ȫ�2dcoY��� ��T�]mc�&����c�E-7��r����}���s����J�Z�T�VT�M�u���˸�8�}zh��P�ӭD-Z��C_=���^�����Ɩ���:Z�8��u��V0 �*i��NU�2�C2�3�y�-I�����Աd���Ŭ�mcTh��#��5�1�Q�ê=��D]���ڄ�EcO61e�z�o�(ǔ�m
�A���X�2U˚@X���*V�E�xl8Յ����� ���7�h�5FV�)�y�@Ӽ��aCl�@�QxU���wHf}de�� l�̆cB�zF�16 �ˬg��޹��٬������������F/kq��K��V�kA�z�,c�F�T��Q��cp�/u�6�	hK�a�˽n�X�VhښoKM[ȭ�͕y$��l�:ٺo]=2\˻E�t�����ױ+X�ؽ"�SA����V-�r�g3b�+$GV �,JC����.���'u`m�Y�wpcZ��S�NXi1���¬�F�-1S�e|l���:�m��[�yM�;Wvq�n��6�Һc(26 KNlcb�[z	تU���ex��tƋ��J`��@2��cwUe\�y7Da���2�Tp��IT�Zj�(��f@���W74��]b��.:Ts�C�Vۮ�I���H���B<A�Sa��!��Wf������BK��n t=ʈ�Zi	��1�tjI�dIm��V�������[�;���>MҖw2��w�SNJ�Y5���v�EF�5���Ul4��\[�N�,Y׻��6�+��+t7TH[��V-�Zh��۶�ۥZN��=Z4�`����n /���H��j�r�Lܽ@���=l �n؎�vv���RI��*������\W{���Ro���ֶ��Ne�����u '�Mu]2�}�)́��k@v�^��m��y��Ś�e�W�Ċztػ�Hiɪ�2��,�j:Tl�±��x<�CZf��iE��,��M���62M9ɶy�s��� ���66��$�D��֚]���W�+�Li^�ب�7�o2Xx�Bƍ��E�`]�Ԍ6q�-8�U�%��4�i���P}kH�e��*�Y�YO� C����k��9gkU*���s�d����5��Og)�ޜ��ZB6�,:ڸV��u����t<Ƶ���,��Z�ːL���o/U������Ưz�)�u���Ss	g��C�L���������5P4�ƞ��WV�h�d�ǰ �8��l"Ϊ�q<{��ռ�NA��|��Gr����� ǚ��JA�VlB�l0�^�CS��ִ(�h�-SdP�M䲾�œ����� �vXV8�Ht���7T�Xza��b��C&8�F�@LԲ�b�7r�t$b)W$��h"�CUe������ �^\����:����	.f����-��"�X;rV�N��{�n�G���2|h5.�e4�66�e:i�9t��W���@�ы34|�tw[��8uhv
L�vQ�ƽ�Z���ʿ[�㒙ܱ6g$є���-���|%P��;NfP�4Ӕ3"�����hb��]��R�d��<��O ;!��c�[|r�������5o`�D�h1��ahM�/����ʽ�*�������J���+��"��y�l��=��$ܭ�R��nm2���ێq��}��uk�v�bNA���!�������w���Wy3uo��>G/y�G#�KD%�����g��-s�m�X��M�Md��OO�[������i;1Jǖ�}S~׸D1���(=�]Vn7��1�M^Q4����#T��w6�>۹�z�zt�s��������P���K;�[jܝ]VO�_7��'2�h٩G��I}H�.�r#�}CѬF�=W���}��{Θdt��iɹ��)�bK��m�W�<69��SbQó:�#jT�Γbƙ$���\��<H"�̩�����[�*�˄\����$;6�ue���"����)x].��:�t���7Af�4lg��%�8�ӂ�kTp�nX���z�=�1�u	}���ޜ���vSM��d8�*wQ�(�̘�9i�z�F�8Vݖ�j����9wҍ��k"u�6�	{i���x����=��ɐ�kE��>�b-p1��mИ�O�=�ZO$1�EN�2<jεysN2�����]u��%tk�^$u�ѕ�.-̦���U�:Q���ENT����"��Ohl
�NO��z�Sҥ�M'��J0]!�td��:���p�`g 3cZ:��e20)���s+g`�	{.�1{n��n��e�ئ؇_��V�r��R<������M��	@��r�9� ����N��L�KkM��v--��tN�p�r�� ��'3�U`h阘�f��5���"�uBg{P5�9n>�"]���b�*:��KRX�s�[9�]�d�b�X�c�[�,oI����]=���m�k�j�]����)�|�(�ct��[(��Ŵi�����n��k�"h�d���*C���%��yx�N��	-�6��d��n�b�8o���Sor���:Q��.����Ђj�Nw���oe&2��Z9���q\�����{l�R	fv+�1ˮ!��ѥ�ί���-A�@�k� PA]}R���J�i<�⼾������H��%46M��Wu�o8�k��<ת��k��b�i.�,9��;��p��E�7������Ŷ;8uF�����Q��A�������{E�rA݁��pR�R6 f�Ewt$v�6�������x:��'��$s8�IzQ��1ʆ������8J��i�`T��Sz����s�ȼ/���f�9�6���t�,�49�����z]JQQ��ҥKvʵ������9�{V�ͧ����F�
�~���j�z$B�:�����o��p�(�iΌVV���N:��[[9����qK ��?t2�N�9���#�9���Mرҵ�(�(��1��Z���������ˆ��Wl*���]�$��6�S�Θ��U���i���lN���pZr�>�)
Z�ٕ��;���3�*6p����cQq�7JV:�ػv`�G�
�IY�6q�"Kѿ6U>K�]胀o���)����3�\v�ķ�ٻϪэW$r��z����A�]��=3/	�;�����wZ� yX��x�P����)k���m��{[�]1��bFF��l!ӹdv`ؘ�q�X��ڎA�Î�&��7N Y�I�ɜj��z�5*�/P���F�ܭ_5([ē��-3�f�ѻ��� �U��ܳ�NFF�;���e�J���{�=Fs����fl�4��]͜�ɛ�4��N����F���3U�pJ+g	��av�oh$�Ǜ�x��kzgkW �����'Z�zb=�:㙵cY�_VX5�6��-�3g3;xf��CKӁi���K��L�f�y�bt஑S�-Nߦ[�u�)0��Ĝ~�*�*�'Q���v`ެ i��Ԣ8�e�aRnu��=���T�s�V
|`��X�i�����F�;��9��<�K���Z�E��R<�����w)]6-+32���J)*Q�U�N���Ws^�\� �,`ųn�8��IY�!��\���t�w�&S�YtK���i��Xk�<O�[�&K'�<�`^!36�V�,Y�{�A@
S�(m:)A$-���J2,��͝�yӊb}h��B�Q������tS��pQ���ԭk����ޫ�՘2���	滜X~51o^ǝķWʐ�XL�%3*�ݯ#Nb��k��N��A����}M�!NKC�EvR���l��{v����4V-�����O�/.>�C�z��wv�A�^�Qa�rQ�L=��ANƴM�f��lzn.�u�����IR��e8-��2�ZV�W\Ӕ�e#mVV>׬���t8ܺ�)Y �11�
*��{�ߵV\�,����.�x=�͵j�ԺԻ"�5��q�r�W�PqR;)eg7��=��fr4.�G�ν�*efg`o�':`�7z)]��ϔ;�Y$nj3��x�f\�}��	�@`*�t��9l��	���JA�9��%`�+���^�v�Z��77xZ`9�Y���B�����Z�X"�6��eX�[�W*�܏i�9b�1���[p���(���s���D��2M{�y�1	X�N�"{x8���w`�;��xe-�+��epO$�����\u����p��W��1vE��wƔp�:�f֡��cT���{Y��z(�6�II�ѥŞ��jlV�q�U�b�wb��w���sh�2ʶ�I#I 6�B�}θ)�-.�F՗1c�L�C
���n�b��j�;C�ꡢ��T�8����:���]��\�&��%�B��:��b��};�b���e�ݡ�zm�ls25+7Az�o����!�4��Q��O����@%�5��^<� ze�gnenEʺ֤��x�Xy��73�⣨в��&����fV ��+�֗i��; ����h�E_��R��|q�z�k�m���+b%�5x�4��1h�&ev�[hL�ix����f�	%�w�K�v��ۓ���0l�F�t^��v���yf+�?8��ݽ7Z��������!Yj�M�⢉{�z7v�sc�c�p�G�r�Nr�wטa;�z�r�8�ǖwB٪cR�wn:H\s]��'���N��՚��WP5��H��*S=����սY�nS���(���>k�s��[�:���k.�t�g#i�R���U/�������V�/����]�-*z�A{�e�!A��A��r"�5-�����8�EՋ8B�E�=/ ���]�>�"d�Pl$�]�j2{t����5�;q�`������B�j�u��@a�{�GGV�4��1˪�&���tbX�G���E�Z*�L����y��[V�&�vZ����#w	��Y`<hihT���rf����	�o�֜:w)�ƶ��I����z��)3/7�6����%���f��c�-�I�so$�� ���-wk�"Y����'� 
�����1�e�D�V��l1�X�rSR�
����E3��@]e�]��}�1-��+.�P\�Qܪٜ�=�	L���mj�(���T��gq�tx+�:�uN���j�(R.i�]��n�zαn�gN��*�ޒ�WQ步�G�/^3"�q��қX�B~e��fQ!��3�ݛ�H����l�O��%��h#S��YO/F��:��Ytk*�)��p����9�
<���ٰ-�R�E����j^u�@�t�RB����*�3:ʍ��Ѭ=��;�=xl}�U���{�/Iy��F��Ռӣ+����')���ҭ����q�&M��wd�]�)�t����1�+�ܭ���M�X0�;Af����4;2^�3�D.�s��ԗ^ŗF)J_���wL�[�ʇ��oj��)�º��� S/vk核1���$HLa��7z��c(�˝t�3��v"Z��3v�5W��ҋ5��fMn.�#�';0�<�6�1F���Ǣf��WW��&L�Et���+pʸ��#�k����7�cS�-���Pq�k����;]��Rٔ�:���;.�b���ʁ�'8(��]�X�p.uk��\E�nM�@�Ө�ۜH����e�_7}J�V����;i*�I�kn����7u*X �v_C�2L��u �قƳ,�hJ���	*h�1a�Mቒ�\7{O��Ib_S�<�N���qy��ˤ]���*=O(��ƥ:�9:��'6�$�&8��݄]
	ڸY�PZ�R����@�݃/�S@�zVdil��թ�iT����W;����S�b�Z�U�����#hIعW;8��F�D��e�� e��:L�^���a�������u�X��L��-!t�K�g�Po:�jW90i�o��0P��7|�4��f,9Fde!er��Q(���2gܡ�X��ϗګ^Q�V�ӱOQ�p���83uŪ���\�G$g1cV�=B�iM�Ġ��2(��6fԾWjK�y��Nh�.`c�
�WAcFA+�$N�M�U���*�H�g-�%6pR��՞f�ᮃz�n�Q���L��ά�	�(��X{o�e�c�s��&Н1�>��BW�=7�7z�"�\}�E3L�O��j����qM��(��,0�m����ӧ�����+�Y�kz=e����7�@��������Z�9P�9%H��R��7���5�ʕg�9{ر��hAR����\��������.���:vV���՞����Tj����d����&k�:w-�i�e>b�ؼ �.0�XG�>.��=��\�K����v�ZN��1���AU�u��5�>Z:�n�V�MP	����h����ka��Wm*��&��t���'*�G9rҨ��,f�d�z{~�3�'Z&�S�,��W���N�A��/7vvu���	P,\�/���)H��y�rOQNyj���.��٣ ��i��կ�@�9�zp��fӣ��]��ɹ�I�RK�`�(��)oJI�u)f�0�=��ڳ[rF"��Z����ɞ}����Cu��*w��A`_otԆr�7��;$؝��K�:�ǚq,��SuTl�4wN}�n�����v�2{4�)�n�����5�Y$]�|z����R�'>�۴��ïj�lժ����b-�5c(q5�{2�0ҳ51�,�������C���P5�k+Z��^���'�\{�&ܢoC�R�e������:ڱr6�lO��L��ndi�/��NzD������=�c�]�j:n�}4�r��6vm�dk`B!wR���.�k:�������o��w����,b�e��Hl�g��_i�#���Ԗ\�)s�T��h�Mu�a=��ۙt�8�+B�vf������ ���,�j���kUȵ�E�x�TU���u���u�7r�s�)�v���v�Hsa�O��I��u�����w> 1t����Ժ�&Ke�ho;��in�6?��	Ti��9.9]qطR t���}t�3u�@NqN��ʘ-�� ������yW;S��8����D��:�1r�ܲ$87{A����3/�β��K8m^��A���U�d��+�VUա��E{�g
ޙ]Ɯ3�6���;:���;uɬ�6i��5�����G6>F�cy�.��O9�KK���s��ڌ�uo�u�垦r�sCe�6���c:�7l��
�1l4	�<�bY�Ԩqq�uݗNcN��$��S.t� qW���z�`��t3Jf���ї[i��fTU.�-�	Yr9�:����E|���y�L%-r�/��ޭI@;�r��v�X��)���$�tX���Y��r����B0t}Mm�1.�~w| ��r,�gv���̻gS+�v�%"@u��W<e釷&�8�<׻C����ŝH+���o|��G���회�����Q�Y���d�,Y��uՉA|���a7ia;�E[W'�A٧B3\h#mԩ��".@��
dʬe��p�F��]yN�-�٫We^�p���,����S��"�%�E]���sY���A��p��� �E�8,�;���2�����V���-�тbŶ�De���9a���"q�b��v��OkH��a�U��ުYƱv3�om����z�;a`�:�ZG�ʇ��ӴQiΩ�2��/���q<]��"�-v*V�"�QWp�ET��n�A=R�â� 1����ϏTZ��q.ا:�Җ{��GdJ>U�#ށ��7#�'�=��<���DWj	�R�G]b���{�*��䣺JXz�h�}m{IJ��S^mn��+����8���WL�WNK�#;Oq�*J��7U������Z3'te��ENw�i�3!}Ym��kvS���tJ�Y����9�Q�ɕЍm�܈ȵ�r�����T��2L׽u�,�#����:�R%��@F��Ӧ�g��4\d����崨�!�i�O��Q�����^���eӾ��A���ek)q̪�(�d�N�;�v�v�����zk��\���YP�=��])�x�ڂYEމ؈i�㉝�]��O��ba-u�n䩎6.���P�xm�vg�^Rw&��Ee��۱�
�'1�i;��>��`D��wnL9�Q����.L�_�T�'JC�֘�a���gVY)@6qJ��TW��ed)�_t�*�����r�3Bmaɹݞ���K]!�-���͖�f:D�ʉd��s��5�h��S�x����D��}�ݯN̉>td�#j�iV�[o�]�c�OBrC��Ú /�iON�D������"$�X]Hb�:������DOd�C&�1�Cz­}m9Y�5Kt䲿���6?� 1��_S���޽��H�퉨��S�n1�L-���)o�+S��+j�ۤ��*e�뚥�7�Vt�T��a��`ŧ�6�;s2-�C��`3������[{6�6��,��];)F��j���Sn�;׼�u��3�F���*ݙ������_I��6����R�w{s*�G{�II�P�
���g�y��H:���H�='f'e"I�.��`��)*��6��j��L^���m�X��hyg��Ѵ���cT�U�!A���>ʽ��Q�e�x�4���z��Sq+U������@嚰U�'T����4��Fv���l�[wՎ��2�%E�"�w>�ZE�Ϝg+��,5���S�˕ց������\��4G�Neo<�i�%x��{$ �r�Nern���t��Z��W�������U�\�hR��`3��|9�ԲZ��]:LlЋ�Ւ_FNvł@�!��'�F�M#�j�p���P�*��gV�tv���m`��(
�@�ք��{�\b��\ޮ�v�;�HO��E��m(�K���X�l�����y��KuRYu��T7�pM��e�:��&�W� �0��Y䫆j� �N[���{n��҄����i���]]�{����ݚz�����'�9Ǝh�s�%_ �Nq}�.ѻ���W
z����=�4��ev��'Y�W#:8������i�:�E�պO)�#6!���?h����a�ޭ�T�T���%I�j���@�
To	J�S�C�e������Yy���F��y5ƨ[�l���Z�o���7YO%C�Y+�w�L�����ՊT�o�u�h�d��bS��ׇMs����ڕ�c��+��k����?���,���(��s+@�:enR�g�/��'Tuݣ1�1��,^=�(ܭL%3��b�����������g����F�8*ү��elV�� �ngs�6�qT��$�Q��`�+�a-�s6��)�	���f}�xġ�*&�
��woE��@b`�n���i�*�Vi�SzJ]}MiB+��Jj�r	X�v�3����U�b���s(c.�爵3jK����R$e��v�ƶ�u8�{X<�y4˒���*��Q:9�˧(M&ɷ���|�,��:�1D�v����;ڸ��0��ΙwH���9˨��9�4a�Wq�����2M|�W����
����,ٛ]��-����@�s����R�6�fZ]����P�����fK�ךr!G�Rw��r��]´�#C�Į�A�Ǒ�Y��(��j�B�_r��u*z�[}K@�pѻfp�q!�7 A�`�U�7�:�˕Ի�����P^�yR���z潱+#A��7.��lVj���)�c�tvȟ3>Wl��I���-z7r�b��X���f�m+3"��Z\'V_i�srtm�M�+S�h��Z�Vꨒ��jAQ��4Y�K�\�F�{���!Fcr���`2��unH]e��{]��v��6�ghK�799�B
���J3YZU�|؏�d5��4�}g,�6E%h�%`3��6�>��t���	\��8IG��Z�n�$Cݵ�H��ғ�f�b�����%uf��2����8��K� m%y��e\2��m�Q��͉�pJ̡�b�fT���:l����X�4]Y�}�nR�)�O�}P٫aRd���i'���^�α�N�qv���_z̋��n��Y�DhǇQj�,�p�Up�`c���&��E���'��T��9�\B�K#Oi��K�E-+ӑ��-�XcǰF����O'��/ �ܸ����ܘ.�[nP܌�V���W�kc�B���s(�y�>u\F�d�I��akK}�p^6�^�')v��2v��N�e�\;���J��L�
�]�u�\�::�M��̛xֆ���חf�0���v���Z/����I�_i�Ht"J�
n`�����J�ћ6�}�͖�V�S�cja`��t��uy�mZAA\�T2mYi"M1����ڐ�;��N�Sp�[UA���]�2���=���O�)�C��Y�x�tI����Z�].C��^I Z�2m�»f�V�{��T�Yňg3h��Jp��/z;��4�J5�ڶ�v�.�ݻ�Hk�9kS,1|���"�+��R8Ǚ�K�v�y�y��7�lK�|��p�XPi�*P�$9���Y��cy]#������);r�B��K����k~�N�ǃ*n3�{�v��.�a�-,b�!�ګ�3�y���t��c�vr��3U]g��=��V7n�!�<�;NO=P���1BU��n������01�S�;�u�K�Ku��#��ur]N��z8��I\S)V���9���2���fM�8���W1ͫV8NV��m���v�w��p�㮴p�;x{ff2�����'HUA\vX��l}V�]C��/-�wa"S2�5l3�X�Ub�U�T��j�|�P���),��/�ɋ@RС��V�G+��{%U�Y�϶ܕ�m�Y(S�Q�݄O<7����̩�&>��7�,��R��=��Ch�$5�k{��&�+0���D w��J���Q��r�5�V#��OL!k�p�����c�dٙ���n�C)u[�3��"ڔ��?b|-)���40�=Z;n�Ҕ�����۴%rG���`ᛪ>mm1�$.���u�}�&B%Ob����m�;H_Y�6YY��J��w�w*�.s���FH�(��A���6ۂG�B�h�����^�v���E���v�{5�J���̞���2�
e��m�t{��@��Ү�'m���t���|'��V$.�8�I�Wi�Kzō��Ԗ�4$�`�@��ѡe�մUvN7��i�p��A��("�xeƖ�VPס���!�u]J�]K�n�(�2���rb�(m�f�.)�t���U������IT �<^$o��Nٲ�4��k;6v����G�[J�+V��'�Z�8:�ن�݄EMᛤ���ժ{F;�d�~���,�W�sǔ�TWnu��`m}�6�D4=,f�t,�y/����Q�3Ҷ
^����BqV�Yq��.i�,��<yӢ�dk��rZaZ�(˺��e@[,kb��D��y��r��9x,��VĎ� t�<x��
�VK�Y)�\`��W2{0�PyG3�m��!#[��1U�T�@�!�Tcym�@�N���hqX�1fǑ����ݻ���).agٮ�f]\t�-�jż����'&�e�Ň�;�ɡ��`���뀋38��A�V����Ქ���m �t5*���z%��Iw�����x�A��@W��8�vY���m��g��X&m���,�<i·(���ZF�@H�kT���<y�rQuٌ��M[�kfr���q�`<��d�X/W|J]�{�J���<=G��ZJ8q�z"�BVq���i�{HܱJ;G���i�<�e������G}5n�`�Zy�:�cI�i�V�G�&n�V����*���6��p�QB.��C;��1��gu<��(7���������J��],�ˑ�]�k)�}��ſY�r��$`d�1N�!�k����\v:}>AB�q*oU���R��3D��?m��lR2�g^k��z
��C'a��kV�����������V��5R}�|�U_uYS
w;᷸����XiS�T�[�j�]Fe(5�|��Vo��?-Ekd��U�8;u�R�;nVn3p�C4��H��SX�0Nzg\�.�q|6�(5DÊĨ�e�+��[CTq�+bx���k�*�՗\��/o��ɎE�o�6�E`�g�E3b�BwF��wq:z�j}�"qɫ)q�T�F����Pb�ܺ̈��亙Ϻ�Ï��Nⶴ��,Q��ʇ�bV��{4"�g+d/Eo�C�����{dW�r�Y���4!���jD%-�� )S8��9�)����c�h����{X�-�v�����9c#Üy� �4;tk�+i�k��]�3JUi2j1�HwS��[2�u®�oM7��i�M�%���p�[���"�uRV����+�Y����c����ÒF�<�n:���t1��w*����B���t��w�/EcA��拭5�K��5�l�
�!S��I�t�,�Q(����w�Lp�H�/ 9;Q�!}p���c׺�;騛��T�s8�7T�28� 4Hv�w�-NS�ܫ�u��^�{a�C]$��hv�Q֕'��Y�e�.���H�y�%��F��v_�x���ڬ�gL�8<���F��Am�R�U���OZ�V���=�}���ΛOT��$��*�;�`Hd�T��`X�G��,���)Jx��ޱ��F����/����̅]�G[��Ԟ���&�7�9�UX�ӭ�p7ە�h�v7Mܕ������Y)]�1>�y�Q�Lv�����JG�.�2��YBro�7�R]�ܥO�\��3�+d}|r��J��Q�P杶q�3�!���n�g�nC��'|U��6f�%�oY��v)NmdrF�[��E][<Ne�pqX�ݓj��k^쑢٥����+A�v�
��F|D</�M�\��5�Ver�h�����"X*N��W�N�����y�@ݫu��
���љ�H�bC\`�c��Ղ@3Y��4Γa�e2y\'W=6�'	ݹ���\JN�k�LR�ci������"���޵j�e�ۻA���eѻ̕�����<���by�k�|����@X��ŕ|�r�i`�ށ��^bB����� ����E�N�&+�M���s���縔�y#'nfm��xH��`�\�ǞNǲ�F,���M��(-���ohp�-���]X�ȕ��֔�١Y,�˦29ư�t�d�$�%�u���|�y��8��:,�I�6��@
���t��(oE���_R�]��\��qլ��u�k��>�Hv0^����V�ovf#�#��j���[p�%�7�����"�A�KE�7�Tz�{�n�>f�f��d���ۧ�T1s�TOfL���&��CA��*��#����(:Ni��G$]<	s]�En�k]�.,��)68mKo��s���ݪ���{slJ@5{���
h��un�N�:�i�*�gR"'�1��'�꒺ŭa�%e�+Z��t�''l��tj�c��˅	�i�����}�9V�6���;n^|z�,V���{w)	{ԭGQ*G}d9n��gS��C2r1���!c�������ۨ�TZ�:�L�!)���&a�y�#r*���n=؄<��O�Z�[y�N��g`��ڱ<~:��|���{/���T���ʰ�ڇ����8�����R1��S��u6� V��,f�Jݜ�Ͳ�8r�gA��Gy�'}�������߄�,"��4��ס�N����D;�t���y۶Ә�@����.��+��M��Q�V�2���6�*ւ�:/^p�;����2�Yt�Q�ȹIǵ%��jY{�m���!§Z6����7@�a�75��4Y���[wf(��mL������v�]��:��)u|Z;�-��B��
Ѹ���iZ�v00�%�6>
�@��&o��U!�,�t kZ�P����7K͛y�˔�������0SBqXzj��Ol��a��rN&l���m�̢�։�qW'��4��Ծ{�W���h��agك�p������}	�V�ݑ�/b��d�`R`�>�^��>z�ŗy]���h�_b��1�ChA��y�����Q/.��&�]����y�4�C�Xz��O��v�V���җ��H\aq��=g��a�YK3#ݼ,�[����vZ\��7����ԭ���Q�k�V��q�9���L�c��4�)��v���a�ړK�^폲��>�i>;�R�ڲ���O�E��� K�A	�I��Ϫ"Bˮ�ә�hx���F��d�t��V# �i��t����%މ�U��#�,nŞ�|��9� ��qʰo�b�͔��В���v�Zi�y��V��Ow�s4����Emu��9u8�L<G����q=wz� ���#]��*�mM�m_+(j�����G`�卓L�61մubbT�ˋyWE�j^�=Έ��0�{P�V�v_Lo�^:F�R	X>�c��ty��)b�6�oseK��ޡ\�Z��`��T��3x��W:%k����ͭzp2�.�M()��L��{���Gt��wI	��V�����&�ًyS'�He,���ڐ
/��0�;Cz�g=R>c�����+��Vcޔ���q����˸��J�t@X-D� ��-�5 9D�i\q�-�˺i�����E��3o�bj/�-d�QM�v-�A."�A�`��b�70�쳅gβ�mwI����_a�.���v����$Q�\8i��0��\�.��b���VvX������Pi��c#>f��۳CL�o\<��<��;�.Nw�i�0��������u�!H�tg#��.��`%�J��3G&��2�����岷m�+]�2nQ0��w�d���r�`�N!�4jo&ͥG�Kw-���{grL\�+����HB�:�ݬ*��dK0�jT�`.���,[ind��J9����\��WAM�:�]R�txl��1j,Yuq��jFS%������X!ң�Ҽ Gl҆��[Rƺ>%#ľ��1M>n�^����xn;0���+Ƹ˵bdWP���q�a�S;����t����S���lx�����&��24�{�p�;'1��ZR��AވfS�y𺔦҇����ٛ�������]K�@�hݦ�V.��&��mݖ��c]^�7m�6%{
=c:��PQ�m�nZ엺�Ѹ�,�5h�2j�;TVE�<���������oG�|~�[.�n�%46��IEv�v�`#�qh8 n"�`�4�K�u�.G�;F��yep��������:}P�R�;��^��N�qY3O;�E0�һ��3���F5�(7ϛ�K�s�Z��&v�Vaܨf��*^wz�������*	���'���*�'��fgB�Aו���J���+����%��{l}���v9�5��+J����[SN�{�o.M�,���r�By� �i�N���еS$t�A������������J�h�7+��:�Hg:�2��L�8T��o�Q�'֝�Ρl;�J��	oH�Wa� e������@n�
hu,�3���8�$����E���>����J�HY%��ɡ���R!�ѵu�3��G\��R�^�:�Z]��)LG 4.�m�^��e,W,K�k�²�7ݫO3�u�nc�5b2���.�'Z05n��'<��6+^evޤm�51��[�9l�J��god�/BGjۡ&������\S閾�U��8����J�z#�UgB �S�Du��[WY\jS�x+�Va��[I�V������z'�w	����*�#`&㶡��SӒ�����#`I��u�j��$�5N㝹�C}Y�Zuټ�o"dɌq��s�eG�g/�[�6�#;�em��o ��%u�r�.�Y|I.����ݜ�4r�ԖYG�3.����;���J�~������_�*�$̩�9��S)%
��)s��IB6�uԐ�鉘���MH�CD�$�*)I�eV�\�U��34T�1i��V��L̬��h�
�H���j�F�R!��fHMD-D2B5K1,,��H��bQ�6���DH�B��Ugf
E�BDu%�TTe��H�Ȱĳ.�Z�J�QM�Z'@�5"-Z	)�m3C��U�Әe�0��2L�-N�(X�b[-" �h��DE.�i�ad�6*U\��\D����R�:XQjj��"CiI�I�Z�$E�'(���FI�B��f�D��������ΥI��:I*�I �:!�c~�e���X�X:�J�dK���:�fӾ�uL%6�v�|cv�'2���L��]Ptm�8�=C9"�9�}�7yΩ#6�]�h�*�X_h��l?�W[9�j��I�R�t�x�]ʚ������]�2Q���y9+G׏<��!ð�5�ԁ�r1�%ѷ���߄��qM�U�799�VB,J��w�1��ʮ敭���������~�Xw��r0�����+)�kY�]Vf�7����I����O ,��,��(�`���?_���^��Rn|���j���I�qS����g�4/�9�}X����k!�1�-�O��(G^Up�"o���ߔ�隕^��E̚��נa�O��0p
�g\�Awy�9y���W���������݆�셙����5�U�,��|W�:+��([�`w`����2`���Lk��������D��U��7�$�	)�'�Em���l�h5(�@ݤ�ɜx�ުel�t���ә!�*�m�u�����|r���LŢ0p�UN��C��[K�z�����m9��~��\��$��m�;Kg�d�>��d��NS�N���!�Y��x�Ie��_R|��Y�З����aT�ѐ�t����S�CgU���9A�)����[|+��r`���M�x��5+��z�θ�J�j��γ\�(h}wD�S���dtځ�.�l�m��<u��PLf��s'M�#E*Ն��Lq9j�fM�8�w�m��NL��B\�!�P���ۨS
������2L���v��],cf��2�C�&�R.�H��ٓ:���ps��@|�+��c��PL2.z���(˫C�!u}�`V}Mٱ�*��B�|�D�M��)a���l� �DTݡ����$��="�;���4K!�Y�|�c qdt�͵	�!,�Ͳ��
�`]�-�v��n�^{w^�ض`9�@�x� ���S����Ld_P]{75%����!����G)hX+zP]�eZ߻�@��0(d7��x�5d����`���c��~���|9Eg[�����&�����-��a�ξ`\F:q#����>���Ѯ�i�_=�}���<s[�z�V�lۈ�ٵ���ާ/ u��9�������9��u�M���n�f�sy�Z����巾-�{ꢾ�0�FN��=�fs�C�A�!IW!����tx6�(��֗�������ϙ�n�j1}��Q�vx	�f�����B��i�{~�k����*�U��[#�b�Ü�޷r;���e�8�W
�.�f��әq�{���ڡ��*�tY��u=�U�O���O1�3:�ɳ��ݾjL3]"󱝮�p-�VJ�X�Vgi)R�:�5�U��Ϧ"�^j�x�j��ZH؛s�����a,��4�kOC7n�Y���������KG��.�.���R���7N*�q}C�~����v�|�3�Gω���A>_z�AOU{*Y���|��(��g�V��iz*Th�9��Ǟ�=�$�9kɛ�g���Xz1�l*n��#8Q(¸�w>+�匴�8���ޭ����L)qT�p؇�t�,���E㟲�jw]D�ͫ��k_�sr��@F�U	�Y���6 �#����yf2��긧�<zf�!�9��k���A����_�ޒ�Ӝ����y�R��U�E��*L�\ĉ,-؄/�6���t���v���^���7�m�O[ �Dg��|�H�p�8��x|;��cWC��E��7��j]�r�'�bޥ��V����WL5�^��m�ϝl����F�r@@��s��k܌+Q�x���8��>��2���xȎL۠a��0�!�k��(ZT���U��^f�p]>!�\=�ԗ�}����ᐋ�/""�E�I࠘��86���{������-ē�{���U_T��W����H�ԓS-�J�<kl�ۇ�3Y�(s�(*��S9)�ݴw�V�u�Į�J�(l�d�ۨ��u��[�Ѵ�X�.�o'w7��>��v���ɡX����y��׷�U�֫B�f��O@R�����~�ǐ��m��h�����G3�%;��LJ�mә˭��8��j5�~�3��ٱHE���U%����U��0�z���Շ-+�1�ԱGHJ��f�Cm���C$H�z"�U�L:b �������ϸA��ӵSOx'�/Zd��,ӹ���$����/8�7�##�\��2bT	˃NF����?P�]�Ǚ�P�?�ƈ�:����-���X�̽�3�AQa��,F�s���Sٰ|pS�<C���'�~�.�\N̠�r��`�;���6�r�q=p�/�j�FŻL-�3؞ri���׮�Ƿw�vx@K$�Osn���q�4�S��c�e��C|���{.��7I��n̵�+H�@fQr���&�����zLI�s�Wu��QQ�]4�7�l���0{޽U�y^�>Z/ȭ�Zjz��.>B)N;�%:�=Aƺc�<��)�6�n�������q�����VI|��j{��~OM����R�o��4xC�xS�h�=u�k��ۧ�}�㩐�л/�f̬8��X�&�=���Ԗ���ԩ`���i��#˴{!.�͍�
�2������3]z��r���=X��NwW*����1�ye�Mk���Z����`G�90��[�����`�o5.ΝR�(jYV�C%��WS
RF�(����qnp�3�UN���DT�y�~+���+�u��!.W����u��;wF��L>Ү+��3C��'a[��l��hl|�f/����%��G���u����\Z�^���ލB�LG��g�����A���~2���3�p.x�&R���R�Ve�,�<������@R�Y�VQ|F$z�&ԶU�r��c��%l��9��m�~�[ގt�2�X�M�l˃�b�`��Ŵ.���C����5�Ժ����=3p2�e�����z�-�2�	ۻW�Ѯ�+n2i���>�nya,\S�te�H�c�'2���j�Χ���~ri|+&���}������>�;�\+d��''k�2��;ۖ6d�B�I�g^�L� F�#�iW���52\Ӝ,m�{%�	d59D���Xd���4�Ed��kT�{�o�y�];\M0��=jl�C^��{R�@`Rf�/U?-9�&"��!�}���N�o��d���kG��>�xl�0<.�g9�������q���dl���U��O:�(�d]���Jl��."X�թ�I��]ނ�fMS���՝������VQ�T���C�e���R����;�|�^1{	��pQ��=)�kA����v��]���@���.�,܊���on���d���H���6�Lq^��*b=O���B�{����܈u]�{��德�����@�[�4�o�Ϳ\e�ƪj�{���}�͏݇6��,S,�v��+r�M�2+	�����+r!�Cf��xi��`6MA����^��)�Ɯ�e��a�y�-:0��5��D����j��Tdl���!L͠�� �0&\�
e��ož!7:�bުB�����z�ŷt���%��P`��=s���K<��ξ�:��z��4�<� ��񬄇�w�o��o�ɝv�}�1���d���W}8&k��Ck���s�6��τO
�&$��k���*͌9Pe��q����I�S���>���5~^��w��;�)��y���� ����OԺ݃a!�RϜ�*n;,a��Ì����[�MTh��!lx�  �� U\�"��q? Gx�ʏk���Y�'[�Q��#�Ce�v���5P$����Cn�K�.��X�WO���5�9������L&0lX�{j����I;�r�U����[h��j5���M��,Rk�s��}��!g���^�%mYea#Η�K��Ds�]Xӣ��� �/:V��By��R��)#xjV1f�K�,�ڵ���X*mC`���_�ML�i�����}���x+�\#�����Do:��c�;>o;����@j�u��+UF��7ao=umѨ:`��g����d�ĭ��N��[����ׂ�T�_C9�ش��z�Me��%p��2��l9v2���$ۍ=jfo]C���u�V�vX����w@�El]K�E/^\�5�z���Y5O<H�0{���;t	�Y���D/#�^�1��Li���wE�>��us�࿲-F�>&��+]K���7NTCB\�6w�k��һ�`�<��dN?�t�]�y󕁑���gVP�ƥ 4�O�#K9�!�/�Ay���ŵ�&��|���D����=�޿���!�FO�Rh&���2��+<�ox֫��r�HE�;�Hbʋ���x��eҜN�X�md3�@�c�~�N_�*"�U�����������8eh�d$?��ηK�~��y��k�������`��Y<*��^Qkjř�\���e�2g�a)��9%����\�E�;yT<B�Q�����2������aU�̝,���n�3������;/['4�{�i�]@E$d�܄��h~`�v2��wG�Z��ݫZXm���;�f�.g]��z!�]��ʣ�B��m�Na�[Zo��a��r��k8YJ�]�%K/)�,���5�i��q>��P~�͖�>�Dk�|��'�!���Z�5tK�\�SKGX=}킖bK���pٯ�oYc~�U����^�ϛxfrl�@K�0�^wq�ҩ�c�;�̝��E�>�Y�i�ؤ�O�t?*��/�g��}���_q���xx>��΍���QDglv �y~!\B��|t%��T!��
�Ds�B�b��z(�j-�aYLf+l��Ʒ �W��hȪ�c������oF��;�ja1.��Nd�:�J���Ou���vwB�{��.��Lt1WKt�זa�9Ja��8�f�9�J��U�
�mw?tg7���V�h�t��yS;hS�(.Y���+�fK*i��<n��b�^t�����=�L�{gz\P�:7-)�K�]k�yM��X��� �-�K��G�u�[����|<j��p�*���1�?6�����6n��a���kG�F�|Gx.m�}�k�aۿ��T�9Ⱥ7,֎�2���0�,;��<'n;�Fx�(����f�Y�u.�c���� �T��=�j�]�g'1v�]��,KddG6C��mϱj)��:��3����c��U�5��v<xv#)���0�f�4n�pe� ��R,�9P���Y:g���6�14�]�m�k��z�o�of�9��7}ګ�4�@���
:�PQ��Lk��[�v�3��0v-ٖ�j^�Φ+ �ٸ́��L�^���@�@V��qTT|.��!���8�ة���t���C���+��ʍV���ZVp�ˬ�+	-��}� ��0��)�>�|Mg�dY��Q�~�"�s�bB%��s
 �w��_��y����߬2c��<�r�
t4w��ݯU�.p�����q;Ӛ��/0H�UP���yS���y>)�@�R��:��GYP�ݔȯFiv�z}S�6�]rq�'~V���hl:�ً�7p;!��e��0AVd��%t�>��%$���?�ĺT4��ώ;�=�!N[~��8�N��D�0�/賻;��J�{�o�������E* ��&����ne""��R�\���	+`<�yՒ]ݱ��!Y�qE5�wm���2�Ҷz�\@�v����C��Z�\�K�����@>1z4�5�%�Wm�{w{~�����:�X����Ltݥ�V%���
9���i���gU���MAU�kQl����=@��%�:�U-���{�ו�W� �}ja;v�؄Mf����y�W��{��.�9�I�T����+��Զ�H�7�����27R��.�ua�$Ռ�&�X��4�����,�Lۼ�b�5�:�t0��w9-���pv�c�wzܝ̺��\�+�zf�dE����O�g��.s�Ji�Q3��ž[H�ڒ�춀#�L=8�쀪�Ĝ_0���v�4$#$`�@Fq=O�i�t�I�O`�ND�8�td�]m�����z���s[v���1�S�`���O��H��H�<���J��rL����h�]ea��}3�x����Kϼf���	��R��+�����'��q�200{����+���~{����}Ȏ�J1��s6��k$��Z�ۘY���*m�2��t�Fx�+���7!D�S��:,)O�t�T���ݕサ�:a����M[����rF�
@��jD�kfT�����yT�iv,[B2\vT���J�Pa���_��u�Ǩ0a�J xxp��rơN[��k�3�w��&0߳�|b��6"ۿ�L䥮�������ۨS	lSV4@�����rqܶ_#�� {_� k�5�$=J{��:��8 �O*�qxs���wA���9sDz���� ��>��o3o�A�4-�;���W��>sDI�0�n�u_SB���n(���U�VҎG�)�(�W�8q_�Z�[���{L�PGOg��0�ӳ��bb���h���S�	Y�qg^�F�����ҲC�&k��#w"6�xʘ�u �2H���I��Y$:a�6�C���x�oZ:Xܤ���]���Vu��k-y���O]EtU��\�*ȡ�ԫ��_9C��Le`��(smh�S2Wn����л1��k2���2%y����X��8��K�n����xh,����n�����;��1ؾyZh7M�u�MF��l޳�����ܫz*�.,�YӍ5C�-���՚���	�-�;�
������c��W�e�T�NX��;3s�Ū�xR�e]�\l�����I�8
F�B�]�j#F^�J��t��;L�*��mk�)���F�h33b�Q�ᦺn݊�n��T����,S��J=��\c�	��â�ש���������n�{s�e��YL^�M3:������%V�k��	�NLA��v�b��\gj������|r����W�黸9`\��7B�.��<�SF)�jJ���p	6ᲫehF�>��ʇQ���m���$�N�qt[t�j�]��"����S!���>廤�s�]�o�����a�k~Z�nKX��%�«��ܧ�/�:�����Y�!KGl2ٮ�ϋ�����[y��,�cW���猵����g�:��Y��K�4�3��[q��u4���th��)qM���5���%
���'�ǅ��xm�'}C8H��^#OeEx�9�s/HKZ��I�f��V�f����.�9�3"4��nZ{�)i�ZJhnC��l���A`_D��Xs������������#��`�哥�2n:e���Ѽ� ձ^-�u�JНg)�[�t0�jY��ޘ�z���9a��4��<�S.r��γo-���Cf�;�Q����[��U�b���Y����"/��差�JWF�<�k5֧�W9h6�v���f�Ņ���}v���Ȭ��0�k)j$�uLQ�E���i(�{Yɓ�gq��H���9�����*	�
{��<�E��� �Mh�Θ��L�B����:�7+��۩��V���k�n#LZ��"����Y��vjCMj
Q�Ϸv5���e�B�̳.M��p��t��P�qQ��͵d��k�;M�}w��<�(���O���C�⬗u�d�t��W�(�`XҚl�)��	_e��QD�ݱ=�/#���7���2$�z]�e|�v�\d��-�؎]�����»8V����X
���]]��A�Q�4{1T�|�'��X�1o8��2�:�����$���m$�.�v��K�t7�d][OE�l������Z�֝2� ��:���,��"Y*҄L�TT55*��d��Y�2��fSI"Q9)s��NPi��Yf����a�I0�H�EU��!j�R��"��"�T��YD��al��9��N$i$"�f�R�ʴ��ºJ��4YFD�e$&Euit�+%J쪊�P2MCR����Qu	SeQƛ2�3��f�-�Q`Z\��i�r((�\�L2�[*��BҰ��-H���*��H�J��h�jQ�d���)Y����hUGU#��er³�"馴SVXE\��,�i�q6�H�-6��Q,���$�gB���2�D�\3+�����FU��I���B2C�ԭY��AΘQE{������ϧƠ�iWH����u�;M��s���'O%�UL7�u�Q�J��e�����q�{
��3*P�];��ƣIϏ�����}L.�����6:!�©��"����n�A��t�_��N&��~�ۿѻC�|?|�T��{������<v���.���#~��s������zˮ������]��Ϝ���o�������o�'�����َ��ڭ������N�a�o^9w���p)��=�>�u�����i�nӉ����x㈦#'��f>����1�Ǎ%�(ǝ�b�;%b�~�͎�g���ږ�v���������n��rަ�=�;M��k�/�o�I;������wH~w<x����m�i7��q��G�+�������LGL|0DE׃��E�:6����-�@��b�S��>n�����~w��!�aW��΃��Bpw��u�oP�q�ۏ��y��ۉğ�_���7i�Bv��n/�n'q�}�L>H}����h}K?u	���f�~�������ڥ|����������{����o�����.����m;��^8���:���0��߼��㏏�8�_����(z�C����6��eӸ�O��x��n��f�"�i�D��vhv�{�艂�8�5�k2O�=��T�G�5_���i��z�N+������x������w���;~�q8�}���!>�_�p�q�޻^��w�޿��0���n��B���`����43=e[�_gydN�V/�bZG�/�xCy����l�I���|=��x�q���ߜ�t�U޸��8�C�����t�}O��B��';\��?���7��!:v��Ͼ�ہM�|/:�o^��z��~�Ͻ���k?n�w�=w�UxpC���lT�ݻI���s��c������v��:M|���;�8�!���:L.��q��x�I�]��&�����\���N?�<�q8����]���ӍfcS��cꘁ1��G�2��'q�s�i0��v��|�η�ݠ~HO���>��~v�|��!��n��v��8��q�o�_�w��<w�#�}N��;��=N�v������|��|�x;�E%�������L�\��W��:�l�w�˞�i�ۉ�n��~�۞������U=v���?!���?���;W~v���}N��O��|���:x���G-����m������֕�?r��X���������W�=Kn=��b�zs�n5iʶux��2����q���n��C�s�Y��fR8��b�}y���>����[��ٽ�&��E�,9��Pv`���I�&U{�t�׻�S�tEk2¼�:�j2�jܵ�{����7�CL�����0�;����Ѹ�˻<��[v�Sy���A۽v�`��z��=q��7�q�{�0t�S�O��xz���N^�}C���ϰI���ۈ�o���^y�����u��ߗ���wӖ��
���:܎;~~���������7�8�q?~��[x�y�Ğ&���~<�.���c��C'���ͮ�5�<����{y������~;��P�aOJГ|BC�����q8��� x���G��q	/�?���~?{ψv�z�v���z?���@�/z������w�<��1���~���&�O��vؿx�[���C�n;��ߓ�!����>��ۼN��~j�ӎ>!���(
(z�����a��t�/v�v�q�;����7��y�n��;]�}���LF�}�G��"=�ާC�����2��iǧ�s'i����}q��xv��'��~�c��B~�{��~F't�� �n>'H�t�Q�x��(��L(p�y�����/���~qɏL|gз��C��;�ݜ��1�L����{���A!�aC�}�|q�v���n��&_S�n{���;�����n�}Bt��lu��q<N'���ߐ����ۤ;�#�N�ny�}lՉ3��CW�w�������'�vU��O�}M}��w�z� �}�I����=<��[�wHq����t��oP������oP�q�?���;@���;<�I��ۉ��ߜ1�v��w�q�Z�7sC�[�k�kG�3�D���z����@����o;�i�>s�����q�?~��&��^&�~��ަ���8��'��8x����Hq�{�t�������9�L?��G��׿?����?V�p��}��~����>�v�;��:L.��u��o�q0�׽��W;N����<N��o��z��!?]���Ώ��7�O��{���Q�~؀�}@}���.c�㾾lĿs�:��߾�������������;��L/g�=���t�r���;��'���t�]�~q�.�}C�L)�:�St�8�C�>��^A&_S�￸|@�'}v����v�oP����~c�ǫ��oL7��3�{15Nk f3O�|���;eǞ������]n���u�D��x:7�q�MUl�����s�x���o�-�����G��x%jv���w����ˬ�����VoJx���J�y��we�X��RA�fn���i&l����Ĭ��9z�}�u���ݽ�r�f�a��u�����;H~�{��Nv�!���>'n:q+���&�8�C��es�bw�=w������0�ǧ;�z��ո�>!&����y�S���5ϴu��K���z#혊���s�ݠ~Iǧ\�I�����O��p�0��ߓ��to�v�y}O�X�O���&���ێ���x�&�������`�o��z�?��w�:�����<�y�nAWQ��N1���=?C��b��b�x��q��zs� �]�P����G�>&m���n������Nt�|�۟c�{��>&O�����c~C�
=Gn�W;_߸��q��㿼�_9O�Yܼ#u_���|� I���E�t�7�w���۴��b~w�]���?��?�}�w��������]�@�ˉ�{���w� ��'�8�;�[�I���>��7����q0���z��v-��:T쒽���}V*���j�e�<Oyc�Rw��έ�ۉ�B~�N�{N�����;I�ǞF���z���@��/��ۅ���{=��$�;q�]��xn�x���������=�E�ӫ���o̒s�M�������	vlC�q0�~ߐ�wn�ޡ��+�	7ף�S��C�c�:;v��N��N:O��n8�w���a_���ԥ����÷�ь}���;[�_�ի����z���6^q凭�羁1�?|g�?t�����q����{�>+�M뾼x�9�1;�������8����w�8�q��wˤ®�(���&,t���q�������aw^�r�����⦽�y5y�!����}�sD��z:�����&�<���#�n+������q$���������M���<���\
o;�{v�s����N�m��:O��;�j������iSsν��?=
���Ko4����c�b"�퟾����	��x��{�ލ�|L.�>s�z�����:�һ�����9���I��{��6�����}����t��#�t�r���
I����P�?v�|���n�9�s�{ѓ��O�	��b6}=�\.�vy�t��~N8�į���
o��8�g�tn�F'~C����|C�=N&��7�]ӽw�q?��t�?��y��&F�OS���ۈ%��uOA��4�,L�8���G!�-���ϫ 0;5h<����-s1�̲V4��VVWR�R&*��8y��1k=
D�ĪM\��9D�:��{�!W����$mT��Fܦ�>�!��f��bD�b&^�Wf�8�՞\���b���kvB�M��>���[u����{�۴:L+����&�]G=�v��;�i�~�ͼN�o];����B���z�֕�����<���ޡy��^�����qǥ�bw�S�8��<����]b'��q���>�����������i��v��t��q����'I���c�G_�!������ױ�C����mב�ۊ����h$��{��v�;I�B|���۴�/:󾩷˫�\�۟�jݝ��W�|�-;V�;U���ӾrL.�v���^ܻ�ҡ��M� 㾡�V�Q��'��s������������>�����c�w��뎓����I�����zgM����{�~�?|�"������-ӷ|?��A:v�����7�I;}y��c��۴��_��:��7����w\W����N�#�7_#�'��=wh}C�r~�����Y�w�kCk�'��?9���S���9����F:WP��ϼ��0��=�v����@���8�I�ӷ����
����p?��o�I�`��n��&�rP<Hv��:ܾ;t��/�A�7�w^\�.Y���o����g艓v�<zM��c�ϝ��M��;�q?���N�ǩ�߻�v�K���{瞝/�*���e�Q�F������c�o>�ܶ�6ɭ�UC���~q4Bp����ka��S���6"�ka���Wɑ��{t���8�����Y�q��1�U�|+��n���83�x��S���)] ����n�nOf�̚�Jf#�����q�yqo��J�_Xk������vP���(&��'4�7��^P�	SJ��sE;2��E<��Նڤx��@�|.��Myc�,��F�ga�vꔭ"oGc�S/���)�**_]Mؔ+�[C4$�:q|�rP���(�}���Ţ��]gM8&�옭9��(��^�{}O9˸�+.iۦl��ݲ�g��4k����V�t�W;(:.���w���2��W�N�<�[}B�X��9��v�l�×������߫m[��(��	vq�ܮ꿺d)�t�ݔ�ec[�T0�fByx�J�NA�aώ��e���S�g.��1cd%r��|�*Ɂ3R�38�؞���������p�ɝ��K�$9�c��AG��6��M�S���W]�p�� o�� ��]���Or�����v��2��D1���8F��������Y�v�6wSF�q���;:R�T]�r���B�B9=!3��'Z�i%N>E`�햨�1��`[}8�]}M��m��$I�8�:Kڄ��Z9�2�66�iL]�R�8��'P��{�pg�/�,p�9.E]E����X5�	޳v��k��)�h�ڛb��2!�dd$�>�Չ����̟x$ �I����z���n͵�sپO��ه.r]���]�o`t��nBҞa������H����C���{&S2f��f�Ε��B�t�
�s�^ÃeFU��%?:Q�M��_FJӈk(e����:jzko�Uϑޡ�
�� �x�5$��t��嶦�=7��1�L��ׯU]	ت�V���?[�q����[N���#Jr�}X���漕o���R)��.���Y�*�s�Vje�-E�L7a+�Uݳ`ݼp�4�<V�F���f��#�F���ӷ�O/�u\Ř�nyk�c*f�n�|���qh˻�+�^�`h�`�4�|����ae��zs�jx�xv�}��.� ̦!���)��*-刅����|�ݱk[���2f\nq�!�hLb���EO���y�N���p�u-b��Q�:^�]�j�zR�=��V���N%dHr��j��<�����j�[睁^� �t!G����9�3m�q5JM UGYw E��,���ȇQ,=�6�y���&�}�za�^�0Q���A���¼	�x��1��ʋ��^9�>f]��"Xـ4�<Sΰ;���5N�r21A,V���˚� �+�T��_jU!���K�~��|,M8�s�6'z&n�������wG� `��mr�e*YS=@�7lɞ�����,�7X�H],Q��K�nE���,e24�v�����O\;�5p����&e�s�	_H��ܔ��XK�Ҳ�i.(Lj���	;Hl:��loη�^���^.���:0��T�t�/#�+khۄ�u=ugjсm%*�Rݲa.�rk�K�}���GiG=��տ��<����Y}].�w��,��-��!�J��Ή8��Xg�=��GnZ)��l���0��f���,T��c\��J���ߪ����Kx��.����Ż��O��Du�q��n�˜uZ�{���¬@H�2 �,�.yo�y-��}TR���x��=��}���aa^[�?W��`i�K���=�Kʌ��yƍm��=:D4Rk.�����qP�e��T�~̩k~����s����죧����qɘ���|��1�;�-�-��r}���b�_^$>G}L���>�}w��kڛ��s��f¹M+�C���0�[�b���t�yS;hV&��n�����`ᠻ��i�<�.³RȚ�=-:ler,������ ɿFܡ���^��,�BrƐT.����_z̽z�U�#'iU��@!��"��9iU�1�q�mg� ��2b�F�v�q�{C�7|��pH��0ytGIoM1���ld)���a�Xr[��߮���T�r
�|��<�yn0�)vhl�>S�
s�"�)���r�Al����]��[yJ�,d��#{�g�HD����?>p{��kzc\o�4��x���m)>��+�w�|Wp~݌e�SP�k���[��i&�5ۄ:Wi�[�u�|���W���@�}����IqB�k@���w׹���vg�Y���s�):�G0X�(�a^G�`���r�� �#LC�͌�${&�#nnO����æ�r����j+]�*�\�4ml��R~��#�l�QxOe^t�)�S��ľn��5��ZCK��>!��2��7�h���>��+�^P�jӬ�����aҷ�Z��s��|n��]��>�`.��`�w�,B�ߓ��oɎ�FqP��(,}y<F�k"� S�9:7B`�=yS��Ы�UH�ċΗ�ۭ�dm=3���ٱo�v&�z���E�1��q��;��b6$oSCa�F��n�m��z����o�K�o�Hѕ澌j!#:&/�μ7+�+��^P}���R�5��P"m���Uvu���\���L���y���r;D��f�:<���DVj^2�K��®\>������Z>���b��{&6f�;�1D�:��g����=ӛj�5dj�\���Օ)b�,E�=�gSW�3C��{��i�Lo��~���ݤabk\gU��H��>�"1�8���2��v��<J������C�j�f�t��}:YX6�r�6���~����R��M� p1Ɠ�}�T=���
��P�4�7t"l��g+VWdPW�Wk9���Y��tI��}N��\)�]��z��eu'[5pW�eǈb�y\UF,�<���o6j[���WVVۑ�p��4�Ɏ�'�.�n?��zw���I��S�AG{b7���M#މǷ+�������WI�� �iW�����DE��*�!B���g��C]5������J��exe/>�sN�� c�AM:'�7�3;�Q�i�/{.>z��#ۈ*�j�T���:v�/�C �u�=�nʆ�o
��k�/3���Q�A߭����6S[�#�Hhg��,��=x�֩�r:��p�f��W_ޫSH����q�W��]/8<&,/��C/�\I����R��I��_*F�I*���lH!��Hv�l�×���<�����0
Ϙ� Xɶ�z;�a�Ȟ)�]����g�TD9Õ*jkc��F�A�Eh���P ��\�=u��NL�Ι�:Z����N*���ky㍻�\:rgg!.x��j��gU���S���՝���{�W��.�$B7TZ��(�.tg��k>̷MfC��H6��Å��%���";��^?/���;���FyFs�j��tJz�-˭��x��oS���N���p��2����s�"�Y��ld�zK}m���^�u�,�W�/
5{�F�f=t��oh;�5�j�<�2��7֔�K˜N�!7�,��q�<kP��gWiDSM���4yU�`R�C�d��b�9vT���N�p��Wq�.m�+����m�s�8ǉ>�0�U)J�%e����o�`��]{�T��{�}}���Ӆ�Hm�,�K*j7�*�p۳!��d�D�ٚ�v�U�i�H���c��rbr�Y��3�}��/O�m@������g��ҩ0(dCn�K�.���# 2o�ԬԞ�7�Ӿ��3a�A�|<z����Xce�esͱ��[5,�t�h���g0)�нWo%ԋ�F��H��!��V��b�����t`�k�p?���j�WY�r\�V��7+~pvY��yv_.wu҅o�g�2���}���8�ޫlW<0�X
vF��39�����f��t�we��1�:��6�����f��������7U\�v}�g�r�а���e�D�H�j��-g�Q�H;J�Kc��1��2���^�P�t�5�|�qP>�:\�y�(�2��t{D40u8���-�,3я>r��ȍ��j^�s���N�X9D��֤7�ڀ���)���`�kN�pie�>U��!���67vW�'����d���5�}�OQ] @���1�ۤ3�YQsW�s�}˵:�>p�w���r��q#���G:���z���%���ea�����m�D���D6�Y[�{�
`��錩X��]�f��X�(1�)+8^b(�D�.zl��ZڷJ{��$�B{�+���h�ïe�F�S��@��`�h��#�
O�e��ٸ^�.���*�M��Gt)]�k���-�Ks�������^m8�ԁ�˗�u!׷`t}:�^Ä٤B��ιR���udв�j/B��\$���-v�`���JYl��&��>��!�]v����%�_Rm4�BA0��K��w�e�����g^6��8S$5����JuȻd�c��é�ʎ�*�ò��f��C@ۀ����uh9��E���oG���Z���{�|�-��g.�;�''�9��:ЗBV�Qh�$�_!\ we��\�5j���j�����[�;A����WV���0m�L'^&��6��J�м�6jF�K���e�D=�	���s�r��#��ٍ��q!%uns��6T�z��J��/��ԩm�m��4bU�Q�EN�0�ф���H@<WnQ�RŹy!O���*Xur�Ռ��P���oW��St��t�(dڸ;��Uv8�6wn-zk/q|z�6D��Ⱥr�����+��w��U;פv��˶�o@0jU����Gk��eU�g�����nrꎲۦ4��<Q��7g:<ͥu�>���>��EM�ٶ��FǴ�;�\�@�l�׺��_T���m�햳�E�\����7���0܁�v���&�Vr����ªf��Y,�C.�X��jr�p��oӊ︄�ފ��"��s^��s�u&x�N�}q�9���̣}�֔W'R{F�xy�W�����su*3�٣OW�r��1���U�8�|�JN��w>�H��K�;���(�{5N�Ȍ<9��S�j^���x�܊�J��ڨ�gqX(#ns�����V�E�Դ��Q�mV���8t��p��"�ߡ�aά�;��?N��]��m-�A�(Z�]J��풮�m�Fk�W8��ޗu���p����Ԍ�qJ�fv.�oM�h��Svb��Zŷ��"��%b囋{0n���%2)DNZ[�W^��V]X7���K˚ܣ�`���KMN�������8a�Y�:WnG�K��N��[Hs�̦r�uH����tmL5����� 1�,������5.���hZU��PX�n���`�N��L+$��L�:��vA̼�M&rQ.���A�ƶP(Xi��A�]S�Z�>;��(Hx$&؝��-�6`�+E���o/�NY&�'��t�U�{�k�H���:B"���ݥ&VU
t����q�Z�
M�*�׻��^Տ�M�M�z�JM����W�J�x`|Zm��%A�J��T��U���TL:ُ����K�MGR��m�)�v�`�cs�Z��u���;�v,Q�J��;��wv��g`br��B*�)0��	MՔ�HY΄!��H)Q-ȡdUȳ	XY3-"!R"��9�!'6�F�#VQBG8\���Y�!Tr�"$�*m**�2�PYG(3"��(U����B+��P���D�H�͔&f��h��k��,"�**����H\)Afm-��(Y]S3%��9Ur
�E����	�L�f�*Μ��D\��"�1R#,�B�5�"�Vr�KDADG*��u,(��)E�
֠�Ñ���JVU�,�*�B�̪�J5(��QEG*�� Eʋ�3��&ʍ�% WT*���IR�ȳT�Pԫ�8E(F����Q��̳�J��B��jZ%�B�T�e�Da&�&�(��U�%RY4��QS+:�"�$(�
��� �8\�Us13$d\�*�˕��i@�J��"��j�
�+/��-�V�DJ�:��J_2�6{6�`����y�W\���v�5#I��·W԰����hV��Mȵ\�aQ��ԑ���}��|;�����wq<7�ͺ�ϊ�?:T
�c���2�:�������7?*����5�i���묞���#Y���24Z�p�' D���`�L�%8�xW*�/��ٙw�o�qf�k��"^E���A�2�����ݩ�UAU�D̡�ri���yIj���!ɮa� ��������U��uײ2xfq��
�U ��3�P�j���L��mh䈙���)�7L���)1��DrF��A�s��;�{��U��˲�ZeY�B7.{;�L�6��(�R_�^Kʼ�RtGDK�.��B-$�P���-�P/����寺b�R;4��<�*��c���`��5�����^�ᒺ]��;vL��A��ɡ�y�ν]Y�.d"$���	�6>��c@���c���]
�7��S�!�n����x�x�s[W7/�"�ϓ�s���)�H��h{m��v�\��}�fK&ɷ,:�n����ֵ�k�#�r��_�~�\������.g��gT	ˏ�9#F�O���8�Kn����$Ss'��x,��緘��E{Q�7XB8L�!Zͺ��;L������C�yJ�9�|P!*\aK��W<����s�rAQ�iN�s�R�%YWgeX��]-���n�[<�m�U�}m����$�"'�aU�#ފȻ����G�r�7�f�+�<e�X�4*g���i�5��2����m_�`���	c7ah���IӉ����fK���0u�n+�jx)���ŵE�#m�aI�Ei�Y���= ��n�Ky
��u�6�]7�p�O���:[�q졾v;�������U����#&�h�fZ����Ƹ��h
�G��EG��!���*%Ӛa��R���B�On��s�K:v��;�C�����?VWI� ��@#�dB�x��Ǭ%���⻌�kݏp�胹�LdM���!R��a�Gc��o�lhm�����Y1� �C�!?_$�x���k�1�Wu����W�x��Ll,k"�S�9:�И/]��}��b��j�ͦńz�+w�=�/ "@�6�(ؚ����	�0a�/��̝V�7����f/���]wNN��nf���#X�S(��jc�_ x����8���N^:3�ZG����ri���n-��[���2��Ϲ�����ɩ�
uDm��H�UI�~u_l�C^k�=a�x��hd[e��"��h��}�{)�n���^���b�>�}O�<��Y�^8-λt}K�����6���fOR���ͭ͛�k�w�y�u��m�<�GN�-�d�jw�\���֚��[p�	fc�$�zԿ{{����ȭ�Gd�(����v'��pw8��sH�n�˥�hmd���畇�;��sce��k}�W��ϫ�B��e�9ߓW�249�smә���7^#�c�*��U�z����H�x�IQL�K�|x�
��]�l4nRu2��d�#a�T���a���%n9㯽�AF�]��V��#֟�g@ �4��j�?@UDbN/�\^d̎�Q��Fqn>��*���B2F��PvX:�g�T>'&�U�+��v׮�B�|����HC�yi�!=|�o�����=��vN��y�}Zsx�@�8��e���A^�|�+��ώ5��tT��5�NS��صo����6���S�;)9�N����+��q��䎲pJٛ.]��cT%`�k��=K�	�ʦ�C.�q'KFx��%�b�.�t�����[�|�.&:%�p�fB2��_OL9{���չ;�m���FUd�K����F^�w��������ϛP�%	��q*���<6�[����g'k�Y�NA��U�ѵ�$Q$�b�)��Z���s����jI*�U�hW>K��ww��]��U�^�
�ҋ��0�����ײ�HF��]�yL�by�B�S�tRZuٰ��m_��4N�WQ=~VC>�tf��QîVX�r˰�p��O�W�D}�i��6�<GD܌�p&L� �jM+"z�b�c~���Ó9=�\� ���f��ܚ�}ܶ�#���:�+�h�r�:(�]��Z��-�*
�\�ɔU�cC\M8�:k\��<h"ʲn��Xc�wN�WgSF��x����^�P�t�K�<�7-T�^[���=�t�9׌��coz�ge��)a�1,����CבS���B�P���yvΖr{d.�T����Î���9Pʛ��*�p۳!�C�d�J���Wj����:��k:���*i%
摏v:=������&�L�eyr�Z�.��̖�U�s�s[�($�1����ɜPS���6��V>��yGGiq�59��w����R�ۚ�n#��\10������&Q��g�]���WK��
�/��WU��z��6<@b5kx�������!��H���������\Ŕ� �s�l����0ۖ��s<�[����b0�3]AN��������f�����p��\�v|��5�x/;Ӌ���mCu�2VjV�81;�Z�,�m�ړ��ն��3�>?m�����G-ZR�����6�����Fo<�mM�rW�<�(�L��6��������ª^�dg2S�y]r��$ �QK��Ɲ��w�_����꩙���~�&���fy]�>��8� ЗF*Ȅ��������X`ܔ�6��65���Ec=z�.;��j팳Q		��TK�j��<�ʖDf�5���M��a���\��&7���.L@vCF(pe�>X���*9��;�\7�~^�]�B�� mJ��֑�tQ�uO�]� |+��J9�3!�,���]����C/'��o��n���P�_��^��Y���@��Ę��(HH�:�C<�/�Z��@�5���#�Kdn��뮝������,�R��H!�۾!�<	N����%�Kj�u�� ���*i,��M��r-Ӹ2Um�;��$�}P'�ښ�UAU�3(GI��glY����7??���*���Ƒ.3_�;Hk�����dco�:ـDӣI�66�<6��Q�@.�n/@U����i�F�LRc'��䍺��0偌Y;�������P䌊ٖk�'������C�����	A�]�xB)GA�֒�}p�����f�K�g%�������<Sbۢ�RÀ��,Y�ӻ)�K>��A͠t�Q�U��.Y��$��52o���d��x��j��Y�Ѵ:�$8HɄ�Xq@׏o+j�t��g��V��..�i�}�G�D˸�ռ�Wo
ި�Nj)��:�	����~�����r���[����6O\�1��+��|��rF�T�%�[t�@�.�~�R7��nv���u���_���Nh�w]�cS�o��h�q+�1��ܱKi�H�٤2;hS�<N0lO�v�v�ܓ��s8��ض��8�i��1�����oa�;"^��|��uT~}�r!e@���M\�\�^�ÖZO؋AKW�do��:���(���!�o�[�Fp��k�rY�@J��;�\o�O�L��������#�/�PK���8,�c�a��+'�ťE�"r�&�ͥ2�-�H����ո��x�(��u�>��hd��1	g���]n)��^�sQ���쓛�AF�=��L���٘l&9D[�-iY>��(
�?w�1p�����ѐ&�䲳Wq�x�O��9�~a��ߞ�7=�d����^�	1��4�
X�76�2��Rb�%sG���Jy�
�ei|�uM�yYB���p�ݒ?a]�����΁d�y�KLI-(��X~�)�X��7	̷�v����m�z8�[�v��*�#�V��v�z6��jTf��^|�;��V��4���������>�+��,2�d��zq�S����P�y��f�دr����D隳&�����Ͼ�ꯪ��*A����, ���>P�PS���x�.��#V5�y�$b��'�`Lqz򥶭�I�\Փ�ݛ=�OA�Bl]�	��)ؐ�}=!0���K��:��b���pul��-���_=}����JCK=��P|�����5D�Lg�/�xn�N^C�?q해�M�����0�qR)c��(�G�q�Sq>hR��\Pf3���Vc���2�#�Q�'����v��(;i�1k&��V	S�0l}p���W���dV �Έ���#֪�r�Lvpgodui6��ԇX�;Y�
`��R�W�3C��7�t�x=C�'"^��>&>���S�W�݉_dy�YX�p�#��s)YCn��Ġ����=����-̚��$���β����֜��ħ�A^τφ/����eԷИv��N,��z#q|����qä�*��3���)�어O�jr�l5��ƍ��[c�!���L����s�^>��蟣l�������:��Ưo���*�}�xg���t_0<:Lk�|n蹀�;q��b�xȓN�7m��_7`p[Y����x~�c��H��� s�oo�"�C\v6E)9jGf�s�[�6������)li��Z�[�X:��{}����R'��	Ov^��,4�VC��^sx�\��OL7J��oj�.�Y[�bG�}]���Z�=�ɟn�*v�y��E;L�W��Ȅ���q�3"3�y@+���g:�d��� �=&)�>{�{>��܈uط�M���:5���\�=H��2�dL�&ֺ�x���9���q����E�p���,�ZC��:a����<ko��s���%}���ݐ!� u]3R�à�=*����Ec#a�26za�uº��gm��,�����qD�>���u(�ઉ��x���������n�ӓ;5C�D�C��w����Ǘv���d@�>�u
a\D�.%$uE |k���ԧ�n�f��-ؽ˃�{4��V��g����c��knB}�t�ς��}Ƈ�"�s���Jy�)��NseŪ�w��iy!N�5[9=)5jTC�h�#e�p۾�ǯ"$c��$c�a<R��wȵ���l~��Xǔ�6���2�㊨`ݙ~�/�,p�s|�-ם��;[�7ӟoq�5A�q�6=3&�h��d���DbO��M\	����̗�}QB�����ã2SS�����[@M�3�@9r�b���v)����o���+��2]��B�����l
�o���5��[��'�a��u+0�Fa\��/�u���c��퓰��H[N^Rt����x�ԅ��uJ�ź�d�a�}t;�m���_�����ޔ���p�3��`�uu0V9��]��ώ���ۮ���Ԡͽ��21�%1z{﷒?h��F�o;A�h3'�r���=7q_�Kt�˳Lr��g+�yaOKJ���n�[��7�6rrnh�7P?xՆ�r�^��Ū�a��k�$v �#�x�f�Ü�T�X��n�������o��˩���Z-�vv&N��t�M�jrQ�?�Gƺ�h�P�f���A�)�]X��0^��
r����TA�ǟ����Ip1N�ӪC��QN%d�,j��cϜ��ޚ��[�ׯ_SQ�YLzyb>I&������^���	��s��pv�c���*&,t�_C�:X}.s<��}���W�C��.��u��*��`<~	�n@j����D�bwE�nXJ�{+�~|��S��%����L�+<~t�C�Lep$$]T����ۿ����\�c�f�maz����쵴Ї�`���
��͌�V�ئl�];���n��(Ŕ�(��N�Et"§!U����3Z8mu�Bf3�P2�jH8*!��C�%)FJb���roq�2ںjc�I�?=��K�����L�YE��>���\�fm�$BQ<�1�( �a�<��f5n1@�j�gn׋�x��n�vl�L#|��#���ic�N�ֻ;P3��1���[�pd�*�dw7jH
ʽ�/6�f	�;d����'�I�vE�}� !�����}CWC۴�����}�;Hk��ƺ����3X&+�������;���+޼ع-ذG11�W���:�]���搸��q�R���A�r*����5��:�y�7�H�z�+�C�CH&��U�Ƽ�g�����.ĸ��k�}�-TU�&�5�:����!}�����+O� ds��D�����V�]��)r�$�4O'�����q���"y�9��I��/ K�X>{�h����]7�O�)�[�ֳ��/�=�����̴.��>�߅^w��]������L:����B&<KVoOHm��4&}G����&�l�N���}���H��\%"29e����L���E?f�f^5%�f�D�u��nX��TI�o��s8W���!���:�CإVX`tX�`��7�w�Y�E�y�	qh�����|�D�����GZ\1��:K����R������V�ު��o�����,��x�0�*�����͑�,k&��Uz����͹C��:�Ѭ[���1� w[�����p���{ך�8�|&f��va�⎅�_R�*�R�b%���:�}��ʽ
�T���G)!���/���������Kyb�{���}�۰P�B���ˬ��V�c���u���z�%�<���SVO(��&h�>��x�|K��]�
3C�y�I({w�Z��_H�l[���T��/��J�b����w�Ȃ=|�LC�g�\t�`�X�K�"�R�.\]y#cc����j�>��M���|�1��8�J�\�畷n�01.r�U�U�'&T���Ԧa�N]��y�p.�Ђ^Ru��Ɋn����f���k��\�֒�K�;��u�%��1	t��{�#n-[��iA0�z�ЉB7eҳ��^�i��cv�v�N����7��ת��Y��+q��������l�=��^�!�F��RH��T;.�7��̦���5��:�!�|Uv�3k�3C)����, ����ot�å�jv�zҺ�U�U�����@i��U���n+;�%���]�ڶ#\�l�D�up(�R�� -)�myh���<��\�abT�n:Ee/k��ަf޺�Ct�gZ�Ж]��kTj���n6V�yi��[�Gsc�����N�ab�5
=͘���W�k����3�3}����[��E�Xv��m�-��7!WoX{c&J�3E�c������d���q��(�,���=�d� 4����w�كV?�s���7}%�z�G�l�Vbʹڪe�W��ڝw1]�qp��P�0�{Xk�VK�]�	�U��l��	veQHp�(q��&�h�:������Z�ڽ�e;�G'v��׬S��'%x3p��s�kk#�����5���l�ʋ�̂6s��.x+�4��1W�>lm:����q�i$��_gS�.�Ȉ�!8�ݥRGQYʗQa�w]oh����q-=/���9P�T5o9�+�b�f��Vq!ˍ�(f��7�6�	`� m�'�8���W�
R]8���r��k���P�5�3îs{H|M�y�C�Voz����-�@�w{����@�c�XflՋ#�b���T�	z�-C��R��5��VY�ײ�^QGc����'b�jc�.�f�ڑ����j������qY �����=R�u�^hӁ��y��(�P*�.�+�3�/7�6��i�5��X��5м0���Ů؎��QCu���<�B_w�1����fBvF1�����7���z�:5b}�e���QYO"�fƃk�{ކ�s��L��Տ�J�ckve��E��BsǷ���tW{U�E}��.�>G4Vl���n������������欹A�_���,ޫ��ޛ6�x�r�·`�e�w&��uy����Xv覮@|P"���QI52�g*�D0����(�UQ��%NDQEU˙-2��)%R�(�YE�$Y0��2�"��j,"���UTQ2���V!J��Dj�J"9�UE�Y%�M�%I�D�2�(��8UJ*�Q.Ut�Qr#�UEt3�Uh�t��91iUV���t�!�QrQ
d�]DL(��)S��*�Q&F�EQY`W9QU�,�U�h�1�\��Z�\�9�"�
�ML����*���h�*��PfVaJ�*�3S	f!��3
T"��uQHS9��u\�D*�*��er��M4�UUkJF�������")R�EP�,�#�PGT
eÙ	3:h!2+��UAp�
�P.)r3���V��&gU(9�ȓ)˿��;����wxOyQ�*�\�4̙w���N�uŢ�� ��t�x��(Т��i�mN�Mv4����w򾪪����SoG,�#�Z��ۣ1���~�8��
������<-��Mo1ǝ��²:�I��k��������=Cc�J�t�t�;��[���Gn�ϰD�+�x�e�\yP�xb��89k�/��r�w1�R����9����]��|�'�(pB !W��[eÀ]�d�<�U}���hN��Y�س�}�~j�ϨK�_��W,�+���ov�w`�޻��V��h��
cGq�]y<B��-
`��*�rxlCt&]�s�ey_�SW�����$��C�x�R��b�A�_�J��ƶ]��3���)�ֿ�k{���O0��}�Ӻ����m���P|�����5�蘏�9�S�+__
��;�e�0z�*?S�w�ʝ�M`b&q���СZ��!P.�C����T�}P�rXm�8Q���SJԬ�e`�9�0l}i+`=���'�`gy���x��Giy�e^X��th[���ز����ʖ��,�1p��s�����̹�����z�^��?���U�b�^O��&��i�co]��O�6��bP�=g��經����ң5ᾔ�I�l�В�G��׾=�-��X�`���z�v�Z�3�qwd7-qS](w
��ݶ�M�V5j��X�r%�t����}�|3n6�_'��}E�n�-�4l�������l�Ԃ��<�b��QXn���p�N�]����Ԏ�(moxӌ�,qt�j��^fu׮��s������6�p�i1���`*��* �뷊����Dy�+��r�	�R��6��˪���:5��b���3�
�R��wƚ/:_I��qe��l�l�6��������{�)jxtu��L�7�7yW������U���<��N@Ff�˓3P��b�m'�NS���W��M�sf�R�P?+�.����5��`�P��-����v�̵�I��1��Л}E�=��,���rFW�{.�U�[=l���{"�9��Q����g�Q!\�!lA���r���bSV��g�Z�"\b8�@�(��'\�)��% ���Ƽ$�G������[#a�2&*39]�S87�����v��X3�_K��o�P`Ò�
��I��d�$>�]w�m��ڨtG}gp�u������l�ڡ�`�>ۇP�"x� I
��$:�J{��o+מ�Lm�vP4�gk���¢�d`U�+��=�mZ�]�
��P�y��[�����fה��"]�nL���J6)�w>�{]�jc��"�1�� Ty���S��
�Z�o���aF��M#19���7xz�%�A�j�ݘ4�N�\�������Ʃ�:�<����R��C���9�Ο��@ϟ<�#"i���*���pΠ��[��6���s�Xq�P�s��Fș鸄��;��!�d�;����|��U�A�rUBr�q5.Q����Y����3eIG)�o~K>sC*n;
�`\6��ni�ں�n�iV��[��zs�N�L>އ
�E�~T�Y��}��,OfC�z=��5^*L
�I���]_<��Yl	4$3�U��Uq�����=����}��Ǝ�:^]t(V���t�]H�>�t"z0^!�������e�;��t��:5�8�zMsW�̺�
�j��l��^#f��~�{|����}[gO�o��^�U�YM��#�^�YI��I��U�+a���=��L������f�Ü�N���n�X���}i��'1sD9������:�.�y�q���Y�Q�?�+U��&mPU���pNQw���k5�ڳ1�����	Oq@�\�2o��.
�chЇ����D+%��eM*eӰ�ȣ#��9��<���}�>r���D�������~[�G�� �����^^�Eݑ��WjD�{o�ne��؅�m�VP����s��[��e������H���珑�gV��X[��\�,��T���w��4֡ޓ�i՛���ܳ�\v�0�9�s1dd�x
��eXal*~�ﾏ���%JD�f�B>�r�i��ә���]K<F:���i�.+:|����Hgt��P���3�}U�{�/y���^��0�ȃ��@�WU���uS�܃�[N��{'K'��yi�q�?c2�N�΢X�md3�+X��X�>$�W ��d$�����y��*nh�8�]�OD�N�3�{g��6=���DF�U��uu/�h�T>��Ǽ}48ɚڶ�z�8��ؖ1��L���B�2���0��ȅ[l��nԐ��ME�)�S�*�R3�r_#�\ k��Q���]�~DVB�>N�����D�Uu�g�K�-V�g7������+6g�L�$`�� hw��5��ݨWx��ֺ��j��cޠxT(\�Iب��fsex��+�C��GK�)T�Џ��*���: �Z-][��y|�-t�Į���
���Pϓ��x����=&x�X~��i��� �]�0�������tM��o�Pg���O�*rS�{����X>V�֯�]1�-O#�sdm%�Y�W��t6����<����e�nzL>��<��;�k����8�Zh6�ta���Ũo:��*�2�e�I�F��gy ����KΎ	
=w�����2ڤC���Ҥ۬h������Kq��)̏�ݱ+&T1Sߙ�,�@(�>����Óӥ=y�j�|�YFa��zvjÞ����jw,R�s�8\7Qrj��s\���Cg7��՜$M�"B�c w\�HT�Ld����ÎD�x%na��^\�Eni��{�p�.�g.U�l)!�d��T�s8W���~2���i��U� a�=�}q���7'�{�wY]���_E=���B��O��:����;9��5��L��rRj;45�y�l��h�6#�Lp<
���W�O�&�\-��𶗅ɯ���{���\��N	W6�o%o��������ct�;��2֊�!�C��1��c_*���Qd�'��0�	�t��A��f,Y�~��t�"�}bWd7�>·ZRMy�+�,%+���� O�<��l���m�4pв=�����#�X��񪝚ؙ���X�l6_���6,߳��mא|�ԏ �*�C!Rɧ�/̫�4�n���������y�e�E��X�Z��W�`�����f:G����>�	����%dpI>��㍺;/�J��n��Ч����K�;����V&��ʍ�ͬ����7��z>�N�\չ��o�h���bp�~u�Mv�O܁����k8����&�
Ϣ\^M����y�}��L��1m��a���j�ꁴS5��r�:�37���a&�,�{�{�h���6b�q]����@"�Lɰ��z�R��Z�؎ ff����ɷ�g��9R�V�8�����B�-�B�)�z��5g��$�}��ϣ=s�X����y��>`��%L��2^ؘٚ�;�u�L@�ۼ+E�]V���} �� �lxy�e���^�*���������W�3�f\�t�x5;W9P����n��65cz��<jx},� �~<'��iH�c�8:QZa�=��OW�Gp��9��h��$�0s���o����n*���v�������Z��a[�y57Ww�Mg��JN����H;J_v��o������\��g�t���ۘ�Kf��j8�b�����=&#o���Ñ����p�m�7�u��'��gb����y:⎢�R-�SL�R;�	�u�����伢>v�Ko}H��!uѥu���[�Ž_[M_��+����OJ뭘H�J��{�C��Nl�z��/+r�"�]̜O�s|����i�۽S�'wc���3f˿fмͭB�RyD����^��'ա�`�)��=-+�]p�q�s�b{�.�Ez��.��c.�+��thS�=���I��%��`U���G��}�z�C�3�_��˯�5
��Q+����Kx~}-�Gϛ6�߬�1��e�ߝ�xR�ެ�9wʄ���͝jl܎{����4Y�
#4q\��=��?}���s��%e���I,_�����e.�wgi����I�4=��OZ��鿞���+��T~&�8K��Y*�EI���r�ot�����G'���9�_͞���u�b��~J�GQf5�c�>'�T��׵G���
�}�r��z�&��e�c\����������/�=��+�z��{j݊�Y�z���S�s!�e��8�;�V��҉��/7�<^�x���X*��|me��J�^�MX��v��W�5'�:���zq]c�t���z&��Q8��^;��{k�o-��^������PTW$�1oq�q���O[{w�=q���7;�=ǻ!��6U�J���լa� ���j���"�|�O9��L��2�v�ۮ�2���iu���L��C��t��jn�t <�+kB��n�X}(���Nk�z����wC�������n�»����Sn��jn��*+�6SY�1�����@�����2��6���ǉS����w&���+���2K�j�f�؎�S�����g�ۧ��yE^�� *zƷ�d{��>7��-���j
�����*�:_�Aob���&����(�3p-��=e��S���%'�{�3���1��w�:���lq��tn�CY��:��E��<){���;���.���%���)��,W=�������%Z�iS�uݓ�tz�u��4V}W-)'q��E4�ꆈy.�P�/�n�~u6Y"�d�Wos��]�9½
����'�̵���������"�#��s�4Z��O��X�b��y�;�����I�C\��fr:�C��]ԇ�*��j�sU&��Z>�p��7ͭ�CM��j�t�S��l��cciL����)bf��#kx8�&�#
n]1ȼ(i�\g��X���J�)y�EZ�ؾ�D^޵Z���dɭm�F�� �^:��ˈ�	�3C���4:;l9;"�����\M��KP4ޥ1�פG2������ۃ.s(L�[7�q�}��C����T�i3s8c��u�7�}��J�="YC9�~��I?�}�}�}^�D��ϙ��>Ժ-���D�W���f�=�'sҼ��d�]������3�]�\1�Z���jh�H.�NTί��g�f��֭ʺE퍇�ST�8ɴ̈́��Sq���bs�*z�\���*�<���v�w�썮�Զya�����������s�5�Ms�k(��%ˈ�ZowKN���m�;_gU�J�jp�Q�'�ۃg�����;��-<i �s���Ӻ�+�������j���>i�GK9�O�q�X'_��le�N퇕>�q�������QGYqu;@�|��59��(��3:Ggsmq/I�����ȉn�m�(f�kX6NhN��X��ko#�t�[���d#��'�N�rM��<���cbca,�i࠸��m`݂��N�7��o[O�S,���{�3�n�c��Mk���)�Df֓�"J ���<�)��Ue4v�A���[�!-�9�2P�����5VdqYB�vZe캼�t��-�_f���"����`0sxֽ�<9ܮjr��P�k��뎀&�x��X����m�{W7�K�W`G���菢>��Z)7�o������IZ�x7���ϟJ��ٽ�{P�~�5�]j����ٜs���wġ),;�k��R{�Ե���}�,�z�k8i�##��sr��?3A@�Rsq<�5�?d�^�7��\���{�>g�W|t�s�z�ۤ*�G�h9��s�kT�E�q���te�]�It��\^1����l���:b�BUA�J:d�Y�dQ���T� �����������-(a�nq�s�h�!����Ңx�q�}�y)ڭǛ��%'����a3b�N^0�D!�������5T�
�����$�l��/m[6���E��E��i��-�ސ\s3U����x���'�K��58����q�n>�\�'�V�d��{ն �ո�5�//���6������^�958�n��{pmu��zW��جPʝ�V0vE�q�� �]���Ab���ox���}]���������/���;�3ݨ�WgC���ڣ���K�"�DY�"�]����jݙ&���Ӭ4
��*�V�]��a0��'A�i�Z�t���m�"լ�u��Y�N(5��2�"\�f��ϡ΋[�hs]��p��.:]7i��nT��:�c�o�nKF��S+��T�u5��AgR�����WY�#BU�(:
��c(9YZѡ��^�8v�]SC��]���B�ڹ��7Y�yҧ1�by��SFp/�2�qC=r���8�۳�Ֆ��G1o���c�sӈ�x��9��������jY�'�ܲùmR��jS�xޞE�#~��}��5���9Q��G�K.�5�$%$"��w�2���s��IQ� ޺Q:��j"�eD{�.ε5����`��':�h����T�N����T7��(F�uU2���ݢ����l۽���ߑ���j�{SRӮ�h���n���^�諡�H�o#�=LI��Q�o);�������	7�Z�Ҿ�r��h�������@f�����:F��XMd��`��T{���Y�̴���j�T�8a���Ņ��Ʒ�j�	F��yu]�.M��+�n"��P5j�\�+.u���&�=D�9+uͶ��ǳ��0�㒸�*����R�����;�X�JI���ak(axwu��B�V ��f�m�)+}Z�otҫ{-�>�5ra�����zκ�� #x$�	�#��8�]��PQ�B*f����c材ncm��VB�<9��M�"]�gj�o-�^�
��>:;�$��cF��BJ��JJ�F^7��N���hg%捫O���Wc�u*�Ϭ+Uw0����M��O.�A�M)�ˤ�v �{lּ�S�'���w���t�\�&.��ڎj���u=3%;8D` �҃���,M9z��GSd�|*�r�N�kMJw{ϙ'z�z:a�beȷ��5��3���EqO�Y:��dSW]�)]�5�]I��ŔcK���eD�9��}��nq�ܷ�jٝ�ϢE�4�8i��6�<�c�\t�a��LM�J�k�Вi�t��昄�Meٲ�A����"<G]f6N��ٹ��n	ȝ��2�E'��'Od�y�˛}1�hλ8,�t+v�Լ�j��1��ƞ�6[ۘڦ�ozr]2�]�B�'��J5�)@M^��跇]���eꛒ�9�vq��V��,���@�sEZC~Q�;���o,���>���*���h�<N�I;A/]�#���T���#�2�m)|M*rl���0TƳ-��;Քˁj��➯��*�!�[j��k5�L#:K
�QX�� _�Z��&�-Y�^�p�[�2O�PƳQ6LW��Y�,J��[�f|��N�.�j
��EL�ݜ�Dqn_u9R�����Ͽt�D~��
���PE�X��D
*�T�GN�"Q���U5(����I�F���E�M0��,���%����(XPEΩ\��'H.QQ���U�EˑFe%I���ap���Uk+�UFI��GI*��&QD���.�B��ED��UD��V�U��VaUTV�(�TEE2�feZȊ�D����J��U��9r(*�l�iHY�Q�MJ�9G
#���
+X��h�FZvW*���-B9P�E�t�B��_��2�I�P��*� �U7"�q�,��aZ��r.-"�EA4��%Z��:l����\�hȻ��.^%�E�T*�"��%bDQDQ�Z؁�&Rs���*�"����w���#��3PU���}M�.|�b�����
g,)�|�b-D�+������`3ɴ�u`�X�X�=:������ZY��{}߁���n;���q�n� ���o(w�[}�_ەl+�v�P��)s�N�
y����(sR�������G>7x6�ݰ���F8\v�8�a۽qN���:�H�!�Ƒ��O���G\����H|Y�x1�!�<�1�_Hj���BY=Md�r����i���eT���'�������x��Ԃ�����%Z�k#�z�[÷�����:Y���%�õs��&��s=P��%'�,%J�f0J5�'W>��q����z�������_\=+��蛓Q�eE�,_��\Qֺ�'�Z�H�OV�7L�%��gK�3��Wr����������;\�I��V���g��q��2q�I�s��e�c�1P�� ��!Hg-��Z>8�\�Ư�ڇ+��z�&�0̼�5�ob�M
+�V��Nܳ��3����=��J�T�R����.	m8�I���o ��ה;ݰC\�Ć�v��rfv�Sٌ?x$n�x1yw<�q*sz�r�GF�̔w��nTQ�)w&sJP��3���t�X�kQm�7As�9��嫀�O��U�Ub�9=Ox���;�Lt�@|���=Y�)��J�6̱*z��]NQ�hf�{����\OlWΐOTHN�쮈�/� �֋�)�}ݮ]	w���J*�2xȸm�<�
ێz&��S��^;��t�Ʀ�%N/�ϡi6�h��N4����M�f�cq:�R�z2㜚��n'u^��s����>�oUyv��緋Q�x�!*}���5������W�/T�Q�,��?I����E=�-����f������4]f�>4{�)��(U�)B]�R	���W���4���Pu�Ynv��9�l� �p��ݢ�;ӣ�ܝ�q<{�to��d�ܚ�J���`����y���-,�w��Zpw=UQ�U@�:G��ޡ�f���]vHV�u���{v�'�\-��l��ǰGU�w��}��톅&I�W��s�8���%T��(�0��B%�ۢ�7Oٵ�k�y���;�cjf�È���T��k"����U�uԻ��0��Tr�<".u�)����[��tΧ/0��8."0pV���r���Ym=����Ck.��V���ꪯ���vy�ڷ磳�n��o���C�|�zh߹�$�,������.����{�{0�-]�v��'�sGb�6�M>�Ȯ���<i�u��.�}�:�M��kT�+����'�{~l��G7ł%���?&l�����!����U.G�.���^�!����&����2�����3�h��qö[{���ni+��3W��߈N�m�*L���k|Z�B��m�-�9e��jj��V��r�E��l.��|���1.Ĵ�F&���%̹e3b�NE�n9��ڥ�/)�Yf,�+����Ȱ��[�X���[��˫#yr5k�v/�N��W�ȿ��[��7^�ڽ�}=�̈́�8�]�;���Ϗ�_^u�Ȅ��F�-w:,i |F�v����*/�"/�W�-���q;��W�c7���܃��v�\7[q
�򣾣��L@��RnU����%���\w�l����:wp0^���p���o^�9t���*nn���� �n��������{�{{�/�_�n��W����*��w�k�9r�X-4��L±�R�����Sh�Eb����p�R�ò���wFeuj���菢4�<WV��H���7&����he���*���^U���Ջ������u��;�Z����i�!����^���s$ڑ��m+���*uN5�vO6��QK0�u��H�9M2��O�����;2Wu=�s�z�kp�v-�N�����J1�oe���9L��3�X3MD/T�:1�⊝Y��+�Ų�#}v�b�k87��[����m=�<��;`��*��s��]|	e]��_Tس~���j�/�RY����Y�U�vå���Ws��q��5����(����u��L�N3��<.�:E3�)mV��'�!��=cm�����s)t�pMm�%͡M�Rs���;�1�{�8t�Ȇ7�s�<�n����_��"zz�Þm9�!c���h�*{z�9m>3�	����k��#U�Qu��{���j����ik�"�~k&^q���@�GP�P�5$��Z�3u���9�S��%��ud��`��֕6���+;']	�vv8$���L�����17ӹ��A?�b�F9�n��MĖ�ZV�U�:�7��ʅ�U����D}o��e�՛<v�Wl�a)���LظI9y8�!�'ar�XgR�T;u'�G�:%�)u_Ҳ��܍���#yu���&�^'$��٢���|������m�5�j1��w�ݸ�\��םx�O�M��@����j���i���/���]��9���J���r>Ѯ�1�k�[���˵��	�i�])����T�n/�0�2x�eQ�Z�)�^J=��M3:���E�T[�����f��;x6ʝ�n����c�[U�|Qyg�"��Q�2)�"�g)���wP�͛�g�~cR����-�KvT�wN��(K>��������o��i��Ul�q���h�Hȼ�6�`۳3�
��U�d)WT�:�l��b�6��Ns�)oU�n?���E4��srk�zT\K*℞,�+�Y��O���w�]#�У&��Yg���Ű& ���(�֨�p����vw�z#᫔v���y������Q�\��ں]�-w
��R�×��y���;�J�f\b�,Z{Y�h*	��ݽ5R����ںJ���7j�{v��z�����bCE��U��'��k�K�zW`Ģ���!@�Ic �lS��/��֍I�z������l��L�D%��gO���d�W�3��xD$�ʔկ#���1�6�m�^�!�s<]4��}���z�0�Np�
o�d��I\�G����Rf[���E��!����id0̷8�E[�f�sg~|�����pp��7#�:r�Vm��S��S�Qc銉��f���Ijs�>��J��d)��	��r�.��/k�]�{�` �̺�d��j�ֿ�V/r/��sR3c��*N���x��f�.��Dq[��D��p��f��q8A�7���=q޸mt�u��e8�ל���o�?k��j�Og����׏���s[��޽��4ҵڟ���sle�}=}�������/ *z���5���M��Þ�W��RG=sت{�>>����ڼ�I@�^uX��Z����+v�j�:X�g�w]d��>��:���$%*R�����
��8B�{:j%SOzr�{y+6�8�dI=c�2�P���K��5ƭ��D;�n�F&4o�G�L�^���/�DG�C����Vס^����-|:s�k]�,gR���==�S��J�>�i�x�nƽɦ~~O~��m�;*�x�8�\���p��qY��T�1Mr�'����$��i��3��r�::����\O,����w�#aU�[ښXI�*&�Й������9M3�3��ke��)Z�g�Lq*@37G?Z����	%û�ٺ���e�ϟK�m>��om�X2����|Ǹ���뢤nXw���y��4u���@�g:br�B�u:��x���O/�0�DJ]7<Z�CM��i�ICY���F��VN�Y�D�ǝ��2�^�2�����/�r)�E�4��=��_0��G�3�(�V��3��N�m�[���I\�	����ݰ�C5�v$:�J�.�q����-1�^B
��C�"Aw��@�O,��m��F�f
ƻf���c��ME�w$�m�厫���ld+�G�s�+aw����o��2���X*Y�1Χa��}��t��Vk�J�4z��&�uee����^j
��"3�5�bR�y�]��n����+6�@��OR�g�G���̝u�^4wUeq��2��r��͋I9	��Pخx&���}A���A���^�����4���}Y˭Ņ;�0~m��yH^*$(���b'�{ճa��~5jn}m��:����}y׍ ��p�G=��6J77Z��}7���3؂�r�)���+�,�Ϗ'y�^������eXճ�Y����0Z�J䋩�����0�s7��=���Q���g�^U�&��y���v^��s��!���k���6�is��T��5{!�bz�i�^��;��\�*�N�7���E�>4��'����r]BY:V����/NoLֽb=��9�W8K'��ӉM��Kq4�E2��ۦʓp�7e��w�k�2���Iy@���t�b������C�]Σm���� u���AJFw8����2h(��UL���ز	�w�i� �(F�j�m'*�t3)d7"gtu	u�y���2׉���o��n״�Ƽo��V��߄���zr���Gۚp�"�o*���Z�ŧ��N]7�]TL���S�]��':f�8*'����n�ͺܕ*�{}�b�y���5����ɾ>�'��*J�nMD��
JNn"y%��Owh˔`{�]�ਗ��Q�E���g���oX�t�|��?_���H�H�a��8H)�]�����<U4��4��ٿ�c����Ԥ��o�}KHT�����7/�O��Y/��񞴋X�2�r����hVʛ��e��P���dw��z��L��G�>%;�T�Lؿ�N^0�7��5/mR/Q-Z]7��`�g�$�r�3�l���]h�y	���«qE�ZЗz���<�C��e/x�k*�[|^�=��\��]�R]�L�^��e�q�����lvC}w���&�'��WX��sf�6;0���8�L�ԲqJ)'�e�Oq'��������^�S�q5V�H�v���N�*���+qm渧JS��U�/����������|om��vU��̧�|���=A���ӄ��%L�=��i�fލby���fT��tY��R
isC4e�V�xk[���>5:�@]DD[�ƶ���/����V�0v5F��]���lɻ0�/�*EV�P��A�.e�W�fՓoJVz�MfVZ<��pꟾ��O��[��S�z���VV�Dӆs��Q�<��Ǖ#�Цh	�E�|������Q��OC�$�y�0z"�BY=MF�&�{yP%���x�P�y� �W/3@�����ڷ�}��)WE68΄૆�M�$�ea7�z�)K_7�������b*��=F��:G����ttLf��y�j9��B�ui���Z�g{�s��&�����WRWxKEz��|�[�[�_�4�'|�"�3�k\�ft��X�蛕s� t�:ǁ�R��S�CNi���8�.d��Qo>��K�4���4l��t�'�W�����5�OH�WU�"�~CU��=i4�f]3`���<��-�\��q�t\<b�`ĥ�=2��G� ��S�:�!���P��SU���V|ÎylT'�p���m��ۊ��/U= ��^FP5�ٝLp�B�[W5���<9��3%��	Uoe􃨥�mc�#/���	�.��d����ǧ�Rs`�;n�Y�:��Q��zF�'u6��㴂@���!��r*|f�J�敪k�Lr߸�Y//Q��6��:���16)��k���,�E@�:��xZE�uj�W!ed(��jfj���l���{ق��WD.�;lOBW��'V���+��n��ZR Ӈ�y-[堝�*7�H�lc�'W ��
��{U�"v�	�����Ԋ�km���ǭ=Z$W��n��NW�fn��r�yՔ�edjۥ5d5����}��n�gÏZ�@%g���9>�����3�enD��֦���f�j�g��P�����_H���T��*���OM�b���7K�HQ�ʹ��o�f��r=�K��M�0%0mQ�ly��r�:�	���Tv��J�7}]�*ڳX9�[����H�03�%�Py��#��X�P����t1���8r��2�P���6��m92��w�J�֧LGX��dn����X�C�,֩L�G�� ja?d�4kz�ă��C�۠�n���۠94��h��w(��aoJ�ރ��:րG>d��k
�v[�.�]�o�j��Ht�}*�or�ɖ���@��ؒ�_á�f���+6�6w�@ ��NݷrSw@&�m��9Dq�Q�S`=yb�[��k�,*r ͤ�ڮ��#�h�2s��"��ѹ�9�`n	��=]l��6"�K��Rq�P;�[�e�}��q�+��Rޭ{C�(��;Ǚ�Ӗ*l��A`60.�7a�2�LkV��as���"M\F��\�G�r�m
؜<7�� �^��z�we#8TW�1學wG�Kr�&�ͷϑ��ܺ�|�	J��1�������:�ѐu�r3Y.j�ƌ�}�s@V�E=�t��	��M�mj�� ���K7\���p�f�Sn>���V����9,V��r*�ݼ�ǜ���fX�|�@�����f�Z�����\�F�+�9�8(]��5�i����*H�����Q[��݀֫S��Π��r>�/~�j��ȉۋ�LOy��L�j�T���k�z̢�E�3E���p��G:�]�)Cuk��U(5�-l'w��yu���Hքm�V����kp+Vg[X�����2��sl��Cb�6����7QCۡ[�@V7&�x�$L�p -U��ˮ�����0�;f�����/P��G�3�RXB//^V�M�*4��N]���-Nɸ7+;L��f�<�l^�6���µa�9�Y�
塚�N�f���r���jE�&����]����L��%鹘�1��u�\��� $țʄv��1qf����8���#[ez��\�Xi�"
�;���nl�u���-���|�:ʾ(�V��nJAr��q�D4L��y���j�#ox*��$��6�*�udkV�z�PU�gʄ�8�˅r��eEEʳdr�LL�is\x�����(Э�I"��\��)�^*�a�9sH�<�*D���	8QIYuK�5"L;�H���!�q���T	��r��	Ɲ����Ï(W&hRgq��UQ�jY
��.���Ȋ8�es��Q<x�^'9�Ey
"
*��VJ�Ywp ��:兕UQt��g3�q�ur� �(H/g:HAr�
.��Q�˂Nr\�Pq"�	��9B�9��E
t*"�Pˇ%bT\*�˜%PN8���%�$\�҂"�ye���TEQ!$P���9Q�9A��1*\��Qs6E�e��xȣR*�����TUN2����(���Qet�E��F\)ǂ�qh$5Z�90��B��VF+"�.�$9NG��GIf�iUd.$�ND�"8DD�܂�H9U9I:$���D�����]]���w*cN5���}��<�1OW���t��W'ʹv�hV2�(\�\z��r�⼸���Ӆ��Q���\�6&�{��D��c�5b�Ĝ���s�+n9蚂��.�x�e5[_L�LJ�ɠq�d�O�f��oD�58c�ކ��9���'k�<�d�E��%i�{����������^<���}��5��N������i�T�����	�;��f7V�X��ê׬�����%��+St����:%�%�B�.8�����텕ʸ�����}+)�w�=��N�'����J�c�r\p�7��[��T�7��W(|�/Vgf��X[(�ʥ�{�oT[Me3��r��::�g� �����%��;�m�k���!����{-�6�ϩ�ru�n����k7���Φ�N{�u��r�ٕ��C*���!�krK�m>�h��9Y��!���77�Q�4��3��I3�FXw�U�:Os�k�,�r�s/���1c��9���1�n��ɉ	qch���=uNv���]{��Wk�|��/��͖xQ����@	�����)ķ�a�Q�4N˭o�t�r��C7R�3w!ক=��cBBŷ�:�i����\���V�|�,PГ��G�oP��E��;�O��m�S�<��-b�6�����$ے���7]��7�l�|t�����
e?%Q.e.��^/�������tZj�R驧���͹ܖ�´Є�4��H	�}�u��͝��=�X�Y(�K@��|g�,ٗ�k��lR�&����`Ν�`rJ^֧�~�˧j�{�,4ߔnY�3b�I9��x��}����*�j�cH}�a�$햪��\�]����7�cyu�7��@�p��n'�2.���s��R"���/���N.��t�=۪{�~�V�H=������@�8�����h�yo=���)�f�Nϭ�¼nil�Oaˬ���9Bv��9!��l���Co���O���Gӻa�D�f��׮=?�� �;�\���Iq�T=e�E�ߩ�8��_��\�ʲ�w>��Woj��ޚi6����L2�+�S���<���OI��[yĺ�C}u����dIS�}�u1vY�Z�W+�� �&��ݚ��]Эޱ��#2�:�[�|�̱��Q����󥩥��k��%��4P�Ԫ�N�4�s�ES��z���a��uA�NR��M3���B|��::�&e<$�Bw$���\�1��PF�+�%��n'���[��g>�Y���n��#���~r�L-��Uڹ*��q�n�,V�87��[�#g^nf���Z��]�-y�Sڽ��?]�� K*���7A�դ�07���C�8�����e.}/L=#PK������\���RL�v�3I�q�D�ڵ��R,[�ND!����鷬kj���UG��Y���k�H�)z5-s������Y��lC�6�\:b��WN�î�N-����'\D�J��^�A��w�"�|�2�r��68-&�xw9�[��퍒�Lu�ί�z���R�f��I��])�Y�M����%��o�=�D��/(.��/h����� �[�6�e�\h:��n��p�eV�l�s񾹉�&�}:�P�^bo�:�Ɋ|�J�c��&͂x�Q��#�m{�r�x����ۍ��!E�^�sk/f��1���搻j�e���u�j��v��p��]�t������x^E�s��dҔ���U`pI�-��
�x&���a��E=ۍ�̎q�V�`�<X$ޢ�S����&�58b�1���Yx/~�&���՝�J2Nb��6��g����F�w�e�:q�o;�q�z��ˎS��,z�\����=�4[�*��+X�-s�yEE�/>�*-��=g!����Ǘ[X�Ig9n>A�kҟ�w �}:���9W�Ý����_J�}�jK?dq�Q����33��٦}��H��>'�Ɲq��,����P�ph��sq`��h���oA$^gk��ȦY��z����j�<�ΩGKz�eF�\�z��k=���k�A;��[܇͜�i�����3��P%�W�d�z[���h�K�f�tv�OL3-v>�����K�����os\] dMX�x���E�8��9{4��]k1٫�t��%�ft�cG绅���g.�3s�=h�]�������@d�͒a�ʯ��uEF���f�t������gU^6q�1�K�[�)\Cu����.����*���Q��/�����#Ǎ��V�-�r�z��s�Y'�;��t����-��v���X��5�V���80��I��l��{~[�K}7����\�a�������4ʡ���D����/gWH��LI?5= ���E���q�I�)�tW�p_Y�}�l���4i����o�7���΍#����v�fV:�Q�H}o��n��2ܸ�P�\�/�Ty��G����_�M�^�u#Ki�K���5@�$�6�Z��;�/��b���9Lv�p�/����}T���s���XS��N��w�oo�1�oH�x�2E]+��]��*q�.���R�5�sSY׏"�٩�Y���f���2�$Eqp�\7;Q)��+����4vw ��^@T�i,�Ntt��؋K{�И׫����-������lfM=�:`��©��]:���J��Y�\�ҝ���k�|_������J�b>7U��L��y`��SR������++�r���+η:�ץݫ0t��"�A�N�c���
]]�T~Ysj�ok"��&��U覊�9LG`��j;��S+v�K�#u8�wי��V���XAd�
"M{��k^r���jܾ���v��ۓ�dJ�.Y���E��i��7��ztu�q�%���� T�-��=�vӊn��.v�Csp�[���ֱ{]�8�vM%���V����HǍ�h��[1�.�orKz�^�m>�������^ӳ��q��N!�˯�����$��.�Uä�>���V�(B�����D�%��wrۓ�1��+�nDwϤ��.nx����.f�C�������]�d�]�{�:7�YK�B�����1�m|�叨%׷�-*�eح5٧�tݥ��O\&��7�s�=���T!(�����}F�0�>��w�A�e�<�5���]�6̼�5��6)Z�hw:H��wQC��=j��KVl��/'���/�\wh�w	��sp��ylqU5����I:�I!�/�/�暾�=����S�f�r��bp��.���C ��;Цt�-������ښY��J�kC͉2���|�Ǜ�����6(��}.���p��g6�*p�x�n��wk������/z�XY��E-��l�e�<���9�� 3��/B��]|�͜Y�����cQ�q�6%={Ʒ
(�0}�wh�.Lb��A�\u���N-��9��C�ı쁳�E�|썞����~cwc��A��s���T����)���r���O�',�B����܄�5��M��ΐ�1�Az=���ڜ�$�bg-A鴞K=��.�\E�Ը�����_���6�m�)�W�ѷg�|�ڳ�n�m�8'"uA��-�}M3�H�'�໬�����B+�4�&4�qy-˸�؀���	g��c�Z��ɦ����{WRSE%<ʄ����7��n�@1ʁ��G���ǟo>��t��*33{X|�y�k�&�_�O[i���nM2"T	|D����v�vA�vUHE��������}/��9�R}>�G��'�{ኹN(s�l�k.B�oVSd\:e,gL7:m�x��3��uR�	mvjM�"����Z�0��U�V5"����khE)@/�{��|/DL�S��������8 4�ú|_G{�/9\�s.�h鵩��'��ױ�zJ���+��F���ᤊ�V�t�w�|�Bw5�Z�f�;-����j�N�A��]�SK�y��loC�4=����y�j��T���s��tk��Ȁ�WR/O�%�9�Ki�2��k����ڵ�4_W�����uĆ���\��ՐJl���5�j��f������3�ҽ�=���eح�����k�g��9̡�g6��#|��J��C�9'�dA��|�Ts�5"o�������ڑ���o�S�Cg}�k�'}�F�_�����|�e��]:��n�M����m����V�{>�n�:�A�BN9���ɸ׵*�o��v�����Wa"�9��Q�P-m�:yA��e�T��7��7{�y(Tmq�n#mp(�g�]�KK(Dj�f}E�gފ�Q�����S�2eS-E��w}�;���{g��Ú���ꗖ����7����Wտ=�sKk��ݻ�Ӟju��(�A�[�ؕ;����6���f�< 82���twk&�J�rY�vI���\�X�	t: B=�
�ֱ�_��vm�#������t$디�:��l��z�M�!����eWcb�̍<m��m���o�����{W4Gd�\����<���X��g�e�������TM%�_��{-�}�C^L�ۗ|��/7{e��qN#��~X��q���ٺ%=?3-_�e���]�����⩉��3	L�(\�zB��C�ޚ�����C��*Oq.h�7�~�Y;�[A�lz�SK�/b�_<��nMC����-bC�����9��k���H|z�i���7ѷ/����\�i|�_��j?��w��ŏ�Z}�S=��V��h��m�_��3� ��ْ�a�xGm�S�j��>��Su{ӭ2���2�|�إjh��qoW�[�7�|ӽ���꧓��e�-�Lش��6�B���S�Oq���Ż�'��,p6�~F�K)d�ˮ�Y;���-���{of�U�p�;�@�O����m`�z0݊I�{v������YS�h�MFT���-f�[���\����H�NT͔�*��'�j����7]4�C#�*/�_kͧkw��
jN�8�]!��3����sbC`5}/�v���rG{3S8�E�JM<�<��/Zګ�wKv�޾��N�%O��N���]�&F�Ʉ_x����v��e�D���W�gp��X�s{Ж����Y�`�=����j��x0���*%������8BC��bb�y�V+I/FC��r�nv)�9�k�A|n#rv���dO1��4���:d[䫏b��J1G9���-�SL�R���::��e,��rv�]�-�&�Y��n(q\�Z�k#Cr�[��6�ϩ���w�7�r���2RK��aJe1ЋOG]�q����>��>���j��V��}8m������Nj_)���CZKVXn�W:Of�=���8���M꫾.5I7H��RW7#����~�O�}16��kr뼙証��X�ew<cY�oM��:�t�B���3&��ug���D��h����^RX�b��=�f^�eᷔ�f��X�MgKXփB���[B\�&��\�"/��6�I=v̢��2����OP��S�^�ɏ�M�c�ԍ[��uY�.dÌ��?)G̖����7,����]��F4+�o��H������L��fۏ"�9��lr���d�n�2����u���y`���]Su&����s�ݛ|WVѣ/n�;S��-�8ʱ|�Ƞϖ���teՆ�.!h��N^���G����{Z}���^#WӇR���
��g��7�r��/(+UtS����r�(V��1II��]tI<�ͧ'����Aֹ���ɬ�l�]������^�� ��)ԵOؾ�U_E�Ko�V$��Av;����j�yY.&S�Kz�G�b0�n�@��Y�]u��YYKv��)���?�+��u
���ccկX��Vj����3�cb��v�T-V��:�w_$�{��A^r��aȕ[7gB˻ɽ��R)̙�,,�H\٭��P(,���
��óm|��g��)��̹��)���YX��q��WPB��o|���bVqŇiN� xZa4�kV�kv�p�,�O���P��N:U���s`6�YV�mҮ��m�V$���<:��X������R�Oo�$ۦ���F���{��.���J�tǕ���ֽj��mts��6>��]�k�g$�x�mG�^�T	�X���`��B�X�R��\_T�d�իoQ�y��b������uرS���,�zD%p�a�J �*��r�[O���î�[VZ���NVsv���V� �����w�lC &�aCu�ȪY���]��|mG���.���e����d�v�[L�����vҥ��K�X�@����j���3�PZ��Ԕv���,mk�_N��ֆ�o�<v��4��WAc���k�����7V4𮔄���9��Q����ʋt��n&-���21�u�{�@�εi��5ӫ~����l��n*�VI����]��wJP��38CH]]��j-�zq�O��Ħ�E�wX\�n�'8gNN�t��c(�\Y-�9�����m]�Wז�� �Y���d@X�IN��YG��x5�:%]�k%�	L#)�00Tw��s��y�I�WA�ͽTv��J��y��.��krV3�{fxT�0���5��S��[ݸ6ݥ����i�+h����gH�����g;���U�M�=m-�}t�3)�Z,�i�U$�s��3��z�e�fR�@���#5�d��F�=�o*���S	�E���K��gP���	Uv�F��ҭi���T �{|D��1*�J�f����$b���u��Xr#Ң�ⱊ�N���n1�֜�7Mu��zR��x�qr֭�a�:�TL�8F�+ޕ�n�:��Q�N����7��@�)UP� "EE��_�5"fN<!R�����UymaÕUE+H�9�9TED!T�j��E�)�Ӫ�#�DP��
+�\�D�K�"e�tr9�ȜK��W
���\�DQJ,�鳗r�)�Pui2�s�x�T�Y*,�r�P.W$ܧ����ȒF,�(�AT\.Jӑx��W�r��)
��\��#�2T��F�$�\�s�.QG+����eU^Rg��\.�8s�#�aA\���R:�ʕe�mĕ܎'r*�H�K�9Ur�����*��+q�˔�t�����sX��Ĺ�B�UDW<�d�"E�($�eW�Rs�k�8Ú�Q�DD\⬦\�V�*;�"!D*.*�9��x��9���.7%�b �*4XUٝ8W
㔐ʨ֔Fc�$�L��l�2�I���]���)��7�Gd����[-��a�"V�%f7PumD�a��jb���M��yY�E���Hj_��\{�v=<�U���y�X'?�
my5�4��济ٶ�_��%�����怳ϷZ�xy�#r�ો�!���z�"�f^1�V1���T F��oa����l�U����F��NI�[��/����\��̈́��	����q�{Fc��y����j�SD^Uyڦ�\��E�{_��]�x��{ǌldӶ�r?hK[̸��3Lu���<�&�'\N��2ul^}�q<���Iy[�~�NOG"Oޯ��܋�x\��9շ�EyB1p�=c{�;���³�ȚS�n���/���淝ɸ����b��WGgY#\togi�g��k�JS�QGYy�T[���oz��^��00L����n>a�<�b��wN���p�Dꊃ��E��qH�#�I����ޙXr�n�i�Ek����=��yR:�f���	d�_pvwb��ty������AQ��-2R�t����^���Հ)����t'�9&�u=�τj��0[Q�[n�xΦ��bh��zX2Z�6������ĀjS������x]u���I�����G�֓g��+]Z�l	P�V E�2�LDʚAt^�gT�QNgju#��f㭅.V���|�oݩ9�ㅽY�ݶg>��{��ɨ*dD����	{������ŋ�0��<1���M=�jZ�}/��u���T��w�x+B�7�J��Fw����<��:L��L�Z�l7:n����q�2��
��#C�4 ���uＴ��g2 ����'4����l�6�I~�c���d��l8�V���T�h
��E���oN��P�2�K� A���un��otˍ[�
���'�ҹ���z����T�a��ڦ�*���%5Z���Ʋ�©�3� ��y+��yU���}�]+;)�L�e�J�����8��V/b�q�>B��	�܉�ۉxv�'#���M�s�N"�l��o-��׋!'}���������ї�*��=��0�/F#�ΰ�ږ����	�U����7�H(V�)&\�Szfeu���s�����=�I�^���Fn�"ΰ��c�b�y��
��E�6vm��6�S����fJ$���)=�_cun���\�����-�j>�BK̟%R-C7oox�������P��V�)����l���I�5��M�ܾ��o]T�\o\a��	�s�cw�������/Yd*nq�frUm,��Y���Say��vg�vz���ԭcޗC:�L�;�8I��o����E�t�'����	�::�ܚ�W�1��ޞ��	�O]`��+j���t�e��i���뇝G�m)�؀]D�[9���n���A&뉵���W�����e�ϛl�SL��R˗k6:��w�{_�
j�_�^�[������)�2��콶���_�c㢮`Xt4ʍKX�p�l-c�D�5	9[��>��Rz��ϧ:����9t�EYOM���'_�k����w����R���8��n!�L���W2x������Oa��e�|�M��:�I�7�R�@/��Ƚ�CL���͸��TL��OD^�m㋂ܼ�x={����y��;��u�r�� ����_s�v	n� �������;�>m8p�6�Ӭ�|6H5.�={ggrL�8��)��yX&`t�;6�]����L3wx���i�V#E��^� Bf��˖\�a����E�>�)�6��6�连1HOD�; �U��]�73(��x��,�ZE\>3֑b�f^|ƹjr)1OD�d˴]v��N�W�����zfѾ]Y��E˴̈́��bq�>Cb��w9fA��W���O%6&/�O1�@���o�>�]h�,����Nm��f6�tyy$Ϣ����|/+޷�f-��t�o�k��/���BT��4L\�80{P�"R������A��,Ѿ�}�Y~߯�ma�:�5<s5k���	U��]���&�������Smt)= �)}�eD�WY[W�1Q0��� �9����v R_��-e�����=e��N�F<;�N������c.�k0�޸�N��a��Χ-�SL�E#����S�ho�y�+J�n�S�z��hԆD���ϧ���ͽ��!��S,�Cm$��η;���U�N�Wo*��U��n�t���bx��h�r`S2�2t�S�CR�F��ͽ�g��X��m����+A��j�>ޅ�Ҥ�H��\�A|�J|��OGu�@/,��e3��S�&۠����b���]�����Q�%�/�Z��|��U�n:�6l��KzŁ���r{�^Nhn=���}�b)�"=Dz+��Ö��4F�Q-G�3���O]g�u��}=#o�I\Dܚ��4�Rsq�$��S�N
-,P��q=x�Yu:d��79���+�%TA���緢U�QK��TֺƎr�5-�8�.$⦖1�ӝ����9�6��'�1�,��ue���W��q��t��6��A�|g�"�|�2��)�E�Q�nz9��Ɩ�����!9��Tή2���S��R�3b�$��6�����K;9r7�	��p�	���$.�yAv��{N�E����fuTF΢�w��p�6苆�s�Cn㞉������;Ov��\�:w2��̊��'Vnz�}����Z�1q��n����Rjq��Bs@�*­��(�bݢk��^�Lm#3���S�-�����Z$���3�S�3yj��YXx���0%��L<�E�9�H͚S}q*�7�����lt��ޥI����%i:�J�1[]�T�_+kUK5�#��BK�b���s&֡(&��Ø�37�k��a.���ˤ{Qq��S���gYyS�I�5�s�7���C,��Q��z��Ӳ3o0�דh��q,�����s�yE}���
�s�S�q��Ϲ�]%�&�@6��5�H[���p;!�VV�P�b�Q`"܆Wat.L������A�E��N�r^Ї*Y�aJ��ǵfKZ��TiX���Z��	#3;_�e���83�`�S=���P�w�t=��39�q[�/r��!g5�g\h'q�������3��7$��߂��Z0�
2��N~�{<�ǘ{�·n�����>}/�!�]�J*I�������^N�y�8��8�{��Z/>]z��l��3�k\���=cXJI�^�g�F���3Ͼ{B'��M������̜�M'9�[�#Cqr�l;1��n�0�l����}�5{`O,ձ�K��v�����~6n��}��&�w��Q�2�4�&�4G��z��|��{�$��z3��i؉�Z�¹�ڈ�;:�`Oi��k6�wj�������w^��K�we:�n�[u.呜:&����júm5N���w=U�[OQd�c��
�5��T���䶻g2s���跌R���V��=��%9�
�z޾�������[l��s�6)Z���	��'(v���YWw��R��>L�j{�^s2G�X��crQ��\�NG)��p��=J��xoq��t/�����E����>�\"�w�=���o���{c��
Ѝ�Χq#�vRI+6Hv�_���d]>*�8��mϲ#Nfϧ[�����g�r_h^�G��5�U��p�"+�&}6�Fx0;�T?\Mwy�����v��fn3���z�«���U8�j�I5�do����i��|���P��ˢ�������-xK�������������;�fa�}N��
�F>�۳+W�)�U�ex=�T�\@�p����� hvr������-i'����/"{��2<�xx�F{!�=������&o�OF: ��O�qR�>�����x�l���d��G���G�>gג���#�C���{���_�G������{�K�4+ٴG|>O��=yiR�
��F#����tq5n����b��ZF��.�����s���J��kF;z�˭m�ѳ7��w��}��������u'�Llõ��«�[��H�c�2攦��sb]+�B/1����������,6�Y��1��9P�YZu����L��z���G�G���!<��c!㼛�k��3�G�������9�<��������̘��c`���{��i
>��>�#���$9��_T�}^���nq��t�y��v�*�r����k��w��>�jk�G��<��_�LO��*L�D��/�j9ϖE��dyS�H���{��YZ/}��]i�Q�{�u'�Ni�$&e���QMّ�&��%���=~yhq��K��c�rSpq����G���H��}2cվn��|.�	���WY�]��G�.��OicG;�o�v_0d��?�<T���z��<��~���b�f�cn`���q�JD�4���!ޅމ���u&.s��h��J��5���B3�߰P~��(b�ƣa_.�F�ڵz	$xp�<B�;P�}4�@�����~"�8ۓ�5���a?fT�k�Ϫ����=Hj�y���(���qޜ����E�k�+�چrk�Bϯ��2!e2<�����9���/51����ك�̥��L�������� ����U�B�W��@���n�����i{Iӵo��ާOJ��[^�q�Y;4u[�h��LZ2��2�j<D�n:쾛�1�MT��W}z�!X�i�vH4�=,��j�pգ6�t���B,hr�WNP:�ۙXWoNV[���ި�I6/wj}�K��kf��K�k7>h����݆��+oaq������ď�c�;^�� �F�Jˀs�i�Y[CHr4oU=�����i����*�6K�Ƿ�G�^ xh��M�.k#��ׇ���*=�V��/�ڮ�^�ÞXQ֪��|=���Dn����9Yt�t�׮R����V}<��<�xzC�����G~��KG��/em��U�w�Χi1�Ղ� o�
��Ċ!�E�y�.凱'ג�8z�"r#�>�Oo�~�Ge�D�	�|�+�wq�������·�\x�׆F 6*���nr.�!�s.)bŹ0�'��t��K���[$�={�������G޷>�Q���P"Q�)b�����#�V��+�*�7Yi��\�)-����u�<6!����>#"=��{!ݹy0*��*�a��V��H�u�JK7�ܻ��y<ǯ���G�ؐ�u]���z����T�G�ث�U!��PFJ�<�]��yr�z؟}Y�2���TCP�eZ���؇��c�Tx���G#�~4���=���=��ʹnW#���7Q�ȕbD�ʮv;^����lOz!���;�,����?�tџe_OmYz7&�+��|ir̷��l�՛t�a2U���F�Sj�ņ������պm�F��g�������s�.1��z�魋�Z&D��n�V���:�je�J<�Llv98sYׇ&1q�#�����έ��M�9��G�N�.�ܦ�RE���=�+���@��t��L߬m���s�}��O��eN�d���En�Q���.�|��)������캑���T�0{n.����K����d='O��1�f����Y����I�P��z�}Y�W��}|d��o�0���|
Y�~Ҍ�u^�_p��J���G���]�c��G�^##NnCo�|?\Ϩdo��vD7ۓ�C��NBi�%�>���foC�v-�Ӟ����u�k���Y�u~��+�z�����G�ج?{D�f���w���߼���⟪����z��t�����������S���_x/z�w�ғ��75�Zne{y,+�L��؏�ͺ��,�������_	�S>G��s6����k����aZ�Օ�;����4��Dw�ٞ#��R��]tEπH����nz���e�5S
le�����a�f�=����������b��}(eYQ{Q�i-�qCu�!dp,�6���+V���N@���d{~#���C�ݱ9�;����+$`	 O�ﾦ��<v�{���PP�O�L�����N�m��@.�'�6����0��ᷣ�JLrXZ��zBR�p<��d{pO�1
�chͩא�\�VU��9�|�KgU83Ax��7Òn��ݭ�؆-�/�r}}��[��J�ӳ��:��¥��Q�=��3y�=
��vw�k����W�:�T�s��Z5�ȝUF+U��*ۤ���̀ǩ#2�Z�]��J*񎹱k��T��N9���*u���|.���*^ʑt�"�@��q�:�cљ�E3�P�4u�جBv�ņn8��eH�9wHh�����W�4P9Onm^J2Nᯅ_���O$��)'yZ���*���^oH1-���]����Vz8�O�D�:^�l<�-d��M��I��Yn���lJ����1kwL��j=���[X#<�7;�$՜�d�Uat��<�0�4o$��iݰT�ApGL�nQyv�s�RԎ�H�/A!�S`]�4��|K�_'��z�iѺL�-ɒ�9���,��"^qR��-�ffӎ����W2�3ɵ!����XÕׁCO���X�@�Xn�=��kL�@XL͵/��e��#*p82�������
0&�0.E<�t��x�WϑfHX���R�&�Ҹ̟X��ob�3C�:�ua��a�u�0*=�u�]43��S�Ό�z�
=]��Z�d�����K�k�+b�̱[r�
'�v��V�t��(��0��sK;c2[6V�T�T�~��Q��B�"��5݌�n�IηQ�6�zm�W�.&�.�	#�Q'��,X�{�Vm4�c3�j���Em<�v��Y�=���KJ��[r�aH�c�ϭov@δ��0�,�U+x��Ge��ue`�z��va	�1�*����
R�
ld������k4�*���u^O�`���sP�+����t���=�m�`���V�cU2AM����M��֠��W�Җ�|��l���e���
��5m`�f��$q��Y���Z`wb/�6r���u����5�tN�[W��K;��&���˒�U�ƙ/ ()6����Wv,Ȧ6p˕+B<qt���L�Ւ���=��
we]�m������}i��[�q���囈���l�f�}#ۀf�šrb���٫�m��+^7v[��VT��P���+�X�;�4��[�.�������E��$J�fM��I ��q�]�v�>�)�@6�vˢ��(oQ�aL[���g]��c����mu��e��,2>�n�h4�^u1S��oQF�."�bim�
�Qg̍o`"�VmkZ��V��݈ �D��
�/�1�5� 8�I46�N�,a,�}CW� ��$u��P^��i1tu�	xr�t�8�|-�:&�c��*$%M�@�T�7y�vVL���*�fq-��aʂ�M��yV����f�X��^̼��F�n���)$�D��V蓺��R�̎�&��s�����]�*
�����B���p�<�H�3��r�ˆ�L��9Yq�^%$�t��k1iETx��T^R�i�0�U�E\#���
A4¢3�]D��s��/)�F$T]���T��Nr]%�W)R��J�RB��kK�RW���p�8N1��s�(���[�G)�����<��#+�&Q0՗%d�4�9�#����P�'�)p���RT)���P�ڋ���&�d�EʖI�8p�<dJ��n:˓3Ó�E��,�M�h��O8��V!9O9Ê9TQEP!��s��9%�DN\��%NsW9�ʢ9Y�"*��/#�r��p%⤻����8)P��rVY�]s�!E�%@y��
+�rBQ45T���iAWr�E0�Y'*
��Ex"�4H�C�TY)�
����8S2�*�UN��ƀA"P�y�ZB�v�׺�e�݋9켋� �BKN>fY(�=�2�yO��(m^�4mH���sOS��ӝ�]Z�\��c��'���tΟ�ܺc>���oy�<��|=�1ޏr�gEk"FHC�v�rk%m��Eo�����L��+>�^�s��_xo��Z��_�ON�g���*{��]y?l����Bӷy�+��{���NPB�d��Tϥ�BvR��(�Ȇ}�T�����㞓�#ܢj*�Z�ݯ�w}�J�:u�b����M"�z͌�SCǘ�/+�p�yI�V�w/�Su��.S��k�C�����������o�)���*[	׬l,����M�.7�ᐶ�Jb�e��5�垡���H���~���5�<��
A�g�S��
�d׏��`J�{;��+d������ǐ�}����(dF�~�{޹��.���mP�5�g����0s��5w�5���D��}�O�N}��9����1�܆���B�~����z$���V{�3��`(���g�Ǎx!Hy���چ�'���׸t����s�9�>����cy�����Fy�\�䋯cc�$�=R;�s�'#ٷZ3��>	��]�^߈�n�Gl#�fn3����NX��.Yx����K���}J�(i0��|�bTkt7�a� \s�pӚ�
7f	��7���%X� ����'��/wК�l٦��u���m��؜����u�m]�ǯ5_+em<�l�>�I9]t��2nt��pRnw"7�V�{*��6��9�0\j�傱u6�=���y̫D�k8��y;,=�������칇�����c���=73�11�����z��0��G��o���l�����^��Cb�ƳM��+��s�u����U=(�-Y깿Z���]�>�-���&��z,щ���^�qޯ ~�������7�4�U~F_0p+_`�՜����[3پ䖓x��O�j���ꓨȳ������_�g�����W�ߞG��+H���UuO�ݑ���|oڅp�Fz��X�3R���k�V����5����)������O��e�k�S��{=m�k��n��-�=A�>G�)#��ā�:�%[�q^��{L��;~ΕX��|_����Ww�!r����u���p��cP��)�rv@�T�t|��B����u��[>5O����Fz/�m��O�א��Z�D{�u'=v��V�̷W�=�,6�G����g�������o�c����c>�Spr�66=U�{�ëd{޾�c�D:�A�Q�ؖ̍�
}y�ᯟr��S���]&:yH����M���z�{���Ǫ��{X���u�	�_{ۯݝ��ݿn�w���Q g�\ʉ��q�����dE�����:wc-�2i��@��2��	)7NU��J�Qn���D���k��m�y&�Z���=�%[r1:t�k�U�j����w;b&[��vn�VkK&Up �n��,�����yL��	���;��3��������(\���?%l�k�'��2�6�b��~�D�r��x_��=�]���K��x��@_� �N�#�OD_��gN�;���ܜ��6\�'�ʞFn��d�{�X�]�����F�)�r=���>ک� �D3�MwY����]g�Ϯ+ؽ�ꢳWI��)��W�����}��φ{���?�-6jܾ+<ڱ�?T�y��/˧�p�h�=�3��w�Z��&}L=��{�>ӏ=;�;�p�k4����^\�Ý��<��#���4��;Ӈهo�=N�}��N&�w�G����V��}�V�aC#�mWO�b�19�B{���5��cB�WN��P����\�V�:���瞑�y����?L�o3���Ż�����MFE>�������K W�nE��eܰ�$��^���D�����{tdMu{=�0x�zǫM��N���іTBQ��w���<�	d�d5�u=��B���I�W��XOe_�����lx؟�{����2�r'�1��|���$w
jc��4�YM�+m���1�����������;����*yW��Y��}u�oh�X�u����Cs�⍯7~2��6������+�^�q�M�(cǏ������l��&l@n����Z�3��P�zV�P��6f�2��ԙn�km(:Fj����g�Z~��=�|�y��>���{ۗ�# W�*��*���{cwy�m,�b��u����I��7��k�,�ȏ_� ����A�G��S��)�!�+�xש��ޥ�ֈsb�^�5�jF|E/<�r
V�k�cb7��<�G�����(��uލw�C"��d��q{YC�H��5]�#!R=�W8���=W���Im_�ˏW�
�vt^_���{w�3y�@/q�7�w!N�ɪ�쉣�.)����7)�W�[�dy<�$�����>�**���!#h��^�>؆2:f��*E¦�,�ۋ���ὔ��c�n�Z�S��k�J��Jb�c�Wb����~��R���$y���A�]H�^\��F@��J6\.~u䅒z&��Ny���ǐ(>ח	���7�~��Pȍ�\��rL��������� uq��o�x�����9��9�^ߧ�e�i�g�qd{i���o�ߢσ�>̀����[�����w��'㲊�w��b��xxuvEW�G�u���U�5u9���HT^9�X4ʟ��[�	�.��}Wvk4[ק��fPg��!�(&3[\�&��JmnMʵk쾣Δ���Hՙ2�n��Hf.�EP�r,�"u�.f��dp�x�s9Vå�f<��X2�;���6��n�u�i[�nX̶���&�qu���Wj&6����&
�ͺ���r��*�0�G��^!����s�M��D����z���k¦��`�G{N�oi/G/1���~Ao��S�lC�<���� JD�P��v�Yw2�n��Y��^��������;�N��s��|��g�Ϟ��8~��45�aߑ���\�с��_����O������(�����f}^����r=�[�~���ed�Z� ��F�FgxWn_{�ˍ#l��}�"ꑯN��.�v���y�6<�x27�=�!��Z��>/:���*�����c�g��Q���Rb�M6�9}�~���W�N�l��C�ξ��v��3����Q��W�����D�L�\*e�f����]�Q��ϱJ�W���]��� �wrӅ��fW��@�w�(�����b�
f%���TR��r�=�͈����L����ʅ�7>��c��z��
���z��{}�N����C�6b!/G����1��$��qӅ��:��Cc��GMg�{ޥ#���̟9���[�V��f�O�S��Vl>�Z+�p��I/)G�^ǝ�iI R����AЬ8�q����1����N���cj���Z��\�wok���]�(%D��g�ӫ�]S��ҦY��LkY͸H�Y���s�7JyIζ
P��[m���a����Oi��,
7�i�0��ض�d'JoۖX66��{�=���(g���
��d�~b�n��r:Y��ϱVwTxӌ^��%�ˠ�l�ݞ9��8�!�ˆ���G���P��z$����'ʶ�U�ڑ⇡�´dxxq;P�}=}/.�ç; �6���3gӭߎ�*.R��;��g��QM��~��Ͱ�/�Y��ۜ
"*�k�CȽ�����q�Ϸ�PVRA�
�ŷ�ϕ�t����+�޳�ת�xw����ͺ�ϡS�C�c�����=�:���c����N��0:32���Qn���5��mٕ���r��r2��Ȫz<��.�}��圍���ŷ~��TG��N'�I�q����xx߮����}��7���H9���T��J���_P���p�躦�2"˹��\��W�=����l}��J}4ۥpr��A�+��h���0Аd)���sAR�+v�x�&��zL�����GIJ��^������;=����=q��!���%� ��w�g�Ȅ�/]Ey}�i����I���p�`t,�4��[��9
9RR�frm#f=/���Gy.{�S8(j{��%��Kf��ժ����Tk��"7�E��������'�CՍ���W\�P]j�ݓfN����-��0Mԑ��j֘�N���k7��3�c���O9\�hd�_m�Rr�wR�H��xϚ6�]V8,�u���C3�����+�T8�n����gW��Ug����B���z/%�_���j�6��/��R@ϣ��9�sL �~�&e��3OU�Y��ޚ��U�V�_��9�Ms���CSpq�cc}U�{ã�o�dD{��3���
��T@�D��Xx��֎h�@�	�����,� d��2<T�mg�{����b�dg��r�o����KH;~�zPu�P�I���Q��t�YJ�z��C�̡��
L���F	�Ϊ/|��fqF����E�G��@j!��k�"���߻���Ny5���[Z9����Ǹm�Nuj��T�W*�=���9�ӓ��u"�5���C9]�z�B��x�����;�9,��id��gs^���.��/�^�����d��v�0���U�����z�A����k_��m#��<�� 8x��j�>��w�a��j������g!em�NG��D[ޜ����j8vmq�V=��)Ys8<�#L�gY��zߎ��}��yj�.>�}��"�3��Sw����p�'��	��uq.J{�pmL�E�:T�E�ȷ�ѽ�N�����n�S�"&��M�a�W&f��"Q�͏J֒hu��9P�]�3f�����O��̳WZ��4T@���u���+��3 �֐15�l��8����a�C�;"���^�t�t�];�*���VD��Hȏ;^���~����O���x�n_y*�5bɍ)��J��s���!�]W���XjO�%�p��D�E}�@��=�>X��2o�w�_�U�S�V��5����*���+�����mR��_�z�_�2���#�H�\�_��G{/�67��b|}�s�IQ9A�H��+��κ�o {��S��積��Ȧ2#��y��t<��G����U:]ۗ�# W�*��*�~�(�����_��8��f}9�22}Mk7��l_�ǳ��Hk��G{�8/w��Oޫb�7�^q2�W�_3s�����甂<`O�BG�FA�)�9�(��2�J�~��lz����Fg���[�lN�`����߲�ď�[��(x�.%_��k!R3�Q�9�q��|pOg�,r��el�/��7*�%����vxh�Ur�x\tM��qWS�r&��h苦o�6�]Va+s�9��Xͳ��Ī��3�VeNG���{|+�'�eh��-��ͪCtc�T�鎇��a���OKw�'��`߱�9��B��g4A�뢲Cyn�`��ucܶ6s�[�tTg�c�8�x�ɐ��ۈv]β���_fpqA��(>�7��e�I+��H�/���؅F�8@M%��g	�������'��_��dy{oҡ��P�~��VG���#�u�mT�U�č�E�O����g�����T={�o�w�_�p��G�⩑�sr���6#��g�3}���ܜ���Z+F�Z��U�����#�#G�:3���Y����lq��qd{i���l7�������Ya
>�K,���(|�~������+FG��W �����.��Lү�o#nf�=;�{}#���������u��Y~h�����Pjʹ�)��fS1�/#���p�'���O[�u�|�xyyGG�����8�fyp��թ���N����9�.�#>�,D�P�/�h/�T���o��6Sk	8%zfק�s"w�����z�����P�3����FS qAx/��b�_�f��q�j��,Sc>�R��]�5��p؏��yVߝ�V�ٕ`-LA��|=u>�f����{�L�*��U�W�an]1���4��o�T<4<}�������&w|�ü��^�;�#$h�@�>��jU/
�4�s����{Ԧ��ا�a��hU�5���������̢��$5���TiSue��b���6��������m{8F���bc �錍\�c��0�a�ͻF����ޤp"�[����,aJ>F�����5���2�o]=�JRa�Ň��f�M����kt���UYJ(��Uu$�gֻ�m� }��Wz��fr�
&e.2#��BHε|�L�ԙy����gKEXE���(i�=���3�w�(��_�*ؠ���ķq4@��F����GukF��R#�~,�����~ԴI�����z�q��2=�Y��z��z�d���B{%Fej3����k<�o����u��!�dy9�)����H�ǅ�fO���yn�Z��~��~�]� �?e��=�C��<=[7\���rׁ��S#>kݑ����P�����\��������mwi��jo�s�T��?Cz�m)9.�]�g���s�{�dcY�?]����~��V�EX{���FyD��{c��Z2�
�jȞ���u�9��dƜ�Ɯ͟NvI�x"F�,WkY���L����$�K��גG}X���sW��|��ݭ7?iLON��ֹ}ɮ��~n־/�u����9���~�����=�������ͺ�ϕ0;��P�O�CȠ���]�7�e��oG�]x�ힿL��I�T[��n�Y��t��qNG*�ǀS��&�]	�p���gk6k�So���e*%ǰj㇥"	]�%���m6s��.�1�VH8R`��Ĝ`0��,��SI[ �c~� V�t�"nكtBz�;��e$����y���v�����i�r��� ɨ�����k�uF�u'��*=g�t��}�%���S�;�C'YPn� �°#Jl���dɒV��-�}0h�'s#�Զ�V#��B;@�V1�l���t\
���H�]P�[�3�c5T�U%�O�3Օ��\(�.����H-�k>���(2��y��ލ]��ˮ�y�)�o�M�I݌��Ô�6��]+���mp���&vLt��5Qw	��si�ʍ$Z��eqM����d�#έ�)Q���3sf�VS�s�Y��sTڻt��2B����J͛v��r�Ve��u7c�2�B�4�{h�z`�c�Nf�0e�-�P�47J]ٽ�Xp�J���U��w-�١�M��������F��mt�\>Tr�i�������9�Ws��ǃdN�Ƕ��Ű��J6�M/2
��7�����v����Z�t�\�5Q�6{'u#�56��׺4���s{�yGm���T�1'2VK�3���V���ՋxZ���*����~V �jn��B�=����*���5 �ڦ��7,Q%������n���:�"	{��V
BS7ێ��N��U�����8�Bj�t7�O��.�t�W�XT�U��]�h�ºq��>M�M\��*�&�r�Sv�j��*�tM�X��8SGn+
j$.o-כ)BZ��C(��Z�7�E�M���o����O�w��8����z����\���u�Mкx�΃�|��#jI�W--��w;]��|®2I���<��T0-B��g]��vEp��(\�Z)h[(Ǩ�(��)J3RaX��e�B[#L�j^���e���a�	Er䓐��[��*�c�w�(�,)=Z�U����`���v��0��3F���5�"�sj�-�9ָ�jP8�K��	��2��Ԯ�S��Q�cU;4��L눝�졇6�wZ��d�j�Pop��'oX�N�b���tU�;Y�䡆�e���K��r���!u�SI�NvD>Pf�(�a�{�*��}�f���	58<(+Wu�:QH�+ڵ/y��Q���֠��^�����N�.Ua���P۩�fj�Bn%�eL�:�Hh��m�F9V����FY����,��b��F�\�j3�����X��|�ys�T����׀�ۡ&Kk�sot�e"U�|���x� �ًn���T���5+���T=({(����c�w��Mf�맑Y�1ƒ�ef��1ͽ�m�ϥX�&r�'wus��Q7\Q)��K/���S�㙶[Ta����d�C�B�qU�K ,��(-/���ܶ�e���� ��
 �C�>�$�]"���D�+C[(�#�Ȥ�}�pv㫜Ex2I�E�XU vd�\���!��:�*�K.f��ffTYˮr�J%,:$.p�M%$�UʔKR�t9�xȼa*&t�)r�9�q��x�ȵ�#��\�rT[��+%d�R�"���58�+#L2%XQ��L�	R�Z�ʨ��,�!x�$�D�l�UTUUZU��(*\�9B�°JLS�h���G�8�P��)1&���jŝTëY
�I�����M�j*eVR��U-.�NQ�#�&�W�$Zk���q�]T�ZwE����Px.U&Ns�����i�Y"��g+6b�C�rV�V��U�R�<��nI�d�+��k��ay��)-1�)�˕�Tdd�R<�-
K0�X�s�(��'C��s�$�)�p�U�Jq���.��w�s�gZ^��1�P����Ml0�L��tcE>�_�9�G� Y�u��oCѮmR,j�:1V^�=�\�c[�D?�=��l���=�Pz%��޿�t�<z#=����dq�ڞ�֖bq��3�2}���Pɶ �UzU�Q�@yTu�r3�h�_�g�Ǉ�o�^�@��^{;��>���g�%5��}+x_��^���q��D� �.����t�C�y7�׳�d���1eϥ��+4ުɿ�G+���G���y���#�����$9����G�[<��fg3s
����f��d�N�?��&
��Jxºz[����Y����A� [�r2���kܤ�J��lj����ȼ�=~Z�a�_�=��jH�]I��ۚ�uAҙ�n�j륗r0�oWz�7�"�t�}.��b��T�o���G�ޣ}#"=�a�Ͻ[�Oʆ��T_!�g�\�x�xz�xdBk�N��,����S��7Y�������崫�$�5���$�)�}
�>�wª=�5��N���}��{	[#���?,���9��F1�E�O��@�o5���C�ԢK���5��s��״E�Mvt�c�{m��g��y{�u��H��U����w�����g�4�Ɋ��Fi�q�n����4NVDl�&�0ئ�-����VG{i�@�P}Y�L#@̼qd=�G��K�����H�3���	�c9�lssj	��X���s��J{\kR63�u�ul�*���M�7g���5ց�-t��Y���#��s�J���o�s꬏z�2/oN�~ցE��cz_�n����>�J��^ZGx�Ҷ%�۷=9ז���߈��
[��=�^J������#ex:#ˏ���9�n#_b��FS�����F�ᑧzw�w~�5��j����������Q��n�9{ogsɺ�\<�p_D+'~���<���3����Q�k��t_����8�ٟ^X�����j#�q{AD_�ǡ�ڧ9�C�dUzv 2���:s�s�[�̬�瞑��k��;�sk�z�����;_c��}d�q�{�������6E�".��dYw,8>��V3ϩ/,��7Z��H�&���'�7*������m���l
�!�C�0��~�J��]RC�_�k���9��T����W��ܘ����Ν���o�����ϸ^h��M �dp
Hng���Y��m��b�oB�Ei�5{�oC����s"�v�źw��:tv>�>#=��y�9qz��x9W�A���'��*�'L�z�n��C�5;֤d����f�y��Y�z���.
=���S�9yl۞Q��E�]��U�A�3��?i����C(���Z���u���0�N��%�v^jSZ���YW,z���}�G�K��+�������S���dM.��@��s%>��4�*-E���z?GO�l�R���^�-Q�&��E�X��c٪c��gl8��
�TH/���FSvddO��tCPϡ�jV��6#~�q�0:�39��[Kyծ��>gw܀Ԯ+��
� cU�7�lM}AyUʷKÔ1^�g��$��U�~�q�f�"�OO����Wx�ؗn��!N�Ϧ��飢/�f�cl5�l�WeN}��(9~mL_�o8ؓ>~Y�9��؏
����2��R7�Lq"��>ʃ���8��kSJ���=�lzS�7�q��׻=:��(dk�����{=2G��\�uԋ�^�g3ygyVe�����i�t��Vϲ-�p��d4;⩑��7!�~�#c��g�7�P5�ˑ�hA領%��k��t�T�2�����������Yl�F�ᑧG��W��ߢσدk�}詘��yk㤎XҬ�����3��
ѐ��W���=].���U�=Ne�w�ǧ���+Ժ�x�y�RjA������T�~�i���YW1�~��Y�>G=y��p�'�gɍ����S����n�������;�$*w���zF߭�-�v����jr9u�>"*�nw�^ܸ�.�.�Vg ٛBdN����N�k{5`Y?uq�L<��4I[�*��x�=rʕ56��H6�cQ=��U*V���D��ל�ޫ�PqiΙ�Ud�콱�S���Q��q<��y���IO��*��=c;&�``�h»���irU����Y73�o�n�kv$�������ؿb�J��3h���� #��?C5]���Y�Ox�+�#�+�H(q��M1���{��p����r=�[�~���eyfW���c�V譮*5���ߐ�5� z�*��%Q��ӿ-˦2!㼛i߸(���؏�z�=k�VjkׯNQ���A>�Z��FH�	�+�Nf^�I�Ýg/�6��SY�j�K8�����~�_�	�T�k�������pY��Ev}�!�NPb�	��L��lМ�5Kλ�b��`�O��c}O�3�ƋK�{�g��Vzv=\s�{޴@�z�z�QM�Z��65b��a���e��{��Ҷ+��/|��y���&[�.=^��º|{޳3���E_Ϋ�K$T���u�6|rWn���w-�		Ѱ�:ɸl{�����z�{޵#ޚ����1}2�
��9uk�u�-嶗���~�6|*��[7M��}�~`�؄��׶����P����:��,p����x�F����K��>�;T/�T j�ғd���p��f�6��l���܇���YH��8"U���ZB,Һ���qTYS���z�4Q{b���{��y��|��c���i�]g�����rQf�0A��*��� �H����#V�խ�k��Ty�q< ���w��}�����y��ՠGN�x�q�ʼ���g\�9��V�{竓ДP�����9��ՔSi�e{O�5���q�E׸t��d�mϳLw<�u�;�� ��o�L��흍�z���A�䅝���Ǜu�80;�T/\�p�������̓{�ʁž<��������w�zv"��;º=�>W�'�>�R�;6�u�}��p��7��^�8�a۷�]�����=nfn!sX')Qn��n�Y��t����9ʺ����}��wC1<���ez��X�\{"�v��1<=�Oz��^��~o�#��誁Uv|u��}Q��O�z���1P �EW����yU�Q�]�u�3��zG��=�<=���S�/�G}�iu��z�>����߅i	��FW�9�s�3�#��aJ��+��)������\�s��o�-'���e)T�}6<}�<����.�Hs9o��T�̓��7�0���5#�=��ž���_��;�o�.�+G���v�NPb�	��'���	G��:��zl�yj]��y��T�}��pPg���z��N����zԐ2#��9�5pꃬ�R.�F�����E�N宊�.ߪ����b�J�5j���l�@)V�P�50�.�eN�b%��	�.��y­�����ܣ��rM����C�i_RF��\�뎙$�篦S����ज़�+��D���
z�2l �9*�߯N���
)�l����ׇ�MEi�"h=sQ�.3Q��66=U�{ã�o�{޾�����NSݽ��Z}�km�����@�HdBj)���,����S���Sps��z�D{���(��Q��r�nw���rx���cm\
�^�7�t��\��E�V�Ϛ���o��Vqn�yn%O�A<lP�{���b��״P
X�v����gN�v;�.f�����F�7[�Ïx��ߒ��3��̩���U{��#������]H�^\�C9]��g�^��î��vv��4s����I�.��ɜ�9���n��ls�υ>�����śu;�u0;۰��ߦ�/�tN9���(����f�xy�z������pD?iǞ��w�[��Kˀy�ðF��G[�~�w�^t#E���>���0��"���ye�u7��<�Wx$wE[��w5��A<|�����a�ϸf�t�/P��9� �7^�ӟ];�*���VO<�*	�/*��X���^�$_�A��_�[~Y_���ˮ��,�n$Qr.��Qu,0}���[�`Nkۙ���� �+�H-���Ťmb`^��9��h����@?]�}��.R��5�����鸲m��M[?_�{Y{ճ�p��k�n�v٘�Љ^��(�[@���䧅,�c{F��Kn8;R��\��os.��@9���sr�% ����ۿ9�GjD�C���{ޯx~�>Z+H�Gn�ϰ0���R�)���X^{�;�F��ں��u�E{=�0�����;x�{ühO�}�c��[FVNPAK -�ۅ����g:�^�hߠ�����D=[��<g"�;��0<��6'�{�T�wnX�{Aó�N�Ǜ�[�<��}�3>5q@���ߤd�l=�o'�ߞyd^G�ؐ�U��x.�W��ػp�[�����r>��#�sO����v&���#�����2�Jߝ�q�QgK���k�g
ѷ�G�5G���d�
��T�u��lH��W;��1^�lOA MK��Lk���r�lM���S�W���Wx��q�7�\!N�Ț�^Ϧ����o��[|�Z.r�sH�̫KN`z�U��/#���N?,ʜ��~���zd�~c#�m�r�Z���T�/�шD�s��ޗ��[]��S���e��׶�)��P���{��x5;W>��u�^òu��>�<k���W�@��Yn��DvW��S##NnC�oلo?\ϨdF�.L�>&�kO�-�~�:ӗ݃젒gb�����g���ٝ���ۇ��n=�e��,�4��m;��F<����=ש�.��3�.��yܿ%�}�z�+8�S�[Ц�d�Sh�bXkse��w+O�)˕���6t#ڽCvܥ9��Q]�}�J��XÐG�^��OWK����D,�@#�~4����:�p�7�ޱq/3&��ͣ���W,��4���t�>*�8�����Z=5�迋��'w�m���}a�"x�2Qܳ�yg��5�G���}���aB:�B��T=���׵|�k4�½��Xx�>Z���6��S6�ؼ*i�_�8�[�[n����9ˮ�ϰx�C�m���(�ٟWn�����ۿF�/�he��Ϟ�&�ad�x'!���ў�>u�S�*���;u=�^�+/z�̉��F{[c,��P��o��P��40�8�a�w�����������o��~�y�����]�L��h�7�=��ޣ uJf���}T�zun]0����4��y��j����=�xk������Sw�a���'��&gˠS���R𬈓M�:�_xm�֦��ʖU�S+�ڕsGn��eV��yA����hϢ8n�=A��0�|wl@^u�{gO����8\y\\�Y�S��<s��9�=��h��{��Dg��1A��&%�؏�������7r�p�^���:e�3��N��'\��<2�;���Y�ǂ����a�GY�w����K}{7mB%w�ؠ�u{U^==ԏ'�
�ی�P��P�*]X|��Ŋ��;|�L�iGOL�Y't[�1��"�uv��=�0���h�~v?Ges����OIo��z�q�]>>�{�f}����U��-uy=��z+A'���t|�����Q�z��n±���r�C󛃉�����jG���̟o�_L�f���y�[��ݯ�A��e
���SBP�5�yt�:��*dg�{�=�]�dF�~��{��j��:�]k{0�Nw�I~sq��"��\%����N��������Ƴr+Ƞ��e�޵�tOF�c�mź��D��{��0�p��\�CQ���׸t�t@�\�|zy��G�^�'3��^��B�͕:�~;��'�Ϫ��Μ�y�Z3����[�SIXg�����A3d�G��ӣ#}��zfo9���;�w�w�g��/^O����f�N�ʘ�dUpm�4իE*;�s�Z=<�E���t|��s3B�NE*-��w�o�۳+W�)�G���;ۃ�[۵�/�Z�%�Q�\�(r����J�t�LvŻ��٘ܚ�	��ʵ>ݼ�>*2/�חa��[C�� �R�j�����Ϭ���!�^K�=~�N��k�s;{��ǩ�Xm���	�W�:�suՠa�~���	qD���O��c���n��j�VK���ɽ�&轰���FyC ���y� P^Ɲ�..�-�V�r����d�W�lZ�ʢֶ\����9*�y��\�z�h��e�WJv�vi�Yo�Ӌp��nx`<=W�[~y[+H��:)�t$�W�U@���ms��+��͌�Kf�>�xHh��^S~���L�O�θ��s�t�m���(�$s�yā��ւ�|�U/T�E�ݟS��u��������gNǙ�0��h>�3Z*�f'�jc�
��R����g��z��h{��(d3�y���:���޵$�z�NG���u���~kc�+��_#�@נ���U�T&��ž�M4=���!���9�����xtz��%P��z�Mz�y�����L��Z�x C��hMS���Ym%H~�5�Y�wӛ��Ӊ��������t���د��/Č���N�U߮�x/)��yn��>�xI*�UE��^zY�Ʈ���|J̡�?`���^�>sQ�G�PX!s�k�"�)�Η�#=�5R���髫@���]~|/�ړ�Y�.S��J�~��W�=28��ӓ��u"�5�h�t� ������:�V�8F�/ָ;�g�Λ�����F��υ>��=��u;�'ix_�,�W]�7��h�-|����_��1��)��[oZ��[l*"�-v$�'��3*�W*M�3K��ѺW�.��.��Xԫ���#��^��e�&F�^1��ecƪa��F��^iT��X���2+�M�%���n�t�c8,���ڽF�Y�2�Uhn�m��86��[�-��tw>�]Vc���;�\�hF�Εv����*���}�UЦ��L/t�I-���.��w��0���x��]ૢ��g� .˕�8�A�I�x�Шj�fj�h#Q����̣���ŒIR�uv�p��L)[ѪN�J�٤0hٴ�aM��w��F�`��	�Y��<�Z�~K{��,���M�Hvu��n@��ݹαnR��x:�|w��a=<Ֆ��6.�?�_��x���s��u���M�X6c���w�z�Hv�]�j�E�O�p<���y��N��]7�7OB��Z����$��f�A����&����ɲ��Oum^��騎ՙ�̓o�+�=.�R7��cI�� rÃ"����0Ѓ�7B�FW2yi�
�#,+{X �J�9��Y�X}t���;c���v��U�#����)j�R}�يc��������E@Wfo\:;vQg�X:c��8;+�>�ɺe�Wcy�L������m�L�Ҋ&��9D��Z瓎4i���Vm�
ύwm����b��S41������\�ڹy`]� b������S�5q�W��f���F���XTHj�uu�P
�,�h^)�N�j`��>��bk�]iG^U�������\5�8Q�����V1�U��6nIF�I��I���|g�D��殨��w$e�:s�D�8i�EE,Q��ѓ�Ni�s-�!s�"�x��]�f�.K�I�[;0$^����w���-���%}���m#�%XCd�1�N��$�F�ec;�Z')�V�6W*c�)�D;[�ȸЮE�v���v������C�eի�y�`�v9L/���˸��C�e��L��7���en��)�T��+3���x�2��I�b4��tL������6�RsM���]E+vw��LnK��B�������kW��V҂fl�Y���w�eT��M�ߕAp��@݋�++4��_#Q��B�שь�\����)�w�vM��W�x7A��7�m����-Xh�}��ɇ ;�[�6���pK��@��u9��s2�.��Nƛ 4�L�[a�������K�u`̣�~L�u��:�B\��v��Wa�AGa������r�n6��M�?��Y�����OP��R�e,��pNɹ�!O����w��Ol��Y7F�0
;��uro�6�+�Ķ�|N��w�h��^Q�h�Qp���%9ts�L�:�Z�z��΢tĥ����8r���C&u��7�)��G�]����9+4�4���1���l����mQӛÁ�/-vvԍkv�k� do��Ub��5�����e�I<�Q�ͥj濃�����"(��
�!��
0��Us1�E�*��\N0��Be�U����H�Ui*I�D),��b9,R�V�E�<Nry�
s0�BQ�rK\�UN!)p��ZFK%���e�9�*�J\�%b"i\0�H���"ML�f1L��M%ns�W�6�%W"9h�*0�
��P��UJMP�J�S�&�i�!Q�&�V���%eU��B�!B+��3����2�Y��GJ�*F�)	N����!U��UAf��b�ʸ��B�
����0��*��P*�F��Q�L�]��V�J�h�DU�D����t���1�B�$��4gj���Y��QBLMZuhTIfR��NZ*b�R�L4���JC��a�%�'9XW�@u�ʒ��8�����q�b�������<(R�f�2љ&�H�����*r��?kW��WST���9Φ73JyJ���zq[;�R� �����5?���g�T����n�!�{@�w�l� ����+�:����y.޹�<����'0�aYF?T�Ε�a|�1���˼�=�N�xxJr�e�T�N�{�w^�'���qYj�3��]9���T�J���΋����Xux[��O�E��v��VNx�g�G���Ez��Qmdq��,F}������nE���9�&�ġ~;J����N	^��>W�����'"=����ǽ~�[�S�
�"�ۤ.X �~p�O��3�=�/���<�b�s躦�{2⽋��^����o���Ͻ�s�(�9Ay��z(��F�sj}˕饡����5�Õ©�K.��ȼ���p�ιǍ����]OGaS6"��G�k��Ƶ��H�6��L��]3Q-ߤdI���f�y��Y��bC]Wx"'#�.�⽜��^�������T�z���U!�P%=Bs�ň�)�9�b��R�{"QG3�o��ڬ2��~���({�G���d�
��T�WP�}&ĉ^Us����4%����H��o�f!�v�ч�1�ܡl{���f�r�����Eф��	/��9o%�ΌX�1�q�i:{�:H�2�@���~��^l��ވ�1�K�؀*x�Z�W�ջWV�9�7�e]eN��܂��8�s'�:�k'#��m	7M�?C�-�`��MϏ�{�R�'�z\�z��xo���~�蛇��
t�GD:X���W��铵�g9���es5~T�����K�-���
����2��R7�Lk�g�r���'���ޑ�=���qq����R�7���g�n|��(f�\ϫ#��L��c�&�]xć��q��⣏��H�ʈ�(�ᒺ-�p��dy*��7!���S.��[�A[��*��̟!����ۓ����pӐ���r����u����e�Ɵ��W�{��vh�DL����'Xg�p
�߳��b�g�xuvUz\OWK��:{�j��'���錹�>�Wb����d�g,�>�Z��GE���l{�m>����=����$he{��?A볕�7K���g���_2�=[S-�"z�3k�/
����zF�~��ݩ�5�ڞ[TA��J1t{�z��Y]�牼W�\=�pr-]��}s-�I��Y:�	��[���s�~�>���f���_������*u����/~���>�Y�HqC}v+�a�q4�C/2��p���������e=����P�7��s]�=2���[�������������/F�sh7�r�~�g)V�{��t#0ā4A2㗷������F�9%�{��	 �M��5�� �<W�طI)���891���3ۈ0�N*,:�1I�(��@u��d�*V�)�Eq�n;����[/�# ��r 7T�j'���ץe�0�x�&�!��!	[H�_�62*�,�,�z��P�s����,�dc&� �P&|�9��T�+"M6�9}�y��o�{f�,ܚ�J4{���p�N���4<��W�ϩ�)��Ẽ��wJ|�;����0�=�.*�}s��O�t������(�ϼ}�T���φ���G�h���dQ�����KfxF?k�^�4�%�r�G�z��lc�Hx��2�I�o��z�q�]>��t���"������K�s˪�$N�$	�#n�,������spq5�����H����>=9왬Bt+�>K�+K���>���W� ̀��2TS7�y�k��ߡ*dd5�����̡���ݍ}�Ǻ��Z;�����y�=�_�b֑Ϣ��\%~6=�5�:r;�M�q�E��.�Y;�ފ�噉�{�a�w�����=��G�V�#�(�w������:z�U YQ�k:�;��RȜ��=���#Nfϧ[��~��Rgגz�n]�V��ݐ*����43�=Y��s�E��N:lq���,�����B��NW!핺lCh���s�T��`M|��?g{��%ۏ�.86S�fy�/`��J��e*���G�.j]4s_��7��Ld�]�u�����gNZ��so+g+�\tT2�ћ��֨��w�������ڬ.�q���yg�i߳�+��>W�'���js�n�kB=�==��uy�W˫�^f!���}-�M��LLw����y��r��Ԩ�C~�q�ֶ�ʪ��(Ⱥ���oeh(��s�����S��W�H5~�]��f�O�߁�D��{��3�:^5|Ձ��qp����v��u���r8�{�M�X�����1�\?:	A릗�Ut�>�gג���<,8��y�{���}^��� �o�^�[~yZ+H��B��2dy4/�gzA=;99���]��O:���o!����O��lx��9����/ẞ�D� ��~�{܌ܘ~���}:�b�g�����{L��޷��ߣ�ߘ]V8,�u����<���'S��'pV=��<wԴ9����M�@=��D1pP�g�"�^X�C�� {޵$w������{��L�#�������
�<&e����ME7fD��������H��{=�+C�c���ܻݻ�R=����o�\:��$	Ԧ�,���Ѕ?�Sp[��3���/u27<_�ْ����~��"�*۽��V_!b=�} �9Q�,&�yž�X9-N�[�SS��u��̵�`��ö�q�e�%�\��X8���-w���Q����Wc�z���[X����$�1cV2NK��tŌY�Uר%8�;�-Ԧ��C�Q@1���s[3α�6�� UB�}&�C��q�"�9��}/6��v��Iǉ)����4$��fP�m����}�\t��!������w�;��++=4=��ڼ�����6���fl�O�u8�R��zd����Ϗ��E����s.��c�X����+1�Gd�?E�����<T��:o/�[���S�I�{6A��ˢ��{^�^p�q	z����:�l�	�f"���E�>��4�24��N�;�p�w�`��Ƕ��q>��¸r�%X=}�����_�>s�����ꛙ҉��؁��mw�G��&�
�y���7���C�Q�_}�٫���SaW�^_A�eS�����X�Ϯ�ϕz�켸ʎ����b�|�߶g}���#�xzF��߂؋k#��ab9mQ�JC�ؑD9~Ѿ�j=��ռ(wy�m��E�rǠ��Z���D������[�[~�>[��G*��0�y1�����*�o?o�~�G�WY����ˊJ�\�3�{:w��xw�	�{֥��m@�]��q�o��E:��NA��g^ኳ�wmT�e˗G<����&�K;����y���c���6���/+v�s����bvkuy_�Ԩ�QS���⧉�s�/����5�7yD��)5����Hb��������9^�����R_�Kc�Z><G��A����ϬSal-̊�Ϟ3�y�{�����b|E��\\K�Ll���x��.����B�S쑀z�Lϕ_��}��~�6�f�yy�y�bB��ג3�q�|��W�C�]=�ʞ�U�W�1(���X�����)�9�#�~�CYT��U��i��6qxF����U!�� �z�¦��o�M���ʮNϵ��x�ɼ�;�=�Y�|�e{�`������W��Wx��q�.�Ej�����rq���3��{i��[�"=�n�nRf�*�����O�>~Y�9����L�l1��/�u!d*
:Ĝx��(Wq��o�EI�ςۋ�o�oey�{�!��5��K󫡏�2���zd��rпG��Y^�>(�D_yO����~� �$l�3�ղ��}�#��@��=9�[�a��DԞ�,�~���fW�Moe��{r��Unr���G�b��=�-���O�Gmкc�5g��D�Z��� �:#���σ ,�߳��b�d!���^��=]/"�lt�6�U��V\�9]b.rڛ2�S35Ʉ뱮�5���e�������ɺ�Ӽޗ�}o�r:���1�4��SZ�%���bn'�A��!�e�a9�/�v`�W=�(���x�-=�3A���!{)Y��(�9K��3�<	N�U$��j� �����gylzv)���GE���o�y<w��(Fvm�,ށP��n�(��"vV0��^�;�����[���GS�+�/
�����^��TE�S�k�<����Ϊ�_�9lv�x>����
��#�mݡ�e��{n�kv%�櫞z���_�O�;ٕ�r�J�2_�.#���>۩�e C�)\<�,W�6M0Yy�������t���1~�-/���a*Ǣ��Z7�[�eD�Uz@��yT=��n�:�.�ǎ�o!{]�)��E��N�CL�=u�#��4|oإ�|uy�q�w�I��_D�l9}�i��+gu�s�y�q=��趯�Y�z��zw�ϱ���C�ϣ���]�'(1j�W�Nb�>�t��sf*�%���$}�П}�I����gإN����;�9�=�Z {�q\��� /�&��{�3W��:[kC�����QZmX�9My����V�3��㝏W���º|G��39�b��\����#�[����+�j�W�D�8<k�6S@���C��'7Y��{޵#�LX���͔}J��s��Zù��%��S�aP9�]��+^?�<�jC�Q�Kk��� N����$/D�dr�tt%K�s�m�;}��Ȇ��T&�
�٘��HFC�p��L�0c]���3���ұ��v�̳N�3�d�}�|���"�'��-Ks��=?�ݕ�"�f��e�� �@�~V�f�o�ܵ�ljT�k�q�\�b���@��|��y�%^����({ީ��b�n��!�\6���V�Ϯ����s�v���N��;�u��=�=�r���B��P�D���l2=´�
0C+���y�s��L\��iL�{�H���>��[ �S��Nfϧ[���~�>�}W ��t���6�FGr����|w^,�G�-~�p�)p�}#��37�7��S�gxWG�g���ד�lS"{I�]��kö^�����)z��=\v
���WȽ��4�F'����.k�t}n�Y�y#:���3����{��i�3������Nr��r2��ʧ��Q�Y~�C>�N'�h5藑=���þ5�>k�	"��Y�h*f�{����oȓ\?:	A�i~�Jy�&�}��൞���m�sގ
ԇ�<=�}�W�y�x��_���$�jG�rav'<bS���Mx/�f/f�Aݺc=���ƽ��;������x��9�<�����)�_��%�YS^ϲ!����T��[+�ul+����V�M���{1����3�/|ν��(h�#��>E\ͭ�ݸ�*cT��8r�\���Ve����4���u3�9�=�YJ�)�˳��s�C���"O���)v7�Kt�iwr����ecڀ��q��h��E�c���{��������3��츯z��nO��:v<����V8,�Z��;wŌr
/cۛ�R�]�x���P�j�d��/�\2�ȼ��j���_�=��jH��e�6�\��z�������3^ *�Bf|�ǨHn��!��l\r��9�f��|iCѽ���o��݀��4o�g��39��|*�PM� N�������2y
~G��f^-b��Xw���T.}��6�ﾏ�||�}��@����U�k'i���Њ���x��\��F&��_��dg����~Y�#"~�C>~�D�o�\tY�h�/����g_p�3o�蛨z�����b�Y�~y��i��ܜk3eΧ�ʜ�~��V{��r>^ޜ�>�B����c��}F��X�u���p���+#Ǎ�z^����w~#y���{6A:�,����l��חbD_5>���N�ޯ�#e�OuC7��0]>��4�3�8��W�ư��F=�O��s%�����YB*��对CU��e1�?�?EDi�L/�ds>�7;������IQ�Z� a�o���W{�v�{�fo>�v�Ɨ�%��]
8y��}*j��t	C���+5����Ϙ�xڸ���7a�:#@wmW2��v$���$:
� �y���cu�L�'���d��qIkMخ�t4M3"���N#�w%y��ޥW�LtE���l{� �������6��>^�ò*���5FV]z�L��|��xO��PW��֢pJ�گR�q޿H1�k��6/���Yu��ˮ����ϠS��e?����n���3�	ž�}TP�:�����{޿H��O������~�>R0��Gn�o��Dt�Qc��r�8�z���b��Ⱥ������,[�e����#���>>�����n:�b��$�׳�``�x�C��*��)�6�+��g"��o=�c·�@����j����w<�	$b5S��ۗ�0p�f|��9����2$�a���O!�<�ȵ�l��b��9��RKi�C��	�
�w���)��U!�P%W�M}Mّ�O��8>򻊞�������q� {0x�~���cb7��<�z��޸�
� A��o$ؚ�<�옼Z �����o�<�����g[`�G��<V	9�����y`������]���)ɸ�6{*�&�؀>�^Û>��駂.+����4j�+�ʱ.L'v%%L��s'!\l���6�������� �6���m�h 1��� cm� �m�� ����1��� co���� 1���m������m� �6�  �6���6��m�m��m�m�� 1����m�o� cm� ���f(+$�k6��(@��0
 ��d��H�|w� P �T�!�E( BPP
��B��UP��IERJ � �@�H$�P
�P
�*�R�)�_a���E
JT)!QH*T�TR
$� �BJ�*%JkDB��$��"�����Q)*��T� �IT�(���mBQ@�l�S�������"�T�AJ��c@T
P�H��T��H���v�*IAT���R��u��IUi��Kx   :�e�T�-���5U�c�m��ZF��4�bEejiUFĘT���`�5���(CKk�6 @	Z�$���   �l�TS+5HUUfSX46CS�4�F�]�4QEQ��;��(�Eh���E(�E4Xv⎍4QEZ�q�E(�Ef�qGEt4��H�UR���(T   �c��;QB�6��T�icM���ԩD ��Q�5**�����VA�k*�ѕU�`ګ*����**��P)Q H��   䪕֬��*�
���4�$PƢ�����PV�����i���ZcV�;�M3���h�Pa����WIUU(1*)U*Uo  ���howv n�t+h��6�Ul��Т�YCWC��4�6�)�Uv4�Kj��f�֔ZZ`�V��l��Z�6�*��*RAR*�T� �  ov�[-m�i�5� ڣR��U��U���:�vk�c
�ke�sm����mm�U�`���t�wc��daZҦ�TJP�c"��D�o  3�K�M�Rƶ��hP,M�]T���0m ��M�R�41[kfM-�F6ШKXTAm��:u��U�����J��
R�x  L�`�-��T�=j���
�U+KJj�\�,*�lw�GZ3v4t�h��*�6�f�-m�M�0*��,�����)B����!�  w�H5B�H5M
d�IZU3R��
��������[�uU��4�Y�©�wh�P2��h�Ec
�T���Z)QR���  �]5��E J�*���Ӫ�4��J�j)�˵�`U
h�CU*�uө�k[MhV�P���.���@�`��SP��T��̪RP# #S�R��  ��F����@ �J�=F� ?ڄ�*�d�  !*S�T*4x��)�Hv�:&TLQ)�)+�z�`)%{W����o��ϝ�u�~���}s�TTA_y����+�����ED��ED�eVUS�����G���[�u��ME�U�Z-Һ�u�1�7����78nAX!uiV���eZ�!H�ݔº��M�f�'$޼��ub���>G�:W\�8P�q�phQ����L��>�2�v��}�E%����Ѻ�@�/ ש�u�e�1��^���Z4�3��Ͳ`�!�Qeh-V�ض�[#1h�m4^�G,?�S��$̦�e\.����m�������&��M ��V%=�F��%�x�[?em�Ɯ�H��RݭZ�Y6�4�-f�t�%,�-Miݬ��`�Ot�Z
�,Ʈ��O6f)�-n��溔̥��ݱ��4�ûh�$��t���u6�&��]HJ�})���׻im:h��m���y�Xs�'ib,f��uz�8%�Tb�B�݇1�C�3��,��\�Dd��锇�w("Qs&Bڥ�fH[�����fZjc���h김��W�u��՗�B��VCo(LVޕ[SͭR��U�Z\�Kط��>�CYi����Y��3[���$Mi�:R��Oe�W�l8��*`�Y#Xo��F�,�:v�N6�%�����y��*���[�0�W�g0��4=��A���#ה�0�\��h���Ѷ�	cf�=���^��^�mj�[�XWdg.�@v��d�KX���n�%Ԯ�x��lsֹp5x������5���vj �Eh�E�<8��u�(T�ڠ.�kKWf71�IT�-e�c�^e��	-�%�J�DS
M��H����`�O�P�լz� �r�5��w�%�.��Mm�-���t�$���R�mf*d� V&"�����Glukde�#sIy�EV]���B��سu%�8K7x��� �@S �
�U��p����.���oZt��ћ-=1�n$�m;�á<nb�[rټB�ۀZ*Ň��-&��Ol5��+zeM�L��Qo0cFe�{L�!R�6�U��^��i�'yv�d�s#5��F��f��Z�2���U`��FP�VtfY�A�[)I��iƁ�S�Q���[ ef�;������J��)��6=������Ʒ�O�����z�˾�b&`ԧ�]��ڗA]k�
�v�hVՓP�wX�]�w��v��i��bm�LVw=��Cަ���W���KmΞZf�����o�ֳ7N�\��,87)�l���V�z�^�am�E��ݷW�lq�n*vkv�	̹A�Gl��B��c�ISB��7]�9��O�.�����tc��� :��3��|�&՗\�H����҃��(�[��5�Kox��z��C7�c$�+�8[ђIYw��Y�R� �ئ�
����FJ�yAl���[���W�)O-!���^ ^�W5��0�A�`����!]�x�Lh�h3��U0�j<;u�l�=@�H���W�F�G��CU�MƕS[K	2[c�V�}�� �4�� X���-�V'�֊(b�̍�5��᳝�i��6��2��gNT��l�m��Sw�P��v�3��ͽ�J�^k�޼�����7��6SŹ[�`EG��qU�
{�|��p����(=~�Z{�'%��;�[� B87:�@�c�
��G�z��Xa&�3fu�t���h|^�e<���ث2��ﱕY�
��nI!���,kʕ!��֋5���E��5B^�� ��- ��ɭ�Tѓt��h3�KsI�h㨪��`�J�m�-��%��P�����z��Ie�kE�&��6͇��hН�S$CS߮��j�)6JˍK�)Ͷ������	6���wj��U,�ƦY.�\0�4�j��e<z�җ��k��䫙[KRv�)���U��pf�r�]G�ʰ+��i<0)��7��)h�ݺhn��ܢ�u3.�c��(8��32Σi�[Mp�t�Qx��,zx;�M���]e�]�0ff����9��f�Af4ۥ���xj�m��t!��f_��e6I�δ��k9��n�a.u��-)��G0Jf°
˧Vݢ�و�V����
��F��I�F=O�p}&�t�u�*cXVOA|��~;���������uh��tqj̑�	��1K L�m�$�ۂTvŚ��,Y���j��Zl*�VO)��e6�b�^�OBcn㬄@��`u8�h�\�/���J�����|����6�Gh�oE�z�O4Q����l�J8��,r�,[�t6��z�1s]�c(J��u��V�����uq�� ���K�+u}77F�+/Z`�X&�	˽%>���7G1�]�,����)괆�`n�n��֩YN�W��fEݥR�9�
[@���ۦ�o/l�GL��V�T�nܔBʾu�fwkC\{�]��$�ꧤ�b�PL��)
|����D��X�oV)��&��]�B+u���r�&vP:��e�{�eK`@�7m�mU�&���ݨ�E*�=���J�I@�w4l��sJ;wDM,7jnێ�k
N˔wH��b�6P�Zr�Wn�'��.�k�D��4<v)�����[*�4K�4����h�ض�_ʁ�֪�}��Zx���B�Հ�Y�4����9�KK�{{�E�%� ����vJE��e�mռ�+v�Ml̪5
S ��d<# VL�F�kb@��J�.eF�L��EK��5"��5:�fz�j��62�ټ""q��7���R�ھ<&)�W�C� |Eh��Y�6>���h�î��{��&���8�PeZcS1�UЦ�V�m!r�Ӡ�8����4(
x�$�"��(���؀3˧��!���E���L�`��g6Ό�V���,8t�&����_���T��
�mm#�E=�]r����P�*`l"�;�1z��sUX{�����GF���i�r�Be`��,�k��:e�m��HT������n��zEdE*��XoEL��-�[���:�®������%�����Zx�9��t�0t�mn;���9y��7]L]���A:�������v'��e����A-�춈�������6��0"	U錐�����N�va�c31�պ rҧt8��]�t�U�Z��ڬ'(
&��{b�� �z�PN�(��t���6����F*yLE�oedh�^̡$�ȼj`׳`�2��^�ы�t�]:�u�)V�K!�e�Bs�t�ZL�Y�����J��ۀP�K�+����i;���xvIǦڻM#��*A𩹋XڻK�h�@V^��E�X���:��5uw�x�SUŎ���ٹ���3X�(v,��Sf�ɹy��ؘj��7�/@��5t�%54^R��[[�dT�[$u�C���ie*�Tq���7�)t-?G�wR��j˰�u<[��[����e��
���t�ٗ�0=�k$�(���� Û��Wen�]=U�U�V�v5J1�8by[�R�<ɜN�	=��+��=����+�%ʺ�WӘ��sB,kCO�X�u��QbUʗB�R���k	P6�=-���g,a�A����hSײi�4�X�*�9h+�1��2�op����Or|��h^���-T���V�v�H��^�i�);�s)*�D���iK�dՕ����W�M�l�m�;v�C�^
H�ӈ-$��r۬��I"�eEQh�-�$K����;In��Xb��>LV�R]Ӕ���A�-���i1�WYV���]\�R�Ͳ���Q����N�Qab#f� A�q츁Z�iÒ���2�0�{0ei�Ш�-�MY�L��Ԓ��J{��Ҏ�����U���`�H'�i������f�7[���m;��thU�繼i����*٥����N�e�)}i�1m��C���.��ܱWE���Sk.�VȆ����cL��n]��:�f�]���ͽD�n��9��Ӯ�>��h��Sz�=����;r�i�i�����AJ�����V��(:ݕv`���)ܱZ�� ��M=(f<̤�aX�H �r�%�.����z��u��kW���L����f9��R���ݎl��/6j�;y�����n*��v�&���eMrȶh�[VK�+p��GXx∭;ks�Ԯ&�4���[t�+G*�A�M��S��lQ��l�*�Ct�\�i
F�C��a�*f�����I�ݺ��X�6޴VYʩ�;�S�o �Y-[b����L���\�ڑ�82�(eL���v�L�����G5sIQѣ(�]��	�[S,̙x�$�T��LB�hZ\Dh�P�l���6_�6Oa�U�In}x�u:܁	�)n��5�����6�v������O� ą��Р�Cf*�Bb�Jn�B:�5�1|E�����in�F�&�X�j<N�i:Y��6�a�6�7 ڻ��P.�
*��i�YV�b�U+��S�Vij��!w6��G��Ik��2��ю]�q����Zu�ʸ�$�R��[�L�'"���F�L̴�jŢ���t.�Ф:��'N���Q��۰� ��.l-1I��;��VN���I����{h�4���F��m<w�Pۼ�3#t㱖�2���ܺNL����9���1�C&���ב�{f\�1�J�dX6�V:MM��6���#X�HV����DF ��h�6yjm�)��wX�k)��i��5F�̭
]�b��SK]���M[˨D�E*�xkYR�Y�Q�����/�%��9��iQ��-6���"�E��(m剡<N�Z,�W�-N�����p̠�wb.fU�ˌ����6�b1*]$"ס#Oi������r�M��уv�WP)�6e1���#���&�'2���,�6E��j�/h�l�����N�m�p�n��osi+8b�؍�3�S2��B+{�ג�Q�ۊbvC7�FQ]�fb����eL6Au��Nf��6�oڍ��SU������Wcvp�\l�-8D��b֣��[[yt�8X�n�>��1,���\�Æ�ޏ��@ǯx������.�k5=���ض��.�V�������]��Ф��Q��s5�j=;K!�v�jYUf�4����v��[��FC�ز����Xm7tk�T��/u��ݗ�Syկ@ ���X
�a�*�+j�ɡ7fG��׏m'�Y��և���w��f����J�]J�F�R��ݸRnT�r�N�f5Ck5Q�m�`B~�/>�8:��S�#Â��i��۳��K��L@�yt�okm+|�%���M�`���CN�8�p�5�Ǵ���ؤO�ZL��HJ�GTY�lRs�i(���o�j`<�"�pn�ٕ%����J��dh|�a�>�D^`�H������i��n�c����kH���s���$y�]ɉѹL�$vs6�Dɭ� �2��ݘ�)h�D[��c�Ա�!�x*d���;���m�,��S�)Tͤ����i�j�f ��z�)��m��g`��d��8��ø[d
	�������W�аՋ�lZ�^?�A>����pĠ�b�FY��S�l���l��AV�8*q��^�lV�>{���aU͚]�a�zv�ww�č,�ۻ7I�C�[w=&��l^#{.*�^ 0^马fV�ѕh"+0I�Z���U#,:��Q饵��w�:��/j�����JD����ef��s�������Wق�n#�P��O4�	��iB��͐�t�Z�!w��:�J�P;f�	$��ki25<U{ս�����r�m���X�˛V)��mH��3b��M��_���k�w^�O8p �\�j�#I;o�]����mf�T�Z�J~x_+�'�/�$���l�۠���IO/6jtu�a�)�%����*��a�8b�J�Vնp��r�̰�6E^`�S�m�M�u 
�Ac�+q;U���l�%S5�������a���op������T��ZNc;ST{��"����"�������-s�y��*��W�K����M���O,�wׁ�\+���պM֌�t�ۼ]kˀMl�µM��(e�z�nFI ����~�{1ռ�*`mn
;"���5y�Ea0Ymd�WP��@��ܔn�4-̨�c�n�aݩ�,,�EE����gŀ���m�#蝬�t��
���zñf�����禎�뵪����6f��oPV��-1���e� 	�2[�y��*�lk�*�#�tc ��1�qi��f�њ[-��V-�6}lSXpL3㛕5;c`� ՜��M�cQ����M��NDU���ດ�^a7W��4q�X�d��o.��Y�����ʺh�nnRf\�kSïn����wkE�]�5
���~s��(G6nL+��i�v]Y)�e�\3��?�q�9DZ�gS�2k�(��-�J�L��J���
���m�N��`m諙����˥���m��qތm&=��VFw(ö�ٺ���3��h�R����(^ ��n|��&��NnK:w���4w�h꛲��Z�f�Ԯen(����߀�61YƏf`������$�|�����j�C>8l�!I)ͩ�Z׵f�b�1Ǚ����Y�4:��6�Ԉ�1]�$�La{G�x�N��F�dY9��r�;N˧4�[�d��V n�:0��1��5j�;(���,����*�݆¡u��>�1+ǳi�G�C K:$s5V��p�{t��T�eمZ��۷9�� ]B��Z�n<��.�6�-oڤ�tf��$"��-�&�Eꐩ�K7�)Y��XZ#wS������qg�o�l�ߓ���o(=���u&�w�jc/E���FY�1*yp�,I��40�i�K��l�l�/�P1�XS6uH��)=o���0��{�J�CʈaoJǘq���NM�v�EL�IIb/� �a��G˜3�d��L�Dv��"z�q�[#Ux�;if�Zg.�Ou,9�8�7�:��o"���Z�.?]o�Ivti���^է�. o�mY��	�6x�a�39�W���ZS_P��)_%n�kL�0FK4�r�7��N�� �Í99=��j.�������&�j��ҕ�a�Q�[B�{c��j�Z�I:e%��_Eՙ�ˠ�멍��s1 r�� mZ(�׻ҵ2�@�-	uQY�u+�Y��6�ʵQ�غ�y�Z�d-�q�&=Y��Xl�\�ۀA�`)���]�h���u�3-�U�T.��]qv�v�u6Zov�%�X�j���\�qP�(&癶=�����	Af��v��27mKb��RZWrOZ�%�:��嶥���r�����!������:�'X�h� R�::��K*�w�aS���"��H��<��p�Lo`�͢ƛF�TH���\��h��ʧ�Yrmu-O���T�n-�w��v���Ljd�DP71p4���h��E��6�p6���6n��&w
^9:ޫ��5&ӵ�r*�;���-E4�ǵƳ��i���{�4��-�m�!9##x��	4��z��u{7;�+�j�H��9�i�Lo%�tG{�Z�D��#���O���H�Ys�ۭ-]嵙D�b�e�/K�j����R��=� ̣�V�oB���Wr�:噢���d��|���Π6�|����ʹ��'^��	��Շu�y;��o�P/6m�����f�R��S�i���2܂�k�%��7\�.�ј�r�Q������V�+˫�X�%�'J�O(���C�>:X[���=��n�O�����A��1F��G[�,+�n��5ْ��AUѻ��\�
 �xu�lk�Rv�k�i���SC3��zN�lہ�J�ž�;�5y�+dO���]c�V�n�q���kp
mDĠ�󺂶��ǹX�i�]�.�:ɏ������IWW!�cCy���wAx^iG�-tΣmZ��i����QC]o52ȩ][��3֐uc�ھ�Fv�8+��#�;��|j�Z�b�z��t�r�E]��ա�U�ubۄҬ	�LQw���L�MΛ�ykk)8BL���p�B��S���,P�]�EIg*"Ž+뮘�n����.Y����HܭI�;zn�3�	�v�}�1ܧ��m�r\�;�����"�֟ȪE��6���%��H��:��ʮ�ە����[���SLd���.�r�z��L���k4z\	�)��v��+�qi�5����pS�Lͻ]��@�Se'�����m�o*V^ڝ:�ݒ�+�	�t���]S*6�,k���TM*̤0�\p�����0�q�HD�N�+z�,��e,�a+��3��}bjok�]7:�t��"=�w�Q�[����]^��uj	3Fvms�KZ�ᡔ�ZɊt�:�[��f�䌚��k��.���ubn�v
�ou2�9�{:E�;fMjh2�B5:1w��jnT���q��kv�-��њ��N#n�pN�օ��̹R�F���7���z.�vJ�hb�����B�_�&S�6�8o�=KMb{2n�C#�g27h���v�!n����ާ��.*ȹ�ݖ��JDf�Ư4����Q�8oS��}:[y[�M�k��mۯ̷bWO�g��9q�sw5�ٖ��?�Ru��bY���v
Ԁ�}0�.�]�f�ֺ��F��-���X&�3��-��ڳ�t��2�++8v+�c�6���o�i��ʾ��<�Y����"۝���:��u�w:b��m��uuŵ:d��-�o	���x˙�ż�c�ki@b�6�4oJ�)t:ղOv�t�Mc�z8˥�ڡ;�'K@d�y�=K��c!�*��ل�`�v��b��fD��#8L&U�\lTyh���ٝ� �H�Vz�����>b�'4:f�1(��̐șUǈ�G
yݴ@#�n�u��;+1�DV0s�f�V��\��l��
�����@n5�
��O)�y.����:n��`N��Jڮ׏��y��Y�Y��cfem�[�"J:�q���@����,�R��/x<AZ����I��FV���������vV��
�8R�YZ(_m���:7d<�V[:��Y���B}�_qT�xe)נ`�NXn	�1�d>�����*��$�)fʉ5KM^�M��ʘ�eoJ5c@��!�ko����ǜgkyH�R�U�~jŏu�e�P�mF�#�`u0�P�������XT�{me>8�0�S=r�Gf9��h�I��vU��"�.=��cR�c1Ү5�[��ջ�:�y��8��ue�8��Klʾ�r��5�֮ff:T�e��i2�,��7P����]E-���T���k�m�ɣ吷�cp�F`5��]���A��I/8^�ֺ\C,�5�nj�S3z�Ռn�I
Úm����|۷|Jt����v[�/vMz�7��+/��+*v����Q��hfs���S�z�T��9/t��ٮ
V'l�1�螤&;�J2�:�f�L?����.	���Hâ�n�7�)"��+z���f]9�XX&U�з%ݻ� ��J���+����	k���2;96�a��J���)u���*�`e^��g&š(8���s�iv��s���l��V�,�ik/E�h�5�q����a���!��р�ߚU1O���9BL`�j��/��9*�.�4�Uέ�%]ZύK���}�4xx�7�|��OL��a�-+}i��3�-fE."�]�`3���
�;ks"-j�д��+�;+���t��\y�q�Cc��bn�˲:�#X��W�[
\��.ehK+P�B~�0G>�|j��ST`��\fѹ6p�&PW��t����8Ի=��#�6K�z�p��k�:R[1m���+��,�s���QU+�&�}upcͳ�\��{MJ39�z2$w���v�܍���5n)ڝ�%�]����ޱ�����S9� tf���0j��ӎQyX�ov�����1eD�j�(׎^���+V���K��e��}LV�{r�,F�IV�J�z�4IW�拪��%�]6l��F�d�������!*�,���"��[�*a�r�`��5u�>e]�@���TmM��ܰ`|�J�����|n��n��g4q�[I�ƥe �D�`���=� �
�R9Js�e%v��u{u����7`�g�؄&��]1�V2>ư��L���\�6�u�Ӹ�������u�����R�MW<��V��c�h|��R�ǵ��+��uʊ��m����v���̇V�c�M٥KE���ו�0�ul0Bx��ۋ��珶������V�����T+FE86� +�a	��Z��ܿ����J-�rپ쳯�ӜH� pfۻj���9���j��hmA�*i�D,��0Q���v��{��F��5���3�MY����ީJBlNy6�_^#���'��]��>�TT�D��E��ζ�]gơ*���F��M�V���/]�x�>�>�λ�Cb���Z���a�1�/���_�SԽ�R��n_�ٿ�'vXP�����vۉ�R�t�e9V�7�����+��$��p�չ�x��oq9��=�d�u��<֓�H
t��Mٛ�L�}��͏A ��25b��*���v�s�J��Fu��D���3@QF'{�XA�)n�i�K�ظ�׃MjtɊ���|Oͻo��mfY�9pʲ�mCy�5Dr� ]O��L�suT��v��]�5V��ݙ/�[\ؕ�r��h�/�)�۵�@���ڧE��|Ļ�fP�����T���h����l��.H��h�J[�T|2�� *@si���z��ɐ�zU9ft����� (��2PӁGVڽn�G���2������$��N�6
$�4W��!L�aWvD�f�i��=��|]��+�R����N����rک������$ZX�wٲ�t���X��:��	oU�z�b�9t,���Z��(���%aMk�������+:�������n
yO)J!J.��:�d�M+�s&ɘs��jB���������P��V}uˈ���7*��#�j�G�-Ǭ�7ip���Jl�1���۹nŚݮ�Y�m��˦K�.Z0�Dy�n<�6fE�Ʀ X{
-�!I<M�}����6����X\�C��n��Txo���b]z[�F��� ������r��&�%�M+��vQ�iA�ӮlWd\&t �%X�[.w9�4q(m35i;�v����X�_^�
���r�S(�_|Ǝ���u�xf���Z��g^+��0l��k3:��]��;)��� _m83tf�=�c@���͹��I��R!d��o���N�J�-7�jm�S-���]��Y�R^��ubI�%P�Q֊�yW�g�n�HT®:ֳv9���wZ�;���X"ʚ%��+]ByYv]bh���E���}Lv�	�����,ձ֭6 ���]G�q
do=3���5���y���0Y��"�b��#����3��"cy\�-ĺ��M\�ላ��(�ɐj��=�9"�h=J�iB������O��X����[��jȀW�O_݃M6u�Xm�i�.�,�cX�<��(�s��-uܫ��H�nZ{ӏs��������- v'WuxyO�*C\���xG&2w#�>[���/ZJ���xFx�+x��;|�sE,�r�����c������3��+��4����اb��� nS��а�;7����k�jʾ�2��4-ů��ť`�OS��@ͨv�)mإ���<���TQnd"�J�U@eٕ�v�]R3-j��{n�n�8�Ȟ!$��1l@���I�TX]�5��S;Wu��۝�����;M�s4�[:NֈB��!3��+���u�{�(����V'�{���#'A�d;�򩶺��@�^fU��������ޔ^%�E��.�v���n-ӜfX꼏t�΅��Vv�q�ަ%�;,]!u7�oOA��l���F�YY{�kS/!�����`H谂�]܆���.�n���.��0�>�L˫��uYjXC*F�n�c���|�-�b��N��+v �jN|�H˜2���[��q��u��XM�;V�Q��6��7纰b��I�tV�3�u��'��k��ݥ���80���,u2�kSg@�v'�E%�趹�F��R���r��m �����jd�))R�9/%��[,�M�HȯoE�f��mCA$g
��s�s�qx�]��~ʶY�.��5���wkf[N��(��z�
8����ǅ���&�Y��"�t���uy��o+������KR��e��Y�4�xP��C{o�rs��$׀7���_�٫S07>ۼ�H�e�.<���ٸ�̬�>{\#z#�����.�Y-����k�5��ms���e�7y8�L��Z8�_���&���]oRַ�2�;����G��k�ϱ���	�r�xB��U��<�l�w�l��%ޞ����1���n��w9ъ#�Nc��6�fX��G&e>r5�E����tnS��&ogk��&m^p��@���%���|�C*ݞ(�Yf��6&��j���I���	�v^�n՜x��#���:��f��\]<uX��&N�t*�m1M����P9x����D�O=��m6�'&˕&��B͊�B�
Y�.��/t�V�Q����K�W�%��.�1O�07�7��h�Ec,ށ]�!ǂPZZ�{:�1S�wbw�8x�Ga�V��*�S��������n�yB�G����u�]��Sj���q��S����1��Ut"��Wnl��-�3����h���NK�o����n�t! H��g,�X����*덬�2�V3
�m�Z5��`�b�q'wh%�b�-qu�*��_.R��j��dˆ��=�SE�Gms��c�5�Ju{�<ʣ��d-̦5�,py{uV��P�lCz�Mj��ҩY$B��L���3�1�m��Rwp�F�4��]BⅮ)|U�����}��v�?��gW;���1�p���b���s��ܾi+�s�3+�&��j����o~��b��Nܖ��:Q���9t:���c��p{+6�:Z��<�"�{�k�,7���i�Ѩ�i�,9����t󟼞�|i���O	�r|�wH7^��tD�ml�1�wy�]�F� ���A��ϗG��s���	�T���3��|5����!��m �ʏ��V8�ZT/V�rR�*�ꌼZ�*�u�]h�m*�y,wY�wdm�u*��Rn�Er�ks��È
޲jV�X�a,|1����a:����Ұ��w��_q�F5�h�$z��.��,����<�v����� �9A��[[������f���譢B��]�o��+5s��]���[qS
��)��Kz�=b|E^A#ɖ�s�5:d�gC��/��G5��}/D'�CYX2<���e��L͒ҫ�o��d8&��=��:��Q6*$�\�x�EoU��0������n�'��'`�x�O}O���Rݛ�`�������u>F�E��+'hq�t�o�}eS��Y��̾�%M�Y�_�7�`ö�2��u~p��ݧ9����O!]�J�{�P�k�<�X�[�\F��-^�S+�� �w m⮧��˛b�?e5�N�	J���O#���]�)���ċ��S�����$�B/�'Y�ҝ���h�(����|�Pݻ�⏻.WbwEsS���s���Mۧ��*���a*����� ���L��:x������ߞ�@QO��ED����^��'|M�Y�?*���V!X��}-<��5���q*B�����}3��,�c�-\1��>��t�J𼌨�w�v]�F�.�h剹�����2��0�>/�0E>J|Ç���cϱ�[n<����[���R�)�f����1"r�@��@.`�]
3u���m�,՗�E$�A7f�H���'sj��QلAԥ*8$���`�K(\s��u1_��p/M]@I�G9����F��V���°�0&y�ֽ��}�E
���hbb��=�4�#F���Oaܷ{�Gw���J.V+����G�J��c��@�˽�iu�|�K�:��6�f�h��3L��j�h����.tq��%����&ֵ�Q��yt7`��gP��yHLwQ
=x�� ��r���B����шou�cT[Y��D+	��۶�m�d�WC����dS�S�XXp�,���Kƫ;B��QR��$���jX-�@�&S���|aќtŗ�֖8RF����9�z� ��G�����7e��S<q#�5�d^� ��N���2�����;zF�hv�Jn>2<۟e5��Y˸�v):�����S ���I��)��CB[H
�Y��&��N��睄�L@��!C�91դ$���+>��sep���r�n�����"lįG)2�U;0R��e����-s5k�@*�C��ٖ+e�m���+qV�Wv:wJ��Ct�! d�8�E.c�f�BM���N��y%��0_�"6���i69�DH���!S��,��������{$���e�/=z��Y�HsO�Wγ�����m4��x�{S�_e�]�z���\v�4H弧�4]E�Ǻ�ӞU�2�e8��tg��9�*��2��ӟH7e-7O(��96��kԙ�j�Z=f�i���&fj�\�<*��� ^m3����e�YR��h4�8!҃Z�Хh���ZϦgSp�ㄾt�ׁv��c�l쇵�
cm����5����d�'���1��՚q��g;=��h�)]h�S 1h4�W�╺Ú�{��U>!�n�Y,�p+qᇜY{��)���*9[{SK�}�KB�b2�e��ܔp�ԋg��;�+xU�oC�WnX���ه�zt0Gݦ�m��O�9����B���VI��]I�Pg	N�����(��-ӗ}�C�9R]�A^�.`�˥��}��%��T���B�*�;3eDZ��f׃K�E�-�2�V!���:�C�sx{��G���_QLK�LU�*�ܹP��N�'ss�v5��'xp�ѹ�4�0�Y�<���
��Wk#�&�^�$�G�v*��}��$,�/GH�L*t�����Z]�яP�h4ho$������Ź�f��-�=ٶf��sI�u���oR���U��r�\����pe4*pG�H�2wIX��]�aۨ}�n���JWt\䓤�[�Ju�*͞�*n�Cu�b��M�Jk��Pѱ��Dm���^�L<%��P��x��Tݺ:���e^��mK���N�&�b�n˳K~��҅a��idO#'�v�ٚh:j&��+d�VN9��j�x[D�w��F�^�Y�[��*X`x��m+pv�M�̺YAP��r.Yl3l�����ݧ�v�L���;�Z�,�m`u�[���\r�Ђ�ٛGl;Sk@2��g'�V�Z5�u��	e�'GAc��L�ks-��c��jRWu�l� �{1�'}e�o
��0���C�l���e�{��+-�T�y��mmo �ܧ'mۛ���}�=�Nt�=V��'�. ��k��b���A(2{0Y4�=�N1V�7su+E71;���t���Z�n�2���(�9ηz����XʀQ�R��9�ۛ�;.�j�ѕ�RZ��\E���\����R�>�1�F�9}�y��>���[�m!�vVV�&��mE�׺eX[T�΀��MZ���-j��sn�y�vK̩ˡ�E)��k���d`����<��$j��f�]�j�n�j间��$��$���m�O�e(K�x�R���9I|�8dV�C����W�Ø��s^M�fh3��v� L�gu����k�aH�;rI|(��%�E�@�"A�X(����2�z7��Hc5�:���+�ۂ�".w5:��a��z7�Mn�!�Lث0��j�mKr�`
�ܵ��=V�w�ވ����g5:yk>f�"�}�����Է
�}ZTU�\Q�+���Y��{;n��r�ܢ5�8UgP��OuG�[���Cöe�؆�y�]��M'���8���,vih�Ř&@�B�M�{R��>�e�N�7�stE�4
e�Tmfn�n؄v���7��;B�Y�m	�ƃ���I��6k3�"v�����k.8�.�	%q]�!�g�Y}r��wp�+�Y���#�N֍u��k���V�T ���{N��^:J���}�i�]�k@�kyN�t^�GWdp���̙��,A]�Q��4�;���h��w|���6`O�~�\p�I�<����|��޾��OR��օO�͗�R�z�ꬠ,DGL�^�Ԭ�wY�n�th�Ħ��r�!��Z3�����0a��[#����n+����E1'2IV�[�G5Z�{�[���P���RuLAr��R4�h駥[�wë7@�y"ޝ�!��i�N���=]Op�
c+kD��m��,%j�Yܚ���Y]t,ܽ�&B��}I���ͮ"L%mmɃ%x"�`|����/Q��d�EWc���e�b
�ʆ*���D��gv�}���2m�\�BI�[��9���]���+6�ռ��V�N�}0��V�F��:M7�T��qX��*5m],YAm�WF���T$���=n�`Vm�\�ܻ���X���ݑТ���^N��k�?b@9�3c#=J	����`�/Vef^��n�	�/��̤�瘬�ˉ^��|n��aH޺o[��g���S����n�uq�D+(�S��銬$xf���*���kB�D�l�.S�\�&Y�lS��SCvU�	wۃk��T$�.��on�����8ђ�P�B����∮8�R��C�T���Rr�R"��c��![����J t&Qk�^��)-PÊX��ePC.Y�bK�a]�hp B�]}:�օ��FͻA�W�f���6-Dc�i�'n<��F��9�6�8�ņ�ʲ�TԆoZ3�If��3��y2���blz�^�:��%�P�{����DQ(5n���ԸA�tث���"���aUκXX�l���jO�7܆l�ib�%HT�&V���%r;&W]� ���M�Ī�ؽ7tZ����b�U]�K}�÷/�Sh�E�G=�ue�@�{��V,��fgr�s���Jj�����z�JC]8�];7m�o0��[��I��`]2���L�+���p¤�P��|���|�k��v��o%�P1gL���=1˄$���%=]��&�!��1�W�a�>;��y|kp���^�_
��첖d�P�(��u��˷f����sx�FP��]��˕3CW��T��!oi�К nu\rl�x�+_*}��w�ǚEʝ.���� ��$���T���x8���kN))C+)�w��;t�7f'��v\�j�������P�d����o5p�,@Ա��N�]C,��9��H�j��72x*�<��8��f���Q�kz��O�;,c�,t9��Ԗ�rn���(e���oy��j���%�
Tsk7��5G�����"�l̛p�l�c��5�V��ݡ��h��W^��Te)a�:)Wv�	���o4!�yN�T��X�� ��yZ���Q�Gk5嫝֑dv.�F���#��#��5��v����<�N�볖D�V�܂�	>֌��9ا���m����uq����S!`<�,�{J�#�o��3q�e�ұ&��l�yB�M��n�w�a�x,�!��p/yu��sΏi�f�}�pt�Y0��d��lb���( \����I�`DY5wc.��x5��0:��{�mM|*<Ů�+�eZ)����u.	���]�&WXV�Ȓ���gM����ٽx+�geuhD{�T]/-5����P̐��sx�Mú��/Z�즷��ѐ�~ӭ�+nN/�/rL��Q�V��R܄�W.-0�P��f:W�z]�����;I����V���@D��-�t!����:��a�,��Z��%]4;f�	1i�N���
�q�-���]4|۫Hk��\7u&Wj����q�FsZH���$E�isΧx�Z�e�}�cǯ�6�ō���gP�����!���e[� ��,�J�pKCq��m�!c������i�D�õ�6��\��`
�9�#i�T�(�)�;Yg�d��kdQ�����`
ľr��h�*�M��`�ɉ� ��u�d8k�=���^n��(��vB{�%U��)�*浏/� �nʖm��u��s#�34CRśg�AR�h�q9�(�`�.��ޣ�R�AN�F�WԠ���.����� �����[J�k�G5_��#K�t�m��x��v�<�ZC:��-��GtG:�X.�a]e_
s�^݊8�$2���	Â��b]alPt�
,�]!Q�yW|w6�W{����]Y�R�y���W\�����U���ؙ��Ź�2R�ʨ5����=t��*^�P�Y�K6>��f���)j	�	�m\�5:�%:Ol_.�����2w=yߵ��p].635cf�V�y�Y�.��I�q�.���Qu��̭Ȼ(�'U�����G����v��J���^��30P)�9r����.��t�;ze՛��S�a�}5��}��|�:�+;0�G)M��oy�ӹF#�FN��j��#g35�Nm��z���7�8mqu��ȭ]�����>�W���{���%+�����g:x�=0�q��"&������s+0�����*b��Y��P�G�L�U�
l��䱝X�R���8gD �n�@)G�S�n�6YO�ɟ5����]��3��!�%xS����}A=�.k��:�c8f"��|3c\]�h�'d\��vM�#��)�6�j�٪��֝0�Z��S&���N`��}إ����g("��8����> �7�߶��C�ɨw���k4�h0(9���bZ	6Û�
�w���u�E���'��ˆ����*���7�,�w7��%�Q����9�j�[��%e���{dp��ƍ+�h��-}�@;�m 9�C�Z뒀:��J8�˳ukib�$;�L+v,�"�$2�+A����;�H�c6OsC	�j6�_�_�鵈�J���������+Y��HY�"U��0tN��bp Y�jH�M�l�������:0��2�s;3�u�o�g6գ���mީF��X���E����;���[I�>�鵄�%*�}�0��8n�i����gW���MV:]ǩ��$`"��n��
g ���/d[�s�έ�\��E$p��*d �KE]t�ty���f#+@��t��a��9Z,�]�pޛ��+�w�Tik[M[�d��z݇WM�7�Jc�Q9s�V����gs�R�*���GKt^�0���|�{m�!�j�2�	y40ٕ��N湛�������啙7V껨(),	�nu�[I1v�.�7:��]���}fc�a<��SV��n�ݫm�B�ղ-�ʶ�kMs��)�X���\�c�v1ug[X���FV����-)N�u3��r	��6/HV*�>1��Mkt��Wa�F��z�nl����`�u �4bĮ����-�h�sWЛ�xr�P�e����)M(3�7�u=RpL���P���x�W5�^Vzd,E��G������]Y�5���󊳽��>����Gّ�ړqή{Cu��b)-2���ի�F^tEq��g����	s��ldf�	��jW%�UC��j���*Qֶ�VU�#�H*zK�jgm�Y+���Ƹ�]�&Y;[s�!�^��{��z�%
���6��	]I��ųs�����S���r��W�K(�����V 5Ȟ��ڠL;�MY��M�b�k1�&i�+��,�|fsP��{��}� �2/�[�T��j�dev񮕟l6!�-ừ<��S2���AڧZ��7O��*=�h��|�ݤ��VYx��s�H��I��I��ttn��M�ܰ��'X�\v�I
��έ�b�
�Q�n���'���ގ��Tů�8y�4��`�`��A�N�|h7�B���z����2nv �lT��벵��E���U�3���hˆ�U�M�L�'��vt��VrOe�58>�ɨؙ�����[�ȡW$6m�Z�-:���7/��������怵�/y覉����]	w��Fv�����ݾN\u�� �Ǔ��m[�-�i^��>��!Ƶ��������$�LZȚg�V�eD.���ܛ��l�-w<A�l�����E�n���ֲ̣j��u�0
w���5�CVWZ��9k�9�}�GT$�j��A�$��u9�9+����b���|&�]�0[ẇ)9�;&��o����9��6��3�z*���77���{Zx*�#[�&R�(o/s{�X�Ȓw���8+9���+��P�B����	,;�JGp���B�6�C0g �̗�i��Yv�ӝ`�'u���9�Q Q����rڭt)=�)�;�2����)V�&�]Эdj��,��_ejƖ���>
�&��ӆbu�:�t��<�u�e� ��r�W_WI]��2��gbҘ�y�V�r��hW���eZ�Er���ﾯ�����������|F�
��I�Jl�]X�ّVVY�4Vd�h䌨�m]>�,��i�.���ƃ�U�vu�{�f�u!R�\ʷ]���;VL�]8f�@sMͺ��F��Q�f���ζ����,�kd�NG��_<��M+�6v��v��]��od�u����Y.^��#�.�΂$���\����P`2���XMw��o���r�%�L�C��V�FZR�3
D�:�D�q��WU�k����,+���t�n��v\+��L��#H�X��е���ܥ���#	��vXcT9�#ۤ�X��y��嵳r���֊��Xt�3�КDq �y��+Z�(E��y����+dV�ikZ��+\�p�R�X�IQ\�3�f�x����J@�o(�JS���OH�4^���zxl�q%/�gp@�% ���3-�u�d��*oT��QI�q_Xé�{�f����m�/ �h�+:��TV����
Uj��uՊ���O[��LK���Yt���X��+t�j�by��>�AhUs��͑Wؗ���v:����:����]_�,P.��-�E��Vɻ�<�ck:_�v#����I]��4��%�܎'���{�#Q�V�ߙW�7y�s��Vډ9��ɒ�u�&l,�x6�[�1�ő(�[k/�`B��9�t�g����d!{фz������K�[$��A	"O��H$ͣF�4��mcSF������֍�U���[Zm�EmZ���bc`ƱU�ͳ[uM�MD툂v�A�"�1���iփMR�DPU�D�U%i�US��lj����j����tl�T�EDT�4m�������64���1S:ͣU�Q���i��j�����j-:"�C�l�UAb2լh���j1����Z�`ţ155�(�gm����ض��`�ɝQF�j��N)&��Qi�4b�&�
�F͊$���b�cDL���AT�53b�:u�9"*���*���آ���Fɚ"�����֪��QV�U[Ѧ(��94ffb-�m�"�f�� +m��6�S��
��͌Q�F6ccEQ���
)6�4SF���kTQ�V�b4X�
JKa�QkDUP�P�T�DU���� ��U��ִ[LRPlRD�R�#���'o�;.�S/z�dՉ2TkM��L���ɳWTώ]-�N��_2��K_f
K	�`i1E���p����M��FJ�+�~ǄVo'N]!>���])V���Y���g2Z��'ll"��mI+���1WgQ;���N��|�g�(KZ\�E�:U�ђig��>sn�	5�e�S����\���	��B>��]#�0�2��q�OQ�(C�%Q��m�2��D�̾�ϯ��'G��Wy].ko.�A�u�\�q�wL	y܊�|e��)�Y:^�hÕ�o7������Y��i�<Cֲ|ׅ�Yञ��ܶ�o�H=YC��	�š=v�~�i������=��($�t��ۄY_���b�}�=�́�nd3s�q@IS��-ƵD���I��|����{����o�p<��&Z�k��[N�+���UcJ����#YL�F���g�]��A��gr�r����|�E��8쒻<� Im�`�HJ��m��"N�ٙNfxt��GSv���8v�����8�>ȼ�$���@Y�P|��V(@Bf\��ZV�e�N�(K�0�z�{b�ssj��dM��Uv�~^���>��P����8r�{���C�5sJ�
��&���Zi���דl��ʑ��(n6B�c#77�*32�Ӄ��ah��˛�*S�n�4��]�Y>����)�2��U�;v�vj�B&H����É.s�2�k��FE���v%��|���u!ܙ�k�QE�qC�P�'�bߐ[D��X�b{����ݍ���Z�]��AF���?�����;��<�ϯ�Xa�{�r�_<��<�`�l2,	f��wkU�ԋ
���	�c�,�{;�� ���ƅb�\��(Y��y�+��O胵DH�.�5��J.�\>��j�N9�Ϥ����Tju4����4�u�þs8�j5���L�zk�g����*��(^:�����Lec�ED���"bumo��+�Ρ����%fi�|��������ó=�j���<�"+�j�g�跬�ED�
G��۰�_ݼnE�'Qk0�l{��_�c82�%$ʔ\n�\q�2쳏Ƒ���H���E�3`��u��{~��� W�׏��~�����{�!o��3�(��JG�f]Á��b��^^����%q�I}|��9�nz�z��Ŧ ��JƸ,+r�ܯq�o��!����	֍�J��G�K|qoq���G�v˳����q^<`�(��+��W�����*֯m��G9�J�Ժ�L���9��C���C�OFe������bv�6����G��q��	Z9n����Մ���N�Tt�V�a�U<Y�F/*u'(M`:�/w�	
;Y�}n��*q��>^����������/���X�0�=�I$��*5��vu��KD�ލ߂}�oq�u�gU,��!��ڰ9�"�o^=����'���,M������z��6��:�
�p�ݖڪ6=U�)+�y�Q�
_l�	Zkb���k��4���8|u��&Ͱ��Νb����X�W�1�q�UC�d{��`�z�Qc��F��vs6d����]_{�;�&�j�5���[L?��=),����J~`/��wH��H�5�ښ̅�1�V=6r>�z�DfƵ�h;�U%�S婎��s@N�n֏l���/U�a�v�#�!1t�FX~��f�e���}�k��X��=Cb�m���XI�ݙ��ǵZ+O���qܹ��V�#�����q���,K�*�]z"1���JV��Ƕ�`�Uq�ѽ֛�@�l�A/D���֙ϝ���+nqP�8I�ރ���̏nz��H�6������5�N��0�/�
+�q��y��%Kn���]2碼�U��%+ab#`5뙺y��{)Wbw�K��/�{���o)j��[1 +�ՠ���|��C6:�=�F��i�ٵ1�R������˷M��n�7�S�{lث ����'�kں:��dG��x�G�{z�*�.N�Qr��=xYeMٓ�kS���m��aC�#�&�L������p<��6��x]�Ѡ�z7��k}�w��j��&�cNIJ׆}%��&
���IP�H�,�\EX�g���窩\$�e��y���Z�;����%WܢG��������y�{@��t<@N���蛉���S��˱ؕXl��V��V��z ]u�.�=9֨D�m��_Q9��9�I3ez��6�����rǷ�"�m�k����{�P�V����;G����S���?�'�A+;��r�=�7�"|�:�-�i�Y>�nxӫ���]S�ؘ���>3yר��Bē}�vՙ������{i۷j�}���cC�gR��oݙ���@ǳMjG�7F�c�q�}��C5J���q4����/�`ͪ6*��͖��g)r�]T� 8|�λ����(�s�3����ᄜ���r�?��^��f�zו�8�j���R��&{l�U�.�ٵ�q��+ˁ�L5G>zjD������x�M��ƽ��fp���-�P������)=�{���H�b���X�k���� 3]+Q� ��Vwn�3W����G)�յ�^K�f^�n:�Z���S�.1��+/:�2P3��'^Ά��\�v�J�.�a837K�����2�pI,49��f�y��DN�;�G�h߮�,zg���r#'�M2�M���i@�^�t�o)���.o��At}G��%��J�M�|��q�&oKm�d���t���`��{meTˡI��O�k�ǧ/����*�KԑR�I#i��'��d�y3��N�[��Z+��.�S�W�͎���j�O8��}�&o�K�ϦK�0:vB��T8s�,�����q�zsx<ܵ�E�N83�����eI�%d��������ם63����;�R�w׭�Ln�,I��2���{��Սv��Kk�5�}ճ�L���^��Q��m��[П9�lk�6{��β��_Fgɼ-��P�]`w_E^���!��t-��~7�
⽊���d�7��`��,9�:W���;�~uG��T|�K~��z�WM���L5�V������4����}��,�ދڝx�}=�3�.�2���*`�Y[<jR���o�ڣ�x�`���bCQ�8�uk��N�Z��"u��ll��2.
��p���P���Iڢ�M�4ڮױ�W[�z�;#�c}L;����v5�S��W��ͥ=G~���=9&������yk7��	�el�(`�����N�o�#��T�]���'��E�{^3��%��;D�H����h�V��������U��5|���P_{\+\���k�pz9��.O;�3Gf�~�\���������v�@\l�;ų��XNtϋ��K��&���\��NVwZ�����2v{�c���oL���r_���=l�+�=�ֺ]�<��[o���~���YVn|��)��{��.Y��Y��ڸd�31��k�2}8�����9�}8��,�GG0�)�8�rTjw����Iר�y���̂wP���^<�/w,ȈѼ`��� �s;����Q��P���|�U��So�����}X&u���`�po��?S��=��>�:k�7�r��F#��U��/p	%��`��Z���
�`���z@;��\�����y��W ��so{��XD\	Ժ����O��BJ�mN����z] ;����̼�r}�R0����Ɩ]��ش�n��5�62�WP+F�q���h����*��k�Sz�yћ�sy�y��X���N��n�v���ȳ�U�EOr���zZ�W@��1������NҰO��)O��g�������~�%���'2��\�S�>��goE}-���;��m�h�_'y}&�FV�}��z�L�k�oI�o;�4<�<��ӝ�޺��a�cFz
��-�=F{����y�;�~��<�������������W�Z�{Of9����f����.w�l���vm��޸0V�nV?N,W��U�5%g=̇4���,?��9��vW�~5q�Ǉ{dZ����{�^/Sk��D����9;��9Yƙ�Oƅ���1��p�.U�
Wr��M8�A�y�w�|�������6��6��SW�Aɴ��)֏�"�_��9���7�U;K�<f�逸�ޜ}��Y��'�]M�����6�q��Y�4p�Ou�ؖ��O9���}	��"�6ʬ�f!��̘�1r�8�I�[λ!}���>z��z׫�vsh��K�w��ʁ;㜜�yЛך�O�)���h�A6�Z*��:['kRdq���̕:F槶�o��=}�o[{��N��Fo�I��<�{�f����1���C-Y
��t�u�;#�'k���)����@g��;J�Ӽ�z�zo\Ə;�#t��c�������my��(���X�y�C�_S�:�{��y���Ny{�๐<������r�޽��pn;��	A�x�As�A���ߟz?���1��2���gwn�N�On����{X.K�,:�+Y�zvȑ��X�	�z;ٚml�ekf'%\xe=�xI=�X��V��i�5����(���<���vN�m�F�݄�nG�S�~!�;�v��v�ղs�SK���&}NP��~�3t&��5�1`8���R+ָv���y8v���vY��-�y[����^���M���g?7��/�Fؓ����o�ջ�	�e�zy�|���Y����'�Q��^7CC���g�^خ���q9Q��?>qQ�B��{���xL�A���(��C���MA|�<	�&un�GC�Gt�]�o6����f���2t:S����V](�+�*�V�I{�c�4s+N�ٗ�@����S]�oeIs!�uDݱ"+���ڄď��{OW��^�p�B��ʧ�eK?�����L�'d�ޝ��U	��s���<��R�l�Q7�ϰІ�o��ы�S��%�2 �>�s���Z�-�=�s�S���+��N,Ed�ߕ�ﻔK�ӢeN��3z��m�z��{P�:sR{Ӟ����ܚ��N����ʍ���e���%��A��ٿ��=�i�&�/{�*W')�Of�=��?2�g��v�����%�E�M�{�7�q��r5<9�(^���?13����s���}r��Έ_o(떇:��c�?t;�.�w��=3�������yx&I��g]�.��7�'���l�Rw�۪�=�Dיh�~��'��;���&o��}Y��r���x�q�	{�q����
�o�]A\�y�x=+�ޝ��<2���eI�X�����ڪ�Ne{����V��6'����[2�����]f��<o�i v��왬}3;T��֜GG���wM=YW��d-vNG~�K�+�Vx��G]e\r����aLG��sy�.�'R&wEA�N��� 32k��5V��.�"/75�#���歊Y��^��T���}�����2ę��U=P��d���0񮎭?6d�=:���"9����؛^��w�g��/އJ!{&Oc��zq��<��p��`��+�q־U$�����!��,绻�	�GR5���&���}+��m?Q�w�U�Nu[/��[�����ۭ��R�`򧲸t~���ހ^��N������g��웷���_��yW����x��R�{��u���� �l� ��m��=��8K��l�Pxj��X�W���0�����[�_[t;1}�p�ծZr�5ƻ�>�j��Y�ٵxxb�W�;�Ef��ӵ�����ِw�e��Nt�ھ A,B���׾��_g?h�To��z�t�Wݎ�鐎~J
챙x�O'K�����N����9��6Wi����l~K]Ԯ�7+.����U��;���뤯���@E%�;�tƶ��W?�b�"!�=+
����"U�D��U{G����tG���[7�W�;2��/Wc��TCC��2`�|2�sy�x�}mЯ{i��rp'J56�fu$U��VXU2��EC�ws���� V�p�2����,K�6��du^;���j�6�
ۈlI#0i��WS����n����J�w�K8j뻆��N��:����rؖ�x�r�6�
wQ�_kb��x�n��t�{�F���ө�df�f�;
�!aΰMU����m�X�i�/�Y�i_Zڻ�����BG�1t�\efj��w
ݲJ5��\��-��;*��H�J�v�ҥ���N�r����(-4�w;��W[��iXz��6�v[u������\H��6��.�&A8Z5�w��4�\J΢S{�Jm؆i�6��֍Km��2fi�ɣ��I����ޔ`'���ޡ�&V��s
pq}X1gvϮ���;Â-|�x\�����.���`�'��|!n�o�V�u3�5��-
�I+7P.���7�B;����/EX�N�ȶa���K�ŌY��u�)�ۇ�V�V�AR�1�u*l���;\���I澭yeޥ$Wv5S,�
}�"���5pW����Cn�k�p�xHg�T�̈́
�{E���o���Vh8Kİ�'�3jn�I:�J���������oamҵt+�˜�Twe�B��d�A��h�C��B��ٛ���(��V�K���n��/�c/FVT�gy͠Q�d�e�����S��Q�%ԍ�	]ic�\鑗yN둾����=b�u�uC�E�����4a2�2��%�h�2�a��s�4��IV98��m�G�m��ע�h��X[�o�J����h-��皒��:̹6}a���r�S��f�P�&9�[֍�5:��Vnʅ�Y�w�=�H�\�,�����M.^ �f�h�q."�*�[@��۬e&([r۹٠\ʸ+�'����;O^(�]���7��w�#W)�a��|;�u���J��d��zĊ�*�j���ox�չو ���)z�|�Y�)Ja�t�gj�c�kC�
��
*��Q�8�Zf`hfZS{�#gB��ޗ9��Ը|�Ά*;(�,Wv`���'q���̧Z)b��9�*��R�U���1ƎX��DK+n���i+�㩚	����td4�ޏ��fH �����ٷ�˨�|Q�{ؘŊ��In�s��-���*�
8�jIg���Q�R��6�U]�'Ś'��t��c�w�u(L�j}���z�\:WLyq�ׯJ)Z�u�Xb�}�m����%v[.vn�Nk�����q	uW���pi�7���aF�35��[Vn�T{�'�"޻��G�jF�u���t�+I�d��*��kZ-f��F(�62Z���C����TE�kS�m���US[8)��chu��cm�5��"���1��E[b� �1j���mDEE0Ulj)�����j��4�jv+�DTA��g��Q�J"j*'F�H�f��bj4j*����hŊh�t8���j�(��J�"�5��+E��"�ъ��1F�AQEL�Th�E��)�m1N�F��(Ѥ����kZ��*6�ĕ[j
(��`�����m���"�'C����MUي"�""�IT�4:sLm�)���L��QV�%E4E����10STm�mj ����%��"6��b�"	��b�&�1Zm����AThqUC5UE4&�"������EAhƍ���LV�A�Q��$�Dm���64�D[(�h��S53Q�2kLU6�*����11Q4�Q�Z�:��l��	�I�ƌ|:��hW{�k�T�8�}p͔7��g��CÓ�������si��R�L=ɑ'��+��k�Tgo�l���/����ט�\�*:��ӑ2��M��C�{�1o���x�79=�;Ӷzc�a�%��cYΩ��zn=i:׺}���Cz�������f��a��r_VL�(��bak{��*{�;t�]�2kr��Fs^J�v/|M�zx�OyT�N��ku�L��W���W���7�cǣ��3;��Ks+)�]�|N����õ75�rM�u��k/��^�:�i�0�[VP�xb�C��lgvi1�����~�g�ӱ�q�ԫ�s:�Nlҝ�O�%��5�ݟo��xNۘ;�5��q�y�΃}J`�8�}oS�jlrrU~�o���%q{6�[��<���1Ͻ5�^N,I�?z뼽��������>>�O���_9Գ�i쿲�vm��޸2�%�/��{�:��΋�La�v�G�d������>��W'QJ�cY]�1غ�л�P��u�'��ܼ�:�Y]��4a>z=�Z��v��#��=r���-��C�f�X5�Ifr�:�g=�œN4��z��ݶ�l��7	�YzeTd�l���G�sd5r%Ш��#��l�	���C��;� ��=��P���\��7ɲͽ\��S��q���w�Ҟ��x��-��EI���}9���1�e�	��[�3���>��e5y6�ɠ/[m�ݼ��na�}E;���2x�_���L���q�Xv����H�'�w�Y��U�^�޸�`VԵ8��^�O&����zf�Ώ`�Y��(�ɹ�7k�|n>�a.��{���@g��;�T�;ϵ��g�aU��	��sϜxv���`�9hs�}N�x�z53�מ+�����<���P���2��w���;!oh.}a+���c^�� C66�{�ǟx'�y�ܵVz/s�%�g�他|�5�4�umd[^�Jʥ
8v�U�����57k˜�WOpHk�ēnX��5��]Ϫ{Pk����B�N*�]���B�=���
&-�h��ܺ�ufq��8�J��{�m�F�;,��T:yy43��?[��xCRV*���	O��nIG��TPe��>�;8ӝZ�7��K�b��>}�W-��+��V��E:�t�32���#���V?v�Nv7a4܏�Ň��wM�=���؟@d��r�)v��zg��z�3t&��5�1n��;�u�T�u������n{__-T{۞��7{�j;���OU��~���3c�z�4�Y�=���`��U��~{�[-�~��Io�u��Y]�e��Z���RFO�7GGlf��|$�=��z��n;���Ѓ����I���xJ�eoK�9y��f�G7i���aM��w)�>�ß�jc���]T���h��K3��{d9�k�������|͛�,9�݃ݷ�ܥ�BSnw��u/,�b��bѾ��.�l�9�':`jOM7���1yb��e�k�\Y�|x�k�_�lPw��l�2g4ǓeAv3'���o��������7�?�Y}(�ttx��c��;��6$��Fy������/�z#g��r#vY�;m�9G��b���"lD0�o^�J͹�NhJ�W���Vn_x��f�m�xLPe�5'��/��)K6�����]}wz<�8�v�w,ܘ�,�s9\���V��2\wˉ�fDGF̗��?UϤu+�D�~��w�7����;N�[Ŋ\��:���[���Kҗ���k�j�r��ztw��<�$�˝v��Cx�As� ����T�'�6��z7X
v�H}����&���7�\��.V���������}��.������6b��]v���e���>q��q��S�%xp�<{�X,��[gtfVF��5����z�݆�^��#��l~���u�%��S�����g;��:�n{�ot�b�ۗN��eó�P����/W���O��S����?��N�<���A�<�ti1�'���߯�A?H��Zn'���������y]/�R�}�P{/Q������/��<Ҿ�ϟ�]~�����s����~�|�̾�����C�?��=�*�p3:;����π�<~���?��h:��J���=��)���:��{��ϸ�����~��r�X���>?}��K�������uNߟ�K;���o�kޮ��#�g���?���?G�3��9��+��p/P}'~�}#�������z��{��d:��{{��~����	�Ľ��~��8��럿z�+������k������G�K������~��>����;�e�h��\/p}/�W�y��;=����W���|K�h���}/]a��!ԽK��<���~�B�s��Y�W�	Kɜ�%y{����oz�}�m
�ͣ���ܜ!�CX7V��n�ھ�e��%eS���8b��*du6�s��J��a�em4�#S&�	��p����w���:iɦ2T.t��h��P6ު^��� ^��L��c�#�?}��?�����G/N��y�?J�z������_`���^��_�O�����'���������������P��������3\~��說����W<s��y���������Q�/���}��M�8=����_����C�>Ύ}�}��?xS��'`���ԽS5���G�}��~���~����|H�y/����/�/�N�?�����'�rq��?��9�J������)#����F���cV��DhHf{=�*�ۑ�~">��G��_$�}����_��ox~���}��,��|O��}��98���	A��}��!�K�rq�%{ B3N������_\�º=���gﾻ���{�!���@}/����8SK���߸<���y��^�̾���>ϒ�}�	�{���]p����X@'���?~����o���<�׿��4��^��?������ל`�_oҝ���u/�����<�����^e�^���^��oǿp/�̼�~�4��&�u�c�:W������7�bo�� �~g�4�AI��C�>�<_!�?�ry������%��S��pH����3��H��}{/�<������V~O}d����W�໯��>���~��Py���x;�C��4��}���#������B�<��	��_����J�{���e�Gû�j��?�g�C��z����️� ~���^�����u//߸
W�?��Ѥx;ǲi|�/��`>���r�d}���{����/�{�R������,×����o�N�B̏ýμ�~�#��;���7���p}�AĿ�����O��^~��W�}�.���_.`4��Կc�O |�A�[��j+����L)l�*f�YV�V���A�Ѫ��\1Vؙ��k�;�&��p."Vf�U�������C����?2c��}�,�v�`�n�02� ��3����e��ه_�v&ةؓ̀]���L�u��nb��"+׋9�_ =[n�r����l������{�����WF���x>��#�~��`�=�%����Ͻ�MP�{��/��~�w쯷p��s��ģ�?`�9���bq���_z���>�|�O߳�Լ��=��w<���<��]O���
W_Ϟ���P�����>��i<�	C�=�����g�>߿�Y��W�w���N����#�}��}�?/��q��_�Q��'2�)���Q����N�{���}������rw��R�?�z��_cJs��R{/q���{�Nܔ�%��DՖ�%�������z�_e������/���#��gA�s�v�s'�?ǟ�;�e����_ �_��?�����=����W���8��e\��g5~�d���п�����^������_%�<���=Hru��K�/���G��y�N3�Q����I�����`�9<�����u;�����J�����7�������8<�aA��x>���=}�e�^�����G���p�_�����'�t����98ϲ�F��r{���?O�p~~^�ҷ���I{?ȁP�A@}�\&��|�<�w�>�����̏�y���ߤ|=��`>���z9��W��9�t�H`�4���<����?}�!�߫8O�{�啜��ޯ����ߟ��W�?����B��<h>���u�I��Ɵ=�4�}��e~��K�����.��}��G�����~~�]ː��kλ�=^���M/P�?q���|�N1�/�{<A�q+��=����{��}/�P}�SK����K��pw�����w�~�u�Լrm��X���zWo���~����G�?�.��O펤��'��w���$|�������B�y�O���S�x�:��~�����M��<uw/��ah�,c���P<<W��]�(�����-��eZ��+�ss�R��w6��ݒL���O�M�߬0x���[t��� ���dae�^zZ�;du�ļ��Ir*�<��9Lй ��u�
������+<��$���=��ǅ;x$�u]_��{~x�"�)_UWĕ"b/.|��R�'1׹'�_�}��ҽ����.���|�C�?���}��������s�����y����_��?}*�� �ᥟ�mC���;�ݹ����	��ￎ�����w{/�y��?p�G���������/g��i_`�=��P<w� ��]���bG��ÿ�|_}�?W�>�w��?Wsɥ���(���#���?J�{�c�_�>]����N�?}��s/p�_�~���^~瀡}���x]���:_#K�<������0חV=�F1���W�u��]6><���>�+�y����|������?J��}��/�w!��'�=AO?}�?Aܿ`�~���:t���;�YV��'ռ������/����_�o��_q��{���9?�>�q����~��:���e�NN���]:��x~��__pK�'�d���S���	�����ߚ�໭�߫&�67}߅����~z����?>�_�?�0�ܟ������}������u/�}��2G��'��q�.��׼?M+������G���6���jê�V�����;�{��2�z�i?K��<�?@r~�w�������������K�_�pu?K�Oa��!�?��O=�}�@>5ߠ��B��*G�q;����H(]���4ǿp���O�}���K�u�J�/����}��0?���4���}~��>��~���s/�{u��m{��_��W�}��x��?}����}��w����N}���)����>Δ��z��{�/G�p��/>s�r�K���/r��`|�����>��|�47�g*+/����[��8�>����9��)x������� ��rq��̯��{���:S��p{/��w\��@w'w�޸]/R���?}g�Q�k�uI�J����c��4��y[���2�!��2ڿ�������ق�t��p��e�;7�	�#�y���*�6���ȼ�����y/[f����'Ce�(N��/6k�֐��,�[Ko)%��-���=l�1�fGk���_�E{�u������DY��'�8��/ӣ��'�J����{/�R��\���h����'�sǼG2>��y���������K��?�u��?}�{	R,���el������׍�#��H|������)�q/��� ��9=����_�Bry�	��_cG�d}��<x����_���Oߐ���{�U�,�4ա���3��/_����_��</��\�����d�4��� ��!���<�n%{�����������Oa�t�!�|&��~����~����6?Y�~�{휥[��0��﹓�w����?w�/�r���J�>q�I�'���i}���a;��}�x�H����d�?�|��'��:A�g�3j߉��Ʊ�<�?�^�����o��yM�~��~��~��%��m#�w/���:��}��t�<��4��I��'p{/��W���Y��Cw�O���X�?�",�>����	�u���R�/�Pt����#��py{�y��߸��I�~9��|�e���H����.���y����埿)n���+���-}�D}�G�W�<��`�Ҿǿ�{/�e>���W�䟸���z���8>���=�}�����?����)���������~�*_��~Y����[:����|�(����{����}���r�d~�����J��uܿA����>��{+���������_��q ���o��<2��]�d�Gz���}�{���R?C��]����|�/����_���#�q�Y��_��O{�W��A��|>���N~���?G�C��w�c�����z^�~}�a��?>�%�������~��~���I�9ti�<�K�솇�{����O��S�θ�p���<���/0]s�>�f���]�?c�^��� ��z�
���9���k�|����/�e�y"f`I3�?[
�G���A�B1nvl�	9�/Q^�tNK�cI��	��hB^b��F'}��WL+e_ {c�؆h	�u���{��|��W�8��׆Ic?���������=���R�4����<��#�ϸ9��)O~�(=���s��	��_�į�~���Ҿ����rq��^o����?|g/�3�~��}/[ōt#�#�?�p�q̾���8�G�4�������޸>��)~���a�t���(z���z�W�y<��������?����C�^�����?e��E��������0s'�?�c����>��������+��8�>�����
G�9}��}���p���:��u/R������Z_���.�o?V��?�
4~�O�yq��{/1��O�z�'����8���h���>��+������=�?G�����}/��}��=��^د��^��^��7?,�\�Z�7o�?���_e��<K�C�?��S��_������8>��?m�/�����}��}��9x����W��rus�c���ߴ�g��G�����_��x�_e�?���+տ���9��h��y8�����d|�G0{+��_����C�>΄k�?o�x�m���f��_ꯕ�����0�̯�^��~�H��|H�y/���/��ܜs��;��v�K����:�%�4i^��<����������ol������߼:罯�gﬄ~��"a�tr��
i~�����!~����O/e�^���W��y���#��C�%S��hi��_cw�=�r�߶����<~�� Y����Y�ﻹ>��>�����������4�I���.��^a���!��?��}��>ϒ��<&��?���t=�s��Gy�ι�u/񼗚�$�����?�%���9������O#�W˓���}���{�Ծ��X>�!�/����K̿���^��o�����2��^~�������p���{b�Ssbo�. ���ŨoS��Ɛ`u���Ά}�M���5�8P��U�b��Iޛ�B�V^{�3�tE݆C��y�����E���+�`]����08��֬q�;;����J��x�h���H�ќ�ٛ+0�j%��UU��|�]��=7�?�id�:
�w����'���>O<_!�?�ry�������~�����ԏ�?p�/r<��?_���R���+�B	eq���S��w�sܾ��|w��|�e����u�<����:_�K�<��|���������B�<��	��_����C����˿^.~�J�r������}��=�쏟]�{/0������^柿�?A�_��J����4�q�_#K��>�}/������/q��m|8�>�~�3���,�=���߻;�ϔ���'ǽ�}#��9>����J�����_a���p��z��O��O��^C�x?�~����.����M/��������߭�׽�e~����Z������:��θy����A��p�}2s�|}+�I��I����<��'>��P{/PS���	����/�}u]k����AO��=�~�~}��ם^wߣK�`>�/r<�G'�=��O����R���z<�;�e���}+�I�{��������}���߸z��{�'�ϸ��~�y��8?y�ϛ��������7m�����~���W�#�>��Ⱦi?]K�s�O�]G!�'2�)�����}/�}�������ٯ=�z��;�AJ��޸>��қ��{����߸��������w�w'2�O����;���{�W�yN�p��r����������?G?�s'�?ϟ�;�e�����9��/�����Kyw�~��n<
=��d�3��{���2�~�����\R}/wp���y/�������C��=Z_�}�C��w��<�ez�������~�O�}���������]sxj~���)�x���}�����wUx���]>A��}<������}/��u���/�p���!ԏW�����>Z^$��2�O��G'�W���������uh�0>�xiֲ�t/�f��ʳ�"a�^	�漴�Wihv�p(�U����%�7��*��{@���Oe����=**r�1kƬ𾾷��s8���{��p���Rb�]Ѻص�x�G&����n�g�ՙ���9�E�9Fv��m9�'Vy�W��	li�VU���h*���:�2�[��׻,_sB�f _wimÍ��`�� �9�'ehI�j�֗�� �
��9�5Q<�g /�B�L��94��#l%�&<j,V�l���+�y�<�"�K{��74�bsn��������L��U�5��Тx�W�&�7���a���ݐd&��bZ	�M��]����j��B�|ؖ��%��\7F�2��j.L�XU2����OӦ�SKs���V7P[d��2���u�#*��yI�+�+u����7��ff��*qV��-,b۝C_0���Z����U��--CL�z3�:H�i*{Ru���2�k�2^�%:hf�O+z��-L,H�+*KaE��|��;,G��fI�n�=#�����<���|�`n]�!�5��2�6n�AN��·�1t�W%�j�{/���R?�n�U�_ExK.z������f�ժFʉq�C`��GV*r���V3)G��v�,V�Sn� �1���,ѭu�{��u�O�fF�Q�4-�������n̤%�jӻ�������)�zO[/aU�������Ab�Q��ܩ9e$ �f�QP�im6�J�zwx��ז���_`(b�_t9�W�m6��os���@�F���L��aNoqNTp�9�1�7L�Gs�p�����ڛ�B4�%�ǘË:���q�x-s˳o�*�ܰM�^P�g^��/WQ��LY��`!N����#�^���/s/�VU�A8/)ٮby&�u!q��+�.����uk+1��r��0��o��� S}�	]q����k��ZKs�b'�\�̾�s!;�xMn��p:ċ8��(��Y��/-7!��v��)DGD�h�	+��P�3qYz�oa[��TX�(�wr"�PŐh�k\��cL�c"O�c�It5��P���p��kYn����g*`�#fT�؄�ݝ�˿�yEؖk�~��v��gU�e]WD�YM��U��tiД��降Xj��yt�U�u�$ts�W��;Fe�-��R�z)�>8�2�L\��� P�K@������D����з���y�U��V3�DoK�=�܈:N��L�;�Y9v�:E��b!��.�h1�".Ǝ���&��L�9��	 ���\�SX
�u2�Y\!�c�Ȑ������j��{���4��(=���9���n�Wl_J��-��-�[�.��Q8..�c@�1����o��*�ͺ:o����N��(�t��)B*��6�^���Uk̘
���8�sz��׬T�;�$fE]�*&	*�"��D�L�:�QE;����EPU4QT�E$UEU���
���"'cQMTUS1QT����q�%EAU2kQLElf��)h�b*J�`��H��L[[CF��T�TQPDU1QRAQ1EET4T�QUIR�C1D�T�SQ����I�(�$�� ��cl�F(��&*'gP�UIEMEDD�TU����֊�&CcE5U%�E$�Zͤ�ATQMM��DQZ�V��M4N���QF�15DѶbh�5TN,Q�m�"5�Jh��Z�h�*"m�I�Q5QDIQD�EV�Έ&*���*h)�Mj(��&�QQ0D�TDUDV�h( �
6uD�I$Q�Mh2T[h*��X"����$��&�1PF�� "����d@�|vZ�a��.�sl�\�%�ٕ���� 4�ԟJܗ!ʓ�L�u�a�ͶŇ�d���\�����U}�]�K΋���~~�*�����P���\&��~�<������O��v����u#���=��N�%����_��˥�C�0w����?S��`����ܯ{[~٧�����y���8�J�����pP��ƃ�}�!ϝp:Oe�4��@}{���_�����~��|>��^�!ɕ���>���gU�ț��_�:z6u����s)���4����q���}�C�q�O?�>��_.O?�Oe�4�'^�4�K����4�A����G�W� 4���?|B��5Wvə�}V/�I}�q����a�<�ҽ���.��O�$��'����G'�G�}� �x������}�)��8��_���ߦ}������ܠ/�夓�r0!�y?v~�9��~�.�a��Cx�G�#���mS�⮌�FǏn�������jq.s�� ���9���$�ɝv>xd-�	��9׀����9պ���6Qu�y�����<�J�v|\��%�e�v%�AٱJ[�������Bx�ץ���c���2�xm���WOpHk��r��Y0��a+��鳪�f�|Ϭ��AQ����7a4܏�Ÿ���~;awnT�9���\�X�'hh�A=�/E�ǡ�׹�]��_K�(Ѹ[��]��n^
ݜݽv�J�/z����܂�2�+7�K;:)Z~�X�m^)�j�5d֎�4�;�;�)�-a#V�k,�.�U�[�ن��<�҇r\і�2j�Ke_]��,�V�O1���zt��S)���-����2����n����}oo[^��߇��Op���:�'e[�R�o��I~�o-��-�yY6^��%#z�ԛ��}/��m��~{�۪=<������h)'i�gBg7���ػ�'���o�č{ͼ^_k��a����X�Dv�i{}�5ygz	�|0W�A�V����7��v�[���۝�<V�-��C�~����Y������[��V�\�����yM^+�w0�Âe:�����N�Y#���a���l�9�Κ<]��Pl����(���|vk����Y�M��h��l�����{X�t/�����O�gL ����α,�Gh��Gc��ة�xy��q'd�<���1��2�oKϦof��Ӣ7����l��`��a���t�WNz)O��\���y���;���d�x.u�v]|��וUv�{�4_�����I��i�t�L�F��P���-ъ��,�8 SmWX͊��ԽҮ�tt�pv3�kn��<0�/o\��/��WZ�}��ºS�|�n�7�R�����̶�^���\&ru���At���M�2j����������r	Z�M��{���W����7"y��_t��%�d�v(Z�<LUbw�7}����y� ����0�;'�r3K���{�͏���{�Z�iA���Ŗ/�Z]LG>�M��v��mdY�<�ST�Iw:�^�`�g�����h��$�I�R�(p젞��TuǗBWH��665?8����=��n�F}_;��m��e�P���8U��J@�kv|�Ng�o��+�=W��Ot6�~�p���|��vd�t��~���=]���s�G����t��T�ۖ5��c7=����U��yz�[����ג���.!�wD>��ZrP��@�o�ދ��&��.��Պ�QƮM�~�7nf�X�-�a?%vb����O^;ߋ~��#��v��_s�G=��o��������O�z�|}���dU=�|lqiZk"�s����xȣ�)�$�$��{o��L6#<]ecB��ovXǺNJ�Y�l��kxu��JԼ�'L�Th��+�1�w;|U^�FN�>�}�W6�N��\;)�c�5�|u�uGg�C1J�*�$��V�m1K1���&��	�W�>���C��;�}�'��{��L�4Y��3�����gq�'�sMt�=�B�����!���8���}8��6���7+������<5��׷�\�fɾ^OS��I��e3�\���/�鶜�^���� y��/u��}{f�צ�
~����_Os�y9>ީޝ���2��~�a��ny��u���6~���|����<|�s=���3������
(yOUk����mG�S�/ׁǵB��޹��~V���܋�8���^y~���{$��=L����x�Nu_����ȹ<��_��;�y��;����L� 2��VM�.��pk=���}���+�E�ϯ2�b/���.�݄��ȭ�a��Fq����w�+���k��O��l���>σޞ��=97a3��1��=7~�p�If�z�m#K^c���R���;�s�it�w��[�1�{�~�Hx�Ln��Y�Vf��	�C.#f��|��l�aF�Ao3�	�.kAm1u���1�AWj�V���\���˼��md�Lv�
����k �r��4��?������<���̲���0Oϯ���6���C�}��j;+�>�S�}�\z��fI��q�z=���+�y-���z�N��v�^�ُ��Ƶ=�vd�)������$Gԛ��z^�^'�F��;D�3����\y�S8M��:�"�j����Z�/9����\�����ro��x$��kȘ�q�d����򔄳8_x�l=r�r��s{���jϚWqbVLى�����ɽ
�/g����l��Ts�q��9�h���~�fl��{R�r���n�<@ShT���ٿ�ĞɦSɴ��|}�V���On��r�B�坯�XòX	s��uw(�@k�{��UT�\��[<ޱm�{�w�L���;�wΈ[Ŋ���:���ՙw�6�g[U�r��E7���^\�+ ���?;!oO>Y��:9��wYE�����]Wy��^�JS�o8K۵�%ʹ����O�l�!nAR='�gR�T��y�|��#J'%jK�N��an�v�&����qVjJ:��i������ŕ`�^9��h��܈6��Ъ�f'��Ůk��ǘ�������e^��������l�o��l���U����	%�T�(7�w/%��z��~��k�6g�|�����2��kGo9��<Sܐׅ�&�Y��"�[�]:�η��Y+����e]4��Ot���M7#�)�уpӗ��}��k˶OTv�N��5f��]�L�����
����c�v���	�b|<Û"�(�Zr&j����߽���K97<�����d��wt^)�M�u��:�u�����l|�������<b���'�������3n�$t��-�o�]Ǡ�Kn��+rXn=������^���;n}檠2�;���1�vUϓ���͸2���8'/07�O#���]�v��˽�R*t�|����SƮ6�b�{\9Z��=�߳,�4��㙑�]�(��}���z��ƾ��.��~p-�J���ߡd�'�[����)��7ܩ�W;.-��F��D���y'�}D�r�N�����t�^Э�M��q����-�Fo��ު絳��4�اr;�hېn�$�;Lv��U�X=�^�ˮ�1�Se�(���j�;X�.�$����*	4�>�����(S�/f��7��t�	�=���������Wcg=g��v`��Rpd���v�+y;��Wx�ΰ�����v;K����+�<�k���Po=��N����M���3z^	�َ�,�D/��c,K��ŧ{���q
&O�)�3T�C��~~��&I��\�eׯIg���=�[��|Ď��v��&�~��s>|���[N��r;�k�a/Y|����z�{��Ө�=������Di\�i{j9J���^���b�rv����돝���I��X�앬��U�Ok}��~[���}y��9œ��㳻'g�S�~$��[�g��+EG���-���a�[�K���twX�:����;�=��9Lo���|���q��sF��<�N����ld�����i��}��kf}�4޸�Ň<��A���:KE�=N���;��3)�$��B;�+�}^�!��G&���r��a�5@��P��8gH�G��ҝ�3��s��Fw+6$3�"/�:���#�:�w�T{4,ȷ5Nm��s�=/�'�x&��C�H��I�o��X3rO�}��_W�W�~.[_�s�=�{}��}1vJuQ�j���Qz_�Cd;�obp^�m9�9�]��N;�~�-��Fd�ٴ�׶@��ܿV��e��]��Zdz��O%�%}9M����7��}y+YS�^��`3�{��bˑ>^�7�ծ=�s|�OX
�����KO�[�b���M��b�o��U	�_�rs����ئ�,b�c�ͮn�>��T��$��K�T�����.&Fo�Cs�7:T�o�v^�cѶ����̜g@�W��ز�{�I���cbK���ɨ͑=��dgɟ �)�:��OX�|T�>�|X��O�)�a����3�������90i�xI�{��7��6;��DE��`���hS�k����u@y\u�kgei�7w�8�������{����;�dk0�˟XA��.z^���a"�w��̡].�b(k�v����v��+��_;ǖ��[z2�����&�")��Y6\�Z�)-2���]�{������}ǫ�meG�.fا֦����/On��g c7����|1|䌇���s/9N�p=瓮`��^��� >�<e�{y�}���go��ܒ^��=L��V�ƾNu�j�i��o��H���j\�T��2���O��,	&ܺ������y����ü�R[1��-���
]���*]��i��������%uE9I�QI5�^����^�����=kf�My�k�c����o2��׌��3��|=Y�����O<�~tz[���_�?j;+�3��Y���oҍ���v�i�S������[���=|��ˇےS�����JH��<^iS���P:�R{L^�*�O�?z7�>GI���hCv� �K͇��ۇOt��XU�=]��9y�s�s������9�S��#�Y\���[nT��a⫋��|�.��\6�,'.g(��8����Ύ+���~���[޼l�n���;Ke�m���e��Θ\~��������|��7^��:4�n:R��h�񷂵s!�rU��R�Գ�F�����.����4+�g�R�;�ݍnu@7˕��s/efd�����grV	�bԵ��V�kT���]��V*+7��K���ydWw����F�c~p�FP�������[�  ����S�=������
������K]�R���7�����W��f2婈�l��=���"�uM3e�Ύ��� vBy������3�	�D��N%��N��دiSz�y��O;�0�:!o(r��W�S>�-��e��K��?�������L������߽����Xλx;!oI:{�Ӗ��&R�>^��t&B����<%O<�K�+7�%�T���a���v<�xܝ��{��C��u�_o�v;�n�y��<��{������s�m�7�>��	d���XSe]5�~����v܎n�u�^��)�!���u�[=g*nM��^�x��Tu����ݳ6,��=��\xc}�v�C\b�p?���Ժ���iQ�o�8�B\DB�n��K$x���ނ�����Ƹ�gd���fۿ=�s�o�P���E(��V�8 ����t�Fo0p�$=�qa��̺���^���,�Ĵk�*�ԭ������IK��/��M���\v��(�">[�ʻ��q�t�^f7�r�$0h)w�&B6?�ӛ��އ,uJ=N�%�;+Dm7S��9��Fֳ#�Y1��\��W��u�33�ރ��Q�d���e��Z/41yMT���ͣ�ս�=�j:�f*4o%-�ѭ�JAtkWA���1�X+�.�X/��N}w�Sʼ� ݱ�[�Ҕ!��$޿)����$[z����6�~�+�-�h�\���3M�9�����"��B�\T,�vI�.�:U�b�7/OQv�`G�1�Q�}e��H����6�	h\���'2��T�G��dqm�ԃ�v�*H��$l7Nt��7�4��2�Q�m��p\�:]��!o8�Ơ؋��(whW�bR޼�٩���t5س���X�h�퀟��v�m�7s��.�ݞ�D�j��yc�;qݱ�!�8�	�O�y��X6�+�ݧ��K�Z�Tx�X�J( �E	gU�Rr}&���˔v�Y�Ob:{,�Q����geb
��^��	̫�K������b�j<��w۷�4lΈ���)�*j��#�]VG�r5S���n�r��%�<)���]�;\�P�G�]0��}2�v�%�twF��U���¸\
#:�^�e��4���nM���)dZܱbf�
����2��SS����0�ru�l)�ۈ��{YeYb����G���4�:	;�e��v�)P�c����nX �^i�Z���w��x�^e=�!ׁ��{����}�m�Uq1������U�{5a�^��h��sw��,�2dN�+A\"�B�X$4j��#���kgXӁЧ(ga��W�������[��Ab�+1�r\'�l[�%c�yW�ӘbчT�47VV_K��b+�m�D"�.fT�C�*��M
�̓���t5m�����F�a�l���v�ӡB������P��Y@�N�3��Vҕ���g�GQ:��j@k2�&�L�˰�>�ni���)�(��F��!Ռ���>�d�w:uIj�巗��X�4�k����*�E�I��l{fno/���MK�� �/�����v��Y�E�m~A����H����9�w#�L����or"�)��(v��D�#\����9�}W/a�q+u�^���8)7�IN}.� a�vȣ���8X��ȊPP��(�!�,>8��q�ٛ')H��G֟^Y����N�)b�Q'���:ne 2��Y��n�Д����Mp�$jJ�΋`�C�eJ�Jes� (�>6��t%ʷ�6�PK��:�C޼G��Ò���_/��"Kޔ*�m�m���u����:�ǈ��܋wt:���;��`'�cn#��7�����d��Z��ډ*%U��;��)�J�U>���1�ѓ[\�W\�TEyfӍZ	�H�&X����
(��W�5h6ښ�
6��MEE1U:��"�*b���KDTq`���q8����iӢh(*6�TT���Q�T΍QDMTCZ5U�LV�:tS6�8Ʈ#qj�3���"�F���(���&*lقb��SUU13U3DLQ4�փQMT�;l���$�S1D�h1UUTSmE\cUDQ�F�d��jf*ֶ��q���&"�-�h�΍QE5["�����Q�����a�b�������b���"(��U1j(���l�Z�ETF�T�C��������n88�jiJ��&�
�""���Z3Fƚ��)`��(**�(��?���s�Ij�ga:�E��dk3�б�Se�7;{]M-�!�l�̠��ܮy�H�oZ�gy=��a�܏��O?�}U�W�X>�bL�)���{���������I�;Qz_�BU{ͼ^I�D)�Y�F���t~�s�i9�(�����vm���-�������s��X�E��n���U���n�=�����&�h>ݡ쥗�O�T��V)��=�w/�E�g[�ai���N/O�l��a��4�/T3����p��["�T��{�?KfߙEx6�A���W3G�mu2vxT�Y�s��{VX�ET�J��j�=���'y{����α,�GG��cC�oF�}�2�߽���or�S���Fl=���T��r���pǾ�Y2�]/�vSLY�����s�C]_T����>���s����e��e-�?g�S{�[Z���q�ꨀC|a��XC��볦�S9��wI���ߛ�s�+����ɦ�ç=^��}Sl!��=:�)����ü6_Ϝg���ta;^
�7�*3������JM
�Ցs����7{��ǊXǣj��uk�92�Uc�H�sv�����}�6�+8H^a�K��y] y75�=�7�K�3{/���_ݴo ��CsH%S�}X��P�*r:ul��Ύ�M�Q�R~����卿9(�t��o�v��r^�'���x�O}��g�����M��¬����W?S�\���A�'�M���+�a{��uIo+v@XR��G��{��>�w���홃�C�E`9l_���n3�I�a�&:���^9���f��;]:�}��'�v���4뀼�:gxϺ��vE�K���rnF&�v��rXy�jg��������[�p����2=��q��;���)�q��Z���S��߄>���m��l� �ɞ��(IfG��=Jg�����x�$v%5?y6�/m�f�J���5���9��}7<�w_���r�5ǹ��o��=+7Cxӿ��Z|B��=����n��F��'����0�=�{ݕ���gk���<Ոo�W����gY�\K:�D��7��!���������8��K|���5�����k��;�W���uY�vƎ���q��es;,-֭�2�}�;^�~ɝ(Rܡ��ĺ�61.�n���#�S.^쵖�5Ȧ�E������>���b�[��+T��8�b�s�5;h`Ȯ^nd�Z+��4⏃��@�t�+�yI(0mv��| ���fT�{]�ٿ�:+��	lQw��6��l�%��'<$��Tz�{�Ow�s���>���`îXC�_Wr�7��;��j��;��ɻܗzs���漼�ܳ<%�`�ϭ��]�����^�ͼzw�[�	Ĺ��t�đ�x\�Ղg]��Ӳ�a��p�k���[~�O�y��j������r�݀�{$�	S �;%k<D��{��=ڨ��ʽo�2��|'���u=�$�OpHk�I���+��D��:��Ɖ��y=S& �ܵ���M��?b]��Kr-r�p<2��x�n�~�oN�亗�stK�N���3/��}Sv ��p�<���ˉͭ�=��α�����NuYR��=-�|�K���微ZU{4랉I����>w�l��7W�ϥ�b��tnl���5��=e�ܷ�	�tUg���a�����n�����\�vŴ�,d٨���H����S���ps[EZd�J��ЛI�]��N��ݮ@�W򔣷�d+��˘�3��jj���^Ҏ��v�ᵤ�����&́�%5G_n�:�>;��BQ �J\�!3puV�o��� �enM:�����~���[��=������z7���&�m�T9�מ���̝��]ݦ��u0��l�k�ʿq�sޖlˡ���WQ7^�s�����lX����N\��?`q���,N^}���(�*V>�Cm�W�Aɠ,�9km�l��qE��Npn�d����Mv��m�Vtx�ຝ���J�M�I��_��̲�ii�� �ox��{��t�Ǧ{���_�'�����{<o�����R϶L�S̚�SJ��<���;��Z#x�����.�*��Ys7zK=S��S�u�G�^~�S�I�/&I��L�v�vG�/bc�{s7�u���|��nq�Ͻ������~�%�T����f>'���3��{���J�	Ϋ��л���q�W��zC�y��C=�{_f�GN��+G��w�ו�K��Jo��41�v�+^d��j�-g��w�5��5�F%f���:j�Oe8:��>��^Θi�	��]nԤ���Oa���H�nkS�����L9d�ԭ�X�a��Wk|!��Ί@UU}��r)�����w�~�����+Y��{*���/�x�7R���U���t{ZLZkɢ�k=Z��X����v;	t���{�ʎ�3����z�pg���\�������8���Ϩ;��m�G�]<��gs���9�N1�kw�G��u�T~W�'��������ð㢳̃�z��-���+���e��3�߯z�[sCp{b���1#^�~�5��W���cI|]y'���7ǝ�޻O��6��^�ޜ����W{0����ю�v��Ͼ��9D�M�}�B͔ߥk*z3�2߬����Ũ����|���#��=<l�wv�XS�am���{��^�ޥ5��qZ{��':cR{>�|v�����o�Cɿ ���8�l=鎧[�!O�f�&�=4�y6g��s�7��v����&���~���ՃF��m㈛�N��3�i�c�_<G6;��O+}R�Ä5m�|h,�a�o��3���ޞ�ͮ�o��<��:�X:�z(ИD���8�`Z6�\�b��u.��x�G�,��oN��TDQ�ڵ�̄�ʅ���������\�Ƣ5d�٪0֞��������Ͻ��u�{��%�WT���/q�M2	���f�`p��,�{�淮��ޓ��w���O�l����ד~y�z1�o�.v�{���3v��2{���ޢ�v������Ϩu��k�ϭ���u��s������3}W٦$�-��*{�s^w��m���"��5�˧U��}����w%��}Υ��ٛ:�p��d��I�%;$�5��z���|��8����{Hf{�Iu/�[�O�j�t����J��L�@��neه�#-}رs�Y���N��z�8�Y;��׊��*��;�����V6T![��r�Z�{ЌѿSe:��R��%���-�Z�:$a��t��ޙ��R�vV�9�aM����y�K|%b�^̤���"���}pzs�\�8E2��=�ǫ,�C3ב3�gm�G�q���0��{���6���{�#=wu�H=��U�]z}���F�ȼ��_���e^��RG�_a�)��W�������ѩ<e���T�3*�NԱ-�F��_��l�}�_=^w��nՅCċ~��hnJ�3F�)���gVo��]`f���~�*\�p�H��s8�J�m�cr�]��^0��9>�Gҳ4��W3�/����ﾯ��s}�����k��F6��^�/���I����Z�H՗�]`�cU�D�N�B��{���v���^2���"k>��fS��ǌ/ǯ��+-��X��	��%����'DTma��/���VV{�)��z�Mg��qX�;!.T��=�v8�t�x��?0��՜7˱v�pߒ��eUB���넛i
�&Ҋ�S��\�i��։���}wWC:��r�q��tD�+84*�d��5<���/܉����Ԍ����w��;�Z2s�yvL{�rf��,�Di���6��2�qvS�˩Sˀ���G9�T�;m��N�$O���Z��5=&x焠�X�H˗h�� �5�B�K�䙯N)\�s*1����)�V��x:��[q��nJ�V筜��&�h��H�@�/�����}Oӥ�s���R�s��`^�r�s?J���2���%LZ%�>=<*�i���jb�����~�*>��{��u0m];X���Qj�ˋ*+���cN	)Z��,N"+x7jj�Z�8���2K�9�rj��G��3s�V�BL�KFTnJӭ���n���h&���������]{
�D�x���{�T�!"���X��z�v;�[J�X�`�O��_�!'/9[[�J5��V�5�A����
ݲ��l�M��'�����k8�����|wK��3� �\EX�f�Y�'�5ً�i+�[����g�`��s���쟞 ?�iyK��޵g�V�����\�u�E.��8��vZ)�d5�n%������7��%N������V���u��]�J��/:���
D���������}ڎ!3en-��z����E��Գ��75ׅ�ԯ���b��f5sٽh�l�)�N�Z���մ|:�h7���y-��2��l+7�NQ��,�ͷ��+_J�x���2�D^�U���{\D�m�|)����z���/�����4�o��5��|��f6G��]D�i��ZU��Mv��=�a&��39x'�K�����g�mm���Ր�.b���
�K��6�DV��]��H��MH�	��[{��4��9Ӛ�w��X0j��� �ֵ�*�MѤ,Dr�ԓ�zMP1���YC��E��R�ۙ�*os�`t{'ӱs�4ѿ�m����S�}2��]���f�A�:+̑[����VS�x��-^�c�wU�������L9K����Ufw76ޞW�3O�
�d�7IR�6�v7�V���eY�{p⚟�����#�g#S=Ρ���3u�q��/�7d�=���38����D<�on;����*���s�_UUU{o���=����|�����b"�o`��*w�<�re#�QD�Ý(�֩��$t�ߟ��fyk룄�0����_c���^i�S�X��{���`�Y��~���)��w^^��M���4��+Z\YAB+����A���p�^2����,��!GT�^�#��S�]:���.�o�Z�<6��IW:E�t�x.���	v;�N�������;'��Z5�ק�1\v}��U�5z�B,K#�I�Y��Mq��]�C�Y��.��tPn��t�mrE�3ӫ۳q ��`2��s�=G�O�Tk���yK�H�3��Ho�+/������w�ec\�T:�3t���<��`��.���h�f�7��Q�g�na
^�c���=��M��}��A�3�q҇���a[ّ,��&udx���p�*5�w�*�ܞ�]=̎;a���E�P�z���������T^�yb�lZv��0�:�M�F�^#�]�Äן�~�i��`���И_)���uO_E��D�v�Wx��<���GY)
�{�V���n=�M�]G���%�%�,���z��V-��V!��Ҝ�+f�����-�&�ͨ�h����t��u|1A��)h蓺�up����j�]d8��g����W�vkB�q��g
v�'��1��lƀ�uoI3�}UU�B�)Ć�(5X��=х���5���@o�:Ey2<��;eB��}�Ĉ�E�<�cӯ_=����Jo0��?!��s��mC��h��f�,����C����z��(�}�z�G�oNҀ>5Kř�R��>�άJ����t����*��ʘ���c/�YQ�۴����!�'���*����S};�dڇ�k4���*�ʯHF�-ss�n�OBɜ�s4[��Zp�P:7��%��4�k��l�hy���u(�{�L^����ʞ|WM�O5�y�㢧޻@�X�\\YA3/َ�<CC�[�B��s���e�L�R���{�z�S�du("$J�_j�W�u2�L��iK���qԼ=���h���G'����<��<|2L�7燐bÀ�N�/���x�ϕMn��r͢�G�F+�/^��|q� ���2�."E^G��p�	�L6l��K�Eꗼ��<�;{��wD׳T��n4gH=�jN�2Jȃ��]�pC�0퉗f~4���Edf���<������L��l���f#N;�t1����挨g)�s8U�o4�Froul��i�Y�Z%�p��7�f��6�ګ1�
��;f=y���Q�]b���V"�<Xelx(*d�E� 9`ui�/.L�tቁIC^MP�8Ɗ8��jûK5��%�����&�#t./�I�*�f�++r��"�ݔŧ�Y�+㍶�QB�o�{��U�}+MQe�d�y��e���� ��E�5�e���3���oTHu�k��Ov:;��
�+r�X�L�ZBu�?�ڒ�]
��ue
ٓ�@���	��Ng ե�vܳ}�"!t�����iL,u�ݚ6�>Y��sf���ע��`<��[W@ܽ�_��)��
��>�� ���]�|��ʮ�&�g�'�`B/�E֜�:�sw_];㇖nmvXQ`�Z�%��ʉ��3�Y��Ӗ���j9�*�K�z��mŹE,�N�gi����97/��HS,N��NUbW;�+a�r�X�}�$�d��Uq��YG5+� ��R]ϛg��<�H�;KF�z��r�q�y,���S2����x�˂$�]FY
�b����b����}�{��Q�wQn
*>�Ɖ� ~j�ۮ��س�%����f}fVcL�էG7�49�L�c���]����/T�)we;�z�85���f�0�E�=���zeY��cyvzәt�-���X�K��xd���%ۧ&�;v=�;jF��61��9��7RP�6}�^Z�u6�/:y���9Q�q�SGS��EY��:�9�9�Nu*c!�(����r�r�L��c��|����*=LWs�7��Ř���r����)�z�]��C�{��@_G����.S6fGF���+*P�.렛�pJ�����+������s��C�ӈ��ZW�!��ÂyKd��xNg�Q�o�<��V6�Fg:�0u]�Ų���ޅ��tl%�d��QX�-�ce<j�hJ���`>�b ڱd<��]ҡ6�rwEG�wEbq]���s3km�=:�1���a�q[�K�N9E`CN���H��-oV��_e�����W�{|Q���w!�w-��Ks�>�f�7���t���r�81/��9=.�J�k�!�}O�q���Z���ݢT+���ի3Y�N�CaV���yRq	fP��u�����IW=ڶ�EY@�\�K�G�]�f�I�8�m���`-`��zy�ڎ�4�EPS��r�辜�{ 1t���:�-:6ff���VF�WeJyj�7�d��P�V<�y��fq�LU���W[�"��o�Y�+HմmK*��8�Y�8O�7����:y4ibgKR�C2Y]�S��B٠C��qph� �ԶCw3��:��X ֹ����#�	r�k۴���k�;i��n�Zzv��9��Ĺ���%-�SXU��z��γ��i��?~����ce�qD5E<N����$-��3ABAm���(��*i"`���*��(���$�)�"�X�(�F��3IADU5ARM5E5�5kUU1UED�LTm��&&��IT%USMD�1D�DDAM1S�:��"��-�U-��h�*&�J6�4DD�uE51G�513Ln8�"�j$�������EQ1UKGPf���*�b�
d�����:-bb8��P�4�%TQUPTAEqe���"%��SM4I�ESE$LAT�QQUq:�X����
h��8��T�RQe�&������b�� �"��ۮ����NI��Ĳ��\��6sy�'3�&���j����w#E-
�1�������G�(��ive�:�� �}�{��?Hz�oŤx��>�P��ma~��{���%�B�|r�Z�{��.'����ڔ���7~�p�Q#��u�:=�L�z��pwK䳜��6V�uh3)AY��f�����ҝ(��ڇ@~��0:�-J�d+��;���.>0L�3��ѝQ��2c�2H��V�]�gX����
2̟/:��z]i�g��1r���f�u��w�
���'�{#5���؆	��my՗�%:x}��@�f���y�#�N��a�^�3)�����Gp��c�����.�����\�)z��Y*��__
��\�n�q]9p�]-�x�Cϫv�ԝv��f���纏s��j�Iz �R�0Ui�����,���'��l�{J+NBar���6Qx1y����]q�`�\�|)�Z���U ��f��/)W���x��H���jFou�vf�_=��i��9+�=�����`~bc*	Q�!���8���r5�뫰�4}�Ͳ�I]gq��Lӧ^�M�ɂIμJ�	��h����U������NΤ��B���l�u�R�C�O�;]��sM^L�zwv<��
��o����Hӑ�<����ՈUJ�A�9p�Y�̊�Y!���a����K��j9c?}�������'�\�uߣ��q�k�~�<r �p)� E!�@%��
:v
u�N=�ctr����E��:{=[�רf�X�,7�<&K�g����'��lL4OI({͊tc�E7Y�=�&�>��C�<�C��\fG0k�y�?B�g�Tž�p��<*����o=Ρf����e��g��e.I/�X�����_�Yk1qf.X|�s�)Z��P�]I�{<����5T7��IWJE�eJ�)!*9��Ň>��W�qB��=y��YDed{�f�7����ܥ�<�;֋���/*�>�\H�ګ�6=�M���0���n�׎�����v�+f9�_�S$��D��yV'e,A�+L��X���
篆�V����0e��9�7��W�Z���5�c�r/�gK��ݺ�-��f�)v�yc}<��=�RT[��O���sۘ!�]j{c�cP��{-��M�g�Pӧ�i��e,�x�P/3�� �^�k�U�����y*����q:�}Nfy8���߆�^ܺpk�u��9Y���V�#E�ײhw���hʖlL�̡W�ן�0��K�>��L��T/ٰ],����l�^g.οx�u��ne��o�������Tc&�׊����Y�'^R��d�`��A\�Hٷ��:ֵ(�тث�(�J�F�(�?�����3�/M���|`�>-x�倹���R#��I���NU�~���������y͜��_����}x�{e���W$}J%�p�`��4�G>zjD��|�ѥq�*[6��_$������K^f���PںZ��A����*0�z�C���[y��l"�k��0`�q�A;�=cH��}�ύNY2��T� �4��9n���:������J[���3��3ޝ��y���<�֮���t��4?0�>��f��I�Y����P��U�7��{A`�,��^k��P�����=P��0v&]�N�7����Y��`�R�iD�f5���צ�{��:mO	w��S/N|ǯHy��y�-�Z���Q�y4�b��������ѡΑiX�P��w_m�W�ੇs��%���a�ڕi��j߁�{�J|�P�X�,<���W|&;����T��G���2��s��s��O[�ax�h�~Ge}�i
�]u��e��i�AYZU-Y^��۩�&�m�Ӷrݣ��7+a���2�-kD�R�U͸�<��H5��B�ȫd�޿��n)!��Y��:R�e+��:�k�ˬ� 5{��4��x�%a|���k
XjJݵz�M)Z�mMT�S����4�Ҭt�E��gn�V�u��5K\f_Mg-�9h��W��U�4�Ik��u�C}�y��q�,%��!F�.&�৩dv�������Eu�z0��v���C�ر3�����Y>��q��1���`���\"b���x���S��C:�Kޝs=�Gm�������Ep�����w�x{*kc�'�X��Ǟ�idֳd~���wV�\6=���/V��T;�R�ު�,2��l�5[G �^��7���ꪳ���O;ݘGA�n0z9����1,^���\X�
cEY��2���]&�K�{o5n[�}�~����)���
s0��A�M�y:��
���a�QX��@�5^��s�1�U��k;�NM5Q`��T��O���ؠ���tQ��aP�`1hS1�������㈡dAZ(K�f%oiE2m��\ڇ��1�;&`�S-Z�䜮���7�Y�,��?���g�*�I
Ǎ�4����Q���hC���sr���5�߭��:�a��n������A3/�͇Z�l5*�[�b���U��U�B>/�e�M��Ȫ�Y��E�z.���ޮ8ga�P�=�_�]��uDP}Lf���q������Ox�k���Z��5ա8�^�U�ؙe���� T�Hňf��$�X�nl!�
��Fo5
9�M�7��=��!u������678y���ﯴuxS�	!�ݠkW%	��ߨS2��iK���
�^�n1!��Qjo�P�^����A"���$��s*��q��5�K�ۙkML��K�C=�5�o`�V�r�1�����~�V`�.�\|�����2��E{�i7Է�ڢ�A�1��R��7�.Ƶsz�^������� �e�8�tb��2���{/���]�ٵ,L�՚0��8A�O�Lv�����J�u��\4uf֙9:�(�����N6E���w���!�FQ��Ͻ�L�z�wK&��t&��帥u�gz�g:I�j�Fa�Խ��yXܨl<��gP��Z�VB��.D��m�F:�>w���>�����l�;jE���^�J�]}B{)��lT��r���I�w:'��R��>��f �V|^�h�!��u�%u�C`(v���i����e���s��â���$�w��!�L��٘)��������(Y�U�����:��b��p;�}C9b�X]5ǭ��e�T*9R���hc+��A��K�)����Z-�$�H��(c��)Vtݖ��:e�&F�;���5$Jf�s�2R�����M��w��-d��\K�,��/l*��=y�m�nI��-K��zcw{�Vb���O��Cp����R�8��r�=C��j�ߓ΂�<ˑe�Ϫ
~�U�ᇔ�&gWOJ[G$�}"mҊڜ�&{7ـ�7ԇ�O~�~�/�z������,7�r@�ļ�6�/)WR��wr$s��'�Uo����u�'�cz>����3�j˜kL���Dx�`l*����.��=^���͊(lrm�NƮ�Aշ���׭a�~�<s҃�be#A� E�0i-�>���W�Om�uչ��w����b�.�c[���NY2���%�0�'8v֑8L(rK{��W���~�|B�}�f���̎`��^jD+�@��-�p�uK�79d���s[�Y����ԢI}�a}C�g!~���a���]ҽ��5�����������}&�c���2�Uґ~J."�U���]������;�|-�x�ɉ�z�oɐm��J$x�������g~�u(K�낑K�Y�����ю? \�T���:���[��rʁ����E����K�
�of^G5^�{��݊:Kz�#��{n��{*�]|�������b_Mೠ��f�`�r�E����o��}�n�ٲkՕ�^JR�%Va�4�_�g[��#!�}��+��+��e�ܞ7���ߎr�>v��s	V�F���2ODN;T'�� �i�>�c<�5��@��G��0{[`�FekՇ���7/��(������]+��X�x����%\��jY�};y�ٵK ����͂��]�,�j��Qմ|:Y����ݶ{��c�<�+8�ͫ��;we���ޥ���k3�u+�P�U@_����s�q3%�����׋١�?`�����=�F�*!JɃ�1r�lc�k��R"��$�{L�̧�����w2��{ӷ�ʾ�^X�ˮj�8������>.�`������:��*�x�ְs�&s�Vc,�c������<����6��#5�`�P���j�l����e/e�G���<s%���^JAP��˞��t��]��S�	�-�E��=VLi��^���ů���Eϒ#�X��\�F�fgN�a�=���[ޯ9L�֏���j�X��g�n�-��g���ei4�i���W�uZ�>=:��9�LP���~Wpk��Kǀ��F ~�ۼ{�q��X�;�]�����)��&`�"];N�I���X�׆c�\��Oq�Cg�8���J�VL��Z-����U��W���ՙޙ�<,��Gez��X��f��1.����@�s�h���ЦkR��>5Nj�L�%(7�L��sM��H�(���cH�z���C�����Z𩗦�=g2]L�w�����7�u�S�(�S	��wH�H���B�.���	�����W�<$.������;��5Aחx˶{�P��o�*K%���B��k���q���zk,��)Z�v��?I�_3V=^�=�@K���h�pS�rWާTC7��&�߾U�#r�ި����'$���ZE��0%c�!F�.&�=K ���
������=Þ�r���;B��e���=e=���}��c�§JK��,'���g�:��o��]y�j6�$Y��u"�_��dY�Vq�U��e3~��C4g]�N�a�,z�����*�����>�J `W��
�%�	�Z�k��Һ�`�|�a|DgU����qb˘���}"�H�˭/#�^��{��Pu〃d�n�tB��V���{��hgzoN������fe9�s�����ܝp��օ�U�W��F٥j��~[d���*cjEc�zM1����P �Z�7�qo,�4)�yu��n�f�8�ޜ���_g�c,���\<*Vq�z�!��=���#;z�&|�.�2�Q%0�D �w���M��ֹ�[�n3�"�îX�ǳ�f�p��*��eq��5Xif'S�<�X�τ����tQ��Q8|�Nb��s|7˭v3Z}*��(22����ĵ�(��F���|��	���]%i���%���M�c���R��4�"���3�y�Q{w�V}�z)��u(��KV���M����ql(z'`��/j]m{o)m;�w�/����̼wf��؆uz�mv�D��+'�w�1}�x�{��)���!֭�C����rP�L���3/즔vʕYG7�z�n9}�w�Q`ګ;�o4�Y�r]鷕F`����!�5G����.�o����)��N��;��N�iq�6Zhdrƿ}+0pjE���^��/+сH ��x�N�w�uT��g�v�9������K˰�_ݽr/}:�Y:XG����.�Ϝ��C-Z��(t�.�rIaRSNMl��7����H�5�B�(;ux>���K�ިBr�,�1��I!=�7��q���]S/�8�FQ��Ͻ�L�z�g�V��z�y�]+�WM���P�6֍��]�KU�>��D#W~j��F9����Y�A@|z<�Է���x���czeޣ:�X�*�wJ�%�%n��&D{�̓�LH���ZU�����i�FK�o/�蓬��������H�+�f�R\�p��'V܉4?S;^������/�l-�R#��0�U.Rb�7�xmoz�vzK�O[��_���b�����6��$X����	+�u�	��G��Y��{iY���� �G�,��_��Nǁ��P��ϯ�l�__�ϓ�ώyǈ�YH�@l�_e��6��q��2C�����Y�N�W��Ề��6)���N��:���=�7��;��d.x��K��1��}⨸*���U	5��Cp���K�L;��t�Ë��*�"���̾ޝ��k��\׫�2���Z<}��Ė�G����m�;�������>�k���^`�����|ë�(=5�*Q6O�8�:R+GJ~l�U"F��r�K�Y��b���os��j=�zߧz���a�W��46��Ij\��)���ó�zh�YQN؂s�f|��Qz��u�y�ְ��L�ȃ��)� E!�מ\�9�{�q�寝yzP���[,���樽P��*�'<��d��{��g0OY0��Ea{��w{���Z��kg��x%��0�(��ۣ�0l�O�B�Ҵ`�R�v��p���=O�B�X�to*R���NA3�����Gk]NHl߱�ݖ�+�ym@��!�bb*�,�RL��ʷ���[}3�;#<� E��e	Ќs�oX�;Tt�r�Ww%�[�:���cPf�Fҙ�z*�`�x~C�-�ݥ�	�j�Aހ�����^�I��K,3Wb]I�[���,a�m��Io��4,B�����r�;ə�t_eӌz=7r:7a����^��eB�[��^��� b���]q���z�θ��OuKנIQcko�TDu.�,D� �9������[.�$�D�c�S,$z�S��nN���M�N,�oH�6�w4�d���Y4�;�ۧx�S��� N����P kk�1��\FV��X����h'A6E09 ���^d��0����7�ڽ�� ��f ��"n��ki}x;ZG!��sU���P��m�V%��y�,U����w��ь�0ֻ�77��������]K3�lvs=d�b�EM��%'��TqMqUӸ&i'���/{�ؠ�3�Vp�3,q�X��;����.��c��qŜ�t�+ɉ�b�\���h��0�r3jEw��#K���ݫq�]\�Ẳ�c���fL,�u�����[A��]!��2�ٜgsl+��zZy�9�:�H����x�[�iu��)����6\��j�O�����/�
0��Au�����k&�P&�]��rŷǤ{8t�'H�j�,C`V�n�p��nk�')���	;�%��b	}@]�]]�f�s��% �����G���\X�v���K����aGrsk��L:�8;���p���S$]n�TY���8��\tp3�]�W�2�w�\�X�zWU����u����2L��N�%|�(�����f�S�7-�Ė\0�McF���L��-���:���gL��S����f��Wst:�;|ԕ|&q�S)d��z���9�FR�[s�9l1Y�=�;]=�:�2�J���U�6�.��r�h��n�&��X;�>���Yad������.�)�滭��,���f�-�k��*}�d�����U��d��=r�7sN��Z����h	wį�2��{s��;�R��E�l"�e��t�nr�c�e����1�Z�۳���Jl�?v"8��e�Ѿʶnd.�N'{	���Y4���7_m����t�7r�3��f��*Զ�f�%r--�$wc"�|�5����X�W�ƞ�bVƸ���-ĹN�ǃy@r&���Dt�w��u�#�̹·mZ��bqVm�ҔY���u��Ej�-�N�t'i�ӣbƻ�n�9��H��i`�72��5[��ڼ�i�-��-��:n��vMQ�t�<��yd&eM\H+t1�H�8gS]���H�K��g�{�#<E�t�ɕ�{S�T��_�mTCM��PDQ2EAE5%W�b�Z�����"��(�`�H��ƚ��&(�m�LQ%QQMS�OMUP�AAQ\lPU2�35QUIqm���*&������mh�"h�j&*�h"h���(����`�60PU$AT���������������!�f*(��J
-lb���"(b*��37MMQLTA\N�i*��%�h����REAU(��$��5�k&j)*"*�������MTL1�EMF�ARL4�53Q��)"���"���gT����wfv��S-!�:v�cK4c�^p�k���jѤ̫�wx���o�Dru6���-����Ω�G��ǎj�移C�V@ ���Р��6�\c��*�P~2���*b�ឃ�DvkѨ�k��n
���6��5ΓJ�Wڗ�}�{��/Ϭ���0��0?d�3֎\�ʩ�o�>>���1�+^��>�P��IWDGY��E&��(O��<`+��0�T4T�K�Aiu) (�-L�W��#��R���>�E������q��]�n�v{v��v&�Ǖ�u;�>��5�wKE^����h�S$�J'��ʱ0q�ENu��O8��E#�~���S���/�{ld^��b�3����x�}�n ���ӵ���+NQc}�ҥ��-c���vg��32��YՏ��2.j추�S;��[�J�md��ʼ�[ה�q�J�F�JK<d�L�Y:�wǵ�A��:,�3�Wq ��v��~V��=
��s}m]���X�
͖��e.X���/x��^$�ׅ@��9�V{xM=�ܼv}]ׁ�5.j�A��>�v<��_i�9J%�&S��h�I!��uT���<��vN�!A�-2���Mm�F�%1����1j]�^\u+Rm�#���;�R���֪�L�uaPQ�EN�5ܰ���t� ���4k� ���J�-�O6V���m)P�͔8�\n̷;d��i�2��X�2t�����M��m�Q��<�6���rs*	���
�:��������{�gZ��������ܻ�����~b���،�=cH�k�p|j5�L�z��<|�n���jͽs��סx|F���v��u;d{3�,τ�<e���e��+��|�{.,n!�z྿|v����vP��A=ki���M^uZ�#���=��p�/D��/)�K���yٷ����OT6R�҉]S1����צ�{�tڞ�h��Ҭܛ�s=ѓ�ӷo�5�*bs�1`�(;��@s�ZW�:���z��L �|�꼚�[틼�����u�����G�ؒ��(Gt����odo	�!.�K�{�nK���A�~h3�"畛�L�P��V�8২�Ҿ�TC7�M���5�ᗘ�������MAI�*�A�6�.n����p�>��p'�;Ge��Ve9Ż�z��=���DA�����L�j��wޗ�>^�9���`��ofC-JY��5���5�tr�`���WR0W����{\�C��=xh��8}��Q8��޲@�u΢�����ti�SI�����޲ּ2�wQݜ���Q��S�7�I��4�Aqr�9��r�N��eµ�Lv	w��%���e#!�j�WCCbp�l���$hu��N�ir�_^���g ��E��L��wy�f8u�F���7�`�oyKBD�WS��^D��E�������Ã}[H<_g��R�/%�`�hܗ���LǶ������)əu��v+������Lw�6������+�qBv3���ՙ��{��z�Ƹ�p�S�e�2��8:P~Cw;�FN�ye#��*�;-��ڏ7ɻ��\�*�����[g����k+K2��s�%�zma����ͭ��c6������#oï��2��J��t����$�(�M�a���8��H��y��ӛ����6)���v�u&��+��U�#s��+!覯N���&3\GI�������><y���dw����ѡ�H�`�āf[�=�C��Y��t��[{�0�\�N%���=PK������l�GRߚ$:wh�W%	���̩+�-��W9�+�H��8 ��rUY����2+:nK�7�ٰlժ�
7�x�?�]�W���*sݵ���9�u���݉ΔU�B��7V��u9�f'�܉S�ӧ�{7��{؆��f�x��\7:I[}�=��}z��%#{���[��f.nd�)����եæ�l�.�j�̉���N��:�
-]���.�|���:�/��j�\n�������Uqw��ġ�)4�X��+0pjE���^�R��̲B�^t�P��&Sڞnu^��Ie-*����	�{z�^�E��,#�VD�2�
�G�)�����u�m'E����Q���c��8{C�eR</��?.7�>ͬ/���;���%B�	����.v�A6i�}u�g�tb�r��`L��:ѳ�Z��j�σ��K4Z>{�)AB��g��Z�m�wtPP�7��8M����/d����yT����dc������@}S����/���G�.>2��&��$��O[Ҽ$��t�^�Yl���3]�����=�)�{�7u�ݨY�R!����n<���N+>8ǈ�����N��e=	Y���]�q�9��+�@�?aWl��ْ�j�Ǖ���V��pr���f'R�e�!��]-��6{�"�H�lӾ��%)��`xk¨���Q(I��B��4;�E��q]9p���v�W9E��z�wb���wؠ<�:��Th^��M-4�|�������m�;��=4U��!S���wWy�R�H5� �Nǘn����rY��w{�ĭ�h��.���|suy�:�ṶzfZEJ3KiܵY32�Y��ӷR� ��g��]L*^�\�D႔�8\˩Eu^�ɫ�����-�˶L��Ɏr��v���m����W�)��[>w�Yj�������x9,9<�'S���NM���S
�<��|T��@�TyL��,�~��s҇5�'�K46��_%�p6ؤɘ�_�uϞ�ѽ�56��9.\��+n�N�_��k��������4*ًč�l��ž�_�}7b2���b[��P����~w5{�[p�ߥX�,	9��\����pl�w���y]�[=~q{Ӛ��Y�����$��a
����������ϟ��V\�o���ScX,{��O.�x�^�{��oe2�0�>�k/�Uf]w��;����t�Ɯr�����CL��D�Ģ�+Rఱ~>�yo�ݣ�[�޷�,�]����xe��H�7������|΀%��p���p-�s>W�O/]+�+�2-3�h��0�`:�\	�t�O��bgzאf�3)�oQ���/C���!���;��ZJ��Z�أP���p^�hÇ���d� j;+�Ӳ>$�t-�T��dU�~��_�c|�����t닎b��"Zy���\�r�zhS}�����]�������s�8R��Y0���X�S�dYɕ9���ٖ���fC@�3:*J����!"�(��탥�Y|Fٔ_�=ǹ�dǲ�~�l�!����<i��I\-��z�环�q�{ {]3I���g��Ipjማ�`��9i�ǽKTK�^��u,��pŎ��Փi�r�g���N��2��?|k�7��U�k�A�6l��k0߸�\�����{�m���Gq�}�k���{�`���N^���^a���(ϋ�Z)qh�>�/=w��Y�u���Y�QP
��8�pؐyl"�s�@Ԟ�3��'i��W�Z�A� M�׾�f��1�
����C����2.�Y�E͇~���HB1��ZT�x�Y��s5���4p��Z��2H�U�oCq3=�N�a��b�L��P��pBV�Ů�ސ/u�2���Gǥ	v�8T�\�#S�d�[]od"[�ʾ2�s"�ɤ�Q�1��8�˗c�h~4̀�5�:Q$�� Y�K��N�S�&�f{������24͖�����'j���G�Tł`���{�M�^�7�V���wQ�_��-euѰ���m�JzA�gR\�\ʶ�G`^��v�c���/����L�B���̝Z�
�Rg����:���c7n礍��؉w|�e�Sc�j)�6��F���7�9�KMp�y%��r�n�����Q��Ң�s�r�_�9��1�����	��KjcO�yp�|e�=��\�E�#�I�i"ǝ������_h�)�������&߹Y�t�]�0	Xax�h��OQ�B�*��$o%��^;���_;r�Q�ұ�����3��/���1�sr�X�5F-0l8)�]�+�8{,gcEvn=�s{wH��0j��z�Jk��tKTI�Rc�\߶���hOT�=1���O@�z��}��w�Y�s�y1�AA�T�W��qp���=�5�U�3Ժ�m� �����T���|,{;f4�M������ۇ7մ��~��\�z\|8fOm׃_���{k���<|�����>���f|$�#��dW|}=ͅ]�LuW��C�@o�`w[��M}6��	�nw�/s��#���]z�Y�pj�,��f}Nft����w;���r�E�f����m��hˋ}�I��'}�R��khD�`�2�8;M2�V�bu9B\��	�~==�-G�No=�o6���FE�GB���>ʤUi�1C��������>���eΨBQ2���-W�w�i���d�[�v�zܹQ�ʳ�����o��Uw���u���Ũ��*(bq��s*N5oLT>�q[�h��� )�*b����T.J��SM����Dh;�v�$BPr1�����ln2^#�p�9f��3�wG�3����W���W��R�hg�(h��RKG�TG_]�V�����e�Û������)��&/5�'��Y���֫]H�`�.$3~�v_��s��c�;�O��s���f��zz��b��;P�'��h<��.�_�J���-"�י�������J��z�s8����L�7�=o�C�A��,��Ѥt�����آ�}eZS�^�h.=��m(f�M�rƿJ���.�.>Ez�J�����nT^��/Ӣ޲Y��!v҅X��u��{x܊r-[�`F䬈1*���������ُ�� �=�X���2��|#�X����BZ��,놛���o�@ jtD���F1gM��{��
�d>��Z$�|w��o�u�g�@�,pb:���ww��D%OϺ_'����Zgϝ���A9C�p�|�G94ʙ��,��K�Eb�tk"^�{k�-�q���#������q�a)�BH�=oJ�������&i�C��m��v��Uc�G�K@^�wq�ج�8�8>��	�i�]Ǚ�o4�r��=J�u�%�����.ʋ�Z��bpi竔�)�ޕԛ��b�Q꽗�Dc��=�k�YX�3����yi��f�x�G�m��l����W�}�T�V؆��m_!��^�������N+>8�<Fo�{�~���֍<���I	:\��fzw��f�Ľ)CV�E�v�Ϲ�
�f'R�����t�a�!���U�L���=�ر+�+�	�JK�K�	u=J�n�Rj'_8�ku(u-�'f[�-u}�y�'���5����F��%I���ϒZ=�
�`^ M�����\=��U���]H֕�\����\���5Q����!aa��.'f���u;x��3��t��'����*[��S݌�P��M�e�N�9�k}8�r�0��ӉrL�(Ϲ����_��y�OOyb+R�L��\��[p�{�֍<��0_�~�b_�U̿DFff�?&9�)'�F���Z@l�Iy��4e��p;w5zV�:�J��\���>��<����5�~#Osk��(��x�ڽ�yw�}ґ'�/��⿷�l3��1.`��3y
��~�[~����:3*;>�iA�O߄�C�'�C,�pt�Һ�GR�jZ�G���nt��Ww0��`n�n^c�i�}����'��G>D�.1�e��g���`*߶U���M9+�V�Z���e�"�Y�%E8+K�K6�Ol�84S]�KW���G3bT��ۤ�v:�j+�oZ6��˼���b��<T�K������SR���x�歫v6.ƜR��K�	���2�Uґ~X*WWT�땥������\�X�3X�'Y�wKIYqB�˶���씼�<���L����#��������ʛ��d��۵��eg�L�-3�h����\@�@[�zb�m{���\��M�����7��].X���!���{^���t���\^�-ׁ����)�ȗw�/A����{b�}z_����υT>�=y��n`g�^�bb��D�Hfo��l9�sO����ɭ����J���-S ��Y���J�J�߻2~Վ��;�����'ZUMq6ŗ"��V7�D�� ��M��tZ�n��K\M�3�����͙���BI:�k��G}L�J���:�Ý?)�A���ͥ��<>wBX�<����gZ�{&�R�=~5�O��3
�#�=5"Y�ۄXNv	6�ߣ5�dʇ���!}v���[yu|���g�m>���K��T#�w�`�M+MC7�v#.zƘq=���ƣT>	��BƆ�ve��O�j���mGD7+�V�1�\cT"�h��;��Y��/�|oV�Ř���A�y�l��JG5R��K;�C�ڃ�(!�Nn�`�7�QO��i�\޽T�*α�g�Z�[���������3�^K˹q��W��B�Ҙ�d�]�ʓ+V�t�9;�����{rQ��K�]嫓�@$��v��������+)�3L�'j�Ӏkeފ��H�%�U0�M���*k�>���U���R�1v]�rX���|�8Vkȯu�ٶ�J/��һ��4\ `��>�T$��T��ʡ���鮘zEؠqQM�*�����ݛW��6��U%�W$����!Σ#��w�qp9��κZT�"F��Q[����Ք��*2*�5�d�K�8�V~�1�Ux�U�h9Pho��P^2����{��&��V�.�oj�D��ǻ\�M��N��kf����Pvc�n�u|�u�Y��\P�e�VV����6s�Xu���-��hÏc��lmЙC��<�|i>�|+������Pr9�r�$r��Ff+\Ի�3I�A� ޭ������d�JS˼4oeZ��ۣ���(.nt�d�
�K�ى�H�9kv�(;�z��Pi��[YJ��\���B
R������ۋUA�:�3�$��'�(�SmR��cVN�y��]�]W$B�v��֦�X��ZZ�����M��������FZ�X�(.� �ע�ݧCZ7��w23�Z��~�.�5��}yvH+^�:}��'uݓ�g��t�<�����1D��Ywz�ut�~�ms��)*���]��6��������E�8A��*; p������>$R���-�C�<��tnaq�*\cU��h�]�pm��✞���{+6�m.�+�u��Tv�����ˬ����x6��F�4�O�T
�ݡwu���%:N�'W��n��%}���vc|@*w� H�eU�E$�YcL���PShP��N��=��b�Q�}�}�y.Z�#[�r�D]�zl|�O(ʺ� ͍+t�l�d7��k�r=X��6ua�f/�n�>�fő�묲�Cce�qC.��v����9C�t���?T�wF�`�b����U��᧧2�*m2%��	���̌.�wr8^��X�Z����ƴV�:�;�s�����Q�zf�k�΀m�	�B���}��7V���>wi��;��ʆ��;Ap�KPR�[�*��卆;�t���}��em�p�n 0:Y4[�:r�m�t�/�W��9��@i��b�^+��\c�Xt�����l���Uv6��`�KtVm
ف�8�b��y��1+x��,�5716��F�;:���5�/Qc��j�5�f�lL�AH�yD��*#[�e��sx����+��ج�R����u��Gs�k��W��a��ïD�v�_��x���yRGz�U�o����>tyS�/�|	**) ��h��$����b���)�cDEk1LQU�I6�TM1EU1k4�STQLA0U�N٪b��S���$���bJB(�����������"��&��:X�*��ц�����J��*����h���cDؤ��h֒���8�I���`�Vت6�SDh�E�R&�LI�1T�`��N���i�"J4b*�����
)6�4RDD�AEhiĄZ�ε��4�3��Th��M���T�5��h
�|>��*��"����6���|/y5J�kK��H�1:�C�]j��̂��iJ��jL\3q��i������[��q)�RzgjN��E��#�����\D$�k�\����K*�����[d�	�l���L�u�q�Uy׸�<���`�J#�!��]H;s�U�=Y:�+��I�{w��NH�y^��q�k�=u�}we�)j�:�����`j2�H~�����޻����ɦw�Ut��u�.�t�Y��*bp�1`�(;yh)�r&.y:ONw�)��^�盥G��f���O�F��J����˶z!)x�P��X�-夾4v����{}������:�o�[��Y�T��ys���F`���U�K�?#�J�m׽�mW���L�&�ﺈӖJ1S��o@��}��7\Fg��V<�EG>2���7G��s�_Ǽ;S�֎ڰ���C\����p�3닃��K����º����%x�z�s��ND�u�d�gVG��͸p�]�:���0����w�xz���6kw����y��o��ܼD��cٍ,ml\��Ӂ���>�X�t����V�3�%G����]=+dP���]�u��:��$�C}u��s�8�zҭDWl�=�Z���v�k3e^2���R	(�h��6���`ے�$�:�+�dʴ:8����Go־�NQN��ɒ�ɶ�X�y�Ή�m��)K��la�nwo	�G'd��b��U�5�M����g�n2�����/j�{��gڵ+�]�S�ێ��kշ���xW����*�g��;�fe9�}����0z;�ػ�}m�<���53����W��j�Gi|�W�[f\;M2�V�bu9C�',x�a�ƛ?M��\��l{�Nލ-���\?,g�Z)��P��f%oiE	��<;=A���fw\��{�y��I1���_�*��zN"���I��W
��)";�v�X���)c��:/^�$�=o����8{��E<��!򷦇%�;����E�qqe�]~g5�S�׽��z�r��������C'��zz��b�:]"T�@��4��?��k̾��֝��Q�l��+��Hr]U0�Zy/O|�k��M̮��8u��s��7u�V�_&�D��+��L�P���ġ�&�M�X��fi��b��dW��fM޲��޼�?Ln������,�6�F�\V
N.��>W���^����ȭ������}}����D!Ot�苨�^��\CwŘ#c�Ā<�'����q?w;ʝ{o����/-.:[�R]�9@f֛��t�����͕��v%^.�pѸ"�-J�S�5[���4U��O�-N�4A
��i���-M��㵇{q�w/�Vՙ:�Z�
��P÷2�ß?F�dv$Y�5�<\����<`�^y~lRog�9��f�$�S!k��c�ZтKGM̻��/)ȑg�l�����߰��d9�;���f�z�A�(j�w�
��nX`�r�֥�.W���8�K�1w�Sr? hR?s�h�4_�؜|jw��>9����y�ˏ��5�%=�I�<v+�10��{%w�ё^��i�{f�[�=Η��G9\,q���CmH�'�~��M���l�^�/��d�.�A�f�]�5�z�ݹ��Z�J��Ϫ�g�,j��ȡ�n�<F���ݓ}����Et���#�Z<\�
�������z�|O��F���*U�8 ����r��_5^V�/�ݘ��OɀcP��ڳp��i�K�)%����v���;��-ݿ{�o��~eQ&v�/���P�A�\���3cZύ���u�^��.�q������jeQ��{�>���Z��y�x���	�5#8?N�9�(sXgںa���X,����~�}JK��Fh���~Ϣ5~���j�5(i%�3{2���ϗv�M.��61K���k<�ֱi	I%�Xy��ĝvE�a��%7r��g烵��V�׉�nu��}a����>�Gz=B������\�Y�6Twj^�^�n�l��ȸ��*K"(����&�����t�3���^�V�#ޝh��kPo�~�b_�s;�7�pj��猿{��#�z�(��%�L�w�֙�n�Jۇ^�V8�9�a�Z9O��Ck6�t\�_vֵ�ᾶs���0�5Α&����Pqo��|��S��y��9����m�|19�Zo�r������qK^���p���4�}ғJ��du/���oK|�7l��p˝:��O�@���d���2�i�%+^P��`�o�2�T:R/�E�TP���Uo���ֽ�����������V\P�2탟9D�rR�a��ZI�Y��ŧ羒t�4�ቨ+������+�S<|e�t�U�s	V�&��7O�vL�-����Z�>򦜛&e3�8T��D{��m�{´���Xxx���W����c��9-��׮��m����v�|O��
Un�xM�oZW�JK��Q��%wT�A�+V����K�2-^�dj��Q���y�ݢX�������>���.K�yx?��OPY޺�炊�~3�>��e�Ɨ��IJf,;F��>�wx����2$��x�D��5f#Wҍ�jA=���d����+{���]��i�3+!�1��܃��S�j[�.��{K(�Wh:����x�ӽQtѵ�P�wt���]j�.���g>1�v���`6�;=���V�y��h�V�m'.�$�;�t�Nǣlث
��k�V=\��'����w�^K�^�x����s��r���)����5{胉��cz�k��E4#-}��љ���X�
w�^W@vq"��M�E��`�.��f2��̨x��ʳ�_gb���J�wu�o��xІ�IإCeT���4�=5�֌�CŘ��W�Yu���7�Oo;'��j<�vûG��5���"9������x�ώ�37�v#
�'��w��̓ۧ����tp�R�pׇ�eˤx�D��J"H#���
���Bᱭ뮽����%jq.gy�~S��й�y�S"����L�@�:Q+�f5��g�oݱeuP��,�z��e�2ؼ��q��e�7�	嚽��!Gʘ�`���y�ZK��t�e����^����Ϯ���`�ޢv.3�yp�|e�=�	kAϮT"PBRޤ׳��,s�ߪwl�y�$�jW��_����r�����љ+/ 2��\	�g����5[�:�-���r�e�]Jp�4ӛq^��q2�$�����I��vֳzxǸ���bp�J�v�o��E�F]lZ���R�9��yHy�y�9{Z�t�DE׊#K)���gc����iU4�� ����+1�f�1��f��l�CeK�E�ȹv�o��N7F窽�u�C���H�[uR ��vz&֑lwL	X����o�4��s��c����ׁ�b����Go�f�7����8�K�;D�I�Rc�W.���NV����u��u��6,'��<�gV}�`d��LSz��B�/��.���@3Co�t�	I�g7�[���p�|#�#\1�_%<�֥����C�o�`���;�fS.�4���{��M��K�z�P�^�>v�{�[�c����_b�����+yd�]j:�UG�����@�{|���KH��y{����Y`���wڶ_��'������}3�f�D�pG��N�~�'��7����oi髋)m�Z�A�f\ �4�YZY��s�>UW�(�˩h��7���5��={��۷����p/JK��*E�)�}LĞ�[��^��Ӯ�g�T���|��wT8��N4=�&c%(�G���1%�Ѥ+f���>��w��Nt#}4�ӷlz��C���옄<չ��"ĳCmݭVR/���c�+��]��qUf��9��K3\�{F!��]�㮆���P!Ɓ��]�_�����p�,��7޾�wvj����\���P�B,ѽ��NBx�UB��M%.TGz�*<����e������iEY-l���x�5/$r2>��H�AfV�pn��9��js�=��?!��nmo�B��=׆����\Ж�"D�v���;j���h��s_U�}�xV���qw�Җ�l�8�����p5���d��o�z�-[F������gu�����!�P �ҢH���
g��q(pM�����J�V�\�pv�fY��q���/p���[`z>�Zѭ�@&Y0�$��qH����>W���S�j�;�N˯C؇����܎��^�<:��
�����fƑ���Rge�{L��+,���I��<����l�8&�	)!k��QkD�����p�KޢF�9+�i9�����F��V�#өھ�-���ҕ��e:�s	vB9���`��U/{�9r�����7��5�j�D�R[�<3��ttX��s	W�ۄ�a�[ҽo*ʴ��L�{Ottҏ]�~��O��v{i�𶸍�"�mY��}~3 N+>8���T����/1�5�T����:W��죧�Yx*�)C��Ga�`�r��4Ԇe	K/HѮ�]�2�8����[��Iɏ]^�q��-U.ڤ��z�z�E)'�S�f�����ݕ�"�0���u(�{����gUv���ܘF�J�L��&��LBt1N�X�2.^ڊJ�Ϧ�Wu�=�H��z�c_pӺ�⁑��{K%�i;�uf.3晚��Gp��Xp���VZ[Jh��R��
�a��a�cx�yT��? ���=�M�A�=��?�����[L?U��=),��$�Ԏ���~��`���M�S��]`�^$[+��R)�@�?-���a���*��O��<���xoUW�t��f�vx���ྻ1�H��8ОSR1���C�aϧ�X&.��}6^�Kp�Wvt�|E�����'��q��&uܹ��Jۄ{�u��խa�N�
��{����M�A���z�=���"O5C����;w5x	[p��ٴ�c\;ިcM�jz)�(���`��W�=l�}=d�L4Mt�5�q謩��������Bġ!�yb��{<�w��t�5��P�Y%L[s.3�	�����I2:��gk�o�WuWf�>ћ�S�k�x}'Y�1qg��r�pIJ׆	,NY��C-$�$^!J�N|��d�}Ϛ���]��"��Så���JIqqB�.�9�H�7%/+yv.�	c��x�S�ܙ����Dι0lr�%]I�V�9�<�.�Es��;RL�;5s)2�{Q�宨x=yW�jn���둭>���q*�S{;z\{�0���ŇY���3!�8d5fl��	ۈ�$��d}��
خx��R7�7&�Y��覓���f�s�c�9�Od�~�F��efT��y��r�1`�,���h�pS$�\�Z���ğ@2%&��٨�UE�8RT	��m�w�+h���Xx{Ρү]�Q�с�ъǽ�9"�^G�B=Zl{	��0*ժ��"��I^�~��jKn�+8�}����}!�86]��>3����N���e��zm��(yb�1r��ؙ�.�Z��9w����o��ߡb7���v�>��Cm��2{���< ]龶ª�� �� ��՘o� �;w��
��D��3'�����&��j4^�Ib���N^�� |*xDy{��:��M�6����k������)�,��]p�P�ӉzjD��.u��Rm3�3Z�ȅo������r����3������f�?rSԨl˸�i���g�N�e�X����&]���3��^ny�m擬�j[/�E�T-U��=
�Pd��z���m.;��ߗ`���d�>6�)ө$M�w�1>��hO�����2��bY�hs��Wm8������/
�z,��v��.� _M`��
�D6ds9ApwC1ɺ��v�=��<��=˵��V҉|*�+Sp�3�B�x/e�j���q�n5����;�Cr�i�dcEL�̧�B��Nû�؇�k8PՋ�pQ���է���jrL=ɉj�D6�G�u�@�'�A��Os����˗c�hƙt�9�:Q+����U2덛9=Y#s�1�4G���I��.�ֽ�L�,��ˆJ���S	�����7�9�{˜oa�(��=X�\�ݖ����Y;,Ƙ���l�BR�=��=t�"�FO�x�U�?buԎ�N�M+k��]���~��Ϩ���v�ϥa���U�Mm�3/ed��o�����=�~h��8��*�f��hK�]�巷r �:�'�H��0$P���v<�L����|�Ϗ�@nAOR�#�1�E�8?��k��E��v�.�����~6bۗ����-c���+���k�·� "bg�@��csn��ua��P�R�`�1!s{�N����z���>�L�^��{���H�pX��X&���x�M�͸po�iz/+��u=8�ܛ��w�WK.}�Fj�������:K�<��(?G3�nJ�:K���rC�v�� ���`kYK��
�u"�*��>��X/m����>�,=A����Nn>>�#+ٞ�k��5�;�ܺM��=3q
����rȥ^<]SH=|J�!zr�#��WP9��f�Zł�:*����)j07����4�R닅ۻ��)q��7���pA�������+P��kH�u�W���s.l����MgE��@4�;�J���e\쵙*݉g��u]:��� >��^<vP��&W/5��qζ���[�&��:�}���Ա�C�J�!y[�h블�Zv� OF����"������S�R��Ԣ�;3e�7cf (>�Y�´�{2�񈝛Ȍ�o��WC�R�7��+����1i�j�L����K	*�����"��=-��ݖ��IY��r+-��A˼�^�꽑0��q��ތ�xkRղn"��:@_b_*Zm[�8K5 l�{XϓV>a�6Ѽ��=�ʂ*@����e�j������iV�a�q��g3Ӌ�G�͐N�mt����&a���J.:�u����n���R^�����Hb�;R�&e�/�v3eu��ЖQ:/y̰ �34�/:�ϴ^�k;�2�Y��J��9l��G���r�ֈ��oiM�L�q+k�P_NC���Fʹ7Fٺר8����^���n�u*�,{ڷG�����8:M��(�ZS�t�����N�����F�2Y��F��@��;1�R�����J.�[�������
�əɎv(�qn�H�hu!�6U����n�oY��ۻ�\��J�-ڻ�/� U���`=�h쫏\����I���R�	U��������*�+K�é�v_Tr�H6����cm�D��ҷ%�������G2WK�ܿ��^X�[YHM`Ad���o���������e���ksyZ;C��MꆥI�;2�����	z0���g�^�;8%A��)$7n�ې�Wpmk��Hቡ����;n>�;/�m�=J�`���x�B`�Agk��*0�E�'�,V*y�܅j�0R���kv�_ kn��&���@�Ů�Θ/:�erl�J�b��H��P!�5�D	1V�2�ZY�ޢJ�S2/�YZ����M�݄�b�N�ʇkW������C��=�Lj���A��y 	Y���	jՌ3��<'�56����E-��gv��Q���I��/�$	�7���֖�t��y÷� �� -�ٛ�����'A5wÑ|ܶc��r,�fȖ��{��x>0�Ԋ�����r��y�
��7s*q�]j�ǄZ�1��w[��V[�Ɲ!0�EAb�+>��݄�p�؎�v�-����[���uQiI�2��J�¶eسҜ��J׺w�֯��e�T��>����C��强Lk]&�1�������FA��HJ�k�bc\ҊagQr�+X�.���|=���읏��iJR]+r�1>�2i��`&n�5��Jt��9���$�alK����6�U]��(�  �>h6�[f֧K1��X��j�-mZ�]�F�&#V(4�X��Z��X��b�T���X�SA�ӡևLA�Q�
B��-Q8-�Ai+E����N�Ӥ�hZMR�[E�-����(s�j�����m-i
1��Ei*��j�M��Z����*���N����1F�v�.�UA��%PfB�Z*�э�m���*��h-���l&�"�ck4�cTѶ������h�IlF��+lkfZf���իjM1��:�STm������IAm�,b��5M4�lm��iQ�����UlV$�T�bI�>"���J
��7N�=�hbٽx��=ln�oJH���f�.!�s�p�9�9,�{�Mm�L_p^�!7SS�*�t�냹@Tԡ�����s�t{-��֏������C�'C��`�ٗ�%�Պ���2�ɥg7͟@�kNv�=G�Չ��cm���FF����=),fe*Ba��Kv�v_c׶���G�yT��Ｉj��o��T8��}8��d�g����I���E�U�4-]1�0���M�;��k4EO���P��yt�QX�}��<�`�l2%7��!�Px.Wo�Ȟ��=���N!=\}�>���uFhwa��nmlP�s���&W5��Aڸ����{|'�U����Q��3�,KA���ϨS3Jh~�F��xw�s8�j5���w��<2�s����������#܁^񨕊\�`�L��޸�8&�M�X����>���7S�h#gB��̌����/�??�z08?� Q�GAh�����|�v��Z���]D/;��L}5gg	ݞЌ���!�U=]��0���lxN��T8V���j|�p�c:� �P���u^>�N�wK	.��	˶�(�� ���`L���yND�#�y{�>�(z��G9�,`�ut���R���븩� �m_s΢�f�]pȤ[��ֵ��㶈<�~�bu�{o:n�B1���(RR����m�{LfĢps��ͽx���v��bcU|fv:X���V�V�!Ҋ�9M=$��f��fgB�ɉ�n_z��zO�<a��P��i+\�,0o�+�h�����v�.���zT����:'�
P�*0�3�<�߳���z��=�I��D/�&���̝�����zr��#���~�P8ᦽ�!��^�x`�����8��ǫ�m
����v%�4F�G��ki }+�`��:p�VZ^����V2�"��7l�6(9N�x��G��>����Jv�x��/V}���+�a�Ƭ���ڨu+{Q�{�����}��B����\�|��s2�ޯ�:���(/	��=),�ݜ���o��;S���ޯ��d�P�}�E��索�r�.[��#65� �AتU[\0�s�j���q�t�HzΉɥ�99����D�N4'�Ԍ��;�ᇚ���'<��Z�%a�����z���K�
���L	o)�R�.��·r�Jۄ{ә�����S��%��g� �S��l�{���N��_�)�v�x�%�L�C�WRg@v�j���u��i+Źs7½�v)�hT��̷5�(����@���Lg��8��&��%5~jxFyO6��H�5{��ߜ���x�bn�ƁšH
�^��ͻ2�:Ő]┅�)�+��ӓCXYfly�;�]�6�/�K�Ρ'T82�g�;*�\`E�=��v���w^������%�+����d���0�5Α&�#��q{}��Sk4m:�;w�q�ۓL�4��O���%^j���E-z�Od8f��V*�J�a�����c�~��]3�YP�q���Z��qg��r��.ƜJV�$�5w�C-$��5��2���蔖ʋ����g�]f�S45Y�Så���JIqqBĪ`��e��x8��D3�j}1�J�I��V\D����/�����E.��8f,��a)�$j�Ǽ���̜{��=����j��zא�8V�L���[�4�����}����*X��(m��˚����{AG���^/R��ɥn�xJ��u�W�D�_�U��N�$�imh�'��M��+_�5شA{cܳ�>6�[K����,i�c��o�z���0�I�%�/Y�^��ʋ��o�k޶���;�}{\D+ltX)���'k�7��U�k�A�7��7�ނʸpV���a�F�A]P��Mvqo�$�LΧ/�r����鴾E�v��L��%���VߏH�&uk^���bMX���k>�����'��]-b�J�RwvQ��Aު�V��:�����;.�$6����0���Y�ڱƳ�-	�`2S��ƚv����:��������T�aò���e��k�X'T�)r�'>ۡ ���}R��L��H����6����3�Y/l¹���^���X�y[�v��\z
�\���І�u't�l����q�����3gZ0ez%�3��m<��)V��Q�>[��zq��2���6���K�v#���c���Iޏ.�ߓ�T���{���/'ϱlOs�g&V����L��h�f���҈�\a��Z~�'���X�<��C�K}��!ߦV��ǁ��]v�{���KU��:���J���&��̳��h��O�3a����p�^��^�\W��%LB��-L:a����)_��}}O� `����3/n���K�޲v,i��	yp�v�x	BZ�z�fN��}^������H�PBW��Ier^�\e໇��� ϟQyX7]�2VZI�^��{0�V�/���4�}�ș�T�pJ�ʢ!vJ��\)>Ks=�K����uĈgg��"EUרxS��T�z>��%�z�e��৩{���8h�_؇�d��^Uqp�� f=��݋�G�E��P�#x�c����t�=y�y��SX��v��W��5>h_&�B�=�O���l�ݚ�w�\�l���#%�
$�a�;�ksQvrett:�2��r�;�b�W#��[.�X�:��YxʥL(�(v�b��8LC��8tg&<#��0wK��(.���<�Ց�:osn��]��>�aͧqzK��l�����;*��q�u�(�u�k��?K��kb�����<cGa�U"��6qN*�O�Y�6��}��9~�2#]Xg	.���C&���ǳ���W����㩻~<�W��K թ\YK��L�*r+�VX8�8��fe9�}����o+^osշ����^.o���yﭜ:,�V3�V��:���ٗ�)��W�w��q�6ߊ����m��f׫�%�=�o���nގ�24:8��Xϥ"�E5ԫF_�H�9V�c-VO��k�IN�Mr�7��.uC�'/��q��ɘ�����i4l�Ȅ�y��~�n�.s{��ຢ6��e`E5NJ'��옼a�'��hm�v�B���H����o}%5�Z>��H/~�v^|��������,����==|ױz �m1I��&o���{ѵ�Hs�h��6�B�L�M)o����U�޹�q�q�F�m֤a�(Q�6�\>��I�Kh;��*�oM���F�_�G&rt����t���Ϯ�]C]�vOJ˰��ҷ���ؑ�^n����P0տ*ۭ�;f��%��^๚�6��-Ƶ��b6�T��q�.����n���;k&�F�݊@wx�i��4��7��o|%|Z�D��5�B���C�e��r���i��;��p;�;����x���"�G.\;�	�K6�F�������v+���ȯ�l�Xguߤ*�w�v;8�|�`FEq�˷����r���f�"k����������^Ty��\hy�J�g�a�N�wK	.T!_�f0p9E������e�8�K���2end�k^��Iæ˾w��{s�>���W�	�r�L�yA���1R���;[��x��/)9�o�J�E�fz�;���.>2��0�a��H�7n�Oa�Tdg�'	K�.�b0P�>{^�t�xR���*X�c�c�CmH��o^+��o�z�^�z8�>:�w�0>sɻcuF���e9�j��U�GX_��
[}C}}�g�-�T�ǝ���k�^�/)����/ɏGp���/��x���6��g�u~��c�kʸϹ�cp��`���X��N]ë��^1�u�,2=`U����i�q���^Y�;3�Iʡ���QA�I`�3'![�h�����>�Ō�=A4A�iE9ޝ���^�=k�>yv55+���+w%N�v��Q}QMiwW5�����w/�	N��M�u�[��x�B�w\�)�Yy}n;������[�L4{����6̩�,�����}�ɯ�2M�ޤ[+�QX�r>.[��z^҂�
�^f�D��Ç�Tc�ۅG�0�SϒN����N��w��hO,�H�Ӽ�yC�a�0߯'�|7{�ι�r��(zDi��&	;ߩW�N�9�sT^�Fw�u��z�N�W`s���0�(u��e�7��SE�2��T���4�
9���L�sQ���8��7{N�\�L��g?Y�GV8�9�a�Is��=l�}=d�b@�_o" �Gm�iWx��q���v#����/Y�xt�{S�����_��y�?B�`��-��!ÓCba�k�&�av\YQz�f�q�uz�et�\�7�s�-a��D�����rJV�2K�L
��;IL�Cv��M�{/^$�)��]P��Uj�觀�e�8;���/>2탎Q#������}\����w�v&�˱1��\l
yX�Z/��"�pz[�d�w����������ϸ��ѻ4�l_�0y���9�b`�^A��[�3�=���fyS��|k�IU�Raw����і�{���-��[��RN�kh�w�s�,d����m��V�M����nE-�7����%V��~F'�X��\��@J4[��Äv��VO��Y􏖔rܬC���C�G��^8Hw�Jܔ.9L�'d�4'�� J%�mg��� �#�E��,,�_z�b�x:Ҽ0��V�0�G�M�'<��#��wW�{S�Ǣ����ٰ>[-��n����:�hs����H���89��:�wv�6�ަn{�>�����躜��q4�:�upǶ��]u�<;:�T��I�	���~��KşWV�c%�@v���]m30S�����"'���0?]{S����ʕ5Dh���#n��@,���;%;8��:�)������,D�w�Q���>�~r�1�{����b�W��GRv)Pٗp7�ƚV��o��z����"�𔟡z-z��w���|j5�L�zĻG��5���#����֚���^Sϙ]wM]��mQ�{�����|����Z7�# @�#��rཬ�ItJ��y�F���Y�Dm	o:&��~O�z:'��]zׅG>�����W4hj��\�dg72z��y�s1F�p ,
�u�\�k�������Z�L�8[�����!Gʐ�ti�ގi���ߥ`/�}&�w��}l�y�6tn.���������G(�]��t����[1⒮@��z;���C_èe3�u{Y�2��0a�c�H#�<$ʆ�s��
ƻi���ͣ4�X땆�p�����-�e
�=��*��~k&z��C��m�]����LƲ^\,J�t#�K��a��}7ݱG�3S_V���4JX`�c�ng����R�G�;:����%�؏G����|v|v�"d	��!���m�4'ؽ�'�n�D7���E��'M�[�����=x�<�Qό���=K ���Vh�|�
�_���e
/e�3Z�N� �]�t�����h�<���-�o�H�=[B�̀���-���oj8F����^+�f3����v�AOQX/�\^�$���P�u�^�,{>{1��M����ʌq��/�)���S8�T����R�cҪ����%;x=�.���d{>{q�7|ǫ�u.3�����Ȼ�C�w������A�X�ܺ ����Y`�jq&�35we����F�	��&ߤ����|�*�=��XuM\Y�-�-:��m�P����[V��S�w�W��
�˰)��	�*�}��m�z:U(�����_%��V�t�ԭ�$����Ԍ�%r�^�h���5����1m���ھ�ܳ+R�#����3��s��>�w�ؠ	�=�p�lR�ݡ����8�����ofrD���Y���Z��>�@qr��ʌd�NC�ζ�Q��|)�qǢ�����r��&띱��(W�էR����>���ꇃ�|���C۟L�x�+��[I�;8+�2�}��>�����ؠU��"'�����j�өEsϲb���q�ȔP���US{�7{}JѴ�V��A31���? �S���lOs��x��*���}{׃�ߚ{�Z����p��=]v��M(��^
��ғ�]�����|H�f��A�I�Oش�s��s)�〇A� ���J���vP�{�Q({��Bu���ۑ���_�{v㩞�R`ۡ�����G.�D�(�7�t������ ���n0&����T˩��-�<G�˃�=�IY~2����0��uF��h�;_}{���c�<�o>x}���i���k���0$�P��f0p9E�R>:˸S�9��{���N]�:�*s��j�葆�8�C����ߗ��-%zభ�r�֤�$�NS��J)����{�}}�8}�˲�?�>U.&8/���<�|G|tX��� ����o��j%�0l�`aTH�Wm�)^�sB{2��~K�j��Բ��v!��ڷ3���*�}F��f��<r:��"^�9H�>�j��`�s("^	ܠ��G�u&Mի���R���h+;��î��օ�]���Z]�U�Je�NBKwY��k]X-ꭴڳ��Sy�d�W���yۨ҆p�(m�9�P+sf3�1 �����y�����m��kǃ	�a�,̺�tFb�pRٲ˸�^��z���"��x��Rq7vZ���U;0���Sܒ,7l�tuV<����J�>ѻ�SSZڐ@�wEfb�Q����b\�p_vX:�%�����k��]���p�t��W՛�VKĒ�{�M�u�թ��e�#Z�l�VԼ��2us.��G_[[̰�n[Nnh����4S��X0Jw��]�V"�P�RN��kIÊ˧�@p>d����óxZ�J�gR}� ���7�4(˂�ޥ&�d�K�Fc.3XҊ�!w�PfM��n��Vg+G+-�N����^��!Uq�P!�4#�����t�<	��#����tw;f�(_Y����x2�]:႖��wK^�̤�Rz1���]
��FM�����
zR�%̮����7K3�A,���xl���丞pEyOs���#�K��v�M���A����i�wWl�^-S^�����-Gm*͂��MWA�pœ�9����V� p�b�x�
��m��aK����:��gR�ͻ��9������,ܹ}�kr����5n$�t�%M�-Y&�A��8��9i�IW�Ƕ]�e5��ʺ�K��cL[(�ڭ��ݱV\�@��t���$�c�v��B��+I��妻�it�ͩ��E��ȏCN1.����V<��+�or�$x�	�|v3���)ɼ�xܭJ7�T\�A�q.�*m����n]7%C`�2��<�^���+e�b��]�͢Ʃp�ȷ)����ʵ�q�6yT���3\�sS������k�k#heu�ඝM���,�]VK6���*f�e��n��/�tt#�#��:Wr�;��43b�����u����]6�Χ}%��x��afM�z5r��C�\N�/�{�&9�X�������%�P���2ue�;j�)E�[N�@m-�7�4Ct3�C����t)1�����x�)��w�Y��0� �^h	-��7��@ʚ��P��K�N���4�u��ҕmI;��	�y���t����y�������v��>���h�y�'zoU�����+|�rR2fu>��]6R�Vr��1_]2��]����C:�p�i�I{�S���O*�� 	�;kt�����-�3qP���[�_7E���l�CVq[�\Ӆ�f+5��:�yX���D]��u�ʥj�����e䘣ެ1#�d���=��kC��5��1+���8�m�i60h�"
L@P��m��;f��ձlkU�[���)(�E�B��:5��ch�КP���-�)�4JB��:Š4�lUM&a�")�gX��AS��ѭ��q%-�U�6��+N#kE��ٶq�m��ggJPh14�Q�V5�[if ڃh�j��a�#[�r�S���-��QZҖ1��4Q�Dc���*�m�kX6صZ]V�`����v��dhvդӡ�5��"c`���h���c[@j`���BS�ml��5m��F�CK��[XӤ�`�Z�+E�k6p�TDm��MQ�F�N�4:ֱ%	m�[kZ �
(�H�b"5F��X��
[tS�Z��4j�F��ŀ@� IG��E�������ǲK8�_�y>{�P�xL)��:�ul��\��=��L��P�Z{���/z�j�W$��N��{�#=wu��;�`��6:�=�u#���kC��q�Mi�"�7��x7��=��h�$�g���o���~G(��1��e�^�P�J�d�y�p�W	��2յ��2&6<׌��`hH���g
w1x��^��w�}r�|p	�^>⨴�JCus����f���Jw3����S�b�0��o��(�u�9��Kz�jsˮo���O3p�!}�_���]��7�ė�G��| ��Gp2��b)�L.[����{3�]	���l�����2ݡR�*K�meuY��/E˲�w"G'�jFp~��rk���{��f��e��W&`�i�P�TF�K�`��M���.��s�r�}+n�d�uf��g�o}J��>��������=(;W�H���0i.j`��s{^�~�gƕ��E�t�����g��D��0�Is�����'��e�Nt�5�_K߯]:�B·�d{%�t���R�f��k|��c� �y�1�)��d�p�
�a�u?���gV�]�z�\�4�Ɂ�]�e��&��JЄ��C�Ao���.��R�`��vrp������v��f�%̀��D#�H�1¦n�ۏh:�s��맔�9�b3]{��=�`�k�k��f�PP���"���7�w�C�;�]�d<sZMI|T}�@ �<��w��g8�|��Y�qg��y0?|e�ӂJV�3�,NA�o�ۮ�{ҷ��7)%A�#<��q`U3����:Yk�i ⅉU����ֆߊ7�?g��]���"������c�w�%�S��J��n�*�K��4��2�|�>��l2���]s���o{�J�<�2AL���yN�>�f�t�ie�J~uy-�wx�q������S�|��;u��|�*ƻ��oc�s�^����(z�bÕ��(w}�,�7*�C�{���u��5���j�P1{c�g���������v�cO��cޥ�M7�O���j�ݴ^1��R�T�J�ז���S���N&�����V�Zv;�uKǋ0��"��]��!��0߸v{���d�a�Ƿ�p
�f'*����X��cai{&mW[ښ��~Pz�w��e��KċGּ�PU�.�"W`^�3�c�F^����g����OsZ�0�~�23[�&T=���Mo�:��T6`���4�Fy5}X���}����܃$]�����/`~�S���������l�th�_Y��]N�FPL����ǎn((X��kA\�aΫŖM��(D��(N괛1�hTxV7�)������w�/���.*]��ˌВe��de:�6��Z��ý����s]̷ު��s~��W����Q��e#�%�<o�����G5:&9����zT����{}�
\<g��،7=��k{)¸��h�Q<҈�s7-׺���Ҟyk���CK�&
{OgD�PD��2���s�㞺��wS���K/(����{�I���3r��Uiqeȡ����Aͧ�w��e��ܬ��1
<����z�W�`�Wsz�B��k�j|�(m��s�ZV:��T=��	v;�Nō3�u�!e�o������n����x��:�.T"��$�k5�X�\e�C��k�v��Q��;����k�e�3ڰ��e[D��=(C�%Q�xM	|1��#z�w�_�s�_��P��u۪G\Fg��W�*"R`낞�#�
�o����g�{�~×���q�fLN2n�}���8�H����K5�aX{2�y3�>��Ϳ]y�c��[��q�˧g�:��P�V{*��2�׸�>֑c\=��ƖM���&�
`��^fGE"r�ۊMkֆD������p!�<)�%�� ���V��R�N�t�Ա��]�K��[�z�`:�#Nj��Nn���:F��:��y��k%p���.܎��<f<��RRJj�Ntr�U֋������ t�x��(ܮ�4��'�s�!�V	oNK�#�{��u5�c�������k�G=v=+�lUŞ*��X�և���oȍ>�j�^J{����3׭a�p��)�
���r���P� �~��T�_�V��}�N��8m��N�%�j!]���7�����n W�#��<�KU�*��e��e�on���x�viL򂴳,S���f�3]�Z#E���,g�����f��T����C�Jb�EK^Ҋ,�n#��T8�_4=8����g�
�\C:��Y�c��h.�>���b��Xv��̆g�TGX��Ƈ���'R�y��L��fN6W�o�u=6�e��9�]�GR,x�Ŕ2�;��݇��s�<d�<����l�5��53�S׸����("�$��.�:y(�S-̴ҝ��x��z�����uP;w{�;��n�˚���$��~�z�,��!�"���_Թ��B���C$ӝ�`¦��q���`c�{轴��gr�@.�.>�ȯQ˗��d�(�5��o�'����+��KH�/���jӦ(`�Ⱑ�j,dt�V���Yŷ�:}���<o�2��(.���7���貂�D�Ά7���iR�f����ׯF�Q��$����[yZ�)�["t��k��w�p�xc�H��Y�r̮X��{�sb�����N��G,#�VD��o��5gF;beم�H�Sj��}3*�{���c��PRg��^�7��ma}�b�t���*�9�����g�KGJ���AF­׽~����w������gś9}.����и�s�ZJƸ,'(1arzqi����i���"�~�a�do�}֍�ia��<�\Lp_Io�e�淠���i���l���~��=X�Q��$X=oJ���r�α0��.�Խ���q[W�m��$��7=ѹٞ���珻Ǆ��ˊ�c�pM������죧t�-,���,j�"8���۹$���l�"}�7|��^�1:���j���F�����+�Ƭ��p�e�|.�R~��y���YW��b�aB��&�σ��V)��OJ~Brg�Xdz�c-�=�N��S��:wc�Yh��T��$�yyu�(I��"�X��W�S����r�����M������7�K5�z�X���GQ>I��]V^R�.�Qz��H��ByOb#�^3��W�J��٣_v��<`�|�p>�vsr狔Q�O���3��{���X�˕���r4�W���k��rY�w��(�2z�OͼZ�Zl���w��=��k#�6=���m�Ӛy�RW
J`��X��8�&G�~����R#su�-�LӢxi[%����H{�m�'lS0��6�ۊ�Bm�^�Di'�`�[ϩW�N�8�sV�ȏ����{w�A>%��6�Q�q���D.)���"��4�=Օ��s��Etު��� ϝ����P��V8�s���d�<����g��L6�D��H��[:��>�yK��#�PmOCA�^k�OK�5�W��W�J���2d8pL�B0S�q�
�gyd�;�����`)rIq���o��/�>��`\Y�\�Ī,	)Z�&ܖѕ�o��>��k��7�y�
��RJ�JE�`�\E$�V}�E�/�ZH8�}U�ldG��>���>�H�c���<�z�L���ז��n�*�K��4��;ݽ�'���h�흍?7޾EO��%X��\	�z"q��bgzאx8V�J�3wב3�o�q�"�A��7���j����C�^����;G����X:Y"����9�Ϋ�rǱ�8y�`��x$��:�!c�������m��j�a춖zm�ݲƞ7�-0����ә݅�n���S=�ּKf��>�B���Et�2ҵ[~����R<�W�o6{�O���[��d�]o��KP/,b�~�|Jz�o=}H���(�'7Εwf٨d;&�cLl��j��Bre;��,.8�=�MTy�w;qԢv�R��fꋚ)5�fؗ��7��f��{��*�X�P��ݙ��q`���'.�j|0�s�0[���KUt�}<�N׫zE�/�F�XVl��IX�'��N`*�jDp=�0��3:��k�;��U��7=mi�j\<�O�����S?a�F�tȦ�
^�0T�*�S�8����*�w�P�^��D�/��e%u���Ğ�/��o)j��\�҃>u&�n��ٙ�mQy�H9�*�2T�IN�L�δd�,ϓ��^|j5�z"7�����tW�o��ㅻ����>F���E҂���\Ɩ|wə����Os�g>�[ޯ8i��-7,�ݻ�<�^����DV���pB�"���!���BuK~ZV��h=�{��n�ּ*?7Z�)����<ּ�7~�^fٟz�Cv�I&c[�ȭ�6Aͧ�w��zp�f����'S��ym�O{y�!FnV�ϧ�	a�k�Αi]:���z��K�޲v,�cY��1~���n�B��M��տ^g�t��@p\�E�%����5�䮝q�����~��o��GW�]
�<9�x�#����*�s�ĩ/t���&�#Jܺ6���`U�w���ͮ��QWF��� ����7�i�t���r�ͽKu����)�ڋ������Z��5|�g��jګ�s���Nkꎻ��,�z-f�M|D��E���"���২��!���l�З»��n���\꙲HTG�Ѕy�8���������~��৩GH�@Vh�|� ��o�l�%�\���Y�q�bg{qY����O��ku؆wK�pXV�d�L�ΘN��1�tW�����{7Gn�m��,�.X}1T>Ճ�L��wc:��֑`k�ǳ�[��o=P6P����ʜ;σ�"o��W�.[��X*u��:\�z��&�Jv�{�[�c�&31��9ζ��Ry���:w[�\��%w)�U�V�qe."�&G�}w"��5e�"�%١��x�����yܯ�A{l��3����=Mڹ���������R8�3ʴ���� 92�V�}�uF=�D�נ�*�����O::�A����ҔdhuG�����ebiN��Y�6��
T<E֊��f%a�(�ɸ�6�P�|��h{rf3Ē�	���0^��觷�,m��`B���d����ڦ�l�q�v�����5�|*v/[��<��ʃ�����a�2��cK|�\'� ��9��­�^���#�����R����2�`f��1����Qw�}�u�{�S�6���f*�!mX���5+�`����&۔3[�V���b��q�u#+93r�����1s�u�J�{,2 �uKW�t��\\Y𠙗���?!�׭ͭBȚ�s�fs�u#�9uy��wܭk1@"�$��v���@|��h&f�����di�+={��%�}�5��q>��u�I����u���q�	�x��:t!k5��.i�ed�����v��>ͺJ��/&�o�-3�i����%fi�S|dW��ˇre�͛$�iqR{�J�*�ړ���2�[�x�ꇹO��6���-f�nJȃ�o���՝}�L�0��^��-2[�^ʞ����z�"�)in��3`�6���1fwL	+�J�+���9E����ݫҎ]:5-�ݲ8sK��a�j�_G�~��'���mC��ZJ��,"��|��WN�卻yעԼ$�����9�~��0u�@�/ʋ:3=sɝ�m�6{+m���Ik�	m�7���]����+�;Y�j<l=yP�
�F�	��o��'t��c��{ݜ:��<�xX��3��f�/N�Ki }1�|�,�62��>2��7UN
\��g2��=��������jip�
��fd
N[(JO!�tԭ�)���s��^���Q�O�EkIJ��v��z幧���L,�V��p27�C��l�s��s%aל���/1�Պrr��R�戌n`�w���Y�f�ͪв�׫�{��9���ىԵ��{��;�mJÆ`0~�؅��dS��=�t���45`S�7�ژp�7�3�?ꦖ:�)�C�)|�gR����k2oLX����5z|��)%�����`�I�ޤ[+�QX�rY>!�n�_���'�E/�]�b�CcZ�mu@ꤼ��+���J���v^w"G �(O%��^�3$� �?^��l^M�/��k	ƻ�L48�4�K�`�Kb�Ih�yͫ�.�7�Պ��~�Ÿuz�'Z4z��>�<��JՉ��ۻ@��0s乩�%��jJw�����9��u>�v���.j���u�CH�'u�=��.�o��z�� �yY4ˉ��ON.�_n"Li�!���-�K�5�J���2��Ϥ��o�2$h��S�7}�[�h�Nkxk3p�5��Q+��u/����8��Z�\Y�;�����J�+��H�}����jb7a�ɂ��2�]/�J�*�XX�^��0J��$����~�E�.�,������=�t�*�x[$=
�h�8�s�7�iQ����f]\�ռTм���j`�on�xa]��Vn��k0'���P�DgL�2��G)��U�vUӝ���uV'g&,��3�Z>�Kn�q;�Ƌb���aP��^��i��m�;������;��I7��;M�]�����G��=�� ^|��J��Y9@�u��%�d�����Q��ÌclJ�vm��rT�̵��nѴ�c7�K�ǽh�C�>��
;N��wVS/��V"�#�-L����H�܌U�n	��dەf�e�����Ag�Z��m7�C��W2M�.��EP50	ifM)��TYA�P��e��*�Mj-��f��yS ��J��n$7�@��(z�j�ɪ�2�^���u
��k�͸t;퓘�{��F@ל���m.u����4,N�{'���c$�G���uS�8S�0��% ���p�Y,p^�:r7�f]m�=d*�&*�߶���n3� �o��{S�wR^փ0���YS�J'C�LśXh����N}����GS�3��T��V��V��Rc����PkB���eL�� U(<ԯ�/8��H����]Mҟ+܆��j=����Ҥ���ٶô*�==�p`��������+�˱S��5��&�PI8�Г4�@bP1�T����x�L��\U%�10��{�9�FwqQg8G;�:�k-�+zp��� U�qQu����+iI���7w���6�vdgqOE�h���;���e]�y���9�0�׵�s�L�5ӧ��Z�^Kz5�X{]��YJ�����t^8��`��.�\�j�;�Wy�����g3L=�A.�7=����?�7ip�2�N������X��3RJ%�h��>+�(��u_IHI>Z!zn��}طp��&R��.�bWkR�f�M����1]M�O���]n�]V��%q�{�U��it�V1Zt�j�5Z�Uh�$޽���u�2�SV�%ĩ����_Ǆ��Qv�r7��K�ܬ�59�(�k�U��J���ݭd�q��m���M�%��ڕ����ɯW7�x<��i V��I��zm��Q`��%f��o����[��]�f�6�Z�&iܸr�E4�WP���K���&�$�K6�0'��^U��w�/1�vþ6*�ւswd�.Sm��-��/;w)k���N�r:a�	6WO=����$J�uÀ�GM�-Z��[�1rķ't�xn�z�gS�rv���b�u㏧No��K.����3�����j��탍]%��0�3GWoj�1�ѭMŪ��6�Cq˸*��ۚ�C-�kP�ιƮe�Wi��Qpp�A�svpRa�ժukr�ԓ�K�����\�t��)�7N���y��Y�&A+vS�)	��%[��L�N��r�$嶫LY��:ޒ�Ww�]�}��6��(ز�փMh�a�N�vɫ�M:�l1֊"�ڍ��\A[`ֶ�m�4�mF�t�X�LI�4S����5�ѭ������(��D �kQTm��m���mQ��ؤ�Pi�MUj�q4��[d�mgmAcV���"�lQ�gE)E%È�%4��m�Fɨ����Ihѫj(Ӧ��E$(��-�h�F#X��i� �j"����cX(v�N٭��4�K�dj�("

N"��`"B���E�]5E)AE��"�Y���b�6�R�LL�b&�I� ��"63[�(��)-��[i����Z(�(��"��6ڙbb	�������ѭSE5QT�5;�)��5��mUTDR5���T荪Y5�-����j��&��"�fj"�h�S��*"���J�
���Q3@�3cR"v��[٭q���>�ɋ;�
��ڻ�"5fNX��il��0���>u:�R����҄�N-�u 
qģ)�M��6�Z��_�.�P�����7]6�'��>�ז��n�)���%�K��nMf��C6�=�U�s	V�F�p&I�҉��U���T�X��V�h�Z���3g�lN/y���R3+X�ڰ���aқ�qzi�c��[�/�ۯ	�-���/
��W��9��a�,�ެ�fw�z
�W`g׵ؘ��E�@|m추�S;���1�v�`�=[2G����m3}K�ʮՙU��B�n�.���2��E��`����)�C��EfC�ۚg�z�a}k{�6*³e�&Ǚ�\�S�5�jDp��V�b�}V_�­��.Q��k/{k�,�{§�C|}��`��qՊ^��+r�4;8�#�x��Na]��Ys� =˭�O>��=6���js*��\��4�:��T6g�q�VN���k���z��>9�R�T3���FOP������KH��v-��W��lnOK�4_Y3i����=�E��j���\Ɩ�fo����b{�2��S�q���G���z���NW�I��1�{��5���4��-s�^j���Q��(�ݖ�H�i���J
��\K��ޛ�A{=yn�Z�%�r�}r`-�2��fS��e
¥f���V�kEJ�2+��������GrZ�X���fW��6����췞�x�����'-/#
�	q�]H>�o�@uZ�է��s��ئ(Eܿ���ooK��^J�S)�W��4:Q+�f5�"���穹{�P��j��=��Q-8��P�PL�x��eLX'�a�hs�ZV)��|߆��@s���כ��.��㷌N�a�Pu����˶{҄���*	b������\��u�^]��ʲ^��n�إ��$��^3����3+u�1�%a��m�
z�Bh�DCaἯoα��|�y��[��������,	���Z�#0wL	_�H�ᖘ6�,���EV�{�`�w/#�mo�G�Х�[9;s�P��/~$����]�gt��`��a�����t�J,�b��Qn'�rޜ��뮷���T>Ճ�L���2�g^�ƼG�;�h��N�18^�H� <�/Á���+-b5ҏ��k��J��T5��"+<�Y�efj�ڿ=����\zs�#��q�3�grђ��=�Z�i�\TJj,Ȫ��[x�Q�b�}Gy}��ڼDr��m	�+���ٝ��&�Dn��w���b@��=�l�kL*����o�n0��ތ�j�sMB%mv�t����km5n<��� ��J�Ȭ���ۘ�qAv�]s��ù7�O\�5)	Kg8j��D�޵-�}"��1v̄)��9Ζ��]t��ղ��d�u�t����u\ڇ]z������[b��Q|�^T�ɴi�d�&��f�p�S/��|}�j�V�eӹ��'�k;�Y�-��'S��MM��/�8��m>�Z|�R�J�!@�xu3z�Qp���`��:��N4=�G�;��s���GJ�2?g�s�����<M��ł���TGuSehhz)��N����14�V	S�Ϸ����������l2,K46���y"Ǿ+��̼ww&eN�a��mV��2�@���ԍ�i�}�8�b� �_�%	v��5rP]L�)�e4���٘T՚;������ׯ�u��F���I���=o�C�t!}��J���u��l���5W�r���p�5�����i���������H���ˇpL�Y��T��GӾ�i�+��{����m���ꗂ�>V;x܊r-[�Ȯ �˷��CVt`Pç]ZѼݾ�ۜW�� ��/��:`�F��X��u����}�X_u���%rT!Xs1�J.�mC���ͬkV��/\m���ae��l��Rӛ�{Hq���)4���蹘n3����#8<��ŒP��d.�·�_������o�b��oH��Pg��Pvؾ�H����Z�Zv���@-��A���R��77h�YE>3��[5���שGv�D؇��]����o��FϦ�*81�}{D���������ߴ�O�=v֌^��ޏ���w�@lI^kR莭�߄��l�V�/3ʥ�����g�ewN�4���G&Eؙb�Aٸ���h{p�/�=oJ�uܳ��L�^]9�V{i��8��Y�~���;?!^��o^����18���{#�v��i���:st՗*�_���s׼�M.�Z��;X�����r{l̬���A�q��]#[�6o�%���\�_A�ٍ���EϪ���*�Բ:��Rj'_8��̇˥�_UJ�e9=Q��7��{_ga����e��rJ81K �κ��G$���6���.���4�����Y���̑\�k����Tc"Y&aa!��%<�u;�v^w"G�����ż_���N����Q�#�ӱ�`(y�98�rɆ�Y*1Hh8U�p�ORd�h�.cc+c��T��6��k@�������>~�<r �p�H�@�<C�l���l�9�ZJ�+�������s5��*�9^�f^&8�]JxՕoq�A�����`� ���9�C�������{�@�a����qv'-V,�iX�ٕ9��	��8-�׊(��drˍ�5��ފtd݆գ�X�6Yv7Ӝ2���YĔ�8������%��}�/T>l	V8������d�<��z�̞�a5|CI	9[T��̷�7��|l���3�<y�[�4|��j��0k���>���$��ow����`�_m��»���,�� ��5ΓJ�S#�X!���9�����z,�`v���5 �����\u�vdz�_�<uT���&
��RJ�JE�eJ�)&t�Ȧ�-���+&��3����.ʇͱӝy��$�;���`�r�Ĕ���a�z�L�3��{��gh�V2�ܣc��yX�S�W�i���"�k�J���.�:J'�U���^A�
�)���^�8���G���q�S�i�r�}�=�xP�V5�{#�/�gK$P���=K}՝N�Q�.0nJwrj��~��o�+�'�x_�U��Wx�p�x��^��Y�Pe��M�g�a�-k��}���(����R��W���K"�C�f@|/k��+ltI˱��{��QV �^�֟G�����
��]�@�XVl���z�Ϫs`>���x{~/�̧�h鳑�Xi(oE#�$���ڗzzV�T֘$�ݱ0��F#����܌ rw��ж���eQ#�vR������g<�S`N��f�;�r�q�=wԨ���vm*۶,b4�M����X4��T�?���i��E���^�oz����%胉��M�;��^VGM]/Z�W�vJ��_[�d�my:����g4�f�JmB99�'��6���j`L�{+,1[T�K����Ib�7H9��4i�{�m˸#"ik�P���F_��4Á=���ƣY2��h���xz�禖N?',�x��U�t��1�7i���wə��lOs�g���y�L���sA�H�om߷�c1�1�\��Q3v�F�+�6C�<�~s�U�D�L��s�	q�&��.�2�]�K�z���;�sœơ�t��K�LưPL��4�m?K�u�tOL�i6�f��ӷo�/�f��1
9�ʘ����49�-+�x�=�@�1z��6n������f�)Ӵ�[��O�]������P��(Kyi!CY�%��Ϗ�>�z�6�3��{����3�wOu�3%a���U�N8)�8%vĪ"xM	o,���U_s��
G�彍V�&�vxT\��I�Fgt����*8e��?%��;�������&N?V4v���v�����V�n+٭����gu��7~�����E���p��]�`�&P�7�6�����^nYi=��6+�Su,��,�o�C�� �cW-II���R�U}�t��d�X��q�=����+SUY[+��I�2�ANY9r��)�&�yj�A�Fz��9�~�S>�Kȟ-�t��SՔ!�ʺ�k�x+#@�Sg؄�s�=���A��+��ʸ���Ww�˞��>���/�Ej.o���M����iA6�.K�j�nmÕ���G�m6=�Ba|G/@��N�F��^�n7�������IvG�=��5��Z2Wr��^^>J��q)tE���=Lom�K�ð�I��tFysJ{l����>�KPχ���Z3��6�VȰ�~0��ke����E'~;��ʫB|���ͳ����i���g
w9C����z�{����PRg�f��F6��|��q�U��
T8����K~{J(�M�a�\�r�����:�̋�/�5����<s��\N����q�`U�`��:�]�V����'R�<��z�.燐��k�����P<�d�a�r���֫�u"ŕ�ş
	�we��_o�	�]"�G���Ŀ;a�n����7��pD�%.�4�Jk����3+һ7�'�]���{�z�bD��b�@����;����քUie�[j����ݻ2A9�n�R��~ �G�����{����D{�VvDq�Y�[�/Hݫ�*&��X�n�ٮ̍�<Rb���G��j"�;B�d9�9g4w9�:Qh1���k�W�ýh���p5���&g�N�|p�� �eD7�_
WS���̕���Gz�����C�l��ϣ�5�Vf�������Ez�J���y��9'>��{�/��$��KJ�^��}v'+��Ƚ:�Y��IY~�˷��CVt������y��ޏ���.�/
G��;҇e�^�6�k���b��a%"d/���e#ݺ�k�������F-R>;�˸p?R�:�C4sK���nx��ڇ�}.�l�V���~����I@p��t��u�W�	��q��}h���@^tyT�U�w��<��n���E��Oc��|���x����5�%kۄ�	=oJ���q�5ץe�g|m�Pz!8���Kӵ9.�{�����j�k������aqQá�x�	�cuz:��{���9��v�p7���9�]�l	��G�j]v��!�A���N��:������찵vO^*޴nN�)zl32��x�E�[j`��R��P��h0{�58��̆�Ӄ(x������m="��R#ݖ��rT(P(,�7k`2[�7^�5�%��4Uc�]al��Sc�*PZ��7}����c̼�ZR���$�wNe��5����6�)�J}��+%/y5.?����N�cq�kbh�p4oI3��|[Ӯ�9���O�Tu­�a�=�Y�Ib���+�-�rKlh�8��w�QU���&յo̮+HS��lA�����������f��'S����՛6%�����������+)��T�~���
k	ƻ���hTF�K�`�Kb���zU������F�=���N���^�V�#��=z����<%j�R;n�#�l#~�y�����#�ķ���(oX��P�sW���u�E�'?{�S?�����ǁZ�_7W�o��������}؈��Pqo��}��]�{�s������Z�<&^����_A�&z&�i�����p��*#])4�}T��W��}��8�>��gˋ=�����.̿wBw��o��C�|�+^$�9`�*�I*��"����U��hj�觅x'~��qm�����v�|����\P�*�:�<�%/'uA�����}�-��=1+�W���oo�\��}ެ~�w��X;���\�SB4N�)�lt�}o*���� �˃�E�(�z��AS�ZzJ�A<,��m��o(̩�]l��On���E���H�[�KZLf��Z��y톳>q?BQ�A��MkG�sS�I[���`��Q�A��a:v�A� 	�R����Or�T�����#3��W.��s'3��G$7� >ٴg�
ߏ��E�{^�<�t�]�Q�ǈ×�wS��{�ڃ�yJ�ɲ�~�X�����,���w�Wx��xǢƠ>6�ifs�"�gi��s�3��H����ӷ{�
�zN<CUfK�]O/ײz���h�T����(��"k�F�z��s/�Ӵ��龶�融�6*ŋ)u���C)r�g /`^�ؚ"����1m��r٢ =K=�a�˚�q=^ɳ,����"��F��^z�(ګw�����ŵ/I��MH��jD�T"�Nn�ʛ�gDf��E*��`^4�g�/�2[�R��:�
׃��}J�<z6DҰ��3|'b2�i�������}2���^�/���Ƕ��Z8b���$t^���oXwə����=�Ş�[ޣn��y�IrY�c3��~eqq壦�vh��J"}�qv��w�1��y���ߦQ��=�:]y�m"���M�{m|��X��`ZkF���tv�N�pupw��w�\w�+��Q򈨂��QQp��+�* �������Q�ED��ED�؊�+��W��TA_DTA\"�
�DTA_�QQ�ED�eW��TA_�QQЊ�+Њ�,g�(+$�k8A���"O�0
 ��d��H�|]�J�*UiL�Ii��(�k�@�U1�kf��ڂi���1�ƩQ(�5[U
D��%,C!��kU��6`����*5jj�m��l���1�V�lz�]m�ljګ	Fچ�[[J��S5�"��[ce��مl�U]܎��"-5�B�V̆��MN�;ѭMKRƉh�5JT�m�ͭ5�6P��[R֍�Md�ձ��L������&Ɍ�K6�ژ6�Ƣ��j�f�����cKM��j"��zܬ�����f�   c� ��.�h�낀;��R�۪��:�`�: W�:nm� ��� �i���:��.S�KC����)�֚m�x  u�RL�;wwT$(Wq��;vN)N��۶��)Jg&� �� ��s��� ���4����:�4ՙ��f�[Imm��f��  3{֚׀�;�OxP�B�
(^{��E P
(]޳�(P
(P�n�w� P�
(Ps���B�
(�g=� 
(( P����(R=(���@�4-J�Z ��m���h�+V�#-mkml7� �zz &�	P)[6u� :�Ƙ5M��v�)��W]Х@�V
��M9����(��Paڃ::�mV���V�m�� ���q�٣AImcM (i�[�
P����m�N�
)ѷ)� vm�T�p`(ڻn �iT;�U6Ŵ��+j������  xP��x�:4���M��]�n�#�h.��:l��p:���9��B�mƷ(R��8���R�NR�����*�Rf�R[3� ��  ���벀���΀ѥi۶���U���Ъ ��j
���E���h
������`"�h�l�Z6-�j�[Bư�T�  ��%@^��-�i�5Ӆ v�ܠ q�;M i� 4n\�q�n�ά  ��
b�lkc&�Vf-��k   <��hn�p �u�: �]�@�V
 u����:��ks���t`�CLe���L٩�����jι�kL�   f��@w. :�V@8V` ��t Pv��P������ʶ;\ �np�o 5= ʒ��B)�IQTd#MhE?S�LUT'�i�` �~%JD` �0a�`L4d�&�"l��� �������h_�������Պ�|^�C�Ӑ��?>8�g�n�����}O����$�l�8B�r�HHl	!I��$�	'�$ I!		$��!	�����O�~ �~8�ǖ����E��O�Jo� ;R��K2jP�
�w�6�Ŵn�P!'���[B�l/LG�v��Xt�
�P�2)<��c�)��b�Jz�%�9y�F�aZ�0���/D�7e�N�*��XĤdwN��{��H�]�0|D�Uz��,qZ͢��!�r�[v����LZ�!;�����.ɚ�	�u�E��V�CwN�b�X�Y�P��"V�X�d1TO6�b�,R����)�Mm����E᥈j�Z���ԗ���,�.U���%�R�� ��B@�
���^�P�p�������j�04@W���n7�R-�Sl����U�[`e�,�b^l��O]��F��.��b�!��4�r𫡇&+:�1�0��&`��Bn��?h��)�A�4�dW׮�dg�����ś�DS�0���Ō6nR�<ʼJ(6���!��1��-��̸ͅ�Z�U���� ��HM ـoP8���!�i#wj�59��������+-P4��y��� �o\��A/I�&��6���V��r՛@�6���f���؊���B�m����&
�7PH*�!҈=j�޻��X�
F�E6���e�
`�H��J͢l��ڹ�F���d���Fd
�fa�$�B����n��E���B�%m�O1>Gw�k�+r�]u�p|�j�+M��N�^G���h##�����%��沠	b�����6]a�r7zȅ��(=�`ڹ�[_B1�9!���u)��{K�7� ����p&DD9�W+��WQhŤ�p���j�k.�(���m���,q���[t���,��U��Z4�ˬI�Ӂ��^zCq��djU��v���7`�����;��e�I�)3���m���CNP 'p�x��3 �Vcu�6����7Th&,2�/@�S�{)[�f`(e�Z�P�[:���@�2v�n*� H�nn@ZW�Ő=��J��}�I�.� @Y���m=�k~#J1�M4��^����9Oj�[$L���ѼN�65�Iø�iA�J=�*G��Fh�b��Y�Ս�[�E�+5����SS��=X3F�OU.,�YA�A��!�m�j�*ƍF��Ň�3b@����?��<��X91]f6i<���u$!�`+G�[kkS�.���j�4_Ă�a�u{�6e����Mڃ)�Y����v�X�W�R��'��B)�1Q�M�"�ǻs^�V�U��An�l*v��Τ̵w��3R��6�	P�E�WQ�U�d�Uk�*³AC�ȩ��Ƹen��u��\@`���;ݸ�w���Զh�	�BbBE#S$Ô��m��z�ƶm9�)�wor��v������%�Ú�yl�˂If,�ic]:e���F��4l �6���Dmb�,+��X������ ���+"ـ��&^�E��&P:.�	�f��m}�ki��U��f%D��v\��g�C+1S�jJãob
�-죸�]��Mar[潩�kҌ�btv����2',�`[y�8�HF]`�]X���F,if��n�/�%�L�j�KD��εB��6�0Q�]5��V΋Ӊ�1�͢�(*��I��ij���ǉKs �@�c6�c���lv*#����0<�`���ŏ��J�3 �y��	�n1���Y�*�D�,�B�R߈6����n�:�,K`[rV���U�+v���űcܧ�I���M�j2��f��m^r��9���d3v��(�-L�	ZiX�����'�c.V�V���d�cZ�w��{7+DT`�{Y�lX�{qM�@G�e@�ٯBP�2�|�U�%b�IƩ@����f$f�����b��y�a�k�z^�}�� ��
Z6Խ��U\pSB��%�+rrl���N{ �L�#��n�W2h*�qGi��B|n��1�����sV���C�l\VݕARv�ca�ݺ�L�"�b��fܒ�+�ON6��7�E�oI�j3�\���t	Slڎܶp�&��N@�(�J��ȣ����p-���ɵ��C�˶�em?�,z+&Ūۍ�.�xL��ڰi�y%-��Y(TC$Tq=��Y��C�7.�kmk�ڸ�TSEa�n'b���ֶ��.�"�Ȟ���@:�і÷�
�u(��q��f����\$�i�����d-:��3F����=R��P�ͣSZf��� ��F��jBT��skV��)�Cy,F�O�a��IEWuv�*k!�jP� ��/7V��R���4;(��"�5�ر��/r�نF����K-���M����b7��{�`�Ɲ[�d��b���ǌ��2�������P���K1*�����BmV5x���t.Y.P֭�p��K���:�%6���ݱ�K�٥�jXP �b���7�6�lDp�r�
3��eL�㹐a�/ouJͻ2Mn����*fSX�!S:tbB�5$���׃:��cʽ"M�ڒZ�E�s#A�5d{,T��
;SR�#ϰX�6]m .Щ����5���	�4�#8��`#-9�p��\�M����`D@/d��qR�n�Kj�0�z7��W;�4���Sy�`��ŢI����:3q��.�u��Wl�r�!�ź�*q�,��agL�*X.*zT��r��t㖭��=P-�ml�{Ь 	��q{�����=�K,/tF9Ve��Fb�Y���r��O��w�
q���
�*�;vTf�6�ƲA	�d�	�ܻ6u�^+.�`$V6T�z�4�+,sI%Kq�}$�M[��%�^L��!��y�ùCf�͊�Jb�oJU���an�V◵e�̷��4Rhi�7sr�"������(�X(�t����krc��ɎL�%�c�{A�$gX�=/�$(5̎e�7�!T��d!�ؤ�8sХ���E�xm�J�p���k^�v
�2*��Ů��,�P������l��֢y���SK+���(��ăU�jɩ%�[E:^k6aDK��B5X����n\�p�٢H�kv��aV�M�c,��ҧQ�
K��3cr�Q�#�T��S�l�K��������.�ѫ2k2T*�F!�K�*��E�2�� �&��w�f"��V�H]�\�G����)��9��!�Ie!��J�@u�:.�a�DP�NZ���dR/���aA0�`-�C.&H8%��Td�K>-aۼ[[�SD:r�<�?�wN@l������)mF��>P�a�0*�WN2��]�n�.�5P0��mzX��6M��YT�N	n�n��2RӬ<t�[��l����9��D^��`I�N7�O,��������ѽ��0��#�_F�/V8��ۣA�[�~I����ݖ�T�%iV髦�*��ܽ������jA�ͬ$ى[��aZ�0Q��0oO$�Q�{	�A�0(sg.�o�H7���'(� MYA�݃x��*c�V^��� )K!5N]'b�XU�t��nS�8)a5�A�~��=��Q�w>z�W�И�)�	����"�1y��Em޽�b8��3���vÔf���s�V�R�9N��'<n x�$��ՕQ3Dz��P �jf���&e`A�{���A�u���?a|���{�~��&�Ϛp�������ǳ$�kOHRbF<Њ�n���˭4�я#�Gda7.T�z�Uclښ]�WQ<ũ��@4\B�A.d�H�������1S�1D�`�(�t<n��[�8X�J��A	an���LmڴFӻ3+p%s#�o~�b/&��c�$
h٘�c��(��Z&� ��6Ҕo���ܚ�met[��II&72�T�
�n�V����V��][�M�w�@z ,�U��ׯ/koJ�4Z��՚s�+;j��.��Y�*��`TPIt����(/6���,Y+^�Ѵ�V�4V:�ݘFdFn�U.��R5`�w���1!��S���AEQ�F�B�ͭT] {���}v�E-5�.2k9+Q�x��M��-���l�S>��߹��\|�QŒ��I��K�&�b��M�����H�3�6����-dl��7]fF�M.��7�B�ܲv�h�:0<\#��A�>ңz�,��������ʶɲ��s5 q�l�ƷP��+�V_m�p��ia9:�:pkǲU��-+ōYu�;.���JT)��G��(ZW�a�,�e3WH�W�n&�޸���cC)U����n"�lն�0]7Gؓ-�9A����l8`�-5�t-ͦ��B�GzG�8�7����L8�/cpA�L�2fF�v�TX�W1�m��eM�w� 
ǚjEi�5%z~�s#T樥�YH��*U�����R�&��m���m:YZ��h]^KL�PTJn�$��г!p�#Ǉ��,c�uGY����kJ8�՛�<�[�#ʻJ�mͫ�l;�)�j�cWSl��-4 �V[J������܎�����*j&���77X֪#V�
ݘ6�2n����iBd��PO$����v�;cb���ХM1A�WAU��
�u�Xo �guF(�ϔ ^�q&�%0��&n4�-D�he��2�͍�@[���K-�"�6>k;��0�1Ea���V�@) /f�ah�S�4@�diQ۽w�n[�;�"%�f}cVjm�p=�(RjXǹl)��)�����1!��Ѱ��Nn�y,���0�ݢ/Y%�-�2�2����ԭU�Q!�U$p#�`�@÷���v�	1^�󻵟d���u��xj0��+���=���kE��R��k��m��T(���c����X����\��Ԧt��ڂ�3e0�$sˉ��;e<&pݧ}Z�m��K��nK)V6��"��C���Xp�YtA��4�e�3(��2��k�l�.��	g8+��'����9�c2������ť�j�+{��	ÃU�ɬ�S�,\��Ǝ�A�4��h���e\��&	V.e`a��LYљC)�r������,ڍe��,2қZ q�'JAY׺�yB݌���S3V�rn����{R�R'��5�掱�+�j�N�û�nN;U�ի�u%P`�yt
l�GX��CD�e�4R�(^�20�iJx�Yv�JˣlE�ٵ�*cl �d���
���Ej�r�md%o>	��;>?#�ݼ�Y,��1�Z�q�Au�xˀ�du��R�Ă�v��fcT�F�
�T��p���Sc���t��~��Ȱp��瘼�{�=� ��ǰq?#���4�oۏF���� �����8<{��#V��b����b{�5O��n�Me-.���J��w*1�/l�)��'c-���NK��ʘ��\؅^1�^�Ge<d8%�P��ԩ�X�:a�b��w[e��N��9H�gwNn�m�I�V+4��p4��CÅ*��kw!��(��[e�jX��12f:�0�I��*ք�:a���,����a�.��c�^Y�;�����d�dS�/0Z4kib5���95Ij�-�d-�)D�ێx��ÜY ��jy�>�f�m_ɝ��{�*Kqv�6wjfQy���^Ԙ˕j� VI.+2a�7��b@�M���d�L���@×����N�����e\��ڻ	���HR�-�kn��N1d�����m]Hw3Un��yN7�I�:,�@ѱa�X٣�(�⎲���,GZ����$�7l%ܹn\C^�4��!��&C��4��a�����N��R�b:��y��Et90� �Tux�ӫd�wՉ�&�4T��ݷ� �|��Z32��D�)�ë��]'W�V�R�e�SW�*����+3$���0(�`��;D�&!n� �M�t��v�z�V�Z���F�"�3h�5U����0:���[sm^JU�E%.-#1fT����2-gxJ4��4�g��ѐ�1�a�}��¨E26 [�Cf��dK;�)EI����
� ��c�Tg
y#�3> ��y�|V�	p��@������� ������4J�bk9J��1����
%jY���j�G	3i�m<��;t��Y,�P���Ɩ�ⴙ׵�橈dxM	�R��
�h��1a�y����Sh�f9��t�Kam�� I^k�3�J̖�d,�Z��D�Q�sЙO*�����@*���R1L���\��n�u:�H6�g^�Q��S*��M��E�����Z6nIf��qЄ���4é��nݲ��SZx��[L�����A0i��t)M{��7u1��F ��sT�	,^d��6�Qn2�4�]f���U��%O��Y�T��d	|��E�j�
�T0⡒��	��q�zl5ytmm�s�A4Jߑ���at�Mi(R�[��a�w+o"��ܶ�%�7kf	xv�A�l�0]ƃ4��`���	*�9��f��kG�\�iV�:&ݻ��	�V����4`� ���BC ӳ8�YU!���,�I����q�����Ak���Ƭ��I�6�m;j�-�I��iLҜ,��(̘f,��v�bI�p�	����*xGF,n�Adk�m"r/������f�T�[h��G4�(&�,:���0�{J9N����e$���K�]�	[z�������6�)<�tP.0К�[bޖ7bF�0o �ݛw��nG�*?JP���b��-n��Y+��fj�藲5��mAn�跹AaH���v�ا���ң�{�nĻ�<����t�-��n=�G,�ķ��_�@�8�dG�^��*19��;�	�g:���zh��k��#=��̝¶4�����q�ڄ�r[�FWb���9<Q��{b�Hf#E�㻷.9�R�˯;���x��Z�6��d�y�6�0Դn�v55;vf��u3+��Zx��]����@�}���b�]J���{m��
SH��K��ua|�3�S�M.:�܉��y���56e+��h��x-����8�wX�|�o�@�mX})�]����]�}�w#�n*n!o ���Y�q��6�`��C �aO��+�� �,^�MS}$뎷��ܮa�{��N�wN�� A�%�b믮.����kݳ�@��g�	�b�;��P�A��d���m9���Kk-_���t�������9Ld���t�_�w,lز�o,Y�u�)�]1�'o�G{mS���PNc�$N�6;('���R�Q��g!�+�5D�2*�xm�`Rp�K8Ǣ�����+���øf׮�=%�Om�o��gL��C� v�M�K�fs�`N>�8)�bY}u���N��}X�V�mp�0� 0�����!�FD|�:hU�A��|vD��:�A�)͵/w�FA��ޕo�j/W)��V�6z��kݭ�joeu}B��=���� ���x%��+{N�	d�-�Ȟ֏_[|{�o�~�I������tI�m�2�U����c��Π��U1�b[�mh�O2���'���7q�7廹o���m�y咼\���ȣm�7�ԡ�GUy~x��t� w6�	t"�tF�q�RQ�����g�R4��PB����S�ǎE�x�$��T3yqhu�:<�
GAj��E&���n�YH��������T�w����*e*_���2"1NU����&-��9�*�\^X�sUBr�%��n1�YSbf�'�g*��-6�&_@bszN�m{��%�����Y��Zm$����� ��FK��a��1Ǯ���o3���>С�I������-�����ta�\�<g�}�,���-�~�^);R��6��4�2]���"AP���г]�u���Z�F#�h&+�я=��Ʀ�$�hR'6Z�!�^���{�2�&zaSqy��\Q��f�'T�D�]�}�	�e��BR�L���t����xg�?S0�zmy�l�1r�Vճă�n=YOv�&�!.����M��@Qɿa��7ٳ���#�<�-f���y����Ȗem���*�<+�A����˒G9���^�|���@)�>x� k�:�ُuݫ��P�D�)Wg�������\�l���[|�N��1���E��a��f���i��k�\�sj������2 ��uW[�݉&��J�xy_7�/y4F;��DRҶ�����{��ܩ�+E�oB�#��<��2^.w��1Չ7@��ޭst��N��l�:d1��%7o)#�[��g� )��ո
�S�H���ņmX�cˈ�P��`��@w��w�T�Į
`Y�QW�=Y�P�M��nG��a]CU�{�m �L�4�	������P/gn��Q��v�73Q�(�����[ǹ�Gyn�	jv�/�j�m��m�g�O���0K{�u��kp�m�3:�b�ZɃ�E0���U���TCk�ɔ/ޥn�'Ɖ���HOv���2m��ʹ����$Y�'��oʦ6t��Ğ;�&l9�'���ʷ)��]jlX���Px.ҡ�XmO}qx��޼�nN���!���2�Av�:�-�1]
aҩ:p�8i|{��рtp~�����
h���,�C�p[C�D�v��9�vV�-X�b���|����	�s[�kF� __���b�V��$1H`������m;#���L6�@�����4����|�k`��uJ�qf {�������$7� ��؊�0v�oSw��uI�o �1�;8�osNt�m�j�	�S8=J�)ej6p��t[c컼wG���>j�&&�:v��ۭ�DEy#Z7��ٍ�=f�z�����f�`a�**[z/�ښQ�W����h��!s	��`l;o��D*P��3�
������n��vu7nTtX��ݐ���W�ކ��n�I����'����Y�t{�c��v\&�(�T�n3�Kz�O`ս��,�D؝B��ՉR��-��On�)�B�a\��q���a��ŖǍ`k3̗���~r�N֝��F��Jv̮��kZ���6�p�sl�����˦�e2���c�ٓ%$���E�*}�S�n)���X�X0���3�����-�m�4F� �ao�q(�j=Wub:,tmt��
��c��8M���D�T�՗a�����M���h����GooY�E��mpN�������U������+�6K��曣s���e>;܂�:��m�W��-�=�iԏ@6�7Yf{n,Ao��R�d1z]ـl㜕뱴��k�]
�k�B9���Y����<4$�R���[Ƿ.V�E�LT&B��|2��,��R#��Zi��6T%�1��us<�y�*6��ˎg�ǩpu�m����>�nEsNms�jıxn�K�G۳5[�0vQ��vnљ����Z�|W8w"ޞ�l3ܻؐ�\�{%�WU�է�N7��Ŭ�&�fy�n�p�L�"4�u��)�>�T,���v���͠�S�c!Z�=�6���e�N	պ�>7���x�z����}���0�*Nn�؂9\ȕn�iӐ�ܭἾ��A�oV�Κ-���i�-���'��u)
��;�vᖣIc��������U�1���vp���f�Ҕ�� ��2XE������Z���G�����}�]�եW������j�_��=i˗6�h�����:.�r���%�w��Z��V��]�7meq�m^�+�*�m��݈>)4�V��Sۙ�D�SUX� �~�ORR�AVU�[۠�7 	o�<�����{�����Ww�i�#a= ���ʛТ�|ͫwX�ل>�б&�n\C5N�wz����؅˜C�~͢�m_T��c���!��/s��M�B�OobD�hѬ <�A�����Yq���q =�r��u��*Я��~�q/N����V.{%���.E��Z͍Yy�Ĭ-U����,9�j̆���Yt���W}��3�ox��4�Hl��ƦL�@�u'k�����U�ȹ�Q�M���-��ur:hD��ln�8�u�k���@o=|E�md�)RՇ�X"��.�P�@� -���t+n��P�wJ��b|9�.��V]4�}q_>�����V�e�x �!��~�s�4Wg�m[�(�F_[�����=��YGv�G��S�t���߼eƺ�=�pJ\ʽ��r7�η_%�/�}�����#Õ�W8j��%D�����f�ӽ m�Y{]wz(3F��X�����.w,��;�4��sz�/��=��d3VR�S(e��ӷ\X9��oܥO/kquٯ5Տ��رSU��-�uj�X3��ۗ�&kL�����o�郉���Դ���{����S�]�=}}�hb��R�iky�`������krniG�a����n���ځ�tĄ��q:�	B�.��8�fldPr�!�t�ev��O��U�J*_hn�l��p��9����%��Y�/+�_nc��9xH@.�2w7�����F���J�-�Ԟ:�>�ئ���Dj�ށ���5��È[��1�Pb*HiC�c���q�L���>�i�g��m�c\��Kֲ�u��~�;����o�
C���ӛ�F3�ۋ���Y��\7�X�or�����ҞBv���`��wżٜ>�m�E�ÊrB����K���b��_5B�6�j�3���!p�~>=-�J:x�}_`��{���[�{�]����A��1�R{P�Ԇ����dc�;b��Rv��i�Q��l؂gc1֕GGv��MbD-�]�rb��ǁ�s��1S��&���;�� �ԃ��G�{��\�U5]����U��/H������wsy�����z�D!ɷ��s��vޘ�q�Y�n����N�gK5���MI��d}��͛#\�o�\���Y��5�;�E�4n3�2l�)��O����W �	D^�[�;�e>���E�E�q�ux<Z�&�j��w&�����=�p��{v�u�u�d�-лQ���VP|<ۂr1&���u<n�[�@8	Nad,��:{Kݥi�9�q�g�K���"��՗5�V��]r��ʰ�ϓ�]>=�]�>�ý��CG��
5I�5D9�h�媔�۽�7�J�,�̳���jUm����wkT�=���g!ᲿdR)����x�W����ի�{�}��b-���Y}�������l0�rd�7bn�+�M�;�.sR���ln>��y:f����������� C�]�-�F㗰�@�V�t��oR;��{Z$���Cv�����Z�o�i��ͮ�^It�nDX� ���;5r�s5��
h�H�Г�5������gJ�h�fh�ujN[�wwo�<����`���({B��=��ϙ�� �@��D�m��#i}-�A\��Q��ݗ}=ouv��z���rdA��e �W��Wgz��L+Ƕt!;EgYX8�Dr��.��xn��f.����4�CtQ�}R��Z0�n�'Y�q�Y�'6��;�I�
�*J�O v[8�	�<\Qq���]�B��6;�<���9���I[<w�t��#� U_����q/*��F�`�O�(�u
��7f���3�~M�~@g�l�ޝ�r�'i���¨�Q%�;����[{�܉Oz�ew_<zj>J���5k<v˲8��D[�|crJKw�c��F=�o���`�̈8��ޱ
p�5de�w���'��p [�٣^{�@'����K�թ�z��R�[e��p^� ���	���u�P��m�)1R �������+��+*Kɇ��\�=�Y���H;3�`੄%�뫈u%LN���&�:&)�xO(�\��l��)�ն�w_n��T��k�F�*㔝�V�U�0����rSm_d����P[.$�Yv���α��7<	����El���qMD���Z;HETn��S��	1���~��).���g��m�p��u89M�}`>���6RE�o�R�D�N�$��XnV�5�3��ge�:��N5�ve�oK.��
�Ib�(��Nm���8��g���)>�[h=��4��3� ��J��\�8�z��nhl��0�;���69,�=9vӳ-��/��Q�L%�T���+�m��5޽�:�)���� :��bv燉�(��d(�;�D�<2j�d~�Nҷ��I\;�F��n���ɖ�;j�r�=]wslTj��
�p�%.�H�l�૞�M��_lAP{7e�쨡�{���H \������A��j�+��J�I�[[%ܫ�L��xM�joΊ�vFt���.Y��w�V��M{���?Lwٷ/��t.������ؽ�8R7:W�5��=v�������,��]G�
+�R�Ⱦ�MѠo��D@���N��^A|�n�%və���6cK�4!�y����-��^���JLu�B�.���ꗣ[����ݽ�^7��l�����^�A�[�sV�CJ����^y��
٣�]�A�S��6wno\a�8Y���a��󼜑��f��;�����<������Lh�G���CRB���G�l|�޳���W�ơ�m�O�D��tPܰw*�/��}��D��1!��-Y�	b�jWV$�&/P�� ���N�-}�~�tJi���!7�回Sz;�67" ������j��ϊ��:B��E�f���]	y�j�մv�eVI�HZ݋�v���̘01�s���ϳ1����r}zI�/5m>�g�S|7YMA��"%�N42���Gs6赴�F�����i��ͧ�i��Mm�p�|x���l��M�h�ws�����X1�,�jz2j�8U�*kYu���L�uL���w�9aS���;�x��O	y�c��Q�W:V��c���ȧ�i��?�fV�}��̭�� ���O
Wn���M�U��!�]:��_� ��V���W��*և��6�V������	��Kq6�t3�8o8����
���^G�i�OKGc�.�&1Ԡ��(�ޭ<�P�.X�{�*/]�ڒ�P,Ń�*H�]��&{�έ"�oj�kX��{�/U�*�DU�b{fI�6_�-�g�S�9�|V�;��C^�c�^���V3LK��pd;^��q1��.S�lT�X`q���0J�{����=LJ���i
qۼ��%�qxF���y�3T�������v���jn�t.���ݽ��!��:fj[.�s�+5�X�����w���|���x/ԅ;���,e��}g%ʟS�3�<��x�t��N�c�����$�X��^��|@1=7nΔ
y-���o��zKzU\ٵ�qW�Tpw�������;g�sd_R�sY
c���o�^o��C:�X���n�Ր���}tq��:�_$��3|%��ݨ..�m-��zx_d���EF������$����1!�A��}r�|6\�\��
�|aԚ��T\�i�:=���a��(g$����x�r��N�<����$�q
�Nn�-�#�^�`ꆣ��`�/+!�Q2a}gD^���L��xp/�\�*M'i�i�]�'�͇=t�?C; �ON≊lr�a���v�j�JT~�?}��HB!!�@�$��?���`�t�~;��R`/�N��ue]���U�����u��Xh�ayͽ3�{���'�b鉕�i+�ӽ����-}��m���u�$��ed��`� >(,���g���{s{T m�3�݋�����E|�~�ݫ��C���ik���}�����ݼa�X(�U-d���Q=���)t4qǗq�K||���iC�7|�la�P������V2�ks�#Nv�V!�VLy��؅���o�ڛi�	uG�{ �J��)Ժ���c�d������M�]�dޚ�`⫰��*V�P^��kV��%!�n�^gV+�k��]uU`���jU�ڂ���W�݋o���,ÿ4�9��\���]jP��>��X�9P��{V z뛌���X-��A��1`|�ga/5L�n<4���yBJV�5;�;5S�I���.t��A�u�6)��z��0qy`�/��wW�Kz���W��򛗴%��]���=�>�/2F�m��]*D-�
�rN��pil��Ū��:�8榀Iuʱ��]�\����)­���� ����eG���$ݦD�Q�
.h��u�_+:�ݫ'k�@��[1�2��6X�5��}v�s �t7/mL��u�]�9b�I�ɳ@V{h>��0p�,�����M�dl3��)����ҫK���;����P�R�5�����h�v4��VL�!x�%��Y�Äo��+��t�
�s��F�J��՝�X�Kjv�N��';#U:��.M�i�pC���Rtܙ���k�xN��`Z�f��b(�n%�нTwnV'����� �Uy]vvw�$���b~�Õ�݀�n�[{�/G'Z�I�F�3�-�nG�[�ր�J�(L�8v�&cHlΤW5�ya��7e���K�x;|"WsD}������{E��<(]\�7syU��M����,*9խw�Yg�v��t���s��`����n�������ʗ��=�r<�f�&�;�;e�<�i���-�y��CPtj��4W��z$�b����{��\��Ž�l��Bg
�*Q��]��\k��cdB��R�ۭM<�k������~�elu�,∂�5�Z��CRˣ	N,�$4t�tM<�96��h��<VR�d�M�m�;@����,���gp�"+����}�P���h;H��U��\'\ij�3�k�ű�7��Y���D����z�i�U9Ǫ�άnq$S�]���Vr����㗶D�z�3N�9E�h�0�.�D���K��΀�P�Q�_פ���}�^1�t��m�=�*�ti&��Ҷ;Y�#X{q۰믻�����7r�|Ž�=W�f�@��XP���w�W�h񫐙�4�Z�!P��Ϊ�,��)�1�ogfA+�;|bG7�'��ۑ��p(�vCc�c<�r�;�\O��(^UnK��wt�#�[M���u2)[KNWg>�¶�j��b0ī���z��b����:��:�(DiF)6�r+��b�zy㜸)�L�s;�ẗ́���[ա�h�eXt�o�����-tB���iN�
4"c<��3:�@S��n�5�F�F���}q[�Әj�s�U��#���|�i6�WS��v�c�hȋ}���P�~�2��J�<3j2��in�RS隖+�+n��9�)�o({�q���'��-�UfټF����u{x�Yq�����*�$M���#�K���e���[kX��p:��%<Gı) ��9i��\V�g�G��Gc�L��}k����XAC�:!��K��b�S���r��
�Fd��;���[��N�c=�w�Ԭ����o�b׃�
rh�byv��vi��L�W���<��J�Է�E��]��ٽ�ìt���8��6S�-8��[�Y��L��j��Y���˹�Xʩ;V��)݊�S̫���B�y��+V갧oa�h�n.:4�{�ŷj�w�iI]炾|a4:ff5�+0v���
�����h�;�J��M݀��]��*�Чf�sXi��|q��o�JV��e�|�I��픒~}��ɹ>�96��:�u�� �&E�N�����hH����,��ש�t��|x<O�S7����i2ע�eY�guv6����n���b\UB��4�e'��=��wGL�V�WDЅn_Q�5��*$�`ߘTt�ބL�&^A��X�]F���ַmS���d��uY�ԻC;%�����煽�*�7i���	�R&a�H��_j�oK��u���z��[����obř�wSk���#7�mc����hիT�9mTi����n��hn�|�\�VD��,�4Mc $�×�3:�Gt��oFLk�Y}g9ﻒ4
�ԝf���N��!B���Oh
r�� �P�z�F�ᢻ^F1Ce�ǲ]���X���7O�	��V���I�<#���ܰ���Ի �|�dB.��������R|_W��Q�����*��UKV�չti���sl�'}R�W-�l��\��{N��w�ѳ�q4�↹�NoK<+]9�P�V�NW�c*>u=Å=8}e��8-�hWx=;��W|�o���Y��r4��b��e"�'�g1���;��͝vt�HY��{�a��<�N��E�-QHm��*Kf�mty�YgGoq��GYE��+6���ĩ|S��*ɰ��e��n*ê����u��{��3Ϛ���;��2^�n��l�r�O�y�&�a��@���ٛY@�uANХs��:�P��<)�g��xtIl.���"�P�u^�G��mu���c-��y���7:�$_ˈʽB2B��WQf0]�g���Y�a�'1��yt�5��2��(�13���>�{����ـb�,u���0k]Oj�nT�-Z�_=�k9_ �*��8ٹ��ƺ�"�u���mW��2Ak���޹{��/CW�m�ý@m|���x��$������i�7�g�:S�}��ݧ�{%��m̷i!\�E+�3�#����&xB<�qe+v���E��lMm�*�W
L0���J,� �]_n$&U��2�]`���S"����֣y��I�`�)T��Q���+C�Ӿ� �r-ǖ[VW_d߀][ΜS�VQZ����cx7f�u�ܾ5��p��}+��v3��b1A�n���&Qc��j�Z��>>?�~������Gv�-:RV?J�уqǼù�x��`�d�Okum�'J�!�-���a��]�%�A�w�b��[bcۊ"���{��Ҝ���j�p�DW�>>� ��WI��}f�ӆa��^��"���]\6$�ZŪ�4> ���r���p���-�9/��-��pl-pÈA7v�(�dK9���h1���}n-(�e���\�t&�c�V����<��SlX���F�
��^y�}���^dC�y��3\��f񏩠V�f��A1��t�a�E����
JZ6'Ƭ�ct�CV�,��1Xl)[dA�3����i,H��BpK(I�`w��d���5ކ�ۣ��˞! �Q�z2�E;��m���#"s`"ཬ�m�ʕ�(XЊޮ����	����r#s�����9���1��r}��h���D���C]B�u�]�+xpո�Y����Kd�KY<������{�7�����*i�	ة��v)K,޺�<�j=ge B�f\��eC�a9C{��-Vѣ���ϰI�Z(��t4���!��>��ZNi��;��¦�rX��z����G���-`�o��"�ʌ�z�}�4�,����C�^�嵢�7J���*>g��hд\{��(/���d��ңJ���3Y���7���1�tKc��z�uRɅ�@Cj�^uE��m!4m_Lf:5���j����
�Ck7<�2�}�s�s~�����y8�=gg��U�:���x������Oh��N������>�RNJȊј��������[�P�b��6���)V���3�]�t!�xm�[�{s2"i�2�8Zj��w�;ާ��" @�Ȼ9�h[5o��N�S�6��S׵�q&�k�tD��={�����SQ�*hH���i�`���.7h�!t�|=3�K���e����9laөN�����4�`�՚RRc��JūG��6�JГx�}4(�mͫ��\)aQǵ�nK"�r�7��U�-�4������է�!z��Vv�/�ǹ-�Ƈgg+�msGXڰ��bA�w/s�ӯ���ED_!>Q�o ��9Q�H�]wt(�Ѽ���[ʱ�kcMk[�5��o]��`��*�����zLu�H��Ҽ�>T�xeYsxG�Ee��w\�N3���}��Aۂ�L������; �]��u�1�ר��b��b�A����\�2
7C���^��{W\�q),Z�o"�tM؝�n�Y=M��ݴ�\���޷e֞z��e��e��+�e��%Vdo���Z�������(Ԃ��Ī�-�i�GcJ>+v)m��ÄRX��"`X���b˯��k��ѐ�M䤵�J�CУhj̄�(��<��1#��}���~z�i���=*׷Ӳ�ԍ9�6,�q�\����cj�R
=��@)�78:_'RYF���Yq�{�,�z�1�,ooͧӝ⹮�ճI@�Ē�©��4���5V�]���wZ#u#1�*��nJeˣD 1�]l��wB��5[ai'�W������-��3�4�Q�%LYJ�m��s���Z����G�n<��-+:S���>�Es��a�5�<f�p?e�U��x���������MeQۺ;�-P6�L��M]F������ʍ�=�;���:DDH�C�ʵ�Qk)��;�����I"氉X����ua�x�ڍ��,�'r�.���!Y�f�̧�ӗ��*I��4w[Ʊ������)�X�~cceZƚvͫ*��cp@��Mے�e�U�����p�9�5�ܩ:�X�ā�B���6g.6��Y�f�����O���,���)�&����2�xES�Y�����
6	��KC!��,`[ć��V7s��۸���ť���>�P�+�%ƾ����Ψm�7V���ASۍ^k'���9�yr��i
=m�׋���B���Z�b+�(�T�i`f�{���28��]ۘQc�B�ԃ5���R_b�ۻWem�&�1�"�C	f��i����,�ƎڝL�}���� ���V���6��l�g�L��m�8%��bC��k+.U�Av;�S*��f���׀A�P������>�R�T�HV�
���z�-�\)����üH$bz��:��!�w��`/� �m^�Zn���O
�}�[�@�[��+��'X�}s9iMB��]��(1�)&�TN�aU0�p�KJe���a��Vu��wk۠[|C�uŷv�wCo� �2ʱ���k<���MLtLZD�-[�۽G����1�aڛ�;4����H�65֜� ��GJ��.�s�H�����}�`�z�iFWrw����Q��gW$�ۧ��;�z���!�ݘ1�XsnƎ<f��(�	��10X�7:�&E�������Wn�&���Y����7��;��Szy]�ϓ����lCc���B+Q����M��oy�+:����8hgZI�看|���]�] i�رA�y��]��c��嚱44��v]a�v�d���/p��X��T�9p�y�̝�L 	�}���(�zI�aUw7
�\�FD�YT��O(��fu��,!��0��ه[�@���F�5�:�A3�"p��Z�Zj#gq���G�Z���J�p^�'^�\4��B *��N#����c�T���)u���m�4q��pә���Ϧ�����r�����r��w˒�:�{��S��IW��1�8��Bb35�*�d6K�q��0��b�XkNZ��(���Q$y���ʕЬҽ�l]�����;��c
ޝ�@/]K#���ɹ���O�=�9cBu���vO}O�Ow�T����ڣ���T}�ٮ�A�j�;�����!�|�8�L�;a�DT-6�>Dpv��7.d����&��m:V�j�]�\����zJd�Kz��a�x�=��9Fk�w,���
զ�s<Z{AI�|7�:�΋��^#I���f]����۪q͵���B��y�E>���7s�b{�Zý�A�7����ٺo��v�k�HX�)���(�\��vW#,da�=�t
<�\W�d���n�7�Q�(�f�j��o=�vƌ�� �\Â��l4S��Z��&��ߩ��ZP����C��pp�U���ӓ����#[�����,��:8��9�;��g�םRl7*�%y�][��͑��n���,J�*��nno,�NԽm^Aq�2�yjn�pǢ���u�����ݚ��#�|�0��~� ���E��Z��A�T���Nxe����m��I��a�|�[��+%Դ��Ӯm�־�F���//gYC���Y�y %s�ܺ�N����a�}�s4�'��p�T$��34%ږZ��OX�1vsiL��F��,%)���c�14=�a�K~����'��6°N\�.�n`5`#ȋ���Z���ɰ��a�Z��M�IBXw$n�LWʺ5/:i����z���� ߛ{6����L����ң�V���o~�l��Ө�hV{�H��2�F���xx{���n<�%\:�tO�sBwE����`[s^��.��g�w�{ �N�����x&��b[���%LZ�����[�EG�̾fu�O0�7PZU�j&�'>=�ް�9s~(�=Nmx��K���3�^:�Z���h���Pd
ٽ�V��'c���J�GM�P�1�]�n���5&NH���y�d���}��v���S���#�Շ3!n����t���;����Fɭ���-E�u�_�R��o6Wkr�ϭ�t5`��h��K�%�����C!��S�>�7�On
	���)��-7��Y�7���'ӷx�e�LzY7�;�׌�r|���DZj��z��ٍN�pܽHa&�H���wmH�06�y�WT�wZ��3���T����j٦�KV�Z�Sv�EQft�᣷��7�����u۠eٽ�^Q۷m#�*�%������[�i'���h殣[�x6��F��4ʭ����\�3�;<�e�|u�}����I��4���6��Ч{ =M��O)���5��kX�����v:!<w�R�X32w+��`����W\y6[w/�R�qM:�ژ��s��ߖ���}T�a4*�¸֧m�8���-�\/J�[bL鈞���xbkC�Z�t�}�WY��rw��g����킚�Ϻ�sɡ�s^lr�	x��x@�ηVb]R�(����W�H]���  e�)��EE�6��r�r��-�X�+���U����E�F�KR֎e�)kl�-�PT[J�kUjTcJ\�%K��Z�U�*UE3�c�Xfa�V��1ģb���U��b+m1��Z��cr�q�b��.fbbS��sJ�R�m�ۙqR�
��\ȍJʫF����"��e�b���[(���m��e��m���TpJ�T��j\���Q�R�h��Ƶ����\[j[V���,�\L�W)��ԦVcEkpiZ��l��U.����A\�X���Җ�[��U\�*R�cSH�8�c��Q�3(Xe�l�[aUƌ1�[D�m-�UeV����Qb�T���U�
"���m��R�EU���*�˂Z�,4lS2̶��\\*V�\K�RѸ�����QU�TˎKm�L��Kj\he�)Z�(5*ێbT����������h��o(��Y��c������v�����9˲]�{�.%H�GGAȄ>�gIX�����g�|�:�\��9~��k�3���W%_+jl;������ώ ����{��`X��l)������t��*����]���Һ�OP��J9[$�V4�&e&��^h��
;�Lj�b���.�N������f���ug"p�I�������|�������U!�(���W��#+'�vdC��k+:mh��\��6�dj��Ǵ71=���<���M�v.iT�^��N�^�n�З��O��^���%vb��}O��h�H��G��o&��u*�Tؿ5�Sn%��mr'�뻝ZY �[!y�Y��u'�����-�f�uy�*[��e��\m���<i5��ۭ�Ro�N�d�q�[��A�9�jK���ӥ�q��HM�Չc}Kw^�ܞ�`� F:V'&}R��8�)C�˭3�y�o(���2�،^��2�zv�E���T*[Gu�EqAe�U�t�L{�6����c�qQ�㴅�C��f�n�7�
�Ǿ���;{�,�����/kނ�j2z�ZV�e����v�ݬ�r%u40��]5�/������*n�n]�OV�>����ϸJ9��yWRC�*	.�T2e�r��0݃��n�t�9כ�t,ӠH�x]Q9Wy*1s�j�n3Es[}*+6����^M�~V;q��؍�O��a��ޕ$��q�UK�حj*���}mX��� ����R�k�]��_cq�`�8h�]Be�����]M��WI�vP�E}J�48�eg�0�<�z��\�S��y�a*�ن���!UhѪp�7r��h�W��j�[��9��������J`>T&w;���{�z�P�V�#V"����Ϭ���|�C��o��F=���&AZv�����B��\��ۜi��f��{a�5T!��v�7A�˙{ok���\7>��̟D�u�B�V��]��x�v�J�nL��:;��)�p�����5��ՁSl]�@��9|�g#�����P���ek�ČCMw�'d��f�fԥ�@F����f�|����*ުS�Ӛ��&���{�Wn�FS	N��6��UzqWU��m�����si���j�"�f�՗4C$d�v R�*[���ٝ�<QWV���Z��Mߚgfs�w�l�QPf:��'@�1��M �dk���b9��y7���k�K{���Π��W���ʌ�JРQ/+��5[�o�Ȱ܁��/kt��P��!t\�U�Y<�g���aо�V��}K*���&��'�N�P�p�mfnO!O����%̊�c����0�ۧa���z����M^uw�S�����S��s��p�N)���PIx��6����8ś�-��|L}��R��	�0$vO	s(P�ʯ�+ؖ���>4�)R�DcWd�.��0/q��x������R�R�Z�h��ݛ�:p��U��<l;�ǹ�t4z�V��;!_��ᣦ}R�RF�̩��K۩��t2q�fBɆ7�\��}m��l�=��S
��|�}$�w,u磬�'xS��I��k�,���.	�q�ͬ�m�2��}�|����-{w���-�LT�TͲ��o	�Ï�ܖRع\��SX:�*��N=
�l���L�{"�kv��v�ZVk�V�
�f�4=%p�����=o	j�}���YUܰkԞ+jl}ʬ;�'�S�sILr�4Sm�^;��9�k���I`�S�W�:J�S�^�����gf��{'b]����
1�7�@��H��b�_;�z�������xMN7F$c���bN�
�}�Gt5b'q\��'»[H)o`�f�	rC͉�<��Z'�M��<�:�/���ļW鼟^7;\�n��MF��:nnVwW:�)�ի�BX�џ&�; ���k������"&���j��n�<8�%�6��[y��_�i�mk��<��ƫb�:���I���c��i>�K��{����f�����þ�7ͬ���V��&p���r�҂5�3�����G)w�[��řU��^r^sۗ�KY��d�N�y�Q'�{n�&�xc��%Lc�~��Gs���WN��
4D�.���˃P�A�y@7�E�;��
�3�O�L������a���,͋ήvb�cf	�c��$5�On�y���7��9Ox�6XB�������*zM��m6d�C��OK{�$��c=@�X3Rڨ��GY����70f�CrqOo!tg�T�y�,���:%FltE�m*�h��U�W��֦9�$�|��@���]
nq�XE�t͹��Q�������ֺ��CƫZ]Bi4S緻Ntt��U͙��j�pϸ˄�Ȯz�"�:�q�9���:bxN�1�6 ڎe_��҆��t�#T#&��_T%��*��n s���NKRn^i�޼R��>-IjcB�SE�}b���󿩚~�+:��Xn-F�'��[��&���@���T�ь�Z�>�C ��,���4pGOu@j5!qW�b랚V[�6=X��Ff��Ya?G���2�# w�(�0z�L�5����A�ڷ��i,������Ga�r���5BZ�=�փ�,� !��* �j��U���fJv.��]�c�C�}�啝��[�K7����(\3��Er�3B=��̹Z�/����%�	�y�;��iSE_u
~į��5;�a�y;��	�H�Y�����Hᶒ��s�ɓg��ܶ+�40��`jB�^u���9�--����*=��������E�2P�Oa��m��q��l��<h�h�l���9lh��GD\�M�ojF�{���y4X�^�.���;;�죝�����WS��f���N�劳�������oH����F�f`vB��9C'
2k׏�9U�����ŷLɯ=B��R�1��%�M�QU�,t��Ip&�HfAÅ������6)�5c6�)����C�&ko4�V3;��4�9�'(}s����J�afEջ��U ���)��tR��)]r�c�$��eYX�/�,�{7���*���2�	���zVf⋱�}q��-6`v̝��:/�K��7��o4��0�{"5xd�'ֶe�e'\��3��ڃ\�ӛ���?L*�K+���#f�,	׭۠�
s�cO%:g�׌�l�yW��T;X��K��Dm�`�+v��`K�o�V���nQ��CQ��ft^;1�׼��I�"T�6}" ��!	���t �@N'���<�]��U&s'qx%�k-�fI�O���w�2#����L	q	H���I��(q��;�+��YYȜ7�覝qe�A�ieJ(�ǂ<;��D0R�T+�s��ʻ�����Q$��c'n/���X't$�H�13�'<�p̗W{��{{�-x^zD4]7|�n��\'2[8���w���K��C���������.��|��z2��f��W}���$wF0� a9����S������:��>,z��p��w��^<�rs��r+"JQ �B�*}2\qDV�	�6���K���&�ߋtȿj��}�E����p�n=�����@B��{=�,psX54�)��F�|�6��;�ưҜG���K����.Z�.2�0!��ql�����٨��޸c��!�L�Ԍ.� �մ̚�ܴpt�;�iE���=�zB��U���ѓ87N�0�
E���)_��%�B����O��Unw\.ӧx�o�ց�I@�t�~	O��SW��f�+���'H���n3�D��)Y�M��c�A��7���@;psE���a�0t<��)��DK�@U}x�{�}��n�	l^bm�/Bz�+�U�ږFX�v����$�dw�
Y4l�B�O�g-D��[:��ֽ�in�z$�.r�r�M\���`�˥���W6�^�k�{rс�.�%�M����)7��J���p�T�U�4�9�>EX;4�ct͸ڣ3!�>u�a�T��������ar)zz�4�qc�}+O7R���(7���W)l=h_)p�%��|�n�sG$�sB���w�B;v��ï%�SLG��=��v[I���N��N���5Ѯ
�:��(f:�+����,*bZ��i}7k)l��.s���Z`��D?>��+=>� Hs��E8�0$�x��ҭ�d1�揌���pV�F�"�{�B�/V�P7���W%�B=�#Hɑ-���P@���k]�����]ox�o�fYjצn�y���e�+}Pu�d<�<rT��3�$���P�`�A��!��Z
-rS�lY��6�1d�~l�*ƺq������¿�#����9'+��y֞̰ J���W�z��͋p���{�^<��8؄x=U��&J�ʃ�[l�t�7|��>�XPGB5��u	�l��T�Wpr�m���J,�9��͑њΗ7Ƶ�@���o�$����-:$$�������*�I"=Y(����F6�PJ�x�8��T���)Aެ��`�ӬN��.l���;\��
��7�M��P�!=��A�[y9/o��cv��>������~N��'�A�<��Y��mVR�-ろ�&���oX�^�˷)���U?m_E^�g`q�,&��(l<0$������u��p��a��6z�Y�f/�	��[b���Rj�ˋNJGG�^���͹[p\ ��7h�x�# =�/��&�a�!��|Ts;��jr(7�8�n�J�ݷ�l��0N=Բd�
�ƺ�s;%7h�e������]2y!~���z��������R�9M�|*1Fnϲ��dR�mAƺ��e�/&�2ᨭ��h�b�h��u��
�O5S���H�dÃ��deGh���gk��7���X-��҅���{g��h�!����7ۮ�l�yMP���8d�T��J��t�9��2�j�[�m��1�BT��4�/-��;������ti�{k�"$pr2�zQ6|���C�K�E���5;��S3��VQ״�s�I����~t�Ϋ����OB��DM�O	ψɆ��z��l���'��pw�;}j�[��Kz�1MN4����6<�B�G�l�b�15Si�ٗ�U{��y����4�((	�U�=J��YåP�4�/�zmC#�N�-_��E_�R8��aY�0Sѷ�8��goۛ�s�уԺ���U>�b�k�dׯ�_TbS�z�U��@���<�7������OM���|`9!B4&Q�^L�}5�����f��egC�}a��2ٸ"����ƃ�_gɂfO��NĚq�D�2T�DBG�tn�:>| �V�9W�����#�A�}�(n�E�Y�[�wsΏ;GL/g[�K2w]�Λ!�̍��4(^{OW����M}6q^��2ܱ9�J����_e��܃�c)�HvR��#u'�͜7�m�Τ^a�%k3�+��g��ܿz%2zf���f$N��(��V�~o��G��(f��{�(Ƀ��L�X�R.�T��ތ��'\���YX#��a���,�U�j��7Z��!���T����k&��x1�_z>��x&�����=щI"�-p�o���W��2�s�"�M��!��{8eRpѺ�2g��R��Q~J���ثn�!�^U�N�6Rj�S� p�3q*�7o�Г׳U��o��uRЇ�U�	��F��j�*���y�ʭǭ�����fL��΋�-\�w��}]�0�\�eci���q�8[��a��W�L�f�m0Saqx���$<Y�0�seQ����[}zn�\ҟ*d�Q�������*�ࣞ�fVU�*��L�q�~��j.�Oh��Ë�+Ct4�}!lny�fĚȨ���n��.#on8޸�9��7��W���R\^L�Q�.�Nn���>���y����(K8���RjpD��w%��ta��&���ʡ}4�Ȃ�n,F�8Y���܆�w��XӃ��9ξ�b���zB��CE���
��sr��-SsYa��6|3�n�'Y���7�owqc�Ǿ;
�6 J׌#ڲ�ܴ���לm#���_|%�n[dk#���\�9f$N/������\�>�wʛ��}&�,��u��ǜ�õ��ޖ�aP�˺ֲu�sV:`�׍*uXhw�ơ=���aٽ��׃;�w���s�S&	��_o��>P\S�g?���E��PÛ�j�S��De^;J+@B�W=!����5w�q�.g�Ƙǯq� ����N쾙����{n�~���o���m�(Tٛ\(;���Un����4�>DI��5��lta���ZCE��h�խ��5�ږ��BXo��2$�}� ����k�2�zw^�b3
W����t)U��P2з����8:Ԭu���Ik�C�4z��n)���;� g;��`s�x`��L�s���Vv���᳕��GfZ�帗_�L�Q��M�T�;-Ș+��9�~Q4�x�3�f�����y��k-�t�K�S� ;�J���6H����Vi3��	���,5�MW)f٨��Wm���os������S\�;��Ƴ��\�*ͷ��*i��,D�6��֛�*��0�WJ!Jh}�zK�
.8�D˻��-W��Ն��C�_wk;�wd��i��l����la�N��Zɨ��yn�����\%�M��|=����	1]I���8]�;V�u��m}���\�=��@Lv�˚w{�̂�6������C/#���Z]��7kJ��|1�
��Ƀ�3�N�
&���ʇ9Z�dm:#M,�G�j�1JǄ����	f}g]Mps��*�AS�j8mG��+
+:�����ݻ�����ˠ]-"i��Zk���'k6�l͑��l3GW,�(�M*�9]�[��k ͮC�N2WJr��nnV�#�t*cx%�i��s2$��R�״H�n��AeGei=���ew����u���������P�ʟ*�Uq_�REj5���@]n���9���>�0�u�~;ټ���G�f�r�6"�:sWs�����C�P����'*C��O���0yc�/����=��V�{���IԈ����3t���z�|�m��[En��J	�[j
y���n�Us�Ϩ#�Ni�^s�L�i:��N�l@��W��t)��&>�dw�ho�����7�Q�_o�*|D9R�ԗ
��n�X4�L�c6����$�3�)_Y�V1̹f�r���t�C(�e\��
�zn�Vm� ����t����ܺ����&v�ɹuY��\#)���JH��M�(�:ߒ����N���6��n�,�۷I�,�dޘq,����wOP��ٽ��SU����Djޱ������,�>L�=�KB	�j��E�qӉHC�ݜj��_�6Ɩ�X��֖��kX�j�em������F�-j"�jQQTdTb�ʪ�-ڭ�Z���Am�P\���ZZ���IX�R(�6�����T��B�(���JTh�ֲ��ZTX�+i[jԌ�m�Q��$��-��XV*�kR#iU�5�,R�
֪�
�Tc-h�ED*[ZUKAH)jV������R��d�,�EZ�cV�#ikF�B��KADB�R����D��1�kTQ�Ae��m(�Q�FЭPU
-��H�Eb"1�Z �TETU���
!h��F���jb�T�D��#mTh�J�b�`��5+R�k)Z�m�e��U�Q-����A[h�l���m����*��UU���PA-h6��jT��ʕ-��ȣiUT��U���*��V�U**����ѭ�O��
��]\��uv>i��f�;2�V�b��m{������Eoyrλ��C�E���ky�Q·�s�Ն�q��ܡT����%F���69jQ�����/L	p�>4-_��|����n5xc)wǤ��|o��:�)���i��q�ꐄڮ0k�΄���K�UDf��Vtt�h$,�eC��m��88 ;�H�z(	�
50%�)P�����~GLE��D|���o�f�Ҹʩ�tSN�E�A��R����G�Y���+��^=fX�Uf'q/���ތ�8�Iu��[����v9�&�S �B�*����u9S��f�
M���zQQ��'�3�Pޞ!�S��EӪ���dy7U�b�r ^�[=}aV�h-��C�M܀�}�y�K^���=VE��\��+�k(����i��;�d�3ӷ��Y��WȬcY]H��² q[Lɡ}�h�%˔I4�\C�0*��d�U�)Q;�w�)���.�Κ.���e+��~5�(,1~���K�8�a ݤ�*�g���x�����My9���^D߶Y����U ���Cq&�C�._B��R��DDi�W������$��l�K/ˠ�7���.0/r�gq��MY�d`�3��>R��}t���U�(�h�7�io:�S�}�m��w�vY�J����E�>�>�s���.�\�{܋a��فg4g���<�l-ـ=o-43/4���-���4XQ�m0FW�=����Z�*��n�{�W��aZ��wβl���74vu�$��᜺%D��*g�%�޿`����D�l��̉r�kQ��BSy�����3��Y<���ҫeY]C�{W�zB"Swh��z�z7Gѱ����0��oLB��^�Հ�!��ex�����k<�e3�U��Ӈ�n��Ϊ�n
aP�|5�Wd��U�0Ԯ�Y>� Hs���0$�@K�!^t�G �d2a�_U�4lv��[����z���ۯ	@ޫ�|��B�q�W°U�T��6|�u�N_)[�9��\�Y���⫤��;����6B/�yv5pz�t�D9*I�8H0,���a��ӱ������.���U�(��Q�d�a�(��N W��1^]51����V"�uf�;��Vh~�����R��\ξP4ӄBw=Я�h';��7P��
�q�]�QY}��C�e�:8�,�ޙ�ȆY���Ws�+n7��Qf���qln�=$��wb1oo��q���V�''c��*�Sky���;cn�[\F���j$��f�c"gkY�O\�x�nmI�o�o�T�\����s����	 ߥNj;h
���>�4�b��M^\���t�����¹�w)���������	os� �$�����@�����N�Z*I���g�xg�䣞������9��s�ɳh�SD#.Z��6WJ0�R
�ixR%a��n������wj��Nź�U��}�y��M(��t�(�U@,�h������H^8(�T}4�9�uE�����ҩ�=v+6E8���q�=%�M\	��&ȭs��gJ,���l�Z�]w��e���Q&�/2}���{�mA��Xb�!�D��֛���jL��4x'�M��2M����$��Pr�NN\,�
��cNm:�e��έ([t���t����u۸�0{6x����ժ>G�7遆���W������� <�:w8:��,+y�yD�8R�[���{l����M�?.&σ�_���F�hӵ<�����w-1̃�2-�,����çl߃�W���ΉQ�c�&�{8@F�#&�#]��Kbs�r6xSNic`K���
jq�XE�tˈ
�91�c���������.ʺ�(�2�kX|l�Z���TW��2U�{l��뎠= �7���!��r��ԏ3'u���@��F���Ӹ�q�Rp)�?�Mr�5;45L�_����*���;_�q�=�os�Ɏ�0{´_�
��p�^ޣz%�鍬wo��]��
 ��E���Jb���204�^�B��]�S�F�s�an3e�i��Į.��q6�)QAQ�ģ���.�@�R�P�p��֯�0%8�|�����i|ru���DH��ӽ�s:em�
�B|cd�`���$���G�+y�8?<�٬�+:�ͼ�d��*�M67��|���A��Y^�8�ߏ
D��e���d�qGda�91�֊��%���U�XyZU���<�5��
�e�ߏq i�haj�X켩���ϪuVq��\�R8,��\'�������5R���n�!�/�C1>�<VM�o>���J��9�e�����φ����RH����,�`ߪ�2�C7pDW)��w�ޑ	���7ө��T����#^��¦Ɓx����^U�vj��	�DW���dF���-�����ޖ�\W��tӮ���*�H׬�5W�p�&�x�`��*���K�����ǾS��F뾭�t�=��x̀������D���W�8p�u^�7���Lo��g{�ɵ�����6��9�w�*��F$_��/U����K'���}���9���X��Ű�+��M�,Pː@���\3q#`�2:k�؀p7�9F�k�/�2o	�D����/�/�ZQ�~`Z��z���ʹw�-8�瀌�RoL��y�U�.��*��A��؟�^�4�>�P�YG�WK�-�*�����CSx;�`���?b���lq8�}�eg�����]�.����J��yI�e�9�c3s	�����ځe��QFS��c&P(��S��Cp)ߝ��i�<q�����E���ޙ}��[�
������H��`�U_M2�,��K�~N�nà�
s�cJt���N�uK����T�y���U����5�C�J�x5��8�B�B0kح�/A�.��jj{�p��=N`]��1��(�3�Fڮ0]a�=^:�u]Nzs|�5Wx�F�A;�i+X����0t�P��M8��a�xE� ;06"@�z �QɁ.˹�YoJ���Sb��J�����4_���3~w^}ܢ�ȃ�=��6��|�{��ze���=�1m	��Q6�[�"��s���75N8o����Ǘ��v�7ty)�d!�m�h�<��曾�]��s��ў�!��O�����P��Q�6�jQN���9����GL�RnWG�l�y�� << {5�3c+�B��0�jȌ��Ϳ x&��VF�s@v��rX��mK%��/E�K�On�y��=\6#g\�3��u�0��Ө��VG��fźF�!b��v���Np�KkGLű��T�B3X�3�5��@;P���ة�
�Ҁ��A�x�hiU-p��5��K���p��;�Gp�qWW��A��a�+�]V��_kh�����Uc��[,ɻ��G:	t�e�Y�Ĝ�ѩ�I�9�2B��.p�΅LPB=24N(��p���^�2�6ln��*��s�te�[���K�U�N}�h5W�66Y��琝"G�3!���U	j�>q����1���uŨ3f�
1��Źfʞ"�5^؉訋!�QH�4ʩ]�+4�g��őbc:.c��λn
��<X.�|�>�N�>�֘��tB�&����~��{�/�QB��xz��NV��?Xy�g�u0^C"[���ZX�od�Sk��#%Fb�n�	��1>%G�`�Q^��p�T�U�4�=�R;4�P'[���3{VLVM���2�Q�jE8�Hn��i�p���0$�B]q
�Z$�٤lO5��Z)���j�
=ɾ�6��t͘ΜQ�g�$�Q��2}"[��!P����Z�r�V��z���6㽒�G 9�LIs��>ͩ����U�b�|+��O����8�6��o����w>'C7�_3��C�=]뱐t�=�g���ͼ2kb��0/�vK��#��DǼ635�z�Ͳ�-c�Y�����%��&)���Sd"�Ǘj���K!�A㒦�4�����;��x=j���b�7ʄU�(��j:�\[���(�r�=�7P�L¸:�S�d�����[4��z�@��C�����\�a�B�ݎ�X�A9؄B�V�CЗ�w����U`I� h�g��hH�B�L�K,͍��(��ۍ�Qg1u�2c��%:�֢!��zl����ߓ�|��%(���UԒ#Ւ��},�֐et�^�X;1�Q���:e��j�w�����F�
DO	d��@��S�i�{�O%H�0Z{Z�<��ӷ�M(�n��"6]�  k�������Y���)=�z�V�w���ƧG�b����u��fп��T�8�zKW�����h��>���Iv$nmI�W\��8�Y���SQ&�77k�c5�DU�۶��]a��#^Mt""C�h���x�	�����Z�+L���A�F22�mNYڰq��vRo���+G�^�\�%N�i�=��>�g):}�톐p�1Znt�R��X��l���,�w�&�ٛV��*��e����
�e V�9i]݋U=w6�=Y����17�1����`����^y{:r0�0w���j4B�fo�.��Z��yօ����Ղ��Z�����ǩΑ~f�&�u�|���xL4�Ua��vΝ�%��ܸ�\�[C/b�{�!uS��A�}�����@�Yc/H��
W���-xO[!�˱��s�/*�_f�5�1��·�U�E�u�n��nu^�noJ�ՇIN�־�U�f�������~�Ա�[����OPW�i�~������N��t�d,�p=[1��<b�^�qN�y���S�>b�RU���}�3��3�2���B�밊�:�s�ep��,��ԛ�������)X�g�O��:hJʿT�J���p������Jq��G�q��uk v��H��Q��B�_�NVg�=�C�4�
:�h�!O�y�9�ϭ�[�V����~�NooVg2p�tu��'p��<�htuD� �P'��DLAp�ȝ�t������NI��fN�s��8o�j�a�E\S�ғݰ�q��"��G�R��=�u� B�s]J�uټ��X9���3ڌ�}R���5U���h0h��D&;&�]w^��X.�L��p���ѨQ%j���`���s�=VW2ۻ�p=D�zz��[�����[Xzm�iͧavT�m�/��K�pg]��ŭ��]������}�=��tw4����DOrdf�yǢ���5�Le,Ū��wF��/z5�s�ڇu�ӟ�;���b���;���@S�;ixM���BC!��8"5���B���v:��-Om�5[���|G����haB�x���^�a���<�'u���ꪌ���e[9t�Hɚ�p��Y���"g
f�0�"`<�u6s#
2v���|��z�=�D��]��\�Y�(5�̚P��n+"w��6��T8HFA×�f|�Qk��<R�Թ&��oϏ�Z��M:`���t�Oo�M�꾉�T.
�?Z�����|َ�{��{�¿]'��^y/j����Tx�;�+<�/�,����bM_�n"G#N��o{��6(�ĻZ��q#291��t��2�F�]"�<��S���O�i��) I8M� �����r��a0�bl�)4�P�N�*���+A`�4�bu�nCp��j�Fj�9�b��������ʸ�ͯ�����嚝�r�����V��-8�+�V��I�L��E�b���G��6�s<Dj�0dd{`B:`!����t ��owf�Z���x�3I$6l�bW�0 ��~U6�Z�*��3N�'3��J��p���S@��P]�t�B�=u}�I�A�oG��:4E�H��,>��2l;�4�ƶ�Ү�+���ܶg��y�K�v+�Z��A��ً�w,��*�2l^E|u��k���C��xE��y�06#����0�F���j;B^eYN;��@�B=�cP�6ןE7(�b=�u;����#�g��]J��:����;]�V�۵�a�6x'؜	6�qW�����:݄�Mĝ)�u-6���3��{r�҅�|4�	:6|���g�H7υO����7�\*U�w�ؗ[��%�ᱛwg]��ƚ�7����"�%�PHF���u��"�Q�1���Mˤ��}ϬjOMN2WSi�����:�ˌ������D�������2h_nZ,��׷t]��&�<�8���B�7�,rM(��)�XXq`��S�zgD�2�,	Aa�k�c;�sY�v�����-���ڷ���<�,	��Iϰ�SW���p��R�bx	���Um�u}�9f
���0��zs�\[�y�E���bܳ�OY��5�L�=g��mû=�������QS�d\�8��de�:�*4,^��R��l[�J���q�
F�غ�J<��P�ȼ��e��fR{J թ�xs�ƞ�c/lԽ2oN�u�`pdW��p�,�u6�	�ol!�{�y�=8��6�[϶�v�9�� .b��)���
�,�)�H�߀q�%ng�o�d~���:��pP;.����3�k[�CLwM-] ���$vGc�}�8�N;�Nr
���liv�:7�[�uxq���znx�gM����d���Ky�ɠAa�zec��8�z������Cg��V��WE���<���Hr��'u0��g;ùh�*2�´��Lb��y K��F>�q�F�^�*gv-(� �H� ��)�<μ\6�^��0I���hL�֋޲�[F�ʶ4j��xJ�k�Q�rw�ʅ�^pwy���ri��~j���H�2?Z�k�oQ�%ق"d�A�C�m�����#�2E�ewf+a��nD?���f4�/gu2$�G̾~˝�50K|��c�r�v�ȕ���L�ؓL؂�������a�Q�8r]���|;'84I����>�qO�@��뮲i2��j�0���07�j�ZM�@�r��g��r3)�j�|m5��C�n��v�f�H��9����9s�sӜ���]U��K4�dZ�PG��@~m=�{[
Rcu9�����h<��W8)R��2�ܐ��f|Fح���47)j��G�.O��L��
��oa=�*��nE�
�jX��gk��q�`mf��]A�ۭM�%�58up���r�9e�O�ˇe�0�}��;]ʫ
	t9Z����X:��Q�Z���X/��Vnu�xf9��˵��]!��J{��I�<��p�6v�r�ಏ_�	o�]e�I�ּz��yj�l�v���+7�Y~�i1,�$�v� a�hT��4ڬ���U��D[�؍�
������ᕡ�YF�#j㷕�Pf$;SR]eA�|䦷��--�'TA5�0�Ӹ���6�����4����Yl􋤾��0��IO:@������-��x�5��8�#�2@��bȃ��f�h�P�oQ����qO���O����2�YOIû+L����b�;�]�mJ<�i �ؘ��[�go:��i��)uմ��Cqp��<S�����"�>�;l)�ļ}�Tf�rd����a�o8i���㮅��Cڳ�8�#�!c��k����wCu����5��Y����Vj)�Z� mY�� 3��Ny�eڷ���ᣎ�"��X}0E�~ڰvw"��S{�����>�<�U7,e�F�4�8����隦�v����q�u0ui.+4u�n�)I�8�T�<-=7݈05|��:@C
6v�P�C�ʘ���X{��@oV��݆p�<�c�U�A��巤tC�Kl�FU�: �������&��m�c��.E�{4ǚ�s��}�SqԺ�e� �cTދx���ޭ2%;jU�0PD�QdS�T�
���֣d�D(1���
��KlT���F��R����ȶ� ���VQKQ�
��E��X���Am*�m���,��Tm�
�jR���Zт�b��)R,[iX���m*DDb#YD@�[KYH�PAb���5�-eAX"��**�Z[aY,J+-��E�Z6�*%j�j
���,�J�Z�P�dXV�+"��V�R�Qi[+Um)JJ�d���5���Vʬ
T
֕m�����+b�J�����T�*�m
�!b�ʪ��E���EFZX��ڥ�dR"��YF�A��Ib"�TmJ���-��*YiX����1�a[iKEib��h$Qm���mATJ�UR��Q*

#3��{�{퉺6�b*�=~�q�Z�"��һ����;T����_.�yc����̸��
�#�d��V(���쥕�� j0�K]��5pg���>���փ:�ק+gq�Ul�����`��Ȧ�9Tn�q�v�O*<}�v�=�E���2�>�C83�η��*i�ptϑK-�[�+��w�g��_0h��g)�J�7"��#r�%`�i
�lM��Z4�S�y�o����K�����\�B��=:B\���ڋM�&�p��� t����vx���u˽KR�_�<O��=�}� ��Ѿ�D��!��{�Myg;����Ҥ9i����H
)�n���0*O��&ӌ���C��r0����4��c?2W�o_���5᫮w�~������
E�'r�N+*$��01�
�<�!��Af3s�}���
�sϳO�q�'�my偞Xu�"�{���8�3���6�1���!�J�v&����n����i�}޷߻��:!���5�d:[a��Gj�Ru
βoZ�T�B�M�I�u���!�R�3g������Ă��0�S�xw̓O��}$Fo�@aG�fݘ=v�({�w�|.wl�c@�+��!�y�&!���Xi�qXk�]$���떋'a�
��"�����&�4���dѝ½`T�Cg��{��^R���=a�):�LI߰�ˮ��u�����~���_^�g|�N%�h�Ax��5�>!R�<�p<O{�J���Si��4r鬕������Cީ2������i��R�<��Z�d�
)u�����s����_%��.�޳GO�����0@���>�zw�m�W�����H,�%t���E"����jʆ!��k��a��t}E�I���ΰ������1=C�s��w'�F�p�	��:��l��J�u(�e,��1#2[[|7�(q̼�Ԡ�Y{F\��@��uG|DcT�<�!�f��=�����Dr��b��@x�vv,L^��/z�n���)�����M� ��⺞hs��+��ӗ�m�6E�B�<��,����=;�����G�l4���l*%C��{�m�q�=�b�I]�����T+4�������aX[g��B��=/p����t��$�4�6}E�r���';�ҫ�s5���W��� �a��;5Lf�|���T_&�|I�1=�CivO���E�'Xb��3i:�g��b{��(��
�Y�w��1
ɾw&�E��:�ۆ�A��A��Kyy����۞�ݐ���ɴ���i���nr������+����t�N�3ٻ&3ԟ�I����E ��=���� ������ya�S���� ���� �}� �H����kkj�]�$`ˣ��&>��N�� ז|ɭXx�
����?X�d�
k�²z��f3�1=dۜ���0��zɰ�����Ag̕���jN�E"�=�d�O|I�>#j������]�h�ߘ�?�R��?s6�0���_%����g�<9�	��?0��|�ͤ,1TY�ԩ�Rc��&0٫1=I]��vm'�Vm�a��}���>��V����m��~��~��
�Y�wh
�N&��oX'�돦����HT<;��O|ϓ~��
�~LCHWƤԘ�OC�)�4�}�X�f'c'���(�|@���=쐴��r͉2���?s��h��(���t��ZԜq'P�<�Yr�'a�=�0��^�T|���d����:�z��>�h9��/�ӽ�l=a�Ri8��?Xϒc��H�	���
����^e-���f����Y��ρ:@��> � 4�����M�	��Ag=�Z&�2TY<?fE�:������wgY9�w�u��<JÇw����%@�օ8�����'��s��z:7�޴�s0|�NLf��S!��|0�A���\�~a�T�Y?e��� i'U����B���kA�q��O�f��8�3�*)�`�a��y;�T6�|��y��<E�aP8����r~X66�S��6�rSo�i����I�EW>�жI�
�a�9�V�W�VN��N�Y��@URa�`i���l���0��B�<��q<a�6���9��=a��:��<߸�
͈�Ѣ�H�6�}T}�*��^5x��
��/�¶ǲo��+�"R��W�
�9��V�/�G��Hm���"_,��9�ѝ��%M:;����Kq��l~��!ݙ�4jw�o���(u�;�X�w��²֎[�{� ,�]5��cO�BA$�?�?g�u1H<���!�,�8�Vq1'�Vk�?�I�a��eVN���+7�&r�'a��1I^�z�8�R���Ru<z�A�n�-";��s_ς���q�&]�s�a�r����;�$u'\|9��T����.�����9@�cr��T�LH)�>��ǌ
�S,1��LxÏ���Aݟ�3�ެ8�gK�Q�
���wxa����O�	�~�q������|ɷNÞa'�>f����I�~a��d=�S�����O�L?UY>a�����}��j�f-�����A� I��{��0������,�d4�: |~㆐�%z�2g�y�C�+�)��T�B�L�]���
��zw�m�6���N�V�n��w��������Ѭ���<�tP����ÙL>a~�1��&0��&&�++�!����H.$ѿߵ<C��1!��4�JśO�1<}�SI:�g�Sӽ�x�Xm���+�d�ĝBݏ9���s��_wn�W�X�� �zL�}���DҺa�(��̕'�cY>Lz��0�j��/(~7I��������Af�~��׉=B�o�Y:��
�;�&�i�;������w<w�>������i{>O�bbC�ϵ��I_�
ǶJ�6�!��H:�L?#�0�J���2Vc%N�z������!S�O}��!Xi�y�u'����O��s1c/��2�>�j׫��t��b;�2i���8������K�B�����Cl��i�<;܆��?!��Y���a�T�uH:�Ϩ��,�
�g�P�%z�a��x�:��+�Q�R^��+෱��v|�gC��I���6�=����i8��6�Y+W}�C�m��P���<gό?0�Y=��&�xϓi�|��Ag�114~������ |G�	>�´���O2������va���+x����?!Y�7�w'�����Co��$�~3�*A�N��ϰ=a��Og{��,��Rnw�<d���@��ٴ���,�e�<��(�a�]rA廟�	�K'���>>�cr|ʁb�+*Y���Y6�ic#fQ�f�rq;���؉���mg,*���Hw9�F����w������������K�4�|���h�����|ʼRY1��7��~��Fp��BGp;��Xz��#Nm�
��x7wo���t��9�~�#H�'�@��.�m*)o?8�z�Ou@�hLa���4�'Ɉ{�4�*J񒧁ϵ��u&=K�:�$Y�p;�}�� y���i�ϙ+�?'����cW_wGײ~���F�zL�}��I�1�u�B���t�M��H)�W�&��w(���/�
���>֦��K�C�1�uP���%�@�i�C��l�)�g�y�����P"��Z5}��HG��V߇�ǈ��
�{̇h|��N3�@QB���4��$�
�j�'u�!P�j�a�#i6y�3��vy�����OyCl�a{C���9o{�^gf�y�{�x>="��1���-M$m�����P������q�S�c;����V,���')����+�n��&�Y��Xc�d�>�xH<���.�| bWW��uk���㊾֌�{�A>��A��`i�'S����6��;�N'�u��+��)�{�ĩ��ϓý���OR����d^�z��0��������'Ɍ=���qRW��}6ؕ
�_���t����J>D���?!���w��Rw�0�<=���[4��y�@QN�|�!���q
�O&w!�̤+�}��o=�4��r�8�]�k(�墑x��3M5E88�3�P�>��R��ē�@dz<�c1�
�q:M�,�>C���R�<���6�!�1�)�Xu�"�0�'|�>M��J�<���OP�7��m���Ĝg��,�'��!$%����5�֨�ﯹC� σ 	F���1�2VM��O�W���%g\a��y��m��l��M�x��~�*)��ğ3�~C��$�,��<M������W}k���.�eb�a[�zH
/y����i�<;N!���P�,]0�
���˦�TY�J�E�'S�ٺM$�}�M{�\�+7��u1 ���eI�%A>��W�+��#��g�`���O��)����;���a�T�Lg�;�i��J��E �f!�i�8�$���wvaP٪M$=�q�L��(�Y0����I�*S�DW�N2��� _G]������=�gd%/f���j�鷇�"WAA��9�e��=��aA�.�����+�O�9��2 �=0p��;�I!�|M ����ʺ\�uڝ�
��ud�R��t�v͘��]?~����K�t�W;�{�_@����I��Ͻn<��4��]�s)���@�Z������hz����{��U
�a����6�!��aQH.'��OP�����E�C5�~�߻}�gBU�]ڌԒ�a q@�=�����;��6��x�?s&��'s��9��aP:����!�c%a��ɥT��]$�w�6��z�0����a�i1���:�H,�{�=ٜ�tf;���������4��*(2��'�~N����%b�|���T����c<���٦a^�'}�!���O'u��Xc
ɩ�s���%E�I�y�@Q2bc�*c%��y鉋���}���dz�1��>���!Xm6r�T�'S�̟�~q'�Qg�VL}@�6y�k�T�����h�{a�Rq1~�+:�+��d6�Av�'���~C{����JחO7�#'�;��*�>~w$�6��f��H
)Xg�]=`T���R�k9�=5g�4���SL=7a���]�ny���AH�0<=�h�VT:��g��$���c�{�￯���������IR>g��xΰ��}��x���C��݇�1i��@�*�S릧Y1E5=��r��1=C�N�rO�vi������{'P��%Mkwǚ����ei�S�uY��>d=D�G���z>�i&��u��5�B��:�jÌ�i ���{�q<C����O|�CI��R�%b�5E:�H�C�P��l���T�Xi�x�����2���Tês�r��_}ܪ��dM�R����R|�ì*��`m6���Ρ���H
/Y8�w�5�
��9��l:�v���C��<O�8�g�>q&����!���_�G��K����U��������˕��O�s�J��wv�Y�I_;d�RY���m�!���dזq������iĩZy߲�iE8���>8��>|�rm8�띤-l>a�NROe�Y�'��9�-�f���6�\C�,uE"�ɬ���eC䗗sv�uP���2M�c<ϰ+:¢��y�i�0����<�3���S���a�%C���ܛz�Ɉ
�黗��}����=�}��ή�w �ӣ{2[�d���
<��R�n�<�E�ԥN7t�q�����<*6��,� R\.f��g������!G:;���8�V.�s�;�A���( ����t�b�m� c׫j�S}�K"q������+�O[��GG� i��<��C�Mg��[a��d��Q�N�Y�M�� ����l�"�L�4k솹HV��?}��3����a��!�*,�����bO3��>��v���2F��|��? ��*=�#�Y�u1� q+����=ݓ��E��W��E�N!X6�d�>aS�T�c�J�8�5a��&�����?g�ܟ2�߹q��0B5<~���"~�g@�!$N�0+:��$�/�}Ѥ����wO�T��';��x���bT8�M$b��˦�TR\>��OqC[g�N�É�ݚ@�R��N�s*k��{�0�B�{�����	����'�O����P�|��P=�0�0�Y=�5�<�Ag+�޻��PR/X=��6��b�S\�+T+�,8��Y���4ΰ�H����슞Wݳ��00$�>G�?3N����'C�����~�6�:Ɍ��E$��`rw�4J�f�9�a��p��
�ffN#i<B���T����`i&٣'��K l����9]�ߑ|3`xV��SL?3���1�a��?!Q|��1�'��7<��8��vOoQg������ͤ���ɉ���(��
�Y�����LB�l�rk�O��O��ìp@��L��Bt��,��4��%E���b��|�1���w�:�z��B���{�N�S�vLg�?8��߰�)�������*A���ɴ����~��6�Y�f�����c�ߞ�{�ǲ��*,Ͻ�;gRc���w����Mj��܅@�VM~��:�P�مd�뤂�̳�4��x�,=݆�z½d��߹�Ԃϙ+���5'|���g<������2e�!u{�G��� a	@��a��m�a�1 �_�m�!�z¢�RcXT�4��$�bj���*�S�RW��La�՘����l՚I��d�X��������S�o�;2�|��A��Vu���`mUI��y�6�Rm�q�;�0��B��ݳ����1'��
�~LCHWƤJʞ�S�i �B�b�N0�M�}ߎ>�!�?��t�� t3��9�.�h�����lmC�j�ej)�ꈈ=�ٴGv��aeLl�n�Ӣy��ב�&$#]��"ñ�5��Wd�8f�<+:�I��j4 g'[�w�CZ� xG�E+�.Rۻ<�r������cv�xxx y<<�kkt~�d>�� ��L*n�$�>B��{���E��0���4���Y*<���d����:�H)?s���������l=a�Ri8��`V|�A?{|����Ψ�;߿w���O�H):r���+^�11�;a������H,����h�z�Qd�?fE��Xu/�胻:��S��'XmԬ<�!���J���kB�d�ă���uΞ��cu�������zLC��ɧ9g1������6�Y���SMd�QAH�2�ĜVT5{���
Ï��L�����f��:�3�*)�� �:§߭CIvN_���w�=;o���/�53�a�O���>#�t�d�{;���Cԕ�79a�����#���a��}5d�:����y&�T��`i ��ў�X��T����|>>�$��ە+�"����]o��ﹾ|��'���Ɉ|Ιܨ�N���m&!��<9܆س��aܳ����Y���[4��°��aY?8��+75d�Qd�>��CHJ��f���2T����s���=��ͿvL���$��{�F�O�=dݓ�����m��;��O{�� ��:���d?%E ���������_�La��.%I�bAO���Ǭ��C�+�~������י�<����9���� �ϙ.��� m+;��;�:�X~嘊u�� s����*|��7{偦�W���p>���u��>���=�(,8Ԃ��*b�H��@��A��C��9}������{措������N���Vqg�*oY��T����H>XysP�,�
����C��|ɞ���(q%|O3�%I��f�w�{�+���H�i1
���wZ�~���n���o��~d�
��QC
K�Ⱥa�������
�Su�LM VVLC���E �k�jm�Pć��N��Y���ßa�N�_b��}>@�|,�ݭ�Z~�h�3���}��Ҧ�<q'�^��״Y1�o�|�HJ��,�%@s��N�$S,4���<e����4°�Rk�{���Af�y�9�z����{�>�@�����S�ƔMO��9����LJc��B�����!���[���۹��&��3��"{6Z`�Oh,Ў�]�S�Uc܎��dDw��*�����N0<vqi�!mt�1�c���X�f��>�x1S��+���۳y������_}_UW�otj`��=1 D��~O��#�D�;�juRW�%E�^�W���6�wf�|��8 i*�<�q����1�'�$٪�hT�s+���9_b���ݣ�:���{�k�x�Y�ӽ�m�E�w�4�RuS}�m$��*o���Cl��i�;�f���!����°����uH;�Qa�Y���R�4�A�����˙�ʯ���^�8����+�~ﺁ���Y��I���6�{�hF�q���<d�
��@���m^���蚷B�4�_	�շ=G�y�����DD�#W��:��Z#�a�}�e`��O�-��R�����ي/'�s�:�Y=N�C�d#�,�rv,d�ͅ�v!��+����,�3���m�F!�ګ	p�+ip�!r��x�w<Oó� �R���p���9S*���./5��g��$.�Jsli�$�����2M���(���y��9���d�}�c��R�*�4-XN��8�j-L���0dP�����!<Ý�M�Y�����sF��Y!��>�p�$ˎ�ƍmՑ����Dh�;���c�����J���P���Y&�ŕ�l+�>�nQE����[R��h��E��ì�c8Ӭ��mA'���볾}k ���t��m�qTa���?�I�)2����X�Ö��gr���,�YY�Tѵ6�}�:޷�rnj�W�����7�@2ާ�����}s{zpu��Z��6-Uf���$��y�q·�u6Շ�^����\doZTٯ��OW�l۪�z�[��3ڧ	7�}\U�y~�N���91Ǧ�,V��Y�����5D�7&���@F"�=b��+���t����{M׹p���(�̕���?{;�b0���=m�dŧ"�%PHF�}�$L���7~0�p-Z[�r1���<�[������x���+�k(��p�>0IP"t:F�58Q��SAN��q�J:�H�X�o� xNl>�iE��	�hV�8s�3o�F(TTN�-��o��7�S�5��(81{��Uy�f��8oЉ,�����i����fpPҖ>�쾢��'���T�u�>��?DYj,TY/1^�:���E�ƶ��2�눨��Nۂ��-0���oKa}	���ޣ��R�3h�*x��T��������uU���+'�G
y�}�_X5�8�w4~�ەht��	p\#���N
�5B��}(y�lD�:\#ul�����5<E+ݣ��j�a�p�Ϣ�Ub?+��1{��M`��%n{�,<^�q缷n.ī)iG�Z�w�vY:��t�6^2���=�*t&�.v30;;�TU�).���3���=q'¶ ����yo�l�&w'�o�J�-=ĝy����p��]�w�!w�Wl���NA���r�j�1Y��-��߇���dh[��9�������4�8X�m� i�������ސ�J�O	���겷q�[��:�k�W�]��2�h����)G&�1N(��tI�	u��yR�P[�>�G�Y�[5�H�>�R�7��i�
(���ϖ5C���|�*��to���M�)_�9��;$��$ YلwH��Y�ҏL.�p9�(�����g$�+;M�)��L�������6��VcL���S #$C�����j�p�UUX)e���V�^g2pޞ�T4�ŽU��LO��g�(�@H�B�L�dC"E)���×Kr��ݳ����l�lS��'6G_�wyPo�:%I>�p��	�(𡜮�����W���%LQ��"�q�Qؕ"���j�%���+�(�2"�������[��W�H'�[�P;x��ݤ��#T�-Gct��� J�Wj23y]�����c�@��~�ġ=�\i1�E[v*�Z�����zK���;�6	�9�f�C���g]��l�^���#|O����^�Õ��UI�E�-+x�ڨ=�O�&\x���=Or�_�������x8���`CC��q�Xڔ(T{���)�N�K��pM-�����߅%K�j{���}�A�h`�/.���p�_ ����~㢯d����.2W%%��-ٮ�b���a]`08�Wq�9�R�x��9�&JJ8��Z3���r��zr�vͮ+*Ћ	�����{���k;J�1��Z�O0�Ʃ�Ss�z�)�� ~�ב}p�qL�狔�6{�Q�G8hWVoL+PU��Y�M����ܶ-ĤKϥ��t��6�E�R���/#S���,)�'��=�0��Tm��ƌB��{l�Dn&�S����Um��lNKuJ�Z��I�3u1�O$}�!��U�>�oON�i�lx�P��$mxC���Qme�e��:�f��
���/�;FMhhw�/���4�]Q�.ؖ����Cܭ�M<�����Ь�Ƈ�5WH�r�2N���Qں�ppP��!��/W7�Y�oS��vk���`����G��	��u���
�A��
}��p����R��=&��ќ�0��ZT;�.��ӧv�2���]V���j�k�+�fU���@���x#T�&��Ï���t����W	�w��2oxІjxfw��ۇ�'�QƸ��d����;܅+7C��f���(q�ۍ�����h���ѡv_ a�܌�Sۚ^��R/M�3��+z�'#Y_	��7�L�uj4c�yӺ�!����Ȕ�v�M1�
#b�v�T+�%;�����s��]�k@C_��#��P������ђٜ�����|��M1F�.&��p���cOEMwX��^��Vu��̈́�ƌx-�p�Ojr��a �7x��}���jD#Gxi�Ɩ�ߥ�A\w&C֧7W�(�>�b��z;��e:��^)��,��n��s��Ey�ԩna��pξ���hV���3�e��h^F�$�u]�ּ��x'#W�p(�q��[��7���q=���PVh�'<S�]�j�vH3D��1o�X�fY�cx�
�+�j�9�%]��pb�Y1{�=y��_/a�15�3����g:zw��4���٭�t3�W��Hd��p� ڕ0�MA�8��w�У�kx�aG�3�2n�U&�Ҟ�bAy|��4.��n˔m���Vzk��g��_o��>���-x�v�f�)��=s�X�
%�����0^D��)��ui�a"Gtu�ɗ�{��&�:�{f�x#�i/���t�}�H.JI��=�.i�Ԓ��y��r��D*
�5���'��	[�F�)~^�`s�.��/[͇������.��ވz%�_����u���m�«�hV)X�[j�J ڌ��6�X��A�EmAR�ŊE�����b����ʒ#`ZQdm�E�����F(�T��Ee���Y��b�"��Y(�UA���RFаb"��hʭ�U�"��J%m���m�J�IU�
$P�H�(*!Yb�KlX�
�D**�"* *��cmc�-mT�Z�-��UF*�1U�mT���-�XңJ��V%iZ��+j%@Z�"�[J����$m��T�E`"��լ+Z[X
EU��T��dKjH��b��H��Ȱ��,F֤Y"�(Ū��T@DP�	X��,�"��IYUd*"�*�E�,djRЬ\�0lԲt0����˹	ʤ�����*��|���映��f�p����lĨ�ɭ�3�ǳ�[�;��[��B��{���0�V�ѓ+F���4��?��I}����>~�f��b�oEX�v��6����t7���E����iDJ�����ߋ4F���H��oΔ|�]��5�q[f�����9`�}XP���;]8E��15�.&|��Ɂ��6���q��L��Ư�o�Yl����e��R�mV����p<obM�M�E�-g��/+ڛ{���gz9��B=XqY��Z'G2��Ī�"�7^v�ؤ�^���:%C�W�H�����qu+9��0�z��A0�]N���t�"�-��Զ��N�2*fdJ�H>�Ȗ�MG6����V�v)�C�m2\ D dt��]1{�n�T�[)��s�m9�m�F��\��c�s(ۇ,�FC���R����� �q�O=�*����֑wyP�s�z�c�7Bt-E�˭2�x�I��S(��Iw��FF��!�A�s�,Y�����}H�yY�;Ͼ��Z�>�u	5���@�Df��ǩ���;��n��%sBK��5o%��l1v���ƅZ��=W/�:��]��X�����;���O"�DMD�4�w85Q��Z�\��U!���dY��1��e8OF��V���sz]@�D���_3���]X����}meN*��ӻ�<=�a�F���L���R;(��#��:�5�;�L<�*��vx�Ǵ(��f�]�3��o�Ǌ=�L�4&��"��]u��jB6Y���Y�w���qn1έ�K���¨�륣�B�q������o�Om���J���)���TC}�F��́pDW9�5D@�<iQX������Ҝ��>�+��l�4�!�=���_95S�����t��f�k�3|)4F`��bb��ڮ���'w�#!�݋�)��h�z��4���Ha�FJ|'*s{c��`�C��Ep�Õ�H�yqK�����U�6�l�CP�_�i��� 5�y]x%��sJ|���4o��μ'g���<|ЍQSEl,躵~��T�-�!���)�y����g�pf%m���vP~�P�W��LP�#ܝ�ɞ�]!�b�NE\�3�zzh�K��]oCr<�n���ڢ�C֔��S����G�O��$u㲖�a��!;iѧ~�F@�6t�o�DgcѮ����}.�Q}�8���������N�B�u��ۘKnH�x�5�n˿�ĸ�oXV�|��݃���������\'�W�F���l����ۓ��}�h� i��������l<�TL.�Ξ]�����*7{�0h��_ϫʃ��
s�cN4���^12M��嚝�zܢ)�v�eB�q\��<��I���3\+�V���q��XS:D3U6X���y�P��	�Ƥ�$A�y��O��@��V�5mЃ]����,�2M8ƌ�mU�Ád FDH��<ghB�,l>�|�3�F�����9[��YC��
�Ϣ�r��n � ��T�l�΋�^�w�I�ho��ǨL�{��B�T��oO(�q��`;��<����d����i��n��`��<ԇ�&��P�|���O_�k"��B��E�T�}�ۙ5x�<�%k1"t�!SWh��[��n�&�P\
�@W>��#
qh�&v����Z�R��k 1���/ϥ���qr���t|��|��C��.I���*/Z�Y���u����W>��A�MZ#�R��M(�7 HM
���b��B�+�G��E�u�
j��}�躆&+�e��8hJ}B��XΤ���I`��
q�<��Ŀr; q٧.3+]p|��핵w~x��Ԥ%��1���Z[��dłfN��-��!-�����+.
_nTY��!�E�x�6�}�t���Fu�,xa�f]�٥
���3I��s�����EP��;�ׅ�v�>�:aڅ�˵�6���������+Z�n�51�"�	�	��`��$^b�8uŨ�4Z��CNY�S��b5L��N[��|`�f�IO�#���64Kq^�݋"��f@��F^u�pTh<X/7j��
\������Ԅٯ.�놠WdЕ�n�N�W��*��!��ҵ��%;|騎l���n��w�3 �czz�J<)s��G���uƠ���
�8�`��)FO%\����R�'/���H�SH���>�Q�K4�i�⽺^�;�|����'YRp��P9Ѵ�H���0$�OS!X���d0�Ϙ}b�Zn��c�
g�$���I�X㷥��iv�Q#�dq/`��0dZ�V�St�r!�ϕ{�۶�<=����FUtS����]�5���J��F���gj�"��E�,���0�¹��|xVKVʸs[��L���:�@����Q��i��2� Fc�cJg�+�c� "s}Qz�r�8��t���q���B7窲�0!(�G��=�u�U�#e	���\�ȶ�;�#b������}��\��Q�[ڒf��p.�ê��ꂳ�N-�Vx����[��=K>���VY	(51�Ro��}�~u����&������+a�5�� {����p��Gl���a�"�k\�A*p��Uy�J�bK����x{�"k�	�M�F��Xx��;n���!Nl������t ('�
P��r����Z�F^`X�V=�L
�DY<}G{�W���ĩ�h�fP76WJ0
YK��DgHۘv*Z�X��Ȇ8N�>�ӝ~�E�`ح�n0(�4�Ij7�t���f.5���(z]3��꫿1�d��b�(LS�"��� U�b����U3�0��|՜�{)�tN��,l<���y|Vҥ�`�t���P�r���׎�"�n����nk�u�T-�/���,C,����057�6Y�4
�E�_��]5c�ʔ�Y�@[z6�X�|���A�Ձy��V�������k����'�TG���`��1w+�AL��*sC;_.��2�к�gN{y
e��@;r%F��Kt�v;��4.+st�,�pHg'����"T鷕^�5��ɔv��#�4�ؠ����ۃ���༇��<�j�9eqѱP�G�0�]N���t�"�6-ߎЦ�u�K�w0Z��o#�����tM�&�s֖���p]�f��W�h����au���+���ܛ�z}L��Q +#��.WEZs��N��9񻫻?��[�X�z���.���@M�2n���V�����ޮW��=HY�}�.06q���&�<���pZ|�'_%�����єo��O�Ӈ� Xk�v��Z
�Z�	5S�z��ჟ��ޛpȦ(���v�3ۍ����5�����G8�f5N��t��%�b���d�&�M�����hHWd��R�a��!v9Qu:�Û��֡�C�G���p��#3g�l��|����L�>�mر�[�k yY�;���
4�CΡ&����@��]Q,4bF�{2��y�-�'����x�?7<Q��CQ~p8�w:R{��5���X=1=�2��Dm]��N4Eѽ0T3^�dV*g]o�Q�/���ߡ�,���%/Xm�ս빦 �ޞiփ�Q��CQ����Ƶ����u�lR�DWr�;k�D��&�UC+!��8"+ܦ�Џ"#`�6l�
�����
�����#ISr��+0���#o��-n�#���t��1�D��hׁQ�L�6���7W\�o"�vCM-�������4��5!��2h&�mE�7�7��qh�������s=��(^*�~K'>h�E���:ܾǹ�f�_rK�l�P���8Gw��ŝtQ�j�~���$Z�[9����m6��v+z_"��;$=j��i�wlJ*I�o�|+2jR^]���F�.�%DLR��٘�X�uU�g~�π� x�������=�(뺯a�ܬ7����m0U��ҡO+�皫�J��+���or�Z�&!�#��#\TőJ�#
3uj�~Ϊn��qB�*�nF-B�1�5�!V��'�oCno
r���*̢�O������Cɞ�]!�+(���*v�e�ԅ٘�v�M������F�w�K9^�4�Fĸ ��g����������}�	x���4��u��7��<Ү3�X�䀃+���.��z�Ybݡx�Tg-�T2(�5��+;e�0%�|U>�>z�tN3��G&�*u����'zsA���d��t�E[S˕�Ts!	���B�P�^쐜>�p�2M8�h��m�ȢWXɜ�FJ���44TC�C������R#�<�cP���~��ξ?x��{�S�̜�$߽��W�{�1T3�᎒�����|~��^��3Ɛ��ף���gt�/4>GN��u2�q'R����|pl��e�/s���mh/��o������+�8a��2�g��e`T���5��'G�>���S}��	z�_��Bqاl�X��ɂ�H��.�������_y>��Ӱ�H4e�"� 7�ށ�*U9���W�uB��z��-���n+\d�:�����U�L���Ի�xxx	�Gu�X�w#�9�"�û���{CuY1a9$!<
�pT>���ϳ&���Ar�@����c�B�i�i���"��dsrG	kl��p�>1�T��痯D]B�1s�s5NjY�!�_�]"
��dp.\��M(�܁)�X^x��b�:1�дE��\��US���ϳ�1��tGJ}W�Vj��M�(��O�������x���DY6�ߟy���4��AȪN�M��=QdH��zs�\Z�c6h�涃����7�ډ׷��`��e�"����q���h��7bȂ�V�#,��񖋨�6�X�O%'�����	W�7K"Á]�F�ܪ!=_�]*��<�>YL�k��kxW��7c� vHgN��`}Ly,�v)�>��n�y���7c�q�"M��R�湇}S}ׅu��E��*Yy1,��3�Vĸ]��q�nE ����Lu�>�4��\A��}��ͧ�7Dr�W��V���Có���Qa7Lߌb�PF�K�5�L̘��|zF.��L����ڥf����f�q\�{�<qP��O;Q����B�5=�{�֊�1���^�yz�H�4����]����ݎ��s�KǶ9%o!���`&����l뜩�ۜ7e�s�B����z�I������%���+*;�� 5�%Nđ��#��)��C��n}5��Ō���Sd#o���:o��]=�J e�=���J����G�,튔�M��=~��3:�@�*{C�WW�̽�D���&g��k�(���Q��1��YY22D8���c�d(�I�U�9�X��:��ؾ�E�s�U��qN6!z�*,(bP�g��jD2��E�n`����0Y����+���DL�t�9��ۍ�Y�Nl�����N�	RO���R����
����x����[*�I+%PWH�3��JQv����T�`W��	6g�ӕ[]��
l_�DK���8�U�E�0kv[�}�{$�Ѭ7L��&w]��9��rf����dtLF��_�KP�~8(�N{ҝ���g?�:W2wi��!Y��8}�o*��p�@�4C�y|v����W��s�o��*���z*�JQ��_S�zE�M����]a�d<�7Q�M����DH��' X�Sǧ���-�)�K���j���P�_"�!�x����Xg��jčw{�(�I%7\�j"�^k�����{��2�ǚ��p��v�R�4��Qu��u��=����%�!��rd��˔���v�{*�~�_��{C��k��ZҶMAIi�%�{�� x�v ��j�F�ŊƟ�����,o�
��� �t�Θ��P��>G�`3�S��j�m-�%P���=WN����)���B�
Q~��m۾�k"J��+Bه��5������<��e:�ة
�z\H��}���h�td�
; J��/�;�cX��O)�;��j��=���+�t��A�b�C�(W^]���v�^t�"�-�;B���]n�T&�N����1����2�q��Gd]91��)�(u�2\ J3�VD��j��Ta����{.4�(��|hZ���U��qÈaF��MzP�Uԁ����Fr�7��n�^��a�V�ۨħ2���҈~N��p��3�6ļ��#�9�{՚�H�k�(��} L�}Z�Νq�V}��7i���P�C��'�y@��]���u�*^�D��+�D�B�l�t�F��CQnQV�ғ���owf&�eFF��{�����=�psǶ�0F��"�렍�Fx���jB7�7n�y��,_�-[�B�(r#��������.�\�u,'�P��F��Â���04�W��R��^��8Yժ�k�v��D��2��Y��Cۢ٤�2��/�`�/����|��N��*tF�OE�Ӵ��K�zC��	�<���T\(~~�`SvQ�y�u;k6��l
��L�u���p��.+���x�XPg��/)�$�c:�Պ���'�˫�GP��+�'cX-�2Gn����YtP�"V�x��*n
fcG���XJ�v������s)��n��[�f��@D�4/]�]��8� �n�&�.ЬKw�9ڵ~�Vq��=�#�{7���zYj�yӖ�m�!�`̴tL����a�SJDЈ��WB��ģ��Fv�+&9��8�fVW;QĦS��]٢��|�ZQ�$eIa�
:�b��w��8Hf���TB��pUww}gUڤ�y��s�s�{/�a�O�1��W}�]��t	"���p�s�k�=�ȹ���ݮ:�v�WX������xy���=BS�lJ�fHܭٴ�ȷB
��ͩe��n)�p�{2siP���T�ȼi�*��J|���ܰ[������+�=.�5�w�{G$ǍɊ]��j��e�jgڄB�,�M^�	����I&Z��Ʈ^��9����2|R���ׇ���W8mMg:�V$��-l�1Ů_e��vK��.���W�S�,�M�>�������t��=&.��Ḁq�1��y�W�Q���m5�f��ڠ��;n��1-���D_)3�)&�1g��Z��
��Z��;�j�� ���wA00<��e�����ʗ[�S����0�"�s��>������u�(�_;[v6.��,b�L�8�!$P5	���1$�4prC�"P����irYh�糟����>Q�1`��J�C��Mm������N y�wg=e��<�r�O�VØ����Kw�����c@
�v�Җ�tFN��sz�U�e�p������7]��Y�qΪ�}����ؐ�8��_���#�(������D�r���d�7U�����_YdBD�Ӷ/��CDM�$;�s�()1�N�[��b��t�w7�V����[����g)IXfv�yg-� �������k��gt�UUM�n�����y�p�>��T�`�V���P%�2�p� �p{����W�*����Iy�����ɕ�/��]+-Z�`���ڔ�W|_X�7Z���H�Ӄ�)e֮��.�X.$��6���z�Ǩ%8pmэ��{w�0�s/�2|E��gH����DV��<Bn�V�`^�Ǹ6��Xަp9����W�j���Fs�7N�A8����4�ȁ���k��g5���N�]oiZ�1�5��+�\�9��y��e�Z�����_E䤇�e�	�Qls7��������_s�$U �H�(��*��Q`��E�F,�"�b�,U��
-�TP�*
(�@X(�J��Qm�H��h�+YE,�*d��
�+RTkQ��AB�Q���X�,�[H,�-Q�X�+*�(

J�Ő�U�$Q�+PQ������6��e�T+U�V�*�-d�Qb�V�
�!D��YQ@�m�i���2��Z��QT
�U��j�jDDeeE-��QRUAT-��R����R�Zѕ
�X�VB��[*ZQVE
���*J�m� ���+T-�Qk(��eeJ3���52Y5 Tl�]��܋-i�E����u�yS�s���TS�q�U��U랍64���蜃}3v�������n���kn Qӿǧ]����`��#�@1�t�A�j4T���n7�!	�ؔ�u��WeơkyW���u�	G���o&��
8G�*+b����80���i��Vs����������t�I�[��D'#Af���T�d�#
1��K�ۗ#�]�����0pW
b�y<xɫ�ł�M8�jIa�FJ|'*nobo��#��9�����^$��a��Å�����zsa�3W��`�n��ҙ:���sm�;{&ݫ,Z�_��LC]����*�G�	j+�E+0�"�����8�P�VVp�t]u`�6��J�����<.W���P�U��Y�P�D��)�ܞ�ɔ+�uK"���I��Y��2th8�>�J��f��F/`dD�\�����JE;4�X�Qt��b�U�`�Ǵ�d�yG_����p���܆�ps�cNx6������q��T���e[{���ou
��K"��!�o�4헦�V��}��tb�Ih���z�f�e��ȟa?��S��gx������ �_{%41p�ۙV]��Nħ'�5t����
����q��U0�7(l
��lu�<�}�WDr�F�5��O�p��ú
[��[�{�4#�P����a���)-��7f74m����=��v�f��~���ـ�Z�0o��=p���2M8ƌ��ۼ"i�o&�D�F���a��K�(�"2�b$1�z*a�L���/y�Ŕ8ʩ��l�|��u0�E��T%_=jOP��/=T��n���N��||4��ݍ��k��|�f��6�Ip}r-���$��s'
�*����lBpD��S ϐ�d��ʚ�߳��:�}���\\��M��v�y(��u���DZr !B c���(�S�]�q�ټ� q�`;�7fJ�G�Ȱ�y�X�W�1�<e���GP�E�މA���}@�ǪVW����r��6mq�}��^(N_A2��s�hhV�.p:p�i������x�ux\��'6(LS��L��G�U�U����<�,����k���z�F־H���~>N5ph���T�u,��6͊U.��î-@�٢Љ�9M��sZb���B,��Q�����*��W9�������3R3���²�/#-X���剴T�h����Jz���f�az���[��(��U])^��kq{��wKu�s�m�����K|'[��&{%A���:��\Vlx��	�< �B��w:	�'P��5oc�������Nv��MT�5��Q���n�#����T_-�X������m��g; ⫃��X.��y
	�ȿ8�4l=�f�|M��o�C���Y9v�5�����8���*�/0QY�L`d�)�;G��+ݍp/`Mz�H�.=Kyӽǖ��:G9��C�b�G`w�no_Z�#ֺ�������i�1V���������i�mGsEl�d0�M�EtP�Z����J�z&Y��S6�Ҕz���m�����t�Qr��]E�>#Hɑ-��q�]�;��i�Ҧ�F�D��پw�������3]�&(��b�_��-�I�r��1�$!�L i)�YDUdÙ�E6�����)�
�"s26��_@a�(���q��Q��;0�ƙ�zU2=^�t�J\ܹ�lgN�R���P3b�",;��W�n�49��"�M�w�	0�(�A
8��C�%�$�ݳa;�]��H�"_�}�
3{\Y�X�R�(S���!s뼨)ȁ�:�q�B�;�h����V����Z#5l���N׏�}(ޣ<�`n�x�E�F�KVT!�n�̯#�{�d��Et3�'�R�5�z'sN������u�B{F��!�!� d�~��Ԇn��WL�ӅR�92��&�"�o����ZH}�p��I����|�8�ˋw����׼��rd�E�4�؎��x{�5��6�Nb>��xt�[K�*$a��7C�C��O1����v�<�:2>���u�Gz�������eH��51���n ʍ#&Dշb��R�y��`sAEF�[�߭Qۆ��V�sph'(l<0$��}	F���F��k��Fl)�����l"��)��^�YAL{]�pZ�(e��8�Ʀ�f�,��ȑ�r�w��*�/�2e�^�K}ݯ0F,����ص����
��`�V��읛#��k
r��>�r��膬\��}�U G�`a��U���#�9	e=T�uf�`mWj��C�@�E��ܩ�b���]1 ���%z�U��ҕ�	�� ��lGɔv%VY�ל�8�B�+!��Q=�I���F��+������j��T`����:0�]OPV3���-����������4tN�Ҭ"�:fÙ��=�WL,��:F��p��@��)�M꽊�p��v����V�atV�!�2�X�V��U��q�20�ڮ14'N��%��%#�������<�t�Z���v�W�op�<����E���ܫ@≰�U������t+��qi/J9��m-�Y3k����bpM�}�d˻��a�I���P��� /��[쾫�- �y&�l�v^�&�s����*�x���k������6�7�P�>'L�;��V��pߡWc�99��.���O�L.����C�S��sE�!��*h�2��w&�,v�g�V}
����Z�>�U�:��eM��.��0�o��6#�'XN@~<E��
WT+k��'��<5Hj&ÑǔU��ǪJ��w��:8�s�̭�7E�ϻДA.�&�W��vu�F���h̊ 66C�}�L�ڹR�}����݈=��xG�{&IJ(�d��%4��^7<�xS��iǬz{ְ}+=g��ߨ��C%ň��4f�y�5鮬*�O��,gN»���E�5gX�N���A�}&�vy;��9`��.���:kip@x��h"O;���«K}��۟Xcԍm��5�\8 �gJ���y���d�M
ڋ��H�Q�{�K DY-�*�Y�P'��h�^�#HÅ9�Y�^��~�w��m0U�Z@iL�tno�EN<\�\P�q��u����ܞ�\��>/�K�.��O�*��Z�^uSb��p.S�wMd��S�{P78<�J��H���A�-H��U�:jr�F^��e��LC9R@�>]�{���k*r\��ۙW.*��n�-���;k�f����CD<�b��\c����#�Z2�x��C.��LC�'�6�L �RpJ�O���ﯻ�����٬Ҿ�5��Bا�ykzn
��u���D��)f������0ع�����&+%<v�j ăe�R.��+���å�6"n0�{����iH�٧ �i)�q�N�˒����(���4�bu�w�A��X�ڝ3�mx��.0��)�Zo�	��K��W�)�l"�QؗL��`K�o�I�>�ъ1L�ق�G�k�+��Q"$�~C��3D+�H�\`�9w�Bp�Ǧ�' �q�ѡ����O�K�WJ��S]�����d�P�`�S�>��E^��61e*}���2VN���2"��k{� X5�G8���eJ(����1��3��U
q^�>2o_(�ռ꺑���;/Fqd	,;u��y���'[��Wh$�]G��U�RC�G"��C��x����1�
�KG0_WcT�C���QV=N���[��n�$E�"�%PHD��v���<^�Y�/���TC=[�QS����G�Ȱ�y�X�W%���!�
<Fںl���9���cw�K�"v�s��QއK<vcF��v�rg���zd�6&�P�%Zs2��]n�ܭk2���u�X� �
䲺m� �N�<�ɾ�oe�	�U�|�n�w�b�l�V�F$Vm{j��}��xVc{Nn����Uw��7�����}���n�w�s�E����SR0��
=[Lɡ}����T��I4����Л/f_	}�:4�u6�Uշ��d�m
��!1�qE	�p��8hn}@^uZ��T�D��F�ꮥ˗��"��F���P�p�X�/�*o�`�L�7l���+�5�(�����)�6�f%heD���[A�wS�W �{`�򈼣���K<Z9�
���bݣ��{�DV`�܁�G_Uj���<X.��y
	�Ȱ�Wdѷ�B�x��(�Ap������9Sá�83��:z%Y9,��`e��HV{z�.��ȧt�W���l:��f��b&fp��֕�W�2JԃtD�p1�P�:UeM2�tϑ�]V���6�7"��W�d���*z��S��N�N�Ħ'�D�lp�qB`In�*+�W�*��d4v|��f�c��Ȅ!��k��t�c���!��x�# Cp{*�}n|��1����&���:��a<L=�i~�gα�E9���A㒦�4ĎH��g�4���3����bpc{[����1����OS��Q46�m~<�����Fu �*^nq�&��pGf��My�
Kn�0��*�A�B�H���Q�����3�8�W�(�;�]V/#��� �-��K����ǯ��VGJ)^2����2��.\����عP�/�i�9(�~W��Uj픱�l�Xd����è��q�����]8�Og���
vaX4��* y�3�-���m�jIǷ��䱧�>�L�!��¼���;��7P���D�Ӎ��\�^u�������i�u�"
�}�!kOOxr�mƛ)E��#TZs�+}w�ẉ�΄�.#��k*pl���ފ`�u$���}@��F���^9�p��{�f޼��o[��s�N��)F����/����7C�C�����~����П(��K�z�5�p�<�r�I�h��	�j���Q��/LR�"�D���S:�v�
3�z�����(VE6�Q�=%퀜�	����}��W	M:�GL�N���6��&������5x�"*�����8�q��wܦ%����LI�/9|]�f��[��f
=\�]N��X8�S�)�`�j��`7O`Xk���[YiM��#Wx�(��Ҽ��nG
�'��s�;�V^Yl��o!L��@:�ͨ��q���tq�gh+U^	ֆbt�8e�Eʙ�j�.TPR�9Q;�cۻ�պHW;I��r��]�fM^�Y�	B���o�j�w%Q1�jf�"��cj�H�]7RZ���`������5b^<�R�wg56%�:W����s�js������}���|�On����?�Q89}
#!�]U�3P؎7�AGbUe���Vmnd��Uި�/y��=�Ҫ�o��Z�gD���(G�|8HFHɆ�c�-�Κdk�a���ӑkv!/ ޲�Ss��XE�Ӧo�dvF�䫦xl����&K�$FJ9o"kr�U���P,ٗ�kf,j�p���\+�jӰʰ������AN������M�u��Asp�+҆��'a9��K��n��p�>��v�Zt-Ç8e�\	�;��C�V8�fr�|=\�Q�Ѻ���t&B>��Rt��XV}
���7�>���r�:���|��QшI~�ʉ�2T�dX�`�b�Vס�6lGOoڤ5a���**�9��Q�ף�Úy�}��q��PP�>B�w�(�LИ�BqP��B$"#v��Dqj���ؑ{l0��n�K<]	yx{�dB�'��2v�F>W�!�W5�5d9�����F��'#��,�cw�e`�n���r�3Q�Dl:�Y��j��Y�`��Bu�'�k9�me���2�Cߑ��s��ާL�����T�VQ��d��:�t��C�n�	�[�<Ky���F��ЯY�]��F�[ٞ��J�*mY�_�m�Kk\���c���7e��#��[Wʍ�#^p}2K�Ⱦӻ���y�y��[���0T}x��Īϻڋ�͇�jbwS��e�5ș�E�s2�_i�|���F�`��x*l�d�̚��b�yʭǬy�%�n���� Ϡ�pѷ91���W,�=[���E��$3'�U{�������ݦ
��i��4f�.5A��K̽e;fK��M�n��j¡q��b[���)X���V�םT؅3'� �Z�+�n��I���*#��M�	���ȭ{Y�&���'C��4MM�]j�-<4)�p��l�u��2��<���,�Sv�M����9��6"j+V��ǈ>TXz
ۭH���-�=|�[��t!���=��\lӅ�ש��pb����3�mx����@�M��P�w{�,�`�SV��<�S�F��;e�.�ƅ�;g��8�)�>t$=^O��w�����s��ǯ�!1b�!6���t �@N=6�c�M8z-��S[�`ݻ�j$d����ndf�H�z(L Y�6)*W��M��f��7\Cb�hc�&S_{��L�S(��4gP9���=��֞�[�3]�@پF�up�☠Ւ��c&�<�V�";��Z��}�^��g�ŧ�e(�a���\+**ZK<��]�$��wPV�4�S�/or���A��c�m�6Xwy;�:7X����h�i�B�IB
-ӶCT[:��-�4�$.mw:O(��V,����)�0_�(Μ�)g:ub���M�B&��u�(��|�u^�)Y�ȐQ]���^3%��S:��������u[�JZ�6T�ѻB��\a�v��|l'-:Z��mX���0�������Wrǘ�t_uޛ���4�����Y^É�U���f)�R��s_b���}��ʃ/����� uo� ;ݜa=�u�!|�n�������]�D.�yƴ��o	-���=�nZ�5P#sr��K~�Zv���F��x���Β�s�뛓�+���jM�kѭ����39A��� �v�M�%�@.�S��l��z����7�v�K��ث���1.��ev2�v�B~1zф��xא���۾ܫ8h�H���zn���i2�K���)j�:��{얫6������l���̀��_fĦ]u�Y�n1ZT]�v2��X�C�/hu���Du�R�Q���kh���u��1hl�`|�طp�:�E�ٝ扖�#���1��w'�����ҽ|X�0��ܜ |��ȝ�yuN�D��Nf�/-�.�	��L����/��V��m��Vy�{~�/tu�o(;�՝\�W�F��E룭\n�l.�5�b�ApW\��xvb�yS����jR�������8�s���ո��'@����)M=���v��Q�¶��Ӂ;�+)�3���Bd��5Q�4F��-����Ƥ�s��3��d�^jTHĮ�}'F]>��}{�G
Vǃ�Ϋkr�C�j��t)��7y��B�l�(��Uvv�*u�B��O��4E�2g����l�uʳ�y�
�n�S�ټ�7�����Ѽ���$ݪA��) ,�ǐgY@���K��x�#z(�XH�2W<f��e=�:�b��u��Z������а���M|c�m+5$���e�x�C)n��;X��-�z�{&��5����YV+�����.���}�RWKE�3��Ƃ��f����s�����)�o�����\�\�e\�"��8��m[Ûռپp�C�=�uhC��z�����ɔ��n��if�7�+��b��%����.ȴ�Ruͱ�٧��5G���P�#��.�Zz��P"�A���%��Gaᬅ�'����:�A�YorņyC�Ą��
,���8Y A�CO}��t1�N�A�g��j:x�3��u3��(������>^��^��Cj���]�u��]8�ŽV����ڙ=�7K���4���<}�4�y�v��4���*��UtdTJ�K"��TDb��Y"�ʂ��,*AE���+ml-Pm���"(�ز�U
��`�(��eeE��jJ�UB�[e-��Ɣ�5kk)Kij��V�ET�� �5�+��ʲ�
Q��EeT�"�-�J�YEJ�R���*�	l�
��
!P����YF��m�T�P�
�"��Ѷ,���d�i*��*Ukb��P��)+*V���T*�e`�)+ Y*V@�UT�����#Yh�Ue
�VڱEXV"*TPF-B�*IYm%`*���jVV(�U�0
�YE�(�U%cJE�����VڴVQ�F
0�
֣Z�Z�,Y+Pkm��j�Z��aR��R��[l�JS5�~������`��mu#�Ե��kW�+M_H��T�ނ�T�[�~Κ�����\Aޥt+�goB/r�D�N��UW��[�ݕ������fx��A��R�30>��g�	�
VP�%O�ܚN�F�|��j
��{k�P$�w��^<�u'[�Q'|�B��0��~�0 �ˊ8�֙�y.�	]W"��t�����U*��[���d�NJ1"�&�ț�a�ރ�v����$i�9���"�Q��y��5�"��y�X�W-m�p���S�F�(�՘�U#�F�P!���L+ ������g@�so��P�y]�۸�ѽ}��4��3�t���SE��Q�1�]�������R��35S�q�"^�
.���y���b���}c���R�x4v�i]u,�P{�}�]aK���*0mp�o��5C�Rޥ �M�~Nh�#�8f����{��K�|�.�(�=��9H�+�Q��;��}Z5jįۆ�dnmSPz�
b���r�7���ɣa�P�4O�{���f��]�VN�q��y%�	�Ĺ���Ti�J���`�ٲ�Ld�)اh���+ݍ�	�����^���+S��C���k>���`�x_S�%��93y}n�>���cWX�a�-|S�)m����%��^�絺L�^���=�.?S� p�E�
_��/�M�@!���RUqS��J�7�yk�K�sF�gw�Ϊ�V3p����Wrn6Fa���q�B%�xNK�YS�W�T�(�G��]V��i���S��މC���9ܴ�Qt�~}7�m��\�:�/��iz2�WO�WN9Có�xIwR��n�LU�hM���N|(_)�y-҅N8J�X*ҥ��WP����MO��Ҳ��ҿkL��e�g]�D���.l�l�|�cV��T�'�ʞ����g��(��
�ǃ� }��(������D��[FQW��@{iGxB��Vi�;��`˕;�j�ysA���<�p%D��1W�Ӂ��"���x݄hs��F��g@�Ss�e�lz֑�y|��#c�#��iEݎ�(�,v�
)ENF���!
���Y��mm�il\o*��t HRO��E	��U�����@�Ҏ#㒔U���<��fX�0S�ܙ�#N�:���`0��D/��
D�7ҩ�*/�c�����M>�
���(��c잸�N��D l��sT���O�KqS�H���R��Y�L�;�Sѻ ��l�[��`ێ��!	܎���7�V>�毸�&sl��M�;�9�5[n�4v1�Ī����p�6h^���]�W7��|Ռwu�-�:k��G�������zm���l^���5b��۹oFj];��;]�m�W#v�S�:�Z��p���^�spi9Ca�&ȡ�}	F���Gx����Ĭ�ժys����1EݯM^;����-e�Y��x����f�Y�����)P�0T]*�W��>�!�!���ㅂ��v�p�vf�/5XX��=�`�t�HIV6{L���μC���S'�J��W�.�V[:s��S/�պ�<-�|6�Ʋ�)�N"�W��� ur�ě"b,pr0�X��m`^�"��g�iuq֧�̉3��x�Ϻ��9�y[�xS�Zy�:%F{c�&�z�p����ŁS�c�zv�[�k��r�
��0L�
jq7XE�N����[����Z
u���<j��<鯴�[b��|���a���Ә�Snx˅a�jӰʷT�8�20�ڮ1�]"��MѬ�HE��G�-X��V�P��P�P�����u�㇞�}]C+�NE8+{���'wO*(����0�.�N*O^���rtB4 �aG_�h�!Mo;��;F��+>�y�����(�F�/.�~?v��-h�
�SWZ������[��~;�V�S&]���Kʸͼ�4�L
��"v*��S��xe����7-��O,p�t�F&�{��6�Yr��\�tk�~�)�^�V�#]V¬Μ��*�����q�F��ռ�-�����A�>��BO�>��fJ�#�"!����V�:F���j��LL��9�yX.�N,N�9�#�)��.�����Ʋ=^P��F�ДT�p�L	ء8�X�F*20:�n��n�au,c2��Ƥ#u~�x�yV{Cu�����b@�<UL���'2m�Ɔ+Ou>�jW>�-�Q��0El.�o7~��Vf����4f�y�>�.��[���n�_��<=�~z2�e�;J��j.�/��-�'u0�0p��$��>W}iG��y��+����ګt�!`����Y�W���q�Ԓ�y�FL�&�0ofA���;{�3c2��s{aO�$m��$"0�ng�v������ݦ
���[�ꞩ����A�Ue�C��6`�]�iNs�J�?)G�6��})U���"��rbژ���Y�ƈ9�b5�!�}�e`��^}5�_�K(<�	���LR&x�X�Ь��(j�->���Ű��R\X2�Et@Cp)�W�[�x��5s���^���{ċ��:}�y_+M�wtWT@�����Li>�:����R���Ty�l��cS��^��cƩ��y �]$�$R���/f�(�Ї}O�ҥ3Pݤ�oeŜ陓�����A��IKY�:�����x�	N���֬]*�]�0t��X���Sf�u����n�ǔ�+�`�sh�l��(��lӅ���;�pb��Cj��v!N�R/d�=Q0+��j�*x��-J"�(��;e�!�O�W�����Tԑ�7�&�*����Dq���:k
�����b;�Bj���|�A��	��;�e�J�ɬ�	
 �P�x�۫#��
����d�P�@�S�IH���LX��,��fr�����e��k�	�E\7z��쩵���}�|Y�@�`U
q��Le+����D�~�r.��e��/��#�PN�!_��q&���2�# ��<B���p;7���zQQ��M(�N�~<�z��F�<�Eջ�*���y�����z�Fmeaw9g�Kv�����/����Rz$^K7`�<�X�z���]<�,wA\X��˂�B�DV^�j�� a֯�CYZ�:��X�j�^>?��p�U9}ʁ\fxP��$!I9��(���ax�9ș���QBb�bf�8���:�E��]������޺��������g[�ï�Z;&(��{�{����XU�Mկ
6s�����恓ku�|��J���Ps�ʌ�ۻ�GI�[�
7\��]<�r�[��p�D�f���
��j5oWnz�Y�F����p:8�'pg6��ݻ�5��^�}C�w��MT��^�5q;��W��H����=Q�f�1&6�F�ЩRX{Mn��(f^ie�[�y�E�d��`�yu�?���Q�|���@�^G :�N$�^`�Q�11{�R��ͻN
�ł��y
N�E��4l=��׺|v!m
�zW]f�ތ������'��	��s�j�P}(yoS��dS�v���W�rj�vM:é��	�0�QגE�	6[J�`0��仇��Jɉe�#˦�45�6㇄G^�ݣ>�s��`i���Z���WG�0��Ю���Z4�te���b٢�7¸�Z��[��&Ľ��Ŝ����Zo��ۦl�)��3�B;�#H�D��U������B�Ƣ
��7��*���a��7�^�T��=3�]|^ ��$�S�b@� d�x�́�־彸9�R��M��.�<T"�F��iGTg�����ᮜ@����0��aEn��i�����]!���r�ՙTm�ؙ�f/z���ŸDX���v��v!UeB�*���:�k�B���`��=9o:άڵ��G>v���="�ϹІcO�;p�:tp���m��]�"P/CZ��^f�U�o�3ӏGn�}M��;�������p� b�X��ޭ����;u8�X���LV�c�wvt��� �wB�a�dM���@H�B�&}��e�����;n7��Qf�NF�]5�D�s��WU��&%���ʃa�'�I�{�	E	��U��DY(����lj3�ϩ��v�.��U���h�R�5RՁ�̓��,������7C�T<8�`�j�(mm��)v�B>�8���w�7LЈ@�w��s�FV��VR����e�	ݬ���j3IT�5�+~�B�U�q����sph'(l<�&ȭs��n>F)n��Tsu)ބ�]��l��V�ƭ��м��]T���2ȐOl�r��׷�o���/%�6c�AH 4C
F���p���j��6�Kٴ�MM�87O`8x"�ó�nz��I;�<BQ9Oʅ�ϑ�#700ҙ��n�Ú�����&��2�i�!����uC���5n��A�{j�T����ׄ�o�3�Q�gs^2�o��zc�(d[��"��N�ߓ�|V�Y�*3c�$P�\𐌂2a��m�G�h	�Ky��Y�d)��ʮ!좕a�9�d���*��C�̟8�7�맢�}������R�3�����.���3%nE���|��̝E|#��򝦀����+����L(B����2fJч�/h���Ox������w6�ŷ�ga.`U�*8�͊%� R~;B��7XE�Ӧ\@�[���������ogwr���n>�j��P���U_M)���20�
��'a��Q��Fځ2�6#[b����U���ǾYKG�@G�O��ɡ}j�Fy������W1PH��u����^�y���+�`όt�Ƅ�
:�M���6>X�w7�+/E�V���V���cz>�g��P��(U�*x�/�����Gτ��:?�-7�l����ج�r"P��aHg�S������Ʋ(F�!�J*`�F��$�5�+.�13ϴ�xT�R8,��Q�/�<Ԅn�K<]	yxy��`�,�B1�8�7�X���O��;i�>di_M_67k�f��+b��,�`n�U�͈s����oB��ǳ%�P�n��/�UA^Pr0צ���T�=y��_�+�����3~}&�v ���',#��]q#�����{�����7�T�:d�Q�0B��9Y,�&��b�x9U�A,\�R!`޽���x�[:�s��"��w+r�x�����a)u)�X��t�&*M��Cn�[�7�Vx��qb�Mp�'�Ŝע�}C�Pv-��͘�y���d�7K�?i���$�0��\�V���p�@�<	�V��q|�����gJ���N�Ew�>[:��!��S�}����+���pB���^�"������ҕB�^�Ų��3�!��ƕi�2u����4�>�u	YG�(�Ĉ)q�<7�j�-:3x����cW1c�a����n����b��fĚ訌��n��b�F�[C�.�R�e�:�2���ɔ6�C؆�S�k4�}COz�	N+������7t��B��k��q��&�D8��B�i��` R��N���:�q��s��hdQ�&{f矕�U����?$4�u�ׁ��.9D_@E�t�`�[�Bй{��3QҠ���y��>c�\b��F�
�����!�u!	�\`�΄�����}r��3ovv$�@&T1�m��,8���؉���S#^���:/R�f��g�$Ù�[����jK��Pflu��~l�*�7z��쩰���@�.JF2U�\�uj�j������ϩ�n3T�&�響�y~�:؅a�Why)�P(�f
Z8ǫ�[,Cl�y���T��k�2ﵨl�MB�d#Q�aI沜�S
���D�Ol��>�'eP�̏��x�vz�Q�]�+�V�K�o�x��ʳ7Pc��c��(���tӔ��.�u�ܻ� g����=�����x���s}\�5]�42F�7����s�4��Y������4��|~�kc�^�����9�/��ն˜B&�O��8Ϗ�ïT���F��<�^��dX]<�,�
�B�ݓ�eM��V����v���c��:#SR0�� ⶑ�}��E���յg�C���y��8t�PӐ�hV���c����#�4N(�1N�3g�/��Om[�t����N�t6��n�C(��O�	ϰ�*j�ll�S�Ȫ��Hp������S�"��-�:C�^� �P,f��c[A�|^��S�{��K�(�P�G*z@Ş��vָ�w%�=����0m�魪n@��N���r��4y�P�!�$��D;�^�����:3��a�kZ�j���3��-�`�,�wN�k,gD�W56'���^�d����J����>V�������T����Ñ/��]�qJԆQ�<��MH����dNǰ�,�J*`I~�2�WO�WN�L�j�E/�-���$��c%q�y<�yF�%OȽ��`�b�+ަ��T)e�<�w�7�+g`���F�et��i�%r�ülЅ��6�$����j�^[�n�
dLͻ���/s��_���JM�@�RN�=U�5���?Q��⺓k��j��=]�U���Fa�f�	�\:���#VxAӳ�g�v�k�Fb�=�+�k���D�0�I`��օH搲�a�t�uHZ�@���l���e�w����n�	����7b��:-كY�˗]i��V���<����
쏳_+{N��b��o#ݵ�]����e5��*�&�\ɨ���yXֆ/����E�K�O5�Q�\ֲ���k� d��xM�)�!���{'n�uK�ް�[N6_um�i�q����̇X蚥G��}db�z��ۡ2�%f��P��.����.�c��Y�mM�+ ���GEWڶ�W՗ґ��r>��]f�0�m�̐ڮ�5���=�Uǚ�t���7F+��.���<�(nŶ���t��]�4�Ò��n��ה�hN"����{���&\�]�9|8��kB���[G44G�jy��h3�>���s;Y�BbҢ޻�xP�.��1}���0�g��kt#x��=�>u�G=��}�aX-<�:�+�(��yI��젴ҙ7NA��N��B�?Pt3Њ{Xf�L��n\�[�\ۨ��gn�
�)�+�H��q���Ei� 0
��u)է��U+�{��yX,��C5s=��a��L�X=�i�`Y]]�*wZۏ	��z�O��&z�	6�K�ٰ�Isv���^ڐ��Q!ٮ��Q���{'u�pZ�.(�Iijʵ��`�t�㋕U�̫��^��X���<�;��5�t>�/L�	0���b&�j��Z%=���z�ǵ��*�G`>�Y����+�����$K�b� ���y�5�3r���-6.��zk3��#��X].��MX��#��Sk�x�R�_M�f)� �0�|P�KMr��L'}���*�D(����z
>�zc�mHPU�v.�;���Bf�������r��=����k�8-~�L��j�<�%�˾{zB����Su3�@����7z��21:�ӳbM�WK.�H�;��{;�u����̛��9r1)I��{��
=�1I9��b���m�9Q�E*ͱv��֞�̀uŹ+�9YW/z��b����өCV��-;��N�W�;e4��M|!U*:d��;�v�xC���<�|�>E.�Fw����#n�>��6��w�!���EgREf�wFS��&^_f��iv,�.��_	����x���g<�b�&I���l�Eh���*|ep3���Q^:q�[����u|��7�����&��j����҇�4]�vA��V�$,����2��,����Cl��m�N_�B�2Ƀ0�%aX[VV��Z#X4��YZR���Q[b�UAd�TX�*2�"�	l�"J�J��
5F�*�H�H*�#+XШ*�T����DT �Q�ImQ`TXZ�(�[(%���aDUR*�,
�
�X,R*�%T�ł����")YQb�
���Q`�YR�RAIQecE�T�)�DZ�"�@PYm�+TY+X�A`�,�UKl�TjJ��QE���R)%�"�k� ��*�R��KJ����V�
����)m�h�����
1R�YFAAdU��l%��J��#V)FE��TA"��,��QDPA��O2��z��5���֍�؟p��M��k�w=gz���h���;&��k�k��y���.�cA��5�#���N�Oʿg�o��p��L��mB�݉!(؉#H��nL�B8O^P�*���Z�~�5�l�(�岦�F�|g��RuKa��<rT�F���i��h�\�tËK�j�����X�T"�F��Q�.�p/�Ek�9��FL!9~�ؒ��q�iO#@��;�"1=(�޶�fŸDXw7����{��B;�1DB"��d���>���FJ�{Lm D�ć`B�3��U�\Q�9c��A��Y���5Y�FL�d�Kw���r��p�����B�I>��%0uʿT� VJ>����8��:���Gf6(����(�SDq�-_��u��,�(8|%1c�T��񜓤�m�e�x����_<�s��G����K��n�%E狐	�j���Q���~��)��p�����9��iN��YĊ��y�-�X�L��I{~Nn����#\z9)�\fP��ܫ�9�u�:Y���*3b�nצ��E.�n
�kl1bd<��/z`9=u94k<T��*e�b|_�����c�͌��<�R�ϳ����2���]��8�����<y�R�:Ck�&�cw�*c�\���*M�E���e����/�9pҒ���~����jV�J�lqP�W��"1s��M����,�9Y2�4B���3���T���v�R�S���O=Wޘo�5S0�VEeft�҅����b�{�P��`����Jgѕ�Μ�B�c��B����@�'<��d���Y�U����`vP�i������q_R��:����:�
��:%u��l���L�q��Ydcs��U���_����!����8HEf�B�����=��r���܇S���"��-����M�aӦm̎���N�r<cAٌr�;)��P5�z���lbd��r��U�*aSnp��jǓ�ʰ���]�՞�=��������>S��MJʿT���p���T�`jq�����-�@�yeçU�����@��T-E�˭2�>1�tG�AG_�h�d#���M���4���rCF�Q�E������7�������i�S�bM
�U�%@�E��
V*�mz#ds��7R�br���b�-����q.QI�q�O���Y��B�x����Ɂ��w�U�9�Y�k��)�cF������ �V
�q�y&��������/��]�z�7����	�3&t��"��5�P]L���S!�V����{8����^ݼgL�s���:2]���=��^;�)�=P���)������s��>��k�"�E2�oQ�/�����<]z^^��h0h@�!�5l�/e@=6��?/�$i�>�F�U1|��}�H�gip�o���U�d��XcH�JiV�D+sR;pˏ2!�P�	��/=R\^s�[�^^��3a�������F��v�ZVVkhɚ�p��T�
f� Fg��+�M��e�;yذ_)���\�dU�1��<J˩�4���؛��č��U�B2<p���>V�\]罒`�&}���X�R��� W�U&�_^��5W�5j��h>��A�%]�����F��ެJ���{V��1�4!lq8�}�e7#=U�\���
V�J����^u�6���z�.[��!�<���1�I踆)t��Cp)�v�M����8H؉� ޺��E�4�[���R��Ԡ�\��G"\6ULK;��@�#f�,n�M�n*;��}}ީ�4睋�z��Ӷ^s��.0�
�hN��nQ���cf����"8(��p��L�h뽸8fm+!s&u}A�1��P}�GsE��xkg�3ʙЗ�=�@��{if��o�$¾��Dxxӷ޹w�O���Д�k�[���/��գx*.9�i�]J
�nԝA�ջ\f.lRx��3E|Zѷ����J<���O�������>u������GeW='X���*Bj���/�&�U�j;�!֎'eSBM�����n2�ƍmՑ�8�#b0p�=P,���ұg���s�%����v�1�{$�<��UO�G6eb�<�z�uB50(�1��x�7O�֬U�p2�'��ཡo����b�'�7��9_�!+�^�y��'[�9
�JQ �[=8�Fߢ��m�S��X qS�2v�5�	Ȭ�B�E�T�CQ�y(��U�p�[���S�H�$���c.��k��Z����bB�B k�0z4^J7`g���*v��f��Uj0����"�0�N���=p�>":J����MH® p+i5}��6��	a�5K�hQ�T=9І�ax\�1^�B�(!0=�qE	�pE6���`�_#��YÚ��^ݦ�>���T�|���%�#ɪ�A9�MD�33�E!j=�yg��<Nmm���}<��1�0���m��uŸ7f�B05��,��������K�|�6�Eg#��yu�9�j�;�m��۾��A�^Uw�6�v�Vf>���JQ$�Ii��������,�-�7s�z��X�|��������+��i�A��'33�������|��$Ck�����/e��j���XR(��ϛx�rF�}��>0qΆ&7bȹ�qB�Yy�m�P8�]l��	��dO\� \��<l�>��l��X>1�%��.���<*4�];�XΤ+�0^C"_nLݲ���f������pgO�u;݆Ed	�s`�C��WEqt�z[X9�[OÅ�j^G��T�WЧ
]Om0h��c�t���i�������O�����)EL	-�Eqj�vh1n����k1[ג�ijj��6<���gg��dSj;�gt�S�8J��*^�os{��k��*�z��{>UniL_��ӗ����{B��_�p�%�}č�J'Q(O�s�j�tn=|�/��~����JE�B(\���}4��0j�p-�(��J =�4�;]i�h7���Y����;vc��������@�=(�{����+a_y��1�����{+w��f�#���*,8az��B�5"
#�~�Q�;����Qo�Ѝ��e5�{f4N��t�k��s�+}w�����@�J(Lr�	��G�S[�{_�\�'�Y� ��[c�Kp��d���(�y�ͳ'���t�t��
���.T;�H7�Y����4��{y�֖o�-;�*����	�>f�6mʺ�V�LU���l�vq���}������eA�(j	�kN��5mNJ.�8�/��n�y�w^���΋��T�~�n��,�2��8J"DA��3�5#
C�9��߻��f>qf��RQ�G����O���f����Wo�`��X�Q
^3�c�m�c������"$,0W�S�Ҝ�u<\�9��1Ǥ�����r���`I�+2ꟹ������������{�cO�=Q�3v�7��"�ˮۃ�m�,�֠S�U��Sf\-�wܑ�3`�CnofB2Fh�D��jrq�ʜ;C;V9��w걛Lֶ罕���<ήbl��R��ӄX[5�5`u��#�}����5a���y�n�υ����9gY{�`u�i�
�ѥ�ڮ6�d�Yc/H�*W�����C׽�R�a�yLR�ϭ%x����p�֕Yd^7^v;�i�)����^��#�2�*|)��4��{�f��ɍ�*]���-�;B����N���Gdi�J�apxg�Ut�HF�S�R�EY����铱���\/��ōSn�p��I�e 2s�t��@wSX��4��4t�Ȋo7���;����f"#ݞ�M�fn�(�9�B��|��q��SV���q���a;������R��r�A���|���A��!>�W���@|E!k��یg��܋{^������E"�9���Z��Į1�2��@U�'�'N�bS m)�k�dкT�cS�b�5Y\*�3v�60�O1yn +N��p���'Dq��ЙEЙ�}[���F�8gxGE��ᶂ�O-�������p>窄�T��2T	�dH�`�uB����t�Kox��N da��)��ƩD�r8򊷕ǭ>�#�dQ�s�B=�:]�R�3ٝH�<Rqww�t�ئ�6��7����j��R���7Z�.�_�gF����p��F�D��EAQ>��U�M�j�"�/˄�|�zK�hz��JS��}��U���P�X�da���cn�T�h:���ף�p��3���n\�A�)u٧U���3Ή���6Hr'�p�h׈�L����d2̝�`��D�3��P]�����L��'�S�KM
چ�'GO�'h�^�!�z*�����=���pqc�b3-qj:ᚽ�`�m�~�h:�͘'�<)�:����U){�}��X�e��^��G�EFl��T�5[��/�[����,��x�}aϬ�\\%w�U����#b��Mn�;ұe9W{+���4̩��t�8平��7|}�3}+M[�[]��3ٶޓת0�;H!so��H1�5�<��;�q�j���m�yݡ�t�v�����ջ�t�b9GÊ�VV�i�{Uv=����id��*�<����ق�Bh�o 3�Q@�Rz,�@����Jn�i����79��\_cC���}z�;�62"X��ģ�6M9�.+}u4�g�
Q`F�8X�z�#0�[<�[y��,C5z����9�q��^0&K�5¥��@��"���"�ĺe����S$�{�Ug�Ɓ�#b��hZ�ݳ�q���~U��b�>��WR��A����7��k/ކ����(��D�#\1�N�L�`cF�6���8��<6OD5�qSõ�p�ޚY��ͅX��T�Z��-��oP�6���0�-Dok��\x4i���7��-2E�{w�˲�H�,v*�tP��kz�Fj�p$����{XN�!8
�H�٨�ב��̈́��"φ��&K�.�kb�X:"/T�CQ��.��� ��]�O ^U�lJ<��VH��jD	��($#`�\*�=��`0�8��Y2ᙧف�����,���
ܕ�5���O1N��/B�JU��I�{6��:�Se�M\�b��0�4Ӂ-�:�G9Y��}�-�Fۭ���s�o��_#t�Ҏ���s�TG9��NC��?p`W���WęZ#Ƌ;���6�lwV6M�JU!T}-m�Ń��GIP"t:F�Ԍ*� :�FI��XH�7J:�*�U���ZY`�Sa��J,7!�4+,�t*b��D��&�+vz+۝3�-m��$�H�6Yx��x��^��C�D�
j`瓟avT���0���uక.��jJJ���۟,�ъ$���W�ދP7bKB]A���<��)��DS�!�2v��;m[���L1��N���F	�Q{��۶�X-�W���,����їyo+1=H���E+�z<^	G2�vvv��F��t��c:�,���0[v�+4E�dGc��zغ2G&)�>��^�hp/(l�C��x�V�����$�c6w�v�v�H�>�Oܪ�<��f�`��A�+�0��'�z}�Hq���)E	�%��+���-��T6��~�=l�MS!��4�[8��LٌS�1L�tj�0>wH`��������]�W?U۟*��S3�ӗ����>3�C�VT�D9*r6��Wq�t"�}�Q^�6j�Yjͬ�Ϝ��<����6�2�ܝ�
�+������ʲu���K���kZۍ�]lz�T=��P׬�!�����o����lr���w]���!�M@�-�3V��y�Q·�sa�ƇY���y	�H���UR��J�\2���Q��Ek��c��um�|��{�@��<<ՇyS���ʮ�/���6{ư?�]���z�uઢ�	����.!z�*ah"Q��B�0!g�}��T�qG�����j���DJ���e��.����
�]�A��@�$��R�\��I>�g�Kʾ�Wv�K!ȽD�(�	��^9����~����@Aȉ�	D%z+{xV#�[MNkY��|�*'�������� �;u�?OP��yU ��M'���gy��/+/�>���Yą�Z"�s�S�T���L�q�/l'7�r�����oXy)�F��[��^YQ��hO���:�M�o�v�4/�E_�]��on�9@�f��U�9���X9Q~nofl�:!�>�9��㇕8w;U�9����"�D���O���m��
˳Z1�S�bxS���UK�������7c�}�Xu9<sڻVɊ���xU�K��!O����2gm�	U���wJ���H_:��cp��Q�!�)]f^{H��F���������{���O�R���������Ը^��ͷ�:	jL�}鉩&���^����bY��3��i��ƴ{H�<׌��ބ��c����x��^���F����K����p���9�F�/�V��e�9p��R�J���Wb�B� �0ep���̭5�EW�d�{;|A��|*ٚ�=BqVv�@��{T��ܹ��n���kb�D.�Gb\ 9�8�P妑�o��ױȖv��fhuԹ	�:H!��$
Uu�,��!yW�.�� �2��`sM)\Fd8n�� s������]��_#g�R�o&����m͒�It֋�0H75;+��i�XO
R�XM]�vn��u�uu��R�w��h�ЫR[k�+'��Rr�(Q�����͌�fB^r۷�4`bT��h�����r"�#-9|��Yf��������Z��h��Z��k;�o�n��(��뉁Y�ýKX�D
~�hVQ�������)����,�m�B �㛧M�Դ�޺�D6�dI���=������&�5K�|h����w���҄�"㢱�r�w�K��%+�k�����Zdm.�R��U�ŋ��]]{��h�m�4���w�wgxd;k���<riѧM
_Z9�����9u0�xT�]:]yN��Gu��}M�4`�9�N�GK�u�8�Uڞ��䘨�Y���%�vxdמ��476ĐT�v�	�T�ohT"ڭ}7x�����^`�D]^~�w=ƌՙ�F�IU���y>���=����ٺ�}g ��[��k��ʺm^,+~T�c&�u��v��-�p�P6�y�CЮ��[����A
�-�[�.�9��]��O��n%�^�r��&{7K�I^^�B�w	�R�M�'N�>�Aǚ^^K���u�,Zp��Z4 ��v�C$q�����q�}_z-�m�{�x���j������`��t���vJ�<�s�+��&[��Fo�po�'��{�/[�W�WF��rCXc�y��]��ͪ�T@e�/�V����$��u�K� �졝q���5��I*Q,�!s�ζ��hl�}v�nƧy�7�\E����ջM�F�L�G�u}��R��|r��Kf����k��v�Hbm�5��#pˣӜ?�i�7��܈r�=%�NHq����M�w-F�ky#��s�v��Q�@��dg?��˳cB�:�A��]f��]ʷ5䮦���c3�:s����|nE:q<��c�a�y�WO���{�ge�[{��ÂلSܡb�t������eÂ��)��0{D���n���%mG���혥��EY!o���^:{0�s8��u�`��Pq�� �V��N���3�����f�S�i��m*j��In��7Ǉ|#OZH�|I�$���ڡX������+R����m
�!Pm�Jʐ�E1���U����(ԩV�B��Œ�X(���K,��B�T*A���H��Ҡ
�YP�,�����@Y!P*�(�U�`���+b��*���Kj�R�Z0b�*¡D�Q�P�[`T�
�V*
@Y+*-AdU��(Q�B��J�QH���iDJ��U��e�"DFUH��(��PK`T+*J�B�B��Z��*(�e��(°�����0��,5�-��m*Ŭ����*�F"
��Em� ��-��T�+UTEXŊ���B��R�*"*���
,�ŐQTR�VT�����߾<u�߫��@k��i��ӽ��b�{6<��|��:L�j�{V�r��~%��:V��t���Vᖾ���>=�!����'�!L�R^�VmF�q�ջ�A�D�וX�����"�qd�v���r;�UzL���q��AGbUe��Ϛ���_�j��Tg�:"/}����7�]��ٶ�G��a	d�����gM2/������n����J�U�pf3w~@T�:�~�����;����AT�]c�����4�1�)�!�2�[�B�`0lЌ��ea�ͽ������.OP�=|�`�C*`�<`�d����u�8<]jd�[=�.r'MgG}*�t@�<�qaˬ2�x�ǽ0�����>�ӑ8V��1>ђ��h,���^�5��+>�y���
4���&�P�%Y��Oz�R�'Td��u�Uobun�jF�FR6o��oT��l9yE_�W��n��?��4u�~�/^s����[���ǫ�.��v�5o��ߵ��05!����З���7Z<
�܈ww��4���(Ą'OP�;E�{>��;��j�"r9p�o��O�R�!��b��P�{����Fk4t���MIW���2���-cO�,�mu+��=�����L>kM������eƝC�v�F�UcS�������'})�~�of]��T�	y��[��-7F��c|r=�?>�S^5�S��±�� *�޾#��������C�lx�]�PV~�F��=xV
���
�J���A�Df=�j6�v8�`�Г�wQ��3@�k�S�Q����+6r���2c���쵒�-*O�P=7bߛ�p�X��)�9Q������LH�.W�HFAÅ��[��#Q�0A�Kok[�}e��zsa�#[��MNJ�����x��5]�@Ͼt>����^�O���{��ʆ&�a�W���M�G�a���U���kϤ-����j��w\I����=�Uk'��͢� �֏R6�9=�e�.�7��k4���i
��6���DK��8J;Z��G
�F�:�?�]C�����	��ڭ�	�1�gܘ�@���-��=��\Y|*Y�N��"7��FT���m��]�%�T���`J��Ȥ�#��:1F)�":�q�Cc�lGX�HCV�).#Q���4`��hA������,�M8��~m�~p; +��ϥ<���==2�����S�j���#�B��)�;cd�dX�۳�`]ϐ1��_f_�LMG��bS8�\� �����/]�n�����i��%+��!?�ks�4����v��&��0�N�d�j�W�t����1����J�J|O���]�)�5Q�9v�Zq�送��B*�,�x���u��a�(��7y����jc�sN7K
�jb��3^�ףOP��{��S��������	-�Wx��':7�E\#$�>m�rS���W��3> 3�2\qWS[%�c�R"�M�5J"�v�h��jyj%۽�0�s��=m�d���P�bB�B3��p�T����نy�����ؓچ�4E�#T.��
t��Z�.2�1J|D{��>��R0����K+y��x�E�:�k�(Nl>�iCp�
�Ë4s�S@!F�M�J��WS��U�k[��9�7��B���S�a�Ħ�������]s�\�ֳ�9}���!��1��ŵ�yy�4f�U{�аֱA�We-��s",��nщ��i��3p��C,p�s%d۽Śm6s��^�|�r�;ׄ`�x�_���຾ڿ��&���7r����o3�s�ӨT�����Y���{�e�>�9Z�)���c�#3���� �W*�&�r����J4�j��%s�u�-�"�{�51꣬��u�/�_�X�����^��S!����uf�O���PN��m��y��ɝTby�#F���(nŉ�u�Z���7�{��Y��ױ5x`py8%Lc�s��;�u�h���9��u�h}a�7x�;�u�ɯ���N��^R�{���I�=�M>�Չr���*��kL6�;-X|�ۦ��k����'����E��@��%�*}��cjP�\��QYԛ�z���Ҭi+V;��ht�9�y��-��V�$�F�ō˄B��V�Һyu��HXɞ�����{i4`ܙ{��WNo�\ ��Y�lV�w�ڞ>�3`�v��7y���������W���JaW�Q�\CK&vD5S`�E�S\��L�w��]g0�-�~�c�������}7#S"
=�J`kB�f�E82h�X��s)�Y��Ǳ���m��Ϭ4��jz���)�2&���^�1�K��׷H��#c՝�������[h>���C(��0�=}b�	�t�L�}�z��Lu����eok,�1�ծY��}�N.���^��#��g�����7wݢ7n��:� K0�+�fݕi@ye v���Me;ѫU�y�vHge�:�8-���4�\�k��5����u5��*����D�+�U�7�J�:O��/S����N��������w� ���C��Gi�[藎��H��5x�U����B���7��b,��D��A*ȡ��C�fJ]i{�
��<�C˝~�op����s�T�T��
�հҽ�{]�a�lMuH�Fe!A�YHTE[)ocW�[ٷ�6��ëwJ����n�}{@]��v�L؋�k&�2�wv����̮�93S�:�]~]M߱�v��y=[���;U.��X�O��jV4^Ȳ���"2[��W��{a����ɻw�M�YK�*,#3�b����b
�V�.��tHܘϣ��o�ET����eq�\���⫚���&z��0�c�����=#rD ����kQ�G��Dh=tƨ}e�DM�O*��5��h� ڷnC�t�0��F&㦮�jk2<�����b
��h])���*M2Fp�`���|�����PښwgJ�Ԯ�[u��p�ض6��b�֔�D� h�!c�_2����n+��qB��z�U��u���z�NY�eb��S�J��<�\�0H ��^�N�S+��d��1{]��ć��lW�w�wu6���[�s@%0����͇5��7���*�]�ʴ�~�R#W��=Tԧ}ʭ�u'��ϫ&�D+Y�u��q�4��WC�&�g�7��3�ꎾW���i+��>t!��1#6�̚�/�4��6��#,hN`ku#�
�Tw[�zs�]�FͣA�#rh���+i�JfN��a?`�9��O�{���v��Wk�X�"�r9�����>bW'>�.��s3�����&��|72o���Ӗ�Nk�47*_��tݴ�ډ�|2h�"�����<1r���f/:����O{��*W�/;4f�ucu�Mc҉���V����¸��9��o)�'�C�̞�N96�󩰰o0�_]+Mk�WFM��{T�ك��.�1�y�k"X�0���="-Ҍ�-������4-�i��Bl���6��G��-�}�`�u�u�ڜ�[�OWʶp�Ťy[�P��En�N��"��:Y�%�#�ķ�h
#��n�݌(��V�!��n�쾥�&v4pj�xN��cI.����:�u���	�@��Y�/n���|��i��q��Dr�򝓲����W�bh^���	R#%��⛙}{%ss!J�ܛ�;-+l1v�ϩXt�y�,���^!��>�Bi�=���2�i���8�_s�
�������A6�8�ďdo.1#r`6;�-�YV��t&s��+�i�mE�I�=MX�:ƏPm[����oE�f�]�f��þ��2��O
�%
�gy�_Z�UO�7}�޹<�Ú����9b-k�;6���"�X&Y�n��b��y�r�������qp9��ɂfOo*��ȏ �w��`�ن꽱ܯU�AS�,.����w����r��:�:��d
	�  �pJDj���+p���َk�UՏU����`����˰dD@��hh��E����yoj�=/��i�� ���+�6�B�`��1<U�g<Lu��璶i����N;d��vڿ<t��&��CV��.�d�R@�ݝ��dd��h�]�A�=jkݩ}oEm����;��V�ڠ��9�.*��M�qO'������}6)��B�%��7}8U�ʶ�%�{����9�}9���D��=�W��Nݴ�ѐ�ʛ��qmn�,��n����Vhu�Q^�}�XU�,�f�U�-�qV�k�������^��;�_�b�u49��Fe(���Ŷ3i��{��7�M�B�'�⵱6i���V�ؚ�Q��}�̥R�嚅���#�R�x� N>l+j_zZ������&�py#��\\;��DD_��檂��N�0���n�v��Y����:�����E@Q'Wv4�HXn3\�U��KL6�C媓t�y�,Xv�h�5�"FɚǨ��t��'Pu�ٯ bwK{�������g��]|2�Fl5kSSZ�U�3�8nH�P� RF����]6[\܋'8��2ԭИ�sX�ES޴�Ӑ7ϑ��iyUઞo���1�=���9���9/XN.k�О��8h�F�T��][Qȱ?��r5rힸyx�4�7�[]�wa�4�=��g�=�J��9ŹN���6��}� w2.1^���]�Z<T�ѝBs�,R����4���j��Z�(�_76ț�ɤ;FU��ު�ҮzU��S
�����	���]UL靆-ڱ*�ff�
�W�V�c�����Oq>���L�AGy!�H�:�C��yNw+�;%�GEgU��p�4�������o����N̝��aOov�h���"�W�(�q5�݄�����[jKBݹs$��9�"i�i�����i�4&c�d��V���Z���	{8Y'ro��٨<N�v���qAEC�'Â�1H�x�	��y�j�ڭ�G�\;�O`�������v��r�)��M5Y��}����>���M�	�/������.��HP̝cs��k
�V�4���և��4:����w8z$Nd��lj]˳��+�-�����un�Xmm ����Ȟ�9Ր�*!�{�e�8�\��e�'�ӿNLԶ;
x.�����>����gf���"�Jt/��j+F,�cCOu;KHe��K�|iV��������r$R�g˦z��6�>��9�C��·�y��V���/f�OF�$6�p�Q��2&�*�����^K_y�]�`>�)��fE�P��8��Z%�b({�qxo!?.0$+��\��n�1ʯ���a�;-XM�S�OU�n�Dۃv'K�CR��0:1��K�X�1#r}��K���TV*m�1E��l���s/q�t�[�iPm�nV;;#W��"}X��'0�}f�r����z���a���/���ucG��n�<�`�ᣊ��6�lUr��q�N�v�|�w8�3M��SS����~m*��=W4�TZ9�\�u�z�h�囪VXN�S;0�P;ܵSR������k��MY'�;�'�	R�� ?oLΦvDb�:�^�Ϭ4����J����4�孈1)4�A9Ln�ub�;��=9���Yܴ�w���q��&���7T!�:9LOcCSؠ9�����2������Ռʤ�B������'��ъ}�@V�S'ӧ�=��QuhQ7��9a�(��ӛ��Mf�飹 ��ƀ����q���Vu4B�Y���ͺ[����r:@K���|;���eR�۾ko:�V��nV�5�3iW�ΠP�eUwt�cz���<'���9P�B���������u��ѵ��=���9�ݙP|U���u�r��V�P������/j�6��yk�;��0�Ó��Wh�9��+sWB��>L�o`Z��{���p#z��������]�W)\�V%�h����Z�ؗ��:t��N2�(L�`#˨\�Y�}��
[yv~S59S]�K\-=�
��'LO8��pZ�Q�Xz��}�öu��Eg%�X.����[/b"�P�Gi��.扲�lX�Pk:'���ڎ�z��s��EV���+{R�#`a�ҽ������x�ǅ�ᵼ_����S։�y�wt��9ͮ;Z�q�'N$�KG8gn*W�UӠ���>�Q��R�_+������{&��9��B�S��^����{(�;h�C�<��9�/*� ��6�๒�a�Q�S�U�q���F�QN;�v��K:�{�l����qoF��.@��K���S�[ao1n�'����ã����^m��:%`����g]��6>�NS�Rp�M���U4�o67CzUI�o���U�Av�jA����T���B�����rA;�[ f�Ī���C����"�Ul��^�FGv��@��q�Ë���yA����x2���ۜ��b�;�"�Y�oy�j�C^.�`񸎌����9e� &�D���:�p�݁p��˸H����G;�7@G�=��{]�լ��uB�J|��V�Ntn�U�K��#9@mj�4%ر�d4�K��C��A ;b&��y��폮�m�Oj��R5�(NYD�����^oZ��@x����E�m����8�+�|`��=A��1���vv�%\���E�7;ׯe�S�sB�V��U���8v�J�܄D��2��vVZ�l΢���hn[[�J��r�%lLMo{�f�$��[�B���El�8U�m=��z� 9��ܻ.����(��ܓ�k�;�K����_��������JJ�}�ɜ���;I�U���wpze��"��!`ud�G`p۟�Op���>�>���^�N�,;+dя8�K$����D��r�������2'��}m�($��X������D�U�e�3j������cM5�f�����g��V������sk���N����E�u!͆.�B�$�|ڻ�b��g1�4{��9E�0��f��1A�Z��9�R��e�.��>;���!�	Ԡ��"�h_M�E屗��75���ȗv�{)�˾�6��Qe����9�́�y�]��epդ��:,^vq�j�+��vڍ�uS;����V(* ���JʅQ���j �Eʅ��+JPm�mXVV��F-E*"�J���j-Dd�FJ�Ѷ�QU�H�
0���T,De�kR�ذ-
�le��,PeF��-���-l�+m*F��k��HUe�����m��5U��� (�ԭJ1TEJ%��)R�E�XV�
�e��dYYR�U(�KmDaU
��T�ER��R�6�����mB�)Qj*ZV�F5����1`��D��m��-X�+�� �Z���5�Im30q�Ea+�(5���h(�����Qc-R�*5�Ej��Z�S)q�Y+b���EX(,Pr�)QA`�Z�DER�b�T���Q�U�#Z
(T�l�B�+&e�E����8�m�Ԫ"��Qml�Q$UKk�ZKJ��R�RUBڰ�5(�Y���+VګJ[m�1�"�U��F��mw�(������#C����δr�	)�f�ꠞ�}�o��ز|4u
��\q�xr;U�2巄�����Y:�[C+���V5SvO�Q!>4�dV����#�us7�\ ����|=��R-y�O���߫��r�?wZ�����Y2�(eΛ��Q���Fe+�Ssk,gSa`�a���=�o@�����j�?u�������om������[�~���lu� ��0�)�F���{*�Fy)V�vj�ȗxx<�K��׽��%��~��`m��k��a"�\�`&�ۦ��,����vC��	g92�1���
�����UCj^��cb[x�O��M�q������X�SY�|:���y��sϕ�
�1(@�̊Ԣ�e&�KI��ڷa�d,�f��3X����h�:[���%�4t��ʥ����qWֺlv��e*��%�t��%��7�� S=M`{h|���%S.@�Fk{�ⶦ��*�1�o�S�B��~��b"��HQ���X�hա:���5����u�_�{��)yt��"��}dfp	�T{�i�ӝ"��fu��S���:�d�G/W���C���������շ%Ĥج�O[�,[�t�sА���<#�^H޺3�T��\Y��U�ha�����	(��.!��&vD7Z{���0�'��-m����}��ں��3���@�Ȁ�1�"5��SR���KV���r-s/uj=9˹ږ��5a�v�"`hjtHuӳ��;�ܠ�n�jY�-�$(�Q5ڝ���a��ڒзe�25�mY� ��^���܊�cS>�����Y��M^u��N݆��є�c͑YUH���R�m�WFv���28c��n��M�-���U��h5�B�f>��M��;cnU�n�+��$hs>�c2�͹�Ŷ3i��Q�f/r-S�[؅�l%�P	����V��&�Q�$`nDfR�94�<6'����֦����\�3�t-�w-e�n�^���8<��.�q
g#��VŬ�;�����������Ar�m{�`:n�b���c�f��︛���/۞��*��o�݅�em�^�w����em�wS����^���"�a��
��w0�]�	�X�f�)�C�r��J�%\��3���fFza�M� ��;��l9���_�.��4waa�L~���9�o�r��$���:�k���p��2���{;��%+ؖ��i�݇M�q�t����L��*�&[��e�;�s�YMe
���կ��QYԛ����*Y��{��&��Չ(����^+q�
Ξ�!���2kQB��I��/�Ar!S�1��9O����ӝ܎�5����p������/���5�z�-��]j��7��j��isҞuJ�S
�B��]0J�r����Qej�皒���V�m��mvi]]=I�rL����Wl_Glu�P��J��#��c�U@��k�>������������\�ة���X�`1�}qT�X�w[^H*�����Æ�9�}�������>bLؼ
�c�bx#�D�+F@m��Z�85P�#qV/���0�-���<�u�Emrھ��~�Z�]��]vR^z�1=N���
v�֞쇣�-_h�[I�e]u�a��1����{�9]G$[@��V^돀���_h���f��'9��+��,F�*<}f�L�|.w]�@4޴,�J�w%3M��2Wo���ay!%��vP�Wz�qb��ص���H=7L'Mk��K�4���Q:�ł3��C{�>��hB��A��5x6ߵ��ͦ���aPjؠ�ǳ�Z��׺�`X���.�F�TJɖ�\�sL���|ka���B�\��+mmy�-���ؘ���t#�k٪��Q�$�+�!.c+�5-���Z�n�v��D�9pw�3����\`��m��u昐�|8J�FKpym��ca������'������R��y�2�{_�gf�%Ь�F�ȌBi�}*-�5�+:�"p�őIx�g2�;|iRm�r��q�aq��p��B�#h���'c8t<MT���6(Z���4�F�=�m[e�1�F�b{��oF�i|[ʴ�z�Q�lV�*j{���m*��=W)D,��9�[;�^u0�Ʌ�R#B�;"���>��U���V��w��{c~i;v:��g��t����%�m�՗gqp�N�9k�P9;�z����~7�3�<�aY3Iz��zӥ��^v���2si-����q+]�	�9�`�.�ٍ��;	�ۉ��0���1εhu��<�'M�֎[m`x��Sw"qꋅ�R�rNwllj��Dy)��T��b�:�X�y������y=V-K칖p���I�
�b5��x
d ��G)��Ԏ�S`��7��F����m��7��9����P��;.��9LO�#CR"{�!�
v�� �-H>+۴py�\�o�zVwXnL���e�25�O�)���'��$�fJ�y�����;��y֪�Sw�Q '�%����s�ޘ+��tʥr�4&c��FcW7�/qm��n�n���b�J%�vR���^u���3	��w�f�_��0��Y��qϮmft�9��KY�;+��!ڷ����c��U�=����c��*D[�brg�-���71���ⒶʚQ�M'�s�NU�oV��Ȟ�8<�
�%����a^���	z�{��W:�4'ge��v7A�,���^�$p��yRv��B�����y��+;{v������7u�qe�87c��	����
JK����$�^�}��`�S�v�q+��Zļ���}�d��]��Iqu����+;F�i_Y�k�aX�f���S�n���:��*���5#{��ܶ���k��Z�lKo�j×�������p�C]/K��S�DBV�u�Xڔ"��E{��xz�|e��u%�#�F�cz�d�w*qrc#X:`1���X�����]=�v���K����ף**l�|��,o;�Ja��}0�U�1���+T�tOX3�\�����y�y��r�X�zS�S�(�.��L�n�7i�1[R�o��X�ڭ���h�]����Һ�S�B__���I�#�Zy��71Iqk/u=��)�e��j=[k���j���y������Wjh�r�ڶ�<�f�� l�Gz�S���a��ڒзc��*��1�"�Ns�S��ʠMC�3dD�QYV���:�X���A����œ�8q��E`��w����C��9�L��#�	��^b��v���4$�ʏ5m �8@f	R��S
/S7Rīg>X���=�so�#��a�G���}͡ذb�B�G0ܹ�d{��Ϧ-'۪�y��@z�Õٲ�DG}�2+��dH\/v^۫#���NSθ��M�$<���
��`��'�e⇂ۼ��('9iRNܝ@�A��D�evU�[:���xc���O��\��=�BDc�(ڊuլ�]:���)���m[�ؚF����Z�r��(��k�������l.^�a�r�KXܬ���؛Ã�ɨ�s�`U���l��g�s{3힣-�W�%�0���Sv7N�7A�,����S�6��N�]Q��{"�b�댖�Lr��J�%�����ۖ�k�����1l�j\�`�����XZ`Hܘ��B �ί�E�I����97�uOqfD�L�g�<�x�ە���Cp�(>�(RF�kQ/hM���Y��:���D���M��kg��Z����o�g�]v��.�:��u�S\��`j���+jo����C��A깤����v��WƲ���G=����v��������5b��Oq[��	�QzT��v�Y�h����q��YED��2e�8�Y�o��:�4���~�v�FR�J�F���r���Y�ۚ��'!��E�K����z��ļh�(��]3�=����w����В���w=����#��KUޜcX����e#�a{�}{�F�c�_+\9�������\�f�y1���NEOA<�R{���h��4��ȍłC�Q;����w����+�6OU,ކ+E�I��TE�gCwؠd�s[��HFk�⑃r�v=�K�YZ�vr�˅�\�P֎�[Wʨ�_��]27�&����Fwc��8��?k�ņ���n%��j�+��$hs<1N�R����,�u�R�>ט!^17��X���IՁ�¦��,߼�-��1�6�>Jw��]��e(xrD�����8���^rg0ջ���^�͍��JP?3���3�6ǂ������^B�Kvԡg0����9��]oo��8����x�Y�-��]��a��f���a���mF2��n��ٹ�t+� ��>�܈�$S� 
d�ʮ[�9�X��#T��k3':)�RK�oq�!m1��.���۞[�����I�iGF�����4u汚]y���x6p>sbw�Ľ�v'�]	�m����^�t.���>wt�&8pNU�^n˵P�ٸ9�íېb7������v�Wj�㖶�+��a��Lt4��0�jܬvvF�\`Hܑ>���1Ƴu�%�M��P��i�mE�Nl:|���Ӽ��˸}�v�ÿG�4�Ts�n��Tp��3����5<���Ҫ���o���)E�ls��p�mD9���?wO���gg��P;ܵSR�w����y��V�������2�N�[#Q�J`>T&vDb���j<��4N����w��+�Orb__��gɑn�O�j���ւ�'�`a#�?t�Cz��*������0��1��V�=�����i�=M+�Kkb��f��ap��ܙMv�g\��R�ڝFz�+�| ^223mrܯe�CW��!��MXͻf\9h�J��7��fe���U>܄��hQ���cqY���u��0�1M(%�9:��n98��ly��Y{ָ;%�]��se�ᾆ�;���ö�"�+e`
�^4��٩$I�6AA��ǘ.�m��2��F��Y&���ӶG����6���[>��$�ͮ]�V����SI��;y��]�+h,f9�9#�"��5۴�u�4��Qa���W8��6�:[��ck��;j�I��#t�&�j~|��Rʷ��4:�`y��*.4T�:��3j�Թ�=��A�t�0�}�KԜ�,aV�yb�젳�z��{пs��u^��te���%T?)�vᄬ��ͺv�q^kk�X�0$<�ǐ1�6��u�W�+~��5�P����ld>Zg�.����p�A���Ql{B^C��V_��3B�.��EvRo<z��ƝcG����S�S�/���mL}�8y
Θ4qa�KI��Ժx+��c�h�QUHEA���cI�w��ީԦ����U2�9���5�"�����aօ�#*�Xv�ջ�A깠�����(�����4s�ΨV��K��Lj�i�UJ�*����� &F �	@p���ٰ�йΌX)R�X�4�[O��hb�Rz���2�s
}�_VI`P?^"-C�]��7hs*���n��n+�"n$�-�",�R�����p�U}�n����1�^jn� ��I�s�OA�vqF���xȳKب͍x�^ܫ]��òJ�E�v�S7�ڧ�p�z�sk�8@��PS��<��b\l>2G��Gn����8�^� g��;�[n�q����|�u�H��s�G4�<޽B�'B�o�ܴ�ڒ`��j����?'�r����<�>����ԧ=�Y�v���t�F�wm�8d����A(�<�=ؼ&v8nP� ���p��<e��+���Zk����a�f�SvN��p1��n����&)�,魁� ��v����.BإY�Q�ڝs]Bd��X\4æ�a<��94��%'5�N�O��<��m@�Y@�<7��y�ۻ3xS�[c� ��tM�@Z��:?!t
��c1н1�C7�kNR}M���E_R�CVFT�Y8E����ރwB�.'��J"��z�u��^�:L�z	ʅ���(H�P�������k��i*��,DM�2������PO
�W���*<��!7KX.W��+����{��O[��e�nۏN���v��{�ذ5Z�Vf���Z�u�7�[���#�ٽ�� ���^��>��\�C��Ԟ�O�Z�k.�ls�R���{�"}P�4;v�p��ⴰ�]���]�JF����� �YI�i?�u�47��u�Š��#V��Y{i�y_�O$۔)`cqt�;&<SE�"�ӓ�[L$�3Ա\ޣT1�j�j[��o	(@�r����bBiL3w���5�6J��+9�&��%ֲ���7���!����B{YJ���7���ы��&Ǥ��8B��V��d�׹�f�Fw�a�]�f�ݝ��t\������s���{��Z�=K�:p��WI� �޾���X�������s�+Nw��R�50�3�P]���,Kh�r�ex�='�ࡩ���l�gooa�m����t(>�����x�y�ѓ�<���؛.�x���E��Y����˰B������j�毝�ԕ�n��d�P�OH;� �캑�;�/�=�+���p����}�ף����M4x�e��	R_#u���*쀕�t�h�o
�Sﵭ���^g܎c�
��ދ�ˣ)|6�"{{��s�}��q) ȷϳ
JN̿��];5L�P=���	Wދ�=ʛ�쐃��6���M
�>[(���X��KL��LO��y�����NF�Wc�On����)��U	�ί�E�c��r���4[�rT��H����o{���'* �sU��V���t�b��:_i5�z9�fT3�»�[޼�|�y�7�{��
�Z�l��TXTKUm��l���D[-�me+KmJR6�҅Em�+(�d-����kER���E��d�kU�+TJX���6�b�6�%��5m�L��m�%Ah�YTE���(�EJؕ��ԣ"°mm*,�Q��k�
��*6ȫR�E�J�Q���-�Qm�Щ��E�V�U�V�T��Y�E�AAE����YYm(ł�R��-im�1.KkKZVѶYEZR�`�-*��h�Q)J�2ִ1m�T�(ִ�Ʋ�̣U���ƴFU�eJ��b*�V��S�mKFԭ�m+���
���J4�hƪ2��cm��ڍ[`��QQ��JF�T�UbJ�eW�Qr�9�*V�-X�P`ڵE��)�����Z

*"�0J�l˃��(���(�KYUJˉbe�m����b�U�j-�bZUU-�*�R�W<���k��aT���\6�<3�2�A���Z�K��.���զ��ס^;]yS���v
��XuF�[�{�0��sw�\\�쟄���w�j=9˹��j����7�]��E��ѓ)�U��݃>��Cp��`��V���� �ߟ	\��B�GU�.����#���[���~ݘ����������y֫S��A�r..m]'��2�����w���y[^K��T��)j]�J���M.�c�4�y�f7ha��-B�q>y]�mV�xs��xc�̥`M��5ݏ�E�w��.�^����1W0�w0�_b�׵�V������"0E�ժ�U�|�0J�bTȩ�rX�aշN嬯7Ku�dMY�9�\�yG�pz�l���iߧ�>��Z�n�7N�7N1fᒲƎ���I��|��l��OˌHY p�1��Z��{����ϝ�ã�M�=��Kd^��g�v�XZ`Hܘ��,S�}
7�:�w���[5ץ*�`��W঵<;Xu����%f�7g,���yx.c6��	;�����X�v�C�6�^��]v�Q�#��cz�J�k�ڻ���������ϒw�T:τs-�
����kV���g��U|6�M�}"S'L�[�MN����O^�W�+r�ێ�V��P}��$C��;}XwC��9ջ�HW0��\���h������_��C/|�D �{�'��b�7�u6�b�����6���6ު��T=�J��撘TB[k5l�|;�]��������b�3�	����5[]��WW�z�=�o�$K��A|��S�q�֨S�H�=��[�$l
�U㯕���J�SU����L)�J"�$Ѓ���Z!pr@@�T$:�+u�H*�Wg���o�'�M�h[��Qѣ�_�ҕY�����n7:\�h*�]��]���*�V�󇓒����i�T��K���VB��%�ܗ�L�54��S׊h^;Uz��a�b�mļ�MVE{]D�r17�Wz��r��O�=��5���E�v�m7W��j�֖W��f��>�w�wW�Tߴ�������n�].!e� ��;���;:#��蕀5Nv�'ƌ8A;�WgC�s�q�7�"���������w�>�ݫ��6��M��%�p�XD�������ҥ�N�W&�}��Z�\�W;m Э���܎V\��!�c2���qn�9���;u+[[9O N���w��.�sOZ2{w���bj���0J��X��-�������U��WQ�R��zغ3ɇO)�[���:�LHw��o�9P���q��UJs�olG?��n�n݇M�q����B��`Hܑ��i;�r؞3n�B����c\�c��=->2�K�r�ۈ�5],e5�r����^7���.�_1(Es3Z�W��9�>��3�1�ͪ|��5l��]��8.�E��<�	,!��0r�&\�3��q򦧝��V�T}��F�e�c-1��u�s�jZҸ�Ζ7&6�]��!��6�U�W�V��wܩ�c�<ث�);���U���	��%���W�v}���Sp��MԾT�҆y#v��r"M�>m]K������+up�ކ��j�c,Q؝�(z�<�#��T2�~]H5ęA+�����O���ҧB��P��ŗ�,W2�}���F����|5�8$�u�U�Ѷ���|�BB\IF�W�b1j����,Q�a���hO�1����;�Sd���$��r�R�����f+qQ�T3���]:�U�͎�r�d�J{��5���_�UB��yLOt5D@�<"�h<����5���될WtMvۿoN��J��Mz]�:�-]���3z���f�Gۨbq=��&�E�s^��UcU6�c��Q>O�L����՝�k&6^<U�2��?j����c1�������^k
�V�7y�%eF��/j��~�a�ؚ�Q��L��g2V	�qj�:�
c=�4���9�8-��������U���5�``y8%L[�brw^V����0>5ϙ��#p�Z�0�ۦ�[y٫���M���W����q��ˎ�O���ߥ��}���m�v�1f�k�^i�X�'�#s-�/)sj*=��)�bE>WЗ�m�;->2�&�ذP��-RFv���޾�&2�HǤnL�P�)q�֢�}I�=M_�ܟ����QU��ϪXW���J�I�>���.'h�"��`�ێ=��.���x�v�X��A�4�o��'f*���ve��j�:��Q/L�9�]!�/��������F��砉|w�Wc���Z�u��Nu�E���^3���}I��\���_.���(��`8�~:xh����� RF�x:0��E�Ǜ���&��λvd�Wz����R�G s|���e�r.ud�ʍ�KRw�Ncq�T�<W�o���_��P	�T�sA"!��>]����3�r�ל���Է��|�;J���ȼ����I�d
�Y�3��!P�ֻ�>�p���+\�G�l.�k)�-P{��e����&�"����sC�|��9;��(�&�[H)i��ڴ�)���I��]�т�*똞ƌS藊�7�x�м�Uz��7NH�h�/�${RA�#)p�Tf�J�J]c}�e����������5�S�vn�t�k��Hy]�~j�(s��d�3)%���Z��UU:7^�oV5x6޼{�-C��B���ǳ�[���&�Q���w5]�=����Փ$�����z��LˊA��vWqB�Χ|�dpzλ���i{}�aW:^TG�ؚ�=���Q�r٧��d=�,��0U���rg-�&�Vph=��o-�⋹;�(.��-λ�9�qY�kN$oRԒ��KWX�5+�9��g0�[t�KYA�[���'�����.ɲ[�����Ya��!،t�qH��װ������n!�ո���6o��z`��oϯc�٦=!d�1���r��J�Ķ��u���S=�9���F���]J1b��ִ�7lv	B=O�_J��f�1�7�����}���pSɀ��ƒ^r��q�
Ξ�I���F󔮽-9� &�zv
&���-K��.��4R��w�޵`��^9}�� ���Y�4�&�?9�w(�Vg`�F}Z��MJ���^�S�sIL)9wc����`����x냟.����t�6w�X�ms��������X���n�$�.5Hz�����֨HجUG_+�>��V�錱��BY*���7����#]���|��1����V(�+u�K�t����Qfs�lo�yCv^,�n�W��Sy�/|��rm�[�w�g�ur�,~-7�,w;�c<EJh�c��6��9y��%�P�p����,�^�V�A��@�p���
%/{{$`.������7�1n�������m�d��j���oRW4:���(���6u�Ԗ����v�]{��[}^dW�P��*Fp����+��S�+i�N�Brrd&�;�a�)]����3؆�2\��gZ���+��~�͚�v�T�b�K�-M�{]E�V�ꤞ�O��:�y�1H�Ʈo/q���uy�*jئ�Pk�F�	c<��'��g�دW��r	ou�rX�aջ��[D0������18�e����c6�ؕ唫:׳�,�T�:��Avuۥ���8�qݕ}Z�0d�[���yA=[���:�LHw>�*c%���nY�},:��|�B��89?��7n��s�4r]
��bF��n蘜��\�'|�%b�vo;r⽊�y��վ4�&�p������%����6,T7z�9>�<+�
\lV�Ҝ�}mXh�PƏSj�n*0L`�\�Z�72_�%�����d��,�C��� �l�a����k.��iy�>� ����g�v�t�N�ݴ/�C�N�mvi��h��}p���*Ky��7S��=r��J��ϧ�
﷩��1�oy��WP�h���oA�b�-�J.Olp��ƅ>�T˟BFEo8���7�w�SiN�a���}_}͈5&~�w4��TB����J#KS��r��ڝ]���\�)m�+��N�ʕbK3��ɤ�AP�%0(���N��'�WQ����������e>�4�Պ|�����x�ȏ ���rka)��d]s[��#����m+�z����R_Xo��
��[\��W��i�'Je?_k�~�~�[�#kT]v��.Z|%spu41�vQ���[7W�Jwj2�lļV�M�syԫ��O�P���[�V1�}��/�S����:�(�	{�V��}I��J~�t����:#C��{��!e��'��*ؚ�8W����%�q{*�T�e4q�~IQw��em0��)XMm>��a��OI�$`����/g9�����jχ_<�����!�)���:�#�=�/n:ޛ�X�Sd��F��a����q��8�H�+틹��9��U/man���-	g���x�!�����79�Eo���o��`[�}P��j����|Y.I�u�	�H|j~��o���w�r���:my.���m���e7�{�ؚ����q�^m֢EW#ݩ����S���� \�v�^;-[n��n�b��6��Ƈ��9�B�)gqw"�B�P��F1K���KL6�;-X|iRm���bI̷�����L��[k��ˀ���
\kZ���&����-Y{T��F�_plQ2��M�n�q�i��GL ������p�5�"�B��˚Эe_Kwz�)-l� ��i)�@�{|�a�e��|��$C�'�8�v_,��MK�ަﺼ��A깤��ywL:j�/F�ܭ�zG\�&x�M�w;�|�;J�_"�'Y!2	�Swoo@��+�{��~��<�߲���C_>�V��\�MQj�����";��5�q���L�D�+V�����M����f����tG	-Z�"՚h�P��́�[�\�B�RX���!�h���y+{E�ʡ]kՀ�kP�lr�<kS�d˨��=tknOq�<��#c[��ݕ�1��ө�S�=�ѝ���b����絜j�F ��H-Yd��-=(~�`�TE�ƌF(�����U2r��d���^��%ꜭC��h�������s�̎�D�w7��0s+4�7��3+_�����MkX��K��V�s������2&*mf����Y��VWZ���9��_b�ǳ�Z����V��}vw���UÛD��oH�N�'&jR��A���J�.��0rdl�O)�4c��s�{&�%��X�*}�ߧ�s/�aֺ��ct�#r�1V3���-x?w����j�'c+�%g`X݉�T/�-0�Cr��n�ђ�o]��~�֭�u��#��L	���%
|�e��H�c�*��ֹT�s��<=M>2�cIXV;��CNp�}^��ȼ����]�k�re*����Ca�)�	7�~���{�py�B���IO� IO��$ I,	!I�`IO�H@��	!I�`IO��$ I?���$�xB��@�$��$ I,	!I�H@�8B����$����$��$�	'��$ I?�	!I�	!I��(+$�k=H� �[�
B,�������+��7�����G|��U��+�4�I�OЧ��54hz��Sj�����2    U?�S(�       J��D��@�h�h4 �  ���ԙ�i�4�F� hh$��I�<S&M4  A��0 ��h�.���n ��"G�l������?"P`?����� b� 5��@�EdX�`v�g��\a�O��<�t Xo�Q'C��`�Tm��XZ�n�+�`�!+-Nտ�᫤	¤�����C�ed��p*j)Qh�4$4	(�K�+A� ˔qT�'KJ�6{�cǰ=%�N��2A�#���K��(_ü?w�W��T������:ˤ�\�;K��H��W6#;խ��D4��S��(Q)e���➽>�pцF�l��^���8nHnŷal�`P�]N�ز����iA�dI	�D�� #�%�*�H�|Ha,�8�öԌ-�\3���:3��y��G# _���m�^��%Bul�Ĕ{����U�l�C�Q�#��!*���w.�;q�9�<V��f�"*o��N��� �e���Κ�g]��f��-J=ѳ+r�5e��:�mYT��r�ڵkԊ	Nȸ� #���֜����)1�]q��WMZ\���4�d'8�<[^ÀT�3zV��ԥꊚ�A�7�X�P#�F�q�f�����15�p���M,cX[w�d;	4Ȓ�!^Z�V�*&*E^+���S]]X(1u���d��k��:.�����T)aU��y�d� ����X�#���u����v�8��:C^�0�D���bc�uqpֵnؑ��E�@e��C�=<ػ%!ݙ2Y
RS���Y�
���)+���H�2bȑP��J[n��.כ�����3"�ke7[S% �,��x R89:�����4T72a�Eiu
�q�qQҮU%ա8���!���Yɕ���yi��obD;�u�	U�I�iA�VQD�j�FUvb��v�x�W+�-�M��:�)p�,���Vp �#]�!�T(�YpP)u�!�,B���-#.P��tvbԊ�l�M�s�\̜	��/��G���i"I	%��Tm(�{ ��Zv ]��%0�P"CWj��%���
dEu��P��֎�jJ
��ܐC�(7G]����K[P|�<P_�I9���s�k׶xgƻӐ[M��V2��E�c����'��Ry0�@(��`8XX��/%:@^��ù;:�0It."/�B�}��bKA�i{E&�U �=P��kAR��$���^�T(3m \�n��A�D	 �6��@,��@�f�\����W�Vm ?�*�m���=���d����u��]�Ǽ���m�ڸ\��̓�*���ț��#���j�!V�~�4��wRL� ��P%
��B�U�b�6�!�ɯ|�S	��ү-E����
�(���8C@�a�C]�]^��g�(�j�N��4E�:��Nǥ�Oj�'�@t���YV�;��i�TlL��F��<<����P�kbz�<�! ��6���y��V�~$[tL�Vi!������` 2��i$#7fā��j<&� F.)ph@���0�66c*��2��X�\�F�J��h\�����>S��wt��]�$�Ti�T�Z��y���l�V	�=��*�Gf��顋���BO��u'P'AjK�Z�	��T�7�l�F#p���ت9���/h�H��f&u���cS���²�<˖H@��tW_|ʇgv��m� @���^_Y�u�8��[�Q�9oԜyrInj���ÿF��`�'�t��X�\�ՠ�& 6H�������X�o���͍s.S8�BTΠ���c�R�AƖ�����! �D��Hv��\�rE8P�d�:�