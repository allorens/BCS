BZh91AY&SYY��s�ߔpy����߰����  `��h     �j�4   V�2�             0:P    8��L �� H}�|[u���]���᧦���`1�v�0
�Y����,���݅����w������/CW�޶=p;����=U�w�Ƕ�(7lE^   �`�:��f5��n[ٽ����}��I3wog^�P7��f)�J������<pֹ�]9ڪZ�C�s�ܺ�gZI�w^��;j.   ������vw`V��v:K�gYm��-����Q�P��^���v����ۮn���S�xn9�]�vS6�;��   �pV�}�v�s��Ӽ=O{/fzwi3nڻ��V��7���P�u�����[��{3���7���Z�׾���|��>ˀ  z1�{�ۛo��y'v�vp8��rw�F�7�+�w��(�yz��0�}x����>���g��6˻�w]��       xk  ���AQJ%BT�A�      J��7�U%���`� �����i�OЈ�UH L  � 	�F&�Q*U00�CL 	�L	�$�@%RP�F�  i�0 @���� �dS������<��0�m5=M�SR'��T�` L�0 &&C ������T��D*�"B�C��<0_�UTj��(��qQ�QA�����T?�� |�J3��_�7�
��A d������
B����j ҫ��  &FA�`	��K$�S냨6���j!�C��/�7¼�_���;�lQ��ϰ��s?�t�g�8p��!���&m'~��k�&�sG�3���T�Ѣ��+f��r	������10s$��2IgK�:�N�N�:�:��NhNi��/���[5��vn��M���z��^gC�c'���YFV��փHm��:�S�Bp,�(�)�i�BkIB?s$�JG�|�����I�1!�'16&�2P��D���3�'DӒ?"L�aLa3�'XL;�10�����hJ8�X��IOI�Z�~����4S�}�Ĉ�����	B^$Æ;'���Q�DDD�DM
B�tO��;����"a1&[�|��D��+�'4"b"I�lMDM�#��DNi"#�
�%�r���E�"t���v$M�	i:"q�0�L'�N&�"'8�5�5�,�9�':�#0�h�$D�$D�h�4W�DN"#�t��hX����0�4?m0��Dp���پ$D�}ӣE�?lH��""t� ��z��1'3
l�7xM�Bq�p���8R&��8KJ&��V���Ė&$����I�bq�lЖM��hϨ�	��8����a��Ʌ"&�H�q$���<���%D�tFL7S�9��7"S��g�9��Q����7��ު&�Sbn�^ԡ�;&�D�g&��al�fh�U�D{ ���\jY*i>�br��6w���G�0rLn�}�IQ�T�6��N�S�r��+z�ZJ9C�+�'�>�ݚ�����<�\؏l�C�Y�7E؊�t�ꞝ��`��gxγ��8�Z�����&�p�����a����Q2�m��d��!�D�їQ�LD�'��nj&�sxh�bg%C�����;֦�2ac�DG�n�(J�R�lM�Y(N36�J�D[��4Ϡ����b&��}F�O��TDrAژ#���y>Dd��WQ�K|���Dl�bY�}KЈ�j'M�J���b%�Ɖ"#��t���a'DvH������DG������oyQ3'zt���t�5R�uueD藹
�D�؉f���D ��2�a���D��54v��� �"X�:t��"fN���!���K7q�ȝw!C�{,� �����5�)�4h�vQ]&�A�c؎G$i+��TL������Y��(��iE[Sd���M��%?N�5MJ&�_H�'bg
&D�N�}�T��>F���=���l�&抣���֪#��i�J�#�܉�۩�;)�%h�|�J������S%$�N�Hs�U5(J���+�*��e�c"9>g>�>�1�|��C�TٮM��ԡ��Fr�;Q::ʈȏ��II�Ȉ�����Kw(���|��Ȏ����>O�}�\-EZ����_�՚j�l��'~d�̟k'��A�Kb��#�L�������Y�Z����/�����>}��i��_���ًe�p���:lW��w���$��I	5RH74<�=��L�J�4N��s�/���=�N�s�JފN�-!�'S'l���n�r��sO'&�N�r���3�w��۳F{.�GML��jU�yځϋ��*F��j<���Y2QZ����ǜ��v��фdbUɹ�jw�3�R�V5��5��eq�8ʾ�Y��O3�q�1�;�ϙޝߙ��g����$�O�U�G����z5�J�-�W4rғ.gZ�I:�WɭM����%�=���-v���x�\�E��=:wZ��'�~�����'���~�$K�{8����+�+�͓��W�%�${:��I9����p�:&t�Y��:"�+"QO�`�D��H�������r�A��J{)�,N���:�_?u�f�SPD�$D�I6A�Dy-ep4u�%��+�r%~��Q�%}�D~�5�JDy䯟�R�&��D�H��\4V�${)9BsL��:��K4?2�#�DؚD{�ϡ�j"Sr�8���L�74?9)Gu,M"&�"tѶQ@�"P�"p�8Q��8:쯟�U�4��'��ǒ�Bk�`5(n"p~DL�N	|�"N�M�R�M�"&�S�'ø�Bu�F�`�����|�D�T���dd��%�W�~�ډ*���fNdN���òp��r�����/"t�Y\�/��&Ʀ�H���\��ᬉ�eh�t8H\�]Dp~r��|�__�j�����,K�e"�1��[��d��ɭ�I��K�w��9��$֥�愷�]��F�T��'G*�0rIӌ��Kd+q��r#S�ȎD�]j��U:�9��`���:&\K�d��Hw�jt��㽭�ޞ�Msn�oM����/�	�%�9� �YTWj��Rps�)�n}�ϱ������չ��u��_1Z<�<���8�y�~uoʝ,�ڻ����y)��ƪ��\�)ɶMIs{�̹��#��$�SrjK�'\����9�78T����ly��s'�>5w~ohlm��>c�T_a������9�rxmO ��/պ�[k���u�j��h�Q3rQ��%���N�".t�w�0�۝�Nɉ�d�f��KvNhN�'4or�&�N��$2�K;El+ED���Ι�:<)�5�X&�&a,ƈ�9�ϋ/{�w��+s�Ae�D�� �����v�u�oa�}wZ�N����t��xH���a �5��T'�s���3[ב��o�+Ο����{6a5w�:��5O��g[���aӹpd�d�b%�z{��;|iӝޏ�4�>��L�{{��]7��}/�v�Ӷ�#G��3'sK�T0Y'j�W���vr?_j�u?i~�w��vo3g������N����<���ޞ3z��n}�	I��;w^���a��G�{>����+KpL����}�g�S��?e<M({�.�3\��ݽ�ᗤ�w#�f`{��e}�����>�{�̒vN���N�*����d�ϻҙ��`�j���� �Lf����;��W;�f����ӽ]���{�6�Z[t]�v�N�ώ=r|����R��$f�������6��w�{���>��|�ק�^��꟬ֿ0ɯ�wXǬ�����M�gԪ�}_�nx�Y��6��
�ϴ|v�o�����7�z[�}�Ռ]T~{;�w43w�z��>�^IzC��I��ЇzE���k�cy�>@�~��}���}���0�����z�;�\�0O��U��}�����M������V��v��������<�a��=}}��٪?���Ȼ������'��u��}�~�m�S����P��rfx����$��Bz-�f}\����ci���1���)��svug��g�+���7W�^lͺ7{� ~|�o�[�Ɵ^aG߽��}=@˛a.;��4�9���Z2���i}ٞ��ǂ����0s~�O����Yruw�u������0�� ���߲\X�?���4�v|\7�ǫϭ�/Z9��n�Y�N�AuF�abr7|b�׽��7�:���7ӳz�A�����ƾ���0��i�dx�Q�����?l�إ�H�S����v�~x����b�( �� ����,�wᛎ��a�;����N�25�תa�~%3oӕ7�:�c9�8��߷���N�X#�{����_��;+�KL]�j�R����j��#��L�-
}w;����q���ky�(��My�V��=�s���Y7Rp��M�p�DY	}{}���������͚tU&�����O�c��k�]��Zk��f\C��~<���&L��f��[��[y׻{�2���Y��~(0��Ϻj"�k�O��$e���*��j�ۋ�;4��cݯ��>�f�|���v<[���d^��=ty~�V��E�>�ϕ_g'����_������s�ןl[[�,�n޶4�rO��,���3�X�? ���1LR�ߟO�x���gǵ'�o��?����>����x��5]y�ޣ�+�e2w.�\���Ӻ}����{�v�ӫ����W��/�s�~�`����71L�r�v�͋1��'ݪhgj�Ϻ���RW���Y|�nh�c�\2�]�m�{�C��׺��k���=ft�������=��{$�ٟ/t��i�e�7H�\������}��1c��N���k�{&}����w�Gy~�w�����5Rw�[�����F����׹��hirv0�9w�e�M_+W$��ž�;���_\fjn����k;�l���ឣ>����Tϻ���I��zo�ս�V���~ݿ3=��{��������f�y����{�1��=�_t�~k:��e�0��M��!�S��1��YV�Cq�9Oz��s���}�A��yJ1����Zz������33�4u�s�㣽�I�ر�'����N��g��u{�j���,�h���]y��<֦Mni�lNc����I2]y��z���p�,}����f��͛��;��_O���<�]������3ڛh��=&O�)�9�Z�X�	�X���b�S|ߞy��g����t��	�_Y!	��6'�ՙŢ�w�/c!5��x[*����G9��N�[�{��{��{��}���s�9�vn�}'���d��=���C�˒��vE����>�??�
�����N���7�ߡ����'|�q�G���W��vI%��m����˔~�o�.zy�+z�����߽��pat_7}�v������ۜ+����7;���߯nd�q�3�(��T�;ܒvcݝ��3�烳����w��x��8��ݓ��}�57�7�\�ot=��ޝ�´K�lû��:�Z�ח5��C/`�m3d��s;�w�&��Ϧ�q�BoG�^��/^�۳�kY\���Y�s�g��YU�Qu�j�zY�g�t�>�>:�t����M��Gd����z�S�C4ҧ���5�cx�'���睏�&��{!�<�����d'���S��^���=k��﷿�,��������������7��{��k��t=ٛ��� +�5eי�۟��g�:��d�Y��љ���OBXK�}1[��R�~͂�7�mެ���ի��y?=6��é���F���r����~{�3�gnN�eow�l׋l��޶�܄j��7y�Í|{t��7p�{��|8�=Xp=�O��s���t�}"���v���Zx�١zN�gF�lUl	�W����f�~�v�ɋ3�0{�f��ɘv�B�}.5&�c�73�Q���w�\`�w\7���o��w�lע�^�:�%=�u�UW�{�ֲ�^�O�{�M5�r�!ʄ~����Ͻ6������M�����K���y��T�(����E^]�ޞ�ʜ�dV`��������|�fjŪ��-0x[>��w�m���3��Zw>ƻ�ۄN�V�f���3�l�Tե�Y��dצ^�V��_��������|I���X��E�ޛ�~�L �N�/kX��s����e��/�٦��$�w��I��A�I'ow�U��ܞ���v�t��ݽ�$��sf����'��?G{>x�sQ=w$�w	�4Rn\x<مS)���=X%��_<�n�ڧ?^�~?gwL/'�r�|���d��y�v����Kwy,�ָ��P�����C����Q���D�u��vNa#�� e;N�n�80N�7I��:'N|�V�{���lS@���#A�B9$$�8E!+U��'
��k��+\�fA<,�Q�%�%S�:�8�Q�ڄ1I+�:����x�'Z�Y�Sr�c�uZ�٢��|r�P���-��)cV��H�*ㄱc$�ڱ�q�XIW�񨭚'��.�,�ʡl�|�dr0j�:4���u4iY/2Ե�ۘ�.�KU����!�\Xک��Ӯ�d��
�r���v�.T&A�u��Ö1�l���d��څre%��&b�(ՊҴ)x�#(>�Q}3���Ǹ஭G֫�XE�����k��$�3eM���eq8�e�b�b�I�aY����V��lQ�
lE����6i�6��*b1��uA���D�r&���n���ջ�FK��,MX�h+Q�S�أr ���V�X��*9Nj�8BJ�!F���ƥ�!��eFi�V8�|����E$�D�V��ك�!�l,M�,)e��%�#�DN���B���1#���-hRDڭRT���Vڄ(䎄t�9[[*&9��6�B�D�Q2�>>B�X�U�)[RV��[FȡJB:�nQ���ʇ���ydP���Q1���V65��1�BKG9��يQ�c�h���
L�I3�\��F�q����t�6�H�Y�8�X��l�,T�v��{�z8xq����Y���V#����̕���u���QX��6�YD�Y\8r��#U؛1�۴R�E���m���#��X��Ɠ���'�����	�Tz��2D��4�B�g�x Uc�	֊����޺tc@�1j�=�#����Q`�pm)"r�d�v�N�i�����,�*%��&6c�8"�*���䥟5���4�ylR���6>�1�̶'ȋ�[����,���0y�<)#�_�<ol�g�ƫ� ���s\��K���d�Z�N+D�gwtzD��,��T*j�+T�(�8��J�ɝ���qΕLM��蟻�td�ڬD-RTfֵ���3�f�}��[��Z�pxOv��5�UPW��P���f�W�>�F���r�L}a��s�Gr2"I@���-~���ߛ��UUQUUQUUQUU�*��iUU�*��*���UW���Vخ�V�v��U⴪�V+�kJ�������UW�Uz�UW*���U\X�}'�} }�� �*Tj�AZ����
��"�BH*Ȳ(H*|}!���U�+�U⴪�U�UgV*���������UW*��*��*��*���U^�*��*�UmWN��*�U\V�UꫵV�]����U⫵V�]���GĀ�R@d�@$Q�T�����ZH�x#Q/J���}!���R�t����Wj���UmUګjҪ�W�]*�WJ��]*�t��UҪ�ZUW�������U�Uw���j��[U[Uڪ�V�Uz���Ҫ�V�U�Y��  )�PC�'��{�崙U�Ҫ�V�Uz���Ҫڮ�V�v��Ҫڮ�b�Ҫ�WJ��[V�U��U\EUUEW{���UU�Ҫ��UUTUUTUUTUUTUUq�}�d>
�U�Ĉ"H(�"�T@�J
H0Y mdRI) (;�%��
H¥(H� 2=g_��|�
�0!d����=_BP;�y�x�<N��B��:"`�&	�0DDç��B&�DDD�H �M�b$D薓xM�Y�4A�(DD��8P�#R"lDD�0DD��؛f�Д%	Dd�2h��Dؚ0B�Nd6hMO�t�""pDL�DJ�N��"`�,K6QЂ �	��F�M�������^a�WO������Q�!��tj�XWmn�4Gr�튽�z��u�$���i�Vۉ#)��c��1��U���R�%���e�䂊����
Z������霞jV���@�Lw�s��ba !7-ԮrTZ_�#O"&5��!׃	Ud�"-n�Em8�@��uئJ�i�S�EQڜm[$`W�+J��-��c��r"J��j�r$^��٬��k@�H�X�q�-��2BDNE$+�&�'����FrI��b��*��av_�V!���?�Z�"�kr]-e%j�|8��lUܸ\1�FԹb]��p���r�\Ņ���Za�ф`�!]����lj)�ȟ�C�HJ��TV	�%�N�an4Uj�:�$v�[*Q���9*5$ض<��x��lP��%�B�9Fz,2��r
q�UD�k��%䶴�jX(�@�N%Y!tV�ʯo/s]5^>%�-WȪ�wwj���'��{���U[���}��������{��wwv������{���U[���}�����P}�:t�<u�un-Ӯ#��m�������x��$n��]���$b0�q�PدN��"vT�rES���aek*�M|�dF���"g2E�X*Z�q:W8�rr��8KK�� ��5,�H�i.��B6_�݄���a)#7�)��S��$3�p�4Q
�n�.��}�Þ:Y��WI��tg'�t<�:<b���v���j�x��Ht�&�WMݪ�.ĸG�j4��P �[����W�/Q�3$��g��S������[��o�[�qn�um�o5���iIoVt��s�������B�J,�P�����W���4k�U�aȱgGۡ7Bn�ͲrF&���9B~�%�ڕX�3���l�c��T�q���QLUB�Ð�z���o}�im�u��x!��.���l�Mp�����'�U-9����4p�Ӆ����Q��6�Usq�)��U�uJUT��m���M�և�23pafl����FǦ͒�Tp��g�� jQ��z�mn�� ���.�Sی�Q2��ں}ޤ�lF� {�eGf�����v��d��w#m�M�.��I�変��8�C&L�8���V��:�8���I�j�������G'"wb<B�13�������E 4E#�Χa(�mc�b۹FW��ϳ�<�+��+�P�F�Hu�)�MM�<C#�l�hҥ�6T�.����B,�p�ݭ��`&��Yz��:���6�:�V��[�]GQj~����8N�Yy�DE�2�U��i�C��UW�91�h�k�J���"��fs���.��fnb� ����0E19�Kj,V�T����K
���㢜�4�Ա,��LV�r@�vKU!h��ڢ��!� �<�>^�����
917���8h�­l�8Y2a7�)�8{fĜ���x��xU=I��*����<���w~���s�Tnn���h��bڐ����G�mM��y�g��l��X4M�Bjt�L9q�؛1��6ێ�պ���Q��7[��M"(S*5�U��z(񳫃,�߇�!(srh�an��X�Z����^1䦩��fry'gLs4曶c���������<���#ܥ�J��ʶ\�r�^�Κ*�iY�x=9F��FX��b(�QI}��TZ�0t�F��8a��:&C�#/tJ���V�iUf�ocpBp]�;6l,�YI8��I6���'J2t��7m�p���{YF�H]х�蛻;�v�4�5'5-S�N/�����*pwS$0jfT�g,��n�tp؈��9\4n����y�0�{Xr�"I7Qխm��V��[�t��]Z������@*�T�S�[Ne�w*�*l:6%�%51;����G �K#��]����ڌ��)g&�{sp0�c��Ś%᲍B�pe�b��æ�ʂi�ɂ��k�������*�`����n�[�[[�qn�um�o��q�������[�ȁQ��c��F�l��{�M�g_&y�	���B��'+��Dj�t�����&����6���#N(�oZ����x 8�sUH0@��%+��n4�X#�U��N-�hW���|�!.-.�*�I�F��A��xQC�:'��"�b$� �4Q��;=;��gE�fsWQ1��/���Q�Tj�Gr�=�X�6XZ���2++��Vڪ4(Z�v�ct5��\/UD�d�a��Eji7Z����:㎺�V��[�]GV��cy���_	=�S&p!��#�Y�f��UVv�o�s�{UwE؝���3��YSj�EI�&<�`!�gPay	c:�4f�Ӧ��'ac���
��-�c�:�7bBl8�yR�`å��VfvbrͰ�fjr�*��xTj�T��ڠف2="�ӈ�u6���c֝���bZb�bZb[�[��q��4����cX�_�>k�|�&'ε���|�O��cֱ1�X�F-��b|�o-#��6��~G���+O�|�M-�m�cY�5��Ķ6��a111�bcmbbb��[�[Lq�ɍm1�U��1���k����x�Z}M���llb>LI$�Df�b?1���Dg$�`���hr8=K��=S¼Y^O�k��<�q-�m�Lj1�Lx�3S���5&"��ԛc[#j�S���OZ���<	�$��6���bz�z�zƫ��<Q��ѯ�\}��j�T��/�sH& C?[�ߡ����w�o���,7=z�����u��~Kr����Ww��=$7�`�.����FJԘY��oW�3�~�}�=V{}���0|�u	�b5nc�=�����1u��ߺ�f}}>�_��U�1��U������}�{޿{=�ޞ��������W��{���z{���{گ��k3333/2ff~��}��m�q�X�V��[�E�z��?d�M9�UV��R��J�'(��Pl!߽��QwX�8�M	20�ɱ����=a,C�C�����-0Ք}�ڍU�=�\���bsg0�P�����4&>��J��V�g�g52�E�-	f�xZ ��ĸ|H�8T��}n&&�XC�(d4&����-�$͛�3ߢ�����M��Q��� �#]��W���L����҇ԋ�����%CpL�7ڶ���rD
���UWH��?W�1믘�lq�m����z�~�$�kU7�j���PD*>C���A���HZ-�v��!����`��\ʸ펒�����T��c���r+9ŨÐ`z0����BHy�"xMmh�0�g�������(0(�������8NR��
Q������A'�
|�K�EC�!�>����2T�d���3�A�L�]�7��3�T�%�(��(D�OuvXC�4$5B�3�N�Փ&gU.�!6�-��-��V��[��Z/(���!y��92Iǔk��= ��N�M�bhŌ��"ǅm�㵋��l�\�y�Ź�UY"�.7���Y̎m���s3�u����f��JG��Gi$v��vH`��v0tAﱶ�m�ҹ�괵��J��L��\��[WFL�q<J��>L�!~Q
20D���0�L���4��X$�����	�0m"ϧ� 3P�BA���,U�!Q'�*M��2��d@����B���V��OCQ5؆�4�V���JtA�&,�����
�
K:2�bf!��2K��,=�>d�
���}�Q�?�?H��'\(W|��X���bn��	Q4BR�,B�A��(�n�31��n�d��0'��E~~|�l|žun�źu�'K8a�I���)�8�i�51UU��7�n@��C�Xe K�z!la��Y��DJ��7.��xd� ���В�8��C	������7cw�j
����9%91�T��rJ�II.kM�Y'��'j@���}U�ꩢ��D�TD��_#PD��*1��x��.��9��\�"�(Uj�vr�\�AVWQ6R�rD/
 ��(��$N���Y*���w�-s2�Wj��$$F�V&i�n�r�4B�	(7��8�!wsV��5*�����t�ǋ|�n�žuk[�t�i�=���<מi(�"�Z�/�UU�WĪ�����B�R��b��tH},�]ni�� �<��&��%�ƒ�Ӥ�,j���&�Wi�,��hL	>�U*���+�ĵ	g��ƛ���,D�Yc��$aLh�<&e�=�N�虈0d:0��	įgdĘ�00�Q����a��(ZnQP.Q5X����-V���;����nd
Z �T.�(lړ^�H�����2�7%�T�q�����E���$=�.\��992n��Z���:��q�מ��癪x�r��%8��0�.={z�j�!ځS$�_�%�9?V]��Qȇ�pap�"Py�c'�h�%�U�ֈ�l��YKyq-�v)�tebduDb��m�Dr�Ԕn���T&�r!=� �4�*Ii�qV'e�a�*Ƌ�	P���<᥸L}J$�1�
�HX!p.�؋�b��Z�ij�P�$��X�i��l
���C��Ua40�J.$����K�(.�t`pKf,I��3�e�`��&�K42�b�1�b�:��źu�4늪��5�o�;dN��DMjZ5e�E+NZ�G��b8�r�lo�5�&�!z���e:�)a��NX��h��@����5e�dQF�
'��|�#,p���m��Jfn�%���r����x��do$j[�������)o��NA�D:r̭P`[P9�cF���M�0ɫyMÈLND�5���!�j�*���M�(�)FdOOb�p���D��c��2��d1�MO��f��M�<h�1I�	�+��Ip�*ƀ5D6j������S���	��d�'%�|2��Kd�
� ����~���LA�};1n[��q��S�HՐ�\�2�.�b]]}�/�Y��*T�&�����̌ܲ��N:��m�>uk[�t�i��4��m�"'<�V;$P��~��m���(s�92`e�>�U�<z!�IA���'8�c*�5�Q�p�7i.C�.H���b]�G2�����bF�"��1&��#�)R%Ȧn���,ذ�bda�&�=���q]ĞLnG	�X�.�7vh�"`�u����YaT!2Au6�1(bc^2n�t]�I����9	8��`�@�D.|T�0;7(�9�uMU��!bn'(X�v����M	�j!��FqE��˛������r!2'g%*S����8�c��Z���:��8af�Ԅ������h�G�A9"ܹ2�.�/E9`���$�� �x�:ɡ���L�z����~�(�dȉ%FO%�:YB!��� haF�G�I�
�y��qB��l�/��jQh��^lRy)�#��P���[��ݭ6RR�&d���[��hC�m�z�=
��L62L��VU���ahj��3"�KYp՘�Ε0A���ꢵ�3�r�y䆏��#lu��8�1խ��áӤ=:p��_KR�L��a/2�R��P���UU�}uaP`wgE��k�d�~I.NC���J�Eʌ�4v`�Fq��(A��gʖ��%�ȹ5F&�TZp��8��1���
(�������3�M �8��3R�d9�dd=�!�C�|�MXm�"Q�h)p��T��Q112_��.���FN����RR+T��������E�#�� b^�](�	��]FW�4r	 �G��8��u-+�>x��L[L[��LcO�i�lk�է\i������i�������bi4Ƙ�cLG�k��5�LKcU���X�q�i��G�5�>x��5�}��>O����x������LLLO�&6�&'X�"���c�m16��H���?5^��S�x��	��J_���(��DO�W�U>�T����<(�<Vň��F&�i�=LG���+�u1�5���b������&�bF5���Ʊ6Ʊ1m1-1���M��	����D�W��
l���c&$G�z�&%bz�z�zƘ3#�0x��k�U��]�[Op�F��IVI�S�6����+�4��su�a�{����K��Ӭ��B���Xck�r��lX��k��f.�!�-olS3v�9�.9��yϼ�{��0�:�B����y��^��h����fV��*� �:��8��ٔ�O+�ϵ/g{~�&���U��A}Mq�(W�g���3ڭ�<�4��Q��c)N�����(�ۋ�&J��&a$�1>�-��=��3cV���ݓ*r��gK���9��mnd
0x�j���Xc�G�\�P˃,MWr���3^�r�W��P�\��Գr��1d�gMZ�m1E0Zn��l�~s�Q�۪���ń���W��bu�&�>��'M2�8,x(�{{c�����;�k�S]׊|t���~>���sa�87���N���D4X>��]YY
3I��361�ٕŞjC��n�˅� �����AI$�Ii9*Pr7%Q�JT�t �n�LRV�PUR�Yب��oH�ǤXW0Pm�I*�#�*�ګZW2��4�,(�GH�$c�qEc��Y#*�U�dv&��D�i��TD�)N@ٜ�q�]�27�"8Ԫ&�p�J��q0e�E8"Kp�ܞ�j��)|�`�E���,R,��Z�������י�.�Y����}���g��{��V/��]�~���������uZW�������UW�Ҿ�.���d:p�Ӯ8�1խn-Ӯ��q�w��xP�rW�Y�!ȉY-�ӗ�����Kc�n��8�u�H���Ym�(f��_^#b+D�@�B;��\
�QX227c�|��m�%���Z`�Tt�-�S0h�Uf��bo�LC��C���nl�"2^��lvv���"lg#%}1�qP2%|T��>�����U���N(aە%�|C���D�f&
��eCp�E��C%@�M��{�3�(�@	�}���K��1g%�vT,a1�2����s$0!�y�O�8pL��4̊��{E����(�
<�t&�쐍zD���2+I+��>��4�M����[�X���C�Hp��:��˅���qUUH1K%��i.��LGd��rQ�}iZq���*�XPЛ$�*`�j�5����>�,3��A��C�=
�*!����i���[��t�ה���C��h֩(�Bꮌ%@���o�2��0p����^f�)�cW]����d��R�6T#3P�=��]��!�c���;0#*!�`p�
�>>��c:h�m�EFVǅ��!�=�ӡ�qo���-��kqn�	���H-�VJ�C�n��UT�x@,�_PSW�;E��P�Q��6Qe�Y@Y�ܞ��'x�%U.q�(@J�|b��Ѫ	P�,������	�uc]TP�:;�X�i��]��������n(�G%8NS!�K%��pkG�����)��T�$�]͌36Pˇ�w��P�^%�W�Ѡ�v�U)��cS듦l�V��4=X�'��}��sҴ��qrB�C{�5
Q��)�T��~J��q��������-��áӤ8zpü񪞷i7犪�����������IQ�g���+�tؠ����@j�!��]�Nj"�r�B��Y ���p�H��C��(a;�c�3B�LX��ͱ4Z�Hv6\*�\����`1�T�b���W!�$FJd�v��{��8����qUGS0��Qaa�˕Ũpa��{�)��L��0r����EL�I�,��!�Fp��b;e:�J���јT2h��h@�£9_�T�U�+�*���[�[�-�'D��t��fYz���HCR�[W�H�ݪ�AUt������qڈGk���7��yH�M�>T�B
�D9$-���c��J���{u�2�Q�I�ZV�M'!#�GZ�� T�*�*���5"e�#]�����݉0��*X��>(�e^e�f*�.�.@���qf��9q��UB0���'%NL�"�׍�o�����332PZ�Mnbe����C�����SE`�5J�/�;���Y��\A��_zN�� M�����r��o5m.�\�W�5W	UP#G��)L~�Hv$ �T�)(l;���EkQ&�����q%\$�ƍ��!to)��ӕ6,:)­���ו�:��|Ÿ��lc�Μg��>�ο%<qWe&.��@2�Ic������T��kF���ac$�� j� ���f���r!p�`���0miXy)X�gC�=��0�.&��VhQMf���כ�>c���fJa��5NK�J�S�C	Tw}�7�7�� �3q�eT��0B%w�NN�&���X�b��RD���n�\�����_:��u���1źu�q��x緯	+�޴��@&�h����3��rV^8]}Z<�e�����e��D�`�pQ�\�tѲ\(SAȆ�!�Y�(0����0:o�s��]ݍ�mV)Ur98�
��(��F�.�\�]͗g���o�N9ӧc�U[.zk�������*�(ؔ�*�K�nrC	�	YL�0;�<�����913��hу�w�SWQO�~c��>q�|�1�1Ӈ٢�	��iA8�%���n�ur��Inf����� �[��j۳s�&���K0������0	�_[�?Z+��n�6̍\%�.�1f1x�\����.�6sdJ�Q������!�3p�e�0l�g��h�rM�ѓ�-j��a���p���Q�s"�H�
���ʰ�2#�(�IBSѣ&�*rW'P2t=	���nb8\䳢cE�8d���>|�1�1Ӯ���cw�ߵ��yB+B!� ��)�L��(��_��1�F�Ә�aS�k#���L�K�HEL�lYaSr�Ԕ�o�1��D�'�(�o�:�T�h*��Kj�l/%)
q��x�-󪪪@�{ܖ�q����2`�2}=�-W�MM���drbO�����ͩ�4t�,��nQ��d� 0j=�d,16�ZKfq,٣�B�4!�1Q��GM�a0�P�!�¬9���٘�rrޗna���bvb`���Gդ�������QoJ��Y�מ1�֟�����[l[��qձlcc�]GxǙɽ~�׺�����)!�n+3.HZB@�\�����V{�4��+�;�!���MC�,ѣ%�/�QX$,�0�Y}12T2���td31.��g�F��.�5};0h>>-wCwe�xj-�yK�	lx"K��l5UB]��}��SV�Q���y�v���\Ԙ4��v#�W����a�&���%]��q6��ih�--�Śb�Ĵb[�bD�4�5�l[Χ�5�k�5�������i�4�b1��1��i����&:�Q�lih�bV#i��?&&��Lk�i1#�ǌy����ɬb5i��i0�Ʊ<|��#���K|�ȷ�1m1֛LoRc&��4W����'���؞,�K⇋E�W�A��|*����S����DLM�ӭ5X���(��~Sⓥt~_���^k���4��HƱ���5������f���Ŵ�I���?'��&jTa$�Ĉ�1"�&&4��x�&#Ԭz�zƘ�ɉ^�i�=>湒o>����޽б�aqڰH��1���<ߦA����)���}�O�Q7w�{$�{�u�E����{�|����d�y�#��_oWsbٙ�����s�e��|���8j��ls���'5Ǣ﷞{.rT�������w������uZV���{���*��oܻ�{���*��oܻ�{���*�t��r���Ν8p�Ӎ��1lcc�]Gxӑ%I�^*���[��z?9N�4XyI��J>ݫ�xY�8�.�6}䎫a��<f&&f|}F���suV��q�����Uˊ�����n�}���NO�O��W�9KN����7�gaP���r37(�^�ݷkWs3%�,��(�&�(�3�>���,��h�Դ�jr��Lp��k[�͸�ϖ�1�:u�q��<�s�̽nq��|�_,��L�UUHirI׮��Ć�6|�#u�q���vɔy��X �K�^��o0�(lqCU(�����p�ՆB��O�bCr��i�r{��e��(����>� ��wE��A�xQa�<�k�`���4�mX2��놈�����n����e~zGZ}Ԟ�D"��t�M�{(�+��[��>q�Vű�u��um���M~Fޏ�E�K��*m��('�,�!�ŕ�����Kb�#�c��5����[פ���"����U��lF7�`�ˣ((��"@�	��=+�r�paInLQ:�����M�(),$����B�2!��K��K�a�/�UU l�M����!�1HX�[*��CWں��x,Y�*�.�>=��|2�152zZ���l*��J;�EK�C'8*�ݜ	���R7eܚ�*�.>4v����7,ѣ"%A.�q}K��a���F{�ǣ-eJ��}�ÁP/U>=2}l��@��|�ݮ�aLymᙙ[0r��%IS�7�A�x���]��p�Õ��Z�I�F�n�W�&˯�u�|�c[�X�֎��"I%��D�����UT�ׅ�]=��
���L���isfa�=5�S�j�͙p֕F�}(�x٬��umWkgL8J���AA$�һ�>�˓����2��U`R6B�
!��&Q��U��U~��p���5sk*�B�u����h�т��y�5T�j����S��Ӕ���Q����8��u�cb�Z:���f�ɾ��{�d��r�H��ꪪ�:k���w����j��2l��zvj\5F���~��\�n�0.�H'�O�	vXvw�z>�4Cw� ���(*�U�%w3"�,���v��&ga��u>Љ�:v�HmYGHpD���	�F���[>���^��g���X(�.˞��l��̢�0�"�\2fnD��j!�����Lm�Ϝulu�ca���8h��-n��T-<Ʉ�.<窪�@�	]�I8x}�5B�����:\}F �L�K�&J��D[-���g��_�(���T9��UHY��F�?`��*�3B�aAӧ>c���A���kY��)0dC�Ie���?Q��MB墢�;,�JJ~ﯩ��Ju�V�m��_��8�>[�:Ŗ�u���#&��Z�yYF��J�����&
7ݕ�U�y�L9�qa����@v6�C���Q�\	grcY�%dQ6+	b�ؤ�(*��7jy�9ėw�v��UUHM.�%إ]�b-�M�;R�8r�[���.x��`��Bm�=��ʳ�6
�辶Y�rP�&0O�D�<^�cLЙ(;>��M3��\���VU�L��&,>.x'�Y�sx�1&��P.�Y$�TB[Um��Q�����&[�~T�NW����n�!�>�����J~[��Ͷ���uo��1��e�m��TJy�S���Ns�UU w�a��Jʲ�FM�M-I��񉭼Ѱ�8T:6y&���}DFC��]"��d���2n	�7!����>⪍C�\��QWo"�� ��7B����q[�&d�-Aqn�b�l��4nbWLɁ�O�U&K2tϗ&fa�у�C�ῗFD�,�{M����rI���ǯ�[��b�Ǐ<t:tN,�!���]�Q��j��$=�讍r������_�М�I�\�J$�;�CP�4"dD��F��CE�ȕC6p%�3�C����I"*0��H[�K��ao_*�j������#cwue�D�Z�����fgh�L�&89S&eϯ{�`ё.Iv�w+�N9r!�nXr�p���ru62nu�>|�c�]:�8��7������$B�U �e�Ld�'�z�.�%��bc~���z	�wRdM��=���P�w�I�Kl�a3-�n>
HH��)�uR��������J 6|��f%O�5[��8%	읅�3,D�a*�L(�PY�e%3�O*Y��)�b=���M�xl�2h�((N�=��KUJ�j�!��:@����.F鲼�l~E�ю��%���i1mbZ1-�Z1-�-11��ŵi��0�cX�bi�����������X�X��#��ZĬu�Q�lii�5X��4��?&'��1=J�bF5�k�5����������XcX����c�Jŵ��5�h���V'������G��c�0�����=�G�
(|4U)�U<'��\>"�h�4��O��5M�i��Q�rY^�]�������|p���zƢbcL�cX��&&'ש�li�Ԙ��q�ɍm+�x�F�eI+#ĉ��b#M2OypW���xh�	�EO	g��=^�ߏڴZM��*�k�`Q{�߲�7y(Ln։ �e�}6\�m�F�̮@��p/En<dC��]oq'����#���Y��f)�՛����S���œ�'ѽ��/{b�s�W�\�ztܢ�E�N��^���`7�N��u�+���^tY&;k1�PZ����fe@�H���Z�ӶN���x�}�֦���~�LI�}U���2I=��vn��qC���~P,��횦���]�������=ٟdݍ�����.�՛8F��-�w��˹6>��|{�=���w��͉z��5��w�����6�3�t�j���e�K�:�>�o��f^d�����<>�!�MՃPF���u_+��O��1}��r�F�5�"Ț��w���x�"�X����������n�!����G�r�ݜOtr�|�zE>����b�,7X�܆?d�<U����N�>����/�y%��q�UTU����-��"�I����Q��i���e䗅j�a#	S��v+ϞD�S�NfC�6�rFW%M�5AK#�UF� �6�C(�Q�̫%b��݁%R7d���RG�K%@
��]�02)S#�"��V���ܔ#8 ��q8W_�E�f]X��PhN"�V��R��?�[;����߷�t���.��{�]������.��{��V�t�~�߽�{�v�ګ�������m��8�c�-��u�q��b/�ë��N�����phJ4�TX�m9-��`+�*�2���@�Ɯ�Lv��|���i�4C��E���	��*�X�dd��S���H'N ��
&$L�m��|h[���l*
�P����b��P���6`�"&'�ȅd�臋4&DD�
|=�&��V{���ϹE�SЩ��&���M`��nX�2\��Jd����S�8p�6|x�Ul�p}����2wpa�Y��А���Yx���̒L�YD�*��\l�Kk�)�W�+�kG���l4C�A�O�nۚ�[���z���n-ŭ�c�]:t��p�����%�=UUi!�OY���fp.��qM�Z��;7�'�C�N	�T�p����ylXRz��w��Ř�:lD��Uv>�3q*ԭdi���lMd���l�r�CE�~�|�cs�drd[��>��
V^9�\��-Z���	�a�Su�3�Yߖ�}&����M�
�06�.k�kڔ��6�믜bض1�uӮ��� ��T2�.QQ5�*���`�=(���e���*T��`LC0IH`�▖���ѹ�!f�ؘ�s)4jjk��ɒ��'��!ƒ�Hy�P�y�O�b.WeZ���8Μ2�lǋ6'a�S8:��z,~<lٸQBg �ҡ��lf�"u�Of,�3BCF�e5E���6��&��#�OFh�s����:�������-�N��6Y�{(&���$VuUU���E(g���Nό�9>������>��2r0�G�&;�ES�����G=���ĽϕG�O�;�f�L�2"�����AK�X5�[X�&�����p��Ĉ�>�,��Ņ"q37~јpM�_���2��*o��eWs�a�,J,�9�)}�՝`PDN:|y�>|ű�[��um�5ri�񣭒0]�E]�F����=[��o��\�P���u���Z���H����y�(D#�L��8�GY�1�6ptu���r(��U��Z�GJ�c�
�⨬w�����m���Ә���[-��b0˂�lSE5:v}�f�E�B9�p�ag~<�;�lЈ��i�H7;>�����	z��/&D��{+�ܶ6ߴ�>��
�+����ڱ>�x�1��@��&DD�K7��^®m�����b	�nt����P�B��?ۃ-IVY�����˶!5�CSԊEE��U��p��XA��JV"��V�.�<]{������8�ϖ�1�ӡӤ8l��p���4�˗�UV����0����!)��#�0�GG�<zdK4�-�t��9:6'j���.-6d�P�=V$�d���l���*�"��e����Q��ȅC���UQ��0���^4YИ0lDM�}ӋT~�}�-�e�!��!��9Z�D��B�\���m��ߍT,����[�1l[�]t��o�L�䬚R� ��*����U�Tp�=����Q���E1&��qC3��=��(��ʪ�ѓ0�Q��>��"�'���m��]�Ԓ�9yy1����z�*�9F�	����L ���}��X°���TP�#�*�b"'��	���=��;T��k��{���u[,Kk�E�����fa�Q�ƍ�qŭ�c뮝um�^��^{�fk2��x���B�O��T":op�>��Y��;,�1�9�0��v����DV���c�z�yL\0pɑ2& �>�c�P��;(D�a鳐��=���s����,O��.b]�ͫ_Cʜ	�Q�,�L�q6&��9��A��h�;(�<i�n���cN-o�[>[�y//!uj��_8�u��Oَ9DBL��ae(�Γ)�-����� ,[,�`CM�3�$�}����b�Y���"��u�*�2�-��L�	w*���Qmv�^>������{q���r�uEd���m�9rEy�%�|u�+�>�X�ӒF��T�V��Ѣ�.%�ݝ�NS�Kbr��'lߝ���b&�|\>5>���+�r��}�r<�)���ڨ�'У"b���%N��%N(��?H��`�A��N@L��QA�a�9��G�#3q���cMLT��j�ʛ�h��|�lZ�-�[��:C�p�c�G��#=م�8�%V���3�/C��5�Q�.^����&��'a��'~`�M%�hD�0�'8��+��wvY��QٸMK�4"YSpf,>4��|l�-W�Q���Cv}���]�m�%�XˢhM�g�{_	��gJ,���(�R���uy7CFD�!�L��Q��e��D�j�HrjK�]K�8iվu�u�un��un�n:�0L:pЂ��8��� ��btD�B`�'�6&�١4AD�:"`� �'DК�D�0D�ı,M��6hM&��4%~ܟ&�!���'HX�<l�,�X���c�c�Z�k[b"pD��DL,�bY��AA	AL��4&�K�5�A��6�}�sٴ�7����C]ᯤ��kO6�{7��3l�'uZ^eo������qe�T^�V�L</�j��x�ޭ]��m�w/w]�+N�}\���*�������Qӷ3�ng��wp��5=�o�=��&(�����0�C^�_�W�7�P.�]~��&n���D��t�Z��7�M��9����W����z���Uv�߹~���{ͪ�U�w~��޿{��������r��{���Uګ����3����m�:�-�[n��:N,�GRHk���$'�k��WMP�.�+��!�TzY��(��͉�q��U
�/D�*]����b���7^t�}ߜ�-r�Ds�ܓ	QYG/%�G,�	DE�}Τ��f�̐���%�8L�t�:,O,.}��0'aS~�84s0l�>�}�S˵�U��Tѡ6d�������1���cۮ����V��Kr/�0��~�+�Sy0gUUZHl�h70�1=7_vF t�،1(��rdМ洿^��QX�UHP���o�����}�r#���f<c����>��pЇ�a��}f��}�ӂ{s^¡�Ǎ���6a(�K�+=��E6h��&�3�p��fp9�E��k��ԉ�s���;_�m�|�ζ��[1lb�u�Q֜m���2y&Os�����r�O+$�,9j��y�,&'D�"�x�d�s;�#Zզ�b�#V(�F�Ɏ���[-N���YYr:�qB�R�^U�I�UZHoz�ʓ$p�K�p�Y�jYf�W ����	���Dz�WC��I$���H
oR:���A�BP�����s.d����2"b�asSsP��dD԰(��I�0P���VL�<h�1��r"��F��_q$p���|n��u;F}9w��4xt��|یc�-��ui��#��YqF7��UV��Gi|.\�a��ڊ�L�P�,ϡ��kK)�!�d�0��1,�;UeVW�WH��:�#f�s�w?I��m�4#�s�q�� �ȉ*�����E0a�ݗs
��cbfMJL"fT9�R�>{�p,D*0\�&����&�+nmO�u�|��:�O��<&0�Qӆ����Mnn�R����ԥ�̶��*���k뭙5�pّ_QQ��0lDȊt�B%�V�7ɑ�&�T���X����7-�R�b]�K���7�L�n|h��a������t�+��\oЯ+��sP�V��O��\=4lN��Jj��&�j<��>5�B}R�L}���a�vpOFy\�ը�ޒ*�Ϙ���ض>[��Ν!�8l���xJ�x�ŒZ�R��UZH{^E�k�Y�2��wt�[I�0���C0�Bkg�*��W5��4���%��2l�x�����Yr�Eb8�:4!�ML�3^������q�992dNri,ĩ���C>ɑ<l!ΆL�S���Afϲ��N͇�W�M���<�=����żz�]mű�c/,^^B�k�TZw;7�Y�V$��7#C���o(�񰔂�܎4��qKCq�ITS*��M�ج��XE�2�T��ԙ{��ƴU>ln�5,,�V�(��P���щ�r�|��].g/���$2�1ٻ.�.���9@�r'X��T4�!�n�Y_�'=�^"2��~rК���M�3�-<�nlD��I�g!�f'���:hM��E+'ڎ&�"I�ٓS�:l��B}MkT�J���bzll*�;�,�������^6��c���R8zt��4�Vȏi��������)��ku�V���-�[�κ���o�^��$�9�UV���Y�6�td�����R�}�\N�L���B��"���0%u����/��M,F�Qӵu�F�Hg���;���֍�#�`�u2'!ɐMK�ʦe�bk9��-�q�W�D���ߗ�ۈ�={x�!��e�X��&��2x�X�-�[�κ���o��5���k[UUi!+����ƾ��/���7[���*}˝4Q�(:vQ�#jhᒋ����-����Yk"�>�n�����˭��++�y�8���ϧ��L��b:T�LCz�M"�E&fA�N��M=�6D�+ׇ���޺�6�>|�1n�:�:Ӎ�qu#�5��s)���\ꪫI��;GMϽV�h�l3��Bn|w���1�6��W"o���ʁ����QX%�U[���+������K���,M�]���3
�;�eC���\,%'aYm��P�2X�څ�E;
��jM͈�'���E��%�~��?'���T5����c�n>c�>qkun�Ÿ�VZɇD�e�DM���:"lЂ$4"lDN���0N	blM�lК �"&�DN��4 �D؂'L:X�%��6hM	BP�!�(������D�:lD��K͞<mZ�ǌc�X�^0�#�g�N�'D�|%�f�AA�	�bX�"Z�~�C�F����z���o�]���>~��/ �>Ej���LWW��F:�}.��i��c��;No�^�%S�*�My�x5֡�mt�_���]8���:'��[?����v�Dս�A9���ȝj��Z!�D-M�c���[2��U�J����;�7-�24���|ګV��*�U`�},̈�	��u�&��r��%eM�#�ո�3�AgP���3���}���a�f�2��=�E�Y`�]�H�L�V:��Մ�z�E�J��m]�R����Yg��}_��sv6��x���|nn�J�����[� k11n�uO`�e���_��(��2�z3���n���K������|�Y�)�5l�^��Е��j�H땅��8�*� )Yc,�a ���hq��>V�S��Ȭ)c�����Zӥ�����X��B��L8}qWx��̊Gl)B"nT��P�ct���u�e#@�+	]�t���>v^)@ȁ�=mV�! <J��m6Ԏ��F�jUB��f�>v
�0f���F6�N�	�Y[��F�������7����j�ww~��{���+�U���s����{�Ҫ��߹�{�����Un������:p�ç[c�ź��Q֜m����I��A�6Kh�_fcHFcj�lj�*��B�2�A�7Ȣ``Wjr��j�G�:��J��P����Ypj4qK$	J��m��ɛS�m��!Hӭ@��I*B����v���C�xtNB�T8b}��*����#D��j*�C�c=O�
80��GNN�hJ&�ϵA�P�(b��w"!S��[)��2dLk<�ݫeq7F6�j�m`�X�E��*�WKm����8��b�؏VIU+O�V�箺�󍶷ϝ[�K:t�D��3^ʹr��Ǫ�UU(K��,�E�.ቑ��&dܲ�� קQ��$ٜ�Da�0�xܱ7�h�C��:R���;.a�N�d��S��r��@򍑨����T��T�O��2f}��0����o�x��s�\��[��r$�E̍4n`4eɧ�lc�c�c��]GZq����h�a�s�����{�Q󽢕����9��'O�4`�P��V1�?%HG�����j�c���mԅ�ʾ�q�(ӣ��s1��=(�w�̦�K��y(���=���uX�A�e�&`�&!�1q*}3��B����L�%�*\��T[o�1�>c�|Ÿ��Q֜6Y���{�^om2�7.���К<��Oqx�,L��=%�=�~���h��u����p�����i�1��T-Va�bn5��H�^�����{�<30S�o�W�9ڊz���3����F����������%�ta�Cb�ܹ�"�leE�c�>�1��Bg2�l}0^C&O�)+Z33*2f�Ui��O>q�1վb�x��N6���y5��j�/.Y8���0��nb	[���E~o5�����$a�0���nʝ��CQV��V�X��Z$�&r�pRI%dn!J���H�,���ꪫB^����xM��e��n[�9]�ZN2LMѫ&Ks/R�Y�F�UX�/�這������Ŋȋ^��j7U��r���	�v89r�d��;��<AI��8w�*���}3���&kТ�6vn�ʸWJ9]�G OpG��"H0X�c,e��Z,�Ƀ0��)E����jl��'�:��V�-ǎ����o�T��fBZ��X^fEW�UV������l�:l^�XF�WW_v�'~��9À�cP�UI!�b�K*aY�#�J.!�Ɏ8�Z�7�n(��Ą[c9Ȫ�E]@���l�Cga����r5�m�]���h�IÉq���>�6�>�1��|ۋq��[�-ǎ����e��nc�i������UV��0�vyU)��ɠ�9�s�4	�Q��j��`�-C�͂X�@������F�-�Y.ڹk/r(�jPHM{)M*��������t齂t��e����G�M<��>~���ɩ���Z�=�[���O�b�8�uo��:�:��e�u,^K�^:�DѾ*��'j�>�/�އ�IS�^�ܙ5�Q�`׬vVP�PR's�� 8�aA���H�ށO�eQ����gvWaX�w�af�"}k�|YSaFu#CG������������FΛ9�Af�+<_4�8rp,�|L+��~b�>u�V��1n<u�u5ժ =������i����`�u����X\�cY�ű�A91���.H����N����X!��;��I�;�
(�B�#.�dƠ�ծ�Tn��V�Cj�T����c�xk2Y�٨�j�f���;ꪫB\�U$���a�BI�wv�d˸A��	Q[�tn�.�5&B�OL��Z}O�aG�B�}0��"��.�[��D8d(���l�O	J���:4��,�����sG*��|�.���sef8P`���r(7 �#" �Eq���Y�o�|t0jz1�~���v��8���~u�|��Ÿ��Q֜m�r9�Κj�i��f��UV��4}�!�M�����H����'C����&O����A:d��K���& ��9�)�� jK%����+�b�T��0��"Z�11��l>��|r�7^j۹��������F��N�a��%�H:ǧgs6UM	�Q!�~�-�=�N7�O�|�X��[�un��`���D�ӆ�HlD؈���� �M�艂`�pN	bl�Bh���:"tЂ$b"pM��"Y�ı,M��L���:CBQ�!��Bp؉ât���~zǌ-h�1�ŭո��Z-�c���X���[x�,�B � �"QBi�4lM�:?]ﳒ�`����Z�7����؞�o�H9�=�%V��>�?���_�FE�/u7��_���Y~�L-4���n�`�|\y�͹nâ��w�L��.|��-
x�3��ߖ{}�^�s'�ǿ9�=j�V�������Y�����������9����v9���:�4�w^g..�s%�bh�T=�{ߚ٣�u��$�=��>Ҫ��������{�z���ww~���{����*���߽�{����J�www�{�:p�çO<x�<xN�0�Wd���UUUU��uӈ��l4`=
.�T7�"�U��J�
M���a���"�['�AF�+@�lYż���<���v���StC��h���E�h������+��:�C!��̒���*������>[�c�Å�:C��6Y����n{0�P�s���a0���pX>�2e�FT9�C���2n{��X1-�1�&1j1@��V��87#��� G:�)��0ܕd�;�6`�}>�g=�&�L/иp<d�����.?	�TC����Q�h�J�aA���&��0��Q�6}����5;=>�~������ku#��lu����1վb�x����j�}F��jYor���1�VZrخ
c̷�ī�@��X�l���:�*,ɗ�3-әA�m�.��wT����-x,� 8�$n�'U9�lY0�5���Ͷ�o�w�F��B�}my$�30Ӛ�"]��a�f5�v����&{���[23�aF�="nb{5t|>c+�i7'�+���_:;=�w��8p�����飡YE���M���}H���F����h��f�����4ȥ�]�Z���Z��|���j@v���2:�QB�Wǵ�?-g�+��io�[|���q��Zطu�u�I���N��Ʌ�w�UV�F�]�l=6kǎ�kn7���0���ߌ@aG�ÓG�:k��S�]�-��8O�C�fQ�����fZw���l�1�6��|6X���B��f���K]������fr\4g�������Us��ʫ���8�a��tç�Lç�t��$�X��,�8�C�%�mUU�4$��|_.�5 �MMLC��:\�d=�������ݎ�����Pl�'fs׉�����	|*���$S�㤭�R)In*�Zh����ɸ`�;0�u%C�P���KR�CC�K��w��X�\=���8d;u�k~|��1n�n��u�u�I�+����=���o���	�����r��A���t������gӁ�ͯ��u,�e�d�,W2��+Fk����8=�H�.��4Y�zvd�h�g��H�ɑ9*o�~�fO�'�)T�;�{���oa�b`�1P��*z�͛Ob�S�6x��6뮸������u�u�I�z���0��4��[E�A㍺�+�h� 6�m8EV��irZR8�Ƴ�K[Q�Lݼ�m���ާql�,�W����*�[0p!v��"�Q�V�`�,�'U�$��2QT84딒V�9�UV�2bl�����d#�m-��m;�izU'���!^����c��4jt��Ȍ�����a��\9Jo�mD�u��cd��X0<�3�OVh0t�x����8h�_�����P�}��Uɗ/1���9ˋ��1�/��g9&�l�ɠ�}Ki�?�IRO)�5)ݴ��~q�qk8t������8V�F;�����i�Ϊ��4hhB�GڢϹ]���#��[U�1�2����
�|[��m�J��
(�~,d���4��pࣺ
�a��ꮦ��Z�K�g(�6�,v�E��F�Q�<o�.gR�F�珮��홛��Q����a���I't���~�I:�n?8�1œL<t�C
� 1�����u��UV�UՍI'�����#��n�zD��l8#S�a_C���Qaڻ%�oR�Ѣ��g�mgь��(>P�8 ��R[��e(���djQ�!tɦ���Z�OfCYOw5E4�ٓ��p΃��E_Sg�8���u��n���ź����Qָ�J{)������]zj��jÁ`V��腟h��J��b�QpV��qE
>�[�x�ԧ=�S�Y�>�2d��>2rzr�)�(RS6}�S�Ȑ�S�{+ᣫg��ƾ�F���9�N���*p5J��}���b��*�,Hu!�6^�l�b'�~:"`�&	�0DDât��D���B�(D؉�:'DDL�lM�lM�ДADM���t�H"&�D���tD���bX�f�Д%	D�O�D �'6DM��b'��Y�޾i���1��Z�[m,��ַ�Z��ض1�q���?<(�xAA(M6&��W�W����[���I2F�)�>5j�<�5��������2o����s�eB��ve�)i	�Vc����P�T�S��{}p�Y凥�W��RL޻����O�����{=��=a�:>1��p��VX�l�>���~�>�ۦ
*�(��J�M��7�2l��=[�f\��a���
8B+deZU*���VZ�" �#�	����R<WXNYc�_����;�E�I�]��m�Ejg�]����lx�B�8="�G�Ga��QWU���&L��֋}ܫ��{|$�6C;'G����	'���c2��O!]	mFJ���݊�=FJ�@Zg�w�5���H�&=3ڢd�������qaeg��Pgu�gZu��^��M%� �W��(K�ȣ�%~�T��Q[�r��˘���+����qBEJ7D�n��b�Mڥ	mu��RXF�K��R�!��9F_�!�T�w���R�c*�vR<Rc�M�Si�yB�r4D&����Q^�1����̲Jѥ�/-��4ȷ%e���q�R�6���"bn�(�S���$�Uȸ�
J��Ec�\�$j��,%��Cn�kd�7��7*�՝�s���Un��������{�q��wwv�����{�q��wwv�����{�q��wwv��Æ:pç�b�Z�c���w)���4k&Y�HQ�����"$��W[# �������1�
'���$CpN�弪F�; �EmtC�JP�W�, �؈
��0�YQ5�#x����m��x�=i�$�dR�9Fh�*���0�H`�t��+:�]⤸jvgJ�?��(t���TqT�C'tr��C��l�}�I�ڮ���i_?Un�.�G�[״���p�e{g�}Xl3��Z�H^d�H��e�H���釺���}����g�9\m�?6��1n�n�qu�TZ�e|��G%n�d�ch���8BT=,j�0�tDwXh�ȩkX2dq2`���ңa�d�|j�3�	e�ڶ����؅��j%�s�ȰV&������Kf+�a��19G��TI����4�q24`�`b}E� �ɠ�"�B�G<�*���I�p�e0SJۯ����:����G]G�TZ����s��nY�k�,�"s*��Q�8Yc[�J�JF��K0,<1ӛ,�5
1�����N�2rgM���х�19&��*�R[Kiv��E#Q[����wip�pHnQ���]e�}+�>�zj�o�<jJZ=���@����,w�UQ�f�fF;5f�UR�邎օ�GۓO]x���\Z�Z�c��눵mq�ffXcl7�żk��@*���a�8�S��^������#ME�U�2!&�k����Wju��G)]��բ������;&MϧRx�%i��+���?F:ۧ9[��d�e�aч���@斝ҭ��w_p�*W�]c61R	����jJG�~���ʯ�6�έn>[�[�quq�orD�<jO<~�pE���O�m�\D���3,�Ǚ�%%R-���h�Wdm��ΐ���X�̘덼]�)%�M��P�O�W' �d�V�*�3/� qc!v(�b�u�K#b
9YSV���~]KU_#�
j}�2p�t��l0Lqh���4L�73�5,r&2)0�qvh>��f
sk�/����0Ѱ�N�s�?���"���5Ʀ!�:�vv��h�<~���6����u��`�����a�GQ�P�k.�^l��7�U�<W0�!�3��̖{���b�\1߁pn9>B���Xt���k�)������g��8�����ՠ�'*D^�~�K%bep��� �c*�|�ؘڤm2Ә(�<ca��Ne*"!��2�0�P�!��g���3�L�j��O�&�c��������l:t�Nl��Q��U��9$�Q���a}�۫���]�й�h���}�p��4ڱm��7��/`�̛2�l=���)Hڢ���JF�U�r/��\���xz'h�G	!��@��_��5Y6d�U��7d2l�0��9Պ���96�F��9e�f���G*����s����8.́���G��b�Z�Z�m�]G\x�i+�u�\��X�݉{���U�<BҮ���d��91Q±�F!�j\���D�Q-˳f3�.�i麐��d�I��Z�s,98l2`4e��)�8z����'ڕ����:vz�>�Pfap���cf�����N�lq��8��L8~!�M'CE}[�n��x�f+�2vي�p��]��zm1�h֭q�ls����f�Ssr
Z���(����O���X�p��W�
dO�hQR�(�!� 8�.��k/�uʤ%�!���/&qj��q}�O��5v]�;�<�й�X��(<�X��MI�P>����R����$�h���P��ң=��n\�ɀ��٪�	�l��*裈R�q(�I�d�
3��|
._Й��h�y�?9OΞ�8���1�-խ��0�4p�HP��=tl�ʚ�/'|��g��k�ރ�C��NO�ò���Sw����00L�'j���S �����|�LO�\O��_LD����y�A��c�-����G��x��/�>,,���'�A�X6��jf'���SM=s����wo�i��|�X�&	�`�&	�"&��"%�6""'�B�DН8hN����lM��6h�A�܈��'
D�"lDN�"",K�؛4&��(J:S$ �!A4"a�(�kmŽG��0��1��`��p�D�,D艂&�cli�i�a��Z�bhMdM��8'϶��ޥ��V5�;����H!ւ����U�_?��^�n^�ϯmcȤ�n���^�snnX��o�9������~U���o�zI��\��[�����s]��3��/{wx�5w��07*��_>�ϫ���{�V&=���i�;c�����t'}ߺ���);�l����}ȏ{�ۚ����>���ο?.�J��GE�h��7�ټ�Y9���U��89�_k;�VjM��'���t�8��;�]�^Y���ob��s��ߤ�n�O�q~��Oޛ=V��l�_����w�>s�Un�������{��wwv��{��{��wwv����{���U[������N�0�㧄���4zgJ�͗��^��/g��.d=;�p�3^!g�~>�Q�͇�D>��qY=�6���\X-��XIV#�d$J�(̦϶p.�;9�k'�2x���}�d�1������e:�u��Ii��f�b���5l�C=��p���n��-խ��u�uǍ�������Cw�uUa��LL�bfL`�r�:7E�d�wp�ő%F�/F�s7��5C�~]�C����P���KNCӓ��sa/�K���=ق��mF�Ns>*Y��RòT;��5]9����v��<�j�4�6�q�uku�uq�S��,���ٸK��Xg1�4w�b�CW,#E]�ʨ�[��Lq�m�X� ֧]š�Wy��Z�X��s6)V���:m*�M�&cLX¹��֜��Q�N8�nF�e�Z(�]L|/���7�J�,��(��%U:�RU�WG�O�C��n|`��|��̈́ѕ5rX�8��6N�Aٱ��C�#������l��A�p��L�6�a��v�`x�0��=j���~�ˢu4�I��
8�Ey 
����!�(*)�B|Y��|�帵���������T�Ş����I�oV�31�:l.��4pU`ˠ�A����)Z������Ю�����IgǬ��8�FG���z$�߀;D�)S�];_Q��	�W�{tk7v�-�X�`�Q��m�.�5v��0�����/1��N�v>Ӿ��
&�#����b��ۋq�uku�\f�2pDIuQ�yF���e�R7L��t�\�#�s|p;gɂ���eJ��GM�G�T[�%��lԨ3�h�A�,��F�<`���V/a�?{�����zv̛EN+mD�W��>�wǯ�q��un�L<t�N,�ֵuEUϷ��0њ�P�UI����t�<>3�WTY:j`��h�'�џ�[Y�ƫ8�f`�W����36ۂ9��Y���cUf�MI�Ҧ!����\�j�;.;ɓ0���U����3%��T>��d�U�2�p|�-�jf�O�����<|h��g�N<:|8C��4xp��#��e����ֱ-�6�B�2��U�W��q���h@֛�!�,iꪸ�!�F�|��Ul����+�-��8��69h���h���*���weY�tV�V��0�LΠ��\��(�
���gd�*��}G�J>�O~QT�MW�X�T�/�}�D�5	�M8d���fc��Uʈ����y�O<%U�S#W��'�w�T�� ��:{O���sܓQ֚b��q��[�|u�q�����U")$/^~�KQ�ڪ�f<zx֍�_+[=�p�9��'����[V�LN3ᩱ�!��h���Y�ګvYd+tgw9�7��<�Rp�F4`�3�h.��㒥�K.�2@K�H�I�K
��+;9����ٍ�W>5�&L
�r}(�3�z��m
ο}���ӕ���?:ۋq��[�|:p��l�'}���7���!���Uc&!�cتDh�>==2f	�>tW�E'a����R��Frzf�>�l��v���i5%�zm$.]���ڐ��"� �9�����Y�Ӵ��q�J_��];����T/L��5=�jҌ�3�aF!]6��d��]vN	[��4af=cb�[�a���6��u25P\�c��AWH���� Nj�K~UT^-�a�t��L�bT7(��M�[J���I-#�Ѵ㭵-Rb���h�.�}F�������g=p�)�pK������SBϴʒ��NUJ�2��g������8wfU/�8p����k�;��R��VL��q6�)9ٚN�_i�GzB$"I�$d$�D�
*��G��~c��M�����,#�WňnQF�PpDB�b�@དྷ�7�f��"�)!��LDD`�`���F �1E(eb"1�0A���A �b0I��bb"A�	`����� �D`�F1#�`�D`�`�b"0A�2a � �$`�F" ��#�#" �`�#"A���Db"1H1��F��$$`�#Db ��b"1"#�F"#��1$D���""1"�B�.�0DF"#��	 �"#"#��0DF"!�#A"�$���""2$�"#""2$#" ��"	�(�Ȉ����� �0D�"2#`�����Ȉ��"20��dD��1F#"1 �2"#A"�FD�Ȉ���0D� ���#A"������A�DH0D""0A�""2$�0DF�� ��`��#`�`�����Ȉ�DH0DF��`�"0DB�J��DF"#""0H"�"0F1ČDF �� ��A��DA�"A���� �bAb"1" �D����F��F$��b"1 �D`�b ��F �1��DB�L\(D""DDb"1 ��Db"1"Ă�D`��DF#D����ȃDF��A��DH0DD��1��DH1��DF"#`�`���0A�1��bB1$`�@�$�#����0H"0A� ��H"0DF �DH�Db"1��DbA��"1!�F"#�DH0F���DH�Db"0�"0DF"$"�((1��Hj�A(�EA?���*�J)jU	J�UH T<B����*R���AT�A	 ����(�) �ʠЅR	T �T��	 C5G�P�E@BИ��d��H� �U�U �J�*�����AH"�T�QPJ�A
� A)Hj��A*ER��)PJR��+JT��JJ�AA*�"�QU �T����D��U5I�jR�T�R�% �A*�R
�A)A*�*�T)A*	H%AJ�"	URR!*	HEBR֊J�B 1A� n�
�F! �)B�T"	HB��%B���BUBA�dA�A"D �"�"��"
�B��%!T�A��" Ȃ �2%D%!��!*��%!)
�D%!J�BUB!�P���!	HB� �AFD �2 � �A�	�ahd@�!JB!)BR��D" Ȃ ȃA�%!P���!)BR"�"!DdAdAdA�DaA2 �AD��"�" Ȃ0A"�dA�$A�� ��JB�B!*��"���BR�	D!	HD �BR��R�� A�����"A �1A� �dAH�2"!*�D*R��J�BT"��HD%B���D �F �Ȃ ���"��BR	P�%!�BR)�%B�"�H"����� � �12�JBJ�D%!JB��G��JB!* �� �B!*	P!	H%!%B!*%!���"�Q	PD%B ���D@b�A�AB1�bB10@`��	HRR	H%!R�JHRJ��A`���D"�JB� JA*)�����A
��D% �J�R	HB��B���% ��R	H�(�D#�� � 1��@b@bcE<�% �
��*	H$B0@A���#D��JA*)�D% J�JA*	HP�H%A)#D!�d% ��*T	HyT"�@`� 0A�1����DF 1 b�T�% �!�% �0A �0B1H0H�b�b`�D�`�`�b�A�"1F$b"0A� !��0A���E!�~�BQ��N�6/#Be�7��HOCJ�*
�F(���o ���ZN�ƾ�~�mo���D��&�]���t�{w����_7�6!�u��n0,���6�(�?����Ntu��u��'Xں����	�I�?���N�(3�ӿ���N�EP�'g˨��?��O��� A?@��>�"*��T��D��$|�/���t<D?��>�"P�'�7��<ǭ�X�:YZ���@v�o}�<�B��i[�4"x��(?W�4�q��O*On'��Ĥ��&��^�5��w6C&�D��daLWgǾ˄�0������9=e%ܔPE(D
lD@l��P�KDE�U+h(� 
0���
�Fp-%A*�M���on�Xx_���Ǒ� �T@U@�TL�A� F ���E�� (+ B�K�Co@�w �L�?I��� G��h����`7G(g��?�92|��C���E�_'�A���4�#@���G�d�D�����˫�9@�)�py�[�R?W{�2�<��	q���:��~`�
�C���Ǟ|�}

�=�����!�%|<1���q��	Jvn)��PU���~�H�p �&	�KYO)`����7W}�� 	�\�/e "	��qD��f{n�ĳ�D� Z6��h��p�� Xc����dh%%O�)
<CJ:P�Hae�` �6���|�#�M�I�l'�; ���s�{M�	�܏�z��p[�a� �jv� :�P�C�����w�}��Y �8jv���#�O�� y�O��@Z���� �ϴ~��G����aI�"{��}���GҀ ���A���;x~���n�:'XvC��`��&ϵНX �H2�B��� `B�:���(��-�B�������HX7.f�Ǩ�g�.60�����PU�I��^�z�^QLeD�����P �rC���;���M���v��
5��a��8?��M��'l� �pv�=��@�M�����ht�@�� ��a�5V��e���ry󙢁�<C[�0�����F���$�uk����.�p� �k�