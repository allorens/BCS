BZh91AY&SY*KW�,߀`q����� ����bI?h                Ȩ���D��JEE$H��DHB�����eU)J��Z�D!UB!�Skj�D�`��6���RPJ)���]��%4cf��*�D��ݩEITm�T6�IUU�E��T�PTTJIP�U@�$��X>�����������R�7�c�%N��8e*Uu�][h�Ҫ)N��8h��-�-��*J$eI$UveR��j�DP�liI�R�eRl��uB
���y�   ޛϽ/f���e��un��v������:���ԭ]5�s���e���;YV�Y]wF�٫u\仕�U�gk��rWgVm���Wg0uBUR�)&��J��@� ����^٦�S�ڥ(�ǧu��Wzz��K,��͐���g��U���w5
Uv�x9���%Ѫ���/j�[mh]���QJEޫ{�R�EU�[^����U*S�J�@hV�Z�@V�J�)�ҕJP�x�.ڪ�¾�y�A��=���>ڪR�m˞{�{�S�*���o�����m*�M����J��Ӷҷ�|����v��[K�4�%U)��u*T�e�O;�B�T.HR
���$ ��J���o�J+�k�s�y٪T����}��K�ѥ
�O����G�>����R�'�����\�n�}�W��I�_w�{�o�J��l��y�������t��P��uR�EB�D�*�t/��4
 �no�UA:ͼm��S���+7�����:��ܼ��UUU�}�Y��}�PR��|/��D
����v��m���y]j
�O{�UU�%מֈ(�Mmj	UR�n�(� ;۾�J���S�v2��������UWYox �� :��w� �N׼ ^w���� n�p�j��R(I(��B��$�!�^})AJ �^>Zh����ո hs��PΫ��=	�� L�{�����qAT�3�� ����rP�hR-�2*�R�Sϥ������*�z\p ����Ɣ�ޛ��v{<��GA�w5��W�i7��A�h\Y��4�ٸ� ;�$TGJVE)D��=	�P
�t�� [�ޠ(�z]�� ;�v���\{�@��N�QZ'���n�(:�vlp ֻ�� �,�V����P���@���{�w  ���D��0zt��Sͽ�� <zN� �pX e�� X� ��}        ��JT�� h    S���MQ� &   i��� ��P d     4���Hc(4� �4d�&�!�����0�ц�1h �Hz��*�'��5O5F��dd��3S��ߟ��Oӟ�~w�JS�O�4:�?z�W5����#KQ��ҳh����;���\<�����DPU�
�"��p� ��@������qS�TX?�ʪ�ϡDAW���?� �������?�9��q�������v1�xq�gƛ�q��1�g�1�g�1�c�zc�q�c0c1�c�q�c�1�㍌t�3���1�`�1�c�0c���3�c�3��q��1�8�3����1���q�鱃1���q�c��g��8�3�c�1�q��l`�|c��1���8�Lc�1��64�1�c�1�c�7Lc�1��1�c�3��1��1�c8�1���0t�1�c1��c<g�1�`�|lg���c�0c�	�c1�g�q�ǆ0c�3��3��c1�v�3��1��`�1���3�cLclc�c�q�n1�c8�3�8�3��Lg�|g�q���1��q�gǷ�3���1��8�3���3�c8�3���1��8�3�c8�1�v��3��3�ݶ1��8�1�c8�1�3�c8�1�c�1��c�3�8�64�1��	�`��1�g�1�8��q�g�1�g�1���1��8�1��q��ǌc8�1�c8���3���3�c8�7�1�g�q�g�;q���1���8�3�cq�c8ό�c�1��c�3�c�3��8�<q��g�1�c��1�`�q�xq��1�c1�1�Ɍ�1�x�3��ǆ3�c>1�����8�0t�1��8�><1�3��8�0c��&2c0c'����8�8�8��2�������2�0�Lc"ʆ0/L2�2�2�l����)�����0�0/GSCS&�T����A�Q��D�Q��GG����P1�q�1�� �SGS�T���!�����)���"�� �(� ��cL��������#��������U���Q�D�q�1�1�q�q�q�q�q�q��D���T�q�q�1�1����A�q�q�q�q�1�<g������������$����8����ʘ��ʘ�����cc"c �*c
cc"c#�La`\deS�
q�1�q�q�1�1�1�1�q�����������
c� �ccx��d\dLed`\daaaLe��A�P��1�q�1�q�q�q�a&�������T���;e\ed�SN�eLe�SWGSS&���T����1�8�c*c*c �x�8�8�8ʘ�8�0� eSGGq��SSGGGGS:`eLeL`�SS �W��E8Ș�8�8�8�8�0c�q�1�1�1�q�q�q�fq�q�q�q�q�q�1�1�8�20�22�#�����L�����c ��8�8¡�'L	�+�
c*���
c(� 2�L.0���c*�#�,�2�cʸ�x�a`eedq�&@1�q�q�q�1�q�1�ed\a�1�q�1��WY�1�q�q�`��2�0�0�0����3��7�c<g1�1��8�7�̘ɌɌ8���8�3�c8�1��7Lc3���3�ct�1��l�8��t�3�����8�7l���8���7m��=3�c8��c���1�����cq�0c����c&2t��8��3��>1�c8�M���l�3�c8ǎ<x�3��3����M���1��3��1�c8��8�1��3��0c�3��8�3�8Ɍ�8ό�8��t��0c=�c&1�c8���3�0c�3��1��8�3�v����0c63�c�1��q���`�d�q�g�c0c02c&<x�0c8ǌc3�c8ύ��g�1�c1�g1��&0t���3�����zg�1�`�{g�1��q�fq����c8�2c0cx�1�`�dǷ�3��0c7�1��<g�8��0c0x���q�g�q��g�1�`�g�:c�`��&0t�Ɍc0x���q��q��d�q���`��1�q�1��`�N��g:q��0vɌLc&2�.0c1�0c3��1ǿ�Iɾ�Ǿw���~��G�}�1��`�*D�ح
+ni�jK^(��A���K�ҋ��Y �v�7����f��17��:�����L4a�fTf#z�ȋ�������:�In�͈ne�t(dBN�Cg�Lɺ�*�QZ��&�N�L�+t���W	��-#[Xl��X �kv��mZ�xc�m*�l�ۢ5�݁\[�s!w���U-2�R��B.�G�Ȕŷ�4qݛ�6`H�J5�����6p�X�HR�I�9W[)���)�"��v>���geJ�\W�ͩ�B�;�SJ�cUE��(fQڔ��Nۣt��˹y%��Z�su$n*�J��U�([�n�Z�SSn`�m&'�1u]�Q*����֠&�mނ�$d�NhYfm�
1�܀GF�]�sF%x�QO �MJ���T�f��R�ж��%��2�����Po����X]m�աG�e4��J�6bs�Wy-�,yZ��H��j�y`M�!��TGX�[E���&��˙��#;�B�UhC�l�6��j�]L�m��J��&,�Ɋν�
,��x�n"��ʨNf�f����Z�ٲ��3$*n��"�6�bb�
�Ű��ʷy���.����^��xwF�;��EWOFk@\����G=�[JQ�G ��b�h��ϷJ�x��3����Y�"�R����LѵZT(RݳoP�q�R��ي��faSR�a�z �Sm�N��"^UKeEAf���3�m��}�[�ss����k]�[�x��P��"yE	��;4)L�&��3�@�I�ɿ�*�a[���6�n�3!CL��*�l�Ч&@�����L��6C)my�CV^�lg���i�TN��f)�ZeY��Lam�3^j�\ "Y���h̊�1����ȷN���1��^$ZT;+h��ZSyڛ�N��\gɋ�=��ܘ�&.͹p]�	��V���de���ʶ��m�KF�vY�T�����֗5�^��v�"����ԩK%�����J��MR��i����gL��pP��wa�r�v��b�cb�b�rPT֪m�L�.�	g2emQ�i��Y�+svm�=�������jV�P�mf�kaݲ�T	^JM���ܲ���+kNy*2��w��4"1��ֲ���N��h@B7tZ2�d�-;P�F��zr36�v���C2S*��ōಮh//<�۹�6¸��/r��8pM�U�����;5+neGk`L�V�U�]\�[)i׹�A�I+e��!
�Ma.J�`kjh��L�7Z�,���K��L��#��N�-� ����6��m=�V��v�b��̕O-�*�J�C�m�`Zn�JB:sh��f��.:��M��D]�LŻ��oj��#ȯƫHo\z"�ynkA)��V�TDuy{���f ��Hk+�ԡ;gv���\�{V(䭓3��ac�R¶�Jc.�f8��J0�3�fK�
�u���d;[E)b�@�e"P��5�M�0���X-��SթlY.ԙv��Y{`o-�
Ym�Ռ�V�+o
ʗ[gpc�l�lu�rTlc�b�xh0��9m�3Y���t*<R�e���g0�,�C5�Pc�3pv��-�ŉ�`#p�]��~H&�m�0�b�b�[���	���u)J�3�ّma�o��5�;glZ0-��#F٤�	�Dw�ck+�E��Ȧ�,W�Z@���4��EѡKd������-)�Lܙ
Ʈd~kٔZ�-bӴ^�f�xR��A�V���X�:��U���!j��d�lHYi�j������u�x�:b�H��d�Ϛ��!|��R�N�-\1�5{r�Z
�=�Kӈjl��RZb�)*���䛶ǘӢ�4�Ui�n�\��u)c�L�*�����0�ip�ʌ
h�RLwW�P��6C��X���4n�Ց���&�X_����[��BM�:.�rf�3w.�݃��Mm�eOR�&��]��ct�����j��#r�p]�@D���!ap�@	�Ӝn��-D�9��� <��'@ު�(�e-�V*�����\t#Ν�%�ݳ=r��1�bOr�]�f��E�	��So7c�*
�ډ��d��<�R���MJ�H��]&0X��$,e�lm����m�t�`�n�Ef�2�`���-x����; 1ZZ�ZMi�ye���N݉�.
��;��A�Dљl�-���r� �7�>��t
eE,IJ��o�S#�w��3z�n1�b�2aܱ��>y�-�.`�Z���)�D	X�Do,�q�e�Z�R�LiaF�vTt�ٷ�ʔ��TV��◵tMEF��p7��V��^d%mܣUr�B��M۠ݶV
K�W����BJP[���HVj;h]�}Ya溼OV��S��,A?7�����4lKU{�^�y���^Jk*ݶ�#F'�{7K�l�Ql���!9� �g�`ѯ-�R�R���{g �1olދ���s��raM*zp��1�/3%Vf^4'�jy*�7��n�*�@��An�1˧d�;sfo+$	r�Ǒu2���ذ-�B*dV<�YXPMk�Q;7�2�h��X�M��!2�*�ֶ�&�f����0b�3T/<�R���Sv��X�E	�(Vv�e
I*���R2�.��+Ɏ��[���=/�Q�Vk,�d��a��V#�Kѵ�A��V��X��16o���wvY~zi!0b�Yn�1�w�[u�Á哴�%U&ְZ�1b:�#���7w�n���vU�wwFS&&7[�uL;'I0V�t�شQ�����Q�Ɇ�PQR��9���dA�K2��c���׷a�L	V�n����9>�2��V�2����R�p͛��c���iZͳOIA�Y�� ċ� ��,�!b��'s)�W�N�M�䦝hnUhmH�2�Tlр���x��bmk,nY��4�ܛF���0ֈ�l5l3���ԫʹV�^��"�����{$ͨ�83n����ܕy$z��䕗�z<�6=�=,��(b��cFz�h�\�f�*��S�t��u�n1�]=��,���]��gD�f�*^I�4VLŊ�)e2�^F����[��"5�����e�Ez�����"L�������r��+/#W+M��nd#��p���ۣ,Xܺw�WbS�MBm��5�&�VG7skda���R(�®��.�=�Y���d߶��jMAYߠܨ�oZ��*�KHc:ֽ�r�؄�J��8X5D�L!��W!���N�0�#��Լo�LL���B�[�7�E��ڻ�r�ǰ�E��E1��Uc�2���B�
]�Z�Y���)���]hH^�P��#ʙF�F� D3e��*�R���Tr(Q������ʔb���(��êfy�b ��ֈ��U�Ł�r���s�Q̷���h:D+��O-�齨���M�Q�c�#ۆ*�I	�����'[����o4�[���ņ�lS	h�%9Na"����k]��Жt;�|#� �O*��X[���^�d�j�e�ڕq�*�Q��)�L����$FAr�g��h����.d����ъYYP��;ۣy�=�ټ�a��xcfF�'���:���=fe�3��52�6)E��p\J�hf�s.�VS�j
N1p
ck$UA� �ᒚݕ{���c�����U��P+QT��vY%���U��6fl9JE[M�EcA��6�;;T^м�:k�P�x��KF�R�y�P���٘�8%��֦S*�-�sٵ�ʕHՂ�؍$�{�ڛ[��,
㵮��1���	�KT�(�t��lA�7[v����i�.����h������*v��]��XopZ�$ڹ�'C	��,��Z]2ѽF���Bj�+��D1ݐ���6��$�۬Z��W��i���*��F���+)�s<�
�Ө�tܪ�\U�̢sm
ʐ�vn�C�zj	U�U���	C��ޣF�V-��
�^l+�nfmm�(9MQ $bē�9J�l-GM�2p:�Z &@i�t���k�f����E���D����2�ш��mޔi�hR����R��5A�7`Xr�Uz��m�b������ ԯ2���r=KS�Guҩ��P��h��N�6�Z"Ӥn���{LEtpl�)阥�v�c)�kM�L�������j/ڍ�V��t�	Fmǻ��%��4YԶ�RL���M 6�%䘎-e)����wv�v�@�تe�MXriCջqU�b�	��\�ف�j� ������-k�Pgv�%��@���A֗Bl�ث�Ԟ�LH�4^�Yg^M�݌��\�PYp᭧/nkw��.�f+5�!M�"��;���*l��mt�=ЀY��+6ˬ	b�$��ʷ�,�Kn4MÀV�Rl�y�bڹ-Ve��Ĩpn(�;$�-�x�*Ь���I0�i�D�cٔ+I47wve�&��[��w㰷F�a�n^,�^�i��J#"��b�f�.���n��6�mhdX�A�m�5ڽq84<4Fh��.��D���t�;���ue��|����ՎM�l�V��q�F�Ҵ�D�h�����L�*�ڊ���ܠ�f���A#����j6	˵z���/bn��=�P�%n:Ĥ
)���ݳuYh8؊����2��z(j�h�N���B����c��*�j����^��X�㭖��7��6���r�Ï&���ƆLr��e�jQwg)ݙZq�2�7b��1
�����+2�V�sT˨�X��*�a��b�Pb�L@�#BT�B hc,VGiZ�Vƨ�G	N�����$	ODq���������9��rũb9&5v�H弩���
zA�Wu��-j[�m���NC�&Ңh�C�汤j���F����4����!*��%���vRv���{�f�f���xm�;cH%ޑ�-㪙19u�H�Ϥ�u&�f�K%�!�,��W��U�0�`�����-��a�cR!E�`n�v]4�����+6
�����t-�z�`�WO�ɷM���M͙�		hf���Q���^��^Ú*]^l��nDF�6­b�4r��PŮ�Smf��u���2͋]5�����:U����b9u�1m�UlG���BIu{	fc�ō�m+W2�F���#=8e���J=z2�=�z��th#y��2�܂.��Z��&��d��ԡ��Z��;�j�+b�����Х�}�~��=ю-���=�7�t�h���ܶ�׎�VD���
��=�z2� ��ͦ��g=Û���p�������V[f����;d���C�5J���^���]"j�ӊ��Z���w��ro��|�b���|�>�K���Vr����ٜiH��@z+���te�m�������
ο^�����"ŤPM������+,ާ�U5���z�*h�1Dx֋���B��o�rj��2�_G�9��-y�Bn�59]�%�z:��h��Շ/�wO�����(��z�q\���j�ӡHn�s-�g0�����b��6�ȅ��@��g�|<WH
��G����/�,|!��[x��b����ՙ���)Y?.r�$��bRd2�����L�n��if�٤��TŲ�RX��D}0�ʼSd��S�+,��n��.Q���%s�P�wsI���"��a�J�vgū�Ә�]�25�D�/4�,�ۖuF��J7M.���^q�+`/�
�C{�t��x�&�/l���ģd�3��4�6^Bx�ή��J��hq��vU�����KW7��H�yս-�4&��]k���+����L��XTL"K�6��wqU�ʾ	{�q�3V��6���|�v��Æ�8�(]Ǥ�+]Q��u�^�Ln�*��s/�ZT��20^�n.���*yr`U��Ǹk�i���n֩Ԉ*+�g�Sv��Б�����Γ��0��Ⱦ�8��<l�>be�=�v��W��ƫ�^Ò�j��G�.�<�Z�m����15�頎wN����N[�+7'N��za�Ýj�(�����X�9���t��_x�\�5Qg�=�^���|xW�n�K�жXn<KϽr�Bv����'ńt-�,�,a�٥J�i�:�Ʈ�ݖ���9η�����ؗ�u���Uj�X�ؗuʤ=�^(���<�IVZ�j{ѽ,�v,1WZ�Rh�³x*��Ԍ�p�#��H�ui�0�;��.��ڼy�J"���]}\^WL��ݼ�I�t�f��3`�VS
S]aU�7h�eu��h�V�9��!"�;�*ç--\�n�μ}����&R��r��-+8�#}k�F5��W��kIq��ȏ^���h�Uaq{�ޣ0�W��fD�`�<�ݼ���.e)�$v�2IFc�lw��K6[0�%.��Iܻ��!�;�h6�:Hi�>�g�V��8p��ϱ�Aa�beFj�ஆu����8ɿ�fh�A����)�!8��dX�&�]��V�f���w�b%q�����5pg+���tŦ�]�F�/zU�o۹O�l���ݻ�X�^K"��zz։�x���2΄F��@K�w��n�&�b�r�Z-h,�԰�f�y9ϴ�A�df�e�c��:��>�J�䎈�����!��v-�v|����"p�l|�z>��#�Z�ZU��s�ҷ�}j�{έU���ś8��E��f�e"�e��UN��Ȳ4�^��F�*T����y;���6������Ӥ�9����Վ�ŗ7��"���`��3���h}�Ĺ�aI��g_|��0�m�	�vDFV��uQ�}-6���2f����-�P����%�pʊ��$�M��3�.p�y���,�g�sI㷃0�ۨ=$ގ� �m����]v�h���ό�Rz/�vZH��E�,`����~Y�_�'9ۛ�� ����q;�k��Xa=g�����VNdF��O�����>#	���`e���8I�H���y;���i>Z�59h9�	xsCo��W���o1+��F���Yîb%����c[w�tG��k�gna� ��������B�w���Կۡ*���r��n�R��-6��GEcSG{ܸ��vV�x���n��g���]y���U���!��F�ʃ�z)}7F��=�vR�!�s�c�	x�MΕ�:ui�b��ھ��b����}�v4�B;w��{NZפͩPo.�bӻ�so�T�"l\��Cܕ�mb�$���\��R�����ugy�'�����0J�M��U4;��B����:�.ݞ�#K�{ַ�ظf�����]<fL�-ABN�9�.dޖ+jZ0M�1p�\�`n�B�h��nv�����z�ԑ����-�<�-�i�n��ؗ��Mԕ��˭�\�#;ٽ�4��aE�u}K�l��:s�<����5�æ���8M��p՝m77���
��W�do�zj�ݧ`�K'�:�[����[�inz��:UU���j���C�+7��8%�ހ�C���ƙ;T���'1��l�6��s4ڃ����Ht��gJ/�Ֆ �X�+Er2�M�27�"�XG�,��crֽ�ȝ�_z����X�˙�w�u�;d�TjV]���M��uvP��M�*���np�UƱ]�R�Z�՚	�\�Lpk�>}q���L�8'S+�R��,�h"�Cͫ��;����m���6b�9���J����f��D���qv.��km�Bu��Kzʴ{��᯲͝�����:{���sw1�f�*P0a�l�_i�&��:�r���Dw�g����̜�T���D���PCu���9l(�˻���,+�8��6��(�56�`u�Z5L��EH	�Nc8N{D0k�.=�m���1�6Jo���z�4Uom�wŢ��e]�AT�,����(D�Ǫda�r�d��y����=���T��Z���x�7�xK����}�k����u���5A���'^�˸,ֹh�vk��]���S'ܱf�����F>�|����A��;]}6\����B��}1^�a[�"�X���:c���s�q�E�;�u>��E;��pq�U������#()G�gTVgbf��+�*�q�Nwm��2+x�5y�q��*9*��{����T��+u��R_]��TzfW>ou�i¸Z��Ć.�2�ә��nm�a�E�!��_�%Ӑ�_c�Ue��E�6v��k�07��C8K��ב',�O�܃��"��{uΊ�й����"2���аk����r_T�qO��ףqV��74�l[8��;}�e�=%Y����voiN��Vza`�3v%C��xCe�):b1�Lqb�\���Ꮾlܲ�u4�礲.�2TIS����5.��pB��=��G�4��f��CW����l�;�޸�0vE��N�e�(kL�빮�"2�����Ū(Ef`�;"�)�K5gk҃���_.2M�n�{v���s���
t�ZS���SP�ם6��\y�z]D��̦^�]�/w�7��OE�۶5[�C]J�q)�s"y��vf[�U*��42q���o;yN�Z*��2�3���Vb�u����܌��oK��O7jL3̊���W�ft#��;-K�x�Q�%�|!}�˹��C��4o�9�,�<��Qܬ�.x�$�Z*��oQe^��u;�xz�9)@�ü	�7�LŪ��c�Y�ԝh�{]��V���������Wa�4��W��FZ6ص\8��o{P���G�w3Nr��c���kD��֭a�.)l�mӠ�UZ�ɠv�;��hr�[��������x��xܮW���u&�4�Y�_V�č��/ywH^�s8t|�����]��)�qO�l�
m��vQ��ע�yh�3�T,���Kf�uƦu��;�7{�Ɲ���rݳ�Mb�0�R����D3��4��{�-}�}t�̢8������:�WW��]i_���u��\|�H�<�"�7|�_-�ꆯ/s�S�]�K��ɼrx0�k��6���o�J�^|&R�(M��꺒�aq����E.�'i`}vd���o6��Ъ�/S�ݨv��y���pޝ6��O);��u����]\�j�PC΂�zz	�kwk;�ƣ��H��U����"��xJ���t�v�WAh�84�;���w��E��ݦ��oof2��>�uUl��-n�z�<ܫl���X˰B�[ln��&�Mw]���ېZ���84dR>���h�)JN��h�8�}�����2h�s�=�B��ף1�D��f�vU�
�Wβ���/3���cjh�ȧ��:�S��^`�M�L��\���]"�МMڻ������Z\�Z��M매NM���Gk��*�F��t�6z���]'_,�[�,���}O{�*�������ͫ��1�-M���EqQ���*��S��j�����q����	��v:�p�n��{��� �Ճ���
�f�D��zZz�zG��i����g��J�2.�:��/Xu]xkVҙ�p]��챪0�dެ���1LBp�n1�'�vt�,×��Y�D�c�:�^�EV���*p]_z��)sܶ��1��\hM��.�v��F="�-����gf�r�eKb�܎ڂ]��iSu�xW�EF��P��#�u\��	�7p+:x�;�u�5R��ζ���峉M���V�Yz�����6JkB��X�S7���,^V�ͽ1�[*�ld��r�.�����g>�oh�J��9�b�8w\��s���փA���]cPJ�,�Nb�=]'+�Vm3]�V%u�U&���˗��1q�&����\;�;��2���DVٕd(򺬃��Z�Ȅ#�E�l�g�F��V�5�.J�]B�;4��v\1���*=8F�ǒ��X�qg\��Xdψ,
']g����u���zZy����F#��3n�oV����D��@c�F�R��f�В���l�����1��5h�6}aS�Nv�ڱ3��lu;�e>U���4MA��<ʅ�};���;�;�oW����{��]�R9�2�g{>�#�7o:��7�v9�#�ՎOng��eE����y��:�>�+�U�YPӻ�)��Y���}���8���;+���f���6M��'q��]�$�].��M�[����ש*7�j&�6�v���f!\���Ͷ�P/{�0��1�y���宏Ch��oJ���s���3�P���3���{�Fot��l�m�
��]V�J1decu�Ml��]��R.͸�AvG|ʺ�p3�!��˵�ɟd�I�a�����[�׵]xl��f��kXԜj�v�������Ks%Y䭜f���zI\|�->=���� u�Ǣ�v
�cz�Y�lĭ��q˨eeӖ�9fo;���x&��4d{���gu��`W7���Y�5n�|�=`1v,��v]�Z�KUܨ^��ؔ[��d��J���$�',�$fdO,��w�����3��#�V�k�n���ֹ+�m\�)�]�fե��x���yI']�zv��Gaܡ�'�3s�yuZ6��n�p�Y��ZU9n�kw�*پ��7fp#C�Ǔ��̭���n.��-yy��L.Kܽ#�0���M��;�O���t�v�����2�յ[��+z���}C���&B`��.�0Eu�r�\�9έV^�7M�b|d�z�.���Tz�Ӟ�^�Օњ��f�$��.�U�h�����7:��x0���\�,��,v�ȭ��T�-�́B�0�q��pÕ��Z�s��8蝊�����6�0(��h�;�=���ޝj�MqgR�t`��O�J�]���\�2s�"�μ��{i:3A��&��u*M�Lu��ЌnQ=W/tF��Ӹz�@�oJ
�:��x�V �����9�k�B�r��ތl�7KZl���e-��I;9d-�;��Ų�x,/��j��5�O9h�|K
J��ڸr��J�#��s�ufh�n+R�5�=c3�|���!^�N�Bǰ\z�����b1N�G���)u��ì�2�̐���_]v݇�Kצewc.��@��a���aG���,�c�H�n���u�έ!6�9�Y�n:��)mx�s���o�������*�&��(8g^h=�kγb���xԼJ���pиi4���mȎei�
��q[^�u���v���I޼�jw*����טy娪vF2<�Z���w
a�o��U��o�LGA�p�����wv�c)��Xޣ�t(�r;㛲fEc����j��R�*���J�|<�
,�wD����s���N�>���iI�>i���il���x5�|෦���b^����B�q����6��Y[\�r�ߏ�Yʚ�i1YC��\j.��*��m�˵J+<��5l�wxm`�Wׄ����<��C�W�!w�/�dr��b��Y�)+k�[O)�Q�b\Z�u��7����k\�{j�VfM���m��sȢ���30IV'8��L*ue�$$6xM�IV{����X��9��7���*�lR��q�U|j�sU
��
�L��*�l/E�*�aڳI'+�D>fQCt��/���i3ic}M� 
�|�@^gp�T���8�;7����_)�AtΜ����oi�}2�TJ5k����W�&��L%�+�W�nػt�Ӧo4	�����^�q>�÷T�MrQ[���UO-��5ӆs8��ҋc��v�S�יy&CS1�[�LItF�1��i�1vՙ
[A����+.����u1�r�k�O*�n?�e�qF=k� ��ǃ��L��b7��T�
�i
�;
D^���Y4l]�W��nb��'��^��:�Y5�����묖�x����y���ܗ��f*ƸJO$���0����p��2��[7Eu7B�a��z����+��Xh�g��ɕ��+�Y���`}�֊*���,�Luŕ�+�����փc������9C4=GG�.!�הf�<݉G[�g�r��v�x��(uAww-����ە���ѝ��R��{�Gm�m�q��B���L�3Y\�@���B7�.��^��J��w��4�'<[u8��El���6��3
�#j_0�ڵ��3��L�@{�����Q��}@��宑u��hP��Y4�V��:� � �j(���M�*M;��K[ڵ�ڭ�j���i�+R��]�AV�kW�H4Δ����7r�uH�V�p_q�nC�g��n�����̮��E��N;���N�	VVE�t�!��������Lo_)�u�!yׇY��JI:����K���Jo��Wd�nq���y�"��I$�$�f�Ul���K�;fɛ:�����o���l�:9��J���huU۲	�V7C:q�+�%Q8��
O��r��m��_e�(�5F��$Qh�R�CS�Y.ϝ�Q�,��޵p�
�9Q�O�!ZA2��`�٧W�Y���y�w���Zx�����E�&.j�!N�t��"�����%�EDi��L�HNL�R$��ѡ~b�Xx�$��%�M������K�)��(X��,R��9e���&mPO͠[Rz���3��Z�S�ʺ ���I:��&�@Sd�Z�u&
��އA��Z  �E��,��\1�&z�m�E i��d��R�.e��7`�"-�eВ�ee�!��U#����=ݛVâ	�HP�6N=xD��2�(R)�@���O��Y�[C����E�����$��&�!��-2�pI���3Mݾ�7e�A6��B�v\�m�_��`�P���:a��z^��X%1RDP� ����n��wN���JJ��ݸ蠩.�xae�T�cd6�!YR�T��4YC�v��өjl��].�§��e\��%�EC).p�$��hQ{!ڰJJ�#rX�vU��*��u5Y��*�ULq�I�*�%�� ���HP��H0lպN�T��X�5l#m����L���i�U�+ZPW�ZPF�
+�h6JD�d9jQ2�9H� ��jP������؆��d�A)�S������T�j3J�������N�a�t3���-KL��d�щ(U�e�L�Z�l��O�\\=��N)�K'ϯы��$�h fXtA!�I
's�Rz�W]z�+)���D1Ti�U�P�3�[}�1����DhR�꨺l�V�[ʝͰ�UB��iTQ��D47��[\N�l" ��E%M�f�l )�I;*l�^����Y�i�h�4�a�A?6�l�eoS����3$Z;����D�I��A�AT�5D�MtN���SYQi/�
�h��(UD����)�:���(i,�A��%H"��N�@�]���ӿYy�Ϊd.H&]l4�R�`5��^����Q>e^��Wb�ݨP0�T�D�J"�5DJ�]�mA�%6�:%Q-5H���BQ�A/RJ�\[�2�\)�kKW_�! HI�~��_�h
�)�o�����S�g�(������~ �$|�?�?-��<��5Я˯z��Gp\�/h84`䫔=wtj�9*�*-]��T�n�z'KA�9����C����
��-<���yܵn�2D�њCf�M�(�M�u�*<�˧e]�x�����ڔkF�Sx2SV*��\��8q/B�7p��r�N=�w��bTv-�͙W9k��8	�uN��^;��S�5]X���lKJ4O*jr��Ro_	;��^Dذ�y市Z��hunī�2���-��~C&ţI�oF(2�T�8����̕����3���W�J�ř1
�OIȔnqr��kU�N{�z�zV����!u��f���Z���/�G^�,#X�i�!�R�G�F���hYkkkQ��:��0���tۥ�Y;�W-�JKuf�����N��G�ϡ*�Q<w~���
��޾��W-�<3̾�=ֵ�X9�Zy譍��a��WC�3���y��8�R�s��r�e�u�U_u�|�U�'�����[ܨ彘Ѻ���-.];,>���7�Y�b�S���*�����V���W��`x3��@ˣ�3T�U����ѱS�YLܼ&s�����ȸ�ȸ��1��κ뮺�:뮺�:�N�뮽��뮺㎳��뮺����]u�]u��뮺뮸뮽::�:�N�뮽�뮺�뮼u�]u�_����]u�]u��뮺뮺�u׎���]u�]u��3��뮾:κ�Ӯ���]u�]~::뮺�~�_����~�]u�_����]u�׽��w����'�L]Hm�b�suo	)]<;Xzֆ.Ꭺ,�E�-�%q-��2-kw�}�q��2n!�z�!��.Xq�>��5�8�WS��U��M^���N�v�^���p1fK"V��d�ڕ��f�ne)�T�Ug:��z�i�� ��9�!��h�ͤ��f�p�7�G���LoE��V9��<f�
�!о��aY;�J'{pc�4憻�����.[��YԲ;b��SƷ�gURSd���)s��0�5���e�q�l�(�Ι��w.+a��c���J�W�NP��oZr���g�B��W!�R�vY�֔�W%��֫�g��9�_|鹺�I��"k��3Vލ;�r����:��Tǝ�C���t k{��b �f�t
��RZ�����z��|�ح�UlaVw�.`��>a�]m�s^f�k
��<��D�$�f���׫2�k9�d=rͳ��G��ea�mh��e��n]wi�*@򲔇�؅ŝTʥ��X�T��޵��kֽe	2)X-S"�M]���d`S]����0]k��c]���U�]�S���Rrm%pV��5hj�����o!Ul� �$�[B���d��fSY�un|���}�ǷǷ�������]u�]~::뮺뮿u㮺뮾:뮽��u�]|u׎��뮺뮺�뮺뮺�u׎��뮿]g]u�]u�]u��]u׷]u�_u�^�u�]u�]g]u�]u�]g]uק]u�]ptu�]u�\u�^�u�^�u�]tq�Y�]u��~���~�_��뮺�:뮺�뮺��{��u����;|�k�7�^�ּ����C��w�йDb�(�
!�\@@d���Ѹ�0"�^�w��m뼘'�Af'˗d�T�哵w� .P�4B8FL��Z�!����7�bk[ұhb��z�F�.�ګ��Pݾ��B�QYPmY�Kq�r�&g�3A�`p{�H�mYVd��i��8��"۹�t���3O6(�
U� ��"L��
:]<�;|k:�^��*��ծ�r�rb|Em
���b��`�ǹ-���ي���$�bLY+#/����-��C��x� $`����q�0�4@�(�����C1.j��2��C
�$�O(m{hhپ'n꾪�i�,h�U��]�j4��{zq�<�\T��e�/k�'���:�M����:�!�"��^Z����b*ŊE�7�\��S�������jz�m]T�wN�Y��DDeK�\�kiic�rd�.�N���5����`C�[�.��<�F��܂Nx�ūo��D�y&Vf�|����zvm^@m*�����d�NT�]�$���UT�U�󏰞$�&�܃K��5�'k�-=����M�0(r�����E�`0�۪|�����N��E��uN��Ժc�.��[��:�B��*QcQn�H�-��B��
R�<ԛ��BL��.���ć�Q��5/�h�˸#��#���k*�(ʸ��f ׼�jցWM*�N�;bķ-*���k靎QR�y��45�#���&��N�`�YP�Գ.Vd��Qם8�ۯ��^ߎ��Ӯ�뮸�뮺뮺�뮺뮸뮽:뮽:뮺뎺��]u�]u��Ou�]u�뮳���뮺:뮺뮿u㮺뮾:뮽�뮺�뮺�㮺��]u�]~::뮺�㮺���뮺뮿]u㮺�n�뮾:뮽:����|~�?_�׷뮿u�G]u�^�u�JW|:_U�1#0l�ۃ{�w\��i٧x7�*���a�D��.�G�у\]mK;���wNod 7V�]#��5j�Ӽx�g�bA�4Hr��v�wX8�eΤi�{�:��l�U@��g%\:��ݧ��K:N|n�L�*.�yCm�6 mGøv����Ѿ#eU]�(ɜ��]���~�j�LB��РUH@�έW�8Ys\���s$�!�W�㘘��A=���̪��Iڮ�R������O�������k�F��&mr1m-�3�?�\~�6N���=�Keڈ9N^˪�&�0�
.�U�=�1�uVXM��r�2���Ln�+�6�_�7�"�cVp=�U0��GK�����������:�E�j�[����I}��le�5Hf�C��6�sS=GM<�ow@�X^����աF�vѢ��P_7�ĒSX�<�)]H��[��:C���-�Ѹ�sλp��9�'%AWY��;��td����x��S4XY�����% ͐�`��a���*�]�ؙ�IKÔ�gCO�u h�y9�s��+�ÒIN;��b�9���psl���o%Z��9с��bA�Yf�]�]�:��}CC�e�*��
�E���u�(�{D���B��ܘ�u�M9Wxň�sy�|����������]u��]u��]u㮺뮺�tu�]u�]~:��]u�]|u�]{u�]zu�]u�u׎�뮺�����]u�\tu�]u�]u��:뮺뮿u㮺뮾:뮽�뮽:뮺뎎�뮺뎺��뮼u�]u�]~���뮺㮺�뮺�ۯ������~�_�n�뮾::�뮺��뮽9�>����ʰNm�6+ך�!��0h��N^gG��[�4�8t��\�H9��p���;c�%z]��5�j�!򻪂;F�X��}�Cs�8e�
��*(�T��K��%�l7�o_�w����Gهt��+�U�S��wL�Yۗ�I:P�m�����CegK3TG��"}���V����	�h�z���T��׭I�;$֮��WՅW�V�J��o/�]���mlv&P8��t�O@"���a���]qUJ<��0�>}t	�bݾ`��2c[���t�k��y*A�۲�l;���]��i�^�۵4���Ɯ���M*����e�Q���,G:����5qK4���ER'|���y�[c��jS���M��ӵj6�^�2s����f���UK)�T�2�J���o�׭��{4��8��]:�C5+��%��R�M�#����Z���G�:XZ�<J��զ�+5WG�v��\t��Z�Z/�͔�F
ڽP`v�q�a��:{�.��pNZ��=�c��V�k���ŷ�!����eP��V2N�Fҋ���u�'.����##cc##��GGGGGEGGG:�뮺�뮺�:�:뮺뮺�:뮺�:�N�뮺�뮺�뮺�뮺�::�뮺�㮺��]u�]~::뮺뮺�u�u�]u�_����]u�_u�_����:뮺���^��N�뮺㣮�뮺���^:뮺�����z~�_��믎��n�κ뮺�u��<>�QM-MT�5Q�PG��7�5\[g(ґv��;}v�WX̭�đ�*�y�1�j��p��k@��I&f3C5l\s��wt�!�tU�.�t{wUS��ͫa����y�[���ʈ�4ɺg;'l�R�4D᧬v�0��v���Җ7ݜ| 4�uI���s/��kE �������]w!�u��Sr��P�*��X;!�=���FRFک���fY��<U�yJ�lj��"n�5�|q]�������!,�ɭ�o���'�^\���.�}E�n��C{���I�ot�샘��Y��v�>�Աl,�D;�&�֐�S�ǃ��>XT����S1N����YWW]Ӻ\���	�"�r�8귂��`�ڗ3*�����>���+�4�ϣ��2F��P㽫��sr��we&�@Dvƪ��)z�E�X*qP�K �8�m�����B����0V�]I����H֩��U��Bf޾�����y���S|��xk��7]nS0����5ݔ-�d��Y�Gݧ����g]��lz
��a��֧��W$�sa�����������~�뮺뎺����^�u��]u׷]u㮺뮺�tu�]u�]~:��]u�]u�]u��]u�_u�^�u��]u��]u��]u�\u�u�]u�]~�:뮺뮺�u�u�]u�uק]g]u�]u�㮰��]u��]u��G]u�]u�_����뮿\~�^?_�����\u�^�u׎�뮿zϟ9Ͽ;���*���rk�7it��o5c}��Vu�u�9bK��XJ=W��!��J� �a��c���y@���_Ca��5�dG�v|����3��iv��̝�䢍�#a���鞵R��Xǀ�5��b<�iу2L�vp�q����l6�&o;X���y[M8݂I��k<xuG�oWC9�uI�"�ʴE�ҭ��wT�_0���B�8[&�q��ʞ]�Q�����]�Ghn��4��]�&����X�#�A39lU��:�,S��������m;.�9�Hv�9u�p���O���X9��:k̬{ ��tT-&��:�R{�>V	���V�:��!�]k�/^����C�����F�����Mqsz̙�Mܥ�o��e�0L�۽gp1ч
o)�a'�� ��M�mJ�x49�T�a��^�FT���*�gMt3<R\��,,˖��E�*�D���3�hd�݃"�Z۹N��c���u��F��l8���2���z*j`��V6e��^X�淦[�dI�UX�A�ּ�71�ѮE}v��l���p p�E�&<������:9N$��͠{gH]%LH��r=
(��;T�)gF�
��������T	T�a��0�{bU�]م��{�}[z�{���v���-\{M�8��m���m����.Z���F�wᚌ�a�-T��s9�Ww�����
�J�}0���!�Û6]�v+���̷�wn����.eӅw���{-d�wm��b�k�]֦�����%]������_��l]eK�.�N��w/�.	�M���ZYJ�5��+��'1���[+Y�aJT�K���ܾ�#�u���a��P�-��t|ѽ��rY�S�R{��i��Dc+բY����R9Wu�IO����G��`k�fXZ�#9oz��\���[��+;�:�u�9r��f��[�Nб.;��ut�H�q5�*J鹆9n����f
{�.�׫��^���� �fj�1b�_P���^J�@�ISj�R=��Q�o\)Z9n;�N42��n��m�<���&l�*Ѻ������jqb���n^��rB��\B9v��H2�ۅ7�أ�Fکk	3o�T�ˮk���X�^͙��}�f�ꊕC4�p�n�]��:F2z�f�hOJX��l�jG-[wV{����1�k��יE$8F�U��%�\���G�`�q_1(��Вo.`}�F�f��m��Kڶ�9a�����70�j�j�=Ҧ3}�UW@x:��mv@4�.�K�V�d���˘���i[��5��/�;Z3��+��,�f�sWu������ђ���u�[Ԟ_>�KZ�`�8��Vů�e�}�o.w��������54����l�x�hvFjh �.�[����H>l�Ov����tW;}���j���I�M�3�P�����u�R�Nx�%9�*S�N �c���8i�*]�fۧ�h�;<����ɰ!� [3�r��`�doi���q�ti;ګ׎Lwq5���-T˫�վ=޾��;��SD�����+m��G���87�<�SK� fqL����Ehv��SmL����f]h�4�=R{���v6��%��@#�{p�zJ]���\8�V��� ���l��qs�/l@�q�9uǅ�F`��,^^���" xq�/w1������L��z֠!��R6Z�"������u�,�����$+~"H2�^�[�鵶���nh��BW4r�pO	�fE3������S��V`�˯#[H�F!�o�
%��ѽ�c��bU��ChJ��/^�Wch�4��vh�뮙{�u�_iz4cJv(��k/fN2�f�P'�;ف>mvZ��z��T���oQ�ѩY@�\����lV�#�<�A��m���s�󩺔�Z��Q��͡����ٻ���;���O;�.�:�sY�����$_����9/Az	wz��S*�aX�[}���Su6�gTtT��Ιg]_��j�3u(�,�X����Lvյ�^X��eЏN�Y\3GVF�Ң{�s,P�EQ���]:_�.��7}Ɨ`f�5��b:{ґ�3��L.��]o@�ѐP�-.*�t9����AgUX.[�5�v26���WJ�gT=G^d�R�C�C���䙓lrΚ:{ڥC��;P��yկ��Y��Qpdr��^E����R
���F�ּ�bh\�/E�Uծ����e��[�5r�U�ɘ]�;��*�!�d�R�僸��sZ�V튻F�n\�]ml�D�M���-!Ӆ��-���kY�Ә�l�5�}>w�u���������?� �*�m����O��~��T�?��G�H���$��9����_�,P$.(����e�_���i0KQh��w,�s͒Ԗ��9M��Be�L�I�*L�h2䝜w�&�`��S!55��h6�l�}uy6���ϖ!���ɷ��]���6Uŧ"�*j��|��hY�c�OU���b�S�+-o\ȻlgTڛ:m:�/L����r�8,v���ޣq�y��ǫ8O�.�G�wv@�k�xZ�� �.V�Z*��u�wi�
��IS\�Q�����a���3�:Y�
���%8ц�;Y���^ƺ�Rgf#�n�ɧ&_ҥ�	C\��#	��W����	so%�}ȭ�ޭt��jں!���;+Y�}�'=�z����ܙdѳ�]��H���H�ǍMV\��m����paQ�v8��/cO�-ǜ�6nE���wi�]M�_K�����Տ3u�CuZ��<�=�os�u�m��T�0����Z%�[ۜz�9��j�ݙ6U�>�g@/kmq��p��Zo��V���$J�ưNԇ'|�uw�����d<n���ǜ%e��I�ܛ5l��w.]��e��nۓ'{"�c�7ͳu�̹U�_?9 *�F�!5�K�i˕S$�vВ�up�aVMFK.��[��7g0�M/US	��]�ۆ��#�mV�l´�SB���LKe�DWE۳a���}DJjB�F�P:�[�ut��4��t$IB$ңv'K.芉�y$EH;B���W�p�Æ�2�P�(%&���DV���I^tȥLԖ�l��}2D�B������������Bo�&ۥU��ҔaR"
�o���:ʤ1�X��q��1�+�R�2%e�k���^�����~3��g���ҋ
�)im�Tݳn�E�.U����%,�""�*�ZIS-�.2���E��5`���U1�||}}}{{{{{}�gcC�u�� ��\BI���&0�ĕ�P� `CI+!��.d$E	�U��4m��+��b�AM0-�et��c1�
�{�X"������&$Ŵ�:�i!(����@U$1(o.U8�W,Ȅ��S-	��d��vvjjjjj|OggcgO�#���l�m�L���L˗��$Y���]s�`SM
*����}�i2�N"$E�)�Z �-mF�5�)n����~������njjjjt��N�2���9��Fv�乄Yr70p¸�yf(�V���*b`�1�LȖ���F{723ss�ٹ������>���e��l^=T�����d�hv\��*T�3M2T,.R�ƫ�)�
�!��#5<�O�榦��gџNN�2�T��ъ�#
��� �E�U��*B�
�Y1���j�uf2�}B�����B��VT��Re�J��dYB���UQa�X��e����*J�S9$�.�J-<d��ud+"1eA��)�b�b��ƂʑB�X6�,dP�0L+�}�n�nb�f��V�i��>i����:��۔W&�z7���N������j"��,�Nv箝����T���J�F�"�R�M#x�����l�d!vF&XXh��w�n�<p����lH�BT%ԁJ1wP5&	 �l~�i���t��$�F��P��;�gl�����Ӻo5>�2�m�P�^x5�T�3 ��y�+�D�`��yd�1���7�B-�t��{rTUzmÌ�$�Th �X�KT\�����HF���k��p��)���F`����k���V�3/з:\��1��nڷ��l��f��/���b�ۀ�*C�^kfG(��I��3P����SxL�aaS��
^�C*����e3r�yGBM��N9/���>���úd�q�3O�A�_qf��A8VS�D٢�8fh�Xd�FǭV�`7�z�3X�4��J�k&}���q,�%&H���!��V�j'���"�=��۹uf(����-�5G
�G�	�{`Z7-��e�/e���������]Nq>M�ͼ�|����<�᫏��YX3n�X���;��A���[<;�}��f=�n󦜶]h�{I��u�p�B��D��s&伽�������&���{Cq�ڗ�l�Kmf��C#!ܺ%q�JA '��l�oP8��N
�x��ڃ�zU_eϘXbٽ���y&�m:��I�G=�T�l� ��U�M�t��
���� Y�Ku��dTk�9���)��CG�Po��"�dX�T�@�k�{���cv����x�Bs�p}�t��]��c��2��vMN3n
���^]�9X��њ�ӓ֫{��z�S|���]M��E��x�G�$�fҭ;�-��r��� ��5-Q�zfz*���ނ������1t�_ǈ�{�$y��%��{}]�@���2�3H6Ja�A2�2�����tj�s�:�ҟ�!��L�f�5��c��s�	�[�^�q���������Z����5ƺsNn'ڥ51̗�i���1US~+�-l�[�(�k�7�GRP0���rI�GѿZ�k6B'(63l*���"�d(Xh(Q��Ǻq�tj_��Q�� ��-ye��_�wk�����ѻ@�^{ø��?h)5R ���x���l��]����A>���G87�&�9�c#9����V�}�3j�#��u���7M[�H(�$A@@�v��u��iA�:��� �GL�����;Gn�ѱ�{C\�=˼w��;�ո%aj����طw��EI��B5�Ӻ��k�{��k��>*�'��l�Vϧ����C�X���n{��/�O���ne�����y|�X��.ð��k�����
��X@�VR��,����t'��(��)0[e"�&p�����ȿG��	���ZM�Q��4&8O0��G�+i��%-�����t&=����J�n:w��7��T	~��F#8�.o�>޶�l�H�2�Q3[�,��w�}l�����{)'@]�	�S�6�=��vΓ�t82����H�`X�zbȾج�9&|m�j�V������Rҡ�̳30v���-dvXS}ꋀD�Qz�&
�"}e���*��N�%,��{����?c�\;�Q����H�]�x�q�y��H��.��yZ}������]u��zg[�L��.�m�>AX��A9/��4h�ܩY�DW3�>uNe�C+��{/�^��f�s˧}c(�=�.���w�78�� {=໧f��o2t���
�^{ĳ܆E�Fa�|'�(��Q����:o��r�O��`U��(��{��첈D[!m���A�*V��3��9�3'tl�	A7��@���8�:^/ik՝�Or���[��֠��ݾ'NYț}��IMϤA��!���&=L=�ڥ�(ҥ�)M}J{2��Ү%'M%�B��CJ~����mA:�{��O�fϳJ��:Tb�/b/p}6�;Q�./)ġ}�طӻt9��#�+�姹��5�����v�*�R��ݔ�K�x|�P�!�y�v�����9�A(k&�3�����t�FN�AtPpoX��Wr��SA쥐�T��הݝGb����Jn|�~���#�[�Ĉ)�uLE6ߵ �j@�;0(f-tۆ����۷�K��>���9�-Z��'h	1R�-��?Z��Ы�w��㴡����f�yiw�5]v3%�7mb���R�^���i�<��{P��ʻ#�'Iy�&�jg��ls|����1D���-�2������֯,[E�]���(h��n�}�֪��%eY��C��
]JB���B�&���-(c~�@��	���\m. ��@��~|Y�`!�Mb>���׍�тL����u����mI��m���~����e��yv�VRc~�rl��dp���|��yδL�V��C���V���O$�;���4]�{Y�J��0�34ԃ^I"W�ё���l��ru�萞0o�%�y�zh���Q1*U��)���M=l�н��gx=���7wt�t�+��붻7V9<�3�~�3��w�m����ޱ��1�IS$�g#Y��RZ,�#�b�6�3��
�m|�I���wt�s��e�c��]ݥlP˵�n�����y��]�
DTX�����N���lsdQ�����Pr������󤈐
h;fN%s�j��:���^Ǩ��4ʧziS$��Y��kjk~���a=��Y��	��w�M\H|�����&r(i#7��9*S�lx:��h�u���$��ۼ�'H2TU^��K���}���������Sm_�x���g���I1P1�s�m��k�d]�ښ=A[-��i����m����&/�����<��U;%c	��Ybj(v����ӾCO��s7��I�+�В͠М<�����Pe���X�'�T�;y�mz���1�j�I��H��Jj�1�&v�w���w,Jm��=��P�q���>�n�[4�^�{�:��J����a[�l��<�T�J��:���b}9!�fF%sVSg���sO����׹U�
Eg�su�>>׊�/�y���K=t]R��\��c|"Hż3F��+M�������e��}��]c� gv�<����k4��2uI:�A�����й=�2�V�;"��	��2<]�Iɞ�g^z�_���خ���Q�O{�$̢���`�N�CXiu���7y�ެWx��Ψ�"`�����l5�DV�� �C�r�1Z*r�$�U�a���=��L�z\��^��{�F��4̡5G���A��Qd���!����[$��\�7^VGÔ!�v|��#�W�wOr����r��"/H��r�p��v�w,��I2��ɲ�FD�oR�75���է�_c�]�X`�q΀(<H���4վ�K!��n��#��i��`,�k�ӈ2�K,�>�{��R8qͽ5s�����YF��fh0z�7ؙ	i؜x��{_Q�T�,��ͤ�L��wfjy*xl�[��du��1��U�6����]���-�B|��*�j��K�g4�s�����p��S�t������Ϲ�E2R�m FǄf���j*��Q��Il*6��mʤ� �њ$֫W�.���t!d�u:�vb[=�n�AR�*!�J�"j3(�1t���W�Xi������=U�=sO��&槰Vx\��v���^~��\K �Б�J��1l.ֲ6��L�[������������j��
�e#�I��Y�JtN��c�;�{�;zۺTT��z��J��/N�8"X��u��>����{y2@[j�׏�o�O)�t�X�?m3O�˂��c/��ǞAb`��;z���,E�Xe;y�7��t�n�3�
l��H���}��)q�C��OF��(ʔ�Mu�Ґ��;GY|� �u�a�3�GowR��B����A���������9�Fэ+kk͎�S��e[~�ڨT�,����p��*�7況u�#س���O��X@������Ryc,scԐ��\%	�6������s�����#Eޅ��ʽ�@����:q�I��K<�3y=�{l�SE��y�_���� ���k�y^�W�*U�ɝ�s��Nd�:��UŅ���_��}�7Z�b�y��7�����)�{6J�LO�r�m.�Ê�}��*57=qr�WSx��*!���K�֚u&�"��%�ǩ�q��C�w�;HVu�.<��F��������b���m1�<֖X!�^�����F�����O{f��5ű=i;��������0v�A��d�m�)�/K���]�3vm�1QP�)��nь�B�(���r�l�σ2mYj��*��۹Urq�ҡai��D�;ʩ����N�`�<D��i��-�	)��ܪ��ӷN��c^)X�N�M�/��a�c7ko+�3�M�#�&�c�Q�i�bEL&g�)���DUQ��bS���S
Y!�� �l$�a�
� D�IQ�=��fM{|7�j[�<w���L���I\��#��[]�k���lw��~��H��73�VU��Y�Q�f����@�1�&A�-X��#�C��W�E�ճ>Օ_}]��{���V�R����O�]$ �l���ncK�Z�-�*�5��8�����cvu	a�E������V�w7o��ŝ�F�	
�EO���9-0�j���}�[�uvuT%[�e��#A��� �{pz�W�mc��.5e]]��3�����
�މΔ6'Yʐ���b�����F���z�hJ��æ"F�iy�����P��ZOh�6&���g���X��U����/V�	$YE�A$��9먷b�W]�t��-��Rhd)Ł����^������Y���
��#�S:���[ַ�nr��*�^9�S�9i��xr���^/�����z>&��z��ʮ<� �t�]a���W<h�R��Z��-�x�	1�F��@�4�����w�|��3@c6u/.�r-[0WV
)�Jk�A8��7xJb�'	v���1�e%��$�UX��G�'Υ���R_=�K�}�K���_N���o:��g{�z��}����{#�faU�%��=s�N��^yP'��l��u�35d�n� �i0W�i*�d`SF��R��<`��fT�5Zf�-
�&�x�!@ƶ��dny�h(��ej��f��>��cʝ9p�`<�ʍ�I��^Q٢�	3���-������3Zf!^�fI�U� W�:��y��KX�ڄ�s
�(
�Y�]����eH�̒�_g%��b�}���0���&?��_�O�L����!:��.�W�1�-G���E@7so�Y�٣�\L�����7x� ߻{jjB����Ř��em��}��{tu��5����ɁP6���6�H�6���E�hk8�}�(�C�yD�YaNnTl�����^���f�q �/>��w/RĮ��4�}D�����c���剸�̊�+7�Ԗ��]:Y�}"�Prvx,y�� %�5���&gN�:�۾:��ws�����F�k���^$�)�eJm�Y�}�`k ��1u
	�o;:�f��y%[c���rm�V��{MwkL;��F!u��V��έ܃e�43{bY���f�3m^&�ѭ1lbjYF���#��퀮��hukPM�w�ƸG�T�\�\�?��˳�d��,ǖ�^�.9�흲�n�ti��J�R�w�A�.t�c\���9Q��}{�/wq
�I��Һ�xK��t�����u��a�_T��Z*oa�+;�V�YK�Uv��:���w0���ǥ�a�:�,j^ށI�b��u�y��ŝ���ܵ:�\t������&��aM�CT7�O�"<b�#t�s��W����ߘ#J}��-�-}��f��;�t�5���bMAo��̮�#�5X�g�22��~tf����w��F�t�G�T���n�TWC8�l�� �4fW4r�+h�Kl�˵�g'�y�YI�[}�lo�0O��>�I��{{�
)>Ma�;��yMY�.ž��<�����o��ˎ�����*�6(���� ���ZM]J4�u��H�߉%D�Zx�*�N��+"�hitt6���j�C�kF�)��fUꊼ5m��ԉ�yJżڑƬ��ۺ����F��cT�)�}L�&Ua������ v�r���]r�T2�+(l�~������L�G�����rW*d]�T�+nVCݷP�ܝ�Y�C�Q�g
&�����*�!�8���{���/���w6X]j7���w��=���9��;�Vw5���S{����0o^��Y;���o��|�*�N`�ԋOi����a�w��P���Y�5LQ�q��7:��3:o]]������\Yy���r�o��n=zG@3�-���M�ꏋ�3p�OEFf�ܢ�]t�5���:6:�3����b��/�)Jw7�`n�Z�v�����N�rwp��@P7o�[��W��}�j"![R��;cU�F�.nԒ..fluF�Wcp9{�yn�7vd��'I3Wh��]�D���.b���f�b����I6������7�%�5Z� �Γ3� �^[ùEg*�ʎ'��w,{�Jw�κv�]n�I#�V��Ym��kxY���'`�삢n�j�P���/�U䁽�4�O���A�&�t�<^(s���Ȏ��UXv��&�W��G��:��l���Ӑ�K��ˠ�Fބ0^��:�[���k��ܾ�� H7��w��Ac��AO6��!aP,����ז�`-�����=�?__������_Y��=����
+D�[t�L�����ʍ���F��a�m��k2ܵ*)�	�_�OL����������~=���Y���UV(,�d�R֊}��褀��,
����(���9`�Q�}2df�ggf榦��I���ge�8N��V(�-������«�b�;s�q�-)�̣JTm*���%����=�:�����ۣ���gק���z�YV��Jʘ�d�UkT��2���eA�i�͓Ř����������=���e�p啨�l
��Vҕ�.��XVkkE�b�E�f�2dԳ���ssSSS�vrvX�=�*VV�5��@��&5P��I�����+AE������E5��Ұ��̕�Y��k[m�&ڋ�a�8�J���֊;<���40�1�ʘ�3e�Q8�+�T��)�*�R�غLpQ,b�k1��ʞ��6���`��4��A-/	w��[c�}5��ISz�Q%]5�����uE���}o"�W6�dy�;��uΰh΂��+���?8<a�f�W�<��s��R ��Ix��rq1���`�t1'	 w�<�xĎ��V:B�Q�a�{B`�Ml��v�}��� � #�~,��s��.���A�����w��Di�����O_�;�3y�oWN� 6�~I�2i5��&>p�@7%`�=��2��`,� X�A�������4�g��d��Or��>��0���������8}%�R�qf.�b,��t�jv`�g+WWklw��z`�4F~�7��P}�����3F��֦�~`U�3 x�@g�&�����8��ʘ�:�.��D:xj�7��mxx	�x��w� ˼�;d	n��>��xg��ɫ�Q�4c/*����!g��2��ؘr�.�M�t��������<g���t�p(s�^�޿d��T���߾u��>��pR!���	˞�L�7F^�nY��]�& ���H�A)%Q<�H��E��Hj��<j�x_PՍ�C�NC�������q�|�{�����%����-~�=dzU�	�� I=.`q��zp}�8^u	��}���[_�VIs�����5c��!�>��_Q`a�5�T'H�$g�?�Q���Xdk��A���?=�<���9�T�v�w	�]W\���ݺ�};0bU�SM��ǹ�����ܑ'�o�m�Q�"�`@�q�I�o9v���EEMpr��Z�	�����`���(5��{�ǜ�b�c��-5ئ�4�ȡA� �7�ǟ�<�3�����u:�@� ���R^��cߓ� 4�˽b��Q|� C@x�ft�����ۤ 5h��0>oH�LB����	DQP{�Q�|RϷ����l�0��-���(<n�9�4��x8�$���b�s�Xo�@U�1#��"���À(XD��XH�Y�j�gh�
i��(�L����%�,�����c�`T��_!F;T
 h�F��C�:L�y���Ǒ��k���͹���dk�ޠ�-q� &p�ۏwvH�T��e��T��Z̖��*�L��>�g��p9B ��r���:dA�]_�G�����Ƕ��鿤C�B��l�=�w�tB������<�08�y��	���)ジ���E5KY�A����;��� ��^X�����ʻ��}�#a}:�	���O���%���� Z�A�BS���U�L/|��Uo�l�X�cή�2����p39���������?{�F�o����ͻ�nz%��9w�˧¢_Vej�����kc�1Ԝb.W���!K���^0M����u�~�0$��t���T�dr�T(d��9Qw6�%=�x����"w2h�n��J��F�Kv�b�̗��ܓ�9�_|�ŗ����ʄf�טB$a7��Vg���c�6���^N���>�f�墪����Ǝ[۸:���`�/�hLL��t�Dgc�-g�l��rѐeeY�$7EJ	49�]�iu�~&D�HČH�"��w����H ���S�(Z��ۅ�Z���C��s�
���s���ׂ�;��<�p-g]�̛��s��<�#�Ə�PM�H�R�l���e0�	�.g�u��FX���	�y�w5���e�U�ʙ�kC[Ɋ]��]�X�ϡF%f8�`YG��/�`�{�o�Z;W���>�������xN<c��K�$�{���m	Sz���_b��-C�Wq������/�:�N��u,�}�p��������~W%�$�i{����� ׻���*:C'k���X!��)�
s��;� ���W�_ Hw�~W�<j	��>C���H�Zb;�.�0$g�� j��v��aX��)4k�2܌I��s�a�5�ܰĘ����J�ؙ�_ z��9 .p���;�J5�!r���q��>h��j [�W�7�}�А��C�L��yDK[�D��0�q���0��)�!14�'N���2s���Ж����d9��S�;;Q��n<A���P�z_3�h2���6y���FP�C�
0�T��
�:�y7&��j����@��2�o~p	�����*J�
z��L�~X`P Q���+�Y_��_��t��6Ʋ�{A䵌�#%p�,��[W��'�a���o�a�V��P�c7|��l��GTXZX���������f�U�k�x����B列�/�:T�.r�qv)���v.�.��;5u_^�jJwڜ���B�h�A�!���|��;�9���/C�~�����Y�~a�w^k�<�(zr������_zBd(��`g����A.�׏�?$���k��J܌ͨ^�t$t��z�a��G�zl���@#p$9�g�?[tj�z~���FXu�M��/��Ὰ�wbƿ����+��+��8!����2���{���6�JԞ��`,��>�A�3�j7��B���1����Hξo��R�w?l�b���	�p<]�`��_W�O�9\���z'Y`m�J�cm�R���)Y��D����;H2����&�� KVyC0�&�.|�E�s��mD��'>�"8Ǯ���d���h����@H�����@z����њ� �(~����F4�.�'���H�FM7(tӏ�hd\
3�f\t�P] f.�¾���!��0l�5�~:@����v>e�l�ׄ�$7
l�`�L�{Z�矛º�@M��*۫�<��C`/�B���PθV<�a�(>�
�&R�=o��ݦзQ���[���q�<���j'�d�LS�7�yۇt ���0l����J �(xQJo�fR���P+�=��A�VFaJ�;���B>	�nO*��=$��I��]J$i�;?SU��mW���1��9�0Y�I9z��o:Y�����V��!]��>}�d�I�ņGp���u]�Z)o=�Mpr�o�aȎ9�݌�-lf����R���%�N�Ø��59�O��y,�	�),�%�YH�����Θ��e�j�o��y���+�~(z����`#�_��Xz�6��Hh}����f��WB���Wؽq��M���� ���V�1����]�55;�A�и�_ҩ}��Y�G��L�uܿn���M�n�Μ
i	�+�y4����X�p���� �f����Z��HQ<@�)��xyy-�</k_�7O���1�k~�3X��SM��'��;�I�C�Npį�=ĞX>6��N�Nvy��+B@��&H]x�zG�|�ɧ�w} t8F[�F���;��7��g��&*:����#�.�.ce;�?6�U�=N��H
,;q���{�ډ���!���@�D4s=�@�-�6H�WgtRꩀ!?yo;&f�(3�}�	���	ʲ}�dE�)��d��}��:)�C蝴2�]��
f`���	"���$��3�����@�6���	+��� '��G(	�P��8CX�F����ؙ��G�{Y�c�v�������*I��՗���.�q�*3�x�֭����6��-<�^�<�������� �ɀ�I\�����6jTJ�A���Z��qc2��>?���;�+���xJWS�Y��yM��r����l^`M�Խl���}���0Ý�8.� pR�����&6�K�VҦp��t�ޅZb՝��L�
#�w$�
��Y�.�Ir,�3O.��w����xVM�vܘ�A�"�8b���! ���̞���hW��Ś�:�=��c�}~>�����ԊcAt�=�t�;^;���	���׹�ro�����4zD����R��X������16�Wo�:���h����U�;T�1�~�z�=��}��i�)ph�q_�96�b�¬��7O�Ĝc��P-���Z��<���>Ϸ,1*ED)jD�͍���2������`�	�o�n`.�!ϟ`"�GϏ�o�Q�}��t�6L���-)��ՋDq���y�z�}�k#�X�\�f�v�!�y�j|��Z|��J�%���x�6Vu�g:9w�;�oy_������T��>�Y���Z���ˍF�%��"~����͑�ޟ?��J����t��ݑ]�%�U�1稛C��hc]���QB�/׿��r�Tg�h��}�?z��	Qe�D-�>�	����`S����V�����|��T.w".Y_$x��7vk�{O���;T�*T{^��������I��lX/t�5��ּ3~�ɼ�'�p��l���7�n9\�"�^�����Mlf�}��9�����m�l�����ݗ�6�����
f���n�.�k���n��:��7����ݛ�w]�}��e�ã�q��_tm�7uAQ���DY�l�̒y{8Wu^`ۦ_N)[z,�����b ����_�F�]c����\5�r�,(VY19#���6�S`�t@�H�nK��JM�ҙe�B&L�d| ����Vm�ݞ�\�(��$lN���0��j�������+����狀O�b�a��}��m�-ܺ�G ����8�t��C�ld?H�鴽S��5����Ɂ"2(ytX��5�b�wr��gL;������-~��o?~<j
#�����nқw��Ǵ�)�b�<-�,��	��/o�؅>�o��[&a���SР{�G�h(�^>��]c}XE��������ȪA1��m�% aݷ�팀�ڌ!s�T�~N%҃9k��i���D�e�x!78����˧;��k��A����6Q�����3t���5/� �B���������w�&2+��&�{[��6\X�~û^����u�a*��DB�����:�Q=��"7jNa���9|.��~�_m)���]؟Nd�Pk� �Ҳ�W�������m¡�>��=�lR�spj},�1����U!�#<�F�/s������%��O�oF�z/E١�sw^��TB���� st�V��N���^���:��"�jckO�К���ͅk�&Q���{ߜ��i����u@rM����n�����j��i�s�E�)m�����:��0��`�~�i��[pMVS�`�S��4xd�]W)Ev��]2�҃leԏ��v����d��.ޞq���S3n��_D������BD@�ϻ��~����F�M�A뇜�n<c�}�.��S��E\.z/����+����5�u�*;�� �-���`�(|�[�&���g�w<c���E�<�G"��њ�	�.U�fS����Tj�o��W�@����
A��H�m�a�&�5GE4�.�qKǧ6h�3}�L� �s�_��{��1�R�ҭ�P6%�������\�9`RC_-!q�-�k��\��P�(ug����SK���]�Ā?E��1��xebȪ*�ش�{q8@`��7Q(N�."!�T�����#��+'˶���I x�����0V4�4'�0��/�)0�`�oe����ޣ�@(� *!I�#]���?�	��^ "�ˁcIF1}%�<�x��?@���FI8%?8aso�d�_GE��N��F3S�ƙJ��v}!�a_	���53O��W�`�.El�_�����0���ٚ�����P���ߘ�#���:"�zG0Fv.�{����ƌb��'�kf��]�b�ܔ�~WB�v��dف�U1�U�],�p�
��$���&\��K�"g^�	�lA��S������7_j���YN�].����d9�bR�O޵��K�%��I_s�����u.��أ��݊q͊��'!�n��Z�F�.$oc{"S�PJ� ? �P�$bF$fH��|�>���<�7��&}�]d�0��<�/TM�@�-��02��+��T�y�F�¶��5q�3�G�F��\�s��ս��I����fܙM7uϦ����b�s�ǪW������
:~�2bB��M1�4F9��Xt��a3l�N��9c�c��r�;�WeƵM[vI�E���!Y��w�_|��~�:����q�|�����+��/��=:�6�u{:��)����'-��6�Qze����~�hZ@�${ՙ�&Q�pw�S ;>Lz����X�&I��~��;��ۥ����rp�3�&�����>�
�CZ*an���dT���OR�f9�^[['2-��{�sw��2��-��e�1U�RQ���]�����A�O��lS�;O��^�3�[�O_)$Cr����D� �l��=Q��<�36c���Bk�ꃡ"y����!�=�H�i��XÜ3�0u�8i.1㸇�2�Ii"�ot�-1�V��G#�mݷ>L�lj�\�/�{�D�r�<��O>48g��?���]��J�����D��j���}8�~u�u�A�(7B�W�ϐ��$�C�{���̅Ԩ� ��0�a�tr��^Z������3F*�@�MI�f�;���\-��#��M&���Uh�A]��J��F}Ie�D8���D$��������� �x���Ĺ�񔰒��"yI����5�~��������YCg����'fm�"HJ���,'} &�� )[f��P�q4�����8W0}#�"�-6�3׼�}59� M�̪Ҹ��<L�a�O߱o�k����L/�v�*fSw��2�����Uk�M`UY�ݦS��u�b��z{��x�¼�[f��1�L�RYT��P���(��ѻ�O$��@?y�J�OgX���v����|�@�LFS�\l��L�������^�S�؃>���|a]���ҍ9�.���De.��{ɱ�>ay���~^-�ȳ����DHՄ<ݏW��|�d����4lg����_*`�;�;ؑ���Ư�l�E8�������-4��~�[5���3s�M/�ou�iD�^�bykY"�����Xѹ�F�e�h��D� �s����>9k��v�B;Hr�sgo3N�^�ny��yu
�ߝT�9Pk��?nhI�Xj�R���Sk%z�Oh=��g�:>��5��XD�s��T@{��.���q�˯����rwr��(H�AO�0�1�@� 0����&�o�N|2��p��lT6zqr��ݪT��z*�<������������\�rݡ�Wf�v���,e�I�i �䫸iA�<�	4Z��c��,�$ܱw����Υ�]j���e�E%��M%KqN"��v�h5��$�xe�C�J�m�ʓ�k$T�3���%ImU�Y[���(uշ6�Z-�j�+��0[3�WO;�Q���4�3Iϓ��<8.샦�:�[oI��N�!߃v����6q�y�z' 3��I;M�R��;�4���{��-\�Bo{f�gB�Lu�����7607�յ�4Z̻�30��Ѭ�H:�t M����pҹZH�.�W��0t��z�/n���9X���&J�{�W�U��@�M��c����MkU���=�&���\�[R�>��osΠgsE]]w�1"ۨn�h)qnG%�Tm+�ov�D/�틣�����]���}�	5�_Z��:[s�rö�@��t����7u�1d�;utK��Zb�3��j���(�X�w%�u��ΐ����r�Z�DSb��f�<e[��W�D���}��N��:u��(*��o^ �-��.��f����෷����k^ߨn��;�?Of	b��$�霟%W�����Ps^P&��`�.Zh��]�k(7ql�[��19Bs~h��(�T
$U�tۂ�s�Z܁��n�]x�$�C�[lB+���yT$^-F�adSUG\�B��M����/fc�3�x�ue��+�	��=Ք�r�mNR;"Q���]5K�WH\�x �(�nwfL�+�"���2��t�З�n\�ѕ�/����-^u�v��+�鎠�/*¡��6��[z6�$h�Q��ݡ�bF2�c4��×ƣ�s%�\�c�rP#���ˬS�޾�;�����>R;C&�-0�j�U�߻������2c��y�~���,p��F �Kz�VAju55O.��>�5%ܨ|\	s��Y͹c����S5�Ho�,����雚��z�+�2�1�.���\�6�}e�����:�l*��v.ˁ�5/�Hڜ�IJ1qۼ[p]^�T]ۤ��'z]�b�mw��;�|�`�$��+;U��57��M�T�� >�2��0���/�.�մ��5�F[F󰰷�b��{�Zd�[3.c�����)J˽a��	�{+0ࡲ�֙�Z�]�o�1��칄��2�:�T$j�T&����[31��)�2�6(�������:��|��\�y��!ֱ�1�j��,)yu�iDm�m�ڔ��e���>;z��S�5zrZ\��~�Μ���r���,%�̫�x��27j[��\J���{g�t���{}v�����NZ~b�y�aj�l-��^"Z`���бJ�v]�v�I��BRA���a�)�Ce�A��2�m��$�4i�T>.���`��J�a��@�Xn�0�UMR���Z,)i˰ik���)�
,9���Ba)A:5&ZP[�-4(R=�BJ+�h6kȲzBu0�TAL�)RL�	�W�tBM4�eO;� -E�KX��T�S-UNᘔ�*�t��sY��F���ǧ�ǧ����Ƿ��G�_^3����N+<���f�FШ)T�Y*�J��������B����W���o���8����u��<~}�+���a�6���N�T�ZYv�q̪��"�n����-��dɩg������u��<z�{l��D����%X��+
�*T��������Ǐ������믯���Ǫ���#Y��*�X�B��%����\�m��e{=���������G]}x�
)||�mE�h�T^3��I�����f�YQcl�ɍ�
��S=��^����������u��<~}zP�Q�D�5�mYm�P���S{f0uTQR�a�VBYF[E8�1�V!iQ�[mH��-��(4�����X���Z�R�q��a�DGIY*��kSv��r�,��am���W��$IE�h���͚Z�
��1�Y��jm6��ߧ.k1�M&j���Ğ�ĥܞ*�]E��{u֘�P�g��n4����6;SI�.��1N̡h�2Zp	P�B�a �f^*��Q�[u����n�d��P?�#��RA��!�����|��^V�r�E��B���l?���R�o�<\M��(]�vR��E�=��=ӦE�6����t���^����j�d3y�ņ�t�%ƥ#Es��D��gɅC�ñ�l��
S:��߲���>�����ߣ�I����@y��'6ϛȔ�y���1�[�{~�;i�V��f�&s:�.����-}sx1�z{�W�gu�P�O3�oql�j�jg���Z��"�^&��l� ,������-t�3;+/��xzn�`��:�x1�,R��1��Y�	�.1��FI�	]�˞��C���/�vwg��qQ��R���I���ƅč�W��q:.<�C�c�ڑ4�-��T�<5>՜濣�YK踧SG
�c��(׾�%�]��g�O������f�d���!a9&�I�}�c�y�7�>����P�3鎦Ī�l<�c�zg���;l�al���Z�������p�}5[��_f��)5�hX�d�J�����W�H_)5C� ${��$᳖���~��6��7y�g��>L�-��qy�_b���4f;�̘cM;,��)϶*D���h:�e�}�+	�x��Mr��W���f۽z�c�m����c�A]Ј�m�'1�啻��'/V�C������G��y�|��Jfi�$#h���-�08V�1T�n%�{���rÃ�ĩ����W��N��Ue&���As?�d�T��$@�"FH$H�0"��<���߼���+xϟ1��t.-X�{�̨f��YW)co`�8��M5�ٶ>�����z��V�J�SsS?t^={5�L��O8�^;�}�+��T�d�O.��/>��40� ���f�Fv������5Z����K6�&�p���7B���.�ɀ�t��1�wg�EȞlSڅK�"�:�	|R⛃��G5�@������?A����GՏH�:֮�WN��Q�xh���ݟUo�:~�D4��IC}	}9S� ���vw�5K�x�M{zj�*~i�w���1��mxL�6>��<M!�����%{�;2/ᢂ��&��I�E��9=	yl��2�C�b]CM��r�v����L����[+	L��	,}��K��=S}@3�{��x��Q\��'�a�5|FC@7��.ߌ|g'7>~�~J�qlG&���(�5O�1�zU<�A�މ�K,N��W�X?|�({������e���I��U��R��x~a��z��v�H]�q�Q ���<KΔ�楥�^.`�G�x�1�Pֳ9�GA��[[�8\�E3p��{�1\���F�o���i�P�41�����8_��m�������ʙx02��G����C޹�A8%l*xi��s�'	�5�J�n�&/.���Cn�!J�hZ9k>�f+��;�Z����Z��NW\���`�9�BbY.Wmr��;��s�mcW��\�C�[��bwO��~s0���J�#�@pa`aIA��!���!(�����{e���xk��[4?w@�{W��H�$�kŴ��>@�[^�<m~4�m�a�������T8~�"���Ԥ��B�S��T%�G~�&��(Y�G�ɘ��=�N�uɹ��߳�1}�gZ��6��P)�`%�Ä�PQ_�s^ë;~�u�[������r:����Y�3�B�{�n1Ǿ�v�\@7i9f�?r���iQ�v��k �������'��5
�
5o���D���#a�>Ll�!0qq�T}2���V�۫�+2C3�t��eC3���:�(��Y�|_}�+.��}�lY�6Vz�8�׭y/��.F�/�UnL�nF?dŶ�=6�*:ϻwSu�V����8~�l�j�R�>.��B�L��W2h)�-_�9�f�9�n����w��T���p���t&q=��,���<����G2�B���=\D����'��% ���o8�w���ֻ��?�<hw�\�_��E�����|�?�;��eP&�����jE�*�r�k� MFsל{����d�ȱ
�03P'w]��d/��i S�����*��7��ɞ�_�d�3*��B�w�C���ӊH�ʓ:�^�a�ZȔ��;���Nu�;�W��uCz��<s��{��hf�s�U���9e��|]�E䧁E�.�����$f��s���JO	�``HeXdHa\�����xo����w����U����ڴ���|�?;X{a>��zg�"|��C�6���ǝ��g&H�ƴp���3O�m��.vGz^��u����{zu� �6N�8#���moW�G�|�Ѹ���E�t@���a��`���!<��`Y1>o<���N� �:�W�i�oԨb�3Ǜ�c���}��Z���j��Ze,G�-��haˣEv�^��<y�JT!�O�#%�ۙ�6[t�\%]m�	'����ӆ���ɇ�e��d�%ަf'��M�[z<[nǀ��$�B��ڻ��d���w����[������r���ڤM0����	в�1n� �r�Q�Y�*�]Kgt��"�c��	��)Tl�ft��H�\|�{Ԉ��vۘ䩻�
�HxO������f՗����i)d��8�q����zp x�qoއ���R�۶��1�;?d�L�Ԋ�~�Z+҆w(���0Ô=1�~}����[hp'�Zq�����-jtLH��Ӎx� )����kNc���5����&�{x6?M�%���0`}��G'�1��%Y-z���k�(fI�/<D�5\�o-���ŋɁ��&�	(�@�â<b��d6�f"��*��榡u�R�A¼�>�.��k\�����a��%�����wr��~HI���=���k7�v��k�tC��\;�73�����W&Lגby�g	X-٩ռ�s\��3D��2�_T9��BBK%"�&�zۭkN���6]:�=H�$!*C 0Ȥ2��#"�J�w�땞�XӀ�Q��L�P�(HW�
������d�v=؁&\ZV��}1+�)i6-��ﾝ-R��f짵��Iˠ��z�=��ζ��3�}n=��ۊ�S�L��þ^DN�"����0���O�ǋ'�����W}�4�5��U;jQ{>��=ˢ�拏{���N��"aA]��2����d靵��x�q���H��j��l�lOG}.s"�#�"k�x�c@� 5�KT��W4����xu?���3O�=�4��±�lw���`U�jg�6Cc�S�Y늊z�k*���jZ:���$q>zx�G~����叾�$�󌳲*]�d^d��@��GuDc�a��u+� ��]{�lc&��9vl��=�Ϙ@�J��y�yF����{��6$�!���^��,�C+~�����ȱ�r�zR+�����z������������Ѯ-�v�I��|[�.P)6�}���I���)��%�|W7E�W��t7�i��w]�^ҧXS�G7V�I��[��!�������
צM�_T1�P>wș�WD���ɃW�_�r[�3�
��v��ϞS>�����ݷb���DT��ygVT6c��o��P��f�ᐳ�٫�?P���h@�I H�.w<Վ앂���dӶ�X��<��<4��i7^���:��9�<���\��g���Nw�]U	� G��G�%C�"���#$H<����ߵ���4�������N�f0�5v�M����k���9@0��[��ж���_Wa��P���X��~>���O"WR�>�m�FsIL�+�1�"w�_.*L��O'Iw�x�xa�ò��� vwE��g�+a�������"�<����,�V����ضЁ��sRa`\Y�`����P��zs2�N��Ď��f�~�U����x�)�q���]$yg�+	����RE?~�{���>v~�}c��;�K�?�_ˍWo���#)��{'%���������g���eq'��Y�E��b���a!�q���
2棹�Cn�%��e��+=M��(��˳[oc��_����%�����5Ue�t�a���[Yw��Ѫ �YR{��6˒�̠�1��fq�ƽ�=���ɱ�u�I�I�@�\�����|"u1\�_�~Cg��>]~�SF�z�5;�1WN0���%.gXF)��4v�Z�����i�}�L�-#�Q �
���dmq���=�|��8���=�r����d��e�t�w�3��
�au��ekdg3��!�"ӌ-|�ɵ� 0	Rw��M�G�m��8�Mvg��X�s&�ԴTE�_���T�\�6�FPR�x� ��c��<�!�W���W�u����6��@�K�p��1:��Q���|7�3t@ꆷ�J����v���r7v*�;G� G��/ a�^Hpa��`@y
%(=�ww?��O�o�p�R����&���#��F��P\�]:Iu�=��Z{�[_�**9*=��lZ���;�*�6�i��I�*�	P�hv}�K�x�2����K�C�վbT����'��kxN,5�A|�P�F2	;B�Lj߯ώ.X*�T8*�<C�/�r��7;Wo��]�Y	> ��񙷿$nq�w�'��J�ޖq ���#���v<.7���Ø�y9���>�����6+��SPzg� D�jBM�F��K_?}!�ӿc�C�ق���E��x��1S����	�ۥ$�G 3X0`���ޝwzn�����f~���ei����[�m�>�,��}��^�n�m5�0�/���8r��cyP��L�+��1ʗ����[`kkHy�eCP��9�瀶v��wm�L�_��GN �冁,����)��0=әc�����F 	��R�R�d���Hu�eοz" '�������z�iQ.d��,@�Z�`:�vV0��e�.��e���+���gU<����}u��}�L�P�@xῢ�
c3��/بj�(�>2��.��E|o��Ε0o��YK"�[x����&ô��%��/\�ej���ȸ�*��9S#3,��}$�jw�(�-В#H � �"�U^��c�̬T[6�up�76���N�`�o{(Ԗl�����d��5r8z��Ҕ����G>@���dN�ʡ��ȧ J�*'�(��!)ή]�ލxl��ӫ�5������LC��q @M��;���AO^O\��Sa�]���ZF9GE�5w����'���� ���,�F(������1PyH�H��cRY�����8�w��;�DïQz.���fe>)x������O`�X+cn��8>_}-���~��{�k�D%��)�Lq�pWE _N��6H�
�	#$i Ăf7ȰM!�[�#�t��:�e���w�!�j�-�?	��+��������i�e�s�R��<P�,ץ�g�w ;eR��K�4dQ����G��]j�Q�����~R�2>��\M� �=[dHYb������	6�����.!���������b�y�>�w�Õ�w%=����4�\����Y�'z�p��� ��Z/�F�އ�>��D����l3����P�Y"������Z��~���P�H��"����y�( �Ĕ{ �������Y�L`��Z���hvg���y��v��τk�I?xj RC��#����O�'�C���$��7�0�y
�J��oK�]e阯fE�iaA��ݪ��am4�up%KlD�\�����7�r_�����"�ޑ9m�d2X�[�d6&H5R�;faJIqZ���7�ѩ���*�y��TW3N����\Zp��ZL�LS+�<��wX+A(���P)/6�m�$��d����H�)��.��G|�����d�$ �ȡp`P�Td�UN�HfJ�>�n���V>ʶ�J'�	J	��*�j��s{l��~$�����J�7��fe�*J���uhТ���MK�������#�ƪbH�>�r�	�I��B��m"����=��6�ј�u&tk�h����Y��h�A0�h����sBhy���7
fiq�܋�ꅮ��f٫�tŦ�U��3gU{���C�+�Ϯ�?EY,טּC��2��}�C@��Ӈ�P�R��B<��U�/��.��|�4f���r���S�Pc!��8��bR��)��Hi�)1eg|��N�Wi�-����;�-��W�����!���6"��5
�⍂����m�!55�ލ~�
m�<��k	��P0l�/ׅ����+�s�'=�M�C�֑�BC��V]N��9$�³�)�^==�i��y���Q�.u�j; ~k&�>vLO�Z�l�kA��E���/���P���}��{�C�8P�T*�E��{��:D�|`u�;����O��H��,6����8�Ws�P���vZf�l�{����֋Q��|��p�PWyQ�H ���F��T���w�y�YE�z�4�3�rj����9����L��(���Ս/������JdE�q�h�9�J�ȿ^�c�ۖ0�/懶X�D%T�w��ӡ��kV��(�i@�޼V{�L�m��j��9$�9�rr䓑���죝�q�����S��F Hd���R!�B䠔(��  Lg�Hq�a�˕Zҳ�V�+KĂr�]��8����ǜgM�|���6>�8J���p�w�G|���`-#���"x�$�,Z@3�޼M�[���fvU48�2�*���G����Pjq��(�5�ْuRY��Ґ48�'�蒽��~?]���u����dz�$���!��(B��14��G�>/��6L�H��M��_ͯ�˔oH���8��>1�{����*�V�� ��#ʲIp�@vY�	 ��K�����=V�}�������^�� jRR֭J0y���A�K�M�#�Q��ǖ׵����|v��9�m}\��o�ݻ�}�JoZۗ��I�s�
X���!PQfh|��G�����%,z*��]]�O�0�q���B��G��!YN�(���af6�Q�8�4����O�����a��_���V>ǌgá��"y��8ݿ����%���hu�6뭫8�;<vW���F���򰧋�+|�>���wOy���/t1�o�v��,�LDfN�߾�.aNOۚyT��!�R��V;08�YY&U��e^�V�A�c���B���G��@�U.R�
'cw�hO��n0%L5��T�,7S�P�C���'����A�X��/8:�i�D�1#�o$��m;��]���҅ٵs+q�f�>�y æj��Pg)�Q��!�
/�bD�o�8�RR�l���n��V��U��S.q�M�[�cT��m���z���NC��b��(	��Y�K+��\\�.�uv⡙�;;zPF-nuPG�ffsˢ��H%��]��N��e��+�u؈�:r��d��=RwY�u����Z6��l$$��-��+��v��:��W0m��WX�Ba}ZϬn�����g�r�{B��͓��V��]g��;��]�~��F^1��%]e��h��X�	~��}w�X�v!Y���Ć�!q��K������v��&��B!�bj�;��t �|��V��gZ���#\��99��]�����z&��+�V)�j�o���U-�Y0S�-�0sֶ�=)�Kv������:�k�$]+_e�l��<����%��b�]���p�x�D���6�M�B�oMܬ�	�n�wM��Z�>�A�Q�T�w�D�Z-��߄FNˢ>,l�h����e��.{��P��ݼ$�x��CVQ� �eܪ������Q	T�̆v�q�Uep^����53z��q�i Db$���X���/����+(M-���2�[��GK�5ͱ
}����up7��2QX�Sp����)��-�sr��k��ܯy����:�]j��}���4�[�����j�f�p8�m���s�r6�O��#����B;PKǕ�q�a/4/�Z�d������lH{[��;�#�Xr�	D��o]S˷f��2�@v�59��M;��Tt�	:q���-Y���ɕ�Hm
���r��N�c�����8+��͵�읫3���ԉv*n�Mh�9��},��7�;�/(oK�]���sD�Z��2��&�B�|i�>�vW-�Xnށ�fno�Av�|��|+�NT�3-���f�2�xc;��}Fd�n�A�m�����,��S�;K�=G�[�y6)�"���u7�\-�*҉��0�38��$"c֣mŨ�Vv��]J�2� #A�܃p8�frF+�P"�n�%pӹ4p�����h�"�������[T�Yb�멅2"���;S�LhW�X���9�s�M�\O��}S3Xt�d�[%������t;X���U�eu��';��QS���w2������ۭ1��>�h&v��j��/�鋃��a⊨�G֬uc[
0F#���T��ĸP�eZX�C���������>>>?G__^<x���kQ�+���kB�"ә��T�DXm���+*i3�z����������>>>����<~�0��K
��Iƪ��2�7�dZ*j�q��=�ML��L�Og��||}__^<x�~�\J�������m�J�j1m�kYY�UP��IG�sS&��N���g�ɹ��vvvYe��H�<qkf[aU����&��c�(�7*]W\{z{|z}~>?q���}}}x�Y��j/(Q�8���Tkd�4m��"�o�V.�y(��}~<z~8�����㏏�����Ǐ�޸QB���m�2'/�Zn�U�.cU�B�ձf��UQ����[.Ij�_r`���>j�X*���
���ar��Ҩ� �Ɋ(�T��/����\�2]��$UR,Z9���S2���"Q���Tv��UU+U����dX����"���G�7bd���u��C�b��ò��+�ˆ�Cy
M�4�I]�^`[�6�9��5�h��N�o_ȈC�A!��� Ha��L��" �$'���������H�,�.5��vB��= ZKɨ���{c�y��n�tn8�ƾ;/L�m�*�d��az7���DǠ����>[�P$�� ����/%�Q���~���q��FxD+eW�Gxx���?k��ϙM�1)A��!�P�c��b���v����ۆ�\�&e?Z�~���>��}Щ9L���8����pdR`/s�U2��Bt�?N��fz碳�^�NJ8	��{vxd��"��ْ����P�kHJ-��h�>����ǐ�a)a$\�l5;[=�_�̷��<~������:��,�a�P�H�ga��ԭw�AW��v!W�Y.���n���h���� ņ;�𰐆��!��g#���^7��K�d���������U��o�*c]��B!}�BgΣ�;���	�a��*�G�9�j&��y���7�gk��:�� ��<�[���R�9'5mv�%}�����1@��p����^�o����L�'�����M�VG������{�E{�S��f;2�F���ϝlL=��QP�&z��x��}��u�T4����M�G|�'j����S�W�)��w�3E-��tڋK���J����}WOf,��kؼ��ѓ*b�mͽ�25��u\�O�OD��.u۹)��1r�����2��~@�������d��!�$)��LD��������""L>��`���@���|DÏJ��mO�\4ّ�1ъ�z鶨q-K21�s�Ͷ����M���H1D��� f�~n�+	^ˏ'�]{G��f ?CĤD�1�4w�#���V~��}��ţ���% >�%O8�4�.�Ң�ǒ��L�Z�����XA�q1F�E'� �7��Ÿ_
`z#��H!�T��\�!�\�l�|P?,�{����k�t����z8`���[��^���G���%3}Qb����  �6v��:��r<QkH��C���l�i��e��/m��HU.�n�::�TْJi�])Q����C��0C=��r�P� s�UЛ���m��ھ��A�����]^Q:ͯC�-�k��dLdo|BƄ�͏,�B *�V���xX�R���P%��N���A|�;shp��qY�Xq�*F�cB��0M[G�w�㙛�b}4�f>:Y~�Ϧ�֔H��ִ���\��Nv���6{ ���|	F]�*<<=3 |�9�<3Ʃ�A���*�kQQ���h �k��"��2=��G&䣰��d�T�^���V�V�,�Ux�U�fbƓb[gK)��uz�X_:���N�^	Z��J�$�S8��`��3�.|�d}y�<y,Kx�^��C���zT���򆌖�j��Ve�G��rh���W���b��mu��!!�	4JƘ��lӏ<�ה�j�)tf����$���"Ea�%82 r82�B����  V@�ߏ�����{�|�۹e9/��Bbp��x,D&9�~�B���(b�\}4�Z������:ő8��FY2�h���o�K���S%�Ϯ�
�BG=���F�p�a�J����۠&�5�5}n�`��|��kj��O8q� _ �H��F�¶��Priai�z��:��{и��Be��@������D���9�������z�3 �cQ#�ߝ{�W��D��-#k��1�c�n�_݋��?}g���ڪ�7�s�Ũ���%�[���(���e���mI�/����|�r~�)��q���K�"�9"�h��SL9��dp05��2@�Ll.��,A`禟j/�=��<3�'�����Ҹ��o�m}I0U+A��|zЬ��ؤ<{����ޮO�غ�<�����:n�� �H�ذ�t�ȍ�+�����b�� ~P��$<��_���IK����f�(�D�ф�.����z1|~��P��ُ�^�ډ����"��_�vO���U�)�䆙Q���ݓmCY�O}Ϙ��><>�]��]g9���$/��p �ʘ���py���-
<߷m�m�d���̫[6Ҡ���k���s��E��� ȣv�i�v�9����]���, �;�m�!M�b�ڑ�;w��r�޹k2WrA<���?�Q�d@�����!FI#��s��s���F��8y���xhَ�6c����p5�}�vX���8���n��1��`����Nb��z�T�0� xy�(��9�>�6�_�����q4�?�r.})�眝s�z��R�y�i�=�-.��	��q��? ��>4D	�jޒ��M����=Z˝�� <�q9��~����d�[1J=�� bD�Pʂ���.U��[?��8�0N2���[K��r'���g��}=8o�vx��|�ET�*�L6y�H��P����n=��57�vn�Ǻy�&��e
F#�u�y������~�����y�G�' �b�LJ眘��{ӹ5u~��2������&d"%4� ����xk�d�rE��V�3=�1�����������BiN��a�Aa���w�㼔^��=�`G	��l��7��30��ψ��>6=d��}#c���+߅]����_��{���[�T��a��}�fm
7hX�J6|Q���^/�-�B����ժ�\����~~�w6� �]6���>B��_0���H
!�@�oD< �~7�w�c�ԭ��.v	 k���R�a��!kM�޽����m��_w%�F��-�`qV��}���3��ț!�;�Co5��Yì7���7*0���8J�9,Ӱ���+s,��e�֕���I	} D~(� ~/���@!d
�"I&2I�<��߻����m��wB���=|"��:�k���c+>C`�9b�+��3-�!�����=���Y���<p�C�ϋ��^�����1v�x_ڢ�L����������|�Z4P�Ό{k������/�)��":%�+��AȘ��Ei��}�B�엊��;�<�q]��`gM��X<i�xe�~c7CG���|�����-���/0�st1(��Z�ζ�Af��*������}[�,�e�Ԃ�4G�2��%�MIh6g�Ʒ^Ax>D~�����Oy_TdyߘGu8�|z��g�GU)��9a�yfl8D��=J{�y���� ��L�R#U@ʇ>O�c"���*:��0꿭�׉��sz����9�y��1u�ֿ�z�q�������=��>�~u��*T�UA�|~�f�{K�^�^���;��Or6���4hr'u�#�6��;Q\�Uv�{�8�����v5�����3�������x��n�wP-��`����8j���A�צN=��B���S����Oݰ 4p���Pԍ[�$j�%�����P;�;�ݝ �{���)�߉���I�֬�����E����b�[�Y���]=}U'J��YR�+�K�}��WZu� �G5k�i���h��{f��W8��2�:��k��O�'Ԧ�$.��,ݾ���]mR�x? I����+��aFT�G�@��	�W��h�|��|�fx���V�}��#�ȕ�Q3� _����m�C�k���G�t�_�{�"��U�T�����Y��DC��f����F#�;��'���2?�:4�c75���Cr��rˁ���mI�|/jU@��WOHm>���w��!�1�FPj������~��mN}�|���/�b�1�H$�]"'Q9܈rv�[B>55��t��UZӈ5*��]�jx����������se��O�453{d��W;I��	Q���p����w	�s��^ʜ�;*�_y�xtx_N�c;k�a���3F�S�N��yP]�*�2�|5����Ǯ��ꝯs,o_#���Z�˻C҈�cgP�Ǯ��EQ�+�n $n���`L����`�H�\nEfi��8�O�_�u*�ԅ��b�!�B��Dd�����<�E���6�Xp��r��y|Z��q�������v�t�H"H3:���m�]!�|��lƗ����}��/5v�z���s�w�����:���k�S���p+��_0�@� �,��-&~T���n�l�]J��k�Wu��m������:���Ģ��������K �(��(�ʵ����^V����:P�a#tE0��Kr嫪!������2�����'-ꡜ��ø���od���wYݴ����x�Ț⿗�$^��AHA �4��v$h�DBA�`��E֮ytg�W��=a?� J�)BȰ��HaNB��H�J�t��3��l�Od�Y"Z$;3�ż���S��,�e�GP%�t���`kl<f���n|��=�����K�[W�\s�ot�u����Wl��p����w�_&`��� ��S���d@��.��׋
�9���<�X��vf����*��	8���1,�$T��U�R�oc�[�Gd`�p��B��r؞�/E�����(����ン\��3WT�#�#_5~�qü��/�����ݘ����g�jV����TZ��icp���aׁLIƐ<��Q8�n��@�l�� � U�ɏ#�A�$��d���H�։p�홯��
��2FT麽~�>�p���T���C7��q�eG�mI
���u/�b���)�C��BLs=r\�@���m�ŰGT�z�2޷wi�rD�r=�������!)�>U����Pz�~��7T��p�u�;����)6�E
~��)g��9A�!�:��
@�V~�I����%n�J��g�[�O�<W=o{���z�4q5�H���"�07쇂��ߐ���r@N$jd5�eS�Qo�X���m��Y�1��ۭt�f��(�M������b�	V����O3�I���d|���{���i�q��k���
�"��i�X��[�$����F\�{˹F�v�y�k}OI�Ӯ�U&��a��u�ң��@�6+�@�H�# 0�0��P���Rz��"I!�!��~�5��xz��A?��ę� u�?zA<К����"��>��-6�ۼ4Y='��s���}�H����&��Xw��@�ƹrQZ��^�>\�vAn�{}A}���{zQб��;��a���mK�
�or��{#��X�|z�����(B3�w���u,���,��m`����7q*���*f�-�>^��8U�G�l;��v7���v��5Q�1�}�lm�|�:w~���?0R*���ש:��z-C�<I�n��A��h<�Dz(���_���^��u�ʼ.V��~M��N��s��J�H*�!�m�S���V���6Fg)�f�}�3�kUi�K��[�ƹ�F�n(Am��=���Oގ�:֝��y�r}0�mK$��;�Q)��nNR�:�_)�EW�g�z�i�q����q�m"�>�h	����/ ��Cd���`�oU�\N�ˇ�d�J^��T
oc>�h?i^�zQ\㹇�-"��z)�|k���>��V)��'�tB�-ã�ٻi��:qEm��v~��[J�ŉ;�Y�]�3��E:aU�d(G'.v�V�����n��ɡEl�;��m��ly77xJj��m�m�]T)�3���ώ:7�xo���2 � }��9pd�J�eC����9���7��h�����O���~�1�#V^�a������-#��s��tE�]��]ѽ��C" ��"ώi���}���\^�G������嗠���d�j��`���;��P�1�y#�K����ϏWG���S����)4>c��&j��qk`�+ҍ�P.<��ڇk 9�]��a\3�V���~7�HMt��?2����T��(�V"�@��MT����2]GP��I�F����ۀ��d�=X
M�[R��C���'��p���CO9Oue*n�<y+�7���w����N�����7?0��'�ƈ�h���D;k�n<�)?8�o՝~ɹ�ξSu�� t����Bk
 �mtc_dx���4��g�ʚ�[a�J��f5���8�׷�~_?��������Qި}���\3�@�g�����ˡ�r�5e�d��!ߺ���f?�KVB����2~"��6x��V��+�@���1�����GOb�9�ޓ_a�k�C���]j��A�Ɖ���s���$W���q��<���Be���tL~��lu���Ǳ
���ʰ�tcU��eiYu}�q �]��q�=������-�=Qħ4z��h�![y}\kP�Y��7�	e]�>��t�Ὄǝ/���LLo�=�6�d6/��{z��4�g� ��� Ab9>��(N�A�!80��R�<�x{�8wRY���0�s���8�'����D��G	q�>��(|�B�/����G��Y�b�!�q�w�\)+���^�x�![�L8�
�5�vu���&nGޯ�"�
��,�U}$�;A��#	4	
Չ�}��<���7����g �[����*3��cNOK�%��{#����`:�Ts/46����Հ~2����ߐǤ0X�gyWS�l�A:�xMMF;�93�}v����??t�dD��d;Vy���$!�P�Lb�<�p�v3yXcW[���pur�.�D�eG4#$r0�a��aA����G���v�ύו�.���[�u����l�O��$��JX�&tb�0J�!�`T`2	�8�l�V{r�Uߵ?�n�Ƙ��U�wO�8G�`�кk|�W�H�$��>��\h�4{ѐ��*�q_'�uSn{��=��[{zD1�O��hw��d��޹mO*%&�-��WE�-�����1��B��/&���`Oʍ�b����ǽ8buu�Wv弿 ��<�湧w���:?`��UOf��\��{,T�;��0�U�2��M���̵\���%r�h�b�b[�/�t��e�V���ӥ�G+�����h�,U��2I-�3t�� h���rj[Z3睔�0����];�.oQr�+M{�a�s�������Y�G7\�\wf��h����t��@�X��gw�������7q��iw��OrU>gv�9h�%������3Y�|��93�5D��A�5�z���ʘd��⣡8U�*�
u%ޖg]U�j]�SP��S��4Ō�\@ǘ���ŕ�����T��;E�n5��3S�&:8�!�йL�����FJ���t�W>�;m��tb��9S��[�7�k�۫��M����#��>�.��CzhiW�Zv��U�o���ϲ�g:Z�0��)%��*�]%�X는�z�6\�㉇��s��2�+Ulu�v���y��x�3��y��m`dM�/9I�v:�̭�tA8������x�P�U�D��a��(�SM��Cd[{kG,2m�,Υ�,YW8�aY3b[�vS]3k�S��m��bf�Wb��b3V�n�is��f��5J�
4(E**�fq��*��y�d�W��ʹE��i]NK�
k^��L�v���f�����ku�G"�]^)+���h�*�x#P1�����g)��	��_c�Қ�S�Yy�z��H�T�f�50sbwUd�S6�x�Ve���yUg{a�-s�MD�N��u*R9O[�an�v�sa��E���8�2�V<8���E4�="oU��T�KG���e�U��.��^JUR���@w��r�}w�")Gmv�R��X�W�{�˩�o��4TI�Ә�y�۹�]�I��l��&⾣Α���p�Cn�t�]/���0�9�"1����GNp�8̼�n��淳6��˂�	z4٪%ux�o�gk2E��Kw�u*k���3��o�E)ca���ڔY�b��m^IG3�Ǫٷͧ��A�)K'�b���#}�����e���NT��B�}��"`���e�\4�yp�[݂Je�oE
D�}]��絖�z���S�5p���F_m�h>�L�6&M��������c],�"�3���U�ewq��9\��i���o�\v(+zp����z�8��N�X/��m�6�R��8�O*]J�f��c�}�4�^�h��U�#ޚ�0uu�&�6�v3WƷ���i�Pھ�}�]�����d:�Xuj�m��i[�����윺�k�JOǵv�W�s>�)�~qc���Of;���{ב�Uä�9�-�Jdm�B�I�iuyL� J�Y�E��J��[UV)�*�2Y����r�.\�N�&Z�ݠ�0Y�N����y���$[BIJ�D�I��E3%!u(Ei2��l��t	�R	$�L5��L��t��eT��T4.OD�̖Ȅ\(��Jån���T04�Q�D�)�S2����e͛���.j�N��y}<Q���,�j�ʛ��Y[j#�S퇆U��5ʉEmw��c?��fM�̞?_�8���__^<x��FAǩ�yO0���*�X�"%�����AiYU+��a��Ǣc"�"��s���ge��}lUNj�j����֋"�mDb	�q��ތ���7��Ƿ��o���8�����챜:�h�*1E+F��2���KiV�XS��j�db��Q1�vnY���٩ٹ��y<������3�����(�5�+2��+��E��#+Q�E-�kmZ)S�ٓ&�gǷ���8����ϯ�ҹ�1S,U�-���-*(�R���j�U\��37;fM���N���g�ɹ�;;�g��T�*ew�1�yh�1��n�5��Q.��R"��U�����J��$��A���o�{tb�uj���W!��@Bͥ���(��DKiE[�dY�U��B�._��˼��R�J�E�Q�Aq�(�ib�U����E媢bPCV�j�ii�x�.�����B�2I��h�#��;+���s�5��E��C��r���w���l9j흠���C��\�t�E��'�IJ�5DJ$�d�BSa!,n����� ~"$Hd)�H�%aH�2+!�͢����VT���'��/�J�F�Kv���ly#i��nw�v��coe�<���r�lx���L�\���_FC��{���z���Qe�p��D��H��=<����ʬ�v����Ӽ7�؜�mѾ�aր��CГ QW_K�%�c&��S��=�i=M��X\kq#�0�a�y����\�a�����5͍1�͕{���!�2����/����i����7�����L{�Ϭ'��(���Ɣ<�M��P��|�fD���Ij����C��5�B�l�`5������Z{�mV����y�^oƄ�:9�p�}C[aD��Л*�}�VG���Ji�N+��ڋ̎��l7P~�p�#��	����y�@����*������klЛ����K����Q~�����=jb�R@ʢX"��3��������f�D�:�W����$tRz�Lg��y�&��L�u��]l^���-�'<�7 W��W��>cVy,��>�������q��|�=�#{n�K�pD�R_Ոf���Z�@��jo����;� �+s��{V,��t�2���
����obc�@��z�kHz�ʅ���qQŷN�����Wv���;����S�a�"��ܞ2?D A�$~@�#(C#�x2$1�H� q���Gq.����>�uO�H֍�P� ���pߝc]K奥�ʽL�ܵ	�x���wصt����s��(��A����B�?%����Ǥ��OE�f�sy1"�7M��s��Dp���叾S
HNE:8yP�����H��ޔA�c�b"�k2{�?:L�X$l��;�m�]!�(��/�R+����t*�_}TӪ�gG�kh��T�;�H+мО�_�%�	�^�?�mb�gf�V��Hk����6g̶|��ÞK��" WNb���4j������4�Ҡ����0��^��ز9������Ta$�I���~�aˣхO``�n6�S{���x��sޫ�Z��h�cF<�;��;�ٳʯl4t�����7�	��V�&><_�o9w� ���0=r6��"Μ��t0V�r��#)q���?�����Pԧ�Hَ�%����؇r��5D��M3Z+.�{Fp���O�Z��.�$���S�0��1B䠟����1[q�������r,F�]kc�a�L��a؋NȂ�=����X�ˬ*��ĝ\�	qj���'�H;��NkJ�U�H�@Oŷ��S}^{�{<le���T��[s}�g3�r��N���M��.Ǣo
��7� �V�*��e����W��FP��;!82D� ��bB������������>sп_�J`�kAa 0����/�ߩܻ��wf*�e��zD�8�-dc���ϡ��۬s�Ô��boCۏ�n��`�a�'-]�{h�<��&!���y��/�g�.�.2�ȶ�S��ޘ�?A��X~?�p1͓|��hc�g�M3�lv���/�~�w�F���	�螬'��+�����D�4��j�r�g3����B���\�ϿQuҟ0�2�H�|zb�����au�/��tm��8��!WK����O�%���dx��&�,�?L�p՜�vX��Aɳ��ы��dp�0(��=�ʦ-�ÏU�l�ɭ����w��S'�Ut�5�(�pƯ:����!w�.���9�Io,��(7{��~�}Ig�� �~�����؏�@���̻zj)�*�/^�9��n��fi�l�>ŧ�#���O=>1즚�4rA�vn��P*'�E�}�r5�{���1WbV�cܓ�,7��H����uH�K�1�͙�[n�7FE��a�2�Y�dslB1u������f_Hg�8�6�V��U�c����2�����U@��uC�C��\�����}��oq�C9a+^�/&wu�8�6�g�n *�
8�H���AVmt�r�-W���m��}�}�����1��@2D��	J��s���{�Ϲ�����6��#P�o!x��1��ŗ����S�N��ۡG�T�vw:�8vMZ�{�Z���Ag} Y��塠�&C�ϱ[Z��K�zn�Ġ/7[`�p۪b*&�k.�cN��M����}{��0�f��;3D��p�=��f�� ������o<m�2��op���X�1���
��(������p�
a�!�#~]�"��ZR��v�[�,;�[�x�NBa��Ǫ�1�;:j9jM�������XU��n*n
L�kq"{��������+�#���U�}��c����k!��կ��nEwL'����*-��1�%}�k����P�{��;�鑇�x�XC�&kfU4î8=r�5u�M�p�7L!aa p�H���ʢn�=~B�����@Q4KF\�_>�5��@�1F�k��#'ܾ�KH��<>��N�$$R�(w�`�Y���}���}��t�ʒg�k��Ac�o��Ȓ�Z��T`���AP ��SՕ�=�7���ը�m�x�d��k&�iUC�-����leqX)���Ƿ��CsB���q�b�雽G7<{M)��b�'3����򘒷��yO�ӛY
i�':��Ы1�T�.�y�ow)���Hg��-$�M܂���$�52P%�l���m��{����a��z���  �����K�v���.�#m�Y�d}|��K��G����Ί򭖱P�Yu���_|�� �\�O9<xp��.*���-{Ҍn���5�4 IK��=�/����Dg 	���)}��g�4�+���eF�<��S�M�V4����˄ێy1�x©���)��ڶ��3��02d�(d8��5�KP��1윐��4l�$��H~?}}խ��N2�* 3J�]��S�p����\. ʘuJ���W O����\K�LD�N�L��>��~������j�ƾﲳЅǼ��7�7�I� o�FPp9�S�hW"y@���u-A�ƽI�o8������6�74ʖN7P�N+�/:*��_�kB�	�G�|�1�R"�	��^��pޡ�RzOC�-5��l���=�f��r0gx����:M߳_�'ŉĪ}}?R"V<n0�r�����"�Kzm);Ӆ�˓à���3ь'�=" �-��Jw�]q�T��.¹��'�Ǡ;�Z�2�7Ӱh��6hdnL��W�л�x�@�#,�DA]qW�|��ߠM�/v��\�`#�m%��sꜯ)��f�H�ic���J9�C���0U��w�^}���6���k�T�m<ҹ��b
L�9>���zBz���8jc��Z��3l�ؿ$!�	���NJpYXJF	���`ha�������G�>_A�d&�a����*|�5(qa�l�{�cƃ���k�Z��i��D�cf�Ά��.D��W�*��:N������[��.�E����+��ڐ�Y
�Kwfsif�O;uF���E�_�����V7C%�Ώ��Mg�s��畵�vuƽ*C�?U��t47.-�5�C���r}�,���3P�/�b0a*��"߮uD)�{�&'�c����I�>D�ҷ1E�{A��KP~8���nx��R�U뤀�U�����~������.�9���y��rbtКvwq��T�֩�rY��OF��ӊ���*k�Mx����q��+��&	�(����+\Y��T�{���D�����L��,��I�)��9��:��ë�r%�X�-�<�����lQb�4�Bw�=���}�j.���2�|���'ѳ�����^ � 굾�7�.�*s�ja�
4��z��;�l�J� ��`?N��g�˭Q�>]7n}��J�]�ўq�b��f{�|�y�\0�s>��]T���;�nVnp㽖Z��̋��2��=��`I�(#��x�A³�RU�K�w1`U�PT�ݖ�5[O��L��@B�{79얈8�����[$� �>�e7����U�e0�N����=E"�"@�?PC˃!0��P }�����1�����^Ǡh�6��U�/���hZ�}}6��P��N�vm�]�za��U��v�>_v�޺=�$
9*��)�<f>]:��pO�)=sǷoˬ&�ڑ���[u��o������
��^��jΔ�8O����}�D��k�1��\���<UK�K{D��IM����p��#Ѭ0������Esp}"|�/���*������-�Z��=���{�C�	�{['裦g��d8��9C^$XJ�(�/=K�~��֚�"�i��θk�ΤO��ù��=�T�:�f����f��L���	�M;�rR�@�lm�<+���9���Y���p��*�I�$�?����Q2��Ed��]}|� YZ�L;�2DaskXO�{�;�FւK�э��}0�a��P��V#Q2S�wEp!�e����A��?�~���։�<�j,�[o):�28�>��\O4�ސ��ۗƣ�u==z[������>�!}��
S_B�-w�1V���?	�x}|.H�DUZA��W��1�ؕj���r[��u?ޱ�5��_�T��ӂU�^YI]��o2�Q͋Y&�6�B������=�os�x�)<��!ħ1���r�o^�2BM�݂��ٷV�����2���B�@�'u����^n���g�'�� V-#%OS�%%%�"	�9~���M~���/�~���6����"�J�"C������hmO�����O����?�}���?|�z��:���lW*0�ZQ�|��n��*WQ�oq�y��-��(�p˗*���ù�yѳ�F��R4e4G���b�V
?��#�ϧ���6r�l��(��>�~/ظ���cx>�u���}I|@5�D���>LI����9����7|��_nK��vl�\��4���A�Eo�������A]�E�d@�Nl��}FiS5?�+�.���ƪ�{��Uݗ�[��E�͆~�/)��B�p��ػă�!���v)�����v��}9����q^:�w����ve��[Ӌ��)Y0Ŀ�'��&��_wH\��#UK�vvSoG��B���v�}s��2;�c��k�+�4�zO/>�t�.}bdkjO�s������E�۲����=WR"�a��Z��*�+������Q\�Y�6D��m,7 ������z���=Q�2�t���/���}�~Th^�vu�`��I[E8+���gv\�"�?��{_o��(ۯ"�=�f:S,+
�}+�
���u�r��u�]B�Y�I�UJ/4	��P@���L���ȴ��;nG@�Χb�6�Rf;�^ �r���K�1��4��V6�v6:�A��o���D$ڢ|�Kɤ�QH2�ti��)

� �A:�^m����$H��B"F��h�s�q���<B$�����¥��J�R寏�Í��]7Y��PƐ�^���{�et,�w]5���9��g)�3#揁�ȎA�o���C��M�MCPn2-�%�I�����,�k6Qcm�w:���$V&��BxE~�G���?;��;�S[��K#Rjt�)"�˦�燹�'�d���'��)ħ��bcd��1b��K��\�c���Ǯo����ջ��~�� ����!!���Eb֕�X���$@W�(�ޯICub���w��6����b�B.�"~\�<�R;��#@$�hNN�^�]}+�ʯ����� a���Lè�'dV`��D����`S�M ��b�xG�gg5�[�7�&~K���Ӓ!��1�HW#�"B�%��N>��lǧ��m�3%�hd2�7Uy��@�%82��Cc|7�^�Mq'yb�<�P����kϕ�:���˂����:fw��%�0l�Z��^X�J谥ѐ�E[Fs�
�H��������$i���7&~��`�Q��x�j��z����U���0�Rag�^mHA������#β��R�G��u���cGێ;��@�M��.���r�^ͼ���t�:\KUt'���Č\�{�Kjw�j�H�=��4�"$R'�0�U2�����w���}�K������΍=�k&�8�מ���)�yF�����6.H�H�G��|�=x���	d�s�lT8�����>�s���+k�b�h&]4{�����wC��{d����7^�f�>O�/�7�_t���P�X�x(���E���]�}x[ۆVW-3Pb�j�;Y�A�[6�zn���
��UN��>�O,9�;~���y�a;��էw�P~`0l��a��+%H����$�֙r�,�;Y�f�z9��5��\h�jH�f^�l��u"�G���� q��8hj ��gX��B�_����TSrzǮy��Z��Г��~iq���ٻ\��e�&H�H�{W}lz���[��g�M�ì�~L�)�8����Nz�Rf����,��|�1���f1pSzF��7&�:&1��'�"��O���}�~��0����{f^|��Ψ�8<��\@�S�5� ��;�U\�m�\l����1�}�U�}y�[%o�0C��33��%
�ѯ׃���y��;�rH@�s�y���S�-[a��Jwg�c�X4�HJh�/��]��g����D�:;��)����,��ܥ�onWgU+JW�F����15�2�,�T����o�;,��ۍ���e���1vg-����p��n�c�D�/�=���qםrVd��q�It���K�R'IΗ��4�,��.i�x�Jz���=f�]�s��j�ͺ�������O�e�&����)�キ�eX��M�[2*��|�5���b�G�
�5z��S�%�F�Y|�v�\B�9�[|y��^�=it(7zsCNĨjI�����xi�`]4w�Kb9�]���_{���Fج����b�6���Whn ��\l+�ՠZ�F���Z��3�Yٗ-S��Vl<�	L<T)���_[�t)�a����C�4Q����1s~�bذ&T�#�w��W���G�Q��%I��]���r*�u�+��s��#�b�t�Pa�6���ɓdWv�5.7�]��3b��d�N����WwI�j QN��Ů"\���ڃ���25zm�#w<؋�
M�W,ȁɈ���S��ޡe��f��0��c���٘�R�\�Q~��8,h;�z"�,��i�`�ùW�d,~���燱[Jоt��l���:�[wV��$�T>��>��cd+#�a��J�om��^]��>v.���������Ñ:J��3�U�&�R�9̾'kw3��4)H��i	-4PM2NNN�s���A^���>����d�PڿV@���z��u�n�a��;��ݼ*}�����涫y�247�A����e}��8{���N޾�l�QS6Ԏ�m�ӕ;���E���Yڧz�)ʋ^L��	�yud7�Z�\����h���ȄVJVz�U�%,��8�5�o-d�M�m���O7�����h�a��̪҂i�Ȧ{.�uX,c�ѥ��PfLn1�嗝L��]�7j5�Ť!�S�s1@�H͸񫭜)u�]�M��]:�zss�WO��ܷ��T����nj��-YU��*�����]s<s���w&�~����j�٬_�R����I��nɺp�(,�f�ʊJ���s�}�(cI5*���Ե��Ҝw^Kܓ��nJ����Ԑ�n�Q�N�2�_p�W��<Δfk�EB��0V �}��"��L����=b}֩��gs���J��m�7�WF2����q��:�7u�_�pR���Í�L�n�!��j�5�)���F@��� /�_r�1u��'���݅I��2똽qDZ�I���XT�l�o[U�HE��t�7,[��^K`Y��e�\�NV�Z\�7��h:4��:�-L��ĂC��J]f��*�X�:�
"�((�Ȫ��ϧ��57>�������'�s�vv3���}�O��*�`�nZ`�(-)*�Qb��Դ�QPt�)n�8ª���Y�N8��||~8�����ϯ�+��oa�^Z���+����DT<��M"�l���m�k���_��
3���z{~��||~8����>�~��.���f6�TV��R�-R�Fɫ�J�R�cge.����ޞ�}|||~8㏣��3���EEQ�������\h��LL��W*P�Z��.��-mh���M���nn}9=�����q�G_Y�]>^���TEE{q#t*����Y���-����!�ZP��T8q1Q�訨��ȸ�����gg�Ԩ�3���Kh��fB�DSį֊���YX1뼔����k���:v��ED,�n���yj(�2��QRe��aQUƪ�n��<����"�+�.QQ*+��#̦����X��8VƵTEM�ō����k���U�uB��f�j�FbUQ[�f5uKƓ�+���yu��	}ljlWHr�{��:P��I��q��9�ArH�MR��"$kH�R0��{�w�s>����y���U�6�y\ӊ�$g�q�g�(QL�Й�.���s��0��jM�t$Y��5}_!R"{��Ǣ[ϖ��9���y"��v��H�zg��g�x�:�;+��E;v��ꑬ�+�:oQ�TY#3�o�Y�Fr 5G�NA����L1������M���Uϻ��]�yh��:��δ���׾��Y��U,���d�]����>��y53:����ޝfe����	�	�i�S�0�J+�%��z���+R+���@
\3�mcV�i��\��-�_�k�,;����[o�s��p5��uko��	ܴs��%8��sXά�\��hF�L'��ok+�����jd���aG���<X�.�\z�F�8�Q�w=�s�	5͡0�r�ҧ�]�K7(p�ـ�D<6541`f�Azd5��d�����rޗޡ&�n*�9sY����kn��`��:�O�<䁕��,�4��2����}�E9m�I�`K�iSw�t,��}�%��\gЫ�~�"�ޞ3~f�N�v���,�G��X~bZ1��Kջ�Yc?W�x|}��o��j뀺�Mh%�2�7�s�9�7�d"��vE�Zٷ�x�ܸH�i]�$��F6L�޻y̭��&��df�6�q��0G�S�c��+�)�Ք,���.��ս���u����	D% R^e���,��w��}��3R)��̌ف�;��C,�i�>fIN�N��� �v\c����3�q*���;���3n�.��8��`�#���>��Vd!��]"t�}��&<|$m�99��{��p�I�I���LLe������ ���/%�gc7������]\pv����]�I7B5&�L��/FC�S��m����$7��b�V�fmO �jմΦȾżF��m��k�^d�)ߵ�ع*���?�������/��C8��t�����ϻ����+W���`����>ITwOa�r��t���f����tZL�Y9y�oh��za� [���	�Or������l�PV݇�����}jvee���_�8�3�K���.�-L�^9N��B���n˰G���
f��V���ǚHW�����z"=ޱ�Y4�"�q|�=JD����Ɉ�y�Z���D�H�Y�����$+a"5�|rm��B}�ب��^l��?{G|��Ǻ��FÕ��U�T��Lw7���<����!U˄5�����|f���ys��Y����MW��1XF��.��'V�g�$��H~ fB�\0ۧ����������*U8e�EC,�j��q����EӚ/���]����<ԧ+�5M%a�Rh6P��R�&I%���H��H�Ӗ�uT2����D&`1�������bJ��H�C��������o�ߺ��Yi�L��J2�(%���y����}�6����Y��E0M/�s�b��\�ݱ���;��`���e��X׻��ך�WHv�Ggf���;�VRce��H_t���<�<���h��=�⌟51��t�
'ѹ�鶙���1o燈�y4� eY�3�w�#=W�3Sﴙӡ�c{�8�}l'�:^ܟqP(_��*�u��L>��#u#q+[8�d-g����x	�K�M�L�8q���1�ᡸ��o_t
ˍ�����#���co,I2�B�Z�:.T0LA�B�/�����XkM��>9�ac�V���~x���/��uAU�X=S����#�@�t0��)�H������a.bا���˭��w��9���Sg�đ��~�2���
��;/WXn9��L?��!�����wGH��ѕ��4�����ӲİT�2� >�sCs뷻*�"��(;L�l6K0{�ѻ��0�=��Q3���l��x�=��o*��_q;{��u
�}��Z�I[��WT�yU�`�;��W����q�v9���6����[�[Vd����ږ��ef��4EG3f�kv�*��kJ:�PE%6��e]%�k��nwD1J�m�7-�tI���蓮7��-R�Q��#���<�3	�)����9uwC�&{�F-����e[��>�QF�SW�Dۭ��ھwu2��@�O��q/���^��b���ۂ����H5�gofz����2��w�
��z������_.����g;Z�ʖ�	��B���̺���?*f�5!�}����ciu{{�1�`"�� ���nk��g?��S��){��T�u��s�n���$���\*�۽�Q1��e3ܰ�O��w��R����v}�G�� �v�0gw�a^�9NC�}��;^4�y=��*
OI�º��|�W�kCuن-wXR���Y �#���W�;���**5�ݘs�|j@��s9t����O�q	TaJp�
KT��+�6_�{4�wuN�G��M���W_U=ݡƞ�^���N�;m�
����f"#\X�'���s[`�����_��=���M\ѧG��n�� `�J�n\X�]��w�N��2��7�T���]�c�O�r�L@�j	�ID�@����@���i��tS
�r�i'�=��z<�]��WT��	�O'vl"�����rk�&���U:��fvv����q�����w,U��M�^)M7��^^�=�,�0���V�]WK��}%~3zx,�ˌY��^?��Z�����1<�J<�;�0�lǁU�����;Ŕ#��gU��vu�y���
{�KӤ�v��2�+xv3�h��c�_'��~]�6j��M~�Y7#�8��3N�U�����*74�	6���(7�u=���2Փ�Bn����o���ę��}�=Y&���No�Ն<a{���z!�+�Q)���2�+��gk�^U�|6]]�M$T\K��t��	T�n0(l�s�)���]^��̧����2\��f�o=�;�l"i΄f��%�s����A�����l��0v�v��+��]f��W\{h�{��h���g]�[���5P���ƹT�?���T�%��q�]l���V��!��k�;cj ۛ;�	|���Kf�Y�ꒆS��6�oEY�>a�����P����d�}WG�$(v�j1DD.|�UC���&��9����f
��~���}{GFꗍ��oc;�u�U��:��)<�ܸ�;���l��:����g�I�F$LKi��k��k�B��}�W� *�s�>���N�GǱ�4�V]:u��=�Z�i���Ἧȥ����/̙k~|�>����}�*h���W���E��zs�s�=�.�BRR
jQs)�HV�;67Q��>l�Ͷj��)8��lH�Q��땀��W��i7��r1�P'pϙ�G���A�ke���{�����KpQ�Qئ����sc֬
���*�{��
�Jwj�%��zI�ӍP����/r�)���|Y��ϘＲ��d�3�,D�T�P���W�3���(�qM`m!�Zj,Gg��S�����T�W��l_�/�^�g`�m�u��S�~���c���#�,m�qV0����a�@��+�D�f/FT소�]�ā	�i�g��L��L�r<�	��
�@�̇./�Ugx����|�~����}�r�L�N�Ou1y=�w4��۫}�s
웲�n�S�]WD��]F"��3���FrKΦ�glR��V�F"6*c�<�;�3.�\��
��)�P�e�|s�I͗�=�m�D��Y � ��&d�%��i:-$�&-!R�y��?�H���%II�o���u[т嘳3�A��\�UQ���3��6.@�"�R�<-��s��ٲ�g��e鎈��mt���@*��"�{Q�IRK��]�b�/�L�b�"���A.׻�޻���;r���R�Ǔ�p���M�t`���)]�������Y�m�#FN�#�i:�����;O�k���=��>Į��S��;Z�Аs\��/׷�Hby��%�`­�qݞԉJ�c&�nH�=�f��i�X�rZ�������g�{7�����I�-w�*��ϵ;�R��sFN�F�.D3�.+�_n{`_Dgi����[�t��hNlD�Ta��#�s��o\��J� ׃����c�-�����~-�Y��=B�-O�kC�صSK:���kg��e�>�,ᡒ�/��~�1��m��*k����/	�6�RYއ�&Z�Hs�1㑃[c)�O+�jo��R����c?��I �~U��	�;h�j*��\�G�{��FSӦ#��eg}��	"nk����V�4�jس9o%�u�0�}Y�d�om��[�?�HB"	��$"�� ��uf����a�.L�����ȳ��5�G�]�n�j�=�x��2�vWEC8niy!S<���e�5e���ǡe~繮���f�j��0�5�>�#}=w�ْ�`��7i���34�O�=M�
���;u�Z'Wt_��������Q�!��^ES5�L�R�֩�m9Q��y�57z/�*��Hwwg5�D{��a���OXx������w'�5��{��ײX�2��d3���57���zt\�ٮm�`�5���D�\��m~��10(nT�E� U�����ɟ��q��Ο=�5޿?+�\�u���BY�z��Q8�\r��1��=w�R�u�{a>��l�7��Γ{_3���wa2z�iBނ
^��9=�Kv����q���P�s����[j�3w�c�����0Ɓ׋�}����q|�~�~�YJQ}9��]�[B\�Q�N�JOs��%pl�p>puer�c7ycݷoc@�syt�۽Z����$�\��ge�}G:R��Y���8�r`%�`4�To*�crB.�+3��[�G\�]*���@�A�B5!!$ �Gno��:_}W:>�oC�`�oc҂y�y�c+�1���.�*mEv�nZ�����S?����-��������m4d6&g{��3�[�؊���:���.*��wy5{f��Mk�Nsa��9R�+N��C5OE�~��\	�8��mv<�T��o"w;���+XK3(Y(�;��ϣ�b@(��AbPi$d�).�,���[l8�}�:sbG*������x�a�ͺ8<��ņ�ף�v����h׻T� ��m�dgy�A�{���P�իU�!ٻ�k��lZW~�Sy�}P�P��P�Q���`h�oj�NCB��K�p.����N�G�ӊ��]�C*�U�k�5fu��;�����3r��F�<d51<��O��w�]o-�z�j*&Nƭ<ͽ�Du���~��c�CZ�xx���E�A���警̻�7�H��:v��7��IY��>}��V�Mgu����BR$vl�^�r���CΖ����m��(�b��'������9in�W�EH�a��t�K��e�utU��$�U];�|9��VRWǐr/��!�3��31惜u.HE�J���~��X�x��C�?S�7L�̬5P*-z΅�sR5�\[<���.<G�m�,qIX���u]�7��_K(�:L�S͉���{G(�(P??�߼���|����W����7�k�̧+�4q��z���fu-���,:��Bcӽ�Z�^*�3Wl�~�G�A9�֗Q
�Q���Mh��~ɍ�5O_�Q/�����[Ғ�V�[n��R���=��Ke{��� ���PY������-<8����z7��*]��f�Dj�Usņ��g�"ToQ?xc����)�U�{�/m苍�BUw���9�N�)���\nW��'i*��&�i�oc@`�CE��9q�'���˳�쎬��V_�b[~	Q����7UCԚ+֦�{�
ݭ4��Lgʲ2�#ّ�=J7ӺV�^����jd�qJ/�!u+�&���A�5A�}*@�7��G/GzЖ�c"�wo�k�N��:{Y���8h,� ټu�����i� �U=�2ܳ�N'֑Or�+�Z9��Ȏ���t;?͓Oshoa��[H�=�z��C�*R�"�뭙f�hq�[/����	L+�ڸ��x�({�Y��'����\)�	�޶���%�o9rv�nk��65I�JY�j�Ô��U��ۻ���=gX��C�{Z֪ǅlN��35j�5X�5��w�jwd+W;�r��Ј�*��Io�#[|�Խ,�@m�vB��í7k3a����<ہ+_��b�����\��F����U�A�kB+�R�#��)M�F=�l���S����FmvEB�:�q�ݹ%����Y��ة�C�0ͽ#j�����.gt]��X\im��A#�����N�����Ml�33{"H��w��/��$c�L�N����a�|���,ǂ���s�w��k��˔����(���q�K�v�I�Xu�|%��Ok��b�2�l�tѫxup�4�lS'-3l'��%𷙘2W+^�=�Z�ͮ���*Uh��"	��#�ڤ��rǭ_T�K��L��z��NϿ�b(ۍ��Ej���#�j�
� )�v��G��:��V��>C�R��3_k�`�A�,VUk�G�0XQ !I�M!owel���8��M�K�an�vj��9�{;�^	�㚁w��`���-XP512к$�tr�/*���j�)��ʲ���ע�c�S�W|
03J_rr��[���X��ԩD�;��>�,�t�š�iw��4��eZ�ӓU����T��o�o�x�c�Et���*�Θz�O$��U�pjpYR�W��ufKV[,�N\��={Ю��ؙT�����!˝�d�E�[:�B_>�+�}�ud!^�̅+f�����k���f]�Ny2�p���v�
�h�S������ջ����-hGA����PI��N�	�7yu�lޚ��h��f�U7jѿ1Xw�צ: Ʋ	)7B0��j�����-f����xE����x�Wڳ��ĨE����C�%)Z���J���yZԺ�k�#!������u$��\k�"��pΔ�Q/d�����J]�W&Q9�Tz��/"5ɕ�nQ��f��n�<�o�iJ�w�{Օ�w�f��YcOeXulK��E��I냔�����53ц��o:��M��_Q�^M�Q<�&v�K�:6b�{4b�"�����^M�2�+�蕓*�a�$2�ʶ˱��Mb��J�:�q�tc�E,w2��non���f��]���ܥ����Q��'J�,�r� �P�:�YB*��`U�D'��]U�2���*e��n����U� -T�"P-132�Ze0̠�r�lMSn�TB0�	�mUH�i?&ä���-UEtT��U .��8�J� ėD��	�-D��9A�jh�UL:HSi�M�1��%�iJ��6C)_uԊ:�I ��9�s2��{�A<���X*n�k����T_"i��3��n�Qj
�Z9��\zz{~?]||||~8����3��<�]ڊ
:��l7�ER�U3W"(�4�Ko��7�0���p箽=>>?������~���Ϯ��C�hc�Uc�Z�GmV "�����a�����dD׮�z||~������q�G��g��W��YV3��J���^Ю0]%J�+TF&Z������~eQS#
�]Zcgg�̞Og�SSSSɹ�����gf�'b/Z*KN�ɭd�&�EPQfZ( �-�t����+�����=������}gc�ީ��3'ւ���Pթm�]�8W�F<�"����Ɏ8�{{{{q���:�����^�.GTZ�.S��.4PQm��X��ѩP�*�QR��Uu[㊊�(1ެȰ��b#1�.fb�əE�Z�Z��@J*
��TAb�J5kcZ,[o�qDQD���B�.�Q<hm��
ʕ1���"�0j�[Ym��AS�ĭq�ZX�UF?���5�Ѫf��%�k����ok�3���	up������ٴ��J�Z�zI��x�5REm��Gk,֔�.��Y-%9e�jS.T�șRCP�NJ���"0�W �[v�:�(�I$��	�� h���+F{�w����	�@�
��o�\^S�ܘy{�[��?z����	'�'Te�c���;;"�͋�V6�	�;�#j�T(`���V>��&�<�6�}���L%��I����0��z�>Ez9�O�MrX=��K��>�Z��i�l/>�t�ܶ����i�M����aHG������퓓�}�V�C3wrƄ�KtQ��Os[9$�U�o���$V����Br�.>���$�8(M�"�V�%y�M�{VLV��g�7W�0N�exGXGzd�h�I{q/j[�l)߶Fy���Rm��1�Mܱ��d��:�nt��̽�=���[L(Kn�ov�܇�1*e�Ǥ�p�x�A��L{��y)]ē�k���]s6�ZJj6S��۲����dց7��v�{�-هC���s�=�>��a������~Rv=�b�w��f� 6�,Ӥ|%��k�:��Ao�3o>�l��|q���v�~�]�W���
^C�l��=���7�B��u��͠���x#{�]�F��F���,!�hx���ĉ��i�"8x�x�#֏]��m���$���c������ެ��j�f<&��j50��7����;\�gi���.�ѽ���J&1���������_L۠T9�
}&mύ_vH:�����#��k��F��ے��(Z#�ڙr���{J��:�v�^D8�7t��7�;�u�Ti�2�[HN�0q�H��D�0��[F�dٛ$�|������ڢ1��x��\	ޗ��E��57��8ޛ5�jv�wf�v�"��;��h�G�Bט`p��gB�Xs@u�i�f��s�i��{��oz&J�XXX���+�(t�y����e���,�݃��@�<d2�>��F�	��VF���ʆuq���#�� �x�+{�;�ﲾ���--�JȥV6M��HRϫ�5��ث_}3>Ԭ�T���{Q�&�����"Cp�굘2���em���+vF:��{�b��\��uv#�a��cU�W*0*�^vMr"A�^8r�A��vֽ�˳{G��%��I�.Nc���n��β��Bٯ�o�|���o�o�x���j�̓Gb�5�
0���l�і������('^�v5��3�D�{t=��V�=���^��oe�K-ʝ�Y�X3��"�����gp�]�:����_f�.z�o;�z��
��ݙ����Y��FvV���l&;x�l�z����j�
����#M�R���0xf��Bȣ>k�^���r���y�Xv=�
�LF�XW�%�T���zv�{��x�2���o�VDV_iܞۭa�����<��S��?��z�7�Ԅ\�L�fkt����t��,Ö��a�Sܐ%�.)ݓ��x�I�~}�e��(o�f�5�`1�"�fm=��{:O<3��Q3��.��Օ�d�і�c 3��!f�˼�s�&�&��W���L��7��b���@b/��}��(�9v�mF+'���Ğ��\�?!-#�k���9�?G���=�q>�f\:�9�����E�o&�.� �b�1M27{�����sm.�:�չ,_ou��i��'X�ͱ���G��x���t����>���˵w�Nx�5_���� ���1�{F�q"���[g�V.�\v�35�GFh��7���sm������lSܨl�{�{~=�7]p|��AQ�.��;i�������`+�|��w.���ں��U�s5G
�k��Rr��0���>�`���s�
�����]z`��z^V��<'$Kɵ����P�x��v�`wj'Od��Ɖ��X���%OLh���NK�ｧ���#��.P���	�U�˺��dw[	m�~�5���ƾ6Y�횧[����-�z�ۚy�0�c.�MM`��b!��I|���q=���V���Z';��a<���b8��oL�O+l7T�0$�ʃ}�\�:��o*���ߴDgJӏ닛5��M�J1=��w{�H�M�iy_s����[�����_��Z����td�
�of�o@;���̫W\���=f���Z-�Րٹ{H�f=��-ul3|$�.U�d�(1(�.�T�Y`�Bĺ�uui�N����OUՇ�Y�{��\����.�V��yc�%����ܤ�����@���T���$)��Ե(��ӦvK���(�6��+r��uѭ�fU�:�릿��4%��@5�g�g�W�~1�8=]����P�g�Ng���,��[ ���W��Wy���C�j���+TױoU� s*S�q	�+�lv<�a���G^�ٻ�R�!z��0�Z�Tt���j��u��P�{wm��9���i�U*x��q�n��ء�Q�D�H�ѫ3�K�eu�5�c�M�Þ[���IUm���І���^�c�53E0�=B��Q�b�g��e��i�}�D�ǵ��dz��e�/�������$SV���%�<m��ɬ�܍w׈�U��Vk��Y��]����UE=�S:3YHD�]/�M��6ö�ck�x���Y��NcB�C߃�wk��m���Z$Ca�@���l�i�o�3'9^ �|����<�3P�*�J�Q[8�$[מ4l5݇L����"�֪7�˙![0�Oj�ć��PA���G'q=��r���E�!ǹa�SQ(��۬�h���쥰��$^�ά�q�d2ţ�jRC�� ���'U�)H����[�5�3\�7�+:����O���<z�r�"��Q�B�� E~R�B	H�D(P`���߼$T�G�]�@���lH��7�C���c���C3��c��q5^ &��z�BW������iwc }j7law'��j�R�z����Yro��VgL����rc=J:��W^J[�ɣs A�p�"��K5�d�Wvl��-�B�Aj�+�i�g��wG%���\L�xv��bЅN�'s#�Scb��oO��
=�����p���$%{^h��Q"{�e���Y?ezC��@����;Ms�q����rяr�А�v�3��^Hg��h~p��Jhw��Z�#�zb:͓^�f��;'x�ƭYmX�{r�=/ۏ��1"�5�+ G��l�(��Y���U�9�x�cv�a�k7Y�����Lz��ݗ&��2/3t��߸wf?�`�^Cj7�2 NL���kX��WEἚ���z��Ё�x+��kOvҢ)bq�5j�vMY9�b���@q��n8QFZdS�Lqbӥ_]f{3��|��oW_̋����u8�`b�N���cA��ã�t<d���]�]N������F��V�DH�J/���#Q��tz?F��c�cv}c�C+H�\;2�m�ǡA��Ԧ�{����K���/y���)my�mt��!�x�?FΎ�>��\��� �?��d�Y�2Y�s�3���^{�9�5vR�a~jn�y���&%Va}*`gO�t���x�5�H�d\[SW�z��)���zH?/� ���D�m�����6��L2m����d6�M��Y�����<@�/O���a�7,��*5Y�cF%޽�y�b7���rhʘ<��K��۷G3�`�1��{��Y��[�Z��3��L�R{�.�>[�B��Z���~���qbg����e�v�q9^�~�8���v?�����}��y�VL�~���m�ahQ���[��D��H����S��%.�I�4b��Y��l OYMp������^͑���I�Ԯ&�U|��1]{��4�`��<�0X�ޭ���R�Dz
),������*=�ȧ����+T+��;u�Y���u���-�w��C��x��ڇS� ��҆�/���Z�2�(L'�$�Y��p��|��B
$��_|'�g����Z��_��t�X�	�3�Ԧu%ݛD���Qw]�0Z�.���;����<;�d\n����J/�� H����pks1���������m�-�����:���+e�@�=[s�zd�@&����\�x��U��4� h��"��07�r�g�v�q'٬[��)˃�Q�12�������_���1�\���A�8hRn�҈te�#i�Èfb=T�����,�8����9�^uED���|�V/��Ȼ���u3>_�� �`��=��-����@?��?D�ٗ5Y'�x�V�ykʮ=�;���@�γ�0���U:�Z���e��U���f��\o4�I�^�x�5�܄�^B�#�5�w�3첽9��0�QE�ߞ%�y���tè��m�9�嗮1����Jh���L�Qh\������e%O6��6��]$R�J��ճ����U�>��a`���u��S���.�*��z���ʺ%�	�P�7�lѡ<�}n��F��^�ǈ���r��֩�F�ǫ��ֻ�������zs{ &��7a.u0И�=�[�:U&Sh�!$L��h�W�]i��ӁMU��(�G�N ���� �����,a�s�?oݝ
Z� 5- �Lj�w������^wJ,��+���'�,���0L9�CU�m�@9�L��{�7nA�+��2�X��
���XJ;o�}]<���D�	gKz�#��lx����D�ʪR㥠�o ��̚��ڪ��d<k�nmwr&��]�6����w�FF�ϒ�u.֗A<U�N%
�u-;�zv�ul&�Q�'�n�4+ѭ��MV&�/a"���5�{'�]�M��Vx�����8�Ѓ}�s��wtr+yhe��.��*��Z�ym@޷0ou��U^�Kh��w/�꟎�m�A��0�=��>{��~"�j���\�^�k�o�Xi�ic��>߻�PN�f�H���:��(~�}�~b�hh�#G��e���+�S(��55d]n3��uؿwO�;}co��C^�!Z�.?&�Q�߶Y\�x�o9�pp��ήjͼ�5t%Z����Sz5hv�ݵæv����J����ݍ�D�U��V4�҅g,����J[�Z{R)wq</�����؂"H/U�V�I��x9�ۛ��P�7������Cg\v�~5#_�h�b�h�Q5�/T���	��x���b�}�l�����^'��ԑ}�1��v�޸3�����K8a��r��Y�1�v[�ʕ�x������ ���Du��瘷�qj�q��}h�U��$�>�دbzJ�fcs�3��F�y�t�`p�ol���n%��kk��!r&������ye��;�d���eR����lX��-���v�<����ń�����IeI�E�������F@�����������3S-�i�M43�m��u�)�����5�oZ9wH�9�����y+�h�ؓ���q�y3=���Rjnp����;zk�
<dl�u�m��{\�d&"k�����g�+%��wm�U'b�+ӝ��"�9{�FѪ�s��l����ۂ�����$V���ku��0Vp��b/��e�T�D�H��s:�9̓�%��E�����s�0����c���U.�fT��jU���e���S�]>@՞U��/���z��j�3&,Ԝ�f+�)jB��w�M�#��]Y��I��6��vU�ele�P`��5��>�&�,�c`�ra�c��:�hGkX}���gKd9�T���{�S��㫅1���o/L�$oi*�R�|�q�Jz�*�3qRr�����&0Pb��Q�\V:ݨ-�Y�i�u4��ȷ\U���V7ΡO����rEi�[C0��8��G�4���G������:��w]��S���F�Z�6Q�g����q���gjg6����0Z�M[5�Y(�(�wϦ����ol�y�t���6�t�m�b�[�Oxs�۬|�-<#w��˩��n'��v�ˎ%����y�)�=���(�G��6p];��.m'ϲ����]��	][ĳB�X"��0�C&�X�؅6�h[؄��1���
�d�憇q�Ÿ��F�
�����v%{bP����T�����wk���i͇\\�U�|�)L0x��+��H�2[H�+�al:��ۦ�
zv���8.��_���#��ׇ&;��ƈ1"	�`�x�;�B�{y,2a�AH�8�r[,�s���K�p�Vخ��	d��c�PCf���J�eG�J"�^���, ���O~�Vz땰��S_��֢�cŌ���ԛB�s�ѫP΄�=+���{T4CRh�x�ʉ����VW�r��;�rȦ���R���"�\K:����}s�ל�:�}� ;G�l���:�m�뜦sV�����VkmnA2\��{qR��+���{�_w�%L��ww����z�cmԕ]�8���'Ov�Z-�\+h��m����e���Ia����2훔�bu�c5Vn���7WGu=����;� k	E��ʖ�)|�g��svI�x[��c�d�#,���D{�h��Z���eT
��s�]�'P�o�+�Gz�Y��[\��8�&ϩ��]�[r��W)����]�j`��pޕ+D]gv\��D�J��hh�7Af��d�3ڐ�mߜ�u�s*JnOZ�Ű�Qd���v�l۫��I:ƽ9��$��;�YكF�ͱxM4ތf]�	��x+Hr�VJ<��S�yݢ��s�nd븻�s)|S���
l鬙]:Dr�ut�\b�-(s�\�[�Ռh��Q�2�j ]�\*�yhw���=Ю=o�I��7�eJb�:�F���14����
��R��r���HH�R�9P$����+
Ԗآ�ϭTbe*�)iq�r�2�5]�E���<z|qǷ�������g�F��LTN�kT�**%e�[E[�`KKm���{�hv\���=��>��������_Y��Qs�֡�Uwۃ�E�ZcS�PDq�UF
e�+b�#iUTmhV�����jr3s&���SSSSS~���λ��
��<"4Z)�Q��E#�X��GME�cֈ�\�x3��
���ɏ�{{{{{q��>��:�]I�h�dxKP*VVUk:�E;h�i������"�5T�S����������������g�_b�e/0|xΦ��AEQEQcĨ�)Ԭ���R����� �s%����2ny<����{q��_Y��T4�UNܣxr9j"*��#�5�u���-(��tʻi�A����E2�Q�T*Tݫ5JLq\)J �)1��҈�2��P]kI�1�U�AVL�!ZEU֛f"�h�2�j��i.e˴�dEPZ�1�.�R�N5V"���+D�"�ۑ"0E[jiSyGQ���80�;�4۾�����nVu�����+�q���ȭ���[��	v�����#�� � ����.��t� �+'F��|v��\�+��и�p���O$ɲ`�i�u���������1�1�s�!(�>��m,'�(���M�7�Z��(�B����{^��*p������9�JB쓻KI�&%@�����}SFa޸����s�<f��|_�)C�j�����y����[S�����c�B#�"�Ͱ��|��4�98Uz7����s�I����7����8	��=VqTժ���2���Z���e��	^Ō�3i�F���>�9�9}"y�Tix�~������+RӘS�2��G��sU�(���L�MOO�R�u��;�^U�JX�Q@XZ��$�;ݖ�;f�504��Ygk�c�{��f��r��LWw8Xd=0��ǩN@QJkkԗ]ϻE��o���)����J�m�v1fA��\t�d��rk2խ㔮�����Gnm ���aX'�ɃF�TP�O�4L|�f/T��Z��/נط��JZľ����;�rL|�-2����5�k��ݜ��{�q�^�T B����oL�J�	O(������5�l2=1���t�yj�*���t^��mCM�l���j�����N/:|�\��}Y~���^�+ҫ��'e�`�TL���a��x-`�͌��0��>�N�&/ZBo�O�͙�Ú�"���]����n�yj.�}����̌�C����A�s�D�c���a���̕4/%�Ϋ��ծ�Rk+��6�IqxG���J��n�M����\x�t.�fFu{�JI�D߷W�[L���H���=�&3��A��V��J�� >��ݖF�M��\w�
)wkS{Z��sgRK|�[˱��Q�RW�m�p��M-��6j'k'u���;E1��nz��_tصJ�U�OW[U"+ϙ9���Y2�k��e����
G���z�\�v�^�滑7ת�]:�[�N�-w]ɁO�#d��{hjckc�9�����h�&�db����	[Y����e[��]6�9H��sjW`���3�DK�&��������E:���K��*�@�|;��N�٣�-�R�I��Bz��}�l�v]H�BABAPj�FYNLL�6U�%�mL��D| D EQ3Z������F��>�7�5�o���}�{�Re�O�6�i��^�ض�F��;5S�n@�܄�ҧkm�3�V�}>��K�3�^؈���~i��Vz�0U?\���&	�5��z�m�,��G���a_1�a���HO2{h��[r>�R�J�6��z������q��m�GP٨z8��j�U�f��l'���v?
^WFm^׮������v�k����V��ܷm��V�RKVFmh���fY]\���(B�cբ�;!�P�������6�Q�P���Acn�������>�w��M������)=E��1�/�߈=�o{ݗ̬�:��r�����.<�+�3��A��y���V�6�*}jQoBv��q�PzHL�0
�ב��[("q�i���1z��k�k�������L�ҙ��9�/�u[�S1�QS�F����fM픛rL�5���&;hm����nv�;�1Я�@�%NXj�{~��X����}���PC�weǜ�Ѧٶ/;Wm=qm�[�r�'v��k�gh�Rл�J�hs���o9�r�����?�"�H��ϯ,jU�w�<��Ϟj�K"f�>��tr�{p#Y��m��*�5jdg0���sS{�����oD����>轫�5���j��ݸsk%럺~�X9gwh�gDp�\d��0�� �����:�����F\�AvMSj���ź�ki�������"�~�U��R�`g����0�[��|RlzN�g�1��U�@�ew���TC`��/��<�mZlD�5G�я]�yD�s�q^$̘(������}�6M����<��D�nX�y���
!����t�Ժ��k����Gt�g<V>v����9%
�fk��ݧ����[m1V{�ZȚ�����>��be7Vd�Kv�YR,��ˮ�k�a���ʸ}W=�Yv�n3�ճe*1d6�zxs��isߑ]]��r]��[��3�n���|bUR�ة�VY�|0u�e�V	ٕn��Y���Y+�ju-�Ǌ�툳z���[ʤ��o},Z����e�n;u��ع:���mSS���0��ѹݮ��q	��t	�+΢��V�9�����`����ng�A  ��W�����j��윍I������	<�� ��E`��&��(>Ļ�FP<�wZ!�"LG0�ӲR΋jw�y�w���vѤ��	ذ����������;�u�o-�ox�9�5�(���#*d�Q-�)�2<�����c7����`B�v���vs���P�P%�^�}_}�	�ߠ����|���|�e��70�����H5Q���=���ݎ��n/�"�P��K�f���������Z���#�ּ�ipᱢ�2�>7�ӰM�6w4ٛ� v�Ζ^��6�j�ǓLd�2l�<L �I=�<x1�/:/r;ה�n+$���nq>j��P�2Z}���p����l������#K�p
_y�S��)0��u���t��2�,� 5��wF�	��b�g8_}hn��ߔqb��+;�76�c�
��Þ�ih)��+w~��<�f�kʲ�{^Y�z*���9E��i-���꠿Z6�e0��>pEP$U!Ch�/��b[y��2�v���:mv�-;隆�e��&=�=Y��])7�7_�! �[����n����vo���G�ܐ'��)뀗�C��4�=�UɓU���cbz�*����޺1|c91R�Ұ=?����ַ�3�{?! Z(����wy^�@ 0��3-1�0>��(�W]�	�����$�����W?+J��$ܚOm��6�H���j�dܷ73�f��*z|��v8Ʌ�l�wR-d�g)�箣���+�����-��x��].���,�����]Nxv]�2��.>�9����o��i��s��oO��8q�t?m�L��q� �]�M���G�}�@�%��隆VWZ��3�Lh�X��c�]��n{7�y���5�@�*.��P�%��#���������h$�����?P�#{>Y�b�w\9K��O5��V��)a��[�/w��uMn&&��P��r\g���E�G^�Q��}z^h�M!KM,+ilLU��$N�Yu�|T��}�_���Ч�R򶄥y���@*���U{r��"�j*uAD�)�[��VI�#��5�-�_� o��ɹ�L��1�<�4�pt���w8�܃&{):ɼ�t�\������ڦ�iH9!2�0Bj
h�ѓ.Y0�T�T���cH�H�gY�n��������{G�a0B������w�/��ȟ�}
J��m�ެ3��r��L�U�(鮽���yz�{(}Y�f{1�7v�ןU�,��Eڌ����{[�E�]�|>�Xc��=P����\��}��/��*�Wh���E7t0�<��n�9�̳AB{��~��ޡ˲�Ceu�r�x�rg�P�`��]o�7����������>�կ�Cf�j�,�Nҍꚥ�sP���g�=:�����EH�"'Q��w���d�=>��{�^z ��*�S��&�d��e�\Ee�0M��<D��"i���������5�-�tw��~��e��ͺ�c�l�* $��vWrr�=­��b�j<���kF�{��V����V^��tI�F�*�?]�̜�	��(�߾=רW��1��֕��,�U*�l�nwS9\^�p�}�/D��'r��dޙ�|��]�T`���X)ޔ���$G˕����}��2���_Ɗr�WMg�R�b��X�U�5��O�3�sP|/ �g�sJ	|!$A>jV�0%* �	w�(���fR=:�w;J$ukx�?M�=���(7��SK�KLOe�/i�=���ω�>NU���O7��b-{l����u��;=����X���`�Gׯ+�������E��&�NΈ����_��G����w�i���-�;w�u�̩����N����f�v�H�����Y�y��&��ؽ=.Te��X%���I��L]�r]J8��ɯ0\f��y� 8�u��^\��=���㕭�g�e������
���J��/��߱�Z�D�s�A�hCE(�{�S}qr8&1���0�:6���ܞ9���Eb?cW>��xY����S�ڙ�Z�Ң���8�H�u|�v�+S8�W<�#x�0eH�P���6�{��%Q�k��霭v��\S�t�Һ���L���P�؆f`�y��h�#�>dY��U��&6Lk"�/��U��%'���a�y�Hp��+���w�@�7Lf� ���]��'&\8O%���'IΊ�q�3��u�`�.�T�ųQc��=(.��i�
��JԖ�l~
��1{#�f<�zD����1e��
z�Gs��Y�ݴS��Ƞc9�����V�E}룱�u�qn��q��iT)[�$.���ôX����W�[�e��[�eQ<�=�տz=f<�L�Z�����{�{�uT|NΙS�c`P�����K�N4i�A��!<���fP���}ُ������zl�we�{�f���VfQbqOysk��k�O˻V{7g�����Բ����v
Ɏt�c9���}ݪ�x���oLv�;dj�)�c���G�.��E?��jf�@�h sO�x��+�h\9�ޯ:�5�*�=�I�^Һ����~f4b̍�1#�?A9��L��`�X�暅�_�[�iB�X��5ۇ��A9 �sg��#�ϚO���@�YF�����嵮�]Z�?<�A6���A���L�VO��<�/G�zJ�ŏ��)=��Ӡ��+緗˼ߨ�7�1R������B����-fsx��t%�ab�7�4��Wf�J<::Q��5�,�A� �;Fvp��u�$ϮFC��7�}�K��*'����]JƓ��Md8�js�W3�+�;`H��"�gp��q�$�+l��z3��7�oD��_u�$��ɲ���!ԗK�?��{�H�Ŷ���'w�Ia��.�h�l�{���5�A?|� p"L����x*?R��D$�.��]��b��93G���ц�G������&�k6^��6;\L���K�Eſ�<x��Nͦpپ���+S���㮣�������,��+U��_Eww���^:Q雰�,�J�K�s%��Xs��n�.^���o)�UT����p�kM�W����&�@�W
��٧�!���gl��;�`7�� mw��]h�Dۈ[����˼J�2q�\�[�{�'�Λk�y���C��T)��wj �q/T_���cy���
����{O�\��ϏEX�5:9f͡	�ٷ|�O�Ɲ*bl=N[�J�[y���;���f�b�]������1y��j�ǜ��}�N\�^�+��N�4�k��<������n��c�i���p���t�t̽�j��
@Kݺf>�e3��� ��ӭc�=�c�d9s�q��	����Ǒs�:����U���1�vy�a1.���m�muCu�c w]���|��J�x�qWu�v��5݇��/��y�X���J������ѠߺuK�lT�mC���l�5cN�XgI$uB�a�sj�c�U<Y�������Wp�ݖ7�k_0����r�ӗU�qUޭ�W-��ǵ��u��F<�.n\˫u�h���y��!�&!\'��v;v���<a��3Xʶkxc|��X�_E/W1p��ͮ����N�5����H��F��M�W9�d\��3@Sk������y]�$�f�G�ѲM$��#W�'�h���4nR�/�4�v�yVy��'F7�TSE�K}�aY���Y��(���Xf����K�v�m�l$��������H4m��.�r&�c��귲6�0�&���N��]��d���٫\��p��J�­��HK`�s�*5��{;�,�XCSr-��©y>N�$�j�Y��j��Ǹͳ)���R���~K8ᚣ�}>a�򔶉���6����Nlz^�q3:_�߻�7�o�Rg
�5��.]!�Jp(��O���%h��H�ߜ�i;QJ�S�/�7�/Y��F��n�e*vʑl�u�j@�h�I����$DmH`2�](s�˲�
��$12wf��3�[ݜ�yCi�y\U�ܒ��T�a}bu�﷓gfA.�2�;j��r��[=��G�����n>j�I!��3��;B�����s�;��������m-mL���ŹW��Z����޺Gm�x�`����Ƅ��N�
�M��o=�]�]6��Fr[��{�0f���5��/Y����O�wo��tC��^'8յ�#X�6�����,���E�޹{�,�]��%<��l�x;��[�5�9o1p�7,��ni{ސS���k�˗n������}Թ2������6��fKX����v!PWi�s�.䳃A�:�T�1����ܶ�<������|y
,��f�9�0V�fݝB\�oc�}4C{�#ģӢ��"�X��Tt�
���@+�[+����q ���a쩵�����㽩+��O����,=B�A��l�ĺ��@M�����$:�M��cr��qb۹pn�Q��ܱEڨ���؂�fa��e�p��T@�(
.�H3\�,"qB�1SQ��a����%��H��ZL5^5UN�P �P`�Q��ۂW�ڌ*�f���MI�(���#����E�Q�@�5Lכ�eʍ��f#��4\B���sz�"�EUW����#�B[4� �쬗��mX���:�2UZ�q/:���e#D�v�����T|����tCa�\��JtT�#J��\9�D^7ւ�{��bm)Z�Vhq��]�j��*�"�1��E~OC�ӎ?����ܟ�I�v1�8�4���r�$��1� �QTAcR�̂��n�q);4K2y7<��{{{q��>��;��P{lE(*�s5�Ru�c"2�Pq%��*wo&�fM���MMMMO'gI���s���Q��:�2��Nҩ�5B���6ਯ�-��]�3t�b���%�5=�MMMMMN�gI���w�F"��D��̌cv�DX�1��lDA@D��'�	�'g�ɩ�������u���Ҫj+�<����b�(���m��_|���XaR��%������������������3��DRuZ����hYYԊ\K�
�Q���^�<�.Ip9KRM7a�,1��$D1\Օ �����J��Q+y����A+l�i{�PYm�)X�$�.%T=�f����t�ATPg�ETX�J�F�,����DLaP�u���єԹ��51i�Tr�A��ћ ��:t�5���۱��TVrh���wTӸ�Kl�5���l�ܚgsB��l�z#��(*�Q��MSLZ�k���E%(��D'3ASd<���T
c�^�f\¹��I$�DF{�Nw��o�z��'TN�;�q��v�7Fi��2Nލ���Qo�j����z;A��	u��A��dt��c�Y����g��}�[3�P�Vo��v�L�s�3���z��J��3\�<���P��F_�h�@ͤ���K��Nq�&�z�M�"����n�gi.2�K��������˞lY���p	�	�x��[E���A�k$���/:�d���Ȍ�q�j<���|�e�CӶ�~�C��T`0�#������8���&5tؾ]�Y��zV�-�,�]ϛ�@@���oo�f���fK���"D?d�{z2I��%0�`ga�\��/w����"+���M��F�S@Ϲڐ���{;�I߿�ϕg���k'�x<�W[�Y�~��`�}�Z���\��Qz��(9�ג�k=K�˰j��M��@���ί#mEv�tM,�� �� Q��M����n�o��A&�]rP��v�g&�kU��k�c�4i��0,=�q��3��h�z��_~�y�����+~=�!W�bBdo��������0a�2KU,����<>���5�rs�|���D�NEXBg�i�e_q���c�x�SM�]��ݧ��f�;�^�boy[�;R�&zo�i�powܧ�V.=)B^��͊�`�"�z�~����7kw7s����e��*��Þ�,'�إ�'�eÑ�-o~����'� z��m�=e�J,t
��j�9=�X��r�|��<s�/�a�b�8p���j��{��v�%��I�&�_p�=�?k�ϫ���V�ufoc������:���Fr�д?��w�=�0�h7S8m��3��j�fdn�":|�U���[[��[��'/F�
�Z���}P���ă�S\e���1QD�eY��ܜ���gf *�wӊ�N����vMG;�+����Y�R����u��݁��E�y"��ȹeM�z�p�	�#d�UJ����"�Î�A�ܯ.�4���>�W�|�c7���#����Uk�j>jS�u7;d��&��{.���~���#�݄���DB A"��������u�|����2�1����:3Xu���$�&����攘��P�[������b�\�x�Y�ys
����G���W3؝�t^�F��G{���c=x�2�}�5x�I�s�T���W�
��ys(�]��t�ں���⹜"����C"�zt�
�T���;�Y_��H�|�S믨A�����kޅ���Ӊ���b���(�M�Gg}10 i���U
�O>,���(��}�~)R��%�m��ũ*}%�
�˒T�u�����o5� eY�UM�����L?w;	`/1���{��0n�*�*wǫ`�Ɯ�'p���������z��
"ym�x[lytt��	�U��WWKU�z�]s��
1��W��y��̓0�*'6�wj�c�m��<K'��ͧ��5�/���[ƻ�Y2�x����)2�S�ݬ��%�]p�d�-c��h�;���l����dtqV�t	+6�1\S���G�.;]�g+���[���Y��0��.������*��XޫSrٸ6$5Qs�g��A�E+N�K��������� jH�x���0��8��0(�y�ێ��Ek�)\�r��m�C��ֵ�����%��<��X�>m��7_�\�0�9uJ� �H��{>ߘ�<��%{���	��#0;ovǔ��U]xl`���5�ܠ���Y�z�.�C3��T}K����)�:Z�U��[�_"�A��UϹ�^�XY�����^�&<g} �fP��ɭ�ܽ�Q�{w���1��0̗�s�H��=�&���,������DM�}h�f4�m�p}����6���n�ߡWw@�>c�9ocrZX���j�;�Zd�
�t�7@��Sć�{� �G�\��(1��������G���4�|_�h�l1���MSOY�
�毨т��*�F��K)�^>��һ'�gg����z�|��Ѳ�M���M���=�����-򓶀�
_]���8�yj��>�C�~zUl
��<6!CO]6VUL��XD1��O�vC�N�c�m�d9D���^�^6*��R�Z0\�{�J#K��m�1p$����w*՞���\���5��L���"��#�D��� ��&hQj�
t���"���"�B�*���fS�
E&�#*j��W�핺5�0���/��T�1V��	�aIwZ�du�:�fj��������Soo��=��h�b"�0��!W��u�
�y'k���4)���P���r�}�/c*D�N�y�h�����%h��ڍ�J�Q�vޛ��E��ja����E[��7��\M{�Ësؓ�z�i�8F{Z���ݾY~!˒h�[�<n��;8�l_��ٰ+�[cwz����o4�%y{��>�q�2�0c�YT9�qX�.������$���27="��ӕ��0�Q��hNN�7�:��a��������Iݠu�Y�~[��?~�"�����Y��V$�e�w���v5��Jw3%'S�o��~�K߽p}ϱ��={�L#�a�k/�utF�vmt�|�-�#"/��vU&�}>�-�_c42�}�VMu��ߥ�λ2ܦ�`/s�M��y�FH�w5|l7���լ�����+�	�<�����+4��/��(f���7w�N/��,
�@`ȫ��r�M��X�-T�w_�A ���kz������^F�y��ು�8n�Η�ߤ�sn8����m<mq&_s�W�d��>x�A���.�����}���q��0�'_U4����C�b�|�A.-�x�Z�g6e^�Cټ�Ԓ�O5�����R������x!��@��f�Ȇ�Z���[>��I��1��B��۹��j��;��FX%,��0�8R�-�{�j0��ko��d�ܶx�m�T1����Z����۸^T]��ň`���G����}��Y�d�l�]�9l�~1]o۝Fr���7� ��=u��\We��%�PK-,t}�/)w���]�����H�HM�#5d�������tOʃ}�/z�b���]QΎs7�P̖p�uO>�v�<?f�}`�� ^�+���2%��0�w����2e#h����mnM�yG*����������J���t��v�����j�/��	����;�\�a��N�nG��}���y���IÑ��G&Sgz+�D�P��+�i,���P"1(�D vT׺�RĽp�@��kq��?O�I����V�a<����k�NfM��i���{�>�1�õd�o��ȮU^�� ��J�<�b�m� _Jܟu�s83\l���=�����n��E�N>]��]F�G#��s���[*��=�E'4����Q>]�?��L��Yӻ�0�BI� ����W���`b�l�VvhƓ#v���dj���Z`�h�S���N����ǤX��o_�|��jw��p���5��]�R;��H=8����\��#O�[���WR���v��0�������(�����P���$����vf`�8QI�fE.���-���Em�(�LM�mzwY�_�G�#�珶��3�}'ґ;uw���]&t-c��-"�$�c��P�����6�-�i��l���p
��m�F;�[�R��8�_v���귑�Q�7Z� �g��D��0+~�,xn����6շWe%���[�([�}f���1��7�_1��z�ͩ����uk�,�8��0���/�����LoJH|"��D�!����\���Z���>L���!u�z�w jу� �UhI�����GG+p��a��w�X�R���1ou:��=����1q3W8��>��%A'W��1[�s��&'x�,cվ<�x��#3h1~m�e��f�����.N�j����*�N��h��:+Mwv,8�4�Ӓ_Ӌo-kr��.]�t!3�ݩsr�U���
��`�[{n�ido��)��j��ʦyU�v��'pğr5ro��["D��u�lTg�����M�{Brtm� kD8v�;�7�����^��?f��zQ��|��H��#s<z��?�V�I^{Z����p�PE�y�}<����/}J��Z����Պ�����?tȃ�����n]���b�G���M�z|kz\(y��=�U~��AjC[���V�^�r�`�Cϩn<�oLӭ��d�Y��}S�:;�(���"�F;V���C$� ���Wd�EH�A�ژ-Kb��;5pH���=�p�jA��L�Y.ow4��{�k���>��"�؛4�{:�y}¸�0A�ųB��:��&*�>i6��.��ؚ���9!����,�"a����0" A"��J��Y��{��5��"�32�s����(f�B�L����g�`��v�ތ��f�ۓ��&�h�0�L[��b��Ȼf�v��l3>���#T�4eE<uE�V�^_�]l��<�l���Zf��-����:7��]��;�ź��(��+a^�=�s|�8�ZM�]�)j]�utAcU�1Y|R�F@�D�
��o��4�T���<w �L�=�9Ѹ8�!�΀��5P�Ӄ���hY7#�UT���`��!�� ��P'}V�tmS~o^�ol�G^__lV:�����X����;;����=W=�1ӈ������H��߰O����Mr$~v�~[�JCqXS;C ��cx�VŜK $oWr��n` ^�{eK�?D�2�7{)���6z��uz���1�+�ϖ��]8*yK6,_�͏}89������U�s�2>[�9ɪ���K٪d�=��.����Nz�g-��0q��H�&/]��u��]���g}�t��v��������������ׁV{cYV�L���}3��}T���9����� ތ�£�v����/�{����_�Z}�R��o��h�3z����_(�˕���b��՗�(����s�yқl�E69�/��dsv�3r��3s�p���׍Q1f���~�.�ή[��*�)Hq�@#\5Q���7b���ki�����ø�im�bQ��P��<��<Ѱ�#v������Q3�F��̵�u0Έ�p�� jϪ���3��>֟>jJ�-R^��]����a����uyW�E
ߟ�(�����n|����w��h�愶a`��J��}7ʽ M�H������9F/!��=�:R���˺�߮C�?{�m�Э@?zd=�L�\�t�퇢Wt�w�Y'N�
[F_%ŷ��Ͱ��s2;�b���7�C�E��1h�[yt&��{��{�;Mֈ�9��0Yh�k'q7�cʏzfļ=5�UC��z�%@5�y�oϘ`�4+�Ҩ��16�78ݸpWr�+M��u��윦��`vn�َ�n�6���ʥzEV!���<j$Y�Vs�]B����1�B�*k�C�r��� �([8��j�����3�[��4*3���x�)<����|jTfWu�I�mӍ{��r�7hm'��ڱu�re^������%7Sw��f��So*����2]�]�#��e��9�M�O*�T�[z*��N�nX��ٕm#�j��]F��9�=9�-�q-�rscN�:���K�������V�4�VN���s�wA���u»3A�ŷ�ue�F.Zp�se�Ȕj�e{(r̘��@��]�G��PQys�2p��t�*T��b���h�o)��X�5�����.e�B��#ɹ[��*�����Vҝ֦��k{��w�8���mv��!��i�`��{����7܁��Pi�Q��9�b��+"��`�)jW/E�_!5_w1����I�
ڽ2����:�����Ϫ��6_���{-k5uK��\'����)��U"�)������t��8h�6O
ѳD�7�Z�P��jKg�P�2.����S	4e���uxřu]����5F���	,I/p�u�D4yۉ-0�_�y�^��w��ˑͿ|���
Yn�9����Nt���/��hbDN��ц�f&Z��ۇ��+�NJ��ن�o�����u��Lí)v��ݗ\f��}��s�[�`���P�)��Z��G���.u1b넾y�6.S4rU�M���v,ݻ�{�H���+zo8sA�wTR�%R_t����Hj����^�Yb�g>�̲��n�0&+yo&r�ك3u-jM���n%�a��yK��[y�>�/)t�@KKD\�6��Q�|�(���	er�u�W��Z1�N�Rw�O /Eƺ����Q��������J��+�t�9v���ڦ�}�y/��{G�Z9q��:�X�lR��Z���C��w�����mN���f)Ww�S�}�cW�9�T��|X�cc��[�E'#Yv��h.���ó��%�Ȯ�f������$NԻ��sx��$�7hʂu����:�h��N�-�ڣ�^v��+��җ�N�ӪvWE�����2�.KqC��%r��Z�^��-̵U�po�:�Fݭ�D/Yw��]�]�mN�u�|��ä� ^��(\���^~�z�*���E�(���z�x��.�ye�C֙cJ7K���S�sɩ�������XΓ���ƨ���Q�������x��8�� ��<p�ŋ�	fMM�f��������c:N���/l,��V*�`)�����C-�*wVC�9����������������G�v��*X�4�X�U��y��E�M5�iU:�Ƒ@X��w����������������]8���1r�j���I��"I�e�Q��*��a,ɩ�٩������챜'g�rurd�Q&	m�F1fXPF"�J�V�Ϧ̚������������vp�'X
E�{ltXQ"�ё`�@�m����PE
��i��0�0�!�WL0V/T�*3mUb���*�D1��-�!P1
�7e��]���NaP��LJ��Ex�Q&	��\t0X��Z���Jʜq!�ֈ
�Ɓ�	'�$�S�[JVŖh��`��sݫ��;�=[��#�v�u��N��<xg5�7�K�".�7%>TW���E	A#7����׹���;���u|,�]F��*ۆ���+�����H�m��:F=Ǹ{Y�wUy5��2����˭�fF��S��h�!�oA�	�c�{8#K�8g���
��E�v�o/t��Y^�}��3��D�w<ik��|�;���2;7Wwl{3U�4,��X����V\�p��=��H�H�R-����P���X�k�{\W�9�f_i���oh��y�zX��V�$��T�tjr�|]��� �1��a���M��&�b��R ���������s*I�Ec�th��Y����-�c��Ŷ!��+i:Q/;�1.�Q��!\c�{ц(��b�G��'���E�+��Ϫ�;��N�v圀N)��O���/�B�ӏOU9;��WAA݄��}9�5V
�'�Y򍬆7C��]��#�ڭ��Oe6�H@�7��'3Oo�����/�T���.I,�"��g�{F�?�0Ň��W�8�/�k��>�|e��YK:%v��{�K��V�k��{����T�J-]���pv��C�H� '�n{�޻�:��G�ި��}:�v�D{Б`8��<z��#oN�"'�꯴O;����M�l3�5���G�/e�M�Ɂ>�.b���dL%H���;�i�ɺv��3-F̹��C���x�_Sd��~����^�4i����e�FjķgT@f��L�CU��дj��2R���mU�/*P+#Ś9^G�H���uA�1�=Cm��K��v���T{
�R���V@ɖp�䶎�܁��)Oq�g����h2�β�%k���%)m�l׹�Pٝ��;{y��@�f�=���Y]l�IT�݄T�[Ue�Y�;H2;˽��޵>�q�K4�CE�W��og�j�0��i~�-��0g���)"i+���裶�2��ͱښ%K����ܒ���M�}ǵ�f9�V���O���N�>	����hn���i�g���W��-���t��`��j,�ҡ����a�'�IH�t/6R>n턩�e�D)HbD7/-	4��D���� >��k�^{wW�˽yI@$�G���ch��7�Kfdɑ�-N��Ր��l�_[����@v�J	��'k)d����梪�r�	�,��2��N�B�{7���8Z٤˟�ě�$B"T�t������NE�H&مu������,ͩ���W�"aX�lox�N�=㕛X�\�;|gDV�Ak';�;��;��B=m�A���Q捚DUj�tۋ}��fM�Lv}�@k�G7����e6�T1;��ʂ����t@��<��nŏ���cc�Pm�=�39�M ^��?��66x�QǬ�3��#��s͋��3���]O����N���q^��u܅��%�pU��]��c�򮦷>���tc��Rnv��[O��+E����/�Fs�1>��\'U=N�qK+o��Ɗ�Q��d7}l�ES��FvERͺ"�L�[R��i`�de�}��dʩ�߲�=��A�����j�c���:ZLp��r�����;����5L�L���������3�=���y�g�4�o:����P�d�$�{kr�[I\L�ǡa��U��Z[�R��ف���ه�"��O/JC��a�G�@$X7�FL�D�q*��ɴ��[�d�R��'�(�۰��m�|,.|s��c���8�3G�<��{boS�e���f��z��e��t*�)|ST�V�V�1�M�f��5g��U����D�0a��THՇ٠_����g�c�Ӻ�5�'��Q�eÛU5r��[�eLtwo�84�c�wq�^�����f��f�u�����I��*�h>�����Z3�ͽzA�a��]�ů��'zSD;�K4�[�ӣ�V��*��>Z��M|��{�ߣ� �O��m6�"�$�Pv��2��6g�q�s�ѷXg;�=G�y���p���Z�����V��A��p�~߽���)�����0 } ��� �I��s��)Xr�x[��<uz`v��R,�@��=������Dn��3m�Zo9)r3�`b�֛�⤖��c!N�P#�ny����������ö�2'����2>����H4R'~��Cf��<�Q��U�νi�;� }1k�7��`p+ͱ5l����)�����h�v9����j���{=�7����`�4C  LA���yST��C(W�ۗiR�zY�k�q�e7��ʝ��e�n𷎬�t��o}o�D2 ��ݾ����]�k	���]QC{댎CH3���Rј&� Sd��M����p�p_[�S蚩�P]��^a�����1�4��J�,n�Mf�߳�0��ey�*G��zd�/���`Q��d����u��T��G�0�"}KX5�O
����]���9��*����c�L+B��ۙ�xY�0<7�M�Kl�H�w]��}��葻"��W΄��j�L�ހU��u���5ԩr7q ����T�f��K.՗�Q�/]��S��׳ݓH���̲�'�bx�ی<��j���a��q�M�|{�, �Kr.B������~q��f�_��im�n���'l�|0՞��$vC�l�a��<�a���6úm���w��o6{�Zxl�[�jZ���;W�1!����Vд�=EgV�݋���V
Hܟ:��ˣm���7�������2�$9���&+]�y�-�@� 2#�$ �
�Ne��'�6�<p�E4܃�uwOr��]����U	�YX���}sf���)�'Y��y��	"E'��]��/��֧󿸺�t�
l��I�0�+'�7p�eɮa���p���ƩZ��������N�u7�enEl%FO��(읈=-����c�:��}~�q�͐�@��)D�P�)��"�����oJ:�	����f|�	��T��)�g9ٽ��-�Cs�l��q�1�ر\��V�`��\Vk���h�������X{/S�I�`3iM=S�-jV#�L?��q}�E�)
��g��u�����$ ��3>]�.}�('�M�L�a��1�3�5&]�"h��]�l��J���Jf���q�V���,����&[�~���^�;�6I�I4�3t���ُ�!��F��(	��2���Fzk��c�V�Z��s����Ȥ�XDϨ�3�q,R3��a���6�ꊣ��՜p6
\6�|u�X����ԯ;�WG4g�_����{�G-B����;|F'�є�@}=���7��c�4�tƐ��W��ۘ����e�1�l��d�#(�6p�(c,�n�	�gr���[��Z�RWl�wL��c'f�и�����,���%�Cw�8���]�a�l�V�Uc wZ4�#�ݐ�a�ֶZ�Z�$�Y�4M�4b��sR��""��	�v�'���o�0�;/ա��"nۨ<zs�O�<�E蚞G$^0�U/�n">C5_j7�Sa��5p
�bUQ �'���̽�M�`�����M�B*�Q��R�%d��p��䣫;���-����Xke�1�?�1V�s$��bk��P�:G{���9A\T�����m���c���_.�����y�d���S�fdbc<�=��u�*kO���ح�G����ƨ�6v��!7]������{l�0�Z�G f��S��|�,Vb>���>��.��<�����g�Pڻe��M�٩�_h��7qFv!qy!Mo6zZY�?�8��ݘ��Օ����LV�a`# ��3ٳ�&ql4[&d��m2S�k���q��x�����
�B����q���Gq��a��	U�fC��sw��Y���u�A�ϩ��`.���E�2{{۽�`R���ڥ�]�T��1�:�֚Eg�)c��ߺ�D�˧����X9�߰d�ty*��m��� ����"�'Ogu����CQ�s{wV��^\��]4��(V��rp����ʺ����k	���Q��p�Hc�Q�m�jKLs�i��Ǧp+�0I�f�A���[��:0���u�U,!��v�Q�1��a�h�&R���b�ҭ&�J1�cv;6�CV�}w�`3�������ޏMwF��#a--X�i��"���K�����27-�4-�]��!�Wu�l����f`���'
�V��yuG�/d
�RU�R�xw��}OU|��y��v�l�Uvp�`��&5kWr�H���8�{'ʅ�W��\�� �@p�F�L��s���38w�z�V�&��CLs�u#�ܧ��D���`?�|[x�g)��=�o8����r�0Ë�����q�|�	u�!Z�3�]����C��u�d(��ٳ�=��3�
��[t_f�U�3n��
@<قZ����|{��
�����+ԧp!��|Bz?D��j�/c�Uu�-nw���s�4�-��2*��ǭ[��#&������\}a���&���X��z7}�7�U�;=%%k���g�v�0[�[�{��v��p�hWW\ᣖ�UDoz���������<'��j�����m!P7��>�m	oKK;y�����΃�Y���Owrۯ,�L/M�/�6|���-�Fpv�x�4(���>#�4DA[�>�O��M=���R붝.��2}c��s�5HU�L�������+����<����M����?�$,�S)?UW���[Z%��l4-�2s�!�u߮�(��MD��#C��9�\�[����F�F���l��� 5sz}/g��4�Ug+��~x�SJT�j��Z�2A������+h�,�^���'}B]E_�V���4��v/��1q.��t-a��%r��+�u�f�27�������Ҝ�J��v����))%�t)���v�8m��^y�m�����L�fx��Y��j�zm���x�** �N/��fGQq'�bk�ﴫ�i:���i���t�y����t�)u"���b`�[�O҅�H���6�l_�Y	����i�*�u5�7G6v6��G*�κ��l��0�Zc��l�8w]:������xzX?���IO�֥̈n���]��~=��L��x�e�Q��il1�u,��B�OG�d5���#�<�����7^vԼ��"%�gV�X,^\!�O^�El86&{�ꃜ��"0�.������^vK8T�`6L�5�گw�A̯=��g�z�	��z�!�!p�<(S���x�z3O��^.�g�����Y>����h�P�Z��k��ZZ_�z��{}~����ս;�4E	jS'�ʺ���aWԫU�A�k�/ ��kf������zAS)�6{=�37�Z�^�NT�s*G�\	�d:F{;�P��md�;\L�&`�;�O|�����S&�:&J ��T��H��ՔAʳ�ĝԩ�F��er��E�O��Dٷ��~��^n���<����?��g�?E��q�U��` ���?_�_� ��
����΃��@LH`�A�����!�@���+P����"�J�!�����*<Ua	���XBaEB$�3��	$P^2,H�%Q� BD�B @N��{� B@�W�P��*)�J�0!����� �B���8�*$B�!"(@�(!��Jtʈp�P B�U���"� �J�!
�@���J�!"�@�"� ��
H
��(�� ��
@����������!
0! �! 0!(�!0! �!0!0! �!*0@�@�@,@�J�J+*���B#�}@� �������������B!*�!0! 0! <�p�A�T�	�	T�	T�T��	�	��q�<���� �� 2"���~�=���>w���������������@��?�������߁�������,����AU���������A���� ����?@���i�����p� ���?g���t�s���O������`s�P�P��
��x����"+J����
�@��+H�B�@B�B�(�@�(��,H���B�L
0J�#H,�L"ċ@��� �J�-"� $�"�"�(Ћ*0+,��H�*2ȱ̫,�Ҍ��J0-"�,�@�(�B,��"��4�2�� P,���,�3�J�"4 J�,0,ʌ	
�0,,� (��,"�0,)"�+2,@�H0�*�#�$�*ȳ*ī0����@��3� ���,,�3�$��,�$�J0@��"�,�J�Ȳ��(̋�2��,�Ȱ@(�ċ2��,*@�ʴ C�"̫*�,�,@�J2�2��H3�0,�,��@�! (�,@�ī-(ʲ-*%��0J��,H��+0
P-����@"P@��"P-�+
�K �HR��
%  �+�� W��
��J����C��C�������pDQR�PhQA�T(���9�����g�
�����)�����*����������������������_�AU���B~�^�4�*"
��AU��?s��� ����z��Q\��?��5d�}��C��׸	����t`v��*ߒ��?���"
��>%��7������?C����������x�*����J�����~x�aI����8~`\����??��{����I��x��*��0A���'?P������/�����B�/�=�p?��^_�������_�C�O��PVI��]�r��p�v` �������?���%DU
I��D��)�R�D��*��A*��D(DT��!T�T�()$QJ"JJ�
$�T (TH�(�E%"U%HR�
"*��B��( T�)R�����(�@��(B�%*$�*�R)Q)T�1
�ETR�QEH���E	(UQ
R�
IET���%I*UDT(U%���Q	T��
()	B�R�L  
�چe��F��%��Q	��E5V5l[e��0j�jjU��-J���V`fm��5�bU�kF��`Vک�5��e���٨�TT����$8  �P�B�
;���((P�B��Cp��mqZ�����e�
��,f����(ڶՊ��m%���mT�R���Jb�bkMV�b�L�1R���"�**�P�
�H�A� 3�h�%[6Emm)m���[b��*����h��E2V���kI�j"�V�a5M-�V����EUUP�H��I"�
�p  a�f�6���%hij2��hh�Z��Z�Z�S-���ҍ�RV�Q�Um�L͚�Ҕ$����
�ID*P\  ���UST2�@�YPT���j�ʓcbm�)���U�%QVa�j�Ld�	R�e5D��X��U"�����V�TQ�  gQk����d���M�504 %��P@B  cK
К0� �YXR� ؒ$B��TUUQ(H�  8�CM�CP �+  mF 44a�@f�
 cU`��Y, h �F  (�����EEPP�B	QJ   a� ��( ��h
��� �  ,L �4`  Vc 6P� 6  �$IT!"T*��  ��@f�
 Z�� ,��P������X��id-�� V�ɂ�4�56� �ڒ���*��J�%UT�  �*��`���� C*M e`)��,� M6��  &U�Cl(&�  4m��   "��M��) @��a%%)� d��	�&i��~%*(� "�L���  I��hʩ4 ԪR��xLn�p�MA"����B�	TX�"�,ֈ4{���X�?�}U�$�o]_� II:$! $�� II?��$!$��	!	"HB I)��?�/�?ͯ��̧������3h���,���^�5OL�W7v��C�H�	S{���]+;Y`��&���hKr���+Ѻl2��S���=��/[ص��d��Ь�3\�$�QLA	�S;��a�^e�h]�z
�sE��5���wJQ��nP�|h��aiY*�J����k���z�۹��;�F]�Ǯ̩sƢ����h�
aKp���������q�0��Ix���h��XȰ�Z��'��au{���=ջ�:�R�q���-QlJ|ܢb ��n�ʓ�m�ȯ�q�bii��ך*�ʊ��ҸC��ad �$��5Y��ћ�@`O1ИCtC'�[
�Ɗ:ԃǲӢ���p�r�Hi�z�ϋ:%It���o]G}���'�]�@`w�p�(]+$D�k.�Z�W�S7j�G㠒�Rd�N����V�bN���loR67/ڽzvU�;S6��<˨%FV8V��d̀e�ԙ�̊�l
��"5���aC��aʕ��A���y-�����:KoH�l@���n�I�O��lF�fQ�Fbj����!�Lr�-��ˬ��z$�{�Лm�ۤ2<[�^n�v�a'���ט�t��i�2R$Ȑ��4���;�7�m��ʺP�z��sP�vU�dJd�[�n�ЂA=f�*Gu��ڭ���ë���qbZ��3�Z���(#����Qz��5]n�9.ݹ�����>���fA���h։xk`]+N�v�QBV'����ޠ����4�(�Z�(�%(A��I��3d��/UE(F���b��/];b�QGa���G�Tt����t/\��s-6͵�H.ʬj͸q��4���ӓy�[�coi���]�	��mDOm�bVRSv��A��a�/v�ŸmSøvh*s C	ܵt�ZE�^���YT���q�B�&n��lX�R9�hZ�E�޲��I�aW�!����s5��kĊ��Q]j�I!f��F�����sP�3Y[�H*�ӊ���ĄnZ���&Kk#Ge���tLi��t�7MVB��j�5J�aR!�Mg �,Ĕ�D��j�ێ)Q��j�ܽ�bS| �q��	��b�6��sH9���t�7,U��h1N���c2�
��i�4��j�k\R�B�-��V1�3[a�-�bc3L�b����;����F�H�F��0�� hÊq�������J6֫I]@o-^��Kv�J�mV^�aˍܤeZ|M7:�k���vCm[	�ʒ�!�&եV5�R�S���
tpKh≡
�5�"je��C1�X*E�nc��§F�ɒ�-��K:��\9m���?�fC��b�wvw�u��(�-�6m��Z��P��*����ב4P��W.!g%���­�>�i&a�3 T&�X%�����AZ\i9j�)XlŔHUխ�Y�^f+@h�֫K~6ʨ�[ܫi��ڗyhiKTYpVȶ^5+I�v� �sD��.J��4���F0]�шf�&hLK:l����=Z�´Kw�H�4�,Cm��է����ɩ��H���E�*e2N�'hF(�#�V �^F�"�i�[���V�HͨD)L5xwQµ
-�U�񿬐�Z�t��9x��D���2�
3v�oA��T�XP����F��n5WZ��k(2�V�tQQ��Vѽ��q�ǌ������ktv�&ڋ��(K��9LJ&;��8��۠a�Le���`��6����k�Du�Q�w���^ފ�W�(Ƃͅe�d���r��O��2�7c01d;.U$�)��[Ux�!��hЩ��ʼB�8�@5���XƷ����nR�2�RrP��K�K�g1�,Y5e3J�Ҫ!��ҧz�Ly(f3f 6;xY��ҩVR���V�0���B�Te����,
H��Kk ^;��sZN'��o\x+I���vö��!ݼ��C$�n�+��*J=F<Jhm�=F������ L*���eeGkIW0����v�!DQ�3�ot�I;�1=Bہ�?1�ݷ"�p<ݽ�kW�`sFc�(ݤi��d�Fe��,�+F��B\H[yL�f���mh��Q�� ����l��bd����͔­� ��Q�T�ۏ6�*���V�'2�@���.��ٲ4��M<w�C����B��
�?(�#b`p���;�l�(�f��Z,J*)\��Ųiѫg��W jYi�$FEhb��r�)֫
�,YN�n�1�J�͔�<I�ee�sݶ5��P��a�t�5�Aowr��feEXlm�Q��n,�՟8*4�
 �4K�(��K���,�zp`C20�&��ԱL�T�˺Fm�k�@j�Zjm�[{��3�`9B@�5���@�N�dcbOg���PX�@P�tVdʕ��.�`PZt��/d2�㳫1���i6�yK.�;SA��x�M6DX�c�Z��H��BZ��)�f՘r����w1(����<���4B���{��f'W�eO���+ңvݷk�V�Rx��OB�V<�
S/3*���3Wt2����F^�#tv�h���V��v#2)���jېV�*��*G���,0dаIv^܁�Uhۼߗ)�;��R�����5��ku�D%a�A�C�4/�eJ��0H��z,=�	��6ܸ����N!t�t��c���F+��6b
�W�$��N-�+�0Vًqє6$
�B�[Uv�ƷkC�@��U��lS�>�����#��=};��j;BؼW�TǓ6k���4H8�ȓ��D���!騲��U2EP�bچ�]^��h�U��(]<�{�1�@�U��(mĉ�38� �_���Hj���l�F��%���G�u �[Wi��j�h�(�Z^�r�٨�b�q*+L^��S�� &�v��	�7s2R7qfn$��q��2c�Ā�yj��h�!U�N��q�l�W":�t]l����L�f�CPQމ!X&b2��$�Ҩ���Z���S����5`u+mR��-Zn�'J���0,���m�"��5�,�H�Nb��wk��%l��Z�)�kU��U�em���wt�J<14*BуN8�i�҃Tu�+��X`�[p��� eK�����˥n!`�N}�@9Y�]-�����Z��"�q�$cNQ����6����߮�ʻYB��N�B��#�!�&�o�pC��ͽ�J�SCa���b�j�IҥN-'oNa�-Yy�r�ă���dI&�������5,�uKC*�h,�2эLL5�\!���I�sfKV\����n�ˢjvRun5���U�NYP�!��fǔ�jm]��/7(�m%�^Q���])��J@���va"��)$pc8�m3��s"v��v�0�MY6]+D1�1SZm��<
:���n��V�Ey�PW`۬�&�́�[��������5��:1��3)�o0�w��`�n��sf��bn��F;���Y`��)q��˩H��U������TSA�)mѤ�ͱ���P��My�&���y�v+�2J(�b�@.T�B^�F�q-�B�E��֠������d�%+[��!W�p�x0
��7I ȵ�M^Tb��	�i�:ʒ;��ĩ
��ұl�6�4w쥉ZlVA��-Mכm(��Q$
�2��t�7$�x9���oi�s2�F*9*Yw��J���.eD��r�JM��2���%}�h�ܭ:�4�9Eƕ-�g7E��v*0f]C^�#��e�o.��w�U������f��B,�3%Ħ����KRݍ��S&�f�o�V�f�����xFؽpb�i���)��˸CX-�i2�U�9Op@CSY�tM����
ń�ה�Z����]duhl�(�+���i�G^�`��Z�4�Zz�J�ͫ�ФV�`M̥f+[��UnM��>��ebOe��%Qhՠe�a��|5���͍�`��i��:�UjZ�Y�*�o6d9#?;P`&��n6���R�(=u2�Q��񉸱�rh)G��"Ĵ`��Qvr ��#)k4��#w�`@�ڬhP��&�Ô@�0��N=��.� U+�����Mm�m�/+b��5�ZF���ޜ�4(Y܌'�Ѻ/B	�q�0�m��9[ڛ`6%*@�wb^����Զ�C/e���F��Rɋ&��/B;t������m��)VwI�A�_����){�{��Bq=q�MarH� �j���Λ�e`!^L�n��"�V 
�a6��+ࠊ��fH5mV��ea��lj�*[*d�b�ݤ�S���X'���������[2Ӣ���hh��}�t�)�3Nf�\;��dǑ�r�]�=i[�XLyqҵR,\�̌iZM��sh,��ȱX��d�9�)�h��n�9�d�W�)Oo^Q���b[D��6-<�	YrV��^;N���mmb�Q��մ�ʌs2HFYVX���Z���A�ۂ��%M)�D9I�'oQ�@�5M%��yn���v��%�*�@�[��
�<(���s�wr�
�D�F��2��q*�W&ָ���݆�����A��v�t�֤u��ܣ�J�����D�Q�����+�#&F�.�Z�6�ɲ�ŎF��g1KV�5�p�xsm�
�啌�#d1�ݓ�G%:��p�)o2�6/kմ��� �.��;Wu ̜����@�� moT��YP�f@գf��LQ��ؕdf�;2�����K���Ol�V!�N	@]��aze]�+Z����w�����2�̶��8,��!�`Q��a1d��[�i�Ɓ�-*�ϱ�j�Z	Sy�L��y�k4 ��fSu�Q���e<*Q&;�i(���F�
�4��L����1��g	�8��U�fP&}�L���X@4Ćf��%fM80�	�X�qo/E��O�bF�0�J�v����L�o1^��;R���b�)3y!��4�2�U�N��Oj�ī����Ɔ��-	�������T�n�;�w�h�l�����t����>�?
��+���L�8\����Q��Ԣ�S��S[��)��̬���IX��ae� h ygY�H��� �@K�`��{f-a��[r�9oh>�k2(��X�E?��޷*jwB���1��k�����,�+V[�Ӡ�
m=Ȫ�8��rct�W�kݨV�W�fe�W{XpT1F��n(Y���,���n��)e;T�7������lռP55+�a��P� �,�Y7jo)�-ZrG7bO.S@e���f��sr�d4A[j
͒�,��28Ek��F#G!�E�)n�Ad:c"(/.���g�p�p��A�U�O+/R� �7N,iJ[n����n���iÙQ�Mh�b\j� �૵)m�U�����d�%]�#CJ�S2�e��Y���ʑ��p%%�����&�e\Jݝ��&�F�ݥn��W�N��ԙ1%��3V�1e�)�X1��k[�鼍eeU��R&
T�G1�$�{H4Ѻ�@����huj����7��omQ���c6,�����d�Śo[�X�3�J��-)�ie �M#q�Ôf� J$䡗����N����Yuj���lܺq�d�N���i�űnj!^JJ9x[N���v�ڠU�f첮S��}2��Ky{%m@�2�;k+���1��q�7��wOJ�fi�a��W[I��T��e�o%�
�@Y��ZM�ѣC%mk�W�B��dN��5n`�#1�u`[�:`)����X�l�|�Vc�9�̘@W���M*�j��V��F%/r�
wW��0��]e���I���jĤ:Q.%m��x���.����B�'kR�SٯN���j�M�n&��V�mf�m䶫��Z�2���{�:R�X��X7FU=� �!��c�$�m�41d����ZĽO^ M��u��[���PY,<�ڐXŦ�;�v�������qfBi�ٕ�yJb�"�2�̼��ɢ�Pb%�%%����w�m�y)V
� R��b\E��"��ф�f��-��;y�$�uTr���Z�)ʺ$<��{I}hv_�D$I��pR�1WwH-v�p9�	��Ȏ:ۗ����=ztL�f��8$��1�4��e4`h��0f:��^	I����)�D��Q���:4g�IsL�v>ُ�"�"�.��X)��t�v.�0�۲�#�z���M�>ݙ���vݟ��j�ʗ��8TF'����ð�i*�&�$AU�d7#B)7]d10���U�\Sn�Ҕ�C)�n�m'z�2b9vXf��^�x�����d�V�M�5J? ����l���t�i��3dA/D{�h�X�8�ԡj��%�"~.�P�XE�E�h���l���ҩ���������2�:�+a%5a$NV^��F��K�Bӭ+"a�͍�z�mT^1��5	��9z�i)�uP���ʽX&�z����Q;�J����F��X@�KtV �u]�����Vb�<wE��Y�5i�
֕�ǒ'2<�)�Otm��9�}9s�W���Ի�
��Ʊ�^��p�+r�p�C�ROa�ҫe�Rӷ
�C^V=B�;�M;��KM��EA�6�n�]L��) ��{�`��h<�jm�Sa\YsC:�'t"����n�U����J�5aX�j�[l:�u海eed�沮�.d�dU�����ɭ�Ѥ���Ev tNXoQ�K-�_<ױƅ���r;�/&��=��k����y��R!�@dWgF�rķ��H�:7�𤮥�Hqe^˄�$��w5m�3�)WM��x[&�W�°Rv��U�/]wĤf=a���ru/i�S&[���E�Sr)w�.�/s@̈F�h����B$2#�,XC9j�B�E�'U݌�,�[Ռ�Gp�.(+ ��GE]3��7�/kuXGq��v�еX�n�Mw2��&N��n�Wu�9��i�;�*$!�Ŗ�[ռ�m����M]�wk�3��S�+��*���-t�J��o/����)TT�4;���щL�9s�ɳ�nJ�k����9ł��u�V�sV{�:��%�!��\+���y�z�����$o���"���|�+�*"|���	��F^�fVT�Ɵcɡ�YYW�\w���
��{ûby}�U�f�^�P2�(��a��`f���-^�X�{��i�ʒ� ����D�`�pK*�-G�2���.�r]�Ll�{B�����+�����1�R��
o��T�x;xt�$�8/@Ħ����Xox ;^�f[x/-�Id�K���9��W8J�1EO%F�jK����u����^u���8�Ǯ��h�0+S�n]��g� ��F��>�U��Պ��� ��{�:�\;��3��ز�
N��]jR�g8�]���ݢ��vJ����qb��ٹku�˹�{MW5ZØ�/�P�X��S���ed �壨�w`>�.�I��J5u�ۏl�z��d����-��w�גw:	CF.΃e�Zs�".t2^�t������u\,��oFPƕ��H�1V@X��^�ږ t�÷�q.�����,c�]]6�j�ԯ�2m�i�G�۬�}�j�ث.V}��f�B딾9	�w��ݐ���7��Qw� us��͙1Ӊ��E��&��S2�i�;2��.Xe��1�v,�ƶQ�0ù#��9�h�V�Xk�c�Z��X0��Gy�f>�{������B�S�1
�v�<Y���K�Ʉu&I/.��xi�G�W��Z�����J��/yB�!�掚�Q23�w�X 
;�V/8�&t�z]0�%*�,�k��U���+x��^�t�|Uu�|�R�G��C��M��w�Q�ސmР�h�}�t\���d��Ph���\t�V4V!����aq��6sz��I"XE콱|�s��.�rf��c��DԻw�wj�7h��X�(04rQJ���nq���ߵ���޼m�O0���cɣ#���ʾ��[�AA[v�4k$�8Gov�i����M7M˽�;{mSMї%֪�沯9Kkd�J,�G�YC�ֱX0̾�9a7q=�`�-���O����m��μ_(��5u:t����p���
���e�nd�F4�pD�R�.����E�ʗN����
ޠQ�9/�Y��:*�Cm�e9iqX`��:n�G��a��n��"Δ7w��)"�ݫ�Ja��9rgZ�������ͫ���0���t]F;�du�+���]B����[>o�����V*�WI�Wڴ�ҰV>�u�ܥ]d�W;p�m.�|�;�Ϟ9��i��]Ҹ`�����p�,�������
�f�E�h�͒��(��zl����)�ɂnxn4�Y;�^+�)���)ʽ/z��(��f%� �v�>ޜ!�e���k�1Ve�.�}��^<�5R�2�B�#��ս�r����6�92,��{wb��j��m����w�J��#](N�|(� yt,�q�D}z6Z�=I���f��Ju8�-7��x���T�T���1jh/�r�|�u'hg-�����9�[R�u	重0T.�ê�-=nm�en�D�p�����E"�58����out��<����h�$�H2�-(�3@O� /�;oiP6�I�����"k��_e������[�}��"�f�[�휍nf�u,E4t9��0���ݵ��fR�P�*��X��IpK�n�uMC�u�;���ڀ���N�����Xk��>��xz��Zvmۇ���P��L�})��(S�XѼEN.��\�Ɇ,���*�f���J׳K�s�h���x����@�0-��ut7"���=V�u�^*�P޵��%.ۄ�3Cڻp�	�^�[[]b@�/���5�*��9e��{�Ȅ軔zJ�t^��l�RC�J��w����] z���OX��
�lՌ����@v��[ee�����+6�.-|���T �JT���բ�Uu1
'#R�\ioC�Z��`���6o�%gT��w_
B�<�w���$4�me���ʆo��o�ε9n�SQ���R��R_[33�q������X�w�ܳ'e���;�7XŰ4\s��T/�n�N-����pE55�kNm{�����q���q�=;�rK�MeMQ�Av0)�+��]�����e���SM�������G�G:�˜SW��]Ѕ�|ZO,�JIU�B�����Lr�)�0˫[.�0f�iJWYA��&���� ��ژ��N�Y���p��eM�R����%'n�K}�hb���h�v�q+��fS{V �Y�9D����o�v�`k'bPc��ڳ�6��Z%��ք�:Yֱ��WNh�ۛ����{���[��\��4C	�^��8�jd�Z�z��1�}�hfub��+�Kl7� �6TY�ዞG�]�F�8۵]��]+��	*���v�G ��꒺�_}��j�O�`n»��]b����Y�p��'lt-���:���@�����9��WEX�=M�%�,�4E�t.��TG��*��iqZ䶬�>�{J��[�6B�o�@���X1jήqq��;�ڷr�m*���؍�Nq�m��*օk�t��j930�X6e��4W|�ʉJ\��8��1-���_ޢ����7�k��ɛ�#��u5�+X:�mȞa�+�}h��r���ol�� ��=+ �zkV2��p�G�R�y����FպU,�c"��pjX:IX�4��[���{:�B�顉H�p�gVHk�ø��kkD��9�\�S��&)<��t-XJS}q���Y�6�*�9�JO�OQ�\jq�zv�X�0�"�����9b/HT����n�H�.x^�;t5`7��#8gU��F��`݇Q�L�����Rږ�[b�_4�4����o��4��t �"b�X}�c������B��O��6�_=��̳���2�˙kT�=��{w��S��w`L��\� ��_'��V*Z�;�ev.�)],juD;;4K
Ef�{����FPv՗�@u:c57�T�]^<6�4��-�4��|7��D��9��P֤����ۥ�)�3����؏��i+�%@ �x��f��Hmt��^)L�T6��#�9]�2˰�}�w4{V�.����O���F��XU/Q�(�{�t�uj!��%����/�
��/Ly{۷�)N��Bi�d�]\Y�5�t���Ӿ���B+ >���.��l��㓙qzh�"�_'u�Ɵ{eƩg
(�8����z�Lnjm��U�ز�֭utXL<��:v����!l��ݫ̄%q\`�l�ӂ�ηU��/f�� A^�q�S-��M�iW�S��+�__hr)Z	�\R�m���3�̳a��ܣZ��Sx=��J�lw&���@�.r��"�(V��5;j`b�bݸ���˵c�' ���r���pEi9������%Kc��K H	��L�2����]}�w�1����,Ry��ر[�Vn��T3Y�q���mΠ�:���ՙc�V�_.|���
�.|�g1�)HL����8�.�
In�4��|l��k22m݃Y�5AtbenP�"`�as��4Vt��@ڰC/5���A/7�]7�]�͂��5�]m\o��W+\>O��A�p-&�D��U�����3B��.:�73��>��Z���et�N�cQ,�f#Ù��:�w�O�䎺��
s�XH�ǖ��f�޷�yK�^����t����VY����I������gZ6�'�f�i����Wp�8����mEH�sd\��:�]nT��K�)����y�W�����j���ٱ��������w�d�U����}��^���۴��Pb[NWEO%e%Y3��5���^P��kF�c���o���tU�>�{m����v6b����4Q�R �8h�n�VTٯ�7s������㶁�H�n8�ͻ]\ժ-�RK̗pԇ�*̆��wS�7��,�B�\/���i���&<���;���;kC]��hiDm�d���79S
��M��W!��d_,҈�M�t�2"o��X���$�ѩџ)�WL��@v��dԾz�SX6Tz�E��TP��"��@ufp����ַM��OK���R�������d����t�D�ݼ�j�qط��$�t�Ŧ�V�롍ԶNP��w%NDcvxK8r#���R�GF��O���F�Ǚ��3l�W��eӸ0����;_��O��(H�S�Cs\��(o+��j�o/h��ܸ��ފ�Bn�xֻr�ݠ�l$�mw^ee0�9Z2�qg) л�J<�R�{q\Ķ�u����݀�qޔ_w[�{���tCf�ظ��(��@�;Q���,%�\�Vu�;�e9�������U��*҉	tpe֓
�X۹�b���K���79��8Jj:SH�"����rG�Gg%��t&��2��9ɕ������]�������-kc��-��ʌ�JT:�y��GB��;2��7I�'��L���JQbU��o	�'$g���Y��.E�
|#r�gZ� �9+T��ۘ�"��򘾑�"��$J�Ւ*�QfD ���1b�K&�dM�p˜ml(�[�VWeB��JCmt���Zf��{"����n�^�j���.�+K�wz`�]���Cy���+㲬!0��g�egSЉ)!�+"v>�e�%uY!�J���'U0e�;�5�`��Q�o7��a�y����F���a=�NB�fl��;���D��46"�^�WS��F�m=w\�AS��_��ތ�]`�xJ�N��Oɯy_Kc$G�kg��qک�o;f�N�+�]tpC&_1j���r�sb��R�G��ۙ�e�Uq=̇O,3{�ZHrA#(��WPY�i ���I�u�t-�\�L�|(e��n�]�2$�^�+�N�'�G�i�Wl�O�"�6��w�h����W�[�t(2�v؊i��z�H8������EZA�|��U���=�M���y$yݘ���B���&��{�n��]�1���M9{��lx�@������FegLَ�KȆv�w�+j�l�����0��b���/U��5de>�Q�u�W��-|V�`i�`�#�{�nP�����t��v�P�e������}�}�ūs�:�ך�0��+/�*m��_+�'fS�tk=��eEK-��N�*��d�ykr0/r����A�QXiK�Hk�a�� um^��OF�7�>E�}�,݅ӝ�iL��L�Xr_ٺ���d�@o�5
N5}j�T�LQ�!B�U��e��F�_ni�[WŭqQZ��@\��^r�8)�쁐����K����f�a1�����c�_	��i�祛-	�֧������c1�>[��&�)Di�g4�3�{L�a*}@5Nʙ��ۮ\1���[4�T0�rY�ڈnhѱ�F6�9�t%uz;�.�ױ�=d]�8���Q,2��O;�:�P5z��T2kW�@�-�k3Z��5�c�Vq��.�����E��������0��}y��]��l$[N��T�G������AA�Gݰ���W�͞ݲ����k�5��*�bz�}3����/Mk�l�#yT�z�_t�4b�8�m�69f�7�u�r�:���a��i���kHef^�"uq��H`}E6+i�o5ԩ�/�4�^�n���$����ݹЕ��832�����H�is�٭��E��C��,���-:�!��߳.1 L�]aY�3^J9�b�O+��vs��:�Quo��e�J���eɀ7��i�5m���0�|�W����GkK`>�\��Yۿ�/�V�oa��n���V�W[#�j� �߯�wWG�WN7wH^�:L�^�Řw-.�[h��r�e���w
��[\��.qopD;��w�	,�vf�T�e9;��lTXY�� -oc���XNT�8Ҙ&�⡏��݉�����i]�����U�&i�N<ok��-,��ݰL�����:c��F��˝u�pTSI�n�:m�ES�z��+�<!��᪁ҕ�0��4S��N�ǒ����װZ�cG��0{Flc�ߴَ��*��n>�B�<��XY�׃��͕�tx��"�妰�Ĝ�u��&ŉǛ��
��	5�ˡ+ ��ޖ���غ	�����/��ѭyxx�AcH
ɢ����R:]˘6�-W�Os(!���Z�iF��;YNヹ㙺�N�g���兒��4�h����iWW>NWQB�ݺṪ�-�AX
���-���[�rȻ�2	E�%p=��~�X����n��k�
��n�k�tm�Ȩwoq �O�[dc��c_ml�����sо��Ho$�fa�&1Q�J���j���мJ�l�[���*�q��p�w���WJn]��iK޸���.3�����oK�ܬU$���(�:C�}�����c5����hf˭�ݓY��]AlG������L�B�T2�T����gU��*��yS|#W@��N�%�N��:�N#��a��ٴ'�%�wS
(�C���"��'��Em̮��֦���m���J��$bH���b�b��+����*7JY����,��Nw,|n�S��A!U������s�)ݥ�T�������w[��� ���.�F��G�5_	��i�W�ݽ���T�wR��30�Q��#�+o�-�޺�ϸ���+r��h��U3�AK�L���9���R���BND<��*�J��}֊�]�oe��x'wE��hkowN��Bj0!�u{׽,|{2�EY��d3��]�lt�#�Y`m�m:ξ�b�}X�x
0��:�M�WN_�������꯺� C��	!	'�����_�������]��V�3�;�˚qC\7k�a�O^t��d��H��iX��f�Oj��>�H�1�w�^��]�R���@�L�F�t��sA >�P;�X��D��o��`з�!@�o5/ul�7N�uB�ݤ��,�0嚹����F�L}�=�ƁGGc��u�p&�Wl��V��)s,���M�>�����jdX�ظ"R����e�z;�9׻�c;H��"���C��j+SG��� ��,�Z�M��$'jy]���z����+yk�����	�kt�:V/f��U�݇1��Tz,�o��A4[���t����I�q{�o�fL�:xi՛X�P�5�:١��I՝r�+r��-Yt:��!�3��o��9�{9�z��t)�T{<������p�]#1}�;jK��ܝ��(i��y?���q��1�_*�K�2�`<9�j��`�T�w�
x��nc@V]3/^��E�X3jԮkJ�VC
����f���}��(�t������F��� )�ٷ6�Í!�@d,*V�֩���S��B�](`剃d�R]���oDΗXn /e
�SF�훽|��k�$d����"�;3��p)���]�]�n�0�G�rf�Y��P>!\׆�n��9G���2���d���h�MZ�֣V��;���^C����&�A_S��r�ܳk$1е��&�u^���8�0/V� �R}y}ۥ�JM�/��8S�J,�2��oy�_V]�[�	]��Q^^��[ڇd��Bͥ%���: ���,/��*eDeZz�Q�H�E���V��qΨ�fv�bCy(p��];kTyӠ{ۗAQ]5�2� �u�ܲrS��n��}{A�	���\�v���m�s(P����J��c%��Χ ��%�nu�44�VOº|gV�<fXu�7hR�zc���$(䷦�9Wc�yXN��ܱ,�d��>K+�6ƕx���6�!lx���(�\-�o�nT�Ѯ��ᢋ��B3h�Qu0^bFH(S����Ss���>6{2�-^P�d#�*U��d���;�.��k�k��Ǌ��U^<�m�� �<��B��末�J�8溎�5k &��/�Mʫm��`1s;��!Rv$�(����c�b]��V=�Q_e��|퍑��/n�u�`�R��۶����u����ڝЂc�]����#�hs���&@X��[�b�'f���݁ �m6 ��l>j;�rr�аѵN����!u�`�t�*Hxf����w{���1�f�@o�i�e��l٧�w�IORӥg/��m�����g�[���V��[)b����5ڥ��᫉]���\\mb�W>n��+��r�`gC���Ckf���B�"��AjQd릛��sesJؠzc�)5[`t7G�Ϟ��镥���T�ˮt;HV�CV��`χ�ӌ��]-�h�F��I�D����fm�e�OC�q��PIw�.�h�Y��XKiE3Ey�21�eh��cY0�FA�+A���ŷ��C�ݱ��yG�{:�<R����u!�ޛV+Bo 9[�ao#r�u}`�1���#si�J�gtݼ���n^)�3:���7��W5yoK�b�ғ���3Cͫ�-@��%��K��U�o��y�G�T.�r�U�K1����H�ηk��CZڶ�b�m!�i��n_A2$p��W%7���c�Y��+�\͓Q�Q �W�p��nT���s����3h�cjp�x���T���s�]���.�d�Py�aΗL�3�����F�f;Qd�1��uZ}��]J9�i�T��fCd=����!�(��ѽ�*#�g�!7AEyH�:��YJ7^۩ܢz�E�]w�pxFm�[(6Rr�z@u��-^�Ȟb�&qv�wV�l�r5��i���<FDR�O���<����lݽER����{�v+蛣������!6��XR�k�Ӕr�$��>��Hˡod�й=��|�)ue��Z��ɷZΛ&�����[$r�e�]��YZ+e��~(��%���J�d��5�[{�����p�Ab��sQ�myg^@���H�e�ݒ�BP��+�������\�.7L=��IW6���	q��/�&��ee���B�_�/�Vq)WJ�$�:7�M���tI�bƍS�r�v�B�i�2�M���6�������k����! ��,V�Ɯ�[h`b_r�V^�5r���pݕrQU6�MSjfT��M.��1v��zN�a��ˬ�ė����2�e�*�Vt�����wW �x���w[�G�R3�r���G/��0.�1�$�m��f'�	Z�I�M<����E��N<.q�tџBqY�}$++�vwp���pe��ɛ����3��z���ºn��ݛ��N.��OfN\ˎ�Z�k�+u�=��;�w��ˇ��I�of��Fћ�,��A���n�Շ �cZ�
�P��]�:Y^���er�m-WƗ[M4�-o5{| ��v��Y�Z��i�ŭ+�nn��Rf���;d��W���S롛���/z�.��U����M���s��V�*VS}��1n�.$f��5�Xt֛�&��Kf�M��EW�du&�:`���ڼ��:�C�F���V-,=ƶ���Qͽk�&�sU�7b�M��ugN���:_a�.��Z����n��y=��Ɏ0����Q���D<,�Z��Ab�;|cS

[ġ*�u��F�m5�JkUt����ҳN�//9=�z���!u�g�q]��8PS}��ʛ�r�vZIk���I���n�v�˕�;]�˻�F�&��w[Y�U�a�ݧ�%.s�XA�-��W�\�cH��FR8T��#^)�4T:��ʵ�It��&�rOl[ߌ���_j�qje��<�ݥ���*#z�sܒp�UM����n������v���x��D'6i��j�MEi������*��]������s�I!y���D�X�X3[qC� {��R�b��>Z��;�Q����_-㔪:�`�-q�Y�C:��Xx&J�����>t;E��O*�n+���R6��td#q=z�'�+&�u���+�=�j=S��6�B{�Ш�
�%p]�2�7`^y���u���T�%[7�ؚ�ܦ��U����Պк�5u�(wl���z�(�3%\�>I�����w�^�t����&��Y��V�,&�xt�},D�g<�#�P��GSP�*A�/�f��U��f�pqX�P�`�镺6��n^Q-��U��x�}��g���I:�@n[���ߴE��]r�WK�b�h�¡��Cں���I|(��۵���&����̺]�RʓkZ)�Ѣ=��{H���j]JEx65��CO1�R����A�§kw�;�c`�!��b����&M���ᩒ��f��n��������r٣V]`����>)����#���=S,�=+.*�/h10���0�iu�-]j�]�,ګq�kEf�����=�3�v͇[����	P7���#��ʆ���f���nl�9)��Y�U�t_#�.l�dV�2��`���_
��']����T���/�
�n� [�,��J�����oZ���������Y��֑�M��;)��2+9�/q�@˭�1���NgAۍ��fIWD���w\��s:��^��������|]%^��]�i�=���jX��ۼ��:̾a]��uxA�Х0�X1շ���H��,r͑|���2I��&�n.��2�Ùc�ju8��M�
��B,���,_lu����k^���RYXu]�(-��0�M�G�@ 8Z-0��� [��p+�C䪃6i%��lN����z���ۈ'M��w��4&m�ngB�-��5�;y�r��;�41���^ڏSkyX�ۼ�����jLF��ut]�mk�ښ��>ٺW�r+��*��]�G]f�hj�qJ�"es�Ö
����,�M��BRI�k�ثb�P����v�Bk��%mm���%VqQÂt]���z2�ŶD{��p�TWL�����I�u�f��8�#�7���G��f�>Q��.����o�M��E�YY�9�}hlV���c]7B>����@m��%n�6k���WLp�"�7�JT�2vk�}�;I���7t��Y̅��y��u��,�x8f0�[�p	�㙆��.�Klv�>,ʷK㚣���Gc��*=y9���7�vk������d��櫆˝;jL��`�k���Z*r�%�#)����vou�k]5�������e�w�'N�\|�y�Gi��K
Q�o��cn�J޳ŭR�-��Hm/S�(q&|z�-M,�a���S&т�Wfo�A����#�f�
����u��nQ�|��Db�Z��� Fe���
A�Ӽ���ҵj��lV�t[�f�]1��cZv@�u]�WOzO��7Y-��2��`뒷vb] |��4h1�[{�wg	�]�i⥋i��=G��@�7u^�z�n�����I��mv��Is,X`<�n�r�n9x1J"�]%K.st�]�wM&���ܬ]�X���-�{K(��kpf�%��3���%n�	��;�s%��u��Us��6n�:H���nc/�1���P�)�ՙ4���uN�m�.���t2v�v�_̆��;켾MZt�dB-
�=��r�d� Y����M����}ݧ��&g!�9�&��f�Ff���V1t�����V>CP�*�2�
���S�Q�tQ����[P �OX�ئ��X��b�'es�ufjv�\3o����1Tk�#+j���dO���K�Zqs&�I|GFEY�d�on��4@�j�9���Q�yu(��.�v�ݣֻ(��oUb��KvP7��!�\�/�0�sxF��8k2h<�rL��/����K�=�}٥tz�ԠB�˲E���4:�um��v��m=$|�2��=���@�E7Z���d�Ӵ5V[��"�\�֨_v���M�ul�c�bm�;;z��r�]G^�\9G�vr���:MB�+ɻ|��z�m�I[޲d�1�e���f��t�x�ثy��
�J't�L�ǻ���\Vt����E`�u�BķP��M��W \؇$���g�S�h������j�W+8xL�"�j��R���벋���w��൏운�v]�lF�e�}�c����k�ٵ�^gL[b2I��L��jQ s��:��A$t�Y���hk��U�׵&�b�v����k:�	�|�^�~\�]&�<���*$3m��f�utI�9uD|5�eV�-�`u�]tI��C2�YE��C���+6�� ���& &�A�ɛ�NR���m5F�C��#6���\��KkaYY�۬9ɛlb̠��ܝ�W
Es~����C���Ӗ��F�M�j��|+ �.�]�������mi	L���������N
SS�9+)V��s�3 �w\ݕMuȔ˔5*�:��gO�����&����Vj��[u%��L��b Ww��c3
�<gL��M���$�P݇�@�V,��:"	��gm�[[�:�)�Ji�B�u�ZK���=�N���&��.��A,x�L�������J��)Ib��,/�R��WY�_ gfn;�a|�[תkM@LY�����SE1PPM�y�y����m7��.ٹܻ���*{7��a�!�0���V�G[��jm7+K�E`\a�sz��L!�$��i�,��S�u{��d�O
����)D���u����]Ac����,��Q
T�hU��[A��vҐ\��Ȥ���tf����u���X��L�Y˒�q��8vj��Cx��Ӭ�JfL�C��-aį�GX�k~8��.�#����(){x�#��X5��Ǳ|tm�2[�y��;JC�El��X㝎-\��gU�8�`aS�83���L=%����N��NGa�,���!��h�|&���҂��,p�1r�c�\�����Iu���o���1*ٖ�^��w]p	jjh�!. U��L�YW�k��zq��`5��7��w��*^�W�n5��ˊ&0�cx����ZS�=ܦ��J
�^kR]�Θ�:A=�]��X�8p��N,u�43�0�v�f���H�ջ_v�i��}�JWfXgc�gwSn��W6��Pe��V) �5���}k���$���\s�ɝk(�B�i.��w;�Һ�R_b�Ct���]Ԯj59�v���j#�бX=�f���v�lu��G��\P p@�?b{����8��y���Rz���P&*�Yұ����Һ�;X�_i1� w�<ا�uVs�b�;�[m��� �Y�y�؁�j�\������K��'t��H&�}P *��e*wV�����jm�k�Z̉T���׻au<DI���W�n�X	Zv�6�
]Y�{�s��j!Bʶ*�!�Y|�.�����ҽ��Y;��/�n=`�K[Ԯ�7�t�40�E7@�wj8�;��_2�;(�꺺o���z�L��"P+���Onm���RN���Z����P�@�J��ϻ��%1Ɠ�g3^�Zd�8UNQ���c�X��Ź)�Wt].�z]U�W���ϊ�q�v�[�f0����b�%gX�FK��ᗰhV;R�ċ)=x�a�WthS7#p8gc����¶�}���{]���t�Vc��]j�pT��`�-�ʠ��Z��P��^Ѵ����=)�7�w��˽绩��wV��V�kˣk�X;���h�ի�Jūi�q�-4":4u��c�n�`z�l�ft{ܷ{;E>���t3H&cuo���TA9.�4�I���
�7z]���`HL?1.��(#������v����M
������ݧ%��o��o��t�3a�S�;�:U���6�U�=��z�u�v��q�n 8ԡ`�e��JI�/h	��O���_}�}_}���i]��Z+������݋`�6SL���2��P�6�?Z�	�M��i<<�텰��U���M�@ug]��]#JD\�����X��{{*2 �=V`���q����`j ���x�	DU��7r;p�ܹ�u���`�u"p���(���`��g�yc�׼SHG]��=��ƺ����1�e�S��H�Ƞ��=w�x��G\ۈd��^Ҙ�,^�yԒ�^	��\�Z�GsP5-ⲱ)��_] ��ݣ������-�Sq�m��KI����K��5J��aA���9}�о�
�� ��L[�Ƕrr��w��5,���o���uґU�ve��I�[�U�O�aJ������]^dK޼u�B��t�5��֒�@�
5��4���d0m��+�m���Ӱ�!��J��mu�{;�jM�j$BЬKO��;������ ��} hu���R��6�3]r_d;cVǆ�$.�9H5ֶ�48ޒ��s٢�g������a7��}��'h�R�+/e�mf��n'WN�-�V�e�G�Mos���=���jj��9�7;�;���:Tr>t*V�t�)�W9�+*�^�E��ͫJfqM|K�:%nU�[]IGv4
����R��Y�C��HXT��p�'Cz��;[��m ���Fq)���uN�����V+��@R(�+%dY*T�L�~C��+ԷY�E��R�T�XV�F�B��qY.��� F���Vq�ER�m���U�D�b�E��űb����faG2:��B)�$Ԡ�V�PY3%f�Zͨ�fA
 �'��R
EXfJ*H��(,�!�Y�
)���H���%J�"�B,�TR]I�D��×��/,��5EQ0��eTyg����QXj
�P.�L�2
,��U��Lʨr�8� d��f-�PFr���PX��q2f�XreHT�.���2C$ͶEZ�ET�B�x�y��*¡mF�P���ڤXJ�UdXaU�Z2<����h"�����K������Q_p����6cWk�i��o^�n�.�
��%��D����:����5��3�Ws�,�P��ժEI�/�U���J��Ŷ�[��bZ��+�#yR�>�����yUb� ��P`���}�ނ-�z���ր+�_�����v�x�����1�.�mAw]A��Y�2ou^��4|\j�7)�_q`�ȩ[���C8���'ޖ�
t����2¯xo���i�G��3�g����f
��lNC� �f�q
��Y�2��.�F��{Z{6y�m>!i�f��?S�ab2Բ������G�^[D��[��FL��ZV�[��˄9�����(	��D
�|���A�~Xk�߯�~~��Me&~�=Թ������q}>X���傽.=� _��� ��r}������*��{���<�_?x��,)>��ϝ��い��퉊��v��k������n�<�8���n��޹�~���p�ҙcB򓦟�hC"	�`�ǉ�{��j����h����{#��Bg�Nr}nU_�ӧG���/\�Y0�"���y����`>3��f�`?��aDk���)[Yv,!{��û[oV��I�0^0�t��o�����{���/f//�+���,<]R���S��c�#gx{�6孶z>9�,%�2wP�޹[�C��jK����wg7���w�Y]�7(�e�ݝ��[<��V:���k��9ǫ��9~�eK���U�,Pm���r��5j~�k*�p\�{a���7H���Ί�
r�Ohs7~�9Հk|T��q�P��2�{_�9{Nd ���1�U�>�3;���R�aX���%t;.�F0�`FkAؼ;e������3��Z<'���l���gA~Jt���=�7����+edLx��Ugb~���=�`ܭ�c���*�J�ż>�m��b���I_�q�Z�u��U���REF�P�LL!�1�Sw�2 {>�Y��;Z2���m��v�ԥ/���2�rr%�M�"�UD�Q� -#ɽ�@��|q�~9u,r9=�������Ja�'��u�ϕB~�Ke�w�7@SYNH
A�O��f#��k`���a��=שҷ����\)߬�P߶C�����Tl��o"T-x���Y��F\86!�����TN#�>S��l]��V�p���MW�ǅ�6���%�7T!���[W#���V��Eo}�]z/_�	���y���F��w�X�����ԫ�W=�{�l����]'[ǲ�J"�A}ԯ(�ay7��LE��Ͳ���.�Ɲr!�Hؗm7ϴ=���(#Ut#��v�.!ދ����S�V���3D[��Ӄ����@�Uή'C��� ;X��ͼu�Z��s�3&��\�����k����wT%�x�θ�Sw��p6�mze��#q�>��y�_��*�x��b�xo�uZ�&Mg�0�k��^���z��W�Y��h���;Y���9��+%y�#��*�,�Vv�8�h�q�3�+^�(I�~̨{p'ek���7ٓ��t�+��EΧ�⾭�L�ߩO��3TeTh!Ù�8KҔlȏW�L}_y	BB9؉ݨ��'�:~~�G�aS~Z�Tv��g09/�w�[������p�bc��;��}����^v�x���b��0�s���ij�����>�5U٫�B߽p	UqoV�
�)�~ƴi�~��41G�b��=�ԋ!�Ȫ��x��:�^�J־�s�PqN�R�Ww){o��0M�f,����u:ՊW�l������j���B�e�`47�J�lS9��AO��X��[帒�I�y�47k�fyצ���b�V��1�]����i�^�`�(���p���L���t4�o�3N�����zRX�T���T������+́���;Np�4mo��p��cѧ2[�#)l�2⬹�\3f�^Vp�4+*����1P��n� Z�+8�"з��	/�j�J̈́#r9N-47��S������i\7O�n;��}�澬u䡝��	���7U�[��D����ظP�l��/F�ң+B)��0E����nP��J!�c7&������"��Tɯ�\��;~����|����y!Z�5�^y�'�"�lp�,�|,?���1_����lL�w2�ɭ��92�|F�'nh�>��
��+�>;��a��Ķ�S{��+��w����^>�y��3δ!��Fo}�ϋ�(SuLM�ڱQ��7�#��2c��麰�윯M���d����K%E�)c�JrC�~��d��ŵ�&.˞��m�W[�yi����V%P�n��'�_�
�O[>�AXۛ{kP�	�ӑ�:
f#�0������W��m
�d?�����'k�|��r�/{����ש=(KdV[�2���?_�H?#A��^��`���{
?O$�l5�ٙ}^ƁZ|���t�^t!��d����
�X��r��U����<G��m���=�us�:1����u�7�@\���N�9�*��r��F�q/�S3���m�]l�O��~����O����+�;ق�}���^�����v�X�De��7�!''+�J�$����b���0;9�7ݜ[�y_��:����Tp���V���u�^�qK9N2��F�_v+:�_pa{�X=�w=��L��۞Y��z]3	�E�ǀ���y܏h���Ț��G4V)o�j��䈜Swˊ��Vڃ���zwZ��c���ߪ�@ә^��2�J�v�|w*Q܏*(T<�`-�#=�g\�7����M�k�'_���r��)�pb�u��L^���>���r�:ּ�4{Ob�g��ڲ �6���ͧ���8�y���|pdu�H��z�T+�;�L�u��~;ƫ{���7L�u�Ӻ�u	W�\�z�b�����誙,`�.V ��M]�<<�dC�
χ��{�}wފ<{����&1��E"�Db�T��w)�F{V:5ru��Mx]���,�^�m=<(�-�;4%ߚ[R������P�5tZ�r�+���������~�W�eV{��LeE�q�?f:�������P䶦��5��@EF� 'R��F�~�dyuo�m�¸G.}c���2o��,���fgE�j�}1�1?'Y��L<���#Y���4M����Q�mM�Ln)ϹM{ϥ�C�{��\�c5o]�6|��51R˛fB������4�ˎ���$m�+[��z��u��,LKV����� ��> g������}��Ql�Y�öE����\�CE��<�Ľس���pC�|5u.s��<��tbx���1F�[�	A��h������`����טR�֍�6*���n�lw�ͺ�I�\U��76��_.=�8��{�6�n'����3R�i;�>�{��/�O�@�Є����傽*��`���c����6��>����7yzʧa�6��8|��o�+}���^x0�~@[�O��p(���ʠ���������J�L i�!��P�׹GM�z�BV,��I`_u�YV����?�y�I�T��d-���د��;F�z��Ơ���a ���υZ݀#�q�ߞ���Y�z�f�����*_G�w<B���Cr���_zل#��qN�@��+gQ�J[-��b)ݳ��.�O�� �5�*�q��=�V����>Ӟ"�yyW�z�f�d��������Hv�b|�������Bv���ݚG*X�9��*����a�V�������+y�\�a�o��~�w��cԃ���J��U�k+�L\��˱d����	���"\p�{��y���)x^�����u$J.��.!He�ɡP��-ތV�6,0���'����}��V}�3e׋�u�AɍJeI�T����d
��� -TiG�5u�s�۝�S��m��9KT���;���鋁sϻ�E5��n�껎Y��o�rN��)^Φ�<�r'c��mE�]��z����}x���72\���Gt��&��Nf ;$�ŧ���a�_��'^9��Z�'5i�O8_>h_<Ǜ:��{;tr��u%Y��u$;����_��B��L����t�<g(
[.H��/c)A�	�v����n̆��X�U����c���Z�<��]�8�jU����t�ڵٚ��&{���F /�}��"��~F���x��Ƽ���L ���}�%_.a��}�-K�4�\�{F�Cx+�To�<;y�����y����K)^��x<?=�ʼ��� �M{eC��}8�*��W����@��B��^H��k��Z^�k��k�T�R�	&���:��q�Z��l	p�@`B��/���>>�X=��yz��@ާeX�ͥ΢�F|:x˭��*��U�����V��g�U�����{ٓ�U�t��J���b;f�ۤ�P�BisDD�i��V�3�0C&i�Z[��Z��u���[(O�n[�9/Lz�����%�[��pߞ!u4<�.�X��0�OI`:�ϰ�*Ү%�}u��4�
{i��ȣNFy����[��^�X�.$�1����*���ɯ렟�p	qoip����e}K_�z�K�r��w]2�[dp�f�W� *~�^)Γ;}QE��Zl���-5��[��.���1���n*_t�Od��z,Z�t�f�].7��Z�:}�xq�i�"ѵܦs�Z���<��a��##�V�˺b,�;�@�_V�7[���r�ٽ�8��1E�')Afs]�٣�*CE�:ypFєV� %5e �l��Ί�/���Ww*�<�kX#7�������Ý��@B5�pTE��`;���������4�]�b�=<�(7�h�J3�b�y瓻)6��c�@k�`���x��\!���4k�ڥ��_�8�IS�u���̢| �O/��~�V+��fD=-T�W?W�U��J/��ÒR�)���W��]�#�}��VZ@A	�T����2�.��}�E����5y~��=���y�����?n��D{�A����(��=�^s	�Ԋѱ¼����X\+|i�DʿrOG?M�Y��[��Q�c� yx!O�h����O2W^c�.�X��WxEF��w�qyz��x=��ڎ����h��x�U���
�����ت��g�:o��^o��um_��s�ydt����17+n@8��aL�n�xQ����mߪ����zz�\�ٹ~��h�]��p��Y�]O{�{-�4���_a��>�}�^�ݨ5� ]��e�S&���/[#�'k������.�'�1�p�H�;��a����<C��7@Ь����-<�3�!�q���`�Df]>���ɩσnh�A��vm�����=U8��[x9>��R��SG�]���RX�\��y�:/�L:�@_b#ך� �M�"��_ɫ�ց�$(�W����ETo��]��+�'�,n����po����ʿ +�ؐ�y��������DsN�j�w����'�{���q����W�6��M��vyϩ};�R�����xOU3:봌�o9i�[9}�4p�������+���^ ?��o+f ��U8^��"���_��du��IN��0��e��am굆�a��l�ˮ���9�L?-`vkh[3z��Y�����ܡ�70�VZ;f(7Q��Lj�~*<P�
���8�rP�˨�����I!yܓ�+��㴖I ��m�>^�}Fs����g׏�f���,:��/�7�U��`voy?D[�K��A�h��H�	K����j���X���=�ѐ,۵�"������@o�n�����J�>�����r�F�I�n͓^sૅ*��< �۵�|�͸����]"�K���:[��:@iB�k�y}�9�=��eUg��N9���;q��W�9+ɘt*;��կ��:W>�R���6P�j�{}�ʿY!���&s6p��A]�pw�Β����q�C0%Qp*�f��S�˾�C���Y�\�ǚ{��`�p46�(u��
����7k�nӨe�:��6D)'k$Y\9s7ە��j���*hçuue��E��gc鳮M����L��\��ܧ@ED#@0��g��m^[��x��������S���K�Xefp �D��p�If��0��g(
��`�5��Ƌ�����?i�q�Ԛr����D��C����EG����ǩ�1jD�^)e���qWY��
�nݩEJ��d��]a�B�[�y+D�ڼ<.�XV]_/
/ ������[����O����k�=��r���L�W�`�vZ�f;��E���yu�n  ?K FyH��n'}���E��3 �T{�Q�v�D/'�or��Y�v���.�k������h�tX���t������/��`h�
0�"��4\=�Z.!��BT�V"�*�iw5X���¥�{ҳ��ԝ�9�]��i��)XP������Y��^�i��n�3��#*�B�@n)Ү�z���ӳԑ`w-�=����ZU�����.V{�{����xꭚ�V眼�Gaf��u��d����˾~������[�Z�4�c�w�}����|XG�ny��#(3Mzؿ�G6�q^�G���V���f�)(j1�F�+��zJ=\�l//�8�5���E�O+r�@��]��]	�u��$�wu�9m.��q��D��V�.�z{i�Ö
{LΔ��	�kbo6<���Qk%�����F����sy�G�)D�N�X�mvX
����S&nhNB_�T��녋3U�j'q�������
Ar4:<W�Wr"�p��Uy�@�[��4��UD{h�l;
���N�$c=\eI���-��!L�ri=v��t��j�u�4
���-�8���ã�7�3s������7��$@�*�v����gn��E+����6����c����fS��*XXN�'ҳu�X�3]�wrޤ�՗
�˸���6�ScΘ{�+Ou4�&�S�7����y�ws�|�!V�X#�����R�4쇛V�������xk���#h}�J�����9Mx�J��d��C,R�Ţ����)qj��]:�9�E����z`ˇH-#�G}�^��@�Tj�t6�⊻�3 {ϊNU��s����E*��)s:SY���'G[,��_|5�Lx�s$��-鰫��/���C�+��M+��SW��,�0�-�,��W�32�s R�l�8;��PjS���zم�S��`�37zgm�|�k��΍K��S��0�`��6ur���u �I��ФH����Z.����^Xâ��ǆj��J��-��Q29Ou�1�ұӻr��F�gzZ�>d6$@h5�rƳ��f�О����}�SDP�P)��]�P��vf���/h��Ο^Gu�E���ެL�d�>�]���(W/�)���MM-݋�v�̃���n�`�]Gg�T�v�Ы�.mn[���֐���4�
��7���S'|�w��Ei-�����p��R]6��<��r�pr����-M1�x֕�eXUa[���V�4��[	�Y�B�<�[�F��!Jlu�y�xp��1E�1�[qj��h'#�{z8��p�rqآ�i�ƀ�����n��IdV�\����;5o��'v���q�.kU�la����W,�U���H�T�]�Iι\���z����l��:���A,VZd
��[�.��������݅
\i���{7��<�e�w;:}�1�WM���]$Q�.e����1:B�
�*��M��͉);�0d{|(c�b��1�vk%�&K�0��mҿܰ��
�\��qs��i�������qY�b�ґv<˼/GoG��ک�H��zY�uG}�����y�(����\�nem�_
7��o�0^��G �gu���B�ўÕ�<�gf�ŭjw\�1d��.�pwP�ytoH) �i��h�㫭���#��g+<M�G�bwq�e�g&{������5V�{MUbfw�R��7u��<��α$������^yYs�`�Py7�I�vl�퓴�������!�_oT�'\��ŕ���N�я�Rh��͝e�OI�Uׄ��E|X)m�B��Ņo,栫80MV�8���P��jf �*ʭ)`��k�X,y[BfVǖQ6���(+kl�L�@��X��
� ,�U[B�l�SR��G�//���X��9��Y��
�L֌AH��V�ڧ�a�qyv�-��Z���ĕF����ص�S[+�KK�5��Z�X�\ʬ�L�u��[q������Ԩ(���4��+m��*�AE.�!�g�a3u�*f��yN.��X�-��l�����m�Q�«Dex�d��D[���G��JթiZ21PyC0PUqJ���,�㕆kvÊ���kkU�������օ��dm
�UZ�eT��P5�QEmNm�+a�9+y��Tj�kɈT5iu�q3����N<UGRڈ-k*,m@R�!��nү#��.b\厘mKP=��\4���YΜ���Kk����*4� S���]�rc{��u�]���)��%'
���i'���:=�?���}N�|����>��s�<g�> T�|���T?0�7_0qԾX~C���Y�%@�*ts�=I���>�DF-^�E��ǛǞo0�DH�"��ʓ�v�NЬ����~`t�2Vt{�\����'v���ʁ��¬�����~�4=0+�|���C�v��T����Y�3�}C����>� ��|G��⚣QN�ɢ�B�Ի��>$(d�,���2{��ĝ�S?R{���g��_��ߜ��
ï79
��!Y���:C!�g�����'P�/�>w�"���^�P�}`����'�|��M��5���X�ğ��Ϻ���'ngGt�2t�U�I�d���}��S!�������%eg���'>%d���qY�T��9�*J���2u7��'I<N" �^�
=3�U�s��^�.�h�YY+���v�;d㕀�>b}C��>���ݲd=I^����Zt�Y���9퓧��Am�'��f}�֓��P�>�� T���t�YĉDߞ�$k���g����}���P�¡����W�;N�~i�Y�%@��;��W�q�'Ai<J�i/����a�z�{d��Nus!�K���'L3�� ��{d�Rx�I��N�,�@>�=�Y�l���k�ȝ}߿�s��P3���L�N t�~�kg�<g�����>$I�>n�C���_�t8��~�2�'}B�x�G,P<J���힐*OP����0㼰2�nt��|�M@����!�ZTm�����#G�w��tΙ*
����+gg����u�B�a�������ğS�~�� �ԟ\��i�AV|C�d��>�C>0��׈|>ސ<J�YS��g�����[Ǹ�p��DG���~�:Vx������t��+��M��J�v�:�����Y�%a�y֝�I�O�VO���p�&B�2}L�Ϻ�����������z�������8���z4��������+�1��j�� } G�>�?X�������:@�Y8Zx�t�P��y��Ԫ��*{��Hq�W�>��|�V}IY:��nӤ2J�O��{�S!�%���{֓��#�j�����jSF�߯�X$mM/JȎ�G��������Z{r;kpV�W�7��,
ޫc��) �;�����54	~�����w|Ux��␘��wzoes��XU�@�N��1϶U�����\��̛��5S�uԒ�-Sxr�_d��)��t+;.�}�u�s7��3]y3����a��|b2V#�^��%DH���L��Ѣ�}�xɒ�����*A|a���'Ă�~�|g�=N q+�^���Ϩx�!�翸S�Ad�>�ӈd��`u<��_XTz��"}�}��W�_;�������zJ�ĕ�<9�H,����$��V'��'G˒!������;��<aO��Ϩ~Hfu��}!�1����Ə���>��F�R&�Wr_���Ͻߞ�I�����N$�
�E��<L�����;J�Y��ι<~��J��8�!�Jà�x�x�'�;�N�����<M��2Ι+9>S�}N��O�H����}��~�|��wn7}s܀�D1X�#���mǙ����J���u�8�Y���
q����|�H"Oω�r����7=ǩ��*�����̟�w�Ğ!X~a~q:C��|}�ϿO�'���\�Ԗ{���x��C!"���v�߾c��P���=��D:I��?s�$�y�d<NͰVV><@����<d�Rx�~O�hH/l�}ǉ�q ��_(q��0�8���|������ޭ	����{��^�rרr�?xDh��$I�8�P��=g���̟;�>0�,��&�w� S�;B��z�2t��Vt��&@�?'���0�+�k��x��>��I�:d�)��߿�������F��P��}} >�"7�B����z����;O��8�Y�;x������ }J��:���d�2?������t|�N��ęĽ�y�qV}�v���~����L͌���R3k�#�>�F�s�IRv�:��@Y�3��~d��}�Ȥ�
�ßi�:~�+=I��N�S�����l��8�g����(
���?y�b���������jŋ�_{������{C�t�@�S��ZJ�Y����L� x�����*�S��;a�gV}�,<N!�J�O��l8��T;B��!Rz�{?S�Nu03+�L����ğ�p��t��|���Ӧ�/7U��G�|D1�eR��Z���Ak;�օzC�?&d�nn������Ͼ���� �_,>3�v�C0���>0�/��i��Rv����������/^�?y�u�j�θW��]f^E�C]�����]������^�CA�<sCn�&���x3B��f�w��E�㡲���2�ˑp��r��Ѭz�,�1�إoA��79���W<.vo-�H}D�����WyU1
¾�d���p�t����{ށ�VJ��vR�ÿ:��fz��`|mǦg��^&�Ӵ� �Ƕ�I�q3'��2�v�&B�ﯾ�`�3>5ȥK���t} H�4DH������Xv�������VJʬ�%��'Ht��+�w��t�ĕ�3�S��,���L3=L�2}s�]s���_��9������|���X)}�����3߅z��}vi���#�>����+�LA�ꎸ��@�>��|1�����e�^��3<������hOO+�Vu�gk����z��k� 뼪�ڬ����V�/gz-��� ���I����[��rp�Kn���.�vPӜ��yj�U��cC�+_ qc�[;<�w�C��Dk_���=�����/af,f�K1cK�t%s"��R�]�0/���7���N?E��ג��L���l��J��~�^Х7&,#�������l���,k:���d�3J�	�^p��M�C^�N��T���/�����0\b��ҫ�Mx �1�Q�j8s�:<�]�s^���R�Q�a�ҙ5]�c"�������l��M>W����.YY��{Y�'���pX>��EYH혠ު�1�j�zs��ۨw6��CU�cH��'�೓"B<>y8{�|xef��A�A��m=v�g���0�����YM����E&�����בxT5�lL=7��8Rq���a��4�V��
�3�:-�8J:�n�SOM�o��d�zt�
̮ȕ\yw)�S)J�A��wh[R���}6��X]�op�Mb�ڱ�Y>�عX��V���m�i=��ߠ�>�bf�TV=i^�µ��^az��x�?C���VX��_����}�1�/+B�i�����X�	K�+�+4.�I��է�ʧtx�1[⻂=e�jCR<�|�e=�K��^���u���0�v����o�^K�<�
�]Q��P���T�@���+�~L����˅����2��������e��@�sthֹY����F�T�3�tY�<����dE�="D���[�\�:0̿�P��Lb��,�;��R��
�5HRkH�xO-Ǘ�ϟ����q��%��o����Վ��N������UJr���c9�[dߖIӳ�ʚ+:��|�厼2��|�(��4� nz߀qW�U�X��ۄ�^���#޵_ee`[em���E�8�b�{z}q�3�����vܵ^��/]/+��I�^�x֜����
5��kG����ܴ0�g��S�ݧ��P���Z�Avc�%&��&���~���0��Vt�g
ڵ�{�,E��a��vOP�Ck,�ls�CD��-eé7y��iPV�z��G19�}��#��Qm��ч���m�Ң����W^^���E�v�ͦe5������t�q�n��Iu�Z`�}�nZ���v�E��*���n����*zaP��m�CE��:^宅��u�h�{ZeF9W%����݉D�����72,H����RɆ)�p�@gg�����Nv_�{������a*a�(��n�O=�%�����G�b��.׽��xy�g�j�B��&g_>�Ϝ��?_S�e��rP����G|Q¸��p5:o�O��?4���8vqE���<��E��-S�B!������.�쿾��w���h.����r_�R�e[P�׭y,ٜ�Җ���%��~R�j
��]��b�,�J���_���t)M{���R���-;_Xq碡�l�6��"��|+�����eu�K*���D/�L��^k��Y/VK�S��~��
��ʒ����Ȩ��Q V� ��si]�E��3=��ݵ�kQ{�8�??���e�<-�k����J���Q�_�6�j�1u��٬�����w݈��aV�
8:����V18X�u��ަOZ��>�h��G�Ejr^��x�����Lķ�ˬ�����K@��T�DA���]�o�`��r�!��kQϝ^Y����-qt��H�b,}�'Dk�u��aG0��]/���z��蒮p��;�F)���t�֎N)T�\'�����!ӳ�(��f�D�/�ˀ�3#>�%�܊��X�!��U�.���ʸx+��<O�W^t�n��Yܿ7d���%i"�W(�~�-�̝Y+�e{�,̟J�J�����n��
�j(�E-{#��qp�T9�@W��bYb���nb�5e�5<�fW<h\�M���z�8n,DǺy87(DZ/�`f�<X�E��!	�z<
�w��8-z��]���%��:�p�ܖ}K1�>�����)�)�����W�:{2�/Ǳ�{͟�W��oȼ���4����vjU�Z���V"ހ[���?�W�U��=z��Vc���]3�4q�`gܥ�q�~�;��4���o���2�
�ygޒ�s�aBZU��K��ǫM1΁}Xi�ە��<�3��"�t;u���(����Ф���Wd�_�AS��l��K�h�رG1�!g��ݵ�o���o[��;\2��t�}�� <�~ͣ�j�S!����m�^�}��m�3	�T��Ƶ7�_V��8���6)Vև�D����'�*��4^mk���׮]�M�2v���ۏu��Q��� ���J�X\�v�8^��E����V��W��Kw�U�Z�ȗ_5���.��hْ������R�J[]\-�ޥ�xg0a���F��+�ϧK��o�{�̅����>�e��x8�|&[�Z��>=�d�����E��X�)��f�B�����cB
2f�XN��`b��wFμ�;0�֎,��=U����-��]U�b;��>�gճT��وJ��.�m"�OF��J�u/o�]�T���~���-�,1:� ����2��n�xW��OI��{�{��)�k������,����g���m,XZ���O�Eh��}�0+�9UC�O�|�����!�~٪�� k,H��RYۓ4�<��ro}��!.�d#���:�e�Jؠ\)��QwH^̖h01-�0д�{�_��r=e#^9��fum�jss�{^���-7=�y�i�~���oե_&w��1����%V{B��$�~�!�n�����ԗ�V�^-�~��l��Xvg��g���/���G���L��5趽������	����C��HW�e�`����z��K��Z���}�d�| Uŏ
�}k/���I�"���"��яA�S�V����?\��Լ����B;�Aį�}~@Wa#�r&�VxVƫ���G��}O��ׯ6	x�i;��V��u3-�ۿ<�6T[�cF��Y�����F�o��l��ofዔ�S�ܱQ�S-p�p���#�&��*�\9��Z��f�{]��N=f�٩�f�t�H���Kz��[�z��:P6xa�9���_}8&����~W���y���~^��T? �o�˩��ϫ�}S�:WD��.����ѽ{���w��_�e�25�#ϟ)�����ױ��zj�<�3�:�G�Y�j�s����{�oCno�0������7��b)*��6̣��"�vG��7[x�(5w�Nm'��EZ<)�C�vc���tƭ��x~�ژmLT��r�Ñ����g�'����x{�/x���
��عT��j���i�p�=���÷S���
����>z�޹��vU��}���}�N���F0J��b	�k���P<<�=x:��!�Ҳ�j���i]z������~��`��yr���W�JU�}q�xIX�_V�~�_rӇ��B��Vg�iB:i��E�d
�"�~�>�]�sA��o#%B���b�Zd�|�ӐLX��0�>��͛�����*�@/���+c>?b��i��߫6kI<s�}�n@}ş��k9��i��?h��z�,��a�3�g����WD'1���H��4QJ�e�wc'�vqx2�(��`"�S�'Rʻ���#�;�3w7{̊�٘�%W�vk�:S�6v��*;y��`���7}b�q f���+Ň1Y�M��k-�)���Ү>�ҏ}�}���P�Ӭ�`�:�%鋈�ǣ/�X��V<)�����=u��Mv�{5�#0�ܖN��z{D�N���v+���+E�c�6�
��w��\���ٿgW����w�������)�s�=�A�~��MByX-�x�Ӌ�Y��X~���:����`��A�	�SI�^: ��@����g�MM�g>����֜԰Y�>~@s����/ܻ{�cO�e.dx�t��uwh��X%��� �n<�	�0��Sb-�<6�6���V�M��#��J[���[��.��o{.��KΪ�+
�����^<���^�i߹���?jL�X��ױ�9�x���\CV�9�́4�ikJ�1����ǩ�;��ӓ�&��o�ݧ�Xgo�e��j)ٸ�;@-�����5�*�q������M]�>���쑶��١>��{���Z9��y}�O�{%l�h���lփ�0��&3�5w��rIeG�}+M�S��d��L�������Ta���i����v��?'���]��}�qHX�7(��ko������հt��o��?U	Y�z���n%�K��B`j�_=��6o>���k�j������M����C��5d26�úx�"�:�����[��˃��X7��Np�}�Z|jd�:"훘�+P��6��k~���!�2�X��7����D�fTm�L�d3���XE}n芈E�tE��2�FM
��C-& ؝�mVͭ^	Dy�w��,Ä���{_����'�y���{�~��=��G�)Iev�B2��}���^4���~�}f��z˭aW=^jb����ڗ�:�����so�5����dֆR���uc��h�����:l�P�1SC`�+���s5��C��0����n\ �225�jn!&���5�k�o���p���6��>��Տ�$�0`p�J#KߜȆ*���^�n^o���j��ט-��X�Е����'�<j�y��TjZ� A��V�^���/����P:�@���=�r�\�Ż��M���3��o�k3Ѫ�p���^*Tj�$1L�J�� ��a�[���2K��]��8�I�Y�I�wu���"O'�e���g!��x��*���2(P~R������~�tJ2�|��s~><�1��AJ����U����.���9���wT̺lz�S��㯽u�~�G�.�'uEIvވڴ��t7�tݬ뽈��t�#P��s�Rb*ޭ����Z��L���)��1�r�is&���Їr�[���R�灃���޾�^niP�;��YS���p68Q#��bF�����t뺦ob��`���`mR�]��Զ���k��,��A�x��k!��G8��n�کU���,���9�º����I�>�^�Fff%ͧ�
��sܳ�]KuZ�����e$-.�7;u,��3�uէ���# ��놋}Ϲ�����8g%���m�����Hέ�t)e��I}V��d=��� ��m�����BJ��=F�@[�Wʳ�I��e0(9�1W&\�]�Һ��],�{R���v2�XDT��z4P4ݤ��Ow��֊B팬�7GoTt��.}F���蛋-���n��˳��~�\v�z�Hn�%"FJ�]�̡�����ʧ�� �5`os=�=�0f��m@$z�H{�iW����0L��V���ӸX;�L�(��6���?�Yv��V��єf�CvR��C6�ʎT%]K��.�\̳�PJ��FU�[�f��h#nv����=���ܝ+,�W@v����� x]������c�v�N6�P��'ە2R��/x��*�v5�j�_:sDޗ}��d�z85:��fiU��ޥ:�9 �������]�z�b�}e�C�X�*L��k���:�g[�v]�EF�a�L��
��Y[/�\�V�swo���kȬnn<��/�i7���5'�n��]=��]�BT>Ǒ��])lC�?���e-E�\qT+*���H��ZI�䂺�j��5ZEbӲJͲ��Ū���86�G{�LD ��X�Up�q'�5B���R�ܘ�}8�@k�T��j�yzwr�@W��:���;޵�&�R
=d�K��T��ws�h��&Ė�Ypf1¥�,�� x@�ܩ��X5�t����X/�L���׸�N��H$���8R�'�"���A����+"P�1��֜�i�&4:tT�C�E+�su�à���u�U�/S��;�]F�'�u��e�+�>�4H!z�'[�3a�����E3\�|S���*q���G����М���@�(���Z�=�N�V�����kyL�8f�Hh��iL�jT2����RfrX��^�(f�u��vt�D�7&���Y���j���N˭�ѧ��) ��=�G��5�ML�ͽKw7S %�thO�ڝ�!�s6n>���en���!X�=m|lkr��dfaJ���ss��ڤ��#"�n��Rm�9eޚ4�!�<�qx�w����v�,��wU��Cp�i��3v�:{q��4Lu/u�����0'�:q��`��N�^�DJ�b<7v�2[���S����oQ��˃��T�^]<�=�� A�֛�5��)6ա�;�nEY��/zs�뙛c%��՜��p]�u�6�R�җ@n޽�'�}�}�w����X��{�����Uj�O�\1VT/-rl\����S32)�fg!�3
�-lU*�+�欴���1E��(V,�-��DE0�Kn�J��Q�L�)g9�RQkTj��mg35l��Զ��j��+[X�F�(��
�q�X������sx�2A�J�-����-9�Z�Ѷլ�,�iG$/9p+�#(�أ�q�jZ4�
*ō�8�ek��k+��j<�J�f���f��DJ5*�Qԅ�
�b �mn�X2��mE�l-%P��*��XQ9l&�ʹ�Z
�N1xǉp�kWR���3%�,-��B�mjf���T�B�ɐZ�tAh���(
��H	$��䖏t�Kf�w"#�-/m�/w����OR�!��]7Ȇ+�p#N˹�o�k�.\�����NÇ���o���?�W��	9Fn�&�����6�<�Q����L!_-R�%�9u�!5�~�p�^8;�����	���*w|[��Sk�яEC��8_��������Wd�]O޸�8�ُ!\�a��G��n���s���Zg/��N'�qׂԇ ���5��P]\}OT��$���ط�-�T=���J�U��>����/<�u�E6o����n����B�@�n�4zĠ���ُ��k�z�6)������	�^�����K�ϸ�
��r=~��K�e*00�g��噽�f�Fƚ5�8:� OS���B�횺��1��8�S�\�yUŖ�}�dS�}����ʭ�i���������^��áLH��/��
F�)�d7�N�qq�cgs�]:������	K�!���w�O���P�����M��eW���e��ysb(a~ej^�XAC�,Ti�� k��t��ذ{�Ю�q�{V'�+����S�b�q������SEs��
Wc&5wL_�2Y�� C�S!���+�K��~$���8����#"���h��`��w<1��\��u �}9k���4q	��B��1O^�4��]�9�tR���k�r����9~Һ-K}�z�RV�"��'��v]�T��޷�VvlҚ7��*��Lc8��M��CL��c��r�;�C�������~�S�$�k�g�W�,1��T�^u�N `�����N���`53Ӗ��F<KFz�w_[nj��x�>o��V�|�yM<%U��ʇ�}K\���X���Jr��vn�h��T�����+�W�������yj�w��Dz�_ �or|�V��[ù^T�s�n���b>�����G
߬�e�"(F�0<w��̊���n1���J�O�-���؋���ȅ��W=7�{��_7�>��d�G��6����)���WёieĻ�w�o�H�*������.5,�z�
g&o��χ���u����讼@.t�y���d�������X�́��\E}f���AE3q�J���׆Y�˅:��</�V�Z��^�R�X�>3���`{.�#C ���41R:"C~�{�5l���[}���>�Vӊ�5͍륖��v���F*����T��g?���v�|�<8)2U^Ԗ,5g��ͼZ�fǵK����F!2���1:*	��dC�����Ŗ�MK<<��y���2n��*�5 �T�lT5�)���{: u�f��ֳ\tt��u�ڵ���#�^ݚ;�q�%p�{D�]�C�c�J�fs��[2���Ϫn1%09(��%����Ǵ���Q��vk��LՄ��"9�LWR��\�ƈ
���ԿG�}�;��Rz��:'e�����vy׺{��
�T�܇�J�m��M
*�z%i��<��紸߱
V��*\JR�nMi�*X�E �:�6��~�����'��ni����Ƅ�%fk������_q5�Y�W:�����%�$���[�v)��{�	�����0���E6��ƫ�^Ι�;�\�z�7� �X�y�Iq��=F]�R����{�Β����/���A}K�P�E�ּd��d^H�{u�@�}qm{�X�j����ci�qW���Ma�;gLS���8��ef�y�+j�Q:���k���f�T����x��W�{��A�N�~Oj���=P�2<T5��OWd�`0��<;�O՘����F(X^b���fz��0��W�0-�{�-�+�h`R=t[�^�V�O|}��tG�9x>PI���kR��o��^��ת؀P>�	�׷@hQq���[�3/Ղ��t:J�Fw���w�CԀ���Y�|i,st��һ�mSW��F�"���zi��S!7����L}�zٸ�S9�l����hAlSӆ�c�h����^j}����K�4�\W�}��F9�C�wӷ]�;�{�����r99�<u��]��~�����T��W;�l�.62��x�N�y8����ȟ�����V��Z����Cm�m��I+��_��w���>���e+�0�C*2�3tsr*.���i��E�w����;4��;>�?H~�~�=K����;�̊]{q��ۓiq1*�{)�?#�����.ҟ�3h⟛���(j�W*u��(�77%��aV�x{x�Ow���}��k�OE��o�w��[�e؏���e�CgS�vմolǨ�	���i��1�f�_���M��S�4΃b` �o�ԀE\�k�`����v�~�P�����w��lȪ_���w�j|G�V�n��il�vE|��/�s[�`��P�|�,d��d�6��=��UYL�1zènq���M=gX�u����5� ��oL�g,>�2:s�ַLi'��q`�#:�V5�����aŐ���:$��t�-7N]��I����#5e�T{l���|��?��t���2���v��0�.{h��e��"ܼBgP�p�ޔn�����doVN�0f.�/�
f�h��_���G��>�v�x�#*�5�9�c�߅(���E��x�����w���Vwj���8���RI�,������u7�'P~�T��=
ͥ�#�=� ���^��v%B�ȫ���Z�T]c��;߼�S��q�Y�2�{i���9|��6zC~�.���˥Պ��/�o�{y��g�rJ�dZڐ�V܋�i�}5�������\7�g��8��e�n:#��:��*�!�=o����z�-����4��ם�����Qj�-Ϧ���jR5�S��Ӫsaf4u��SU峉�X̴�4�[G��|:��?n��5{_I��ߝ�PqxsU�}y�3�>o~Q���ӯ������;��S���N�8��
3]������E�]����ǜZ�g|b�bn��W�gll;�}M�{�]�T�>ej���7�U}�ڳ�R�-�͕d~d��Rї�d�2Y�C�1u��cFҍ;�׆��q�q��kR�룁�ك֢ţ���"���o��z֓g�Lv9q������
�b�-��6��#[�<�=�cwu��`e%YY�V�f����[�k��� 3��^�Ih;k����>�}�F�i���|7+�x�(����\�kia<���w�xi��E�ں��텚�)p�ѨI�q�	�J�s#�ϖc�sW`�C�F[·�<}3yh��{�G*e��2��|�{�Ot�/X��VG��N���f]n������p�Nc6�
s�'�-����t���"�-���e�`������3.��1�gx�zTZa�!���M6̨�媶��)��$r��T;ؼ��'��o��ϩ}3�(�/W����:�^F�N�E��=A�yud����Khײ��[��\Q{��/o��M�Nɒ}�c|=rM�ܹ3Z�������W~�3>��>>��/�0���G�[4�h��^��ǭ�)��3��Ȃ�zMw��^��t���G���N��[ǹղ��Mi��:[*b(�m�ݯ:�z���M�-�m�%F���-K���<s�f�n�_�%��Ċ�IR����2�w�{ǯ��}Z+Ҽu�4�=S����b�~��L=-jo",�WR�ެ*�1q�kE%)���m�*�K ~�f�1!��ns's��⑲3�"�{�0Efs���@
4�舏�"!Lݤ�u�����YU�����;�T�MSp�Ѫ�Y�V�7
!(�����fs(�RR��2�J�5W��~�2�����=��8�Ҟ�~�|3#�V�t�Z+}^[��p��EI��W3�š�9�?��m�fi9g������^���l浍,��Qr�z")�$E��Z)nB~�3������ȹku��[�y����ꄚ�B2)!�Q�߭[Zr��|ʧ0S�C�+������F�c��kj7'j>	�PV�W�7+���4�����iF�ͅ��T�i��
j��i��+�������5�ˇP���T-g�o¸qA���Z�<��6�|�v���>��_eT��y�R�y�L��6&F�~��ď���Ӗ`ޯE���@���:|�e/�{ƱC�e��Zq�����qz��S���G��f���b�;�h��V�R��{��.8�6�����"�Mw�#���o�;�D��%��Kr��������F@���K(� �h��[*y��|�5XM�2��V��u����y;-MWJ���yNv��܋�w �k3�w]�kguȲ�Gl/�u�:K���T�I-�]���w�꯾���w�N�5��S��L9yji��jǲ�e��>˫u�g�mT��l�XƩ���-�ў������?+{y5��SX=����#KҶ��PR�	�Sz�Z�3��5g6�J�C�WP�'�c���R�[(������zK��^���]�r�2}�0��Y٥ֽ�x���M(�3��1����1��ꎞW�dم��io����8{}��s�4�o����?){�<V�]Ӷ��=��}�̨%D�Ҫ�r�;=�{�'�ܫ]�T�OfS�܆oOf+�U�=�w��'���a*eFW�0�QW�(����w�����#c��h�����?r�_o���}�P���
��*)5P���U���{�y�/1�uQϭ9rƺ�5����^�O�*�<��/�V�6g���ȷq{�>g崳�D��$��eR���Y6��y;�9�j�;��Dun��BRÆ�V�G}�_��H���k���@|v���}�h����g��4p�FT��oM*�E�:��h�a�CVf9@U�&���gQ(kAL��f�ՖW`�u��W^�R��;,���q�Q�����U�����V��Z{���;�y��H{�=�0�YO��́�O�<��ޢ��W3{]��oghO+s�W��̣�~4��0V,�u���ŬsQ�/Hjwk,kM�s�uH��%8Oѳ-��?5L�!vw1^c(*o>y���;�ͻW�eS]��^>v�@g���3�����׆��Ny����h)#=x�NTg�3�ǥ��6��y�QӓQ�ם�ׁ�GZ�Of�.�_�v�y��+��Ŵ���R��_����{{�<��{[g�M���{�˯�����$�����k�׎�]K��-��*v�o>�ˈ���^\�a�����=^�6����%p�u�=�o�/T��-�������_��^zZW�e�A���^�~~:��AR�D�KME�Xf��ʟe�<��Sgt��T�r��F�{��{Xi��o�goݒ�����w�x���Y��+Z8t �Z��t���]ٕ�M��D�z&��J����r��c���Tl$�n0V������:�ݼ�Y1г�4�aH�e�ٺ�Ʈ���ꋇ�� �ih��F����^�ػS�0V�V4v��z:Dg>�szfpm���}��׮wl�k.�?:�Qe�z���-����1�m��Y_<p����Uv߃���"庝�-�T]k6��^�S�ꏙ]K��x�l�s��u�����@�E�l��.��!+��qh|������[�og����N����y%��W�Ƙ���_Bڥ+56djD^Aon��/��co��×��ݔ��5�ǂ~��mCNE��T�kTF�댨ɻK	��%ݢ���"$�p��l���cfN�h�e��y[1��q|��*<^Ջ�W���q��[�׾=c����j���
|�θ�_l�u�#q-[&���i��7������9��?RLe.Vq=!n���N�[�v6����U�5��n������c�~	/��N����u2��
&-0��~9��ҽW&W�r��y���a���}���I��,K��}B�gT���Haܳ�X�k����n���*8콸���V����չ�|�mv�=�ч��L���F�i��k�Ut=R�`�9�� 
ܣ#���6��,HwJ�fXsV4�J��"��^?������Rv�[���ʔ;ƀf��}�n��2aTGe]cj�l�u&���\�G��3�f�	��x.���=�/k`��X��e*�P+��}�����O{�S�Z71�]�:)wnT��,�|��֡�l�:��}c��c�=��叐�������t�N4�¨��ɱ��34m�[��Z����^�z
��Zy<��1���a5��&�r;+:!js��]񩗤�u�%k�jT�x��D���f��{}Y7T�u �+��y�kA������@VpB�u����E�<��}8/�n=u�P��1m�];���@^��aR���w�{.��CG �������~��R���o�%d��ЙFp���p%ݗƦ��@N� {/Ok��<w�l�8ե{���ʺ�k9+���cﮏu��y���Ou��7�S:�(��-@(������B/Y�;J�"+�XsBҮ6��n�w_�R�`��&��1`-;V`�xM-&�G�����㷔�]-#"uU���jV�������w7s#���y�u|mu+m���j�3l����qKBn�S}��>T� �	.a�`!5�μ�U����/]I���QV�{	��ɷ�=[�o��&���g�ypTde�Ego.W����DK���Q�ә�m�޻O5nW	�n�U�3'W-�Z��/.�ܶ���<�Δupܠ4_"������hxy+QV�uh�N�y�sQ�r�}�grĸ�*�Lm����P���uQ�t,��/{�YHk��Qě[��L}c��u8@��k��c�e�0wP���i�:���Ob���(�ֳW��#vޫ�N��CH�5��y�p�(in�Vҭ���U� JS�髍u�t�ܜ��!�ӭc���X{��]y�WF�{�ܫ��{}Y�D�F�L5�G�2�X��j���N�WNP���GY����k[���=�F���|�܉JUcz��)�ly��ά����.��4o97�uN���s��f;�K1b�ھ�̼��9�:{�*�Mm�Y���T�d)�k)q��#���[�H@�E6����'�z�Ӹ��k/���)����ai��y��7.\�	F2�&���H@�o%��ven-ӑS[�xei�:����x�]d˥B���֟neż*r�E[��ۃ�pl�fH7|]3��V��X����ְxƯ���r�e�^��1��0� i[��;o5�v���w:��WD�wz�,��M�C�Ak]&Ͱ�dغ5p�"��|�����ӟ���A��/��*,���B�j����9j�4(��k��Cfə��+�*d��yhX��[[�.�I���
Ų�J�-P���
����-�欵-ejZX(V��X�R�%��L���6�mB�QDk[KUjRҬK����r숃���QJ�֕��
��!��35��V����5e��س�l͋˰Uh�kQ��T`WkR�TUV��Ƶ�-��b0k-mKEne��EEe�����iEj���TT�Zƍ�EkUEmn�b��)j5�)Jԣ-*!��-�V�1��(�2ȡb �������Q��r���h�J��ѭ�KJ�ՊJԪ�XŶ+m�[l�TDV��c}^3��9G�v�xk-��g�w�ϩLo��[ު^��Jf��:"t�F�l�����ͬ���gwd�������\�lG��@��Q���ѯ��߈r���t����_��m�`[H�ڕj��D���L*Fa'����6�r���W��8{X��x`�oƛ���,�sQ��|�'�S��{ˡ�Es��t��\n��l������n?A�Amz��!��~"O;��r/N�[��7a����˻�M\����Ey��3:�}Ү��C��X����UN��- ��%�|�67Nz�T~��:�+��J�򭣳�Ot9�u7����m:��BG�1�����'��?z�e:��R�1��Pٯ�b��J���2�[����J��VJīu��ڈk�\c��(�r�_�a(�9:�n-���������V����3��,�m/�K���A��W�Lcp�|0%��\7�-V��~�����Z&�	�̻��wa^�?A�ڀ�4S����LR�cd笿K�Q��.P�J] �}"�gm݀��0M"��E��+�-R�t�ZϚ��o=�g��%��x3������p�h�6P���*�R�y�eq�iq#����[T�6ZT�q�ΟWtd�5ᆻpp�U��x�X�\f�OiQ9�>#�V��mJ���U}��aގ{��n㧉��������͛�L����)��^��C����#S�Z���g;�*���Uҧ�\�{[��&1r�m?,���U��>���h���S6�\;��wT��3Y��h$�'����X��u���"e��5����!EkA�2�7u��&c[����b�˜�=(1�ggŰ�X�qL��έ��/���=8���}�,z�߻&��K�llC��$��u)�K�c~��:���J^-�;����M��wY��1V���=�OG{O�RX��z��0��Q�Lyo��k4���=s~7L-b�a�٪�9���|�鸡�ޡ���=���^��^�ը�U��Z�>~7NCۅ�{�w�W����rnҖ��ek��0"�����j�={�=žȦ�C����p�J���^ٸ�o"�.�)�u�Þ����؝n+���5�(le��
�GL{K�R�͋�8��c/q%�g,��՚��M�G�s�C����G�׸c�ȓ�,\�n˷Dx�O5�%���O�e�7Wt�4N�,�&>�z�P�t��St��vJo6�κ��=t-6 �Z��n��^�`�m����Y|�����_UU|�Cjw�AV{g}�[���׍y�n}�ЕR�W�nW=��9^��:�M�m7oOd����d�����o�Y��6�?r��t���r��GX.��=��~s;���:��>�ſy��A�y�K\�����A�.�-f�yJ-օ��{|r�T���C.y����zU{�%����~�"��[�����u��x����w�D2�ɕ�����Z�nu��{2�|=01ccDo�n<�ر�}�7�a��y�Uj�T
λ��%���o��wPt��R�����ۙ���f[����P�=�eݝ�K�Z��D�1@������`8�mS�Zp|��B��*���v�覺9<�Qz�r\i,Z�������|���/��D����ߚ��d$�XKt��A��F�9��%�R8��R��>�:�������觶#��.i��[��-�%b&�����ޥ39<�ժ7Cy�,w���/��"i$^���WN.c��>�Ҿad[��M��kd�E�k���3P��o[�3\@=V;��Vz�]BZ�Cd�W�9�or��Υ諭���T���~|X+#z+l�:�����^:�.��LyW���DZZ�9��T$�\y��#ig�F�F�c��k:�U�4�����n�M�Y���2���4j�c^�����g�B���γ�q��k>�܅�^>�}7�+��up��v�NBM�7����\k�ɼ�&�ήm�����o?'~}jwt⢬���>�Zv{h����k�R{��p�����^�33��,��^Q�;#��b��
�Ϸ����M;�"Mq��X�~P�g�q�O<�E��, ��Uu�U�׷�|��ހ����h~��F�͉Y�+O�<��Z�O�m)��Ê��*s+qo��D�^�IU��2�.��5J�C|<��թRњ�,����V�1%0��ߢ�=1v�l��-�z��{�Ϧ�\����ܝ��:\o�<��v�+d-��_�n!��]��-�l�qT��
�7cR�#1'vڀn���WSwmɟA��3����x�toTX�H���eL�7%���{Fhw䍩�$��+����-w� �w��Eq���)Ӽ]�k��}k�]�g���s����']݇�I��1v���mj⹶����tQ�l^T��S9�W�}��U~�L�q�М��z��¹�
|��k�vS�0�4�v���E!�^ɽw�%��c�g/\�n�g��c�g��B�!���kKy�>�R=��-��cNwF������G��3�������?;�����~N�(p�[|c��l�:j׌��?{�ڐ�����o���R�1��L0_{��O��U�mV�����o�]C���ymP������<�sZrf{M�b��uq<[���pAN7#&!�T�O�W�Q��$�����»���6�<h秊Oջpϝc�U/<�5j4�⸆�k��ě�u��a���+���D+~���Q�#VqTE�����Φ7�-���;��%*sE�/{ʉxy��<���(w��Wq�(�/v��=�o�c�u��N�ع��x�I�^i�^�Da��63���?z���T/\mdMydUֳV���S	��N̰��}�Ĕ��,�=���n�0$����jQn�*B�����h&����b] à[�,�omB��9[hr2��/;��+MM}{`9f����ˡ�a�]�\N�s��fV����,���߾�"#�,�1�oVmb�i�^$=N[��ᄘP��;9P|�*.����RJ�voz�����F;������W�?.5}�uf������Ռtܝ��׋�N�
ܯjb���cs^�8�@x=ICU���0�=��y�fS��>P╏U8�FL;yp��lk����F`�T�����J��~��;�]�I�K�W�м=��V��)��fA�j��k�=G�W��>ɏ�,�� GE^׹�+~�}4|�{[�I�����R�|=��܊�m�jFTn�Y��V6�Q�4*=� s���f�	.4���c�)wK	�'.,�k�}�dY���n��=~�����lu½�ȬK���#�3��CzO1�P��m)��^s����LU� %~�5�}�vf�V����Ӥa��x��ſR�^�}JuOg�Ww�B�k�[�w�,�}�<ȱh؅�Ȱ��d� �kSrVq�A��8W^Zީ��CC�#s��Vf{�8�a4��mu��1��&3Cl�:�r�	>�!V�s����oa��j3��Yc�H��慍�Ƴ���k�^����;&V��/�Mΰ��wvull�=�E����v-�}��ﾯ��	2w���������n�lc�(�Q���P��Jޱ�oY�[��F�N�����.O�ߺr�}�Ov�B�=8�1�_�ަfJ��J,z߷̮�\�H�%#ﻕ�k�go��{��T���w��o����^L��/Y�T¯6�^��?����ַԜú�8��������?Sy�aW5jb��^��s��B:ߥ��-ڈ�{�ƽNi����HWw�����"�|���od>�q��
/j���{���OI#��&2ߗs�'�˯��m;C�%�&�{���U!֧/�,�>���ty�jR�7���oǫ�3���:ͺh �.���C;��^��_v�O��m-���t&U���߷�n��FY z
�^�>Ԗ���5�W� ��
���w]�Q�y��ͣ�n�c��-o��2���o�#��P��I�J�sC�>X��ػ�����V:�1Z�ڑ����gT�Xщ�PJ����{2�,�5"&^h�em$47&���M�[��,9��kc �j��`Uc���'A(eGwyM˨U3�� ��r���c��]m.���n>�U��Gѕ�n���OI�OB̝��X��8�Q�-�YӰM({$���o�B�|���n;�=Z+2����7;T��!�p��^��U�a�e&s�;޿y��Xm����h$��K��:]C����E���S���S��f�nmy-�5���63����v�7��8��R����ά���Q�o��9_�+X�S�f� w�[g��*�'���{���kFw�m���}����L�jҸp������������q*.m+5q�����` ��ק��Zw{^��j�^�P��׋g�o��%Z7ή�Zc(���Ͽr����c}�g�x%��S�V�"�u�u���םgW��/t���6ʫӵޞ�Y���U�����;;h��<��#]���z6i0��q�5[F2h�UP߼v|��/4�y難W37�4����4�e8ި���b2>Ӕ���e�
.{����~g޵:���f��9�� ��'�3F��&�S����Zմ����lQ�V�B��xsM]�뼐��q�dkWt�]��ReggM��VJ����7)р9Ɔ:�Pɠv�Is�)uB-��Ɵ�����ߏ������+W�kf���woԄ�gۋC�k:G�5&8,<�<~V������~�b{ˤj�]��������U^�H]�e��c�^��Jq��^f�����j���-�݈�HD���o�S�YF�o}�9~vI����fd���iǘ{���Zh��S�?*�1Q����{�0it��*g2�vL>�ڙN@Vz��tZ�g��������2�,Q��<��=T��x�+Iq��~�gۙ
�����R�g�m���z��Z+k��_;C�뚟�k��}U��W�0my�^���z�f;���}��f1A���X�*�>�=۲�r�\��y�~VmT[�~D$��X�w��1�0��z�9Cz��VU/E�j���މ��܆�;�w�xV[�"��
83�{!��ae+�O�ld���T�$����~��Kd�>�r~\�H�.�B @y�^?l�����J�����7��5tWfu��K�}������4��1'���녽��u�*�0�0���C+0������̫T2��iT7][��t��zW��K:����c���!oŎŉ�i+�}��}�˟�}_}U]�z�C+Wa�!E*tc�i��G�û���-����n�@��~p"�I��SF쉶����4���8�=X�:�׫f�Ц湖IJ��$w"��=;:��mz��6��;��j��}ʎNuDt���v����h��Ɇb�z��{�����E��c�e�����ؚ�ȫ�f�-��KG���%�1�X��\_��v��gd�M��K~�0�2��鼃�q+G��W�d����yq��=��o��������)�5
]:_%Ϛ7���Sf��Sχ���ɽ�,+��o�/v߬c���9��ƌ�@���:yc�^}փ���+id>F�7]U�~ad��p߇z�=oS���K9�ݛ�@��Mx��g���V��U��fO�E�r�-�
#O\�'��{�_?r�Ϧ'Q��{~��U{��mL�M�|����ʥ���z�_Z�߹���R�+aU�P�9�� �sA��Pj�y$�eh����Y9|-���n�{9<mZ���+��b��S�M9Y��;x��EX�#��#��p�S��V��\�j��e n��>��w�wܘ�����.L}���}(�\��ٹ�eN0���Y��l�F��'|�Mh�Ԉ�*b�Ԗ�g�������@橽�E�=��W�A�~C(��pt�Msm=C:p����W�����b멆vi���*���T/��g%o��]����6�u�����rFF��
��'\F�i���dj��q�.WR�����n��S��9�f�SF�[�Aʃ�u�U	{�-�$E�S��j/�]����_R�__�e ���%���vAQ0��Uw��[��+PM����K�}[Hp��Y|�>B�Uͩ��7�W7¸��$����p���Z��нK~r�Tt͎�:��pv|v	��Yƻ9w�<��w�aAF�k�q�z�m��ԓ�~�	J�;�K3��՛�
�Zw��qJ[2U��غ�fR >��:@��N�%���Ԯs�cʧ[�.�a�n���efv4 ���2�GJ����%dξƞ ��JS��S�.��_g>J��vݥ��l5��d��#{�0�|3�u�F9���
V�]b��� ͙�u`E�gKς��]	��ڗct�����H�^�[��$�@,�7�E�]��]�hgj/�^�BL镅�7-�lř�n�I5������/��x��x�9×֯��\���-��o:ǜ�1Q��^弱qC*���B�x��|#κ}/q��)���S]O�#��3�Z�l�F��8�j;��,a�6�·�S5�V��	z�EK{\��V`�;q���om�� �:af���V>���/]��0i�{6ٗeĩ�z2��;�čp��˼��i�5��9ଵ�l�ǜl�T@�v�u!��/���^/�Y����g�� ����u����|i��^�Nı�*%Y����s���%��[y�h�����U�8U�அ�m��Ɋ��!�� ˮWY��;j81�RM�	�Ά�\�*�f6i�Gi���S���<<��e��X��ə՜T�Z��p5h<w��$E;�sW �U��<F�ݤv�TwG-.�#�R�ݸ��{,QyO-N�Κ6�[�=�γ+)��z�RD��*U�����V����N��yϮ	��5�їO�_]t�֫	FE�f�RR]�+�hkԲ�6�j�aJʥ����>"�c� 똟�j���N�uIz͌�����(u�1��J����� U�!�z��r��V���ޒ���9gvq�0�� ݧ���]	�9�O
�N���GR�������l��w:cw1⺝�۩�[/���&!�	Ep��r��+e��FIy����񒶈7�q)]
Z��ڗ�q\)��pS�pF��m��eIp�V���r��C34�Н.?�����o!�Ęn#���x{�l8�nṳ/��M�e��A<N��;�VJ�շw�0�sY�fJ5Ϝ�y�"	]�>��N�GPuVGŶ�Tj6�[EiA(ڨ��D�QjU���[�AB�#����Mj4m��Z���a�Au�!J+D��kiTP�laZ �Q��T�֊�U������WR���]p���*�(%[b��6�E5��kmE"���V-k�V�m���TEZV���Va�lL*����E԰iWZᤱb[X�֢R�U�+�D�E�UV%�Mn���b6��EQAij"ĺی#�UUE�
�UEmv�TYU*��i�[U�TTWXVշcE�6X�����5����QTb*�9��R�D�,�,EB�]i5
*��)]�*�m�Z�V*ڥTb� �:¢�QDMJ����uR�\kkc�E*]B��KJ�)l��(P�I�MS����KIu������F��	�Ƭ�o^]�7�k&��Bf���Ug�wb���^�$��A8($)ny/�G�G�L��zu��д��{	��#�?5d��X{�e��#�� Y��y ������c�sfU�&��o�םq��P����o��o������I稖W��Ŵ��k�l�Zm���ה�\5����5����ٽG��z�0t�\4�-�u/>��������Ӎz��c5��e�cy*T�7Ǧ��S�m��QP�gQϏk��K�v�[O�N��aL�za����q	�Ba�D���\�J����~�'�B�i�X�/�b��X�/^���7��=�y�	�S5>�q�u�������{�7;=6@skf[�����:lN)Kg}�4�}�)'No\��ĤersW��W.򽲻���}��]���e��S^����c~�������O�o´�(xX��K;�
�ik�_�[ȫ��E���^׻X���8�r����$6�Z�2N4�Y0�~L��6�9�s�.�*��4vE
o��fά'F��*�j�ɧWe�)�i����)geJ��^���+�n���<��skU���ԤL�D�@�+���з��d�=I�gu,�z3��c>�|?}UU�W>>�u{���.�7O������΁�yZU�\��+��>�M�/��T��V�^�4�!�� �a��yQ���@���9����V����^���牍Ck[�O0����i_�y�[KO������[^��Z������ӯ|5��8�1��+��Nu�������>�����s4�+-���y1��n!8�Q�-¸Ȇ��J�І!��(�8nq���BgN�/3��b3����[$�'��M3t�B�/Ԝ�jc�EmS�^%��|=��)r ���K�<��ի�~�G"���#��nq��y�E��e��qh��+�G����*gWg����<i���k���	^���U�,m'{���	/t�U�g���/v�R�~��G'�p���O-竕���jw�����f��W��J]Q};�잶��/�bܷ�*nP�����A�WKVC(�>���_���uj�1x��#WS2��(7���.�46����d��P�kJ�����,}�p��ߵd�5���f��!ջ�ui��i�%kn�'Wc�^Y���Q�J�+���">��A{	�Φ_�<�m��j�T�oe�܈O<�G���{޾�QR]ΐ��M�k�/���Q�5��V���/)�׫}�I:�s{�j�`�r�]��3�o����^ֿLu�kګ{�#��������]����y��ԚQh`�7~S��N�=67�1QE+��\�[7&�|�h����4�e8���4;�)Y菆N�o�^h|�U�K>�kv6ܫ�0���M�WJ-6�׍�lZ^a盗�ޝ5�������Gپ��*��X՞�NOŽ�X�t���o/TN��	L{�C�@x=P��V�f�p�u{���V���s��ncXt79zu v��̛�y���a����K���y�Q������t�_�|�^����\^f^:�2���>�X�^�o�]l�w���Bt�'p����F��%�ۓh~^Ľ)&+	w����/n1��⥀�}I�?�Ĳ��w�^��cҦL�xw�I��ά $Y����29�k���{��0�vH�A<���p`��L����׺:�F�L�/��δb=slN��go:���H�ɱ<�3w�] ���u�<�9t�y��W���s~��/S�W������#K�/��A�Ǘُ�ίk�s<sK�yGc���%��e���N��ɭyux�����ϞY���7(0��������0z*{:�o�L��^�k�����Y�I��:q`�ҽ�罉�;���q��(�V�M7�������Dܾ�O`nx��A[�̲Po��s��`ڍuN�<����P���n�$.f�t*kؚ�JlW�V��J�i���!�D.�#ӝ�G��ǩJ��r��Mh�T�#-����k�;_Fͤn#k"��Ⱥ�QDt���>k4	����~�W�}�s߫�g�7�׽^ݮ\��Y��U��Ag��y���?F�k}6�R�Z��nʤ�*ӏT9Nk�	_�5O���ڜ�	߰�]N�፷3�]8R���L�8t��ko�Z_�Q��^8ɧH�'.U�J��K��Sv��~-�0]�8��y� R�Q2i�k��#�֟�x1������sY�5C.������>�G�.��EC�^v{�;�g1d�P�d=k�C!m[O0Cz�%��z!]�p�ړ��.ùK^�+6������ukU"9�)Lg�Y;�G�DC3�uk�8��u�*�]d
[�q��^�8�}��j���.�JU��)I�;&����Q��oF{���'��O��Mv���o���g�C�X>H��<�񹆻��reA~���̽�s�WS��(tUZ���ԭ;�]�Udd<y�O��������m;*6=0|�{[�,:\��_w���˪&�z�U���x�t�M�U�[]�J�m�^��(��co�r~���c=²?W���5;T�HQ6�uμ���Q8��>'~�)���)��ō��˜�oƾ�-�i��E�?^MCya=�����T�A;<�;��[�`��堞���z�P���o��| e�P4<��t�X՞�_{��p���Q�=�^k�v�1�u`�<�ﶥ����SӁǾ������m�䯺�M�^�'�B!v���n�٭�`m*
�^�͛�6�b"���E�k�ABx�\��
�t��Ա]6�cBқw=Kk^��Y�%<�Ӡ���c����jgeIh�w|��3p�f�A=Qδ&b� ]��;�{�hP^V*t�γ8q�g\���[P��h��S����UW�{1��>����s�9~Ӳch�+��MͶv"n����́X�U��XJnSgگԕyU�-͊I�9�w���p�J�*���YxŚe���׆�#	�{������Gt/}Ϥ���O[گkq�)t�P����#'23Zr<9gۋC�G;���RMw��>~]IІS�n�ϗO_����g��j�WO��ۋC�O׽�yZ�ڠ������v�|��$k����R����Q}bUʝ�=�HT�im,�yW������Uҧs�9s��){R��9ڔǵ����2�������V��I֗��N����+'<��.�k�\g7�6*�U���S�鞩��U�O����V��
���U���%��
/=O�x9x�U.�l�v׻<��*�{�#��IM�	u����DJJ������ɻ�P_��ޡ�������'(�u���fAT��V�P��X�2C�* g�+�T���#���	2�/`���)QjI`�i�!�l,GH�Eb�7�M�5���(��q��K��RH����îa����bA|6rq��ػ>8U�z�gN��1�齚/m��`ĝs�����η������h	�a8�~9��2s�����1u{{��]�[������z�rz{l��l#�|`��+�qo˩{_V����ߛ�����\�W����+���V��z���l����i�b��h��J��scm�႟�s)�bU31�M0�ګŘW���Qz�G\����g�)�[�{����F9k����k��Ƨ�B���γ���Y�{��Kۈ4<�9g�*����5gU}e�c�j�nE�����/���.c�K�8��eyN��z��p��[��}Z�������w�]���#c��6̵�9�yOQ���x�]]��:��P|�N�=�N�^��R,M�Wg���.�պ��{HR�b5O�'a�(yz��KNdEt�jk�T�޳����o~�w*"�:r�d6¯��Uc���T��C�-��5a5���B����`�f��{v���<��T̼)��Fj�L�PEqn^���|�魞�6�(����$n:C�QQ��4��>�b��x��x�����7��{�.���1n4�oh�QU�y�G��C���.q;gRW_<�*���>��Μz[��9��7����{ʠ�U�x=I'���"�Ij
�
�X>���ΐu-���]���oܑ�+��0�7'jh�Fˍ�O!�g���R�ԡ�'ڗ<�W�-?^NM�{+I������2��2��{���׺���G}��t|������`�*���w�U�����P�����g��M�3ʨ�8�L=������\9z�g��8��R_����łD�n�jQ�n��ʉrWѬ6ʜח_y�>��K���v�o���e�ya�S|;�vT�����`���|��o�u�y4�]|ՏeÑx���sm@�^6ϵtަ�����Ʃ��(�^q�Qj�j>Jߖ:�1<<c.�-��p�q���>wl>�˱�����E�u�(����7V�_*x�}E��R��-n�����K�C�ya+�+0k���K��ߧJc�i�w-ڈ�]�M���U�V�;�nY��]ʵ)ǀ����Ws���̗]k1N����q�<���^���ް�}GR�\��;���ss��B�_O(k�8��j��=w�{Fck>�+�	D��쳴����}:3.�P��:�����_P{�#-6��M^�Rݨj�{���+T��jj��r����ߨ��[}=˯"Y�VOp���oݰ�?3����Π7�ޯd�\��Z��"d��}.7X��9�k��+d�[�����2[��m��#$����V�z�~��V���_�*"�3V��ٞ*���5cY,ĺF�\�`j����As���/E��CiYj`>���gC��w���н�~V���ٰ�z�<�5 �����u�q������eFL;yw�{ws��:����qo�����%��b�҈������E�i	C�<ɋqV�ͧ�
��6P��L�^o��W��]@P�FˇQ�5L~���*���I1![�79��9Z&��J'�dϥ��͐�_���Ž�g!= �_�9��]��Ɓ�S3oT�V��+2��?W���71�N�HQ1i�P�����d�~|���*'|+e�^����k*I�c�aӿ�a��KB�d����1C��Q)e�gV�빹O:��ߍd���P��I�	����W�E�y�no�U��˾#�k�֙��pb(�DcǧWv���f]�Ҳ|QI��6,b}m���Ho�-�2y�E��y��L��L^����Osҍ��6b}jL?L�e��ݽ�+�ox�Y���.\�T}�Ƒū�{i�,�B{}J�������8�u��z���3o��]��z�Q�ch��x�kA�&�qii�����+��j�;�j�Qo��f��-�,�˴���t�X���Ξ2�I�p����~}�����;jf����M�Y�]�p>�C�r�Ǣ�>�2���xN7�Ҟ�k�>��ؤ���{�z�����5���_>��˨a4s�핛�*ӳ�Gt/}�[����_�ש�7��N�Ws�-�>�`Ȯ��*/}7�|�h�x�(��S�.~�5�^Y�3;SZ}=����=������Ş�<�Q+�Z��f�ln��z�䕩�p�
��5_[����|kj�eFLSyw��L}��b�o=����Q��v�f��5/���Ն�Yn,��}�U�|�T26�`їV��X��X��)ث��Y�9Lx�6�Z<�q
D���cs�����y� 	���|�><�]��Vؽ�	B��,���S�w�{���W��nk�~4�tt4����K�EfR�$n���t�WN���nl��J!f�1ɛ�K�]�o�U�m��d�@|���e�8�73S�rt���d:>��lL��[��Eq�X����Y�zR��Xgrj;��;h��)��?X1��w�d�ЧO�� Ȝ4�"h�}��pO D]]n��*����)��AW��s�|S@�́��޾�t��]j�dÂ�iݫ�G_j�]P�4ؒ�6Z�*p�0R���Wt��do1�8/13�E	��B�Es���n�v�����d�,�BO�Pë��JK*ww�4�{�h���W�M�G8M6��{3��'�;Zi�+/��秶om3M�R��hS�vK���]��r�ܾ�)�h]L4��p$�;������>v^q�����'�I� �˧�e�,T����9;U�5.WK���7.���k3]�:�&����S j�dT�Q��;5�^�{��*�μ����Qf���|��i�h��T�T'�X����߷�-ǭl�ջ��R*p��臆��50�Zh��(")bJ����D��)e�wbYR�=J���!Y
#65�����$]9��Wvs�s��Jʜ1�`o�Dd�{�Wa�:"cC�ӄn.5�X��8Yu����n�+IWU���5Չqɶ���]%�3sg�ӏ�M��gD�F:ŝ�]��K�S�ΜA4�P��qјn�`��t�:t|n��]�w0;��������jG�q�i��<��!nq!Ɏ+�]J�eC;(���+��M!�	��g\�0 ��O�B��wAᥴ"��=r�r�|Yr��*���GN�M�� 6� �sM4]�I�+��S5Ǎw�Z�٭�CNSG&_nU������M���A���˒��`����R^�����pM����j5������:R�F�Q����\�Ǐ> �j�T��{N�d9Q�ӝ~�������Q�]X8�VX��B���6��-�5ݕ���Sz�u�Y�*2R�1����I�4�啷ׅ���|����.�d/Z,֙Z�K�c�Ba�w
�Wwt&z�⛭HN+^��]N�2�5kP��׵�w���4[�E�䓹Q�� �����b�yI͒��cRc~ڋ���[F)�;��{o���'s��9�u�����o.:��h���qY�i>!�ý&s���J1��R�	�+x=��&;Q`��RˬN���o�r,7������G*[���B7�d�U��j�S:���o;p�A-��a�r�	���7s@;Dx��X��Ӈ�����J�h�g�T[j�j+�(�:�F�u�UQ�c�k�R۶�h"(��kUQb��԰�Uu�(,D*Q"��-�JV�1b[U�.���VQ��VjQH�����J.�q*Y`����[j�&�2-]j�%H��)fWku#K-��E���V#�bꖚ� �"�"�&�Uc*QUDEZխ�!���c,ijf�(��*,cj ��V(�1jTPF
��kv4DH��T�-KhEm(���E�DUTm�YD"1+DX�J��X�ڈ��\�T5��Z�VK��ŗ`ȂȲT*Q�0f�[�h��2�Q�bĭ���������m�Z�X��c*

�l�Y����K�h1��5,TX���ib�#XQ�]�X�QB,�6�d����¢9�H�-��lm*>��+�M��q�d�X��b�/���H_ۼk�Zݞ�Ư���{���Y�|&Q;%�|!�|cטN��\,w��}I�����&/�6���Ǫ58O,�+f']��]G��`�O�t���r�!-ax`�2ߗ�a\�~ܝ���]Fˍ��&ۘ���ιC<�����޷�G���a��%^^�k&6B��'�	n�-�5;�,�=�C���� _?U��/�3���V'�*�4�i�yS	��F�jUN�F����@w}u���~v���X��z�|��<���l=�9����'�W������x�?Kx\.�y�_�R�^1U��rK�텷���z+�j%c��ŗ�3�X�9�\�U<�۫�{�*���^ː��)fK�����ܨ���3��ݩ��m�ܕ�~��u�9�Kb�ȼ�j��N�{�m���+��ەN<���q~BE�� Y�3�^��W{Ϟ��x2��5�G�"v��?1ݿ>ܩ�ѯ�{�)=@�w�%����
ǋ.5����3��YSү`D����Ǽ7$h��<�f^����,���T4$6=��6��M«i@��U�{����K��X�Xj�˗�b��"�Hek	҆�޻��AWS�Y������Me�j��7����{����>�R{�7jiT���w��)�����f��i��Gw�wL}�-�7�ɝ\2���8�n5��o��iuv�xus�
�m�T{�<��s~�Nn��E#�z�������ݵHJ�j���>G||o���:��q������^n���:��V�|�7^����a
���]n?{b��p;�w׽���*��f�������s��S�ƌ��;�
{����h1P���6�R�D�檫�$k������ޮּ��kۣ�cy�}%��R>�YJ����7���lN^N���/���K�z�xћ��.�{�����)�w�5���7��>K�ߍ$�%��؝E�v�^Tgk�I{?�
~֠=�!���5�>qDw��c��
_�[�Y�D\�u���k��}Π|j���r�ח^x����|�D��^mǹj���a���
��X�.�J�p���޽ȱj"^t�"����d�y��N�+�>��ײ^�f�;�֧5�N&{^`q������pgi��o������|ZU֫�ҡ�y��1������.�0�'�2�=BC���)���]�������|�n&�5Y�Ň��ʉ�<��}��.ۿK�i��X�Ӣ�d�ǌ�b��ی��pV��}�f��^ߟ�e>�S��k�Ϗ���{���t�wue.S����Ciz�%p��S�������y�ը��
&�i-,�\a��S�[���`J���6��B�#Ӌڷ�=7ǫ�=o�'�:�:w���~�����;k��7"i���[�31�v�;�S9�6Z�R��v��}�����{6v��W�^5+�����z�p��]���^-�W�qsݮ�kV��=�㌖�e+�0�P�3���� ��؝?mF���tJ�}C�Ts�uG�}>od��*���8]�.���2�kղ�y�6��Ǧ���H|��dz���Y�
jr��T>7�0���s#����PS'q�t/N.���|�Y��S�.�ŋ>�܏]�����2�s��M~7(:	���=kO��XU(���cgb�9BW+�=���w_�����^}�u��r��q�V����h�g��[�p���e�9&�+�5em�}�vlU����;�V��'1�!G]��m�[�+6��n�9׬+r�9�W��P����?�O�S=&�R��Ge`��]DZ�!�pz�q�m���~�B����;l#U��=�n��Hq�޴{���pT���.�����s�$
�By�f�������(�\���S0���u�F��n��12z;gC����4OGLdC��I�ݬ��
�xMH\O)�����V�wO�C�=^�����޹�f���
Wu��*�d_ޞ�����{�9ʱ1�������HWΣ�ش�GOe��Sn���뇑���|}>� P����!l�<uT/&A��v���{(�o���S���D/u�#3�n9{*�|���bZ�
���3�I�ο؉=:GG� ���rǯ��z�O<�7�bz'��~�W�n2g�1~r<�gzdk�������̣O��@ⓙ�����fT{yz�6�>%�{']TE���� ccC�(���̋x��UB�a�3��Ḟ����S�]j!<ۅ�QF��H�6˘���Y6���w���L�9xdvL�8K�Ն���M�[�:����Vq�=V2�����o�e��w��ۺ�Rd���#2�c
�uc�S�u������х��0�V�,�/v6��]�W�ߩz�>5�EB����8΋�S\o�3m�C=wy����y�ֳX�H֮w&-�٬�(K��+�5#�׊��Zs�#�S������ډX��f�_��� ��@��@{�L�L���۞��G!�����wU���c���,Kq`��W}U�Q܈wMt΀��+����yt���L6�6���=Ւ�w4+��9\��J�o�Ke�8:-[�3��]E�x���LJgr:62U-��w�<x)k�]�;b0/ߴ{�R�t>�����i(�#����d[�RX���\�|`��qv�_u�`qm�����>���	�4��X{���"gԦ<vu9��{�O&���KF��;v���5��z�R�OŠs�C���7��wc*!O�x�>����q������7��y���%�Ԫ����O}�Wq�=��&}j�'���zX��P�)t�5��
j�q�n�9���dy�/n��}���ڒ��3A�ȕ�\<���׋�3Q�|UT��d���ƾ"�'�Lgc��5F�E_ |z��Gexۂv�A?��У�6�~>W��ڵ�}��^R�ο�>��c��ﺂ;/#�,^9��3��~�G�l�
��^��F��?Vu����m<P~?,w�e}]�λ�1�[�?RZ,�c܅���g�Y�g�8�J������'���}�m���e��8��;���+x��@��r�Hu�	�v:";�e��������p��<CfΧ�s;�8(��]���c�v��R�M\i��%Y��g���b���練.2���^��%Ό�u;�[/:`Z�{ӑ�*&���~�����$-�O�J��l��^݋���n��T������H{$vl����_��u�o�,�~�:�Q��:x_��^��V[��T6�Ԏ�ɟ3�@MDmHc׽V*�LMÞ��Θ�O�-o.�ˎ��-�]<�<��H�=�:�������Yq�S7�<%��Պ�ҙ[W��}G2�ݱ��L'^:����dr�+;h
wi��q\�
�~��M�7�e�͹���O6PS�����nߧ�?��W�CN�������\g��
�r�+db�,�J�a�C_�$=tj�������GV�Vq;�*1z����_w_\ug�WIc�gcӴ܎����O#
�z����<��aL���bp�)fևL����ҧ�"��D��7#�'���\�@�p����Gxe��<�x0ܴ}�	c������|�w�;��̂9%��F�@��n�EPǵ+7���9�Sq�=�T��˭9�/���a����(��烖<TW���5�ʆ�'b�`Ṵ̋�Q��|������rg�P�1����,���@K�xSL�n�o�?P�s��c�����Z_$,�X�2��t_n�L��)��#�.�$��M|��q�7(ɸ�n�%v��<n�_9;{[�r��wDTe��W	D�r���h�~���u�v��� _�~��[�����Q�#��\wѷ@u�ѓ��ӄ�4�f��?9�o�ì�M�Mk�0^fH姹�x�@����*9�t��tx�s5ZϽ׷��=>�5�c�d���ѹk7�Ʊ����OLb�ƾj��1r����ط�O�w*��Ϣ}^���>�D�����ח`�1�,�|�z�]q��5Pw��]�=�G��P�u�9E��}���j^����!$o��Ղ��C�A���2=�q����)�@���[NOv͌��ެkW�m����Y�[��ؖ����n��:\a�/e+7r��k���]��q����<��{/�g_+����4�ڲ�`�=�'�	ӛԇ����1��O��>�~.gI�ޠ7F�w�����t�cĚ'ǯ�y]1�r9����Q��ޢp`+c��
���73�1q�<���n�h�1���,����Ŭޝ>�b���K��/�}�C���G�����Ȝ��������������/T��+U�C~>�Ҽh%ѴŊ��|[/�C�W�,��wEu��.�z�9���F����\rd�SOP�#}w+�ܤ�2���a4#�`��ֲ�o����+&j�����w�4��չ�tv.��5�5
3cNjz�զNR���u9s�nZ��jg
�qm�D`���9�V����=�۰�o. ɻ����&8�s�FzI9�8;n>�/���n=��eת�]*�X&��J�}	�br�F������x�yr���d�U���m5H\ju̯}�Z6����������_fǼA�#��g���Z�Y���6�K}�	�\�f�x5q�z����':9�{�N^1=�<�g��n����.�;R7
���n��{9�4<w��x�j}^�|U��;�W3;���;b��r��z's[[���������\�Q+��`@l��q�����.��2'�E��cFJ�B�Y��R���v����zMî��z�y3�G�Q�=t��n��E�I��}�]�a��\���m{�C�S�=zW��Tul�)��.�'�s ts�Y�ȴ����Ջk��ݺ��������t�t��9�u{_��M�#�1�Ҥ��c* Q�	�
E� �s�-��#�����X�1��&�;x��K9���%�y��Ю넩���'���>8f*63�Q�������ݺ�+��U	;�َ��[뇑���|};�����&���~d���-^E���(��t��Q�^��܁�ۢ��훖���*x��=V�Pz�����O���ΛX6�Sl_7�a��ܤ��n>�/; ��38�mc�9zq�Iĩ弾啚.�
����^�3`�dI�=Ԝ��ǣuʜ���2��Ú�v�a�����(W`�B�G"|d�����UӦ�7Iz���Sl��whouτ�gmΛ����ӓ�8<�+���W�n#&}��'ޭ<+�/g0�S�##��P<����{�r#�޸���8<`{�g��*�H�4
�)p袷K��O/$��3�o&y�����b�5LM��*U��k�yObe��Z�o�����M�I�[7��w�/�a�d�VL��#j�f�]`��e��K���8u�Ǫr:�Y}w�{�\����]�T+����UǠU�z���L�,4}G�q��7���~t����隗Z�f�T�j�Y�;���d9�<_�������9<�Y��~�4�����f�K\�JlH�5r��z��Uk^����y�C��k��{)���q�L�T�î�Z�BzH�r�*���N���uC��v�����.��� <�%��.=1:���ד;/!{�mzl��j+D� �A�����[���V�Ly�*T9��r�3溈
��D��98l���s�/n�����T�~��y���@�2��<*!zi=!t�*�[�d � �o�tN]�ʫ�*�G�y`���Ȫ��xﲐ6����`yb.N�[WuDu+��P��F]�ikSÍ=�%{�-�b�Z��JZ�2%lV@�ө֣�e���'@*�ws��Q<0,��lv#j��3-]o�u�#�T�u���;E��+�*���J�B�jD��������̨����Y�W���ܥ$�o�<�_�,G+��r��`p��1|r�y�=♃�{�t���7Z�i��=�O�
��R&���ۓ4;}/޸y�t��~&}0���cϴ͝��v�6�G���U�㧾���9���U����]���u���,Ƀ�U�)���R���E�3y޽�nVN��}���Tm����Ӽo��w��W���;��O��J_�~�i����Uq$$��j����0Ь/�=P
��i�逽/�.9eG������N��OH�����r���V�p�g�غ�_�����xd:�"?I�� �Z��N7\�b���o�錛�����
�W��U��g�����1�}��ȸɟq� &�jC�ޫ��%�����M��������uo�����BXW�vЧ%����*1�dN�ܙ��̰�]X��g�M���w3�:׵�>��S��[V�U��K*�;v���u\�*/��Nv0�o�+�C5GT/a�~�&wgyY����[�x�+NwOi�W�� ��gr<�f�] �'m��x��_W�i�_���\�N��Ɠ���w�UN�_M����z��2�edR���6�������r:��\3���n���ڰ'v�\LD�n��V�Of�$l��8(Vn5�n�[g�=ԛ�cX�,�}�K�/: �����C�"]��}�#��n�ȇ��k*dyu�saS��u�w�Evy=��"�
Q�`��vԝ]@�&4�\����ֱ��1hӝ�^#��Qa���oMtއQ��<�#�{����㠐b=
��0�B,�+v�S-w5aʔ�_ױ���Z�Kaa�.��!�u����ْ����ۺǄ��)��#� ����G�&�v`��B���z���R�
�q�Y��f}�GjV։F�r�]�gHa�V�����S�Ȼ��-�=��5�f�k�ӱ���t{/����N�+͜��.�*b�1�.�%擿nrO���:��/ei^�������{�|��).�U�9�T�<���Yv{ F'YN�j��f�pGx�é��XZ��r�YS��grc��V����n��A��H�supQa��W��#@�x��#������Uobt����Oo#Y��3ms٧���R����;�ި�í�O8��ό���ܡvo��{B�a�T&LG7��s�t���s������b�>����A�wq*��]u����t:����by��ae8��X�[9]�V3C�����T�k��`P�AS���f��5
��U[�h� .���8>zh�Wx�x��^����	�S9]�|�M��>(�ӝ�m�d�ua�k�-��\��ٶ��,�]��e�eT���Y�k���J{.Z��J����N����	�d��Y�`�Bc��&i�!>$摐m2	H�u�<�a�+1�{Z�U5v϶>�Q�c�/��g)u�����M�^��.�����
�ș�x�kSU��>5lR0�g[����[����ˤ2���1u^j#����bf�n� �uo �ɻ��&����L���!GzEt����y��u��� ��L�K-���z��W����s����������}hM���اYV�#�y�tY��IJ�x����3��T+Z�U𾋨���v1�\�f6�hX�.���{ePƎT�Ė�����.+�ZH.�/q?'��m��o;o��n7��L�8rXt�p��F\Q��ڒҍ�\fna[�����_	6˕�>�#c�fu�5Pj<8��\���)3y�}��7�x����Vr�����J�q\��ita\��^`�M+��k��|;&�ݜ�K$쾄�n5�I;�R:���zA�n��U��s�Å���������;���c���/�R��M��SE�mt��&��ԙ� f�Ն�f�b����+[wc�e�p����mT�ȥ�",�2f�
<����6���:/UZ�o���%�%_tz�Io-60��RVJv�U��2 ��mØ*�4���L<EBԂ0��Gh��!��U��;U�������v�H|x����>�|y�b�AUb�
V����U������im�{�S^���`��B��6DsX�H5���<�A[�QD�j��h"*�+�&Q!ETTr[B���R�eE�
 �¢�b�E3
�e���+	l��F�J��j�R�Qb%��+3KB��҃�hťFڢ��-��,�"��+J�E"�D�k-�iyeUbŮp�PY����U�1E��
��*gjd�b���Ar]k"�m����ZS0��"�®�bְ�A�Q`((-e�k�Z��Rą�Ȫ�<�""����D9h#
�-,m��L�J�ł �$E�$\ɝh�V�V*�+U�TD[j$m
�V������E"1E̬Aa���ikT��V�
�ҩX�'Ň�5�*�Z���>����38ŧ_u�<�l���v��@��x头�L���M�a�9\��bt�D��:C���?��꾭{]6����(O�J��&è�[�.<���20�WT>����0[5ޥ`wM�Tn� ��<���j�������Nx��6��Ke_ٵ���i�p�t����}N�Gt�[C ��hR��k׳-X���(N����׃�G��;vt1���nO��n��
V��ʛ�Ò�W�|���xT��c�����2�ck1�+���a��o	�K�H�V#����ѓ��_mm=[9}�HS���`W�3��S%��0�~÷���F��?@���S+v9�E*����{R�ѽʍ�����l2�
�y]&UI��5ZϽ{z?a�*^�t�������=C?n��C2���T*B�=1Q�O���v3�}�?ed[�'�;�[���_�d0������(~�����:�ޮv�ㅩ�c�=;��co#��EF����-_\�,��o�7���k�����k���f���l�vO �.Olv�Qu����"bT.��jn����[���Ƚ������徆g��k� ������a�3n�W:'�~<��l����齅+v������*>����#�>��#V�f/��lJ�g	�ԫhQRw>���5�q�I�"8�%����hǡ�����ܷ�0���o%�8�"��VQ��&۞7o�ݚ�D����ch˫v73p�!�nU���/��iȮgq+[Z��d�8YK�us}�T<^�R���U}����~�?ǡ����oG�%ʮ~�s����S<@�F;܉�}ӿx�	�3?[�=�~o���
�r�8���\B�Z��T��7�V�}�E�������+":� ����7�>sE�FUQ�fu�N��\F��H�r���|nZ��dwX�;h
f��Rr߀�
|3X1�B��W���He��;��c	�Z�f�wv�����ϼ��)L=G(�;��ȡ d/S�q#[�U���s���p��__Wx�yr���Ke\d��o��!q�y�Hý����pY�Q�/_*�i���i����e��UR0z'_���h��O���,.;���^�y����}���/jָ'���=���e��*��(�#��~���eؿ����>7�0�}?as'`�R�7�f�_��R�W����;,��uNH]'���)�������~�y��c�4�-}Mw�(�z���G�oT;U�tl>.MC����Q]��"��٣�[�{n���t�g��FB^ы��rhwl�;��P�zzTǏH]7*z\q���I�*��`���։^YۈH0���d_r�C�v,�CkEgf9:���%P�KM�h�̾�L�)~����ǽ���?��QlU�긡<��Q�³&.t���밆ގn�|7���%�ƹ�=k�;p��|������f�l�����m�<~��i��,��;�Ҽpl��O�U�p�B�%�R:�����h��9P �}6���	���
�q�6�=#���ʝɺ��9^�����޹�f���
Wu�Y�\O�3;�F��f�}9�R_���S�b���Yy�W{o�?~�k�	�f�����{�ki�'�U�£/����yw�_���҈腷lR9ݕ�y��ޛ�;��q��e�u�Gg�+�q���Mgh�u�4���mmk������9�E�u�Y�Y^{�oE���F���Y]`e}����#f�
ݤg��F������{#�7�B��\	R�L�w=�9�W{��~�g<|Ke�ux>�9�P���Yd��fE���;��l�{�{,K�t��U{q��eX�s���]��Q���G^ڜ�ӝw�+�t�d_�d�f�&X]�V7��}�M�[�;�^����k$�LY��ד�ߪ�u��|ǟ�
S�PT�(���`_�r��ɖ9s�딍.1����sw<�T�K��Jh��ކ��}|1NQe�ܯ�e��r�\��@��}3y0ڞU�j�_�ۆRc��v��C.'*'2�=`����3w�����&�Gn�K���p���]v�|�vՉ�,����,��J|q4�1��d�e�kP"�}�N��F����VF���`�a��w�����L��R��l%���^#��R눨��6J��3J�|��/�G�hץBO^W��U���h�}�>���=E8�7�|T�3�:���W(�}�=����E�����Z|'��j��}=�c�i(�#�Y�dT<�tP��^����|��nڛyW��@�|���U�>��Tn֎���)�.x��n�Ͻ댨y5�@[�{o�}*�)/pQ��<'�w#�`xVgz��O��b�'���5�.�ڞ	5��/$\�w�z�uX�4m8{}ƠW�TR�fcݞ������x���?�������~E�W���iD���#j�љ�A~�9�T����q&hv���\?d����f������I�)=aGm����/�w:�f�=�����^��X�^5"iu/NEV���˿'�^d�J�������~>������\;Fs�}'���}���zN�؉�=Om��(m;@B�^���yES��f���t�)������s=�0/䩾�ۘ~�e͘�}�/Ȧu�͚�����Vgާ`eDgU�C>�Nٿ9�d�͖ I�p�N�K��X7vF)3fG��k�V����������ޥ������Vמ�����9��������n��x�A�Ȥah� �.
ʽf+Õ�����\%,�}@�S�@��y��Τv<y՚��^;���[rgS3OgN�87P(���[Ԏ���*�K����������@<��WeF7�"�g�n3��6�1�ޫ�S�r����i������Յ�	�� ǐ:7�;�T��*p2�j,F7쉸�)�����̰�LI���<���z�G)�+}}lp���WὒY��mN�`=�W8_?d�&Ӕ{:qW({�ZV|��O1Z���5:�aߠ>+��;���W�B�)U�������Wt<~��KœY�յ���=�@ttޔ'2�M��wLo�[ONG��������,g�%��l�����[�a�S�Vp�Oa��6�	��e\Fmhw3�t_�uiR���;"D�(�.���'��In�Юb��;n2ݕc�������	�Uc��~�b'8�O-7�~����n��)�{n����n�q\��d�9뉏Tf?ea�%����0����xU���-�v��v���G�O};Lt�u�q΀w�*��!�S�V�RU�2r!��jgPܱܶ^�Hn�Z<�L*��+������r9�v��.f�Y�W�Þ-�1��0��F/�F��Ȱ�\�k%`��Y�f:X�x�)���[}��z�癭�%���(�3��]>�mCY\{��{���S����K�����V��J�v����2�a5����{ϖ���nb���[��0�]�e���
v��(�^�Z�{�I����c�gÃR&9)����>��wý�(
���3#��gϪyk���U��b�~��=�=K�g����:�z�=Q�������^5q�ׂ6�<̘����(����U"T���\��Ek���?g�~�`L)�@���l�=��h���Xsk�X���=�Ղ�?ZH�9藷�׷#�J��y�� g�����\ۺ�Un)Ǳ����L�x�s������Y����?k�;3�.��U�f?�X�_x~�����嬹p~��R���W|�@Lv�,�Þf������H_{�Cy�O^����mdIF��h��̫�[Ƨn㚹�s:�sL��z�R<��9%�uj���G���h
f�e0���a��L+�f�������M��a��1��,֞�2e�ٳa���,V7[�::])����f5���K �j�=F�Y}>�����?.2�q��%���̨jP�=�����-R2����^�����g��F����ǌ�s}2�v���"�dU��*U���*������&��G�`{�J���;sn�V6�
�B5pꏖ|`[R��3D��z޾��)7����]\��ca�9�Z�z8x�%�)wRw�V�kYc��v�/���-�H�,���5����cȝay]�Rf�ú$��2�c�s҅Lt��$�S�{T^�H���麼(�	w+¢��ȷ��p�#�Csp}$'��G\����{0g��S��T>+÷:.E����?�yv�偳hi�a�*އ�J����������"��T��u,\A�����=Q}�ᝃ6&��5���L���{Q�>�F���ɷ]@+���O*��S$4v].;�=��s��7�^�y�l��JC8��/d��=���b�P�zT�F�P���<q���t�/�Y9=W������uu�Q>�I���y�V,�������?�2|!��}!tک��满�^yY��Ӱ IuטkN�!��o@2:=�R���������#ޮ�z�A���1�UOJ�Y>���(�pnj�{A���8N�zMƚ��^Oe��{Y�0�zٮ_5���=oi� rS���r1WO��N����d�#����7�^�q���s�S���D/��Ԍ��܎����=�}}T2�s�Y�7\������f���p|_�*����QvH�=���w�ޮ���CX�����k��8���=�;���7����p%K]2.�y�Gw�q���Q~8Ke��j�<F)��j�o�O�ڀoNV�zc��)�C�PW��^Q&"n�������u��	��Ҏ�)X�Y�bd5�0�,�Z���v2�_���z������;6�3�r���>�zIW5�3���ݜ��VZʷ\���o���+Y��;�3�\x%�P�VY~{�vFTFuv�>f�&y��!��mp�K�[�)�N�rQ\���f����>1]n.���s���E�~2/&S7�d��h6|��M�Z]ݚd;4���\u�Yhhȃ�z�s��f�KꚌ���X�)��&Xh��s��h�˃��\�צ�]{Ig���;θrޮWW�Ye� '+�� ��(��D�Y�&�L�pc�JO�g�^6ל�L�^zzʇ�)/O3o���=]%ߌ��񃬹���v����4�دO}�\9��>��7�����T#�zxw���1:{<n�[�rP���f]�0��Ta����nv��
�U ���~2�^>�,un֎���)���Nz���&-��pe������,���z��M�%��£1����X�S���l�ҝ�ù���l���֍�4�/w�]	{ łj�O#_uU�.[^&:��N����
��'�M+�K�;�=�w�k�:u�5A���@Ts��q��W&hv�*��WI��~&d胾���g�l�9];Y-η�N��\��{��;���a���먽�t��χ>	���=Os7c�<�;�����j�F���_[|���#nrR77�[OiՃ���oz��f��(.e�9O�s�sW4��������m���e�#��C�Q��T�n�}Gi�y�o��{%oo�'J��uS��t�x�uS��X�BH�C}fKӑ;<6�s���3�����*7;wš��a��@N�\u��� y��*#��®z�^������vy���Nnk�+�oT���->1��n���N
������T�F�gL�O�=F2^v�ኋ�0�u�M�<��f�o�GR=�'�}]`ec���#�;f��=�;=��	�p�N�K��W����yצ���s�ګ��h��Y���>�>�+")�5�\��&}�8����1��X3h����:��u[x�OFMw����YO���� �dK�.p2��� ��o���w&x.*o�c�� yp�Ps��zg%RW�<��w;�q\W��hp���+�Ϸ�E��GmN˦��s�TE��@�
�R���&=�/�{�d�Ќ�ۘo]+8�}��n__ �e�lG� ��K���f�T�"�����և�^߀+ׅg�8�z�ƻ$�3��-��뇃r�� ,B5�O[�w:<���6{�P]T���?m�q<ʸ�6�;���:.N�7�@��h������`�Ps/��l�,�z_~���է��M;r��0�1�`4�^��kk���r�e�[��j�.\�%��mm�(8�J�{<k��7����U�#4%��Y��iV�\z�"�{��B��[+Lzi�ў�@�Re�<n�f�ay�hl�U����	!P��%��%�&N۳�~�ʴ{�n���jd��U��^3�}�]�T=�&���ր�+�&+����Gt� oz_޸������.��%>��!)�����˄EM��JG!ݳ\o��æ�*� �]��@Z�,��3aqݩ�^e�9�a�����_{ئ�)��U�G�'�j��u�t���xߗP¤����˩<t{隤ϯ������!�sv���!W��ޮQ�<fkǇ)!L��}��CU\;!��+��(�!J��{n/��63�ߦTV�s��J�nO��/=>N��g}L	���T]�����o�U���kk�K��޷�;[�Fy����7�r$�\:ێ���:��>�/�T�~Ur~ o�^����q��d��hE/���v��пVQ���VY��W����h3�����y5�A�� yc���Oׇ:�k�7]%��;9V39ʞ�F�ë��C!�>�u�Ɨ20_��{�73�i(3Ӝ��q���tcR.��ۺ��r;��
�T��e�s�[�]�>�5��yU~��ʱmq�<9��K��ת����u)�뷻�t�{yo��џ+�*�\��iy2�<�G�����;W�)һR����1\�-�T�"��V9巁T�s�s��	S2��M^�ާ�����FS�s����>�$;2*�>���R���;t�ZڹʶN��)/la�C�^�6�SoS�����]��-�"�oe�
4;;C$��	SBrɔ7��eCt�d�����:R��)�u�]�Z۷�oR���kҪ��w'�q@(�h�v�oM(������5R0>�Y�[��tΊ���U�WV�!��
�D�(�R��+267�S0��]�[WI͠Q�@k7x�#W��ԩiȹ���R���Ii`V����zi+ݮ�[�C}�M!�h�V�Rp̽Į<V�<�@U���׽�1����M���Ƌ�wKl%Xa��de<�6J�fS�Gp���v8���I4���	�Sk/Viju�	S}yl&.���v�b��W�gB�݅��=��X�J���,	���y=��:�_gw$2P*�!-B��]i��Ƭ�D5\��7m�'��1;g]�b�k\�2�����s�m}r$����7r��M��zM�wn.���p���5Z<7�=OF� {pD��6t�j������n�o\�����f����S͆٠lY��\��"�1X����M7I&�wzoT�e�J�T�oKy4�d��hV=��l��iݜ�34�f�������v�\����\��'8[*7�0
���mD�$v�[8�{�30o
��t�-��j��b��2�2Ft4%n��Z��Of������Àw=qr.u��铈�+tD���+�H:G0z�o�:��0<n�Yuv���U��ӂ�߈_:8�1b�-�Vm�.�b�Ěrv604{�_Bm�\�Q�#Ef^q{�n�-���yA&ʫ0&�Oz�z���8Ig��鍮�:m�apE�d���TGn_ݜ��1��ս���r�!���f�7I��]��v�3['T͕v1�
��I&Nj�q�ӠM��e����j Qx�ρX�ۻ��r�3{�&�Jf%�0��-�!=�B�N�e�_j��腣HO�$n��3f��]�`����'��+2<K����YΕvqB�S���e�:�1�Rq��j�*���o���~j�R"��W_&����JK��}�ƚ�,�S_i7C�r��7w������u��HPs���D>����vh��&�ղQt*R�(�-4�^抚}��6�3�X/nf��牞W��%���	�!����%/3@���$��S5�gX]�`Ӹ�q��H�>�j��0�v�.��hg鎖r�Q���u5m��Z@ĬI'�!�	�Fg�:�ƷyN���w>�Z��őG�EI�q�bN���4r�ī��}]0d�#�r)�����u� �C9�ȯV&�����ρ���;j��{����I�>s��d�VP���K�^;�~��
�TJ���D����Q+QVT�DF(,QTQ`*�����[�e@�[��,�����*T,AJ��,PEA@��e-Q���ְ��`���@��0QI�A4v�噙"��H��.Ni�Cb�`�X)3U�P��8�g)*��Zлl����r&m,L����(��XAA`��X*��AH�VIP���X�jTa�(�5���!QQ"�"1�X��R[W["��UY�*���q�"��Ur�q
��TR����59h�X��+YXT�IU�q���b���AH�QJ*)22���(�YmXE���P�,�k%v�@��-�PP�e@YY��#lE��q
�1k9��"��X%��
VX�F/5��md��W�Qj��ʅj;E�4�*h�Yeq����U]�}G@u1��]V�ڔ�%�K���.Fd[#n�vbWY�ýч�{�m��t�@��o�ׁw(��������?eY��ؠ���]��y9Ts率��=�r��v�H�5�˓�}�}b�2ɴ��3��2yݰ*����H��2���f�w��+�����V��BcyRU�x�L{ؑe+�{ƌ_F��f����={O���͖�١��j��yt���l��=W���7׹	V]�P �k��@��T�
�j��-ܞd�+��=�;����b�Vyy,�~G�����}n�\>����2�>��ι���w�� ��+E���+��u+}�N�^�ꎸ�Wq�=>[�85�vY�-�$T��Ō0u�eH6�1�S�#�hY��^���#�s�^�{j:�}T����q��"�yU�E��>�a�f���9��a����x_c9��Tf;��>�XʅB��l�)�����H��U ��'�t�׹�۽nHB{M�3U�{�;�����^s��{\=P��b�R:�������z���;#�t��X���0��f��� 7/���7I����������΃5�8*���������E��+�#h��pv��]1���h�>�%Y�u��J6��v2��p�Ah�I�U��:�f��}���v�'D�w!��P����4X���e���Ν��$�ޥ]���rZ�ՠ��qk�;-�}Mӝ����6��Ҳ���{�����L��ꇸ�2-5"iu}ӵ�b=^��Ȧ�X4ǿ	�Q�ٛ����qe��ր�i�	�"���Oۜ��ެ�N�gU�m�Ԍ��܎���f,�K��z}����ܿ��<�������o��놳��o��:n9����8<�z���=���/qn�Q�X��~3y3�1yH��#�z�⦺de�7��\<��(�lyW{�Ovf�U��%lj��:��-ǀ��"e����K<e�����H=���b�MS;��o��tL�4��ҥ康�k��}A�튦\�E���~���y2��ɖl�l��u�a�C��`uB���v����G�΄vt1���>��:���\z�e�˔����Y+�.;�}S��㺳��i�F���Lx/����B����!�Q�,��
懎��
'�r7''�g�y�`徙�\������_�������`x�<�� 4o�LKg{#Z�aѥK�u����@�hމ�ρ�xM�����������=��c���ge�_<�tPY'2z�Y+���I�/�e�ff3����7���t/�0�_�{y�x�iɌnJ]h�ӫ��)������ş/s����k�{n���/X�(���P��iV�1����yDҭWݣhv�c�K�]o���cv!�md̆����]�mP�S��Wwl6�s���\;���փ���A�?̛���]�T��n�ƾݝj�n�.!�;5�W �Wr�/����Q��͜�I�i�A��{�I��ƾ,N�^�����<=�,e)�؟�w�?KwKڹb����gj��y���{ ��P=�<��j�_�i�_�-x7�<��57��q;�훟��Q�UT֠�ԕ�ܤѨ�t�©�㺽`[���td�	gb_�p�#ޮ��;C�d4�u�ۘ�Nǻ��ɞu�P�鋅2x����<{�pv�9V9a��Q���Ump�l86]��_IÓ��綱_���xGz����G�}��p�� _����uV��Ub���4wL����߼���t�K�?��������prx�Y�9�,	�S�=�0/���9eG�8r�Duǜ^ܞ����h��RΖc^	��}�T�>Y�W��zxz����<�H��F� 'S�MoyJ�۾�;-v�ΉJ�ns��c�
ð���/�Q�5��ȼ��ΐ�ڐǡQ��ݍ���Z6�ݖ��_H�~�&����D.���r�Gm
sr�+������VL��LY�|#ܿ߶̄�=�
r�&m")nV��
�+�x3�'��, ^Г�o�)e�YE�%�'Iz0,�y?͟z�(8]��׃f��\��Uvx�ċ�|��^��'�����V��K��R-�u�oTL���'d⯛�t:�ƛ2�+^�딯�r�Gqt��|�XZ懡t�V�-�:mV
�oPe\G%`O�{�\h��j����,���fs��*G2���l�F�9s޻Xn<_�;��۫��eK;� :'�*�؍}Y#�ؽu��s�5Qw�z��wC�=��/�G��d�VT���V������=�ާ[��#w3��-�״t3i^�@=�vZ6=m���K����g��]:T���1��5~� �Lސ����9����gD_�r$\5L�?<�>���������7-z}�X���,?������u���AS���o8��\`�t���t9��}$.�ȏ\Lz������]�$�v*hV���5
��D��͊B�e.x9�;\ W�vX_<�)UU�q��}t�s��٦'�+�{�Eo({���{*��Ѩ] .7
���r����WI��WG���	�]�;����W4s���Y�z}�j=/���c�
�CJfzc�8�U\9��Npx*�P/Ǘ�lү�|p���'�;�[lnDO�~�=>����3_z�=Q��P*1��mw��'a�f̍�=��:��9[TO���)L�D;ge�Vڔ 0
2ԏ�[�����'7��X6�k(�G�3)���n��|Ȳ�d�̇���Tu�����vo"��\���n���I	���Z|�
%ܣ��t쭶����.��ݓ���70s����͑u�~V6h5����~�k�A�־o5����a�뼮z|.�G���y"�]��p���'���J�M��ݓc��V���>/j�Fu���e+7� {���8����6��su��{@����m��n�K�u��o���ߨ�܈��9] f:ۉ�
��Z<}QO=���N�@�{fX��oP�&g"��y����k��}����.�<
���1z|rw$�Ua����dM��>s��q�2��H�r���|nZ��vQ㵅�1��a�����L�c=|����9���U�~"�m.#&Z=�6��c�;�����<w*���S�˼����j�Uw+�a�='\� �B����@��\f�[*�ls)�@[C�����3��eL׷}��M�u);�w�0�.��ܨ��UH������8x51�sƻ������Yץ���h�u�����0L;���3��S�����\�W���e�򺭴�[�1��8�<��W}
��{�b}\���w[�8<�)̹#zO;��)�+8K�.8״�2�͛}1�=/���������}mm���Z�Y}a���,K���.�.7G�����eYds���ԩ��^������)ޒކ�7�8�a�ۡyñr�k�9rU����\�'PN����{���@)ou��ǩ�{��n7������������9�/omG\O���L�.NDK��G:"a�]�#sѕ�����z6�#�Xz
��x���M�^ѡq��@/*�g�L!t�ҧ�t�����'�%vj�'Μ��ӷ�OyWm	h�3����t����s��q����,b���8�����r�<���=��u����n ��jE7�eN��u��0�'�Tk�},p����q�Oo�skW�v��,�ΤO_uP�s�b�xԉ���������=lוS[�N�CN�Nz�s#�;{9΍OB� �c!L�ki���s�}���s�M�;��p�jF���7S0\���̟yE߼�;���À�>t�.��.!���,�
�eN���#t�>.B����"����ջ#z�Xc�V�WXY�zf�ɟ)�q������J�g�E�=�=�*=�h)y�=��5��ۦx���|N����������"�ɟ3q�<��C��p�I�b_Px:�@�����}Yć���U��r�(Ư��S7���\�G]���ȼ�L�L��f�g'�v�����ӧ#ٲ}y�����d�%;���ҽ���,u�}d�}���Sq��,e���铂�ֲkOF��X�;�l|w$啌_CYҬ�/xoVk��ƌ�[V�Qv �z��A����جQ:"�sX4]e�D�=��V�(m�ն�t�ɂ�o�"��J��M�_;����pV�q��u
sp�XT�dE�z��)����rz %���ޝ�Mo�q:�E��9H����/���R������@?N¹��s1[��;sA�^Փ>p:��7���f�C��RF�^�g=�>}n�Ϗeu�2e��M}<��}��җ������9��x�V�L�+엦��z�\um�8;IF�U��1���#jR�,�^ZϳyQ��bu�LJ�����_��n���_n֎��R���Ɋ��Ù�;+�6w^�S�%쉭ɥD�By<%���`xVc���s�wc1O�������AS�n;c�Y��w�yˡ.t0u� �gM���Q�73U���c���}��z��:8Uea��ui�v�BP��&�|�@])��>�>�&�uȻwG� ��9+޸q]�>����'ׇ�9�]�{�/��}�f��pJfx��P�>�𖦇+3"R�<^�����j*�����Ng1��_��O��~=�ɨ�`O�]q�d{��������UϾ�.��;���j�U��/V�Ne�N���H-���w�!ŀ���r�0�5`e&���|xn�.��,�7����shAu�>r��� |���].�`̺A���x�XJ�S�����j�b�j��Â���i.;U�/㇍O�Vb��[�OT���pz�R�Uf�l�J�C�[l{=U�=���~r=ӡ����G��j�o���\����g=x��d�F.���ϖ	��Ԝ)dS�2�����d��<�H��m0��(�H�
�_���|0��=	SҲ#�`���:a�����
�]��_cyr/&}��3��)���3u^9��ҭk#Et?U���W�r*{ǯ��q�
�CWnص9'*����"f��\���w]�����j�?YD�k=2ø�ub�Jeo��/���~��,��Z.�eh�嫋Y����Ms���k��2�㑷0޺Vw�/�Gѽ=���2��ݨh ]�j/|��SZ�wxjVl��}9@sȪ��>W�a�xN�Ke\d�z�`��o�~j���_��ȰZ_����-៪o���:��+:�yw�׉�d�,Y��C�;>Ń�%�8y>�{�yf����"��/��ޯ�7���P�2�+����wCE�=޼�h��� �"=�7��Z}3���{�--K��:v_����w�<�#�雁|�s���!v�z�c�����+��4�2$ɒZ^�ep�X�����ͫ��S+�v�*~�st�b��+���鄳Dlx����\�AS���ӆ6{ɾm��ppf�ԥ�����"p���+6�o����4�b���n"�k���EMj�/�sp��z�v�<ڹ���/ڃ��+�߫޼�{�7��烐��_e�_<��.�U}=5aq^���(q��J��gR'��~�2k��Zp��H0���4it��ڮ�9��3�y]&Mّ�>�β�݃%Z�>�W6	��9�{z�i�<0̨�Ƣ	��=1��Oj��Nw��&�A�~'�ϧ��\�d����ظk�grv�m��{ǳ���M�N�5�`Lmu��!��A�W�뵠#C�e�Q���cݧg�����4���@�/���k�����T�W�����9i������o'������TyDt����|��s�[�OH�뗷umCQ�g�������
��)8	[8 ���)��n�KȎu��n;|+Cy'O�z�<T�WHޭ�L;��=��=���3�|:e}�<=� z��ۺ��s���vO��d��@g2.�'��h��������ˉ�q�ld�'9e��걣��E�\w�V�=7<$�o8.gn|������f�΀�7YL9�W~����.2m.2e�ٳa��b�7;��إ�|�n���i�PZ1�����+�T���^`����;�Mn�����BG�^O��˕��N��{v������3Gp����(I��uK;Ĭ�Ոc�+v��$:aF���V|P�Z-\5�_kNQ���&��ܔ�Z�䘳�o7;��;���'l��sPa���ڇ駍E�����]e� ?l+�Q��@���\f���ʿz�s8�����y"�$��]�&���ʛ;���øU�x��*{�Wt<.u���-�<� ��w�o�Ǯ�Q�c��Å����9��#�`xW���@��n���}$k�ι��U�4�Zٛ;��`ۜ�`
nr�=Q�k�ݨw򭾣q�:
�f�py�DO�꜑p���UOv��={�"���7� g_;�̈��9�5���u����_&��P
�����\�{��c׬�Šn���.�#�TG��t�ݩ6�ߤи�=�rc1P�~=*cOH��b>ٙ����)�I�Yj��Y��@΄n����d���L�:��=ޟ�Qs��{\=_)�Xg#�*<��_M�%6F8�6�h>�g� W<&�.'��j��=9����o��:�����ʥ��ٱK}�4w��.;j��q�����������؞\jEy�#�;�z��"��Er�bv\����F1����;7��
zxdB��"�m1<n;r�G�&ǣ��>Ϻ���?D}��ꟿ5.c��K����O�Z������v�]+��^��w�	��P���F��y��WwR.*��][$�b�o�V�h|���5u�9yԶM�:&��f%1I�*b��1���a��=��|Q�Ϝq��n�oK�����+��(/��{����9��pn��
鹓Q�v��͏i�������2���P��Si#Z���/����ܡN�{�8�I�+'M2��I����gg#�Q�Z����5Y�0gp�7lg �*y�o��{T*�RT��VX䢫�W�ԜF��{+g)�;i<7���˺���m�����W/BY�*�s�SL���rPǊ����v�b����*{ư����}�B�v⻂ޱ��\S
%�qs��:���j��� ùC>`�ܖ9H��Ӧ�{�� d�Yt�"�ܯ0*U�Pf��W;"�Ī_5�y`�S6�	-E���O��qc�,�v�Ϗb�x�V'|�R1s��md��ս,�U���'k��u u����k�z��e�4p�[8L#�Iuę���=�U�s2uᷫi2!��)��ê���^���`y�]���נIh0�;i�����O9M�k�+��pe��G@j+;����h��0��5S�#|�Jz�f�e�3��w����n�4�&�s�-y]�#\I���:��
a4�nήP,θ�Vf�����.��SA�Mm4HݬF�L��9r/Y|�����b�E�lW��R��3�&��t�����P����]#ڑ�_s�%����V�=z�g��{�s���҈�h�<mkU��˒�n%�ݛ{AS�z)�c8r�d�YRO�FvμT�����n*s¡�\�7�������'�WW^pC��e�ۖ�4eɰj���SMe8s2�7�;�m�0i�I�*��2��vN��L�N�C�eK�	�H�ʺ<{ż���5{��wn>8�.p 8�MMu	f�K��!�:+�/X�.�t�h����]^9�j��]�U��ү�v�����~
�-���J�PT���TC/m�3:e�١h��m�V|��:Vn����DT�%_J1)]&��\��w� �]�	�z)#.�����Žp�fh7�6��wH(sLac�t%�{H�&��	;�~�3�ܡ���jt��Y͘b�e>������Ka�77oh��:���p�;wR:��"Eg1��C!w�oޛX�K�b[�H�fG\�M�����|�S�l*m&lսN�!J�GLz���w7EKS�<����t�үv[X(�[*gdQ��m�u�m�nN*���-��"�ݿ��7�+"�,]���K�v�v�B��:�su�N����)�h.;f��1���W��m�:P��e��Wh
�VEa��X�Nj�f`[@̩dXeTb��fss`���i�1x�L�`d�i�QdY3�`�H�P�mm�K3*����^$R:�E"�6�3 f�J��Z&�Y3+*u�sI��(��"ŐX���b�Yy��8�F����*�"�5H��d��V���
������T2*���T�EDR���"�*��2'2�P�
(�ܦEҫNr�
�Tu(��aQ�]��V0Qd�I+38�<�R,s�I������Aa���YXd&b���ʐS�8�.¢��8�B��FC�X)�E���PU�*VT� �V�TX�AER -a
*T(�J� �G��Ԭ3��T��b�̇U���DAX�%@X)++ ���T�fd�]i�� )Db2%�0�Vs��=��Z��+�ܮPRI�Y(-I�ˮ���z�O*���'�uһ�c�sN5)��bU&��n�\�T=�ѻlҝ;oA������^`��Lz��K����՜F7\7�}�,y�z��7ޘ�3�S��F�:nx�g��b�z��n��iR�,��}�C<���}(/��]2�7��^�*)���-�{��J��9]ѫ�x���_Oz�
λ#+�t�ȸɟ3q�<��ِ��k��팏x��0��ǻ%˿&�����]{�+�ƨ�
��]��q�=T��/��)�ɖ{\�9�"K������k��n���بǵ�������8aX]��H�)԰������Xv�Ojʁ��7u�l.�N��m��R*5���cE�U��ϥVYe��d�9;�^�×�^�T��X�{��r���Ɇ��f�C�]I���Ͻ�>���c �WQp|��n�{��c�yO�aF����Y�|Ԍ���L�;/ME��
�����%�G��^��R�1�1[��v�����:�����C���W�~9XsAc�v�u������.y�ss�L�Q�D�e�Y�swm�{y=�PF?d��]DT%�g����0z3���9Ố%��~�������d��ב(���./����e	2�����뵈�����u�<������e�j���Gm��Q�O���2r��i7\�-����R�y�k}��vu��AA,�C��_Ka�ݭ��Y���Vgni|�yǷW�w;�2U�z�V�
wn)ڎ�r'Gr��q��>�8�\ �y�7�Q�=3U��^&:��J��j:W��Y�����QX;f���S�*¾]&�>�\T;�|�(
]�t&���L��;��m�z_e%�7/�y��MG��3Q��_+�b���_c� �޻��4+����[���u���RJN��c:�xA�U�r'޿��W��Ǉ�p={���@���x�v�xQ�'TO���s۷䏭����2w�'�P�����Ͻ>�q�#�7��0��=}0*��T��(��:��}�.7ý[=���_��8b���O�L7�� ����d:��y����e��s-��:u�ڴ� 	��'�K��U���1����D��Ĭ�p0�cyr.2g�i�^�Kpv�y_/ON��5r�z�Յ�X��u�=��l*9�P]�%�˜���.�ޏuT�[����{���?����ɟ�3��,?k������r���X/{�Yy�@Se{!ܻ�Fjm\�'�g=��*������m9����sna��k����=Ǽ\�S.������aBdvu`��f�I)Z��u�l��
�Uc�[�A�r��r?��0���y^L+���|�h��T�=�+:�v���:��f��yC.��Z݆�AOU0��:텞�w]�k�����y}����8|�O:o�ê53X��(I�xy�-������Ĺ���I�;ҟK=�����܊��A��t�n] �>Wt=q��G��l���s��(>~����WQ��՞��ހx��n7 l�,_�1-���G]�������m�y<ʸͭȅT���#׻����jx��� u}}o"E��\nx��7�P{����{��xܴ}�\��/6��{��V����Kw���O����w	���.!H��䑼�=q1��y�&�}N��w�6-:g��g��0����xW��H�x9ߊ� +��`S��-UUk�洁4mĀ��gq��=
=W�5��W��5��{NA/B�0�7����x�к@�}9`_bq9��~v����y��/��=�'@������O��DzX��c�P�u
d��>�<n����z�����P���As9@T~��Y�p�	����~؟W�{��q�2�L���&^��,��=z�<��p�t��Z���#���G���z�`^��k�_�Z��X/���A�W�o8���}^l�5�}����O_m`�}��s���}=#ܽ�8n3�n;���_���kr�݆MT4�^c�M,�Dn�ۏ�k}�Zs��*�?g�����n�ňA�Dc�rgL�5�@4bgE�j_o[jv)2��#yh�Uͩ��2�K�d��s�#O�!�C�u�AP�>�̔uBѪc{�z;��e 3���7�n����Y]���:=n����_��B	�5���-�=c:�dM�L����	�����ޠ%9L�ú��{�օ��Q�I��=�^��'z�nT����;^c��1���dϜ��L�s�i���P�<��8�_<�%�/tU��3�O��*㒰-����+�_S��M����G��mm1c�K��Tw��r?�|��EÁ�_�)���j�,�f7�'������=��@���\f�[*7�I�i���:6���д��Ljs�덟x�w_\p�+�y�!���U8�H��j�=~}�����*/�s>��2u�����2�KӺm9��>�X}n�_ϫ����2��B~�<=��y}V���F��=���6�}Y��{�g���A��;p��8r��W�Q��Z�Ͻ߇��E�ֵ�B��|���t�-u�d
�9�`����j;ģ�_%�H
���al;*���%{�s��]$l�����;荺���I�����2�P�u=Ja�㻲��Z���$/�P˫�4)g0�&����֢��
}����=M�h4���̮����]�{�3V�EXU�;����)9W���6<���}��q�t�C����-��Qw�;띃rWQ���9�v�0X����{�m�s���Fw8�[ѤY���G�c5����I6����?u{T����$���Ϧ������*��v��I�*���5Z��]�Ͻ>&�����M�o�Bt�%v1G#s�A��wOĜ�G�-�T���d���&�Wˤ~�t������oA�~3��]&~k�WB��z���X<)]��OQ�:�{�dgnh.^5"iu��շ�Gs}*hA�k�׭g�q�����O&p��>��� �^��3�Eƪ`�r�m���s�S��#8��U纯suN��˾#�z!VԌέ�J#ӕ��t8���M��g#�W�o���>�O?ld_'�x�B?z�,����V�W���`ƳL\y��v{]���Mt�'�t���o���u@�U��ݾ�y��4�Y-��8
ߺ쌨�O�ɟ3d�"�fC��V�)��/=��5~]�GG?S}t�NC�W���(�퉖T��\�]���ȿ�e34��N�R�r��Qֶiu�Xh�k����y����Q�w���%�D:���W�4q���Sjf��u�
üuγ��h�۞��F�\�;�{���}|2�^x�n}�;"�eo������7a�i�] �,ċ�2߅-	<�$�:M-vK�)+@��K�'d�۫:�����uE�y�H�ӼmP\�����j��MhvfZs,b�D�ۆ���v\ೕ�f�r�sX��x��F�JX�O2Xܝ���2/�_�c"��.����CM��ʆ�R* �^�g��A�0ﳱ�k�(FW�E�^&WKć�)+�� ��0_����']�fl�7=�o7jϫ�������X�y>��]���4𲹬�+�ʥE�1<�Ǧ%��=__u�`�a�s����ȥ^bۨ�Lf��~��5�w�=1ѓ�ʑǀk���}Vh�{�:L��~��b����s�w�rg�� B��S%q�u�n�H\�IB��4��N��[�d	4�@�TyM�f�����i`W��G�7����:�J�t������I�>������_*�B�4jH�Ү�q�r�uH���2wlyk�{+=m��w�)�7�C�OM/\nG�NMx�5�|j�1jd�}@7�U��^6�1��)61�^��ݟ�8od�m�����h���޸���ʞ=x~c��L���q֌� _�Q�v��=wbc����k�+�޼�nh�>������o��c�?��`xeVy���|��B�!~~����,�u�ΙS}+�=�*=W�d�x'|w�꓇�"����zxg�Ű������W�V9(f��f:�K����1�$�Aܹ޼��[�`zλS>��DFgwQ�V ;��6�j�ӳ����Ddf���������T5�c�)�|_0GQ��ˏrbT.�h.�[}$�o/W+x��[�stѤ���E�e���w�j�z� \�N�H.�}�%Ў�?�����1��؜�=��ܫ���(����=.yf��,��� ���:^Ԣ$��w�z-�3	��|�@]{R���X��5LM����޶�P��T�Ĺ���x���ɪ*E�~�S�p��7~��~j��L�L���ѳ,=sAq�w�-���b���E��+�����U�y{U�g����@휎��*-�d��Nn#��kna��f��s�����:!���v��|��K�+�]w�@�;Ҩ���z�u߀�ɴxM�U����#	��P=�Ox��{}��G���nG�G;��+��������T��;/�A�HM��+�Oe�� KƩ�����sZ��C��Ō�:T�[�Ƣݫ����p�<by���(=�����^7�0R��'����z�u�R�,=;���}<����;p���;2�t������I�}�m�/7!�ok'��h���e՞�'x��a����e�u¦�6� �;�����u��b�Fkų�|LK�������?U��#�n�M��P�=�	xk�Ba��5���u��r?���C���ؚr���S�;��|DDvր8���%�k)�8�xwVJ��V�8)� v��Ƭ�O��Xv�Tt�/71�=�-[{6G�A٘��KO7h^s{�����m�[��T@��+Y^��g��6�	�ͮ&�n�(\L�o{�oGgޟi����3��z
�����B�ʨ���Xf�ٷ����a�OD>��)H�����'�;�U��nD���������zt��0;r��7O5�似qǇt�P+:�����������<G���_�\��k0~�{^�����b�ql��=�1ޫD���WЖۣ��*��9ެ�^5�9=#
/j���#u�̟'[yժ�<���л����t����k�5�r�����X=F�;�~���5O��c�q��=�}Z��0�������)ig)��;�j_�O��b1:L�}S��ݯ8\���S���]�o��I�=SC��$�B���WU -���3�1y3��i����v*��Q��G���ɞ�s�Z<]��|������x�����ne0�߀����0�,Y/O=�ۜ�E(񬚥���]B��{m����nZ��*x�.��5n���́;/HGx����g^_7H���7{t:���Sai�j��y/u����9��~7<N��mT��"���	��}+�~����!�={����ww3����Z�j���2�}���L��[�t�R�GE�Į9��t��X�+տy�o�W�cT)u�K�)\�������x�C�ɽ o��f��q#��=�n�i<f�l�Ѳ:��b~�x&�x�zk��j=������<��+t�q=;�ӝ��dx(�__�t�wsA���=���>urӦ3�.x]�z惹����M��yP����w>�dq�;���e�w]<ǔ�z��ؗK�IG[F���#���:�w��;v�����V����o����}T����g������mJ���q��EF�4E9=Wk�ة�V�dи�=�p2�P�~�u������jsӎef{ս)Lt#�o�S�:�8�Q�+��j��$��y�^�����5s��'�gv
�^+t;α��8;�:���J�#�a�\	5�	��I���]Gxd�<�۷�3Bڍ��;��,i^��g��A�����U<1L�Ec�'���{�5n	����O�2yec�y=��`�k:���:;ǧ�����{���� L*��)��/�lW�I���X��7�m"G�����<�Ǉ򇼕m���4�A����g��eF�c\�"���<�ދ=�v�8G2��V�[�~4�+���o���#t��N,���:�3���7�G��#����,T�s{��Zo$aW��)�R!�!�$�K�q���@3�n��L:ݵd;}�ce^*ڏ�	��^�n*�|&���6�(�����g9�c}���`�0_xP�.�dwL�����gA����_SoN�͸D�<��(Ƿr��:�:vL�|X1$�a�#�~S�����ey~��=�����E����,���K�^�.�b�������Z�#k�^�	��NB�W��eY�L�K�e�G]����z#س�F@�p�lx�2}�-��޳��:l�l�sb�;i������}aw��T˒�~�^�W]���ُs�qD�F@�k��e��y2�G"�+��r��>u�w�뇅u_[��QG��J�u&�+[��\��7=��=FFz'_����Ɇ��nT5ґ^/O3�{�|:ch����U�o	UE{3�N;y����*��~23~��gs��z�]�fl�7�ܦ�v��mm�%;����BQW��;���[_��D�ߊ��]?���џ�'�ߦ%������V6�x��l{����D34+aZKR��'��;��ͮ���#;��Mu'��/q��p���d�`uw썓��lz뱙��A�nvϥ����V:d��(�힡=7O �u�P�ƠS�]���B~}�;ħ5녙W�U�m���i
�D���+�׊�U{LxWʄ�K�ѧ��*�ws�|�:�O���Gb��'>��W��_Z���2��b�v͛U�Ru��pt���� z.�ы�w��u8V�:��H��CH�/82�aܘoZH n��D�n� �;}�1�e��!c�#;A�y��r��t�����wRh���ٔ�.}��uH��2hB6z0
|�'��}V��d
�2�;��#kK1!JPtIZ{a\��j=+n��1���+��	�t�zf�a�g鑋����U���X#�aЈ�Вi�K:��M�K Qe��qV�/Ьh��̲�ĺug5)�6Kv�����j��RG�hR��I�k�CmAǝ�z\+Z�wK>ע�TѫCۙݲ�z-�E�JRW^���[����x��Oh��p��B�G.��)M��tt��[A�]�M�S���g,l�S�0�ÙmD�;�rI��<�"�T�q�����Ze�]H�C��c��oؖe��v�`�k�oWweMp��{nR�Z���xT
t>��oV�핹�fsf�����6�\FF�����cz�*Lx*�]���٫���Ρ�!5q�B[W�N34.�9H%Lݵ�1K;�2)V��Z���lr��YM��yJ�Њv�xT�k]�cyA\�7��j�;��w8���� K�W��b�q'��Á����;�Y(� R�fu�����[��4]�vӆmRC����ڱc(�۝xZ�|��v��.�	�]��g@{��o*����clB5�Mr�,#���t!E˗ty�9�wݱ�v�g���:
�8�9�7g%�A����pZ�q���&�C��)�F3;�m�k�j1��:���-��N�:��|�ī;Y����}��g݀2��YXq;0Vu�ʯ6��Yl>`N%�j���՗N���%�.�FH&�����5.���g�׼v�а��ݾn,��I5�r?��:�ZW��*rn�,F�Ͳ����ϴ���,��Ec�VU�[DJD&;���ۙDe�c�C�C.�,��\_U�6��A �۩W�Ȼj�^J�ŀ������
���x�(��i@c�r��
9x�p���Ԇ!��%Q|���fT��Tҏo���v�$q���n��:2Q�s2p�7�ҫ�,��ݢ�� �Ӱ�Q�C��ՇNZ�-ֽ<-�Դ�F��ps�����&��,�m�R��j�ɲ2]�ٮΚ,�r^(���x�#F��
�����n��
6�fr�'';.��ՙ��ܐ
a,p:VHt�o=�Dp���v��F�\y�FWin�;�8��&]�S����Y2��gx��^�j��d5{���a5m�ʒ	R����{��[)�˭���[�.�+��>�Q�f)��Y��ή��n�(�Q�[L���[i�,�(����q��(g+���:���jc���]0���2��SPp�ΎJ�I�)�:I[���\/#�&f�t�k��k;���f����h��[L��2u�`qt��OspNAQ�M	���Y�Y����m{nt�9rrt J,i�I��%|��U|�U
��*Aa�1�X����5
%I�!�H�b �X-���T�TU���2s�d*T�EZ��"��s���Dej���`T�U�0�XV���d� �B�P+3
�0YH�[Q�//���!D�V(���j���d3
��xэ�XV��X����%H,
�CZ&c�AH*�dր��0QAA�`�m���b�8°��b�kUD�rkE��H*��%a9�Ț�b�m]k"�dEH(��AE�� ��X��YEE�
�V���,��1J�d*q������E�XZU"���X��Lɐd� ��d����`�AIP�L��0��
$Y6-H����C�L̀�������u�7�������/��n�����e�vz�*x��4����WS�wL��� �r}������	ڜͷ�TO�;�|�cb��%u�f>E����������%U<o�ƻ��	zw���޼�[�kN�#<��?p�{!�W�NVy9[7�����u�Z3��ފ}9��=֞���g��������O~eY���Ɏ��jU~�[X���<w�~��������PL�2��n�Q�U��@�u����t��na���Nׂw��]�뵫��?["h{�-��rt���`K�U#޸�@	�;�']�����C�y��1*��6*�ƭZD����W>�9�y�読��;���Hc7��MS�Wx��|�bPW�bԫuy��Z�-V��|��~X�3�#J�Up���쉿��f�g��2��4<�S+}�Պ��8�>S��S!f��u��mN�`=�W8�ˁ�No��s�ۘn��k�x�+NV�կ ɏu��\n���n��.;ם���>� :5�e+9�3Ӯ�i�-�q6;�
�t�47�^��B�aEU�ͮ�1���N}�#ƣ���,��ǌ���]�����pa�HOlT��3��l=��hWV��s��淦,�T�{إmmY�O�殏D��|rd���z��ڳky�耭��2��Ӂ�����=��vѷ�k�=5sؗ(�[b�pM��7��ow^p<��Ӡr��l�"s�;���PtT ��s���Qe���y���mp��g��\t��@����D����=s�ს��]�њ�&cH�	.��UW��c83y�s�}�@��t�p�. ����w��U�f�_:�v1�3�U C3���K=�V��s�3���� s9�&�x,2��u��A� *��`q�{zm�8}��5n�f/u������	�ڐ3��6�_��*�z��t���+���E�朷��Y��9�*�)2�K(l$���~�4~��z��,��u�Tof}�US�����O�;��K5�v�E=�jY����*���r"}^��O��7�:â3hu�Qkv�8��E��h����S��UǦ�hz���_��m�zB>��ێ�A�{K������I��r��ߊѮcz��wN���@L)� Toepe�����-�������Y���<�±qf���;,��!��kɭ��X�_�\ �}���'Y�q�x�Sc(��O�l-ǧ��x3�Y����k���WHX�r&�g�7��&ofxz�7�	����;�e������
f���g�a/j�t�,�z\z�6r���PV�ƻ�,���X��+�F('��ݣ���}o!Zܞ4p�ۂRS�9/8��^;Ь��+ȳg�C��΃�k�\�gVic�[J�o����:BT��X�]���n3x��Ëx�v1Ǎ����\m���\�Nlf�7��=<n;ޢϋ����
�o����Y=�|I�{0u�|U�|�u�N������nU�r���*��޳��ݴ3p�)�9
��_K�=6�2���Λ�˕t����{�Y���-k������J��ʖcr#�+��9t�W~����pU�^�FE��&�4g$w�v鞇+�_��`�s�
��]�}�@z���áTu�h�=���:Q�	/����Thxw�����/��a��x��t�s��}�<*��ȷ��p���UuG>�`{ ��o(�����A�#�g>w4=q����M�>��T>5{��m���u�@p~���'׽��i=�9��=״E��G�A�:��]�����2 �>����G�j:�}T����y�q��}������6w��IS�w��dT<��"��TCF����_l`d�;E���P���,������y�����s��/�=BzP���9`[�� W��*t�A�A�>�������&b��MZ���M/��='�m)����b�H�}!t�*��Ϯ �xMH��H���5����~�<H'Ob%�;�$�7a�������C��YM����޶Y�"P��,5��A�� 3���ݼ6�<���\街;���C�k��2U�+�"e���n�#��Rw���gq�bp�My*u���"��t������ҧٙ*l��_kޝ/W��5�i�3������K"��w��wUI����r�MН���w���8L�%s�B��?Zx}�ƿ0��ٮT���ߎ��� LB���s�����r�Go{�=h�������#k��qY�_��n@׷E��lܴi~1W��k�LzǺo�.��2M�;���N�S7�T�o�,�
�[��\�ר��:|-�Ex{��x-���*U���O��g��?^�پ�XǇ�&�b�RL��N�NZY�;��̋����79z�6�>%�{']TE�t�ȿ�g��hE��J���ܽ�(���{{LX�\����uϧb���+�J.��8���@wS���|���f�� �>BE�h�������6�6u�ޗ���1�Yhp°������+�q���+��{ϱ���q�����q�Xh��烸�I�N�5ﶘ��]\'�ݗ0R����μ��o+��!)��S�2=Q:�@��}3y0ڜۘk�t��^�g�%jѶ�� qʯR۫���1��ڴ2��/"<d���L�G���~� �(N�+7j��LOp �ߐ0�_V~p!�\MKa�v��ݪ�T�\��;�vK�@Z�}6�1qwc�'�����g�W� �Z�~ܧ���������9�*��:x��@)�z�雨9�v������ϧj����W��~��Ǜ��:��Q�3t�{|V��H����{?���_���������T<�tPΘ�f�1(=Ͻv�"���|m����!��tg��筴w]x�5R�����������b��t����yz��l?���W5����`��G��7r���'��G�\*�\>�@�����)�	r���^3�����_Kӿ�s�^���)k��x�zX��P�).����
j�q�S�.)ߖ���	g�o��{:��:���� ��k)<�_���v��	N�׿mxq'��>�X<���yB�}>�MQgݣt\����P�/NUmpܜ�.gO�X�3_x�'}}�ō�>�
ꐞ�7r�v}��K�@��o�(z��x.#{�0F�������j���x�X/�o�u��#GFN,����V޽�u�]/��{]�<�c+}����·NuI��N���<7��wW����Hk�]�=�z@�\mH^���u�[���l{�ڬ�����%Gx�J,N����ZmFp,���3�n#����1�ޫ	�bo�u�=��l!��)�������Z\�Y��_^a�T���m�5޵۵K�3����q#�i���r6���36���O\C����mөhm궒R�v1Yv����[�,ͱ�j�{-�n��:]�˖�����곳{��u���]dQV�g=������b��za�a̫fX��Z�e�옮U��*#�D�L�L�\sfXw�w��eb�c�88�G�ag]"�9_�ּ�VѪ��ʵ� K�.���W����3a��NDm�7���[p�50�T�{��S鮟���Zo���aYR�� ��r򪑇ΰ6�	��[)���-����^��u�!��m��׷�}�a�����~.O˨�� =����v�� � 9f��o���/.�݂{eqw�Z����J�� u_[ȑq����O3	A��ֽAM�<���D�!��{޼����V��b����ޭg�� �T��9+t�[o���z�L�h^H�=�ک�>�1鋾ܬ9�{��[�xW��H�s��S�<�E9�ī���yv�*7�� �F��@�����~�s���۷�����y��/���y�ޣD+q���=���ϴ��O}���y�7@T=��4�.d�5)�g�{z;#�4�U��J.��~\a�[NK�F%8���*�V��G��K���D�5��v}�9@w�fG�������=��_�gޟ�}W�=2�k̿�:�s�1MCNh�!tTM�ven>����ވiظ�F���7v�V+%�����?
�_W?�>�2��\5�wKT�
�����1�#���A������j*��x��y��5�׉�k��#�Y���cW�!+U�w9 z��ɝ�9�s[�@�uh
�ዅ#�c�=7�4=W�?f��3J��:}Q�,��ި�?w����SZ/ڽ�.��A���X.c7�mp��z���i��ٱ�}��V���;�8�+��W����c8�W�u���e+7� {�6��r/:�3�{K�U���og^����z*=�紭mX�;�~��qS�\�(�ec�Ȝ'�;�x�	�ٞ���a9Lɟt���1�W���Gz0��h{�t�{�Ye�lu�Q��"o���ҙQ�Cb�Vn/w�׺�V���_��9��v�=qܬ�Y�3n��s�B�����4�rOo��I�r�J������E���bG��������WAIf=��]e� ?l+�k�zn���QJ;f�}���׺���3e���M�e5((�s��{�W���0�.���2�/>����������[�*r��3T�=ް2�Fw�\FV�b���H�C:9�gX֮G�{�;�*g�r�O��f��.fCsq�l�w��(&ڟV{k߆�6�~�{���?c�6��`�Z�Y���g/x��}DM����R�=��ԅYBaߪ�\L���F<��F`�q��k�j�U��<�0�@���2�k$I׳{[ǥ�NԍoR�6N�̰�㕬<�4�&���+�g���G��ve:�O�vwN�}L�vMĮew�=��(.��ȭʧD''�
��w=t����2�S���g��w%��2��;yc{�u��x�Lԛ� '�Dcʮ�-�ѿ�].;� f�;���9�:X�מ���k��W{��&7w��BaWJ�1��nT������x�=���fn��~&A�={��:��J`�(�n/���ݳ���p�|���P���ΐ�K2:}�ۀQ3"�I�:s�z�}n���59������г��{�7>����:�z��J�\)�Ȩ�\O\wUq�j����埳-�7Y0����q�
b'����clד{��=�L3}w|������*5m�<|�Tj��7uV�r��h���{���%�>ϡ��\�ȿ}�{�޹�>��`{�����	ɹ���Op^[d,���F��/npWG��:M~��r���U_����0aY��Q��G��1����ٱ�޷��cr����[���]22�c�]۹�YEޞ'��6���!W��ᑇV(�Y�_��{�aw��)�G�6d=��CК�%���Q�\ovQF7�(��8ˑ���ۙ?��3�f_�k��p�Y���Ófe>W��0�r�'w�Ec�{���ϻج�՜�c�����}{Y���b�/��}��[s�%�[��&�S�T�C�q��ʷ)>љs�B��b����{��{����ᦕ�V.m��N��[�>�=`s��J�2��ڰٽsc��--t�\�C�����<�?<�0_�a�71�|���NW
��j�@���d	�)�2�gc&Xh���w��:�����ѽ{���`ey�������]��2�5=�(���hz�u� \e��70ڛ�ܨk�#�^�:��ˑ��g��>)��j�1�g�����8`�v㮨+�u߆dl�7=�v3��e��#�t	7b��s_���];M��J7�qw��ECʧE���o�����`z�����uF����֤t���{�e�Av�h��gԦ.�;7���^tѢ����Q�9{Qdz���TT^_jR@����������;�Jx��4����o�S�+}�*gM��W�[3D�q���Y�=��3U��k	��2�&����^��K�M����� �^�y����|��k���uȻ�Ȍj���Śٯ*o`w�:{^�7�wL\)����ù%�m��z7z��>=���r�\k��O�EV�����2r�|'cŁ�=���3���Ք';��ݣ��:�	6)�����*�.)w��0Wm������u��k��+c�z��T�j���הj	nӝ�"����Bo���sW^B�C����Y�vK
����.W1܌V;�F��5o95�a��]���ke�*��D��M�gjî]�(����=��'�%��:=��p1~�W<r#�|&�+�{ޣ'|r'�P�N����Gg�¼z��ۊ�=>�c+��5�hn�?u+�[/:`Z�{���2��w�p��?
�9�'�E;{���+ϼ��-�;���;�U��HwR;�L0��	N{ũ�x=����b����1}��������w�ͨ��������3�o:@N��1��w�E��w\�.�cF����^����꽥���!}�WM�ONVDu\`��"p=�㤰ֺ�K�2�5P��k��=R��;�U�U�s���<9V+����<Vv��`=��s�U��@�ɴ������T6�5�;��^���^=�z�V�Un�aܩGs�u ��t��B��㮰FM��]�{�0��[�][�:����6���H�ƽ�ӟ{�x����XUt�.=1-��N�z�Fu�¼uU�4�[;�Ѿ��Xbn2y��:�j�2J.n2g[�q"��q�y�þ�^GC+���Z���j.����v՚�s*�9�w���珻������?}��םtW�$�$��@���@���HBIHBO��$!$��	!	'�$�$��HBI��	!	'�$�$��@��b��������$�$������$�$��HBI�HBO�@��	!	'� II; II?��d�Mer�\y~�Ad����v@�������}\ �"J(%)�%%(!B(�&m{*$T����!J�P	"PE%)kU�d�"��u��PJ"U(R�@�QT���)\��e�Zd���fU�Q�f�2Z�$�Jp:�X�mmp �  g` ʝXճP�KVd�5�!@(�nV��YP
 �� T1�t
6 2	)U�0 :h��[`���m�vV� 	 
��"� 
�� �@�4B�hS�Vl���h�H�
8 a�2�"�MI@ʹjM��f��3Ua`��PH�rv�*��ca�l�m�P��dm��hH�� �:�Z1(���m�m�*��(m�	i�B� ۔��CKY��ě�Eb��0�!BD� �9l��ձ**4ʕ��(���Lސ  ( M�C*TU4`с&�4�0B)����40L�2bhsLL�4a0LM0	�C`F�~%*���L� �10	�(�@#!��4�#S'��h�ɩ�i"4*�J0#d� �� #����t��j�OF��`R�c�K𝊨��-�(�sET�~�2PQ@�UT�5��(��P��3��X�O�Oڡ��`4B��AU �~R +$>I2�!�*B�I	$�Huv�t�kz���S�PUL%m�Q�Z�
|���S�����~��R�^�3����������!&ML�h3�I�׎�
E���na�]��ZqPt4���.�&7,<��]�nCo��8Kͻ��5�Nb�h��±T[݈,fF�/ �n�����B�l�b�p�h"��n2\�%��*e4&hX�T+��Pm��k@�T�R�`Y�K�W�We�)��j[�T�\m�IӘ��.��ql���+<�-�-���p᛫��2��=�^S���a�8M��*z�cEZu�v�Ť#�%sd˄<�GdvN��hI� �3�6K�Xޝ��M�F4�v�擡_�nSD 7Q�)��+R�n��Жp�A���kN��FR�EZ)c��IJC*:��c�^��]�6c8��A��	�V���`ufHs$6D/�f�%�4�7nv�	��u�RE�?'jGj.�f])Ղ#E�jh)��)RU �7�L�r�$��/*"�mBkrP�S,��c�Vn�_Z̭4M��el�|�Y��C��|��5���M�hzS�L,�y�����Aqhw7�F$�c8~��S�������N�;Tw��%�h���0�WV]�U�Űl�n��n��zmPtʪ�0���j�e`�A<2�JHI��VӨ�H�ܶ����mC����m�CU��]On���{Aط"�E,p��S33:���Uܖ���F�҈R�a�cb�:��u��j����E��1��Eh�F7ou�v+!����:5�T4a&�Z�2�v[��x!��Dؼ������YH��H���J�Cɪ��|�b�0�����o�����XP%	�좎���.2�Q�N�Lƅ��E�Z��5-^�m��ϓi�	0XwP�[�[�5Xt�K������SS��r�RI�zHg{���l�"�a���p�]�v�ލ�5���z��-�=' :n�ƞ���1�a"�T�5Z��r�9pG�Y�"���.��9��2��2�m6n6b�V�Z�YFW��V&<�5�*�r���N�&���8�xnͼ36��$��W7l��ieť����� Rܑ�H����$|O�PMO����8U��n+�r�6�e�ŤU�;��zu�ՓN�;M�ق)�{\��ea�8K��/.�=,'r�.²�:uq�M�6c(*�!ͧ,�Y�/�Q�k9srr����6D��:�N�8�4+M�r�9�rEm�*�ƥ��1�V��ѣE�%9���4 '�Ei�f�Ģ�w��2��N�8��NH�5�X�E�!��S�{`�Fe���=ׂ�w�ZU��e�Z�V��r�d���4D��f�9j�F2.�m�m2*S��d5�-�ˍ�ݜ��,�X��r�����"v.E�؀��w5���K�v4�"���C[���l%�$�>ە�	�\xp����Ԛġn�j�"ٖ�&�#ݢ�v��l�X�m0T�`�B�~�a��Oe,�ɉcw�@�1�T��j�����Ucq
���e�@KX�[V��Қl"3��^��l8��d{��a�L����h;9`	s/e�BM��.�pP��!d,طJ�)��r��lB㸆js.Y��=b�t�h:�&�D�V�@� L��K$�4aˡ6+zeilB*�Q�����yY�ue�x�^G��E[��ڡL���<���s2脉!�˓UirH�TF1s*�5�ӹ��oqX�K5��֥���������(��F3{�r�Ym�^3�Y�#wK`�u�	��1U�*�ŝ,x�5���x�4�w�r�P��ݥ�PlCu]������I!Wu���
Ń��ŝ�P��sTm�Զ@�m�`N��a���d;�!��K1�G2�ŧ/�%ճw���je�3"�y2�� %�!�0՗�
�4�wj���˫y{���R�D��r�7Q%S�i��ss@���0��S��Vb
�Ln鬯�Lq��oT#B,����f¼�y�F��,P��"��Th%M��aa�8�.�nnZ��Ħk�.�R�Z����mehr]�FڳW�D	3Je�We�&TZ�ˤ��w	y��5�4�kDK1F3�bF�Xl�'��T���&c֭-�[�ե�t��^b8H�y���%N�}U�ua!�P¦�C$��uN�f��&�
�Q�b)�g�CY���^`�Nn��2���!R�k"1������][N
k�*�ǩћ�TC��6s"N��p��Nh�5�o0�b�T� q���-!�7PB7�෻����۸�"W�bB]���NQu�[tZ@�P/,�eSyY���:�I���ư������7r� �gm;��TE�3^���a# �n��ʦ������Yu���r�tf@�g�d���iF�D��u��ĤՇqָ`�\���E�����F��Ff�3In[r%X��f6��)N��SB���;7G1�L8�nɹPdi�I�7�v������G{���ț�p�-n\l��.�Pt��z�\{���7�Jucյ�U;8�XFGq���MY�"nd�ق�*("��c�Ũ�ʹ#��Q�W���g!�t�`���c�M�x��4MH���f�	&Qq �;3Um$L��p͒��&Q�V%^F[�n�Hne�xK�D;w#(�ׇ!����Q�&i�4�ԗ[��\���\������?[�?��蜧BFS��$MZ{�L��X�Ǉ������o<��6d]�t���cW_e+�c����$g�FҪŝ[���e�ů�jK;pd�6�25k��ʻ�k����X���Cwn��Y����B�3��H��-o/���۶G5�m=��PR{�^��<�v)�l�\�������Un(���h�P������$k˟6���W!vV��J2��RyS�5o������	�ùEUsN<��7v_@���V+��J�F�`F�y�q[��6ˑ\�s�5�t��N��Z�UԪ1��Ƚ��<g�|���C6�S7�E֬�R�4Vbԧp��n��ӪY�(_g4;6Z{B�ӷd>�-�̊��L��_�Nt��\4�������7p)�>A�;�2�>z��|��M�Q8�V[�L]��׸x�PX����LPu�JQ�}P>�q��kz��(�KA��4w4�up��f_

6q�e�흛{K�ܜ�gĚ��$���w�#�8�EЬ���+%�9�i�����7���P�֪��2��z�U�Wk��[/6(ݳ@�3�UukpU���J�9;�'$��1Jõk�����6�K�oZX`��N��+��G.h��+�͛|��\�K��wu�`��5f�0�!w]�8�I��gjA��tks�{��Ҿ�Ъ֮ch(Ž��;8��Ʒ0�vj���/YXK�Řa���pZxD�'v�J��w-{.�]W�I���Ho ���x��at@:�N�d�}i���"p�,�h�\U&�U�DK�
�*Z�wCcy��dջw7!νq����of�pZogSPa��U��V�����v�d�"�一R���D�bn CڰN�cl�6a�����Y�e�vy���;dYl[g��E�c����qF�	��y��U0����/.fv,giɪ�2�UY��.��j����i��5#��z��d�e�D��Cmmg���#>3d� 7���-C&���w���m	�:l#1B7z� ������=�y}b��%�en+�7�"�,qߟn��y�{�c�D��;8��yלq �ͻ�e�ͣ.�DJ
Lȴ˫��ڼF�>BQp����W��+���X8]�8m��ʸh�BP����PL�#�baC+��bޜ>-Jm��� 7a]ـ�����5�U#'L���i�/��
���!�z�*�1�����a�+�����	^ރ�iQ�+b7\�wC�˕k�%*�$��O���Jg�P]�Hm�Euf�Х�۪͗)\�3H9�VCOe��1$��L������t�U�KFN�ƒ����Ҳ�T�u���)g$,Vs�9i�-X#2��,u�;s@�%=�;,3�B�)�i�÷w.�BN�[�2X9a�]-	��J9�oyXi,Z�ޏkVW07�y�fW�f�,��R�&�u��L&��IݫH�K���̔8�<ؗ� �K�m��n:���Z�S�Dqڅ��V-9fI�ҕ[O&���㯘x֢��A�v�5��苼�0�}}F��b!:� �4�P͈���:M��7�
���7x��i,}�2Z2�F��bC����F.�\�Śk�<�YxF
�4�����,ծv�V+xk�jӬ�d�i+��&�8��JƓyK�ɩ�9\H��� Q-H'D�Ìr6�1g�.v�p|6�0d�O��ֻ9�V!�b�[x�l�sI	���.?2)��iy���:�(_^�]�$�&��lEY��¸B�n>�x�w3®��ff�0'��cV`���vO,�Y8=#�.��z��6Џt�2��Z�+�!%<p������ʴ�� ���;th���*Xv:,��j[�|�y}4�ٔ ���{ l��o�f
�ɽ�UiT�;����j�ݎ�����N�pY��ζ8,�-�:AX��8�#�ff�CW ��K��T)n�F̼amM��{`Ϋ|͘�yz���_P��w^E�Fb�Z��"��o�����z*�V����1M`VԤ���2
޽-��hX�������2!zR2��gz��o�NE�"[�iB�t���qJ=�y�{[��&��S
h�Z��n�B�ve�g+k��/J'u�Ǖ3wt����G����s˧I�R���Iۙvn���FtRC���V3����`j�����R���;�к�ju����g*��fsonT�]���`��b��:e�n��F󍥼A2��j�WV���]��sGq�;RcY��d�ѼN�q�3�!�s)�)s�;��֮;�m�YQ*�Qخ���q4��	R�553�}�E�V�ɂm�h8NẾ��O?�{���9;�g����D>�1N����O�j16W
R{u��,�W/u�f���c��}�\�խ�e,�uq�+fӿ�9n]�H���F�oF\\\1���1՝q��]C������Ig^��H�	�=Y7�[�b�)�TN��Unxtz�1ٔ�[O JX�l�Z���/d�`����s�wZ���<Q0�훶�`
�7��� �X)�
�l��N�^��ŅK�/4����!��f��C��8�'�C	���q��7
�ЮR@Ƚ4[f��C��z�@���KJE
�T�o+��)���m䚥+����b��VuL�9�w��8��i=��Y���f��;j6Y8��ܣ�+q���kbWVWvm�oV��YK���zCt�����1\mJ�0e��Y��wfÞ�F��H�&�b����V�+d � �H����S��!��4�}7�f�֯DI����pTY�Z(���s6�6xP���j��. ��n�U"r�t�Y��$ؓ��Z����Í��a}�Xz�;Gz���n�g3@s*W
�J�	��mپ'�M(��eYUK�e���i�]���Q�E�SvW\09o�0D�ضl2�6+r�eZ��y��j-!VfWe��_��gT�P1|��h�M:�����VX�<�t*bZ��vSy��ٚ�6lP��5�����%�����C�;�s���L��e��;�VWD�`����a׷���ծ�z.�vѮ^.am.����E�u�Va�K�,S��iGvi8�͝E��`�	�Q�f��Gi'w�8'�Ү���֥.Ag\�@����j4�8���n��'�n�޹X�흛BmZ ���3�`v��8��ȳ>��oqOh��/3*cr�2ڐ�_n�"caLu[��Dh��;��U�X!���������-��C�gh�$���63�Xm*'y�s��ή�L0�*�JR�@�̡;�j<�A��\�+γ���w�+C�t��l�9Զ3�d®�u`�r�۶��g��'8=��p�o�u2����'Q�B���9�S*��ٔ�)J���G���D3.���+/��Pia��G*jݮճ֞b�b���f��tY�(s|.�}ҷQ@q}K�_q��,��H���GaV���q�J4���k�q�Z�]6�V�qo.��@��ӢiT�u;�aA#C����7y��34�x�M;�B�����gU*�ʘ����-���	'59���/�*;�Y�"�3��N��ġ��cz��uҺ-u���E���U�p�٦	+$۸���{t�}���Zv�&��7^�����3�_U�!�v�iK��h��ONy�]w&ݗSdW/�	v�[B��c�a�;��t��Z:�\n�.rw�fn���B���S4�9s!ݸ��z���$H7�#튲�x1�wֻ�8Xkf�ѝ4�jʵ����J�M�f�v�d�%k��~!Uf�0�C�+i�wM��ۢ�m��f�;� �6��NS�F�?5�U'��ٕ"���	W��Yʤy:��u��+-˶��+WqJ�1Z��� ���Ѹ�Βv��cB)�~���*t6��%+��[�^gaͪ��,E&Bwǂ�+BO:�Ӓ�=Ʃ��`z�ؖf���6Fv���|H��7�A����B7n�_t��9ۋWJ���ZѷmT�u��@�VK���2����aQ���5�ٹ0=�w�q����CFfR�u�QX�2([������r0;���;uX���':�Y�V-o�q��co��hv�o�c#n�����If�X8�=���1�a��p��Z q��&m��K]�6�h�ܪ��g__S��mp��ϰR�t��������>l���T�ɰK3��Bᬬ6�>��\5��F���9�\
qj�|p'A�ͽ���n�
�b���pm��y+(Dzhr-�]������*PD�i1w
�m�woI*5��d�+}�d�������Z�K�B{�q�-���	���Ne;��$�qV��f q��'#W��M!���y0Hc�ucT�δ1l���*��9�5�Q7��ck�uۭ�i3x"�m��dˊ���@OU-���K>D�����a��G�����Q&6�"1
�;�%#19|	�q[����q���v_ӥ��z���(����A|��xv镝ئ�8>ӆ�ŏ_u�o��k����t�� ���)��s*�>:��
$NʾD����t�(�nB�V����ۏ�Cf�4���L8}yA��c3��������֜/�vb�-;�x�d��v�|��2�ak#�%�:��*�)u�L�M���r���΅ӠY�%(e�83G��t�u�諘k(��[��L}\#��Ƌ�C�6�ܭ9D���d۲��v�x� X���w�,��ҫ���5�	�����-�㓰qְ	���qw
x��ռY��Q{:���=�Wt:{�u�P2������<X�3�C�R'ւ���k�����pd�kh�ȸ7-�2*adyyYp��IÝ��h\���鐳7�J�-,J�6�7�.�{7rgwƁ�y�6��%�2��s�������Һ�ǤV�NF밧��� 3V񦻞H���i�\�Kr�Z��̼�KL���H�;aI��u*�i��*j7Q^���xU����g�Hn�;o��,�s���<�ۗGp\�5�5�%��6�ooVu�L��|�^��W[;<�c��Fp��c��²Q��V�]����ɥ��A6sx�wK��A�c��v�����,-[�Z��"��]�5}v%@����.����։\,�uY�V�$�|f|��n��&P�|��`�O�9�/1�ZgWe-������O+��.��*�D�4�ݲb�G��Eu.Α�����e[�M�q��Qڙb�S�S��o��#{��xd� ���i<�����[u���3ī��f�?U��q��>�Ks��!.�*n��"�X=�����$�+6Q�D���YC��}֎���i1�ig����.#�xl݉�&$0��yji�ٝw8�Z�M�Ud�X�|�� �x�ڦMF8˙[��2VS�F���30�RT��qlsHYD�F�Ls�~�\�_��S5E��T� �[�o�ιNL��`�dۼ��:�i{y�o��?HIH����K���G����D�/?���6Lwe�9V���d ��0��\���Ӷ%Ed\��dՕ��>�=�X��=ڥ��Vh���b�{�\�⒛i�w�[y���x�����;�*����#�7O�2:�ֶ�CH`�̱��2+ͣ;�>'�!�2��q��v6���%$!�M���O�X˅�xNqjͻ��w�'YJ���aT/h�!i�9�c�v��� �R�"{�����r�˝R��.�=�F����ۢ�!(�gt�Z����@�zq���sI�A���V������vt��՜h,!S\�/&u�u�B���C�Cqb�v�Y�+J3�Ng���/.��L�u�-<��Y4����ڋƵ��m�|�r�ُc�R�mGU�Lq.̘.�,cuF�,х�
�3�E*6�!�V
е���d��Qvʐ�T���4Eĩl����m⫕j,X�����2ɂR�Դ�����Z*�K�J�̶���nYLi�U��t��_�y�ؓ��N�dέ▻��3���rՙ��Yj ��ި�x�M9?����=��u��wI�t�4��B�n�W�^�������G��	:�ɵ�`�y�3ޙ��G;�[}U����n�(㈀�X��ET�v�Pʀ����>Y�R���h�\K���u�We��#gu�(-�}�x�̊�:q�Ӭ˚���t~�_�}S�B��s�!�8DҪ�~�L�[��S����'X�Ti��vWvu30.2"�r�G�erCXu�&v�W�틗o(X�F���Q��<�3���HX�j�N$Z�H�k��t�SY��az���u9�"��۵S��������K�Ԑ�P���.C�B�Y��N�Wwz�5�hy��/@�4E Vwmd�s��b�^C�%���Z����j�|oSس�u��IV��J�"NmY�J�����D��v����!}εm�ԫ#�<����퓳��M�ˬf�Q��q�C�]��9�WtQν���vkWN1sX��,�-��'dK�9���$	��^A����5n@\½=���(�k��l�46�.�����+��g��=K�����,�b4��;����j�N�;]ǥ���R� P��Cw+����~ȍK~�Y������FP�U{6X����Y�K6����Q���~����%t�ٽ�),�]Zjm��7K�Z.q�MP�x��V�_n8����aX�%�"�1}C���zJ�'��	1�����!2�2u����iG����]�/m��]Yjk��
�ï���m�!}��!G�4]�w�7A�g�~��s�;<"���{��c��6��mT�kޙ�����!�M"q��K�Wu���8d���oW����/dpo��~���u{�VYx��m��ce ���7�0z�q3�]u_d��NaA!�9���Si
,�ؑo���˰.\�ؑ/k�^��l���ʴi1^�گ ��c����Sć�� 9����-.�Q�<J�B��<+J�U�g�$�����"0E=�H�ٔ�{Z��f�-q�W� �������>��ձ����B�N�oUCu�A�+��(���F�B$>�J�}�u8����N=�|#���z\��hp�����b:�~�LR]c�x���@��7�.�f��z�#!�_J�:��x��{��p����{ �|�<�x��8�/�$z�����	�5���Άy�m���|*x�p�*����3ֺ�:��R�eN-�-]-�;KK�)�8��^���>�y�י�m�q}I���{�ϵ9X<�7.�Eߝ��^V�CQ�\�yP�1�j��U�����pq���b���O�C�l�]���q��M�#�m�3{5�	�������v�:1F�� dK��;^�����ɱ��VΡA��<�:�3	Z����;�Ϳ}���2/��#��y�=�1K�+$���3�k,FUS"�\k�%�1V�]F�H��UmGv�spdsY�lm����
��[��R�GS�D���q"���c&���j�u�{εixZ���wMJ,fj�Ί4.]���NC���%�A��#�f
&EC�3A�:ce
qI�n�F������&� g��ִ�Tڎ�y^1<h�Sg���[έD��ڇ�^��X��N�Fd�u���-e�1Qw�(IT���o�qˇ������ X���3]x�j���״%�j��}�]R�>���*���]=�ޙ�&F�í����/E�yR�7^x�kgP������'/x��!�4��Uo_�(�F��X�B�x�q��Q��޸{�%��t~4O6��羖�')�+�eV��-��sc��l^*a����U��)����7S�ѼQY۝f�+�!A�s����R6���=�;
��׹
	����ܸ$~dW����g�y���ݦ=�����0Ђڋ� h��ǖ������KG~�ًl\�:A�K�N��ҏR9�}]��Nr��hv)��q����lZٞ۴7}�����g��e�������}�2��^�ϸ���3��h[�Ή��7��gq�#?A��N8
���֨\���vvaCݓ�]�����Of��2��*5�=�mMeP�s=�ל�,�ok} ��.����G�@ꨏ�u����n~��V[�v�O�b���wH6�2��H���
���e��u���|����Ǉ0�O"���p�,%,hwG�6�I����e���&<SQ�0d���n�gV�J��m 9Y�A]L��Q `TQֱ^u����2`V�F��7E�&B��Q	L��{%ĚD��jӴ�߱}�OmNư2�vLT+a6z��h�#�uE���i^c˦��v��*�Xo��n��&�tp-��&�bLÃ�mТ�n�/�t�N�	oS�Se��QO#s�a�ee���*Ӳ���y�P.'�ٸ3��;)wqX�u`������#����T#�?b93.��K5MH�K��NT����b*6����!�)Ve���Co
c+�����2�4� i&�V���,�F�T��uʺAX�+�D�M9J��[8h�I'r�າj�d�J��N�?U�a���r�Tt�ƙ��<�j�/�K#Vh�M�i�Hw,1j�8���cx�7Qҙ��hEt͚PY���M*�Wb��lc,��Z7i����ۺV=6���eݠʶFTR��t�vPvIs��)`y1��U���E�Zd�SI�)T���eml�[s�Q���*�B���2�D�(UJ�Q+Z%m+G�Z#����T�Z"��i��5q��iR�̙PI\�]fZ�չpPf%e(�،c�T���ۘ �V�m
�4�k,TAW.c�E�V�Q��`���UDZ��L1��*����
�[iR�Tk)+X�kU*]�e������Iw�����'r���}�YC�jt�h�o)�ڛH�(~b�bJ�́r�N�lX��]r�W����۴��룮o��g�\ɂ��O��g��9�]���VAE�W�#���L��<yw$n3��h�j��Q�n�GP�/<�s�1)C*H�׹&кz���p�d���8�:v����,��	~U��F,���A!���}�nh�y %ڣp�,&*at��Ɍ�^�8�>��2h��|\��NШ��S����.�}{�|\������D/��|ਆw���`���*�n����^��-��O����x����Zy
NfԳ.5��<c�<cTa/=m�דž�c/PE�<���L��WY0��aZvլ'pb�w�%�n��/��y��y�5-�_�zd.rp�"�w^e\������k����1�\�o!��xl��l��ż��YI."���\��,Y��p�g�Ga\�jU{�(��~����mJ��ZQ�u�=y|��~�OP�ڰ6��{@6ɉ �C��m�{��z����	�C�y�$��>d����t�8��2L$�+42C�!F�Mw{>�[׽�N�
ä���C�E���=@<dz�C�Xa3����u�:�=���g��	*M��ya�E���	״��C�� x�-��~�}�y�:쒲2�@�=d3��Y$�N��0�$s��3�z�k;��v�LÖi'lXm�>I@�4��!�$6�y��o�v@��z�@�B��P��N0��$�"�a�����{ߞ��hN�;�i��'�!�4��!���$�dRC�CZ��wN�{����V�R]�xlq�4Z�<�X ؛L��O�З�z�����w-uN�jb�3{K�(볡]Rd�)̾���� |6 ,��������L3�&�>�	Ht�z����9�y�߻~>�2I��@�0'�P�2Mn�x�g���:�B�`�P2kT����!�M�4�8�t�|Éo!8�d1	���ף>׾w� v�kTL��Hb��bI�@��m��a���!����=ߞH���2Hv��d�c'��Xb��6�t�J�j�m�����o�o���!��A݁4�<}@�I�	���Aa'�T�큽}ׇ^���x�@���$o� �{g�j��I��x��M2C�1�;���o�ô���$�a<`gT'��i�%By�N!��L�dk�מo�
�v{d�d��1�1/ف�I6ȡ�PY<d���&��a��ν�� v�|ræCl�I,Ę�I1��NXq m�l�����ƚ������_�x?t~𾓵alh��/ї�N�Ӣ�d���*��Թ5#��|�v�$M�������6+�X�ߝ� s7����}RC��܁�Hm �%�(�CL!�&!2�$�����������$4�l��:CH����Ha� t�2I�w|�:���o|��<H�i��ā�I��x��q���$+$T� �W��ߞs�M2)!�=� �gl�a:d>Buߙ&�	��P�RC�����t}{�I2t� |���+8��I�C�b��I���z�{�ۭ��~xHm+y2� |�OP�I'���!���'���/W���>�~�Hx�+ d�$Et��8�OSH�>C���w���'�!���i&�O2|y�HfRI��C�Ci�&�������{$/t>` O����$>�CL&��6ɟRAI���=����p�/Ͼ�0f4��*�����1uK�-<���NjE����XW����K=Xw�*1s��j.S����u��Zw*���E�+�7��ψB�n�܏��=*�7�,ro��듗5ug�Ҵw���^.c�Y��AX�Dz�fҸ$����k'�:4�<u{��@�{����r�g�7s�Y���@��2�գ���{;�R��I�+c���c\�
��r��,"!X����s<o���X<f�/��;4� rz��]�]IL��W1��v��^���n�Nc�y�b�-�=]n�r�F!�������'_���z����%���W�:1����T�GE]�Y�SeH��5~�g�r�9��h��)�K��f(U�;8��S7i�v�+���'�/�Z���zyWTp7��\v��_�k�����]
�F���{�;��l	���[L�I(�k�a���'���V�C�ށP�:!2G�<7t�M�!��4>4X�ή[;����5F�*.��Ċ���ǽ��Ƴ�A�z�~*�юR�E'�N�C��L_V%��>}c-k]ŷ�E6�j��}��#0���-���:^�;���F�Ch���̘���gS�oWB��}��a���Dwb���E������[�޾u0\����.����?{%���E��Yc8oQ+���nθ�ub�Ӑ���r���Y�h�Saի�V���}�QƔ�Ǉyk�v�����I�w3㹼������<h�P#u-�}3�8M�E�
{�]���{;�M�[�K�e���*,�	�tj����V�c=lpN�0=���ﶇ��FvHv��Cd�~����t^��՚�������E��`��N>�Ȳ3�x�H,�9��,�oF"��Y��ju�U��KJ�]�v�<�O-�=s�_W�3�i�Jf�~��ͷu.c,w��nj�әG�*�cMq����5c~�{y�+~k�#�Gn:y�8�mgL���[U�<c���݇6�{XU����@������ن�.��`�'��K-���D9@���\3�(��g6�7�\�K%^N���瑻�ٵ6o�G������N�p�Ij�o?N
���1(:�j+J5��HTJ@.��^Y}÷��Qr��KZ�����wHn��NF�$��N���iyϷ� ]�l�E�(1Z���1�TU�\{)-Ntq}ϲLllɜ
�F	V�����Xu�a��=vҺ��ر+	�����؝'n�vth���8��6�-�0m^�i�����R�F�Юf��d$nq�=ӓξ�Y��hD�P��]qJY�����Źs3�WAP�h$T<�:��9M������V�*.F<�{Wu�a$vk۷G^����6"����f&<ʪ��LD�Euc(ӫytn�˙�]�D@��5x�n���2�)w!7�ںU
�u���l*TLT�wNWbf�.\������*�6,�2S˷Ӓc�m��EBY-�t/��ӳR��Z�;�	KaŖ#�E]����K*�h�SF]�R�7��.K'2�UjbT�k��b���Ǖ��?��~I䥦�!Zk��/���(��J�]J�42����D�Yh;�ƕ�B�uM��'r\��l�E�.����Ř�=�O���Z�lKj(�m�y٣ tƅ��TLPE���Z��`�������UbT� �EDb-j�J(�-mp�9F�
�f�ĭ���l�ND\*�Q�F���n�1әlT�m��R�Y�9u�QZ�T����EE)��j)��m�lXb\��բۤӦ)���*�,EZ&%��T�*\Jj�]&ZejĬ�1s��,�Tֱ¥�]eS�SK@Q!�IA&{��������Ѯ�U�'t�1�r�v���j���=���L����ХD��dӪ�e�+~����Z#�3��QI���]�PD3}EB�v��w�{[�:g����+���C����5��/x�x�gB������F{�F���b}~w���:;!aQ&����Jr��	�
�(3s��W��?��Omb�ށmp%{��N�����#,e���_e��P*G�A�Ы)6���Z�%��+�ވ�Y�mJ��Z�i��#��ǒj�C�P��~�2�� �Ӿr��LI�r~wo�}4��G{i�}j��Y�Q>O�&K��{=��yHz�=���[cxSB�'���g���q&���nlq[��'�	a5ï���������5{K�ڮw3qu�����tq`�+J�]���N�vaj&�����I�>�����+�k�OT�^U�j�*�Ww7�>��`����fcަ%I��A��_W�U�g߻���.��[٧+�f�y���4;O`��y�o�<�9Z���
} EMq��`е�W� �4����o_��E҇&:r|fڌ��8	"c�`6n��[�����a�-�c����a���5����B����=\��0�6=�j�e�\y�\(��Q��=H����^-c�Ǹn*"�d7���Q�����U��>�!^�8�:��d`"�-��O�c�5�'��F49�4�~����;�M�x�7t�
�������%���^�"�ݽ_��0�+��u&��w�$-��m ���>�;�5��W���*�㚀����h#ƹ��
��jX~�`4u�H�VE����kh"egu�k����#m>6E�j�߽Y79�Ȩ���hY`R$if����=��]=^��~��_+5-�IC�����wÎ�m����U�����3�\(ab ��Qdm��3)�����0���H����X����}��/V?A� �+��&]߯~����O
XQ�A��D;B�l����_�(�����9_:8~o�E�*��zޛkP>�m�GV��o�}]=�d���j���>~�}����������8c�|�Sy����=��z�s�dC��+��h�b2�L8�"@3��;�G^�w�#O�x����f��XY����l�J����Ad!�q:���y�*<l�Len�����h��M��c^/��8��U������x�8Y�ύ����Q+�omܴ+�"G�4@Qm�qYʕ�&,�.��q}��9i� 8B�l��B�Γ�V����Y}~#91$(�(�_�i�ʐ���g�Ŧ�z��2��+���R����p����^+#؅��A�߫W�;M�)P}{Ŕ�렎[�BY��;��=$�5�[���p����Gq"�oa9�Q�ї�;U���G���t��L�8Ѣ?\b/��M|t��:n�}�0�0��CM�����X����L���Z;�{��1��C㦚�����(�>�?c�t���{V���k;0�{b���p��䇨sx���^Zl�<��	^���B~�X�~Æ�H,��va�!������i�܂. �4�`�$����V����Np�1��a��VGMr�<��ݽ�8�>5���#��<�DN̓�n�,$���m@(�0�FF�Z���;"yɻ�˧L��Y;"7ݻ���&'hg��7�]��!ڷ4�j�'���Ret�g�������V9�W��_!��X�=hiG�zy"�!�
�=0b��0r
�s_�6R/�:)r�}@�><F�U�x�ҭ�f���:ݲ����&1�B�&`��Z���o�Ŧ�=�xn��,��X;1�f�񻌘��w�׫a�1c�F���F:@�gh����V/��n z�.V�rbL����g�pr�e���ǹ-YdY����%�_�y�r]f�_D�㚂�b�Hx��,��#�e]g�3�$/���D4x��ma�B�zS�{�{.�N�C�`��2 �XK6bvk��9��5��g'��ާ�go1oU��ج���{��v F���\%!*]�����y�s~�������Y��6�[��ׯ�֍Ի��8��ȅ�e����M�0X?e����V��y
8D�֎�˗xB͒pyq�M���ƃg�=_Zt�VJ�{��0�$�.��ҝ.�	���/4@Sm��q�a'���#ؾ�Ԇ�ax�����nT���:A�<Q�,�:л�d25�����T��av�^/����f�#Ɓ�G���oY[�Nr��ڹ����wj�����^��[��G��;Ur����G�PÑ

���7�,��`��%�R�e_\J��:뭁L(l�|>������TC��?���ȣDB���»��T\�1��P*(m}�Y���퇖�ڽܽ���D**-��6�v�Y]��6x��b�~�鐑D{U�?aC��hQ����z�he�7�H�✨�t��F�����Ne�q��d��م0@�<�ߓ�����=yM4~���c�|��:qcUE�Əv����GjFD['�"�.:F�}�n+��m��Ehx���"��ƭ���;����qHw��E�Dv��*�I��ǌ�*�'D�Mx��fRn���5k#�4}���4$y49���RP�6�[���ߢ=�DC�OL}�'�4���!��#�r�����,��r�G��:� �+�״��x�'�_^/!���?YN��ə�~���A9Y�-}UN���!Df���A�c}_Ʒ G��?�ɟ,��ǎ�9KK��#W��ظ��K$��a�!慝�Ǎb�м����"�a��,������p�CW��WR��DC��O1� �v`��?��,�G*��>�׺�j�g�F����?"�NZl���·�/~���D4p�0�I��k�U�r��j�W����[�2�����^���A�k	e�C��r�'w<*���IXg����-k՞�լG��� DgOmf�R&��1���N���Y3�ϗu�{fW�x��v1$s<��K_m����;&���^cW����ms�"���6zܑQ���
��M Mbq�(};"�v� ޢl�X+�T��K{:^�R�k�F�R����]F�T:j��d�gN�fr�n�C�sv�ch;��XV��+ST�3�mڝ]h�¥\�꼋5@�F8������9a��t�6��f�7R���^��ĉ���&p	匣�;��(��U��ST@T�]��"&9��7�,��EGLÆ��I�lZb�[�1,�o^�)Ej�X��n�
fa�lr�Z�WD��c�2���-;�j݅�Z�[�6J��Q�����N��&�v�v���Ƽ�KT鐒����{�t$���b����^����X�zp���2��mKd�,�4L3"sٺ� �J��s�v_�͝QAUx�+���s-��m�t��V�j�8�㬮[t�0�*��2�e�Q�R��֦%Erю\2ԭʨ�-"ELj��(���8㎵3(�Y�lmm��ܰ��GB��L�ciEAr�5�""%jbam�0U���*9rk�u5�LәG�1h�uq�E����.Z6�U�c`�Z����B���r��ۉ����堖�bkV
w���G��- �E�rKU��R�쮋W����W��yS�k����Ղ.&ũ^"�6<�~Ӌ��u��=��~v`!���=h��-1��%`�Z=�t��}i�iT^0ѲhQ�(��fN '�B����(�C��_=�M��~�/BD)lkVp�z�=�w*��M�Tk%[���"ȳ3�N�<����a���C���#Ɓ@� =�q�w�m,0�e�;��6G�г���6j!>9��o���ۺЯ�!�`�eY�h�5T�ȧثg��F�Qh�J��{̈́F:~�^c�-^������Sb���9�K%�!<���I�{����/�8��я�����W"dj^���oW���;3^M.ةΎ;�����.���>،���)V��)�Z'�`�.��A[���qՃ�kA�t��,لY	����^� �k35ȟX2�ʉ��θDi���9�����O(x�m�E��>4t�XF��]��oo��=����ɡDQ",m��x�;��OI�yG^ ~�Q��I{z��#5
���4�X��/)a~Z����#ڄ;����I8kPY�t!�����nɺ�|Y|FET�$XsP��;��ӭ���3�@g��P"�7G����|��0w�1���1f�Q�3�k�G��{��|�����5�
4F��A����s�-T����v{.ՙ��a��f�0��f�Z�]������������fZ�#�<�{���.����j�b���"���FȜ�1��1�,y8aW��u��O�ʎ�?Bߞ������d�~ľ�}�ap������x��(��Q�RZ��`U��`��\wZ�<�R/��h���Q�
�.УO#�X�f>Ho��s�9Q���F�8[N�P�A(||k��z��xX�I��L9�;�$��g~�Ze��{RX����!�U�la��=�=[h�r��8��NWnu�.�N��W�}_D���l� ~����*'?1���q8��~��}˼L��nag�!�b�@��?i��Akxz}��Q~C��x�\�Z���)hjv|�E�: 8��#��-�7�Z��Y��#��x�6H�fv
̍{�D�C����KMo��V�����b��,�ԍ<Gx�?o׏���^�<@�����§W���CZ�<YJ��{�����>�i�1
ǮT��-���9���:q�����5��6.X&7A�0#'��mx�z���:fY=������ֲRt��vΚ8�o�n�T���h�燯p�ݓ��8�N�?z"#���Р?Z�b�,#�>����D@~��`��3�Sί�F!a��Q�_X"���6��ᕹ�5����!0�m�z���̵�̎I�ǭ4U���R�4�f�6��c'_m��J4ChQ��4�)������=�zyJ�M(f 7�P�C�,��� |��O�exv�"��Y�M59Q@DU:�[��3F�!�\I�_omA��!�
>�ݿw���Ӥ���a�vw؃9�������?*��8�O!�Y�-8~�L񃐺�~�T�f�H���ɠ��O>`�����S0>��Įm�S<���1F�'U.��ؔ����l�D��N�U᜸́�!��G����_}�&�����Y���g�t����hzo]��ڵE���h��o�G�~�0Ц�hY�Ƈ�z��x3/k�í��<B>����U=L�ݸ'px<�Mv���l��vx¹��X�í��2���!�_d�3�̈rС����W?���x���Li���2�"��(��_b�f�*h�Pv��~��DJC�B�>:[�y�NGR��#͌���j���YҞy�zv�z��yhQ�����:A%m��]}�����=��C��7����i;��t�����Ť)=����7���e��_BIv�[;�����\��Vx�����}ix�8G�珍��(�7h�<p�gu�Pme�S���Ay}��ύ�̣�B"%�YU.����r��N�>��?@l����W):j�뽡&�h#�W*#>!_;b�itu^�@����\C���4I���v����?8�������GM��$����W��J�D��jf,X~�Q��!\�&��E��#z�dz��BC"�yQz���6���l�-0��ϖa�Lv��B��y�{�dxf��RԹ����=��&�l�k� *��W����1+{)"�_G�=᫮��FZp�$3�,-��$,�[�;���G���B}-�:��P��dp�5����(�i�Ϗ"a��ʴ�o��Hތojn�{�|Fj�I����]ӿ��S��@
*z��D�jW�!�?q�D�c���q�ު�����V0��qu�
�?i�z,�~���A��EB8�*6~F,�
ksy�6v��-�C��8L�D;CA
#�4G�κ���A�7�l����t�_a�a�n��T��dY�[Z����	�aHC<�B�C��Q2Ε.�b�I��YW�s�:���kSX����)̣K���;����v�p���D�#N�#O�s&�!�z��#��F,:��x2�~`���T���Xh��VG��C� {�F�_yiӾ���O=���}R�>�GR�C�f��K�����a�!D*Bj�=�d�g�M�D|�,���P����Ԩ��;Q"T_!{o��ޑ�w�Q�I�|~E҇�Ӫ����?R_x��>",��0�I�K�+E��m0t�Ah0E���O��Uz����еٜ��L�1p/���8;�8_����7�[ԝ�ui��yK�ę���Ki�3s�{P�1_b���.M�����E=߾�ꯣ}��������F,%�A�Q@�
�<��dV�X��rƿ�i�0��㕘��mF$��.�<���PE�C��3j�]?V��y>:o�(��5���r�[�Z���"Ϗ�C]l^!�.o��=��#�P�/��hcB���f��s�_d�u]���7Hw�����(�<E�I�c�=��c�|�jU��ݘ3���3ٛ��M�<j��k�e7��屦��k-���=[s�M�>6Yƨ��6l�!:a}����]������%�_(�KDM툅��`{��\��n��<���Kޘ�֗}�^���f�q���r,��~�(1��k��z�)j����*�_7��u�k"Ѱ�n��SԷ%�-鼮4�V!4G�q4˗+���
��'�H�g�P�"�z��/����<��7gBd��p�VfM���ͮ��uz�|�	��U��l�
w:�\�9c�Y%�&^�d�.ND��Ü�Xp5�]��.�*L��jՓ]#�2$�j�Ö
O-�r��wC:��bƙ�ȅ��w�u�xp>A��� �}g}�H��$Oq�6�M��@�=��슬Ҽ�2%���<[�����*8�������eI�>���Wm�n���l�÷Ի�����+�Y�e1ec6,^&�/�0�elZxX�uk9�w)<z�Uk�Ò��g�sC:9�|�9�g�דp�~��<+1�<FW,�gv���;������=�KnC��^���&�`���Y���`6!�j�%�e^k��Xu}ݚ�5����Vc�٭+;y�J�;�)VL|.bt[:�6��Ҧ��O�;e"�����˷]�h�Z�IZ�Z�VT\r�eE
��UV
)E�b ����,X�et��ʠ��m����-Dkm1ȍT3-��q�V�.��Zɪت%�Z��Q�eɛ�Ve���]��T�����Lr2����[v�-*�Z�n��H�ۊ��eX��2�K��d�RRe4�7K\Le���p�F�e.2���ˊ&�����f�mZ55�bQ(\�&EֳM�[j����5
�Zݴӗ���u��js�l�i�����m�pze9���O��$��מ�������zz�9n'�5��-Bݱ���G��VQ�O5~�F5�����|�E�.כ�&z����C؇F� Y�_8��V��g��scط��dq�!Eo���`�dQq��5�1���4�^"!�3��������hbQYl������=q�a���
Hy�gk�����@�B�a�zs�
W{D��\���@g����؁�oȿ��p�[�C��a񲏈X�Dt$y��wd{���F5dz��X��a�6`�N�V�@'i���2Q�3x�4��BLUgD�4�V�o�$�λ��ʳ�:g$P%\vua��V:$B���ޏ{�g�c<<��Y�??�!x�?=w��,���Z���R�І�!�s��X��`�e:)ґ絛��Ɩ~����6F�b�\A}���j�ft�ӧ�yH\TP#Z�#v|p�B�| �۾�����;�~e�(��
6~R�&�w�rB��=����:���?9��]n띹-0����ƆiCk�>��_���OT���q�"&:k��}z��QS���U�<�äY�
#�t��/�M�^k=�_.�Tx�������`�mX��K[ӹ���vw=T��G�,�N뗯����O�^]խ��Rv��dI�r�*�﫴��P[�Q�}w��~���x�E+__�U����3�_��|I���� �B�����uO��!�N��DbF���Ffg����L$�"���wϩz��9	h3�r�lC�H���>8D���Ŧ�z����d�.޴<E��޵�eV^O��r����U��/e�]�;8h�6�e�;��.�VC�f8l�0�D<�F}��ha��%��ә>�LCH�+��I�G9iF�ߏ�u���(��#��^C��C�vg�����WL`��7�h�(Jc1�wnYN�����zN�7����o��WwM\AQ�{�b!�|꯾�������{de��Q�*��C����K|'����C�?j_i�(�訿.?a�-�jcP`�c<��BE?+B!�r��j���H�dq�o�yܙ�b~�V��[��Z�D�j�1@�:ZUTY��ޥ��ű��A���@��W���l@Cx��6|P8q�EZ՞#^0Ob�;�-�[���í|a�H�͕;��+��w����A]T��D$�p����x�o(=k6Y� ��#�����օ�d�b���uY�<d��.2�����3��+2Z�kl�7y�3���Ƌ��%N�]�O�g�o����l~�ք���� ��ta�	,�#��s�{ۯl���?x�f*��"�Q�T$'����C;kH:s��y�F�׬\�0)�ݯ��{�kؾAS�X���"�r
����~���C,�G�K�a�R!Yt����ZC;�ŕ�H�w���9��i���$|p�X�.v\PSPꢚ�錝7�:~Q������!�������l!�|D<l��8�{\���|�`_w1�����n�;ϯ�(#��1��(��5���'�,y/w�APa�5s\�[�쬼c��L�w-����W�9\fwk�G4r�e�Wd�$Ns
	������ѫ�/�e4(�sTxq�t����vkr�C��_�"�x���1Y�>�^��h�4��<5�2�G5<��p��0�Ց�C�6
6@ġ�p��!�"�	;ɑ�ʾ�xG?A��^/?=���gM�j쒧��	$z�)R� ��J�^�C'��]���ԕ^�?K(x�/��l���u���N��j��6~�b��/�*7s�ýy�Q�o�z��,$�fC����a�Vo��ƛ�9��MaLd�����tt�F�Cf���͍�p�zG�Q�n9WTՍ��+JXn�I�&�����3�l=;���L�{SH��	��t埾�|���vƩ8��~9o���1����b�i�V#��B% iB�x��	��X������~Th���iaf�
���	3,C��ll��+{FJ��c�'��,�|D��w=�[�^�#g�lq���!�ST����zL�f�fM�_��7U����
��#@ У�:��7꬇O�#�j�#Zs/V��6X/��-���"#$vTV��D�y�e���<)��D<Ig�Yӄq��i�Bj�?o,x=�W�t�J��Kʨ���:��Y~�p�<Mr���-sig.��\X��hR2��$'�� �ty��N�O�f�����@?�U�,��>#9���!�hd{�F��r��GHe"xW�T�
i�2f7>H",�*�w�˨���^U�a��^�Ba�r�u�o�Ģ7����
Ȣ�/��Q`!��0>��Y{��Z�~KH桄Q�FI�GY.�w'y}�.�gM�!��g�h�����^���޼�L$��s<��CAh2!.��{���`��:t�f��M,>��&`!�~��G�<��CмX�:yَ��Űf�'�d���;�c�Q��᨜c_��P
>��7�F�C���oe��߰�N���	����-�}bK�s�Ρu�.�Ƕ"3�|�Wӫ����Sֺ&����&f`�b�Vt�t6w��ɣΕ;�+-���y�h���6W���W�>�9.aiwǌ!�^�쉩�s^�cj'Cd�w��Y��] ���/�dH�����s3�U!�haӻ�n!\�<Y�exu9���b��G�q�,��U|��*�7�*#*�nmhq~V~z/�c~Ϛ����=�]u�`�fz��*Q�9���val�	n�B"�1g��Z�����_i�*��Gavׯ�,�ִ�$�ț��#�:EhwG���a�b�خ���(.eɹ���m�Ś����,��eF�����y�i��iw`�j���V-Q�e$�)�#�{fN����Ш_k�sSÌnl�����������˳7�Q��4r�\i�ns��Fl`R�j�欭���C�ɛ�ײ�vK���������8����5�6��/;�P�$�2f����v2���^�n�bUh����1���0���1+�q���[�;.s}w��|Z����r��B��"2�I$��U���I�å��[��u����|���tҦm5g��9�<�z�9��&`��f3�H^U�wQڶl5���/�񫝶�d�ܯ����Nr�"ܥm�
��m�V5��%v50�oU�y���Ӂ��Rv�e�u�l+�\Np�z�Z�ķ��8�d�^�=�'V`����X�%/��oZT���%i�_E2vn�F����!�΂��PSŕ��Q�>�S����D��T�u���L�K��Js"�����0i�X[қuɬ˨"Y��ZC�h�r���,T�t�,�������[ׁ�,E�r�e��WJ�꽓�\�թQ�;��Ѩa�� y��ٹ�?��=�`�#(��U埰�1�w$�*�v�]E�q]k!�Xti�e	�qWN�_Wv�_E�0�-rJ%�PWJ�S��䴙���/�M\uU�� =��XW]�5bGh���=[4��n�ui�)_1F<>�#g���Vm�@��;0��9S���QW��z���VK���:�,�N�k	�,��Vʨh�%�A�q��n[��awوv#Wӹ�d)S߮��tZ��)��?�;��l��i�Tԉ�0��{4Z�e�w���ǔ�J^��"(�3"�U�SL�Ƹ�V8�[n6*����ʊe�A�i���@�ʢ��DKaU\����d�9�p����˃1ı,F2J[�v�j�*n�fn��hhVhJj�37�.]�X�YC��U2ܵ\��Q2�J����`d��e�b���k16+UuJ
���(��i�.����S5���1U�*��;�2���k]y߾Wԗ�fN�l�
P]�}ձ�L�9���}Y8?B�8S��P/H�W]�w��w.`B�A�o���b� r�c�a�1���]��.%BB�򩃠C�:\	�Y!b0��Ck�h㕪]6X��.�#�;=z»����S3=w��B��f���#++Vc�<�V|0����AF���a��a]��vx��
r���9K�mB�o\�͛޵�{o�U�md��TUz1��<�J�<;����E�� ����ֳ�t�r�S��==˷��Dj��=]^	��Z�U#���	G���%�0Q�n�x���͏"rR�b���͞Zi]��r����b+�y����y͞O�=��ya�zda�]�z�ʰ��WpgT��Y�<��%&�!B.a��'s:������
}MW7�e��Kt��i��{�z�O��w*WX��ќ�b���$䰗�i�h��[2�N��+b��R��	�2Җ7vH;�Z4C��%�WKVF��	��y%�'nc�g}��}׬�F�=6c�c:�H�h�H���𮔠�s�[G���8烞u+���Icx\�}p��Ht���r�WL5u�/r�z�f�]���F��Ê��:[�ŉ�E_Y�y���"��{��^�0�B�@�0[��"���r�;|8Q>�Þ�}~ת�n��>%M���?�sһu�P'9Z{V����ѹ�U�1�}�(�����;��u��KW����S������ᛗ���E�Jܱ�K����S����3�vM��$R��\�<���)�]�<(�.����y��&5�}��먁�w*wt(�0��Y���w�x�[#��Ӟ�w��ik\��y�-G:j����嫳"�ڴd�����s}ȵ/k�%�V��i�����-^J U^�3�:��m�Ժ�r�N@���Y�����9��2�WWWG�D�ޱ+O>�@C��Gq+U��د��MB�� G��w�+��YQ.����^��J�A[P��v�ଈ�qy�6��.%)�0+�j)j$O�dǻu�$N�͎y�#^�CըK��e��@�KĈ����1�ύ�Kz)�9Yae�Tȩо�>�g+�(j[u�T/l{�w���0�__�iu-�7�DH��W!Q;{��)N�=��o�V>�]�(lW~җ���	���J�Ǣ;y4D�,[�����:�����t��9ѽ�j����K�!b���T��<�9�L��}s),�霶\=�n2�6�N�����kC����7�i�	{��wq۸w����>W]�4W����F�r���l�Ƙ�!>��y�|G%��+�<��3�͊��C���V�@	�����-W3qz�eH��<Ij�py\;�-.S�jr�I�ں���{������=�hz�#�{!VZ��u)H�E�9MoT��y~P�>.��~���`کw�W�$��H�2Kţz��i�
���fs�����Iݶr�kr0�i���]öy�� m<UY<i���i�;9�9.���)e�S��u`�1<�z��%�6�W��{�I�|��H���;�dR<�׶
U�Llų����Ic
�Ӕ'��v�h�}	�����b�;:R��{��ۡ��yHTwƠ-[����nUQ��w�v�A(Ip{i�ϸ�R����OU�풟v(a[f�����ÂO.cE�y�L<yPw�#^�v�2��V9LO���Z;���a�cPɻ��}��1w�;��s��/��f�%ߙ��Oɠ�+�V!.�q���������t�$;ч�Ͼ�H1�a��I�B�'�۫��zȗx�������l�w[hWK������;��G��{�"7�l�Ci�{��H#x�FE��c��N�X6�-�
^[�,m���뷏2R�｣;������wk
5����ë{�fr"�cs �ǭ�<M�8�!!F7�y�}��uG6�WT�+[y=J׮2c;-�E��{ʸh�}'�:|2��=E���*��S�_��Jsp�_�����Gn|�1��}��{�o��q��/��Ǣ���N�;U��ۼ�D�땽����/Y����f1y�,m<Vq�
�A(_P��h��S��W�+au�/���^WS�8���\߭�m����o&�����5�YuU^D��v-lv�T���R��_x`>�)�:���9t-�{�X����ҫe�\=VV��;�":�u�6����m��y��*���KE�;<���ꃪ�`�����_	������-컛�1�8͙�Be�3���e8��IB;�HІ�g(�6�!�_Id+��c�P�C+�t�50RLne	�ǖG.�|�J�Q�J���@�̓��W�<�J)㙣�T�!���Ńm�����y��.��;Y������N��2�ާx��4췑�v�헿N�1E�����E���!w��\�t�qZ���u��ɥm�=���{G���i�(�y��F;B�:�yc�S�h_�5s��%m�H��s:uG[HA��jvUv�F��{7S��>V��'���\Wp�ɦ�kX��n�*��u
�
+��w�ײ��$��hڞv��9��S&b1;v����vicUp�6q%���_G.�9>��`�N�M%g.$N*j��K ��Aj��NXO�t&*���܉�*��J�:����B5w!,-Cm�t��q�Fٗ2��!�����L�H�j����(��m"k ���+m��餬;Wl�@�Ŷ����XvC!۰�=��n�� �4�j64q��t虒���@�dFfeb%Ջ��%�kb n�?�'T�¥;��|�$��
qa��]����<-�Ԭ�б+(�l�\j*� ���""((��L�
%����f�f&[R��L�#FT�E�2�-�q�+bQݢ��)j+5���9j0b����E*���ҰQH��1v�
:�b�`��ܥ ")�ZX��a��ɂ���V��sW;�g>ng�߇7y�v`Ab���r�,s�NZ�[|��Is7��;a\��W�vZ#-���g�f���|~wYSq,�ɬ���o0'M�
�x�+91<�۩�jⳠ:���g2���unW��W�Z�{h��uSt�
���R��b���Z�Ժmr����(4�w��7uOr�eA����yb�������n�l�:нy^\i���K��6D|32wDpn��sz!���&i�9jC������I�B�M��@fĵ�<܆�Oo�IG��|S�����TV����{�t-�S��:����%�B^�Or�ۆ�]��'Y�x��ܰ��%6�1R�(��h2��ǐz�-
�f�oMPM����	�WY��H�J���}=%l<Y5�t��W���|]rLj�6���݇T@�z���x`���]&}���҃�I:ƅ �J�m{8�;�����n�[ק*VA}{O*�-[�3f��p����)�RY�r��53;�����&P�����s��{rI�nS��1sjV]qMV��p� ��`O��n,��{~��֭�y��B�l��~sP��x���Տ�XǱ݃ �cd��ɾ�]��ͳ��G]�u*\�育9R�ے!֛��/@pJ�Ef�]��҃�R��3�\�̑^R�����d"ӓ�G��@�ļL�h����E�C;�v�ץ��hZ3c��ʜ��K&�Nwl;ڠ��w���wՕo��*\�	�ﾯ��C����@�JnJ�Fm��&D�ʇ�����O�ֳ<gX'X���Ǘu��d爚}��&�)p��{��ğ]�yς�f�������S�`C�}f��\Y�����|�	�eN��su�s8>�-��f)N�t'Xu���X��= �*�v�؃;ݰ�l���+A]aovy�\5�-�{X@@������
l����`��V�RrjX��⠇����梅X��u<N���-���yGApj'^[�g�bq.b��h�Z�~�h�ϴխ�@�}�·}=n���h���^��<��ტ�f�W�賮�c�V���*�͘�x���ņ�{�m�8ֽ���1u��L�A�Ý�Ge�K6f�jV� �=�k8J9��X����P������2>���^�y�q,պ^ܐvN�����6�f�VM��$��)�Z��r�j���G�n�3诜V�P�������-J��zes�н�s�n��[����+�|��`.dιΦ�ֲ�U��d�oVl.[���L�8}�F��|�a�VV�}�S������o,�Ts���wZ2��H�
�뱥�6��;����jQIh\kF��'��X�y:~o�Ҹ-/x�U�7����xbUxR�6�ʗ-/-}L�F�L�OPJ�LH�%��5����w�����ẺW=2���y��fr��k;ֻ#�i��r��˫�q�7T����R+�0*ϨMB*��,���;;ӭR��,'���yY�jqū(�>|۬�Mu[աq�����g���\�ȞA+�v�������|ޢȀӕ���H1Pu�Cqٺ�qU�yڣ�����Z��#���\ecz �;U1���:���0�r���S������'A�.�-#�:bN�>՝�3|����\�n���W|�y2WNޕ�㸹"���R�+n�����_�}�}��G��{w[�"���1&�q1�Ǟ�v�,L�V�c�(�7W��N:�aG9C�坞}�&:���;>x}�������D:�k��e���[��\�(ymY�2��*���$���֝��p�����byob���Z+%k�w���s@�v�6���>�:�}]sb]�����,���v*s�=��<�a�s�!����xv_��B3/��
ǶUQ`m��;]��G�UU������
9lb���]b��9k��sN�I�u�9F�y-�^ +��ֱ@oF�y*Ν�|��΃�KK�P5�q��u��5���Y��e���M�w�8��~AF��T�mm﩮��:�뎵]��9{i�r������rO&�,`��fyök�Aİ�DX�ޗyܡZ��<}�ݵ�˟[����tx����i�B'kgӆ��ox��f��Ic|׏���.i��0���46Tv6���^� �_o�����}<v�ʃ3� 
&���[Z����05�-Y��B�=��;50�ҴR(3x�.�F���c\�نn̪��>��Щ��;�qc���b!�[����+���~D�B�$�^�3k(Z襂ڦ��ɩ��2�ص9��䯮-R��>|9휧�w�Ou�¥`E�n��z^��S�'CڑvVt�_wX�]|W-.��)�Gy�u������ۄ��qY5]H���6w�9n��&]�w�9����k0d���AXiv5z�����,i��:�*ڒ�f��茿�˻[��z��E���)Y3�M�#15�v�G>܄��k(־��@
�|�h�C�w�Xs�\�(+�Sԍ]���音XT	b�ה�E�b7�����ڣ[�,X7]��BLp��V0HDm�&���ܻ�);lZ`!�6�X����J��b�9���("��B������cB9p+�l�u�B���*��J+nɠZ�Fm��#�U�DX�t�Qܻ�.��&la�/("M��e��w�~5�@E�B�0@�,9E�2:��eVQ�ǆ�cw�@"�AAt��c�P�Lb��
pL��Y6bS�u�*�G4n���^��V�����ei'Z����F�f�����b���HE�q4ɻ﮷���Z5���%AwiU��%UEb�"��D����
�#KeiAEO�Ld*"�b�IYZŭAF$X(���-�r��Uĭ�X)�TU�TU "�#1�KCLȘ�.�ődm̱E��*�iTd���1R�Eds,���b�4�,P\I�+q*�R֨�R�e������0����$H�;.)��:Y��w3����5��?0+�:xn��#�[���=���'=�f�VW���F�|���e���i�ތ���f�V�´��|�`k0��ڣ�6���+���I�x�����r��6_]�w��V]Z b�����"��=�����i�=�r����6ٚ�w~�|%���6`���������1�G_��6�4��w|t��&.s�����t���¤���w$�Z��(�++��J%�,���B��=�ì�Ϳ.5�9G���kT���	�ꩨ���.=ۯ�7��q�kD��R�Q�W�R�:�%�e���s�WZ��)e? ��n��zx����6%����y=�f�aG^Ŧ�s��+�5�%�ۼ�In�Nul�pXE�q�m)��٬Ȝ��n����<j����t5M>�M�t���x)�Hoj랖v���u�W��)�出�ܴ�U�]�4xk =�c8�`f�/Ըt4=�N������M{ôFB�x=�-���I꽂�0��f��o�-�]����_B|��"��MP�Q��Bz�%<��{�y�
j����'}l#��RZ��e��B��3tQ�(n�t�9�ax�Zw�T��������E�u{;MX�[��o���p4f����<��gvr�	&�Ï�*�+�����v��5��}���}���T�}���Њ�F����,!�=M��^�)���)�{'���`�+�nֹ�W �j�o�p/k5��\A�wn��P��2���U9n��^o�'�K���<Ӑ����	�m;�u���$��<�)��@�s��iݖ=:�9�A�
��z,;E��� :;| ���Vﲋ��&���DsÊ�O]�)Ζ��#��pP�ڋ�α�s�t�S��ݎ<�����"_�Р��6�f�<}�mfj�y7AĠ�$�#j�-xŎ�nTSL��\����C977T�}V�AZ�է8w!����ƃ)�r����K�P��������
u��L9|<��
�tTaN��d���*�5'�7�!1�Z|*�}�wo^;��x�+a
d��Ty����ba��2�bIa~���aR	X�Ì]wZإ<�h(��zNU@�ƷE��W1���h�;��V����b�}���W��T���m����%E�z�X�{4��چ`�Z�᪞V=�Ԧ����D<����;%�&D,={B|�}���\^��^4Oy�n+\�y����t��c|�]�
��}7�t���Q����Ɲa��%�vN9���61�Z����>FKK�l{F��e�U��1��s���+Ѱ�Ec�y9���L�ݒ�fh�ֽ�@E�$���������-t�ǯ����/8J��y�Wh.��:��·N86=��jy#^B��G{��L��=٘Ex*l���3�݁�8��30��i�a=�<"��#�	���d��De2�Llо�����z�[�<:�Y�ʥk5Wh��8ʸ�#��F��:P��)Q͚���N���圝TKǭ<���[�{S���v�F�^�4!��b���7	Q?oh��[�s��WaZ�n��S��J@���at�ۧF8+�]EP3�!,�\����2_%`���~�o3�KI# Ҙ�T[٪��*�F[k�'6�S	=����'p4����9@7���'۲�v�Ǿ��z�'l��*�
'�������C���'+�q�:˻������۬�[k�,�b�@�\څ�Cح<��i��y�vĪ�K��rݛ��_@י��[bV�i�q�:��j(��ڤŭ;j��'��u=�,��M=�<�y���֏YWFi�:�U�

�,��#����~�G��5�{�B_?yj��7��^��wʟ3�D��<�n�y6�gz��
�7�wM�õ��3^���w�L6��O�k9�	�\�3϶���x2���p��&>Գ���ۦ:�Q{'�>��N���9�����g�'4yU���v�g�������>��Y�iGIV�x	�VS9f�N����/�
�.�L�s%ǽ'��q1�j�K)�:��r%�u�9��l�wk-6���`�D,�4;/H��_J��Ǐ�A��C�Z�ډ��v�he��<��L3��y�Fj�[^�O��+5rTe$�kp!D�4�j��!�/[�/;3�;d˯=�=���u3�a���!�s�ud��r���!*�]���Xr{�8Q�o ;�b�)=�7x���vm>w79�.�q!�eۀ7]Ò��7e-�T�h[���s�fe2�$wY��zr�����(L6u�����������R�r]+[��\�+U�~Ů��޵��͵��Q�q���-C�v�5��T�Tm�Ч;��mp��W(���9H��x�_6��	�j�t�c]�X�p-El\o
������D�-���,����ݓs7:x��
!���O[l�l�1�hcγ�(��˸9��2ݖ=���}�++���j+�w-ѪS�Xbͻ[��f���`&�e��S/U�ch�0�wu��8�Y�IJ�W|�Cb�4��$Z����*%+�$DJ���.�GJ૏�]6��T��e]���Yi��A%�x$A�$d�����]Vr�P� ��X����^�R,-�����DL0��*�irӶ\���df�t�u*��$Z-Q�॔�^J�nȽ8��YvK¶�x�SnV��e�K �Z�ʊƥ�f�`�i�j��TL(�����aQ��q�JfR�5s35J�k0F���r�F)�(���1�)E`���R"��AA��֥�M2���Z��#�f)�X1
� �ŕ���h�q�e�*�f���$��!
����U���캵g���K�2d����֓�g��5����]Ū�w#���Q�|�j�i�iF�uq�Z�� �8p�T�[k����yIT�P����JڞU�}�Od]mţ�1��]W���Kܔ0�-�)2Hc.N�98x$���qk%��(܌TN�&C���ku�^�[�����	�;���N�"�i`||G��w30;�������
�j�[�5���7g�����'v^���B�Y4t�Pev�mZ��7��c�z�v��woF�ƺt�.���)�����X��ߙX�oٖ�$���R��W�N�;]��sޥ� �Q�塁�{m�[�m��� �:.��.V�͝��X !�Uytw>u0�쌇��D��0q��y��[^�0���^qRZ��Ɠ�]um] ˱]���=���<��Wzٔ�+��c�7�0��^��1'?O%�-�e*��9�<�@T�
Q�*k2]W_r7���GF�B�ͽnm'Cg���=���3���i�ĝ�Y��o��i�^����k|��7�D��Xy�]�F��g��.A���
�'��}[�Y=���.��]��;g�b�#��5��]�j���2�d�MG6�������)N���BncxpnU�B>�:�R�{/��e���N!�Y���v�n���N�)(͉��:�r��+��[k:=�Q�[��weG��Ym�~3Q�B�ژ���9�W������ާ���F�6c5mqm�9=��Mu؂;�Z�<vo1�s��ןX�{�.j��~��,�!W��ȠӔ�\�K�oi��V^�n��8Y�Y�5܁�3�V�A4��[�Y��/f:�eކ����7v]��g�ϳQYy�Yvq���������:��a�}\�B�U�:���3o�tv���m.�"��퓹V��Z����5$�R���;���_�c�j�\.�Z^l�9Y�6�vzE����������u�)��p�=`xː���{$�}lC��^��BT�hb5�x�>Z�~��u��`�����ј��JKԲ')Ő���-��K7+���U��35
z�c�GTP��t�U���sT>���Є[��n��d�(
u�sz��K@e�Y�3�Y�K��gK"�X�6��ø��^�+{�����T#��n>�ڮ��I`p$�1L�I賏�f,�EEy��34;8���
��7�~+o}li`i`x <6ҵ��K���v�/f�sG�}qA�u�ux�����f��<Z����<�g��v�e�[��+Qh����L���E�|d�@,����;��3�;���|���m��;����	r�R�<܇��)vC��x�t�QT�Xe*��=�0�c���"{�C���-s���L.�vҳ��40ή
vF�ԙ�ki��W�p�6Y�7�'oGc�%�ע���b��N,�d��=�|�\g0|��j��;"+W%��_�e,��۫�7%�(@�u�{�nN��*[� %�Vʎ�\�������Zػ�]��Te��ק��T��H�p���e�͖j��1�c?P��,Զ��ܞw�Y*�ݕ�Q����5���Fx�^�"|�;Pw���E'�G^��%H"�N��}o-7���L�Wp)ƶkη�\o\�=����(���m0�.^���+n���=�w�iфܛ�����jۍi��
#Ƙ0��0��$�Nn���3,����v*��~�B�0w�5{7NV�!��(^��FA�D�;M.|�(f�Z#��>�T�!��λ��ׁrȽ��rm�y<������������>Yx�nL!�����ʆ�5�&��t���u�{�a���sZ?�I�?90��O3pBY����̶�{	^+yW�ũ�qf��7�iuyun��+�K2��N0�g��{�L��s�=��:��R-M��d�/(�AD�]�LӞ��n^���ϼm�r��q�76%�W��q��r�\�yT�d|Z�{�wuX����u���N��u��/���b���*��<��7|�ڥ.�{)�MqݡgDb.<�:�8>�U�8�;�+=�,�}�Q��
�k�˵6�-�w���C�)�K.	�z#Z��ȷ|ﮥ�s:�o�O�0r�V�Χ�B�����
����-ڶ�֧�͖i��A�6M���ic_2��0������Y�ĎF,�2Z�Sð�Ƕ?nӼѩ�-Ì��v�	�>E]�j	�+�nVIy�/o�V��t������z�;,���n@����k~Y
��3Dۨ؛j>Fu�^�U�?��6�!���&'E���M�g �˾�pc�m*��b�7O��[����.}��i��{vp�Y�Egp�*��h��Y�d��q<̭o)�Л<N_��Tu�:�#ՂmK:2�_v-;EQm$��X�g;\R���,씌�ग़ӵ.^�Em��c7���+SA�|��׫�UN��(�[]��a9R��r�M`���o.kU��k��%A���8�d��H��֮�S�4*��´���3��U*�P�kVgk	L�|�e�o>�iZ���DݷK,�{��ןoz�efmdF��E�0���"�[�d�}�vxx�Ǻ�&��>�X����r�k��ge�.�wq��.��jS��X��vA��f�ǹLoa=��T�t���#.M�I뱦ó	��hp�|^��&P�O�)>����;A6H�Y�S�a�����{�kL8��C�Dxgv��V��u�~�Ħsُ���xk9��;�蹅H���l-�3-�f��IAu����U�ņZ��*i��!��+�"��W�8��WM@Q\j�E(ʔ�WV�CHWNfd�ŌE�X����YP�cut�Q3WC#��X9nX���P��T�%kY.�b6�u�E����o]�O]���֫���ܱٗ��>ql9ٓ��\.������z���mv��Rf��(���"i��s;��o@��f.^�1pӾ��\��)˰���l�"�um��۱\�uE!�b<��]��S�Z��N��~^��J}ςE�;(�~��H}�=���=��9�$iUkM�P��\sp\Q5iF�-��T�r>9R��(�}wL��M#�wRs�=�I�d��|,���gfub�[rw.K�����_;~�w�Ӓ��mb�l�K���溄C"�SG*�$��qm]՚S@��չ�Jӗ6ڬ�(�����6��%)�hD�`�׮4��+�c��4y�9}���Rg�B�i��%��{�\ݾ!D���E7q��כ�G��{�+����=�o=�5P�y���@�,����՜a�X���1����T�s�;Q}ȳ�,�.��\���.\���I��}��`����>i��Z�p�2Q��������dT�������q0�X���y�}���U�Z���}��XB�H"X�v��q�-ܜ�lyfu��M�4Bp���\���L,���]�WS��dys��y�! x�5��r>x�G�`er_a^������bW	o�;�p�,��|[wr��"{�i]�X!p�itL���HN������%[7*A�R��!���?-O�q��vE���S��;��R^�n�s}Aw%��@��9��r�潙��*���Q���\T-���T��a��
��q��:��z���]g����q�\�/D%J�'iLcS]kE4�Rλ`��nx.��um��)̓���dWj]�L�����._G���fN��</:�]��9��|������_���F�Y��v�^d���Q�G���<�h�xG��[�C{.QK�謥� T-��`�[���ԅ*�������E��H�2�'����Ղ����k��T�,����Z]5���@ٞ�Fy�ɹ�j���s8`t�j��'��ݩoT�+'����)�SH-��'��鎸���&��E�"xoܱ�sk��ut��oo1v�[�A��B�/<�|�sπN��rY���6�� ��{�*�Mح��&^Q����1�{/<�KX+���ߡM����L��]�g+�:+2��S J��͗(s�%���쪫����M��ou��4h��ٔ���W�vxLٻ�p��jӛ�V�;<Kw8�I��f`��I��G#S��hvo��"<���tDu�������z
q����GI�4�K
��AWel�+<-r3EBs���7�	]{��I�Y�BWPT�N�}GC���K C�Y��n��~C�&�99G�=���٤�8V�+2U�c>�p�á�7�*���\�Z6�	�8��6��0,;F�U�3x�_i(h����O])�y}�A[��5W�_I/�u�9�ov�>]t�+@E��lN�m.�o�]Ӯ7�7.���]wDT{���0J駳�QE��*��2"Q�Mu�dþ���
�w{�o�HWKE��Lް�����p
���	�a�')c��V���%S\:f�xa�Y��W���$PңI�<uc�0���"9�U�*��������)[8�e�F�7�̂���i�I�a��Nx��6h,��}�i�~��X�2;z��adU��g��À���g^�/Z��#.M��Wc����3�W�۷����f��e�3]�]��ݜ�o��s�m*4��{�s�^��{�2#)�0sxw]��s���������Ղ��ά\|֎y�A���zV��z55-U뵔.gv�hwZ���B��罸	�73M�T�a�>c�n�ݑpo�����������Z�؞�����0�iC�2pr��Qú�>�C3x��O��{]���o\�ݜ��DV�X�	eζN�͈���{}bd{0�/671A�ݩ(s��ʬK�Ttw:��ޒ�f��o�7+�{��+�<a��It��e��ڇ�xk�����uc*��o���(ʫ�#�&������02�(�4*ڔ�]WL���ƒ��]�ڕB�8������������� I˥j�����I I$����$�$���2"��f�C����(�6%�]�,�O��M����z�I�B@=@ ���]��Q�A�i��"�`OV�a��Q�Y�)���PUN�#Tey����}v��9���>sK��o�w�4�.%G�{�Hay����#�hJŊz��*��~C��x夯O�`�&�AS�7TET��x�	+C���Ey��Cx����|����L���l����8�
��c��~�z:�`��0�����w����d��	#�Ib�����L����f��ӛ�j�*=�`�ӑ��.QR�\��-��j��\�,�
��Ϣ*Ɋ�D)��ZmD�B�)�y��7MY�Щ��*
��.%�$�ߚmz���[S�=��$=���*�pD�N����O'����_�}#�i4�dTR�l��`�CԚ��G�x�������풎�$	pG��'�E�:�,E�j���u➍T҇6�����l9"��k1����~�&�&&-�hAޒh��`����UK0Q�T��oތE�p�����Pk��=N&�E4�_&���\.k)@@����)3�

�AbF�+�� �6M~�z{��e���@�zL�{��0�er�����$>UAU2hf��2WroET��H}R5����	�|4�ᙣi�O����X�
r��J��
��9�=��'�x�w���L����PUN������F#�fI ���R;QAU%|��c���<̶�Ǘ�Bk.�hj��{&7�'�9*A �q�F����� ��@dC�~;�<}�9�H���(*�W{[&]AM��)�xԺbA݀I��[@כ���$Å�v%���zR��� HET���`��<��#[��UN���]7����dXB�S�T�����zB�*�fi=��rE8P�C��