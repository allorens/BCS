BZh91AY&SY��k��߀`q����� ����bF?            �W�*��j�AA$�Q��f��em2Qij����d�ba[j����ƫm6�i��!��V�dRس[V�-i�e����Q{4�Ֆڭj�fim�C,Ų��TeIel��%!3X�X�lT0Rȃ[X3F��6a �����&�2+V5-Mx �P��[TC5� qεUf�ִ� �T����dEfhdm�4Z��B#-KKj��4ժZ%6M5mZU���Ml��Z�[4�������%v�  hs�@  �/_V���6��u&��wM;v����6�K;�֕t���wU÷]�d���Z����Z;�.����uN�Uѣ]����Q-��ʫ6�T���"�����_9n�h*T�+�5uk��J:��.���u��֔�j�(�PҗU���3�ҥ�l<����@<�cZ5D%c,�c�k6�|�  ��>zt S��{ǧM��z���5O{tUn�{�T{5 =��\z*R��Ǯ�4:�tJ(y�����&��m�e�{G�Za��v��լ����-V���   ����>�m�^�� s�Ov����{�u�G�3�������u��Юq��/b�����((�F���^�T�ڶ{�!��#Z-c#*2��|�  ΁�h(����Jz ���T��V�=��A^ڛy�/�Cݷ�E{`)O{�=+���f��S�
V���C�A�;=��w ��mM�ZٛX�jh��hj�>R ]��O����9z��;ټ�(hꝮ�`2�7P��v�ݶ���=���u����;�ht����U4���w	�;�����,�*���1���@=��� �Wp ��{�z
��u��Ac�o  ;z\  �L ��q�u�Aۃ� mv���X�le��&�6����� ;��C�A;��A�ͭ¨룀� s�  9�n h@�@�8t����h��: 8�u����k3a���Mo����@y� tv����s�pӠ��  졊 ��9ƀ.� :ns� ;�b� �wkD���i����5���LV�f�}� w�� gF4 i8]�]��M�
�v� ��� F��������B���Mh|          S eJ��      "��Ĕ�*0L��& T���U?T       jx@��T��C&�i��%?R���Jd`&CF #L&��CjI$h�SO2�Q��$�!��������~�5���$ o_�������;�-��]�Y�s<'z�d;̞=���dV�{���J(*~���vC �
���	�?���?�����������V��I=��@_��qCЉ�j'dQQ|�_�������)X�`5�Q��+X�`5��)X�b5��X�FX`5��)X`���X�b�`5�V)X%b�V	X�`��V�FX�`5�VX�`5��)XcX��V)X`���#X-b5�VX%d`��VX�F)X%`��V	X%b�`5�V)X%b��V!X�`��VX%`�1�V	X%`���	X�`�V)X�db5�V)X`��V)X�`���V#X�b���)X%`5��#X%c-`5��Xb���#X-b�X�b�bb5��#X�`�b5��X-b���X�b��F%`5��X�`���#X�b5��1�V#X�b5��Xb���X5��`5��X`5�VX`��b��)X�`5�`��Xb5�`��Xb���X�`5�FV)Xb���)Xb���)Xb��X`5�VX�b���)Xb��Fb��V	X`5�VX-`5�V)Z�#�R��k�B�J�+����Z�k��J�k�F�J��
�+�R�J�k��J�#
�k���+�R��k�XĬ�J�k�R��+�V�
��F��+�k�F�Z�k�c��Z�k�R�Z�k��+���k�R�Z�+1J�k�F��k�R��1
�k���k���+�#���+��J�k�1+�F��k��J�+�h5��	X`5�V)X%`��V1�V	X%b���X-`5��XV	%`5��)X�b��V)X%db��V#Xb��V	X�`�����)X%`5�V	X%aXb5�X��V	X�b��V!X�b�VcX�b�V	X�b��V	X%b�`�V#Xb���	X�b�b���+Xb���)XcX�b���X�`���XcX`5��X�`���XF+X-b5��X�b���FX�X�`5��+X-a�b5��#X�b5��#X�`���1�V V#X-`5��XX�d`���X-`b���`��� VX�a%b5�VF V#X-b5��X�`bV-`���+X-b���$b��+X�b5�� VV��XX�b%`b�aX�V `�� -b�� -`�*�b	X���V(�b�*�`���b��"�` �X�5�b#X
5��X(5�#X"���X"5�#X�5��X�5����5��X����X�5��X 5�X���+X�5�#X V"���X�5��X�`���b"� -b��
�b��$`�X-`���)X�b���#X�`V)X-b���X�`���Xb��`��� V(VX�`5��#YX�X-`���+X�b5��X`����#X-`���#X-`���X��X�`5��#X-b5��X�	b5��+X-`���#X�`�-b5��#X�8�%�}�����w�����[�{�!��Q)�.�5���z��PZN*�켫Z�;�+�m�����y�X���1���`�6��/N[	���)��vU��F�` �?,���Э�I��ܼ,I[ �`ֽ�Zz0@Z�dђ�TE�v�����
��a1��œuO����t������I� \N�ܓv�L��j[Wj��i�ףrl9nY�q�L"Z�p��y6�+&&�����\�{�*"bmV�Yv���U����[0M2 �\GS1�\��Jȣ�^��qf=�(e��;Zb�#*��y@��N�ãNJ�t�+yJ�ݍ�O Շh�.�<��۬I�EC��m�v�_=�to�/-Q�6S�sX �2����
��ȥ�����0D�:W���&�<�DM���`�bݺAU�g�<��;��p�yԖR�jn�9k�[Q��,��B4�U���H�+4RRY��21k��mn��ݔ7Zٓ) ${����L6�mT�Hl��K,ښ�R<o6)̵�OsD�L�U �t��6:���*���ne⛻0�#�)M*`��N���`zsiM��3k@Z�Y����`���m=Ǎ�e����.�Ѱ�h�*�\be��f���{ô�nm�l��cn��:��ђm��;�b��n�A�q�V�E�Ԏ[r�c���͔�7� �.�Jˇ:��U朄=���N:��x�#&��Rd^�z�F�)\+)K	�����\�(�70��
ك&mքj&� nU�w�N�RXͬ�� ��g&��=�#^��YX�Vr�]d�Д��[NyT9��WF��]�.(NHɚ�Y�on�JE�B=�b�n���gb�m^�E&�nLFh���6<��%6�*f�-�i<�v�X�Ћ�AV^�mn�p:�s�չ���,�{+ 맓%^�z~W�*�S��	���PQ��w�Vj�BG�l����1Q��[P��֬�컴���{�.�K�Ea�u�GW�&&�Æ�n]������v�˛"
f3�"`]1�ى�*��m\���W��i�����7Xsr�h�1� �q�O�َ�:����W�͌#�lv��E[8�
�8�:�sB�Zi��t�-��%�D������3����ጜ�z��a�V&�Sݲ4��	|�Bi��a��hQ��Y�����.��*\�ř-��ť��f�2��\t�F��n+�*�� ^�*� ��
el3][:a�Ҧ�W�F�lm�Q���j��J�mf*-c5Y��l��u=����!�-(l嗹�{���h�,=��Oh��v�@޴�̍��n������齊��ͫ���K�f<��8e`�wW�	����h6��ǴĻ�7C�k�ut��SV�㳳�6�f��!@�ۦe&���d��s1I�ܕ�FMuk-������0MT��,��vD�bvo�g74�׮Z�qn��gZ�`�.��IJ�D��X,��u�����v�=�{Z��և˔�h��F]���&!�7fB�;iKUYY*ŗ1�-SMJ*ى�;�}�E�!����Hb�ζ�ٰ���he;N��*\���kC��̔��r��*���;l��1�T7��\ʧgj\���wB�ƃfD�TԲlG�<;v7RhKr�ņ�^�2k�R�/2���	Cu�z���o&G{2*�F�YfU�1�e��bE+M����=��L�SM�X4���P�Wm��5�H�^!������"����&��Z�2�8�A����@��#(��*�u�bi^�&1R���fm��Tlk�]0��d*;fi�����m�K%i��(L�,p��Ϟ��3���&�d�r˰���VEl�>x�Cfc��!�z�H�5V�4�je@���D�aV���B��Y.}�0���u��� bI�-�j��>��6"^�cԛ���9z�Ȫ��ne+�q�V<��Z��7�F,fk�y�L�3N]�R=�O!�е�l8˅Tֱ�^�TX��ZIE�FK�u�wDmn�:��%MQfTa%��!i_�E+u��X!�L�W�.<�;@	���h*�bjm�p�-[{�rKf���%��E��2�^;�֨v�����~��}h"��
�#;B��9C#*:��i�w�rb��_��v��ǳm�cq���xM��-�r �Lm�w��V�B�y��а̬�q��g�ϱĮ^`��6��dd+�fZu�����3�dm�8/��p��M��=��mQ�#e�.��-:9,QChf�vI�i
�uja1��µ�6�����-�Vz�1��"�Tgnã(S�]��4��B5^3#���o���U�����dr�k�K��TZ��4*r��f7SdA�[�6�l��웗�)�����P�>mҬO:�B����)Jc@��N�j�-�K)V� ��Hʕm�T�@��$T�+�GB�M�l�Yj�7�[b.eYŌ��|\�J�w���&	z�$&������U�n:��Kˠ}���ѩq(j���RDPb�^��
�Q�`��c,P��rW��+b������%��6ɍ�Rj�Օ�5)�J�m+ٰU�Y3���xU�D^允�Yq���%+r�M�7Ton8t3f�*kKt*�0�	�ȴ4l��ʻ2eF�zD���] �.���&�e7y-���T�b��=͖���F1��lCc���"�10c�E�q9,Mâ�X�#w��&ɀm^VH1ZTā6�2f�q����Y�0Bѳt[(`mX���;u��St���+����)�f�0�,D���1�b��'e��n�2��V���d�@��Xn�a�3dJ��j�AO�fR��n;�sMZ�j���oe�)9K(�Ǌm0ţ��X)nfx��8oi�s�z�O����S�J�B�;.��hE��ټ��ea�(9eb:2�]=T�5�;�Z����)0Sۼ��{x�8e(�ɀ���S���tkh�W�ؽՎ� ��U��b���\�7�d"�P^K����V��uX�Usi̱)�j���^��@Uj�lʳ�i'��vn��QlK�k��D��b����5�M�j�]9+��O�N�R�a4Լ�0�Y�22*܂�zl#v`�/q�[���7i�T)�x�+4**�.M�i�~3n���AC�F�n�K�3�k
��ĵkA�F�;z��n�iޅ)ԗ�0�u{����N��N�ݒ����O�c/3iZ\(IvȘ��{���X^*E\�����676!��USZyѺNkN���-޳���۸��Y�C�8�Pm쬺�A]�Ȧ#�I[�]ն��X
8nF�õL���u�]*�n�ad��[h�rI0�,��́ĵ��Ehçv��L���70^��Vܠ�]��t�n5��:[�C7��$&�g"R�ve�J�B&%��d;a���%DI{z�Mc�MJy���\��\�s`��;���Zޠ�]�)�͘3s#Á���ɸv�ڔ
�<ͺ��un��Y����J,
Tz��l�-]�Z^�%��;(1$��ݥ�17q0���5��^Tйov
)m��b����FzY�W5�A-"�uۀ�S��WZʱ6$��29M�� 6,�(�m	��sӖ�n�;�����v�!#g[�XJ�nm��lj��l��ı]�fV#�R��UU�V���);f��fVjʄ�����)
���Qe�����W#aR�j��m61�oHǈǖ���6:VkS�&c�lT���̚M�M�a&�\ul��Ф�w��V
/]��$ͫ������.���E�V�Ы�{.���B�� ���3J��
$�-I�����yݜ1Bj��/RjXss���^�y�1nn�L�R�W���Vҭ�=�Cz�&�k4n����Tzwf��8d��m�W��/��=;#�L'��$Q1�OM�����K*$l��0�ᕕ7Y�Z�k^N��a�޼�������*��V�Jf� ��j���^��u�X���J\�.�a$5�ӧjH�H�'��.�SdI¥n>�d:�]�U�N�p��ѱs���7;��+��T����u��� ���)�eֻ֠Y�6fd�N�jd�w0�pw��5���k+K�w�lG���<M`W��61U`yW̄�x� ���F���M�X��TR�uh;Çd�/��c�� �Ln�m<n�c;uyv��s�+����R�շ5�Z�ӷ5� �Im	`��-S�#"}q]������A�������SC ��t�8��x�p�{�㷹��GV��V�U)*Ȥ��n�,K}pHS��u���-6��4& hm��0��M�W�RI�+4㹮���nκT��(�ĹKS�l1n���7�H���X*�`��P�q]�8��f����QZ	e��S���6�
p�jޢ恷�Ktj&%�eV�p�H����������ea)�1Q�M�dV=B�ۨ�r�ˑ2m�݇R���JLU{4���MNĻ�(%��!��qԬ�U����H�{w-
��e�$1扛{r+l5�C�yV�VV2�ݶ�L����2}r�Tc>Y�[J55��"���z^�Z�!ݒ[��: (uթ�m��Z{�
�SZ.=ں�X��h�J�� efT��6���چ�	���Z�R���
��t��1;[#X	�D��[�n��66�b��-E��n�]PU�
�9St]ӷd���c$�1T��.�SIĂlX3i�\���LSkf�xƛ�C!�w���.A2�5j䆅UnԚ���D�3mԪ��<��ɗ�S̆GAU��Yx�z�#60%��M�g�n��s�`ZJ�L9�S-�fYL.Ĭэ��W�%��E�*�V�,c��
�wv�SG|Y��@�A�2�B�h[v�woR�u�1�)����ʨk,H��,^�-٫OF�E�/0aXlVe'x��n�ţJ^cך&
�s^}�0Al����#D6v�"�3x�I6��� �#5ܨ�&_ĝC#�WC�ST��!F��*�	��.U�2�kVZ�ʛo2�'{-�ƨ�,9j恕kc���ڹ6��*��f��OL݋0R�ȭ�[� ����SBmL�+&]�R�!�5xr,�I2�P�q� ޓl��F�Q���Ŵ���8-��5�(��*�YBڽ,n@����C̱��V̢�8C�.�y�����\�3�$[�xާ5�)��r�tk�Rܵ�Ë,ދ�E���UG��%<Q|�dђ7oN\�����k�|a_Re�[�"^U=KX��*���E�q�����-e�ѫ2��&�ɘ�Y׎b[v5oU����J�Z�ɆWt�Z���U
Pa5�z�f6nT
R���x� �I��8�d��Г�T)�:m�S�KVK��u0F�:���1n^!�RqëJ*-m60�xa��S��7�*Z�v¤^U�r��zw]hp�r�;�+1@�5��H�4�h�h�VX�Ҟ�!���V%�ܪ�Ӻ`�[��:�fK{��[�j�skv2�7�v���X�a���Q�ɑ�p�i��5� Д�����x�y��{�H��t�.�������'h�l�J����e�.����:�uQgx��U�����)/��i�˩����l�{S�>4*�Gm���.A�ҷVЬ���1�K�F��i+˷�y-�G�V֤!����v������$�K�Q�V�M�O`�p��/UC��U�zM4rbE���lmZcݙ	`P��!(��d��v��A���CD��Jq rW�E��۬hHs^c��\��hs���-!���b�K��Q�o2䛶FQ�m��]ʛ�*f!#j�r����7�<i;�%:ŔPٔsk�9�ɗ��ݢ���n�9��"a{��Y4�(��D��%H٧�sV��{u��Vr��C��lV3}�J���㨞(+��ޛ�9`�ԁ�T��yt�����-m-ؒN���4��K5@[YIyl#kM�=���G���=@�7��60f%J��"�5o��i�n��t6�!t,T�^'O���#�2�"а�ڮbs���v+b~S�;]J��L�Y�*ex�a��q�
��N5��d"����f��%ɽ��i�\�r�]4�-W�%�l�U��Q)��^.z0�՞&��/��۩�����qDp;���W���KVR ��*��Ȟ��kZ�e��|����>$a�K���1VUޙd���xrw�3�=d2��zo(�u+W�Y��u-t
� ��%�1$�)�Z �XiZmZ[}UR��Q����GL�Q(�Cin"W��Ӟ*O��[��e��$�I'ě(�x�c2���������ȉ�)'aǧŜ�S}yt�P0���Nf��gI��,���<Y��-(�"#�R���JeY4,�̲t��e�l�,���H�t��!l�95��'������U*�E+!ꚮҭ:�z7]ob�`�+��\F���ڲ]˭_+�x�Ȍô�Lf�c5�3x5p;�v�D�3	�x�6m-�c9�����T���i�sN�6s�a^��i��Z��cG��t�2k(�3���4
�fL�oE+��BY�'A��s�r�M�|sM�|F���Ҕ[�p�vq|r�ݦ��Vr���MA���h'T�:NȻ;��k�Q �w�;BiZC6*���t�=��}D�4�繍n���I>�vv�E��qa��vΣ~>E�-T��iO%�)V/mjj��:N���(�M�I<C2��0ݔNav�#l�n��'�FiT2Γ������Z�Wr\Q.[�R��y˔�&��+,�(���4��2Y�W���i�V�m�d��$�fɶ^���,.�Ei�+
�M�'�{t.���V��v�˩w'K�(�HI�!Y�����?�H�{�~��[�� ���?��xM0��?*'���o�W�ג�.sAf����:��Sצzg�;�NyS��D�Aur"벟5�SO�u�4D���-�7*��G4�7��/`R��V�妫Sh���؆�����5���6�5���&[čK�2��ѹ*�Y�T��g�KܓH�;�7l5��ݺ���X�����I���v���U��h9�G^���*oNv������r+�u|��ũ���x�e�D%R�}�j�V"xR7�@�t��dc9��!�7w7H�2C�M_c=@����?=�f�ՅCʛoo���)Ni��-�Q��a�浚宝1͝��`��R�Xa�P�%Kj�������\[��3g)19����kZ�ŽΧ�Ҡ��:['={���9��ڪmm��C��K�zmtj�}��sV�=�DR��j�;�)[ۘ��V��͍�5:y�$��֯�e�|Z�ҝ�!�汻Q-�*؊�m�[�ogI�u������lR=I`�U���z�(x�[��I����=�f^\�C��$i{WΣFfU�I�M�e5��xo��X+
C˦����v�jjx�u+�B��oyBU�P�n��ly)%Iˮq��gp����*�s�lC�� ���������\L���pjšY�g�\A�۪j��BfW�:��<�;g�&{h�j5��a�Z��r�q�|�k�J�δ�5������u��Ы72j�W|���o�&�n�m7��F�;�w{[��G�%�K�,
�ܩ���k�%�ȴo�c��m�eN���}})�C��ؽ�w�[W��0EB��m�r��c�r�guv��)U����%g�;m���89r�M����Y0wfj񙪗;����'�]&�}���E�9���U���F���B���4oq���:��"���\�;����s<�u����\����ޙCl,�6=�Y��j1��G��P[�u�ľ�X�e���
���ĳ@���7�ȷ��k�fq��(�ڐ�;*�lf�2&�$�����1�G�*���[Ww�qa,�R��2(ov�}�i�n=0V��m�:�t�a�=q�X���gw5Q�!V2=�k�FTŸ�a��%9��U2y��ugTJ�������6�M������1�"�^��ʋ��hKQΚ]6�حn�o����$�n���$������L����h�Fa��o�/�z��wS���0�����t��n
U݉�-󂤡PۦTGwn�&󣗘3�~�P���)�BC�pr�z�ZR[HHL�����X��M�nܣP�f��9@��i4Ml��6���;��|��}9�j��[5G����@:��;�O	"�����]��,v�J�ޭ��r�����.��{��b�Sfrˈ�ZX��T���ye���KחW7TJ0�hv��2G���_Q��nh����)Doh��&�|�j_5�{q��)�9$�:����{�s4n9F������paER�s�b"��X]F�����إ1EQ��B�vQ�[:H3���D3A�{*qy��ɽ�]L;7�Ҷ������`ۧP�M�Q�5��P�_=c��0���S��x�R�����k|�����D��n2��#�l*^{4�	\.3Պ"G��䴩�}U��ۯ"��8
�����y�YM��k���]�1]�:{�
�Ҧ_e:�c7l�[;���ں�}ַ�Ҏ�+/�^�Q�u�;�OF���%p�.@�Ӕ�f�/�<�(�t�6����&��ưcV�!;��&pJL[�.�1N&���]����j���KǊ��#��O[�]��+D��'ҷZS��=ם\&��	pg �_$�ovB�Eo�I-�Z�s��i�e]�w+�:�g9�B"3�����8v�ef�G�����皻o^S���<���6�Ͷ�ȉ����*1���?og����s�c�|-�h��v�޸�˴g���p��%g�weMə��qm�_`��i���_A��-�X�Q�Z�td;��=̖�f�=�9�r�t#ÞMG,XH�3jY˾�uӕ����{#�������(���uDJ��hBUԙ��C�'(�z�v���гN+���Tl;1wg>Doe���utz����Q���!�}�}��,�����7�uU+ڻ%<���҇9�ch�]3�dU+T�ޕ�Y��f�2�c��<�I��T�8Ny��i�� �>�eG���l��!���m�B���+Fɭ����C���.����tv�(GI�M��ϺB��n�K�IC����%G5 �,jb���B'.�|�˹8VÃTo��ɯ�X�f�%����,+t/:��d$��.�v1,h9Y�\5�dz_c0N�r�ޤ��:���|��s&�뇟_���\��$۳�U�K� ��WW�S���:F>�A国y�[��X�tM�Y��>����t�e�R�E4S;�n�@t`���kL���s��^m��1wʌ��1J/���ha[c�^Woo1���5f=�mt�/��S�is��M6����8v�X��\���qP��ə�+fcnX��O��JB��h�z�k��eN��Z4�[�v�׼�k����]�
pL�]�)yc�U���kqM/�!����\�L�ՑI��z�×5���67{���hl�睊��&���>�̨�S}+�U��Cx�%칌��`�6u.rf����T�2]ۓ6�6�(�n,��w�-�TSgb5�֢�t�T*��AZ�7�2�ü�
r"��q>ʇm�c(��a�Sn�r�69�(Q5-\K���t�<��Z4e0{{�f^q��,���'[(F����PRDF������U��/,n��Ά:7�'X����f\rol�����N�V���H�W�{Ӛ���kWM4��tr���,�ib�4B��/�aއ��M�n�O��T�	,����O�.�|;U8VYV���5c��YQV��kC�i��s�W��ԃس�ꉂ)K�T�^��4hۓ#�on����B��q��\�;��j���3�#��2��2������ƍ6��}]��U�} #��r�'��_g�b��
x�d��#Q�A�{I��݌��y��Y���V�J
tƀmn"�����-���ΗUk�5/wP�e>�֗�[	�i�.ݹ&H�Z�R�)��������M�v��.�P����dwcV�a5��n�R62����!����-qh�z��ʼww&Pa_T<�4k��[O��1ȸ��Sn�U������<L�ѽ�ՂlxV�Z�6j�k=}+F䳎��U�`�V��|'_7���l�r���i����a6�G���8gmu��J�uB
��L`M_�ݪvy}�Q��u���ƶ��z�1oA�:۾m8$X�0$Y��K^�3+��3�Λ�X8+3�O�V<�u;/T�w�'�-]丩vC�e.��L�1��	+6�'vc�H�X�(��n5�yͫ��v�5W��Ոܗ!��Nd���{�oL�t-N޽�T�+�=�j�4YCT�s����tv��q�|Ӎ9b�gufb�-�g7�8�V�6woOښ� "��_h�ciRg[�m�3����B].�wCu���GS�ܢw�i��,����.�n���r��
�c;y]G�p�#w�]8�	�g��\�򺶒JX��lV��ԓ���\5�_�:�j�-��b9'b��y�Q5��LR]�d%���wFaʎq�1"�����u�m���N3jm7�,����cj7�_Dv���-�|q���ms!�.sݔ)u:zzbQ�ʮ��v�!���<<��ػ09{Zi�X#�p=�K�b�j��h��d�뙩ս��c`���j��/-j���LQ�����u�l�(k�f��r�7ˌw�5�G�őEM
-�[� �L��3�7�7�ͅ��Ϯl˰�{������uZ+}8�qUv��]ck=5n�|���w)���Y�Ǡ��<b�N�5v��̵.Nk��]�a���&��}0.�/$���x���1���޹�̋e*�������Z�I��wL�JKv(�Vއ����J���윟כ/z
�d��%]t��7�:�1��^(�'����hF�pmN�;3[�ō��^�>��3|�S�86�SOd��]v��M'�3,�������u`�wY5���bzR	�u�n+��X���Zؐ�G0�R�+f��T%��W#QE��!�p�o]KӬ�9v��_Y�����ZcϽuf�6ݬu�e���JώE�����I��I�n�Q�e�)�EY,���2��(xS�]��)�%h��˨�VT�I�s���b�Y�7�Wa�����ԧp��b�M����I�.m�%��w:��"}�\T)-0��>KF��i	Zlm���܍��%�o閊7��m����ٺ����L����t5��E��1���3���{Ro>�)ł�q��á�R�-�l����8�􊐴��:�K�x��?�oq���b���k�s3h�m�|0�F
V�u���m��6oD���]�-CK���PJJH���Ys8��)`Яд߇c^��SLZ��9�%�]f
s.a�¬��	�	4h�i���Z���!�E#�˧��ύ��ܻX��p�̢ōn]�r�Ŝ4�V�m�ʾ�O��}�)�ro<�/�s�7s��B�ɶ[H�w�z��9/J<���GN�����$b��	�"��a�cg��a-���H��ǐ�(^��ު=��k��燞.�F��.zF1NwS���n�չ7)�׮��wA���u`�)p���W�P�Z��V�*�؝ �д�@L��2!Ѧ�G|�X��`��(4�7���·��k[׈CN�!�g��ea!��
�ɦ�E,j�ڈ�]��dv)ʁɢ;��3�R�@�sy�7�;�9�;��qFH9�h'�V��>��R���s'ܙ{-���{�i��)�Lc����v��֌�L��:� \A��n��{F`Z+p�j7n�eUpg	��f�<��������� ��S��k�ǊaǮ�V����g���ǈ7wՑ�;��C���ѭB�oZ�@��'h=ssǴq�'��;{l��k�2�UZqlޫ�7|����-�0Q�:���,�Z�z��\jI����8桃�WI�WÕt�n�n�hk�����$"`)�6˻CqU�r���et�n�6�WF
v[I�<���nA���)�Zt�k|gfl�$T����4p��!J�. �Q�
x��jk�(�UV;L!��Wt�wj�V��&`�\Uz�'�����S���ӗY�Ă�v#����y��sx�w�Ѫ՗5`��f�}5�iiS�M1�])�0*wMc�3���u�$�]+(�$k!�'l[w$g]�M��3a<��a�t(�ۜ��4=堄����
�&̛jkn��[���q��w#[�Jy]:Kv��k�Vn�.��VY�������V��������2��k�8:�V�7��#lP����Hq�KW:Ũv��Xĭq�U&�!���ΫO3ǆ-ˮ	U�y��k.ba�slEz��n���a���EB����d�qܠx����
}@	�1K�v��Z��]9l���/a���kF�=�a=��7Fv�.�2	�hv�kH+wC�|�=�#����g>
�>��!+��:����v���[���&R��E!����@�D7Ee-�R��ګ�"���Z; ���uU��9{�_Yƫ�P��W����i��{�\�$��YR����:h��I+�\k�W>e��wH�D�GV��	+s��WOb���7�m^��ײ*����}@�����"��!S����'�U�uܗx�U�[îԷr$��r]9�{�6)f�A}z{o�-��x�"�mt
�}��L\A�Ս\ͼ�}��E=7���{��Z�6s��)�1]�=��}�]�/��g�t�ww�:��2�Fg�|��8q\�����k�쏎��ə��]�\����Y�3�wL)�R��v���:�\��.�y�������ӻ[���+��[��r�xz��\�t�����s��@26d|����I���w���5z�=��<��'�[7z�^S�����^��j�5��8h�y�iBN����C�޻��O �A�)��@�!���A�}h��$��*�y/U�3Bȭ�q{#��!:��ܰN����	�Ȇ�2/[�5P��k�u5�u'Q�(��tY��p�z��.�Ԁ!ޥWP��ղ"h��@5��dފ����ב�IE��u��B�f�q]�5��Wv�ܹA�(����Q�+�{ԩ':�C�&D�*u!��r����?����`� ��ې��;���?x�(�"?�����?��?2~�?O�_���Ͽ����-%���fm�~u}z-�ݴ@4�m/N�0��p������V���Q�U��aXm�����;Sri�����NYp��#��&��L�Ōb�Mn��\��Lqy�b��#�&���=���9Z���)�ϞNr���i�y�jgN�hsM\��L�׹�B��uԦ�x���k7L��Z1=A��j�Ѣ$�{��;�����YWl�w�6�t\�:�[�}"n��=�Q���;��}���a�͖kq�-ٙr��Ci��]�)��B��.S���k$�4 ���Һ%E�|4��֕v?��vn̛ٚ:��}�/���������&��֥��H�M�g�MIN�h����<"ywٝ�lo5�s"�V�de��o%�;n,�fі���>ic��Ǉ��b�E$�Z����˺0�!_o%�r�)'�Յ�w�ءm�*�/qx	x��fFx���w��x�."��6ؤ���[6j�pK���y]��>C4Ŧ���:�����6�#�����ss.���<i��[�ڼMVH4�(�4���K.�_M�ya�����I ⧇ǟ��T�V�QY�\(;��fb�O�e�]�䰝4���2�^�=��JH���nѴ��8ӭ|zuQ�H�c����ܩʯ�N�>Qc�V,k��AC²>��*D�ō�-Ȑ�bD*[���±m������7v��qǧq�n8�8��8��q�{q�8�8�n8�q�zq�v�8��q��q�8�8�ێ8�q�8㏎8�8�8��c�8�8��c�8�8��q�q�pq�q�q�q�q��q�N8�8��8��qӎ8�=��q�q�{q�8��qǎ8�q�q�c�8�=8�;q�t�8�n8�q�q�c�8�8��:q��M{q�8�8�>8�\q�q�q��q�qǎ1�pq�|qƸ�8�n8�q�|��3Z�}�����&����V���k��(�͹P�8D#�%$��{3y�<4o+��lo�3Zw��a
Χ�vkKwn�}�r�>�W�e�9�\o0��n��:��ލ����D|���wt��P�C��q8�+���F��5�ӯL3b�}�P��^nT;!�ݡ�c�pm�����+b�\Uqȩ�Sڼ.��˗31Oz�9��:�Z�m���æ�&��ԯ�ܸtl<ڍث{�*6D�N鑊�1_fA{��*��z�-��t�X�
�}G.��#$=N@w�JגZ��<�u��}��[�v�MJ��Q�P"�
�[��]��i�vh�xs"�ײU���}����;KV7�'%�E�A��~7�4u�E��ƖN�F���o$�[�����4�@�C���fSҳ�fR���Y�ʈ��m,���GN][��$r��p� �w�S�8á3m+��M49�]�`u�,���]A�k(�17L�k�Q���)�i��������%���ō��`j�uՆ��JJ���;�C�X�5�Y�� f^1r��`�bfe^_��(b��Z�q�f���뺾Mn#���T�	s�h��@Z�����Wtk����B�*N �Z%�yծ��!	ʼ�dh9�cc�H�Uf.�.��śR�h7Z��t��q��q�q�q�q�q��8�8�ێ8�q�qǎ8�q�qǎ8�8�<q�8�8㏎8�q�q��k�8�8��:q�q��q�N8�8��8��q��q���qǧq��q�8�8�q�q�q��q�qǎ1�q�q���8�=�㎜q�v�8�ӎ8�q�q���q�qǎ1�q��q�n8�\q�q��q�N�:q�qƸ�8㏎8㎜q�q��qӎ8�=��q�q�q�8�8�q�8�<���y9�}�/�Ư�_�!j#��,�4��E�yʊr��i�O�d�:�U��C �J�����Xe�ӯ����p��Z�7����6��:��p�5h�υU\�Z�%��(�N[gK#*���u����V���d�ٗ�q}+^��0���b�=}Q������ؗ��ys���ս���*ޱYg]f�P0��-�_P{r!w�%�5��տj�`c<���܎9W�y�p�!��:���a�YΖ!Z�#f9�g�5���*h���;��2#٧��m��8n�a?r�[V�q���LA�� ]_<ˡe:&�e�w����ǀ]6������9��CSU�����b�۠�`��gWȌ�9h,=��	�s�ꮦ�>�<2�Gs��m܉v՗BgS Kz�����*���v�S���f�:��jN\�����.�hR9ű��v�e�R�oMlkQ�}�A�����|�WVa��]��b�S{�>�ֶ6$��/l�����^2��ńk�R�u]W!�j�l�I�˳P���!F�`W�LY�����oH(-I����c���٤�\,̩�i��%]������S�Bj������c}x3������N3x��˘�,;�*�t��`p/�#W��p�B����g9%�4b(oH�ޫ�D�<�y-�ksy
+s��܋��!�7���Qc��Sژ�]Uo�_5R�{״�S;��<��=��-gH�s8���v5�*�B�l
�ْӼ�N��0\�HΥ�ɻ�q�2�yH�3�����ڮ{��
��:q��+9�V4#�,��Zz{��%Ct�Łϸ3w���N�t�${U���2i�v�g�7��+XX�wO�.�U���	�.h�k�:��0����J�(7�+n�z���6��٧�"G�Ċʽ�0��J<B{M��/-x+/6��c�x��3��T�8宺N)5�*ӄ���B'����! ���Vk	�͐N��M��V��u>C���_`�&�f�4��E؞b��z6���ɻ��	�볍��p=�v�t馷��w��;�/�u�����wG���좺��71�{��TXc��0�b�·n����z��0���`sF��74m��J>xS�c7D����.�����d�c�Q�(����u=����˗e$
�o.�Í8+�c5gN�!��R�8��x�g)3t{�ۮj��e�ԭ	�Ë6���؅�^�ҥ��ndUV�icte��������M�^?���J���2��
VM�+;cz^
b��f^e9��؟mB+Vs��j��V2�V��x �{3uZ�-υ�ض��5���_S$�C�T��&��n���UH�ǹg/om3v:P���	g�ڛ56)��Ėi4S;	�OcɃ�w�r�Eܖ�X���+�Gcꛚ�\��S�u���1��LIb��n�D�Mo����ZE��>���r"�N���eǶ�2�W"���tҧR��!|�������u`;�<t�g�܆��sj8)�y�n�A858̺�(w�T�����`�P�W��8���wa�Տ��]��݅�g)����2=k�����j�݌@�;�^�-��R�Ws��'��8:�7�%T�*k��W�7�l���VC\Ԥ��	|j1d��Y&�j�P8��7��6U˽��nXb�(Z	�S)	��P�QU�SCR��O;����5���&%��^S�RiF	�n���q��N�]�HT�(0`x����'Ww8�(^�nG�}��zY7g��B�6�-�����L� ���z�l�0��wt��k3t��rVu�9�7׌
y�.��\u�i[�5�n{�G�P*���WT��L�g�:���.v����LKu%*�*��e+�ެaE���G�\��A_^��i�ܙ�!yn�4cl�
�QeuQkW�����6��.�/_�>F�ntbө/�7Z^�ɑ��;u�L���r�M4���/V�S5�!t5�)�~<�'n	Xrξ��*��*5��9��U˩˝��@�ڿ�]���k��k���X���P���{z� 8Q��!gk�V�n�Ι���������6�ȯ��\�9,)��.��/���+Q�U����r6�$�je�y�jR��*�m�E��i��į���b��%�d�H���Tt	,*}��OD4��_Wl�K'O�5��S[�䙡`�w��ɔR5�mVZ/{����P��Z�:��<��O�FU��K��I�[1���b:����w���Jܹzu5��fR�uirQ�(�~FK��d�ש�l(���;�b ���X�r_P�^��Y�]s4�eB��mq�fwC����RY��\a��W��c��S���K&�ݠ$�n���)m��u��v�|�\��`���(��a�Rm2K���(<���L�s
�-�.@DT�B��-~���]ܮR�ӎZ�y,�Μ�;�]U�OV�]w5۸��j(Ȣ9u��1�7�8�\|�� �����Me%�l��`}Wy{�2}�YWRJ	��v�몆��НVcz�r�}��dpM�����k�0��c�$X���T�t��k�댞[�z�S�1R�ǐ�jp��a��!�X1K]NՈ�7W;�8��O�*hwqy~*�"ʘm���/��B�v�iӑS.YI�{
7_�t�{�wl˶p���z6����o+7��.^��N���t���mZF"P�6F���M�9���P�A��5�R͙xQ���pՊ�I�sL��3sy�U"ͮ ��ݴ(�2�6��U���ۑ.�	�*P&�VE����C�	
�-ft
�d�� ����M��1R��KG���[|�ik��+�7����ݒ�;^���x.�����Ժj�Y �ӳ:C���՝N���^p���k������Wb�^
^0?]І�;��e�S�v_9EU���t��K��e�Z��x�������
�`q�6���#V3M;�)�
t�P�&f'SUR�nޥ����EU<q���N,m]����ˆ,*�r��l�}�|��0!V����CY��kk��;Y3(g��Ș�P=*#�A�QP��t��U	�3ӓh�}�v�[�#��P���0�Q�����mL��6�qR��<�i�S�2����B��v_ b.�\��Q%�nv5u�p�E'��:V�Y�o2�Cx���n�P(�v��g&��qL��+vq]2��K���Ծ���ˎ�\�f��p-s]�[Y�1ձ�ot�]LU�R��҇V���5�k�65ŕ˷�Z���V3A��\�Y�@�[u1%Qe��ܫ4���
�'F͵x� �>է�:7���Q`��M<J�	9K�e�iʌ�6��
B��Z�X�g$�A!�9�ٵk�-Ꚏ�.G��j��B�.�>�H�p;�5�����ڹ�(����k�'d���3����!�ǁ�4sUs�suEFҾ�cr���Z�zm!L�49xE됌��V&�}_<��M8%ņ��}3]��@N��Z"���N�<=6n;�����������]�u�I��]*����n�f�˛�hqt�"��9&�����3;�ʥ�̾��L�1�s��e�\U6�]���TbVoGiذ���{g��Uz��Y��`�.�O��2�ѷ{��e�����tvV�֟s#�/�pMy�&uU�]�gM�� f����lVin�]����4�V����y�QC�ڐe�kԔ9&a�Z���І]*��6��v��@�Vn ����*!�V<�哈:�VSс���2ȴ�
�"x��"��w-��*��fP��sSZ�O�^���X�!r��s;=��W�_6��Sm���*Ց't���F���.��̸��Cyn���@�z�u�]���č�m����J�`5�� ����c�� ���^sw�ĭ�����p��%�3�ykm��8ޮ�m=�	��Tޙ�vQ��hZ���]$�w!Uq�b`-���k�P�*�g�@��Zs��elA�m��LA�����`\������r��vY�|�9܀�'Q���JN�n�*�2�6Dԁ!!�c������7��f���
�X�]��,��Z>�EC��r]�Go��F��r����ٮ�����&�cNT-�{|sHUG��z1N�c�Y��CK��&�LC�Ng�}�Oe�.�u�+����b[Em��(Y�,'�f�:6U�����A��\�}6�>���8����JZUC����2�7�_5�.�x�N�E89��N�HFnl�}Jw1lR�d=awM#A�'T�4+�g�M)��z�������|�x�%,v,4�'uL�60H�-<���%O�ϭ�l�κ"��J�\C�['M�q��ӕ��w���eh�Ք���N���br�@м1w�Kw��.�b�Z'�}Q��U���VA��NX"H!�.7�eEQx{nUͱ��x�͸�Q����]�Y[��_������6��dkX�*,^��8˃z�YU����².X4�Z�)Y����qB�2��\�x!�@��ǵM��e.�[ܱF��_A�xډһơ������ ���W�]R�p�ˎ�i�Ms�OH��V�Z	$�{�`�;�;U�ON�y��A�U.���Jaz]Hm#S��wF���t�f�:��v��z}�'w�|�1�<�y���Gƶ��m�e�uM	�M��b���mDcm�l��E�U3v�*o���'h8��79����5��gT׊��a�ju������xB�Cg=�(p����{��ĺC����4���1ζ��ƶ�Zr\�ȍ켦.Ȋ�imQ���[j��@��WzH�v�ъ��+}]1�cyV׍���c�r�x�NRĕU٥#D�H����7��G����v��k��34M
:z��]�ld9�RO
�VX�cHyA�n<�Pa���A@�G��ә�D�\����t.���F�N�}Vr3��L��V`;����u(T�M���������_�]�7���(��j��}�A9�wf�ͫfu�4t�ۢ��9w�k{���?Ԩ *��C�?���w��g�����~�}��$���k��)AĤm4Bh����a���(X^l�À��TR-�EP�E�( ��L$��Eh�T.[`�H[�Xe�Ia��%棒@Ɇ(��I)���rX�)��!B�H(&E�P�lmRE��T�
�!Č.GP��R2'TPP��00i��9(�J��4��7��KlR,6��L�1h(ȩmnH�>>D8�&C�$$b1�Ox��_�o�-�~[����,�����2����P��Yx;��WLb?q�8��v��M��)��!c��w&���cl֎�Z=�n��(B)wm<V�w\Ᵹx����S���m�a��j�V��f��v�ŋ$62����dJ�f���5�p̈�*q+*��" ʨ\��DQ�ޢ�x'��r���j�Xy�x�m��c[ZY�������TnY�9e�Gq�.��lv�u���)��GK8k�k/�c50�s#;�q��Wd�3��\+zE��M9l�ض5�Y�K]&�S�}`7�FNn�Ʃ�k/M�4ۮ�SB��Z{�0�xM��[Ɠ�M�-mU����j/�W���8Byw,+t�r�4Y�/�T��"si؃�#7�Ɩ��Ap��^�.�����t9�`�N6������v,9�p��:�K�۝|�K��E_P����gw�����,�P�QcX��G1VǬ6o�O˫2�����L�(���n���t���極֓"B�1�w��+���W,�x�]�{V�\X�����Ÿ4㬗]���[�.��9؆���s��7�wG�83]Ֆ]�]n�����Z��m��RV��]��Y�]&8�O9퓻EF���N�J�ѩ�!P"0�C�,L^r$B@C���2a(B���O͢�~b6I���B�q��AL�	��S�$�0D�I8Y)��!�O�
�HRa�R��JE?5
,�C)��~�)TȪ�L �n��2#JӅ2�	�q_��6I��**G��F`.\r$��L�P��h'
I$�"�QH�#�Q%���~0'n2��4�$"@�5)�K�	&$�"a���#�C	!���i!*�%*!�D�L���%I� C)�I8�!	�ቲ!fQB��!@�,��	�
"k�@��@�j$@��˒�02���y9,�����(NP�(�2�ny�C�*Z�U�	b&QfH#��H�&ʥD��@�
,�$:2Q��"y���	=���8A����]��Bߓ3�F��I���L&�d�g�
�	�		q�����F�	�	`��o8f"D$�?^���٧kilm�����Vi�3Rv�vv�h�[�]񮝻z{|q�q�q�q��q�nݻv����H�`I俽[Z�m�vMd8����j�U�K%,��!5�:v���Ǐx��8�8�8�;v�۾�]��������d��6����{��Okq����y�W�"|��=�6�o�(_n�� {j-=u�gc�)/��)�0-�[헗����Oi�pm��n/l�H�d����n�{�����Z�g(T�ۅ��9){XV��z^�E���Nv5�W��%�2G=�L�8��2įo=��m�vn�fA݉��zNN�W�����,O���gW�qG��휖`q�T�[�����Y٤����-ȀO<�,��,����bu�yi|���d��fnVn�{�ֲ�sx�R���޺Y����w��s�-��#��������1ߞ��-�&�Go+=�U�vk���]�H�f��\s���=����ȷ漟*�)%��&,L��1E��,4�&�DR(���@��_�$U�� �E:����:3�����P�6���k����Jt�vlrL�}�uQ�����S�~���*;�Ee�
���4ɂ6qG ���H]����qB#(�0� �KQ��I �J$Bq�������P�ЁA!�#�
2D q�l4�Td�Vc��U�x�� �^��02.:�M�TZ�hz��&�՘)�f��Q��Ŋ�և�����p)gY47�ߘ"��>x����w+�=�t�����dǻj�^z��z�x���>��ap�w����JO�R��Y'@�����ݢp
�k�e읅�	����I�a>�1��g� ?uI�`
Ώk�{v	��'�.�'�no��}���'x w����ܞ8��Cٔ}�����7��O��`�V{|sz۸�$GPx޲,����ȣ��ڞ�� ��
�L䶃�,�o �`�.�}�sQ5%ף����t��������T׌������({E��z6���o��6
=�@�w5�=ǭ�_n�罦g���yk��}����Ol�m����߷������mOy���ɟ{�yuuטץ��u�m����m��o8� W�c���F@{ٛ$�vk�zG\?�>�"TC�Tg��Hd�X��T��&)tO%�ۗ��3�3n���3/�;C�Jǅ����f^s�),�e/\��Ya4����Ը�Ћ9�(���C�
ک槹s�ކ.�R�8Ѯ�꺛�ì��mv�����|����8DJ1�*�����rEӶ�h���8�x�����}����]�W���s�o�U����2֔g��tfO�
yCު��eחb��bpp�����ż�O�ޜ�4�h��w=�{ù��'��Aʨ�*4�P�����}� u�/OZޫMWw� ����vQ�h?�w���G�,K�U���>�q�{ˣ�հ����7q8��+y�0�5��,���r�tj{���ά�y�������~�P��M��S��;�.�y>���O��Sw��"_M��~O��̢{=�g2]���V=ۄ,�z	���?}��yU���������w��J�{�$^�?�P�v­�{�Ϗl�rf\�>S^i��ǥ��]����W�M]����]��1�t7��P�C��3���7yUTzzt��/=��v���4w��홾O�+]���0�M=�ڼ-�g�v�H&/.�h���;���W����7���u׻ǌ\[wd�S�f��g���=��>[qxq�����xǕW����#A���\��'�c����m�>���uƃy�+r�c�s)�`�P�[�W&���l=���x���:m^m[�`�7�c�N�E�>Ρ�����o[L��<I�g5̾_O���.�&��G��7xd=S�H/eW��wz����߽��B�WY�0�EEg�+�(�Gfz��ϩ���H=9��/}wX��E�Ͻ�j������#Q��׽T|b�恪*�C�*��;ܾ��׎I�[º�_�<Ě���K��wy�Β��5�¯,�8{���y�.S;�zc����>z�<�.��_(�{%����|Тh8,m�5n%�ۻݲ?u�B�w���ϝ��(z=tdy����8Wgc����^��.9��8CYX<\����>]��:r���0�@��?yE�7���&	}��3�r�o�\�t�l�!!B?fϬ��7��y��j'OdH�@�Pۇ�^�U,���S�<��u"r;�꒚��xV�����e���(a����\��s+ǰ<�g�[�A����C*$�7\p���Rv��=���x������_sf�:;�*�f�U��k�����&S	`�F�Y�q>�x��r}��>��ε�����[�=g��T:�xܴG�r#υs�z�"3=�$�����6|��W�^	�}����|�+������Ol��}-5ػg{��ԑ@ϥ@<3}7�_v�����Ѻ�4��m�wSr�=��3���"�90x8n9����^�b�;�f��뽐�dq���_{c�9�p�1_�mw�����O�׌�o�s����]��~�U���P�:���7�yWU+�}e빢��=5�ra�+�p9]�o���v9�^YӷW��{Ӿ���������U6j��#��,cn��$����6}G��G@�{���x�+7�Xco�X\���a��n5~�?v�*xg�޵����ϯ���LB�����NY9��"�4���[��DP-6f �מ��q�у�3������dZ�!�ҡK�W>��ɯz��Uo]�S��m7\݉{��kHK���k�B8�ӹη�%��DxJ�^���ί��a�ph�������//Z�eI�;b�S��ŭ<�;h]]�F(]Nq�B��U̙b��A�%�H�m����u��:J����x�;<kRU�f����OӯlU�fY�ˀVB�ٶ�l�~
�9���PC&����_��}�}]���ED���^_}��c���9��t^�b��,�u�����Fl�U�Ǿ3�9B�q{ϗ�;�E&A��������_����P~�N�A��y?fC%���g*����Vk�c��z��Go�{�K��ɻ㕎/y�i��hx}k� f<U4x��xU����i���d}��j���N�z֞{�|���Ϟ�E]�K��}�����(��o�!=�;���M�8z��Y��l�z$��V�.fr�鮃�	��hsǢ��s�vk�� �w���i�T�4�M�=s�~���>�SSL��|OF���+�_������7~��K/�m!�,�2P�~'�|���˶E5�u��^�ɪ ����5�'����ve?�ƾ	J��G����3�
����#9&�v�h�~e��P:���]ߺ��E�sr@��c��������E�xqw�Bb�@7�.a�H��c�P���0+��<��ðڂ��.���Բ��ɝ:��2k���dhq�}�Ų{�����̤�U�����ӽ���E������,�v�1�2���u�x�Og�}��K�����5ݕ�� w_�����sN�ϻI;I�n·޼���K�
~/�����sl	��1sgl��N����y��	:�uK�%ޙ�0G?���h���#���/�~̞&��{�L����l��Ǿ��o��.}D);�~UVC��}mv}K=e��^�e3�زs���Gg�_?T�^&�{~`f��}h%�9	-�l�� ����Ñ/u57<Na�ވ�R��KcW��nr}r�k	��A�Uf��h�Sj��hmr3��,�K�&{��k�gu}�é�t��Ë�v�����h=^���T�[B&���������d��nO;���}��ٛM.�}�o��n�W�g�L�g��{xZ~�x{��<o���c�.b�U]c�a+�҇�A��J����i�7��7��f�s�N�0��ھ��U��uv;v�"�j������	�����pmW	��6+���G�f�n��wnd����4�ll�VMzᩑ���~?0T���}��
 ����<7�(5���P=��q�u	_:����o+�wd�}�t�<z��&���x�/#���V�3�>�y��z��|�p�>��*񢭮����;z�ۑ���o�s�z�)��{�z3z���P���)��=Ѵ;�N����|�?L�/�~�����'���c��#�.�ws�{]{(Ha����vMhz��NKf��	�=W�U�|�v7�8�O��:����&8lS��������{��kN�׽��3;x��Ϸ�`�U#�UX��W���J�����W32��oOm�+�ڟ\�oYv�*}x��9a�󽓞��cD>��m�;�[,싎s
�7M�������3׍��5wQ��E�-�sǯ�=��+�{���5)��ꮧEϰ�����z$
���f^9��}U;L�}�9��,�GS56�Em���&*������\z̤�y���։��=n�Ge
?|	E�B��O^�.����;3��a�4�m�l���tLu�r���Y»39eH��v��m��]
���Y7n��}z������7�j�k�57���;�N��rz+��>��5<�3�Y�ɍ7��1���-~������S���[��@��x������}��|r�f��s�o2��[��1�JJ�/���	�4qj�{�%)�����{ҩ���߬kף=_*�3���N8�S��]���Y�}��-�ܻ>��}Y�Ԯߪ�k)�u=���}��9��d�俞+��밪GM�\2�t�����^��k�Y~ӳ>̷x��:��(��z.����/Q�} �ܤ��şfS^���o�r��۸�������7:�+�y~����y��9p�=��̺r������Y�����|�5�E�n�j��R��(܇'g�¸M�?I�s�}����Y�ע�qj�}ϥot��S�g�i{�>��Y�F���轝��ʿzoK
��9F�K�ښb�]��]��<�7�5\zK�r�Bz�����6\�,5����r%�K\�@�'[�BK�M����Nr���v��?s��RαN�����UΧ-j��r����1�UL7�7��
�{�v��	Mw����p;v�j�v�h�\u[n_=x'V�6@0��9�ۼU�0�xi׸�A��Oi���ӳ������qP�m�A�O��������l������NTa���4����ݤ����+�5� D��>V~�p|}K��|.=�͵�d��uO=oL�ޑ׎g������Njo��w��6{w��wo�F�3>��n�we]��._ժw���rܟ�G�5��3�[�wC2z���F�C/����I�6/N���e���0��-�NKI��N�=yn3Gҷ��^�X>��1�V=�1��[oM����ksGv�5L��
������\���O�������r��fO?�O�pM1�s�W{/�=����%��Ouw��l�ژ���jp͵W$�Hd�p��:���;�(�9;9�:p�����:������0��6������^��v������>��=ծ�b�@S��`v:�6��#iJ�!g��9̎�!���v��h��;{B�Tޚ������Qk�c�ux��89@���C�:��(+�񏻗	��U���Wc[�Խ`��\���k9�ߓ�8C8�q����;uH������_v�d��ϛ~�n��=!T���`��I~O��Do�l��������;�B��F���O�1*��@��g�������(��P���OfY�E�ݭ��iM�xMl�sw5vjC6����E�M5\筲� �vn�cf�� �8ϻ�n߽6zf���ηF!�»�R7�؇���]=�u��U=��2��2�9�m�g�����͡^�I�^\�wh�ͽ�:{fk�Z��#��N�i��ux�߇�b4��%��z�D��r�f�p"��䃦�9f����S�{�;��,I���TM�/�g�w�V?Ut>즀��Ѩv�o?@յ{ �߮�Os�������������=�O����(����U���<�c�l���z�{��I�]�ݽ��E'�7��̩�?#@�W`���?D_�����7���9)�_���ԅ�Ɯ��fe˶�/<|���C->��n ���r�]a�6+k���i���ۜ�p���֦ۮ@d �(�*�gLWB�m�Q4����Lz��v���B�&R�@�ַ�m�G�nF�T1}ב��Y��%�r�^c��U�D��ghק{4+t,ߦ�³`����!�ww��r�@f�m_Wn��Լ�.�9w�G�#S��vGs��v�/y�Q���� [-���mDq��(\$���l�S��,�b�N4OBU������j�e�K��-;��J��N���3�l��wr���t��qw�]�������f{7���OWH/^c�Ħ��8�;T�"T9�r��sj��Λ�Q��y�C�)�M��Y�ڥqZ��)��9�|T��rێ�稬/:ҮfvM4� /b)G����ל��9�\2�X�G���8��q��RGsn�Ӈ��L��#�z�֬�{ev;�	��e����mN��-�j<���CpC���]�/�9�6��NXcv��,\@u�jK�Uv�θ7���,e'GH�SeR��<[+��^L�n��y��YH�魚͸��^Լ���\ӆ=�|fo�W�,<�X/��5}z���|�<#���YW��'d����9*+�^1ղ����L��a�:H��gq���ӲH㸕vq�
�9�R�z��2�(���©���Mc�*�R�}�����;cO�]�EԂFIŗگ*�`�Cm�r��q=����hQ�a2�����x��[��^5*pYJ����:H�we����N1Sz�t�t�0Ih3c%��e�c�2�#�p��W�:[&Cǆ���w*��y�Kyp���ē��;]S�]�5�$�Ŝ]�b1����@�4�-�o��m����I�`ۺ�s�x�zf�y��L1n�x��t�~��3�4�T�X�3k�^�0�b���c�OzX��vE��L���T�eťGĳ�I�,';�Z�.L7���V�[�h��i���JY#k���.��(����5�(�ܸ�܀w4T�G3ĸ-s�"ަ����Ϝy������9�+�r�>�3}���cN�!�CI�&R���sA��nf{�ۗ[��["&1�ܛ�aN���}w�m��6�ۤ&iк��$6c�);�=�S��v����4�g��vK���75nv}&��i��]V��t�:��Nnm:���W���A:��dֽ�*ni���C���x�y����NX���8zq�T�2Z�b�'A|ܭ�|�o����R����oYn���Ӯ�h5]�v��>�๣q�lW,�')�1��z��ࣷJ�<ر�wazq��p�O�&�{C�KL�zm�k3�e�v;a*1м���Y� Jf����R��W��7/��}��7i2ݖ궄�������f��V���{=u�x;�p���W�֣���o���ȓ�t��n��m�ە;��=�W������b�������$���}kӷ���^8�q�q�88�:t����5��Vq����fq���*���79�[�E�<���[Uo-��Y�����.lf��mm�)[5u�k��;��޵5]iJM�j�$c�oOo>��}}c�8�8���qӧN�}x�8��Z�j��W�Y#�{{�?K����{q��׽v��2���?+��w纼��vf�[����ۣߞ����ۛ�g���y���P���#y�I�wve���ve�_{*Ov�g�O���{�n�>�w��m׼՛���������wz{��y�۬kG�Ӽ����,�3�֕3y{���@\GF��g���J;/�y��<H�8��ޯ���gu��s��#�(�:*A:�N��qoU��H2:�՛q�w_�{Zwv�8�˻.~n��/2���V����,��pA\D��쯶�a~/:�g�˛q�۲N��Y��{�@�h�$���7c�;�$��:Ύ	;;-;}�}�s�Xp$W~>uz����	>Y�G��;�͢{qvC�'��;0��@ڳ� �a$lw�#%�ۿuߦ�<5k͸{1���1�qj\9�6������v�(��wa5���+!�{��a�Mֹ���ַ�״�w׹�!ᙽw`*1	���24k�ll��rz>��z|�x����I��w|��
��|�6��bQgKsc�3�!��vx��BO�21X�v9��oqz5�4H��ASe�x���QN��d�@vf�y���y��{]��V��xy�-&~��q3��؋�`8���4]ô_�d����1Мh����6.��]��zoZ����5�P�F���~ZU�R�������b�G'.�v҆�ȸ����=W�,�ʵ��m��uTǔJ�� ,���$��au04�ˆr�gٕ�Sj9si�r�,�0�&�=4ɻ<�e��+(V(��W�:����ȯTGS�Ym�l�Fm���x�����|ʋ�{�7��2�����&��{=J6�*s��qx�˷���y�+<�OT�TI��7o�y����"m�hcO�)�tǅ�J�πj�NL�T/mM����$�=z*�e��6=<�yk�0=���G���Q�sc f�}!��)��k�F*`�'���xsA�Z�OAr���۴�0�z�mP�+hCO/�x�!�>`}ʽ�x�L�ewD`����{&p�z��玳�B�5���ُ�fm=W:%���WT}��e��ǽ
�k�%9�μ�J��eur20��e�RZj˹U��)V����p�B��#w�ٱѭ���k�H�n���%M���i���'������뽻�I��=-�\���k^ r�1�欍3�샨D���ǿh��9@/�#w�����g�.�u�!�n����Ϗ��G��L��d|�
�C �"f��=0��Z��!������Cϲ�5�����N0�h/G ����r��[xKh��Oè�*�[�VP�5S�)͊��Dj�{�S�g�l��{d9�U�<b��Qv�Qj��i�m���#��3R�=[�H�"}�ߨ\y7�����w7"�����y�ό�7��{;[�&�����#�2!��;�*�T_?_�W���H�=��z0Ŷk?����g�-�p$�8e~��G#%;v������|B�o�	��ߟ�Ǥk���W���}t_;��4�l�M��C��\,��fOŇ{$� G���]5�{�!o�x<�G??�lAPKո�ɗ�u�y�/���3A\ϺE.�h����t���@�tVzD�������x�szY���z}���C�a;��1)]�Di-{p!�]z�[	��=x[��^˦�	]
��[uC�Ϝ�f��?^/�V���aݶɚ?
��,W�Jj'��9ڹe�w-͖�\���qCכu�h��S�@�L�*�9S�(���TsF��f��������k�φ��#wU����59G��hC�Ly�6�|�H��^�}���~?{خ�fɞ�~f_,����p�쓏K���$�s3�ݲM����$J|py<l���y�HTD�c_>�osP��o�P�	Nc��w��EGakquE������|=1�G�5���@����zm�\��̤T�&�/g�P肟
�-E��v�����_>���Ą=6��Ђ��vT��w�q!{�v|'�߮i��7Ր~�0Oo͟io�H?r���ٚ�\Bc�z�c����۞�s�b�=��'�`~wΠ�.&�����Px2�L��k�dGNc��i����n�mh��x�a�W6�I���㚕>~��y����?40s�r��,6�jX`�M�ɷٻ� 3\{#�\
O#	�>��.	�<Ò2X���8u�m�\���-��]2��U�&un�qP�[�*b1��A���G�=hШ�j��� �D'Q���ğ�Xw��N�w4�ت��+L.b�0���z���%�ɖz]�2e�C�y���{�9�޿�+tK��ȰvF�B\ x��u��>���>v97N�	�>f�Մ���1��w��B���:o���_+&��	}��u�{J�^��1�{�������g�ZV��B��: l�N/~s�L���V~[���O�8R�u�T�7�m��r�-�#j��x�3�_e��v�u� ���t��s,G��x�ѹX�9}�1>�4d
T������x�l�U��yͯd�I�e�;���'s��G��:[�o(���bV����`�:xdﺳpwj�6vD�w��?��<�G^cI����G�|���cL�R	{���r�,^���3㚈�
��r�K�>�77o�u,��ފ�<���\@��4㕾�j�Dk"��
`�b����>w�̓Ӫ!�)��G+3;vsFq��mkoMMx�6��9���S���X�9�+"x3-|~��5A�u^�$\�oM��<���/�7z�gs���+$��wj�%�����)��o�9��-��t�p�g�`� ��
T��ͤ䉷=�(�ȶ�}f���:����Ιc��h�*J��VW�E��E�C4aی�s'Q,ޭ�L\zl�}���=��l�9��lY~���8�߇�\me�[�]��y��^jr�)G�h��g6��
�!P�S��+���d����wf2X �-��@�\�Smy,�aEFd��y :��p��R.��	��a�)��t�U��_Q��=,�B�ȝ[��z��It��Mܔ�oz������v*�4�e�����a>��{�䯿W�2<�G	6�@-�g���R��� 9�EA�O�iG7P*V�0*�nkwS�e��͛��>)?_cK��+���TTҞoM�5�J�N������f>v-[P�_���+�%?�)P�s_eEJ��X��6������	 ^^{7@T�dE1�w�6�
�'nqi���q%�[�������3P}��O!:��_Bup�Σ7C�f�wQ����s�D�f,Lq�����[�̾�lL�v�ĿNu�=��8���Sfwr���=}���Ra��G���F�o���Hv�g�_�mq��|�`ur+�z���왚���!��0��02���͞O<t���?��L�@|r(tǝ(�謖�<0���,�4�3B��=R�#���O?�y����n-r$����0֞	�~_}�"H�3���7��es��(�k���Z�������+R�kM�,(�����key�Z��3ꦗ,C5> ����^��Bȼ��&�۷����;����@R$��ۊ�ǅ,mWy{�Zuy�b^�O�G�l��2�VD5u���I��{��)ò�)��pR��f�7����)��Z��X����
�.���1v�eQr�\�M�k�o��T>GI(��3���g�v@�'��n��x��j�I���QrU�f�<·�D�9���_v�?�9�ѰR)�B�E�'�5���и�(϶�P�Ǹs=������[�g`�e��b�fס�H�}�}����ҞX)Y����%[�t|�_s��\%�ꉻz�-�{m�'�p�8�Vי���2k[f����7�r���VU	����wQ��Պ�kK'$-�ɪK0)WP�uى���/}:�9V������q��=�����txX�:�F�G=vU�`JQ���7�/��Mop[ko��ymgh��+����-����j"k�s��ͣ3�,o��o��<�|�fj���S��}|�}�*�����|Һ#I�	lҧ1�Ɔ�y���֨�躛Y�TQ��y}�/ǆ�>�	k�~���w!���~[��XΡz���?���y��BʘRh�d���ڭ���v��o�x�����d�n9f���1t�6��a��|�n��׹洞���U���v���`��1|�����(�x�T;����HD�F15�x(�[���\�����{7]T�a�;��#R"�y}�u4�.z��܉osB�g������qr�q>�^����9>kaE�bFz�(��'�]�Չ`-|��׾;��Q�Ի���zdmq��C���4\9ז,�)CT���Z���i3�'!��:���f˗O�i�r����W!�	�3�:j���cb�Ȏ�� �/�uj:_�ju�q�h.�T�k⌵�mC0`-��7@�D5JD��so�:1P�z�3�#�zU���&��2e�����=|�
,Ls�����S��k��E���W��L�= ���[c{!;�'�e5�"�m�}�І�o0̹[��<�s��ݔ�Ac"�]_!����0�գ�բ��b��yX��KU���� J��v�/^�hq����g��xs�����J�7ǚM:�B�8NU�W>G9�9E�i����|k���Vz�e�[�N+H֗N�B!�f�i.N&87E��F\�~�ˈ�fyXb=���)��[Bz�﨩�����9���#;9�0/O؏�R�&T�e�Nf�w�f`���~f؇� �S>g�3��^��r���v�� ���Q�1��|�5�unqf�q��ǭ�M��@�La�r��ʽ�D�V���T若9�X�0߲�3������#��v��Y���y�`Z�̸�}"�X3r�%�J��rCѯBe��W��U�)��rbg�^91I=�vvwRk�p��9���s�~�<y3(��>R��5?��Lu켧W�e�u�ֆ��u6��*N�����dOƏ��|oi�fx7��Wz�-��j%�oA�#LzK��Z�.6u��~�����u
�@_fP�o�iW�,>f�Ռ=��Z��A��)��]�ͪh�b��3PՕ�z˞t�d�E喾���#��R9Ck�F�����.�|�]2ש~��<��R5M;��u!�����u�����-��9mff�I�#�������>�cӸ짣;���Cʞ��qu�yO1d�B��ڝa�KT\��BȦƭ�gy�GQ��S����~c�f�;�n����N\�|"ѕ��]6x����B�ܹ�~����,?Bi���V�o�>���n�8H����ή(MZe�*$��M٠�S �Z�ɷ��YC�I)[�.��Q��#)r������������W���7�0�o�\&�wo��_�4��\Ȅ�i1��-),3s#����}�?��ٽ�}��8~�Nt�=��d���uoBf5=	yeQ���EO��&v2Zzd���8׉c��G��D����C������������~��<5{e0p���.i�H� cT����l�m��ŵ���M���V���&y�^�����$=�۞��<���=y�TG��j���pi�漝�n�������������^�~O}S�w��B���L����g�޺��.گ	J�ԏ�x{�
l�w皎���^Oֿ|��U���D�1M�i�6О�L;{Z9�2΍^��m��z�U;Ļ�O��?0B�������OO�C5�cZ��\��R��i,1�"r͝T5D�C�Ķw��3�P��b�1L"�8�'��2�}^��$�y��Bn��;�ҮOqC^s'�ͼ~���������Ω�W�
J�	Y�{�m	<���w��1{�P���CUd4�s/����Z��=5���:����+���mj����D�@H���,�w��!��0��G�*����S�s�o1|�wrAY�St��n��O:��@���7]�-��Vfqʖ��`<L(���#�~Zp�T�J��W۵o���M次��J�K�n��twuevհoBz�Q�7����z�o0������rv}��5۠��ӠQ}��Waʔ����p�ۤ����2���S"���۬,�`S�L����\Sנ@nFEc�Ws��Pϗ��oP�a-���5s�-�\��]0���1:�Ԣ��tGN6K׋��������;p�+���۪�C��ח�Ђ�ng��o����T��>���z)?1[��t�[�k�oJ��WH��z9óy{��Q=�&!-4%{�:�bg�+�	��$�Xv	TK�~lY��B�����#˫_z����k;4�FC�Lc ���v�>m�x��|Y�/C�޺����o���{�6�/�nj�m����6G��tT/0�Z������C�)o0��_���څ?Ͽ +�L__�ң�P/7S�#��>�ϫs��˘Y�<�yj�r��"������c��i0��}C���ݲ�A���+��<�1�YދOQ01��G'���`:�,a���5X�lrO�@e~F~�?6�����yI�x}եJ����}���C��Xp���xh�,�͈���1^�/��½��"s&*ui����zaݯYٱ ��W)�_�1ٰ�ʜg~�0'@��X�$O�zR���of*��FT�̴9��i�s�Xe��cr��;�w-J[2ΝsoD�]n��Z#09�Z��I8�����;��#�>D�YW��7���W��մ�F�Ql4��{[��Qn�|���kG�zf-x�'۽ܪ�+ ?���}t��ӧJ"��w����L�>\�P����Z�ZbL��J�&v~<>�x��ݤ@��ߠh�iC5��~W�J�w!�=��f��מ�W��Bp(r'~�15E�����})�����Sj�!�(c3���o;�=t��<����3�
�l�{VS���9���Ї���ʑT!�r)�c��TSɞFޘWd�ooN��o7^ځ�Hox�4��K&V�*�l��
��1,X4�pw�zEJ;�i��zr�33�j\1G` ��[�ml��}�	�{��i�z5��m����ـ��ifW�=������C˞��G�ڢ�ڄj�>�&��x&�p�
W9.[�{oh�z���)�WW�l�!�í��!�&/Q����}��V{�~���?-�|K���))����cN
�T�۰����hZ !���s��hsQ7#@�:vİ���xD�J�lMy�nn�C&�0�+g��J��]�}�WA��as�g�oz��l�	�.��9�>�Ɵ:�c�%�q�5���f�v/��0
�
d�TL�Gk��1�)�����;p���h����v��&�Pl�7����]Hټ��]��)
��A�z`�9�Vh���q(�u�q]���v���R,��k�n�v*�6�'NCWϦN� Yy�� Wܪ�ӭ�3���lիX�Q���Kc6���Gz�S���v�`K���oX�e1l^��[��Np��X�^�"Oh�pM�>��� �h��-�M5�D�l��	t�Ȕ7o,;JLG���S7y	)ۢ�46�z�p5$&:�z��+�msך�{m��ku�F�Ng,h�g�];5*ͦ�NK��c�cko��X��YA9{�U�S�gb�w1�����:��P}����շ��q�<�m�F������tf���fY�+c�u��i��ͦ-.�G��Ļ����D�_uъ��0��.��I��^�������9��������.�ݪ��c��ǻ��J�>{�_R��=惀���48��	�}�	�d4��ƫ'!K������4(6�]�"�S�qɾӔl0����ɳ7�G[�Ί��k��Oź�O^>{fN{M���M�<8�٪��c�5;jＯ]o)3y�t4R:ԝ@�G��9L�C���uʂ_T�K�4���Gu��#��D��e�ϱ������.�C�SG7G3�N��vz�w�V��ֺ������	�C��kՏ#���F�Z�b`��B} `��X�x9[�tvE���(^�5@ѱs+� �$�f���L?ȓ#`��/6�o^$�$����_�6��}�M�>�:n�/���G����;q�up��݋���΁ǀ�lͱZ�o+6Z��#�OrlB��Ғ�zya�A�0ܮ��-K�E�u���b���N;�
��Rax��:�H+
�ۇjҝ>�6�a����`��ɜ�U�����`�o���6���}�+�B�4T���j��;�s`�X���W,�#w��'2���F�;�J&��w۸�
�W��)'���N�h5�*�P�7W�c�I����ѤL#�E��iRU}܆����jP2�\;]�5���stt������|$��}z��̮��Z�e�/�q��w%]m�mp6�طs |�A��rG�;�333�c�\\q�Ё�X��V�3+cy�F�;s��Yjt;Ɣ���[�
��v�]��d,ev�{8�y��j���ӎ>&�
N��t������7ү���ɔ���l�&�wb�gv WA�\����sk��R��w��oE8F;*�u�S	q���g\����pG&�҃7vVzX�X�f���4ֺ��x����-R�}�>{�+�0�/�ըn�`�0���	��cq���v�	^ԛ��m�C:EFrZp9��G����c������8ٖ�P2��r��b�C��U;���O9�90RvM�m-�]7�-p{�28U���_{�I 	IRӷW�k��#�n�{GVS�gppqw��_Aŏ����x������־���������8�ӧN>�x�BI$9jXXQ�Wy~��/�%��#���*+���S��݌�BH��H����<x����5�������׏���:t�ӏ�$�s���kT�����Vڼ�N:r���;���η������Q�Irte�D�P���/l~�gI�gm�����*/�EGveו���\TR:Ĕ\����������!:98����"��8$�ˬ�:踋�9"�wdETGq\ApT���.󼐏;���יAIՙE�%qwGw)q�Gq�q��Vt����*2�.ku����wY�\\U�uOT�Ĝ�O`�w|��R*;��t�;��+�9��B��ZqDge�Yu�uE'qw|���J���>$@ ��]�- �M�Dh��n6�R�r��MȒ)�#!�Hm[��э5�8/2��߰�$w�)���B<�-Υ�d�)G+��R*Z��K���l�+��`��cP��S��˷�-n15���jM9>+�H��7B �!(Xp2$	AQIP�1aJh�T*e�DeB|"F�DI��(B҅��g�4�����5>§�l}t�WLt��9~���������=ӵA+A��{k��$���MeW�����L�χ�ZH$j��iż���{�I�����
��{5�p{ϋ�R��Ў 7��z�5/9_�t�wܷ/��f�a.;΃w���C	&-�����#u�qd�bs�Fѭ��͞�Oy��Ŏ'��C���:/���݀c��ѝ,���vX�n=��#�i}9^�i����L�myb�7��E>0+�%��=��>@~&yu�`�k�o]�e7�m�j|��� o�q0�r�o��mXCۃ��3��k^��X���5�``i�ri��hO\����O>��i��Q�S��M7�klC�1X���(z�(�v�o��`Pق̟�v��g���i�)�uC�ͪ&u��?�*��0Hf3k6�z�H�o[m���'�.���+�X��.�j���m��EC�3�}��ˆɊz���ٲ�y�z�+�T"6�z]K�=7�N���S�zSe��-�R0��x6x�9����y�~bH��i��ȫ7
ϐ�\�

y���Lu켧؁*:��C]<T�iuX��M\틷𥛵$^C�t5g�*�������h?�����|�~z�����E
�Ʌ��������ʬ��*"_Y����)��~�^�?k�g�,�E4��?h
��5� �2��]ʋ�ǇzOiJ�ܝWy���u�'��;����X+��t)Gi#�e�q�w��c������K^�/db�_l�ެ��uש�����������]1ӡ  ��g\�߿>g�������*G�7���ڻ���NK�c���[�q�y�?[�9�Zf�p~�=Գ��7;����3-�=-���/�8�xa�e����O޸7C��u9����M~?�D#�0Z5�c�}�Z��ڙ��}z���}�T Xwf�tZe۟�ɵ�(}�qxk���:����I-�U>yjݘ�����x��U�������弗�M��8c���U�,$d�X�7���m:�uR�Ѡ�z�ߵ�;���$���,%xLB	U��.��}�Ъ�%?�~�z@����	|h�~{���f�=�7���ȵ�h�f���Y�\;6��<C�{^Y7�FAo^"�b���J��3W_wQCױ~w��v�q�� %^�	w=�?6G�A�(i�~�C���M�\�BP�|�S阰��n��=�,���N���~|kT~����!fd�Ny@M}��^~Em5����9}�e���w5S5?0Z6Hg�Sv1�iP�K�\�f��*5K��Pߎ��R��a�1~K�o�	�X�#������׎u��,Lǅ�QLu��b)gp�~6ȼ���\��Y���"�@���혺��k"�䋃G
;���a�sڪ$�L�6PW���F�&���z��z#H��7�BJ�&P�2^��m���F��e`���iM�pjh�A�ɘ��ԇ;bW�5�][ʬ��ۖ(d��*��(�W�&w�μ���O�P>�1����z<=��<T�$��C�,"#�D�7�:�`슁�Q}���eH�������zZ��e�@,h�B��z����[m�ޛxw����~���pŘ*�(���6��>��Bh���v}���"���o���(��ô/ٝN�(цLmp�Z����A��`����u�v!�|g����^E<2�ԛ�I6�/��f��%#��M��ynY|�����ݓ�[[��qt�`�<��; �F��rʹL�N��Ӌ=����[4�����1�YY�Pj?>�d�����������1�s�G���Y�5A.?D�L-*���W�o!����&���zr���*���8�l��<�%�3�D�O�Ȏm��O�i��<��'�5<]��p1��������!{�Y�u�M.����wߠ�I�|�Q�i����~�Y��zE�y^%W'WL��	�4�'/I�z�!�;߫�R=x����.I�c�P����b6�z6w/�#n��t�n�ד�'��w_!���:GD�g	��0��5�[��>&<�7Ty�S�p��*c��+���tf��)���u��/O,X��h%t[���TG)'�YM�"/-[\"ҲX�L��`�l����9F�q��S�ł�K�rf��N��mLy�|GW���b6Ot�q�����9�gp��޳���8�J鞏@��=�}a	p�T������ ��OH��d�A�r�P�I����2�v�dDh}��']�1�zee��a4�Hxھ�_(��&��Wܘ�,�t�m��zw�ZZ��lrr�)Or�w/�6|���f��8��D��{�+ӣ���@��y�4�������6L�l��GE.K�K6̫��^CCx .!��C���ԇg[	�K�] P�f�̃�WC0T<kר+os�%.W�l{�u��=X�H�}�������Q-$��
�L� �?���}c'����}�y2� �W^���=�`Qp,1C��;5�Y�w�圉ߧ���j�أ��P��W[��恂�ǣ������1FG�6�$UC2z�'�M�9m;	;ވy�{/B;�~ǧ*F��kAF�^������[\ǇK�^z��Gr�k�A�u��M�[`[vyl��a�7���6z�A���\�f(��<�mh2��:q)�l𼁳�ؓ�;��s�(��u�M�
�Ǽ��ت�D��=8���fò���QMmB�6�O�1�'�~�K\�[���5!I�~�A�f�|n|�ս�����e>����]|7��uvwC�}YOEL�r�G�c�T�e\x���6+s�,��mTx:��YyZ8U�o\��w�i]�7��h'w�k=rj?n�G�Z@zK㧄�v��ǽ��w�y������}(�����HWL_���=�Y{-���U��{���nf��<��rM6��C�s��7��q�C�j�X����%Yҷ	|�_��*&F��n��jӒc�F{aT�\�O�m�s3z���vV%R�{;s�r-)�4v��y�t\/?E';����1k�:}g�<��������~��x8�TSp_�d��w�<���;��ۻ*U�^��s��$b�ӭ��l;w��-�=ǆ�x\�Bn���j����o^hC��Ƒ�3�N!�����˙N�FK%���y���-��;��>ew�%�0uB��[�򇤷�<�.���%��<����a{�:О�͟Y7�����Ú��Ʒ�Mgwk�l�7G��?%ʾo	~?7�ɟ0��Ĵ5���F/�ϝ=�	�wO'��
i { �z�MU��v㳥o}�,o|=|��ʋ���KHp6�S�0[�x\y�)�xKW-��Ă]�\�.1h�N�z)��<�t��9D�O~�ϗ9zZ+�=O��X����,�\3Zr����]L��\xޡ瞬�ϙ���j��Mr-�9�ǣ��hd�o��z�ܢ[�CM����<6O�G���ȵT�7���;�WE4<�k�犩v�,1?3#xF3H*�7�u���u�4�{��P���3�����aJ�!��b�����I�k��ya�鉽����`��Z���5�o��	a#Q_3~�) _�sڱ��zz�On��
!o�bV�?;����>��q�8<ђVA���R�K^�Lٖ���t�=��~1Ӥ@���Ѐ�����k����i���O�ڮ�����9c#� ʸȖ�����<��7v�eYNθ�U��ͨz;}�]����T"-�����"��T.�5|���z0���Zջy�ۻ̈́{�*�%��c �LC��e�ʱ��K�r��g���Z|���:�B}��J�Y�>�3����}�=�V������ŵ&��Sŷ��\�H�%�%9f�Jq�J��jE]���{{{��V�!xq�%�(;��ׯZ̡C�NKվ;�SH���Z7��2�#&%��_Od+��L��u�C��!&<�Tv�ٞO`��\��JG�GZe��&]��7�D�(lx�I|���Z�n��v�l`5���e�O��@�d<�SxO��Kq|jSu��n*8�Q��Xg��۫�/���ծ�x�)|�����m��m�8hș�<\Y6���`�-����ف�Y9x]ˎ��=>�ge�]���-�F Ҧ���'��ţB�S	b���l�z�˃U�]����ۙ�{��\V�k������v�8h<	�X3C�iz�O����̔�^���՘<4��E������K;޿C��Į�ڗ+ӎ�W�'�������);DY�{�f��`[3��m���|�c�_�E/7����-�ᥰ�6�D���l[�ʂQ'��6�/cCy�z����nf��M�&w��2S������c�B"����3�}��>[��y�vg�TdW��I4[�L[v�>x@~]�_��u�|'�
������N�|��on���v�r��>���4��|u��P�0�� Ny"�z����g0.a�s:������.��]0�a픋24��k�q��� �]�������oSs;d\%��PP�7�]G����<���!{ޝ��P��2OC��[�U��ǟAb���M�bK��xʤs5\�����`���큄C�>��`8c��&��E��t]�v��Ahi���Lz�;���m�4��{1�1�㋿@-/���p��z6v�8r�SO��OR㚤
�nJ=�4�t��ۓ7���!�7�E4WG�n\n�c�խ"s덨 )+1+6_�慠!�@|�;�6wi�d�ƈu�����M^�oJ��m�٦��mz�8��a��b�d�>�ݙuz+����魙�$����W��9�G��Dߧ$�|~+՛����t���Wl�ި��	O���Os�')=�W�F�Y޽�|�H{�|Ԯ<-D��o���<,�<�W���E�WR��<�n��o�WU���7ɝ�Bo �}�=�{c���<� �_4˫ξ茖��>n믾Dp�W��ۼ�i�%�1v�랹�����'�,f�T]j����ޣݽ���;��D)bR��1ˏ�ۼ�7�B�D��p�� ��7��]p˗�xk<�<�H��N�Z�?0���]/��O��剚�!�(�i���z^=>�jM��5�����J_���1I���[��n�ӆ6�6j��CٯMK��k��1��y������'֎vokeϢXׄJ�or0"�sjF�/Fr���-�=:�$�$��Z��矨?�h	��|����Oچ2�Լ"��-����ꛧ����w*�twg!�W���;�0��n[!w��^�Z�"�������<����y�����v�nJ��~d�ɤT��`cg���B�t"�����x��@��dgv���V8�~�L�p!���;�������k��|e�g��|�r�W��^�oT�8�i���" �'{�{a�{z� �/�GS|��~���a{kcjض�6#��@���䊅b6Ͻf�V���z�� b,40��fd�y��H� ,��%ƕ���^c:���\ԟ��xkQ�����K�1��ş���9�*���d��/�2~���^ONU��/��.��rW,�C��3+��>��9K0ƒ�=x=�O#��t	w��Z�o��[�׻��cYjz	n	t�wX$wg�so svѹA�i�R��W�!���a�7���3�ΐ��~&�5�w�f����?��q��^�}��1��9*`Xئ34�l� sּ��Y��(��W��T��V�jn��� =<}�ТWLt�����s��w�j�l��?��[�ݽ7�ݨ��T%�p���rLCE%v�mR�y�~��-��C�_W�ϱ;�Q@;' �ۊ��`���p����ƨ9�|Z��i�h���x��hEȦ��9�]G�x
ޯ!-B�G��l��Lߊ�C�<3f|�b
F�{7������u���\�>m���]�oH����n�cω�8�
��cv.��㣰�B�1��d��[ NL5�#���4�5�*|&����k	To8��*��u-gҡ8�j-�ln�z�9�:ۘ)�=��:��^0ְV������
�~�z/����9��	��f:��U*�}Yݙ;^�\��*,:2���#�%���"<c�>��)�0�):��!��ӽ:��xS 'j:��|�� KL��v�["}�Ry�7�Z���z~���f��`�*����\���wX�<(	�R銬�)��xW��GF��e�d�2Y&0<��Z�c�qY�Z���ݬ��Q�l2Pa".8�z^S�{� ��zg¯T�����{�Y5 sk�Of�r��k �/j��xO���@Do�ڙG�T�\b1^��Rz4τ�nAN|ېz�6Ll�nJkg�mm{ß��������5�:�^�{�U���H�o]S�)��cɃ;��}�:���k�ՠ�@6���⛓���Ѫ���o
b�ڒ�B^um����&��3�n8R��fPh��Sx���M�n^�}��ߛ�9��T����JǛ������{v��۲�;3P���T4��Y��"�
f��Q�?D��,-�á^��k��⑭j�ĩ��9��sO�`��1���`^E�g�5ٴ��8b���F�'�X�	���ѭS3NK�}��� ۉ0���_�����Z�������M	����<h���N�l��꫷z��p�	�����y�]ô
���栟���<Dc4�t�T:��b��X�˷�T�M^V�|zt��$B��R�n)�����6�0�(A� �7��[+Tۻ�v\�m}�e	vv���P�ǢX�%�0o�Mn��(EԥW�����k��':�}m��a���_�N��,������ӈ��k�#g�u4v���]�@��}T>��Y�v�%g;�ʶk�-�t�?	��k�͗��o�Ch��qv1Vܷ���4v�zq�=q�>���Bp ��]�#���Q�������7��ƨ���yoG�3��~݂{��Vq ���a�~vP�>WL��Y,�GS]�d �f �]_���Ss�JG�i r�؝5�Q`C��� ��]��>������n˷�cT �cհ�9MV�4`�Q�gl�زJ�$k9�s�|�7�
�J,3�������q����^�v�v5]���-���%�6���ڊ������݃���s�t��@�Ұ���]����O��J����˙*��1ȯYܐ��q�3������:�K��XE��wtMû���ѪS���Rw(D��]�9�;�^,/^=�T�94%�m��W��k�Po:�ٹ�c�]鹔ެ	+YyK��`�2��/�u��j���A�ܵHY&�cr��ruּns���9�Jr[s����N!h�+A�<��ݲ�1^�z�0gl��.�X��s)F-`P�pwp�F\	��ѫ+d�:��G�\�tNV�\|�|1.[�f<�Z�88.e�"�BV�w���;��fS����x�r>����:\��j����ܲ3S�覰�Tl�m�ݺ�C4�w,̫����ቱ�f�Ԕ��Ϋ�9ޘq�IV'RL���4��-�ż�I��쵦��9�z^\��X��ʌW�T�b8b��D1��u�.1�:��:�����C��D�J�UBn�=W�wY�ر�q�Z�UW'c��(��[B}d�vV�O��+�7Wv5*P�;������(0���T�l]\Y�ha���o����x卹l��/� ���;LW����Gx.��@�จX�*��9;�,HְH4�7dK����<�{:i�f��]�@pR/r{�B.�����l|�c��s�13I���J�͔��>لV�*h�Bs���%5MM<����6�Ļ��X�^%�q���0:����cg0��5s7+��o�N��L=�;�{����zn❔�ʚW��a���f4gPY�f��f�T��[��!��a1���b{���ξ&�(���jV��0*G���e���n�dr�2`�E8���/z��G*���\I��#�"{�X�$8������f���yRh��*lU�1z���쭊����J�&�'ZY�fAhf�\����A�Rh�7���J)�(`r�e�]8�v�P��d\��p���/Uq�ǝ��FHs(<؍������7T3�=�:���Y+t>��̘�Mȯfͥj]�(@r�G����vG.�t�rtk{xKqX�s��3Նw/�)��b��Wek]ǲE *�)E�+��.�ԫ5�o��4mY��	Qۢ���+2!�?��t'����fZ�?ظ�虳�H���78aǼ�,�UhA�2�n���uC;��:]�ʥ����:���k�3��]��Wk/uZ�黈+�P-z+9�E�L�ꋸ*o���S�t�s_^�"�5���`T*�7����������grW~���8��
.�Z,%�1�t����>���q�q��׏��}}}v�ӧ׏��d����9#��6��m\qߧvu�tqEyv\�Gq��Z�)'ק�oO>��8�:q�qǷc����N�:}z|<��!�W�����~�v�$�*��������^gAW̎��ʲ�3;��:����R��j���m��k��;��]���ud'Y�E�2�8�..��;���
=;*�[w����(�һ;��"����"�����:΃��2�-�n�,���ep6�.:�����^w�S�Yf���qq"tۻ�;�"yg�ŕ�P\D\u��iVu'EH� B]��vwI�T�Q�qu��u�vFV�죨����Q'K���*����!G_/���|�8�8�8��u�J�Wa�׿���aj��ب��;��ƈ<w$��7`i��fX��TsH��7�]k�X� �n�A�m@���,u��5�w�q�����>���+]1ӡ@ߟ9��� I�߄��0�k�M޸,��I����=��M�����SVvתE��.�9�˶he��z�M�w�'x�m��d�<�2$
�<�,,ҞaA.�n#U���>s���o�K�E�`���5b�w��8<=�m���=������N.!�ޞ(-�n���O���Q.�E�% �<�������Dy���<�!�Iz��O^U���V�
��'!e�unwn�l �/b�C-.�ǯ��oH���ŀ%�6�dj��hD&
iTl�>U�*5�#Щ�6�z���50�j��?!;�����Z��
��ãӨ_g�3kǎmO�9��#I���zi�{�}������B)j� �Y�/�D7c|7���~��~���w���R�0�_��}�u������P��b6D'�����z�?ai-{���~>�
�'nz�0Y���Vݷ�.+`��Eʹc�w��������rT
Qk"���w!�/=	��[l���i�d=*�̤��լW����$��64@�Ԝ8�g����cBˉ�x]~�ꪧF~�^\��+���z�eh���]1� mn�i�X Or<��s8f�lSo�Z�-w/oFn�0a6�t���+�.�wӥ2�_q�m8� �.����-�EL��;A��_�Ak��#��"~���Ge��}��?g�?*�Ӧ�VD﫽�ܖ�!����h�v��Ȝ}V�-Sm?~H�$ѣ˾���nH�?-�Ee�ns�2>L��jqK#豑�R�of��,]�[@D<հ��= �1+�GѾ g?��ݺ��|A�N�y�16�Q�
�<���p%TȽ�M�ԛ�6�
�ɏ
s�s[)�֍��Wv��O�p�^WB�g��c@ǐ�G�d�T�z�]0��Jn��Um��3�p�-���=k���9��*�����!��] 
�?[���v��篺#T�qA�������xU�(ގ@V�2�2�y7�k��p���h���x�Z9�_-�Ҟ�?��m��Quv0�����(wu$����]ndm�`��3S�{�$3�pa����6�Xu�.���¯Q5��P��a�	jI��m�d
)(��Q���02�0 l :�髯(Y���iq-�2�^|�+�Z���gހ%��Jm�25��^hj&)�K���H6ņ^9���=w�.I�a���)l&Wy@׈�1O�c�����-{���ծ̯�,��.��1o�ɯ�y�x?+7={���o�� ̐]Y���8@:K��{y��ݩ�FE׻%f�U.�G����
�=5Q�E�X������{E�YR�>Lj9�)m�1.��ͷ��oz6�$G)�|���_ї���xy�y�淛��sϲ��t��Ht龏x $ӱn������o'�:�{�&�D��3:wfܺ�Xh������\;�����}�������i��0o�+�L#R��P����sCT���=���j�pd���\˙�]��R7Q���y�{b��xf�c�
�0%F���k'�<�D���QѢ�Y]�����:�7� j	97�(t[�(94��J9
�T[���*{�߫*q�[��N�챩�b�z�40O�h/'A�Gf�������\�ڤ�:�5o�>�(݄����g���ɚ��3{I�^����}@c�_O��w�]6�^��ǡ�%��{R�mLXǬxO����q��4u��Ⱥ�l�xX0;���J����1i�ɲ�'(
n�b]b�i�42J�:x7wmR�'.cC�/p�bC��o���D*�އ��W���X��;��u��I�CS]����	pg׳��|��� [�c�Z�^����xtט@Ol�ߒ���D����v�N���γ��w�WOX���f���S��5��c:�q�{^}���׎��Hg�Tz��w�u�2�n:�Ω�Y�D�f�f�u���Gc���wCs�|ĕi�r���O��5�E��z1���  �~F�ܼ��;�Xhx�u�����]����0۬��:�&pᮃ�5oG{7��k:m�^��N�;#��\��Z��������K]��E�-�#�#ܰk�Б@�&�ڥ��n�x$ܖOV�6��3���o��3�?OO�:t�H��W�x���j�w���Y��i���i@�T�W9L�֌?g�[`v�*k�z�[<�6M��3nw0�v��1m�sߥ����8���,�Ѽ����eC&*̖K���B֛m�.-���7w�g7��0i��p�A�C�
9�0]�k��EV��o6vП�l�X i�G�(Q���g������l{����p�p�Å��{�S>=um߸�W��=�xK3˳�}���*��5���
�G'mq�ȃ��<��V�H��~��Z���w��s���ë���彴�
d��W��~/�|�� b�ƽ��bB`�a|�z*����h��~�p��{/7b�a�����i�f�(Z�F(���C�c��H\��m	뗢��W�Lb�tsф�&{�6�xV�SS�&&-�{��$�k}P�/DI/�?x��
�Y��.�PNC�[q��jm�fV�����Ѐja?c��ʥ��B�]��_�؋�O��B������os�ٮ˥���)C���p����#�b�U�� Xk� �U�?T6xR7_X"��dK9ߵΌ99;$�ֻ�����yw\_J���n�4i�9h�8m�Ρue*���s|�w]�}������
�i�,�n�Μ���Yn�\ob���7Qcr�UȔ�^q�ը8T�a�7Y����$Z�T®h�ޥ�['�!���]Ӧ�PBDDח�UoaUU�:6b&�-��k?ƚ��_`��C/덭�r&�Y]���O���>��ݑ�p&%��Q+�����_�s�yN��W^J��c�0��v=M�ڏ@��~.�h=��>�-w�q���ꕌܶy�0,oL���+=O�xb���������Љ���Uor�r�߿�;M�w7z.�[!��@!��f�Pe���蛦fj�\��O��+,m�3�1��%����E���̴̇xA��A�Z ��Ƙru�Mɐ�SxwL����t��خ9��Q�v�ګν��y;.'��0+y~�Q_�ŝ�C'����g���q�k�l������4f�����޷Mj��A̦ŷs�8�[6��i���" �������F��)�u����XȜ����"1t�|f׊����r�3k��������s��f5>�E�x��-yÖ3ykJ�{q��c��@��hkH� [��m2&#�1����$,�фt�����WDb���ƭzm��ɘl`98�����hׂ�8Șn��ރ.�RkƝ��xA�jBEb��.��"Oc��6"�ʩ�U�W���޽��'���?`q� ���#l!�r�䎌��г܏�]�������Oc��r���ϖ�8�t"^�(V�fm]�p�tr��t�f�&�N�G�_ʪ��}^5�t鮁FAFD7�}�ާt�[���|#c���vo�,=�ƅ�W���7��W�	}��~�k��T����ӗ�����ǿK�<��-���O��N_�4�İ���b��x{�
T�ƘUј���([<3<q�`��h/�k3�:,�b�C}��R���x�]��W%:��h���j�z����I�C|߶/;H&;�(��G<R���Â.9=K�sR�S7�_n���q���R�>i�9�x�L�+��V>��O�⹈~��xijgk�-�M:��q�{0�Egjԇ�<
��a�����[�j�OV�u�(��hO�]�ڈy�ڟ�~�J��V�]��.�����z�S�Z��9����e2�	U2^Q�f;��|���a�:[�!)�	i��g��s9��٭~�t.|X�?7kA~���i�Py��%�Y0��Sw6�癜x�Wu�;��5#����c!���\[Hjjyaʇ��	��5�@{�+�Y�wx�&���n�u�*�A�R�G6y(,WG��x�0�/�1[E��5��C��EUK�)g3ۛ���fn�g�q|%�N�����M�oMҳ�C3|U1k�[�����ׅ�����v*;J��,�M�w8m5;�VrҼeI��TV{��d�����dq�� �X#{ZXR;l��{'�����W1�$���w�.u�}���(}��鮁c�Mt��`���>��gk+����3�қ�*,�6��0�!�q��~����'�:�e��P�{�|ni����@3�pj^9����Ό-�����K.Q��������SjD���n�
W�)楰�ƅ�R3\3n���B���o�'y�S����ϕE>_�,�Y�����c�_�{'��7���>�6�7������J��;v�z��֕�m�˰��%���c�w<���I�ɟSI���� �kyO�[V�inwޭ��皪�+�<�4��&'D\D���B?VyO�a2��l����;ۈ<�Ȍ��1����l�:�"��w���b�ӟK��������C}���"���}�s^�U;���Z=�����o6XgѨEy�P��C7�`�� I�yg�	�{;�C���s�Z�=����J��4�v�^޲h
��U�Y�͍^+|�L'�w}2뜷4����V.�9��=qI�o���o>N/J荞���K���Ҕ�|��J%����rz����w��}��vg�ݷZ�|�Z�U���B`v���"|T,z��5z�K&��Y!�~s��~&����ꮧc�I�H�ӷxҜu���+�q���򗲲��u!U3�������d;�h�~l	�������E�,ub��ۇ��}�:��.j_%��6��2��� ��zV�}�s&oqV�����g�����z=C0��<U�整��ȿ�3�3���̜ ��	愡�O*�75��׻�����O�ȫh���;����u=!�E5�l%[�mel�^;���yƘ����%B�9�1���)%�규�J��7�����:�:�@n>�16*�_ă~�3ǎ��:*�~�
�3�~�/���)����`��	���3���)�)�j�������i�r�ͷG*Ot�h�\��)"�)%S3�:�)�2�2iY��"�S�r��0��Z�|����W]���&�#�L��Y�jwЏ���p��W��{�:��>���?k�]�dĘ,�r�E�n;5f�,������;C��TҀطp큤:�o��/)�{�os�^��
ތgJ=<���k��_e��>Κ`������[=����Q_|��g߻�ƫ�@�ີ2��ӟA��D쇥��֕C��b�����Ϟ�~D4�:y#��LV�m�j|����dP�ۻ�}��*�QfGvzO���L�if��	�}�vs�"]� ���Gѭ	�<r�)�\gٮ�
knfD˔sS[�@���WS*b9��7t�%�9Ew'��Q��9ۮ�%|8��ڹ7�z�nn���O�u�Bu��f>K�=�߳��n�17�^�������gBi��>�S���ݗ�#����J�Ӧ�E������ܖw_j�������e���-�Y���``i*��-�=s˾��ޥ��o�zD���BY��!0��fbؗ�މvg�z�Ӽℨ�b䇶l(�خ���Yu;:z��Bwr�G�?<ߢ.���ܽۋk�F���0��\9�E���r�0j%	j��wtIɁC�kW������U7��湫���΍e	�Q��Ⱥ\�kn�l�c��Z�c@q�����6*�����k��mi�����@PS�-�CS�`N��;nT����ځ�{im��k��n)�������O-o�X϶�٭�P7�O��v[��a�׋��ܪ���p����L�kk�7�Rmčy�hV�ҽ��_-���}w���c��v�jY����Zf��>y��7Y������zg��=6�z�yT#�\��4#v0�_plQ�=�Y��bN��T�]~��05��K�����œ!�i��{�Kq|���ؚ��TN��5�8��#=�*:�K�V;0�gM��0���^с�c�����pR���4���P�7�X��6r��4x!=����:��5�Ľ	�-��b�;�!�������y��|����Q�n�W+��R�t��`�sf�Xu���?��M��r��U���&��VH�B4^�|�M���u��>�}�t�BӦ�IxxN�;��Ž�Z��ܺK%�9�a>Z��9jH�&����_�]������2��Q�X����){1W'���p7P����H�M=<I�(g���D��+����F���i�y�p��.]z^YL)M��.T0��������o��[X.����A�7�����<ޣ�
�
4<����t����W����&y�^���b����k��}+��o�C�k���렏�*�B¢_�$(�7�q�����=�h�s��*S=��~���z�M}M�|é���W�?�*�#�]%d]j������69�|�����{�{��[f8x�CZbG	&m�Оza�j�p�x����ɞ�����|����s�"��Ч�����?bҋ�x���7��	�޷�dM��x�;e~jg���k5��@ܷ�9�{�������&}�?4_	�5"m��V���s��zw��{kd�lTّs4o�'���q-S�w�ؤ��fw��Ζ/B�7��vyM���4+Jۘu���l�q�rӽ��q}ٕ/b��T>s16x���m>��2X�V�tWV�J�M���il�[Χ"����f��(��-<22闄��WR��h�Nq+��S�&��Cc��/{��/x�ݼ�r6��j��g�
�jû,�)���C�Y3GXI���hη�]]�^|JF�i���z+�u�-M����u�&,Ǵ�K��1��J�b�W��L���v�sro��"J�9V�ro�Z Q��F�]�3`�3���h7q�ݥ��N'�/l.�iͭ���=p�od(�gA��k)Ugp��w��A�p<+x˱��>V5Ӑ�7MU�H�U巄E�uA�y�:�Km��6;Y������K�����:En�Z�qJ��:�-�b��U`���x4�(��s,�McB�V��Џ+du��os����e�fv�ˌe�����F��=�v3&���ڹX�-�Zl���0���+cxjd�nu>��i-�Z����
�ޥ�+}%!�,��ݛ�O:�����왌rk7#��\��㸲3&��Ǆ�#]i�E����P�vj�3c�ZZ�N:V�,�`O�ܿi�eS�$j>�B]l�}g��WX�x)�a��dC B ݁����#��#/$�rb��P����+쎯�Qb{V�
�l�t�9��A����سV����z�EDE�V���w��6U����'0�ӄ6�l��;]�YT �
��M]�k{1E!2��
޸���B�{c6�EY2p(4v��b�wJ�3I�ZV��V�|�p�-���r[O�}���tK��Vv^=j���x�yKe|"f��Ԑ����;��Sx��odDb�!^�o;��`�lf`��u�*���AKǛ���oV�eh(9��
Z/of�Iq}�T��i]!J����ͫ��s W�	N#�ʷ+̭1*�﹩�f�`��ew
���{Kq�sf���*hh��{��;�T����z2:��L�Jf�8{4�3Ki^w�=���Μҷ��MV;$��ΦQ�J��wf��צ���BY���5@���<4�5^7�čk�)%�`��KQ�2�r�n˰�n�׸��)Ĳ��G��u���m�r���X�\�؛�]�m�ډD��`����E��ޓ�8Hw�x����9�َj��x�P����W1��c�;����Lor9q�X�6�ji�����k�Ywk��hU[�$�qJ�����k�w��23�d���[���3Q`ޜ믺qX���4@�f�;�V�N[U�;r[z#��������;��;}����CS-�U�(DNw"�A՝�����-\S6���f%7/�������k�W9
%�tr�\IP��ː�����-�r��(*��7��9�U��"un�x�(��"���(����wr�(����w�Ett��8ֺv���8��8��q��qƸ���������IFd��
:~��fWH�gtw_�^�k��++#���Y�5����Ǐ���q�v�8�ӎ8�v�������+ Ȟ@�$���N�/Ӳ�2��[t�GQ�]eYG	��VQ�vd���PDG]הVW��QGtI����}�.���;�����Yt^Y��ʼ���D�8�;�gtQE�yX�q���nw��w��w�]���}�ki�j��JJ:7�K#;;K���mU�VTT���qkn�:�������vAS���������Ί��q��Y�3QSc�(�c�m��%��^������l�����=Ȑh\Q/?�D)���K�C��M��&�Q���ii��#�^���7L�����ր�i�WM�ֽ�^�z!ш��/js��ȃGwko-�y\�n��<H�z�+�d�$-��P��l��D aH

F��dFh��O�%Fq"�,�!�"Yp�a��DrF�"�h�d ��$eѽjlֵ����(�|t�C GN��|��<���hv�������Jv�s:�D��I�F-7�m��������f���p3�ӄ�Z������*�E�<�^&
��:��G�f��4����d��wU>������65����m
jO=�x.��m�)B��j����:���=��Y���o��ug�*W恤����~">㵌|]�@�.���Pّgu\F��}���y�=�c�h%+_��@v��+p4x��'�OCk�wB�v������!�1�t,η��*�O'��5��t�פ����
\i֬�_B�Zn.`J�
"��?�بSV�sh��QiAc�!@�,j��66���f~���\�G/f�(1z2$B�O	�d���ϝ�1Bl��օ@�yڤ:�8'����I�ce^eV��xgAk�mn�^��!�!$ώr��+�0�]�K��?���A�>5�-�T�{�}b�"û��ez�������������|B;���|���cP2�/z��\��i����=qH�^��2�OH�f����gCws���d����fOƢ���q��=x�Q�������:��"��]�_h2&"�6���Ѿ�L�]�z�i��5��?j��lY,��Rm�lb��s��	i
E�`b�-�y�D4\�M;�։���Z��	Ұ��L�N;	2��V	ܞ�v�\\{:�(�h�i���#���t�t鮖IdE:=���jS�|)3u�,נml��x�{��8��	�>}Wɥ��v���o�<kn)j���1[(���y>�wk�w����-�5�!��zTf�o�t��v�wiI�m~WBˌ�<�`;����g����
��2{ �6j�v
���gg�&"��d�U�L� )��נ�b~�}[�o�r9^�g������W1��1,�w5�CK�6Uvc�*.zNŞ�ȚTֽ�k«:ry�/#4z7]��X�\V�M���#�x c�-mt�m��j��R�\կ���%�Un�6��V��i���-��
�lO�ۅ�Β9��)���-��>�a�`ˌ����&'�͵X�Z�d����O�y�m#6���ux-oV�sJn|]	� �!�:����_��_�l`E`f�p7Mȶ���[q��.f��:"��2��A���Y4��a�Y�F��7H����1�X��m�Q���CGouT9��Ǯ�"�ݱ��}�d'��^]7��6�KMto;v8�L��^U��j��������f��^.Y�ӎ0�騥���H}ѵ�`"�'�3��s��&)6�6�N��� ���-\�-���ji5�>_+���1���M�����f]_u��]�a���z�Y.nԼr�r��^W)�j���Ϸ��nu�{�ѮN���}'��t$t鮘���V�r����{?���^�M�VCj_�פ7��U�}�].,^���^���P؞�<�C;&"Wn�VY-���]x}���{�Z��g�#��o	gX �ȵ�\j1^���Gb�Z�m�js�ѝ��/Q�\e����s�Fh5Z��-��W����\�#K��
��ޑw��Rd�ɉ�u{���1�H���r��]�q��f{�X;Ȉ��5ٰ�����tA�O.���2�a'��?<}��ZO\��>4PQ�/Mw������T�����a-���~m�����K�Ks�X]�9>�xׄ�����Q~t�~������=�&l�ք�]�摫Nu��_�u�L�>�s	��h�l�=	z�����f�C6䗵�`Qyv��5���.���3�g'߼�$�y���b��k��/nx���n���E �vG|b�+:9w�by��٤��$o�F��Wµ׋�G(V��Z��&#}^�������@�;[���4�󿾝g��X<�x�rV�du�[Q:��5�.z����s�,m��fy��?�{�D_s�s^1���b7iH��E�Qr�h��ڐa�E|����|ev�.�fs���tT��o���HEc#x��r�mwz9�y�ٯDt�^���`j�Nj2�'(�ԇ�=ǏN�t޶]���8�i��C34]s��Lh|��v�3%�V�B���y�7!>����]Ӧ���	$VDTI8�����m��K�k�i1���7�ޘI��uyq�y��c3$O�\���%<R�1	i��{��b�=�*q�� �\3F0P[���3�옦\��O�'�GA���ݜ�0����^�ۈ�֠j�"p����|�7ߘV7��A�R[��c��UYӜ�G�c�I�I�������w�ı��F>;����>]k�t�Tfmq���u�٢��#E���<�B���k_>�ǡ�3C!��Ň0���.1�1��F��4�Z��)y�|�ۊ ��'��w>5����y֡�ͽ>x!��3v#���MeV�=g�nsA2�M��}��<��?[ɧ�>*�Y1=9�\4�#3,��������;f��ݻ���C��-���"�����?|�E�����!�o����R~`�uj��@�su�;G�^(n]�uݛo��ߠ��~U�������Q$�7x�7��i��G��A�w��s��Ȥ%�g]cWA�iz�}sQ�>d�D� �����O�B��>�n�����%<�M�oN�N'�˺����
u�/#�f�an,�g���Rt��rq�R+��r6����;�v���4���0�52�-�8gZ�{����Ѵ���aE��EӮ6F����x�&Hw���;�73��5u��3��_	�5��N��BHA���������~{޻��9ݫ��������N��:�^���$`�7~p��q�=�}vgl���q^�o"�D�+���]�v"��ފ���_W!�l������۰���FH�6����-��Gϩ���[٣�����8Q�7�1u.T��m��@�!4����c�d���2�)�����Rkҫ�훣m����i�Zӟo����ڡM5n)b�f%��J���Ve�>N���J6nmM�eNd�Q�g�f���H�B ���{ɑݤ*DfU��v`��j�|W��x�Ϸ�J�xD�&���m�gS���64�}�H��˩l�a�t�G*�)≠�0\�u��Fi��Ͳ&-�\�������V|Ϫ����^��n��Z�zP��X���t-I.)ɐ8���)>��RXص+_�z6���G��'�t���WGl�MxE<M]��]Xk��P	��/�VN ޑ|���W'�Q�[~sCm��k���1��Z��y��Q#���{�.��4{i��a	/��=�����/�[<��:�	F���`BƩJ��LYܻZ�#��E7���Q�򭪸�=��L���|o7X��J��Z]X����|�rM���79�%��C��W�DVa�/�l���s�J۳GF�]�Ky��PA���i}7mt4�Fk^;Ӟ���y�o�9�>��A㶺�@��5҄�0o�vA�|��a��H�A/S>g�Ƣ�J�p���P�ǧ~��+���}�gΞX�V�j�A������h}�,a'����ҟ��Ȇ�~Ox�6�m�֘[����{N厼�����Ԫ� �P�����@��� k>����|���C#,ξg�+�P��ǵ�&�Ll�l��W|�(;���7~S�VƯ���Q9C��_[��);�}�|�!9���2R+2��%\�x	�C���ހC��'����Y�����;k��W���Z@��d�cXW�W�a�=��N�!�f�Qǫ�E�����a�>lL=���vofS�u-��%�ϐ)�.7^���"��l�g�9���%�fd�!)��Ĥ��gq]<(�v^�onTS�`�E�s�o}�Ȫ�+�|X�lQ�'�OJ��[flşrVP�ǌ���[���l�SRӔ�o�$�
����+�N5P5pjO��1�b��=�6P�� r����<�s�>��u�)9��/��n�b�ֆ�u�e�׾�~j��v���]�(�my-�I����b
�ך�m�ZW�%v���%�r�'N���'��]�r�[�nN<0�>Z���o���R�G��m�LY��Pc,Ʃݔ�p��c�|�%��w,9*�B�1����.�7�xH$���8��gλ�Yּ��~�t�Dt鮠I	���;�^i�J����7|68��N��}�w>P���^ׅ����&1ο��vN>��n!�
�#��2��4}3�v�Ju�>@�a��p34%C�E#�4�
ltݎF�W<�ʳ�e�j���{����<)�Wt;d^�;�V��1�X��wT����~My���ζ:���f]��2��#(k��M�FH�y������~ʄɻ�L�o���e+���+�=�'�?f ���p�ׄ@���y.��sV��*�Wu�y��}(�n���XJҚ9��6}u��4�����ql��������oߚ�KT-����Z��7w��:���s�OH��������z�ה� ���:9[��{��iw2,k��<�5ݺ2�y���\��-�CY����8�j9�������~��z�(����ڕ�gl>0	��N^�;@��zC�Z2}.َo��1{�`��1ÌUAn�\�������.��]�/��ڢ[������Qo��zo��G|dH������fG�2��eK��#[:��N�_���ݓ�L_�OR6��6�h?�-�E����7f,{q�X�ek+�[��0q�U�[�f�����^��!�a*D3�R�qL�7z).�(%Z�2�t��r����î۶t�<��ҥVm쩸�~��G��P�:k�	$"�@�7�`��R�׮Evh�
���tOM���_�1I�7����hY���}�i�f0�5;L�:k27n���FU�_Ŝ���I���`s���}���$���p!�\�������/8(���
�*Qm8���Ԡ��M�y�/Uk
j�bz�;
�p��������:�Dr)��\��h��\��^�H�����M^]�S�YCk�*s]�چ��W	y|`bu�jKEޝ���6��zc�u�%9f�S�Z��H��2�O��Ѽq[5�ڻ��<c2�V�����
�,]Ĳ{�§�9eՒh`3Eb�/[1��˟���7-�XYf꾫/J��d�>G0�vjhb����L�ɠ��	��'��z������ݹ4��cЄ+�,��U!���_�}>�)��"��X�Hs?��f�5�cd��Z�D)x��m��V�R�?�&�*�R�V9�W0P���ϩ6���{������RqL��G_���ݏF1�z�ɽ�*a�qq^!����u��y���M�0v�+��D
<7�����n�nK�[T��Zsr�GQxeg�T��@�z�߀�l�u$��V}�'�gw��[柆:�Z��턌�AM���OX��E�B��j��f.�R����Ǌ�۝K�2�8��%ŮL�u�}u��L�O萁�MtH�c ���$Oي�������D���so��M��VIM�w ������r�gL����4� M~����w2�z��ٌ����1B���8��<	��#�[x�+6�m� �w(��L%<_���!�̠���}W4ɤB�i|RXw9i�g�e�AX�ʫ��Y�zD����# �����������8�^�w�K�{aa��=jq��S_4F���YU���{����-}9�'��]~;��%�k�+U�G�Ƒ*4��N�Q��lzkٗ)�Dsw-�ݝ��,��1X��F�r,aF��Q�gO��o�,��Ȩ1�};B�/Rͽ�g:��C�[�v�b�����=��?���"��9�3�������֛9�����X��.;��N������^	�G	�x��X���G�e�Y�P�z4�/���ı���e���l)��AU����%�Ζ/B�K-�����Ozj��/�Nb���.����!#���ȼ�ջ55��K�x(	�l��XwD&YI6�xyvO�4�Wdn9]ȵ�ưylH�s
*3&z�ϩ�>�X��P�t��0����-��ez5���r���F*ib���^M��9Uy�s��?+l��e��6p���3L���ܶ=�U� T6�;S�wA��~?�$�"N!g;�{���C��4M��x:�������;)\��k�q۵�ro��Y��[׏�9�����a�� �>��/???/4�D��I:�|�����y����W"y����N��
i��zY�3����j�3�IQ�0D���ȕ^+���L.ބ)����{�S�/a�I��~m�k�Bo8f<���4�JqdָQ��*�=j�{m��_*L��L����������4�����9�ۙ�EF3���/��*�FE�0�l����D3�8T$	����*e�����7xc��~n��0����Y=z�	C`5��\@j��TP��4�~1�t��p���C'/����,�n��n~�����|E�x~�7��0�����ʄ\s�zO1�1���K�y���Wfiܸa�y��O���	����=jZ��lw����	��`PauÑJ��95��N���{��-jV���@6�	�����26��}X^�����@�m�xf��;4=Տu	M_��l�6���\n���tfW�H���K��M�0O��^���c�_(�[��*c����=�+53=;� q��דӔ��E��+�PC*iĻj+C��'���4�H��m4H�7D0�gYdu�W��_8f��v�ā��$,�ۿ�����N�������G\�9�]r򤊉״;v���["�0sL����FP�b�/�[��D�Όs[��������i'�G�b�<8V�f�Ǐ
.�#J�f
f��"�tYAN����Jv�n$��V�h�lfյO��C8�{V��grB�}|����q_�1wf���*J��na}C���p�*���t`�6fW�<�tZ���÷(R�>޻�����Z�y��<��q=�� �љl�!��@̆?���q:�X8�F��\��L��8ʇ�9	:Q�!��Y;+h�۳F.:�3�w�l�p	��������M��ء9ͥ�jt{L�ch���m��u��u���;���[����Ƹ���ޠvAN�s;��ރA�U�jS���Y����_{�{��Mg5T%�\�@���0��x+G4�jcf�9�Ž�R��tP����L�E/2�fM�����Gu��7$ˮ㽲����Y��
���'uX�1L����YQ�R^Z���є1q	��Awj������|�u����@���齀�+�8_^��Wo]��/���R��y������3h�����p��˾�4	|9Y��K'L=3gQYX�@^q���M�f�RM;�|]�����F�r~o�g����YÒ�hq=C�?���;!c�{-L���QQ1�d!U�KC���tEP���Ц�$s�/��wL������nn����v��VW]UE�8:\��Q"Zm0� �c�RO�	�I�]v.�X֧��2��#��	g����XQ��B�[2`b�)�u�ܢr�RB<���t��:
6�ح ���t�n%�{����q̱��q�+A����1��$3�I�y:�C�9�Re �=�;���M�內w��r��<�ǜ�Z7|N��0W�T~�*ȧ��:�Y0�Z���S0t��Pg��Vz뒻k��v�s�Ȯ�V�����M�]ً�|�	U�t�I��V]����#}V�!ҟi��ª��n��w�{`��D�*�K8��4J�rb/>�Qu�cv8trv�c\��WLGդŲ3FnXYV�'�]8v`XZ�;Z.��޵X��q,�1��U����uv���B���T�k:jXI6��YY!�ouμQ�Fna�֮u�.�&�Yy���<������	��4�w|��r��̺]�>,mԸ�
��B�Itҕ*����(`��ʊ��z� �C���'�[�jsV���E���p�:b��&�`)��vNV��录�J9N��/�-�u�q�g0���R��S�[���}}J؄[Jd!��ߗ|����h�[�Y������Gܴ��
��>[��X�Jа$��t�������q���8��5���;v����y��k��'|��#2��u�`H7U����k����o_]8�8�ӎ8�q�N;v������~�_��U�v{6�i9ۻ�Q�k���˾U�'wȲ>V�p]Ķ��/{I�S��^GgQ�t�mf;3�H��΋��6�V��.�.+;������ݝgOv������e8�Z�dt��k�v��^XGt�#��|�'dyvqE��k�^�\t���y���Ŷ�����ϧ��'�nD��I	v̾{R�gY������{f�ҷb�ߞP#ys����|��r��D�Nۚ��u�$�ҿ}��t�Ӧ��HH�a3���Ժ�����;�=Lt!uu��(�}E0��3��C��3'�U����q�᳑+�Ok�Ӱ�L\D�{/��o[�r�U"��Ɨ�j���S���Y�{o�>�&d��t =�~��f�=��9�YB�
������w�������R�n�3��7ɟ������
�O�zy�{����dSmUn�'�v^�y.ӯ�oW��ؼ�+RW�W5a���w��̽Oa�U��{�PxR��t�7,�^ڛa���mm;���ns��dA�w�����N���>�f�_Hf�Ju��ހ�����C�E#�70n��p�<V�<,nt!���^����9�mb-�MwK��f`��9��������@|&U_�mwM��=ې~�U�v@�˞7���y�KMto<�����本3}x��owfd3����I���=�X���<�xD��]:��ylf7O��g��7Wv�n.�t)jy��y����e{��+��?J�U��A������,-���i�+��V[��ʇ��]\r�[z���������Ε��
}�.�6�aq�,�y&�mq�ο��ܾ��[Fz�T�:���2	�Ki�^k����p.�`nT��W<��n	.�k�W��R�M�tw��j�5�S���a����=���t��oy��u��8qOP�/1-%�-�7��P�m�x�OH�7�#:g�5`�yt�N(I���>����9�׉2����{���l� �͌��TLs�2XH1Bc��N?G61*fWvwd,�~f���:���/�)+��~���͍ӊ}[#+^8�x��c��Ļ�d����g<i���U�%��Pph��:�L"y�g�W�y
�|����Ǿ��k���=k��{f@�#��_W?�����b��^�N�n��ԩ�6��Ř�%毑��`�������p�#�ۻ��oC�3�hD{!��N�j���B��ᥙy�Y�3��|����</b�m�c5��LI���i�3�:���H�6o{?1��o�:�9ݽ��L__��+�^E�Q�	��ې���C'��,��
U��3v]�<&r�S�'1^�5c���6��rXF�	����8���6g�s�Oz�$oج^�f�K��C&�L8,ӧt�S�^e�v_3ϰ�_#�=�� f��˨fz���5�?[�K��{q\����c������XQ�.���ݥ�̝���N>tj�L���zޚ�QAqz�b��K�۝���J�/�-��Z;�ޅ6<z�J9V�	��F�K�OS�9��}���-�GbƣJ�,m�`b��ٚW3��;�y��޼������U�h�7�ߟ5說7�����v�������0c���Ƚ�Yjd"�ѽ�@^c��ʝ��ڻ��X����~bjF͈�6`kA����ߠ<�v�)����խ��27����ƶ�A�Jn��	���R��Q�0}�z�g�W�Ԇ���K�n��^���b���x��a
i���P�6��ZY�E���w��wF763k㸶h�cv79#����i��%���Io&����B�T�qo�NK�{ :JK	Z�:��ͽo+���לe����*y�tm6MW��$~Q,��1x��§Hb^Y>�oX�*���{~9�z�Miv����.b�n �c]�oK�ƀ�Hy��L���~��`��%F���';���ucx���Y6�/{z��ޚ��l���'?(��~P(F��vO�&�ۨ(��	p���Q[[�Իn�,!������1�x��-%�ׄG�#"&wʴ��\�Z{�;�6w��5����@�8�1��^w,�q�6����Bz0���a�|7��x�yo�~���zs��-(@e/H5����MM����,������L0B����G�a�؋-c7S
�-��^��Cf��7~;�z��;�x��/ƺv"��{"�+Hf��R���
5�˺׻���B	  R���#��֗s�c]z't��u_[\
�郎��"�cB�N(�9�d�b5��7�;�P���������������"R�,���驤F���X�	�E���)���a����bԌe\��c�խ>�8���i��m���띎u�j�����0�K(�e|�}.��|���=����o:��x�"X��i��v��C�?��QRw�r�:�V�M����L���P@�L6��/����	��/[g{��k�UPK��Sm��aQ}0(^C��w4ԋ�2kV?/W���veV��������v�r���ۤ�����v����y`k<��h	4zv���T�Uс}�V�L�Z��-xX����8�*@���)>��(�����7>a���'A����}���+� o�z�X��>g��Y�����"8����s-�27^�Q��r"��K깬&5s+w|qh2��
�;y8��z�S-�jD�-�m쀡BO�֡���q�$��'�7�V �j�PV`3ttzD��rz��t�/-���-x�6n#)c�z33o��	h���fh=^���� ���qm���y�P�	�6�zO��w�	��uQ4�׷�(q8��J��TiW
G{�׳�i_n�;����6�Z�o��o~ �eŢ�r�]H��ꓰ�`�I�9�b7�3�-�բ�d�Ғ��g]��ؒ4p6�]�m��g}�;������2�=3;���_�����������Ne��Kqv �7ã��^�x�ok:OoFZӼ��'��g������a]�.����h~ڔtƟ��K���}8�l���ƭ���	�b����(tö�<3eC��v.�l�U#U���p�Z�4���͵	q��������ع�,w
�	_���[�*����-ys$����
Ĕ=D�X�l{?]�yi��O����L4�&D�W�K0ƥ���\�J��*mq7�����:Kj9x�N�Ш=L+��Z��k��ú�D����&�a�§ι휪ɩ��w9TҒb����_��#=ߝ��*+��5e���
���o���	���hy��Uf��푬	.�A�X/�h��ceG��׳�39���:�Vnx�� K��i����y��lll�R���<������<��QI��H��*s��q ^Ezu����$4�o57הm�]'�0��l�#"؆����Q����I/K1�T/xZ�a�U��ęC���`�C>T�*��5{�9aO�O�:�/���]�q_�k_�#Ñ��>m�C�����V�c�EO]vlf����]UQة��o�6KUٕA�һ�
�U_���Wdj�˫�Gg����Auv���[�U���W����~̤7}���au�m�u���ëPuvA�5���O3��m���e�2`�4�\���}L�뻁�}������v֭kQ>�do���]s����6|+�"��}M�_�>K��?���ߘ}����v�w{s�`�ۙK��w�T vD  �����~]�C�F���:jr�E��Ւ�k�*�d�r��؟2/[�����x�gf�G�Ѕ���[XčK%�gб��l����!�3'�!F�עaˢ��f��[��a��|�sOH���f�U^��Q;�x����ܾ���d��d���i�|ڽ!�u]R��K�k3��ye�q��@c��Exd��oW�
qtN�����j���\9j;8��ӱ.IkYr�ow%�?��&��1�0�`����3�{��������o����G��]f������6r?N_{�;�0y1�2�l�p/�5��5�U����^8��GVJ�lM	�ީ���,�Pd4��c�4'�gO����l`Lʛ`}@MN1O��2�Ǭ��p!���x޾�GE�����1u˼Ӭ�\��Tzn_��<��EC�<��!��|^�ų��k[r�Z��[؅��v��ѭ��Fi�ej�wy��8�ꗇ5��I�Z�+��S����c���O��/�ozf0���gk��l��W|��]hشyѭ�Gv�u�gO7:��O��3q�v�y1N�C�v�#��ֳ�3r5��ڍd���#������[k�w`ra_u�d�'|ׇ$ׅ�Fp����ֿQoy���f�bu�)��&�GN��5uF�Yn��J�6)h��=������v��b�m�y���_Bm�Kz�V_�P}m���kR�Z/:��y���l����7[�����I�tk�jj��q)�}O6�ز��*s\7,8<5��7ٵ��/fò�m��P����I��r�Tksk�٬���s��>�&������y���|�μ�#��G2�Ɍz��%�?{$Nʜj��&G` Ԝ3vl|�B�"��]�X��{���!ٟQכym�Ԓ�x����;�ݨ�x�e= �l�݀���ݯ>N��1�pN罹�vf�u��Z�a ���_Ԧ�H�cj��B�hh<�v��Wǃ��p��H��{zvj����!�K��)��2&�qqDڮaj���k�0X��׷��y01�L�I�Nѷ���"�Q��1�b ���{bѡU�x���l�z	Gs����Z���v/x��.�����}���Χ����h��"���#K�C'���bJ�r@�Gh�1�2^�"V�Uf��"Yy�桮A�5C ��!����n;>.�V|�58*.�:�M;��ݳ-o�M�2����++��]n3�f׎�)?>Vm<Z~��ge��M(�.��3�� h�C���,�u\��|	1�z���/&�$F�K��ͪ-�}S"�f��wR�0f+
�(�eڼ���D�5����{V㏦�v��=�^yyxx|����C�$uTц�����?ޣ8���P'<�:�_�0�k�+�`X{dn�T��osM���0�����N�)d�6pK����_�=���z�k�*�ky�?~���~C�.����!�"U5����Ҧa5����*]�|O�Cb�$`���4�3m	�t�y�%��-���x�����W�F"��^�=���E�p��r�ܳ�Q��o	�f������,7+OX����\p��~�ڪ}�t��	=K���)O�a�'��ʉ����4���ɅQ�]4�솪���b���ZVl��ve �������,_g[E�.��uҽ�5�:�!�5��oj�9�|ٚ��}����5�1�ޚ�D9׺��z�6.�oi�xa�0gk����%ۢ�	t�c�fYs�b�_��m-�`S���^�Y�*�v"61�0���kk���X�l��S�����L
�M��J���[�����j�{h[�ҋ�l��u�������6H����:u�|�A��{~��؟��+Z�)�B���ۓ8���\�3
�x�Ӂ��VHӼ����F����'�f�]�Ok���MV��E�\px�ӧ�T���u�MTd���Bu@gG���Wûn�[��S��xo��fP��4	|����u�n}��<���� ��� O*�ȫ팚�w��i�~h�D�S�Bv��o�Jy����К�]����ps#uڨ����}U��|����%�_����'�O6�;�l�j�W�����p�Go&�[W�\��pѽλO�v�����a�3q�wF�$?���򨦯�E���c��D�͒�m.���Ka3��]
���:�	k�#���#ޠ�����Μ��}-�$o��Kh[���(�P�?�۟K�{�z�{JU�7����,��2��5y����Q�4��Y}�t&�zF�O^��e8�h��ٱ\���f��/F"��\I��ߺ����<?%�ܪt���\h��MB\��;6Q��>���x<�� H�]X��vKF#O��=���>?��`}x-��bx�uV�����v�E�~�o��?`��2��ߪ����vu������2����:��ȝ����(�]�qz`������GWU��;r�j"vbs�{nrlxX����Õ�e"'|�9RW�Pj�_|`���L/�K�۫�4��*S<��ɖx�rJRM����������Fx����g��%<��y��y�"8N�2�v�@�#�g6C�<˗��p��5�{��G��!�b�6�$���Y�
wY}�[����.��a��ɪ���FJ���� ~��yx0|������<��y��a�ҟWYJ���X͎MVbY6�+n۱l��k}Y/-B�21.���;/n��NZņf���qK`&��d��/
��Cv}]�����%V���`�Q��V�dna���Gւ�������U1���%�_�	oMl�l���a�a�\s��Z�LJ��A�E*���m���G�9U>1uR�=@Kw�O�)��yKc팎f��Ky���j؁�ŗ���0��門gZ�釺����C�}�(u��L�s�^���*��=�U�P�������A;�Ԟ~�O�������Lc���(r�١#����>0�kq���M��B��MڏK�z�O5��w�ȉ�w�CYnq=���-A.�9��9�BƊ^}��q����5���>ŧ�"���qB4�����F�W��|�
o@�PXY��ٯ�{��%��k�Z�V��kI�����v�^�5�g�16����i�B6|hW�`�g��C�t��5Z_z�ג�vkBm���[1q���9@��v��ȑͿ[��Cu�E�;�Ӓ��3�@h,3m��󋁸+��=nE��䥃z_nVӁ��N�' �O����7�p��L�&����G[��2bΦ�6��j�9&�Վjhޮ/.���]�#�ِiZ�`X��ڽ��b��wJz��h1��UvwL�ܶU�"uqwb�E����[��K\�z�q�X!�3x�:K��IeWb��N3iR9��]��6�;� ��/vmh�]��]�6>}���{�r��k��mo�b/2�E����g-\�=)�<����;e���J���7Z��LAɘ��g-�wȥg��p�*Kf��3�չ��v�y��'�QW7�6���h��sN�%�s_p"�lX=��-��K��;��0F�̮�p�sn>��lZ�y-=�t}��s��ω8�Xj�c\����a�zz6��{nc�,�[�].
�bVpG;uN̻a�V���Kj�N���Fයv^�ڛ�u��c�m�s�J���;���UY���s1��l��y=|�ػ��GW�5jZ��ŗrP��hqt�݈���L�×on�=���!{�c�o������f��>��Դ�6���Ϊ��d#�U�4q��0`��'+�Q�#S����l7�of=�]%t�</�$��ͳֳwS�����2Q]�}&;��+.5��ޠ)����vpV���1�P���/Aǧ-{�'���/��k��kN峍�E����a˹!��gUڻLVZ�Y(�K"Va¨�&W�Z[dզ�ܦRFkȕU�\�e=�,��7�cmm�W)Փ����P2�k���n_p[�<e�L��8�l#v��j�sܭVq�*�Tw7Wc������VEAo��x�֜�!
��8E]��늚�7'01ڭG��Gٍ����s:��H��k���ڳ՝B:�;�;��l�%��>=S�ɋg3�����7��s�w`�Bc��&�xb��K��6�3��5��t��!���aй�h8I������O9�Z�-��d]\vct���ȸ�f��N������{;�A���A��i�I8-l�v�Ǘ��&���h᪛������B=|3�OV��F[\��3�L��Rup��B��n��eY�$��p(+u�w�Rt]�v��{��Y@.� ��7�w8�р�<4�o�.��u�r�qo�j��I��+�7��n�A��r�v�e�o���ݲ��̈́M�*�B��+��eL])^���c��W1&&̰��[��8d;K����Pk���8Ո���&�ة�����t�h��fö���Fg��a����{/$����+Y�u4(W;��7kAe�h^�r���^X�v�]ۛ!*BΣ�g�Fm�`t�����2�
{5o�>ڤN̖�]���[{��C�x�N�f��ȡAH|r'G�ڎ�e�HY�:v�����8�8�ӎ8�q�N;v�zv�����B�JB W��!I�(^���:v������N8�8��8��qӎݻ}v�׮�	By)����2�츯�����^�q^����λ�#�嵅��9�٬�#�6ډĉ'm�GBG���O��Y��⢊*9��+['qG�������m~�O�]�O���$\���	%F��+�s���r�ã��X�vgG���Hr9էy[��� �O��r**#��
�)�
9!&HD*<U0��AV!��&����ywڌ=6�a��qu������3��:�0�n�����SQk�=�u�} �����D���pHIuQ����B6�!-)� d�@h�o��+��� Ih��cI8$f�@�"�q�a0 Km��R�F���+ġ�}����MGN�� BBB'����}�?/�{���;���!����j�na�΋;{�P���<�����pG�Z������c �=�<��dm�4�Ӂ���Qם�U�1����ύ|ݗ���߷ɍ-~���L"1m��7�K�s��y�P�(�����v>�w!c��ƝMk��<t6 Z�>����!���V�4��P���k�^9h27��X|�%[��]e��>�+��^p�����Y����|�GL�������=@�^*S��]�O�����6c��:r$��՞4�ɌM��}�VaD��+�Z���iˁ�At����a��u���]-wj��Z"�ҿdx߱�:Y��f���t��Sw���v�L�����x7]���s&��nc�-�j���|�ū��Ck���T�o���f`ͼx������6Kyu#[�n��4���'Ϡ�ʫ
��ˠ[ёS����y�I��tuW�Wc+�hJ�YP�N�0���5��\�eu#��n��cW�+r{9|�����Gv�`������g��E`:_�)]�����-�ψk���2\�BuvM#b8i!��"�f��v�@ƞ�L�j��;n�n���MI�[Ր�:� ��7����
�x��I�.�[[d[�����@���>~�?�7�0o�`��J�SL�~�FyA?���(�t�Ե%%�^W�kU
�OY&�fk��!W��@��tz���3��q{�D�+IS<���T�շ�}�E�P�a!2[�Dg��-7�ޡ�W�{�أ�]Y�%���2��;q����H�X����}�4���o�䲹U*���k�8rsOk��XM�'�$A�F�������h'cE��+&��dLe�8�����C�	�ʯ,���6d^�9�W����l�k�f����6���X��g��;\�f�H#�&�8���i����ƾ+s��9�j�>�=16j�.:�֗�����f�R��r�ۜ�y�!���-l��-��Ut$��O�&"Y��#7ӣr��
,��������D_�Z���f��`�Wc�WНU�]Ɯ�+c����_Р
��+^���I�Ƈ:�^&��P����T�.ݺ��Vy �1"e����xϏwj�U���o�dB�S��ƺ�1�ꬄZ��%y �s���i-ʰ��t�]�l��,�S�o2y�|~�<v�A:k�#"�ι�>?I\������/�5�;�=�QKv�{E[,n�jTg�}��w����Ɉj*�Z��$�����q9ⓩ��1hw�ìȑxʧ��f��S��h~������SY{�M!�?���e���52X�"l�}B�6z���9w"1�ņ�����1��|A܆@����6H�;��+]��߳��Ћ���j�3-�hoʟ!P�wh
�.�}_�`�o@
V�r/�ZPeXy�����3}��WS�V��3�pό��5�צ:lER�s�����Oen��KJ����.q��d�-�\dDjQ�{D��iì���nwH�잛��_����2��)p7�)=���W�z�]����}qѰ��uH��k���}���c������f��׀~��Yr<���ο��U¯��v��!c�j�k�^x��4�-Ze�_tg͉����4Ix��y���Z{�����n�Z���a���w�ް���C9��ޛj�%�s���,�H�ٞ�D}/�go�m�&رv�.�0���u^t2�JA��M{�2]ap��B���\�W�&�t;��Ϋ]���ro�^5�:j�y��9�wd�pϱ;�2!�%���I��{�����������y��F?��<�D���U��W'���loV�y[�{��&+kOf�<�y��}�쁦P:ٓ�S�5@L)�*�2өQ5�d��ޙ�w����:J����O+w���/N�KWf���{��G����ڏ�����W}�채J�=�[rnr�ɼW�����r�c��G���7Dȭ�2/T|���Rv��W�\�*��LV�9[�������)���~B��-��� ��b���K-%�B�eh��"��z��'N�4��
̆��7�s4,k���z������"pp��ϳ;u��vT�n�Q>������h���\��͈��^q���܌�-�#o۳�K�s^Ȩ��sw�n���O�4�wD8Ob �[o�yv�R�.�t�Wnm%;��ɻY(S9��>N�ɝ�ԋ*�k�9�S���$^қ��ua�����k;�v�9/a�
��g��9Y�;r��������Ǚ\��{��
}=�jִ_}�]o�'0��Y�&����.\�}�κr{� s�U��ƫ���]9�.f1�&%����j�7)j]�m�0\��xf��e|�u���k���hB"7�{9�s�o����ۢz57�}��Ht\���=ΧL�_I��-���!�8�m���H�P�[��ª��9`�y�|j��|���*������1����W]rŰ�nFi��^�]Se��eUq'kAq���k��q�O��#��]
1H�4�V#��a8��{�Gv�{���v�%�Fk�#��k/�1����Ch�"�z�w5�X2S��yr3�\E�T j�Z�SO�5���ڐ��	�.0p������j��^Ϟ,����Qx5c4T��dW,myc�h՞}�ۛ�p˂�A�z}
 	��#Q����7���Ŋ���b����gf��͛ws��*���T���P�����S#/��f|����A�����(�Y��0a%you���F��3n�IΠ�jq镶�-^��$�͇cs	m��.H[נ|���`Řk��Cb�)m�x͠Ǝ���ɽ���$7L]݁�n�^b\V�Y��{:��)0����Z���<������o������{��^[��n�k������^�C6:�:8����'��h�����v�t���o۫��j���]�ݟ:�f���}[>�*]�y�Ki�7�5����y����+zG�#���R��.�h�T���0��fh��,3F;���x��������0�#.�<y������'\��>�蚲�{z�6���Tp�)�dD�#�6R��\�Y��%+c��幻Ymªn��ٵK.�zߚY���>.T:�r�	 lZS7���s)Q��~��Nͪ��פ�}=�r��y��z��]�F����!���R*�_z���ַܴ�}U\�sZcǲ4�5��cS��#~���쒳M��ݛ
�kg'9����1n�^�ϓ�:\>���d8����0��l�����6s�Ά�%�dU�a�~�ۃ��<mù��^ ����MC,v��|�Ơ�����kJہ�e�Tv"�=�^����!�����qmn=��3v�!�8n��o��w~��=�Ŕ���)V
���zo�\p��9�c���_Sk��>�����o����O1��������<����\���	 �����Lصv���\���	���?�iE�N�5�û���w��jar�f���w�|���X�츋��ئe'^�vs{{qM�2#o����g솠4Ur��>��	_��S�2��;
L\wv�O����N�6Z���ْЪ^�}Y![�Z������+Wv�U3�g���w�f�vK4��X��=Al �My�4�3M2�]H�7Zcr�\�� F���+4�]B�䓞�V
�ټe"��.m-j����[�CTs���g�c��d�F�`�4LdѼ��]�Q[�a;��IYޞ�
my����;"�E�4m)�2iޠ�+����#g`��̼u��3O5/33z`��w&p�f����ݧ0%oH�E��8�j��i�{=�Y���ۖC����So�`n#�,+Ӽ���R�O�T=�j��.��%��)ܹ*y�!;���g�7�=�3�g:�d�ﾱ-�n/F1���-6�ɻV��F�xu��$�BJ�m������К�r4<�r�B��hc"���i�CO.Dfi���m��k��t�:�=B�Ч��������^^^���}�l�ob�Fȕ���*m6F�p�`{��&*cRKf�e�bB�A��1e�fs��V�wZ��N����t�����Z?�I��w痫�%�w�=s�}�;�gv�s�UN���.�w��ZUZ֊��i[eɶ�4�9)&�ҁ^�g��s�9��1��ǭ�]Yz���:����Ȇ/����V:.��j���kԫ�K�<�=�f<뉆7z��!@4���⦀o�M��U��.�c�A{�ʶ�oU�,�;,���CU��k�[%[4i�_�ϫ�y�#Yn~6�{=]���+V�������/��ȞY���~PD�X���~��n���v��q+6��^�xZ�S��r�lC��B��M�f��Sj�<4Ǭ������ݳ��I��g2Q�y��kp��Z��,���Y��ߣH�f��o炇.��3l�$���w2;�/q^A��S>����c�/5��d
��l�*I3��K�	�[����]����-�����y
t2s�7}-i��3��q�O�C].���%�g.U�5�}R�U���<���ﮍ��Ho�ƓQ�U���z��h�f���5�A�C
�kk���ޘ�9�ճ�G�oq�@�
�^.�	ex���Ӕ�bgZ6��m�W�ڽm������̂�*��-�|U����2>-��=~T��,� �_�����P:���t#��WC[�	d���o[�n�p�8l�fb�����Gt�u��$o�ۥ��]�.��u�����T&����9ݚ�:"�(P!
��৿H{y�����;���,i͸�>x_�d��:�q/��gw�4�xEb�����d6-M���<j��wtx�VM�s��yYY����a���l��k%C�Ā���9���X[����w�k�O[��;0u��Z4sT��5E�Ű�m��6f>����5�n,�j�R���?W�Y��ǣ/�QB��"Y���h���)U��(�\���ܪ�CJ��l3�0���e?ߴ`�/�b�;'r�gʘA���G'��J���^�����nGC�RFY��m5Oh��VU A@B������*u�`-�����3�|7N���Wt��ʼ6.�dXO�s����e�n�bƊ�K������// ���~��#׋{�z�r1_�U�h�Gͅ[��6�}鶮�q=b�捝YdV�����<+�.��U���H������|#�짬��b��9���.���̩ ܚ�M�+�U;iT_�<L�^Z͗/</g���j#���t�~��
G �W6Tz��:�@z[����Pyڰ�*���Q1��6�Ww]�u�o6��<*�T��u\yɹ�!�K�O���m���ӻ�+s�Gv���J���}w4.���Z�a�[A�k����CM^K�L�������vo�طF�x��&�n�+�Q g{�I��$�*�++�Y�~�vB�NB3��ќ��Q�`1����#��s�b9�P�/R�{��g4<`�!�H���� �b�鮕��K��{�Ɨ:�PL�~��ׇ��j�P#̷�a���4��Ⱦ3�iӚ�|)��	��O�����H��c��e5w;YU�:��X5���f��
J�)He�d�5�rH��N���	�I_g�uٓi�2ٽ��Lɻ��3j7/�.֍���
�r�oj��>s�Wz;xË�}.l�K�f�+���ּ����:�6=��ѡ*)Q��4 Sv�.-i\�v��G��H�:7��r��vi����M���F^=�e�Q��݊[Z����^�zP��9�O�
�]��d�g�_�h�`�(�;ɶ��Je�]�ӽ|�[�6��Jǹ�d�w��*��(�2m�bg>����1�7�S�c����Yu ���YK^���#�U.��å�XsM�٫�tkZL��r��A��k�Ƴ�gs��I��\M�vU�tRT�[M��;��&F�nc�E�0y�Y,�������s���q�]h���%����Ow�k��Jrm�M>+����W�(�/tK`�`<��9P���]t�U��t,c�_	p泩JO8s�wk5�4"f*�/�me�hf�o��ͭ4pv��`S�FKw�C:��)�2
��v�V��b�h4c
��"�)Av�zx���d�C��n������Tc:�h�)S���y1㗅qÑ�H=�&��k,�tK��/뒣_fok�Y;�4s�z��:�M��p��xQwQnKܕ$�l���e�|z^��E����\{3��ޮ���
��-�L<����L��Oem��ym;���[�q�唁.�Պ�/E��8S]���c�%Cu&��\��rQ4�b�4"lv�a,^��ZIeT5�Ўl[6ِws|sxۗ�՝WZf��e���$oI�wOj���Vl�o;��b m�K��I�����U���ݭ��3��cf�7M���x���[�ۆ%\z��,�����uۮ��d,��c�Vc9���㫽��&=��]�ei�*#N]�o�r�����������Դ��;�B�Fh�xLʗ�jZ���6WV��Y\��r)���|���fv���G���
�Uӻ
���T�
kk&a�n����mͷ=��{��:��-����ƷEI-V�Ù�Z���X���f'�{�B��x�c+O@�,*G9����ZJ��8E�_Ε+§��ǋ%�L�c�H���Oz�Em>������'F���y��u����CR��+�a��s|�^;��T�ۉ�5�.oeԕ�]"��`�i�Z'B�9�\���ɝv��n����8[��a�#a����4�T�V��pL���37��9a㴀�i3fn5�0��uh"ܽ}΢ԕ�O��Z�Ů�f%|���M�Jn�*w)��}�ai���{.�i�� ��y\�۹V`�;�x�=���6�q�YB�n��gh���7���m�[n�+)�Y���
��@6ƺx�����ָ�8�n8�q��v���������"��"�XGV���N1۷o<|}}k�8�8��:q�q۷nݾ���<$�!#yl,� %�����䣀<��m�aYW�g~��N�|�Υ��޻������y�Yg��V�{�__jė۷�ygE�t�����O;u�Zq%y��Y��߻�`����N�u,�"�K�O�Xwӳ�lq_4���*(��8��Q�ehQ��qǙ�Q��e|���,��,҃̄�<�U7�镎�^��yL�I5'Sw���g�U+���sV�jt�):�.<'2�II��ιGF��I2����q���Ǣ�kML�ݸ����:Ӷ����`���{��0���u7����C:*%d��^��ʾ/rl���qW){z����o��3��h�@���0ao=���ܧx�D��������B'N(R�5��ot����lY��|���쿸N�o���$�ç/���r٢�h��c0vZl�~�o�E�`�޾9#\�"��fr����ܪ{:�/����Ş�rr�Dٻ����Z}��mOFo5F�C��MT��F�:�P�hL����w�]ѹ�}�ӥ�؋M�iOv�f�
sg��Oy���w�6�޸�r���U�a%b�4�n�c�z��v�-��j׈pΊn���)[EfUb�x���P���{_f1>��w+rT��0�WfչR:TR��^#v�Y�A�}���R_O���������U��,��\���.�Ɛ�<�QZ��tU�3aYBFS��ir�}^�>��#r[��f>�men��=_����#��A�/�hWgz�t��T�����ܤi�غ@�� |�֜GMEmG*�+`��}�����Z��i�=oUT'����������=�';�חR�l�_r�v�g�%KU�[4�:�2�&�ĽL�ړ�o0F��u	G�pY>�Q}�睴|�y�D5NZaU��/��M�r�+�(��m{����Q#r�<�YQ�b���=|���4/%�E��٫n2n|_����*��e�a��D-�ѥ3H����k�����ves����=֌/S7����X��]��5�!�q檉��ۻ�+Z��gp��R*<��r�x�z�Ԃ@������ېۥ�n;�]۱]�m���ȃf}s�Hl����.��[��x�钯���3��ML��?�)y����A@:�w�Ê����ݫ~$�Ҵ�,펁��_��+w�ͮ� �S�ؘey����s���ѵo����y���q�г�6,ȡ�<��Ԯa/��m�����\���*�m�U,�i���5;�)¥�oϗ�l�^�^�~�K��2k�:2�9�k.t��Jŕ��tL���}�V;�u�����\E�$�� u;z�Q_f��<��x�t����U��͊���0m�΋:�wzP��>���!����ѩx��}\���2�㝻����܅_i��;`��)�d�GL���
��/]$�����|U�@�N�bg�h�{�`�k�C�{�u��VU�e�����9 �%9��y[�CYi5�Y��Z'*e\U�}8�Dސ���zcJ�U�Ƭ��	\��~y����T�
S�b��O��ͱ2��l
������e�:�䄜����K��e� ����u	'�׍�{!�Z2C¼�]���K-(5nqyv:Low4�S��/o���4cݩ�[状!mp�5	�d���{��3�;��:a9j�L�S�x/^�F�ps�a���l����]��K;3{����nK��n�o�ёb�ߧ�H-�6��=�w~va�A�>���j���a�𖥻�ߔ,�;d�2�af�e�M�=���~i��I���������~S�?��/��gSg�b�~�B�� =	MH�]��W��Ut��I]�ԃ������A�]�W��g�ovR�=A���r����[;�C_h��Rڡ��` |v�����xݷ��:#Kn��Sy[�5�v��=U�1�q]yׇQa]�\We���(��r��?}�o�y��{���q1���P�wC�vA�"�2�ڍ�Jnپ�p���yc�a�9��DS�5�ٵ�׶����l��w�G�c����|P+�S�C�JeDl�v~����]�t��!ٞ��"���n��+�4��-0��m/2�D�A]%��Zܶ��õ�ͰGW�e��%�E�W�49�B�c�g��?�؅���	��;d|$_)w�{!��U��y~��p��)����-Z�_o���ک<݇��;����{����᷶�M*�=����1�:T�j�lVq��^��ȥ7wGM��,�t�C,�ڪC��] �zj����x����Qŷ���7�]�54t��{��x�g���T���c�z�,���kc;�)ujg��,�WSF�e�.{5����ɢ�b���{���e������d��f@�)]Ϲ]�U��>����~b6��~�F���*ւZ1�-�C���2s���#jּN1Ʈt��j>��An�-�t=�.�3i<�"��X']���ib�r.���Z�^�@����nc�g�2�B�$�25�Y����]��<����x���x�ǟ��񨓼�)�-���GԾh��}#�ܵz��sU:+*��1�t�Nݣ2E�J�z�r|�u$��M �nS�G�����vyM��݈�u��`Ue�i��p�޶ >ǧo.��*�*m��zV�H����>�$%�����=N�똝�֑6��� 7gL>ǝ������25q�k�ݍ5st��Õ�[P$���s�q*��[>��6�緳�I����GP��������V��Kԑ�&:,����;����s���Kb1틄��|�c�].���7&��ϥOu��_gњ_<ѷ�5��N5�̃U�ev��׽�"h���:ԋ�Ż�w��~=�������z�B�Xrk�6��m�`��u�˞v#Br�����rƹ27���ɇ{V���/1��l��d&�Oka�5���%<Y��a�f�.}�d�G�͸a�e�ٔ��5k��Y�sj
�ܙ2��PZu�_W���p�|�^&o�!��N�+ۻ��r��Cţ�aV=�Y�R(��3�mUq1>˾����b����m���4�c��*�Z��ȹ�n�o��?yyy///I|֞�x"8�C�
f7������2!x�������ͺ�Η�Z{z2�K�[���֬h�N�6�0k�4L�So�B�3�u�Vd��t�;�=hžԍ��Y�c{6�V]V,w��-����T��Y�^�9�d,��;r3�{��t�R��MR�w)z��b^έ�1��0�5!����Ĭ(����y+����{�*-F������0���ݩ���Yn �4<7�"�����P�|�j�\ycW�3��T��.��3��Z�vL���n���ErJ�D"��r�f8l
�+y�%ڜ�����u����Ƽ�N�~�⯎�>�Y�;/ӑ��cp�B��[��ǝ�cb=Uؼ���.�A/+i��`n�o�d\v%�go��mu���茵^Tm��)ݠ-��+��}������	CcY��^�x�R���׫q;*^ݔ�.�����C�y�d��u����J*���%����y	�d9�0\���*�x~�A��swhޙ-�弍�t=ud5ΏP�ɜPn�į���5�ҍG����I*k�6�C���q��tj<ޢ|���~?OXѨ���m��%7)���$�xQ��b;��IR~>��o�����.K��r��ۑׯ�:r�h('f��5{QEN�fӈ���� ǔ�>��Ϯ�
��o3_��P��0è5��J�<�pE�t�^�����s~�W��e��<�`]�S�>]n�z��ƻv�{����b=ƺG=_�붝x�kǁC�˹��'��B�^j�c��^��f�w��+��
�hS��v3(/��`�g!��w���5��׶@�K�Wjn ����b���V�-e뱰d=#�S�{�?��5�J�{c�=S�J��/�4%s�\=���ϕ�y��nE�F;��l�[@�ny��Vm�\���-Iދ�zވ-ه������2����=�z�i�᦭��]^h��]�K�ʝ��ͫy���=��cǻ�YoVH�Ky]� wj|ֵ=�`��^�Z���h���}�$�:XկV�(�2���r�(t�{P�z��ܝz���v�K2gk:�;NW@��-�L�h >�d|T�&˳�7�Ϫ�Eu��9X���������i$:Ҧob|k�ȟ}���A���%@����ƅ��yǟ���l�s�����5q=�2�lv'j�Fх��cW�%*e�lшx���r���b[(�@�P���O�G|��)u�����ɽ�u�Y�ӛo���n��X(ԿYvů߫ӷ��t�)]��V�w�g%ꚲL�<���5��ɝ�z�<{���Pfnu~�7^�(ק�R�	z���Ns�ݰ�;��DE��S�Տ�Z��^l�!��_��C�­��j떗����ٌ�n%�"��>����{�c��3y�y���7 Xj�]"�%$�8�.k+�xx��Sׇ���I�n���Ĩ� ��,ÌvE�2���s&��/�+2�o������%L�evў�{/��~�~���X90EL-���'�&Ԉ�GaS�om�٤B�"�x���a�cZ�u"�7.��Ӝ��g������5�}i�ZO��{雕a���M��}*�e�{R�f�od�fHvl��VwQ�x�*��e ث�i<�2�CwD�d�K3�ɱc��9U�G=��m�X_A���2Z�u��Ϋ��m.ű��oK��:Zf��}o�����<)�<�9}9��,��ğ�^~C���ܮ~���v�I������ٌ��R�jc�=3����wy�)��*ұCw"f��;��&,��]��\0�MT
�~oJ(�3�Քf�����NY=��w���a�J�Ux
>̻X��hk�W���`�8W�÷jx�F�^I��a��~��,N��Ur)]�lf|�U�����[r�֗|,�@���yK��riGa�9v�ԵJd2�P�!4>^V�4�nn��Tx�/E>��
�%�ܔ����XB�ܗ�d;�6;��na�í;��?NG��s#Wv9Ǥh��V���{�����VF�? ��hi�s��w(�׻db3o�JL��sq��6�\ż�������VVϝ���kg��q��R�>����g�ڧO��Rn^=ݛ��D�=��ճ̰�Q"#�?����%�q�$�óJ�y�}r��js�t�էi+�(4�Q`��1=�W9�z�һ{�
���.+cB��i�oe�;mt&v�:���1Mo{�'r+��� ll�sF:�4VJ|Е���Ww-���?��뙮<L�c�Wx����mך�7��tώkNzDlÈ(�7��]�8��>h�g�5mH�Z2c��o{=����Xқ�c�_]-;};� 9�k��O(Xn(��`t�^���Ls�;4�9�G��"D
�L��}����*ٮ��������mِJKW�俦��ʾk(�l��K5oS���ag����_&�rٍ.P8��US���mR�ppkǷ�E+��h���=�Ւ�p3����Av3A<���w�Q:8)����y������5geq��X���
�C�OQ�z5|e�s��ee�˭�H��C���H��v��k��:�ffNNQJ�7c�������j�����pV8H��䊕�$e�3��ؼ��c���+e7��o|�,5���,
���Թ@�*�Y��U��a�1�1����4�g2�k�V���n�� �f]U�v�.�6+{���S��.�f�t����&��O�"��l>�\v���o�V���_v���L���t�7���s������{:�������y�b�S�g
�X���.�R�!�18�m�)�2L�c��3�Ӹ������uT71��yӺ�Nk�'g;pcsJu�PT�����ݥ��0Ȳ�̋nk�6�2�*�u��pY�J�3T�%Nۙ�nZ�s��WvF�+4�Ӑ`��YT�͑�p�������CO[����ru2�<J�V�E9t��Z65f��k7]sҐRކ;��R�V[�̠jc(#.�Au��ͥ�ps�]Y��23A�0cn��X���\��e݃N�T�]��.顝�<�M�{������cYc��L�}]i�b��69�Vp���/HdV�˹���B��}7�B\��T��"���ǝ.R�{O�8pL�7���w���t�����շoqc�f1����B�<��ox�Y!���`��J�;p�Y)N��b���yq9�Oc*\��qJ�ۦܷǲ̣װ�JZ�ܗCo�D:Q-�]��e,0��&���b8k^�l�s��Ȣ�͙X{gr�zT��g8"א��>ç�W�U�W~|�,X���,�!�s�zƓ����8���]�����g�IƎ"m����,6Ī7n��\������T#�rr�GY�$����t�&)m4%�p�y��&�a�[ʹ�b���}���7�ݵ�a�ق�������X�����Ѽٯ��E�`C�N�zPg{E�)��a@���t0�ם���q��*\R�8;�Q꠯r�;;7�Z�/M�;�[ΏF�b��U�c睤�PBN�D�]�h�v��
o��]���#�r�V��9�}�#+fS��Wp}ћ)��=:�Qxf�dvf�A��k���˼�l��)"��В�k�v�@�a�1*|o3�[֝ba(Rq\[VJCq�vc�o]�T5�!;�6�[+yi�ȽD˷{s_oܝ��G/4nRئ/�!#��|B壚/��5���9{·����������	��-@��̾琍t�#j��x��$8.J�B�j��>�.���w&�����f\��MT{)���.�6��B��Y;$��rٗ1�*�k�nL�%}�p٠u��Gi��$��b��ʣW��NT��$��Rh̔57��܀W`^K�|*��HE�3�k�!BgM>�Z��Cs`�R���Ɋ��m�<J]��Z9o��yl�{�fG��m���I�%�e�9�*�,�Ĵ�G���gЄ�$�5d�&�7�0��:�l�z���ݢ#?W�dsv�����Ǐ�q�q�|qƸ�8�۷n߳���2C�R �G�%+�eם�d^zw�؝�v�w������8�8�>8�\q�v�۷n>���U��F@��$BL����,��Ȏ����@U���z�>����]�ytw��{n]g^e�v����e�����wbgdW�ғ�6诽�<���y��e��s�1{w���gy=i��Y�姛k"i�����:�����^�{��y�E�y��Zݪ�@�f0��|�<>���oE���œkmݽ��:K�S�ȷ��=���3�m�rm��5��}{���������#!<R��
��&? R�-"D2DYq�	HP��	p����\�D�J�wHL�_�kxt�8I��<�κ�m�I�i�}M�6���|�����*�E�W�H�|�t�����a�#����� f^>�10�AyD��P�1��e�� �	�1%c0�a�P(�3į0�00�1��p�a%�Q$�Y(�p�,Hl�癞L��) I�dq�My0�g����|�_/���E�Q`~PG�]N��U-x捍dU)K:�&b�Z����ڬ����Z_K�3����q�u� �0b:�o0U�+x�ӏ{��w^b]���%�,�ْ8��5�x���޳��(9���a�g��"`�������U�J�n<w���F���O��mU�QDK��F}yT��|�ī=���u���qj�k����ٽ5[�N�?�uq��ߞY#1V_�n�>�؍�W����X�a��E�e*{��@���G�>��8an��1�Ȁ���03�[�q�ɳ�5S(i��.*���;w쮛���S��Xey�?���Ȭ�?zD��+tF.���@��*y�˹I �:���d<d5����a�ͱ�1Чs��{�~O3*���w3���ɱ�
��>�
�k�N��1C�[��ϳQ�fVfG^����K���I���3�x������Y^�wn.�߾�ד��6,���sir4�Ig��q�f���r7���5�����s��ǚ��d����\�:��W3��,�����]�������qS<O2�긻/�����rG[�'h�����H]ïxW�w��������O/s���A�3�� ��rd=*���3IT	{B��<at��Q�S���ݝٴ�����Ѿ��K��̆T5�W(y�Nk}A��O��&1Nݸ��}w�B���=���'{2W����eB�Z�ܺU�s�N�M��l�g�S��oȞ��D�5f�ɣkhr̉�ݩk|*؅�yMXM�&��Μ�k�Y��2H�c+��=+�*3��>��;��%Q�鹍��ss���
 ��\�n�޿7��G��g����T�J�=����ߥv�@U���Rc�� �*n: �3"�[�=r�\�Qn�X�7�����ќ���-��<F+7��y4�^�Ľ `��s�sjw@�ʥ��/9���c��j��f��A�9ui�Y�\�ZU(���Z2:�#{��r���7�e��gg�i�{�`>y��t8r2�~�$��S���l�wۡj��HU�0�:�Υe��w��<��g��zS����&�^��fɽF�v{%�?��1c_˦��I��mj��B ���	Q>��c:]V�1�ɴ{me�~�z����隔ʵ1��h��)V�d�4LtE�
^�0�y�f,_q�����}�dwi� 0�~�gc�E���*���Z�޽�n\D1^kU��{y� w� ��cP�إ�4�w�]�ߞf[��s�|j����mtT�Рս^��4��Xa҆�45���޸ܚ��M����Y���R"k���ś��-��{if�k_X����uP���6˙�M9v�nr��4�BME?��WhC�Q}6�O���sfnlk�&�w�	��UX�ߡ��U\��G��Qg;n6(C�d��Mv�ӹ�#�6�q��1�*��ª��gO�t����mZ+�H�z]�ޫ��r���sg]n�W����aW�S~�[m�79S<��Ano-ד����=���,�ɣ؎�m��+����%O����^���k�N��3[�1��O������3���G��?�%J�ʌ�S���o@�'�w��pHj�]��d�p��E�N�?]�|S��(�.,�����x9��1V�ұ9p��,�
̴�H�8����}X.煰���Ǫ��;V6%v�&��~�|+���z���}iO�:��X�m���	e�����b�ﴸ��2�\������|s��r����m�-���W\��!q���W�����tW�5�,陮e�i�~�G��J֊�������9���)�rV��戻Zw:y�8� aܰ�C8��_�/�mØdo'��}I���'���UUYާ�#}xůT�fE�@uq/|��i�� Aq���sN�����&f��ӎ�-��20�Ԉ
�ܵ�[�܎��6D�G_f|�+�Sh��ޝ����|fY�X'ܺsү�1`�]3���{�{&,<wVHX[b��凧�jj�ͤ�l�gx���d��6jߢ%�$�-�ܗ��|�9�s�ey��ǻtv�W�T���a��x�h�f�L�^����T�N��&�8�9�J&�+V4�p�*i̊�[и�j]�K�פKZ*+���
��&�x�eYhQI�ѝ���K�V��ۑo)���������*�>R�/����C�m��}�"	0���r�Ф�Uڶ�Ɵ]�F[V��Q��e���V�.�Pɼ9�j$9`��ah�N�bx�w�;�̢}�
�|>]iH��y�!͵�Lls�P�ë����$|� T^��5�K33��өS�vZ�p�^�����x��G�7*1c��ǙO�';qgK	��|ʮC�x�'񕧛��)j�߳���;Q�X�5)�wy�c/�	 NdK�2����,^�v H���#cn��#�;7Z���zz׮�zu
3��n�8�Ϟ���pY:����2-p})�.I۫�{s�����&��'�t\����fX-�$��}ɨיT5s�s���B�'�W*�-�MٜU��9��!��]-ۙ�^un�<�ޔ�列Û��Y���%ܱ�+i�M�Z�2j:#9b�:�5�'ϸ�_�Dm=��U�n2{��߿e�z�s���ۛLҦ8w�?;�l��&���,�&��z������g�wzfX����۴����R��[���F��"�k��d<NO��g�cǐ`���dW9�K��E'�ݣge1�<�mʰ!zX{�,���TI�ҡ�J;gD"���y}�+ݵHU?Ðu^^՚玉c�v�z�ޙj=���(��\�#�����{�#���{u�3�����{�0~���7��7����g$�d|v�ț���z����3���z�j3e;I��ŝ��6��݌tg�|�$7r9����b{>7,/i��PVybg߱/v���øm�����.���kQ
o8-*����z�آކ�nF�|��6u�Ԫ}vbnf��A�f?���V�ף)�[MI��}��kN�E;���_Hzb^�]	�L�0Uw(q�fV�G1�ּۋ��4�8{#����;�3{n����}�T�G�v�.g���D�\h���D�_vG0��w�k��jw(�[@�~����Hb�M[v�f*}t*x��Oc޽��w]��ۚ���5����a�
�K���g|�N��#��k����E,��5{K��o	�C�ӗ����[�[W^Tu��{����c�5��%�6g���gH�
�-�
k��
����7�v悎\�L�L���2"k������$tl�o��|�Y�o��VԮ�!���8�7�{J����xu���Ɔ�=h��ς��0����Z��V��o���˲iR�^9���AS��S�{1G��Q�GF��0�F���k/�Sli]�no#�j�7o����x��������9>yt�h�l���x�3��邜��5rT��Iv�����V_����yo�$՞���`7g?�]���W�T��if���ا����畜U���o�mc0h�^��e�`��J��g`VK�Y�[��u�;��;9�|ga���{[�_'�m]2���3�K;8h�OM7�*�<7�f�ݧhA0^���gץ{���/��e���+.| _�H�k襾�9�9��&�r�i�n�6YQ���/yi�Ƭ!��� �jDM�T���@7�E��-@7�^N�n�Ӑu=ȼo'~��q`�����uX���Yk%�fX�pib������pn�yzg瓽�5���k,rت��!�sT��^�s��~�Zz�9����\Z���:[c�(��}+G���ϋCd;5Ӥސ���%7m��v�A��]��::x4鸻*��k�'򏻱�g�mj^�g.t�ﲪN����u	����f��!\=�l�Π�������%f[γh��x��|�����Nf�gn�)yG=�n�c�Q�\�M�j����n�׌�]�v���=��=gn���/�|��z5�����J��'�һ�Wqj�)�Dti�"�Uv㻳l.ۏ}ج��8�b���Xz@]��s��X�N�)'���m}�5�#g�S���}e'�Z3���<nL����Eej����ӛ[�a$گAO�R��dƭ�u옵�1�Hz��
��ݙ1�������%�PYX�3�X>e��n��v6����jF����7�׮vt��x�E�j�0����7�}�Cw5�H���=�km�0}w쩓��Z�^�OP��h�xwl�f���%!�?���goep��ū�@^^:��JfX\y��3�u˖���X�{����ׇ��q�����Vg�3�����v�{Ws�?���U6���M㇝�Be�_��{�V�>��?Y�_eI9ՙZԲJX`=]�2��$��ʡ�@l��E�uҗH���h��y5*?���Χ;y �dV��9-��W3x>R�j���y��[������W���$��P[��/Vu=�ֻ�UT��B�Cp$�(.[�.)�Br�j 1���i@s���ȼz�*}b���[�-ob�Wݸz�$߳��{t�xH�)��������ں}Њ��m���n��g���OQ�Ɓj�8��7��M�@i�a���f�T�&�2���o�I��:E�J�
�<��A<�)~���,Ӻ��Qu�}͓P�ϒV:��Ȇp�cb��MH:b����N��4]Y4������ՉC�u5]Ś��=���
��Ur�BJ=S�;\y�ҡ(�y�X���޲��3k�+��U���x�1��r�ѢR��m���r����~�K��N)������ɡ���/o�*<�-�8\<x��6^^����T�3�C.���͠�6�����s�A/ �l����!w@��Ť;V��-��pZ{���-����++��f���f�=+{�S�Wnxe=�O�x������F7���C8�{��{�ʺ�o���7);=㹠�G���Ev8V�)�,�����4bZ��+xww!��9� ��p}��b����	I�碆�׻96��jͼ6��!�����{NV���J�jc`R��9�ء%��\�h����t5]��}�4!��ˢdDjQo��lK(f2����$��ڬ��I��=��5|FU~�P�k`��g(��ᬕ����VRyU��-�Vc=��{jiZ���r �Y控�l0���Q���!����p[�L��w&��7-��&yv7��[H�ca�ㆠ�����ڪݷƃo�R��M���BQ}�#���>��X�5��zs;�^�����\�~N<P�`]���x�6�So��M��	�**���:�=k��[�<=Oz��^�3���W��+=B�`u&#L�<rAH%����<���뼎��o;R�MD~�w�M���Z���-]5s�K�ɂ���ź6�W܅�w����h��7����i�
mR�q�5�2(�a���wV�R�����e*�	��);V���)�ʓ���ʜ��]��w��b]L��-��n������T3�ocO��#�B�v��La1t�.>�r�e�ݽS��"^S���ˮ��Y���;MppaUÓ�J�K��ٴ$�ia�5ܚ�1hIh�}����!�������*��ռB�c�=�,�nǫY�c�k��P������:�)�/pH���v��]��i�m���0VDIKr���w�V����[i�-m,��~hH3��ؖK�u���\�u�4�N�ܗ�o-��_:��m��2oJ�w+��fv$�8�o4傯%��Ք@̩{ �t�(5	h���֎��[�祮xu��.�@���������j�=t!|�^&_�fSS'\d�$�u\Eދ"�T�L���A�v�]���-�]�ը��*5N��	�O�j;��˘�`)ᐎy���6��nT�G}�����ƚSyw�1���2�eQ�{gKl��u!��a�묡�^�F�-s�h�p'k;�{��X5u����Mư���"���tK{ή�.RB���R��a�TUӉ�Q��طuâ1W���k��	n�P!J�l-^P{Օu\�e�|��٘�{U[0?�����%)�]˔k:oN��źJW��iYŦ�KS[:����X�v�Kc`{8֋̪m��҄���&<����O	�0<�p��ݚ��|���j�0TJ+3�13�S�����N�:��� �]�=�D�N/:��\ܧ��LD��o�n��7������K�<��G�[�x�$��ίU<���1P�9؎���w_[��C:AYՎ��7u^u��d�O��W�ؒ�ģ5��p�f�	ͣ�k(�b�$��ĎpF�/
h��Ҏe�w
"����W<Ό�v!ឱ(m�K�C|^�b��0R0�kP^2�Ӷ+ɶ�۠1Ѳ-w1p6�w�{݄_LJk֜Ӈ&������.<����I�<��>��8H 9s	�	�v5��}M��B��c�th�eV��u�G{y����'AN�L��05��u6��M��#���0���j�o�޽t�{��G����@ޞ��1�J��r��w^4��R�|:�2��W�T�U��n�u:�0�2�2�u�?ruo�q;W�ֱks9AӶ�]_���gf+��/9֬�����ь�f�P�N�9��	�S"��!�F��ð���ٮ��fm�D�ތ2����s��.�HpfS&�yQ=���l%8k2������&:\��Y�]�b� ��.��م.�1���d���٪��y:�gR��A��ʟP�d͙N=�">�w�E�:wr��b�8�B�WWYH�Uy�H�	x���GS�	$��]�]�p7!&�M��$k�ooo�pq�q�q�q�q۷n������A��$δ	e����;-��s=�L�[S�m��Ǐ��8�8�<q�8�;v�۷GιY'-�2�d�+�H�^y�6i�n&���y;Ϟ��mYe�{�o;eC6[���G�~���}�Qߟn���zޣK"Z�[l.�6���<��lY��lYvf���Z�e+E�p�{d��k��66e��Z�������[n�3�����י���;n����y��!���>�'���כO}����|�zۛ�9��o��[�=���V�m�=ﶞݹֶ��ke�m���_l�by��}�Z֗%��>|�6͸���F��~z�y�Q��{=��;AnvvvbL�����H"~ ăH����}�5#��[K4��ʓ�#����&`��5
��F��{w�ŧ�)��Vz���TF��9ʹ_Q��<�lKx~��>>Y�T}�絺Z!��vh��W�f�삛��E[�[u���(�
%o�{:�;c�z�,mZ^ҘW��1�zWn���s؞�c�݁\�a�`N�������n��vl��id�|=H��R�З@�o��*R't��N]����;\Y7���]w4¹�xq\S�綎���SSx�0ѓf�3��[��zCk�a���t[x�O�0x��E%3�����˜�0���fѾ���ˢ�Y~z�������o;�rz����;�v�Lʮ��õ��Ó��q�<���G��M�|��b����t��bD��%�Ŵ��CYs���z���j��lI��/��:��w�M�'O���wp�0�!כ	�����Ӕ6|jGu��/�u��^�ü<���u�Y��!:��@&
FW����������m�0Y5�_���gTu�g�ˎ衱��5���Zʌ��]�H滫��
5��={���pE�۵�V��l�F.���
OE]��K<9��ػ�k����/P��j:F��5�z��*.�ο�>o7�{/�J������A�<���
у�M\n�׸]�w���]�����D���~�ؙ��a��S�{������}~˞C#�2g���7�����k�z2uVy�}������ *��ni�:6����
��p�z�v��}<֐T�<6a��.�nM6��X��K7���7.��Cwg�ș�ɲ���8g����0*���q#�fV׬�%U7frnۦ.D,��Ҟ{_�e�t�p�XdV�k%D��@�[J��c!k3O��ڞ���:5���d�[d]qi�wY��e�b��Օ��p��ٵ=�y�ً{���;	z��^rJ���^.��	�ʺ]^��VCt���ݞ�qw�`g�6}`�4��~���S�R���r�"��r�/��6x�0㚩"QwN;��r���Ƹ�6<}ƹ�rh��l��6��ϯ��w���>KG]��rR�ԏ� e^��� � ����1.��n�t��8|�e�ͼ�%;9����0�u�_kBeAu�#��$��ܝ��`��dMc_e�Bo".��5�VҖ��wq����>�Rr�2��;"�gj��>�-f�pn:�Rt�Xla��I�]�+o�X��|oH�ԝcN�6 |C�`i��2���k	x�f��5b��J�ވ��؊�%x�ZƘ�*΅�b_+;:�j��q��E�T��t��z�|��ë�։�ݞ7D��k;E�\&��ְ���<Ra���Fz�Wߌ�/�ʂ~ˬ���ؾ��d����?�S&\��u�k��h:���9����A�5���C"��ʑb�cS	��l����.�S��z(q��8۩�m��<��觴�E��1y�׷���Fc�w� ��6��o�9�v��ng�����J����Y�y��<�^7]oz��=2T�^Q{�*	\�iƁj��5���I�}���7��{I� 1�k��L'ܪ�{��I�J$��O�t۲��;�������ix�Z1���AU���$�V���;Ҿ��|E�|�]L��ٚH�m���cm�ɃXŨk2�c``�v�gM��W<aU�{��X��ڷ��Ë�9�NT��a�d恰&sl���Vt]NX=��+[W�a��P��f�x^L�;yMǵ[\5ӛ[:a��������Y���-U[�L�3:���RW/�ƕ/�dz����>U���1��w'��F�u�*��'�������T�>N�ߞ��;p����L�Ө|-M>�,�l�;��WUx7Jėo�uE��}ͲY0�U�t	��J�՛d�Q�c��K?G����3�z �Rgْ8��<�7������e;���p���»fU�-��� ����P��s+5G�Qґ��_'�E����7��t_O��3�T��C��U�m���i��D����?z7��n���o�e��8�K�����'�8.�J^i='f�O��;��;�o�E�+���|�ӑ�A�}��,#���g��Y�*.#VF�\w{Ӑd�Hȵ��pI2b���������7��4�a��2e�f���3��hmr>���lUw�5 [��,]m>�c��r�=���u�����U����]-�0+�l��Z�Cb�j�j��j�h�>	���~��c�NA�;��WA
�w��~���^�I;���f�f
|�k�Ṩ��F�b�S�+���-�w,,���ok<���/2m���9'R�>��J���w�������t�[W��V�����B��V̠��� �-駭x��Ncƿ�:2<���Ez��\���ÜrA@S�ں����s���=��9��Gu���Ϊ��V��w<c�.!b�SB1����{�:;��E$3�v�,����N���]ǘ�7Dϐ8�y;0]m9*�.8s������@;Wʶ�̪�X��x�+;�*�A"\�R�v�r���V�#�H�]��^$���d�F���u����Iѵ6�v�w<�oe]�#��N���#��sO�݉\�R��1^�s���'�/ϛ�ً��?��7��>�#����զ�u�-��vӣ~�<�����n��fzk(�A�����Srװ9�:㞸جLP;�ms	�ߦt^��e��3�0�'�,j�f������-�]#"zެ�	�B$�<[�x}�%M�n�[��&��h��,f��8a]@����V3uD�'�i$9�hL�ڈ��R��W�N�C��,����a/���ٙ|�z��Īs{Ul���=��V���[���M���2�c}� ϧ���Z^�qZ�n�^M��L��[�uטח7�Nm�|V�e>jesRl_v��<�����*��ٽ| ���O����r:��(+k��hw�[5c�[X��}�a�܎�R;�� ���q�ny��3�m.;��M�
y��8�+���9��d����,��9��=]];̪/��S�6S�+/�+6]���އ4X�pI�\����N�P�x���G�P��A�ܹ��{�)�Mu]a�%#�w.{;�_S�3�����t��&�,f=/^�k2�!���٪jw�W��Y퐖:sksoN��}��͠�D�3�St1b��ߡ���������}D�Μ��d��M�@VB���v��V��ꀳ���װY�Q@]�V����b�{�S�L<��ה��C,S�~��	e�Q�K�h�Ƀ����C`;�Q,��V¹��W�*%���J�������B����S&�e�T���w{�=�3z���4Q2�9w�E�f�f槽�zILV*E�f�M�Bl�&�t׵�1c����u�:��t��^�HJ>��kЩ��L����~�r��kG�]W1�^v�_Pth�WU�&JժT����V6єμB�u۔O�6�ݒ��d=ш継㑴1������;��=q9��S�yt�'6���<��r��q"�t��S
3"�*+O�}a^�Z�8c+in�� b�B��9>n�`��F������_dF��wDL훳���zX�%�rAww�ϯhpѹ,̳k�;�P}�-�<�����tU|�B�MJUeN�5n�ww��畘Z�{��T�����`z"�����ސZ�����N��bc��*�ǧ�mP������ڦ���l�=~�?6X_�9x}pn�B�	��kɻ:2,LJ�c�}��}��a���Ѻ�_����?����a�`z�3y�Y��oӸ���>�f�[��8^�ƻYn���Xf.<P��� 0h���ַr,��9���2u���r��-n�����w{w���;�O==Ntץ4Rr��t�� �fI�ơ�G�9}]ą=y�ˮ�q�yJ�kb���Z����������*
K5��h��Y�+c
U�f�}��r��\UX�]W[�����lt4�"N�w�K��vn���V\=�CS��{��/�̂h�]ݮ�_x����/��ei���sY��2�o�b�sx\i�h�Ndl��c)�����;�6l�a�="�6|�P{�(�T�&�;�P��
$1���\�V�f��͍��i��+6�33�� �@�mMV��;sP;�__���73F{n��f�dQ��w�TG,ʯ�w�`5P�[��O+��k˽�3�*��'�l�v���3�f/7j�X��`^��`[D�߲��c1@�T(�}���^�;�����O�حu�*���;��G��\~�O�������MB˹��w�7��3�<E�\���F���w���լ��)^��D�ݘ:$5jb�k�<r��цR��B�1A�V��^Ir����ϙ�p1�+IP����%넵x�z�i�s�z�6(�Y��ХG���E��g㹙Q���f�a�sIS��v����� �_�Ҧf���߾�u���s$�6x(�y� Hb��"����+l`�2��2ʕ����,P�lwk�Z �κ�b��=���U�V!I��0�f����^έ�+�.d*G�{��핛��-�Ӻ��,��1'0�w�l�mg�_I�b�]53�Uҹ��n�/�||}Sm�e�݆���E-����-P;א��y��R"}�hd��Nj���Tѽ�:yKydr8w�]����cz������݉��b.t �\�����U{���ҽ�@��>��~R=�b�G=27=.�|���˞��2�S�u>�Q��n�Y�}��{��=�w�S�X�~�ʢ9(y��U��o^�i�x��v��#�ס&z�G��&=��#x,0��Z��]���!�v^�^��5*�"�<\�����_�s�gZ�`74�M�g�@s:�;@�>�1n��o�D}�����=�[_���T`��QC?^E�Ol�woHY��PJ�(����wx�ˤ5��jtH��ҝ���e��u�m��l`��ː�Q�ױ,�RMYU�
̢�V-�/\�0��+�o:n�1�9�Nڥ�𑰗.7��e7��L�����RĐ�۶s�웚Fw�pߝb�/1 U��S�Іڥ����O���T�=T�h��H5�s�P~���q�ݽ�;z\Qi݁�1h�4�dl`���Y�/Q�����`t��9���G��O������&��7 �Q�vşd@W��܈�Y���fh�F���n����B7q��oV��K\�=u�V��W7�B�;9E�.bt�������wN7ywb��#��py�}sO>���ʪ�ؤ�'#8�U<���ik��^d���2�́BZ�߿1���@e{!K{yܣ�؃왖W;�6r�?/VE�C�?5�z�����5�ъ�=���z�dв��k��Uod,}03
��7�9�|g`q��������-��y��V��f�����}�) T���ٲ*�|�Ε��ۍ?��z�m�~ඣ)���~�-�8l\�gv�(_�\(���@��	W�WG�tg^N�ˆ�]t����i��p��;\�k����t8,�²�|�=Sp�"���+wF�e�κ����Ehl1��t<8��\]��w�Ͽ����J ��
"#������2�������)�
�C��wv*-$�$��`�(`,�b��(`���*�� A��b�(`��"� A� A��b*���`�B `��A� A��` `�*� A��`�(b��
����
� A��*��� b��*��
���
�� A��`� A A��b��A��b��*����`� A��`�*��+(b�
�� `�*���b `�*��}t;ځ
�� A��b��
`� A�`� b��*���A��B
�Q��`!
���`�*���*�� b `�*���b�
���B b�*���b
���*���+ `
���A��b�5��B b� A��b� A� A��`!  `��(b�
���b�
��F�@`(&���EP��UTP��UEP���D�
D ��@P ޴!�1P @ 0P @ 1U �@�E@�1E-F���"�!@b ��A�`��� �A�"!��a kZ�
,
0��b�A���� ��@`!A����@ 1�ZU��B   1Fw� � ��`1V`1V`0@��XU���� A��b��*�����������}�"�� ��b ��ˁ}���<�?�~'>���?����������g�����0���Ԗ�����n���?r ����?�����^�� U�����@��	���������?� ��)�~������A���'����������?D������"��@�AYT$UdQP�PP! $ �@10@P � "A��� "0
� �  � @ 	 "  ) "$@ ��A �$ �,D �$ � � �DH� #`$U��(@!`�V  �X�@�c��BQ��o����� �"2 �$�  �H(�?�?�����G�������?3���� t�����o����?���Βp7���G��t~�� p??j~_~���
� _���D?����4� ����u�DPW �T�_�(����a;
?�/ۤ���?���6�@Y�?y���?R���� ����?Q�?�ó�j����7��?�A�_���$ p��R�_� @v9�8�a"U���?X��P�����A� ���D��� *���||>�P?xl����8������_�z`P�u����o�n���0�}����e5�`�WP�e� ?�s2}p$M���,�lj�R*�J�مm��
�+mA��J�)$�bZղ�j�T-`�j� J�!J�Z$KVdĕֳ5E+i,�5Q���5SEj���U�Ӎ[Y�m�d��mFݳ�m�k-QlI��lca�SY�5:�s)�YlƖ4�[h֥�KU����Cv�ڵ(�jٶ���lfZ�m��[UZ�P�m��`Smj��e�4�+e�V����
��5�&śM���5M�imV���l�5�LU��i��   &q���6ͭ�(��;��kkt]�sA��`ij�j����)�jSY���%���í���Ul�ZM�m�[V��Xs[WQ�n�v�]���Z�[m�ֺ�kb�S[o   BB��D�
�=�(�(�B�
3ޜ<�
$(P�B���l(iiv�]�lh��Ӯқm�TM0b4[*ev�5vuu�Z]�qւ�պm�S�h"����f�5��Y��$��^   ү(�����r��-mX�36���l��( ]fv�.b�Cl`3TZ��S,kjP�5��w0٩E�L���j���\Y����%I�Sj�V��Y-Um��   p�h$V�cU6�z�U�MܻB�(f:�%T`j���h� ���v5	7p��Ҋ�Ua�Ts����6YI�fͫS-���   ��)���$�f+ 
�*��n�4��wrpҌ���4;1M��U�@�j�l�ӶTBl������]tu-�+�  �=M!j�(��N@q])��Օ[n�t3�h(��ՊTUE�w Pݚ�UT
B�ѷXrHAKvHkSL��)�d�U�Ƶ[<  ׀ �U�� �  r;���:�  Yu� g\�P�.E` �����N�:�I�cM�F�l��ե6�#x  x
 ��uP (Mt  �S  Xu�  �8
 �0  6��h�nn  6 ���֦��5��2mf�56�  �  �  zg �F�  n�q�� ������  ��n  �i� ۻ� ��f4��kfFZ��ēM�  �@ �` ��0  �5�p iۇB�7-� Uv��@ Zs��
�k��ݵ� � E? 2��  h��$��#5 5O����J��   E?� � ɉ�LL� �*D'�T  j?����G���g�dC$���_���Z7�s֟C��+���-JڱC����������K���͌co�  6���6��61�m����1�L  m�?��?������VO�"��Ln�Q�҅� ���C.R�½2f�j�yB1"cul��^M�����ށ<Ŭ��0�<�k䵲k �/]8�E3I;��2]+ܠ33h�PU�'*#1]��9�C�V�I�o1���e�E�+ڙZ��� n��sZ�#��ʅ&(���T)eՋ������e㭆^+m
v3fƪ��^F�^ ��pű�D�0&��Z�W>ynN�����*�5wc����RF�d�@�,�sj�>@��&:l�TS���5��x�c�A�3�zM��V�z��IgK�28�Sf[Я-ݵ�lC�1-�Xh-�ϱ��"�VDQ�p�eUGu�r���W��Q���ۙ�@-^IW@��A���{���Vm�ț+Pwt*�f��˴U:)f���-e�,��-{Q��=��D�!�1O�eyJyR�l�"VN8&K[�l�yN��[���X�����v��[�1���.�-x D%���4��f"�m�pLm��9��!aԯ4eY2ܺ�M�4r��X9t\�y���[�. K�h]6��D���Ȃ��l2[{��F�$�rZ30U�����aƩ6�MŎ����ͬ03J�1��w��8�W?�r�-��5�c/K�Ņ��!Gz�������p@���,Oo�5#E^����3n�����敔"���Q�0�^��x"NP������F�U啶@���r�3W�b��2�iKP��$�k�4V�j�.�T���R͕^�B���+\Rt�R�W�.��tu��44l��@��cڰ+U^��&���1�g/h��m�"0Ȣ!bi��[Q�)w��n�7ë�.�\{��FeX��tda��/L^�Fŧ^� 1�O��ZRڬ'.�)*���IS"i�	2���˸�P�ިo[�݌���B ���лۛH#4�H�{��an��tʹD��m��[��k/#wu��a���v�⽑1�b�,��>�p�� ["�&�AyC3N�-�X$�j�3�@�"�A�h��G�V���
�V�����n��>�V�ouJ��M}�։��ђ�nn��e�Mf ��ݽ�t�wM����0��̭r=�Q1MECPی��U��ʸ]�b͗��Z�-hFh������W��3(��b�S)b,����N��Z�;��B�1"����De�cLu4 ڽJ�JW���Z���rH��Y�.��JH�J��6̳���nc�/N��n���wN�^Rf�c��-���V��KɤL�� nC.c�r�EcE��ً"yN��<��[�;��H���0��3k"�n5V�N��u�i(�( �Z��$����(zt᝙�'��C�q�4�'paN�1f�f��(�)�J���c��Y-SNI"�-�S/E-�h.�Dތ���J�ǆ;��d��nS��U�ѬKU=N�n�́-*��лت�l�����l�f�-����U�pѧ���±��ƭ��Ne���[�sX�1e�x����љ5�^j�Ԙ�V��dm�tq��Ơj{g{��R&�嬜�U���=��������`J�*X���섷l"���.-�S��܍�q��6�e3	�c�M�Q�D�%:���Q��ܚ@;����-	�EŸ��2��X(7i:�	Z�%�.�+ǲ�r�2���V��,PBɸ��MtJU#/6�e8r�.��u�_�˲�M�Xa�qn�Q��%�ua��@�`���n�1]����ĝ��u�>+i&5��7��C)�r̗��q��]�X.�7L�*4r�X�B��-6��q˸���=��ֳ�����Kߙ̩�'��������|W�6qF�۬��"A������#p�JʃI�+fK�/fYJ�ܠ�I�@��P�:�pX�N��b�,�ǶƦw��M����^
��k���4Vds)^��<�]��2�U��B��j���nYӉ�?n�H�,݋b�
q�{Z�%S�l^�����=�:y�n^"^�t��Лv��Ô�m��L�+	
U��7{ M�������^S�n�Z��'�0�{�E��FɠQ
9�6��@*b&�mf���Nզ��E:{�ʡ��D���A���"�]���sn�1�����&�ɲ1��˥NQ[&�4���UTIR,�gF�̑�CkZl��&CX����`
Iiһ\EhI�|�!�MU��2i�m��>�"���)A�^ٱH]Ah33]h�V ��w�KNE��wt����Xڶ�nQL�J��#*㐁G�x��)��np)q1?֧t�-Xt=
D���@'��ts/!pJ�bZ5���0^e�t������;���O��o�u{�j��[&Ǜ�%�m
2�C���YWb�LT���MQ�*�YJ�{���cm
��7DM�a���7�ے����y�J�rȚ�UփfPq%W��#WB� *�n�h26-�_
J��F����ȗM&��75����gM���YI�b���9��S
4-2�ju0ȭ:��ҒWRi���*"%��%��P�/Nlj
k�-�է)���W�Rr�����;�i�9�;t�3�B�6��Kʞ%��l�����4�b���3ss2�ʍ�D��;�1v�o����h���7t$�����۰P��d�A��=
��g�p>� ��g��1��[���/`0ax��鰎Y&g�	�2���Lsj�:�ӇL�����f��Hp�LK,�ӹRLy����$P0�l3��9n�)ZZ�;*eF1;���dJ�mTH�M2�0]F���N*�il�L��Y�L9!��^���h�s2���W������^e"��C~ eo�4_ʁ�!���hT�Z�ڛE�V+V`� ѷ��U�z��T�V-�ږvEX�3 Sl�ppJ�+J�R�
nK�
�0U7[
=�V�4N6m$򅼿��p�q���q83@#`ԳB;
y!v��0�!��Gb��owS���v�.���GFV�8�MP��Xh� �I��膶�;����NiT6a�N�L�`Tg4C�Nj��i�2`���{���{X$zؖ���aV�Nݟ��pGt+%�m	g�*Q�M90�nt�Ì	vJŸLOE����M�L�^��۸r6A%dw�� ��ֺ��ٖí���l�d�#ẩ!���a{��;���r�u�iH��B�`�+�k�%�v�1�N�=Cqi��'oqn�18�fk`��Rx�lJ#�a�d$��j��Y8�t$����C)e8	��˛wm�L��a�t�U�Ȗ(��ȁn����jkN��<��桉�)>�"�Zh��$Z��rE�Se�h����G2��Qj��YpF���ۄ�'& p�=�1`�(�Z�:�q���#�w8v�n+ 4ÃD�ą�0���!(f9h9�`�5���j��ٙ���E̗Y �`�@�����e����[++im=H������͂A$>#}�|��'NRXw]�z��L:�SPG*ݒY���V�,u��>إ�K`���U�`�D���oٳ�E�k���i��Ƕ�9�^���E^�jI��0"G�8^!>��wBf���5�Ĝ�u�X�Sl� fi�r�0AOA\�]�Q5��lP�����j��A����d�{Sy��n���E��b8�M@�*��P��;P]�'0�&�L�3(���6�� ���	���7���q�1�� ��sr��v�H�p�cR�BĶ��F�k��%��PBh66�R�;ص�2���B��]5�0Mn�W���a���&��TUah�P�1 �-A�"/��f�mɅ�o+p\Xm�X�5Y�j!I��%��vj��Tj'sr��B�	X>�lT�rVT66��G@"9F�#*»,��Pa�[@�
�ug"�HA_�J@Ev�5%"�!w�ެ��)<j���%�
¶ͳ�2��)llj��(������5Lʠ��U�m7^lil��0^�' av='SԲƝ��l��'[�I�Y�\[�O�(q�����Y������HM[��g�5����Mf��Մ�e�f^�w��&kQ�3(^:�R�L`gVU�XI@X�Tؔ�;���1��eL�V�+#&�t4n�;�i9-�KMn[�%,�Y�s,��R��dZ�����NU�J#[b��1J�Q�O]1У7b���t�3&6�r)O#Ɇ	Q��ȣ��V�^�гl��\y��K��d�m=�q�+6�'��#�j���m�}r򒺕0ݶ]����.ޥYz�[H�$Cˠ��}�f���^[P�şn���A�&�*�E��v���5v~Bh0�nyk洦u��̘����j��q2�>gV��u��]�9��D^n]��T@�er�ěM���,#tV�Z½˷��y#�a�j��j`1m*�`� {	��FS� w��]E�K(���n�\�]�V�-̒,�N�Y�4�l�j���y[X�ꬩ{*9zN�"��M���\���.J���Z�q��(F8!E�z���	^��Д�wa{A�fc�n�r�!Ӆ�0�����{�a���©������V�^�F��,�ɭ�Ǜ3�h0�u[Yr��F���^��,K%�e�m'�%���S3m޲�[U�J+ud�N4T;��y�웽f&ֶ��݌��J��+��	�i,Ӈwǹ�I���m�&1�)E�Yj��� ��Osr�Ы	����]�;��3J�S)�G �tw�[ �n FbQmk1Z��"�EU�,���(5X����1|>N��OtKCk&��[���F`��;R,?��(V@e����[p���e�D^�m��`Ԉr��ڌ�J��k�u�.ӕ'��ߙ4еu/6�
�w�b��
ͨ��)5t�zKF�۩�'�V�[+e�JAB�b���FiEAT8����YAٽy�x)Y3
 �[�t�u�F�bo5(�c 6�l�ݻ�)-ڲ��9��2�����J����c{n�Kp�ma��X!��7�L�{3n�Oh��#�L�6*�7V�3(�/]������kbP�X�D�R�2�5Y{anR0ͣ1��iFB�:tE��`��`�ʔa��i|�ڄ�x��6��C�ݼU1m�V���͂Tz(��� ���<R,u添&�ܱ��@&�$����s!�ܡd��$eJ�[@X/U��[�����kR�%��ئ���#r���� �x,#R�qʙ�vQ��WZٻ��K-�j�3a8)�kK�MڔE8���XFj���^��Y�Et2[�_��&�ϴ�4c��A�	��Ѧ�`�5�p�JЬ�y��O��A���4`����H����3.nf���`6ۨV�6,���l4�M��ָ���iL���QSH�31�[YUh����]^���`��鶪e�	���nҖEX�G��f��Q�ܭi��sEC0m�0Qh<��e�x&�-G��M����n���% �=82�p]Q�҆���EZ�Q
��]��9�V�R�F�X�Y����=�-���^�ڒixf�A�L��T��Em�
N�%#X�DO,�5�PU���QG2%�kXJ1K
*�y�Z��,��I�
 h�s^3DF�Ҋo0�#�pI��7|�)�<"[�q��Zj�l�V.U�x��P�ע�ݲ���K�co[ܘ��	�xښ5،<܏�)A�+v��eK��/��ޣ�/��+#{F���C2?l5��3o-#���6�CV�*�)#t[P�P���k���t�C]K��
e-ͼ�r��G+V�ͅ�.��q��|B��n73��f�:��z�յ0�A�0%R�t�X�t
;��,tf�nF�aFS7��Elߜrm�n�K�I�z�+�˴&ѡEȒu����B�J��C��-��^�n�Iot��wr�w*:y@2m���X��0����9�(t�0��MC-�N)KYm�B�6��-��i	/)5h��j,�DN?����E��A5.?�k#LY-VA��O[�v+.�����q�v�*i!i�>7�	OC���:L�B̳0�JƻI݆mFh j'�&���F��r#�A�7[cpH+FR�Tު��|텵����.�Y�&n2CqV���4L1Pu�C�l�V�����@�[71�2��f���Xci٨�B����-^���YM��x���3[�C[{k0a�ŭM�tsw�LYk ��ֹ>��DȠ<��ow&���+nW��4僊��N0���<�̥aTɫm��6�����)Evc8*�Z�<l��4��_=�ե���<v3�pɸή�c%�Q��6c��V]66"rV�cm�:*��&Z�\-l�;v�0�26�D��c�QZ��(0��U*���Q|4�sN�C��#O�!VJN���)e9I%/1^E P0N��T��ېZ#o+qY�j���M�/]
�R�2�W$�բ���E�c/\g43o�vh䫗OV�9���v
dM�U�(���q�b�����k�R,;�t�]�1�90�FpTv�-qU�F���h�E5Kf'l�Qi
�[m깒��4%X��6*��Vk*�h#B:��Զ#`�:�5C�HEv��Fb�x�.d�۳u�ٓMh�M��:TSd���dͧwN�YCmK��ɱ��$��2�6��v�2V)��h��\��[�#��n餚�8M��'�pȳ�ɑ>d��#��5^�&��b������K"�ґ��髳*�
�-�w�˸^|!q�~�̰ͫ��d�QJYY>�Xg���zL����~tUn��E�ZmLs��������jK	�#��n��n��5�q�V��s�'�iݣ�H񅹜�oNL���+n�+�ɋ��va�'\���d8�Z蓁���w�����m.���Q0�v�i�v��1�h�O��i����t��o+�V�RQ���7l�[.l���r�$��ٝ�79H�N,Q��E7��(�qE��q*��}*�Y�Ӓ�Ї�4�D!x�	;&�ԴeHF\OOw1:�ʴ��e;�jP����ڡ@,��d�kP���5f������,8"uWf�K�G%�B�V�� EC�p]�b��8���黲�Q��'��q�CG�k�8�΅IKŻ��%�SZٓJ���,�}��p�IY|%EӔ)��@tys�ݜR���C����e9k���rmci\(hk4fvg|�� ��\�ɋ�0�}��N����:3��TN�E�^��lM��_[�e�v"ei��2	�i�TZ�Hѣq�D��wc�鎂cx��C\�.�k��PV�k���N��U�����)�z	f�>:wm*`Ƚ�˴�R�Fg���Fѹ�4Ч��޷�M�Чa�`��{�ڭս���ٵr%y�^A����|���p���&�ca<m�w/����o~����`%	G|��[��-�a�$e���� f�r��rT�p����| �۹q����fl;H�.�X:f@�;�y��)*۹ە/.�iKI�y�zGwN�ۡ�;Yב`���*��о��b�	���l+=�]���6�'X�`��,�6^e��T�J]��1VoK���c�=�|��M
�3Z[ƺ5&��K2����*�밠s�c�U�h�� 2�뛰N��de��tҵ�DK+�H>o�M��VP����0�1=��^��.��ޏ�/vPU��vT̡
$�|ٲ'��`f�J������q�(�Fn�:O���puh�͗�����8��p�/��y�SϬ9i�C��zqU�޴է\�͠E���Py[9���}w�w/�b�b�4���[]ǵ�FAnmg�X�T��$�O8=�&�EP�#��6�t�7;{�\Ga���i����jX�A��*�l�^Y{(�8�N{ K�t\5�j�]}WC7.ւ�9����E��ͷ%5�Aի��m$\'Z�IiL8���7Wk{�;�DQs�!p�)��>L��[?`�
=k7��Qٯ�_=u����΄��1�4���<�S��*}\f>�'zƴz��D�9�ri3{9i��ݢ�;��G��v��Wb�+.����t�:�$:��_i8]��kMCِk.z�d��u[A�¡�ێ춮�T��o:�q(��Mwi5E�5i����zT$�V�Z���U�\?H����,��>c��"��g�֕�M3��8�G��L�����V"�	;J���i��k2�ck%��5R��6�nq|@X��G�h�b���F@�,�s�$;'ږ�AP�P�U�i�d+���Yǹ:�}��6�༺���,E�K���8A��41˽邮�$���x�@��×`�kf}��D�-����>[T�Bx�n^ Ȕ^�����v�J��dۊl�b6�x+e`����^�[=Q��m*��b;齺���L0��iQɯ
�E�!�y��s�$������1��l����+ck�o�T�����Ù��n�@j�u�_;+�BkB<��E��u�	E�UY��l���j�����c2����g�^���ܼ���=Zj�#ZQV����5z�}w>=}v'��1�}�;����9�v)'qn��&�mWI�s�X�r�06޿�>t�Y��J�S�b����f%��f�c�%����ȭ�����k��|�����i��1�Ny�1�jﻅ|�����\����Ӄ��k��Z�q%7vqC!�#&�k
ٳq���2�ݛ��Tx���Oxڮ���,��g��5��s�]}F���	܊E}�j<-*9��xB=�08b�59RĘ�j<<w�-��oif��W.�8� vOgk��噷/q���Y)[�jʣN�Ŋ+1�V�=/U�zm[|zN��2�A��̕ӹ�r�� 5̦u�s��fkjJ�]�+ZP���	�Nէ-���F���N�>��1˰�Ĩ1[��}�bZ�]Ǭ_���)<�Ʊm�G��o��˚c�Ts3#Y��5%�u@�e�6ɇ�P�w�t�����Yu�^-�~��Ŏ�VvgD§��f�#t5雀�������x��_0P�6��컝�Іk�ܪ���*�H�8��J�㖉i8�3ƅ��Y���d����zt�q�<��)�):H��o_a}�����ۣ��H�����ȍ;W�׻�!R��
)�b�E>�#d���ۺ���9�b�[5գ��Y��o��	�8ã�
�����SPЉ
���fT�j>ǚ�gI �m������|��B������s�����H
3��Y��2�Z8��uf���:_S�w�$�b९{w#�;��ۇ��E)��vT��i�(
[����1L���94�����ѝ������Y�sS��Z�K��T�`ltκ�DZ�ᨾ�w4��u~"�0#�t�ё��W"
P�Og^,��k[��6hK[��rW;哕<3��ow�D��"�jw�^��}��O�O�����$�n���P��D�>t�����s+��M��-q��s����;�hH�������ޅm�_FM�)�U�C��a'f�*Zrut ����y;-���Q�f�0rK�X4��e�����Z5��α��rޱ�`�lQ芋� ����Yn���8hS-os%b��]q
Z}�*.bsǻ�ˠ�D��nCo<�՝�KV�������Ѳ�0w3r�J����T��k�rǲ���v��u��]��F}&�υ�DU�����]3Q��K�t�L3�i�W��c��g�W��v�Ӛ�[�6�
��-P����d���͢���Vl�1���5������F5.�;(H��j�f9�衒�Z���F���	0�mY�+��R��l�X�}���H(�b���R���}�V:0����l^��6��*ĩF���:p=�pq{YLԢ�D���5L#��#��9�Z�8���[�j;˳��\q`�dn b��q=�GX���K���&m�l����sr�I���	�ՁT.-�dʅ*�3m=�s��;�
0�; ��T嗰��.%��P�X/-�'F�Sj;�WX2E5b�M�l��m�h9�g%4YG	��zj~�b��&���N�L��g�~c��Qgh��::��{��ke�/�X��av�6ކn�0���0�l����{2os�Ī�p����%���|\]��zP�v�)��l:�Z��1\|�Ð�4l<�3����w���L�7��uq�ok��!�X����|,X�/xt�I짭���)��qv,�`��n#���U��su�=gӌ;8�N��`S�ep"ޚ[l*��ӵ,"a���u{��=Y�.��:�����7j/fY:�QNۃ���7�\Ƥ����঄h|G�5Ex�#�xt<�x�`"of|�=J�hA��A��XU6ʱ���pI�F��%ٯ�ʽ��Uxc�q��ʽ��d��Koܥ���ńA��+�7L�u�������8�h�̱���ח;�$�\ڬ 1�V�/�νȄA�l�䜥����zu��v�6��վ8�����ܾ�0b �n�o>�Pq��z6wv��9r�.��]������[iV���X/a�S9���f�crC��,Vg�`(ޔ;��K��t�oõ�0�40ܨ����n Dw�x~q�s�%j�, a� ����W.�M����y�7�.�3w�ı�������V���ie��}�[w+=HǴ��1o}i-g9��-��hj� �x'�Sm�ֻ4c8^��m�s'E'8t(w���x�űB|Gc�ZC�Y��2�1���GPep��+� 	�f��A$�[�lB���{�w[n�����&�JJ�x�qj2o:;-�T}}����i!�N��<��f���ee�Sj]rj�'vI�ڳ�r��Ņ�r��^���ڝ��B7qݛ�F�t�����.x�,>}e%�83؉���10�ի�S��оy�r:�k�oak�-ޔճR���ڷ���p�*-�3ˬ-��A���N�b��;��r�Bn|���)A�����g��~�5kW������D!!��Ft��9�{y{;@�ܷ��-p��͛j����v�WX*=�y��JF��D���f��0]�������򄹶�V�U���8"%��9%n�e͟R����R)���f��g�U)>��8<�z��V`뫔��`[�.�uݙq&�a��p	�:�͇��ǻ����MYt�Km�,l��\z�d@��]p1��k�OVg:@`�a��-��	wm�
7Q�R�k�vF���t_V�jŜ��-8�\����Z��u�A_d�d-3��8osZ�w>�s-���,�`�KwN�̍<�-u�u��k���;��Kw��K�Z���Dl���4ɽB���6��u�1�	n�V�ʀ�Зi6����g��w�ɇ�OSf��1�s������`�ۭ$�@�����yXx?��Z�Ҝr=����H��o�e�=��4t�E��zcY(�}���:`ȍ4����I��؏b�ns�o����=��.W�'���Uz�Я�Փ���T��ڶ%����0��KD�t�\�zLoQ\�{�V�Yъ0��VS��fڻ�*Y��4����7�JmZ�oD57xrq,?akvgr;��*[��8�i��o$
�VsG�*��g��Ы��[�iZf��}��g��|�!�Vmㅾ���Y�gd��,29�鑃�u:��M�f��������Rh�v+e�3��'���S5C�҃�#����,pff8��a�J��g�n�۽{��M��\�ݧ9�Չl�cA��VP-p��QC����#,^b���u���9Ưb-:4����5oqqԞ
����z9���Щ�<� �IQ	\����-(��3�X$=�o��3P�b,��CU^�Xg���&�f2�B+�R9��P)�v�ڤfP��4�W|&���;y�K#%r��k�*��rM��ץ�%��v���%ڭ�Zl��m��6�4?)nD�yg��N9I�]��i�y9c���n�d�WN��s���i�R�k^�0�T�tc�;�9ׅSt�
�<����s:y��i{j:G\����4k�5�o��A�8��^����f�Bz�!�Q�5O>�7<z���7@�ZʼC6İ�[���0�2��L͗�#����DΡz�̶jy���w��9gh��]�'�����{�_�-��E �Z�t�B��bz*�lն:�gA�c3��,�o�َ1��Ƒ��"�j�^.L���U`�@�X]��^<S"���i���|7�<RּV��KI��˸z"�g�m#n+�L�3F��h�T�����{��w�#v���9A�<�֎9'4�(�o�2�a�}1�e܁��nn�I�����Ԅ�b�]2�n��}Bf��7�}-f��'��k�z��Fu�O��kW�<�G�p���Om�P۾�O;7��'�q/B�u�}���[�>�1��9R�jj:lC���<Ù�wwm�{aֺy�:�-���a��5>u��ar��ڞ�]#X�_i�<��JM��G�[�^D�!��i֛��|�U̔�|�<|�4�����.��<Zn�IܮW�����<�徖�>IP���w��q�-ͅբ���o3dNk����N�=���=�eLR� u+:9>���,�˩��b۳Fqn�E�X����U�]m��X�Ts7	Cܘ~��*e�j��7g�N���k
������f��eS�8Vm�fwa(�,�/(-W]]{�8��մS[Sz��Y����{%�秔ӻ�����8�)ږ:��;���U7����Iwهzwla��i9^�އ�/�c9�/P��r�J;S�)k�9���YAk��G3x��GrRf�C�7��vo%�?h9���x�ۻWb��P���B��[����D�εlN�V&	ء�b+4p��#Xj2�'0A��©Ws�.�u[3 �l�����!w�($D�
�j��߼{���	��r�W�kJ�p�xg���q�9}K�ʙu*�ӗRw�ƳD#����̾9y��3�`m�������q�F9�׳6�4�ԖGdp�{ݚ�^ȼ�o��|NzE�o�S�B��#4f�5�GkDut��E�R�[T_j�s�*�{[|�WL��0V��_/t=�3�j��u�Y��U�و�{�����1u���2���!an띶�v�Ffc�w��95��UU��C�e�:���ݫ�n�5֯q�Ǆ#�륗�M�������z�����P���^R���[3�H7;m(3R"9�]� ܝ4y��V>����ӛǊwrI�V\ݻ�8�{[Վ���-���&��kB���f��t�^?���"$��x��'�D���3�f�[�-(��fZ�#�ުx�u���2����WG�l"������v�L:M���j�r*e˛�����N�	�++.�kw��{����Qi��ƺ��Z_Go{A��f��	TNd��kr��P.���۽�Μ^P��Ȧ�}t��sح�:�?G������<I�0kљ�v�t�rT�Z��Gop=�K��9lW���L.Y�>��rQn���Nw��z������u�����  ��m�`6��^[r��@���@��kLKb���R�{?S�o���;VJ���7�/J��w�
jA�H������@I��SCr�a�z{+�s.���$�/,=���h��I�@��X��T��tHīd�AP5�˪3����FԽ�	u�Zp�%�ڇyN��Ñ�N�q�ɷ|�X�eq������4��ōv�:oE�Ӻ����W`Ĉ�DʘK̜�$�<���������js �69H��R�]�wg	�٥�I{w.�m;��SG_WP��,»Z��}��Un;�m<̕����A�+uP,%&�,�ٯ�*�b��zZ!��M�*c��J�|O7G�O[�xvꬥIg�TS��h����w�������^@�v4��YC�'�ʅ�r�;�v�:�՘N�
��91�� ] ht��H�v_ҡG4��d����S��+���򚽹�]�uϘ�գj���[o$������\�����ͳ�P���p��C٣�9���v|ZQ��U\��(����Q�D��d�i^�	�����	{rѠ�۬�f-�C���?eH0q=J�֞k9�Y(�3��XM���>�o���8��!6.�^Q�u�;׫���W3l�I��P:��:�j�(A5���l�+�1��6�u�ɥ�p=��u�+d'O	�v����1�x�Rӝ��D�><So��}*���mQ��Դ�GnT�a�}�hO�]Ù�Gq�F�Q���v�������!\y���u���ۜ�W�P���&c��x��$�G�u��7N2ੈ@���C�+zӖ��x�>E'���Y�I;zmg�7��%��;�u�ˤ2�4��$�v:��X����;�PB��[,�Qs{PJ�b��&�p籋1Ӗ'BG_=��:T�;�C�tc�A�}�P_�o1�v}�+3����TW�����[ە�S�2B����'oy�nT���I�B)_��_q�-�wC7�挾��m�p>�ӻh ��h�tm\��A�[h&ur�e ��8��j���O�U�*�&��V���S@@�v -[�Ǒ�[�l6��pԴŦ���3��J����9��+w2�O<��6���уg�
&�4������"��9Z>�]w�j�ǥ�@bX9�����d�BU�z��@��h�&���� �n����U��<q,H�VF�����(*n4*�g�P;�����	��)M��q �u�T��P�e뿡�b#CY�4�d7"ۡ�F�qݒ)��t;�hX\@��7��[�.��5���|�V��-��!Ĳ����E�5y!o6/��;;*�,�Mr���캏����רf�z�"j�U�w]m����ڧ`��{v�Ȥj�Չ�ܖ����56�dHaln�@�%�=��n�8�"t&^-y�
��0��N[��r�pA
�HPԺ���:P�JR�:b���v�9R�@�bU��$в2�|�6��p'��������o
C͵�u�Z��T�t�"(�6h��b�3{�T$Ѯ�ʒ��X%���k�h�#�z��Y���{Ws �{�Q8Qt)�3D���G���6�}����C
�p[�'���nz�_'ܰBF�qh���6�cLܼ��gǌ���n���;0K��į8��Ss:��j��6����(��ӚCU+���,枫-oa:,�v䌧�����b�@�v�!s��xhq��e��L���F�ˡ�И�DD7P#:)9m����&�p��:�e[||6��<pp�ˣ�)����6�=σ�!(@�zX� :h�����W�
��7N-��[�&v{��OU�R�+�{�pd-�Ӵx�BKT*��g�LJg�:��������Ċo��\�!�:�^��+O�P9CU�sb���uZWr�!�j�nҔڼ.s3	�x�F����]�(�F]gI�����mZ��F�4�"r��Wuއc\�eZ=I����B��.l��<O	����I�o`�&��nv�i^x���xn��Y�X����#]��'���L��⍲�rƍf�hk�p�)[8:�D�����3Iť�/Ε�EG�]j��xeV����<�\H�fV���i�E�6�h�_U�1ea�v3���z��Tg�F�L�Q��e�t	�Oz}�#��kb�Z���4A�IU��w�`�P���R�Uܾ+m��c����Os1��)��eXf_t�lk���t9W}'rg譹�l���c���(譴��SO]�F�)��1��u�՚w
���p�19�(��Ѭ�t��ڻY�՗uv	1l�4�.>�seY	�k�M#,
a�<���AiIt��	�%�/=vnw�n�����Z��5dD��vt�w5�s��u��Tes�0�3��z�o)k#��4-�֋�pD�vig~2^'��>nZ޵X__n�LH��s�3�9��ܥ�v��x��n�V����5Þ���>6�^,F!�۪w��x_���vWgu�5��)�\b46˖7g	��	uC�e*O�	[�b��VՁ���+��L *pK�N�u!;{&�C�ue�38�ح�]�躋/��1�k&�:c:�Sv06�_Q�#B�����.���Ys�A���:�����v����:�c$�V��k%$>��\
���K��W�q*��]J �w#ͼu�Of��vF`|�䒲�0CºV�3��+s�]����t6&X�$��������_G��U��7{���Fi�N����N)x*TX�!�l��m��m["(oqu��7;G7R�}�h0!F-7G������Í�K�S'����	R���;{}��y<с����ŇG.��Ӌ&���֙,�x�:|.��;�g!T�1Bq�G���!�Y�ȵsW[�o{���9%a��Vupd�
�ˬpf��(w
\�k�c�C��@�۱�i^b!�\ٵp׳Q:�x\B"���\wxi(�
/xA���cz�/{2�j�a)��n�|�}���p���ـ��c-^@�[�#��/�J�骉��q����}��Q���g��jW���Y�N��j����mi��#VFopؑ�ِ�F�.�`��S�n�H���H��&��o30��t]�0� 5Z�X�T���t�b�8�)�iQ�z�gm��9�[$��0K\�;Q��(UG%B����wz�iUt�:�xN���)m��c�]u���(�W��t���Ww&�H��N;cv�u�L����KJ�Y%{[ԉ�%�*y��-�w��N�<��Ɨp�vme��ZhMQd5�E(�Z�����e-t�yi�^�C���_���TM�kyL���<�h\;��،�%��nJ��1�b3Y��b�5�T�Y=�c�����7}�]��`��fK.{�u���4�*�7_�+�c!�16j��܃��l�}�E�� ��a�u�PU����/Z�(�(]�'F�NZ�[��vК�%�1�|�
�٬�������}jbK$����4ݚ�T�)�ꕈb�\3�B�k�`�����̢'|�ƨ�K��qy��x��j[�Bĳww<�n��k�t&����}-Qϱn�
֝O'�/>I�zȺ�'+��v-	.�2���͝�����,��!���|�u�Z��=O����/v6eq�V+�J^nv�U��}3'm�`���1cs���1�ij�d��E���PU�g�����)���yA5�k��2.�����Vѭ��e@�J��z�ig'.H�Hn�n�n�5���UrSv-4qh��ۏ�vN���[;�Z�[V8*YB^%3�����hb(�K�K��,�tT��U�q�nf͍k�Zg�wK�zQV4}rL�MX7H�VI7wbm^�;�h]p��Z�(�1�d����u�!������ ��.��2���].{�{-���&'KB�[�޾՟ZzUc˒]��ε��f/��aӦ���mut=�3yC
�7�8|g�>���[��O��al_,�WF��-��Z����yn�n�N�Z���V�i4�=FX��݌�N�}l��v���F1�xv*3z�����������Rl]���~�{`];�sC�1Η��{�"s�F���K#C3��>Ȫ�՘�\zs�U�!��/&c#���qv���hi�D'f����^��6����1��gm�{z�HE,�ۇ��H{���h�We��c�v�ר9)�o���$�)=�Yeb���B�.� ��qY,��*��i�I�&�]]�Q�5�,��	ݎ�9�$6�5M!�� #]NfD��#��n��M�Y����rsM�ˢ��{Ds]3�u�S�Ym��J�8��P�:�T�so{C�������5�!�so�n�hK����(U:�ؾ�Z��そ���Ǭ���Ջ䵋]�Ʊ+D�Y�C���ǖ&���Me�9��K]�h��jA��Ti���j�ݏ�<*�،�
��w���_=�+�*��ê|3��1DA��P�lZn��B��bTo��h>[�jD��lyܳ�����X�)�6��٦�M�@%`m����fW�F��FH��%�X�����V;,PUǍ�4�Цپ��ˢ��}!��=��\rF&��}��q9�qO킧��ƢonF#�*\�ȨK�w6r;�י|zM]������(N�y����J�j	κ;�a��4��x��\/&>��j_jҎ�n'N���
�	�wxm�u�rK�l*�ʽ�ɬ����+�-M���sf�2�˛,���ݝ]2R�+���p��+�Kʼ�y��:%==�Yj5I3)=<v5���T�A*��N�W��WxC���PZ�"c���(3���k�%ۊ�Aĭ'��v��v�y��qW�6Rv6r=A�F�b�x*�X_ x�2�F�ߔ7k:����@�<�_IPǝ�Z��d��ue
`<I�XCu{��\�qyVs��39|�9�E#UQ���T�Wv�l�#��A�)ӈ9�.1��t� �d�t��c�)���[ڲ����PJ��<���K5�jF��'�{�.ôvr:5s</č��}�lefu���U���o���V���;�H3St�͚��N�XNp�T�]��wb2]8�2���i���V1fT�ИT'3X۾�l6���7ʻ�K�Q��LQ�<��y]9/���^i�^����9�טQ4d���7Z���|�[���hG&��H�k�`�����ye�S�;Y7���ݜD�L��}�No�
����{>԰�q*�L�=����Ӻѧx3�;���v�Yva4�8���p�f��;�3�e;툇N佊z�����G�̜��&�f�x�ѱʣ\9�7n%�
�yU�;r�LR���rS�5ps9yO�G�V� ��*[�(�ǥ[�K!�ƵԎ�:uN��}�4����Ц�t�����-�$��9�X<�����	@��(�y�u�kn���׼zS�y�Tzr�w����:��K�M�7�u�U�l�IJ�c�����.����O�)殀ڊp�H)ژXf�p��G�
��[�D;����~O���fu�p�iG؂��`���)���Z�d����β0<}8,,>���f�i�[T%��:N�4�������L�C_l��Rw�,�Z��Kr�õۉ6�k⺉���Εm�o��$�3\�V��N��ѵ�4uj�Ywr�gI3��.M�GP�#�%Ep�;F�&��,!ɫ��^�o�� %��d��;��g�[ú����-R!��RT��B��/HQǑB��V���ցW�z�������2f��ضw�}���q�5�q�i:�5;���2��4,s\:�z6܍-6�:}���va�ۻ[�X��!}��h�U��g�f<���0
Ȭmg�ls�B"#���[���V�[	�ZF�n���*�C!� ��k�T�G���Q��hֲ���$.�5ڽ�S^��̿g�t��AݛHt�9�'��Kr^��X�%o˦ ��Jv�Z����u���xkiJfʵ8ٚm��)\sk39��E�Y�Kb����@Ҭ�7�Q:�Y���<�7��kQ���f[�0����@&J��Fq��C3�uf�B�I��J�7̚;Wݺ��K���΅Fnhڇ��3����8^5�.���f������V��)A�n��|;�'੍GxvzJš��Z�0Iy^�ڒ��W�]
}�9�r�Ӈ^9V��w�X9�u_:s��	��BK�XN���ɀ-%.z'֍��K��Sa��*�t�{T�ԥ"1��D=ڤ�G�<���L��_b�G>��<A�|�5Z�����仧\:<l��p@���k�-=�>Џ����&�1�OGv�s��Ss�&�1v����q���l������٪+�@OuK�*�'{��ɐm!:h~�d��a���_QÝ8rX��e\��*���9�c:G�&�G6�b|'�`��ki��W�ܸcqoC�M��	�0:���}�%r�xN¥xF�6�2!v�p��\�̼p�lW���<��s�l�F<4���%�=�H7qn=yjc��]JOy�űuz!�Ȼ5'����wE͍�
�'k�.����
u�
�:n�0=t+/�z��ʊ�`b��ۗ�ɧ�$a�a�k������f6]ԕ.�!*��9���y�6��|�b�(�m�5�����Q�ܦ�=��i��0Ϋ������P%	��u���;0m{NB�	��}�;��砾/\j��a|&L��鄯�Á�R��Ȝ�BahnZ�ۙ����1�uד�Q����1l���e2ا��x�y��-U?jNa�!��Ƃ����g�� �Yݭ�1o˵[�j�c��������
}�G��������}_}�V�o�;���"�>�8��E{�н�X9��S@t�!�fjaF�ڶN`�uep-��A�B���js�*97��-�1}�Nc���浊�[]3ls1Ѷ��"J�۠��^��V$�bhD]��O��j[X����[��^�g��{�K��x7�ɐ���;"ִ��9޽2�=w��KVy�==`�ţ{΍<�MO	�L5+taAm�w%r"� �{R���SP���Gj�zv�ܦ����zq��Cv�N9K�ڔ�{���7�/����J52cpW&�^�w{�Z��Pk{0� C2�[w�{��[4qcPS�:��J�d{�cہw��TO�����*���>J/>y���h��ƶ�(VVep:��I�OM��i̚'��޾�)ŃIy�	�}�5.��61@hr�x�@�3�ofa'�j�e-���^Pֱ�dO�3���-f{M����q��=d6��z���Ze��X�.v���9�[x�v�p�ze`��7��m�~[5�$��3
f���y�H�i�(U�GJ��4��0�����q@�	�Bg�s���\}-�Xi=����(o"K�_hg������	gs��M�/#�j���D�=v�ɣ�Ѩ�;^�{�P���rI��`���XH�s6��c�ek\�Z��6q1�y {�t$ϼ�cMMl�:��i�U+�E�p8��&^]�P�Iba�]�9�g(B����\�8\�s�� �,��$����ĩrćF�����BE�K1�]2ֿGđaZ�E�i�֥A�t�XM3�a*$YT�^���D]2(*��QH�*9I��Ppr�I�q�9C*q��W��n46U�(JP���Ù)�i�p<�[\`�4(*�		�=r^�J�ˉ0�rC��	ĕ��\
���M�L���tR�Mi!+JJ(��2���kET$�;��Dr��S#Yf�m��:^1ȬYv��0q\��,�Ȓ��r�08��`�8�B�i���$�:gd�bjÔg
�X] �r�J��,3�&�D��&Y��9��ZS�\��b!���p�����g-NA����˯�:>w��tP��N�����y[h��s���@�/_G����y{¥a��)F�T�����Mkɀ�s��=��_Yj���_O��;fc�tE�U���]PU�������҇
��T���~�S��g_v�;�\���4����u�����#�O<E����h�/� W)4��w��0f�x1Ņ���l����S�+�`V�?3��'�X%**q��/x�V�aJ\�\s�����{���<���N
���d=�'�B�r_���Y��u�����σ�ӫ^v��Eq�X3YH�Wo:���r���s@�'qq����0Eh��i�`��R��m�pqa�a�X�'DaB}���<)+�{����V*��D&�oG�кο��o��n:n�پ�����l�K����s�eP��xU��`V�~6��E��]$s����
�k����_�w;�|�/�^�k�+u!�u��<o�z�C�K��fHBr�.�����S9?�!�ۖ4\F��+N�M�_�Z��XH�D<RV�b	����{5gf�e7�tY��5)�%���:�c/|���W�C�>\�V��f�=ί��U��%��>�O.����B��Y�
��}?9l eͻ;�x^v���Y�a��+��tj��ά~T K>m��>���鶮�}kv6��R�WֆM��n���=����nۊt����2(�Y�*&[\�N�ޮ�rBڱ�!���r�0^sT��t;����n��k�G��6��7VO��aO�;F�=�w;ט��![TV�ڭ��{`t��*������p���N�{gӴK������0���z�$�����ޤ���;�ET��Cp�w�T.��lj�ie��!��zj�;�fa���ʾ���eꩼel���N�U���~�tOqɋ����|�������wV/L�{rkW�-�s:�D?��R)
H��2��?X��ON3�x�:V�%�Ԋshefo.g>��8�p�rN;�5qP�*$
��q���[q�$}�~����L���7�o9r6�_u
�Qʝ�����T�xD�/3��U�'ɺ�w���V��y[�"Y��B�u���M4���L����O��0)�^�����}Af�������W�q�袒z�2C���$TF;�O�\^�i6�҃'j�[D�!��{��3_�K���}X'�DqW�ϯ���ux�c���N�|��#W����@"Tsnu������8/�f��g �J�s5��e]�� ��{֑Wi�k�p�:C��8V{�B�V��{�Z���t�[:�RQ���V
��9W�IZ+v�	�8��&b�Hވz9����w*m�:�d;]�^j�k��\gvQ��d�0;4��]���h�n��v32�x����̙���N�d��s�%���jי�T�n�����K��<�%j�p1gqO�N;ˉ�/h��o��c�xGQ;=d�B/;�qQ��7KI�����u����Y�<�UI���߷���K7R	�Z�E������M���74�"1>(���̤o&_�2#Wu6~Q�%��a�ꌶ��؁�2�nMEqL76�e[�{ݜ���/Sp״�V�pq.��Y@qb�͗�9|J�����<�����i�8T'�t{������ʮf��@���[ǯ�CY��9V�������o��n��]��'��ܿ/-�d<<U��P\����O�#�g�F�+�ھ��o1Kb�U�ػ���^]�����o�p<�Hq{Q!\a�7����ȁ���3k�sX�z�ʅ�^rY|��M���;�}m�c�!P�p�C� 7���1718L�$����,��>����LP�,��b]���B��Szm��U��&�Y4���;�+�P�ݦHB�2�{Kj���A�4�G;>�����K���9��J�y�}�,4��,Q[c3���A�U�l �Q�)K�T�Һ�ه�r��nݧ%�3%��q˥�һCh�@[Uyn��òk��y�,��޷��?ڟ�{9*�vL�C��r��v��@t�.��{�l�����"����R��@s��^M�=�xO��Z68W�}������:�>����FY��N��'o�s��Znݱ��a�d҄��L�۟���ٻP�6���d�g��	���`<J�@�����\��.1� G��U��f�=�
�7&|�Q6E�V������,���X��{Z{s:5^sx�^�����裢������r	���r��,BWF26-�{.Ǵ��u���$f��j���`R����x�k��q:��NAxwLZ n�\��ȭ�ݨlQ4����h1�0�(8�1B�:@ŲC�δ �h<1�Ύ�{|;9��0��]����T�&�H7eĹ��&aY��QB�g�� B�B��a��2�`y�fmGN+[E����+�h�BX��PiM�lq뉯��V��9��c���U�|5���r��.�b��pOujSʴ�:t�W���@���+�I���W 4Q|��9��ю��OݽU��C�	�9�Z������+NdO�è_ ,0�|W�R���ۘ��
���ܵ���9׹������T�}��V#%�Z�/L>+e��SM̹։OsT}�QJ�a��b���oj�E�����^���yW4��7lg5<3ea��]9z��EF��.8���);c �ԣڤ�H��E�ҩ �*����ֱ̚o`�0��AZv����Ҡh�	����N���JDj�#�R��C[�MW$Tu�'����8S��:���TP|x'��Lc k��\BeɄJo�PN��_/\w����5S���^��Q�'B�d�1�
�jB�X�f��ހ�� �	6�Y5��G)��F+t�r�6��[aR����&\)S��~���sȮ�8xi>9��� ;�06NlR_pܕ������#�Fk��s�F��֋��[�m��Q���(܁�U͛j@l۬�#� .#ޏ�뺨��`���[��^��g��J0��|��x!J7�\��V�Ɵ't���ڒj8�Y�R����cZ^������:\�Y��z���%˧Ӡ�e0;z�C���-�s�p̌��#�=V!y��tQ�����>.u<B�K�B����ٶX�Ѳ�����3�@���@�˪����J�U��놝�w�����d�R�l{7���g�g�>���`i �{�7��04_Q�k�
ެͮj�z;iؒP�0���t+�+;պ���s=iWD��}�$g>�� f���g�ʹ�81-�j�M����W��B�T�a��˕j����q�M>9�O!g/�b
ܞ{ �<~ T�@X�ؼ&�U�2�S�$�"{�>��f�ӭ�B^�w�/���g�����#� r7 �2z�X5�k���L�yQ��M�7�-9CF����bڐ���Ń�M��=+�ZX~���~�@��!��]��&/�W��Ͳ�Zr"�Tp�q���Z��%�]HA��9�k,+�-�#]M�{���レ�ʖ�5Wʠl�pd2�)���V+��vWL�{վ g�v�#<L�Na��;�� ����U��ow��'�c�J�P7K�F�[ǐ��:��ش�z���w7����lWi����"0dJT��1��L.躍R�]�0P�;Y��g�.�kP��լg.���%��ׅ4ŏ��O���=�q��c��ݘ[��F�,��^�-���f�p�$�̇D(RcAlA��p~X���S�J�x�4��[Y�6*���/^���B�e��{@l��q �n���s�;�p��ɠ<F�/�TY�,�x�[���+��ґt�F�+�p p�%k��b���(��������d��#�W��,��]�����GE�u��b�6��o�3�&f��K�uYv6�����-km9'��[9L�Ɨ��o�èy�%q�Æj�j TRր���#^�ZR|�,���V���t����ۘ�3��>ޏ(z����y&6���4@�;L�>��\����7Q����A�Tic8�(dG.b���3�cB� ����O6�}�A>>�Y�mG����t�U�/�倦�����	U�!��0�А��=[4y_s�G6g��׹�,�8��K�~Ҳ�����X��e���{��o"�쳫���h:��T:� ��",:��#��y"6̪V�\��䭟Z��>�U~6��� ���m�W&mbѐ��`^������&#�JQ�������6�J���'g��[gO��y�L�G�򀜯R�+X�-/�^ћ<'�"��7�O�r�����~^�`�7�-�΅{��a���T�&q�&{�Ι���?\cT���c�F��O�x�β�stE9�LWjj��V<8L:�`F��	iWO��t��U	��~s=g�[w(f�>�JT�J���*
R`ɂ
��Y�Պ��>�uS��^�����eKЗlȐȖ��^�(�a��'w4k���+�5�����*Ɏl[4m�˜�dx�W�i�T]�)�إh���dz�t[[<���R�����T�w�UhOط������]B���s�-^C|��Z�����q���ˇ{*0�:��*�ʵ�Io�מсM��/b8�v��\+����q)�ċ�Ed)��Ƨ����45�;��]�#\R�q9�3�ֹ�c~��%Hy����g^pѯ���/���bB��	�����HR���h`{J�<�i�dZ32�T�D��og����w3��L�A=�������g���j���=�˶�Gs��p���Q��s0Y�Xb��9�ȇ�QᯕNV�y_�W/I)=������ϡo�{�I�yBh~���=�9d��ډ���JQ����mZ(�eI����y�FG[�7T�%��¨yc�9R��%[�~T��VxW��X\}�|jpUẞ
i�j��"�q�=`n�����o��rģK��x{7j���֘�c&#;KR]]u����D�p��lsG��>3 #E|�V���ٸ��a�σ��&<7ߴy��S�Xg�mX�ӻ���șp�b1�T.�k�����m�n�LX�@���e�5��ܼ�\���FZcNzu�t|�^��-L�]��j��3��V���O�Ʊ�`�S�-�.p5���[��~���U���E�܌g���<��#�}Ny#.����:��[�{8o+d���1J�-�t� t��c-��7vJŵ���$bw�������靃&�Y�{��,y��34��.@�L�q��[w[=����;8%^�a�|����e^� oݪa��t*��84�T跗�dT�(k�j�K����p7Q��"$ňꙅƠu+��o�
�fBk��:��u'9��]�Ŧ�7gS\;,'�-��\oi��g��j;)?���:�D���%�;ٟI躷Gj����~�N��)�Y����=ա'�B�UAT��9@��ʣZ=;Uꝯ���Ę����WU�(M��9J��D1�m9b+��	t��;3����:�BM���Vz���������,���X��t��K�B<#EE�b��%�2lR��^��^����\��d]ր- ؄�a
y(u}{_*(></����ȍr8��U�d7,�qg�s7��֍O}�K��VQ��t; .1z
�������0���p�id
��.R�����|iN#dH���#aAhѹ!�,�w��B�ı۽zs&8A���q����UU�q����,`�<�)f8����7'���%�#Φ�E���:��F�{�>I�A޵w���{tVb���|����t��<"Ɖ��nz�������N��]��\n��D_�>cc���oe�Lƾ]��gV���]	�fy��q��|���*�~(�ρ��^���>�Fѻ��P�^�e��AbC:1�kV��d���Ӄ���ӓO�e��:���d�v��XYi�{�s���wO�Z��.�}��>0 UV����'�X'����ܽ��i��k=�"�1?4g�u�I��G:��qQ�����;�{~�Ɖ���f�K�΀�fY���T��1{7��ƶ�?��Vr�S�����yg��TEDn�G���5r�+͉%i�����-�t� m�Fs�*�ib�	È�
 h�@]�m��`Bf�w���Q�v��8N?�R��D���Y�K�:��k��{p{+�3�X�)�����'ÿ.�ߎ���\�u���e�'�mN[�5��lL��.���^���4�5;m�e�����X��М-v��;�#��P���Mq�$i�U>䰘�b�����w��]�f�v8�x��������2:���e3�U����Zu�����W(Q��Nᡞ��N�`=ja,�c	���W��)��:�q�e�W��m
�Mz�eߎ�v=��)oOw�٧�G���I�t�x ����x�R��c����D-��D9�0}�}�Ț�w��۽�ǐU�Gä�Lg׆�?tP���(��GZF+�ٸCTJ�u�\v�Qf+�8; �W;�]l�:����lѵ�)��'��F��`����؊��!O�h�PY�V�͝�Ht���T�Ԉ�9�h�|1���&���C&<[r�&{m����g�ǜz��C��r������B�$v��`�y]iV=As�[X�<�5�Z�ou�H7�d㛜a�E�-�p����xJ
�jsa�tp'hd.���
�Z��]4Z�m	)�k�g
�Ʈ�Qo�=�����v��u���ש)9�A,�MDR��HM�y�m����ʧϭ��b�� ;�s�+�$��m
י��2wa{x��G���(ig��J�H$p^x���AJ�\h�긺��F֊˧��:eֽ��+5�`�q�жd��^��\�Q�*@9�a��l�}�+�f.���|��
W��C�wOv���}�]n%3�'>�1��~}V	�萄iS��2V���Z�D�T�<��kO1`�Y��	=��w��Q4S��)Ԕ�l��<5ڭ�ޭ�c���Ӱ�c{a���5\s+H���ᬾ���c� Q��n�J�%-�}**G70sZ阵\Ւ��Ort�Y,ـd��H7��8����-m�qAm�׷������)g-=�ǘ��6XҖim�-ݕ�$�,�g��V#SMJ�'3S=d����>T���O۽��#�J���Ҍ�SI\�ڟ�f]��M�P��A�ԓ�㢪ᒅvT.Q�A^C���0�G�s�#}{�>�C�4�� S[g�B�ν�3Y��7}�W� 7��j�.b�F�%�fI�8�:�&V�U: n�&`;�lQ3Qp)n�|'��Dh8u�梶��O4�vg�>XB믦��m5�|LNf�I��`kĔ�͆�r�mhj�9�טּr�����F���wbĦju�]O�V��w&Y5܄�\a�e"��iR6mOV���I����k�e˳��}�=�.^�e���Ʈ����x��W������siK�<`���5'9�;� �̓����4�����1n�pM8;4�՝0��
p�z�0D���^R�oSNvJ�H����pv��N��Hg�:���ft�Ze�`\�f'��Ũ�:n�Vս�B퀛G>��uaT�SH����(��-^ ��/�������z�"NUC���Sw�������<�U7�v�3��c�S��Υ]�/��*d�ݿQj�!`<�g�A���A��7��e�,A���y�Ū͝epA-���/6���季ٸ���'�:�yG�$}j��Hc�g0��<fTx����t��
a�_hZZ :�E��{�YR�f*�҇zl��(���eHV��yay-r���jβ{*׋ۃ+�ߞ`�| .y���,��՜z��f��&�P���l�˚�;��}�ê�3f`[�lW���3��{8��K����J�]�t�]�$�ܬ��"ggt�F��((�"��Q���\q	.X�ʳ)-8U\�TDr��9p��]V�1
E+�g0��%�`DV�"�r��(g����\��Ȑ�����0"�9�J�����
��ͬ�\���	Q��%��XB)���gJV�r�L̂"�EV&R�;�+J�����C�kH#�&�U8�SKJ�E2�YUf���U�QT�W$�D��JGT���Gs�F�Z$r#�VX�fAUn�pʯ3����PXHQU�T�ȡYl�d��r���aY��G:�Eu��(�q�q�T�%e$\�I$�fE:ar� �8hUˉYBlR�գ.ADx����NZDu@�(��s��U\9gXN%�U���˪UUs�D\(9Fj,**�G�ET*����ו�1�E�Ou�NR8u�xӺѵ8�k�� ��_iP���1�
ݬ��t7��n��t��ǵ-��o7�������8���#��m>'i�S�l��|w^����z�S���p|g���x�i�n'������OP��}�v�|���.�ߓH$��G�}��c�DyD��88;}������9����^��C���M����o�N��w�}8;wNӻ=������0������I&��?bW�8�>�ON	�t���ӏ���M��w�x��68؏� #��>Yp�b;j&�վ�SZ�3���F��#�b=�lň�>O�n;|��ω�o�I��7��y��;��W߽��t����O�X8����$=N>8/��]����}���Į�:�C��޻��n|9��?��G���y�T��CF���$�A!`�~��q:L*�����&�	�ߝy�`=N!�ӎ?��~N��N����F��N�7�st��i4��BM>'���\����@sE'U��O��;믿ǿǡ=��ӷ��I?;~x���7�>8������&��;�:L.����������&�u�M���w�[q������}�;@�pw���c��DH�#�"�Ⱦ��I ��J_=�nn��_���P}DV
B��b���C�{�ݫ���?'gθ&��ӷM�H}M{H~?X�oP��ݜ��wq��<Mv��n�q���]��y�I��@����E�>�G�B��)!{�<��yM��z�z��>�#��|DD����8�ޣq�!븇��v�&M���C�|C����}��{�ۈw�A�t��q�9@�'���s���">��"/T�c�,�" ��.o��}쎹�y�ܦ�{�"!�!���ъb�۴���_:���wj�]��(s�&�ۏ����8�x��|:�ô��}x��c����w�>�|BM�}���=C�~zC��v�'?w�·��O���6�KW�h��DBDG��]o����4�~��7i�BzO�n||�|M��'���[t���8�yo��q���v�޸t��O����u��:C���>lw�>&;�������8=u�a��A�`�[�x��7`��z�@��~�������!��?��Iۺ<gv�P�}M�����U�v~��A�����Þ��W~M;w������O���Ͻ{�
t����N;1G� ��|�B�fي^���IQ��Q��Mh%5Ӯ�����������y��[�����l!�=}�okZ�w�ƞ�F��ds'u!LK.��ˤ����`�4(d�݌Ŧw'z��06���m��R��&�)���r�d�u\���2j���鞂�{K}A���������]�~��,}T�V
��a:����0���I&��]��L/�>}�?tx�S v?���z�O�ާ��:���;�|<��A�|L.����!��C���q�Ă�_Sq�W�)����xT)K�{����U}?��ձ���>8�m�8�w��ˉ����>~�������M�yc��;����q���w����������-�;y�K�=P�������"�}�!�y�O�o��:O�ݻ@�����\ߟSqē�}�ӺC�ӎϗHt��'�=q�p���q���v����w�s��z�����}_��9���9qW5���E���A>�վ�񏠈��O���[w�v�]��=�N��|N&�8&7��qS����<C�	$;�cק;�9����;L.�>��<"8DP��(���p�wL*�_=>~������w�ӏ~�擤<M?��ǟ���!�5�^���i�Bu��uל1�<O��t��Ǥ��v�M��x��ӿr<O���twC�>���!��[Y�������w�k����Ʌ�!��OO�xo�����!�z��[���ω���'|BOǿ~u��w��׼�i�	7���p���|����,����8�L���>���D0t�A�z�=sٞ���o���S}B����~|��!��|O��N��C���~dާ�q���y��I�BO���<v��C����ޱ������7N��7<K�se�HB>#�˾��b�ԧ�]��X��DX��!=����_ �n {ߜ:E��w�i��m�t���^;�[)�B}q��~N��	ަ����<�������ۯm���!���@QM�����[�az@�O\��d�ڗ@�.����"� $�޿se�ߝ�O�}<�N������|��8�z;�~qڻ�ӻ�c��SO���uc�C����ě�'��8~v��ノ��랦�ӏ(Gۗ��.�=��5=Z��� |��I�}��Δ_�;�=N��������!��q��{N��C�u�8�L)��Ǯ���q����A}wH~ߣ�M�����;t��C鞗oO�P?g�s�N��*�ʴ�K��O��m��7ޖ���@z��xU��E���c�E_�0��[5��(yN�ZI2f����qѹ���zC�J'��4�}5�$�Y��uL�[�L;ǳF�wu�+`nv?�o�
�@�{���n'��m����8�i�?!�q�s�0t��C���]�um㸮>���7�_�ߓ�r��������>��?'i��?7���z�'���� ��D}"#��r��7�qx�}�l�f=�G�G���1�Gт"8A�8�;��n o���v�+�&�<��v�i��>��9��q;C�i7���.���;���z�x�����s��'��������;�����ǷۺU~�}���E�}l��=�1����Rt���W!����o���_S~�8��� Iy��X={w�O����aT>�=��;N���>���c�qP���ۀI!��~��������ٿ;ܾ��@_�����Dh��D�{���]��?7��۪���?�q�;I8���ξ�U0�������0�������q��~sz��t"::��""DF��@��;�Z��n$��L����z�}#�"4F�z)O�Q1�}}~ua@�$����v�v��?>�뎕�w�x�N'�?~��:M!�������:v��[�v���]�w���o�_���������ϵZ�����֏'�D���5X#�OS��>�}M<M�~N8�׼�J��$���պL>@|Nv����$��GN:w���q��N��J��~��t���'�����g��}���n��En��f��3� }|G�>�}߸�z�;|<󝫁M�	���m�������?yѻx�ߑӷι̻������0������ݦ�>c�q��O��G����;����//{,yj�H��+�E���P�� #�T�q��C�M�q�\q]�����!��y���ݠ}IǞtN������ރ�q������N�x�='��8��I���L*�����ިu�ET�@y���$}#DP��@.	�x�O{�����aw��Q�C�>�?p������������ζ��$���������}�ӧi^�'��y�P���|�n��红��f��|e^vdt�jaG��#� �8�����:M��t���{c�W�}��o����t�pO�����<�<¥� h���w��*�:�=z(Pa�=0O���F�����Ks5���Q�F*o%f���V;�ׄ��B���w�6ˬ�YO*�k��1
�F:L|pnɑ���ݱ�{Z�Vi\7v����y.��3=F�Fs�ǘy+�X��PZ����Bp����ތ��/�3"����j�dv *�2*�S=� ��.�P�ί�|�([sa���m���r�E��V���\���T����f���tݳ@`�6J����҅��b5lYr62�6�Yw:�T,��m��z{w6ʘ�jCSq$���	���պp�c2�L!�c�̻��[R+]���l� �^X�Ԁ�~c�����!�_V���a����,;��t�e��vϪ��m�Y�2����+@Vq����뿢~���6�:�]W�z�?��F��~^c~^��18xi�ߣO��P���`�|�Y��h�j�<��R�oG�z����{8'�Ԑר�h�j���+Ek�rP�u��9Ș�g�J���/w'��or��InN�� ��DpÓPxP�p�b� ��B���s�`]����;��Nd,[��[ sX�|,�92�W;�����hq�����7��� [{L�veҾ���MH��8�ڐF��J�F��F=5�G,�ӹ�{]�1h�[KY��/ў�f��Uӵ.�f�@���`˚W?f9Z ;���.=N]�ox�B��y�++m8�e�1#�ή�Li�ז�YOmK1~9nW�J]XCS=�k���5ŀ���f;��Ȗ�:ݠ��fC�Õ���Q�A�fq��w.��fIg���ڎ�����.ûsp:�!��l���cr��S(`ߣ^��]�A'��^@��3T���b�A�O�2Q��>S�i��L�7)��b��
�+�{�C�^�{��m�f|���>͹�Q�L_5�!�]����G�s�����ϵ�eq�^��I_��#F�S�j�ս�w�r4#�tR�pR�dUXa .�y�YHD�9�������^��+�g�I}����K���;y0��^�!���U"�JT����P��4 t�s;��p�n��V�V��P���#E�\l>����8ӡc��R�AQ�=Ҿ�5=�@u�x��xb1z8S�C�Uk5
��&j!���	�"�]H�!�����L!��l��+F׋WN��{��ΰy����s��-�6���o��`oz43�� �t�r��IS�#\��js�	`W��"`1�~�n�n|
Q�b�\%N�b�g��*����28�ElI��R�R��.�a���ϭՏC���c��a𷩓��.c���QX���X;�V�'�H��ۊk���.��r�\3��7�wb��=�B7�����̓�w��lYG9��n���_�Օt��#yJde�쬈�٪d��i&�.ap�nGJgX�>�r�B�h�,H���� �.��xl������]na��u����7�;xe��b:ջAn^k�v�[���t��{q�VWʸx+�:UR�,��oU��Q2wHf�'�"�2�B�w�G��l�Ê���c�Եa_x,񘃸�w��)�m��y4,����f�Ҿ2dTBrF
���f�:����Q}�{"�VxV�'''���*���V����"x/S��']Q:tF��Μ.'���[/�a�{��'g�<�Vc�Q��lV����ʯh͞��I������fA��=gTd����ޖ�
x|�݃��-ڦ�q��|V%T#�;�����-��u�C����ތ�������g�t3����C�i�)�k<xJ��������(Y�c����;zwMa��ұbݼkVo��Თ\����ʲWy��U.Un'�e*���+"6���	j���8����U0᮵�Ǿ���j�ˆ3�x��SpK�����H�����3�׹C�4���D^���1��9H��Dr7D�yJ�&$u�qPH��qj�yG0U�%f�7P,^)t\==�x�AA����"�{ǯ#�%�(=I�X6�Z���� }��E2z�,�̌�1=Vh��}���H���V`�3�	:vhV�{.�}�p2��C�DtH�p�wW����
��b.����Q�����W=6G�b�ԅge##BF�%񯯺����I� ƓxW;�%<�vXQ�A�դ��j��\�0���&%YU��0�����1q3�l�v���������!9{���S既���K�j쉇�[��D-��9~t��QBiU>�H_���X�
��s�U���e��2z�̿q�C9j5`w�s��g��ꖿa��G]���9&�
澍�0#�e�F����µ�a���X�4��
j���&9��]L�ېf��y�P�6��5��8i(A���Qn�ǎQ�y#-T�6�`B�N��v���6&�XVvL1ܣ#�`���-�:� 3���Ui���ff�LGt������29�(�i�?RkqO�`R���]rB��z�3���V  ��^z.U���P�_!�Z8�Wq�����s�q�Q%�w�͵V�_ZZ�(��$=7*@��B��3����UcC�*�p���׮���n��%�l^v�aU��1��ˮQ�B���jϒ���k<TJ�e�\�!�������X#M��:���ن�ww.]v�(EH�oou=3�z�z+}�ܱ�~�����f^
cn��#����84���慔��v�/��%W]Y��c�\���r;ͩ���:�.1��V&���vo;��C�;���i%���J�΃@]!I�R�us�KS�ݙ���V����Ͻ���t����g��/F�g2�Lq�O�/<�Y#�P��d�|��y�`XZuQ���7)��rƎ���z/!*":����v˾���<�g��=R����*]�����:�c�-1��=�r�W�r��Uo���lT��~���o��L��v�>�P��x��Rp48���
],hv��F2t�60F	MT>5�SJ�3-�O.�]Tp?�b[7UY)$�-��7G�xI��1}�G���O'��ySWv��I�z�@��?*�[����f���Gf�v�2pz@t�X��њ�u��t�|��#�3�ŕ�}�)z͍g�νwt�t�Sr�9$=*��]9���3+{	�K냒�.��֦j�4�{��X{��KB �	�4�܀O�u�9����3E�suj�s��7�{ڻ#���\�Aq\@��s�Ë� ��8 �����G��o°/|߲w(m���,�n�
Cs����6^'���l�f*98���V��L�f-Е��e���t\��w�׬ ����^�>B;�&f��z7��_)�A�w��
�ʺ#��e�ł�g�*|������g�(gi������&���z궓����C��;ϱz���s�n��^�c'�����ۤ�����F1�*���F�����R��xvz��80+8��\�3[���޷��|�j"��=5N9�o7j��vm�IOr�s��z�;���Dpʜ�B����V7�_/
/�\:6!ܯ_��݇3�LU����޻��ˀk��_����j�<��{p �=��B���A 1��6PH��]��U�!�� V�g�]p���/���~֛������QATem�WpyKs�E8��-ˌ�G���%��zf��CK��o��,Fi���jx�bڔ`#b��@7���)�g�D��q~�|jY�}�.p,H�&u���L!C��Rj�Ya+]z�]�.SՁ�À\��\ ��1�N�,�(vL�j��@�L��C=��N_��"ѐC�WwkO[�[_P��c����]@.��2���*�6���8�<���k�[�f�9���Z���E7� mZ�����C��p�6���b�zm��[I���j�{Ao].���}ktF=9��ؔ��F
���]��+��(q�T,}��|���{�
�*�b����)V~&l6��tT��8պ2�Ғ�����m��0o��M5Ӯ���?�n���'�����&x9c�-��oɯ1�������S�|_W3jI��&����<r�i�L,$w�]�Бg<z�z��Ǳ�Np��楙Fl�_}_}A��;��纾Bb:��L�f���{�8EC˩��tB!�,��9�l[����[�sI�P�'0��� ;;ϫ�+iS6˒^H�'�!��H�u:��Y���\�OS˻�����DU}q�#�;���u	�Q˭��'禡T��砻����=ڍU6ҍZ�OI�[j�\M�\��X��^�p��X|-�d���0bX�3z�*�&��:Z�l���^����t���;^k�v�Q�n��0�&��S��}0����ft��|M����py�E�puO_�dC����@A�ۢk� iy���X�H)��!N�֥oq�������*\m0Ś���UC�] x��2$X��t�|�H�7�䡑�l�r���7��%� �ת�M��5T��V�)�)��iy�p�EDsʑ�xF�?���o)Q%?L�Slص{�9�B��/�ثb�e'Ư~8�;�\��w�?(�+Fޕ�G�6���b]��՜�X����1!��q%�J:dF�.��׍SA�Um�G�T�}) k.+���wHLJ�:[���0��J���d��ۑoL���p��y������(Ȳ/bIbap��
�#�m�=ت�	阄�\�	[\�e"3-��ۧ�+���;�2��3�[|Gk7b�����-�d�Q�^�:�&�Ͳ
͵�3�8f
3	�f�[�)���&�z�@�NvUC�`:i=�.�s4gݗ"�x�ݚIp��E�zkGx"9�&<�$���-�Zv�G�'2�y���63�d��d� bo���q��u�tL��� X�)�;kwo��D�d�Q�n���xEwZ7��t�8OQ�<q	wK��qt�ɍ���T�ڬ�4!3�}��eoe�;H�؝��Jqfgro�;%ּ����$�Y
�r�$|�]���n�Q�6!�i?KLg�� �N�9W#;��G3®��DOMdj�.2��6d��[^S�P�h{��4�z�7N����'��[���.���,���C��6��ӽ�p���_[����e9N��n�`yC�E���Y[�l9m����<8�;�Nf���2�j���&�.�#K��X����VJ]@��S8�b٨+X�p��y�ۃ�m�,���o:��x�zS�2�X _���6�r��B"��M�eK�f�g�i;�67��V�-�8ق˧R�kv�6������*d�U�SL8��%� ��Mk1�oy)�d��d޾w#ٗM��f�+�[5S�s�i�����2�S=�;q=EK��������%Qx�)#�4r�4퍙�m\�i����[Ra\����cx ��m�L�a��$ֲ6��\W���s����9W���K�C��&Pb	��҂����iڗ����6h���Z������g>Hr}��0+�yIv�
��m=�[x��`�D�g(ʇ\��,bgr͍�h��Y
݇UA�+���������>�C�\����w9{��A>ۯFց��C %}��g�)0��ކ�YcY2��x�	ŀ�s�sV��&;�VwPw-�[��������o�	7�YNqrI<�H�v�΅�F�K�t��WZpt�eQ�y�'[�|\8K�.E��yq��e��F���*[�r%�BCaR��I��H���w�T�o}��M�\f�OMY�O��ڽF��(w7u��d��t�fh
C$���HzVO��5��	zt��<=";���/��|h��ԟ�U�8���@��u�o��]���*����^�]�$Q��)\g�?Aw��G8��e2.���+(����1x�<�IY���u���4<�9o2h]�󹒶]s��VB!�vyn��q���)�{I������ ��!��ޓ�%�N����	#��G�/��[=
�Ω��^Ɇ�j��9b|��dL
�һ�}�[�dO�P�y[��=�;�o�ZL�K6>�Na�.DS�)��1�9��Ss!@��������U�9SFPBa\�*!���SidTU7�E�uK�D����\�ITP\�I���
����.ae�.�Dfɐj]��"K9.J֒x�""�q���HUV�d�9G<dr�.IY^�W!�f����HUȨ"���
(��VAT)uB� QRg ������Ϋ.����A.�q�r�(��mdEQa�R
̹\�R"�r(�է&G����9QL�PJд��x�t��f��r�[L�R��DE��9QAh�
�.U�U+NDEE\��
�(�:�YŹ\dA"Ң��uB=r^
�H��

�������P���T�eW9�̃�.�-Z�D�Rl�p�
e���i�#��]D&��j�e\�PW�+�!ap�t�K�gI��Vh�DZ�U ����92�겺�5���=<���]~���6�6��M᪄��=��t�핋@aح��^����7��s���k��^ۄe�J��>�,8�RW���Ua�i��t�����##9��ו���8��5�<%ZU��K���Y���q
�xt���ɲ���;}3��t�4_���Y;̾R�r��/�)P�W��pp,��Jy�KZT��{�[Q�u?Pq��5LpX�!���|�n��k<zP4;���q�H�ǳQ{���t�u�vL;�v�4T}}��}	S�����	����祀�bG(� r:v�܈��X2/�J�}�P�.M"Ex��5*�xo��V���7]tK�����M�߽��]��R�����&�����Vr���T���KGe���ׄG�٩B�yMȇ�r�ʥP�kǗf�NcNM�Z��4%,g�*"c�b��eI�ľ+E}�h��[Q#xs~�1�]uᮭք�9=/JӒ!��<��5�;U�HՁ��>��yJ��i�Q�d��~���I�(C��7sC�r�K�H!Aƻ�&bBd�'Wch����F c�~3a�7ji���	ȑ;<�{d=zj*u����1R�e,���'z�oUa�"�BuL<���q��0�zg��[�|�>d����ֈʊ�����-�(��:�3B�I9p^rK�Rd��b�RU��g<Srd���l\��u_v��_��HH�F	|.5��#��d]N�Pg;A�J&�#C��ծ�r�E�둮�L���7��[޻��y�cH�'b���}�U}�RʼJ{;��h����=s��d����N�Ω�d��b������T���5�/k��^��rޝ���5���ս/����ʾC<�V�b��E}�/��9����� *ɩ�i��vou/Ub�l��Df�W�W����/ʘw��d�� Y�uyn����HgJ�g�F��V��o�ȎTQ�ٗ�>�#�f�u,�f�l�j������N�NM��ѡg*X^�P�˛�W�k�\;T�RDP�&���0��h
?ӛ9�/��\��9��¹���j��۔�vS�8X�B}<#��y�HS�v5c���Qk�w�Ǧ{��B�}�Q�Q֧�9���P���=D1�m9b�Llڔz/�d�f��n��ܦ�D�"$8+h܊�R�W1��������\r��/���خ�K�ȅ���;n�}�{��S�q��
��Hc���l��^�ژ������.8K�'�N������n_ڤ����)��N\�W��bZ7D��n٧D��0��W(_Ur�V�}�t�nQ�UB�P1y��t��%�"貍�g9rP>�>�yVs�x�c#K;M��E[Z�כΚ���>��8�k}����SY�W#7f���J*:#&_SG��5&��/:��r��j:.���V�U�]���U���:u�e����}��_W׻Ϝǚ��`@���ˋ�Zx���\Hߠ\����5#	
�c��V͉�Lȥdm�7����Z�O�0�Lo	B�mZ(ܱ�
 ��Wn�����5�� :܃�}� V��D����#�,E٬����
��sa����<`S�yrS�&���.)'��mҿ}{j֕�2#�u���1����LQ�ެ9���'/OHyY�k�����]$���f����R������+��O�|��o!��B��]��0z�en�eV�/�)]J1��ء�8eNT!a�B,6�\F�'�sٰ!t�wt����[l��Ъ#_�Rxk<����5�~7����}��~�YY��j;mg{}��Yv �����`1��;Iֈ�y\$\F=5�G,�ӥ�==P̳B�#[��"�;�`N��$j0���!���s�NF�����P������r��wJ9�*��S|�o���a���S�+��?eC^�S�+�Pa��nS:2�ƈ�ً(�; ^�6_V�]K)X�Q�����	�ӆ�^�����Nw�f�.<82C^�]F��n
xQ�l�}�6n�%���U���A��38�K)Ke2�ײ�zx�J��o)~ݚ�@�4�����+��w��S̛�i��V8���b��V����G�Y�ܵn�5���Ѫ��J�|�SY�?���Mh��o�0\5%��Ц2����J��ҀN�o�p4Gʄ❛<���U�11�T�o�<<)x��7m�yi���WU)YY]�?���:�z���2iW���4\�r�E���w�1��:w���F[�B��7�-�\�0pR���p�`�
��
t��,#,}��A��f�0�j0-së�Ft�a8忶�Bkv�\*�l��r�ϓ�8E<���
Hƨ2�X��Y��a�J0�N��=訑B���r�̀Wӟ��s����]p�6�ɶ�A�Pn8�}c��I7/��,������n���F@C����9�
]B�r�Nc����܌v��۪N��f$�\�'���*;��N}S6&�}n�s��P�~4��[��᫝��'5K-����+�S��W����h���9�G�r(��ٮ�Z�au��{kk�1on��z�{F�c���40=�(��'��b�N���xݺ�Ŝ{\�^{��^��o'���qX��^٬:N��������+��W@R����DCR���lw��C��o��)T���M���v~謹��p��\�?�u�w��>�Vc]]6d�"\��J�M.�l�%mz(�uL��G��qN�N��R0���%�)���UD}𼥵|�f��0��)���;HP%���k�2dks�E�
�銇2Ga�_1��K����{�-�Ԁ��2UBq��gDE��T��VYb�Ӊ����CXG��ig����Zi��Vg)��mrg˩X��!V{>��ʳ��Y��o�3���Ww���N*E�ߗC&�{h�X�w�[�8յ,�,h�ɳ@��1Փ���n2e�\H�[-��Xu�L�e:�d�t61��z����#I�j�w�-?J�
�:'Q�k<xY��g\����n�6�r��O�{z��pXq�RF1�Ƣ%upC 	VO�̾Qr���Aw � ��.^ל-l�V�A�xa�U���X�Q��Z%���������_�{*QX���@#j8e�B�*��jaE�/�+L	���*�j5�_RN�9��"9�N	K{z��me��FQ�=�_-x�tS��p	�a�M!H����B�o�����g��'1��{'J�7)wl�N^3���J@v��A0����[�XLҘc�=�. 綴53Ԧ2�������Wn7Y��v��X��I�-���`�=v��~�?G��DЅݙ��NW�|3^�t�xPկL��B.m3���岇����y�m�����Y�Xn�?'����\����u�`r�2��|GR����QZ��v6���D�Z��Oeӻ�:�l��U���U�}U_2te����x��qUs��%'֟�U-��v�������}��u|�3.�.fW�u,���v��5#F�MIpԇ�E06�>�]'����[t���o	���!0l�yj���x�DV>'U���Z�
a�y��M�񿁲�|��4�7/��g3����9֕��f�wP�]��ȿ�X���w����2#�u��X4W�e�#�6o�މ��;��/ :�k�Φ8�@]K_�+pu��l�a�����5����t^�}�/."\��.f�9{���<��X|@�m[�V�+�Eaپ"�����+Wq�O\��zrpQ���������]�W��W���/�
��*��5��1C�I"�iCf\�c�z��=�ŀ�a������os�b��=�����U�kQ�u����^��k什�p��p܎�oNj�c.)��^y>�g����"+����]쭟G�)X�]K�b���8n1�7�E̱����j/�7)��t�����T����G�a��_?�z}l�+I�a�kXǸ���_�L;�V� BV�J�{t�)�ݣ�l�\:-B�v�f>�>�	�0yuEV�F4g< �Ḵ�3�5��Ʃ�ñ�W�k=��,ZEb�Dތ
�Vh;�b`""Y������,�:3���꯾��7s�>�l������T���S�DwyO���O��R���e��J� ���;%�\a�0=��tޠ��׽�",_��n*�mDJ�E�ph��:�|Ӵ�g�K��}Tl�o&�V�Mp���Y(m�3��R�0�0+"H6���ƽzG[�/~��6�w���S.2+����;�8:��1�ӣ A���x�V��Z�h���˩K9rԪ�����yٛ�.E��Zs��1c���
�{�F!����F���W���C����];\ؼ��P�HfA�#5	b��գ�)�b�J V�\��c�Uf	otV*�կ'P�/���*#�/�d�iZ_&,p���l�r�m��܊�YK+N����^���g*�X�<-Է�^���P�3Q�j�}��1�ĔI5Gg�K����sj����\7Շ�_qbXnK�rX�eo�s���s��FR�����ռ���Q�+�e�"��=�U����e�u<�!F�z�".8^D�Be�B�	�X��8
Y_%�/�]՞��=�,�Ry��zY5=^���J�#�[����L�W��.���k�ł�s�ݲ�Z9��V��md#����;B=�̄�A옰��Y��z݇�gA}�\�Pʟ���9/v���}ږ⬄�����lk�1@P�-i���]︖�Ҡ糴�W{菾����}��Fm���<tS W���� ٶ��+���xg��8v�k�B�������"ճJ�������X�Jg0+x�y]额V�ބ'�~��u�e���bΡK�!�Lɛq��'E8�w�Y�f�@�n>1��2{��LF�P�Q��x�U���'��R';_:9;"�*p`/"*��P����E�|���J����7)��b�Իp�p�$�+�`�8N9R���!��C�z.q&k4��^��}iV�J�s���l	NhK�^w����=��<�<4�.5��rV)�����S�e*rLj� ����x�WHbˣw�Y�&�t.�q�pPO>���|q�s���3��U�q��Ar�=Ȫ�`�(�:��OMM�a�n��niI�Z�2{g:���Wʝw�C�{$`�i	ӛ��d#��d���ؓ]��ј��±&��˂y���k�'�5
�T6n �����#A�5V^�z3���n�J�Ru,7�WeeKd�gc���@�TOY{��\3�Jx�^��o�'���3���ŵ�� ��,�?
~V������k��ݠ�ǲ�u�g&E��r��@��o(�t��6$λ�_H�����i\o��u�&M��f��iJ�cT.���d��敀�a9Ե)��}}���Nge�KM��r��AN�st�nd�0�?b/A��݇χZ�D�.��AY�m9�mq�{^A�K�rn�1��E�S6���Yq�}r�ɨ`b���cF�jgGUg(��Ƚɢt?��s��G%V=�*���g���Q�n�+�])ey��yhô�G"~s�yc=�eK�鰆�h�<�'�L�c�̿��F��;s���c�=�C�W��yJ��7��8��Xu���`��T0/] x���L�NH�Q�8��7'bIX�B���yr��5ȋ���q���NN�g�J����V�9�gK���O;"\
M�8P�7��}��Xq}��.&,��N�Y9�W�Y�z;�A����w9��c��3i>}�Zk�������5b����v�~��1�į���@.�uf�(|$�C=��V�[���p��9��MvR?lC�!ȩ��ju�0�B��
��J���i��׹rlv>W��=,`�{�ь�,qW\:q�u�e�Wd_:�)V�`���}ݾ���䫭T��eX����Oo^�b46����_$>��}{���.��_��wKd�1�(�p�K�U���o��0u�z�s1ӭ�}�:�ڗv[��K�>"49k�w��=��{WM������	��v_[Z����I_Z|���S���ﾯ���g�9o�:��~̝E��}µ�B������/��U#B�ǵY�(���Գ\����l��.�ĕ	�8Ó����Sr�#j5�������C�"9����V�c�3M��[n�c�K��ċi�7� w�F����j�W�״�7Ut�c��U�ʗ]~B)/�٫� D_���1�cCվ�=�|h��T�w[vJ|���G�ƈA�vֆMg!�7z��^�f��YmO��`�EM�1
���M|�iѻ?d��}�������mR�79���#AQ�Y���a����'�yU���Q���b~r��Y���voR��$��*S�o��y����zC�bs���
g�U�Oga�sѠ���Gr�[cz�wr�
q�ͨ�fq�8�L�ΐ�8�o�G�[��"����7�O-j��o���|���+��c>]C�7�|�?uɓ؀5rS�3���`�O[�<��]*���\V�UQ��+�����lΩ�mpo]���4��<�V��#Dʷ�*�5���쩶����ӑw�ʘ~��i�B�{��1}6@�]A�ˮ�B�!C�O"�﮲��z�K��y�].U��3o!�R��Q4lK'�	���j}�!b���ݙ0Ǖ����7=�k\�,/{�]��j�l���`����2+�䬜���2|CpB�μ�Gt���̵�����J`���Z"�w���K��هi�VY��ᜱ��V�a�^
<�0NN�I�_-�5w�a�x�?4�����F`�%B�l�Mv�t��Kz��8�.�o۾:��ܳ�l�"�>n�
�L^˗���_u��>��j�a���[�tE��w��y����Xٗ7��Ӆ#�ŐL�{f_.�xIne
�ZZ=��f0�;'� w.�I 	e�Pԣ�\M'�o8VSnP2��)��Em4J<��ݍB�'���G5�\.ofkk6N��pHí��=(=�F\Wu�4mf�S�tA�.w��nWH�Ճ�X�3k��ͬ\��^�ܦz�/�{���0����&�J��>�x��WW���ۏ�W��w�z��֗-����e�{Vy��G
{��@�Fc���-��.����6���|���xs�D�e�U��*��O&H�:sf��U�~ԻƖN���ϻ���[D�6�����v}�+],h�]���%�q���4��ө�4��4�q�f���	��pMa�N}�A�K�s#j�_ ��,a'�x��
9�>⫕[��yj=(,�C��{�ޮl�.j�ӏ^���¤�'�WJ3@�<�%�mg�����z��.1�A[�yJ]̲�5�����AxfO�X�vț,�a��X��q��-���h�Pr�ޓM<k�LNF(��ֱ����ن��EWr��{շ*ZժL�tʚ�]m�a�dJD��g6���v��p�`U�xy�\��7���_93r�w[PF)��ӭ�4yM�7p��ZX��Xך;�q�r�V?�o��`{sB�jɞ�^���ko��[ݬ<��e�}�Rjʈ�vz��R��	�쵸�f[X+��?n��&Q>�o�J~�TM�]�3�t]�-7�L���} ǈ����?]�L<>M���`�y��|_0js� imuɶ�N�9a��W�X!i]�|n��\90��KA8A�'�a;�?��&ZY]{�dtc��|0"�K1E|7��;��b�����|�cP)weM�r�q�a�w���H��W=ӧ���P$M���oo([H���D�!��N��W����H����V���[ui.���Yr�r��'NY-u����$�(e��ܖ+;�zpn����at�Rn2��z)U���oD� `�혞��W>�������s�*���UJ����Q\���G***T9s�J����QW8A�gI�E�؇�
 ��Eh�!E�B�I��PqQ���\�Q���2�C���Ȳ�:DȈ�ʏk2��2�
���j˚&IJ�Q�bQr"Q5�.�2�r�d�$�rI-�*���)g;)����V��Y��!DWQ5J��A�Q�B�N2�a��beZ�8,��V����@��G �^RD���Z�T*�9:�"�^"إ�YUĚBY!Q�V���$QQ�R��s�Au@��t�9�֕RV\���Ch��r2��+ȕp�PG:�b,Ȣ�TV\���0�"�\���2+�x�,�t�fD\��TJ�Q�d'J&QErr�U˒�E��ESR"�ǜ��h��p�.[q�g��(	mR�O0����l.h�r�U0�8�#�e�s�TQA�@���@������[z7�z1��`k�h�;�o�A4�Q��o`S�,�{�>�����oSip;� 'C�h�\��7�D�V9ꯪ����]-o8?{����8h>h���#�T�W1s����F(��u�4�;���W&o��N18��M��k��y�q�OW�,vO+��u������\Fo�o��6'{	��_Cu�e.o.1��)��X��~bB���ǮV�:�/Þ5��w����}es�R�8�{��5ҟZ���W�}b�}��-��r�5#ザ;njӪ)r��ή]��>�M텓;T�q�B�w-��UT�:;k�Ъ�>��&��Mw58��㦩�|̌55��N*F��<g*�ޞ���������HT�R�:��'�7����]MZ���p)���暝�+���	�͇t��9r�5_�������0#��RZWgn����r��.��P�慐�C�u|8�D{��J��zì��t$�-R�Vr���U�\Y��5��ej6ٲ�:�;җ�'�E\+6��ҥ	����^���ﶮu �VU'J�`^��z�5׋�^�K�R���e��Mi��� 9��߬�=R�S�n�"a�u�%���6��2����Д�r�E㡹���.Ro�X9�mf*�MG�����q��^��uS=�������TDD}]u�[M<iFU��7�q��vǏn���
����8n���I�i����Xn�(PN�9vSڈ4��1W���VR�A}z�hH��O��V�f&~�}W5{=�h��W���.��{n%i�9�b�G����^_W�gi���������#��8��ޫ�y�X���w-.l����_u�.1��]�^�;�ϓÕ�<;��^U�!L�:o�8�%��;+�g*���5�Mꉊ�oeS����Ἓ�ݘȑ�/	��CމG�ne�b����uK�v�x��Qm>܊y�	�ٮ��8��vN�e��,G�{�u.ϐ��\1Pb�����wJ���Mn��Au/�eùw��a�r��G-����>N�,�UO���{}>Νo�&��lڞF5��c��d��_����3�@��nT�i�)D����5���Ykt܍��0�r����{�l�鞘)F��76�ig���b����%����ЎƦv�M[N<��owD�zLۉ��<���*��ͤ�Vu_&��6:��$W�w;9@�d��������ˎQ.fĮ�_\'d�nŎ�ު���S6~������l�N�g�#S}�4��n�����麳�*��q�����)ws����W�W�K������z����r��&Қ�9r�>�	\���NN�9�Iݶl����W�\�uj�n��!檈yd�j�q�Aڨ�թҍW0�ݍX#�lM���ٖ�k�Em+�l��'��p���کv�>*%۳1�.b��>ۈson3΋y'U|r�_!����!Wy��k�fzn��C�3=��~��<���fz3��ZR����6���v�ίϧy��_���e3}\�>��3���<�uT9}��o��R�tl�	�x��3�E�yލl��]2�Qщ��Nq�Ў���e�A�ߍ�<�u%��.�5�
Fywb�qr�!w�Y�*v��v�Z�V2���n�˜Ujr�1F:�?_(��v�dB{������Hګ:�Ѡ}�xjɐk�و�������P�P�'g,3b�22PY�=�����.�Ÿtô��4������O��nfz��m��"C$��K��<]d�\��K�NS1��/�qQYq�M{�{@Q}�ﾈ��*Ufo�[<���X]CH6G��s�]�B��<��U��|�.]�a=��g5���^��K���Y�+�/0u�K��/�U�Ue��͗Y'�e���@��9��I�Ȧ�*�O�b����ߧZA��+��tE��>}/�N]������7�Ujڝg����B��N�B�;B�QO�?�s"b��y+�5ꡫ��h}�V�v�u����ؚ�N��Xc�\���f�n����<�����u��(�ķ;���n1YЦd��9ȱ��$ܞ}v;�}1[���}�hD�դCp�����,��n3F�{,���O\G�5P�Ng���j�$j����]T�ȧ3��h^��N��P�)����,Ĕ���~�%nO*/��[M���	�1oTu8�৖Ҵ\=��:�;�Wnb�=��f�L�%��LH��{T��s¢��χQ�����&�e�Y���t�h���&+"�ˮ�ov�q(�y�_:"��a�ͱ��`��v�ޫiV�ٷ*V=��W�АPs0�V�rP�w�^֙��(o`�:�E1�ڠ;0!WV��v�>1Y�c/�m�n�H��Z2�RWK҆	�����}����Ե@���?bΚ՜B���*�8|�s95��'fT�{�F���w��ROP�>�F:*�¥ޙ�~S/Չ�ڈNq��o�f3����b���IF��?8��[���y���r��^~������^���0�V]/���N�-{Ý��y�~�M�m�����\t��@�]X�T^�����=��4w.+:�=I�O�^AO�����r�.�禠�V�1��n=X��»n����<�������r���76���8��V�]�z��[C���;���Q�e|���ƚ܊y��-ׇ���%qJ1�:����w]�ozkn�9�4�TE�V>�T�����kZ����:�NmPݮr�R�W��(�k^�.��njN�LE>U���ƫT5v\-�2a�'�FK���\�
�¶�hU_�ie(��jo�]?S�/
�Zs�(�����6��4h�t���2��A�7<�o�{�+��Է^^hO�����ӏ�W�<�ړ7��Mc�Ϛ⠰l�U�r|0�9x�+u�ǉ�_V�L��^nT��eT���\w>���&�L£�y@ilќ�;��W�}��UI�x|b��ֵ���v�ܸm9n�w9W���XD�ǟ]�\�MX!��>S��-��f��߫�&�y0�����)���U��5i��g/��SS{}9�sS4��%]Σ}����g4sy�yeYSCY�b��:��]*0^��lJ�	f\s�ï��5�-���[uޕʣof�P��R>d����rS�-�O.�﫰�,{s!N�5���-&�\���i�w!��7��J�ߍ,���QoN,�ﳨ'0��
�
'm�����=�D���i���'u��pu�D^b��{Q��*;y�r�w
��*�-��W����
��;O�l��ˋB�Ϫ�����&'���c~~���c�~�3�=�ץ����lײ�Hh�o���w�q�%l�K�}-�����5�Oת&�[�����q��xw!���Z�=���dH�Т3-��dP���+n]��פ��X̿ �����(��6��Mf5d�.1��h]�;d�-����A�{kA�Gk�<�Gq���Pk�J3�+�J��)�OԈ���fGہ�;�
�O�D�|���C��Q\�D=��#�舳�5_Jm)7~����U�\ⱏcr��{q�ث�����6i|D��E6;Sݚ}�\n欰�]cTMA�֪�+�}�*���Wf���][�-�Y�\��Iu}�����\U�nv�c�����:x�|9��;6E��%횗���}�vCx)V�X���;��mDN��K�L�� �x^_t�M���}�b)b��.��<�Rq��q���P��k��˧3O�Qr��W�e����U)}ܘ\�iܯ���*'�aTWKɒ�j�%��0,W&�>�]u�bs�n��N�3�:��=Z�'7�Ҫ5��G#���j�ƭ��ek��.��^������Y;�g^,��R���s��*��a��y_^�+�q<��+8w/p����"ˌIDv�N�eCۅ9���v��/������[�<$���u�����%Z�DʛR���
��u���LD�R�\�<�;��#ѕsQ9������ۧK{wp�ԨL��t��.u��W̙�1�Y��P�ֻIkyZ�˹^�gܼH�v��s޼d-C���/�W�UUFy�t�Y{��ws�;�B�N�3��G"b9�2���4��b�J�b��m'3�	@��R���g��u�!EF&6�9�q\ݧ�o�t��{��z�|�\d�`U����uD^NV7��T���%*��)��0���MS�7�<��gVq�R�_.
����7��[T����԰ά��>v�d]�^��v�n*1y�xq�����҈=��f���;Q��D/o˩v�y�N-B�a�����8�o#���1V�s���䯸��W�Q����ڼǏVS�����̚�zV����"�૮���J
����'a�Q�0N�}qc1Z|v6�J�p�}�U}gܵR�����k������7�+SJ;��[�R\��$�Ӕ����ҳzw�$��Hk��yE~��`�G\���#Ф�wmZ�C����P���S(��MM�.��I4�C�܇u1N_�aΈ�ڌ��\Y���!u,X,�{�GU�#ﳞxN�g(���ڐ��z���{<�`ߢ�F��ӄ�+lV�����b 
���c��(J��}E�N�᭶�9�D>u;k���N�:�K��ܒ�GJ���"��V�������9t/D�%� �J��S��	T������5K�;J���g$s|®�2�5j���8Jaݙ���V�5Xc��P���9�\2�5qg�bL�#~כNv���1��*��bU�zeØ{Wc'�j�&T8�w�]���s윗�n�W<�于�p��/!>��T�*W���ݶ໣�p=�$���U��E=	kx��1��jɈ�
s�������p�G�4�$�ٗH^�sI)�q����y�ዕ��J�ϝ)ޫ��u)�}p`On'V��3.���g��t���;�y���b��mV�,��T��6�g5�v���eOTk��NGe|W�>}��uj�l�[�e��ڣ��Fo�nC��n.5�q����/p[mOoT�������u�.gKf�?;���]�r���g<^�<�~Bo}�J�����e�0XB����̂e�uϲ*C�iR�|/���&m:Zs
�a�x�0��Ʌ�'l���s�v��j��+;��-��VP^T�ѹ��0\\�F���
̂��QN�s��l>6�����a�2p͖��Y�Ms7!!Sv.���r�����s]�&�'k۵�gD_G-
�7{����z�[X��'��t%U���.�F'\�;��1Z�Y�V_;�T��jym��"��r�I�0�1oB�ď,�q��|?�mvJN�mG���=ޟgNc;n��]т.��Wmjs�v��-cw�)c.�8[_IДOsS}�{���X��)�׏N[��|����N���+��Q�6$��y���j���=ӉTm��g�ί����A}ԛ����wJiK�K��K�@���R��z��s@�+v��ˀ�n��S���掿��u�ZW쭱��0:�JyG�'S���������o2�+�Fr�X)�_ꓱ��D��;�q��S��y��S���ƞTE�u�m[�U�r��f���]�M/^B�ym�׸wT�������}<}�nz27��K���\�*]�Wңx ڮ�TZ�^��Я;:�(�i�@��x���P٣;1�1�xmu�����f>�b͜%:���]����C��3]���?.X�!M����:��,�2��S>��wX��j+X��+6��tnc�ͩ��;�zm���p�`5��ϧ|H��!l;c6�l�)���}�J��Ԁ=4ᑑ�T�i���M����e������:�h���n�O�em�䫘���ow#���N0nn2��{wq:�-�c���uo ;y�CD�&�����J��5v��o�8첥�{P=L�#���hnR{�,�"m1q�����lB�q#ȱ�X��T�q��{1)�r:���Dڭt�āəi̠�Y�&�5a��i��4Rԗn���T��Y0�^�,�:�����h�qwv:foM�҇�c�+{TT��׆��c@��`�uoAzK����qM��������z�c����f������k3��y��o���9�*j��1��wD}"�}:�𷀅Z��e��w�t���,��sA��h�C������ÿ%��y��"��c��׮N����q�{N;瑎�p�c��+;��ugy��_u��}`�5�D��X�^焮qT��G�GKʆ���ɹ1�)�
�61]���4����LZ!D�?_sh��������o�E{��-<ּ�ح5$3��'�y�^�xa�9���$�
Ա${I��>C��{�P߻�\��/H55�;7]O2�P鲭��ݔt *���&�Yl����{Yҭ�ګܪd��Ns̗�D����;��i���y�v'��I���i��c^�~��
���4h�M�^�$�:�
�q�ݻ��Vd}xz�O����M��KD�͙Պ�ӎ��"omc1,���7����W��6�;��~�+�K��ޒ֎^�d��Μ�l|�kɕԔ��������`㢗^C�����z[�%:�;.^���ђ͍Ϻr��hO�1�����Ɯ��!&㙹��g����I^���QM|��.�R��P
����m'�I:L]��L==�B9��7����]uNm�/�����G���۴M*�rL�n���M���w�v
��0 9�sqC �WVʌ�2��asmu�Jq����}v2n<�N�srȇ82)f���K
Z������=��\s!�J�)U�O���BJ��)�W��~L��u;|#@7G9�6Dᷰ���>Ջ ��9wk���i�yH�x����m�63Ћ��v���1�s:)6.�"ݮZ�W7k�����C8��0f� "B��k��>�;Л"Qұ�*"�nu�b�Yv�$+�m��8a����\��D&���y��,��<.�<n�XO�S{P�f��(|����B����z�a|��\�ܝ� ��O3]�M�zT���eՑQs�J���rAwWM�K��ۏnP��l�xr��R��y���$�S�4ؔΉ	�/�aZ��[&��� 
�TŲ��eW*(���r("�s�I� �3���B�[4,X�Dl2%i�AgB��r)E��jTQ$�S$����TA�V�H%��D!$$�ÊA(�
�QE�
"�� ����ND'(TG�˔AJ2JB��"�YQ(���
#�s3U�"��PJ���$#P*"�I"�r9ʪ�R��p�APRt*N�.r�(�kN�DDU3�]2�#��QW(��UTTr(�!%H�(��J�*�U�:*�&�\�J��"�4'.9ES�����PD�JUr��TDQ�IDA�UUVg.\�2��Df�
���!YaDG9UE�LE�B,��J��\����\��EZ�QU�$Q���8��[dgB("��R���d�@DB�) B�,$Ñ�R��T�eʪ�B9 ������&&�+��$�V�Z�j[P������y].4�;�+ӽ�ӰVt	و�&œFTW.f!;�b4v�zr�%�w�������]u�o.���Y%մ�s�!"~����ۈ:����W����L��X��i�ͺ�Cu��HqX�ڄ�s�z�ml9��v��R�3���B�6y�>N�JȀ�yә�(讥�������׺m�eG<;�[";�z���t�gj�'�M�Խ����Օ���=�S��f����/���s�\�!��9+�%\��*�8�#r��sb�-�ꃐ�QyOwl�˓���|��BO�!�j�%p��C_�h��G�����"2Wvt��M��:�����[���U����(*�*j�D���)�Y��K�U�k��r�CS�zm�oh��Wt����Ut-��j^}J�ҙ�;�MojVa��;
���.�t�uz5�ݝ����r�θ7wMʕ��-M�ƞn���Yʉ�hw!�o�\F.��ԋ�Ln�`���jޞ���3�\���$�:ne���nO���*�3��܉:<C�\a�$d��v1=���KL�L���6���ْ'Ě�,'}J�s�цsHr�8�q����]خຳ�u�Ӳ�a>�/sq��j��8�G�1�ﾪ��3�ִ[ԪmK�0s��M���.˼Nc/J���/4#�]��0�c5F��Lt��u�LL'�BY�bV���|����>�k�EIR�#ʦ�x��9쭡+���"m�E���7�T�=��"�����O9j����Z�I�u
^@��p&
���4���w�㧻Wy�f�`%L�8��e�}l�W�����VO7���-��^���T��P�U�^;ǵ���s�(�1�����[Tm�ʈ��n�`��r;6�gL^�+��0���7�=ؽF���%q��릤}��.���A��mm{.-��Sh��>t����x�1 ��ͬ����vA_�'8~����sn{��qU�}s���:��[���h�ڛ<����ͮ��VV��LU�Z��cü�V^`�w})�M�G9oq�X������A����0	�`��qq+�X�;yt��b �i�,\C�d�ç��tŎ���:��xm�S�ɹ��<��|cx�X���u	ư꺻�$Y2F�2��po��p����f	�9��z�[��5�e���')?}UUUg�p�X���ע�'wJ����7���X�!��`���H՚��2TV����Ճ2�j�ues��V�jyoy�Ȧ��*�_q�˓���U�)�R0N8��;n&��q1O������WIf��z�^�r3�α��I.�UT0n��2�����I�)D�W&��un-�I�/�Վ=X -�6�٬�<1[�8d����	E�X�M�}X;�|B��!���V�H㍤�c6�\4����YVT��`�Y�`�+^>���Oe�D��vwH���9����U)�H[��*yfc�{+D��ײ���F���g��^q+QVU_BPNd��[����9崭o��q��k�S�9���Y3������yGW�5#I[��C��~|������n��S�3�����~�%�Zh�V��j�=�)Ԯ�.��^31���O�U�Hh�~S�<%��˙�U�y�&�;�-^q{ՔZ]�ż�A9 =�!��omNn�MYAh���=dlV{@e5��Jrٛ�}	C�H�ifMf�M��P�<�����w����@w��h1Z�dє��'��Q�|{Z�
㵚�B��b�_N���a��)I�����*���������s�p���J��O���2���bߗ~������U�G�Ĝ�r����Ϻq����QN���n-���|�J�ce;��ב;�.9�*{&8�)WE}ܱƵ��,�Ǉ+�ۂ��[o&����cz�_֕V8�_iyW����[��ڨ��Q��Z6���zDYع옚F�,��}cێZ�.o/kr)��5�gzj��qs�Q�̧k�k�%�hu��֪�*���q�Tjw�ZmJ����l��i���Ҁ���q�������Ύ��*�����h��tLՇ�	���kUg8�m��*n:�Ĵ*��-�5?�b����Z$遇uR}�k��4�4��J�Ƽ���C��r�G(���&���Wc'fTR������2j�@�Wx�kuR��'���T�\��\|�J�`��4�ʾ˻��]%L��E,���6h�^��ni�H8��D�m�GZ��Ð�囔L.����Տ�n�Z}Z\1�ኟfRYmU�u'�e��>�я����z��nƶ��˭5���Q%R����}���]�TX��G�����2�}��esy�mf�Aܛ�ۻ�Ml�糫�R���y���VsH�y#�����1�i_��f*|���R������\TK�w�nb��>�v���v!�����/��)>�^<q�٣�~m=�6�󄰽�+���=8_m|iu}y�O��\�J���s��p��{�1FşR���Z�K"�U��G�.Ӳ6��B�cޤ�޼�ՂS�l��Q=)֩*1��\�ߛ�Ρ��Ge҉Ó�XХ��un#9������֨?WR��n1��^Hmw�Fw���t0�s�`��V�P�]���K�y��k�T���]�Ք�{��4;i^�<��Ņ�4�{DcOf��o����z_{­�쉔ԱQQ�O�yNW,eHb�?17��w+0u�5+Z������Ii�Q�YI�����ƈd#�{~��jyd��D�����ޏeװ�m����X��~!�2ʃ/[T��T��W\5�cb�f�P�F��#�"J��YC�RX�34�(�pTus\�1{G4h�M6��-������/�\����o�舀iovuNM���᫮� ��}0Wv_��}xĪ*�&b���LK#iU�ע̵�1�����������W˅���uA([W����{U��{yp�VcT_d8�mM�.����r�Zo>�C��w�����J�M�2`ˈ����o�E�yq��/J���1���ǳUyMԲ Խ߽*v�x�~B��[rnJ}we�}��
��:��eJ���Ni�.��^����U�r�MCU�9m�ؕ�����+*ft�����N�t���ɣ��:��L�AwP�����Gk�'��J���j��9��++<�ʎft���1��*W�{jr|���;s��e��Yx�F��ۻA4������:�3�*ݜi8�6��:e�B_��^�}�Ȋ2�~���դ�Pض�OJ�i󱋽�M�j�}K�i��xozM���Ӎ��H%��K�*58W/4g:�vH>�����	��+M�XJ�x�$ϕ���:,%ў�49&�
t�|���pN�R�? �U���RϠ��Q�p��Vg'�����l2��� u����+��t�԰-˞�l�����.�j�\���>|C�#���-;�p6�H��>����r��_j��ݤ�\S�u�F�����RU�.�u�7����5��|�e��B����o��+c����n�v1���Z�V#�k��5�A��=��4=ECY�(��<�O�x�dK����>����b�[��1K����}��o^`J����]��l^e���h�-�(��R�/��i[K��ƚܦ����Om�z;i]��Cv��Zf��='�ݚ�Ǉԝ^�}󃧋��PN�_WN�E���v�
�n �vP�l��]�׏ԣ�����;�"�%y+�5ꡫ��h}���������SM�c8.�����@jܚ��O�\��]�[�3�Ʋ���{h���u��������ݵc����tXԶM�A��as���~�' ��HŜ�>��熜F�T^�N�%�U<��~5�uf���Բ���:��J���U�{K�`ĲW-��t�z� dWқhQ�\D&tPT1kp�m��]�>Q�7]Gw6��a�x�<mݭ�gr��	�*�oIC��#Uvқ�
��苛�%MP{���x�b��>���5��ﾰ�}�K�L�F��Lv�S���;���w+)bKP�@��B���b�T��^���i�g��ɬKvdG0�ҸE�ۂ�9:��teS��s��ڒ{:Q�L8;��������8�ΫȮ����N��'U����:�][Z�İ\>k���D�i<����R�d��|���$X�w;�N��z�kF�����J�|���ե���Z���U�����o�iy��Ľ�����b�hl�nD��\�r;*q>|�����HΗ�~v;ԽK�O�V����)��/��y�<�dz����	S'�w��s3�l��{�<jR����el���'+�-^�y���/��p�*W5��I�js*���}g[�UVW˛�ƚܧ��s����`8��K5���W���A�}�J�*�u�MEk�D�=<X�j{��oS���,` ���F�L3��y`q޾WW���t�ʄ��3݇Ɲ��<N-��5)�aq�|v쵋�
���+K+�<����4�h�ft5(9�l{���6_N��,���]^�>z]Z�S�P�[�����]N7�q\��*������E\��UW̑��Λ�욺~��zh�����^1*�P��w���)5G$5����)��,���<9���5. �ܿ�.��5���N�a[kB�j;(����Y6�8�S�Y}Nd�*ܓ;/�Rǿ4�|;s�z2~N���+�%C:ɹ{���]�-5Dgu1�^.��Ҫ54��
���|�yr��<6l�בmӋˤ��ٽ(�څo���0���2�'۫J�����&�l��M9�d��J���M��j�{q6%n^@O2dkc�u���o1�-	�����%��̇O���1Pzۇ6�,=���Ƿ��Z�	�;+3�{!S��o�L��]�\)�t��:sӵ/��,���oL����9�VZb�{u�Ǩ��]��w's�'�Lm̾�:�ꓭNθT��sי;ДN!����81�M�j��1�����f�5��f��7˲�`�>�+�<�q�re\���$���z$}�:��EypJ����y��z�
�csd�(���V�ix	���YJ��nHo& u�MD&V;z���;u���.P�j���`��p3h��s�-�4	�Y���Kp�/HY=8��^��>���x�y�ȫ�j��ߊſ|��6�R3z��^�N>ڥ�lo[*�XK[��vk����ޞ����и�|qC�u/?QT_VV�>y����<�69�n�U���3Q��j9a�~&���{�^��;X��2��ck�<a�X7`kGj'pv'�{�,�kg�3U,f.������^�w\�c�q��2o��N��w�i�Ȧ����L>�
ү���O{K{����!n-�xa�oU���U���~zm�&v�g(ЯS���T��2���p���v੡W���e.JqwS�_]ִ>ۇ�'�鸓1='��,N���k��|�#V��	BP�d�J.)kw�~���p_u&5����1hkJy]�,����!�"�9�;��d@��ƥ�I�)�����+ug �^dc�u�YUx�����g�r�)�j��-��y�ƽ	��F��Dc����ʍ�[�Ҁ�jץ"2.;�T�S���������b3&��Em�C��`��r9���b�����R�S�����Vv?)bI�\cW����ڋ.��
:���������{ٹ��6_�i�ah���6��v���L�}�dUGIk��n�HMʒ�~&q0QәZ��3�;�����"x��\�|�Ĳݭo4e,��d
l�V6c�"9y�Ztv���LN/^=R���nf��kz҉�{P��=I�Ts���XU��uݓ�'�"DAA��IXr��L�ѡI��ۍ*À�@C�c��૭Q���.�X����A��=/s���e%4�0�lc���ݧ���eNH}�K҄�w٘K����S#�r㲢����+m������Y�3��}�58e{{����̓����T��J�,��O���X(op�[�ň�T{�!�*T�-�������2�X��
�@D��{�
�,�Jo�ky�C`�RZo�CInt�}�=�(��v�x*H�Fr�K#��l�O�C�(�iѿ�V�^�t�֑>��l�9�j���"���KW�j���x��o�U6s4�ݙ,nS�Vy5�W_d��|>�X�wjW�l �&N�F�*��;��H�^��z���{��*�-��pS�SN�-�fv��E���cwL�'5�O�y%H���b�]5�v[�k='t�#��Y<u�7��{*���a�읶*�*��wND�H�a~�.c����]]"�mJ�4�ls����o���n3�O���R�rx4�
�\w��W3�rb����$�lWQ>�(��V1��`Ŭ�j%F�C2�ź�#��nt�{�w�r��8tn�2[i�.��ꙗ��*̚�m̡]9Xz�Vu�\�$,�V�]�+f�
͑�NF�e�v��z�7��M>Q�pLҴ�V_0�,��eZ�͇���Z�RԘ<8Xz�VgD��b��ّϟ(%�xg#�0P�}�9c�RD�)K���E��1f_s���.{���
f���#R�:bW
��ޒ�i���\U�6_��0�O���aC����n���7|����H�����D�N�n��RV-��M8�Ƞ$��bb���g���J�ǘ���/�V/�e��md�����؆��$�&ptaYk�D��uwZ)Ww����m娔j�;r����;f���å���+�б�D�4�[�d�[CHOO5��K웗Q�G8F�S1B=���u2�S�Y5<�Q����垕9��[,�0ON����֑��#���ӗH=�[�|�Ah�%�7M���M�ǭј�������p|sa4.�T����pw�nR���4`���$8�Z���ԝXj��s�>(�s�WֲS{���rM�U{��޳� �&�n�`�Y��5e�:o��d�M�#�>��:k���e�4��_�6��h�(P��
�Ej��E��t3L9��-B���UP\�P�B˅�)R吵XDh� �r9\�T2H*�����9p���I""9���""��EU�t"��*��EUAL�H�(�S�P�E��ZЪ�:m�D-aYЊ��$�(9�<\�S9Q
(��9x����PJ��ӥp�\�Z\��p�,HI9#��*�UQr��DsYi�K#�(��U���J!2���T�e��Y9��� �N��(#�DEUȊ�V�Uh��QZ�aF� ��*L�k:m2�"�C:H*�Qr��4��Y%U�3T!�W;��Q&����GR��q9E�iʮ��I,L�--(���%j(�s��]5*��j��EQ����s�������_$[�d��!�r��h�}�{���O���k4Ƿ6�c����d�ͮ�*gK���K42�.IG,���|>r%�՝[޳^Ǜ��(��-G'F2�T5�]��C��R<�]٧Z�Ub����R�un�V}��:W�{p�!�7��+~Ѻɚ.�� ˳�K	z>����ͫ�3��kɎ���K�N/���C��+���NS�@ܸs�nvWט���}�A��#��gHQ_bcnѲvC��3�D�'���a�W5�츴.:|�Եn���_՝E����]^����L��jN�����L��T��G���S�l��eſ�N(|
�Լ��V�4�Ht=��5�q�O��Ԣ��}����h=�A��i���Q��V���	�	�3��(�p���������19��^`蹭�15�Qn��%��H��u�����r�+io3Zor)0�V|���]s�q��\���-�T���r2�K��3�U�V>�j�jx��j�o��M�V{�**oVZ�~Iho>�%�c�5'���Ѯ�K�c��J}y��8;o�����s^b��������ޤ�ݵ�Ob�d<�f�s���;9�R*��	(],��E]9/ay�G{񊳰�Y��f��� �y�z����S�k���eW��ڄ�����(�ʢ�m}��������	�3T����,�{��&5s�[G���R���(j;(���Sq���tF�{�Dm׉Z\��qx�>�Cѓ�J�<r�`J�[I�<�����:�iy^��,,��ޮ~�V�hX�k�uuǊ�a�FKf��̋��P�Н�����]n�j���v�Geo��p��yG"˟���Щ��{"���z):�T�S��7��%�7]�x4�Q�N	�-���<Mt���n�;�� փ#�T�-�����9�Փ�}�z�CM�^��ϩ�v���uH@+�eOga��g�[TR�+�+�]*�p�J�f)��>A.������a=Nrn���/��}���;�qSTٞ<J;~mq�ͺ�u��N8�hM�����G�]{.-�.1�u�]��	/��F�����W-�2ڛ��Ɵ]��7un�#3�w �cm�8mn(s���w���vǴ]���	z��=�:3�6�W��;�{V)�]f����Q�x�����('->�o(�7�2���Mу�I��G�U:�I���_��p�*(4秮�,�R�)�>��z����[�'>�4�US���z��A?/�7�ջ�Lǎ�R���-���v�c�yͩ��J�GI��w���}K���9�Į�f�����;jL�j{��{���|�K[�ڴ���w/�r�K#`���C��1Z�E�Ue�<���;w�NL�&Q���yɮ����ˈ]�u���-����Vo�r�U��t��h�^�莚��o[���nn��M�|U�W�լ�����m���J�٣ݞ3#�0��yM�駎����>�p�d�M��r�%=O���e޲dek��i�)?R-Q��>�IWڞg>^ݕ�����͗t�E|���	�j��J9T���`�\|���/���ꨂ���oD�h�f0:kί�<Y��Op��Q�����|�5P0sۛ�.��K��dt��:M�,��N4�i�Lv�H,w�\��ںf���8�[����9�P	ۚ�k�Q ���y���F�[� R����>>9*c=+���e��u;�f�jٳsw�A��V�r	����'#̈́؜�}zqݱy����^�����+� z3θ�hv�eh��n!ͽ��b��bǢvifnC�!�	ڍ�O��g[�.�}s��>�9
�g�!��8ʢ�9�W��*���'�WGd>�&�Ay��.�_}����8и~�f{=6I���t�'?=�ɧ�GQ�A��Pb{���).*#;f�s�c/@u��и#^C͇��{�n�������<��R�1�>��z��O/S�[�n⪒�],����g����mY��9�h��zW�������7��6�e^I�^�(T�˖��R���-s\����4<��Y�.����:���PSA�o��'՛'��o����~��&��;�J�͡U�ݗlڰ�����H�8�X�M;<�����֛�Cy��qG�����=uo��W�F�N�bپ�]d8�n��w�TO��Л�*�\q����^�W�Pͩ:T��G�tN��m=��[��x0�&M��g)��(��ţE��WF檮 �NF�n�Yϼ�nf�I{H���2j��g'dܩ
�ў��p�b�]\�4O���j˾ыz��脽�z�/
;z��]�z�辛�wI�d�3�#v��-��w58������ܡ���v^>�p��,��qJ��B��p�؎r�DHJ6��b��[��j*�|�5���JԹ��(b��m�)�N\���	P���`8;К����z����:�[�1�Ɩ|����aAn\@��踕�6`D�9�oS���}O+�����ڂ�Z��l��N�|�\���p���@sX�����ꛆ�u�5��aW�y�Z\= 7�y;3�&\�ù���{W�ru�᧶�Oh�K���s�)��d����֦qڽ��21���[L�V6�j��@ʯ�Wh�uv��wڴ�O�]�t�a�S����#gPUۍ��Tg�����j�k�qZ�G˴�[I=5���Z�j��l.�a���n_8Μ��sW��
�궷�qm�~8��"����WzZo�lj�_MJHk�U�/lU�)e흩Ղ����d�G����t��!U3
���=���l�Ή4�����F��+Y��,��_N�%�p�ð)u�W�.�ڙd^���>ʣ/o�k�ʹpF���}[�O��� �D=Z�[=O6|������_Ԕd�-tr�	⯣3Q��y=�����u�^��:��]�,�Or �)Tc�Z֨��NSͨO;o�zye��۴z��pc�����s5������ά�Zo˛��3�kq����55��0���ԧ�9�9�9	uU�njӭTX��GO>ޖ����tٌ�E��՛�su�]����[p��E([sPe(�s����{�>�8�/���X��s=I�z�'}��=���*t�U`�����Z�vA680e�qbs����!���|��Ҩz7z�hɇt�Yl��51{������Tһ��%���S�]2�U���	F8�P��¹S��5�E;����A�)�<�no��w���D�<�֊�4���o!T<��
�<�n]u-뮰]�/��rهc]#)X��9���W�>Y)|����j�����[X�,6�������U��3Z���q�>�!�_`��,��*S�䄫����|���m�j����1�pޓ�$T�q�9��"�>�ש��P��h��޹3�-��¯�;鮙�Њ����nޣ��m��6���g)GZUi6�{ꉽ9��D���;�J��FqI_eo���ٴ�)�ǫyD��/)�|�v^�w�r���Խ]�S)���O��ʛ���%�]��fq`4�*�,����*j���Q���Nq�#��?zˏO���l^c�����_Y��o{����OS_u'q�V���Y�	Ș���5��d+/�:T҃�U7�w�5 .��su���(�Q��R��x�߹��������e�9�׃����)7n �^;�U��;{;����GR���m�n�Ou�O��⥁�w��7/9���uĬ��Uqێ]VTB��nt��!��o�����z�c��6�,[q�Ou�!(*C��ֵc�ŗ���/c<�뤱���e[�ܻ\Rsi^��g[�]pT-��1;СN㝭h*��FZ���k�J1m���c�*۱�V�д*��`�s��4hġtn�Ħ�h�u"Y�!��E���,�e9�2(i�eoi�e�˳a�$�������Q�8��I���kG-:9qC���C��A���.Q]�j$�z��\�JMa����~�s��<}@�c�.����e��f���tL��'��c}S3g�:�\U��g�Ի�)㦚V�	vF��r�@=n�<���d�]+6oq,恀ad^�50[���b��P��\'�����վ�-݉&�X�;�tr����Fj�ZE���u�&��PZکՓ��U5�Z�Z����5��eeB(����!=��~���<�
�N=F �[�Pv;S�Dk�U��f���:���Wn`t.�son1_�b	*d������ί{�o��S��?f���'����:��N����F�u�S�T%$�Ч������;�������:B��d���o3oQȝp;<*S�����h�^�2z�n�|=�J�W�k�נ�(=��Ϊ-����zf����J�vk�/�z��>��k��u�oU����j�Ԣ��x���q��<�<����S�;�$7��9�.�>8���Ϋ}U�1�k��h67 V��y�Ǝ��Z����yu"��h�vp�>PM���*��w���d����^���.�)K��`t]�\)�C ��Vf��&ノbfI��m�ݎ=��b�&iğ�Ҧ�e��x=�ڸ��o'>�(�nr߉��\��*�8Й㉓|C9�u���SY�ɩ���{�YU�9�<S��.f���G��&�͡��s�h�EV9Ҕ�J��g=)TE��B][���[�M��k7��+�*�u�U>Ǫ��_�Q-���VW;�Y5S�p�)5����,��+Ms�����|P�|���	B�Y�+;�>�=�it����s�5(1Ȧ�,�����+�ijC����ᄨ5nMLAJ&��q�~�ҏ�STr@ܽ�R՞ș�q��8���'*^]*�\�~�pw�?_Dw�e)(���>�{��]��f��nٽp��P��J�aW��ά�vE{ɪ)�	�>}��6e�s���ՙa\��QҺ��cf�/!TC�bK�	d��멅=IIɶ�u������5����\�H[�V���7k��Y�F]�w<#�bZ<��O��w�����Y��_f�L�0q༘�1�҅�&��c0z��y�;43�>���R��O�7��&�ȷU_ݭ�g^��ז�+vz7k����8���b����]�5N��p��Zl"�yZ{I�}Y��_7�ɝ&�y�څvdi�;G%t��Cy�њ:̱~�.�'r�jS��-�/1ս3��kɌ�E<��p:p�9��GsD�ޓ�=�@�6Gf׳ё�[�K��=|�b�d���Y�P��ayk�7�c�t�P�jq�8j�����죊��*��s�,���j�s�4��7��ds�q{�˼�~Vrw�6j����)��ãO<ɥ�-O;�>��Բ��͞>��Myxj�g�l�QS�����}�G��yf{��r�<]�S[E�gռ������kg�P��'�2���vH��|��Z�XĻ��U��Ue�+isy�>�M�`�˙����x���<�j�-q�J���3Z�<��+�ƫT5<��֞��4�-	ޭnzqs�l�ZS��]�6�W=�C����DG��5M�Y�Z�}��U��R�k��=�z����v�0�U�[rh%V��ݑ�e����8g���]xT��Ə"��Fr"d�M�7�}k+�*/�g�i:"Ț�{�Og#���o.��M�<K�̮{5�`{#��dN<�d-�ZNi�ݙ�d	:kE��3�~���]�LnW-�]�,��hk}�D�������.�:�7�����;\��9iY�K���[o6yҿS=��~���w��@���#�(�����ؕ)����l_^�Z׼�n%-o0OQ�WN��9B�e�!qv���.f�fn�yٲ�ow�[A�E1�x�,�%A�a��R�/����A{=�/t��H���Fҙ̶�}��*l�I�ϫm�os���(�AYڬ�;���~���P[���#�fa����.��n^��|��}���>��
���o)`E�-#&HhGu)A�e\�>Ӈ7_�wփX�}x�Տyx�ݗk�b�&9�%��W���h}�Ȅn��¢���n�V���Y,��o&Cۺid��G�Q���8h�־�^�I�_j���|n�N���{��W�)7^j[;���:�)e譱lZ��zs�yc��!�m[gC�GT�0֣�ǗV~ǔ��"���Gy��t�w;*[�w���q���N�JY����%md���=��|@��rZH�ν'k~/;9-ٯB5��'i� t|v:I	�����a���b���u�5�My���JϪ���-,��GPƻ����f�=�䅬�t�p_a�5|�-ï��\��:���]a�̷Ԛ_-��
l��˅6S�����z��ΦN�V�|~�[}p6e�-��}���g��[	���"#���=`oC�U����S�z�59\D؟ ���f�< \�z6�KvV�Йm�g!�
%{i�`��&Q��Oi�=3�ֽ��H]K�I��̇���}����h�c��x��`�	ad}^��	i�JiT���×X��a��j���]]hk	�DX�.!���J�*h������a&�=�T�΍ʳ��Y�w��������.�Kf:��z�f�e��ô;�e��e���Nd�N��=�̠Az��-T�S�"Tf<Ӳ�۾ÄoIk=<��{�2j��+^�e�W���:0nhm":ILq�
��v��p�ǽ4|W�
)q�R��[�wM�xv6Y�n�X	�-b�41�U��dۀ>V��/L��hֵ�<T4��R��{�3��s�<HwV�Z�fB�q$���Y�D�+�ǡ�F�*>��Qu��2�c��D����b(�����++����~���!�0M׍]��23�G#�T���s���3�Wu-9[�`;���e�b�"�����ƶ ಩n5��'KN<�
D�x%F 2V���^
��d�4sq�:ֵ�z���w�A6nB����I���{�*^p�N�G=�<֗�B�Tu���%WW��FX�+R�.�!�7\v��Q8)�o�g{������_~W_���fDS(������Փ"9\���9TȨ�jȹr�]S�%Q*�g9\�p*.s�t��
*�'.��TG&\�*��Dr"*�"���QTT\�A+H"��\�UW(�EES"����*#�AE0�
�
��* �rĪ!D(�*T\"�J�\9Ef���"����ADG(����J.ʮTU**)��Ur*���˅�.DUȊ�*�*"���Qt�p�쨸Dr-iU��We��(��Ux�<IAʨ��UW*(�ʂ ��QE�.\��ʢ.�"�p�QE"+�r8P�]�p�(�EW*��ӓ*N��Q�� �b�})�l�fo9�-^Vv��w ][��V�\͙*�
��B O��6 vQ��A"b����>��[�fi�{?�uO�}��I�֓ю�-���@���IrGU�mdv�eM.yª�����c���V�ҵ��y�_ю5S�*ʞ�`l���I��H���w8��HGn?��������Ĵwr K]<<WU��;>_�~��+GkEVzl���/(��=��
��y�A {MB�1?S��7���A�gW��W��[;�ڦ&��Zl�יs۞E/��v��<�+��
�ⷪj���C�N�؍/O��xn����qZ�א�
�\�C�cvl�y�̒ly��B�W���>O}7>q�Z�S�y�v�=:zU�쉢�.���p�3b�UU�UE�k�I��?Uh�C;Sf��~��ӟ�x�OW��(L��i�خ��u=L��Hg��+�P�7������)_�<3�o�Gz�Sq��`߲���	�3�g(�I�����]�f�Lm�2�/6kM���7å�����{+�o����k���y���2Wy��3z51��i�q��:���+j�z����@�}R<6�9�i�x�U�K���<��f�e���Ŗ
�����h�ʗ7eK�SM�"��壯d��\�C��z�ܭ���5������4�t���-��_��ʹ�磣���n���v+fRE� Y4�|�ԅT^��-�ŋSw]q�3�O.뛙���s;���@�h,�o�TjK����h�ޏ��5�_�u���#�3�B��c��Z4���n+�w�;�>����c]5AYf{ݖ��x�W\�U,����)��1l�}H{��(��tE0��uU�1}뇄�1SV�K�&�n����\�ѦG�T���+�q�_�����\m��|{?"��s�7 �u���e��FG���_�H�d�0�x�s����ѿs�S�{��N�Юe�OD�+�ݾ��j�Z�4�7O�_%Ss�z*�Y-3�)�Y�«�h�?;c��TG���~�\xN�Y�哢frs3^⡉g�X�3��GspvTvUH�W�Y�Z>̈چ�7/��qґ�~��Ê��=�9*���6��=j��Ζj=FSgd��r�����9�-�ơwT42Cx:���s�W*=��j��}��S����q�ˑ_<�tE��Cŋ:%x�Ee?S�ӹ �ӽ�{��,���w�y[�>}�P�5w&�ex�M���=�~�2FB�;q���Y�n��BǱa���.�)�J�w��zh���{ 2�T*=\��s�~��8�v���^��G-��u�a{<��-����st��7��m�Ԃ��|�O?G�V��ۣ���+Mn�� �a4�sg���{�����6:Dbwf���������Uks,R5$��NrԨ��N����j����8P�C��
���%��:��FIc�ϲ1?P=7�>��ۀ/,��ɸ�6�>���Ogt�=l��:�d�B���0�6���<�� L%~��T|E���O=�&�k�� ׊�ٕEz�1����5��I�ꢎ��vv3�P�fp�~;+��&ջ��=ޞ~ʲ�i�Z��O�����Žʑ�����E��,_em¼�+����NO�yJ�Í��y��ͬ{�����gk��9^�q7��M�ڑ�O�p�LeFMiy���:^�I���}��)v���b��M�4g��i�2�v�;��_��w��2�N�ٹn��k�aP.�</i-V���	�{�H��������yי�W�����r���oy��X�r�
�Q3�n|3��BǯO��qS3@g�<�nS7�L��ά0�J~���u?W���c�bM���yG/1vTԺ���	@>����M7@U�^.�j5~ڇp����}��Ϯf���HN�mks����o��u��&YO�2�����Q�u-�
�|}써h���>�$?ʅZ�Ç�gR�cu�De��z&�]U����\�J,�f��<=�z,Wƫ�tc��Q��x���^wl8�!+��+�
� �z�jx�ɥM�g��ʝ��G)�\����v�Fޥ x��̙�9E��l_i�ӒUU^�7J�|ݯԿ�����Iex�#�t{)�~���d͝�쩑�ϑ���톞vf�_N��g�g�����=q/��9��Q�~��߷.E|����|���J�b���:�4�䙕��<I���KӰ</b;�����3s�L�^���1ٟQb����~��f�R֭�G��9��ܜ&'�r��χv|%��Ud��e��>�:�r����M�_�����Q����h�
�^Gs蛨���}�z�Miz}W�ᢕ	b�]U>>ݮ��f�?���*�o���23O��I�F��Ux.���d�������f�j�L�z}$iC��[���#t�ߐ�uS�/g�Y~�������}�G�ʯ͑�b��w�X��ǋ��`�Ν�>���>��}�,U�l75� dw�o}�q/�S��Tz���;Lc^W�`C3����d��fN{e
�o�j���k5=�q�^�Lz_��q�����:��݌���ZQ�o�_��߾�ᕓZP���u�1�콦 v��#[���u����	c�a��&���q9�G�)�*�q�+;Zru>�nŷ��<��u������@����L�[X�R��>�Zg6׫R����W�Ct��ܭ�����F�]Y~�K���˝ᣍy�n�K$&V�w����.�v�cH�B�{��wR^�1膴S��s�J��Y�WLa:�dςy�!���~ӑ�w��=x��Li����#n���*wH1���cH�ҧs�5�]뇀�{&X^<�a��x�~?g��9��z�ղ5#����j���z�8)x������ϟ��v]0NQ�&"���ϓ�Іo�EU�ch�~����/�*��+�<�#�����|W���ȫ��[/>�A�P��R.��r[���{�{G^����ҙ����U}Z��lǐS̿t�5�w=��,-���ٿ��9�>��[���P��U��FT�qXG���ς������`z�.<G���s.(c���}ݐ 0�z�N���(R}8bs���WO��@h�p�=P���9�y�ׁUh����[쩕z�ql
�F{2$vO��lD��#q�=��	�};G��Ba��>��W�3�ӑ�V��ݾ]T�O���z�kO����	���t�/�ꚰ�nI�9%Diz}E��x����[����v���׾h�>t&:�|�l�/z��9��y��'az�%�\ׂ�7>�8^�{�G8�U5��N��1���J<ԯ�2�m�K�8d�����G3�LnW���{����h�,��5���NgطJEnB/i󙲯n8�ޓ��Ƿ�V��p)#������^h���U��*WW��b�X���-bQKDL]�ڔF�`鏯o�U�џl��Ύ	UT<���x��V�(���9�:���O����g�.:��ib���ή���B!߾X�X~��6�	W�<69�� dw��;� ��\�cBؚ�}>����k(���T�;N�v^R����i�@�tGSw� b�W���R��Z���9��f3J��Z�<��G��kE��m"E���P���[P�3��o<��Mh~*��	_��{�z��X��YS��=>�s^�내����4���jY�Uhҧ(��������	�ʶ=}^��'˻ul����ʶ�}��W��\�|V��F��n�o��Z�v]``�������Ù��F�������>�=�<wf=2��#������/ţ�~�"]��ֺ啛�"��n�}��՗L��Lab?����O���c��������ᄶ|��p:Z:2R㐟�x�<�G�ລ��e��;�ؗ�y����揠�h�+&[ TZ���6�[���y��{N��#bV:z��O�іtދ��z.��f;ѦG�����H���KA-fDmCW=Ŏ�^������>̀��tS.�n��?��kF%
tg�����S�8FT5=m��v���̂�wZjۻ��;7WCf�'[(��Ǭ>k��bL��2�vof��t�Δ�c3����)jh�rH{��vG�`V�Q�0�U��V�u.�N�q@^�U����ɼZ�Vw{A�}�dp�y~���zni��6vHO�(��Ȁ��Ba�ѭ��N���Q��؄��D?��}Y?`?G��*�޽ ?mԍyT���ŝ�znH�s�u��b}1gj`�[������%a�ba�ڤn��������*ez��TG�7^�Q�Ό�z��u[���,=�G��:�d�b�P�϶��'���=L� �s�.�� )��7<�����3�!���f�kbY�0k�;[Lz��M��>���@��/M�N{,p��o���(��D[�;��U-��vN����7��f�6�~J�~����K��,w���Ы/z��ݷ��o�ك�8����f!̱�(3ћ�cMU�K���j��=��|FG:`�o�nC�����<{>�U�o��c.#+n���s�\w���������ss���(g�5���ߋ����g%�����s�Gi���AWLg�2��c�6:����%N��<h��Ǿ�HNx��k���g�v/Ӽn��EU?C�����r�Y�qR9�R��E!����D0���0�uֻi�(&Ʃ�:�뽚�w[�O�7�"�������`.B	��H��:'�=�rC|0�˭I8��ço�{���p�[@�iG�ܹaBá����]� �܍�Ȉ�y҈�ZS��̒�|�;%&�9�f����պn������~�ϑy�!��~�ѱ�^g�._�D�ز<EߣzT�a�����5ƌo�q��ȉ9��g�ʞD
��)�ɖ�]�ǟ�F{���6���*�O��k�1��DO��8dB�㟄�����"j.�7@U�^.�a��������53����wiZ�����r��|�
a��Z/�W����˦^���>��9FEԷp*._zK���۞�{\�[�Uܳ=g^�/}�v��~��g��[����%ޙ�4gz�Fn3쫸ްU�~�Ǚޫ9����l�j�����㞙�%��E`ۭ�r@���7Ի�lXsN�#r�ӳ�ܥ}�^��&��pir��|ޞ�u]nc�{�'� .�츟R�pt��vhU�qA��m������؝g��G����bb���z�ú���bצ�g�=��q�������d���5{O��a��{���Br��(��*�a�O���kK������:z�z3�3#o޽b�Y��^�>�tY���9�*�T�W�z��vA��f�C�ͯq�/���;�AVw�κ��pc��Ȳ��JE� ��^jQ� �PI��ư>�s:����]{���]J�������yMl.픚�|��7`�D�%;��1�O�h7����kh��w�*^3���xb�sK���]�:_q~TS�aI]s����Y��f�-�.>wu���vY>���:j��z$���!a8X��V�ֶ��&eA�+Vwu�׷Ɯ�8���-S���5� gy�F�۷o�s�����q�����;����<>��^�Ǡg�w�:k��>��5��M��F'�*�{=02"_�x��1=�s�;��߮ �Y�k}���/p�}#�*�ʌ������� c��ζ �Mߑ���h�9��_�
%?H^.�ى�=�`��kƺ�JD��Oz�=���t��L�7�>	�����z����:M=g�j����S�E��0�%=�8l{��Y�ӛ����&����\;�)�%��ց�۪������{�7n+ҝ�9+��_���_�|VԳ���N˦�@Kupԡ��5U�hkҹg3�x�N1�F�T;�s��>���_��z�0��e� 6W�΀}(�,�"f�*�)c�L�IC�^�\}r�l�l���ξ���3�����̌3�p���G½U<s�}C*sޕݽ����4||%쪑�2�V��^9�l�*����x���������e�!s���&Rt�g=E��X�RMZ�IE��'�g0`g����������4E.i���ș�"y�%w_A�DDV��d��E��	:ê)��AŚ松ve�b\d�o�i�P�;+U�N��Op�m>��Vi���0����Hr?zv^�Բ3�V�ï���5
щ�7���͓�>�i���	c�
{���:j�Iv��}f���׷�k|�s@߸ր��#�>���U��� {M��1O�h��ݐ&���5��ނ�5x�#�<�գ��@{����~��g����P�]�TՆ7rHu��"��*v�+�.��W�ZUF�Q�b�_��l�BO���gG��P�}%��D��Y�.�4�\I<>_�KWu��:bke3:�����>��~�<m��G��v���?He��к#��9�ٸ�S����}p�lq�����~��V���o�}���ƿU��#��d��bT/wf�{���Lz/�.9'<v�v��y^���l֛�\���`R�d	{o�baH0��'���ʎK�be~�)y꼿��k�]�6@���/�k�j״���z#\������qXf���9��(g�;^�Uc=^~��N��{��hn�tz�*d1��+�w�;�G�5,�Y���û��
϶e�����NF�_��\o<u��;�QW�w�
ʫ}0��.��:6ǔԎQ�cvmZ�a"7�f�O/�-��QP]��ZU@-³�<��Ir<q_B�%��+����ay9Ծ6�ݪ���,��ؽ��A�gQM�al�Ŧb����Ӽ��<�'��dk2�],���Ç�����".��
FЦ˼�b��yw�Q�fZ�q��Y&��d�K��-��`K�q3�U`���-a��C%%���1�M]rI�fuAA�bP�ЭZ���+��֓�DP/��>(�[�����V� V7n�$��[-n[2Ioz� �]�r�c@q�9J��F�j*�D(�3�U��惦��c��ӟ+��억���g��X�%Ө��C�sp�%Dʉ<'I��7x��j>O�6��(ĭ��u$�.�:9�*���Ա�� ��t�[��	�(�b�z��x��ѹ��᱾᏷��rnЮcc[G󖁱��K����P�̅�ǩ�"s�@$����+ë�\+�,@	o�˚�~$�̢�$�{d�����e9D�!�ՒB�;��˸��F[��)lZ6��FAǨw{���^}��$W��[2����7�4�[g!�z� ��D<�F���u��V��B��|�Ke]VOM�����U����m`��<�D���r�'�0w!b���k\��e�|�wS�g�g#��E{�hV���Ǫ����\��I۠�p�ĜvuamݍZ���/�nt�4��z��#�N�v�ŗػW�weZw�f�4�3�K6`(���=t#�_���7�ҏ�^��ko����^�c)h#:�]��4X9�帤"�s00ˊiO����Ϗ�_l��`�����X���Sl��ъ�q��m�!�8��f
������4oH��aHe����K�����n�E�0455[�>���b�I�4kn��tc��;�Z�S�dz�����=�)F7%����{X��	��eqm\�=�|F-��
��ʺ���Sk>���c�c�-��e-ǲ�5�����έ�ې�;�Ռ�]�|���[X�H���a;z6��mWr�{"�sqfr�����=�N�W�������Kt�fQ����[5����~�J��c_EL���.��݀��Fj�:���uJ��Vw�I
�v��Z�×|�T�|=�k
j�p.��7)�w�ڜ3)�M����;��%M��=䉂N�S1sc�`��N"l�ښ�n!/J#�q��	g���c��)��빚A�{�H1�A�sm����v� ��}�e�IhQ.���ݳ�ٲ5��f=���&*u��V6c9E�{!�9W��m�r�d[ �g�#��rQ4��@�������u�-!EK<-[V]�΢�ჶ����T�j��^p=u��:]ߍ�d�Ij���������r[&lI�S���#��` �t��Q�x���Oa74PJ	V�N1�/el�(���WV�I[��ݧx� fՒn\�R1��ŕ�6⒮�x�:i�S�M�%�����%��ĂO��~�r|�Qs�s�r��������QDQr#�"

dQp��Q�eUgB�.ʂ#$���HG"9�r�Q&U��U.Q!dʢ��(��.TDDt�vQ����.E]�t8\"�YӲ+����r�PTU�Q
�E@U\��G"*)���(��QD��E�N�ȮW"�L��(�\�$"�dUs�AQ´hE�X�;"�".TQWU�R®W.�U\�Dd���%vP\�((�"&Q2dQUW$�r�i	TG+��"�U3��8Dr����\�*��.h�Q"�UvAQ@\���Ӈ&QWHr�(��.N���~�����}�w��.���&Yt{\#�oEk�9��j�^���϶u�O[ŏ�}X���9��C�|����W���*�b}
8��Ι�1q�>Ns�2U�����u�Q����j�=��H��7
zT�V�[���j�>��H	��"�Z,\d�g���C���>|=K�?O��~��L���[U"f�ʶ��/|9zl���� �@>ʩS-�*"ԯ[,%=|<1�����~��qu!�+�7<Is
����ދ��#�[���9=���b�W�a��ɇ�.���q;gM���5תG��noux��#�{-�����=y�;$'� ��}�|KGv�i�R�zr��]�����M�sڇq���~7<
�����r|�Q�v<X�0{Ǯ����r:j�)j�K��&��Oi��'���^�&=I��8�s��s�{@+��\��ؕ@4x�����q��l�8]<��|ؾ��w�=�C��zdTo��;>��B��MLZ~��>�N@�D2�bD=����:����I&��]N��7Q�ͬ茟�_k�j6��)�X]'��������)��Q�^�����ձ���FT+O����u�V�q�^�qޞki�%+��n{=�����"oGu#0��0���F��@c���V��Ϋâ���\ֆj3y#���N�R����{g�S2T]������ֲF���#|�wRć%�zx����S�ս�[{Ɂ�OW\j�a7 ���k5W%)XX����o�,�x��d��T6O��X.#�x�J,�)~�^?'���c߄�~�N�?eT�i�e�-�� {�W���#�}^��9g��5�~Y�9�tZ`1�/���%ÇVצ��=��/S�>T���t�-:��~��m{U�ﲧ�'�<xg��kq��^�H�0R��]SI"}��5��3���B���#�a�d��I���8�C�+����}0Scx���%w�:9�|}����U`L\���:��ϑy�!�^����:�=^�q��0;��W�������n:�QF;�kL���s�U`Q�@ȿJf�&X^Χ���<����������v:�krG���>�:�U!�p��X�G�7��܁֥x�ȍ�h��>]^����fj�3/a��ۊ�s����}�4?W��,�e8�!���`{�>�"�[��L��\�7�%n�o;M�36r���|?S\j=oԑ�����?D�e��g�\�` 4{�[=+:|��=�I
��G�I��7�x=9�����w��㞙�%~���n�;�t@�z��@-Q��������凛��1N����� rP��oZQ��g�_<]c�Q�\��|<_��������-���6stw�ǁ�kP�7�RdO(��r�V��wb\��t�%��xoP���%	���0J6�<(Z�Y�#y2���7�������FLy��g�XL�9�tdJӹ�/oz��:�u1mO�3s�V����"C�yYf���1Y�}�_�߫.<�kI�������fm�o�'��~s�7�m�a�z`}��{��9O������z�5bUyɺ����a�g���z}]��u5�����p�%���U,���P\:��m�����eJ5��fǴ�n�;����A�#�����F����71h��wH\j�,�s�t�?Uh�3�6o�Q��QM���� ���G�_y5��q���G:�7���f��	�~��D75� gR�#���q>Rl�~�'��N���n����n��w�/�O��_�5��2P�7�F�n8�6������`t?V��뉎~Q�,h���Y�19��zi�,�8�����kK3�:��̏b��`	��W�n��q�C�osɅ�Ӟ�c��L�F���>����*��k��L�8O�k�C�T.��˰����_�|�ך>����߫�\D��4g��i��ӛ�s��ɨ�&+�p��NLo�'$�
����?h.V����C:"�{o3{����J�Mj��t���p��|G�}#���.��ׅ�y�(�s|w0q"nF�5���Lث�x��YȧB9B���5�+G\8<�ı����F�{�����Z�w�f�w&(v�#�Z��T͕z�� MrC�O�O*=h�~��x�ϯ�ǁv���TY�~W"�A�鸣�b��I����ݡ����>�w9��O�_���I����=����>�_��,��L��T�k&ĳ9��~��b��	�m�>�_����a_N�ߩ#~a�����k�e��2�/d���1����>KuG�1>f�:%vET�����r�s#g�T_Wr�P��\����ۆ�䛛���O�ؤ�!��;2$vJ���x���ىA�͓����s�c��W��)o+}-P�j�f�l�0Z~��U�+�p.U�ā�;�>���_�s��[]8�6��D��f&����\Ϣt�/�)�t�6���>*� ���^z��C�nTՆ7#v�t�V��E��}��!��G�d�G�G�H1��z���~�<�:���2@ߗ��Nk"�z�{[w�S�Z�bԡB���87�;�5>�d�ic֮��US��D�6�U��d��|�_�z�;ڥ/��I�I�w�OSq����N��z��3[L	����=t;?H�Y��/�rI�r��Ӎ���Da�x�d/�k���f�u:�ֶZ(��Z�) Z�$�R���@dH�41�ۭ_N�/(�D���h��_=ʵ���T�ʳ�ku�H�PA�s����r�ٯl���V��̇��죯r�YS� ��]:ߝ��.F|b�j���T�v���yq��,\f�i�@���� ����+�j��(v5%7xkJd��=�^�y���i�����O�a�3��V�;��u��r���^JK�j��_���3o��������N�ǫ}���������H\cږ{=U�J�f�+�tú+�z�{���nz�b{����
��%�ֽ~ӛާ����*=�wᜤ���]V
ج���y��HZ�Ĭ9۽q�3�Lar�tѝ>������x�����s�唻�'�X�՗;�Ԍ�����]�V�O2,�X�[>�$�E\�4tc�J�o�M7���3�w�3P�r��
}^�ۻ�P\���@72Ed�dEx��c�_�G����l	��|�\����\z��<2�I�;�G�A[�yd77��PeT�+԰���l�X�}��7u���L�y�}kw�NG��k�cӴ�~�<;���X�K5�2<�����������mUӃ�?`Y/צ�klUSy����	���Tz����=9\
�z� �ۗ"��S�<�x��x���*~�H�PK�͹���̤�ݙL��TtB�_�@���:Q㤚M�
&�.��oP��c.����es�w�G][��C��Z�eJt�`\�5v�<�Q�+�����1�A�׫"�U�����6+���Ǚ���N�+�"jv�RZjn�������U#�����wH����O��Ϝ�o�����yP��sDy�S&|�kֲ���p|����/CܒE��"�};���/B�0��U鹋O�<�N��[�����h���<Q��>�JOaȺ��d�Cܝ��'ä�k�vX���X��}q5�F�#u���"����o��/���N���VM�ЭlW�'��5S�K���g#�;%�Dʋ��)uא����/]2zߪ�ɵ�5���'�_ު(�هgc=��6�Lϑ~kTt{O�
�/7�M>�e�>��w,!9�{�@�o�nE����'�G�Ό�N���������g�:��9�}�*��O��7}s�I���7�F�^�q7�۞7	�H�<��9���+�t��r����}T�VMiw3�b�\����>;p׮_;,���;Ɵ���k�3�7�x��O�]�G���/�"^ւ�������b�ɝf�&|�Ι������y�J*}1���G�{��I���[8���K>��q�ˮ|af�U3q.q�9V�<��L�d��7�zѩ�5o�݄Z��6�d��q����S1^��}�����̘}�2�w�����4<�����r�+F�Nx������eH�a��'S���Ts��a���X$��5F̄wi̝/jl8�v�v����CҀ������5N@�))��-�ɋq�k739q�y���#ؽ����A�x:��~����`>Ϧ��SrE�^.�s�'�C�ڼ~6w5����Gќ�ǳ��#=�ݐ���_{��𲤲�i�����=ӟQ�~�@�T��.���_�\��q�j<�_uC��z�9���S9����e���3�-Di�5zA+��*����{�*=�nI�\�d��}��k�\2�zO��x��:]Ƿ.A��n�pY�u�YQK�yҍ^� {��f�bP}��DӞ�џJӹ�,ew���W[�Ϝ�{�=�m��Z}78�g��ˏ�n�'ݓ^�P|��z��ݑ����5[F�\��`,eF*�X�W}���Uq����Dϯ��T'f�� ��� �����u�{&��en�w������Lm��c�nU�FJ�Z�C΄��L�v!{��9���h	����7~��]�l{M��C���C�;�����]�پ��g�q���ڄʪ�Ԯ呟r�G!���5&��މ(�����0u�ݾ�u9��޾P��c=��;�������7Łj�q���G�V�v�m�ntwպ-�����W��We°� �&�A�x�eMj��������ex�i)gX���س<�]B��/�H4�%��2��{)W�7%��X��z���dHI���7{՚p�ɜ^GBGK;��{��w�x�h۸�ƫ"T�28�Ѥz4\��=ҎeY�_#�F���N%ػxm2
e�_N�k����	���^MixX�;��鸞��jy����`/:|n.�y3�]z�ay{�~���}���o��)g�Lf���L�ƹ]�T�m�[ _?N��@z��NۉvOox�׵����������b���}���T{}��'<w괿�q:�����r]��j���������zy��;�c��f!���_�����I����p]뇒=�錁ڧc��r���Z���d�L����s�i�t���~_��[VԳ��D������b�6=��/,�s/T= {_\+ޞ�!q����:H����.;��%�|:&V\��uО��bnw/1�� |���T��O��W�)�3Y�¾��RF=��T�ȏt��A����3���^x�ulf��'��#�l,��h[���	TT�8��gB*u�4������{�{���?H�*��,�+�LW�����W���	h���	cǩ�9��S+��^��Eʚ����0VD{��;�ndHy>���*�Sq�=��1�O�h�L/�*��N�\:3�s.�ʟsщ.�t��/3���le�)
��bQѵ:�չ�z�LX'.��:#�)��D<;}�D���\W����[��9�>R(�A�g��;�B�{G����0Z��v���9�����c�z2��Ƚ�[
�_�paY�F���,�P�Au�o�`S��ԏ�f��W�J��3^�gv�*s���^�U)5izU���޹�q	���9��y���}ES^ޑ�Zbs��������r����Fj6X�3Q_���y���c�N�����K|�y����{��io��zG��}�'���;��pNg�2�i�?%~���9�R�͂��PBHȞS����sEϱM�u(��z��I(���C���.3f�޹}u0/*���Y�c/�=�������`{���#�X$Tg������O�aՑUFV�;�=]e���+*=+�ǧ�Ε��ܰ�:�1�ՁQi�x�l{��\/m��>�q�/�ǵ,�G��iS�X��w3t[�����$��7�}}x�,f�ׯ�r7��_m��x�����Ef�"���?%��g�{�kRޚ�`�W��	��xJs�>^��JhM}���9���|r�?�9ˍ7?
w]�V�6��Q�˺�zl���^7� �>��&*yW>E�ɖϳ�`qţ��|=K�U�C��v�ig��.<ĭ���\�K�F��]Hx,kl��:�A��2h�=Z���gY�ShM�H%iP�t{+D6�*�4��.�u�4�|�"�B�	\��w�rVS���vU��c���]��O�W�t]H��^�Hj��@�p;���FT��r�G��w�Գ��;7΀}�U"�l��Z��5�,-�W��"���ǰ����c"w�<w)�� d�_�����������PdUH�R�K��*`�C~:g�o�wvWw�=~���b�N�9�H��#�G����5F�s{2>������gd�@j6���g]n=Ο^�����B�w��I���@�	�Ｈ���uN����x����|���o2z_�����rG��+N���9�/w�ǩ>�g>s9��9/ho�`/H�ǀ2��O�7�O�7*9y�dGzn��n����EF���X��b�ڟm�ZO�%I��^����ym��iW>d��~���?�ڍ{O](��-�O�~��=:��d�;]�K���.�ol��ڣ�/T�����gn ���%i�T�=1����0�#6�����Ϳo���Q7����oh�f=��=����gz�Y��.�~�74*�7�?~���^��k�_�מ,���/D1�S�I�l��p&v}L1j݁%����`�q�ݹ�g���A~��Ϫ�S+~��x�"��g?�w�zY_v��F�C�����Z�L�� ƪ*�Yo��)2���V�n���9�"dP�鎰n;��
�V������T�1P��K����A@�n���i�Ry����E"�����S��f�m ޙ$\ƻ�3.���1Uo�-�)�o���XA��{�/�;��bdqY`؇n_<(��|"ו�H]���OrC|V�m7�����^!���<�l�r���<�rr���ZP�+���'�H��76�1BTpV:n��U@��}�#";��K�!{P��-��e��;Oh�H���q]Yǩ�q*3}3�Mӹ�KǸ�2gê�;ݽ�-��n�zUbyS_M��6$��;�`�0�
�8�ht�ȸ����[�o���m��~9��M�g��۸�
`7t��2:��Hrnm�/���������_�fj��ҾBں>׻��k�P]h9]�VMbIP_mt���b�At5/��T�o��0tN���]`u�*�;�S]>7��*��V������ݝ��>;�c6bo@E}��h.X���"��4U�28*�4�X��=[N��\�k-��h
��w�rOfy��/e�����Yʊ�j]����,=����\����;vt�s)�Wb	$w�EC�p��
�bخ� �I��W��\� �A#49}(B����Q�ly��{د��Ⲇ�o��k8��'vQ�l�'�R�Q�)&g��D���J7v��T��&V����f�TΕg�e�7�H蠵��ڙ���u-軉�Sא���y8�iq���k0������ƾ0�9\J�l[o$��;{���t�C��;/�Z�����:A�`�1
D�=�.G��su�O�C ���x��yཀ&�p�6D�����5+��P7v�K=�І�|]�����;>m��Ɋ\��v:�����j�Y��4+V�=�@F��Q��Y3�{ԊM��Wg~V�c�S���:%�tQ��ĺ򻯼���\��!+^I�}���U��Oy���А)�Ǎ�v�wD����5g;z�9�gp&Z+�o�R�[�]�`Z�z�+A�ͲY��ǎgb�#�S��cr"�}��rٙ�����u��^D^��ӷR�]B��2����%W3ά�p4������mYo��K]hA�8���u}��P���Qg^omE�iKU��ط
)��ur�&ZWO��55YV%�nerU�ֻ�Kk��f�f��x�a4(�?��Lg$i	�Â�C��Fԣb�A�g�h*ֳ�$0�`�e�+e�r��۔�[�cN�;�fM�%*#r�ؼ�w��Ewl�qs�6�|�c8#<��Va4fq������%��f$U��� > ���k(��Eːr*((9kNBdQATUÕ��\�r���*
(��J�����Ur��W*��8UDUPUZ��쪪(.\���(��J(�TEL��HUAW�����r"��E\�����M�yN¢�.A\��(9QEUS**�"�]ȑܥx�DZEÑ�U�$�dW+�q�j��y�se��E\�B�
"�.8�s�H��d�Atɇ�<Hp�Q�,J����$RM�X\T9Y�;M8�:p��,�j�P^D/x�)0��F��������Gr�,��A�����)!���L�R`R�uÙx���8T��*�O9pA�4U�'�(9��q�$�e���~W�a5Z̦����;=H)�� �o�m��������{\ꥑ���)}�X��oGH����,E���x����^+�Y��n˨�%����o�@��@/�S��U���2����>�G=���!�#�5q2�����gҕh>ʦ2�kK�ɝ��ƹ	����*-�g�v�;�dEEuG�8�/��WU<ׇ��7Գ���l佭eU�?\���:��L��2��W�pz�Wz�xN~V��c;�Y�n=�w��G�:��n�Ϥ�.n���ȁ�E�S7�,/F���#ݓݙ>��c�U�V�{��{��K�A�p:�p�G�!���&��LSt]%^����Mx�^t�I`����g�mEr����|d{������+n�znj��L�f�(s�9��.��x(�
�K�g�O&�P�z�8�%ϸ�t.��E���/�S�������g�D�=�22��^G 0���ﺡ�GSY��o�F��������rTe�V���n�y����� z%(�3���W?S��ѐ}+N��Tw���W[��@�uFy��}u��v�.�^}3蝝ߞdK�>�ʉh�z��ݑ����5[GY�݂��1S�tF;���)��l��u��sʮ����[:�ޭ�;nT��/�:zC��h��`<�+��ĭ�Vu�C�em�����N�ppX�m���N��o��.P鮸p�x�����p|c���y!fo=�PIDJ�4� Ξ�m�iQ2j2���2e�+��|�#:�Wx�ݤ��=�9w�'��_�uzǔ��� ������U�{&���[��z�NE/@>{�LS��E�W�(9�Օ^�ᢡP�+UQe?H�j��㝠){J5q��fǴ�lk�5Zb̿la���;��/Gz�ǂ�g���һ��UQd^��<m���{b�ٸ�D�su�s]3�5��_�,}��O��>�},e�*а�����̐�V�����/}�<n7۷��X��yb|�k/��^�}��7�����^MiW��Zn5��On'�-O��:�����_�fK��M�ؽ��l�b>�o�&�V��OMw�,�滛�3��'<z5��G�2�)�W�L��JQG6���X1�|k�:?e�y��a�	l��ӺJȪ�a�WL^L� �Z��0G3�y�{�+�����$!��'~ӟo�y���x+�yhm���(-re�}.p'9��X9�D��ϋ��q�^�Գ��?Ќ�7�?�g9�C�<���"<�_��a����ʖV?Q��BټRN�׹��ƪ��dȠ=�5p,���!q�za��#����>�������Q���̿vK5s�����a~��@U]��ԝf���u� ��.���>?DO��_L��5V�:��i݇DK��O����R�ܤ�fԴ�¸��9�m�����8Lե�<�����[}���[Z�7�L�<�}˃��3t��8��湽M�/�m�ׯ�����f9��M��C��	��� �*�]D�`YL����8������l��zx��7������Tu�f�|�x#�v�:8�>`�#Al��ex�9\�϶|}}\�s�HE���Q�mIW�>�83rQS�����Ȑ�\�/>E��(>ʬ&&�W��ĴwEC%�&o���\l�k}�����/��^�d�W&��*�����/������� {���1��uK���>������K�>���=�a��LO�'�l��}@{�����)�z��T<WU5%5��g�����m��7	`�o��
�Vɯ��>�q��R<���8��	F���~��,���H����tؓ�|Z��'+֝��o��^<�Z��?�xaI�������2}1��'L�v���1 �>զ��k�9��0��jl��!��?T�����:���>âp�k���F�a+�G�૕��T�R�{�Ehͺ�/9���m;�S���5���1_w�w�N3�f�e{��p�F�}�!n�{g&,�ov�T�ŏ����~ {�S}ާ�g��.#}��/a���>��VET<9;0�ͮ��Q�H(������)Q���M:�
`$���~�e������I��X��lH�X�f�h����}S�ϻs-�Ŷ��h����Z���7rcۤ�IH�]L���Đ{ف\���72D���ݝ�ʵ��j��h��l�C=΀���<}[�_q+ۈp���lgۢXۏU!�N<n*L:�Jkf�*���i>�~���;	�6e�L��ׯ�w���w��玴w��EO>Q���Uϯ�{�{�e�����#�b���2e9�'�Ҿ�!W�y_�|�i����(�^+��.k�_�oѮϊ�j�[9*@}3�eO"*�ȱq�-�s�@�h����vh��������<;͟s�q�����,�f5�E��dUH���l�QjW���i��"n�w�ؒAz�>�ǳ|������{���ǆA[�y��͝��UH�R�K
W@Jlu���{i�L��z����P�}u�|-ש"���~�#G��[��^���dy��l�	�����7���j>mzǎ:zp�Gw"ǼjuC�}~��NW����ۭ*�b5��v-�z<:z�3;�ܣg�s��Ee?E9�;���t�/gxTz��S7g<}'%m ���"��9~�<h;�sS���^iN����<��z��;#v��}r�ȯ�\�g���D�ϹW��9=�O��4�xM��,j�hIܻj*�j������ޫ.�-�y�w����qf;o�`�ݽ�6��}�t����L�Z��--p����Gչl�k����Py��6�뺓}P��QN������{��j]z�awː�6<����ṷE�?I�]�y��琝�ԦH�0qaޢ5�ڤ9�c�5b/��:���ڿ���b�^��G.���}7P��K���Q�t����������{���1��|�'G�Q�����6�5��d���?�?p�&��ikb�~OA�Ĉ*_�S5��yb3���}��zPϵUE���O[�P�6���_z$�ˏUv�'j򷦽���/��[<��F{UV��=��q����ǀd�Vx�z|'JՕ���{Mh�����t����w^mn����?g얍-f��������������<z��9��W��MT�S8�a��v)��W��Tb>��{R�����c*2kK�w��Bs��f�^�z�2�d���ׄ�1�4Y�����}��{#�jܹ-��p�V����:���>E�!���32=r���6����P53��xz5:�=���7/���\��Ϸ©��8˜��&����)�o�/]���o�f�����<��(~��>Gm����>�bh�/_�}���.P��Qp5g,�vh�/1W�=�f��Vw��mG�����8NR*	�=�0tC���2
ږ^F����F3^*3vO>�])����Vl��F�^�U��>�wX�޵�F�w+�,�?(���epJ����kk��z� C@�-��q@Q6�j�Y!�2�;�E���F��by��������:�p���>��¬Y0�s��jN}����O�s�2.���T\����ݘn�cgO�QL�����ve�4z����]	ԛ�RBG��zI�K�#��,-9���k��w���x�ޙ�%]O�@K����q{�Ǎ{=�"�*�/�8�3q��슬&~�=��i�_zt{���G��Pn�|�y���_��ϧ�wW�&���(-���G�NMVѽs��D+���yU:�v=����/)�xTF�U��9�t�pxU@�����^E���8��ue�Y�X�QK�/a����i�.��
��Z����~�<��P����k*Q��Ux.�%9�J�2��N{��(������g�z8���ڇ�J�/�UE��|����G������6�6�`���_���8[�!a�D졗�C����{fx0_/l{Y����*,�HN�N��{�5������Kȣ�z��qxL�OO�~�!����1�}���˝
�ܗ���ş��Y;�J`z9��[��eO��5�O���[�����ZY��� 3ߨ�4��r{A���n;��M)��Mi̓�<T>�K
sa�����:�q��n��3[�����WFU�BԵy2�%��vvns��C\.z��p�c5L{:%c��2:Y�j�s�b>�h�f���qugr�ݻ�ڀaurt�N�)qW�� 4�u���V|������׽::�����F��ȉ��=��]1��J����Y~����Gz�����L��t��z��#|���߫�\��4g��i��S7�����河Ѣ��{��@�]����g��d��>�yP�s�i�t��{$!<T�]2��`#{ԣ۰._S��rR3�V�:l���1^����'7�B�u�����#od��}>�V:��)�]�����tr�X�D�U�#�@{�ET���L)�3XX�ա�7�l�"Q>�n�3�Y]�[�<3��I��C���3f%�ptJ��F�U���x�Fς����`����a�^z0�F�6��ǼQs~#,����NnG�O���P}�Ua14����:�?
���4+s�.������yOqb�u[8�k��z����"��znʊhߦ@���������ߧˢ�CP��gh�4�{�Ǭ���U��}@Nڤ U���C����VF�ؙ���c���������{詫7#v��['G���DqzT�"z��~�=�C��^ߑ����l��i.@��ͣeV�f��*�C+KGA>�ơ���)<sM)7�w�������;��E�[�֎@��^�Q'k݋�����WWB��w�e�*<�WEws��統��F�iwE	�⸮w$f��;��wT�թ�>�t��Q�����ی�����cʍ,z�]�;�J�}1���wAvG�ny���Ѯ��[Tl���zs��?�{'�����>âp�k���}���;����m�8�~<Oo�Q�^�3���:eN��/�S�Gz��I(�ɇ}^��i�9�1{���X���$��w[�׀�4��W���;��ؕ׃F{�����7�8R��d�mx�\�Z��l������}����} k���y���N��5��Wk�hp��B�ǵ,���]��U�����};~�eO����T=���7��72ư�^¾�K��T�����y�tb�����X��{<�h�G>��lx�U�L_z���2���L�zs��CU{��/�q]��y4��>EnJ�sw�S��C=(�}�����>+#}DS7-��h	<�苟"���g�ΰ3Og��n/;|&�N�܏z�C���[G��K��XU�L����:9�+"e�E�^.�|DW������3�/ܩ.=�;c��T{������G��D��������$Pߢ0���H�6k��W�Ε�����Y���$�Q�T���8��e�v���0�bw=�b�p�ҵ�B�M�����Vh�׊�6�7v'�d�����'Z�W�tƖv�Q��K����.�GN�oʆ�q�����߲�x$}n����#(�ux����\���� �y/�Ǖ]w�R)����a_��|3����;˚R�և�:�C7#�rz{sq%��dI{I�|3,L?��T;�__�sӕ���=���n\�+�7�5�/o��E�w^�#Е|.6bS=��E3�s`�r	xk{£���n^>�������r�V���=ۚ"�RG�՗�7h�U��"�\�d�T*�'���mw�ťGF,5�N�&r��9��v���+��QTs��=�D�C���/�I�p�����fЪ���+��'���}s����������ށ+MǪ|6�T{�w8�4����^��+ں+z;c}��ϻ��f�i�&:�xj�,��^'���ɿ�����I㞙(������Knj���U��>����U������`T��9��^�
9��*E|��hD{7ӂك��j��鳯阼59<,��f{�(k�.V�k�c2��iph����ہW���}�{s��#���kAS,^�Miw�L�/\���k�B׏����|��Ƶ�*��-����(Y�O�V��A���N���A�Y��K�[���|`#�g�z�o%���ڰ
���~����R�1"����sس��A��	tC�q���G�Em��`W7{���p�����D�f<һ��ю���:���d! �pm^q{ȯץ��jw��z�;c�\��9�-���������&�X�ɝf�&|�����i��+Փ�}��ɾC}ë�v�GF}�>gs��{�ĬW��uό-�eK�e���	��ק��ryin~�����n�F̠���,(<�z3�'��?W�\K�A�S��s�Q����{s���_a�P�]�T=��-O�]f�4ks�p�r�q���ݿC�0O����d�>ި�tSs�;���f�w���|\�NQ�u�\
�|}��j5��T7>����(�s�'E�AV�J���K`T�s��^�/���Di�7D�=�T�ʗ^G 0��l���w-�����K�\˚���^��k{�?.&Ͼ�ҿT���]�q>���6OE9�}+N�b�mNϲ?ŜN�+���*�cޝ���};?]D�3� )Q-��G�������h�S܉���P���/3���_����P؄�n}Bv{�9�=q�w S��\��麇�&����V���.g��a�9ӓZ}���xh�BX�UG����C���8�h
��(���c��.��鑑�3zXf������,|�WS�Ü�#.�1wl�10Sd�㥾�b�턳V,�W�!�'D�f�d��N�m�U�)��z���m�Yj�U�����o7\L�]�8ǖ4��a]�X��%�&v9��Y��8�]/"ĄM�2���M[�c!�O�3��f��K��[W�X����(��WC�e[ü�c�<�%
�2K5.�d�����״5K[���05���h����a��O����[�`.9.�{
V��#���^Gq���9��+���2�t�+��g7ƕ���+QűK���H<y��d�$lC.ؚ1���}Ɖ�.vL?Y|[���D�ydыDuv�c��T�Žwm�wxە�ѯa�*7 ��_Wduȸ�4qo���QEs!��ǣ*�󾾒��Ӎ^M�Ty��qEbVB-S)��v'7oPˍ!Ҹ��ܫv�ۨ�(ѣ��}�3��;L��ti��S	��\+��"�0nձ`��;0L��$ۘ��G.�[�|�[i$L[����3a����-7����G}��N�ư�&-�մя�yس}�9���/����C�x �G(Ȱ��_`�&�rL6ZG.�����
�j�#�=��od�m��!<; ��]mf��t٭�/��m���#���V�CZ�b�	��}��J�1���Y�j��_;Y�F{�/���2܇�^����h���]����D �����4�a\�.�xX}��m�]/+D\x�YJjƱ$	�Fq����<����V�*��]K:��pU�C���D�c%
t�wr����m�tq1�p2�3qrp@m�w:Qv����;^u泻ė0 7�P˻ԣ��&��ճ,�*f��*�Ӥ�7`���[�$��K�eX�q#�ϗ>�[���z��@�:2������0:�흷��juuwGvU�z�W0)��x6��]0+�ݾ����� T���;(V
Gs-�t�E�r���M�����c��hY�[��,�ёܚc%w_aw7������A15�������M�n�>Bu��=���=� �6)���>L�NY������$s���"���+nt���]3����"
ձ�6�^�}xji���TB����\��PM�M *�1�d�"С��-pS�(�xz�^�'�ݸ�&��G��=���^/�b*;�v���ܰfR����7�M�|�ny��m���/
	Ⱦ^k�'�um{{:-�	sy�-�ˣ�Շ��WtZ*��9W���c9T��䡝;K{��y�����ZD%�x5�;��@nH{��x�T}��a�1�t�ya�ӕ��-t=]�����r'�ӈX¬�b�c/|��-��ɘ(¢��eyL�-��k��ݶ>��N�+Lȃr矖zl\}�,ɛ{J4M�zl"���;7>��d�CR篳2�4��C(�n�I�ʇe�I��S|FE)庫��sNG��l�S}��&D7�|�9aY-a�h�y�}��Qt�:Nhl�oh-6(�EG���
�VË؎��u����
���Dp*�:fQ�5ǎR��䨢W(&W���WiP����sH�,,�Q]�]�V�A�6��UY$��2�%��Ǯ�͚ʻ�W�xND��9��(�2"��r�x�u���JQM-D�!
և"ux"KJq�8�P**��VU"�9sp��q�Ҋ�(	*L�*�s�jˡ��r�j'4O.nr9��䭔Q��qW't$��D�H���9l�p�	"I"E���d�%s%���\U!8�g#2*�"���$�e*��\N4��<�x����¢AI���%9�TU�I'1l��Rr���Wq�Y]Rr:I�i'fIʳ��J��͸�N ����RBe帜U�ӗ�)4��&�����I� ���=�|Q�{&�	@�Ǜ��e�N�!�]���t���Ŵ�wlp�/!餆;F�9h��!E�t�%vc�=�I�����7����ނ�����ڇ�V�/���E����|߮�W��㽰��F��3Z��{���-9iX�T�~���ީ����4��#͙�&�����c��U�L�$�u�[�ϣ=�q7[s��zA��~�(m��q�ZU���Zn#\���q`lx�9�$Ե3����gk�=�o}06>~�F�z�w�ۤaC�=���HESQ�ZX��g|sհ��&'9�]������=�!�� ��{�(�V���;;�r�[����*��o���>ꧦ�a�z�ϊ6}��t�f�g�>��k��;�>G\C�\��e1��_c�S5��	BK��˿j{�N�l�蚄yT;2�e���*�u�>�W8���!q/�0�g#"�.��J&����y��/D'DW����6�M�
��'7�B�q��\U�Β7�O�㷡^����o�ݾK�<}��ה3�[V�ߠ#�@O��]K��ϙ���
��C�F�ER wd���ͿTҹY9O�ǵRg=�tײ����Qc"6b[#AA�ET���^+|\�C�<z��$��;:Dnis�Cɡ1Ɯ���,��;8C %HD�p��O�U5*{��ڹ*�����b�n����Jƣ�����z�����)��hs�Nh{r�	��3�*+;�A[w��N���y92��"�Μ�5�MJ���\��|�h�KŏY�������D�x�����y�0x=��&�r��-����۴�:}�}�;��	a��|9�U��v�
����w�ȑO+�p.%Pjw���=Qu<E�����6Ͼ��N������0��	�[8�`yi� *~V���
��k��]}�T���裡q}&hxf�����l��/O���^��Ba�.�͛O��}��^�pz�w��k+_!���� �Ϩ���\s���ͭ6|'�e�35�ic��OX\zmFOL�v���)�Y��t�|��{~;f�~����O�Q=_�\d�a�8w\�pr���G��]{-�K1N�@��q�ޜw����{�k�˔c� ��=RQ۝�yy^��C�N�';*�ϰ�zY��@�_S~�V�	{+�o�i���	�i��k�� !v��-���8�evqs��Q��~�u��5H뎩p3��p��x�o����_;�e�����\V�*D�k���NS80��6�]øɝ��@L�,f�^�i��K�}�~��'j�7eRuTs��z�Pݸd5cp�sq{'�[��g�$әH'����dE��gB	�3��Щ{E�*������s �;1��Ƀ۪�,��L7��g�P,���\p-���4Ҷ��Q�ѹ��
�bg�>��,�u�:�.��X�r�V�R���sŇHᬾ�8�v��xOծ��e�
Ȫ�&���&S������!Fb�x�.���<[w�9�W$K�y��3ᅣ��ѿ�*����嗾�%�-���b��|��-�򃃯�z��e(ՙ�X�|:}�F}����*^z�вe���\S�p|��U"�l��{���I��M�8����=���\=[��xg�鋏O�=�H��~�c3Q�1-;.�+�%��o�n�\�oFL׻�G�P+g�� ���چ������ԑϡ����u�£�n�[�zn�{�塞sf���圐��w,�l�"�������ǒU}-_���?���*���r-�K���o�B�՝j����Td��ϫ(�g���T��w�Ǫ�o��\����rLQ��X�/�J�g��wh_�y`T<��q*�h�}�����v��E��"�^ׇ`,f{;�N�{"���Q���#����Փ��J�?��ITjK�ޛ�{}�z�O�Ix*���!G�0��w��g�+�[�穒�B�.�?H;=����c;pzXv=S�VM��K�=/��yT�7�<���EK���ew�u��we�D�u̖;��x_ ��+�Ε�FotrDA�j 6lӇ"X���Ц���*m��_x�\�Î�gլ[7��g��x̮��&:�iލz�S���2�`�NO�ŭ��*�L���Y�+��������3����x_ڪ�#y׉��U��46;�<vq��G���5���;�=�s�ꇆ�T+�ڭ7��=7Lj��B^���`�_o�nA��_��}f��y]v�$wTr-�o��ǽ2E���c.2��\d�\ޖ�nz}n9��g���f�:�ȝ[��I��Fq6�\O,��臲x��eSY5��d��b��r���e��1�⻗�Ny�ٓ�����>�N��w�w���;%�^N�*�	���b�ɝf��#^�������#~ِ�h�~:<ϸ�zS>���m���r�#v�I�\�W ��~c�ܘ��OEz�׶H��F�&|�vXPy��g�O����뗖��u��}s}
H�T��^^��[ޠ����e2�}��mC��$r"B���ᢾ����l�̈́��M�MN<���6w:�×��z8�nn��r(Ⱥ�%��e���mCF���q�i��(�^��3>�`D+��׻�<ǭ߮����d��S;$��u�r��/Ƣ���3����j}��Ǽ󑵯|
b�Be��g�v+�b�;�F-sƤ��69����Rci�@�k���`v%}O��X'_���5���S��3y�ʐ����(k��Y�n-�he�=V.��������9�ډ��w+��ή\�r��Ҟ[����;�o�M{4�6g,��ޢ����P����|��Ġ�f��s�:3�>��}�KvO�'�|\���7Yռ��g�{������_�r���'븘W>��+�z=�����K��ߗ<>��髲jg�t����M���L�P�NK��7pB�znS�wј�U�t��(l����
��S�x���iz}]>6Պa)���~�=�5C<qN�w�/���.uQy:^��}~�7���~���&��m{�����?Wu�z��#\�&���i����^59���0�d�CQ%�U��N��a�����Ǻf�~�Y�nf*�9��Fɩ�7�hRt��(�����S��eF��S�W��n=BP۝�2�kJ��
�z�o�m���>^ۓ7�{�{���__R�02!�����}q7�K�kt��F�����kLO�v��K��s��Y���X=v}�wR�g[ Wֹߑ��
߶��G*(�D<b��>��z�w����s:g�2�۪M�'��}�\/��o
	�uHcm�_��o�y���GW�Z��]����Ż��b�7��}�[����<<�,�p�4�.��ʕ����7�Ip��Q��[�i��:�s�� ��+�1'�)ѭ׳u�PbOˋv��>��G]�yJ�󎎭?4����
�qz������z�_ʘ�����q����3���׻���3W��cL*�	�v��d��u���{�x��u��ޚ��>�g��c��E{嵼}�@�E��ȣ`M*�?W���2;��}�q� }����i��(�_����Ox�h��>�q/=~d�=����g�R.���P�3d�ٹ�P���||�vSV��h�Dc^���U���,�7��G�l�>�b� 0���G�U��$���ōy~��o��i�譭�U�1�i9���w*>^�7#�'���(>g=��$�װ]S��x��e�v9��@>G���3�W_�{�\�+�&���z�g���ݷ9=W�����T�6df�	��բ����0��xO�'�l���au��X��-Ab�\���}kTr��t@:Z�۟~N�2�ڟ�"���4�5�0뗮lٌ��=�H�m�w��x�����u�^6�u�_�&��7�Ҋ�Z�o�>��e�2j4��ƌ�~���d�j��;�	���{UQ����z(���gjE}��^�S��=?��mh��8?i�����S�>�<���9R3�ؖC���iV�z=x]���Q仇�i�\Р���3��ka�/h�zֽ+�T�����'��}������E'�g9:��6+��_J<U�Z�����Yܙ4�y������tK2�{S��u۬�ZV1��X���<�`v�o#]��}�Sk�=��C�T
�R.m�h~˔b�;���&�˜�y����ӏ��>����3�ǌ���ӣ��Z�d�/m���0�}��C����k��vK�A���֏5�6l�Tjnc=�]g|@��uG��:b�;�]�Ъ;�Ѝn���y��2s�\<��O=��ۣJ��,fL�˙�M�p9'��x[)���D�`�\�.�����ѷ��z9uJ8�e�6=3@;�\;ɖb���s9dt!t��~��fZ�7������/Ň^���:�my\��}DS7���U�1SȊ��"�`]	�������r�f�U��L෣��_���s
��(��y�;6|��1]��WTcw㹹�;���X�H̞E�mx*��V����2	�=�{��~�\xqZj�	N��`�X�>��Y�P�\
�DUH�{��0�fDmCK)"�u�l��<<��F�������}0����;s/�f=�U>����2=��"c�y%��0�juC/��*=9\
�>�
����¯ң�>�=���G�k�h�bb�q�A����C�V���s;�m;���'ţ����4�j�t3B�Fk�J��K�.fvSKjv�8����Qױ����N��S�7u5:���h�� �_�n+t�Gj��w�`ouT�NL������{nEvU*"�����ġ����)N��|��9K�Yި��;r#49�3>���L����#2o�@U�\<��\����e�v}�DO�{���ǎ�����o9��-]�k������o�Y��{�=���x\�=���K㞬;^f��<o)J��~�e�r�Y���EI��O���M��S������C*�u���V�O��P���Q���g��*�����f��|灚چ:}>�K#���C�P�p���Zfl�zh��]�Q���TQ۝��7�c�yU���Ҁ�+�ůNx���	G��� �u�)'�7�^CϷ��B#�zd���챗��
�=T*0�3�z\��`>@� �S�5�~q[�zT��S�ˋ�1�Ds�k��@{�ܹ�ح��Z՚ǐ�G}�C)a�[wֶ��wp�yb�v���p/U/��8�D7��d�=�N�g~��L�e�x��^�����gI'�J��^8�x�z��&S>���W�pd{μ�l_���K�q���":�J6������ḯ�.[wf0�����{]���d��-�G�Թ�k ��w[�z'��-Ԟ�x�۳C��29Ӏ�' }R����;A��c�E��m9[tC���r�{������^1��Z�����O-�p}P�K��ƓD��H)�M[�< T�:�1��� z#g8�_O�o&X^��xX��ף#�W�^S��K�G�}p�<��w�2��	����JO��As�jϦ��M{�E�^/#f5�v��D>�=�{s0��������ZVtr�X�D�U�6KsJM�&ET�p*.W������a����*2��9�CV=�D�[��)�!�s���o�S�.����l��;>����C�s>�~3��쁑<M�տtN���J����ӎظ��8�_���G�.ECʧF.<�|�����#)�x�01�VM�O�fe�z�v{}�{� �u���=Nb�ʯq�N����w�� (��{�����i@����d�ް�<I�Dm�uE�ހb�:Y,TG/U�Ϥ{d��8~��*��p-z
1E�#s���]�vl�W��Χ�"����+_��*_U�����+sT�fV�2؀=�U{{�5x	��:n�UL.���f�C�ͯ
�K�f����T���������+��������%��E{Ag���L�߻�%��,'���ON�~$h`o�G��in�>��psJ�eYT�;�Ϧ;�ܻY�.�3��̰z��t���pQ�ܿ#ċ�B��p򒉓��\iW"NV� ��7l��c�W]���;��\Y��rۄw]"v�sV�6��vR�n��v9��Ww&<�`�.���Pgc��'i������O�]��7�#�{f򩳟w��} ����EߧB�
�TM^��]mw�,���Ͼ��&-��_%O=02�x��Ѿۑ�gp�O�a�ȪC<2+���#bt��S�:W1�&=�[7��5�uH��u�Zu�3��V����q�mr1=�Lz��L�_t9��3:�=�����,�画����ɝf��'%t�^�i�}�"�Q��Z=��R�u88�gVz�5��w��^��s���1@Mo���xU��^<�8�>����x�x�V�c�nw!\���c�����Y2οI�t�}9F���P(����V��߆��=[��V
�<Q�A�h�a�wN"��O�߆Dڔo= 6G�����E�D�`T\��g�3=Sެ����+3q�k3�/��A߽�l�G�T���/���>�Ib�b[7g�쪑x�oc�6q�ێ�_���P�w�_<��nօ}Jߋ��>�ٜn���z��,���}�s�\]Q�*t{�w}5�N��M-���g	�1Ӻb�:e�jr�=���/[ϝ�q�#c���F�1���c�����1��lc��c�����co���6����1���cm��c�����1����6��6ѱ�cm�61�m����1���1�����6��lc��c����co��1����PVI��r��@۫` ���������8�>�Z�J�JE*��`"����T�QM�*(kET�J�$�T%%UJ$�JZB!UE+M(��QU�I�ٵ���U��l�m6�}��m�ci�#m�QU�mj3fŰm�H�dѭ5�*2��e�ڪm�ڵm��3Zlj�V�6��:j���L�ٍ%��`��4��T���A�Pm�6�kl-X�6Z�Z�)�cY�Vj�Rb��V��31���U�3kXi��V�Qm�(U[SwWFI����M�   3^�.�ջ��/=�zn�=����뺡���A�[���%UZ����]77�[ީ��t�+/�=�ݻ=��O`4z�`:����������fmU�F���
��    .�}V��=�^�AZ����u3W��>�    5�q�=h�;�p � >�����|��=  �_8Ѣ��4z>�G��}�@h�:(@}�}xz  4{�%�k�m�)J��qlm�    -�կ��em�h�+`Z��k���;a�{�{y��S�8�{d����8����7�^���yޓs���hg�y�R��n��:�[ۤۛ�=�9�e�3Y5g\魥��   ��˵t�wJJ�<n/-���m{R=�r��ܳޗn�I{kuܯz�����T.נ�KV���s��Чy��w��֯\�Oe-�
��u��o/b�B�<��A�mXλ�4�J���  ���uMf��ݳ���7��^�^qS�yZ�]����
{����U�x�z�{���%��k��v�s�<�u���Jkg���k�u�-w���Tj�sey㽯Ov��i��{�VRֶ[L��kf)z���  �墨̕�U�Ͷ�^���Wo=%��N���M<�PP�����{j��mY�;���9�Y��涍�!�w��'��v�����^���z.��{�&w�#��64KZ��%��4�� W|;�+��l6;�޲��i�����ww]�s^�Mokn�����kP��������ڭ��z�=�Zͅ�^���S�Euݺ�U�;�n48����U�wg{ڲ�c#l��J5fՈ�m| ��
뮻��k��n��u>f���wm�Y�ڷ���t�'9{;���ڰ���;�m�v.]y���i�uٽ'���C{���{g�ǛgF���i֊���{�u����Zm�6��j{�Sh� ���W��f�3�z���i�t�;�Z����s���4��{N�{QzU�;�m�ڮ��j���޹�6�[��8�G��I7S�=-c�r;w{�{ֳ���7^�63J�mf,�L�jե���  ���V�i*�=���S�e[kpy���i����\��J�^�9{k&�ݡn����mm�f��{�*=��FK�J;cn�;�//m�m����ֳ��� �~!6U%J� �S���� � "m��� � �JU#M �ha�~M	�TT�P� $҄1U=$@4�I���C�/���_���?��V�ʱ�p�>}޹�|��}�K���~�$�	'���$�$ �$�	'脐�$�ID�		w��y����3�}�c??����zC	��21{ȝ(���C������5��Jf�Չ4�-�V��&�A�HN�i��#�vQ{�Qj�@���[�]n�u-��wy�T�ݗ�����),�.�eèMY
��Aٟ\�m�˗O/+ �l��f� ˦�s�4�.�����0�pEh�Z�Z7=�X�g�}I�����غ);h v��mAZ���2M)["�	�
�ET[�!�Bw�X�z�!�`A ٺ��3X���T�Z�+2�v��6�.ͬB�}���*X���z���B�5/6�s�o�<��k~l0
�;
�c-5<T�R튽-^�˅џ-QP�ͼ�vLd��u��#��&��z�p��{NQ�j�`$X�-�0Q��m�yM�MJ5{����pG�]w�$b�]�Q��6��7�\I�r�5�4^LYN���{{#/-h S����]cx�=���m�-ֵ*ө(��b��nʅ��s*IQo&�f-q�޲���	W�e\��r�!�A��n�-����Y�v\-R� $��S*!����iZPoaUD�څQh��-lN�&�+Imf�&T)B�t����Z�Vx.dֵb��2�H�d�7mM�	1��l�x$J�.�:vĽz��v��ӽ�Q���Y�̠� Vh��l�w,a�S��P0$@�O�

�8�;Sr<U"��X�II�v!��3HRf�	U��(
��CI`�kA��)��x���TL5�+n'&n_���P<@!�T���[S*�8��͔v*Jk1Q����YPfM-���S��b����۸r���b�n���ԍ�.��^`�@l����4ۺ���b*�9Y*�{�m��NLu�B1�0kK�]��n�Jn�Z�"�|�%��F� �Vk�[1��J�k܆h���ءJPax�ɔkZ6��n�2#�2�)V/���X��.�e܈},V*�;M��=��ͼ����u�3u҃L9�v��є-e���ܫ"c��u�m+F��$�N�n��4ʉ滔m��[WrD*	{S\�c�į>�*�Kǒ��k�%ޡWO	e�m�Q,�u�-Z�X����,Wt�[��͸�L�ōT`�a�UE(݈i�8Ɨi�^Y�g	*�SL�r�ȅ<���Պ�ì�����XͳR�;�ee��K.
�Z��ܥ��a�2���QX"�҂h�E�̺��M�.J����4FMQ[Uwri�Y�,�#P��N��i۴�Ǖj�2���>��.�`riQ�O6J��<0�ތgb�5&Q/k2�l�V����0��kNP�&ebl��:f�l��HEY(n��M���id�tuS�����2ݰoVK�k73)[L8��h���X����f�ƫ3�z(�VD��.��#��$IRh^P@�!#��+E:�= �X��"���-���.�x��:���鍾Vv��Q,�$>�-�۵g7)nʭwm@&S�f̭tS�x2��DTM#�;�q�&�Q,�]�xsR]����^
Ub3_�"Uo#��n�� �-���W� �d$�J�Ӻ��R�¢ݣd�$V��GP*�Qe�6��4���l�y�v�-Z���]YI�I���8�lr����2�YB�E�b=��N0�2`@i6�3WC�'r�J*еHVZ�d��g2+�Q�Gy�0�7j����ƶ�	�N�w�f�v�"4�9s�:U�4�xmȞ6���KJ<���k�������t�aa�ӥ(�a�@�wV�M�J�uʳ�F��y�j w6�:��B�v�Km��4�(4��Tj��:;��*ӏ����P�	|������b[��ɽm廨�e���ڴٹ��S�V�G
kPVS;�3$.�:��/5m9���j*����Y`L %Mf���Ju�]���ҬbXx`��0��
��ό�/m�
��۫�@�b֚Zn["���\��Y��h�,dr�[�"��yL���5.��1�h�5�zv��ЖɱfU��V�w�"94�'�X���E�Z)
DµwP�ح��R/5��;��S���ת��,�AN5���0��I��&M����
���
ŵGi���֜.�U�����w�R��[IH� 0�̖�
z�MEO!�Sv�a�Վ�j����5"-�ctJN]�eB��v�̙�R�F$4Z.\X��2� ��,XP��=ܳ�[��-�Z�@Î��Y4m^�÷6�+=8C0&�`�z�����I� �f9*+�͖�M@X��U[յvp�+iء�����jRm�o#��
��-I[z�ek�!p��YAc2YW�9v�V����{/.بv��۠N���N���p4hk�Vi�V�[0��$�jF���c���a��+Mh�aRj�71���n͔Z�VlKt�Lc,�b�b;��qؖ�X2�S��H��E�aTQ,�d�ӮSLGtc,�*(�9�r��yMҷ������U���%`	�:6�	m�)��p[@:�h�Z�M�q���NXtujE8��۱ZGؕc�x3�z�҄;R���-P9E۬�9p�Tr�ti����Y�SIR���@���d�)�9dk���r
�D7���!��lrե�*���#���J�M�f�j+���1ϳ����%�<�0�Y��+�6�T�CN��wz�i�gS��!����e�N�yy!Jd�y�V;�WE���F)ƥ�Pxscb�ێ����ɒ�����2a�C,�U! (e�t�M�,�WxF��x�R��f��mMW��&U-0�P\�U 6��jKc%�C(륅\��NJ7
��7oX�)X�bbi�lei.��v���K�2�CS��&��;> �Q�i-ӣP����'I�+7{Y#�r�J#T0eeDR<�u1�͂� 1A��a�Fj_�7l¡��V �q�MZr�TЭ�o�ve�j�����aZG!q��P�J�r �hXr�ͩu���+�.���[[�;�᫒̨��Պjv��m=L��V7����H����\U>ɕ �i ��W���k/*�j�
ң�JJ�?���(��WN�]�ᷥ
����5yALt6������'q&�S_f��z#�m�Y8'�n�ܙn<�MfԳ��ys$��H�oKu,�%-�0��*<)S�P]-�"t@��൛���'M�r��%ݽ�c�]BtbZ���hiʲ/fi�&�=���# ��i��7ux����^m����1�&�i�v�u(S��}����6�6�lZ��Dw1�`.���*�2��yUn��b<z���B���˫#]^3��Mv��Jθ���ѵ�MK6� -�R�ҡD��#ҡA���V�n��of�	��Ą��to"��C��
��)^�5�Gy���fc�t�����+��R�>.���0�b��Hiv����V�Ax��Z6���^"�Yp�v!6��a�I��Bmln����|�<���˂�b[�+U
j�h�u��JsI�)EM�p�{+N D�ی'�5ne��L�z���.;Ö�8^f�&�Ym�V*�14���ݽٴ�+ z)ܩ^k�f�K[X�8�P�E���h:�������^[�fÛE�ڈL2���-�P�BgE�QKj�;����op![O!� %�Z�FlV�b��`�Z��r<8��C4�ѽ���4��q�&�-�Y{�L�C|��@�V,�ks1ֹ�r��V���Z�a��=m�SUè�e�JN�t���V��S"ȶ��t�Z3���-��t,u�05OX�Gؼ$�c�6�
�"n�mJ���
6�f��c\��YS@).��[��G�a�W�$�;��P���2<X� �GLT1�ݶ���m]XƂ�����@^a�0ZF+��b�c��Cj-iŎ�}���6!�S��vF4˽�`*����� �K�SX5lTz��XmJ0�i�W5y�Vs]fZd*�Q�em#W֢yG�Zek*Ŕ��VUʒ��Y1Ч����̹�0J���6%"��˧[���!vj��GH��zѕ-�0엨�!l���d�[��͕SH^eiV���i��ԩQ�wY�m/�
٨df��<�4�-d��Z�0�>Y�2��Sb%�H`w�P��Ԥ�M��v:�*�q����hR:ś�GU�`ƞ��L ��K��(ƞ�Ѐ��`V�V�:)$���Y6����v0��ԫ�c0dkNFnaӚe��k$%Kf�J0aY��;A�Ź����VΫb�<�f�:����B6F��iP]�xH�u�B�"ڻ���x淘v�W�\�6lMn��5�襔X�f�D��@w@�)�
Ե5s1)�����S�m=!M9-��e덝w��~y�j&	�0�K���t�08�Q������ޙ,�Fچ`M�:���蘚X��j,�N!Yj����7�B{�g,CO6�Ԩm
#P�&�f����H��R��Y2-&��qYw���:z���mݤ��W6P���[�VR�t�q�̮�}��:����Z�+,*8D��U��wz%4��҈�7L5���a��&^k��A�zmf���?��W�:�۬�T�R^VL1��ؗ%hw��km�˙+M7��ɳ��#BM�������T����sJu��ue% yb��{Q���7�B��j9���޽��2�mZ�.j��q���2(�j���e��3L��և9�1��ra�p*F���Á�M�V�܊�'��5V�/5��l��6�v�`�ˠݕ!%�Ԇ�V����-f�3�\%�ؐ�ɭ����NdIӊ�hb �A�X�i �`@�z�ӑMw��HF��5^��μ��$rT�y����y�I���1���y���(�x�u�]�L^޳3*F�s6�.YȂc03eC"��)b��F	VD��Vu�f�p:a�r��Kw3j��2��P`��T�(�T&�MTHz��!�i:�w.�߲:�Ŵ��/��Z�b*A�aU����XwP�$�Țɛ�����Q���!e,�cU��3w2��n��)=��Z˸���f�KiH�)izV��{��-���gC:�sH��r��Qe����(�$`;WQ�zn����ǥ�솊P�B/ay����u�,�"_b̭��@Ywkr�d�[.30VHC5b�el;��^�3�B*;ǋ2�D�M@Mӂ6m��ZW�a��T�q��EG�Btٳ��dM��V������
� ���K)jl���E"�eI�{����*�e�81d�B��5%e;��l�K�P*KoE҇m�{u�Xs!U�F��8jS�F�UlC ݗf=9X1��B7H��&��8�U�衱��9zk52��2�X�3ʖ�9�Ӡ���n���A5�Đe�Y���oo4�%ҡs�z��=m'��V�eE���l��W�=��N�F����t�Zf��ND>;�TX�,�]3��Ji�cF��P�����`�ͽ�u���%C)EL�n�w�qk`���G[�� ĩ���D���
�PX��in�XUۺ�Ue��e�)*�Mj�ki��Yr��^&��y�(��k(�?
�\�P�v�mU�KB;�A0U�%<+P�NRGR[�d��]fǯ�#�4��ʌ%�S�˦C�C*X�����WqO4#��iJ�/�U�:���
���l4���e�=�$��"�1j�M튆Խ˖�ivZ�f��뽬�a�P�!�JVu�b�����;ͭn�~s還�Bc�ب�IH�>�j�0�A�^�MU��H�e��h����3F��@Q����d�h�DK"���5M�;�Hq���(��M�{(m�VZ�#��=ה�SM5��F����/U������ͬYD�*OYlme�\~T���1�wi��V�a�g+un�0�	�ň�=֍��lY�jm�WS��X�ԭ��	L�<��Jī��t.���H)����ügh^���En:Q�[�M]�ʾ��	�}dY(�wRT �y[�2����d��D�gN�ׂ��Ǣ������+^�|���z�����YW/�dm)I�Gv�*틤Ҳ�X��8���i���V ���B+N7�&cն���*�e9�#.���Aֶ�R5�<�(]ɶ�{l.��M͛ /�=��Y��0�j�"���qMѲw]�*϶�{t���2J�6�J�%�XaBqj��t��ʲV\[&Z��k���kJ��n��r�%&��Uh(�6L!U�CH[�����{pn]�
ɼ����;W3)Mz��f[�fR� �vh�am�eF�+G0b�m���-�˪Ylf4aѨa�,$_�{���I�塢��U୨����`�
=�[7�B�mYV����+xr=&�t)�tP�k1*�,��6Tq���ncè��"o5M��ʖݰ�l`ʱ{��e��9iM-5,�0o^��n�4e궤	[�J�̄�`N�+SŖ񳤝/8o�ŵXE�ɦQUm�G!���#��2ⱳV8�ں�`��-�l�{�n	��P͠�)0�@ ����Q��f��ɕqVQ1m��V^���l���uyDZ�/n4BB%+�J��;��ݺ�����5�Ecŭ�֫[�K"��Cq��
WH*wH^] �����ln��8�R�Qۥ���䌙&$��9�*�g"D۰��CvL4�E�b㘜r��D���PmN2��Y�b��E�qIW��@dX��\�� ��"O�+���:j���Y�d����a��{����&�Jȥ���5ɻ{A������˚�8D ��r]��+)�Ι�]��i��;O7 �����4�:��y�jN(�Y}�W�Fէ+'���kU�&{]���v	M�C�fu�*4�_>�T��x�V��2��m�j�83�!�r�AJ좖o+}K؎fRŤ���c�;Nlw6����e®h񠷒(lӉl[L ^�s��d$m]�aZ�ƵL<�*a�W75Q�
cY�[ kp�����y��fdG(��,�.�S��k��P\>�I;�,a���P���:��A"���f!Iۭ�W���4�\K�I�
hNY:7O%��5>���B�ӳ&_��ڙ`��2v[&�}�;4a�;�����ڛac��L�A]mp{}40��"�Υ��{N���L��)����:�Y��G�ێP���5���j6k���
�e\���;P��ܡDk�p[�_�Q˶M낯C�tj5� J���n�l�#�=�Q��I����7a��pV���F�;�҂�0Vvm
��v�Ut�Ԭ9��0Iz^�͗��s-�	6��[YwA\ʣ�rY�cy�A� *�.������ym	�V%b��uޜ��iX�[u�u��T����umG�S�c1���9��#ZT���Cw4&J�;��c�}�2٩Ƭ<7�����֊�'Z��Э���ֲE��,�����e���6��3�$t��ϦW<=��E	��,l���QY��������Ӈ8i^wAwR�v�٬��=�z��'>�m�7���Ag_TO�i��5v���T�E��ӏ�u��Ph��_ْ��;n��լVp[�Y��ch�r�'����_FS%K�ޕ��i>���2�휲�
ȱ�b�_c�^~�Kq��{'�Q��^g�r�] ���;p�6�tJ�@w��B'(�Nl
���]J܍v�ǜ�_
t�űE:�D=��v��Y���eC|���$n-bŎ�,E+^�B]��$�hU�i<�MM����4o�F�N.룵Ѫ�A�:�a�2f mqH=J��@鎎��:}@��v���/bɮ<S�P��jK:��ɤ>�[[CYB�Y5S��#Tְ(�vM����{x���^x�3�(�;����J�w��v�؊5��*�a������k����y����W��@5��֎r��zV��]ؔ�V��Pǔ<맨�Ɛ���V�l�)H�������(����+����p�g`�vu!�)��A�U�6�C�j3�P퓰:T.�����6�ˤ�Ku@-v��y�NX�1�&E�u�yhk����T�t�s;�9{�\$:����B
Fe81 j�8��2]uDc�Kr�s�0`k4�.IS6;�k�ӣpG�Ԟq8��sK�ǻL9�c�x��dؕ����k.�3w�sh5J[���ε��$2*�7 ���4b	d�uЊ��o��3dA}������:d�å�1L�9B��."�&v�`�:��z�+�5��x˅NWǅp�SRm
�D��a�n�ޚ�_s�L�Zv�d��!�c���z��1�hm�R��hw�P�9��ڼ�C�؜�l��ҵ���V�ǽi��)�{XJ\�����R��ox���b�ʵē��=��)C���-�FG��!*�_�a�8���q�Ia�N��]f�K{��J;����u��v[�@M*t�
Nvf�H$���nt9�/���IGy�;]�r4���a�B� ��#��5�"�ub�lz6͙PЬ
�#���6d�{�����S6q��
�Dܹ�7]nf��iE��F�K�W(h/>Ob��K��h�jך��� ���uo��2�JT�+�����}��a�k1��̥�҆.J�ź9��ʴ�h}	�ڳ,'PYۙ���
�U]1� Ļ4�orc%�f��sS��YET�T�����^B�M�_K:"D1��L�U�g)f+�h�f^��Qά9T(��ȶ��d\�9��PZ��������8�k;+R{[.�z�Z��&�D\$�x<}�d�$l���)r�)�Y�\9WBY��f�#��D��Z{�z�0�fҫ�n�7C'	])�ulU�� (����Y���t*�'Z�X#D�6�p���n��0-�(u�7��g����;H�b�vV`�Rؙ��i@��Ğ��a��3���2]v����%3��
W	��n���Xo���yN�oV���pB�vq�(N��+s�֧[�D3�oK�����.1I̡J�M;X�w� 8E��,Q�:���7� �8�J�d�w��̇X%+՚7��Y�[���Ğ^o�dz�
�PPu���e�f�h��
�̰��|0�ȋ�Mv�Ճ���oj,�"ShN���Ģ6*(׵ږ�p�8i�D&s2V`���� �t�.��S���
J`ݬ6��\Z���4�}�[�b�-��� ��n�TkZ�`Xov�/(�.�Q�ݑ���Vm";��!�G�u��O{W �M���m</w�VK���	��:�r�|���L��:���SY�k��b̀W_"�ט�.+o��j��+����ԛ��:'�Z��:[i����k�xۣQ���S�l_7�f��9�\��zQuJ��^��\*��?=cl0�+x��C�vV��-4݉��rŭ�{�I�YG��o(�7�6q EgQ��!/�9MqO�N�4�_d��$Tx�c0�b��i��Eϯ;=J-9;0��b��+^�����x���Y*�6<��=;*6Ïo�B+����R�9Y{7}�Fн�ªf=�5 �`���"��s��c��=k�{�[�Y�⮳�˔wz�	3-�b�Muy�k0��T�K]n 2��hJ��*dѳ�]������;���2�qd\��ny���Q��S-c+0]�V-��- ��Y�MJY����Pu ��J�Kb�w�L�6��^�����v@�L`��c�jZ��%s�Z������12��N]��6�Ӿ��+_Ӳ�)�6uk�\�B�<���Y���!�vn�Nۡ[�����z/�tw��W<T�b���Vs�c�$;�xMh�/tB�>�0��Ŭ�qr��u6�>S
f�Q���)Vl:�&ΐ�Cgj��:WWNV�!���s�ðQ��Kw;G������ӽZVr(4�ѽB�����d��ݽ��R<i��[�
d�jŪ��j�=O�`V�b��n��c��嬵8`�D��o��eeC����R���u3�&2�f_i�R�;�L�xY�ޫZ]�ALM��N��V�`2��3eb�8q#/�U�׶�Y��c2lY.�bq d��S)�H�+	iuah�VN�*�����R]Ҙ�)N�W���>�X�|,�ʳ��K(L�]����h���v)*������s����R��u-�=Xyt�)|m�5��a�swxV��t�T�I7h���=&�,ǽX"D[	�-�̀w�˕p@��d��O;�����%��.��M�rp!�R����bΡ4�5�;��nIJ��#qݕ��2���)c˱��z�.�@�NKe'��j�b��N�,N���z�!t۾���t� _ru�>�k�����2M��f��x��uG��^�h�M���c�c�vhb������6]n����Z�A�7M0�� k
�G0k��.b�eǍ�h����#�W3��9��4��u�'چ��E��`[�ҊN�)`zrw���r/�5%�:³(ǣA�!u,�d�lop�p-!���ђ�m�y(�1��VRU
�u�]��d�������s��Oݜj�gM����M��ILh�����[���"���y���"�	�7�� ^r�@���;�]���$M�� ^Q�#9NY����HV�ˈ��)_P.}�Q�7VAW�	��+�o79
#�7��������۷@^���w���I1�+q�⮺T!%�U߼k����%uj����6����nT5����Rm�� 2Ƹ�ړ�U�Xŏv^�hӖ+�.\bZ.�gf��:6~���u��#��Ef}v�Ҕ�ת�3'E�[�Xa��YѴ{w/8��5ޔ�	��W�77-�Y���V=��u�ժaSj��2�����''��t���D�k;i��	�Sj�\���!XW_�.��R]h�rĺ�R��n�h �y� y�
��]$0����{;Ϟ�.�����.�ݢ��B��l�)�#`��fə�����;'sS)n�)��K��[�"˥*u�&��E��=}��� �d��cB9�n�{ݗ�׬���o�F�h9���ci��L9Kv���ʓ)e�S�/R��s��L3X]Mݱ%�ν�諙X�RO����RX\3�XP�j�J! Ȋ��� T�!��'=��-r[f�G�uv���ayo���T��A��-9���D �ڝg����9e)`�<�gSO�6���u9x���v3[q���zҹ��<����+�:���j�M�i��������d�w���#���R1۳,C�YŦMAt�xq����`V*�1����.�s �7�����-��NM�	��.\@�c�j0�����F����=���#�e-�D�u�7��N�'{J���AE F�U��/��+�4��YbI�2�v�c	bMR�Z�dV�ȥ�m
|p��*�$�tٔ�
���\�q��s	@TKiJiZ|���,A��ޝ�Te��`�Y{�|i�5�t���q�y��b��T���9��(�T����t1Z��B�hnp��b��f�ˁ1�Y����������n:Ѵ�*\�Uɹ��R��emC�wDs��%Ǵ@��0W��q�d�jM����;�����i-����,�:زuEa�QQ����Z��;x%�cy�n�g"�g$_Jk�nlGT��fЙt����d���<����Y��!��7ë'��p�^�3z��e]�Z�e�P�[JDE�(�ol��v�)7���|�XOe�nS��/!�&��W��7���s�%�i�����;�$&�]I��#h�W�nLd�)�fձg�%w�D��)���n�}�r�Cctx"���
yYJm�󰾵��r�f��۬�;[\:k�;8n�E���/���ҕ���`���YxN�4mr��5�����5ڨ���0[׆;y�JG�v�h�.͜��[�w�v����#1V���6I�V'bc뱒�F7V`ʃ�V��Waj���"痁�Rc�L�w&���M�FlC7�$ޫ"id��|�Ҁ��u�%�����p����yc(��+Yi^�	�	�a��U��F\A�T4�={6c�2^pF��u�Y`�T�U�����Z���:]4K�r�6�b�"Wn��8�_m�j�Z�C��b �`�ы�_c� �nln����<;:��׺fD�a
�Z;;�Q���|�:m�n�ulUv�E����L��3�d��d���`�׼+Q�(��)��o7������کHL�98��]k2��uv���(AǯO)r4����&\4�!�ݣ2^bԶ�VesI�}vƈ:�6U�V� +��"�]��8Z!��쇡ȍ,2l,[X2y�b��E����٭�=��1AMQ�W�d�ibZ1F20���p�ga�ww8E2�U�S&�-;-N���sj�j˵lh��o7ip�ݓ�9��hʙvMs҈�>M6#.���'s�@��x�XA�Fc����O:mfQ��^)wH1�[�j9Ū�}�Eک�wVE}4��Sy 	:���eZ��07�v���hW�ه!)�23,�N>�A����W�<"D��a�;�F�)]��I��;��ٱaO7밞d�Ebm��N	S<ur(M��w�$���Y[�P��0۝�}�)��nJӎM�hn�Qz�kqd0�m�Պ֡�Ͱ�㵇!k���k�7:�VK���j̝�;�P�Wi'DH�����Һ�,�1/��{�N)�2s��wz���Ok������R�f�wR�l�I��«5gm6���9�+OswV@�]�c�:�VH�Gp���D�X��}ו(u�8��xL���d݉��� �t.��f��	M��ؖMD���Ȳ��U�U��t�r�sn%D��`�J�2�f�H��Ӡk�^3�B�\3s�ev��B���3.�M.ْ7�s�e˻���e�x�r^
̥@M��"�b(� 9J�=u��b$�ܼ�1�����ا�1�{r��h���aG�s�z��c�v�=4�ڕ�k�U�HoI����;8�V�̑�2��Y��u�(m�V�ݺS0^�v��ώ#�dt6h�q7�i�?N[�M��)�l�h��USn�Eb"�c<1+ǔx��
	�YD��K�$b�[:&�.o���n,nO4�P��iΓ�f)�u���iY��i�1Å�3��j��l�HK�s]�wh�O4�:�/��:vH�@�K8p�f^r:+5LD�C�̮'��;Ob����k���C�dŗ�B2ޛ�ik�64�`���8��
�j�{w���}t9�A=s�}���u��<����m H3���#��B��Y��ҡ��W4)�!A%�P*q* >��v�$1$v7qψ0{pCS�iýܮ�p�ױ�,Z�m\�� �J���O2j�!<��w�TgKɽ��������m�5��[
�"�qborV�!���-Y���o)�p�Mw�wm'e܍��P-VnY��O���=�y�.���,A-F��{�i5u�b�R:`��k�4/�͖�G���-V�ܩ��)��{�&�pS˘�����9Y#�2p����m��(#�7 0g<cY2���7:��ъZ�v���vw7�<z	*��S���Ia���w�Đ�HH~�$�	'7�cc���n2�'#��fJGu�sa��eRBT"R�{�IR��8
YZ�kgn�����;r#�Ő���X�>JXǂN�X�x �l�r��S����}6U����.��^�n��Ƈmfѻ��n����N6�m+��m����tW���X��g$��#ˀ��\y�2@Ɗ<�ޔ'�ʵZ�6�u^�ec��w&ުu%K:��{i l[V4N3*Xʩ�o�Sڵ
=���� �u=�𝮻��_�Cwz��t(!կ��4���3��r}��s1Wl�a�ɡ<*��TTAe��z���'��Ћs[�����Xmj<�
�������[�z��pL�V'� 3�E[����50l���f�w�퓩�0O*+��Y�<mV�td$��5��&�mn�Z��-��WBơ�pf��H6�i��ֲA��O��N$ʺw���Zn7�E3�T��͍�+U�{����n�ŧ�f�#�i���A�q�M�Ȯ�t�����8�N�d�°�ʰ[*�1���<D�e9���2\��n���!��9�v�;㎻uJ|�Kmt�)ŷ&-�3 ������>V���o��F�!��Uj�����u�T�5�K[�QH������Q����\OzS�#a��^�sV�"f��8)�l��,�S!{�@�f8nM�mY�8mI�����.�����)��ھ3v;��a�W;׻p��2!؍�^�j4Yj�)֘z���<���N��Kv�4��Q�V(�ap6��M�I��ypB͆ڷ���	�I<Rq�PV�q��B��E�(b�hQ(d��z;=E*�s�u�[\�5��Q��xvo���+��4��2�PXyx����ŉX�t��[��.Kr��<[*���z�,��nL�7�mNxQ�!طnܮ���A��D|��H�u��T}B�
#j�&�P�M%��f \�b�h"���{��p��J�Aizu���N��f��4sYe���mݶ���v�r�����f9�h���Ee'�9Ɍ����tIK�B=��̵I^�"��yش����{f�Q����:܍��A�[F��t{F�U�3�ǳ�0�[�DRtN/d�5P
�E*�S��;�2��@Jԣ&�2|*7u�]`��P�A"X
0p�7L��_=��W����'ee۾���q8*�"B#I�1k���:OP
�`�!zrp5c�چK\��B��l�3s!�(�/�@���%���z݇�P���ڑ\�X9��
��!Ö���\]�yS��u5�׶H�+3)f8�] ���$QYr�WL�����j	Du�w�j�S>p�ӡf֚W�h�����@i�
�g�ir�r5���{�]����9ܙ6��?��08�|�e�DT�ێc�&�pT{E�5���s�e�ZYX"r*��c�c2]<�COR=�ڞ�(��3�kh3{�w�wRP��{0���ʹ�t���A��.��J�qhm�]�Xm ƢH�U�{0`�ɳM��*�ءǲ��[�]��NR��Uj�Í�J��,�Մ�p�u���	KU��Yx�0^m���t��7W���^�H�J<h��C��9τ�_*�)a;�6���ර6&�R�h�m�HYf7T��s$$�~�?kF�*<�.Ԇ?�p�5�g�Jt˂�j��`�`��V����䐭�wL�L� b��[��,��b�+4���}�qe��Վ�&J.U��繋f; RʶhU��0E����E��)M�T�{rX�ήaΨ7��1x%��m�G��5�P��Kc�P�j*t� n�1�0s�*K"�6!jo�q¶�*��ѵӣ�bͣ�."�˳���n>�V�*�⩶��6���,=��X���FL�̣��-�$y�{�6��B3��rK)�H����c��%�9��w7�u�V�me�ʹF-�e���سg2��.��6̲�12N�SV�B�aS��W�'�f��K�qJ��.p�	^�vcӪ`�o0=����#�֦�-Rm�Hqv�X��Nz��%��J�:ϛ"�!�Ʒ �I����1�PA�����J�1�YE���4��p�s.�۵e�9Uq`��h�]v�bER������ڮ�xJ^��]�/�c��9�lO����μޟ1d��Ƭ�m�Ǚ�E�@ԯ;:T�l��
�7M4s�fS���i'B3F�vu��k�,V�1\��G�Rml<�;Y�����V����{|U3��V��m�X���,�Z�8f=2�^�ns��Ao����Sw�)Nׄ3Wcl	J�y�fLZ9�O�e�L�
���kQ�Rp+�ǰ�K�u"�����u*��˨3R����e��\�[�f�^&+zMF!��f���[š\��B2��ېW�/���SS*go_M�L�K�#v�A �6V���r��u�J�g*�-�VYzO�`���|p�k?�5�	*���+o�]�VJ��y���40��ד077' �O�C���SŎ�{�'mC�&h�7�vT�v�b�7�ܘzӷEv��'�`���]ѕ�B��`�/(#D���Ҵ���yRR���8o���6���J���� �C�TEǵ�CѼ���gjumTOr�}j������ox��a�[�T Pq]���6i�y*�m]2�]��ak��x� I,�to(��l#62�E������t�`<ݷ��ۻ�\1�d�_�Lw*G .$$ȶkxv�>�2wm2m�]v�
������zq��E�ij,���󺔾
Y�B0x�.�9Ql��<�wL�I�e�v��>\)
�A�{#Uَ�;za[BWt�d
(�a�i��
��;�"�<V�.���`(�:�5j#-_Q*�Ʊs}I�^�$YZ��P�枭(F�7[2�c�*J弻�}�ky�� ��M���M-���6�^���m�+�:�$�Uܥ�@Q6"ol��IVԩ����u|^]
�kc�����W�2U��7�#+�3�y�8��zkl����5���v��M������+$O{���Z����\.���d�6��E!j�-�1�ѰٟCX1���p�/�����X�k�	e#�-���ی��w�o�N�PAeԥ����5up��_P)�Z6bs�;6�Ǧ���gn_V&y]�f����`��"J�	A|������j��dR@mԟ;�wP�'������,���U�EЋu��i�h|�����kt_Z\���u-�av ���vs�visU�.�+jeeB�����{�n��K�����h7�ZlEm'����q��d��bb�oAq��b�ȭ�9D�U��-�GR(P�WQ�s���O�2��)���zq��O�2ͥ� ��K75��VV�YW[ju�:\�*)X|����}ި�M��)�;lh���8We����y'�ƚ����(�.������$6��a���`$.�,�ѩ��p�^��H9Hǌ���]*��\�e
���씲�*Zwt]����.bzF�c��tG�+2(���Ո��/2V�ck��>���MڙL�ϭk��H�(ڛ@�
%ٷ5h��)�|F6�ZwvZv˰����̦��H��Zad����V\��˸T��v�:8M��R���,���6�T��tyԃ7bGw��+Q`w�9�V�6�##ā���w�*WET43@������b��1��X�m>s��X����V��6�1���P�嗈n�C)�eTR���������jf�T�t �T@QHZ:��w5e������Q���c�\���y��to\J�)�;��ܚ��b�[Ac�f=Բ�i���e�e�Rn��9R�Z)6���D8��yIA,Н' $�n�K�*�qW"��tq�*��
�+n�[Z��/�-� �6����~��rt�;�u���'�X�JcB_o*���1�k�u��+���2�BM��6��.k�ƺ_j�N%��F���p���r��w��[�m�SIi:ڱB�'%���`0�����}s	qU���y��C�t�����|�'8S����t�lmj�Mmr�BTW�0P{��2�v���p4�v���{N�� ����|c���*�	wѶ�M����à�u���`5|e�JLn��h��f�{4�OPR��Sr��K+L�4=�6��uP*̉#���T�u��v��]�
�e�M�tӸ��Q[��w2m����}�`	�Fƻ��Ҍj�E���C���� �.rkIy����ά`K�r�h4�5������&�=�)�[�h����ԤSkz�mĶ�j��j�� a��}��4����*��i<���8�E�
<�t]�e0N�K`�3i,��mK�Y�U���{����"0u���S���c�f9�j�1���+��K.������V�pk����8w���&Ww	��!ɾ��s���O��С<��Lj�V�!�(�����pS�]|��`��jY�^� ������c;9��B���J�4�T�7�iu�5���k���lP�*`Nq�}�:ZN�4�<&�S���8�����*e��8��Vf��m�DX�J���lE��ή�?t�A$��o9����,G����EJ�>��@,�����zI��;wr��k[�EQt��ЩJ���!y�y�Tq�P�lDWom=y��]m&�Y�����:8=&U�P�0��zNW(:�*@nL	�����G&���L7ra� C��aĮ�YmwdF�f�c�ä;{w:��jau�q��^Z��l�T�`�4���
�a�����ѼKYJ���/ock^��r���VV�q�Rk3:qN���=A۾���-"���#���ܳd��;�ro5��Ә�,���{��-�v��(Q��&7���ǔ[�.lP˽�M����6�*>��F0P�q��5i
��sr�]��`8y@��X-Pp�+�U|��@�))�k��"��3�4n�y0�w���'J��r�U��L\n��W6�.(-E"y�� ��G�N̓�A�Gb�;�ȴ\3BVI�4@Yޔ�4��3������R
���Ȝ.ԋ��ю >�N�Azd%���_���6���A:"�v�l�\�r���|��v��)i��h}X虗A��A�1�Ӌ/sl *6fY�8u�1=u �rإѭ�D.%.�l�]��l3�a��i7/��2�����Ѱ�w���6�q �2��o�&1/p�L�$Li^�Q�$,�qQ�n#���ԕO }�tuyM;�OP=�	J�rv�pQf��'�#[�Rݜ%�)��u���� �h<��YS$u��cE�48?1XhC[��X�y	pI�um��F�,�h�J[6���ni�[rpK�[��5
�6�'b�]�^z��C;��ƁZ��K��-�5���gD�ȫ�A�g�ݖ�n�G'Nm�|Bn���J���0v�	ij](}U:���im�S��BQϵU�8 VBY�{�ocgr��B�������2��Akl�?��ݱ�չET9H���F�eV�ن��[�#�8!�$P9���Z���%� oH[ܤ�'k(����o�M�$�`�zo���]R���\���[f�Zۋ4�{��J2�M�=��@n�ĳ7�.ӫpʎ�%q��XF���#6�Cto�DyGԨ�B[u���a@�
��cZ�H��ж�'r�2����̓
Tީg���AL\��!�r�E�I�wұKmEf>y��Ϭ#l���e�y�w��wbf�C�V�m��PY9\�.�Iz*#(����Wtq� \]۔[�h��g������,�s��p���b�p��Y��ޏ�taxW|�Nec�YV��z[ǀ���p����0(��L�c��N��^f��Ƴ�I�XqZ���,�����\�?G�Z��mI�j���N�2�T)1I��rTN��P��qj�<�����S�+���(���K%ȳ[���4��m��Z��yk
I�k����l�|�Z����E��|
�N�"����3k��X�е|	5x@����F��}s���:��]33&�+)��lz����71;lv���	��9�N��WƠ�i����QT�5*�RF7KA�\}��H�M�9IOSt)�-q�Q>l䫰֛�7[�h���R���1k�I�e!�V	�nb:cj�@�Lz)�Z�`�(#P
gC��1YU�R�WBS����B�H��A��F�g��4���2�A�/��b%�@�9hvn��*�j�߀�kH�rr�滾M)r�ҙѬ���1j�dte
��[�H�K��wR�-�X�,��b��z����yB���L	i��U��N�OA<-@]��O�!k$%:�Rn��&��f)[�p�gb��`VVO�>�tM�R�kQ�5n�����!�I�Q�4`�#��b;���6�⼷�n��^�yܥFA�A;���>��[�k�I��
��T�`�4 ��u����t�n�t��:��nc�D1�{KP�ҡ\�[3*RP^�#�Vm`#���B���QtE��)ȓ��v���gL�xN�Ȱc7K��8r���d5���:}�#�+!�R� r�f$-�6�u�Zu-y
����1V��ڵYw���vcD *[������U�cbϑ�bdQE�vZ��bS�s��J�/+ r-�9��[�h�^��w#���������|>�σ�q)L;d�B(���P�z�[zī*�_�r���|nt��I�e�U��N��7�)+h�j��di�m+�A�"�B����,K�1Y];���ͫ\x�`�K�r�������ة�n���*��jc)]X^�Ɍ����.��t�L�x*$.x#i�ݛ�5	�Q.9L�<��Q��Z]u��/�(�F}��Ƌ"���h�y>3v�������m�?V��sWקa�4<h�4gbV�D����δ�v�32:���~Af�˳��1�{���U	�^�9dʏr=�Ԝ�h?d����d=�{��v�[�<h�n�h�Gj2X�H�]�:1�SF����d=�U���V{OT}���&^xC0�>�%@���R��ko+�è��=dGPZ�i��J��V+�w����'ݪ�s��i���[~pvSJ٦�҅�G����(�����N�-����{��t�=%#�E���7�(C��u�f�=�`�R�ȨG;�%���ݪ���j��]׶"�&Xĝ�p��i�z�@oX�2�.�
�˨3���2T	�O��Q�|�A�K�J�up%WFJ ��"6��E8�,V�0�J�[��ɓ�ή�
�sXʻ�׏P��ۜ.+����U���9m9�n�w2(�MjU�g��M*A�v��F�jS/K�s�J�V@���	uq� �KZ�w.�#]��j�	����Ŕ�O'd���{x����ЩM�P^�Q��E���;[��[�q���{S)�e�Z�U��"�DP W�X[cH���Z��֢�&ł��b��
�!m���+QW1DU5PUb0KBѵ��#�PQ�V�YR�QTF�QU�QQH�F,Q��UQKF	lYY1��*,F#(+Z
�E�+U�����ֶ�ͦ(ڨ��iDA����EQ-��R*��m�id[J�*�(�Q[J��-,dL��b��TQ�EcQ���UQ"[TEX,J+[F*"��U����1Q� �b*�UV��)A�-B�Z���J��F5�"[F �Ub�PR�UPUm(�Yb�!mQ���T�b�"�����)TAUET��-*������*1�"�E�+mJ�T����PTF*�(��
Z�6�#,(���k(�@X�0��,QV"��F(�0EAb[H�
�UX+����+*"��QUEZ�,PA��-�X��eb��S1V�TQUF(��A���(���*ё�ѭoթ�5�nj�u�°��	����n�²�:�R`���c�K5�k&�;�vp��G�2�d8{�L���Q�y�`�����D�j��&��ר_h�}�5y��Os ����`�L^"�{1���)�yq٫���Ϛ�^�`����0,�9��p_��t=��K׶�g�����!h1�d
J^jY��fz�t���`Å�ø�澫���K��ה�>�m[����ALDu�׍���`*9�ծi��*�Z� ���1zx.R���q��]L�'�?f�:�����9�A�Yض[�w���/��(�.��������:ߵ�%���>	Ge����$%N�<I��9-���I��'���=�B�s����t��f��q��s�s"ڧZ��r3Z-ᜁ�C{*^�����d��W�^t�\��u��==���4jR�ni/z_�le�n��M��}rm�)T/'3zu�ү~���nfP�MK%����M{�ޟDj�4��`M�e�d�NC�j��ē�7s
��X{�i[t�Ss=�Y�s;	��ߏ`�_7V�� K0��,��q��3w��N�f!E�׎��%�Ó.�6ݧ��z����;2�4�N������ۺo8���p0Û����ގ�S�
�v^Rԭ׮:ڣ���6~�n�ǹ�h3�_g������@�Q�ԟV*����pɞ�u�/*B����7���s��k�B>�i���z�Wk�Tx,�py]㣽����.�����C�������^�5���Lg��ڍ1*s5��-��̏6ls�P�^v�������d�o{>|"�o�\�8`�]�]{�*��V�o��ر0s��&��+r|-��?R���\��}z������a�A��XW��ɋ|�~�A��W��g��}���b�z������G����dW��x^6�&{��4}�s���^�O�q=��mqןL�ښ)9��h�T�D-goGg�W�7��<i'.�\�xL��R~+���<�������[<���;���&�QJlL��x��8J]q�>>�t,z5.\�i9��b�WkL:��)e뇓��W��\��V�ڎ��$�,��/gT8/�N������3���n�+>����+�j�J}�0�m��`9�L�0�֛��pV�W{���̜�VN삕A]�wq&��K�^-qZ�t�)y���rl�5[Ыrm�/e�L�V�gbi�d2���V$z�����˴�{�n��~���,7ҝ�_Ӣ�/�.�:+�"k�^ѯ����7���>�+�_޺�{���`�@�wL>���<M���_�d�[�i\�q�c�"8:�V=�R]n'W�%oc����^bLI�;�s ܢV�?z�}��4Z���._�\�'�б;%�z�ֈ��f7�����L���Ƞ�N9�j����ج�OZᗝ�����N���`�{�ͻ6�E26�����g�n�����V��2�0���{�B���v�"����ק)�͘�7�^��wM�%���o�s�,��>!{]���\�\�%�?n�:��]V�cy2G/�9̥�[M�����ԡMr��ķ�*�㝵�E���g6[�6�ꞈ�<�P�3�<����s�����f��<�]J���9d1Q�N2�׹M������,6�	��������n���x+sȊ�k��c��w��{F	�#�V{�X=Ջ"�UGy]G��s��G�B�gN���+7����D�����3���W��ͻ3*�Cu>g�u����F�]o���0P��%���f��u�§;�zK���<�c�5��|4�֟�SŢ9�Fm��}��ȇ9=�����W/�%���k�&�2�u�u������gk��~��|Wg�&��d���E���E���nm;�z>�KP�a���A�χ�&���,�����t�lͫ�1�e��M��ޏ���/��Uq�f�?��u�
�S��1ۓ �¼&��8�L��[�~w��F���;`�f������\q��� ��;p{�
���㷷'��3cO�iN����Kӆl;y����1W[>��:Sŷ���e�ɼ��9g����w�V��ۯ:�.�(�4)�Ԇ�Ol]�~������U��f�,W\u�~��W�n�!��J�!����}�g[΅�(�j�3Q��z�I���,f�D�"F1[u��]K|XhE����.�VeZ<�[At�Hӷ���Z��Rձ��-��]���"ս��˽���-�˧��³;�-%�Z��}��N�S�Y&�Eûi�f>�v�\�:�:�V8�ы���M�t��I������:z����p�sEe}*?�A�����;��sD�,�r��~5�َf�s7�������S�k��Y]��x��������_ 6�_n�88����C�zs��x�Ӧ��с5�{]���W��<��%����v���UϽ�;�d��}$jx��w�R
�{��{c�h��>�D	���,};��w_�P��g�ÿ=闕nL5�Y>k�tǧv���z|Z�/0���c~� 9��҃בG�l�S7~��r�Zl{ٯo��lx���+�o�x�]�Ll�~9ۗ���HSe�8�G��9�j�[�H��5)wC������
]�y�>�
P4��E�U�
5����?F����^Ӄڝ	ृ��m��=�e�TW�/��7�z�����\@5�[�/:z5]��8'E�7B%r	�2��r�8W-�d4g�;�Dy�ɬ���=݊[�i�oF�K(�,�#3z�)�{5b�8A��[�o��u�r�`�$���[��\`�Z����8���Cז+�w7���A�v���F0�O�Լǯu<�}Mp�RW�5���s՞�[��uu�gK7�s�1v���*�:�K~؇�F�OfeZ�<�+�6n��?m�b��|�^��]sj���ݞ;�i�A�S��W/Z�i�����R�}2˯b��+��H�ɾ�*;�̓B��y�w��<m�_�Y�JҚ��:S�QӬ���ɹ<��^�5ʟS�z����t�ޜ���<�J�u�r����|��]�ng�z�brpި���m���}�} {+��%�{޿�LLF=��P�E*�/c�ޙU+��ٮ)nB�nߝk�'�fs��/�=�<}�WЊ�돩W�j|J~�7x��v3;��㧠�������z��5�_\ST���l�����)�<C�����%����S�����e�����7���x���s�z	�YT'��0��<&��]
܇oP:�ǑU�wR�@�#	��Ĵ3݄U�)i�T2XY��)٧A�g�����ti�Y�R��>Y���%��c� /�=�M�3u�p7Z��K��(���Bz�mAo�6�prF;\�c�^�ҝ��T�@#��r�.-�/v�5�o��lfZ�.���РɎƽܝ�Zӕ� ޴���r��=���=��L����s��s�^�7LC�0�󓈁M�}��$���T~�y[���|����v/'�ov4w��f�>�@�����N;�gԜ��E�wxK����xU�ۍ��b��2 ׷��
̀\��ҽPs�t:���<x���v���9������řn^�L�_��/M�JwL��G/D1���� 4�`vbo��>��Hg�}s*M��@�	C ��g=�Oj��7[���(;]��E�͎5`M������mc��%��u�%{���f�{�uN�(|��Orou<��3*@^�8f��[�s5e���՞pyr��p�'��B���~���N{�Ӛ��e�y��=�����g�3o�֦к,9���O܄��"y/��=�Ny�<��<ݹ*�Y{K��=���{k�Z�G��r'�����g`|5�R�u�N�d�rB��Dgesz{%��JWQ<�sK;�D�΅�\�c���ֵ��|[�U9��h�ڐ�~HE��Z��M5��M���z��Z��ݢh���Fk���S������������rI�麮e?Y��%����Ytzm�v�9��}�>3Uʖ��W��UX�L��3�ʅ�,���3��3�^0���������]���P|��/����Sy��'�y�|��y^_�K���=�:'κ(����ۮ<�2��)����Y@���"^��D�؛5��Ge��l��u�P�є���~Q��ͫ`i�������,�zLq��S��\�-S���R~����&<H�w���^^���vH�^?����$�mz��5t�Q��xO+���Z�ӹ��]fwE�ܫb�̻��_{P��2G
�ni
��lT�F��������f��><4�9W�b�a�� ����c3��Y��k�YIzo7ha��/���q����5&��	�N_��E]aPl�Ll��n�p�R�����bK��=|0gA��>�Uܖ�C�⮶۫�ZGy�VXn�b�#�.�i�(�lI����{Xy� �)
�����݉���tL�f騣��R�:�5��v�az*wm�wm���w]�i�����m���8��S��3s��|3z�^�b����?������u�1{���Kp�m.�Ҿ�b������;3+`;�iT�,-�����{�OC�_��G}m�꿷#]�o;7�پϻ�n�M9��vfۡo����U ���zo��w�@�����gd��3غ��w<���(m�*���=$Sw68ӯd��o�V��ۮ��\}�����ܑ��:`>�H�?Z˚5f�a_b�<�w�9Y���ʿ�������l�2dr]w� �o�ocП{���������ʻo���=�달��߶����ֻޔ�^��u����E'9����x{�˨��W�Y���vn�L�u�pPbiŞ���q�����ݦh��e��$�6�X�jJ���Сڼw�W�i�xzyE/$�K}��m����s=�7��j4i����Z����+He�sUӭ�I��c� �����L���=oQ����a��6kn��J@aqO���ºm+��� ���"7j�Ѷ;$R,���U��׀`G&,��_@S�ǎ�2�r���訩�
��R�R��Nôy>�h��� {Ԇ�ׯ)L��'��۽��r�)�,Pf�e��t̿	�u[��S��)�Q��r]���!s����>>f�uk�ig����R 輪���T�F���[ͣ9��i4��� �]qn�����(\�J1�*��E*��^����Я[��t)���{��z�
���LYO�@�(xr�A���E�c���K��f��s�`��Yums�nOMy>ϟ��v���cL��7�e�0'�]�U�fg;�y8��N��z�����u"�i�
��5:��\��\��4�d͹۷@�]顂^/�y��f�v���k����^|�+��'K������>WG-��g3�w�W�����]ϻ��~��+���e<��VQS�NK|�i8x½н��4��T����|��ʞ~�Ϟo�����<k���A���&bW�G)�q�[ݏ�^����k3c����G�J�CV�+u�(һvx񩪹U���v�!;zv�k��>�����48>T�mr�\K�O^���%�j�,�n�M�]�YxΉb���Y%��h���dz��ݬ�k�]w
��|��]��4�����������9�@�4�,����.�ݨ��1+��4���\�RE�����f�#��<á�]t%�g^Lf`��I��W[o��H�7�+3���]5�؈�ţ8�覃����1�΅Ă�[����xD9>�:̧�wz��%P۩��rշAone�b\��a�y�7S�mhY��i�Yui�'3:ԓn.A�Y���nz�HvՎ��&|��������S+(R��2e.��]l��B@�Zh���[�o���:)�L�:y�K�	�������c�YJu�V���K��iV�7�j
蜂���f�V�hѻ-�h\�ژgV�9��-Y<�kT��3�I솣�!y��r��3�C;1t֔�{�	:�-����쭬��qA��Z���+$B��&<88'6t�CG����V�;u�irk.]�AF�D/q魬Ґ��js[@8�)��g��r�����w!I�6ZH���hMt�[�[M@#�jW;S�]��S�����,���-JҚw�+,n	�c�.B�ь8tK�+��a�WY'�;�N�\/�J��Jn:�a�&�D+�K]���-�0mn�{ϧ�Q�]�h�/�us�-�f�[Ks:����N�y[M!�+=M�J���W��W+�d�`���z�xea�9]�/NQևP�,\�9r�*Q�^F6�Pcv�7&�p�몜��]}���R�:N��EC5�ZŴ� k!��[�n� <5�]:)j/O��R�d훼�d�(#N��RQ�t��R��1�,R�2�a�g{9TrG�!��Z�(Q��w�Y�00r� ���-xN&/���I���C#>�wR�xFV�.��N���ջ@V���g(PxD΅2��ʚw��WB=�G�%�4R͹yt���2�1M]�b�]��%4L��;�n���m����m�!{�*��ڰަ���Q�V1�-�.i��֧8	+����ջ�b��1�
=z��U�\M	�X�/qǲ��k) �G᪣���f�z�`J�l.u8n���U�С,�M��iȈ]S;�^��O�[<��8\��Q��e%e�<���B�Lt"T^�2r����9v�v��>�M��>&���\7Y����h�,��B�,�v��(�-PvS
��v���{B�mD ����d���!ޕY�^$��i�4-ӥg+2�b&��T�r�#�O&m�����z�v��É�u�n��h��ɐF�e��A�䮠�c�%>�t�RMc;�]�o�ʋX(��x���Ԋ�0эQP+[j
���Z
���!l[Qb��[l+Z�P�T�ZUX�R�VEQ-,B�kUdEIQ�2T�(���e*�lm�5���(�*�VR�R�(,m���iQQV
%�Kj��,ֈ��D���k`�"����b1PְFР��Ԩ�G�b��S�c��b�-R�DA[lF""��QjTT*�Zj*#dUUE"��PD�(���#��c")ZۜQW���b*
(�Ycieee�(���ň�5���E�jQ��**���ш1E�[J�%�*Ȩ��c��iTUU-�+mAke���R�qi-+���"$b��-�qE�Rҫ-�����-�1E�Z(�+V��QQk���P�J�Vֈ�8I��cmQ���R�e�Kj�0U�QTUUDUEAp,��QVZQB�B�U��\\`�9j&)*U�UFV�3�0֭��m)Z�*�[cZ*V��,�"����X�(VQ�b"*�DY���`B�Z�l�+**��QE���
"T��X���U��PQDV,�*1Ъ"�JR�ԬYm�T���k�Qh�խb1V1�E!X(���1��J�yCA�o�6LC�`�O#����kTv��f@��e_S�	�7�֫�#��i�E��5��O]�S7y2���14E|���"�^Yie�"�>����4���5��*o�kdn.!������]�w��=�6�E�딌_q�e�Rߥ�3ݳ����ʱ���S�Y��B���þ��]S��2�~��4�W%!xv��=��_z�{Cr[L>ս����|"���=ByF5imx����e��+$s���pxwǻ�'�_'eA�+�����|�2¾�WT���������sJaRｽL//m�:�����-�9z!+��$.�vfg�������[��]6I�X����I�؍}|5��n��ń���f�srv�����O�J��#������t�N�	uY|4�1��V�w��{�u��{Mz��)�Κ��U:1q�{�hXҖ�-G�~��i�EⓍ�\ͣ1��陂�p�$��#4�/o�֠�o���O���(�6�;w�b�+ڝ_��l���}Β^ZE�p�s�7�Ѫ��U�[�w�H��=���Z+����َ�-W��n F�i� tZ{q �w�%�v��ɢ@m��b�����,įf�F��g��� �'��0e��c�9��w���>��^:��V��W�=}c�Kme*�Q��3��.M�ϗPێ�y����c۪�Գ[�s�C2X�ٻ=0�i�fG��&��ݻ�Ra������ϖ�����Ǧq��k�N�u*-�3�6'��t�H�<��;d�����	t���7>/=�$�O�o��R�Uka}����;/f�o�=ۓ)���߽N��M����(�ʲ⫕ʭ����k{6���tʦ{�>�au�)��w��ܵ>U"���xǵ��W����ﲩ�E� �a�	��
줖?sW�=�q�����'��R��mP�Y^�g�V���\I���y�����Y�>�j�dt��s]g�b�v}�BOx�=�c�cU�����͘��C�qnK1��vF����CD���>�|4�uۇ�)9q4N�λ�@/km1��}��N&�0�7�ٗ@	2b�sE�rZ�S��k�fP�������V�������Eޢ�L�ݶ��Ŧ{�J�6D��Ww��eD��YzZ͗2`����/�D.�P�ٳ��)��ݚ��-�{�����Mq�N�����Uΐ��S�4[%&�2�c\����[O�����cҗT��{lk�����I����]�o6��� }V�t)��U���>7�<��b.�`�Ĳ��]x��ݗ��{�Oz��.M�n�I�Z���3��u���]��eԚ�c0M��vS6�]^:28���i�r�I���ў&���0|3x��}{q��Jn�m[���3��A^׫�ұJ�R��M.vfU�zCl�}8f��nk������o��,M�������r�oxd޵;W/'�w7��<��J�2b����^b��N�����ϔW'Y�y%f�	I亜��������%���X��ɗ�ә�/"�yb���s��t7��R�������Q~w�c�X�j�)��7s�7j���<��П�� i�5�
I�L�sv�&�Y8��`}�2��~���<���3���.��K�(q"i�p�pUڧV>�.��\��2�<��&qBMb�b�j�{��MY�%���A�#(��޴���M�����G�MG7��"}]6f�Z�CoZ��N��7l^�p����Qn;�E�9�s��NR����K
k�����~�w�Ʒ�1���О06��q=N2d��C�q�d=;z�q��u�C�����p,�g����Y4��Xy�Ci=dλ��6���`�jI����^7_^룬d�gz�t�����&�l�8��L�f�=�
�u9�m�Iԛ;��>d�8�[	�
��ef�N��Qd�'�ͤ�'���(@��|�w�?g���������睒x���4��m0ɴ�z����8��m�� VC������d��@�l�C,�C���!>eI�劲N!����m&Ͼɭ��{�`��o�����y�/t��O-%�P<d�1�N�3��'N'�l�!�>`hǸ�d:���{9C���9�3�x� xk��hi��G;��IP|Ź~�t�q�{���u�7��9RL!Ӿ���I3��hd���`x�+�I�}��x�q�3I�<g�LY��Ms8!�I�s�OY����i��Ư{�5O�sq�w��~;�1{�z���w����2c|���8�Ö)>k	�^ |�	�L$�'�~��r���C�z�q�����XMf��z¦~���?cW.����~������&��e��X�0N��&f���a�s�$�w���N�i+�'���Cl�3�p��O;����L�Ng'o=6��y��7g�=�<����&ӽ�ROXT�,:����1��Q`jw�
��&-��u����09��d��"�I�	�`|���&m��g�ߛ�~����ƺ�;���w�c����X<a�OĞ��0��\���N�7a�d�Ow�d:���<垠xɋC=� VJɎ��$�&�+'̇�Z�\�~]���m��{ݽ��6偆a4á���C�&����q�I�'��I�]��N'7�wVI�js��R|�C���i�������>�#ꓦ����_�9]�fD̬��u����6�W1H�qsk/A�Fj�#&%�p�p�n�q�ڲ����^'���8�3��*d���\�8�4�c�3��}�[K�\���^�#-U��Jiqcs�� ]��Y`���T����+�RN��'��W�����w��x�&��u�Bu�&Y�OugY'�>�8�����0��,�{�=IԝE�Bi����j�0>�?W�� �W��_���un�s���W�}�.�ӌ$�6��!Y��~��+������L�=3Bz�Y5�I<a�ĜVI�=�:��Y5�'�8��y�O:ϵ�w�����{��q����c��XM�����Xz�d;�=`z������!P�b)4��8��'��f�z�Y35�dY'�4v��RL�U�}��������P�Z.��_2�	�2nӹ﹐���ş=I=C����OY��s!�3,9�1'�&�},��C���d�4�d�O�E@}��+�ΆK���ߊ����IK}�6�dղM�퓉;l|��N'��bCl3S����</1!�m���ROY��m�|�ŋ'��!�Y�_`��(�W`���xO�k+��&�������Qa8��g����6��x���`q&����bC���{��Bu�C�m�2e�}���+�+�c�|�Ժw�4~���w�(��E�$��XT�=d�g2M�kě��״6��u��hq��=f�����d:�����d��0N��&��>-��3�u����=$��O}���=C3��Y6�!�x��M�{l�<d�[�a8��;�i�I��ֱ&�x�0<N0:��m5ϰB��ν~��r�G�Kc~�{���_1U������L�g��VLy�
,��d<����g������<���Xi4]����OP�C�CL���|���3����zxs~o��I=gӽ�xβM����>f�3���&g��$8�P�{�E��L�8b֒gY�>a��O3d�Ԛu{�N$/}7�g'��Mvr&i���'s��� ҺΚO)�<�m�i��t�_�&���
�r���4���q�yW%��QF�a٩,�݄�%.�{��u:�:tX��ol�*x�S����]�vP��(\),�ٚ��~Ӝ�o�o{�er�z�C�O���d�<3�6�*�7C�u$�{��L��CɞbI�&g3��CӖ8�N0��`Y>���� m�OR_��w߻���Ǹ�<�����|ɤ�fО25�g�4èy=�u������|�ff��,����C�����,:��L[��:�P��ń�"s����p���^wI�k8�~ί�;��*M�I7�� q�ORa�!�g����SL:�Hq�����:���	Y*bs{�uISG)���w�*�a�<�^W�{u�z�n~/��� G�f�~a�\��/�N��`|����:�Vy����8�x'�0��u&��|�,�GvH��{�pE��k]�}n����[���w�g��'��w��(0��s��Y+&�5��&��bVzϐ�J��|`zg�N2OPיĝC�M��d�zɤ�d�&^��\����|��g�{�s�z�����O�8��o�&�9�C���CÔ�!�(h����*<���y;�zϒxé�C��|y�'Y'�h�8�����×/�t�߽w����y�vD"Y���U1@i'>��9�N u5>�!�XOXxw��z�	ϩ��L����O�
����
�19�l6��4�&hOR�����V5���=/��~��Sr��)&O/�6��`j{I�08��y�� u5��m:�|û�Ě~Bo��r��Y<d�9�ɦm��>�����>׼��u���|za�OY�t�!ԙdλ�d�$η�qo��d�<�����2�|��rc���a����8�!<��̇�|�!�cxþ�>�}���8�}��qȳL�Iَ����5��:�L��
��O=�����d�M�=Ĝd�2yC�0�:��$8��4�6�!:�����w�s\�V"�V`��<�to�Mi��L�*ݠ��ޡ#�izzQ.��#:ǲ�È�	Zw��б��}}y��9���j���*xI`������9��S8)�,�Nǭ;!]L�(���7@;�¸��=��p�����j�N�1�9�~Chi�$������0���dY�I��Y6��'|ɵI�,��&��2M�h9dݰ�fg��I����`m��i{�������|�o���~vY߯�'Rk�ĝa�L!��I>B�ﴬ���ŊO�B}l�O�<�Eh$�kx�I�UG���W����e?ׅ~�v��Iy{�wx����!�=gS��+	�y�^�<f�;�'e����:�3�p(�N3'}�b�h�4[�?}�}�� ����"#�zW���n��y�|���xI�{���	�x�g����Y�Rx�S�o��d�9�܆�>CHv��2Ʌg{Bu
�����q&O;�d��N�����=�����~��M�yl����=a��y�N�3����:��l�C�|��xf�a>a��s8���I���CL�"��,:��L"��	ĕ���O}����h�ϼ�����N���x����K�����x���'sd��M�Hm���p�$���Xu&Y���z�L}�C��	�W^K�b��@W���:�_�%V�LIy��w�s��	>dš߬��*1�l��5�`Xx�a;�@�J�ə�06�ɯp��PY�L��5倦L����*y�ͽ�r��5�y�ƍ��[�����^�h�O����z�C���xɋa�y�@�fc���'Y�I���ذ>g���Y�!�C�e��ɦq��򞡖N���/;�sw8Ʊ���>1�7�����Xz��zk�$Ru�C���g��1:���w�
��&-�y�d
��q�+	�GtP�<Bq6�6��&<��	��Ͼ��O�k�~�<Ǘ}��y��i����<C,�E��$�&��o�N����l��9�C��[!�S��<rû�+%I����0�a��w�=g�N�w���w>ſ���0瑱I�n����x� �k�4�U�Hf��C%�2�z, )_Z�@��A�í*U횾�*�~ƶ�-����ݏfs���kv	�nk"J�yE��3we�.e��h��do*�V]�����~+�)6����S����n:x��Oݧ:�{�_����פ.�>����0��;�Y'�c��O���J���ny@�';i�v��O~�C��&�{a�'̇9N0=I�,%w���>��U0=]���?oO�,��J��k�~�u�E	P;�N3l�g�y�!��fk��a6��Y8�I��:��(=������y�O:�;�M�I>em~j�
�C}W�S5�ϤA�O7-,�۸鴇�e�N�|�T=u��Y<g�s8���'�i�L�Xe�\�$�&{d�,'���$�'m���0������AC���NB<�������Ϛ_� q�����?d:β=d<C��6w�0�3[��L�!���d�b��OY3�`RO�k�N�$�����N[w�Ǟ�2띾��Ly�|�����I��߻��`u4c����y�`�M�l���:�q��u�C�����b��!��Y4��XT��x���3ޗUY�չ�~_�ś��O�v�W���z_�rɶ'X�8�:�Ǭ���u1����Bu'�� ��2a�O>�s	��gN���ɴP�[8�����w��*�i���^�4�{��y߻���a&X7�I:��w�ԓ��l�$����ԇ�6�9�@��S'}��6��4���:�Y0�^M��aPϼ_ �}�T�Բ�WGe�)���z������z��Y8���>@���H�m�L���Cf>�4�a8�f�i<g�b�2C�|�NsYXe��9������W�B���	�޿.
>���y������%C���1E$�n�'֒s�dݲ{i:��&�c�'0�z�q��i:����Y��O�����~��e�*�5(��]z�3;�W_�.i�[�8ɤ�E�3���=�6I��sI�XL��8��OY<3I��4��N2����a��%!����+��]o�<ں���x�� y�ڡ�]��XR��< ֈޕ��8�e~;���V�|q��;�]��p�b��>z���;�6%mҾ �y���m�� &�7��6��Ȋ9>��ڀd�M��&��q��w7,z9�T����j;���z��:f�}��UG|ǜ��s�_�2OT��q�l'S��s��'Ȱ<9IԞ��,ɞ`�P+����6�Gz`�N��@�J�ɜ�q!�a���8�k�^��=����n�۾���m��T�Uh��}�0=C�O��'�*zo8�U�q5�`:��,C��TY1hg�ćY+��6��.�OXNxc>C�z��c��9nq�7�w��2a�7��d4{Om�L�O>����I�O9�C��8�/0d�М�q*���>9`x��1�c֤�d����~�,��?z�����Q�S�D}PW���XC�zɬ�m��u�Hq	�i2u�I��bO�4���$�$�y���0�'9����h�1*�<L� y�0��:`�燜�]K��U���aӾ��0���p(zϐ�k	�i��|��$����$�:���&8�'Ǵu'Qtn������Ւa��w]~z�h	������_�G��
�����x�󸀲a'�Ϩ�<``9�
��O�a	�a���ROVN+$ϔ�d�,���m�������,�G?%?MO}�}��}���~f�縆�z�2�����a�{�>d*�x�M0����6�l�3Ha��2g�Y'�>�q'I1s�^��>�Ǚ��|�}���7l�hd妦y�0:�cx�=I=Cý�8���!���̇�|̰�bOXO�Rs���O�!�,6�Y=g�y�l�Iû�-g?������^����?P}��}>�I�ѓ�9l$�'Y4�Ou�Hq��k�3�N���q�l�{x�x��kβO�F�m��3��X����3��\�����M�z���:�ԙ����u�I�d�u퓬<x�״8��M=N�d8��s���'Y<;�I�m�,��7�m
�y����q����it����8��N��`�D��+-�w����@U�[P{��m��X��n[��Hҡ�`�u������:9ԅ^I��^��.�J�y��<��½O����н��Nn��,��q�^ټ7�m-0@���$$1�6h޳���3��CI&��ʄ��1:�l�����zɝw9�m�F9�7l'}�m���'CL�8s���S3���6��d|��\�������ޖ����}�����>���&��!Xy�(�N��y�d�,��I�O-�д$���o9��X�	�i'��6�I�G��!�=f��w����q���<ξ�~�s����0�O��]ěCL�f���N�T3�p(�N!�9�d��L���m'�I��@��F�'��&��:���k���q��\���7��M��q�'�'��<�3��'=�M$=f�<�1��&f���C��v�,'Rbk�Om$γ� m�Y0���2�<������_}���s�|c��Hvw���Bm{d���OY'�Vo:�RN���4��<��!ԟ2ajg�!ԕ&q�G6I��0,�[	��y����ƶ������>�9�=���`q�M$�l�0<Cɬ�!6�h�3�a�<��Xu�)���$�
̛��E�W\��'��3�bI�&-��<��T1�{�n��i�x���܋��_W����B��˩>��*z���m��fu�q��yM'XC�<=�0�����T��uI���O-��9�����w�0��<1�5߾�1Ш$�P�>��V��&�=.�)2���V�i�2zfÉ%f3�I�q��i�d�:��2z�G&�$Ru=�Mkg��y�~�q��E�8�_������8g��W��?����L=�q�;q:�m]ƈ��j��t��o2�W>�מe���H�=B.�*p͹��w.|<�3ѓY�Oyfx_X}��Ns3���#(G�c]ڗ/I�K�b7���i��
���j����@�S��'�W��2���\�*w���h��+f�
�һ��rn<ȩ��xƼ�g!F�׊��*�զD2S��gK����D�v�4��2�b��m�*Raᗫ#�6�5�$�%{�y�w��p*"�5IeiX�F�9�e�E\�xq�ngv��ԧ[���d� �vO{f��ص�6��#;$��z����к�ٺ�<<{�b�w�TZ;Q�&p���_؛ǯ;u��}���%Ô�09�5>�C��-��(:�i��Gw�ۚ�ڏr����ʝ|2l{�9�zr���"���U/6.#��X�g*�M/1Kv��[�S%Le9�s��Y%v�ᥠQ�]+)�\r�-h3�!�DF�Q�љle�;��,\��1gzl�td���s{m5Z�9�݇���8���ѭN!�X���u,	��Z� �hk�VZ.� �)��NdjX��XA�%c�ɛ'p�Z��[�2Ј[=�����[ʵ!*�k¾m�b����U�c���Y,s��m�#��\������8�pm�=Lk꤃���n��J�i���mdW��w,& ���ɶi�Y��Q\ 	�&T�w�`�	]n���o�����"�P/�ѱ�3gRt�Ct�V���X)Wfe�w¬�+�D�9̊WY0-�M��r�z�]�0������J��o��W�}9r����z�6���*;+D�ެ�3&�}� u0&�;A��T��|.��h�l�*���M �\�3�Pm��K%w������K�;%γ��b
���Y���r���92�P
P��+RK�:~w�X@è�2��
���%,z��E�#����,�M\����]����������IV�t܎��7u
��i
b'3hPۗa9)d�oi.ʥ�1��t�Ǐt�O�L�6���Y]�eBN۽��A����ף �H9��^TR���r��j�+�or�:�8w� �O�S��c��Yk���c� ō�ot�:-����:�����[4�4IJ����^��]Z�S��B�W@�b���C���&�:Z6V7�����R���Ò!6§Qt�-z�ó尛�;Wp+wWqŜ�T�� ��ļ'��u�ڧ֞�)�F�# In��E`���� �A�y��k;��6m뿚�
�s�+~)ŖL��d࢓�du�V)	�2�Y�^�wD�`ξp���s��ryr�p��I1�&ʖ�fAb��C�ٶ��Oj����p�;�a��).�c6,���-��{7*��&��&s�����y��:l�P�$������^��2�[�ЉBW(��:�7K��q����dEPQ�X��1�����"�VڑTQ`[,���+b���U�ZDbIPQ��b�Y��*T+R(��Q*��QQR�E
�k4[H�b��*L0�Ab°�m�!iEDPDQKJ1����e@b

��DDB�R�����
�m�6�
�PPX��JAAAEU"�+"�(ň���++B"V6�mAE�d�,`��J��Ki(���,R",V[0��U("���U��U�U��*��P*���1"����ԶJ�"�1EX�DPU�B.�&Z�"ŘB(VAH(��E�R6Qm*�DV2*���PU��*��,�%TDV(ZX��G	#J*�X��6�U��R�j"*�E3lR*�A���,���(������QUŁqaE"�����*"���"0Q��AAE"�Q�`T�T#ڭ���d��m!DX*��E"�b���� �L�qRЫkJֵ� �
�*�-���X�h
,P�b�R*�b�
6�F6�Q4���08�TX�Ŋ�4V ��E�R���TUT��Ub��X���VJ�]�ϳ����>������zx��&p���l�����2�gVK<��^;�L�L��[��:�8K̼��V�Z�����|�x:�Z�I�Y���ί7[�-r�}=��Nwv��ኦ���޷�E;+�5�
����M��A:K=[Y���b�<��oNy��uw�7c�/�vp:s�ЊŞӎ<��U+'��W;�Q*��뒻���K~�|������5��Rб����v��1��M�\�Bfз]nU����2G==�>�X�v�zQ��D��3;�z6n���j��W�YG�U��T_l��en����9d���<�{�A2{�|f��a�7O��ǃ���v*z�&�J����/�^DT�Kс�y����7���2�v^P�U��|4TS�CYX�6����{e�_C���o|����z���^����/ז��Y 9>�m��vz�F�<��d�:�p�;��%=9��m���Ksʔ��5����bV������9)���\3S˭����{Q/�hU�$�#�ė�+V>�l�܎� �v�8,Vd�i__�W�Sʋǖ�AD��^�L�$��d[
��-�ͩ��eя�.�I������]��k�i��Y5]ӫ��̺6�70������1�LP	��d�i���ݼ���԰��y��7���ꯩrߖ+��Z���wv���8tZ��=2�!��먹�,)E�<��h��9K�״���9u��h䐞�0
޿��1]��-������6e/3�1e_��/���J��#F�I�z�_Q��'3��Kʸc�g�5<]��5�W��參�.���^נ��r8뵷z�h�ޏE7�Fj��o�[����p_����f��i��m`��a�y˽>���n�,���׉�ŲW��>��l=G��Eײ����5ߥ=�N1��՛qu���R��yU�]����YIN玹\�!��y�8��\o���&V������v*�1]gS���#`1Ա��n�N��!����:PR�,/{�ޒ$&�ޡ�1�P��V�o9�{�鳹�?|d>׎����I�ln�ѡ�s�E]S����B�����~�	G.����!u���J���l���0WWsU(;�k�fW@A�S1�.�>�_q�\凊�����V�,��n<�O���1���i�S"�r�&�@�wL�tp��WU�wN����*b8V7�丵�U�e���~_����|՛딼�{g������XwN��.������e�=خIg�����wrɵ������L4ǾU�c�3׼\�;]�2��83~*�'����^�r�ӯnw�u`�i���������٪;9c��s]�?/ɳ��Ig�{�۟H�$�RRwC%xY|p�*������gd��8�=ܞ�K�Ъ��eB��9�E��]'ug�_���9��)��ށ[�۵������N}ꃘ�;��tt+�£:�^gO��ّ�F���=˱z��T�9�㹕^��WT})�sDbȌ �aC��u�C��R���_N�I����(�6��V��b�=�U��Oa���X�G"�'e��6I�v���t�b��wF�8���p��r���qo�+0��z�m�ގ�Fl��7mz�P���m���M�9+
�Tpb��hi]h�QWXi,A����p�fl���|���z���9��K�V�ʏ(��EW[uI�k�y���E�zw�]�=�[Z�S��n�^f��XK�C���ʗ'���:_*�Y�4�IZ���c��vz�]��nhÍ��{�c��T�O���تs�u�� � ��Qo�{�˭?�.1���sg.J����ե�dŵj�t/0k'��.�q,W��ar���g0���.�8;�$����R�o����׷��}w7GhD&Z��O{b��A����j�cʷ�轒	?�¥׷��f���f�^{�jOj�u(��>�O�k�ߧO�R�����y8	�m3:^y_+��-�M�T�����WY|�d�o{�uv�ŷԋ�n��N~6xZ{�w�������՟x������|��r�<�-S�)�L����+��{s~�z�b}��ׂ�v�n�<�R��suk7 7���ͱ��K�.��m��S�vF����	S��4�V��^��,t�5q���`w��6_��ٟ)�zL�z�KCt4���`��g�-����:Zv}����O:��:�Z6i����f����(kg�B���f����.�%�`��c{N_o��i��6�N��D�N�9�f�Xdk!(��x�0u�	�Ɩ�]�|�W* h[�#��o�cV�}v�.-Y��o/��ACiؙ��]}FR$�7���0�A�Ұ�3��EfBԈ�e�zW��{ު�2�������x:]tȽ�>c+_�\�by��Lu��q�l�O�~��PM�=]��y	U�-�`W�G��]Icr�U��V����Jt�۱�+zQ�0lc1\�#����O�f���Y��s���S٦����S�j�[�Ҷ��z��/1��۵������}�W��w64r�,V�N�zx�H��ٯ�m��I�/s���ǻ�V�rx�N�v_�%`ă�"���.����{nR侲�����lZǳ'Lbo^�f�)����8f�����Yw�л�+�j����˒��ו�]z�[�>a�̰\7��P�S��&����]��r�S����������ڪ��+N�l��+��I/FR#�u�;�_���Gx�C�{+�+�T��Њ�X�&#�[���lM��H�;�n8,>S;������C<fx�/�å�]K���'�`�� Ou 㬳���U��-�V�jQ᭡ [�X`��4�]�9\�ܺ�u+�o6g�)�PR�wz������.O)�gv]�aus�\B������{� 9�r蘔��U�e��e'�E��{4�NIq4g.S�)R����vn~�����q�g�w���x�N��9�u��G��'�1ӧV��}�w��~��m���v�O�U~��g�����M�nU�f�������;K��U�nemoF����G�^�8��u|��?�L�Y�{��#������Ѹ�q��ƺ�?��y��Ϭ�����]�D�f�ԂZ��%�{��]�����B���G�8t�u~��:�O��k*&Z;\Qt�gX���oMoI _v��`�8�3���ҟ�o0���E;�m�lV�x��&��ԝ��J�������ށwK98�5��(N�.�V��$�>�9m�m���ْ���.��$��g:Y��pǹ�pRS)E�Rn��5����o��z	���ۘ�Ԙ��V�x\��S��/'iY=�p��pCz��r[�w��@�Osm^{���_՛%o��Ù\���5�������QP4��uK�aM�:���{sʺq�v�YQKad��WOu�B�%�k�����{�2x���؊Åq�����&:x��m���g���H�,����2��TP�+�KgVX�zN�����j��gXf1<���/�W�U_R<-`�w!���^~���;������S_�Z�6��?uk��ʇz�v�`j��o���KZ:�t_��m�TٻW,f��Ҽ�X^�|4/L�xVqFJ+-��,z}
�̙�]�g̾�#.{*vQ���)}����byo=�1HxK�r׎�_\��2���ú^�R�;�TW8fy.��%�nl����3*�mu�|���/[��|"���5�X���6�7;d����*����}�:�؞�e`�M�;��aUvkg�M�����\�v����!��y���O`�n��,}��ڠ��GVd�p7}�O�??�s�o�A�]Ƥ��B�㸞�FY�ͯH.|��A�:����)����
����8I���9���!Q�����byܷ�ޙ���}�=o6����R��6�F�p/����
�p�|�Su�o�8*�	�k����.u�No�PpU���"�Xz�b묈)Y\���
U�.Dhb{�E]�k$���/���a��_�l3]�]��"{q�\��ZA�1��0O�ׯ���l�Iu}j�lz�şs�s(�5�͆Z��].b�s��<|���eg�lI^:�k8����6:�Q��4��ޒ�.�h����������M8��8�>�^m�-��\͊z��]gT�r���	�ȼӬR��~��C+S���h����F���K���=u%��P1��_�W�6��o�jO<J�=�)�=�1Е:ʡ8f�N�e�;nM<6�A�|���X���b߶N>{��㽕Ȧ���m���fͿz�E�nQ��X�n�y�Ώ×T���O%�Q�ܞ��ٙ�{�-�{j�V���gq�[���ZvG<����J�:��p���-�nL�^{��y޷�7f�k/՜�)�.5w��tлn(�W�1��[��Ɵ0�9A��&Y:Y��ױ���f"��7@�U7�*�u˝�غ�~}�oϳSy#��=��=wm<��R���o�9�>m1*w������{XKۨy���%�{�y³:;/�_��sǛ�=+��f�3��<���յ���U�w��{R:��ub�����$�#w���l��b򂝢�
=|�SWJ����(٘�q�f�����3L��KT�W�"}uݪ��b���f�ѹ]N,r�؝�[�8���۝2�0�����W�^�,ܭ��~s�;��u�ܴ�#��������N	S�7��ulnS�tm��6�f6�I냆v�5��� ��:�oV:�u.���ӫ����l¬g�l�r�sܱzT�=��r1�6�Ӿ���<i'��h�1�����_��W[�L�����j�����[}qo�4�ި;��8�6����V��E~�"� �� �z����B�Z�.[��1U8��nT���V�X�ڦ���ƣ^�v�p���/�Q�6��I�ϻ������,��{}O�g��U��[������ԟ��_^���8; apY��:���^ɉ��7W���ͽ���OPX�M{�=�l�,n���s҆�;yyA�_�B��<�����V�{6�6�������M���kz[�z�������x�*������T�I�7���n��I<c�Rf��ůwI��С��"@[6U?��v�����|� ⧦�-���e[��k�����Mus�&h��.����%�2kЬ��5��**�B>9�J��TB�ox�լ_
r遮��up��mN��܄9���+���1w�{�C�U{ު��d��d��s��)]Wt��㙿.K�u�nJ�l͘�����r�YW}��_,���M����mvנ�ڽs	�:��xE�2�G�f��2���6�z9uFs�>��6̡=�u
��`>�r�B,!��]V�-Z��.ń=��k�����3L��J_q}��ۦ�rI�ߥ��?>���(�(�����/6e�H��}R�>�ԟ�=�W��Q:�����\����F�1~>�^��fY��b�~������*#6} ���w:a��t��x����>g
S�1ab(%Vr>0xVx�kDn�!R�C0e*�;�h��4������c�=4,8��%
"1|Δ%���`5�,��#fk�Ɛ)��y_J<ynv�;гXd]��7�k�.��B)�T�0��*Ǆ������j.�.�v�ܩ�.\���2a�
���}�@�X��bCZi:�
5�r�U�ڣOJ��^�o+B����0�|��k��̴x<�˃�ЖWA���[��n[������	���ۇU���8�y�q;��m�('���7�-)��qNNR��y5�Еh�>O�A�v�ե�	��U���,�P��0�Ĭ��q1>zsZJ�G���\V9�0RVc��|f���b�j���{L�n;89���+�p����k�^�wK2S��C3���f�駉����/2b������s"Ih�y-��9��6eaDa\"������O��W�2{$eT4���e���&�+�X_!G$�E�o0.�� ��*6�čV��w�r��Mm���ym�
��7ë2��r��'f�&��;X�����նk��k�ts�8�v��lk�%�k^vԆ�U�ryM�}���`bT[�u�u�Ru�t�+��(��m�㋭�h�²���k��23o���2��
�>܌
��!�?3G9`�/FNdW?�b�`�$񫮾yjfct�ۉ�NP��Z���WK��}�;Kxܠg�[,o	b�����&���/-5au��ś�6]d)�}��7},�խ�˘��
 ���CO����U�ח��+��/Qٕ���n�����]\v~�G��;z�f%}%�դIc��Zv�",����`o&�Nt��؛q�[��[{8fhyӀ�O1Wt��N�}:��O�A�2�z�xhr]ec��f�m	�Om���0�\2ǡ�<m�Pչ쬦
�S�dQ*X:����sQCu���2�e�9:۬��ƆkM�*yF�c�[[�����V�G�}S�)�)��bg0s$%����&�г�=�2���Y�Vͭ������y�l�;%��6�����'1���U(=��6�-� cz�cRӓ+jA!c�����t��.@���Eƹ��e�5w6�\�l5�J*���Z�4�	.�#f,��vZ�{z���)���и�KI���;	[/��*(4]:7�y���a����xS�"8���J%f,���]��%�وw4D�ޫ��i���Y\%�{i�!�ˍ���i}��[��ӦbܓB �{Fr�
��=*;�G6���tyl��HʺÃ��P�r�S&��PV�B��P2���Ә��S�$��������;#U޲��8J��7%�GY1�1�eԡ�J�Ƚ̳���WJ���.(�R;�lQ�&P��.AC u�u�T�-����i]�.�!0��1�EmJ��;*�AXooT]x�b��2���4A��u::ǡ�]�_���r�4�iJ�q�a�(�#�դ�I	~=ڍ];��gE��C��7xzP�a=2�Xh��;��E%����2��o�ɰ�T��C}j�����B�p��ۚe�Ts���.����T�b�����J0�V�
�£R���B�m���V����e�"�ER����TUU)hP��,A��V��Q�5��`�Bڢ�VT+X-�b �b�҈*��h�)1��"���J�G#*�JZQb�1+ie`�ʕ��m�������mV5�Kp�V8J�Y[*YF�$YikQT�#""��"�"ԬD��YR6��4�(��PZ%J��%��mAZ�6�im�EP����5�Z" ��@���T��TF�D��Z�)#���X��ki��V2�U��\Akkj��±EQ4�*�`�c0P�
Klm�Q(�ŗ(�	EAT�(���hQ��V%lQU���T��U�b�X#�ŕ��F�Pb��-)mm�(ŉ*��F[%U�
# (�X5���-cZ�YUE��ZQb�͕Qb��YR�-V�УPUTE
�*��H(��(��A�)i+iX���YR�jF*�`��(��#����c�
�e(9�0Ũ�b��I��#�9a�CSB׫u�P�����r ���������â<"�j5V�.�,�<���]$F)��ov���;�?��UW����L��h�};m��m��:��l�^r�,�y8�}�F���n{���F���O�wF@���7޳�^��0��Va�è�Y͐����ݱ=^�So�^�8�:��������'6�Q�3�c/�FD�m3�eV���:�E���<�����'�U�;�$���`� Gy�jҫÚ|+�'C�P�,q���q~�bܱ�nz��,���Cᓝ��[�������Ϝ�-���:�P��K��X2���ne����)��?s"Pp_\�M�������Ձ=�ux�5�c�g���7'_��VV)8{&�.���x��/v��"F�ԅ1���Y�C�b�vC�uWwV�C����ڻ5^S͝LS��t��:�$ǆ4��(�/<��]jd�F15���*������ur��lLm��g�d���M�~�S��2�E��ݱ��f�,V����&��N�¬��h���Hv�#��x�7�bE����V�U����^�����(��T�U3)�{F^��nJ��qE�G\�E�m!�����ɶ��<=5d�d��&o��L5ln���m^�.Ӧ7�����.R��ћ������A��?�n��X�_#&Y��
*�\tJ�k���tl���Kjv��N��S��e�}��,�T�18n�d[g�fPI9��e[�3^�ߪ�����n<���>��o�z��q��Ć®��X��ֺ@R�`�	�r�S׶�o��f'�$w��ExH��M�߰����T�������XL\��f�[;��f�S9she�o�u���+�f�r�q�I�:�K��r��Gg�
�X<�=~��4/(�!fn{��Ez�b�~:M!�� 7[��.R��VP����E	,�y=�T�g��P=<�崜�2�x�`�>��*�׌����:�g���5 �L;\+_u^���S���)g܃��F�YT����n�>�J��[mY�S_R���6��%|�U�]OYWM����F�i�������C��01����3o�����u��\"e�-Q���`i�g���>�k�+σ�-�p��`�����[�٬���(x���X�V"�tet��iѷ�鏶�U�1rᙂ�3c�<U�ޡ����|�GI�����@���i������ߗO;��Z��J"5��>&�9H�KޒZ}��Xe�ӽ$s2���1oO��,#�_��9Q �F�Wc�`	uunb����{��iW�E�Q��.�\��������IQf�5�n1��w�W�^�P���Ju罰U��Z�n��é�Z�<�K�(!7��j�pv��h4�`���{vޢ���V����1S�*���c���Zp/_W%���Y�ld�bp���1��2zD��xF��jo*䙀��͟���l�9_5Ƹ�<�B�g��V�V����] ͹]һP�>r��{�ߢ��F���/_z���a.8ש>^��&��އB��-����z��l�7�v"*dbڿ���U���E��}P��
�L_��S������E��I�B���<<6b�G��g�:�i���|ʧ��L��O��r��wj���9�*�'��f=Z%
�X�k�r���\6du��(B�QV�"��3�)�B�w��NU�T��)�����|�T��'Sf������X
��C���Y0Vj�*�ض��3�z��K�r��]MץiFj�'M�|�����N��@&zq��϶���;k��9�xA�@|b�i`�kM)B�.ƌ6�z{>��|�Ep�W�Wt|��}�y�X����f�wF�H�:n�f�_���C��*���ם�S�#���ujЎ�I��)���`U�(v�L@ZF@7��
%�+;�/Lq<7���Mc5�����{�*�W70&��:���hr�ŝ[��g�������W������4�����՛�A�J848t���ѷ�= �* ��Oa�*����*Ì7�},�s]y�}r�bw�KM���y����X��Z�mf�H���
�]��
�����#�3�	u��_�e'~�tx ��G��ڪ9��+�mC�t���V�q�SL��<���7Aʮ�H^��u���+f;��C���xq̛��7�;޺��.����]_y㗉���६�P�!��vGԳ�������rO��C��ϝ��l���h;�������/��rI2�ҷS�08}b����5��+�E><_��({}+�v�\����U�����&x��)A�O�A�D����7�,�b"��y�lz��c��n�I����u�:�I�{��F�+t��r�ػ��`������USZcR�T,K��	<z,�o}����=w��O�a��`��H���Y�< ɨ[:^Z��B^�HBF��gC9�/r��[�R{K�Ji�'L^���
iy�+���:�����U�L��3[%�	g�u/Zp��������=�o���7���^�&��ߝ�=j��:��A�\�u�Lv�W��G����HG1��r�5V�E+�2��}�Ǽtl�p�&@.��z��ngg��t4�h8F�9��e��	7i�n�b�ҳ3�̒���z�ު�����d�me�PV
V��]9�}�I�<�IT����z��/S��L���ר\r�{{�#V;T�t���а>)�B����B9S�g��T1�<1�W}�������d�A#��S�C���l�Zi0� %��U���v�1�����w9G7ػ	m�S�K�{��v	�i4������U��jgPڞ^� #S�peW���.���h��e�������hm&�~;j�OQ5|�z)�9��F��M��}�B	�Z�����w)�����Ņ��q^�3��^�%i���F۹�hsG8
bZZ�&���퓞s^��l4,p��|�
_d�Y*2'�m3��ܮ1_���Z�#ʽ�yn2��o��-y�Z�`��V�]�l�J;7}yj��۪�z�W(�P��>����[ϓ��3pC{ڇ{�]��w����~��0yұ�&��?�in�c�{�zE����z�z[�w�;Ю�8ޅ�U[�b�����b�zAg�z���ɋ��fR>Q���<���b}(>{A�ܺ�ʷ.ngm��Yfm�(���|�����(�
�2u�U&\��@e�u�t=�c�Ƴ��hwj�6���V�v�J�_7�ԡ&��Z�1��'mY�PPw'-�h�wu㎛U�j·G*kǐ�.���	,ܥ���pA\W��I��Ҧ�p}4^b*^�1�s�0�����U{���2��C�nm��B^�e�?�0V&ŵA-l���[k*+�_�+�L_�KYK�;����Oy�w-u��򱵔�/�lb���j�֞��įr�U����V���x6ǟ�
�Sz�iZFW�A^������$����k��ݱ�(���f[)�g��Ȟ�E�1���!{���Y����Ī��q}(R�R�A�I�K�C�mo�祃GΜ���ޔ���I��������vha[��x��D��aV��뇵�D�k}�"J�/�����y��Kew�N �w]����д�?��>�R�_�:"��%G#8����ݿT��X>�aN����jOΡ�o��<�WT(�p��q�	ޞLf�����xMyr7C�k]�D�^��h��`V����C;sV�h�<2�*��2�&V����0��-�x�B���C��ee*<<�������(w�r����ъx�OtW� T� o�%T~SF�@Gf�\U�i3��,�thBP�\�Wc�{[�/�A��qS��8�2}������nK�T����Oj�]QQ�QKU�2V���c}�-PG��t����w���4
1f��qu,�5z;1a�L��ĺ����{�v�����W\�7X�۞�r 6Ӳ��(8�z���AM��u��?��7�^ͻ�)[����S�}^�f�@����>�F��|��M��҉V��)������p�w��ʶgW16.S��4{σ����Q[���Q�77�|�N�p��w�:Ӂ�����+��5vd�4&ǲ]�b�%.Xԡ�0��^���?M��c9�*y�wZ��#S��x4����Y���znZxw
⇱��uX�%���U��[�>O��7�{����%�MZ��JF����`�CD#^�/b7x�.K��l9��w>m��1��K�ξ������E;:�`�D�ǥ;��k�U�4S�����%�]3�!�oa�ް���̏-1��;#���0��9L���A����Z��%�����<؍7���=��٫hۧ�W���ݱ����9Y\�}��ce$c
E<;��N/s'9�X�E
�����g��5�r%�x�<��t��|�
�ʸ�r�%�Q�)���Z�[�N��"�M6=��0�5��Hۦ/�������ɪ�o�����M�;��ҿ�<R�k^ضoF�I�dco0�ӷ\�����cʺΩ�u���*���b�zf½���1V��P�sn�wn�uT�s6d��U�Q(9]>���e-%��
��Wz��x��b-*���g'��������r���y�-z�@���C�w�Cd�p�~V��?����ˣ���|0G=ox'��h�n���?}��=C>�`��P��]Nߕ>���]�u/>���h>Vg?�IG���Ϲ�oLD��FBAUMJ]5/I���F��"�u�<�oZ[g%5��-c�ۯ=u3�e�^�oؽ�5&��^;e�r�
��DtV��������	ᕦ?]m{���ga79�}j[Pxe�v1��@�Ť@��<�}/fǩ�f�~�F�=�[��x�I�|���2�?w��:w��zlc�5C���K�L^󕝫ת��ܴ���֦qK��ةv�C�ѷ�B�Ţ�0U��r?�p.�_�(ba˄z�/=�4�v�G�{�O:�Njc�FP�4��Jb#���P�O��4g$l��[���}1]/y����&11K��F�H�㎦���ApxeP\oh�<)\�����_�N:͇��IkEνh��\�����pnS�m����D�_p���Q�v���x��D���o��j�Xm�<�M٤�ːM��]�'�I�g0�+
���Ӝ����2�(�t�P^�+N�:�h4��C��9K?���UQ�`{��5��w	���=<����ZU�U{$�^F./�������;�®�
�B}�g�t�	R%�%��(z�Y�4#
{��!O}��I��p0��SPAR�����CN.`\<1��pn�a�F�z{)�b����4i�IȝL�;�S~]k�}���#��z:]A5-�Nы�2�w}��;K������Qh�|:���Po����t/��\����Z�!�)}�ϕLhx��שX^�*~���3U�Bw��`����w���p�X3|�y6�c(N����|�+��=K	�O�é:�zج���SI�N���V
3}u�����ߨe�7V�t��,AX����n�v`��V���署{fE��)�� MO�TI]Ү�mT0�m�*��\�K��9��n�s��AS��+>���sZ��珗�a.f�Cz)��/R���K�'��t�3�S���<��̗j9Ca�u�d>�yh�V4֐� ��=c�2��F%9z6n� �k+�(~��Xܸ9b�HV�5����*H�:H1q�a�r�W�1&TY���ٙ��b�#�y��
�r*����e�lZ�+)5-<���:5��o9���`ęM�� 4E=yJ+i��x�Z���ﾯ����@��޼)_��7��w��ǰ����>��P�|�%"ћL�67+�\
���FL�u7$��i�Tkw�)6��9=lZ�� ��sV����w��Юi͞�|�}^O;rG�����yW;3~\}�{�7+1=��ē����q֗���}<2�g=s{��R��
qTȹ7���noU3Z�S�tut��&V�e�u�y���=����]z�/��h�h
�-�ﴱ6-�i�)�`ڦ���E�;����ì;���a�_*^����ߩ&<.�]�ad���g̻3>��#<�W����uQ!�����x�eĦk�KwW(_$����k�LyE�ͪ��
�֞�����#빵�m��ힾ�g�:S�x��1�/��q�����Ϲ&.�,��,�G�46:�x�q/�e-w��������7��(`2�_c�A�t�78�Jv���q=zs��ޏV	&<cl�唢�Ҹi�w�6Ⱚ\�р#�:���I�ץ{[l� ��C�\$�����We��W��$w-���2��yu,�V�_�!����dy�RV]�n1F�>�%�`�g�F	h�Bmf�)^��0����]�]H'�6$�m�@��0T�;*�qښ�3����7Fҭ�΀Ь�����צ�&�Y�HX�Z75#���f.@_���Ik��|�>����!��y��̩��j��ç����/\�n��g]ͭ'��5mǹZAD�	d��ܵZ�y:�\�8�*�ѭZ�($8��c�7�����Y��l��զ�[��2���.��:#6�	���@�ɺRΖk��r]���a�P9�����\��
�C���:�'G6:��oQdڹ2�F��i�A�`
��շ �a����ɵ�0�=�F��0�YZT(���r�#���TW��N�@��
�nFh�ѐl��Q�.ߙ<31PY�[�e3ʎ�,��
a�(�y\'hx�:��ä5--H�*FA�,{6m��1���았����9V�ȹ<ޔ7;�L3�QPڮ.�
qH.�m��Ś�V*-��*^�Ύ�������Vd�BLZ�2�ƾ��`��wE*�ڊ�u�b�Ć������/��(�|��*$�W���z]r�!mg)@h#[vvf{÷4���t%3S��͚���FY�K��/E��>M���'��x�aŷ�c���pfU:Ư��k|�j����h��� ��׹u�W�t�P >'�q
����MD<kD���$D�ۻ���I��a�Ucs%M��N��v,Ƙ�K�6�y�[�̳�ֻ]��X�v�P�R�fJ�"��G;��]�*��G��=T��aTpHkphh��`1���J�_E�ה_iV��Q�$�OoJ�L���jo^�y�۾�]Z����E�x�=)�'�I��.�\�g�k6v7nЎ�4~�ݢC6���I��w64t̘0�a�<�8��˒�{]:b�XmG����iB��)G[�f8���[K%km�n�.��&��f�D����3���Ĺ��/�&[y��n��1�X�AX���lYdS�-��sq$��r��,%TW�ʲWA�/�T�x��b{ή9u��[0
l���W%�h�Ȋm8Z�]���K0q��_������z����.-2�֘��-ok.*A_R���5]�a�<�\H��	���=j����L��9���M:c�̻,�Wa�&u����ӡ�?k�Y�KF;�ތMP��%wB����:�e���e^c6��&�ti,n���Mf�n��k5t�C"ٰ�Wob�����2�q���f^N�o��kg�v�n�*ӭ!�!IY������r�S�M�q���	� ,�u�����=�кw:oa2+:�k8���f�R(%Ч�ј*�y�D��Sx4��+�����&����K)�7�ι�9+t�	�;��T��g/!�}��" m��ZQ�*�,v�(�b�A�slYj���AZQYmAQ�"
�b��[�T��1`6�C���DF)��#�V��DPG�DJ��"�TU`1UUH�2��(�F+�X���.+d�ŌQUG4��kE-(������ �1T��8,*(�����2ҫJ��ł�c��(2"a*#���QA`�**Ŋ�E\Z��TL�$KI�`QQE2� �)2Պ�mb���PU���9j���j �bؠ�A-m�si��X��a��0Ū"��DD�R(,DU1j+X�-�
�("�.S+QQS�Ub""ZUPF
(�QQ���(+�� �-b�����X�V"�#�F*���V
���E04PUb��>B���{o�f�|2�kG[P��n��c�oE'k��r'up@�$�ۓ��$��)�ܤ�Zt���⻻[���l��+�^�"���;����kB]^8�������8Ƥ�����X�SU�(��K��O2ԬzR����mx�G�K��E����A�a�h���J�]P1!B���({��VyᏁ��#3������.�x�tK9O��<s��8|'��YC���w�, 5s���P���������h���`���qE��v�J~Un�*|^�̇jѰ!��~m�,S;����� "�\i>�*��u�W���u���v�cdp��IViK��d�5�0�Ժ�5�YG�N�b��Iˆ��6/�e"wV=� 4�_�)~�FŶ}�lΝQ��5{�	oiӫ�^���������a��{��?<�h�^��^E��}QY�y3��Y�`����6�'��k�2�,m�z���0��}�=�{��˼��U��ڑ�����~ka�n�z�qu=���uk�Ļj�<�w�ޖh{Ϻ!q3yĕ��yx�"�NX�y�0�"��{�K���2XϽ�w�rZ9���/q����ר՝�����-���l�z�edv9�*�\6�m���3ͣ�q��w������t��Խ�9Nv
�O1�;���Z��sP��t�B]��֠�t����Ǭq	t���U:.ڋn��xb��ID~�{��3�ǳ�,/�e;��	��v��Ϛ�<��0�|��~B��cʮ+��b4�l~��w�N	��3z���<#���vk>�[
k6��K �(u��������}O-�ܑ�6���.T�ǩ+�1��_���&�	؈�*�����!Vϔ��<�VY'�����8����L��M�ъχ��Q����P��O�d�#��Uu�iR���p��m��y]�'�}lg˪�1yhVs��@k���X�^��债��t�Mw9ڥu�o�Y?��q�Q�WɊ4��:�*wQ��0gێώU���;ᢂ7�*>%��|�*G�eŏO���0A����*����Ҋ�]IץV���KN&�W��<+V����k|��R{w���O��#η���֥�9�ax#r�
z�Cz�x3��A�)|Ɉ�l��^b�d����^��ʟ9��C��Z��@��P9N-&�F�T� �P� ]6�:�n�<��{�r�1�I=>�ۃ�TPn(�ڰ�<�=�=���~J�=�5��i��hz�yNҋ���+][��҂v�����Q�A��;[�J�iǒV�%���ۭ\Rb��F�3+du�V��/��f��vN��q̖�m�t/��od*)�2�����28�ǜ�Lo
���eވ���r$��{�����7$]>ܦ-�x/�|<�<����]�+=A�,y��TP�<���wl^���ש�k��l�~���=ċ~�d.Ţ�0U���*��f�����bb$�ì�����]�OMp�<��z?y<���x�?]�lR�L�#h8�>9f�\�e�w�������Of�7�e�Z)�WF���Ll�с�,�+(���6}6�11�~��p�>>�CX�|�ή90(��Ny�����*e�XʗK��N+H/&��{2�����^J` T�੊��֖;9m>f�a�aJ�B�51�x�CsX��靛;:̐yQ�|�q��09����������kì��B��K�a%���*� �գ�fz�
�T����O��L�^<��a7���%^��Et���uK��wb _jV����C�Ԝ9��az!���Q�(]w��aux؊���ͬoȍ_?Es.OGd�ir���D� Ch:qx*�v�����y�0�����l�Tn2Ϭc��;����#@�l��$2��� =�?.X��Zjr�Hj�M<ǫ����A��d�\x�.�0��d��;8��,ͫ޸��W%6��E�j# gz�M�m5��rvƥ��y�B�[zfv���Bۨ�-U� rpY�着�f=6�==�;���>� )������ߨe3	�F��W�ز�UCX�����?=ͻ�c$.��;�dܵ��,z���r��i8����]<�e��H�6���o�'�K��m���G)1^��mh�\�|&[~�Q�h
NR���x��)pU��:��k�֝(�Bp$*��=K|^���`���b'��Xa���&}6O���O�b�Go��M�@̊�tKv��4A_NшX`o���*�c�ܢ���|�:`���^L���	/����nƱ��L}��mU;�N�Zu�=�,�^��f����]C�[��K�Fk�2E�}�Ӷ�A��ͨy_ϯ<'�ӱ
�7��S���4�����甬����*<��@wg�z�Ԡ�P�ŧB�K��W�f��1wL���~�%���7x����R�6��vJ�Yjy�*����+��r�b�����\�!�אw�&ھ>��kU�۾�Wvr�7�L�"y�ľa�U��gB\p��%��`cYvgN�&�Q�Q�n�{��9�/]1G ��(f^)���F@�!�q �X��ngQ��W#�ڌv��*�ovbrZ0�Sʘ]�8�H{���z:w\�h�sz"��,1\�:�PyRf�f��*0�W��
:Y�"	�]�cdЩ�0�4GV��fC������R�r%cG�S+�)�-۳�"��:��g�7��2X��,foָ`�+<��l�Ƹ�eW�������M�w�
��c�+������E�P��v����$�j�4?	���4a���a�>�-d����7���Pf�/+~�,�����þP�$�^���X��,���^�1*���ʥp����Wsz̝����G�#�>�g������Mi9��U�{�(��Hhbv�kf�}]��,mY���_ߖ
I�z�+HW�:�"�џCY��E+�s����h�,_�����74g���VH=�V��f�����)���&ӫ�0�Y�5.���S�8��2��@9o�ֺ��^c̓��r����"�
��#��D�X�9~P���V�`]ɋ����bBv ���z��5��T���޹��`�.@�������u��6��Y'�4^�/���h��f�Wc ��03[�61g(,!fVy��7��a����@6}SԈn�Uk�����5��;7�!<���Y39�+�
�eKޑuge\���\	TR!��~�V�c���.��l�Zz�tJ���ؠ����v��K�	�[��.�)�/r�rFʤ�Uͤ�a#i�{{Mv�GNp�h6�ﰊ�Zɏ�V��I�d�I~��Y�+�vnG4SO�a~�.R�*����^=����J�;��X;�~>z�܈�ފ�hN�wr�~��Nӎ=-�9Դ:�^���xcp:�p�]�z<�^ݽ���(X���uS�G��}:1�:�3X��x���k-c�2�.��������
�������`3���)>���ƛJJ��[�3z�����K]��	��z��6���X��;�����@a���>1��0��K����>i�y/�ݶ�?cU�u�0b���a�\�#���^E��Ʀ��Q�����y'�y��d�ʺS:h��[�'�I8lq4�O;)�ֻ9g���]6]e�5^�ǜ4d����S]��O�0h�I��`^����3����ȱ�_=y�bvo�^t�y�9�;=��~(O_X�V�CB�I�q�X�z]�8�-�^N�nz�-OJ�%��ۋ]���N�w��yV�@�ꄞ����OI�s�����>��/��򺒗�7S��P�e]YG��hw�����!��%N�Z"���]�^���v�%�C�
d�� ��,�c�����Ё�vѳJsC.	�ڮU�T�i��o.E�h���/��g�jaU���C%y+2gb�7Pn�P�9����*`|uu9�ާ�8?�����(��� �fԤ��W����伶���%wy@y�lB��e%Z�{r7z\\!u�d\��8:��VZ#�v4a>Z{�0v��\�ZBN�kZ�g����k)��CcV5���{`tX��+�8�z�@��n>�Y]��s�����α\'�|b^�����c��˸� �P��讗���q/�VKmZ��}D�~�8�0��F���u����f0�R^���C}��_��|v�9�xoZ˷�;N�}�s�mW����yQ۝XB��²�
�U\��>�N���	��[��9�ݕ��'gz7mg`e+���O��b�OG�'�cӶ��A��̈́z��
�	yj�b����v]����]5	��ܠٹ1�b�;���[����Tb���'�}ěx8eh�"s��Hz�A 5��l�֘�g �����x��x�ʙb6�?�Z�:����ٴ�W\���݊���t���a�-|K3��"PQ��Z\��^�j��Z�$0V�Z<-H2P�ݜ�	�cB��{WK:�\"��.�7m�Cy���_ +!��4Zö�ͥ;0��Z�)8g',��-��������rV����P|,ݨI���X�����F��Ѽ������b���3Y҃�Y�GL���W��o���kr�R'�o	|2�e[��&<h������V���Y�F�z|�o����'^��w[�O��\<]��|��y�/�Q�ԱJ�vT,_���g¯�%�l�������os��ȴB���^\|n���"�}B;�� ���0����
�T�����*{̤�3�jl��VEE������!��6����_�0TT�<�0jun_&�M-� �L�?b������.Pk®��\�%[.���Q]���)�~O�i��ң�U�nw�أ�#Pp�'n�a���٢^C�x�ig��'�!�eX=8֚Qn{6b.��4X�:��egۦ�XPS#�!�X�C);�|lnS�gޢj���1TJ�ӻ��	|Z�U ��x�:ͭ�g��҉�p")�0oǩo��K��gE�K�v���O��{���7'ҷ���柁����ַ��N�%tw����_m�aQ�?P:{L�.�z��1`t=��8�����7�yH19Z�{��knu��ѾwkCZԮ���d�X�
ѵƂ����l�ހ�ڭ*f=��y;���A5�v[��H��:���3�.m'wr�fv�B4y�;uo�̶wWv��w%Ʒ��q�e�����t������zц%�{�R1��:�ۻ�� ����~���^����MxG�~��!�Y+�g�����tuH�xV��t�W;`�>���gO>�:�a��w�;6�]��R�����]��~�YuV���xl,6rz_�Y=�w���^]���8Φwx����W.��D�b���b�X���Z5��>7�Wg���;��;�B!�<�����gF�I��1j&OeyVZ��:�/3���+T=�$�s��
��l���F
��T�C�'��55�x���Qg-J��:��64�R.m�'�;v0TmM=�����R��>S��TϏ҅~�D�(q,��&���=�G8x}��\�V������yI��p���vhZ�_dd,g
$PSވn�(�٠�}پ��@@�?}C�x:�2x]3��a��i\5�y���v�V(�#5h�*!e>�陳��<|%Q}V���mu��ߖ��nJ���5'�P��JP�Qȳس�	��5߷Ŝ«���o���P�})-R�r�j��\5��ѥ��m
�m�S�k����T4�2��G���&�V}�T�PTwp�WrE��=8ޘ'nR��on��Һ\Y�2X���	3m��N>{^}(y��}�.�s{{\9w�'S�ͬ{����<;�S��nR�O.��y�o�.&�'��/�M��sSa��u��G�_[�R�IKF�*�����N��ʣԱ�Oҙ��_�x��Z�T�,"�ܝW�m9튳�ԣ�	A�j *�7Q�
��J��(�^l��?*�L6E���&��v�^�-�X����aC���aVu]^�0GZ�%�OnC�6)P,��ct�t�>���'�L
�N���7��Gt�3�t*��p��XѿOX�
b���uӚ\���y�dy�]��u��qæ���j�=>��C(��^�y�
���ӛ�ͅ);��p��u��u��-�բbXʝKC����& C�x�OWv]�^N�Z�8�b�_y�v��*)�����u��﮻(�W��øv���txz��Kϼ����˷ƫn{)���eGz���Վ�/�����2�."E���Lǯ�c��aܔ�
�	�����6V��x��xO�w��C���/�����.P,e�Q�<�P��mE�q.��z��P'��2��W��}�Y<�^q���]>���'�C�"ʩCFv�-\��F:T<EY��"'@b��gG�A�\�q,�`�8��Ο8��f�C�1����a��xJ�Y(oZ�lvI�Z��i��[���T�,4�9S k9w��Nޘ���Y��rozed|�,YJ;q5�6�A��ā׹3kl*'p�d9���/r��;�*b!K�qCۃ���x�'Q����E�5��=뼽���R�ؽ.i��*}J^,�I�\��L�Q�n;y}[��")Iˑ��n� p����V���c�v'p���6�u�R7Xx.�v�X��y���5�0�J`}�f^+8;���cTKՂ��)�
YO3-=��p�dGx���#}�v�BbBu��f2���7b#%�7ϸԝQ���^�0�����TD �E�'Z�]�e����G]�4䆥:��e'oF�j,��l+9o.�!�k����l�Nugo@B���[���w�_r,�}Sh��e������F'�~�&1.vSt�:���@�(Q.h��Ѯ����[��w ⻔5�&�BWd����/�ܒ�ɶī�C�b�$xw'�+w�Ŝ�!l�6��M�x��G8�W�:��yڋ�	�`^�@� �R�+	7.�3�����Uff�#Kݘ�b��WBu�a�6�U��!s�F�M��c��щ:fW���6�b�WE�+��0�K{\�k6�\��G��bP��D*� ɥ��q'k��E<;�Փ2�a�yN�t��h�+b.;�� ��zc���Uff��7��^Nj	L]����}[�JӍ��t���^��QF;��۠��k�՜z`[Ӽ�t($�C`l{�	�2uH���Ql�e��l�7q�Z����і�U*}L�Mr
GQ7�,n�.kYo�qV~J<���ޱ��BG7S^�sk���sz��od4݌5��4of֫G5��Νt�Y��K�g+�
^\�Pc��ъV"TG�����s'N�%�U�J�lY����v�h�Wm�B�	l>��\�1ґ�M��lw��
y�cۮ]�)g
\-�WR�uDO\9Ƕh� ui��R��~UleWY����a�(��c�U��%u�9")�Ws'f�PP�R����*4�ka�@�m�7�ST�8�<���ƝZP�Y{�(����z �I��6�W�nF�B��Pwj����;�s"���-�DxT��Cͬ�k�W>�����㐡���e��ҫs���{�O�m9sr�`˨�Ʌr�J�s���7Sn=��3�������]�4���׫���T:����#%��y�4d��C�B��혹ܻ;�s��e�&�ȞJnîkq�0l�5��]P:}4Ջ(�v��Y87On��n*��mՔ�}B�������H��ΜE�B��p3�"��n���6�`V�!�C�0���"K+i���a��nG3����P��oȓ�-�˼�F���jv��u���Ě���K�:����ক%�'h6��F���Ļq���HS��)�O����TZ�[yM��ΟT��|V1X�"��Q�X�DYP��,@QX��X��Q��EU��(�J�T*�F"
�DH�0Dej�""�QUb,V"��U"��*%����1LP�iU"�UU"�P�I�b��*�cAb����V1���
��a+�"�"�(��",DFa�"����X��1UF#AT�`��V,\0�Qeh�`,�+�"�ĊШDTUAX�X�AU��m�8�UH��,*���W��1b�1F�`ֶ�TV�թTE�Z��ֶ���QUPTDU�|���<=�j�
��Ȅ��zF���9�ņ�҇r����h!�.����9"['Y� Seе��U/V$0��Ѱ��%/���RwߟK:��[z �k��B�/���~w�z����Y!	q�jܭ�RV���m�2olwx���/p&*���ŏY�eZ�>ϒc��{�
A���A���wle3���_m3^^j�1�?���`d����X��IH����5�9�w�h�_G���*y�g
���!��
u�;>��;,�p+�aɗ7�	�g9O[�wL�X����+����=C!������]Iצ�f*뤴�XZg_Pٞ��+�Lޏ^�<i�|n�G��,��JsR�����F*����ȀK�
��ꇱ�+V��ع�P�s>I���S�x�e�^��5P�U��h?��I��F�^�����޽鰢�T#KG���ض�x�鱎8o��p+��Aaz�)��qs�nQ*Ҟ �9���,DPX}�������~L�zt���p/6�����O��r�ez�=�28�XC���f��~R������5���������FR�#񱎸�������*��s|[k-$3,<�]�y3�5)��Ƨ5�U{�R��?��^���j�Z+N�%29Ӥ��wPcDn��Z�B[��������aP���U�V)�q�����z���l�fm���a�rf՘����X3⊋�_��K��-�:���-\z8��PC�{7²r�rzޞS��� w�1��6)y���^��k+6���F������P��Plܘ��/´tn�?I}ط鴠x��|76�5��vS|����װ()B(8(B�=
c]�oZcf���ۜ� +���}�/�ץ��ۭܯ`r�7�!�=���-1�Ę�$W�_O>3�,<����j�ո`�{���⻡��G�qu�����y���^|0�^No�p~�]�a���Co3�S\�'V���#~Gg��m��e	hC�%��P��\�Q�԰)Zlr�o�dwx�S�$�^�W{��y�R>���Z ��y�xe�à��BC'�#�gJ[�^��ui��Ө�J��M|�8������&	��1��WtG���r�VDJ|ƃP9c}���߰_[N����_3�U�Õ+����_<�)?��7��{B�:R�7��IY�[�q�{���Y��5�i6���������ϵB�PIW��u��=|�ѵG-��u���.���%wAh���)�,�T��&�V��ǂ���9tU�A�����:��f����Pu��<�x-�I��i�jjJd��a�����(uu�v���B_es�s�e��˩QQ�A͡y�ךᇫ\�)\��,�*�=�$��ћ
-���N�����N�oﾬ����|�ق!g�[�g`�O���X��\<���˜.�QME(��H��}[wSv�|��I��F��������#�u8"�G�{3��0+���5�r��*fXs��w:�;��h��D�HQϩ��&�?_�kj4AU;F!a��PgԎ
Y9տz��9��Ԓ���5���`^�z�u	���lO5,��������.����k�}yk�/9>����=��u�"��]���C���0�w�j����<"nVbz=��lo�8��3���/=��a��f{�7S�և�.�uֻ��V��,��.�zc���]��}/�Hh9����o���������Xډ1ᒏd@W]jl���vb>(>�[W�b��˿[�M�����R)��t�ʗi�8��ʮ:XP�6"�Pg����{�f�Z����K�?��DK�lL�wr�}�i�u9T2�.���|z���.�ݰ���8�GO��4YӞ�F7l�SZ �V��ϑ�v?��3+��o��q}�)r��r9b�r�<�kyt y)!�u�(%\6}�Fp���ͺiN�jG=��(�n�-��=W���{��ȥ|ѥ$a��V�Qj�;����}Hi6��84V]�9�i291�j���k���Z�[�i������|1\�g�ٸ�5����;R+
����� V�v�ի�����۷���V*�>�p,[��SfF6��9�]4�m��c��RYn�}�y�@D �M�����D\�Pm���ʬ��E��т�{.ԭ�&�տXQ���P�n�P�G�R����c3).R�5�ֆ6��/�
�-��9(���SWd�/4R�e<�Vж����$�J.�xͤ�o�S��_<s��s|/ٿ\4�m:�-L�Bf���}(��{���J�����Z߅Կ�F��ߑ{�֏Y�3���sx������L��`"W�� ��������¬
r �{�!�T��f�M���91)�B�8/]��qvSߖ1�1��x�(/�,��w�ب�W���Zl�eX �\�5&os�%b�к,6�kii��6\/P�j��rm/��$�J�:��=Ys�{��'���Ɵ�xS��G�㗁�,���o� ^���s=�½��G�� 嗒��)x���2�c�f�K�m`�V�� �w6��!� �_t��:�7�����ӫ�#�C���[�R��N���I��*5��f���/��Z�f���ֽ|����K�]H�(��'t���d<�Ls7.�l�c�@Vb9���e�g���3�tS:����<j�AK�k����b���u�B]���s1,�uw���Ȯ�	�5�fL�����*r�Ƚ��	����a�/�jY�v�oN,����m��o�]���>�3*�3����S��6��s>�*��^�᮹��k��y��y�f;���oMK� Hi�ʇ.�%�wՑyE�,�L�f��v�6��,�D����W��L|���hz�� 3O#LZ��Omvr��U<��+���Q�GL�r��=�'
�|5�A��0%��^>Vk�e�W�5�2�{6�
\w%]!�}<xW����n����N�b�T�B�|ǒr}P��W�`[�Ƽw��0b�={y4+*�z�I��ܙ�o:�gA�R�A�$��mAF���j'J���q0.'K��&Šu9���;�Oo�-1�ˣ�aCJ�7��p��w��/RU &�S�u}�ˤ��ӫ�~�)@�ʸ�F��+�(�4U���j^�����˨*��h�y��W��#�Y��ï�S���GW�&��
�]:Ѵ�����N�B�X3K�w��r}��k���J��T��C����@Vr�5�m2��3.���y:%v���^�F^��C/��:/� O@�<��&am�xKY���v=(Q&Ff��?{Յ�������V��^Ŵ��q�C��k����8p��K��p.�d#lk�J�kr�.�� �l�8:�=1/Z�9QA�e^8*U�2��bf$�&�5/ܷS��R�w�`�tm���Fߘ����r�NW
\�J{�/�]q�=:��&�a�ʅ�/|�l�e��h�>�m_�e*G�$���������)�ӰvPzx2e{��\�!��8vz�׏	����LzV�@o`O6(��=Ȃگ��Y�N^����_��B��(0��t��[U�8v����؋�Hum_	�^��+ޮ�k�;y�I�-H�� �������W�z���]z�kLl�P1���%]�sG�b��e(�Xe�wIж���%��ؐ��|.�|�Lk(6o�S�U5��"�/=H�{�Iţϛ�G�����*2���lx��A�&=H����a�&C�{�-�5�;�?�/����L�X"��ꔘ��y��"�ǉ��e���H�K��)+���}HՅ��Bwf>�jೊ�rJ�nʐ6�n��=�w��yk�s$���RT#	��+��fK2R���9BY��ჳ�O�9��R=�n���S�V�L(���)�.�,��|��f]B���Nb�r7+����i_M]� [���kN齰m-��}4�wۮ7�-K����*s��A�6�����1�ZF%�x�}J��u��z����+P�9��(g۝5�s��S����Ϊ��{,��V�2W,u��������*�>|4EM��Ny[�~��{�������m_�x卨F�p���H���-^r*>��E��\B�8�o�����+4|����`ݤ��t׆�����㸳Q�+e�}�@�CJ��fj�Hn�����3�#ax"`��OE�:��k!�xy�o�B�}�jz��d>]P���OvN,
�t��t����Q>�"��g�o�'��V�dY_
k�����"� �oy�݃�*��X�&W���Lz9���^��tX����tN=ׂ�Qg������f�٪�lT}���>��q��<3z�U2��>���j�ZV1=d�Z��+�{]��d��;��Q���bۀ��Ƞ,�|yU35qظ�uYɯu\�n��c��lxe��d�N��@'���b8�U�-�x�-p#�et)�F��3�r{X��H|�۳ZUb�L�X���O�ז�~7k��h6���ݚ��p*ꔝ=cGgD�Msxb��C;�8'��w�r�;��E���nu�4NT�Y�`./YC&\�Ҡ�=��f�����{�9��������m�ã>����|���*��x�=W]�hbcD{�4=e���'�ڭU-y�+���tc����?j�8��ʮ:_�<������\�_W�<w�9L���"���]�Y�.f�T+����-4\B��m.��n��~��������Y�ܝ��	J����Zz|����g$�Jx�%�o}C����^}u��Tva��*���by�(���p���`L�����Q�~w���/�0@d|%�6b>%Q�n-�gtPBOR�"~'�mK����a�˞5��o�;
��l��}�]��v���XU�Հ��#��:���D\��p�p��el�k��i}�ʄ��4t!zע�52��S4f�������/qT���R�wPt3�g�p#��#�ic >��13ײ�����ހ��}-ء6*������8�U�)h�2�/�Lk��Ι���	��k�E��[>�C� GTxJ�@F�w��%G�u2�F�AEمn���\Z'�^`�N�fN����v�q����zz=<�����FlyX�V�k���v�-��j�[$�8*��q����Y������^"�k�Tww�E�0��6���IC��bKٝi��J`�έ�]J#ʺyȰ��D�?{qWD	s���v_��t�貶�{ņ,@�D����L�R��i��5�ͬ���S7�-���C_4Y��Ǡ��귑��lB٭�7�,�Y���(m?K�Th`g!j�s_>��`�h�k�$pN���֗r�ø�a�z�gyD�}c�KN�
��9)K]KrzUs^0o��r��V�w�c��烺N??���,��}r�,f�$�=Q���t��sѦU���|��m{~1��{9��W׎�||)�~ka�m�a��Z��Ȯ�ԥJ�뻘s���Z'��1	���]h�k��� ��i��񐾵�e5]n�鋆���:����[{��)��v��]:,*��<=3ފ<��u��<vg����(A��ј8OZ�����w���i���E�Vz�s�xJ�[z(<�V��=׌�R�)꓏������7s��@���C���s���6�&���t��g���[���ը��x����kH�^�vWYN|%���}P��A^H(�m�Q>\FR��m���,c2B�HO%��tc�Z�x�y�p��l��bSބE�!�0�����-ќ2����y����/��٩ff��珐���u�MN/���%߉yqf�e�e�����n:�O��`�ʶM����w�,�e�L]�|�\U���1�k0��D�G굨�6gzY���3%O+�͈�T�tɺ��ŝ�|N(�-9qp̠i��" �r�F�rq�d�*���+���\�*B����(д��N��ϣ��|%�gJ����cדv�m�}�s��
}9�c:�V0([C�W����v�H���f�N��6��{�z��N.�7�	�U���|���<)�T�Ϸ�Y����A��j^��^�]sw�.�{e�F�;���@kG��U��m��uӹy���:n���U����u2���4Oݝ���}�
Ź�9�c@�z&�%��������E�(W�C�ålZ|�~mֽ�n�OOJclv��VbÍ_�#�o�~L�cb^�6�_P�n��&tQ���;�{�?�Zp0��	{���y�������4VT�R#���R�M=��L]O�oO<Y�۹�5�&����WQ��w���<�����|e�]/���
��[#�kٜ��^����i��ρ񿷫�{�&}r�˨�6=;���������˴��m���w�V���NIO�^b�2��[.޹^�D��/�樇�^�*ѻ�#!櫨�W�ܼJ�������`�u3.h̕�N�ث�R��:��.�Uwg��F
�=n#n��b��6�Yha�O��� ᔦ駲���!��m
�U�i�z��*�=Ū�{fI��R�)�}ǠY;D>�K:�ீ-�����AZ���w}�9����j��ܖ6���v.�����5��K���a�YCf�R�#(汔��̧:�Gfs���ض��3���2��^�VG��z<�xԚ��5�s'N�WϹ2Y��ʡ�V0�J0��VK���k���!Q�H7/2�s*�{9k� }
�2��Z2�v�+����m�4����wj������hX��u�N�1؛{�t+�p�ژk�"*n򂨬]wH�љ�V-֕Σ���l���Њj<�m�[��ZU�TE��.�LҔ�J��^V�vT�bkkQ}�U�7iY��R��w�nA�b���
�`;S��^�g:�k%'uF���흀-�J�H�:%y�� ��u���5�72AbD%��'�7V�̣-^� 9}���3�K۵+t�q�,�!˸�{;�y�B�p��Z99P<�Im�l��.��bS�Gb�e]�9�EN<����7,�V�����d���BL�U�4�λ7(t��"����۷ab�.�v���R����u3A���d��o���T�7��;:�df�:x���_f,�<�<�V��9]\ef�r��ʼ�q�Ȧ>[0�Y���#���!�#e˖9�d)W���U�+-�	+pv`���5w��73�r�rV��|�n��3�7%��r�)sf��@>����up|)���4��:AA�G�N���߱Ĩ��]����3[�ѷV�����b�uU�4�;�K;��xv)��q7I�V��Mn����t�!wN5{E�[��0�n��W���Ք���i�iT֊bEc#�2��c:���,odW��o��sz�]�̉L�a���.L���Vr\Xi�(�C.���F�U)y�l�w��;�\%kYه����d����)�'b��9X8��0��V\�B�n���\&1B_f�.Ȏ�raif�9��2�����dk�{Y�᣶UtoVCԜlUd`AĎ�ͅ�o*�v��bP�"u&�n
s50#�dV/���VM�:�<U���:W`d�
0��.��J"��O⵵r�ĺI���gU�w��o�UĶmB�&ӫ�Q;�E�mfc�2�J���
�����j����LiW-�ͻQD_w]V.2��N1��e��f�-���I�Y�U�7�����5��Υ4�:(y&�XuwJ��v��.���(4��c������5da��Q%�n�nGZx�F���Ӏ���S��m������(�(��y�9yƹ�}�Jw��f5vCu¨D�RUQAEPUF
,ڪ*V�DTQE
���((1*UH)TPDX���*�(*"���E+b�TEU��PTUFETQS	X(���TU��1`1T`�b��VG�Z���T��,�QU�UjTQb���iT±T%F�A�Z(6�,j�l*V��)Ufc�Z-m�R�,X���Qj��1��,QdPYD-E���QC��j�-�UE�*���0�D`���Tnl��0Ɖj"J�����iZ6,DTAF*���+b�Ū�(��Y���U�/�9;�A��|B�몘�<���B�s;y_#C)�湰�c.M�_�pۦ�tSiv
S
�3t:^��
�q�G]Q�n'`��e趴Ɔ����,F=���F�*&t���X^?����R<)U�U��]k^2s�X�`�U'� �ew{�V<��6o�Zެ�M�
L���wJP���ǫRc�H�_'����ֆ�4+w ��q�ۈ�&-���=bsC+G_W��UB�LjO�|���>:�$��d��F��eTU�`(�ٞ���x�GO�L����fm��sB^�J|Gp�AJ�K>
V�7�X�<�����x�Ĝ�T�Ja������Z ��꼸��b!��P��t�>�͏+7A���"D���4��?��|6���2|�����x���BS�<
�>|�iW�d�k{�>�Wt��+�t����Z�ZP��:���jD���1�����<�hzm�<�>�7�׊��Z�:'�A���2���\w�y����J�1X{�k5Wy������ɵ���
�.�xS#�!���\e&/q��qI�B��l���%g�mo�dkI�
}!}�
ꛙ�r4t�n���z����Ybq�<�|8���=�&��jKXiy�g����%b��uv�(��Q����7[�0�LQ�{�\��F��
�U��}Y1Y|�μnV���XL͹�_>�u[F�b��އM�&�N!E����Q�ʂ�C�C����g��)�3^�<3�W�͐�ù�(_�'��ש�%};E�a��PnpAY�j�yݹ7���<�Z��<�g���\b����r�+*���`���,����=eK�=��fb^�/ku�|�2��Z�?�Ey�Ǖ���L�������4̟[�++<�Rfo%����z{���WS�z�-ځ���o�]
`�D���y���>X�U��p�;��|�$_1��������ʙ�O�:7�&�m5\t��~�D�?�����S]������8Y|58����i��B�x�9���z���EF��q��� ��	����U[쓛ո���qF��=d;��!]ܭ�Qi�uP�"��6�.Ӕ%����-���r�w;�|�C��Yڴ�
��i���D��zpu�b3A�Uk��h�	�c�m�{UX�{џ�:���/jb�p�z�(/�9�3�鎻������p�Oy��`ӑW�ʸ�����wP��V�@W:tO��5�6d�l��J^U��^4�u+z��W���g�%}�Ⱦ�"�?#9T6�A�h艗X���:���Ob�͐4E���}�g[!e�-wJ���N��eN�]cIi�����XӖ�e����n[֋��'���3\���_�B�Ώ�n���_ªh��<�K����g;����������.\-U��Ma�򁷣������]n�Y鼯�\t��7`�)���q��n �7�%�\�HXc<LE���P����~��z 7���L�5����eL��Vи����&��̱���ϒ�7ݔ�W����)7kq{6On���}������ؕ|���@�PJ�1��~R�y��oI���8��]��~=�D�.ͫ��]ɏ+jE�4`c�OP�9j�q-�4|���LY��SGa�[�Z�ϙZA{�!	N_�%�����%�^��B�_��ѭW��A�6�p#9x��F��z����2�� �M��������P��ٴ8������O(ݫ�>49C�����ߵW�r�E�`M��)�:��cO����y��r�?�R��yz�,к�[�:<x�ϵ�0���VX�_'�6��MS�����Z�g#��m�bǜcF�;�ή���߲���2{<����>�|'�h�2�А��g�i�o*US�IS��d��ҳua,��W(,CĴ�4]mM�)�RgofC�=ː�q����@�F����ΧC�\����Q%ܸ�[�n�� -A�c��`3ԳU��C8v*x�;U��9#�JS[�$�>;�{3F�#˧9�lS�a��&�G��K[|��7�4R�?}H�6rU���%���a��L`ϧu�7���U��-��:<}�!��Q9�u,����f�t0d�R�
\��P�Pj����%�3��0o>�>�M�f�L/Se^�3�s&OZ��q��s@� >>�s�$���ԇ��v/_+�5S�-�S+d������w�+u�WfT=evp!~�&,l����.p.ê:�1��y�-!��9��-���,�q�	�Sȫ���eXˊaU�>c�`I�B��+�1n?Ձ��gDk_���s���}+���+G������>Ð�R���)�E����:̮߽՜O�I��=z�V.��Va앆��?�N+-�t���z��d0x&�% ݾ�sΉo��;�����B�kn�Ӊ�U��d�W>3�!t\$�R�TԽ&�	��+���u�m%��|�p#z��Z#C;M��v@��<i��u�0�=SU�>;�J��Ff?FV!O�F�N��@�Ţu%�|�1��r��j�Dy�E�-*
	xK�ݷ�۸��kSX�v(��}�I&OC�d��v���ڲz�*]^u�}�G��]]����rԮ9o6�!3mrM���H�]IW�0�Z隕�h�0�pPಧRBE����8���B�������ćvYȐ�2��D�NQ�Q��U뉪ϞD��;��������T�����PXfz�과b}x_�������0�r�b�֤�?<+(M<]j��U���n���9�[����O�v׈������Uyۡ7�����Q˃6�P��b%�P������p�I�5C�鏉ͺ�i��=�V̑����z����ҍ3_8�>6���(n8�b��Xto��>Pγ.�Hҵ�9>x2�5�����K�P�z<��l��i���b�J)�/��w\��mf�D��%]�yɐ)V�,_��:b�k�c�H�
��t���TIwV��}R�q��^��Jtj*3ܠd�Fa��x{O�6#�����>������s��tk4C�ތ`�����b���h���͵�І��JO�C���TR�2r�
���O��{�Լ��v1)|3�lS������Q^�nJz�����VC���O�J�szQZp�T��������^��0��̨�U5>^)��������P������=H�0���ܐ]^awJQb�u4�er�uWNX�˻��֨�q�n�_3=�-��.�Z`������zJ�XYɜ����ʦR}M�o9u2���B�bV2���Fw�-U��_lǷN�'H[�r��{����yZWX����H�$��f����[mi���P�~9</�b��Z|T����d��c��}:�WP��]?O�0�
c�-&��p�_�ɍ����	����(|���j�eA^��	)$K�=Ć��WPK�?	Tv�Ҩ�Cm�E�L���B��A���l����w�; �d��!�'�s�U���T���H�ǰ�O��Ծ�^A�^��_�v5��Ov=X�k��gD�����Y塉YT�ZB��9���ϧR*���tF��N��S��ɒ]n_��ܰz��ƥ�R'�L�67+�W�zg���5�:l{��s.�v�8��1������|���<�4o��ֵ�<G�W<r(��9o4L,t>����=��;�^�+��vg�y�9=�Y�+�>s���SԫC��Ю�.�l,��w^X6��7u������]:o|l��5��X���*�{��gB\|v�.Q#�<73=|�[�yw���A�3�bb���5�E�wV�C�c}B��|㳣*���l�Kk�'��s�䒄y3��(���*2b��YF���xu&��φR��oM���!��Ba.&b�-K*u���k�{��:����ox*��D��%ԫ`n���C�n3L1n�����t��^r�t2�ڃ,r�v!�l����y�H���e��@yxeoN]ۧZ自��0����KZ1�x��u=ݧ�B8��ur�����C�qOמ�����E�LO�X�ڴ�
��i���b]Ov?��38�l���a=��o���*/��-Z����{����T��|�L��om;�S�pn�R��}�aM��c���B�|4M
*�H
UA$�7�r����a	��5�b�5`�c<��������]�w�6ڰ�U\���s�a.>tE���>\Ы�ڵ����t����ɝ�/�.�7R��q���5P��8Qt�j�^(�Mr.�� �8U��tn���7����b83� �����uuƥڈ��j�ZK����w�8՝SJ���=��r|u����S��Y���cB���Q2���j +�V o������~Vk������
��^,D{|���۬Ul�q��!�(J��_V��(1��p������u]�xIM���^
>�
�7B��u�c�sj����6!f��Ḡ!�i�̍��7έ��'���(��]L���v?u۝Gٗn��YViR� $^ V�V���S-놻��wtb�:]�1�HM��/(�ˡ��^�^�l0j��/PN�vZ�L{/*X;p/-X*E��iQ���<*Nr�]��n;�^��.�oE]���%�n�v��BWޒ��D��hߙ�p�OR!wV=�-�����-��;�]C���#H���[V.Y3g�9+/����{���퇓�L|��Jͳ�ɐ-U��b�.��F������ve	<���6}m12�>�^��Q��ys���*?Z>�0�8���a�z�+��7y�u�Q:�2K�PBn���ֻ��R��28��z��j�A�9J&��)�S���`���3t%R>�c���d����P`����;�~�<vg���"���K�+��ij|v�1�ݟB��GqP�S��\s�W�P{�<#�<�j�o]�d��6��q��7��S�4�(u�'| �X����vS߭vr4��v̳:�[�L���}śa�O��E�ŵ9^º����A{)q6<4�b��<�/n�8���ܶ|=�j�˩�u�>̫nY©�d��>P_�)BqE�i9�"Y��e��=��?n�9�w�П
�-ͫ7�1�.D�*�@�0IҺwZe�|]�鞻�J�U��2�SP�	��g�(<qt�tR�VI�em��:۾.���؃F���	�6�	��F��H�}��n����h�f���{y�\z��s^bv'��wA��SXz�nu:��YҶeʓ�$BӘlwu�iT��R`�k���T���'�f������*_t|��A\�l�6�C��,�������^u:|��z����G<���q򺸪+��A[f�;�#/�,�����*H̙M�s2��������(=DA�z��u�[x�<1	�<k>�W��8�P�ᝅ�h]�Ҥ�7�c�34�E	�F����a/�Z(�u��b]��W����g���cp�ޢ;�Y�� ��6F��y����_l�%`Ň��R6���^?^�X6��W���Æ���^��9���}p,z��a��P{��k�ݾ��r��h���!�=��	͞�B�e�h�r��(]o���ܠ�*�h�ܠީ��������z�(75ԥٛ)�.R�����ʱb��g�A���\�f�9%�1��0:����w�H�Y�ѝwz'�ncg.��x�(.7�H�[V�W��5��'�kLlVj��T��[m��{�Ĩ�w�oY2�,eT�N��/>W�\1ąht�C�5o5���&���������P�[�k5��d��&x�wںvG��#��Y���5Ҁ��Χ���k%l
���y:܇3�M7na�r��ը�5�`�4�I���{	�y{Kmɥ�5����3��F�]�(���Lw`dF
�eXТ�W����� �︱��]91-{�.UB�LjLN�������PA�,�ɷ�7��y�`�7R԰�>���4w���ׄB4!��Q�F����5�ӣ�p^����sTLa#�E���lS�%�|?��SZ �s��B�T`�(k[��y7qb�>�ż�߽Zǩq5)>��.�E.K�^��<2��w0��W���=u�Q�v�I��߻�T�~ڤ)�;����|�Y�b�Nxc�������W����/={����K7�|#W~��'B9�?�0�	^5D��S\511{�/!����E�1x�����z�jD-.�(v��=Ć��b�Wapώ�b�V3-�Giv��ݙ�����띊߄����R�� Q�Ү��w<Th�D�B�!|�(.�R���/CG/B��gy��Y�ա�p���[��,o2c�j���Pߧk�u��j7	������X���1�'�P���#�^ȫ4�!���g�1;�/��*{X�����[��O�����]�*]�Ӹ��l`qdv��qө��n��f|�G��e�7�س�66�,á�0U�w��d��}q�\BK��J��A��ux�74�D	��nwڵ��Ϊ���gRv;��{�(�U�3���U:�ǂ+�C �[ܨ+�5Qh��)�3����W3u'�j���Z��C��*�)n�1��,��A�^6ʭ�e�&��x昢f����8��&���eNۃ�G@�\^�GpH[�Nu��m�ڑ�}]�]E/G�f�%���^�݁��(<��zF�K�x��� WЛ���}��޺������)����|���Un�=��2Z(=���\%�e"�!�I�{��(�Fl����t�J!J��HHH�PU�nը�D)�nS��^]�n9C�a��}��IZ�Ե���~6�krslJ�I�������$Ď��D��R�E�4��S�s�XlWN���ٖ�s+.�m il�e�&�%�^:�+(j�}8_k��J��Q�o��T�͓k�s<��6���K%X!�K�*���9Ǌ�x�S[^��tL;�	gk��3Q�#f*�0�=��3/����.1^��uu����7�h؆)I2���;�0��hR�������+�ӭ�6�Q��q�n�*�F���������]2�h�(���+V�*�LX0�X廫[]F�Z�P9N+�&�g\.���nFI�Pk~e���Ek{J������'�(,�#�[���j�KͮL�9u�,�ǁ�S�ʒ5�hV��-��F�ҹ�$o�Nky��=��"����P&���*���X�H�j7SW7b�|��;�{ٹ�h-H���fQ��Y�A�a_V$܈�	����7��ɴD�y���2��.��p�c�aJ_K��`���^����.5��g:��R4T�j6 "Sh�1�:-��9	���Z1��F�*�tģ�K��YX�E^�*s��o��MYZ%]���vtzY<u$(�-��:7��ɸ��{
5�ݐB�t�_9:�n��"]C-j��h���;�ڑ�F��)�s�N�)n�Hh�;G��;G.�t���ڔ.*s�.߂���[�v k[�Za�W�dY� j�9��b��]+9��TM�����)����!���&�1���t(����P�t�Y�Q��u<��D�t�++�f��s��6�s���#(ۋ7�R�E*�Vwt쫔L�6ۗ�n6�m��,�ł
硑����F�u)6u�6Y���:Q��Tp�"��]��Z��_�5�S0p�x��]ܬ/w�(�3+�� f�U�W1�c�Zi�J#l�[3K�}�Cn�E-��@u�d-�PI�c7	�WY�j�B��=���	|���f�R�9Q֭k�[��Ŏ)�]a�J�4�WL���ld�[��OH��$fJ��;ƌ��5�VP,[��{�ܷ��jΥӨ{-����M���5���"�͢1E�������*ōHШ�DAjTF(�Q���X�EE��Q��DE��Re�����,m�(��UG6�-�QֵAEF%l��ZV+mPU�QTUQkQH�K-�b�P��D�[h�
�lQQ�Kh������Q����*6�+b��16*�Z�����`a�*���VA��*UE��fёX�J�UUDQcj�F+"��F"֪V�lm �iE+V%�[��(ԬR�Tϭ�_.��|�t�V���q�
s�+q�C��dΧwk�%��:ثTo�
s��������KMĠ�wx�H�Tۓ��Hw��W��yc>t�k*��9�¸b.�mlR����U��1m��C�/"��ܾ���L�,��Ӟ�zOtpO>s�ks��DB�*�x����R�i5��ߦ��>�6����8b�yᰰٞ��]3�toLMX�t�Y)p^�(H����k�`W�]����Ƞ�'|���b�$^S��1��9�ǜvtk�=�];��Jt�s��	U:�QB^UyV/Zxf��"]T\�
��l���ѿ���1��R��)�0�oͻT�����}@�BX(���k�
��Kzy�#���H���ix�`���īs�F��=�&�����h�㜓��!�j��WR�����)!�Z=5r��o7��^���K��(�U��.�����<72�Kw�V'ySS�����d�,�6l�X넊^C[%�Y�r�*Q0p�τ�8Jo���e�|�hīm`�\&�ޚ�M@.�3�k*�2��GCU`��T-�*�x�/��(��[z7q����g����y�<#tz���R����@�9��ec����ڎ7O3�7\+��x��`��'*���PSq��w�@f2D��ř�����EH<.�������T��n=�T�u�x�v�IWt��:,}�����s�q�v���s/���Y����qƌe��<R��q]z�S:5q�It�X�Ѻa�����)�m�������y�;��AG���&P^0`�Iq��|r퐚�v�j��9����2o�S�Ez��R�mXP��|���"ϵif�M^e\�O.њ��8n���ಧ��X�W+
�;-/�C��%����cr�B75��ő@��<����>�������COO��Z��+5{�f�6o҉V��E#@w~�t�֋�7�=�{/�XxJ/6��{���=�oÕu	��1�W�=��Of��ۋ=��h�&�p�d���c �k�5�"�]���/N|�ؔˠ��� 4t,���bb}6��`y깼Ǽ�f���[{�sK�=j�߳:sѷ��e\V/씸_��%���A��?��{��T���3���)s���|.���ړ3�U9P��V>�r��{���ቦKP�;=S�	�z��=}��!c�|-j���E�w�8�`ٔ ��5�rw[C=+�uŮ%��[}��{\�^S�V�®k�R3�&�|�Π%t��9>Tj�>r�^Z�~ϖ�ټ�����wp�x9Of��Z]�͍c���1՜��%n'YR]l��Z�S��i�YVU�Eæ�h	�U�3f�8ͨ4�C�o �Iwn��8�a�3���>����l>��1�=A0g���t%-pIcGLm)��ҝ�,%͎�K��y/'���}���ע"�5Wgj��+�;�O��K��:���Ӏ��\���x�����A�x��uص.;r���v��T7�s*�>0/�R�0��l����7�'��9f>����0W��-i�"��أE1��fD�*�@��G����=�{%����|�?M�Lkx>K�>��C��������
�P�T<��}ʡ�ld}ն�;�J9�I0V��Χ)J�&*����o��G�¥VL�ͧ,��ض�zX*���:8g�Չ>���q�E|�0��oO`	m���N�����n�<a7���Sw0P�ۧ́~�g��44�]$'�åN*ͼ�z�F��!k�=3W�m���J��+��tn���ڳe�*T#�_�1^[���+5�$o8�>}�9��w.�S@��9��A�Z%V���LJʯ-u��j�_��O�p��^F����ª9��2e5V�(m��d��P3�5���� �\_E[IE���u�j%}��GSxe�]�'
uE��b=ʸ:yX����,J������
;�,N��E�G
\:�tD��	��Ǘy��` ��*N��|y$�Y�/;�S#՜�*3>#)P}����\j����,nȩ���zX�������\P�{{�yhr���V��M:�S��k�V(���2n���Y1������ٞ;�#L�:����u,(yJ\��k��WK�Pp#�����ϒ(ۖ;�7���Jno�}�c�qb\���{�g����`�T]ԶjLz�!Z(j�sC�>i�fo6�~��O+9���xЌ)�nUB�CR߽���WP���pe��_^EӲ~Ôg���o���?�NnH�{W��{��4u�w�o�h"R�R��(z�;�h�go���oV�n��tbcI�ˆe���X)�]��)54��Z �����-�Tg�[��9���}���n�C-v�7�sשg�V�C�_�j�����L|���ԡ(��ә����>�^���*��DF�<P�[�ڣ����.PO)q��v&���ͬ�N�,��,lW~��>�p��Yc!�<N�-����v/N�%���A��ɱ�Dm��t&s ��v��n+���e����u��*Xj7���7\Î
�4*m]��с7N�� �kS4d�	4;�Z�w]��M�k-�δiC.�FڣZle��.ٝq+���O�s6����ǻ /�Q��E��b}K0J[ar�9 
�}^"�k�D��i����2�0�jx�P��l6�����ݡ�k�޾��g��|�������J�6���F��M�a�=WM;�w�^�:��hL��c{���ڎ��[W�����"����IŤףw�Z�N��5��Ȟ/o."��\A�� ������\-�x�(u�����fs�*W�i���V��m�zE�Hh�s��M���V�d��F�����>���p?d2�V�0�ƫ��hy	{==7/80Ƴ�S�g�mW�n��v��Tx4�D��M`nz�huP��|��n�A稫s=&b��A�ؼ�~�7�{���\{��g�ا�pM�S�>pe_ԗ}����]�4k��[^�v�~0N�F��0oK�aچ�����h��[]b����W�*�L3}�NY/|R�#�_���*%��d��Xቧ�J����=�W��Ѣ�ếi�{�=�7}-�EO���UO-J���|�,X��kOOk�"_�ݏ�e��9�x���xvo��x�y�]a懞"�v��I��Ɯ�u�zVnu$p+�V���N�������*�s��놝�ĩ���qf�EW;mG.�'���c36"�8ț�;w�M= b Y��u;F��r�Iigm������]�]4NGk^�f#�Ұ��X�������=�D�-W���򸡿�Vi�Q}���W�����]�'/"�K]~�+�1�s��*0}��/] )Ch;D�-�2�lǜ'��HE,���Zr�;Ǝ���XV��Ԯ�a��p*�.f �]/�MQf����+��ٯ]��f�p�Ej*�]WZ����hz��*�P�'Wl`�3�,�6��B�o\磻,Qb�n�A�g�3k��\���2�U�/��������j&�M�j��6�����Jq�KE�\~+��>���T0y��� Rr^��r��о�v0����8�*���yA�|��{|���K������=D���G%�]�y���:���n��Xβ
������y}vӽ�^�dׅ?�^gPBm�'�=g�f�g׋��(a��+=��P����J%Z�l��د�.�C�U�7et�fEt��;�6p���2+�2�ל�
�2	��C�u�Y�r�� Z��o۸R]37<&��9.|6�Q�vD9�¹K\y���k[���#Uv�R���l����:�f�� �[�^� ˙3��#������8 }։�Ff-�T�{ز�J��P_Գ8���Ǡ,ɤ�ݸ��;�����u��YOH������$]�ʉ��cy�����$�.�-�ϼ`�`�,IE>�^ߢy�'��u����wk7n2�v.�/a���H�7ex��:�����/<�����V����Hg����ZͻG/6sJ���R�`ߡ�ghg������]cL�1z^õ&��2�$��fL�wBo��o�|������\�|`<u���?W1��#�S�Ǭ
wı�y��=9Wn�^�FxM��N�چ9Na)���}QKaMf�7:����=p �ಌ�\8�UԔ׿/X,f/N�goE�^���\boo����,�\^¦��!�����M����Ya����Xԏ�������vX����,E�lZ�WS�2�(e�I�d��� ��{h��a�ֻ}5���??՟?V������	�m_��Ҙ���p�Zr� EGk&��u�bȻ��-=U&��J\K�쳗�>)�|e]��`*��P	����\+λ�i?vZAЂ <x�.���	x���Ӊ�U��O
w>2ɥ�������QR������qз��]\5Xμ�P:_M�D��1����!c'�g�t��Ou���+��(`��EgvM^�o5�ܽ��MS0T|�>3n��-�3i1�u�F�ua�=#�kw��Gܐ�qV���Ǯ�iXܭ��{]wq��Tuk,�}���Fʆ�ډ`Jok��^@�[{���vͮ{�d���J��\���G��
Qi��d���v�/"���;9J�{�Jn
�2K^�c���`z��CvE�dX�N+F�N�_C���xNK��x[+�?ZMû�]�ә�{�d�M�L�^��Z;)Of��?l'�Ƞ��H�O�*fKx
�f�4|�ޗpx^�FQ�چ��	> �*�Lm�e�Y��}�N�<<7)[�������-��-jv~�vܾ���&!9�PC�/E)޸<���ja�b��b�e�ْ^'gG��y>Vp��x���3b��`�k�T�9r[�P��Bm��;���{�S�kwOJ�#N�ӒV�&]F���x���P�g�C����� .��8��:R��2}�<5�\p=;)�x]^�Хtc���t��!:%:KFK�)���0�m���:5ú/il�|hG���p�J�������YR��ԥGf!}���d�����oc�b�>=a׭KCؽ}掱��k>����><�-����R�[n�/^��f=�'sK�O�.���9*]�c2wf�HV
3��cxQ0����5���Rj��oۄ�Dy���� ����Ͳ�!�6�Y�&&��Tq5q�X*U���:�u�pd�>�$�}5A\��pgY��+��a��t�g<Ҳ��!�#�x��;Z�� ���C�븠���R<��2�_�j�i�L����{��=E�[��^=�����/ʐ�NC�mǧ����#@�u����;oZ�˛&+$z �I��Pؔ�g��I���u\a��W��돩b߽)�[Rw����K�����x���iW��J��U��f_�d�x#& !'���ԬS���Y����D#�죾���u��Z.�e���O|6��D���*������u8"�$R�';y�А�Q���/�M��t]dY{U�^8 ��k�s�<����h[�W7����7s�޵*4AU;F!t�#�K��
�+���LF����y<6�7_;^vV��h��p�GleG�=^�[�Z՘G�[|g"��;�T*�ob��Yg�}:`����p��|2�;�R�������T��y�e���R�� �6���ݗwk����qtT��
��_�+A8/����(�y�&&�Mx�j��R�7�ӕq�j�<{ �96�z�������t7X�u�$'S�\�Q���ɋFF�v9,�r�G]�Ȱ q�j��6�`�(��e�:7X<�,���':N�ohWJ��Ezz��1.��7�Xl�N��U�b��S��Ϝ\������ɋ�@v�LX,?Q���U��o�,M�
b:S^��E��چ
b��Ӻ��d˱�����k��vL��U]�1d�c>Q2^yV/Zxfκ"_ӞT����{ڥ@�F�~OS����Gي��ʥK�.I��I��L[33�L`��Z�=��șw��Y�ώ��WDNo�J����ͣ8'�*w�B�ի�l'�����O����r�4��{F�jM�H��I��|T���X��P¨dd�t��>J����瑒�6,��|����{b�x2T5���;�^YW.f ��p������sBA��s,u��[��u�3Z1��4�ŏ�\M��AO*��$G�W5RPL�yu�dβ����ޚ�J��\� Y��@({ꇁT�VTϙU�$b\չ~��������r��O�C~7�����^O���`���̢�S�%>�6�/��̱�F�װ��x=�"p��r�[b�"�R����A�Ū�dJ�����i�2Y�4[֑�R����Ӿ�v���֩��b�.M~1�4*^8γ�-��a-����B�^Y�g���k��#{r�6��j��Q�o~If�:��1��fpG�)�iXd�iL�	r#�`�T����̈́��+��rMM�����9fK��\�ċ�����0��a��s��,)��դ	�x<G�v����Ku��nkL�gs_@��C�	�ۮ���;H�t�>(��Q�u�b�yn�H��Z@����v���K$�.��D;U��0��s�����b<�ʝr��9p_N��y�T;��u�2�3F��]�k46��G2��e<��^�t��$��q��V�%³���h�OQu˩�MkQ�Q��v�F��b��cqқsax�19�E��1�&q���祾�չ<�^NВ��:M���\"v��HeCS Z���)C-���N"^-,�t&���>,�u`�)�'ZY��F:�8+�a��(R�j�p���Tyw��cL�0L�n�-cxVB`����(�\�+yT��7���n�� �{^���q��,������4�ɕ�L@7��T�z���˧���|M&p��z��e,�j�b)a ����iw���f�5R�7��c5���̧ɭ�{4�I
6��=�e̥��wy5[42���Ǒ5��TczV�7����8X�"���c�d ̸�Q�#tU�(��.S69����hcܭp�)Ģ���<�����:�w1[�.��(��f���f�"��ʬ�B�4l�QB4�;�Pf��Ih�p�ۤ�f�����e���m�oqË0&c˼�Tڻ�!�E��7�@eȶ/��X6��;�F�Br�>';,�G��2�1X��z����>��]��^5�%�Sȯ�\q�;v*��t�P�-�iaA��L��.��.
j��Q�{��׻�J��Kv�R�\�	l9wg��*��:��5�I)^qƸ�Ԯ��b�2:�����<a�3)��3��tfhs�Bh=yH+�Ti��7?eI��s�������0PN�_7ݦ��Ñ\��Ѓ�Y�\�䭺Ũ�꼸�g�_Q=Kqsȷ[�M��`�<�T�&݆u����u��=��f�b�F'B������u�#Uh� �V��c1�k>%�����h؆��ٳ�w����,�wi�X�����T��I[u��5#��l��Q�P���T��(���n�S�NE�@4j���íw
�(��Q����Ғ�������,��]��@�VV����٭]��9ۭ)�E,M�Ӌ�:5Y,[Q�
(">RTQDF�"���1|��h��b��1l�&�Y`�*(�TE�T�kU���0����Ŭ�QTT
,T��mkD�[)jF���Ъ�j��R�(�eK�c�IR-B�Ҭ������chW6�AE�0bD*%F�D�ڥ��+ilIidJX+D�e�j4*�Z�V�h�Q�08�V�Q�
UJ��l�� ���F&m�UX��J�ԭ!Y+T������Ԫ���B����TJ8j�	ZT��}��}��lM`uܤ$\ͦ@L���ݥ����L��1R������^�MlG��-}]��r���7��KC%:�~�6�� ����q"|�K�п(6�{喥֊,�q�2�>����Xk�uf[�����^��ppcI�F@���A_w\!�o�=�K/w�Y+��������"�~��qNf/xD�?Uh3�E��fg�Z�vǾY�6%o�U���uՋa�k!_�N�;/:�>5硈5Z�����T��9j�}�^׮��r��6����$�#����zsЛ�WlX��.�5(^�@��l�OG�k�c9�*y�wZ�${�;cμD��tn�l�WbEZ�Cp�S���:��8�V�c�>z:U-��\ѹ$���ܐ"�|��K���֙%n��0s�\X��B���{�X�x^r����ؠ��#G�óϳ;�>^yx��D����[�F��ut!?E^*���t	���+!�}��!^���7vlG+T��2"~ߤ�f���
<6��BP��'l���ڴo��a��nn]�����^ؘK�7��h��A�`I^�^Ϗ8h��C�d�2�w��	�x﭅�I�i��Qm-��k���;azW�¯f�]���8��ӎ�h A���1+�DO�_;���]P�3햠��ט�9wy:uhX�m3Q�|�����m�m��>M�^��b�����J�o�=��U��\�O��+��ϯ1�<����s*��K�@�IL�Bd)kD�w/���9�!T��������F3d���SΤ��-�e'1�	~j����݆G��ɐ@x�����C��"��C�yˆ̉�Rti���{�S|��Lhyj��z������>�����:�&1:m�V�.�0x�̧���6&�Um�G����?W~WP߄ I��m'N���U�T��N�*�L���geM��/�(=����9�=$�"�:��s�i���]�l�ޛ�7��GU��0\4���=��L#�T<`ͦxXB��z,IΉ�wR�#�Ex#)cjJ�5e����z{�w�G�0��|lnS�i� ����_K�Y�73��N�����"�i3�a�V%��o�'�=�}���K�E��(%g�� ��Z'�T���Oݞ�>��#�9,��?�A'*>ʮ��_v�Γ"�5#Ӣ���Pû�V��
����ko�<!�e�6�L9���,N;�8t���W/�*�R(*�Z���0J�^'���H�ٗY�W�1�</MK�8d)�hյ�Q���j!�Q;Ǎu��ōg���R-�5���si�VR��&_`�YJ\�:���H�;,H���
�)������6q�ʓ�z�X��z�킘��y�q�����(L�.W�r��V��3�*�n�Q���z�p*��%cPl,A���*����0�e�X��j[�:Ǧ'����>K�Η�$S� ���S�W��dO����Q/�ZYT4Oez��n�*o���rǃ.�-��JE�(���Q���֌}����!��D8Vc�u�;'U�0f�C}¼����X�i�a�\��ico���Uօmcc6�F��^�������p����`O�_-BN��fis�痂����SW���2ei�ƕ��'/� ��z*�1�����R���ʐ�:�O	�Õ`5�����~$�/j�;�nם]����S?-�Z|TfR�8|ջ��)0a��<'U%�����g��x�\ܺ�N����������P�*踶���-�bt���ˡ���Q_���N:뾪X%�
�Za��]�Q5c�!|;�0��ԧ%jɩ�c�.���Ҳ*�+т>�p����B�؍N�ɡoWb��zT�%7&�tߌv�A��d�%�͑�%�hVf`e��7r�d1a�H���;�����]byٿNW#������Ru۵�Ty0nT��ݫ�t�͊�>�̜��Ū���68��0��%�侦��X]ʾW��;3`�L�U�����o�3���5��[��Rĭ�IU�B�@7��~#1v�ȟٴρ��P�,�)Π���?bS��o�ք��:��Az`{Ԟ�:�=�>��̕uȮ33��I(�)�c*�r��Լ��|ݘ��<\�<"������V��OY���5^:�n�y�<h{�V��kXw-��emp㠆{�@FE�߯��Kӑq������g��^��y�P���>���}-��h]��T�X�_��+�&��53�S�*�̀6�Ǿ�
�ؾ�F+.=��+eYY��nR��𼉋ș/<�˳;��R����Ʋ< W���^l�9[2�M���ʖPx���KV	�e'���x1J�.��׵r�z"�ƺ�b,��4�sM�ڽ�A%z�����1���G��#��;e�oD^S��ze:;��U��닪��Iľ�_c��|��ù%�Y��e�^�@R��@�^�~�U�\��S�&�J�r�h�x�L��}��5e�F]����suy.[Pq=���X��yt����IƉ�x:L�+<V6�QՋ5������ޕ�܁&�kg+���\@'���ƥ'�5z�=3����4�te7r�Y�v5�����_(�9�o^ً�C�eCYT�fv��U�EF <'Q�qx�xu��}��%�����=�f�T���Z��g\��mڂ�K����Ue[���ة����g����{��6�q�S�yD]OpKDȳҨ���b1t��{C�Z���խe�="�XA��MӤ�������J]_U����p��h(���L�����X�W��h���B. U�K1��T�оPmR=�J�4����	`��w��]v��J-�����D��놈���ƅ��H��78mx˫�]{U��O˛b���VC7�y�V4��\5��,,��9j�����6o�J��3�V��ߧ�[�Ozv2�����Npܳ�/��Y++);��C�wXȯ�k����-��M?�W�1=ȱ�S�-{/�q���RY�v{8nm߅�ȸ_��w� =��l��>
�S'sq`� ��<γm�슞W[^����esY�t�0�����^1xx�Y�������TYu�̭���=+�R�٭��]�t;q-�z?^����;q}���ܼ�qR��|p�2�+�b'�=h�r����2����,�.�YU�hZ"�M]D�E]d��W�uQ�P�q
.����{u���N��.|w+t"��S� �fm�V�?�����|U�Oz��j��y����@3��Q^���nj��vug{�F؞����i���W+�k�pu�׍!(?��gQ����ceCzܵ�=(%�[�^q����;'%Ҟ�2����0l�u��?�s��T�7��q׳N_ec��:��-\����:#ka�5���o���������L	^(��8�� ��u�KS<��);c=D����L����y���Gz�\4�_H�
�j7�	 ˦Kk�onp�f_s��O�ta�p�b�Ǭ�h��%�l[A�T�����ɃO-�vT�g�����u�^J�����^KjW��^7`�ƃZ���fǞ�OQn�W��.�?�q����Ɵ�h���X�A(�Q��v8��>����ï�.��e�]{Tn�P�Ծ�o�<0K��A�4>��S`l5z�%啡�	N����8�tz�䘐z�#Kg�
�P���*�$Oƕ�B�[F���B[k+k���R�I�[v滞�Y���[�W��BU�*��HS�	�B~�A�
�U����L�"�ғ�����q�Vyz�r�lZ��N���Kշ�=//�� AQ͇��c��|.��T�"��8�\��
�ӥ:V��gQ��%8�&��CY��7rL�]���yB�xg��9(;ubP���*�n�"�vEB��Ըذ�'�g�;�A���+ﮌ
��,�_ٌ1���5e�L�z���C���OsDg�!���=���rb�v���$���R���U�r=7�]�z����&/zJ���vd�wuɖ����lzW'���^�\փ�J��.���:��ί���Ce[˔V_���{��,t�lBׅ`�H�1�:_q���J�{��qQڳZ�.�G�t�^?G��c���P�|�����劇�����Iw]�6�N�Xg�;��5�b�}�����Rۛ���2�Ixc�
��O��Щ|�p닟R�3��>�|���I�Ȕ̽˽p��������ĩt����[&�a�c�ϭv�I}�}�	�{��Z��؆��M;r,���d��	]��,J�KG�>f|�S'�|<��{Ϯj�K�e^ھ�z�氉���W�����!��P��?>ل�X$^j���̿Cۋ��E:t�7M=θ�ѧoD7�d�y�F�9��p4[����t�Q�ٻ��8��^t�łM8��J�0<Y�ȣ�٫�J@���U�SZ��b4!Y�f��(V'��M&�ywtT��[د�!���-MZ2���R�U�QZ}fw2kl������xϽ��	O��*\�^t�zr*mY��r_9�p�]m�t�m����τ��U��L�"�%7���h|�N����V< �kݦ����
N�kY)�W/�y�X�Hl@�z
�Q�=�)\aD:9��6��y7ze��E20�j�i�^��ˆ*�D��z�����]��_l�Ƚș��y�mI-i҉�S�!	��Ax<�K��X͜*�X�̱��,u�W����
z�K���#�Qƞ�R�����gJ���'6��_/��aQ�?�i�ן{�u�QZ�w��9���-�T�pɕ���0q����kZ`Z�g����Ɖ!c>a����X}åu/,.�T��]�&�y�abܰW�_��9$���cB�g!�MX5��sګe�S���qQ������~0�
�zo��s#�*���ҝ�����ѥ��s]Gp�r����Ud���"���&��S�f�;��ٰ[��ڷk٠�2A���iT~�dui{c{�:���O,�M�6�w%g�p@�i7;ynZ'˔Y��>L�a�~���/x�@�cƇ���a�y��FM����6�[�Q`��������G�dעĖ�Dy K�eZ)=�;�u!׼����u��䘪�ګν3�gq���X�p��.[%�Ƭ0�xfκg��~�Y��=�2�K�F�WJ�=<xݧ���PD!�P���^ՠ�˗��K�,N�&0R�z�sXG�G��ҽ�D��[�X#>E�q\��V9�_x䵕i{�o�k�=*�|a���Y�	^?<u�-����c�Lׄ�U����
$TP�
�nzEpJ^}���/[��ޘ�r�U�x��Vf��ɵp�U6�;��^Yr�7F  ��1é�����5��������['ݏ(���
�CG�&����*��M�H��ʍN*����4+�Vc��k#�Ipc�`��E:^Q�T�Y����������ў��f�:����C]KEpn�^����\�*��8ʇ��Ee|�a�R��nOH�v}G0��UgQHUڨ.��t���@[�)�T�-,1��c��aO }�9�y�\}A�Xjd(��C�z��Ex	�h�����0��L7չN��WA��k9��N���gT�os��N=@��Kc��Mm��(�cu)$\
�㼳z���A؀�g(d�J��2��F=7W�:�=�&�k`���j�'��v� $��_2x�^�������LT��8�j�=��3f�ˎ>gv���\++~>Po�i��9j����|s��,D�?R#���|���R���oE4�#� ���c1�C�b_����s*�L��ݔ�0:��Ԩ�{�)�?{�S�#��/zY�^;r�/���^��f�~�Pw^:��O�#+2��/X���Mڼ5�.7-{�t�0���症J���sM1�m��EU����z�P:�S����)�c>qFx�n����9�X�,aq
6��ھ��t{[���|�=����n{8��ͨ0c�&��b�vu���7�(@�F�'u�0}��V�=p�۝��]9q0_ދa�,9�GҤ�f�襳S9>)�<х����|FY�ٍuV��V[��ړ�&���}@/=��{"�55��H�'���T=evPw'��dk��M��ղC�bOQ�typ�E�@qb��m�t�	�h튮��`dy����.��ڷ���D�
s�O�7Խ���t���4���&mA)����M��!�Y�'B��P�j��\�N��.��� �W����8ҝ�'������7zm��e�wV�\�ݑYR�8�e�Љ�N���)���Y��5���ӭ�#:�%��A"�^����es2�ˎ�o���t�y�2o]ګQ�W�L��V]�K`�hoJ�p-�-�
��c����=L�M��6��0."Yz�V��mKQ�ά:<��(=d�Û��n:˫�׸���MS3�j0>YG@3^�_����]=�u��e['�+���kf�Z��Os}M���}4��g%ai���Kh��1�j��sYSø�4����1;3B�B��NfmN�.�c�EQ�ҩVJZ]�:Eۣ�b��ѯ����w��
y��N�˔N�,�.Ә��L��}�7q�䩞�|3n�Wm)��������Yz�6���)���z֑���P@�;�Gu��X���u\��e�e�O4h�f�T�m�q��M��v&ݻ�l�|b��-��{���Fr��l������m�`�2NM�A��є�OMޭ����U��K.����ZE���wj�u��;�02��u�,so���)�qz��f`s9	��#]%;�,��1���~�|��X���{�۱���k�/�ŕ�݂�j+�(�z�f<3^��J�����pd׬e�����v̬�剻I��N�+u����e�J�vL�igGq^u칣33tҀQm�#���
��:u�Ax��%R��y�8	Â��C�3���/|�_c�-^��<{+9fa�ݛ胁�"���Zy.�$�F���I�kc��ü��@���l��hS(w*
�?L��r�/Q�`�ֆjk��w�tt�Z�Z�u78�K�q������H;i�V8�.��d��4�s (���>"�G���r[M	��/^rw-���Ti8Fu�a�%o�8�r���k�=�ܱr��ɝ��K*԰��ؽ�329��__EϤ��t�]�B�n���6�4v�r�,qm+���`�Zj�Xz����A}�Ȝ�=&Њ�GTcz�uc͵`��NF2kJ-	X��<v�����FV�X�y��ˡ�^;�Y����6��n��B�;g�n��(�^��f�wU���K.��c��򊮏D%>�'\��=�<Rw�M�v�����ݨ�4��n�U�����|� \j���=�KRC��em�տYru�鉏��h[�8AZC����,m97��U��\�`U��{;6#��l�3i�u�k�pnbH�VBuI5B�mwP[��S2�!�_B��N��'���Hk��VH�� ���Y"�q;;u"�8sG;�8Cl	��Z�c�,\�.��I}����J���I�[X�a9Â]���DNaJeuvI��Wd�Ց��e1e���5=坍çG׻���2(�R��X��*�Ŗ�E�-����Ա�ѩR�*�[m�����*V[QF�H�T-Z�R�ҕ.�����-D�Eݦ��Z�J�XVP�R�E�AۜQp���abQJZ0�YZ�J+V�R��X�TZQ�j�J�iikZ��l�D�\b�R�e��b�5AkD+VZ��[F���bŋYTV�����X�Y�QT���ʂ��D��5*�Q�����+[ZKim(-eJ�VTj�
����r�5�Tb(�EF�#iEb0bĶ���F"1eT��5���AED[D�T�T-*2*��V(��J��" �J��F�*P� 
�@}wC�dce^��0�}F�N�:k#-�`O���
����ˣ<c�kA�C��������=�]��b��dd�ჯ+39.��я�P�8����98*~��P���Xr�����_�J���m�u�fe��z�TZJ��=B4�P���U�Fb���Ӊ��W����e��/ Oc���~��;�^�K���:r�*�T��1`ߣ��s(�T� �K ��ˏ��[�{���ĉ��W9�kb�G���������E�18����dx�� Bu�*��ؤ��
|f
�b���]�p��p6D�r�����&���[�˖ڑ��Iy[�nl�El��3�"�6���4�KG��o�	r?	X|=N�`��Z`�p�a{;��m\��3�z��eH^r�qA�u��Ad�h��&Eҧ#�c��������4��CK���V���l�zX�wJqh;)J��_fU�E
�SFn�/'�e�.�~���4���q+�T����7�d;�[��7~��P\oh�V��ٺmi����dI�_Q�5�~~I��C� �x�j;�>iW�VF�L�g�^mZ�����~!���Q�1��z��W�V�NZ�(�/a��ݚ�zi]�{lV���r䷌�{�lԽ�"ݮ�b[�.�Y���(T3܅�[�Q�4��wwV��n�c)}9'N� �g`���J�M��s[P�iY�K��9EN��/���}9�R��.�U�]�=�(�Wx���X-�d��o�K�6�<:�_�Ic��O��:��2��z��0�9�4tka�?l8��q�ɳ�Fw�J�^�4���$z)W]GW�.��ǉ����pg�-���X����x���N��=��s�奲�����7�d�1Q���j�]_�GI��_�-xeC��{���^���[6g��vzz�7q\P���}�T|�"�Nc�Q�6�Vs���nF�����l���-�d>'%��U�`�Z������m;X�g��M�f<��x��\�0�y'��S���Hl@�ށ���G�܅x#�'�{=�M��gK�!�{$e	���Z����Z����q��]H�� ��]�J�J�+N��������7��$]�|V��tK������fj�d�~G�L����f�x;�����Y�K>�UI��x��)|��aQ�Z�'�x{޵�����it�X�d��:D����<㽧|@CV�@�D���w����X<U��1*u0�Ûj�Z����EQ늆j��-�S�0e��R�C6�;$S�o9�x3e�^s8U��5��U)nv���7�sR����B%N�b��M<'�}�{j�����A��kN����ߦ ���S�������� �\˞�פ@��o���k�W���`�傞��6�;�}�5z"厼��G{bk$��XKl�5���N�l�#>�Ц�ɿ_�6wt���򻿇��JƷ�O:V&�zq��*�A{�iEcؓ/%.K%�\�jc\)��I��qt�꺱�v�	�v'����A�(Jc,a�9x=Z�Y�2^}�X��iឹݾ�PB�C�4]9�^E
}�l�%�B!�P�
����{V����������A�~�'up�B�q�d�ٽ��Y�R�X�h����#�z���^)���%}(UԻz��O�w�H��;������gI�.�X0�<=O�C�/�O���t��ù%�YV���B�
���C6�Vף�&w{�����B��Z&?8h������D0wu�����vh_�8P�bC6�T��E��3��^I����,]B��c��T�Y�8ǒ|�č�(P���#���(f����RFw������wN�޲$��ޙ�f=}mr<.��Y�e�:�B�A�Y�Zz����]�o������븳�\�i�T�c�h��;��N�u|�]�3�(�����ƒ5(n�uٛ�n��]X��q)x�v�u�u�wx̗�p�^��A��g�����ނ)�Qb�kY�#,zW������d	���y=Q��Ф��НB�NuD����!�S�-˗��|o���g�r+w+bg��tg5��1�ʡ$?�)j�5A}�TσB�A���e�Gظ{vE��ŷ������Kh�ZPuu���\_5�Ϟ���u�T{�WA���ǻ�cś����8c������wLU��J/��X�P�~��!�b	Y��~��l��D�Y�L��^���(r0z�RӮ�Mぇ�C��4��wY�P�,g��~����i���')��JMy��q,eNZ�P��( ����N[U&^>�����1�y|��^S;�����U����d7�O-��x�s���a�K�=��iU�v]9{��Վ��8M����S��E���u�A9����m�n����7wȔJ����M@�<#j��12��b���gz&�B�lmj�WC�ݙ�ݭ[#U9���-ӈ��]���z�ȭĸe-��y^���-^2�ɏ`"uCi������c	ଝ��[�{��`�g.�7<g���_�����+��ֺ�23J��PR&K�<�Z���}5<��܀�Ʒ��Q6��p��[�JU��2���З����>}wS)\�K�C{9��9�}�S+��6��a��c������G��a���N�h��� 3�u�����l{>z�+�&�	؈�SUZ2��U;l{W��}e͛"��c��l.��h��/���3/���2*y2�9�0����H�{��~�e�P�O��AQ'n?8*V��
h=5��	�mM��ȕ0��i���9�K��|#7�9mAF��j��:WO�\L����g�o�:]"Ї��;p�m?r�)}�<1<`n�Pm� .��@�:*�z#�U֖�@�XS<�[�^���\��傰Qg+F]t�t�j^��Џ�]xU��xU�w��v�Ϻ�f/?s#}���[�=N��B��lCcQ����B�󔐷�F�cVb��s0]:��"��2J���O�U�[o:m�ˇ �P,:D���~��Q�M�V���E[Vdޔ�u!�Vm����l�迢�5\σzt��zlc����`�Z �]�K�ThQUf�Y@��p��b�6�WrY�t�䇹"��K�˶x�M��of���=����9~$/�A:d�G;:mGO�+ǽ�jNř]y��Z�ɣ贙:G��Y��m���ۮ�����B��sI\�ft֥ڙ�M���f��o�Kw�Gb��s}P���{�+����ZCk #Q_\��+m:A�˳ɳ��S7���}�C��|*}\�����N��7��Aȶ��N��JbU#l߃]}2�秽~"��#��{��vׁ�>�Q'��aʹ�LN�V��F񍮎cv��tu��0k�>�ے��d�Տ����8�u�
__R��֙>�;���53����/��u��!Ǭv��6C,z�����D𼨐��hu��ƯK"ڜK�9�]s������	��Rr�d.�y1�1�Ǯ��MK��R���1l`����fѦ;N�ܞ��)%}�֒#e>R+��1�}tzOKƯ�hC~��SHC�@�)lx��c���M��)��_u4�מy4�:}�ʋA\���*9AKgʝ��`�kw�p��#>�&qb�q��{&��o�k���U
���z&S��r�DX����aUջ`�EHS����h�1�4:�'�b����ލ�+P5�n����;P�Vب�&6����l�ZhWT(C7��;��3�U����t�y��{5f�Ō��;�� ��Bڤ�i�W{w�`~��V #a[�Ԯ�7�$���pZ�_kn�>̛.f���*G7܁Y�$���R��� 8��s*�ddl�UΗnŻ��&�j
����".�-"�V�f��4F��ƍ9�kL���j�pz��6RZM����f.:2;�3h��J��u�G���_�������G2�aZt�]���`�a��:��>67*Z�E(��H�â�m�S[�d�̏�=J�P��|�:Q7U D/��`��~,���8֌��ٽ� �����n�Z�R���8�`���"�73��Tan��%�o��NmC�)Y}B����?��</��,��OX�O+�{S����aYSXç�+-^�=+�J5 �^Z7�T����a�������R�(F0��?�z��\b�����{���7Մ>���/�쀵C��ppy55��D�f�X�/-�.����u��C�)T�~&U
|x�v��ۓ����͝)~���1����蹱�w�L3�>pd��1u���
�m�`ס�{pm��ƹz�B�-c}O|<Zm����TU�[u��a�~peZ\0?��pu<����;r����:[J������%e�Kbb\�
}���i�p��󺾡u�>>�t�`T�|bx<�2��8>WsTB�ו��,���{�蚖��PT�2��RC��'��Ts�Y�(�� â��`��[���ihe��i�[�rgP��s�e��$n�2y�Ew��Xj,l��n�hNUb�x�b)�I3{�c�J�S�wԢB�l�}K(���N��4��\R=}�N�eL���t�ԥ�)���u	_x_jv��V�r��{흼�wDڳ*%��p���}��O�Q~j��%�Si
�����1���rՙKkf�RH�3��	Ṃ]A�r�ﭭ�*�7w��iz͸�*��Y�j~�$2�����~(�D3�Ԩ7Gmq�)Kc;W����Ur�h�[�9��J�j�U�,���.��	m>*���E�)Wpg���3-p"�5���G���������z�hQ�?Zٹǥ��?�`;����$���mAW�%�t������f��a�9c��{�u-��s��lc3�(;�vA_���PW])j��@m?���G�����d�RP�g'k=0�˹G��O���5e7�L���G�6�zB�cՅWӖ���s!�s�?�Fx��ๅ빾YW��ڕ1Yi:�!�,t޹��l�U�PV����RϞ�9q�N˲V)<)~�Լw�f8t��f��X�����l^2�������ňĽJ�.���Z2*��=9L���콝�yfR�DҐ��Ǎi��}G�ނi|���J:R5����!�����$��kl�</�Ǘ�CƆg\+C�S�-y�k;*��Z(\%LX�;�=i�)��o0��C�3É���;�'_��2�}��Mwe�Ԭ����z����잼]�5�`�.�g����0˾��/>�����v���b�>�U�h9��g*mlۛ���0_u̷��ٹ�F�l����)��\3�G�՞sU���y�����s�\[
A����S�0�������O?�P�����]��~%�O��q@�?lǭ���2��d�j�<�u��l�h�u���ٽ�jB��*�_q��>U��?]�{}�2��SW�-�j��g.��CQ�m�g
���|8TS�G]w�z�_��ۢ�z�$�=Wh]�}���9���i	!�d�P�Z�%�O��=9�]*�pB�w�O���ݝi{9^���G�릠��!���8c�q��z]�;/����o�2<[)��i�O2I
ں�j.�p��/c���23oO_R������v��`�HW�TJ˱�+ya%fv�4���V�n����I[5˹�n�x�Ⓒ���&�b��R<�a�Dg)P�@֩����p��As�[xf6
��^�C:��k�{rv��Tp��� fA:�k����^{��i�)f�3��)u�bp�҅���3��J���V>
����:_�8W���`W�z�2�M���r�Ss@��|U5G��Py��
ɯ�Є{���ƺW�>;-��矝[��}�R�k�+ء�Yd�|�,��۳��wi�.�`83�*�A�qno�}��L��:�a{י�my��f����\���^O~�����Y�C�y�J�zK\:����ӏ���+ڟp��]yzg9�~}$���o�d_z�,
��f�w�Wy����^�;�����Ά�͜_����e�;��ٻW,f�Eaf�h~�l����^s�N���_\�/�A���9�$�2����������t�
����%h�n���hz��>��|���`��4��K��`�1h1�y�~����ŇyS=~���Ƿ�x���w�B���$���$��BH@�RB��!$ I?�B���IO脐�$��B��HIO�!$ I?�B��$�	%!$ I<IO����$��IO����$�HIO脐�$��$���$��b��L���[&`�� � ���fO� ĕ7ǏR͒laIT���"���*�̔�"��(�KV�)$%hh��H*�E %AJRIV���$�F��+kU3Jś2[f�6�B@��SjY��CU�m��ZRd�ڬ��*�Q�m���15mjK ��e$�$�r鑶�ڭ�-k�V+Fٚ����[6�&h)��[���j�D�m�M���4Q���FճR�mK55��ͭb�V��R�36kkN�K���P��   ���(Pг�p�h�6:��Nۦ�;���N�!m;wvt�[`Z+4��]7�(����F�ۦ�2�(ێݴ�M�ݗ;6�e��M�mVʛ5��V�   sޤ(��qF��.�ju]�iR�l��j�M
�]�Hm��0��(����[�³UM�l��JS[eθSTP��z�U�6�U;h�m���H�l�   =�(P�
((P�{�@(CB����(�B�P�B���
B�C�z��
 � ��=�x�B���
=�p�B�CK��{k���8�M(.S �]�JCn��Jک��R�[x  �A�ʡswb�ehR�n�+�:�@�ꛩ.����w ��Ws�ũM�ۦݗ��(X� r��黥�
��f�2�k�i�d�"՝ir�d�J���  ;�=tJ��a�P�t7A�B���tւֻ�٭�;��Eܭւ��Es]\�ST2FXSM�����mݔ��d-�ӻ%SZ�jY[lZ,٫Z�Q�ko  ���`1]�:۹ɭ�TݧEU�յ�8�mK��t:ź�ڹ������T�� ͶMں49����m]��)�eP2�	�l+F�� t��P�:�*j�m�k���F�� �j��;�5*�2&Vh�3f�3T�S.��ڨ���E-�pN��ZmZ�jն�kͳ[d5x  .=��*�&�sBƭq�"�����������q�G7@t�a��F��k:�(S�Ϋv���sr4el�#U�#mR6�o   \�S�]:�5��v��ZjWn��h5J-Q�A�%� &��ww3S5M��@��vs&���VƵ���YS�   ���:�ms�$8n��J�j�k���j�s���j�
]7t�-�m�[
ŭ��WN�涚�m����'�RT� S�0���   ��i��@ �JT�� ���4j�" @M$I�U)� B Wb��� �5M�I��(z%��SV��{�=V����@�$�s�s����H@�}!�����$��H@�8B���BC�:�������P�c%���n;���SK[ZL��`(���ͬUa,�1���mB�VV=�-
�%`�&$�f��
�����%�G��$�\�ʤ£i梲;̚��-R"��B��5�&:�q5+Fԓ ��!�n<2����Y$v���N����x�M�m��+ϡ��s7`�-�̦�3u �ph������Q�6YD�L���ch���U�����G]��M�i���	����� �9��Qn��RB�s�ZoV��f�B���e��K\�}�۾��X(�ԁ���oa:��4�Ͷ^1T�ZlY�MO�/�	�,ց�h�*��-~� u������ �Hܔ�&��[����n�l��7�%7P^A�*����Y��F��8e�r^�D�!��A`�b:�M��P�'+Y��Z�+��7�]�VJpc�)��T�����´�s4DJ���4�뭤ً0�uY�L5~]Q�L�e�/Yт��\P\��v�xM�5�DP��ď�q�Z�y��ve�2����]cx�VE�`��|��H��ߣ����VЖ���ff��}��q��n�`ֹOa9Pm��j�E5�(�1Z��̡�jr�0j�ړ����Pb�9Z�Tx�M��L��SSsi}QiE��WyCL��	���"�bn�[U�.�xN�`�2�ȑ����<�69%�9���.
�E��e֦֒��gF���+@�0b�X�ɗr���x3,�pY��8&�B�[��
ڗ�k���+�!zU�4;F�v㊀e�mw��S�і�eM����p���Și��*W��m-��mH]�̣��F����v��@�r褭�h.�ڼo�,��XVA�z@
1�r�_��c�*	�](W���b�ZtM�Y�����#T%�J˭I��m�M�Ϯ�=���S]��Ꚑ�i�W��[�Q���������sii׉Q
��-j�L�gȶ27hh{K-�B��zl��f�� �B�<KcY&VX��R��%�C��2�Rԝ�dW�!fIh�T�GiX�%X�V��6�-WmA6�m\TI5�lM�)j�Zj��ܵ%�f�d�-�ĶQOrP35���'T� ؒ�rP���j8)���8n�"3CEh[y�[X�A]��;ahV�ezúu�qB�X͹t�s�[J<��,^2@�ּ��ޜkb�T�A�e�H�ʌ���յ�n'���mD�â��x�P����z�hY�.so+e6�i�E�HK��ea��"9�,q�u���,���ɖ����̙�]�:ݙz��ݹ���sT
�^�)�;��â����zq��Yj��6��h:��d�ьYb;�MR0��nⵈZM��WX[I5�۵rZ(i95m:�$jVv6�4�-��eȯm]�7W�YQɸ�	ʸ��wRkŎ�����lc��{�Eݝ
�9�f�����\�m��\E���8By/wc�2��l[���+I�ۇY˛I�]�/o7n��m*eڵ� ��� Lތ�V"r��ˬI֑[+r�\R�h������#Ub�a`(Ф�b;mP��y�VQe7XpV��TKjf]�$�2�,!$�Nm�[�B�,�˥�&AGc�z͍k[��4S�z՚a���VSZW�E�FXj�h�kzkq=�i�v�T�pbt0Q��"����QllTTq���4�Stɯ+(Ҁ���L�j�e�5R`��M��H��K	�R#Qc���lV�P�����O�CV��wB��@ie1Ę��,LwCK˧3_��cy�u�rٚ�a�Omn*�Tݣ{����Agw({���W��?n�INͨ�{.1����6���N��g�/MޒDt�B��k)1vn��reY�T��k2V��U�)��s*X �c&f6(퓚��Ų��P:��+����P�T�Z�`ġV6�J�\#)@,��?��D���Q+&�;,l{���l���t�V�m�X5mPG�g�P� ƬjƻXi�Am���X���*ܩ�헐���eM��`!�1tWR��G)\ۘsS�5��jS۶F�Ml/v�J�I�*�lRX-�21La��Q���D�e++.��nV�[EJ^�m��%E�4�'�Wb��"ɽ�-�(�S�[i���wR��F��%Ǯ�k*���W+4^N��	���VE�ɶ ����S���%fe�r�tK���76G�r�Wr�:�.4��V��G�*�(V�v�3m]�ɵ�K1��B�n5���A��ofj��k����e�XÔюٛ�ejb��柬VM��h�20eb�McYaEW��JL'2ء�/n�_<JQ����MV��ڌ_фC����:uMQ�1G]S��,,^T�%ͽ��՛���;Uo%-7�O[v��޻�U%V0qO]"P�w���MțU�G���!��;�%�YhH�ʛD8��&�qcc4(�6F�y @Y{����Y�,��4�6m�Ì|�Q�,�����Ń�	J%�pKn�Ju!w�����˄،kOIaI��9z��-:�ha׎!��B�%�B��j�ܢ��}�ɀ8j��"��Wx��3oa�NU��Q�iT	\Zn�j�B��a�.�GP�v�d�CI�%��R�*T+J�r�@�(�b�qm�W+3nSL5i�$��lj�-���cdR���#�E	o3lŗ5Z��GRU�B���p^�*K@���M�)�l#]e=���bn6���v�HZ��A�c���ek
�5y�<�����Xb)T�*
����HQ+�2��˘j<��[2+�0�U6nT���W��֖�z�+�f�*�%����'C�]IOl=��ûCh�'.-8��R�`s"���Cw�*ؔd�!�CoJ�V���@�a�Mi�z��Ɠ6�����g�rUk6��NwI��3+`V8�2PW�n�ɺ6дe�6� �m�WZ�/E�қ{�spBW�Q�`;�P�t/p"M<�5�-������d�{��Y�K2�$������/l�#VV]�f��[��{�ßuP�n$�u���jTTNk�ިHl�M��f�ҫ�	T)R��(�
�L&��j+3��v̲Ip�5��:q�,�Y������v2�O%�6�'��9P+��Z�0^н!.�h"�^70}�vI�X1اvӵi�m�K`�w.����aU>���8����ZJ�ߔde�sZd�spX[��o%G!�w�FTx%û��Xd7��vլ���`lsD.���Va���z�*�h�Yܚ�1u�E�o-�b�����
Bm�v�*½��V�Xe	��
�Q����{f�l��{@�b��]�D=KH��;Z�H84f``�ǰ��LY����q��Hd�;��٤�w0P���o���͖�%���ԅU�7��.�1�x�l �)�B�SEV�ۃ~�-q콰�a�O.\���*�6�`����z�8�k���,BГT�	ٶ�ema�K`��x�����NR9H����聘�!�(��
�Ԭ��(E¨�kX�VU�Ў�u��v�x/�2��Cq�h ��Q�l���u	φ�5���Ls�H;���ef��:�W(�N�bkk �e�[b�j�)�f͈���U��|/n?,z%�e�we]"�%G�՝�W�`E��D�L��M'u-Q�A�`��.5,	��6��y�TḂ`@�bm2��h���u��y�5�q��m;�+^3fձ���˳Qڷ���eI�`�r��q��Hˤ��v�[X��V�;y��o�#�+)��p�J�Yv�[{6dCh�D.�в��j���x���v���蜙t0i1�oߙɰ3��"���	�N���r�g2톝��h(�e�652u�U��{C#Bt�,�pe���T���SA��E'dmf�P�x�ˊ��쑐NJn*�J��,:��ZW��k!a�Y��?�f��)S��f����r�iu\��5T������$��O���Jв�C� 8~���6��+�z&�� N�i�:Rt����$S��Mbs(��}�E��ܧVU��Lۃ(h�ׂ���-vjP�Nb�ì��m�]fJ�+Z��1e"���6\d�9.�c�a���Ր���:��1����׻w���/L�Y� Q��"OT���*0^�Wb�) ��E�ZQ2���?���QY�n�A`��	���+`w�۫��
V�A�"���#r5�kJ8`N
����Ŵ�LNa�mv�Z�,R���i�ݠ��hQV]���ȩ����Tj�K!�����x���雮�cL�a�w�� �Gm��+�[;4(�a,n�d��ʼ"b�2����Cn`���[�c��RN��Zun5 k��n�m�-��sj���6��I[v�v#[GPve��f�^ۍ�3p�SA��vT׈ཎX��`�-ҧ6Ҹ�{�enlt��;o!����6u�f��U2$��z޹V�m��&� ����
�w�0b��oN�%@+Գ)�:MGks,�RS��h}�VoB�-la�,��5���r�'�1v|�e[Y�W��]��9A��M��J�\5�!1�ţsk���mU��ra��b��47+j�5��N�D�J��M�Кd7-d�p�D����Փ(����ж�fzrэ�t��/o[D(TygsQ�B�z�m̶��@/��LJ�wn��"Z(u#Ճ��PKDl�ȫcM��i'%��T4�-�ʭˬd���q]�C7V�l�u�@�+*�8���d�uh�)-S7x����ؚ�:�'-+@�E��f��LF�.¥�]3mM�zX	�)V�,�v]���KU�mS,��T�)b�0UȀ�n
Y��e��r��K1E��@\:�����잫Ք�)�w����&4n�ݫ�^�����sRG��K�d�uQ���)�gv7r.![����Ex�,��m��Yy{s(Q �Ji'\��V�v��e3�J��m���!()�\���[2�'�!��k��U�]�ƈR��$���i]f^\0���FށY,(S8��lD^��i���Z� ���$fE�ޱ�z����6[a�HR.�9l����<����#�}2�8�GT[J�6�Qͺl@��=�"���8����ޅf��n\��p��u�Dl³��q+�eZa��7��q�m�Y�r]㿥-���-̣W�Ġ�M9Zn��	��^��9��y��ec��^^6��Q�kizh�V�`짥�܎�d�kf�a�ZR��x8<�
��T�"�V�t�y��
/
��#�&�5I����	���];U�!�C-��n��c��Ly�`Ar�6�ejY�wV�ʳA�vr࣢G�[6��R�:����%G�XA�&e�J�5����˻R�8^gؓ���xaj���V�@*c�B������qK�&�<�(�[-�eَ��6 ��YQz�:2�'��hrG��]����Nl�%�n:���(QU���m�md*���[�.g2�.��ځ�n���^Kq9j���]�d[/	��v��ΌWs6YUm步����/ǉ"�0�i�m�:Z�T�8N���h]���. V�Q4��p�dP�����ݔQ�����雏4���dm��f��`�]n](YL呔�h@X#2݃4#MЏIH`T^�ƨ�;ykf�
�2kV�����W��7w�:��QU�hҝ�2�
�@�M��Yt6Px۵@ⲙ`3���x#KY9A�.+Nkf��6ܸ�Q`yr)C)��L�GL������m!�Di5��.:&��7�F-1���Hi�e��nb�Lr��!�{d�	�j��b�h�7��l���`�3����B1V�6iJ[/!�d�pv|�gSVŪ$��UcE�!��m��kIp��Jj�-ۧr��v��GaS.���ְv�ß<P-Ej�Ъ�F�VVZ�b^�c�JYVF�	�M5V0�7��!�u��#w��^��lY��O�qV��EO�'@�͵�-�^�(�7�+�#g-ˬ��kw6���y�K��� �h��:��x�|�C
�J��+v�0�ۭx7q'�&�#ˣ弭�7�kC�V�7MD�j�*l��Yc���a)��@m㔃�CF�N+�Gʥ`��!�H@���4˸t�ˤ �Cf�V�)�D�J�Is]���-K��Pv�ٵ�4V�`���	����7,�Uȅav�J��Нf�!Y�+��M�����\�J�.��;[�������H�ݶ(�v�5
O�[�%[�Sn����O�͐���Gz��^�pQJ&C�Ad�'�Xս��i �K����%:�:�9yCw��ڊ��8ӳn,HF��7��e�ecv��t�nZ�R�{J�J%j�n�K(ݍE�4x5��CkZ��QLa�7f�tV��JYA"$f��iʗSs��wOdw��2�c��Sf��] T���
��f���I�,�A���֫TP�����nT�H������m�"�D���p�6�:6%��B��F��x�jV��y��Z6[W�U�E�� ���o,,l���pk��V�1csn��K7k�Bq3�TI�䣹Z�5z.P+[Ide�gf��]c.<i�z������Е:u�)� �.dW��M�JvNXG5��6��t�a�4�;D���C2�Cbã&l�^[�b�y��U ���<��ʥwι4�����������U��+��� hX�5ѕ!`�\���_W@�'����ë��:���K[�C�}Ժ��I����/�S�D�f5ԩ���!>$���E�yїo����U����߰����Z[x����E��Eƭܰ�@�_V3"�7�:�q]G�����Vٝ���@RƜ�S�벋�w�HEۈ�5��2̱W�wD���o���Y�9H�!�ܮ�H�L��y�t�Vj�uʺ�����&R ��]a�il��n�[�]o���:�꜖H3vŶ"S!HJY��!�.`���`�+���~{��1��-���g]�;2H"*Pkr6���urk;n�q�/�*��R�w�ө6=	s;I	����;צu5�@Њf�r�a�2��{U�\8�!��Yъ^��jR��a|��9\�ܡ��դ�:�w�89u����Yjf��s̀�ڻ2�0_uuG\zwm=�Sȼ�5Mgp���̣��s���y�i:����^Z���5�[���l�Q1��}yvf��Y,e �U�� ���ۿcGS��,"빉�'Pߎ�����v+Y�n�Z��4��N�S���Ί=��Ӣ�N��w�����e�T��)����ǲf�w��1����� �-�B������M5U���C�w�5�7U���ܨ��yu0K}]dJ�wүl�C�KS�������f���1Qy�D2�QS�έ�zX�o8z��RR���	b�:]��Ky����5R�m�J��&��k�ѣ���-n�N�<���;�h`�V՚x�	�2�gE{��A���!fpͧ��N�_-�g�fȤT��-Kil)���J��d�e1;j�U��A�ۭ.�4���	�.[7�[�I���Cl�&��Ro8�v�\�,0
�۴�1�pzR�om���m��l�zw���T�M=�u�]ѽ4S�B�"6�A>Z5|%�{�ru�U�饽%kb�+2����V�C�Ge-����m��ލ[�v�����r]��lA�c�����7��o��*X��nq�	�\�oq)J�`��Ra�Q��/sU��C��k���'���U���Z�,ytYZ����ݕ��!�6���TA���#�i�ciX����)e[���.3��'׳����S�V;���5ŲQ��rR�ԡO��h�k�2k���p�V�B��%$'*�ɽȕ���`����V�A�ygU>�C8�U����������z�s6�P=�ѓk�Z�1�z�۩���:����2-Z��i�ݍ�Fl�`YFN�A�d�TɎ�����ׇQ�,�F�p��r��R���o��ꪄX2ٜ�IV�qx�J�ۣK���
څ3F�3���5�fVbsc��h�\.��s�0����x��]Ș]k:��-i�o�Vk�v2<���"��Z6.��<�(8Iw6�U�%o*�&�M��Ɵz2�nr������;����"��w�6�6�*�q�}�ٖ����T�n��z�:��\N����f-݈юh��?��g��y�C�5Ov����@�}YY��:�pgLWY;��w��6ݬ4j6��X�	f�x��U9�A�S-�J�c�h�k��`}�ݣ�m��3{p��q̎ʞ���Z��1e���Z_^L�ip]�
RɳN����έ�)��Ӵ�u���vtK�Q���Y�e�wM��^�@f���dC�sC�'�Ɖt{��vs&���u����Bu��"^܃��Ւ�ɹ�M���2/��Ww2�V��w:/n�2�hԎ:�MV(I����k����0�y��pZ�ݘA@:6�9�<ud�o{rZr&$0=+��A��9���*��]�}���&�1�V�J�P�_Wp��i�6r�+�`7t#q����D(��l^<�v�2�{lu��6�/Y���'�Ӛ�u*�Y�Χ�@��1<�TcD|t��(:�;�:�f+�v�0P*
��5��9j�^vY�����qjPt��Ix^�4^��q�Y��6�h�/��#Sg������`�f�PټV�a�D=�V<b�ǘ��]agu��vN��q�K��l��,�e�$�EN�k���FҼ(	0��f�Ř)8��������䡊S���Q��b���K��+��l�Ar��/>j�1U��WF���1�m�џx��bx@\q�͂c�̸�ٖ�_Wi#mdg�L���L�e�ڱ��O�M����e�}�u=#�V�i�|
W���|����[�	0��g���#�������U~K[̈́xq�ZY�m�y���H���H̕�\�j�\M����:�,gB"[��V�m�Yyj:κ��U�:��Y�u��Bᮧ;�����{,6�SyK���OsY\�:��i0� �]�#Q�����h�+�A��Z�/�2I�B�$}�tA ��$:˕�o��R�<�,b9xb;3��g���E3m�je�K��-rͥIU� ��2�z���	����h3�0zq��ݗ�,d���d!q[�)B�SR�w�W6�ï[����ױ+�ӭ�u�A�5s��6�ƾ4�a�G�꫓�:�����p�Y��+۠k8E�0nov[TD���k�u��m`Aܗ��s�3՗�pz\�D����ɖ�=��h�Z��w��k�uiKH� lέG�IY36��R���XIjݬ}V%�LeXM�\gR`:��#�OG*�:=���Lb��^0OLZJ�n���|���M�B�ɮ�H!�1�`7yČ��'�(ZX��k�R�.c.'���v�s4���.GB�njcz7��0,=!Φ+N�6�P�ם�ْ;#B��M*�{S�8��v������;9��� t�1�N�v�R��b�e����P�z�/^���h	t]ozނ3�!t�9}�`�ч����W{E6��K4U�Q��f�6!�v�c��$��Aͣip.�� �ۼݐ�����bB1�Db�'0�::sA;Sp�";�R��kv&P��xiQ4��r�b��a2��M9�ҩ�F�OM�s��Gl.
Yx�e`�=�df��j���M�ˈ�n�y	�X��oo�آк�o�b�=�Z���s���ۤ�M�Ok�YG��x���EWz����k�����g6Nl!�n�̢��s�mme�BЕ��7���[Բ�DJu��x���N�}*��5ݬ�c3��䎉l)XH�ַ*R����v�V�*��Su�˼���!���Y72` �rP�*�ы:�0��hѿ*3u�ã����)\ҵJ`���v(sn�A�h�m]u��#m���ƒ�/r�z�ޓ�"��ǔ�s�yX`=v3����]�է�sm�X��H�T�Fr|���W����1�y��a�l�{���5���@�C�Z*<!R���.�py���0�X���ZR��6�E/���ִr����,��x;� �Ǌ���{L�Cw�j5`֑�P�W��J��CJ��YIO-'���ګ2u�DmF2)�sb(jʧ�TI4P�ᝏ�tV��u-��C�W��!�r ��]�>�Z�J��v�k �:v��8��T�Sn��u��r����Rd"�]�A���4�G3��_�N�aUa�`�)�/��[;ٛq_+n�2�8��¸��Mv�v+� ���J�b�n���Q�ZJ�N��e��nEێC}�*`6��#7�4����s1d�=�k��
�E|])l���P\oM����и6�=P��x��|W=�33qdF�p�*kf�K5����P�haT�U����n_l��7��'[��7m%G�L�uغ�C�FbGe�l�E���R����,m�9�~pu]���\jr�~,U��>��ٍE��C�y:���>T��n8��ᶸ��]ԙ��3�E��Qj��H��⤟f�w�^�D9i�r<A�Bޥ��Χ��GX�t`��R+��u�b�1�p:�Q��{dnA��Tb*�v7�#�WMV�Xr�'�fm=��5�S�`H�Ǘ-�Y8�����ޒ�`
~��=����L��8V(����7F���sp���v}�XJ����>@R7 `�D��\=S2�ײ��ŻM�c�D�]w�M�Y�w����e�w�L2'W�r�|��Ơ��Ul5.���\����c`��@ ��Gw���� ��PG[�nX7�d�*��eXNުS�6�i��\�����c(�����!�3���!X��D���"������u�y6��8 ��v�'<����.� RB{�Fo��Þ���]��9���Cj&m��u�/P�=wcJӢ��w!�����p�r1E�{s2���=�(X��D�Y��9�m�1�4��c�Jfʚ�:4S�4���"���q"��z4�F��hm0�F9sf�wn�"¥а���{�n���n[���	WB�!d��{��um��;_6X�ŽVu`6�bw�-��å\wΜiٴLw��9�Z�بj�}Ίb�v���k�G��(�RݭĪhdƩs��w2b�E�H���X�5��h"�Ҿ�ñ�Y�#�jZ�+VKΨ2Y{��\�����u�ܛ�*�f.�v�=�t��	3z�"�Z�j�ht[���z����3�	�a�eh����H�`��;d�:����\#���wٹ�S�ƥ�RM"�)�x{��o8�J���Q���6ӗ�풞�jV�K�Å��Zܴ�м59������[]&L$�7�9�u��Q]����a��nq]�e����3w]��)��e붨f1=�[Zv$L�=n�p�r���j�"��Q��*QS:��r��SN��ۧK
|��ћ
��8��ŷ����b��q�޽.E�{�
�� p�,.���&�Ԛm����l��hOr���.�M��3${�2U(�WF�'p��壅�� �1��3�B�ꕲ.��q	Z������
ɍe�D�?�!�12��<�<��c^��rR��;s.b���@)E�%�zC�-�áW�_��dݥ�c�s�(�n؜Xa�MT��R;��(��Zr��G zb}����7�1�cά�t+���H�ೊ�3M��fh��3�0�1=�4)Sñ!S�ܻ�[��˧6���!�V���4�U����Jf���r�,�Fu��+q�,��'�R�d���"��5��)�]ϛ[�P��!��X�[���bwm�V2�;��V�%`�Sɷ�Q�����H�}�Z�eMzx�`	Kf\�y\�,,�4�v�j@csa��݌(��f�ۯ]����ҳ���l�4R�/fXt��cm9�>�9�R�÷v�mꜴ��b�VS�ʴ�ɚJ]��n�<��W5Km�i�(sw	��N�������+o`>O����`�%~��j$̫K}�`�Cx�:b��ށoylX�}9��5n�$f�I\���f��(��c�G����3r�f��s�����;��%m��e�읬rF���J�����Ǉ�㱝\�zE�8l���2s�Y$�	�$]G��
9BR�CN�*Y
�9V�|u2����6B,���B����t$2K������Ғ��_^#�@���S/hdi��L�'$�J��o�7�
QΫ'����G$5�[�׽!�$������7��y��;�'���mӯ?o��7y>x�R�X�z+�R�e$�-�ݮ�`���!Em����1Ͷ�5;o��],MT���`���I7���������YQ[!0��wp�|�m+���l���4ke方MWO���M܂��q2��1����c8�[�Q:��1�L����v�gs�-v�d��s�ڪ�z�2t��w�c��K�T�9頺p���H�ʵ��K�͖�V�z�U��P$�(��'\.����u%�]\�����x[�� {�y�{(�L��4;^�f��a����k�Z�Y������F`
���-�B�r޸��KӋ^�B��ϳ.Li5�\�l���ɪ=[�Z�49X����9�θ�LZ�x��F�Dj����a��!�p6\���0����r+�վX]I,�ﰼ���]қ�3+��k]�6y��Nu��mG8>�65�!�vK�	j�+Y��^��\+(OiԄ�A���;�������v�Ӡ��n�%E��
��<k���*)�5=J�*ą�خ�\�c�JT��1���R�f�&=B��վ^Y�g��rz�ȼ^�ͮ�t�U�� ��b�'w��(���N7X���DUHҘ�"�ͧK�����ʕ}�+(� �ǚ]qnA���:m��9�c�3�N�.�n�;5��ɧg[־]�H�1��ހ���2�I�d���m�uEm�o�
���gV�R�qX���h�H�ˎ��}ݗ��"�Rc�P�r��1Q�%����k�I۹kc�Z�qNn�,�ʔJ�x��M6�n񥺼�Y����e,�:jеp���F��9��\b�W8ͼN�A2��
���M��Y]7vܓ�u�+T=��Y��6����boT{���	w%�ɷ��P�-v��.K��0��]�NA9�pt�[RZw �e���Za�����_KW�1�AIdZc:\�L,��ok0�V	t!��4l�%�̬�58��X��{O�V�G�o� N�0;ЀT�v�{uv�"�<�!c}2��>l�v{ii��d��sQ�=MX;A�7j,q�5i��ؕ�V�)���ڕ�C_-�s�FX�uC!���(���rlk���];^���9hճ�M��l=K&��<�}��\;z�X0����z�ų(Z��:�nQ�^lJ��*�ԻX"q�Y�Ao��f�;��5jup�d�o���~�B�HH`B����oL��p3�m~:��sl�T�(  �c;&=*c4�J��`8�)�<(k�S�u��*��`�L<
� �A��B!�5����̱�[�n�BP��&��׋����z��k��<䢡�W����s%ڊ���r_s9p��+)XY�pq�1v��鬵�����F:�r����Z�'p�|�T&F��X��WΔ��DzP��5��o*;�����,;��!
�`��Jq����fŎ�����)��n�Y��m+����6�{m�/SC�o�:����
���[7C6���ɑ�ymT-��N��o�r�ȫ5�k�*��zM���,Ё�˛�+�t��{X�BvT��w�_Ca�U�oq|p��7h��VL[��bQ�|�z�V�v[ue�=ζK3S�x����s�X�1865q�;�_rJ�8��&�qoflw�Ѯ|_V�ف�#�iC�4�:� �̸����яh>��p��$�i��)P��6�R/zd�4�q)LT�H��Hz��@�vV���ɚ�
﷾���$�|h���5�V��[�&�+�M⾡��i�}.ܫz�������ϵ�{���Y�f�ܿ�HJ��ʰ�ۼ���괒�]��b�`X�I^�e�Jn�l�i�tU9 ��.�c�ۦ�@�;�z�v^F�'f�~�W����@�4r($��Gb��t6 ӺuQ
^rvB��ە��μr@�����T��|+u�2[I���ۖV�& 5�;�}mY ���W̊�
�Vmk��7G��r�D�NT7G,-q��B�p�i���T�}�)wP�w��j%��ǧ1IOj�mP]X�M&�Q�3�N{�����n�5��6n���meJ�&���m�S�s�ks���-ѩQh'n����Z����	\���q���;�,�0��0�|��+G�5��T�,E��F	1��r�a��V;9�k.n��LbSŠ[T�Eos:���:�S��fskBai���]B�;J�v���E�7�t}c�X��wWNV`�5�+;9NT�O'4~�u7]�ﵴ+�8GF�WP��ٰ�_h��.�އ7M!2>�gUػ�qj����2��v#kF�Pƞ�$�6�l¯0_M�s��(f���QS��޸ԏ��fmb�`�h�Iv��g�T�اƗ5�tp����[���ֳPW��=����q'���(��#ui����;z=�OC�UTGN�=��U5Q��K
"��K��B�l��2�c����."T��nr�6K�a�yh1;��ؖ�Y6����Y!��f�֤�ud�4�9���sn���{�Յq��%�I�{�}�c�}hWMI��,��'�Yw�(e�Rn��hkE�����$��B]��L IyW�I�ܼ�˞Q�dJ�6)��q���2m_%z�֝	�pr�]���8����jmAs��-_hf";5k6���Ju����m.l&� ��{��RnY���E��U�^ɔ�H_r&f��]0oN�Q�^p|;����]���d�*J ����j$b̓�.�KS��1ꭱ�C��Fe�qX�&���(��ό*�|6�-�Cq<9�)׽Lp8ś�CV�s5&�vՅ��.O*�ɮ�C#���Őc�8�E�U<�ė�;��,�e�N쩓�g#�Ȋt�6�%e�#�6���R�k]XLɛc��2rD{!�%L��/����ޔu]�Fbg+��
i��wwF|z;��[��&Qv� N.�q�}YӰD��\�>ح�e��}�Ie�&dk���%u�6�7u�t6��F2\�v�%v�������N������m˗9s���g��-��}�l��ͽ�d�[��V��ɻ��֍RiƲ%o0)B^�}z�'�,*:�e�Wn.��uHvV.:�G�]��t쩺��d��e՝A$��d�����#kȢ�WL�ܸN��wD��jXVʨ&>܄�}�AJ�V���6�Î��A���Y4�6 &��ec6�hu(T��u��ۮ�j�JM�5������+R)���m�
ν�3)�c�m�h&obK�+��o��a��sΏ0vID��T������jL�Hh.����ן�U��+[�V��Ь[��</�Rn��"Ya,j���5Y�i��l!W5��Gp=Y���gʙ���-i�a�1����"m�/Ÿ�N�K]{���u�������I ���������ɚ�hD������^F��6؛m����ۢ_VIĜΰS#Q��X�|0+�oN�lf�|�:QVb��Uth�(�.7NVM���iLrx}�hj���9�-!����!���31�/����]}�����0f�Nם����G>ۺ�r;'K�mjT�K���J�7�:1t���TӔ�*NI&1<�/_Ww��+�Q݈CtZYRj��d�tv�YM.�^�W,��GvS��'�wA�����I�{(�K2��|ɭ`.r,��i�D�3�[��	3�*PWf�d�Ty�J��4�kpDҭ6>Y�� ��C���Y�5ݬJ�oZ�s^��ID<S=9W��b��t���+��Ɯ��bV,hrtѯ7qFܬ�x&j�3��6�볝y֖y�����$��N0e��O��*��2T坍��&�X�<�I����3�BJ�|��]��@��j���Gw��/;$�#]�n��&�]Ib�/l�=�����4e��ؐ2e��7����(t�8������cc�9�#��*�I��u�U�gF�cs�i����sUۻ.���r�
��a&��%ru�l�\�̊��X�L�u��Z=6i�7;Gj󸋣H�aL���|�9hv�w��n������Z�tZ&N�[N���;���[�	Ǵ-mǶY�aB�bZ]��D���խ�N�jԭk&�h��s�ǆ��92��s �K���"[�T�� �H���f���FT�(q
K=*ʧcpS9tc�- Uw�Ո����X�Zz�����v6��I��}OXk������.�7Z֭w�{Y��k^�U:"��;�j�J��;��|�Y�#z��Kt8i"�+(���O_Zgk�%n�R��B�b5�0�M���ϡ�T�U[�F�MU�X����A*S��!7�=�7��U�%ah};X&���s1f����|�au��맦���uW^'$�+�s �4�.i��#�@7g�R�vĠ�.*1��]����$�7�u*��Kl�ײ��yx���l����	]�N���CLk�*A���-*G�tn�]⼣*>���UεdYܹ�4Fޝ%u{#����6vZzp\3(�������P�E2�F�'z+n��q���e�y���;�&L��R`��)	L8�oۃ%G[Ȧ�vd/_U�(uо|t�̻��XO)�).'�(Z�vQ �B�����]�(ov�Ν*+���z:Z�#�Q��zMZU 7dژ�n�ʄ�˫�oA�c��j��F��%���9���vY�t��
.���vDT�x�-Nz3{�"�i>���q!QS9�5�]��Ճg5���;ĵ�7�y�� E�q�X�� Od8�J�s�#c�Zp���m�	�u�S��sR�/�I�	��%
y��,�{VM�X��)�8��{Y�aD���Ҳw*\��9�OS3!��Pa5��o�or-��hhU����:�k)ޕ��:f���p���pCLF�ehV�� �g�-5gX���������u��F����tR�'�ɜ1ņ�^v�Ƨc������';��;q���T��W8��B�����)=X�=�Ք���}Q��}ڍrX�P��k��W&���5H^�]\�P7A2�n�tm��Ȣ�P�k�XN*�7�ok�׌��fguG՛4j,Fh��ЮU�O`�"�9�xP��#"٤���pm��zdLU��lOb
5J���o��܉��hv�s���S��._-O$�u3H��h�z���m!vR�#/t�����)�H̹�VcvU\\ho_N��F���M���r9���tk�d��R⎒EX��O�\"�pt���z�4�ku�wRn4�x�)q/��kf\��T-��A�geL���
P@I�uLǰ&ʽ��J^\j�����:Qf^ٮ���N�g�X�t��,泗��ϴKZ�}6Y�КX�6�WIG;Aǈ��Ktr}׏��l��7]KA'0K�b����m@�+7D#2��̭rZۧ��ɋCU�:V�j��ϭ�nYH��ڌ��"���b6�+:�t�C1�Y�wwW�|l�#�Be�mm]�`&����'��(A$�NѾT:��4���Q�%�d7R�Vn����t��}E!�u�·��n�p�s������`^��Y�������=bmu�����#KhL޵EQY��������7h�m�\9�>N�����.�Z�<�[׭�p�E�P�(�����T�4��+W;�§u��1������0=��݊�4�.��zue*d�i(�7h!x���ɭ�%��M��WH)V��L<���rK*se	Y��wm�6�@o3�ëi�p�fd��6T0�&V�#G�
;����a�m���h
8���Yi����v�G3�3�u�"�GN8�K�;.�5��,QG�*k�u8K��r�����0M��F]��֎w�gcRu;S!c�]Wi��[�2�:XS�kz�w�F����b^�6��qbib��9zH�$�{n�K�Z�t�[ȍ�R�q��79j�5�2��*͘'_:qtΚ��r���E�J�84���#����9�0�q\�Z°亳-����n:@M�@JJ����ib�9�?S�tb7u$'vX��H���́�:�.9�(��y���	3+/�g>��^B��Y���9�)��$h�<g���W�1�{n���{wY�Vs&n��:u�a�ByF#D:5xN�v�tv�wf�l�EF]��4"l���W,y	�X}Դ�V��c��GM���^P�vr�����BN����W����k~<
�������ɛ1h$uQ��	���0�ː��E�@�ٔ;�H���s�Y=��\C�x(!lv�)��ٜ��c�&<֮��R���-��6����G8n��:�C��`��c�S�n��6�%��,�R�/1��%�Z�]�(m�K�EwX-:�Ҕ���@����v�k�^�\�m�s��&.{�si����6t�,����9���`��V{~�:U���:hmZd�F<�yga����z�r�}z�޹ug;CM��MРMeY
iEeCf������ż�zV�׀A�)��2T�x��E+4��ʘb�LT;�[��qS�Uβ
�f]34���$�b\�tc�N���2��F8��u"��ڪ��!�ۇ�%n����C�p1�Zx��X�AiҿiʧT�Ƴ�㘶dES�;a�C�y�+���Ź��S`��Σ�>9J�b5����e.V]���k�xӻ5ua�Y	\��Eh���)B��/A��ɻ�wWA�{�2)�_m��J}o�S9�%5�Ez�/��W��(��Y}�ض�F$�{�%G�HR�H��̫�[E�OZ���7/2��4��p�[SG)�&��]�U����h��D���U��hAU.�7L��3%�iU�6\%�n%��ۑM�fnŨ�H�<zx���W�A�Ur������]%���	`�%;����[�5c�p݊q���v�i!ƶaMڑu]p��K�ag�)�KiGY0�{�QQ��"-o6����;D�$�����OREp$����%-w5ס��B�
r'1�N92n<d�����檦;4hV�	�$���Z2����;�"͙� �t��W�ە�2'E&�Df�����W+�up�}�*<-َ�ښEi3Ʋ�Pן`�J��dI��M��҄Mq�����0վ}���}kb]���0�D�&^0�m��.
��y��^�h�nE7��o�p�-Yn�5�j���3�CwR8���LWXD��j��&��%�+����:̉���i�����KL|�c���V���D�
�f�o���Wc{A��N�Yqc��^Q��I1��v��Ef�9i;�r�c!��Q]c�%!�-�c3xhy;�dN��l� ��a7� C����nU�R�tgY�fe5>SM�(��+�qs�C� &�8"�1�@{z�=T��Χ���(Ѕ� '�H1+�� �C{��8Hgv%%���[Sƻ��4BUGy�Am��U�w��[m�L��)����@�&d��k,��1�����Q^��h�FlѼ5��dI�W��f�
�J<H��F/:��e�v�o$�3͋��<��Z(�����Jжc�7[rY@{�x�;���zS�I0��m\ֆ��T۶1^�z%�V4�}ΉC��#5�s�5p��sI&�8�4P�d��6�8�:ҩl�c����#�`����	��I��	�yϹjWo1����v����C7 ���\:�N��U�ˬ2x�����\Xd=(�w^i�c�hShrQ��c7[#��|Iv�gZ&ҭy�ձ���],�\[�rq1,L���q�j嫫j)��vX�a�p()la�'hYw¶���Φ�/A�i�8�u3K��u.G�]�٠�\����v�4v�څ���\}�t��f�(�w�͋	�odCj�n��_�_���N�V������.\�+10�$@_XPN�N�TY���&ޤZ�h�w�\{#�^9E+N� S��k�R��jvc7������u��`�]-ܺ��)�
é��ڸ�-6���H+�4�*�2�D�v#kJi���y����K�'�\�5��$�	'�<��<����=A��*@��r��❥]��uY-�	�gs-���ܴA�Q��0�ɸGSӽS���f��U!���9�CFq�r,�7��������4ҥ	�n;�u����m��Vs��.�c����#�ӥm�\ ƕ$f�MS�����Y:{z9�i�܏Z��L��) aZx��WZ�6��������p2��'�awT�R.������j	�����I��!�Rf��t8���K#��.���f�1�`��(�!�	�{���VL��wv\ܐ�4���-���9��� �iR㝘7No:�|�7�)�8�M+�Z뇠�����ժe>8yM��4���l����� ұ�������uӶ�X��!B��#t!zj��s�u#�Y��X�rfpӬn��p��F�+,7ħ��g19�CT�R6����J�3�[�|(%�!.֬��.�4Y����ه�r2�6�[oK�|;�7Z�N�Ąss��Psdd��x5I����c�����@H�!rjă+���kj�2;���Ԫ"�V�9�@Jw7N��װ�� '}z��2�8Y	�1�C�ZR��雾���ఔ�x}r89�~�y��qWW%�2��'S�Z�f�5]r�bkr�o 
�\E���S�'ܻbs���(Z�j��)�:;WL�Q����7�A�]ե1`h��9�;�34P���͚�A�5
�Z<��Y�Ll�ɕr�A5	������QKv��e�W�!8Oc��]�u_>�=��R)�$��$�@K�Dejڵ��X�"Z�*2�,Db��j�F���Ec-���%��*T��Db�j�J���E"��,QJ��KlQ���j�"�m�(1��2ڠ�[UEF�*�%��F,��1DA�kDV(�R�"�D��E�QTF�Q��aYZ�`�EAX�X�(*��,AFX#UUDkAV((���6V�`,-��Y
�DTTV(6ʪ*""����DF,��5%E�J���$AZ�E�,-,EDQEQTD1�DUYF2�%�TFE-)-(�T*�R�"��1J�b-Fؠ��1���
�#`�ł���e��JE��DJՊ#*�����"�*�QAc��E�E��
�V*��cZ��*��
�)FJZ�����eU`��DX�� �QdQ��E-l��""���jV�X�[EEAG�� �(:WM��{&�b>������n.}2\ڴ�Y*s���<E&$���0��\��JG):���S%s��\��d�H����ڳh�2�����VW(z8&cI�C���s����Hc@��x��?�������U�=�����xuG
nX���Z�!W[&X	�w��h�Q�_��EuDc�,`�G��u_�p�8�z�����`��Ī��	�7X�F8B�]2�7�Z�ET�(\<f�T^9�:/gBwC)3��>��0�vV�{�=a�b��^%{$���4p9ee����/�W��j�ǲ�};"�7r��XZ:!a�k�y]^�'������T�!\30�Ta��¡i4)�P������Q�����(E�Jf-\�O�s��=p��
�qyQM��u�V{h�1S�،��sB�0��e�d�����g�`�����q���5�߼zh���qۂ�gc�Z����O8LMMe�&�f#�Z�˳�"+z�b+М�a]3�:�%.s�j�{^xQm;K�ɕ�z�m���E���ӡᨣ�^V* ->�-�͘p�y[hq�;�KWgdK��D����d��h^���duF��1�pUZw��\s|fܪ"'oL��Ԙ��q��iE.(�:��OP�W�%�۴�{0��s/��ˠ�W+7�R||"L������}|z^��ڤ�2��uQNNR�;zYӧ�������uu�)��q�
g�����U�T0�|���71����ǅ��uo����}�mؘ���s��f.�T��K=j|2w�c<����U_�{e�8tb�;F����.7omb�z��VM�841b��������T�\7y{G!����@��'f`S�+Y�U�����{>�R�3���.$u��+�c���t�UiZ3�^���o#7Wъɮ�n�[�әJŤ%�t�h.��q57��@��wT���j/������X1(0�jb�%����w�qҸ�C���3��<#Q���	)�g����$뉚�Qv)���R�T��\xs�T=T�����ePZOQu�p���:QBq��Ln9��Fv�m�'��Ԋ�`��{����f��[(C����r�G�R��rC�$r'�)��T�TnH���dM!8�L]���1~Ξ��ߐ}�)��yFZ�(�M"�t����]�Z&W i�."j'��|�j8/�%3}���,T�Q�3p!�N�6N͔�w\ ����N�ht��L���v�] �HB��a�E�i�-d<�ɛ݊�җ%a��C��{�����]o�V~w�e��Ž��t.���Bl�5�mr�}tp<0��0s�t^�:�ᙜ��ܐ��Q�}$0������¥���r��X��mk흯
gk�#, `�Zu�Q��,=�T���=�E��Z��MM�Ui̶��ǎ[��o�'���#��:X�K)e�8@�W6*1��	�qK"�s���s^p�n��w�kY�dX�p�q�}N�;����֐b2�}t����#�&�-���t�b��1���y�QJoL������3�`�7�:�5Zن�����tj���E��!�8t@w{,&�&}~�o*�{�M!�#N�N�,��f�x����WQn��:�H��;fp�ٻZ-\{jFg�N����$�@�Y��١]�� cZ���l�5EC#������F('q����V�#n:|�:�c�
�Z�R��q�{z޷�՛o5��`�D�����o�)��k���X=�D�[n&qV5T���K#����w���[�w���NP�L����*�5!`�O]�Z~*�[8Oe�9�Kyyw~�8R8yV3���Ktٌ�3�d�RF�3H]��N�!��A[�&̓٤M��9����W��x�qP�p��r`���X�'z��!�V����K)
i֑��q�w/	��J��{dps����Aߧ�����b�%b����������O��e����s�vG���
u�f����q�F�Y0s��ɼ3s�Yj��`WÐʼ�7G�2x���:���'(�:ۨ|P�yE��`��B�
hglˇG�"���k����2lGI�qn���0��t[��7,0�FZ����[������r.��N
�Nܥ�U�h�U@d�n&-[_G�"�͸}��`������m�L=[���U�{3:�m-�+G+�8#�%P O9`�<zA�炝R)���x�x`g�g�kA\���1�׽�hb{Զ�A�Hl��T���`�3��"�â0N��7rT�V�DjA�ΒG�]ZC�XW��eʏ�^V@���ؑ�Ǒ(N=�:X�8Ԓ��.�'6w9�.F 	�B2�
G�`�s~J&ÿBs^�b�kǶ�*��
uH�q���S�9�����s˚����W8��tF:�"����0�W�NmQ�n��yN����5�7�i�e�7\�ؔ�MF�hXD�c�~Py]�����b��f� �U��u=�>N�M��$�;}�U��x��Z4�~�Ud�3V<:E�S��c>�ϒ7��9t��ʚ�̻���F�9�����_{bo� �AųM��;�^�w�=WEV�Mܴ��Ş*�>�֤�˲LסD=�р�O{hrot�)���OV7�웢t�\�
��t��ۇ���7zq�r�v��MN[*�;��N�3���v��7{J��+T�Z4b����,.�ϙ�@}JȨ1�DK�i\MU6��]�'���X�9�j��ʐL�c�=ofK��7q~VY)Ѐ�8mǱ}�&�y�]����E)/F��#Q�F�b.8�5%1w��p�s�x�>� �3Z9zt*�K)K�(+О�>̭|U.X>�[��a���JnP�u�^�r���WQ�כTF�U�uq��:w�U�KYA����@��Hy�U����>�b�*>4>�5�p}�_�7�+�*ɩJ&�-x*q5�BɇxVw
B�����$k��o�}���
�"����o{r�
�&��IUhA��Z'XLR1�'�ex�<�]��T���M�<�G�9+�gL��{�z���/��5�(=q���)�����V����"ͣ;��4�^����꧴[�iL-��{]��臅+TŪ����(���0DYTB�fa��1�Pȱh�\15�a%����{�Z��~Sa��yg��w%��x]_�<b��d\'&�%���p[�$d��ˤ�:���%�[��K1�qi]�h7M��$���k�qc���䫞�^�i;��^qnoT���`�Fhg�.T�0.5%zu
� @WM��q
��(oZ�ۯ���ϳ���Wb�)s�OrG�y���ځӷ�/�R���b��0�xi�X;<*��\�1�=qZ���e@T%k�)�>3�+�N�xJMA޵U��ӭ���/a���T73=�Rkp5w�(?��;�<נ�F��ƽv�"VTv<�?*�k�\� �k`���~��F�qt&5���Tl��н/�>������,{�K6��W�0�9��n�n�!
���"sfu0s�q�^[��&���5�:6ٓ�	�lGE��J�e��=�jWwsQ�0 �`�6f6����ŝ�n�+���U���v�Uw�{x[2*+M�X���-�Ò�(�~���t�"�,B2K㏦��vW�Q=�w����Mf�5����<~Y��`�^���p���}
^�*��:��|�f�	���aZT���:��8�m�ͷ+��Q;Z��m�c��E{��:ey/��g	T����G�����mWI� a�{+$��=ãͧhg���G��lN��|Q�=�W`E��~��
K��v1O�����'Pzz�e�u�� W�=��t���Pu�8�T,ȩ�v���Բ�89�yw6���Sl!H�R��z��4̚���������㗂�-n�nB�ޢӀ�.��M�Wt��y}W7%"�ܦދ��䫬i(c�tQ������z�um�r0�Q�Xc�+������V���u\��<J#�A2G�%�"�W23�c�j��9�}GWj]�?CJ��!�5�3��� .�/�UObWS'�� ���m��rq����VW.p�P��b���v��-���Z�4=���S�;ldF����i�&Q4q%m�>�xe36���O�_���І
9)��Gp��b�)�php��:؉Hn��~�Y�)��^=>�^�Q�W�W�ճ�FU `����E#� �����o��/���g��R��Z�ҽ��V_��JS��X����e;�!a��wh���@�Y6���xuw.�ӆ ��ډ����s�L��,����S�R�-�)�8,X���};/���)��4�BT��n׌�M.�E���b꼢���@��P�3:�;c�.3%��\�!�]\�)тv/)5��Kpk�m�����=���Ѳa������󪛹N̽L�X	G�ATlpV���։��|��MI;�E�O���x\$�V�H$��qS����ڎ�z��L��c/E;5-�"��n��E��q��sՕ��L�u3�g�����]�qL��nE�9����r�V����
���[�j
�:�]�I�Ϩ>��Ͳ�t���g_�V�|{
w�ʸ���t�ۯ1�d��ex�8��g�����t�+�϶��ۈ���W}W��&R�9�
ކڮ�A�+A����8B��p+g+�f%��OU� y3�F[��CǶ�v!���v5�N:�zk��YN�N�r���8%��V����Y>J�
T0{���&�7�<��ʏ({ݲ�`���x/2��n�1��FɿrTGk�t��ӷemgOu�W
}[�mB��8��F�J��u��8V�p5�ssO���g��|na�m�3;wA׺��{�>�l���mA]�T��v�w-��Xa�ф/ڧDv��7�l�����s)Ң[36�+�Q�-eՈ��uTk�F�hН����l;Vʺ��Ί��0f�{�����f���ACr�po�<��oH�qT�3�P�Ge2k=��rӨ��;����1C1��4p��R��~E��"6ty
�TQ�9�`��h�֡�+;w��b�� �f*Yɩ�5��;����#6��X��wAu�z@�8|>�>
W��>m�ݽ`�D����cF����Y���q-G��Qޚ�ڷ�]=.#8�2�mY/�Z��f�T3����A��t�����m��v9}âq�|Es��K�S�2�{�T7UYJ�U�Yb/ �|��Gm6����=9��M��{�E-+p�3�������b�pӷ�T]*�t%��r������ٙ���=ZQ��ږP��.98#+���m�)��Q6�5�b�h��ɖ��.��5��@;oŨ�0��'aqW89�GP1��H��b6�P7�Ho���0�*��X�eUn��r5-y��'1�1[zj�q�:��1ae�.�0���R�c�yQocܓ}�ȮѽJFJz�۩��m��{���57���F�/Պ��Uп��	�� ���bVE�
�,t��)t�#d ����ܡ��0��v
�<����RWƚ6y]ǻ�*#_U���-�������z����nxp�}1�ɨy�D�Ø̢4H�a��K:��S��Q5
g;�5ƙb/��	)��N�F�U�t��kGv��Y�n�	�x9��*vX�[��.Z(X���)�m׮���nz�i&��\lؾ�w�}������o��x$��Z���*C֜����`�l}�Dwf+��.�x|>qX$������pF8S�%2���;b�A�I.W�����a��Y�o�Y3�3��Y
��k($���վ��Qk���I���vZ���,ǚ�# ��c3ئnv�Vٖ���o]*9�od��5��Wb�6�n]�"bbu�\�ɻ��t\�RVuې=��q�Ѕ}x!0���:�E#!@�K�O�v�x�.�	�j�����o�#��!!<Gz�uQ��9�Mҿ}��x���<�Xdu�$
m��q��d힍1=���R�"�\S���ܗJ2q<}-*H��
ʭ�)�Ş�{;��tL�eQ
���4f6B@�B�3n���066��{�a�,�4=�O��O�;Y֜�	�oL���Kw��"���({L|e
�9հ.��4e�l<r�^��ׄsg{�v��ms�&�RNs7a_���T&5����\!~��	��h>��"��1��e�3y�0Þz����Wr�H6��&���WɃ����+�_��VY�].�u���)�)f6�}�s|;���Pm5D�s��M�a.͉�����duF���zM�X��af쫨�ums�gf�����A?�z�ܯ*L}2�ߍ�vφb�b����6y�Mw�p?VM�98!�1����U���rw�c<��6��Ȉ#c��ϼ�c��EcC�f��y��A�ɝH���&[妷�V��M-jV)���Lj�ð��y�y\*�f.��:$8�F\7o�Jg+0���;�E���򤔭śB�>c-�Ypf��@�v���=t��cf��c����ݢ;�Z��h`�efd����ʤ�.��ɗwZ��g���m[�-���OJ�8ۣ�S��ڿ���&��R���P�Bu��E�N3W��Uݼ���R�ٴ��v�sF�J�9̗�ca)��;��rٸ%Cp�w�X��W8M$�]y�$���s P\׉��X�t
����E�nr��`Q#�N�0]��+.�ɣ�=��m�2e��έ�5;��M9A���K�}w*;�y[Ӄ�qR��%�]Û��rƝf�fk����bQv���MԕBrQu���Ey��T�	36��OB��wۯz���|0#`^e(R!Ҧpe�.�A6^8qP�7f����S�]Ou�z�Q��* ˩����2j�9J�҆#Գ/"8j59b��v��/�.��"�u:�pV���)�r�%W9�e�s���ұ�h�;Ѹ��kϢ+^�e��:l5�_�أV� NۤuJ�����J7n�:�O�Z]e����Ġ��S�n\E������٠]Lx�q
i��]�*���ԫ��/��z�����}eCQ� �V�c�V3�n�.!d�O\G��Mp�Jg�ރ܏5x�� �l�u��6+Xт��d�1��J�_�@РhV�-�)r�J��3�O[�m;�%�Õ5f�V��$�M�3���5�髧B!:&�oL/��\��w��5��n�s��';���/Rr��[�F;8Â���o���e��۠Lk7(�֡Z�]�SXͼ��*�j$S���(�㐦���T�[*����R̛�w%�U֋�����áE�H���|�����֐���Q��ި��q���go�X���Oy��ۅ#�p=ٵu�e��3	��m��LCv�1E<���<Pz-�s2K�dU��A� ���2(PH�� ��R��M>uc7$q�Wgk�V�N�DV�8��g�l����Ѻ879���V��'���\�*��e��P��(���،U/:�
�qUܒТ�W]�� �l��Q�M&��&k8C�y�������ɜK"�@?r������-�/�ef뻁J��T�s�T������Q�X�umf�F�s˄���j*�W�֬buڥ�C&jx�D�`r�O&�7l� u:�:a�B���U���,%�6�7��G�b�wW>��H\�#��J��tIY~�v\w�ۊ��
�����K6�v��H��˳)�a�Z��l���Qô�}YL�z(��
�EUE�em�EE�EA
*�*X"��",UaR�UbD�R(�V#UU�� ��*DJ°X���FEm�UVDDQ�b,E,UEkb��DU�-lVX",Db�*%J�**
�%k1��1b���1A"��("�"1�b,UdEQ���Qb�b��0b��b1mX�mD`�b(�"ѕ�(�JX�EJ�F��)E`�b�*�"��
�X��TAEF ����EEb**�"*�"�(�"�����Q�FEIEX�Q��"��QEbV� �DDPDc����
�Q���X*��2*��b0X�(�#
�Q"��*��1Ee���DH� �V�Q����Tm
"�E�APV*(� �"(�V,V"�1Zʊ�1AQ
�P@UDQ�D��߷�O����~��P"ޛ�G�;��[,�0�0q�z�8�d̆@�e�3v���\WL���M+�����Z^�i�uG*块;���u�>?ơg���Ǌq�`�xa�-Κ
���1w	֏2��F�r(�<s�vAY�5�X8eW����f=PuK]���*ᢻ�j���fK��0��X���D�lkj�k�ut���b��M��p�:�!"��������T�h�pB�W�2�kW~�p6����hg���G�b7ʫ�F'��N��
�J=�?�z��
��w�,��������b��t�V9מ�ZRw\�<J#b8�
���"q�T��:3t�V�C���
m+��<#���7(C����z�t��,�&���pq�N̛�u����d���fxG���U���e
��mL_���K+��>C��a����~u�����
�|�}�,KS���,;�iamO�&O���f��<�wQ��f���X��#͠��N����
`��
�z�|�9�l�5���?�>�f�o1 j��$b��EQ����	?8J�����R��R������|\��Q�i����+����`bμ��V'a�NN��8ٹ��ٌ_���c�}�_�i��wϚt��v�h�bP����+5�Ъ-�;���@�v{�YkM�vr�v�|����:h��M9F����s�Ӆ�Z�0����K=����D��|jr;�0�������M���`(CAO�����g)�)�[�W��*�gKr+��5~��{��CG�H�k��O���Xj�}��fVꩉT��X+���j�t|�a`-W��hK'W~����\�;�:.�X�>م�Kpj#�m�����=��� eS�z����=��]~�Tdʳ~��ˌ��H���>Bk�4y'z����47mG��{�W*���c�����-�:�Hz�g�B�����c��y��|*��|�Is+ݥ�켝5{7�R'���V,\F��k+z� h�E���f`�;����`]uဿN��gz5fl먮�ũy.GD�Z�X��$�ýn�����}����GBu�EcJ�
t��e5��>��%y^t}Kz��L�����(�9T�7�n�!p��
5^ܫC~}4[K����j7S��nb%'�ly
���w2��nb��p�	һ�]G\7P�����[9y���byZ��O�T݆P��L��NR}��
�P^���r�����)�j�a�ǜ�2`���8�o�+�Y'��`��$j�����4������iG�w+w�S��m�}	Nf�O|]�l�xl�R�����-�>��qC#�����Nj{b�ju�=Ѯ�.�^�}UWm�e�R�yX�c�Gځ��7v;�e�����v�ؿs�#�+�����X�Q�-TЀ5w��!p4hOj��y_>��#��5m��Sκh+�d��ۖ�ǝA��բ,̛8�&)���9��IV�Zx���Ma~�cB�u������l\<��8x��4����3��=Da��.�������E��F�1�v��NB1Cj
e��.��]}�������l�JK��+|G�����!5��8�ΐ7`،���S���l4��a�����D���m�e/m�o�����)�f�OK�op6s�s����;1THͩb6(�D7���X�܉�4E�'����N{��{>�u�bR8=�S5]�=q{��[�D<b��|�,U�JR�w�����<MJ����)Y~XC���,0��+�-9�K'bە7ڛ�뵇��,�[246���AѼ5��`=Sn���,TuI_#a���k�1^�r��|��������W�c[���R��|���k�ˇ����4�:��n���Kγ{<�����iy����݋������ew8��[�˰��촴:+of��I�iY�	��S�pV�5�̼`�ֹ�mֵ}����͕�|#|��cɇ0lU8�u��n��B����nk�x�Cf����JU����⿡�tRy��E��,Á1Gw$4xK,G���U'?J��^��5�
��8*��ln��s|������沀��C֎��n�BĄ��BS�ߛ�UC�9��t���8�{��<��� =�sE���~ݪ���&�)��G/E'H^���>�}��ڕ��N����n����c�O��U��X*�j
�[�y�W��˩��t�uEvKF���s�&�ro*������u�������V֎�n��p���������ii��YԈ�uP$cZsRռl_��+'j��g��P8z����*tG��z�Z�S��Aq���1!<��+ޙ����S�ݖ�{�Vn!_S�����"F@]eQ
v)̡��+�Ս����8��	�X^��u-\u�"�%��x]]'�\C�������4TE����شU�|��Tf���7V5d��)��`��䧄;��8�Q���s3�٩Ѷ��=C�N5���g�&���)5�j�����H�Zh]>��N��6�E�j�$��|������������Y�K�mwgt.��*��3��4�ۼ��u��Q���+�p.�v����m�Π�;�+���]�Zɍ��vV�&���(��2et+�������tN��ڶ]	�p;z8�S�4X (P����XS�8�H"c����uW%�25�.������!+��<<�Fع��.�5��Q�3zkMG H��Ω^�'҇(V��ϽZ��%���1��T��{��s�rV�Q�lн0�l73��1�����]f��x��D �ʀ�@V�a�<g�߮ȇ�L�8.�l1~������n
GK*��g'y�2�1"^�m�S�P���B�m�ӲGV��8�$踍/El�"�'����Z9�頪�"v&���5C��)vt�FE<�(;�t7�����}
^��:�Z�$;�:�>�9Q/*�8���ɣ���vf�yYԅ�%��܈WZ����ǸN�#}hdU	Ⱥ��e�)h�Ī��N���g>J�*��+@��ƨ2�(�Õ���\��G�����vl��%�vюE��𘽮f������G9��=����X�Ģ8;��uN���Wש/�-��|UT�m�OE�B,N�y�B�*�k�+��i�U�|�����9������y�uXk8�5��{i<����K&B�v%/�ۥBQ���7N*����3C�a��.ɫ���;Um��|���;�<Ӈ5�.�\��xk��ԛ��b�� �)�5�*���nV���s�tjY���"5��c���̾���;�K�9�<�(�^U��?a��Ę�U��>��.�[S�<0.�G���1꾮v�-}�ُtF��r�fy�7�t�3ض#+��j25�r�EM��}�+ cKM��ٝ�8��s�!߱֘+�(�OExS��n(�0�� `�N���6=נL�+uv��*ΰp,�j��U>��7V
��^tg})D�X����cu��x��'E�x�S}j�V)Zb�HL�(��9�g �!�>YsC���11�7"�ÂmQG�6�:���YҶX��b 9�|a]��}YPu���}ڜfWr��p�>t����d��d�`}����w 5��㳫��b���վ��n��;���J��tLs@r�-���♣�b�];o�}�q�}~n�*ʑ�Y��C���l ��<.TŶd6"�=U��R6~zs.�xpn�Vl�:*'%a����A`+�<2m�zͩ��U.Y�F�&���O�ph�l�'�r����4mv�Ui�W���uG:��l��T�q�9lʌhJq�E�ٶ���f�N���\�wjM;���3�'S���ɧ^�nLz�y;�c\�]���2���Tռ]�F/.k����zlãQA<��MG	�=�^�`�ai����م���aO����.�į1����^�5�,�V=1I+��N�N�R
m��x���iO�
�h#�'��w�P�Ň�j-uA��LEq�y�*m�nXC���1�΍��I�q8��]�é���ړ�{K[YBhk%:<�D��a��nc)JP�*ƺ��'Q�u�!D���[��M����KX=�5@^�/���L��$A]�}���	>1�P����q�a����ʞؘ�Y�:k����*�1���^V����Nh8@�dZجG(�9Y�$�>�sȧ�����VVI��$�7]��jXC�譕|�PU�/�2�o�Xu�R0�,��$��i г{u��p�w���q��Z����S��q��l�0y��dM��0j=�{�����mB��^�f9����\��Q~��6J;�G��,R,1%�lIX�X������\9$z�
�OT�
��Sq[ m�>�S���l;��P�T��{�}s�&��'�·t,�Ǧ�Ƴ�pN1ڱ޺����xVP�7��ԍ���^��nԃ=nN)ˣ��#��;�ى��	fhF�k��q���ՁG�̿��L�%�x,b��"/����_In��Xܤ��!�XT֑}֬��"m�7�s���p^����8eX�q�J��ng�V��]gwtM�=}-P�Ow��SV-�	4�U1�h�	n�^���Y�*5.��WUڭ}��yVM�	�5y�F>���p�u�1=��j�F��~f��-��b�� �t{�����&������ �ֶ�\7u�S~np�@�V_��W�����/������y��)g*�w[[m�_pj�`*�*��?+?�}��f��f�A�W�Ѡ)�W�
�i��oP ��Ǽ����6Eb�EQg��ڊ�^�[x1�y������^CU�eş[��Oi9��q)�A8���*g*�!#^�L�
;%1w�N�F�u���b&`��P�vb�|�e��uJ��( �O~fo��P�ǭ}- ���S��sꉂDְ����pn��WQ��4���e��4�M]Z��}�]��Y�;[sS�D�>�c���C�Y�XW�N�}\#DW����f�!�>�0�Q]Q�Ѱ�jؕ�*�Z@޻��G�X�qW��՛q�����p���R�Ҽv�x�.����ΏOJ���YNy�]1�j.�C��7u�y��/̠p��*�)�Dz�w�B�' C�$Nk��_9�ȉ��»Kʔ�[��Z�}�C|'b�ΜT�h���[XrbWR̾�e�Y��pػl����S�Y�����ؓ�W�f�vЕ[�
-�ޏDG��w�Is�	9���R��-b���}�,ள>���M�v�[������	j{K+��P��3�h�-����֡M��
~xm�u�
Q�M��Q�[)�0i�2S��ѷ^�`g�����s�xP��ޔ%z*�$|�v(-}V��D��Ҷ�V.��O:�p+2�f�h}w����f�[���;)�;G��T���΂��U��&���:�+P�w�z�UJ��%�9Qn�ECj�b-�W�����	�Ga�W�D��ߨ؅��"�U�B%�w7��cG�5|��1@�W� H��΢E71��
l/UX�q�s@��o&E��u�ר�M���L1�+u	��\�+[����5L�y����Lʤm�}���m|d��3��ٰ��דQ������C�����S:����x�ZWFZ�����Hy���h׶�ʒthvv)�J���ٮV?>�����7*��'�[B���.�5=�c�.�JF� ��{L��~��
/�+��aQwT*e[��]^��1D�zl�X_1���v�{�ד��E9;����ܖQ��^wq�-��BX�D����bi+���̙�a:bNQ��ڛ��6���k��ϒ��<��ʩ� 1@�s�vz���$��������´�G�*hou���t(�+�t�ھV���Ln+�T7<��p��o�	�n()���hm,��{Jcw �j�GܡO�~z���-�G� ��jK�Q����C��c\���>����e%�h'����Y��"�]S�����r7�6� 9*B�s�K�K��u�ɱ:O� �:4�`r�	����CHOwuc�����HEz�aL�r�8](<��*�;v�;o��z�Q}o̍���%�^���ȃ:};H]춦/:x`��s�֢n'&#c1�ŭ�i�7	,��Xq��hf���O�W��fm�F�u��qVqCx��=H1�S.�IT�Y�lh�^��8_����֘+�(�T�xS���0�� `����=����gtt�fo.�S�p0m����%hc9FC^��Bȇ41\a�WFx��e]]���d��&q����.����$��1���U�yN?��MI���i��d��-P1+8�a���ACL�2�g��։��:�?�i��E�I�� (��}��u�����!�n�8j����u����z}���4���M�̝��!�z֧����R��%g���=M"�\d���'Y���{`y�8��͟fAE ���ف�m�C�i�=d�<Ǣ@�����MS��R���3��iVb]q� �ΥA��!�zm7�����xt�-�	�����S�F������5��O�(�8n�q�E�]9���byv2�Mי�Vk���I޻����V܍w@�oH8/�H�ȹ��J�
�{���f���$�L!��RՓAì,�x`${:�t�a�E�P[���si�$c�=�I��uu�����aYb������oW+�����4R5kl\�fU�W�ͥ8"׷z⮞�EK��Xn:ۋ��ƙ�鐩-p��Yk�Q���R�ތR�[�WH��%���5h��Ī�	P�ij�V�9*�a'o�Cή R5�k��j�4;a�zu|3�l+�I5�0h���g>{-XAIC��D��^
�w<Û�ÿ��Zk�<����ՙ�f�oK9g��s����[�õ����m�������ٖ6�tCyݠ��>y���f����-P�H�$���'�j���b�)i5�pe0���F�o b�q&�[C����ͣ*KU������f�'��\Ճ��1�-5rޭj)��i� �����ky��f�7p�&EB�\2WH/n����L����ΩӸ9jn�\�*zr���3ӽ��ɘ���g����+iRt��|S}F���mXU�Fhc��f�ư.�t���`�e��bҭ��{�}J���R���i�l'QD�w��y�u�Ls@B�c���K� �!��5v
Ѫ�S9���4�<I�G3q��*���ضM$��_*̏��P�B�t���@ڽ�c�����kd�$��Զ��I}�J�&�*�Gpjݢ��f����Y�t��3:��iʠ��������Q�/k�`��-����ܬw�4[���6��Z��^l=}5a��iVi��Ңo]�� �Cc�𑻜Ean��b� Һ<��qi'��y6Y4Y�I��,�+)v�PS���n�[$_犣��Q��,E�Q��[�Tf���>��c�ʏWA��4�IӍ3[�SI��N�bZ���,�/0,�e�-g3ս��:E�aw����{��=���R�:��oK7oV�l{+E9:8鎱r��$�Y��վn���2�L�d����p�7�l ��F�]j��^8;��P�x�k]:uQ�:�w�;/V�I��Bpˣ±�S	�MZu1r�v�NԜ����]���\������A���Nu Z�i�*�cM^�vwf����;o]�����V9�-�s/m 71Yn��]2r� /wR�z5�,z�B��mB-�]�����K8K�8i�vAX��ݜ��r�浲H�ִ�
���E���w�f���T�Ai��A�$Ӗ��۹1����E��6흂�X}�wi�v��:p��M*�gGb��R�u��;��$n1"�B�.���;G^n�-N>��k5#��ۻӇ�j�:k7��)v􆥰��/BfA��q���tt_EXgq'w�_��_~�� �VF"	����"��,U��U�TA�E�iUb�D+UPA*�#X�(**1F+E,U��
*������Rڥ�V1��b�U�(����Q��DU)���"��"1Q��PRڅ��PPU[J)KE�Q)Z�Z�cc`���*�"2�U�#iV((Ķ�EJʑJ���kF#�(�Z�QA�*��J�V�`�Q�Qm�*�iQEV,���b��h �����`",Eb���Q��Um�eb(�H���(1X��� �"����+`��*�DUAQUPU��m�D�Z�E���#*"�**��UU��b�Z�U+mX�Q��m���TTDDb
��#amDEQEQT`�* ����m�Q���*�"��Q��d�Tc"TX��1�*��m�*Ĉ�"����PQ
ʊ*�QE��ł�D@X��UR����k/����Y��1R�w7��V��Ñ�w�ʗ��;sf��*�7�K��N%T,p�]0e��N�fLc{�����j�ژ��1-E�K����$G�I��1�@Qa��ُ��&$����RW�X�n�iXq�l?�g���0��a�H,�Or�bԂ�y7�$�u�Aq'���?;H,�=���sj��.����0����p���;C��0�$�b�����������g�L@QM�C�g<�b��4��~�Ԛ��0�°�~5L@�񒦧�u�EY8��L�����/�Y��'rq^J��}�b=B ���>h���Xc�{�=O_w�y�&��O��L�&8�_S��Z*A}@����0=jꇩ�q?0ĚJ�����=�i=B�x�����vB���ƫ�_f-k����#��DG����L����'�iE�dѾ}��OY*OP��;��6�Xy;��Ciԟ;t����Y�%q��K��CL��^'����6�A}aPré�4�-s��J����w�i$�g�#Ѥ���%x�QH,���0�g��d�2�ϙ18ϐ�ڐS�o��OXy����z��2m0�9Hw�d8¡�=s�>��%g̕�K�6��<����{��޿}}��[H,��SC�-H.�@��u�xγ��1�'SL8ʋ���i�|�L�@��N��s:°8�N}��s�o�& /�z�g��������7�?����?.��!���
J+�E�C�<O30�Ĩ�d٭d=eEY8����i
��̅x��1�<��d�u�A|�a�'5d�Qg�,�ͱ�#� w�b= !]����>=�����~�{Շ��1�ƽ�'��:�a�sT1
��'߳&�q
��y;���)+�a���I]3�%��b�>a��wg*O�q��ǌ
Ϗ)�'Y;��M��p�Ͻ��3u�vo�]��r\��c�=����:�u����Sh��y��D���&���g\Hn����f�R
h��6������c����8��,��R30��& (��������Nr4�,����=,E�zG���EC�+��;�p�T8��9�h���J����E ��y�E
Ũ�p��LgP\|�Y��Ă�|�0>M����j�3L<La��<�u���un�n�i���FlN���u��� �u�ڎz��7/#Mڔ�,�ރv��6ІH�L�1V;4�Y��4F�P*�O6�5N�Ї>��i����s�Ԭ�+]I��rVY��NڭK%�I���x����0��g-�S���{��7Y±bZ�F��= �y���	^0����ϙ�s�Ld���)=B����sf�*N�];7�t�>aXs�`~v���?e�UP>K�u��&�b�s�&ް+#�ǼP���}�E��y�B">���VO�C�T]��1�I��7�s�6�_Ry-1Xq�`{��JΧ��s�M"��Vi7�󻆒u
�Y�ؤ��q��{�x�c%�����6�iM^��o"k�x�� ��}��%I����m=d�ǌ
���'�N��{d�VJ��_����R1&���b)�m����u�C��dI-�C�wZ�@Q`=Ϟzw^y�ϟ�k�|�������g�Y�+1�!�ٞ�v���=��i���{��R�xɈ
l��z¾'1�n��i�+�����V���ԅf�+�i��Ag�6LE1jM�|{��.��2�Ժ�G����"��ٛ�b1 �>�4~a�~f�TP�ZE�����|.d�Av����f�^�����Y�����Ɍ4ʊM�Y�(~�f�~B���Y��a��������T�[�U�)����GDD��4��**ɣ�sFٌ�&!^}ܓ�ot�C��a��M&�$�{��~d̡�m������/�6�P�ֲ
���ɸ��@�Vq?0�����{�>=�7�}��\E�S���>a����<i�4�J����m�����s��O̕E������,�%I�}���zɧ�y��0��M2owO�lg̕�����*Ag�sO��]�K�Z�jNC��d�5L�Q�W��M\|`]�w�OŲzԆ��v~��M~��(V|��>�.�|�'������5����i8�Ɉ�0Xx¸�d�gh���1%�eOn���}[v�����C�">�}9?;����Ʃ�m�O֐\�~d�(u�P�$��N��Z'���a��eE9>�c4É�7/9�!����Û�����~��a�VN��ؠ�hnU����{G��Q��{�}��)*��7���<I�&���O��a�
��C�iP+3�&0�**����i��T�͞]=d�c�|-0��u�i$��'r��O�g��_~���Ͱ����DR�Qw�D�b��I:8�ioL�85a��mϫ&�U-í5�ǉ�J�$x����A��~z�̕�$��R.�\�m��<OV1sR]݋��\���� 8�p[�̕����Z�8 �@8���������3Dds��W[��"= {�{��'��Ă���d�VT��0�hq�%g��;l�A@�}9���>a�8�g�P�4�bÎ0�d4��Y����J�_D�'ug+g��߼5/��GkxU�[���",F{�|Hc���'<��׉�2W��{�>O=wXE�É��o�ɧ��{C���Z���üު6�Xn0��+8�;9f��!�%9����]�P�z�~�p�z�Cg��kt$��2n��z��'�0�������XO��M2~`z}C��,׹�>d>N[�'����ݟw��ni�j�U ���z0D�C���=#Г�Yǈm �!��u�E�aP7<��d�������4AI���v��6��T��h+��a�<��6���T
�ì�a�*��g9���}�oÝ�z����'�"G�{�G��3A{Dc��[Ͱ�����I�d�P�jϙ��͡������hbC���Ua��1>9�I��f�þ}�x�P6s���z�u�xxg�a�ϟ.�����53�o%5،�{��P��=���<iiY�>�0g*��`��O�g+�O?8�{I�0��1:��Ag�=-��O
l��zɷ�:����c����������u�������֤9�}���,��������CR|�7�m?3���^�����&3��!��?n��b�?��`c�Wy|���zc�G�TS���O3�b��O9��8�2y�N�}ɦz�QC���5���
��ڟ�_m�q���CL�La����Si���f�=z�$i�o�<Ax°�T6��Vs����=� �Ϡa��p��w�j�q�O̟$��g�c��0��1���Y6}�k�c%a���d?!Y�J��m�2i1�O�y�L6�������Af�9���|ͤbo51$G��#�N,a峉ο��$��H�V�!����@�Vn_9��H,6�&'^�bO��{M2m����/��V�ƳG>���2T��p4��11�H��M�S=q������"��1���5_\s�u#�j+��!���r��ޥ�h[Ԣ�%L���̲m	Hn����s��.�M`�!��Zͭ�������l:y���|�՛Mynq=QD�ލ�Zޚv��PK��Z������U��q񤫌�EP���I2��wǧ�=�{��y��u&����z$�#��D~��%�!����%x���S�����݆��g�Z����Ae@S��a�b�g�s'�m ����{�§��@��i ��L��{��������y�������쟑aP��z�XM$��C���04��0���WHzî~�*xn�ɦx§mԘ�̕8��1�A|`l��:Π������-f�u1�<�M"�YXs�}3Ϲ�;����u]�h�`B"Dz��{�="!t³s��O]�c+5��N��Rz��a�g�&$�
��
�=|@�=}a�6�)7�g���Y]���8�g�J������N&>����v�=����wn�:d���P�ZyGAg������$x��7�7'�E �{���8���c{a��Xc�l�a��@�W�O�@Qg��M3���$���d���x��1��_|�����O��~�g `�2T8�E�d�Y��bM�S�N󙷌
��<���8�:H,�?sy��\�d��ri�2Wz��w �0.��3�x��X~5a�Y��9�o�����wu��fV���K�s�= y�G�4y�4�\Mv�!��8�y>��I>x����������d�'�~5��{�|���T=C:`o�޶�2Vc
���g̕o���w�"�'vr͚��KVqH� ���=#Ҟ3h.3�'g��6é���u�E ����i���O���:�Ax¾g2O�l�2��9�I����L��LI�~;�m'P�] c��k�����sfy����������r�k	�u���v�EY<J�2zaI�+�'9O(a����t$~a�'5d�QHjo2m'�$�hc?Ns$�,
�:�y��l5�������z��y�����3I�@Qzs�'��u4��èm�^�O�Zq0�~��Y(�2T��&"Ͳw,���E&Щ��뷌
��{�:��뤂���1���>��{鵷D�[?+	�Ň�E�h��c�b>��Ф���ϼ�'����Y������&��E ��Sgs3�uH.V��1<gb��q ������Xue_S����*_�݂����R�7 A>֯�7nɺ7�Nq*}�^
�9�Up=92��i�u���,�l�oc5�t1pF�gv�s���\^��q��;H�,�4�m�|�1M����{aCh��{u��g��)� �X����N+��FKУ0�[9�"#��A���Ͷ�����y���;~a�>a�=�~�y���J�T���{ ��J���*Az����6��\gy?fu�Af0�g���|͢�Yw�sP������O�D �D���	�L��������!K����Y4���m=B��Y1'���I�+��'��g�8°��\O�y�Y�J���EY1+8���5<I��qI�~�u�Xm�嚴>��=BuO���j_t��o�O3��~���l���%eI��~C��jVx�|CL5'��u4Χ�1|���iY��|��P�M��f�;�o�d�30�Y�%Ԟ^f�YY>�_m�����gk�w�n����'R~B�Y�y������[ɴ����$?M�Z�2W�%�J�Y�J�O5�B�5��݇��m|=�<՜Aef�̂�Ag�3BǢ�D�D.��;4�v����������>�]���bi�0ǹ�ڐS���a4�����4��dğ�Ụ=a^��1<ݞ0����z����l=��;i�ɯu��� ���d�u�Aq&���~�z�w��ǿs>ϻ8��Y�:g�V���_�SL=M�����s	��Lf �|.`,Z��l�f��Y1E7�?!�s�&!���$�����rx����8�5L@�񒦳���νty���{}����3�U�IY��톒m
�ɳ�sG��
�_'9���|�H,~�I欚j)=;�L�&8�ɴ��i�����5`z�7�1�O�1&��@�Vq:��i������;����wi>B�q���Si�Xb!��u�����Y�q�|��<d�<B�鯹�����a��'䞿:@�}³�J�%򗙄1��+���>� ����V`U��{3�N�ؖ����i�ٿ٤��ΪJ��Ɉ�u�y�Co|�2~e�'�bq�!���Ƥ�o��OXxg;�m�=dĞ��̛C�/.�,�C�"$z�>t2�m�e��K&�f��{��앛d���?fM'֐Y�3XTP�R�큉�8��7�g�c7��a�TX5�É�>x�?g2�u���{�u�`q��k��8G�ޑ y�鞇�rzu|�bZNZ����_-ɪ��:��	]8C�Mvxd��rלּ�窼�'4��l�3x���Jew���d9:��O��}�Cݘ�so$�h�Ӽ����m�|�K!ǆ���|Y�Q����Q��7!en�PC����/ս�J6�GG,ۥ�X�6��E9��t��E��OL�������U}�}]P��xEZf�o����{���#�1DP�p��Ϭ�s2a���ᙇ�%@��&e����'��k�I6�z��,�W�
���5�'S����y� d3�H���	�t\�o�|��}o�������Ï�c��$�6���P�P*Vx�O~̛I�+'��q��J�C�14ɧ�
�8�Ն�Y�'ug*M���0Ǽ��=G��}��I߷�J��>O̟~�I�sL�%z�N}�$|�_;�B��H/���p��é�i'�7�N�$5lҰ����AL���X��x�!�~7I��~C��m�H�Dz.����;.F��'o��G�!%@QN3��OY1��B��%~哽���q�C�<s��4CL�%f￵O� ��y��E
Ũ�1��3�.>������Af>{�&�R�Wu����|d�^��D5e������c?3n��f'O��OV����1�u�6}q��Y�,�sf�*N�];�}�0��a�;���Ĩ�a�{�����K�>cޡ�C�]�ڲq}_,���Z'��N<`V����d�8���Y<�'�E����m'�ީ���A}H�Vv�0=���Ԭ�~a���a4��Y���y��I:�d����F�=�s����?}To�_?7�`~k1�E����IPY�l�d=ݟ2T�O;�OY=q����,1?2w�L�=�c+%}a����T���7n=a��R�`f�8�f��@#ф��W�zP��P��IIf������,�+1����9�i�c&'��w;�m��Y<5���& )��{�1�|N2c?�C���=��
¡��x��!Y�J�"ǢD|Lz �p��o�̵�FWG�'�?_��옊��'N�M`T�=C���^$�6��^��x����QC�icz�m��]$�?w3h/XT�Sɬ�z���d�n�E# #� �{���0}f����]g4��4³充:�*f���p6��TU�g��L�J��>�ot�Cӽ�o�&�n�xw�g�L�'�|.eH,�O�'r�����?�Ұ������0�����<ioSS�8{w9���� ���R�]���a��v^Ν��"��u���1�J�$c%��w�Ay��
[��N�nB^������J�:�%tz;A��"c�ꄯ�""==kn��f�����G�C��T%L��8�i>B����3OU�Cl�i�����ӽ�O̕E���'�ٶJ��w����4�v��y��z¦�7��ö3�J����#��̶�s��x&�e%?D`��4Ά�i�É��75q�����8�'�d���8�~��M��q��3�{� �a��}�5=a��X|�����7;�,8¸�}����\�w	�!{��-.=�!��8��VM0�¡��3'�~��0��i�O- ��2b(q�P�/�J�`T�8��N3�0=��6é�:ʊy��0�c�s\CI�=;a��+��T��U�|o!|�;�X������7�>egڲc<}��)*��7ߵ�x��*M'�����|¾j����T
��}�i�YURo�q4�Y*Lf�.����_->�Ͻ��E��']83�uW�gw,���d�Y7�3H�m'�u�T���$���&����1�{C��1+?'����h
(M��jx�0ĜB��1�J�}a��ΰ��hg(��(��n$�}�϶����e����\d��>d��f�����r��hc���N�~׉�2W�w����)����"�a��Y79��~`\���O���֤<���7��͠(��¾��"�`�y�l�`�{�b= |Èt����XcƳ��LO��cQa��8��y��|�C��៫�z����>��	�g�(2���V_<4��;��e���j"=�Qb�ģz�*�����u>�י��h�p��*�@�L�[;`>#�GA�3�^D���
Fg��^̤�����cO�0�9�m�L��}����W�TD�b'm�."����ؖ�:�Y�{r[0%T���zW]��� �Z�`���9�7��K�]9���dƗg�g^����;��w�`{/l��r�6x��	��Y��ͻ�o��ח d�-�����S��*��ܾ���Mr���a0]MZ����Mr�r��}�r��ޟ�Y���Yx�I����W{
�����{�j�S�^�w3t:��V�rz��T��5�d\;�F"����Y�.:9YgC8$Z����s<��N%�C�=�t�z
�%[3����NT!S�a9�I���l�\7m-J}8�U"�J��2*9PEF�Z�����r`�*\r���G:�*W���t+e:]M)���6"��!�|Bf׶l89D��Q"���\#@�p9�|
���]kg�7#�i
�.v��B����{�u
U����w�Q�j�TP[Z�"�/�q��kv�;���z�gՆ�v�V��7�6<2͊�����n
�%��K�ړGb#��}��Ld3xbE<�"zٯm3'���7ꝫDg��&�!���W�r���<�.[ϡVQO��U�F.�;���/h�44QO��\��mꃩ}�M�}�R8�1$#�A��!3�:l$�
=�^WZ�nx,{��#}hC��ˊ������x�M@r}�&)��7�!J�5X���Z-�G�FT�~tϗ�mj����76�ui��ε#������5��+S���E�[�a]�J�]y�r��6�,r7�d{��`�\�('�(�p��T}:�&Y��k7-�c\j�(ik�m�4r�繵��s#M�'����-���R������ܞ�PF��_z=����k[YC��}�Q0�gn
Yu�z1O���w�m�BமN���(�à�wS��4.s�˛%��x��(+�3�A�ع���n��!'
g���.M�S/F�_3���X�İ�9���":��#x�x��
�<�4Ư��V/{�
c�؝��-V��WSV�N5	]���;��q�c���S���0o�jqe��~���=���0Ŕ�Y�8�;�<,T*u/����q���W��o�=^��2/�o�K}��ZJΐ�n�Z�L�b}iת�G`0�a+C�2���BmU���b��Y3hm`��L��{�go^s�z�/Ry,TDC�6 ��ZʑX��!3Q�
���γpL����ѱ=�ށd��Ky�φ9Pe��?{�WL�b����_Ei���P+�Br�GMqs����������3�<M�p:kƼ�Y�:���S��bl.N��5��qj��任����n���G�#��6��0�F�`�>㒬�d��"6�Z�l�#^Ƞt�.j^�uy4?��I�LR1����uɎ��@�,�Q�r�+M�6�S:�m\(����I�I*�|�w[����M��tq��h8Ӿ�N��l��C�kit�Xa9���nԨvtx9΋t,�,<	7\����V��=߽����z�m��S>��^��u�����y2"��l��f�DT3�V�e},��%�޷���(1"ӇZ,;�+OIb3c��b��295hd5Y{]:#��
g��:{=�z�y&Tr�u���ۧ��Y�[0ځx|�,�q��5�vC�1I+��N�N�R
c��Q��:� ���P:#A�'JPj-*�^�LEq�y*m��B̡�r��u���][��k0�M`�f��F��� �ZV>�ꖧ�( �����R�=�PI���y��ݬ$�3}1�L-<��&�L���[�@�fM�[U�9B���V�^%�p��w#��}��ܰ�.1��I��s6��.UQ��ߨՖ�c'6�o�9�a�t��l.	�>\y���Bw�è�jX]��:�Tܰ\<���MVk�A����p��rf�y먶j#*P��3��4,�U�{\6�F�h��T�5+WwUԜ�ի�3&��J��bl��g�-�m�0���,<7�,M��Q��|#F(9{�J6
�����8�sus{6f�0���t���xhk��3up\���ug���2O���!���Ul�q��4^i�]�͆��)K�$KBu"��ZJ�dS�2XR^���Q\��9�y����f�MOR��v6�ا]g�a��ëX��SK+;�VGƲ������C��)m�j�{x��M��3�o�\�xd�U3��.I�m�T�t�����3{�3��c��YC^pؕ�i���R��'�An�;>��]X�8�a��w�1�u�JZeɞ�:Zc*�;�KQlq�U�S2��*��G�R�m�q�fk��q�o.5�������4rwq_
{g.��[x��Fh%`î,���ʗDǔ��������/N,�F;ݘ�O�rQ�9B�!��b��2奔h�0gR�y/�u8�`�*þf�Ae
l��N�Β̙���M^�T�eb!�v�823vei��G���˼6���C7CVݽfS˵Ȗ%ZeK���_ �����kp)w�ޕϋ���9#σǕ|�qf����"�͋���0ON�wsr���ԗPN�3�Үn7-`�IY�R���y�t��@a�,C).t,����f�t�Q٤ga�XT�Μ��$Ȗnɽ�;M�}+]r����|������<!�[ۗ�V�O\9�ֽ��qYG:oh�Oīg mu�,-� t������t�mҴ;/[��ڿ���(�Y�ɞS,�)�/y��'N�.��!��u�Y�
FY ��*c�|�N�u�X8�駽�"Z��1�NT,g%�:7�TtHPk�iե����1�0�Fhr�����@a�M�U��ԧ�:	���T=u����k$�AM����*zc��3�ug^��[�Нqr�Sy8`��g	�����Y��-qKO��l����n匷ݔv��e�,g5���AnT����#q`0r�c�v�@�F�3w�6�o*�ܪ��Ŋ=fl�9�lM��XD쯟=����r�)a�©a0�;�{Y��
+���� ���m�(��n��z1uw ����/�"�N����W�$)P�BJP���w����і���|��xv�b��AJ�&]<�yIQn��tn3ZB��Q�JX3@٣&s��{��Nˠ�BP�Ȋ4`���Lw�q)Y���1���p'zq����{�ơ�gF[r|4�K��ۺر<��zjV��Zp"A�P):~��讷���e0���&������x�ݻ����`�����lوM�mnt�7p�A:��
���S1�*�T�ۘٺNѤj�uj�iŋB�
�mo�j7��-�.�%U�P嶅8+Fv�����O-���|��2���z���ſC(m5ͷ��wLQirA��hHh�Ra ���̘
�`���Ywy4�F�+�웚���-Ս,ƚ�%y���N�5�n��yq����i�Ė$G0��إO:Ǯ�A��.��ȫf%N�P���^B�YDDUT�,�TB��TEPX�,b�
�T2-b�m�Ub�Q��F	R�Q� �1�QF1F,T�kl*�X�U�����U���F+-(��Eb(*1PdQEX(���YQ`�1F$Ub��cYA* ����EU�,T�X��"��b��TX���"�[PAT*T�cP��
��)TU�Q�U���Ŋ*�PDAE`�*(�F1TA�0FDE��T#�h"
*$�Tb�**��mQX�
�""�*��cUV1�`��TF1TV���DUb1`��UAU�"��������bFDDE�QEV1TE*��E1V1QQ1XȊ�QG� ��Ӛ�NM<.`�%��*�.Mw�®G��>�sls�F�@��.�7rL�q]L��D���bS۽��=���".�����݉���]s�F��e�*����ۺ�,dTjt�8#+���m�2���[+a;]
��`�hČ��L��$��*�A��'#ު����pt�;�����*��!��=�ylG?������6��YH�w�S�^.�0��r��:㷂��MrȹX���`Og��^�t�^���RA���m�l�ߛ�'��"'9Q����U�T��Y��/��.�B���.���Ss����п=��5p�`3�`��5
���I����_!UO�E��V�6e�^��\F����:'n�%�K������s��}O�Ȱd�f�"U�\:����� �",�j��!#qYb8I��f�����wv�����Nک�,@_L j��p�֓�+$ŏ\Z��C�=G'n�h�f^(W[|��7��N�F�(V����k�'�j1�vTFk3�@֔�����A�����+w��H�B�Z/ѫ)#y�l}�s�C�����Z0��o�3lX����U����=�8�Z���5�^]��H��mz�y#u��V�AS2�ͽ�l�ݩ�T�N*߸�n�
�r��y��<�,D�09��;%�*2t(�SƳ��ǑΆ�_���*�}�YS6�������o��\�R�r:�ɀ%[�oGV�&�{�T�Y������^�/+������]�LK�����ã��cT)ѣ��
��֎�n��P75����o�s�^RE�o�Huk�V�C�֊�4꨼sw�gBy�<��}HW�Zdr\�T1+C�ʹy��7d�/�xn��Ƈ-͵�b�r�mA�c{�u�2���j2(-TA�ѝ+��=ݩ҆@vL|U,����B�Po
���Q�r��yR��E	��H߸i�+�sE��jZ��P=�NLPK0zD��j���Ϊ���_���{Uo^	Ɔ����%<!ܹ�b��E�8T�*���*�3S�U�b=���r�zw�+c��0b�T��<�; DW*�L�c`���/A�����H�S�8��ճ��*��f�c�����/�X��ӵ)���@�	��H���0�T�`�����A�Q�f������1�i��;��Pc�R�
r����Ѹ$����k�j�D��[����Ҩ,�Qӓ��6f60��Xf/pV�4�M��-�bm�w��D�fa�W��gy�0�<hĶ�g�kx5C�eӺ�wnd�����#%�)��\( �R�K��5���!x29�Z{V<�Zk�Zd�3���.�Cq:ɽZ�wi�.3��ᘵT9��۸��r�,���<Aa~���������r�sJ0O��|&5+Zc�1"�m=p�{X'�����v��t0�p6�_^�c���}��ߞ⁩�n��p�ޏ\7y{E���)����R�3-(��KX�u�����kS�=Čf�	�q�a^�r,pk�6�������/3��3m�ՋDGh����X2n��}I+�p��J�ڮW���Z�|uA��ʦ�m��
�)��-�\��¹��\E�.���R]�S5�|&���!�WW��μ5G��ø�^}ƻ�n.!�������DTq��3�
�bE���4:���^)B(M�ɛ��fa��d�vo�!����gO�1])7�N�q~$r&��.O�ï.�{K;3 Z�������َӢ�w:\Cw�)����\��>P��`�Ün*���x�Sk�h	WJ���q�Lƣ��JF;�3�煊T�8Zs�!�c�0U�PQ���
�\�I�7�sɵ(J�.(�0�r��IϦ�g 0�a�Cȣ!��|B�������%KW�1ow���!�;_2f-Yqe��\|]U�w��娜��;T�Oc3CV�F�g1�[#�*�-;"r�J,�D2��X�b��.�uo;+x7
�֧�ȏ��Ԏ�*[30�ޏ�33��Iw�8�V��vC�,��֚q�nVM�\��W�_C�qա`z���ȇ*������Fڹ9U���ځ��Y�z#���	c�Oy��<K����K@g�r�d����f/�$&kܐ�䱝JI��[r.e0��<�"��k�Յ�Gi�3<�d1d*�:|�^�1���ڛ�����ߞX��-���ٖ]��>��~γ%�gC�q���{gEײX����9��]u��j{�={6H��]{��mIہb��v"��9&��˅-^i�b��p����:�r�߭B�{Q�=�40Ts�! �}��!'�q�:�dE<�&y����à����x1��uvn.�Y~!������X�]>S�L�V�{�Z�j.�Z��z�j�����pb��v�}s�-��Yn�7겇ݔL����<X�BJ�U�8Α/*t��'5�+���͌��������1p"`�AH�طLEi�<�ASl̷Z�Y��Dte����Ѓ���?K�+V{�LG�����,
�}
�!�A>�M�Ue�-���!��TM�cEiWy\,�0��p�Ӓ��8���G*�+���d���b�3��K"m��e�S"O����n���֍�/LZ��f�H�����	ǜ&�`��#�5�x�ӆ�k�vD*��1�ث�y�Z�u��7����̛�%9��ĝ«nC;n����x<���ϣ吐B���P�-��r�q�ПssJe§D8ALE�D�[����ڕ73���6�޺C6��ub'�JG��ԅ���è�j��W��@����&��42i���p=u�ϗ������"L��S��CE����'���O�.�[E/�	��(z�9$g�ޚ:�a���ץ:��
��_�5ݔoiW�Iq�[�a6:�er��!��d
|�(ϹzN�~w[���9�oH1���[>�}�k��V�k��^�֮U^��4f}��@(�4���#)�X
�ND��[3��M"٢qILƃ7!+ܧᕗｹ.�(� 'q	���7{r<�'_���0ł0;2�s7�ʍ]�r�x�T �N`zWn*&��ǧ{�!<��Gɯx�th"����3]z��d�O�iKd+�s0��@��fUz�Cs��/P�>�ǃ�yX��o�1+�ovr�(�ˋw�n���g����rJ#,'�)3s�g����y�=�\���~j���o��r��V���x��A�o)��0w��W�͞����<f�1��֞j����B�V��QC���C9�<iE⭕Vw�ܚp�2���Y�t�z�6Z�����2������_v9|� �-o��Z]�wN���&�z��L�)�������:�=��KӋa�c�m��༓�Ѳ�m��I�ժ����U�;� %Ҫ2+K�˵R�(���LYJ���j2���1��8�â��z|>�S�����QuR1�*��H˽���G�#�)�m׮���j�Q�z����n��������{ 
����	ޮ}x&aW)��)#y�l}�s�C�>�����0!Jg�Ō����l~���Q��@m\��&���e�*q�0ƫ������Z;�wr����b-�y|�u�B`?Flț(tQ��Qz�.��!zt&���7���,�vd"23!��v�=�{�� TstDGq@�a�²*hcs�m�ɿ��B��%�g�_�Z��2G�Z��!O/o����bPRG(f|�;9g��FY�:��0�Sj
�|�l����\}��u��׫�$x�W��M@�d��K0z�F����s,>ò�n�E����'qi�)-�C	Ow.j�s�L�SD��ؒ5���[ň�9�=15��&'\_���ř@{9Ͳ�\�\"X�����oi�vuz�[ ����g;̌;��"���	���\jdI<����3��c�ʢ�o��'���[hmJ���S���(��#�'�A�Ժ��
��tP;!�`�D$�z#���a)r�5�ȸ��\�`�s"����%�@b��Y}w�^�#9��y�f�f�W���3��u�Ft�7�6!��`b�1N̦j�tXp9F.u2;��T]";"^��J{c$�0;PI���5�ʤ�@�L{��}颐�xk�b��H�)p�#�P�K�<�K`�d��5�PD��`����	㘖q�)��UY�\쪜'ʆ���GLf
�yV���B���\�3���/���׃�HzZ#ד��(��/YXZ"&��k�����Jos(��~���l�頪�~T�G������c��%7�E��׈�6t�V���J��k�ٰ��W1�C�&sMqiZ/�k�Ue�,W��3�fZ{VU`�|��Zз�ϸSF��g�� �{��ڶ�z��PU�����t;�b�V��:��o�݂0O%��=�
���bY�b���v8�0��]\�WS�C����8�\s�^x�����I�p8J#�A0}a#-qsC����b�<d��˜Ӯj��[��r�.�m�z��wCB�<Ccb��ar��C��뵯pD�U`�]CR����Q����t0�+f�6ɾOn
r��������S�q|𼏙�u =�
�;��8��4��lT���UG���q�K�M��������x���7ʰL��:�������*�%˒2G"p��R��p�p���U*%r����B���S�<0Z�������1ѯ(���^1^s��M"�@��X�ݺ�Eys�U�&:(�.;��̂�����p��@�x�Lq��`�)�B�-��;���j�+�F�㞢0ïNP)9��hVr�[V�3 �6���(��^Ks/Jԋ������3��ץ)T�ئ�g�e�(��h?�˰��x��Py�ޞ�5_f�q wE4����]{=5e��؍�>Qr����?{�V�f��='?���V+�W�Lh�/=��n���N3�]��=�>�fu�3���gˈ��lT���ˈ�?��y��e��_	CA
����ʃ�y�{՗Vw�ޘp#F�2`�h,�-M`�.��̰Ov��9=c�bj�[�"�Dk�!<d<Iނ{���i
~�	[<]`��Q�M)WX��[�����JB<N��u39�tPueq��#n:|���9>�	����r�׫��pi,v��B�wZ7`uBH��=��x��sd��=y��jKWr�(�'�A��ӯS�x�]f�XC�pE��i�s�tP/�t�j詼m�JpDi^�A�����D>�ƭF6����)ۺk;n}Ъ�ˉ�у�Ab�MLy?W�W�W9d���� ���o���O�/ZoTBU���p-+a�8�J��)ΎRZs��F�3��k��+GR�/ϭ�r	)�7fb�{CPr�+�nX��2��b�qs5#-Mj���-��8��R��>0���;�Q�� n �LΏ x�xP@�����
yU��h�}�ꖴ��Nk�]�P�i�V�ÝBNcB��ӓ~U0����I�����V+�W�%��!$[{��wg�3�.�}=�\�8W��^��˛R��s5ϡ��36cOv�V�嶂�!g'�4"��G��#�F���/�Q��1h�<!f�lT��n-:�V@3't9�ۧl*Nt}�x*R*��:�-]�>�U�i�l��a�R�y���Su=��tƏ!W*�W�0t�=5#�9)�d�w`�s�+���V1c������Ȣ���Dw�ϕzN�|u��[A{��� �}�<Q(b-zcq����9ϹlR��~WM��`lly����N�*hA�3��ȫ��Jw�R�|�%��w-���F�8�ved�\��V�8�yI#��Z��.�,�7UЛ�Y����,(��L�wh�a�޸�\�,ֻbWVoe.���^���u�ۭCkQ;��Q���+�2�=�q���P��G�{��yu>���\�Ā���*6���g���9����ȋI:�t�\��/���k�n,�M~�X:��Ǖ�izdu9p����DX��P�S����7�n�=%���o�n���4x���3f�^W�]�Xp(UA�npz�sۡ�Q�{�weV2Ԛ�k�V�U�l��$Tf��F��+���vW��=CnUc���[^
��'�-K�iu�ڦ7�����B�Ή�'�s9Zy�YdX�Bc?DL���b�i���䱮�ZlC�:j51w)�h��uä��.Y���iឪ@pc�қ���t��k���|xA	��#l�6���Lg+��[�R2�!תa�(3w���W\KL�1ǋf��P�<l+�<}M����+!Ճ��P��醙j�e.�vd����
;�!��朞�2\W�	�_��_\D�hX�Gl��*��`,p��f㰪tl��,��^�Z�/)�ʫX���z�6�+YA3��Z\�u%_�p�pw��:��x�n���d�� ����t
+��-`j�K3�7���5���W�����
}6�d�¶ެ�ǪvN�����5N�u)�8�w�P�֡P��8N�k���# ��e�ɾ���=����}�#uv[�]�fq��SMk��x�<d^+ռ��r}|��pK�ueMK{5�r�a73'PsP�XH+�cK9C������Ewh��� �#�ل�w���4���l�RX%��G�ն�TU+0Iwķ���Vv	�p�E#�\�Tb�Z~�[Ň�&*v���eb3��IID�ƚ���I�r����
�j�7��[y[��lz�!u�N5�����i�m��˙�+�(��)pԶ���V� Z���{�{X7]֏�A�5�ɮ��FHwjޠ��^���*��N�g^���t.��%8μ�Z Cʒ�M($EI]�}WJ����չp���U'2�F���A�.������54�yHm7A��)1�$�@��Vms7j�H��L���;��1�8�"n�J����-�Q����p���	X�V7���87��4u9��LK\Bqr�)]D�Ùs����S
ꎤ�vs3�]hu�9��К��&w��@�>��)�ΐI��
��u�9�[���ɲ��|!6���H��I�َl`a�㲜=+{V�9�{o�����[6�Aj��8fr����(]�5���F�u�!��
��#Is��<����W0�3�U'U���oD҆ە����VN�](>큙�j�X��1�c��ɕ�xx��N�~d'��rpX��[U��U�7d��b�+J]a�Q��5��=��m����������M3�S'��t3��8>	�x.]�Q�ݼ̖&���I"�M�++�&�|��X��j�h�H��E�y��S5�x�ֳ[��N��ʺxK�������A���ڇ��nЌ0��N����l	�}L�Q�[w���5��Msʴ��$���,8qʼ��1���N��*A�'�r�	x7n�K��-��8�{�v�۲���]%*3���F�6n�S���s�fD%H����d-�����#�-�@V��qY��*p��e,�X���cf� 97�e��i0���L�Ʌ� �Q�(𿕹�@	�܌#z����qU��]!D���u��N�t{�U�v:=�zR�t��:�*��8�R��+eDxn|��<�9�YYut� N�;�ֱ�Aec|J�
Z����x��㚑���F�o3A$���rШ��n`��ta �shXc/6�Ov���}�P��j]�i~�)��EH��fQ�f��
�Mk�I���"(���0b�UMZ"*0Db�UX"��U�
��Tb"ZUKJ,Q���b���EQUV�dATX�Ab�E"�
1YPAF,`�b�EU��DAF
���A"�"����b*��b1�#�U�0kE���*�
��b"�֤��e�`�mDdUX(�E�m,U��DB��QUX��Q�*�6�EDT�Q"*�IUb��Fڪ"�"�(�TUF2�� �ЬQTb�J�b����AH�V*(��"�*"
����
+l��"��(���*+�U(%�b�@��E��Fګ�1E"(�"�@E��Q��F�5*�[(ȫ��*�-��F �*�(Ŋ�FV�jc͙��G�T4�72��`߲�����#)[�gb�`�k�[�ױ��f=���Y��MZb)J���u�g��u���G���TZx$��-*����h�.������6�T⁬3�VT���,�WO�كj|��O<59c��dd��j��]^���K�W��![3C��P��|̳ұA揓�5g�:�����MSp���B7
F:���'�s����v�=��Y�E���M�To�e�,�#�;;Z�XI� ��)�z��`2���;�5[�Ⱥg ��S�Y�۰�F��OY�T��ĿMmƂ$P羟h6��W����"9HF�9������� a���\��׊�αQ\x�����⍈Y�a����cjS44Pp9@��يx�r�t)V(�T�Hz��Z9>�8}tc|���c*M�6+�((u��6.�=k7��ll�˃q��ɧ�^2j�\aX��7䳍�O�خ�w
��������y{n5��q�(ϕ󿄮�5>�i��B�^/�~(��'��=��e�S�gi�x1Qy0Ƌ�r�_M^�l�ߕ;���.t� �qx8d�����{�wtrtF��s9�y��$�&�i��yU��^��C���k�'��}s�L�9,�$^��� �Z�s3�[Km�D���ۊwO:�h;��^o1�&g�P�܃� ��[II]"O[j�xfne�[d�\bUY�Z�t�yuC�� <1� rG�C�B��l�q�q#��a3�h-��i�Tn)с��J���4�c<�V�#�l��T#}hd��
���b��5M�Y^T��kԭ֡��:���.�&I�����3���>�%�)�
�j��K&%����U��a
��[5�kƈ"S\��o.��}v.h�����%K��vp8R"������ �Em����-�c��Q�0/��"��.F��aH��-u!QUu_�U)7�N�p �N��L�Nڬ�"�*C��<罞� w�`o�%1y��¹������1������u71��Hu	1|��5���]A�G�|�j:3�vS=Ǚ�CE���^7B��<�.�I/R.u��5�ʦ��9>��3�FU������Xx�!l�Q��oe�{��6c�z�F�n�~�L�t:��N� IL�a�eH��9�b��6�O(w���ܭ����PB���}]XYGi���糔l`���j�\��w�ҙ��$�b8*�J��b��{U�o�M�؞�=o.gJ�R���	f�Ht��p_mJ��r;�8�$;2b)O� k��f��������q	B�jЭ�}k��+9wV��&a��5�J�ci:ٽT��сI��$������g�TˎsH6%�Ӎk�Țxc�:*��-^���Wo0T���9�C1}����%7�QDhPO���g2&��|r�#���2�ڼ�].��~�	����7)�����y�{7SG!��&�:6��<|�K�NDVҥ礛�n�{[
���b��cBì���Vk�Ӽ�^I���y2!�g��3��(�����ϕ��<!��n�b�y:�ev��xVJ��>��k��A~�b�
��̫�}��-�k�G u��+�[����P�~�����y1��H�q���c�W`,d5�+#9���NQ<�� x�8R�n��\���5I\rǗfU��j��m��nOqp\�7�\:t�Óc$�G%G9�+~'h���-jc̏G�{#�ݱ�}R�6�Ǝ��s
���'!���w�e�U0.�k3�5y�*����;Ia[.��k(r��|�֫��|P�-�nXb�.1±�^��7V�n:!�s�c��˖��n�ղ."WDޗ�RȚ`�GՎu4&�u�v���ϠT����lݞy�I���w\����pk����]yA�9J}ov�g5[YXR�vx��W�5��s��W��#1�R��>�x�|ӎ�kl'kO��5��va��.��','�>�'��b���ވ�el%���˃�ab��-�Faׂ�*뎧�G�qw�i��&81���Pv�
t��L��ڛ�a�wm���!�*�W�0t�=Daw[�ܴ;��*�/��#���tҟjD6_��X��c|�+ R�n�j���X�I����=��d�:�G�V�x�/����;��V�u�0s���sp���3>�f6f���;~eU��1�����<�[0�:랉x�t�u��ӟmD
i��s{F.��~I:����F�Pj��Е�}a�R��(S"���^҃���N�x}�9�,^���׷��/�b�޷�~���哃��Z^���RUк�XafO�g�ӬE�T�C���[�BXǲ���{��X��V��P��y-,�uJ �5�՞:h�j���9UX'��&����³�'wVVA�#*���Y�{[�	���`[8�<m�ۤ�WA
�D+�>��q1��	P�S�^Cx�5���Jb�u1Cuä�M ^x�>��N��Pdb|ǲ�z�������E�����\�Ivˑ��k��S��
۽ػ�tX�����s�3 łVn�X�L��.���+@.��ΒU�d_����S.3��S!2l�)�K��[|_u��>ӿ9��r5������*���\��:���ݎX����,��Km.�~��KG����ͣl��հ��7!]@�ܪ���u�q�&)�w��]�����sSq��[4C��N����\V�c�$�Ͼ���F$���$_C��6����]�s���(?9Q^�A5+�*��8�9�v��@,pn6���N�'!�'�X���P+��=���S.���g*sʸw������s�T�g�y��ۂ}���ð�X������ ������3ڽZFh�	�V��$�5}��rٞ��}~�����RB�f���o
�!��nfr*��"r�jjb�'Jl��@肞Z���h�S�_���t<���z=Tk8ȟ(��s��&��T�Faq�˯d�����py����#�z\�1p��]3�*h��Fj��T�ѫz���5�LI���hXO'��In^�(��T^Np19�B�Π��a�b�	�zK�������)Q��|���n����[���a�c^�s�Lz���<Y�|T��k�����avLIv�/9�W%V!5$�T�sb�>��e�4�\�3��Q_	5��Dzߒ���7�^+�^��9�o�c�!%�Ȩ
��s\���=�c��eX���;�R֮�3�ZEs�L��r��N�m�g�3.�����"�Y�F͸��e���F��;�t���8}���5�ʤ�@�=Ƨ�S��:�l�Ҋ�j]��Չ��S�ʒ#B���5��ʶ<~��l��$��llV͆	G�[������B9񘺌�PW�̫u�Q)���yQ"�m<��u�8tl����1�sϷ�w�Ǉ�VM�7�Cy0Ƌ���_�h*�l�ڧz=~n���3 ۋUw�rK~ԟ?�s�h�m_�b��y����.W+юa
��	��Am�h`�/UF�.��h`f�k|��i�U_%�9�C�(f��:����59 �(]����+�*�^aA렦���*H|7F�:��A�k�Y�\��8J�Z)��hW:K%�D�>�X���ϖ�צ���;�cFM�Z�A�1��� s�TcT��wZ<��GGϼW�t�HN="cv[�莛|,��'[MD��kTL��RS�Y�)���1�u!P�T��*�'�:!Œ9^�:!�k�_:�#O&&_c���.���S�b��yʯzy�r��F���O�s��/m�TT�9[�
��r�e��%��]�v��F������A֊>�r\��-��Vr�{�����wvVUZ#����U����;��j<�'ɧ�ͦ��-��X���n�)龴���7�e��`�RL���(�ry�`^���UTn��=ǀ�(~�A�ת����G@ҙ���tP�Cb5[�C��M��9
6���Ej�Y;�z�N::e5���qߍ�,�;@X_N��D
���˄�f7�U���w5��Jj�w+�>sD��9Ewv�X����Z��Q�^�nj�nZ=`pɬ���ܗ��/v&þSZ��pCȀ~�_�^pu���O�{�V�,K {llg�f�V�ݮ��P�����͹P:C\g�ߒ��(�Cگ�Ϲ�����s�9����,���S�K,K�B�L8p�"7������D7��^�x�Xv�"ϳ9� �;��J]$��rz��J�8)w��`�|��t�u��ݨ���-rMȘ�sy��S83a �-+J��Fc>#���Xn�PN��F� �=%�[>SI�:�(5x�y��^X߽�y�X������/E�
>kiꃨX��;����.�N���*N�:�X����=[ʽ�Un�p��+}h: �(�3���;�y�����fKˡ�r�)�� �G.�Y������-\�7!�p���!4wd�{�zK�ϕD����)�Eې��=�WO��~�&>}�jׅ���r=E��2is�Gz޾�Op3���kݏ�3�]�}$�	�U�)D.������y����]�?@8R7��h���N��d��;�Q��pOAQ��,��k�=і��wytf�L�`���7�Ra
ң\��w�{O?cH�&�Z[����q٪�ꄎ���pB��9��B��+�)�,0���1��niL�M�ǣ ���1o3�gC���1�Xy֮$YhȎ;(z��u4'o/�QmK"p�a��ݥ*�|�����*�b;|�
�7|�î�JEC}q��#��<���)�ɫP�����v���o36�oEرR�)-V�ٍBʒ����i��9�0芌�j!9�Z:�T������[�P�<�P���b��d
Y���a�-�;��9�,L
}3�Ыy��T�)�ܹ &����} �sp�M�q����Lf�M��UX�#Q��,�
�Zɝ�y�<�-@ؼ3F�� mڬE#j P3H�Bs{F.��a	'Y6�㠗'A�?oM�r�z���bR9C����;{�Ď� Nl���DP����MecΖ���+��$5�wb��g!�/�#5o��{16��y��et�!õʥ�U��cm+tYJ�� ���Bc���n3��^�y�$���������/5�΂�k��S��+�$�v)�7�ܳ�ݙkFY|�7��n�ǘ�[��-��U��K���g�7aZW�3
�����%]<:�|��Nu�h�
�!U6O��\o�µ��;o�;yv���721+r�"�����y-�FX�q�7>�4g�ղ�[W�Ä곙{���	�����m�l���j��݉9h������MZ�X ލ�2�W���C���S��%H�58�5�i=�������N�F�Cuä���3Z9zx[{��NZW���^�:=F�h7��D		���6�Cn�v��7�i4ڢ7^�Xͦ]�����>ԲE{\d�,5euPxam�H\u�����O!���d� �4��Xފ�K�rTH�,�i��?(+ڕ�&Kξ�����aj�
�pU��Z��ؼ��$��uSj�BзMhI͓�P+�2��}"+Z`j�r��X����!���lK�ob�D�]HJ���e��J�҄�Y�z@�m����v�ة���E�Gg�p����[�{O��[�p���i��cUmy�{S��ɀ��U���"��7
j;�s㼊Qӣ�f��y��:��T�[��j�kTW��$*�%�cq�;KkY�{Ii%xg&M�wذ̫ҡ�H�8^��*�S�}]�	�+)m��`�i���nVU���+�3�q*9�[�����Ľe\E�m�Mi���:Ս�ۗ�wj�W�1o �-֯ �+�4N�p��ܖ�Z��uqI�v��S0"y=�n�E�#sve�Ս+D��!��g���(��L���tA���I�a�ynT~9�S����D��j9���{xM��d�i_t��4��\.�Pw��Dh�Y6+�=��ʀb(D�S���N�P�]U�x�<����p�}U3��6"�M�4,>�)�7A�w��}GV>��n�D�q"ᘼ>�����<F���,{�X���WS�M�=�=��	~���� �cy�����-��^j`w ΍�bn �|���G�S�e�'�zI�VHA����d�q�gb���'y�3���LPzpO1>�����.�<�LwwZ��M�x8���t�#}:�0�
ږ�磦����]�*w����/h�չL��(��n���/f�!p�6�H.�q����p"��a
�	��ARU���>�<5��WppF�^WnN��^�p��U���Z�6p(���AU=ڃPӴ-\���bj4��8�Y̾81`���Y����w)e��·�����5�����Sk�jjf���B��:�Wv��j��S#ڄqQ]3{�ғĲm��+�A�P�b��puc��������d�;�|�M�7�i+]f��;l���uc�����ʻz��:vIQ45��3�PG�[�X.z�C�F�`�Cz
����`]�R퍐��BnS��04�|.'9��Ӛ�#�u���V���ࠖP�&&�GN�eZ�8�D[��2r۹�����2��	1D�ַ�XoB�ZwB��\�̾�G����u[���da��#�KvmtR6�R�9`%���{n���*o ���VgV�S��7+����
x�%tt��b���]��atm�8=�����D����y��ە�"D���.6��2 �LE,�Ŝ2��'8�.F��ݥ�ͬ#:7�=���|$� /���H�Yݬz��i�ջ|��;��B����e�������e���IԳ�U�֙GV�1d�$Ȅ�����B0%����O34��G\&N�y�i��k��YB���y�CE�P�}�w������������8�rK.R��+]@چ)�48e��
ڒW.u��܈���wyZԫ��O;5^�1����K*Un����7�%fÖ5�Bn����b���}tĿ�FrL��N��j]�{MÏ.�t���b�xû�qM��	�H�0\��{$��L
��F�Y��UMR�;��cl�:n�XA�[v.⾲�}!;1l��ܘ򻄇�d�l޴�!�H
��a�T�z�G�'�]X�˃5�7��tv�NҰ�Gu��S&�0�`f9��`;^T��:���0ʁH�1%�������Ɇv���@��-�op�Q�ń��KmP��7\9�3n���m��t&ܦ���ʰ�Vn��F�����ک�=kC.�BJ��-�\�bL,�֗��F;բ���x���cl��A�"+eI�H��F�{N��~۽�J�Vz��H�����%����+l>[p&.���Q�+di��OdY�3�����d}�@�4�.�zRYY��]����[@��ż�-�fWj��cI�����w�;x
��f�Qv�z��o��<n�]��b�k�A4u�ը�Aҙ/����p��PĲS��V��l��RV�� ���DEGn0x�Vś{����9��sR��tC����TQT�v+}x���l.��������`2��sDL��-�4��n�m�1�&+��u����6��h��6����ٙ�����0���7d��{t�=� ��i.��zqѽ�+�$�hKi�z��;s��M��N�we1��KdWB�F0(�2�Q
pob��L��ƧV�G�3p�Qn	�Fp�*�-�ֱs��pet�eF�]�
��Xl��"��]�0< I�F��Nݨ���W=u�4C���ݝ{���˫V�ɡSP��P��9$;��	 虺���0�T�Ԏ��f9wk�.YN�@ �G�A>>Eh��A�J*�+AV,EUA
��T���X*�"�U��Ue���(�(����(*�Ҋ��`�l��e`�dEX�UQ[h��%aYm���PTF(��

**�YR��UAb��E��UAX",X���R$ADEQH�,V*��V,�������A�H�QUE�[j�����(�0PDAU���H�F�
���TAbՊ(�֪�)mX�Z�UTR
��*�U1A���� ��,�Q�1TkQQ��TDX���D�IR�k+T�e֌e�ɍ������}ϳ�[6�s�v��Y�N�{�������d�{�p�i�<�;��D��ݕ��Hp\��Y;��ʬ�탙i�Ͱ��M�O��*�x�v���)�.���ψ�!z��z��&�>�y�\�T� �T�ķI��45S<��S�;B����u�*xʮ?�L��S��EZsC��>,��/�\���/*�V��M�	�QǩϬ-�)&Cںn7������	�Wx鈫5�3���!���Gt��I�ʒ2G"U�P����M�iݗS�L&�����\����U���om�-����т�·V��
��v��r`\M�����vzoZ���g�#��qű��'B]�+uo�]4@럝h��{Z�-�LA��y��B��fQ���:<cZ��w�tȳ\�aUN����J�}F���=��FT��v7�Rʙe�(ht{_�t���Y~t�wҔ�<��T�O����;�/��|-��5+�ط���<�����H\j���9�g 6!���'a���l�;U�fEQ7E޶�wV9WIk����Uj}��yo�'«�J�{�����ؔ>��3��їC��Y�@�z\U�c���軈(E��8g%�5����g������z�b�Βc��CL�V�
�h5O� �:d��v�Efc}w͹�0�]�`�i��c�]�=�O���Y{h�\ԍ��_�J]�һ����
`5�n�32n�|M�_KR��*���$y�@���NK�q��A�F֋Wj0k>Bx�}��A��\�Ƣ\տ�#��h1Ԗ���ˉ
�ℭ�]`�g,]fS4�z}o>�O��#k��l�0hY�C�۰����|Ҵ1�������+�g�g�s���0kҼ1Wr�
<�hL��[�9:�Kf��W5~�l�}ǑѼ���8����|�J�u�.?g�w�Sӓ��)�ق�tCޚEY�m���-ӧ�2N�|��ġ]�x���=Sy�/s]�:���Dyep3rۘ��T�\@B���:��C�;}fM�[k���,�5�U�sI���]�+����x�6�WO��T��%Q����H��e��]1½�Qֻ����(���QQ=��mv̿uu����O�lV#"l��WdD��}:瑿�y|:�U�`_t�c9���	�Θ3n��xuب����~$p�,����:{�=�Of���*1C3f0h�k�{lKU����x����ea[�WL�8)՗g�=�^R�j鷞�f�V�	�V6�)����I\�ٕk�u�H^d�c�0&� �tl洴�TZ|n�! �j>�s��YZ��9��n��wn;�*&�;���c}�f�7hLV�m�ͅ�o�v���]�R�^�G'3g��:�Qʦ�*�Α����kl�JbĄ��+ Rn�e�*�;[ׇ�cc�n���\XX�j8�ΰ�� s��� ��l��Q6f}��t\	f����)�Q-t5S��=�*�+5�	��V7׬UW��xV@k�o����\7{r!��l,.�&q��+5��]bI�`�V�b��N�z}AVE�Q��Ȩ�Z�&�e�N��`g�+�4�sA���b�=W��jo��(H�3F�a0���Ŭ�����mˁ��c��Y��Ľ�t�wi�g,hl���$��ۜ�Z�`3�p�xu�#GI_hՇ�W����UlƍZU��,��W��=W��v��ڨ�ʿx+w�(����{�M
z���}|��.�a�ީ6ov��rID�(���rBG���p(�)L��u6ۤ�>� �3��Jp��dH�[�<�}/�=�/٫l,{��CESq�Ѩm׮��>��R��j-U5��;����7ڟ���h�f�sz���\>S|�M�qX?������5��n��*�����Ζu����&���)Ԫ�'v�(h��Ma*��Z��_�,OPK6c�0��γX����L��B�^�������/i�Vb�� �tz�2�a�1S�ݼ�;��"�Ҏ]c�	�J�u�Q��V�cD��K�#)�b��xY�Q>�PS�-�x!Qf��n�AJR&\��Fv�������B��
��9�B�:��A_��fd�(l@��b�TZ�[٥���+��1�-�	d<�plt����#����s�#��w�gp����>��-�������>��7z�	�;=IJG����Nz�X�w��Ojt���0�$-fa�n��g�L����tg������:�T�)����O�-WI�v���[�=WUڧ����(��|�x�6*�3������Å��V;"��$�yf��[6qάћdo\nV�܅ZYSD������4��\-5x�`����E��W[��N-˚�Oq����Ռ�q\4<���s�^5C�TpBˌ�T@Zb�R������mU�����4���9F.u��ׂ�K�	����L�^�41�)Ws*��v�.���7٤Q���|oG�`�ҹ��d�S k�gF�OgKeyC��q�4�d�j�P���w�E���L�4�TU"���s�}s��w�r�U��Us
�k���#&��ǹ�_T����x��6�ZF�4��HO_g��cS5-@���et�T���i����w���;t�ZZ���b��2�,��.���G"���8+�R�[D+�o�d]d�qȁ��[�N�k3y1B����Q4�T��'J��|����a���aϞ)�%Z������q�҇l�U*v���m��=ʶ_I!c_ik��gQ�A�ք��i�xnuXQ�W&��
������"�<�-1a@���S���s��1��6"jrI�>��MSFB���1�W�ݍdM���m{ED.�mnZ=��#7.������x6�p)��8B��i3t%���%�O�����t�5�َ{������.+a�hrlO���&���Ђh,�,%�N����(G
Gh��S�Y�)��r�8](s��>Os�>�h�Q:�N{�������@�"LZ*��;(U�l��/���������}�6����7g,5��i�`8ΟtW��#�새�b���1��S;�<Ί(&���WFf�Ӯ�9F�
�����̡�E#u=^�v���0¨��u������j��r;��P��I>�%���u��Jw�L���
�k��`mdЌ����]�{f��s
�տ�-��^�껟h���'R-ħ�h���e@��J�~��"۳ٹ�X������bHb�99X�S��)�ӻݘfn��t0}�X׋K�&�]��yO-��xW �S���v`�#|�by,TI{�Ŋz÷3Wf�*�{���o'�ň������m��d؇p�q}.�V������� g�N+
�G�n+�H�� �U�1�nh^��o�>��e+���U	Y��z����Q'E쏼�ӝ�,}�n��N.jp^�b.va@�>�nF�ۃg���w4���*�,*� ��;�6?U�W��I��fp��',�,v���C��Le|��;*"k_Z//
�M�˯�p�s��q³�6���n���B�`�"�=�:�����o���׵b�wup~k+z�<4p"�'�r���zք:�����g���{'S�K���ƴ��*��]^�A痁�+�`���Z���p�#R�p�����ڰ�wC�:�FJ�A~|�{!�4���2�C��O�g���:n9*#��.@d^����K K���*$�J�nc�OP�*ƺ�Na�A�J�W��C (c��
���&6�����K���;u����v�{�5)Ff�(c�:�h�Z��o����T�w�p��8_`S�+1��B��_N��Ɠx�	�٭��_x��U��h#-q��LT��Or)A�o�u|c�S����lb�GY$f�B�U��LUy���ɱb*}��
��w-��,0Ů��] �=]M��'h=��Ju��7�ҫs6��.��[h���M�uw�J�c�qz0�Vyo-��:���b�v����P Kr�po�������3G]E�BXnk,Yp@�M�V��ܦ:k�cB�u��ևD>Ȩxa!�r��l�0n4�~Ţ�wJ�1���^���f�}�:��ꍰc�����,MAL�Qr�,���Qe�*���$o9z��[��%q�'1��Q���]/H��f��߁��(4Bs^�gE��@4v�ӺQ�(d���u��ura�N�3{kX��R�k²YU�V�����ɍ���:�!�a�[v�wW�r!�J�f+��c�������Py}k�Pd�t�/���N��%.��$��mж��jn!�������1U�\�Ur��©�v!M�ƪ��͚�5͕��,�O���p}��ƃ���\�;Z�kF�E��+�N����=k��^_�}v���pv+��(Ivq<�v�؝��۶���NgZ�,+��6v.�K
z��ǖ�����:�`�HP�2��@9��R[�,��hI��ʤE�o\�}��s�^eowW2zu�M<�,'+Ox�K����tx�ǮC���X��`��p^�W�Ƿ���/�X2u����|%����ke&9>�	��5����#蛘p*=gw�!�Qƙb/��A%1wI�p�s�x�0,hV1��"��&���ӈ����1p��5�D���:z�����F٨m׮��P�cmʉ��t=ʅ��2j�v:�}���˭/����<-��Ξ�=+&��:B��+������ӓ��L�Ћ���M����ބ>��\#qJ�G�b�fذʉ��	�	Z���h��1��&�6'2i%������đ��#p��T��8TcB�v7X�c�(Ja���r�F. A���j��a�/[|o65-�b��m<�pv�R�b�$e�G����)`�&�N�l����>ְإ��ͳR��Q�M����BX��Ȋ���'�(���0YTB�.v�e�����s�sV�Q�a����n�uTuG��b3f9\�Rx�×���Pc�˥��3��S�h�^����9c���c������)��`��<w-���N�R��e�n�]���o9F�I�r���',�k3r�+�}�^�|B=�L���n!oH�mmD�S���g�.��v�L[�`͕<�=8tǛ^їS�uddQ�F�g`W�4�/������&�t�)3�U�ز&�c������Io��V��.�gc`�����o(��(�"�F��S{���hN����lc��)+�͌ ��o���V��*�#Y�ӹ\"jx�`�:��}g}�@�Xع�
���(GHݐ4F񰃂�K����bQ�=^5��p,B���vd\���)�����|k�}��acO�l89D��Q"�ꍒ��н.	���ꌸ��`�[��+�]���rʝ�Q�lо0��W��l
N�P'ye��P�V&�Ѱ>�	߁Zvtۏ�����z`�����A\�X�{�{�@�fa[�
�N�Lg��1#���R��b���>ú�O���pJV�eah����FCmKGpt�VZ1F'�R�4b1_�:�r�����UAR���Ѕ�Ϳ]���
/ӕ��a	�	�QGM=�d[�����-�	�+cxK]Q����:nϸ]Ho���G�B=�GO@� ����d}��;����+
��F�Shg���;"�Fj!Up!O�z*���)guEϹ�̱L:�It�\<�	��F㍳��/u�jV��֒ŃĢ8KN�g0�����I��=V�S�1�l��jUn�c�U��[.�;�E�	~f��u������+��7Z}��v�;�ӗKf�9�ET���B��g^�%��fE�Td<���.�R^�XS9���u!��Od����Xbwr�$��Ω&]�,|0�V�Hg�G�v���mLZ�Hhȣ���~AYu�����w''5�1���8�7�Q�^�>QL�3�ӈ��O�_���ƣ�c�;N�d���t8�FN�V���s�';�W�n1�R7=^�c9FX@���{z�ؓ�ذMlN��א�Y��T!l��b���
�p�V_��JEc�����.[���$"�oQ�o9$t "��~�+LX�	�Ph=�sL@�B�>jS����r���p��9���%
ߓ��#�\ڢĆ�dS����&%VE�4Uu�k��#Xu&��YI��j���{IO��	��ev�M��)�����>O�]B.c%�5�n�gG�Q�@PƸ�ݹ�LИ S��v��	�ڇ�z��<�cB��<���jc���8N�T��:T���~�$���+v�����w[�FJ��b�y:(.�8A9W���S%�v�C�ݬC�OPB�u��m�bd&����Îj��wc��%��R���m<O��Ǽm(��`���Q�;�:B����ٙL��g^W+��1l�݇lң[��=lu޶��H�(�OKo7���"sdǩ�.u��1i[g|�K�,Q�2.����-�IVC;���G|5՜=�{��Ҵ��\pf%�/nU�����>Y�g>�����$d�95)4�+�}m�q�ȡ��$u߃�X��>�LI�w���Y�H!C���mک ��0� �'*�Ψ���o�U�з��"L����yB5�������Bu\Y<�C��P^��� ���W:�gJB�;�y��baA�+2���3�|c�cSݢ!����4�nF;��6�"x�j�"�ږ8�*cy��6R �+-3��:-��4aQ�uY�4�!P�)�7��fg	Y�(���h=��U1-�v��I��>�6�o����e(����\�����M���a��J��M�|�u��r�l �NK�<&c��{`�1_-K��l]�#y!��V�_\�WN�(y���z�*{�: �����NS�jD79��:�N�2�P�q�ZL��5��ⱌ�[��L��gT:$fh �1!�0pj3�w��3}��R^���B�.\�h��7ƙ��N�������c�E*�1^-�F�Je�뀊<���Z����sE��xήꠉ!Y���s��Ȉ��j��پ�;Oj�8;��I��Z��ָ��IS$��Z��5Wz��d+`Ƕ�UC4����2;a��܁U���f��t��҆����؄��-�}r�k��-�q�W��q�v&�>x:�������NΥ�h��/��,)��՝�t@�����r-u�o�c��	�k�4�B��:ݭ�IP镥�&���8�w��7ʐ�X�l	l�K��4VTRmq}��Ub��ĩ�b�}�1<��@q:2��'��d���WtU���%����A����"����4��*NaݝWx�r>/��$a/�j3)f@̺32j�w�㢲�:%��4۱ۯ.�����O.63/69g�F{]4F�D��i{L�f��W9����z�DsM(V�G0\�'�Td\��W7yT�t�p�s���n)�9�lZ���D���I�,|�7,���<T����p>��{s�c�1�������P6��Vim���h\MA���昍��NN=Y-3][�F�"��{w.+��T��� ���Y� �r�р+`R40Ve�:ȫWZ~n��@>5'�d5)�5rD-���U�KQG�JL�����F꜎�E���j���gY��mZ7L��2�̙VE�������--eF�C�AAm� �0�K���
,Em�"9J��*�ʈ��bH��41ĕ��X�,TpcJF�V5��UVj9s�U,���ZZȫ*U��Z�-*��iH��D�DJ�U�Kj��r�!D�%[J�-QDQ\m���ֵ�����@Q�J5
���iiiT�iQE�����XZ��4�-�%ih�Ym�kej�˘b�̵����Q���eaU�
���lmj�F�+Q�4��*E)Z1�j�UQA��F�Em(�Z�#ҷ32�-��QV*���[P��
�r�	����'����4��juWU*EL�|�cŻ��p�_wj�̓1��j�9�ٞj�ulʃ�hVe
pȂ����D�N�w�3�]$䳔i�����*�c�����ީ���lvx��"T=kB@6ȷq?ov̺w�ޕ��l�+�<�Ǧ"�W��N�NeV���ڟ��W��^e��A]���F��W�P����j�T��LEq�y�U��a
�N�0���;�Q�%�����v�e=沄�������*O
Ԡl��7�Ra
ҥ��u�<'J��>>C���޹2��}�P����ʯ-����tk�HVx��EܷӍ�`2��HM�]T�۽0�����˛R��R��N��2�˯蠥Q,�����y����_H)���"���mS;N��U�r�pn:y�����l⩊f� �^���HZ��0� �v{���'��o��@j#gG����D+�z�7�{\�}7'#F�\�O3e�t���Ջ���f�:��)�ã��ŉ�)�)�V@X�p�X���j��ꖯ@����N��*�22pFT��߁���(�Ӛ�00C�	(n�ي��ܣG-XAY�B�#���ˤ�nr
�*�w@��p/i��1$���ҳ;��y�60{{m���8�
�B��15{+��`��K�B�pqqKEM���S�M�Ie뼆G��C:�UCp�-R��v��Ц�;���q(8��΅��+ԍg�:)X�m�c����!ՑxV�F�������ilwS23U��X��.6k�^L�T�pD�*��^%R8=�S5�na�� ��Z�]Z��"�����w5G�wuEk[t�i���VN�-h�V*�IWB�X���978t�KpM��t�v����N���A��{Z=p�Ԋ�̭�MM�=3ْ��WGs
DoK��F�����a�\^MD8Y�5���*����)��OE�<6\n���d�����Tv��Ò�H����蜘p*΄�$��{�2�\GF�Jb�i<������wf�e�4h��R�������U�^��-^9�E�(\		��m�mׯ3\�UW�˵�#՘�s;l�^������߷xa���
�<<<�N��i�h��L9�C����ӣ�5Q����F�8��#±c6ŋ�*+���EuFSF��8u�^�/9`�W��E�9\@�h!XX�8֛�nhЌp���PW��ᗄu�]��$�o���ؾt#RE�����ڣR��)�7G~|��V¦"��<�]q�W[�����W��t�����s�Q���)�r�l�Ó5�9��+���e��� ]klw[��y�և�QAE����Ok'r�6+��N��t�&��t��Pؾ�w���ӡ4����3ԃ=jl���H�{�P&r\k����r�8@ΝqSC��6�OO���I�â],WG<Y�0��� T�&uc���U�N�W��5�b+�cp�qPo
�l�u9�"l���l£«i<c��!��4�T�����qپ/P�՚�Ǝ�3pq��Z:=C{(�=j���c��w^�@П��_��e��Ջ6���e�����U$k1&r�&�}1Zʑ�A)v_=�U�̷�9#W�O��E7@1��b�]]�x�<��]>2���F }1\��6�7騮��;�����j�l8��\�$SsK���L�Gk#�7il �vtR�|&^�5�z�h�D�8X�.-��b��������_�P�i�s���TZY�"ys}(�C_��G	�lo�mXc X�1fck%�+��U���N�Lo'WMn��A��.��5זbC�TD��[7��ãge�4�ܝTa�0m=���S6���������5(���Z��f��>�:1D�[��Ԭ��d��L6ͩ~L�O�p���>r�q��޾Zm[UC�Ԕ���Kj�2���3E���(���K�A�H���Î�W�4�bV𓁌�.����1��2�jG2�;Ѡ���b�k�}��H�q��$��I�q�Z=\�t� �#Z�s�~���x�Q�9Z�f��^�;v+����\V��Q�S��W����Z��u���3aϸUB=�Бp2O��;ԗ]ks;��1��[T��+�r�
��y�V�u7t�o�j9P���Ù��@�u�L�1s��65^�;��7uLJ/�LZ�G�3q]\xs�W��\V��L%.�m����}Q�B���$�^+�>J��>���V{p���XS8ܡ��Bު�>��7u%v���^߽i�Q�X��<a��L��8�W-���-T���~}��)�ѥ�����:~��6ô5ܘj|����0l�8���
�C��Bx(�����7��Y�gx�Ov��q�,)S6���1֘*��7]>�[2�[���]��uF'�jv�;�L)�?G` �R�C�T����B�n��X!uws[x 	���^�9�l�έJ�a�\"],�ͳ ��oD�i�b��@S�Ɯ����$|�.�����{;ZU
�m��;�G�Sz��to���1��d��TTl�a������z.h��%+F��Gp��x-��~K���/��	�#��Go>;A�M��!��6�i��ZAgzn���xd1�t�:ߘ[��Q�#�u��0ѯ\{��*��o�Ly�z������y��0`S��}�Ĭ��h��ڜgk���f��E�o3-�K�zt���>��?�7]���\x��,��b��������f�e�*��_A�!�V:��5���##����As��;~� �Y���4���,dk�!<�)���{U����5	��E��ݑ���E�5�zᚍP�ã~ǜ����4�پ
�-��l�;�7���{Ӣ6�:|��95\\�Կrś��W��o��x���H��:^$�v�Ǉ���8'Jވuc��I_�s�syR%_�M!<kp��5�����=��rkupH��&b�D�����{1�2�#�M�q:!n_��nKx���u�qu�:�	跐�{�T����3��T��w2�&�7�j�E��ZU�uk �o�}��M����ޘ��#@N�ҟ>���tk�_O>Q����"��(�ը�mc�N[x/���888�8Tj�o�!�>�.HqЌ�O�lV#�kYub& �GҔݺ��2�S�M�,S+����P1�n�:ҧ��Sχ�i:����
�L�Vb�� �t�et���Y�^��eQܙ��b&�=�h�Ӆ�� ���gg�mi^kM��7�;��sKp��ê�b�މ���M��v��JB�<���������SEJk5.S�qZ��44�u�6���>�[P`O���q����8#A���WbG���ݚ.��`��/q�k_*�ĺ�С>��l���Z2���N2��R����D�������v��F�V�S����Xxz�PS,W��d��	��P<�=b�M^�{Ț��.����(t�N580l�W��϶Nv������yL��&�a�rS�p�Q���'Ŋ�s�2�	��V;���5R�w����ub��&��t7�I�3�s�ݘ�3��\�Ml��J�F�BI�~b�٨c�1ad�Xa����ܼ�6C-��ݜ�#�|��0o�zv���tkw[57��	�`��4�H���f``ael��e�U����P�j�r���Ճh���A��npz�W=������j�^KF�E���WiW��~�2�lY�����z��#���s�Z1�p���6��k�Pu甬`�x/%�W[B���/@�����D`���l������x�51[)�h؄��5`�����	Wل@MI����jņp����O}�r��e�Ej��5����0i��rD*{�1��N�ų�r�-����(	�9��!Wյ���:n.u��4�}�dBH��.[.0�4��U��#XQ���J�R��Zd�r+z=PR�w�5�>��0X<X�Z��Z(\		��q�n7_I���ccy�e�K�nB����܁rW���*a�t����]h����K�c�(ei}ڕ�����hoϝ�鉶e�yVq����Έ�[O�K��1��c�Tf�	5�C��#��?3�q�5G*A
E����n��p�zel�V���M�2et�!+�7N�k�/��"鴮3!�!1F�v����g�6z��!D6舋��덶\��v��y#�X,�9ꦘ�g���p�������
Xn!\�5�md=�{�:��.is|j�I�����v寈J���K{T��G����Zs>*� URƽ:P�S�"�U�������X�y�5�v�G������ٛ��VU���k���\J�P��E[7��
��5rѤ�!_vXƯy+����j�$����!յ�'�t'0��p�p��fz�γ^2��3������N���ڸ(V���n��XҦ�.ͥ�� �W.�i��}R�M��������
A�p�|D,g}�)���;����3T<�oiL�3�96�:�ۼ�r��.�����cQ��3��z������+y�3q�����{����w�^����ą���ic8���Z�;)���zYᙑɓ5�G��ZgSt��E�s^�����=��)��ö�Wz�aW���k�j�M�	d�~8���o*�����;�G�w!>�PZ�C~G)�t��V_���Ъ`�N����Y�nF�0��x�`�Jkt���\ឝ�6z�mEW2�qRct�:��X�k�v)��{����d�O�"���y�j�w�
_��ǲ�/.f�a��KK��'j1�w{�ȜHEo'Vҥ]ʶ!K��xu���W��j7B����ӝ��;-�q����r�
^y����nC�Ƽ��[=U�<T���*��]	sz��G"ߎ\uD�>��o����j�j��i��d:�vw`��o2�7���Ժ�x[�z1_��J�S5]�WM;�i;�kC�g,Qbu�����㉥lה�LTr6���fڿUp�:���3;��m��͸�%X��vQ�t�3� ɫ��S���];e�i<Χ�>�r[F�/L�Z����"�
�ʿ��eI$f�!��o=�W�RM���5ҡ���x�Wv�{6�Sb�.����	Χ�}p��T"ZJ+��w�oeCհ3d�F�쉕�r�+6�w9��p�n��TסS��a�=�"�t���=�bqUM�����VU�=xЄ�,��nwQ	u��n�Tb��*�©:)���$�OTW���Xcs:�D�E�(��*C�'�����󽰺)�r�.8��S<���|��Fq"��w"����eF�.F�iv@�gF�ev�s}U�8�Z�g�Ǘw��i'|���Sޠ��{����z����ѧ�`mJP�rj5���k�q��f�Мk2���L�{��j�Ɯ7X�}��ؙ~��|�.y�j̵�L��d\Z�R�u��Ģz���nZ�|��4nc����wT�\������^f�Sʛ��؍YJ������jߦ\Q����]m���AOws�w�*
&Y�{��d��?l�t���ku�:�]��]ѫCPR���o�R�5�e	B��^���Ӥh�6��1Y�b�x#�V>�mj�o�]U7Q��E�ڑ�,���O�PY-�Ԭfќ�~]��pg���Ș{n��mNFҊS�Y�d��T���H��wNA<�����}j)����5p:|ٯ5�
WDR�P�
j�{��3F[�q�g��U=.�������c`��J��@�4��Ka+kw��N\tg\2���%�=6�U�+�!�#^�&$M_tYn��v�G�C��
aD�i�kc�͵~�Y���.;�AofK�kat��Wgrs����B�w�ن�q�Ǣb�_,<��螕���+}����?����j��y��{���q�h���^k������J���{M���>���WZ��Ie^{�^�(�z��`2Pl�حyj����q�E�<��,JmK���9F�+s))�����x)P�Y�;͕s�'=�����c��oF�4���Y�3˻����cV��f�߂������a��<��VO-("�ɗ�Y�S�0WzL�%��;�-�Ys���[_Fy>z�[V�ex��ݘkuj��Y�q��)���|�Dy+3�4�ނ�����z���f��l�|*+x���r9�J��7�����f�c(V�>�Cf���q���F3{)p���+'d��mf)���&�������E�^Փ�$�����(�ٌ��[�A�S�v;sliս0�=m2 lܨE��bۜXS�ev��f�3�����ob������}M`ќ�S{X�������12�F����3���̸���M:}�1Q�{�ջJ)̷}2�o(�
��ê��&�e�;n�nrf[L���*�ʳ%�7�ň�9Y|����v����4[���N������׳pa��c�u� �J=��4E������[�!�4���h$�hv�:�v>�X�uY�Ê_�\��]�0��*%s_Smҧ{���K�Е�� �G`˴�;��w
}���╢M"��kKK��5B������}|��P���9+$F�kh�]W��P���^��Oz�i[��]���{�&��Z�����s����l=:MlY勀f�3+K��mm�B��o7ʝt	�D��%%HZ��V��]}%���v���GH��q��/�5��tTu��\���)��|����{�,1�	�=�Q�^���v#Li&^�.�[W��34Ɗ_h�m0�K,=�vٕG�#B�W�_/���Xd�^�b�������+�e-Ք0v�͋���*�[���|�۳Bq��`�����,�eL);�:ZX}Ia�u��=|��5��{P��k�%���K
���8�s�K/��h�P�*���D���.��1Ջs��P���y.,sST��rʶt�[�\ �WC|zv��H�d�\�;�1h왧R�W2wh��oQ/W��K.n/�1��<D�T6��1����[���h��;��Ą��aX)���_r�b�������c��ba�x+d�Pf]:]x�Jon�������7R�ꩽ����)$®qE�si�5Kh*�k��c��އdZqvˤ���m5t��J�;�k��Z
�c��[1T�4:�p9�-�{�Y΢�H����骺�s�¶J�o���eQ���/�Xn�zA6	O�Q�Q�3��Yj)����b[x�f�b�����]ͺQ�VP��t(2��!FC�V��E�y8�b���q�S�a���켆�f�N���WR���'�8����׺�qT@�+YZ`�j\�Jĥ7��|��#x�n���I��:�	6���nh�ĵ�Yw�6Şt�5�M�E�s�gH��B�|ja[�M����k���Fu���r�g��.a�ۣ�+�L��G��R��/�Oo�༭PS�*��X�X�V�G�0Pd�9��ޒ�,wt�[�Um+T�{��^��Kෘ}����H��6H��Նh��ף��R�8��-��<�P�����q�%��Z��=�`��/�B� ��"�{%[���F�fL��x�J(H)%��m�*�m[h�*1�ڲ���%hQ-*J�"����D�Q�+*��5AciQr�YT[j�s+j֤R-ecQ(�5[Z*-j��Tmib4jԣP����Ke�m�Q��kklm-�+PZ�b�++(R���F�̨�.aV�2Ѣ��ض�%��T�ڭ��Z�
ֵ���X��YPH,��a���х�R*�KKR�Z�Em��`�Eb!QJ��fF���T��5r��XZXڪ�J�ZD�L��--aiF�J�V�E��e`�iB�ciJR���*��Zѕ�e���V5QTF�Z���1%�TU���T���Ymֶ��-��Ueb���*	$�O�'ȎźvLR�R���%U�ܾ�����0�$`�鏇m�Ma/�ȱ�|e.0��w���}��
�<;=yx3پ�˓sn>���dU}���\�q��MP�`�x��@"����ף�w�F���mS�C>|>���|�k�O4�{S��
���|#�=�%_'2��ƥ���;*[��ɟ��&��xVߊbej�Rӣ��N*�Q�aQ��j��^F�LW5g�\F&���Q��i]ʔ�����Z�f�y����Ô�������=�Ͱt�{n�;3�� �9N��{�1�Q���^��a��������8+��s���ao8��J�}_S�����5�|8K=�9���"�єo�l�����G'�}{ϥꅻ��&�gw��o�������v�1Z��ֲ̮�E�):�/�c�1V�B]���P���+�56(+ܻx̭�#�N���i��V�{���C�dTh0|=՝��]f9��]�t�4��u%����}�=���R�$L�dc���e�f��Cz�;cRyd*"[��|���`����쒻P�t��)�ҷq���:���{�.顽kV�pow���tk�m�xH�RЍ��]�K��l�{ܷf#了Ϫ�Lsgq\L^*�S������i�`Y�YxV�+����L%�	�)j�����UK���;�uh���{$�2����������ꃐ�Q5ʩ:�9H�w:+3�|oV��\7��|�w#1�f�Fu���')�se�R9��c:,�T�dq�5�u��iX�\�>W��+}���f��5�����v|��w��=��:�0������������c�e.�����=Mxh�۷��d��i�ꢍ�j�{��ÿ�w�Z�ד�qlX�:�����m;%�OUt7�͙
ʮzɟx!m��[�`VFɪ/Nnbf�ޅ*���r}�\����"u˗��(�[�c���M K�47�6�c�Y��[p�RJ��ˎY���ˆz���%�T��cIEM���z�����BF�>csh�ݫ>�$D��7�P��k���X��M��ԉ]dd�| �׼�7,��3`���>�$=�3��+d@t�w]�X�� ��o\�ΩY�"{y���K.V좬��vt)Aܔ���/j��=�|�U�B����o�<�q�B�Ň/(!�|�n;�V�5�+�t!��$���1|�u>W�ˍF��mjV�_g]jd�(<-^���ˌ�\R�3ш�K}U]Pɞި�����U3��ȇ�yd�[G���ه:㝅^e2c�E��s6��a�U�}t6:�\�X9\�{ݲ�5�㭩��QۻjDcIEC3פ5�
�8�������v��K=�u)��3��7��Wo�y���EL�u׾k�,b���_]n�����u^K��n�c삙��XQ���Vc��_as�r�_�2�Q��H�+�,ܦ�K��י�܍i9uV�t;=��#0\�:�س<�.��3��{eD��#Ω3{Gb3�c �݁��^���;9*�`aj�d+=�9�yN�_=��EյƳ}�i�+	����e���{�%\0����<��ѱj�P���z��Y%2^9���ˡo{7��v><4���{������>4��
���;+�{��/�ɠ�eq�B�&�7z':�ݦ�T���A�u&rT.�OR�[C1�1�ֹ�6�^Վ�^��2>滹�c��:Қ�ΰ�CV3����PW�0K�.���8Ԫ�[���_vGMGK��
\��ՙj��y:\fU/�I�Q�Z=�����:u=�=�^�Sɛ4��<���v&�]Z����k�Z���^5Ϻ��yVs2�6� nϣe��h�J짻�w5q�WfݐGl2�3�6����QQ�����w��M�Z��nV�}f�V����=�^�5�N�h�M��3]��=�{������0���·2V��ռ+��b�m�f���ќ6�G�5K&�Zӷ�9�������v�1ϩ���݃^R�}����D�W��S�8e��:r���MvR�}��O+�|��-gym�m�ǣ.V��	yU(c����Oa4��C�j;�׷ue��5��=�x�BAx5o{F�����p�=S��ew&+s�)%+���Z,U��$�T) �ì�Krǳ��{�?M����qf����H�`�����@��_���$�D�����/��蒿�8��xq�Av��榕��*�T�Ϻ��XN�x/���7tj�_'�o�*��~�LN�1W�t�{���I+���f�1�`�tNݍtѽج���'8�:�F+r��W3N��)�1�/y����0b>��Zns�'��cچ����6�]D�"2�zrӸ��`��ѓ^�p���ӎR�)Bu�N���aH�`�S:�חV�凱���N�z��]��<�w��#1��� %sɨ��CT5�3���Q�%�����j���C�gi��~{�1���s��[��㎀�uC���8��҉Z��jj�[�5K;���������i��k�'Vr�,OWاB��|�X����'��Yԗ�(�ϩDĞtV��"��T�.�ڭ�����c5��[xjf�a��G��>�a�Wa�G�e����t,�휘{��ks�v��ⲡ��G޸3q>:��O�V7
��|V�)Y9ܮ\�ڷla�"�K���٤�%)c�ƌ�Z��A�V��ҙi�.e����ܢb}�|b�9���!)Ŋ�=ĩ��H_@�t����Q}u����VbRK�q��͘�C:G]!6�gqM����y���d�B���2��4�x�5�`�K;1�7����bLϻ��bM.0t���]wx� ��;C�-�T��}_Wں�v�C�E���[�A�#��㥄�����M�k��=W໔s�|�;{�x("��Y�F�B�]��}ؤ�vTeA4��vҜ��U����l�z�{�x�Wr�를�z/��b��y�͑��m��o���W��S/���+Y͋�%h}L�����q��U�Xb��g��E��5YEM�o��T���,fwd��<:W��ץ)O.�~S��TIΧ;���^+�;k�=�L:IΌګI>�R����a.�~�.�����s��؝uFr�XG;#��0o$��_N�j���b��on{�b�#�G��^��9��Y|���ȷݣp�B��������*S����ڪm*e1�~R�>����W'U�{���(��)-�=짝C>]A8n��4MG�i����C��)��Mb1���7�t��'�l�F3��)����]��*�Xw�E�'p��i��r��Dk��g��N��1Y��Ɩ0���WU�����la6G,�g�91��,��/���Etg��Wk��u�4���Ŗ��sJ��݂��n�>�3^y���S#7HU���+c�wW_Ft��;[��q���^�����[5y[�}��Y���xf�1�4�|�.�M&����>������W~R�/ܰmD7�nឬ�í ;�����#=a�n*;A�i��(R�6����^�k�V�{����jDT�tL���p�BP�K���1|�GS�p9q׬�"�U���8�uejS]��:�iO^�׎��JwJkUT^{����$��Vl���˾}�t�S> ��ϓ������:�\���i?t��G5�v8��鵰!����'u$��\�i��ͫR"|�QQ�w��.�辇-ڴ+�5�Y���9*�ݺ���5)�B{���Uf:a�@�E���.&�+��3>B�ѷ���C]���D����P����mp��r���N����X*���<ăAv������*�MHN�5ܖsk93��Ԣ�tXʍڀ��W�I[��v3;n��qrz�.�us�S*�&՜-���(���v���RF㉶�0��ځ���7t�]x��\�q\��x#�=S]�c���6Ⱦ�|�r�yRTOe/{Y��MAz�����a��+F]ks�i���9��I�j��5ΞŬ3M�F���(E��{�`�]%v�+��;�S�'W��J�sW��'�V{%'#�ŦPʗP���ܪ��Ev�`���أa<3֙���k�r|�ڨ6��㞡/�2�r�Ѽk��s9O��g�~vc���F˘���7�j��5`�5�o�-`^?O7\+:'\K�[�Lt�@�/E��el�O����V�;}ݚ��a��|�a��3�5��Y���K�33N6Grږ��$��S-�QGK��C�M������٬4(?u�[��<��T�Vp�nP�!����wp\G�61�2~�'o����Q����^c�x.�Z��-�:�'��E+2���|�[]5��.�[&;�f�j�s4��ٽ:Q9��4x\��]�{ @6����~��`�7)�E�<z��z��Ԕ���"��)ҢJX!�`|��Δ�o2�c�����V��C7�R��OkTj���m���ʖ6ٴ����P0k�hW�ڎ�S�9T���|w�~U�M����t�)@D�5�h�-������xg�Z�Hm-�v�V�U{��;i_�)x�u���3��_1�;2o�{��	��<��n�ݢi��}��[��W9�'<�J�n�;�CҗRY��f�?�	r���3o ��\�)�@�z�o�.��f�9�"��{2�N^SP�
�D���r���CT�����y�s���m�-.։�{��9Kb`�#j\���<j���Rຕ@@c���a/�5� �glН'8�M��|��u�:�1��n��K��%@�p��ӛL�q��	��&��a��k�g�h��:�v��}��t���WBW]���z���q���b�p�H��b��6Kc%o�FU�=��Cz�T���;���%�eZu�X�p����]�S��eh�ƪ���v�׎98�p��V14Ar+q	�ih���䗃C�xQ�I ;��`��vjY7rQ*���tLC���͛Q�`��N��!�*܉���gr��e���h/�V�Ҫ�(Z��Yn��o[��;gkr�v�4�2�Uus���5����b�c���h�5|������J��V��މ�̗۝.F'�+�+u�ð�A��Z����tSTs�S�%��{ݩ.�l�T��:(�-TC�+R7p���S�k�Ԏ�=ߪ�kP�tsۯ`�k�˜�-8V��M\J�C����uCo���
��ٞ�]BzŁjQ���Z��Y"-����.�ȋ�U��X]��s��˹W��_���{q��eI��d�C�n����=D�u���UV�Tvjw��3��+V؍��t��d�W\q?%by�⣏!Xw���Ϊ���uU̷zU?V������z���7�]�Xb��g���(��}�����	i`=��KzzN�Umn��v�U�N��~SXꓝNw"��2���}�
{Mw�����<�$����L�\7��t�C4�K��R_"�'<|:���f������s6�<���K���wb���}�,t�Y��|���x�Q�@��� )���ٛ�8�Qr�w��M\���F�k�=I��'gXղn�����:��v��[� &�h�\�[� ���v(K�"�T�8�bm��ZF�������V�,�����yT���spKH��bK�s��f�:�d��M��r�;�.S�a����(��Z�Q�oa�eE'g�Z
��*3�д>�Ϙ��ǝp�I	L��D��J��0Icv� Am�շoy�Y����YҘ������+�b��)F�u�����y�ɽ����t��g�m�9��ܶ71s���e,C	!�*�7m����ۙDST[VpI�pf����t� �D�� �s�[�)�,fp�l�Ʒ�d犃Eή=!�;�&k����D�B㾼�e�ݬs���.�VÏ2�NL�Mw\����\D+ܮ�%[�+�r�ؠ�5ޝL��|;D�4����B�޾�2�a��Oe�.����:�4��rw;��BG�>�s��,�-��Qj�V�&�(��U�7�C�D�n��ޒ��5��smS�r�q�L�+�37k����ɕ�VE9��ۺ�s��M�b���!'�q;u�-�j��La@�0��4L/�M�����4ʳ�"(CQFp��Κ\��꫒fd�,q�I[�a׭Y/#;�����r��B)����6S�uҚgevX��<�%�&k8K�[�i�2���.۸gf�-�	B8Z�]ٳk��{P�L����W��k�ν�rR�;V�vWC73�U4�fJ, �4{i_Xg�7�u7��3�X�!GmŒ؏H�JS�QvQ<�R���7y�I�5{�\��* �*df-�r�C�[������w��њ)��P�4��ed1,����a�A��Q��N^�ѶȬ-*Ҿ���q�a�tV����L8���59sRߋ�613�yu9�Z�w�Q2Ƌ�1��r�w)��o��+|C�#�[�ݮV��Ɠ�I�.i��q�	/1F���Y1ۥ��f}e�&�	 ݨa�X9�7[�sJ`P�e]`J��v=�]����o�%N���Om�,�j�
�v���n��i�l�Ӣ��a�jN/�'g[��L<fn�6�؉N!Hi��։a^�B�v�+���Q�m`�1"�	���1��Sm^�t/�0y�@|��;4�!mj�;�4ƛ�9Vӈҕ�Ӯ��pLPWW5ݾ&h�ё�A|1��6��%�gZ)\ ��Qϡ�7)_
HT�R<�ۂ��Z7�T� ��zr|�U��R�î�U���+cT��
I.�w,Ы����PY��3�r�U�b�ۣ���R7�"�U��z�F�m=w#	H��P> �T�Z�Z��UZZ�m�B�m�W��0`���X(���hV�`�+E�Z�����mh��0�E�X��Z5�)l��!r�qJ�B�����J�ڥ(�R*�+ն�ұj,*��Am��S-\fe�+F�-T��m��PFT�+m���
5�-��TX6��YP�--�U+Z*�iE,���iQ��*ł�-�m���̡QF#Q)(���h�F
(����(�
(�L�V*U��DEj�XT(�Ԫ�`���DE�T�����(���$UEƦ6�DQ�E��\�U�R�J5(��b �[Y�PkE2؋2�(ֵZ5��-B���J����UK+b�kVЭ�����R����Z�
5EJ���U����[iR+*y�{�����vNz���W�X�;%�W,;�lp2��gwZn�2*�ЬՆ�3�d���us���4F�K�ځ��u;{{D{���+��j�p��MO���i�5��/C�^jGW�K�u�v5���14 ���<�6��0�-���w�\�z��X��Wnff6�L5�s5��	O�Pq�5�|�𣧲��Sެ�(T|s��>��[:��AtN7r���4�6��z��y�ھ̩���(3�^��'�iVU�ulqj	ݝ���͎�{S���\;C�n�2�a����}Kݳ���1��'Y�x�8ڮ�lסC6�����7�����S�hALT�<f���/rNܭ���T�yw��[�͗��g�bbs^��u���3׻7��t1u9އ���<���T��-��{�rfE��ݗ�me�o��ܰ�4o8��:���m�l�+����E�z��� U�]��K�"��=���]l¸��V��M��\j�Ļ�F��,r�9 �L̎z����񤭺X�9�1�kU�{�� �5�`�S!b!5�Ϋ�]���-X�`���G{��0N��[$jH�.Ńٚp�������}� w�u��E+J8!#����S��-y�;FXT�,"&��8up����ѹa�r�iIu�jq�]�:aס�)�z1_�m+���j�(��ʹ��tA��Ҩ���ws�s���5�,8����)����\-W;��m.�<�ɭml.��z�[^w�4�*�����ۊ��X�S�|D�\�G�H��U����[�fZ��[��v�\�^�B{����B�((�����"֎�z�o%h���޿��s���1^�j�뚔��s����]��1=Mc���o��
�v�F�Y��ۍ4�������Qr��o2[�-%w�����my�]q'Qed⟽�+t��{�w|8S��4g�5٥$Cn2}�漕aQ�j�\�^~[���~�<�^].���E���w�T���2)<3���V5��k��и�T����ݛ�{���8�ʟ]���^��I��f���>6���>�|f75��c1f�q�ݓS��c�v

�Lݸ�,�f	{6�A���I;��ރ��#B��|�)�����L|�
Aj�y�i�ɹ��;�7/8�FE#N���ݽEN�y)d�R���%\_u9C�u�%$4>	%̭��l8���&et��/;�8^{�㘵�7��+��ɳ��w�������3�+����o0�c;ӎ���Qy�{�e-eJ]]0:{x\Yԁ�ί���]Ƣ�7P��#y����j&"����܁����w:g�^R\���|�ڔ�sʖ��Y�l�TB7���#�� ��SAV%h��q^��aol�s���WLBo^�F������uו I;1������%��y��\�ԜoL��Qt�_��W�T=Gz�ރ�;���:�+9JA܈uI�Jr��7��-��N��;E�z�z�ف�Eͷt����j��E���⹛~;�(��i���K��g���>k���]���f�oi��9N=�b��=f��FV��[��j���^�'�3�{O�f>,F��	�¦��j�y�g�=pZ�{Z�YE�Ҥ(���m��^Ԝ�+1i��~r�P�K�(�)�5��]p��R���J��y�Vk�� +:��w,7�ؖ�+��k�u�&x�/U`/�J%�ͫqo�pu�ǦNI$^�!�X���u�	O�i4�L�b��(�x,���0�ke�WFo�c��+q�7�2�l�Z�� ���*�,(.`�5�D	5��
��!ßt�{C�=QL�b�ia�P�X>u��^t��C��9u�j�#q�:��5(Z��������\W8�ԧ��G��.'���f�3E���p'��gE�0�U�`˳��SJqc����1��i9��q^��\��7X]�C_ZL�^��q��6�'�/u��.Jji�2��]@�O2.M7ղ�Ψ1��Gj���)N�F�� �����B�ձ|o�V�����E�O:S鴀R���'���O��3�ͧ��9;}�߮ӵ핋z���`N�Qsh��vt$�o<�вS����|���7y�p���:����K���(W#��ڝ�҅h�ýY�����^�OzV�$��e9�Y�ތ��g����v���4�|��<����]xͥOtO��j�W*W����-����<1o�q��ם��e
�T:������HO�oTu>W໕�}QV�F�'31���T����)q�T���7�Rs��6�jF�!Gf0mʵV��0�>7u�Z�I���M�)F\�Ѱ_�܎��i��oa���3;��/�X4>���ܷM��ӹ:���Ο[u^�ʻ/S�4�9b�N�L��q�QmM]��ӝx�*�,8�<�FΟ%=Ѻ�Y�=���n�9��4��J����m�'ʡ��x�F֤b�11gm_�/FSyQ��k(8Цڌ�^��n��V�Q|��7�ʃ���+��'BJhɸj$��8Fwn��I>�b�3Q������Ĺp����tDYaL��=�t;��O�r}���^�l�da��}�f�	N��S��N��X�T���\��s���9k���-�1���Ż���c)9��Q;Ш[���t�J)������ٗ{Xv¡���c]�V:��[�Ve�ǽA�M[��⏟�����ݠ��d�C޽��:�w�wXB�lN7���I��dMA�����÷�q?-q���]���0���}xe��~�M�3o`΋�
ɲx�F�����f:�~v��P�ך*h��3�@m[��v��z��Tˆښ����VN�YIޜ�G�)�7�(W�̛�o�p���7��M�s�.�ЕKgWX2_E���#�7)��D�m�%6M����d˕ˬ�NrSy*�����헼��~����?-�t������>�:���,[���cD���F/9�����V��D�O'?b�V�m<���P�AT�M�e�f2�����z���3q>;�M!�ڟt�V:�m�UO����r5�_w_]ku[��V�rCq��l$v�W���Cb�uԹ8Z]P����U{��`J������ǯ�k���F+��J�zm���]V�CO�G.�\�-��X��������n�E��M���m��9bUeW5�Ѹ
�[��r����UB�u����MC|�!�4����{ՐOZ��ޓ��x��"�'��L�wT��VƧ��ܷ"��Kޯ'���D �`Jc6[fMwb*��.�U43pq�q٘�G0��኶������^�t�m>��D��}��*��N��[��-�Dda��A��	�S~�8#r�[W�`���ޖ��ru�_�Fbf���|�F�Ý���<�x�ֹ��)��Jf��Cϝ�F
��y�I�0��=&�Q�Y��Ţ��b��B��6w-�V*�GpX&��ۄ����R�=�ЌAD��wm�֐���{��4�i�܎����JӔ|�j��粩���ҩ9ޔ�����X�����eVs=��#|��K�|�JSet�����<��XZ�Fz�A�gY��.��?Z�����ϱ8�@d-�no&������06���[ʳ5�3kUv��;��8�^d�]��½�r��P�콫3�X;��8��8p(c����=Ӵ_?|��ڥ��������z�e�O��)v넺��[���dӍZU#�P��ٗ�%E_P���Ko�S�N=�k���i������p�{��ڍ�ߌ߆��S]���	2đ�R"�{:f�.�G�gZ~u��wnR�Sxv�N�>��k����S�ħQ@�i#;s�=b�(�oiR���j�m�܇X�B���T�Bu{P\k�A�M欝����9VWVC�R�o�w+����n٥<l�h�ش����p�����3�%�Ʃ�����{�m�(s��KҺ�J�з���ͺ.��|�ֽx����3��Qˍl�n�I��:�U{�/d5iī�G�]�$����̚�]�ooДwp�����ߍЩg,bR,����ՙ6�u��ɮ��_-�_�7�����t�v�o�}}�����!g@��rҘf���V�����b��&���V�w��V�;@j]&�p/������Ӫ���*�(*g����bܧ%��Ve'�f����g��>ԍM[W�%'��;���r�|5�z_�_JU3�]ZhT�L��򍛻uw�.�T�έ�5�t���0y�t��"�TI�j�gk2Ӥm���1S�J���]�;�����3����ާ8��͗qu��yqL�W�U�2�wz;��P��斑�K�e=�f��S�����uŬ�L.�R|��a�8Z�^ߊ��Gr�Ne�������t��Ê��g�ҽ�oR��e:΃=>��mz���qo������F�iV՟�0%]��wsJ?ov
��K7^M<�z���23h뺉�QxЏC���&�Gk})�[4j�!�go���$�圓�����:)
�����2񥮬�K�鬫k��^�'}��?lmu�py�
o��`s��Mj�!{u��D����cԋk��h�"qo%ԛ�Ժ�>�H��^��53���#��#/*���B�g;*:\�7h��n�f��7P��2��[я/Z�7��\ݠRi(�P�h���GJ{~�U�9�<�w��ވ}�v�S��md ��Tb}��$gm���8�b���MoRU�W��%p[���# 1��~�rz��t�cJ?6ҹ�y7j��U후�1I[���X]��s�('����ܛD�f�Z�R�����}t��j��s��Tw�Sz�'�z��3[e�Kp��5�G{��^rÇU�x:���)�֪�XlL�0��x��{���c�-՗�z��*���w�D��Q^�z�^�D�bp�D�Ic��Me�s�O�'=�ݵQ�#�ߞ��ל�:��S>ꑽ�S]<���.K��}�tnz�wJ��W���q��r���C�*�Y����z�km� hc�����6�FF�Fq��)�E:Nq����f]�5|�S	� �u��379�4r�w�F2�/E��N��Z5�ݳ2Z�j�&�|����2�x�>��h�ςU�l�z�S�\�-�+h�<y.���]�������-hˉ� /��93 ��i�3>;"�w�����)waQ���b�zzr)�^���~�x����k4�*�!���ͧ�X�'ӶbѸvG��l�R��}��9�'�uL���7��~t1q_��Xw}��:�uI�T���Hr��t�Wk�[6e��\f(dvU��o3y2)���ö�)8��f��S��N�<�ǵfzX<��3jvm@%�>��,k�o���n����w�촮:T�yw�O��^l�7,W<��&��d�#'9Ӵ!�ԏ;Md�V��D��s>����	�6���e]��]w5ꛦw�(z��h�v�f��L���Wr���kN�C]�˦EE��V����*ѵ��:u�څ���i�l_c���X���T5��TM�?�WWjnu/=yQ
x-��U^g��fҺ��<�g{w5:t�Nk|�;�f���4�v�gz�eo�����Ǥ��f��|F�:�]["�ǲ��a�,�fI���v�إnc\�X��1�;��㯱�A�ؙ-ՂJ`��#7���H]nѷ��z�rP��F��6j틃�B�;�xdW�˂�94V�����
�6����`MFϋ�;ю�n�[S �F�<� {q�˩P�y�	U����W}��;�Q�Ƌ�꬐u�3(����{�b�M�i�;��V��
b��V�E%�T�m]�'{�+��`��Սq8�6�]������j�8]n߂XŽ\��]��Y}Ac����G>Lf)l�X�m
��~E��Z������c���,(pQ�����ɳEԨ���7_=���2�)WP1���g8�:l��=��R�_s9��ͩ�4�Z͎;�+�j�o�Yj���ɽL+,��)��j����2��[�ׅ��MT�L�Q́V��/�]�T��
#�J�عY�+˒�Xy���2��v��� -g���x�e$�-�;�9�W��V]�%u��b��3P;j������&�; ����Kf�Q�1[[�@�┠�Y�����N{},�r*kzC�ҋ���=�2T�vvf����$Urˣ�w�H�my�v�ʴU��X�e��X�qe�R|���Sp��H8�ɴ́n�`��]�l.��2���ý���9���К3K@��A�8��	qƱWb���fuH�ɝ��7!����
.�겭�߯�k���FLa�C'�^Ͳ�K�����v#�h#bR;�S��5���d��U�}Z�mE�3�(��h����[8}.��dX�V�72��ݡ3���gH�h�ܜt��W4����!k�"���l�`J��	 �}���ۧ�[�4�wY��(��!�o3��֌Ŝ�;pd�˘ Xho�f�n�y��I���p�*j��t*5����b�H�,T��WYe%YyS9��v�� ����*�AyGP�欦��"�\'~�/M5Y@ �R���֍�Eْ�WV\x��p<V���5@�I]E3J:6�°��"�Q�&���kXƜV��9��u��ʥ�@�!��˷f�&f�cE�5EA��<*
K4J���٘������.Sgo;�qg+^`1���6���,���Ž��r�/���``��iu>Ze�[e��6�-��Ak+ʳ�U[�I���t�ӥ�:���#FN��7WP�Xv�uN�\�+k�1X���͂��`��IQ�4!X��c�h能*�{�hl���W���g���R���Ld�iXW`�Ǜ����nF���gҒ�ėr�5Ч���,����V 6���(Y��7�5��6(�7��������������2,���hPm�����[T
Z(V��Zѕ+""cH�bdm�D[im�-FըV-�EQTQ����"�Z�+Zł´�F*�Z,T�q�1`��*��&5Ƣ*
,Tb�E�J�AE)ZA�-��EV1-�HT�nZ"1[UTDYb���bA�bVQFe

"Jʪ*L���Qb�QKe"��b����
�
(��ֵ��b�,U+1��,b�m(PUQUEr࠳-��[b�* �A�7
��DdDADPDJ�TF"X��Ȥ��ZQQ��X(*\�2���Ȣ��e��,[kUH�*QA�Eb1J�-*����U\h�
�E(�e�A���j*�ʮZ�d�bѭb�V�,TEDEG���ZTDA@Z���"�`bbEn%\��QDdQED�m�m�����օJ[*[
ʕF-KDT(�j�j%iiA/�[�'o;�%te:��{��̩���.�Q|���4��+V�-�]]\	�mEy��[ʶ�W�#ߣ�sQO�"WN�R�ޒt|�(�������N�w����*��w�1,1M�]��.�O�o\�|C�Y�7�e�ձ��v���+I��w���C����Pڬ9�V��u�?����=�5�졎Xv	��d�Cގ��#3I�D������[ܜ~��:
��wӪ����0ūʀ�����e�u;ڧ[�=��Pg3"y�*pb�q�eW\I�A�Y�OcYG1)��z�M�;�S,�m@�����%XU�����6�y7��< �݇�n�1�x�T������\�=��R|��.y4�^�\:�w �y���}<�d���]91�2�=�\v�DR�>�y����BO.{4���LZ4f�\N��X�p���+Ce�9��2�2B��N�{K�l�`�d\jǼP�dv.���G/3ͺ���� ��Lۍ�ن�;q���R��Va����r�\��p�]ۿQ���,SQo%u�wT�G�����}�q:��t曽�W��d*f&2H�ք��k+�c
Vq��@J�y�yR�6�:��׺�K��諍.�G�]]=J�\�t;��v��N�3�9�ۗ9��th�z�v�썾�B�z�Nݪ��^�|��q�)��5a���;ny�6i�^p�h���s�<��m���ը�mˆg�+�Fj�l�U�x��p���}�Z-5]K�)n7W&�eäB<1\2�LA�y.a�'��!qN�U��.Z���j�+����+σ���K�j��K�j;�/�Pذ�Gk�R[S���U�|��Su���T��h	�1�7(�VN�n��j�'��qÐ�;��&m���n7[��W2�P�K3
�Wvun��*jm6��c�]�u�ׄ�� ��e�ʇ���#XΐN��-�}�NtJ���}�߳��r�\Bh��{$�u����E��罺�\�e��^�o]{zi;��e���P:F�(q�ѹw0)��>���jx�5m\N�ϕ�7{��b7���M_�ş`�7�bX9�G��K%��Kg|��rM��R��p�V�T���oL��5�K�=FRR9A�ͭ�ly�sN�.�u��:ob��>s˩n�1@@qz	�k����via��n�mnc��B��{����0��ב� ۫�X�fp��1+_lN�J���|;L�6����غ�	���f9]�f�-^�Љ;&4�6����.Q�Z��圂�/�A�YsV��b9)�{i���")<<�z�َѴ��ոj2Gky���qY��3*b�=�Qs���*=w=S}U������ٮ��)U�U�+� ;�㕋{ƒ�W����oMOÓ}j��Ŕ�W�^��k�Vmy;�P�u���u�NR�\��964��\��6w*#e��t��M]�{��l��6Up}���2�����>y�iRO+5�YK���m5])��R�IXMnr��z&�+>2b4����)U��"n�]w	i��ˠw���H6��q[��.^n_��ɏ�59�;/�M߼%vѨJ�SHdR�[O�.�.x�V�s;�K}u���8���K=�!)�)�S�n�o*�x,��4�&�}����^��sN۔�V�^+F��⣏!�'bSܖ��m��$�g-�>q���)VN�NN�f��,BJ}[N�tUY�ŵ��Z|*m�����e#�ssm�<�0�=�On�-.v
�/V,����`�q`��R�}�b��2�a8�wwaG3�Ƨv���Z��k�Oz*}�]�;1I(��z��X��;�Wُ�h:Ev�Y��Nb[��n���}rS�Ords���+�n��%UO^-]�բW���V=��1�׆���%��\����oov�4K��*v�5M,�e�jϪs~��ж��{j�!��3�m�	N�E:��k��i��*]�J��l�ۥ^�:�A�xf�g���1o{0���xn���N�D�Iܬ:��j��j��CT�μ:�D�,�(���]�mUR��v��j�Yp� ����{�ms�3k�m���6�P�P\^
J;��j�]-]��
��)`��'
k��%�By����D<�z���\� �W²6��-���뺉��~��wd��J�ҩ;�Ouy���7{!CC�k[�;�꘻x%l�}�z���$����kϕS��cxS��qW�Dͺ���@Ć�f�i�S3l��l���*���v��l�vb�V�c�X�I�e�ܤ-	p��s��3�V�B�TW[W���W�!�1��G9�7�a8X����{��-�E�0nGm��;:�c�*l�c�lq�S�a0��nms����n�1��w�k�M6��\�䮜.)ڙ��<�Օ��7q�ۑ�MrCr��Rb�	\������%�{f^�֞Gk��mQS�&��Z���޵�^�K��8��g��fҭ泬������`ε4�}��Ɠ�۵Y޿7aבa�G�ާ��Imh���8Bb��fҹ��5L�_+�M;��7����V c7P��%��^�=�{��3^��N%�%k�S��՗�'G{��)�I�S��� �����n��+ws�(*�y�ø�V+��L���i���RVM����z\M�Bʂ���,��$�"���b��FFZ�X�|�l�ofܪӽ��a�����S�N���t:Fס�]q'Q�3��&�=��ɕ
lٚ��>և����׶%��B�jm*¬t�Pd3�ux[���5���)��P���['-ա'��5*X3a�s������=Mxױ�R]:��u�$X;l����1�龌r��:lk�l��t�f>��ΝW0�nM\v2��kٗ�{-5�)͍U8YƯ^\s;p�4Q����H�+&(_N�>�p�N���3��!l��_?F<3J�q���\�i����/�W�@�Cn�qMՙ�-�
�,�̩���Ot�O�sS;ua��nTo�7��zFy3bKm�Z6�E��!�C]P��H�WU����ȫ�ݲt��!�PͯG/3y����x�[եL��P�	LoB����''e%�t,��o3i�f����S��z���3q1Z��W���Y˔�H7�>�Mߺ�m�Ô�qVi��ܶg�+� Nik#tjt;r�j�:�?D䪋\&-�QK��Tݍ]P�c�ھS�wUY���ս�X��H�aCd)���Uk�E�����zmy���Z���w+�]�S��j7�%�y���
+�\��#�JO]⪋|�/u7]�d��s d}�4�>;��İ�G��9�ø�&m��郪�7SɌ#8c2�-�ѨBY8���R�����q��@?yy��N<O��ĎD-b���ވ6W=���U&BP� ��P�pN�/YyJ�8.<�Ɩ���M�c_8`�^�
��t�Ks���}td��H�s����8�<ذ;����Z}|���߫\�����a�{H�(e���mk�s+�h��x����bMR��r���+������¿/
�O�j��<��O��t�f��ZԶ-'��Z{Ci킚I[Q%��^���Z�;�T�����{�P��V8��gcv!e�w�%D��7P�����g�ҭ�=[�ԇݥ�.���Ӱ�yS��������=��}����9Ӻ���g�Q��NcP�~��z�ۯ�Ѿ����v��Y�qZ�k�^�uUr�˹%v��d�{xf�����w5U,�(w��ex�����5��ˑ���;��Q�[2eT>W��&}0����z���#6��!���^-��y\r�5�u�/+Ѳ��J���ߔ�ۆ����Ў�������P����#+�yQ'i���1M*��+i%a4Ԯ�Ƕ�w���H�鲼�㮽$6�^y`e�,����0R�
����b���.�yl��S}Ҕ4�V��t�.�Zۊ���&^ߚ:A�w/�a����e���Պ��X���7{�(���(�q!1�WG�z.{�Wś�>"�v��+�a���sw܏��3,OS���gk���/+���K����Ԕ.�������"�=�W{Ϋs1�V�^S��=T�B�5	R�e!���S�l��$���Oc1?�s��P�.Y�k4�����S��Q3I\T����'αI��X.2��1�粹�R�J�I�7)�j���H�9a�q�0m���i-s)��<�)�lWs��djgv�;���Պ��7ʡ��w�D�J)�c����';�K'�8p�N#qT�&ۨ�s�hj}����O�˟l<܄�Rne *fv�L^׃P�ک���j��-宧Q._^��:+��B�W��K�V�{���$�4g-\ȴ�QB��K����b���d�� �،��n�;�^Nu�t�wຉ�7J�N�Fs��EW� {v�;En�@��t�G=h���-��B6R�+|:���3��u�����_.�H�f�8] �˯G��h�u�A���8v	��J�E9ҸR���EW�7z38?�5�^�5�DK	�٬9W%�:�H�vt]��o����Vˮf=w�gH-a�B��0V̵�{q�J�HG�8:d�ӕ]r�<T�U2�w�{��@��^|�WΣ��f�h�S�ÿ��k�Gr3HM;6K7}�����Y/͝�jF
�>Bx�y	;�E�O�}4pF��2j�#2./<��SFo1�:v�U½dq��-�)�c�-���U�}���ܫg��j{�z�]x��[g8��Ý�$���+뾩c�X�S8��c�z�z����*�n����������9$��Jmy�t�v���0�&�<n�q��F t�4/����bl�A�xx�꼞X����,�F��r��>1��tl�JM��T����V6G�iCޱ���o9{�����q��p��*r�t+J��:ۨ|P�w���%u l�u!t��E�Mʴ�$�G�w<�oAY�k�U9肽��]�}8�1~]1�^��ʗ&��s�FjY���Y����Y��o��C�k
YWdD�j>��s����è�6�����i��R�Y��y����ڇA�����ϯHERq�,g��(tߎ.��X:o��G����!<���t9�&���̧�E�e�i��a3#�KC�ڬ�퉃�EY��骗�[z6�+���r�#3@3]�y�B�oݜ��+�G��(E��l'��c7{���Tv���ĻP:]gf����{�����հ���-�98$Td�H%	,�ţv���y
��D+g_��v���g:���t��C���V�E�u��r��Ԉ"l��$$X���i݉Qe�q,N=�:XȊ8��o�7����ލ�'��q�+|�K�pa��<�R���9�S:.�q͜�x�5�i��N:j2�Y�i��'p=j�s��H�s�
{z@U�k(ť{r"�p�u@1=6"��i�n�=	Z��:�F���/�{
� ��}�ˁ�}��^�x���r�������c��.�0Ŭ��+�ڵ~�K=#"Ӭ\5��P��b�1\u�=w�n��x��V���V��@Sԯ�?����l�c�}>�=Ctxlv.�b�ř�I�Օ�y�ʹf�(�z�v)�z,JQ���}��oV0�Y��;Y�)����cP���,�@Ԍ��u5�Cd���4��bbZ�շy_Y�Ja�N�{�:3����h]	ˎz�IY���~��jx{����y�;H@��	!I�	!I��$�	'��B�H@�HB�� IO���$��B�� IO��$ I?�	!I�B���$�@$�	'�$ I?�	!I��IO�H@�XB��$ I?@�$�����)��Ne��l�0(���1%�{���R�P,͠�l��U6�Y�jD�����ͳT�l�j�UZ�fm���&�f��[�뭵�MZƁ�J�Ԗ�-��6�5�J�2�4�T>تJ�E$�lYIDWn�UIIRU�4UU* )R��IU]�TB���nڪRDKF!	{1�Ī�4iSE_g�h)J J���T��������(Sf% D�RUEA	ze	(N�PS}nT�)
Q[b�m�J�M""J�{�A��P��   5u4�����h�ESKh
�̌
�l[Uh�JicL�`�&UF�{�RҦ�M����m�Vi�S[6�["��mV������   �    q�V�R��l���1�eMEm�@�55%T�L�Si*m���Ab�l�&jUX�2�Z��Z�*�iaJkJhڭ�)M�T�T�R+mBU%U�'��    -�i����j�b��,iY-hj6��٭e��U���B�dUV
�5YR���t���(P�@ �B�tN�

B�
q�(P :(Pn�TقT��  �   �8������\sp�B���	 �ܮp�B�(����u�nA@N�օSmP�j����r(��QIդ �eUQ@��C�� ��|  �  ��UV�k[`hѫm�4Ր�!��� -�� �
�2�JJ�X�#&P +b�*%UI)�Rf�S� ipU
�- ekZ+(+Z�������E4cl(��j����)EM`�R�d�H��#�  <  �=JUR���Z��5U���)JMR�ZH5��ش�Z�Z�TֵYM*��u�+Ce-6��Uk�)*!���)V�R�  �r��U��&�j�i[j�SB���5[)����[PZV�Tmm[Y!Z�k5KV�0
UUj�ڥ6�[�[mJ��5)j�J�VjiB��R��     3�-�j�V���+m��T��3@��V�j����jT��b�,)-Z��d�)��`���i���$��ҭ�Z�e��ZB�R��RV   �  ��Z*֢�[U��m��R�ج��X����	����Eekm[l��j`m&�6�Z"�V��҃mV�Z��[J��4� jf��%* d ��a%)Q�  "���*��   �~%*Hb B&����Q��&� i!&ҥ)� ������Oj�����oֱ�_�;�KU(s�zH���31�C���������ﾨL�wĿ��$ I9!��� IO�H@�hB���B}�������G�A���qJ��g�g5�!�f�!�O3C�l#2dP��z01��M��x��Hr��[���z�����B�)�m
Oߥ;*���E\�A^8��ӌ\�u۫C^5�*�meDa��Yݺ�MIw%������ q'��Xta۴���b�Ve6��6#���0����f
룯,�`�F�Og�)M)\i�u�G;x��ù)��w+q�WN��X���L�@=Z���;;��{���r���|g��1	��>~���<�g�+�{Gd�}�]S���@A�:��
��yѻޱu"�$��ّ�Cd1cN�"ͬs*�)bY6��CP�~�d�P<n$m˰�Y.ѬVj�H4<Q�x5��6�P�#�ޡ�{iuճQ�"^Z#*B�)z GQZj���P����r��@U�i��i�u�ÉP�� ĮY�f
dF�𭙎�G�S���rOhHܦ�&��r��oHjFY�+��tjQ46��ʜ��>;� l�2���w`��כ��)6�;W�U�K5�C4�b���4��i���cX�,]�Sj�ݰѻ��^�����#�۴p��[G&�ݦ�U�VƊ�앙ky�>����{(�=Z��bE�E��w(㨈�Z����԰��ʻצP�!PVm��8z�=�����^B��u���>-J����X)^L=��W�h%t]5�}��j�GצK�N�ɠ��=y� H8s��8�{F�M�[M�;T�M��Q_E�q�C"��E by���t��sB�XVF*bc�]K���t�ֶ.��"�(�ЙCe�x�GFǵ6v��L�Xu��`�/�<"�g�Q���N�����?&�c�rMwd]�P`�e�T��u���mT��Z��I]�F�*�1�^]�����Za�4�ۓX<銎p�Ē���|�'���2�L�ʫQ�flR���]#{z�WA�P��# Ŵ �p�os �[�F	t7od��W�,E	L�Lmmf�i[z��j#�QJ��E�7�(n��4�0�P�)1�$ae��x���da�1�bݭӱ=tr��P�����n�v�<�М�!b�=�ީ�{�5wzb(��,�XJ�E��+�v��U���Z�n*��,�`e⹍��&b0�y�BP�	�y1��9kya�K~O�B=��oY��hV��]���n FU� �˚>{T����d�N{���f�1CeD��ck%:ɒ��u�1���qݙb���2��3k`{Y�śK�������eh�t�%�X:��չǩG'�A:�v6�T����^��nqVX�����S����ӴI)i򣚯6������D�i�X��\;h�hɭ�팤Emt�1�z@ YǷw�ө��s�@&��&^ 扯X1J�Em5	����nL��Pz��n���m�����ΥǱ����Lr�ԊBɨ̭Tz�c��+b�Ia��.E+�U�N-U���(�{��]'"8s"��	 �ZǷQ�����R�-rA��e5FM�Ђ!*0�-�ǎ-��K��&䱳Qs�t`
]y�ms�W�AO�m������b�XU��G*�������s,=/wM���H�[���P2Z�p�:��C&�V�N�Պ������)á��B��M[�,�})mX`��a���PM0���ݑ8L�����}��~!Hk�g�e܋o.J�7XiM��Y��IV�:�0%�,����=9��i5*(����͉��m�����%�Uz��V�q<��yI�
z���fd����Ħ������.�6��w����d~^Y�y���4=Q�R�v^1��v����o.W7l�]7�Je�q���[,T��o�e���_Xk�e�*$��S�i{l��zC�w�^�j�/up�o���8[-��S7ѵa�h�l
�;����HSy0�"�����s�G,�"�q�p��i3��"�Ze�7�5�{��^3�>�	��7R�w��/: _TS�מ~�qP���Xq򢱼`Lylԧ�B4�jS5Lp�R�D;�ɑK�h6o���y��N�����a�$ų�*G��A.�Tt6�CJKs���w�]n�sI�X��j���f�N���݅@����.������;�e�G�їP F�W,mnR/j��o �XXe�+n6�����o2?��"TV"W���wŹEc� 	��-��v#����ugƽ붘���g���;�˫s�	���n�79��q�Um�� zNBN�ۦJ���v̛t9,J�1��>�37�O�Z�0j]{�.C`T������5*�_zz۹7WxxM@��sR��x	F4"Pޝ��[D,��>��� �D�zŠ�1�G�!R�e����o(e�sA�:��	Ь-��W����^gׅ��0��[�$�Oڊ����C�ʥ=�V��H*�[��o1���Q��e`��լ1h����x�D���b�~�����z��1�s0��z���۔�Uh\���FҫXn�u�lԑ� m�i��7���a�36Fk)@��u���i)u�m�Y
���.ZW7|ݓe��!�5�zcy/t<j�+�z�+=f~��� O��b�Bz>�(�	�
V�M؁�0n"�SXP�{�n��oC��������.�|�D����
�J����ڧ��W��ԝ�4���K��fc�W�֖Ȣ� C����}�
����srf���M8��2�Zi�jf�z��T�Z���;�7��3JuS(�֯e��2�o�#���I��b$��uY��p��g��I��V��m�Z�]����hwmy����r��21c�r^���.��(���\�e��K�_}��Ux�:v%x׽vӃ��U�J��e��L&ʗ�q�,�ey��}w!�-��y��-�~Ȯ��[)�FE���%�e�]D��G:x����>�v '��x�����Z1�6Э�Yn��)���R|z�E���^����^�Ct�����Z`��Yz�,E�ׅn
���X�<+���a]̓���|��q^M֕<����GU�m�W$������\˽��:r�,ik�~��v#��2��
lXT4`y�n1Kw�J�Щ��v�:A�FV���Cf�E�ja$�n��uk�6�B�*�+6��2�t�fLs$�bZ�I�K~��k#ϓ�E�^��>���7�u�}� �u�c�B��G�uI[�kIn���T�Ż�v�S�S�$&t^:�e�C��4��cd63FVn�Q�y"��=�݇�X�|���Ք�&�rC�sk	���Z�/v:xDz��~;�b��i��nb h=�?�gH��K\���օt)���Di�������Ṡ�D_���x���"�q~i��1JSқ#yW�c*۩-^�qݧrn�b��e8�	�"�6�A >�:�FG���pR������e]A�b�LX�*�2>ԋd�������g��(ޔ�V�T5�/s���cIv��1��*݃b�	��l��-ݶ-E���bh]\��TED�u�ɭ�E6�aJ��H�:�Q�qQ�[���>\����}�Y�ޝY��ˇ�XQ�h��ކ])C@9)����՚�L�v�y�*+�3��\L�S�!�.�����|0@�y�������eS=b��ޡ/�Zoβ�M�]xE����M��\D�.3^���H6�N0@�v�[r��`���v>@-�[;L6/\��D+RѲ�T�[�A�S���vݩ@Q���X�	*����ǅ�{t<�7(�J-Eܓ�W�"G�7�����;f3�0"�y�&�y����_C�"�׷7f��Lk�Pq�[������W/����F\�0��w�>W���S�Wk�
w�r�tϣ`KR�	�18+
x||�!�*Ӧ�Zsv�V��-S K�M��C���ڔ�b'��=2�G6�!Fh�2-���GkhI a�94����M���{��Q0bP :�栰��δ+Y�2fF���!H����B:�[�e�%��u�*;m���Yj90,
R�C��^�a��w[W�GC{�+L�OuR��ߥ����qm*����V��JD3�l��h\���Ľ�fՋ2��4nѵR]L,��L�!�V��2y.}:�[����<��;w
� KbY6«�h�V�8�'f����KA�Y�����n`�q9��,'�\_e۟j����&��P���������W��E%�7xu�޾k���E�g%�6Ɗj�͋YD^��t6"(z[ۚԴ%y��!7-Dl��(��U() '�s��zv� A��(���&��GO���Rܝ�=�\�� ~^�:ӞC������d��V	H�U�����΄�U��˩����R'o�v���� 4�D��A9O
��N�)�l�0`�T�i��N��U�-�׵w��S���BQ�(�F�y&�2�+TyN\	���`�@=�U��T�t2���ϔ#�=y>�":����tx�N	�D�R�"
���Sn�:��Hh�Opy6bA�j�G�{]-bq@^���+���!��NIwR�j�d��֟X���e	<!��t$��l���~���g�va���+��Z��[���n'�j��[=	w��b���@��x��<���]ɠw��������t��Ҕ��w
jͩmh��#�2�$�(�G*���4j�;ɘ���W�MtJ���f�����pl�M��,�e����/y؈�Oy�Ү���<T
��3�;�x�7󽽣�Q�4�����2�sL�R�l�x=�o�e�p��<��2���{����Nʾ�x<�}�>����_@�C�IoG�)��PA��������sF��+|�fe���Mi~ϗ�E�sI5;p ���3��}��[�HFj���N9�D�ªؕ�l���J����RK�]gq�v��t�A�K^ZRU�F�Y�s3�V )�;P��3jf���8�@3�3]�ܺ��x:y{���H��[�7z%d$)�6.���vU�z�V╡��
4E���n�ع��_Wh��K�<B�2ε�V�Za�	b/hh"�&jq�Wg#A�ʧ!4�ϥ�[����Yˎ&�i��Lo�=	��RP�K�X���ȫY]&'��R���D��ub�fV��_l'�V���y�������a2�(�C(��.@G�8�c!�t�"^.�e 2^
�,�J���1��J���V&�p�9^הC۹4�{O��f�rHN'�j�Ify�+�|��K����́޲\~t��D	|�w޽���8WR�,�t[��L�.Va����4�{úҐ�e+hjU��pfH�6]֙x�lĠ;=igB�fB2�~��Ţ�3n�^lzΌD�.����$�����b�=�	�(y#��A�.�jᨄ�����Mv�O\�d��>4���O���.QC<%�5��;���֜P�M�4�^V7D��V2�ᙹ�h-�#/r�3�y�@���f%�/���l��1Q������8nZ2�E�4�W�j�����֨_�D�9Db\8�����׳,+-�sn�eA�LܤC�i���k�״���t��J���L?��.�x�r6�)v�I��ϵ�d�eC6h��3���ח��{BL���~�����>{�x�6	�L�Pv1��R����!����YS��H�f�)�q��Q��-�,
[q3G�_6���Voe������'�׌��EZ�"A�x�(=K<����a���#��I���Ed횼c�̫�Ƕ�?��ۤh7E�7�����J�t�ׯ�\7#����9�(�O5�4\���|
���Gt��j�c3f,��+d�V�ck�T���K��0*i'n���!����W4ީ��zbn�8.� 2��O1�˙���cM��*K�*9su�1�ґѱ���L�K�Zk!2/��c�Q@1d�A�rB���iT٠`%V�Oy?���D��u�}�*�}�
�|O@���<k������Cl����J�"�L��@h�Q�Y�DD�Lࠒ2du�W���\�Љ�yi^����֚k��֨�LRk`n��Us1�3EB�,o0M�f�6"��,Z�Q�a��;�����c�;A��{�I�A��[c�@��(�Vd��$��{��%����Jb�!*���̙�� �V~+b�$����<����"K2���,�V��BD&��tr�@����$/p��)'����,�+�>$ni��%�>jf$�:.�\���vЯ���1P%�go����rp<⤢�ps�[k�3��п	�Ӥ�T�i�4:�����Ic!4'ņ�R&�RlY�0]�N�֨9|:��
���NH�<.)�-�
%TP��y5��ց|7��7��oƱ'x,S]�	�YJ)'֐�v6Z,�LhQE��F�l\H�[!��M�r*u��kU�c@��n��M����z�L�<�}��7�R���<���](CTn#����Z���R��i<�k���~S��e���9��{J�(w���J�X��:��@���+�ؕ���oM'�Ɩ����y}�t^�Sgi�{����̿zf��;�WD��qs�ui�O~���
׫ve�K�vM�y�]L�m��n��4�孾Q6��q�dD>2���aP�(��7�Ӕ\y��M�khk�ұW���+l�.��{��JQ�Ff⾢E&���JN����Iՙ���^9�s �DD��V��.|�B��ɇG\4.�7���lۢ����P���]-V�_ ��d�Ω�հ��Z�t���Cu0EZ3�.C]D�ʲ�:�M��S��9{�Q�6���f�'s�ޅ=9r���n�ѕw��ZǓ�)��k��HҺWl*�յO+a���;�u�������vo�xuV�G��Q�د�������pT������Z�����TVN�C���MӲې����d��ȏ=���X�R؅q{/ib�O��k���.g��E�P���I&�;(+�V�����}fh�52����5�q}2���6�.�x�w�
����$(>��Ꙝǿ2<��!@�1[���o�m�W������7��P�ǋ����><l[���3
X����}�cu��u�uj�d�����*���UѾ=ۺ��uN
*��}����ʓu���j,o\f�\
�WS:UHf��A�T:�c�GW�9�SF-��Jfel
R�?5mJA-���F�3��E,�\�pc4�2�_g"���v�z�B 8a��o
[P�o�{��M�\��1���K;�n�yE.��_e��ѻ[���c� q�M\��\���h譨iS��v��
��7GoF	"�U�#)���T�t���:�:F�ٹ��S��ŔH԰��{B��
+�R��ܥ'���hN��+uQ�4;FM�E�����n�&��뻆�`Ki��k�E*bX��1Q�^����6��$��.tG�˽� A��ޫut}���=/0�W:u���-J�t�+�c�!PS���#;2�-�!�6d��m�`1A�C��:U-դ�����fwf)W�\%�ݼ���3c�4��9L����i8�^,��.��iHu��i�x��8�Q�6�@[�EMUNޗ��˗�'�������9H� ހ�Mr�jjjv2Q�3e7�r�7cV^n���"{�J�Zn��+��T��� q��K �l.��t؋����7���٠>��%yA��KG5�޷��W=�C�h�pw 5тՕ.Z�e`ӫuM�ł	�C��<��Q����r�����|(�\m�yC���*�3��� ϓ35 �pyKj��݇må/���}5��x_�� ��6m��b����߬Z��0�.�\93��jb��Ճ��x������U(���LE�v]e�x�;���ZF��"��s��Q�K�4��匊�	�\���������Ѱ8�{��D�5ug4�Y�����O��6�:��E6�̺��N�<�NtԬtM���n�5S@�&�A<�4���1]�W�Ud�p�M�11�Vv�]���Quk�m�r�ҽ��wG&���Q��� 9�*Z��:���u=.ӧ�:��GA�h�m���<�ʁ�轭��9�n�F���uPy�˃��Wr���Ռ|r��|A��c�/�EK�U���;��%x�5\�k�J�n�nq�h�Ċ]8���;���R�*�h���{��X�������P���S�7$�t_b�Z�J�����t��/IQ����m�8(�\a7T��.�l�٪�0]�x,	�n��rTc��'�kp�<�=R]ٲ��L�Z��м|���Շ���[T���r%�%��s��ґ�l��6���yc������މY���c{xqP:+ui����A�<HmV[]���Vϴ��;���䡞���8�ў~̒R�����J��VJ��Mfi�bEABs��u��%�w����v��J���� �Ѳ��p�\j¢�.�r�WeRH:�U�G;��t��D�+뽏{{y��tO�_�[g�+Ƭmq@��ʷٹ�*����N��}yoY�w˱<OiJwR�6z�b���tU��τh�(#���U	�n.�� ���=�&��7[�Gu�e�vqq����%���5�\E%��)��Yn)SNm�S���L�h(�w,��;�$�� ��䊳}Hm��3i&�4�/0��x!�;%��k�%��Y|3K4&0I�Κ�<5��Z�/�L�z���wb�,�ݴ�!a�ĭ �ӂ;0r�ˎC֨	�t�����n�7vy�M�)�6°���Y��Z��4�im�E�:��!{�h��ޑ���JE	F�5�І�r�b\���"<����u �(�����&�#�;�t�ێ�U���º�[�� <y�Ȁ�u�Q��hb �>ɴ�;u�@廵e�|��P��5̞5��Yث�M]��)hi�y��)��tO%�W��5B�,�Is_ee��<fhj��%%gQt�kp�RT����ͨCY��ך���aΰ��ш�.�z���l@�t�:(����bY�H�.��7�o=�+6�ij�oɎ��_Q�93l]�����>ʅ�dJ��h]����z����_2�]�����%��7ip��Mj�<�A��{������k31�k2��u»*���øw2�wzf�F�M9@��s��15���Gp��e�#��4�`hk,5t��e�����_
r�%���]�-�2q�]j�ս���܇,C�p��7lc\'[�fR=��2�[�,�P%R`'��΃�����/�EC�n^g�sy6\[�7�ؚ�cm	�H��v���2#��Z����㺥�g,$��Wm���FP�S���J��7��(�.F�: g�[�H��MR4�`u���[�U�bm�S6s
:�Zu}��3��´��Eq�z�<�X�:
���3�ao��J ��wf�`�e�AI�+��Zf�,�ɍ���ef<n�
�mgE����s��4M�2sb���z.�lX��u�a/��4��t���X�+��	?���*���9�wG*���bF_j�Y��+��~(ͬ�� ��+���:���\Ů]��k*��'vm҄nMR���M:����FN�緧@�+��F����qQT+�h������f��x+K쥲��L�{��ױ���s8��[�|�05K�b�j�Ye(��2Kw���{J=�@>���[�+wsB
��.ugW}�	ҐSuv�J��P�Z��+���f���v��GY��c�YvS��K��OWijL���/��� ػ$��P2�{��o�xҞ5����x[6/�V���%E쾘+F��{��v],�=:���%�ݰ��?�Jf�@�a�1�Y�ss{9C+�N�����V"+�ث\{c������k���r���S�]A� 쵊%X�7&����o\�7LW]���m�*3Bgw�.��Ǽ�����W����m����.�4�f��Y�d�}������+�q�e�k22���N���\�s��V-�x(�Ӡ���9z]�\�.L�\/2��\�(�J�T����뤙��[�\�r��җX�̽�yӨ<�o1�eI���� ����o��4��W8��6{h �]��X����>}^{�=0k�+e��A儱�@-ۥK%x#��h��Ŷ;H�e�)��|´�+�Y��shR��r��"��c(E�'���W�DrwjӲ��	��h.�d����eiKnYp<s�k�}>�ev�=}�hDbG�}[��f��&A����Wɮa�6�e��7?/%<E�8z0ݧk���.5f��녭��ӛ��J���PnN'���Y�ǉ���m'2AJ�e��9��od6��j&؋X���_�|�
�(�-]iO.���JƩ��nS
}�A����jXV�cm������#*v��»�٫(P�ۉ��#5�F�yt��K��p���,��u��W�]M��-�n�ܫ�ﴝ�)2��
ܕBK��t	簔�6q\�T�j�i����80wuv��hV<M����n/�)��7�q-�u`��+ T�%r�g.��F,!��]	�p�ͱ��� ����-�i��v�0���^8V�-M�'�ޠK�~��\N�KK���s���3D<ޗd�.ՓCE4n���aa�O�B9������F�"�ֈT*����+�YF���_5ԁ�.�v��d�=[�:�J޲�qi� �%`���Յ�]�8*�#��5c7�e�/xa�n��P_?��S$heԣq3���4�5�g]q�[��KW2;ƣ�Q^�������߇v�Sӓ{s��u���҃�c]�N�lc�J��K�F��hB=y�.���qZV�E�{tWT�Z�4�Y�����u��憯!+���wav�B��ՑbՉ��t�~V�NW��q���/�]��:=�u5J����ܮ��f�	��D�*V�v<����vK�y�R���KqM��� �z��V��+�%7Y�iS���+u|h��]l�����a�l�M^
�|��1� ���9�@G#{�PW[҅v��,�gX�Hk5S�*���e�k2��w��Vw�_Z��ֲ(4�ۏ
zQ͍�^��'e���Í1!��5�r��w,��	B��W+��i�[ʷ�RUܓ���ݙ(�����ݕ;CЍ_aYdYS_G����kv������p�O��O�5�N�^��-�]��0_*޽"x{���|y�2�`��R�)�g"+w;7^MR7�>|���E�Mei[5���π�[���E��3I�9E��3�ft�㽫�7�ߥ͆,����f=���fǌ�<�sڠ����2�j��Hde��j�8�v9x�z�,*mV�#e�����+2�v���Xxs,�:�AA����|��О}�\��GyD�=��+��$Op�)جԉҲ5�S(Tq���t���=���)�����ri;W�5e�X����<�rg>v�,�	SY)Z���� �[�wF.�ݥ��	*룡k+������Wr�'�Q�1o^��oCs��Vh�Ŵ��t){z	�D�)H��v
�U7������/�y�y���qr,��(If�`�7��"�Z��kK�ah��z�f��ǣj�n�E�����Ay�x���t��{�Tc�jo|%gA�)��d�3Z��KwedH'������l�<�9�9i�m�[x�RڌR�5P�����Wܕ%�;�lJ�-|�g(�Onb�L1.�:u|�ҕ���;��8_'HCA
6eA"���=s^��QW�KK���2f�}���G
����p$I�����FV:T�y���lY�|�H��)/�P=���ƞù�X�0,s7{Q6�j�����ҭ��"��;C$`GR� ��6�ڬ���o�gg�@aG��w��+f�"P�uS�L}b�s��R*�{|�ҝ�.3�2�o�ŷ8T��hl��
���#z�\�k���[����S��N�^n\����d� ��m�\�a�22/XWn�3���A�!�Ƙ�k�Yܢtؾ�I��*L�c��du̾����D��C��x�t�[�b�a�@�5_\+�Qו/�J�i(Z�H_7�:�u��6��ǎ� ���*j���GY=J`�=��M�o�i-�@B����\��쑽��g^{uu2�rqSn�����{�H�65z��Al__!�2������n��U�K�u��WP�J�ǹLv�;Yډiӽ�E;�aH���Z"�@�Wc:��-�dIt��B10�ث#�M�ur��	t��b6�F1�;�<�B�ռ͡uM��ǂ�m�ʜ�6݁�h��;.;�ُz�NJ�l�L�,	V)YcV�|qWIjP��^\�/��泃U��*��KK��-�u��K
�IB���8��Y�c2��,��RV��]�@-���xh��Є�-��힔^�.��S��[|k5�0�Yv3w�jL=���r4��:s;Z��"��a�H�kF����e.Qa{צ���^"9]l��ާN������֌�k#j��& ���t�Ӥ+s�c��b$����GAu<�n%���:����k˺����a�%�r�#;�;����w�ɽ��/(�#���Ig6�;o�uի�=����8���2��o3h��q��s�qP��2Dbv�x����u^Mc��,��������;��+�I�y�8�h������AW�_]16��[�l.��U�6��]-�O(b�	����]��My[k'SbgJ�&Tˋ��ͩ�+�r5c1��e�&���z�d�}���%�Lޕ{r��5�Tq��c��A�|���,t�j�\28�nv�P���k�&s��7͌��j;�r�}uu{1x��NR�wjJgQF:���Ӛ��s��Cϕ�{��,,O��zG�DF��ljd��"���$T1����0�ng؏��G�����[�3k��R��C������(S��S
���HR΃f��ǎr"k�o��W-�>��ډ�R�]pi*��C��
{B0��	;9�iZ�)�{�I��Iʺ�ڕX�'��|ɯ���;�/�s�n��;�YE��(m��إ��c�IG����+�KU����P݋TR�e_�[�� ��R}{]6�ա�V�z9��ۢ^�n��W]�^��5/���i�4��Y�f`��i��;��uu�ܬw\��RL���ru�j��M���g�}� ,k�B���ZH�^R�Ӡ���Cj��(�0m;��{Ov�Mv<x��r�^���N�!��R{��Ѧ��#�	����6irs��Z|����Wf>���nqf��৻6 rE�1}�{�b3PO���*�!��V0�W҂��:���%��Q��Z���L��j�"��%_��!!� IN~���=ָ>W<>0�� hw�Z�AG���{S��|����]�$�R����콡MT�d��ޓd��G���gB���őm�&W��CJ����iѧ4|H�Y���U�Y�ɦ4�^Vp�G���n���L�E*��2TE}�KҲ"�eoQ�޻�-�O��<� ��7��61:r�wXf����� :,����Қ���doU�i&wp���o1+�ʰn��UU��շۓ������0�����}Icl�6K��[֩�l��\&��2�d��Hr�v�M�6�eF�Z�	�>aU#�׺��2U��p�^�_J)�M^��jKEf ��}A���n}����q f� +_3a��<)���c��p�r���n�֏lr�_ru��?�=Ւ� �;�WY|/�Z�8[˥��dx�PU�l�Bݺ��[]O&wʏm���'���nI[& ��
˜���ˡ�*R��<4�D�
�Md,�Z��E����eh��:�tr�y�u�A��Z+�5d^��O��J�JY�+���F�R�\fp�Tm�C�͹cZ˺4':V���Sm]��Վ�S4��Z]4����Y�r���n�#��E�o���xRg"�U����hJ���UO��:)�k]�خKu���j�[�*��]����\�A��ZYN�܁�â�+0N��l���`:�l+D6�ӗ����\,0gT��ݶ�
8��!2M_v���%�+�+���v]�1�?������YNO��ӳ�K�V��"J��֔�c�]�ԟ_L�S�tI�]�;��QJnu�\@уa��c�sP�SV^:�Q�WϬ�z�H���p��2�o_Ɋ��'m�ƪ�T]��=8u˝*�/�wG�_4R��yo����Y�V�
�ōf�})k,�V�v�+��g]�耋�:3�7��oVV)sz��,ks�J�	:��n�&lV�n��5�	'MC�� �VwZ;�e8�.;��R1;�J*����k���8Jށۛ:|/.���)J-�r�NI�.���e:v����;-.��V�-K4J�m������;O	1�\����|�v���+��g�$��(�D�Jy@����ms�[������}m��1�6��۬CqVGQm�ό�Rv���^ �@��B�W|�^�-Q�6�Q��Tk�%�l�{�6�"�;��ye<��;���__D8���|�H�4��ąۮ��4��S��\�Ƣ�7�C��f��6��Q�]`L�`�MV����&c'9ލH�7wh���|�U���ǐ{;U&T���/%;u�W�HK۩0�Tu�ai���fvï�N%�kU`�Y�#U��ږut-����j���7l_Y���V��82��`u��kk��!Ψ���]��ewo�3^K]�7�3��89�D�(�]��/���Y�,I��������]P�U& ��� �P�Y�S��G+7.��MU�+��`�R:ú��+|�G����~Umkq
5=K��vt��a��o�v(�ߘ�l$������ۀə�;L���B����[w�Mt�g�
��D�ì�C`��Ë�['z�{�f�WK��Tr�n��J+�!Y�K�a��iV7
���E%`%q57��j:�� ���{��0�ͥ�1���:���;]fv֪�ܐ!6l���$�/���D@~�ݧHp��mB��>]np���`�w����������9nY�ֵv��|�� U=ײ�i�g�&��ؑ��������N��MJ��A�!�g6$T�A�5��n�}�Q]��e��$ͤ�0��vu�N��M��[QHMȢ��YV�ܲ�n
DBq؃[�`�g�b�;��Q�&r�L�u9)\�fWA;��
M���Q��C��{�%<Ē�媺{*Ȋ�]�{ Vx$�N�pZg78r�7ZrW
W6Qb�����m͙B���J�6Rz� <w���q�3k~�<��f��h�cn+[�����*����j�3w�\.ɽ,�R��:#Ze�Γ*�r�Vi����&T!Z�W��s+/b�<;ʕ_w�K˂nh�v�gkx��p����ڙ�Q�r:��h'��{%ZYJ�����Y���vŨT0+��R���t��b�.�hi!������VumȨ�dS`�YBݑ,M�мT6ݲ��q�N��(����h���5�J�B�n+����U�ō�bЄ�p>�x�ؾ�w՛m�!l��oy>]�'X !���`���z���M��z�un��=ߴ��p�U��<��8���͇'46e$��`Ɉ�]�W4.�U*F�[wS�j��ە�r,z4U��n3�m��)�&HJ��jK��{&@�2�\��S��R���)�Lc*s� =��o:�ӝ)�#��r�D���Gp�^>޼{,DIP@�r5/Q�t�w��+j���W8g(�E��r�	_*Q�A���.�*�v�(,lJ�i|����-D���M�5RFJ����I	s�uPt�]<�%;��yئ`I��}ؐ@�=�qJ��b��tnN��Xs�ʘ�����o/�nr��S~R��-:�RA�ا��* oKD�3�Jc(��������-]�/�\��n�jIv((WpY�y�A��<�K������+��cV����w�G�J�^l�Օ�uuwvɺ��B=wC��hM���޷�K��{&�����������SiԒ����u-@�F��CF����Uz���^��'Z��c���>_H��h�ͭ����֫A�s*:��0`#$+�S��H�2@Zt�.�A��ӕ�[g��#����*�:����41Tmm '�އ�+r3��#
��]n��1��iNY��\*J'�U�{�>��n��v�-�gk�ۚuh��I��u�����/0�U�;״+��l�;�v��3R��� �uh`VH�չ�U ��t�e�u�e��ޱb����;�N��	���(+*�4��㈻���˗�+�mTBI��W.�	tveh��W�չ�5Zn�:AT����:\���m��G&�ph��7�q�Q|1�� ���Z�{����x(q�xb�m_-)���V3->�Qu ���cV�l"n#��)�
�����3�m���UuDsXz�e\�`L��vR���W��ݐ�=k��S��޽z�+Eڳ(�ݩV5C*ޒwH:6\��j�u�n�r���l�c�nhS�գ�؏+��A�*!�E+��9��Ԩ<tU�Ǐ`7�cD�`s 1T�b\r������sz�z��@LMݳIb=Lj��B����1�VW�Ǣz���}���0>]Xk��Nͭ�&X)��i>��:ٳV�1��MŖ��B��A����7�+UJUq���N8�lPn����u��Ժ��҇�;]�v����c&���+u�O��N�v���U�SmG+�]J$�UuhA9$[��r�Ia�C7*RJ@�@]���r�wKP	wR��{�+2����]�ªoCI�F�yZ_*��ڸ]�ȯ��dt�꛶2$�@�b��%>���s�z����m^P�>��7>]��-O�n�^�4��]�f��"[;�\�aݤ��3K���ࣲ�M��Y�`�s+."�̩��HH�r��le4*b�lt!D��)^��C6�)�J��n�����4z8V+�t�ξT�i)C3U�IQ�²�b�tj�ً��T�����`���:GV�`�>���u�|��R���*�e��.L��z��/�zũ��|�wIK�C�n�K;�{n�U�����o����v�e���V@�8K�B�w�T�X��!	�-&]�w����n������E����WQ�b4v��2�˖qb�tk�Z㋹v�K�aZzH�w�펝�^��&�N��a�h�+onS��o����P�(T΃X�r^�%�}�ӧv��zr@Ft�,R��M:wk�*,*����hT����o��*�&�wLTuD{��7���S���#��W,l<K	�mf>����|&枺��)���y�)e���U��sT�;ՁՊ��S&��wY�u�.��*N�hє�R9JY"��2���]o���D���ޮ�����X��@q$�Rf����V��s݂Juڥ��}ukZ�(���S�q�X��y�]H�ԫsۙh{:*S2�y<!�'�+5�ޒSB��Iʗ-�
�y�,�J�V��f�9�"�S1����P��gK�JWZ̗�V3��Ŋbݚ͛t$��(�wzChJ�J͕tѽ�p³�&-�X�)��f��a�C(��*��ḟz�
��[i��NwoM)�U���˧�q�O�h�r-�2�P\wl�"t��k�i3�8�<Bk�P���9|��JVMh�*𗣞3�Iȇe���z0�wm�m\2Z� ���@��w�5��mF���:�Q��W����+~���o6���)��B���w^�.�����-�2��a���+�;N�63�������\2�����"�*�����g�2�,�m�۱,�jHT�p:��p��}O�Ԃ�L+è'|�ĳn�,�Qs�WJ�WI��"��P�.��r��-B��[��W-!wÌ���&�Q\�t�ñ�V�n�Nь�
,Xa�'5�Ǐ�X��x>��77
���ԞQaad��ds�ޥ޽���kTPQ��{K���%�ծ; �20S�&�/�3'��%�{��.�6� ��s(�1}7��x��b�����a�͢�%G��VLQ44g)�o���+�"1�_^��|0�:�)�B�͚���_�Sm�*5��k�����쫷9V��S1S�!�b�<�4������1ǖ�S����:���f�n��j�d��
!i�ը/���N�I&�;%�o�*��8���i���hT/�Kk7��I�Q�&�����C�7���V;"�N��]��Х��h��Z�n�e�� Zc4���^�j�U�^�v���Pvv�1�ì�,ʸ���E!�#\���w_��n�{�2�v�[�x��z�K�����s��a�Ԇ��}��,��9�r)Y��ي��S���j�KA�·�֓`�v�7������4�U}+#X�����R�4pv۵p1f�a7�jZq����m�4��XQ4[Cjl]��쩽Fj�;z��S�T	c��ر6(�J;۟G�o�k4Wҍ��GiQ+��C��3x��=t9z�RH]m�qޭg�8,wk���aR��ɍHD7�'D茣[�o�9왢��+�v�l�/tT�р�5��
Ϝ]Cau�n^�n�����YMU�;)A��jC�P&���s�N��e"���������w]̎���C9���G�uұK�jM�����6
�a۸�,��Nfܒ�^�ǝە/B�<M\�]�P}]q�Z\�)�G�ͺݪ�`�/M�q��ƕ��5�N�TZ��l�r�^�x:�z@��q�OlB������c�2 ����)bҘx��X�@�w���&,��@�ީC��j�J{h��tWj ��yd`��eV�B�O�����Y�nq�l#�]�9Y��Z���V�5�@%����(�j����[���4��Ø��KE��x�Q�퍦��o]*����r��
q�igi��͠��G\Z�u�z�������ݡK�e�r:��v�����s����V+�Wq�]r�������<�]*��eK�Yw�� �	���J���b�,�iU�R�P�]���F�d��M�=x�U|��9�I���lC����w��1��ЖY���Lu6�`s���j����`���,5n�����W��zw
y�m��]�<��Y����;�X��צ��o�y`�A5.�k�hr�Ռ�����`����Q�5�P���ԛ��<�C
�Sy^����Վ�f: B��E����n��]oe�R�������3HR�|��)c��\��S�u	���d��2����-`T�|7�xd�Z��N2�3q��_a�y�0��������ab��5S1��n<j��Y�鰙Q�U�m��)�)�+�K���Go�ݱ�/�'}����p�'�}�\��80�������-�yf�=+;o�*��"Ε2�S@���J���=��LDU�����Vǝ�t]�!m�R�Rr�oe��[�+��W��>�Ab�W-��0���x�M9p�]�Tp���	w(�R��Yz+0
=�h��Z��Ӹ]m�ȣ���A)�tV-d��M��r��U�*VM�U���&᩼ ��Z�n��XD�ᓍ��Q�D�L�8�oh1�c��K�tl�=��Vty��W���1-�_$��F+.�MПe�
ի����%W[F�q���-�m�����)1w�h�6�_Vc�ړX�_Km��.���JC>9Z�Ѷ"�n��L�ݸ	���+s�͐�����=��՝NR������B��q6�hv��V�7�xgJ��Uї�+cU2��Y���w":n��qf��WFU�A鼫�Ue��uZ±���j���)�|�˥��8v^�ӝ[@�&J|B�#x��Mf��f�P�0Co-vTxӣܦMw��p�4`�JS��GF`�O��t�4��-s��
����N�id�锾�m;����s�}��Į��`��r�sm�����a��N��Y˛̭$�,��[8-�z�vvw={���b]%�KJ"9o��x��6ۦ�QC���%K6�`�x��\g���2>�-nқ�V��0R��7�k��"9�G"9�? ���Eл3{���[Zf~��CC��b��_օD8:���K'3oU_8nkk2ŭ��W3�����v��k7Wk��&�Qĵvԩhn��R�dL�U�w��K.���NE�B�,w��;��j����R�ut}e���}�l�����&M�.d|�u�򶺗;&�:��y�)Gl��h�bo]�,�v3�䀭����� w�.��P�s��(5VMʹ�+(�]�V���<J�u��V�J�m����e|l׵t�B;��kE�͝���dm\@*��/��qGr��b.�Pu�*<�K����W`4>(N�0.�7�4ʇ`�h�5Ƕ�r��f[]�c����(F/A)=����596f]�-���öY���&3���)K�NYZ�%W�XL(d��.�%p������ۏm]�
yʇ*�&�����a�ӕ��vB��}���]CG��ijW{�6�S"w�J^t	��K��c�\�w�hև/_���.�̷;7�,��&ܭi�6�Îg�Y;��fk�]�%!,m�h]���P��]�4��fF�t�/pv�4i�$�z�k���pM�>K{�,2���(�&��t�y ^В�p�寜��r�5��yc�|�MM�SJ���+���5�1��t��ڷ�+F*H豇";|�utY�7b�a�a���{�����r�T��՞���>j���7c��q]�Y��o��	)�w�|S�3 w1��P��1͚�uer�ܫ��۬�{l�����Dľ���� ��]��瓅���b���̭tu�+	b��y�ى�nN}��#b��걲V��1�Q�����m��KjfY��QUQkQ�UQXVU��aR�iX��m��(�R�b+X�2��eKkF����m��
��JY,F�EJ[EU*�(���*�h5�,UT�X�Y-
,X[��V*
��P(µ�D,�ʡR��ZT"�V�
���%���E��QUX�(�+QF,���ƨ(�,(�ڱJ0Q��iKV���!j%K-�
*#D(�TEUdUU����X���b9h�E��"(�+
ŕ��TX�(*���*�Ub5*
�		F�U�����F6�H[*(���(�8�"1TU�,VTDeB��-(�Բڢ�Ub*6�Qj"G��Y(*�ic�1A"��"*�F���P����""��D�U�J��mX�V(�մ*�$X���(�j*%�����h�*��*��V�\eĪ[b�Zh��"$��mDDEEXn�߾���廝��C}Ws��g2��vⱴ��a��Vq+r��6��/���f�����L��pV����ydGX�c����{@�B�9�>�Z��{����X��o�^�h���c{��H��]�)`��3�';#w9k�����$ �w���V2�[����E��r�3/S"ã���b��k���=W�#�]	��r6&�>y4ٸan\����<<L_���L:�J������m�W�s����8vic&�hN�q\����	:�#�	�B��g���9{7U�J�R��е��s���gN�L��	�;��9�';�)9���@��p�Sj�Q��il(v�F�W=�2�T��Jȍ*�^;��K�	Xv�*��֐떺��|=n�A԰�iҴ��H���4�뺥��.��cN�c\<j���+�fz�ƞ�4//Cԧ��6E�w���c��Q��fU������o��[ܽ�
���mv�0L����0���zg�� ����՜O��gg�1��.��D��Q?rk��9���˕8��ǳ��}-*�w/���2]o�+�cz�9e�,D���6Q�1."M �=�U��C�NM���K�]�����lK�t�Ԩ�(�9�lCn�F���6����?Rڎ�*+��Z���_E�z��������k�eS�c0W����]���W�G��A\�O2���̩y@��NS�2P�^VDA�+M԰ <��^�S*+��������q��8n���M��
��n4;s����vǼ����]?*�/�=d����⃄�_��ߘ��C���{9���V�y�Eכ�'���U8V�t8Ż�ŅP��MWP#<k�s}W��3�:�#�m����\NFܷ5��26�g�Dhu�<,�y����rb�����e��H���~i�s;���OV�W&6�X#����Z�yب��d��4l�Z��vxq�P�G�3���S��\%�i«?r�|��|����ܱ]?E���������^�$���خF���~t����W����)P��>�]I�`g�<��Cq��,-����v��7����������D����P�k�f
��!�!D�.�_*a��6%lZ9�S3\6{���C�xux�>/��'�󂫥V��%�(F���Y\k�cU���;�t6��RZ{�FR�j��X}-�劎�*iO9:~ v�Ubq�:kt�U�;�y�Pn���o��0k��o�#Q��$d��aE�����FszS�*���"�:����O7Wv�����%e൯P���糳k61�#8X;G;��Zl��K�
eby���nP\�ڮz�����b4�oP���P};��L��D}���ز�n�b��'(����S��l���b�S�a�,�b��1	H� vU{`�?�>5���n�Ak���z���=�5��aQǏC�K��׺X�b2�n�a�W��m�
.D�*�,�����I�UXz��C�*�	��w��C;����fÝ��n�>����UH��Ay*y�Uz�<����-/I�qVv�,��PY@��d���Tᜒ. �c��Hq�]��Nu�*�}�^�|W}E����MJfF�@z4�k�P�L-��o	����w�vX7��k���Z�;|���=��P��x��ᾛ�E�,��B�-r�� ��SϬ���=B�:�7bW�[��E��״�-�Hea�-��sz�����IéH����3Բ��G_(��ڧL��ѸQ�&�$��B�;�$ym�)^D��͙��w�;���±>��-���c��|&�}讫ڬk��H���@f7�V%a�yKs]�8j�-H5븪��2Z��x\FΩ�AH�!)y+����liR�j�Q���X�S��z���U�2G%q<&'[�~ey�r��}M�~ޑf��c��b�tì8v�E��4��[��yK�Rutùΰ⅌�z�����=vU(l�So]v��4�V`���&=3e=�=��fH�GM�O&qf�8��Ϳ)V7������Vl��y�{()*��8B�\�s���L8���<:�#'��a']���<���WX'���;1��t��ož��g�ڧ�o)��������uz��o�.5q�����=���P��Xn8s)�%�揸�9�K޾K����9��Jy3:Z��٩�V\Ş`��~��fxkV%!��#�adnQ鰙fD� ���ǫ  u`B�����%�p��^���z����WOFj��i�A��3svW;��$8��t<��͓�]{�Ÿ@��Ѫ�J�n�_���e؈�%G���*�����_3��Y�k�e�儁���Ҁg�����N�/fB�ip��"zr	�֜N猸��~s�Y�^Z�P@�{��Y@j�θ��V\P��|0�{ANh�i�^�}q��J�)�|����Y���n�>gp�L���H�9�'8w(�Sy5�J��g;`Q��/.�V��s�W��*��|���!NP,�!Ԉ���3k(W?ve���z��l�c��ߘ�5㘕udN�f>�5"ﵥ�à�kS�1���*�=:�V����N�ȷ����s�����^~ZM	:�)�CԹ�압���t�hF����qn�ګ.����3��V�I2����G8�}�����E�;	.=1��Wh�mO�NGw�US �r
�P��Q�3��:������ �{(�?<�v�I���O��]�:
�0�[��-�$�ʮ��^��_"��1fmyL����r�����j�c�G}!&0�P��^��]���
˸�ĊQr���o˪�\I#h�bϊ;^��c4����	�,yZ�]�[�p�t6�}Ң!ē���&��qOv���K��:*�����Ln�4E�;͌�m�+<r��|����`ȁV��Z�{�����AeÉ�q��69m�\����Q�����U4�����5������A�r�Z�WN	�e���8�W"�<���H���V
��eJ2���9�3���5M�������~���%��d�
��x���p�n����zs��O��8P �����}�3�0�b���:Uy����*�U�\K�	��Su�_^��t�p��7��ӹ�wfS@�o��Jɧ!j>s0p�Ւ�Q޹B5��Ƹv�LWf��q�Moq��v'��˔�U��)�^ݫ�r��b��ќ�[�+�p�=���ܡB��B�e��3�V��'Z0�|��|�\�:.�a(�c���c������ԣ��{u��+c�j�E<�r�v��s���)���m�+o{���X�5��˚��[�Ɖ�X�.��hv��e�N8��p{���E�Y|%{�������7� ��H�����Ģ1��K�7�湗�+��nj&0B2��h��t��-��U�k%��Fv���[X��u�̓��OGP]]�3��*��2����.�)�S���d�U<��������]u��9�=c٢�m�/%�GjT\�����n"�o0E�V�����9203��u֪�2b.I�����[ق�g�	u���|J7���(���d�4�u����;U�a���%�ډ��hVn�.5�r�Y)����� ���E�vbݻ�~�g��|��G��e�.W��:R:�x]�0U�jŋ�(s�!
wv��3�ҫs��۪�c$(zOE)�91�k�и�ޫ��"㠳�n �Δ��N�P��܎���[�wB��7D��Ӫ��]��|j�掿+p�~��\�P:�+'0��h�|���]�D�Qga�����02,G��r�EiY.�\=F�[[���P.�s,G�L��qKUF�8�Uь<�,�X��R�45g$����*Vu)ԁ`y��_+�Փ�o�d�1�Y�XѼ��`�5x5�<G����h���s�N���`�t�;\˼ۻ�͠M�����i�9_ĒaP�N��4�^u\��{�7�_G9jCMw`FЭ�P���q�G-3#���RsN^N�TTh7]\�7˔�9������b��o*�^�Q���Ih�r$(�%�,����`��ND)m�zϛ~�n���ݍ�R�o�M��Y���T̤HG2(O]2�78꧹]yK���@}�q�ɽn���'wvM�7ٸ*3�%M=ׄ:q���-MD�':��W{�O6Zk�6c��� B�IJ�\�V�dך�+��R����y� b�U��Z}=����t�W�! Dz䭛/����t(���M�T�M^#@�!���۾X[�m�yۛr�����s�m�����ٮ��G�[^N�����3X��@]ln���f�ȯ���e��hz��)��Ō�j�� 	�7�Y(�8�Ӟ�T���9{�碩�~�.�|PC}�dЄf3Y*�!T���yq�L\mb��L�B�D��b�j#^N��A3a�ȝ#�qpp�M٢ߖir�}`�QZk&T<&��H�Kb��,@$�۹�2��u�2�W����I8k"�gGE[b���qg��o62��`h�w3,�+�
����Z�^���A*�WWn��n����v�3��&7j`��}�:��^�K��S�T����Dqv�$nu���=�)��ჅK��CUYɩ�n&�C��녃5b�P���w��m����\U'�;�e����*��8�D-%�=Ƞ��͍�� �":u3�x`]v�{y���ʞ�
��V�W��V�rc��|�m�>�k��R�� .S�z��$��jx�"�X�3 ��vA�]�VHY�A�h�>����b1H�"��{*k���u�&_e������@K�_zM�;��+� ƬU��Vxϰ�
�$x]7��z����V�oy��Nf�3�1�>�p�t=�����W��7���!bߋ|>�#�k�r�=��A��CJ�H*��**(t�dWA9�W�5<���S�����$tZ���������a�L���hm��|��l���z��<B��T�e��09��(�Ӊط=�k�x�Ԝ=�'rb�k��������)]=�@���in�q��"_D���2v{/���o=�6(�0��^����Ёt�u��ܨ��b��^��~��n�7�����;D�/�OVn:��/7s��r��,��#f�kE��̡�,�2�Vu^;�O+e/�[IY��u^�:�[��9�Z�}z�3�yWw��_�m��n�+�h�]�si)
�sBW���ꣶћ�u��9�Jذ����{�-��F�ͫ��V�U���}]���*r6���@�{����;#|F<��3B�p���Ƌ9j9s7�!N3�j�j>�<��Gr~/���1 ;��J a`�D�j�qWzS���a��I���=����ź:������(FP���x��(�-�#�N*E��i`�ٳX�9�|]6���͹��v�L9nD���b�F`�����>�屜����{�f��lR�;mA[��Kz�8b�_h팹~'׳�R�=�b�,�!�DAj���<)�J�4�f�+s�y��<�e��w������N����FX��W��b�Ɯ�� ��'9���ѻ�Ib*��8N��G"N}��z�v`��&׈���B���ϖo7�f3O��ݙ�~�aN��(��' ��'"wٴ�"\��q:��2�ܒ%��5\�Y����������#��x�_�v�=ZlF:��B+�A�� t݂7+��yw~������w>��K-�)W����(�3��b;o!Y�L��.3�-�u�{����!j���EʇB>}����o��l�ʎg�>��y�;y�+��Kdr0�Φ�ސ=^⶧�lv���X���m��{���~�o_�=<d�}�x�		Sȝ��7H<��8S��Q�;����@>���i1�'a�PW"�<�₝��}�5�+�����H����N�1��ת�7`���dK|l��־�i�Ft����%C!W_@��kYy[�әv�wktu��V�´��2љ��!J�Ұ��)/=�d���J���W�x]�}�;�����ssN�Ю=���0p����xDk�vJ�'Z�c*�,��k����U���0�E���%R����?3>��V�u�EzqVA�J�1Ր�'/z��O)��b#�Ď�J_L��v#f��	��y�R�g��@L�A�}x�淅��7��:~���ܾ�*��6tE���Yp �DB��3�y�>J��n�0���DjϷ�Fh�Te�Ne��%'6x�E&�U��6�"rz�>��3�
�}�@�t
5�>�1(��7����n�2z+���	:�q�Ћ#k��n�g3J��S��m� ��8��3ܟ�k��|��)�ײVL���5
 3�*^��X^\�p홅�mGV[�=.2t��헺jcMxU��ǝ��� ��v���n#J�����B������\�sn�	|���:�i3:�o�*T:Jʺ�ݫ%�x)�w��p;+/�LIr�y
�iwo/������6��S1���d���Ć��d�fλC7e��Va[Pk��O!번[;!Q�fo�ڙ�k��F�������X�W���rja�m�t�<"|ி��c'u��@@Ʈ��t���dͭ���=l3�WK�K�ΐL��_t�qo��)�*\t̼tt���xv��+\-����8Hۭ��١cjQ����g\���6���m����+��f:���Q�w��uc���d,rǂ��"qk���Ѷ�]l�s$������_���a6�*�P���i,Ǆ�@�;�%n7W�d�(��T�Uoy�CCe鱙��^˱{���+DG��.��Ewr��n��ޕ����b���L��X��h�v�efv#d�����h"�� �Fۡj�. ywHZ�7n�\;�@����vkV��|qa�b�h�j���/��#G��n����r�R��Q�q���O��s���U��^��YK7�0uF��L�|N7)��X˝[�.���x��چ� ��jQ;� h���ū7A��+��q������vQŝ=�i�n��A�Q%�X{�,������}u��W�:G�4୬\`��[ĭ<��8;���;YD�z*n�Q�ꂡ��"�m�۳}g.Y1+���5~	.�'��W�=P�����r8�c3���	��b�u�nH"�b���ӯEP��+�:�X����4LW�q�+���e�;c6
�*U�/��&;�,h�-�@��s�k&�`���rZ$�
dXŢ��W��G.kA����t�E�VAj�&a���AS'��F�u�W��u��Y��M؉�C�8��z�z��%�B������Hȉ� �������pA��R��nfn	��nf^1�r����r�Q�0�,`�~�7^����jq�v��[�KAk8�I͖��@�Rb�fU䦢D{q��n$0�%G���Ƕ���ñV�����v捂S��G(1���X�� �"`��;:�B���4��s�ގ��+^��wE 8�H�����c�׎�dn�a՞3fXܜ��8��Y�1w7%1s1*��nֆW.�l;`0� �6; �G��0���.�+�貎�Q�6�e�f����rlUb3�iB�(�5��e�Ōih�����(�p���Z�dV"*�[bVŊ,DQb�l,UX����J������b(���c-
�iQU �b
*")m�b���R��*,Qb��DV0X���"��* �J�b"+V*��%�kA��*1(�ZUcZ��UX�*QA���h�QDD�A�b��Eb*ȌDTQbAX�*(���PUQQUFj,QL���Eb0TE�-k�����E�E�(�[Kkjh,bDT�V�b Ŋ�*��X�#US2�-ETTX�$FҨ��0b���0H��1Q(�UU"*�QTTEAE"��TU"����**��E�Q\h�"���QbQ�1EX�[X
��h���**
,DQ��E��H�QE�UDdUQT1q
��(�ŋ#H�F(֑TX&5�jR"�UU*PQQ�`���TVV��E��U�V����(����J�j(,T������J��+�1E�DF6��TQ��Ԭe�Tml�AT���U�R.!E����n��ߛ���[៍�8��"̧��ھ�=�x	���{Ά��6C�X.��: ̔�ÍA���ȼ�9[�"���Y�Û�%,�3zc�#s��_]Ǩ|�����4zj��~>G^�;�X�96nz�C���3Z�1�jB���^[T�眘����i$�ϻ�"J�^^�-_ .�z��XS��G�J�c��,y�]��b(Hv�wv^B�g#k�����;���Fɩ�e��Mn�oOn��ˍ:@�Z{���|����;o�x�ς�\=F�kk`>�=<f�Q���:����%p��ѐ���ce9���4��U�����ι�xr�Nk��J͘\^���S�KQ�;�b��\s�**�i�9���U�+p�\*�:�xo<hp�+/�����]�js}Δ�~�s��ni�|l��_2OJ����V	�n��;'�e��ĭ0eu<��s��o#w�.m4��6��^�״�z�F�;�Q�uW��D�ĘEr����7΄Í PH��D����UGخ�IǸ��
���!�t�^���ΰ��0 w�碭>Y��-�:���i�"���GUml+�/��>�P����J���3#�Vr�+��+���ڇ���r�dt5�e`ʑ��h7p>Jۭߧ-㕏o3Y-��X�4�/g@�c]u �3y�1�QJt!�B.f�Q�u1�q�/���,.�07�t��[ag]�<�Z���%���es�[�4��oi�G�g,�u3�vu6j���J w~���㋅�w_�r�,��,��
e�  V�W��p�k2���3�l�h-�7Wj@Rv�� �3Э��}���wV�-T�Ǘ�{K�Q�bED0�8�T;`�B��J� �\ l�]Y�^�5̲߼�C<�e�a���1�c`L4���n��E���s!�C�`�	^��B��m�U���[���O�{8��~B[]����~���dXj2�(9��Z��l��]Ѝd9voVj|J�QIK���u��2kH=��]3(���d(1��o�66/0��U
���^�XpЊ�e+"���G"�oq���AF��ʧ��G��Oc���/��C=�[��w����ה��g�2��@�,{�@{�"��9��q�5���\@�v��[�Ƨ�p�����H�Neޟ���%׽ܷ��!t�w%��(@9*e�%�f��Q۬N>ح�~�.�ifRb�e}׌��pww��[���v�t$g�:���{Z:�e�w;r������[��ǯ�����i-LF"���o1ܾ�k��X���$۝\��(�s�pΝ;�(^t��S=�s�+3v�t�Y\�d�UeE�H}��]���A�5�_*V�Q�}�S��p��5-ت�78�Z⯥D%���x\Tl6�-��������dB�|�<{Z����"q�fV�]�[X�uV�M#`�t���}��V�n34��m�-�X/����,Ș�:�we^�-o��r�DS�0O�[dF��0Wq�7�a�q�:%�'��4���������])xyv�\�X�t�ٞ���M��� �j�#v+Y����`�{{��k��e�|�ʻ�2�/$�Ǜ/���]���/J a`�D�j�qWz7�!6N�u�:�����*w'4���z��������'̡��q=�P�[�C�c�x;5�ێ-o0c�N�VU5AX9T��r&TD7N�/T��=@9�k�7�`!P⧗2���G�X$��1�B�8O��e�8'w���:"�L8؈j���*���U��H�ܟZ�̫p[���,��E��[�����"�9:�̩1z��p�Uݹ4yv��י扢l����S�Z̚�y.�Qȓ�C骗	0XC2��_��|/�:ņ;��noM�6�P�;�=��sy��G?���d(��aX�T�FS�G��Vr�}�V�gNS ^�t�m-3M�5��b;.�|���֮D3�IY�X����Z7�����[*L�q�t��ș��}����;.D�g��a�����+B�,�^��5Wf�ꍅe��.���|;���%�a>ͧZ	Y7��i��i�o"�,=��^l�d������W]V�
��D\dO=z��&K��<4C�Ȉ/�����t`��4z�L
���&b�˺1)�x>�N�e�7�Lnn{�i[�%�F�
�,`�Q��κ����_>�~l�}u=+'&z'#!��T���}���KaC���b�A^���ΏEt�E� �Mt���=/JY��3���[��S8�x	6|'U�ވ��,����|֟-�I�F)���C��͠sR�}R4���[b��q��̞S��>�Ҳ"� ��Q.8e���MWQ,{R;�ayd��=+kM�p�I��2���t�Z��t ��A�[���N�}����c��Ş���t����eg���*ϼH�.���f�x�=`:�s�%֡��êM��<�=�y�9�s`��C�>H��X5؍��n&*�f�!�� �@H(+�=���7��~b�֧ĪC௹�E ,�.&K�k��2��c��c����+�fyI�U��X���[t��bEor`�k�I�ŝ�֕RZ��oB�w�̄A:���J!�/]�f�]ԍ�e��\}�/�����#_���j���v!�MN�y	ۿ�S�١�r/�%¯>��S9<T9び�>�yeӰj=]�3��z��&�DB�c.��@U7�������:\��J�M�	�z"T��L&w��p���,�J�S��=�
�|��J��F�gJ��DS�/El�g��a�oS2����yj���U�\uv��=�Q�Ϯ�C�^��C�W��������)�W2g��pYG6�5��ާ�j�!���4�D_��i��rh����q���
�z�`���C����2�W�e/�kҫ��������:��@�����&�����]u>k���g[���E��UW���_J���q8P�W#mz�T�L��w�h����m��[����ΐt�vu�g~�@lW�O�iQq].�J���kk`u+�� ����s���������u�n]�U͎��\1��3���}�
Xs���:�rnϵC�I��>��=����Kf�{����_]K����db�B�S�����C��Kӷx�,�m���B�<�[��{�\4ͧ��l��7^WGl���ǳ^MO�dh��4�\��Й&����h����W��fR;G���-�����𹹔�]n�<�+l�t�/��_�LώV����l�R1v�Km��Z2n){��9]"�8���ǖT���07��EN�,5�����$��n��j�H��)�L�'��ِ�8͢�X��Ns87a�۫���=tT�S�$�2�!q olw
���>=]��ϓ����k���Pw�\�Oyn��� >�w%�vGe�BRN&�v���������d�~��D��L���۱����y���� -����}���Up.j�ͬUx�'Q����PkB#��
!���}���a�p{��[Gro�G�Dg"sǽE��]:�H�	
noI�Qs�``X1be9����pp��"3;<H%y�F�"�a=B��y�U:<����g���u��Є�]�VxW�anq�^^7)�[�����mAb��TBy)�׼��"
�4t��S'����i].rm9{Vn���<�+#�d7�_�������	]>�g�=B�=�A�Dpsq0$���t*[�jٱqbNVd�5��=.gr@��w�&Q�:d8���Zluј�4���˛�L|�Ӧ6`'n�YM%PT��wm+�d�s���(����ƴ�&�,���
]Y�����v�WE��ս1�G���/�3��OT[��~�%�vY ���Y��z��j�7z<�ۧ_Jk����R�wȯnf�������2W��ǂ�ڰ����vj�8��<���{Ŀyn?]�ȖA�s���"^�0�$U��IӍ٭�ee��vݯ,�ؘ�]����c#�Ț��e��B�g��VA���g`+���yw�R�dF!]��;@B�8L�*Fʬ���7����C���u%wY�
��׌᝘��HX���|>��􅇎+���tA���{������P�\ t�D렜ߕ_X��
|LO$k!BKlOe����R�X�;�9�W�������# ��w��W�+q�4��a��R[x�^�%N�̮�.�N��۹�dL1eTB�:�ؿJɃ>���Э���|�꥕I{ô�A�˴[~u��,�A�����!�eҢ4��jm��
z�*p�c�@"�*#�����lS����*�\�z���m������ύ ;WTH���@3�(L��/,����`N!���ȭ[=W"���jy��^����<�Rc��1���xϭ�!�ι��{.��Ѳ��l���5�4�:���nN>tq��:ۗ�X ��F^�b�,V��k6NN�a*���0����]m�[����5[d9��Lߝt���-H�F��3q�d@9ef�0uL�1Wh%�P��/H�p ���9cgeMX$wÊ�b.�7J�B#S%�� k��W[O��3�R﫚Ω���_<=i��	�f`2L1_���=�z:T۟��=��a�A ��Dd䶂�r����)ț���`�Y�gh(s����7o7u����7�o��"��X�>�� #����b��ntE�*"$5���5l�r L������{�1^��+=�v+�����:ާ���E�s�L�(�c�ħT�}���ao^֙"X�����1�o�b
r��t�Y𩜬��:�!����*��mJv���^�)�^�tgv�L;��9E
������\ 77	Ȟ���P�U$�4l��U�(��j&��Lv�~ �l{�g����yj����@��E��ÿ�������B3��f�պ�@�"{�DE�F��UN:0��2���f���Sʪ"�o��0�@f�瓞�ə��׫EwC�c�&�V"��AC���@W�DD�x��G��,��L�$��ܶ[s��Oc��}ucEA^��H�zU�r.+Pp�����VB>>snsO̊z�� @{�F`�X�b�<.�[�b_o�c��U���X�7��wz�F-�.�z���\.|�IJ�M�̲�X�q����-�t;;�G�וn���d}�l����L�=�tx����̬�����O&�/�7�G��2m�J�eH�FH���YJo՗Jd����8�	���ͻ��۠���p�Y4���dҋ��$]y.�۬J�u��Ar;�Y�X�a��"�U�]���%]�cQ��1����O�T3:�B���)g������o�t3�vg�Փ�e�F;��Aq+������6((gR/fVk�4-����ʚ�h���O��!oGw�����*��˖�t�K���uv�FOx�l��X2`�d�QU)WS��w��Ҷ�����񣣲���F
�j/gD(�\��\�w��̂y�By�r�^�8�ɭ��Wb��D���	����DQ�V͆:υpw���a�b���F�gZ�&f�{�s�jDG5����z*99�/Ԉdj�ƭ��vp�����s�<�ڷ3=8��<���#���WۓFx}�8�z�`���l�����ڷ�y���C��RhV@b(�]$(ZK�s�Ll^���I��H�&w�yi�j��N��uv2��s�mRK���7tb�뫧2��ΰ��8jg�7,>PaL̠�IVowUż��6���ۛ��ig8ow��R�*5�|���D_�<E+�l(�D��oII@�Jsv�U��)���C{���jj�53��U�/����z5^�4�kr∼��N�u8g�H�TAJ�@t��P��6VH�ˡP�b��#G��-��m\��t���0��-t�Q;=u��+9X����̜���!���e�0�\͖�O<�7s��9q� ?weK��͇G2l#J�^����s��
Xs��].����q�=���O�p߸�u��Vg�Ol���d��E��P�H�K��7���[y����!��Ɯ����� <w�̓��n��V�a�I=�h�f��� �6{�>�����f���n�����q���pn����8�뢦���I�l
���bPwGN��/[wXv��+��b��9#NnH�M�F =����L��-�ce�q¶1q�\���/X���� c��`��i�
�:�n7R�9=������Σ���n�ў[�U��+�Γ�C�B� ZЈ�U�g��w��G/,����Hq��_[��x鶗IW�.�&{p�¶�`��D�j��`i1.t�8�� w�ʺU��}ck���SoM���$��Ƴ̮�@�F�����ދY�3�s2ԠpI:�����`����=k6��4�=�U�m�<:^���Jv�g��9���Oc��gl�(v��ܜ9�4�Sy�b�d�m٣��(�*+)oL�7Qʗ�ʻ�;:c����V��S��C39,&M$���%|Rp�$�e�r��iù���[	M,c�u���(��J�v��ToGc��5�{�on�q�*�>B�X�νn9*�/��ٮL�;T@���[��bk.�8��P�oV�n�1�o1���YQhŢ�ΧϢB�d�N���ᦐ��B�v���P�gMu�X���^�f�X>Ͳ�×+`�s�2 ���Cu��E��r�:CnDsl�lA�wi���4d����9>*��#%*ؗK�����#Xx����ī��'Wtήm<���gk�xЬ�$&��,^��kg�N�]�Ɇ���/���G�!�`VN�2�q�V�3ZVz�僓"D��а�vjk}�R���'$�(5GNFFR�Kvr�%)�&�X�Ȯ���l�M㢱;[x�)���mÝL�l����	ܚ:�m=�6;{���Ots��qJџ]�|66vm�dR'o׍CY��A6j�܈�{�͆�K��׻�F��(>r�Mt�px�5���9���\�' �Ηj������}����iR�>[��
���0�׆�u��j����D�dx�� ���j>z.���ݸnv��F�Gh�d��@;A3�SUz ���ZU�0�e��;1#����7j^`�˷'%��Fղ�-{��;@q��
�<�n�Z0E�%# ��
8��*���ĥJ�P�m+f]���.��K��Vv�Ԙ);���
�����8�^17Dp4h$��f�ۆr�5�N!u�i����
j�-˥�d��@�XwpZB�т�&&jbq;&N��T�'�B�U��/�M��*v���`�6FWNX(�ud��_iP��mmD��f�r0־s�F�!�ލ�u.�w�#ј+:�X:j�+���_V�����r�k+�Ȇoup�H7YO�tz��XVd���zK�)!X��h�L嵚����#�m5�5�F�y��w�L,�SZxpj�u��D�ǣr��pЮm�i ��ADv��{�O[*��y�����n�#��MϠ说��I7�ʮ=�q(��ٙ�d{3�ڞ�q�6�m�

�h�+�:gҴh�[*ec�V�Q�N��1��Gַ&hu��}��0�ÿf��dT|	>?/;.��C����$j;�v���t��P��ihv��U�j[�A��g%R���;�zE(-�X9j��	ݨZ�o�Wk�{���[-y&h&�u5��	ʼ����K�Zł���9.Z�t:F�m�[�yEj�M̢x�5�z^�TF� �̂��'s�	�m�ʰ��}�i�1w6�������X�<�Pi?������:�;
�9g�]�����q��xm�U:X�ϯ�f�c�����->�[yeh���[V�]��x��c���[�(���n��,pO ��qW��X�.,e`�c/�=K��M��CmG�o��T�m*�m�X
�1QEUU"*��TF,UEU�*+T(��b��Q�r؊�Q`�X��H�Q�Q#�-�V("�V"��1bȢ�R*���-�X��(��TcUADX��FE�*����X�\�AX��EDW)`��+X�b
֌QEQUdcŖ�PPX�F���UE+�"",1
�k��DAjV
�G-ERe�Q��1Db"��b�QX�0TADkDDX��c�X�PU���TX�������D\����(��`��V**"�db([Vѵb(1T�E �b".R�UDUb�*e��
�EQX�*�%IQ������B�a�X�*�UUD`�* �X1QX��dUDL�U���2�����(*��,Q�؊Ŋ�"E��E�V��	*�TT�EX����0X-�0�"1D���EATA�X�X�9j��Ub���")�(��b(�#X�`���
�V�TTETq,b�*+No�~��~q��~cu��zT��ǆ��h:D����VoQ�xk�����j]�Wej�:����j1Q=p�%3Ys������[|��Cެ��Cs�0!Z0#�h��IBt�
�و�0��MG67�/�
b��3Y�[�[6�l8����H*���ty��"��zS&����֐
��<���=��8����x�j�0FK�]QAT��.lC�4J��p��Q�b���s������c��;�	TD黜񮭇��\d�P��!��e��L����$vc9or;:��O�f�ո�%H:��:$��^a��\�
��.�1�3��'[�x�����=�O&��/Z� {����
wdd��[��GDc�\@�YNqQ7��{/��������l�R(?��M��=��ظY3��W��RB�b��w'\�82��Z�fj�c�B��(X��V��E�u3����6����a%�c#��w՘�8���T�GWU��m�#��g�ru
�7��c�K�t�Dt�����=mQ�˜«J�r� �FJ��i��L.�`i��ԭ�f��vm��R5�G����d��&1�TDX��Y;��q9�X_b�ťW��GA�Яv@t���Ӄ/zݭ�H�xx��hF{��a����sY�Ú�<�K�[�u�zr1�]�}���m�'�	�<�[�J�&kq������gmZ�"t-��{� D�X��ۿ-ņ����X������c_o��]�[b�(d��sԙ���λ���N�o��-��@W�d_��)M����Pmu��±�J
�w��Bl�9��^�q{y��/��Z�E��1��^��4�Lꃒ�F���@3�D�O�.Z�c���ok-[\�$��U�B�ҁC��*%���N���Ltz�0�^I��62���{vҞ����=8�
�~�@^

�:7U�s�9*"3���b�J�\͂@]��s�gr�槽ɒ�\��o2cCLο@e��v-Vuz�x�#��>�����O�w7/V����G��l
 ��u����c2�g���1�ȅ1OƗo��ey,�Ǌ,{�$C�q��
~��Z�1��(:��@A�>�IB��t.�t.�9k�Jq��;i	ݜ��T��w��9��o�΍���QW&C��r	�95���ii�)����z(�]�a���eީ���y~�4<�VE�����DvQ8p}�kwU|hg״��H�I[w�Zݭ��~8G�b��>5h߀���Q�1	]�#B�z�uJ�6�ް��3,�L�b�<H[�Q&^��Ĺ�p]��+[{����^�u�+w��qus\{����rs��n>���A����%��=�x�w.C%�؏����bO�����ЄgV�b:D8.t�1��e�
�v=��d6���n�VK��{��N�Ѫ�<O@u!��K��n�#�X�T8��y�**��s��z�-���N�sE[�بC
�	�ry�<Lt���O�QWn�!FGw�((|�N
�3Vu�4b��B�s͡*^J�P���!���$�ʍp�3��O~���l7�3/�X��T[O��ᑆu��}6�o
�P4�L��P�aR��*",yM�%B�'4��WA�l�����a��$�y*�*[F�Уh:�r�'�i@���y.���u���8�@���X�Ѫ�۩*
�����r|/�+ˏBi�;�وPD�k6��r�WgE��o��9gn�DB�pX���� tP;��U-�^�uC�y�:\��:�ǫ�o;�G���4�B��!畟=��>F�\h�r���u�Z(,��㩹���Vk�ݷ�צ�ɤ:hLEj�94y�@e
�`�[��&R�oW��X���>C�V�ԝgf����{��a�Bt�N�V�iF���"6��y�˶i�5�ok��W��m�K(�{�ek��kK���$�,��;p7�k+��#��b��̱���Y����>�%`��qb3�R��wYFN���k�:���/P�K8�p�؏K)�93���-fFղR�U_}��U�ƹ�4�D���~�)��
��Dߋ�4?�k:}咈���>u�
��5����;�>�睷&ga��54���G���� =���O��)Ak

�!Hfka��TH�«��oT����-}�W4i'��/��~��e��E��B������	��g]pdd��#��Ů^/KH���u� ��}��J�u���J���C������pm�ӎO��}~��{�Z޸=hER����ٮ�P��y���t\Z�����3n��.��,b�{�!�3�4l�\��vz���eg 0`��U3' 9��/�w�(q��~{O�N�y��]ѯDΙƬWa�j����S�1�6ߴ�zb9Vр���)+nc�Ö���fL��y�R����ѝ��ѵ}��8O���x�U�#Ȍ��.��{�g�KiI�`��<�n[�F=���}����\l.�|�=+�����c���I\�Mef�Ԯ����JC�񐍥b��2y�� ���~utX��*mOD�0V	B�LB`wIjS�Bivm�
�]�m�^ANK.Z��Y�4�]�!�ñY�/���ɸ̃=�0�M�EnJjf^���E�c��f���͘��Y��}�eZ����̮�쨁��\]���:��\���D�Y/_[�\�R�n=���Cb��MN�`���}�U}������ OƨPxp״��R9#�[9��OF =����NC��*�D�\���W":���w�o®�u� )q�B����ţ#��h�;�/�K���#8��{O���珈��9��c���/��	�fE�~!E �+���M�%@e��̝^+�n�]F������L�)�`7@m�Q
ȍ�U�U����E��'�o:^��{q`3��&)��o�Qv�鑐29�U�f��: ��=�1z�O_��p�=}�N
���"��gnqdFta�!@�:�ڂ	p{�TBx'���d��J��nǮ��������W�K����'�k}�5O>V/=����
�I�#s� &jj6�a�Ȳb�s:�0���DG�H��1,u�
�vn��m�K�j�_�zjG�v%��˸��p������g��ve\Xl�$�ڡ347Hu��QȤ[�7��6�q��g{���(x�����ފ��|pt�v ~�a�h�\s'N7f��y���� 9�Z��+Xl�� X�5��w0�e���,�7B���E^y%S2#Y�0k0�;�StG+l�;�4�š>Mgv�s�0�Ν%�\4S�!�3U�&����h㗂+tnu�S��҈<ye��+�]�+ςz�<�+�fZr�VZ4��(�/����m[l�G��^�/xRӕK�G����U��;�w�kf���oX�@�jj6:i;l.�㻿����⼵KK}�r�]{�2�n#�K�*F�K�\����ccD,�����P
HPV��'m�GaW=�: -����Q�E@�H�į lX�KrT�NBVL(ʷ"�1I��nVesO��ih���l�~$��������[N.,C�ATG9�[C;��������+����z4;,/<�~�X�l
�=�
&F�n:��n34��m���_���/�i��qQ�[[��O�@p����I�B?o��s�4��ոpX�5F�^��f��hS؆Jx���`F�<E��`�̱�LGN�r��H��o��Ly=�]�3����lR�rXL����#hY�Q�l��V����bZ
�D�ñ1ڥmNzF�ݵ�1���!���u[����	����z���X�P���܇��7���K�����5�߽�D2wa
�v� �ǑLD���^
=!͓Ӟ�)�Ł."m嘰)U31U���Õ�8�e�~7�"3L�s�\=�VѨ�+�/=F��U���=��Ⱥ��qAxV��M!o)J#.��	N�1ۡ�vz�6�3N�p�y�v�a<]\u�_p��;�9�3� F��V�;ƙ�sup�]:�s��_W�}/$�K^�~e�t�����L�+��̿�����V�}�!LS��=sޓ]�����ڶ��c�Bw���!{���I&+�f&�Ǯ�a�-������y�=��o��Y;0xGV�Tm�����󔺋a�Z�d�]���;E�c+\���对\��J䀿0��پfDKs�L�<�q��d5=7ΪaP�����-tgZ7*
��o#9X��\b�VD[�B=*"�no�S��|n�<ȿP�Ln���U��+�R�]o*�O�Ct���T���.�|���5P���גW���T�ڹqļ��;��9,��A�<�0:��j���l�Z�Z����?��~Y�>a�R��Vc%C�x��!] {=�gY�Փ�Q=��|�����H��~�Х�g�\��~��,?5��6�\H,�}�T���07����1a�P��w�i񓩈/٣!���c=|I�K�&3���q�C(/��x�H)����Ϳ{�kξ3���d�Ųu*u�����d�I���s��q4��PX{풽jAu��u�yd���=�OX�����S����Y�AN!X��>f3�ua��~�Ӵ�1_ױ�Z��C�t�@�� }�1&Щ\כ�����"��8���+�x��r�P�����=`T�![�8ɚ�`V{|ʑb����g���:�R�����X�������Z2~�.�&�����
[�R�\2:yRxt`�Ѝ�leF1��؏���L����/;�0(�W6n�T3$ �t��/j����F�z� ��;������� �g>��i�ɽt2����}�uŚ]�W\�ӍN�-�Y"�l�T��
7� � [U�������ܺ?���M��+�*��7M�@�+>C�<9�%H/_X|�!�z�0��܆���1�5y�`V��J}M=d�R���oퟘk��x	���H<&<&ϼ��|���{�|����5�P�8�^�2�T>�0=M�HWL+>g�wVO��0*�N��~v�Y׆�4�>OɌ�����?2u1�?!������"�#�c���X����`:�ܸ��o�~�3��b8S++�:�>��CI��5�RT�K�u�B�L8]a�R��39`bOP�Y����X7�1񒾵���4ξ��>����c�����ݞ��k �h}��>|g��7�v���`Wgu��rVV|�!�*�_��s{��
��E�a�R;� u�|�_���d�R��l������G��oc��0!�~5#'�u��(��?x�d�/�
�g�H�C�|��߾�8�̕*O��H-@����|�M$���ʇR��s&��:���S�(bT��g�8͡�mg-�z��1�5�tx}�~�ۯl��Zr�ޮ=����޿��ߡ�%g�J��8����Xi�h��ܟ!��~��1"��y�yuĂ�d���O�9�B�g7�&�Y�Փ�^����Aa�.!�H)�?x��s|�y�������c|���Oc�pՊA2|��
�`u���3L���}��?��J���9��aěB��]���:<d�
E���8��B�Q��@� }`8����|�V��73;巯9�gz���8�~3jO������&>!P�2��K�&:������`m���_���P��Ӧ�f�����J��+���"�� { 	���*$EM�*�:�V��Žt<qa��P��a�5����̛@�*��:&�_X��+�2���R,P�?8���gY*T���x�Z�yb�É�i!����ǀ�q�>�0#V����§����4��˟I㤃�O�oPP�TϽ�ݜ}I�bOP��!_x�3��i"��Rp�04�2b|�a�
���:���W��a��R(~���������y/S���j=����1�W\�{�q�΃G"o&�;�b6�qb��ɉe^��Y����#����?P��i�,�2PwN���"}�,,Z�n����n���9;��������ĥӛ�s��>�gVT���_F�rn$/�<�(RS� ���+#T���� {���m�]��9�`C���
��Dg�~OSHo�ru�0*>��t�!�bC���*��<LNϷ�i���;��q �d��i�
��ޤ�6���1�>Ld����y�/^aq�rW���w����{��~B����1�zɈ)g�3�l���OwI�%OX~��8�����N��\@į�
��i"�%z��ﷸ,��r��W���񁹼�� `xD8�:���0�˷37G��O��S�+��4��Y�=O�6���%v~��)6�f��c�Xc�*{���6��C�:���?%vw2~Ir���l��>Cn03/Rs�ɴ�����������~3�ݲ��ػ�7�������&G�.- �0��v��>7�M<`W��|���H=��;��q%a�,1�'����ߩ������}�8�"����{��m4��pם�U�<�?o_�R���G뤜B��+���m�"�u�l
ʇ7f�Y=L������gY��i<��������]$��������*J�>Oɞ|G���{ �����c23�0I?,Y��N��Ax���i�
�����%eg^�ǐ��u1���f�ߺ'T*M�`/S����e�OS������xɤR�����~x�����=�  k+��Y8���퓯4Y`�_/�����Xx��g>ÏS��'��[����y��PH)�+7�aLZβ��@�P<�4�
�I�Wc����<fȑ� �`R�q0~3�h����g�y�|t�d��j�_o�Nf`u
�̙��}�&�R,P�o�>��Af�8��y�|�Ă����|�&�o�d4�zʇ3�i��H>��c� �*ǹ�h�򿡑G˯�y��<���=t�L��xP�A0�75E�jE�ֺ?{��O2b!��0�ΐ�kI��CS�o��PR){M0�ۦeL��MdpO��'�c�=��-�ܪs��y�2��>���l��tzb��L{�\��Ș��8�g��i���Ru97M$��Lw��$����*�'���Jʟ?$��͠x����>�&�bJ�C_w �&2b;;�~��q�����L����3�öv� hv����iҦ:���ͬaZ\�uܷ�X�^��o�Jp	փ�(��b+jK^�,GV�9;3b����c�k�i���1̀|����C�3���SK���~���}[�+�kW5���'���~�� ��QY���=d����=Pc�I�f�*䩣�Ԟ�}`Vn�?�=Lv����
E��y�1�a�c6{CmM$�z��&?3<���f�����W�`m�o'k�s��/b��:ý��f~�� ���8��+&3G�f���ǓZ����R��f�j<g����w��?$�_P<��'�V~d̺w��h))/�>C�٤�Lz� �z�k;��ͪ���Y��G�6����`x���i�K�I] ~q7߰�6��P8{���I�ACI]ϳ -I�1�צ�P�Av�������w��N!wg�LNRu4����r{I��B���=o����p�q�l'���0��
����&���}a����p�����x'��x��w�taZ��?8ϵd�bJ�<;��~LH.�7�a�|C�̇�m�
��z�}���9��ߟs��������8钲�����~J�SϮ�Y�LIP��
��>d�}�I>g\gP��i�d�O~��2c��N^�x�8��1��'��m"��ڗ���|o� JS�w���M�~��M$�|�r��ě<���T�7��`i���?S�:��*T6Ohu4�
�I���H/̜�s���槽�tx¼gY+���=.\L��2%����-�ʧ�� ��'Ǚ���AH���	�.$|���'��H�S0+�S���lt�����>J���7=���Y�u�ACO�Ă�'��]�O��@��Q�Ϫ.��7A}���Gs]��=��ԋ'����M!SRrk6��Va^�5�bN!XxkXW�Af�T>a�X�f2bC�Ϭ��ɧ�
Φ�^��Y>e|d��4��}��1�>�|>�2VUV�1�xg�*�̳I�m ���_��6�O�c�{���C\a^�u�J�κ=ߺ'=J��Zɧ��&$�Ӊ����S):θ�S�X,���=��çJOO]%:�m}�v)V=��N��O\z��}�4���c�x~�nJ��}C�1���0��yd���Axw�Rz����I��PS����k�<�3��@�S���z�`�������/s��O�~��f�^t��Y�*�[�^�JA
8U�Snf]������S��뙌��*S�+}��y�^������%���f/NĻy'�v;���O��&iEu�*Ӝ�'ww��ޒ�R��ڼ`J�[�<��aO뮲YⳘд���u�g@�I3i�V��W�%�G��� [��P彉!o�]8";[�%$���茉ݻ �����pv�VSR�w{�i)P����c����=H���P'(a��͘�q�՚ӄ���G`��hTّ���\�y��R��N 8�#|]�{K\��&�e���HC,.O9�>C9W�]\�7�}�^��릒l̰���1zQ��@jd���/��N�4���� �+Q��qd[Ǘ��T�C5�*�j�ή�	�FX,Q�ƙ鉡����]WY|��L�z8�X�6sk��9�q�O�Тv�币��/�<���y������a���7���|����wï�S��+Х܍ˣ@�sYj��I��Y�sH*����<!�����s����5}�^��;�%�u1���Ry��b����Wmwx /'LY�Lm�m-�s�:�k���i�(�D���2iV]���צ�oˇ}����+����J�K�U�IVi�f�;`U�IMɲ�����ړT�t=��Z�vS�,33Y1o+�湊y��f@/���#OH�: W�l�Ҳ�
���o.N�)	"�Xk+v+QV<5�\�<��;Qz-K��A����Mq��`j��i��؏�9�K���{�O�����t��(P�x�ҺT�ǭt�.d�z�+��!-)Ӛ!�8��p��E@XR}��	[���ص�4��Um�qp���7ŵ�����zqE���ᶜ{
_[QAL|p V�@5O�d�J�N�\M�E��-�-h�dF�%�<�Cs��:�խ��cM�
E���7�Ͷ+���&\���i����7:���ܹ��X���:�6íE!X,(g�n��p�H���
�8�5B�Q�X�e�q������D���Q�2�	��MmP�R�Є��=Aǡ� �M�BE. ���n�r�V��/d_E��C[���5Bg\3�4�[�'��9�*C�:�K>K�p��Tg�� �K��ê<��c5���@g�!)(z˚8.ˡΐ���
G���j�$��L�ᴋ��WE��t�.B�u�O��λ�Cu��1��VT%�]������
�j/>}Q�F�@G��K���.!��Mx"7I�:.S�T�ZL���E�u��P`�l�1\%�w�#�*|zL����^����\�MѤc�������B��@\;ɫ����Ϛ�+���L��Ү#����V���-!ڝi���y�k�� 1��E���X,cF("
�Z���D�U*QDyeb1�!UX�� �QEX�b(�1H"�cPr�TFF"�1H
,Qb0b1`�b1�Q*�V"
���Ub"�*�b�[Q���1Pf5"����QDTV*"�TE���D�+ �B���

��UYmEUT��X,FF*,X��ܰ�����aF
�UV+"��*���Ub+�c"�[i@b��*�$"*��(�TADU ��Q����R$X�DUH���,W-�*�TQF"*1�F�UAb� �QPAUV+�Tb�AR1`��R��Ur�"�F#EF"EDUP��UE�DT���`��*�E`�E�1V"�EUTDR�V*
�mAVT(�b��@TUQ"2"�AED*����b�`�1��U��	mUQ�F��Dr�[*��UE(�1E"�UE��R"���,G�c���dQEUPb�(����y���:��]~7��z	ږ�*��Hm�2����x��$>OsiR�}"L����hv��E%41ov֌�Z�l��������r9���]1�n���xDdd lz�X4C�J�8ɉ�������z����q%B���kz+�AH��4�츐YΖLJ��]$�?}��8������Ak���{��o�4�;�Ρ�V5L��Y�3I<M�$�:�����H/^����P�{��ğ����r}�N T��ɹ�7�> bM!S��1^�*������=d���3������˱�;�j��n���� �`�[��pX��잡�(|��`�PXzԜOǅ4�Yԕ]��|�6�_�ȇ��}Co=���O�\C�}��ƲVT���ě@�T)���><���-$�޻������>b�B�!#��u���ށH���q���I�c%a�gS��<k�'=��u
���1祁�)����MjAgY��C_Y6��`_n?0I��c�������d�%��Ǝ/�O�c�0�r�+��G߿}���6�!��I�+�+4f`i
�^���}�8�eH�b|�I_ɶL�y�u4�`_�Ӈ�M��
�ɸv�{���(hK��W�臵1��*w����N��c>b�<��Y�%J����>3�N����i��Aj�exʆ%`c_�`e��=f�̡��A~I��5*'�c��i��|ԋ�I��Yn�y[�Q�W�	�ۮn8����a�%g�|~�O bO�^�0Ӗ�Y���H��q�}�Cl�%C���]H/����1ݓ�����z�XcR~?Y��Ag�7w�1��`xD8����C:��Wģۜ�����?%a���ܤ��'S\M��4�����=�M�I�%NOl4�>3�Ç{�7�$P^'�?	��<a�3�u�L�%g�w!R����ǆ��p<`	��W����}�6��B���������/�c#�L=�_ړR�|�7I�,6�I9��^�I��pt�^�-OR�P�
�?0��m�!����f�h%}B����m
�]>��Oq�T��s_���s\��c�1%'v}�6��P�%��zo�m
�Y5���PSHQ���JβT�=|M+q�_���?'S��6{COYP�+6����`�
�����s�j���K�.fī�w~�����r��+��gH��]b��ؖv�:�@'ȳ�qD�Ǝ����	�T�vw7�{��ҭ�;��R���ꂌ���5���m=8	��j{�vh��ax�:��(��
�1NewU~� x{�.�3����	�x�_Y��i'P�M�y�O�1gZ���֠xԞ!S��u�hJ���>�@ĝO9M0�
�l�*E>d�ǩ�~�+4�P�lO�_H� B�����|��5�R�¸7Ȟ��VN2��́�~eC��a�z�Ag�w�iY�=L`zw���LLa�P����|d�bϵ�Cl��Z2i��$���Ɍ��u&3��D�}��9�؄�<���7ۻ_x$�<a�n�ퟙ+8�^Kd�*~d����d�I���;�8�z��,8_~��m~jA|���&=M!���i�����}��A sY�C����~�MC̠ο�=L����QQ��1���������1&ЩS��~��YR,�0�b$���s]�T�C��xo��I��=��L����̩���I��`i�dB��YF����i�o��7��>�v���y���Z����C�x�H-g.�}eOP����l���9�q*Az�������c�XcXz�?2��>�L
Ԟ!w���M u+'�E� ��������7��/�k���Ysw���[AH��~��l������)
�CXu���~q����T�T?3�μՆ�'��1�y�{���N�0��T���{`���+g�o�=՟/�o7��5~6�`cX|_p�1�:I��|a�J��Τ�لPĊ���~ԕ"�Fy����J�0� z�?2x����@�N�_�ȇ���AI�&2=� ����������*V0�RL�V�Q�/�\{�����@<dR����|��$I5�1�i|�\�Zγ�16k���T�%~C̰Ri
����q�
G��]!�J�N�&�:���~7��w�_���$�;9t�̛���ϲi"�'�\C>��l�a����Aj��5ğ&�\�MeC�X~.d�bA�gP�?d�%H?���� l�zI贔�c��jX�9/����E�!�^0����{�4�tɈ�a�
��3������+���wH)8�s�
��]�ܞ!�sT�t��ma�Փ��{���
��^w�wߪt�W�5�TM4���en��u�[���lH�k��I<�@z��d�';�%	Bq��u��84�Q�ً�2����ֽ��(���Z��ݙڀ�X<�`�y�� [��g@��5χ9O5��y,��GF�Z&��4��U�A�������N��Of���(�� ~������1��,1���ct�����g�+��ֳ�hi�f?$�;gɦJ���&��aĜB�P]�ｻ?2x��g��g���%f��g����w��כ����U|��L�{�.�x	I��f�ԟ���A�%x�^5������d�O����"�4Z~f$�6~��� �P�8����ϐ�}p%@�+�־�Ǧ�������G��{/ވ�`{��A�C����a�5RWs����'>J���o�
��7����� x8��b��\O+:�R��4��AjO�b�É��C�߯�����W��mm_1��0�� (�Ͻ�p�Vm9����P7�~�gY�����3�HW�!��u`i�7�`i6�d���L>a���+��CL+
��~IPR(|�������9��n���>���y�ϥ}v���<q�q3�B�~�w�6��=C�Y8��PY�}��������p��J�:���o ��'��9�o]C��'��h.�V[��4�L�������o�����Ř��܊���&�j>�P6=�ey���4�HT�d�L|N�b
E�ì�u��OwI�%O�:�jc�����6�d���O;LH��^���}����.Y1�i �`oϵ�滟s�]y�����_S���H)���=eg��x�@ĨJ��p4�I�+=d��=a�S��04����N�����d�R��qOX��Cl�L�ԏ�����5����]��5����0@�G���`xD{�J�ְ�<x�Z�7a�����&�9��^���K���@��gP�1IXm�z��b'�߻��x( �{�#"�z#�}��'w��uw��4�������ܿ�˯��B����?�2}~ͤ��a^��uAH��,7۴��Cf����g��;`Vu�C��ya�4���.�hu�OY댜<�M2�������>懝�Y�f����^��uu���������}��1���߹��x��@�>8°��Ԙ��I�c%ezϵ�i*'����& ��j���g��M��H�O��v���'�	?k�]_�+" ?ٟ%�t�Y�Cú�X��Y�n\���nE����r��@���d���,f��b�ʰvGvF���qۉ3傓QѦ���f8�Ԟ���W� ��vd��{{ۜ 璗(貯�X��Wo���D���Y�\o��Vɤ��,�{_&<�΅\w���h�8�2�7aj�:4�Q�v����Y������bn�cm�LA8h�D%N�����ž�[]�����=<��o��ͺ?�Qq�l<��_�Vz�5�2�_�ÝÏ��At�ߩ����1 ��Pz�ga氋��gY��� T�4᧨V
LB��
�����Ƿ��u��^}��=���C�P��|Ɉ���_oX��`|�g�L��8O��m �C[�z>x�Y�N��m']:H-y�����>M&�yW��Pz�ǀ10<#c~E��[�ױ[w�g�|��{4�Y�%g�Y1�OY�x�𡤂�����,�%`|�^�x��o�����vLa�
��$�+'�}�~��Sfw��^$br�ChT:�풄��u_���O�ٸ�᳣����Q�#2��\{���I����&�q�$�7�Y�sV�M3S�5�z��:Ɍ��d��׬8g��t�HE�þ��3��o����t���Ld���IY��Nw~�|g���S�Ox��=��3��?%v����H/�T1�R��_��54�^���L~f n�&>�D����߇Ys70�qkʰ�����絔~ l(�
&=����f�Ӡ�*��_��K�
�vW�u�a)�Y��%��m�%��.U�W�[:N�j�z�qQ�˸���$�":Hgv��ۊ�Y9&�o�X��ވ\9%w�Mwf�`z�1K��D�o���]�s��R.������N�n�m����Yz�zp�z�B��eچ���)���?ܽǯ��/b���`�����&��w,m�7Gj��E�.�>���Hx<�0��E�u3��c�#���RX(,a�����)��VY�}ah�	��[��U,����7Qej�}k)e���v���g;X�z-
у	�b��z6����{���u�w`���AY�~�ŽJGl�BFip��8MB���Eͧ(���޻�	���-���ި���["�j@��=�$�|����;O��ʯ�xZ��pb=�ן�%�l�N�gJ����Pf���Ge)�2&:�\�B�]�O��|_����Z�[�P]�7�]=���À���*B��S%��X��ċ��	]1�]���~�;]�8��Gm���Tn���k]DgY�Q��̍�R��b96��c����r��Y뻍M��<�߲�l���ӁB����F�.Ɉ���fr{��~��!_�2���E��}z�T��!@�5�c��2�!9D��X��4��]O��YӶ�f����0�5^�\_��-�!��xX��;�Q�*�vS�l�=���-������훰�Q��0�b�x0���e�f
UD�\����bcmpW�}l�:�"����˶��Ȏ�BX�E3�&,�b*UȘ�-|l���d]Ʌr�d\�9��iK�ٮ��˥!y),D�r�Vf��n�Uv2{f�c3T,◛&�i'���/f�s�t+OU���\�d*:��L����²G:v������RG��7����պ4{ayn!/���Ν:.�L;*au��v��%��ŧ[n7ض�5�q��Y팷�9�� ��R�7��rG�c�;�;�W�v�g��DR���a��֠�ThkfiE[*�LV�!5�W�),�{#rrM��M{K�=M�M�ZS�m�W�Q�>���F�l\�&A��>ʹ�0�rѯ:��no �1׷P#P���Ձ���E<�c9n^��Y
慯$��������Z�u(�ɾ��<����:��d�@��O{_+֧�;�_*�++�J3�VԮ�e��P�u>}�WAi���)ul�>iүq���y<�D.F�ro&GZ��fm&a^^��2Tj{�){ۿ�0��<�T�m�� �w��=��Zr9�=X�5ջ�\��)*�>ӗݻq��wj�gZ�۞��Z"����+�겂��ˢt!<����ܐrPq�~�ޔ����=��1���0�N���
�#��RҢ���SB9k�}���R��"�N�ν�f�:XO�W%����)6N����\Z]�+Fe��xK��v>���x+���f:/w��eZ?�n��ٹ�*Ud���˰��;Q����H�^vkT(��Ѣ�p�Ժ7���`�fe�>��d��������+�����¤�O:���������ug�����YS@%��$r��������ԳLv���՞�6y��7&/�����n�EȯO��u{Q*����S�H��(��ԣ-{(�[xP��*�k��C ��L���v����f���ࢥl+=���d�a;��t���5�A�7r��Z1]�Z׎�2��1�\��ڸÉ��J����2�t�]-�OE�W �K���ۙ��{�@���K��X�Gq	��o]b�z��kB���η��{Gp�ٖ�F֣�u��Xa��-�T}\ޛr!�Ѭ��:��9�d��r�g���MY>�G�6˩�@�|�.4��؆&��o ��d�Oj��w��~���ch,�[l�R��x��c�v\d�6��ި�4�x��j�K�k'ܵMu_V��duJaR6��V�Ñ��t�k��F�wJ�m5cpj���H�Qv��!q�1�b�o!��ʾ�,�*�PSw��iy�s.�&�0�wb��d�v	�곖����h�k��V����^w�z��zi�P0�[$b���+wWo}�����꜋s���֛3�qM����w9wdP�P�ڮ�WG����P���jyï���و��A�Ȏ�e�\���D�W~N��w���TOؒzډ+FT��Η5�h*���C��KlS�\���9�hJ��s�\�)�X����oVS��#�	��j9u]v�3yDa��:n��N��6l�7�B6��K*SEM~j�G*t�s��9\��ǁ�-�J&r7Ƴ��9ۘ��j�'���E7s@T�:���\���7DNv�Fyr1Vz²�2;N��0	��r&���y+�WUHYpRxwf�z�����(	��&�s	ؕ~��q������xU���a�[���u#�o ܳ��Ys�����2������6��sg]��snm���WrCO�gu؂�5��ߍ�K�E��+��+��aeb�\�H�t�*y1{ ���xȋb��~�"p>Lb��N��q����>ց��ȭ�)�C6gb[W���,p�Qv�ֵ���+ֽ���ݹ�3X�:n��*7O�*ii�&�U��Y�����]��Q���Q�#'.w�����!��g��}��7�E���hl�5�O�dz\U�ߍ��� �q��xY�x��ʍ.��J�]�ctK,���E�oM՝�� 87���V����;�ⵤg+�X�Vp�Z��۫�z�l��6���[or �x�����=��淑}���1;Q{���:h�3���C�z���{K��7���n�g1v����w��lJ��+�Ր�p�D{��)S}�u�+��.��7�&�lc;��=�¤m+�eL��-* ��坭t{�si����ǥ�Sq�o;��+:�Rj\�R��ꌨV'����#�y�K��rGJƝT�[����_=�Y�G��J��q�5�3�:��Fn�.|V�I�Y�.�Ѽ���CC��a�Jh6aկ%���
6�畷]ͧ�w�Br�c*Xo��N��Q��������x�½�*P��xZ;{�Ʋ,|45b��B��lz���cV�СAҝ�7[��Ƚ?D���E�ۉ��kb����1؎����9ۥe�x���	9��gVp�t��U���).��)VX;��V0Ab��I�K�f�g*��2'�Tb�t������[Q���R#�I��ά�3�ٸ}�0+:���UjnyFӞq���U�j��-������H�'��k���2�����+#�+x�n�3Y�l!7�
Qv�'�9� ���F��b���[�A��f�R��w�ղN�;F`��&��B*C[0|������2]Gfd��nq����ިhg^�O�7"Nbt(��V]��ך���g���.w+��QKV��[�E��
����Z�K}�v�]���Y����u7=՚�s�2��D~���,��no������B�t�E�3�Ъ��:Vj1����>���e�!W��
��Z��,��&kj������^�|s�/+3S��4{#��|�2���h�R��Ur�o-X���\څ}��x�uPy�8ڝ�N�x�!)��3Y^��R ��N�8u�}��̓+4����UҲ�֒��y��������w�N�NOh�LPݮU ��.V��:\��f�j`�\�*Ū[���&��s��w8Ћ
K���u��Tu�s39����a��3��Y�m��t�o{����\��{u^$-fXp>��]zf��A�ĚU�]<�r��k~��MyL��c/�κ�; ��;0HN�TNG|�O+;��Pe��GYa��ޔ��ΰ{Q��ⷵ�:r5��:J��\���i+x<�jC(��m�ȳiUҝս�{��>#�s���8��L_iX젂YY�P4�I���ϳt�2�&PS��k�-�@��u��C��%�9��T��йV|%o����������vK���Oz�;t��2��Y���Xf�!^�,>�n ^�A#��=��m�4��%o�����x�@o���ga}a-��An�]S2(r�-j�W#h�9a�%�{�Ѝ欃�T!o�d���F���'@':���P�WJ�	4<��ö��� ���t��"�9��,���)����y���]MfA@�p�p�l��uu��6����X��T+���4�]��tw�GGUgRƹ�N��Ev5��:x�T@��f��{{�>�w�ɚ�*t[&p�E�ԛ�������[7�5��)�|�r�V�s5�/K@_o�s�;�E�\\7^`���Ho�bv�Y-�����H��E�[G&3rC>x��_S���:�=i+�7_r��F���4G,�6��$�o^v<Ӷ��+��Y��f�+�f�F�V�-��
$��� `�^���EO/��kV��
��� �7q'���BE}�l]j�b�g�*Β�D��mb�Sv1�g�+���sY�7ZL��M2{4cw��6~%L�e(��i��i/-�0v���r()��1�G!�-�V���
,�:���S����Ea��� �U.���̜�r�L7)����ܛ� Gj �N��`��2�Ǖ�U�)N��GïT����4:�x�J�ܒ*�*	Z�r}�Q��z�ڜH���43y�]�ɑ�C�X��ӂ����pɍ��BiɄ�aqh�:Ac�kْ'T��9�K��_:q��zVP�9�(�򪻄0�X ΍�ϓ�ܷF�z�țU��-���.]x޽ y>��auW�r���s}&=#|]խ�fi�3�@��H�Ҡ���W$�9��'7�"�QT��)�X�a�Z��3�.Z=}
����kP��x����IZㅱ�Q]P�+�[f��k_�����/T�X��"(5�EQ���X�DX�(�EEb����UYiDeh��W�Ub*��"�*(��DPTUX*�1De�R�b*F �Qd�� �q�EQV"�e*
,����
�EQU�PT1PEQڵmEE��Q�
�QPPT`�a`ڪ"(��QTE��X�-aX)-�*(1UbV����EETc"�"�DU�Ԣ1b�b�k���DF1�(� �������Tb1Qb��(���J��EEX�H�QUUQE�*"
�"
�UEbE���E"��L�"�0E#�*�,+D��#�֦!TQQ��b���Z1`���br�TTV(��QQ�
,Q�X�PPb�-X�*��R#b������V��2����y�(f�>���vE����o�h�f5��X�1�N�)��#�«�oX���ӴEy9����zP�����ْ��7��GN99����5�*׻j��I���gmvl�p�ߏ�
��uWW|����9��˱G���R�jE�n߳���lu�τvJY�:��u��j�j��up2،AS<n� y:7	u�"=��5�b�a����ٵ��ꬴ$�Jx�b6�����D;"-lЎZ�p;������v8����qf�9�/�Q����T�J���r;k,r{A�z���o=v��mQ�~�FQ��-��K���\�s�{Qi8�Ä�<s�*h�����Az���Jϒ�{W��Nī݈z��/zd�"�{U.yq^}�"��^m&��Շ�aok��"���|�3"����v3�K��O�l�D����J�̿IY�¸�O:�P�B���~��F��oB �����Ɨa��m���h}���BW�^y0@P�����ŕ�X�ڶ«�"���o٦�f̽���>+�pbs'M��Į�� Q��ۛ���f&��O��/���.7��_�����%qh�F^WWd�qr+e��8����Շ��	��bI�N/y]Z]J��Q����%�Sg�c�[{�њSV�#i�o9�w3VV��c�6���r�V�Z��9��T��Sҵ>�<�"���n�f,�)Ѝ\�/��YL�sv�Qr��i���G+s\��m��h|B����gX�k���P�Jrzu�%��y}=FT�c�?fT��f��O�f�+�{�����vf�[rO=/vg�h�^5s٣ӝ�ݍ2z���!w�z�1��������}ٵ���Qֲ��Ҳ�k��_*��N���vby�s5�77TtVͦꝩ��f1��X�r�t��h*x�b����O3�������7�&����^g*�F����/@n��lץg�>��?ye/��.����h�����{�}+v��MC۹.��l��o�VH�^8��,�c*<�{����y´�4�g0&ڨ���E7sEQA��%�e�~}�ygV��O���N&���nF(д�ͼV���>�38�N]ܚ�,�7iA��̵kzLM�\�6j&\h��%hf���Fyx��/�,$';X�nP}��uЫ�� U����p��Cc�nq6�*�pprQVb���h)��U�^��齘���b:�4�����:��s��^�F��
�bݚ������(����iQ<f��*���#��E��m<���������YC�5�>�=^�MͲކ}T�Tؙ�wM�w�mk��W5!��΀s\�{��w��c�
Ⱦ�T���b.�-���U��6J֍��}q@��h�]*��F���q9��0�ƾ��~�.�Z���u��Y�����y�88Uܴ�}��pw2�Ƕ����,��]�<y��WsQ%������;�A[��4�] ��t�1�9�v �js���A�^V��nC}�IobU�#�g\�c(V�U�ҋ����yA��3������x�/�<^ئz��u�O�P<��.X���w��6r��=]��p�9�Es޽~x��d����Ctq�K���Ԕҫ�մv˭B�5�6<��y�ݞm_o����"��q*g9�>ޟa�}�45\�����0��E��ԓ�}���jc�i-�Y_NtGO#^��,Y��h�cR25̢� 8q��ٷ�-8���C��[��5^�p���,ЬA\��4/�®�
 u�˽��}���Z�����{>�UV������k��:�PMK�����Qt"�^�Pג��ޔ���d��E)?)^l�K�{��62,X0$|��U�R�5�;OU�öl8yb���P��s:��z�����R�����g�̶��Q"��L �]ԴvFN�M\���r쬴����;�q�ob�F��s�ˑCJ�R9hv#U3��(
νu8{I��r��+'}Ϧ���t!��*a�J���+�ӓ;���ߓ���r�]�rOg�n�ƿw^�����P>j܊��K=or����
'Z����ʹ��=z&����#za���Kj�ؖ����^�N?o&`�`ym�;=�WgZ|��gm�ys�E�:a,-է[^j��g<��=�'���ޜޭ��.RwQ��.���Bx�^�]�oos�|���a�8]��<�2�Q�b�Oy��<a���f�b,w�����x�}ן���`��k��;����Ǆ[ܔ���I]��<�	Y�B�^.��e�t��u��:\L�ux��t&�!.�g [�NlYqRg�<}��Ul�6�r����j^����߀�WL��d��Օ�+Ǩe��ϫ�~;���H�&�Χ���q�����ݴb�j8�V�Rђ�U����\v�9:���jd�#���~�Nk�Rο7����M�闞���G�����=�=#�ns����p�P��6�w�'�ԱD*�W��a��=D�u4pp{�LZ��{X��M�"F_��b6�$�KbM�=vәwm&�,Y�[� �k=8��>z(�٪�9����P{�z�:r�s+�����~AW.�P<����'����ُ_(�n��'�e��-��+�Y,��C�F+�#�;�}Gu-aW��2k���9qW�;�_nt/������d5�d��,
��,nAj���ǚ�7t�������@�몵�Wu�n8����(�<S�νgb��M�N��V�d���;�\�nD����S��Q07B �o�]�s��|6�3�t���1�T<36mޕ+9x�Ą
��I���/�=5��ӧu:�j�|���>��7�������r������{x��;gq�q�v+�BD�'���|T�8�[���zl%ifo=��e*���%\��
�݊�� ������bX�U�0���=xhc�kV����b�EO�Q�md�dvq�ݽ�n竖�52�l7S;LN]��x�e,�I��@t�+��~�ԾF�g����N(uK_u�hޱ�T�L��|���g�w1`�(bq$b4�V�-�j"wU텫m�c�w��mb�8�"�0�n����=Xr�!�"�D��ڰ�XotJ[�X�!�r�X�ϯM=Ⱥo#vً!N�k�8���y�t^�*���������;�r�<�'�x�2�v��=�D[=
)w��/��{3��ͭ9wF� ���R枩��eTO��]8gl���k���;�D�IM���~���R]���U����oDr>�iX�ؑ������hݜ��U-�"��{�uzg�KKE�N��#뜻�����E^�Z��T���}�L��֣�:yd�cv�٣�(D;�3���_u݅�M�7�5�Ρw�3����臱T뭳(�J���pEGi��K���Wi}�����H�u������9m`e���Oe�v�ػ,�]��zׅ��4�N�^��η�6�t���ޥC`�;)v�܎d��uw��ֳ�d�;�T1�{�^�M��ud�=U߸D^)�]����O��,-��Ok��szV�y�в��*��.kּ�����'8N�yGl�ƍa�6��-�{�fڡ�����M��EH�Y�nj�%��=�5!c�Hn��DW�����^�Y��ÓsҬ^2�=3g�*��=����ц]�a�4�-f�-?���+���:�NzLL�Z��NB���Rt���ו�q��7�%S[�bK�7�q�bc�p�Od���_b.������$�X�}0�𕡣���	��3~}37n��e��F�����T��*��7��oQ���F�˧<./��%P��6���]�����ֲ�f�Ó��t!څk�^�)ս�4���j��^[!9]�v�S���r^|���n��$��qGCW��ꂞ�= ��Vǥ�!{�x�Z�t��EBZZ����խWmu>_K���2��,T��F�m�͉�F����Ń+�!ZN����|�Σq�uځ�;<�>��r��Rq�$���k6s��h[Z��y[��>zM��
�)c'��\_��7��mp�h��~:�]z]b@�cgO7�:Go�>�5��N/8c�7'%}�	^K/�بT��--�����(�V��hvw��UL�۴��;��XȦ�:��W�5�&z� _)Nf���KfN�-�6����"q��̠��k��딚��ِ�6�˴])[���B}NiWx��O��9z�E)5JW6WR�����=�g�%�\��6��r��V(��;J1���uO{u緅�&�C��tnx�{%v���y
��{%eZ�貓'1P�}B��{@�Yʥ:�}�u�i���T�Et9��h��l؇٪������L�7���g�8��в����z,:�Qr#�N��;����-x�>��u�2�͎v�__Z"߇�I�~���są��W�M��x��7� d��ՙ"h���Zz���z؁wN�������' :|\V�v�]H~��n���͋�GnV5t��9�}O�2��Np�GǺr'O3��u
�A�P�K��z���ּK�-�U��弓�Y� �j����w*�n��"8=�,����ͦL�Fv�f�i�Y9�3��Y�z�":a�.a;��t�3�������㔂u�)����Q�~��%[�Ց8��S�E����6v�Qt���S���Քr��Ws2K2�u�eFc�d���^�Kw�ml���h�J4i�q��.�}��D�\�����b]GΟP�>�y�!]��g4i^ltg�ս������mo��7l#@S���-4u߂�;E��}�6����P��:�_�h-�]�����Esk����y嘲s�\u}Ԫi���N1�^=�j�Y�k�\�yh&{	���!R6���i{S��}ߗٸ~�QXc��}�
�iUz�f__*�5��uʤo0J��yt�M����~�3)m_��#���#eNl��`�@��u���*DB<��O�����,v'�@�6|�g=7�m�Y�˭U�L�ʙ�:�-wTv��hޑ�-if�t�5-��ڜ&>�ވ��R�Y��xv��})U��J�v�U���v�n�Z�啬�u�r�h�e��0Uj�qr�]^����:���X�Z���.�5P�T8�1j����\smp}�첺ސ��1E<��'[Gbts�J�����ʙ�FL+����}��_���y���b�V뫲ldZ�]QeΥ��$1����[�g(4@��Td⹅w��.9/^��d=�^��m8�����.F	຃�έ9�<��Y�Y�Ϫ����M*����{Ts��6�T�r+�1nh�A��%
��x�k��&��';�����l�Շ�.q7�9�y�oczɒꦚyxRյ�a��s5��u	��bf_��hbȓx���a�j��y���vK�6_f!�D�ݥPE��&g���<8���Ughbq$A��#	�Xa�H�륮Wn��:m=�)�����}wL�.wU�9���X�zeY�l��Z���(��7@�|x�����7��lŐ�Q��=�
����p�D��� �N怺�خ���u�mB�Z�Ыγ��-�G���q�{x�t�;��&;kt-<̍m"��d�}�v��}�"#ya����*��C����M�o:����� ojR��
E��;�1M���}�tp-Nh�+NV�8��[h#�Hva�᭳���`P�M:O�|�.��h�;�WL���DD����)����S��|5CS
Tr1vM9V'R]�UbY�S�@HL�x�v�s����˺���;�1�� �S6es�#��X޾Q\�y�n�Ŝܫav�����m�}Gy�8I�����{�)��ؒgD2K�a����莜o�FD���zlOy��f��BIe��η��;Y�x��sC@ÑM��̘G�ԽW�����dJ�kK�U��[��@pv�9���:b-�kEo[��Y̽��{�a}f�.��=�m��Iqn;_i�������(���e����j��gw%�H&��8�М��蛭�[��l��\]+��T5����w"⭌��uk��j#�h�5���v�e7-�x�D��Ѭ�=#ҳ*5W���ۊ�q�;u8�R�T;I��E�+n���!b��۾�\xN�VA�*�b���Z�[:��0ͳ�9]�z�!r]�36�t�!�wkfXM�|��êg|v�s�d�w�m�Ey������V��P�C;ri����T��5z�sk�Q���g�Gr��^U�P�D��1�,gQ��u�����z��E���R�m��W:7]Jț�����7�y�G\�V��A���3�i�]|Y�9f�ݰ�0�_L�`�+$��7�m��Ϳ��]�r�]l�0iFѹ��r04��!(m'|�s��1/�
�b��z�V�����ͮ��p����u�m<�ꄪ��h��r��.��!n���%�i�y+&�n㘀WAg�d��5�S�B�ڜ��廀�a�jnѰTN���h��n���D~�m�xPZ��own1�OMe��v�s�g�s�������	Ȼ�c��ڛ}[p�����9d��z�,���	
*8�f�g��P:�>d��1�D��u��H]�)t��"����E�c���	.�i�]��5���w�+b�|����-��Pާn�u�>+A��KN��ս発���-���Xyؓ���P����d<ޞD3�VŇ#��p��%G��hUҺ-�uo(�	�>�b[�l��v�YĦ`�ΘaQ��cq�\u�^S�C��N�ǫw���Ꭵ���v�۔l؊�j�c�ə��U5�l�!
&m��ӕr^m�S!��2���M�������U>2�}�Vau
���0-�بz�._�J@�Bѽ��z����fo$@9K�UK�̫wGE�qq��xe�ϵ�K���HR�M����c����At�ޖ%�G�ABh�klލj�v���{��}E���c�R������
\�J��E�6�:4�QK�p��EhXt�un� ��v0��+�����[$�-�C-U�t���8����ڇFin�M��	��/]�ζc6Ԭ��v�<�j�����J�X�dN/��\�.$Α�=��9"�N�L4,�Ȭ����Č����Հ�,Y)�6��D��������1"�F"���W���U9h�*�� ���0R��Ũ(�"�� �kAX��X�m̱`"Ec
��PdPU��V�e��*�����b�*Ȫ�[
��#Q��Qb0ATjQb1�Qm*1cEQ��AE-��b����*"�X(�EQ��E���""�[)mH�����EDb��"���EEP���ATX��«mTV+,V��V*��D���X����(�P`�DU���#R(���B�P����zGAp�e�W\4�1�:��]c)�*�#�������4���˳@_m'�Ru��l�-�뗰��o�l@W:[-�S�!��TL�隇9���b<.n�`"9��1S�ݺwT?6�KZ4un�WLR.����n��_}f�.���gEΊ9W3�Ȑ/��,�ʜ������+!+����Tdp�tn'���uж9P�Gu�٪߯�n����Uh�pu��X�U����G0ͪrVY��&y��}����h��7a5�m���L�}O5���y���5��Hh�E�);Ks���r^
�Z�lv�oS^n6y����!ܸp�J�2VY�U���r�kEn��7v��|WsG
��4�Kv�{~�1���:٥����;�������q���ĵ��uK�ί]=�s:���i�,b�+�A{Kϩ�����s=~����7�զ#A+�Fm�z�X�m�Ə�<�nƁMܶ/�gT��כ���}��G��T(A^��:#�z��1V�'�0+#\#�xrnNlf�'0=��FnF��r�a ��5��٠�41c��YaNN��0Z٫J��@��6l&�*u3���[��cf]X�XCE��\;2��'�]5�;�|�����oe��'"�W��%�J������Ѭ��E�nf����\�٘�.bx��2�H|�-�g�J�[��c��	mM�W0_\̟'����;�O��TI�՘�v0�-Oٹ�_��]0���v�c]H>��4�r"�'#�qz�>]��tn���a���u���l�����E����}��y��^,�r�9�:4й�\ݠ�8`��}����b�<�[��[���%�f���-�n�FʝF�WS��Y/1
�x�lշ|u+�w�1�9��U��߫�ۈܒ�گ�Yqq����N:�:��z�G���q��d�`L��yo"�>�5�~�֛���w��5�3S,�R��;}��c���w��Awy*�wo����6}�!�ٞ�/��Pg����u�X{�#B���L���g��n�,!�n�R��`Q�[9+����V��6��4���~���u.�=����LKG5�Ƀ/����G'��,'h\)=y9V�H��,�R���/-TLFU�FyŔ�|�J@�uMLgs����(�,���ʠOF}����Ke\�)��!n̻u�nuA�����]X����|���9�r����|�h9��c;���m��kh��[�2i��uX���k%��U�9S<�*ok��OuE5�Շ��k���i��s�R�{@�}T��cL���ߣl��I�-)	`���{yݽo�f�ֹ¨mEy��[� ��T�J��u�;��c`!�s' ־{��f�h��b���AO��'���ȯO�&J��Yz�3[��+l7�F{8Z��m*�(����Z�ߟ,�5�+�n�#t�3�������L���W��q���ݫ�
���K�Vlg��6T#`�#��E"���=x�fw� ;<���x��Y�Q�X��!���_.]@{"���6���:�ݲ��}��a�~��]K���K�^QཬR��Z�;�CͮI�=k�d;�n�/���8��Z�;��U�"p:�ڹZ���D�29��90[]�VPQ��i��=݃��٬a5�@���h��2Tiis�FI*W�\������S5c�I�i4�y�!���H7��۰���CnO��C{��b�W�Y�#ef�"�H@�*qT�
��zlM ��޳�/J݃]_ #/^���S-}9!�S�7�`7��du �!P�@���{0�y��I��JÜ�Z=�/��,���ɛv�rx�}Y�Z��T\#B�]��r|�m^�qc$�L�w�S��#�����bF��vl�ξ�u�b�o��ݭЭ�*�#
�fq�����L����8nOG���h�J��YN�����4�업�]�Pҁj�������<��s)����37�ϲ�eT�&+Q�,�\��Ad�'�y�&�{�=yu.�]�4������y	.mu	�ԟBX�u4TԽ^sb97J��·���zzE���y��Yf�r>[�-�F�'���h� ����d�w�Li����t��'�z�=;O'#�VF�dv��ʰۡΣc3"�,ܛ����M��5!͆���r�/��Ŏ���Dk���vh=��.�;n�#b�yB���06:�z'KɓPΑ��vz��Y�.h9��]�2�+a����gJp���r���dݼi���]e)�����C�q�+o����N�3E��]K��.L�h�'>�`�nsg�x�ֶڕ���k������r��EsӔw�>o:f��3�L�e������=�;���|5?U��+�qA�b�h��?h8��\̟�����Q�N�8��E��λ�]�Ѹ{BB-��)WgF�F��ư���͝49�����x\���Ux����~Uͼ�~��(�b�3�S����qM�fw����_�י{�wS�ˣ.QNǍmm�ţ�w�<��O5�A�Ɯ��Z����ՇW��ey�������Y3�ב�#UOY��
kf���{KY��.���r�*�6�J�{��&������ˎ�)�T�0���=�kr�璩�V�B��"g�Q|�盌�����=�sm��=�Vo]�ݷ����6��ԩ�xYP��ںB��*�Gl'��<��ŕۤW��L��:����O\�����C[J��U�������{(�kW��������*L�e�e�����r�)�mN64�m
����;�2�`�7�����V�k�����ĥ�z�=z9xF]8�umF��z��:�]��=���.vTr�ν���5�����h�Ѻ�O�UN��7���Z���*�D�~�9�94�{�%/Ͱֵx���9���C���V�υ��t�sB;n��e�f��ڙ�,��K�zso1+'-���bt�l%_Y�bĨ��)޵u�}���[RL�V-��x����GR�W��~�#-�� :��8\����hW67\��\�d
�0۽�˷rcX�$XЧ�Pn4Pj�ДP�)�̗xp{��D)©=�=XY[��1�lč���E+�9p
�Q�7/��a�[˽�3�,������q6�in�L"��V9��=S!�L�JT�E���X��P]n=x�ᨧr��9��6n���hn� ���iE�z^uf����҂��v'�s�X��XPf8�Ѧ��qsbзC8N�����%��k��2�=�\����9�p�ͬX�֏M�ur� �ʟ���E3�ͫ��&/�LoZ2��[��Q	O��nu�$�x�1����/�ns��31�y�ی�znC4j4�d�ީ)`�޼:����[��zu�$��̧Y�k��y\��:��M�&m�Y �8�9]#v��q�k��3�����f�ĮCؖ׆v����Uo��ox��f�'�������:F"}�y�V�͈��'����3ٰ�ym�W����l�ndܦ{��s���F$��wbh7��dN�=�ݗڍ��Iywtd�B�D� �o�=8�tŢ�m�+�\]龮�T�"g�����u��Ǘ3�����P+�꾉�{u�G8��hkO�o��u�����(��C����N��N�3���������4��b���l���F�-�w2�N4������[;V���T���q�^�n�.��]��(��m���(sq��<��!��ຼ�;7�_}��gGK�)��n���U�<�s	ߧ��CU*x>��N)GS����_���ڼ��|3>ډw�ݽ�y�$k�W0�)�E�:�W����Ř*�l�M{A�N�*[:P��/:*���л� ��t�$(���-��y2�����U��W�rT��s��Eeu�x#�^*��s�}hS�C�9���f�z/�U��:��2U�08�l?a(V�1�Ms�4�l�ei�R멹�Ζپ�O����z!5��ʨ�[����{2�^:�$�i��[�e�f.D����8��ku�K�mU��d]Po&x�<\�w1`�9@�qA��f�ː�gN�z�.ݷZ
�-�{����b6�:S���Q���!���U�4�9�f��T]-��T��[�k���`�q��+N��G<�8��;K��\m
��xg^��j���y֞f�nNJ�׺4��^�.؏ N=��<t�i��[G�T�W�%[(���˓6������%������.!0=��:3-�D{�_ݩ2f�{�Jn�� h��.���ͨ�@"��ǲ�b�x��;ڐ/�]˄��ڧ|y.��¬����i�d���|;4�D_ڬ����Ɲ�){3g���1��W�9�d�t���4�U�ʙ�c)
m����9�N��/��7.��<�B�-�[w��^���tfj�5e5��ȍ�p���x�f�&�&F^���}� �z�����t���8��*��m]H5�;{H,K+r>�aoum�f勺sט�]]}p!��t��Š��7l���7J�0u,���۫z��#�B�B���+I���WP���Q���|z��3)rr�7�2�qq�c@u�\�y��bW<�|�l]�O7��W�e3*h	z��r�!�E�9Iv%U��ێW5n��4C�"-����z-��01xGD�e�]�uɖ��ԅ��!�v����P�(;g݇�G4�P['�o�H��ȅ7A%Y���e�ǎ>4���W��g�(��k:���#�	~��[t[��{.�rG�9"x=�L�9˼ �f�,��۫}ceF��}�7���^0"�}�V����+�s3�}�gu߄mFe�ǣ�xc��K+V�H𻉻Ȯ��|���6t�o.�յ&����o8K���g3{bng�VU���Õ����҅{r�<�˺���`O#vl�_v�ݢ���Os]�8j)��$M�/k}��<�5S�+�Ϗ�#t��q��h�4�L�AB�ȵ��:���+v�^�=Nko�t�]������
��V��#��U����������xMe��^z�eL���K��o�d�>B�qBƞNv��B��Toz&l������lm,	R6�J���¥M�����;�Z���,���O��������ܰ�J�<Q
�)P�Q�%���8���K�P�KV�[5�*=_,�}�)<��weY~3�s�RG7p+6T�j��J��}~�y]�|+�{x�&[wʆ�J�r�ngJ�ͧ5�i�͛��Lu�|}U�9���h5�X�S*yl6�j!_5���Ō�U㣕H�}R5S(�sP�e�L��=������}����I��Q�}��L���<8�끪� ���n
yt��d���û�,�Gs��c�����36ð[w@J�"���<�sf�j��6���;�ɬ�J�rc�x۳_,�)��LsV愠��J�����]N�+�c�n��.�$�r��za�a�h�5�������E�f
��zj��}/d699��Z}��tv�d|��v���Z�`o�㒌ۧ ��d�ޏ�S���0h˙m�{nu��Ebj�t��W>"��6��89�\����KE�]�{L�NM�9�����dkl��wX��F���QYX���jUԺ�-yS�t�'j��9����ER�X�:���������e���.�QT��;�MqO�3��f�wr���Z�
H�u�4�Ŷ��n|�ɳ��S���v�kvoh�,�����
�Om�@w,�V��Wf�w1ڃ��c�s�em>m��xV ����I;ctc�b�������- �w�����=��9ԝ��8�n��#�\f���:���i=@�ݝI77*f�����4�m�ϰ���cK����x�w �A�k*[�Waݛf��8'[0݊�@%�5uM�Gr�s����qG!��n��wNv)��M�N@��&Q/"3M�Y����T�Ʌͨj�y�yDXk9�:3r�u1u��[�yt�!i[5���u�86��&��]�b��� ˤie�ɹQWpm�ݓs�'৶��)�]u��y)���&X��Ż~�
zO�ա-�Ǯ��qY7�IYhk�:��u�n�+�Y6U�*� �hӧ��tv��l�J֯R�BݻR��OAAp&���Y�IP�.�imw*�d���C�R���_Y|f��et�i�F�J��9K�J�k�5�\X�f�H_v�u�b}A��&j:�wRE�hu1�f��Zj�̱�=�
r�zO��O44P�ӓ�|Ju�j�W[K)x٦[�(��* �u�;q[H�Lh�|u�����V��i�,`��$�n&���m0�J�Cfu�N�ȥ�l4�~\����ˎ�ݶ��q/���NF��{H��Hv�v�G NC
d7��b����c���cyE�&<2��9�z���tG9ZFN)���L񳑼˭L�P�72᥼9T9G�>SI:�k�[���c�o_����E��ܜ3_U̩&�KM1:"ӔZ���7�v�
���c9�6=�ۗ��S��!v��Ӑ||@�0d�/=X&�	�7ɲ���mgdX��\�k�M���( �����y��OAY�X��'o�\i�%��cЙh��cq�
mD!�B�����ϙ��B���θ
o�P�nKyI�|j�/S�� �6eG^%ա�$NH	�O�j��N���v|�^xg7�<�;�bR*�b*�Ab�DUTAC�(�,X�D�+l��*A`�DQ`�"�*��*���Ȫ	P�� ��H�#UF,X("�Q��A�"*,UTX���EU*��PTQAU[j�ȌA�J�EA����*��A2$c�**��
�*Ŋ(�X���""/�TX�������""�����ĪcH��,�� *����,H(��"��X�,U`�(QPUE��VDc`�U"��DEb����@ >@BfnK�b�(w7�u���%�Vp���Vy�@8�Y��2�(ֶ�����<�
��!j����sz���v8h��.�=����T�A͝����-m�ȓ�e��Z�����Z<�i���� ;��0ߍ�\k�m�7��Κ�E�wo5&�+��kڴ����E�cr��qS�h]A�q������ވ�4�^8�s#��Y�˷z�\��lv]�S6|�#G#�b
d��xyfv>�{�պ�p>����o�~�6���{��T��8o=�]��V�^1�C�g{y�\�5�~O$�=(\?l���{S��&{����L����J�I݌Y�w���Wc/;�tSZ����h����c;@K���;�3B��b�Q�O�	7���R;Q7՜�ɋ�S�� 5B�ﶝ]^�[�{N��>u<ݚ���؉Ŝ��w�c�sǀ�"���\����>���}��Þ��rV>�ׄ�[������uy��˕.���IN*�.����%���f�����(�U�g\���;\=��Y���VwS���\��KZ\�R#w��<�|�k��=/��3��<��+���E�n�:ox����u�9;�����`�X�V��1j�YS�d�{)����Su8EM�Y�a��b�dd㌢`�U�d�������f���=B98��6�h�ّb�<շN;�N�,��+���?J�4����S�n��b��5NAA�N��d����Z��6�2W9��g���5ac\5�&���:\�oua]�kL�w�X��m!9�*�b���F�*�L3ҟ)�6z�*ɽ{6R�B��k�����ܙF�g�n�w1`�(N)�:��ˇK��x�mPzx��-�=��a����y����
�f�Iۛ�)����OD�&X���N��]�u��N��t��\�7љa��ǃ�[��1�:!ó��xŽ��u�B}��y�XO3m�GR̅����f�J���]��U�V�I�z#Y�V���˓6�9�cB���E�)WT��Yh������<T��F�5!�3)�[/[���JU��>���Wǰ���VQ�Ω���.���j�]�\�nY�S�53�o;Rɘ��W[ܭ2Wa����[w�;��'���v�Tv����Urt�:��y��\�Yoy���V��t���W�����hzx�+�Lݚ�[�IօPy���w���2�$�	ܺ��H��z�LЈ}�&O,�/�Tc�� ��Ÿ�7��(�k83M؎�U�Yt��<����5qpv˹�o/�n��c����|��r�T�K��w� %Y<���[�Z
M�&��?i|�>��CZ����S�	>�`cLŴa5撥w,5��5z���t��Mjȝ����,Cˡc���"�W�rq����贸*�T���,p51g`�q^X�P��x{~Be\�z��b��`<�4��qO986�.�EO*N��2]]ڶƫ>�}�>�+����v)��E�u*]�v�F�u=���L�S9�`�f��"VLrW������������}���G�z�ų��>}s2COhL�;v]�d�u�W�LR
��$��J⟍�W��=���%-�Ҹ��wt��ʾ�ʗ�5�7 &��ߧK ��b��w�-iͭuײˍ5�o}Ǟ싘ǻ�PF6�u�t�>����3r.'u�v��W����Y��h_�M��C筮��y�EW�r�v��B��B���F�b}�:(�,�l��]y�[Rn��2w]�s[�ˣt�bx+c��P�(e?l���VW�,�!����1&�{͌�Y]��b�s�f�����l=�(j�4z��J�q�".1D-�e�f���p]X���l�mw��5SȰ~��Q�uhoW�Y�ÕQ6lҶL̽�ʵ^M�.ܾ!X]\mS���g�_�vߜ$�On��	s��{i{��).[c�:���S��R�;�2�WFѓ�� ��ټ���-�n�vt@}HF�/��M.�g��ᜐ�Yʣ��ts���	ŷ���Ӷm�yb�뫦���F�wSyV�6S�s��f�q�x���qpٺ{��{안_���[�J���kZ��f�D��uӮ�K3�`�g=%K8��z�{9�U6!���ϩ�ֽ�;k�*��=6���os����S��8�9���вE^K}4��wm.��u	�vR��=G,������Ac^�7���J/�j/Mgz-k���(w�0c�s'��@;]���Z�b�y�WP�/a	��:��f�z�N��h�+��kF8js؉0ƱWX�������ƯQ����hu�W�٭L�_���O,R���\
��r|�ogE��]륛s�s�Na���Ԫr#���\<ܣ�:�L��㐲¦�������t��Y��Dj$��-����%zm�MZ��r��}���1�i��8/�4��W0�t�X!����ܞl�OH��wg�j���tԓ/���"H�:Z��D,,��gz�wvsj�2�v�f�;����i����bb�f�֞��>��Aӱ�N��/�Z�s}�m�:u�z��yM��)�3s���PB���[o�Fˬ��o����-�|�Z�ϮO�\co�gxT:�:��Y���nË���øHh�ͬCo:�x��=^f��W'�+�:w82<&�O��]y6V�R�x=�=
m��K���:�F�,'�E.��8���7"�k�':.{�q3׳s~�K��N�\���x��:m�kk�]���}�Y(�#}�$�e��j׊h�J�f]8�6��=��/X��Z]w]ǅ�we;�y��T���)d�0cy������jk��%��Z��[�=�gr�PΔ��Y��N���.o��ߋ�B�߶�ĝ߆,ŉ�+������������e�z{h�F�D���ο
Ɖ��$��G�����U)�,��9@�t�>��A�t�\u_tq��03�'(#�i�8�v��;r�c.x�t��䄩�������N���D�oZ|�H�.�]���68ӥ0�KA���Yظ��xJ��m��0V�l��W��Yҷ�vy�Z�jq^n��m��/]����ȣJw�3ɾ���!~�=9�Ns�u��Ɵ�h��`� �4/6݉�������O_di���J����>�����Ϻ@߇�z���^��<�S<�n����P��츠Ӹ�����ffX+�q812:�\r��ouL2��!�K�mg`d��fx�-Dn���X+V'�jL��<Go뽳��䊜Q��P�t �u���Ԅp�7�jM�^�.�����72�O�T�R!��[�;��ɡ�����NU�T�ݎ纡T1���ӐڳbU�)�����-U}����lH��7s��-bʄ�5�λ���č�V+����A+T�bos�KJ-���;ޗl�{.g���I>;����g(��s�H`�W������{��o�{��n\�n���m<BX�g�ݸ��4_�E;�=C�^�wچ�sɥ�f3�����x���g���k�7�����9��'���Ѯ�Kt��u^�ɛ�\fA��QO�ϔ]W1����	z��%t�Z0�C�ce�P�<�3�⫰{����Z��@gw�vJx�"��=�&z�/�`0����8rH�;��#IcU�O~߈�_w�ٹ]v�ZtP��` l5C��%Fs�
���X�O��K(�p"{��v"�@���M�F =�M��Y�m����u{3��Y� 6k(V��7yGX�Ш����{�E�1n��ܖgȚ�ܫQ,0lu%��<�̟!��K�%`�����d���_yfʲv��q�=a���Q�9���L���d�y�S��wi�_��ŵȊE�{@묣}F��3�ߋ���)���^�s���:�N��n�k|,���SE��꽆�8��r�5�,p�5JvL��Ģ�Vܨ��z�C()��������|{o�����45�*�ZZV�啕�6�q!���I��K�ya�} �_5��sL[�f��õ۲�h��&V�8�Z�r��{!w�!�;�e?����=�+���_\.e9�Y@�8+$�	lT�.�d_s�|i��9\�q�p#���8��Pw��[4!)5�*�
�ѮeA�C�OC�}ں3�vٌ�>	�D7�UdDS���>O]���s��\(�k����zl���Z�s�SZ~y��(�l[=J��P�Q.n>>���>Qf#C���'�P}6	�1��;����|���R�u�c�u�ٓb@�d;�eKj���C����YW��	 �.���+)*�oW#[�m��-�z++`u�aٗ��T�|��ʰ�	��w�}�����S"wB�@v^h�U�i7�[O:a�|��^?�w�)�N,a���=sQ�����[cgzwv݇ج���7���
Aڷ]!O����Å�l^�9$ڎZ�R텀{5xQ~n�O��^
іf�]z�#���HV&cT�ڂߙR�Ъ���e�J	Gj,l�u{6�\_�� �WC��꾱������J��d(Y&�!���e��	ʂf$�"I�$�c˸^_�����d��Z��x.!òN��jNg�u��l:{{��z�Q����nr�3�8�9yݭ�Yu�}���������n*��3�^�=���=�o�������!�t<�=/,���,O�[d#��b��q��g.ӣ�BOG�Ct�#����K�;�o�+���襼|O�VV�`?��Ĉ^�fGmU\�
7f�a��aT����vJ׾ɸ�Xp��0}�<M}��x����@:<�!�N���qWzSy����(���º����;޲4y2�W����D2�pY0[�#��b��ܼ��[�eڛ�|�5j p�F͒�6[�*\\D7n�J%��$��g���+�޶|7��}�߹�"�E�r����¡t��>�� 2�\c��NQg�@2�I��L����Z���g'��z��a�|/>��`��53����mj�� ����(�e��,G:s�A��|�eV�2&&�0ٰ	5؉��bK�^�r$��P��n�B��<��e�U���� ~�f�y��Vl�OF[Q���%z��vU
˳�4]}��Z���i��V��d�"�f�F(wB͐�RkA�;Vl��6H ��b�� 
�q�A�Լ�v�:���LL�.�O�� k��[�5���I�̂�q��(Ꮇi��Ī\���4��g)�]v���ח�D\׋2NL�$hl��|�h�p����oV�y��}��~�6��z��^��~�ds'�(�V�<���/֬��ҷ+Ŝ�*����d�DSa��4_��'����DF^�����7m�׉Ȫ<<p��&铺�b�죴]�l�lE�b�#uX����J������^L����}��[-��;x}:����yd��l�ҰL�3���RE���k��W*�Ύ��QxۀɲL��ۗ�g�cWƧ��'l�H��i}�c����0n���xkE=���.�Ư�5Vn���|ک�6!_��UʤU@^[����k"��n�<�jн��޾E��mp�W��8��<|,��w^K����� ���]�^V�Ws��w�=휚N~��R�z�>Ӟ#O�_����/l��,�n@�4��E	�V��YV㸳!�un��An�g�n�;���N�U�Ӷ���z�f�@�57�-2vwJ�`��/���;u�8o�P����G����<T9㍝^����LИ�����!�R���m�(�]�X)}�B�* ���ٺ��*^�W%FEk���=)�.̵3��jD#���������ζ�-ӌ��9�^o2!���kv+ЧQ�m����R���#g���+$�;3{L��:w"b�������5�� .V.�6������%�B|���J��V�^]�ح��Z��]��:�6(�Jr:h��ɺջ&-[x��ҧ4l�D����J�xE�"���0�����X�-	^��+��w��9��dJY����V����`��6swmi72�\��b�u�-�i�T+1���,vj�QmKxo2��&42�޾�n��:cT�p�u�{V&���4�/�3\��km�Ց�p�e[�	����cL7�����p[qk)�����x�I���o�c�����;{bU�D��G�jw�/���1[9��:�N� 0�pIr�Esȴ��u3z�oFX�8��n��<�I�9Eά����ɩ\W��/r�y��Ld����F�c�����v3*�ZO��}�T�K7����i�e�u�SU���6�:�G����c3˹��>u 7��|E�{'��{*͹�S�a�k��"�D������"N���k��
'�u�4<� �4�T��+p2LrmB���v؆�H}�]�f�iT��o`PU�u�l�C������{�iҎ�n⫆<�x0@��F�49&�c {���,I�.��H�{yg+.��E_c��r�h��tb�*�x�)��3Q���7P,�U��k������L؝v�)�;��ݾ��@v���u$b�Q�c��+X7zi�F̦��������+p���plז��XIm�`-�������,�l<���E�g<_m?�J�OQz��ԣ.
W��Ӧ���`R�fb�C�B��]Ki�얢�,�l�q�Di>��tI��ٴ�����[��|4��[Tu��!�WFu1����k9�Z8�b��gOm�pz��5V���G�vt]��䜝&�_Y-i��� ���(͌PV�Ztݍb��v������̪6�tc��ֱ�w�HC�Ț�n�YQ]ĵ�WbgNċ6�nR&CWP�֣���l,�оp���uoP�Φ�]l ���yE]�t�f�SJvɨ�Y�PRs��<7>�)J�{k ʗ�5H ��ں �C�]a4Ҙ���X˲5������ޠE�N��v����Q�Up0t�
��Y����6k"Wֻ�[�1t���.ZB���;��ԕ���9cj뫶��.;Ns\1�C�Y��=l>'��6���u֨H���	GGr���[:#��_$���f��t���*��^�l��%s\�tQ�#b��1�#;z-PKEj�	݇��E��+z�c�F�vf5�j&�C��y��4,��'bdKH�*3o)I/��[�DgM�8�o\��Z����J �L�A�2�3�Z�(���"��pv&%��t�4T|/Tr�K�ޟ��KKc3n\&�h�\C�Y��mWV�'bc���P�M����-],�R��0l��'X��gS�r���VJ�˖�
1�X�X�6*�Ċ��風��F#b�#cQQR"�QVEEQ��őT��Db�
��b(�����DEDDX��DTQV�r�)���1�2�*��QDX�(����1TR*
��F(+"�TDX��PB��*�`�Tb*5����DE����.f�#1Q""%ecAV"�P��1b*��&R�����J(����1F
�h��UVڭ�U�ª��EE-� մX�Rڢč��"-�С���=����3Y�Y����գ�b��X�V��ܡ2��gh֥M$S�Җ���m�"��M:����y�b�Ա�l��V��s�g]u'/m+ b?��q�P�f
{��tJ��8��A�Q��\���ozE������H�.�:+�&F�glL
�l���e�ᐨx?�|�0�s,P�Y�	�.��6[�cv�6���N*�"����)s��,ݚ\k�ݞ�S_o���� z�F?+�Ѯ6��0p�	wr���܏`�>/�h�ՇT�Y���&�o``�##E��h�ɨ��ͧ�!:G�dd�6ƈ#&���,%�9�������oX�� �j���Xr��j��nZF׳}� �r&�v�^YT�7�:�&���!�=�aC��FRM�@�����ͭR��gL.)��Vjz�v�^��&Yq�65��g̍�Q�al�8%�;����w�����#B��1+�]�+�<xخ�����@�xХU��}\���̤��G3ۏ*���89��p�|z3��3��
��_J�ٮ`�xo]cC�wnw
�G+.A"�?s���C`w������I���֭a���BS��5�	ǘ������`ݠéH^��A�y�t����^��(�*��G��������z��؝��76G�='w�j���yL[�wW��8�rʬ�2rx��2�D̦9���}��`��t�kd�Zs��u�l�'#+h٥���6�FYKv(�[ev�J��������J�}g|s/�+�g�u�Ƹʮ:���+��T*�~���a#����;TC`Q�R��nG��+���bټf2_kǂ׬����%72�Ӣ�E,o��\�l�/�� k5{�|e��5��_OSu���ezݬ��tɸq�k�9|��#W��T�z`����T[Ny���vkJ��y6��jr#9��ۗv]�6��U@�V��D��Q{����\ȣ}!tOxܺU��!�q�W',R�ܘ�S4��J��=�,l�ˡ: �N �]�=P��MB{�f�%&��`�^ɇ+e�v�6��N,^@��a�ʢ�*�"(2��4�:��b�;7<ǓIlm�E�V�#kk7��#�ڲ�/־�c#�g�����.F����� &~�>q�^�`"���״�J�KU��n�� ڐ��N��z��lɿH��;L�)mS�r���-7�'���N-Mw>�u$�������+4�Tn+f�1/�W��C�+��gʁ�l�U�X�u&�V�Ҏ�t<���T\v�z������y����mf��gt�yw���G.3��M8l]�y6�,W9�Ǯv"Y�D�Z����3�#.�v��J[��|���:�l�g����ʰ�pecǕ��fr|3M��n�.�C�am=V�A�2�}�J��N�n�m�<�W����xGx�:eߨo�ը���O�er�1���]� tWBlߒ�h:)Y
�t<]��]G}/���}E����1Q��cTE �QE�7S'��,V=���t��u���3Muy�N�zS������;ʰ��c�=�i�ň|�4���U�����
��S���Yj�iV*҈���4H� w��-�e��<~���jV�0i7f�e���u��;(�[7�ݏ��.ז��S�ȓ�f�CEL71�]}Iy1b����J{���#Vt��W�#�z�[��f���qNŨ�T��K�ϫ�z�?�k Y�@����
���\$+�Kl^Ɓ}ם���E��i򸍡f�G��Ez�0�x��}�΀&��N�*�w���gV���ͫ�����S9]��؞�o�F�"�S(p���C�Ҭ�7������#���x3fy�n�h��Mܬ~t(Y��2PY3Ӣx�"a�DCn������@]^s^�8�2��Q%n��/%E�<��+���݂�j�2���+Xͽ��*WB*��M%/`W2�&�!vlCu3���{�<��H��G�Gd��؟!��J[%����"3ܲ�q3�o�#��]X��s�}*/u�q�Z�/zb��9������dgg4k�,��[���o/�p\���Y�P�������b��pEBh�Du1�[}E��Z��y�|�Q�3q̘A�&
��X�g���k��͑J�7�0���G�99�
��qV{��eQ�^��$���bCi���W\n'he(u�7r��D��K���s�D+���Έ<��=��̥PV`^�vٮ�v �㽬�5�זd�]���]
͍�g����lg�:i�9+���I��|��>����͑ΉÃ梱Z�70�%��&�{]�Q):I��\`X�L���EF��uN:1������h��T�V^\����u�}��2fR܀�HJhd��s臛��W��q*|�����;}��h,=2�"h���%���[���Ǳ=�G����D��C^�פT4���ȸ���\\��y���^>��i��A��A��:�aؔL��D��ľ�b����xر����x(V|G�#��恞��T�e����Z��Թu�Ρ�)ywmp�0�O׺�������W��
��.�K�V���
T��(
����E[��;k��dˀ�a������+�:�l��N�UY��4.Mʷ���)n����0��3�T�U�B�0�͜s=��%��BU��+��Aj'��JqǤ6�<�B�P�/z��+��9�v�xF�.�TDA���n����oE�G���%D.���t,��p���]OQ��驍[ݳ�cޫښ|M�ݒ	���	~@X>\'��"o� p߇��*��n�{yqZ���hs�\��H�5�t�.%w�Ӑ:+�v��C١+��2��fI���z8���`�5<K�Em�\�ߛ0}��8����u:�^9'��<p6tE[y`�0�˾³;�w}�/�.����t��B:� ��[7�����*2���H�J������J�I;�o�q��l�؆Ђu��
P&F�;B`iwYSb�w�'�l�#���̕�{�G�7���tI��1�]^?;� �~�%�{���]�A!F�W��C�q��v��CI�LIZ�=9,���3=9�*"%�wQ�m�;��4����i�xm�0Wq*���T^ⷋ��Qx3�EFGI�Cɥ!�\/���~(`N�Π��px�0n:�hc�w�썷�����Q�P���δ�3�9�Q6���Hv��P���#+�+�nE�F���i,l�-�*�d�n�I��7��uP)R����+�`��V���+��+5�Z�p�3P����|ya�8ޫ�u�7��=b�ҔZK�}c�YRX�ϳ:�t�,�7���o�L�ׯ� b7Xu��Ʀ.G���a^	�",��­��3��NfJ���W�<�l������i5�+�+"�Yq�+�&�Q=�R�����}�ڙ�%i��[�Z�-_W��]���WV��w����c��*υ�U宐j'����w��B״��n҈�;e��/Q���K�Ǽ*�#�EA[g��ٕ���:c�'<j���U��|���Ȧ໳�w��"E�ݹ�;+zC�Q�5֙�-"!E���EeI퐲�,���4x�8�V�{�s�o5Z�Qy[}nq5��x͎�8��̓��n���/��2���}�)��~�aј��e˖kY��ʅEz�9�j��^����EM��F�҈��b�%�u5�u�s�j��� ������S��?��� W���4�^��A�q���s��״Ӽꋊ�����yk�&�b���˵�V�ʕ�/g�
�3�{�+s�,9HÅ-voL�Z{R����!G �+�� ]D�n��;�0�RX=�z{�9]��-��Зz�oT��5��J����^��IJ?g�ϕ��	GE̊j��!>��\O�a��*���Y���ŕ�n"Ct�
�و�P��MBy;X�`�E�d�c���ۏ�ĩ�
[��"�z�8	���i���;�b"/�0�㾙tn��L)'�zsսݹ[X	a"���C2Vu��V�f����g`Yה�<�l/�UÅ��{�y�Ә��>h�2(���٨Q��I�v�D��[�d���]�Nt��2�.uE]&\���@��Y�E��h�ӱ0$�ٰG���`�|޽�ʭr�%Pq��pW���2hf���t8�DW��:g81�����m���v�#K��C�8I(9�|����v3pvpE�J!I�V˹q�ҵ����]�}�{Ջu���s�jC�2ϑ"�q�k�uY#��T
��b1�ӈ��-�jN�V��n���n���A	��`l���: �'O7���+� ��V����#r�!W�q2��1ڔ+Dd8P�볘����gt�X�����&
��.j�z"�Ì�é⬢�`^̹̿��CڿUB���iC��!��� �$''ʷlryF<U1)b��ޖy58�Q��X>a�����­J�f�8ݖ����u�6�tU).�]1��͕����P�3|�)�	'T́G��G)����+���_	U�LN���X9�����-�\y�Z�i��ȥ�����ެ��:�͎�_][�K���Պ��2��[ר��:Jk�uϹ#}��+�������o`#�a���&T����*��o��x��ڝ�q���=���CA�+7������9�싁���[yJ�%�N�k Y�@ZxVҁV�b�;+@�A�8�>���H1�X��V��D����M?�R�b@o{�t�&6x��n<�"���K���і���!Y�P+����n�6��O$���Q��CǬ7��oY�z���/,<Y"j���Zp"�"�H��
�QA��Bx�"lK�����1~�U.f�$�Vf�z�|M#:�$W���y2Q/�Խm�=�����^Q�,@W*��]P��,�T8��.�UȀ�z��w`���k�#}��|�����Q�T�N)��.6�T�>���[�L���!O�͌�=	}:I��NFd߅J�p/iVDՕ��\�^�wV�бw��^l�_�X����]Jݠd�����+�^�4**
�}t�&jc��L�(R�ܵM��2"���09�i,���>͒ڊȶ��N��aDl�zjn5���MN�_s�=t�	�G�"��
"'��)�c��h<˘^��3.��a��wS��(g�x�8�ElL���Y[{\��J֩��Պ��Z�E.u�Q�k7lR/[x��Mο�t�h����ȸ��<�i;�]ԁK5��f��2�)�]@t�����
��n�;:���;tg]��9Q�����͗3����o�u�:�Ro�bˍSl{��HW�ݟz����A�8�q4��6y{�k��H���ybPg��̵�;+�0~y�՚�föu䇮$4S��r�X�k�������u��m�3EͶt�;��(�L]�hJ�Sˑ<esWƧ�v"T���w������v"��OV����D\;Y԰O'�b�N��Vh:WgX��l:�P.9��¯�<�5�6}��dET :��eZ*XҴ���q\S�FnS�q�����.�����Y�/�>�.����[(�A�ٴ3L�O��=^om�7��	�pk�鱬�K�sq���fo�v�����p�@�o������{��V����#�-{N@�wh)��w�/i=x}룦�!��2	��0��e�6�[��r:!d��1gc�s�����c4磠l��EN�x�L�u
�0�L�s�Y���{�P,�1."����H�`��r��YK���/B;R���;Z��K�֍+�/}�,7C�|nP��K��oJ��DS^�ق�σ���ߖ�����$ceu�6;_:)�@�e��JXF��V�ߢ�'0����k0��O΅gu�GC�%-�p%�΂5d�;�o�v��B}��/L�~*�(���������Э���f>�j���7�6/����%��owb���s�����b��o��a":�N��(�����ѽ�`xJ��������~�(��r'Sb	̐�;���\կWXD�Ռ�U��%�΄0a'O���ν����#���r��SX%Ӱ�����U�X1��n��å����\�׫B�j� ���B��:�ʰ�ˇ�a�GA���>�\����B*ϔ-S�g�z�Q��9��-�%;J�P����G�W��z��]��p����W$.��O4s�
W�sP���\!�V��A�J"������ĳhaҜM�S��m�5�L����'���0}��=�ƶ<t�	�4��|���DSJn\�	�}ގ��K}>/�A���|hx��~��蝊���"9ԡ�k��Upwz��Xn6��g%D��=ۗ�����Ni�>شt��K418�z��zW=��.��ѩ6��Յ/������{+�1E$o$�.��+�T*(\�;���lWAŉ뢦��L#�ð�5�I���v��5 3�m�!+�i�X�ձ���{��#��1��:=�2ɼ����{��2+�i+Əi4��6����B���K�^!-1[�P7G�g_<Bh6�n�d�������)�{ǃmk_[2w$+���/=n��sP�.�[�Ir�=JQk�]Z�n�o���'w��}	V"):U&��WW)���^��T�E��^sZ<�S�Yb���(��N�w P��qR��.�γ�9k����w�R�����K�R��z�g�(����p��H�����N�ݩ��M3�z�[[�����ٟ>ʲ"",�ͭ�lE�e�
��$��)�����t;���͋��ʹ)�@�fʘ���幺�4��V����0�g���>�1DX�ʼ����j�fc-��kع��!Y�r�V��>�����`I�^Wˤ��[|��G>�!L�[��A���
6;��y�J=���yu��y��ioq5ݷ�Qht5��v���9*W9�bdxN�8=�an��W@��U��^U�W˯�+BU�շ,�z���/A@d�,�k���YEE��-j�AL�����}�ݸ���[ǱJ٘�L;���x�]���������sU=VNL��Ԙ�����t�̎���*I^2���qh�}1�����s�+{vօ�[��-%�dWD��:�j�*�c��+�Lp�c����� �W��	#uĺnU�g]��N��2���J�I-���M�Q��ml˰�;Z:�VU�pY��P�4b"7Ն2.X��(�X�j�±��6��a ����Y{�l���s�e�S�������{e����]Wf�e�N�7n��%�p:RՇX:#tR�ì���Q2Ev:�Uҟ���\T�Ne�N��DfH!6����SË�� k��6.}A���_��	ҙë��o��뙌�rSCUP|�9T8w"#�V�i]���;�lN S.��'!�%t(���Wײ��toq�u����x�s)�h�A\PE��oE1��/�P*U|:[χ4�۷f+��`|	�H������U��Er���1��	�%K��Z�*�l|>�(���ƱB��=��U�6\��}ը1ґ!�&T��'δ���S)zt㐤��- �!��@�����5��G��#�p2���[B��&ц)7p$f�i-ì����G�6Gn���Ō>>����5H\+@�8WE�5�J���Ն���Ehd�(�]�J��<� NM��W�!s�D��Q�6�a�cCP��=�;:� �	�(�� �0[�]��3wbq2�MM8E<�2��.���q<�M�̎C��ӡݙ@GR�n�Bg�<�̨ O��d�ռ	�H$T c��;W`Ȗ��7$��3��
$c�$� �ܜT6�xN[|6Bv�W)��!w�T��ϬL�)��=����k/۸ |8p�q��Q�mh���"����aZ�m�Q�+[E�e���Z��DD�e��V,U#j«iPQV,���UlKj�j�+T�F
㍶(�Ѱ��+ib��Km�1b)ED*T�*�)Kb�*U*���E�E��Zҕ��4�T��(��,U[m��R-KJ��K��2��mR��уKUQ(�����*J+J5�ԭj�(���T���X�Z�ѣR��Z��"[h��Z��Z�kZ���+*�Q�Rа��-D�kKV�&4��E[JV�UER��kkJ�e�+��{�<z��<onmҋ�4k�:�E�m[b�r��5A�e�%�R%ץ�צ����ڽ�+¶s�'���[�n��Kwo8�_Lb��ڃ��3��8@�^~�Tȥ"���y�ܨ��ut+
��/g�
-�Y�c�J������X9,��~5�ڥ��� ����ᒾ5��yf��؂� �8�;�<Sc�.͠���7vҪD���d2DB�r�Y`��e9�O!,�]�ux֥k�2� �����yˋ8n"[���*���*�|0�yU<�^\���@4�y��R��X�ʁ���C�l!Ը;��O�VDE9�����P�0��r:�A�w{����2�����X�˰�?@E���0B�s�>�����Y�F��"�]Y��[��ݣ9�����׼bX����9t�ɒ��"����g�:f{5�i�[����S�{F266��6�B�+�2W��du�
˜�5j�3�V����AJ�8E繜nfp8��8m����zb����f[��p�y�)W�I�ݚ��HN O{�47~���w�e/
��;�j�u�ȹu��2}|��+ч@�먬�Å��WNm�u\��!\�DY�0��k5<s��W��n��~GK��
Mg�	�0��q�jZ�����b��^�Ԯs�#��>V��/���Gγx���=����
��9
U�K��Dv#���C���9���B�hh)f��|0�qC9�E{��E�u3��V3��gL��v�]+:�˘� >���Ͻ��1_ެ
�P���B�s�­.*:"yn,�+����^χ��db��`��{�'�a���;-%��_#�<#(w�]9_u���:7e9p$ü����4�ګN&���e��}]��h�S__ڠ_$�H?n}<6����7��:	s��y��ʪ���E<�Cr�_d����EA`��ey/P�Z��,� -<+cU��;�֮����Z�QRL�0)]g��ox���FT�Q�.dP�$o�LG&�t�Jq�H�y]4�fvB�*n�O���[���8!9؞���m[��D~[�R���s�{M��I�����FVu����j2�x
�=WJ�(�^�|{��xBs0tD6�u*�f��{�I�U���<r�dB'�x]���Z$\lD���B9����5[���:�=-d�ǈ���|���Ҁ"�#L��s�Y�ڜS��S��T���Nx��ӮO���1{]1����ܗV/�>�V�6�e�]�T��WY�Y��t�E�(�][۴X����7�ӻ����Պ�}4f�3�;jL�cv�s���n�\���'{��ҫtx+�]��Q��)(��1����W��4���R����)>��rC}P�`x�*��]x@A
��{T�����)���S;�\<0y�e���{qUsw}K�R��Y;ș�G��Sd�kQY��Ҋ�0:n�v
����pt�����I���\��;�Q��qͮ��m����qA�3��T©���[N'/)�Ւ��Y��Fr�U�7Dc��EB����6�q��jwq^j��f�s][�T<�wf��2�LT00�u2�`\R}r�5C��T#�C��|�r�W�q��w7v��y�8	�cm;8}��Q�䪨8OBBɎ��J�&;."�eD���*
89����;U<��sWƧ�Mؔ��</��+�ڷ��ss�n5���M�Ǿ�t��Å��R��R������z��G!Gʕ�`"�"�)K�!V�ku"�.�.ukr����p�M@"ڭ�f�.7P*0��[�'�iE�Ji������N]�I��oj\V�I�B�����=�}ηgT�K���dT:EE�U����﬉;�
��+�\���"��B����K�3F]��n��Fm�sor֌�Ӧ�e�&�W���q5�0�[[y7���N�4�*=`;�]��[M��Ǆh�)R���Iڞ�g{���R��vc0F���:��x�\7�B�s�nA/��W0���T��o�t�]�f8'SS)NY��ք�Q��Vf4N��0n��)v.�*s���t��Z��oAI��;�P:�{��M6��Y��3^��z�X��e2΄�镛-����Αw�\i���ɊL��|%��y]��f*_z]Q�s�����3��λ6LXЎ�x�Z��sl�we�9١q�u�����]yR��V���`��r�n�YL������<��i,�Y<�]!�huGMOC�>ޛ��W��;�0	��_.`h`�[��,�E5�ퟺ,e*�,��E���<q�w�Ϩv}=4h���;0n�CF�=W����#�Z��ڼ�N�Re]�O ��>�3�6��q2悗ۣƢ���.�55E�5�V�/I��Gs����2����+~�]A�^zUpu�����Q63���>��zSۇ�i��:�~Y����ӈ8se�gjv�m �lB��T"ćl��P��;+;�j���Ӫ���fRLj�[�z���{؀l*����)^Vvz���g��>��>v�
��x8����C5�3���i<�{�QK�A��q��ey���s��1�4��U�;�sB�P�*�,[�9�/���]_p5��A�� HqV�Y��3�e^o��l�a�P��a	ڊ��H��+��Ǟ�n�ŕl�o�|ZR�+�B��z[�ಶ˹Q�5���D(�)
�V3"s�" �N�ӷ}�s�{)'���5H1�;ӑ`u������L��9��&U*�9��W�p��2k�.�Ә��.����p�%�P�v�~ɨp���B��`��	�e�����u�(�k��Jdxhkp#�����suHJ� gt��v��V)�[�tϪ�D��b�2���w0�E�9�u�I)cEs�����^�#4��Z��]09O9��Tu���W��yd�._v���śQW~��qw&���hԩ1���4tv�mp�5�d5��%lwY4�7�Vuf�ni�r�*6g�� �zJR��|�	�c�R�>�>����~��2�7��1Z�q3��B��V�za�~V|�0|*������aɸN��)��oA�w�9dn��Lےz,�,8�/������k�5�)T�΢�B���f"�!̂E�x{���v\�n��،�51��zml�|sNJ���}g�^���iG���?P�����8��I*~[��ŢJͅ	�+,�.P#��a�z�mD��UCM1�
ܽ�x�ex�78��ԇ�K#�{X��s�� p�i�O_G�yˍ��^�eJ��3�a��edO�m)��������Me�J�HK��f����Ι���4�Yɐ*X��n]��h�>��l��`���:�3�ׅ�;��T�=�2hiE�; ��GgmK�:!�lQ�ۤP�vG+5$���,��x"���U�y8�hm(�d�O�^���iQ�:z�E��]G���Ƹ�d�=�k ��p�4�8��n�E)��Q�E���W���SR�]DZÑy�E���!짽Y�^�Y8s�}.���W���<\������[&��V{�W�ǋhW�#�e��CQP%+R���˲+���L%Kj�Cy^PV��l���=,h�/=�/�|�yH�f�L>G�T�ˊ��K�A���C���c� ��QC,o�C��˯R]��O'c�YL�uI*�Mi�@v�l�c��ױez��NY���\5s;�:�z�W^��W]|=mx����6�s�XpЄ~��+t�Q��w�$�J��j`���t��J+;�b�^����郎�"��Ua��x�VME,�R�2��18VLD���VE���D��tB��m���q�P������Fh�Q���̍��a#�1�2�D>���ˁj�E�F�zNZ���Gq��ΩМ[d ��G��B
��
d�oB�*��WU��75�TM^d�^���ɸM��͠���K�v���ձ�G��vSk����>�h��{y�Es}���r=�>cs ��'vN�fGf���JWgC�$��Gm� ��xCdr'vB���';����t�LX�\�=�L�=�J�"7��{V�I��<��Xp�]X�iP��O�k�f@�A�7v=�C����|oX�[���%�4G���?��o2!>}o�Yi��~��\�K�7<X��MA;妕P�N��4{��yC� ���E�.�@DWJ�d�R�yX�e���5�g$E�D&b����GyE�r�ڍG��#�ʠ��܇�JI1^����C�W����̬�73���v�����%0XB2�'U~k&�ŵ�4��L��p��3$%]�u����U�z��1x65K��"kK�<iK��q��uW�{^�:9�ӝ7F�f�r�sꈬ���+X��
�ܹ��t�36l���c���gJ���x%T�Fy���.EOtk��M�Y7"Ɲ�c*�u�.�>�Q��0ϷU��*J�;�妲�W��b1{M�]�~�˕6��U(X����ai�{bCE8k�zV$9��z�Z��Y�*��^e�{;;�쳚��M����,.k�'t��J�4`ו�ϷEo
�sS�`s�z��+��x=�M�1W��,)-�A]&��kۭ|�MZ���˥3��x�uok|>"d���I�����spb{�.S��r�K�f��t��%�+ �E9�;�92'��3*o�Q�"�4�D���j7�n��|�	��J=+�B�I�z{�F�ϖP���0�-������~��
ḥ��YdB�F'`Du<���i%z�vtq773���j��`^p.7pو��r���(��4%D+��K���M�뺩��x"��X�=�	v
ηgT�K~@Xcϗ��hf���v��t�p���U�_��V��^��V+C��AY!��	�+��ncg���s+kČ��r�#���Asyi�#Ĳ;�.��
v�p]��U���t:��2+�k�zn���|�5eS޹JU?&Et�_�-�m�X�k�P�8}w^�s�K��9H��ڰ��2T��,���
7A��"��FDd�t����0(���������3�un5�^|у�Y�n�2x<���x��8��E\D'n��>(���]T&�!l�}+f��r饫O)V�hd��&���Q\L����C4��Pj.���U\�;m��Ҁ����]I:l�$�Kq�b�̣4�D��L���627b�Ts�WZ�]y�i�=���˿YI����gW��߇`��Pؖ�������,��9!|�F�����}��5����d^B�&�]��1�B��6��{�N�}X�m��3�l��ۘ�99�W��o�P⦻o`eNFEd�rhe� �r]m��_�.ͧ����Ƶ��ٱt�X=��<����fO��ɣ��o=�s�*#iP���C**�&���{��gն5Ttt>W[`3�.+͜��7捗�-�H8U��y��X~�����{=��)��<Rj_�N[�r�*MD?i�ĸZ���vt���
G@Xg���Jq�8J��x������"��[�`h�w���Շ��\���ច�":���NiX��y��z*t-���jn��l]) l��Oh�F�0V��bVţ�74࿽��/���<�<�j�������&Fj���V%��Q|͌�
X�*+ؕ��I�]�Iu�`����%��n��ŷ�.l����51���RUD=�E�kt���ݳ�+x�M����}��)V-��O<�����r��u�A��Ҁ!�5}� ����
ќ]C�p`��8�:��q+aRs������}d~��b�t٦d^?�z�و>�@���e_�="��ϳ��J�<Q�4mS��iA�u�ڻU��t���D��n�� ���Vx&��.���0����mX�`�T�9�+�Z{YK�Oz�V:vʽ�칻:�Y#�
��'���i�Ƀ}D黎v�ૻ�s.nR�W>`�m�M�ugp���/OQ9��\l�&@,�T�mT6mc�A��[�z-��F�Og���
�a�et��!d���]1ȸezH���B�>O΋��q�y���	Oj�||ȃm����fA��/��
��ٔ��u��\�ʐ����y�׈d���j2�s���D��<�gj�F+�E�����B���ڂ��O����
�7&w���P�!o!���2_��kn�����(״��� uHn������	N��:]&]^L��vu뇽���oY����p�E5�qo�A�r#��wl0t�ƫ"�p)q���ӡ9������r!������T��#��xH�׹�wł*��ʧ�[�cR�/�=v&-~�R�i_�s.�?=뼩����
>�ӑ�����`덇i�k�#m���ĚSi�bii̺5 ���QQ/�Eib�3;�����V�]�];5�h�LI���6Q|bO�%�&�%��-ךG҆ٮ g�T>G:j˃�ȃj�':=�5���h[í^L�:��xv_����*�e����M��m����Ӕ
�p����
{bL�;;0��A��κ�0���䵽Ϲv�p.Ŵs�Yf��
4���G!8��;f�t��g\�z�i������@�GEKz�8���Z� X�^�˲�
V�q��Yrf�D}��x��7xR��=�=�	m!��ǘ]h}��a��zCC�sv�n9����.�EkDL�{��7oq�������ڗ8�O[9R���@������R��AŹ�#��N	���Ex��Æ�3n��:��S��V>� �3	٬low�Zg� {OK|�`G�� �Hk:q�% +����Z�Wmn��]�b����0>�@�I�Zs�KT8l�kiQ�jr�F�cu�pnԺ��GhQAY0Vb]n�$d��Pwqy�]dV:�|��#�k��;[��E+=�n>�vTQ�җ]��\��"ބJ�]h��C��t����"gbV2�㬁�})���1蝍8� }�G�"��'G���gr-8��{�;z���q����Mē=]�V蝘�ӈ�6���1U��u�U���wM
��ẅ���h�X��-��y���Hٱ|Ɂ��]��EbM� �lP`�c�L#ftyv7�q �)���	;���d�Y���Ci`�ת�����[t��5m�D�(��`덗�t�Z鄷S�d�U�Ea��N��*%gT�@VӴ9]]�v��(%׷�N�u�l�:�m>9���	��%k'�"֖��5��d�g�,vG]�b򱇗Nk���;.�ԡ�a��xv��ݺ���,���P��#F�	�uxu�<xʪ+�څ@n�do���Op�Ą�혋��m�b�fSX{�]�������K��IAhWu��9��k	��1�we��ZU*=�I�-��j���	ԤD<�2��F�N˶�Η���s����-�'Z�"�Y7n�|D�9�!��3h��'J��Ǻ^�!)"v�c�Z�"���T�B�V�HL�;f�����a�|���7�.���˳cxI�
aGE�4�J�	yp_	�g���#���C»��ϧ�L��-��tU�����[�d�٫sx�M����RX�V�E\b�*nS���m�6�x��Q�S�@$�,t]j���y�&o)��U��])d��H��$�\̥���2�t�#[D����9��n���no��E\�0�
�z���ۖ� � $�(r ���V�m�-�YX-EeK,kE���J��-��[+m,K-��ڊ�e*aV�JZ"��P�k[A`֫[U�F�kkl(���Z�R�ѥ��ebԬX[J�E+[UDKe��Kj֌��Q*V�Z��2ce�Z���T�RҪ��h�ekh#KaDkr�H�UKJʕ"�#�E��*1�2�J����e4���#��Ѩ[J�s-V
DE�-F�V�(��ֵ��m�*��iT�h�E�H�+,���[Vڪ%Q�F�4��"VV+iR�kkie�TFUlKj�
�s1���Eih�+YBֵU��T[R����J"�����KQ`��Y����qmkJR�-�Ĵ��6�m-(�����H�m��k^h{ܷ�5��n�$���o���nRw�Ģ�m�ڛL>��V8��$�D���ꂯ^6[���r�}�mAl�~�ݩ��7-Gd{�p�*�B��\{E�Aö�fä�����O	@�����c����i��y��
K�=����;(�NY�1�G!�ב`�VLX�s�R�h��ӕ��.Ȍ�NJ62���Ւ�b^Ρ�l�}ힼ�R4h���%ЧX��f��C����:n��d��V��8�27V@t�p����W��6��G�&\ȫ^)M�1���ސ������6j�Y�J7�O.#=R���])c�C�8Ͻ�:�~��p��Sف5��{�vn��&a��\�kz烺�kE���\)g�ץ+oL�d�A|ݒ6����|���3�Ɍ�yc~DJJ������V�"�+��bP�w���j:]q�a�F�C�kΣ����v�a�,WA� �4|I��x�b�r�욌�vXJ6ۀ��3-�=��q������90��}P��[w�ۙB!l����h��3&���1�����m�� _��sѹ�C�N@!a˶�l��.-���~�����A�ޖA3qt`-�+�E�v��(q��AY�7��A��]ӥf����<`pS�%d�;�A���M9�`̵�~��l���{{���l�\��e>����MP�;rp�����w5^�����#�b/"O;�&��w�S�+$�w�����@H���E�wt�c	ɬ��&��}Ɯ��s�����������Nth�ΝH�[��0�o^��v�!�����;x+���j|���Т"�;u޹ٗ���D���h�x{�y����גZ/��f�a�-�ħm�ڬ�rυ��tL����uu���-�=��q《�{n3�ޜ�B�+�����"�����^e�\;���I����R��`�<�QY��~qg��ȝ�r�g�G�$�a'�T`�yNW�@��]�"_�a�.��Og�o���\a�Z�ګ��#��@��L��������q��6:�V��n�W��߰�L,R���T��\3�w/�N�c��4��~v4��oo�	R�~�:�O/Pڽ(s�P�xxDk�veՊ��]�|%_�����Y��->��Gԡ���9}Pb3�j��D�E縫�{��q̯1���j|�uO_j�R�=꾡gۊ��̰��_s��x�*�5�%t�X�*.���.��n�~���V5<#z�����~tD"^s �=G���*E}\�p
����3�`�Ժs6�wj�K�V@39m0	��Wd
��2v�-��/x����T�3+����E���U�R�+G�^p�s'6��J��)�o��>e�U�%e�=dQ�qiO�Ļ��t�y�e�Sd/���E�֜Ylq� �u���;,�Z8Iw�r�bK����}ֹ�}�8��շ��V��xu[���)G����������B�Cb�Z�*M�!�+�1smI��{���9�s�Tl����F�)�x&�Ul�%r ��g:��DT�ô-�5�w�f�
*S�]r��*f����6���+��=S梶"(5��T4t5�d��������w{�D��d���{$,�5���
/��4�����QY��:`|u.�Ф_1�Wn�sF�ξ�eQQ�9 Ԍ�*���C�ҫ�b^ǰ;;�Y�,�7�6�=[3���m- �=U�D�rDp��|4���[gjvƐ1�Ң(
T ��{\������y1�E��c�v*^�s��e�-t��'g�����;ʻ�'���=
n������w{���4:ޣ`5��,s+fT�\�A��%P��lW"�Kgk�{z=����o���!��0��>�.)�[�p�Ԩ�g�w�����R.�jKĲ.��%���\��~ev��@~���8<�Lh͊��}�v���p�N7��J[T������w|�4i�	^6P۳�:{��P��'�6�$'>�fB��F�Q̩�Y4���3Z�r�ax�P���wE곴:fq�O��	����	X�s��PK�}�ݪ�ex��c������=D����Ճ�v5��A�:Q�uPE���{��3	"�1����Z��x���z�͚Y�� V��Bˮ���X�hWX w�]DO� H�b��p~��fe����N��K�L&�Wك"�gO˸�N�V�{�Dcu1��[rY���qXA�Q;18T	�L���]��t���xvel�54&\d�[t��7J�"�B���b(��y�������M&�Uuv]E��(�	���yD8
�t؞T�^�qݾ�*��� �8�_�����[$q�U���^b#�{Ք��u�*�G3ʠ� w�- g��w����K^��x�#��W���������7f�O�4���,p����G�L�t���jUK&�Y�} d}�ڥ�����*�0&Ǥ>�	�,I�̜�#�{2kH}���Q߶9+��hq]���>&Q�zʶv&6J�-�Q2Pr#���+ԱX��jò�:�_��ڌA����y{D�pz������V����n$�Ļz,�;h�;#.�ty{����\{;՞�,۽����:�wy�G�5�dC4Xκc��f d���X]]��Q��-�So�(4��fg:�8rV5�݃5#��_=A�����G�C�ؗ3���ϡ!�� 3�|�"�H�>��^-[�ɾfr��j�\A��b1�ӈ#�)���[�A"�V���f����vs3�9��@�����9�OT^�b�>+ �Z�]!Y�a�Φ6<%}�@-�Cjn�f�t�	/�PN��XBϷ���H�_���M5΍�`�w-&iqQC�� �yn�t%Z��7ۓs��&=4�MAދ.�c��7���`7����ZD\].��p��1�J�������-��k¥�;î�T͆��-�7��2&!#�����*�2}�V��m-v���4�)6� q����̮���}=�H[�ߣ��E��l�ut&=��!���՚�)r����LC�����;d8ݗ<�t6�FT�Q�����a#�{3�Ŗ�����6��yW�f �¬DT鸘�K|A��
��
��p(Cs�=a���eܘ*�bwqo�1��(��0��8z�%�t�qu����`!@פ= �WM�:�Ǝc��K�J��+�5���V��,��w�cyFa��	�YB�K%�	�-(�TO�f)��̾
 ��q�B�TV�CES��UoW^��q]�:�Ϭ!���ElS	��(V���Ě�_;}���f��f*�x'����Y���|�M�|�R�ܱ�Ļe���g�{�4l���yf0@j�׹͌��1b�͚�)�F����\l�N�iȁ�n���P�}E��z�
&��E�r5��Og�'��љ�槥{5��m�KƆ�U��w���-�7D �F���d]�Fai�����_�_Q�^��X��l�k���ݛ��%^Gҽ��O��؂W�	|"�y����z�%�s}��R��w���χ)p��������]U����L�y�0!�7:f{]<��wxe��TQ3�	�d	���W�et���&�!h��g�u���������Uɲ�k�5����/V]�+ވ���Ȱ�oF%;o!Y�B��G�gJǝN)����Ľ)m���$���]3U舀��O	�z����XŰ�$h������]Os>�/��<9=�|6�މ-[4��\(�-ȸ����zE瓡;4����sWƧ�M؉)�����}��o�g�w̟%u��9��gU��]��EB��A��!VA~x*�L�73y[�w��6kfP4�p�wX�;���wINW���6k$����Ea�*�ܫ�B��wʵ�]eF��,�w��r���-�\ũ�h�ۦ���5˫iv���@b�B�k{0Wz[Z�]�kx��Wkk7977���Juޠj Ş6���,R��J���w%B���s\�n�#k��j�wk��ױ����K��t �GC_:�q�����[���i�s��2�A��YO��n�Ga��mM���H��u�XaVA�䋽9���~$6o��%��s�X�ƭ��쀆=�x�B���}�.��]��X.�_�Ҹ{������y=�xj+��p��X��o�����q�h2C��B ���{�Z�I��ۚ�ٚנ�Y.�c����R��� �p=�IC)s�J���B�5�&��p��!z�O99��,.�װ�z�M�*2��ʊ���I�@a�^γq|�z ����n�[��r��͔.;�0e�|���vj>U���J���Ї�˚R�"]�ӗ���Ɇԟpג׋Ըn����.�
BVxx���[�l]qs������l�4CV���E���۬#8<I/�2x���6��V*��a���mݼ�;���$W�V��U�Oi�}�(3�x���@�bW���!����g�EOdRݚ�}�QU�ۋ�F���vV�D� |f�F�t�Ӛ���P©�w,�vk���t��m5��i�9C����2L��-�k.���ӯ1��tR��ur�y�P�u�4h��:�>�P:�yY9��Ѳ�宐uN�Y��g�#b*��-\x����C. '�������pnT=F�[[��鰙q�'��7�'қ�]y��cQ���w�Z�l1D�63�G;�0�uϫ�TZsZ�A/��������7�;ł75rڽ����̩+d<�9p�C���L=9�Ƴ��'��r��ٲ��Uލ﹌���=O���v�8�����4�3]��o)VP��1��}Ҡ�Y�ɦ�u��<�v��+al�7����;�C���}mq�xɏ> t���Ł)��)N�ܼ���
1�T�\b��1s��vY@�yd��ň.�}����+.�	���:h?OJ}d��z�'��jX�¿�z�n�Т�3����P/$W���0��\���r�߽n�L�Kg�.֏��
��B>Y[2�a��2�&z۠)��sT�&ڨl��\r[�L��ܾim���Dx]L
�=�(`!e C�����M�yS�bEDct��p!��m*�� u���Yb�,9��vOt\ɂ�יy\F���W�a��w�|�V:x8���+4�ky#�{�P�K��W��c^�:�fUݦ����w*�R���G�5:��:�h������9���s�Ѻ�-��K��a:ᰶ]%�'��7�����a,��8�˿P0{~�7	�ү����3�%@z$*�PB��EF��N潃ـT��-&h�=&v"4@�5�ז��b8��~��E���.V��`(|`���h��U����	}C��)������u��E߳�O����R{�*��``��Y�f�0١Z_�-��R�΍$����&x�S�e[:"c`�����$��GI�k����QI_����X�O��s$�ޚ�H�y.;IU-Ց�.�b� h�n��ј���ό_m��O��.���J����{��ciDǔ�PR-Ƞ�{+<ݾތټ���T��Nul�v	}��g=�7���Z)�j�*�8:��(x9�����n��/�����[�b�7�u^�~�ʕ6�ja,������ٮ��'P��zP���¿�'��xS�h�]��J�K+=L���\����O{m
�6>O�����=�/�E���{`�a�����>g�wJQ��J-�V%:!��wl,��=7��2&(JU��\o�6�}��Z��"��bxdy���q�3�*����<��az{@d�������z8���c�ˆ��)y��w��>wyD����{�;8����6����YOu��
��4]Y�����{Qu�B�'��GX�lY}ӵ�yߕ�fW�|.��?b2����l�H�WR	���R�tf�_Ol�z�8㍔B|��d!�Z=�O���w��8��� O�.�^�#��T��Нr��t"6�*<[.g���b��ѝ��ef�����X^�Hl��J����M@�s�B�������#sv��y#z����H����!��Z�A�zXT��x:��{��^���*�D�w�FEZ���s2If���� �o��2��%�U��_��-�D��.�6�Ѝ���,u�P�EyI����-9wK�L߇d����h`�`^����-`xS�%
�U��0U��ܖ�|����<�7�ʽ5sLa��L���!H\�&x�Q��e��y����Ը���@lt�پmo>��a��&.�`=g"Me8t8�ˋ	e�@�@oM6n�׺�Y��`o^���DY ����h�T
�,�a�Q�QȬ�܉�* �4�Ŏ'���]���L��dE��p�~�N��لL`�61=V�|�����7����~��ۯo�$�	'���$�� IO�$ I,	!I� IO�H@��	!I� IO��$ I��$ I?���$��$�	'`IKH@�rIHC�� ��	��IO�H@�hB����$����$��$�	'�B���PVI��Bz���5EW��@���y�d���F��xE 	  ( (*�� (P$ }�U�
UBP$I)U
UQD�ERUDQOi�@�..�JH �UR*�IT�EBKѤ� TJZQJ��2\ڶ+C2`�3"�4$e����5��V����R�%Q� .�l�a�fcF�V�[2�A�E��Z�1feM�T"��HY����jKm�ȡmm��0"�e�+dK"HU � v�"�a[i��@ 3�    �0   �;�'n��v6�r��T�DC� �����-9�v�Wl��hjK��n�Uifkv�gmZg[NU]��Z��ItS ��3]"n�k�c�ոۡ�Z�cD��j�j+-�i]�:m���e�۱��[4�EAUC� ��R�f�4,�nn��vŶZ��u�wu[;2gsws;fSsGff�h1d�T��p s+T*Զ��RQbc6���X%*ҵ�&�T1�ܲ�5%��kZ�fIk�F�����mZ ���*V8 ��(�-kYl�6�3llQ��j#fъ=�   "�&6�JQP40��b S�R���C@Ѡр&�� 昙2h�`��` ���S�)U       $�M'�=&�4L��#A���R	OI �(�`��� L忇W���=\�­�e��%K��.X��K���(�PA�?H4�\�*��b� ����ĕ ��މ.�y�~l���G��2C���@H���X�@2P�iDDd�D�HtA�	�ه�}�\��������D.(�`��Z�o�o�7�U��l2u���i���f��m]5ȕ��Ep+FJ�*�D���.�n��:<w�+�.��\	�q˭���wtpiP�.Պ�<ZBM0�#՘^�d'�Ȱ�&�!gv�hë0^^�����gT��WA3c�s3e�]�D���p�Z�L���5�.f97q��VX��\w>b4�`m~���������6��5��J��x�C ���ۺe��vZ+�')�Љ��$��x��Y�zs^�[э�iX(K� f;Sv�P�2�������{Z��b���f결PN��h{�r�}�8 �4�^<v��ӣ���6��qm���Fĥ>pĆ��*���(�bM�I�T�#��"i����X�2���\T���ѣ�$@�*"k2w�TJ�j����8	���n8�P��VM�+)�$F����� Z�;�]]���L��+ -e�օÄ�s^���@�F�����2�9In8i^U���,�MKd���`:kUëH�nPy�(f[�C�k�4��^:/������^�#���yq�Pƾ�{��Y*Cv��KSZ�4omB)��!�Z�Z���v��u�h7�Vլ�wXM�yaY�yہ���\�kmW$t2i��6�4��.�Źn�iO2U�Cr�yN���J���)���휢A#��7���M�a��y����-m��.����*0l�t4���0#���5N�A�7���۸B����p�m�$�\�a���Q�h�Mfkywya��F�˙�3<wz]�K� pe����vTׄ@b�,�̸w~!
�n���E��8��4buma�q��yP�f�De�5�P�W��lKvvLr�7����M��j�eZ��GH�>�0<8��au�C�����x�O�Ov����x�;F�N<ERe�YT�����x��"�fU���R���6�IvbYR��K@.�U�U0�0�҇R[����`�$5���7Kʃ���)��B�m�9&ҭ:r�$�Z���Ea�n�.�#-M�F�҄X���l��U��F�ܭ���j4-l�1&ooV�z*�)�׷+Ma��e�I�4*�����)�3[�0�Z�&-�*�Č�x[m,�X�),gU	�*X�!cT���K��F�`�ψ{�M���[V���L�����4�����t��xJ�ee�(�ae��	Sm�6e�B0����@5����X�&�3i�ˑ�j�t�JwdK��r�)�h��m�+`j�{��n�kC9mXG!Rͼ�wl�tմ�S1jZ�bəW��	o�ҍ�/ki^Q��_,�#.��)��V]꼼Q�F3�&ކ�ɌV�Xu
���!�чeݑrb9����sPa-�o+6��5�k̴�C4��M;��VЖ#*Re�ܡOD�e��Za�[Qk*:�n��c.��u3wRU�(�ܘ��7r��3�oP�z2��6�=۽���WF�.���i|�ך`������Ҳ�gQ8W�
��X�]�f��v�H��3S���J�v^aWb���*;���̘��A��Ј{L���J����,�Ő	`S�m-Y�*e�mś��lkQ/8�i[��sM����!v2�!J�u��\lͰ��Vj6�+uݼT��|��7���`[m��+���j����	Me}�a!t�d��6w��XU6-��r�l9x�n�.3��n�ұ6A��XS�=���*��{��a�koV�ۋ[F�ӽtZ��a���^��l�D��e�.�/C7�5n�FT/e^��n9�K�4�̗k/6^�_Vb�#^�Ď&��G{u���)^��q��ݫ�074��f�y�Y9Or�ҞMv�F�?`z3.�L��R#)�چ0żZha8sYlD�I�F��؞se�dR	�3�J�-Wz���+��$���L�@'�5L^'[�A�Cz��Y�W��l
 Y�Ε�|��.�4�Uf^�[�EP÷%�3�mhVȰ��Rd��b���n��jœ���R�Ԥr����kU�9z64V2Ry���&,������;2�b�YQж6�k�kF.���Z�ZM'$D]�j�G8em�tO�	Y��˽7V(���x�R�©R�mb����Q<�#v&�0�ֶ&&vPBM�g�N�q��8�#c��i����-��X\��v���]M��Ѫȷ��%��Ooj
9��P.�����F����F�[6����%�6�E�6�;Ϭd�X �,��n`p֝���	��f�y�Wf�i�G@��&�š<�nhҒ�Z��H�{Q�l����,%�N��t���$���RbVX�1�z�{dGt5ٽ�YϞ��L�W���ho�^m�u��;�; ]��g�4V�g�u�k��7��P�h�݋�)V���j' �ԅ��!����˭���Ԁb	��Z�#,�ii`�>B��)�I��q3�Ú�ѹ�e ������Jw��+�K[�B�����Ci:C�5r�e�u��-.�5q�z�4qOm4��GR��ŠƝ򼫠�h���(ݗ@X�1pN�{\�WHƅ��]�{n�Sm��W�D]�]�4۲�� M����N�ctފ�@"H ɈR�[(޼Tb/*�/+-��6�
AM�Eؼ:��(��cl�R�.Q�r8/O�R�
�q��'Ĳh�e��e �k(�kۢf$� G4$�7+�>	n��˓p��@usm�ͱ�mcm��,m�=i�G8s�#:���5 䱆6�Gt�.��&�n��*�ZU����R�`����ҬJ��u-�{h��tYm�J����6�p�7vbzU�LX�&�(U�P�b�V�
�y��"!��<ԑ�u�w.'�a�T�77W��(��P%I`(�ZO�$�Nf�Yv$*J@{���12���Z�n�CfB{�c��ʻ�ncM*Ęgded� BR��fP8卻�I'!Z��Kvt����ͅ��ă1nI�k����$TT�m�j@���*[���N|�Żw,�pKF�Sv�u����h�q-9sq�ŘM+Շk,e���%��I.����Py�!��E��F�lfT�H��Hf'vv��x��6�ڻ��;;NQhʻ�����j��ףIV�[ux
��G�OK�F�2��Xۈ�
�*bZ�|�����{��E޻��m�K��a����ƴ�QYmj�w2V$�G�K����o{s4}�G�?3�	������`�	Q��f�[f�a�RkE0ݿ~&�e�3�q�6�Q56
���c��!�]֋�"��7�4Ԝ)��r�u }wjI)I-����jiVt�������E[�pbұ�䓚���k�Q�%n�˩�4�B�r;죬�v�8)^r���1�O ���znY�۷�����;���,��|zc\N:o%��؜{&GS���e8h�\/��<W�(2�����ĆY�je+���aЩ��O_vᨨhmt�-��0ʐ��3{�@9��-IKok:l}r��꾸�܊0�J�Ӵ ��<7r��k�X�C`\V�3ԡ���k*�m�.\���P:�i�{�;����ɳ�lbh�wG�|c��x�5YA6���l��B���u,D���Sa�􂯑�6�v�r=�	6��6�]41Tg,_]κ�A �:�c���y��,����ڨ7��h�HѢ\Y�`9�u�Iv�/r]BN�����M�;t-��rYL���fN-������f�~�t�Ch.MJ4*[��y��F4N�����K�˻�Lrs۽-ǃ%��n�!5��Q�Q�j�b�h<�f������qOR��\
�n��I%LP��3��,�[Q.�r���:[ǃ�����=˘��u�N�g���[�ɗ+sE���u��b���a�ۣ�������:����m>ٳ�;JA*��Ia��H�5ǳP$ i�{q�@��̫��{�3e7Q�w�E���h"�;��bn�.��a�ʆV�6�1hͩAT�Y'$�59s��n(��[t���Á�1[�bA:�wP�Se��U��S�L!�b�.fh�x�F�/F�=�x{��]��Ðۛ��Hw�y�V�V��o��x�'*A�E�鍁��m�4�<��_	CΡ�����rnZz�^P�@lQW� F+��"�D.��2L���
w��"�!��u�v�u��(��刉�� xvS�;�/1���K/����k��]+]F���V���2'���x��淍��ٵ�Q�}���Ve����0:BR�WI�W�ү��Gw�w�͔M�B�J�tF�hl�����9u�A��h<X3�eW�w�\�ޓݹ�e�4X��� ��>gs�f�.t���Kz�,�O����Yx	}v�.}ڗ:�nu�����J�����9���]��-_W\ԨN�x� �a���UН��Y�M���j��:ۢi��+���ds+h��z�[{5�|Sԟom=�t$�p�T���8�ec�)�	L[\*�.��1]B�;}���ަm�Dm%�+׀CV��!F�����\������5^C�S4����q\�5�qt� U&���/���OV�&�ݧ�s���ӓ��<�@��ߺ��v]d5��j˖ް�q����
͗2F��Ċug�gU��}�Z�hP\E�JYw]�rQ@$���ix�V��ɢ91��z乪��J�״Y/�(^��������>ƨX����騮LY�]�$��nVQ9�r��\�`�Y:nΩ|@�V1=�y�v	*;��U��UtD K�]Eu��v��~a�Uv���0��2/z�u�ެTħ������0K%VR8v+�n6e�*�Gط��U���6��4ӈ3Z���^Q:��e����Y��3�� �E�)��0l��=����Q���noi�y,�i\��ud��x�;�s&Ij�q����S�喳+ ���M�]�F5-��]Ek9X����r����᲻4�vq�97�x�Y���3	�T�ihh���n���yۏ莹� ,A�]�vWc�eէz}Á��KNڣJw:��=B�y���*õ��Ԇ��.�4�EwtY!f��­����u`d��f��-�v(d����x0jZ%���g&�V4���f��=eV(��{XB��LKn���8�� dT�)�8�F����QǺ���V������S���ؚ�m����Q���*9���U;�t�Yb*�/��<e�uy�u�q61$|�6�����������[���pw�e��m����"���%�R'72�qq���$H���Ŏ��{�.��)ڰ����1�m�A����*��x��콙щdЇ��;�͞#X��Bf뚡�h]:����ԍX�����Lj��F;� ��]@��39��j{��N�z����e�H7i'�7M�����c7L9ul �ې�W=��`�-�]�~����Y&�8�y.ˎ9K�wt��{�;R�^����٩���K�U�8���X��U����d]rNbCe���$t�Jފ.���Y���^�B�]r�ΰ�
Ky,P�q�N�j��;S5^�r`Z�q蚋�����SLFAg���FX�,P68q/���2m�
fb�� 3�K�\*�ֲ͗G��])�(��m)�;�W���.�3k�����)!�i�gBm�]|e��)$�zڥ����ہ�+E�ԇ��:9�����u�t-6,��vk�ޭ���G�`�x�! 
��"�A�۾���ظ��Pt��X��y� "��>5c��;8嫜�R^��e�E�m㳻� o������ɫ)����mB�Q�7@��r��8hY�[̳3�o\��06���5�fa��Q���Q�,�Ԣ�|)vGYm�&�ќ)&ΥlZk�����B�t���j��P����
�NJD�Jx��N������5�s�����ob���W6O,)�����<��;ub����l����s}p����S�ɀ��37(���06&�wAL�B{�EfW[x���I
�:���M�D#�8�ڥ�A�M���G��PYv帻�!�j��B�LL:;F�pw U��Orڷ{��\VI�#+{K'��x      �t²9O��/�|��&ђA��$     ��@�� �5�F
R^nI%�h��9�C��ŝ:ӄ�-��.ap�9ã���w��[�`O����&�3��Gqչ��y��)<�gӝ���gX��Ʌc�k�'.Ly	X[��hH�[�M�
�a	&��r�� �a\�R�n���=#]�e^s���Qs �7�P f�����P�R��3��E+%gs��t6��}` �  b,KHնI���0�mJ�_iJ��ΏGkdEZB �8����G�Gp��< �85.��,F�� ��� /�p�#�� �  �    @ ��v��T���R��E����RI����?�����v�ն��0�v��ࢊ���D�T���;�wa���3�IQ��_Q�G3��ύ�xݩ.�K�]q�wg������n�Ί�,YJ��t�fI�l$�2�����]v��6
�PWIyf��4JV�i��)v����݋�C�t�����U��k�n���8^Ձ�)�I�BKۚX� \���]��>���3����69`�[�T�j�a�1��u��aM�ߺ�Be��:�0�2�2�]+�����w|Z�������-k����f��ꂭ�+f��\��FT�u�윾�: ����[�ؼ�4sl�l��#oV�kL .u%^;w�(�&n�,P�[r���e�ce�##���^T��aU�ʭF�2�%��^5�*i�D�ٓ�=7)��E;x��C}��G��\ZYY����P|.cYQΈ�HM�\��ԶE�Y�1�vp[�=�/:_+��+�����6�XE�"K���΋�E�K��|��+JMk�%�=54�[��t>|_Ңt�g=`e햣�6�e[��,3��b�����0�[�bGT�j�Z��)�)�ܗ1x!vm$�Mt;R����k�&+��\�0p��'�b�7�Eր�^3h�[ڴk����߯B�.�Kk W`��ʲ�놛Lʳ��=��j�ʺ�����+��hI��U�OO"��Y��V��s�Q ��Πn�8d�/�����i� [����/:���Y�n�f.�r/mwSŰpü���C�ܔet�:�����e�<��o`����āۼ��R�ʊAձ�d��V��^
cD�>[��i]������J.73H�.���37X��!�P��ֶص\�r��͌cwJ�hu��۷�$�Jմ�f4ֻ���.�n���
��P��*=7��b��=׺m^6�R�y�[WDs^ޱ�h
�\L��8ڤ�nu�u��u�XnL�&S�z�ҝ+�J�&�&��O2�mZY��L[��v]��GPv�5��"a�1
jU�G�o��o[�r��D�"�Zr�ns)l˳{V���Oe���w�D������G6�*)���x�C'M�1�#kB�J_L����nP����;0�\�1\#A�V)hv�t�A���S�_K��Rf�R�W�&�ɰv��ٕ%gϭ�L�8�,��r��;@��x����C$B��4T�\�U�]C.��샢l�eY��7h?��au�|��o0��f��Rv�R�F�j��,���,ΰ)��78h'�g�V�}�X�p��\ՖY�.c�5�l%���f�_���C+�Rƀg]kSw�AԻm��{�S
bSf�[���9��M8V�v:b��ϣ�zz��W(��\��vn�q�%���^S
b�ο���q�d�x2b��7v�o)β�����a�{;&q6/z���u����Z�tW,֪!]�Ԓ���Źk2à�xv�E�+/�<z���Ծ��1��=��]����t��^s�г}{�ȉ����	�����ZA]:ͼ.S��=���m�,�x�s�f�ѱ9�}����kV[����kv��d�o����u�r�tu޵���/W�Y�.Ķz�c�])$��>�i�z��"��t7r���Zs-�S�y���77>p
)�u���2𢡄�H�xFM�ś��u�"�cY(+�2��Kl�r��,����wM�C��t��I�����NN��s��t��\f�s>�Ru���5���S(�fVe�Q+�A�E�d�4��Y�nT妙5z/P<�.وj�U�*�.�l̮ް������ ^F�=M�{E�=�[�ޣ�4��f+aݚPM3��*��Phv�f���0:�)�PmC�j�a� ��+E�p�3���w2I���	�J�+�^Px�7����۱�2����9B��ScÈ+���h���d �++nno3uZ48n��h�-���]e�)X�BB�|��%VVU�p�3A��$��L�6���B͝v����{stN[�7V���e�����
���	�Dڤ�)ri�;q�lG|�Z��o[\�FZN�t<��z���G�vPy�V9Y�w6@왪������dSK�X��D�6[w�л�=���}���WW`��"9qz:����,w6̒_q�=�gHz+�"h�I�AIGxd��1TOP�n��PS��kt�b���
�tFNRi+l��������C���d� �f�	����k'���)�`�8]�Isj\�W��0�=q����*�V�҆ZeR�X���F��)�:��i��m�ZfE�я��8X�N���u]�g�,������:Rȅ^���i��Fu�X�['t��"-�6n�̳R>VRL�3J����hӫ,�ҫ��{N�F�z*�_�	��oH'7�c�C�m:-13�P٫�������uA�h��+�0�/8�7���;�W����Cn�f��wj���r*f�KnS[Pp��`��aѹ�A�1Q������h��G�X`My����Ezkv�c��x�K�V|��j����z�Vmi��lo7v�:��Q��n7 �Uf뢝������]y��^���B���]���:tT��>T�9��^�TK�lm$��|pd����Nݥ[Vw{�(���
�^;D�U��8f%b��x�U�1�ˠ����upE�k�N�uesR�"O�X����rvn^>��$�zj4�p�� ��k����z�����.��	ۅ'��9��՜��G�Z]�k�]ཻ(�_h)q
]��.y��+��TR�қ�͗m�u՚Ά`�����|��Ю�f�ۢ�W2Ŭ��������b얺l�r��b�7�S��U�Ptj����LE6�o�a� 4m�)��Xn�
�p���2�mڙ�HO6��eᨳb-ފB�0� �>���a��pVҩsUY�5�|K�Y�6��we�Y�Q��������k{%���֬��� �iwU�	 ^�m�gjn8&�=�%�2�Ŧ�}\Ӻ��M�]([b�*ɂ��o3��g_&�˷��3Sn��q"Iޔ�U*�:^��3i�� ����ؙ���3v,�6F`��,˾�"�X�t��t��&�%�ނ��"|�+\��Y�E���UKǷM]*Ʃ������nՂf��:*=]��q�U-�i]Sc�.�(�7Α�[8�n����S���SZ�n�?e�jJ��4�E� �j�^�X�e�ٙW��pn�
��]R��8:���J����ue�j���q��%�b�_WGaoV�����	�����"M6��+�e|*���Q�������sS)��;0�\��G1��m�y��j
k��q� ��r*N��Ǧ��&3Ed�[+RZ�C{΅orU�c-k��S�Wb���w�U���^ʺ&�T�a=�];�J<{�r��m��^.5�tC� �B�@3/e�R�Du�˹�H��i�۽3@W�u�	eDK�7��n�}6�w�]�7V� ���/����%Z��}�6���N�B�gY�����d옆�k'I�!R�eӹy1��;��A0r���?a�u:��(Fo����p�����8@� )� ��=�E�v�����      �Y;�--a���7���D��(q�:�.D�F�;r��\1$�*�B�-%��(��Bb]����$���.��1 E`�8����Ii� �ܑ�x�aY%+Q�wxn�K�e\���iT��4�E�V�A�*��弒�s�3����VZ-*�d�<��TE$�H�ձD�#B�UGm�VҰ^l��������F�w �c����?k�{�[�t�޴�����O��.��q�d�n5��$|i�������@W��0�~nEk9�w��5�=N�V�T����R�de"�����F}��z��mُf���D1}�=0�9���^_	�.��ǔ������O���A6Y�е��9y��h�ݷ=�-��W����\�O<��I�{۴�É���ع?e�=��s����
/�`$%�ޝwS�vMc��KBb�ߧ�x�&�~[0�h��No�Z|l�U����l�zER���O�jD�9o�H,������m�&�	&��s�RQ�h\�;�]8å��J���/5{��rm��x����9��{����ae�(���f^'y��y;��t�<X��χ�����S5R��z�h�M=u��ޖ*i���5S�ǐu«�+��]�}v�JI�]ms�Ĝ��=�R��m�j��P�����7�W�Ԭ�������P�n�U�뇵�vy#J[N�A�mIEVǂ����-�W����.�e�VPQ���^AݬJt������gWn�wb�6b��g�����2HI% ����5�V��3v���37nw���aQ�)�)�k��0;�^IB���D]G|�%{����oޑ������s5���/�hȵM4�ܮ�{o3%&��fmr�;�ssK�f{$X�%�c��.�Vy^[	�Z$��=��,}��~�_י��޴�ߗ� )�l��.����,���T��כu��r���u~llT�|U�ڜ�Ͱ�о�ѕ�8�e�WP�E��j�a�2�r�nB r_B����#j�tm��#��JJ{�Rm�Q�*$�0�-��OgWdW��I��:}pb�O���;E��OP�T�K����L�(��$��}\��Ug��)��:��,nt�v��s�&EG���iz��*Z�g[�u�=Vck���N�M����p:�.�<�׻�ov��4Xq9��Z���H��,�z���Z֡�%]�����<䬚5Ր��_�6=	�XX�e��k���a��Qc�s�����1�B>���
��5�?��̳3X���K�q��{��<�MT�+�nu�=$9��%�$������=�
7�߉��[>���`���M{H�b����"�b%�>���r�z��_6��g��'TuS����Գ=�Tҷ��~�D�`��B	ȳ����EK�}������� ��F:�r5�H���lf>�}���V筌����I*~b)��φ����{��RQ/��}Y�5����f���'�O�F{�eW
=�s#^� ��]s+��w!@V���<��}KHg,ef,{����3����UX��x�k˓s������nC��$�ĥ�Ɨ�F���ׯ�,���?5���ܩ���h/u����k=��X�����;��ӑ����kVz��5�674�[����Iy���ܱ�,i����>���Nb�����c�$3��*�ř��S.ΰr�^�wp���i҇������&�ت'�K˚s���U���F�u{��]�	���4,�nG�g�\�^�O˾G۪W���fm�r-��	88j�OB�gy��7�b"�_C�V⥰ʂs�����u"�$��I)A*q��l(���3�}����q�&�4Y�C�z���ߜ'}�gɦy��՞ou+!5qu�`g��+@չ��+3����3��������i��kY�W@�~^V��`�5�U.y�x�O�{<=�N�zI}�5����ͷ�!<-�鿎��gv�YY9��|;g����-OScS�Ǎm�F�5�;����[jK��o�]0�������n�S���n�@���^[V�W��1��eҕ����l��`[�P��S-�hL�!6�J�=M1F�-�6��a%6���s�N�&Ua�6R���nA�jN >�M�(���������~�&��<�6,�ޘ�U�	��L�T���@ׇ�I�ϩF^{=�lS��dt�ҷ�H�8r�����۰x�,.t�׏��k��6�Eزg���;�'��^xOw�)�m���Z�6�m�W�#�}��k�����P����z��$
���S����˴c�W�U�.U��o����m("���%���Gr��k��IE�0��J%%�z��t�x���~Z���{ǋ�?��lX���_#�5�=W��y��RU<��%j,�k}�TW�� �~���v�N���-�~~��U,�^Ϳ��<��C��η4y�@X9��`�RϵL����<u��sJ����2�����B��y��mu5�u�jfC+�iM�寠�)X�5��A� R��}�I�-5��,��n p{qZ[����d�o7�qZ�E��u���y���L�OF����s�3�zpv��V�5+}p�*��o]CX���t�Y�����Hf��R�\B�_���7/[lu�(K� ��7'&��~�1L>ۢ�����&��FI�D�v�F6߯Mz��x��^�O<w3=�`I���*�tY��E��Z
Ca�F?hC_{+b�f�z��܃]o�ȩ�(�z�w^�Yy�NA���+�C��bZ�1��,��w�:��7\��7鳗�0~Z�h������'������_��T��ݻ�x��Y#�+l�Q'��]��HLx���X�a���R��������4l1:e��[j�C�Sm:�=
A��y��-B�_d�{�[�p�U����nU��*C���Ӵ�aXŻ۴rwh��O�O����0�fL�F�ud��_hv�q���X�T�c�8n�aW
����Ȱ��^<E���Ɩ�q�*U��/n�[�.�:�a�7X��\
�XGK�Y2��Һ��;"e�xOe��t�-�Z����F�*;eu[ê��#5p�˺�V �ǯu}n���{8u1���? �P���(,
k�̚�%�;/�l{�˂S�0����W��]}|S����!uMעi�:be֍s�r���t���O��҂��:�t՘�=�q�c��Z{O�D!��Ч;ť	|�u�);��՗¥�<%�jVB��U���)]��'i�;��3&��4j=E��{�����r�e'i�ٍ���=��)c]v��F%�㋨�@��^��v:)���l{օ���I��T�/+y�\�y�2���;��Z���Cyc�-Sܐ]�hA�=�	�KgX8mظ[핸�� �l�=�+xG�:�eiN��֠B��V�RG$29b �B4Eu�@Eq��I��p$ �  �?�*�蒪&biJ�Q�E��U�mU����Ɣ#Y@��Kh�<�
h�P�-G)E�Z)���A�Z%C���%���U�U��miÆ����jVZ�Vƃ	F�x�$�L@�B��RL��L�6ť�.	�ʴs�re��9�3Q�	��1a��UH��#UƫN3(�ƤծR�E�TbI3wyKJ���mF���a��B��JP�D1dК�K��e���
Z,0���~�u�5���!eޢd�^��B�ɯy)FI�Z �9!��~�Cke~z1��>]����獏�y߿�k��+�5����n~Ԕ�=B���4?V����S�V^~<��Y[�8޺�Yq���W���G��9}�to�T��Q��t^gd���b�f��(p�±&"��ܩw������gj��P�~o����2m�����g� vp�Oz^	��-��x����֠������C4��Gʗ��T{�����z��л:���\/��}Ě���X���V����a�����9�S^�
�޾ �v�gd��ַ3"rL:�K�?�锖�r��Տ�#Qc�ꗹ	���;�+�'|�	��'OO~�ԭn�W�?~��4���7-r�������c�����)�vk}߳�)�~�uOǂ+�Y��,X�����r��_���߅~ּIY�܉�w��?����N���x�l�íԟo;�_�U4㚨J�R�[�����'��q���llw��q{qPsv��J�5ըO;�����Ro�����c*K�[����⃫/73�e��X�%k��(_���$'w���P���V#jS/f�n(B�$��w�9Ըb�4|A�Y�OAǐz|sV���M�����z�t�lQC-ޛ�uV.�O��L���yG�F��ىHJ�=�"j�;�Z&�5���S=�a�u���:Y���^)*"{^)=g��i��ŭ]�G����f`��U���=1�⥬���:T�������]ۘ:5�n�տg�<�.���x��:o;�ѣ8C)����W[��$����[����[갈��d�]�Lˏ���11~'�G�մ4�g(�c<Ġ43rv�:V'��rq<R������k#��cžKx繖��_K�B�`WTU�ww_2;�0�ows���n�
�{��B�2������N�e^�<^��੾�2%.�|�]�����jM��{�o��D�A�L�Ő��;���������]�x��� ��L��W�+�m��`���⩍��a�{!�~�]�/�Cۥ���ٛ�v*���}����
+e��F���{�XR�9%Cz¦��@���+��\�56mxx<[��mFo_7h�S#ޒ6�u��mI"$"����ʼ݂���0�'e6}��_x��Y����&����̞~(c" W�EV��3^�U���t���t���+hG�������k�?3����]�=Ͼ
b����-�^�S��f����\���b;�n{\�im����eDe_G]%����t�מ�*�ѵa�,7Wyfc
��K
����f�u�^���ӭ�K�V�����M��C�����}���(�k���@�}�eYֲ� �{yrVR�ܭ©9_��L�xO]��ǳ Β���yw�Q��i"� ���[����S3�\)��?n��X;��z���0%=)|p�>-qdx�e{=ꑝ[ji���8�Eښ��?lQg���`�^~�l�I#�gp�]WtZ!�o�;Q<þ݌�ud�wq˞����xل��B�i�on���蔊m�yT����Â���f�l[}����BT�}�әY�������Σ�;\5~�k	�	��U�v��蹍�V:��3�Y�B�"���p~��`�T�әJ]?t�o����x�/"��5ҥ\�s28䳼J*�����)��r���]�<ҵ�$��wϭ��jU:�9���<�u�ͷ�M�Co#!=ޗ�U�/���󍾿|�6��~���,yx|�Ǳ����9�w�^~:0�,w"���7O�ƚ�;����藓S��׺q�;,��j�m���\`����m{㳢�ĳ�z�$x���t(�8��q��bcǘ��%����"ʚ�{���^7���X�h�m���d����ǌ���F���\.LY�K���� ��#A5`����������d���S��qmA_���ԽP3ݽ���P&�����(&o6�r{�~�	\ކk\4�Y^>>�U��xhi.����U��^����<����w�J��<�?r�����3������;�����W�L�����eo#���ֵ3�;��{\3�!�ӝ�o�e�Q�g*Hn8�����e4�緓�;>��%�J.��b���RK˶)w�R�[5VwV�w�,d�v,����.l5��mG�;�o�ڥ���TM0���HOd:�[��FI	�IY�����%�1���x�����H�o�;�� �E�8�oIg�=�2F��+;G�{��Q�/i�N.�k/�\�ӮU]�5�ؕ��7�>�e��y+K�NYVF��L%b�:�Z��O{���L5��
��5����,���YY����o݇4�>�컯���`:G圶��u\H���]�ae�x�M��dk�� ׸��{r�b�	w}ܔ�;u-�U�!��2�֙A�~�h�{+����l͢�Za��1q��[+���s1�$��Qi� �^��s�6C`d�\;Ow��H�v�A�Q�޶������#��z������I��:�6��G3�,���^T�-�s��ֽX�Ȱ�����	���SS�y���~��%j���7�h�{��
{���8�P�=���^ԟ��ַ��j����Zȥ\Z 7����
��qsW�L4\z{��ե^g���ޛ��f#�{�������7<��2L��1&oapdӮ6���H��:JF^�iia "ܺS�u�gw��z�nf��a*anTTT�����]�B.�+��ŗ��P������T[�v�dݘv��6���{G�3��]+�P�B�����3'1������x����:p�5Z�5c�.����Z�u��0���bL,A�.�eN�kQ�Wp;�EKl�������ά��T����3kt>�mYwa���%����?o�uB���|��0Ķ::6�a��vW>�T̜m����@�R��hu��u�-ܨ�𧝕wZ,e�c-�,� +@e�����;r�΋e�hD��Y\*iV[e�2�w����&�;�`�Ld�PN�8�w���v�?����??��#d*9yz� t���mD�5�L��% ���y�X�u]����p��`�]fXj���"������Eͼ�ʯ9��3��%�@�l�*ƣV�N���Ѝ�%�v0���tU��������Z|'e�vN��� Y8�`���P�qڔ�.�����/N��N�u����j:Iμ �'��Q�E|�ܮ��b:Ov�H� ����K\WnFs!ٮ�Q��K�
��Mx�pcy�M��3�4�)H];|�U�ݒ�� �6�7��uAV���9! \xX�]�����D���@  ;����w����~b��W�:��	KQ+lo�)�0�1l��ܱ �a֣X�l&�i��QS(����`�W%%(a�p�u&%��81��k�Z[U����P&e�#!1�V�"-)�Ir�r�cTZ�	�DJ��Jµ@�A&a-HH��")�+	���dV3n`���`ū--l�cL�J�)��
a�J-���	w"k��BH��m��[���Y�Q�.�����
�x��e!��ܲ%�A�(-��6�M��������<�]���L:w�!ΆS�F+k\�,��̒_}�E&�g�~���]-����Owf�_����{���>��8��hɄ�:���[��^�����V,�Ж��إ��p.�/=�9���b(Qۑ"y18ʰ+S��N�<d��q��C��*�����M:�ͽ����x�wI��,��{�t]nW���������쭤-�!^#����׻��z�*�x;��)�ttѴ���)�c��۳��㒿���?H<�Y\�n����F��pS�d�=}�����[�K�EkZi���+\�9�uk�F�:�ۙ�?��Dv��I��q�w$Yf��74��|��3]i��E��T��}���/ܒ�q��w6C`{u�hR;�^��������D�.�NQ�5��0d1$��.W�E�8f�������w޿��W���0̮��i����Ә
�]o-A��!�<�7�f�m4�k��ާ��4b�����
o+������Y^�]�J���s՞�m�6�6����D��\<����|�ʒ��k�뾘T��n̸��d��y��`�7j7j��Df-�6�j�DDF�䔺���V}��!U�{����a�$�?j��վ��>�y$��C`�
�p��5��;�:�{_l�^�i����^O��cc�+ײ�
�yI@��]
b�5�.�@2���R)_p�|�v���e�T=�U`:�~��x%�E�Ī�C�W�m���R�n�_���<��R�]绬!�o���&��Y\[k���g�|P6LW۬��f��p�A�zԜ(,��<��"6����ee�ct����vm:�}��[�cfI?W�UT�I���N���Q���H��΍*~�F��G��>���s������㼕�����2rV��h��H������0��1�V����� ��O��fHl��2��7��{�%y3��u����eh�չw�L���V��,iPM���D����/q��}w�S����->�����g/?��K��_kU+N�]��e{�lW�=\������i�[{�@��7:���/j������;�*�+EsCdi��\&Ԉ��ʄ�U ��cnI>�_}U_4[r�wQ}�3z��(SU���2��~x�i̪�_nN�|����C
f�3��wi��`�fj�5V�B�z=�A��=}+����A׸�| �V������.z��M�-����ʷ�������䟇�� Sَ���z����q{j������*�>�ȃ���k�Ns��JqgDߍ>S6�-������Uכ�V��5��d:\��+DwB���۠�g]&9�yZ�5��{���+��K���\N'�`^2�0� ��46d���}�}E$�~M�s�ʿ~4i�(4�z���֪��j�¼�z��X~ձ���:��C�R�G��p9�-�_HhQ"��%�y�>RU̎'č�x�D}��C�;;�p�)z.U�(�H�0��z�s�y;�\������^�9u=�Qt��wq.	:�[>KO�Tf���x=��뭌6q諺��F-hD^�����&��cToʓ���O�r��(U�0̃n,���`�\��b��}Xs�u�pwlIn;o#��71c��Q53[rO�_}�}I��y�طU�9���kV�s�~�Y0f#��TEz ��j*�ָ,6s�xL���]^s:t{�I��:Ba�o����o �Ϭ�Z.�s1��.�;G���Ȫ��*�^Ռ�a��8L���e������C!�F�O�<��4�1T>�X��V�M(���R�keC�b�����w:Y9u��7��d\�f)����|�z[�tӴc�^���D�4��u���5�ȯ��,��s�*6)g"��f�1=���[�]Ӥ�6)$�_UW�Qi6��Au��W�0{!��=��	���w�
��[����>�}�g�َ�XKw��޾��;�T�r�F��H��4Ma�5��q��f�3��'~�O�v�rCP��kӼ�׷�fӺ�b����x;in�?]b��^�b//c��bc��J�*��y��֮����mo��5��;�Oy�O@ͫ��v��5>� �^^�J�ۢ�xwp�^���γF{�ub�8)�
�8��7�1��#�1��|�'"��eol�t2�0&� b&vƦ�>�8CfI?W�U}�Jo=�����o��GD�{z�|�[�������?dKz��ų���c�Oo�p��ˇ0��M�����0�+lEg����}�Ϲj�nx�����6�W~&̚�j_�mFz�����+r�-�~��[��ϫ�S^�66:��Gč}�p�<���y���*��]rP�n��\�m��C�c|��żm�u{�S�8�ή	�ͯva4�g["���s�L^Ⱝ[<q>�F�a�=�c�!M�h�2�t�}����n!h��2'$�Ͼ�������f�����C˲h<w*��c��A�����*!Q�~�����}��O�{@^��[�����_��]�c�j����z,]�o(i�L����K�ٕ�~��ۙ��C߼��1��-���,�ɚo|Y,��xܩm�K%!N-{ʐ^1L�Y	s�9ת4	��;�z���`[/��l�b�M�����'DI�za�~�b��;D^u_�G�=XG�@3��#׎��kf�������sfm�Z�gq������u5^�*h�Ҡ����uo��C6ܖ��7[Tʜ��@�|����Cb~㚦eN�]��n���د�|FVimK�]a:y��f��ӗ3;2,��p�s8��p�+�RٵՇD�ډ>.��z���⽣v﮷ZL��~N�f�¸e���2Q��4�_A�CFT
�&��%|bfU��CG&��$p����-��u�� -��5�C����+uje}0�4ʑ�f��o��iuy���8ʝ�
�ƻ*�3��a+{� ������T�ݿ�wq����k_K�u;qYSQm�o[x����L��I����T� ]0ݳ��,�~y�Y�\���T�M��I�L�YyAm���dܔ�����nն6�Q�ԕI��q�\z��U^���*�+e��&V>�Y�w[o���+�)�mP����:��9eV���b�{��w�Q�	S�j����˙Q�8�y��hs�>�)�q���l*q[6��x�s�;��ܳ���w��L$P��i�\^��E}����X��a���2��d-���)g�:X���.yau(�#�9��MCceA3��i΀+ˉp��g x�A'nU��Lk7$�Dѷ� �8� %�G#=[�D��������   ����}�=0�j��ꘪ����TJuv`ĩr	�0�L�E�Wv�����%�--��I$T�K��n���m*�%��Em���Y���ܸ�K�L1�����m9�K$��p��ӈZK�̱¡�"Iw#q#H�n.\.
��r\a#Ilq���X#Q0����࢕$K��m�i1!�(�V3qJaZ�-Qlb�p�V7c�K�j4R�T�Lah�[i,�*%JT�Vюb̛u����I�!JD[��0�$dp�a%JcPd�����`�-.B)	SB�Q�.�\�A-8o��:�'���Z�y�;���my�jw�&d��+꯾��m�y���7��������gSc�Q+?�C����ơ��縇U�7[T�ͺ�ߗn�W�.����n�ߙ���&CIVn�"u����/3��9j��W�� ���|�����z�q��7}�{�����y׽g��ws1ٮ���y|sF�lf��s�$�%��;`��3����^I���1ggGz��߮�/U7�S�-ej��ns�#S�+%B��2�[��L��ЯOb��2�X�7��Ӷ��_lX�5��O�)��핲m���r~����\�l��i�?*_�Q^9ʺ��t�ku�T���.�P���1�J6��ڸ$�R}�<z���6A|�x���$M�[]��qr���>�YQu�3�抾�z�����M?d;!��L��ּRΨ�W���2�y�_��=K�^�K�w�/eC���fQHT2���g���J�	�����m����L�W�G���r��w��l�-��S<��W�Þ/�xt�/my�k:���hi�W�
���
�^tlX����;.�V����z����׎���٠�qa�{�$���$���_U|Zm�#�����W�ڏN�a��� N c�}gb�=SE'��{P�!��Ґ�O�y;�C�v���o�Ur�����^���7�|ٖ�:s�>�<��Tzk���Mt7J3�tR�~țn	�W�e��[i�����f��0�ǻ-ʺx`�5���Sԯ[̗dW�pwR>���=��)�mj���޿W}	�������Ϧ�^�vx��<�'ȳW㬷�!�]���5]��p�W���7}��2ZME��&��B�g���C�p�y\��>�����I6>�W\�ڗ[�9n.��[���ۇ����+lb�熣h�5�\3�u�\�]8�5��֖p@��s'�'�c�1.��e�b��dn��g��[�{�����!����[��~�M����
:�i��; �W�.M}�5�GR�ڣ	[hw��w;���(�A���'P����V�Z���uT^a^h6�c�Uu���ƫ�F���{��}�~�g��A�Í����U��� �j����]��G��]j��s]��;���Q�A�.J8��+�F��>�^j�����Kk�Um� *bP
W�J�7�ɟ�Yߧ*��(j���(�q�5A�h�PC�J2ц��A�2�Zj�J��ZW��Ǿ�\����oY�f��K�����^U�U�(u
U��h�I�L�8�D([��ත���J�Sr�� p�����N�%���'���UQ\�9�s��>B��
�:j��~NJ+�_5�)h8�;*��@�J�vi�8��U�"r��E��c�k�h>h� �U9*��U��j��*�@8��h3�EN&Z��_!Ġ�aU�2щs�}�}�OUQč�Qbh�UZ�f�1�EL�U|�ģ�WZ�(�Ty1^�Too=�}�sܞ�q[iJ.��4��E�[��9UF���ƀ�U�\����hs��y޹�<
"sҪ��|�E�[B����҃4�4Q y�� �+��Uƃ[�Q���l�9�N�a!^J���iU��ZPg�Ti��]J%Q��	�*���mZ���ε�{^���������ڭ�@:��Ъ:�ƃmw
�FЬ�Z�*��(��������a+-W�5V�u�3�UG��e����T
[EM����
�T����U����w�^��}�Tpk-j���V8�u�	�J�!y�iX�����ʪ�V��W!ĠϾ�~S?]�\��m�Q�Р�E�j���*�B%�䯚�hVkR��(���.�8�=���	�9�#�es�s:��ھ]׺�U���y�Ϳn���2aU4�C�4�a����}L�ˆב����ߴ �}D}�fjIO�#������?
Qx�Yj��h0њJ�k���U��U3
!s몢�*��q��޻�k7����|�J>��G�ƈ�CmPk�@�ҸզL�-(F�#A� Zv�B�7*�զP#X3Ma(R�k���{��s�1;��P�yX�戔/۔�ֈ�>J���D:���A�!��6�)�֚���)O D�Fs+	B�)��i��f>~��5�����H�戔)��l�U��P�Uְ�-b�
[j�����
WS�a<��5��-(P�aVѴ2�VO�ZP�iw���|�\�P�"y�[��!�*%�U���)FwvP�
^O]W�Q��ƈ�u�;h#8��A��4q-2���5ۜ���~εͽZ�U�Q���iB�i��UiB�--R� F�mD�U�҅(Q�X�-ܢ�4��Q0��u���QiB5�w��w�g>��A���G�
$h4��z����Z�-X�ֈ�d�-h��0���mD5�*҅�ZP�������8�o~Ϟ�(Z�U�@-2��zk)B�cҭ6�gТ ZF�5Q(S-]5�a��QF��P�cT����%
V���q׻��}�e6���ͥy�/�P-C����-MWea(S(\��Q�A�(s(�p�(�\(R�ᦫn��k�Ϸ���w�Xh>bW�F��@�iB�/�ҫ��e!�������J
P�촡J�} ���L�;
�UƢi%
Q߱�����_��o�%��o�����v��^`X�I�1\�\-]�v�
���=�K�[Ҥ�F�on7N��*��'tfR���r+꯫�Is��e�X�)�@�᠍4D�v��5�e(R��,�h8ƴ�v�B��@��LN�d�j��JQhD�B�(ӆ�4D�������ﵝzt<�-h�#U��J�B��Q4u��eZP���7
�M�Q���-�Qi����8J��QiB�{���俷�s<����j�j%(-V��ݖ�u�R�᠉B��"e5XܫJ������a��%F�v��P�Z2}+W��Z	�����5�ޔu(nW���(Z>��؅
R'��6�F��A�5��4bU��҅(P:�-8�V��UƢ>�ZP�Z�߭���'�J��-(ZZ�3��j�j'��eJ�-D�T�(rz�-�A�����Rq�%
P�B�q��(Z�}Ɖ�����j���O�P�V��e�a�/6�G�J�B���V����͡Ĩ�)�0Cmm�?J-(Z�F��N�C�>���2��P�Ѫ�����m(P3R�B�-�)^L5[j!��|�J��u�R��iB�)g�6��5�+�F������=޵}��FZ0��P�
F��iB� F�l�J��u�iy�g��>��v7�޹��ۦ�6��&�æ>�3��x���<I�kͬ繂�*&R�0��)o��έb�M���U����ȹ�([�IC}%��`�ýD<���h��Rlj����z��J�b�Ӟ��H�K�?�}GŦ۽���W1��*Ǳp�`ګ��>���U��vl &Ag��A� ۽}���eh�d��|:��&T^�x��7�AxR��*_�{��]u/鳪f{ύ���S��vz͹�,�[毮��D����Vڠ��6�邦k)�Ϩ��ۤC�j��~����œ~� �k�ze�l_<�m�x��3�:�{�{�m;��rw��)���f$'��)�N8c�����]������X�����5���ۥ�p�;۲���R1��\C�Z�b��os�F����ן����_��Sݛ�S�M��oF,��Ͷ��ܚn9̯[���Q+�ud�#d/a\�OBҡ�mn�!+e룕}G"�T�7�Aa��75�$��fI?}��_|���ɞ��/�=�.����K!�۞z��LX�ku�&Y�~�Y&+Yy�X�
���iɢu3�=5�w>l���;r������p�ͺE�"�`w�>��{��|}g������9�3I��	�Lz��f&a�Eߴ;�\�n��;��w���k}��]W]j��׳}	��R����Q�/n�)<��_W�;|��}	��'�.]U�];;���}�V��1�}Kz�N	�w:���vs�M�0�<:Y�S��|w��I��K�I�DǕ\��)�5���e;��qp��:�i�^��^��h��^T
�ͽ�(��u��B�/�L{[�+=Ch9׃U�WP����/i�U2��%��s��]�lE�4��V9Q,�Lܚ�ú�J�w	���>�#��䒊r�?|�Ӓ�0��]K�٘�]���D�䇼��b�{=0��[�3�m��uc(���]n�g�/x��j��|lZ�}��_^[�Ja���:z�N�+�>7Y}j��@@)�x+(e�
�{j����B߅u���R�u/-[��7w\EY��"d��
����A���>�vP�V�`���f2�-���/d�m�����=7�c�Mu��ds��/�绗H�r���65��弗/B�vp.�u;u<u�S�^U׀i1������t�$��N9Ƿ��ގ��_4i��z�Bi��r%m��ߦ�յ�oGR�9C�η�k� w��)�3Yք��t��1v7oe�B�Zr�tfJ{w|C�(c�f������fZ�N3Fn�`��Y=�љ�A0�^�b�۫BB2+cBykM���>'l_Wj�'�}���K��a�>ݰjq[�K�R&�v򺵯 8V�<��u�jY�=�%o@����cO�".�h|��
t�5�3�5%���*v;z8�Y���w2�}wO�z[���v�W]d�S�w\0��9�'�27��
�K8jV��Y]Q���>�|J�	��ʸ`�JCV��;+^�+g��k�YFV�h��7}�#��'�t�e&������[��E�4`g�*n�p�#GiӜ�6�mjr�-���]/,s�\-�h˂K�X/p�G]vʒ��|��X�6���=�%�c�'h\�ٕ���q:aJ])��oPݚ��ER��vU�{j��[9\��Kd�J�Yݝ4U��&���ᜠ�1N����uc5-F�	�L&>5�9Y�сSG{8Xeu��Ֆ���m4���lj�����[�:��P�jrO�֙��e�F�܎����.Nv2�ݞ�� Μoj�e�.��ھ�{�]�'�]����\���H��Tw`���x�tʀ�����GK��\nM�L�� ���s� �D �GBι]\u�N�ҳ�    �}�a�w���4�-��Jb'��\X�B[�,�D���Y#��\AV$I"IYJ&n$�M�#3%��p�1�EBS)�-��e)��Kj"�*F��5m[��B�&!-���0�%U�i1Yw˻�m1�*�&��M�čbH*5����Knp��jK�%�QKY	��X1�Qi�мB6�T�Ҫ�Q��.$���m�*Z�QU�.T��mZp*�4��
"-a���42۶��Z��0����۬%[XE����*ڗ(f�&��&��d�
�?L�s5�D��-��Q�#���ho���DD}��%3�!�Yu����3!��e��q�sz���'�ͥ�q0�~�m�1�cwzO&5+�T�e��Ƨ��D�kf!Ud�uE�d�e�̯_����ⷀ��z��L}��j��8���VzV/��8�N����w'A��o��W�om@n�����������~޾�3r=oЃ�%��i�sX<��������Jpw�w�:���6�ZYPӘ�W5���Ƶ���vT��b���.���+��ؾ�qZK� �d�^��P
����|��<6�r���]�^�ؘu>�V������`���ݷ��u��?�uP�׺����׺8����e�G�\�u��|�(�W���"�k�3L��؊s���j"5kem:���a2�֖�/�Dr�@�������j���6�ߘw������f���{�d�X�~�N�n��]������>�ƌ���_/!�̸�/Κ�Fq4ǝ�}Z��3<w�Q����~gi���u�m��ɩ�K�0���u��=}/fhv�J�����h�}eP���lV��̣�x��ݻ�}���#o�엷Y(y�{�%�Tܬ��R��7�)����WǅW]{�x���a�j�ݎϥ_��ktQ���3��ۃ�J:$���DU���2�w��]�۳t��
�)�Z�/�
����ec��(�Z�]�x)_X9^���Ի��Ky^��v!���fȃA�9ХYaU�E�zfW8��3��l���q��ͮ�y��j ����ѫ�AF�?~�1q�nk��hj�|6��]+��K��9����f__l���Z��{�M��1d6&5���0�z�>����ۗ�[�| �>xo��Ԟ����xR�E�l����t�!"��g�X"���ۿ���V�Y�����yj�����9�i��[�$��vi�pÇoN�U�vg�7vK���+�����LUH2���Ee�w���{���wf�+��A��J���]k��޾�r��xBB�]�[���"��U��\7A�1C�^�\��jtzðַjo���<�8�s6._��ys�����)X9iԆ�t�����g:܃��v:J������[=��Y��]�����Fh�$�Y�O�}�W�$���W���[�_ݶ>����aS<{c�#;��Ưv��vVTCl,Z�_������4��n��Y"m�7�#��o�/~"���
7�z�:s�c�Զn_]�V��଱���/m].�tSڏg9�P�j�����N>M���v�уy�{~����w3��k%�7�]{3��d-�a��w�45���S.��E|�ɹ�~w�z�ev)L�g�
�z��xP���],+�"��N��^�r�w�2�����0u�{$��;ɇH����g3Lw�{�= U/�!ڹ��xed
�vP:>˗��*{�/�c9�� ����-\8�4�]
/�vE���>�a\�[p�K����wK�:�ۙ�G'ꯪ�I���������w_���+`S�mAB�^/��1�y����E��ϰ��۾'{�>�9:��7f�L�sA�~�*\�M
�`�o�ݫ��.�oy����o��O�Z�4�Ұ�M>vV*�fw�y�OOJ��:��/���cܯ��+3����>e�^���v/j
��7^����~�>��"k��ݛC�e7�Y�;}p�p̂���~\���K���B�+h���1]y��8o^ǹ9N>�y��u�Ӽ�͹y��|�%�7�mS�}zx�̎�6(U�2�P�F��kk`6�y���y� �}�#���eM�
�7,�G�(
���������u�����S��ջx�tt�@�5;����·��6$�}��E��NF��w�|��&�;k	���3�mA[Y]��'qVO�om�MyI������1ә_)��u�=��J�9�%�C��#�o��}�0M˒}�ǳ�nUO,�X�xr��8��O15��ۿN&�5�cY��i㣵��NQ�yGE
���v;��^�(�����X�mǎ�n�|���7�^�]���Lk<vG��p����K7�V��4��Pͧ�C:ߤ#ְ�^s�y���;r�8|�s�F����z�^"�x�B����|�{7�qӱ�M�g�y����3���T4=n��b��o��Pa�ze{�^ҳH�w�"�Yux;3��Lqw��B�a]�ofJ��P��p����8�7:٫E�1䠤8ْO��URl]~��(V�߿b̤�)Y��P��{�g���e�z�*z��G#]�6�>�vT9��;�;�cZ���sח�r�qr���/�!��R��{��;��Q��q̩d�b��ں�[�����b�m�SVQ�u�;�����u#��R!�u W�B��Y^�t����X��j��l&��\]��cy�Y�g���C�V�>�`�C��F�S�c~�/>�ELрV���t@�����'R'Yu��<��z׋�u���ӄO]כv�d��!�3�H[�^����=����@l]e����wYu�w	1u�u�f����i,�}�_z=.q`���/�e���[�I�&"Ef&��_Bz�D�q���$K:�U;�i ��Dn. �.\I?�B��
yC�,5��&m���VZ|�]���$|H�f��ŪS3�*q�$\GL(�2{)J���^}$[^�^]e_L8(g��\���c�-�o�:��yj�R���_��m_��YwJ
oq_���#ݛ�GއSO�6��3�U�g�ܗ�Ia�*f�q�=��{u�%��B�__�쎿^_�GS�r�[�0��9
�y��n��u���^2��)嶽^�~��&�ߐ��
�}^Hߠ�ˢ䥎Ogw�wx��x��M��/.Ӊo&���a�1q���
�];Lm�,ޱ�Эں��[|�3v��6ku'j톘B
[aϕ���([�R�U]���8�
�v�{�k[]I))JC�{f�;��r+����@?}F�I)����jr~�$(U�Î��>Ò�yl�P7�.S[u��<��YzB�"��;���S��7�-t�ML{:�K�*���צ-����j�׵���{{����D>�=~�t�Y�*��C/�V\���%%��b^V�Hb�O%�q}6�CG���Ko��1���*�"��;�i;�h�*z���J<w���{��B�>,!��Ю��*{v�z�Ǭ�g>㥏S����ɦ�?e�l߼>�WBlǅ��>���������3ٗ�̆8L��5o��{zۋ�T�Pb�ז���@ؼ�2�¸~��n��wW��;�̈́�@!bV�+X��k�.��SHGi���N�nMu�����G eզ�6q�NI'��&�}�F��TE���t��`7M��엷�W^K�q���.�*j
�ͯ�w�[D�v+�iס�����ˏAz$|�����I�y嗹�����i�Աt��wZ@�y���ˮ��6Y�`����<o���Hl2�];ǒ�ʺ���y���p�)wOw	y~b�s�lWW�B�콵}t��>y�Gq��b��5�l�7��z�ؓ����P*�*ϩ_��u�2�^pˬg��T�ˋ����0f�)]zψ��������U��<��h������
�w	de~z�ۼ$}�ކ�_���_��{kN�t�)\��j����}���U�z"� ��.�m�,2���Ќ��]+
6��N���*8�*-=ש�u�r���)��oV3t�m`��\*;t+s9؉�]��m��e 9�Z��!%�u��[!j[�9_��Jƍ�8+�r�NXT[�,,n���mN��B�J9x-�$.A�.�O;R׵zH�N���X�qrrm�̗W��u쥗D;�E��3fWf�0�̀U��֋��5ľ�����X�J�W%Lvq�2��/"ڈ]�4[Ttkٗw�5�S>��r����05�:�4{.�'aU���l�Vq8N�u7B����*r�����y{v�T��9�����L���{��߶+�6�ZQO]׭b��U
:���c�92�3e�ul�x)WH�fL<��S�KGt�/`"�_BFd�#Y�r��E3������3��v�2-,�h���K���ۡMk�s$p]
�X�y&W"���']B�e�[z�o2���2Z�jnϖ$�;����KF`����8�:f�u���x�+tѰHwt�����; *e�=8���s��pܡ7pZ����:�"zR�_I֛ɚ2;*\;���H��y�<�����έ�cϯ��+|���ޭ�E�I��� ���{����5W�3�t޾��  h꿾��ө���ŸH�D�FIm,j#W��Z��M�1��(-
�DU(Z}���Z0�e��H��E�H�$��1��U"fB��!2�s -��
�H
)lG\�!����T�����B�*�479�+SZ�.31d1�QTt�UQiL%J#��1p�[KM\#Jx�ҍ:b�i,K$]B&_���cw��n�;]憰ur�p��q<�D��� ����w%jR���uT������u��%�ںWB��6,�aw�-mO	Wmy������\�L<�6�.�޲ov��.\:�N�iӞ�e)���ӵ�Uu��e���ҾaY���n��+��o�vo�~k�{/}3낝��hy�u�
V�<6�5����<'���;LF&�۞��zT��r��׵wK���+�&�&6}u�L�eq0��
��ַ�S��̢cgN�ڨ�	�Q�WU�~��[�ϸ���\��I�Zú��)�!�����W��z����ө�M�e��<M����nW8�����uy+��,z�F�J֯j���'\�L��ްƹҲ��]�q�*g-�������fI?}�}E�[t�P����Ê����X�zGY5�畅eu~�����r��>wR�e�^�S�nG@��}��f�|)\��6�:���
}f�Xr{���l�����&&fW����X+om_1�a�W�z�\t�!R�>������a�=��a��3�x����H��]�S����r�BE��1J+=Yu�J�`Z�vq�����Yz��ҍ�{Ⱥ�.��7g1�{z��t�zKkژO>Mc[�Yˮ����Y��̗/j������˩���X*���{���م7v=�{p^޵�O7�G�_5c�r��鋞�9��7�JpҜ��x�{H5�H\TK��s6����1uu	%0d#7:3)��Qϡ�RHvd���;�{�.� 
�b9O��>�O���b�Kp_����8.�����+�g�-_�7F�n`��z���o�G��
�5�~gFH�V��v��u.��j�t4;ʨ>W�Z����z�|Lxz�}Ɇ��Y�s8�G9�qמ�w�2�Ҷ�}���f�.M;Ϯ�"�5����ѵu�J�u�W��>�mY�O.\��sx������þ�8�s����
T����U���~*�J�oD�f�w0�J�k��箋���Ǧ�N:ܶ��w�,s^ǜ1���8����c��خ����J�̡ࠫ��X��:������}�o.�������m]W��������ɂ�s�3Zp\��1��iĪm\
�xJ�;�;�=��u�B���UG}�)X�d�G[�����IJ�s.��F��g��d�/6�^���E�Ʊ��_�vlikP�}~�u˓/��2�ʿ���^Z@��b�1��r�]]�_���i�y/�_��,U$<�����R��i����_��G���q mԺ|>>r_0������Y��gOx�pg�ϳ��K5�,&*��Z毨a8��q�u�j�6ㄭq6�fo��_1��6���y�����u�6�]a\�k��1+8��������y��z���IHe��ܿ�_��lS�p赢A�v�ws��P���z���s����N�-[������wҕ̗x �Y��lX��(�n	��jCy�O>{��D�ռ1G`N��J�m��k4��x��:R���r~��E7����/a�tX��۟�e�t=����<�gzl|#����k[�f[̴��E�~�ߦ4N�;�|�';7�ְ�u�YnjV���ӏN8�[�w{״�N����M1.�((ٱ������ ����[t���;��a7u�-�u˱6��9�&���\o�{�x��؇YȻ�,�epr�L<v�9}���KH��jV{zu�{��t9e�.��3x<<�w���~�{DU=n��b�����vM��b������,�9z�Φd3�a׷uf�sn7�:�u�8o���lt��G#)�{*Y^�C�/{�1�y�xib�Er�ϯ���lU����3rN	�(Nk���WMR1&���3RI�猪�c>���]+���߬[�7�U�.����3,[Vvb]�>��C\"ùN�2��t+��5Z)ت�S>�/`q���eψm�f!3���/s�笇'70n�|���շS����y�(��ea���ӽ�'a����7�ޕ���J3g=u�xP��V�pe�d}S�e���)vW<�{�e�4���Xk3��;��9�|ŝ�ݞx�.a�g���16���d������Lʗ�wm�Uɫ�;x��c��7��kI�����;������z�L��C|�Vؾ�_8g5ug&ճd���y�U��N2:������u��Ш�y��Y��ϓy�@�,�����Y���roPN�J8ۙfT�pL�'�����m�dCɇm)�|��5�M�]z�'-v��q�؟����zmm����2��}/�(��qΡ.GYw%���ه0�2�lWI��>�̚��j�����S+�"���o�W�Q��3�r/"E�[��o���ٷn��m1�oR=�CY��������W�W��:Ż�z2���������!˻;7�{�f_&gmc���[tjͻ���W��c��Ԯ�V�\�ޱT������1U��w��d�wwW2��h�[�TĴs��*��w��Z�A�\�b��t5eeG�^��6����ǩ��?e�"1zľ�5�<*��^��0U���0���붮	����M�؟.��;7�VR�q��7�z� �gn�Js�?��d��ja��\���u�Ю�v���TIiyf��ٻ����
勥�?;(xõ���k��{.�N^!us7HkD�W��������;��35vk��08r��u���u
&!��
e,[7매�Wrkef�lm=&�ǥN��y�y��=���p��^<k�yq�i�q��4lߜ�D6��fN>v꺯�p��6�^��T�5\{$�&c!�[X��i�ry�g�Z{������d�^��!s�Az�J-ݓrL9������q�LB������s���#}����.c�.��u�h����W�U3m�/��v�5��b}"�R��4X+ijYs3QW���過�� �7
{sx�v�2�������ޔ�μ�mHwR�O�Sn����j��Ӕá"u�����I�{�m����]ל=��v�&32�7܎��rc�-�{-��]&J����F�;��t��_��������"��o�+Nm��AZ|:͝��KO�tP�gL��^ھ�
�P�|*���%���Y�]R��em���z�6��p�����K��Yn�ZX.��ۣC*���SW�;^�ԼMru�'��Ԭ�kf�g���7�o�6���(Y�__zm�w���5q[7����eg�7*Ȃa��S;�*T�;��2Y���>���*z}�v/�aףG^+��/��p�j�0���#�h��=��_e���ħJݹ��<�o^mmur�[xt̆�'ݨ����˷\U�;�q�H�'ꢉM�_�_�ۿ��]��c�u ��yW�SxE�yr;{^%I*�<��M�CO^;�on
o��{�x�wT�졟{����qٕ�Vߐ�k���L�Je��G����2�����U�x�T��6�a$�g����sW���a�����i�@sfy��	�خ%zt���_�
^98ko�W�^��=�}r�z��R"��w��w��W.ϝ��!�s(|�A]�����ɜ�nBzrռo0�|�^&�\ӽM�x��9u=��L����YF��ĺ>�ʳr呂��W���^�����ܪ��0o�ZER�)[��V��� K��v{�����B냛 Uû�mأ)�.�g�6misKlP�f����Z,q�]��6M���pK��V��5H�)�e��ˋH��H�E������S����1UnRU�� ��a}jG3��6���͎�|�"���3G1}�;�T�;z6�dP����b�{Eu�9��r���q�ژ[���Ǆ�j�	�-y�e]a��Wt>��;o�� w
'�)
��I{�6I}��EX��P�Gn�-�o
=|s��.L^p\s%B�;�hM\���ח*2�.w�|	����ݦ�U�V��N�;���i�*i�ԍ�^�_گ:��� #"�B&+�s,P�����9�_lM5�@��SP	���Gn���q��m����椒����_s5(�V4��8�E������:��镭��ҕ�R��1	v�py.��K�&�#1�������g����_�����|��M�u�]'�̋I��RZ���g5���O.=�W%.ƞ����r�3;v��7d�H���cѕ�)I;�a�c�-�K7[�2�J`!�b�����Nk԰�O�Z��r��L�O�ǩ�zX�+qJG�;in�]{��F�]B�Y=WH�A� *�h���+�/�z����   �  4���S115?DTL�M(���e'#K���JnEhW,-��*I1"��	�lV��
���Nf�!�F�1T1%*6Ɩ��Tn�0��Z�]�a�"Ҫдካ$�"ZDZW1r�p��p1q"����%�ڻF��˄��D�U2��,�Dh�V"J#H����ih�UkDF5��X�(��U�UQ��H*(��[�ZE��ImB�UEQbf��J��T���H�U"���h��Tf�t�͙�[�L6�� �9dmf�����#RI=��}1�[�+Eh����6��j�|W^�|����e��{�[�O:k|�Cڇ94�-�Ksz��6��}�+����������\k��L�k��0s�Ě�u~�B<|�j����]��˥�s��g�Sc��|%�wB� �We�P�'�vx$zŞ���805����=Դ��ַk\����^���4�mҺV�hW��UJ�����}ï@=�/^��Uer	�J��Ϛ�'[�"a�]��L{���{��t��ſzՔ��!]�6�t/H�U'b~冽���\=����y଱����?�J��Ifi��� �,�Gn<�r���J�[�9v�Ż�X�N����#�]��u�X�sq`I4!�����R�
����W^]8.��]M̧�=�v��C��������{�+�b� w�EU�W���n+�v���S��{��`�_]^|�{�bZ9��
ˮ�Z��emG�,��}��{A�!Yd�ul�Ǻ���&.rvrbҼʽc�����ۯKbs��+����m�{��'��h-��i����5�v����������Wz�a��-=C��8�;!��	Kw}�V���k:aW�����Q�����p崌�<��=�[��Ƴ�w����9zv�n�:�����n�ם���v��׳�=�N�׎ޫ�ܕ�̹M�m��o^��G3�T�26󘗈�z+�I���5Nu���I�ɜ��(=_ö�u��ݙ����N��(�Q��1�=
0I�?����+�n��K�����6���b�y��r��Qň��;�7�t��o~�M�C�y��v������'��fP��P�/n����D��b�����1Y�;��Z���˭�ۙ��5�ڈ�e�oѕ��e��jb9��Y�ۜA�BD���;���3��^�98[�J㇞;{iK�o)�p����>��/x�;������oP��]ÿ��w���M������Z�c6�cE/C�}*ay_˪��fU�j�w|+��]�*����1E�
�B�t�V�� �L>�ιܣn�(�C�L�W�^����y^Z�����*�����%������uq��,��)Rj�Ҁ{.��nk�S��_3�C��~�[m١��e���(z�ޡN�M����>����`=�D+����]]�g����r�e�]t���"�oX�� �{q�}<x�n��2�Ӯ]#��k~���	�����Z�WU�]�Ok���Z���;���A]]���y��v ��*A�uH<����ս�B*Y��%BB�i<�۳P&��8�onw=��g)r���7��Y>\Ͻ'���+{~�)����d��u�m��_����çɇ"�����}�2��}�ms3���\�y�m��\1o7{�2��7�s�+�wK�_�EyQ�p�(�E��F]g�8֊wW�7� ��`�Dj��f��ZE��(����_h�2�fQ�ӛR��Dʹ���W�z���yGIp�HG�ݦm��U��6d��E&ÿ�Uv������t��`�u�;S�Gd;��\�'�bzBzs-a�i�r��%�U�C�=��dY�]zW�}�KG�}YA�u�f���,���x����c��Tf]���~�*��Ǖi˺'�-k�ӕ�hw���y^��u��-v@�/3�����*vz]]����sb9R����9ɴ�m�d�w�:p��+��B��N��󿙫�tG�w��>
����b�.m�-��J�t=|��szƺ�W��8L�`�2饩���z��]T��쳧Ȅ�|.���nW��wkF]�}�����E�]���u�杈�48���N#�#ܤWk�bsh+�|ڻײb8�q���wUf�]��?F�H�O����^ө�\�Ǽ�{:�i�o�����S��|\g�J��MI$��,o���6z��_q�b��ɇ(c]��N��lǺ�QQs��o��xĪ��\Ø������];��NQ�em���H9sV�3���Y�Si�	��&>&{�w��žkMa��^&��&�y1�R��Y��F��
�W��[zN}�7d+3>�.���::�XW���=~�˗Fd��X`��*�t,��Z��{�u'��}r�+.�9�/.�.��9�qYs{��z�{��y��^m�'.�IPĦ<%푕�}*�!���F�e��SzwRk}{G�4z�Yh�x�X�+ސ]t�ycM�S�.��H)�X�E;�8'�޿)��m�(�&��_�χ����a����ʌ�wO�T��B{x�vR�qvq��ˤ�J�-,G޼�s�kr��k��t���'.��Mby�d��[����٦�x�w���weߐ��]��>��w뭽���xu�$��ۂ؃�"~�'f�s�L���+$��9��uG�R:O'�I�=��M5����l�wƳ���.E�G{��<�jڿB�r�����$����;�6�L����|�]��^{%��Wp�"��x����TV������o�WU�V�˯��.�j���
w���ɗ���1���a\�L��}�s��w ��J��{eu�z�~N�2�{��ݵ�x�[J�&�����0�����#�#M�m�w(���q�2I'��&�o����
w����_��C�]j8�};w/���c|��G���W�z��{%�k��آ����/���.��\>���=~�(|@�D+[�ۤ^�����|'�C-�u��ܯ\oWNs7=ީ�7/����	Wכp,^.��3���m#�_��m�˄�)�4���70�B�h��U�y3���N���e�>ܦc�B�los���%�Дw�����<����\)���b[�
:����9�Nn�C�	���:5�t'���%�xw�,�u�Y&�� w
�q]]��Q��uZ�YXy��XƸ�^�g����$8b�O�|ZI�ŵr�_W��7c+b���v�*h��\?�8�GL߼�kw�ʛ�4��o�i���z���^��y��hx�ޤ�ѥ���G�R��`�'�L#k��h-{u;�W�Q���]�����Z�^��~w�fo������o�b����A�k��=��G��'��=�a�Q����0�_m��/XZ�u���j=~ֽ������Ǧ���^����^!��Szq�7�"iߚ(���e�7��=�]��4�gS���qe�J�y�(�Ve�p\M�ا.���s�WIL�'�)60~���ki�k��^*�Ohy�/�������ʻʞ>T�)���5�����3�������c\�\��+آ�>qk��Hn���_���ޭ9��ց<FI+�5/[��=��ͮ�I{<��9��}��>�?y��Wr�Z��^�i�ܻ���lSQq5�7Sﺭ�F���N贚U�}��)8_�˷wV����
k�{AG����g�?���0U�v����if���\�kuyʂVe�s���xhҗ�F��s2p�\�]K�Z��� 
�J G���!��:�_%͵/r���P�`��Qf������B��:�AݞU�:Z��B Y��̩[ˍ�p�8[��y�.�mBp�\[[��Rۮ�4^Yz*E���8��H����w>wi ���v�@ԥ�
]�{���6�����{��q�Y�����v\"�%��,k���)�zPv����޾��w-��P.������R�:*V�8%J�gumt{�ze�1���2ԹH�C�z�"���ƃ��f�T�O,V�6�J�������40�-�a���7X��"Xi����em���:�mC}�u�m�g���Z�8��<��r���N�|-��C��Cz�x�wuuc����ً��k%Yq��V$*��a���)��mL@��Mwo*"Hck9@.nd���5�8t���jF^�����{�s3�I[ᳶj��"Հ'Wԋl�C�x`Q�<*�F��Pf_B�:��N%���g�&I)�t��b��f�M4��l��Pwǐ��նX�f�;Mq��H^pf��\�>��=�P`�+�/�ݧX��K��2�)K���.B����rA�  T$����I�x��H��@�   �{���~�ȏ�Ay�J��H*"�-=�Z�V�T�\@�R��"��Z�-��4��YJ* �4(�"-4��4�B"�"4�"�(�bvJZE@F�Z�UU�h��-*��:���QJZQ��iU���E�iD[b*.X���*��Mz˹DSR ���� �e%�BP�i�UUPTF����5$UQ��Q�(ċ$d�����Y"12ڊ�7*����H�I*4b�"[��&eD����H�F�.f�ⴢ�D�#W#lXл���n:�g��ϘDŲ�X�.�zh��{.�@�#�O��`���V��N��
C}���U�h�(��K�0=������t�Zc�4�o];���z@�r)�k�Zh�&¿Be'{L�W������h��^R��`G�c��[��|2���{�gB�S�oJ>��Ν0�)=���A��B�ԴHG�k�U��j5�{y�3Cݽ=JTB��Ux�oź��ٞ׳�kt�31|�%����{��zU��oz\-�\r����J6v)qO6��n��(�u7�j�V_jWr�'w\�5�܈Ku�2�b6�6�o�(d��}UI&��޿�叺��z�o��>���K��Za:���w�+���?y.}C�b��>x�z�1/�j���5�&FM�i�,K^/v-��}��vTN�;��#��3Dה5�ᕫ(9~R9+Y�+އ}��k�,�.��!b���0���*�C������JK�|��b����d�]"���a�S��!�c'���
J{���ּ���&c�%>q-WPy< x��V��7�Ҭ��.��c��Îy�ʰ���e�*��,#[�mIrT�z�t�m�z�]�:&<ĶJ�☚�O�U��"�o���/#���י�Ŗ�6�y�Y��q��{z[}(��O�;1*�Gy�����s��K�ϻf%����#���~9ʥ�Jq�N���s6Sooi+�JUΣ6��]�Q�_�����;�gOO������}7�On�����N'���:y�i�o�N?>Qh[�I^]��{��淳^�5��/���;sI����á6�o�����^�PYB�Ӻ��/��[���lcrw���W{E���<��A�Lfݲ�N�zHJ��s1�$�ϫ�����c�~�C�h~43�R	C�J�d��?^�L�i~���=SJҲ�P�K�_�����G5�bG[Y��B=�Rg�odɧ�{�eG0'w�zsi.M�Kd�:˲i�S�&9�:���o�� �#+y�v��.ȹ�\1�t�Gz]���o��k\�h��އ���ç���.^��ώ�B�\5P�)ޞ��C<�z8��F-ݓ�f����sq�Ä85xp��.�O|e��Yg`�	YH����E��*�ecf�����RI�3$��ﾯ�)63��﹍ֳ�0ˡ�+�.9��ǚ.��(O��<�ҽ�+y=K�0pg����z�����-üV��peu{�#�S�>��?Kͬ�y%=}��ܸ�	)��lvx���g;g�e$5%��h�{r݇�λ�����^�r.I��_��s0�WM)�/�h�Ow��-�]�֖q�>x3; �y}w�o7jz���I��;���V�`��B��~�؉8�T��l��]K��snd�X��Ŷ
��ig�N�.�;�N*rM�oE8�t͡R��J������'ꪥͶ��G�:�K���|�u�^�8�:ZV>�yR�[�뛯L��KY�]��ޫ�E�'De>��Ň���vH{�ͽK�.[~��\�s!��<��g]�=7~�.��b�WO��<������˝�[��q�w�	󛎽���&�'�|���x/W5c�(u����������w��Ѯꔜn���w���oih����yZ�>O3= Uj��0�ٽ�S�b�x������[E��[���ݏ��4��'x�bh �;:��R�;��!�1�?}�wwn��ߵ�A����!�G��ۇ�*�ם�啂�J��{��s�!�+4��A�h�v�1�
��O=y;��l����Y�����V[O)SN��vY���6qמ�U��xУO�fsզ�|��{�����<�_�l�buyjT�o��m����F�y]������;�vJ̞��k�����uŋ�"�I{�|�ug��y̯i�[}}w֑ؕrV̈P[���5�SWE���9ҕ��9%H�]��!��9�a��$���I���f��>is��K%���"�/;W=������q�>N�
�8�����7�ի:=�LwX0SAg���ҋ={�X3(7r��! �k�����-�QL��V�
�'Z�޼�z��>��rP5�G�Ħz�b|��Rg�W��_	E�i�=�eL`���ܗ�b��~[��&��֫��sru;�������7GU׽��#�a\kGxZ�w�(*1-�����v��V;��܂{]�P�������U;m��2�\A鼌�H�I ~�"#W$����Ɋo�'����d{��Z�^�!�Q4��!_���+G9�Fo��@|��@�m	C��*/u��k����J;�ol�c({�y1w�x�ރw�"L 賞7`����n@��W����~����W6�t{ʼY�(�=�K��)�v��1i
�EX����v�)�,u�%+�>p��>�����:�*L2Ot�ܮ�Yh/sWb�K��{5v�2�ڲKu͵3iҖ�I�R��[��j�V���t7�ԝ�x��m�ř#Й�O�U�$Rl^��߮���}�4޽k����㣞�������x��oZ��>��/6�u���o�\c�y�,��'�"�&�`η�]�nF�m��u�[B��>ެ�W0�^�zb��t��T��wlwO�k��Sޫ��-�u��Ղ�g3��=���<���(���ZQ�M[�w�S���|�r)&4����Vp^�C��z��WPв����W�%PG�r< �D V��tB��֩,:8Q���h:9�.����i�d��v�B.�Ѣy�W-��fX������#v^A�[ݵ7���HZ����U�K��X���筱c�q�=�%Sd[�3B�މ�^�*�$��Y3:,��˟D�����zr�ͽ�r�=����+q��ʄ���»w(�t(�䋐�j{K0C[�f�Q�Q�m:�@��mޗ���2�j"t*�z�����R��K�0ۥ����,A�8������+Mb���:����jOi��ʅ�\��F�/��v�(�V.|�Qe鶌�ʐb�Q6x[]��=	��I\�9c=��X�4�vE�Q��fK�h�%��a��.��!�}��rɔ�� u�����7��:掚�Κ�r���v��pQ`K�n���}��X�jąN-�:S]��9^��krR�B��KN�7�R���l	��q�9]P��m�=�-Je(,� �0a�7�M�2u�ӏ�;��"m���*�@F��%�uNn��|��q���_����L��R��R���v���_Vw��>OY���,V��0�4z�L��Y+֠.L���*j�}�&��X�A�稢��� �4@ �K�A�u����H��p � @  �n�333>���J�2��",����Z���ƒ�M)%BEd�GHKŮq��.DÅ�R�X�܎�*�!QF�V�H�KX����QR����"B�(�"���"li���60�.�QP�`��+.�PUUQEj�ĒAD��iiV����B*a��"�r
)KH��Ui1
��DAU�JTT̔���TF�ب*�VA�DnF���,<n��L�3b��T��6k��S��F	"�!��#���I6!Fִ���l	@�79
��T1*�WȒ��=�}G�����{C��ݹwY�y�s,�R�L���}}oi4:���I����S4;��
�9�rn?3�ߏ�߰Ћ����XOn��w%?QU����j���]�d̷�z[��k�������dv���1�{$F�y:�-�t�{�DYQ7�ѭ�{<h�`;�z;�o� P�����X��Eۇϭ�{#��8��O������/6�a�:����a���䟪����w~I�9�W���s+��
���vV��B5J�k���>��d��R]�P�WM�qֽ�^v-�a�V�a�Ν�i7
����]�~+|=g��}�L�����֖�ĝ5��;sqW�&L�(�L\���,����}O�۶�90�z����4׃�u��H�9��+�eߍD���*.�c�����:}��[s}g���d\�/�d��k�͠�V'N��>o�
�|�q�4X��w�_H�Q�靬��#�\i8�1ʷ"�̒>��"Su��O��8�Pkj:`�oz@��OgS;��w��F{��e�	�~��Ψǐ��p��(٨���<��z��SRV�Y7J�~�V�a4Gg#΁��y�KPQQ�p�*��d{p����^b'΋�Ӧ�[^'�v:��&_W��v1\w:QN1H��,]�2[��˅�����y�5����{:!�b�����6u�7ҷ�⽁8.;O�G-�1-m��\�����l��C �[�H��x��o����&s0�.�Otɦ>p��-, �s1��>�w$5_��c�2ŗg~��ҩ��"�b�1S��Օ�2u���xjЂLÊ��So����1]_4��[5fSy�����R]>^�z]�����1�{��"c�{�s�C����_��"���Y�ؓ�˰0��,��5�
��y��IW���>$�;)�b����3�WP/y��)��o:4�g][�v�Z�g���ocN�\����g�C۽��}tH1��.�g�V]�(
q�z��]��o]�{G������V�jZ�|�v��̒~��)$ؿW~_�Vw���W��nv��ۨ���S��^>k��t���nǼn�?I{����n�{��;�Cx�xj�s�VO�K�ژ�u۰�&|v��^��XtU	�L�*|Plz�x��i����м���S�����@�-"��A�<��<����TY[އ�]Z��':���X�ړ�X��e>l8/��M�����׼z��eZ��]א�=��w=�����G����g]K
X;,�u�g�F�f��[q�K���z� :�ۙ�G'��\�m�G�]��a�f�=
��d^��x�1xD߷R|�U=��C�����Wv��uE���W(���zq�{*�e'���<j�D�W5t&����Mz�l�F���x�o ၢe���4�&��ܩX�����׽�2�b��\-g�D-��^��-mL{$�/ݐ+*kK��5�Mk�s������� ޅ��}��7KE�y�,^9E!��~�O�n�l�gA�.k�֎���)R���}�`4�)�l����:Hsb�O�UD�۳���S�����P�ޛE+�u=�n�;��}�mz��t��{÷�p�D�.鵽���WZv�?d��7��`QӞCW���ۃx��'���p��>>Y^ڔ0Į�q��/w��V��:z݃�����։�mf��:_di��7��G�jMY��^�W�q�{��^�)J���ru��}����'�kg~wR_�Ol����(,^�d}SD~�y=�~}�V�v�J&�u:�y*v	ͱz̉U���@fG`'<47ܕ�C��$��|Q)����S����K�J�o�����(��N�%g�6�2cg48|�gs���+˗�>�+�uly�	�H��xr��Ug��pޖ��c`E���O�K���0U��þ^�V������,�Z��|�;������]����\[B��@|�v���Ə�׳�7��_�>�빾�t��}���}����s���o���U�:����ݦ�|>e��CY:�m�D[��1��w>��j'��na]���Q��{$��Z-�Ȝ�~���j9�e��_������_��	��?~!����3d6o#{�I���.�V6��e�)%Zn�x�a/=�8>��g����I䦆�g-���쉦�呐J�Ҷ��y�w�g�o}�Vl؁SlV���{���Ʋ�ۭ���q~�kU��f���C�{V������6�Ao�IW.i���Fu���ی�v�X����z�.ޤaCr��X��o.��g)������Y���S���E��ԉ�eEis�+hj����n(BfI?�UE6��������[�$mi�>)�y�H�Wu������p��]��y���xj{˭=*�V�V���p���f�Qo��f�l�nxP�c���������;I�B`�o����e�xֻ������g�^�`�^K(f��e�,U��u��}Ec����2�Y�"�˳W^�<��δ7{��+Ba�'Z;�r��d�C�.ߍ�����~Yϕ+U_������>��w_e�#uEc �E�R������w!�J����W٘1���B<K��:۾{e��:����j������v��ʗ�+�D�g���eΛ9�C��ͽ4�%\ bW�1�'�t{2X�K<3tN��A	sw�̴W8���S9��Wq�:
$s�*�*Vtm�#9�M:�G˷��t0�lj4P"���;�h��4�a����*�EPݛ3��紉'�:�.4Z��ĭ�Xp5�v�QD���ZfZ�,���i�:0���WV5��E b�t��0�ŸI8�J͉�V�wQ�T�b��.�Vē�1�F�����lg+g(ioE�u�yh�wω�@U�;GM���Y63�dF�wYO��9`m_ځZ��\ٹ:b.I���S�6�����8��2�;�gb�|��l�~����vk�z5b!�$��h�0�թ�:� �OT7zxc�2-X멮�r���"�O��h�%	7�p��n���8������MWlE�Ck#	&6�t�����&2��֬�C��p[p4f��e����gs�z��<�� 胹׫��%���0c{
�t2��˥ô���L\��Wo0���]SI��U�z��%*�.�۩ժi\�ٺ����.�w!;�lTWj6�.���D�4@� -��Dr��4��7�Ash9    O�~����)PV�2�Q�n�JzUQhZPR��e�)%)�PR�̈�rԄ$��,dx��� �T� jD��Jd��4���F�l�m����"X*HEi�e�j"�A�Ԃ��*(�4��$UĈ4��Qi���B44��e�$E�����=���F-�Cr
�S��DHe��2KlCr"ܨ�AV�Q�.$�-�V�[����������pMt:.Q���'�*+S�j)��$�UURD���#��~��]zw\��6r`c�OӜw���8s=�I�z��xҫ1��O�h$��O {7<:
��Oc���s�;�>KA�]:��"��x�E|�O���cg{cX�^�%�}���ó�=�J��I�r5�݀,s=�^�9��]�NZ]����$}{~�<L�*I��,����Y@�n��~4VU����e������%V�U¬KwCn�AG�q"�g����/1J���mި�5�lz��<�3GGf��zI7RI���mߕ�� �[�����coC�0��iCޞ5Z�{�y�������m��,���A��)��}W*'y�3I���`�b*��Q
��Ma�dwJ{E��r�0o|�<34�Ű&9�3�޷>����,���v
w�?��gك���u���Q�y�w��� �.��s��[v����w��$��ek�F��L�?[���o�ǹ^��-�Ԝ�S���L&�:ף��a��oئ 5r�^����e��7�1	��
y��:�}0����y)G���Z ~�M� �����8r�p4f�k��m�wq�or���<C^`�ͫ�j��Wm�r�w��U��
Q�,eW�����)y�ӹ��Fkc�uV�u�V�C���������O��uW��C�qR��C+76�TeTE��У��m|��)�"b�Iq��j��ʂ��x6>���F���V���*���h��ϫ��o���k��13O.����zz�/׵~�W�z#��
Js�$��C��RB@j��I����/8F�72.����=�.�F�������֘�uz)+l{��c}:O[�l<}��㓇���	oS��O���L\ϖLO����W]����ǖ�U�L���%�_H���M��K�˼������5�~d�����2���c�ܒy����-|��|��Uf�F.����NrQ�B%�x>h&_���}�wWR�)�z&�n	�y�uVFv`!�J���E�3"���z3�ۭ���I����{�g;���[ޤmu�[�:���zI'�۳���}!���c'���]�zY����o�*D]ע��_d�<�i,!�T���R��~ى����2]�E�#���9����V��3�jO���z?_V��nL~�\��:�>z|&k�b�;{�|Ѥ�{%ʼ�g}��y*_z3��s׽��J����N������Q�o��O;u�KV<Vg��!�Nr%{}���+I�R�,�v�K���/R���� ��I�%͏���d͗�+�*��ؘ�T�R��]�D��k�x��̥�7���'JK<�������Tr�B�(h�0��@L����2�v�6h��]�oe-X.���#�`k7�G�N�d��^Ԩf�l���N���Yy������� �o��O�o��"���W(W���/d3��S��N<G�L�Li��� ��Y~�+��p趼�ϣ����3��p��ښj7���n��%^����#���\�?����_�,R��^f���ne|V d'"KY]�z+�݇�ɡY{�J�)7�jpoe�m��zh���ev��K�3��I)���px���N�{�x�͘jQ���d�����V�ۜcLQެ��E���f2����{H<���U�yt^ss�@��H���������ќ>��8V:�F]����^׏��h��͘!��|oK�Ƽ���s�*�og��������{��W��ث�=1m ޤ:4PjY=P"��Qg���X�����y���o�_��!��m'ƴo�O���N�Q=�����]�����5mV��ZAu�۱���Cne�rI�3$�M�{���z�D��S���%W��%������t�}�70��d�!���<.�tڜ�7����p��Pn=4�Ǹ��OH����F�(�Е�=|R�	��^�ܹ�Q�&���ٰoO1�Κ���k=3�����{ׂ\�ѝ��mC�1�� ]-��r$|Wt�A�'��7�w<��Cޱ둴�C\i�w�`�a�~r�,�;�ei�w���^z�~ ���!5���#u��nf���$�s茂aٴ�S�t��B=` �fowI���i{�O!F^��z|�i��LK[.�lx:�)����~Jڞu�ԯ�d�j�)m���k���*�m�����n���x߅�%��0��ގ���ڊ�9Rq���D\ˮF��
��nԣLy
LTA�f{A5��L�(���/IT�
w^Z��;�O"+��^�Í��ݳHX�^ח�'\�,�킦�Q�|��:6o��#f�ٚ�J��Y#&����+w�R���ic3^��gb��f��-6�oJX�_rfC�d�~�n�{�w�1����+���7ٝk}=�ȏC�A�ā�ؽ�^��{��oֽ��6&�5�ȭ(:/&��wނ���y�����4���3�o����+���(F�����(E��\^?9�ҷ��D�moL���ɢ��O<x��ɬ���<�����j����LNV���<�0��6P��R�s"�>w�d
5d�l�1���#�����C���$��'�*�@Am(������|���Dcu'���J.4��m�j\�%�
�qq�L��N��?�^D��f�kT�B0))&�1�V�'��B�X݃Sm`�-l��|�� ɷ9��\s�v���8�]���Q��!�x��2������ָ@ނ��,�B���7U��e�ޣ!�����!��xj[��s�����@AP���/�P$�Kc�:�ܻ�MJ��B��C���[_�X9'���^�2�~J  ��O}|���a���,���YD��؂`����o/Bf��Qyh�_��Wil�����:p#�˥�^0mft �W�"Rp��%z�3ۖe-��4"X~㐪�[�"���<���ū�����p/]��\l=�  ��
`BI�&�x�v��<���V�g��Nixn�h������и�=�Z=�۾�΍y�hT�X��B�pz�Lh�9�Cw���G��Xt��>»�t0��y�^��?���� ��^� ��<�M�A]�ȋ�W��`G��[�#&� �}�Pw�,��5B]�DD0��Q����B���b�%P�Kٞ���r�a�xP	��_106� ���	͉����2������E���q"q:��n�̶�,-R������Y\0i�B�U	���\dٓ�^
�`�:�Y�h��N�YpOy�Ɉ�7�����=�Q�CSN�~#�C��� �;C��]C?�'�������'�=�6�M�]���2�߸�^���~��I�QJ�<>d��"K�xa�̛�z/�� �S���7!����;�1�p"8�$=��\B,��:���>J�xg��M��\������f���ok��\9r�L��ǫ�%�ms��2!߈Q�����\M�u(ǖ�"�.V�ܗ�v��H���l�����P�o��ˬ�T����"`7��r�C�}���rb�oe�0jH�P���"t�j#�����ܑN$y���