BZh91AY&SY��!9��߀`p���"� ����bG��               ��#[L	$�ID��	E$�$P)Jm�QQ!	6�QU@���B����%�B��"
UV�kicJ���Ҥ &�L�4�I)H(���f�V�͙m�J�T�i��HAJ	R6�P7�Z�kZ�����Ek/;ҥTR���H�*R���M4�	�t�̶�kp�B��K l�R������*�T���[j#mT����R��K���áG��$(�����o��PX��Q���[/g��\�ݭ��u����ݛR��붳5�(�{w�^��N��ֹ8xͽ�j���r[ڨ�nJ�R��Ӕ��F��JJ���{妩(p��_W��mAT�[<��)�O���o�]����:}/���z��{o��x=��C�����|�{��U��-ʾx����1S�y��EU;k����i�*�<E+�P�>��(P�P�JR��9���D�Ix��x���I_>��%�J�o�w��W�uJ^_<��|T�vj�i���>���СF�6��:�,���c���=u[�7Ͼ��4��ٮz|�U{j�P��/f�*IA*i*���JT����U*�����=����Gw�Q>�}JF��w�/��UU]�OwC��J�W'��}�P+�}�����o���[��|w��3��N����T�5�n��Uk)ob��B��b�R���ԓ�Ғ�(���_j�
��y����@���x�]7�YܺyÊ�U{7���'�f��R.:�ޯMT*���v�Ԋ�����_o��+�.���UUI>��PT�k��J�J��u�̒q��R���U*�R��W�xW�=�g�=@
������׍`: ܞ������7���@���Mz����P�Q��V�d7��R�� s�o�l}�w "�Ma�� i�ݙ�Y�� t���*��ov�@&��� �i�ҀSR ��`�%UT�F��JR��{�����P�-�q�xt�ў>��*������6y��7������� ��� u�n��z�R�*�tSl�f��	�!�JJP��_@hgM�i�iZ}�!�Q�/�x >����(���
���z
���ފ��`V�vaPlQJ(y���� ;��� q�.��ν�8=]o]�p�w=��@{��;]�=� ����`(��i��         ��2�*�@� 2d�)�IJ�� h    �L�����    ��L�T���h    )��% F�C  A�D��zQI'�&��	��i�ڦ���_�����?M~��~����ѓ"�}��+'7D����q̛��TU޷��[S�X �������?����AX�$���_X����QAo�~���x��m��`~�F?��lm��-������6�������`[0��-��%���-�l�ؔĶ��%�-�l-�clm��-�l-�lK`[1�l�ac�[clcl-����m���[�[�[ƋcLm�����[dalm��������c��m��[�[alal-��L�6��m��-�l-�������cl-���6��[g[b[`[`[0�%0-�lcl-���F����[clm��L�6��m�����6�2��alm���6���٦���������[dcl-���6���cl4�clm��6��[�[8��Sclm��-��-����clm��`[ٶ6��:cl-�l-���m1������clm�al-�l6��[clm�ali��������2��alclm��-��i��l-���6�������6��[al�m��-���6��[alm�i�6��[alm���6�M�[a���X���acclm�������m���l-�����[`[)���[g�alm���[���cl-���6�cl6�al4���alm�llal-�����[alm��h�alm����al-���-���clm�lv�lm�����`[al�cl-���6���cl�-���cl-�����[cl-���6��S-��-��a�6��q����6�alm������Al`[�-�l-��i�6�L-�lKcl-�[`[cl-���6�6�lm���6���٦[cl����6���Ƙ��Ķm��S��#x��F؋lU�"�m���[`邖�`�lT��m��V؋l�!+l� �m���ثl�*S-��V�*[N1ثl�"�m��
[
b���lQ��-���`-�L�"�m�;`���#lQ� �m�6�[`��m���� m�6�K`��R؀[ �-���[`l�(�m�6�`��[m���[b��V؀[`�l� -���#�
[m�6�[b�`6�Kb��+lA�*[m���[b�F�-1b��+l�m���Kb�أlD�1���`�F�l�[m���[`���m���b��[m���b��)��b��R؉�*[m�6�[`�B؍��Kb�؃lD� �m�����-�B�)lT�-���b��R؃l�*[)��ةlA�"��[b��أlA�Ō�)l� �-�6�K`���#lD� �-��6�K`���+l�
[-�6�ٶ����� m���b���`�1@�*�m���b�Kb1�6�b��؃lA��m�6�`;b6�`.��lU� �m�6�[b-�c-�6�b�F؋l��-�6�b[i�6�`��F�)l��-�6��-�6�؋�"�B�+l�"��Kb���l��b	l -�[#m���#l� �m�6�Kb��m���L� �m���B�#l�-�F؋lU�"�m�6�[b%0K`�lT-�%��Kb	l@-��`6�ؠ[�@� �B�.�[bl v�[a[��clm����L-�����`[6�[`m�����;e�-��[clm�����������[��clm��#m%������6ƙlm�lc��#m�m�l`[dalm���6���aL���6ǌ-�lm�l6�M�4�����x�l
cl-��-���%�clalm��-���[`[��lm�2���ǌKcl)����-���#-�lKclm���6�Alm����clm���-�Lm���%���-���6�m�[0-���6Ķ��6�٦�������e����`[t�lKalv�ؖ��i��-��6����lm��-���[2���alal6�[�텰-��-��[c�6��[clm��1�%�-���6������%�m�c��`[clm�h�6��6��6���f�[c�6����;alm����[clm��0-�lKclm���F6���clm��-��i�6���lalb[2�4��[ؖ����F��6�������4�ؖ��퍰-���alm����%��6��h#`[clm��m�ya�DG���?�Ĩ���w���u���}]��ل�yy�t]�r��.��kp@\�]c�{�B�P���k�������i�"Z{��`��{���5F�]���z��GX�u h]j��K3�ԑbp"�wqM��X��e	u1^��K�(�%�� ق�r��6�.H�^f��z-9�b���oi�W�U�.�u�v�e�f��6"�g�Ld�5���w���X�ĵ��K�\�À��[t�ٕ�b�Er�,с�Ǯ�����V�ط[:b���z���&۷D��-�gu�ޫv�$0[6�f���a�{�%9��XˬA�֢���^��A�9���yanݧ&���P��*&Gn����+lYx(a�����	��Ad�]�C���UK2��D�E��3 A�3i�&ϯQ��0ԪbۉĘH'/J\-���r�K�Sv�ڨqS��L+D]^��˗�p�1�r]:�m�F�q�+%&;�"S%����b��3��-��s��9��dF#� ˫v��C0Z&�(��(MӒ�e-q��1Sp����G>�/S�2f�Z�Y�P�F�IhYwo��Uyr��!:��1��^$�����J�M�Y�,���Σ0�[Q�9�ɛX��MrAr<�V3l��w�Y�^%N�9��h ��UV�2�VLbPe�T���E-�[�*��LN2I&�J�zvC ��(c$-�l�cʸ�9gk��fckS9T�1�����YJ��l�VS�9�	D�D��WSY�R)�0���j�s&$�WCU`$ɷ�ۼ��
ەkji˗R�.�GbY��kd4M��Vj��4���է+.k��&ޜ���x�X��l�P��w�7v^�	2U���aӨ,��!6�ů�vޛ��(p�a��H��)ɣA4]]�c2�
�Jx�Ū��Z��7bm�i�vCʋ^	2�V�����ub��ƛ�W����^j��X��{�6�n�e�f!�J�i�ƝDlU�����r0���t0cy����*R���ٖ�SdQ׎�Z��ͥ�e��ИhYb���E���4SH��
�Y����f�mD�=gJݧ�7t\�v�f�d�`�a��։�3�k�[@�q1�^�Tb�^��Ah�F������+�QS0���a���J�+aInô�,�B����E��8K�r;lcٶGM�w�sEц̲��I���l�l�N�	�7�m4�,���&+ƅ�ٔ���#lEwTS�n����)u3d�7W�Q�����Z�T�b����R�MŘ	jGZ��yYT��[Z���M扃5�@��~�#a�jSnh�c�d��j`�HZ����i�\�Q���/.�^@#��E3)����.L;�5[j��Ʉh9/f�44)e#�z�)t�Y�f�R�!��WB�Q�Nd�n�F/nd�4Q��-ݺ�bєuqv��&�HT��"�P>A+0[E�ij��Ѣ�C(hywo2���Y��6�V���1x(��6v�#�z�;ͩ�2�:R.���)wVK��J����kܥ�ছt�텹`�S3^W[�\��̢h��5��E'waIz�osM���ʆ�MRǹ6J'\�*T)E�!���5`��e���x�*�j�b�! �:����R`�����q��c��om�j���ئb�� ʿ(Lۀ����+��N�ڡdK�&��e��j���ul)AR1n�MR9Uz.�c�n�y �ee���W[��t�Q�mV�q�eD�,t������
�����V�i�XZ��hq��UV����Ǻ��m:ݏ��E-����v[�[�@��������-��z«��Zԩ�b�^�2ˀ�K�9��u*��!F�N&Um�*)�e�^m�@]3��h�w�ű��u�,2�6��E
c����ض��eeYv�QD,���mMn�i2��ˢ�n1A\���A��iZ�U�)(闃T�M+�6�r]
TuՌz%�����u��bB��:�ώ!�o�a0b���x��Zjˈ�t��PGy�v��V�UmC�Ko6���#^̞�W�����6���t��L�����嗸r�Ǥ���&�8	�سlA6��-�T"�H�ʶh4�`�ViS�*����-�6���c�{�.e$�e^f�*TN��-�YgT�F1���L�H�n��ZT��d92 Z͹���	� X�'v�-̀£x02e:�ɖuE��6l��b���� ���+��z�VF6Dcm@�ղ�wDw� �uk2�$H!�5�ơ��4���-җ��'�S��-��
����Bn�X���1p�Sqҷ
����E�˪�`ǵ�Nձ�MM��Ԛ�,�e ���N�Į��-�I��-b�˫�ZUXi=�"v'�]���W�'s� ٧J�2���
���OF��`Sn^��f'j���+�t�3Mݸ�$�M]���ħ�E��sc܊6n�٢X���d@T��[�*/�WM
&ً<�i�U��v�T���"���%fTr��3��<��c4.JcL��݆�RT)���V0[GcI�E�G3"չV��2yYN���8Tx��j��x��[N��)�J�V#+N�+�ı�;��w���~��r]k`�*�me��M� �h�+w+HDȚ�E��^k��E�ye����	��ۡ7#!S�ɘ��k6*+}W���k4�x���I[PG
����#ul	��6�6i��cȅe���ض��t5��6�/n�%N�NV��&m�F�^%`T���5��*�hV�����7�j�6�JhG������#v-r� ��ښ����#Z�J�^JH�.�l��D��J�2	T�a�;{�J���6}X��X��ڬYl�W�&Vx�d�8�!��P]�@�v��k
�Z�p�'�-:M*vMF)r�T��iM�q|�5�����f�1K4�%9	n8f#�J87l:�an[J�Q���*%���>L^�î�Ghܠ�V���,�Eʣ��V�{kK#%�X�x��n�JQ�2�v½XtVT)`�:h%y��1�ܫ�l:RV�V�kLm���ww� �1�Y��V��n��Y#�x��!�vS�eі�U�[��ض�7�TuW�EЛ�S*\�xs\�r�0U�/}b�t��#6�X*2�9oCr�7�欅I���J��E�<�T�`[��b�����''"7LF+�n��9$�gu���v�
����.�T�=S�U9`���!wDd�/aB�x�[ziGcL%�PV�Dm"]�U
��h��զkZ�Iu�����Cbz���ٿ�aW�aW��f�4�jj��k(÷L�Z;p͔Bvj�WCs���e;����lZ�E�$�l^a���� d%,ݒ+Hћ��Ĳ�lSȶ��k��Ms��*m��6PV>��I�k����hmi2�kD*�� ǙF�2]��D�YA8�ji���z�̆^�8&d{�����r�T�3*�7!(b�m�~1
���	��1�r�T����3^nj���;��i�	*�c�skǚۖum�X�8��Ez�mGf�W�cY��y�I)����A��k1�ݚ�t�������Wx~������A�7r���EPNm��u�mMS2^��6�����u����:M���n�p���l�=XL����rSv��f̹�)��Sp��U0*��4٢��d�)fJˏAj�9��PAR]�BbF�e�a����2Y�*�oe�12�B]�5��[o]G��#k.�wA�QQ"�f��ݒ�<����elm�u��7Zw0L�v/U�m������1�8U&���$8�r�0��u�Q[f���Q�I64�K�Zц ߍ]B�ԖA�=��N���[@[xF�e�5nMkZY�F�T��t����
�̢oպ$#�ӵ�X{J!++	@i�h�b�;{74x:�)����fm�W4Q͂T�n�	��;튄ac��+���l��=������q+�[V�M&��Z���	������q�B@�`�T���`�c^*苖.S�z+��X�a F�)˳2�Gukɥ�wWC)�7@1�°SH��].R�sI+�K)C���M�un�$ˤ��ַ&�f����J�{Kp�Q��P�8�8��nl�f:3f8w#uzE�UYoe�T��5n�����{[r�H�$x	x�+q;�2J��X�F�#I
J 8�u�d�,^4��+%4���
�eb:�O�F�ˆ8n����Q���^��Z��mh�)�*�§��l�<
�U�eS)DV���̺�8��j$���AM�J-��fƩ��m���)��*#]�0��"���A�Wq͗++�N�#zf��L�gF42ʽnU��^�L�aך�X$�P�~����%k��3-����f���b���%�d-���$&%��A��yor��a�y/^Xz���� ;X��k+i��*�M
^�!䛭���Ɩ�M)MTP'��R�7{���bN�l-�[Z��F��CwIw�N^k�z������a��lRH��,�`�a	
5�ظ�� ��h=9�Ȩo[��2!�CJe̶�D�WF�6	2�K��oC{BmV�����U�2g��ZiE4h���ɩ����H] ����"�*��^G��wx�u#5'o&Ì�5FkBPf(��ب�j�����uęD���Ѓ˼J�,K4+6z�*����n*�vn��t�[f�,7����l�µFc�q'���Tt�UL��,�'kM���*�,Q��p��^�Z9ub�v�鮺YY�^�0Σ��Rٔ*�-�Fњ�ֈ��|ru5?��t7)���&�A)[�%h��Q}�aR�X7�F�mX�UAtj�:ܙ�(�bh�q�7��d"����`@��إ�Y6�&�&ItDʭ�s���[�O5�r�%{����0U�m�w��9��2H�i"2֊Z�T��-Ǵ�8Uɀ��n��V�iJH#�� V�n�^̂m-�mc���ս�����G��:V�f����x�[��Ma̼C���*̼�f3-�q!�LRj�@W����B0m	�d-^��{yw^ �[��KoTgh�)l(�),f`�tX�tj�X1���z�E�n�DF���XuA\�Y,M�R��Ď=-�;�zwU���6T�n�m���M,�Ӹbl��@��*8%�z��*�� �Ҟą���m��;��z�Vn� Bؓ7w�Amk�M��k�*'C.AhU���Y��φ�^U��6�ٲ0l'j��V(�wV�X2�*��;���0��iU�K���G/o;Tl���<}G�WT�u��l��)��\�2�r�IT4wb�}׊�/�*���T���9l�K>ڣX�%yL�v�ܕ��ى�qZ�۶\���*���"��sGp�8(J���e����F	ΟV߲k����Y�*�j5+� �j����ya&�cVD�+4��r]D�6���)��d�I(�Q7tV8�ef�\�G}*���v�n�b�FK��H�%����o,"���*!oje���+&ʣ��f'���ĞV�%.(�!t��iMRI�7&�Z�!��6�B򌺋0����A��L��aW�Za�E�ʲ��r�d��y�9j!]�r��%	vwȲ�1��l�}��D�ܛsx�����y(�ǎ��Sw���=N�^�Qaֻ�YbF�T���5&.w��R"�J���ōF,��Ĳ�ʼ�I�q�2�T�A�䛷�˞β-Aʹ���7��.��ͨM\ݺ!b��D�[J��m�I���ǝ(�b����NV�Ɲ�+b��V.�<������*<�g��敞��CΫ�5��HJۼ���^\+z� �1y�����}e�KW;��$ͮ�����1��^�/�c8����4UDb�7V 0�(�k;��yA�X�����E#Ȅ�yaډ���B����x�[�I��$̲ܭJB����7�4N���/9|���l?e�D�o0MWJ�Su&�r.kPX�x,%��+%A5JE�M$�FŮiW��!��q��2�B��7�EӰڽ���dg˽W)��U��:�k�5dSa��9c�H*Wu��&!O�_
Λ0�t�����LīE�nn��%�l��^��L���-��^�}�$Yhׄ��	d�}������G:Fm�n;��,��Ҩ�9#職06Ŭ��}S�d����#\�ص�΃���M��B�GVb-�75�id0	�D+��Pi>0��R`���p��:D��͖���	.��Ǎ���[�X��$Q-Y*JhD���v���%1�beB��j/-ʩm�A"��ҁ�u����f\j����%2�^�	�K��I)�E-mೕo���B���/`ua;7jR-����%ZqƢ��m��rÁ�ZcQM6������T�;Y�r���e�cv�H�-�띜I�3yh�E��Fb���y�1/_u��}]L�}}&ι��7:dl���eޗkb.���]NnnFH��pcUt-��c�����s����3��kwr�iֈ݇Թ1*�u�콩�V��{٩����nG׹ԩ�i��B��l�d���i�-���Hu����@��
�d w�x�.���$�h����n�څYk�)����"�a�	���I��lOc�U�(�#�#��:�`]�����eNf�HF�W˲�BsYkb�
(���X�F�+�Z��:�K@Q�ϲ�TL��*�<w*xu���M�{x���G���a��a�U�CU�U�4cbÜ�Y7zh;]BE&��^�CK���V�;yo<��$)���T0��穵�:Uy*U��#h��˔�5�ث����AA���g��M���c�15�X%Ig@ȃ��*���n-�GI[]�1�33f�Jȭ�e!Gm�Pd&���@�3�PQ{�p�=���&�8o.��W��Am��Π�ˑ22��)
ӕ���y����z~��H��w�	��R������wwwwwww\��oOvewVk6�ѩ���3�.�{ܤ���v�l4��N٫,*w��h�:[�՛���b����m�#��Ӭ)]��0f_���d�p�&�!���6����z���F������9��{~�.��󠻙�c�x2K��oګ�QZ�{�X��۽62�\�����z��~㎻|y��U�]����!B���N�-��ѫ�Y�Ƈ<����h#�@��-�f`���W���Unu�:�p�a0�9N
T�4u�f����2xV����(��2� �� 1ҠR� �5���I�����U���ȷ��M�̍�1en�G�����@г\�|�X��u��A@��̳4;��̤�㭙���oN<�=T�}�.�hs|7�(�Y|mU����Ⱥ�r�;��o�ƨ=�v�=���WwqB�`��
��-=�]l�cǑ��-o��u_S���-CG��������J��M\g9�3q�f��-ܑt�i6�gB�B����Y|z���q�3#�^�8z�P����T��xbd�[�P�:����v��#����p��a�Q��ڑN�rng*��C�������gy2��ji��M���v�_*Wfm�m����f��AI�wa��Ә&-�g����ղ[pD7#�n\k)���s+j��'(Ӷ7y0�q�2���ryh�x\{:U)uxXYI��a���_g$�ā/��ov<����x����&�j�K��ܸ	a��_�4��=$~~]=�W`��Kt��� ,�CJ�|���fRe��3�h<�;�v�d���|��+]z��Y���t�Eg���޲��E�ܴ��0d��+�F�kJv�ں�k���Ʃr�̳�m1n��}���re�
wЉJ����Gtg�X���v.��e�g��W��ApdVnT�;�B�Jת�W�b�,>Wy�-��R�U��6�m����1N�t�W�A��f�I���`Į�]d�B^d*\�Z:�AYzw��f���0���=
�7�7��܀��N=d�2��s�2	#n3��vq�1:Y$�=y|mJ�m�p;�_e�KF���wc�V���\]KR��u���{�en�6���o����;K�Fa˧Ρt�PN;٪�tژ������	I�G+I�-&��!pQ#7I%���|�u5��-��c:A5_!�}�N��tJ���w-�b�|�۫��^7iІQ�|y%�]s��MĞ:V�R�4+�n���w���t�#u�4�B��Z�]̏��,칷����6ڶ�B_5�Bq��B�K����x�ͅQ�JؘJ�����.��^�މ�*b�;+�a/��.�k��g�7�-{t�8X��횹q'���7;�0^#�C2�e]�S�r��Qn�t�G�=Ϋ�W^�;�7YI�b���"5z�!���H��m��q�h������[�/;�cW8�zˡ%���t!�̡T/�����uEfnd�{];�+n8��K7��R������ګ�� 3)�Fh��Gm����ŏ���w��կ@��V��� R޻��s5��G�^s\�Ÿ�B�ѣtA���Ge�إh"�HR�;1�-+52Ru˖�o^��L.?�H�{鱮�*u�L
|E�YݲK:"�}���e־
d��s��J6��!�=b���H�)*\l���g���4i�K���ݗ��oG-a꾕8�l�WA�z��e��3W��r��A�쾎�sͿ��xm�=���<��d�)W�v�;i�K��2�[�&��"yj:Qu_0��inuM�R�b��}��f�"%�T	���l�wX��4��X�w��؝�ֺ$]��b�B�ܲIa�I���&m�;���Y��ʳwJ)��F�Z���Wu��oWɡ��_�հQ�����Iti�eN.��"1��7e��FΦ�̆9T�����U��4{X�j�cw��C}���V�t��<8 �T�vcz}:�r*���tJ���]V��0�xZ�r�x��C'.˭�{\�*��r=m����yRnn�hm�0�5S+^Өm\�w0^�ܠv(����m;,Z���a�y��!�z鬐R�Ao�Tk"҇d��#���׬9���n]^H�uG�G.�y�9�E��u|{22z�fgM�t������9cU���%�76sVj�)M�)ݪ��U���1�[f�6A.�w@�yF:p+�cu��D�M��#SI^��R�nA燗yvX�u�ݢ��c�wY�z��K�}��U����]��K�g��l��K^兼_0{ik�����:��o"����Υ�ͻa��[;���c��O��u��c*�e2��N�!��^;�M��>��p��b�p�)���}�wtm���^J6������7d�M<��|:.�FI��-�W�-�S����{fХ�+�3�^d����X-�.���=�gs�#D�ƭ���Z�q�O;��k&�-��-�tc��pB������73��"���!�4���d��LVJ`�h�f{W����']8^��g���95�7�h.���Xp2[60A(��]�Ud�Y>��B�iݹ�.��s-�K:o����p��73$�b��p Gw>�hs��i��ʑ�� �32�H�]��l��]��)���5`J�M�ށ��A�lY�Vp�{մo ��%�*�[P���Hi���%DsqX��v�����xR�*mNZ�#E��\]��3:^�\��ܹE��`���D�8��
�Kj��Qm@��e�{Ӻ�y�BD���L �FQ�Ja�9�K"i.�̧����U���KO
�J�aĩǙ�&c��#�����L^��[�΂R��dƧR�u����WG�|.-�����ZEn>�N�^ޜ�wF���H�Jՙ�]1h�%ٽ���UB>l�*q*���=/��R'��U�;H=vj��h̉\U�S�$��úŤQ'�.ZU�N��]/Q��0�r��C}x�vj�D��Ua=F��T6d�;��-��oyh#�[\�z�֞Wt��5ܺη���|���Y�Z��Dђ-�S��f_:�il�Øt����0�F����y{�΄T��&�9uȠ��w	PCs�������i�P�5�Yf��!�b�p^̆�+T�F��&��̷`�/zٹc�D�A�REl�BV%��P�o-j��æ�a�wx񒫑�#د��\���J&�����9���Ƒ��ِ�Yۡ
��n1o_L�����ِqmІX�/20�Ü�˹���ݏ � o:��ͱaf�\��wX�F^K�YahS� 5kD����`�q��'2]�J�u�{#��n��<�vXG8GƢΐ� (�Τ�s�#�B����J�}���;��]R�%fAa�H�3a��%puݦӮA��͏4�B�<�ڔK؛P.fP��,��Dk_)\r�ý�S�9+(դ����U����kQ�+��5�Ép�X���tY�<��>[�XVe�ҹ9�<Wʒ�א��t;�H�11tenⓧPM�YN�핖7�7�y7�����+#Du.�7�F�X\��;���Ǯ�͛G�۾�]�8�b��z�[��J���dEx�t�`������vy��hwK�����=n�j�H��Fs�J�sF`�͓��j���A;Bs���u��u��-'�;��n�.��<�ؘ�rEs�i�:\)f���[�)��]�q�F`�ɯ�+���͗T��T蹔���Y��U�N��V��ݧQ�ĵ�}�!Y4�x:��|Nއ�[4R"����Gs�d�s3�������zu���_��/���n,�87������&Ҡ{j�Yf勋�/-=����J�f5
��E2�\]��J��o��JN�=�����ݾ`����o��:$:�՛Ê��r=����3��;:H$��fVk���unD��]�t�u��f\��z�xb���u$æ,�q(j���8��G�2���G�%]����h.��fmM��6(m�p��맬��Zu]�sB�Y�9�2�H�8��e�r͎����{���M���ɜ�p���۰U9\�a����sC�����'e'�(�<��+3;���y��
W���}�P���M�Xy�A��6^q���H9,}������-�ܷ�Ht���Rz�B��A�'��du(GH��9�<�ӻ�v��I�j(v0^Z��;���&��ku�ԙ[���kƩqr�X'��@�j�7���]��9)P�k�����C鄣W&���{�;�P?c��O"�t�����>�n�]k�|���늁b�'+����������{ے�U�B�V���N��oRsS��Q��:S��p������{+=�:��t)^�BBꔹqWr��.�����3�P��(l�F1��/���k"��j]wg�&�A�&��[�]c�*��G,�9�����ʗ��oݺ��t
(���V�2]�h��υA(��N�u��y�a^N̥	q�N�w0��;��t���ݝ�fp,�WB��T�X�>�u��h�q��j'�6�LӾ�o���K��VR�V��R�<�+�{G��U�3-�p9�,w�wH0���3/4n�oI����R6��<�&PÍ�8�Sγ���k\�n����KT����3ip3���si�4�ͅK
�VB���.i��3)�>vs�S��M�͙����*�{�j�$�@�9v��S�Μ�<So���k��ܟoU��4>��EVf�Tv>$���7��m�o�ף�]z��ӛg�uRR� �/4^��גn��+�ҏ���@'�V��&+z���d�`x�s�������
}�NN�#}f�/o��Hc#yf�b���k䋥�:��ڥB�Fz�_3���Z�hp(����AL�����:�Oz9�Ϫv�ڼ]�\���C�1��\�֏T������<�{�u�ڎe��^�RY˅'.�h�$v�҆��۹g��;}��K�\�s��z��>��)^��Ǐ\����.���,[R��K��8N�25*年8�ER��Hk��M;�s�B�φ\������c�1��4��m���[y:���d���a�p���ȉ�m�:!m�жs��$c���i�Y��L�t�����������Ғ��a�c�g6Q���zwe��������]Mv`�`�͍���u���JN=����ή���E��s�sq�v.��]5�*)�D�M]Jgc�]�pq��Z$4��\;��%vc���[C3�U>|��N�lz����n�;.e�*���s�2Vj�>9�L�������Ϋ�w�wwI�wws��ӻ���wwm�wv�$���
D�\q2�0�Bil�i�����l��V]��e��[�id��i\v[��m�����������;i���M�]*��l\d�;3�<�d�کD��	Y�l�M��RB��e��M-d4�Mӑ�:����i�Y���xm6:���YX�����!y�!P�ƌ2�����.��yh_#!V:����R�rF�q�ZD�M��kc,X�Uݾ��u���"�D�	�#"��	�D�I
lv�*0�Vm��iav���&��O8]�/��C�5��.����v�&���&&��X]�#i��>m�i&\�S���6j����#u�]�Xٵ��wnٻ4�4\^�4�4�V�f:T��X�.�&�v�.���-��[KGy�w��$�Z�,�H��q��P�
K�*�LA|hC�R�nzu�x��L��!T4�E7�-�f�����!PRP$($*r3` W%���դ�l�Ը-��+��p���m�
��3�IԆ�N��Ǉ8�Rh��kf�6��Hnɻ&���[9��#��7M5��$���Ҧ�[��j�nCu����I�B�&�M<n�e��[	#,e�6Gd�j�G,��*D( ��欩�w�c�Y�GZ��y�a ��f�la�]��HF���$�]�V_m�+D�,��q��P�
_%!T�T��n*NoV�9��&�v�.���-���a��i"��N�4�T��Ǎ�Y��č��v�cf�7]�ƤP4�3� QM>�����+�	6"LM%Ұ�L�v�����\�[h� ��a�?0��܉6,ZYd)�۰��mY�F����[GRPI7wtH��g�I	-P�5	�p�]���m1�؈�$j0�im6nY��4�d���9\�Ud}�<v���^Rʼ6�M��jl�V;��m.�I�H�S��s�e��,�,�TjPZlZ��f�	Y�l�M��RB��U&B~O�jk6e��ui��y$&R&�������;i���M�'�6���M�埤iM��&�ryV]H��B�%6�HY%8��Nu�a��,���bK
����n��30?_�߬��"(�����pS�EAS��T?�������|�_�\�[����凒jy|�+�UD˽�����dn��EhpTg���l�rZ��w��E9���gl,1�0>���^ݯ6w�=�B��K���oz�>����
��:xU��S.U�}K�;�1n0e�0F���b�~/$�.���R� �H����|I�B�q�#u��Pt+v�5�f���"se���2h�D',�F���T�����2֨�8�Tr�
�]eui���}R�Y�14��}.�=H���z!ܟT��e��f霮�P�'[F^�ǋ̶ٌc�vv=��hs�g���:,��ܬ"�\fv��"����nv�$��^o+2!׼nG�U���KY)����d��m����1\�]��Ԡw*�Dԅ���e=��`����׾�}������hl��whձ���Krt����Lr�9 �Q<������: �t8u�\�w$6��M�����.V+�"�Φ7S^�J*���W�h�1�;��������@S��=`[(خ��*Zf�q��h狂��Q�M��eIv�-�5+���pp  ���.��wY��5jc2�n�o<�U�[���s�����}|x�m;vӎ8�8ێ8��q�n8�<q�t�8㍸�q�q�\q�8�8㏮8�8�>��qǎݻv�8��q�q�}pq�q�q�q�q�pq�q�q��8�8��qǎ8�8�8㏎8ӎ8��q�x�q�q������������q�N8�z5�/{��kU��]�C��X;t,�!scu!��K�}sv��^;���%\�C�p�\��ۨ���>O��|~�����K~OU	�p}��؊���5�6������<b�z읝T�Ӛ7��_R]�掋��>i���r���}xʋ��gR9�"�=����^7��p��7��[�S%DS�F�#̑��nn�Q�M^G���-,Z�5�L%�E���E�QM�4j0����κV�f��7N�P����a�f��\u�\Z���]��X���U��^�^ӈ>a�v�ڒ:u�8*�
��i��u%�*�(������NW]�p��3(-��w�+�m��Y��LuٝA��,�PZꓦK�}bb��K/a��J����P��������y��$��'	�
殪T�!S����|��4,�'�L�+R�륆�2Ó���ޖ�>Br@�r��O;���+Lb��X �Ţ�9�#D���&C�ӛ,ΰ �U���bZ5Çv�� <3;f�ӏ��'�5*ͥ�וwB��F�DQ������(5J�����¯�uE4�+��дu��m;q�t�n�;c�8�8��4�8�6�:q�qێ8�q�8�8�n8㎜q�q�c�8�8�냎8�O�q�m�i�q�|q�8�8�>��8�8㏎8�8�8��8�q����q�q�c�8�8ێ8��i�q���G������q��8�s�7��p�UkpwS�����NW<\4{'��f�4@sOm�\�arF�UWsof���:�:� !�	����9�mW��ʸ��� �\�h�t�tq@��pB�Gmh7��l@�ξ�7|B4��VPb�y���x
a)K��4�W?CG5@D�� �!EZ-{�{$��7]{zh�Qy����v���������������o.
�5}���H��񳵩
��B8�]~�a�J�	ґٳ�v #ղX�b���%.�"�x{����S��}w�D�=�z�a`�r�5>�\�@XŇHޚc����ZD�#Kk�Q��f>p���^)�+�uв-�sC�w����mTu�� �<
�NZ5�W^u�K�LJB�hNe�!Π��Gm��L���]�|���e_c��d�G1Y .��6���B�CH1�N+}��e�:��`T�d/c��ʇ� q,o6�u�۲�����S�Twce��N��_<T�
���Wϩ9�nb�S g^Uƍn7�3��v{� ^).��E)�i��
�)���(@_h�����x�j�iI]�)���L�x�QR�dSN�߽�C�π�
��40���P�+w6pf�]���CܹHLD�G�W9�ZՋ)���G��ww�/F�K�� xoI}R���.�n}�J�K���DT������2�Wm����j��J��wQ�;j^��ÆG�>Λ|qs�Nk���\��7����=�/SW���m�m��Ɯv�۷c�8�8㏮1�q�q��q�q�q�8�8��q�n8�;q�q�8�q�m��;t��qǎ8�;q�q�8�q�m�qӎ8�6�4�8�>88�8㍸㎜pq�q�q���q�q��q�t�8����������8����w�ң9^x�vÙK�tº��U��癆��Y�w <�^8C�s�Q���FQ*����U����)w �.��L@q�.v��RL�����v�G�w{��Z-�FS�+��>�P�U�8��;���[x:�Ƭ�`�z����5�t��dXk�W7��糬�c�<0���`���,�*V����ua�n땭2��8j'Ol�^|<	 �x<t��VFfs���}�$V�y��)��q^u�}�,Sٲ�c�1_wp;��X�B�M�6��6���w.�1���M�"����G�������vw���W(oQ]�|�8ĺ�qI���jJ�5���N�t�D�n�*m��Co�~����1s����]��M h:r�/�]*\h�����'c�Oe����Ϫ�9�vͪk&o�*�6�[2�&�b��	�����U�2+�]q��s�N�pUQz�/�m5��w��lZ�dk�-��`�7���3u��9�r��E��I�]:e�, =t�(٪����v,����u&��u\�$:�$7�Z��e)�5ٷ��)��G��W�P��h���tC���׭N���,uU<�/:묡땲ݕ��������z8�۷n�c�8�8�냎8�8�88�8�>8�N8�8�n8�q�q�qӎ8��q�x�4�M8�n8�q�x�8��q�n8�<q�qێ8�q�8�8�n8�q�q��q��8�8�n8�8�>��q��㏮�__Z}}}}q�q��^n^��C~j��y7N��Vf�|������xv��+p�1�dϾ�z��Yu��zj�ؽ���bg�f+���v,H��	T�����:3.���]�f�r=�'��$�6{3�9�|z�s\��}#A�կ�r��h�l��zŅ���3�2�7P2�W��QiX�Y{O�[=���UFd�W��wsU�{����J�=�uAX�#��#����Cu;��Hr���A��_K��RN�w�w�9[�ԛYl@�6����p:6�-r��`����3d��iݜ*ΓSB��bJ�+9�n�,VTg�c����K"�
9q�^)�7�)1
�T/(G+��\2<�f��D��V���[��QWPD�{��1�T�`<.�[��>�3��k�,hX-�z�N�J��5��5�h��X���pK�M;�m�5��x+�E��g����0p����e芄�`�L�����<��mV���n�B6���3d����U�r�Oe⊸+a� t�A����/�N�o�%]3F.��v&VN�M�c<��G;p^]�;��u1��fv�ܺ�͕���z�B^[�*���>��q��v�۷n8㎜q�q�c�8�8�냎8�8㏮1�q�q�\c�8�8��8�8㍸㎜q�:t��|qƜq�q��q�N8�8�n8�q�x�8��q�n8�<q�q�q�pq���8���8�8���8�6��O������_\qǎ8�h�\���g6:�/�_����M�,���}���"6�Tçҭu5jE��B�KڒY��wvm6&�K� �Ɇ�7�d���X7G5�R����;Ij�Ƨ��ᳺrU�����O�ƅ�
�n��7O�6#��I7��b��-k��i��9�n�9�s��xs*7+�4���Ӽ1rݬCjꊫ\�&?[1hÏ:��f�󎜜0�{ۉP[J��r�r������5ctIB���v�mH{�>zM�B�n
�v��,K�v�����/�Q�z�P�Ԭo����{(�.XN
����|��b�3V�U͏�7�Q������VliTUu]�NP=�y�w.Wj��#ۣ1+��Y�KJ{�|��:��*�Ӵ����ǆ���zuQ;�Ӟ��S����Yy���R��vfP��Ԓ:����&��E<�^�����\�.�=��c+�>��E��5ٻmҡcW�`A�zwz��66�,k��I�_WNa����L�@�"/z+����$QUa:	�C�E� frF�*���[vۏ�6��ݻt�8�q���:q�q��q�8�8㏮8�8�8��8�8��q�v�8��m8�:t�ӎ8�8�8�>��q�q�\c�8�8��4�8�6�:q�t�8㍸8��8��qێ8ӎ8�8���8�6��O������\q�n8�7d����+{eR<��Tǀ��р,����r�+����޼�hy�G9�y�u����w�1w���%a�W9h�L����ʔ��\4w����SΔ9�2����ӻ8vv�-1�40��6�썞�]"��p�]Ji������J��N$�6�Y|�s��ӋkK4�&>���=�T)��~73��,�Ղr�N�w0g]�Q�����v7�Ʊ&��_Xyz��^M�7��\�1���d�f.ۗv#ߨ��L���=�t;��XW/z�v:)�7�`��N�����ƻ{���8Ȧ N�u�]�R�+�e�S�W��e��nv2��Z8�L��ot�\��]q�jOBX��Nn��h���v���F���^g#.�̈9��&bz0+7�m�u.x.�T|�K��CeN����ܡ����:��11m�w�x�6���J6�7��s.�n��@���1r�q� ivv��	V��.\k{� �XV\���]����&���f�7N$��y��ʹ�LJn[��F���y+/l٠��M�E�ׯԋ�R�:Z��gm�S����W}y�2`r�9RMX��aʏ�\�6�2��2	](�$V9��u�h���WvD�;d�dŕɎ��\�A�m��A�X*֞�㾵u{ �*�C�'�b{ύk�n�ۈ#>2����+;��[31��oz�"�C\��BE۩�C�u0̭D�mu�ygF��d���(�p6	t�.;���<��w�Ӽ�:6��m��W%�(�I/6\�{� ��;�$ϻ#�'\�/aPv��W�Bס�}gR�hͼ..�ȴ\��z{6�h�}x�ucb���B����eU[����J��6��EņY����9�.�c�:p0d��T��v/�J��pG)if�&5)A���d���V���9YaS�����V���@�%H��{�m�n���t�o=�s�����_3h����"�߷�� uk��>
T[d��{�A���.���oaUz�p(���Vsޗ���)T��;t�F��$��W�y�|x���ET:9�	����k:�)J	�]`o	��`��ӛ"���5S��J�{���wpc�*� *-���ͦR_-ɏ����ޮ;ڸĸZ�ݣ1�$÷5�U�/����Tq�d�]1��iˉP�E�kj��o����l���G>@���tOCZ+�ݱW�(�Q9ky���<�����Z֌#2�r����@��ݗ{�rM'IV�b����med�J���p�ξ���=|s����"��:)Da��#�u�&	�Sl�+�ɜXE\��n:�q��(*m�|4o���;s��BV9�&�G�NR[&�ó{�Q1��lɡ���v��F�d
�:�ǁ3}�n��Xn�����:[EGr��{��ty�6��sv-�2J�kWq���9BD	y�b�����Î�N\����s�}�/��o&+6��o��bY��m�9��X3��7�D��7�eދ|��/f�	c�GYGNUn;�tl����9�^?i�4�q�1��P��q���Ng��Hx�����k:v��RA���P�>�����샗NWu&��j�\y���ˈ���o\�05ٸe�ُ�EZ:����m6��[�LCMe�7B��~�;Wǖ��R�+ =31Ր�;&k:vV�U�!�m;4�����v?�����Ǔ���T�Wg×/�Ү�Yr���/Jn����\n����On����f��"b�K���P@�$�g�*�e�K�[Z*4c'�%=��L׳�u��r��R�lpΤeV��i����ٸm��x9}��lN�u��	�m�wY+[Y�u
+q�;Q�5�ѕ���ϣ#�+�U3p_F�k��ut�j5V���
}i�1�׷Gy�]`�bFZ	S���(ʰSǸ��3�FM�\Yrm��s2����L��BM��d�Ӻ����xs�R��15ܮW��F+��lmɋv�u�8-����3l1�W�� �;-Sꙇ��!��:-\z��U�}����kyhLU��"i{��wur	TM�����Kod�.���W��4,	Z�G0^)�(+2�4n�÷mEH�q���98��,��=���w,n�Ƈt� ���n�ڔ8����}��.䁣Ժ�ƍ���Úî���a|1��:��^�s	��i�"wfw d0}�.�[����ZTW;����n�L���}���[d��:�
�y�i�q���&����A\UI�u泛(��'���y�����O�
*�d�����>�������W�V/�]���Mњj��*0ڐ�����(є��i��m��Պ��A4�Up9!�ѐ�Y5���ɰ\���%*݋vn�;d�H-M"C��uN.�F2T��r�c������A�����U�?A��t�j��n�Tn�0#x�V�uʆ�xN@⻫%st�Z��� �ϫ�H���UXe���U��
�`�U�j8��z�&�Q:t=�.���<w_k�NfR�p�GX����s!���{[4�ɛQ�E[�����]N�������T���퇴gP��$�E;����hV<�J�k��1���p�\-��zs)����y�UG�)�eѫ�|k|�����k�f�nBj�]n3fr��o�t�+\����ΖL���>�]�J^eՖ�2�@�2e;�M���َ�<��w+/i���F;H�+���_]F�u_*ɂ�3Aru��q]u����=n�ue#�E�Bq�Q�27���$̇��X�%4ȯ�,������]��*,�k&�%�(�Zpk�W:X�f���+bF�Ψ.<��v��hzjl~�����C��'.�����Ɵs#1p�����>�_h�5o<i:�7���Ƌ�Z2��4��;6#/�i��ŗ��%��Ȼ�8u��ތ��~���N�%��q:��.�};�s��^Y�5�r�p�E�%����u�,�`��4+���9��5�6Il%.����͐��m�eӦ�NCXF.���f�wF�3j��	e�P(���6EZ2��A��\�ݱwf�M�:�MI����[�6�ʹ9rW7v����"��(ѽi8o7`I����ۭuݳ�q%N6l�t�&��I���UD�:��Nj5 L�����*G�n�m��#rN���$FD�H���f�&))&"�ɑ�X.V�w�UE=����.L��W��<x�����1�2Q^V���P�I�"q�f��'�����⫊�g@ԉm����M�:�	�J�'��v�F&�DHl���Bttӷ��z���n�G��Zc�C�9_�����9�Y0��X
BHUR��ME��D* I0�%AL
�8b��2"�8I3
&T#���\̮D2��:�Us
�� �J��C"�$ș�\�j�$�1I!`�ds��X*Ct5�=���語J��m�:}|x��oG^����H���I! ͤ*L0��Kh�)c��R�X�L
"5��R���$ΉFȰ�IF9ř�V�	4j�2�F��"�ҧ�d5*P�n1ӧ��<x����׬�>���Q���r`MH�Y�2G̍��s-,(8V��k�8���\(�/д�9Y��j���t��n�z�o�z8�֙����E��V$�g�s)��!�>خ�F�J�iF�	�*�!"HB5��۷m�zۍ���o��^���r�ʎ�$h!UEHH����E5��$�+E���G#E,�-��1H����.��&'�VC��h��Ĭ��FBA#�'���&$c��(��A`�BG8֤�V���������Z� �!D�Q�E1D���O/%�=ͱr1��*��AǈɊ�q���w׀< �Ի���jjחv�)!e��.���G�)o̵���e����Y?��{���ɍ�o��\����q��حΰ��I[7E�f��IE����)�G<f�a�$\u4i�3�3x�=rƖ�/���S��F�Di�B(&(����1�P���e��n��TS�R�MѶ����m�C����~���{8�Rk\�3WuX������z6Q��[L���f�y�9z[���w��U�-]��w`��яT�-�"oj��m�9 ;�i��i����/7���z��Kqx�<�wD�1�$ܟW�c�z��D�ΚcwX
�����8�&����w�-r�q�������f[���2_c�qz���ˍ4o,�y|pe1�7�g�z@�9$������5�~ٽ�o}|��{�W���Ŝ�����9���xη��lv��6򧏶���ح�V����亡І��������P����5��{�Y�4����^�� �׶{�,�*�	j�h����b�y-�����/Ӿ�/>����n�m?O1]�w��r���vaX�H8v~ݞtE����gyg��f��x��y{K�Y��G&@����奡��z��ɂ�������θ��H�7G��W\�>����J��Ɋ����,>XI܄_����M{�vm'ݹ�{`>D�����ǵ��v������e�>��zƓB�#ddq2�u�M��2rjq�{%�}b�=w��l=pf��r�s�0�wtmvF�ݗX��>Y�;������A��;�B�"<�^��q�0W۳;{�}eT�����wK���][��hP_r���3Nj^�{��Cڜn��;ݫ���.�����:�����O[��$�l�K ��7��^�r16�������w�.����ݞ��$K������fƖ��i�P�J8�p�W�&=��J��T��1��_��U���k(P���)=�p����؝핃��k:��[������~���?=��^d]�u+���ǹ����i^�c}�5>~/�I�c�xv�76xÒ:�6�K0��zkgW� �9u�7M�S�ҝ톻��,�����}[�'{��Q">�9O�T�h�q��sۏް��ٹ5�k�|��"�
Ej����Q�;~9j'`�s�L߾�T|���>�R��:"��<�/���m`6Z[��^L���w�!n�Ώ��\j8�N��룳$�* Q�����=޾��g���5V��_wh�A� ��"$\��a�yy^�%�U'���U� ����9���+KF���GFcOv�	�Y�s�����ҫ�Ͼ �BV���\�%׺_�]P�o�[���|��^=���Cs��д�ϕ�*4�yB������7^|��,Z�������^�wz=���50CO
��o'%�z��f����4]O���/�u�ܾS�c}�{e>�v�U�Dq�ylyx����c{}Y�O�X��Z[6r.��$��-�\gl����;m7�M0я��5�T���FĂ�p�ç�sS�{�1~ Q�l�9�vؿ���m��^��ݹvӽ��Z���yj�߹XY��~HC*�O:U�:�EUw/uI�\�y�@����VP�����T�	좾�M��7�����3��V�5M�E=����^�=���^�~�ϺS��G���V�n�c1�ʅ���jt�)�Ts�d�q������6���嗹���.H�*����!���~��N]Ϣ�(�׃�� �Q�Y����C�8�0s���x;�9��ȃ���}�]]{��g^	�i���Ն'w�5��=7��~��x�g��{vՅNR> �A�����h�z���GID ��|3m�|�>>u9�߷�y����¯;@֫ޖ�۞b�)���5��u�^�fٝV���;�0��;1��&��o�ĵ罧;�z�ӭo*+,O^��[�+7��z��;�ϲ
�;�׌!��^"rqs��u�zv�<\UyLTm��|��3�{}�Su̞���n�O=NN�g�s�g��:��ɼ��Y�4ѡ]7��7��[��V��uW{;<�s�R�;k�����[C~k<CT�,B�2�V��?L꙽��o����q��K=:O��ٝ\k�[雕X�5�M�\|�|}^�&} E��GE��۝o��o�ؒ�ܘ(y�%�{3A���ݒN������ד���>�YlI�N�c���y�8����|uu:��ci$K���kH�Y�Fj�k�$)&�t=�OX�i�lV��������f���~���ӻ�$�V����x�M��Q�ۓFYuF3anݔm�Yev�m�Uiu��1p��c9���{��v��ڊ��� ��5�����S�n��Ns�o���ھ�b�~<�ԃЭ��"���:�`�;����O)�Nnv٭����n���Z���{l�^R���h|k[�^qr����J�ǝ�n��m;y{�L�3G;�fg�Y8�~3��.dc=e[5�n�eȌ�r��w�`�rxoP�I�d�(b�y�^�K|IGކ���m��t%?���|�8�d�B�su[�2sW*�S�	�,�L��;�+}�<�Q:G��a�����	�1�_�bX\�݃6�:����Bkג��iϜ�޴��/����}(s��>�ћ;��<H�T�>r��潃�A�P�#&�3��������\��p��k���j%���N���	��U/އ�` �r���<����P 
[AUo�7�Q����Uv�p{��0&��L�N>�lQ+:h�<�:v�AIh�Z&-�&G���F���P���Q���z�m��6����f�9����J�\�\���En�M�5Ҙ��m����S��L�1ƞ>����AU}Uָ�h:zc�葧GH��z���p4�vհj�b�
���7��h�y��������@�����m�>9<�9�����h�p����}�,�JJ�]�z��o�O<�>�/�곘e{}�@��;-wػw#����]���F�u���]�e۠�[�����8"_z
����c]׻7h�{��X�1q��C��pg=��}쫋س�Xv�-E�r��险�ק������r��:�j��1��tz�d�T,�g��}�;P`��3�]�zXߏ�v�n��C�1�ް�/=�*�{��^El}(v;^�<t�]�(q�1C�Ǵ͙����f�Տ(�����o���˛V�Ь�r�����2?j�xyY L�5+��s��z��N2�^�B�~�7+�u��(>����V��neM.����P��y����G&>�����ي�nJ�ǴT�e�֓�6��X��WO��>�G�Vae��
����.��W]Z�პ���/�J�7t��9Q6��].0�u�Qnt��x�+jK��\�O���Klo���ù����n�7-�{iI�r%�Y�@��I��}^��|s�{k�Y����O|���a;P�}�?>p��'.[{%��ӣ�{�.&k\�ޞ���w���j��O����i�"���6I���q��]�t�77D�i���'+�s����ݹ�o�����Uü4uuj(CJ���\�����ɽ8���*�XY(����4\G��N���4s	�5���IK�h�-n{���w�=^�3W�tOf�=��a!��A��[��eA�{αK�]'o}��}��!Oh%Z�ty�}��:k���3yn"�Q���`��\��wr���s�Put�.��{k3�lzY�k��j��X'�&���	���I�+=�,��@�������
ߺWϔ�}~�Uvu��=�5��ƻ>��Us� (vsr�o��)�l�y���/���ৱ�t�g-R��7�1Y�[l�^E f��d�� +.��W��ӡTة� �GZ&.
e$;�t�%ś;�p��z��ݓ��s�a����v�'��"V��ui̾qUU�wee���#�L�����H|7�d��*�0O9�T�{.K��U.��ԯ�j&=R�$pzǒ�B)z�ώ�e�qE
�5��!���ÛC�pM�@N.���ý��~@5�&�bd�	ޤ�;���0��Uyc=2��Dw����_�k^٤Ru<(�ν �k�/p'�kZ��zIRT����1�I�R{h��{O�8�t��9����o�����H�N䷲�/w��!S~c�����j���x���K*���E,��{�;e��|3y�U9�x�>��7gm��vrU]:��5#d����m����s8��58���p�7��^���t���D��4_����פ������^���]��B�͟KޣY'��w<���[�����ŷ����}5h���9�tD��j$��@�K��na/�ϭ�2I�:G��]�=�Zׯ��5�Mh��U��s�Ę0���2�Nds��2���䓙���
^�#�q���G1B�Z�hN�EAQTU䈪���݅sa	+P�ԩ�"��̎g\�\�[6�.����/��G5t
�۩��I�A��W7�Z;����V�6�+��4v�&��A�@A "��D�-���K����i�2a.��@r8@���k��`{%���)��� �4'(����>q��C=��;(�c��֎�yr͙�n��1�zɛy�;��F߹�ҫ���V��S'h�yƉ�k����Wq����8w����XX���s���W���ѪzOw�/��.�Q"	ݶ�c~j�߽�gv�.l��3�Nܘ���:v�8���`~�ǀ,���\~��ʇ��ײ�g_���ԭ=$�Ms�n8��-�>^�7t6^�x@�y-�t�ˣ��N���s�}l�!���������]_g�uT���,�2�/���z� Iދ�~�� �;���{NU죺F4Y^�o��V���|+]y��ߤ�� ��P�"���)~�W���;<����ذS5���&o��J���<o~�>��ɇ��7Ճ�ej�h�eMX�ė�X����o�����ۙ���>cIX���(��ڎ��1���a>�*׀��{� �Y��VE.-�= �Y�m:��^fs���C ������Wa�Ϊ���7�X�M/j��<A�y��i�Ȓ��n���{�Psә���'_40s|�"y�U���$�U���ӓ�L|�����ͺ/ە��3���{޼Z�N���w'�_����%�}T���/�^ٺ�IG�S`>#���O�)�ws�s��q����`|�gs��=�Dwۜ]|1n�������8�7x�����sd��+��L����w��ϵ��ON9��SGw@��5��W����c�|������fVkn��|�C�s$���ly������f�Q>�N޼a��s~��tz�+���Oz\��1���^��3�������.��4�����K����<q����g��p|�O����,q.��5Eۧ{�N�]}��"��?i=�������ζ{ݦu��y~�+^������6��~AW=�c��̝���<�V�h�o�g��˓2����
1��b�jt���S�;Et[�u��M��9*N��MzCY�;y8Mc��]��zK��c���ܘɓ(Z6�X���-�WuqUo.V1�wo���+gq��@ȧ*���/ 7�}6>v��]{(��Λ�tj}�e��2�B��f�Vj�����T�hl�a��"�mْ�d�F�A��T���z#j 7�Z�X/w{8f7 ��ηV|6���rTJ�t�ì����,!B�n���y��_|�r[�z���J�6l]	j�Ud	:T�m�k�����t� 8p�c)�S�i�Ux�f��x�dCcp[��)Z��A!��ܺ�-7��l4Z��t][�Q�*8p��}x�l]K��DWlv^�{;1l�<�	��cK��S�՝3-�k�-���w��2��-�Cu}7���8��dy�n?�d�k�xN��X��n1{qk��������8$�U�sEoM1Y��P�>���Ň-�E[�l�хGG�t������snZ�ost�n�)��i�}͋Qt�f�vC�03����1�
�9㓫E�&�3GU�R�� �ѾyT8�S����l�x�]n;b]Z�=ha@�ۋ�:�Ϻ��ϑD^l/�#z�9{�z�7qZ�����W�c�B�/J�<Qp�V�
!�@����0�Hh�;:��^��]�}�����\d�7��o�E
�~��Do�r���h�f�P��5sWtTyt#����Pʾ��r�����:�7��J)s'.�������Y�J�Z�[h5�^]� �PJ䳋!PX����[L_<�/�ѕXU˾b����R��Ռ�[�c��ob�k2*��t��뙲c{�!��]�Q؜�[3�'��\����3�esІ_,u��kP�,�K�Q�p�c�>��,����Y��]�3^Wa�F���v��%��h:�u�cц@��e�R�J��X_*J���&��1!����������񋷯�yYx{���cMj*��ʍ9�1��6�����1D�62]�;Z��R��v{/M]fr+���g�VtX��_@����k�L^ۣ�]�Mh��x��	�-D�"J��%۹��E��b_M<j*�\��8άd:!p�<0�ٳ�;²��o(m)�\��P�ge�1��#M�Y6�>��9B�RW�o-��}p�����;��췕��>�ӹ9v�c������M��v�sX8��w{�볮��~S���O&LT�EX���iH(���DQu�RI$�bG �1����n�<mۏ���oz���J����*�"�S����ܬy#���DM�D¤�`�#�EVkZ��<t��n޾6�m�z8��M>��(���싐H�<�E��e�+��F*#�T�P�QU$��BB3׬iӷ��q��m����֚{�$�QD�DdHB��\�����LA�U6e�i� r�zƝ��㷯���oz���5�G���QpT�D�z�"	��T��b�����kD$�8��;v�n޾6�m�pq�ܙ3����{"'NA�W�#���
�������jન�i�:v�o_m��=�z�O��О��5."8�b�#��8�����ȖG6E���ç�H2L"F*�̘���(����Lc5�"���p�^�*⢪*�A9=�E�UUc�R⪊��(8�q��Wr.EA�NB.8��QW�#�dO\� ��TU�6S	 �=�PZ~�8�k����>����z�a�Sq�p����r�S��ql��Ӿk�6a���bRJ�N郺hcn4:��0j�����񂵺�k��������Y��{8W��� �q�y{�� w��<�L{�m"c��W-LN�|�4`����1�����.����p~� �vl�s({�1���M����#�\�����|q����ȩ�j;�{�|�N�|�W'*�@�ĽȐ��͏���� t	��}\���D�1c��p���h�"��g��1��=��{�0�c?��ԁ	��fb�b'�D4���qr~�{������0�0�(���9�Ul�rR�=ӻ%��ɿ���(�a$�z���~��A�A-�yJx��7k��-{� U;�EЏ�<���>XIį+w�@x�k�76�� ��5��Ȓ1M�����0��y���ۂ���F�Jw����L͕G:xx�����{'�k����E��������;"���W�����!��짘k���� guK\^�M�(���q��}Sk�:o3SSϠjj�Rx��u�-R��kP�s��SI�fDh�6�'^q�[�;�&=n��)��il�Ju�����# a�3=����X��^�)�S={�a�r�+��1\��~�5�q<�º���k�>�n�D�;<�g3#��撽��W��AZ����)W;�f���>�\84�"��7A���"B�i���f=Q7��L\�OB~tɡ�f�Y�W�s�6=ǲ���}�������pibaNQ%��W6(�]1ʐ�X��;���ڂ�0c����u��5�}����P��* ��Jo��<������o��vk���c^ f��y��ߐ�8>�c��鲻b��ۀ����G\ci�����M׮�Rt��$���1�����̞��L��1e]Y��/m�V��,)ǖ�3�����?��sp�w?��%�;�W�y�V8vR���@$�< ` XggS��#S�}����B�Dk��X���ީޟ	ۃ��e�ȶU��?�J�`$��L,��@��
{]����K�rji'�{�}h��PԈo�@�^�9����@ai����q��Q�����b�놞T���2�nH^����f��zR&�����m�/����O}�O0�,�=����n��8v�I�Jp'{.O�׃��C
��o�)|oPH�\�.��o����(��>�`�!�"���w��^��8��f��r~�m_�yf�� ~��]��p~����\�Aļ�S_���� **�,�y��ֻ���6�6�o�<n<9(}o#��W�c�ì�X-� x�SƀX7���$��.�v�[������kK�lonQ{���S���^@.R\�� 2��da�g���C�3�$�v���iU�?���$�F_ԡ,��%��[�P��R�+�9���c#���?_h;h}�n�O��dV�!��A7@�2�$��M�%�cX��˼9SE�tg�&�!���Ѭ咟m2ƛ���ô�{�����6j��:������w��-���&�Y��m6�ld��6llKM��7d�1m&�bs}�F0`A���hu�Wʩ���r]����u��F�`�`q$
��M~��F��U���P�4�kw�5�	����#[Ŗ���5�f��^l��Joy���m�:XѬ�P�����y�%�@k�B|�����S`�����6�@�70	=�0=���Nu��X׳�]܋��^]#y^��-�flo\5<� {��o~h=����z	Ȟ�Nq���;!dl�q��opsv���o���m��x̆��WW�T��0�Y̑��I���ۙrx�B���&ݦw4 ��
�x:���0ܶ󁣪*�n����.& 憸��y��_
'�@�I��^>х���?��,�'���������&|&�8���}̉}�d^����B<���`e�A�R-�g:'Sڞ^f�m�oQq*� ���.[������;�~~� qo�
~�[z�1~��,��iaa���OiUk�ec3G?���fu�-��<�p%��<�_�<̒�7���۟c�IlT����x��������3�5�Xo��p���������?�>��*���q���Nx�xu��Ϧ�@͏���.�Z4y�{�D��wܱ�ߍ\����%���eY���I]�\�{��~��9|��ҫ��ȧy�����x�$W���x�G*��v������t/���$,�����^���=�;��>n%gUyR��u�����ږŧ�:��:nAr�6�oJ�N�U��� sw{+nJ�@�z�-�o�4�O}�G<��yd�G��M�i��M`��y�D�����#UY�7��[�����4���P\��!/��QV����]^Rgq�13E))뭮^�������ZI��xt�3�g��@v��y�0����>�۾dߥr�N��,y�w9�ŉetOom��z<.j!�=k�\]��k��A�!��z�lo��ݜ�DZ}+�{{}�/��YD�p!�����(��d�%�9�EM�L{�7y����x�O��\��U��Mw�}�6���a ,��- ��;|,�^���ߺ���� ���CN����_z�~H�웻�rǀ�.c���r��*��7�<�n0���֔ Yb�܀�?V�?_�͠7��
��KI(��=6��;�hyc���̰=#���W@c
�Q�fL��F��8�S�n�	���>��*"�U��(P��`z!���%:��x�'ɮ|�O�Q�󹄸�%��e�����3c4_��2Y7�4[@��a�F�����g�<��C�Q�{>$�� �����J|b\mA)k���)O���4�,]��'�:0�C��?�a�Q�� 3�{1��Ȑ!�	��ɥ%k0h�2hfoQG'��X����zGE��t�֪��B�5�p}S�	Fm��Y����.�kO�ұ.���ڣ��m�wǌ�3FB��q[���3���aD6�*��>�*�ng�t7)�j��5����|��<�2a\�H^.z����u�[�^s~�+�_��:��v�Di�ir�2�nS!���}�y�����?���K|�v!�~��;�=>{3��[mG�04�L6���p���׹GN��]�zoBw�<��|2�ǃ6�Ǐ���_P�����9���j��w%� ��`)���ZF���Z�R	M5��9���� W��1�5���O��sa}�D��C�نN.�v>��y�#��y���1�X��7^�c6Bt�\>�D����=<�Y#�s���}�\%{���=��<�חᒀ���|���&���@'�@n�}���� MP �u����\��K0mEj< �oKrq����ɪ_������������xC�.铌��h=�$�	����������CG:	��~i$��w���!,�uw9����[�_�rM�ntes]]�o�u��7�d7Z<:}k��0�����@%v���h�;�aa�a߽�ulr� k2��4a1,�<{6"��s�|��k�<��y��؀�qn�a��*k��<� /�Z���!��IB]�����@T��3vٵ}o�~��4 ����7��x;s��qɦ6S�aT1H	�}��~oPUx�'f�o�b���������3���_��R��;����j��<͝HѾ怊��f0cˠs3������6۽7y�hG��b�C�:o�oY����^�S/3��]ϣ�`W%ݗ(t�V�_p\�w_<7v��F��uN�@�N�����Ij��y|�=硧�h��?�o��� y�ކ!k�!0\�yoK#�Y
�dkʧk���ʚY�I�Y��r�(y,�`��L��H��D����f׌�a�Nn����S.[�Z���VP�nsvs�T>�P1H�
�����|�ɭ��5�99�^�uC���Mq�߿_P�;?{C���L �eT����1�n�u���.!��}�fP�˙p�7Zὢ��.x�l(�����x�ku��a��>�|���3�D�e-�OK%�y�f����D�2�8W�>'hxN��~�����>H��[9�Y�vP��v�uҬ`8;8��Lc�[���/dH�,h�(lgz#�CA�@9 s'Y�ƈ��O���f҆�{������>&fn�@=�ݧ8�͇dg��u��[�<�w�Q�N�08�vR�<��G�&H�����0�n�i��W��L857�����-➱鼚cL�n��(�S�m5�8��3_}�-��;���L���T����0�Zg�wiu���&]ٻ�+\��q�7^�E� P�k�}k`n˾�dȬ��e���ǐ�}�>:�sp�9�LM|�/��ԇLd\3]���)�i�^~1mS�m��s/�V�Pm�8f}�{��ˇ��K�9n�Ρ��x��33�(���������{�u�hZ�	I"]�F�E�ITh�����Zou��Ry���mu�S/������4����ջ����.�p����<"ԬFq�t�I�*�����+�<��M�l]n�$���j�$��o�).��l�>��f�"�01RR�Z���<�2'Ȉ�/���y�;�oɢ��Zk���w�Z����;�t��n='�)2�����w`rzt��[r{�o0�X�]�E/K���\�%�Z���\S�Nj'�\�wҚ��/�EW����C�1�U�L��v�|�[H��Ȧ�O�ӗW&O�x�5�`�1�u!l�w�3p�GL>9��`[x\��qo���uo�>]�'y��-��-t� ����x�x�kW{{��pnbsG�/2�j���C­݈j�>|V���Z��@_�r����Z�Ӿ^Ù@�634����Gm�S��ӈImAԏۀ�<c)�-v-��d�%N�dd@�0Z�M�O˚�ܓ�݌}*��ax�Ք�����*>l�[E�OKa�zm\xw�)�����,���Ň��ȕX���2��0��,u��3�4�X�g2o�o�U����@Gg���̄��� �!Nϻ���7�Hȉ�q���I�0�?�zS	ي�������jIr�|�V/@�w��6����>Ꚋ�(�u��� &6�.��Ph��jl���w�r�H���M{̥�¾�+{�xʐ|<�.�}{^�(��=�2��=��u�TY�`�q��`�����>�sQWK�9��fonj٣�|,� 	�xh�_W�x}�+������?Fד���a�޳aO�6Emc�8��]��6�X���aU�,��of����u����%}C�#�`����T Hhb��C�
�P�M�P ����[zP� 7��ʹ.!� 9��_����{�3q"�
z��qtL�����
N���F�!�[ ����.����lo��>-|��	�e���kH�G�Sx�Ϝ���!D��T��7�9)��v���<�l��᧶+������L'��o���,�0W���ݯ�6�7�̱�!N��?5H���Г�Ƅ��@�&�/�-�
��j\��ˤ|�Y�T��kC���r�]��5�8���8�%@�_H��Bf[�����_�O>7��ܵnd�_�&�o8>��/C��mk>] �c�g=3e��f�R��Qf׽��
�����=g݅��XL��Ζg��]��q_���&��&ϊ?���8hܪ�G|13X��j}�S�O���FlC�Fa�:�D�D���ܞsN�`"�J+���\&Qقz�`�g��2�a���o�gf
�z�it���1w�f�|0�s��psO�6��GZ{�F����ih据���勱߻M�$��q#U�U2l��1�|�:v��}�>2ەX�������*Ӵ�uJ�8g�8�Z�8N���̥��( F�8�.�zƪ��v�r�U���k�j�:0)�zo���+�o�E���٭NV��{CB^>����xa��r��H0Z�0��P]Ehb���j x3t�HN$,�?y<@��r�kO@ٶVN0���`U�:��� i��!����ׅ� `�́s��W���u�ױ]^��uE7o�J���e�k���m�T۠�sRqJY���r-�&S�4�XBH(m�sy�C>\_�N'-��� ��)o,�e7gz�T�<�m�vAt
�h�0SQ�"*�ѩ�� �֤��!�\�E��.[Y"8�>�ucw!�I�׻�w-��D��8�q�<m/����^Gs�$;Et��<�>=@|���$� ���
�&�A�L�p"��=Хa�m�',NE��q�X�	Xq�܅��/��WKSWƹ R�ΫĖ��V�Ҽ=*m�?6X���W.sƷ����$��a|V����<<�V�m"w1T��hl�E��a��o��Qs�n���kd��I�Q7����h��~϶���=[� �s���ء�߳��г�%��dn�����F��ޭ��.[���T/St�1TC.����f���ƄC��\����>`G^���m#��ʌ���k/]��F\���Y���\d��A+M-�uJ�-�����@��u研�ߏ�=v�{�r���g\7[q%�~8�u2�ٗV_m�J��zu]nE���f���>��F(`!	�����QB�*C !Q=���{���r����3Q�k˾瞼�2�@Sa'�����o+�n<=����.��k��O�_�����	j%7ҷ�׾�;[|(��\s��mN�K��'S����R/�%����|���uf}U*�Ѫ&C�|�χ�d�1���.�>~�:�-�ޚ���h��Ec�7V&������T�_�������SO��<�<�b|��߸�S��e��S�1-ᑉ���H�FT\�*�#��l|��]cM�_���]����F��a]X��<����ܕv��inV�#ʞt��@�k�O�8XY�]a��o����x�����H��l_��q��rɐ��=xr���=����Idȫu�%Y�zr�Oe<%�pNj�����,-�W��mC"�êi�b�T�i�7�#�g)�����;���{{"�Ϧ5�8��y��٬�#{_C!��k�OB���A�� �:�vc+ķ�_đ�Y�2�xMx���mV$�s(;�|P%�zRs���X4�ϕ֧|#Ȧ{`gaH>��3�c0�{��x@]�[i���N8d4P�x3�&̑�桦�e(�u�wӊ�Z��:C�Ja���V���v���ծRT�����k�{�
�N�K��E�P�|�����gw%�3�d�ޢTw���r K��)�:�cZ�L���z�o���&���aQ�,K�+`O%ˬH�_u�����Ud�B�0��|�����X
�ɷ%>ɨݏWNP8:���9KM�r��ې�z�J��uB9fP��}}Unj&��5	ocΧ��e�{v5��G��؟<YN�f���P퓻�[_;8֌1�+A����j�e�з4Y�z(Y��:�]�A�5Y�ҙ�o�q�%�L7{uF���\%3u��"��	i�-ڝ{�7W!��h�ǝ�y�Y�P��oT�ր�Y��4;��~�ȗ�x� �b��fGF�fWՃ.�(���}�W��г��K�e��:�v���ns7ϕ�[]zrS�N�#&�cj�猗�*fG�t��8�8^َ���]����0�ݏ9W��	����%���7�𕂤o"�e�8�L��+O�m7[BwOG '�B��Ǡ�u�qU�*��qYW��w������ۗ�cPA��b+��*ڰ�`���w^Bu-aR������D�Y��c1Br�<�Wi�S�,��z��(��Fex�*R5Gb��3�Kڧ�v��#�HEQ��-�j��F�R/,;A)�e�H]*�ʑ��y�ѩ�j>Býn��7y�"���W���~78�;��C�vT�bT��*m<���D����˵l��J0�R��^��n{/���q����>Hƫ�v�v�!HN�Lviq����rd��z�K�9ݻ�Pg���/�\(ݓ-��Af�B���M]���@W��{W����+�]ښղZ�x��������W�C���Ӈ9����C��[|�9�5����St�gV��<h,��6Gr��\�ne��7^�G�f*�l��ɏCi�:�G;���P5�[���ޝaR��9M�W���\q���S[n	�Z#�!M����*p4+�0ӕNu�V�C٤:|>�N�Ko:f�ӭ�E�y��1;x������a�Ӡ��-m�)�9�4$�d��;�_Yb�Ӯs�Y/���{Z,9c�d-����5AY8��vJᙨ�������&anmܤ�)��i�h�}]Գk��&�+��N�h=z�+�J�`�핝�{�S:Q-��u�C�8��Kp���z�wU�Wj�I��w*�ɝƣ�b��BF���=���+e,��*\���5=	��p�W�|L��V(k�q����묎�6�e���iݛ�^��r>^�W��0�R�a�9��tɥ�GyB�L�Q[��[�+l*qғ��t�WS.�%#&���:�=}J�d�g[�w.�z�G��l����t����6-�Pv���jG&�����(��6��ݏV��q8�ŋ���u�l��cM�3]Lf9*��H��*��		��%���ݏ���N9��+*�m�Q�H&�	8CLہ�":eJA)m7&��j�f�ey!i��nh�q��66���(ι]�J�cJ5kĄq2�D�
iM�&U�N�&�t�y�h�S�^s�yyG�&���"s�N�̼&�v�͚���= �!q�	fD�8D�'i,>r���'hGaH����h���NPm�<v���Ǐ�����i��ò�<�UD!�H*8��dA񋜐\X�AJ�a:�$*Q$��t���׏m���c֛�N�R�	.A��8�N�*����<�e& ���$GsP4z�n��z����m���ǬzӃ���jHI$�z�UT�b&1"��Q$�$�C QoXӧ�������m��׬z�޲�fJ�UBI�Qq�-&�1X�A�2(�$��j��BUW�ӧo�x���m�����p;��
�Ȑ���\��Eu��l��*�$�I�*�櫏X����z���m�����=i�vHF{�jC�*�S$:�G 8�
���0�.=�{�\CSƵ�*$HI\qA�"�&z3A�EQ��ʊ�-�"�f\\�E�`�*�ш��O,��\\"�`�[#R��{ĮW� ��f/MTUqV�f"
��d���%s+�td�I�!�f�]�ڎ][�f]�Y��+O&��{�Ceޛ8�/����.�mv������gco��^F����"�3i⸅�X���r�&���m٭����M��\bB��Kl��b�:�XU����`�����"H1P �B�c��]�Vwm�o���l��>k��O�U7?oO�Y��ߓ�8� �{��T��2��������Ot�H쇷��;?d�Gm+g���D:� 3|P�Vyx�"����G���ѩ2H]j�Iޑm�W���? LB|�G&��j���znb�/V��C�=�}f�M�l���F�i��i�NG�zދ��:�5��{��4�>ȅG�݉�߸�g��]�`���E�l쿠g���c�fh9������r<N���8l���L�᤯
�=:F��x|޽o�=n� �~�Q�L�@<��Kr��y|I�o����zo�5��|9�
b��o���>�{�&���.�j������.�B�r�.Лr�A���@��H+�������0�q��c|�`K�3�j[����.�}N���Pod\l�nյ�����|�$-`(ֿ7d��[%���cL�sb���d -���x�����_m�20�L�� �C������g��Y�
�>>G�D
����##%�|������c�y��6�De0{
��g7Bz�W���qY�0��!}��{C����s���JH��Q#伊���}t� ��]�3�������e�<����m��ūS��h��[Sn�-���.�nv~����i�u�M[�.���p�ϓ�]g��y�0�F����M��R˃�w^	VH�鈲������,����#��sO��u^��ٝ�����yＯo	��1�0�0A�Q繞{��ϞW�<s�{�G��9b�еyB��&FTE�;Ϛ�����8��dg�A&�`s�h��;P��1�񉋸���t����%>R�卹3x�qt����i�kR��T�u-���Z7�!r�	���U�#��a���ϽP�PԨ���
V��wmR�����.O}~�B���r�wM͌g�K�0/�@�/Lv��F�ÿ{\�(r��M�3>ťgaOf��a���[0�>2�v~W)��G�FDީ�q���z��y۞�i��>���u������ �\��>�c<���R����)$�|Њ���_~*F��O�Bh|��i��gh��w�6e����Q��/�9�@����}��ަp�y�^+ȃ�}�0�<�A�;�`ṳ*%�x�l(ֽ�OU�wު^�Y:�a{�Z��i}�qqB�X��s�y(5�Q}�+���������'^����}���@���D5�P�y�f^FK�fѯL�pb#��	�L��FU�NBe�i^�����@�`��$��aa�k�]=KǢ4/�q�Ǚ��z(���l�G�Z[U@��©�o;F$OQJ����]:Ʒ�r�=�&�jf�J��ټ�r���%`91�Rܫ{]��-�6ʤN�9�wS��Q�I^gH�*]9���sM�ls����HBD�K��.7���w�,z���G�O5��y�������]�R�A(`) 0`"�Cu �7�ϟ;�|���y���֕g�f�3�F�~�B9��P���r�4c�xh)� ӡ�̀m�/gI���"���75��rMf���T�G�UD6x��2�=����T�ـ���^�C����t����O{�����ÑB~�}y�v�S:x�a�e�~�Y�׼I2-�T;�v�衬�Om�)GOu�^ʸ�s�nU��-{pf{k*!ꅲ~��\�&���|������, ��G�� B0��}�Q�^m,9�^E4��)��H	��\&��������E���c���]t����Wg��G\�p�S�N�p��9���P�p]Ƶ�����v�y��E6��7^�P�>p7@&z})�I�]�G�ڽ����=��"���������Ŭ}��|P�,�<8�}���l����wgr/�����t�Kܟ0�zsPd�;�es�;75���9��ҞoH�F��G�I~ά�(��gPN��u��ݾ1%�r���2�<���/}Y�)��gG�6{FF%��-E?US�/��Y�:�1��|�`\jQA>�˖�`f�f�q���h�7�(���͟���%._�R�SGU��%�$�W�.������/�޽�[�X�z�g-���>!Z·�\C	X�c��mNj��q�]�ػ��`}��fE(�N�,IlV�'kt򵞵c.�Ձp���s�_x �1A �P50��`
� ��y�w�7�S'�>�h����[��� >��������+>Pq>p�wS8��7�"g��k�g���x�԰�[|��X�^|��kS�Wgkѣho7���ѓ�XD�F��0��w��F<���c4�!{��z�	l�W�}ǌ�s���*]k�Dqb�Mu��z�h/����O����oj����x�v�gf��0��zۚ"�kCǟ���7k�&�``i�v�O���������/�q�1 �E�xh%@Wu3 �<1�䳿.a�밻������-p�w��������Bhv"��S����z�&��g;Ek	򏜹Z�/�U\��y]�g�}�z�^뮆|�Y���X�
hah>�;���_Ė:���_����<�w$�bW��v`��k��J-�'�����w}�v>� ���5�#�Ωt듁�vg]�l~b����P�o�YP�ׯ�g�R�	�����o;z(�M�@����CK�t�Ʌ4��Av��K�]kz��Qt���Sx�gt�h>�x���R�������h���So��uL��z��b��P\�z{Ǿ[�鿖(f��U�6��4��e���t��y:��}�����3sN����O������"eU�s��0B�J��)$�ce��^�Ԃ����b��A ﹮()��Cm���뺚�1OP%����:�ᙹW�t.�}]�zȂ��Om����$o.���tt:��ޚ��e�(h���n�r�D�9v�"lt܉�k������XGU�wl�)�4N� ���l��0�X0�U�Af�Uz�J�w��\����h�Re6��s��� Jr��c��9�nc���{a
�Hs�O��Q�niI�N��"b����s��V�t=l:�+�����i
�P�5"�׍���&�^�$���k�X�!U{]1y�1�����1��&e�pj{Uޱ�Ͻ�a�Õｖ4��#�Y�.���^ϓ�y����w�w}>}�Yl�]��3Æg4-��F��M�C�ׄ�S�}���c\���,0�A�kʑ��Xqe�9 ���6z���-��m<���v����yտ*����I�3����]9�M,j��^��s�nN��В�?��֣�~�|;^�ǣL���$�/�E5c�t[�Y;8VK�m��P��˒����y�k�� )�������Y�${y�Ϭ#����:��:  �nV%4�Ùk����.o�#͠��V�����c�EuO����e+���a�t�r��J��~s��梁�Le�PI��_'�Ƥ)0(s�t�����9ϕp�|*����n%�?����Ƴo@��8�v~s
�����ē;k�4$I!�8��;�>3���`VK��	,��>�}�¼�bYL��e?�p����޿�n�9����h�A�VUr~���)�A��'p:s�Y�-�u��lb�r�p*��MO����:G�\PVȜN�fB����ё��O�ؾb�B}�uf��'=�Lه+n��d�p����=�ל���}����b�1�X1  �T�AuJ��w�����ё���W������Ԣ����^�M[�O5\����#'O����W-�.�҅����"*"ϿZ�'/���V�@{�J�Q�Ƕc��t�}�B�ӫ���#���u랐��3݊)h+�q���Ud}K��e�C��>dL��G̯�����`ʪ	��a��@٦�Y@�3x�ןdg�����N'g�S��>�>G�Eӿy�����-�~�;�W�� #\"cy�:<WY���Zq�B�G��j-��T���|���><��Ll_c_K���ʹ���P  ��n�pZ8���tg����^��ϔ�~��A̱^��u�\S�Y\��/�c�=^ř�����#�����p+����@C�������FS	1���}	�5H�EJʆ�4(��(S�*���Y��z,2�]�?�q@�	���'�Z2/V���a�w�Ƹá���jt�^*��V��xj:O��!ݗ���y��G�6V�dÊ�t�mu��9GS�5��g"2o]v+�[��2�4!p�ְH��� ���5�")_)�>�*V��>TP�����G>.���Z��.��ۮ��62~����ɛ]�w��9H`�RCj��{�*���4&�0Ku.=,{ȶ	%k�\��tyd�:�-}OD��Ud�33eo��Kי����KX.��j��_V�+	���9�?p*�`(A��
" L=� 9-�%�<.�dW��+�x��7�gO�Q��@��:@k}�+��E&;F���M�Fen�n�uor"�����}In�  �H��'1��y�<���6��g<���r<G�cm���;��l���;���j~h��?`X1|����I0U:�,�>%�}4�k���S����.l�z��2�P2������'g�*$	��ʇHK���M��鰐/!t��nS�S�[�� FC3F)����Et]qA-4�x�A��<_��H�(�~��k�|�	N��v�5nW�@��ϔϻ�:_e��z�����`�tϐ|�Z�E{<�
�*3�¦t��-l�
\��>1�P�����0�y�-N#ڭ���@L}C.F���s΅�������Vo�-��0�X
�  q�{S�H�3��ɒ��)���D������X�k�A*���}q��� �}���ډRDZ��"�Ƨ��9v���D���`G�Ȭ�@������7�L7'8��*�`ȳ�h�!X�I���e�_Lr�����h���XXܮ+~{J�M^"���׽&���y@d�� >�x�v)U���aش��ݴlZx�g����mr�?P9fu�%���[h���:����ѻ�K���{4J{fa7��f�s-�����͇Y�:҆��w*WR(�K{#���E�gkS,᧖q;��jWv�y�}A~�U�����������D@ddDdA����ruxm<5K��jmBJ�L��x��,nlծ3T_���&8����#1��}�oYʴ=���|@r�9k��Ǟ�kB��»βg,|��;����N;��T����,I��><�q?	{�X�:l�Pi��pz�	��/{�r���=�������̤�|+��|+�7>'�D �B�CxU�6�n��́l�(ML��D`��ӑp`i�lh�� '&1@�����w���ӗ���ﲱ�3m=��^�vz*h� ����r�����{���ց�P�>�WF����(>���C\g8Xw�5{z�o�خ��W|��z�����=��l�Q �~Ѧ9����:}S;3�������@`%�#"$(����lccuV���#kR.�D7��2~�J;0��;�X��҄�� �b$0��2�a��ɖxD�`������[ >�oG����)�G� ׽��Uk�Z_Ù����6-��\�U��Ma��r%]� p�Ol��L[r?Fϳ��H�ȅ���{��w�;޷�Ӏ���������yM|m�i�<ST�a�~N��EU1=��R6�lu��Ce++h;JK��.�],գ��B �1S���ʽ�|�p]o6�R���b����@����*ƚ�g�{�F�ݣ��Ba��a^���if�']�A|�m�˵`��A�������s���u+�T�6�펚�e��[&Gt��\��]���fg��3 fMD1�Q��� �`��a�ˮUvWs�FT���@�pϣvSpA���Z�5��8�����M�>�g����/��@- %�N�\k�Ϟ�h�M�d0��<)��!�j�U����Ƽ��@-��2ݾ'(V�xn^�ы��zW�.g|��&�7H�0��}C�nU����P~O�}^6�ߕi�:�����}ܭ��yd��CA��qq�����tl�Ϥ'��_"�j=z�ۼ�<%�-���2r<���w1���SAH�=um�3>����+�ao�|aӳ��V������{ �X�\ҥ�r��t9�Y'��)>{[�����k����M�/@���y���V��ۋ��"$)aή��%��v���2��]�!��=~Y����zD�h����?D�������E?I9��:���F�C5x��������^Wy]�����xx���뇴1�!���G�����K��ҹw��3Z�]�!iGt�>1R��"���s���}jF��:ۓ�cz=]ѭ�V�`>J"4�f��B���;0��hgQ!}����@���}X�2Ҡd>e8���;o�x�2�6S\�ʹ��s�[�*��]/^��+�|v��U��p�'�q�oD�L��
��UsN�R`�K�	�u&B.]̡�k�%)|2��`.����ěɹ.��I`W�}l���'f�o��k2��\y���T�X0  �F =��0�* �  "Bxz7/7��6�����Q`3�5�V.## ��/<�qw�7���k��w�j�������\WT!V�B.S���}��p�H���'\+�q>;�^�zC�B�`�g�+2��]W���C���k\�!�[��*�Sp��� }���dai_g��|p���8~Bg��?!���}>y>��Ǫ�ڛ���ĬIc틇�f�k�|�mp�y�Ҡ>bz-a(6"Ќ?��|&p!��K+`��2pY^,���x���-��"�>Ͼ��:ݟD��%0����P�"�d�}�[�DW�tZ�Qc#Ә�N��^Q�I�Ҫ?w���i)��,��ο��9�7hϗ';�S�M�U�~\���UA��o�u�%�Vŝ�w�����Μ�X�s��/�Q�g�ˋ|YP�CS.��D��̷Ӽ�G�!�]�*ǋ�_�܆��`9��?����ao�ܪn��I�,��'%����*]�>r�dL�g�S{�&��ڳ����.(2���^^��3�B������ϔ�wR��My�5��z%��qQ�a�C�~��Ͼk�����[��W&s�"���N
��0�Nd�&�n�1��,�hsSӹ��d�i�HQ^7�\.�\Z�2�[���A��CUhFf];{|�)�9�0R���ɖ,��n�r�aK���d�"���3��+*���uqgQ�[�-N�����	���-�Z�]�nX�e��X��Usp`�Mq�'[��]�m%r����E�{���|e�axop��e,���u��W���Vk�0�ň2�9�{���#i������(Z�y�Eۓ�e׭]�7KN5��G�wj�3n���ge���9�0"�K﷍�a'm�r��곰����+���;����,+'
��lI';2)B�e�'���:+���#/u����(�8 y[�-u�7� ���Tj�p���؝�LyMgP��mn������n���n4��#�;|�Y���sn�EڷR��ݝ�k)\&�J,��4vV[
���FS��P�2��a�Wcuu�՗/�1v4G��c�T��l��[K�KV�aX�q<��5yO�0�� mA�r���DH�jB�y/DCn���3rjZ�j��L�GtR�f��v.����J����wfco+a}tR4r��Yu��50j(M������&����	��9� ����|�dv "dO��>Em�e�W�y٠�ݾ���"��O"j�h!Q�u���#j��TV�QG��a��t�P^� ���e�fM�N���_.x(�]w�I�6�+9R�:�z0�6��a���p��c�b�Ʒ7�P{�����7�5�2X�Fts�Ky�\�۬���A"�;f�VpZ���؝���*�u�T��sȝ��+�Y�SX2Z9'r︡e�4���(3�v����w��a�+��И���ҳ��n��B�ݢ��ud0���3�F��޹�.�#@��q��}��&���KM���u����㛏�\&�����{+'{���Ԩ�K	��JU��s�6�mv��P9-S-��MP@���i�(��G����}+�ť�j�N>�k�kw�.t44��a��7�f:�o�V�f�'jj���vlb�;�cʱFҏ`����p�9T�K9#ќ]��L�}f���H���uC%�b�c�kq<O0�Y�؈����}�'A�U�b fܬ�zvwS���\�wg7�l�*�V���O}Nw����dc��Y(��qPpqŌ�Er5(�!E�$x�(+�a��;�&nko��>6�m�=zǭ7�c5)ҩ$[��\UJ�[ny���fw�OdE�����9�s_z�����m�z��ZzvƣnfB�`���Z��"�N��m�[qV�Dp�1�ǬiӶ޽x���m��=zǭ=�HH0���(��W�S�M�b{b�(<����AWs�Zt���Ǐ>6�oG�XǯL�� ������q�TDW=���R�FID�
���g�X����<x��m��=c�;#.���<��NAbk��ETuYĎ:�����]Aq�Ky��e鄑�jn����z�nݶ�Ǐ>6�o���q���$��b�!�b�i�r��q�y��z�qUUcE�#Պ�e9j"b�s�X +!6dMH�ީ�P���D�p��l-6�QUUUB��1�h��A����늶E�;B"c\I�@E���8S"�yb�PP1�9ej��"`��0�N�#���9��y��p��H�L�P�$�ǄeGZ��z�v2֬.v�+7���מ~J���*0b� 0b A��� �|�����y?;DD��l�u������ ��[����9�(X�q^Ƈ=�P�u9���[n���קp��q�� ߜHO��t�2����ma>�[���t��z��]��Z���|��[&��w�2,���:'��^W��\�`���f�J�3��h왬.������~N.�3��}�ё�kG{���'�|�U�ld G�<�{yR��v)��Q�էt�v��K���N���9�f���#}��P�[�22qf���$����p4�y��?��K(ώW�0�Y���!����Bt8���V(K볚��y�h���� 8f�Oxе���]&0!)�l��o.y�]�&a9^��6��W5qk�(��)��w^�+�!�{~���
�������d��3��@��ٙ�EcZzN ��=�~�:yA�ܰľ5�wy!�[wDX�5����y�sО�@��%ѷ�F��9P�����싮�	ڱ�Cw�ͮ�Z��N������P��v�"�"{�3�+ӊ����<xp�ĩ��Ue��cɲ�b��׺�oe�A�Q�Y��Sw�yR�֧W\�	�����̜�?4x�"j�	�gA�u�i��߂5���ݼz�\��{�{����wV3��u�;V�9~��*��` A�,�C��C����f {ހb�x�q�[7��� v�-D}��'�l�b��6��%`ąŪi���-W��yR��f��j@]�dl&5�����r!�ﲆr�b�}�{�?x�����{��D���6(�Z�l�"q����wZ㬀���
�<{�;�t�O����Ȧ4
���ɣ!�Tn�>����.� V;�d��1_q��r��
BS��Fx�جs�{`��n?�@��V�3)���]������-M�L�(k��`ϔϭT���eN@���1��s�}����cz��I�|�3�r�R�u4�ΐjh��^k����f��	��_�F�a>6�QM�5�dH.�-1
l��Dv���,W$n��I}w�%��k���z�_� ��U�""�Y�YZp�ܻ
Z���|Ӟ{�d*�@)���ds���A�	���t ֮��2A�_����+��x��y頋+ş�y�K(��Zm���E�L�o4��k�85d����Y��"�fa!?s�Kǋ���g���̎O�X(ױ��pW	U��w���9��ٿ��[�ks1*��r�b�;[�jlaK;�z����m#�gZZ�s��w�#��w_9T9����F裍v��q���mՑ*��:��QBU%�2�Z���dm�Q*�e)t �rǒ�ErCz��:�Z��p*��-cK�k!��U$G��̺��.��,j�V��w���ؒb����>�EEu�<�7���ҷD��$��ouե���G\t�%0�$�f�n�e٪L ��L3Z-*P�VC�(���g�ȍ�����Ϋ����r�u)�#�(�k��5�a-�~���W��CGGW�G<������C�$Ϗ�o[7@����\��l6��n�kvA:�yk��7��Osd�������e�sς���v�м��[u�>����H��Fu�U[O��&�<��������|�r��k��1�L�z�����T��r
�i�(��ò�6�,'��lw��g��h�f˜3+Ҡ^<�ʃ�y�����%�9W
~r�2�gK�Bu�:��z��09}>�M%M)�������dS�`w��?l{�\:ͣ�#�ev�o{���V�e���=;.�X��ڛ���۠)���
�#l͌�nU��LKG��Ǉzj�ܤbF��%:V�oƈ��q�C㖻�}|~�9=�H��n�YM�L?!^`;LU���Nf*�}��q�NX
�\G|�t�_���,T��(�\��/ߟ�
���N�w�r�A��g�:�<m���7c��/��Xr�+ɦ�r��z���g)接t�����q�6�Z�
^5�#2�Gd�����P����zOxL�ʺ�a�H�tCu�u�Gd/�����v|w�u�ic��J򟮌�٣��9E@w����F}
���E��Wa|����
�K��+�  *j{Lk9������r�j�c+xa��-tT���&6�n�ϛ�3��.�}m�!�o:����.��<=
���b	*b!(b	L�-AE�7s��}�=�7>P�=��f���`$�"F�-~�ty'հN`���,�L �H��!��,��X������N��?.�>o%���)�`�{�����Bئ����W1��.��vOk����6��_�\�O��킫>�O� N5ķ囌r�q�}�fXv���v&1�z��5q����c{�M����ǜ0w�y�W����2ƣ�q��&���:�^ދi��/������� p}}k�\y.�{1�ٛ��ʿ6��/!w��n�H���͸'M}�Nz��#��TTgE�.չ�t8݊��]*����i W�=�u���q��8����1��~���yOs�P���?ahk�觢c9,5�S��y�qM0��[����DÚ�s��t�����3e3�>4�[FN,
�B�'
zɯ5	P�Խ`-��`�.�ŝ�pka~`����y+�ŭd;�f������O�|�J���8a�n�"��?�@�!xc�����>
{RbL�U/���#�V��$�=Eۮ�n�]żtw_]Xa�VRr����Z�;ҳ�����w��!�k��.��÷��]tm���^��Ɛ�����q�b��#�#���f�Ϫш(A��b	"��x �=���=�vb�D�Q�!sw��M��6|W��o��9��N�Y�/yz�c�(���蜽UQDCax�8�o+�I�;��yE��jچ����w��eE��Lz�r;�ڼ�&�n�G��KN�1������=>1[T):Ur0rym�uI�&�a��V��.��?,��%3��v-`!p450�O��QT���C+�C�>J�|3	�����g5��'�z�h����.��k�#��c��I�T|C7�C�>�F���p6\��˹ڻd�@W=�/��j�Ӈ.�tWk�58~E���;�t��*��.�ނ�.q�cXGjhL�ض	��PSw�?���tp�ՙ��\�t�l�0�IO������"^��+�,[�΀<7N�����-n;��*��u��u;y�~��\�znQ�':1�``����	���nz�e���s�;cZ�<ޟj2.�>�΅�=7�p��v��A�ϹI��3f����p5n�r���	���>�l2g⳨sڷ�P{��O�|��H���jµ��6S���ƕȻ�a�bm�S�Δ���F@z]G���
���/�(��z��/f�}Ʌ]	���f)s�����7=��e{��pw�1��o��P�0L\5Xd�Y6�Y��Kh`f�1��رb����t�*A�rC��C)bP�Z���מy��y�������~������
���N!�z�y��{�?�2[g�N�K0�������x9�%���_69�|�o�z�/|��n6n�Kq|i崚⪪y3�M<��;:��~���I��B~!����|�p�����1�;�U�ސx��T�����C�вI���J�,v�<��_������v��=ޢ'!+����D\bz��:��`�4k;�8�7��}/��|s�u���	�+��C��n��N�g�S��/5v9�c<���DR·@�c�Ꮸ3֝��ד:�_�񤮼*�n�uٵ;w�S.�3+e"�Us�zf�3iyNg��?�u����曯)����� �:
������b��g�{�zr��ˈ!�Ck����r��8������o���>�S��P�x�j1��s�VU�3й�L[j&n�Oߧ�� OT7�1~2�PnY��Y�n6ҕ�.�`����X��y=�^�}��R�#�~���+z�/�8lb'������．2�Fڙ�9n��i���@�/������#V0�Q<XU���'�7>�Z���9��0��]P¨#�+�\�q)�//F�Tۨ0]p����*#9��[�H��OGFV�wר�u��������l��d<D�`))��m��$c	
]��+��T��?�gHg�13�&d�(A�b�AY/�/��Q���n�m�9!%���O?�}�C���-ʽ�hm:	�mw���jg���e�pE�n���N^Ko�_D7!fw�M^��}W'�ϭ�� ����5@�,��n��d��gwt�ja���^i�P�ZgM Պe�nW�Xޜi�j�jg �F+�֝%��^�G��ؑ�@x���,?yW~�L5��w��)`�k�����??~����o�}�y��,�$���I���#]�p@�����������<�AX7�TjOս���)��?��7�s�1�i"|ØI��u������\���=򖉿��][`�M,��x�o\��6|�?j9�ToV�I>���L�gǷZ����]a�t̶�=�G�];�u��X�4-$�?j�	Ѿ�~U���LLF޺�z~�w�㌯���3%L��l6B0c�MN�m�Y<���\��Ѯ��g�|W˼�M��>��dw|�39~*��c*�����@r�Wz��(��^�eP���3 ����8�޺�û�z������@Q�����`�GU�4����ϑыl���L��vI�$F��3qP�/*{q��f(���}�L�e>��g��Z�s2_!�L�{���c�I���V��1eֲ�<�}�k��׷���3�҄A������)C("��Ĩ�����&w���7���w��@�iY�19a��/����0%����n��UM1p�8ש��_���1�5W�����RɆ��}~��i���A>@h4l��C|�f��}��=����l�{�a�Y���r�����o����^}�4����~;���;�������]�ƙ���gι棌 "��>e�A4�9CnL��s	��E�ݛn}J'޺W�]��W�2��H��Vv�{@
��c��l�'���%vX����>�c����w�}&�%��& ӕ\�	�.}9��9�������[�O��[#�J�X)*k���˻�tФWB�cF*N���'ݷ��Y���Pf��a�:�|k��2+G8�ا����d��������^箘{N��9�H&{̃Q䨲/�E����>��-��D�y�8�UQ:�="�}N�^s`w�"X��B�(Aw� a}oՏ�-�=rK�xK�Z]#9�J�p�����꜅g(cdz=�m	���h�ͮv�$��L���>^'��"[
�_��W71��JU�.�w
��r�}D�,\[���(b7/���H
�cB�r�lD"#����}�5t��(�����w3E��5�Ĕ՜�,�����S���Ĺst�-���o��<y�?��`Ĩ�C �v���8�*u��y�Hl`���"�}^�����}�L���Z"�����&Ts��Í�@��0����L�1s�p��+�DF��ʅ��H�9�w�<cC�?�gP5�n1���ɵ�7��肓��Ǜ�P����w��B͝�vڗh�L�/B�Mf7L7n'��\e�/�~����ݮ�#t�|����1���r,�D?�c�;Vt�ۦ����y������I4h��%q6�i���i�������jpO��{��F:��6�h�p�7�^k�Y����|��w�K{��m�9�%��Zy��3�Klu��^y��;���#<�?�f�>'ƇN�û�Ў{#0�Í��p�� L[���ʤ�al������i�%��닗�[�0�����k�v���z�YSmY,"}���a��y�}���\�,���D_�)Wt3k;����6Rګ\Y�{�j��.*;�D�a�}oI�G�r|(L3K;h��	��`B}�Xڣ���ޞ�(<h��:�
\삼B��`�Z�'�o���x�}!Ce��-��6l_o��)��<$�."��*sh�<`��Fc��t� �O�#����%�yDO��E	��*㻥�J�;���J�4�O*&�h�(0r�,B�EM��s�39.��i}�L��wB~�C�43�5C�� `�)��
�.��������9sϜ�N���H�(p��Y˄>U��o�7��6
{�Q�`�g�r�M/HI�:\Z|�yf!u�N?t���K�s2|!<LQyX���O7������|[{ʹ^w�ٕ��Lĵ7���Cr�t��#�"���-���x��P���`�\�Ӽl,��C�yN�6Z-�L|�K�ʏU�����鰺���<�yMjz�k9�lq�7�D39ڞt�NO��H���Z����!f��c��>�b����
Xp�3+Y�f��׌��_M�c�\�?0�ǳ�{���ߗH�U!�߼<_�qv��Y+�֒'ys$h��Of�5��HX����\�%.���1�y�r��{��. +ܪ͝��X��>���� Š�Xc~�m{�H���{�'	�a~4c��/���d��B�t��3A�8��56ُ,B�-/��>65	�{W�p���jj��ą2�����pO=�M�W3��;��.�ӕ�q��'L�x�WB�+��@{���/5p����v��O�V5RUB�ؤ#�_Wqko��{�ڶ�pn��YF֧b��D�5�G|��T0�חv%��n��o�}:����J�f�%{K�u��5��n��=�R@�j^��P�k�Q��r�{J�v�ڂ֞����xd|���<��{oJ��[�9}�/�j'Dk���puR�m����+c g:1J���RSu��n�?l�ز{�fe�W+�[�QWB��P�Z�6�p[%1�u���՚9���ə�)@orm��k9D�6���N�r8_y�qF���)v޼�Z�ϐ��[�޹0�ǝ2������Um����dT��tMl�Ҩ�����kN�_�
��G!v�Ǆ�٫t�.Ug��5J�N��;�H6[YpKJ�����L�1�A����vݞ�:f��t������k��F�o`��]�*���^��D7V�Vu�ٶ(AZ�|թP[㵅'}�Ҕ�WI�HL9�j0_y�s��Y�vh1؅��{{���J�%Y��4f��y�y@d,�L*[���r+/���|v���O\��um
l�MW�O�/� �ri���W�T�"���/(�����'
�邎KBל�^�'zﯞ��;�����zS���$OW#��Sf:F#DNu.�4����\D�A�i��JF��� ��ψ%���.�TEJG����SR&��jOF�����g��.�6��W0ز��	]Q=�\\�:{s�����,��s#�G�#$� ��Kh�0�"[y��L+֑2X+t�6�x��G�Z��*ޙ;Rag�$��5w7�h��2�S{��)���j�7B����gS�]%$k��f[�����k�{
g�r�a;)27��Ƴ)�6��rZ����,��;١\�״�!��Ր^J�yQ��u�'w���	��r�6����@��EvP�ä�vW6��]��� sco���UQŘ���;���-�W�5r��mZPv;ل�X���焆���ť���+�;Z�ʕa֋��u+Y=S��79.����K�e"��ts;�D���1��1���!�n��ͤ�W/��\tՊ͡�M;6�T�g��2i%rq/�L����犬�]�[�����M��:�|rQ���=T�\*��*]��.�����#z�g�0��t�kb��;b³]��y��u_;Ph����uҫ4����f�N��jV����8H�#���bYݬݢ�Ύ�	��Ў�����g����ZC$�R��Q����`p�KVmdͧ��t�++M�;p�;�Avu�[�9P�ݵ���%�����B��B����`�v���.����g��]-`���ee�T�8.*��ݮ���l,�)��H2I�%:�9�N[��E�k��ҍ�M�A���c��0��D�$��%��o)N(��I��o��yy�3|�ׇ�m�����-X��G$H$�M�J�&�,��n78JN�l�E+�,Z,#�H�&����+3v��t�6�M�]�6�!M�dw�8k�,��M�n]��eT�$�"*��j��q�C(-L<�Hra�W�
�b�ڎc�#��"(T#d;3��L���x���Ǐ���=z�:����N�
	'��Bȼ���.�}2"�^J���w�v�J�$�����u�cN�8���Ǐm�z��p�5�qq�D~I܈"ئA�1��+��p�dKg�D��ޝ�Mn�=cN�����Ǐm�q���Uf�d;�)��$�s�|��I�칉X���V����w[�Z�۷o�_<x���G�X��}�#>�*��n¸�"����'�P[ ��J���2��]j	4=c�N�z���Ǐ���z�s�s�rB���ɭ����e�����+R&�\]g!�N1�O�|x�����}z�9�� 9������������Y	�`HjT:ry""-�&�sQQP�!�9���v͕ʫԜ��lEX��A�X�r٭Q[0���a�E�U�H�b��ʕ�W�ۅآ8�"�c����	�'���[kǖ
��m�1���Oe��b�'IR�")���)���jn��K��Y�]Ivh����n��9Go���k��c�����kz�c�in�7W�O���Jp}�k�;�劅M�����thл6Ni �Y5�ݑ��V��-Yd�u�,SG�V촍8�h�C�f	����"P� �H0=!���'�$�@���u`��x�J�l6�s��Z�(����ꯐ���zO t\b����weC�������ي]�'cb�ʢ�`U�:`aZj�6>!���3O	�}ڂU��\/��Un^��":&�3_�c)cH�l{ �,��V���&�(V}9�;)�Hb�u�Vd����pF�/#K��>�H{_1����|�a�`��_��ǌ�U�Ȟ�;K�J=)��^A��(�~�L�5�/��z�Q���ߎ0�>Q��c0�y`�m]�R�1o�;sA]2��<!�R��>�|l�f q�FT�_�;*��מ����v��B�7S0r#�@�^��:j��ցY�M��^���\�07��;�wJ��<�ݴ�:,�W�!�܁�σ�P����|�����b{��SX�ۺղC�/+O���R �o��W�+p�8�	������������m@����ᶛl�;Ƣuh�}/;��lsWD@Fp�$�Wn�d���W�]��d{���|�PH�=�Z�Mڌ�{S�1#�u|Ӝ۽| �6����sW.��&�Κ�IA�#{Ggy��{�<��v�T�e���,��2Cǉ��Y�,��a�oFfE�#�/�^���|��/��g�a����&�}�	$$b$��g�>|�R�_$�����<�P�#��џl� �"�z�K��� N�8o��&|��oq|�|�yD������x���8�����g� ���.*��cy٨�kR׀�����|�˯�.�bp	�N�|$�����goB��G����G)��K��w=�bʼ�c9j#}'�����}k���U;��	��yP��� '� ���!�+Lu��t�����/*����X��Tx���
D���0�4$�<�?��ه�fL̦�p�\�.x�ի_Qk�\�_��B�4�%W�}��a��;gS4y��]��ń�?{Қ���^wR#�<$�$xR�RK�G�s�ܟuX�o�O��KBʶ�U7/����v�����ء�љ��*v����v^0�+��5	��j�����'�	��vGQ���x��2z�!�)�a��|�2�`A�,�Ř8��5wC�z�g�e�=s�'Z�kϼS���`8�%ܡ�Y�w����*�G氌-���A��<1�=���|؟��8���tɐ��� �KDA�]ޢm�ց9j%���MwV��ӏY�����2�)�/6�֒n����aW�g�����zp�-��u
���ztY+�����Q��-(����3bI�/����Ʋ��-��A�=��b��A�	,TQ�=��ξ�_{��[��Cc��<��F�ԝp����X�هx���<��-�c-����YX�������w���D��;�0�À��Y�>{�^?���V+c��/��� S*qޘ�|�.wO�Y��o��X*���>)�2�}��7Tz���s�͐g��:g��]��+犜����X�J�~��8<�][�z����t�.~�r��)q�e��oiT
��� ���)�x��6�U����3[�xcjs���*0���1�>h�c_�����^��H'��lb��!���_3r@��9y�B�s��L�:?�W&��W�N?��L�V��e
����e���1��=G����q�$n�A5�%�Z�TM}C�|+��(�{�z���y���:V�L��c�>���ش���.O�>�����V�w��GX%�]E����g�M��c�~�=3�{�a�_:N:'�E����}.hoe**�Pbۆ5�d[{x������UL*G�wW����ҫ��G8D�Η�v��v�T9��8��va;��b^5����t�]3�Л�.�;���N�+/Fn.c�n����\���^�HY���ܩ���k������P��)$�0GD�o���ϟ	���;�t�Ʋ }a�¼)�'�c1G�H�ˏ5��W�(r��y�\���	v��'�9xVFzd&�p�kʝ�>�2o4��c��^���{��z��Z�dϒƧ��v����.+��v��:qD�Q7	eĝS�Tg��g�=�k�cF�>D��l�8�n�`_|���^+�rӊ5�>-<�wS¦+�z�2œ�����yM�@{�-�2�� e�ǈ��<�@��
��$t�n�爵���,(�7*c=L�x�����Ѳ���(�!��r�n�v0Ԥe����S�20�rDϷ�hMd�79�;q���析/��'�:p���1�|5�8�J�s��k�8�<C�<47(����R,k�����zAҷ<|��S\�\#ֈ�C뮕0^&DsE^�����}�"��#�@t�Ә	!}�Ȁ�F/|��������}.q�w��Icik��xx �����>h"OyOԬ4bH�g;N��b��3R�Vj+}]��WԳ��?sծ�&��������#ˁ/��2L������e�K�R鎾�X�ڥ�����;W�ҜZ�f�p��:-�Z$�ku���ٟV7B4�N�ۺ�q�iP"m�#i���sɊ����c+^����{-Z=\3`v+�z��V�M.�42%����j,"��Q|�ƒd��P˰���ݏ�^0��&'�gb�i��bh8��a�����w�n�h�M���Ϧ�%�ǂ�8���r�&�����ȁ�����I�T�Ucҳۈ���/z׶X��m�}�m�3����A^���"���x&P?��Fcq��g�3~�%��t�xl].����;z��ϧ�<�p��/^@%��rD�|��w�3\2�w�%��g-��G|��o]�_Q��w^p�v�[�4�e�,gQ5�XW�}w���	]
 z'�X�3:דi�C����}fj���p�����x�7:��Ǉ.�!Ҽ�Z�Ȍ*oN�a�sr ��v���Ӻ�f4��[�L%�4K�#����M��R]Y���U�Ƌf�m�_M2���]ߐ�{K<�T@|�~�p��1�C�0�a��1
����bg��wA/@�'}U��g�?Z���8y�p�������Q=s3���WP,~Ye���"m(0h�av�2��u5���&��9�̡�^o͖�(ƶ����#a��M�]���ɽ#fd�xJ��ɳlt�lّ-KcN\?|����x61s���:�ϋ#6��v�?�����_:��c����1�N�����X/+�{	���
WfU�6�o.�Y\c+���0c�[G�������c�����z�3w�8w3I#�C�x���:�S�9�ά�������d
�`U	D�4�:�N�{�W0����}
��c??�TS��Qg
��ܮ��|��-��K[�u�:��g�&0���JY$�!����b�K����s�ꮯr�6z��� ��"�}���-ƲcX[d�7��]��޳�W��~��cG�T<e�~L����`��,vw�j|���T���eMEdmj"�d0�@ׯ���~�{x���<��ΔM��o�0К��:���B-׋�7}��Po,q��!F���� �� �U릙�@�Xp�Θ�cv��+.��S�&1������h�͙�Cɂ�4��Pz�E��]�q���v`d�P�'{�W��+V(�|M{���:�A_ܞ�\�W9(�E���Ӓ����T�f��o3�m
,�c�R�*����{���4x\��C�U0��ќ��p���ϼr�8��n�w�v��w\�������Նm��@P����8�G�z�W�|]��M޶`v�n�n�� �����~�nw�f���<L����ow�o!�p��� �7]��b���]��l�I:;�q��ռ�n�]F��������z�Pו�ࡅX�]���ӽC`����eAv �I��No5t����Jy�p5g9���q�p�b�7gG�U8X�ٴ�ǳ3-��^�?�������Ph``��HR�|�}��ϓ�7�=_��P��^d���62�����>��Z�>ԁD"�z�d|7v1���R�rz�//Fzn;˴��Č�kxr}���M���4�
kŔ��l=P���%�
(�a�2��#Y3��Bj].�Q�u���te���<�S��.l�D�e�]��Uo΀o2�ڍvq$���ٍ|s|��v��\�ϛP�1��ޱ�� ç�����5�-�S�/������m�n��A��ZVC��ig�گ���~��ɹ�[SZWL�`�}d��#�>ޜ���&1�F�ļ�la1`!��j��XKE�]��ۇF��,0U�<3�������Zf���� ��c�A9�{�͑��X���Z�I�HFF�z^*��/�^=<r�X�G�H�^�<�%sV^�Yo�Wh�oo�?=�!����!�=1��1c����W:Y�sV��HD��b��mm�@�ۨ����,M�ʖ�2��ƞ��@��HF�����h�Y�.A�=u�����q���V��Ԭ�{�M��e�'3�U׏�ĳ6����TF@OQ�n��	dV�յ
�3q�U����/!��z�I��"��sVjͱ�Y˝g.��9�����0�Ŗ���W��.�45��%��'��}��oz�wݮ�/��g�s}�a����R�,i��^��y���揘O��86n)Q{W(�O�ְ�^�}ȫ��l�g�l
�=.��u��6���������9�}٭,�M��V�|�O�Jn�@�y�g��<�B4����=�Ɔ�M1��J2A����J�G�������<�:��޸ז�U���?��li����2�4�7�מ��#S�Ռ�?�1�>nw���Eg�L�T��0����mI�V����ښ��o0&�i�Z�G84��ב/`���r7.�^Q�2C Jg��=%�Eê�L]�%��aSmP�}p457�~��}/���G>S�[?SM��x��Ez<��J����0g���8��?mEq���(�;����́�(L9�b[�[���5ͭ`,z/�b�r��n�T�p��y�����^��3=�=x�|�lfKP+�՝W˩���<�_åF0͏F7-x��f�Z���!���L\��l�@�W���-�jz"���=���ך��I*�ʹ>u����ǧ�q�q�r�v�#�!�6���ڿ[1��>�C\v����Y������z.8=[8R��c�wt��춵�Efˮ̥�聡E����:�\�Қe��%�WM�p3����M��VvugVU����{'��#vj��ֺ��F�W�V���/�����6�s��f�B
ʀ�a��CrNR	�%�*Q�F7v$�9*X��^M���󚯯�F�R�41 ��+�P�G>{w{��d`�u2閁)�Cy�W��cSԻz\"2y�#
�t60QA�} ��^XY�>-�"A�����~*� ׵�,/�.�?��4��r��;$���)�>�Eb���^�Մ��]��WF� �JD�[�3��]�F����>:	�� �ge�:�
6�U޻����U���/]'�G�����b�2�W��+��_:N�'�b$��+��QɥOMa﮻�>s�R�OO�4?�+��@-X���L�Րfo���a�%Q��3(���}=����/��a`��n��
�n�o�wp'-����fv���x�)`!��v!K�������E��a1��3�{T��H�s�N�%>��\�2���:_i�h��W�oһ@1�'
��ѯ�O��Y�5c=UҺk�8~�5K6�I�x�!:n�ʠ}�?���6�Q?y@��&���T>p��]c Ŝ�|~i�~��¥�5�mj���־t,g��l��*��?z>�H�6y����4;r����������WY��0�K_v0��>�S�r{փN�`��
hإ��	�J�6K�ь�\�Z���|U��1N�N��U[.��s�K�]����� (��N"4웛�����o�,~<#�4<�0�`y�x���j]O�K��y�L({�'�����m�Z�k�����|�������!��!�4�j�̼Υl��	��c���a��I��(>�o����P�w�T
��ߨ2�33��A��Mю[��g{��u��9��^c�E��`�_�=���viQ{˃�A}���;�Ƞ%�R%�tk��$�9�v�ENga{k���5���r΅ �g�GFH�HL��b)K�Q.��
5ߟǵo�~�Y��Y��dWu��N����S�7�R$k�F<c��!����9T���C�Z�{P*ܶ���:	)��s��=!�IK�$JH�G�~�Z^��'�OPަt�(=�z��Έ�_ˁ����'3r�䐇XԗOy��"�/5s/;����}]���'!D�?�"���?�)7]�8��NB�R��'�c���+:���v��&0���لNr=T8�I[c�,yJsv���{*�7�v� φZ���Oݱ�9�h�.lr�5�wzA��^����5��je����]2�g4fX�W�G`�Ծ������r[�Uu�-�B����-��k�y�$��9u��X��ۢc��Պ�b�i�
SX+R<�WqTnSЕ��T���̊�ګ��-���L�4`���:sOn�#�����g�]���d�qb6�4,��ʋ==l�-��
f��E~g0�z`LC׷�?y���L��c�ёV�s_3y�.��Pv2���y�",�0���KO7̈́K�5�e#�Z����G��6��T�\��S��:�yҮ�C�^,�9Ûwh��[�5�\cqR�+Vc+}Z �yj�}.
Pv�}�IM��2c��rM9�Kps�Lٻ}]e3���i��s�ⷎ���FÜ�]Լ�|��	��!�3n��LkO��r�p�+[䭥�x�,;Gd�T:��hI�ү�])�rê�5�z���9\��ɯ��b��5���f����f>+g���#/tĲeT�u��}��Ӫ:�x���N�`�+#���;ɭ����ڵ��Ջ���)h=��o7�R�x�\lo����n;�a�D�땼
[{w{�	W˄�OǭT�M�W��CM��ԯ|\
��{�[>���O�˽$U�#����:	&V�@��a�i�KN�z�z{룚�q���Ep��O*II(N�VT�Ą�U[	d�2
E^/�R�NL�"���︩6�}�����%��lz����R�DD���ɨ,^P�}�^W�N�;��KKQ�k�x"���t*�*v`#�/k�M�ֱ�k0V:��R�t#���m�qw����'+Ȉu��k����&��%p �Wn�zU��d���ЂQ̍�̻��0�k:���pC����2s��l�	�ed���A��+T1���\�g-Ļ��[wGk�V*m����+�W���k
��l���I��V̪�nQ��)��)zoҹQ�f�;��=]2�Z��5���T�m�C�ةZ�S���C�k��7A�|vB�OduG1�_^�C�Ԫ����Ok��	Kjc
p�t�Y+��5,�$Լy��\h	�s�Hg�����\;��]��h�LT�,ݛW;.��Yꛓ{�IR�`��"�\|�'3owh��&U�.Mk[n�<f]�9V�hε���t��&f�,pQw��L��5].`�x�]k����{B��=��Tq����q���$ػ�)4eP�9�"^�G.'$�;u�):�mK˼�k&\Ջ'�lA�{�N�\�f�+��3�{�{�-�/'}�z�Au�*b�ヰ��
�X9�	X�q��e
l��3��I�M�Ų2����v��^<x���z�9�}�r5(�O��:C�H�NJ�R��Ǎ�@D�3v��9����>�<x���o�׬c�=�A��� ��΢��J�%*�2A��Q��o��N0i��޾�x����ގ=crrQ#2�)$�Y���a��Eȓ�i���M�8��Oz���Ǐ}����VA>a$�5��S�˓��Dy22L�A�-H����c��X�i�Ǐ_^<x���oG����"�����]"��*��=�͎Z.P��(	�jT�w.)�pi���_<x���o�׬c���20Ez�ff�ɑrI$q�8�#$jX��dTh�R��ٛ�q��H� ��́�mT���2|�1VLb,�
�u���Tr�*�2b��ͷ�l=�."b���\��5��ș$	�"̏��=J�8�S#��2�	�ɱm�"D�GNvC'{�1��c3��������>l0����T:����? G�HQPP�Tv��9����k������Y�:P�_���տڪS�R��Wޜ`,���ZS�;6F�����y4��y��bU%��+)_�K�o]����%pQ���+�)����B&*{��=o�$��n�3�z�ŷ�������y���g/w����7����	�Ie�<vU�ݒ��M�������w�����0pe��ﾫ��G�J.���\q��f��U0���6:!�Nef��͑�,0���LB�6o��b��T�}�!B������yړ�#G(�0gՂv��'��S�?�i�9\n�0���;�Eí����_���Us��S�j��k\`7�rz���l�	�+8�c��$�P2���\�C �¬=��>s�U��$��f�g+��
k�Z�`ϡ=�[M"J�c�[N5�NX|w�@��Trqpj�Y@�ǆE�P��E��N�R`��s5�]5b�Ύ��Z�y(,W<{D�_�fõ��{!��`��$ �z��Vr՗X��.鞷���i��i�`�=�������OsU�R� L��%q�0u����l���ػ�%�=V���
�����B-�
m�8�h�m�u����:ft�ڀ�4:�*�}:�����jZ�����9�����s�S�a}Z����ң�1^��*��w��t���Z�޼�^�wW6B��0A�T2�hj�d�0��~��g���{CK�qza�W�5[����¢���v���ޫa�E6����wf�����U�y��ߠ���K��/E.�寙�<9�Vz��늅Gڿ���yh9�������ȅ�E����o��>L-��|��[&���s���Y����V��[���QT����a����'U%w;8"?k�w>�B6w��p�4h桾2k~Qm�s�**�i3��R����zjwz���	9�g�c�~uJ��y�a�=X�vB.L�����=���q�۾�}�PfKhNls��l7ΰ|󆚰7���g\�8)8���vU��^�ӡ�8�T�Q�k��`�l��l����:��q��a�gwW`י�3�<0�-��-m�`n��;�N>k�|^�
b1��:�VP4
U��7!�0ں�ڕ�uvw�2(4Sz2���5��&p�;��O54�Fy��/���A��R�t�w}��w7��8�N$�v_Ķy�a趸p����~y�E��cK��0F[!2�wҼ���V������v8\ތ:����.�cV�S:.���.x�Ӕ*���8勷D�X'l(�p�0�)��n�m��iV_k�X�h�r�7:���Z��/�]�x�;]��7U�:H�ً��n�Y��e�Wiؚ-ly�PCM#wvmM����+br�hÎ�����ꎶ�"��g�ɉ�c!���}�z`IM���Շc���a��$}���7�ϯn�y޳Ǥ,VՖ"��.w���hϖy[������~�7W����7��Z��1��r�(��T�@��xa��JM��g���X"~�ʌk�Qm$0.cN;so:V2�t)\�ԧXW;����8�2���K4?;�ly�Z���W�Sy2n,��]ìk��\��yl;C�F���'\UǺJr�n(��#�Ӎ^�f�#��"�}���Y�-2����g����c��C'����JE�G'�o3ćx�Ҥ&̥݁�N�`�ܮ�"0�i�K�@{�V�����	�mj�-"c6?&q���D��.%�M�F�:�A�5�"gdHT��{�6�G�5Z���������J1�t�gP���UFG�W� g=����޹	���YM����?Nų�����h��D�I������f�4�D�I<Z[	.,������R���7��[x�l�|�[��U]D��uҼH󗌸13[\��Tc�Ϛ[($R'wuN-�[��|	�����<�͇5~��:L*t�S:m��3'4��CRُ�*J��5ժ��g6�f+�������:���s.Ծ<�쥮�;r��_|PzPUw]c�x�,�$f�rj���5eysܽ�W�}O��hbA��������<�A��������d�G�陆��uN"g�,��g�/q�𻖓/$�	�������;�,��f����Cr;�tU��s���y����c�]����3����[�;� u'�/���}^��M��[���3�/����+/9k�T��-�s�kAX}������O������֋Z���À#�־��ْ\W��շ�®y�-�j�v���s*�q���] ��s�oJĖ�F��=������&p���wwM��-0�
A$>��c�ܫ��گ@�˔�fI*�Y�/���p1z��Gg6�fg�u��h��L&E-2(��E]ͅ,�4A��<��Y�o'o^`v�����y�"D�a�J�g̩������٫���~����ڿ���b� ]�R��V�q%��:7w�z.fD/��ѹ�`D��Uդ�`��oT`�f%Y
wVǶmw�H
�А�G�Eu�)�3�{����LQ��j��(�gfҫ�]��	N���u�6���d�F[�$��,=������y��1�����Wr�9W���ޝy��fy�5�m�ͼ�0�+�����^>�~�~ţn�לch�����fy���ͣ1��k��F��4��7F�{>	��X�g��s;�z�mX5�"�`�;O�R��h�ti�^̰�`��,�-^����y�N!�6�0�3��8�lғ�}�/F���߀�=�x����HGcKOK�D;�n��k�7kx�Ό�m����~v��-��C����}�ﯬOy��o�-���"�7N����^�c8�OzZ�76e�Kf������C�X�R�a�	D��ިu�,|�$�I��'`�5$om~Z9�i���a���X�A��1������9j���R�γ���\_�)�Ֆ�U՝,\���ˁ0�D���K���Wd����c���@�/�q��d\��&j윌�x�}�w	��|��䦮��ƻ����0��+�����P�k)�U�ʳ�-�gm��.Oj�Κ��y2�0i�0��nK�o�Z�c��7�(�y��^�u����X4T��(a+��Y�N�ק��ec7ۢ����n���W�����S�s��������N����M`1������|^oL-�1I;�c���~>f����o��H7�$.��lᆻ��|^4��C�=���k2�zĀר�]���2ѐ�α_ki#���[җ�Y��y��=u�y.�����H.x;́�Y�Z�d�z0���i� �+�f��+�q�0z����w��y�?w0�@q�3zc}�|�ٜ|ˏ.��vK��hy��g�������΀��r�>^���QB�
���ow�;�爯T����К��w[W#-�Ѩ�S e۾�/3�"h�|-��M�dP5��K�M�.v���q�s��7���6�g�j�Jx����/���5�;�^Z�ǭ�^6�k������mצ�3��X���>f�)����5d�Yڳ���]�$��x)iXɮnU�$��0͝k�	UQ(v�N�p��?/�}�bBB�.����-YTE���n���;��V���;+������P�N�|5:�r�n�%���8�4�4�J�a��D+��nqd*Zs��8n뒲��6~3��!I28@�g����R�=����b`�[|d�NQX�U_���wn=�w˛�ROϡ�����C��9���nwǧ�&���O1������qF獀d�{gf�1460��k��wH-�'�˹-ɻa!'��\����\���Х�iq�Ww�����]t��᭞����o���	�zJ%|�O
cgժ�վ�Rz�Ä�}���ݕ܀R�𙨾��h��w���8>��ssh�Ne� N^��Gd]Ϝf��ڻ}��W��q^X�=>n��4�fԎaѭ�s�W�m���w`O���čiW��0�曙���mMM5��?Nq�v���\wwX�����O{�Ĥw�6b�q���D
(�a�>�����;�"!��-��d�kzb5LW�K��S��ΘS�A���4ܛ8�'���6v9%T��<��qa�#�T��[��%��\�t���_}�PWẼ���ۺ/���F���:۪ܳr�T��u�n4�Z�^��#����u����2����<���N��_��t�eV˻���7�u�v�՘�y3d[j�3��|��Y��2ڦ7�}��{#�q��\��������>�t�k0"ػe�>�F:����2� =f�oL�eS��;����� �Z�8�T��~�%���r	M��ȸ�]�c���GAQw>�Jd6x���b�Η2w����[ KD郯�\�\`ɖ��5<Vyu�WLީ�b�᎕��-p�L��c��_�~��� �=>l����S�c��d��G$7_��q��h\.ӡx�3)�
^���9c�C^��58l2�t�t��A�N����5{��kc3;	�OQ5h��s6�������[��3R�^�Hf�*�y0��S��$�����k�Ԏ�2�Z�
��Y�u��je�ܖ<�z&o�����K��7��y�{Q;��&ԅ������ �\5O���,��1��=�*ޙٓ�qZF��ݥ�+[��$k��&z7���d����_�����[S�mf�$��Se&\��oT]3j��o�YS�TW�+|�d�0;�����;�.�4R*�-��{b��O*���'Y��emu61��BEb�.S���"��;���~�e8A�f�<�χʚϳ�:���Z��V�&�W��G��V�^�_o>D	|�-��;L҅	[?�r�^��S��[��u2f�久��vkYw��������@�9#s.q�3��~3sR�U�/:Y�����u�ͪ��z�j�N� 3f������Z��C{+�����V�-��4v��o~����\	G9\�/���[�^���luv�{�v��h�@��:��rc�.���C���{�د8�ֻ3�O�}���oKz
���I.�Q��gM\w��i�K;�D�h��`��Y-�2Y�=�,�f��}���V;K[6�7~�Ӣ�d�``7��*�-}B����ÆH���]f��ɀ�b}ӻN_��T<fz_:<��hM]́Wv(��;Q[���q'5��+��/S�6�~�}g�/i��a{X�:���}���jށ��|�2��>c\���X"�P�Ѯ܎iZ6���{�	X������U��"���D8�0�ͨ���N}�Ge����bu�`}�Tp�68>�x��ˢ/��XK��`�������5�5��{�o3�|��W�5L��$�羱���I�,����x�r����o���c�q|�w�m�WG1��A�o���cA�&̔�� �v&-����ZM�tx�i.T\�$�أ�{N��{[����! Rg�T�$���|�����{��[�ޓt��P�PR�OR}�ܡ�Q�yή��8�Z�cyZ�;���*�ӧ[�}қۏ#M��==eb���dh;m��uӶ=��;CQ��f��x[��joH�`;S��^)�z�{�
c#N삫ŋ�W�&���9͕<�3�9�ɸ=\w��-i�>]E7�w�z#X�97#q��?e����~c�8k؛��k7����c�g�W�4�M_.̜��Ɔ�5�%�7��vh����Y{-OT����].˃!�t�[Ⲡ��������j���gD�u1��#����2��z��Yk2]����9�^����Kv ����v�m��Fl}�e�x�g&�cz�����٘�s���q�&[dۋ�;�u��{�#�׵t�t�N�h8�g+8i�Xj�ri�Nv���	��j#�w����%��7p��6�#U�ު�"��XfiS:����v�[C���`ʺ���a9F��q�Rg��j���HT	
�G�4]��bl13d�H��97���+��ˁ����V�|�L�<�̼� �m��]!�/r�f}t^]�϶�Ky��Y`�����<3n�L��g1
�����q�g5�������w�f���8���]UX��Ⱥt�n�������l�����P�gE��bd�U���-��I�i4H����>�s��h�s��b�u%����+q�R.�Ω\��ȯ!}v�|,=b=2�W����B�w+8��Wꂅ�x�`&щ���}2�D���TMt��D�\6؆%�Gm�mi4��n��U�^��h��/8ӨsU!�  ��vukN��b�,س4M]��\�]K��oYM����-J���omX�}xq̮v)u�]éCʥD/��E`�퇆��{+���yIܮV�i�.<,��7�T�&�eM�5�4�A.�q��A���F��C�hv�6��FXqĸ`%*���"�qQ�]!�V�u��V&�Ā�ٗ�
�z���oj3��h�ܙ(".��e�onl���LY�Խ"�S\5�[���6����,]�/v��F��q�H�5%wڂ���� W��>8_p�
�����wS���4�
j=*!�!!�)�yRaaL�O�`�g�+q'S)H�sT*��C�u&�ͽ�u����ʲ_7-�F�A��S�@�fY��E���
���"�&of!���wß+�]��M1
���z2�G�T�r�����[ަ�v.�-���A�k���1z\hEU��I�,2�5�Sp)mSÅ[�����6si�'k��=0�8ۙ�����7�Ԑ�ynl]2��g/���>n��7vGe��ݺ�^��ӽ�V/b[��mG9�k�b�s%Ү��|Ў��|��v&j->�p>�1��	�4��Y�n�t�nb8�|F�P<3�o7��Wʷ�{���,OC���L��Lm�ޑE`^h�Q܏���� ����Z��V��x}� �Lݼ��c��W��pDuIۆ�2��\�3�3�f�͘BFi���[�3+�ܛ��	qvF֣��8���\)�����ɵ`ѻ.��%�c�����oU�]f��r���v�;��3#h�{���E9��+ju��;p��ʧUMSR�]���^[�m٥f=�ӑyu�Ӝ�5M5m�5Vl�h�l�lh2r��d5�pH�ZU)�(DOK,ll*6Y�^I�Ndf�eƷ|��
plrl���"mF�.�kj�t���Ɠ��w7{�%��Q,v:�n-�lՆѳ���p�)�6�k�ʺ�,C=�$�I$�l"�ʃm �\P\��P� �-�c��i��˗5�<x�����G�X����Hj��u!���"���X�կ4W�<�rY��lJ���C&\��}�x��Ǐ���^��d���ڪ��]خ=�35	��G,"dAr8IJ�+�x�$c���&nn}�gyǏ<x��=z�=��AQ!RQP����.E���#�`q��q���y$s�V3�2���ɛ���ٮݻv�����1۝��Tԩ$�5�z�ÿ�E��7K�!l���Y2>�r6F�`U���W��.q��nݻv���8��q�'{^��IN0�cfd�#�������� D�2H*���s��}�����������g�±	R���N�{��5�	 �.$h������1)���&t����k��[5�Ҷ,��¹\�XX���c�qV�i��.�gN�Dq���d�3�D�Cdu��4E�Ķgoi�f	�N�h�"�ԇ������T�25 [K&Dr�2H(�J�ٚ�	�56��'�����Z3k,��vןfu�:WCt\�X���w%�=�E���]��&���-T�犇l"�yt��(ފB��E���	�L��ck�V�'	r��%ە8�DjX۽o<^��P��u@j�N�	��� z��! }-�)/����ޡ�}����* �]�G�v�6���c"�E��s�w���zW��:}�?��$�)2A�}Pp�\��.b�[ �Z�E�q���b��ۏ;�p��<gz��chlù;<<Du*�.��M�_r�.��;��I�^C��7�Z �����ib7�@<��͹�t��C���6fe`�k��#{&�ex��7 <�lw��ssS�������}R�0��b��C���Nq���Bk���;e��&{�Ұ����鴮j�=ozN�<�ծ�~�� �)6cwf��7sA��ϳ���B��p��i�������������z�ԓpjj<i�y�������&�I���I��e��C�ۆ�6�]�W;}t-��\����ک4q��-+y-��Jo)E�]#��iE�=�}~�I�=J>UZ�ε��nY�-������l��.��fX���]u�w6��:��9�so�]۹Kx��=Ttsb��F%#��}�[���3Z���!}}���ʲ��u[�î��w���G���nQ�ƙv���9}�> �G#�y�y����G������#�&�ϵ�l�eb���@=;��{��?D�P�!���"!ݱ�9�;�vU3�5'��{*�g�V�7��۲U�K6�2M^u��[�3�>�k���
t;cϪBj��	gh�bU�q�9�H��4���z;Uw�]كV6���&���/�U뇼�3��*�ߦ�k�3���^.�71?v�^�,tk�$0�uF(�f�--%^�!�}uفM �r� ��s��j�����`�~6��%����߰�6IR}���H�;^f�X����G�GG���<[�ܠ�j���
ٹ�ط�]Sg��VN��A��-��؈��.��A�kXm��]���ff�L���	�2ga'����q�:␆�W9��/��I�Gŝ�5�HZ̸ĽMO������&�;{U���}�ˆ��y͝���[�o"x�1����]�5��RW��Y�_.�K��fhwP���%�� q�
sq樟n3��ޭ�����ue�97�������].z!���}���۽b��x�~=���X��uo�7ُ��I&�즨���ᦣ��4��;��==:��n�чw.y��P=Y>�%,��j�o������ɞ:r��gV�W�|y�O^C�y���/Xo�ԑU�ڕ��zO?�ɹ�Ղ#��ת�>C��ɳu�%��˫�b�%~�	��++F;Ϭ�rKy��J�PEMP�k��~o׀P����WJ޽M��������7S%f�/x�Y�����c����W��Pj}Tϒ���b�r"k��kg;v��H��x[q�l�@'��j����4����/�:T���>{�ڮ����~�1ّ��+͐3v��ȥ��L�b�t.��{w��[0���/��8��r�������&}���跤�zD�E,ɾ��A�P̀�T��(6��3�߶ ǁ�T�U�B ��S	U#�6��u�f�Ky�Xi۽����<Ul��3p�N
��Lا٬�Y��I�q�D6o�9X*��K���{@�#M�>���	Av�a��=0;(�Vs/ێ�1�k9.zc���d���+`ƫ�}�<�w8K�cC���~��aW�П��>�G��5�\��>�xrdM��԰�ѝ�b^g!�6s0΍�16vx��z~��E�k��(�%U��f}�`4wE�p�dP�x.}����&YY�3�8]�ez5S�w�4��;���7�76���U����z<i���[(Ǫ�Y�q�.z3+��'0�X�������8���ͩ�j2��<᷉��AŔq��on6���o�32-�ǈ|{+���pSS �y�Yۮ{4k��~ 2q�P�����Vl1����	�-9+t�v]�=9�	��D�B��>���YZ+Ӊ,��X�-���ь���%���ڧ��v�N����wx�O�~����C��#�8�֘��jn =I�6�GDV����V�Һ�xx�b�7~����;�����k_3pX�l|:��V������Ep�\?E��w�\���Uw=G�-X���D�m[���
�'I<�oQ<�����ST��%P�� ����ȳ��ռu�׼ț�ݐ������L��g-}e����#nk �K�"Ȁwf(�<��N�&�ǹj�l�l����G)1��6n��5�"�e��I��ˢl���0�h�R�=��<��T:$L�-��F4�r^�M���r����=�ك�ЯG��3.��Z\6�*��E�B��Q���23#����2��;rF�7�'�[�9ټ�/ދf�\?��|�"=H�����([v�����pG�|��k;n�sρ�C��{nM+��Xa��&uSp��Rx�I�T'܁�@r�l�e��`���}8�T�f��ʷ�XyTM謮�wYEe5_5�+��/x���_j������4Ot���>2�72yH\¼�L�x�0ޗ3������)�6��M�֟u�����Ze|~�z��;��7,.Sʈ��*�I�hOb�蟒H���$~��ѯ_�*c�������]�^��M�����#�ļ�p��6�U@c�>x��:���p��{��էcR*���h{t-�`����
^�"Rׯf>][��em^S�;ݦ�T����!�B���/;�҂�.
�(�,}�� �M�R�bHؾoa����ul����),�|����D\��j��7�P�fb�xU����������Y��]��*U�~�����|��;�z��n|����L5]{����L�ɬ�ӎ�ͷ�'Q2�D�vw�B��v�$Uߜ؎Tʯ�z�m�F-ʣX�v�ޮ�2*gqJ��5q#�E{��Y�!����c5�=r걝|��l2@_����N��:R��g������I����"�[�f���H�L�؂�za�&Ӹa�/��t�G;N�g�Φ�7����r��Ձjâ�~^�*vom=[�H����7�[����Yn��X`჆;s�5$p.7��K���!7�A )�հ�k,���YwD�f�\o{`��u�@�l���S��\#�%�,|��7]��	�e���{��;`l�y��2���W�V�QkJB�����ڎ�at����e\6�^�!Y��S�����޷]��E��,Ė,��qj.vT'{{m�$�,V��k@g�up
�5�4X�kiA#z\x�ea���j�%��Ƨ(6;;�H�ݒ��}�uN*�^rU�z��b��;q���F�쌭���`<�4�n�3�҄^�L��w|p���b�-�tj��V�|ܨ��-޷nL��b�/B3��MY�*��Z�O��u42���ʬ@��N�;��!�2ZSi�}"^`	�Qf9,��aW���	x���3��kݝ~_o�,f�j�ߣ��O�ίf[Z�IK�{����y-��b��E�4+(�mz|�^��� �mK���.��mKp
��+مS���s�Γ&�����G��O�:��5j�V�V�d0�ۡ�5(�����t<���>�h�'o2	4.��$�]����Qp�+/wy��E�����|�aW�7�gа_m����J�Io���-W,r�ss������Js�,�l�����0)vL[�'��ym6�ݯ̬�M&�.��l�P�I>����e�{t'�s�l�x0jkOO(��䆌��C�K�m�6m�����xe�wK�]M}�q,�ې��{�l��x�ePT�w_L��e���}�3{�3ה���;�\67rHܕ��,�5�u����,=&np��Wh}�MsRy鿃pA����|�������}}��XC���2��0�G��(n��o;��+2�Cb�e���ӵ����{��S���˩�p���?9)<��?�a�h��~��W��������|�gξ�|�5���=�S��ξ�]���]#ƍ3t]M��h�!���B�g�:�X�=k{g&!��f�P�2��܉؋w��
���h$pۀ�᧝��=~n�<A��Z�ʖ}Η����C����ȇ�1��*���`v�}�i8��w��)�1�gmSN�z�u5u{ˑ�qs�w[0�	B+�:���6���ٝ��E]&;�dk��v�-\N<�n���g� ��.�S�:ZK_��
��f]B�Q�0��e�H�m���7�v��̋4�[i���_z��ꊚ�fH3��^��.��h������:���Sp�f�DDc4́Kkm����PGNK؛Ƕ��&\��Dn�E!�']�՝��S�b0��m��mSiЁ�4�p�F��]6�k^4�n�!��m�fj� ]]�(+Tt��i]бa.C�^��;X���.җ$_����Cx�T�e�z#�1%�ͷ]6�ٻ+F嶬�����KYYb2��uk�ь5DѴ~�A�?�:��rNy<����w�w�_H�nq�
'>G�����P�޾3^kf��6�w�n�ɞyR�?v�t��z]�>��Dɦ�fu�<&�+/�t���հ�7�o0���ɟN�!���=fk����)χ@���Ip�xJ��<A���#�@���u��%&���ܟ���h|�������n.�n,\'x<��2m��v��6{7'��# ��ާ�ޙ^������ѻ}���AQ���S�X_�1j��kס�
���i�1��ʪ�Eih�[ ������ɕ��ikfW�d�z�.`�77~������?kc��42�(h���N���ǆ-��z��@���Ȇ@m	D�9.ow3�]�+$�,�$gk��q�s>c&�,{�_�/\"=(�^]�هo&��Ĥ:���Y���i��_�5s�z��h�+��νۘ%'�4��X�^1c�*
*�m���t�R�U�K�f��ם��d����̷"�.��3�<�@W��Z>����4�����<+����Cv[��h���=���S��=��z���^���j~1LS1C>�^w�����Hr�3��zF�����s��C>[m?��.Ӛ�����q�&��� ��=?��p���;9��>̲;+a�K�������{��U���<�)@�;��S5~4��2����"�=������a��U[r&��/l��:���R�A��o6�l�`&&���K݁W�kJ�w���v��M���ͺ��EY�Kү=�w2&��K0«����ۖ�@Ņ
���|bL���S3��ķ��y/\����2�������qM�w��S�Ju߻̬5q�Ȕ�iޯP#�wwfv�j��N�k}	�a��x�˨].�G��r�]��,[��ffnP�����6��������yQN`
#�`�{�~��q�m�́j1oO�2(�!�X�í���}��G��f	*���z�9"l��0B�E��b���d� n�)�+�6�P��c����b�5�EX���Lm�<k��K��Qmi�*�1��:�@ӴUwbU�S���V�����7}�Eu����2�5*Z�3��b���&o4U��n[�-��qQt/*�ЏQ�-Эb��de��+{+'oq�Szs[�zL��s"it���8���n�3�!}O���1ӘW)r�a�VO0�p��V�<Uun��S�bq8f�>Xu�l���.���^����Bb���	�60���.N�WJ:^���V�7[�@���AAۼz��i�#�i���|��N�`[nF��\������� ��������&x2w�t^&׺˔H]�˩3���]�{f�]��8n��z�F :ܬ�0���B�
iq��.PW�6���r}Im��5�eڼ�G��Zs*�J�3��vI[sD�F�g�tVں�{����#�=�N�ק�������R��N:g)���O]eK�b��Q��z�^nN~�7��SN<����c7��T��_J�j`�H�6���,1�=�k��>wV���͜�)Z��gq�Y{"<U-S��]t*k0f�Ѣ�������1e�q���j�c�R�׮�p����T��<F�\�$1r
�2�NɌZo���X�#o�a#ϴ�<ҥ="�A o:��sA����e�]:��2d� ��6:�Ue�HZ�\}B����?i��wG%Xg%ł��p��O2�;x�Ǽ��Dh�ଽ88f�'�<����v0>��f�D��;±�v�:f�xc��E�?�{1g��w�^�4`����qx0�q�-Ԋu��U�B�V����C�gEy|�V�^4
�T�9'�]dQvv8��d�M
R���TRo3�-�JR]k�;\�£���J�o���B�mOcg\:"];ʘ@>����o���5�D�AtwW�p���0J9LR���R��̝�+i�^ڡ�@}ڮ����9rKu������}��0\AZ�y˦jb$K�x��8tm�tb	vef/�*��n����k2�]`��PZ4�ӠU�B�/ir�Z�u��SD�f�G�0줍���/p���E��ys�K^�����͋�[S"X�P��&M]�^]���������L�������;�2"�)�I�oX��(+�iʗV��fh�B+Z]_+�z���,���.MR��b-p��)�Xﯖ3d�Kn��y�*����V�$��΍�N�n*�g*�)V�|�Z��;�h�r���If��J`���=����ɇfȥ�v�{���sZ���BmD��2� 6�$2E��YqCDi�\����eH�w�r���#!3��e��>��v�۷��^��a2T�Z�բ�����Y ��G5#�"dbG�"1�Q�\�<�g3�ǯ�ݻv���׬p�J{55U�֨��^�G1���m0�(��c&Nc����%neq���d2�z�۷nݸ����{:��TI*����#$,�r@��T=�{��Ȑq�5�A#l�	�Y܎4;x���nݻ}|z=z��ޔ
���D\�t��2m/v�s>�a"O�����#<����r���x�۷n>=�c�=��4TH����"`��b"�!lQ�y
ݵ�����0�=ɜ�78���۷n޽}c׬pr@P쒊�嵘��&9�}��é1�0�+U��I-�#�࣒�B�V8�-r#R�f:�ݑ�.T�!�Ɋ�H��.!��8[	#$R"*HtĬH����J��LEp\dd$Ū����U"�� �n�Ɖ� � �%�_�f�o/�_Rv��r�|�}�1��,k�ڹ�^跗,'Me��uԽ:��H9�{nq�o�4P�~(j �_{�{�T�}����9�,f�9i�>��JXM��3�o_Vm�e��������9UX�(�Tb��&�����M�����z9�M�	1�����ߩ�g$61{	��@�u-�d1ʊlXQu's�m�^���}���l�P����P�+Ͼ]����b��{��I��\�A�O�����^�*�����Z���88=y�����RS�<�:��u�-��C>
�I��`��f6��!�nٛ嫮8mv��EفV���~�)^�ױ��zno�˪Mu-�Y������Q�V����`Z�
�5��f(*��a��,�SS�N�f�!�-��3�I��Ԍ���Ҍ�6v�W6��T���e� ��s��~|!��&�S�#�R�/w�i��!v��}s��E�@�h���s���8�3vP�̍^��ݭ�3Þ�S9���V�y��l9k���Ju���w�������긋Vn�Y(�%r��f�4�9��VU��s^�kx�L�}̌w:�0������k��"�z30 <� ����U��������۸l��YNIG	2�Wy�*Sw;����~��@��T��YM�~��ޏ]�Z\s��Zm��5Ո�p�ײn�ǹ�&P�c�p�H���0���(ѽ޸�����tyg�Y��-����9��̈ʬ�
j�I��1�T�u����O��/�``���[�%�5p�u��vr�Wfr�m���0b)���zI�m`�l�w*��G��g�o����¸{h^r�����i�fm����ywJ��U�z�\�|P39]�oVq��/��s]��	����/x�9����4���'uF��X2����,�^�|��pmF�okt泂�c0��`�u[>�*E��-@��n��V���xTwq)�3�@��m�;�o,��2�V��7����T_��W��f���2��K�I�[��� ]��]��c��g�wu���՗�u�?D�"�'�,�J20�$c�.k�7��DRk.����N�]��P��:`RiIuyա,�&v�Jޜ�|w����,�V��z�"o2��v}�q1���vu��ԓP|A�hF�&䉘J	ې�Kd�k"�Y��r�s���8x r�&u��SRe?_��ڝf
e�T�J��&:�&X���ɛ���.7�.dv�����Y����f�b\��4/5˳,�u:���sX5�'ه	,��cC��;Y��X�`�T��>o8k�>|>WS� L�Rf�l{O@ީ�$�j�s����^B�B���\}�������d1�6V��y���s�-�n�^c>ÅO6{:n㷩�#u/\O��.>n�j��>��Y�d�О��Ok�7~pO�p��j×�D�Uʎ5�^�yƟ\��]lz�8�ڬ���V4�!�b�w_L^ij���D��n�Ú��uh>�Y��`:��[f
�k,ڎ�ޤt��:�A��3m�IHշ�l���"d�{},_w��{�=�S��x�߷��Lb�0������::(��ݽ;)g�W�_�/�	��ټn�(/z�rF_#	��6���r�W���Z��o�2���^��lv5*�0Z9���t��4-�h��Fܐ���NL���Rn�Rl�2���V%�9Ww`�}��9��ۜ��kC���ON�NU\���oaή�f�P�N ��i�XJ���2;�h��7w���\��z!��4A���T��Ǔ�3���^�/=�tdGj�y�Rz,W[��)�đ/��ʝ�W���؀@n���lT0f��*9��Sq�CJ��]��{�"n���f;��J=}{�0"I������A���n��!Rm�m���$=��z>��f����ޞ����dg��8����/S)YÄs�:Q�f�&�5Y� 9 x-Y�c�����7.���T��<(��Y]�[�w�ǲ��;��L���FY������ou��a�
-��;�~Y��u��c�U�OL�BY�_w��/)��Rˋewtjm�v�~�7-��e'(ﲰ2ԅ&���)�,â�:�x�[�(n��x�yXUs Z�ɰ���V�m+��:�<}v����ќ�{�������+���!*��w��i���-���l�Sp<��c�R�|����J^eػ�nP�W��<4�ɶ&��[���Ĵrt0Ss������wv�}�אdF�I#:v&�]:/9�F�;R�=���k�͙�V�E�CWv��N��z��?i��b�����A�5;��燿;W��������ӑ���y�~*�f�;W��M�,���
��}ά��l>*���X`�Q��ƌ&�]{�Ҕ�����ׯ�������A�p���ggP�ͬ��i]/���z��Ҙ���vb�]�Z����s��#����P#]��5�s�>���z3"-�
gb��xeL<Kd�b������d��@\=����(}���^z����F�}Q�D��,���$�L�Cy/r�|�z6O�?I��Dߒ`àv�ihd�M�>:݋+o� ����v�����3'����:����F݇;�����/{�<��݋0�^�ʹ�`t��w����fU�Km;e2�7�x@b77
l_Eۋ'$k����� w�L�"Ǧ�Ж�����:���6C=�j[>����}���<
�np��f�wy�X�1��+��z��jP<�1���T�H��B4(0�W^	�XYաiηh}�e��"� B�4~��tB=9"P��U�Wˉu�8�n�y�]�aTG��h��h�Lt�a���~�`�1�TP��P���s�雷�������z_l@����g��4֖1(�Jʜ5V��3����ﶃ\s���Ɲϧ�����P�4�4Zjͽ����۝�v�鬩E�IE��(${��$Q�� �����p]-s��c0{w��w��;-���&;S��>��Fx��duɐ�Z*�m����Q�]�����9^x�d�2WZ)���$���<iJ0��7<
��4�e�(J�(6�ɟ4z��b2魻Et�mt�}��gb1]��ˍ���x����,K�.1+�	-<$��n��Ң"��W�{n��:��XhJ�z�3�l�����7�V�]���V/nf�5v&��+0�+�}��w�Ƌ�j����.�s)w��Ւd˻k"#�T��8��NMj�e��"{7���;M������A�^��g0ޒl#��Xݝ�w���[�.��ϕ��x�Љ-he�X.]Z��΍9k^�6��uE�b�|̈G�a�p�n�j�]���-��2M�W>��_P�l�"Ǖ2�۾#��oW7G�]4*b+8t4�7�{8��A��K(eIMQ� �HZ*BإR2�r;��� �<�a�[9>|�>|�ߜ)�����#���O�_��q�2ٳ޲�v�oK��PT�45-6��?�/4�7�P:�щ���\1�8�&�8�����B��� �Wu�~��S���I�ұ�O�{�R���ep�21r�v#qS���؈`�����+�g~�j�k�~	�����Zާ.4λY�Ӟ(p�W(gD!��;�@��~3���K>k���]]�v1g��>D>Y8_������TEg�s7tqn�k�~�����k����9z<�q�4>ʩ]c+�f�;Nt�9p���!��,{�直T50�i��΂V޻�ʑxAC��kۣT���h$\mCu��6��M�
������M�
�x�kn�z�Y;�͉q8k{T�=tF���U��jfN�/kе�h>�сQ*� ,��}��[���٦6�q����3����.���S]�w_J��:"�~�!�zv�P�i��uD1,� �n:��/��K�����jr�����s->�Dy�v�\�N��:�K�X,0�V=I#��8?�<�?N��-���߸�=�T�޻}��4"�>k�l��Ռ�Ӧ�U���%�_0��k�6T�zu@-ҏ��%�L<�w�`��]�0U�{��s��::��6R��Զْ[{���B�ʝ��k��ސ���$�s�H�����=�K�6UO)�'�������J�������A����fZ��:=h�dn��i��jd���"�1���_x��{�CW��j�`���n��kҖ���©U��^���Ut���}]k0e~4Z�
�D�\y�����E�3��;J����<;��וpӱ���7k��~���X��djި�S�Z�ޭ(����Xѯ��a�K�G���q�2�B�-�)�f��SLCg�yLy�;�4��&���I�Rg\���ʸ{K�D������{�3So3/ XǴoH#����ۗ�!����nի�N��mw$�8�;�}�H��#¢ q��"�^B��o`B?H�oы�S�e�]Xt�����n���\�</F�]�dfiκtu�R��?3�xQp��8�w��O|U����i�gp�/�g��o��H1��$O��5Y������_�uyu���ݦ���d�*����\k��Y��d�';����VFo��̡��8ax��5wz.�O
۱���m�+sN��W�0�|f����,6�r��jBUr9[�ձ�hͱa���=@�����5���8�&㋯oM�p%Y�쌍2J�%pUVI��6+�N�c���;�hv�<�lxY>�Bҡ'9�Y�:���[�a]5�n�۾��WQА�8Ν�� Q/��
�+���.�CٍN�UO�T�Swܪw���穧�v���+�'9��N��g�{����~�-�����vݓ���2sp�I�v���q� �h���@rt�F���gr�0��˜���l��u#x�oq�~� olv�Ʈ��xxl!�#�?�m_��l�.Teӳ�����e�z��{F̗���6����zz�EW
Zxyg�n���t�'��"2���{�޵"i�/k)ۗ��|�ý|��uoIe�X�2ﰕӷ���11<���P�A�o�;�F��t���=B��ffc��t���v��̓򽸆-f�έ"Ć�~��5旽���|��v+;/z��8,�k�T�_2�l���]�9�TJ	�]o
�n���J�~����a�i���j���E�k��bQ4��]����]-�WX5�����aq�羾�U�_Gn��s�Y��a���6��F�>�ќρ�R�f��+Y�mk
R���%��=��r1��F��4�e�����Dc;�9G���O���K���x��ȴ+<[�X9FRYU��.8ge��k��&����Ƭ�W3�~ͫ��ɾ!�w�9�������,���ʅ��V^">3R#��{Wk'b^�?lv���ӰG=|-�>�M��/E�	T񵚷����^��^���î&�n��[@$��=7K3�q��E���~�jU�:�::1] ���,���oxR"�U�M�ӯ+3y�H�z���a��n�#uiQ9�+ �`�۬j^a{#3��}U�O@p��U�7�]ؒ��p&֐+�^�lj�y�p�� ��-B��ˬj�XD9��Y���9��%�I��U0��6�J�wov+��Y�M�O���z�bbq76v�t!�Õ��� wE�P[s�;}�B��Wq�et��m�5)������Fz��ڭ##�gԒ��wXGd;��}.����Q�0鏻.�AW����r�	iWz���!Ft=�np�mvP;�i��D����^Y�s�XΏ�X��+f�V���j.��l\{�����>�]iI���;�,���R�0𼾇����d�)������S�d�2wu���[L��6N��[.���e6ǝE�ȳoe����)�I�g.ݼ�wbw\=���gL6e��:
�uuخ��=u�AYu2��m^�Ӓ�컩�N��xhZh����l�e���s��aKk�ќ;�Vmb�p�t�Y��.�y<u��NfK v+���J/6ɭW��+l[yw|:�i^�4B0��<�^n�)�Ŋn;��5u��;`��q�u�œY����9�"�H�*�D1I+��)�fC>�P�����v���t.&���P<#�P�A���tƄ��Yl��A4���	��!2���P�@Ul�a�O�!�U�'K'���4"f�Yo]H�$�W6�&^��P�P5,!2�a�I!��y�1#~�U��!�	����Vs��j�lVF2V�t;�"Y!�vD��E��}xGM�@��2�\����ku8C�����Ԋ�޷J�r�.mB���zEI3AUVK�-��b~�譚�5�s��M�Wqrwk�ۥ��z;�}r)J�r8���$��&�pƍIN2l}c��,ɵ',�]�gL)��w�tv�M���9�ʝ{��N��P�g%��I��(&�:;4��������̤�t��
�$fi�N/��7X6�R�w5���:��G3�cM�IY��%S���`w�!j��aL��7�ɜ��'�<vz��u��[�G)�� ���_�s���9Q�Ҝ/�|�S�>\��Z�b�:����F�h�U��v�S[q� �̾�2���Bz�!8:���s
��m�+Uf��6]������ N�f'��c�`3kf93�Z/*�ۤ4�ޏ_T�;i�g#��v�V&��"�a�
ʗ���7�ht�jN:*l���,d��9�.ܖ�©��d��눢�+1>��!εÈ��d�1�2��gj��ʜk$}SXoJц7��4v�z[�:�ڬ�*�L4��-���k���a��Vͽ�!�1d>����r��ċ�7���N�6"d6m�A
��!�1P�dݣ�l�qg ٻ�V͛,E�&�6�m��$7]�d��K+Q�ݺ�6�p���:؛6z�Uȃ2:<T
�қ-�h��L5�8�A�B��jK�QU$$5�-+4YI��00��BR#A3� �j�TwP��Jd�B�R(�iY�v1��[�v�ɶ�Zh�J��)2id�/�NχX�ń�~wMh���s#8IY�-��ĎDX���s��\��m��nݿ�����>��{�N��*�$cS�:���D�A#�6il���A<ϳr��g���nݻ}z�ǯX�����!�.�5��^�Q1AV�2�ܤ���^�$���:t��z��nݽq��^�́ؓ���T*Q*%1+����=��6�DOXd�#�*������k�V=m��ۏ�v��X���w��u���451H�Y�ש�dH8G'&E����9ć2x��61�3㮚PW�v�m���۷n�^����8T�\�ȓ�*�<�lq�B�(�$�9au�}5\J���nnGm���nݾ��ǯX����T�wF�Q�j��8��bH�Y��id.��E�!��M��0���vf�@�"�#"��DLQ�iadb����:$wn-ǖ\VO �Z�`m��MwG�qN:�A�v*�+�r��"A�A��$	 ���eG*DYյ�c��1
���IE*�d�e!2��ӻ���Z摲4'Ι(�U�/�xm�Y���#�2ccCD�9X3z�ͻ���4y%էy�st��YкJ.ؤ}c�d�i[���G�#k���v��L���,����5�,�Ƶ��۴�h���5 	�#�H�}�v�|��y(L@�jgj�q����ɳ��>�l5���d�@�i�SY���Ǫ�t���Hq���n�r�љ �v ����v���K�T�%�eY�Om3�Dttz�}-��)%=�ʌ �Fj>�
����d��-|o���v�}��J��
��{}˨�����#Uzd�����]|�)�_�b��I�k��,���*����)6��]
�gfۡ{}[V�a&�-����$�Ҩ��[�����+��0a����v3E%�j�|M��^�bD�|���3=�}�TL�dGj�^F)Wbc{@���rV-��&�1�am�< -�f�2������S~�ȣw���ج��_�*e��3�yh��>��P�'K�z<��C��cz\���w��v%差���W{D�R^}�'�F�����YApv�sm�U��c�����Bb��^|E�	.�Vǘf�p�ٷ�qо��n1��ҁԕw�)�D6���޽ee��{����qΜ��|�ߐ�s��ޝ��jR���k��[}`4B�����yٝW�x��*8	�����\ӑ���o0�� 8�0`�E"��Q���dc�Q_�ߜ����!y�7,f���)�L�%������ĥt�~k滀�^�4��g���35<�2ݩ�����Y�a@g�q��{V�3-��0`,sD�7��3
}��ieǋQ���L��4�ͩ�==k֩e܁ʮ'ݙR�>���=��)A��k�eCX�w�mq���F2��5(���z�FmF����j�L�k�i�y��e��B�^��y@�Y�� .�t.�F�Ʋj���4��m�_TϽ�v�R��x��|uZ�(<�.�n�~J�m{ys��/�輓9�k����W�����a֬ ڑ���"���,3W�Im/o��e�
[�qL��7p	ѯ�/ͼ�˞T��!���r�sf�V�y;����s!Ǡa����{���y�N��B�B��[���6����І(�`�'F$9N)n�v�,�Mk��وAp!&?%(V�����`<����Λ.=�Z��mj㾬�Nkw�*���<��7�8�LP�0�X6��d�y�P��=�0��z�*u��3��233�clu������"��?��@Î:���D��t%����#��,�j��b����v5�du5�F���}֎6����suN��+�3���d[���u�[�3q�Kv4�:2Ne7h�w�M��!�[��`��.��>�Y�u�wU�j����6Dˣ��3N��(�3�>Y|��?R/}Nލv�'ʣ� c-]	�{=F�)��Җ����T�t���\i���桑�N�I�=c�d��W� 	����=�~Qۇ��3Y�,��o|k�G���c�S�ձ
U�<h���5���B+�兲Ǣ�$.ە�o�r[IYE��D%���c/;�����ۗ���Ok '^̅0(����
/"]LJKWl�#���9�^c�����:"��!Y�[�{_�p��[Oe��xUV_����j<�϶����=�'��`h"Ь_��F&䆡ޖ71�B�쪤h����y껫���������t��nK�Tsr�嵶�jWһ������7��*Ny�5�����0`� �O$��{���mm�ϡ�o�i�@0�ܦ������g7w��d��7�ޞ���=��<�O���ox��}��M^=.��$b�����n~?L�J�� �,�}�f06O���t�f��p�f����08mp��Lq)�VN��!{��+8z����Ӵ_MtD8god������/���m�����W�6�^�}���>/�/~��}wY�淓��w*���uszy�Zk�k�fy���	2rg����&�������;Գe�9�}��"�x[n��q��h��nZ�@��p�#���P!��l��0��N��g;tX���3�y
k��o�-���^�뻆�b��枈�����5�L��Wu �P2W�5�SJ7/�s���oF!9�D������p�SNh_M�t����̯�CͼYS7/ܜ2�����iw7S�A.U����J�B�V�񕕾2%�UrOQ��,"O*���R'�ذu3�Y�W7/%_z�8k�WK�G]�]J����p)���[�����v�����R��Z+\޲����|'}�ozK��\��-gWi��o)��ywM\�M��m��dTU{8r\~o��醾]�س����ђ���9��1V��
��#>\q+U)S�z6���]Qӡi�Z�*^�>��S{�ܾ�O����P����=��LFJA+x���m�Ė�*}�?���$����{�������W]����b�qH��aP�\����:o�_�Xq��G��,������IĖ�H��~|���AL�fv����ˍ�IL:�r�t�`Gi� +"�x<�ym�W��2A*�X|q[:�q"�Ta��UQ��	E�zWzj�70��Ĥ�i.i��{G"2ӊkdP�ɳ��G���r�V����ʌ>������ڐ!s�S�����)L�2�S,v�0f�굀��B4g�^�/����+����y���Q̗��&�vL��T1="��<fv|�+q[tNz�lq<u�z���ǂ�G�mtհ��o�����4;er}��iگ6+wjif]�&�y�z�S��z���io�0r�S���n#�r�ܔ��h+��x[�;)��i�Y�m�f���7`tS{�ݼ�q�߇,8�$p�V��"w���s�w|�	q$��,.[�wU�#J�x�I�'WVw��e w�u���g�(C���cvQ߯�F�cPw�����TF9x���L�g�ǃ掹�{yz����D�;���]�������\r���['"'x�8\�z�ߠ��SK��?Fc�0ײ��n3,�7֭��L�f/�gv������$s���rՓ>Χ~�}��Gz�x��O �9U3�[1�$d��r�Y�L6��^M��%f^���R�/}v
ǋ�],v{�q
౥�j�]0���o;�(�^�
b����YAq�7JA�SH��]�U����,��tEB��q_�	����.F`&�	P��eFu{Z􇆗�М5��v�/V2[�<CǸ)I�m�]�+{�.�ƴ׿y@�"�{j-]�"X���z�sT�nu�R5�r՝a��4<�N�&�M��\2�^d�7:��
��t`��zd����ɑ��s2�L���wxv4��x�����8W����́ٝU�EL����9��`p����M���[����"����T
Jv��Yً�i�#CF_�����}��
��8k�
�ȌCR����Jԩ�������4�4���=�,����N�ŵ�N�~&���	�1�ũ*7݃�^�H=�#�s�\`q��Ox���Z���t��~�	�G���+n{s�U�&	(�i��8�PI�<~��w;�{�3y�ܙ���5���u�p���K�G�6۲No\D�Ԟ�oX�]�>Ռ ��W�߹�4�nIV;��������y��v'�_�K�����X1�T��`Z ���-����"g��sG�\��X	���{�Ȋ���-%��w���>�������}������4��{�%����;�@d��gn��ٯ�o����^LG�ay��􅇰˽��Y_�Qt�v���S�w�xGۛ[B�0}�V1�}�R&�H�:�g�m�>��(��޽�|е��s��uo�g���W=8a��{��,��%M/;�!;��Aޗ����w�͊N��u�;+�����Z&�1��:�K���\o;�����B�P����e�ϕ5��.�ǈ���8�\s��� ��o�,.��7l�ƙ��-�sYc���Ω�6���K���A��$��UC"�T���e��zT��p��@!�fD�d����߁o,/r3ʽ�C�u��rr4�*���6�B�J��n��S��/�d���Ṣ 
}@��g�re,Y�;ں�{u�GV6��3�|W���c���j^=�/m�a�J�T�d݀��3Y��WO�R�8�5�##2G��n�W8o�@��Bh΍��}�����z�Vwu�]w+����4m��:��ο�E�����q<:a��~����>²F�-��ά��R;ۣ+#��`4d�~[1QK	�|�"�?{��OcZ!ٝ����v�[������NL�V��r��%�\?��!��w�T8Tj=Q��	Y�w�W��2��6�v�6�|�4�tQhZ뾰���J,���gd66-�����O�[c:��g[3�>p��w�MpR �$�qV�%Kv�u5׏��9��j�v�țm�]���*� ��:_\�ۺ{u�4���ݷ!�r�[��*�m��ܓ�kO� i:�T�f[$� ��Kv�dŖ��	�fm#�2F��d��1x/��#�]u��;�w�û��0��#��o��yl:78��a����ŏ;�{�)hfWâ���k4m��f���a��z�����x�_cz��(�a٥���I�Z=K`A�k���6_�Ft<^0e0|~�O\q%T����7�g� �v�$��� ��x�����oS�����8���5VR�3^�ݕ.��=����TՐ�p����x������*�Z[S�������Y�H9U�)d�{u�}B��B�4��Pg|�,^+Ia�7zi zݽ����gg���[X��aU��S;*d=-����{k8�}���	�2�UO���͒�_�T7��ߒ�f8Pj	�.�+�-�h i��?ܟt��φ��?W�^�s�����2p7vîg����wu�	��|[B����Q0���l����%��uY�+4�{Gf�3M|����ȅ��Lsü2G��VdUsbŅ�*�'dW&��%�A�;,��w��c��sXX��j�Z�\� Yr {�ˌM�q��ma�T�ۀoN��omθ˰����a��wZ�S53|]4�tfv�n�z1�OQF]��mn�2�܃�U���n��ot�-P��f]ȥ�t�#
�}�j<��{	�%��G5f����4���5�����g%@�a����Nes�nj�ĸ�Rd��nF����22��8W�}4�����4��6K�,5Q�afx�[\fC_�$fh��_ o����g����	�om򟼇��b�k�U�^�neg�E��wfzF�n:&(�P��e�o>�>�^m"Ӷ6 v� I��`���>UH-��Su*����庙'6"�1�6�z�o�Zת����ۖ�>"/�/���t��N��3x{��=mݡ������>�G�j����12�LW!X�ĝN^�UUT�>�e�B��y5��� �t5P*��g˔^� P�j�x���k-�<4����0�͝�/k���^���f��St�*���n�x���lb���c"IX��3ˤY���e���M��q�Gps:�a4:��iL�g�O�n�4Q[�um����)�<nR<�p1��c���� ��4b+�\��*@P"�A�n+]�9�uT����f�L�[R��Іf�\���Π��C�a�g�)�q&���-�I�9p#هOq�v����*r�����0gudb7W�{��7�~�+Z-9(]�8.�'��H3����M���˨˸r[�}���n]�k"���V"�7��lmk�|��V�IK�lUD�X�h7��뢬�S���'�z:)�SIΉ=�z���Eu���}�u̫����FoLg_B��S����vqwH-s/���c1Ί�������"�$!�V�G��*���:�ڱd���;�6��*+��J�y�b��Y��Z��/���5)�XH��j7�sM77���(4x.�Uڢ��Z�'E��X38�Yke>���r �!�Sv��a�j��f������x8Ŕ�����bvwof��oU�-#����QU�^!Gm����0��
T' �dF��WNv���T8�yn϶��*W��Q���`l���vWee�u=��8�=n	G��*	E��k�>��2��_5N>Z����{ܨ㉁v�=Sn��t僝� ��U���g8M(��)fb�P��s����Z� �=eW��Yz�uw��[0�e�}�"�aގ��[�7Mё�-�!z����Q]��^��\(���
�鷃ML��"��[�o�FG�ܲ�\�hSM=V�/W+�%�Ίp���!w�ͻo/u������v�ޚ�vړ�&v�	�N�T��U��ŗ����2����(��7�2�ۯi�i�V7]��v��b�����`�iH�m�ŰYؠ���!侜-����ad��8�'/v�Su��8V�k�p�L�� �5.ן�!�����Ң��!��<��J�7.��x.����I!0�/�7��X�.����y�MX��wc�h�m�9��z3z��P$��o+XH���K#�ɩa�ӆ�\�.�%ը�G<�c��mƊ���2��Ox���qv�GU���WM̒���^�5�`���t�F��OBMܙ�Y[òr��:d�p����E�8@��ܤ���]]ϻ��t��k'�a���>w��:=�&D�y2��"&��p㓐���� � ������l=���d�~�t��<v����>���3=A�f{iy%��
)R��\�g��o���M�I"�_��7cɄ�M�&�Uq�N�m����nݾ��ܙ�k�E��FA�����&�il��.�-��$W5�5�wb�f1ȎD��=˛��;ϳ���nݸ�Zz9�]r���+�[���v��f<�2�p�lr�Ŏx��I�Q�m����{ϲeβgY��;v���1���(��*HT(ED���9$Q�����a$��5�I9"-H�L��d�=t��M�>�x�۷׬c����2%��d� ȸ�&.����\����f��HŌ��&�s����N�����ǎݻ}z�>��������p�%��EUU2$�Ԁ�Eq�LVc�d}��� +~�^KdT�LHH@EX�U#S��X�q��Q�$&I��jrX8���8�W:kz�
�0��J�f1�!B��J�I�����X�,�$"�-Đa#bEǮn�#����#���(���BY�� �H��]}LM��e�7��.�8���e���=2�e�8�o1ϛ���R��S7';�<�Fi/na�_?䇨�=<�=v͍�ꧧ��?UZ��ݔR�6U�[-���%���xε͖�ꥷ"�h����L�a#4�=�ϳ}�M�	+��9S���>�����P3���[��8E$�V�}����>aM�<��-��0����=*�b�ʚ�k�7���Z1a��+�;�roc,���Jun��S�2h|R^��w���zzY("����O+�4cC�zl.l=ǜ�З�Er��~ޘR�]��ao�ҹں{�����WEnFX�kv%�=����<�㞪x�4�����	�/u u)�*F��4`�\n{a�`���4�a�@!������Y��D�>��g~;��ڮ�g�1}��y33p0cղ1l"*:4��F��`��v��g�[yN��_Ͻd�{b��_SQ$�v����)�x��|�&ᷣx8[�����e\�:�Ö4��X�:�v�~�5����kҘ[�,�m�jl�-��
V{N�4�P��T9��5���n�1D����V%im��zK��-�w%Y4i�z����f�O�ѿ�o\�{ʇ��W���z=�8���Mt���i��3� Ļ�'vk�K�,��=��P6Y)0b��W*q¹{o[���ؙ�>w���D�-Y<G�'�Y�`a(���~���0}A"������>�wUqNwmj=���>��}-p���%R$�y�K�Xf��O�V$^���2a��g���j�VnV���<^��+v����g�����ŏu�]��ӑy��6�w�.�@%5
o��u��	ȯO�Ͻ�it},q'��%�mF�صi�yd=Ax8�)��>�r�t)������A �uϗף��+-t��vy��P����'M�w�=w�"��,�1�>V��-y�F*��U���U�lnp�=�NH��׵!��u\����|6���T�������;��n�x�9s��� ��~����:���X�g����0�/���q5�$���gr�}����{�WUǃ���S,�]=V�ڒ��,�>q��Y;r�7X��H�4 b6�ɋ��QL�8⇎���E�zq%���iyf��l����#���k�ڟr���(Y���	;dW��p�Knm,e��;�p�})a��Ꝼ�����t����#)u�c%ݳA7q���1LD�^u�ǌ�i$��?����;<<ϦC���~ص�L�*{1]1'2ƌf���2���y98�U��5|�A6=Bd��v�Y��8׬�쁼Z�[�/���{7���psֽ�3�y�}0�w�Z�#w�[�\r,�{��-w��v��o��O��Z6OWzB>�јcxe_a��.Ub���y����4��{�R,M��o�s����dQI�4�~��1�Ł�	����X+s�ƶ�3��D"��֘>5�y9�Tf�D�/N/]W�=q�Ŝ3
8�&U)��lz:�{=?oW`�1�UZ�B�{+x6�����Ɲ�$L`���ܲ��B�k�pgt{i�m�T��$���OsR:}�n\�S` �R�q��l۹�b�r�\�99��8�{x��A�X5U2��k˙�6yq�_3d�`ے����jb	6��;��u�C:(۳��H:[OE��F���i��t��A���Wwb\v�Tp��i��<�����	����׷uq�j���o ����Vs�
3!�ۛa����k��ff�=Fr {�ۓ���]�w�V���M)*�*ۓ_��c�W�K�.���i�<�PK����}�4��1�$j�.'�����[��C����<dN�ꮖX��7���ҧ+	L$ow�&;�!�ـ����󳞃�i�%u����e���{]W&�n�壣2A*��[=M��eK�+N������z��7���Z��͚䧳9[@�����u�&+�i��g����fz�.mIFǴVuM%uz��]�̘��<�ܕ��V�YJ�AF��i����Ţ������~�%0|u���|��*]Fvov���ܪoTGd�6_�0�3�f|��=>�L;�\HQJ3!��{Lfi�D=I;�!���#�Óސ� ���m�ɠ��jeu7SW�\v_�VN:�@fK��b��MPh��{l���o�=�E�W���Ý��W�.��r�x�lm×}��u���U�*��Pe����R�C��4�.m�bvύ��G�	�C>B�"5ȗ�S��{���J>���5��u�V�ՠ���9��])oHAv�w.��y~�dxa��eIw(B{�ӕ虾��쿣&�F�\3�" ;�=�6�Z"y��n\Ұw����,�-J�ZauwW�p��V��4�1n[G{Ev����6K��{������lZ9��T��M�j��u��Wz	��d�O�8��;�� 5m���/MTq������ZXX\�&���\Pm���0��4��]է�����	U�x�|�e�%kݓ�_!V�j�o�Dڌ7�P-���?�P���E��@��?��p�[��5Wow;S0h�碟��W�RYxys��ה���X��K�y�7]Z��� ��43���\gӑ�慨�4-�u`ԡ��-{i�9��W��ё#w���iq��#�;%c'��~0�u�d��n��ƻw�l(99����dC�J���GO3@p��vqx0"�6��%��R���u�q�͙�����9U������O�_3�r���x��PME��qa5�|ܺ���{��G�xj�w�-��9��_X��O9%,���qqM�q*����	2��wp<��1f��x�ʯ_�n�p҉��oX��kp @����a��v���!d4['8ο8e7���z����n��&:���0up ��)]<D0�;+{�^�,w�� ��|'�B|r��c֮�v3>��
v��s
|��m�%P�Z��[{�a�`��C�2 �y��2�p��X��nw�e���R����fp��`/��2�+0�@�R,�jޟ]\��5T�R�ܦַ� �1�"o�E9�Ɍ4�2@h0�)9l:�#Ǝ9�36�����=�	[Y��@ޣs~»h����_~�w���T���.ӄ�R���������<d^�a�x�Kd��8�,D�*��_�R�/D��h�z,"w�y�D�����׫wqꡚ�����Ip=�iQ>��ƍ�I����p+I�	syI�Hs�3
V�Թx�]-dˍwg1��ڱ9B�<��z�o7�s��]�'�;��ݮcW}ّ.��L��$S�6���u-J��k�Ȫ�L� y����A;okwr�Qъ�"[���1e��7�Ug�rV���~ss��n�n���si��zz޷#ɱ�J&�v�M$�6�b���;q�Sr���`D��xwMlsVY�<*C�nK�p���,�Ċ�U �h�
��T��8>��||�=C}�9מ�����񻼜�Э��=�#Fo	��y�P������F7����fG�ᮈ�K�OIR��J��zv��nC����6ѕ!� ��Rq�$��G�۸`X����x���q����Ր��X\@��N�����]��7x�1v�V�	EN����i��n6�c�gq7h�Ź�a������A|�	�J��좨��F,i�ȎsW�)Im;{�������v���y%@Ga�\���5�,��	er��n��c�˸`��Qq� ΋`��D�w��ϠU�n��iK/k�����gg��,u��h�{&�,ƈ��;�^|���c����$��W_�/^�r��v���������5�
�W���\W��Y9���(k{Q��	�`�� �=�?]+��X�tѰi�Zݬ� %L,��:��MB�z��4O�X��!y�w3%h�=�����m��&�#����V��W�db7�-s$��=ٕl�t�t�c�V��ϷZ�u��n\��r���33�~Џ{!Ǚ��#f�I�#笮�s�ji��.��[�6��h��	��{�	j��3�Z�\��ʅ���ف�.P7�/N�G���׻⻹i/l&�'�R�����}w/뱚`^O�uY<j�H�љ�l.6p[�ގ��ۻ��}��*��x�vUG������7��}ڧk�E7�GS�l�ݸ8MZ�U�U�;h�-7�'��c)f��!����YZR;�7����;_�CS�EE�Tg���s<<1�պX�����x���$���v���.�>���{a)��W���ǲ���������{�`��|��R��6��3�g}x��y�
WV��3N�n�-����	�b��5�~��
6��ͯo���������}ǩ��}퇷�&�=�1�n��9)f`W�RU9Y�^�`�;�μ���ܔo0�i�ѕ}�R� ��u�K�;2'��vg�{��Ϋ�o�_tb^�ek��g�<���=�1�+T+р�kp��^g��K�pn�����IM<P�9va��b{]<:����zN>ɶܧ��f@{���9�K*�����ꑛ:Z7|��������Y�RQ~��woug;2&Y�����-�1�Y>�}�;#z{�X)��>'�-�#�-�{
����^{/��Rrg� �~x�faf��ǟ�Y�V�����2��#����<�+)��X��.,���#���vd]4�"�o�] ���5aX������OO�z&�P��i����o(㐩�e���;o�Sz�u9�h�ϒԀk�~R®��c@����SA;�t�x�N�0�|��x]Ov>.�=��k�����*��w�w�˺�϶���p�M9)lڗ{��U�g��hL
�����eI�x�:���ב���fl��h��]o�-��P;f����ٌ��G	>*'˯դ=V\���<���ʃT�w+�@�|_�n�X�
mӷ�"P���/�\���8�-�l���ۂ_3�Y�-���)zO4�<�����'�Υ.��47*���)�����Nu�ü��W��V��kN�X����۷0I�:x�|�+y���J����E/��{���?NI)�2�~ϧ.g� U��g�V��� f�3+�v�+�4_	�ژ�>��lT`��/pD{@F�K���S+ګ����'G��Yjoz[���J���ig{��Ψ�)�OX�Y�}p��luqop����f��8�j�����Ot��g|<>�+^����_�A�R�H/���Lz�;��l���M���8�_P޵\����q��W�v�Gy�n���Uw[�����̞^�^��#03�/�q]{pr+�; ��wx�CM)��!�n��yobi���{��R�f8l�#�Y{�ϬN]p��e�^���\V;�g!e�zP(V��w�̀m�7�SZ�,ɘ�ؙ3f��ǯYO�i�q���;��|����K΀��ruU�%�&썷��#��=����lF�_�Ϧ��?w����y�ꑤPAV�� 
*V��DO� ���*���AF�  �10���T5C�"�@B
��$ )��B(�����B��XȬT`�Q`�Q`�`1��E0Z"!*�@B�銥� �P!T !T !5��C`
������*Q RQCt��!��! !�!"�!*����� B"�@B"�@B-�(�����(�(�(�(�( �"� �0�"#��B 0�� #��� )�B*0�"#�B0�"��4�@B0�, ��B(0V"0B"0B"���RP��B 0��"�@B0�� #��Z 0�, #��B(��" ��"#����`s�\��*�$b  �* (����u����<�o�g�ʿ����?��C�����$�?�o������A_������EP_��AX@?��������>?�?�( ��_�}�����D�����?G���`W��?)D���@UP`"��" �*2",�#"#"� �"��"� � �*	 � ��""Ŋ�"�
�
�����
2
0�,B ��� � 0� ,(�"���" ��,�"���`, ,���0�0 H ,`,",F(��"�(���"� ���"��1"#��"����� ,"�"�H�"������",��"�R  ,H����1 , ,��",�0P ,��`(ň���H����"�X"�� ,X ��`� �����`,+���(� �����"H��0"��"Q�"���0H#("�b��P��(��  ȋ(�� B �"�B��������� � ,�� �ȫ ,b"H��(ȋ", �2�
�"ȣ", "�""�� �� ,�H�,��2
�Ċ��@d5�B�C��Oԟ�TT��D$AY P�}����_�� g��mL�
��*�?����y�	�ω�*0?����$��~��
�C�'������'�U�@����C�`����  �������*�
?��c��O4��O��G��@l��
��~H���X( ���`bH�������~��B'�?x�?H������� l?>!��?5������������.`L�����A^�����I@�6����|^�:����Gl
�تS���x����!�����e5�7� >x� ?�s2}p$�|�}�V�	j����Z�������j%6�J#mm�U��b����T�����m�ڱ�2ِ���4hc��-�eU����٦�Zj�Y-2M��RZڶ��`�+@����m����(SdL���UZ����Ո��E*dj
�cX�+d�����ұ�������
emYZ��M�@�Z�l,��l��l��mf�j٠�"i�j��m�*����IcjdS�5�&ةJ�&`�ai	��٭jպ�U�Vf(kp  �>�f�L�[-m���(b�����1��)CLv�Y�[lՋ����k[+iU�U�kf�'�a�:���V�1�a�,ʪY�6ٛEmY��cl�m�cI���  ��@$B�
;��B�
(P�����N�U4�k�w6٭6�j��Z��֕��jU[ive�CJ+UփmY��]��P�n79�"�j�u�ke5�U��i����Z��   ���6�Ҳ[K��4��dj�����ӷvmkUm�]n`�@k��GYA���Z����Z�V���j�(g`�C\mi%��b�Z�K[dO   -zm�Pښ�A�X����BX�]ڱ���*��hmkk[h6���T�77��eUV̦�κ���,��Ғٴ�[F�m,�[-�  �U0l=�EU�X6�kZ֭�3�N�r���Am��kj��Wm��c�U�F�muR�H��n"�D�B���[L��lC�l�  �ժ��c^�;aUh�H�ݷ 4 6p �����q�(  Z A7W h ;K� @�N�F�R*�[FkkY�x  �  ޓ� &� �h`
 W.  �L4�k 
hݳ� ��  �L  :�f�lSe�Ʋ�4*���<  �� K)� n��  ��p  ��T M��  �� ��0 @ۗ:  �u�� h��J�khj��fU1Tm��  �xz (jj  ���  ;�\@ �֧  5`  ,��  v�  ܶ�( �� ���CFi�lҪm6�+3o  n�  wn  f��  �  k� �Y��4 5�  �sp  K @&V x'�)J@ �)�IIUC#����#J��  )� ��   ���D�➠@�E4L��  �KZ��V\eG%�i�S0-e%�֡�XD1�Y�(h�.�Z���}U���yz���HBI�!$?�HBI��	!	'��$�$�!$:��t�\Z�Y�Z� u� ��!���J�(��[2����>ǉH�"�ɶ�IDe<qP���L�SD���mdsR��]��� )�X�y-�Rl�(�n$���*h5���b0�Ub��E&8�]��\-���B��J�� ಣlJ���̼��\jRP�DV㼼ZP��(�ļ�����X���1�9S0)�X�2�խC��zP�:�׿l��,G�8���b^;'ʐHT�u���F�2M�?B�$©�mݯ�5��7���q٠�P�� RaF�pk�����Y�m�ޝs"ߠ�hݬ�]�/�J�v��y�$&�q��@�L�E��r�ז�YH6kss3*�!f&�T.�S4f<Dl�i��CE�e],ĕ�q%((��5�e�M��w��2ua�7����rG��9�L�
;�s�뀚�}Z���H�̠f �Zf��3t7Y����Hg �w`�ͨCv�PD�x���,n+�Z�7JSM�xh�g=l�F�=՗x͠]]b��L���2h��lBB�y`��5N+'�,��t�R�E�>s_��1�^�0�;[��e�E`T&��f$[edbe%��J��GVWz�&� �R���O2�h��Kg>��#�kkf���p�fiE|cɓV�ڀ\t�NP�ӎʡ4��ɍ���$������ja[���`�I�@��$hB�sU�ְs"�`,{��t����T�B�nՕn�6��'��<��������|��̮�F�j\9�tmݺ-0�ѽi�� ��ʍ�[t[�RM�eQ�M��r�n�J�mJ�yOK^K
��u����:��e^*@��G�azA}�"�ś�*�#sv��CU� �ѳu�������,�&�;X�z�YaMjƕJ��@������5+"��O����4-�Uuy���pf��P�En�ZKt��v�ò�Hj�U·m�t�r�淥e"���������P
v򡿔�{a���C8[��� ^���q6��8 ��kRX\�rBX�t3�kkQ�7bxP��A�f1�u��F��1�h�*鈆�O4��Lyf��0�Ԭ&�n{CHT�N<�W��� �{+��.��:��u�hB:3<�z<I�=!T�	���[�e{�C�MY&��b͡l�|h�W!Y��[|��v�@��� N��*���I4�U��ʙG 6;XңZrH�q��E1�Z���-�5�h�]�H��cM6S�f<����c���ŰR���p�z���`���e�z]���Ɉ���4��m�eb�����]�iA1T��j�9����Zʄۚ�̇J���p��x�+N�BA7�f5��d�&＼}-�cTiͭ�i�d�v�޺oj�
1�74�L��ejX�k3+a4EJ���*/p[t)Dm
�³*aA!n� �ݵf-Ɲ�B2ƒ��wF�,Vw��]�:Cu�EdK"��Ѫ��8mY�]�W 5��)����c`(��1�[���b�u`5u��w.���Xԁږt���9���E2�[7��4=�X!��U ��XU(�\��D���V�k]�t��#h&�Ʀ��"�������k�fOU�
��r���N��XrQ�]J�g-*���-���)L@1�j�BɉG�%�x#�v����N*��d�r�:LdR��<���0c_ۻ��g^��B%�,V ʦ�Xߥ
�Q�^n�`d|}��F�]Xl��k.	��LW{����QiW)�Ğe�޻=O�@�Qe�_�lE��1aVzA�Ȃ��[��=imԀв��yz�(��z��v����)Qli��ȅ�6�!��M���n�o1;��,c��F��Ô#t�����6�M�ln��L�4�.h�t�)�,�	 +�@m=��ˆF���fS�Dۼ�t������JD�c����f�yRF�NP
;�7�α]��z�ݵP�#	e�aD�5XS$	��/J�s&P&sw*ٖ�$%�`ͽ��&RK6���iw�tɦ駖��
���J�Ǐ)���T�h]D ��C`��nc���٭lL
���QV�\�5��Ŗ�75%�72S�sc�#6<��	c��nL9�k�
��K+�F�e�Sr����Hd��^�_M	f]�Tw5����!u.��e%+B�cn��Oً7R�1��4L�qƦc��+i^��Ӯ�!w���a��2��Yy��`n܇I�#r���r���cy�}�!��ՈS����E��F-�3//F��,b��	�r��H�ڌ7�h�.�]@+N'k*�Wp���#g�j�B.j�L˶�x���ۉ�T#�� .Z��*��/��`J�ƌ�k�L͚V�7�.��0<���X�Y����̲xM3D�էt-+�x�e#V5dó/Y7�����t�$���m�pڽ͸�2<��v�MҢ��qR��z�V��GC�*�.`t�nL�<aӺ�=T�tnW��ė�:��]��m��◊&��6 1�;�榶R�KE^�+n:�+1I4R�!�n�ъ�0�d7 z@R���M�$yu��~z�%۹����Vcl������շQ��rV�71�N+��r+�@v"�tٛ�Tƙ��*jg֖I}�c����x�$�U��J��P:��[���$��nS�9dY�m':��,�݈�ݡ3*)mX�
��<������u�uU64����PDh��nlFe	� �X¨�&4/�"�%�^���수�L;�3�[n�!bٟl�M-*���P�d��*R�Z�J�_H�K�3/B�^QI��[��Eݕ�5L��;�zAh���7��0��!�7&A�l=˔��ہyfH�eIM�N�Cٖ6��h�A��V��ص�5m�6���
h�k(㙰�{�)L�`�fO�����0��@�ͷX+o2e4�h�2,ȦXv	��7`p�6�>C���qB0����<���I���wLZ��6K���h4˫��]:���p�N$�Y�E��x.2�f^柖�D��$�hL1�i����9��JV����$UdNŗk�s��0�\d�W�3����0#i�-����4��ou}*),��j�1	�z3	#qY� ��H�\m,Qc�n����]֕�j���zF�bn��,©\K-�@d	]0�P�y�#/a�X~�J N�efޱp�zY%�޴���6[�7f�9�m��iÑirX�k�e���Zx��
Z�a� �!nn&�&<�x��J�Yܣwn�62=T�/�6TV5xQ�C��q<�&�p�K/,2�L�] qZ�ں��7��fɅ���ԍ`�����f��|<��JQc۾ףO��[�;;�T"��X���Av n�!��� �i+Cm�4kP����$`��&�ʁ�����׹t��,���d���sS��F�]5.�^,�6�A��6�%��HN��')N��j�ˤ�"�:���%��+a�-��!)�&ap����N,�`RT�v�V��M��{��6 �7Z3)�2��$7�K�V���wV��tR�j�������/����r��H�:Æ2�֦����\�TwK�X1��*VhSDj:v�-��-܌Q�dy��c^�d#s¿��LZ,*�a+� Ě,ֹ��GN�D���AW��C�Z6*���w��L�njݘ%	3AC<�S�Q���G|emhH��ĸ�{��}"��4�a�?�CyxF�.c����R5m[/�P�_�
�K�9����<^�]��$��$EP:�ú�:�f���H���mISn5p�v�K�&j���
�j͹�X��U�;��7��(@�� �-���{��+��� �<�i���eD�!�����ϛ�a\$�+(�oa�.:8�5vƣ/�K�B'��kqJ��d:: ��	���Ħ�a�;��Zӥv�VLF�X"�p8�[4
׶���{�,��������Xo-LH���R#L�c[�5Rc�zjG|�GYtx+a(xݳ_�T.�������a���b�X-1xj�ǛJ���W_�����8�8���y�ak�ʘ��Xt��J�̕�����*{�2Մл�N�C��F�q�k1ڷW���1�t��~��e{�#���l�G���$�
�*OXE������L\{wZ/tPq427���d�U5z�XR*�WX�ræ�>�uҒ���6�-�^aA�A�٦���w^P�Q+�&�?1Rݚ{�

�5�K~D�t^}m�dԊ�����͖�۷,,����)�2�,�~�(��݌z�X�M����ڴsh���O�i�f���cP#�ͯu�ڄ���[���;��n�;|�M��s�~&T�ֱ/����&��w��j�wd��d�2��Z����Z�v��M���,3�>�;�ڈG�+��A	��n-x�i��q�+��7/��dV���mp�1�^Gv֗#Q�ӑVڎ麹������V�
�����'Y}��t`���G$I���E�qU�r�+g^(FЄ�V�H	c�ϵ�1��m;�'�Qbtk)R��oE�0�n�ɕ��n���Ձ%V1�Tu�m�׵���z%E:QG��"�*�r���'@���:ͧ��h%�j���}C,�vҦ�2��F0b���-�7o#��d���SSfEvӉ՜�T����{oM[x�m�V�482��P�M�by.�4�V�r|��%8)P�啁�yYyE�֝�a�P��U�V�) �E+�X�1h
�bjn�j+lZ�i��{�1���3^E[O������U]Ŷ��ߢ���#�#6[�i1��tri.�IMV},!��/$��e��f)E���Ga���#C����&+Df���xn]��Ut��K0k%`�Wl(�B�g�-+�,�n�$0���c@�hV,m8-�g֨^|��C�����x5�dj/6��MCNv�W{�X7�6U�
�P���1�&X+f���cb����m;6U8�����ȥ9��&ލ�.�y�ڥqfZA-'�Rgض���Z`�kd��[���V�Kx��ɤk�R���n�_nb�676Ψ4���%��H��RD!1v*���
�Q���Y~���r/:b��k��YV�m7�+��J���c[����/
1������	���46nb�}Y�%`ʁcmŢL��/R/" �@nV�E�8efS�����f,6��b��T�Z� ,^5,J*�X5�@1Qдk.��{j�1aj�4��"�*t�IG�t�	�rݡ�([���f:"Pnn��[◨�X�6�7�݇*�^ci�cU9��d�4^�ˢj�ц��	Ͱ�M�L��&8\�0��b�]d��
a"�&����H�jU�*��Z&���P�)"���Y�u�����P�J4T����(eC�4�i�u��h롆��;u�D�XQ�CKy@E�ڼ��ۻ�{@AS/4* �y���gM\�,i��L�<��bSj��uŐ/m��6��4u�#F
{��i���h'fX��r���5���G�-�����pw�wP�ez�ǙR�/d�Bc=����`Ș�0���nx�7w7�k�
y;&�{��PAX�7m�J���2|V�^��ܩ�b]�����QAu΢(���:�.��x��_����ء���5In�D��F�6�k�{I�Z�,���l�,T�pB�Z�F-���ZkK�po������@k�Z��,�f�[2�S60�T��]�$ut$
@,�u��ƭ�*�{H�#��h�T�ONX,�T�JyXƨ�zE0�]3��<��ǔ�F��]��Q��݊���m��v�Y-T�.�e��[���a*��%�&=�16��5.�~�Ӊb��4���D��9�&ۨ�u!��E�\Kww �6��[1m���KeF��k^7���&n�ٖr�b�qcZ�˽vU�e�ֺB::im���I���f���zH:qa�dհ�>�T�|e�M�V���"im�Ni!pSz/CmM ݪ*�����e�[h<CkY��fT��RJk��Q�o�&G��Q2��)�3������,��&�Q3.\@�Q��T�f(�h��GhÎV�ԭX1+,X�S6��,�W.�ϭ'Xk+n�%��R�"+s$�����/V�T~�(��M���Kp�2�ջ���M���S��xp�m����:�Ĭx��)���-d1j�B�e�{͎�^"u�ou��E�(;����f��GAէ�%�2����]��d>Wq�o�:\/4`��N(��X�i�e	XCQcV�ފ����,O��4+Z�E)	�}|����/����� ��(�+�n�M�W������;��	�D�i]��1V�`so���䁍bc���x�cD�VƠ]�3�cq�*j�wWjbŽ+0�˷D�e�C]`gAd��$#n�+��P]�E�����dǲ���Ϥd�}G����ӹ ��$F���)�Ш�F�]ަg��1��-�n����uj�fvXi�z+j�Y'V[���!��-���9�5;���%�ME�m v�@ufQ���t`+�2n/L������p�&�L7��7v�Һo
��)4eXU���2^�
�n�z�lZ�M!q��إ!�HI�F�yy���&�6S�/
�ݬ�\V=ےT�Bů�&]fAF�?1��e�$�݌��'���nU=Ebp��{R�7�Z���8죌嚎X�$X��a��7n�
��6��$��Е�r�=�Ip]�e�oV�fc�G�d�U���ێ�\L� ҕi2���A��%F��_��何r�8'j���Y�|Q�%�Z��w:?m�CS$^�Ms���2//@�k˲�hJ���ҤYe'��\�K��
������������F�m�#�n:8���.h�kw1&5o�X+�]����>��y�:�g���� ��k6�X��^�}�,�p�W]e�X��w��6��If�����לUo�+�׼'��Æs�6�mDo�-�b�}�����<�9���:�q�n��:�F#op��䚏=���y���WV,&�v][�s��f��K�.�����^.�Da���R�hN�,Cnq����H�ܳ�`�,#:\]��#rEҥ�	��ET-[��ں�8J�G�`:�W]��M<�-�@c���b��K'!GئK̘�jZ\z�wd�/f
���ok���1��vN��H`}��B�v�v:�4��:op�ވ$�a%�jqY�c֞�VH�ti[��=���Z�4��r|����hnvT�e�X�%�ĬՋ����]�d;��%|Sږs�2��{ʰT�r�1h��9�r��k4�En-j�
�l^���<o\�y՘�}pwVL]�5u�٨��q��ⱽ�s@�5�A�X)G{��c��w�T���H1 ���g5�E03�@���s�͍Qm:b�5��w�\.����h�SW3׸����Ì�Z?,�`��EC�Y��ҋ	vV��;��}6j�C٥�Mm�������F ��7 ;}�K}*r���]�w��f3o+��_ �{��
�z7OE���-��$�m�뤽�r���5���Q��k��[�7T������V�S_Z�(6��-_G��l�q0p��y{.�bdab�v�r|��b��^>�/.[bRE̷sl��O'�)
R֜��0��;��j�Վ��6_v�\^]�����xe�)�j��ѽ��҅�o�U���k�����u�Q2���G��e�����-{2�%#�N����\�!���Ɠ���l�ic��עfs1RB���zι���P��EGU岨��O��&:��T��ne<�ʕ�[+n��5���Q���R���I�:F%������8�n��q^|`�O�fY�o�Qtv,����3LY}Z%g_"���ٜwx������p	w��*��e�t�BW��`)ݑ���HL�3ZSn��5D71��Ųv���=�7��ئ��\ڪ���#�����i��{;.[[3� ��}�K���m`��8���f	��9`���3�d�>�6+��x�]�T��p�]��w�j��#$�'v��w��'�,�j}���Erܷe��"�E4�X�7�=�:4�,/�h�`�6),�;��%�	|.�Mn9��x�5N�����{ٛBɹ7%����.�&�u�r�Uڠ�=��u3=�R3�;��HU�' �V9��mvS�����0+7�ЫH��,�M	�Tq�Eޛ05���s
\�u4�}8>w��^Bu`��9�5ejyE�e��(^�@�&6��]
,vq#�ݬf%���o]�+�`��Yٍ���e�`�NͭW.��c�h@�}N���Ҝ�h Ȗ�O����lq4w�g<��uV/z��x���	���`Tj��O2���v.L̢�﹕ustJQe�p��h�K2=�j힝i�Qp��+���쮓�
֯l��q^�:1�[Jӹ������\���o�ڙB��E�&�|\�:�z**E��L��(;��7X��" ��w��;^�J!���|��4�Bw��R��o}�*n���YQeGv���}vW [�G�y��gm��_q��W�Wy�(;  ��ڎ����H��>�]��)�C��d<����\��v�1,U{q�]�R�@
-0��J�ë)G��J��/��gɌCYKʯvy��q�;��/*K�������,�BU�M�=K�nf�t�es<��N��2�\-�#}}�N
���v��N��GyC���}�#���Ɋ�pOOo�$o�	��a�r.9B慣��L�T�F=�V�1��5�_
K�zM~	�#|�E������č�B��o`�Eڴj.��Dֽںw�F>�ȩ"@K/�J:����W��K�-g>�m7ٽMa�v�;(�4�s�C)ө��gH>9}f0�eXHĬ*��m���K���ڔ��#������8\vA�y|.��rr9��S�Qȩ��AO�bU��,a�vP�U�̾yN�!-?�c�|C�\=���{>�!�Mgэ��t鯕b|z�:�y�V���.�hmcU��Oj���4OT���R��N�vsv�˼��ba�j�$q��\�܆glP����q"�_5����9�5��[�*�=m�@���V��v����)j�6FT�Բ�>�k"�>ŭk�ƣx>��L�Ij�w�8��[�=J�co���1�̷�C�����6��k��gxY��+^.��n����#���H��2�`�ָWT����d��6�k'B��A���W[N���wq�f��(��ӭ�3���9���$���#c�c�˾ݝֺ�mQ�/d]O1u#ލ��˷��#�����|DO<���1f;�ǧK��(��X���!��O�|��o��*�[Gb\2s���T�ߠ�+sM�m��N�ne���ޣϷiY7�K��l1�g�W͇�lR{\�b���ʥ����<W&|��\a8�$�XV̢�̈́S��O�&�wٷ�jr#]ۯ ��S�혛׷u+��
Q�Ѭ����A�f]�����m�|����<tP��vTz)Og'Wz�lv�(b� Ȯ�3�ݎ�ɕB��Ǚ$�ڗ�|��{�u̝����NB�.s��5�.�EE������#3P�����b*�ոE�m��i��K�%�HЇ.�E��8�]�[Τ�u+y�X�E��u\�$A3S;�i�Wwŝ�Ct�rfGs��[N�:�YZ� ��Gq���'l��-�u�%������<�c��j ��#�V�rⷍ��u��)mLÄ\7]X���M>k��gv�����t�+��d>"��wq�����]�Cǝ;؜�:�HИC)i�Xݭ�w��5�e���ݎ�-���{P�ū�D��qu^c�_���W�L��h�;���7&�a�\QNx1�^f{��N'q4�O:IJ|�e]��yR
���Ω�A�]C�� ��x?�g��
Zh�AJkFm����j)�:���ow�8.M�o�Z{��'I]��f1�ڻ4� �O��V���S�+���^*J哹�dn�%�/�%��w�����}�����e���n<`�bV���ebl������$���n������u鱛t��Z�_,��J�b_R�ȥ�P�����p�������͍?�X��Wo��V��㭩BP�;I�l����:��!ȭ�vo������ԯ
}�th3/4�l���zU'_�baг,��IZ9j�7�A�)eA\�R�@8�o p���
���^��:y�ol���{f$�����8�w����F�&%.;�Ի� }�e3z�wD.�j�MRpv�ʶ��D�v�>�':Ń��C�KK�:��<w����f1M<���-T /Z5�tT�
7WM ,B�b���6�v��ҋ�;�^jf-+�UT#���:hX��w������AI�O�5��'��Ūc*-���ewH��F�'a��+��Ԧ�> �Hγ���YG�j���e�2(q\�ض�z}��v�師�90O�
&�cE$�`������(�|t��
*`s�5pf.��wH��t{�����fd	N�z�;�,!� 6ɿ��Eݣ98��{Z�	֧%�:�n_.�F����uX�Ǐ�Cx�C�gt�b��w�'k���86C�0���r�Q�s���O �R����oqY�Q��U���GW�CKP���tk�\��$��p�³��¸�;u�ZGSC6�vD[-#څ,�iN*�;e�"�w7�Y%��N�b�h��N�Y�q󹱥�V�gWt<F��Z��J)��2mu��as��
��z2�'��{��2����F�>��i�'��	�^�������^�E"�.��S����y�赜+��-�F 
��3%Z�XV �4����*��O�5}��I�k��7eR�:@�T�iɫ��`9`IKxc���n-1m��.���7��� 	�����h��Ui9M!�Yq)��:��ⶭH�N�O�^�垠�O6+�"��Wywc� y"��������zl�wg�<bJY�\��}u9����Nn��MZ��x'!{`��,�T�3I� ��|�]�)s׮�,e(������O!Px�/�9�N[�O#��aj�]ܼ�Yd�[G�E��]m�u�uzV��k�_,1vJ��nt�e��"Բ�d� {������#"\����,e��E��=Z���*��Yr�ɔ%Y�wB���u��D�zy���&��v$���l�;�ZYQh:�
}ʮ�u�Q>y&c2o��.�at�����;���	��� �n�b��4.<��jv���Xd-`Vٷ�8�J+2���"-���*� ���P���
-���]�rA�d8���6�bn�p��f�˺׵�W���64�s���:J}���Weu�ҧ���V3��0պ��� 젴o'v�Zy)�g�1��e�C��ZP��ɂ��;/YjݗA�{ׅk�8L�౹���'�r�9�P���j}�t�[4^=B;�[�4%m^H�ƚ�>�0x�-Q��k�9�D���*��S ai��{gg1��f�ϝ�;ѝymKݸx�1����®"r]�g��m��1αm�aJ�ĬmS1���xVS�X���le��m��}����3���0;�0oL��X�Q��bؤ�>��c���:��$I�8�4��]ݙI��UnZ��͵�y����A���puc����Q:��WW�`�ի�טkV9��v5wZ������ΜYRh���*ۼ5��]#�ΞÚ�2�ak����,���둮ʣ������`;��p�X�Y�4�`:߭�d\v��C(:͗x����M�5�34�Ò��,f�tg/:,d�z8�}l�wxJBZ�Y�bq+�bƮ��菘��.ѬH@�V]���5.�k��CA呫�5$��9��Å�!�즋�+-LU39��R��kП�Mk�AT7q�i5iW�#^��OQ�D�g61�[�L�'��֯��W�Ҟ�t��Q0Z��.�Մ�r��V�#��M%��}&�`���t\�����1R�R�jm�=���^ ʧ)��}����h�Ƃ����+ �ihlѰ_�����K�v��(�R
����2v+�l���V�[d��v�͠����i>���m�oz�r�ݢ���ژ�]�[�~�{�o�7Ka/s-��I~�i^���Mg%C��K:&���wI\���Vh7���E[Zc	�^ c/D�e��n���x�ְ3h�p������ea��9_[]^!oGP3jˬ�P�>�ˈgflkmXR��|���V�)�\��xqʗy��Q�N�f�Gt�S8��S�^������,_Vʊ�$��ھ��g%�d����|ydn�V��$��Vo����y���a�؀e�j������/3<t/E�%�8cܯ.�b��.\�dz����3����֣wP�}i�X��&l޶��k���@���8:i�Z�g�[��;(qS�(dɳ,6���ى����_�5��	��Krm8�����f漳7���4��ۻ�^^vP/e��El�T���k�vpb�����u�^��F���)6YV�x�nY�Eb�؞�-һ���c��N}�KcŰ�U޲�����u��ݳ��1�y��;��Wa9�8���*֟���;�Uլ��rS\XΗ�x�B��w���ދ��:餀��v%��5E��YiU����^B��8;f��Mjr̺]ɰ(	P�A���]KV`ߟo_�opN��l�����aB�c{S�n��p���
����u|_^�.�ju׻5F�M��V��;���
�K�{ʌ�I�����}��9y�������OT�w��rC��5�{��ʛ�@�0������B��kE�y��7��w�.���oV	��z�Da��X����k.�:�\0��[C*F��n��΋7Lؑ
���bSy��yB��	y��uK�R�5v�\����F��soKޤ��d�L�s�R��)]B�V�vƸūp��\��rg����/vM��/��K�1�c[�N��z�Ig�r�6ħ��E�������8՛����s�)�5���֦74�}Xy]dqGZ�f݇�4��q��P�m<)`�uhὒK����S�=�cz8t�}��[%�Щs���ib#R�9�i�Պ�*�;�܄��W���V:�\۷i�p��.N�#���hu�v����-gD��o�g�\���A@�AU}R��8z{$��׸������Üy�5p�qİ��y�"�[��u9Т���"x��p+�Y&��\���z޶��f��(a���9��+�jj���N�B��	/���Ut/���*qx9)7"(���S�ps˚���Yy��0����{��?W�l�=+'p�����x�x2 }w�����uY��F��w��^�`�]��B#3yX9�ٹ�G����8EWho���f�3�*�/Pє~=�eʾ�K�����\�}�.�������'�u�Y�0r��_Y�O]i�[���u�u�}3�{���gOp�z�Y��h�Q��V�̗�m]��Ӟ>ÊgF��\}G��y�5�u����e���o>��޿w���I@	!��BN���w���uu�����5ۖ�����jhg���䦐�l�=�ՙ�q`��e@����|�����C����,u�w;�_;q2a9�!wo׋�k�&�w�{�W\��Jd���"z�f�;Wv��
�nl�q�t���e��7�n�f��D�]R��o(�d{�N% "��{~��{�qc��R�k�>�o�+.�F��,��z8D.bV�����J͢&��5��X���9�o]��GpZ��%�-�&��v(���t&pzzD����Is��ܡvQ��+�G) ��3�ڸ�|�P){��]����jƯF��2,0�.i����N�7�Qd��It��m��e���f�e�k��7�3��F��������K���K!]z�ի)���kH��m�v��k�tC1��%����q��;-ZX}�En�b��k$�$���b���V��#`�%���M--ϸ��-��mAWF觼��n���)PΔ�'��޻�{u�)kq�U v������)���X�w*�K�	bJN�+0������w.B����<@�]k�f�N�%�O8H��.��;%8v����\ؕ;�@�:� ]�;g��/�ki[I�x�;���t2�v^����v��ym��r>�=�QϹn	����Ղ��b��Ξ5p"�/m�E��$.����;C��8L�Mx}��8��G�UN�=�z�:!U��&n�O_M�w48/aS������Qf��s*��g!i���6�Z�\9V�M��nL�$��ﲶ>��v������GH���OW<�7YSR���7�^�Լxe��ż-��˥N��g�Sj��"�ֶ���u4�#��A��e!��H���yj�R;A�Ԛ�.uquo�\��� �ي�;*N=�YA�u��t�t��cQ?3A`K�>-\�j�mg�O뫛�����k�t�4���ݭ�f�IY�3(��mf�OJ\�
��l}9	��^$ļ��h!L`��G1-�����rb;G��Q8u�'D�7�C);���[E^d=�f����m4�[�b����w1F-�����&�sa�Cy�w�������w�K�9tX�4j+�˷H:��8���ӭH�o&
�(��N�M�M#%�T)V����W��A4OI8Sz��Ӳ]09b�@8P���ZCt�1R�fl�g���U�Xi��=�jnVv��d7GGtsmmnou�ĩ�]��K�01�\�e�E��Ozܳ6aN�,2#�S�d6:��Xǉ�@�];�m�H�s���H@>�EĶ�n_`:��î�.rU-Y��e�ۤc��]��
�����!k���+�l���)��}-ۧM��O���0����Z�D�ѡA�;b�ft�����B}�,����KX����Q�P����1��FywD��3�nOUL��e�a؅*A�����%��F�9��q;��xL&a�oR�;����2Uٴ[��h	P���K-���*���4���Hq!o����X������E���Ç�A�R֛̤o��r�G໠)��Ԛ���n)P�[�F�9Q.n�%��k������`�
v��E:Ĉj��Y �l�6)�կ��"�;c���	S���깐����Av�9���'d�q-Q.���YM8�t�%�3�c^�dIV�eoL�˻ծ1��hg��7�rث��q�[t��nb	�FAL;I���S9��of�����C�ev��zo#�m��wlv]7Y{}��>��.oo3f���9S:Z2k�0%�j쵦�0�ٽeл�U�9�б&2�V^т���݁^vB�[�΍\�Q���k� �H�����9��B���'�!J+�5�9A�y�y]�
t0�@�= �&�#�h<��E���	۹o/)D��EF���4lI���u��껍g)|4T�J�x�5�G[�'��V���݉T�������\[w
��8Rk�k����J��@ q!���]�Mփ�Շ�քs/2�@�i[�;�'�LX5fu���gυZv��N�2��V��Ԯ��Ylu)5�׼B?t:����:U����פ<��(�e�3#n�)v�^ �g+ߑ�W�m��'vf�4c���#X"�9��gM���H��|�T�M&K�2Ѳ<�&�2�(���χ{�������zX��h�����9-��+��]<�mR�3.������]χ'&x�9l�����l^���������A�6QG�N�)=0Ok�u�=6̮6+�v�CX��n�c>�}��E����48�Ǎ�$�<ܐS�s�`�.f��KԺ��=�Ǚ������j�L-m��dż`��up,����*���|#c�_�|���tF�*��	]�ב�F��!�N�ST���I�}SԻ���F �����t�m� �p��^ty�+X���W;Ḳ]2�׶`��m��9C�oW'�q���i!YK=���/]8���wCF�����q�^P%�1�{<ǵa���ź�R�}3�j`���%ם�9Z��SZ{;�
R�uD��t<����`�U���a�2@�*��ջ^�Щ��|�
$���� �]떥�k�X���$�^����}����u���[ʐ������T����GlM�W����nfA���r�Z6):$�2q]�ڼ* �sX��S9���\+�d�]t���\/h1ս�a�Tέ�F6�Wr����r���7Z��L��r-�Rk ��vۇ3/�F��qPt!��|�jv^e��Y���D��	N1����eX��f�ek<�`�zk��(�1�4 �D��c�+�x��5r���q���BWc/�٤�J�Q���v+e�[]��Mrr	�>�9ʨ���ۃc����a�0AG�ڴ�BWvӉ��Luw��gv�;�.��Υ���]� �K����E}�F%�o�WVX|X��{\ӹ4nx���^VB���/��K�=�B���`Ĺ7�����g�W�Ws��#gd�!�Ѻ�K�ᲧR,F��(�c�@��5��k��N�=�run�mv\7���[el���i٘�pQ��"��h���٭�K��gj��c��}4�m�<[�{q�5žq��F��úFۅV�vl���aw:S����sS?��b��WZ��VC��GU$�X뫸rvԡ՚ؠ҈�&�R�s��|���:Q����Zx��g ����^��ޥV�O,=s����0Q��k�����E���:^;��N̫%��Denq���H���H��ˬk�upp�v]p��k�$��m6�z�(��ogaOٌ"��Qń�B>c�C�E]b�P��>����lt�;�4�eջ�������N��л��;r��<]�bt���o5���l�20V<�hӛ��W4-��,3�zǷ¬ă�wa��	�	�,�:��Z�JXjgr���k���%�
^ɕ�n�	��#$��3�6���ٜ����R23�:W�\�/��FX�9׫�d䄔����:���Ŷ�2�庶��w]�q��BD�^�J7|K#�v��,=쭿�4���[qaj�^��@kܺ�Z��lJWyaK'��;��+�o�1�f˗����kM��ҩ}�'^�7}���8��-�}-���)<=��,v���v,���nt���4⺛�,��اYUý�j������2�Z���c����B�K�b��C�����oa��G��H���xݠ"!=��6�hv����B��ts@V�=lf�W�u�Ivӿ�'���=]sjG/�Pb�b�W]�u�]Ň�Y��������*y���u�1 !��,� 2�<X�3E�ϳ��wR96J�,2�
��qi��}��5v�[�ք���N�U`��{�o�%.9�C����R@,���z�]Y\�o!�'0:��fKOy�E�I�|�zu#y�ǧ)�	O5r4�����ԛ�0:�U(a�{o�������]]���G�I;wn�U���$WoB�迀�����l�y��C���z�mf
�l�����̌�U��VpQo�g�#�%�W��Kx��mww��4y{�ꔈ����;��A�̯M�3/>��
��,:�%Q��2ݲڼ��V�w�������V�,+)U���*U�K����#��@7��.%d���p�G�MY4܀* ��]�ѡH���]��\��_pn�S���c2��NV-췯�G�뉌ku'S؛!��e��f[��T�xĮ��aA��r���|�!���P���l�O�h��F����E,[������M�{2�B۬����n��6��+��^��*@�D�I��܇oi��/[�f�S!Vع�nf��tgo��^����f:�5ۯ�6�A�������A�C����|��v�RwD<Nj��&Sr�1s��g��6_��j��^+����{Gs��0)��m [�2"ǵ���=�H/�d�n��U`��T��G��p�Vސ�Ǖ}�۸�}���R�MT�Ԥ'[R�S��B��U�(Y���cln=.��D`>�|,��cT��a�k����Iok����׳V+����+���!{�P�r�|�Er����/�3yń���J��;Di�,^:Y�I���7%&������k"4n�����D$(�϶@�W����/�}Xޅ���h`p�ڝ��Eۼ8�;�B���)ǑB8ƎN:.I#f�	\�������۠�SDm�!	��X���⩚�Xh�4I����Ȩ%;^l���?��t"���G/��!t:P���n�M���& ��u�Vԛǧ./P�2����ԃN��X=�ýk{�3Gk��Qt�kR��C���������Dy�WBT�M&H6p�47�ч@��B]0P�}�:�+4D�o9�υi��>�V��~�7ܲ���Srzfއik'�m)����:���{�� D�j�p�}�F�0n���{4�3��9��`ۑ� ���a*'{�m��%6�S������])����Jۛ`W �5���P���-��8�*�Ls�!������2�x'��%�k�B餬��h#z]e`�1�Z���	����L��KAG
6��mf}�U
�&��CYغ���=�	R�p�8��t˵4�fIX-[�s�=�:��Jw*���=Ď�rz�_n��2c��RU��Ȯn�;*���)ݥ��q�d!p�\#E�;WIu�[,-�et}��9I�A��f�pD`���'uwǠh˰el��Ĵ�KK�4�s�� hD@x��8I�ۇ5#a�p�zq$k�3���.U��1q�݋*�	�Iw-��8�-uf��*%��eʽʾkQ�{PN"��P`�NW>�WfT�f�5O�=�E�X3�}.e���!�S�Hf�J�jm�/�)�d?LgU�u�:#�Rh˝�gr�����YӪ�[襕{�W x)S��a���e%��;�B��W��{:�EL��2�C\k���=nɅDc�������hǇ�,ξ'�!�� u�Ü�.���V.�uGzC����{-�W ���T�6�va7�i}O.�'52�'x����2U��N������>��cP�P�����V`������5�ۭr��E�{׾����NL>�W�v�G�c'vWF�X�CN�_y�K��(eS2 �=]1�k~+,ve���]rr����H�e�P�}�i\i�nجo�q��xz]`]�N]�������"�8�;�b�'r�J�o8�o,�ܼlVF�iŒn�vz�H՞�S�:2n#�����)�������A�L�ۛ81��m��3�9c�`N[Р3`Vò�y����J��yB��@����u�	t��h����D90�vq��V��Y�.bv�A���{�d��"xH�-]ۺl]��IgM�i\3���@�Kv�t��Q2c�U�JbX*����ƞS�{��qs,̘�uԉ�R7�-�> ���v�bU���7����1Jcf\���
WR�Q�+S{o^/�$dH&�h=�*��������eۤс��-ū\��+E7�L̳�\v`!Z,>��N��υ��k5r�ֆ�#3oI�>��s���]Ē�
;C��p���ܻM׾χ>ZC���x@3��2[��d�s�EϷL�y��zg\��ܝ[SL�f�}>�k�ys��:�2�7�1֜n�'�8���/�c�@4Rt�RM9�I�cIv��Fr�<�d�^=��Xײu�P.�9d��sRCz��������*̷���x��+���� ]C�v��"ʷ�����J�!���7\�g$�dۄ�����j��nww5r�c�v֬�@wR���=̭Q�v5�bӝ��SF�+Rw�I;����=`^��*���`�8s]f^|�ӜE����gH��ʘ�*�{r�ݘ��\����=1���ű��@�6��-�V�c�}x2uCE\9ܱ��Ε��Sj�Ar�uXy���v�ݽ�ie�'��%�1���'�T5|���A���>F�#�����:7{6��{��Ij�4d�J�T˥��g�hZ��2�"�8���N:����݈w/b����m-Um�_2B�sxjO���<���P�������`�	����N�ʂ�����
:�mIWuhcz����g.�V��+��u�m���=��Q�f[\e�t�\-o*y�Pn2�N�� ��~_,�w͂���L,���haf��n��խ���Wv��\SeN�:�V6��b��s�u�ԕ��%v��o�#�ٺ�m��J���0����Ӽ/|;׿����BN��<����=�r�\-��t8|m�\oPݩ��0�cܽM{��{��.5��!�%�n�u?.L�]L��IX�����k8�����Y�-$z�X����s���YgpЧ�`��,j�V��Y�;$F�ZQ��8/B�2uu�Őz��Up�q�͹��t6�-�e�C.��q�����ڔ��n����R:4c�R�;2�kA,�g�t�4��a���'o��;T����M��&���-��ΑP�yάv&+���\�r���d��
�y{��S�b����m��-�LWx�g@��ۤ�-�%������ې����ՌV\��vv�bo��4b[�� ��7��C��<��m�O99���9����u3�2�G���/"��ht8+7�UNRE����'��B�ұ�.�9�7%��౴����ܜDy������� w���Vk��|�]� 0o�tl�-���I9���N��V�Ò�}8`{ݤ��+CB�(���ܥ��$`FR�V3�1z�}�Yٌp�݋�� �mv\۫�}H
5�#"��w�,�"�jRɕz-�mv�=Rv�]���E�5�(��Y�b��jd�B��tR�ǹ��#<����]��)LC��O���c��x�����0�
B�+G�����.�vhp�G�B��i/�5C��Y�(���mU��6�2�	S2��D��9U��b�YD�m�5����L��Ĕu*�G�[h�e5,Ac)T`�+[j,EE[\a��u�e11�Qumu+�,dUQA\meJب&�2�(�9ewK\QF���"�`�T�6��m��1E-��UE��B�Ԫ�(9J�����+"�̲���k*��b��!���Z֊!�\�5B�TQGm��ծ�YQUԕ��em�DV,TX;[DG�1Ĭ[Z)�X��Ll�1�k��*n�c��m.��X�ZT���1�ҙ[X1�v�i**�V�bTS(�U1��DT[K,DEQ`�FJ�73w"�h"�1��`�`�QW�mLĥbj�.%�8խ+DPCI�AA 9�ܕ]J��完u�xq@�M��I_|�͂]���wu3�O^���2D��BY.�����d�ԸD�D�U�^8�c���f\���π_�v�)���\`��,��]iʗYT_^���;�������8&w�s�ѶWwT ��x����`�ڍ�\���F�1��ʂ�N�36�w{�$ng=�q$��W��OyY\X}�ȩ�=c��A�s��z�²�pk���0�Wr�'�m���m�ъ)u/��ʠ�i` F�XZ�!����K�K�1���R�S��|���Ҽ' �����=��9��.�O��K�h���<2���$]q�������W+��)��@�����E��4� L~��/��uk��{�0#�֢�j�eV�wF5Pt��G��=�hq��l�w^�c:8~x� ����<Wr������P&�ig0�G�����WF7����.��:��n���~9Vz��}~���v�M���2���^���X�b/M$�h�'+����� �+u*³�~�+Ӱ��}u�wN��y��Ϥ뵵�C�y~�h_���p0R��t|v{��QԘ�l����� �fX�;.:���O{�2�D���B�}f��5�g��K�S
�R�#�����o��=y[p{�0��s\p��-�����K�}my=��{���g%�o'�h�(�x�z��Ꚁ�d�{@������/h�������U���#b�6�^̦2Y�����"$�,�$���K-�^��^dN��1yn>�:�,͵��|n���ΰ���k���=�ok��Xk�?�T�d0����1����)-���>=C���_x��fo��?U;`2P��T5���̶k�B�D���Ǻ�o}m�H���5(U>y�q�7>wc���^k{\{����&�I�=|������t��I�"�ltYb�*�N�P�H��2��͓�mJ�s�N�֨�ĵ˴k�Yk
�.���/ 5׽�C����: �/�L�U����ު���ny��,�:�Cc��i�>�a�0R��t~D��htJ:����{2kW�$����=���v}U�W�6������^�
S�-�<�;�h�p�G;���c{F�Wo���:��9>�V�Y���p�b��� 8x��(��P�y���'+-����2��n�y��%R��7X�'Ү*���x�� ����jU�(wNH�wWC�4�Rt����4���֔�X�ս��@�C-����gB��m_ecv�t� �cݻ����4�9�Kp��h9��-��3;��b��r�Und�Wk)"\��Q[�޵0�t9�j�ފ"��c�d�:*/m��x@��C1.�fZ���$o���=\�/�r�u����Dm�؈�W�^��Qo,�Y���+\�
�-��(g�7�6�
$&O��W"��/ڪ�7KԬ`> ;��aVNyW兟6�u؝�X%�L���d�v�X�Ĉ
���6~4�� ?p�u�g��x�i�j^�w���g{�k�睨�5�/��v�,wp�p����>��x�Z��;U���|>�V��5�"��'�����T�"�^~����,O�*��\7׎㢐����k���8�xEc�z�j��tm���M�^H��N,���g����[W��`Fs�Z\+Dy�_ܫB�|�33畬g����>�Q#��WGǥjt|��W�3B�䥪��/m�5�z����Ha��w.�3�7/9��pz�Ԭ:�\����!Ҭ�;��@�9+ѱO;(T�ur��P�oշo��v�S�:fW��/�+O�6:��rJ�AB�X�d=�g�E-Y�ö �*��r��/�x�{f��W�,ǃҒǪ�^:��U������m.�)��ʹ���s��it�RX����K���r�3�!��h�[���w�F&2\��m�ܐ��:�F���G�rf`Á��a��с"Mѷ��!Q���F�����012<��.g8ֱ�jÎ:�J�l����A]�*�آ��e��;U%u����X{�.
~�́b��|x]��p�F�+�m��V/0��
��w�Խ�j��@�v��<Ϸ'^'��6z��g@|�Ū�e���~r�]��.4P�E0A�j bv�&�^���'o+ɘ[�f4m���!���e��bJ[�ܷ�pU�7V��^���+n�<s���L�~Rg�p���.�^�tB,ۑ".��fN8�2���e�$)��������������q�x���Q�c5�^Y6�ቋ����j�u�8�׷F�O4Y�?���6����KOs��	��g��>suJ��yU����{����VУ\.��{�]w��o�w{6�(vӶ5cw�i/a�'�ǲ�0��~��d�_ �X𧼽���U���k8V�l��!̖�u#c!X�J�7F=� �W�/�
�$p�Y��{�����>☽��Ef/{���7�ݯ�g���A�!�;�K��U;��>$oQ/��xV�&!�pc|e۶�J3wi�$ZZ����E[p�}�`>�ą06�ӥS�o((��+�W�uj�:��o���ܒ�E@�q��n�!2��#��1�v֬���r���(�.o'Kh3�G�rN��Ng@����)�E�8�����D47����a{��$Ng�KX�Z4 ί�B]X���J�.��<������]+YV��0��}�RR~�x�<vCp��a�R��w�u�8�2�@ܿn��3���q>��q����>]4ZD�Zu1h�c0���g��t������q�s����b�[PM�n΢����^a�/�T]�o�+�lv'��ZX�,��N���̰6�N�Q:BMI�C^II��Yq([>�	��Z�hX�w.4XC�@5�۲�ه������ϩ�p�ދ$����gܲ���*f���\� �
��j��)��׵)�	�@b��M\��ݳl7C�F .�6�L,�����k������W�y��og�')�+��w���z�v(ea|].��� �5�R�<~�-�J����K:�+;���r�d�@����-���}L�m��=u�l6 �ui����dY�&���m�V�z+�B���u�}��j��W*�
��f��E<�r͊�K-�c �uP\��MoLX�Δ�N� V]�xQV.}�����D,W�7-8���Yd��T��V"�ձ�@�BO�7�rp���܆�g@�u���&4�k����`�eYe扲�3�p���b��.�����U�����Р�봶�7oY��]q�R��"��V���chT9r�$�ǯ<J�֖�f��Z|��y��A��G��ڒ�~�Ͱ}��B�w�>�u�q�5�	�����s���+Frϻ{^U�|���v�8W���	��t�V�΢Ŝz��T5<Y�zKR45�i�B( H`*��VY����� �߫�)�	�E#,���,���WNF��ס@�6�����ܕaY�|�;�:��n�ٽ�.�"�x��s�=���R�ׇ��Po���� �����Q��w�U�*��Iü�ܳ̓|�_��ì�ʗ�}�*�D�	'�4�:6=l2Khk���R����}�K��)B�'a��*�q����{_��}�.��YT��ʽy�4�Q(�"��6-����%��>'�{%l�h����փ��l��`�Q�6ٯ����n,��ʯva54�p�c�������q�>��+�LY��iZ�ݏS߽yZ��.���đ]S&���k�O@�iP�?�PS��"��gm��](�4��ǻ7N�Ԩ�܅�_�<ɝR��yOo�AeK߀�u̳�2R� C4�`� n���@�:�0�S2��b%�8o���;��91i�oo��[Z���Pg���l7I�����zfD��w%��Q�pK���0�`�j�]��nԖP %�]W��c��:3gnu�ؤ��i]�bu�p��z��+v��ؙZ3X=zM��k�����.I�n[�u�R�[������Z?{�[�(h�U�:�)����"s0X�@����X5���{�nn�����N3�a%��M;��X�X�c�����jd��<���q�GUxzP�����/�s��Ӑ�������4��YE
��ceu��<jG�<O�א�.�����Nf\�z���L;���r��e��硯0��>��j�:���h�(m�8��^������5h�����0Z.�ʠ~�-`����Vs�h��ʞ-xX�^��w��o70���
�V�]�w�i���k����b�����]�"�
o9�:{K�KÈV�����7���r�^�0�����:PZ�|���_/z��~�a�-A�L��TP95(��xJ��U�$V�2l�F(�L�A�w�4N��$5k[���:�����*�=��9�+�2kEC�t��ߪ�Ѥ=C�i��,�}e�iWO�ヸ��LOb�5�)I�����w���{��}⊛kG��pS�Ar�ʫ�-(/��p	W�
�1��δU�u�G,r�����Ҥ�{���ߔ��[�^>%٧C�4߉��6���ܥ��EZ�+d24����Yn���Ӣ�(5"�Hp#]e��m
��/�Ͳ^>f}�����c8b���'�7i�y�!�/�����o!��ac�<��E����O�y�ci�g�Фw~X�;��+�.d��~�e����s�k����]1��O�_ā܇�Ʋ�j�<]QN�R�ws���g�Z����-�I�/i��E2��@*vq�E�� �j�� 43��u��N�����\�O�����{�*�]q��;ưV�9�FFu��𿼩W��Z;,t�0'�.�o��z���@ｻ>���j�xyT̈zQŪ��~<���T�%�������X���0�sd1�#A�Ԫ 
%Qg�N�����"1>39dEa���1����u�[�;�˪#ݘK��R�n��|����(��^V�A��.����ߺ�Z�J��}�r^h=G͏#(`i@�:B9��Z�w�����'0�Z��mF4�E��6�DӪ��m�ɻ	���� dwA-5'ˬǏ'Uxv�e����������V��V�ء��'�0$��E����*t�CQ(�ȋ:��7V#V%}��t���7\}��;��ݺ��}o�B�3H�^��.n�������u�X���i���Tֆ�/�8vP�-��5�\Z���6�zčF(
X��{���
{ �:��+����y�u1:Y�gpDq2��]����Q8���.r5���):�
G��y���+L��ػ�U|-ˎv��{6�L���;
����}9�<.��0��@_JƇ�k�ـ�V�gg��ŷ8!�] �������1�Ld`]mә����ڣ����ty�֍?i����z��#�7=�>��~��p����Y~Ce���n��v/O�N�)J$oQ/�."$+Bh�� �ӱy��v����χ��[��������sK��������U��x�"���q���;�m�K�Y�g*q�ǐ,W�0}����{}e���>�)�@u�����g����o���p�����#Q��h	Fl��f�,5����EY��Ή�<��:3P�[u}�O޷;��H����W)��6�J]f�Q��NKUǴ2�b�=�y�k�v��J�h��ҟwlS����	�*Z;n�F0O���%�M]�<<�a�)b�C����R�����0E5��w��O�	}%!�6�UJ�>��(ȵ�pũ�'r��3�UO���v� �`� ��𛶩�T�Ҙ���� ��R6�)�	��d}h����ޫ�0m!�z�^��ҍ-`j����f�r��J���j7^��q̔��H�mX��5#Y)��2��Yn�,R�l_=�ɦ
�<O{gY0{I�Ĩ���t�!ze���ZF�Y�W �/*Y�q|Ae��.�w;�yL"2�f���e���ʡ���h����)�5uwL	{��<�j��]�o)�.Ӡ����V���v�Pp�Wbp1}PF� ��D̲�������f�s�6���ɱ�Y#v�kx.����΍������ģ[�*F���,A��aa��n4�'N��O>��c��=C,�Ɩ+�O������B��ó;4��)�{/�h6�M���=��-�oS�:<��{��p�KrV�%��Lw���E�.}�����Dz�x�O N���o�]�5��z�-Vg6�p�
�۟c�R�S&F�)G��׮b�	��NM�
�ȕ���E�t�f^��WwDp�R���U��������P�����_n��+���.�!fG'w{�*A��{dl-���!ze�}H|����<�X:��}�t��N��L�y6�ֶ6|��O-e��
�|�S�����G�:���}K���!-�zfVbU��b��'���;�����\U����<=g�㪶k\�t&�E���ھj�|{X���Xk� ���^��l�i���z��!����-�闗k���w;�c���}��mQ!��R�]Ñ}(�� cteνÂ�cv[����{g��'l\jl���5s�,�]Cb�aA����PG����i���x����z�bmv���:r���$��ƴKqf�f�;Gs��Y����i��>����ە�����B ����2���[G �/g�iݜ�[";��e�,����[�^�	^���F:�k��-V���V׀^�5V����S�:�eӎ%�[A]��NΔ���h������0Z%e.;L.C��t�r���Eu�m]}���\cVn�"���k5�����@�urP��ux���*]�KXd�[�(��V�sՓlv1
5��v�d�@��Φ�/5^N��kI��|���
`Lᣔ.�(�FU�/�q����x51�1��٪���ܺ��//$
�M���9u���������i�Պ����*;J����s>S�t����G���ܯ�\�o.�{�~;ܰ0������k��<�X���K2�N�����J0jC��h��������~�Ԯ���&qhy��+��V-��Ooz�ϛ(W:9:fu�ƽ� 9z�W��i���zN l��墽�{��ؔ�*�oAS�:�����;A	2�;�0��i�`3�*�QѩI�k@|;�:9�}J�.�����J��p�9�L�Z36s���x.[\/y/q<)�w�Deh��Ɉ����:��,��b"KF���~˥W�"�[�f�2+��:+�g�橃3��@M4o���D����'�W5�;8�{
�\��e�s9�z�鶓X����� �ΨU>�Ñw�^��{D�_��-��'ݽ|2w���
va��L[oG(ç{pf�X5ծZU��/�I��&̑Wy���8C�M.��G���	�
�b��d�]H��5��z��o�wGp�wg�n]\s��'[��Ш=uzdn7[��WbS��݊�̝��m�vuA�ݵL1y��:����V�wB�E�3��64�#���&IÓï��Suv9�5Qt\�w&�K6�����ψ�B��lZ~�|�)#�֞X;OLҫ��*5k.�[L�)3���|�x��ۮw�s��2�sF�"_
O]K��pJ���'!�E�(b��jlen�ӍY2����{Oj";�5�����V��glǥ_q���Qg| �vC�.]ۗ=ʈ0�f���[\��h� b�/
��jg8�fR�����2����+�m6�[Z�"��4���XNeM.�����\Fa������ﷻ�-V�X��:wF�w.V�m�b�kVlN�hb4t@{f�P�R���S�Vi���9��T�̴�w��[�v
=7�˗o��7Y�U����|�<���)�l�ì/�giTi�}�T��HV<
���q]}��83� Y�OI�0����N��;;<g�*	���/�w}�x,5��<ҙ���
����!)�w0��7Π�(��]��Y����=|���[oMW���9,t�[��L΋ ʱ(�O���w���U��U�(���ʠԪ
�Ub�Q�V����b(�ic�EDb�K��ڦ� ��e���I�Xd+\�X�#`��bUb����c��
(�8�1���[���[J����V
�m��bVQ�j*���#mV���Q\����KD���1�#YUA�U���+dX����YԪ���1�W�Q�A�(���,q�(��V���ZX�����QU�*H���@X��sUТ *Ȣ�Z�feƵTƪ��%�E���VZ��d++	m�e����5UDm%V"""T*�UD��X� �m��eh�Q"�h�!��)Dƌ\���̭��V�%���R��L�Z�Yv�GSr�UYQJ�&"���+j��5(��&+�jZ��V��dY�AV"�ZP�G)Q�����`�Ynd1��
����Kl�V*�D�R����(�F���&��T4E;���Ykn6�ow�%�w��X�g7�Q;���i,˺8�vIBX|�f�h�㛑6ws��g\��x�Y�&#޶E�:H*��H�>}f$�g��@Z���~� jV����x�*T9�;CU�*L�sP>K��9��Y�J��T�)�M'�LC��^{~��w��?nox��ja�k��s��oZ��^��[��k%g�nC��=N�%I늁�{«0�<M~���X�w�Y�'h�I�e��P����t�yzH*��W������U{�a����b��f��aE��8fY��Ld��ĜB�=���s�+>d��Ϲ�t��:���v��+:>�'HT>L}`_3"Ɉ(z��<��H�gi���:�!^2~�;)�~���Ϸ������zv�|a۩;OS���'g������ ��v�����no�������'��%eg�/��:@�+'>ܚ�ĕ%f��*<B��p���=���8`=8�����I��J�h�X��d<G�G��s��gbMqXG0�!��!���T>I^!��i�����M����jAm�'��c<��&� -C���� T���5�3P�
�4�ߞsۗy�Wx�������P�
�٘j�W�;N����g�*��(q%|Md���|��_�C�'�W�����q��z��?~��~x�Y����� oC�� �0<��'��}}n��p2)�UEsPo033�K#�3ҁĨs�&[?!�5����R~N�(q;C���ϻ�byC�Ԟ!SC��(�a���P*O������\���+����޽;ws�ʚ׎�͇���b�38g=>=���%ACԼ�y������Ɉn����L�0��O���N$|���d;O�Y��q5'hT�wCX|�!�p���VJ�j.�``�J*��f��3.��J���%xy�N�z�q>d��V~a�bu�ߺ���V��;N�Y<qY8o�t�P���&=�P�%{N����v�Y�;<���:|M`o���C��t�e|-�j�l<]�������l
���|}��:@�Y4����!��{�t��UC�>�C�5�^��s!���VO�^&��+�vɞ������K���$ԕf#�����{W2\����`Wf��6w��H��j��c��]{�l4�.@2y�
�@��l�nު���fr�;]뵔˧Y�4��56zw��;W5�"����qw%�j�ϹǨK�gq�O�����v��",Lì&�M�	<�&����X�tS���?w����6���5S2���Ԃ���bT���풤���=N$�~q����5R�{��;C�jϾ���q �y��C������ ��Ԙ���<�7W�?zo{�g�]y��t��J��w�HVOӞ�:I*ua�9���r�C�<g�8y@�I����!�S�<C�C�����z�L��������=�S�v�m^�b��a�bA~>��)�>B���	^2z��SS�}���d�����z��:J���b��:qI��>a��:C�*OS�����2Vo)�<I����z����3��&���.sq�ԝ!_̟O�sΎ��*I^�s�����������k�bN���C��$����T��0߰�<C�*�Î��=C9��Ԟ�X~axy������}ͷ���cQ�\��mG����kU�$�>�ϓP�����<�� z�_w�tC��!Y�������1R������_����R����쁩�<�z�&$��5��y�4f�ssѸ�g&9�n�,���� �gHq��O�a;N�
3�b�����1��Agϩ3���)�;B�S����qԬ�g���Rz��y���+�<2�&!��>'���H��f��MUu=<z�����Z��k��T�`}j�g��w�́�����P��t�Y�6�=$�?&09�����N�=�5��&!��w�{ bVN�{�gL��& z�����̃x�b�m�6�YP�Q�:߾xy��~����zN&m�B��8�N���@Y�J��3��?2v�;dRz�~a�S���Y�Nm��N�SR�<��N��c�j�Rb�7����� ᙢ�a�)�ۥ�q�W������~��HbJ��q����3�J���+��RT*�W=C��ԕ�r���>I_���j�P���ԅI����z��38�3��#ͣ��j�X�Ȕ�
����?y�~��T�:~�� �׼�~LN$��d�=C�c'��:H?���7�hx��$��;gHbjã�}aP_��u�:@�*Nн~æ�j�Y�|��}��3������]��..B����S��ջ��Ma��V���/r�,��S-���5�di�L�4�`�u��O{a�#n�߯$���V��x�W�L�4���,*,t�����aw9�6�e�μ�wι���{��XU}@�>>���+�����z�C����1�X��P�}��|�)
�3��ϐ���s^��?0���;O����a��O�S:,�d�*LC�;z����L���9��U*Kd�?7�j����ol8��V�3��& u/�VJʬ�%߾�t�I>B�'~�{'Hq%gL���j(5���0��1=d�ǽ�v��+�8w��l
��W
�]Y�Ό-��8���@�77��>x�l,śCt�K� ^�t[�����~�3~r�o�&�^�~�j�{�=��V�P;7�/���R����V������)k������[	W*���9՝�0���
���Ns�CHg���d���xT��^�����}��Pmr�6{�ۆ�q�^���Kʬl�7F;�B~3�
��h��o��duL�/���y���Om���?�:�Yx:����O��8�^�R��%)�#x�|7���D̚�L����#fԆL��,9��6cB�'&��/��c��π�HS�:UbԏC��7<�F{=��/�ze���к��^�"Cg�eN�6�RpűJ �C\U\m���c��*2�PMH��$؀ ���'t����6sKf�,6="�%���G[���ǷMrtq�eu�i�f��(���M[[�j�v��#ܗ� U���R�r�w������>�6���Xl-x�U�O������溏<lKX�93�uy���:�S��c�Xz����JgQ�̾�?$�;wo��Һ_HF�Ԡ��ӵ�$5>��X���,}��ќ�0���^?��Ӣx�� =���}w6K=IN]��^�v���;R��w���Z;��$c�OBD����B�vtc۠�$BRBK�[.kKܩ��]���q�||Ҭ����[��/݆��s�5���kTz�?\*vyn��T5��^	�W�=0:�c�6��6��<�O���sS ?�+�vL�Ϯ����{��ӹuu#��Y�|M@��r�9�w����`W ��Ȩ����q�KQ5�'�vY�n���1����,��Y���}��-�����U���T���g�J�Ol��Z'�
�E^���k�P��S���S��,~��9T�/)�&1�����k=���W��K�3��h��#!Dŝ$=҃��0��&�B_(��C���d���2��Uwx���Uϻl��t��Y�K�Ob�o��> �:��7
�Mݛ&����}�P��췛/�Ֆ�Z�*ҳݗ6h��F��uZx~����О;~��c��W%�ӴG��������S���rLs�Z�R�O��Z���ԅg�ӣֈ �{-��u�\��Xiםt��f���#o�+�>'��р���ƶ;A��1޻j�[K�Y$�F�%Ej�\Y���+�{Ko����ڗe�f��.P#��XyWƼ&�fI�`�YPpʼ�q���� �)��\Q�zE=޵璤r���q��^�S�(wE�Əo-gjr����}�t|vW����_b���y<;���XMXb��$N��jzâZ����ܸ�"$�p�*�([>yk�M7@�-���m�HP��v��g�o�ݔ�S�X q��³�V�~�:g��z[g�A5��e��H�-�Z=���������j����f��YR����Ӿ�[�D\�'Kۙ�7��>�yh�~�"ư}2!(F[i����ͧ�/��
������Ƞt���t�_�~�����*��'t�ѐ�xq!}�cǄ��R�*�U�kH9f7˽ǖz
Y�w���Q>���k�ѵ���<�]�ʯz���� �i�6��n^�5{�Y^8�e��#L����.���a�=��O���j�O��mEL�KۂB\C�8Fl�w��Y]wb�t��+����P�c���L��:}�8��6-m���^`>�CdK�\�^��X�m�`Wis�]<Mo��!���dq�Rz@��Ȳ.{��U�FWo��.����ف�'�r���^`��"|�1DgX��c+� WBhN�<sx��ەwR��a�.��ҵ��J�
��nH��ܚ��'�8�_����-P&�)�uVF�7��L�ٲL8���rқ�]Z�f�}j���g,5\<ת
]�Ͳ��Y�����M��X�	�Nᐆט�y]p��@8�>u�^a�[�qZ��X^0����0�w��B�v��@>���c�Q�dS�Քo}�n1^ \!�=�/��eE���1تY��Y�hx�H�R1gT{ �e	DK6� ����P�j�6lS3��n���R>���cj������2����z���U3��O޼�B�Wo���.�^�g���܂��W�=�����c������/�"����O��V�+ُ��]��mp�yf��ѹC��lF-~��3�|g����ʾ����_[�,J���'��q��tRc-�fm��� �,�;���+�x��xo(�p�U}�-GMV��N��}H��Vg]Kݟkk�]{k"*��K��n^[�<mBv�4X�<���^4�
�|O�B|kW��C@�Je�N�v��}#���J��<����~�(s�=�	VxW�ʿR��|�Z�7��;�$������:8j�Y�N8)�'�=U]t�{��5�I��B�RqB;��NybA9g7�7;y4�m{ut`z��-�*�uZT���-=OK�P�f���S�53[�&��ލC'm��RV��AxB��p^̾N�Ys 'M�����`��i����ﾾ�ׇ���Պ݊���	���{��|��5���;�:�ȽU2���4�N��wN�t֯-���CÕ�����/��횱]�D��G����eWr/
��u�vo?r�(W|�� z�����*��!N^��\-ѯ
�[i����[�y�k�{ݪ\���{��\χ�ԫ���t��P�[�t��S��]i�^X�A�j�pι||��d�wt�j�xXg���	�0��ܼ�K����I��,n�W]e�"̤���;9 Nh��ny=*�>�*�]��	�s�� 2	;���j$JVc�=�x��I��ڲ�-_g�G��e�m��(��]m�a��'U���/:��J� J��>2�#b�z����5b�%f*��I@�	$�2��:cVCwcE+���*�̫�3�V���b^�T/Wo��[^����uδ����%}u�]�]̊εPE��|.�-S�}*���3��/�WxF�a�)�a>l������T���\~�Y�^Ucg���+ /�w]�2���h��kJ�n��tMIv�u�ݫ������;��/nH���s��5�v�t$���\o��.�U��L�oE�ܾ�m8���4���D!�@w�]�������y=K��V����XhP&��}.�x2]��YV*R�/�`&���p;�miƍ`�a\�o{�M�[Y�Κ^]�m��6�h��`_��~�)H�v/O�w7J蛜3[�P1f��٩�]<%��!�%g&�o˯�>��l���s"���zj�@=��8�J>�JgG�sM�H�U^��v��=�,f��z@��xe�UܸV�~�m��/P�E�祥�&�ї���5����N�5c&��ӒZP�;Y��qՙ����z5[��9eX�xR�{��~�Vw�9�
�$��X���|r/q�x��F�ù�����^o��i�<���{�v��U�y�K�eGm�H���ӞB�{s���*��T�Yjw�֍���pP9;�UL��;2D-|b�\�Ǵ):���k�+�L�ߩOu�zVNkm�CC�`z
��c��c� 5�� �u� �}�_����ˬ����=�gs�o��=��c�@Q��+�g��U��1 )n �ޏȥ�x}�]v'��&x�<�HyxP�h>�|���Z�S���J/�<<��ʴ��ޤ|_ݭ�z�����W~����q��w�w�L�K��Ø|Π!c5�"�F�rR�LC��g�1�?x�%LtS#m=�niCgy�udZ+k�f�{2?-W���N��3/Z�	l�<Y�|*�J7�n�鸥�*�l�il�kv؛���Vd���bB�~�����j"����f
/�t�|*��jƂ5=Ѱ^_@ƫ�L�1�fy��S�?y\��GZy��#�:�|���{�ܺ�Z%��J����+.��xQx��� ���j�"����W�W��;��p��ε�G�޷b{��'�C���t|��Q�A�����:�_3�*&��=vQ2�������yb�&��?�5)8w),uO���<?K7 {�����يti|��6)�i@�i���v�t����>�%�Wpt���РsI��n-6([�/*����J�l��R�a}z��!/�xVa�y�(���5�
�TNe�jխt�-[:��ad�Ƽ逾�}�Y�xm�Z=*�}�����{�p�{��q�@crz��\	]�ے��q��X���{X��XU0Ʒ�J��i�㽫��|Ϲ��[������El�
^iR����c��(2�>bS��F4M}�	�ڭ�Qxv���޲�E
&ksv��D��gQ���p(@Q��?]xP�LX�{�L^/\���t�<�٠Y�|@r�n��WA]v&g�$��SVz�Ż�F�U����ro]"�aa��W7�}��݇�z ��u�DcӢ�X#�[{���ذ^WJY����^%�k�7d�V��K�� �`��C��Y�,�ՙD �?UU}����ˤ��d��˿3'��U���f)��n�4�r)�PS�-���[[]}\]'c�C������c�ڭ�zB�*�\�����5�o�TK߀��k;���\"y* 	�w��[ ����Vu-�/  2
�Se��
�(ӟJ*�]�^���j��P������Vޏm�Gd�u��k�s+f�\��Hc�L]�*�S-aQ�no�E!��Q�x'D{P����:r����아q�_wJ��~�KA���(SIZ�Y����]g,:�\<�5�0��'�����V�f
	;�"֝%K'p�F�G��(Ì�e��硯0�����Ԏ+�ܭ�$!oxnn�zM%C������*��|��-�U�u������f|��T
�<N^�yׯ����{*z�m��U8��{����C���\<5�"�CX�-�"��Mx�:��B֔� �s(Աc�/ #��>���J�C<5�W{-��w^��U�V�k"���i�����5g�\j�w��^�`�@-�_:���2�/i�ԅc�������e}�{��� >͹�
��(�v�|���D�&to:v)�j�Y�ȏ���鞠�Z��W�Eв���W�Ȃ/e�r:0�Rv��Đ+��C��fSv�ʼ��!;����G��0������%V�I�5��SA6F�����T�8>3A�²\��%�xX�赥P��j�|�{	�;�j�ի`;����5xrSq�j�޼�!�-�YqQ��y�����`<I�4��(s&D��!?G`��[�6��5��º"�їH�k�.���0;y�ќ9�6UnMv�Z��!ܨ ک��t�77r]���3+^��7�Dm9�z��-E_w��1��[\�����MX�⎞9$�w�n�3z������S�X��ûBr�5c��"1�5��������U�Y|���)̑�[�W�ºhI5x����:��܈�ot�V-�cq˗"K�Q;������{����|�)��s��|�W����~�^}�"�
��r 9�GX�١���1��]�k��Wj;`N�x�;�U�)IԞ
����e�K+��EP��vV L�bؚ+^Á�̧KHB_��J�k�ۢ�v�EbJ�ե:��5��
^W��2��+��^5�{�(�W�]�س���nZ9�2�V���[�S�h�wd�f<���W(�-\VBDu�����O(ݗ����ے������������X�'��ǐU�M�dT$���f�Zf�T18�.�v:���󍯕�����2�I�����¨�>�и�\�s���4=�Ŋ��v�oeC�4o���̣J��7y�����>	�]Y��t%�x&�r*��Y@ڲM����"��}X�J4m�i٪o�	'��cދ��L�4��51y�	�������ӫ���,�D� �?}��3�<��NҶE����s(��9v����ل/fr	iÞ��j<M* �ei7T[z�g&��
�y ���f/��� �΍�ʙEB]��iwv��rWN�#�%��������E���K��G��uO�q��
�y6�'6�RK���r�.�f���J�,�[t��Gݜ�Fn���u����%4˺�N�`�\#�j4
�J���5ǜz
sg�����͝�!����%T��\&���tuَ��]��gL�y�k�9���A^р�s3$P6��о�A�����p��F��;���:fs@鋳FpjR�#����ak,�C�,���������ם�����"�Xx�h�A��/�<� uo����v����{������N�#�=��/cч�ܖ�<�7�3QP�t)S�V/q�[�b-g>���=�ٕ�Д�	�x5v�ٗfڊ������La��[��=��X+�b��'1L�S���bz�|\2��R�k�*�l����kL����܅M�v�5&b��;���JhwZ�2�Y���ޞ���X�4,B����b�dUPD�%��UX �,����XV�n�*1�B�Pb1TKm�
�nVҵ,DE �@��PQ�XcP�ETYm����+U"�jPL��,P�("+h��F-S�h�I�m��"��YQT���¢��A"�@R"Ĉ��j�)AQJ�J�aYR)"���h(�+U�ʥQ"	QZ��B(�\���Kj1"��*��E�KJ:�U�"*9HҋH��D�V[E%J�����R�E��� �"*".5"�EE�b�Ь6�����eZ��QJ�e+��
�X
��P�TB�QV���� �� �QTU��2�K��F �ɻ�+TH"
�E���w%dUX�QA`�m����UEYYdQjTjR�U��b� �ȣb��V�LITI��Z"�@iIPQE"����U"�����J�aX�b!m
�9�:���vs��������3�!���� ي��[�}�X�^+g芴�"����@��Z��ۥ��AQ'�m�_�}_UW��ãy��,���v3�����|>�V��#�D�טS@?����%U�\D�o�ǝ7�뱒2�F����HlxbINik�
D�<,�uVN���ʫ�|�T���������su6��<4�yד���0�V�PT�Z:Vs���Ṟ|0u/G^-g�B@�O��q����Ѣ�x!�����&�um�~��u��W����(�5g$e��('�@)vq��@T#�,]佛���X��z6)��b���{�K��ӫ)�������*�@�!�8��ڤ�ʺxx�CK�����=�I�-?z} \���ʦdC�����a7(���I݂�-�F���U[���O���m/i��xVKl��4����r��lׅxi�|�#"�/�\���L�΂O��.L]v�]��e>�2���{T)���^�|�EXxW���6���|�+!֕�W5�rL�=��@@V�sfBsB@wP�@G/�&3ڒ��oXo���k2�]���<����EZ���G�+R>.����J!^m5%}f<y8⨖���^���5�2V�;K�h�V9��W])T�L�^(���E��d0;�j%І'W�30d���u�1Y�"g>զ�����k�Y�w�.�GS/�qeF��%v<�t��Hn�(c�P��b��ܠ�\�i���F�����!��0F�},f=��{�o33V��k(�Z�w�����-xX�b��ex��\.��Z\)���XCE��jn%�3�fy���<�D��h>qp�V�}�jf_!�SO�U:���B}��|�z8�<x��{������]�+x����^���y�>Yj�u|���cC�+_ 5oS��v��0jUFƫI��E��)���䝍�އ�1=�{M�PV��tt��!	��q��A\��h�緛�� �m��c��*�d�����>�����e/O�};��ˏ��@�+��?wt��צ�h��`�7�p��ra��[Ʋ���;���g���u�s�����5�b�d�|�ڣx��*���H��Y�L�<����;j�fl�ٮf}ܸS��|%���s��\{<�_���b��@�=G���[�������[�=�E!��y��Oo�_1򾩘L�ǁɻ��<���9�̎�h~�tuX��qu�Ϯs��iu�&�=�����B�J�{��u�Z�-�$�(ixE�QN[q����A�e�)���!k�ԫ<=��w}!�M�93u!㏎�^iC�)P�n}��1�C!�Onm�솒ǆj��L�$�+;e3%��¦a�/p��Y9�o�������P^��Xg@���ĒPvڔ��[�3i`{� ˵�q}��ォXF�^j{)����h������)�������������ĵ���L�f|{��<0���=҈�r�{��(��#
�(Q�t&�C֏�<�;Q��_l��bw�
�R�^m=2�/
.� 5��W��m�g���q�E�9X����P��lb�ó\�����WP�}z��[*=�>E������duLΪ�Z�˵N�j���6<!>�Nێ����!n}�Q��[�[;q*��w��H��sO���|�b�y�o�_U�&�Xl�}8�e���#p�d�#r�.�F[��=r�Nq��{m?|��p���s��>�Uw�:|�+̬��#��m���>��H�i?=��:�]+�Vx�:��S}�K=(T���y�B�iy��rT�K:i�/1�w$�ו���C�L�Ȥ�AD�k=�G5b�[O�R*=�Cr�V`�[F�W�w�9]Q�hr���B��Dzq�c�{1�rNژZ��o�޹�[-����Z�M��ާɋ�S1IH�4������}G�ʯ˳�&�Z�Rt�m�Nn��2Ro��Yٽ3�����r��vgg�n�<״���7s<��9���Ƀa�}��Xt��r����
��v�ku�D�hnfo3y��/�8�Ω��}�δq���ex�;;o��l�]���6)Tm���b~�;#������Vul����Jq��N�u��G*kIڽ���ښ۽l1;��nܵ*v�	`���F���E|�7~Ym|L���"�q����eX�k2v��M(��t��l��{��ƽ��h��?f�����]0{��S��m2T/u���a��Ѡ���f�8׃~��y���U�$��^~�2�����R-E�/!T�X�=J��-&�ZY�v
�2�T���<��f��f�?{O�b���Ha5�g���֥}�R�m�|�{W��P�<�����l_��L��h9��7~w���ac�������lu)Ye��'kf�;V�*)?l���ޮq(��ޜ�T��ۧ��<2OJ[L��2�kd�J��kl2>�1Fϫ���0�ٳ��
i�	��աK7܇0/Z�h7��3
��Ģ�ZTn	�[���:5
�X�St��^�D�r q���L��h�_s0/��
�U��Ϋf>ɴ���F��c������H��������+���G9�=R�;��f�y�V*��j�,b�lM����F�V ��=�UN\��d���hck]�/��������W�zG�R��S�S���N~>�f���%E���=Z�!�~W�����Σ�G��^t��;�T��T�_w�B��s8������\��3K�>#ܹ�v���O*��m��}:�ͧۄq��)b��FVH7�:�������·J�ǯG����4�4�O
Ժep�Ns�ϷkO��7+��Gڷ̟2<�Nܤϰgu��3:�;�����XȦ�P�dVF����1	����r��]K%��~Gbu�`-m���]�yw�w��R�;}2�]�l�Ņ���}�gR߽��W���y��^T��+�����(�׾��ל���7�(M��T��_���b��o	�`;�KM׫��v�wj��Z�}�O׽UW��m��}?�����3kث���œk�ڽ��:�ǲ����M3�����G�WG���̼��@hufps�����[��xzu�(���o]fJ���HX1���s�=η��X�&�^0�N�[��r���:�3F�_m�@�)I]c�W���u��_�"��꯫�B���,�\��T���\pV}�]6�s���Y��=�]_�L��L�&�M�[�]�̯ �^!���K<l���Sʿc����l'KU۷�͓��mh�j�J���k��C�&�c�Ci�[�|e��im�PY�1X�V�r�N��*����S�(m2쾓���$��l�g��ں������J�-���z��X��P�u��PIt�H��U�7L�`���j{���v�r�?,/�8���>��άk�ո|smg�ל}�9��݊ko�"�:�����X�MCh}��(��R����h��Z�}	ŃƟs�Ӡ��W�OX��?qK���_3C�\5^�8{o>�}�ڔ~�������oν8fN����y�U���O����+�=9_�f�h��y�����5��{g>�O.Wz�o��S��*˨��_I�٪�N'u��뙗���'X�z�t�<�����y�^�\'��Q�UP1�׶ vo%�wt�e(
�l���<�g{`�M�X����
�\U֙�z�$J��6pQ���Q�;��+h�Zww�5���[ʷR��rp2��_�U}_}UXuE+��^,36���ʶ���Gy	)�N�w.g����۔}��\�s��Xq�{꾮{�f�5���n{�oiOy�>c������y��GԽ��\�"����f��m�Tw��>�[��<����̅���Z�6h҄�_���k������T�T}픻b	�SO�;�WCej��W��%iC�eB�ulzT�l�e��.dU�;C���>=ه�t)���R���!��0��6�Q��Sx��L�6j�V���o������O4����˶8�Fq6(�L�v��!�����x6A�)�Ռ|������|�.�Z��ƿ����f\�Mon���0��U@k)�@�B�ងf��&��zE�� �`wWA�Ju9��M��s���ų�}�l���V�;�h�@TPR�E��˴l�S��X4Y��l��hx�'��%��R��K���qɗs��|@�X�@%7�^���howpt�|3oR�56LR��Β�kn���΢�4�N���b"fK��k(���a�ӂ��
YeG�о�Q�`;����V�͊}�V,�������܋�YQ�h��1mz7�N�jG~�+h��_CA��k��Ȝ�vD�	������[�N��jv�~���M8ꗐ{�V��x����a��NR~̣�8x���We!㫨S�ñ�t����R؁a9�4%��y���RVw�%l�ݡ�ߧO����|�ܓ�\7%p]�^O|����A��Kz�[ȫ&�\8�W�����t������oPd҂d<�Ɩ-���:򽚶(�yl��I���ʖY)?t����K�Kv<��a�v�v�k�^Q���T����H��-��Zi����wO$�.�ΔGwa]�Mw���
�m>+�͵�I��
6<����ۻ����.g�޿�;{~�5�U�2缾�λ�Y�X���T���OPƭ��ש��kܯ�Ѕ�޺�ym,���M[��U��v�Ꮋ�]A4�j���݁ԏ;_����}ȗ��*�߱L=x��2��D��J>彚�f���w_�Ѷ�yЋ��ui��*(���(4PI��1e�r��#�C2�斜eb9�j���-�Ĭې%�x4�2���]X��׶��u����ﾪ䧩����뒺�Q���~em,�<�m�d��o���32��F�-�\�����5����B�,��e��^��Ψ��*\���sNqT8w����Cg�ҧt;ؕV�t���-�M3�,���ڥ���7,���hj�Dk�_j^`���z��hؽLi��U$��m�j�&DK��#��J�)}������tV���z�6�Ca�h�AB���0�I���W��v�dG��\^�?y!��#�iu/>�S:���������û����=���}�2��6��6�� J�������^�.���O�N�=�k}apա��zc)���\C��2<�ÝG(�my�T�|M[+Ìo�em��Iy�p�{�؆i[jYn�6ڳ����I!��ci��sE��auI�� ژ���l��𝯷+��ѭ���Ë����t9�:W3U��%E=J�(�Nv��ꇈ���u��ٻb�r�c)k�#6�kP�]6|�M�0>6��`����3\�����MKW�XUJ
͠�2�X�:`ԕ�KO3�IT���O��]��i}31Mvu���`��Ϋy�/R���8?M��ƗA� �����>����3y��1S�i��;|�r᤭Sq�{�Z��7�)J;�M���N"�^�������hࠛ[�����}N7�>k�����v��딺Iۭ%;���Ӌ��S��J�>�:��t��_�u<�(����X��<�G�s�sͤ������݀�>�X��k:>��o���W��Za�%3��2sUa��P��f�ؕ!ۢ�O�u{��R�γ%��l.��Z�N1SI��kkw2XFؔ��j�16_�K����[!�\�s.��e�/ۭ�{x^���K�v��b���{L3�l�a�c�FH P�a�n���(I�՞O�,b�aw���A~��~Ҕ�њN�n1���ɴ�d|�N�^�1{ۣ�S��f�cn�a�Ө{q�?.<�j����:'����<��;9 ����/��4�-�]�R��>��[�/���a�¨��hfnk��A�
����x���Ա�&��}b�A[��X������]����t�lj�p��Pt[r�'����+dk&N���f� ����yR��5D�'��i��<��|�h\V�ps׽t���*��r����"�޼���S�6�y]FX�w��6��R�v.r���ӭ�;+D�`R�.f�������VӢ����nWv�
U�ℋ�#��yr�ȑd��n]��&�fp�DT�&>T�!��=�ds��t83ͱ��}m����Ch�����=��i2�S(5�������? �#����V�����AR��z�����Ջ�p�p[1�]�:b�<��wfP"ybW���+�i��zd�YCE�P���le��@ܸ�m��zcy��x��s����t��t/a�b�1j��
u�#	��e���y 9��DfWT����� !�a���=.A���Ҹw-��b�a�n���uy;{���_Y��C�=�j �6�ۘTTAnE�tE�3F+�P���F$��k�J�K���۲2��<��/�*W8�X��]����х]�g)�Ѧ�(�2��ڊ,q�ǵ���\�7Y�5Sl����} p�u��^���mf�����,���]7X���.�{��-
o���UL��f��ʁgϋ��_S��ˤ�w�EV��3�od9l'��;�����\��.��D�*����!ڸ�W_>�C4w��AZ�q����dβ� �V�WŊΗ�25��X{q��v�{`���487� �^nD59���'��{
w.ʕ�WP+�_w���\V��>靍�5��I�E��}R�tj�$�EY:&9(s�n�+�U_.���j�'B�iڳ\rܙh���Ϊ�)��	0��*���uB����й؍��7��Ru�d�j٫������f��8�$=����>�89l�l�';.3���h�m�u�d�^BQ�&l;�`��	�ɽBLޫ�9c���u�(ػ�K
(�"�5c���eT��9�0a5��;��Ɔur6���<J�'�}2����Li�7j�5�藴8ܩ#XJ��#.�3��:81��X��O���.<{Yv��LɗSv=^])��o�=ʁ=�Zk��W%�2;�}>�FQ�qu]�3����z^ܜ)LR{�8C�`Md6�ں;Ҷ�2^ai��fA�$ʔ���]��#��N�WN�u��Z�ӱz8f�/��㬜���V�rA��J'���ۢ�K�&��AOKZ)��	uz�0oH�\ἵꖪ���صKl<;��X!b���[��Z�OXk��tH����ك�������zKY�W=�v�����{���Y-ATQ@U�h�Ym�Ȕ��b�V�������+"�X�ֈ

�C�\chV,"0Y*AV
�� �mB�R-eQ�Z��
,Ęe�d�,�,�""�1U(�3���`QX
,���TQb$QLIF9J��
���"�d+F
 �AB�#X��*cEV"��aR
 ��DJ�DF,-���b�X���E��j �1%E�UB�9`�eE���XV�k
�J�EdP*��FchV�UDX��$QH�²V,Zª��X�*ADJ�X�U����V[d��h�PT�+�aE�Հ�U�UF�QR
Im�"Ŋ#hE��U��1�����UU�
��[P11��EQ �"[m%AEV��H�iH*0Y1Kem��V(ZX��72�b�H���U�Oףws�y�ǽ�:Oʟ�+���V ��s�����{��e*e�!A�J����"�o�;��0�Kѵ�(�[�}���Up�|��O8�/[��{U���v["�|S�������3uu/\𲦌�c����F�ϖV���VS�]ޜ}�f� ������Y����7ԭ72��. ���N�[j�����74�ꭔ�rY��M�W�G%s�.r�>�d��wg[��mz���Q	�x�����^�ث{�1��Cҷ67�_�����Q/���շ�t_�����9J�:�ɼ������9��]ws����r���{���<:����c��%-���J�|r�v��ε��>Hs�q[+��ףy���^�g��@o���*���f���iރO�>�*�MJq��.�s�����^��}�;����+�m\�~���b���\>AyOf[Ɋ�5M������J$��,�-�;�͙��dVR��+�7�W��%F��*e�^L��V��>G��0�u6j�u�yU���Ҩamyq�]�|�)�>�P?�h�owv9ƹ�l�݈^�@���I�m����x����x��1ӻwK&NF��uǩ�43���w%�s6o��&���WǮ��z��E��/u�\b����`Q�f��k�7����h����0��V��N�������-�I��}�8i+5+�}_W�}v�UhԀl�wWQ;%�R������Z=Sξ�W������U�8rS�k�7�.�_�wYT����/5�OƑc)r�o��*e�A~�+�IA&���I���Bd�{]� ��5��V��|�;w�fo����|V,O����Ȼ T����{z@������k�#�-}NRJ��sp�f^Z����yk���	��B�2ef��G�@e�=Qh�ewp�l�6{�WI�n��!�˩v����T����|�}���������k�g��}+����[����.�]K��-��	��k�ˍ{�1�t�^�M��n��:ͯsW�4<���wS�/��������{x�y�b��5���cǍ���<��7���{��I��؝C���L}�Jn�'�����Lܫ��:���d����l�g�g��Jq�z�}x�C=|���\Q�J� c���W].�[0u����޽=k�8����2�^ ^�A�a���
���];��G.ɕ�����#����(�c�/$���$xM�ٜo:�	�\��3�ɰz28�-5zuB:��޸b�~X1��Ȟ�!��	��Ő �S
�e?�}U_}�.~�=��."y�f��g��e��¡(�c��=�W+��ܟE��S�=F��钳���lm{ű��6�==$�\��z�V�{�x(Wv�v^�\�OZ� �z��b����[S9g�my�M������>�|n���X�?Q�.r]an��Jx,�沈�=�k:]�m�j�ɿ_zޔ��:ũ��!/�|�ycSݺ�}�o| �BW���Kuj��)��d7��.;Gut��I�����osE������7��}���K�+�lc��{IAr�d�;��1�sor�U-P.��b�8�Ki�.�:�-�u3�y���E��1���k伈�� �ZȅBv�L2OJ}�bQ%k-���Fi�KZ�HJ�FF�-{�5����auy�mT������^x�~�#f:�_
���ȰǸK9�ݑ�I�^N��1K��+Z�y�X��=�T�s���yW�p<8[+�r�
�US3ߊVf�8�H��N����s���d���/�gASoLSӧ�&΁�ф-�=q��Sܮb[�a�;<i�u\od��ˬخv�^�[�t���kFcs�@,���}��}�{������S��ӕ�GQP�u��~(�]G�1�7ՙw��������	V���=�sƦ�>!lJ�?J���G��k���{����w���K<uI����z��|��N���<�ϩ�	�gm=p{ir��
�=��o׵�3�r��32�\��NnL��WJo�Z�`Wׇ`�$84�k3ɿ������u�FM�Q>�Gw��ؽɏV���a�J|2��c;��Bf4O{�7E�^W�.Q�/Jro��ݏ��n�S\����Z]Y�YS�ƵI��\���۵��^�&Wl�50�w��v�-��<ߊy���Ŀ˧=v}_�M���:}�,�(�m�C�1J�DnUW���+,�����lK/��N���c1�6����?��[,U��[���QHA��Sy�/�H����K�&�}�'�ox���R�J��x�M����O�
ƹ
������ ї6��1���	��m���9C\�pN�+)���a]N�M�k��n��[�ƌ:��1Ә�{���<�g��W5���E -oh�Z�(��κ8�v��n�w,\rݥ'�Z����sZ��BG�>�-K#���I��65����΀��ϫgmb�Zw<��O�[|��f�[�,�[d����H.�u�!K�8�kAݲSb�Lm����Ne��Wm���XjS��dmUg���c)r��ʦ_d��_�WGHEm�ư�ZT���o�"3[u�~Ma^5H�{�󰺘���R��=��ʽ�\95Dm���������C�=��~�h�|���k�V����W�%>�t��&��Q�sO�al���J��k�:���=��)P���l��L���cf�3��{+f�=J��T#����}t}D�6I�K;ܽ��h�Gr=I�a���Zc��a�V�[yj�B���_!�w�q�^�*��
N��uI�^dzq���~��}3���"n?Q>��#�j��!��W��i3���?c�y�T��������zj���-�6�[Ʃ%ZL�n�ܳ>K;E�zc�iݮ��"��[]^�q�H��i��cV�.���c��tc�����������r>�V)�b4㺓C#�Ec�"������h���2�=ӍsT�U�+BS7������<����`R��t����Wy+��}�}��ꍚLo�+��MY��F�E�a��Vjn��*�z�3���.f����s���6�+n�ed�Jf�Z=��Qm�aC;'���v�.�Wj�����x=�y��w��K`*��T��ص���+_�o�Os�ޜ���Y���Y�ȟ��'��Ug���2��W�{կ��*➧6�m'��懙͙^�m\��=��y֝Wr6_��_֟6(���-A���/"׽;]w���p�[T%t߬c�����*���g�U�ڀ��i�|�����sp���[�E(�,�[$����u9O+�>o���k�3w/�-m�Ž�zT\�T�H�v�ABOJ[L�,�K�PU��y�Ar����[��J�Vu���F��>��zM6�jR�xe��[$�IM�j�N�l���2� :l���⑚��ɩz��ԣ�z���[&��{+&�)Q�,���T5~^@�Da����ǧ-��:n�/�Rc�yg���9�U�1]t�odyT���Y|�ν�D'w�Pm�kd�<L���C+hB��x���V��PK�\�U��{��s����H�]m�������n�
2��'aF'��Րz�]�qL���&�vW���v d>��M��3{��'���A��u�x�Q�=�o�/.�Ω�&���<'o��S��Е3��攔c�p�EZ���F����+���r���.7�Ҙ����ۘ��� ��y��ޜ5�9	:\���2�zWNj��z�k��ul���zs�
��r);�����Ϊ�ǽ�{�{�Vo�h\u+���)��gܲ�X�$m)����ej�T���BX$n�m�X�DU�:A�&҈)����&z�'Ş��}OySo���fD�� �Y�wb��ͳPB҆^ל��t5�<�R�=��ͣ����R��ǀ�^�JS9�j�u�毶
�ߐ�̭���L��ʪ���|Nd6n&���F-�[���X`��&SFfJ,�V��j�v��<�oǼپ%����z��6�w9v�R��؆&���g�l���d��Ug�����=���F쇛WW��y^�\o	�V�ӶU[#���Cܑ��u$q�ҭ��uk��� �;��w97J�.��}�x�����=>�e7�������5C�U��q�{���8-�X��\UW�W��|9���a�R�����]�C��6(8�Ki�vmJ��e��՚����t��QQ�cRk�b�{gMmLԖ;��	�:�$��m3������1m �!=�xu,Uu�z�w�;0f� _լZ�(�d<�j	I��L���?ư��&�=�����k��3A����8�Q�}C�X�}J�||s�鋷�tOϬ�^���\�߻��hz���wؽ>E�TǕ)f�s����S�,�e����%;j�Sʳ{R2����N�]T7�P���I�<��=������rzp��<�a~�7γ��p{Z���Y<'�?*]�"n&D��ȓ�Ŏ��<����o����T/��:����n�7��������ig�ex���̎�{ݿ=��趽�;���혧LY��g�S�����uM��g&yƴ��Q����q�Q�w�sI��F���U�B�*]�^�(�6cj\�˨fb=}Ϩ�cvI��Ūc���M�ZپPӫ�\���������^���F�,�Yw~��(��7v�a��{}�O]��Bk\�˭1��s�׹T�t�X��cG�m�7��Y�}�v_j�Z��oy���Z�n0Ꙇ���q�p�u�E�/`�|�6z>�1�����F������&_�k�����d]F����h��f�ٷ5PR��a����1�ާ��q�S������5�ʅ�n��iR�gK:�[aB�Ϫy)=4�����)ە{�u\�Uک�O�pbui�M���>�-v@����G�x`F׸^��\έ��m{%̪�A{�W#e�ƽ���M�be�ڳIrѪ�q�]]C��Ns�#�VJ}V�{~��}}`�z�X�A�_z��"���E)�̤hf]R�g;���e���F=�ݷ%�Z�iO�z�X/�ֲ�)�6�>D�Y^O�\���7��'��A�G���|�-]�9/���Mǂg�4guvZ���wX֥b�W
^�%�,DH�ϵ���yޔ�^Ϋ� ���֏��{i�X��g�w�w��^!��V١�[��7;/�(�|/�he���EX��u+,�=����w�:�pS�z�~���꽾�Jr�Q��E�V@r�6�>�*���5�|�2f�J�p��u'R���"E�x�t4Ws��U#�_6�\�9�6C�X��{��{�m����n	�����a�����m1��#��S��}���~b.}|
�ה"����o���'��wa���*͡��0ms#ӏ�wo�ۓӦ���w64�����>'��RX�ϯ��γ��psMex򣳙<�S�R�F{g&׫ݼ�zNY�՝��Z���N�:�����W1%/��ZL�=�r�h�"�%�\f]n���\�[{�\�j}P����f���W�kSJ���x+�p���*�MKyRQ7j<U�m��5&��cTB��ۨPԤਖ਼�tu-�%m>��̹�a���Eފ[~`�\n�ؕ!���������U�4+d����!�t�4ъ�Bəa���A����M���kVة-^�����w��hW����>���҆�����:�����$fU�9&�e^�x�lmt�q�ge��Ce����_g��E�\����Uq�������-20�|ג�N����8�?\��a�Q�w/e��0�46��Qj�Yk�s �$��69@V��J�{O��o�c���X2>�B5��8�b�77 ��
�F���Q�e�����ސ�����i�s������B�����y���C����<m��)6�X�C;��5�K��mg4�l�\�_���L{;�"�r�b�
R>���a�L�\^�lm@�i�Zb+�OX����u�50Mɉ)�s�%���C��'R�3@���,�Γ�Y�v9��Vj)K��Z�͵@�O�%�0o�m���un��鬣:��n=Z�Ek�����-\��׸w{C&z��6"3��w,h�9E��`�R�V�x��^�S�eE^��r��4�K�9<�S�����||�7����˭7i	���\���W�[F�J�VAչ��d�t@�u*ʕ����2�[\��_A�o(R���+={�sN:S-f�1�+����p��rXK9���n�Z}�t;5�*�2%�cm֕]�n"
���u)L��ޑܭӄT�r�W ���YzG>�7���U,�κ�ń񝬇�r����m�v��}��^ؔ�|����T�m+����u�um�z�e���)i4+�{.��la��}�'�0&��l�=�t���,б����P�k�����f��� }2I+�2�P�֥(� �w�u���t���?eH�JK��Y+e���2��\B����]�D4k3
ߴ����~MUJ\3F�;Ǻ�[��U*;���{c��ȷ6���Y�)ѧ��Vo�]1�)[
��V�_L�4%�+7����&Ι�:�9u�L-����s%vw �z���eu[�hp�}��\�H�2ēTC��b!��Ѩ�T�2�3'�����D����n�],uo���G"�W�������b��0N�)s��	�w i0�p g8��p�J�X똦�\�ދ�0�I��OokktWB�S�/L7Zx����������̜۾{�V��SO.Ĺ\�I�(*���]a��:-w�q��* �D���\�Z�ʻ�on�-"��̴���ӌ	&1-�iA��\l��wl��T�x�u��h��%��D$��g�9�S����B.�4S'@��������]��
�Ԫ.̻�_
�S�.��V�"�����E'9`G�'q�H�N��W\�^�t]b����J���;Ȫ����@V9B��K!'�K�3�<��=y�Z��k�Yxk��-�c�k�v�U����p����l�b���j�`�/��ɶ��M^��Z�j�r5�o`����Z_x�{�1X��sz�e��`WH�b����.�Wѡ�Y������Է��G�!��oZ�t�C�Wy��^YCgG�7b1�j�⶷ӄK³[!Ю����6��W��&�E��b
KS1_[}s�WSCq`�m�ĺ���K��@��sQ[$�<2r�\�C�ϯw�<���e�v��ᗇg����v�(��%VVdP�m�UEUAE��إEQ��Q�h�V6�DF1�X(��
��e���ȰX,X��+E��)*�Vj ��**(
T��b�E�EP��RV&5L��IR�%J������lFDb+Z�Pm�B(*�eIF)R���KB�X,EHT�(����"�T#i%)P)��,������J%��R�")Y+ ��DQ�l�(���T��F
A��$�#l�R,X)R��+��2"*��\d�E*���eD��cb)Z,X�� ��@�(�+*Ek%`���	Z��#h�T
��*B���eH�T�T!Y*)r¢��T%�������QchT�C�J��J�,Y�U��|�Ǚr� �;�k���V�8�����SX^5Y`5F�����x�L�F��`[�zn��4~�	i���0��
����m���d�MB~DS��f�)F�g��$�-e�%�T��l��U�� ]o%�f����OJ���W���Ѩ-d���zo,�K�ѕZ�8/j����B��\���:��)�~��{�_��qҏa�՚2���U�	���Npl�mh�*�wik�l��^)	�ؼ���jMKi�,�:�=G�ӏ�Y�1��E� |�Φ������4:�����ǵ�!yu1������U�Qc{6.۾=����x��9�ܓ=�䯸�<�Þ�{�*!v����9�#���Jry�W�V�G��=���='8��:��Ǹ���6��2緻(���<�ԅ�%޾��sy�o(k�yW�u����֤ϰwnY�X�Vb�5��L��Ew{ 9^�~�;н�m��f����j�a��-E�h��ɦ
�s�_�l8�>��.��_�ƣ��]mQ>��=�K=�}="��>���|.7|v�P��S�� ��;�nv���w�#zh�l��Gm�et��3�%�2��g�+�謀�E�-3�EBт�u��1���h����^-��\���>L���N����*'<�t�/�F�"I�80��':��S��UUU�n;}���f~�[΅��kۋj�r5�<�"���W1����vE�1�s����i����u�7]����yU{�*�Jm��%��eeHN[�՜ę��y��T�m�N�q�#�\�?-��y�=��Z�Ѽ�׷�wM̥�r��N���lwSl��� k;V�O3j­�]�����c��v��>��0��r4���%��<]�ni�n2=bs�W��?#�a.�UM݇�
�0Q�GRF`�ȵ����q9��CI��:\�5�{��ߎ%�[Z��i��X#Z�PA���*.չx�_"봶��7�.;���eţ��~�#���_�u�WV�Ǖ�i�o����%{L���X����35�Z!=)�|j�\��/��bd{^<0���,��勞L�{��ݥ���J�q�QϨ�tF0��� �Sşo5,�/����}��R���Xj�w�� X6 ����l��vk��˄]`���6�5)�y��2��ei��Ϟ���0u˃���{\x��46<�ۛ�	�W\��3^jsj�F�	��tJ.ܝ
 �x��#H�$>ذ��]���՚��������6����kP훚a��R���^�w�^�:�RHkdV�>QH�ج�F��D��-��i+$n,k;���vś�Q����)d��
,�$j��R�.�2��2���x����o���v��uw���� U��8CM�}�|�{��ƌ�U�I��� ��߉�{����ң4n�Whc�hׅ��jt�)�H���X�r�0��D՞�~>��U/�V����M�v���v���*��pl�R��kڝ>Ϩ��ѵ[�h��kt|B�7i\���{(��j�wz)m�T.7Sl4�']�k-��W<����Tu6=O�d��R����BZ�f�6_ւv�|��Ǎ�m��H���~��<�׆�a���Z�<�2�`�s �5�W,6]� l)w�ء�&G����W���J�J�Ւ�ڱ��Ug��7[@�j�7 U����
��!�	ѧ�Ypeqe����M��`��qel8`58�B.tV@&Ɲ�B����B��=6�$+�1谺�&3K��K���㗊��n����%��o8�7;�|o7�$A"�jh���y����9T�5��!�3�N���{��,�yY�j6魁�9�����1ɻl궧�SS��j�ź��g/ 1���*��&�$�+i$e�تVI6�Sem?"��Z�U��Ҍf�9������w�v�cN�%m>>���{j������A��[��`��ɌeH�7��>�e/)QZԡ��S��Y�emժr6����ېl��'Sy�X��.W�o+��r�k���uNߘ��~�S����ysK�4nv����j�{���毼~J��ݡ�H��Lwm?nE�݊
׳o�'#���%��c�k�ޗ�U�D=��5��ʶ���t���u]y��n�y��y�I�;�5��}ٳ� �ZL�n���j���Lb:��ԋ��P�1e����x�v�VTN��O���l,e��"�e[��1m��^��
M �&Sva�nG�n�
��͵��oУLw��O��t��{H�c�ǔ��YE�sY��Mz�Ȕ{��n�<U�\@�.9�������V!:�2E����_c7��Ҟٰ4Q= �����3�E�����'bW2�b�۱g���t�� ��`�	���3�zN;����y��^����u (c�3(z��Rβ^�S�]襶ͅX�e���3�r۹;*�����W0嗓�V�lW.�P�K,���V��>@դ����l9پ�z4��q�Z{G��L��=���Oii�1Q�6~�92�d�]�i�zx���d�jM�,�Sel��Z[cz�y?E�\���V�uv���LO�ƕ��!k:��Q��+L����k���h�2W�A/F�=+��|{ ������u��
�y�2���l�%�z��{��>,l�i��wA�8&��vDւ��6�P����}Z�_����=�Դ;�ՔR�ֽ|}ذ���y[=�:=��[�˩{~}K'P���mwy��R�M�|b���R�ݓK�S�=�wy܈�|�QT����U�����4���OyX�.)���9=�\=�J���5�o�v;����QN�`�c��箵X#rN�P[�g�ݶo&l���ڿ8p��e��=�[<�$֑��Mn�`��ޞ�d<��4C"�~���¥7���W�Sk9�g���Kyr���jY��咁Z�� f*K�!aQS��>���Q��6��u��Q-�Wy����5�f��v1|͹���nk�m����gmP���R���+�I(r��ui��=8~�ޕX��g9��J���f��s>�gh�fE���/_..v���,��^��f���m�{�S�6���5Q�=������y[ޖ���rT�s�46��^��ߞr����tI��zL���������7+w��ڽ���4׺ӷ��X9ٯs�X��#0���c���ԥ�i8�Om���L�~蝍a��kn�J��'Ȳ֡�Wꆨ���t&����!�yZt��lq�S�u:\�b>���\�]�����\U;O!�1��cKY�c���Ը��\�Jjm�l����6(8�5C>�-�q�C��R��| !��=��/�<U^^��{U�6�K�V�*=�-��e�������{���<-@+'�^����4�m���#a��:�$��i�w"��fD��msGe����j�]�7񃓜��aC�k��S���ٔh,�֬�ź�:ý�l�[}]��v!���+pk��[5�����������츱]�m����<�Aj��g�%�zĬR��v�vm��Wfa+�0�{��������������.@{����,�n�6��涠�z���c�t�5_Sc��h1��^w�/?{��^�_IsO�cͪ���@Hײ�o�<��,/�PխJ��E���T^k��6�2���W��^�f�/ v���?QP�Q��~(�H�Zr�nž�Y��1L�S��!27P̯+=�T���C��T�L�|�z+�:�/g�v�=��j9�;Y�t{æ�T�9o�ەS���/�}��������Iw�p%Y���W/�'����c�_n}�tu��a/��]i�Y%O�w�䕇��/}~�N�J���[D�ڢ;�i�v��iw�~��r5a�K���;m/t�YJ�#S�M�U[V��x-m���b�NM�u;��ɠu�v�Do<����S7�#myjŕj�:Q��>�7�d��ŝȡ;��"���Je�I�Q��	b�,�	��;w�d�+�(�ѩ�5�uf��[W�B������k���-�.��ȹ�������m�j�^�Uѡ-4�볝+*��|��z(kC��s���7 ��%��Ԫ��WJ���t�b�r��f�og�K�2�v�0���{ݤ���<2P	+�pg/���0�R��f�Z��Ekۯ=�����Z�w{��T.wS)f�3�:Yٓ�{�²��[k�[�t�c���W��i�fF�T��kA;{)�<5i�8�5C&�/�;��v0B䗳����ў���j�' *�:����V���f���]���Y�j�]���ֵ=;]Ey^��� J�������~(��X=�S/�>��ůyľ^bR���aK�#e���t�&�/}s�y�Q�v�SO�BҮ��U�e��ʆvL�&6�F ��>�b���M�1��r��ǥ��F�,��x����OoK��%�b�c�Z���zT+�}S`T�QVtQ{l�oU��a�J~��ݾ�1�5(����c����e^U��T��{�ô鍚���<�og���s�p���B����~�:pڬ�.�,:RM�z-���?x��g�_���5C��izR��t.��>ޘ{�y���	����k��t�
n`���^��{��i��Y�H��;�N1���`�C��m����{2�YF�uN/��ɑ�~��wc%b���u�g\۾�4'?/nƐ>���a������
b�ՄN�'�j���U_r�$�%/� ���%��+n��md��}���j����[�����@�n裪'1.�v6!�i2���W0�n=��2NܲL��s?d4�m�x��{�����O7�k��v�zcv3s!�V\�&���J}�����YY����xS�3z���14T�d�V�2��6�c���U\���h�p��u���l���D�ɚ�Z�=Xש]	q�U�š�·.������m�W�{���u.�]��,�f]z�B�Wu]R�.���Y3>/j�1˃Ѝn4�KѾ�����!�=��߽,v粴J����vK��m���g��'s��X�ؠ�eF�l��q�C���'�T��;X�/{7��яwz>�i#��YI�ͽ�]��3�>���3�^��x� ,ר4M�6�ӕ�B��ҝ����ԓ�B�5�PZ�=)m3^� ������/C�v��4f�������1)���jp�OoK=����q�=���{�к�\�i>�[-��;{�m�����:���w&��G��^c��Nڂ��F��LE��Y�x1_)8���\W�Pn�`���M�m\yBh
fNfU�U���Yz��8�������i�Z��)+0׬[(l���״�Z���(�ݛ�ђ�AJdF�+b���*�iTx퉉Qjj^��Z����N�=��ġK4�w���ޕ��׳�v��ː}�ڿV�3�r�kD/.�Θ��çxb��Kgbu��Uޖ�z�ږe�Pز�KT�ѩP�y��N�b{|���j�Ҷ,z���KFxF�)��t�0����&�:���p9�]�ݻ88n�hW�$���,�I��-�|G�{ݵO��F��W����w�~����~Y!���T��������[�kN��#����I)��^����{�dc��	Jʥ��l���Z�n����;O9V��{��{g��\�˂utu�:��� �?��!��v��OW���9U�v~
��U���UY�4�ϵ(֌�V[���U*��Vm&Wc'YnJ��e�(f�;K�1�7*���.���cS*+u;����w�_�������	��Bv^XFs�^e'��˹|�������{}�N�Ѻw���G"9ܚغVv �c^���1��5���b�s�m��չ� .Gv�WD?�a[��%M6�����rB�������҆ᾛʭ���ښ�V��=
f2�ësG8��;*���o(�d��H��/t�kc{}t0�icu�0��0����c���$s��L:�8]��bS�L�[��gX�'uY�#��^�'E�]��)�T�fh0��	��Gn�kU|.Ո���ks�&�[/WVfIբ�p#Xp]���o~2N��h�6���,F_�me����9�E��ĳ��WV�U�ct�ʖ������b�]�^c�>u��"�H�:5j�l��|�ne�i"�+r����P��1�Sݾ|'��Yuw�
wrr��Z����p�� �l��0w�VT���II^^\뿆":�[�dc �C��}�W8�$�vmHLG1��Gp������G����y���K�0�ޱe��*,��r9Ӈ��M�+L�jĔ���g8�Ǡ�O�R,�����T��E��awg%n��M�˱��"�@�= �C������ϫCy����׵�r����ݸ�a:BX���vo�o�̪εE
�hY�q*���!ڏ*��q���P=�<o���n��F#n(��So��������u{�����7��s�8������+��/�N��S���Ĩ���U?�[s�t�3r�-�ۨ Rdm��4������#%��:77)̎�*x�kI��te˝*��x�E�'yid����V]f�T�a��:U��v���V�x����+R%;�/���k8:�@趍��գ�h]���G�֎(=�=W�3���dr�:�r�椝�W;���eo!ty�f�]]qH���r>�q�Xc���&���br�ܬ�7��_!��S��Z̭�/��G��^#!�u�^��n�u_͠��|���@f�YBA��F�6�mުO>�*օ�3���2O);�S���_vr3���u9��U�XJ�ò��Ut��X�e*���Y}vD���7����>�tgny��`��Ȝ�Ԗ��y��� ;�/���/�2���{OwR��J�n���x(0��:�#�/9���j^1фܖ�Z����Zu�;1����6�ѿ��vw���sy��#���V���;�ηqs#��}W�b�wB��Y�nQU,D���;�6����N���c�L��Y�Q���.��8+xJW��&�;�n���d�٪NM@��Ց7���WW_^n�	�3��s��+D@���/�[����6Hjȫn�e;&�֬�pV�5Z��H������D}0�5�	�Ax���;��'"|���v'{�6�$1-��៼Ϋߋ�'�
�1*�T��UAVE�I�jTiLf�Ld���m ��B�VUMB�X9J2
����2�����VTX��,��]HV+QTPP
T��f\ea�,EP��HT�5�m	DU\d�7(�d���-1�81`�$�,1��F��v˶�$m$��Ԫ�V,6�Z�[l�*�QB,im`�P��t���,*TF*,�ĨJ�LJ�d��
�6�%aPR���`:�[aP�Z����+
�j-J��E�1�-�"Ԃ���2�f�b]��Y"�aL��[AaX6�$r�& �UB����bZ�La��H�TJ�VJ�H,�R�-J��)��5�6�m!Da���Ad*JR�*�,2�b ,�*������9z�2��*������nVc�4_V.�a_K#a̶��ˈ毮��i��	����#�;b�-�����Y����}U�wz{����?��O��^�lR�3��k-�+ڎ���Ec���9�}��,O��L�.�)|в�S؆&���gh�E�W���ѹ��y���C��>�<�ک�.ԩ=������Sb�%(�mmV�����=a�7_�OjِVJ}�2�4��Qv��_ի�}�'�N�	�5i����[�a�(�/��zw��S�;���~hi�H�]���ǽ���nPQߓ�y	b�zs�����-ȸ�)��M��\W���~�+����������e��/.wÖV׾�ޥ�����ޅf�����c2Q�Kغ�����rB�/4-	Պ誄��鹦1�a��C^�������v�K�=����%rm��p��WѪn{2����&}S�1�i�r.�����Da�˳�d3���!u���J��t������R����;��}�}gv/cnVF�:���*�^�F��V�m'Y��%�|o��"y�:�Ǣ�� ��K��,��3ĥcfʵ*��Ք۰�t�q�of��e���A������)[�)�I�8��i1l��'z�Wukr��L�3�|ĎO���w�כ���7���ͱ
b��jɧ��Csm����7��ƴ��Gw�wJ{�z��W���nE<տd�8֣�{T�����#���۷�g�v�>5�g��{��o.�ۓWwLC�/R����Y]���\^�(Wv�jW3����r�f�Z˝�G�f���/{ReC2�lT2���S�J�,��n�l�f]�V]A�s0�� =�l�d����m�����B�SnzT���ѓm�q�>"-*��٣u͐�������Tf|�*�C�xz�q�]�*�w��5�.�׎D�/�-���_����S���,�M&��ҹ8F͠�5���Sj�$�&孵����0�岉8�-�{ڧUjjl�m�Z����m�/MN��M��%")�Y�6
Q�U4|�{��ύ��4�R4��{o��毽ޏ�`�c�z�㛄k<�	#/M��d�ol�6T1V��6�
#��B��n�7e��V(6]i���6V�nN�UL���+��d��%^�Wp�:�S.�R�:iW�{�^\��l�:�nY	�BZ���[]��VRBh{!6�p��5��-ŗt����N�l�;��s�1��,�ԖC����<r�g*wM/�}_Zխ���B�;�/U{F����E�M��|���2�vIh˛I�-@���6�&ڰnW�Be=�5NDV�+M5zųa�.��{���3�����N�E�/�Y!{��f�%p�Q��Ɛ���v�ǖ��	Ӈ��{f�o�o��׍�����[i�Vm@�	mOZ7lǤ�ĕ�-gv�L*)���*k0��R��y�-P��x�?*���f���[����_1�B#s�<Ο{�-�}^������h�s�͝�K��K�ʹ\�$�C;����\�[�j�:iKM��Nٔ�f��s!�V\��Sꄧ�hnϨ��[d<�c�HF�y��5+�S�~��NOiu=����=�~��J�u_�zzT��Kb(4����i�C�_qq����^ศ|�L�{��e�s�y�9��ʵ���h����={�7�8�e�$CuD("|�(O���r�� �i�ô̜%Q����m5C�y���y#�� �Ѣ��pǿ]s۾Uk��1�Y஖![¹�H��K�>�Φ�y�De�o��Ue&��4�1{.c3p���S����2����j�"s/^������� 
_Z&�e��K��R�Yג3W�4I��ۯr�7�A0������N.���(CJ��"|� -#����8����O�r%����։�8����n4��ˤC`î�ǜo<�?0S�`�QĀu�iނ����Ǝ�6Y2;Q�Y3W�[j[�C�l���,�.^	��:s��}xԍK�DÈf���÷sc�lWNfyބ�`|L���⬷W��7�b|��3'v!�z�c7t@�4��D��'����)���Y�M�S�p����������gC\§���X5L{� /�%�޸��@�}9|��ݼ�����yR��y��(j�D�e�dS]9M�uf}e|�0�� .t���5u�N�㊹�Dw�B�AB���/�Y�\�O1�Z� N��N�w�v�Zqi��Ȩ��
��e�+<��{�qZ�ũ~����r�^�:e�����?\X;M�$TR�E���Y�4\E;�z(鍜��M�Z�'�s�����c��{ke���j��ծt�k+h�3�פS��O�!��l��0�Th*��{z�w�2�N�oS6D���'�]���ʄ:z*p�,��J��^�2�KA~�솵~���.U����K�{�pW��
^n���}�k��1;��s�&����)���c��[Y:�ܺ��f������(����*��L���}��&���/������^L$s�3-��(�ozh��UT���rS��={׵�zn�o���������=|��O�vS��0�i]RA�s���Y/�NJ��L�����D`�N�'Tpj�F��b!�S���S20�`GsǏ>�����XmT./4얽d�,m��1t��7V�ͷKV�>խ:�Ҍ��L�#�zP�O�Uҍ��r��bϲتf���V�_�*�(-{��v�w�N=Y�a:i�H�4�r���9b��S d4�M��D��K��蝛�κ��bzd�CfF�w��ib��<�����b��A���i�<Gc��ͯ�K^2�o�R�h�(sv������9@�Zx�E��t�(�{e�v��&X�i��4-��5���u�S��D�n�y%�Y�"�Ş��9X�
��0˜��؁�rj�l����?��W�_�۰�)�z�Tu桖]G9�*�{v\m�f�O��FlVV^�#Vҵkf�E�2��֍D�mˇ�C�����d�\�UoQo6W�,�/)��r!�����uv��&���^��-|��vDX��/����ptQ����KS؋/����G�dG��dT����7��J�;�wX˺k*"��ic���U�ҕX�4^�L^6͜aV���F��pPo��]�,θ�����b-}�W��Q�v@�%�$h��3YW/+��
X�V�	Z������{ϴg�B�NJ�u��}������U`����� ~��������,��g�j���˰��9�7��R����/\���9�OZ����O�f���9:�T?I��M�(\��K�iev#p���x�u(�gД�mm�cӄ�z6XQ�5.�q-N��k�X�!W���Btz�co)CE�+���vY]"C��W��OX�[9�tX⭞@veK)�Y���-N�7�3c�
|آD6��;�{_��*��}L��j/Dt����r�~;��:�*���T�i�S�Eq�6K��7��&�2MmEB<���F�ġ��'B<r�����\��ŭ	,�`O�A�[x�h=&S�5����ytP�m|���ێ�Mz��.����r�۳�d�@+�`Q��R�	��w33zG3P9��k#�?#�Ց�K;���u�Ԝ��T�?<2ֲ����`�ǃ�4��#��_Qn���0,K:ۚ�e�M��:��(K�G9�q�q(�WU1�x�\u��Z��Qۗ�tû`bycnF�z��;;D���^%q��eF3�����2�?����M�{�?*3j.`87h��˟�;��N_c�L �[�ux21(Տ��R���R�QK�?e��e�N�s��Q
]�����bn�-���Lm�h�3��nY�i��ғ%�lB\R��:�iҩ�Y�=��)a+�
GIY�e��{L
�y�ҷlrQ�5�_}^�n4���@�_� J�� �9��F��ɀ:��K�f¬�f%Q��즁h��<�.�=.��<��k��As�ݷy�Y�8�ʣ���D��F#w��^��/n��~��ĊSL4�we�Op[&ݱ1(���p�f
���﹟�r����w�=�S<�c��k����gcs���Ϡ�z�@�P�7\�a����M��2%�̆��&.��m�Ys�4+p��ER�0���/K�8*Kѭ([��]%��8	m�Nzo����.��N��k���ܐ��ս��D�$�ۆ2z��W��dͧ�[#���dg��2�<�L���ǃ�P:��v�����8l�裮�@�QrΚ��k)��>�~,������}ۛ��3� �"�/M.�:)��O]9	�(M4RUL�N�������43+=�7�8�kU�sɾnؑo��A�+�2���V�px���:L��F��df[mqeF��^t^�{2d"o�c�J[!	Ԕe�d�aO�e��L�x� ,Sg�[Q:�)<���o|{h%�����@`��G�.�l=Ȧ���5�s�{�b�nߥ%^�:�*wpj�P��{9Ll�]���^����p3�t!�m_�����D��A/y`  d��E6�i�o�h.�l��j�qWu����.G���BEYմ�W"�:�=av.��6G��F�3F7��l~7�o�I����?��h�R{K�:Ge��G#:�4n��q3gF�����>׊*�z�sY�vՖū>���7�!Ĉ�B���/�O�l�VN%��0�89W@'�E��%���Ψ��p;ְ�)��ɷ#=3t��|�L�{��e�=9��^�[��'� �t+�T�bv5�h7��@p�1BY;�"�H�1b���L��&�����D�2�l\q�֨���r��9��#L�+Js.� �]R�S�9� -2zcx�LsJ)�	m�kKf��U�d�u�\�جp찧�m<�y����O�;��܁�;��F�T ��B�w�+~��6Gӆ���'1z�NG��^	B=�:s��:\wg���m�ulT= ��dGt�S���2�9�e~���m��7�AO���G�G͟)���耸��̞n�x�Zvj���Q������ ���%��n�5rʚ�"��\q���']눕��
����i�ۙ�Z�]��=���%Qpg��	J�>��#lˬ�*�2[���-嬦�p��c��>�2��j����ī��h�#���Pb�|Ѥ@ɰ_d�]~�u}�[~�t�� �E�5����.Zg��=nx�l\��9UWw4�n�NU��R�f+�]0�v����s��5��_VS�É�9	p�X/i1G�@�/'jL4��|�o6D�.�C8�t����|8ܮ�4���/i��
�R�����|�7t|]f��,l�E��j�<6_������y�(=I��[3�N�{%"z���n�"��x�[�F\\�b����GT��wZe���J�6;���$G�l ��
5���l�W�����v���@4M#&z/���Wn3�ٗQ�@GTuN�$���$$e�TP��Zn�;�8Uj�X�mg���4��m�����$g�2�??:e>�Si�Z��jwAi��~
[n�lO�r���j변c�QQ���4s���{��X!'�΀X��/���	����N�k�]��'�]x�$�GU��\V�>JXx����l�ƇL(�Ɲ9��e�H�Q��-���SH�{��_[3����QWaf�nΆR��Y�t�#��j��Ntcs��3�a�,�\�m��j&�_�O=�{�q���v�̌/����֟���~Ol�)x� K>��c�~阊�Y$�f賾!H���M+��4���t+O��m�L���t��e����ܴ�0b^Ŏ��%�U��å> �̭�7���]:�X������R��y�f��U�^�U09��<������̀B)C�;8�H �6�v���.a�-�+���pn���M���]Bl�*�{������t*s� S�����9k��,�Ҭ�n��J�{F�Hb�-�7�u�kk]b9f_�8���6+�u6�Z�-ͅg��
{"�q�6��~�J����5l�S���~њy��m͇���'��Q�QW,�_��d�5�.1�0�����ø2*��vm��4c�*��ꈀ���H���@Ⱇ��yqSaW��-��]ּ0.DV���WwQ۴졇tl5K,x� Vs��vt�	��ܮa�a�=�,�����>�%��P��N�
�N��}�#
�)?a�5�0�c�s��܅��ݵq7�OE��X��^g�ovd��I�+^����e���.���(�8+�O�fӁj[!�\�B ;n*�Z���6���e���e0���~�y�q�2]\U�'Sݓ��Tk�É&��1[����j�A�u���w
-�������N1�)/�}�����Yϙ��Ӵ����2�~��h��}��)lQ"!��'�
�����>�֥t�����
n�(���$��b��,ѯ�G��S	��O@��Ԍڬ��Wy������NQ��vγw?a�S��ã�֠&O(c�8�|S@c3>ҝ���I�t��VZ7ut���-iz���Ş�5��g0���@"�s��*&[�ABcn��įi)��u}�%�w��kn����oR������f(4�]�p�6�݊���l|�� �⠼����n^=%ҏ
�5�x���*$c4��8J�Z�{b�G9Ww��i^�ɾ��:>���r}��p=VJ����-"�c�x�i�t�[�̢j%��Tw��f3L�j�p!I�֔����o-��f&ĸ���Fp9�Y%������\#Tn�j��v����c[+����}J�;P�ss%6��n�U�K������N�έ�χ#6uZn4�$��6&��e˾a���\u��w!H�c.�2�U��f��1] �@&�2V�7�Q�|n��Wh7X��D����+pR��� �auk�ۦ���-e#
7�ݕ����:�tO�-ǑNG�(]�4��t������Lm�|����V=#.]L�3pr���`��V#F*t)��6�CP7���e6A�O@u`-42�S/9��Glb���#9�<`�sö�^���/i�3G�9vts޲��d�Q�e�@�kw�]�b�R�P�S�ElE;o�2r�a���	�!��v>I[L��$�F��K�*���W��З�����դ5����:!H:~�u��T��fR`ۖo�݅�+�H �>�+�a:� m��t��Ÿ�2J�{���I��$փx���s+��r�N��Xoz_nV�x�g9���(�n"#S���}K�`�ȼ�}K9@F�O�8{��F�y��Cʎ��8(1.<����s��Wp ��:f�,�m�;}י:]����9�I\fU�^0V��Q����ET�`mm㘔B�h"!v����u*h�dd ��\����poR�X�zM��yGZd�<csf.�\?�o�xR��]F����҈�`�)��m�f�$��`ŷG�@�	.Z�I�y\��������V&�In�Ŋ���^Zk��������>N�[e��r���׺�b'v��b�8�qj2]9շ�Y�f.k`�22���iŉFfG��T�b�.�Ph%r۫�0R,-ݣׇbN�]��"�K�l��B��|}�<Ÿ��
�%�Ҥ�r�e$,gf�u�'��7g}�w!��Ϡ���;�^/;�rF��̕����p�=�d�f��u�B�6�R������D���N၊u�+ &�dVR����88�r��}/�RX���n}f��nc�����`��p�V�p̟X�Pܩv���GeMK�KS!0z^�i�ܨ>�G?[��+e�kswj7��r��͈���ڬ�}�\��8�#�r��:�V�u:��79TRU�pgY=�������]��q�JD��2M��/���&6�U�{�{x�GK��w7z:���땶��#i_4t�jG��*U��\��t��3��)�0��tWna��z��f�R�̼�E�܈tO��d��=�����Ͱ���b��)�!i؉�+k5��n'�?
��h��,�K�״]op�^��h��"���`
�bk��E�ZAHi1,Y��c*
�W���TR[H��T�Z�XʢU�aX�77MAb�ȸ�q�� �U��
R�G,�JbVT�`��Tr��*��b$���R�b�1(�11��붂��K��.�"�V���h(4�*#�ab£���R���˴P��\�l��L�T�0�,X)E��7*�[Eu�R�dR. �3ȫ�2UE%JԨ)�S-�fJ���`����.�SmACXVf[�Xje���]�fDQ͢&1��v�Z����V`��pB�n[���J�
�3PݡPSQ5���1���5+\p�aVЩ�����F�$51++1�+YED\��P���UB"��n��"��]�sS�$u[�SY2�C�)?��r�u�gl� �{�P�:Ӱ7�D�c����7�*7qJ��RߏFC�s��y����mՕiŕ��݌6.zJŊF9�H�֐x�|�Vd]��;s�wj�툫4������VFOa��χ^��zU3��������;PVWjP��r���Ά��8�o�sB���wl�|c=�#'���d��Z��؛�Dn4wF⋪� u��a��$��$�yf�gl��t�h����f��m�N˘l�X���x���3R�hO�Th%��@�U��K>�Ge�s��9y0C4�IsU��LJ��▣P�S�b���]�s?yd3��o�����ʣ�����K�b7q�8:��t�dШ�ز��̮3ie�"0t
.�H�l��IN�˙�e�9����L:.>�?#{猟�ghl���a���c���k'S��}7̞����^����5�ԣ�=�<�n���ۤ�A�܄�׺��t�0�JW5�V+�Oo�|l���%'���m�s���Bܪ�)]Lf���1�n.����i�ӊ7,�%���e�Q�fӁ}-����Sjy��8�2j�x�1)�r-s�g�tX=.�͡W�SO)7�m��ׯ�n�'�7�Ug����z5��9d�>S�F:�"�*r��]pC}�ً+C�hSB��b�;�qu��+�x�w ���>�r���k|�j�:r���j���W�}��j)��.�v��dFPrp0f�a��m�ǘ�Į?/�7�(\�f0K%b0e3�X��Q�R��{�{�k)��-��/2�O]Ed�eNKfO*��B+���Z_���7:���Ӑ��,���=IU3�;�v��!v��Q/����T�~���2#Oj}�R�q�(����]'��d�:�О��f���R�R筋��;�N�&GT���N��Sc�J[&P�i>��5�XN��P貯w4t��1N�V����s7:����ל��@��q�֠�gVƉlO�r��Y�]=-��t��:¡���q-�)]V���F�_"��N�vSl�
��@��Z^}O�m�c�5����r���~V������~#�TP���)��kɷ!,zn��s�κ�LL�{��e�s!�h�lwq����5j��DQ�o��@ग़����rq����\8s�6*��5Gb�a�§=.�#o.sv�+����-�듺�� t�9"��H��㷓 \%xGj5qW���,F�7����u���EF��Xy���8�y}~a�:`�)�r��/�w/ة�I�~�٫"�A��y2h(`�YH6��B�����5w?0;ѷ2�at�|S�!*t��U+mpog��ݦE'"���#�0�#����,�jP�+J��\����I��|K�`%����f	ԇY���w����,s�_GM��o[��1|�:1�V�%#��Z��:_�Osܰ	W�����Ͳ��ֽ��%8�{ ���V��v[��;�b|���l�34����O��'u��[M4���h�u�.9G�^�D�U�p�7/�-�j�YW��"̵�� -�:8]
mh�ࠛ�n��tE���Gyt�F���2i�m����r��aY�u�EWFKv�ޢ�l�/��0&�	1�˄ճ׊�oiۥ�f8�򈔣�#�/B1���	or�#0�c"�:@����Q8�%� ��?le�o��v��q|���7��y�J��O��R׌��8�Y�R%wE��:����lv�����Z�⻔*.'��xf�֕��x�$F����9�Y-u������k�8�����������=�i�~���Q�>�}F�Cz�ұ<�j셧!:�{ i�7����^���y�d��Y�����+�xl]+�:��\U��3�K��n�.
[n���}k��;ڌlkG(5ͪ8`���ᦜ����I�:c�m���KW��Y�{������­�H(��F�C����\�J�/]���n6C���m*V�Ɋ嚡�s��oN�2�PY�)��u��!f��4�_o�5�b��>ܧw]Oä�r�wB�T0�;W�ޖٿ����=��[q�%�
��	<�	`��B�Z�Y��U{�N��{�3L�?i�9f�uJ�8��e�H�>\v��c��:RKZ5�*��ζ��eVJ�-��C�zb��y��;��t�'Ut��!A�M���ɰ�!{ ��7�*�W0���̛+�z6Ͱ�ۙ:Y��5�X��>d�pL�RԨ�AȊ˲u5�퍶�Z�n�<x>��k��zi\�f�~�
�j��xX:G������g$,�j���r����S��́���=y��u�wj�=�3UE��*�D�!b6��K�O�����ö�U���Ȯ�k��(ˁ̕t�wN8�0w��k�rʙ���Ǭ�%�qW9K���n��p���6nþ���lQ� O�~�^7m�p��qVK��y�	5�E��R��S�#_+y߸Iw�8�t��izD	��x�;Ћe�4%����n��,�G
����*�.�d��tg��E����}�[
XW��y�K6�%�M��Z�����Z(��_]
�[�[n��W� TR�]>I���Z�d8뜄 }S|�v\����%��%y���^�r�7H>�f]G�}u��W�S>�ҹ�$|;�[i�ܦ#˦w������"uk���%�:�r-�]fcî��*E����t����7��bx`*����q�`���V�s}c�-ɇ�b��p�Íl3�s2��w�*򶞌�E�fqzc�����{��K
1�J�ĳS��W8��!r��"6��%�:����j|{�ܗ�G7.C�}-��e�^�;O��y�*�yj/��<7�����T�/��<f�"9�v�ù}R�	�D�خۇGk� �,T =F�Ԫ�Q�O����g4�^ʚ��;�?{��T�J��^�ٖ���5�=0"cbQ�fN�c� %M0(�Xr'�O�w1M:ݶ
�;�Q�����h�Y�v[}{��׭8�]=-�6㠡V�����d��D�;�^h8�Y�Ew�fK3�+4(�F������0)�a�,�z0�י�OOK8�ssV.�ΔJuR��We]C�k��v�D0�׍S00K?u�
�Zn����l|��#,Ǟ��BC�NS��Q��j�k�X�YT�CuBya)4r2m��ǫ�v��Һz .5X���©��Ն��k�̡�!j<�w�zb��
}� t��8B+\�H�;��s�D�8���Cl�E�Jɞ��M��<������x�>��C����8�����D��F#ws���ғ�Ȣ���r�^���)N�h��6�<�Wvy�������4ǽ~�6��c+�8�*�K��y�Y-kiVx��&����G*���6ܻ��ZGB���3/'e#�R
V����v�Y53Y�ɷt�F8!���U����q���;�ꤩ�����M~L�)~�<;\;uk��h��s�<�&xu�?1���4s!�?۱�*�kE�Y�Wh�QeY��q�>���GKp�k�)?|�x��sA�d�F-���;o���1ܷ�O\}p���Km�yIz4�{}��3��m�Nz;%.�j7nrjk��~�?}<�Y���$'Y�h i~2Y\���N��p��,�Lˡ$����'�����_��јU{�P�3}e��c:v��+���n��K?)XSG7Z;��J�����"��`��(��?F{���f4O]�	Q��`?{%-�����!���=��{�[���}\���R��"=��>��N�����]r�v� F|��U�.JKn=;�}�ۈz_�*���Ύ�(��F5;�?V<��ЁmIFY�-Pp�2��R7!�l�R-�uM���NV�0��S���Mʎ��>�yjt�Ϯ�"��z�������C�ՅN[������n����'��)���}a�M�0(O���N���?�Q�P���%�������w�c��ܺө#��*�B&����2��^Yv��CwgV��av�}��X��ѭ΁>�i~��O�l+�H�>'�(���V�*�ܲ���k���b<r�O��y�\˳ە����o%Z0譮���w�.�V�m�>�ȝ�3�v3h��nR����ˣ�YX!'�6�jǮ��s�κ�D�׸��\a�˩�*jb��gmn�/�s�Δ�F��J@५�H�U��N8��6Q�k�᧺lTsK��=�m�5��z��'(ǳ����#L���9+��]R�%Ds�/��,zcx���x��y�uALd��Տ�O{�f�����9@𨭑,��>�Cc����7C���@޼���1�*\���.��G��h˶��ödc�������V��J�:�8�ygׁ�됽�nO(�����]�������{�w-�NJ�aR�z���F�up�٘�-����\�0�Bօ�}�Y�U5��Q�a����u� F��טOS5��X,z޼뻶W�w�2�4T���i�i7}c�ެ��@��ʋ�+�(O+0�n� ��,� ��j��n�[�[�9��٥_Y�u
ɺ[8:��~�᯶@�F8��Jx.7�ً����$]�hnϣ�
�͖��9�b��ۺ'o�=:]�ۚ�ŧ�.:�K���w�_�=w]�eg\��f�H�-9��~d�o;Yr��.�2�#���Q̦ng1E ^X�:�Mcdj���G�v�j'��V�t�Q�@���.��"�V���D�x�N��n��ש#Y�m��){
�2:�|7e#�bD�}����˖���VCM��
���� ��"�pT��WW%C|�?߉��GQqD��;��X�K6G	kaև�a�e6�M'{[�����sj�-�����Z:tU
�	�}F�C{["BF[Ȯ�Zo��e�k3�Q�|��x��ȩC�1Tz[)��!gN�YL�-L#��RԾ�4��Y/�Wv-ʆ�&�)���QZ��a����<0K:��;RQL��~���h.&2�	�����6lR��ɭ��Ń4D�vT2�r��-ea�k���#�R�	<��P -(�|G)�� ^���Xb��6-���Z��a���u�nݷ�n=��RPx�Y��,�ӝ�0����m8�� t�N6h�
 
�JٱB��m��0(tfF&�]�<m�'�
Y��X��`Wi�Կ.Q:y���z.�gV?C�:�&��M+��H���Tk�<6��F���ޮÐ���T����}<���~J����L���~�9�{q�(��Ƿ6�U���B�lBx6��8at,튵`Y~(�[��'�q�OPr������:�6�\��~s�k*�z��N�-�s� T�6;����Y}ˈ��݋�˶���I-?��/��yM[�Bm���.�
vk:^�F-�O���*�c g�N���!�z���L��˩�����6,`�U�*�f"h������`8n��{n[:�XWG��e=�"���3s72i���7L�	d�p��x�wDp�dj$D��"!�t�+>?�����Y�w�c|:�+�ZQ���x5n�]����
[�D��x�dE��2��OϏb��E��:�N��𫅙���&�'a�_7DW�!��Zq|��P�
XCc�s��ɕ������OE����#u�h��7#�I�$�� U'�<2��M�,l�r����Q�V@�l�^�q20;յW\RƬ�yk=c{r����]��5�t�d�4)aF��qmN�Ƹ��[!�>Ή������GT��U�[�h~h�Vv�t�!���FodO,��#���-@E%T�4_Q�w�kaOb玚��ܫ��z�sg)��Q��*�8J�ٱ�N���� ���F�ԦX<�##�j���u7��<C�#��6K�,Q�h.9e{������v���kP�'� ��y��g�FOs�֤O!<��@Q�:)�;v�k��[r�ޑEtt2l�Pxv����s'z�i�i�ɶ�$�<����S�|�f�1�Z��٬�
|��pN��ןRp:q��qk���㰳��xm�J�[}�k���Z�vkgqW`.�����1.i6��r@��e��mr�Lҩ�JQJ$����kW��1X������$�-
�M�k+0��C�RGq�+X�jZ�d�b��_�r`a�����Y^]�M=66��s=ҳ ��f��u��T?V{Ke-e�#-nρe5���,��4+�]i���tc���.�r&7�ft�N��}{ݲ�:�O,%�@�y�#{�坮����q��eE�A�����G�^��fn�v��sv�i�ϡ<��p{� ��=.��xs��9m� tMT�.oʾ	����z��d�]�G��1Y"#.i�z ~3��O�!��9xhP8��/�ݹ�A�+m��tu�i��";�����B˼Y���G���.g<a��p�
��ɇE�/��̶@����M���qY[z�5T�ܰ�}�/�"��5��8�/���n�T0�~�~�x6s�\�v��fq�g��1���yneA�9�7,�%���+
�t�fZ��ǖ�@;k� CgTp��-�c�Dv�����?k���TP�3��R(��⍕��M��rYU�l�D
��G .��:��~�d�,�'E�k1�s2������E6�a����:�C
{�B���3ϩ���o6�m6�=�z�r�o�'���.[v v����(�h�v)��t�u��1Qb�����=�j��_�9�h2���z����ޝ��,��k&7HWv�l�r��-����,��Z�v�\]mg[��y9�ݰ����oU���uo�����N�c0S��R��Z�9���n�\TE賜6����X�x�ʝ�I|킾�9]��[cK�����A��::���pE5�3Mյ罝�B��*s!b�N�Tyx��+2;�\����m���R�/�C+;�ҶJ\��\Vu�6��˳ON�7p#JN��Cq-���YG�M����f&@e�6�ڎ*��fثas8�PL}��*�I�Y-`=��3�\�z��r7�aW�fΠ�X�od��р����@u�bYp��wˬ���E8�g���>�W�\���ݠP�O'�-;6��v�j���*.4�T�6��fܼ��X��r�<R�Wni��>�Hm���Ϣ�*`�� (4,u��]�o�؛w2IF�A�W�������VWs���j=}b/@�����2�_(8Ï7�e6�2�Sogp�ꎮ�s���ؗ�&R���j��Z8݄��.�r��sysz{�/.����ÍU�:��.�0��*'4GT7f�Z���
�O�.&K�-6	��U���ʷ	8Ae����v�r*����qv�����w�s�R��J���R���V;;[{���.�Nݮ���S�i�wt�C�m���eĐuc	1��mf�&�L���GChA�	����OwQ�'-��$_I����,���u�f��s����_|���A��˚�����{�b�)���SѪùW�n��DL=���wq��T�xVVuio+�Aև[����C�,M�NT��.6��9���>c�.����F�v{���}y�zo�e��R�E�Kv��I�Im�8*�mm�g�1#�9�DK)�[�K5�۲�ín�7��@յ�l�].��q-�9܋�3Ye�A���U�� ��E��P�A�}�2�|X��ů2�&�U��%�O%��wGl���\�ז5�![�9؎.��"vb Z�A�]W�љ�j�@Půd��d2+�)��;'���h����3Р��m�1gopj�����փݴ�X��36�ú]�B#�|�2n�v��.�Wp��{J�P���ǩ�W+���]������AL����8���d}�����̌�&9`Fo1�	R��>t��R�2��,ެC���0q��G��.�n�;N��f��N�oK`-�/�;��!n�-��E  �mZ9|��o��1t�,�Ǖ��r���IT3=�#��"R�?f|l�:�*�lT`vU*��+���;��ܡ�¥�=�6����׌�;�v��lh��
,���B.�e��+��3�|7�q{=�X�����ٹ�pT���ܙ3=ں�}%c(s}�6��6,t�
��[m���`۲j�ĕ�ʁRר�q��Z����khP�]�����,*��`Ȣ3n�a�I�cR��B���b혅����G)ET���.�CK��b�1�0C�`�������`�ܶA�CTY1�n�r���
��*�i��ѓZ�*�3��S1�nnF m��&�QVc4��e���,aR��Z�X�U�LJ�#e�ef���54b�j4��f[��Ԭ��H���I�Q]c�n\Ki��cAB��d6�&Ҭ�ˌ�AH�����+i��3S3	�CJ�ĸ��ʵ�e��e-,YP�*���X%�X,�1�٘[�cZņ����1J�]�
�%c�qv�]6��,̢�f�s�s2k�ݡR�A���-ce�n4[qr���IXe�+UTAB�~�g;����9�fй������|E�.�_kyq���eȕ�/1�e�b᷋�r�9vt���9����B�LJ�����]�T����ֻKS�jz��)l鑣�>��4���Pם�x�^I�)�r��=�[Ѕb�g �ꎲ(Δ1��i�ǐ�:-�(�4��2�'e�z����UM�f�����g�g2֍�p�l��P��-T���#�O#�կ�q?i̺�~�������)��7�&���,���F%��h�#�d	�u�嚟��j��T��#���k�����a	Y���5U�b==*\J��U�.ycnF�~�⭟:�+^᫤��-����#m�nc'����,�q���rY��8)�� *t�_B�� ����0��]��Xb7n	�|��6aHc}s�j��cCt��F�bW�p7uK�N��[3� ���kk���u_����g^��ـ.&�m�
�{�	����]�ƺ��9�� ��l�ϼ�����]_�����ϚAw��p��u5�si�tK6G�mx%�k��\F��<w���o'a�gUۉ���m��L{����԰�K���v�S��uך�*�*���,؟xk�8G�f8.9��� H2� p,�����x5p�RbYK�����K'�#�&lsќ�Y��;@5��uX9���JS���F����*v%I{Ȁ��2����Mh���y�J��0̶)�f�%;�b��u+���X�ч@S&q�<x�ލ'egL��le�Gnp�ܠ�~�o�<+kѭ�1��f�J��u���zC�u�+[��9��"+c��>nʋ�><���n�#l��D�E�v�5��4T�ջ�u��?2<���+S��c��J8b5�Qb&����8lg�����T���/:�k�c\��_�������I����,n�=i廮�g\\Umx
������<����c���ݞf~��r�L�QJN��ӿiU�w'�$F��aF��T�.׻3J�~��S���5T���Rx��ƈFY�֔�4*�F���jwCz��!#>�Q@�a7P��3L��Z����O��㔛�mQå�4p%C,�	�ӠS�0�i�j_Q�PZd��{}m�qf��ݭ�xkT3��3L�?�����Y�����r��B�G� ��^NB�aPv�#���"�-���g;n���;�;_s��\�q�:ƝY�7��{�S҅x�=@����^�QX�!����1ݡEv�͊�i4��=7p�/p���'N�'Ut�ʢ�-�`��D-y��t'I.�_���yL��u3�Bs�[���6�K��/�A�=�y�ƮJw��3����SO]��t>OB����˴CPB�ov(_�}V ��pQf�I�k�x4<��j��=�#VjPqK�k�hW����m�c���b�Q�m���|>g��wiG�<2us����@5zSE�K�켦-�U�\��Q�(>ۈ��+��,ԟ�e0t*_����8�=B����]�qjǊ��
�����`%O`u�c�x��w�~�r�5Qna�ʳ�,�X-��»�W+m��CL�p��={���8�2��r~wq� ��`uerʮ����*�����ċZ���E��p�C��k�Fs�x�wDp�F�D�m�p�ܠqXk�0�5V�������i��6��|`�eQg�gB.�͑��-��-����wD`�nؑܮa�a���o^�ꆜ��g39���=����<.��+
�kzfm8�|�R�������چ�x׈^M�@2�;�}t[vn�:-ݖ#�ӧoj�U�xg��$ͧ��!�\� �~���;�<ԍ.�im��~�m>Ċ�U7���A����z�!��5%R≾8���l�\�_igMW-.[���svt`y��g���P�Y�cF׻ BygOA�~��!���g�������	�)~"�{��ft���	�+N��p�=���t��_=,���w�Ʊm,�K:sb��&�ܲ��:�@���>M�J��9pN���h���i������k]��\��w3Azɏq"e��cV�Õ�uu�?�:Ϟ>�Ƙ����W���S{��G����H�m��w/ʥ�B/�
;ٰD pn�ѯ�.��UA��N�v���/�;�P��#��r]��b��,�W�]��gΧ���tr�@
Ms���"�c���|Ŷ7��蹁R�MF4��N�٧��63^n�م����[q���(�Fgv>t�������'� v����M
2�C�S�;X����χ\��~;]�
�9���U��'���sfM�8�-��ʽe����B��qC<��4���L���؆���۰�4��Q�{%�*�:���C*���}�'H޷�\���M+��D�7rڂ��"�o:�5�u��n�#���?�r8����Hϰ�a�#8��& ��O�7@)F?_X���r���׉�:ದ΃7��,��!r��/-��g��M��WC�T�U���ic�d�G\�T����Ւ���!�6�C�1�0�b8u0U Z��ƴ�/&��n6ld|����3��x�C+�6>�����|����[\(aJ8�C�:�~�����w�HP6�:�g��E�{U*�e�݋��80�9�������)q��e��zj3ۛ�r��� ��Gq�M������;f�iU���
��F�z��E�ݴ"�PCv�.dX��k��φ=��sOV��6.�d7j�c �3�n_�[���5A�Mf�_���57�yK��]���Ӂ��k;�1�o�	=�\��6�������{�����h j��y5�A~�/���j�!}�έW��� �݀ݏ(��Q�Ur�Y���	J���g�g]��6ԧ)�[� m�7v^�V�5k���.2���g@��Qzf���wb�͉Θn��	�P;��69��9��a��=@-ٖ~jw�v�u����ڟ`�Ju�|��Z�u�������d����ߚ�=p���G=7L��P����(KS����y	O�e
�>Q��a猝��k�كy�_�LK���3���?A�+ �b@�u$	��]5:Ge��r:��E5c����#/� ���f�����(�,���I����E�+�'�N���?��]OKĻd��vӻ)FGy���]9[tA�OWS�d��t�K�Z�H	c�K�ӝS!Rʎ����aڞ��[.K��y���E�g�7�2K�r2y��J@঺���Kr��	6Q���r���ȩM�\��
�v�rY­_-$�v'�(��̅�K<	��+%ụ������qR�Ҳ@�]��ܨ�p�9�N�;hU�4�B����R�3%�q`*Ym�����Ŭ�w��j����)�0�����mo�뮖�5;q��g�ݻ6*��Ti�Tc;!�Y��4�5��)�y�@
[����y�֞�Usaɧ���f%�D��o�
v���0&��P*�6�vQ�Ѯ�ǜo<��0��	��^�m�����ڹ�呄��t�1x�v�7����c�����,�/K��k����򌹕�,�_WaS�\2���`9�Q�����S<�u�S��er�g1>��pL�ln�Ͱ�k�u�M�ٝc���ԡ�����/�lÇ�Ptܳ�Ku�f���T�QK�\�1��\�T%-�ٜ=u���6�k�q{3�QpWSȾ�Ǘӄ��8� �x�z�9���ݝ� �C�5w��,�@R|\6���x�fJ8b=��#��/�y\�b��Z���6-a����bHn�6� OR����w�v�����<j�0vm�G�ģ֞Y���g
���WY, ��nuNs�M��J�J;'W��Qq-N���V�;���$j�A�`P����L
��N�gk��4{"�Z�ܮ_Km3,h�e�="�����P���jw�f��ެ�	|m\�B�o_��yx�ϐ�.����t%�(Rs����p�p���z$����+܆m>�)h��cE��4��Y8s.�!;P]B��[�nfgbM:}�1�Et�}�P��,5d�]\�kh�(.y�r�pׯ5�r�ɣ5�"9�7r�ӗԤ�}0�-���!9E ��e��z{�@���Mާ�l��r�<�d��ӹ����9Q�W��kO�2�O��=<&� "���}c�:wM�~�b���V�D�0�eQ|^�.��ʆR�Ѻe�����5�=��(��+l�	1�]�	J��޷>����1�aM����y�Xbn�_�{M�t�#��uI�-.ېY�<�0X�%=U�����L�v|FM���q TwE	�L
��;��]��~8�b��o@��ޮW5tf�׎�'����3u<l��9���vS\�"i\�jO�r�
[Ouuyå�-����_�Ǩ·���`"Uq��k��lWo�n[�����YVzǉ}�K��U�b�ph+%�o8�v w*��B"��m��f��J����t�Sc��LD�d����C�f��K��n�m�����3��<�8<�lH����*��ι�WL]2�u}�!�K�h�y�F^��΢\Ŕ�GKt�zD	f�~�>숱��{��
������׭jˑ�^�/)�b�SQlq��Bہ#X�(^-F'H�:y�ͱ�-]�K�\�x�0s08��x���Y����N�	���zr�.��Y���ؼ��௤M�$iyҥ��{ޛ7⫦r6�u�&���%|�n�ݻ���5uR�zw1��S��s:�B��p�G}i���a@Vǧ��3m��3��E�]�K�ȭ��/i�{�YjeA��DI�u N�WD��^�|�6�R�:�! ��eT�bug=\�A�tfM�(\��K�etl���,�Xц��\KS��p5,Op�{��-c��W���$g-���A���ovR/�a�o^A�}sA��m)*�~�ռ{�u��-��i���|�6;���D��}GqL!�{�vlvӺ9��)f*�L3�k�;%pj���hp=@w��S	jz�z�}�씶)�2׎��7���_z8K;�K����{�iUF�E���<s�c� v�D8�{��%��t�y�:Ge��(͌��{���Zp/޹��Ӊ��5!o.�ho�r���>z����K��7���\�K��(������s�:�a�{�N�n7'�����α�M?y}�GK+���ǋ�ڗh�5����S00K?u�
c.���t9qll�g��Y-]u��������O`�<�j�"<��	��ύ���r��J���X�]v��N�ŴS�i���q��ֶ����K!	�w+�μ��6��A�]�U�ʷ\f[b�Of��Ǉ.0�fA��F߉��ætx6;�B�!�v=!}�:=�te]༻������%��V=f�"�`qz ����
��������Ku٥��Ft?��Ɛ������#��� ��g=7���Ъ�]�+^2џ�ȱ������pe���OQ���:�p7��p;���Ts���W���s)�0�.�Q���� {�]s�U�a{(Yw����vQ�睡s9�[ç�qf��ܾWe��7}L���Q�g��Qg����g>���GKp��
TVv��T3a�m+���m����e��'�q>n�,�Ɍ�=tܿd�]y�ⰡWOf����@	`����d>���Wn;%�f�Pz��E��e�'��4���:�cFZ�rY\���ּ
N��x/:y��vv�p
��4q� ;jy��v��Tk�1�Y+��)��ŝw��p:��O��]�f�s)��\e���[�\�: v���ϡGF�;h��{�-�pBMeN�;+�Q.֏NqQ����LzE�}4z�U3�;�;M;�����Ήõgh�~�Wu��C��f�c�#�l�Uq\�s�� �2ΪOM�43uB�&���-N�OV<��Ё=�f=�'&�v�fl��(���r�!�
XGZu�k��t�so9_&��ȩ�y�u�],眯K04����_��^̻�}k�u����;lN��aorbܪ�F�����o2�Q�����Wܥ�k� hG.�g�H̷�W�rL]�Q�R��BKJ<��||omz������$$�+ƍ�2�Qj�x��:Gg�qC��y
�U�ى�v���������78맩���v[�˄�X���0(NB�Y��ix�}lu5d�{h�ڨ���-�"y�'�	t��[S��W����.��q�R�\$�m�ŏM��,�J�9�*9�ຸz�Ʒ�u���8��{�k��g1�c�O9�8�QC��t��!Aݰ8�ב-��u�p��jU�'|���`�JSb�Z�f�Ta����qd��9�] l�.�p�%�*0:�S׽[tv��k��� Z#a�̘��Jm�	�'�9^
���|y���?>Ė=�ơͤpq7�uuZ�߭�З����~gXd�F�o�V{Zކ9�Oc�V��W&O�_�?P�wi��A��~�j���n7^_�u3#R�G*&Crq��L�2�u�x�,�_��>�\on���5�q����{yT�b�t�P���M�Y�n��S�x�FH�d��Y�%��z�Y,�y����T�tm��r�p1貂�oo�}t;]눖��nʋ�,ˮ(O+0�o���/�.�E�jj���N|��N�1�͕�j�[��%6�nS���r�Φ5��䓮�<� �{"̶pG���V��{(����>кt�ۑe����ݳ�����n�ii6񯽱#ؕ;�}	�G�p�� φ�+,�)^-��}6��s�c����!x8�U�w���Q�Nd�Krj���K�r����i�Ts<�U����V WMW��wF���[�\��Ϩ�}�Ճ��G�aY������e����X�pβ_�W{��(�^{�{O��V���t��O9����|(�����ٞn��!���z�+ދ_ 3o_`�Qʀ(��tfa�o�BVQJ���6�����w
]P���,9lVa"���5�ޭc��!)c�N؟v�[�'��>hW½y����xP�\���n���N\�3��ڏ'�3:�;Χrd�b�K}6��+�[���?�ި�[k;�/������n�I��ٗ���[b�&7���a��;؅�o���qH&w�r�U�:��a��2���N��*rmBP(0�Ge�ڝK���Y$6��?�I#�۷��쳊�q�l	uҒ}n�o��Ϋ������^st�M��c��f��5�@c��*� &o��'�X�3��LN���;�� ��G���՘mt�|��@m8r
��u��{��u����;�D�{]�4SSd���tEb��wr*�6l��,�L���ɉ^�#���� �y�ܹ9D;V�U�2��k�a�f^+���F���9����+��v��X���������0��_6�I>��|.�5��x�*���/v����%},�~�I��D��Ny�h�%]-�{��n��N	�Z]��dg�Ǥ�A�͇sr����� -�:X����54�o��ӑM��9��Yf�*�j#r*˛7�՜2v=��=�����%��ZaЍ��-�Q�R)��n��u�$��f�,�=�[��_4ΰ�`�vuM�7p�ȃ�e5u�IH+e�,zIVMR���=�t:�U�̱'-�u%{����YG�|xЁ����Rc��~<̃PNHc#ha�޴�Z�oK���\�%��]����ޱM1W��������*Z�^h3E{_s]����n���Mˑ��$cq�JI��Cx�m�4����#�Kmu�y�4�h�i	��4��Od��33q^�r�|��W����Zċ�[��C��Z�K�(c�r�2-�{[b�}9%�{�HC1���:�aԵAi��w����Bnj�Rb�|�YL\�uw\1��r)Sl^9Ơ�.�Ǜ9�e���{��XܖI��{o�W�`|�Q�6Moh����ad���p��E�Z�:�_�E�\${�̡��yfWd�a1oB�{�"�Yu��;bn;�1�7�WIYU����8k���h����t��ƤY��)R��i\h�����,v�L10m�����V�Um��3 �X..�q��X(�1+D�1(�֕�.
#l�30Ȩ����"�Ĵb��\�űV��R��b�U
ˉ����.��*چ"��.[1�JȎ1���L�Q�6�Jդ[l�AZ��]n�Ckk���R�壙n8�\�-��q�j�\SR�`ԩQ��R���*���B��E�Wp��ЩZ&3,�1�VҋbF���e\j[J���Mq�J�5UB��V#P�R��+73+����V��R*Z
�E�JU����.E�2ٻ����
��Xe��S��JVŊ�m��Z��j��L�Z҅�9mxy�V��o�5���q#M%O��Ӗ*��l�V�p"nݢ��w<�VvoL�1G1trbΪ��w�G��L�1�D���m��1__7)�m�z�yk<���L*�@��~�6K�r̳��M)�5"ƭ#�e�0�զ�����~B,n�E
�����|�6�Z|u^)`��[��W���@���2(����K�y8��r�{U�񞷲R4���L�PԡQq4�h�;����y��FM�c;=	�T�v�(W���A�кq�黱Kmv���=��:i�"�Y��@�*�FӾ�D���\�E�;W6�غ�a�EY���"�!i�U��DƎv�����YӠW�e���LY�sx4WD����sk&�L�M��d�
[n�lO�r�����¶"䢭�	<4�BS�u`d[��2.Z�Tw\t���Esd^S
2����ךʆ[Ϻh+=��
ccGx��AZ2������
�S�B8ӟ�F�J֦�P4���~�y��e,��t��Y�8⪘1c�bY�1����UwL_+����ن��x���jd���B�eFٻ`P�����{�v�T��6�<_fF�]l�:�#o���-]T�<�㠁>g�u�O��^��,Dҹx2ԟ�c&�t��Rf��WC�pV^L�7>.*+�r��V5��y椝X[v��{F�[�Y)d��
�3K"���D�f�̓���7vsݫP�u��#؜*Wll^W^��b��a2�}E�.��;�R􁊆�1����j�BfmK3s�,�:Ȥ�.P�J�P�A��y���;9��L�f�x�&��ל���iU�XM.c�)G���'d���׈�u �7�u��G3�5�b�,�vŋ�Џjss��5�wb� �S���@�K��y����"��p��_9��Ts�
�{�n��0����0��<a��g�4��0��r��0q�������U  �Y�<(��3[�[Ϭ���Ʉ��Ku02�K��nȋ�:�F�!�M][d�Y��u�9�.�Y�PE�:��t�Xz�ބY�Es��aK�?W;�o�l�owwS�e�މ�X��ꆸ�kWOE�+�k��(޺�&�p�|�-i��>�q֠�=���S
h�����(� 9,�����O�b��l���̮�,4��d�t�1IT��w�1K�oBD�F^sUOV��O{���ؑ���ϡGY���J�8>��p��=;L�-@SD���#fy�O���7_�i����|_t�;�5%�����s��t֡u�[v�:*�� BM���2��S��a���td���z��E�\���vJ}�v����k�����tZ���l;fVȄ�8_Rp(�9�G�rqP���{+��������iw������S�+�3��ҮiZ�I��k�Py4QCX��a-
�P�q.�9:V���h�+��YP���+PW�P^�܃O�r[T�{+cJ�P_ß#���M��v\�ێ��%��+�5��G��7�ʫ�їO�s�l�BN�f��/�h	�<����t���P�Q�Z<m\��j����+N�B�U��mt�
,V�cj Y^�,�
�
2�C�?#�Y:�#�Kf��zk�Nk�lw���s���=*�Ĳ��Ue����B�k��`�THV���u�X�x������]��+��D�t�Y	�1'�WT����0���9��r���Yx0Q����Ry$���?:<�ޛ��F=�?��B<�; �n�GDl�c�@v��u&��՘�w�h�5�0���1EY�4Ī0��Ft7��?m����@���Δ��PTe��7v{\�F@s�9�5�hY8:��|kt,��YC��2�O;.bx�j�ήj�<�ٕ�b��������T�����g�����U�U��[���>�p�v��n�)��*����f�.7�w�{�O=7s�ȟ-�ܭ��sHܳ�KuռV*������ǚ|�\W����n^VF�NnU��In�4�9]F�-��ݑB��.��<���f~qG%�d��-]9-��{�<��s�(�B��b��2A
�MA&r�}�Y���Ow�*�)�؏�ƫ��m#����<jXCU�o��O�'��T~s�L���]���$0���t��u�T܄�n]��e����Үk��m��٘�ړ�����G���_Kdh�8��ϒ�«�M��W5P|>u҆���:��%gge9U��.iGH��d�3ϩ��嬦���p/S�/-
8Z5݊tVu���g�ަ���֌�y�-2���=,�B�=IU3�S��i�;���.���ڟ`�+���mir%��7}�-z���x�f��+\<�I�GT+"Z���-N�Oa���*"�Ѷw����K��ځfu����6��<�ݞP�WsGI�)@)�f���T@�;��re����㰱Wh��8W�(Bwz9�c�e����P�}e�O>��L;m�!Ĉ�[ oL���kX��״�����c���t�f���[S��W�����q=��YU�	<�r5c�zq�@��[3qX+�G`��WT)�������C)�=�"8�9��P:��(C*�PCܠ��T�C>����̓D!�G��5�pӽ6*���׻6Ī1W���7�%qNgκ �ɊA�MsGEp��֩�P�C�s���H�P�%Lg�p+&�ۖ%_��;C�r
����J^Me~��r	��s�	o��͖��P��:ݫǏ�2��L�s]�q���a�ճ�����u����?^�����\�ٹ���Nљ��K��MʣF�f��U�V�'�mCl��:t�t�LJt3�@&�6�Q�H�q��վG��#L������@���7�Z=y>_q�Z뫐׌�<����t9%�^osy+4x��|:`nS��{N����*�m�si�tKdp����0��v�m����,���%���O��ǫMC����N;_�7U��U�U��"!V�tMV�5e�
Ί32�����4Cd�h�mw(��OK7t@�4��D�ه��׫��Ku�t�Y���kF�j�N�o��Ӳ�G�g��@j���P�<D�6<e�_l�w\P�Va����:��iwk����|�QG�����e����P�8S�� >����wݵ!�Pv'�s�^��IV9e�3�z��	�jQ8^Z�֜Zyf��}�X;m��w5��!������'�{o]�f;V?v��*̓�S�)~��w���
��jw�f��J�w&� :�C;������A�{���4t%�^Q{-�ˮ_Koc;�Q�:飦��eP���w�V�[\iv�Ko*';���n��rTP��u����M�2�A��A�^t�Tϲ�#I�&���s�q����~���ӿӐx-��[�����0K?OO
m{���Yp����z�l~f'��f���6��;�ZŐ~��3&t��^��-�6�.�.�(,��Նv�v"T�����C�un[��˪�<7;Ɛ^�6R9��t�7��Y�I˵o�ҥ|���0���޽�r����a3Ӏ�x�i�̡]0�z�w�5;%�>��e���X۬<��1���]Hn�}$��=PJl�WUW���N�͡Fi5�t���Sb�GCϩ���!���8�{	�PԂ��b5���Y���������Pt"Ǒi�d�OtءLeFٶv�d`�G>�,�UL���:����aצN��v�]Q/	�)x>��h�(<J�x3I�fd�Z�{Xt����^e-̖�'��I��_M�q����ϗU0s+�0:��CZ��N[�(�a����������|�y���,G����
��ǽ�P2·� ���<�6�dL�p�l���mλv�Z�茹eMu�ʲ^.q�٘B}����}�9	x�F7�	�lּv"��;�S1�y���+<dh�y�ޢ��]�� o:[�K� M���]_T���R���ݨ��͝sBwVL9�&���~��uq���z6֜_<�a@;6����z~ɪ��y��u;��,ׯ7mC\_T���V#0�3�7��RCWD��WO�m)^��w���Dmϳ�m�G-�僣� �;���L�˽�Ȯ��EVp#����a]ty7��`I�.=�H��Q��N�6ԃ�̱���>�ɭ�=��fe��a������Z^���XP��e1s�b�՘�[^
]�_Э��u��4���/A�n�Ae,}6��J"'�0ئ{O�T�lPYY�O���؅�?=�)ݪL��p�EVv��z�ن�(I�ѻ;��Z�R�6〻�*�:$j�A�u��od����ƍ�gtwΞ�:��o����|��W�u��j�嚋���~�	An(��}Gr�+�8ONŎ�wG&Sb��b7#��7o�/9n;�MZk�y�1��;�����UL'���娸K�2]��&��k�����3n^��̓�QUB{Π��NA�� ,}�o�h	��<�Gu��wj��ݳy��G�W���5�TQ�N,�t��S��(Yb��7���L��|�f�Q�柑է���3�B+[NU�l�G!\���׆iN8�ON�8�~xeA�iMnϡe5���,��4,�R�3.�0���]�j2X�ɕ��t6>a@��p��9)O �����U	儷&�FM����)�V���ݺ�X^�4�5sv��Ѧ'4ݱe&�8G	k/�1�p�����2�#ʧ� N59��у�Xs�̀����#p���0���1G���*�6�vQ�6�e����]S	�5uu��1��u���E��X��'���e˭�188<���a[=v��w�&9	�ܵ�����x��.�g&9�{wyj��s�*GWftި0���n��ܹ�mc�zz�W�Ǵ�8'=R�<y;����XK���<%;�g��^��/e.�e���u�����{��ayl�7�{{sV��y�lB=��������G)�'��Vz��}�s�x�@NI�!����x��mlј��s��J��1;�4}�d�A��s���%���B��m\t�
�^,R��ٜ.�k�t +^4�^R�6�ʃ���C0������e�~qGgβX��r!�,d��m�.�!zNsWuGI� Wg�#����O<^R�«�P�7�_2W�M�P'*Ah��M��LT�6����FK=���<���Q�lw�s� ;6ڍE��s��WP���V��h��+T���W�.BA�h��#�IU3�S��i�~��KY��D6���J�ky�T�§3�Nt��vDt�ǜ���+��� B%K��=�47T+"��C)�i�ǐ�v���hF�# ����V����r�[KN6��u��<U��n�g�0�V��"@vɅ�	j��/�w��Kl9=Q����D�瑚e-�؟��5�p�z��ןB�R�\$�y��e{f`P�y2�v|d��V~�Bx"4~S�mAb�C�
��#5�$��,�m~�{����k���m�Z*�֋p��U��{�����Ck��*���e��<���x��}��*��|�X$<��U�9�٤9*Ѝ.��cgr�_pKfΫ�<����9}�e.�}L��_�f���j3
���[S��^��#��zlW���MK�Z��g|�\�+I۾�(p��������D�yf�e�&�K�r2Ǟ��d�
k�H�SS��!��mȘ������z���v���r�`�Otت�3��d'�!�^�4�\S���\Ҭ�;Ӄzwo"3����=��4D�@~���'~=�4�=9%'�9L��Q��Z�iȳmG��uR�l��ǳe��ݻ�v�G�v�=�c��/���|^#�����oCŧ�ѭ$�,�)kvu�j�k���	B�d4o8�y}x��԰s����	��n�jx�,�1F��s�1�z��M��=���\ �6��	mw(��OO�� _�z��f<7(^�(b:�C�s.W-5�^y��m��l�k��3gQ��@~~]눖��A�כ���.ؠ���@�hp��֨9Y�vl�y:��ʌ3���عeLb���8:������*�;�U��Ƶ��ǕW8�"�v+�⺜�����B��#�G�D�yjw�v�����#��K��{�`]ᜭ�k@k�;��v6�yҟdG����wE�;)zs���ͩ�բ�Aen�z(���)b�o�^�W8{}�{B(W�B�X���}����,�������h����V�c����4T([��j��F��T�OX��lfI�\j�u��ku�妵,ӵp>�N���{�t�U-y*���~��v��d���K�jw�f��Ji���7i��ۻ{.���yt�Bw]�Q˞�/e���_Km{���OH�~�K�0*D�J�`�����6'�O{��j��	F�Wd-8����:8Q�*[;��t��+�yƃ^s�$6�Mᬺ�i�
i`�& �~�-N�-4ӕy��cj8f[(�b<�=(Qˇ�Σ)� ԓ^��z���K�x���y��~.&�#��M=.w��k�eC)m��3ea�o��� :(B7���*:��3��*l�����{� \�)�U�iG�_k2K�Oiۼ��ܦ�K繜��Q���8~<��t�̦!A�M���d�})�d��"ٌ��7`���2����e��ۮ]���g|��%>�t�0[]R�<s EԽ��p������D�\�-5�N�I�ˎ�ɵ-]b�3�Q[J�f���>Z���,2�0��Ga�/ڭq�l�x�f�g9Q׫#��Ovܗ1�9gb}���lB=��ys��,v wb� ��=.�ͧ7�Ur���p�Ec�������98P�	Y���5]�g-]�K�K_f�wX8D�X*r=��&��sy1��s�_u��%խ�'�-�K�f�~"�nL�,�>�0q�!��I�:�a�wq]!J`5�.フ�����*��y�޼�(Cqj���|���Z����t�G��{�c�T�S፧�+ݦ���e���8�}�c�H�7���v��8wǻz�\21"s��+~ͥ�d�Q�Ϭ �z������ާ[QփrM8�jf��z���k���Wyܳ�YV�u*��$��)��J!�(+c������z#P��Y�N�����1���Q�޽N>��)i=��>����쩗�M�������#���nRK�볅��I�Ǖ��Q鏷�mj�����n�*�-Nܖ�Dhv��L�WG����]OP\!�_Iwl
U�og4�U�Ϟ��
�#S#�m�}.��鯁>�R/�q�{�w*!W��/t\t�<6���9�,]�[�˖��w�v��&������k([l�È]�y4���WPrЭgw[�����IJĲ�K�6J���j��T���b$+~�YA�C��3��歵
/�f���Ya�c�f���}�HoR��Ai�۩��2��}�յ;[4_a�� �
R]n��l�[��7Vu�0G+�>��h'f����U]�vo���ڜ9��Ʃ�:D���:����*�u���� Wj����T���ؗU�#Xj��|������˹V��r�o0��Dx�܇rS��T,��O-����+tp��g��(#H�,��&�u,VL��G��-�h�4m-t��Ԭ��`ͮZ2�h���Qv�XNZ��z'�2��@t�M��1K6��-ʼ�`�/1|.R{٪���TGv�pjk��v��5�Qp+~�(F�+�7�c�Ӯ�g:�-��nNoA�-�JP�k�_p��=��<�*�=�����L
U�<o��/^����J�Wb{�~���������m3ǔ�#8��f����\�b�8Ob^�	��~��pĮ����r�mXA=1�y��E�Q*�L�>��N��T�%fM�)��#	rJ7�kM�(��
UqR� �y�9��� Gj��nQm�ٲjQ�%�6��PC�w����ԡ%��z�r}V�<�Ι7��&��F.j�NW3m�z�<vt˾�p9nA���f'_q����n�z�|e��Į&/��YI����s����\Nt`�V�f�s� � �WB�,�]��B��X�x��ٰܹ㨅��cb�tXJ��t<�
����4�hy��=���2�z������D����e��ò�O���G���t�\�]�$��ڕ�au�rny�NR�0����)n�{��=.uV
��kr�����<�*D�Y���u��Ƙ�3	%K��O`�.{�Ѕ��;#�{1�|[|K�<X8�`9q�3��n旦��J%�OV�\��������S��h�j)Q�a�%#ZҘ�1U���P��B��j+o�QW܆8�ˎe1r���+kVYcjTk
��hѬ`��)A[�9B�ƫ�b,���ڣ+L�*�R�9�e,���Զ�S���[��ws �3
:�`�kaZ1f�)u�:��QLJe��W�q��V�j��PQr���ͩEZ[cm1(�fe��j��Q*1��m�" �K
�q\qws+Tm�4�)���U57R�[b�\qh��dT�4lX���Thԩ`�""�D30�ۉ�"���b����a��R�n6��c�Ѭ-,h���X�)�T�ʨ��Vܵ��n����\�e-,W��-FjT�u-a�b�h֚�Smԣ�i[JC�%J�6ª����QamFTTTih��Y�eq1�EAFe >�{m�S+��31�8#���<����,��#d�"�G:��@���Tc��L�O6�V�\�%�3$���� 㳽�"��!5$|����wy�l�]F��*�x��.1�0��v!��x�r���2 K�<�����1���	���$N��Q/O�5�b����Ǜ(qw�����n�/H�Z_'�Y�Q1W}V��NI�2y����sBV�;�ئ��埲x]5�V�zf}i���OR!�B�u�"�qi5<Ù�#*݅ylv��d�+�e���YH9G<���J�(Us��O�_jv��jz{)���8+��NE�| fà��v\��e{:�����?=�;�d���J�[�V]�?>^V�����q���s��[!�-�!�l �ъ{Z�+͈>����:��ux&x�&^�mvht�E��}��)t�=�}�-N�7�6;���D�m��w-�T��[�vl��֗�*���f�T�j�[5SG�g,�#���ǯF�ԦX[S֧���.z�vJ}�v��Y\w^e��K��ӱ��R�+s#�O6�VT�gۉG-�����5k4C��g�8�<���R;�O#�gY���ʷi�y1}<�,���g��Z[�yF��a�OKu��(W���2o`���K_�س<�/-��/��b���g�ް^����v���eǛ��`����y4{�ol7И!ڋ�����}��Ab=5�VMO;�Gt}o�c#�9cCO����׸�1���6_W�T�>�,��-e�ׇ-l�le��!�p�*�Ce�S�&/�;V����0�s
�F�;���ï-I��i�T��Wq�Sr��8KT� �}O����++�!�^Y��a���6>aB|������9,��
k���U	����s�ُ��#�M=*��Q���D�K�t�s0vTc8?m��"��O���ݲ ������;�`�suV�b��# q��s�#Q�hp+��[E�QV{1*��,������x�f\f����qT]gf��
�8͛Q�^Z6:'����Gd��k���P��me��7tZ�!_����[�歗6zJvT�������N�w������G)�'�qg����{9���c͜�2o:^��^�nT�@�*��x����<���x�2۶Ɍ�=t����x�(>��i��r�W�F���|TY�n�C[#@}xDΨ�%�!9��W\P�Wfs	�$�g���Ʃ�5C���l��h����u&Z����� \b��W�O�T�l+z���r#?(.�Uu��/�~^yW\d�?E�8��U(�g��{�)��-��.|��������-���Xs�+���zu�se٬��FF���H��y�c	н�(h����-�W�d�j��W\�<��yIr�ouw�;d!�~��J�i�CG���Q��t�v��cd[1�	K�k���.�*�϶uU�;dm���ձJ`�k��SG��ښwx�i>���u�Y���贩���D�~����N��~���×�I���=�S�gA��yß�_�{"6��3�݆�f]r�Uy� D�t�D���
ȣ:P�V!w�G:;#��T>nb��n�W�H�j���7���}�;-�6��l�掓>)@)�f��l�T@����t^Wt⼻�=2_��K]��ӠR~�}� \4��2�v��:�,y��f'�R�<Md��?h��u w��iy�Al��0�/Ϙe�>U���OJ���OV�쨻#qz�����󑹏M��/�d[K^�ݗĭRϹ<煃��8#|��i�9�۩��.Зޗ� sO\�"S�(Ch�z� ���M��g��ͳ��c�c=�i�1�ǆt�m��[U�*���9�[ otÈN��k>�L�����S�Ժ0ex*[+^�K>UꖞI`֡���}�v�c��i�G�@��@��h8g�B�h�V�1�uc��=��L95�$��d�u���E��x'D6�Pй��ϙ��w!0�_�Q0��y牖�k�G���+B��zһ�ugT�+�\�L�p�W$7�ޢz��8�6=�i��+�YA�*M4kR[�Y�܄,y�� �����q�a�Հ̯%O�b�xS�^!�����x1��X}6�c��H�p�<H�m�(E��:�kJ^���$��:P���N�:;���z��f�kUӅ��T,2؟x���6f8N��DU��z��1̭y���\>tY��F��*1ls�E��ϝ-�m桕K�k=�r�:8N��,װ��>쨸<�h��Q���G"{�8��2軣\��2β�f����kz�y���|	�[j���x�M�hDX�є�_h^��
���j��*I�C��E��"�G�D�y�{�ikN-<�q׆mtTF�Z8�bUn���P"��[�k��*�����6u��od�i���ވ"n�*.&���W�h��{�j�l���a��q�-��F�t=
9s�(��ȯ.����DB:洧���2��
���6s("��T��L�S�X�:؞Ev:�z̪�n��+�v�����UZ�8�(b���x_����ÚR�Z���;���d�8�t��qС���xChܶ';#K,���2��uY�F]<s���"��N�X���[L'ާ����얼�eC-��;ea�y=�N���_]���)�o�}y7?
c�

���$e���s�wy
lUH�yf��ז��e�׳|��9#�C0���pҦ�r�v�v�|t�S~�&�T�Ø�U [����C7�MN�l,�/tl���5�!�(���YM^�o���uY�C�)-�U��qg�5	N���0��3sz����qҦPb#�;��
�Ǳ���5���WK���B2���U��Y��s	�>����k���!A�^�g�d�}*�@�f��B�ʍ�o�o#��d��7uqۻx��N�w(��q�'��U1hU�}gZG��=s X|l����kOe�ff=�o�?<�}�P�mtOm��#��s��ĺ���U�Xq�����p��y��<�m׎s]�y�m�l�]�saY���B�lBw���7����m�P���5�6?S�Ş�ƽ��[���}($��$������"���%G�q؇B�]�e���K3�5�����mI���;�6���Va��2P8�4�2�b��UDa�YC���VOSt�/��:�$�"mn����DV�kw�s�sB[��������'�׮"��zބY����ɝ�]Z�s��U�N��n�1�s'��a-����چ��맢ܨ>Y�~qF��H�8xN]0ކ����Ef��\o�]n��9W����x=2��*��(gS6l�,�C�9��'l����C�g3f��n	�.���J���3���>և�J���u���?>���`�γ73_:u�XC��鵤�ؿм]ײ^f�A ����Y���GS\�i�]��o'Hupt!�~��x_��yl�CޗL(=;,\+�{7+�S����4�*�p�q�.�!1��:��^.}�v��vy�t�?�,�PQ��E�Zd2�K�{�t���pSJ��ƟU���G�7Υ������3N�7�6;��H���׭]!���n�\�����7�&e�w�FiX@+
�'�נ#�J��K�9E�\���S�]�k����ٗ�۵5��9�Y�?OO
;p��5�I�y0*Y�M4��:G[�T
����{nV���bs��9���s�{�]�Uu2�n��jy��)�Y=3�� m*t����>��yO���WVF�;���ï-I��i�T�%�G<�����ϭ��,�z�7��{��^��S��N��(s>��
2�[݃ã���	���8y�A���,C�uO=00T���P�pI75#m�k��
_���F�;�ix뗒q�L���l��)�'�; ޞB�"�#�v�^��Vt`�|��p�Ӝ�<��t�Is�EY�4J���3��uQ9i�׆Sӛ�i�H�Y oy�!��9~�� �Q���������Ւ������Zq���5}ͭ���5�&ݻu���߇c#P}.踿���r��'�늛fG�f�$�v9�F��*(���dL6��{�='�=B7���l��'�|���#�ԛ��5��'��%E�n�F.��.�����9��t641k�)\h̬5"f�fi�ةN��8l>�ރb,Հ��F>O/QF����]������!9�0�Ҧ2aW�m-��
��<����n��:[D�!��q��x��T[�c��$N�=p�B�����"RV"7�m�8ǝ����:�}xDΨ�%�!9�ǑPoˮ(Kr�3�T�n�}\���Ӝl��Whef�w��Xі���T޺��6��~ U� �j+��~»^B��\��u�#�4ݵZٹ��9�\r�T��ШjS��-N��>��j3��/9��j}E��d���&Ջ�yʻz���7,��M�p�g�wN�Ń�45%T�4�iڏ>�`���	V������5<s��`ק�3�[s��/�k� �gΪO[3@CuB�(Δ2z�.�do�7��19��_V�枊�΄���~���}�;-�G`��-���d��>Ā���)u����̺}n�Oo����?q�09ձ��7�����nvʖVI��vq�{�K=Dj��w�;��]�0(O�+�%�����?���	|��(`䫤���qjO=%�)Iuc1�n��;�<k@���nF�=7K�����&���5�.0ә��q�Ϗ=��2o(I��/;�+���i��͔�<�Ml)�{:�-I�̮gO��J��5��=86�8�k�
KEL�n�C�юg<�rkY�hD�Fu�%�=g�B��|�y�p���\D��{{�WP�aB�б	����fi|b}O1zף�6Z������Y3{�	��������P8�>6Qʹ�.{����ת:Ī0�|a��<�{�4��79&�e�n��ڍ��Þe��uI�Q�K�i�o�`�4қsi?a΍�uY*Z�n^�-˦����#]��8�yg��#� 1�Qā���e��XWm7���4����sb���9��|
'#EƼ�7`���8�yft�9�rXe�L8����&d�=��>�p�P|�Y��VYS]F�O���-�f8i%t����Ɠ�H5�g'��E��Y��g��݀S�܆�9늹er�F�8��m[=<(��+6<j�Ԝ�_n6����6DҤ�޺��,���ӹD�r&z.[��Ql +�=�0�mP���8�)��-��M���GwFG�^�e���Wfg�z� T5(�/4�|�6�Zt^A��U���#Y<�nCn���qL�z��wfSu��ҫ�9�&���Fw�B��z[:�Os��3G<N��lRl���Q��;��� ^��aG.ze�غ���ocD#,���7*�zB�A/7-o�#ŋQ쾓/e��k(�FhMt��\�]G}-yS��]�|�O<�L@��J�ݖ�画�I�ge�
�Z�Q�;�N��	o�ֶ�wۆ��7yӀ�r��X���Ż �K=n�SSP��ԓ8H{�(we ���ߥ#6���Th=@v�*0%���L���ެ�	F�Xo[!���8O:�����8�x���5��.�X�{h~u���<4�GvH��e����_��Q�quѢ§�zݛ�&�f���ؖ�ܫ�z��� �Se�'�}c�F�
��UL*]qy,�:��e,�Ѻr�i�D譇1��i��ܓF	W=<r���H`���L@��d)�T#�査_Z�|�.�F^��m�y��^��;ϱ�e��閤㊖��"TB�����`�W�2��M�u6�
W�;�ԅ�@Ι=��̌.��,S�ǔ��R��La��& �>�+I<Gn�s|�n��D�uv����Ns_���߻r&e��9^`P�m~'�6�ƙc�7�|ϯ�l�uSҫ���uz��E[�T������l�*)�n�]�sg��Kd!b6��`� oa؁�i�/L^5�n���R�\�̒&c6A; ��oMw,��u�,�%���t+��x�ݱ�9�ɡD���t��<�D �K��vه���?�<�F_�eq.b������,�#���?��ǫZO�3��?3�V2�Vv�A�en>?��~�i�@��O
�e`�F˱���q�un�鬎�DL�2IZ�@gypm�U{͝ggLQ��+5ȍ�|�������Cv'�p�v����w+�!r§+�/��k���0K\r�ƹ�îؑ~�w9f��g�MqS����"��!�D^2�+*�j��O�t��a�����B�z�k���z-<��@?!t�|n����y�+�X�p>��}=dsu?I���ruϲT?�%�W��̶��Ү�,!�����I������csmS�&��e�]0�I�3�K��Ή��x�(�=M�����; �ˋ����ƭٹ��gyl�?=v��Z��jJ��h��G����t�b��Qۊ�BxƼ���Ө�E�ǎ�C�'f�r�~;M� B�� ��^��u*�gS�(�<ӕ��v3�9͂b�ín��G,��feO
c��/�Y�(e4l��|S@Q�<�9�.��>����J3r�`�=�y���ŏ�k�������9CZݝ"/}�ga��'v<p�����[�炇���O���F,��E{y����z=,�;��YXcÛ�{�\��6��OXx^e3�]�,]��3�,Y��G�]+;����:���@I�@��$�$��BO� II)HBI�$�$��@���HBI�$�$�� II?��$!$�yHBI��	!	'�	!	% II9BO� II?�HBI�d	!	'��$�$�ā$!$��	!	'd	!	'�����)����Q j���9,����������0�m����$JJ��I
H���QUAU%$U
��P�D(J�"�JRT�"�H�JH�J�J�B���&�I�U"�)�sr�EP	u�!IR�$�QIl���E"�I
T�%UB	I��y
TKp �kAP�mF $0���RM���� ��PE@�1 �B��
�B�!� �0�� �� �n�� ��n��V�	b4	s� PW  �v�l��e(1������
i�lZ��V�+`4�R�4Y�fKl�5Q� mt$�lJ����([D6�֍���ɦ�mQR���ASYV����SP
�[aT-� �aA�64�%f�-�������kR�R�JٶQU���LJɠ̵$V�U �6d��V� .젡�YJ���h����-2��i�3�j�Md���@���dj�[`�	*
' �P �+0Z0QkD�E l͆R�QDZȐY��2�ʀ@ � �(�
� �6�i���j�ka���	��M��� 3�`Z@B4
�b�eFU����ԠmH���*�� )A���**34�l�6ʕ�@̤HA�o�    ���JH�� ��  E=�	)JTd�&C F&�F*x(ѠڃF� �  S��*SU z�@  i�� D�'��dɐ#)��f�A�O5 �I	��J��р   +`Jl3��UbE�'*X+,D	֥�F"Lr�"�/���u�����Aj�="���
 P'o�������⡈}�� �C
6��O�RB�L�����E/�����j�ו8qق�(�Y\9P�ZY��9D��S8�1�K$�	���VO�~�9N����N���f��y�-M����DQ�`�b&��.F�Y�Π�X�⺽ʼ�"f4�V��M����f�3FE01�V��]͡��U"��Z(D�X��uBG '���`k��gE䈘Z6�&���(jb�QVe�����YN�c:���ԙTY�\��"$��c�@���on�#),1l�Tn�CO���̸CV��"pg���W����܍cIɷ����^nf����2@[���֜�5 �2*��v"rl��iM�K�p�V�cR��(jѮ���*MV^ڙIˎ��h��PN��n�kBB*Xݵj��%DEM���;��
��ѡ9�vr^%������7P�GAt6�ll[o����63uڹ�*:eR�K+���;��$��$%��;:�J��r��1b�E��Y�,�9wyNa�I7[����t��F��[c]Ŭ`�O-�z�Lt!wNE4U	��&���R����Rm�;��G�v0���J�����j���Q/j'MQŔ�)�7o7`��Q������2�)�Թ���.5��Kk��۽���#A�ҭZ�K+Yu4fmi�0!��	����%�����[T�M$C7nҼ7jJ�ݐK��l.<�Y�O&�/h��GBG�ih�c�ݽ֎qSܷrV��V���مѳb`WG$Z�xN�N�]nJ�n�aj
�*�V˃-ܩ�d��� �h sd�r�(��ҵ�8D���STա���DXm AT���Q2�1E���S�t�0V8JЊf��),��]���-)³ө`@$.���7U���r�j���k۽i�l�i�I�y��N���ǥ`��plB^��])��5���RwMTx$&C(D�u���=Y�(VVK�4�L�f�Q�Z�yR�EL;%��Cz�7����Y��2����	�����^����֠8�H[�͙KKĵ�mt��ڥie�7ËK�RA��ݛ�oH�^��v���c�˹�,�޽[aŒ��<��׮�-)��،���kjd�!�^7f�c�ȠV�)ݱ�ʫ�v*=��yzeS.�ӧZ6�ƛL-Z�4�����I�ME�I�J�����	6�MX����5fAZ*!f���f��ؚ&�27.R?f�M��VY2��f\��(ѐ�Fֳ�o[W�R!u^-�/f�"���Z7��m�[��û&�q8���wY����[w�!���n�����4���Y�J�}j,@���4��w�e���0�z���I4�ZZ�]\��ce����'J����2��5�.��.e�&�r�������Y6�T����$%ټg�NM��`{tm��K��Y�Su�ܢ"�'X�%Ϭi�FCom+�6��+3CN��)��= ݓ$�(�&m�3`�lV�7��mJLdWWBL�I�&�����&���ЛE�J�[Bmօ ���Wk`�ɹw��5�6K"�͵rj&Uv�cPz�u�1h��J�H[I��(�K�w��=1�� �Am;�����,��6m� r6Y�%�ѭ���5b�ڸC۱
x��˲k4�u%�[q���wXw)Gtb:M�d4.�pP�T�GM��*jGA�'Drܥ�k&c�n����,�Zhǅ
�{s�ޜo��VYz�aU�dSU�	��5�0�ӏ$
ڗ1�FBplP���clmjrLT�FPc�F,��k��^��÷0�	�	6�^^`�)�ٷw�*S&P��ȋ���2��6I	YU)�m閮\�k�nm��*�<qc�Y�kٰ�j�5enF�t5!0e�G�*)�ފ	�Tec�������Z� e��I�tE�Foi�5:w��5��,mcȡ�4���!YQC�Ub��rYc�
�����7
:�6�j��fݧ{����H�m7ZU�2�x���Fd}�+�R�㷅�Wm�i�+=�^j�L/e[bn�H�nh�̘��ĺX��\�+@=P�(�_^832�1f��>+�`@�������/]lt��q���v�K$�H����V5���W�:r��ݓId��lU
�m��iت��Ӓ�#p3wB��N�9q�����j�L�5
/Àa�AM�g2�Q�3b-+p)OC)a�Z�ֈ�U%ۗ��]���������1PܠT���2��b��)���R��Oc�i�Y�]��tӵ��#3D문�㱅�������Ԭ��H�l5IRܼ���z_W"��K�z#8[*���J�j01l�V��&�X��ɫ�.ڵ$���%SyOv�ʫ�5�`�R�+J_CC���km�!w�30��=��iZ�`)���34�I��*T�c ��-�"�>�јE���dͧ �$�w����[Ո�!�]9@��vP��mO(K��+�T��K(3�!�n�Bƈ1���G-lh��h��ap�K)PĮ����ZoT���&^�Z�F��ءw��1VjcZ���yz���A�6��3`�*c�nX7V�Ў�r���ma��"�庢ofM�%�D��s��)R7���bB��H�UG%Z��5�
�Ƚ��3[����D՝sU&�)��B���-�e�dL��b�K`z�p�q��������h�Km[�)�RC*��Y�@�#��2����9Z+i�+�;�W��w��Zĕgj�ͬ@��P���P�D���pXٔ�
[1V�E�T��w@�V�J[D:�oZ�D�e��bۭ�Qf�M��I�,�xii�B�^;!��a���Cv��a
j�J��۔�[��/&��a��A����vu��!�ِ��7q	2�v't��b��k˅n*�(��KuksrlZl�Y��Su����fů�ŵ�����V�0Й��f���0K�r���� uf��I�����B�ʡ�s�S{$�Q����u���W��]�3[5tKU�ȯ�s4K.ۖ�Q�1��;������%��J�6�	��,\�ѳC�l#s*�	�i9��n���&ڃD��^�x���Z�����@������f:��J�P��!od��%�.6[@T�ۢ�I/�5�����F�m"dU���ϲ��U[5�e�,o��˩���X�wf��eX8��Df�h�ɿYE�L
B���G0�Y�M�T�7GL݆i׵2R�T1��za�V(�)�U��ڔ��]�Z��7�]����V��0��^lp%%�9�q,��ZLq�Q�(�u��B����s ڃvԭ�̺�t1CS��P�2�9�� ��-�-�v�2�K���cn(hGz�L7wC�[6hJ�z�tsK�����j��&ؤ���Z��$;�k���� �$��-���e�mfksL4��Gw�V�cMk�e�V���4�6�Ul%�.��h��2\r�7���Ytvƫ�q:�W$�[�� �k�⳴	K1`ol��7������n�c�;��$TX�b
e��ه7f�ǆ5i��#B�vcŃk����(���X�8��s3e0~W)\��f�وh8Ժ,h�C/UȲ�&D�Jw���婡v�5�c�X�)���R���,�k.���p;��ܕ4����i��[�*,,3r�C�_c��ֻ��M*��r�Y��O^�`x�h�#�H�2��> ��uaD��W�w�Jhvh�fs�O��)��r�)�Q��*ukN�8N��h��cX���)i`;V^�i|�^ͪx�n��ԏ����WV�^(튴�D͈�j}�y�����pP�-��Y��l5En�h��!����!C�*��b���P2��iM9f����ޫ�ce���ꯪ�3���!�'LtP�օ�(l����ɳaq�T\~�����I�҂I0 F �JJ	$� "M���� � �$���I0 F �JJ	$� "I)($� ` �$���L �$���I0 F �JJ	$�wdP�gu���Y�\�eJɳ�L��}Fv��"�=���:b͹0�֨$%Y�Nu;"�u/�w2q����u�$�͚��[��RِѼ���-tS�]��^r��n�x�p����P��N�Eb�r�
���0��dN�<dVY�9Tx�}$$�J(e0ʙY���K�{.��ߜ�k��� ��������dg{��$-��N�;�[����c{Uw3ـ��V��)��c7��k���,wmp�zdKxe��d{f�Bo*�/��pf�3��N�����.٪�H�7]x�!坲j=�M;8DB���_�=@�\�z�P��� ;o�}f+�`�����ɩ�Z����7����8[����yQ�6��|�Yr��Umήcz�(��Y����0p���/�B/�X�Fې�S��6��y�i��g<|MT4i��_��e�ͽ���k7�S�OC,�9� �Y.��˗{��e)e�(@CW�|N&�4����ڡK�EB�����9�톻e��,'7I�҄�*��F��H�c��ޒ�,T���缛.�r�>.�_�ٙ��o;��x8������_B)ߔ�̦f�|�b��G�����C�����ɔ�abml��d�`)V�n��oݑ��JI���wbr��P7�Js`�.�,�������*�e}�rv(�Ѵ�Va���Ȳ�s�`�`��ܑۗF����B+�ـ�`ݙ{�h�}	��ռDഘ;D���uq�s��᳊�m�˂�̬��NL�q<9!L�d`_��n���Ј�Y��r�ڎ��Uَ�p�����g�n侑z�={W��$VɎ�Ss���Hgv��6���DU�&�j��*�� �ֲ�뽍G$++����/��ElZ��`��m,B�T��v���uқ���8��5G8�����4�|DՎ�*@�7/h�Wζ�}2���w_.�w6��2�1�����ַ�{+�h]<�۩4�VA.��t�%�]�q����Q��y023rm/�H��ٰ*�ۖ��wY�7�_[E(ʃ15�Gzw7
]>فr�"�ܤ ��q$qv�S������ݺ��L��2���öIm)vU]���9͑��Q*�"32�A]�n�,K�Ӕ��u|�g(B�J�i��:�Hq��k�VТ;m�k������vu�����4S�rۺ-LU-;�G;���47lG��j�Y#*�B�\+"��O����u�]�z�e�+K�!��llƃX�:X��H�N�.���q�]T���'��'~S.?5X�>s9�0�B�������B���Y�L�&	;W;�雚	I]W��I�hnY6����EA�금�u��r�h��T��k�ׯ��9l�12�[ʮ,qz4�R�1CWb��h�:��n��х��*s��D�GSf3��n��v�ĺV��Y����lۖ��-y����a��4ܷx"�ȆX��nu��F6�O��c��J���8��.;;�t�ivTe�*GKhƸ�J#�e��z��c]d-�(޸R�UkF�@�j�i�zy�]֊����Çe��%OTNmL)�O���y���N�(
v�辮��vǼ����N�����i�T��{Z��]�F���Cns���q��q���+��4�Sk!��AoP����g"?w=NÓ/r�4�ʾ��%�ʗ��Ƕkq=��|�����"�ťuuxH�r2겸��ن�M&�n,=/���i���S�*f�� �o�1��K7��ѫ\([�ٲ�;Kh�;�[6����b��ozM�X!�6Zո3vN��`�ܶ�B�%��L�QW�3eVui�io6v�m]�"lEw]P�:�P��2*���%s����O�����e�p�����'���S,����d��[::�=[J-�آ�܍��Ҷ/K�QB�$���Q3��f��+�`�Ubmu1-4�cKzV�.�Q�6�R�'-�f��B3r� �7h�tu���V���ڬ�:կ_u���7:��u]H��L�>^�^���=2X��A|u���j�=��ؠ�֮��\v�]�Ϙ��)����xTַab���l<��H��	�%i�`�|c0�׽������}�Rˤ��O�����D*�F�VC��m�V$:�A}}T�f�\�&ՇS\�b�����c�#vf����W
��,��
�.16�M�%���Cj��=-�=���[�7ܢ]��8*�a�ih�$������t>d�7�::~����&i���F13]��tc���h��׋b��⁞Jm\�{6�^�=O�Y0kܧ�'h��X�;Ε���!��L��0�~��p�=��Km`n�2��{s~<�d��v���u���y���Y����@f�GÖ�q(x^��Y�t�0��|��<���h���س_	[�m�qsÝ\_ڸ�C�GS
��ٓir��^�b��/�Y7�;9t�K���]3��R}��'m�J�Ҕ��!��j��������Ӄ�k�X���oWb��em���ي(�=�Kr¥j�1ieaP��a"{d��'I�/�勬އ�$�f��\�	>�3��\�(L�����q=�jv�v�8��f�G�	����]^�(�^��/4�m�Z�AB,�x�N!w�˼�x�ݒF���s�w	I���&�]�eX�u�ْ�O��Q&�iG-0&�8�f`��w*���r4�]��|�]�í�龆γ�E[uWhR�.�Y$YK"�`C�c�>Sɸ�36Š���Grպ�5�|%�b���2�iƱX�Qu]�f��J�(A[�%�ؐ�yy�n;�Z��;t"{�}\��{�lB�V^��t�V>5�qP ��K�oosFav{z����Qf5��8R��ļE�[pS<k�E��l'�Jl]�LM�ss[d]L�0��\��N�u�st����2��*�At��Y�BWY
�s����3�k�ϟJ
����gr��f���W���D��{V��ה%�\�X�9�)`���;�mJ*�^q���w[Il���U���k^0d��'PDv�n|F�,`��2gzh�ul�6�8��{y�S/(���-@�O�4e�**�F�<�w�wwQ���Q�\��b�Y��]�M�B(nk��W��{�ٝ��[�+5�9D�^��<���Ⱥ뫛0������d�˵-��6�YBf��dT����t�;!�z믲#뾺����uAA�
 �&��И�Z܎��ԝ��FI��T��<�9�Z�[�l�n��s�\8�o��Z-�4Ӡ��x1\��n�g|m�ֈ�20>��F�esd�����{1T��#EH0S�'J�����]����)���M�{�f ��w�|��6U�C�Z�D�;��t:##��7r��:;be�ō�YڽBMdq�si�-l�hOֺuu����O�Z���9�K�����$��SU�Ϗ��"8�k�X󯔿�Bj9��`#&���t`z�
�j5����Ⱥ�a��GN�U�,h�nn8�w�w�3������Y(�Z����u�g�u��ednk �H��x���$�^���_]�Ε�I)���+!A��Vr�y��C�����N��+�
�w>��S�<�]��jo+�K�N��;졦�N����|l-�ֺ�n�-�����.ICj�`	E-[0�6��"c'	�掻ѵ)ʂ3h&�^,w>O;��§[���42��Nr��P�6$���+��+gc��š�띸��d�vZt�����s���
��39ed��oI)($ r48"E�2uT��r�%$��L ?�������
�y�E}�(�|Rښ�aA;҈!�d�0��(��;Hpw�򦾋�*FɊa������L�d��^+sGq�]N_D�Ġs2�� ��wd���G~��12{��O�$dc׃��toov<�$�u���o��K�]�NY8��o�UW����XfT�8�B�����H�{����
r��g+N>C])ս,�ɽ�����{����v��Ю]�)�(��V���v�3:v�=Y���soN�)cb�:�gb]��/7i�xͪk��\w��;�&0a�Q<���^eN��	�aN��tٲ]�ٻȈ���[�A�����B.�7�n�p��D�m��wE?�i�k3����d&j��/�wܵԎeidd�Й�ض���
�0�m$oC��3L܊�ݗ�0��o�{�˩Ǟg|�����������'$N���e���Č�|�؁
�ZT<<{��Z=�Y�8f#������+2�f�Rc�I�\4/��Ќ��C��Cݳ�W˸8y�I�]w��qǗP���+32�K*$�E���+��-[���ȓr���KUjH�����c%S�� �E�u���u+v��N�"��V���W]ϧVӇ].�Q`�&G\�X�{h�)u���3J�ˬ��I�LW���YlO�h%�aQ뱰�[��F��*I�<�=B�v�T��T�/6����)2��'�A4k��|��Y�{�wpT��%�so	�쭇6Bz��n�gݶ%o9xN�e��y.@C�M�����
�b�FT*dykP��u�ʼ-��\�jdr2��q��-��7xjڛ�����[r�x�f1X��7)Ajj����Q�o�	��c��,r˧��5�a��d���Z�hYc�3��.5��i��p�RjC�V11�F7�,�fR˨�ܲ�@�T2ٕ���$�����%��(�$ 
�Mo�y1�GJJj�[��&3�v�Í���G��ιeb��.�Ť�B6_&�WW�Ȯ�k*�<s_ۚucew)E�k��Z��n���0!��Y��Cٲ�e<F|u��]H�,u��!	Wl��.�@3�\��F]*v�*��Wk�����i�.�U#��[�d�PkI���fX]b�;��k��38�q7{�|yS+i�׽d�?"2�_q0;�ơ�팕M�\vn,8U���;�6p�o��x#@Ar� �����*�䔖�����5���!�:�:���L�ҹ��;�$��2�����r�/��u���wC0��W�\��̲&�I٢d���lH5w�W�r����qA��u2��� �b�X���ѤF��z�
eS;G�r��"����\﷗>Jr�(�b#��W�j��s=hoh�s��vK�A�L��E_%J�5�d�YCx��K��͞b�)�(F�%ٻޛ�%��2���*t.�m����Dn7�D#@�Ճ���mu��T�7�":讨���]c��'�Zz�����(�pC3�E��P�{h�0];�Ų_[�W�x��l�x�����e1�v
��R�����&H�����)�-u��̫tfX�5k�;���+���i�4M�s�H�FZ��Dޠr©t�T�N�5.9y�iC���Ǖ��	��C'b�;�vX�͍�Z�&U&6�r�F��Wգ�j��%l��^���I�z���r��8(��Lv;f�YxX/3"��N\�1�Z�f2��d�+�(V�25�7u�'Yz��ǆ��\�`��8�l�>��ejo�5��8{,o<;ݓt�Z����b��d�R�hv�G���xE�R�n�qv�J�*��U6�at�+�������r����[��i��ee��U_3�i��y"��Q�2�7Ϭu��%��*'xJ��x�]�� ��,8#�-�+����7H�%"�֎�AKg>ݩ�e�+T��s_�,�C�>�k.��� ��s����JԦ����ƥ�fU�0����U��R�
���.�#�FC��@��v�?b!��]
�'���}� �u�i/+[����w׽Nդh�O:v��n�1L�`��0�yґ����A�ވV�Ӹl��Q��`�Q��ː�׹��#9􀏦���|i��dCN����Yjɭ&Sx�]��ʷ%�D9FJ��;w�;�i��Z���ٿi���ʚ��q���9��d�jK�\EU�7n�:��!�VeK�E�^�F�E�gm�<7@ݒ�����*>�]L=p>/6%�v���˹��gF�7ZpR���6^�Lk�0�p�(��-U�U��lҋR�;���Nơ��	�N�^'�����APV���+bTj�n�U�]�k;3]ͱ�L�ĕ�[��<�����ɓ�>(,�&�e��(�'�[��t�dPdr���zF�Nh��բ�v��p��ػ8ol�`�:��d;zfY�w����!6�R�r��˝�ze��I} \�Z�*�>L�x�	��]��m�u��Ǘf|�3���+]�u�2��m�t��pҙ\��v�]��c�1�e�N{m=nd�V�+�����o;b����7�j�ɱ�VJ6�l���Ӳ�V�����g�N��U��j��Y}���g-�sK��EAT;Z�]n���˻��@�	�t�Y�bĮ%F�t��P�d��7E�G\�vZ��J�B�B\K�fk'{6�-�S������l�Qw8X�`Ю�jL���w;yC��]��Q$�,��S����r�j<�c��-v鼻�'���wu��U��l%b�Vݲ�0cX�_e�&��6��Vw��wsn�j%�t�m&��w�L�&�m7�J�x�*�Q�o0a����y���a�=���
�S*2�λ�
���K�igۛE��u�ӳ�Fo윳Jɷ�xO'��ԧ3m،֙�z��g���6��\������sOX �6A}��l]�sX%ʝ��2,R�ZJ��=J�G��g!�'���%t�M���WNm��-eY�%�j�d��N�j��̱Atyz��5iĂ{�D۔�����g��\��#�6R��yh�����c�<��_.�Q�(�[hL���$/8Чo�VUws�ս��r�g^�}ۺf��dl��F[�XK�R��;z�X�p�}�J>���tԐ���(�U�+L���*�"�a!��T�S�/N��S�)�X�+)]�6k	���YJBj��c�u�ٙi���aj�8)ƌ��Y�+���	���t��q-���K�Z<��*>���\Ғ�����=�����N�m��e`&F�8���W�g <��m}�S)0� ��p�Ow��E&2��Du��V	 ��2���r�b	F|�v��B�eɃ!9u���; ��rb��%GY���(��*y��B|U��X�u��dS�lE�K�}{٥����c��Z.ޡ��}�Т��{Q�A$�=��z0\��o�_��u�v�xo!˱D��R��͍g��lZ�f�9;w�Yޓ-n��*'\*}V�[�N�*s��L�}Z��pR��]"��t���^X�@�*���ncYXD�Ż�[�*��]i}�d��U95��J��������[;�d�_s�c�����U����U�޽�٣)�h�v'4�I]S!��^�U���{WOd�4$�Rv�гS)��6����*-�uś��_
J�bñ;,��l�3v�]�,���~�~ʺ�0>\gr�˂Q�h��6k`Q�ܬm���I:q��i�`��4�j����^�q�|M�<l��T�PI����I*q�Rp�K+�іm�Oi�E'��1�}Lõ�s���L�A(�t��ܽP���&��=�h�G����+���xse��� �Z���C#�t�k9ۇp6'+`ե�ic��"�!�||�N�9;���f8�&�Ƚoy�1JW+�2DN�� 
  �E�@Y����!��#����E~;\���+]YFF\�.�8cY��W^t%`����'���2��S�k�¤�{�mv���M��m��;j������դm<�i-L}:���e��,m����3$0�=6x',�u��:f��;'��]�ҽ�;O%�o���h�k�FI>�f�{j1�5�`i�6`�/���^����ꮱ�ӻMu	IX\��Iq?j������skf�
 ����*��ݥ�@���oqAk&������ѹ
�ry!�,:He�s.�}	�-���.�l:{�������5�tڢ�}�\`��M�5Qf���gJ��UrW"t��nc��z�v� mz6i����T��<|/vg�v���-�|%���x5w!{�6���{0Wr+| *Wq�d��O;A9\��w,�3�@��n�ly� ��]M��C�8��w�؍1��z�;��>;w���/�R�zx�ݽ�#`��Q�EO�J)`����
Gg�5�z�����`�y(�F"��J�P��˗�{�VǘJ��n����#��C��1yLCX�&��h��2���.#�i��MZ�*<�1�6���n"��\G��V
NZ�Q�Z3CJזQDb�we5�1x����ՆJ7����E�����{���J��W�ٕ�*��r!ī�ሢ��,ӡ�*^\D��i�M�5e�.��=a������Oc1+hٖX"����j#i��qrYۘo.Z�j�[x�E6n�3��hQPt[v�Tt7e�ֵy���+U�J���Lb�U��Q��A2�'�>���h�����z��[\�nGc�A�v��|;�5k�1�����
q+���7$�?�W���弲凳;D�?B��i��<�/m5i(|�ͺ�m�(�	Z�0�m����u��ܖ]�h]	Vਨ��\lȐ�*R�E�V$���A�)͋�[�@���)���gCkZ$ܮGP����4�*�]H�0�h�>���*&���k+�S;#���:Y�k�9��N]��:�me�Z��� n���wO������(N�7P�螥���~�?�����+�����>�2�Om���Yt��
pB��%K�hf��*�qic�w˖u:���~��F�A������uƻ:8z.N�;��y�d�1�X3��)f��T�x�t=Qb;�N�X<�WAP��^��Xyؙb�<O��U-y��l��u�f��k.��&v�i��R�ujй �[�S�p^_Y�%�������g\�w,mq���&�[�3���1_N��/
�����4r߄���dNtN����ʰ��zP7ɖU�L,��+��[`�M��\������Ժ�.�f3���T0s�S�2�)�f��<�	�W�~�{H�0��K��gͱ��6" ����<V�ҵ�"r�w��y�h=�k��EM���K�Ϊ��IÖ�e�l�/0��8���{�9��݃am���f��E�w��+�R����e�'�|>�;��x0�h��W(�.pF������5j'���Ź%ޖ�����NB�!���Z4�� �FVۮ�GU^>�N�Z��b�+NJ�f;4F��B����5R{�DBp���x�1��Z��6$�sY(�t1\m�{�4h�F�v�f^�p��Pw���j2-�j�Yp��z2����dovVA͊{[�w./_�$WFc�	��HCT���#h���CCGݦ��o��������C�s�؆j�S;uYk9Åd:ڗ��p���!Jﻌ�qKo<��d+�bO�T�C(Uݍ�t��h�طʤp����mu�C��yB�k��8]�
�Nv9�hv��*VS�� 텒��՛15�*㳳k�"�X���|����A
⁑�֋���&�WhUܬ�o�Y�`�lD��r�X)����o#���f;f=W\��-=�v���~�Y�x����,�{7y�#6p��COK��Zn�j�+��'/Qp��Y�XN�1,����0r:�r����S�n�6{�7����{��W��z����)���i��N��V)s$Ɏ�:m�wcK�7���ou4N��[59�<�}[Oxs���ЬT��b�ܮ3��"�Ў<���f�S�,6=�(51:Z����3�l����5$C��Rәi_]�gF{�޼�PΦI-�M�+����[~Q��`����&�j%��d��[��y�ȹ�g,R�i��7����Q��C��h'�iU��^���D+`2�)�;p��<���NrD6��nvG6!e{�Yt�7��]��{���G��ul)�L�wHe���<��P2��AXW����<~-�
v��6�"�'G-ߪ��8�]݄���p}���y8/mL�-۵��������n�!>�[�6��^�1W~.�<Ri�c,�S�7J�}
*�ö���OFTPn=)�M����ݪ��AJA�ޖD�0Lg;�ָ)z��8�]�h\t.�F(A1� c!>��q�e�s<���_Vì]������%0l�q�*ϯ<�����ƫ�SP�Mw�6�kݡL@G�]�xGg���z��zq0�f��W�]�ЩM�W�
���B�C��y�=�����&��z�:m�%7�T��|W�l.'OF ��#��=�F���\�Fk�وgSHw+W\k����r��ح��;���m����q⒫ʶ��ͥ/1�s�EJ���(��X|���y��x7w���G{�ͧeu�D�,�j]Aݸtۗ�U��RV�ͭe̮��w$*Tw>�W2w}\K-s��&�z������&�VQ�H��$=�>Ѭ�K���s7��fVNZ�3f;�����T+�[��j����q��z,W��#4q�8�X��;<�ǝM�\$�b���8m��n�W �5��;�zb���K�2fK'�8���o���32"�v/a�b�A��!��z�q�����N��r��0��sӺ"��ט�w��Ë;7�N�4[�z�^��r˓���.*���XA@���dӳ�
{P�'6�m�]z)EK-Ue�@Mذ�>��uKS;8�0p#R�t �Z���A
Y+��f��f=��py��yOr���G��F*�p���fJ���K)�$5���.ˀ6�	�8���򑜜e:9��.-�k�{U��m����⇣:��U9
%ZƤzo8��.�vs���wsXim�pk-��'�I�v.����Y̖flS�ļ��$#Q���Ӑ�w]"@�.�����iy�RЪ�+p�|�e����Y�������Tz���*�aqS}�:�}"��7�k���;�D|j��7��MGY���z��j��h��(��U��M�G����]�σ���K��0�<�;c�a��.sř\w7ˈ�Ckgw0��]�t���Ȟ/�N�Rr9ݦ����eQ:ʾ�a�)8����W�l���`VQ�b����f��̤� X�o�����8"ݳț�x���wpo�S�lv�R�y�6:7<�x$r�C[i׫�O�z8O y�e^�Dا��_	����x1��m�p��5`d��Ǎ�%_#��շ��2&�H�ݘt��)2��.;�-��ZA��!c�����S�UEf�n*a[�Ĭ�K�n/5�Cb�����T��	���．ٸ]��3�!�)� +�싙`�q����,�O��j�kI���s�� �r3
= ˜���/����*R1sŪ�g)X٢�Y���̯P�)ygqz�ڙ��ey"�f͜��.󥦅�Q{���W��h���\��lqYr�dۻ�V�P���]u�F�(BoN�!A�B���r�<�����&�ϵ���fl-�#���~�����{��]C�G"kj*j�	��M���'�W�Q�T��^^�fS�2$�A�ЧLH�V�-����=�E�9=��l���\,(�]f]m��W����]����E@/�n~2�ݲ'�y,���h`k~��{�u���3��o.�O���Q�k9��Q�Yɸvْ��`���,��יx��r`m�mW�v�%I�X�Q�NP�:1_;�iˋ�
�3ɮ<9���t�e*��c�R��-��4�f�=�^04Ag��ʸJ���|l� Xt�����uu�҈4�+�����%���t��;�;3xZU՗ӳ[�p�$Z;OOC���̭���噊1�ڛ�!E57$�e��6���Z�U�Z�waܕj)�;������:��(��K��	�nr\Wg9�Ιw�s�/���e�7��f;���W!׽n�J�:�o��-�1���t0*���v5%ýn��w��f��Nl�{�����ܠ"Cwݶ���t2�襇LWg�?�U6�ǫ�I[9�8��f����?~f~��8�l2����*�sJ�e�,�
]UE&bUA��}y-$l^L4�a�j�ʁ�BQ�)���F���!3yA�.���Gk�'�@#�w�P����3P`�h�x�ҧ�������z@��a�`���2X�ID+੤$%�T��V�;h�Բ�Eʤ#و�!T�\�w�	��]*jah��[*��x����j[W��4#&�16\X�e��x���,��+]ʻ�3F%f�[N�2�P�1Qt�#�%l�T�i$�t������Y�-���͚�JU>t���-�S�Qf�*ফ2�U�	��}���rX9T��N}-EQe�e��PvZ`�hV�Y���i�m�,�J�6�m��m�[�y�[dP��Gٗv*��5�Q+~n��P��� �PB�b�k�QF!��oV�u��<��R�3J�UTUe��4�C���*UM��h��iVң�"���7eEUV:�t�q��Gw2�UJR�t��Z�����w(�t���,WM6��*�RʅAUլ[v�nٌ�&�Gn�9X[b(��b%�Q6ܺʺ�U��M����\Ebm*�`���j�]T�\8�)��UQ�UQ�j��1��U����m
��3-QEk��2¨�k3*���a�������g=L�[���fo0��E����(hj/�;��^V�C�}M�a����%�A��obb��&"),3����w��c����4�%fG'7����
�۷����Fժ��9���>,�E����.6�|~;lg[���۟Gʪ3��.1W�Cg1Z
zfwT}�w]��VX�f��B���.���5��u��g܈���FZ5[1=ѻlUѱ��������S�5UG�#"/�0Ui��BW�V�#�}u�|��x ��b1^�+5~���������\yVz��D.�7?p�*��(�ؐ>�e���O�� �u�b�
��7K^`d������]�|���+���"�\u��y�1��]8�)���HK��(��Z<�odّ�ם�����1вe}1�x�\�Xq�qd�M_���E4Y�c��A�&��΋�C��c%��;�:��y���|b~Hf��Y������k��D�������qum*�<��_�?��]j�W�����O^�[6����)�}�W����0�I��>�	e}5��ϭ�3�ct���k۱w���֗�w��}B�u�e*5���.I,7�G��Hf���64@�����o/x��z"3�ޡXFcʴ-� �	�����Z�Ny�����fx��nӣX�w�:����G�d8+U�����t��C��n��:����ȭ�F���8�3�����ޥ�̿ȉ�G�=i���_�U%,kQ��J�(,�\KE�^�8�7�P�_�K�U����튐�oJ/��{&=�S�9��1�1���LBu!O�i�.�J�䇌���Ԑ㟾�������������? q!��d�YI��s,���x��I��dM0���HLI�!�y`,1���:o˿{�Ͼ��I�=I�l8�>>��zȰ�ԁ�0��d��4^����bC���bC�'�~��י�ǿ]�w��ԁ�I�?sD�'���e���E��!�s��
��RB���6�=E��M�י�~^����<�=����&�iHz��b��!���gl1$�����Rz��@��Eϼ���Nl|�Y���t�~<C���Xq��Yd��2O�@�,'Y��b�������m!�C�5�ǧ��������~C�Ͽa!��O3^��4�� �&����>@;�O:Ȧ�aX�>��}mr�K�ß�_D9�D��Hc'�Y6�����Ci~�������`s�i$�&�I9�'��l&����͞�;����*�,���(hPi�Q��U�F����/{U�F���R�='���\=�e�Dvb|D���F�t��B��[Նk��]g3�����y�=￿|���=���=����&��C�O�h��6�ɩ�=Hq�����d�I�O�!m�I8��s�_~���s���.��~��>C��=C_�C��,ԙ���$�!����t���Ԭ!��<I�0ߴ���>֤��1$8�ğ�C�N!4�����N0��I����,'�i�8�����b=����� ����A�G����8ɻd��m�~M哈yI?!������X~Hz������ԁ�>�-��O���������i$�>��I��u�d�I�M��`l������"��~O����h|��˔���J�޹7ip�Q i�HQq�.��E����O�=d���Y!m u�yI�Bh��i��\�~�s��tj�7�6�
@�M���ā�R�Oz}g�CXI���=Hq z�l�CL��k����Ms���}������ē�>�q������C��!�'�4e1g���̓�,��(�9������~������!��쓩$����Hh�z�$�$�yh|�f�=dP�� �&�Y2���L���w~�y���}�<H}��C���$4��u!�Nr�b_E'��$>a�"�{�Y=�	�?�=�C��t�_�y�#Sk��m�I+��	@�i�X�ð�ڭ�E�لz����|���V��\8=�X�	� M9�|���[睩N�'�y��H(k��{�~���!�w�B/l����'7Hu	��H�@�O�<|B��Af}a�@~0��3�{�~��~I1!�!�x���i$�'PRN��H^R~`u�hO�}a4��}�;�y߷������@���M0?!5�@��p�`_��OOXOP�'�Hv����O���<�׽��~��M�)��Cl� i���=a:�z���M2���$:�g�<Hi~����M~՟��>����}�����M$X�O�8����?3<�� a��R^$=CH I�x��C�X�{�7o��y�}������l!��@� ެ'�:�Y�:�7ܒ��m$�О����Rz�~f{���-���~����x�Oa����2O7�E ��F�x��_�!�g�l��MO�?2~d0��ǆ]=��{��~	��4���Hz��:�o�:�ē^��gل�aFo$�ì��Y����L-���Z_$��Lz#�]q|&�=`'����3�:�3^�2)'�ɾ�B���-�h=���o�y������O�P��L<Hu��!�L;d<d�>�� a�������i<x�u!�˜����������L/1wkA�ٱRz��|E��ҮO�w��c[{M1
���~��~��^��z��u^)�"U���NL����7�DTiݢ�m���X�^�FϽ����w��ć��'�W�q'��RK�솒d=`z�w�@�	�)���)&j��	�u�ч������z����1$���Y<a�!�)'�z͙I
ya��^�u'�&�)�zʄ7��/������3�C�l0������C�O̓�,6¡�G/P��ya6�!�dP����%�ٮ��/�	��2OXI:�Ԇ��B~Փ䇉5,&06��'x�>��{���[��~��~Hv���C��&�~I>dճ�C=�8����m%d<BhOb���0<�c���7�~��B'߬��w�YHz�~`,y�H~�ܓ�&'d�'�ӨpՒz��������e��}d<d��i=`g���ya�<���0�`z�ԛ�H��i"��S�N0��`q���ַ�����B����O���z�S'�&�?&�d����=a5��!�@�C�\�*��	�lgϝX�t��c�s�"#>HIw@�$�'Pj��������0�:�N�P�'<��O��~w�����	��ߨu��MN��z��2�ɬ���i'��d8��������]���S�^fߛ�L��1+�N�x-�]G�-q���Sx�j�ȋ��Io`7��o
j��wP��kI�w�v>�����Њw7Ƿ5�]����CO��ܐ����$��i��/�<I��m��Hyl�wI�������_wR�!�?���:�k�=>�b�>�!��yN��>���w(�_N�*��͞"z=I��� Ys�ﶤ�Πt�X��U�����1�
[e{ଞo!g�IZ��df���sڳ�[�8��!��zy՝�ԉ,E�]"���o(I�Ǳ��4�(��t�E �w��f��+����N2f%nm�F���� Ѓ�Y��w鉊�v���[�[b�GB�F*1��P1�rq ��Yk�<2v����w�%K�fp�N��ssfhǢ��7�����w^@�K�a˚�P6Ҵ�e�W��V�$��ԴW����}�Ev�[��a�ɘ�O�ܮ��x��S��_I��{���R�����$:\
	աLL�t�k��oEq�3�L�C���z�r0s��w~��\�ynkJB�{us+�pxu,���-�U`ظ�Vg���ӚX�Ǽ���O{q�p�U�;��X��滌}q����5,`�}���D��J ���U]^ݬp�O����s%�>��]^��7�s�v��ɒ�8����}�K��+��7X�`�y��N�zYa�;Yy�(\qRF�*�S��EF�����t����UL�foh}7zd�R-�HȦ]N۽:��w�"h?z��|����������w���HH�BE��H>����h�J��CV�ݾ��\S25���5�1��TI��>��OB���˴K��Zw�����K�Y�fP�Xk��c*2��۸�Z�t�r�(3�9쉵�9�4@g�x:��O�pE�15��(Mq�$�{6`���/Li��|LΥZ��;�bJ�u1Av��AC��m���-CqR<���ü޺GK<�.��%��b �y�P]9��4ټA2�6�TV�X��ْ������I�.m575�]m��9�,���9�����W-�ɓ=�voP��]�0�FI��r9:Qa��gi3��Ǻ����w�x�|�w������E�BBa`����E �X"��u���{�����YH�鎞7����_�m�,���SY	+��YJ��1-�	�he~���[.Nj#OȌ��7[����$�I�',s�\��$~��)��'�ܤ���i�����@B0lC�ƃ�ЙZ.�:Z�f+��!\Ppv��5��/����/:`��x#���tQ�1�&�}���}�7�I^�4��)�I��vs�*���δ{��$���J5c����o�z!xN��5�����՝r���0�ub�?�>j�p/U\P���T��xN��c��k��R^�HM�*�G�v��Rf.�.�u}v�k���oゲ�^�P�;O�)[NdZ'}�/Xv�2�ko(�Zst��O�Qj�-f+�4Ĵ�U��NVk��%�G���,�v�����X���V�0z+��3iXO���荧�HU�pU��p�U�o�m
�w�0��Wɖ�yZ��庳�Reۭzs:�85o_�
}ҍR��g7�N��y��Jv�h\ۤ��읡����T�9��C�p�eX����VJ��J��:���=�^K�{ŕVN��:��tTN�Ӯ<�b��٘"t���F���+�:A�[������/���	M2�A�[��ڸ����y�SD�c��.{@�E���c{jD��V����জkT���OyO~oo9�~a��-�X�U��������r�9UN���%H`�B%bB�WL�����d���i�B�����P� 2�2�Bȣ)$E��0�c,�hfTiVEX��J즥����{R�d͎m
4/~d8�A��/>�K!UCeG���U�jJ91�ă�o�춪}hX�) ��n�)�I@�Fe���Iɓ*��4���X]Ϣ��R�V�
�ts��ǃ�
����H��z�-���6V�X�8��w��©\2��	Ev�Gh���Y�w�Cfg̸�
��6lZ-dp*
e#��$Ħ*�4��m�4fV������L%I�J&E<�2تTlQ_���P�!�;J����m�V��z�,�ޫz�Kx�]�c�����b���~�}�$�	$��~�X����b5��#S(_-EOܸ�<���j�`��7=���QFu���0`�5�T�++�lY�v��QW)c
�%B���֌T����a�ر]Z�#��CH�Kݖ�T�f1�Lƈ"*�<ʘ�-�N��Q�`�y|����V�dլ�|��6آԢ�6ԭ�X�KUQUO��^yxj���������i]ۦ�:�ժ�M2�/_�"<M�0�۞�a�_.[7�_2��bC�a�4t�R�抰q9h"�e��T�[h3ī.��7�:�6���3�3��_R��=����M�@f��g�C{��s�]�̑
҃Fp�p��/�=�z=�����4�
�~��*>*o~�U �?%�L�F�^t:z�$:z$���Gt��^򺋕z_��\1�<�`�8ፉ;>����^+,��Ӕs���a���cFzbp���D��ݩ��rk����%�����Z��EZ��	�S�B�#v��ۯH��{�G[��,�qN糮�+ca��aM��N����Ƙ��1��0󋔇B��\k��k3f;	��8���Q��n�S�c.F4�׌ k��s��<E=0��w��[h\��;�����+]7뺅u�N��������,;kq�=�
���C�*������Q��	���Zn�\O[ܰ\��g���09Ʃ�V0n�#����K�"*���]PD���@��@3�鵸����k��쭅����5 ���B}�F;Tzk�j8���/e[e�b��ܡ=8yt>}��@�:Zƅwf'�U�9�b$�s�Ⱥ�x�.m�뀸-aGN�mWWW��Sy��ɘ�A�*���I�D_N�^���nMֱ�٥�*����VZt=�㼞7���ln���t�x�n��d����wJ���5Q��wNZB;��}�M�2f����S�W(n!�jr�UЄ��`� ��@~z"=�z�x�-��ô�Ta9��OgSHr���E��i�H���O�-S�7I��_E	9J`z c�Iw��(��Q>�])��.. _֡�4�P�-��V�3۝�8������CH���?q�R��^��OZ�NQ�P����"�%�;�K:IMCf}�v^q��5N�{��=�b��ㆼ�Sl*C��'M�Ԓ�=�@�H��i4$OK�]Et�
��-;eqW�����l�8V?��?(b�<<��!��9��H���D�k����z1��`��r��g���1M��2�7���\wQ:lr{j�^�t���0��򣢲/yR���l�J�,�w �h%�p���lL�rut��v��1�͖����'b껒�8ݛU�=�(dm��Ó����'�}6u�+7���z=�]^f�z3_�1V��C��N�ט��W-Y�x;꿱�Y��Ej�U�N�9���,4FV��BPCژ�4����s�-v�maƎgi�7���-i%�?���9��L_Q��Q�e�N��;5��>�?Rz��a�,���:w����/��N�ڬ�Ri���8�͘S8�N�c$1z��gydb�9���O.�������,���8�eռ0o1p���ڷܸ^�b�!ܬ�}S��~���ѳ�]>ّ�'�a�K������v'd�ʿ!Nt��毐�Q�A5;��`�E�_`�d�].�#���ڕ��H�+ɻ�)S�AS��t����]S1�P�㣕��p�.6Ej�o�x�ۯ��uj���L��!�|޽���M������o7�����f�-;���2';3�Y~�u����pPJ+�ۜW:�.)@!��(�ӓ�(�������:�}�/J���6�jq:D����^R���W�tmfȸ�V-�� %ə4f&}�t���PO,8JNwz��m�kb6B�i/�ü��C��!�F�p�%Qs�;R�_�C;_[n�Yä6���8�;eY�<*��sۙ�z�&txS��H��Lk���r��j'<*ѹ�5`�X�^iZ�⢪�����K�D	k���S��̞��g7����5~C�&y�Ť����I�2Q:��ʽѬ�%�V�6���(ڧ�l�"���2��=����o@(�����+��za�����.���gJv�:�j`ʕ��B4gc��F�J���/��b���:�����᠆�Kok���{V�9�0L�N1Z�{��hS�D=%�!�o)1z*��ܺ�c���h+N�J�E=絯F���en�|#3P�Πx^������n�p���'�h�(�p�S�r�5.��Ӌ�-��]z�s���J��j�O��(�TFq��,�9|��4�}�B}���IxUx���a0b��iF�$#<�i�֟8�N]{�n����!�?s�<�Qد	2%eF�l�w��Z��ur$��:w�1�[8|~��׎�#O43}3���d�Q�����M)f��ɗwq����	��T^i�	3�T��H 2��X��z��_��Y,�V�D-?��T8"M~;V�;��b���t�"s���i껭�{,q��5b�k|�!����5�l�<��1,�����Ğ��N�0$U�K�k�����ف:���[`�ERK7�sz����b
n�7��7�>��m1Î�5��qu-�B���D��P1���vS��9�t�˒�LF̼���K�W����Vj��vc�֧�s�0���ץ�7�b��"�x��^g�Z*�#�7���_O&t�ko���#~�
���WO޼<=���"�<�<t��p���J�S��lG(���PNnvFT?4N8��ث�Y�2��4�-�c��WP����޶,ժ>��Z[D���jÕP�n@��*O�*��+/�>ˬf⎱�LVt�+�͊hi�kK��a�aX��S��H�o��7���:�BY߹�-�%g��C��w������Qb{g�DΜ;hi
c%����V��ʿv;�W��_g��Kk��}�<�x�.#O:t���II�����go����hz�r��>l,C�Շ�;�$=Q��nOa��AIKn�92n�R��rJc�o�	וظ�e��u�4�S6N:V�]s�\��z��cxc��L�\�B��V��ڕdda����|���kh2S|.�n�Ǻ�ҕA�Q۫�;eɖ͘C`WVR�C�G����8��}P%�����e�~0]���+�=\n|�u����p��+y5a!������5H�:xA�z�t��U���O�/����<N!��^"%df6!�,��=�����`�$�Z��"p���6��U��ɭL�'���ݧ��;��w��#�g0�;;\�����g�����f�x�Y���Βp��BR�����]>d��fOw$��b�x+��˻"����bW����{�T��h���O����.�i�W��"̘���=��0�Α�b��9�Mt�D1�!b�c�ú�c�E��2����W����Q���\r���.#G�c��ɍ,�6���=�Z�����\c�Z���,W�8B��kR�q�KlR����}�y��ɶ�O�5v��~[M�ꊜ5ӆ��N���ժ}vˑ�R:��m ��߶���Ux��:yJ`��4�=tc��	?3]O�!�����>7>�2�k�������j;�"\��j2D�S�4��ԉ�\�)�֋�k.F�C=�H�,�8�����K���Ѷ4�k1�N�qB��u��S�޾clrxF���D��H�9�p���Ws��0'�a���-a�|h����7p�{���Hԁ��O�D���(r�z)ec$~�w�������QۧG��1�#��g���ir�lnw�9���	WR���z嫗oٶ,�-v�|%�\�Ǯ|E������a��9_\��(��YMa-�2���*�v����#�Cc��ʶu��s����u�؜Q/K�|�r����^�nH���~󭓻b}[ד�4r�@�1��+���Z����e.j�K�T	mKTry��P���
7�W	�ר:��d��f�zJ��Q�z��n5QU��#�����M{o�}�ŋ�͋"��ʣ�y�>W�%{���e&�����ӫ���#%�J���߫&��|;"�r�=*�:��I�#�Rb̸f.yӵB����a۝�<��ۗ��n��}��5��7���:Q�o�XWbS��n�7�HI���r�[��.LLt%}8��� Rڌۮ�3/�e�%/+�DK�<v���:h���㦍�p�%��DQ<����<�W�J�u�:|d�UF��'aY���Q����_ve��:�^�to����bl\hMs�$�c�����[:�{w�:Fz�/i�k��,-g<D�^�j�/�s�2��`�/-`���7w�Mơ���1ǹxn�X|g��9��u7��)f����;*a\R���^W!��^b۩�8�݁aiSU�lC9����5�qn��GLk�PsR�IK;�Oe&�I�SM]�a�mG��V��b��_}�{%��+L}2]G0eMב�8��V���ev�9���r��n�=»-���g�e�&tٜ��uBx�]|P��w٦�*�&����u>���u)��0k��k+���k��w-Z,���2u3�*�cn_swR�s��m�qؘ5Q�w�ӳ�^(.tu���ڙ��^q:<��w��g�zQ���O�"t.m�<��x�*�Cvŋ ���֮l   	�Vm�'uc,�I1�U@�$F:�1Yue�0�y*�,[��)]b�bSJ�IX��S����S��ٷ�cAʅ;ɖ1�U+�E[^^7px���Lm��B�XÌ�1E������(ћ�6KQ�R2�L���YT"h�E����F��t��v�g�4'�24�F��٢[ϋYdF�Y,��U�����#�j���]�8���HP��1��˺�	Yx��N�u�IW���qJ�����F�h"�k(鲯
�խ�,� hzT)-)֛.����m�z�m�z�-4�]ZtnT�{e㈭�b�:̛�t�(��˛ME��Q*U�yu[�]81U�)����(#�E\J��h�)�f�&����yn�rq8�#������8�y�.un�is35oosWas��PSVi��Ly�X�A��2�0��7K�E�a��c�ATQ�%�Ef��X,c_5`����)O�exְ�X��U��&r��b�r�Eh����V[Q4�r�`�Z���� �J�ה��PAI��NR�*9u��V
cEQ�C���QժL�TQE�4X�VUkM4̲�3�$�A���z!�oh��ulT�vۧX�+�2���V&^m7�����눺���|> :�������F��~;_+����
��Nb�L�Fn`����H���>�;2!1i�A�d�!�D���;8������&�4���*�MTu� ��O�uZ�@�/Q@^��Ta��jpݦFS`W���KEd�+�MJ�`*2����:���&h�j�VL@�30lmc:���B�3��c��+��ϵ}3�7�/��a��8�n�=�<,.�o�x}Qp..����8��C�a���P�>�5ˍt�h�b0!�U�g)}����Z�ή�q�R^f�X���Vf�/V�h��M����	�\�"����3���yUs�Cw��嶠��#LooP�{+��x+����9l��j���N�]8�]��J�*�F���ʣ��5��8q�|epή�x�55���A��Y2Vq]DU.�\��S:˩�wP��]w1�#�-��`�>Z�cc;9zr���L��UW�U7|r3�M�1N��x�R�'����7��0�C��8���x(b��Qߵa�4���{���%�w�y��z"�~��	
վC9��g.�:0(�{��R�p�S�������w�K���U*١*jA�Z�bC� �Hg!DQ�����"�^7z�ŧA���U�遖_pmdKU��\N�u���q|b�,4B*�>��+{=��#	6��3�cI�7J����xCء�*:/ ���
3�f�f����d+�2��}�B5zɭ@���7}�&I���Ƙ4ǘ�P����� k%5}.BA%ޚ�TL���T���Gj�CK�ckJ���4{�Eŕ{X�!��S�M��^5t�!l�%��=�g�!����DpES�|�Y:��7�W.�i{�B��گc�B">���s;}��z�DCva��!>�ע�/�I�]�5�h6;g�� �ϴddwZ�Di��l�<C3�Lc$^���8SE<�������=\���0"�K���)�cO�)���{��w��ƼGn\��߼��]+/��d�cl�k��{�?{Q�***��^B���zv]��*��8�bZ"�q�8��=�3,�7KJ"���W��z�@��nz��D����Kì�1n��󣔁3�^�5y.4������7|^�ƹ��ZGe'��GH}�Iyv�;D��Xl�^ɝ�.T�;3U�}�P�;�d�χ�R�x�=�j3Q���#MD�8���-�л����nu��Y��c�������̑�.��-M�e++������']\�q��EC�'��{��}��T�]$�5_�/�GU���dx�:�rȡ�I���c<;ئޯ+\#4Y�13�_s�	�@��O�D��-P����#K�уʹ3�
;<|Fn���a�܏�{�t�e�9Sq=���+�1�dH�#��u��MwlA�>�Ю�r���
�U�q�:�����B���gWn����Q#ma�W�x�O����#3� g��,���l��H��GN��<E�|z���7�����[�r^�y[����P�cG1�0T�YC�T�w��P
z3�P*ٓ;�QnQ��1���O�(���;�M��ì��-8�I��t�3�yΌ�F�%dX�)�#��L �%dv��-�K9h(s^u���^����T���s,�K5�:��E���u��D�U1�C3!eq�쓵��̜�ʹ�����G��t�[[?C�V0���L��8h5D4�,oy^�K��{=^#�)��3��0��+��Nyh�UQ��[x�N�Xf&T����}gN�/5���Z��F
X$�W��X�U�rH��^�h?i�bڵ&Sܴ��m��K���Q�QҤK
�f��x�@W'Q5妎�]��:_o�(�Zz����1����CˁK.Q�����(|a�/`tҭʇ9&�H�����#�����e�ԋVW�0�ڦ�q�`�m0$X�o�']	�N� ��I��z�g�f5�R���P�\l�bo򭘍�.cS���Lxm�?{�c��Ǧj�1���/o���s�Dj"%
�ގ��Q	ݭn�z=2h\V���2U��~齚2->1�n5�'2�:x��u��9�:���T�e.!17Y��tU!n^��Wݍ\V�U|�]�o�WWo
Y��eu���2��[����/.,�,���ϳ��@t����B�=lq7F{=��u�|Q^Zl�B�h��s7��>Y�����dLt����WveKhQ����J$�O�8pD:��̱�.V{�s�x�"�]�;k�44�4*���x`i����6���nT�NY��G+�Ք%��V �"��I�aU�^q�2����q���0��!Ld�����@t��Z��:��X�\mB�gk*�R���sb�Y˨F4�ZW���a�JD�t�ќ��A�cmq�W��c�↬<{������wR��#<����6qҘ�s��@�%�'2���)ژp�,Ԉ�+96G�?��,4B H�2���좭#w5�9��/�''L�K�p����S[JW������>�:�g��Dz>����f%?	K&@����ɜ��#7��v���%�(��ԗ�yi�ԁ<;Y,b�܉�|����u�=ˮ'������Qz!�"����/ţ�%LEq��]��b[�[�V�)V��Dx%��?�4�R�������af�\K:97�}H�OB���5*zL���|r5T�ZV����ʻS-_��^��|���עв���vL�7ۧ���^�)ק�fFx�r��i���!��f�&чv�vy5�ӷ!T@���OO*EڟmP�;=
�^��'ei��q��P���yFa�#}ҝ-��1�ҕ	��n9�b:�P&B�� �7��.���Z�Nz||���{�ed�K�5�˽�Z�]�Z��S�3�NgG1��3��16�j�='Qݾ������M[�=�ԧ�os*3fʮ�w�"I��+�����V��E���;X`�`0ۧ��CRb�����&�J*n�OP�l�I����0���@�p��_�ի�/wk�Ug�޸}��0f>1��rcg���S�TD�����������=�k�b�d�R$̇u0b}/�AT$FR���e@�0���}֙�ԋO�@�w�0|B������NE��*��뾲�l���Mș�����O��*�J#HCB�Ӯ�2߯;g�G���
�fb�R-4QڧG��n��*%U�oٝ���v$�x\3���˙:v��K�f�Aw<t��I��4�a�mw ͞�õL��Ը�Tf	w��0�CHk�fZ��Jru��*�;��Y��(t�^lY���?!�PH�*�J��Lt��5c����^d�n�z3=��[�YM\꩎R�Զ-	Fw�]�<�мY�Y}�N�u��6Ĕp7���}�G�to#N8e��u��Ü�y
9V���9o->(�C<���7s��}DC~��,��j�!�FzV��F�W���pwǞ�Н^LY��b�_a�uOհ����Љ0z3�E7ut�\�7�Bb��˪��m����WN�׾w���W����?\�.s�v�p�T�����A���<S�ڰVC���'�1X����G�a��7�"r�Ǘ�ud��m��u��4���1/��͌c�����Zw6�0l����g�����j�^��".)eL3UQ���ۗ� I�ǥ�|�>;�l�����B�DΒ4�u��p��(�\p���C� ���l3�>xŎ�oY��ff��Vx�ə̀M�O����͗���_f��������S�fez�]�4q��{y�s@>{C��*�U��g�~�����Y����Fg�1�PyF$�C��bn&�+׶�lW2�C�`:��Q'�<�Ǭ�(T����-��ʫM�],ӛ򬗂�`:R���P�أ����S�z�]������~\~�#V��b��}�8`�cf	��aͫ�}U~�Sxg��_��ȑ`0��dY�ۆj�[Q�@.�q�9ӈ�L��B�D�@�1x���V�x�]*����9��X�lW��\���MG���6&�cw��Z��&w!�I�'=��W��EZ��ϱ!X�Q��~�d���(߳)H��1p��u�;!kr�X���'�������TC�%��xh֡Fo�3��D�J ��N�w/-��}�w���+X���W�tD��ɢ^��l�M`�')�@N\�[ytT4uD3D��t�G��#���������Xx֡1fIGd�[��X:*e�M@�L�yJP��z���k���h�*J�+�l���ǹT�*�yt3P�R��!�K�3���b��[ް��&�;$8���͎% [�[�wx)]r�R��0���[/_sn��Ⱦw��ӹ�q�P��^m���cgp���4�m���جM"]z��yE���cC�zkO3�`XC��s�=��t��a�j�)�2�ߺa[z����u�Ȭ5�Lϳ���fu���4o����;W�K �QAZ>�m�����䂺��$,�n�}U����˝�2�bq�nۋK��`�f�����4���{ \0��t/,�,�Ł]GT���W��*ZI$�I)Ң��*.�S�o��u�����`x�<�+�S�إ�PK]��8{lӜ-VM�mŜ�l�;Om^R�!;u�ug����y*
���#�kI���r��h�u1��,��ns�zO,�:�d��l�q�djS�Z*�P�4�s��]����e��7'��2����t�}V�ˆ��\�ն�e������v<���Tjp�jz�t����=��B���ݓF�b�y}���怺�1�h���FBͺ�{p�EC�v�=�\w{W,�ε)�C��:�]�ε�qpCp�z��ͫ1j�f���և��k�GA}Fͼ�;%H�ۖ]˶����.T͘x�]l�z89���cOD��|�
���I$\IAV$�Gy 
Ԓ��������DQ�[|�0շܘ�X��,�}�X
#�\eb��Oua���t�LĶ���d�UE����a���B���q�\�3�3��I�Y��.#��=K�Z
;�+!��Uf Vq+�ֵԽhj�X�eUXV*4�ی�b�� ��S�ڊ&s'S@���1AY��@�f���PYĨ�ՋjP嵜f�����2�Yt�ePwa��4�VJcG��MXr��B���)$J�Y�ujU�z��zA�8��l7O�,�����r�is$��@�G�"/;��3���S���b�T�c�|�Tm�T�������7�e��"Pj7�F�ֆ���|��Hv!��b�1��=��\�>k9F��C�����8`��EE�w��K���G��Ho��܅(�#E�XnV���=�{x��t�S=q���̘�c��z1cWB����Rwί|v�l0a����b�s'1q��C����8-�+�%�
�������die��1X�"f��Gg|�w����墉�.9j��քK��~6F�yN�R��g�z�q�N��~^;\�T#qC����ZX�����Z�n�[J��=�%����o��*�`Tj���T4���hYs3�~�o:�ޗ`�q�ACv��Qo`<{�V�z7;WX�q5��:����ଜ@�����\zQڛ�Pw+��)i��h����x��iEcq�Jo�#5g����R��w�c&�	�P5=vf����F��ۖ��<0_>2���.?f�Q�=�S�u�S@�"���>��#��Y�c�:�ct�EMFV�c�b�{� &4��:�3,�51pI(��������JV�j�����u
������,$��E�@mTH�+���SNN��i��)��n��M��h{�7�pޯw�����م���Tggf����	����,��6�n����ݙA�h�JN���ϸϗ=0b�yi��cg<+p)��J]�o������%(A�G� �-%��2l�S�lo=��vC2����7�.)}��'��d�E����Sr�o���[t:�+@�Yqֳr��m>������Q�Gy_,y}�L�۷Q��M���Y�f���K Z� A9v�� 7Uݻ���_1e���z�Ti������Bp���oO>!��8�%��C�u�jB�x飤۞Ν���E�[&a���H�a���N�+*�0{�R�)i��C�e��+���=����C>�6�E���Ӧ��P�Q�؎�j�����TeGj����}jݸ*p�yu��'nɼk��u���x!Ɵ��l!�E��_!���W��k�
��Ԑ[�ꢓ��lp��;��6o��py�;�
_�߶��Zx�\E�wM3V�]͇Q��+!Rح�!u��u�ǎy3������N�K�f��j��>L�[RV����kMb�Ӥ��g1's�<�nz�;�n�_�/i�E$u����*3��+0����9��QF�"�K�9����P�ʳ�O]��B	�y=�t����[v�	��w�j��������	Eg�~%��档�W�1��:Ff�p����C�����+Յ��V����yg׬jH����}���t�C���qq���P(w��V�2�׈c+�ڊ2�X��9[��"�"Οeo���M�W��Q����� \�P����@MyX!�ax���cށ�0�iTSʎ��&�51B3��YDe#��j5�2����@����M�F��`JX�7\il#����f
^/T>��g��̹�|�&I�6"\�(<�M��C�	c���z�x|�]P�7.��!ko}��{�^4A=j�##�L6t�E��p���Z̭�m���%%{-��:a؅����g1q�p�Ю��y�`��U����D��ܡ���^K�F�����г��_v9Qu;e>��Nn��č��8�<F�K�-��Bz��]��w}��:�Q�n���<�U��<#L$�Ǐ��?���F��������dt�r���n�qN��bx�xD8
%Y����.��%�nӕ�jb���>�V��L)�K׵�U�V1����)XB�՝y\O�ѹ�Ŕt��CH�d������Bz���f��.}oi+�Z�5�2�γ��2ǧ��=��Q��E���!�Y��͍=~��5�D�W�-��N^�WFՋLy�sE�6"�3W�wE����9;����uY��x����1q9<Ch ���3oվ�OV��Ǝ��+���Q~�Uڂbk�����W<����<��V���b�"k��:_܂
���]�ɴg����A�U��j���A�O���s�i3qA�l���V���9؆���]����h�3E��=��ٝ�S����>��4����l�L����a��P^"�@�pS���Uz-kܹUw�c���K�b�hh,b��	n�1(Q�n�m=��B��j�Ⱥ3�n(u�Y:��1�#I.��*���+ˈF�����kzaUA���]GJ�[��4�Z��8n՝�����o�PCMv�G�f��Ҷ5h��^��)"A�Ǎ����~|cU%�j}2��c����c�m�u5�~|P���5�)���G�v[��-���f�5��Y6�~���ZTkWZ3�\�ךSg�rw�tLxK�T��=$�Y��©�����$�w�9���u�|��/V�ckY"��{��B�����Y�� NS��6��v@�\Ş��N��L�k��5G�ۭr�yEeP��S��ގ�-�v4&���}�����A�-�"syrѳ�����76;�0B�E���4>��s�5.ou��&:�ZG8�T�*]1Cפz���+�`�������o��O���o+ɡv��=��u�~ϵ[� �p&(ҥ1qtf]@���R�	l.������:h:ڡG�T�>t��2yd������pd{���Xbvf�U�E��d�d��PX�1���Y}QF�\��F�I�-� ��ڬR$�������s�Y��VO�!R˵	���ñyWӭX�oD#�`�f{0=#���,&�b���7U�5��ٍUrS�9�5���kb�up��/�gC��uqD�j�u�_y��OK�W;�v��|�׈_E�uW!����P�D��s;$,ˏ���T?#��ڊ�zFƔ�f�p�;;9�&��(��8��&o�\�P�43�H[8��wu8��;<5kP_DD^�I��y_1p��4+7�a�Ȁ�P�6\Xw�x�®iej�@�;.�T�ɞ��Y*���˾�ik��C�T���N&�P��6��l�]3����ٱ�Y�2<_f�{[�<��Trb�<t�ڰ��%D�#}3��R��m��F����F�nu�t��j����_���Uc�6_y�V�rgg��Bˎ�t8�]W�˵&T�OC���)�&L�Í6�ӂ!"k��uZL���ξ`С��N��SÏG�.���oL��=�&?��~�^���%xV@��#�<�Ʒ��4�J��ʎϣþb��^uY��H�-5�c���|�X���Nj�m@*/����ӆJ�Gc��G.��[Rdļ�ԝ�fR�KCE��Vw�^(�[o��sjgh�2��*\�\��ss�����+j�������ꯪU�g� �6��f�8v�6E�t��z�4�3m�ڿM�.����=��SG�.�&-
�o/�;w�58W��[��٦y|՜�C���0�כ�)Bc�H4T�Wi�rU��q���=71�3�Q#�c�\�P�-�J�&�Rj�^�;6@���65im�:���K��u�����#g�o���ci6x�����t�}p�9����O�V���񖾑a���=~~=�侏M��kEHeU�y��K�q�V\�=U�Q�>|p��ՇL�x����Fw2l��U�8n�����1�����ոPs}��x�V���KI,���7��Ui:�XUt��\�b���J���{Z�=Xﯶb����ޣ��"�����2���&[9*w\\�;ݮsԞ��LN��;6s{�M�{v��� Fb;�G�y�-�	�����H�I!c�������Xt����eg�6��DĊ�"iL_��t�e� s��F�'�^��#O�C�>��)���о�ChsZ�4[=��9��I��SU��V�^c�-Tȕ(B��54������A6!�]��k��\�r�����V(Q������Ԭ��K�|<����g�rÜ����ZIv��YR�;�߯ʼ��<u���;í�SR禥Nș�\J�E����]}�O_APy��ؠ�+q�غ!�P�b�KI�{6��rv+�|i�*k�@��p��~��;3��w3s|�,#��!^0�;;����_>2���|~τ"Ķ/G�*�:��|��ʸk�8�A|~Yǆ�	hL���o���)�\�Q]}1�9�J�^w#P������V$a�!u��6�f\r���e	Xz��v�wW��}���c&��e�pU��,W+<�iF�>�i):�6m�S�t�B��I��x]�34�3`��\gvl��/�Wj�!��*k�4a����1�Ԃ��C{0��H-;9NǬ����_%z	�xB� N(��|\5p6���n�2���{�lsؓ sw8s쫧��0�ְ�,�<�	�,�$�u]�~��3z�!��8�ml�QQ����i�B���p���(�m���!����yEl�9]ѐ-��r�u֢͏)`�!^��*��{�#N�ӫ�Q�bV��Xm�^۩�M��.��2��:��pw�N,�ot�]ua)�gXv���� CksOf��2��fi�\U�MB�v�V���~E���k�V�%k�[]\g�;4��\�gCݽ���(Xm�:x�*�Ur6%cK^�
Ͷ��4��5j�rp�J����b�fn:�����w���K�)[�n��9Y�k�G6�jF���r���6~B��E|U�z`�|iNC���E���0�J��#��7Ju�S�#u�v}��x;f�S9���m�r�\��3v��֣�s7F�X'f��84=��Qvn?X+��FC�����vsfr�C3�u����m��.���ws2�lH�6��w��N��c��Ƕt�nQ�7�$>���[�(�2^f��n1r�eYŵu+-�x!1]�g3���w��=����N.=J�`CfV�q��"]nW#Ҷ��Lʱu�c�����>-!K���{�i��w*f�T�H��5W���Y`�qs?wf�a-�W'���U�a�Fp����Ԗ�H"d��;h�F���ݗ��3�����ݔ$���@v�������W-��Z[��U���*q�N2�Y��E���T7j�H4u���v�r���K/l�f�1�m�0^&eU��'�2ֱE��5[�G#�Qc���������R�3�k.��&�\�׮��jT��.���Y��,PU5{��f8e�S�.5�_-�9����Jm��(ۭkZ���B�Y�T��L�r�3+8�C���]Z�(ܷ	m�A�����8�2�R��\""�ݹek�B9A)F��ЄHI/����>��Jz����h�7t� v���E�t";�Y�|�hCZ#��{ѹ��?>�=�'�������ȴ��b�o�^��b�]������³^F����bҩ��Jc3h[Y�`C�"І�@	3���o)|��>焟����,�;�V����}{<r��m}�򳓤5����G)�K&�)U{�<Q������|^&x�����ɍ��;)��5�S����Q�)�������;3�&eј��C=)v�r�N
��ޣu���p�_xNxp���@�^!G�`:N��o{՛���\��qq�Μ�p�O�!�Z�L�Y޵�U���'ƍ�����?!G`>xl���i���3~�S�+驹�NX���1���b�]�L7\�!*�|�l���;�ye���$b[�Vn�v��|힛ܔ���f-�v�Wysҹ�<�>d�4��E�/�O�OV����L���`�K��76)2P�,��?����͘��-{P�m;#���9Wӭp���}��bTEjhw��=�=]�GqY��؞�\_��a���z���M�ns&�q�g�z����Ǖ���n�q�� �E����(l�}��A�'D�V�\��ͷ��Ȓ��a�b�Y�B�p�~"-��gql�;�i#���
�4&R��lˍ6&�\�a�8��C������?W�28��c�<��/�����H��NA��:�Y����!�c��!���bg��ʘ1tb}����v'+1Ĵ�U�����^/R�[����Hg�Νho_+,�熾E�rT�^��[���I�Yqv���IX|��Ѝ��x�0�,�c�
�km�0<���j�Xo}��9�W�'��l]��;S�����%�SxI�{N٘&پU��܅�����D���:i��ףz�S �5a�*��O{:!��Ϫ�Iy�����M��-q���P�\�wU��l�����!��R'�UL�F|fyi�_Cܡd<^;���Ҭ����,﹓�cs$=�r���ҋ5Tv�j�\�wi�y�C�G ��~�����T�59� �X������d!��*֘x������Χ��sSe؉M�]�޺�L+�P��	]t�ѺL]Ը��1,xT�%'���6��km��9o�G��X������{���.�B\)�j�n;�֊���ϊ:tñ��n/�ג�ܧ�COh����f�6��eÿY���sλ��5�=��X��C�TG��\���!�1x��{̩r�A�V���Տ���L��������O�}zz>�����{کbC�e�)}"���<D���W��,OHE�Y6KqK2�a���u�x��h<Ce�AE���YF��gu��!Nd�/�C�t�����m�Lj�jᕏ�m8�<K(�=JaI�0&e���&rz&%]�4�����`ov�����B�����ƷT����"˵Z>��%����?�dk��ῲ���	��x��\y#�C�Y�q�U,^���r-զ�!$�S�k%�_/T+!O��y��6_Ts�X�6�L`���4'��y*fD�J3��E�������U��ɭQ��=�&+(�V]���%$a��'M�a��kg�r�:�����ns�LI6�)�+��$�H����Z�8:txR��k܃@V*Ծ#��7��}�B9ضL39h�Ä���oq�1eZ�]�:�s-n�G�/y�݉?��7�	��3P����ȨbU��SMX����*�=�oyL�O����l��gb��n8kˢV�I�h{oݛ��"Y4t��ó_��ƚ=�\��4�*��Ry�߽��W\��$_!Ӟ h���\��W����b�uﷶ����T|1
z��C]������p6;�a���]�I����bpӿ����K��H�D+d��+p{��C�1���qʹ�>焟�����9�����g�;-i�|ozAm}��ü�ì��s���A�&wo�p�i��͑5to��x��Z����~~#�g�/G=d�AF���r���W���:M��O��j0���g�m�e%ZKd�"H���»:����b�խ���ϰ-(����S����Χ��cpJkf�Vb����3�4m��Ξ,��� Ku�&�<�������3�|D�B��Q�����o���8���9\^<h�ZkP�_c�	�y�*�����G���P��
³��y
;
�F*�Κ���{�a�<����b��V����[Hu���*[�Xd�tim�A��n�֡�*hv�ʦW�mW�u]�o�R�:��0���ls킌�� ���n��X����,Q��s?jBE�\&����3X�|Uvu�/ƹ	��T|<���y�B�.����u!�S����m�g�^�;sf"(�`�~Ŧ�u�P*2vz\�ۅ:hNɺp��M3V���l%�pڦ����{n�����mKo
�:�u�nC:f�G����A�9�qo�hҭe���+�[�m���N�ծ�M	���7���������;9��k^V��[�u��yӎyr�\���T�6��3G��p�V~��;���(s���B��1ݰ��p�O	Zl����B*\�Q�eɛ���X���n]Lw&BjX#�O�����:^s� J�����D(U��,���7}�ޞ�K�nں�@j囧oە�@`�4d������6|F-�:���L!�4�ܼv}�҅�5�kU�uw�����⬇��8|F��&�����#�I���}M� ��O;c�� и�D��F$�]�40�,����Q�q�D'O��7R+���� a���I|��L���un}�i2;��+��ㅝx�ˍ��fFS�<F"Y�șj�٭u�+�d]�"�1�.�1x!����px��Rt7��J.��;��s���;{pqi�K4J�N]����V�w.��m��_G��Ƶ��W0Ϛ�Qp2�L�Q�$[�Q�f��P��	K0y2�i�6�a�o[�R_n����W�� �_1�C���zet���o��6C���5����3rg�	�ڃ#P�cˎ�w��G��8���H�<W�n��a���<�a���i�_F#ò�����W$�m���&�qolD�qŇ�0۳�k���M9�Of�篜"�B��}��<��G�1��S�r�9�\�
�3�O_Lr�/P�i|�����6g���scw�^�ѭ�����D��cbp��({�Os3,tU��1��|cM(�󤪦�Q��)��=d�7��_oׅ7;l��\�.V.�ќ�
���Z�)��V�ص`xwj0*�{��;��{�xC��d�u������@�p�j\>�gv�-�0f.����=L��'�����Z�#2��V��p����}�<�!L7�bBE^X~��`��d�\ꎨ{�<t����X�H�L���@�&<���k��K՝����YLy�;5��W��|��	���ȥ��Vf{�,,�Bx.:^�����!��T<Q��xJG�ޛZ�>�D�^X#���'������vsˢ��W�o,�Rdu!�j&;�só_����*`N+ZB�gcD7�0�FK8f!��d�|��gr�G}|���c�vev{�5=�i,7�Α3�&4�6�Ү�7&a.u�ʞ�w��C�·F8;^E���������a���Y1Z�<���V\ݶ�"�kr;���l��zCd�9��/�w�G�b�VA��.�E�W�8�{Z\�{�ËqżC�O����s�"��x��h���o+�&�9a%�Fا�F�^U�n�\?D�+tr��7���x��Cf2C�z^Bo��9��ݔx�|C>7��zcM,�R&�H3J|
��.�hѓM�~����U�����yQyP�
�}EE;3��&B�M�%rl��ϜiY�9�R��a�E� �U�އ�����w��>������0rؼ|h��jw�˙D��5XS�{���V���.���jD;��4`�R-:�������<k���=L'��{���:Eq�Un�&�����
�+�Y��์�3Q�lN:�;�Mɦ�@�ϵl^#�39�Ť���b�kh��x��cIj�k*�]����8.�h��SUk3=����e�ˎ�u /��Ƹ,w�Ԭ�r�M�K���+��V��㭐q��p�A"�q�h�Iv��u(�N6T��1�e*M5��^�(K����r!����.�{^���u����)�ָC*�&峺�\�5����WTeu^�L��S5���`6�L�,��i�G%�@P���]�K�.L��"k6�v����v=���p�ss�{��K.�-�9d˸��(_�Aw�y��Ŝ�(U�Z��Z���w���t��3�f�I}Xm��ovr������|!Sv�&�&�v&ay;Bj;7/���@�S�,^����}�`�]y�Xx��G-p��6'cF�i��d+��5��R�V*m����k!�?��=�0�a��;��$V*򲨧���ʍ�b�Ji�Hd�"�,�h�!˺�L���q�[hT���W$�WM�.|�VJhf;1��4�9�J�q��L�+�V&h޻��R
A�(��w�l<)�UՂ�j�:f�R����uB��F͚�8�Nb-gѲ*�ʻ����i�B��O$Q��.�]Ŗ¸a$�J�`�wN�_Մ��!wP?�증�WW_e,�,� j����yHIH-����wW��	e�b�-��F��/�C:+5�IYn����H�Y󄖩5�2���@�T����w.�"Re��A�b���]��ǒ�ϟ�Tm���n�9.�JY����nem���D�a�(�4�;��i�m�M*8��cu��6�i�i�N��R��j�lEq�,�DSL��p�̦ۦ��%6�EZ̕.�Z���\��rYs��[m�`�)wnPWVoV�!Z�F��&��Km���E7l�E>���󏼪�,���+�e�J��V�2a�is2.T����&3H��t���5q۬��b�6��X�Jn��=v8!km���֦V֊/���fbg�f�e)�G-7�ț���2ݷ:�eekUP��;�eGU̸��ی�|�(*�F6˖�"�H�bD2���Z0S	���wEM����]��R]���{�]�wiᷭ��]���*t}w���F��į�Q���'I�[ݱ���B�΁�(�r�|��y��Y��(��9��]lY�
u.�|h�����'������6l����3]���D0�/��!l!�r
s;҅Y�������u��=��C�����ٳ�Q'��[/κ��HY�1��\k��J��=�#5Cu��8�kӓ�]wn�F�|Ej���G��<����X�ZEר����U����p�0���5Da[��s���,�ܰ�{��Xw�����0�:�<k<2|�Z^/R&��zC��Uvl�`��vxA�����Z㦍�*����5K|�]�v��y}��F3�(�JH1��ǯഠи�ҹx�mH5�~��>K�/��5
�u���F��难�ܡ�
����Q_oΦwm7z{/4��"x�ة/[��^Ý��N}�@��a
�c1de;ȧ[;�qs�Vɱqǁ�q�1=�t��Mmz�U�:������!�����ܧ"ss'���J&_�쌘ݮ��U���m9�w�u"3�C�������k�؄>�x\��7.�Y�ۤűR�E�����_�����q��U�
��K�
��H���\E&7���pO4��W�x�ѐ�ʎ�HY�����{��l�a
}�2Sܽ]e���Lf����;a�Gy]��Ow|k� \=S#(h�v⧭l�%�U2��G�4e�3������NӷҶW�.���JN.R�h;a�{��׷+m��7��=;	-�S*s��*EE�}ﭦ��3.�4����|�	�5������.M俕_n�d���d�.���G�٩�jf���mw�q���^!ȼ�sfv��-`ڦy_��KWMӾFE�5r��x�B��w�;��)�te>�*nj�0�gsc3"��h�38r�D�U�˂V�7<gk �WUu���!�q��7,	����Ey�
��+t��.ؼ�ݑ�6:Z����W+@�����g�.C6"M�[D��J�ԉj�>�B��M�0�t��];�b\���6�<U��x^K��m�h*X��}����;�������|ڝ�eou�w;��)�,{�1;§.L���d�E�D}�^o�T�� ��y
{�Ԅ�S�N��N�{���i�e�YT�l�<k�˞�.��
;!�9��&�7��g��賙Df��ťi�ԎM�)��pc:��	����6.�4���k�o;7&NʥL1Uzb\T�* ��ЮBFF��e�7hj�7;�/)	D!-���e�Ai����L��o�wL�͹�Y�o2�ŉ.;��B��z�\tVC!��W[�I&�{����;v�бY���z�L���wa��@��(�����{�C��{���7��H�����������a��ԩ�*+ɒ4g�q&Ϋf���8����yˢ���3*��lބ�&��d���i	���N1F%���ɺӦ��� É��9�+��do#Cb�x6pU��n��bX�V-��r�ޘ�ÁV���j잩E۰�buP����QV��4篟o%�� ��X���16�s$[|�.Z�~ŷ�3B�{t����g- ��3��r��vпC�q�7���u����9�����מ��U����]=9yk�fB4U�R~�5=�X8x��M�Z��3�/&��H�U��;1�J��n"ݘ���u�Yu�} ��nMX��f������Vq�|7�E�wWGr�s<N�������^�{�����&׼qT���o�q���j���a]{q�]� %�cC�r�LR�u����n��"�t]
��m�t�t��Y��&0��!��8��]ͦsi_B�c`A�1�5ׄL]]�4�s���z�r�~�wy�:	�>�J�Ev� y�g-�N:v>'���	���bV��^�)6�3Y)xjuSF�����/�r���X�ơ�j��7�Rq�1���A��j���$�X�U���\����	°6U�ݽ �w�y��B6X����}Ń���v�n;Ģ5Z�n64�<s0ᶝa�lj%��_ꯁ�vzJc=Y�Q�����M8���e,�'���ލQ���#q����Hn��*�#�1���gi��x��]KEΜ��f�Y����{�xp��W�r�j�q<��[w�9&��U88\B5�	�Y�*��zrE�ٝ+�G�J�z�O�`�boy�1<��p�E'�7(���Pn�*�5�e�1A�ǩ���e�1}����H�y��9m%�ȵ�[{�lF`b7!� �Q�W�-ټ<ʋpqe;���k޲z���̐���ѩ��hZh��1Uj�j:�v/Z^�ݛ{��YՓ��X��"���D�f-�*L^�5x�8R���lZ���#�ﰔ_Oz�-��B�}d��ȼ>�$U��x�(;��)�����z�j�+U�n�ݽf�)3d�k6;^�<��{B�ΒOo��V/*��7�s=���ִ0Z��M���������:q�hɸ����c1v$sm�`V�Q������<�w]�K�|:�R�qb���[V4%�F�T�'�/Wwl>d3�[�Ll��w�:fv.̚2,����{�j�@�n�Cm{ݱ��\���Y)j�Њ�~�2�NƊ�ӥ�~�ȓ���yt�u��U\O)Xz��Θ�a0�7QY��N��x+�s�1E]�7ʲ�#���WT�N�z0�9H�1��W�a-�=�_�>z�ƹqO�D.�%�wQ}�K���� ����]�w�/:9�c���a�/QZ��fD[#�kc��m8�x����8�ߜ#=�;���Ov~�<�
UrPpJNo36���g���xs���s���e����7�≴(��Me��xa�3P���Dr&�8��'M���U�v�M���f8�X��Iв�m3���@��]u՛�8kU�� %��8(��<�Wk�c:�׼��z����Y���� �u�}騫���k�#fݮ�$���˶Q����a����GI�:o]���=���Wr�gۢ���9X7o��:��)b�ށ�ځM}	��:�Ƒ��^�iÚ��b�j-~�#1��V��m��
��>�E$Xgq�V)܌Wd�k��@%;�wN@Gm�rj8.��Z�SUW{:u&U����T#�`�l��x�PuȖQN٪��H|�lVzj����sSԝ���bc�`˧0�H��ڐ�f�16oΥm>�.ԵP.w�[�u�S�e���Z#h^t6`A05D�:N�Ԓ'Y��ec����^����O�!�q��l�7�;s�N�a<�n�M�x��=yӆ=�G)A����js��zٺ�r�mm@��و�2�U$ϵ�̙�]h�nHE�W�.#A�t-n(��#�Y��w�����؛r��X�1LX����<w��3��t@��JԮ� tq��Y/+Ӎ3�(r��B(��7.�o_�¶��/c���.��F��9}0�$:���mC�/�]�O�+���c��-���X�ڵY|�tf�>xX���+o��K����2�5�:��ft��Q��j���f���<p}SM�y9&�e%�8�
)����]�`���)*z�vީ�1˹N[�t��Ϭ�THum�s+)�"_ ����`��w9^YB��G�Q���wOv�oud���)�G�|���of�U��6�;/�a�Owqf�S��\il�l)0A�[�{�w0��'�.������JȺ@�7�S�P�|��$�q6�;4n9T̒J&�x�YN�1N�lܒ
l�~3$H3v�V�Wq7�#S�ŗ��C%d�q����ʦ#��̔oY�+*%Rb̼2"��TC��Ihf]K���I�,��m,���9KĆKB̶�ٷQ��[��(,t	�J%�7�Q� �R/1�p��ǔ���K�-Q�Y��vq8��3(�ڣXe�b�F�5�uvI���u�E(.�H����P��f�J�)$b��՚��V]�I��&<h�0��M��g3ElY��0L��g�s��/X!:�027-c7�
8�  
�;�Ͱ�Y�n�j��Q��"!R����1����l�i�-������@]��0|,�m�L�nVUJ�Y(�-��Z��̻�k��>n������1պ�(�ƌ�k�bܢ�Ӵ��sF���ښPĩUv�q*1Qb��Uq�6��2�cF�����[��j�]��q,r�j�̕����T��j��a�-�`��
T�e3�2�-h(��T���2Ʒ.��]v�s���0fQB��3O�uJ;���S1*ZZ�m*�	m�-�� +iWvz��°uh��%V�(�Ll���w��*��,��Tm�\�0����Xy��n���n48ٜ��&�NV�[9�j�����)'�Y��9w������tT.����kX��n�w�[{���']�7p`��Г]̳
��X�-�]A�Y0�E@ه�5���������Ŗy��j���dm�t�v˲5�\��}lt>�8�¹Ew	�,����Æ��21��z�$��f��-�S�fƘ�ў�~#�Sʐ煼�^Q��xJ�b�s����zwFh�F�j'b�F�dk	�cU��%�N��?`�8h��̛�7.pZ�뉡�#y�
�Hv�i.�VܝuɖѶ��[����23��ƙ�5x12��I��xoL�xVl�Z ��Y}t�� �Lgd������f��(wR|�f�ٰH��G�&굹/{e-�x#{��c7��B�v�L�����a��qn�E�۾�3ۥ2�_G�;/��#��{�û�I�"�� �����0��zB1N�>{�o*����.�~��z֮�&��n����kZcc���n	�vs<� k_n�ŭ�l���3�km�es�Cq�L2��w��kn:,� 2����N�e*ɓ�>�3�
��5cBt��9N+���ɯw>h���J�w׵[]���gfl��lqA����39�v��n�������靇�p���^2��:�舺��I�-|l�HC4�\ F\�a�z���`$Kƹ��/t�'f���},��s6l`L�N�XF�bҳ@�ʶ0Y9���H)l?R��cf4ْ�X�=�ײ�iP�4�BqW��5W�N;=;x#荍����%�<_̨�7�/:]�J4�"��z�@&^�WU�̋}�<��7�c��1���c!���I�ƶ���{^q�36�u�-����#	�a-55x�OV���O9k2z���y�^z�6���2�h�X���v��r��t��d{{�p.����dʱ��4`��r����^�"a�V���AS�S�L�|�5G�k��G���4�$��=�Z����u�>��"W���t�E�8k���_̱�g��Kµ:SF��^��1��~�n,8�z/k:L�i�|��b���H�!�{!���]9�;��Б�5��K4*��@sN�_�J]�:���Wx�m�����/��;o��Eo1�����S�\�~�Ks�6�������n ��of	���\<T2j�]���ki8n��,E4x��0��Ż����ݖ��h#Y���N�Ķ�F�'���̭�5�<D�[�f��;��P�v,��9�V2[��.��Q|�V�z$J�����鮮�Y���.p9P��ݽ���܁*��y>U=���\����9�7K3/x �k�,��ã��2�cSE��d,[K���e;�m������#<k�.Z�(��"2�����f+cfa�D��A��,B��2�聵1��k�͞�oa5Ū�M ���zǴ�ßIʅڷ )x�Иp^���gQ��Y���"ђAHqu��,�DZK�&!����1VPkt��������2��W���ir�f�.o� �w��d7u�ka��fFw4���l&(��x<�¦�(�5����K�blv�)�N��{��>}W����﹮�0s��u��(�ȲA�w"����!k����8��/�y�T!\6��UB�E�ôZ��ռ֬O�$�]h��і�Ekյ�6�͜�'��,c���%`?C�TG�VgD�93�^<�A5�M��gWa��\�+t���Z�E����XX�N���	����Y�n5t1ib�lR���;��7ya�9۪��KTTt
�+�+�ci��ʙ]5�<���ZyǏ8��$��YȔ]c'<M=%�X�n���0)�<S}6�K=���ȶ��YKv&댵8t�����`���p�	C����l��B��pw�6�}�:��0L�y���u}E�R%����W�3n��Se{e�񉍧|+V۽{h�������"�h���@�����X���e���x��6��v⯠���PKi=i�cFjDb���$M�ְ<�Y�냣��H��#8u��T	���> �oX�q;��GcԐ�#z��˥��+Uk���
�U��iH�
|AZ�z���U@/�Z�R���%��η���Y�17��=�_v�*kV7w-�tQL��y�4-q�2ƛ�����m�&�Rg'�ĺ/�˫�hkڃPƄj�M�XR����/�x��s��S��q�f��҂��ܹ�G������}.c�
Ѣ�-JV���.vI�pV��*NJO�MqzTK��0�wu>ȗd8?�}�Wvp��ʇ\�D�n*y�����q�v�a}����f�>u(s��À���9]��?!<�y�c����櫙�h�t�ִQ\D#����~[�h�6�켚%��� �����}��l�>�3�['8Z��^W
[=��]�w֊a�B�q�������v�س��v�2o�h~�r��l)HOoܗd�B1e�9|��>ٴ�B�KFIέB�ؐnF8;N�͓5�q﷖�oڰճ,,H�O?Y��0�k����7������vz�S��z=[�Q)���{�p�����!�8w���K�O\dz�%�]d2�:��ɻ�
%�N����;�p�t#`��v�n�Uu@c�{�h�
tJ��9��maY^���F�<�o�u�5���0.����طiL��	J�<�q�����]�mȃj�\'�;��{w6͡з��[+�s��y�����vhL��тe������0*Ls[�� W�|5��gȼ�4�k\+ˁU#cY� m6_7Eb�X�PzJ
�>B$�P�_,�b��P������X8�(=�����ӿxw>K>���z����3�K�ӽ�#�"�Ph�����G�{�Q0��ۛ������w��q+�(�I��45��e�]��F��γ�L"�+�7ܚ®,Yu��k}����v\�'�J)�و�#�Z���	��w���A��1 �'��)hp�GnTP�n��4[�v�E�����*��Ȯ��Ѹ��󷙥��[7ۊ�n�D`�'����;�����������E�U&ӎx�ԛ��}�j����Sz��bԘ��D6K���&�p����ܱ�8�ۡ�B?g��Ԝz��])(;�X]��/4�����X�%ֲEw7�Wr�Y�A�̸�0lu��9�����H�X��..	k�H��������k��+�	3 ��2;7��DŜ�;��Y�R�^N���t����DV�Ar-�_�H�((��"�ws)&l�g�����+��Ki���
6�I�"��L�:�1���a��lU*�\�T�o]J��fLbp�q�е���f=}�+��_U�9�-0�-��G2�goVf�:��Q��5�
�l�2�KB��= 5���O���ə���7�>�35�a���.w
�����.������A�7]z���E�zF��wp���C����ilג���n�W�vIlz��[��ȼ�$緤Z�:�7���ed8�V��:�T���c��dp�������K��:V��E�h ���m����C�*��)�YKo�	�V�LR6Z�k�ڨ�i��j;�̅�"e�# Ö�Y���8���5�Ƒy�LU|��`U�@[�x0\ɗK���c����1�U&�;�2VQ#SY"�#3�5*�]:�(�T�+�-42�3���CiЬ&SZ$x�B)Q#/U��J�a��2۬����ғkh��
��j�-R����-'jTUU��ą�\�X�U�L�
Ŗ�J?G��mˆ����FS�yД��U�m]ET�V�bK�m^&�bt.�Ȉx#�jQ7k]��m6Re�֚,��Om��.m�imZ�TAU_��3	�M%�֥�U��Z���j(�+4ԭ�0�Tt�QDPE4��cs"��{n�eLƦ3�������kZ�e����*�ieJ��q��y��F~�4�7�b���E[q�ӫk
Zb�kXbi,EB��U]6��8�L4e��E��,=�l,G�]�6�j2U�[m��q0�Uu`UF�Gv��v�eQVƥ�%��m�5t�z�ޮ#j�jQ�Xƶ1Z-(�YAE-�CwZ�b�������e�c���b)˧l�YF�UZ��K�xf[M�n
�~AE��������g��}��]�R7�9vCt:���[y�8�u���`�;��^�Jk�DW����6y+�����;y3['X,��}�BTR���4ߢ
��͏d�逮��kQ�\��T�@�,a����K�q�⮽��8X���Q����I2�2d?�6�Xh��VU��Ѓm���sbV�Q�"�׸����w`�z�Æ%0n��.� �y[}�l������2��ά8��X���I��E��6P�Ɩ�O`ˡ{�]u��	-�V�9����8��1��֎��y��Q�e=�s��F�Y.��Ըd���������p��� �Z���C�d���@�풎l�6�s�JI�5�c�_��v��.ӭ��a9҇�rܚ�I�o���6�0����4�@ѝ�?#7Z���fo�����n1���ִ�`�z*�]�-��{��}�,�w��/2��;X2�����m����xlg*���:+8��xs4`qIH;uIVS&�|��k2��y�B>��w�tsx��@R�jV��i �Dj���U��C�tK0x�U��GH-�:���[f���=c���Ogf����\sw�'/�Wln��;��%��M�-6��-��ޫ&�Ut%ǝݕ���{^���V���Ê ��pVr��x��F�3���K9�>�DO�m���k���ol�Uu���b���)���%x�]�9>>��ɺ�'GhN�307�,�����K,�>!��S�=�@��U�}����ѝ!�M�49�o�UY�[��q��J+�	Gm���Vbz��:L�C2�jd;��eeѲ�N5�#�Ak}~�a����t��s�z]�HRmc�!��DO+lJ�9)����ף��IwpuH7<[�#̀=]s�S7�|u�R�b@}������U���U����:��]s�X\�')�mk�q�J<�ZN�&�Γ�;���/e����zvj���KJPIK :
�4ej'�=�^�ԋ}�jt��/��l3!�ӎ��dΥ/�Fk�%EwG8�7���X��i,޼�<�`��B�N�)W��F��69e	yǵ��� ���|͇�Ɏ�YӀm�R��)��k�G����n�ׁ�"��19=�n:���w�z�����r3a�Yl�uR�ʏTmZ�5�'OL��D��C���;7�h�&��"�Q�ĥ������r���U#�u]Z�A�����O�[*l�j#��=���x:� ���DutZ}�:a"R�3B��B����j�.��muJ=y�,l_(	
k���R�9
�Z5�vO;�������ԟ�?VUQ�v2��]�twzq� >k�X�/`,���� �:*��! �p�T^+�{f��`t#��곣�M�\CA�P�	��yI��g�F��y|�=L�r9�DQ�O�]�E�䪻��m��~�`��qU`���ɪ�"�%͙���-E��a����n������b���p�	�⸳s���)C,��"eQ�y&;N�F����yow�xݬڅ⪇�tE��.��t}�S�`V�̼~��y�E�ъ��_�G){f��b3u��J1�x�S@}[�TS�蕊�K�Ѵ�Q�`Y�����m�I��t�["��N��J����f�j��8�ĭ���\�L����?}�Ro��?�Ev��k"�d�fm�U�ڐ�����냋3��ud}y�4pO�c��3.��(=Q}�!�"9�ԇ�P3�NNR�T/��
n�����M��<9�K���@�b���3�u�����ա!eo0���=��ʼQ���PS�}ťs[�O旇�_����*0�^3|�&��oU��� �b;A��A�s�`N��r!".ۥҰ�۔y�e�=�-8����Cy�پ���Q�X��
Yb�T������v4UA5ں�f�����9	ƾ�5��}앂u�GV�� E8tY0�o\wu|�hd`��y��ᘠt�(SÛ�z.g��g(I�ل۝ֵ4��x�9pI1|0#����2q� 	$C��^)Фh�V,��d���D��i�ڣ��C�Y�Y��[ҟ���a��\+Jr�ݓyMԟ X��.�y37��S_N��x�!�4L�:Rx�'���Ef�;���_pW��^~���n�qM�w��`�<�k4b�.��,K�Z)��Y����?:k�G+V���l1�"�ͫ%u��h+[���.{S��rN[+�W��J�t� �t�Zo"PRա5���wl��1�'��U����}�K�WB$���ue)���d&��+���Q�z����>{��oW&�Fc�w��@�����r$�$��*a�4LVز�eu��!�dm9[��[Qp¯wG,;�f݆wh_C��C��YM���[|�0a��������v���q6`Q�c,�؀�T��al��� K��ܴp�~�f��3�� u�H���H�y������x�R�ld����p&ߝQ�����ѯ��L�OI�7�[��L٤����Sܣ���+�l�_pW/LUTM��!$�^"�cW�L�N����+���N�trn�M ��,jub�njH��k��d����Q��������%FՇ��	8�C(Pc��1�����]�@A�����8� �ʡm��6�
�{NҶ�1�(賨��F�L�	�v�����^U�jG �	L�6���7�����|��8����:jpp��&P��R:*����z�4*���՝�&W0��'���ym��P�{H�l��QADh�(�[��;u��Q^����)��:R}g~<A��x��_���!�NDgr�D3�H�m
�]3!vݽ��r�K��*e��;n�&:צ�M��ݷr����ޡ3B#+�D�`�ޥ��#p�	o>�UN������������r޲�O%��������������ZoSQ,u���6Mz;��f���[��.f���;��&8B��{�[0���@YȬ�m$�ˀhs�dZT��y;�/jGD�i%6��p7�z5]�'Q�O51�2�i��Ta����ֳ	LӠr��=�Ɣ��jE5�6�jDmt�T�O�ԸL��:�*z�c8c�E+����� vΫӃ�<��QS���9���b6epɺO�#̜Q�Y4T�y-����%ۺ���w@5�]:���\�5�T��do.B=��h��0.����w}�4��[�o2�:.G��<HjS�&��	<0O����Ґ�Y�ʢ��j���燮�hUk�n�y�m�3\ ����/*�k�h�][[��cn���v�H��tk�����L�fE�)a3��N�8��:��3�v��;s�Za󼙭ˊ7�t�E��7\�.��7�9����$�ؓ<X��q�w)���.�>�����v=�ftDgD��/֪����ɩ�ox��\q�λສ�X*���c�����z�S��,�Uf�.]\�S�K��voM�u|�����.BJ8o��5��\md��p�,ugm���i���j̺Ӫ*��&MS�)3:�m�̇��	�G:Mb�2���h�I$�I$�pB3"��R�l|�i�	�s.iX���;�6�+Xf�kE�p�<H'���YX�S�E��'3�H'��|Y}u-}\�C�ݠ�a�=Z�V��gsr�d�������'����^����cڣG�S�	g=ߣ����Q�!z4lhWSi�}7R�k���w]��M�5;��iXP��f�o��ϳZ�b�|��j���?�n賈��Xϥ�h�˦�d�.|,�����&u��G\����#1�qCy�˞u1ˋ���X8q�GX��<��Y�\�29�n����8b����Om���|:q[G�uPw9|��+�lé`JI�
�ìH�w�YNa����Pb�u���jJ�q�/���E)�RKJ�\�	�Q>�1>��U�dS��c��{v����Q]Z��j�1Ur�V2�,jUD+Ki����g;E`�t㥈�4b�*���SDb��U�%�%�QA��^aX�
n�+7j�[1�J��[֔V(k3!�0��<¸[�+�T`��h�m��1���1U�SIX*�\q�Qv��33;MH�R��E[J*&����X��*m**��"����یm�T-eKe�&:Ѭ�(�Ӥ��n5�c���ڱӘ�ʔF� ���lU�n���ox���q�Wj�:f��Q
�5f�B�4�ut�l�4ʂ���1��F<����Q��+��I|�3g���=�a�7�;��X�f��@���ڻ$�,���#;��w�ދ���hmΥ�C5�*ދ�36��n,ч�'�kreW�ne ~s{�_�#ذhCϠV�*��ݍP:�b��~|��ZX}2�̮[��y�b���sp��^�8��z�y�^�Ҏ�/h�e���f�����02�S2�Y v�}ܲP�{#Z�3k�13�v�y�M����n.~䍍X3 ����=��X��.徊�Z�X�]��z�2��(� ��V?Y�Ί�O{�Xuqh�.���>��ʻ��L��t�N�')�Q5u-U�^��ybt��~MY����=��9��}�ۻv�@���d���+�E����7`�c���ջ�k=����T��F��ؘ�m�Ϥ�of�R+0����
m.�95]��ڳ*.��>Oe�Հ�nM��^}:9�Vdo^d%��^�tI�\�iu��j�D��hV#�U)��'U6�BIY���[Z�-�*(��q5�v��Ú8��E�W[��	�ȉf�Z�x����38	ULL6.��c��V�VΪ&Z잆�(Ӆv�Ͱ�mc,1�	��fw����Q�yX�݋�<��A��Cn���`^ߞYUqd�\$�8w��iBM���U;���g��W|�;J���om����u&{,vUnO	b�=#w���-��~��J�%aA�c�=���Ƃ�N��8���A��i�DLȦo��֊pA�s&�����i��b�\�K(��}��=PpZ1U�������%Ӛ��2uH,Tm��6�Հ��I|�^AvF�W2Go�d	�v�|:��JgR䫜n-�Y���:���fS��..�^8B�V\`X�6
˲�tW^�z}�+����E���XCX��{%I�j�Q^c�u���q3�q]^�Z`V7j�������+����a���N�<���3w��ٞ*,����]օǃ����GiK��嬓����TFgXH���z�p�[�g7%/��M<�%`^��`��S kV�N#��9&ga��.�{�D�1B"0Q2r@;��`��X�������NB���F٨B�� �bf��L��ʊ�7���@IGh���B�XEuBGQ��ZKk6g�y�O��8Q'v��Ĩ`����u�@�=��;t&���͜�=�^�}TtB}�pɭ��)��]p���	�IX�v���_m�6S����� i8Σz�G����@���s�!�7���Tݎ�h����Jc)�TΤ2�ˑ2��$�� 2:�+����m�(�#��r�r��k�9�dv��,=��V�w[���ۊ饣����f%��0�HP�ĕ��]�y�y�Q�c�H��H1]�<��לYMPO}�z�����D��C%3��bVF
�����	�7G���Nݾ	+���l<���(��x����ٖ�.�3Ɏ��R!\P0#��M�p��$��/2{cz)�3��C&�wX� �����g������� �kR�e���26�����} d�.{P�v&Ɯ��vv,��tǵ�%�e���v*�wΩDVo�_]�f0jD��;pU�J�69��m�3��j�s�V�e���7#���x^r�o��/�b�&�V�����c�SQ�.(��*HksV�n�з����HM�A�\󧙳�ؽ�7��Mg��%�u;�Eڎp4R�ԹL|ٙ�%�����d�!ZFtSӽ���S���ӭ=��&��&:��`%�+c�_J�Z�-�h'��m͞7����Y�B�5~���z򫫧���<!#h���j|.�_���b.�3���]���hGw	�3���*n�S��Q�J�@��1�������i��n�+��R�����yH�Ư���y0��.����T*�{��`�v1����MoٌsK���C�̂��i���׉�;wX�n�gs��Y���'v�q=O2�b����e]P�������)��@	>�1�O6lyѬ���w���P� W��9r�ڻ�4�e�kd_����P9�p𒛮�A�6�v�&m:����a���-�q9�
%��`�oN��u��E�s�Y�K},��zpB��w�"���|k]܍��:�$�\<VMB��Cřxa~S��,�]hce?z����Ů�ۆ.�e���h��T�����u���g�0���#�ʮp����J0�8)A/z���Ah�@g0��]��/�����'(��K���wen;/��]����՛�0��*"�=|�}3��U��U��v�ۅ�Y�no0$�vQ��R�Y�ۯ]�B1�l�U������!����j�f*���ñ�vs�tR��8�N&lz�u�7�`��t��b����CS����ץ$�p�0�T�=���0k��d��b��\�a&4����yV.�ֿ�;�NPq;��~9�U��#�+�%,]�W*R�df�Y�.�Gh�˱���]���b0Uv�zc�*�#ޓ"}� �g����2�f���IY;;�����C���5C�mT�$�ks����fT\�'�ٶ(������Y��f*��<�_��Ƥ)���-�ub�
Mw=�1;s�����ũ��HT��B���;$m�}�7̵7^��w�����s�,����Y� *W����u���
%~+Zډ�cBDh�u'la�<����Q��}K�#�a�1��j��>��dKx�͍��y+���)���"�=�k�湬T���V��̇�"86�����ۤl�͘�f�8X���Wh�Z�xu��,J<�!�Q]K�$脾˞��3��&QT] ����n��zǮ��6
?^��li�'�h��	�g���uE]�Wc�͇E3۠�{#*iv �ɱi����K%��{��y�Ǣ�c!�Y����4��]�̋}}Y��M�U\���K*.U�@�;wmت�����mb���r.Yط=�s]y�O�hl�gX�@�\q��j���`ų��vA�\)�F>s��nUl�.B���Y��#E+yB�Ix�+�:�_�qˍ� �X��u�,�!��o5�+i���Ί�V��W.�>�+{��CƩey��H�r>��M��U�[�������ȹZs3�����G��\G�ELDDDw$J�(��:�� �p˒�(��Y<�����J0͉g�,��z���k��LĄ *��Q@�	! �����^��A<p�SHE�4�<e�m���,�Ή�vRDDA�2���N辻g��sMz)����R(oXiYq�����$0�)�-K�F�Е��p�p�@�GG�疚���� ��x���0��((��&�bV�#?��M���/��=��fO��c��8}���O1��r�(���	�Q��Dva�!h)n!B�S%����)#��R�޵	��]m�q�ݴ�"cUy�����r� �eh�\�;*zir�
��,�"�@L��D@9Xd�6�8B�)��n,���L�� QKu/;���ו���j}���#��\�����X���U������O۶���)4�e@@�S.�b��<SU���8��+'�w�4t,�.��O_e�:^$E�j�����;�SJe�yw.Ø�(��8�;������6Lql�B ��M���(� Y�=J ���4`�-��$Į�r|	�P�r1,)����5PA@�\�H��F�l�����QDalH���w��a��E4/I��RD`�`�4B���!�$�e�kƁ!�*
 d�:w�GfJ�M� �W��م#[խ�G�H��4m4��4����AN|�����q_6|����;�;M�O��&_�� Q��v�a�6��w� �}��G�@@��_��Z$�2ۙ�y�t&��������7�`�qb�\� ��H�<�@۹y����02!��7Dw�=�40r��F��U�D\�lr
o�1MSƥ��H5��چ�ވ$�L�p��İTYJY^��d	  ����4�Awǋ��lp��@�;�I� .�p��F���\HB�S�G���t�A� ��J��Ҏ{\�.�p�!U#�