BZh91AY&SYπ/9ת_�`qg�����*?���b_��p                                      4(�L� �*  @�       P        @�  (   
 
�  ,�ȩT%T�%BR�$�	U���%D�AT�!E"PJR���
�%RB�*�@)J��J�� ��BD�@�*TUI(�
IHiM��*�b�3i6������T��0b+wu��H[���:wIw9e�h� O}{4  �� !݀�:' n����v q� w* 8 $9 R� {�y �@ ����J���� R��J��B"���| a�� ����y <�z����'�k_}����}��^G�����R� ma�z���!@�j�	[�d �t|���� � 2=<�@�`=� y�;� <{� �^ �����v u{� �� PgЀ ��(�%�D��$_ �|{ 9ˠr 9��` <���U^��=t �Xw��lrh
:�� n�z<��=��  � _x�� ����@+��E`M����·�U�8��� =�H8 b8�Ы��J���^�{� B� 
   w�EIA)(H�<���ӽ����{:�{� 8gPR8 2u =[��ru� {��� ��� �{-�N� @<�� ݃�z'�P"� �8������:UE����tD1h(��Q@ �� 
ԨH���HR�
 �P7gS���wp9DYʕS#@;�ur"wa�KuAR�JC�
 ��U�� z2��	����jT��t�պ .t�;���݇[�u!�c��>�    �?MhT�T`     &O�Ĕ�%F0&L ��&�LD�2�Rf�( d�     4�*D�QJ�Md�d �)$�*0�0F24��b`�F�$I��4�Jzh4)䍩���i�<)��C�����_ٯ�o_Cmh*���κ!�N97z8����AEz5�QQ[QDAS����O�?��TV��¿q��������O��������T�O�X(*+�c��H�("����w��!~�
�h��AZ"D6ІC;a�p&`��C��ІИІ��hv4;�C�� !���M�&��m`�6��	��BBC���И��hLhq�&2 B!�M�&���C�!�pC�#�p!�cC�4&�!�DB�����T(��A"�%B�"�DAP�((�T(�QP�0C�l���Lc@@J"��B��DP��DUaQ(���AC;c &�&�**� (�
�E�
�QF� $"�EEh���@(�
�U�(�Q !�6ІЛhpB`Gm����8�mƄ�BcC��1��Ё�B ��(���A�?-�/����s��[�*	a�6��)�w��=�e@f�����a�g��,8��ѻ�^�n	�o��_�w�����6a�F�ߵdC(rF��y��|�gU܍�3ͻ���kP�>Ql�os�9��}ػ�	��y�8��f]+ag:(-�';*�=݃�a�Uؖ���E������O{.���jos#��E�����os~<8�Uy�Nɰ0�yV �z���Q�x.����Sb�k(�V^����X'H%2�Wq,��ۊ��N5�o."躪���qۥn���_6��C�e��d�v��gP����bsM�m�A@^R̊�N��؁���Y5 ���V��b�V�e��Աe��y�{qeB��;	�pP�d�Pk���"7��ŝ�y���[��s�7�J��6tX�'�C�E�Y���/J�.���;^-z��1-5j����9܃q���+7%:�¬{�:��K�>3Iв���4��;���7�,ʛ��W��j5��x\�q��479oN���Aod#��-=��ޣ�a��Hc�n�A�p՛�0��#j�jǽ�M��-��V5�q�`���I���pK1��Ōtٖ�}7@���8)��Qݧ$÷@�7EZ�@	�^I�4��B3�9�� �˗��h2`8Ns휦�x�iC��I��E��GE�C�y�]\Y���OF�y;�Đ?><�͈-F��-b#ř�Ï�~gڧ(��� ����{�l�zt]��d�L�ݚ��,[�	;�B����	��"�y^��wN;X��K����ˆn��QYˍ)���"̱b!�;ؔ�&���+e�0��k����L�ݽzn�滞Ӆ����Z�$�[�j���μ�ճ��������wY�z-�Y�swz��8D��h"�1��c'�v.�6��S���f�'q�g;�l��1i@���^�_�W�6��dzݖ�0J�g;�$���9j�}�O�C�p���9Azo7�Wh�Xu�$�^�e�Û�B�̈9�C����C;!�_f�{��k�g�FO����lA�0!��F����!ۻ�݅�^]v]լ-�� �F���w1
��]��]oOs85L��Fm
�D.�v��!���tm�1�u��i�N$u�-�|)+�o2��n�ID�.&���h����������qb���+A�!��v��~���Ѫ����7S�5�y$T��h��}��;�F嗳`౩��X�ݠ�Y�u��jP��X1�����ev�	����88���D`�P�N�e@�{�Q��V���t���g 4!5&����ǽo&%�Ћ ʋ;DY�Am�Ѭ�Jcn\��BZ�6. �yot�� ogp{ۅ{�{v�93gEi5wq�X�f��]ɝ���WB9k���e���-���2�����Ƕ�:]ޡ�=^嚙�`�y�ܠ��Y����ܒy���Z�V�ٱ���M�#y������Vn��+�M��'D����m�.��3���� cу��҉�۬N����&�z�w�u��a<5n\	jBڳA����s��h5�zZ2,��M&�4��H$�Z�;r �����L�BQ���=�(O�Ѳ٬s�8v�?��JW/u.�^��ح٢�7/ߩ9�3�9!gv�I�,�.��Z�t}iMv�T6�|@ձ���6@��8���^��v
E�)���@|��t]$��pQݚ��O7*Q���9���bn��,�^͙s�p�wNjS!:�]��6cEÇ:�]Y��i	�C�9����H�����;�7/Dz��]��75a�HWÁ�,�=P_	<��ī�վ:��=�}ƫ�UΚ�1���6`k#�I��k���H�9w��\���|��W>s�]/����r�m;�v��u�����i�R˂,R�KdQ�U8�[�����������<Y]ڪ����c�vZ���VY��8�ֻ�7>�Yкz1µ��4�2�p�]��r.��=��������7��U�9�IwK��DVv���K;����V��ǳf)R���97��:�<hN qմ�$a(+�#����̌�BpfR�߮���쒓�v�]����AmŤ(1^Չ �J��9�Ų\� �ppwO�``S�h�ދ;Y�X��%m��D���'6ۜ�R�-]�Tg�`�=(��|�h;6�h�lY>d��p�$n����u�dv��joPr��pp�Fh�]䣙9>P-�\����!�dÄo'�A��2wi�ؐ�m��*V�o%R�[9��%�Xjgw!]�tOsS���⬦�c��������OԖVS0R�I�����Ɩj|����^�Zn��D�D�L�GH&�k8�i��ɒ�����o�ӟ>X�w��n�Ё(�E���p����k�ϣ�T�Ů4���0���:5r黼��X�R!��#��y�ri��z��N�ӆ�^��6��2;�㧪����Nn����3� <�2U6�!��M��2���+�_՘�1.�E��ߡC4��{�prh�/v��x7J�����t0l�3��n��(&���K��U�r��L�k#u����Oai��wi������rɆǥ��G�Q-Y�M�/�[r���Ö착g]�Y#�7/+ꤝ9̎ۂ��;�*��v���v���X�䊓��ņ�9���|4��t�ov��̋Z�/�2IφFW'��ur|����H��7���Ee�Fmk��x+4� \3^�"fT5��_,SF��Y{;uG͊)�=I���r���s�n)��|�dgN����VA��?��1ۃ�æL�K+B8d��rN`;�f���l��p����[�B� �:�Ugq�;#Ը���v�μ��é��L<s`��U��q�Ў�!�iBi<giA�/�	�;LJP�v�y`�QǴk��C�s�1H��4ar��
I`7m��V���_f�N�L�.�+�&Ϻq����"o&n���x1i5��N�^[y�T63eY���j`�gu�%����q���jF�_F�\�-�s`<VL�-͘5�.�F�vGv[Feef�WN{��̙0,qb�m�x�ݜ1���f��.57Y�F��7��Ճf�t�-�ڱlJm�Y�#Vnj_o<[F�/�]��9� �/n�fi9�ŏB���t�N�M��5ucj��Sɬ��;?�.#��W��k�Oga�$;q�X��nn�޺U�DX{=�gh�#��>�Gj��p�>�.�M�u`���T{�_�oT��ѹ��8���T�z�p.��:�D�O,l��z������e*p��&2�� �N?��S[��\z�ջ�B��<-\YOC��5��<�;8E[��uI��p�zЀ���Ҥ)�W�u��aTJ�9�u��v��M�,�ʳ{wM��	�~�j�S܇J�rɣ5�pU�i*W,Y�J���r|e�㗋�/��M��0q&��_uC�4�Q�㓺ؤou0B�Mc �Ȫ��reef���7F�0`�E��o�ځ7���n�J�mSF18^�v:�K�v�h5�Z�{�S����	5�n٥U�on�>;+[R!smkn��^��;�ڛ�jǽ�Wy 'r.�yn3�E��C�Kwee�Ό�qN�؆=n!�W�$�ɷ@/{2��8��p��6VÈ<�&���N�zT&��bI�4��Nq��@�Ձ-��c�\�Ɲ�E�z���칤
�G�Ä	\����0�O�Q�������&
V(���|�]�r;�]��y�;��x�Lr�.�KU<�r�щ����veZ������˳Jt����p����ϻ ��c��P��p)�[{�t��Մ\]$
���ٝ�rԷ �V�V�����J��XW�n�dÝȊ���4���9��%+��8���)��[0��'1>I�Ӈvl�{��$��;c%*l����Ǔ:]=b�aN7V�J9���FKܷH�QŃ�M��t�m:�;���ˀf��V���l��0�N�
�5��vf\��;�܊1����`�L5e[�Y8<i��n��D�<ut�j����t�+���b�:�w�.����S&ԣ��K�U:�ͪ İ����w����l�M���1Ưr�5����.�*�jزCDW�C�:��⏌�u���x�I��ݱ��\�)7:��'f�u�Ν�j�o&�%X^ܼ��*���><c�H��EH�,Ⱥ'F[���sV�e|R�u���a�w}e�MXF��P��:;�(��
�]LV�g��˴����g#��NrŚzi�\��x��D��BX=�A.�i�0�D@�0��ܿ�Hhiv	�q:	�\��1�:�&pˊ��5v�B;M���Dz�"ȯU�7a �^�w*k7`\ɐJ�jF��
��]_;�(:g3��d�'Cwqwy��]��m�& Jw-��&�2��VsK��U]�_w\ߵ�v0���B�ѿ,��&̉W��Ӱ����X�,�9��~L�2s��1����xϛ��k�!F�5���]�=�A�����wn�'�Mְ��N|��p62�ۋcZe��h�!ܰs�N�h��H:r=@Ȃӣ-]]�Wm/Yޭ^��R�^�ߘ�VB+ȁ���v�L��c�AhU2�Λs��9����O�:-xa�E �01X���9/�ٶ��z����$Aƨ/1��6��Z���Xx�;�oK[�Q�A���p�X��B<}ۅ��["�6�^�Kc�<y��	��qh�
�͛��;U�cj ��sz^Dl��}�$ޮE��g����;{���f�=��2D�W9�;�0�7�q�4O��'GrQ�4t�j��a�7�������x���gY�dz�C����WkT/)�LnX0�on��s��]��d�ږ%�;�����N(�pR���1{���6�W6X���W�&qbg"0��3w;��t�k$���3�\.^��F�$%ږk6k�\�����/J9�$նж�. +��m�q��xP:�o83Dʷ����]�E���ܙ��%dG���������ձr���%��Ve���*#��)���ǯ$hdxc��s�9ɥ�g6�>�C{������W�'�YQ�\�NՇ*sM��گc��xh��=9�U��.�2l��f�Ǽ>W=O�c��Fr�+�Y����9��۳$ZV���T�xkhF�]wP<{
ʲT�Pa0'k�g7�C$��]d,�5��=�9ki��D��T�sK��e��7��]���.��!k�9�:g�s�wNE�h�K�B����R��?qG��ܻ%ô>x�Zq=E���;:3�l���	���f5^5�Hp#����h��&-��yC�UH7\#J�b�p\'d��=j��rYq�+y6.B'������^�v�ƫ�f�c�Б��2�g
{�� ���j�j�t�ʀ|ӯjS@��R�M��oYʽ�{V�v��:��;îU����Ց0�k7bѻǆ�v,CS�����a�Hz�{���H��ב�[&!b8R8D�s�7K[nw4^��,���Bk�y%�c��mq�L�T�۔v� e�S�.��[gd7�^˺N-�]��vuF^f3Sѭhr�ڀ���҆X�G�Ms��u�3U����M!��M�f΍c�z��Fo��R{w{�s��Ƨuݳ��雺�k
��q�W	���n���C�|�,���#hc=�ыf�صe��kf���<e<�;�a8��:��rO�a�m\*���]t�w׹&x�Z+Ǌ@�]�S��M�/[9ecD�<j{�Q&�.^oFni��u#
��jB����I�Yq��I��bpU�FI�X��rS"��1jý�S�ז/�O�����N��K,��9g�����ii��v^���⫚��SW�t���;fHC�j+��J",���w�<hw"�U5�&�@-�ưi{���p���$R��ЗZ�iQjY��O���¶�q����`k�[կv))�-��b�!��x�,�pr�n��:.t��O4�a��r�Z-].M�!=lz�Z�m���X����d�U+	6��`�f�5p������yҍj�׷�]�)����
����噸{��wGP9^�[���lE�7�2u�n]���p���J��(��a��;"Q��Iyi���s��]ذ��;�]U@T��Kt}z+�a�S�|ز���K�9n�sf�i����S�ٳf���<p_!xG����7��R>��U9U �ۇwN0�H�ꋹ#���N'��ٛ�V@��t����,����tލl���ǈ��5���95��0�zF��]sZ{�ES��5��,���twc� �j�}E�hh��z���e���l�e,�O�ғm��Y�M���XD��h�Y.j�d�rN�w C�Mg[;��$�h�26΀���Wc��,[�&������5�obӮ�$�%��������Ż^m�F�vi�@R�v[���jh�p��ǌ�^d�h�8��'�F5�6vI��\��cZݣp�����e�_5Zs:���.=����3Px��.[�0fkzD�g�g�`n����d��Vv�� ���>1I�r���@E��\9� /��|{�죮��Q����4�-�#�2�Q��)���M�[q<8iF��f�L)�g?���i. ,"j8���&�6��� �������c�/�}��8��~PD�@$IA��YEdE�d@�T	$@	T�Ad$	I@I@\�0���l
���
*"�H ��,��Ȋ�
�(�"�(�"��"�"*2�H"�"�(H ��(H �p��`q�.�0���H�� �H����� *ȉ  Ȣ�2
2 �"*�,�"Ƞ� �H��H�2���
� H
2(� H
"�*�ȩ"
��H�I �Ȉ "��)"����2 ���"��*2 �  ������B
� �H(�)�ʏ��jV��Spӛ�5��ҙ��{�Y#�Ub�)>Wɸ���|��Y�����֩�i[6a���/� �ǚ���A�0��Voܞ��1�A�߈��d��8�k-��w'r�����W��|�D@ 5��~�v/�~�Ã��X�+���������g���+��[�|��ٜ�w
����Uc)�=7xw%���b�{8����[��{��"�C���{PS���/�������/�`9z��gznr�3��]�+�w/�t���;9s<�^�����Y��{��nJT�dy�>}ڒ�����F4��˛�O�p���߱6bV���w���c�W�o��N�y�A�|*��|0y�1�a�W�wd�+ս�;9{\lOM㒏#��(}b�qݍ�`�zi7�������O���zj(���WB|l��#2�N����ǻˁ�2�7f#�xќBst�B�o�W��O�s�gI���|/s�^�f⫤��|�{R�qm��(8��i���8v=";~����[���LO��	c&z�L/}��f��蜭߂�3^���η�սx��c���k����ƾ�X%�(�:�s�^������$wLA���ﾓ�N�*��{=�Wrb�����zy��3e~����LE��4�VH��A0���u�)��M�����uk�����y��	|s��)Xs�v��c#j�.'`���'q��z����ڳH����@�{B��oI�ɯޜ�b�����2q���t�dŤ���4E��xXG��8.=	��(�����5i ��|��`G�?,de�T�VPw��?xÂ����ls5l�0cម��xo�w�L��\ĊP`1��0`���0`���`�"B0`��0`��0`�c0`����䦓���ѳ�}���y#���w��+t�f/���~Y�^���.�=/�q��;�}�n�W���{b.є�2u�yޝݞ���	��Z�K����矼��uf��Z�'9�.�����*�5��g��>�oNi%�F"�z��e�:^-�P_Y:h|k�φ�^��-�h�)�ά~��tB��w��&}Ѭ�[�h��(�����{���z{���",^1�.U|���/j=�\��O�.�ӻ��-��ߙ{�y緗B〗�9��S�w%PY5�D��:������Z�K��͘�F�^�÷��9;�x}��N�F3�gW��<��[[]��3H�N�����j�S�qݕg��4V�Rn���0�{��<o�f�S�K{5�1��V=�����~��vx�{���ϧh�=~�O<4r��m�9��3��D�{��ᘏ/��o����=�]�v���pPv�'lFeeYF�1���N�l�bէ
���}A�/�����)#�<:��'��Y|(4��p�g7֒��0�;�R\��>,��o��+���{�W�L#��}�����~~#�ݠu�h�N�=!���o9�o웃�//����OvN�;���T���ٹ_nF�|6N�c܂�KHc�p�6\
h�<2��w�=����Q`�aA��n��2��r�����u`����iDx>:�"��u����ػ�_������0x`��0`�����$H�# ��0`��0`����08�� �]��O1�w�����Y��<(��9�]�M�k�}������L�o!��d�E3��7�s��t�)���M���?f�;7���^Xe}���{\�/E��L���^�Q�r�]�����<��ޜ獻׷l���N�u�c�������&|e�N����ُ4h�a��3�OI��w����+�gf��lX/QC~��ن�����G��Π)�G݋{3�I9�gw\>�a(�,ݞ�7�n?Q��.=����><�e��}���ޡ�)ݤ�6Ӭ��xl����K*��A��Vu;�c9unc�W���w�7�3'�^�n-~����^�w�,�x�۳��r5��=���랣���H7�1OU�ݷ�{�	s~�k7^T}{�U#`���;��g/����O�� ^0[�U{A��?k��N��s<����>67�#�&4�]K�Z;�{�o���'�i��_x�
ɩzOa��'7=M�tvEG��dzaܧ�qQ��C�@�Y�X�"[�v�b��|xc��{��S�y�����s<��5�.%>��U�C��P�R�����wӶ�P'l=�1���+�����dq�����6G�Nn�÷����z8��}��qA� �뽞��}^���N��=����i�ǃ7�t"G�X�w�V\!�Ӊ罼a!��y�~WP�ǲ��<�6\�[�ל�7�}�v3O������5�y�!�s�y�v׆��|3v�vEx�j�{0�㩳��"0k�34�ըi磷/�y�,C��=��W��B�V����xs[5���c��^<:޸��Ǵ�{�yޣ/m�
	�C]%����ז�E˗���4�Z§)�~Ι+�ƶ)�Z&M��^�VE<���򫮥�}3�O��Q�8�V��'N���k���I�D�{p��]I{8����wٹ����*(��z� ݧaK�^l������SWI�����ůL�r2�ҎY��ޙ<�Ƨ�n�Z����}��	fq��xg��f�\~>�y�>���8X���Ń�Q���'I�]F�곥;�A�.�h�(�<n�%��7=)(ר�v�����s�(�٭F_L�VP3�=	|�ҽ��t=�`vY�.L䏽�.����[�wu�LW<7��l�GOQc�k9¶{� `���a���)�D����ξW۲}uW7���Rr侙�k1vG�O���.���鐬Lq���j�^�ԫ���}�;��Ŏ��βo��tD�����������M?VJ�=���Rs9��G���Ƞ/i�;�Vc�rX�^,{��L^�����Q^�
�� �>3�JG)�g:ے_D�N���;"[�}J�ۊ��A6��F�t�Ẽ�� �,�w��G̯���O�f����`�����X�Y���X����{|��x�������{w)��O2/��
�<�pI&��(h��Ua<��jo��Δwfs�t��l��~s���eN{�g�|c�.ͷ�>��U$�fx~9F3cCw�ʽo��u)�s��Yw��peq�
��q����W���u��ݛW�X��ό��u�m�L�z��6�C���Y���%�>>�#�x���ò%�n�5^뾋}.�cx����=��L�C���%g�^����f?�{*桑�;Љ�%�����Y��~���;(�c�4�6�[�fh�N���.!��$7��7�����]�]�b[�����v��+f=�{ �x!a��㜴&OM��ˍv=�Oj��Ӝ4�	��js}��Kk��N5_?U���o��+۳=ă��˞�����vFsr���4)��t�/=�Y�����x�՗�����:4����n,�=`=!�R�����t�gK.�5�J�p&�r��I�����ۀ�N�d��e�6��l5��Q�;���{��s�<O����W��
��)�"���Vn�#�o�h觧��j^|��2)"�R߼&o ^�i+��7�T
�Nm�o4<��e�J|��I����^�dɐf�����pv�_z�T��.�ݻv�{��z���;V\�(����'����������P�����CS]�mx�sS�@vu���g�[��nw���zՑ��8�~绞9�8j��o�^!�vc����w�g4�o{;X�*^����re�K�{��%84-��9uu�7��y�Fw�ǾS=�N�2�#q�36����/.�Q\ǧ��E����{)��3�����d��L�v?jYd�&w�>tOJe3��.���s�P<��}����z�z�����5)�v������uBd>�_o)��8�����XQ����r�������:R�z����6�x���zf�O���B��זq6oL������4��M��z�t���:���{41�;4]�fypp�X�(��͎�����YB~��{͙�gz��E4��X�>ي��%o�����6�1�]~p/)�༂��}�i���/|�!g%,�A�o�w�&y�v��}�Kמ{�~7���X����LFnLJ^���[<}}�E�y�xe���z�d��hђ���O.L��Bgݓ�#⧛g;�2}1�f�����F�q��tb7W�yC��K�f���B^8���*u��=�3�H������Vsͅ�M�;}K�i��j3����7)~�9 2O<����Wb';�2+��ڽ&��/E��9�Cτ9���;��2��P�%���\3޾뜡����W���ew�:���d<�r��3�؅Y˖��a�&s�����cոE;��x�(��r�p�>;1`o;������m4+�;]���fA�mg~��;�*�G{��:G�-��Iz��wڼ`���5�/�[l5Nկ��\�caC���b9��6}��8����L^�}�6��z�fn氧r�r��b[9��e����T�ί9�w�,�uP�(n~G�e
�q�^#T��nm̝�:�ѭ��]!�ݡ&�����W��(��j�Sم��;����_NH�����{77ە|���tm��A��%�z�'���.�2��f�t8�g.sq��Ni&��H@�٤�:���v���.z��.3z-������k"�̳�X�j��w�B/�J�Gx�U8��or��swۄ?T�����g�)��CV��}<)��no���s8˸K�vv��?yk|i�֝Ou/c6�d�z��G��i�m�/"��"t�}�W���������f�0�Uf=��d��j�c�}�<�?f���yE=gb}��%Om�n{�ʇsv�w�ؼ�i��ٮ�
��u�ɸ\]��h��J�V�Lç��<J�t}��_&q���;���=٬)���}
>����x�t�mV���������p��]�{���'/�޶�׎91��0S4��Lc���g)A�����u�p�0����{��o��~�Xt�p\��{:�Ֆ/ޜ�&��0y��:�Q,}16�8����T-ӵ�t�N��!�G�~�'{��0�^]����c��|>$<v{���#��=���R���c50sy�m�wH��L9�K��(m-�0i�z�i�L�;��b�x��a�Ǥx�D�����4t���j�tu𾕯bI�8��n��=�7<v�|�<U��z3fJ�z��;�%�_w�#Z��<��3;�i� ���ݷ_�I5=�1W/�}��.��A�p�"m�����~�X��:�7ݝ�r��ǭxc�����v�V������w�����4����i�/|7�e�v��;&w���c��l�'UEf�gn�}�Ei/f�2m:<̩��@;�x������C��kd,�w<x��X=��ٝ�D|ߌ������v.{��Z�7���5x�Ly�|�ļ@qG��y_�gM�S0�C����d��|4�����4k��/�i��n�!s'/��qs���}M#.�&�7�����d���7�3����J������ޣ̉�{4�S��=�Q��tLs�[/�4�/�#��q��Fۀ>��[���&��yw.]�h�G���5���7�9�クe�D�4��dA���_oa`o��`S�O5����'�������=��@��s�Fs���sLn�������}�mU�b+��.��Wu��՞��W=ji�o������mi�����{��wzy�D=E}=���
�В���S};�cB��+^��Jg���f��1/k=�����w=Ox,\x��8]��-�Ǟ/?X������M�ğyS�7=L4dY�>�،�
&��C`�=�"�������e^^�x�ܙ�;���e�f&��DΗ��e��yp�mR��������uu=az����uvlP�y���"��=�+��:/���}=>���h���w~P_N���r��ێ=�<��B�t���.�m���ݚ��� Bnܩ��]��tE:�\ ��3��. q�wg���S�?R�=��<Fr���yv����9�?7�{a�$W��k�׸v�8����vףޘ}r���������*L�8|Sv 3��{�����2Cs��I^�9w� ����۶{_\���o\��{Y_�b�c��h�|��8l��:X��De�Ў���\ˋ����ܟ�_|��x����D�h�SF��)1�	�J1e�b����l�I��28�u>�;��5,a`o8,b#*ٽeBML�5i��^�>4q���<�b��f�q���x��ۉ��I.{ZFs��9�����;|� �g���J����|�s����Ox}ǧ��	����j�fwv>�����F�&)�]�<�-�l��ƺ (�8G�L�k�x�	�Zs��p22�}��F�/�C�  ��c�o�΋|x�P�hk��|��s�Ϋ��u3�[ƀJWF��j�;��]7Z�fR����yg�=�2籬��y�Ӿ���,T��9q�eԩx�z.���]�-����;�mXo�=��R��@b����o����/#뿙7��L�nPÇ-�t\?l٥���|еܾ�c6<�x�/=Q:7T��F����0ݹmS�n���v��GK�͏囖���k��FB�a�^��ln��)k��k��k�6�ﷶ'�^.�;�qi�Ζ�������i>1�/u��O0�1l�����#�V�'��ˇٮ5/��y��W����o	J9���;�������c���%�ȗm��(�rx�c�4	0�+�8_U��`�_�Ty{��r��x��(7y����8��7yg3���k��E=�NU��;����9N���qg��UK�H��B<O"�p&��x��9����P��!�E��'d��<�}��z"�=���"�rnX��7&P���3s��rM{�p���*��� �J\��V���+<8>�{��b���b��q�<:��{��Uj�<>��LY��'�jp�&,�N;�l�����"��ӎ�~��)�&��ݨ�e��7��IKs#���Oz��l�o��rW��mu�˼�W�Wō�7}�gY���m�\�#"��K���,�g���ɶ$��S��8��]j��gS����AQ_�??���_���W�O������]���(��ޯE�u�R���<.��9�.��/��[Bf���	�����\��iude&�UհfrY]V`L��u��n��=z�X���S���η��7�q���.����GH�n��v7�g[Kt�a���1l�\Ą���\`{N�i�Bn��u*�� iSM�^k��RX�HK1D���-tle��h���/�-���_�s�v������mjE�гR��\���/Qb�PX�s�8�J�.%��(�i��P6�,#&tnl�gRVm�.�6VRXF���3\��������K!.u��+W"�Ql˭e�؄�Pf�i���V;-l[���-�tH����pbh��l"���ؙ�����`0{kG�����`*�.�׍6)��laVFm�œ�� ��� <gC�L褌�&d��%�h-�2�ͫ��5�QҀJJ�*�d��Ј�Я5�S��ۣ���Wfs�l6��A����%ۚ�uC�i|'8Qb-p�غ���j�6�h�.F�w(����=jK���ۧr:\��Wjzè����9x#��k�3&ÚU��WX�).�Rg��	��٨B���[�YpubJ�W���|Ov�ںtq�Q.��h���\ñ�`��f�ۃF邭f�Vv�!�ͫ���s.s/\!lq�\Un�f2�]AR	[��9���{Xk��[<-�]۠���P	����a���AK��;,�u��&�,��e\�s4Ԫ�Fn�A��c��m*l�fʶ��D�WW@5ل������KVLu�D����X�J��q��;��zq�+�Vu{oG:��Iv�U�|u�HvE�g]U�[fuU�e�e�˝Y`WA�2J���mv|�ɫkƲvi�S��m ��p�
����o���i��T��n{�Ss��\�4���HYtk���ba)z�����d;t��3XǬ����u�V��4H�[����p׳�2�mf.]8�Χ�:���\�4'N���9b']�&�5�米�J�[n�7^WB�^��j�f3EV���55�u6�S9����o=���n��.�Y�`
I�'�q�b��X�h�\b�$��x��k�v3b֞��!̷Fq�"n;A��l��%����۳��6s������YU��ør�W0-���MEL�)�s�W[nͺnΧ�>�9�{�q���t�R�U�oG�h���xWl�� \��.x��6{;1�ż��h2�ڦ�k�sAQ��1�\��M�ۉh� ��뙣��`���ܬ�:5d���h�gÎ1&*�%�6���j0�k׬+F�%�^��U|�ݍ���Z�fiq����n��t��fʼA�h�K���H���մ����(]ͳ��\<�]�C�׉�I��Xk���Wh���]���ʏ�<���k�.юR�ظ_W����VyL�JԛA�V�+r�k���%��Gl�O����f�bL�%��f6�Q��\����v[��q9������by�ܙ�^n��j&֢K1���[��p�����y�����[�̞L�v*��t��%f,W=��3,�b.)p7,Kf��}�t+���\�m�HD^��\/����P�{[�ݐ����Q����n�y)|��S���9��G��s/v�Q��=Uv�\%v�j��!9��]��6tL˥!�5\k, ����p���p�=]�'���|{��~sm��Aq2�v�M� -ؐ�2��q�+��n������m)�n�H�9���R��ty�g�m��iI�Y�:�G<�Mv��qv�k�.b��u�8z�Jz����[�v�2�#<xREm��X;�+��Y�����D�;b-H�wd�r �k4i���m�,��q����r����粌��#rn�p�-�g��ʇmmpЁ�l�cv���6�`y���7��ֺ���<����Ǝ��˝��QëQ�����㫩�u����G��N�.�1���)�T�YZ�j��װ7\�YCX�&�.�ؒ�����By��r��3Շa���ݓ��lt��B���_<t+�f%�CL"%�� �kt����O�v�K���[4mKYb������$ڲ��m"f\���B�.�I��m���"@4�ƃ����tX�(�:������+͏9`;4�cy�l�Wi��e��"���.���d����hA��#�!X@���,2OS�v�h�;�e��Uۅ-vj2�l���1�M
D�
�)��v�(��A���z՝ᙜ��v�r-ڴ�ovtC���P�ݲ�����S7f����=�	��>��2��Fd*w6ζ��Sn�MVb��l��u�#y]� Q׭�k�^����+6���:��%Z��n��S.:e���5�J��ѧ'���L��;m���y�O�s8�]<�iXԖ�pX��ꂰn5Xm(��tN5�n��6R<����Qm�n#���$�鵌��ݮ�!��Q܎�c�n^�^,l16	��v�[�eUJ�rU)�C���� M��N�;Wnr��oV[ٞ&���<J��+�v�I�|{|�Eۊ��#��
���g��ʯk��Rb:0P�mՆ�n�8ܰ1p��uPW���sۧ�۵�r���'vn@C=�^L�%�y(��c,��5*��c(�*6_Zv�^&=	��7F���v�ϐ�	):Gs�+��ؕ��Y������i+���Ky,s�#nj<���M3)��gu�q�����-���ە�m��ƸxX��3$܏!Ҷ�����;3J��[��c�j�Hs�l�Z��nϻ%��_h�\θ�Xn���ZR�������2<��g���%�v�6��8�BMz����&�Hۧ���3k�n��e���1ܖZ�[e�n+����UfnFj�f�c.�nN�A8l۸۪����+�`2�6Zpr��M4�+�r-P��nf�L�:&c
��X�/�^q2PSŏ)�e�%1�B;��np'J��4	��Mf��`�uz�8!��+�;K��+-�1�Z�I���>�wsb�#o3�]a�CqDn̫R;S5t73M�0� 9���̜��^�ֻqgmzĚee%y�
�5K���ի,���'�Y�X��6�{d���;E=��lG/FW�))�k��=�V�,s�m��3��@Z3z�4�3�+��/kŜc��r<V�7#�
-f��V]���r��Gn��s�Z�^�[�⇝�ܢ\�
k�]�p�m
�ۭ{���!�N��oluL�s�{u�lv��U+�����L��
=�[�<�*�n5���-�l�{t�]��E:2����a��+��6ݰ�xhr�s۱���F'��Z�;,�B�Z����j(�GD�,�ml뀙�:�cuզ ��<�Š�L���L����"��Qf	�aXh�ݴ� #�Ҫ��ib�ێ!GV|[�2;��R�KH��zv�5�ݸ٪hy�7cK�v�u�.X�r�9�0�seh�����ͮ��kC붴���v!��`Ξ�^�R�[�i1�g�`Fj�����)�<]��Mð��W]ð�����m[��R�s�FS&����,@:;Y�o7�UBۮ�͵��tڔ�W/iJ��)yZ٠4��YZ�é���-���)�])�k-2�un�,�dB��T�H1�q]�R�<�:��7]B{�$6����v�]qP>2���6�1��>�+\r��0�a�x�yl-eV�˗[+���$ֵW[��ūv1�"B��qO����"�m4ۣU��H�R�;q�Ü�^�n���>w:3م1�xЦ��萉�b۳yTD#en�1)��0 �N�a�i�g]�tl4F�F�'�h�_&m�%��f2Ё>l��b�m!�F�md�(�-���lnE�����pp���ԫ����W#�gcVP�b�5��u�R\�������\���O��k������AK�2Ϙ�e^c�g�v�q�!h',�;Wu�]�)�3L%��ٳYe��ڧG!s=���t��,d�uz�8�ĝ��JXx�(��o s�s�&yz�Sv�"����!˞B�yۊ�v�;W=���<���yKn{\���6�B��:�g6�璻7OW6]c9���by7��Փ�y6�!�I�'fM�hv�m�>O<,<ZF��\����6���7Hu�G�7j�d�s�v�we�Z9��2m�u͉3���e��k�ru���m�z�]g���+�< b(�O
�t�S
D��6�df�Ґ�[�� �y������\mI��\  ���$B]�J��곹������/=97��\@�%�32`l&��-	T�E!a,@͢j�ͪ��2x�4/b7Wi,�4,�R�mǓ��t�O&O]��Eg�s�(����"�{Z�n�h�c-�w*��895�u��7kg�݋�B&��Ǘ=�����GWs�y�/<ܝZzS�^��jc�����ml�b��%-�ѵ]�]�m'��d�杸c;��P(�c1]6M-�z�XCWXEKGY�3u�a*a�������9Z��ٷGB	lurU�*�J�]�L2�62�]�3)�����9::��;���Q��.4�&0���_>|��"[����wa��,�%���q ������XM^wH�`7[T��:�'Uu�5�G@X�s��܃K�#�TM�Uu���B�����xܖQ�3;\󎐪��S7%�^�8].!U�������v��\��7M�n�tI�E�u¡�E�q���Q-g9�/`ۓq)	h��q�ٺ���=��"i�sSC�k���Z���m]<�ɉtnmU�B-t�:����fX�7VuEY�EMs�UAj���e��e�����n�gT�\f훍V���V{a�l�ˀr똩M���ͽ[.�Y�\gv�cL���^9+(p)n�����=Ͽ�����rw�t�e{J.�n���A�>���C�r��;���[�_!ġ鄏Ӟ��'���<c
s�h�Ҟ���jc6�@&)Huy1؀�B��)�]�'�ru(�8����~7���7?�3�-2�=����.UP�0��AN'����"�q�X�F#*�y�eħx���V���p��L�,���H�e���W����g�AG"��'"�B�YQ�ǽz�;���D���^��%Q7�z��&: Q�ɊJ�p�N���&<x$F-9�ؼ�����]͖y�� ��?x�9�N\��G����z���.(�;kҝyC��JX���򲸦�dO]҈7�EZ+���:����@,H"ddF�๤hjot=|�:�Dw�t�u�P搄E�'bF{���p����R7V^z*�r=��d{�G�����5V�"4�9�uU���y��:K+$�H�#�����LuQh�F���-iZL��9��b�_+��/�'I'��Eعn��ix�j�%0�C0�MX�=�fg���N��SE�p���Y�O/^��vvE0�;C��n�4��Sv�=��ۄ��dzj��$�Qcq�:��[,��t�cai��bVgkI�h�"��Ѥ��i�<��:�l�Wj�1]s�q̌������Շ���m�z���P彈�T1I���ʺ�XKA��ӯ[���U���ݷ\���&�X6�ر�IL�tƩj����fv��b1��)Kj;[wnm���C��]g9FĂdv,�k4��[��� �U�����64��tW<rwg�y���Ys�F BXS��5��2�a�#��n�����&��%��!��K�g��n��X��-�F��v�U�JjG��Ҷ)�����l�6b�vN��`J����9A��jz뎼M�9�&��8��δ|�]4r� 6m�[�<;�V�3��q�p��.P#*��m�M\-%�G�u��D����]M��4+�"��NM�2ᵁ*HX����3d�홳tsaQY��c�=�Ǎ�2��n�q���:$���Kȉ�z���0�ݴ�VR��Li[C��c/V�h\M�6y`�c�!��rus2��FU��͛f33�Ж�)��K�e%0�Z��3s��D-:�"�Na1�wB�XV����t5�ƶ�0*�pڝ].��1)J��+E�T�b6�c<��a]3Ԇ��^��t9�8s����ro[TV�;��鍑��h}���>�+�0m�[��ڸgs>7>����=���R���uVǬ���$��z�Ι,L��Q˫�s���ͺ.��k��w`腼�����������v{Z�4��Ҡ���W
.x�*���i�m�4J�JK�ꋠ�밭��e�7/O7V�!�i5vײ�q�!�ڮ9xg��(��1���f��ɳ�Y��'���Z#��g�y�I�3�U=�{�;��gm��R��VQ��k"�����!BV� ���(�/�*4��<��	mbJ�l)ZJJ�H0
�*҂��͑l�[A�&�/q�r�Y���)
�Yz�m��0���6��b)Eba-Z�����B�E�˘�{�R8�W/FЯ<�*K-�V�Jش� ���|�_���S�n�+l{qZ\���<tsg�p{��벁�In���H�Kp����u6Ֆ�d�w��Ohw*��d���7��gC<~�j��u;:���(3;�\x�g/cfk.�B�|�Άz�	�����|u͹��9߹Z~����7%�����3D�?��cSA˥�����+��]���/n1����ɼt.��������h}��KVSo�Y_ T�~Ζחp,��.�Α�B��q�5�{��>b��٬�i�ڳ�w�?3;����q����m�2�2�vcub�5�ce��4lұ.��6bdʘ�F�Ȼ�.� �O�se��4�F)m-��P�!J�/��`�)��n�93n����.$?n�r[yC����&��9ô9�$v�Y����4=吶���F{��ԥK�{���:b��|�F٘�����_���_����D쿳%��M���ֈ���wfwj�Ne�����a�����5k����B�.���r�mV۸��DW�H�@�.�do�n`��юf��1�)��m�%�	��ͨ]�p.�]ߑ�1�)j��p\��༿o[-��v_���[n���j�?�8_��CpnGCH�[��]XUאf�Gi3taI��1k)��J�����z���л�.˳�êk�[�e�s�I���r�nL����9��i̴�b\�b�e{�lg�Y
W�������F9�	nc~S Sh]�z��a�/ȍ��_]�������p��${L���p�סa��\�6�D��5o��Ӟ�؎���>�]{�V�a�7�}�=��V�r��u���}�j�ș���묇i��el+u.���;/�j̴�rڲ��?�}}�nG�8�� WhF]�[5�٘Ql\�Q����wz=�ؓ�^�d`m �M��@r�1�ZY]4&7Lk�79�%͉����OϪ��[W��{�����g60�O��8�b� �����n^�88cNB�R�#e��`�2�Q1���ػ���������h��E�s��{�W2���[Wh-�5dVz���l���F-��N��F�]���m�L:�~��� >�?]9�r̶��ic���K��2�د�{���±�
ܝL|)���>���C���d��\�s�~��w��ꝇww�D쿲ڹn��;� O����G�L탺=��\(�j�ҩ�S�T�9wY^y1�Y��!�,t��Q�g�z w��T�{�h�u�,ٹ�OR18a7=fujӖ�j�q���ٶ��f�6/�b���ɘQ�\�j�@��.ƽ�9e�7��y)
�ˑ�5�ah���,�]u�][�u�iz]�ӺC@G7�(��������Ne����o����nN�7g� �T�^z�T}w���`���@��f~Ǹ������O�=���wn���ChSה�Y���m�ۣ�'�/�~#��[��Y��˿���9mYi����ܟ�W�^��'��q�63�6��jX�1n���y.�a���v��"� ۋ�_\]����Pԉ����ֹ��h�;��mY)���[i���� �Ҹ���FK��Ռ�I�v�,H/-�����{sTXu��L�L+�~�e  ?!v+����n�|~����׾z������ptaZ�j�N��	'�1��y,Lr؝zx��Siu��,��a��]1��j��hMf+=1�qGN�N4g�8��<n|Y��u�n���J�6V�v��qE�::ˉ�m)��m3�m�{6R�����9�k�8-��q��I��vƈgk���,4]f��c��Z\m�m*zāy:r�r�Ɇ�NY6B{uN���K�@гQ�-Ň�����>Kn:K&��]��c#�luӷ;-�bYt[qj�q6�<�%%*�-f(�A��7������ճq1�\����엉9��_�Ch|�Z-D��ɲ'}�6�z�����y:�K�0Ǵ}5U�	��R�DP�/� L��8�]�ݠ.�d8��/ד�d��}�5��Ǳ��C~@z�!w�է�Mc�;�o5�㖟*׍+߭��\Le�����x����W:pt���>���w��J�pӏ����#�p^m(�/�?���]�w]�un�2�����w/�Ľd컟^��Ų�4	�l՞=�Yz�!�5���)-t�}�����Ve�<Y���Mb��?^;&t���������n[U�Ӈ�����=m8d҅����/=c��+�u�ћ������;<]�M��������~it:����i�
n����I�ܯ�P�Wݑ�dW��p�:�6�Le��P��쬑[w�ӻ�4�C�@]������*}q������e��(����~�`t���i�Ӗ�,~ů���������k���ɝ�;���:9��9o,��Zs-�-�^8L�f8�����j*���D�x9߄�wv����L�����=��ŸF:�R`�azq���{M�ݥ��Z�.ƹ���,k��qwh8�з0U��^��Ɔ̶�<���}__�����2��̧2��y��{�{w�ڟx=��.��T~�{���f,|~�9��Zr޿��{�����eo!8J���K�~Wo}�]��W�:-C�k�r���d>r�zTa��rJ���5ۏ�琈Ҋ��3�5W,���䵿^~#}8*[������>���5��(-1 n��ݧ<V�}W����w�럠M�y?K�{��ne��'�g��3ߞ`e�P��.���鶧�w2�n>w�#�e�>�z�2���f�ki�]�]���.�G!vb6���f� �()(D"LĹσ���@]��p��n��Nn��A��ū��;�s{��.�����whg�R��١�*�hVo���+s*�1+ׁ����N��u�o�῟n{#��9����~��{~���&W>������?6/�s��d����әmXE�L��D����/j�\wj�eҚU��}�g<1o�j>�j�&2=:T��)ӻ������x<�|�l\��W��mx�T��ў�qξ׺ow�e�iJ���W@��Vr������_d��O�՟Zr�{�~}���AY��|}5�[ʁ�L���rtc��ڻ��q���g����H�߲�h�)����o)I�%��=��q]�!<�"�I		�&aDJ��ܱ��u�������F��kq>�ks׳u�(���7��[w-?Zr���|��Q�g���.���>����o�������6ݙlܝ�ʁ��T|����]�v���;1�0����i�9����O���c���t�[m�A�D�R	���֜�@�׽�G�v5��x=�	�㻻�����J8��~�}i�Ӄ-��~&���Y6�77�-V�55��� �/
�5���볏J#*�mz��B������6�Mm�B�ǳ^;8��}�u�z�g�� ��;s��y�^s��$6�36zK(1(�K�X�"VM p�퇠xڮ�u����Q�r����;��Y���ս.�8��v7k^��CXnk�&��.8��Ջ��*:�m�+l�h�]�����Z4!�f�*��v��\�9#�\�(<�7<�:�h��d��sn�V�7�E1dc�.�nN7�1vm,��3�G7i��������;���:d�ѐ�i�%�k.�Q�˒�ѳJ�V��;�8���A7[��/W��ف;K��C�!'k�&,[j������ߑ.������lg���l��b}x�y�j!G�}��JrӖ�i���;���y|��Z�=�;ucm�W���K���mT����`2����������3��h��w�;�?�oqw�zx�=�}��֜�m�`���=Z翶���|r��ݣ�<f�kd=��e�����2��VF!N�_^�ܻ����ݽZ��뺹�ʿ3�Nv�n�e���{���}w��^,�������h����5|���E�nn�t��:ٮ�IṸ�!�nn̴}}�d|ޫ������O�u�VA�fB��������f�
m}w]��v�Xu��+ua�w;{���!ꮞ�0p��];{5iO$����o�S���h�ߴ��qɶ˩�0b캍d�Y��w�ɔ|"�^~�5�1`��GVٖ�}!�T���:1��s�3yYQ�+�<d���� �����^���Ơ���Ws�ss;�>k�6���疯h����g�{�?;�&��!���X���\md�d$4�hO�w���G�6�}wv�����[f�o��زW�P1�L���u���:8�Zp.���S���L���!i�����^.�mt��Sۤ����Ϛ��>q�)�"��g�@z���p��n��F�X����߳j�&�.�A�n�~�s-�����F`��Oi��y���}�q�ź�+ ��K~����]��s6��1�wF�A���ÙNf	b�|^�����{���_�����/�mr�~�[���(��Gۦ�<b��~5l�����i ��:���\F듔���f��/j�9�O�zk�����>��Ք�C�o���l�7;���s�~�u�x^��zڒ�xm��r��0s�c\]��kJC�t_bu�t�9FG"0F��Y�|{���=om�}��R5������V}�Ii��n����Oǐ�\��7�r�0w���_-���}��n����y�ĳ��K���+޾�����T��u	����������g���y�{bA�^OX*�l���;f\�\`/{����Ҝ��0H)&R�=�p��F_S�w�gw���x�{��7R�p�g���C��h<s�皏����y�n�ob{�r[�	md�5'�²�|V�K�(į?4����>Y��#*v��=t�<}�u���Ċ=ՙKn�D��?3�l�]fr����W�;��ˮF�tC�^^۹�c7I�Ù�/C��Ο%�4-���	[�Bb�s���Z�Y���S����|��lȫ��sԏ?+�g>���h>X�x�t3�����.�v{ �t��ʏ,]���hC#^
��ou������sϻۛ=��(XӾ�g3�"�N����Oi�A�q?�9-���ڻsޏ=/37z(����o������G<����{�uomջ�(0z4�./o���o�9nA����ܚ̪4&Â�ʩ��S"e�R�_��os;�͝�ץ��KO`���I"Lġ儙���#%ĸ��n�
�[.�G�*=�w�Bc���.���8<<<��|����g��0��)�|+����w��ϞP|$g�l�	J$��f�W]�Y�*YI��'���b� HS�ʜJ��[.��,�ن͘Ueh�jP�i�K�IS��hV�F���C�AN��I1ţ��g��{������� 4cȂ��� �����.��.�+���:��py��E��Jz�<UH����!Ⱦa����ۺ$���Ϙ:n�"�.I}_Z�>\�s+�
���Fz�Zp�((�9>�z�SY�P��-�J�B�.a9�{����jcK2�̚BI�2-���9�%E��*=�8I�@�����	"*(C8�j9���uqۡ,����Yz$�EIa�N����.$$��N�%R��rY=^Ey�UD� G,�,�t���V\*��ݸC������n+B#�TEeQk-�V��pqwr�&�d�$G%���zY&�U���;
"�$�����u�r�?';��;���)K(�K)P�)&�Y�7tU�XYU���YH @Y���g�-fc����8��܀� ���	�� Cp!���'�ϲ~�����@�AP_������s�''�:���^���?) �	�"��<p�g��7IA�� �����[���s|����5�p��Y�z'W�󎬊���ԯ��m ���[_]Ӵԛ+����4ҬM����˔v��>x�:5���O8��� (��6]�s����|�zo�׬?�/��ь�{�铬�e�=�Ws��9�k �{�@�A�g�� ��_ۑ ��"2
��"7w�V���H��h�����u|˯q�n�
08cC�q�SQ�Q؁�p z���Ol �m����Ќ����a{�]/E󍬊������^��6��?���!��r3`rfT�ĳ�5�=Џ͵?FN����S���O�Ȏw`����;�סK�1M�z�����!eʻ�� χ�؞p�ׄ�����zaR��Vu8G��o>�#o�wL�_��������c��{��ّ��|s`"�A۟����_c�C޺�2�DK~����Ջgb7�gЮ��߈&}���w��l�q`����&��F� H&(3�^��k%�ݺ�m��O�����i�u�PS�f���?a�z�$ܑ%�������^��Y;���(��Y�^����Q�y���g���[������>��ʔw�|��>D�Qժ���U��b�^��9�� ���$�\s��S�Ə�Vy���A�|Am�k�6��w�N-Q"������w����׼��_"� ~m����TFx��I���ܹ^�D�K7�7&=�:��<���A5��vNm{<�Z<C�/��|�p������k�q�S̩�G�p#�ԁZ���+��2g��8������p<A�x};�(W���r$H�^�P�?��|p?'�9s����������^q��`�=�������=I>�}�$��iyf��`AbD/��bz�A3��v�N�0����'e��s�hM/��g��5��AL��v��դ�x6�e��ú��i��aL�øN�e�>�2���s�Yw$^���,!�b�"qo=����Iۢ���:⺱�E#�%��Ssz���O)ф]�5���l1De�,!+3ڊ5M��{u"k���@-���M,���ۘ˜���j�0����f��[�=�~ϥ�tmR��I��颕M���]�n�OL��F4q(�Q1�3�q� ΁@����6�Z/i���:�ħ�t8�:���&�o��*D�U祭 ���7����Hn���J)]*��� �@d�����>��YJ3;������ ���6�yͣ�gN��σ�E/�݉ �~_Kk�q�-��9^!�Z��*����113�ǣ"8�`:܉��Ch�R-�,����"`"���'���Cq��{Qo+�u�ݩO��q��{��9@�o`Mov-�|q�?[�?�|�n D��n=f_j�g�j�Au�j�[ϕNI����L+�$@mCn@��q�Ǔ����зH�C���85"@sN.^`w8귲��d�m�v�Kvlr�&���������Ӹ�E�@��6�ժ�3�F�s0�X�dG7d_Y�;ք��� ��An#�輍�dyc�#i��UD��H1B�Y/�7jBLc�v@���)��yN��Lfc=��?0z�j��f�g���l��it�C3�'�g�e�����}Qo+�u������p?W���Am|�-�P�;�'7Q���Ed��Dr$�m�'NF�����MF���NI���k��������7�qf%o_�v�j�A��Cԁ�������#�50�X�dG|A2 @�s����"�D}5�O\ � �m���p�6�����9�ޛ��������}~�0��q�yH��� A���c���{�l7���J��k�4vi���Mu�r��q��]s\z�qP��tK������8�Y/|����p ��ozڍ���s7��!�"<caO������o�'�_ [��m���ͤ�ts����	���|�_)��������Q���"8� /�:�����ع����: �����}A��?O���սmq*)Yr��^st�*��z�����0���;jRi�P����Qw�Þ3�u������zMҋ��`�Y��ϋ����,737L߇�0c�wձ����˿td}��O��-���@��m�7'�;o����7&�A�܉:�h ��mj1���s;�=��z��ّ����8@�����p�ؐA9�����E��Pt��-c�<�o��k��&����J�V>��~��H-�J6��s��J�ɻ����AVx����٢�.ՙ�ƣ{�[�N�9���a{[9IS&4E���"ր@���?�ˬ�+y����&[�FG�8�z�]�[꥿b�{�mI�D�Aν��mqZ�X̅��s���[����_r��9����zh��s-�$�Sg�|��n �s�A��n?6ѱǪ������>���;��}X�dG|@ �@D��[����6������z���@��#�Г��ˬ�+y����&[�FG�����.����?�y�d]On���#dq�->���_/&��g�����{�v,]���/'�}�I/��|h��V}��eG�Dp ���8,!��@_��O��iw�ϭ"��xr	z���Q���s;�d�Mz n m�?_U탻�:
�^3AF�u�2��K�[3�E5+���*�A�=A����[Q41��� �� C��-��mH�]�ܔy�/D���/T���P/� � ��"A܀�n!�2	n"4H��T'._w
���H��d|��;J�w�G;����ё��~������}�L�d��k���{�� �r$� A��%��N��"��{�x)�9��9���D�@"<���m|�-� �`�D���0A�=@=��ڑ�v/orQ�9镙�"� �a�@�Ïڕ�Uf�9�4��"mCn~�~-��� �_iXki��k��9I��r��;�}A4��Ck��n��]h�G\#���ײ*��z�{�2y��P� ��3��U�7���=�gx��v�=�=n���6�?xvkWT�^���	~���f{�/����g�c�I�z����aV���l��~��v,��Ŏ��N�5�ez�7k6���*1i��j��^9.�:�C�9��<�)+�4l�X2�i6�б�Mrm��R�E��R���,���s�^5���7K��U���%�����d�d�Om��R���υ�۷z��v7gu��m�J�H0�ct��Ϟ-k��Ky�g�:l���p���}}o��x�l�����vkz���h44���{kr�x��e_��Gߎz��/2~n�-�g:��J=�������#ӹf$k�<�h G�ȟ�m|�p� �ڒ&Uz��^��9��ԁ�z/�t(��ʜ�q�=��[���������U84E �#��� ��!�3�q��2[Ȕ�|a������;�c#���-��nڟ�n{g��}�m�Z�ހ'3�H?n�6��.�Zx�{�x)�/;���A5pu|�z���{ق~:��	m����m|�-�l�w�dM�c� ��#ʮ7��t(�y�ʜ���� ����� !�eT'u� Q�6p��D㭲N�]��Q���zAw%��@�z����@��I&Q�Q1��ݐ~9�Z�����kbW�;�;>�3��G|F���5��_` �/�;�����ǈ?�
@�uÜ3k������/��
�Z���ys�<2W;��~ѹ9�~�Zrgxl�ٓo��O��<5{���D�ϒ%��y]��<�l������Q��qYFo;�x����C�h11����X��ٚ�ߵj�}b=� �u�I��[� A�_m�􉞁�^��m�Q�xr�^���A�� @#7tP�d����Y^���@_���j~6�C=�J��8<���]��~�q�����݅� �֧��A-�D܉�� �f�������� ���O�G���e�ﱮ��� ���Ck�F=�u���)HQ�c�痛�z��>:׋�s�v�-����mC��<Ƙ�Q`�g��{���p�ڑ�v.3wy%�y�u/�Dp"m���:�f p�� �@_� @mП��
��=MwF��`O�����;I����Ȱ�tdpW�$�ǫ�3L�w��Rо �t!�"Kp������{�Sz�a�7��*�]ga�`���X������n�V����֢?vGDx��{��,�������8�a#�6�~I��ݙ�Sɿ��s���,> �H�
��\�f�FMG�;�k�}p �����Ŵq@�\˻����Ŏ�A������b�]����<Ⱥ��">�s��<��������� ہ���[������
N����w�&��(]9ܭ��(1n�2;�	��Am|�n���	�^��U�`�T$k�Vn6�c��3�4�����6-���������%p� �Y  A�s�H-�_Hm��O`�{�c'������r̡�۹��>A����mH"~-� �����a�W=�O�k�|G���S�q�����G�_���=�����́�Y������� �� /�A|Cn~�I�����7�d�ʚ�s1�1L�~���5~R-�� �[jA���3r]s7�� Q�r$���	um��}=�ѓ��g}�w��� �=?���7���.��nr	�F#<j<��t��<�a��h\Ë޻��̖�[�������	��f0��Kq�TT�G��~#� �l� ()�����.�	Ex�=�;�Zaߖ�9欄��Г���-�g�� e���l�Y
���9�EC̏T��Nz @nl��|A�r���tBC�
�q��;;�;�7Pm�E3=.��[Z[`�{t���j��{[9��+D{�H ��m��6�C�ƶr�x��4���FG��5�E����V���2>_ڐCpp�c���8��/�Amm����q�s���� �\Cp!�$Tǻ3�o��y|�{�	��n>_1�?6�ʫ��"����7��⊇��|2#�㞀� �l�-�_[Aۑ#È[��V�j I�R�n���?�;���L��!�FGMߔ��C��&���� �����?7 &܉ �1^�=UV0_ �
}z�c�w����Nw���<m@@Ch/���~n>��� ��f��;�O���6���P����}�m���9xt�ޛ�Z�rt��7:�н���h���zP̈́z�L���b����=Z�/7�Z�{�h�|ݐ���|
�<��1>���E�_�vn�D`{Җ���:s����}C�留�>ʞ^�q�պl��9cU�_l���~�{��sq{���VkW��q�>�f�G�۵��Z~��넻�W
�=�n�C0�/y�{��j���h�ۍ��a�<�}��z���&�m��V�����lHw;��[�q􂬻��^�𼽝�xI���p��OÝ�p������3�xL[:	rL���d�a�����r��=9�>��▧�������`�27@��{�æ��i���O�ƕ�ş{(u�uz���MxvN�w�]����͑n�u��}�}t����ٽH���+'�K]a��ч��Rz�\�ҵ�>٘��C���Ep����.G����k[K���N���>Ia��>�2f�����<�~,xu�~��{Fw���.�����V]C7L��)��VڦW�3�/��{Ӗ1�^��%��ӲG��K4�9����hs4���	�[�5��:�0pޫ��.~'q�x�h��ɞ&�F>�w����x�|i�7��Dj����U�y\ ��v���;�����'I�5���z156?zo�@1�dw'�����?�>��2;E��s��������&���x��5���\�V3�3|1�z��c��KoOU$}��!O�h=�W�0!م�W$���OZO�_~���3���}=���n_E�����=�����U�11�����8@�>�%$NRMl�iE��ҚT��%�d�����~?oɔ%gT�{�W��{��,I"����K^w*)̩$ܲ��IMc�T�*�I�����l���@�T
��s���Aa^w�����EF}��.�����I�yZdrUIZO���}���/%�\�$J{�}G��K޲�^Q��g�;������%<;����h��e^H�ȗ�ϋ{�s̡�Ԁ�9��շ?0r(C���r��$\�~m�\0�3��)�{�|�?%%z�W<Q	d~O=�H��e&c���& u5x,��a܄̥�1D�R��Ž�\�5��֌�
tH��kn9'�B���IJ�_��y�U|�Е���^�IZl�NS�,���p��UЭ���1l�qJ��ґ����pR��>�q"��1)Nͼr��y|�)�ZB||�m'��@T�!���u�Q�B1�y����r'�)��
�[�=�b���Gn׼ڴw}G��^�.-�(����A���'n��s�u�R(0
�U�;E�YֲV&e��܄��>�}뼕'���ꬊ�&W���Gd����*�mtc�!�)a��\���?�vC&b`۫�ȡN�qͭ�֮���X4��pu�j�u�D��9DV|C�5ۖrV��5��UmٶY��h��ɤ\r�&��9s�B�<f5R\�q��E� Y�\u���n��୴j�s�DQn瓌���m�7b�M�ǵ�,��{Aͮ{7\<��<�'N��0�N�V�<�KSZ�#i�H���7n��;��-���N
-���zbp��=��gq�-���[��eۑ���enF4�����ƅ�\�E�6$�r]`Bz��kl�6\�8��^�X����e+��mw2�,.���?��X��)���	Z��aҷ��x�u��[��L�c)q�7bq����zp���6Qݑ��sSKpvҌȴ��\�� �7R�z���	����亞GV$4���E^$�.Ë�`���f�k4qY��W�g�Iz�eH^7.6-%�ir�h�d�n]��1�Q�g���|v�;��$�4mf4����9k��jj0j˰AL�GX�â͝�����]�=��w<�t7n6��b��j)�hh�&V;V�1]����h�`�W��Ϯ{EÍ��ܘL]��$#���Ef��\��6^�D�V��v �kb�Y�lA���5Ԛ���e��&e������ɴ��5�۱(�=t�v|��e��[�S�,�ت��Ya�+)5�2�Znn�u٬r��nb|��]L��)�4�(�0�Me,դwjh܎���E�4M-�b��R�TF2Zr�]6H蹝(v���t<�[=mr��[�ڻ{{��[��sm馡�.�l����v�4PY�����2��0�m�-�-�Ѩ(]�GJ��-���:6ST�5�)��`S�^K�����uٻV�,x��]wg�/]k9�����M{����r���h�ca�3H��Yl�E��=s	�
ǃ\�F���������#q�m\�U�;�xI;�T���Ƴ�G�Yx8�͝׭k�/K�y����>M�!�����W׮ؙ�u��P4X�	$!	!FE$	R16l��[饉{X��t�%��j���ںxq�'X�e�v0�;��xܧ[;�F�2p��l$��:�\]N��m����&�`�ѭ�����uܽ:ms;��=i�n]�tq�Ed��td	��\���.A�[���kp�tX#��\��ީu���W@s1Q���{Z݌]���t�muз7o\Y�zۃr]Ӗx�u�sYz������J~�8v�\�@�t�AvAfh�F�]5e���¤�`
F�Xl�������0�>��{j���mHɞ&�wc��y���"8��o��d�oV� h ��?n���7r$[���
�=�lΪ؁[w��/�?O�����ؼ���L��#+�#��~R?�p�j,���,P;z��p��6 �ۑ%��
����_N�uFTϏyee��k���k��w|A�k�6�E�@���7�<�%���C����mj\M��G%P�#�/A��A��"6����~y��p=AP�۩�q�m���>OݱQ[���!>̏mN�B��q]&��H?p-���mc�U�C�0��C8��BD� ��� ��8��Kq�y����at^kp��V�3~����aޙ�?^d�#2>Y�b��Ӟ[]i�����k�V\�ú^��^��ψn��i��Kp�q-� �|/e��*ښ}<!O]!{7kp�Vfl���r�����᰻��ػ%�<�^pݫ4J2vW���P�w�F����W�3��ه�Ea��RD0D� �dERE�֨���XB2�~RL�&�t~�j^d]K�8�=�����!�A7���:PA؅|Cp�� 6�'��n����������w�>������?�/�p-� ���|�XXǻ>��e��6���� �A�۝9�֡�Ǔﱮ@��{��r���G|Gv��� p��������]�Bu�>3^R9OA���ԼȺ��dGΠp#sP�Cr�[B{H���SL��R�Ke(_0w�˺�pE��sۙu5mn�\#[�v�i�}}��$�{��As?p���R���*}냕ё�L���!9U��v'��9����o���wO�P��ƊD�{]5��7˽�E������H �\ !�!��n�f���+c�� ��R`-�_�"-��`����ң�R.&CW�CV=��ٙϦ#��k׎����=<קq��M��J@~
g6;Fs#����z���q�U\�\�뺮w诰!�R ��(e62���q"�  �$�2 o|�WY燜K�R���@�s�nl�7����!v���p��8��'���p=�e����*}�ձ������|:{\ǻ�`<c�	�� �6�l� Z��3�g����lhA�z}ٴ:=��"��ﱮ	�e� ���V��lm�A�`JJbQ��'�$Cٸ�(c�ꎶݚW�P���r��<ZW�ӿ?�~<q����A���~-�?r�y�;��x�T��}����b|�����["K8W��\ fbp�Dz�����E3:7�6�}=B�:����0�޸=]~��ha�+�,��8uB��V�( ˨�9 C���Ye[C�~�~���s��ۡ�v}�%�2�����(Ch"m}?2���`��9��*b�����j�� �ڞS�/7Gp��yj��f8G���:E���Vj���u>
)W���f�R��=?Q��߷AX��;��n
/)���{�mv���_����S�2�<�;�.ڨ�7P6����}�=��H�"��*� �����$"H�H�*��;��B��Cn~�Kp�[� ���_Nǩ��4uő�==����N�{:e)�Y9[A7~_N5�����md�_lx>�{������������Mb04M��g �X������Z
��6).HT50�3�G���C2���p�At�^��mϽ�_7�n.��Դz@��ޘ��"2�D�@m|�p�?ڒ`��x%we_z ��R����z"�]�T>c�w��y"Ae�`���Y��B� D���t�D�D6��2'բ�{T{i�#�YO6eL��9=A��H#��~-�$7`��^��{0ڹo "͠��{v�5\׸K�e�ۋ�k��#�F�����4�a�?!?G׋��-��6����(��mgQ+�ȱbmO֧�3�F�ML�.���8���~����Ѝ
��g�X�T���5+����w��f��f��o��)�O��ӱ
NQ��p՟�t���aO��uT'1+`9��_����4�"���
�H�B �
� ��,����`!���>�N��\U�5�5��M�;u��Ύ�x�I��d��;�D�^�|��Qv��=ۖ粧I���6�LHq��n5�L@C�%�cs�vqt�v͢��x_@�nI^�ie��]f��L��=N�Y�ŝ�sٰ��z�હ#j��>e�<6iJZǙ�6�x���vC[�aV&fB�[#nJ�.eFЙ��a�gh_<��ϐ�_����s��8�tmS�`|�������[�Y�52��~C�/� �1��m��Ck���2�k;�%M]��ё�~� �?l��oڜ�=�oa|A ��Ȁ�?7�L`�wHu�p�t��u�^���{�>�}�����~��EުX�?�$�d|���e��-��mg�^V잻�)޼gT���>���@D��$�����h/�m̌Y���(^�a���#ۓ��\2<�Fz���b��9팎 �w������Q�=�g�q� ��$Xq@ �/�m�?Yq��s��%{r9�����u�|>�u!Ə��D6���׷2ߟ����s���M��z��L�cnm����L ��p�q�u%�,v]�u����;矮'����p����0�A���Ʀe��O�1�Ͻ�P�����=��&�,�i�`8hQe��.V�l���V8r-TU��������[�����|}�^�F\VJ��Ԩ�Ӹ��0�������r�i�\sֱ�+}��z�\! �!Qp@2��q�\)�65���߾q�/��~u��ä���s�8�ߔ�B�!�>Y����z�Y���>S04�`�|Ay�Ye͡�1�@Z�U_���\�Y����۩���D�D6�~!�!� A�<�z����In/���L�G�ٞX+f�nn�����)>�~;�꧐�V�[�����9џpn��!�"~n ��!��zOG��V�߷�$~|1�o�t�UvN{��K�/����D�K����������|\��k*iF�L�ݞQ��݊����IEnꎱ�X�)p9�m���'��!���?_d���h,�{r�E-��O��w۫�!U#���w0�3�m �}@ڐC�͟Z���Y��3Z��;w7L�L��)>����H���ׂt� S�,��`�3@�̙�����p��ފf=�
�z�3�<�����L���n�t����[#GQ��2'�o�O�߿A������`��dxx{YQWncزߌL�8}����HEBAP$k7��<y�Y\*j��C���������|%����"���.勇��ï�$�hI�������E-��]�ϻ���A�j�"^P���.g��|�B�n(����m �VW�X��И��T�Jz�f��2���dGN� Cs$In nV��>O�4wx�zg"ǽ��QQ)��0e��k+pK��%@�v�{h����{x^�x�������� _f��!�"~!������g3<*j��C��=�킛O���7��%��� �������WwzǏtA����s}Kj�V�3���H&�d�1����m/��>�߷؀�� �>R-��-����Y�Q�*-oT�a��N@�OE=����j �̑?��6��?H�!���v�Ө C��?�����o�O
��'=�� ��� ���[SQ�ȍ�$��e���yDs릷N��g=����{e�=��u7���Tj���w����N���+,ֹ��Y}o\�^��@ !VDX�d@����5d�ؤ�/� ��BKp5�=ڇ����&�3<$c��{��Q޾�L���] �^��?6�m�O����mWnI���o1���߈��#u�Taub��zm���T�������E�ua���;���~�|��1q �Q��G�h�Ʒ��OE=�{1��q�z���� �O��<A� ������tJ��/d�࿈�j�Kk���v2�ݥ�
Ub�{��|~��Am|�q�]gE�4��{���%�A��"Kp ���=�ݫ�7�μ���o��n>�R�@@�����[_"� Ge;��ba�Z��d/�� %��FLh��[�L��"�1�j	�F\�(Q���\,�g���m!?YD�ۨ9��a��~�޶�o}�\�V,g�}�/����! [�A��\̹�+LϽ���z���eUƑ����/d���f���M0&��H����y�x�(�w�zD�@h�ww�����Y������F�l��:���:�s��F�P< ,�!� ���\�S�r\��ѭ\���ʗ[N����zܶ�5�']a�	i?��7����lۃٽ��2r���4Rݴ�����`D�2�6;��R��iu�m�-�W��06�Ŷ�R2����:E�FP���n�v�k��C{ ���ur\�j�a�8r�\�6� �����(��,�F��Tu�a\f��#�\>�	�������;@�6V�M�4�ҹa������n�et%֝��t
޵.cN{�^Ѯ��������D��0G�e�@F�� ��~m����>�·	�߳W}"�=w!
����V�Qdh/�w�'�p��-� ����o/�rj>쏬�S���ѻ����OE>�#�@����H��n9{sX[΢��<���Ar�An^�U1�Z7������x\�L]�����An-� ����E!X�w�TVy���X��t�_Ch �����;|+����5t��Y�o�Ss�D1�3rg�t�[�͵0 2Ȑ[�{�ŝ��@`�5~S�T�����"g2�*|0��� -��f�KB�_A��S�߿�G��x_P�l;M!cr`/7�YF�'%L�6x�RA���W6��u�O�������^'8ۙ�����ŷ��L�tsK�W���=��EPu樂:8��P?6�R�r`�d����F�:=qS�����s��K�_�}R1���{��U���F~�o�b�?g�����.���c~R��v]����K�@�3��WJǛ��(��A�A�=�����C��c:xm��L�����G�m �Ð������L���ۅ������� �K1���,�=�l�3�Gg�� �@_w2D��"�~�G��D6ڸ ��"ۙ���f�-~���SSG8��.ԑMV���:TZߧ���x� ����A��?7��|V�#�K�f�(��_	|�|�p�Mz ��D6�~n>Uv>�{?~O�O�:�Vm�&�VM^4l��54C�Sv���b�v��亹�f��>�Y>o��	����n �mH����̝�&s(��G�'��������"M�A��!�"A-�~�{t�w�Y�?O������կ���NyT͌��?�� �_ [���{;�V���q7S3z�� �z� �Œ$� A����s����5��F�x�5��GV�������Rǫ�Ef�������8"����3�9�R���'�H 	����tc7�9��*ϱ����C������ ����~y���<>��ْsx�h�!����1��S�Q��c��ޤ�rv������=����DǶ<���u^�ҳ��f��.Ӈ�%�v�7�V�K�7��f�����<��bM�
GtʕMn^�">K�~��'�R63]�K$�l]H�� 9&3󽝋S�x����$���~�Mr�>n]TŚ�{��N����ݽ�.�Ϟ�m�~#��/��U�t]�cf���%��0��л�8צ<U5�MӔ�l7ڠ����raͅ}����%r���6�a��Y�w�x/o��Ad☸~��~��O�f>�퇧!���擩+}M���/��O�nn[DL1쓠�r��yi�|�#�mZ&����9�Oc����S� ��M𳘳�̹�u����wE��|#�-:֟͝:R�O/�����j2�nl�cDF`*�Ӄ�� �1�<ۅ9�>�_(=�au���
��N�q!Z��Ťz�\<�J������ k��M���z������F�����i*���3�ۣ�粗c}�!�H�DP>�M<�K3��&�T����[�|�ׅk�GCs=�'�S��--�����]��CM���z�����J����/�x�'<��=�R��ac�۞���7�߼:w��=�@��}�q��]s�:�Q�l�s��p�j��߼`w�o�'F	��b��BK-�����˜�t��� �E�:T��BiQe:�[���{�f΍�`nY.T	$n	E�]F�%���B��'�!X���	�(�]�'dh����p����s���{����}TNH����[z�m�"2)d�V��J�Ew�	�k
F/Fb
�-h+��z�w���}�pN,�q�wl��ݬ�����,�B�[}�E:����E
�',�NU�'�$�#��8�S�"����U�
U�T���rn���yВR�QET*=��9z�B~:ہ�O����2!3�,Qo�>� �N�9�\�:�����C:��i�W9��"s�V�>����@F$�"
=c�E��\t�nWq(�-�<]�#��xwwV�Qa���9��i8y���@�� �S�N��u@��ϝ��X���ňC5��U:R&c�XV��-g����
��	6��8aS�y����Ke�Hf�b��Ř��dF��dAHDD�\���n��o��5�=_��Mz���p2���~̏�̉�J�ϡj��W��A��ԈɌ�9��t�d�U�2#� �o��D3׋��N*��w5���D6�~n ��h/�m�z�� ���}�)|�/�s�qt�iM���'=k�ƾ_�	m�q��kz<�,(�%��Bn`�V��	E��-�4v+tF�"r�R]��u���ٵ�E�A=�ܑ ���vi�������j��3,�z��I�DCƾ����#�mI7���^G���~=��Ɍ�0�~�Y�qVpȎ �|7�HЂ��%�4�L>�`���"Av2> �A Cn~�m}P}b���Tl�My�s���qq�����}�DfG��_fG��㱕��|�'W�'��r �h {sb#+���k���.A�נ"+	U��^�*F�D��9P�x�y��|�����_������ؽ���	����Q�W{R��ῧ���jI�e��-�=/z/&��BkН`����>���G��"��\��C<�Zg��s�j�I�<ވk��n$Z��½T���☩���i�d�S�2#�'jnb�����6{䉚;����.h��Q0Z_jy�.�j�8S�ݑ��[�쎭v�[�.p�[����� ���7� m��{2~��{�Oz˹�	^��\|t��=uib�����"3aK~S�����s 	���mC�[�{`h ���n�����5��w����� A��a��V���_�8��E���@7%��P�ɇ!+����I�S�2#�;P#s�,�Cp!�?Hb�ee/o��k��8g��mF�_O�{��m=�qs�^��������/mɨ�|3=�y[dH>�_@>�Vf�Ÿ��Yf���OL��r6�O����dW����p��b�O�[A|CnD�C���k�ar���2ܾ�;��CB�R=��ͫ�q�=��K�K��1{��[
�e����"Q�^�$���y���x�t�k�K��vIG�v�QOH ��*���͚��Hk��j1�9�&ZV\���8�ɤ��V9��ܶ�z	S)��Ͷ�;K	�s�[�fF
"���X�u�rv���uWl��ݭ�7k�w��.ق�ݸ�{^��mkR-v��a�cW�[�0+��{"uuF���]��a��'�����{��^M�1��գ��9�xzz���OiE{nn��䠺���g���^˯̍��}����~c��ۍ�+�@��7]���P���)v��zez��.�N���ȉQڣ��b�#�E�~-ʐ�Fn������S�0��vz�>���܄�Y��A1 �?O̳�wVi��!AT�u�����q�����\ֈ�Xz\p �v��2��n�V:>��w)q� ��[r$��Ш*u���ܢ��lM����w�	�e|A�����3�q@������T�,ߕǈD�%��Ԅ�3�����9�w�	ʀ-�3�GG�T���$����	��P ��mɸ�u��:�}gH�a{���qsZ#ް���8�Id2n�4������~zО�a��AH�*!D�qs��s���1��M�4�:�CF��.vm�?����>� ��~e��z�=F��޳Q���8�+Y��w���h";�~��dp9���f)0\G4^��q]f>遷��ڷ��9�7��0��%yy�v6n��F�)um��˫Y�2��x���t�1O����vS��v��z��ȯ�s.�tC\Nz���_�V��="�B 
���uϗ����
����%Np� ��}��$�Ϲy�P��z����v�<�<~n|CnD�">p�;ۃ��!Iާ�����ǽa�q��qڐFB �H���� �}���]/����#�`an�	
�~��!�ʪ�d���:*w뇠O�D�ѯt�~�>����O�d2���H mH �d"�D�3��z�8�Q�z#^��a�9���@@���ȐYe@m���f�bc�$��wX�e��SM�=M9��[��u�Z9x��Vj�����$x��A���܉���=�o5�y�\��{�!���̓�mN�G��@��Ŵ�C,�[���ib]���l�Dz�=|Σ^�o3\=]����?8沶���;��a�n+�.��\2n ��Yr�Ff�Є�ɘ�p�gj�v ;.����k��;����m�o�%�j$5����Dno��7��u;�Ί�y�@C�*"� +j*�Ggt �a��?@ ��7vp��32�g��*�R��p����1�3s��,�n�Ϳo;���z���������xG���ff�v�A�� �Z�Kp�6�H���A�q�է��EN �^^
����Q���dgH?8QcAۙ���b�ƹ��\k�od��}��$�9�&�Q�� �K,<r����k�A�"eJfbem8�A;�_3�{�� �ԥ���7;��s�����u�"�6�����Aet����@6��p4�'Ѩ��>2��H"��~;���M�o;���z��� 㹒2q����+u�;�TT�@��Gl A:�Bb� ��=|2i�s1��찫ލ�5'��,C����?cAۑ2���|[�u�����{��LZ����@�mDlfh���Z3�Y�"8�T�lR�g��*K�n��G{�~�tz��<�����?����?=h���}�����=�_����#�e�N9��_5����Fk�z2q������Wh���Ag~�z(�x�� ��!�ވi�A��>�ߜ���}��������X|_��	�j~ �_"�"	m����uT�Oa@BQJĦ;\��E��f7\���$��r�9�I��l�[��_��=��@@���%��͡��tT����kD�~ŝ>!���Z��~ƀ_��~!�!���S�"�q�aO���s��n��|ڑc3Dvwh`�O����@@��_2�U���Tt���y2(����m�?nk|�K͖�=m��Y���� �s�O��>n+�	m���|܄
�9�\S1��H�1� ��_-��gD���<+���̮���_3�*`\Z��.����ۀ�n��R��@��Xrk<OR
�iݕ"C|5gp����w��ʀ���� �C�L�g��=זw1���?�������*�飏�.������\�u���wf�T�N��s~�4�o��7�>2r�lG�۾���^�<��<Se����Q�TQ����������)�#�l�L�f�;���:z˷n{JiY��V
���@���vfe6�ؼ����@ݑ5t��u���Wc^L�n.�stW�8�M��=<��{v�s��LUu�휗$箱�G]N��ݻt��@b�u�-������B��9z�w��5d*�(Q4Z&�2�0ެ�E�v<�t�1/r�L��&;S�f����v3چ�Rg��?#�&����k�^�����4�qϮ���k�v�[V��ءlj]M�w���v���I��)r'�[���woc~����K�eM+��2"����@KmO�#�� @.�
�
�FJ�Z�}��Y�Ή��[+���̮H?+#���}[MeJ�Q���@�o9O��p��[i?x4�:�}�����µ膆s��8 NT#wdI���A|Cn~ ff]���I�c�H F������޵ݹ��?w���|\p"�Ɣ�iM�n�)x�f�
/!~.� ߂�n@n!���z�_���Z�U�_	�>�W.�}�fWH$VB����?[�Qobeaݽ7�
�10�lV�4qF���B��]���[���h��˵��+�"Tn���o��Odp�%���[��gp��s��8/��~��=p(]\�=������,���G�!��T��T(���h�~�.TFcɁ��h��j[�xS�T��!ϗ�fo�����F'��/=�_���B��ihͭ���D�" %���铞��sֿv�7���+�a�q�v���8����0��,A�j~?{P(G�\,@��ND�YD�=�>�D���os��Ͻ��}�d�	��D6�~e�Ÿ��,�>�^�˝�����{?��R���+7�1�g0~s��S���eTV��A�@���̳�mm���W�=7��n$�7����o��W�����S�!��-� ��"��#�������a�$�D��&�ut�0�d���N��]u.�N�j�n�6vm�>�}�U@_��OŖ~_6��v�h����ºO���-	�h�3�؂#1ȟ�m|�-�ȶԂ<<���wŀ�z�637�{��FDw��|��BAn{�Lg��@e��2����_f\�Qr(t�$�$�ve�sr\���)��W�k��?����C#ӡ��0sY�ްo�h��n���-�������^#��l"9} 2����G�;?g�}���������z{�[�|��E�q��<Ԃ5���mO�7�S�o��5��0���{  �	uݬ�j}�l����Np�@5�k���8��F�����>_�Ŷ���ȷ��h�Ћb�J]��f��sY�"8��ۛ"~-�DCЅG�s�wב�cͩP
QRP@��D�LH�\m�6�9���D��8��i���0�u�U���?K����Ph"r'���o��;����нt^����}�U���-���|�t A-��q�A��2�*3�uE�͏��W@��_-����g���\=�l�k /�-�q퓑#B�������<���) ����~m���]y��p�t+����k8dG| �͑ �mmȐv���qw�+�Z���������������|\q皒�LDFR���vE�y���/#�9W���M�o�����6h��D���-w����}�У%���wr<�t�������������$��(���zEQSZ���wW�{���d?�&� C3$H-�u�O�O.�6PKm�т}U��1\+���8�P� ��@�M}.���eUO�	�� �_�)u�3�;�㦹�󇭨�S��MX酒۩��L�L�[~y�?C�!� ~m�	dgoB��-泆�S���*��Cd��	ݑ �¾!�
�n�h��!��vl�:�PoE��u��FG��f�����V)�q��g��~�d [����,��:��a�$Y�n@_CnD��?6�=��~�!j��z�ݒb�V�=�"A"� ���"fH�~?��{�t��O�|A��#�$KmO�d=��Ĵ0fMg}��}�]y�*��U�z��7]�w��,���!�A9�ogw�dQf���v˺��J�S��%�) ��B�� 6���8S����/��9�=��'q�o�T^�2��k�^��׷���*�j�.0_id�:+}�ag=��n{��)�@�3V��zOcgے�{�|�)���������1���ƫ�3�9�2������yw-�H�������;��Pr���iM�
!0f���at=4��ǡ�s����y�����oyOg�(�}�-��N*�#o�vs$�v��gq����N��c��w���)wv�[��w��kya�{M�7��s;�/}�w
��׾��|��K���o��}�Խ���7u{�O���<��7͏t���݉�/g�o,D�v��n2�\�UgQ"Q��M���/�g��+�e�M�'i�s�w��i@�v5"�<�?I�*��ˌG�0�\�H�ʋX��>�ZjV]c�M��|�ŸUP-뛳�����\996�ۓ��֬�]��X˸5.=0�:�, ��I��}��:e��>��i  :b��b� �u{�{���+�Z^!1UW�5'��"w�����I�x�`xu��k�'��`��fj�썜#�8!�Y������a�Q�V��Sޅ^������v�g`�̞xA��X�=<���|E�b�/�~Uz�yH�
k��۷yxB��9�yd�ݺ��5HȘ>���YF(<��t��.w��������f������0OF��&�zq��V��n7y������C��Oe��7٥ÁYR�_7̞��?�|/9�V�׻;J�XCF�	�?�ţr�ǥ`8<�y<���Ԑ�y�m7D`t�3`�� �pp�Z�2�t^�>]�gw������~��}������U��g�$	Z]T(F���9� ��e6b���R	{2�᭽/"
۷`8 3���=�S���F~�:!���>g�{�FTbDQ�(���m�W5jвJ4���a�D�-���IQ�Q]ֻ��F�A�3��gdTUp�UAQTW��.\�g(�]�O�(=bQQDA��Q�"��EQ�+����i,*��9DQE��8y�QE��*ѠUE��z��G�ṭ�����zh�µ9Q:4*9QDQ�E��S�dU×'2�"�8���B9U������::UE����9d�Z�pw���)�juz�
�ݮ"Ir9DU�*�y,��G"�Oq"�3�U�E=�9y�^�UR�y����.uJJ"�#S��"��̉=A�D�|��\L�c.��s�p �ź�ݘͮD
3#�`��Y�U���Bh"�Ш�5�3����tӶx�.i���<�Z�=��88s�|R�k�n%*r��h�%ݧ�s�b*8�nʛ�c�lsE�\M��S��yn.�h"NXޗ��|����ٛp@�v�`�qB��\::9[�H@��2��y:�y��r��-�s-Fi.�@�i϶'���uZ��nvň��le�ݔz�^Ϧ�^xYݰ7ny��\����S�lh��������cs<ogi�$f+9��:�cM�k\BSE����8���4U�����p�F(m����GS�̉5Y�Wc. sX-���������6Б�Z��NT�m�{XF��2mMرn���ō�C�..�%���p=r���\�<��=�/|۪�Utb�%�Rjm��Q��MHTGJ)k,9�L��n�4sn�R��G���9���>v�n-����uAS� Պj��f�)�Z5�/-ۚ5�|��|P.��nq�y��b�{fyix9��n-��[�)�uZ�� ���8�eѺ�J�����sh�u������Y�GH��m��Sh-m홖X�.�&��܈�h`�Iɜqt�.���ӉEmǵ�;opӁk����n�C\��)|�ۮւŉ�q2:�=���rۇ��������ь�\��׋�@OW5L�pvjg���4�����=��@��-�jc��ٹ]���mY��:۷m1�x�������9�oI����؆����w7W<�R�K�MV8�AA0�lT��1,e�0�M�-Ֆ9���æ{t1���-�u��^:���,����A�k��玞:�ns����6�A���+�˺1ں��v'�S���3\u�%V�a��ز���'��k��E)�oW����qv�u�V�/�=g���ܙ9�Q�	����yjၽ�t)����xv����WOm��.E.&z��]iqn���ץ&�Wuw,��)�DT�{��j�]�\Z����֗�/d�caZ�'�z��b�֎�g�͜�]c���gK7=�6H���q��z]c7h��6�1��&�SY�+%&ep�$Hk�9���>����%Ǆ0�EGb�Ñ���ݒug;i6ݻy��J�-ד���[��h+L1,�3B��[Y,�X���f)W M�v�2毝)�x��q��'���٢j�h�� �P�w��w�������	����ׇ��y{]ź(��y����fu��*��	뀈��Ie��pY^��`����1\+��ޑ5�+�UL��� ~�A{��C�B�@�m�!�c �n-������?yƐO�T�������0fUg1� Fz��Ȑ=Tp,�'���X-�	��S�(���܉���!�����.�ۜ�W�ܻ��iU�|\q�� �2�[��m���`�e��
�N�o�p(��c����Am�Zk����鈮�o���h�_޹M�#�}뚽����$��~-�I�Ÿ��ؾ3�Ǘ*߽^Qo�nip�ʬц:��@���,�Am�3&2�ݓ�{A �O����V�PL�Ҙ���^լ���ƻr����.�Sn�1!��331�_J�Fjs?�����}.��b��A��~dc��9�� �_ s!Am�7�[�2�l9���h�߲��U�q�2�`P�p��u����?n��-�e^��z��|�����{�>j�����ß��/s����Fi'S�(�P��0�
���zN}��;��s�nG�����=»���k /��D6��q�4Ӌ�\�(�����.�N>RAm|�-��R"��=>���	�`�����T;�"~-�@�ṁ �go�//���A�@��<'�k����n�K��f������)!?v�8Ĳ��{G~�����ԀCp� �[����������
J=��ln�G������o���d �
6�~?�����9�ʛ%-�P_�n�F,l��]d�4�Fu� ,�kC)�]l��HEI�Q�ZXA��A��[� ����Fot.�����2#����ּ6�|Ai����Ar'��	���(dEU�cC̑?m|���c{r9�^2�����n�}8���9�C;2RHg��	��`9�����|A��}���)�����5��}��*� �W����$<��&g��=��Ⱦ�0������y3J�����r�|�I���7.歷5�B]���>~�> �������u��{뻪߇=�t@�uE��Ak���B�@���}�����J��W�p�ڈ����{C�0d�=��9p��x4��ޏ�3�Cn~-�_6���os�}9g��k�y�㽑���QT�_8�?]5$k�p� ��V=�����ڏ%q	S�vv�^j�.�t��g�㌷�n�w'�v6gn�e%�24��ꀈ#�Ȑ[�����E��z+�q���w۶��{��D��s��7s�~!��-����R���\�DO[�l# �9ܤ]�yos0����"8�9 �;;:���Ϸl&:�qnd� &�@���?���u��ђ��uƵ�w��*�*��p �~RA�q�-�8 a�'3�y�
9�������P���+�Am#3�y;������=���h�G��VY�9���{�2�`��&�ȸ�y�3���T�:����\q���X�tu���){�ݺ�x�q\���@�����xEE7�=�<�Zx�B�s�7j~ �៛����a����|v�OЮ7���r�`ʜ|0�@ �@@��Ie�HnFt��������X1V�@���s�l���L�0h���3Iq6sd5X�D(R�M�go��?'� Cn~��p�@{��{r9�f4������}���z�3ʾ#�H@�B���Re�In���1��a���A��^OA�{O5K��۶�G
x�6�.�G�{���{_}"���:�O��ᐋp�?ڹ��씂fI��>��N��X�a��� "��Ye|A�����P�N�ٞ�p����;�g��B���}���e��b��G|~��I�a�^�Qs����B?m�,�����,��<�R�[W�c=�����{8#���	���H&�E� �🋆D���W�MD�EvPSb�<:|�ٚ;R�]f-�[U�؍�:sF�ͣg����{ղ<�xj�����3�`E�5�t��~����~��w���y��0��zAE�g{��,�����l'	�vx8�����r\j�̻-3"BA����:j��WH�y��)e��u�B���}��mk�@�e��v���Ŧ��)�Ͷ��'L�%2��;���d(݇I��.�un:w;t�1�㜓q�3#�6ǳ�u�;r�h9�;��nP�N�����)�	���\SmxBm���]�/v:���攰c���.�>�?���g��sc���y�lXj����k^]2�E�mv������K�)>��ŸG����D-;|{gc�K'+��|��Jr.�q.� ��?� ����� ��p4�Gۙfs���#q���/V��gwٗ35���G��ԺI��ȷH}��'���$fB ����nD��6���o��y	*W*4�%�{�5�h���e��-�&e��W<�wy̼�@���!���o��G�ڑ�h��;���8������苡1v6�׽�{ w����/� ��D6������Fp����;�_*�ܸ���_��_8��U�����ʹ_����<���o奚x&�W�9��k�e�%w6�K�d��E9�.�����>�����=�B�D�[��n��-΅���u���Y�2�s�v����A�@�ݑ?��|[���2kp�S["������o}�Z��mJ���NnuQ3��9�ţ<��.�����Є��!5~�Lu�	e�\�p
��[Z}�z���:��s\��ֺ珀��EU�-��{K�=���!~9�~�\ʜ
q��yF��%�=���+_9.	��g����Av M��m�����ҝ=3���^�{�T��=��_�W���G���Z�~!��|p�?ڒ�����,��H�^S�0,�=}"n@@��
��:�ù�.�mg	Y1��۳춰����־@�KmH ��n!]ftd�{"خz	��"�w���$�c����A׳$�� �m
ܧ�N�XM����e4��S.뙬���'V��{o^�%#�A��ch6��v6��޿���?�2��?��I���[_Md��\޻���U��|�^�ؚ�������Dw.���>"1Ta��9a|s��AGg�s��^���g��� ~2�/�?y������]�{}/�ݶ��V����̶�fU�32�\��{O��p)Z�;�a��po���wm�+��?��ec�l�>�KF�r4Ys:�&��v}�vj�Ï�Ɔ���s��\^�ƫ��Q���+z�w�s8mpy5*s��� ��^ ���������~˽��J��sם�>�3)|n��[=�8W=�����n#�&}�!�S��t��5 v� E�"��]�@��[�7;;b=�D$����wZ��Eo�� L��� ����v�3��/p{c�>
*
�`I���`.�������냞�a�y���u6����[Nl��� �TX"~�@7`�B�w8��R�1�ȏ���n�fפkۨ@?k_n���h�@�f�ޓ"�����X�$O�_�����9¹�O��{qA|��҂$�w5,�=����gGd�ul:�mgt\"fYyRd�p.��$�}�+�U1�[��T�~���K(@�Aw!qd#B�|��1s���;���&,���bl@����^i���/&�Ncц8@%� ��o�s5��«ޠ�/�O^_�3�����^j���M��wp\z<fvT�&´�Q��x��#=x>C9Q'����c ��99���>�HD���y7.�,�fX@�l�@���F_��Ʈ���h����f�+�d��{�W����|��!�Dn�$�=�1��M�+��SA*t��ؼ�mF�N8��u��l�T:��v���&fR\ �} ��P<��l����Ș޸Ŝ=U��uJ������WXʖ�ݗ��Y&e6Lʲ��y�'Ԙ�1~"�\#��(X^i�ޏ9ɤ�1����A{���l�"+2Ĩ��,��6�<�_Y��"��h/�� g�i8��npv)�������#�ϡ C6B7q�7p��7��Wwhf�=�F�㥔A�AF硧��[}q�T�����2Y���|�t�opasm���h!S*��Sl&e�Lʲ���@���!Mv����5
s��~{� h{"Kp ��װF���պ��|")�L�*�vHǑ�s7���>|ޭ�R����)�_	���m�Y�孭Ȕ5��	���1��뽜���OH"(]��;�j�V��Z��'n��Mn��k���Z�记��U"9�P�GF�։&祺���*��XS�Y� A��
�ۣ�r��,#��F��[�Z3kV�m��ˌ�z�;O^��eT綳��Z�v^msWn7��-��w�ˡ��p=�x�;�����tj�f��^@94ݓ�%����Kgur���,�ێ��a��皴mcX��N�	������fB��ۋ;q�\{L��=<	���۴��n�˧UU*�5z�x���N���(��e7�m�����k�,��E_\G�A\ƚ�1�5N����w�XL%Jʲ��p�﹝1���K�=p{�C�y4�z���~�]��\Ah".�K�8�^�ϷZ�pȢ.���|��W��\NiKq�����fyTL�>�|^�_o@��D��@���k������"O�>_]��g�4v�s�s������a_`ǳ=}x�m����`�qC-���n�"���M@��1Bs_r�\��{޾�N�k�����<� E�}wOu��t��G4`A'�$t�11J���#lY��%�.m��r��]��me�n��]������?�C��}%�@�pa��sw��F�s���=�c�Ԣm���v _��z>� W�h�_]�Dg��^}ң��e9��uah���g�f�x|Ϻc�#=_�"K��ˢ�������)�V�¨<���E](�9UMӟ��?�����|>�C�!��n/�_�8~�\��LU��qϡ A���^;��-"��o�\@#r+�v���_]�v��5��l������=wג�Mw�|��p y�O�2���ZV�O��f����G�?�\ `��{�7{س�iNc�ٰ�����p��w�)��ˀ���#3(�L�,�eֶ^�F���;_k��;Ms��k=1W���"=Q?~Z��@��7qz��Z������<l�#��rF��W�6��[��u��Fh��i�K�
b4j�?8<_]���	��i��z���nf��8�~ܕ��V�`o�W@t�]�.�����#[:m���D�
2C�����A�9��Dq�6 �mn�Z~Dww�b��g/�'z��v�"�/��k��5y�§dzs������u�>��;�~�C��|J}e'Gwz,A\c�eў~ث.���ޞ�t>��r6������S��ݱw�.���q��E~�7π�[٩���57m�wAw��;o�ψj����q�o�q[��\��y�v&���m�DcR;�m��̚6KGb��K>w(4{ڙ��ϯ��p��ټL���{nc������ǌ{� �_�%6�i����D�y��ۜ���&���.�q>����
��Bz�ۨ�\�����F��|�k[��@��zO6�H��Ӟ��Ê�6;�cw���"���3����~�b��G����(q�O�w�ۥ�qW7ǧr�9��s���<ǔ^ת���F#<6} ��މ��w;ʯ;:/M���)�Q���܇�Ƌ@���R���V>Қ�[	�W�-���N�oou�C^ w/l���f/x"�^k���=��m��K�>�\�o��η�>��&	�/pwx���U��N���I���vJ�#�^�}��S�[��	��=�۴߫�]�~}���Ǧ���n�k��{��2���I$�x��n�m������ѬOU3&��񧺶����r�޶9��wz<����Q�kkw�/y��;ܷ�@qN��NR->�������x���g�|u�ޣA�oA���X3؟�=��y�_`�nV��u��I�%�׍�w=$ ��b�A�	�{Jo*w�L��)�Ү�Y��|{���_}r�Gxo	�*:̐M���]�r��������'�?O���ߗ��	EP H&�'/�bG"�Q[���t�ʖVb���dT:<�8�q������TW�M�D�G��E{3���^�;efI�8Q3ԯ~>?��ĳ~�F�YIG*�46��yT�Q�F[o��I��2�@	|�+1ӹ�rR�Ӝ�I3�HUEFesD��=YNe�Թ(����3*�B*�:�"T9�»T"�V�Ru��EQ���U%�tI0��NHDz W$�F�+Z{�xsP�V���I��%���r��H�W4�-S� �wAܪ�N�F�=Y�aDT��$W8U�.f�Z�)3·rN�djr��<���@8UU��y��Ur�:��]e�l�$�7S���tKCwZg��5 �֔EE�L��U��2ǘQr�%\�i�����oJHAQb�M�Z#��QJ9{6`PT*5E���AA�}q�O<�v��LU��~ �� C��w ]�!�'�C�o_?*�t;��8E��.�i��z�o�ڪ�� ~2�
�ߊQ��{�y�d3�{�2��eY�m��g����;����i���-7�ww{3���>� A���_E��]����WjƄ�:�&dX��1�'�"QaIz���Wt7���<�!�9��	a͆˞��U����0pqE�}f�]N�Gi�g�1g����q��^�ߣ#c�#���Y��� �軍�x]�|0���h.]��ͳ��}6׫����2Y_l��}��{����^}���!�/��g븢 @w[o;�*t'��3ٞ�4�1�� �lA���ٲ�pk�;O�D�e�.4G�����q��Z;��g�#3�j����_��י���Hz��KŜ�4���vlZ���~7��7�~�����c�:w�� �}�y��{�xC�8s�x��B��n����f�	�G:���yG�zA!�Q�u�B�j�.�L�,!�E̙?vfG�����xRAyy�]�.�|�������W�4i|n,�BB9l����{�*~�g��[�6&���[��!u�ݹ�7=H4h��])��������$7���������7p�l�݇7��~��>a�{TX����h s  Ah E�n�Ž�f=\�{�*��>���~���3�s3�)��8A��C��w4"�>��Q��m� p(������<<�⬾>�X�O�e�<������.��G��>���������� ��C�w�y��ٞ�|�1�Ȏ�� ̀�Cc+��]팩���@��-/��".�/������舞�Ϸc��~Y��3�s3�)��8��]��7p���V\�F.��ˌ��1%�9���N�]k9jۑz߁��
z����1���ڄ�5��3�h	r=�vo׆��I��C7p\�4������"��R�fy
�N������MλX7Y�i���W�'�r��eQ&l�V ۶���٢���]���Y����I-8�ks6ͦͻ>}�N�R^���<�s�[�ie���eu#TfE��Z��a�k6wBg��i�s&��+c-��񩚤*L&ʜ�h����4��؋Vw�8�w1d��)��u֨�oS� B
�m�__������:IaCu���� L��Ri��vu�u5vm��7;G4c�l~��r�2�@��_n�B;����~����~�|���J�"*��3�/�z�_������p��T�`�Ʈߴ�|�\A�fz�yecё8@ ��	����f�fH��ď��_x@�� ~8� AmE��v��>��0�!�묆W����gk#�S��3Q����7p���"���F�W�>"����Dv����Y�*�k�<���zc�p8�����ʾ�}z83P_z��Ҁi�}j̴���1t~���`�O�}��>y��+3FD��k�Ah9�-�К�Ǟ��%J32dD	���cT�tӌdŲ,��mc��뫫U�������%� ����_'���;�g�#�S��C	�͍S�� w/�������D��ח�ˇ%����Y��q��N��Fn�����{=����y*}�KM����^�yP�8�]No�r\䞧�H@F��I�T���#��g�^�U�?W}��.����7o'���چ������l/�?6�F�>@�ŌMq���b���f�<��4�/,���|o`/�-���Q���P��"<��W�質"��YP���q�ge�<����c�O�#�j��d�u,�Ml/�'\".� A ������f���`{_Gq��ޣ��v���A�ˏ�?z�!i|@�_w�ɨ�����GAr�-��Lvy�`��6�og[�R�4e��3.�.S*&U�>�(=Q���A���}#s77��W�����r8��u��wM�T��.s��fYz(̣A3�,�f��;pn'X���#=+k�vE���_Fy6=��;�	��A����~�}�	8wpd=}Q��Q��� ��7p ��+}�S�9:o���!ק�_�+"�Sv��b)��0p��]uwE��x��4f���"M{deLOg/ڃ(��Z�^~�fd�ʬ�~������@ g�圴m���e�w��?P �Z���]����;>�kf���.��	z� ��@FH�۝�O'�yefp9 ��@�#�Tze���r���Y̜s�_Zs-8�e��T���a1$��5��wy�����l�%��p����e�ix0|-7۳����U�u��I��+��b��K,�:-�]�%^y���]ř�~����{��Oגּ����AC��3�5�e�w�܇Rj�]I竣��w���u����|��w��{z%�y�z��t/��ם���/I����";�7���w�#�z_T�a�h F����������������g���v�^C��	��}��_z6�@���p������w���?w ���A�@���4e���.�~^�&\G�ܷ���T�@����v\<���ۛ�?X_�����=��=�ĭ��7z�4��l��uV@�@��6og65��~ɓ�J�A���/��^es���Tx��Hyݶ�4�w��|����w	/ŷ����:+�P����u��iefhȎ?^@@�ڐ4ZqZ��׵�І	�	����[�==<um��Ttv�G�0[��֝�J�/V���@f� ������]��i����+�����\�'7݊/7!3`Ȣ��b$��"7���4�X�\�m�]@@�;�B;���8m���>�\�\�.���&��!��j���@���!||`�}�3�Q�z&7�Hٿ�u�U��Dq}b��6�7p����  �I�l�z&�w�<Ez ̯��������u���B}q~��C�d�Cw��=�{`tX"�>@��D]�@�Ƃ�׻�1O��2�w�@X��.�r8{\��}�"�q�}h E��|E��b�i���c{.�s=ܗ�d����w͡�0� v�Ŷ=�?���w��y?d�03��s���bk�$q�w�Ny�8 ��g��:��]����L�ʦ4�����\�룢v������c+��[�,�0��n�k�8WgѱR�L�rO&���*t%�uk�uF�ڭͶ�ȗl����v�:�.��])���{v� yrqq�v�Y�nخ�g����Qh���=�����vn�4α�j=aeY�����9#,-Kn8�����<���|)K�m�1��Ꭽν�n�D������߮?��s���/�Eny� �\��4�Z�u�v���6��e�5�7Q��K���߹�#�3q@��#�_v��u�U�y�"8���m+6���y..  A�@]�@�wuZ�5�E§�}:����㗙}��L��B{qA3P�!���.����ȾD��uE�"����"�_�4�=��t��,e伬���P8ˀ�"�E��v�F��P��f�5q��;���@7q}�/xno'�G&�GQ��H�0���_��m�_ A��.�����[;��_)���z8vL��^��� Sp��7q��3�Þ�}}����=A��~��	C\ŢPԂ��fc��54M� 	]mZn�0X`-�\KtG��|�m�����p����������Ew�A���7&&�=��A�!v�F���r�+��ӤL�
Ы&�Vh�ү����I/��E}oPm3��������~�x,^>''h��i�1��9��+��I�*/��ty��s��?�}"B*=��I�up�=���}w�����ɧ�2#����A�����X?1s7���R����+Ve��j�Oz3c�ɓ���w��߽	��A��B��@]�|A7p���FN;�SN)����A���?]�����r����{N4"���\G&�����Ϡ]��_!i_bӸ3i�fO��GK �\�ȷ���}142i��������`�j�䕏�xHp�����܍�MV3X�ш7B�"�w;�������v��4�^���P"�]���|��8���;��>���;3;�9f�����<�s<�aUYNep�32����W^gz��"�/�Ǯ�n���Wq�]�Ι�"+� �@D�r�:�� -�;C��*�v��s}UǮj��l��ls*��q�׽еdLD��iԴ��⅍�=@���;��/��}�iU44��zQT���l���Ts+'1�["Т}�-ȶ�>4��������#<�o�LM�y�"?	�~mn�/� ]����FK��G��� �c���;�����h���s�˚w�Bz\q�G�y��2����ʲ��\3*��E��e��2���ر_f �Y��r�z�Og��s4W�-�]�e9��k�5�g^@��	�l%�V�$l����h���/<y볹��O2
BT�+kc��P�"�>@�� ��� e΍��t)��/8dG��C���{��AlE��k����������൞��}���_c��ۢ�ga��4��	��f;���2=�V�ጿ{��?iC?F~8����X%8�?]�[�sD��[57]�iM�TfH�pY&���̲�f[ls/�9��wם��ʃ�ˣ"�5HqDwt�{{�<��L��H�;N�B͎�ms�}��H�=�����ҡ��ދ\��v�����.�[��1�k)�f�p.�F�ܪ�;0FВ����Wv}�W����E\�����~7p6�"�"I���?]����sՂ"�������f�o�>ɦ��>qA3P���7q� ��fb?{:aŝ[��"�fT"�&dJ�q�]pv�SӃ�d�D� `hD�p�д7/��~��O�֜c-8�>�7����)��:#2D8GB%���� �������|n�~7p�����%^���"	�C���l���2#�&���m}w��f�]�`��"Z���.�_]��{I�����&�_x�7�݃�nn��f�|A�@]���".��^�p�ܫ�Q���@�.�_��E�#s���{��S�Έ�"3�@�p[.�}��;�/FZ������� ��D�� �������Z�������#��}�ю���y�"8@5����������g��L�Q��yL�5�E]zp�|��{޹}��&V��C� ��V��cC.ण���8�
�V�V��"V�ش8V�
�tQ\��а�y�/]>���.����L
�ǊPW��ɛ�������Y�ȗ���Y�޻�";sO��i�����ُ��yg�. ���g�Qf�s}�߹V"n�x�'�~��zd������j0]�o��o�Wx�\���}	��[��_����6����MaF\</�sM%�q{9=�>�-ܸ�[���Ic>��ܯ�����ُ�`� ;��[�ӰN���]�x? ��R�әݾ�u�G���X��Nv}�A�_p����=�w����}�9�8	�<l\��������h��wN�8f�=eֵ��q�fS�Äe��߉�%���Fz�)A��,�i��� 	F{YB]� �(���<�G�ѯ��t�ά_�n�#ñ�9�ُޭ�Z�:��ڽ�� ��_?y�� �J;ˇp���tL�����V,(b��&�j�z��5���]W����{<����om�t�xw&{�h��|���)p �Z���0�8�l]�Sٺ��;�̜�������w��8������G��μ������Q�9�D�L��0^ïع�>;eu�G�+(v��57�����t_M��E�ｌڰ=���h�jY�6�W�0�n��m�x����wc��٠�Ǿw��rg?6o�Ў;Bܷ�z��;ƽ�Kק��i����};|�������o�7�z���l�����7���AD4@ń�<~����'����R�':�w"�<�V�FB�B��'q+��sD�S�$q����G��7�f(���V��(�B$�Br]�J��#��{��y�j#�����~e\��eh\�JiGuu�����%
=D���E��vT���	Oϝ���(��"�wr�:9�ꦺ�Ր�T�	�U��YY�"�*NV�s���9�L�*�YFIZ,4rv�2W>��|�(�!V�{��g��p�G��B�(��k�y�t������%r��%%U
�8TEU�	����+�%�Y.B��9c���bXW�׫�UIa�T^I:%r���Tr�GA���
�r)�]qZA�e��EW�ȧP����Qw\�E2	�<��|\����T�Ȳ�@pO%��{���[��Y`W���8	�	��I���Q@2�tr&Z3j��Q��J<��l���次8�7�,z8�]Y	8�$�m��IR\�,���x������[��.�ꭼ�A�э��9IR"�m����cg�1AѦܦۢ\�s�TP�Xit
�ZJ�l�:Wi�Q�r��p�]��G�����l�X���\0�gh�!�GB�nՄ2����!�Ƚ+r�]v�4��8�.���r:�U�^�-�������5���ðWL�ۍg�N��j�JF��yƷF.!�]O;��W|���ue� �]X��z�����3ۉ��F��m�]�@Z�%��-�[Wv�:��:YY�v�R嘲1�4�ה������H�K`��qť�m� �ų,�f�a�����6������B�5�R�H�t��7]Y����}�(�,���{s ��yk0lq���]��[��\6f2��T��Z��z��su�3}���#��pc��;X�h�2I��p��i�,d;G]��S�� ��	�0=l�>5��wby5u�qn�8�SqѶ̸��X� v�Xz�Z�=f�VSs��h	#�1U[v��p��u�qv�&�T�VWh�CY�D�k]lJF�4�[����fMҪ�ZX�L�i�U�VVS�����,�0%J��e�Y�hCC&�	p�
�1n��+
պ�c�ώ&Phڷ��ͻ(G�f��1����C:�� {q�વc�l-v�,i5]f�,��^����cLV0i{ZE���ψ%��9zF�WHu����L�q�e'�rϭ�|/k����4��
wwlM��h���M�^�Ss6��<��:��s͡#�m��4�1�(�2��<i�m��f�.m\�m`�xݓ�N.z��P��F^g��ݥ՚�2�J#����M��,��8J��j�ޭlH��i��2��u�sq�d�_I-��*]�7���'�������v��s�=�k���k]LEH]��MO]u%��d"���C�w���E�ԩ�`�L�ҁkc5��77͆��#v֊�κ�j��6Չ��Ȟ��g�E(�<���=�c��Ѐ���ɦ�秡����xu�:�f�;#Ӟ:�6�ڋݵqA�[��ʩZ��l��.G8+��-�׳tS�`���u��Xe���d�8K4���ȳR�^ͱeF@���͎�%�!���oZV��T��\�s�ٷ~�����}����r��6�`SZ�{X���ֈ�1ζ�I�q�:�U�>��<��ﮠ�_v���>C�^�j��>ɦ��>q�`���|�z��K9E�G�w ]���X ��e��.#7���A�A{�ns�����gDc��e�@�v�]��tfc}�I4��5 �;��?f��`��Z^`��u�߽,>�+��z=��٨�u�2#���m�����7h�B|��>���$��4���.����r5��O�ϒz�8A����->�9g;+=�[��^B"���D���p'���5T
���rwk�W��9FzDg/�� �.�_6�_������w�w���ft� �����)BR�����r����{y�d��'Z�ι�k����o���_~���"7p�ӯ��sF:Mau�2#�ʺ+݃E7Q��{||⁐A��D�}p���N��uXvh2o��6���z��콒��xc��Jz_��_j�I��j�\��/7�Kл��Ј�}�����8s� G�$?|G�>C�}�}ۑ����O��$��q�U!��@��I������aBfB�����@��
�
��g�+Sq�
�O���{3�fs�1@�.�n�@������������Bhf�� ��b����p�N�����kVpȏ����1۾\��!Ǝ9P fYl3-�32�a�E�39�<w;�y����.�c�g�L��҇��U�#w~7q�pguO@+�0A!([��D$�W��:�o\D"41�M1t`��-�`IJDx`Q t��=�� ݤH���{�}���9�� �[�Ω53�����?@�A�@gG�.���� �w�=���«���w�q� �n�G܇���SȬ��@h#w��nt�V��z��w`".�".������ñnܼ��3�������TLٱ���+����L��J/�߽��(�~� ��d|-9��j�}<Pb\E�A��~�����\2g�.�>ȏ�$㊲:����&�e[wߘe\�q��*�"�]�Q����>������������D���#;��ݷ3*��U�������vV�ߓ|3+/kD��[!��f�E.�k8d@
`qy����p=�X=�+��S�Ik�>��P�h�y��61 ہv�`Y0��qٗn����L� D
J����z!�E�|���p��׺�eO�](}�$@>�O�˭�\[ds*�BfS�\#3(�$W�xDe�CU�[:,�#�`�/�t;s�5�}��ɜ��Z�'�A��;F�!ܾ_�@�8�]�.���N7��0/<}nhM�y%��>�5}h/��A�A.�{^�ˇ�ں��u� � ��KA�k��[�ϵpʟ\�P�";�	����z��QU~���<���ֳ����+�S�[�vC�#��� 5�ad)V���x]q^Cgo�20�ó���\'�~Zy{	�+�f?~ ���?A{w ]�p,�v=���N���/�l^���\*�{�N]����.�_]��{���=�Ϲ�|��t|��-ʙ�R�<���6ܬm�kv�H�\���6km�_�}?Є��z��� ��@��/�ӏw����a��">��5���u������#ފ@=� ���
���@��u��0�k FZ��|��u�o���}� L�����s��lx0}���P������Ah@��g�{$��2�;��T�݊r�b��\ ��A.�����(���z^��ACME�n>@p�&�Ct����.g�i�Ȏ������9�>�E-�΀�"� @7p ��u��t�=U:��	}�>��}�)[����'7����U����`�a���jޏ6n����_��U+c���w\����=5�[�T��;�:�:����Y�������~voG�~��z��<��BF_i�����ae1v�siVm+��C�b���u��nͼ��q1�#�� ��q�8{L�;[���nTc�;wK�'<lJ^�w��5���z�nB56�x�
C�7j0��s�{:�.ȼ���i�c؍�a1��I�u+m�>7Gg:)e�֮*�
˳nȦ���R�g�V��y��;�+��J*�8뭞��T3L�V�'��'��]a)i�Ŏ���%v������e1F���tZ�[U���'���!8���������d_f��4�݊r�b�1�=��~p~̻�?�|G� �7h����"'�`wV�����D�4;Ky�X���"����P ݠ���2��;�S���A���2�/�?]��i|@�_`�	Z���Wң1�~�F`ʹn�'���� �wP7p�"� ��o�t�+:s*�h/���AF�כ�4�݊q���}.;�v��ڑ�B4��k_!B.�H �� �n�����K�okb�+E�wЃC{�{y����"�� �@_�������w�q��e��|O�;rE2���#m�=�A�ku[�O:�$��v�32�f;����F��_]���Y{{�/��D������v�Jk���+?!���x�e�6�_紒}%,�2����,�~wy��x�]�䝗�Wa���~��p���������|,��_%�W���j��������R������A}���b=�;�v*̡�ph E�Ug����,��H@�v�F�>@�q��<�𛕏n="�c��Qk]�E>�5 /�����v�a��Yލ��N{�4�ւ�`=�!����}٫�\�u	>ȁ�x� ��3�G_��h9�_0��*�VB2�a�-��s�s9��S��+��7�p�tGx��z�2F.��4[	�eQ�v�̷Tj�M�~-�����Hˈň�V�w5"1�uf�F��v܏5��{W0v�ֹ�65]���?��Q��@]�	���m�=����dS�@����9���n�]�@��HD.�D]�������Υ�3�բ�<�_���<���\1��ta�Dp �uv�@��Ϫ�j#�ɑ�k������ +�7p�]���N�Gi��ƏG�ʮ4��Ӟ���
w}SZ����އ=���i��^x�3����e~��6�,��B�hʋ�������K����]��#��2�/�7h".�_����w�9WL�Mn��G���p� �w��ݸ�ۼQOFDq�5 d��ۧ~������ A������ �h E�ϲZN�m:�ϲ��B��ww5p�t����uC��7p�&�)�tKo�>�����WrfW��֫��[���k�c���Qm`ٴ�1n��?�q��V1��^��A�@�v���x�{��#"�d>�~I�/�2��we���m̦�fU�`�����繨���r �}q�:�<��F{�E^~Ҧ5#� |C���Xd�Zm��A E4�`��_/��_:F=5�J)��Yg:�	�Dw���/�!���Dwn<���O�[�6�@��� �v��u'�k����Y�1w�����/6'b6�uđO2\�'�Y�>E�a��p.�=�'���R���N=l��n�}��c�݃e�o~��^ο�/�X��S����u�Q�W�\BvM���A���>S״�L�nfSy��J}�m�{t0|�Z�����QO�Dq�@D�h �A�Bz\8'�﯂{�i��[t�خ��5�� p��[!l�ø��6�i:���v1v����|��K������_�_.톞�o]F7�M�}�C���F*�o�A�U���n��>�� �n�""l,-��ހ��wn���+����fH��9�h".�q�]���y��9�g~S�O7�l#2����$���3n�*.��d\m�(��"8�f� G���8ߐ�#ܱ�����5�^ �$��_]Ă'{�?o.��~�r_�p?]� ����S3%q(��t#�d".�~7p �v���l6͚�5V"���Vh؞��̑��?�����i|.����c����G�Г3�j�j�"�3ba�~%n�n��L�K�}����<)�DN�a��u�u�E������\��;��I�2��C�MS�j��l�w�Z]������љ:=��n{��ē�M�)�({.xҧ)�-�m�6r;��=.x�j��у����QƻOOcHbZ^���ݢ�xgl^�4ol�ڥǓ�����y�FN"���]�4U��\`J�وiM��I�m�#���l"�����t��.��Z�N,Cs�3y�ݵv����7C��RnΡ	�h�3�-Շ�?�O�����ґ-�
hb6D�9�۷mE�r�q�g�D���t�}��B�W��w|A7i���{���w�<�dG��k��s�Ӌ`a��@D��D]�&� �ڴ�KN/�n$�&���|�wo9oug��w%����>�"�������D<�`�]BVB{w|n�v��9^���c�c�lK~{�s$b��2�"�i|n���@�R���4��rq�z �� ��p8{���F��^z;RGA�o�(����k���p����.��� ݠ��Q���V��W������V�y���_���B ��|�� A7q�å�(ر�4u"m&.l7�B����+RJ�����N�[�0�#��d. � ����G�hJ��k0lO?>�9�1r=S���L{���S� a�Gr_��n>@����/��*����)���W�lCTMz��$ɬ
ac�(�^ޓ���Z�nחw���_��R��e��8�=�"��ZzN9�����L������w�y��8�\��n�s��ڭ]n}�����|�� ]����_+G�k�A�>Y�&z`�?rř�λ���������fZ~b҆Z~�����B��@�́ �p,쀈"�1n����<<����H������=O:�г���A|C��7p��� ����)�˚�7US�'ކ�*.'�wǻ���^��>��?z�F��3oJ�M���L"bLĉ0&`L��x����:���Q˩�CJ��6���K4?^??�����w@���_��˳K�Ν���;��/���{׳rY�,�|1��|/�J�.�|�p{>yֹ�*84��7`/��;��T���gD�H��e�_�h".�kѺ� ��~�������wa.�����s����t("dH���Ju�d�z
-����nA=�	����D�
�����)E!Wg5����S{P�o��]��;�4���{�V���f��*vv�=�����jd;�nH��Ǟ�D��UC���A������s\��aJjy�pۣL������z�wQ��NbŤ�e	��2�G�W�	�?*��Y���o�����}�{���sЊXHw����ɽm|z��oe�\���b|H{��8_�����G��d�;�)񇻞�fz�x�_��%�w�<�g�g�ob��;�{y��}~x�W^�\��������Xw�u�Z��^$�{V�:k�xѾ���)g�iqoѽǩ��G��#�E�\���~��=f�SB����E�1�e���E㿊ǐ��h}���g��u�w��ao���'��cGo�z
(��� L�=�ǳ۵���> 7���{=�|Ѽ�^��_^��{'>�Evu�3���q�_}��ޙ�R�v���W����^��6���
4��ⷮi�{�8L��y�_�m�&K1�1a��иK�|�-�H���ۯ;�����=���S�^j+����Yq���{��wO[���\}�4��}�_$ӛ,7@<�]�xv�%w\�	:�Nzi�3u?S
�o���A�5zb����sŗ��XǨ#�������J���Q�Ob�W��k+�������z�����SN?o��Z�k8Q�6�%;B����U9�����+�"�+�<%@��#!�`߇�_p�ׄc�=��~ �|2��ݯ��jq5$w��K��u%i�Bl���:�9��.r�ͅ�付n'�����.�%q���G����	&@��g��Ԩ~�.WԊz��P^��DA^8���~?;��\T,���PI
rir�ER��Z��Y/�YG|���"���>u2�RĪ)R(�9y;���&I�-Bҋ�8{�./]�a�B�2�A-�Jr�B�3[�����S1ww*�9	��!��\K���<�N�t��R��uХ3]p�/"KqCC�m�!�%#HG�����z4<�縗9s=��9�t,�U�D�$�5�����uYNv�,S
��ˤSV�Yr�G,��;�x�Q�23�q�&��/A%����q�E\�G%iQr�1�<=��r�T�(���S�fE���8@ 7���]+�y
�Dg������]�D]�=z��31�f��@��!�폮����k=�:��ז�_dG�_z���(Ι8�w�ʅ��]� A7p�E��wb��:h�%��k������ݝ�F._K�� �v�]���}�.��D����#������F�r�E]U&���eՌ�e�T�3b��Gku�_o���x�|�f����~7P���K�5�=�p��dG|F�.�d�k�SH"ms  Ah/��_ M�G��͙MU�y�tK_{#��5��[��m�X�Ȏ ��Tv�_7����z/�v�������Q쀁��?]��F7��G��E�S��O$b��ˀ�7h�����}".�A�O���������8� ��X���{=K����A�@@�g��n�E��8�3���O"�D�䳈�)��� �8��;�9I�u��>�l�z�{�Z^�<o�����SU֝�w~�C�����m������>z���|A�@�� ��q ��]��ʟ������~=�s?ӏ�n{uV-�p.��-�.��p]�Ƿ�I�a߇c
��Xic�0����mW]I��(�q��2˂��9�T�1R�8+���A�@@�v���@�v����`����ОH��3�ŘFD@��C�>_v�C�[�� A��x���x��kЏ��b�v���]�p��dG	�@y������ٽqf��e���Y	�[fYd3,�2�(�fR�;f"�Z=�:�+1�5b��p ��]���� �n�wG�^�G�Fgt$������	��{X���Я$b�	� *� ז�``�i|F5��iX>����W��!-�wu~����6(��=�ӵ�����~�@@�����BH��B��7&Nh���R2(6�ں��R
���؈"�ƯZgeJ�~�.wvG����ީ�e�{j�����9.�뗷���(iv����o����N��B���Ǝ��Ʊ5˵A�Ϯd�����氻v�^�C`�w9��6���a�+��.����p��pɥٵ��y۪.4t���a۞����z�L1F�U3{��(�mp==��<m�g��e3�	[z���x�[;�7^űr�z�V�G���7W�9s�W����3�������d�.l���ڍ�g��Z�Q�����f#�Yfv��{�}���J�ؼ��shĕ7k.̸p\	��T�͞�W�*��n�M}����x� !�w_/��_'Ù�݊���n}b��p"��ul����Vb��Ȳ����&�>����
ֺ}sG�u��=5/�"Zz�V����t+��8p����yV��٬��ԾF�#�� A�@]��b����<�n<d��7l�OV8O�2#�!���� �6�7p�]�D]�]:�,��w@<c�}A|@m|��/�N��fS��7�#�&� ��'�֪=qDL��;��9P� �� 7��D��	]#�#��^�r'�~�/B���}�
�Dg��i@DZw/����bnrs#�`(ѝ�7+rW�s��<B��v�L*���yz���u��kv~���!��C���x��~��>َ�3���S���B�����Gj��Dv�]���r�>Y��g�T�P�����e�"|*Q���J�c^δN���}x{�g,���=��}��b��/�]����}���ȝ͜������H�K���_o��n����N��oNG�b�C�����f����͛�Dp9ĐM�[Aw�C<'=�Q��**�W�Fq�<�*��h��h�k(�fYne6�2�7���c����GB�ذF��O��@������;��N�2��dGO�oI�;��o������|@�A�p�e�j�ɿ8%k<.��e裏��v����%c�u�7�#� �@��돨��Ov��گ$(��(D�"�H�B�����v�w���� ��$�uV�]k����?g���P �_]��A�AfOBy�ytz_gB���_i��N�~ א_�A|n��w ]�ֺ�M�ޚ�[�3;~>�C�u��܎��Hi����A3ph#w�$�_vʆ����
s�@�㘻�!�����f�>�����乶���;���,��'��{�iCܮ�L��Z��xK�r`9F�joH�2n��nSb2f}ps���+m�^仯Y�ȏ��k!|Av�F��n�?�qDh��sp\EΚ�왁`�\s`"�h'�Оd]��Я$Fp@�p!4�5�;�H�� ��_ n��n�|E�|��8[�lFſ�Ď�X\�������L�Av���(�-�ބܽ��>��K�6��@�6�v}��Qv�a�gGP;�k/X�v)SFkuؿ{��K��)>�e��i|E��}�4wf����.��o�#�!mWٴq������^ۏ A�_/�l"�����➼��=�Tr�7��<�<�=7�Я,FwӍ	?7s�a%[���Q���yw"�л���'��HM�]���zU�L7Y�4�g��7�]��]��4����)�T�sz�~��ѣ�622_yN������]����b�
��}�=��{q�|�����Ł�:W�ד%�����x{��w��, )�PŔ���$��r����	� �w^��w_]��qwe���F*��W��o��q^Ý�v��~��pݹT"�8��>��}��
S<8�]2��Қ%٭����=�Xѷ+b���D̈	Jf&Q�|�}���|.��Gt���A����G�k8����ok���ݯ�Lr�q�5\�ˠ
�C8p�úv_b���-� K���w�}����\�r{:���wwt�a�6F!lU��Z�(�y�N��wqwk��s$[r�o�/�*�x�O/�c��;�7�xv�1���	���7Ar�g{(j�^��!�.����r�'7�F�#ݢk��Ѹ�x�]�6�������+��]�k��S��u�;��b���7������C����h�}�'����g	�ћ�D�=��R��ȶ�>�&܀{7���i����k�tgEH���]Z����n+;4�P�a���2k M�<��v�^��/s~�U��l�4v녷������ý����{Xc'j�
�l��*O�n���a�XF�9�p������o�r��Ì�Z�E*HC�n���b���]��b��u�ۤU�}'1���a�YfiKq\X����c6����1۵�/�3�3��fQѺ�'1Ʋ�����LY�v������}�`�q5"�m\��X����.�*2����1R��~P>ˋ�_]���e7�м���(�9à�5���n�`�_pm|��˼f|�r,�e	q��1����A�v{��|�������or�UY\8M��޻����{#^�Qol><��~���'?r������ߔW���=����7�&� ��K0����Ý���Cڪ�vl|껀.��wwxu���j{:���ɗ�}��N��]@����M�V��3��	 �
&!H��R����WLYu%�St�£fщƹ��u��m$��_o���H�]�w/���_NL[�݇�B�5�]�܃p>��.��&����k�h���Z���f1�/�����s99�N���>j5(9���|�v�Wc���C�����~�m������t�4�9��[�Q8r����GH��Pm�w�\gG����qve)s<r�9ݢ<�lϘ��A��=������v��}wa4'0W{^d��n}n�
���_F���&�݇�'e�l�ʋ�������N��w�]��ܹ�����J�^H鷜���-|.�]��ۯU����m���ܟ��Sܡ
��k��q�tF���@��6���l٦*-ұj����g���/����}w���t�p�x�t��g�Ab���%�Hs���i̶������w��T�:zc����p�-��d��S���}vh��-B���������]�����=u$/�ǋ6:g���A'���J	���2};�vK�#�m�;@�;�|)(��B�)Jy���TW�z���V�%^V��	����"i~���w�o{���Nл����wwu�}+�.傻�8��)j���x��v{��=^�� ��W6=>Wx��p>�����S�/+�ˈzw_b���@N�+��]��'&�?�s����'��z�kVlM�Z$�ḣ�[ScPcҽk�G����|�ޟ?���=��,q��4�=�g�<��{�9�� ���~7�-�-9lW$��������CC)r���x��v{���}�����&n/��r�%�_[��y]�������3���0�a�y�F_��=	�ܮ�����Fdw�K�3�b ��m|�nq���
zS��a�;^u�--��q�&v).�m��K�q�y,�|��~F��e��S��[��PԜ��꘡��cb�V�ۉZ_�7�oq�����.���W~���;���yrͬ��g�v{�����j�g�߇�� 	G���:��rЎ}��3�H�e�wE9K�ahG`��	g��p=����@f��A�;��H��݇��k5��M�/���]��\b�Q���ݿ�����
zS��a�	��]���(�v��oU���}ށ��B����/��W?O4.EJ���xCt�������W�]����vr�l���>�O�Ȼ�;� ��ؤe�n����C���X3�}��wB��}w|6������iC�8b�K«e;ވ��b]��p��}�#q��+��//N/���h9�2����j��jO%X������Uc�+�i]����|ܤ"�u��a/��߯��8�I�扞�.�_�5���֮�Gy1���w����E�o�L�3̤���`C�yZ����]7��r{llr~��I��9��"#(��eͬ
J�P���mg�s�>Y���}ǣRxc�y���2��9�����l��)�	JFkU��i�>��vK�� ��+i�Z����-��o]Y��$Lg�fB��ǀ��`��̙д��+��}}����iȣ�7���&�� �{��0�KP���cE�u�����±�#2��r��&���_�FfW�N�D,7�s�G�VײpL?y�(���t���/e���
Z�lZn7���o�{q^��K��av\Q�ϸڥY��w}oL��(a��;WN�e[U�s�v�t���_���w����p�ךǬ���`S�W����&�n{��8Ӿ����������6��� <���gf�ɮ���ӽÞ��}G�Bq8=������3�/�����^a�^��;����`��O
��A�<���J�9�;{"�Y�[��aٯVD�1��I朵�V���7Z���E�}2�f��z�@�,M��+y.��	����_���d~�rg���S��2W�0��(Γ�k{f�{�H{�\쫽�����c��@��F��Y��]8�Tؐ{��]��B~cq���m�c�����K��#��]���c�w�$�=���ѭ�h>����-�'^[=�br@��m������ة#Vx���xM���慞�Pkzn������_i=УX���z�^���~-ţ�8B�N���D�4�c�P�x,�O���z��GG�Ndp�G"���V^d;�E����y��Rr�͞�?������ߨI'�Y.Q�s�U谢�W%P4JT��K��eG.QE'h�
��p���$^�(�B�y�"��bQWQ.\��u�Np�T|ʊ��9 yN�TDUÔQ��|{��Iݘ����B�������X��s��(�ueU\���+r�Μ�7::ӏx��r.b�ݪ	ӥ&�8I���u�T=hNdG��YW|��6D	��q|�i\�U〯<J��C�1�Sy�u[r��s�9�S�(r�w2(|��� ��x�r�(�nM�� ����U�a�By8�ʠ�洵"2�x�B�|ϻhKevu3VZ��4���L;��GmM�:��m�'�J[�b�nx�h#R�[5�MJŽ�)'���p��ʇC�8���s�a�<�i�q�i��5�Gj�e�).c�s�6jX�Y��$5��oV.ypZ�Ű��-��m�l�n*Ն��lpsCTV-nwk���(DX�\�Yj��J�l�{X-�{V�ڥ�p�xx��6�˲E�e�s�6��눶d��ړ$�q��D"*J��"ę��ųS��,���q����2��5����y��:���t� 饌,��f��k7"\�8:�����h�<\g����7^KC�M4rfkX�5fq,�5���5�$�K�Nn���f�U�F���fwF����}�w
�Jfv4��Y����.Y���e�!WY���i]&5�l����bh�W0ڍ��e�
�f�fQ���-��/�_�g�'j��i3W���v�s�ϝ�vz�M5Y�`@af7��#��ؚML�mia+�iJ��^sؗEtc+bG]��>��9�]�Z����Ȑ�����[�;9��<�rJz�'��N����y�C*q��Q��8-�89��[X���5Rl�ٴZJ��eɉ��r����!�i��Ց�g�S�0��[�Vm�]h�^��g�'�b@�;c�m������Κ<��\����vA����B�uƚTM՚�,��Й�s-ݺ8�\�\�S�-wa�v�;F#F��&��6���`���j�[4�V���=�mҺ;Fr��]z�N�Oi+.�D�ࣲa�g���q�17e�}�1S5u�6D��#�R��l&�x;X��uss��9�m�hL���X�i�pm f�<�5��eۛ����\���umPņ;[�;���.�&D�gmgB�{F�9�^�aB�+��X��U̞���pA��@r�\ۆ�vF5ƚ��OM��ݣ��t]\��m�Y.6m��v�≤\�]�$��6彦�ՠ��⑖ݮ���m��˧=��`b���ڮ^Ԗ��n-Øx�g��I<O��li@4�tlDm�r�cj�ؘ���<����ez����#,Wl���k�gf��%���5��k��i�7H"S���0�si�lU͌5��V���\=q'�^6����=Q���qv���������WIc�+��,�p��u��Y��:�A7�gq�y���s���}�뇏���ؖ�b�-�\7���'dV�����	L���
��⻫����t�x�"��?�������:w�H~���M����ף�7Y�n �j�;�8��#/�v΅ǧ��M$&��?����y���r���}vm��M{�N�y��y��*�S����pN����Eݠ.��x+�6cDq�PVUU��ػ�C<�t�z3CȷN�w��-b��=����.��Wq��C�h�ř�E���U��c8���#/�vΧ��Wp��e�}��p�%L-����ify� �ͧ� s�᭄�5�;a�Z�-�?���6����wDKg9Et˽�Ü���.PV_`돳�}wh]����!�ޙo�D�˝<1±�K��'w��}<��y)��.<�e׳xg��Z=��;���=�#��M}�􌯚�I_�!�~�R����嫧�ڎ<V������K���lT�}D�~���C�w#뻸����&��x��g������+��]���&M�:ＡFy�r���	��q����U�2�x��|�:�,��$��M80O߭Zrھ����?V=( �q�^]/6�חN���۹����	���yJ���|�ȑ%)&D�"�0<&d��<���Ck6;=�m=��j�5y��i�}���~ ]�v�z;�Fq�}�G��v��a�*�7A�}s�Y)̴�e����_����Z���؇/*�w�b�;B�.��dr�)��{\]ڻ�v�5����#^����+=5q�s=�8`,�~����w.<l�W�����<�>�ڷ���/^�B��ye��9���o��%�1�yv�u+��|�����O��j�.��UW1����ہwhv�у8�ɟFzn���	hp��&v��~�'hs��t}whz�}ww{�ﻡpQ�ȃ0��6�T�Jw�b�'h���]�A�׳�{~�-����}�пқ�U#M�u��9�Gu��&�JMu�<�B� ������D�D�lϻg��֜���\�{:�feӧg�����ң���;yw�>���Y���~�ʱ�06�|�V��ѷ����g@W`!�&�c�}7�����.>qwk�gac(r��`�	\G���I;�1x_|�������л��NNcv�܈���}�vt�.�θY�t������r���N�N�է@Z��ZC^
7a��{n��.�(�ٗ9U�T�:^d*{+Nx)�E)�D�PװN�auB7��@n��p����x���a�?s��՜�Ep�{��e/Fzn�" W_�]�z���_&����'���TM"�]`���ޭ֌kx��.�Հ+[1,$SA�&R��f,\���3���n�C��vz�;�1x_~�A����Q|��G�����o���=w��w}���g@�=���gOr�����]��e����_�vM��G����|���.���ã���W��r6lT_+y����vί@+M�ڱ,���S;���~��֟�ߢ<S�x{�/��g{��3T�i�ӱ�U�}��}wk뼯wQ��;"����>�k'wM��~r��}��򸻵��޾��d���Z�ߋ����oM���?��;�8)����L-9VZ���)%��ݴ ��>:"^G;�}�ñ��/���q�my��a��_2d��E�u��1�[�M��j��躥�f."�Ջ����݌M��w޷�2��F�Gv���o<��X����f�b�P�b�X=f����q���[]M���񩌻��\����[��ܬ��#��r(�颅���q�����i�M����\�v���.��K#������h[].go�f�7;�2�[.�خh}�?�O���6�lL�طG9�Ƹ�#elZD�c�{nf�r�]��<���߯
u�@���z+4dv��e/b��g~�Gޢ�=v�K�m�ݏ�����U闳�9^p��}���f)ٞ��������ZU�\���l{��yO�rھ����#�#En�����v�,�c-=˷.�pq�˻���r��PM���x��	�}#��΀.�|�Vp9�k{){.f�
�Ё��މ�~q��06���]ݻ��h����FODm^�����!��B��������$!9���b<
/��7n����Jn��Rqv�K[��3�'l�n阙G�#_+�p!�Z�{�7�m^�/=V�I�����ww ]�Kv�bgqH{�O��=Y=�4���ϗGA���K�4(�G�IgC9ض�ÊU/ ���R/�Sb��LnԊ�{ZR�T#U�\�n����f��';moe/e�ݳ�*�~�.��c�Ĝ�uq#odf�7v�۰]�j����6�p����N׮>���_]���N��~��n���)� .vR�����]5v{���uƱ�~���|+9|@��.�����jK{îC�)�=�k{<��3v��/ܾ��߹���}�~�Ig���S"�sƇYly�����pz�X���a��v�W+�tO�~���_ ]��]��z=�ݚ�����q��&�����ǝ�E�򻻠.��ud��G}T�$�ȷ�ir�}�onZ�=�J~̜m�i2j�p�L��g?9�2�.�]�
����F���e$[��*G�&%���q3��.����eϖ�n[��&̽�,D��5隢cpOg���2���x(Y�'%';+�\}@�e���{.g��Sp!ڻ������܌����H�1�>�r��7v!���%��ox��UNZ3N6'ª��B�.�ݫ��ȝ#f>�k���l+z���8}���wh]Ԉݚ���(<$L�$)�lR�����!�Ls�#'H�ػA�pJ]6�[I)�X�]�v�
�3��g���X�����e[�u��'�.�]��]���l=�P6�ޡ�����٤����_��o��fWtE⡛�4����j>�wj� ����X�{�l����e�l�r�h���O���^o֜T��n�0��wu���]��w>���yO�=
`g��aUR��ѯ�6B�7sU�_�͏x�z;;����f��s�4v����p[���oc���ࣇ�������g���iy�|��}����k̴�i����tz,�U57h��//��tC�k�Ֆ�����u�,6\�Ly�;a��<�%b[�X	-�Lə���p������F�t�LD"�&R������} �� ��\������V��t}4��{�����q���&�i��P���ˡ����[���}YK=�>��f ~����\��=0c�-��qϭ���y���ek����b}s0�C�����~@M��}wj�<ƃ��"+bo廮���K��w�-�8�v{�޸���j�mv�[��[�wjn�ˑGr��gw~�
cf���Y�)���f>~���>�������>3�����S>{�&M�4�B������GI��I=[a?w{��yt/�Os'�������wcj�1~[��AIYk���7
u�|�Ox�*�t���q]ƺ$�c����<���IźQ{E�;pcY� ����,nK*����vm�#�:�F��]tl뗰=�&5��m�8s��n��r��6�^���sM/c�.d+��N�0�=A�+)��"�6�5=O��}�ۉ`Iv�r����"j���<M�\��;*a�l�{6�+M�jL%��خ�������������%ݛYn�A�BD9�M��^˺��]d����p7.���^ݩ���_-g���7�+���B[�������뾹Fs��{3v���q��peB]{Ǽ�M�������v������b~��P���~w�C;�]"|�xw��y9K=�>l��0�}wz�6��Og�Y����?u�S�wٻ�S�J:L;�|�>���׍���.��vc��� ��wj��ǣ���kZ�p�Ļ�u��z�P�p�ݯ���Oy@X�
�_�	�B��P��lQ��zX�HX �D%JGd`�Hq���_n
y�6��'�)�gW�7Xb|l��_<�/`w]�p=}��p}Fb�;�w{}ҐyJ�{�x�[	��>�{��3�nvۍx��y)���ES��i���~�ƚ鞉���)hkЦFo,�7k�fc�ý��C����������8 �V^M෨y����ھ��n����]��Rgd���e5���q�qwj� ]����
rCȖ1sk���Ѻw�VS�z'��15�T�ԕG��m�� ]ڻ�.���}��I�Z��);ǋnR�1{����z��z�]���c:�cb;"�U2,&`0`���2�Ξ�R3ָn�";Q򘺎�i�v��.����G�� .���%�7��^�\z���9�WT�s<�Ր;����������Kc��*��^��������:��}��S >�.���|b������wwWz�g.���_�3�/p�M����g��+��,5g�d@�<z���'�Fu�pw)9;�v����7��Z�pt�pF�[o�<��/�l�g��x1�|�
��7׻�ӽB���xm�?\"Aӽ�=�ݣH �#��"�iy jL9�j�d��m��,8�t̝��*Ϻo{�������?�HG�BދmY_�^*�Q�h��ȳ������=�DQ�N�� �B���&}0"����_����>��d�u�W�D2�6KՑ�����=�6}����c�Y�n��x�୓��}���V��z�F7�h�m`����y>}���sw<��s�n$5�������M���/�OK�����ָ�b׷|k��;.�h>�s�4���h�xN��%�CBcٕ^�[�k߶.�eW�ˊ�*�k��Wm����\8Ix<-^ܧ��)�t�x:����{��J�[�u�� ��Eϳ��7'�({���9��;��-�i�:[J�n�1�rrQ�-w�ew6'�zǣ�o{`��7��8��Uv!Nx]O�Nt֏l$ǜ�����7ކ�{^k����M����/y�ݷ>ƾ3gyӽ�p�>}�o����>,x����$�������L���zs�������G�t��F���R-�3h��S�y%�j����5t�x'��Sڄ���_y|}�����pY��Yb��z����s9��o6{;^���I�I�����9�w�C/{#��Y�<`�a���Na�<�9��k'�>w:��T#������|�~>?d�0(ք<J�뇜�Of���=��H�4���ЫZ� I�nY�޴cm�����y=O'���VtR�(���'�w�-�w�k�5����
[��!.T^�'$�ʈ�R6���L�]
$��	(�j�E��
�.A���l��X�UAg
R��R��I��쫁U:��wA�A4Ù!9�$��qX�^@�����fd���S�E�HQs��~�UGs���N ��&��&�Q�Ɇ0�S��Kuqu3�&m*�O2z�]�wGjW��T����wL�C�"E�;����B�<9� Rؒe��H �I���P���g"x����	oY	m��(K�h%^D�A��J�Ԥ	��:��6\��1 �Yu��ނ1LP�2���:�6���R��Mx���8:$�ǠC4�(Bmc��y癏�Y�;����+�Kh�<��C�=�4�>���Wq����,���a�շ�.�VT%Ѵ�^��_G|/�Ș���d��N�0���v�&�=M�7e�/{ynVz���^�0���p.��PJx�}�F#@n��D�'/�5η�,�Jt$ƛD�{-��V������DIJDP��@�'�����w��5e�S�w2�N��T)�Ihk~��W�E��л���ؖ~��"��T}��=	tm8�מ�W�����nU��nfqv �����@]�����a�sݾ9ي��$zǽ��+���mh
c���.��w ]��y^O�����G<�q����.T���]:}u�"�2�h�o��F�)I�mK;64lL��W���0\����-�]K�|��e���Q�n� ���g�d�L]��"����V+�ꥨ����h]��pݯ����c����ide�����k�B�����G�����UwS�C�_��<�4�!��k��m�Yl���%���&�`�X��&%D�3*aL��{Wq��v���7w�=��݋�mk3Q0�njlXF�_�ر����_����&���R�Ş�D��ueҞ�w=��C﮳�wx�
��R������ݰݡw|:}ޅL�#��Q�0��j�QyYx(U��*��@]����Dt�]Mo��2;�����f���Ywb�[Z�����%QY������_�i�M���ӟ�:Ø|s񷯱_�g���\�>X��� ����ɾ�S��}����%/Ip�7;g��t�y���jq�%����M�^�Ic~������I;��v.夼�|1Ȣ�?>�D���g����D
�ݸ�9�r�wd���2�-غ��kp=۲����>�v�ܶ�.���c;��9�8���f���r�uWh������`<�a[���u�7�C��pth�C8�-��[$&u����ǫ�ĵE%��Z�q�� ˌ�%]3�fkpM7����ʛ=�-_���f�N����,�n��QϨ�s9DI������^%���W|������
%�N��d��G<m�v��W��3!�6�,Gdv��~F�~ۺ����-��m�7\�lv��%?>���Zrۯ�ز����g�ʻ��7�=�۵���ǲ]�9L��[�G+��*l��gPn>r.��P��^�������z��
�2+2yh|����wj�/�-u*�z����Ȼ��w�(ݣ���7V{��F|u���lo��q�ݡwfg�W��N��wwV)˻�t�L���w�p�eh���"���7=��>�Ri��ݡ6�7aY�ы
�D�ZXA��&k�"�e(2�ce���_]���ۯ]�<�����U]�>QS;���Ӗ��Zr���I�C�m�'w5j�ָ����mu��轛��#&� �-jZ|�'�*\X}��\�y��7YmX�˻Q �|���2%���w��;�lo��Q�Eț�=�O�7]�D�t�V�����Z��qw]��&���Ƹ_e���˻��o�)�����w ]����� �_xP�;=���=󃜾n�>ͭ�D{��fO-��]���67�w��j�v��}wh]��:��$��|P��$��\����>�������t�*�7A}��k�$����P\޻ �y�s.�-@�-��(����sy�g:�2a.�ߧ)}�w?]��zo���
ʺ^��~01��޽�w����Y�>�S15��|�W���=y�[>��#��]:}��qv�3��k��׵��]܉���������NO|��u��xu�7���N+牆k�^�v���D�F��*3�lllP:��D٬�뉦V��3�	V�05j8{��ݳ�Do6��{.��G����mY�i�`:��=*m_�Y����ݧ��{�;�)�1�ֿ-9�)
w'3�b��s?u6�����ҙ%c�KFrA�c�{'ѷ1��]9 ��^R����]��~���f��A���<��],suK�u�Ez�뱌�\�Z����&`DJ30�!�k�w ��X�ji=�(������o����9���=�C�pݫɊ��>9�b��t����ܱ{/²�)-~w����t�;�ّ�Bǯ���|�wwjwfE.�`L�q����'ї1���g���=qwwu��|�s�[5���plg�MUK��r���w�Q��\b�~�(Y�F���/�y����/<�$dTU�Cm�s@�9��a9���$G�2	����Wj5�����n�o��o��HD�x.=q�P����]� ]��wP��	�cٞ�z-����;��yd{/²�+D���Wq����nGkU�{�a� K�maS���`�[�^m䇫��ݬ��N4e	����%)s������m�g��t/W<�NY��FOu7ϼ>݀���j�<��\;���}�9��T�s�ZF��pP>n.�b�g�~��V*�����𻋸���ou+������B�o�d�e߅9���f>w��.���z�=��ʹ�Lo���8��+Ǖ��>S�{��_G����_l�J`]껀.�]ڻ���tH�.��s4�ۺ<��Y��j�v��9k!k�Im���uE�W�ё��;�kϵP|ya�	O���,y��_6�ݶ=���^�Z0�ʇ���Ͻ�3F��8 �Z��li�qaG��� ��C�qpۇ4c6uM0�y�2Tt��k��ù/�T7Æ�T��%Я;ev�0��k�n�S`=p��p���ݳ؇���\�Ԝ��is�CP]����w[4t�\�!=�NW�ë������F��=#�=�׍@v��Wjv�\c�����v�m;ݫ]@⮔���KU�ӑ��7]6�}}Ϯ��:��U�rV9�e ����v��T��̹���j�aD�&b&L��+;��|��������v{]�S����G�82b�<�#�m_e���&����-����������~��MV���{�����fd�M���V��DG/\��]ڻ����w�{�u�M�2��l�c�6Q����b��2־�N����F�ɍ�;#n>�v�����+{]Ч7K@S0�YI��*��kݜ���6�����߇�"{�����O�댶du�/k���� ]������Kc����S��2p�a$ș�$�x c�ќ�Qѫ�YvpJ�.�c&I��s����<}|�g����}���=�*Q�Y�����r�=�=�ܮ��.���·ʺ,I���ț�t�B��>��߼�o.�w4��}�M��X�]�Z4�����b�_�<>t�~#�	�Y��j
������|�f���ⷰ��
st��0�B�����S3�5Q�:�	�}��7qwh]�d��I�T�Zf��vMb�~^�����Yi�O��_�ߛ�l�?6�c���1�޻��^��h�F]��50�d��v����w��[�w��}���y�j����W�����]Ч7KB�}Bn� �-�"=���q��XEPF,	�:m�q�դ�n ܨs\:�76���"�	#*&-v�{���Z��kW[��>�`q��<j�'On\��N��������;\y�ugG�!�DkٯV{�T�.�w�Q� ]�W�:�z�9|.���[f��������&nӥQ���%n?^����J�p-�b��\ӏG�g=�}k��'핸> �$U׾�LǴ�"��&�j��t)˥�L;�.�.�ݠ�=�1�I��˨܅��Z�+W��=���}yi��ZݰxO.�����iϭ?[U����=��;eS�g�}5��n��e����n�����w��?OP�К��5ͣ,����7t�j�%	��F����%# �2$�Ob��,��.�����=�c�
r�h��Ǔ���mS�6��wwt>���iq�Ot�@[�v��	��u�����|�?��r]�N��[��jᶾ��w��}��R	�X(�+��}�ֆ���f�{q[Vm9��x���F�`s��wk�`�΃��c�������){W��;��BBI~{O��䷞�{2�*�x92�p��h�2�1u���cW�^ʶ�1S�2/!{G�r�mexj�	�J�1�Q+��^��@����}w]����I�Aq��9�1U��w�}���.���>��.�$w�����}��!,��#�,}L�6�^ɶ5�$��mם�u!fe�=k� ��u5n����߿߬�����z�k=w�#N�p���Á�-���_]Ʋ	-|�ZpkKe����B���O:y�z��:�N_O}Uc�w_�'���3:�s9��Ne�e�j��U�ؓ�1U���8��_]���.�]��ݾ��񋻒��S�oW�����v�6j��)F���5���4I��@z��ݮ7�ث�m�)���op����77K~����~���~�c�����O�*+_�TD�����TD����YA�7 jVVAVVAVVQVVU"
Q��(�[�� XF��"� ��py����,�,$ (�����HD!�7E��"�����"��"��"��"��"��"��"�V\!�
AAAQ�
QTADSDTh"� �"� ��"�v��� � �(�(���
�T��
��*��*�9�a���T� � ��F?�mr��s��ϓ����?��l����s����0�R��
���3���ٿ���~3�?(�*+��?3����ߘ�?2�*+�@~7��-�8|��C�'�?��}���	��������-�0,g��~��)�� (��VAV@dAVTV1X0AX�E� E�DXE��Ab�DX$TE�EA`�P�A_� "�����P}�������DAY R@�Dg�>)���Y���}!����"�*+�߾�
��ǂ��t�G�?�l6t>ނ
�����_�g��Ø

��
���~d�?-��
��_�=�����~�S�t��)�c��G�͟�(6j><t< ���C�c������AQ]82�w����>?�������~���AQ_���>�TV��t��1�� �g�2������CX=�G�����TW���$#���G����Gǃ�������X���m�| ���?w�������(+$�k(z^b "+0
 ��d��C#�                       �             >� ㄄�P�D�� (HT���� %TU*�J $
��"���B*�P*�J���($U�*�^�E"�B�TIB�B ��(%AA �@��%!B����PEP*�UR(�TAT�"�����)J�A*�$B� 47�_*�x��<ڗj��ۑ�	�ӭ)WxJ�;�ͫW��iw��^6V�{ԡ�6�t՚��p=)ͨ*�ӽ�^�J"�
�  � ��t 6�TP��
� =8�� � u`;�r P^�=��z5M{Ԥ��֚�޸�Wv�W��y4�Jm��z��h

� � �|IE(@P*���*AJ���օ��z�Nmv(�<�N�Ŷ{�=R���UO�[���m��m:S�J��ׇz��w�����T��[��Um���@��*C|   Ү��Tz���Ug�!Η����Ū�x��ҷ��95{ۅ�s�J��T�������o7u��z�^��{�=JB�T��   �T$)R �(RJ�
���4����,R�]
�uynZ�U]��h�z�{�E[�xK�N�� �w :@�8U����{�*�=�  `���������g@� �7`��& [ n����ʒ� ( {�  }E
��"�@��| �� �@ � r�*�	���9v����TU�9 �R�UJ   0{���©G v�: �����w` R�p r@ 2  �� U
/�� }�JD���*�R�TK� �� 8����9 �R� � �� f��  ӝPI���>@}��RJQ"���  F�}� |��4
�����#�݀r #� j�p M��{�� �7X ����IT�2F��S�1%%J=@�'��J��Q@��0 �d���@ h J~�%Jh��`�LMD�B��x������������XI"Hc��y��F�?F]N&ސ �p՟_��I>�$	!!�$$��@�BI��II'�I!������U����������X�'ۢt"s�̼3� ��#�وKܷf&j�^E�v����^��:.��mE����p!ڲ��;3�c� �ӟ�t�Y%���K�6dK�pc#�;��\Y�iY=��cdI��e�&TOp7{?B9�޶�*6��A�)�Jf���s����Nq7H��*g^�ZmރM��^�o.�vvk	H����J��C-�F�u�4�tn�t25�5W�8g�<
�ҳ��w�oe�^5�.�o���J�S���\�u��=��(�'��mٸ�h�s�B���{qh�a/E�.=��B�@�� /w+�Z`����c%��-(�=l��x����)C2�ƣƧ1�d��Hs�,0�XPo@YV����3�U���U/y���az+ׯl�
�.��W]�ts�ذ�vΜ���>`��D�i���#E�y��!�� ,=$��b4��8DO���(���12�cn*��Uy��_o8+1�ڶ��q�6���f�Κ��΂8����>���u�7I�\�:W>��7 �`P��.���2��xj�Q�r���0�Rwx��K�1��2.�򜜍�x�TV��ys)�>bɰ��}>�8������P����]8WK|��yq�"�����Y�W2�4&��0 �l��N��)1�wi�{�}�;��Y$��
"^�7�M}N�}��"ch�w��\&ui�����b=��+�T�����n��C�Y)�s�HS�E��w�sgvNނ�H]h=#�Qb����t;��M�e�������H�s~'6����j��hM�Q���jLM(\�����>pl�U��+�˖��<��o�
�]���'��ac�Ɓ�����gV�M�μmz~�(�/#tAnw"TjZ������.K*���j�bG����o�gP�9H�2�#q=)��4��³�BF@�V���n�/��d��\7�X�姰t�}�����Ќe�'uex�4W�{�6a��\�	�.ʪ�u�3RLp��Z�QJj�W3��6��B[2��wF�s�{��Y}0S6m�ñ�Y�EK��dP�BSS����dl��2�A�p��\�R[��Ԡ�i%r�NR�צC�L�ms	3���F����t� ���]٥rNm/��=��禜��;�<�	
�#U	��7,ۜ��G�m墊
��^<!�bZ󴞜S��Jy@�i��LT�;�񝆱��	���v�d`�B�h����:��Qf�H��5;�7�_nh�pmp�6�4�ܞ=�4�ʳf;����-���
�E�s�C�ˡ{ᒙ���-�Vjxn���A#�2�vMn��U���z�G�gE͆�(���Ċ�)ۧgv��o(֜P��ʝ%#��A��gBã�[T�����#�������-�}w]���]����
�.=���*ya|��N����8d�4���@�η��={,IoRn���ѥՉ��٣&������p��8�X@���*V�,%�����������\��`D����@Zj�T�����ݜ0نi�Gp���L&����3��ܜq����(!��:9�M�%+U�qL9n��i�۹.��b�.'�Up��z�"���x��(���l�W�W��&ph��|��u��wn�)���6���#Z ���x�����>��9��v���e�.�"K��n�{��d����ݗ)�s�]��n��A�q�>��)��7;�l�qL]Z����ص�.����0��5��)���mZs��ec����^��f�a���V����H��!㔌�5�S��("<W_/��4wm�]DC\��b�Bb��=��E�;�Z֨�w7vW�.\�p�+�7�bnm�:�w�^�0��6&:�ǘ��+޻�7-;���(�v���E�z�Ź:�f�XwOp�9�L,$6�$ls�u�|l*x��K�:�G+�%.8�-M������,K�ʳ^�&_$8_Mr��J,�D��ru�F!@[ˋ�(�+-ѩ��,b�W��'qU�M�swUSͥ��H�\65v�ܳo7vӬmե\n�EbO�$=w��
�H$�-C:�xH(�H�D��bOA�9�4eb;�p#U��]�>̕��Sw;p"t8�9�T�jg���6n�hY��Y(q��xd�ŗC���� kZr�4C\9�R�8���C;t� ���՗�?0y$����w� u���)ۊ�t'�p�-ﷲ>e��8��=�<V�Uy�*�壡L �w}{ݓ1{G��G��t�GL`ŨųOQ�Df�6|�u��!��Ga�,��	�Z��%��mz��7����1eQ \�2զNr�s�[gi͇
��Ũ�I�-�]�
Or��OY�sm���@��In�E����g������x-���7��;N۹l���q��kša⺾!sl W@�J;�i�iF�jg�O�nk�̭��:�h�1gpx5l��R	-�M�!�'d�|�c�Ά\��ͩH�n�*���;{7v�PYkbz�Xg'g�S��f�sa�+OU��	5�B'�lgIa��U�xὗ}y��.l�i�=�5tqE@���@�H��}G
~�
�޴v�Ι8 ���f�CT�����=˲�%����L�y�Y������ �S�ԗ�w@@'�_<lM�����n��_W��a����.��Y��ܗ׈��'K��:�i�9�i�ߥF�,�K옆��@ɝ{xL[���y\A�0�͏���8F;{�n98{����f��<ZѴ2�.(iw6������ۑ͹��ʓ��jHn�7^%�9h��b{=\����N/%[���(U~37�M`�����L<��7��WnsU -���"F9^��
�6]%�n��{�3�vrm�gq���rl������T��j��Mۯ4�Y���sw4�4�ne� e��;	���Yq��� �F�פ�����H��[���v=ݸy����%*y��y�]vYۭ��Ǔ�)�7dN[;��������7���dѺ��SC�usǷ��M�YɌ��a���ٯ��R��̢��(�~��	�pל�f��fI�{�˴��䅼�u��Ҿ-�b� \t�(2�vS�ݗ�;�zv#L�M�,a.��M�$ʳzD�*+ͧ�����gF-� �IvM��ht�cM�r�^O9h�'s�3[�gÂ!�遍��,�<n�7咍Z0��ݚ��{%J���3���.��S��s
�(�c��cCHѷ�R�3�8r=�olGo.7f��T�:BT��ڟ(����J|wV�7�G:鰲�f��`�_M3�* �˻�݈�s��Hu٫�#�V��vۏw9�rL9��R�ӻ�fٹ˸��ц�kq	�{6�����x׽n�t�B����^k�>yUjIq�YIo�扡�Ms�����:��2�"��JK��P�	�w!�� p[g=�ޗ^�C�*猥0���8�4ܼ;*�shʀA��^��N�KX\rۢ����-�;h�n=S�:�ug"i��S�t��Vt}+��E$��9Cs���Z��R�J��yO�*gbX��n�E�~D��X���=���%��m�h�&��Z�:- 5��5a�R�c����'��c�M���Om�'���w_L���-҆����"�w����4��u����N���=n��:���MG,������C�wvE�,又��d8y�����[ݚR-�w��r"�	�Z�d��1�s��^���|�q�/4qy*�P�2�t�sF��k�/r��s��=���Ru��Yyvk�ߋ�D�6�Ü-ٛ+ׁ�OڎV[��Hժ-�� nn,��^�7�
oe��֐k���ҋ�b�=��,|Ry��Vӳrmŝ��C>���AR8�3����#�N9�Vi�4b|�ܞ���U�����ә�k�Hi-����ޥ)����ӏj&�ɗ��pAm��s�Q�ًQV]݂Bx�W��պ���Ȧ�j�tc��Oanr®í����wM�;sC���<X�EkC�!�!�n���k��sLi�/v���ss�� �9��]���7��s�R΄�h'tG����R�r����rs������D� �*�B�B�;�yr)8�b�ڸp���&�jT)��ٕ�����b"'�q�,=��j�%l{Zn<��mt�M\ɑi��3�Ru4F�y��f%f\<�/X�vb"�oa&�cp§ ��N�+T�3� 騮�#���N-b������ɴ�ay�Z/������:-�X>���qDN6n�rf�p��Ε��[,��`���l]om��y��-�Nܡ,���I�ے���$����Q���GZ{r;m�ŃsV.�f�&�3T�1�Ev&��̪�x�s�Y�Gc�~��z��|�v�܎1��vk�M��;���gZ�k4<݁V9�=oh��e��ph�d�\��:f�V���1.�mS�Zx�)�O�&�\[P������ہ<�;�i΀�懊C�s�]��ַ��S�rN�\�>	g�2�yׂ[#�vh�g��٠n�:�Un��2�����j\� ���n����ɳ�LQe�hc;.^�h��O��_��ۼ�lh[�w{c��ҲAV����E�:g7[�_��#��t�d���%�_A�����yi��WF��7^��E�R��h4轗�.eͻ�C庄�K}��s~��&���))`�����\�]B(Ov^��Jd�G�hz��<(r� q�i咆 ɮ�uPfʒԴ �a�:Q*�Q�d[��*�bi���|i#A|:�z+f��%��run"EѼ�q�^�;4�9�z�܏�LGiŷ.-�^Lc{X�+e�h�������݅^�:�ͯ�v<=��ZB$q0c���w�(A(oV�-pδh��X)ΔK�999u�As]�#M�N��Z͙N�8�&�m�0ᄳ�׺٣�0%V��㪦��_CM��%'o\��LH�o�f��s h�����%M�ۭ�'sޗE���v��F��1ݜ�n%�s�䥧��.ܚ�@\�~C�%���ъw�'DF �u��Nv����_C	`j#vj��~�1yaii�ϓ5�٬wn��i:�����;��q�#� �)�a(h:�E�T]���ɥA��u�O�&W���'R0k='Oq��n�3�m�Vmuqg��9ݝdf�O,Pb�v>���)Y�wW���:��I��r�U0�ӆq8��7��\���&t�_&nP��N߻�$� ^��k��7QQ9�h(gu���{[��B
K�]��:���i�R��īZ�T���1�u��=����F�3��B����9v�g]i�:���iE�S޹���Z�h��ŒA5\ܢ��c���,�D:��;>��؟:@�n�%��bio-�8���T�=����1]z�a�e^jM���P��e�#�����&��j��B���Pm[�����j�j�C��B*�{���N��{\�P#k�T�`�V>ws��Ϝ]��n@IZ�J��ٱ�y��vd.-�h�;���TV�z߆�x�|����Оk.��\@s�n.fm��i����G,f#D�w9�6����8!A� Xһ@���p�o9�in0CY/�ޚ�ij�{��>��#:|��oT�����/���'u^4�9��'�Ku^Zr�X/l����;s^�����;p�2�a}7vU��&�hc����PS��V�0���]]сݼ��!ݜ0�ŝ�^3�0^��h���5on�=�m�n�uN5�����+��ŝ��*R��3�G˝T��3�����x j��
�Ng����{�$�0M�9,�-9	E��gM���{��J��unr+r��������4]Z�-�SP��S	���K8i��ہ}����� ڀ��@*{L�vwG\��&�p�f�A۵�We����c^.�Ր�q���CjVn6���\�tH:�.6]ܻ�F���6
�����q����6km������{�g4��Q��m��nh�VAp1{������kf'�-{�oܙq�����!���t���q�H��9��
f����6���ޕK�y���O��u��f�7 o�p��jkl�����:�u�:vDh�7��3ES��N<�w^B���Fa��O�~V�#p�b�%>ǨkM�0�]D�
�g]���77�:Lt�1�䫔F�{m�+J^Ӻ^��tk�a�u�B�
+\�U�u���aJN;`b�@Q�]�٦�x��we��Od�v�C\��{��&�&�3K���a�&�HDےS�8<B�gr���S�s��:wQg/C��������yv���h��BL�l�ti�M��Gxf����k^� �/>�_UE��U�q����Gx�Ki�0�ݼ��;I�yk}vӢ�Sg�v�ow8��>��a��wl�m��Rv�q��lG���up?>�婫R�����僰l�c�w�����)�T0�����I<��ˑ�gA^�a�K^��j@&ں�M�͆��������O$ ���
I	$�$"�U	d�E 
 AB@�@P$��H� �	 �$PYE$�A@��(H�+���������������H) �E�$���XH
H$�"���X�H �B(!(d	$P��H��E,� �AI$Y , ��A@��I��� �Aa$�!E$��$���E��@BEII$"�!H$P (H��d d�E�I"�A@� I R��H�,� ��$���@R Y�I"��, $ $YH���?�	 I	� ���w�u\������黪��hJ$��Q��7��<�[S�	���Fl�lV,�,K�y/vt]�-#^Q��3DTe�r�V��1��A���3f��>�sj^����tMD;��[«�]{����:es���8^{��V�޼c�"�M��1={��:��Я����xw�>�]9q��CMy�<:GW�出�l���\L+�F�6m%���ә���W1;��ٲA̛ݑ��Ù�<x?C=9��i�=�)\Th��n�`x��^�E"�����ﵲ��ƺ_sO��h�r�����'b����%G���:���4��0�J������d����!�T����57d��wHvv�8{��,�n������8&�<�������z�-����E���ͣ��	n踯o��87���8�x̓����F����̚M�F�*LC��������P{�9���rT�k@[�H�N�xж��(�ܻc�Y'���{z�ޚ�1w����ו�n��~$��k�5M�1#dn۶��^�7����m��-����fz�ޖ�A'�j}�n�����ٝڪy9��G�v����b�R$]�&w�6����xr�o�)طp�D��.X�1'`��{�<z{���[�J/�L�ȯ�������=���vIٮTOLʑ67��>�_y�����^���4�)���c+D�q�.2�V��aρ~=��}�`�Dܾ�>ӫ�F�:��G�p>���Xw�An��d,Gf[م �/2ٻ�u;Aa�֮�1��.�	��r.9W���\���,���?`����l������r6��;ad�A�؊M3LiI��Z�3�^��6d[�i�/��.�r\/&8�)�zf"�8<�Ӄ�����t����,y�����K�>/L���R1�'"��ۉ̘;	e�ƶ��b��S�Ҡ���a]|��W���j����� �|13��F���s:�{sT��i������g�K�Gw��	"��/�"k5c6���{z���WAG�kWЌkW���v<hk��	Z������3���R|������y��.�n�y�+S{�w̧���B�8�]�b>�ٻ�"�����ɾ���B9�g����F�Y�mi��*M-���7�uy��v�Ց�m�ıP-��	#V�r�J�9r����n�D�λ٩�ĳ���������x�mP���ʖռ0BNn���2_=	dO��{��^�yFh�13���b�m�DT�-nbٚ���v	�˛K72D�F�e�I�.�Fa!�\������9�V���Q߹8�{_��Բ���� ������G���9;���s���Z���5o�C���tӢ5�͇H	�E��s��N�6����$�z���Nq�w��RNy��;}�4[�Bi�`�0����kY�^F����v�`R�n�Pgc��SP��03v/����\[v����y.�ɕ���|;��"��~=g�_�;�'��� [�b�U�`<!�Jnz����L�� ��{ݽ�z/R�k���ty�G�znl�8�}�GyOw�ɽ�y�M~\��V���N��� �ֳ���5��� {Ħ��ݓϥYܥ\�Gğzf����8����c��"������ȗ�=��^ƻ�/��n�L�4{�f��v��X蟣�n����x�Hrś�vEZ�ʶ�ջH$� �g(���f�ݏt���r��i<�`}͞)�d�6��Z]��M�(9�ۤe�2�סNS�&]kp��=�gO9�A�����傑t�{���	/�E�iD������116crt^����6܍���u��q�4�S1\����~�7��=�4��-+<��B��8{q��s�Φ��Ny��� �g�}S|�j��1����gt�/����>~>��-�GOZ<�g۫Us-祐�ڒ	�5-�]Vi؍������>������b���{z2�	�f�͍��کe�XD�1���;�7��[d3 �Cgv�nչ��w�w[���^:d�`�R�ܹ�k�A�ӛB޹�˜˙�V��@�t�L�ܢ6R��u�s~N�Fm��S����e)Z-��҈�ȌS��<�FEeFs%>�ޭ.z��{�w��{z^�:�64<��8L�-�(�����ŷh����F���ݣy�I��F�¦�}24\�f1̚�7w�ܹ�'\�Q�3�Kԋ�n/r��{T�����"����V��<ӛ��0D���gM��v'�5�	fz{�Y��������KݍL��-�H�A�-֝�)� d {��jwP2�ɼL�.���d"B-����V�:mȸc/�>��V�U��^Λݷ�6S�go����#���������f��L0�����}�s�@��=M�9�=��q¯i��F=2n���
��ǽ4�֕�^i�c/����R�%��מ�ixr;�Hsה��8cI�#����Fy�!��.��N�n���>�&S�\]^o�4��L-�M�}�M1���d�o�>��zp��v��W�[����Kp�}{�_h�n�ܻ-s�M�����{��{ō~�Ǥ���z�NG%������x�&,�yA�(�7.��P���\�W��� �3@��['�;���X
:\Q�N��bNn���TEe�;��mʅ�9�MX����a:����SI�w�C�j.M�s�Jql^h�4w�����a������P0�&vB�e	�=�c�I]�{��+�r_*ѐl���w�^#�ԻY�aa�y#fi��T��.��lE�hf���ʹ�o�_jLx�W�^��_w9#n7|��̟�\9�}U���tozsͲ���xp�y�}x7	�;��^�8��O��<�{��ݸ׽b���X9���`g��4;�����VYm�y_�}<|�nl�w��Ck�L|�������zxj\gd:��]�����q���փ[4''
;�4T*��f�:=����r�z�h��Xk�؝�VtA����;aQ{R�`���C�f��s�ECw�^W�J-�}��P7Y�C�N�M�&��X�ys#�؊����g���V���Q��i����I�Ȑnj�ڒ�Ӝ}����6Gմz:��p1c�21CF��[*�ɦ�vE�&f �]��}�{{A�6o�{�o���{��EӇfZ�Ң㪯8N�����W�$�BF��Lƃ���a�n��!�!�w%���E��YQ��v�gӳ�{F"��I���HA�kgd�̆b2��Vr]�^8��4��Ӯ
��G���KN4q��y�Z
�����>U5�1^�f�2���v�ٹ	�A+<���uw�;uPyoH�.�O�ǹ�eS1�ŘA��1v(a,hx��n�ޢ����X��<�۵�O�����`z�T��d���9�{���6����F�7p�`'���h�cL�ѷ���h==����v��k�v��c�#x3��٨��4f�D���/��u�����-�k�{��k|2L��#t�����S&"ꖸ��^w<Yv��YO׫���QuI}~Y�J{��q[os<�_a��zl��䰦�ÑC���|�V��c)x��q_���u+7�Ov�>��~3�n�ky4(��=�ֆk�3��>���;7E�Vv	f��lO�8���avN�$�n���������:F�zor7�nj�3:s�!���_�)șCf6��:0)q�vۘ��s�Ҧj�a�#r�;+���T�Fy��3|3^�� X���Ǿ�KFZő�d.������w��i��]���޵�����o��&�Y2��{��̍��-�NKڮ���6��ܼ@���=诰�sJ�WFv�y�%�����kW/l��}�7�1�Afmn��[rc�ڌf�*'d�~>�$�m	Y�o0����� �Sl��X��/�ڃ�b�}縸=;�{��Q��M�N��@�>�@���㐄�tJb��M�IGJ}:����>��j;uf�ӣ��$�N�y{���U(�S��/��ۖ�Qƚ>"k�ޱ�����Ͷ����H����:@Y<%�7����9`7N7X|`��
/����Oq�޽aN�y����z6���/��nA��s��U{�Q���ܳw�`��y�뵮DlE�K]�������Z-��puU�P7``�u��P�Y��.�����ɘ:oZ��N]Ы�^�?N��۾9��=w5K�ޑ��T��8��XdY�R�*�Pƭ�g��<~�Ⱦ�wϴ��.�����T�t�D���tJȼ��`��>ۖ�����F�_M.Ǝ��vv&�r�.�7�}q��D��L�<G���']��2nL�e���ݽ��n9��`هu{�H�:��}4ɫ�+;�����4�Q�.�q�����<uFCݹ�[�sX�x)���q�$x3��UЭ��f��bc4!s�(\5dLT�ћp�������{��T���7�>�j����g (!Q9u;Z���su�MC�������X9;U�y�;-��T,�ݝ����	)@����.�ƈ`�� �`Ͱe�@�{��l�׵���+/��Ǿ��]�5k .d�w�|X[Ι6���IF�a�{9�����.f�u�ǻ�!�S�l�ꭌj��:�N�17R7\�#)I���m
IV��jN�9�]�>I���X׳F�i�謠����z�w��d8��:0䞶�Y�n�lӴ��<�)�zQ_c� ڰ���;h���w��L�5&��j�vg�NLؽ�T�ȭ��%�TYxp��-���7{��Ѵ�!n��aM9�̲�w�pS�.֩V�B/Th�3o`�䊞�$�j�e��g�t�0ԋ��C6��ۢp��j�4q�_a��Y��C�`���c\]hsB\�Zq�/Z��uJ+h��(�����9;V�,��y�!���k޵���G�)��P�Ag��Oy-�R�j�5�~�����'7��m.`����~�Y���*�R8���1:;��9����E�ypn���oa���$^�ý&`b7�ل�P��̫+bڈ��^z#"lų(0�4|`�Ǟ߅��yܾ��e��WZ`7}���o|�|��_��z��2���w�)��Y��q+�]��G\Q�y������[����Ū ���C�F{�Q�̚�փ���N�6�g��6�v����\@d��]8��2��#�����u�׺L	�&cD!��I��{ wgo.����!�[vvD�Rb�kFe̍o3" ��^��xH!�&�N�/@�+�peo5O?�0z��<�w �拦Q�7�U��+J^�9@���иr�!ܷ;&DN��:6�[�)��IT�&"sQ�N�)�#[�d\T�͹�1u[��M�Fo��Ӆ�=�e:A��-��Ovv��%T�$iW�& F+k�73X�z�6�O��y�}�����6NI�ۋuP��p�B	j������rN�
���S0M�u�9Snv�e��5r˾s.� H<���#ݚ�C����m�r��2���{�>��	��\�t��
��mК�z��^�
�[3�4X�q;���t���)�&��ТB���*�5_m9��s��7�f��U��n� )Jۍә�����nIZ���%��!^�r��z����Q����OK2|i1B�ElD�=�-�C.�T�ٸI�,]�9</�����.���H�z)�uyb�8�:�R��썭f�w��W9�����F����d?`�Gsg��m\��mM<�B�6�w6jy�íVD���q�;�-l�)%�l�n\ڲ�i:�ͷo�7��� �k�_zxg��i���y�Y���cPy�Q�!v'sJ�f�\72F7;5�A�0.�ӡ�dܫݹL<� 9;��<��=4��O1�}�U��u��ջ�1�����T=�^�����_L=l{��z�u�t��\�v
�g��fSIW��w��]Io�k�M>Po���y�MŜ�MIi�	����osk۩�ڭ�jbJZ����.2�V�Fx`�5�T��^�:��'�W,VC�b�ʕ��6f׳�wOS��G��
껻�R�P�V�w����N�6d�M���,�P�x�;��f���b5���KBԺ�4\��
�]9��"gq�{�ckC2��ۀ�LN@�[��,ȧQ9����R��ǟ�N]s_;2%�y�k�Wr���G����1w��	b�S7�9�QgsN��!y��7=�wUz�`CQQg(K��oF��ݻ�E��z��93�z���y.����Ks�͂6��;�d��n�:�.B{Q�2�%�{+w��w�����7/]1LFCk�w�i�����E}�9��!E�}ug���������Z�9��.����`�M��d�:sJ7e���#3�W<"��v8û�.����;�Ձ�X"o��D�b8˯�=�07U>=w��2���c��*�o�	��	����pc�|�����s���Gu���p��'x��PA^n��*b�!��2wK�zN��hV_^�s��-gnj���թ��8����Nr�}�[=��~Y�͈��/�f���iUZ/g/vdE����k@��FO�����u+�)=����iiא^JSpj��Ϊ�Wb����Q���;pk(Q��=�mo�H�����ó4Ӌ���Ã<�x�wG�����2c�b4�=���;t3-�j��c=������M���roMYz#��޹p�ď�f�]vH�r�p��Ӕ]m��#��"�oC2���'N������u�!f�=�v���);�{jB�A���z�Q0�e��0�LJ���h��ll��Y��)�v���cN��]\�k����,؅�fc����Q��j��7;�Bk�{�Q7��j�����N�d�U�S��n��＞�^�����| ��M�2fK�;�,;�&��UAf��P��4-���wuwEVC�[����}�< ���� }��hK\5��v�i��[Cڮ7E0�n���/nՇ��ݸ�R�2��h�:y�a-⳷bgrR���tH渎y��z�I�[ �[��m�����/r�qu��y�9�3h��Ӱ�ZRU-tم�s��j%ћ-��L�[Iu\A�$9ƫur�v��&6�]�n9q���������Fβ=^!a8�]��gX���[4�[Y{3�n�Ga�nz�-�w<�%%ֶ�s\���GOX���q���+tc�O8{%[v��,����N��I��c�D*1�,	Z�b�L^�g"��F�4ilV�^���tl��#���ݹ8�kq�.�tz1yvx���z�q=�p���̏F���ӸwJ����o�~��C��1��	����5�-�(x�%vN��b��1��<r�.�X�
�;8�x{\Q���;v�Ű2�L�8t�)Y�K�F��2������ֺ�Zݵ�"��k]5xV;s�r����<f�zG8�sm�6��˴�ipůj�(+C�n+�V���Hx��¯���th�8m:LH���;U�z�-�5�p���qu�N2�S�5��d�B��=�������nJXљ�v!B�4$t�mz�`�ǡ�7��*�Ξ�v�]�ky�i�f5�`۬����ڹ5����cV6]mle]�M8��s�a��֗���7l���*���M��vC�.�Kzw	�T��ە����b��>ɮ�=ZUm�{@tv�1���2�+�[����N{
���
{W��,f�X�Љ�V8h����b�˜<����SU�8�F-`;+��]\D]����a^���Ŋ��[�����7F���8m�h]�<�xݎ��G8�N�vn�;�t��by5mvB먙]7�l�ei�l��M����Ɏ�`:;����S<�\8�벲���!`^j���v��:����:��k�Q�n{�Z@�Ea1*��5�3�3\Z�gB�]d���\�25�,�R��5Wm�1��t��Ûz0&%}�'��m��Ƽ8�z���Ǘ��:�zA4C�`��Z���p�[��I���ZͬsM.�YYe+3�����>Ҳ�׺�ŭmv#�ᗋ�Y8��O@�'0���l�h#3e50 �[,j�.-v��4����mi��/fn���h�X�t��W��z��<����Z�9]�b���X�bK�P����t\��sb�rnN�f��s*T�-�����^��b���ތ��}lV[X�"4٭oa�xʼ�l.v��+��q�0���$0�K�m�X�|����2p;���O}��v���w9�v�y+���i�)�z��)�L���l��|6��%��#��q���gJ��8�%�8�f�4f�,�a	f����3Bi�5��!�2�!CD�]jF���5�Ǒc�y�)��g����!��;Pn��X�>�=b��rx���q�xWq�*�&{]�y��e^�����k�]��{��m;��!=Z��m���E�ecjۛJ�ܡ���d���ɦ��G�����6̰���JQ�V�0J��@JQ�u,!�%�ڋ���d�Y��܋OQk4v�Ks�v��Y89�v�'ly��B�k�u�I�)694 npu9U÷�M���㤀T��6����٧h��n;����wF �����p�vҰrܩМ��+V�t�ū�%d�l/l�W�+n�c^����'�l��f�Թ�(�51;�qz�{u�՝�4�])����l�<�u�c!��-����vgP�z�]c�C�\����9o\�<v�m�x�MIې���
���Xu�m��E�\\���Xݮt)�UC�1Y��6�^ng$�����z�΋i��ܳ���u[b�f�]��I�i���6zL�;�����`�^"�$Y9����.��z��uv��(C�(�i���^h˖q��y�GE֬q���H�+��C	P�í�\�a��̣맓�uk�I����8���u�:ڶ�!�F[k&�l�������s',K��t`�68bh���#��&c��k�cu�&��)��V�v��;�eb������)nQ���h�{`��*����މt��77Gl<�@�d)v����k�=s��<���9��\�Ss����m�;�ޢ�I�`�ͱA�F�"E�P)��8%�ٵ�	�����Y튼�R��D1��LC��:��������ͅBm�ZE�I��\ݒ��f��h$l��c�5$h��3�Nz�dJ�ְ:���s��ݓV�Ub᧒��E�l��`�;f���c�y��ʶ�7m��s���6��6tk{W</j��Y���k�o������{Scv�=�A�-�<�
�3=�uiHn�"Z��j,�2b�:+uˁ�f��,��k��v�f���a;2�z����%�[(�v���)��HǑ;�ʾ�:�]��Ty�$�/����M!\f#�B��9������W�X\f���Q&��:1�q���.G]AѬg��e�|�k�3}Z=,[���/+ČSݽ�4�3�y��`�ꦋa��U����K1؀��pm�]�Ytm�ͦ�s,,��v�s���;�w`��vx0�GCZ�Y�a�+	�R��hR�.��Y�i�j�]�%�Q�ܝe��!�9�a�p����{\V��S��CK��\�����7'n6ɸ=hJkh���ԧ�\@^�XT��h��td�Y��͒Nr�q�y3�9�dN�I����r!k���qΓ��.�vz�ɽ����)����\A]+!�ݣ��n�vN���v�,a�t���A}�X7���`����y�{m�@:�������� )[knTeEz;x�pG)�)�gg�p��9�<1���]v�i^���z����V�C�֯���i��,�h#X2v:��x�v.������O@��I��:�jEpL�ka\Cl���	rjF�Vj"b2�&YI�W���C�n������Nytl�:Ƚ!<�MQ m�q�3�6Rkm�8ͷZZ��EAl&X�H��n-%6V9�Qf��%�N,�m��Wm�n�e������\ӈ�:W Ǭ�vأj.��Y�f$!�Κf��4�h��iS$U�8��3^�b2)������Z�%b�;�Y�irb"�ݜ�u
'[n�j6`:x:M�y]AW1�dz��lW�,�)�h��9�m�$�3�:5�����pmX���ۀ4i����a����rhD�n�Y�����-��H�/<Lx�X깻M�z̒��a]W^.%7��MM�z��Lp��r6��뱸�G:M�0څ�v7l�n�>�݇��m�D�;5�m&9�O`�k��Ǝ��#%��=mۮ4�jdН����G�v�8����u��dd.o0o��֗qW�|����㟗�Ŷrn;i}!���S�7cU=�����X�[q�[V8��M5Ŋ(�M]*�&��D�^0��T�و��pqCn}���G�6"���u�݅�s��m�g�X�b����Qyϲl�d�(�fr:6�۴�f�u.��a��άy���BNF�M�kT�W%c7F�	i��ّw���c�s��jpن:Y.��=��;n�+���kGw4��-��,��5vts�<����Y+׮W���wDh�7fEn��*�{A�Վ{C1�����/%����e�a�#,�f荸���;r��l9��-����M/3'Bc�P}������n{v�ܺW���q���0�t^5v�&��e&�=B���*%��bm�2���8�-=I���ܕ�ح�>�$*�s�m����&�x����ٍ�hr˞�S&��[uE�9E�<�c���3�v���T�.
��$���v��D�0g*z�p���íam�]a��R��B��s�L3�m�z�����&땍� �j�l=�F����V�V���k�D�lNw*qY��/�����sn�Lc�iW��	Ω�+M�fZ����`���������Aupj;޲Y;��tU*j�ȶ�sʎ{6������YX��uH
�^e8�D�����$Ҝn�q�֏ky�6�VXk�h�m���[�c�/lP��4xƲ���	��V��srg7FM[
d���;f}]�x������jB�C��mΠw}v�wр���{0
2�]�mI�J�	�mR��X�f#X�l\���)�[�����j]����m$��� f[�n%�e�
_�c�/mӋ���Lq\EpnIs�[ٻ(:^� 6=߭�O��Z�]c�+�[��n m�5�ô���ZBߣg�f�T���ռ��hM�J\�Fg2ݜA��q,\�W�c��˺֠�C����ٹ�	�
�K�'i�i�غ�8����Td]�`���7Av0mY�x{sͮ<��pزy�kY�y��t�d	5���J�U���f�#�(K΁a�����c��3{+��5Z��3I.e�-#-��ћ�ݡ��|`^�\�^hl�c�fu�g҆:�Y�mtk�^�ǘ�z�r52�(�)��ț�^�W^����^�\%�!6굺b@-�����&,l�Zz+���nCtp�+6�X�tH�nS�bZ9lE%YbJ�s1frm��ك��/^�ui�yr�'&f����=]�f�I��Nvke�-����">`��Ƚl-s�K�����p��rK���\H^fq8)FU����a��\[WJ�SKnl3�:&�ţֻT�gL�p\흧���[�ع�	� ]=��<��Wn��m�i9��Z�����ɍ-��I���I�Nm�y'Jm�;��<��r�oS��d�������==�z�r[���8x�1����:v�ډӮ�С�j�^�/f�L�핮�\�����\�5�kY��1s��j���Qb]�lJi\��F�k��A�t��ax� R�:��XDFY�Y���D���G=�^��G-�8��m�n��s�l���3̎�����[43C���-�m���k�=��i�4�i��Kdv6𕲔Ie�tC��m��l��K,�l[n�6�Y��٦ɹن'eM���,�cf������l��Bf R)hXAx��Ρe�������	���/;n�]�1eon��m�y��������{w���g����<�.q��&��톄��Ưz�۬�̙�M����,�{y�e�f[am��i������z�ͷy�w�gm�--��g��2.���e�z^e�f��5d���&�{ݱ���<�̄�8��Y"m�[rW�Z�9���x�$�OO�X6��4�d���̺y�s\\��m��c���¡u�"�o;Csɞf����I�hᚈҨ�Zlck�l�]����m�jK��t�5ɖ���d��镗-$v��3a��+YC�i�ݍìnw�B9/gxxZ�x�.-��p�AK�b6mcuSD�4�*��������\���(��)�7�ca��l���&�*�[ȩ�q�;&:�����zk���vιbL�prx.�u��Gm�j�[�l����8
v4��nS�Z@��)Ys�;M\H�5�m��]<x8r_a-I�g�]q7�)f�����]aٖ��,<Nvqr^`��U�(w�S�g��U�{q�묯I
�vw+h�BfY�W9x��j��rA��r��0��K6�S6���ɰ��ܵ�����kb�#KVb��ic+2a���eܔA��\	�{?�>G�|9�nݘ����[KU���eH�Si7��,n�!A�n&17c�7c��Mf�Y�Ws���E��Z�\W�����wN�7n�2ƹ�����.�S4!m����X.5��`GHA�\5P��њ�ʶ� t�ZV=Y�I���
�[:�;Vżq�X�8�˪K�u���G^��<��S��0�k�s�<=��?�}���\�#F�U�x������n܃'E�l#��M�Z��\�m-�bq��=s���ڜГ���ֳR:�.B#�4j1۶����m���tqvwn;�:��Gi�yy�Z��ι�pv�v��2=@6��7L��x�Bx�=�t2�vtF�B��$P�JІ�%��8����o��C;�M���^��g��k�b]Wbx��:ɺ�ݺη ]�	�.D�t�8����6ۭeM�6�iM�f�-k���w�&��{M�|�3��L7��q� ���v�b�qWd����{�v]uN��Ӌv�	��5TBi�dl�b�WC(�a��h��H;XÔ��F�+YF��$Z,E��y��D�)B�maYU�QmX����ic⥐�ah-��6[UDZ��)������<F�ѫe����x{M���{{�&P�ධ�Z�y�z��)a�aՒ������Z�4�7i*V��X�P��R/߿��_�U���4aQ��5�u�aJl9��B�f܏9���[WzD5�]��a��9]f�D��<��<��>:��0�rе�M^G�;��xFk,�O<��fYq̫E����Y��v�õ���1pb�qrN�f��\�t �5�s ŷ�U�+G�z�|�g�V	�E��WfQ�[V�jn����X#YkD����}�,D9�,ʱ2�2�����1��]@^ �@s��و 6���ʻ��FU�Q��� F�	�܌������Vv�������Qh��̉��6*2P㾍�~��{�ڃv{oԚ�=�-9r�ʴs,�����~�{��tG�L�r��m���N0k��@f���S1Z�̺���,��*y׽�6_�X�3!x���K�L:��k��SF�Y�|�cr: U@/�G���b�ӈg�-�->�=�{���JO���VC���c�����;�W���Z�{�%ת����'��O�B���rwV�8�>�h��{o7	>�s6�ϐ^�cS���]�lVU�Q���-�����؝ٳ�DͰJ>ʁ~5ub/=E�̢�2���{�w;�{7��B ���8P�6�A�qހ�#�9��f �̄C����/a�]ITg�"�Fl#�3^�]�b\p�ᮒ4MLw� �@^#A<�ٍ�=�E�@�: ̠�9�f/ s"�>d��C����i�粺+t͊ʻ�j8�w�����G�وm��xv+������ńc%f��l=�nz�x"�u����F��DP@��<s�ꚕ|�eFw,�̫��2�5�p]�qݳa�0E.'v�� �\���s2�2��T�������Xw+A�� .����s2�I&�8Ot!�9�n�N��2(�@Dn�b�(�L˖�U�3,�����w�|�;��s�������Pꬸ=u��f�B����|of���&�A zE5�>������ܨx-��M�����6�U�=39ձoLج��.#����ic�O֖0�s?�X��߷
P/����y s  'E�w�z����0E.@��b�+�*�Z�~�s!7`�̫�eZ32�2�Z8��Wu�_�D��18�s2�Lw�>=���^9���@�l���UO�Ea�s�p�d!�-��yx;�m���i���3m��nh��M�y��Qh�,s*��U3�g���7�����F���1��mf|0d��R��-X�ZP�-8�d�i#�v���?({���w����"�d�@��@�� ,k��Cqp�=�/��͠�=�� ��dP>>�Cn�V˥]Y������̲�:k�W���E��YneX�s(���!-�N�/��u%H;���Bf �U��5�}�M�ʲ* ��54�����n��S�x�<�E�D=���S����� 2+�O��?n�3�<��u=�O9��v��lQ�5����+ �V~�_��,�>��,�b��~O�Z�N*?��qw�	�y��;f,v�)r�c^@�B �!,��t�ݼx^��O%⑙��#*f�4"DéAt�2u�a��3��u������A�4��Aus�>�?sL��EɻQ�$[j��.��(`�X2԰Ng�G�z� �7}@������8�����"sՑQ}�����!�0�"W�H [�Dy���[�V"9�}Z�>�{�^�Uh�v�`��1cp�K�>;�����jŃ-+u���z0�������|Fb]\莗<9�P��j�8��>�|E��<��D�@����,���ŀZq��Kr�Y
��)�qwS]Ì�\U�Q =� �h"3!���o�9ag$P��F:�����2�Q��4'�����$w�ذ���"s:ɱ��u�M��a&�(�/�&i��n/7��`�&y�Ё���{�����dUb앥�N�T�l�_]�sM��5�d]�%�R�G��9��=�4���m=�y�y��� +��h9܎;��F+q�Q���)����C �bRR�
�[�n6�X1V�R�m#2�WmWHv��P�;�&��]��frF����#�R�Rݖ�Vm��k�-�<�F�%.c�Xͮ]�kf�I*.�[v�&^��.s��Mv�6��Ͽ�F�\U掴F���k���D{g;�0�(k4��g9ݨ{�O$��}�"�̏#�zv�C��6ʱ�f�������k>�g�F���,��G2�2�E̩I��k�ֵ�ʻ���U�h]Z�;8�s��f��Lp ����b��g�B~<8�F���֬�K>�c�C�g��LB#&��9��3u���#�U���Lʱ�b�B>'��p;�r.�5ոCh s�q2���ڮf{�gv��c�O��1ހ����)�\pW[�W~����0e���b�i�Y;��?i���f��%�Z9�Igx�Tw�'� A�)X>��Ҽ3����� ��5$���XEW�	lA7d�e˲�2JBvWێ�$v�;�c��Q�@�� ]���2f �5ѝ=N:/��yqVEDx��Il�8�Ah"=�L�,ʱ̢�s�^�W��ޓ��C�I��h�c9ϵ��)�HKs�rZ�/
���ǖ�ٯ�H�4����D��������	N/Nو���sh͎�0E.@��q� - 秊Es/�b|P�=J�`�V,iX>����J.]�����.�ʖ�UTq�@@��#�@�@��ƴ�S���@duǑ�#1&�3���E�/.���� ���,Y��"�v7yGS�V1��,s*\s(/2�e^�ߎ�R4󀃾1x�Fh��9R���ހ��Ȣb�n���V�Q�DH�p���/i���Z�:`KU�WjT�0$,Y�[��땪uZ[/���.�G9e��V��B�7�Γk;"�jj;�b�V�]�q��y�Q���s�q�Qi�E��\G<�p!T��˱�0A�Azkql�8���%�Ҹ���/u�3 Қ�z��wK��-�jX�(,̹�_D\�+��qu3�:q��0dZ�r5��Mo��}�f�GsxBm����G�zC�[@��7`�����S�f��ڂ������K;��NCr�ι_R}~�}�."g.[�V�e�&eY��Jo�o�"�y|}��K�������sQ��El�e��yV#��2�c�E�s.X9�2n�v`�����(Ms[;Y�Dۺ��d��0{�,i�V�쒝#�Q"���mB+Nm�MV���1s���۴��9Խ]�/i��Z��_�S��Qiܢ�2��Qb�DEޝᬩ�9R�!��=-Vu:�(�g�X=�K3,�̫F9�bww��ޚ�s"t
q���|�I�;�sjk	�M�G@=� ��@�E��cwj��E�=E����,s*XfY�s<}\F����\��dgin�.D{��/u��#2>̀����4N��tM��'|A�����8P�f"�N��T���)r�@n�G4�+���#�ۢ� "��{�u���W3��dl.3��뾛��Gr�_�NA��cEB����PqK.�_B ���>��eX��Zc��{W3y����tn��kX+}WU ���x�B �8lB�'�L%z�u(S"��&�xKF�U�z���E���Stm�[���OC���z�wE�f�r�V"�^��+���:3{�n�.DqC��t�76w.�YYe����2�s*���wU���Y�����Y��m\D]��:ʺ�Ȩ"+��;�#y���k��:`H�eX��բfXfW�s,��W���7�����m�T�����8�t#łҰ`�i�2Ջ9���1y�_��3�U������#2��='x�����Z���"fg*���ŢȬ�\�Yps*�.e"fYn�^�.�� ��xNdD]��u����0DW Oz���.Yʱ�5����f�j�}{�e��<:6��x{��������{\3���k*;�OB��ND y���γR���6�����Շ=8Z��{�����ܼ�;������Ԇ�PQ�[��<ɻt��ش��Dϊ5�صUi˦%lm�Y1��j|�z�c"�̜�6J
�c��������lT�l�T�͗@�H5k<���7l�����kX�֡�����0��ǐ'���0fΑs˼u���P�Zc��8�2l ��ݴax,wk����v�ġ�-�z�ݮ�5�\�lR�tv�����/��knsl�9�Lly�s��W�j;N��`��i�;:��=���%�[�9�3 
�b�K�};��2z����Y��a#�d���"Z��>̀3( À���E��]��_B9�5}='8��M���*#�'��"3#^�C��r1t#�����9�� ��N���հm�on#4�}�ޠ���̯�32˂fU����d�nM�����̊> f ���.畱�9��'� xܝ�e�ro��Gݢ�̻̢�̰̯���yuY�;hMc�+�qǾ�sqhTGxOt{\
^@��G����������n�83�����u�M�.�Z
�/�C�ރ�ڪ֦�����s(��YneKs(�}�1]�M���d�"����8�/�����ږ�*�s,�3*X�U����׋x�h4�F튽ʺCs
Cu#S��'s��ϮwW�{p��äY��xl�Z�FDڻ͹q�$����614:7b+e���m�n �z�����4����U9��A;�����#v���Wi@;�-3�[��љ�,s*��\��bg�6��9�7�;D�sqh�}��(�̫�S2���Ƿ���������ɗ�,���Ӌ����D��{�";���ر�:�ڮ�χ=R�z�Lʱ��`��ZfW������64p/!ۂ��n7[�7�x��ِd���ͮb�B4H�b*��WkN�jT&��`�2��l�V��~�b9�X�=r�V&e����7��sqh��#g.+�5t���T�e��U�2�s*�2�����r7&��� ���W�����`a�}���/���X��h3�a�'�U�$yʴC2�Lʱ�e�H�`נ-������h� �����A�,�tj�u/y�
ܞ|�9^x���Im@i&A�����=)!�dK��kLS�G{���꽔�~}IX�eX�Rvk ;$I[e�ٚ^
7]�_D�H'ml�n��F�H���6�N���rض�l�6a��]�"�c�g3�OA}���Ϋ$f�+�a�}�iv:�{����8=�/��27��5<�?n�1M���ӗ��/%Լ�3�%����n�6�N�j&�����$ه��4��zcYZң3��/�e74W5�0y�5��ӯ�*�����z��8�-2��&Ż�A�gs^^���1,����P�ًkoRf��鸡�T�ٱn3d��5��H�f�ٷ�,�9�~�w��1��s$W�����U���˚����ӫ\�εT]�z
ȑe���|nb�;�}[w���w���[Ul\ܩ�:��@�0��-��j*��~�ȵS$��p�[�h���.6�,q�5S�5vv���v�P�s��0V��{�	�f؃��Xf������ ��x�-��Y<���nÈy��Ʈ����P�h3��_v��(Nl=��n�U�-���i{��z����^]�N�۝�Wy�����]=��x�e;��珴�c5�<<�-?g����Y^��+���|�����V�kR(o����_]��e:��gS�Qv)Z�kG<q��ww��#��K[���X��<�<��<笔,F�'x��ץ����t꾿���?�k.6'd��Ay�6�Ys���<�y�<�<���޼盭%��QF[q6������l�ŵ��vq�k5��6�k5��^On[j%�gE�fض˞��l���&�7M���n�l�m���Ŷ-:Kv��lm�0���g`���s�Ǧ�lͲ�3r��H+�l�"s�tw6��d۳�i��km5���dܛ��6��!e�ݮ�9��Ynm��IͳB�j+k1��4��+4oo=��Kƶ��L�v�[[5��ז��'L�vfkj�f�gX�;l�#�[�c�s��n�3R�iYLهmY��,�^��9�嶔��f�f���fp�r��m�[h��ݜ�M�Vۧi�+f���mvhvٺ��j��xQme���&���"�]Cgr�U�Y�H��d�߮�(hRAaS��i �r�I�
H)�.�(�r�Dt�RZ߷U�W�pn�H<����n�)4 S��l�d����Qi���?W���w��i�ku���Ak.��
H)(B�~�P�MFRA@߹߿k��ۿ�=���?�$����R
A�C��H.� s�Zh) ����r�����XW9p�Aa���Qi7�|�~o��'�S��pw��|���{o�^������ �*U��ZA�Q
H/;wH)��s�f�) �s�ZAa���gy�+����ݵ�m�Bc�ض֖!:e�k�zۣg(�p��,ښ�?�ygK}+'�/B�)(B�w�H)���q���p4URr����3[�V�P�і�����#� �<	������^��ݣ�i�]�R
Aa��p�Aa���Qi4!I��S�]�P4��Xs�t�R
9E�Q
H-����w�m��淮����XgjβRAB���Ѥ��E[����NC������JĀ�#X~�B�42�
�H,4�^r����f�������zT?v����H��R5)�������XW9p�Aa�0�r�I�) �P�y˸
�?s�q�Q�>�?��U��g�}x~6�X_��$����ZA����;�@R
h@��B�
ACB�H,4�]��
H)3���߫;{�����{�0��d�e$e�Xi ��]�Ԫ ��s�$Y��㿟����޼�ƾ��e��) �߮�) �`Nk�v�����(�^����
���p�����ó��@�u����]�ޗG�����T&�^�mƭ�Ge�(ǙBwLF]w2k��T��_+�E+��U���o}��8�XxaH��Q
H,��r�ZAH,9�������r�H:(�$���S@�L9ʅ��=��]{����9���x>��|>9�V*���с��KA����̨��� �fy�y���[���u��ǚ�uk%*"�Fan�V�0�Q�����&�#�Φ�Ya6���@��Yђ�������XPg�H,49�-&�) �����������gv����<m ���?�
CZ��tuk߱����@�TZA����~���AH,3�f�) �s�ZAa��^r�Q��
JB�s�H)۹]���� �8�A{ʁi ��*�]�N���k{�[�Չ��dG� "(d�ߪ����
;ˆ��'���g�N����g7Ww�m �v2�z�Z���C���P?v�H:��Z�.�
i�s�f�) �Hs�i ��_j�E�&6��-�vb�+��
#����H))
a��H)]�H,$���R��CI�`R9E��) ��}���_o�ݓ�����$��ˆ�)����) �������j����V{o���������:H)
�ߨ���!I�o�}����}�H)�
aܨ[42RAB���4�XhaI�(40�AIHSr�l������Qi�����������w!n�G����$x7���k{�����5��@�(�� RAe���@�4���i��
@�(��G�>��-ǀD �7����o��V��s���g����A�ǽ�ì�}g�s�?x�ҕ`������뗉���m-�0��'���و{�������z>�������ЃY���7�X�7`K\�u�C��љA4��LZ3kye�RR�]�v�gv,�����v�l�+A��ә�gJ��YE�K��v��u�T5��!�σ4v�ږx0���p�Z)ׯ]+��l=j�a�˂���p�wW��/G�i���N��m��8;H��z���������u�u��4��xpQ]�x���H6��n`����:�Jr�cR�VS��	Mf�5���؇l���f�#bӪ�QO��Aa�A�I!U@w(���D) ��kP��Xs�f�) �s�ZAa���~=���~���/k�6�[˰�
K��;��s�3�H)^���I�.�j���h*�CI��9�-5) ����r���RAa���]_۽�H,1� }�-&�) �S)���(���V�s���o�W������i!��ߨ���!I�wZ��ЁL9ʅ���g��m�{&�
��
AH/]�) ��)��P�M����Qi����]�R
Aa�T- ��#�t�马��_���v�l:�5���n�H)��)��
RAaGyp�Aa�9�- �M2�r���) ��(4�
C���^�Wo�߹���R
Ay�kP��)�{P�i��
!�Q���M<��Ǯ�]iN����dx�/ H�R~"���ɦRA@��s7�߿��[��$߮�) �*�P�At0)���B$��p5RAaS��i ��
@�(����yN��~�}�C���)��� �V|b/^����"�`�Y�M@:H)
*����H) �wZ���Ü�[62RAB�9�4�oO�Y�������]���!�z���^�&��V�pި̰5.���d󥳥��/AH)?!L>�B�5RA@��ZA`j4�^r���
A��9P�@�>��ߍw}z�X���q e�Dx<	��8Gw��]�V��y�^ �$�$��$aH��B�R�]�P4��Xs�$�U�QiTB����p��_U���z���E6yf���݃P�f�+����̹��*6m(m��#�3F�`C�cLh�}�����NFƚ̊�	�H}E(��������
AO�0��FJH(R�H,5>�=_�>�߭������H-�� ���0�ꅲi��P;�- �5H/9w�������kd��T3u$C�>��R4�Nr��R��I����Qi5���L����H���<ъ?|Q�s��w����}P����T��ZA�D) ���P��Xs�f�JH(R�H) ���lRAIw�����_�·�~�P�N����_�f�M$?]��TAH5P�*H/:�'~5���uaW��.#���g��O�]�P�RAaG���=Y�R�E�Ѕ$JO{w@�RAa�Pi�AHUP��R
Au9�j�Rr�l�;ʷ���-޹'R
C��I���~�߽����~;\���_����]��$�Sߪɡ��P(�l�A`i���p5TAH5P�*H/=�1����������R�ʫc6�ԍ�V��]�4�X���LKK7T٤^���Gݪy�|�O�?X�YL��p4��
�ˆ�
A@�(���Y6�y˸
��Ʒ���{������}A��AH^��_?er�w~�Qi�!I��j�Rz�l�%$(C��I �����RRÜ�[&�RA@��ҷ��i�����XH.�wH)ECݨi ��?{}k���߷�=��_ߠy7E���*2S���	) ����i ��
@�(���&]�s���w���&�S}���i) ��Pj:H)
*��h���D) ��kP���Ü�[4��P9�- ���Ѿ{߾�?v������!��t�~ޜl�L��q&�n EP�3 ����A^��]����ݘ��3���iZasg����κj�]�ú���,�V$�|RAIB��ꅲhI���M$�����
Aa�T- �`R9E��) �=��7�����&>���RAa_�p�Aa�� ~��HRAH/9w@���o����}�~�������?GI!U@~�E�B�g7����~�y׽H)�0�ꅳQ��
z�H,4�]��RAIHSr�l�e$
��H,$���]���귳���`G�txI���}�;���u���@��i ��%?�]�R
Aa���I �s�ZM�
H)���%�C��^�_���Ϙ�(��&�g�8C;Pr�9���.�:!GWSnp�kec�Rk�,۟��A��AH(��uD) �{��H)�9P�m��
@n��O�����W]�|;������%b@|| �G���n'�ꪸ��G·�L7���~I��f�
AH/�]��Q �P�*H.���Qi��
Ay˸
II�W�^ʽV�üK�����c
@�tZM!I��S���P7�k�g߿7�y����H,5���AHT���- ��Z�u�
AM Sr�l��~�y�kY~�vJH(hCQ���C
H/=wH)5��B�4����Qi����]�R
Aa�W�#���yrzU���ȏ�)�uF���� f���I�2S��� ��B��)���i
H,�2�r�����Ü��t�R���xr��w�~����H:(�$���H)��g��2RA@�(�x�>�������.�8wUS�=�?}��7���������V<_,O�;�:�"�-Sۙ��ɩ����U��YV#U���3��Dۑ��C�{M\��u�[P齚�1��B�d:s��>!���9�-̢�L�-̪M��=�k�=�Ӯy�)�o�}LP���=� �k��B ��+��9�*w�DF��M��E���h6I��xl���m�٭���e�F1SZj֋骯"=ʸ�9e�̠��7��:�]�Tk�
��;��n�3����*o��0s(���\s(�&�\�_w ���Bi�oS�����R���8�ty��fc�N��p���z��=@ߎ!���/���5l�~���w�������b��<��ƀ̊#2 ̊�'Ҭ!��{P�̀�����k�qo��Ok�*��;�� S�����}e�~�D{�-3(��Qi�R�2��o+�x�m�H��U ��C�ھ���M��"�V�9e�̠��+>���iټ�Ά7� S�;7l�ƏF�J؃Q�"�	�<΄���+������"\6��P�q�Zp�H2o�۫���=����7sN��e�i�x���0&$����̦���X)�uҭ&����h�Zu���l��B��.ob(��N���v��t���K\b'S�C7n�B�lml*�TF4R\hn}"]�ҡ���ۇ0�Bi�v�:������r�B��L���@V%([M
^0 �`^�5����E.�ed����#jѽ@�0���Bk�Jm�%i��`WWDَڥ����~�g�l����±��c�Z�C-������k��P6�,k���}_����&�e��b1̣�����{)��nء3��p/b�����mǖU�Z~_Jb��s��K�G��Ƀ7� |s�UϨ��}W�z�0���q�,G�s2�ܬ����(��Yb>�}��̊ �/j����;;ٸ����П�**h#dq�A�k�2���AJ�e�_T�n\h��E��c��Uh��=kV��jر3���Փ2n���=�;��;�,�̩�_#�e�3[l�:�U��D��zN�nu^	����U�bw�dG�e�eZ"fW}���nx��~�z��������2��h��Sh�m�twF��o+٪��f�[B]q��z�c-��e���2<�b�ק����OAoT׮�=y�c�3sf���}4�ݫ��1{2=^#2�"���켙��0���f˵AvѶ��p�8:a@hQ��b;���t�k*�#
q`�l���؉�o"o��"�Fv���ۡ~7��Gt*�ه�Z�v�U�bg��@@���Z�:�w5��Oz˃3�\�*\̰�*<Fb8������tz*��a]{b{���:���Qne\FegŞ�=�]�7�,�/ o�Fb݃��_ڈoTк�w�x��dA�0bhB��	�j����V"�Qh��[�W�*���x������Z;r+����QpNr��2�D3,S4f�w��fg
b�ۃ�ZxH0��E��K�j���h�T�u��JMV�j�w�،{�Zo����uK��ឳ�.�8�sn���r����=V"�Qi�e��EĦ"�J��/���<���n�s�w�z����h]Gx�� A�h ̇�"z������_��,G2ˎeKs(�d9rN�H��əe�Q�EOK�9=�X��:e��~�� v/y��m�wL�J�nh����w;�V�~�@�ys�~�����*�n4v�V1aO�{�/�,s*\̲�2�O���k���~���A{���o8��י
�iȗsA;�I?.o.5nZ���G����Zq��Ol��i�BZ&O�mf���N�W�jf��q�z ��dP>#1{�^��6wH��yKi�!)9�9�ۼ]�/$ah�ܽ��/\'�����\���^Fc:#�}yn=���
���$�dh�ȼb��t�q�[>���U@�A�����j�2҆iC��z���|E�@���Ǯ+�y�D�9�c� �@Dms"�]��lDt�����Qbo�.�As2�2�FfY����;uJ�ա_7y�5
��Lк���_��)V!iC%���u�C������Gv�@B����=�4v��aL ��Dga$lMӎQ��ꕧ6�RN��qjn���b��E�T�݋�ȫ�:{"�{]�E��Us�[�q:z���Q��r�Z�S� ����t.���:�?HB}럇��D�l���h��/�Ve�����:r����2����~�N�{p˹� ���/fEÁ5�����������[����s��C�������v�Tu�����iI����t�s-���K<�y�@�����	���t�W�ff��{p��kW��}���GYa�W�fe��U���xIw=�8�9�c���� !U,l��Ӛ;n�h���'� ��yȝ��긖�K�9�9����Q��B9��zQ����{�7y{�f]�qy���.9�b.eg�k_l���� �� �/#�Fb��o>��W9fT؛�p=��a�7��2�jŘ-(`�_j��I����c��vGv�-�xg������@���Z39r�̫3,�V��}�;Uˢ7�\�x���r�Gp��4=�|����� N�%GDq[{�*��Z��6"����n�5�!g�`o��|����
�Hoݯz9;d�X�(�|�\C_i:�~�}ע��ͶF�	�&�j���NS;��fN�F�m�����n�ovL�Oh��'����������ƕ�w�{KZ���?L�q�#�2ԩ���Ӏb;����{հ�7`�x��9R��2�r�k7#5�0�*� �=����>cvM�u��i����H���N��3ٸ�+a[܇�9�N2��;bI@�dԊ�2T9m��TN���[brFV6��TF<=�o.Ƿ��휙�l��yFoRx��,�!1AN�u^�&_
�zrif{�����)�^+Y=	�͗3�痼48���$�*��i4oV.E�Фf����G{�|�^�yl]��Fe��ƥ�l8Bu���@�z,��������V{�xk��c��By����$x�qg��bzj�i��<���s��2v���e��W��Ϣ�Gz�x������
��5qaC�=1nl��ח��J�'=|�gBE��2j��^��f];5�ȊnuT.����x�-lȖ��@�T���V�-ݔ����n-�x����og�����w�;G�T�%���%�[���Daܛ8������h��67"Fлx��4����B3_q=�&&z�=��j����[���z���r��6�]Pt�r缻����%f��1�Ǜz����"kk��k�֗h�ŖA�c-lڈv�m�l��(kgGn��BI�G;4��z���Y�K-��2��y�ms�ٶp���)�{�$s�����,�4ֶ[��m�LͭrY�Z�i��3t�bPVv��淖��F��k�^���[cl���7e��l�ٽ�"<�Z�8W���Y��a�6����#��Vr͘I�,s�^e��ppIaXe�P!C6�v�3R$gb[i9�;[`6����:����k�gZ6đlnp��6m$�l�ͱi������i��-h�d�7��Zm��u����mfVm���IJ3��mv[`��k�ͫt���-��[Z��	�V�Y�b��9#�,��;m�4fg��=;J4����jӍ��;��։�.͘&�ps�ͬ��Y�����{����zʥU"�UB%RVs�S�Ӌ��V��]y���ɴ��u����Qhāf�rPU�K���Li<�Z�#�.�\��]�'�n�;uֹųEǎ�8�1ъ����m\��-.�fne��K%�RT6�̱e"H�(�a���l���Q��e<�Oni�r<�C��贩6FB8�cYb,�GB�d��Ʋ//=�d��4�c(�ˮ�k���N�/����r��m���h���F�e	f�y�h���I���n8�{8��v\��/[�<v7`'nc�"��h�����G	�
���e���ȖƎB����6Ǟv���mV:�lN�q���/8����.��z��]� �ɧ��,Z��T�nL%mNvK./X��D��x�6�n2�W������� �`X�ʜ�t{uF҆5�;���ة�{uqc�����Z>�0譲�uKl�ԗ�\@q�`-�9�70Z��q[@��vt���G6�'����l�!i殆1[��C�.��x�j�í�:����ѣ��۽�䱣+Ξ='W^��ڴ�z�X�]�V}�v��.�lGOH��0Ձ.t��\�L[ŵϛ�6x������x���;C&��e�;*�nWuY'^h��{=�1��/)��_Aˋ��}�;Zue�;�Y��X�t�l5���0n;j�뎭Հ񭕉\���h��s ����bWst�v�E͚��P��n�̱���6���X�V�����'Zz;�0��CE�@��)�����⺎����=��_}q��0�+c3H36��E�5����}*���]�1��d�C�ֻ��U�]s��K��A�^�<>���n)�u�ۥ�-�If�̺X5�nuH��l��݄�[������{F�^4*0w%*�i�b4\��u��{v7i1&�(Ӛ��J�����+l�WW4M�R55+��3H]�c����#Q���յѱ��٣F;�n<jxzD���x���/SM���R\Eɛ4�lnJ����5�-&]�lԴ-�I�I�w��Zi��fV�1����"8EܻK��JJ��Z�f�5ל@�.z;:
���cn���5\ѝ������}�tRF�'d�3�듥��h4��ٍY��2w)&�e��u�Zvi鋈Yk,Ϋч]mزkf�{P�z �L��'nM�6� ��ܥ�^f���6�8�խ-�hL���e���e�y嗬t8��k�K������bU����;Cs����r��ot܌�M�x��n��Z��Q)S��/�#�5̅��3�{�+���e^�6KYGdF.���8�u�(�v��"�ӋZ�֜_҃��b��)�߻0fB����Gy��p���2���w� �B �1��ÓB�ō�sf��6�C�U�$q�,̲�ʴD̬�k{��l�:;��Q�Ή�ΗW9�¨|q/BҰe��Ջ=�S�8�8��{2�E�8�}��*�ٲZ��;a
���g9�=ۯC3�� �p��H�xf@����ݣ�+FU����޼�W9fTߦ���Ј>���b�Օ����g�&#3����uGB��ӝF.�@MK8���gq{l%��.&|Dt � �/fEA���Un��/�����h���^����Qn���� A�"3!@9�����1�����Ǭ/���ߧ��[AV��b�%X2�l\�DR�A4�E�I�h��f���z�)�߭w��-��>e�O����[ﾀ�3~q_>�q9}��/&8>��-��̎
���%^��>��\�y�̹c�V�̲���;�;��ڨ����7r�6.���"mbi_�8�ZW�9h�UnԾ�6���H ^� ���S�2���w9�¾{` EOv�Βm��ڥ�7����,Lʱ̫FfYi�[y���Pj�랏g� ���V��.k8a�7��y�@�^̊��g'6Wu[ɓ���p~��y�2�v��#��@����O"v�Ub��m����T5<v���ts,3+�sB^������6��6&�E�伇5�/�{n�x=���2��eX��Q`��rj[!��v���QЬ��q���놇�T�谯���Df�/�Y�wl��#.P@��D�"3 ��b����(�Aea+:gfUj�����T�_ib�O<���n�n�o�ʚ�iW���#��~U�Uâ��K�frI�Y��̡S[˭f>�� ��+:��u��V��كw,BҰ`��Z����6?ߵ�s�#z<�m��'o��}��u
�WBn8�ޅ�3»8�ѹ����:���!��1d���۫x�j9���x0V֍����a_ @=� �5y�C1qtuV%[O:Ş�C��}*Q�.^�����s ����J1�u[���u�5��\�W�#�j�a���&d#�ᘂ�8���EK���q��=���Y����>D��ݫfe&e؇2�#FZ�N�GUU�sA�!.�j���V�ºq��D6��#2<��8}l |���b�C�N!�ՈZP ��mfn����'��y\8VN�9���k�6^�X��E�gnX�U�a��-,}g��\5x������|>��g;�W;�/;ۆmǻǜN�ޣ��y���ظ��xxOx=&�21"��8F޺��Fd�m�$bNl�]
��ԡ��p��}�};��P�±�M띾����$B�ɿW�}��3�b9��^@�F��;��1��S�\����I�Tcx��>��:�X2Ұ|-Y �E��g��A㈝@-��,�3q��N��;k�ʛ��`�x�cJD�[�F۝1���,�~|#c��B ���g��s��z���a\
�Wu�b�G`.��2وȢ9����Q�[��������q\��'*=�<�"md	+�=n��~�wG���h�\�2�C��L��12��E�	qܝNf�ʙx�|^�ȏ}V#�Yi�V�3,�s*�޽ȃiNf�b��yA2���_Qч�����_@3:�r���ݛ�rˌ̲�s*XfYc36a!���9z�ܠVj���E)��6L�{�����@�^�m�Q8
Iʁ�ө:;{{��	��6�pMZ�ι���DV�ĸ���P��p̢�.4Yy�x��t���gc���:�$ A�x��SF��N�Um^��an:5�`;%�A9&Z�ZM��Y���E��Fhh4�E�K,�L���S��L��5�F���[�1��#�o��8���j��$#L��!�X��	��nk0˗u\�_B���W�ݺ�n�l�M�r�Q�!H���p��QN�}I6�����k.:�.YM�%LnhЪ��#ہ�9f8�h� ��ݚ:����>�[I�x��0�s��^�W��vgoQ���u*�.��q����	̄A�A	���=��2�E�y_9�f��;a��Z��^^9�#��E�"_`9Ѹ�o��[��n�eհp�;Y�¾{`"-ǳ"d�3�|�l@�}{x�������՝)3�y�c_��x΅�\R�z3a��G�΄A��d#�8}�Hi�y�F�N^�X�s0"�vEFb
]Ƶ==��2�E�3� �B"Xn����<�`�6�x�� s!x�s /Fb�D�:�sjȑ��G����87�`��v�E�|�=���҆ZpO�?i�{���G�"H)��8�^ƭnʕ�X�E��$�u�W���K.�����WM���#̫������.k/����S}��NTp ����V�lí����\��U��Pf}b9�X�ћ?r�������/Z���Γ��JhyF�VOi��ni�*��j�1�c����i~��&C[�}�#�wsڸ�mU��N�fm��~  ����мF�	ێj~��څ2�b��p ��\G�e�eV����w\��Yn���Ń�����iͮ��{��3M[����Ά��aWy{` Amy�@���#2!\��l�dFĐ{PDg@f!9�+�R�ѷ���GNtjS��Oay���̵�N!����&;����T�܂���S���P���{ѽW�#�U�ܲ�2��e�٭�:��~��W�%|��5��1j�����V^�CR�B��1��s�hav�4�Eq����e���2��̊ ����rc��5��q�(*�7T��k�j�D}��̲�̫��d/2`gYGf��]@����NF����3z6�8������Ȏ^e
sB�����:q	�1e��-+�'T�S3;�WM�fX���t���v�aZj[�4��9i��7�^���ͬ��lC���wc�'65Lͫ�jt�^�I�����P�*��_x ���>�*[��q�>ބA�"3!㘂ʕ�����ײ��&z����P�]z�0>ڊXk��
� A�0'�����n��o�S|�處b#�V�e��3 DʳZjqɽ����Z�q<��]W�N&� ́�7̏Q̀����4�{���\K�0X��]��Kte�K2&Y�R̎c�.B�G1�{�C��O���O�@�����|�w鉙n��Z�����NoY���˂w*���-̫fe�eƉS��s�Qdw`*��kn�J�]g4PU�@�����1ič%�vZs�b.v�G2�M�[˛)�os��DEOD��=uZ6�8���>=��8�Z~X-8�e�埼�]���]�����^��f ��͔��wLL�w".8A}�9� Ѭ[����M���wػ������u]�!ǫ)�l���^K�����1�G�W~�X�D�ݨ�j�U�u��ПBQ�$��a���Ov˃�V��-3+���3LҚ����Q_���f�ќ��x.{�Z&r幕`�e���^�����~�:T&Xڑu����ʚ흧�K��suq���+�N6&��ￏ�[��e���>d/�2�r��\��En��UA�q����m򾩸A�#�H̄�@/f@^"�2���cV_\TǕǳ�'���]�;�&&[6��_B �Af�u�q�d�Yc�Ո�gj�3.Z_�2Ңеi�p~�_�Z�I��4{������%�>��9�.9�,3.^,���uX���|>�X�����1r����Tq�=%�^U��Xe��j�fQ`�PX�Qne=�{���s�h/[Az�{�;;Ǻ����W��`�����-/���a�@��׾���%|����C���-�ʋ�j�7��2�s�%�fĶӞ�w�4��${���� �[b�6ȷ�ϗ��xx	���K)4a�3b�E�vݵ�::<2��u�nn�u�6����ƛ0Px�4�LJ�1��4v岱�1���\�<K���T5S�G���wg��k�܈݋Ź\�ݳm���:�Ѭ��/5w����nJ4�R�q�9�g���HW�H�����7e�<�cOk&H�ASkZ�,Ʌ6u�U�H��y�-�m�qy�=���n?�}����_����]d,ĺ٤��a�A3-n5�ιݝm�b��г���Y>|?|#/σ ��U���gژΊ��&�+'{u��1Ϩ��*�9�X��,c�V���Ts��Q��f�����K�3��觫��p#�͠�dq��26��\����h�P%v�L�ع�."�Q`9�� f z�퓶��r{r&� �tLN���V�,G��G�e�̹q�\̨��ki�+�DG�1{�(�Fd!O�!���3Ԣ�D���ǜBy�(�2��l������-_e�`����Ѡ�L[��DJ��X�+��~������ZUQ�;a��fEdTb��<����k}��
����i�RWM���5<�z0X2�ۺ��Y%�� ��,pGOG�����_<��s#ِ(S�͙�:;OI�xez/�W��{�Ue�p5��;��f\̯�D�+_��h�q��˳�S��GBqRş��t�.jƽj�64����fT!8�oss��nog%���e��{Wr�(�h�וw"�$������P���Ѐ ��B�bC3�홌�QW�ET<�"8� s sT)t��	����-X�}j_Z~��)�y&;���egM.�ZUQ��X�@�B�i�V�I����93�w_�|2ӛ��6g���6L��+�p8Ё��f����U���g�w���_DS2�L�,r��/����70d�o���>�鿚2�H���p�>-�@�B����쟙�����O��Ɋ+7"�k�#��t��wm����Y[��j��;�}�?2��Yy������U�u��+:ip��)UGx��9����e�5�O �;Ё���d
2n��
�g#2�ձ�n@Bw�6g��|:���(A��_B!��U��\��h��]����H㍉�q|-?,Qs����?'�~�l~�+�o��tZʅ�<����b	��V݊�����V�dM�Qu�Y�=�2$5J2{={�9}�9����=WC��R�J���{gH58j����8�eg�="���>��>���V�65�����=&q^��i��}ȮگsK��P��v-c'��ٽ�V��?5����\Z^�>qJ�"��au�)��%�)�.ĪU���M=Я"��HlFM-Y5S�æ��e���ܭ�� I-���޽ ~e��R���۷fC�f�2�rX��]�y�^�>�kr\��6vkV��{��&y�ҍ�&����^y�/|VYji�a�U����=�[He���e�t���-|�3���ސ>��k:��u��i�=�[w+��R����{b*�L�'E��{V��b��r�wb���*��lh�Vk�*!����=�<�������ޠ��jH=�8NaN�yN�o5��{0cI.b����	3a�7�Zfo�iڛ �G�jF��^����*�W�)|��/�՟�Vw��ɋ\���'�g��P�O��6{77z�wy����y&���z�?,)^��x���ޚ�>ݯϰJ�V����æl�hn�a��wsUX��j�e�����9����vL�9: ޲����RvuU32�����M��+�`����w2�ca���Q�5*gbÜm��p�#I��WN@���G����O�*�ov	�#�`=`��4������/�׎�0u�y�|-~�X��^���s��'C��W�g�k,OJ�Y�����%*RR�����4*��gEY�Mj;��$Λ�m�ؔ�tۓ���FSn�vݶɛ1!r%m�͜G$m����*�����f㱣mز̓Hm�6iL�vetmnP��"cu�[v��kgFt�[dmh�$��";j��6�왛���K;Cv�v��7n�������ls+.k[� �;"&�6k�n�C���$�rm�B�m6�)�oz�N�m��Z�"um��9i''8�Ҷ�k;m��m��!�۳�G[d��8��mn[ZI"��nmnS�L�������m�Ҋ�rZZ��)�+,��vբAL�ݶ�D��E$N)D�/;V7n��6��ڴN�4͵h����$� ��mN��de�1��^��Fѭ��(6�J"����3�tm��E�tA����w����gI�P �}�����qHvޕ��މ_ ����%�eX�3,��.����B��7> ��#�Q�x�dv�=,�)Z%��UP�>Sw�j�k���0�k׺�f�6��be&8��V��k����&�wa����O	��P�}�ݫ9�X��,̱�k}��-��}x��3n#�B'Nj;�I�A�X�v��;�9A:�'��m��ܹ���Eq����Yo��d �qs!8p��1���l(��Sz L�z�����#b�G"b�8B9��n5�'���,�4��w!Y���s��/f"� gO�ͯfW��9y��`��;ς�<��,d/�u� ��1Q��2������_x���V#̲���q3,�̄�HICtmv�V�du�^=��$fEv��G��(��sz )��=�"]�ޚ�ޜ��;{��nl�*�yY��N4Fo��lq�~�0sp��f�j���iC�B^��+Ѹ��R�9�L%�5�r˪�������h���X�˱s#�1��ð���04ל��o�A՘�};�3�Kو��� oB �h s!A�����u���CD�Rnٴޣ�ے�8���gF��:�5��Ṭ���|,G�Q`�eʴs,����I�xz��6įEr��6\�1cu�W:0e��;�����2R�)Z�)�RJ�lx<���h��+�Z�pݐ>�x�E�=�[bj�@�uy{v1xfW��#���uB/9�k��s"6�B������1=�y˙��13*f}ek�V��8$1Ӹ����=��b�1������K���m�A.f����ˎ�e�eX�fU�eL����^��UM�D�ET,�<�t=ԥpqu�����-��fT�fY�ߵ��h�U��]�6�SʽK^��A=�la�c{��k�y��F9��`��_ި��ּ����̚�t������y��_�;�I�翲��4���i0���mÃ=��h�3�Ƽ%1�l[��ŵ��b��Nĳ'�F󬋳�Xu� 6�Yn�k���h!{g	��Mg�6X�;� <������%�������U�A6����kn��N�6�<�G`�1]���u�6��5�0v����'k�5��zvm�ƅ�CA�Od��I3�crb�"�K ɜl�svY���Gd6���<�B����IyY�s,m�6җdHs2;W:8�آK@��cǾߟ�%r<���#2>#19s�/�w":���و��Z,�C�l@�A�A�@�r�X2԰N`r�F���Ϗ����f�[���:��p��%
Q��<��̇z�<'���O@^;P��@���~Zp��1些�w⡇�>Zg�YT���gh3+�fe�2�N���gdi�Q��3�"B>>�AxN\���܈��Q/TD�{�Z���7�cz�X9�K���X�Qh�\�̯g5�9� ��3�5��K΢��%
Q�>�\G�e�eX��;�iؗ�6ꪥ+*cB��-�%�K�����[�K8���W.�w$��gj�GyE�w�,s*[�G��U�^��jyZU��6�@ə��A�-�j�2�̫�e\�}���ob�V�ɿI�x�ە���G���8�9��N����<o���e� Z/���H<C�j����ɾ+"���ޚ7���H^t�&e[��\�ٯ{_���D�*��DL���|A�N{c�����pL��Qh��,s*��Bgfy<���ѳSo��5�P�^D}�̰̯��YneM��n���Np���o�?���Lѻر��踛���ϝz��e��V"�B ���*:w��1���������K�")�SA���̄���E��>�������B٦�B�bmn��F�En#.nX�	�kM
̀28&��w���f�y�@���v�ඵ�&�J��^�b��]D� �(�9�� �@z�~ݳ�M��r���S�J� >خE�m�r�df�#��G@C��5�G��DVB �8Df@@��G�f!��E�d��}w=�q�,���?ʽ��"����� �{O2��Q�Ň�ڌ�� �O-��$����6�J��$kc�_{���������s���!L|A��̄A�-3.Y�G������GQ���L�n��k_�"k�j8A}w	���)���Y=�Hy  ^̏P�3,��V�}䧞ގcu��ѮQ��J���q\�Em�&y{ "�W�9Ji��o5u��V�����q"���մm��S��;�`v:��c3�jt�9޲�`�0A/#�͠�̄|}��K7g��J��U�Q
c�2q]�w.+y��$we��V��E�f\��eC��߹��}�[� �B���LF�k��dM`�,��Ј>x�Õ&�S[�qC}>��/at"b�2Ȋ�ov�Vh�=o���0s�W'[e	�@�� #��D��ِ*\[���}��EZoG��B�1�t�\�][�3����������{_5����i{�B�}��/C�Wd�"��%��<�g��X�����!�cw��ݞ��Ц8VFj�"�t��]F\�ɂ1� ����|]��A;��2�e#�.9�����U-r�kϦ#����&�R����̲����g��_l�_��R3�6��3��g[#
ݬU�<\��I�� �޺(�s�E��Q��xx���eX�㍕����Cݥ��-���AD�;ˢ.'H��C1���D^�9��es�ѷ`Y���*������e
ި�1�A����P9�+cQ|{'c@(ḝ���\D�ķ2��f���W��Q����FU7�QȚ�HZ� �Јy fEf@^9��v��}�6�2j �2�^7��� *��rzݩ���AL�"M�6)M���y퀈̄A2<�DfF��3^��ג�I�V�˝�x+z�Ǹ�{�B��-9�����[�c^���J�Z��V���$;�7��=;��e9ا��b��>>�+�ڈ���,�~cHmة���+�x�L��r
� ��>3ne�d��x�,W9#�\����MN�::p�L/YAk�M6Xitm`�۫҅O/R[\K���Vm���u�ڑt��4e���N��M�:�7\>�^{A!�A��:�`��Y���a:4r�wqě��udeI[d�4�ж`N5+�V����e dQ��sk���v��-q��Sz�tGDsini�h�k���}���\�K��4WJ�Nl���m��I�����G�n0e�>;P[@fEx��
i�Iښ��8TM`�-G A��*c"�n0���V�fYq̫Ds(�߾�3����}x0�^ ��Wn+�����C�٨B���>�-;r�^���������f��O�V"�j��-3*��5�Wnm�Y�]//�Q�6�b�Ot�Qc�Ws(3>�V_�{/^�eN�9��#1=}�vgm�\*Ue��#���	�k���,B(��Ȟ��z�X-+i�Yj�𴃰��:�˦&(P=��u����\��M$��{  A9y�^#2F��p�b�b_������ֵ�^�ݍ+���V,a���0u��������@��c���߯��e��gσ�ِ*�:~�o-�]*/6�������N�Wqw��2Ӌ�̴�Zr�-8�y��5jUh+L�-[��{��i�J����؝�X"�kB+oS2�D�q�Ê	�oϖ���ԯm���j�K����9���g.�� Ns���XA�Azz��N�վ¥VQ�q�/��Ne�e]�g9���5�,wڴG:q|0e�����i�؏�:T��tR�ݞjv&�
y�{ r2(��&eX����U_ؕ�n�D��X&�W� UF��WX�#�E��B��}� Bw;�k;���G*���s ��̋U�Ո���h
��z�ruy�]>���4n���z�Ùe�eX�̼���v������(*hp���X�.���ŵ��GP�z���oL9�J�Wg��	2z?z�F;�,G�e�eZ �Qs��/z|�zZ�����2�A�Z��@�G8�/ᖜX2҆������L���T��r�{Q*/6��Ot��.9�׻i�{�.'we����,-?;VEQ?T��ߵ�z�w����#EK�%*nV�"��ոx��K$o~Pt4^��K�ZO��)���2v>ƈe,X훃��y7��� <Tov�Ozf�� �� ޠ�#2|>Z�`���`�o*�#y!̌����z��+�\-��3�2�S�{ "2Eo-������HG�{rx�8��Df@rd���%�/e����^����VfڅQ����x�p̄�����|}��}�#��K��lZ �i�.�8wL�۵�\��³lvJ�m/�̷�� �t�s#�1����cn�	�L��B�p��������E�`#. �8��19�b.8�Nn���k]֍���oU]����fw��P��Ƿ`q#H@����WBŚɇ�g
��8�2Ո�8������s&��݈�Jny���O�n�M*� �?2��-?!EZ�g����V�TZ'k�q�Ո��kϳ�Z���SS�1�@ �B!�؈U�%>+���7�]uo�t���l��p0}}�#��v����VG^�A�"���@L$%�x�-�ޭ.��;�+��v)me�������%c�,�|�r�@�(s�"~�뛙����3#O8
]�Q�K=]մ�̠���@@�ᚼ�d"�>�zV��w.��d(�"J�5��۴���;��s��@{:���C3Q�ʶf��uYy�h�r�Lʱ��e�}}��{EvZ�Ҹ�$8���hʸ=Z� ��>̀�̀�d�D�S�����3Y����DsBx�1��/��
�p@��qބA�A3 :��Y�;و!!C���`�}i��N9��}8�֠��e�mm!3()�	٫��D��#2=dA�w��uۊ��c���<sUK��+{�
�m˻�p�<Drڙ��������G�x�Fb��d da�d)<��c�zt �zy��V�Y
�p@�#���z�Õ��d
gi�<�qŗ0�a�]�ȉDڷ�샳si�o�������}����g���7%Վ���9����/5�̿+bu6.h������;\���Nx�ֹ����ɝ�t�%��s�n5a|�AL�21�9sw�̏w���0<�reM]��꧖7-w�ݐg��w=�^����d9oa�Q�̠)������&n�,>�j�oKS��a��Kx}#���`>
zo���e0���M3���F��1ү��Mw���>���@�[r����`�m��`H�ګ������{�˛�a�]��sN��[�ǅ��h���
�!�q�0�Vo8*��̭w�^V����;���	hc��+�2XR���N̫�*Z&�����F�؛osbfn�KCҵ���U8���Ɉ������D��׏���۰}}ۺ�������ظ�rܶ���R�ʃsO�G�\;��x��(���u��l)՛���ǒ&|ܾ��\ʸ�=�Ys�h�UX�rfĽׁ��L"o/v�<fbpʷJH�2���0��ط�4�����0Yy�Ib��U�P�:e�Ǯ�:����/��y���a�Roy�1I٥�+\b��Ɨ��ptU��B�߳'���3񽴭�?U��8h��� kdkhgg*���{˺O/a�/f��TFH[[���s����l�ؽ-�ᒛ��Mj��%�,>����z
1�w4Z��@��) �5W83�g�f��yg��Gj!1�M�f�X}��9u$���[����8z/x+�N�#K�'�a>��z�>�3��i�z�wӢ��UE����J�X���w-���^��u�Y9BRGM�mŦ`s�2mP����mZVZD���s��������8��Z)G��ӓ�s�� ��A9ÁC3��A��yy�DG$G76���p@)�md�{g=�Y�)D��5�H��� u�E/j�Eq�b���Ƕ$+K9ɖ��,��	�Q�98DRty�'�I�ZDՑ�nS9�=��٣��m���9Gמ����g`�=�{��8��ďkS�z��tm�k\\$w�sۼ�.}����f��ə���sK&6q'IGw�{�=3���m�m��G �Fd���Nm��J)m�o�9!|����3E�9�h���"q�)�rfI�N ��7[���G�f�d���,��m�ٍ�:/{��9 �e����#�ӛh�ݥ�gekZl��%��������)�Ԃ�ҽ1${c;+�e�v@N�_	�<��<q��e�n4:�c�I�ֶ�f��M��.���U3nα��u�L�.8��]%���	i1�	�69��@�]v��v�jF.Թj�ƚ��j����̨F�#0F=h�LMn�kb�8;1�zSh����KK�ɜ6儛Q��K�y� �ݷ^#��3��[/Q�6ڬ�U�Mv���u��qyY�s�7#K�k��ᑵ鞬N���b����A�ֶ��[Wvy5Ț ���v4ѺZ�О9�< �|�����L�bm��<b�&{
j�z�Xe��Xݓ��h�[�&�v�5�<Q];>Z�Z�jP�"8�A{�J��]ު����kk�n��Ս��:�Wraz��čΟO"����t׌]��QMQ��n��ΌU�;��fA�r0��՚�LƸF�6����nfi�KW�L���#�]V�Sj$�ѵХm�&��6y;�l�[�:�BW��B�鮵�n�n�0�v��g�l]������EɁ�D7��d�*c0\e똇����"���-���x�mv��2vx�q�JHvq`
�2�!�6ݶ/�Ѥ��RV��ڼ��#�4��M�����p��/N�w)B8��PG���Q����%����%�-	���Kc@ԩ0e1�d�C���B��8�	�ڰ�f��v���t�����-�;G3�6'L��n�����˶�pA��׮����]���x��`^v�]4�Q����u �0�B+�����]p�b&��M۶㱔�5�+QE�������gf�
��(.5<�'t�,�>m��0��٥~.��؝�I�!��5�<r0ƹ��"��uQM�Na�v��<�{\�Y�9c���(�ۗ ��݆�(-N�.�����\n�^�fƵ�=e�Mn���)^v"���]n�A��
. �1������3i/��"���u��.J���k�v7��ݮ*�,�t��6����2��A���%�HaÙ��s�<�
z�0v��Kt��z����EH�ӹ�:sqj�im��ڴ%�v�4�k�q��m���=y�[s�m`���n"��Ƅb�f�a\�k�Fi@)nܣvf��/�ޑ��כ(����a�䢵��b�үu[��Y� T8�M32Ʋk�-sh�5첷G]eY�rXZ�0�.�ku֋�>�~���g\��3B�%���M����r�I�[{p7mf�$���}?�[����όōA8p�V�"�	g������&y �t�^��g���V���Z&e�&9e��Nsz����&`�9�gU�^��W��	�uusq����md
��ն�j�ue]Tϸ��Fj��� ���̄f!xG\tH��m�};�q����XQ����U��E��.�es#�)Vj�h�K6h}ܽ}�5����r;�kiQ��3���&GE�[��<���*�s,�1ˡʴfb�9ϙ=�F�]���:��rZ��mU\�p �<W�-��d"	Ç*k��I�o~����8�IF� 3J�(�zu�=�Bu�-An7��4�XHfZf^�>y���d#�̀����s8f�58 Y�67.��{���X�we��D̹�_Fc��g��ՠ����,C�J�ᴾ������~3�a>g��� t3���,�ջ���tw��[�E}g����^�9�1�V�����у���J>�r7�kiQ�����@D�!����YϪ�E�@3T{�sr��f �^eQ�oh75�J�;�}�|���n����Q�9�-�2��^dY��TU���#c@�!���;�n��� �Nc�{z"�^�s�y~ݟ	��Q=�[�V"8�/2��Cg.*��D���fbQ�F��m*30��t9B2f!wR��]���6���|�e]B[2�`Aл �Y��f�-���4�.��vЦγ�����;߃,�?��F^����t���z�2xSUY7q��p���`�g��%+0`iC.G� Q�v��9ހk+�K2�_ ��=�n������1���Dm}��0��.#�V�eǨ��@�b�^�3"uE�l�шL�y곢7ѝ���n�^�z[ɻp�7'g�����)�5(����1Q/�5c��r�)�v�o?�x�-�_�¯��}�����C�\v󭩣3O��x��B҆V,Z�e޸g�����c��i	��b���A
��V�s֢�ڪsQ����Ι��8��a��@�7�L�,s(�#ʙ�˺����P���Av��;���Me��z<��X�ʖ�7���{����u��[m��ۗ�=t�v�GP�L��6�ۜ��شep���껺�DSyWe��T�3*��y��`�����PSOy���uC�5H�����2Ջ֟�,f��{ztM߄�cu?/�U��_��z�7�G�Q����s#u�3ۚS�h���=��w�-s(�2�3(���[]�m*��8�'3��M:1�@����ٙe�̲�ʘs'4�U�_(Ϗ�,X�����¯�|{�#x���x��v�Nl�<�t��6�B&]ft��'87���75WZ���eo[/)���������.����YvA��[5/�xv�x��������𔡖�C�|w�ȿ<��̱b̴/�+^������8�� �{2<�Z|^أ>��\�V(#N��ު��9�ݶZ�r�VXSe�ږ%p�-�	����@D��Bf@U�q�9y�{�N�z㐸����bk"H����#�H̄�ڨ���{�:n
���o�$gD�]eG8|��h)�3�ݰ69��6+f�T�.P^>�Hn"Ӌ�Z~V�����8Qx��صI�J�{5�Gt #ّ@3!xL˳=Ǐ��g��r��#z���V����[���&���=��Q������c�y|�����ZVj�2���&nd��F6Φ1���T���� �l{2(���0��'Q���K�ͻ�ޕ�.�à�	��,2����E�oM�~��f̲ds���0�:��2Bٍ�`��6V=�l��0ڋ������{��?L8�Parj�&���.�#�#�k�hɛ����8��Zh�8��X���,f�jMjs�gV<Vqfr1=t��fW��7�t �����N�S�i�m�&�l���]�ؼ�������hR+2��6ŷ��|K��]��=��p��R��<��'���^8㙷-
f�7�m
Q�c����]��~���tGT��3M�\�F�wu���h����1��-�hSZ�uG�}�s=e�2��2ˎ����]�J��{5EBk;odG9U#*4��[���S2�ee/��^�O|�";F�
����w�o��N�z��Bf@@�3g���Ƶڙ���k�b{�,̲�ʗ2�;�pw�f��������w�̄B\�9��ȓww\z�K��z(���܏P�Ax�E��ۆ��[5@�8g�^��~����tE7�i�v.e#�,s"uLD����/u����_1N�Mׂ�}�s,�fY.fQ��]>�ou^���>��	OT�%	��3A2Z���dA��)[���m^��1%آ�OΖ^��іy����3"^�\,t���0&y	[
�/{n���A*/�b���`�iX0�f�}�Jo�Ig�{���k`~*`�����}�-����i�M���>��?bn�O�Z�Rb���$��L�S��ucs`���Ͼ�����x��2j�"s�%=�
�T{��A�G20ة�7�(�6��-8�Z~��ӝ>' g{�.@���y�~ߍU}Ϛ��#�Ṭ�feK��ّD\Vƀ����/�]/n�x��3"_]g�\<s�h)�3���;��uz�N�Tp��V��fYs2�2��#�8������]�[ۆ*�1Z�8H�A�A����[�1ӽ���>O_�}��w�P�6�8������݈�r�c�n�7!n^��5�Ľ�<����e�〼o!�	ӭ�}�����F=q�{vR����mI��^^!�"Kp�>!�DmL\u�T�H�E%��� ��B{N.ñ;�{0
��K�À�m��DlӠ@�^��;�H!����|r0F/CkO.�Al�5�9Pj�+WT�X;۝Tq�7<p�����r�F@���&�1�.ܨy�0m��73U���\��1����+S��`�}�V��|�Ay����%�|۹0�����܉��q��� [AV�7�)�5}&:0,�@>/�H#؎�e��g�x�t�-��ŖP6Г��;�ֺU��U��J�����ӷ����0�	�0�[jNwҟ�yzO��L8�;��"� k��j�m���ι�d{+����;-is���=�����O�>|�e�x��H"�Y�?}��%�"V�ǣ��_"T��0hF�k� �Y�n� ��@�|ݢ=���nC|�g3W�DS��t{{��� 2�Y4�fe�.�@�r$����t�6�H-� ��3}\*8��Es���r7a�7��g��y�@���/x�ԂmC,����U�deZ��^�6АE<�;�$�\�%l�q�t��<���U�Sz���cT��bb�(�p�xbs���C��^�cu��5T��ˊ�W��v×�#�1�P4Nc�p�{��E�@�mτ�[�k����q�O�:GRAe�7�I�7}%t`\Gx��) �h��m���=]ǧI��� �z$A*��M:/9���"V���k=d�WC������� �@@�7����-�B�r��{�a*�<$�Ӧ�vix�n��^E�^��� A-�$w�%�N��c�cH���}}�
y1=�I��ډ٘�A� ��q����4^D�P�o�H'�7E�������˅bD���w3Օ���iсq��) �h Cp��mȐ[�D���Y��C.r Shp9Ё�p���|6��ﰙ�O	�@DV����ϴ�/��Z�Cp� �פ6��!����EW�Gt�of"���t��vf;�{�/Cݑ �ȷ�mKSZ�ј���W�E�is����c��Tlx�=������}�{bs4��T!�8�:4#7�(ɛ��.��N>N�;{�7�ҳR������CZK���3.��Ջ�闺�׍�TE���u�>yJ��V�u���ބ!ݷ2uX^��܋�pЛF��X���o8�f��NR�V��B���*kYwn���K7=�VT�^��&��y�Y�m�� �gs\�8�����k����M[6kK�c�5���]�޷���p��i��R���Q��DM+��6��������a�Ҡ��]�Fe⹸wV�
��n��U��ejJ��f����M�w���m� ��
{!��C�n�J4����Eo\�.�Z�w���"1����q�p�����-�P�P`�'
�ة�-��w�c*x	� ,��m���3M{Z᪣���E�}zNr���b6�G	�4gz��=�����ډ٘��tAwdIn�%�ۙ��"�H��.�\t ����^5$7zv���C�n�HT�������t�ӸT5���ET |�W��X-�D6ױ�Ǌ-�r�b|V@A��\���VC��1�(��o�"�^E��!������4������3a�S3`��u[K[3C�di(�f�xYE�u�(���_�}{w��hn>!�"|ʈ���&&�N���f{c,e��'�8�/��H:�x�[�hYn ��P&c��kij�|�ܽU���ڹ��b�m؇n"���'a��I���ua��p����>����f��;vs��:$�X�k���e����u��� �܄���s-u{:2.#� ��> �A�8��UF`>���'�x�hIn<�,���k{p���f*jlf��(w|&0��A񾀁Y������Z��&�nĲj��@�����m	4s*"��B�\�:�=Ǐ�2�2�k^��[����m�>8� C,�m;˧QQ�X&�M8�o-N�{:2,� ����A�^�ۑ=7]2����L��f�Y�u�na*�@R�i��Ҷp��j��ptq\<�x�thx[����Vˉ��qE;�1��Ŕ�:�.9��6��6����)ۮ|�kķ�o5T�)F��1<��]���uy�E��
�ٜ���6�m �fOa�4�utz�dV�#�Z�@����1qv.a�����Z�7q�u�-��U�Әܔ��Se}��|��U��6^�&��n"�~3�NUl#��(��,,+uK��32�������Se�l���gt��.or�ol����k٪|2=7G��*�ܮ�2�
C}�W�3�ӓ��%y��!�ɺ��[m��+%=��4[q����.uG+��;v%�p��|��t޾�:շ8��^���#E�As�r�k�M�ݺ�pᕰ���.b7���)��NaT��xo�׮ɽ��V>>er�M[G��@��}�y���a߹�������g��6���Ӻ�2��9�s�_Si�m�g�����,=�'])zJyإ���O�U�C����ᜌ�94m��x�U���D(""��c.��n��!m7Lѻ/4N]KFx������ז_&��5�eA��)?8�\|�|��e�=2/,OZ>[W��	�;�]���[����³ٹr��=x��rj�s�pHNx�Pvw{Ք��3�Ҝ��6tfCҁ�0�6rܕf.\����;�k��=����fM��U}��m�V}����?��Je�#ǧx�{����Kw��~�wx��/�}<wγ��4�k޸��ۀ0����[���3Svi�k+�GG�:�n�~����j��8���G��K�]�{��$�z��#���6 �n cІ�:u�[�pF3�ƋuE57�B��K��\V��`C��#Y�����}Ǖ���k[�;t")�Y�Jf�I/:�y��Ͳ���/<9����n̛pg3���zm�l�kmdֻvۄ��wg	�9��۶����+6�����Rv��:�Zh��%��k�m&Y�,�)(���:s��Ye��#�mٵ����כ���dm���-2vkl9`�VY�b�2�4�l�m��l�t�)�a,��2�gSi�3���N��
3�"\��cM,>��t�Ќ�i�\�Dvڒ�{d����l쓧$��f[v;�l�Ӊ�l�2N���`���N �m�e������;��٭`�XOv��u�;7#�֘��e%y�^e��qkkml���,��/ow��6Yy��֣i�Y�2k��rDvT�(�/7�^�{Y�nIN#�����c�6�8H��D�4�T4�@�L�!�+��}�׎}�8iѺ����{6my��p(U]��rf�Cզ������p�f��.�V%��=*�-��R;�N�݀�A���<۹�6ÏQܷq���1�Q<��]��[���6�D잓����/.wEaQy͒�%�(Ml�s`�2w*k�c-v���F�%*R��q�Q��w��-�|�mO]��5����Voc�w���h7�m^�\�n�k�=�'��\3n�
�|+��; my��/��q��n�@��=͠�6׃oe�����UP�{�%�a���n�wSpi��=�����}��v�nT>{��������w��N5�Zs�_����u����Ou��l�m��oF�9=;�BױF���.&�c]�3��@�R�ɗ��k�v~ã�m��/���m��
��M2�{v�>n#E�[��ZJ�vG��h6h�aY�k˲8@F"DH�J�;<�kڇ�z�.� �I16���a��F�u�?���� Cm6�Ӊ�~�愢y�50�E�"��w�^��t�nh6׃b:9U���=�.�� ;`.�}����Ʀ.���=�n�g[��ȁ��.���m����M�vV.�z�'(l;�0��P��d��� 7��,�bw4NNKqm�y�4�b;ٌ%NSS���7%jڙ�V�:m��6כ}к�`�ͻb��廘�x�c���Le�w����Ǜh�*�ݙ��l���FD���]��UN?�s����Z�zN_Ts�7��S�@ ���{�u��$���}>��I�����|�V8�m��MIr����k�^s�Ce��lck�v^k�J�۵#����[u��6�f�K��Ў���:����ؖk4Il�� GKnL����>�=�:]�GP,�l��7�#l5�8{A5&ҡf���%cC��J��+f���dH����Z�yr���9�%&}�ێh���s�4�p��n	ے��x!����]p��`b�WOMS[�6�����m*��`M�譊�vp&���rV��6��v4�M�hُ��z���h7�OX/�F븄��Z�V5\M��k�RI/�ܽ��6כ{�$7R\>���u}��@orNV��BQղ�L.w��u7�'��l͠�	�hv��ށ��n�n0txU�w��㙭	����{w���m��M��8��Sɲ�by���������9��!K�)Wxv�t�]��h6��Ӑ����bxkǛ6���񄣫eb�]�n�u��x�<n��G��T�0
mU�W��u:����Sڌ����Q��K3�(CBW52`I=ޭ�9�����ר�3\K���e)��qI/+�M��7�z��5�C�Z��fx�Ev�W�c�(���v);{�hiW�^<�,�75��z�' n��+`6QR�Ԭ���6�&�X��_x��W����?X;�8�څ5�q3K��1���r��7\J��>^�mx6�f��}.��rU��	GV��0��^oW��i��pN�v�v��O\gk�o��	�2�k��^�d`f,:��^��y���M�7sNF����ʈ��#��5��3K��ٍ��q;��)���,)�"�fQ�Bf�=n/n�A�97X���X3L�V*������r��m
�Y%onhJ:�V)�r*O��w8fr�t�������5�э�Q�xG�n3�uE���u.�w�݆���e\M�φr��A���y�����-�Zr���F�C�)�J��Q+K��Y��d0�-�*E@�SnC7�S��xrwQ���kl�Ȼ=��UJ�uT����=��7gc��B��:���:�f4i��L'}���~��y�T�=��z�SS�;���]f8�j�v� {[^m��m�p��.�2�e���3���Q�0�]�p}�۰m �71$�b�[L�m��j:��mLʌq���I2�vZ�^`Yr�7f��]������y�^n�j'l����U�uMO^&>�4��yK�wSph���%y��^5	�xWnm(�[2���v��z��y[��/_rޏ�m���f��KdWt�l⇜�+�Q�0�]�w��^��^m�7���&��lDk�w[n'l΂���U�uMO{�����TRf�b�Y����u��3l)+s���g�cJ��lkh�-s��?C��EU|;�g{9�k��8S2�r'r�f+|n�wX>���{��y��k����@�����*36+�h8�㊎7�.f��<��6�x��������j���{��Y�E�X䞇23A�M\dm�g]��fD�d�a��m@�|��i�ۇ����ĺ�wJ���}V���VG����m�GU�[��:vEm4�R��b'l΂���K��MO{�6��<����^�NB�^m��6כvs�_;�<��8��{R�ap���M�m6�sW�6��f�^��n==p���9�ˤ�����Y�3h�{[B�M���m ڍyӝ!�kpB�L͂�i�S���O��6۶�7��R�Z&R|�3;hC����oul�r�ؘ�3K5F�x����k��_��ڪh\�=��sE{IR�5^؁��V�éM��ǳP��^���רz�Ɣ��g&R���Mڃ��]���^b7i�J����ɷ]G��,�!P����T�*�l.�ݝϐ�N�NT���ݍ4SX��I�л�NR���mݼZW��$�n.��S���!j��,�cVmAL3&K.a�Y*m�g\������mu��<��]=;	����j��6u�6����j��Z���ڊ����<��(�G�2!c�0]�d`M��K���`�dX}&e	32bLLL�'�/c��u��hUS�{��خB���¸��/^�W���A�����{��;�[�8��y�uft��;��v��݀��Vb�F��`����m�6�׽kHm���٦���{î1���n m��)o!+���A�U/ާ�+��T��]���&xc�SOۚ��^n<�A�an��U��	��oN��eDp�I��v��x�6��N�ZDܻT�$�%J��а���	kR�k������#'sEE�u,J"c��v!oPn m�U�o��]�D�
�S<g}ӛ��hW�r׆cM�m���a��"��(	�w�TQSQ�L%t�࡜>�h�wv,��b�K�/�[��f�Mv14m#Ԃ۝���8��yvk������2y�c۫� ��<q\�)K��û���b���RkS+'����mߛ޸�񊫬����NvTGYu��v�u�^��a�x��=��}�Ϡ6Ѫ�7�L.�"z�i���\\e5ݶzJ�];=O���͵��A�m���
��i��S��q[��g�\w!{�����6�����v�ȹ�)H���;WA(���W�X8��39ȶ����z�l�m��L	����^m��W\fv�l�Ș�a���n�Y�Ro�`��Ƽi��m���=ktM�#N�3�ޠ*+B�؈��"��i���\��y��2)_M{p��Ɂ�hz�Pnkͳ�w�y��s��eT���}K�+�)G�{Ԧ��S�����흗�+}Q��,����::ڿ^���r(��o�#ſ5_�tP��c��q�la�T���W���6כw}"ƺ���=>뷬�W\b�ӵ��g89�s}��ޘ�N`�T�W�k^nk���n5�g��ټ����z�4-�b'u���Zjg��^m��K����O^~c�/���hZ�]���h��ٖ�9Ձ�KX�Ff�[έ݀��������~�|�@]]�4)�j��6�T���7Z�?	�[���nۋ��#g���u�,s���q3�û�{���6�X����\"�Pn��tw��(���aU3���U�*{� ��vpkD��}{Bc&�4���ں�zhS�Շ�iF���{���ޫ�4nz�VV)��U@���c�'+4�Uz��7��L?l��/�jT
��aX�`B�H=���*���Zs��T���v�>�� �M��m������aد�F.�\�3��w9�&�w��/nǛk͹�Fw3��K��� ��9ب�kt�\�M]�g���g��ʌc� �W����Q�j�ݵ�ּ�6Х�W`�Q��d�V�S�\Wn	�2�vv���nm6���Ӆ>�]y
tz�n��E
��v�#�bxv�ڼ�r�ub�Ļ9x>�y��hc�&.��)Ã���֍�γ2�dû����k͵��&V-n3����=7�t��c�b�LL�X�n����[=��P�tk��m��V�zwf��H���gmR:�Wv�f��m�-'A[[Sy߯�z��܌���۬�uU�j��t��>�辐o>�;�ލ`���9'i�u�W�A��zX'p�r��S���Ey6��|,�(�կ��һ�Jw:�ڴ i����%D�цC2������]*tU���ɱl*۪��ȭ'�����E��ERg���8OO��J�t�����_� ���׵�
��^�0�21c��(^-�x�f�����U������o��mאW��Lf�1�.�s[�y�ML΋jDn��T�;]���(U�'C�3	�T�2}(��p!7tg�_�a7^y�U��+w"�O[�������vbf�7����N���f�,̙�gTT8}=����͍E����ۢ�-i{{�Ϯ�X���J#��d^�k^/�^K,�:^�0���w�i=|�W���;P�_��o�P�ޝ�=�ë��٠���-�8�����vs�*xhk�lqٹ�BA�9yx���շV��{��4_�<���3�o��|����Og(퇭E���2j�m>�γ_5{v�@��
���g�{����1�2u)�;���ol���ͭ�3�c�KO� w>�$5viEu�GŘA�͍P_�����'Y���Ƚ��������\���E�^��.�^��[����7�9](��=�O?j��75>�@yD�aG�
 ����v�N�=��b�^�]Xk���ޤ�w%�������8������4��9�ڽ�����j��������Z���p�3۸I��oԮv<���#=7O���4]9F�)����.�UeU(ƙB��e���6��\�{��ݕ�[[�$P�^��Q�r�쒎�%à�v�HvN�ã����m��˔QÎ�m݆v$�!	�I9��v�X��Pv��"�u�) ND������ȅ����:�ƶ�������kQ�����{[��}��Q=�'Sl��3��XS��:r:,��4�-�q˜��۳�"�њ\\�F�[]�t,-'p�҈rs���t��.A�V�[i9fmthr��C�L�.��QiY3'8�O����ls���(���F�d�wm�6��M��Ü�L�BN�ge�gsm7#-�`E�rIK2�m�}��Nm�\SkR;�{vt	��q	G�靮��+��R]�\Svlc�-�]�e�]���WF�DU]�ZЍ`&^�9wF�S�l�B�'R��d��.z�6�v�ו]TR����-���A��=P(Ca�n�6���9��h�V��1k����S��z@�y��ɸq�η�2	�n�v8�q�"��9�{r�b�6C��s�P]�We����U��Vv���c�c�^���*��c,V@���e�S	�l�����C�mRM�h&qŚ�T�u3�52��@��V�Sïf�n)X�׵��=zB3M����m��f�V�nD��+R�`�TЯ7h����7�U]�ӻn��O�nG �1k�!㸲�, `ѳ`ey�����vuT<q�G��ɍ��؎���/h��J����Ǵ���On�s4[`�nơ*˥�ƢB���!���׬���-��4$	F6��[��k�)^\3����	,�Jk�;�p����ѭ�n-�T��1;.}�Y�;z*�q�]u�M�.��x�R�B]z:Va��s�N����aI�LD���`m�\Iė[0m�O.���ǳ�yl;�j� �p��^T6�� �����W�[ḏ`vvg��Ç��k��v�)�Uv���A%�9��n���33s�^��mq��;〝�$.�u�B�l��b��6��V��Cg��u!���]zɵK�{]�����S�����=ъ��n�:8��c�j��}��tt�j���{kg�p�8��]ƹ��:�3�1e�%����c��:s�2�3�-z$`�� ��\�Xv�x��\���0��c��Z�'c�8rEL���uͲ6j�P�LhicEY��H���f1)X��h�k�9�\�e#u�|&;�fkms��Vƅ�!D�gS�b-d K�xT��)+3]�	
�-0˔F�3�"d"D����fA%�W�MX����[x�xA޽	����l��n�f��ܘ1�kj��C��Y�f��j*t,3���N��'�U�َ�uY�؄�Q"M#9�qK�!�Mg���)m���$�ĳ�Wp9��rIC�AA����ؽl��m� ���.��G��MZ�
�up�%�!��L�TŌ�6�G�()�l�K�vZ��*�%�e�5�ɀ��f+M�k�\ˮ��X���5c�X�-�X����^�TCC��^��a�:�"��:�0[��{�?w�ʑwC��.�J�5�\�J�-FQ��-��K��"Q�|����@6כ�	�0�γ2�dû��F���GX�t{���m�6ז��D�T-�3W����*;X옚؉���m ��B��d<���@�M[�m��o�(��6�(�)�"k{`f�R:�W��vjx6�m���=μ��q��1o���YR�dû����P�����S��Fu��n��^m��b0o0��3��r�&��vKV��U<'�m �M��\��Û�l@1��;.�c��i0]E,�1+�w&+�㷺Z/.�$��c� ��8m��ڛ��$��5{u'T�ځ$pL���e��y��k�n<*v��t���ɂ�f�ثݣw:ټ&����X�9��������X���yy��p�Цo�~%��̔���JnVϜ�{�=�;f-��y�Ծ!�� 7�y�ۇ�h�q��vgCV��{{���M�o�>���.-᫅lrX�b�Kbg�=����� �B���.�Ι��;��6�	��r'�6=���en�{8�vS��鲂���_rm�7��u#�S霢\tT���:p�/��ys�{�{ʹo7h��U��
�k� �
1�vM�3�=L��6�$g��u�^��A{=3u��Ld��������u�G.��ةRؙ�#I�틐j����u�6����x���T�5n4&�Ȟ����N��û����J����Yӡ� 7��m�֋9��ea���Y����nsj��7qEA�S�����e���.�O!j�D��=ʬj�nf�A�H��Jo��ҩ�7���L��A�{�:�,k.x�^�����n�<Ȭȟm5�q���]�.����b�Kbg��ފW��ώr䧒�կgG�h6��n�5�=U��n^Φg[p9���)S�����^n<�W[<��T�g��]M͈�x�.�v�{<7bۦt��<�i�o�aAf&�ɸ~��@6׃q]�b�v|5�=�6ą��x_҆ds��6ۦ�9Yl�sf��w��Tf��]�.�<������L��ckʹѹ�P���ȝ��y���m��WI�U��{sK��k��n�aJ���=٨7 6�m��I�����I�-��~�U�]�c�g	|4�{{�� ޓ:�D\��d[��Bn��bűV��ݪ��E�X��k�-�X�ev��jKUc���'p�3I���B"�t�/MV����A��m6�l�*�rb�s�`.���i<��=:�.��3=��כh��x�uwxd�ULAP�L�B1 ��sUNê2���l[G�3M1���)^��=�������m����-7����v&T��1���_]���[y���O,�2�F^b���K��u��9�cYs�Ϲ{\6��Ovee-�$�z�V�{�W�k���q��MmI�����˗�ji���mߛmל�<Uu�xL�d�=��k�wQ�ێ8����*{����դ8���@���vm���.���̨����S�g�e�>�m�ۼ��Z�v�&����<�5��u`Ej<%O��t�=u�U�.zE�p[�O��.7��]d��"*��BZ*���E�/^����g��ۈͳA�$���{q@s��v���]�u���U%�nff[F5�{t�>�:��$n��c��[����q�\�7��]�5D2f-�#`�B�]�G0��U�ؕ5k�-�z�V�v�f�X��dV�Ź��lgS����c0��	l���XaYu
MMH�3isv���������v5RU����e�i�Nnn.�n7k�9n�o��JB���L �Ҳ���!�`ciL�v�W���\���[�2d$Q��ƣ�;^Zn<�^�K�:f{k�
��R��q'��]W�֯=���ʹmUuIc�)ۮ2'u�T��s�}�q{y[*f{���W�s��*�l�r��5���^n�F�����W;y�Ѳ�c#C��\�C�ᶼ�@7]\.ə�����O����غ]��3���*��K�Pj[�t-ͷC[^�m��pgY��&�\��4�3c)�/k+eJ�������6�˾�	+����-j���.���&��n,�n�� �-�I�u,��)H$3�� frm��n;'c��'}��2.W{aWCwW)X΋^�8��m�� �N������;�]R��Nz"�;g�z��{�3Q9��:��"��(U��w��W�S:��.�K��~a0���i���{y��.�dGL��Tj��K�����m�Aݜ�5��-րnmx6�X���v�oVtug3��e-S�wr�����A��fatڈ)&3���{m���d����b�+�r ����&�if�tk���9�S5�[;ח���+n!�WuM��R�u@��s�����%���� +7�XB+��(i!n�I�n:n��O��9��IG[��9�v�����}��'���ּh]].���Y�������p��u�B����v�m��^n<5v[��g+j��­�@gD�Gb=��3���+�����x2�ҰS��������MǛ}��1ߦ����M�;��6�b���]k�Yߗ���I�����[O~Gg��-�=���B[���c��q��%�y��!���'fHԥ�\�=��ST�]����pws[�w�l7�ں�]�������LO{�����9;�o�v:� �i����6�v`���p5)�\UV&m�OQ*��f�{�y���ܐ�j�g\�$��0�A*�Q+�n����fb��F���q�am�WN�5*!J�tU��o�m��R��t��Tљ�e.�e�M��z7+�����k;���8/K������B��n�[ç�4V��C[^l_^��ʾ����m6�;qO���ӎ61ڼ�Vm��~��Y��ws386�y ���o����uڮ7K��K��
iؕ��P0#1<��Z�!��p��E~<�����7w����3N��±A|o��=q�������q�����n��,�����M�m�6�nz�״*ɝ���*�gk<^���1<=��v����Y1����ٝع�3ue԰�m*�0�1&�t�q�Z��&��`�B	3
��ؿS�n�n�qU�:z�s����ͥΘ�\]��uPƼ�M����9(���w5��t�t����N�Wu@��o^�P�:��F�"��V�35y���{tv���1�dN�dU�θ�7[�;�{^��y�۲��L��ښA6��y�;у��vp��\(�X����2W(����A��m�n��UF֬J�9K���A;�k����o&���p��s�@��w��n�u��)���7�{��v�^~�-'~��bZ�~�b`�SA�/�4	nzy��.��H��K�����e	����>�r�C]���Wg��g%�gv�]�W�C������hY��~���VM�C�m��*k���۾��u�2��r���Ս�0���,wc�Bl٪�Ya!nok&!4W3�e5����닌Ѱ [E�1дh���"ۢ$�L����zLh�#)������պ:���1��N�k���r�]�y�Lu��u+��)�����y��s,�����F�k<����ۈ��tұ�ZR�qF>���^�m���Ws����q����M�mm��P��7�8m���p���bb��1�k�S�;���Qk�K�������42J��u�C�� �A��n��coò��n;](�vw��m6׃p�^��p����M���K��{����cgW=g�h��T.��r�X�j�(�͏c�����m���혝����=wM���3kEK�����kͽtg��t����-=K�� ��!��ucq7�"�m���3���m���2dB�Q�^��A�n�m{l].��y1��Bc� ��,D�������ᶛy�7��k#\�Z�^���(ɉ}���w���^�$�tb�)4 ��0Ր����6��4u��í�s����m�7�Y,\�]�BQ[}��U��Ξz�=F��P��Ou��I�����g@m��^n��׶���]q�rj瘳v�Q��v��ۯ�n=�**L�1N�Ɔ�x6�غ\2'wc�8$UI�� s!'�\��*s
��C���yٝ]�f����Ǳ���sl�\7� �Sp�:�w%WN�$>��ck���5d4���7.���}�N2N�X�	H����P39y��n���uR��f��Q�]v�E��O*��F>^m���`�72WV�<✋]�9�۳K���;̛UQ��tci�d����N��;�m�^m�c�ƌLZ*J�x�y+��@���*,��>���77�l\���K�����챣}q��.r�٥��TF���a(c7�wl�ul-<���q:H3�;�M</�ʎ�q-�T���ۛ�B����s`�5��x�%x"�o8V���i��W��^���4� ��z��f�'C��3��S0#����s{��P�E���/[*���/��h�#ϊ%w�1�}	H_]�n�����C��u޶z���r��M���6��Ou��.�.�q�6:�(��$L5gb�[qBZ���5�>��<k|�>���oŌ���ި@��0R�\�PV:.���4'r%m;��8�Q�闱�Cg*
�ۊ��U���t�\w�O	�d�A��[���"�%_ws��K57��|$���<�d��k��>U���ǥ5�e�󻭛�:�z��o^:�X5l��C��	=�50��G2z����G�w�}<����{7�8�i�כ���f!����^.�fU��9 ͯ��۬n�G�[�z��4h���';"�a���F^�IӺ�qd<�Y�!3�3M�^���dE�ʇ�;;�T��3����$��)L�0��~��=Ʃ������Y�G{�Cro��=sry���l�JwF�u�m�ݿlķec��zx{�{X��3�V#j�Fo��5���t����d��8z� ���j���<o�.�+"j��ר��L'/w}v!<����[�8��b2����o�v>.�u5������~�4viA�E�Vٷeo�^�K[Z�GYbq�b�N����g~}��3��}�|���ó�f����d���6�rVYם�ÑB9J^ۣ��om��{�,DC��h$�,˼�p^k0J.[l����\�=�M���Z�����������f쳬�s�Đr]��I���E��X�+  �l�}��qO�޾�B�oz�^�n,�(�i��k�C�ڝ���{ZDH,���e�
	H[n.D���+:盾V�����؉��'<�Β۬�y�M�z{ܝ��ܜ=��>�I�Ob�'۵8���=+w��D���Ds�8':@�m�y�7���lͯ;Х K�n�V�ޯw�d�2ܗfVG#)\�oqƴ�o
��{����i����y������-�^n==|poQ��Tpʌ�������R�U��P�7���n�O����^��Ipź{YQTc�tch6�l	���
�>BŻ����]��A��b'����͌� ��|�'��0�T�EI݇��@g@�mUխ��=��sxT.۽B9t�V��(���mvǛh6�ő8;z��r�v�2�t��F�
�c�h��������l葛E�"׶��u��A�m��P���ja���{*��w���m��phdK�Wb'�t\��8�כk�ukz�;�y���\7� �;=�݆/{Pa��������"��1Mk��.m��D�<m5�B#���0�)�s8��2���Z7:�=�[v���l]<<��͡�]�;�j�G]�2Wv�����Լꖆ��=b�ܺ���0TD!�L���M͍�a4�bM�s���;�Olv�nd�gJg��k�� �C�ɥ�c����F&�W�j� Mr`M��ᶃm�	L��ð*�{sP�v��u=g��5�B�{{��jmȅƶ����!׉�y��h�-�ddM�V�vt���#A�Y1�Ϲ{��n�q��ig�\ܝ��)��<ۮ�2��v��s���U��1����:����=�<�^m�6۞�7Sx7b�I4�oH�z�U�����[�6�>��'vaKw�IC�.K�ϻ��Zj��3E���o��(|�+���4+͠[6�GF+�y���e{�����4�8�.D�K�w`hA��9�0�w�:������l����i�u��sNf#Z��`�vwm]4�G)	f��S����r�U�����S�Wi�`�'V�ei�+�zn��;v�g�>�u�����*ݨ���6%�5�Ƀ���ܣi�亝kcvbKã"����lcy�c%��a�ı�h�q.5.�����?����D�=0�����ocn����4>�U�Ѝ��ɧq?����{[w��V�`�W��1t4�8{�3��;]�}]r��M���^��'Mi(͔�</5Uq�]�;Mp��DЪ��m��'u���/FT�^����^�m��荊��½��������.� �Pn=��m��N
�ɯM�i����j�84�4�8ܺ��+x�m�����h�n��^m��^�ڋp��15�����g}3B��ށ/wt����?{w^)��"a�IZ  j��s���:90��%ۮn�0f��,Yj������@k����\�;�9�|meU����u���u_���m��^ߝ�)�z6�<j6����Cut�ȸ�1S�3��6��V2����j��-��+y�f�=7��sv�L���U"�L_
�,P�T��9^v�7��`z�{����$]9���-�m��({1{���.��5�6כ�6�"�U�Ko���Q	n��Z'}3B����i���m�qע=��`gP�'a�^m�Y��C��녕W
y� '0MV�p�����6�n<kͳ"�fQ�؈39��oF躾�I��9�����۠l)��-̓b2��@nD�y��/ϳt؋	\s�c.�]��Pq&<M`�h=i�����"�a��k���К�7�u�o���Lfzf�v�pm��(ֻV6v_�l��Ou�/�,��P�=廫����BUE��~��{h7�m6�o�ԃ�!��xyL�E�Λ�n�3�j��ѯ��dD��g9�$��3'�����{v3���N�D��`W��r^۰i���h�8h\o���&�ΐ����7vj�=\�u�7�{vh�oZ�[�ʮ,	�A�ڪ��>]'����{z6pc���ӳ��f��i��m���9�z�p¾�}]�5辴���B����u�Ͱ�.ܞ������$$�A�]�vG��ƅ�q+�׸�%�ZUn
Y)B�/��?z$���n�S��z�<���7X���ؓb%��\c�{����q� ��@C���3Yz~����:<����ů���������^ޏ|3vD�������G}~V�9ڧ�|����RA���5��ݿn1�dF�t5�UrYsp�
~�@��"A݄�����bO����>��G��D��H�n�^����ױ��| ���)| ��)"7�t��\4����M�F���y���<Wz��ݔխ�WF��o��r�0����Eױ,��v� ʝ7,Ee��Z"e���/���)�#v=��X �wdI݃'Z����}$��-�Zί����(�|��H>=�/FnȒ7vg��>��;{1uv�@�)��f9��*;<�n���a.Z��̼*�a:в������zo������)!��n���y��Zw�5�U�i|�
�`�/n-^�� ��}�`wv@��}����w�!vc����$;�g�}�/]}���33���|�/|{@�Ax��Y���lۯ��P�b|	��$g@@��A��ȟ�@�7vF/�6+��1S�����4�7
b����� �#wdO��A��A���0k��]��^}��ݪ���U�G�:ݏ���^M��S��|��?V��E���9W��yǐǲ$��$��7vD���s7
I5=>�W��<���r2��-�5�_���$���'ۺ�L#{����_��;/2g+r��F�5�ܺ��-V�E��4;�sF���{�T�+��"x^��������m�3����DAR�k�#�oE�A�b@�p��t�,hh�MWe���z ��N-V�Sq�]�	��`g3%�LJ��y�E��*���d��f�����ۮ&e@9�S��2�J:��������g��&f0��*�G;��Ҽ���]���6��N��8��s7\rk���mRd3QR�m�:�6g2�QڷM0G�����.`KQ�s�.C[�Zƃ�h�����=���=�v�]�(��1�E&Aut�=a;���c��/Z�X���X���4'���C�Ղ;�"�Ȋ_a��]o��f+���D�Ͼ��[�(kP���������� �wuI��S�W6sF��]�	}��#���k�9+�p�)�����H;�.��1���<��G۲${�@�7vD�7vD����]�s��
��Z�j��_���`�|�W���) � ��H;����G�U����{Gf��x�;:D�{�}��&�Z�����-L�|_�	��@���Κ����>����o� wuO�'wW�n����_i���k.ih����k���m����^+��O�w�BA��}�wd}5�l�m3��%>J�&��)4�XĀg�n&���nѐ�\�u�³4��d��F�� A���ٟ��������_��C`�|�W�2�*4p�����\A�#��|A;����>;���D���om[)vĳBr����͍�c}��.�6�T��4,��v��Awz>Y�'u��e�w"Q�L0q=�Y<����G��}"E����}���6�b����� C�BH�ѵ<(��3�r�����^��wT�N����v��X��.�+������)� A��<�D����"@#wfAڜ�Q<7�*;�0A��G}�>݀����Y���P1�U�_=�)">�}Y��G^��S�[G�g>� A��RF���� ���$���~��T�o�r��}��R�����B�n�#wf|F����w����7z�Z1����<�ms�L�uF-օ�v�qQ��tN/� ���H�A�R�uMg�/�8�����\/����߱s���XQ�JA�b�D6АCiq���}ݕS,a}>��*���|2���`�����'����A�����KcOՊ@#�Hu�wv}���OƱ	8�sf��k��ۣe���½ץ�q��5���XՋ[�����?#���s�Ҥ�U�Phc��H]NC�7�2Ԩ���H>?}���$��Ӻ�;����/��kݷ��X����$��k>i5�j����9s��w�H"�ڠI]c<s!x������n�ݑ$n��^���|a3�Ϡw��<��N}�[���9_x�w��ܽ���>;��\�]�>TF���#[ ���b��|-�Ey�)9N�sv8WF��r�h��9�z|~s|��b>��$�Dn�}�>�k�ˏ��qJ+�j��A}F�%��?F�7hH#{W�n��� ���ϛ{����B�n�6~�RA���W�&��_U8��.b~0>;� '�H��	�	�����D��t�A=�"��ws��Ẅ`٫��Wr/�b�ܟ�N>�i|�W�r�� �wuH#u+Sy(ӱs6���$4��BA�-ݑa��qw�q�츥��� ��Ј�φ}5��q���L��e}p�蛊ۤ9zs�fX�x�"G]��_m�vC���u^Z�Ok&�7ܷ⨛fj�D]�12�b#����Nfώ�����H#u��n`�Liܕ9�ӕ�j����9s�� A��>��$�� �ݑ���f>^b���{�T�+Wk ch���r�)��6�+��{;�U�� �Q"Ѹ��<~���"H������>����ָ6�u+�:��iw���k�݀���H �^ݰ�����	�����~����.�}���Y�?eŨ�����	��^ ��ȐF��7��:�A�(���> ��T�wW�uY�M�����r�1;�s�1<&~����'�vn쁻�$*��A%�����_�@�~^݁�M_G�=�T}�&�b-|�W� ���$wW� �°�������>#u/n�#wdO��9�C�v�t��ᏲZ߫�층�7zA�?}��dI�>�n��������W��_R�������cieh�'pI�>6FN��ج3�	k��PnS7\����k�G=����U�Oݪ��B^�(��k�_Q�7���ܵ<���b-�#�f�0��]�O{z? ��q�xu��f3|���[�G|�ܹ�r��C}�d]��t���6��=�>���m�W������x�lv�a÷[����l�ڏqK�%���[�>��ܒ��O٤���~�I��.m�/�B�D<^��r��f��<��1���=T��G����{�<.:��[c��<�o����c����z\���V�=<��x��W{���zNd5G���Y������<œ���ʒ��������2k����s�ŮM^����1���s�.��W���w�^?Q�@�$��_gJ������$�܅�묺3Z���u�@�~�{~^�q��79=�L�4��<'3�{�O� t<}�(֤FR�Ǥ�+1�/x�ӏ���vL|�{��P�DH�6.�3ue�7Q���(�oe�L���-Z�I�>���@��nQ���!�����5X���Y;-�����Di�6yǆg�)�8��$�R�`����fQɠ�L���>���C(z��1�$����9���,�H���!�p���zi���k�a��~�Y1`͕h�*tE���ؽ�:���=�i���8o.�^oQ��8ow����V�m��������C�_ E�T�����	GzX��'.����-����Wg%�*�8�6 �%~}h��柅�����JRw�p^ZW�{5g t�;�w���[l�)Ӗݡ�qrcjn-%���n�כ4r�G�"��NF֑��y�=����n�;=�9���	̭��{np��i�s<��i&�^���X�AfJr��б�yzb�j����=�"R���<m[���my�-<+C��k��\�>��;S�-q�I2�<�,���
N c���.{^�m��^�����GG/Lvm��F��[�E����՞k�NOkQq�9��KoZ
Ie�i�
��Z/2��-��YKia.��^���9nJ&֙��ټ�y�f�{o�J�G6��헶���/E������|�З���9�w�ݞ_2(M�IHm{�S{���I�UC���*�G�����֊Ck�#��?w}���v�#���U(�l�Z��0�v�pS�h�[�3�t���A��J��6�,�����ih��l�#�����YJ�8�uճ�6�㞞�b�O8ݩ��I^N�y��A�����b��5��-�*��ڎ[xN�U*�;I�XK�F��E��+e1�6BkZ�Ӎ��:�v��mv�A* �����y�J�x\�� �]��.��Խc���;���k[4-� �IT��WY�q�;ե@p�84g	����\�k,��.�h�do4�k�PeiQ-��%t�K��]1��9�8Zm�/�n`:��u�L�����on be���X��j�Ѭ(���බ�8��{V�]�xz�9�՚e���^���� 8�Y�6ɳ���9ע�=#�k6��{:W�=�-B��i,�,��W]��i�PW6;.q
�!�3]�v)݋c�Gm�2�`a6x&#rBS���r8\S� �*5S7g��v��
��*pJ�A�YWXivz���di+3[U�X6�/@q��n�#q�{j��� �n{bY���۠�R�n&R���9�ɪ���f�]��p��6�L���[����
A6yGL�bֳF�ƺf��K��nXvf6���7,�e]c�jp�6��qhέ�#㓦i�n���'e3�瓖��96��ڳ�:��9��WCHX��zK��7R��)J�e�՛D�ôj�k�,�g8����Q]k�\��N.�&p��#ܝ�́q�ݹ.��^q�&wU5�t�/��"�h�D<���[��ۍi�>����*�.���V&Xiv�������j�8]H!jiol���^"��
c��Ş�]��ƫ��.�[�\������d5���p��i�����yv
����S��dqv�J�k<X9c�F��G��G[�vt�u�{]v3�c6�6�۞�K=�U����B��WXI�]Wk.n[o�.�g�����\����Ņto+���fP����k�s�n��l^�=��5ړO���H��"�XMUⳇVn+c0���rn���tȰ�L�u6�ۜ\%Rٶ%xd&�*��54l�x���70�!�a��۷m�(��i�k�i��Jy�%��]�;p8C��:ysQ�J��rv|[2�oU�z'>46|TF�m��h��)���a�\biv0�E�������^�. �W�3s]n6nU.�����r]q����3�U��5��<A;ڤ����R'wT���r��_]?��e�L��t�;������? 3>A��<�����$�Dd�؋�PYG糭p�3�z{���ҳ���lɫ،_:���'�� �܂;�����}���u_ٵ�VԂ/�w���Ȑwc�n쎩�����;��붗eŨ�����ﾅ���n�>>�A wuO���5����ڞ^�h ^�N�y���ھ�E�b��R� @;�!>!���'+����3�I����@��B|F�Ԏ�Z�w�6/cGz������u��d��F/�J���|��܂;��n�Vy�!�G�Ws�TAI������m#��d�R͓���V�՜��q`���~	���܆�@��ݑa��qw�[K���WW􋪏���@�Q� ���#ϧ�u����*��'�8�rn~kf\?�0ޏ7��=�<��<dZ}��9=�����������GՇ���?�ob��F��t�OVdѿ�����=SW�&�>��m�F�����	���D������+�{���}���_�;� n�O��Ci���*��r���ٓ�v29ԯ��w�A��#��H ����G\��ۭ��_j���"o�1�K]����.-E|_�A �� D3��{}���:R��#��㺂;���� wuFЍ���~ʧ7N g	=?)������y�Yu	Q缇��;�D��Dn��=.�����_|�p�6 \�
:��	��B�E�U5�uh!sIpE\�y�日��s?y������ﾞ����ٓX��ԯ�џug۰�}k�#m~���#u N�$m���pyvѾ=p�{�H��d�����ˋQW�~��7�����]=ӝ��ݩ ��^�����$���߇�$)��&�K���^��~G���'�B�'�{�(2������D�ge�i��V�37"h�s��l�[F��u��)o%k͸3�Q��� ��!> ��'v�>���7vD����6�����H�=>;�M�};_=��fj0F��| �|�������M_۫VW
���	ϹI����O�;�"|wb'����S#�9;6ܵ�}g�qj/�j����"�'�n�ψ�B+[���g��}Z��Y��m[6�f�����.z��4.q��ܶ��*�����~�-��T�~����Sw��>�Y�W�.��+��%�}�_ӏ�(��w���"|F�nő��Z�z�W��;PWW��k���uM�~j��>��z{�GwV���w��o�i}�1�	�y	��$����AM�o�&�����g�Ũ����A�C{"|F�O����":pC�e�v��=�>�^���;��]�	��n3쯢]G�W�߾BAw8���w����M���2J�@ɲ�D�r������F�����D.wo��^�[�?�_���\7�C��H���r(,P�-���#��� �� ����ȐC�펅�h�*~=�.�^��{5�u�:���~j��w�^�������-`�7���D�����/+sM��:����U�.;gA)�B��7^6L�	�� N� $f��v,F�ȑb�W�����_a�W?
W��_�&0�gF���/~� ���Ӻ�;��'^�"�.q���L*U����5X�K��7y��~{q�:��˨�J���A��wc`�\L����:�dH^����Bn�#wW�n�]�o3�"GƷ�˚��ժi���| ��/Or�wT�A��>#ux!��3�T�[��x�����D��@��B}b������|�.�g�Y_	��{3�0�p���1���;r@�oG�u_��uO�;� wu���"5����#���3�Ng:��̨�J�{~�=�"A݄>�9W�b]<�`L���#�b�s12o����N��˄*��9���w��Z�g	4�+x+�g2 p5��tR��z���rl���0i'7V��(�{�3�q��t�VU��8�{v닭��A�j�vS#6�H%c.,L�[F�����;�V��N:ڻf3;n:��.u��!�y
ϓcZkso5�W�+=v��/6-���z^,��k�y������m]8�"B:݅4{g���k3`�s3��q+�Q��PN��I+aח��ni7�bjIs.��h�Sk������Itn���OX�E9���w`K�����"@p[!H�O��	ۄA��$���vW��5�u��K�cp�կ��÷|���|A�Ax��$wuO��H���3#�3p�j��:3�;��l��c�_?��fF]��*���B���>#wb��y�~h/ߔ��[�{v=��A�������'�3�3��1�ҖeG
_y��A��݄A��Ȓ7vD���>v�ۘ�_�"A�H��U_����>��d����_A|�[{[��S�7,�w�N}����R�H��IwdI݆��|��S{��Å7��Q��#*�~Y���мCz�������O�+���\O�0}�"�{�\{h_Q=j��S�f�G:���y7_����F#�������@^;��	��7x;&n�ϝ�̘�R�!�ov~��;�(��� �ݑ �ݙ�%q��27���F��{�Kow^nF�X�R,�������Ҩ��r�����Rf\Ѥ��V6@�����ʇ���f���Y��N����3�w��[���*���m��Fmb1�~j���Gr��`�����m�U�!�����vn����ML�&������nde\�«>?}C{"A�"|F��wT���YD��'뽝Y���<�z|��^���ѕ�P�,ɏ�/� C!�|�O ��7�$7vd��Ỳ$�ݪ�H�
^(�����շ����"����{���$w@@�� ���픧�������%���I:4h���؉6����^}\pY��.x��^M�����+�K�x|{��H�wa��M�?
��}Q^FU��*��#����ȧk��c#<Eo!>#�dO��A��A�S�:n�ݟb��W־W��?�����_e�̘�K��~�	wt�v(\��2l�>����;��#wdH#wdO��P�̜�W��}�+�l���M\�R�+��'���p.�5z�5He80�tt�;,��]�L��Lj�W*�C���Cn�j����y��U�EN{�ݶkNδ�l�կ�%���^��d�RF��[�>7�#�؜C�� ��ۺ�ݓ�ܾ�^FU��+/���z2H��{n�l_p�C�>���VA;���7W�u:�W��,~m,��W�ۣ*���dd|*`|��A��wax��B��wqK��\��!�������uu�v�q9�Ok�<�L��*�.�/����߃,����g�ߴ��5��w��M�ʥ�Z��gMy��)�ի�ܽ`��7R�BA��������9yx����Nl A��'�_=�}S����V_�A�@odO��٤d�|�Ǐy}���O��R#uwuzN��	k�_^�Q�9��u{@����T��oH�wa A�"H����o�����nȐFwH�����v��\_ɹ٩_9��� ��^zng�3/7�S;ދ����M�p���ǧ{����=�3�޺RgU��KE���P��X�K���ё	�eD��6.F��~תA�ϔ�7W�>;���}��'�vn�3�<>���'�7��T�}�n�~Y�O�B ��� ��^��)�	���N�d���ff�1-ui6")�F��ً��Y�����cQ�f������WA��S�A�A�R�꛼�}[����~����,󰯥oA�|~��[���/�ݑ$n��� C��H@��f�F��|,�9��
�>�v�~����T��Z����^ށ`�S[�v/�&}�Q��{�a{��$���'�v �쎹���m����{��Ю�~Y�~��� ��^���;��26o�Tn�����#��H'wTݜ����_�O��#�s���	#y�Rd$�~�_1��G��􁻹��Dn�wH���&2����{� �|��m_A���3�1�U�3�|;�ۺ��㻪���m^���.g�c.����[���x�S�����x���[��A\Ը��3`��ͭE^��;{5�o3����vo=����d�hE���e{UWG#�"cM[�<.�!��֪v<ESY��cv�XƣX���qb�k��e�	��GV«�9����\�؆ƍX��ɢL>��Z蝹��d��v�v��p]b�#u3�!�g�����A��u�I���������Sgg]g�C��$s�W.l���
�Q"��t���*�c��%��-�.��X	p�M�����<
<,�%�<�#\�s��>:y�k��C�[��pC��� O_! ���;���ݑ6,p��G�Q����s�Ϥ^��O�*}�H�1�>�n��� ��R "g�����ظ�{�M��}OMU�D�N2>?	|����D��.����V��[� ��BA݄Aײ$�����
�o'�~�"�.���͝����| �����R�uI��%�.� +Z�v�n�,p��c����-\�&���G�����Sj��_���wuH>�� F��K;�w3����#b��zjo��������_|��wH�������v����{���=7�	J�-�r�i��-�/i��h��{)ij�[n�����B�ub9�s�5�Uw꺎��NTu�p}��T����."�^� �wuI��wu	"�gnU.���2�"1b%�NEQ���aY�h�v��f�SND�vN�����輁��~�jx!t��B�qCu�Ŝ��������p�;�H�c�}�>����6�xMg�	�����F�������嚕��e ����=ڤ�������Զ�P.	�6�����lP�g#�s��!$� ����ȟ���Um�u��|A�H�Gv�O��
���v����u;Se�����"p�N��F6����N�)#u N� ��BA݈�,����ک|~yR'�-������Le��V|$��#wdI� O�```����z/s-`K�棃��Vk�@�tAqV�i��������EB�BLG~�- �|����{wU�	��4/��Z؛�H����\��?�Y�U���� ��ϤI��^n��7vD��>��ա�����ݳ���S��:���S�1�v� �_�)����X�o�r~�k�� Ow! ��ݟnǬn����Nr8���9���8�[��W]�!�o���-ك/���>�[�d�~���Q�?{6y���U.��f����b����f��>QJ�W��	����NLf�;S�J�����6j�BTj��tݙ0�m�|Tx'`g���3܃o����f{,��0d����:�\p��̿E�O��V���bm�4fF�V̙4��S��R6�n�{cv��x�x�2��w=[q���˥n��9o�E3`Y��>�����pР�Ǔ�2�oj�N�
���of)����-�;w٧��ӗ�n�{b�f�4b��ئ�~\=�,�����0��u�n�űQ6�XE��z�^���V��ɩ�)R��=��{[�d<�����I�]K~w���Ű �=�ww�s��H ���gw��^z��7����ݘ:���U�ttɭ����Q;�`Z�S��;��F�6��X�B��j~���J�?��}��l�����w,���^G{O�t5%�7|��qJii���`��N�����U�R�cM���z^Ճ7v��M&<�?id�m�!fS�`�P��}���������ލ�^r�3sn&3^R����:A��'KfDG��pGSdʹ2�"���>:�4��Z�yx���zSf�x���1��e~n'��g��.�wy�cX[�Tx�hd�;���OJ:��R��B#�_��d���f�����^:��of�n�Ʌ�R����I����1?}�9��=t0��~�2��\nKw,���nC��q�@��u��Vg��VW�HԴ,Am�1A�:�%+Ҭ��9�<�G�<�w�q!.3vמ���q}�e���ĥ'�z�ۤ�{VW�^y׽ڎA�{F�k�y�N2�;����6���g��Ck^�� ��������bv�/4�;�i�=�^@tQ2��t���"_m�Im�tGwڵ��9/�Zt�ڲ𣓣y���6��7'Ͻ�Ok8��C�"Dr���������Ҏu��z�Y���Ӭ/m�����ݝ|�:m�_m���$�>b�Ͻ�&�Jq
�[W�h�f�ٯzk[Y$͔}��^�;۷}��+ӭ;k�E�����y��&h+�'�;��&9v졙��}o{m���Vr�H��7��!$����ȷBp��ݲ̌{on���������b���'�y�e����0�޾
��H'��Ȓ7v@���;���SWt'b�'+u?F��^�>��>�x>Ϧ���������{7��u�%�V3��>�^.�x��ݲ$�ݑ ��^ �ݑ>#wb�VgO��������n������jc�_x�����ywuH ����;f�~A��?���l��b�3q[�k�J�u��>n��H�5tDsm�ľO�ǽ{�ɧ��onő��H�c�v������5�����!cnw}A�"|��g�uwuH ���H���zR�΍��|sqI��"����a��U���\����I܄�غ�]F:aޑ>#/�H'�=��Y�"|wP}&������w���]��-�ژ�_x�_�/o@�����n�>�ԈϨ90�Ԁ�����@���&Ŏ�o���Y?��A���D}5�:�N�q	G��;��d9�����ʓu]�/����"m����8��1/Z�2�im��x����陑E�&�\>"�g�ﾀ���� ��݀��-��Jq X�t>���|v7>�zn�U���\���! w�D��[�# vг��j`���I�v�*S����.ݹMC;�CA�Wfw�A�h���~~��<�~� �ݟO��e���u��-���'Ge��������x� ^��|wuO��A㻨O�ywÝ!������Fw!b�	����<0Ud���� ���"ײ$��ڋ���(I]��^�AW�H ��)7P@��A���(K������-��������|��o�"A݅�7u	#wdH��Z��z���[b�~^��_am}w�jbt}�k�/n����-��I���BH>���}���VQ(��X�oCݹ>�>ޏ�_�����EO�	��@��dH#wW�ۨ@������byuX���o�<�dE�vK�y�I�����F&k�!(���4�d�9ĝU��$/}�����_c�o�%�O�����{�|�E��6͘�bԧ��v�WE;]�	�nӆϳq�1r�S[��g�i0n�$a�Վ���h,h(�����;]<��8[v���������<�cplt���̶��){Wd;s�3U���)���)A�wB�Fb$FiJm7R2,Ok���[E���c�z�X饰7#�/,�8Һ��6�5kQ�S�ůn;[[�]��>y����Wa�I�I��9���7��=un�L<�S�٤�������_?j��W�u_�'wT�^drϪت�O���§�����>���nw�L4>�܄���;�"|F�̂wax����E�]3+3@�����>�k��w�Z3:>wK����|A�r��왯��O�=o�^��{w��n�;��;�#sa�36��8M��#꿄���D��?}Z�D���'�u�� �{x��7"z�oJdm{{��n�^d|�����3�qQ��|��Le�n��U���8���� �ݑ>݄ۻ"|F���\Q�w�9 ������3���Ώ�R������ wuI�G:q���3|2�`@1� ��/,6.��+�<��L��c�g#ksל<�>����^� �����X�ۻ"E�ٱ����V
��%?xH�f�n~Q�dݛ�w� 7������'ۺ����'��s�O���Ə{W�P����cH�X=_.������O{7u��έ�[=�^ćo��lt�L;�{�{i�fr��N��A8�M�Du�P6��p�.*>?�|�����ϣ��Ücr\�}�L�w���H#wf|}��=Ԭ���}XO�W.�+�Ѭ)��K��) ��;���wu{v���[�NU���$������wdM����5}H��૟�)�H'��Mow���(�Ͼ�>�3�>�;��|wuIn����G�/�BH����������ң��c�S�@���I~��[�#�{��cXd`%7@�[q����3Z�(/l�[X���]<�i�6�J��~�O�@l�#wg�O���ُ�u�7�p�*gG:��T��~����*��A��> �wuH#v;����N�6Ns� ���۽"l_��٫��G�']|"g�����#wc��鯊���\��k�R|��Iu� �����!��N�RP����:	��7�Aq��7jw���>L����v�����S���+&Lj�7�+�{���B���L4�l-c�]<��<w{��q:�7' KM��.&>0>/7�B|wax��������ȭ�x���"��I�� n�����Q���iS:9�/����H�̭ٿ���`1�� ��� ���� ��;�"N�Led���0_��dH�}��/���
��D��A���D7�$�ݙ��NV��V�]3_#�K�����.�z-�9��t[G+ON��6?֧��)�"LG����H/���}��}w�d��!���q1��!1%wϋ�iAnO��ۺ����$wa{�O�8����(�CϦ|C����gj>�|1�S��T���>#�=��>�Q��;q�_vu�G��u*A���! ��ݑ �ǖ�ȍ�� ?��;�Z��u���3���[�F�ϧ۰�� q�]}�
��7�ϯ>^��~)�Wy�h��LG���
��'~�	o���������}
h�ʏ��
�S0�_����Sw�Q�]�Nɝ����R��P�{���9�s�sy��7�uh�yS�����Cw����vݑ$n�_A��t*����|�vt��3�2�t|��>� �;��uY�T�^�����&R"B1*P\�el���1�Ջz�qKZM@��HmE[o$>���M}�I~��yݑ X��1ٴ~C��3u����"�ڂ�a>���D���#w�|F��� ����|�Գ�l�A��^5�O� ���%c�~zb>.&8T�'~�	 �t� ��U[�'~��q+����I�Ȑ|�@���$��>>�C��\ɧ;����f�f}�U:>uK�}��H;�ۺ�A����,(iq�W�
 ���D��wdO�_|#�h����u�������ì�[�d�>#��O����A;�����wU�n,�|�)1�OF�P>�1�U�@���!> ����ذA��H�������w���
�ч�<����籟-(��ãa��fi*ҟ��j����܃�n9����ܶ��'7͊��sU��@�k�S1nZ�Zwn�+��k�����aB�Ȅ�;q��ds�`�̽Xh���R�;%%ի6����@���^M5�N��I0�v9��"]�M2W�T�Q�v�-�7c{IF�D�[�R�-8�9�J>z�͸���wX�JԱ�xy5���5����Ɠ_����k��ACE��cAGXZ���4�+���/��ιm����:���zi���Vݻ& sIvIx�AHJ'�+P�{!x�� 7u{=��ϳ>�f�f}
�G��|N|�~��+�����Ё�mI��-�D;�5l}[�k���5���7>���.U�����Ё��#w�-YSi�F��@��) ���n ���f_�vA�2�]�;��@�3
�� ����vD��� �@��ý�����yE����6�^�j��VtQ��c����+��鿼�s��i��C�s>RCip�mϛ�v'vEs菥���	���Bp�r��D��ﾄ<A�/ۑ>-��ߢL�?�_��~���\�C�%a�N�Y�'�x�OI7��Sk��-[�H�	kql>�'�{�����0�����DGW��Ӱ�}fc�O�
�߻w�uvl	�>�^� �������c��Ze�s�g����dFJU�e�][?^��<<�g���:-=�A�EU���]��1ft���ZxDe�D���}���,X]|>�]3��+�ѧk�>¾t}S ^j�۫��q%�`��A�#�ۑ ��B`��+��s�^��%��pS?zA�s�@������P"w���l��k�+��\<�Gz ������Dv|>�'�Y��T��=�*e��dV�c 4� A�4!�"A-����Ƙ���C������b��.tuL|A���n��n�m/�Q�ТqS_tQf	����!���^l�L��VG!ƻ���Z�u�A�j�N�)���b��-7��hyʸ��Y~����ϯ�B��K���J�����Ƞ��H#�A����/�|mI��ԬF\�� ��9P�'�T�舋��I�G�f>? ��� AvD��s�5$ء�+GD[w>n�6�!�"|[A��_w@����X�-�_�a���r�i�}4�w��,);��ZS���{���b�w�M���؍
{/�:�-�n_�K͚��$�|-�bY%fpZ$���>���A�-ǐ-�$6����ػ�Uy�ḮA�h*������]D������O��C��5٧��O�X���-�͵> ���n:��ܮ���~t������;$}fc�O�@�{� �Ȑ[�A�.u=�?L���Y�������@�wF�3c�l�jwT�RB����Kd��?O��;JlysAۙ��������G>fxI��1�#o�{�߶��Ƃ�{���^n��-�@��)bG�C������;PS_|��}%]�W
��A �Ј>�A۫��"~��������#�������� �mfP�05	�Z�����ZK�>�����}��q~ ��^!�2����?W_C�����_gډu����'GT��������{�~ԡ���o�'~ۼ���i܋7A��욟������4�v����L��^�8��B��{��ʜ�K3Q�r�:�����RCp-�D܉�nJ��('(.�{2��W=�N��3�A��Ds��m�7���F^��m����¬t����u���.�X���^3�\6�,���.�Ns�P���,�������<Ax�<jo�����i=D}fc�S��G��hg
�3�o-��}>�!��b|� Cx+8D��K�=dT�F���^n���m}�\�$��\|A�� ��������NY��ի�p,��ۑ%�D6���F#3w+�칛��_V�Ժ��\���#����|Ch [�ʟLfr����x�+@��j}{�"+~�l��G�j>0>�/��#G��Ɯf������m�����m�o��Ϸ)LD����G������sż=W�G�ۚ���2�ff_�� ���rO��O�HI*@�BI�d$��� ���RO� @!$��	'�$$�� @!$�$�� �T� ��p� ���� ��O�@�BI�I?�	'�� �d� ����(+$�k9p�� F;�B,�����W���&��>�N     �        �     � ��J(T���*��AQUPT���T�P(� $�HPT�J�IR�IQQJ�(AEI$���JH� ���	�*R���x>�(�eFأfS����V��S@\��@�� ��O@=�6F�u��Jhѐo�@ �z���� t� �] � uC�T��������c�ˋ�C�Ft��V�Ωn��� �tP {���tw<G������Ό�A��x���A�ѩ@(QΤ �$���P��W����lj���w=U��M�:�W]�)�4�kPA(�J@���}Α6�Gr���zrć�jn�N��W`´4�A�l�TDs�QQ�P�P���ى�Ee�F�Q7Q3�[�B��}��F��*��;���:)�Α"����	M���D�UH�C��d5&�*�b�ͨS �E��l�*֥0(	 z�$����� ��UKa��V���hS:��J�����(֨S�Gu#B��D��U8w��#�grG�12h����4�65-�^��      ����Jz�b0F	��LɀCS�2��Hi�0    ��U&�II 0� #   �ȩP��@  �h�  ���(�$��&��a2yM&F�F�0��$��H�i�&�L�ɣi�&z����{���Q�>:Όh���s�(� ^��6�� =a��
� b*��aO��U} '���m���������?����G�X����H�D�D������P؀xD���?"��Ε4�P��Y2@@���?y��{��K���i!�>���/��� @ �9�� U���@j�Q���(�EJ���*�T ���DP
��T**%@AdQD��!P�"-EZ�
 \��9¹�U�`    @ �|7��\(�_|���=��I�p<����v���	V���F�K2zz�f�����_X�Z���Si�Z.�eʷX�M�wS"�+l!v�#��Ƌ0���uV�I=��ʵNӺ�R{�j�Y)���o�b�yR����'(��L˥��W��-h;Y��Ǝێ\������r� �f�5WE�[+-C��H�����SҜu��W�n�ܥ�a̔ �ODl�Rn��6��
�6���5Z��FY��"���#uX�M�����5W�\qn���ii��gsN0]�Z��a��7�m�@һ���j�Hӱ�R��u4T��f��a�q:��LB�X[m�,:�5,��(�V*56��h��զ�໒�9�H��U�omQ�uCiɤ�J�b�¤߯E�zDlZ2�9��*�	%`�M�CN+�t7fӢ̬���n<�U��5�RGr�������`��Z��:��e�]�m�UslR��-x�ťb�ɮ3�ה�wM�f�Z����f��HCt���
�z�Ђ ��S�֚2��e�^�&V���U/ �V�%Իcc�p�`�ӣ��¥::)4ݙf�Ul��]�)+�KZ�Իښ䵊��y�%�(�1^�t�!�nm����;�1�#J�j;D��Su�fR��	x2�kE�r�*#N�ފ���әFT��[[�w���6�Vݺ�\��>j�^1�yX�97Jn�ZH�X�c;W�,
t,�J#`���V���Q0����D�vj�j�݁��{&U��7��t�7��ɰ�ko|ܨ1h{wf�x u��a�4(�X�bkgM亣ZmPe��,^�Wct���_i����G���mI����RU�$�!N��Y�*Oc�����q�ȁ�H�]
%n�{����mSȣ��+Vk�W����I{�6w�J�Uy��̥��$nMuzA����F�9��u��oԵ�R]�zNV��
��5���Y+^�C�^O�?�Ʊ)Rf�cV�R�0���
K6��Ux��,X�u��k�Y1A��A�u���^=yS,G-ʛ�i�(e�:+6Î�71 E��r�w�f�^҄k��$VM��V�A���(�W��iTګH'T&�h�pf�6��q\��*heP��COF��n�"���+��a6$����v�v�^�*%��v����7��.�#O+p?��ұ�k��l/��*�ʺ������j���(�Ln�[w����#Sנ�p*����j���.�+�W�5�3j]��4�f��W�+�T��n嫕n��Vbu6c��Jf:(�Pc9�T<v�ø¬�{i��YX�k���u��S�1��C��Vwk.��X+2f�M�ȒSC�x/m�bCbR�sC��ͫ�Q�e�mVeS�2Պ��6ޫ�d��4pm#��$T�Ɏ�f�]�Z����Da��ֱ���cs58��,u2�p⊅�����T9	�@����V��S���5��.�V1[z�m��=��,術HucaT)��2(,�.cT4��s$AU�����&�ШP�cYBȱ�R�N�X��ٷh\:%�)������.�X�m�[��j[X7r�z��M��I^2"��8Ʌ�z�o-�o-=��vv��3F;63c��"+-V�G~zV�l	���P�Ԧ4����ݚ��v�y3,V���#ͥV��Kw�9Cf�@�#va�4�~�r˧�0'���CSu`W2Ep�E)�L���K&��:��A�ey�휘�(�o��]=�$�6��L:l�F�ڗ!.�'���6
�/Qb��31�hp����*�V���\ɉP�%@��˵1�N���7�T�fl��%����]�t2��1��X2����F�",�����r�+�mM�t�j����ݨ4'*�T���C;�Jٶ�6�l̂�I�,�q��a��ə\F�8�U���A��0��e0�4�)���u�H���Sj��}�0+��Wb��e�,�I��h�r�c�n������ܷ3hV�Zb���Z��ni�Ǖ�p��v5oCu�Z+]n
��;o�h�Be��ӛe�QB�l�Sg!�t��z$�*�͒f��ܽ�/�����M�x�%�PϷ�J��*�^V;$Y��O$�(ζ�k�Y������cّK���c�U��*�v]�7��f������#�ޢpV�{��q�vLa#YA�.���q��=5W��Ϩ`ٹ-g0Y��V ��D�Ŗ��4PQ��l��֓CS�4�ys2��+kic�U�Ǔ3>��ö3N�1U��׺��#*o�] Qo^��4f�KbQˊTy{�+K*��X�ԭ��Qkvj��������lk5)6��r�T���a�N ��*�LX2�-JکA���6Գ���,Q��0�Y����R���ӳ5�mÎ���*�Kw�;��)2���핉�ƍ
�Mk9R�R(�7�dr�KU���uy���W���7=y,P�Є��f������I�yM5�d��%\��(�f��t���X���7�m"�ҷ���LxÀ�j,ʅ�41�0�{FZ���&hȃ�)M��n�i���݊�E�NX��W�uɴ��[UwQ��Ufk�ۘ��0�>�՘���]��	�m�"��&K�yt�[ۦ���-b�rk�e�6^e�[��7��Vշ� ��p̫��ou��;Z��@�Vle7՝CYb�����ST3A;3�T� �ʙ�&��7*y�l��_�Y�%�T}wGmjQL��L��W��q
tu�̓�O^]3z������ѹeI��\�{����u�U��SOFB�[l<ۺ�{��"�y��*�2�ۯ�Ѻ�;ߵYL��5�DVff	�)�sT��Ve�Yf+��������Qm�c%�)�F���3����V*�{NJ��	l���:;(C��m�83%-�q+�yV����
�I&]V��ՈpTERH�k�0��[_10�M�������v��
� l^�N��^���#���bԩb��W��[�P��X�YuB�u�X�����n���fw�i��²���6��;lI�:��^�BbU����N��4b�¢�,c�S��hK�y����n�9pY�(1��ʱ��r�*��F\{�h��V���L+h���z4��u�3hU�w�c٭]ɁҀ�[1��"�J�Ũ4�li�v�n=;v�؎Z%��ڼߞUKU�)eoY�dQ�sq#�m1ob�6�)�ř�f�^%�U٪�'b�W��^ȅӥ����GQ��UU�����jc�,������[R�&��k�/�U�-�[�yF��y��QEM�h�
�k륿)�o۹�h�u��VQ��RZZvΪ�MK�d�%ُC3�k��w���1�1��כ��5B)A��Xh���)9y�+{.'�ۢ��X��Y�]µ�[f�e�u݉v�]P�����4
�{G**O�rԬ���ytt��;th���V˙`��Ft���*f����bT���jӽ��hӹ�h5L��Wy��ˡ�컗t/b]X�3rX�yI��He��)�
ЏfJ���Y	tm�U��)��^F�wV?g1��T��"�y��Lͫ�{�(Tj�'$×tf6åu1m��,+�[l^'�U�Õ��闦K6��;��U��]GuyR�1[���fð9xʘ[�Z��ի(ǵ��hHb�`�[U�̙��qeJ��߬�f�U��!��TY��s�U3 �Zd�)�;�-NR�tá�j�:�GhՓcoo;�I���z/a�Me���P��uULm�oq� �͚�f�(+�{X΋�EmȢYSkf��1���i�U��m��Ii\V�p�X���˧Z7�@�:V˻9��V��b{R���To]UW�u�D��>��"_���lά֭,c�s�tMr�H|)t~��x���~Y���;��@�C�_�|%O��wh�"F��^G����:�
B�l�I�M�����1���4*튉"ȨH(��� ��� 	 *�$����2 � 
�$�H��"�
  � ) �H�#"�ȠH
2
��(Ȣ�(�� �
��H2 "��	 �H*H�*(H���Ȫ��*H �(�"��� �2
2(ȪH
�!"��  � (H�"��@U�#"�Ȩ�}o�������V���y�%��xIn��}��j �x���g* |����RT(���}����z���H�E������y{�����܋)���z�.e�c��Uu�,�,r��w�����ߵǃT��\�)F�uaY�݈YYX�X�H�[�QQy{Y
m�F+�m6;e��]�	U�G:Y2�SR�//����I�$���뺬q\�g;��K	�=8��E��$����eh���t��	�+o�G_�UUa+Oy�L�jd���x����I�ʛ{2��f��(ݪ�Ψ���̛�s�w�|�v��uOfWkWp���ي�tsUćJsI��x���eu�Lݤ:��h�XeG��̓7n3yK5Y�4��{��s��BP}y�{��.�w(�\|r�(6�.���m!%j%�.�u�K��˺��O�9�(H�)Ǽٛ��.ݼޱu!�P�w�R�v�G2[�M�m��m��l6ܴ���t�i��o��od��Q�b���{Q�-c!�`q殻��0Y/E։����Y���(�m�Yu|�ee�aX0ѵ���JLc�P���y����"-9����Y�1�Yau��M�w&.��S3E�v5Y��CV��ƕf�.���&AD!˳R�y_}DY���۹:`��+L�ok*.t���U�dm1u2��m�P�kߥ���w'9JǬ�ԭC��|6;�"R`<r�3ճ�jp�Q����י�Z��oS�o!�;)���v�h��|�^AZqE]��)��T�p0�<���K�uZ��]�����mu���F�hR��Ɇ�v�`�i�����y\7>Ci���:ڪ®���C��;fĉ݋�0�f��j�6S�l횻V��\�5\�y����]ª��k�G3u���m�m�m��-��I0�m��e��o[m��$�˳�dz�cs��Jn)�K��Î�ܝ�����f�H��"7)�Q�l�,��5��*�[.�r9�Cf^��vE7���
�
���Z�<��}�J�%�49��4�1
% �*��z��;3�X�a�Y��4N�v��B����؅�N�x�M�R�hV��cg�fjƸ\�0M��SYU���|,�:E�'`dDζ]�9�7P��Hzad����-.�7��7�	��J�
�nS�M�g7+qc��n(�u��f"ڢ&О����,%�Ǩ5�-�(�2Y�)�r�.�fh`�ע#������h-�J���M.�.zo�AW{�5f�L�����^�g#sJ�PV�of�/��	�U�)z��K��׫�����+�B�Lñ`�Cn�J"�@S*�}9��](E<wQ�7\�*�� $��u)��ͻ����t�Qk�MrWE�$��Z0^l��4VJ46af�+j�T� f�vЛ������Ӯڪ���w-���:2��v��߱�y�cY�N�//J��5�t�T��a[eW-�mM��+��ڧ{y�IU�S��Ű�b����G%קV:�=%r����h8*e#��D���i�T*QnvLY�ȷ!E0t#(c�'����%u��B�YV�w#&��ޢ��^k��lI]�S��
�V;�Vj����gǴ����5�Wh�����++�4�
tԹ9�Ud&a�=�uJ/�7a;]���k+	lE��Q���0�θ�^J�NP�����փ�&o���N:�s*%��e�M͜�h���|l�Y�#�kZ���+2JO<���x�q��7��;�-ۼ�T�%`�b��|�F���\������.�a��^1��T�z*�.��#�r��:M,�G<Hp��]ck��ƽ��(=��L$ķj�`f��o���-6�<��6ռ���ᜤ�Im��V�19.g�1�����%Yʯ^���Ӭ��Y�@�[ۚ�i7��&��*�n�m(�r�R�Cm�e�o��Y-�[�b`���+=��v���%�MɴK��1R*Ժ5��s�y�Ձbܩw�\"�6Pڟ݁Ώ8���Ml����j��d�%NlW��}��.�=�ڙ��B�ziS��A5x�Ɯh�����3��5hA����N,�����"�8�YP�@�+q�)Hgq����Q�.WM}wġK�j�b�.��[9\��Q���#rp�V�O5�W:�B��P�N�u�`��i���ѻy.�͘�,�%d�%n�3u{"^�կhݴ��^��''S�����"��!�8'ϫUd�F�ER�pB��ți�M�ɘd����|���_m.�t�i��x7J���R����V�p$֣Y�3�U��֓VB����:E����W�,�B�ßZz��
�t�5���`;�b�� ���ڛVLo���1^�b��1	���2����{y�����S3m�޽�n��Q�����wj�tM�̢Tk���iq�����U�!;�,�pƼ�[8Sܨ�V�h�xaI��1����V�:�v���up"�-ڳ��[U�Z��V�G��V��Bn�u��Һ����_چ6=S����)��b�1
Y3�}�b���N?.��k6��MF�")4��U1]�Z��'W*�3�n^����1J][�wk*���n��D�Wu��5�yCsoj�h�0٨��%��>,0�+���o�#�떂))��z��!��s7��:�ӹ�0N�;;������([oI���ڴ�s���p��ft�m\fkL��K�:奚J��i-�:0����e�ȬU}Z^@w3^n�ts���&.Vvf�*��I>�����l�鲊m��Ǟ�D M��3u�ٙWԳ>sFGH��Ϊ�2����6�:�YZ�u���;�������=8��z�͗�/"V[9�7T�uaY�����=AS� �:�Fe�홺v�g���n��SUb�)TK�r��_i<�#�B���S�`�;��Q��e�-�æH�]�A��f'>���.���R�d�.mc�9Q��Y۷#��J��n��]�`����-��eb���;RO��nCSnX��1Z��yU[w������3>PF�EC1�ݼ���aߤ�5Y�RN�p2�KMaxYj��n�f�溧osp�ک���6�[��G3)=�J���5��3T�D��5iI:��T��v����j���wػ��2�$.%$*���9��Xrގ5��j������h'�";5��%������Rq<Y��h���Pje��J��5,W'��v�$�7w���P�GXJ ���b���F�^v֦̍�Y*��m,�S��֪��P��T{�η/M3���3'�w2�0 a��>�)Wu��nv���W9[��]Q�����J��|\��[�a��!p�˪���m!�_m�t���5]FJ�V�j�s��5���	�;0�m���(�13uYH.5Y��"}�
f_R��GXs��N�N�9&[��wZ��컛"��6T7�k��^MD�E,���ة�8R�G+r*u�Y���͢v�+fn���`����6��P�0-�3FgGCN��1j��CO=}Quy�"�0�~k"˷k3�-��,G���ΛU�cV��ޝ��}�e%�0X�1���g]�~�ҙ%Mdזj�6�}b�P��:��S�:&��ù�.�*G�z\Ÿ�s�WV��gݽB%h�f�r��vƕRR�ƻ�f�|���Q٩|����DY��v���Z��Н8���z�٦�9�;�&Gd�O^���2�Q�i�Q���t%Ս�O��M����Y��j�mC݉����˸��o���
̓�R���A��S8�}:q3���7���[p�2��PUĺ�V�^Ue�}�,���� �p�Ġ޶f��U��6j��:�e�geD=�p�6A��zg]e���kX5�%�mU�N\��f*vv1)N8��g.�r*҇n)[�b}]wo6^��֡�ޮ�j	L�o+S�]�k���(��G;7��&�b��:��+�=�=�֍��U�#\ܲUVZַM���r0�sF�g��j�����ZRQѣ��8�ż9���g�
��/�����TU@"�Y?�>H	�.$��^K������Q��*:5����OS�t���O^z
滑v+���b�)��um��v�*]���Jr��ik�V%�6���l\Kl�ƘT�#(T�˙�K���g[�q�w a����O<��IKmmuژ�˨-Y�Y��2Ml�C(��⠣����.�0�p�f���6\7V� Y`V�eL�Q�,iͤ�;j���v�9���;KRZ$��c�Ť�S6n�ݛ�W�.��� j����p/Q�jb�B���hl�7L��f�T.Ha�-�6)��f���5�9Dqk�]��ЮVl��dX��r�6�v��xb[1��ˢl�Gt�S]-\)�]�D�k��f8KX�-�h�{ �]Ԙ��0�iM�M�d�V�J�!tK�D���GZ�%�F1�P�]y�J�j�L�K*ع�N��b�	��MX-+��l�iKJ��q�t�r�b�k�E����%�V��-���P��&��T�f��ΰ�n�7l'��! �%��үK���Mշ�P�
�S�#(���e
�\az�-1Tl�bd(�9x�S:����1�Ɯ`�+��<4<C1͇���gXD&�9�!eַ145��b[6M�;��+�r4 �!]�.���a���4el֎M�-P�����J �.�3(2�jWE�.Mx��0�k�:�a�W.X�mf�3Ra���]2�vk-�����5b��;6@f�T����eV:��چ�S^g[���#4�iU�l[ZZ�X�,��fͶܤ��Y�r�0j�5�],u�snA�.B`ѻnЩ
�@6�rr���B�"��ZXڷL���(��r(��:��˪�HQ�*YYh��v�3j��vX��5k�j]E�V%u"9cv���A.�  W��b\7 ��6�Me�]m-��͘rh�mD�m�����`P�e8�[�0����CZ:Y�GB>[y7�#kI�޺1C[@�Vč���^L�5D���v��GLc��c��,3t��r��dΰ�n��l��f&�!��(��+C[[��1q/0�l�o]u����[0)�FbW�
Z�Z;:�P��,�j)fWhA��Xюu����H^acZ�Gu�٠��Q�J����Y�c�f�wݪ�=�����,<V������6�x�a.�Eˣ60Z��6�`G6�	�M��X!u7�Ĵ3�:���Z��71�����e���e�)�`�G��필�;.�l����Ж�!��mW�P�a�9۔.�X�M�]�H9�M#fZl��9ՎͳV��h̦!f�,ٍ���������x9bP�lۛ����ɉ���B�#�����m��7Qk��,ё758�(+]2m��H	���eMs7A�kCe�)��fB��Km�6vX�mu�D*a��B�hc5�'mdo4F8�\�h�c+x�WAȅ�k�|*��|�-�\J6*���B��T����R�騒�T�%.�mhM`�qpV䴹m�24&��έGj q�1+�Q�@5!L1�`�&��TM���e�16�1	��`�f[�̬��l"dfX���6�*Y��� kepb&l�ll��\;eN��훖g2�()�&E�4l� V�YR\�րM`	i
��GgSb�7FU����lf�á�h�����1��
�[ƫc�X����#��SePM,�I��L���*b �)�"K��:��%l5ܤys1�(�� bl�vl����e[+jˆ6�LE��L�m���(�Yn���Q4���v?�] 8��eى�̲�5!%�l�X��Vcj���6�e�,̇��`��܋j�1�.�h�g�UWCi����`7����b�A���]Hƕ�-e`l�3[�*�⃠,�Vܩ6���m�W��T��"�҄�;f�қ�"� �6.�*�X`�u�*��`��imBѦX���:.���v�2:�ؘ�f#��t!�-��v�ܛ��7A2K��+/*[�+ySF���%�YJ�C�nD@-&�ٸ�f��iCJ-&퐫j��3t.
Y�����+ZD4Ù�.��5P31�5+A��P@�J�Sa�+pKr��D��"Fۥ��lų5�%eJ���!�ۈJ��e��љ6c��Mp�Z$�Bmvsa�[��z�-��I�52�
4n%��]FRe���i�VA�e	mo���DD��f�,[�� K�Z�Y�H���G[��Vf�d;d�J�5K�kt5SOE�Q|c�,�[�q<\$(Ӈ�Ǝ�%���#@�F%.�&[�� �h����ii(� ��]���p�����6�ޭ���+]�d����˱��[0��-4�-�9�a.��[`X9�-v����#�*]E���H�Ҕ��JV�.��Gh��a�F��E�f!���Fm+����"6]᎙ɉ�����3���Ͱ�$�����F�¬Eġv�J�%�
-@˭ql�fQ�V�&�<��m̡��Al�ZG�3j0qyf�����\M��m6	���yS��C�5����ˉt�X5���PeVb(g]0�Y��]�͙���B��nWPI]�V\1�j�Ub��5X��W����1��
���3c��(��M�Ml]H7��aњ"7U���;K��3e�lұm��yF����mJꍸe��¨������7-uʪ�����yJ����X��n�R5��61��qE"��m�5b��x��e�̮F���A2�j�0ɰV<�(�Q]r�Y�cfs�P���-��Y�7.�[u�e�\�M��1�n���ϟ��w��\R>}8��X��
��IH�R�%�w���{�s���H$ۮ��s����9�z����{aǵ"�$�P��A)i��6���$ ��i�{{w��G�۝���W�]��[g"��]$x8��J�Z��r��{�]vq9�{�y�#�N(ESXAc()�T ���ay���6��I�e�HK���(a��!1��R6�,y�<��ֲp��RC���3��3rA�{��ON`��7 �]$������~��C���e��-��+���b�wLK�$�
*K�eڍ�!Ph�S� �Lckq�mK�x�v��̹[b&��D��kv!��2����أqf���é�9��]��YcMV�L�Ȯ��60Ջš�D�:i���V\��~yh�_6���!��\�B2�[458�I��J��(��IZ+MXk�(�rV�L��x��U�&�Qu@����k�J�e�el2jg`��j���hۨ
[ ��Dk��4.[�e���؁f�R��͂ծ�\ݫ��KPъ�qkpjS:"�J,$0�(Nkse��.�\W�JKFX��k��\6gf].�k6�RG�е-�QABۜ��c{m�u	��Dsض���Ȼ6"l�cMU���c�M��3�IU�H�����)�b����2����.k)�i�v�e��m��h�9�U#a֬x�P�6\h��[�[�րk���S����LX
d��
l��ep�.T�Q���H�(����K���l�<�v�L\��q.,�:2�f�mlekj"6�-A�@����,z�����c�x�m�[ċ[e�B؂�hs�o#@��h6�6�coA !
,�KRZQ�V����>���Ĉ�ٙq�GBiA]�":�y ?�_�"�m�/-��5��x�0��L�ύF�j���=ٙ;<�=���sc����ٕsP���9��SGٻ[�f!jQ�{K��[n��#�w�����^�QͰƟ�T���n[�W�-�9��7�3:��mȪ�T�8c�^��>���m���P&��c��(!JR%L㎍�|*�i��6�����޽՛�H�l���g�*�U	�Xp��8˾����:�s�Pb�E�s3{E;rtUy�{�l����w�m����-sty9��_�v���g�;�������=D5�r�����ٽ�z��ʥ������[M���x/!VzV+��/���*⏪�E�9����#���`�evBѕ�udՅWfA�k�eΛ���>�	��~+qz��=�w�z�8L7C;��5�iT��wM�9���U5P�w՘+��]�'ّ(�x*�}�*�9�/4dUO��ʹs/�mMnn���z�w��|=�M����D�f��6��͝��s��!���ׯrX�Ke��ܥ]�{��v���$M��=2?D�=���-k��� �j�WKV��QJb"b7�UU@J�8/�b92*�t���fe��=��Ö�g.d��S���w/���wc�ۯw(Gj���w��Oޛ=;���țA�]햆��تI�l�����n^�s�S�g��z�sbN�Մ���F�>���P�C���]-�yH�d6���U�L3W�3w��D|�r����n	�.��V6EuPV��	e�6[Ƭ�DYt�L�n���j��w{��PNSRWI�UUU�ݺN�L�wIo^#��WZKJ������am6���Y���N�s�;�w�t��J����w����+}�_s�=�3����4վ�}�d�>�>�����Һxw��u���|�3�V-綯o�̀�	򒜖	[c6y�^�<}���0�L32�U�6���:�l�c3�1����V�pe�J"`ٷ6�lܖ4Τ�2��e�R.�V�k1fڵ��d�|UD���.��mu0�{S:Rp��M6�c]Uĭ�tsr11�߻�����i�hh��d)E*! �H�T~طSB��}�毮^�F�:�[j����S��mF:�o���}�uɸug%F�w&[n��,D��G���>�1A���<Ul���^_n������ue9�1�UI)XiΑZ�/{�����n�)�M>Z�$6��w���6nuIT�,��)
T�+��j��,���k�{��ۙW6��MxM��귪��|:�9�[�l�zzm>^{*uH�=��]�wt�ɒ��q	��/0r�5����/g럧nz����\CxJ~�Ph���>m|�͵o�x{���ʹ}�H̑ݻ�>�4�4�����%��G��su¤߷Sk��6���Y|���ͧ:#��-��.�u+�tg6r"d$T��(�����.x�#�nV={��{z�t�gM����D���vo�:D�,|۠S�T�-�3a+��/�Z-�]S��P�W�~m6�O��{����-��UTH\s&]kʧ�6R��S^���Y�5��wv������	*�[��GV���͛��y������5?l�X��5Y��W����>}h��T�S��6�w�޾|��=T�trL�a]]
d�B�(��JG�uUs][�毮�QMU��z�'m�z�7UP}������-:Ku[_77�G��ʩ����$6���O�u@Ge��j��y�ь�3��pc!��2�)��[�:�U��(TսۉVn���M�MͥLVL����~�������<JBf��n�ܫ���H��%	�mVj�j�q�j�ce�u�<U��2�����x�Ȳ��9;BW��Z����_\#�����4ɻ����#��Qɭ���6���GK���2�%�{f_wZ<}�:^�������;;��v���y�|���-p�e�S��Ψ�9�	L]��D�5��s����e��Fb�S>"LE%����MhF���������ac]-����k��9����CV�e����`ЗM�tT�K���1X]M2	23����P+�+��� @!5�xu�J�fX�x��0�u����4Z�V��šv�kxD��6�|�������UA랬��s�vBI$�=����֞n��7h�U-��[X�n ��4�褞j��r�,��BP9܂)l��=���
�1��*��8�6&*�J)%zF��wo:�̾n��3U	8U^|�wۼ�fW1t[X��b�gS$�)�BeH�Zs�!l�k�r�,�l�k��1%+�S�$����<iX��F&f����f�ܬ¶��w-ǗO��Xc^s}j��i)&��V)I$x�.}s9��<��E���t�sb��m�랼�8k�K��h)�>�S���c����};=�����%��|������zw�
C&�Bd,�*�f$Dt�<}��뮉��ϿC��ѽp]��O�R���nޫs[|����̅sڅA��ܛ)%�@�>=� " ��O���_�ߒYvϰ�2F�zd31ų,Q�1e�ڐڎR��X5'��[�Չ	���ń��UY�\���V��w^���rc;H�-e�͗��ISD�;���]]t��#�T3�ʀ-�C���wG#�g��)�b����ʬ�t���lESe�9ml��ug�櫹�{��g-:�A͛]f��"�[��yD��f�:2�1V��y�e�΋��a�*��N�۽0:�x��L�]���*�+jt�1�\�0S�G
1>��X3D�u;u��ڻ�gN�Ay1.�]Z�gj���r��Rv��P�r%���-18��yj�4#I���*y(�ȳ��n�4���w	d���?U:�#��2�	^�K}{͕*�1W	�U57�)�����$�%V+9�oP���r�"Ʈ�P��V®�]iݼ�Wd�'v	M�y�r�ܐL�f��;Y���>���BWAy:}^�k`~V�C�_�]-�.�ϋ�>�!��6�_�b�n��Af9���<燖��ܜ���ht(�4�iI��(�IIIT��l8s�z���!u	` ���8"R6ke����ˊxx��PIgKy	`<�a�^+IA�`��ZB���b7Kᥙ�kG�^��l�P8���Z�-��A"�p�*�ox�S���d�¤9��	 F����[�����&�6�BVF��6
�W1��XЈ�F��S� �X�ٽ�-��0��_2~�+�pk>�7h�>����m�}U4E%�M=�;��}�����k��"��u�U=�m�`��0X�k��Д8���r�A��~o{�Y��go��q>�/aZEE�̆�G�������f~��GR�����	)	L���A�X�_ܳ,���UR�z'��FfaF��w�g�{N���>F��%k���h�u�V[;�5��þ�D�=���93i��ܸr��޿��Q	@K������꿶>���cO��y��>�ܾ}�g]{��n�,�̻!\�X�ao]ϒ�,]8�i����}�,�='��uNY������w,1���3u�}� �>JM��̏/�QB����~������))��|C!���~���^d>ޡ6�;���hТ�䡮���d�)(X]�$CK��j�mciN.�Ӈ%u�����(�	aۃ���gDXC4@����7V뮅����sEH5
;��/�,D�@5:YvT�j�Pa�\����KR@�VetιÁ���0m�l�n���яYu�4��avf�׭6��3E��"H�,@x�@[����~���[u�U�.�eK��i6ʵv��~���
4BQ=�=��Z8�}ӑ��P(�O)+�"���,�9���'������X�E�����߭dϣMTQD]i��Jr}�j�<������Ï�ɐ��v��)���ވp�['ז��ϖe��>���Q�37�QfA+j2�5Żal�F�0���0֩���gk�Y�c �s %+�o��9;%,��ج���c��U��kqVê��P�D��>���������٦����Ώ��������E��\
/�����G�QP���I�OZo7w�g��~L�������"XT���~s37���>�zn��=!5��J
f'�Q:�{���>�~UB+�z��YJ��QEQ/S6��B�E� >_���e/�|�g}��fY�\�>�*�ȯ���*� ���2����<0�	fiμ��%G�9���Fj�G^|���T8�]�������KI�fv�Uh���}��l�-��7~	�ۙ�}h��5q�4RӖ�o�����}ϖe��쐔���cM��U@]�r6���V���Wӓ}�گϾA�����}XH1��[+�&$Dt÷�Ý�ϖUD���g���"��O]�y#�T���g�M���^�˳����s�|�IJ����mf_�NrO��ک	G�7p�D��s���9�ϝ��������|<?��������ݣ����[&��*�ep6�u�
cͮ��[�V�뗄���j@��C��L�
�,��P\ ��f�1@K��/| �@���Z����9�@�$��DI�D�#�AH@�)u����Ϟ��D�c�X�kvk�.8��/r�{���~�5�
� �"\����u���1�k�� �樾��l�w3(���@1/1b��D�[\�}mDF�
 ������}ukw�w��P9y�"cT�b!:޳֭Z�� �(.A]�j"bTG�,DDV�ݹ�&qmw�U�g[��{@���w@؈�AJ��fh� g4�b f ����;����"o�D���Q1 ;�u��c��h��x�^�58jL������/$E�($�R�8�[�u� �@�����ks�s7�A���R%�8�Qz� b���S�f��$O�Th���:ƴE�\'Xfj�q|�j��̌���_��Z�YwT8erK(pR�ѕ- %&�C��\�[fg�.��k
��Mi���f�J�	���r\ m��6DA���آ�-���re�R�F�F��eGFQ�����>��{��٠�1G:�L���
���@��q"$�j��0DI{�[X��w�k9�@�&:;�x6�@�"NP��@1�@� 1�$"��DInUo����[D��B�P�ε�u�9mv�z�qDN��P��U�| ��;�o4�$�"TG
b$ U@��?��uҮf��� >�
�Q��1 )�� �\�ur��@�#�&���ꀱq)�����|�5���]�6���z���;�%1�(�=b�- 1��"��D�)�D:5��V�o +]�k|�9mq�H�<b'P@�(�D�11W�2j��r!����Z�#��:m`�76^ת��U�
��"�T�$wB"-�c�k��}u{o���p�r"s]gS�L�QDN�HP@�@/z�ޣ��#�IޖD��k+��
�+J�'�?R��yկ�e渚�6S�F�{��I�=+5�� ;�{�| �;*�~���T��m!�@�	���c��2�~��05w
�l�b"܉�����wkB���u���h�A���0RuO"�9� �`b"s�Iު�]R�4 ub�7~w����j݀TA�C� ��uFCGW�� n f c�h �F(��1@Z׫�p�A��u�u�\��{@����t�$��Y�8� s�j���E��^��lsR��g�j�#�D�5�A�w�k��s�ꃑ�j[����h�kT� b Qz@�DH@-�����J�3�"���w��|�����p�r
��"L�Ȗ 8�c;���8�"�Ah� �b�b�o��d��V�{�c�Zj���ۛ�gVĵR%�N���7��\��w�\먳b+�M�<�@	ֵ�|�9��<@���t�[t�bh� c�b ���Cp��O]Y �"�&�y�kz�s��AȉP@޺�]_�i �tdA��6 �b
b�u�o�sFq��wT��;�:��;��
�<�w�.@q�������;�O=����-s��3n5j\�3V@|�ݹ$��s��NK���8�h� b Qα�o���s�
��"wε��5@순���Q@�)�x�A\�w���E]5 +=gZ���Ƹ�z�qDI�"Q�(	�W�*�w�ch=��Q �h�Hb�(��Q1�@��S��x����ջ ��ȇq �� �E� �(.DM�x���u�h� �F�� ������o�׵}� �� M�1�ʿ;􃃈)��ӛx������HJᗛ�g�̇X�E�`����#£���G�D�@���bv�A��k7>����Oԗ���ɍa�î��PR����7A�.��L�R�P&W?NǭBYt����%��V�k�Y%!n�qc&=���k޽�=�U��:�U�jRE><.�������rxi�A]����������od��';���ʴ��)���뵷;73[}{Vg��$����P���w���?#���J�
�eޯ��ŕ:T-2�צ�ghY�bPB�W7���ٳF-J�/�<#MÜ~&�޼2jW��ZީY�U��Jɫ�:�W�`ɼ�F,k��A�yUx/Y�yH�ZZj�OUݒ�5Y�]����q�r�br�ʽM^p�wwК�$�̝x�Y�I����!=bV��P�2�����U�ٽ�ٮ�"k2�-�{D̕d����OM�U>��b�[�*�ջq-�%�ЪkVo��T���d�O�ٜ;�:��^(Sfgf�٥��U�e��0�z�1���.�󫥕�:��g��۝'q>��p������o[�&��%u���q��-e���3��,ݫr�5 �vû�ʻ�1�b�e��̣d"�W1�k{:�c6����.tYx����ů�i�(_b��Y�X�R��ǻy�y����8�WXE
R��~����?���D����ieK�!C�����e�VQal�}���,��ҕx$��!�W�$e㰶��ŗ�����	>����CB� H���JEW/V�RL;�� Ȉ�FE�*�7Zc��� �<�g��
�b�RR �-iE�X�Ƥ�s�iҺ�Y(鷭��ӲЄF����Z-TkZR!�ю��cl�D$�A5��J���9^e|3U͍2����{K8���Z5{��P����(�D$�4eY5�eFҼ�]a[)F^���$J�3YC��w�s蜷�ѥÙ�b�a��k%ߺ�ĞJ�ԕ�Ŋ��i�xf$�&)�U�)��X�39,�q(4��e�k��K�.���sf�e�Z�[��aR��K����8���+]���`M���BP�n��GGPq��qI�
Ń�k]c�KRjf4bZi�,%cm#�Mc�2;m48�Vů*�YeC]��a���i��g�(��ٍ�m
��CKs@Kٛ��;�+.-4�`��Zm3x,%�+)U��бtuK(J���&y��5�F&����e�����2�a�&a��K �f!
�(�L�05K�����l�1��ĸv�X�Vq)��-�u�	��ǖ���%�/Pm�׮A�����G�v�ɈY��R��Z�Tq��7sp�,b�fm%�ж#43�lM����$f�.�M,����U2n��H�f��l��Yl���:C2�,6��M1��h:�q�+[-���A���B����hT����n���ׂExp"�;Jm���ynP���p��6���H�]FQUUF9uJ�&44��%ƹԺ�kn�\��$�N�%���5�#荺ո��l%Wi����F'�M�mX�2�MnXpf���YL��+���Z٦�X<r��jq��P��]�旄 6dKXŎ�WZbi����v2����Wz>�o���2��0�B5f���X�+��~>ue�_�f�r��O
�)���s�}8��K���O���}9�[�V�{$� VG��9n��d�R��fF	���޽�=�4��)���&�G�F�<����d���8�v��U�z�6�Ք۫]��u\�N.�o�_�'^>_zyv�5�n�x�T�P�
D�����t�kou��p�IS���.��;]˭��`)��lC�̴6s"u'��)[rP9N�h��&���Qp�|?{ĀH������[v�|�,�ݱ䫑N�����WG�j7�]M=y���)m������k/����=�Z[ű��$��!=k?s��/���xq�ɨ���멼�w�y�+��3Z�#��7M���6f:�e�O�4緊�{ם�si�A�MY.�`i	$��h�WS��Ҿr^�o��\>�i6���]��m3����D:�t�н��^^��[{��b[�o���Œb�R�i"����H�"(����c�է���{�x^k&�dZ~mH�:�_���q,�3��۠ڦR�{���M����4ٻ����}��|���|�ژ�t�csV����e��w�_Q��׿=����V��"b����y�}�t����y]��ȼ�5N��2:ն�	+=���^o^ݞ��%�EoG�|w6|��}X�Z�=�>�x������+v��n�J�93ʾU�1�e.��\�JXvi����� ��f^����rbӭ��y�^S��{���QldV<�ƣ.f	��dq3���"eQ`3e(�y����Ѹ��8BP�����h��g�8�YO�Z�<8�N�La�ZA$zy��}�g�wSxOx2/!��z���g�wO��N󷟶Cἵ��ހ�B�Ud]ީm4!RN����G���}~�9sۊ0��*�YHN��mɑr��m&�ͩU���������x{�@  ���ײ�!	~h(9vsX�L����e���&5Wk���1j��,�&H�\�b����ԨcX���3F1�b=����c4�I�#B���̪��UE&Ұ�n4��TX7":�oL�+�y��?M"��t%M�t�nR`�EGIK?���A*�y���a;4�r��	/	)�:���9�ۯz�ܳ��z��>[1�PE���WE]<}k ��J[T˘���BP�cX���f�t�ޝ5U>h�eWu��Q�^�:��<5�P�b���{����B�YX����1�$�PbP@�������F)U�7ֲ\-�V� ,d����R/�nγG������w�V�����ƅ����t��.r�����7n�P��  '�� ޏ߳���6�a<�Z��M�j�e)��ݍ-�o�=�=�I%�y�)]fHB6�+v,�Ë#.6�qP�ԡ(G�L*��*9��/m�<Ȭ��Z����ߧ޷�e��ȉ�%�΍�`h�R
������J S[���۔x�X[<��R��;3.��܈�U���A}�*u@���(����PҬ���{�cԄw3+w?Zc��������Y�����Α3A���Y�2%��%�ɯ�߈Ā ��]������2+!uKnYř(����۔xk��Q9a.��w�>@�\�2������7�9��gڹb>����߽��V:ǚ%�u���.�͙���o}|>�w���^۾�xT�a�����J%���+uh�1���k�)��.����tө�I���l:��q�O3���$�7�m�6�%���۾�x3�Z�+`�#b�=#��d�{mBw�a�ع�ʅzb73�{ؠ4Ҝ������'�x=��RI%���34���^��U��{\2�	U�^̟̄64*QfJBB]k��.�!�͑����ב�S����ӘO�u��˼խP���YuNԂ럺o��M��?�<��[E+�J�HY��19i�ƫ:���INϚ~^Q��є�Ooz�	�f��|^o478�n�ٵ�;����Bw�.��E��^H�T�WI�ө��Iu��%LbzhL����B��:\���Io99�Hyy��C�-j*gaٍ5k��S���0d��ca���F�
BlUJS[�#��uaJ���bVh���`:L]R�m���C�rI�l�*Q��+�]��F0%̷Dغh ���WAZe�����O��f��t�r�c�E!!**D���2,�v�y|�gT�Ź��$�Ub���20��4�7&wt����#t�*H�BPN�Sd�+�~}	� �Yn�%����%N���y�p��ƅŐڐU5��+��>��|wkեV�d���T�
K��-�ttcnR`�EGA~r���Y���_�O��8ݮ��CK���|�7���8ed��1H�Pʩ��5#�'kj�˶�m�q��˙�;�=���$x  ��\y��+���U���p}��[���J�TZ��ӘO2��%�OoJ}P�,�յ�N�N�
ܙN���R�)7�"�{x��Vr]�<�	��zc�ϯA~�,]�d�LnIBb&%
�%L�ğe�(��]��Na*+"�v;�i�!%4�t�_yܻ�m��Y<j�d��h\�;P*�W����b����EV��uS'�@��]��ԬrZ�Wh�xq2+�0r����mޟ�]�l2���&��
��{#��Lέޥ�Y2��V~�}5���vKڊ��V^Rn��d�k;���+�.�9d�4��5S�g��X�g&J(>E�p�ԯk�r#Z:�&���v�p,���;;{q��@�{��P����B�W�������;W������B�av���t�rP��c��c
ut�J�y�*�S�z�Y�q.�[X+u�@�Tz!�H��O5%%n.�`%��ꍊ)]��"��i�͡VF�m��h�5�םˣ�.u}ӏ��M`�d�8\�>��_�wMd�m��.!h��m�(��f*�L^^�J]�XpmV��ooN"t��e����a�+ǆ,wK����}.���#K�`n�tdnl�*dU�(L	�ƻ2F�ᢣ��I��iKZ	~ݓ��*x��L�If��
;iK��.�Ƨ^>|��e��X%�������V$��B�6<Es���"�M�ߞ{�I@�{�����9��u-Vޚ�nZ�	It�YC7�N�y�E��T�%8��kT����^!KX��*qH�f�r�	LlBfYP�H��,���<�% "p�*��k�8	QB�Em�à�2�V��RJ "$>20�� �X4�j�mT$|(R#�B�ǁ�pq�l�#���!�J���3l	�K�h��f�n4H4��T"���ųxj�-�"�{�L�By��#)B��1�%.i���B"D�X¶*"u`֭hT������H(��^]�}��o����yST��Ώg'/d.���t���e_fdȰ�v�JRȨ��W^��N���d��r>t��w���|��kAwdwWRؘ�tQo^ϗ���-^�s��K�9�Or��ɹ�,�Q��0�٪�{�9��8UR���S�ʩh����Y�������3�Ф$��O'�sr�e�̶귒��y]�����J��#�
��}��X���\�f�m^�j�*h�[y׀�$��ߋ�#����泮0�v�s�ܳ	��$�^���u���PЄc�f��x�4eB��A	��H���@k��ʹ���7˳���x�]�Q�s&5�����{��U��WϠ2�s$�}x��ǒ�"�\�n,;�����{�a(J(�ɞr�a������Z�y��QԄТuSDQKjF����ޥ��p4��/�מ�j_�4"��ͮ�S�IFM*�̸�����81}1X�3W��x�	E��Ǫ�ꥥb��kڪY�v(h��2�Ѹ�X#sK��s����TMf3�2��\»���-@�!�+6.�VRi�4�� ���A�qF��X�ݩe��f�gXiZ��
��ehU�����~O�j�ex3(�4���k6 Pg��λ|z�����f�Y��q��7AG�W�;7�H���ݫ�ݴ�	�}�LP3 ��@E����v��Z���iDq��-W�l�:j�s��a<7�6e(�(�Q��7*$	ȗ{ݻn�	�w`"��;���z�,ٔ2Pu��͡3���P�$&T���v$��Uos��K��#����C��D]�݀�OS��ݡ=N}76�d�9�Yc$d�.f�j�lњ-��Q �\�ǈ��v���;��,��)u���;�7a#*���z�E��2gO>�wۨY�����҆���GmV}�s�_�`e��	QCO�a��F�v.���[����J�a��L�߬fm�#��Eɖ\��
"%)	)P%-6�,��YWۻ}]�󚎞�W�旒��xp�U��UgcKZ]��8�Yp�N\�{N�S�p�n�A'JT���:��H/ԹکuB����v�1Y�j�-�V4k9*����QE��w���!?���iWS�Uf��r� �:�ܬu�Ox2���"���"K3�;��N_wo%������Ven����z�.M4��6�0\�R��Vo�������tݓ��-���ܒJ�n����V�k]v��s�.�pd(ˤ��!���CeJ�ϒ֓���*�x�2�@���oo�N���
=ۯi</N{�aѥk����*;Sot��UnX�-N�U�G������ ^�22�UT�?��(���u�7_���=ʛ�-�y�u$�H��D�Q��+c��[ă�P(���|��wW��,仦�N1Iw~�y�f�h#տ�xq��o0��D�E �<���y\��<jQAB�3�w�3U<�K9.�A����L�`�uw��
��k��VK�)GƖ�vO��=;��8��h�4crTZ/�`��{��*����]ju&k�/�+"���	��F�sXr��j�+�,BԱ�� �uƥ(,1Z�3f,��$ĳ9�ȉmI�ػ9�`T5��me��HT���(,F�e$6ų\䃄	5y����+3(m�]UU�VlZ����Z2�kfcT�xM3D���k����;^/:��Ok����Qo{N�ϑAG��ۍ*	3���{W�9,仜i[<��P�c����jҜ;.�n�'��JR�59{c7.�D�n��v밞�Zr�3�++b�"<�J�P�i0�s7y,�s�iD%�wYY"�R�3)B䠤�"�p� �l@�λ���]��sݽ�p�'�w�zS�5:[;���7���䢊�6z֪t���I�0e��ke�i���g4k��|@Ax߽�ί�������i�*���x�Q]����T���kI�)/�U��f�CQ�Q�w۟|��|6���;�B>J��͍�Z�oa<�A=�~�w��z��y�*�2]��81
��ʑ2��{֒��]��o$!�)��(	B>DF�y���e����Wd��v����C�`n�E([��xج�U�O(D�'��cדnv2 �SJsvi:W����O����=�~ xx��  �_�s���'�>�RJ�"4d+1��-���o%ø�^e�"�I%s��T'��{��=��Ĥd>Tb�ݺ��60\Q��,�5R6�P��Rnz� �VU�oZ}�����(���= GanW����7�%�%�b��0�2υR���웺�Y����I�i�{��Rn���[�Oy�3kC�;��`��Q<Z�4k;"�ًv�Si��]����;O�}�@���{ޗ�v��wbϭ*��9\�|���f��.��^늨�� LS�m)�HbI�XJ[����*�P`��� #�nk/{�,�ih�"�(%��sWS˫����	�C�A����))M�-m�{�o%ú�UUʕ���AV�#i��wz����h;k�ӊ(������n������{̺�E��b�}��_"�('@ߥJ���@��S�@��·*^�r�w�]��6&�6&�kT�V��Ċo�t���li�ܡU���%f��7��m����O��sT�`mߌ���%O�s�s�iv��4�G�
�q*,�(�,Ɍt̓���T�|�ֲ��1R�{ۢ�F����q"�dg��k3��V�˕ٽ�z�z���/�uSהp����H��j��f�=G+(�)���v@`��3Y���y��e�fZ[R�IE'�sm���9:6�eZ�p�f���Q�Z�MrY'b(����Y�[5�#(H�s��v��7�r������8U	�ʭUg����՜*aGsU-9�Ɲ<��w�kAImų��/e9���O� :��v�X�F����\<eh��k;S�m����oi�Gl�����Kxq��b���- �� ���Cm0�X1���)�`���A�XZ���~{�=1�'�]+�sf��h�nt$�ȹ�W�7`�V�B�~�{����#B7�Mt���z��).u�ә�ï rb�ތ�,P_�]�g�[���g�	HJ��f4&2�Dbb&imQK�@���`<�k5��fQ�%���xitQl��u"�����L�%�ר� L���f�M)aZT�����7��j%��5�-�@�!�$��1*��P�v�Q֑H�6`E'2P�J��瓼Y :�Zg9��icbֶ�m��2Z�JHr�0{[,`�VB��yW�}�ޞ�]	��V�Vi��V��Pv���.z�W�m1Ֆ�1��nФ�E�*���4ʺ�tm	Hꁮ�I����fAcq�ڰ�n��fGU͵Ѝ�b��.��i0,���;�F�������!�8��/X%hYMXV��I2��cYK�:�,��fkt��-X7FQ�+	ZJ��f&l`c:��
��B��̢�Fլ�+�e�4ô*7#,u�`9���.q��
!lP�1Yx3t��;��
Ak�>m㥮tn��#h��f��W��ьٛWhLɶ�0�lH)�d�Z�.K�+��f�:�X'Qa�3\b�Iecd��
\[�K����F�VX��S@m���m6D���	MI�l��IIa��(�+5��jM���1.�"X[v��M�K,�b1���h�p�^V��0u�t�V5m���
D��8Iz۩���͵�fƭ��XT��D���uЄ2��ܸnH���%�fU�%�4����5�hZ�x�������[KW-\�4�]��fjڪ�Z�5evc-xr�U�ܲ�UUe���,��m��J\�6�����d��wt�l@<}q=Z�p��B�ұ2�1��R���)D�j��2���t[���a�CS<0��-�*��֢�e�!
@���+WXKtE��M�+f�m�M�2@�v��8sH���1k����~�a�(.�fGU�$�|��>w�'*�9[�t�7;�3�(�\d�����^s|�����Q�ݺ�9F�J.�'��ά[�O ˨E����w3�T�VG�r���5�+�EY��Y�};�
"��]��	�o�>Yd�g�RI��3���6�j��2�%[�m\D�B��Q���I�<ܮ��'�O���P�,���=ֻA񞺺dr�.��Q�����ׅ�U+g��*h�kڳ���Zݳ��j���<@T�><��S��l}��W>��)>C���I%(ka�����Y=��*�%2aI��%�����샵�*�D�'�BQ�|����=`�*y���NW>�j��%uІ�y�|�����V5�\fՖ�5()�3*|+�������a1����%��F�ʭW�1�c�uݐy�H]��z:X3uC��)����{=��t$���^A�%�s .����q��F�_~�@�'������W�_�F�BP:���]�RU�a�Dt�o6�f�������(]Ԋ����t=]on??v#�?k_Y�E�}*��JX�^��2�`A�U(L�i�.Q2�L�/�������WJᘂ��/�H�4�B>��.��c�y]����a<�L�q.V�����&b'5�]؏��5�[l�MQ�b����_�p���"z�_X���9J/�����v��Il����x���g<�w�1c��[� �Q]`�<���{w�x�润�b�����Y�����CyƊY~a��!p��SL���HX�R���R5��rR)e����$�6����))[�G��"#r���һ�ڲ�V��WA��f�j��cٞ�<G�qR�"�S=2U�#�Q��x�wWd��#�H��GUH�D%�hCuo�^/�c�RL.dE�V;�q+���n�'��ڙE$�@�sQuG�:|sD�����|E	P���ZU^ͪPqqXK,%�c�KfZ�qC^qJ5��&t,i����aa�f�Y�̅�P���3�m��p�ʴ�Q�U �D�!0�in�e�ټ$s1�"�CF�ͺ��Ͱ��1]��?-ߍ ���eؔ�/-`(D))	e	S)�v�'SwW���k �lr��ݵ�*��"����8��>W[|�>��2�n�^�l&�2�J:�+j]�;�K�_gu!�����`m��q�ȇJ��{��n�v�(]@��R�YqN��<G���(꼞�ʆ3ʋ���f3]WR�$&d�G7�CJQ�o1��]B���qԥ�Y�p(��n���%TL�Oqi��L�����Щ|�;Y8)R��y�p���|b�����U;:��qR�-WqT�	�����me��x����@����}�%m�c�s>پ]�Ύ]ݑtg!(	BpwI�4������y�x����2�5�.�� ��6e�*��M\�k���=�馪�ݽ���#����vV��!�"���bKpk_)��n��ʽ�[gyC�;�QҒ���dl�
���	�L٤ʑlv:�U�m�q�J�o�l=ʩ���| $ �m��>�/ �g
JQ�l��8��)(ͷ����uD��UE�"�J�z����|���{:�I,�W���a�*�
�e()H2�%()�3(1�X�$3��w���+ �xt����VT�%�ݹ�{Xa�l	�{�uvQ��ila�y'*0�SԠ�n�7{u�=����JT��(	���]y;}��}��>��s�a�q�̨�da٘���8���9��"z�:'E�qY��¾ ��V�)�^7�^�U�Q�T�������Q�qj #Uʎ��f�1F[�[J��U�T���4�!(��ܾ���{���	)D'��Qj�k�7_e��(7�QL�p����y���w^Q�q�Vn��BA�eM�����U���_g�n��
B�UO���x�t��_�rx3㐔9o+,�����Uv��!�<�l�#]�T�����`K���f���s�I?BIt��ߞ��ƹ���Je#��68A%���K�[\u�FP�:���p-ieR73Z�](�����	��cb��
3Wd�]e�c� %)6��&[�P\�dn�`Y�Y`*q\Lۮ�,�������������;&�j�X:ĺRb��h�{�<ӺاϿ?=����C�1t�
�#�m�1��"����{��g�tiI����0YIHHu=[v�Us��wrxq ��}��i��:ﹺ��%v���#�T|�S0uP����m�t;�,��Pp^�����`�K����5*���%L���¥[����rh��eO+��(�(s�2�ؖf��U�Ś�n�ݸ�����]�sFWejDģ.)S�F\lE~���@ �=�
�GO���:�ז{��2�gGUh�(�([�f�%�ջ���g����"�H�=Uv&��jz��s���O6;�v�2�P�N"/kbK��<o��w^Y� ��>W٪{���3g���nP��k�R�c"TD̘�	�Q�A��T#�1�s����J�De8�\�F��/���m ���ZVpޗz(��.�罻}v�G�>�A�L�L��0�U��-�g����/�?o���U�Y5����ǘ��l���4�PYո��ed�b��>�2�wEݼ�Z�tKRu�YyCk�I-�l�+�H���&-�v�-S�2�j�z'fTګɒ��
�F�*qn��q�!dhKeK6rr�D������Q���*w2P�������yu�t���ǜ�b+�@eUZU2�S%��˛��*cj�Ьn*#Y8v6l��h3[�w�6y$�"Գ�"^��ˬ��L�{n����-�c$掌I�T�����{�dfaĚ����4���b�1��Lm��y�N*�-h��k�	g4��=x�.Aӧ�n��T�'	T�E1(u�T�v]̃V�JÜ��\��֑�{��ܼ�;��/��v0�a�N���}�S��ݳ���W8%դ�;���O�VK�\�r�^	�W�����8X�5�5�Ikr���7S�����R�-��ߣt�$$�K�òt�lm��p3,ă�+�׿=N<'���DH��T8�Na��7-g�=���=�8�f��,��6�pA-����"��`�0^B+%x#��0��m��5��mb�zw����f�BF/@�
�V����� �!�kMX�U8ZK�Q�! ,���D�� *��D9%�J�p
�G���"�H��
Fp�j���ִcm��ڜ#h�k�T�Q�]@$Pu��z�w��8+�A� �P���mY
�ެwQD���|Y�S۾��Ex N��ӕ�����"bCK�P �@0j��A��%����]������ �Ǥ��T�z��ߟ���4�۲�.u�=f֩�/\מ��}�o=��y��{�#�p�yV���&�"e �/�h"�%��]�U���>�G�+�������D�c�,��U���� ����hY<TC2_�F�����]��A>(F �m ͐Ȭ��_gV.BȲ ��8���}]�B�ύ�bv�ҟ�����t�Ή{�pke���p�<�1���#qk���ʉ�������������~�_��!��]���&x�����ȴW����d����<S�]�(@��.�F+)W�!6%3&e@.8}Y EQ;y��w�/W�q����b��?:@�Т5VmZ�6�(��������^x��@;j��B� �Ȁe�CA��Y���^o{��ȴW���"�͠�dQ�����óDL@C���U&���zK��#���%���ϖ�O���2dnt��9`��+��﫲�A��e@�ƠU��aE��ݩ���lm�lj�Ő��Q{���%KfCZ��x�� �Ď� ��A��EBv&h��\�)`hʤXܹ[m[�MA�f-ۀ"Ы��d�yR1�����]1��!��n OՖx��(��
c�Ơܰ��MVA1(����S�î�)�_�o�X~��ʶ�e�J5D���n��[������{#<}&��_kw��$�ྯ*ޑ�~��=�$U@��r#�}ُ����!D{��W��Ͻ%ZP��F��\��
�6�@���b�� �Bǟ<>�۹==5�F� �D����4m}�܋��|~�8�Af��ot�f-�	�!D.�����0C�(������$u���{�*����u�mQ���By�T�bb�M��х T"�h��-;г�ί:�N�o�;����D3�o������|CK�BR+
�I�z�5m龬�1۹س"�$mwm,���՜�k�[��-��o�|A�C�'9V���+j{���f-�y
a�nݠ��Z����B�k��hP��K�s�=%�@i��i��K+��Z^�V��A�䛱~�l��#��)��1g=F��" �m ͐CA�X��+������י'�����v>#����K���ķ��tQ�����b��T�J&����������y~u��>a��{���TG!j�l�Ǖ�>�� ��)�Io��F�2{�g�la�������ۯ��5���h"گ�%�ő]u����}����*���ۘ�,hUXd�sU�(�S�~�#��_�������� aт:�M�֎|C�(�A|Z�=����ե�	∉��ys���� ����@YS�7�Ӽ载����G�>#bi|Zc=99:�%J�f����q��`�í;C����9hW)����ši��~Y,� ��8Q�@�~f��1�����\����GV��'��Eй*��_���wP��?�ȅ?iՅrʓ߶k����<Q�?[A���#�S�0��"�}@�\���6���G��I����gq�pMcƱ�s�
�*�Tж�zK��TR�W,�I{z��� z,~��H���E/�������۟������v��ϯM�!��/�z���mWn��kaT���MEf����o&��8�,�Chx���<�c�B�'��*Y�_P~��CJ�%�B��	� �m���5�;{�o��^_g�__�����Ğ���C��������[�e^�{��K�t��{�mQ���V�Ӵ��!��ha���y����~��+L�&�|�=U Q�>J6�k�Px,�t���]�:�@��@TAQ7A}�in�gyux� �����,P�p�S�igҐ��jK��u���/�D���*����~~�wt�={��g�y5X:�6j83i��3j�¥T�6�l[�-�eU�N#�`�X���A��k����"�2�jV�42�ʆ�e�)-l���2��lt��&�P�MM���Uq,p<F�Z9??7�-R�Uܸv���l�(5��Ks�?�`|9��e��{�?[����?��Dp#g��Q`A܉ �0E �@���9ϻ�p��r'b�w�{t#�}�'�����`;Q���/�V̑#�����t#��<A��h�Т|��l��OՈi~g�˝=�}����Ǐ�K~!k��� KhP �z�m���ˑ�C��\�.�i�� �|CC�|�9Dz�Q�O��Q�X��[r�D�P�7.�Ry1��� �@V��ݴ���/�a.<�� ��x�*�H"�4`�|���r5ywx/�Q��y�۽�1�nޝ��r4&��F�ʆa^M;JF��~ � >Z��"�_��O�T��qg�D�MY
抪��t�#� �E�AС��f���}��G�� _�ͫyG�i˅�~�ƀf��{�:��t/������� ��]
!�	e�X��n����}Y�[�R�8K0A�-�Y[,8ZWWdR"���,�[�f��*4Vugr�p�0�? �
�^�������҈�5�2�.�?n!�"~mY�����ެ� 8�)��u��~|���>��J�`�Т_Њ����;�r���e��3ON�l��%��M[��	���e�M�4�*�z	�^����>'�>���3���ui|~���-� �QӣS� 26�@2`�U#򧕯�}_�0���D!;�B1/��ڳ�(CA�я�ͼ���2v�aм�3�"�,�An�I+{=m�Xbл��|��f��㹳ZM(�A�;�/<�i/���M羹WK�qѫl"Y���mhQJ� �B��y����F#��6P�]�<�Z������A��hN�����t#��<�g����	���4A��_�[�ާ��L#O�h�u[�!�m�C�D3@���˜�mS�{xj�b��z��[�F^J���}����'�CK������T8T-Ь�/�u��#�|~Ce ��<�X�u�oվ��e��A2�q���j�.�#2bL$� �ğq��"6c��޶���H�B�?@F�p��D��@�8�y�]U0�~�T��ٿ�~�WK���5|ڱT"�f�#_f )��(�ss��0)�����//�Ql�D3�h [_^�U�8���g�T���;���G��x�-�n3� �9�(���M�?K�{��~���̝�}r���?��-���{7��͛q���C~<����ß;��A�)I�ً3j�p�$�of�|QH�����U#���ZѥL����%�g��t��	d|V��I����둜�C|L6����;="�ۨ�7�ne ��<پ�j�^dY<�m.���Ўn�M� �{Nn��ua�7X̺[ޔ��l��D�?p4�7Ggl��[So�j������q�����+�]E�_9`��Ԝޭ�]� ԡ\duX�h��hw|�i�������պzU�U�^�
sk����j����ۻ(e����f`�Њ�ʓ:��9��_����h�-��{�'�%�v�uT�Ru'Aa�V!�!���dn�g\��Ρ�oK�*�哆Yɛ��t�t8���(�eM��-ո6���:���mӭ������>�!�A�-���Ž�b��E� 0cȽ�HPV0X�/,��=��C�.�[Y��i��5�7o��q�מy�xٯN�H���<��e�a+b<#���f���[f�mw�wr����B��tba�P�$���l� �� ����'���mYÍ��{�m�� 9����-u^�X�Ʒ�K�Fq:k2���wqk�աD�-N��jKZ�F���H)�@�m�ĢR$ BZ�R)�"�}�ןhJ��[B��h6�ki��
�� hF��õlc����IMA��*�X7fղ��f��lKщ��ݦ)�e�;ZX����E�]FΒ�.���#�k�+�),����8�]6�v-��c�.�D�lԥ��٥Q��3���Ċ�kK�;`���gi���v�a
�cq
��P���\�s�{3Z^{Ex���v��ys6�W9�u�G���d֑�J2�C5Ֆd{eW�Z0n���k+���]��f6�\+[f�efll�&�Ќf%[��/Vƻ2��(�b�`hC���H巘&�D2�$����Ҍ�E�v����vխ����%V�m���!iZL#@���R������e�-Ҷ�JV�e˩B�#F�	sFU �lHM	\�ra�D��Rh�i�u�h�4� <�&�GB�.�1a.��i�t:S��N�Y����l�i���Ƶ��QL ��,���]LF����;�/dخ��W�+u�i��h�SM(��$��6أM]b���mL\�ȕs�.�3�%�ܶ��UUQ�֫�n`����[eW�m�����}�I{�Ϫ�,}Q�A�%���.X��yu�l���bY��+�"F�ZX.���lKpD�"ڈ����Bb��M�k3�5�4f2$nt�%�� ��K
��X�t&�������_������	n�ٚ�;FmuK�����Q'�|��_�0��U"WZz���`�G��q�A9G �g���g�M7��>���p婛ӵ��G���|ϱ�O�'͡�!�D��:�/ӷ^��t�����j�?Q��6�V�C�PGO͡RV����;����^���F����(�ͮ��Tj|��b������>N<8d4}U �]�ٟn�q7����h�\�t�a��b����Z�x�� �����;7�޸��PԠ������Q/�B��u� G͜����55��W�r�qau��af�s�Ѳ�B_�� ���>��H]k�~��]��ǌrP��nj�MϺ�@�K(��ͫ��Yf���zn�aм�~@P��4m	"��vޭ�>̀Ǎ@��}��ڸS�x��c�~U a�#MT"�~6w�:z�U#1��v�SĄtx� ��|�@�=��߷3ﶗ�&bU�m�KV��m� �����}����׮�K+n�wns��
Ҷ�h7�@e���MТ�Q	>��x*����B���U�p�=ǌv���zPæ��@SAP!� ����ڽv����W2Oٗq���v����Y��~6"&�(ݧ�[0�ܫ����F<�|���HA�?�F\G�T5Q$m��CűT.�A������}y �8�6���M��:!�d YD����{}77w9�u_,�1���lz��U����מO���xk���4م��P�A���Zy�9��W�T�Wkk�d�#�@�ގ��0A͑$J��_H���e7���g>��^����CCg�d��1h^C�ą�"��9ޔE��Dr@�(��D4�-n{~޷o3�u�^ �����hY���3��J��DAf��EU�oj��P��O`�G�*�wi��u7in�U\�kc4]B�f�c�(�寸͚��e�3���@͏�!�b���_�E����p�8Sڛ��}�B��!DAP ��3�x�iZ6���6+�^.����i0�(�A�yg���y Q�@�}���_,�1��A�$!1 �����������B�e�y<�#�{�r�I2�0�z�{6<�0���#gk�?����n�4G@': �A� �B�|��W�Q�1#��=��U���8q�C���w!����}G�P(�Q�2�Täo�nȕ����d�ϸfO��5�񙫞�R�]����6=Y�0]���u�n�'���T��s��f��0!���� �����K�)��@��k�ك�P���V+y�c�)R�j`Գ9,K)Y�.e-CBd1�Xm�Ԛ��*4�0���eM@`�uFVmn�[+L�ʱإ%���%�@�M#�u�A��s��߳�%�:Ej�p[�"�hͮ�Y���e�~���
#�E�D�+�S{7=�B#�o��b�|A� �҈!��/��_^S�2#Ơ@�y�_U��S}���㭪=6���b����gY��&�j��/ A�D�(�~g����qY�H� �{.�Q�ۘ�24GG����ؗ�P:P#5
�J
 �@58˱.l
{^vwU����|'��q�D�Ӯ�w���]{�l�kjFGZ�qn�.Z�z���픇��誑>O��1�p�p�x��Ȯ8A����3E5@��!��TC�¾G�39��^5����-�!Sp�i����TX5��3��}�?�>����n��ٓ�:;�$���3�j�܉p2`�9��D�Nu:�ﶷ�V�B����5[TA,���(�DB�"�D�̭l�uĈ$�x�LL�S�E����j�?2���T��������eh��o@�AQjE�8ĝ�ъ��ř֐p.�7H�]�ت�5V�ha��B��h*�n��+�QDC�{���dI�8J=FH�	��3�ޫ��l�A��)�W6g��J짹S�z���+u���w��MƌQ@����^	��(�����{*�a�K|�',�'ʨ���ծc-����U]�t�o߉=ٻ߷���~/�B4~MРC"�Vr��� �P�_2+;���[�
#�x�>�u�;�"�z|t�BRȀ��,��{��y4`��W�y�k����JCK��g��Úi� "�,F�ukhk�.�EثB���OX�2 !�ڞ��g�=��J��д<A�����_�! ��s�N`q���3=�Oe�K�,� �8�(����}:#אQ�t0f�_��ۓn�A��rP�_���ļ�/�?��u�������Ј�� �۞n@�9�x�Y�,en�.�k�`�Ծ�W��:�
�>�ع-�m+��"������C_/��7B�O�v+�̆5;��}�G�>�ꨡ/:�n}��z�s�ޣ�-��r1�M�[)�w���B��ƌUB����\H����n!����������u}�(W�{�N�Ɂ{�	�!DiDp�1����Af>��(�T���k��yjT@�B���-<�����A(�Q��1���D���ӹ6`i�5|ڳ�?&�m{��4 8U��;�y������?2��RP��-�o��k0�b ��I�gª-.#ij��G�ck�zd��)ܸ���3���@����a-`�-�e��.�����+���JLsU Fl:�A��	���08���X�5�p�t�d�֨�ˋlclBئ�-���;�G	1*Kk�5k��1�@ƥ[�	@��єp�Gb#��>��,Uv�35ml+,A�Q������q ��$���}����*#�3.�����#����,���՗��EU���\��<�x@'���D�U�y���e� �(��@���Y$���Vf�]��e����#�U"|E����<8F4(�~d/{���_Iui<� ��kj��1Q��C!����
QP��M�=� �Ǐ�]H�(���;�N��߾zǿm�q��rk6�L���6ѣ�>�<;�>x��71�y��L�p�������;���v���8�}�Pv=���V��w���Bd^�(C:��K*r�w�ܗ�oT~�O��#�>�?N������"�����m��A�1��E��ȅC_3@�����m�+\^�|�(� �/�_6����,Ƃ�;�$�	e�>�՗���+ǳ�w�<A��,�ChZU}����r]�^�(0�[_Qgd嵾���潖�4d�f���֭զ7e�-�G�C��,!���'�2��ռ�d�G���L��� ϶��PJ�ݗף�q�<R�Yη�/t{�E�Ez�+�D! p�ChP!��³���	Nw�c�li�{��3��(����.�N=OL:���7��{!�.�
��yY'ltC��t;�ǖ�P�X��$�S0��l�\�D����Q�����9�Q}�Qo�Lmy�_f��]�2�j��"#R���<2���"ؖ�Y2�U�� ��s�&%��e:Wڎ`�p�q�����wn�+eM�gRp�ˮ�M�<�>�B/;pH���b�淹�^S��S]���Y�p��|�VN����-�T%�!B	���:�y�:�U'�ꖐ�����#!��q�B�s(��������k���s�ް�}u��ʈ�qV� �"fԥk��&",ޡ��N�֠�?U��5�m�4��Wp�ejr;���:\<*K-bU�غM7�p��^�z^ؼ��N�:'`-޸�t�	��ZOF�x��DZ�S�b�&�����_PX#ϲ6!YkI@�,V,HÎo�=z����T�F)�l8�V<Bt�Q����9n��~�Y#�&�\kkh╻��IcZA����f��88 W����V)i
,�=-a�a`�j����ф�N6��ۛkqI�i�qwspN]֛sI��Yj%.�w1��m	�klu��E��]؎3�j�[�+�UX�BW�s�H�C�a8F,����H�8!w���R,y�m�e��Q�+VR�-���9mj�Dmj@YI�Oᄐ)�ۺ����Q�'O����YD2=�Y�Qb�t.F�<�A���_���aϴ��$�Y@��E���N>�v!��w�y�}��@�y
_3�h	~l�n�ܘ�1��YC\�] t����P��� A{_P!���7Ϸ����%�����V>ʁj$Ae���~�9�0x��7�(c��Þ�z,��D������v='
 �mP?2�=,����>����QP@W�6��B���e��s���P >��Ϻ��Q���%Nk�뜌FT"��✙Ɉ��掲b\���(m¾�}�?~>:���?���͡D3f�6�2�C
ۿ�xu{�D�<x���hGD�k}$�)�Cpٗm5\��@rM�)\.#ߏŐv=wM	;����L�*�ע\��2��5� �B�
"M"��S��0Eq-����仴��~X����	�b���@/n����MT��:0�}�)��}�	����~��-��3{ӑ�8A�܉>�	;��՗�:��$.5�Ѧw�2��mH}G�@�E7������#69���%ݥ�A:~X�mYi9[�<�C�x_�6ƚ�i�s�ѧHUJ���Ө%�T�L��ޯ���W�u�E
�|�V�Dvf�
)
��a�:3 s��[�X��2�k�s�k�XK4ڣG��q6]���]��	���۩n��s+�Z�P�i\Z��eL��z��u3��'��G�n��h4�45al
!�4h���4��I#�G�P-\�p��$��T}a�#ɯ�_Ye,Pm�Bm�����뷩�e����F����\D�ص�uB�"�e�h,?B?N�}z�9��suv����FG���0Eĩ�:��Έq���AЬr�{���@���q�I�fY��e��,�C!Pe���6�w:�Yx#�#� i���'{��[�=�٭\�fj��F�V�n�	A���q���d�^ *fS���]�QD �(�gg�p� �>��MTcqG�%*\s6\�Y���u��'\��ڒD�:�'&�ATT�i���/3�r'���e}� �}��
!���-��RoW�(�ͤ}F�:1����ڼ�u��Ύ�d aD6�dn׳1f���P�D_*!4�L�{��J�K�?5��u�D6G�>��'��h�}o>���Sտ6WvH$qf<FT	"���.��ᵞ)Q̱�1X�H���]���\]vZ?QB-�?3w��y�L�گ�#�km@B:}U U@>4|�val�}�u�����J >�����_Ħ�R�-
!��en��^����p9o�[���}���UfT�O%�D�+U�*A��{���@���#���������A��QK->u�Yx#�� 4;����dmaD6���}Uw�>����}��I*�/N�8�mX �Y{�=��s��5��V�q�ct�
҂Q)�)X��{� �ET�W=��9�F��vQ��|�Z�V ¾#NM��է���{�Ͽ<�J��>�H�ξ̝�^P�!���j������s޻�J#���a�Tz�Q��庅�ut��������,<x�:��P�B+��)���57"��r�]g2ӊ� n.�:����3�a�<G/���A|[TA,�A [K��*��VIy�{�&�	���~:�,��u>0�������M#ٔ��q�q��-�o����N���5�>����(�f��GVf �<r�A��d [B�k9e!��X�;����@��AfeH�I�>DI�TA ���mY�%V���{��v�����&~�@xj~m�b�&�?*A��ɠ��7���I*�/ ~����0ΐ��_Q���}"�����2*|�h��>Y����;�}��9R(�}t[�Tׁ��ծu��Z����{i�u.��4l�=�Uƺff@:��Ъ�l#�1�Q�Ʃ�#� un-R�mI]I�J�Rh�%N&R.�e�3`rR,!�6b�[]F�&
GLлU�+�t45�1�նlK��(1�c���P��6�D���9��+B����ߺ�_)�gl�]7b�I�UģGD|�n{/��� �@P	m�wS���,@�p8�D?6�!�����>��mF�����;���w)Dqşaj�y�owU�ЁG�1�������<�fse���@��3�hY|�!��_]U���D�q?2��t��zd�����۔�
JkB��?6�r�f��Z
f���ޒU�^?q�&�$����#�{�^�Q0�!e�D�]X[�e��+:�k�� �(�B���Ǘ��/����@w(Q~M|��B��m�^��������Rue�ӤD&6M�gN�r0����\���{��J�o���r��
 �9ݏ2�-��Y8QJC?&�X���o�f{�K�K�|Pa�|~g�C����Bet#���W�0|��*)c�?a������}Mf�u'\�'��l�?8�C�'�
�e[�^뱝����3��������"P@Ġ�J�A�C������g>}�v���ł�/v�Q8��yHD#v�� DƤ����2f�^�`�t�A�@5�t���A���P �mP?3�f�$2��1_�+�R���*Ӂ�\S@¡T��PIz$ߚ�{�,uwf�fcޙ0/	��������D4�Jם�'�����!Vny��@�ٜ/��`�4�Q �[@SAIJ���C�vq��F��O��R*����Q�z�()�!HAB�f#���n�P.._˿4���(~6b��������b�U��"����i?W����0��
����wv���	�����wA^đ��Y/��n�5S��~�<�����hx��_�mY�3�?6���.����/t��H�=Xط7�*�˳�mlW�.��
�uf�-)@񛵊�
ۈx���!�	e�ި�
�>�3:g���G.�/�|Qb�����J�����R2���f����L��"fLʠH�� �� �H��;.;��>���7�0�A� a��T#�Qŷ��_�D��'�{g�L�y\�e���N��@�~m!��O��Io?o�令�?~TA�2*?B�Hz߳�eD(�B:~A����=�{��#��S$��7�H�����-��P!��kk���?��}罯�&���@B8`U ���E|����>�nw$��^K����9	������9
o{C���ET4��U��Xb�	�G�7�����.�y�o74�=T�$���:����Z��	�Tx#M��>OJ�Ǫk����O���չj�VoUv�ި��76�B/�@[���=�*��1��Ʈ�U�hU�h�ea���Zl=n��t�f�(ñL1^+fL�;,���mX��b����t�{v�:À�1�p�%�­���t%�{��uT)�r����`�t�3oYTm���o*�N�:U)�!J��)�f<�ar*�Wc,�[C�	XJ�)����oW.�-��2��n�V1{���cb;t����:��ol���Ĕ��o%�V�7|I8�_@V�q(��CDů;"Ô^gX�ޓ��(�cGV�����ݭb�>��[�w�Dk�-�/ ���NV������#'��_7wu�Je�i���Y ~�&��h�37{��S���l��|�=�{ٽ��D���F�� r��H��'Z��s�۾���l3Q(p���KT�D��U�в0�o$(Ҍ"u��U�d̔-%�XKb�ED�Fӻ"F���s�m̺�-��k����D�F(Jrp�$]u� ��c	��D��!�"�֝Lw��H� p���nkp���KVsQ�m+�w]�	v�^�_+y��� *J�D��@ !�e�mh�1V#!��B�Hp��r<�@UX�Z�Y��E�P���o���@��һ趄~����V�
bhb��&�e�i�mq7*����x��jͥ�T.�2��B��&�)�l��[5``L`�t`ˉJv�l�x&����
5p�m���bQ��c���Cf%t�!�W��6�nm����
�GU�K����5Kpm�[D���&�ؘ�frC1���tM[���n3UL;kW",��4J��2%�. ���p��3���v�F�8�9�.a�D]�4���3��k�+4�q�:�it�8�"�,׆b݆�%�&�5�K(֣��n��������������6̦���o��1o!n�aÖ�uf��g�M3�͚dJ�pb;P�qs[3�
Z�腂�Ql3��R�͋��-�k,e{>�fy1�!�l5.�CYbRM:��WSV��u����.���6�6��R��f�\�8�tB��e�W�K��f[H�g�.�&X�/�ur:1���bl��L��.^$�Uyu*�����5W�%9]S@/
�.�7h$��ɳJjU�B�"� ����+-�fUUTs���F�mEW](8.�OT��=�ۧF�Lb����FR��hh��j��Fh;�[k	��@�8��� l��-�iTiSj�M�Y�<Rb��lKc�La�7�a��wmZi��h]�h:[�m,\0f��V�Yq�}��ٿ&�l�A��G�9�12�S2&TG㿣��>�#���mIwI~#�:̕`�D�F�Q��iT�_C��K>��Own�qց�	��Ǽ7���V'
��}U������o):���^z:� ��,��Џ|��VРF��=��wr��1}��v�eG�`8��U@P /�p�"���_8��@����t?2<�ه6��>�B�UT�i��؅v���B
��ͤ�>8}UY�����/p��2��"Ϩ�PQ�=�*Bt�e��rF�g.w�hID'�\�ݽ�q�k��5Bz� C>��&�s�m]���~��_6�|��b�OG�P5�k�h����OU��{=�{����8�~g��*���Q���/4eSu��ח�:/����S�0)�@B,~m!�T^]Z
�'��w+�S��9��D�7�A���ܗ3jV5JѳhA��M��Uwbb֡Da���T�ݝ�{����N�|~��ؾ-|ڳ�?3�Ӳ?����B��'{��L��B�B,�ߘ���D!�(�����Tx�/�~��X1�;cT�<��6Z���,�+]�YY�Uү�f���]#�K�|~_b������,�̐j�k��{�h;�F�#OO���A�<~�(�������?���9����/k�4�uT�Czz�Jd4�f�������tY�	R�����"A}�D�c}�=v��6*�ݬ��|���!��@25v��'�tuЩۛ;��;�p�2 ]�R��z�����<Q��j� �F��H��t��t�~�0//��
�4}R$�#�,�>������=���=$�H?c͋9�م՞睺Q-�Eܑ��Y�&nӹ�íK�Gƾ�/|~҈k�	m
!�hU ��Nk�|��R�ϻ2@���'����w��k+�뒙j��mj[���F�������0��Qm ʧ��<�2`^C՗�{ (�p����C�?v�1c���#xG�@�O{�����b }�b���?O����mY@��
�����N��^�;��?!�B�i|�ͯ�PM��0���@2���?L��y]��Y<�:~�B� K(��I��;���os���}dqm �i�K����
�W�(���=ۇ8h���:���w����e�^��������e�f4�3F[Y�l0A���P��q^Z
�76�5�9�ET�Ɩ�f5��va����Pn��	��s�c8��%�	�s�BS�MDΚ��M�j,��m��P�������&V�Y�k����-�s\�k�j�h2�i���2����G>���׵�=HB�a�A̡@�?&�mY����vv�O�Ǧ�2�z���A_G����z�h���-Т�4'���*�w{�ys��^����j�%�CHqڼ�� FQ�T�yOvg�A�>���N����!RmF�5�j{'�u��O]vu;����$���DQDM@����?~hw׳|��+`Ŵ��2X� a�@��|��w%����^-[�;}�/9U/O��=�����E���@��C�ͯxߍ��͈B�ݼ���n��W;�`�I����y�%,��G�H�{����R@'� 
"'�ҷw�u+ �Q�[@3�ju�y��6tف�{�Qr���D2*�׽^��Dv�:���+;=��.rRK���9.ޟ<�A8}DO�TD h�.�P7��=�ʤ��H������J��m9�Sc�3p�e��\��w��� |{"y��U=�=0/!egK�0Aha&� �@;@�~���	��;Z0�?B+noo{��%$����mv^�>�G�!� �$Q�"��{��g%BL�uW�jׯi��w��ku��`�;�;Z�M�u�U ��H���"�G���)��:�����TA,�����zt����x��z�mߴ"����P!�����C�{���^s�}�/^J�U��F��V~e��k��#ILj���#Ej�6�A���h.�+5�&r ��G��_^���ʤ"�u$��܀Ⱦ?5�j���������\��t�{o�y�����(y���.4��G ��7@3��T�o��+��˯%$���A�ŴQ8�)�F��At�ChWd���~U �t��״���(�������f�H����+Y�*ArU��l���~�mQ����iu�lYÖ���g�<���@YY�B�]^3���ґ�l0de�#P�jɲjº��aD�B�/�+7{�G,���r� D��>��4A
���@��D8_�����fЬȷ~n�U �a�3 
�#ރ�"M�I���h k��j�U:t��׏��ϞF�<G�FAТ�N����h,����/^JIx�x�B9XNk�u@~��͡D�dJX��ݡY�m���@<#�`���\G���{�VQ�����bԹ�k�#>���ea��5Ǫ�1��]yD�ݲ%4v��T*�$�f����-�R!�[l�A�62���؂���)+-\�Ý5�+���t�u�ZM�ɔ�iWF�^l���Ke��V�R:R�df��
�j[�YV8pd�Z
[�_�w���e�Aj��mk	���������p�UB>��[��?sЈ��J��~ � ��!�"�0FF��*_r��$q�t�{�Ϣ{	���A�WͫT'O���sP�!��!�6�~�����#�O�2�g�G�jb�24f H�r&&~������Dx�����zz^��΅���!�(�E�X�ŢWI۾�*�G��	�a�d�{����I�>��^)J�`U[�h��ſP'��x�l�E���gg:� ���G�!/�h"��#����k��W���C�e�1�n�=�a�1�$Z��^�굴`��>N g�fS��s�G� 2,�7۶"�F�:~m ��D���l��lI/<~�(���,��BM�D0�9x��y]���FA?i���YUZ&,�dZ�~mYP ����=��;]�5v��i�8�� ��Ae����uk|�vn��b�*�� Jc :^����m �̇�����lI/7g:�D�,�"q�4Q~5� ��c����۲$]r�m�7D�Af́$UN�=�/s��a�آ�EG�������嚱����j�����UFUJ�>ԧ3*]��E�S�9��a����}�oE�m�^^c�y�߱��U�+����:��kr��®���җaƙ��v���W�6�˴�K����Γ5X;�֍u�Gz�,�l��@f���: 33F��޽�o;P���J��[��:�[��C���mS��0����6X}ͫށ�W9���M�,�w(�L��d���5d�1ajf��.rK�4/��C]�yv�`��(�x�Ytj���D�kʌ�o12��F�/�����v�-Q�ˊ��z|�J'�ʁ�)T��Je�I3ue��2�n������U�A�I��V@��n���h�0ѫ��2e�έ��K�Ϧbՠ��S���5N��S(B�H��q7(h+��e,��v"C'����M������ջ��J��`(_�=y�0OOG�0�5�Y��z��{���Xt�� w��z�����7�� *���y���[5�n孜�ڴP.�nPC���`�V8 �z�Ͳ�d{ڎK��m�2q:�U��-�
B �'�U� ����sxU�%Z��D�%2�b������fu;��8�E�� .�m���ׁ,$�08��lZ!�R����WWfK2m`sn�t��G�PHO���I��m�{�`_� ��#E��n�d�|o98�+��8��C��o�ʻbIx��-EG�|�2	҇��Q�
�f���vJ�۽7D�<A̐(��qͫ�����w_;4�����FK�Q�X�s5����=/�̬a獄!���m=+�9��Pz��@�(�O��P"� K(��ʂ�/�C��{��]�$�����j�m��sA1g��	BMM�y�-���t83���_M]G�HUK���~rx_D!�Z�ҡ�E{*��i��v����G&��ʡ׵`�w�C�`�m����<��L�t˴�7�7'�ʽ��q�v������ϊNhR�i�X�l�t6ڒ�TtU~y����n�o��f�]�q���))i�q:�L3��w`�o�����Ȍ�5{��%�)�����-{��d�:|�y(�bf\�y+Y�^�M��� ������RI�����r��{�^�pz�=e�H��l�"���ˬ�L��Q��j�F)����;�Dƅ.�t�H�d6Ͷ��%�� �Y71��9k����9�̲�3�hg�`'5)���5.��qU�ى
mfֳ��,�A�5���V���3����`gL��B]���j,p"�[��b���<�|MR:�6�m�1�
0��f�g�>�ѱ�v�Om��V�Ej�=jm$���j���˟j��m�����ۂ#>
[�) u7͞�IQ��nW@�	-����z�D"�e���x<�ϖ�5y����P�R=���b��>o��w�3��~�z�����h��f#�\���5���6[���8؟}����
`�:S�%(����{	̭p����cݟE�d�5h5w7�����9��jz��k��D�d�	b��2�+�������w�i8Wg׼���fJ>E#�ZF����*m���p{��!���Y�Mt\*K��{}��9��djR޻:��;|�ɟB*b�+͌l�Z�&�\�ߞ*S��w�P��P���7T��G+,`���N�lN����YB+��7��M��A���S�z�TT���W�ްH�b\�XVr��lή�Zj>ux��u�0���um�L�U���z�}fȀ��]:-^f�������X�%]\ٍ�[�% "X�&�ej�ؖ�9�?>~iۢ��?t���� �`�f&�CG8�Da�b$��g�2�u5}��gd�v�S�ׯ�Q<�9�k}�tFd�}�ʠ�]�Pڰ�;Vؤ���X�4��D�>rz�,�FYwW>D:[m���<׹v3�#+V�w�9ʼx+��u�2瑷�H7�Db�u�yuB���aG�(EQa쬌T��wJ���p�7�^<؃fb!	Hd5�BJ�rDG@~_�y�T���o9<2�+j�=^�,��\>ۺ�YW�o�y��φ��LurS�ȏb��>	w7]�N�����T;�n����bU�%`���^v�{�Og�,��u(�BI�kq§���n�^vA�F�!nt���὘���ZuLm�4�51(�*斻�n��'�N����@��0�vɗ ]�č:WMhn��S/d"Vg@�A��m5	�a�jbU��c.xi�a���V��4#/-������h���vˆ��Ͳ��m۩�������DnF�D�ߓ˼'�6��blT%�e�`a��2��\z�D%�c}�C�����0��H{e��i᭴M/�����u_������k%��]�Ac�����?<�W��Ym�^=����qqwև/�����U�x���jA�]��Qᆪ*���wo���|���U�h]�T�_}}��âu��3aH�<��X�vC����6MXUv_���rl����G�5!���TQ�Uft�9^X�rh��$��3��K�b�z���T��]������xMT�Qi�������
�������m����3��{���|ܞ�� ���o��򯶈�;6fv�����=[�lUW�w|�_}�r��U}��t�'����н��i�۰e#&Q��Z�u�a��5M��F�<�U>��\�y.|�����ՊER������]�����ͺ�x��]�__6�s5\�K}��u��t�\�$�q9n�]�����f��v�J
���(\�X��������w�VO��p(��
���YT�'��.|���w���tF�m|����q~����]����3؎i�6�t/���Oz�P�_+*���Y����Z��D�uU�V�k���Q?}��Ō߆���USU6���Pn)e��<���®�&AԱ��{�w"�`s�����y��q�P@6��#���g����v���U�᥎��%�u^YĮ�`i"s�2nn�T�\β'{��)�L��9v�˯� �m�-�=a��7^{ު�{���E\
>Y�*�%�tD�J���Pu�CFgTa�b$���o>x�Oݒg��g�>\���3�c�ƙr*�=V/.&�{�k��[���&���~�o�Ǖ,�І���Zxrw���{��w�q3�i��G4c���#�$��Y�����n�!b��k��Y%Kr���U�����ƛ���7�~����C�c����D\����_��}KVg"�w��9%��*!G�~�QD��*r�E%�?6$#��F����Ō�K�Ⱥ�&k��vߍ�q����p�:�b�KTPE!"�Q��k� `��QH�	QD�*���\�B���*���m��8�DQQ^�DD�q$���Q%DQP�z�ں��k��J����H~��i8��Z$�*>)Z\�-ZJO�>�o��AP	HT���&�3������9�����P��0\��(�,�4�E����.���W�"m�5����4I�I
��"o�4��Y<L���n�UT��x���:~7��8���
b2"��$B؂��C�	$B��� {��y����6�?�_��m�{���W�t��B���Ae�'����ߵ�|��O� �~�TA��?e����9�v`�A.�\A��5m��O-�ʨ:S���X�^)�ʨ�΋�0`�Y,i&=G��O@�$I��|�~|0�b|����&N��(�Q�碜0q�b����/�( �q�:%섽SD�*=%�Ddb%hi�A��Q��X*���?=����f���?���_�@<��(IA�(��*��"���a�h>�<����;=Ǭ5�g�L!V�m_��S�`~$�8��?�a_U���F���?�B����*գ�L���Y�>q�H��O�hvXOh��G����j|��=G�X�p����9��`;���]?�?a�(�>'�i��	�d�Wڹ>�)�	�OÂ~�����C���؛��>(*�C�R��X����'��Մ::L&��!��<����J�'� � �O�
���p}#��"v0���}Р������~`�0/XL���hl �ȇএ+ ���Z$H�x%��Q�B���i��
X�
�l]�}��6.����]���������6 _> :�J��@�~� ��G���˔tē��%��ʊ���������O!r9������I� ����9��'H�F���>o�?�A���<�^����o��?����K�>������'�9'��L
�yҜ>1>�>��A[�JY?\�'�������?�H*������Y��d!�SH���~�:H��*�#p0|�l�~B~`l=ρ�������O�-�1>���jh�����?wȽ�@%��7'���ny�M��C���yF1Mϒ�t�}��{������p��6;/�d�w�y�U ����|�{��j�!��=�����O�h0�^��O��'���x$�,Ro�2Q�:0%�<X�� ���>ׁ�>�,DT@?����?�����������~������h������Ї�"�pa���hr�3�i(�!���ik`�>����AB��?�"����������)��4�