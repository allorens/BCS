BZh91AY&SY[�+��t_�py����߰����  a4���� �ݳ� �(@J�ݟO  ��m�Ԩ  ���c�֨
�*�R�
)TU (�P� �B 
H)T
Qs�@(�%   �>�l4O��TR�T�v���=��n��w��ͽ����۴{���gv���9W��^����� g�
^�}��Yn��ԥ�+��t��p��{m�:Y2.�޷*<z����y�^��j�7&�ݒ�  � ��S�A�К�f��k��{����\���@Zo{�G�O{��{Ow�^ԇ��/z"t��魶. �x>ޥ�һ�IN�x�yЛ{���������˱K�w�Wm��nv���s�zӧ� �@=	;uWã����ֲ��{������{A;Ķ�wq�Ǽ�{t�c�sҝ�os�lp {聽��M\��cם�U�Ov�m���v��f��w�����sGGg9���x <   ����T�w���w{�6v�V;�u���W����oc���wW��<�������9�� �C{�n��yOs�^y6�z绹������u�JO��w{y�n�sG ��   �Xvp�v�19����'�����U����������ݽ�]8 >|QϽ���� ��sc���ݓ]:�n�z{����y=֝���p��    �Z�)"J  �    �  �~�z�JT�0� �42  ���)R!�b2 `M�0CA)���� �� d� $�A	USL     `��I *���4�D�M!�ڑ��O�<@US� ʕJ� ɀ bd0	�'�|���ؽZ�E�,T�{��E��}�`�i+�>H�����(��Q��� b?�� ?���*���/�F[��(Q`�hf I! )uP���rg��h5[�M@	 �"lb�I?�P E�7�����O�_��'��i�\ï�e�%K�����j{p�}&	�'>[�)4�OS�o?t�yoV��w��腱yh��^?����uy_-��o�}���ʖ��|)k�e(L�j�E;�:�~���Z���`�V��'���k*f��n���8������N5ۓ�s�{w%1lOI���[���ʉ߭�<���wV���t��1�5�\ŧx�ڴ�ۋe>���mm�ݧ�I�U~N�ͥ���KeWi����:�_k�-n[KU$�+�)X�KZ�[얥�eJ�r�-��%��s�KZ�-o.��{k^�k_w�j{��r�R%��k�B�!ڔ*lB%�@��І���s+Z؄Cv�XЅ��EC!�,ކ&�*�.!�F�1���~E�V�Z�V�
���b$<R��""�s#�B���wkb�۔-��hFd12�DT?�\C��bT��|�F���ԡSb9B$��~�7���b�R���D�Z�!�!6�,��!��"ȁb����;��؁���(2"��N��\�"Ԣ�b!��׹��^�V�"5yrS��������y��[z_�}��ܖ��j��g>�0��i<���c|Z
���Y���z���C��~P1p�5��x�n}����W����7���i�j%�r�_��Zux��w�cji��2#�_ƾ琮��h�#^���V7h�sg�"V����Ȉ�~�X�^������$�,�uj˖�/K��M��+��k�վo)�_y�fc�^g^���)�7h��^�{�k�1��k����֜�Sy�<��cO1�dD+C��" Ȉ3�:DF��Dn�纎��H���"U���Y�dGP����ƣ�z"4����w�#Dz�=W��Gl��Ȉ*"�p)�t��l�s9޻n�8r�DB�n���F����z����G��\l3��åD��vS��g29�k#""�"5
	�����lק89��6����!H'\�e����ַ>B��G�TZ��o~�m�����|��]�/.!1M��M7s𳗖�g���7"�oVb���޷����m��m��Q#sJeM.Vy��~<����&���T��v�ܛ�Z�I_{�~���w垆�~�^S��K{��O��
����Lߓ�M�{OF��O��?,�7�ŧ)�qI�{YN�7�a�&�RbV4O��7����<堞��N��>�e�I��a�[��޺��%��ے���2Ӕ����w�y<��y9Q�T7V7t7#{>o�#�5)�(OV��[���[����q";��ڒ������ZT����U%��i-yZ��J����F$������7jv��rm|S�nL;&p�ѦZ%yo����yb:�Պk�؄v7i��'	4*%�Ml\��}�t��!�n�m�R+� m�hX�ؙ�PSb!kb�V�P����v�f6,Z!Z9Z��sm�؄r���B
�,Bm�V�P�G6)P��.L��J
lB�S�F*�����x�֝ԛeM��kU�KS/��5x���w%)�y��j�,��V�Z��ZskPǪN2�j��iN���W٢��[b6�Є��E6!im���7�Q��&���
Q�D�t�D��b�D.��&�jr�B�B�&"��7.�p�3IMS5m�j�_bs�-8�����*��<�[W�i���3zO�koUĶN1M\���v��{l�c���}����(�Ž'Ķ<^并��lk��{�;���}-ڜ]ί�54�c����[W�L/�;%��6��y�I)��ix�cR�[�k��j���I�����3Kwr�R�o�ٹ�n��������{Ï!6�누ߛ�����~�������6����O��7=�}�|���$�#J_��}W�|v����ވ�O��n��ۧ�o%,]ϓ1Ǳ�y��.��l��1~[����Ï�>�ޝ^������g�?�/��^�8�y��įy���z�6�nm����9b�6�Bޗ��%�k�Z��$��bֺ�m�T��qcS[ًZ�[�=�����Ҿ�LS��2B�B�b�SlM4&Є�p!h\C�r�hX��B�J�p!�kA�ұU1
p!��q_JU8B慉�������T��BmL���F���m��б�o��)��F�*��-L���r�;R�N��й�br8�*!��KKp!N!5��!2\V!Hp|��6�RhX���ÎT���B�b�
�4!3j��r�B���B慉��iR��B�rt�BmX�����x����o�^8�s�+�(X�3�JVS��~Y숿���v�n+�	�)W�Ǘ�ҝ~��")yN�"�/.n�\B��Q�˹ҍ~^�+M`�X�z�E�r;b1�")r���#|�j�A�~��H�#������.t}����.���3��ԟ6�O5@]Z��z�X����e��z��*YT��Η�N�����qs����ug����;P�����w�8�<�N�����������:y&w�W�>���G���Q���ݭ��/c�J��E�P���p^F}KOi�i�4V��mu��T�=�O<S�W�dG�^*���gDa�|ϻZn�7D�Q1LE��_tF/{���<Θ�܈�k�"#�Ȉ�Do�ǹ���";a�Cވ���\��â6y�sK��2r"q��vDi1�@މ��[j�7P���A���s���}�g�>���1��g>@�ָ۽O
��c�Ǫ�89�'��>�^m��xb�>���W�>�)�0��e�1��|K�}�f�uӈǽ����i��`��hS���co>c���;�g���^����Gߵ�:1�s�e�{N9l��q��%�/a��Ϗ�{�<���u��p�kH���S��DwDY�f㎇�f#vb�z���K�Q��-ҍ}�N6a8X��wc�r'�|}��V��-z�sn�G�B1�V1J��,���q���=�"�f8�G���b�����I��BAN1J�b5š$q�V�1�qi�Z�Ϙ�D��b�z���>!��%8���A.9Z'||k�
v\Z�B�p,U#���Rk�8q�T����Q6���qjT�1
�p!qN9J'��|C�
Jp!a��\r�N8���츴*1������R8�>)��&����q��x��9�`q)��[n�����[c�G�r���g<�-����h�q
~�Ћ���8������D:R؈t��z�W1vc�O�Kh������^8&_�8�	�ϐ��Z�\!8�4��q���u����'m���x"�#�Vݢ�a�7��b�^��(A��h�q�F��X�|ϵe6�x���[b9��DB՘��%� ��6"�e������g6�s�T|#�G|�^�3������ӱϛ����MDĦ✊r)د��#ڏJ6>��[�����j�[�W3����������W�~�y����&�Z���Ȉ�" ��1��͈���{�>���w��1o�a��2��x�����U|�!b�M�eh��]U���r�����_�a5*��?�YO�N��%a���
XIkھ��ZO��ݿ��у8��m�Œ���1��b})��u��W;��yN����?���T�6���@�<��S>�qci�P�i�}nON�qR���5�1e�@G)x����Q��ew;n&/�w���W������ҝ���am�d���W�c���\c������&������^�7�R���=N:!�v��v��o�-�Ww9+el���酑�ʯ"����ݯJ��v�K��l��g�kn'�S���ym͙����޲�|f�'��/�{z�������F���Yш7��Fic+����lnwз�7����u�n_fϣA�}�~����ji��ǒa��,�='Hf�w��5	�gcU�o^�a�>��LzK>�����=�1G�uݳN7] ���x��L�';��(�t���㢱����(����g%f�p��g�v�^�kޞ~��)v|����Η����i��&d�]-FTI<��r�:j�̻$˓燽��S~�dew	��l�6�����Γ���7a�15�w"��N�K���d��v�&Ť��c$�x�;�߬�Es�!Fzu��e{UC'��0-�����͝�kXJ5������{_djaֽ���K��])�`�U��e�gd�v��~���D�.�{V�f:�5�Q�r�&b�ji�}�T_qݙzv��9}I���w]�e��w�k��������]m��w�
Ub�QJ�H��C��ه\%7��}$��釴�R;�s���a\TS��62->�D4N�)�F󿳹se�Ŏ��vw�I�Q!����-�'��ݕ#Ǜ�}M���B��y^ʽ}�K�ߎ�}���Z��\�n��ݝ��&u�����D��/��}y���z�}��p�=�xg��Wr�N���$�/^���>�}Tw���c��-�0A�1�H/��q����=�7�������Y$���;��v�Y�~�roJ}�����O�鳳�٫�d;ƮS3��Y����ڭ�h}Я�K5dDcɋ�D���E��e��{z�a�w�w~�lN�=0ݫ���a�l�n��_�_K[{^����ؽ�r�o"��N�����%��vLw�\1N��\�~:n7���){�U�+�"��o�!����gdlgD�r΂gh�WΖ�E�c�%�>�Sݝ���6�D�.�~̕�ӽ�4f��Q�n�T��#)d��9��`̽W��ݗpKϣ�V=�듹z_E5����	����{�w�ˡ���.��ʛd��tg�ޛo�<c�Cr�,��Y���W�O��:��K_�3O<F��r7A|��Dd�j�s8�c��Xm��Yo�7�j��WX�ԦaTG�z��o�!�����W2�s��B�;2��wn�g.c��>�cߙ����s����y�#`�$o#xڷ�kq��~͈�����Vf_g��s���J�(T�.�n]�V�Ș��Q�jӵ�ߩ�g�^E�h�1�yh̒Ol����G��L�\`q�5�"�,з�ec�[m]�J��.�1�R��~m"o�)d�A|gw?1Lo�	%���usS;�X���ʫuj]�V=��|f6�.��n�xl�����*%m�w����ŷ���4ɫ�R���ͱ��U��"���{>�P_|����th�	0��q3����u�wqn��6|]F���֏^ڎ�F�e�Ky�]4��Mʷ"&XQe��1m�e��'C}}}��W'_�h��۝�T-v}�V��o�T���8�i��^۹��;�z��f7��W���ӧ��Kf�%lLS1�v��ܢv�\�s����uj��a�
��j[�D������,[�F��>��v�F��U{
��&�ǎ4��bլ��Rp];�!����=�ݝ;{)�ٓ��L��7�
����_ۋY�̿�?��v�a|]3_���%�^�2p#�����Hɑ�7�)�e]bdFNd���y����W��g{�*��e4��0N1~�۞��c��Ʉ���fL�'g}�L�����?^~��vw���aS�3�g����?mj���7Dn�C��3��u���=�r{<��}<x�d�u��u�Qؽ%�{�a���VN���gM�<���f7[:J͇.��k����=�nˎ;5����ߧ���P��Y���R��dw.:]��r�R�W��>����ʬ��m�JeˣjM����˹0gr1
/3zE=��i���N�z�I���'"m�ڻ�o5I#�#�]9�F)U����ͧ]��9�.
?C>J���	l,�ٱ��'ޟTǜ9NՕ��j�IW��k��k+�w=;��{�>�Y�7���̏T����Ol�7젻��1dO�ǝ�GC�vaүm��4�w})�G����1kؽٹ�3o]�����Rˏ6v��r�Ie3�+ޙq���=�ﲛe�{!�&o�2{=�x��bq�m��ӕ���F�^e��z������y�WY�7Ue��j���rL�ƻ�Z$���W�oLa���y��2���w/s&����K�2��v��ɐ�6Gmx�����+I��(7YF�n�oݢ�hs>j�	�9<)\�<Y��
�������ɐ��R�ŏQl۶��~���i5��T�T)��D˾�U�bYYz���9��SM�3�92�Mԍe���cSS�^����s���}��#�>��=���xk��w��ǻ���=�}�o�n�+�=f[Y�����~ޗ�\����j�5gs}������Z�}h����)�s�������0�������zc7�WM�!��ջ75���>�ɇ.�*����T�e�dPMT�j���y�����Y�mfU�sw��A��ܩ*sgg��y�2��tV��|�n�dɛ�Z��~�qy�x��[��F�zHf��D�ט,���q7���*���Ş�-�Iڵ
=�z6v��:�J�zvu�g������2��:^�:���,vytol�������rɜ���a��f���Y��d|�������x�3-�:���d������v�v3׻3{�s���6]kL��{{�K6r!E��%n5諰�Bdv�j�γ�$>�d��A��;�K&�.ʽ}��t,��^*o���W ]��z�����z�{�2��d��]��f���L�e��vO���f�O{7nse]T/GZ��QU�Ӹ��;gU2g��=���;c[���~�7n������~`_IS�w��׺������1������_]\㼙�m7Z�v�7��{�:�G�Z��'r��?S=�c
'�!^͊�̳o��e�Y�⽳���34�m>Ǔ�l��������C-ܿ��l��,{��l��u�4-����!Nm�l)6CϢ�5��7����e�����L�=;���o�qd{f��ݧ�;*&���ݏl�Ӳb�_=��O�u�����2��m��vOL6�O]��f�⁆�U]{���ae�'jsfs%�㜓��_S���k߿@���UB�G�,�ʖ7w�/�:^\�s{n�W%��	�y9�1��/d7}�d��d����Sy���CwN�ٍE���Ѵi��n����w�P	��2y���Xz��N����'��:�:C���^����`���;��� ǘ�Kh߻���]����YqF���O�;��}��ݏ�&_>޸ϧ������o%�U����o��&+zw�2�s{G�7dnn�8�U����}�e��Nz�W���|�n���R�.p�Qu�M���d�]1�	�n���׋'K޾��ۺ�);#j�ۙҗ�t����w=�t����:��}{�g�(�߳={�nwT}�a�9�鬉��q2m���w'5��1�|�jܷ3_�o���?���Dj�0O��ꩽ�i�LPᵈ�OW�$}��(�}�>iW��?�h�Q�N�"�$���#*�4�fB
*;X����M�Z��'#�r	�r��־̕�v��lG>?�balM5X����T�Cjq��R���3��clv��A�%�"��@���q���-V����Z+��G-,�in³��j���2�͆�h��d�[Q3(�q�8��\u
�ꕊI�NԂ�[8I���$/��ԮpYj��(��+4����f��6X:SK6�[��kv�+�0���1fqd��i�W�;,T�4<�q�cu�����ĄW%�'�C^�m�,���u41KZ��(��G\�`i#3��r=�1��^����J·�ш#�U�ʻ��e6@��d�l��$
[eNTH���a��Q��kI�1bmZ��ܶ��I��Ա׵�1H�+�
�ecV>9FY��\!J버����*6�OW��Y#���
2JZ�m�ݔ]�mT�����i&J�jٲa�f�ˮ���ɺ�FPceU� �Rɕ�T<=�bBb�PMZ��F�rUTG"�ˉ��%U�Z����o[�����q�j[g�m�7J�e��j��Fһa��]b�[8s�d|̲(�9(^9-eZR��i�
W�5!�
��\��;+	A��wri6iH$u��9#�"$v��\ Tq:�p�u�dNڭ$#(�]i�����>y��(�2&@V�G#j�,v�IK���+���ơ�L���5�YqD4,	QP�\��2��[~Ʊ�1��.�q���7����� �m��w2!*�4�(B4PU	��e��-hU���RYRh	F�Jk�.4�1Z�L��h&
6XG1Q�e���%1�5c&HB9kR'n�U��
��R8�i*��r��9P��f�*/5�ݎ��� ���9N�ŐeGnIUUm�i2X�Mٻ�M�L���V*B�JI����4���j|��#0:���$/+u���r�<eF<11���j�Ty՗�v��m2�,pj;VJ4c��0x�9`�e,E��mJ�5b�ZR@�p��U�Ʌ����h&�x
�	y)j�$dq�Q�Ǖ�B"��>Y(�fbE�ٽ��oc���r[�m�['	������lMX��vX��K�7�:�3�\Zә�;$�l��n������ޙ���,�C�,�S� ���h̍H���Xیs��F4M��Z���Fx�O	_졕�u�vr���*�Y�"~�"kJ�u6�Hu�+���倰r�0Q��eU^C��k��
�CU1�$�$��\R��U�4EX������*��܁��ϑ;tTP�9¤��p������2�}��?����?���0;@�����-* T
�
������5�ۜ�9��$ 0 ��$ 0 @
 .@�0      p�  �  Ѐ 0	 � �`0 �   P`   0	 ( � �
  � mUP`@� h@ � XF:�XJʂ$��FDY"�!!2E 0IP�TP��
A!����1�a�
"��Y�g�+��I��D%�ɳCgs@0	  � 0	  Ѐ � �   ��  �          8`` �  8` `00	  �`  � 4  B 
 ,3�  p�  @  B ~J_̈́��`�##$"�d�� � �B 1�	*(0��XA ���b�Q�����H�i7�� ���       �  @  ,�$ 0 ,�
 ,@�4�� �   �  Ѐ�  �   �  �HX�    0 0	�d�   �  h�  @)/����$�k�D"�	c%H� A$�%I��* ��,դ�d�o��Yw��;5��    h0  � �   � �H �  � �
  � �
B�6�� p� �$ ,�$ 0   ��P �H`�  Ѐ���   X@�  i��}��J��HVE��f��2E�$"�0�J�V@=`MEdAHF �"�(Ȫ� !hh#��$�T�J�,�FpHL�D	@SL �
��B��J�
��+�
�*�A�o����آ� @��B�~������ xN�|���,}��O��F��4m�uN<�)��R�Ҕ��)��QJE)L)�)�)�)�y�]S�R��*yךq�Sμ�<���θ򔧔�S���<�e���L(�)JR�ڔ�2ҞR�JS
R�iJySn��u�:�\l�JaE)Ҕڔ�]R��l(�"�R)JiM)N)Jq�^y�^iN<�m���R�S���m:�G^R�S���R���:�z�h����6�:�<�<�[Sm0��imEQ����W2�ޘ���Z~��D����:D��v�ҫk����TRN���jRX2�v^z�c�+u��\e�#������'kDjʝ�pTT��c��!��<���>VE��HEY��\̋��ceq�	h��;�9�� �Wji;^s���P����uaŬ�K��ft��k\�MV�/-s�:�9 ���F봾��/%���d�Q
�1�;Y��$m�KS��d1�;%��p)*rJ��+
�b�e�h�6�"��U[S��6�\��m��K"�q��-2
0=�Zg�Z�,y	��U<L����q*�+wRY��棯4�%����*��+�U��!��b��9�1eQG��Q�N*�N�Y�Ze��N86�@D��셌n�aD�5%6���v�kh���s4�N�kOv����f&�g
�n)�SQ5ia(9ʫ����u���A��ܣn7mRY6�ͭ�eێ���E��ev�ԕ�[n��X�J�h�$qaB6�X��GRt�ǆ��*�Q�$s��N4�tE ݂�J5*j��Ĉ쉻ij��(�eW�$��"vY	:�#��V��fS9�7����I#ed��d�����K��v "�y78�pT�m5D�a��5=�n��XBP��<�:��׎��B«���R�R(�����5b���уDp��7�iߞ�   �
��<��}�� �`  ���%��%�0 =�� 8@UU_|���  =�� 8@UUI}��$��Z���奲��-J)Ja�4�[m�ab��]���ld��X�I
"�l�e�����nݒ�HU�k�$+F](����h�7��#����DH�6��[��n�V�3aᛷ���a,㱸���ZB��:ݑm�4l��M��]+aI�I_ %h8�E܈� q4�6q�Fe[��cb,d-���؈�MY0~����:�,�X����%i6��C!�L�(��M8jHBY�ՠ�X3�掛˝ѹUE�^�t��r����e��gr��4q>��`�V<yQO&��-~p�:�?G�&�n��K-�����1�t��\�?M�$�|���{�:t;<�S���6�=iig���ym<��
a~QJS�L2�8S��6�
Aط
K[�&Ly�UB��lɩ���uXa��;W���4�G�����jX�zCGgg�A�����<9mj��d�QEATtEvy��������ľ�t�H�}�p̓�9`"LI8�6�\żG?#��RKl��)0�C��g��7|�Lq30�:k�����s
�{�'C�C)��iL�ì"�(�)�4��M�4%6a��/��/U�7pUU2�Qٸfc��s1ː�Y�h�D�`�uC̿}�3)���Nw�{\��ӘhW�"�Q�:�KI7v��R�wGv���f*�V/Ӷh�"d��~>33١<��`�!��y(d�Ύ���L���0p<46zVkыt�i�GI�`��	����[/0�E)JS
i�0�(�j#��A��h��K_� O�/,S�FC�-�Ap�Bq��
�9l�9��;KĐu�ݭ#[VVX����K�ri�\�9���-��|{�4l�S�a��6�jVкt���,�p�F�C��g$"��쑜��R�a�\6ZnNwFMs3j�F�.�!SC��ԑ�/�c�A�l�s��U�ܷ#���&�ԧOF���}mm4�/0���������z'A8Ra輭|ޅ�8��܄�m��O28'�̍�Ν���py��J��B�'��)���<y]�F<u�.K�#���,�ҫ\�6��{���;QE	(�e
�.Z��*$qD>6��s�:�e�E��n���g�oy�� �Lr�cN�pb�!���I#��D ���Vq}ϸ	ɞl���+��F6M��yy=T�ɪs��94{��i}[�h�K�ٷ�s2$:FG7�*������x��@�o	�vu���6���!aӰ�׼2|Of�kKU
1�|�n5�47םD�̼j�my9�q�M��n!�s��!��ts������`�ː��FK(����R�SJF[F�e�*���ms�-B�̥)着�K	f��p��&ܖ4�%T����&���~W!��g�^��92y7$��l�!�ӣ`�><�oҖ�q���ޖ�mb7!}�0�_i3-,��8Z[��Ёp@���q6#�Ta���}0�a�f_I�c$Un�x��C���&	bn�C�_I�� ����uƛe��<YJE)�2ґ��Fe3�����ћҪ��p���{7�R�2����d���}��b)��d8�0���[R�\�l:�����9�A�p��.K������Ķ֍F�͌W9�w�Ҹ�Ç*����=�c���t�JN=,����F�8i�5j��9("!��^<�r��Sg��nY�Xy��hY�������i�y��G�R�����iHp�O{��Ib��{���*:��9⪡M���
��\�\<�7<g��F.��jJ�[�h��ң�����a��D����y��b����s蝇guc'�Y�K5��h�w�m��pO�i�p�0=��X�1lCa�;~h�Sf�K�%���^�	����.��pi2Xɓ'(���R)L��6m����g��(��ƾ��
�l��A�[R���B�4E�y�xbNG6�;�8�$����N#�V��RX��v�JB�X������VS�rj^p��*n��\8���\�-�ԑ��{"9��Z��(���ܷ,�rB�H��V�UQ�� ʅ,��,���h��X�eҴ��OO�܌2g&������N0QW�0�y��N�Q����c6�%��R`0`����ҩ�R�D�a���zup�_V�O3�C�AX���s����z0x�ߎ��wJ�������0>�OU��rrffepcr3-e�#F�h�rK���q"��� N����T���4n%a:��t��:�:�YjR)L�M�mm���gӁ����	��@ ����G2)�x�%�r2QA�����K��4yt-�*(�:q��]�L&�JL&[��h�3U*U�l��IϨxs��z��ے��A��+W1��C�������//&�<U;��;>&�0�䏱F���w���ɫ����l5056y7�E��A|�k�6�8�����rHl�I�!�l��O%%#���)�m�2�"[�̶--�6��'Vͥ��N3�f--�.I����Z4�In1h��"�Ө�Xi<�\�aiII���Ih�u<�G���쟑�>�:�y��O�ɲ��(��+�����������L'Qķ�e,��0�--�-�:�--<�J[��,�Z[6��e�E���o1IrFƐ�->�)JC�b)�JS-lZZq-�--lq--Ly-�,���KKi�E��ih��%�Vť%�R��--���R8�%1�)�S�hq)8��I�nL0�->��q-�E��L"Ғ�b���bu�m,��8�%�Ţ�b׉lqlZyx�Ғ���ުp��c��S���D��<���Ϣ�,N	�?g2J��=�����n$���{S�1�/2�v��������w:��ޟ{�Ͱ�牞��qv�|�#��qY�;-��oL�S�}�ޜ�F�1��l����#Ũ�w�b�A��|Ysd���ؖI��6��dɊ�}���'�2.������kq>A���q��Y���L��`��ʤ����Rv.��)�Jw=��4���ϋ���uvde��#Gsu;����+�7	��1b��M|7�oFr�汮{�!�r���^������ � L̞m}��wtwww�w������fd�_$��;����������������.������=�{��y{�32{䇞q�e�aYJE)�2���㣄)N�&A�S�EEED�h�,<�z0��CΟV�;�@�:$`�5����	��,&0I���{�:d��R���B�DR��0��2K��q��A�k�.~���c�i��[Qݛx��iEV���]b4R噋C聟k�Q��[5��*$S�:SIM+��B�X��lC$ Aw8@����!��la�CPCM;˙MHjYP����H�)���ؑ���������?@,E�i�0'Z$M�(k��=���y��[��,��x�����	�	�EF)���-������p'�$����^�0� �I$(\�Z@.�ǩ!>g���rI�!��~ʙV�����ЭLg,�tmʋ1%� ��'�ᴤ5�[�K�h.�d�	��|l�nP޵�@��Ҩp���jI,`"�H�.��A����!��!�����Q�g�4a�!���<?5@F��R܁h�"���!,Aݭ�%�D,H{�|xl��A��'㒆�a��/��.�AP�Eh�y m"��z�g�BO��>ï8�L:��G┊S*eM�mm��.4�0Wq�l�m�bG[��e�帥uH27Y����e��n��n�KI?e�a��uE5�37"*��DCۘ��]5kLZ��ǆِ�w6��̑tG]%��-n天m�qa4���OQQQQ#7\6[a۩� ��6��ɻSk�9M$x�ksp9������Sġ���("�� ]!�#��%J���OMt�����<�u�=M!���+�DWdp���!	'��.	�e"�:�`���^�B�Ԫ!sŀ�O ZP����` exFP�N��0E�1�@{�0j�6K7H"�{$�}�x����"� ��"O��r���׭O��a�H��m�H�*vZ��mQ�൲l�nZ�k�h�ɐ����
c�<�r�"4S�@�rÑ$�����H.�&�"6��e�����?�)D���i���tG���VSM����PC �{C�'�D��vO8���<�He:�Il�$� ]"6�` \�X��"5�HP� �8Sv���TQ�Zօ�]�@���Jm B�I0�6l��$���gݘh�@��[c�F�����~��{�0��$x��
_@�Er��]$�J0�4���t��ѓ��*g2ō[�ILn�xM�ʃ]��}��2C䌜,'��F�	{8d���(,W����fB��9 �E���_Є?1|}��W��|T8�P!�����D@��+Z��z
�x�t�5�R�E�2��)�Y��"�ʔ٦�[�4��d�ܶ>���"�Eb�S�q}EEED g�`u�ܘ��&	��������`,~��prR�g�Ӝ��� �'���dԀ�F��u*���`�� RA��	��z�n�&�4'�	�5�ƦCB`!���d�2I�$_T�<!����H�[r�l�m�ilvm��;[��+�4H2iv�G�Q�"�"(Sr`Ce)��Gb�ؽHH�Hh�������Y��-�Q������6�!7�)�42lB�MC&�d@�!�ȥ�b��!���//{^�0a��Fb�NJl �-$��B��B�10�����G�CIa`v�Y!��`Q'��p٧T����?�JR�4�Ka����+�C�z����[�i��rE0�甶���P``��̧R�兢� y�#X`"%B�
0�:C�\i!���z:���M�2ԐQب���!,��cS��,���U�l8��wn�88@����=���E�@�)��SE�6���?y��s1�1�1Y����D��\'�X�Sߐ<���D��ivl��082�nRQDO"�}i�B�S��:$��idP��N����6�#�%�ujH�ՑҰ3ݍUZ.�a8�:�����L��d,@��@x��]F!L.E/��X�0�(��>JC_C�{�9�k�#�uM��8��,�R�JS
h�m"�q�r�~�����\}��h�F�co�+FPPTv��\V>�u��k�������,/��Ah�|��
䪷m� �Z��8sG#<�ST�G푨��%�C�JU����n.�mF�$ݙ7!�FZI�u��TTTB�L��d�:KY[��1�PF
�F�E��]	�uA�
gxw���3�W���@�H��R��و~a�IOb�#�Xd�F( �}�����^�ì����y�5'`��:����y�ü����%S�!�,/�m"l�!�P�8
���E�p�0��}=V����jѲ����b�>6�7sBh�k����l܉
2!����a�c	�ʔ�dg�A���GGĵ	����V�EP�U*�ŊҪ����Ʀs�m�zBC��т���
a7X
Q��q43��cn�7�!쇜iN��y��)L)�6i�>8p���>�j�ְ�֕�t�;�������{$�oy�����f`��J�C��s0a���=�����< y0S�LU���x6|��8HI��Њ�FSeݐ��85b�Ixn��7�*��&���CP	�n���2曛 o�W�d5�q"��6��ie���٦�X�ˆ��'K��C��<$��B!� �d7S���0�|t��o	��18L�|5��M��Q5'AA��;�rZJ���9d�H['W�No�-�yl-����)H�2�T٦Q���ϷOLȎ�k�Fw��[KiF �~�2+��M�w�P�����WP��jr{;����]a�̛�!�Ac�Ԛ�
�e�@2�<�b�i(���gK��3H@�}�dy���Y��6�BƘ0�Ҧ�-a^�')w
f�8e�H��l�ۧZNK�I��'�'�Ղ�ZՄ�y؉��jr�>=�O6��'Cr������0��e.��$d.�})<WL�a���VsÇ����!M��{ӆ�N�G�B֦���<K^ϋ$��h��4h���h�R�JS
i�m�en4��r��kl�sT��9�jN%�����cP@"cRRx�0t���o�xj��@&�&�;�hiOi=��&�g���
���f茨3*�f�$u��ns	sa��6��&�x~��G�n����re6�h����h�[Xf��*�p�ߐ�l+<a(�(d2,_�. ��}kZ�b1]{I�覙��h��Z��DO�Խ2}ɫl���B������0�w�r	���` t��w�<Y[Q̚�OD���bl�"�Z.���r}�XnH�l}i��aI���~E"ґkb��JSٝb����K̶0�--�-�0�:�--lRrL�d����[L-�-KE�Ţ�Ӊii�T�b��������uKO��%�'�M1�--)��JG��y�#�&S[�����Zy>��yl<��O��y�:�����~~c�~e��m�kb��iii��R��Y<�>�e�--4��������Kb��I�����Z??0��Z:�&��1����M/3�b�b��s3�ZZy�--lS�2�KKa�KF�am���Zql-[)�L%%�����Kc�%���KN�������RG��JM'iIԩ=�<���&����<��Vŵ�lZT�c�1iiKe�L�iť���b�űijĖ����[-�'�L��K"��ZI"�"�䴉R[FQ��W�O{��c����*��'�t<�p~�l���{S��8�mM.bx��ty�:��^�"^�*�{�����G���k Țo���c�X��]�����"�33z�@�KLvy��W�m^GO{;��a��4�hj���;PgvNj�H9K�J�bo�j�(�ֳ�0�Ⱥ�U|�of�[��s;�� ��(����������ŵ��0'l���<�+l���To!	�"�2�u�"b��4�Fмb׆Gi�C�Ec[�E��״c�|�wT���l5ڣOt�1f@��b����Ū�X�z��Fe�#�;��o>���� ���w5<�K�N������'�>�^����Qf�� �E�q鮨(T�}qa�ob�L�]̆;���p��ط)���N�jk�Q�����Fs�����Pgf*�΅a���^F8�;ﮬ����=U�h��d�h�$�מD��ϫ_]W�_��c'�
�����m����o�s��l�N�\���w=���Ե��%���:�ݶ�A������V�v-p=*��c�;�������%D0�UE�ƭ��9%�ʥ��#}2����ID,ʃ��(�!Q�U��BJ���Q>V��c��|���ɵ�2*ꯔQ[��s&	�$v͌!��J�4��[H��X��-U��E!�U�ۊ�Ƨ,��]ad!	vR�ZU�u�x����d�����#O��r�yy*Sm�k4�J���#l%n�*�Lt���)8"4T;��"���х�E�����7�7%�NT�����6��M}��ߞ�� {��y{����任�����  =����陟r]��]��X��{ީ��}�������H `3���ϯ�V��˗6�0���H�)�4�6�2�-Uy!�q@㟡lCUҁrf9H�,�����Z�&�)|���	�cu��pN[,�����g7���)b#w6;7"����;�Ǎ6�Q�&dlv++-n��)kq�mrXI��0��tnIk�,����`,�ɍ8Gj>�F1�cHH�f��� �#+�ʈ��Uk���B�SRB�Y> ])��d�m�FB)Z�&I��F���%�?�����	���,/�ِ�2��¶}�P�UC(]<.�͔\ xN�<^��x�̛+�h�q�]ˊ4CA�D�&\�8����Ƙ	
 ]"l9��p�N�K5�����*��`ĳ�:d,<��L=���~_sD���'_
�JK%��2�;bpF�jm-�&��!���t��a��p����T�J<q��UU7$t_��)N)��"���R�S*m�m�en<��s�9��z�[��Ƶ�kR�	蟤�l�vd�Ia����+(s�U�r�3�<dH��B���a�L��1cEg���1):r�Ц!�B�&&Ҏ⓵I��Q��������<!��&�vK���t� aN
����jh��`���C����ꤍM���I2Y�i2l�!Fp8rg#�U˸ny�s��nS�S��>�݇J���S��$:�i/�eӍ��`�{�Yq6��������K?c�ܩ�5|�sRR\�K2\�s&�p��oŭ�Tʛmi[�i��D+��r�a�En&�c �mNi�Zֵ�D=�r��,����MÐ�q~�̡��e�U}K��@�!�$�e�x�L��A���c�!؅��e͖��+ѓO,���:X ����,ԓ,ʂ<~���ׇ�u�S�ל�K_���tݳ2��������M9b<�Y�1Uj��̤4i6�w��C��<-��|�Ž�CI�Z�(�3	�l�-�:G)������M�p\������S�C�u����5��0��q��VC���2���F�Ȃ�����<s4�J?f@�]H�b1FL,d��~E��Z�Sf�F�⾤s}��>s�?5�kZ�A�w�]�z~0��#0�!�ZB`Řh;f�wS
S�̟B�q���O�U��H¼�Qu��+�]f��q�y���Zg�F<*y:�"G1!ޒ]n�v���$��J�D 6S���Y�e�0F)��l F��s�BK��ĳN�×0e�l t���,�u4f�,�A��q<�`~e��Y�1��4$�a�4�C�0�,�N�aK�Rִ������G�l�b[K,:��i��S��[�YkE��)�-�kq��\�ZDzOa&RLaZ�z�B��� p��n 6����D ��6��<�1��5��R� �L[�	l�w��_n�t�d�k�y��Vf��hQQIEkDiȭo(�Tj���X1K��M[�F�]6ڷJݖ5U-�� �h��C=J1�c�BNfmp�dV�DF����K�R�n�!�		9���~�
�6Q�&�Ip���$L�����jL�sPd��h*A����Y wё�{��q��e9!�>����!�;�(��z�It�}�:N$(�"ܲR؆�&B�xbH\���y�<�X�� [�6$(�IĪ$2�8Z��[��A2�R�Τ�M��DڞJ^!�#r��]�rꧺ['b]Y6h����0kl�3��k,jhi����t$Pmu���K�J0`^K��æ�aA60�!��i!��C�,��(�
YY��*��V���2�M<�(��?�Z-L�E�Ī�X�-]�B�a�MZֵ(0�=0�0�g?F4t�2'��Y<F�ϳ0��s>�������p5�6�<-��Ot�� d��;V��.Q�G#UEA��'��Y.��`(�x'��6t	�J2k�`y��P��.K�~�:&D�bz���tX2	�0�!�?OE��o�,9i97a6��&���ђ�,,��s�<Jh��$2�$2L����T�F�UjY,�O��}"nP"F���z���s��OWd�I��@���\wR���m��q�ʍ�մ��~a��[�kE��2�b�,U
*a�� �#�U��F2��J$
2z����+�6���Q&�6A50aa�A�pMa�"jL;.̤.!�(!��i��gt=-ޏ��3�u����x�УK�����Ce�YZY�ׂ�����<�xb8L��0؉�50�!���<�t�9����dX�g�5���ς�\����%JpY2�ѵ��&�����#m��p���dC!�
4S��Ry!�+�ÕR��Hl �c��n#�&#]d\�影�>}2�.����?0�~-h||SҞ�)d�9��	�gJ�g2Q�R�*��1�M!%�Hy���?���M�k����z	�MC�Phd9�?A`!�W�4�s+sz�&<�a�q屓35,���-w��d2c�M\$�(�t�8�0�`l�dbXɳ����ѥ��0�.b�d++w���@�r�^��f4��n~!hO��!p��B����u��1�J�[z�tރͣAd��D�Ԇ��2Q��A��R�H�]C�O��S��.�r�=�"]�Oaw����f�)�:�*[o̿0������ʔ�Qb,��~YYL��d$t��*(��ϬXёddM�?��\ta����;s�r@O>GonV��+ƭ7{�o]�U�a��+q�[Tm[,�JH[U,*e�һj� ������*�,p�Z�@(��)��JԢD"hM��~�1�M	j�V��1
��Ԅ��lel�e����.����assgg����~ɽ���@�t�K�/�G{�*T+~������c7(��y"P`#�
eO!�YfB�=��Y��5��pJ�9L	�n�1��#�2��x�\���!��:�^STv�%�2d�n]�L�E�PLrz�f�Kt x}���X̩RQ�"a�ȅ�!AA�Bx>���ID���w��m���*`�j�Ҋ�D�#V:�3�u�5���z��d:�͞��K>)A��Dg ��<�4���4�����4���.8Ҝe��#��kE��2��2���kMgDξ̄ģ]��>�c�1�0E�xZ1)ѻfI)8�	c@�0�a���h
v0�C�Cɐ�d�Ӊĳ���ѐ�pj�ͧ��2�Jq�)K�����ΓG�n'HhL�¹�B�<;���7L�K�rC;0�K�!A�JNǦ!aћ�LɰC������j��l��&�����e��=�	����Ԥ�nlQV1��Ô���21?{@�%�X|_�q�����0��pX���4$(���
nCT@�'Oߋʘ%�29��.N�fN�m�zW-�� ���KO��QH�u:��b[�KK^%�����י�-:�--j��K%�KKK�-�-[q���ӋĖ�JG�H�8�T�JM��|3�8=	��|���
�-L-�c�&���Ғ�ғ�i��Ǒm��Xq2�ɜ���iiiim-�KN��K[
~c���"~}?%��e0���i?%����KG��a�u[̭8���J���:�M%��[6�����[�i�E�l�2�KKal�4�Km��ӫb�KG���JKK[S,Z~E�0�����'��X����\T؟���O��M���є��,Z�)�JVe1��y--X��8KH�-x�[6�N-�KV%�E%����L8�8��)Ix�E��>���-"ZD�$KHg�fw����)�~�o;���_�N�_���n��#~��j��3>�����֏=�X�ְYr|���A۷�����s�y�vNtK�Iu�d5��<�H�f/_}G�gSΓ�����q��E�M����_=��i��*���F�_�'�Tw���ϳ1�]�_�O�?(???,@�몯Z�����z�$ 0����ww_w�@ ]Uz�����z�
 ,
��z�ؚ��.i�[y�^a�֋[*eM�dM��}�q�>^5�kZ��z],�n��H��U�UM�ۃ$�D��L2xd;�ê܁���M��@D:<C;$�cI'_%��.^�<y���:�kJlhk�Xs�y����G)�5 �v5Ur1B�� �/�9�1�,%JJl`�,�!�؁DO$|��p�7��`�H3�9H�2)~������/��L,8G����]���B�c�rB�a.����H����&�(��->�̔������%��L[�1�:lÎ��6�
Z?Zֶ�̶&ƻY��(WN�R�9��iSI�������(!�`tN���6�s'SU��~C��B`�}�Ul���NFN�&�yd�4 ou;�V�)WK�֥����`�N��&!pxR��,X�[ñ�,����UX�E:D.B�F�L)�A`�b��1]
񙙕[3�����XVEa�ɚ>4x{�`�D)��ō�g�#�t�M.m,�b�7$���
l64т.��aN��F�>��(����$.]��N��i,�A�ioբ4��rRE�R%�X�<B�M�)~-h���6e�o�c�c��?o�|W��!T��)^L� �ƌU����Ņ1�`Y�LUfO^M�|tv�����Rܲ�"0�9�&<��1`ev��)!B(Z�@�콭K��DI���Yji�1Աe���v]�I��r�v(�J�Wf*�v�{y�9�e�Ғ���TTW�s��4"�J��)F�C�H2֙crKl�@%F38p�>8���],�'�M����>�/'C7L�p�*Y)��:���@�˥қ�c�N�Q`�c��j5��$rX�q��Nܒ�s�p<���u���Cd]�I��\�!��	���,�9%ސ��HRfŽ	�ݥ.#��K�ɺ����f�O;,b�!��u8�!,Q5�	����C�%&��Ɣ����Y��[Sm�k6�+A�n�v�%%���p�����C�a����ynyC�����2�p�bi!t�L��H�XQ��i��Ű�~-h����e�o�9������'\vYd���QQQ\(!�e=�W Q?l�$a�8|aD<1�n�ܓ y���l!�m/�62��v�7�%Qb�un\�����݅��,ā�"��񆋥8��e�h�B�X0"��X���a���W����[�g��P[R�$hM;�p��{1,&aa��t�.�J,�.f.Q�e���U&��A,�ڮ��#㴺�I]x؄<�),{]��HZ�0bX�G�:�1M�Ѣ��<`�S���Z�kel��L�n{�<rȢThWd����99���>�im-��Q5�K'�80Da�9$���l-ۤ�y�؇D7�nb���Pp��d�&�U0�C��8��`�����+�#�t���51����Ȱ��+nܻ����e��'��A����(�)me�i	�K��[DZ��g�~�Oe�;5��U��<(�2.K����Ԫ��ΎC���'���vd��[n��G���V ~�(��m* �OM����0�;ۃӰ��d�>�P�Xrt���&�r�`��2�!s�|t�E1�D�m�a�~^X�#M0ӎ<���8��ŭ�V�̶��q�"c��_�QQQ\�x#��}���9�fk0�8I�0t��}2t�B����C����A>:�g��o��6���Y`ۖ��:�u�^ͅM��G&K�V�z�ǋu�b���Z{Rz!��BNl�<�@�=Eb��y�����Н�8t<V8w!`�""|z�%'�l��:s5$*n�!A���O�xgF�5�o�5)�L(t�g�MC���m��9
n�M�ŪSat�f�m��*�0Q��2q~m���kE����-�lg��v�6
((i����D�1��`XS��'Xp�+��y��d�cO�,r��Q��WҔ�2En�X�F')`)YU��e|u��	FT�V����F��d�~�QQ\�7�:�$WV�۷*l&��n�܅\�1�P�L/��i�]/���s�O�E74{,������7gg!���D8D�D���=n�B�l��� �ÌFk�Zz0����d%�&�^zu�CĢVӸ^5Iɣn<��L�J
n������[�rv~�&�؟���"a����_M���=�p��z������5-A]��;c�VY@%s�j8iY�������a���PHa�
M���Z�nO�72�N�2��4�/6�?0���Z�kd���a�6}���*Yi���ɌȱF`ʍ��b*�%B��p�y�[Kim���}hf�(��&ƨ�d�����d9�ɓ�z�A= ��<ÿ�nP�a���>̕.օ���;6'�nY���!��XJd6��%ŗyd���T�K��2]�l��<����!��3ò�!	���b���l���ӈ]blA����ü�x\<S2D�Ԡ�
#Ě̛�e8x<z�]�
 5N:K'u�W)��!���#-��-m{���;�w�����D�W�0ӌ��Ͷ�QjFߖZ�kel��L�i#,a�L"wn�{��	�ft�̆��͞f�Z֝7�
	a��|�(�B6�ek�R�I�m���(��F�!��*#��'|<d,!�L�.�:<= 10����c�>���rX�2-+)Hէ��cX��5%�&�HQ���7�7��NL��CBy�B�жS�O����K7in|G�<�HG�(�fr�ٳ�Ce˖z�C���V�|=NON�z25U%BY������є��G=����U~)�p��0��29�>�~~y�F�ml����#o��Z�kekl�h�]���q1�Zb>����$f2W3Z3ta�$�_��-���±)����}��l�}'n����Z2Ra`d!�֯�	�;dU���* E\ᇩ;z�vD�t�rF�Q��d;��2�V����%��g�e�N�@���h����'\�8ʞ*�����Ht�d�ɍ0�Rz~=���.��w��޶��-1l���!)[���0x�],e���0�f�H��&B�8扇������|N�m2�B�iI���}���O�H��]�-�R٤�qlm�K1ii���יų���ص�Z��e,��Ih��\�m�G���->����Zy)<��T��l--lZ0��JG�ObE'���$�ZZR-)��"�a�1�R��Kc�M%��KO%�'������an��mm����ZZ--L[lZR[�ZZ��6�E��-��œ)h��ZZZ-�-KKO%%����[�����E��iĶضX�Z8�-�-lo��KOZb�Ɨ����?����R~F��q?'�ulZ<��%%�����Ċ[%���>�Zu*I�rHܒ=�E�.L����KJ�m�)-$��aly��~o�f-�O'�����[--��[�����%�-��-�-'d�$�8��R���d_�E�O��H������ե���z�+���7+^9uo^ߣ]�;4y7'������,�d�~[}�S�_���78����tC�l�=��&_j��vd2�#�����?���ݞ��0�����z\��w���|��}��N�E�~���YP�m�l׎�yۿN2�S�=���+�9c�1ʄ�9���H��j瞍�z�8l�� 휖8l�Y�Y��Z����O1kh�s �����u�7�{�w��QBs(����RQ0�-˭-�	��������iI�W�'0!�m��>�|e�۬f'9j̹�7z�S]o8X�(�
U��I�Tf]��8нP���?]�b���B�+��"\��k��,S��u�ѻ���ٗ>*�(ta�:��o6դ��#;r\�:5~kcZ��/q���k��|=Ӡ�[>��_H�ca3׉�vw�o}��8���������y>���Ϫ�f�}�f;V���s.d���'��TW5�b�$���#B�>��M�揱o^\j��5������M��2���oWN����Ssdc��M�O���&�W�l�_W�Ǜ#F�^�Zq����Y�:�5���i_��L�y��k"7ÌP�\ˈڷT�z�a���v�`z<��X���=��k[��;-��F�ʣt��EST$�� �EV�]��ie͊���7Fn�r��r��24�"��T\&Q�Jƈ��� N?I�	�0#�L�KF�S�f��RتVH��2��n�NJ�Q���U٣���7"�E,�RZI��M�U��vĤ&��J���G��t%J �m0|�*u5�B::����2��ɌC�RĪabE,��v��P{ܱw.��F�\ �J��\dYaTuUQ3UJ��S~Ɉn:�oǽ@ z�]�����P@�^��Wwwu�{� P`@Uz�������� X�^���˗-\�r�֮MR�YkE����-�i�bc?Tְ�9	��:弄��J�8KU�]i��m�t��"�lmm��@��4Dƫ,dR0��ye�n���7uv��[��5$ݣ�#��*�*�@���c+��v��򢢢�!nq���I��Z78kX�,�D9'�~���'��~�B1<�4F
l����`*s�n�vr����Й1��[Fѡ�t{Jnnt��[8���ǣm�_��Za�8�#��d;�������ÁA�|w�r���/�&
'�F��}8d2�a��^�W�W��-ц�[�	UU��Q1�"h� | Q4��I�d4��tN`�ph��?C��<�'����q֞��)�Y[����S��ִZ�Z�"�,[ï���2b��S�JW-�K�s�_>R�[Kl��'b}8�9��`�	���_���z{�_ъ�s8��N�&�e�'S�
����y: �������K�SfO�@�So�`�1F�b�����8q=�,p�����>�sp�x0O9����a��m�7j���Dw@ܚ���f��Ѫ����D���������:���S��9�<�0Bɺ����Δ�z��r�Ѵ\nt�t����92"��8cm4��y�[�)��֋[+elJ������!�s�l��0j��}Kim-�������֎C�X���'��\8rC��	��S�ET���>"$%a��_4m2�}�0�i��z4!u��	���5�������1Œ��91���JA�����%�%m����.��:��;:��B'aD�QU���4h�X!����7��LcbIt��SSsÂy
X&����~�\�Έ�������|�KES���T�:��5��s�����e�V���u�0��ߋZ-l�m�msL�}�ڱ��sQQQ\�r`�W�I_u���S.�祹�6m~=8l���h�tlL�}�����J�iT�J@�!�9"$rYGy�\4ي�r�8tᣃ�0O�������m<=?O
`lD��lɷ�%̐�˒�w&��U[�L��K���C�ː�
�=c	�.B
JOcF�Bɐ�4s��E���{�GX\Ej����I�g�!��܎�ߘ��B{��L<�N4ی��G�k-h����e�m�ԝ��X^�-v�NG��kM�]Q�Sn�]ėl��:L��|�s��cMrZ��G%�U����^ب�ad��kr�vVfcX��R�D	�`�lH�ʯC"�2T��%`��p�"������S���&�J��jȂ���Y����TTWzQR��UŬ�iY*[-B1��`�&)w�%��$т`����(�������.e����P�ٸhDF��G�\�bU��p�� �'��@�Q=��5�0i��ScDZ,D���rϣ%0�B��L�Nǆ9%�,��x�����铇�
&I��ʍ��Û��-#��B{=��k%m,n�c�X��(��z�	j%W��E�wiŹ��e���QI���37�����Ka��mM�ˬ)�[k-h����e�m1$D�a&������7�M7��**+�C���=<�s�����bᓵF%U��H�2��C�������x�rS@g8xd8"��C�S�e��J��
''�Ӥ:~�����+��k���QsBzp��R�q�԰aH]�SR!6�
�ln�,�Aʉx�F�V�T��	�~��N��ۤ�u.CĜvQ�&B�K�6����$8L��(��6�����ͬޜ�0`��Jq�R)��֋[+em�e4y���Ȣ�'��-�����9c��==+w=���qV�
�8"C�O%˗�Re<`,C���ɓ����4B3u$�/�P����������e�)��l$����UPElB�QK �k��^�r�k���E%���W��=7ٹ�8	�!���d;���ĳ=�̧�X,B'��>�q;�ѓL(�պ��UUQ����8�8h�t�=,�z�y���B��<M$	y�81�]�g�g0���q�����ִZ�Z�2�6Ģ[m�[i�1�**�Fd{r���[aD��?la�"*��d8SD�����8J%�7�j�4�B;eEv w(�q�dfn��i]wm�\��CG�C�Ϥ��m�b�i�	���B�������e�3i�&L��v�R�����uy ��%���ѳ.5ڨ:��,Z�.���6!�Ƀ��CAj
�\'[�ah��k&���6�5���_<��i��q�u�Y��֋[+em�eq�f����k��͠�eD�m��&��|kr�Q���5)&7��Ib��)˷��6Z�T�iT��<��.��2::�mmW���P�j�B0M�s.A�T�Dj������wQ�z����$�.26�N1HڡI,�[v��UvX�8��5@)t���4�ԷL��,�C�d��g�ҎE)��g4&���h�p��Q�h8'n�s&�2��{	:q:l���8�M�2]�S���4�Up0MrS�= �(�!�S���^c�O'��҉ɇ�{�N��Y�Cb'آ~��#�[NJeݹ.B�I#�Z�)��jt�|rv
cļ�t�V�����8\�Ҍ�l���֋[+[l�l6�����5�Ӟ!͌ɮ&��c����"��y�TTW�;;�pc�?w��h��Z
&�t�Z��%�<4�0çN�Cb^,��5�K{���U�w�=��ss$���蝂~�O��,u,�JK��k��0��$�s-R�ӆ��˓D!�0m���O��Fd��V�5����il֊��?Y'a��>3N�T�}("2����f��:��:p8!����0�>П�Ƹ�i�p��<���{��?O��ZSOζ���)JQJS
R�QJyJqM"�R)L��4�:��jS�:�y�^:�q�q�)�\u�T��m�uO)O:�T�mM��QFԦ�ʛS�uO)N3R}E)�"��)�)���ju�4�]y��ʔ�)JR��)JuJuM�R�q�)�4ڔ��yה���SΩ��-��aխn4���]i�\R�Z�ee��4�)�)�)JuGSm0��(��(���I�y�zU����wv�&�[��=�ɯ1�K�[ar�ޫR��w6t쌬�s�dt���.�*�ϟJ�S�7 ����zn�we��Z��ک�5�׼��0�=Xz\d{~��+��ɺ����s.D|��y�����ܕ�f��]r�қK���7�Yj�/*!E���P8����'�j�;oh�����FeWwnIue��+����P�^���wwvw� `%Uz���ݝ�H X IU^�Gwwwg{� @UW�إb�ʗ4�<��"��-h���V�HQ8��{�QQ\'�p{�� N�4��_��0D�9#�HJN�Âw�ѡ��C}|oi�q��ی2x�CW�v��2d��q{���kd%e�-��e#E$�l�ؔ��f��S&|S�X�
��C��CG����KL�827�!R�|�0h.Ci�AGK�����{Gg�)��e��C��q(��]�b%�I��`ǳ�\�ۙ0�A�;��h�BmP�J���Dy��̿6��q��"�ͭh�����6�oq��"��cùg�i���**+�C�)M�͝�)ᢍ0�4CIGz�i��$G*��#��iJ�t�6�n)�qF��&�Ό�f����{�8��]6L�/�i�Ibɖ䱾��a!��ے�UƎ'��׉�h�`��a��	Z�|��/�ڥ43���s��%Va�����L�%�7Cϩ+*Q�x��hD���c��
g���H7�m8�m8Ҙy�^e��Z�kel����8<�Ɵ1�6J�Φ�x������ޜՎ�vo^�f:	�vs�f�X���!��蹐i���H4$�Z���v�Ց��q��6E�����ik�i��1��S�PB��6��6Q�%��,Rdw(�hD�)�
���p�:�m*+�C����zm�wk���V�+[+T"��2�䶗����Nð��T�2'C��ڨ�_�'�<���o����fː�j/��Mo�a���`T8�tѨXh�>��Uۙq�~U�5�J)��4�6٦j$&�pɥY�0�O���l���٤gNIÆ�C��}�Z�~�5�9��ޢl����aY�7J,�!	9�}�<L'%��a4��E{a�I�B�:�U:��l�zp�E6~<oμ�?6�Z-l�m���ڛ�D��;Kim-���<����� �N�x	�\�����*�\��H�0��Iŋ&R�q�;��V����9�i	8hB��PNO�'C���Q���[[�����:�Ol��3*��X�2y�h�<<=)�L�~����Jl��v��ќ!g�	#�4DC�|��L����g%nX����7wNp�8y).X:h�l0B�L���.Z�"�u�}���N��WϚi��i֞a�YS(��kZZ[+im����jv�C�L�kTҰ�J3)d&0^A�C�E�N9MP���**+�t\��K;���'Xp:(&�'��<i6�"i�3A��5ډZ&aOa�a�xp�4rS��܄[Fֲ%~�����uh��e�%��i[ �]7i�,����p�_SF+����8�p�p���2_���b0��K��yΞ1�!���{��Y~á���N%j]�S��$*d��s	��݀e���I"�i�?}m8�-??0묿2�[h�������6�kmX�d>���R�f���������������]]7Y]j�nT��t��p�I;p��S)�M��/�*zK^Z�ԥ���7X�lk&$H2h�u,�0T�QwM�iW������N�6��sI���R�X"u�X��l�	�����Ռ��2o����=��t��j2Rb�]!O�y0n�8X�̦�0d��8�ߖ~m�����Ѷk(�s�&��)��$t���H񘫙s��cͮ	�Ƙ�	�Ѩ��|W9� �y\�ֶh�KԞ<lX�c�M�ed7�wbݚ��33yY�����D�P�B ��bq�2��)Z���*-MB�V2
G��e�[������CvM7kJBl6�y�H���	�7v�	�-�:�u�D�j��n(�-eQ��BvF��t 8=0B<m�Hm7]t��20� �4C��� \��K-�h�\�nu�X��I���4�(��li6�\��X��0h�Zħ������Qd��:`�R0�\��ɐ|�},������46t�|1[S}v�+��)eI&\Iv�R���83ǩ�&���r��&4Y��^�jL|���|��u�4�8��??4�������6�n�s��}0�0E����[Kl��PHrj7�5��I�>�fe�ΟqA�Ԯ&[%NԪ���c��r�N�d�xq|e-���ɳ4�E�Fi5�Q�Q�l��a���e
t�I�fy�J�V�I��E0Ca2f�$t$̳fY76�a\�����ӕJ3�,=�N���F>��<�	N�T����O!��!�rlD��>�Կ���c�=����q��SM8�:�T�,�KZ�Y��N��9�I,��f��u�TTW���~:�s7��3���¥�0Q�8�4�L:B:x�d�jJ%`綅��L�I��ZR�]8x/�O+�ܣX�P�3,�FҚ�C�:}��51Qf�L��|f���f��.��9�8e�\5�X�`�mI,h��a�^-҂�����UD�O'���UDɗ�ľwMV>�)�y�qH��~[KZ��O��)	���Ӊ&+����\K
L��o��TTW�~d �O���Dҥ�({��`��!�igڞ�p�I,��,�R��1��P�XkV�5+�l"�~ ����8��[�TV��p(��~�!r�'
|�p@��BFs�7!87$2<2p�Zz�)�?�G�tU/�Js� ���ZY(4&d>�$�����:�*�LK�*�T�5�.��tn�x���n��uxl�gXF�m���R�u�[R�E�0�)�)O)N)�QJE0�2�T�ԥR�yה��:�:��8�)ǝq�4�uO(�T�uN��y�)�QJuJu���S�y�T���aL�S%)�)ǜ����<���S�:㍩M"�R�R�ڔ��R�Sh��S
)M)�:�T�[y�yה�μ��S�qN)��m:Ҟq�KR�h��kS/:��aE)����n-o-JS��}�6�
(��(���ס��#��5S��J��ׯ;˛���{9�z4>�sS�~mf�'�Z�ݗ�z�׫�QG�T3�R�{��4W���:_�^ǟ5/3ً.9���]3�#G�ƫl|q���L�+O������7b�\cyg��y&�(!&7o�؅��ϻ">�-�nnwuf	��D�jس0�5e�L�y(�)+�����`(A���b��,Q�����V�"�����k.L-�3^9P>�mnO�b�H
rn4T�#�
��Sv�:�El�ܘ�P�g�n�'ɏ�7T�����MY{�OWV���(�ao85+�N�e�]�X�5º�I܁,7�o�jMXל�wۗ(q��ya6�Hаhl0��C{�{<Y�tk �ޭ_^�#�~�s[�l�)�f7l���,���s�vyXL%צc7f؟^���& ���i��&�^U�8*Eo�;̸ߪ����Z&��쌹"�o���~{wP��g>o-��m��ʼ�$����{�gu�>@�Kۖ�2�ȯ��:����*��K�m��M7 �nXYT��WZ-�QGmAd�h��jQ@emR����Pj�g*�DW�.;A'�-����	VK.�Z���1nݛw%�m$�4�"�X-��I���M+��l �������D8�	䓀��i� 5R���B0(�\E�V�̹V5b�	LEh#���:��19�V+��\�����ZU��F+6�m�4�[���mg��O0ӳǤ ,�$��W�����}�  ����������z  �$ ���y�wwwo�  ` UUU�q�y�u�^eY��l-�~Qb&�<�0cX��X�W	@v�(�5%����U�� 쮕;e��j]k�j��M��E	*�kf����tK��u�b��U�n9EC��w���rc6�[� �cf�iB;mv5T�%jR�Ү�2�ySr�2۫�e���**+��s��wiQP�I,ptPi�ښ�H��Z�)R�� 8��]^Z~�m�HHx4`;�p�i%�$�����N���2�5�y���@��~����F���֗��g���|E!���|�S�4l��ӢGé���L�|�r`��aG{"a��j�#332V�Q�n�ip��Oa��S��yD��SE,��cM�J���,�ÕR�;!)0��d�u�dɌ�
޽D���Ze�q<CǏ4\���8C������l����y��1#﵄�� �p��$痈����ha��;77�X6�7����ƀi6�sЖz�����J����s�D��I,�'�Ev}���pˆY�r�j(޷�I�M�� ��e�I��:;.�;N�&���B�m���6-�,��UT�A�"~���g��0���~7۫n�	���%�OD�	��Mx$��Z$�s:Rp2]-$.�ї-��⪮��:㭴�H���e��ֶV���F	��=��mx�a�������**+�C��i����3��`�\�cG���a,��؜(���Ǝ�6m�J2�<�{N'�&j��uVX�"�)�[HV�DY�B).t�ٕ����˓�vd���Tn&�-��a𲞆���jmE3�s�&æ��q�Y��"�;5>��$g!g��<�\�FW>�|�ϴ�l��)N�Ŷ�����Ɣ��_u&�I���'��QQQ\̽~��0�<: S��zi��ĨV�Ȟ�4�]��Z��/���4�����B�ZŋI']�x�(o
�h��Ӆ��s�?�x0������d�L�8,4�<�_�2L�I�I���j˻M�di��'a3ޒ�h�\��)'�$:l���t��m˙�f����6{� ���T��K�+�}��6ӭ��m#�y��ikel�m2�����jMggN�nn�H������o��N�M��� ����m�����-�)#�K�D�1��*�R&)�,���6�a֦Y����`�\�� P{`�5d����:I��ԙ$��L���jp��Z�5F����B���u#��U��"���'/RE�D�S���V���B�!
DCn�0��8�e��~	�"�C2J0���2a���=UUQ�y�Y�Lܡ��nC����2�0k�=E�M���a$�Kt�`�tӲ�\�q�HE�s��QP���n��#���s>/��Y�$����qDc�-�n͛.R;fŋ��&e�+�ٺjD��4zu�Xڿn0�F&�~㬲묢�S�-k[kem-���2�m�8�>�ؓ$�d1;눨����\����ny�y��p鐼G�+GgD��'Nux4OI�S&�M�U"� =*$��I��\.X!̒X�rJGP�g�tok�'n�z7r���=p���r3���*k6l��R�֔�wF�&6USq�D��,QHԢY�mˠ��,uN9l�~�`�o`�m-�J,hxC����.�f��g\��λ$'eUQ6��iSi�v9�uź�̣έ��Q����V��O�B�ý���VZl�g3o֢����x}G���l�
 �D��i�]9i�N�{`�0գE��%_�e����3��?g�<�Ԛn|C�/uj�~m������x �b�
�euGF�nR��C�}��?���8'�}��'�fW2"4ɳ��.��NL�=���I���4n�=`��(��a�
-��o\kMI���\vFō�L�!��O&ໆ�L:�h��0�孵����Q��pX��Җ"0�u�H�m-��F@a��'�4|^C���Jְ��0���ٳ�MΆ���Ҷ��v���p��d��%vK�rGU��X�"��K����!!�㗷��GL>��HK&�l3!F�bS�6<��hK�ĖO0^n��ż&��`}�������,��13N/Jnna��7�>M��p̓z0Y<YȆ�&
<`��(����?�[K[+en4����,_��)���]mN���7?#`�NE&.�ə�\xBC�af��TN�����'2rq���5�fI�E7�m�k	�̬��G:�*m��(D	Q8P��CT$�,�����"��;`��II(�l�Xs]Bć�e+�!���u&ڬ��QQQ\M�e
I#�(9�H��7o�&�M-&n��SD�+�,�����{)��C���j�p%�*�S�Ã/z$��������a��i[j4�/�!8y��qD�'���zq�10�x���|;<�0���dΉ&��K&��i4vZJ��lӰ0zD���� q<�P������oP���В�Q��� �n2 -C�7�K]��J.Y:�6;2;a��w.h���?#��Z��+iki�q���n\0�'U$3m�ǒ��v����JvrjjC�+�D6	��U�Ƞ��l��}��C��~!���K�M��Ab�%8ɧ!6e�����Z����HBu����m��4��j�K��{���l��*�"�eA&�챛kTw[���C�3����7zpv;: x�'Sxރ=�⪊�z�ߍM�K,�L�B<jL���i���g�i��6�<�k~yJyH�)L)JR��R�E�)L)����:�i�^SN��Ω�[q���:�q�qN��R�uO)�:ڛiL��R���yH�<�R�)JeJeJR�R�mN)Ji��uL��:�R��)�)N�N)��Q�)JS,��S�y�<�S�yO)ǜm��m�4�
R�R���y�y�V���
)H�)�)N)O-kZ�qm��х�Q					Pj�u8c��h��Q��Xb��Ͼ('����`����ǌo��/�]N|U�)�㷢��;s����ٳ�qW1.�+.p�7��V���v҅�[VG-4ͽ؃qeU�F�*ƶu���0�>�=Z�le(�;�L_Fc΢#�˓;��M�*-ANX)�c�zaQ���(Ɏx������]%\�0'��+�}iˊ�t�P�T+���td�M�n��4׺�{���ے �/�mE��yj�ͪ������9�e����  ����滻����` ` UUW�������`  UUW�������`  UUQ�Mr�ʔ-\���G��ֶ�[Kmm����2�!$�j**+��EzɆ烅;:����_uu�E���>OD�p�H6��5*�\B�۰�NG	��3��~�K�صa�w[�U�۩,4�cV��вL�K�������E�	�$��v\�2�'��(6�\�4�l��9	(4��SI�@���;>�tq[��-��"��&1�U�8�n�����ֳ��>>:)��p�}����W _��1,Tb����篈���.��La�0�̆�D�/�K��/�R��=�Qr��縱iZ9��5�1���e�Ƀ�U����m��4�]�S�60�E<l�+�@�)�d6����2�%�v��tS���9#TJ.���7;&��E>��v��|�R�J9l0�ܚ06L^���2e�tܑ2��2h<��[�ٔ���s�yƘ~u��<�ֵ���U�b��T(�:�Im����r��c�+D�d@��	�m���I�˶�u�ؕ-�VJԱ�0��%V�)Y0��dN,QZX�`䕺"��(��%E�PQ�-��.>=�n�ٕ�v����jl^VK� �ja G@�h�ƥdi��E��)eA�ϻ�����Ӧ؂6vr;u�/��ә�*y�'��\�r]6,y�u���Ov�4{��'zͻxC	T��xч�r�}%�a��)��?V0��,r&��$�O��'�g$?0(n����
�*� �N�r(BXD�K���,�M�FS�M'	�)ϙ����e�[u���y��ֶ[K|l�8]���)�)�L�`5�u�j**+��dΌ)�:��?a�5�NI�ꊿ�����o�^�0��ۍ90ll�):���T�T�Yѷ�H�% T!��u备�"]�8<�z�Z���ڤ� $G�F�SY+�e��wI6��i��`�̎C�F (/�X�$���l.�II�Y�i��IY���,y�l�_7�t��O�{g�0\�g�x�y��Z���[Kq�e���>�X��K1�M��u����8h����<�����0��������*�c�v�4[�������	T�6l�0�;��C,y񾞢��㕪��BS�%��w]���2��T�Z��ѐ�wKm��<ì9��sӁNg�e��/hᖯ!���Ӿ�N�ɭCpEQ�6؅�lMzFC]h�6�8�a&c��k�2�L�xǉs}K�6p��uH�?����Z�ecry���2C�����QQ\'���{�JW�N���&<�;Q�39�_2~�wuɻ�������V��4��i�M6�n�B�KM��,a��6i��]�ic'�9USL����v�`�X��c$���T
q�e�M&ؐܐ��A�;�k*����v�4%��0���\�G!�f80�y�xp:v|#0�����c-�������G�m����B��~�ϊ�2ń�4�i���"ؐW�=h���N���7z�X�Q0B(�c@F͊EX�T���b�ٵ������L� TZ;6ͨ�,���h��j�^V��[Zj@�������u�ұ;k ��ʚ�8��vċ%�DQo��Ô�NR��X���[]�r�.U�Ij�B҈\��n�bu�8�:�qc�T(��B-sA쐀���鼶,bLp�m%��]be�6D�G�vz�P�xs���S�S�<.�aVa��լ�BE�!�m��Ĺ��KZ����{�N���b�Y�˃�qټFX�3�y�4�4H����3y�փ1e��a�d���`�~@��χ�wP�ibвl�l8t�L<��E)��������8���$ �#dI3�QQQ\-=�P?6M2m3̭����۩?}��=��?Oa�1]��a[KPk�s�`vh�τ�CA��}5�Fϴ�2�n�2e-�%�o�D~<)�P�����̰��-�߸V�����uTWc�
�(G��u%���_m=��B���`.�]�R}�1��K�:�i��??0�)��������(�����#�F!&�?yI&7[p�C�|EEEp��ς�a0wW(�T��Bͺ���6�p76��B�'��7�x�f\8��,��U�]Q�6��D��.C��?N��+��g���g���h�O���Xz	���6ᠦ�C=T%�f�!�	�Y��*pٰ�	s�{�x���N|�����ʝ~~S�����M>>6`�.���b�-����QQQ\.����t(9�s��)��O���@���~Ӥ��KJX��h�V��i"We�r0Vl�Q%mj�&��Ҝ�+d:�7���M�]���b���U�ԵQ&ͧN; j_��m�+�nj'�O���ٶw�Ĩ�����,��dT�8ᷞ&<�!�锲`�9m$�T�ɤ���K/�(`���.h�F�)�y�]u�ה�5'ԤR��)M�JyO8��E)�Tʔڔ�S.�מuה��yO:�n6�SO)O<��6�yJyN��T�yO<�jm�*O�H�)JiJj%<���S
S*eNa)�)���S�R��S�<ڞi�eE�0�)�)O)N)�yDR��TқR�uM���R�y�<�μۊS�qN6�6�je�m�<�)�6��jq疷��
)H�)�)JuO)JS�qn-�XE�Ye�QG���O`�c��n��m���p6`���f�3r;9tm��O]5�o�FBO^9�s��Wh+$z����v�{rt<������<rO��w=��.�����i�ů�h��~O�]�n]gvw�ա$�ˏ�����>��cNLrז�]���l��|[�{r>�s<d��;����RvŸ(��x���x����\�.K+FZ�LQ̙rǖB	�����z�ј��'o�2`��� R�,��F��n\�QD>?=�k��Y����Yy�&<}vl�ݭ/��q�;iy	,���ڶ���E��ǿ�.�������Z�4,��}�zb�dvd�s��40n�F�G�Ŗ�2fC�fȣX�O�*_���{�;��r�}UFz�����z�"�R:8��5�a&v:a=����z��w����,���R��W$�w<�����E�r����Ìs��r?Ee���n�'*�v��O�b�M�UJ�I����p��ڙl)�x[S1���)�mb�y)nX��ʂ?I]�;j��u�>�^E��m��S��F��P�f�_�:�z����j+ƥ�*6B�6�p��ؑ;J�b� �d�(�$9�kl�
�mAL�N�V�f��I�|�#B����*�RA��*�|cB�8�Ӕ�9h����mM��F��+�V����K������J'b��#V��Aq��1�\u���<�̄�멵��ɚ2	RZf�m�n��6����$f	5��B�Gp�}���s2�ND�1�"��SR}w5���J�RԻ[[.���6�wsU�T��8������K������W���~~ B 
��=�wwww�   *��������� � UU������ � *�����-\�B�^y�YKZ�����qm����}=��GT��mk3d�鲔��n_�6\a�Nl6ݒ�]�Q�y������$��+
Q��,���X�j�ju7�,�� DXT�b�����d��h�tSMȝ���	҂QUED6�F�ZY`��%����ꊊ��w��:�v�-�k��l�m�m���l�b�0Xz��n�v#��{4�4UT�hl��&��H�3�ތ�6C��K��f�4��RbFOqٞǁCZi4a��ád��6�h�c��Oq�ֳ�(�*��ۆ�{�ĕ�ד˹^ۇ��ݻv6kv�K�9�7J�la�-P��B��=r���w���lq�����2�aoΰ��O�[�O�|i�Ѥ)�:ڧ$���~��S�*q�'"��Q�q	5��$����{�GJ����F��#�'�x����)jHV!��>��I|���M=N�w;P�����xMxL.�4?^����5�6j�ݛ��lHv�ww�Ԑ�c�	H�����k���xB�0��a��4X�e;� i�䢮�v�2�<����&]�
8���<�����N|Ӯ4�Ke�����ֶ[Kmn4��˯O�����b��(�a���,~֦eKn9�W��1I��),cI�Ǥ���G	�����e��>�/��>�4��=>=�����~�kDo��t�S�B�v�쑌�~?}��0��ag�tԚI����r�M�5�/�U>6�j:(�p�]:щ$MAxy���rَb��s��z���'����<�M4�*a��G�k[>4���Htp�yie�H�Hl�qQa�nXs�����ϼ�o-��a�K(��O�ɹ��j�2R�;��2gA_�wf��鼧�
��])0�6m��FY���Q%XL�"Q�t��u�D��ǩ�� �\g�����ǒ'BŒ��:C�w!�ݒ=��;n�׵��N��D�y��Cp���_�m�)�/���>y�˩$�����4��q�Ӭ�ì#��kZ���im�Ƒ�{����E�Z��*#�Y$~x�*�W%��:�i����`�;#ɛ�iƍM��1��s��a�� ��J���O,r˘���c@��Ք�S��`:[6�d$�ii��p�,��SN7�*Q�&
[1��@��3��n�t�Еj�M��L�L�	۲��{k�ZT�J6d飁�y�\�]0x̓N��L�/$,B�; �OD�T�l.��r�UW@�Nw�cIĖM��=M���2g�p�=��ә��}�\�-l$�76��3d�ْ�n�ݕ�˦��,Qb�R��8Ĥ��\�8r��M��u�URI�p���ᧅ:�#���kam4���8�,_�E�V�G]/z�(���RL����ܕSI��a0� q�e�y�a�Ó~z����G�˗/j�#��I����M�D�h&�z*�R��C�~�k�ʢ���{�鿼?(q���D���F�LB���EAa$�*�ljp���w��Q66R���d&K�5V���M+ �塌���S{�A��NțM�,h4繚�z�^�r�Rx��os�������a�^i�Vì"�?-����[kq�e�_zz�~����r���E�a�ti��f�$��I�On�9����!GBe8�`�z��krG�v���vf@2V�+��HQ�r��-lDQڨ�
��9*�q������<(t�p�?~jdD��j�Ϻ+���p�(x`��DI��8#n�m�z;!�_:���=��O��C?�mK_T���Y�a����e��u�x��kam4��f	Æm��DUDuLqI�_:�(��s��a\|aMO�a��jx��Q�y�~=������ {֬
���&EB��( �0�4]�����!��m*-:�~��d8o��.��!�?
o��bn{<!��N��t�f�g*Z�a����ig	�.��H�J�Y2��)�8�1X�H����M��_�;�33�:������Y~aL#���Z�[m-���2�*rj�SY���d^k�Ǖ눗69�3TL�Y��A�����낶6�|�*�((_z���8m��:9!;s�@ܬ��Tj����NZ�J4(��EQjn
��,�Bja�j��l�#�A��W5�1=l�Ue�В�j�E\\��Q�+U�Jh�Y�D���w��{$6�*�$���v��4�.�g�!�4�_UϛoN�b2�6!�abd�9-h�Xzw��CN�adَI#2v����{O�,�ժ%�~��P���)	gV�hEф�seҚRmsTW�OI��	�<���M1�B��(���u�S򖵭l-����Gz��PJߋ��2r8y7�����tI�������Jy��ʚmi�W��L��t�R]{͛<�Ҩ�U4FQt�a�`���F1z��n`����WY��l۴�1m`E=ˇ�~̹�~��d��9�c�!�nk����j�m!�1�jd��M��fB�`��R}L��=mţ�8���)Jy��R��)JR�R���E�R�Ҕ�Ï8�yJ<���6�n)Ji�R�Ӯ:�R�So:��󎶦�aE)JR��ԤS�mJh�<�)JiJmE)��ҞR:�0�}IJf���%)�O6����$R�R�SjmJuO6�y��y�)�<�]qN6�o6�i�T�SjS
y����8��Z��
)JaJSjS�S�S�u�6���+0��,��u�z{��c{�}��[��9�T�9�2�U���d^<��;��RVg_r�iֱE��ǝ+�S,Cuu
���>ggk=&j�?�)���bӫ�]s�k~�J�2Ґ����~�_�\�^*���.��z.� �_��h׷��w�'i��n21��l.���Y��_�{���:yueҼY�Mz��cໜ�In7��b�A�f�w�<��wk�=��c���ȟ�߷Ћo%�k����g�x@  ����wwww{�  8`UU]������ UUG��www��   *���ؚ嫕.R�B�	�^K�-kem4���Hˌ���"O�5��F��5D�aÁ����={E*X��}?OO��1��fP��<��[M'K'��"Y9�ѻ1��x�� ���,����
%�$��<܇CI� N0�Y����D�L8����I4��&���\��d�$dvPX/�)Y
n�k	�(�r�K(�D6<qk[+i���Q�j�sz�Y�>MLkX{⪡��é�U�Gޞ�d==n�Hi�*�L��İu�
%jZд��ڕ��%d�k7#ZI���<�.l.��I~�&���w�e3IQ�N�Hi�m˦���8$�3��nz�]C��׃N�٥b*�ЮGp�牔��������QF��c��ٹ�����i�O��H~??������[��.2��Y�0P�v򊌧�H7�S�y�9�)�����Y9q�9�tWi��a�f,��Qܡ��fn�{�#C���0� �:'�,��$r���U�� 㣰��3*u�	�ӭ
J�RTqX):,����9%�  �C"��X�{�{^r<q�`-p�M��*��S7h�X�%ݗM�^�Jԓ%6x�,��I$���W���y��S3�|�z����ǡ�.U���h-#�oM���.�qr��	d�N��hd$8a�\�I�e-�)���UkQ{�a��")�疥�M�DLGqj�K��R�k*����򴜸��p��%�ҡL�YX`�]��Z���k���`�V쟾?*�)Y��x���Z�m��y�0�)�KZ�[--m��8˾��}�&`%��r����q�;d��UQ���r�a��TP�ֽek
�y�C��O'�'Z�F,a���5a�Of��mmnC���	O���$&��:��!#r��d�֍p�{��y0��d5�M�֙�����m����n�������<lv��2p:fHZ�p��Ò��V������!��q�:���Ts��=	)#���M�!��6��<�<��R���[m���>�Q�6���f1�djI$�{0�x3��jֶ̜�.���Sfjo��s0Ǉ��L�g���G�γ� ��`��#3�t��T�qݯ7Y/�G��Zo�f���O����%��;'�w>��[�[R���K��b!ћ6��h��ًH������0�/]���~��[h�ߦ��;3��鲞�t��a[�JZ�[Km�Q��g?rg
CHdyUU=(�稧�L�K��5�!�Ṅ��;�v̧�X�l�f��ؓ�T!(����
��-s侯�O_IC�=g'�(�y��B8�Rd2�tH~�G�L4�h*6䭷S^��@��Cy�fܹ>�Κ	�bd���y��\ޞ��q�FB=�\�����tnLK�K��vi�N��Hx��R��V��m����y�;�ɊIx�.f+	�����^Q���E��
�+����ZVF�'��#�V܋b��W3O����]|�vEV=�Ŵi��M�� Z(�u	���+�<*�Ö�4�D�!��v��/!#���� 	l(�e���m�"�U���K9�݊�\�D��%e���|�BB�XӲ���|& �n�BI�^�&'�wi���;�I�ρv}}˗..rL���<��b�^�Ч�-�ODˇ%�:�ꪕ����F# e�l{F�	˯����cY$Ȍ�c`�]�j��k���eQ�yP:"&D�����ӽ�>L���)���]b勚.�2��"���R����-�m��ч
�6���cB� E�.���ge���)�}��ag��7�mj��X����i�	�SM���At�C�UJ!��r쫥6/8\�s7���>V��?XK,���Pm�ӢVKBA^UXuN-Q!sp��2�����ּ*�����,���rlJM|�/|7:����g���W��[*SKe��G��)Jakil��H�l�>���>�}���d�9j�x��r8z{�j��{?&�_��x~�;�y�����*5]0��bƇ%�p�����O�2��eɘT�8�r��
nHw�<L�B{z��<M��B?��J{����:w��TWp����N�8i�f��_-�b�hF6��6C&S�Y�Ju2�K&L=�FNi�TE(�)L-m-��F͘;�p�)C�oj��F_[��Sv�\�=s�}]������έݥ�]�Թ�-)V�HN�.�-O�Ӷ.�������)�>C�F�eI�o���;�ɖѢ��j:SNĨN�w�|�];ԗ󴉅�������CZ3�,X˶�/�����A��I>�$�I$��TP�?����~���e���Z	?i�ر!T@�WC&'�����,�聒
�"�B"���'�(C"I ("0I�( �1@A�F$��B1 1 b��#�A�� 1#DA�H1 $@bH1 Db�B0H).RI� ČA��A1#Ab����$@bH1�#�E�#!����D$�B1����# ��@��'�D'Ј�� �'�D0F Ĉ�`��("�$ �b��DA�1�� � "A`��D�����A`��1$D �1�"	�>�O��!O�D �1 "A	bHdH)�� � O���O���!O�D$�#�"%��DA�` ��2" �H��H��0DA�"2""$��1D �0I ��2" �A��"A�DAF$���D"D��01X" ��FDDD��0A�� Ȃ#A 2 �0D� �A	""#DdDF���Ȉ���Ȉ����B0DFDA""#""0B"2"���D����"!�� ��#A""#""2"e&!� ���������DF"#����"##A"#�0H�$bF �1$b"1F�1�A`� ȃ��DA���DbH��D���F	"��RB�� �D#`����D��DA�� �#��b
"H�Db"DF"���"�A� �0D`��(�H��E�1"H���	"@,EhH�!�A"�"�H��lA
�A$�A$�E$T�D`�	�0$	���	 �H$D�A$ �AH$Be��0�Db1�a"$(A"0H�H|����G�|��H!�H	�H	�0H���"A � � $ A"$A"�A ,�A � H�H�� � �!�0H�A" � $ � �� @�A �$ �H�A",�"��H b��0H#�0H��A $ � �(@���H	��H��H��H��� ł0b��(���`����H�A��b�*A�0b(��A�^L!�F0��	1�H1P�1@�	 �T�DH�D$@"D B	 A 0�"I ��*����� �b!���(A�0 ���"�! B$A�"D �! � $d�$�D�� ����"�"@�A� �!#(A�@��D �� �$adRT���@� �`�1FD� �`$� �H1X��,���%HT �#�Q	@dH�@bDH�0H� �"!"F ��"D��$D"F �""��A#" Ĉ$ �A0H�D��$dH� �A0H�2$A#�$D �0A2$D���DA�2$`��"DA�DH�A�D0H�F	H�"$dH�3(I�$D��"$`�BX1`$ Ń�(bA�	$A#"DB"DA�D'Ȅ'�B�B|D`��A� � �"�"�0A�A� "�"�"�"D� �1A� �D�"0DF"�F�����@D��1@c&%HD`� � �A	��"#� �1@`� 1 "F�AA��!��G��B|��@b#Db ���0F"##��"� 1A�"H1@`�D �(�1@b �`��� �"�`��"D��D�H�H�1"$bD�$`��D"@DbD"$`�! �Ĉ�1 "1" �`��"H1B0B1!��TD�b@�1��!!!$"##�`��0B0B0I"�	������CI`��`���A꒖�X!! 0IF! ���!$b@bA�"$$��1 1$b�A� ��1�@H� �1#>�� P���n>�|�xҔ&Jq������T��ET�1>�|R}_�_���z�w����O��.��Y����ϟY����o���~q�>�������9^(_����l�����|�|E�ھ�s�.o�O����S��)�������> ������o߰��A�j�C� ������آ� �4!(���'�\��?O���H`�X�)K����6����)��|O��C��QE 7�П���ℐ0��4����"}���v7 ]$�1>������RRbk���@�ݜ�nM}��g�$���_��/K1��������l���T ��@��" �, P �@� �(�ဪEdF1H�-���P�����r	V�ߛ���U��O��'�n>?@	*DI $R"
D@ H��4��2 �(H0���K}f �����L|�̏�}���������?�����a�Ї����~Ϣ@���'���e��Կ�?�p��������#_�C�+B?�?�� ~ �7������G�!���_󟫿�~�G�>c�@�~�@g�}�!�<~[~���gzl��!�����"�r}��QE ?����X��Nk��V�}�t�e|�飍�
|K����H(����HC�f~��x%�@EP� 0,�'�l��prwIID?�)�2��6�u�?F�.Y��\Z	��O�� ����(ϧ�~�b�(��?7�2'���	�~�>�����|�l�'���H��_��ڧ�?�>���?g��:3���
IG�#��������qTP�S�T�K+��"�(�~߸�r������'�<X|������K��:IT�͏�ܸ,P\[��������$���o��VC�	c��3�[���\��QE 2�AC�����~.S!
����� ?!��C`�*������;O)����d�aR������4)��'�D݊E�P>k�
~����>æ�@Q��.�˿��R��򠡙����]rO���}�?JUY 0S���7��ܑN$�J�