BZh91AY&SY�|c I߀py����������`�^����            ��($�*�PU 
�T�@) ��m)�    �   �� ��ou��v���Z9oZ��zf�^�>#x�{��>���w�+�������f������v��mV�����}� �@#�yI�Q^�ԃ����u���}u��t}����z^�=��k�w*�w<T�B�w_Gpw`]aZ��Wm�� �N��f��Ҥ@v��{��y���0a�W}���<{�Y�n�۷}k�O�v;�8�muV�7����>�  >+��m�s������-�羪�{���s뮫�>˭>=ޛ1�1�O[ڈ}���{y����8  �`��g]g�[��}�ͫ^����p���n�������{l�;5}��F�<� �D��  "���i֒���T�:��  @    �:CS�*R��b4��4 0   ��BIRTz�h`�	�M4`�$$��HSɪ~B4�S���F� ɡ�&jR jUP�И���0` $@%HSO)���z
z��'�F�F�Q$�U2�&   h� ��a!� ���~�o�> <I�&����H�H�?�@S��r�Ԫ�� ���?���ۇ���i��R��rP����؊�$������3ʿ��Q S�����4UUUNJ���r�I 1k���O���+w �7�Ց�%�s$n�,nS�0ɶX'}�M�����A��A��:�s�d��0)�6�;'Xk	ڜ&L�n�d��I�k%�y�tLT��Q&��!
��2r�&�~��d<�3PgQ�35EM9)��ﵐ_�I8��Q{�AƔ�Ζ�fö��:�����ICd�6f���,�.䬑��Ҙ˛eU�U0���%�j�L�2�ю
�E�����²�˳�e2u0R$�t�51%�*��eh2)�}L��Pj�tS�.�l�e-�VR�lŖ0��-�V�-I�T���e����x�ZI�&�Jh��*,���(���,�a2��ZU�*�+I�I�Al�%4t�&�	`��-��Q��ٻ/l�g^D�J�S ���ZR���d���N�Q�f�@�	zSf)�lɂj�U��n̻)ٷ�6N��L��vn�'0K%�ZS�)Ɣ��Z^2���U2���	�FM�}D�Ixa�M��M�*$�2���­�X��l���h�El"�NJʲ�ƐfIa�����$Y&�8�x^����ݛtV�+\Ѧ��m���/͕M$��[E77j-����pS��Jm�d�$��h��RU��x|��e9�Q�F��&��H��LT
�`�}��K��	f��%��L�(B	
D��i9����5�C�gL�p��3T��p]Df�|���'x�/|q���������:����E�Bh�6f����v]�T��N)��WPUL%D��W欥��l�Z�m��Y:AҖ
Te�N�9)��!�����EDJ9E�*��e4ϩ��Tj�tT�e�M�L�������1e�!�I�E��:��b�V��V�x]��&��e)���QeŔ(�D6K2�fS)i�e\"���8�-��M'	�n�@�	Nil�2���Ku�L�e;:�$�Y�eXR��8�-��M�V��͢�,/zSf)�lղ�"s
�2��
l�&	d�8b該��2N��6K4��S�*\�KK�V��tS;�N�0�l�$���Y%ч�6j�X��+0ݝ�*-�Xl���jJ�Ed"�"��e�"�cHbbȰH�H�E�i�O���:�e�+\�
h�Ej6�N���2g�2[E77j-���F�4S�NJm�d�$�i+��*�D�!�ZنMc(�ӋJʜ(dx�]�e����0���*�*ޔ��*�
��Rb���.�(
���g�$�'d��,i���W�)�lg�ƒ��c]��JL�AQj�A׋�ҙezC"C"<�B�Q2R�zS�U�����UI8�,6Il���%�&��)���Ҵ�dhdo�J5%PN��E1Nʼ8���P�<X�E[���ԃҬ�$к$�$�d)ED�TJLUi&��$��$�MD,CeL2���oŌh�'\��)�*��)���>.p�N�W�2$2#�J)��vT<)�l�Z�є��eP�$�$��%�N�S�LY&��)��)�W�d0��d�H�T�)�T�1�QS`�?$Z9��5�R����.�6�N��iL���dG��l�jJ��E1NҠ챎
6�/,�xS��l�/QV����TR�!͔���H�N)�b��Y�*�m����Ɗcz�A��a����y��#K����!LS)FC�A��
Όp�ed�#$�v���0_�$�0B�
�0�(c�u�h;�Y�>t�*@�D`������Y`��ؑ`�`�^b�L�`�@�`�����Z��`���zA�'(�	�0�>�@����fD�a�1�č�䂃�H,F�D�4'��.�v�:I�)ޕ��+�2dh$T�lXO��9iHxXDc���L^aV�-�V�LA�N�����TTW���`2`�'��,CªHS���4V8)��I�f�g���>(5�2����,�y2�e ��
b�*���3s��2�9$�f���0HaH��A�AC������xH T�Ŝ��A"E�^a���`�_���b-�����1��hV�W��.A���`k�̐_��S���tXo��t@�`���c����؁PI��C�CX(8 �0��&��c��`�R E�Ė�2�,S+p1�6��Ċ�XR���@v$8?1l1���??1lc6�!��z��R*��� h#>�|Űpb -��"��A�A��j�1�p�,6tn�V�O�tV�TjMAb��A.K��8[5m+f�~�dߠD���$�ҵ�*���6�d�NP�e� f<i�4���8��;#r(��T��b��7�^Ѵ/F�ć����B�B�4��4�'o�?_y�|�i�Ɯ&�G���ۤ�1�'0�$���X�I�E�b�y^��p��ʸ5͔���Qj��}x���uN$�r�mc)�;3�y5-�3Y�g9y$J�T��٭r�Y�q�r�]c�m Q�I7����l�9����>Bu�Έ��jSU������o3�n�7����'1����V_\�\`PH�B�����x�wAU���	ڠ�,U`��V�|)�d[�q>dd �	P:hVWb��٪&�l�C�����98/���zJ�i�1^(��/�~��dGb���}�p}��~�R9��s=G4o�ۓrS��z��3���:��จ7�;����s��Dh���[8���}ӗK�*kȍ�^�7.b6�!i�X��w���x�6S�Rw���f��2���t�1p���P��\���N�˧?s;�!q��:"DO�Z�O����"�������#����Y�nTs�����,B�5ҹ�L�.s�zł*.�ʌ�R#�]`��R��N�c�$^�U^��+q$v�p�-l�'�A�v���Q����V�����f����'�s��G�q�M)���_���:Ϻ����`��b���#��gą:>s���u�����w��6��\��1ꃑXE2$���TC1�F�lUώ�B>��.���'�]D)�sMk������X�w�}9�k�>!z��=Y{���xG���"��Q'P��VP1��U�OH���PU)�6(p�]�ū$4A�I���\��n�Ċ���M b���b�R.5?9�Sއ��[d�Z�_)�"�4�t&:R
[G�j_s|1uz��r'=�4��&�}Ǯ��!�9ءOo�'��6oQ쏰f��t�� �*�8Ƚ$���K���m�#_��+�K�~}G�!�`��r��<(�7p��Q�ǔE��H*���Z莾J3��1w��.k��1	�D!��"^�;!1A|�og(�qo)sw�9��p�k���7��i,���tD���;K�y�:!o����a�!�R�t��M�О�%{�7�Q��b��!ǣ�J�1���%Ð.�~)�P�;���е&#~�A��M�b|�Q�'.=�9�ES�o��;.�8q�/��9��>棥}\</�s�;#s���J{�p�#��_�C/�Ӈ�yR=;��%N�\�8�e�ԙJ��|Nup5�CI�}H.t��6��4ἄ9ɺr�,������@�7 ���FH�.S��/t�:8�γ~�8ŵ|L��ZBE�����M�����g{����>3��'!�Orqgs�P%�	���5Zi����I�`9�C��M7˝4��&�*�,~��������"A�Ȇ�'�x$�N�M7���b�)"�|�8��A�^�*���qt���{�%��m��4ZJ2u�pD
�6(E�CEdr~��ap����HB�Q�X�ʠ��Z."(H8vg��K������>��-�SL��F�s��I����}p�������r�����]���{`��A�]*'�oP�J��
&�S|��-��˓�r:6'
L�y��8�s�Eڗ�u.oU���L�_PTYɘ6���!D]]E����9���v'����{��GO�8z'�b���S�g��&��<��*��LL�W��;��Ege��&���#H����1�|<l�'�e2`��,�th��k�"'9Bm�SXE&".���J�����%�x���]W,Ư�<����y��r͓0d��DŞ�H�5�B���R̒(�jͬ�����&~W�$XK�'�:��:���Y��ث��t�<o&��s5$\���ʘ��j�2��������c�Eȓ��$�u.+
E&��k㨬���1B�aD&ENLD�,����j�g7�������⫂p����^���=g��jꝓ��~݇N�4�!��{����=�[m��toՔQ��4Z@���M�&`���jcGVQC�ffMa�#tPS���P/���K2���qUu&��wP,e�R �y�mZ��%sa���`�ˍ�ns3 ���1)��@9;�.6#ml ��Ȍ�FddǠ�MI�U�g'nd]DmhͰn�mP�Y�6���D���	�aeBܝ����,�[0/7�E
���' ��a0���7����(>M���͊����Ey�c�f\���e��$�t2�!QD�"��YDmw+"�NЦŋ91�՝�9/׷z�*Y�ԧ�T>Rz�Rsp�sI׽}ݩ�t�UY���<m"�2���vqbۛ;�9��9F��S��A�E�T��D�k7�,�����."u1k[8�ߊ�[�q�7��y����O�Jﲊ��k��ϼY�D���+�I�[�Ĭ���.Sme���K��#W�z>�c8fe�r�i.:/��&>"�_C`T?�!�:��m�D�+��Y�^���(�������~�>{��64���/̽;���e���pߠ�|g�����k'ӫ���L$3��;"»��ݾ���ᏺ��?�g���4�5L�Cq#n�y�#�VV$	����a�6O����>��h�%���5-E�<���z��{�5�1/W��#�EW�����I�q��r�h�UY�-�JI��UX"s�N��m��m�Ȃ���yX��|�MQ.�j"�\]ߣ^�RE��J�k_籮o��g��fGĤPG8�gY�Y�@�2fG�CF�m�%���{��*�ؓ>IM�@i�>ŏ&Ǝ+�ߵ��
����n�������/iV���4(d>ͰlN���b�4)D/�3�>S7:V�h�{{;�!$�R5�|~��y�dS�U{j�R��V>b�P�ȬD�
�Dk�4+�����b������X�B�nX"���s�Wx�1��`��·N�YM�/č�D��d�ww%�ȜV�Ɠ�WNn�ڥ����5
*�*e�+�۲1��wfq��b�T�G�)[�5���.�+F���:�BJ�Q�K��L�MBq,,�i	����eL��FF�lQ�N��g7����ĴM���ji�J�M겨��P[AZV�O��Ď������)$�F~���"UQH�kĹJ<��R�3W6=�Lh�Ć����U��Z��vc�%�n��׺MI!�M�.��F�Ij�"bI���:m�'t��}�)���Dʅ!&�V�D���<\�Lr3eVNooy7�p�P�"%��)S^R��嵱7c#���y����w��^�޶�M���7����!�I���� S��=�ݭ�d�֣�
���{j���B�b��%x�ej9�lբM�Wd�y�l�;~�9�.eQTՊZӕ+��	<q�϶[i��r�h��%�9����A��&6���h�v����A�Z��r)���n��UZL�K�e>�7MJ��Z�(�,�����庫�Gj��R4�a�p�ͽI3���iL�i�6�lJ�����b\M��3E�N��/
�)EiAB��A�,�Z����rb�sƲkx�*|���#���s���q
���KF�GS���j�4t�Y��!��I��I��fT�,�jGS�K]���9�U���X�l���T8ڵ��_*G�$'�A͉#b[ERfX�c|�iK5��%��Nn���Gi��,kvG��Ȓ��婅v������F��cԈ�۩XР6"��Q6G �bT���$N͘Ө~r5O�H�M1�C����I����j�j�ܑY~���+��R�eG)h�y�5��L�Z�S�,�k����@wy�]��6��/q  ��_Bb��*��/�N̒��?��ޏ��}ϳ���>����[��}S�}���f�i��x�m���m��a��m�-��m�m6�oi��x�M����m��0�m�m���m��۶�6�6�kt��ް���nfe�&�n�npx{�a�   <=�<P�6ܶۖ�t�p�m�m6�o-��z�m%-���۶�r�n�nm�m�m���m��a��ݰ�m����r��������m�m��3.�m�oX< ���7[oM��6ܶۖ�t�p�m�m6�o-�M�nm�m�m���ۦۖ�n�n[i��x�����m��m������ζ�6[m�����a��m�9� �=��� #�+�����m����m�m�m�M�-���6�M����m�m6�m�i��oM�۶�6�6�v��ݶ��۶m�{�wwv�n[i��oL�̶[m��������2᷍���oYm����m�L��ۦۖ�I��a��m�-��oYm��z�m��6�m�m�l��m�i�ܶ�p�m��t���m�m�m�n�����ۻ��<���[z��m��6�m�e��m�-��x�m�D6��m��a��m�m��a��m�m�m�l�m��m�M�-��ol����{���r�n�]UCm�m���j� HH����C��EU���O/7����%�� �APw�xw��?����?��tۦ�v�o[V�6�]6�lٳgm��OOOU^��V�m�m�m�z�o�z��n��gfͶ����m�m�m�zǭ���<vӦ�m�g����;m�o^6�mi�+f͛6��<t�^;m�M���f͛m[m��mѷ�ǧ�g�C�9�S�]�ǝ�ߣ��=$6h�1C��J�tEZR腅B#I���7�Bq��t�%���-F�!���!p�JJ�C�R�D":	{A���e��l��1�/�����݆��B�n�D��-�*�Ő�N"�ɸGH�DD����M�2��#�B!A�#/АEh�@�i��7X�C�@�NI"[��R�ͭX28��+"l���r�I�\�X�t��,��<�&.~���y�w��n]�m��J[�augW��Y���G�:(�ŭ6>��MqM�
����5<me�*2"=�Č�#s�Ķ��[u�
�P����j"���,R�2��)^G�F�bz%����Ӽ���W�����=��V��9��ك��=6�m(G�'K��QL�����DR�u���SRV%H�I�MD5�n�*l�HY��dDr<�̵>�ʚLڐꮧ�.y�޹�����%EU}�W����o�q�s��s���]q��.9$A�˻��g�>E���;�wuT����E"��3��]o{�Ϲ��e
�����⪸�../��s_N�Y�L�c���&l�M�I��F�q�ݖ�JVV�B�H�-I\�qG]n�ݏ).ɮ�Hǵ��V� c�iDƵ��m��Y�5UT�M<L���y��Dlp�����v0���g~5!N2<r8m���p�����)�O�pD-�u�d���+������m�|f���#1���dj��q���I�)Ѷc���Z%9�H���9�$y��u�������h��9���@]�q�AN�� �	$�w,�BH1n|("��o!��4`��!��cx��˙�ub�</5�]}�a�����g�LZ:��t�3���	�b�A�!�z8;<$���a"a����}�*��80������xoC:<a�6��4�1���(�f�*"����|�\s��=�ӂh�cjn̻�m��{�K���$"��7��5�Q�+����>X��w������2�'C�8w(������h���+цm`c�]�t�w�l��v�0�����#�1�f����S��dl�1��Қ�wE�y�3���{�"�e9����r���%͏b�1s��İ�Qn��㎤�r8����Tm�n�m�UH�h�HPD�E
���+�
`t(�$�"���̷Ǽ�w����1��������{���dj���:�te�bX����1�O��o�k�ΨB�lVZX�c�:������I7� ��>�t�1�G�J��ϰ31�#�c�c�ְ}{f���P:F��{w�[{��w>1g���f�9��b+���*)m�T�`���c�;��=z�zN�i�aO�a����c9wWt�t5w�x����j2p�8�5F�& �&P��~�1��$��,b&�$���#1��wd�69y�7�!I���B�rOK������}��=$_SOMo�x8��`���|B�-�<�!�1��w�c�s3h}���1�������Wc�D�!ZIG��BB?�cc��ٗ�t�5���݇s���c޸���8C��k�A�,�c��6���f͔9^;%h�
:d�!\G�0b��G`��H=�ȈBL�]yp��nm�M��E+�D����Ԫo-�G#�r��H0�st��L��\v2$�KU��n6�$Q���9
�+�MI��U
V���L�V�۝���g�1g��/����C�����[��
�%Qz	C|��mxp�ꨢQ��C#�<s��9����Ӫ�iRr(B�� ��-P8��a�a�ܫ����-�%h�
2x��,�Y��w/����9(�*[weU���ðӚVB:1��q���l���CQШ�m��~��m��Gԅx"��W�2��F��䴢E�!ѡ��g�Y�3�8ձĶ_!�$�yz1���A�&��|�!������j-��UzY��U�e_U_1W���˓����W���^/K�������X�Z�+�W��Ǭqt�ƭ�Y���Uڲ�m�_W�g���������q\_����m\_����6�^-]�t�x�x�
�<��,.8c�h���\�
u�PB��p�x-�W!�8�S�u�pVP+�4>#!��Mi��~/��\�s����>�^�g�ی�̺c�3�W�U��^1Ƹ�/n3�����Y�j��r�8QA�Ѯp׏��]dА�Ȣ>��ikc]���a?u��c<���"�s������H�6zX��z��'-?K��Ϯe���ݢ�ҫ��`�v�f7�TΏ���A'����US<9�+�#��;��g�>Eq=˺{��g�>Eq���ܒ�Gwtw]��p��'� w���C��!�w�F�������>1P���ࠑY�B���p�z�ic!C!����`gi
 n	��84lF�:���alb�kl��X����5]�DΩ�
*B�x=ii����]�/����_�C;�I$�p$LQ�Ȝ6Xf,,�!�����,6�r�C���M22?�=�O	C������X����6�M*�vc�4�M;9�n\�=�(��Q���z�<7��Yi�Z��+рq��A:<?e���F�ۗu��D�{mu�����!qD>�`����vF�C��<�������_Ͷ2e������8��08@#�Ɉ��ۭL��8���j$xWGჱ�c ��m�Xv��?3�!��RWN��:�v��}j#tB7�CAC�S)4��|�i��_L~mB�/�k?���Q撓e�HM�[�!9D4Pu�)�B�պʦ�d�C�����D���I�f�����L�-��uƥu�C��+PN��ITL%Q	+Y,c�~n(��)F0��W���*�����q� :hht�z���R�ō<���P�6	��3a�-4V������;r�p]C��U
�QnG�]6�l 0���v��3���`{^r���ߵ��	���@��h <�.:c��|0qފ5k,5�v��p`z����i�����j(%sCx�/$r�$����/�����G����C,��(�(���0J<1
�g���!���~���7��(��D��B���M�<�u��ڪh�?&L���6&0�Ǚoё����KѤx#�� �j����]��>�Ds���5׮r��(���x �ώ�D�G�$⳹TZZ�y��]l���IBb�	|�^�{�)����n�R��ppvWVL��C0�l�h��n�;ka��0��A�p��!ho�n�ڧ�~g^oȢ�(� �t>���*��(t9&D���������ݺ��i�����x��E��R��!�r��D-D���T B��r`��lu�8P`	>{����xr{Gқ�e��x�\�]��.�"?���@l�*�Ȋ������c �q�;=�]$O���<mXz�i��>m��i�B?��n��/�E�5�HHH��o����t�jb�Î��_�p666�=�����*%T��!)�R�p�	,1�Xk�d!`t9
e�iu�B�@E��l�	��.[�t� B�7�����I����5�`H^d� x��v���̞&�٣���ұ�O�4�M!C��zG�N`�EJ$\�!$Dˤd.����,�ԕO]�=�i]�D*h��W�p�-���lIA��(�TY �Á����,�.GF7��ۄ�q)ZN�3#Ώ��Qa��(@��p�j�`#F��:zh
�.į9x�d6��<ۆl[c<:pG���&O�9�#��XU�ņ��v�Xq#�{��j}��:�˖�.��r@��3b��K�{�,�6��4V%2Q�;������g���i���Ĵ�3����ڰ��c���B��";�lh�F�.j��ajF� &u$�5C@8�h
�G	��C&á����d`�l*��j����Ϳ&��m=i� Zf(j�~�Lh��41E���ʜ_g�Ls,+����p<b�Q��	f5��EU}wr\*�[x�Ⳳ3�ڟ�/��"h��^�k��m��`� �|�:1���s*�N�4�f0��2�����k  S� as�s/�IeIm�:�[S�5i��� ]��%?��5��(�y����(��c���m���v�g�]�P�
>���G# �ڌC������רg�����	"^�Ð-$�_���f�f�:V��Ǧ�p�!E�]��H�4��5eet�(F(�l2��u����D.h,��H4����q�:G���i�i���r�I��:�"�:1�P��
�G�b���;E��D����,ҙ1�1h�C�Y��7.O�K�	1��䍦g08pō2Q�6~V:'P��V&�3���U��b��UŮ�ꪾU~d��~W�;jb�{^+�Y�qgg����Z^:d�g�
�����|��՟?3j��V٫km3j����{_�8��W���lmx�,�x�^-^>1�Uū��8��E.�8#Q��;����E+�/�\5x��x�8ͯ3�칞����t�4�f/�ū¸^.z���;z�ϲ�[c�����L~i����U�x^/�\^+��q�����b��,<�"�;(���7uN��Z�X�ߺuw��.U�j����eT!18!�l��&�CP��n�d{
�"���צ�����SeѼ�Y(�6ZIX�QnZ2���,B�5�80������.;���\ḍb����1m�e�N���n��{��P��)�!��1a�iϙp�9FRf�(��H�t�YN���Ö*������9�\kD��)�\�?(MrdHXD�S��$�1��RM%`�4�D��Z�,jeb\IA[g�Q$���9��w��"yNɕ2�$H0q�>�-�N6���-CѬ����z.$T>�ĂĄr�
B��H��U��������ʎYes+D�Ib�OY���c��U���1G��e����6,���&�_���/8	�M`-&4�A���"#��jWF�hLE��q4��]����66D��u5H���[�q�5*�MWI�m��]��/u������VD�u�B����֮j5�,N���$�i4�0r*������JF��q%�h�
�+8��m��RmQUKJT�CP��������x}�e�G<����ē=��=�wuû�L�wt�]���I3����ww\;�$�wwOe��p��=��=Ywuø�:|8Ⱝ4�8i��4���_tΖDS)K�)j��RA��z�@�%̈�d�펶��7Y�4 ����ۯ`�Rersn�]v���RN�jz,x�%��?P�+�I�Tn�d-l�%K���i�x:t9ly�la�HN����69���`N�! ��pi���+�hRi��3�i���Mx���nP��0�cO��#��p6@3�7�����t��{�][�V'��jWd�٤b��!2A�����g�C7(�2�S��m���Wm��ze�+
�1�M��1�G����dHi��څ�)s$c.�w5�cs*W���B�E[�.�fF`b%P���]�_�m���62�ݏ��% Gå>d������P�"����2Hhr�t�$��Q��L�dr憜�箮��P��8���m=a��ݷ����T� <3���3���#H1����P��O�>ڲ�	��Kf~4�Hm�(gƉ$�4�v���-�ѻfcf�:Y�@S��{&��_���P�;�7�O]u�U�3��+,,G8;Z]~}�BH9C-�z8`��#�ޝe�w�n�}9��3�f��@��9nc��>� OY�+?j�����WqA��"c?�>E`4�I������	�o�v�dK�3�s8�	�YG��QWjr��GP�i��M�?�������$~u�}�l���,�ZI�s�[���:��F�px~v�zh��á�B�ϣ&HT�|l�|?���iˢ�9��xu�ڔ�c}~r9��jjY�xڰ�tǌV��c����b�5�D��ԅ�^�5�<,2B�#�����v8ol�S��8��M{G�1���H�%��✩��:XTIg&�Fm2�J�����R &��I��DX��4�K50^m�i
!(��8��X��>���-1ٱ�p8)�,����:�X��-�SMI(��.O�6������x�~���Â����)������ɧ&�I�&�����u*l����GD:!�PNqo�w�wy�0O�ff:M�tρ3����ኄ� ��L�d�'ɺ攑Ғ�*�9ع;`�)��w�0��Il���DΞ���%�2��5�S[,����/�{Uj9Pn:�?��=�>��{@���%�	x�����w���\"X��_FO%������aX��Uiګƌp��*�,pe�Çc�����t6�@u��t������x��!�t�!��=:h�T���j��%ߍLԕ������/��8c�}L�>_�v<�W�s���O"�Q�iD�~dC���(O�π
�m�-n��8?G�Bl\��e�4�'{Og��ⰬW��Zv���1���x�������81�A��?�K"SL����O�t]���ɋ*o	�-pT�k#�_���%��69y��۱������-[z�*�ۇ���L4ذV�B�!! �`3"b��?2晍��������&"�鶘�<{~�ݧsoO�V���G#�(wO��$�P�QdS)|�颙\.ce
$!�ʱA2,�ISN:��&��PVcv2�d�#;ak[��y�H�8�X���'d^<�)��r��&x0�
�� �H8B2��	Ј�.�+�i?CE���zxx7f�s��4*v8?n�g��M=��8�ޝv�@ov[��B�Cæ��	������)�3>�ݘ�Щ���,�+v�,M��e2�/7��nhi0CD?�#�4�:Q�>ٸ���/7%G�hC�9`r���r4;�&F���F=����n����3Z��ʛ=2;�a� ��m�oݫeRd	�t�� Qv�#$hx�L� ~ᛘCo�L_�b`
�~lzlv;S��F,v�� ���/���F�G�W�U��J�'���zq�\^׊��q\Wc����>V.��j�Ut�-^-^)��_-Y��f]�Wj��mqv����/��+�Y��+�����~|Ǌ�̶��e�ի�U��+��㼼��8 �G�����G��=c���m�]�n3j��z�+̼g�ӌ�x�/4�W��\=g
~H>��O��^S���p_��^�������������+��ͮ/�3�+L�Ux��KW���?��U���͜�L? ��y�GR\]GP�z��Vcw1g4^��r��a�2Od+��{u	���<��%7��Q����r[��A�����S�]�w��A�7�y>ݑC���Z���W����%����{�TԸ�f$���@>���R�]�GrE	��˝�2��9z�6JnQ�O��m��e�������������y=���Ywwø�:{������q�t�wwUe���������ǲ�c�+
�i´⫎��!m���9|�1��][��;8n1����[�ǀ[2��L�d��9߄6��I�BB"M�]��4�%:>1THdpp������$�9
!�Kvh^���w��r��j}:z�4�XV+��i�B?�Pw?�v��F&G����WЦa�t=��UU�2��Q����2{�5�������X�^�qg�|�.����ۇ��"�,�,+���q�bx�'����>N�'����x5�����r;<|�5UҜzp|'���z�o؝��+�ګO�_:t^�uZ��<�H��!A!�g��]F��\pd�6��"B5���QVww�e,��j�2%�h�"7��岤\y��n�I��ETh�͵J��k�`�b���e���L�Uʠ�I�þӗ�� ��6�?;u�b�v���H]�ˡ�T�����
$�py�$I|L�Âr���?Wy��NŷS/$040�3�d%�*�+MLnU�#��>�C������<��L2�g_�)�+
�v�Zc��GR&/u�X����U���l���Rj@"Ew*��'�9�@tt��U�9i��7əc���N��}0�}�7�����E�5����#���s};ѥg�S�bq=�|O��F
�F�Y�Kel�n��MN�ŁB�F�԰�2�ꢕNͫ����4E�8��He��ݬ�*V�X!N����1���(�|v�c����p�#iTӘV��[��P'UU��ٝ�{U�,�ڒ=m��ׇ�|�zo�~�օc��7oe�{ܗ��9�W��'��J�OEcr0 iAKDf��",z�h���m���8�)f�����p7O���9��)A���Ûh	�,�^�gJ#Hp�.-��7������3����:���BB,���A�o���S*����г��8B�4Qd�Q`�1�×���*�.���o� ��z|`m�~�<e� ;��VA�u�fTݛ̧v�<*�����;t���<y����Y8�<��]���bjp[�F�����#�xr����D0C�DA�1 z���'�ff�4��;��I+N�Ꮑ�F2�ȝ�"�U!J���a��,�u��Ӽ�$!�x���c�Fc�4c%2�j��GCN���bz���:'�ʟ~J54���aX�ݪc<@��y?vC��1�:1��!,JHf�C�� ���ٍ�x�*F���nEI�(v�������IG�5��T�h���V�B'�9�M�U��d�Ixa	�H;"Kĕ�b�|`k�S+���(c��W(��RX=�����FH~$��9s�6?;ht�Y-�٦:����R2:I#�Pt�|�?��.`���fg��l�|���x�Cc���!��p�L��H��rB�:e����n.�V~�wm{���x�XV+��c�a�f�Y*�1f2�߷�;���鲪�*H\�ض0wנu̒UeN�v$���o �n���sWX�>��VC���p=l�	޶]�\�U.|�L����L�p�20�&~��� m^46�@P�k��t���Ə�V���ch��w��{F�=�u��kC�a���# 3���:Oɉ��6����x��l2ѡe��a^eN��r��M\�E��:��;`�'�G.1���;��066=O�����lt9�l�0:�`]8,~#i�����?+
�zc�Ռ|Xz�B�,t49C����>�z|������
�j�`u�3!����p�a��4�WR�k��R�
 �-hAr��y�8�Ϲ�����|9մ�l�~3,�U
+4����Xp�Õ3�$�ֶ6ȏ�"��4~2'�W�Q~*�e�,�L��������1ǹxÄp�.�G�2�Ȱ�T\(�5x���Z�S���j�U�쿙����6rBr5��{�����r-��a����_eap��WKū�8�.�g強�qx��j<D�t,*#�`<4&5����X\��0r6�"����x�W4�W��\/���|��G#h���xH0GW�p��3g�����V��^��_���4Q��z�^�}YQ�6B��4n�6���G9�"܃Q1������E�%�P�R�L�8��.�������?7���Mt��*8k ք�DS`��,��YF"���iq��(��MǏJ2�����ol�t�4ZC̓^,~�e��#x�,+9��ZN."L�h�7�ߓ7y�e8*��6�B,j�R�TB�Hc��a`��{�5�Qx�q�Tm�ךZ�ൟ�����\Bo%���c޺{y!X����Zت�z���$���k�~��D�)�nN���o/�wv*�';.yŝ�_>E䷒�ڙmUW�h�^���ѭ�Ԋ��(���Ը�9U78I�8�^�`1j�A�J��,C�Q����$�E�1�4��T�e.�	��$���N��P�,��J;E!�S���j��[b��q ���18��D�F��Z��;�I$-$�O���W>xѺ1!�-KB
�<��1�91st�>F����7���Z��]�nX�VKJ���~�ON�ۻ��s���]=���U�wø�{����.�q<0�wwUV]��xa=���Uwwø�{�������9�x��V��;1� }��Z:���a�4�cƱ�f��9�LC��)I&���CT��J4=�&�d ��Tzl���Ʋ�K�1���(�ӡ���\x(H�)��LB$�{<��x^3�����놘�rY�Ii��	5$�`t�663�͎��1N�������ߨ�D�نs�HP��4�5��|i6B�#�% �|)lQ1���G^������O��£UZ6����?`���vA
I�'l�x�C1��c4k��>8z�>L�Z���-��H
�r��l�UJ)����xx?�}���T¾1�@O� �˓Lf���&4�'�mp��^7I!?�u���ߵ3?4]��ӱ��N���>[y1���c�CfBpj�.C#�P�;$�J�!�͸|�1r'��n�䆶;�A��4�d�%=���e(��O��|���"i��s��-���6>z��|C�]�uWE�Q���%�,{�p8`r2qݿ>tg�C��1Nc>+�c;$���%Mq��X9h��^9���$RW!kn��,I.�x�Fx?��D?Ӽ8r��s�6Ӓ��g�i���x�P��d(z8���c�d�>$����J�>�}����n�� ``��m��⁌G��4c��?�����(�Ħt��A
A��@���q�!5�[a1�q6۴mUH���!�@UD�m�՚�$�f��b�$�Z���w"��b$��1��j��Q�#(��-���
H��Y�e! O���_��'S�v�.s}'��?J�R�׈INx��sC����p=���vY��O=O�(�>a��D�2���=m��o��w��a�Wj�t�cj}<�s)a�(XS
!�I!�gd�0{ѧ�[����6@�	2�p��И��t��������@�ӔFڊUF�t��Rf�+�X��<�2�&$ƌ�{(þ�ϼ������a8;x�"�0|801����1��UWW4&(z�f�8(̌���u<8kìa	�8m��͏�t���h*�� ����B(����I�-�iD��	�*Sx�ɗ��$�G�$��(��G��$�eG�h�zn"�='C/��]	��Ƥی1�ګ���O��P�G#�A��6�<�{S\��B�F��[q�ܘ�U�ՋK�A���I���O�u��0J��t�r�ǣ�.&"����!��Ε$�+c���CC���n��Z�=m;��I�u<z��_��1[Ucj�[T�����ұ�:U� 빹J!a�+D��I=�8�]U;dN��	r���ƪ��N��`��N!�8�F8�1(���f�CdU#f!+,eV�ʈ�3LF#=�|ۣ�*��׭!C���öFB_�,v;>~˳Zܦ岡E��~C���3eNI.�}Y�C|�c�ΰ[%շr����$����Aֆ���x}G���0�+�V<R4���썡$� ��!�c2��0:��d|�|hL8(6�[�t:��=q��Wvr���IFk&�ɳj��U�����D��>�x>r6����C�>l������"�>(ُ�U�E��rE���d �=�c���ǃd6W�ڞ���������qj�j��W�U��o���|��+�3�+����������8���ڽ^/k�e�\Z�*������q\]8�;��<s-��m�<a�hhZ-�"��ph��gv�q�^>g�1���^��3���y�q�2�ū���.�����|�=_e�8Ε���K��U�x��8��qq�8�^/~U^F3$0Br4�!���6�w2I6kе����d�M׹�<���O�Jq��[m��+o8���&�X��L�-R�"�s����fю���_r5�}�]e�e�ĕN�&�:�'B���������wwuUV]��'����ꪬ���O=���UYwø�{������q=d���ꪪ��ܷ���1��Uq����/�J*v�K�+"���=y7R�ۡ�g��`\}i�?�L)���{�p�[?�'�C"(�;-�F:GJ5���>�`d-��^�a��8���t�S����ю.��7)�m0�+�V=Uq����gHt���y,UО�=:��S�y��n��[$�zh����06;��w$�>��:<
�|��m����
`׼X}��6r���i�����mU��^<�o��1��=p@�"�&=4M���U���B�ML��C,-%64W`��>*�͙˱l�Ǡ�k�qTWI4�q�z48�X7I�c���4��1����������������U�"���TL@�3�t΂�
qӥMsR�ū�������6�Sx͇�I$�UCd�`N�G�������.�L<׉R��i�~��e<�5�bm����T�Չ(r'm�ضŚ?L��rv�����a�Wj�x!��tCƗx�M0�ο¦pҖ9�$��G#Cǣ��$�R����C�y&��E��n�x�F�������X���������1(��kC�Ҧ�n�l"�\��C4������?49 ��C7���cgͰ�+�V<Um��߬��/��1��K�5%��p� �~|�u��$��t�u�Gp;ߧ�}�B�����ؐ4>�A�?4�c��Aâ�&y�@���#���+$���d�(�^!�>�z/�� F#�z+'�b}zuz�i΄��,l���&{!&6��8�mG�����*�<~���VH3~����47�(���M��%��#��ӆ����jJ��X��6<t4ۦ�<��C��$��������HIUGD��ꊣc���y�Og���}Ǣ�Q�ұfΔ��ګ*��45.���`���+b����S��KD�,�HR�d�+�1R�;(��4:��H[?��ֹ��+JRW�K:������d� ��4Z!�Q
̭�]���&�8�;����u�Q%U5�#φ�Ik�y�<x9x<:8�;�����y���>;�l��{�b�̷_��|�/��j�Δ.-�G&Jq�$"��S��\)��ʦY���'t4=N'�^���f�tz�z�ʬmU�C�l�%�P������C���L�8g���$p�prSt?� ��F<,3ܙ0?4�W�Ǫ��g" ŐDDQ�:QТCq��.d��vd2<��C���o���7�s�ĵ��Y�!i�L:1J��UX�U��'�\�fQg�����Ɓg�G{�x���_��	�Ä��!����3���:�f�#>����G=�V!�X�qX���T\�8}	&�Ã��`<<�ν���:tПm���6:��}=Ӥ�a��ںUc�W�*��pХ�"k�A�0�ՈY��5�I��;i�� ���!��S�+���Z�|J��Fy��&,8��xpx>��	�<���\�.&��Nɤ�M�?^w���0�z�8ڭW�W�U�D|GFe~*�0��8Y_�<-�gیq|_c����W����TZ8d\(�D\*�a���6W�m�*��~z�˧�?/K�_���8�����+n1�z�]ʋ�������#�X�H�1��\\'4XXD����࠸0������<4,��8Z&G���< $�x^-^��<W��2��e�8Η��sK��U�x�x�\k�Η8�^/~U]���j�_!#�@��sw�RҬ����$X��s&�	��e(�DM73G��JA�EQ*�<�X�Zk��Dj0�k�9��]\p�����.9�q! A3�v�(y�P\4� �� ��Q��4�%.��Z3D!�x%��J��9{^�b��臍�ee�5������c�SX�
JHn�M�JIB�l%c!QF*��c�Q��eP�1����,^|��hX�E(եЭDiyd����fFS�������h�2A1��ߥ��3P5}��P���:�+��4N7JwtSG���3j�>g,�m��4D��Z\�h��[&"�[m�U�k���D����Cѡu�hݒ��x�'Yk�l����U-��tm��9Qc��^�n�蠚�A�^݊wu]OK���z�MNA��F��Z&��!�ĚגA��ƑD��M �I�eq�'"����Z�ƚJ�Ui�(&F낱ؗtf�tcHN��[Ub� Y	F�q�;I���-�ʪ��|7��=���UU�ø�����UUY|;����337�;�����33�ø�����33}ø��G�p������s�>�'�GR����(�H�3Fd+r�R�]��
�d')	����cM1	ܱ�H�V�"�Ѷ�␻Ri���<9dMV)��΀N�4TX�"���,��%�ײ��(�CC�<s���ducC�i�F�Z�{���jo_g�C���ǎ�J{�I	�������G���L�2��'�b$n82�y���/�4t6����1p�.�%E�Q~W��z��]ڋ:��d�2~:6=y��͌����+�ă������bg��M�Bl�q��rI!!H8-�z6�a����t��Hh~��>~��&g�PD�>�Á�+�x��ʯ_u��/����
��EV	����o�c���Ȩ\��W!�(ꤨ�UUT�%��<4��Ӟ�/�OJl�6dʐt:4��$��x�ވI����t���R>4�i[Uc�V�߱���K�Sς��>�(��RIp�/H�N1��y���ѓ����^�X���e��c��,�~�M�Ӽ���.盇Uߡ�.��>g�n7�`����Დ��hc��rJ-����6��U��uVtvޜ�N�9���9¹r��p�
a��!���N���V�����q����b�R�Y
�TB�Ì�#\���&2��F3HEJ�E��]VQ�c�`qڟ�9^��cQK�ɉ��e�w$d��y1x�f�zz��k����������a��d����c$h���[OC/Y	%�v1�������c'�?��(���>>x:��;9�Ĭ�3��Ƕ]E��q3Y2d�=Z*���!&����)�c���&��&?|�kmUώ~%�v۱���a�&ps2�J�oL�˜���b_�%���"�'A��bT�E���g��4Ι�u��C�����,���'y		-�<��N�:Ut�qOX�ǌ���$����<q�L
��MPY�*���f��49���ს�;�Dd�j̝FY�n;a���2~���h|#�C��ȣ�J*��X;��j������~f���}�f��=�s�M��ۈ�S�]M;�Ֆ��D��������m�V�S:2U�b��Ps
b
5j�jr���r��o��m/7�&�������8yOg�zʵt(�QJ�UC7�3�r6����B�
s�&�.jcu�W��
�lݸQEʌ�͵�b��8+TÚ�;��vc[zN�O�$P[�H�F��`���W�r\�l�ӱF�3e\�m(6�2�Ƙw{WYE��d7-ε0��%�چv�-���I��p��[ý +��6�T�Y�|�U|�v���aꋹ�<�]�?j�5�T���
R=H-% -At\�!
}�;���6`�5���c�7 l��$ch\�p.U���4�Ѧ���Ɔ��<f��:�P�<���ّ����ǣ��	��5<[_;N�])^����|2q��H�
N�ơ#P����E+(�bc�+@�ʋ!]D���B�)Z��)#q8ܐ�q�NLIђW	J���q'RU��yUD'1$��"�A�b��a��$O��
A��A,�D�2<�c3�1fi-���$S�23�����P��|<t`�UR��j�C����%o|<�|�!��ЈX��������:<U���6@e.C!��Gr�dD�&e}�����.軻�`�rttP�ܐI`2����0%��B��3��QTWD���vl~,�`r;w��cGW]��E$�\��9��C>T
0�Y$���iӭ����>��O����jO�xl�����+n�m��6�[_m�_��Ҷl�f͛zq������x㎜qӎ<��}���m+f͛6�m�M��n�v�o=m�ͱ�ǎ���o^�m��m�o�|�珝���m�1�f͛+�m;m�Ǯ�v�mb�lٳf�l��m���^��=]�Ntc�Y�[���=�Z�P�]��l�8F��D�q9�O@.+�S�����9��M?I� {P}\��u���A�o�]�pFqT�j�� �)�����X湝�|�˞���/���S��J����Ԇ���d!a�pj��� ^��hh�0���{�nn���cDK��+2�fe�0oИ�;��ff{8w;��ff{8w������{���fg��q1û��fg��q1�pp@�c�����X��9m�^��$g񖆬r0OG}~>#��8�k-�%�p,I%��3�?�-�֛x:��ѱ�2��*��|�<�������=xy�Gѳ_�=�m*zW��U[c�1�ιzr8�G���=�(��3�&�1pIn3���3�ԗ���W�e���]�����m����m\���t��2:#�L/c�����d��!����r0r�Em�qU_1����\�.���2���!�N��b5�`�dv�ɦ�c���3Wk��&�+ �yi�sF=M7q�9��rh���ɤ����V�6��X�r��%4u��rV���|���h!E^R5I+�U٢����4Iу1�wP�v������o��>�UR��1l|8�:uzpp��jUO��<��_濒ܥ�2�!Sq��<l�G	e��%�E$K���x��X�᝽1����t��Q�{��\j������y�離�08�e��!B���r��i��*��<�	Bfn����iU�����Á�P�{�=<o���J�ٳc4V9F��i��FG�Ӊ�껶�v��J��½UWL~(�����U�U�b`�����ü�>�졃���F|�����e�|7��������c��n�v~t�nG�<|I#
r��lv��Y�d�U�c�U|���6�W��x�bZ���+�lݖo�;��q�UD��gY�1w'����>/���F{�Mx�[.WX���B2��=���I�ʣ�m��n��pg0`m(x�]l��]]�e�G�Z���wW:e���h(�,cpBњ1�齟bX���"�UR��䰅x� �J�J$V�S����y6�b�Y"�&GJQ���%#sc�H��&�Ѯc�T�%x��M
&"��J��2�0�@LZ�F��KF�#$&Bd�$�d����>B�0�❑�٣�~>`�����69��wI�ӡ�͔ʒ�&ݞ�Iax�Y?F����C��hׯ�oǣ3��E0���@�U"���!#���,Y����\LMU|�⪸�%Q��o-NY��/�ս��{����hy�ꮇї�ņY�F5=�*TǦ�õz��_c�T�Ι�#�A�j6"�F:Ħ�
pLQ�0:�H�4��w�2�x�c�v��	���Yt`A�� CC��CQ���L��n��0�5s���.#�dޔ�oc���������xC[ �j22MN^��_<y�G�VY]�9�F	�;��N�GOG'�M�{Co�5E���o��{:#D!��3���H�E#������$�J�hi����z�d=���~�����)ե,;&&�*G�ZݺY�ĕea(��:�?n�U��ڦ����A�#�,BʵrH�Y<�P�ة�V)�u���7������5���eUQ%0�\��N���u�1�^�?�<W�Vݵ�v�m��޶�;m�lٷJٶ����ǧ��U��qێ8��q��i[6zl�j�n�v�n�v�珞������O��o]�m�;m���6���m�i��b�mڶlڼxӶ�<z�m6�lc6lٳm�b��m�|z||xB7���#���C%�|��ܚ*�h����Xvz�#�<j�|�m���T�:���HsN����q�����p�|ksQ�ۈ�t��9*���5>��t|���1p�U
A�i�*7)Y��%m.�&Q<*	7�a��Ò3c �28(Fu�R�\�p)T�Da��l��u+
�Tpk+�"�*��p�sx��(;���i��ҷ�zv����8�LU.{�k�[��ۨ�%�\�T<����}��w9��]��6Z&�{l�K5��틊�yK��5�Gd���.�6���n�n��F��&�&�훦��1��$�/�i�J��s��L}�J�b�ƻ�{��$�\�j�o}�~�9��;�Fv��/�m�i+y��:��(5fNC|sT�7�%�^k6�Gi-S��8%��Il�J��u�7�FT�5"
bX�%B+��6<��V�lt���i�᳋RI#H��i
�&�n&��]u�)�^Tǩ<MV�IE1DD�7d�t��(H!P'�`��ٙ�������33�ø�����33�ø�����33ݧ������33ݧ���=��33ݧ����+qU\c�c#z���N�A	�Q�Td�Z1j�0EDGH#�̰X܄Ț&I1J�	�%z�e+du��Jm�zn�(�Er�Y��9 җ��9h[�v�X�$�Tcd��������+�K���|����z��^އ����$$�Nz�@`�4:�����Fq���89>����-�PF�s&�HB�\��<N�53�������+z���d�!q��ĩ�M1p�P� ��UJ�=R�1��D�Tx��4G�Czi�nYlu��C��l賹��� �k�kn��VD!��{���$�~���Ǒ�g.C�!$�{�8�#G�0ƕU���8�'Y��4ak}#048�����|�<*dxug�?��=�tщ���k|�T��bC��8?l|�*�q�:*�1·~	��y\�7	��'8���7(8���FGTN �ZPD
 @�c,Cd!L��/p�3:��Ђ.��C���HF�3�ϊV	5��h�[��xbh���>��th��/uA�z�U����4$�x?b���8���2^;�ߺi�Âa���0?�ǌ��i�h4PPQ�G�h�3��L��s�jĿhɢ����Q�<��яZ! �oM6ZBIc��[Zٴڝs�'7[,$�#��E��N�5u�N(*�)�ڱ�D>H�u�{�����d�<�i��]�����h48�\�n[*HKn3/�j�09��J�z=p8<�á�n���L����3��:g3���U]#ih���"�R�7q��Ͼ��S]KmjL>a�<UWlm�c��T�ծ�����c�xa�&q��<��\l���L�b2�>)�7�]�~����E��n~2grgK�A�Y��{-�����mG\��e�2(Ԅ��Ȇ���|%�&�c�\L�Z�p�tc1Ҫ�clc��=����8��Iޒ��yh�<9۰.o�1��4^	/���a�Um" ���>3�30a��MU2��Zr�xlx���g����g�GɆ�5"B_�׌��8�����	Ԕ��Ҫ�3��3Ǹӗ\�\m�3��T����Z�7ׯ��	��c���:x�F5Y!"��9���D�6�� bΏ����o��x��}"��\=�llj?&}������e���X�g��`��#��h�t���q�cn�J���t�JIk&q�4X�ħY¡��T�Im��E���1^�^,m��
i�4�ՂTnY%v(�nV2�9��["�`�SCO�t��:h�6�.[8?=tg1,lt>��)��qn6l�p�H[+�HiA�d����EH�ʄ����������A�����ێSG�0��U�c���a���w6�py�$���e�vԐٗ<Sr3g�=�g1�W<7J)	.�c��{p7;'����%C��`jʹ���rz��3*��s�vO�;��ߨ���n���=w6�6�<����i�����릛m��oV�m��m���6tٶ���������N8닷|�8���+��mZm�M���o|����|�;i���m맭���;m�o^6�[v��m�ٳf;cǎ�6���m�i��b�l�f�Vݴ�A��4@�4��F��'�D��"�,2�+B:`�})�x!aH�[D �K	�	���[b��w�"�Z��ݱ���YB@�ҭӉ[u��C(��F����zu1��{��fg�����{��fg�����{��fg�����{��fg�����{��fg��q�G0�UW������s���j�U���rpv;=��1aM�̹QE,�J���L*����C���颡����O>۟6�Bu�n9��;
8N�����/Ggl0�J���1�|礩������������	R��Q*J%T)�T�D�#N�Md(\tt�GM������jJ�48�#/���X�LNt�ׯ�K����89Ѻh�+ñ��u��>N�0�U�1�q�����ReS�mDX�R,c��F��<T�2�!dJ9K�$-f�i�D�K�\q�����V,ي�-J-{j����R��"&�EIK���yD�t4�&8`��c�Dk�-�gC���}�������\���xo#k�lv$������m�>&ܺ��_v�f���g�\&@Q6�5&CA�ri/�w��o��a����;QE3�r�I�����x�i����y�s���㑢YY�v��٠�T��}Z,`�l=�o~,.�W�<p+�ŧJx������nLصH�1�E$�'<}�]s!�,	d1��t1އ���L��۷���#�4c~�~"%�ils7�s��<���^o5&�LY�Z.��o�䧹dt<6���?J�$PG�JXB�u����!mw�:$�nS:7>2�bEw�pĲ�~x=����V���F��k���}<8�<б����*�ќ�{?s��t3��i���&%�1X�&�����v55$+\�%�r���4��Dp͏������$���CF�4�BJ*�ۇ@Ƈ=t<&��뫖�r��C��\���wg*�Q�K��V��_M�:a��Xh���D#F|1���W�ߝ�Y4���XFi8��,�	�M�e�X�sJ�7��]$!��	V]Kb��N��,�A-Q+֘	��>>$��mi�O���BƋqR��
� ���p-�ZG����77�a�f�}`SV�������GC������oJ0B�nB�$��m��둒���HJ�ꆸk����l�.>K��%�����Fyy���� �C��J�2�Děu9]�EtD�dd��x��/�I������m���a�*��x�1��&�Uq8�<9$�(<_�I!���Y�8Bd}����C���>ӂY���G �Ay%�˓C���z�x�	a��P�v����>�U	?Á�уQGHd�!̸(��������Pܪ�Q������;�m8M����لD���-��TX��Z2jϱT_]����<$��A��Ya��3l#0;��.��H`��!�φ1�u1kf.~��Ve��������rm����^tՆBF���9�2,}�G�%I����&�_'�C�6G#��`p�lc��|'��E����%Q%�UU@ȒI!��^I|��g�`��[>D����B"����B�t=_������4�}�PDOS�u� 6����@�	�$����B$	 0$�����\tH఩
0�$�(�"QP�$0XIE"Qa%�#P����0�*�����G �IB�+0����*Q��R�%QR�(�#�QR�EJ,�Z*Qe(�#
*Qh�E�T��R�E�b��QeQeJ-(��(��)�R��YEJ,�Z*(��(�a(�E(�E�T�Ģ�R�,5R2QJ*QJ,(���R�EL�zƦ4F��%(�TQR��Z*Qi%�YE�YEJ)E�(�����?ቂ�,���
*Qe(���QR�(���K!0�L�C�!0�L
��(�E�YEJ*QaEJ*RK(�E�T��(�E�RQR�YEJ,��YEJ,(��)%�T�
,��*QaG�0YI,���
,��,��YEB�(��C0�L*QaE�XRK(�E�QeQe(���Ih�E��Qe�T�,���L0!J*QR�J*RK
,��QR�(����T��00�C0�00��#0�0��2�0C#0����*QR��T����T���(�EE(L0���L02�EJ*Qe(�X5Ah��T��h���Z*RJ-��,�ʖC3�2C0�0@QR�J���)E,��,(�)R�R�*R�T���Q*R�XR�*R��)R�RJ)R�R�*R��JQJ��%JQJ��K�J)R�)E��RR�*�)E*R�%JT�R��R�--Xe&u����J��KJ��T�E�T��J)e,R�*JT�QJ��J)R�R�*���R�R�*R�*JT�N��*Q*R�T��J)iE*R��R�R�*R��JQJ��%JQJ���)d��J�J%JQE���)b�R�(�Z-,�JT�JQEJ����J)R�R�*��b�JQJ���)R�R�(����J���)b�R�T�RR�*R�T�)EXU�"Ȉb!�"��b$!HbH� "b��b"R�&$�%�"���UUJ���aTR���!�b�"!����b��b!��!�  ���IE�,�)�d
E �Y�% ��XXD�!V:�iR*"��JE�R
E�%"�)�"�a�DR,��R	"0$"���@�	�$(@��p%NI�n���_�._4�)����?8��DYDRaP*���џ�N'g�>g�����j7�WĿ�/�����]���?�@��5�|�����V�j�ϻ�Ҳ���#����w
͋���Y��C��ݯ��Sh�R;�ڲ�z:�I!J]v?^k~�=���p�O���脁���2PI!j���� �i&�/�{Du���{�7������%.ⶁ�����\'���������^=i� �2|�I!�D�����l^�!]p �Z	�('޲�C�[��8����))?ܜ�F -4�~��:��O�S����j�;?�`e1� 0?����f���b! uB	P��TT�<���U@(D@ܪ�����a��!��nx#��`5�o'�����VS��˟��i�i�)đ&QU����U!=�$�YQ���P��"6����y�� ���Ջ_	�z�9����?�C�^`#����P�~B���W�b���1��H�������SsnP��CUQ-<0eԽb>c���������xh	�
C�=��?�?������S�?�S�T��>���^p=}��{ǳ^w�`���{�I!���)�_���z����+��c�S�v��T2����( 
a���DUQ?�����_�|%�����{�+����`��W�:�q|�ѱ?����Q@;z\�
������$���G𥿈 ��@�ۣ�D�9�<�L����Ji_�����DG��|�{�?�����-���?��G�n����0��y�,d����3���~�*����c"����L.�J����?�����u�:/�"w$�]=guG�/Px��p����	�@�Pď ��k�^�����ÄUTO̥���S�V@���������AM%AIAACAM%%IAA@P�CCIAC@P4�4444%- ����S@P��JSIM@SCJSIM%%%%4��@P�R�@P%4�%@P�-@P�P�%AHP S@RRP P��-@P�4�-H��-H@P���H-!III@P��%%%BS@R����-%%%)IKM%%%@R4�RP-%%4�RP%II@R�-)BP�P�	@R44%!CKC@�44�4�S@P��@�IM@SCJSIM)CCIIIM%ERJP��4@P��@P�%-@P�@RRP P��JP�-IB�-%Qh�E��h�["�h��CJRRP��%)IIII@P)CIIJRRRR�������H�II@P�M�RP�����KB�% 4��������R�R�R�R�RR�R�R�RRRR�R�R�R�RP�R�R�P��������%AIKIKIKIM---%-%--%%%%-%-%-%%-%-%-%-%-%4���������%%-%-%--%-%-%-%%-%-%-%-	E-%--%-%--IKIKIBRR�R�R�R���R�R��4�������4������RP�������4P��%%-����-��������%%-%-%%4���������%-%-%-%---%IHQM-KACCIKIKIKICAIKIBRR�R�P��������4��������%%-%-%-%	CAIKIKIKCAK@��SEIKIIIIKIIIKIIIHRP�R�SCCCCKIBP�����444��44����P�%%-K@�RRRR�4����4+I@"ҁCEPPPP�P�4��P�Ҕ��M)M%4%4��SCBP��IE4�	IM%IM)AM4�IIM%4�KKK['�?��J}����������B��I�?�'�|%�C�k�`I%��r1������`I;&vm޶J���������"��'�����_�ȝ���,������2"����9��E��ꊩ
`����?��"����_���۠�W��x�?
���H�����P6��H}FE�#���!��������bC+� �����S��D�O�CP;��ƗO�=��4������ϟ�o8�b$p&	��G?�]��BB}�