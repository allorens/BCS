BZh91AY&SYa�ݲ��߀@qc����� ����bLO�                  �� ��Y��[T�ج�U��Y��Zj�f�mMA�mI-dض[l��6�Z+R�km6�������RLC$�ͭM�L4*ڬ�yb�ڵ��F�36�km[��m�)�)ZQ�Ui&40��Y��A�5kB6kl5���2��W;Q�@ R�
 #��цF��p ƫZ�N ����mdn 8sF�k� ��l�
� ������e�C&�Y���Vؖj�V�m�lͻ�q�L���G�RR@F;����u�۟`�W���V{kЁ������׋�W�]Z���������o5���֯CUt��z�F�ws�w�������6�cjm[6*M��)H�����vj���Ow�YR��ie�y{�J
�U�ږ�=v�{K��PEt�ח��Zh���;��P�������a��<�C�UM[=��_>��(P�wx�RUlT�YMfmJ��|�J�w�Ͻڍ��q��A�X���z��B�:�=�h5�F7���di{j]�t=�W�yޏYhP:�����5F�}�ϓ��Ξ����z�F�����)�W�NM�Y��%H =�}
ն����=���hR�[�[<�=TT�t���Zi��]����Mj��缯Zh(<�kׂ�P��wm�
�z������ �g�⏢��x��%��5�j�D4>I$� o=��P�c����I��z=J�R�O\{f������o^�PR0�誯Zh/�Ga�u��j;�G4�qUT���Gq�w:(�FT�;�m5��fG���H ϵ�ڐ���@��o� sm�@��� 7�AT2]p uK����������zxD�������ek&��)$� �C� ����;��@����� w�m����j��: ��� n]�@� ��w�>�A���U��kI��Tɦ����JH ��� �G{ƀ��=� ��  ��p�A� ���C����������; ����[Y-Y�ImQ��� ��t����� �l��@c�=4�}on�z �0l�� }=� s�nPh(��{��]S+JQ�fڦZҒ��V�7��IB�����Ս� ;����=ztn��@;X�+ٽ��/]A#��x:�`(���|} }AP     #@    ��2R�#)�j6�FF ɡ���1%*J� �   �d�SɐRUS�2�    ��
JR�C F#L�M0!�3Ԣ@�T�       D�T��JL&��Ljjz�H4�)��~��O�~������e����B���6��k�U[�n��x�\>d>=ܛ�~
 
��E`� ���W��?��������v	�G�����������q�T�� U��y$�K�� 
��@�0(D�bv@D@�����_���?L�`��1��u��CX��5�k��b�8��.0u��X:��.��kX<`��.�u��`��u��]b�X����u��Mc���.�u��X:����MbkX:���5��`�kX����b�X��15��]b�X���&�q���/:��.�u��Mbc`��`�X�u��]c��1��Mb�X:�5��]bk#X��5�k�.�u��5����&�u��bk �k1#`���5��Mb�X��������u��X:��.15��bkX���&�u�a�bkX:��&�u��bk8��0u��]`�X:�5�k5����.�u��]`�X����&�u��]bkX:��.�5��5�:���5��Mb�XČ]`�X����u��`���/��5��]b�XcX:�8���:��.�uレ�Mb�X������N1u�kX:��$a�X����`��.��`�X���.�u�kX1���&�b�X�Mb��0u��X��M`����bq�kX����H달`��&�bkX����k����]b�X�b� �.3X�x��.�#X����]`�c:��.�u��b�X����`�5��5��^1u�kX����u��u�:��.�u��b�X���5��]b�X���.�X���CX���.�u�c�.�x��&�u��]b�Xq��\b�X����a�`��X��5��`F�bkX��5��a�H�5��]`� ��u��1��]bkX:��.�u��cX:�5��]`�`�k��5��]`� �3X:��X���&�`�X���F�u��X:���`�#X:�5��]`� ��u��5��X���.�5��#X:���u��]`� �.�u������bkX����c`�u�kX����5�bkX��.�b�X:��8��F&�x���u��`�X��5���u��b�X:��!��X:���b�X������X�`�X���&��Mb�X����]`�X���������u��]`��Č]`�X:��&�u��d`kX:��&�u��Mbk�5��Mb�X:�5��u�`��.�u��CX&�3X�0`� ��bF���u���u�kX��`� ��u�kX�bF�5�k�!�]`��&�1u��]`�X����c�X����5�kX����8�`�X���.�u�kX��5�bkX�u��b�X���cX:��X:�5��`F:��.�u��`�X���5��Mb�X���&�u��bq�:���u��a�H��&��M`���u��`�XF:�5��`�X�b�#X���&�u��`�X����5�`�X:���u��M`�Y�M`��bkX����u���&�u��M`�X:��\��.�5��`��&�u��`�c���&�u��bkX�5���.�x��&�u��b�1��M`�]`FkX���&��MbcX����u��bq����b�X:���u���]`�X:��	�]`�q��]bk�.�u���X����u�k�.�`�X�.�u��b�X:����]`�X��u��X:�5�k�X�`���X�q���1u�kX��Md`�5�k ��X��x�X�0u��5�k�]b�X���1��]`�X����b�5��]`���.�u�k �!�X���.�u�kX����b�X����]b��:��CX�b�X�f�u�q��X���.�냬X��5�kX����u�`����.�u��c�u��^1u��b�X�1��Xc:��.�u��X��X:�� �!�Mb�X����/����b��u��CX����]`�X���u��]b� ��]f�cX��5��CX���.�5�b��.�`�5�k8��.1b���X��1�k�/�Mb��X�0X	��`�0� ��GX
�]`�k`��Q`�Qu�.�b�(�X"� ]`��u�.�U���GXc5�.��b��u���u��@5�.�A� ���X*�`#�b�� 5��X�5���`�X����5��`�&�u���u��`�X����u��c�cX�b���u��ckX:���u��]b��8��.�8�5��b�X����5�`�5��X�Mb�05��b�X:��&�bkX���:������]`� ��b�#X:�5��]`� �.�u�k`�X�&�u��X��#X��`��.�u��]b�a�]`�kX:���u��X��`���u�kX�b� �!�u�`��.�b�X���.�u�X�x��.�u�k �	pM`�X��5��]`�X8�X:��X�f9�	��������w�B���H�z�KN�Q��f�f��ؙ�.K�fd����8݋m��pJ�5;{!PP[��̎�[�^X:1Q�%mi�v�#=$�1Ȧ��ת�Kt�p3p�����X�nfI/!�����0���J
m�7B5�t`&,�(�]�&�
韶���SV&�{�jŊ�ٚ�:���Dm:mືn�*7�ưD�m]�@�cn��K����� �OYvE<��-G��;�Tm�7ST�f+n��4uʰd�������N�ŉw���2������ؓT��Y�����{c.�h�4��3]0��Ij+�c�£*\+1�	�l�-���kt!�ȉ۳�Ѭtȣ Q�m��L��Zt�]n%mL�N��1L���j��d]����GfԼ	e�����6Ű[Q�M`l�ۊ�3&����e;��E��9��������vȺL��R��Ԣ(�wn�8E��u�̺˙1�ݻ�s(B)*v$�6��0f)e9cp�NI�J���CPL���t�ɡ�� ���٥ڒc���X",��I�S4l�uGp����j�Z���+P���c#�5P�� ��7�f���p;�Qh
j��$���U�G�l'j��Y��\�N�d�o)I�&žlԥz2��V8���hn��t\�`嶵+�*�@s�� ɂ�YPڹq�Y�VDBF��V�-�T��4�8�M�,c�N� R�VEh���e��8�j�m�H��-�t���S��*�zƻR�t�KeU/=uJ������X&�n�m-�P.��Q�����f���3��h�Lj��Y�Y�\�hY���l,�E'%�H�ݗ��5�ۖ�"��Sp���%&�ͅ�Գ,���݅҄Gpl�m6�
V<9V7)jI^��^mh�[j�� ^�{Z�U/f��=٫�wL+�#�BL*ZQ8�t��B̚��f�I`*�
��uv���}��P��r�ɉ���ʭb(Ɯ8n�[�V��M���'yjܳ.��HpЃn��7��wA��u܊�I�1j,�x���;��Nh�͇p瘝Xx%b���6�AĲ�M��/}E�/7��ZFcz�fަ*⛧ �p7WD:f���q�=*U�kef�XE3�n�7N �͌R7��j4��,�c	h,jG�����u�4e���w�o	43䱂�[��Q�C(���d�Os	M�������c�����~�z�V<�'��taxw����+fP���ul[�����-���W�Q�����b�)C7^&�o)�aU�t�ͣ�(�1�m�+��:������1s�K�Ol�ݍh��8nBX٫M���1����wRW���Q��SsrL��	f�rA���l�۩��+�-�D8�܂I'��j�e�j�5gH؝���ce'pk�f�"P���a�5�[d7�Z�-z�v���dLc�y���=�e�]Pvױm��ډ�Pّ�ǤRvo^��4le7I$��{LF�B�U�X;ɵU�%�Bʋ\Z�R˔7
z�h��v#�ݸ5Vix�Jބ0e�~p̰Q��?c����x�D��MF����˺d|��q@��c͹j��\i^�h4�ib�j5`�y/[ ��,�%�u��Eٚ�#���t�Q��K���̢oR�F�:�O+NT��ٵ(��y���ס:��rm9��cb�.�ok�r��IY�r�U�`��ُ�[<���9L���?Jͻ�P�7un�����e2�k�HV%3�!d��e=sΘU���b��j৸�*jMei֤�,�V���ū�TILhf�������iٍ�z�	O'vY����we(��(���Eݘ��գ*�̭�NU�2���T�ܬ����O#��X��{b����ԓf�sat�)�Q��-��Qk�S��t;dS[`�nz4�/[o]�8-P%]9�l/du6����sJ��h��i˕E��x�/o\0�,�*:�.���0f[Jː�.��Ɓ.ԭ�n� C(l�l�(�٬�(d7����5{v�֘�k���[J�X�d#PD���l-JA���8he����Xc�䗚�3Y�F�0��n̺YZaVkYܶ�L���qR	a8��(U�^��G�,��.���f8�,ŀtDP�i+H[$�n�\*�" ���.���mh"홦��N�ҽ�A�����ͷ T裲g�i�c8H�AM
�f��ȍj��Bϳq�)нƒ�]̅���
��'�7NJ�\���ةJ{0d��\�6�)dVB��d����ۺ�ۖ�]��y{�0�t*n��cXQ�fm8�6�TcZ�dTU]���7V3v��X�y{#�W��A�q�4\�u�t�]���i\�)��vВ�G>Dׂ^e)A��.M����p寖D(�!
Ć�v�V����m��Fܥ��e'yj[Lֶ�;��`m�B,�5[�m�.�+�iխ�m�Vud�v��.}y�𧑆
���	t�����
�a��&c���
����Cpi��l���І�˶��`Z����4�ϲ�s\j�*�"�۽���P�^��Z���Cfҹ��$;`�W��汸�x�)#BB�gS�K�-���[@�ͺ۰�Z��jM����I�Yaf�P�ez
��$�6�,v���lҗ�æ�U�5)�! �V�nh%bv�b�ҥ�q�%^*��mǹy�v����+��nVJ?��{{
kY4�y�F�Bd�+4��Zq�w���2�=օ]]
g3en�[�x��m��#mM��aY���ߌ�l��r�)N���:;[w����cW�<�R̙bf�{j�n74C��ə�V�&�d�f�j�!U+�n����Rl$rb�/,�r�E
��&lH̔Q���Zu+r�c��c�KE��++M��#z ~��`�0�:e�H\�ӋXb��E�w!ݺư��V��	�,�S�Fx��dA0��%Gga%�� ��VU��d��:s)P�v˚��o`�LFj^M�r���0���"F����f��-4��X/#S6�lJ��Ჵ^Ҋ\���\{J�"�7mI�۳�42���Kww����DT���R���4�CFLR��R�mZ�s��uM:��+^=�f�u���U�`�P�!����(�6UY$Z���J�*�ܼ�j�qr+v`J��Zh�����ږ��8��2mD�D�ڑ`�̖�L`4�5����yDf�H(`0�)=r�V�=�Wq�+<�ugC6K��[��%���I�"\��Zv��H�3m�ƚ�ދ0[���		��+!�������̩�u=ϐ�%�Ϸ�nf	�"�J�*�t�f�����"�&z���P]E��&���^õ&�%����H�b�=!��E�K#ݫ�ln�Q�dn���,Sws0�����Rإbt��nK"����A�೰+�j��͆�����MR׳\�b�me1���r�X᷑,dZ�QP�&kN�r�[Xf	h�۬Ǒ�I�y����!""��R�d�Y� ܎�"��T���;a�ܵ�e��=��i�Q�V<b��ف"��-���(�og6�T��f
��L��7	pͨ�vF��r�Ť�m��70f�ͭ�"�f*jt�]��sPʲ�X$���Y�`�t�+[{���S\Ƿ���[����&8�4��%V�*le��i�
��[.�-V�Zd#�f^�\�1mf���Z� U�r#M�d�d�[xf���I֊��mdM�7pV6�1׳&�Y�i�H'nS���I��X˕#Ӵn����Yʂ��pn���`X�9f�]�y�N'�M��E2��`V�Uj��g���i�z��DM�.F�ɋ]�Y�"�	V]Z������7t�j6�nȈ�Vɛ���Z5z�	��v��X�ǵ���lFV���F��H�i���Q�����L̡{���E�Ǉw� ݡD�7$���J�����ula��L����W���,�v32��NP��r�j^�G�ji+H9��la�	;�М� ٲ#x�+3Q��RD�{ZLsF��ku���Б��M͎�5��),(	qP.�{mݷ��6ȡL�݇�:��w���vM�.��X$�av�,�F�­
�ہ��)@�w"[3�gj���+n��u�<�^F�T�/pѩf��[T�ҷ)�P��ٱ�c��g�&s.B������i�5y�j"֋��3N�[Y�%�X�Mo`V��
�\Aʁ�Vۚ�6�ͤ�5to�w��k6[�[x���m��2d2nmŘZ�C,Fwh91���9�Xړ�N���C �N�nQf��iXyHB�]�]��m9�@ �X���@�b6�e��74iF�p�{b켒i�*9`��1݋p���ě��^�cf��[uےQ�{�XF��{�к��`���J%JE5��i�6�
��{�w�.Hv��������30��zڬ+�Sz�Y�ׅ3����׮S'1�U���W� ǳB�Y�'5V���^���R��LcFH�Y.��#�%Z[udj���;ġ",��4�5��f�71KjnY��$�9YEUy*M��-,M-R�Tq�LYY���h���q�D��vN�K.9��\�p8C �1�Y ��ˢ�]d�Z���^�Fؔ$��(n�M:X�D��(��BJяwp\Ձ�Ưrn6�R�sJ�6޸5V�;-̴\�ddV-\TNFic��ݻ�GSi�*&)����p��S:���bM^C���q���,��U�#���8Q�oP����Ka�F[��swZ��]�2�y�Y���;d�6؃F��MZ���u�T����nV�����6#F(UU%�j�n��$�JG/6�a;�Q�oORbPN������@�H���Z,5���u�.Y�T:I������"��Sc��"2�1�k��酊�2\nT(-�j��ؒ���b��㗍�@����a����0��Ft^� �Kn
�����+km�3`��S��!��oU�����Y�-3���pq�T����8���SRkA����5V�8�c[�	��WkE�P����
���i��l(���TR�h2!��)�
H��ޠM�P]8�E�F� ��A�nc�`T�Ek�l(-Fs�[vFsu�9LVh^
E*�]��.�qD�1����zn�#y=��bb��=�B�[žV�Y��ѯN��"��V
�x�B�mcOض�D�����!n�}�7����+7��Q�!�e�WƳ��Y=*r�8�K�i�p�0��t+E�]v���B�%ܤV�[��b�9,h�]\vKw�GB�xR%�M$ٻ�`��iV�H?��.��o(���8�R�^΢�[�_Ce�f��3�d=՚�["�FVe�x�B�l�D�4�Ɓζ��}��lI�G��]\��t��4Z���T
eî]��l�i/�)������!��7�U���Uvԋ�]tW�¦NCk�����
7LM���E�m;Q Hs4�b�k!S�gAzʹ�d�lBEh�Q��.��Ȭ��	R�x��<V��8���0�4�4��.�+n�k>`��b�ʦ]j��$�%����(�2�5إ�H��[˭�탭B:��}aV�c���WpE��%�5�U�SJvX�)wV�֞�h���u)�m��^���L�Ԏ JH"⩳�]�����%t��+m!�Ė��j�!m�Pڵ!G&�:���V�Z����,L��m����YH(Q.��s��(v�淌�s�k������	,��zcjQ�dȭ�i�d�2�H�8	���������=�`�0���N%�;���Xk��{Dì�n�fp�Z6����+9ǰ�y��9�j�Y!oqw�[hdɋ*.��B�.��g&x�Z�m[�b�Q507�h���8�6�Dis[⦲-Ri&�I�j�,M�3�bQ!��ikKW2Ql��8�Ѝ�ej�.��hi3�n�Z�y��nj�c�I�T��J�9�ݭ���#�u��A�\B��ڈ�8���v�*�Q�X)mXɗԆ��V�-(���MM%h9��ynɜ�a�x�$��=���|��٠I�Jri
"��}�1u�H�[K�%�zqS�q$L&��h(�Ej��^r%%��6�y!9S06��*�m%!	I%�e���t�,�Q5�&뱇0	�W%�&�@�D���V�
��|z"ܜra�a/��ι�Q�:Y���&%�a�5Q o�� ϴ��՘R=��b��|M�I6Z>�V2�5ؕ.ډ+N�ibM!a�ٙW�Ŵ�b7S�\(�z�յ�		��1=��jiH�:	�h�{^�\G�D�M%iEK����ze�ĭ ��p�h�U��޹ �br��iA9ɲ�e8�h"i!b��z%��K/IF�R�enٳ�dR�ڰB$�԰ߢ�UIcG�ڏ)�A��J�J���r'ɳK�8��/wzb6�:�ʨ{�@dܷ�*˷��R�@�K92��0�A�6�&�;hY�=�d���U�N�٨���z����	/E�5��X8h"�D$n���1jX�'HB3o"R�R�qr��Փ\S.$;8����dX�KZ�\b��Q6�M!�X�Զ�f�RMQ��=���+1�3-�Ψ)H��48��8A�m���]�Hkn�x�1c[�D1�����KjVd�є�L9�@Ak��*g�U�b�F�4�F��Y���L�*2�hQd�
*И���#z2�f�҉�mu(ѵ��]2����u�K�冰\:�p�7G6�M;	��s�}u�l����Җ�$I��R�J�i��,�W�� A:��V�T���TN �ܖ��Nn$ڬ�Lf>}��!�W{�ݏD�S�E��+�Y��8�YN^��� �8��ىb}dq&��+�=+�w�.�qc&��;�M2��,�6M]��q�����0·�� ���B��o��Mߋ�?Af��qW_o��(��_y��z��F��w�h�6��ݎ�\��ݵ\s��\�	�R|�xn��A�07|���&�x#z/��7�0��P@h�켉t4�x���(t�ǤR�b�y����W�����7rN���lv�.�+P�,y23%�"۸����s�p�<�C#^�$�n<��Ҳ�P�v�����N����P�2q���v�']8��ő쮝:�B+f��Ջ.��i�PЭ�nP���r��QrVfYGyg�L[�R��֬���28���^��c��/l+r��HZ�������%��.�T��F�+b�glN������z�j�uΔk/��g;��}��kw�7�s>��sE^� ,��]��:}�v$�x����eahƮ�Gs��ґr���qw�x�2n���N��i�`�z�}Q�t��!:a���Zښ���QK�G�%���o�j�p�vp&zZS㗉�u��ל{/0'QT�*F����j��i�Mf�ֱ�"��uVk鏋}�+8fQ���7��0Dؚm.±>��f��ţk�M�K�����c�6/*���=Wm9ZLy�O�O��ׁ��ǖ�{M��<P��`B����H�3^���R�wf��93�d})���ز����/����n^%�L�t��2̀=M4'iwS���w�p�ze�}OMs����N��c�
k�NA�ǹ���(�SJ#�)Bܚ���S�|+'W`α��Y'o<}�),�}����I��IR�šv���>!]sцu��t�K7���!�I��A���f�:�S�n���]\�pLU���%6�U�����u ̙�&�T}p��WJ�{�ʚ-XM�)�P�ês���I�{Ce�`��h��ʡY-���t{�4���Rk:[UYL�,=n�׆�j�o\�JVq�q;���&N���=FL��������K�^��9L�R���z�:7�8�EX�-�o:wc��i��t��.���Gd{n62�<w�/rH�l֚b;��5.�#���V��˒��i���7�D�VT��Iu�,l��Tv'R��3�z9J5����|�xu^;X���A�pbTEY�<����i�ѻ��I�kgHg�1��L]i9R��B�P*vn�;���Ƴr�I�
���L�ڲ�����O���h�Y �Ҍ��+�$���u5m�Y}:����l�����4��Պݖ����r�8��sېj-i�y;b��z��g@;
����+z5\�Ҭd�wm�A-���8���/�r�LaSʾb93�w}r�B�V7��
­�Ky�(P���ՓZy�ts�!b��Ǝ[ivV9y���>�G�t@�j�hɪ�V�~��ٷܠUF��p���a��4֤�\�¢ӉI�n�.Uʲ+�a�&$Zү.�]�z�{��݈7Dv-��6Y]c4�X�ƚ=CDs\9����g&3s*٣ר!�X�t[�ɩ)���f*u�E����>V���3w{Ҥ;κ�8�;ϖfwWD)6��52n����i޵��]F��^�^{��]�Ti<�@�'l��zf�A����-�4Cv��0�I��O �3m��Q��f�tU�R�Z��;�o�{�Η>�{Ң�ݼ�)�w�A+0��������$+�N縔����T�׿>�m��'��hlg�tY[�{{������V����ux��Q2xFt'���{�Jv����3[�-r��-�V�ô�<};��M��&)����r��Lj��2�	^f���2�0>��
h,�뺭8,lh��9�1�4�Q}]��e�񨲏9�v<"�'�/(2+)��"��4�.�<櫁��B�Z�����W�5˾�v��W�q���P���j����++��v��"pb�J�� �q�EtS�ջ����㶕n��\Q����x��lI�1�K��[�Cx�Eӑi�Tk�����C/d@�D̊�	��LZ��N��Ю���fX�eh��;v�2-�s�k�>A�Y�ٶ�sQ-�n��ٗm�ɸ��ˢ7he@�!i���l`Ś^R��첝�_6¦f�k�æ��̮{�$���'^�}�|�x��C(�ܾ��6nNo6-
�xu�\70�7dڼ�[�/^�ݸ�=�u����h�vz�QY��)��Z�y7�o3υڝ���\t\۫��z`�sY#UJ��9C.�rsw�U�`���T��T5��_d���H�H5��H��z2�sL�\6r�Xm�pu7c!�a���͕��+�i�;tV�ӅL�I�[Wz�d���2[�eaJ��p���p/�7�p��8�ǇN���Ι���柱�[ݹu;��0���}�a�X9��ѫ�ǖ�\غv�6����jc8����xG��)[�g
t�ʷ�@ƺd�¥D����{���2�P����i�s; ,���Ŷ")3ƻwl��>ysC;�ɢ����U�H
A$	֫hW.�����t��1�ev�6k�����9��9v�Ngz�؉Y�M��f����je厾s
�ꅠc�؎V���F�x���s�S&�56�4��zQ�M����G��Hq��yta���np�|����إx�g�YZ�ҩ��px慏_M�8"�Ec���up�3\(+z��5�)d=oze�Vs�t$m/p�/�����W��V�b���9h�C��Oj-��t8n�m�_9Š��M����.��g#Y;��y�{盫*�Gn#���*Z&R\��.�B�v��»9^U�	��Ȑѣ��A��O^c\��Z]c;�;�񵘔Ҹ�9}�gW;v .zjb�k3r��\����U���$����\��&r
뫵�}�������7Jk9@k�a�弄���^���Y��I���������O��ѽt8lG���/����e�z�ѫ���J59s����kN�����9���:�����\�V�y}tVú:z�|�J�$B]V⾱ku6�M�d���I��SrC�Y��.�s���އ�l+����2�X�7��`�=��U܏�v6��ܥ|��2�������F�ǹƙ͋�o6�R�".���Ӂ��e�}��ـ�L��cjE�Z�ә�t드u�+��{aՅ*p5vt������Zw؏[h��o�З�2��Q+=����j�Q>v2�Y}�^�d�8�5]��c��B�]�qoP�y%�x��5 \NK�֓'�,��T��ȫe�`O[�9�;��+�I�j���\AR���;�N,�8��gb���b�|
yqڸk�y��c�F^�u5T�!y]�^������Ac�0�S^�>�n�uf�b�Wڞg^�+��뜫��i��WV�u�G #���<���m�ρ�Q�β�5�fcx��b:�s8w`Ǖ�K�u;6�Pq�y�W
}!��[�[O.i����m�a�' a±`�LLZ.�랉g�.,�R�m������{]4�j/]S���X�5�,Ays�)��Y����������^��
Z귔��8�3&�č�N���Q&e.C���1�K	�
v]&������9q.��F�<z���O*K�%%���rl۽|��=;��Nv8�p5d���d�O`#n`.P�0�Su�u�7��bl�"Ы�����^O^�k잱*�@�q����uO�@�j��ЭC��%�wx�J��������ժ�e��o]�V��d��4>�y��i|M/m���R����:��N޾�:;��0Q]Q���P���,�<8�ĜwY��k���*c����5��A�yac�+������TF���Hx�5V��DN�K:��m��hә�R��Ifr������m���,}6��)*��ѻ)'�۩�͆��&��o���m�v���\�Wpy���v�d��NU���(Qxy�ޒFWY�lo:D����kn�Ki�2�n����t�b����d�(�G�v۶�^��%�o4�ʄl��]��lǾ5ثp;>ի�s���y]�9�I�}6�]��������_473@�Ǘ,�%l�LM��nnǅv���7��� �W\B�pe��r�o4�>+�ʽ�wH*Bce��w+��%��-8X�{ri3���<1to�Gg��c�|���TƪL��{��S�U�r�����u�KF�)�ǦM��a}*�u�+S/A7�����É�du�5IIUT�R+������g5Jhϓ�C,�!�j��-�	PqK#�%p&t��ҰdF����j�T`���c=�z�L;�oVF4umi�9®b�rGτxvƲiӝ�ǳp���hթ.�SQ77�c���*嚕����-h��EoX��b���������n�IW-�{H����Y�Ůp�<�Yc�8��/0�#�DJΟCL��5r�q	'0��E vp�k+�;���dU��w��O긄NÆ^�z��y:��UX���=�͹;�&�˾�/�iI���I^��4/�ͪ�~��\o�U�КnU!e���\��C�)�T��׀����BȻʒ�;-���h�PCH��l�Ƶj�Y��)���,3՘ �02(0q�L��#�Ԑ����C���y�W�Ge���^��1���1V}|�|"�� �5	�9��3�V]�k��gQ�e)�D�:��[�š!ؙ�����ʃ�?]��=���fn�c�9kwN�(ʴ��_T^]����o��Nm�w*�Ǽ��V��.Vg�eoE|�f+��W�L��6dX���Y��w��)�ݨ�w:貮�z�CK7T1���Љ�:@�����}�Q�l.X��G�i����P��U҉�z���d�����H{g
(��Ƕ2���w���o-��5�򹃥�#[�f����՜ !�Z{E�ݮ �(�Lo�ii�3n�TR�����6w������Jyw��B1��Ͱ��9���4E�A�f��l�ʺ[���Dq�5Oj�p{s,�a�8_)3q"����&=��{;�L��o3	�vw��H���N�N���I$�I$�I$�I$�I&��]��v��w�p�,�B�'���/�m��^WS��ux2�8�{v_iu��S��m6Ѷy}W����-�.X//����˾ލ��"K1�V����J�EE�b�"H`�D6�7�����]� ��VJ��E�Y�0$��R�W&4�X�4	�I�KP2R1�rb�a훩�b��,���H��I$Ą�2����e���Ym��׉�M�J��!"TFYu�����xXC�0����NDZP��dF���7��pU��g�Y&d�h����8�A�ט(6��������LpUF�;W��BђB�$� (�p �*�"��n�5%���	�N�*�
oJP1��ق2H�pH�J�Â'Â��Y�(�t�TXK�d$���$�J�SQ�ߙ�8���*]�q09d�4!VB^a~1��$��(�@�bQJ�A<���g�QFЊyy(`*A�yEF�0ba����/Ȕ�Ͷ�#H��[u�̩�,"�� d)P4�f�yfvj��#]��°�9���R	����8n�aC�- �P^!6u�t3&Є��� �DD�8�qI���c���I�0N1�P���L�`��!�5K����0���B��T�E�J+9pж�th�n��F]����rk(٢IH���TD�ADI~qA1��S^�c8��ݬ)��'
KL��$�J�SQ�ߙ�8��DE/2�K˹2�=5��`h��Ң4)�G��DBP(��C�A����Ifq�͝hZ1ȐD�(8�p �*�@�Y!?�������3�P��)4��%&m��-y��mĠ'ћjB�y:ʒ�J�a��	7i@A^dB́	2��+F8X�J�S�!�ve���?�-���|Sf�}%�*�~=�M�o`H��I$Ą)E�I�8]��Xl2�HA`���D�%#�8(�FjU��w9�����0 �E�m;ۆ�+dܴI�!�����o����L:��O2���Kmᅄh &�ԘQ6�0ÞprU
C���E*C��lQPF�NU�R�E�J �%�����q��E�䠊���i���u���I8S���J���I�m�l�q�F�Q�f{��53۰�B%H����AI$|��|E�R8!m#$2���Z2�y�V;Q����>l4b�lRb��}��j	�+	 �@��ȿ"S��6ۈ���f-}�髣��K�yy(`*H���GuW�l��8ĳ	z-�&�$��0��L \!���_'y�u�Z*�
~���w��U���	��{�'��p��S��������������o�?ο�;���.ad��gV�Z�#���	b<镼�Ò��2�$���â�7/w�T�*�U�L`?-R\~���F�r�ѻ[�4��3耱��Z��<lR�R��5�[����K��k��]�-�w���ݗ"u���'��=N�v\�֝5���������3TgL���[���2�C�����`�D�0�7q��۶�1'Ȏsw�l$�O������8���%�ÝqK)s7pp��=�
���OAlS��K�|�v.ż4���rgG9��v�7a�2�CW�-�4�5�8{-`�{ز釆D�H�
n��ٸ�:Bж���NJ��JW|d��7;x�ǉӹ��&�q��Y�K�����pVZu���BY�o��j⎛P�u꼜+~7'his`�M��7��]}k$D�� }}��}l�[���k_j�k��V���U��y�������Y��zxضN����6�u�����Y;��9��u8��ƅh�bͭ6�W���+D�m5�1m�v()��5�gr�w!(�}������=��||kZ׶�Ƶ�kZ�ֵ�Zֵ�צ���Zֵ���k_�kZ�kZצ��5�kZ׶�kZֵ�|kֵ�kZ֍kZֵ�kƵ�xֵ�k�ZƵ�kZ�Ƶ�kZ��Z׍ֵ�kZ��5�kZצ��ֵ�Zֵ�MkZ�kZצ��kZֵ��kֵ�k_�5�kZ־4kZֵ�{k\kZֵ��5�xֵ�k^�ּkZֵֺ�~5�q�kZֽ�kZ�5�hֵ�kZֵ�kZֵ�|hֵ�kZִkZֵ�kZ5�kZ��]�\:�w{�;�o�V��sH����:�.:�l6G>�����-�*uȆ�B��7����i*�������g����;�5��i>۶,0z輙[4�r�v堙tVn�s�N�M�QƜˍ�+z�f��^MA�"*fޭ=}���F;�6��>'#8���;�����8����\ޮU�ãL�6,�n0�S�T�ߕ���F�`���+�(�ij��]0�Mj�%քӽ�u6+Y��A9f��9R���˽�WZ�oKZ��D�v�nozb�ܭ�������[)e:���OH�V,�����0�a�
�ui�m)��7����uk�[��Y�+B�F˺���®I0[�廭Y�9��Φ�N�t:ʣ��e�p�Μ�nE\彤f�G
�R�6�]�����\w�4�,�p�ЭB�@P|b<3��:&p�3������8ϑ�G�@�iގ����7���u��b�I��sm�.�f�� 8��]w�����jB���%�*�-��V�P�� ��X����|�r�����Oo�kZ�ƍkZֵ�|kֵ�k^��ֵ�k�Z׍kZֵ�k�ֵ���k�cZֵ�k�F��kZֵ�Zֵ�k�Z�Zֵ�Ƶ�u�kZ�Zֵ�ֵƵ�kZ�ֵƵ�kZ�ѭkZֵ�|kֵ�|zkZ�kZ��Zֵֺ�u�kZ�kZ׍kZֽ5�kƵ�k^��5�kZ־4kZֵ�{k\kZֵ�k�Xֵ�k^�ƼkZֵֺ�~5�k^8�Zֵ�xֵ�k�Zֵֵ�k�k^5�kZ�ֵƵ�kZ�ֵƵ�Ns��t����j�pϞ'
��wu]\J:_H�ɖ2�`)���pw����M��Us�c����w���>��w�֚p=O<9�Z{Z�c���^c;eK���Lr�n�ѷ#���Zec��y���N���l�;o�C����vj>���rr��I��L����q�9�����J�+�
�����Gp�%Ez��D����0��IbX��i%�%��n@�ڹ���h��a��+ef����^��*��K���0�q�����bz"ȩ��$��2bGq��R0*ȏ4#�ki�Wf�|���J�{6ve�
;�7���t�mY��yw�;��Qv�Sh��+�-�/mT!X�y�Ha���3G'�Nh��2-U�H�q��-�}U��IQZ�5kjG�Gx:�#��s�{&bVJ�r��N����%�O�E����ʷ8_	��a�����r_�ph��uQ��t�FcWY�r�a[��;,kk"U�LaPǣ��(�@@�gD�nƥ#����(�Zy�fu\���.��z:�pe�h|MY3��p�h�$�]��qJ�B�]��;�ny���O�_��׍kZֽ5�q�kZֽ�kZֵ�kZ5�kZֵ�kZֵ�k�Xֵ�k^�ּkZ׍kZֽ?ֵ�Zֵ�Ƶ�5�kZ׶�kZֵ�mk�kZֿֵֵ�k_�kZ�ZּkZֵ�k�kZֵ�Zֵ�k_Ƶ�kZ׶�ƽ5�xֽ5�xֵ�k�k]kZֵ�ֵ���kƵ�k^�ֵָ�k^�5�kZֵ�ֵ�kZ��5�kZ�kZ�Zָ׷]xֿֵ�~5�k�kZֵ�kƵ�kZ�ֵ�Zֵֵ�k�kZ�_��l��dL��ͼ�U���lZf���pfi���[���ei�P j�g퇢˕5�zݻ����AC˦[��[d��ec�C�ot����6���_YNrM��:&�����}7�j�ᢖtb���Y�(��N�wk�A��8%`��MT�ѹD�a	n��6�Y|d^	�����`|%Jf�ZN"lM�~����&���^��T�vUG׆C�%ȫrX�5�L���]WN뻞Δ�`�,i�ҭ�ա8�ۓ�Q`�%W�w;}U�G��Υy�i�Vw\�"�K`�3���Xf��ϝh�YEV-��e�m��h�|졦P��{y��q��{�K%.����wh�--^�S�ǋz�T�Q��:���]iM�#y2��g>6�2�;�\�T�Ѓ��.��zY�P�|3��$��X��Cz*.g�:�@�t9A�J��թsTn����1wa�y�38>cX$��Uw�Y�Л\j3uG^C�@<=[��4eNͷ��'*�\塽�;c�\��YJ�;7f4Gvg1��Z��DҮ@e;�(���fWk�s�:�����U���=��|{|k_�kZ�Zֵֵ�k�k�kZֵ�k�kZֵ�cZֵ�k�F��kZ־5�kZֿֵֵ�kZ�ֵ�Zֵֵ�k�cZּkZ�ƏMkZֵ��cZֵ�k�Z�Zֵ�zkZ�kZ�Zֵ�ֵƵ�kZ�ֱ�kZֵ�Zֵ�k_Ƶ�kZ־5�kZ�ֽ��5�k_�kZ�Zֵֵ�k�kZ�Zֵ�ֵƵ�kZ�ѭkZֵ�q�k^<x��q�kZֵ��cZֵ�k_Ƶ�kZ־5�kZֵ�mk�kZ־|<���^d��ϓ�8������6���b�o9H�#o��y;��>��k��+M��,�����Z��f���ak��(�fH���{��7�I�@�t{�so6��]6�$��8�h�;�Ve�l��mB+�rb!�H*��y���'J6�Ud�R�qB��@�	��e�P8U�C�{hn�6�^��OF�[(%mN�1A���66���L\����C�BU�fġ��cw��݅�仭��L<�_vS�i��=ŷE�9���x�1����9Y#��|��:�As7s�r�vBT���Lz���T����#r�G�O�g�y��J^1��k.�`�����.��6�W<�����lQ�S���n�ߩ�/頰΍c�2�������Y�'����]�`lv$%]�=�]hKkT�����vǛ3H��9����-���U��>�$d��{��,�.�;���6�[a���o]�l�.!��;���F�����y�2식�. o�����zbN{�5�C�����b��h�uc����dYM�#5�ɺ*�Y֧K�Aq����cUp�1��h��~l���}���݂�b�I� %�*����3|�=��xAi}�%��8N#Y�*��y��ݷ�x�X� ��.��R�B<+�L;�{��U��:h2����e�w&���[���N�(�v�&	��q����g�{3ě�	A�=�:�\\�`��]Z�Gy�g:�h١��}�
��YĂR�Ҩ����8a�l��
ËbF�Y��1�'n�"K�C�ú�4�7��Ąq����/Q����\�>r$GUό�����=ց�[��Lq��W���qswR�P�{:��0��Sp�/��� �,�cUvv�v+e�q=x �m
�-��b�r!=��_we�(r�b�R�ӶB��BZ�ܺs^����oV,��_���^��V�W9؞,aǴ��p�й��S���*����r0%`S/���^�=��w"�TJ�������8*�Ӛ3(Ů�^j���Qh�G�PG�ddK'ez�Ɉ�Tl�R����U㶹$�g���uT��2;��d�֤!+;�kC��/��X`��ЪP�KF؉��{N��>w��e�Q6Ҟ/��)֓Jp��˸i�M��Aة���<��Yt��e��fΡ�/�d$(2)	� {�ؕ�Ո�:�a��]��7�p�T�P�G��J[�d>�eYΊ��mٳS"B �v8�YѲQY$Ԍ#���ͬȬ_"m����*T���x%迆0A��Ц�(��ae&aǦ�y]v�!آ[����V�Z�q���%��hx>6i�D��\�`��X5���(ZF�%�K�/�V�rv��|J��D��a�2���2����u8���x�M�j��[�|N�O��uk���3�t^f�s���E����ƶ�ַVO`�ٱ�e,��L��%dB[�V��X=�2�F��Xwh���H���#n���o(�)�P���"!Ct{�
��Ֆ�W8pJ�d���6z@���qZ�eݗ�/��v^�ke��N���A�V�x�^z�w�\yDL���x��E���b��v�Z�Q̠�$�K9r���G� �Ѧٕ�[#�����bt�����*/�� R�|���*a>��ufYvVM�e�/�����]W`�j�1�e� ����xx\����V�칧*�G�Ρ�V�7w6���n��*��D�R\U���+S�V3GU�;w��Q��a׭�r�#��v{����F�.��N�����ܣ�}O�+}�>�j%r�₸MY�ѱ_f�y�g�=��_0��h�[�Z�vU�'Gj����)hX�ﶱ{®�::�V�n��݂L�t+m��뀼�YIK.� 3����F��N ޸a��0����>PX���f�Cy,���t�;�w��6Z��w�vپ&��ޯ ɛԁ�^p-���Y�Y����Dc.�q}+��i�q��4��YF�2b�oM��ɸz}9�g2�� ����WT��z�֌Cc��e���������6if��-�C�E����v�#�NQ&w�V�Pλ�ޱ�P�]�ե0\�e���r^�"���M�ZrK�#�θ��5��2� $�����||�]W᷻f��/���3�nE���9�t�.Sg��Li��W��#�:�S�g��$`�3�
�����(ќ6�E��Q���R�lm-z4���%�R��ֵ:�����G��{��ݢ��FjmM���)�߽�255]펏�v�y��j�qr�:��T�t�Y�q�����=G0�}�_U��H�/&.M�?	M�V��E�e��ʉ�i!v��A�f��?bTq��m���Z���9oh�l[w�KR���.����Fdd�4��\�W_d�	�n�vA.̫���:��ٙr��=ϯ���d�Y/QN��#|���x��J��Tٛ7��|���&�鱃���R�Nۛ�����'ў�&�aTɑ�����.�b���L�.�3K*�0vAǪɔ'�hֆ���u_�t��c��P�i=Ċ��b_D<��c.�I�j����}�����{�1�8�eL��:���\��|#<�k���ӣ��z�`��f;����a��n�
]1�A�
�G'ۧ���e�1P�&�b�0p..M�N�̫nv��W-��7T�wSչP+�;[]��)�1O�J���΅zgD���s��H{�j\C:Lh��q�M/`�t�Ղα&�i��o��пN-�s3]c������z�>[w�*-���<W!3�<w��u-M��CJ���l辗�r�ۭ�5�p��fZ�ILٗ����N!�t`��N��l�v]��ʌH�Z
�p�,f��z�H߬�˸�r���lu�t]�+�$1)�w��[ͬ��!,u��q���H_V���!�*�n�G�/V^���%ou
���'�r����[�r(v������0�G_�p]W��5�(������lכYFN͏�9���G�2UɊ��[uL�;�T/S��u�]O\郘�fa�X��i9n�%Z��{��K���a`��x�:a�z�C�RP{JG�(Nl�����i�t��O!O�k���h��,�:'�UÛ��2��u�B0��Uuؙ��3W=ѕ5�_�냸���ַ��\)�����i_(�� %��j��s�P�Ν�'�Ж,ѹ[�W�]�aNQZ��K4��LV�\n�[2�L0���+;{b�A�˞�ޗ����OH3�WD{�<���=����ȕ��b�2��dtP	+ou#�x��Y��^���Y�^�ͬ��]��L�v��N[-�f%.R�T���kkn�yzb�x��ʸ���c]���9��`y:�͝sE����˕�/9"��o�Y�݇5�s���s�.��a֩;�hf��S���]%����5˱��"���N���8�Ix��ùN�ϝu�����4~tO?o�?p" ��d�����G�_��Ͻ�<���C��O��~�J%SM*_ě���52[�h�A!n^P0D*x��EB������تIB'�18\l�-��:b�A2Ct�����*�a3D@D�F�� A^I8h��%��l�R��Je4*�a_����"��+��ysY\М���NWd�VeF6u��:��:eϒy{W,�+Y�ݷy���!�{�֗�ʹVM���5{��M�Ƅ8�f�w���s�^���G�hx|��|E��'��9	ՆV�Nup�o*v��|�H�V�Zv��q�æ�$*m����7�c�琞��;ВƇ�+:rÒR�5-aH�k��1��e�so���w_���[��\��������}sDӆm�9���{*vhÅ
������X�,��9��\��1Wg�����'2\Z���J��:�|��c�ި|;0)J�o^e��+������������#��rhX��b��ge&�k�l�ӹbY8.ըEj{��ݭ�� ��СӺ��ё��j��o��r��kޭa�j�*��u$�����l3Q��&Z��n¥媱�L^˩zg=�!nMunCCE�N�nEfv�Ě���f�f(e��dP�N�ˎ��*t*^8f�־���]͋n��u���]��#R
;(Td�%$h2�I��"zŒͯ$��*� �;d��EB���HO,(ʦ|��D�W��*���e �0��,�

8�!����D*�L�i$�l*�1�x�R�$TE!PS�bpg�*�^$�W�ɷv�7�X0�
03lj�D������IF/+2�(RP�>uG��4(�C�8�0��E'm9 0��6�vj@�m�PIAȂd��(�m�%��&�F���'�E��g&�^���;4�y��.�&a�dÓ Noq�Ƕ��kF��kZ־5�kZ�]u�Z�ܐ��Dsd9��nB2fdEę3 W�q�Zֵ��ֵ�kZ��5�k]u�]k�c�z`�m�� ����շ�o�������M��N�ګ�oMzkZ�ѭkZֵ��cZֶ�������>|�ɑ6mPI�rw�O�w�g1TNn�K��Eʜ��rq��q�Z�ֵ�Zֵ�k_Ƶ�k���~w�!0̓2
�d������v��r4�y�q.���fcgv-�NsG6D�%��;��d�B�!$�ȉɱ!gYx���d�_e$w_���:���,�^&Yą�J�[ń��Nvw�L�fIr�fL�|\�B�$��̨�܂e�9�q,�N�m&ud$�Ki&泓ifY&I-$̱�'�ՖR�m�RI}:�wgy�-�F"���-��
�ux���6i?Y$���%�wbNR&Yi6id��p���I�����N!��܄������"��'|޶g%]볓�{O;�v[��ҹ�9�Ni���9�\�l�=iu��br5��NirsI����I8��	�X��ߛ�cŒ�/����RN���
�<�d�M���������`��>��K�&�A�E�D?��_�k���;Lu���]��EIx��eG;���2Vt᣹mm	����ϯ�f�{�Yɹ�F�#��F�2�Jg�d�!��FE4]�DoN����睇}I;R*ǈ ���`�(���u[����bD�m��"BIGg��`pX߻/.9��xf<폎To��{ܫs��\�
���"No.��	68��Lt��j�^+KX:��(K��_͢i�ئ�z��k�	W��kf�Ś��W{���e0����G�ZEJY�@���p�P�j�ٍ�5�|B���m��]9��T���q��S�mT �|�	��PM�����N������{t�d�3	� �EXr_		e�sd�v��Ȱ7����L�����t��}���wQw$[ϔ^�:��R�E(�i�Xf�A-�Tb���^��:
�P�~S�C���@f��o�0oP7s���}�R��;F!́}�ϵ���?y�����'W�x �0]B��I��5#�k�69�]�N�����[�F���ʗ�)�u����s.`�g����܍���#4�}jƙl�Z�4�e�,��\Z/�]�����X��2l����zt�x>����j�2�	,�MN�&��Y;\��y�>�����c ��}�}��<�}�[k@ע`#W�\
�4�x\���}�{�l3	h��EV��[�O�����>3�X}9�!O�n<�hЋJ���j7
,�ԷD q�U{0lf���h˖�6x��qkϨ��RI�Q~���^?Q>��п����{.)�6�~�>n%���A�C݀��m8�v�T�43B�`s͓�N��8\:�;:7�g,����MC=v9P�T��i�����y�Q^Ql�zy��N����
İ���(il�+�VӗH Ί��%^][�ўt�
�ʓ�j�Ҭ�gI�*@��{,�i� Ӛ���b��$H>\�E]Z������]���J�5#[뇲��Kq�Y�ȟJ͜�psU��K��oK���t�E6���G���mTZ"2�e��r�MӪ(�}��t��)vaXq��k��p��)��z�:���)~*���߇��<�=�G;�������1���e��ԭm�E�)�����w:�R�_fv�;��m��e�=������� \rfoX����~�E���Yf�è�cn�b��s=�4&���aj�ޣ�v��X�5��-�I��K#���{BGY�N�R�Ɋ8�6R�Q�I�|"+o��"�]����HŜ�>�u�(;(�9im���+n��FS8���G���f�sf��X�h��n����85�m5q�^3�zR���hs�G�O~h{�Z׳4�L)OvZX�	�F]²qn�DjX֭��m�����9�@�z�vCP=<d����#B���[��{�
}������U��������m=�@��D[sw<�4����7��k>x��T�k�R��'#<XѬܡ8.wN��nq�`�����>��j�EDL������X��}�	oxkUf�*&l*Jef�ǩ�Ɓ�������[��Im�*�LZ�G���h�;�I-�[ll��w����FmdV����%*�z�X58�bhL�Eu|(}�n���Lo�@>^��qY�0_`�\!�)l{�3��G����g~����&���~�v��������`�3u���s����'{�ݟW�ģ�y��}�����^�b�{��;���F��X��&��[�v���u��������Ʊ���}p;��߶f��� ���p]�t�7�Z(Nz���3N�S$e>Y�ȁ
�*Ro��sM�����i��'R����^H��l�*=�zMo�"�
���Eze�^�k����}�!�^u�G%���[�㷟x�#{�Y�N����$�L�q���3"�N�˞N�c�����b�YA�4��6	z����30�^f	�����. xy���,L��Y�����p�u�<~`���O��Kt�Dk�օJ��%K�t� ?ݺ��v��(��-�=�N�V��K��Έ���<�*u	J�9>g�G:}�;������Y�Ckl�?N��^,���T�N+��W��
>r��Eg%2��{{]��0��D+�F�[�h9WvCV-�=f"m(�u:�wf�H��6��P��İ�/qt��»��̮Y�;��k\�.�S�Q6�L2��"ۊ����:�p�B&V���Ȩ��P(���̟�cČC�>ds������������(�D�ߝxװ3Gȩ1YB�	F��m�H�W��m�w�z6��Q�*����� ��/`D0^f�y�hXa0֌P2aF�\���7wyrق}�/�qk~ !\A��q�}b�wE!n䊼�d�5������Ke���]��+�ַ.��;X���E��W�U�����&���SU���dߦ�؜�}����S"�=��%{�g2�0Ro�O�z�-d�^���X�\�>Ι�?%�� 1�AdOϣ�ܧɄ;�}-�����>�0L��F��-�E=�m�O��WW��y���������*�ߺ��~Mh�=�}�ȵ�n�oc�U��ZX����v�����)h���>w��u�����G�.�f+6���ĕ�3䖙���d��is�l���ٿW���}_KD�y^ՃQ�.�����c�.7���(��f�W�\9�s̬��n�`+��IR5��^;��'�V�ff�WS������f^�3{�Z�@tm᣷+�&hs��\ck+���/�޺˛�M�w�������<����0`�ř$nA�	���a�cfy��CL��OR�V-(6�N��l/9(�ň
��%�!\��&u���I���V��C(�%�M.@���2�t�j��G�׍�y	�u4�*�Qױ{i gCU����/�ˇ��;�kJ��K0��L�I�쑈o����1
#�}��dU-���5�`�!� �U���`eA,�����Tl8���8��E;<N�	��qR��)ʼKh�i��M��Yo��#��/�f�B���,>�[@3�'��޻-;�MU%�����|��A|�+����Aв�r�F\DD�nf��	m��Є�|�3�Y.��pU��q�L���.��S��a�z�AU�U]�>M@4yc�^�������$"=4?v�l���fI�c,Eu��1�AA�	�\��Jo4�v.�"�:�E]!���}0c�������"�t{��;OP���3�y��[�4�gu��������r�Wp�yǤe|������]���fP��b�-��M�:i���R0 �hC�;Oi��֗�E���YCwRկAT��k�B5K�ll*���|�=<���b���|��Z!N��jJ7�#�o���JT2g��$��{���:�`�X;�Α�7i��r���/o�H�t�[eJD��0G>޷�8.��VAR�/�ؓi��!R�L��@/?�Dw��G��Z
�L��핆���,O���Y,���kgT��P[�fbv��y�2`�obܵ{���Ԛó�Y1rcϔ�:�cr��-�Ҧ�=Xgn���ژ��c�%�q���؇ܲ��<C�R3�O�=W�H~/{���ɣ��4��j��v��ۧ��o�Hm��^�C*ɤ��d���S���j�W�D䆺�͓�L�ȯX��l�.9�H�� ��fJ�J��/'�N���q�ꥂ�8~��u:�\ē�0�=����0�bur�����v����^��1�˸��:#���m^�콭�)ոܵ1���5;�ېIo�P�y�gP�̓1<`F`F*>u�o^yp��>��t�p+a��_�,B
}>1���_���C:��|p7���wk��K=R��h�r�����Fŭ�������	�c�wXM�阀�[lq{�춪�/�©�_tq�'����o��"���N�UO�x��I��M��<y�S �BT=T�x�%�E]ZS�s�I���W��&b�5{xc��{�r,J^Ȋv�f[X����rb�*�g����J���u�ݭ�}dS����o���1�i��sL�^���Y=���=nZ�:�Y�2S�ɗs�q;�iY[�iI4%�?���7�j�b��h�l���u,"e����Q�͊�uo閨z�i��5F���G����(׽¸T��a\WInbÍ�(1��Y>;{,1�P�J��������/����}�vN0
�y1P+e�tVY�Y5b�ЊѐӚ�;�O��ynİ�ܵ��q�R��h��|�d~7Z�=�4L}qˆ
��F��x�n��	�f���K����|�}���NI���]��Je��mk��.��ɤ���V�2�����2��B�B��2�5nR,�M��K�I�c1�g[>w���w������fCih�gV!�k}H�5'䐙�L�ƻ@�oD"��O�eu���@�39�M���)*/L�,�KQ$�ٟ\mS=u����{�6��'?t�U�������lc��cףzY��Vo�K��Gp풯�[P:#�6�v�m-�����hxzXn�`�O��Bv��7����������]d��P�E0vf�,��)Zq&TF>^�m�ċ���jZ�R��>ث�VQ3a���c|̂��I��7���^ʭ��FE,,[�L�<)@z*����m�k!⎜�kc}�Ʉ��+�tH��K���`c*�|����s�� �{��&��
�>��'�i�Iy�y� e�i)�H���}B��b��\ڹ�ۦ��4a[,�;�w
Ů�1`9w2�>��@�Qz�D/r�z��-l��;D���.N~��������H&e��ńoT�v����Q�����=���\0d͕���>���\^d#�I	�1�FC	�̗�>{�_{�p!�{��\�hn){;�"x�S��3]�g.o�����l�bqv��]�ˏ��]��ϛ�7~��`F��]�����с5�ᎇ��=�����g.�)֪2���O�I/m�k�\P�-m9�T��}v��03�&���?U��n�;k�eU$��4C'wwgjz�#�2�����&���'vU�ꆚK æ�sd6J%n�fX6HAW�����A���.�n����%pU�I�el������Y�ꥵ��WG-i����@]wdFe�Z��IHKu_��˗�]�-�r�ݼ���7�toZp��l��ρ���}�g�}�*�/�ۙF�S�Pf����kK�X�J�SF����7�]
�)�TX{���.S
��J/��Z��&�Q�Kkdg�&3j1P���pCy	-{�Z�".�ݜ���K��添���M������#�!�1��8�}���=����8s�[��*8��t��o2��I���:�-�+�Yj�t��Ao�
3F���!�g����ѥY�G���WT�%��3�5��������GIr>Vġ7�8c�gY�c�˲k��uMF;��H��-"�/4��-N�5�C8�b��7^�K�˒K���x#Tw�F��3�8ً�F-W���#%��X;nD�A�d�vQHZ�u��EX2N��Ƶ,9�g��c.�ɕ7 ݍ�5��CN��ooRe�|:��a��e`���G0X�\�-2;�����$t�%gr�֜t��e��;��	�����r�2��j c�V8��(�$oObꌧk]���2���G2�ځN��m���{Wǐ�f���ɤ�5R[l'�:*M˷Z�~LǏ�b���TVA�h6��$<�-8F�"��K캠�0�.�o�gX��os٢�H����\�|E�5�&a�虪��=%�1ԛ��;��|�X[[�7;tsm@���i���c��C�������k��ݦw@��O"�zd�͢4�
L��LH�ڒ�7ǻ/���gUM5k�A�~��v@EW0������=Zmu��Yw��V'�]����R�))�	)�,A��}) �
�p[��e�:Gx|%�Z�$hU�d��,`2�1E�}=ִ��v���Tvw�j�,=0��}L�v��<����[�9�a��F],-9Y�1wֵV��F�[B�U�r׆�M�ו���<��0��ɚ[V�&;��8-�wa�nn��{d00a�z)�H��EI��|S0qPѠ�&�=���Ӿ��}���ǝv�j�j�f����f�w�E-�z��,p�&�mo�L�J6�f��B��w�����Ȱ��Uo�����l��v��ͮ��&�8v6��v�+�'�[duC��a98n��2� ���b-���3�9�=�e �����B6�x6k��z�n�� �fF�f9M%�Ve�m4�㎦��r��F룖93����5W�kk{� 	^� �\9�>~��\&;���`!�"�ÃxS����B��2�����g�Y{�Z4)��쨻�;RZm�N=F��'[�k5���c�}���l�7$�%�4d��������;!����w�_M5���8#��d�� ���R�p��B\��;��v^H�/��u�������8o��SL�otx;����:wi0�M�6��Z�̰O�}����'x�4��n2"gw��a���ׇ91�:�}}|k��_Gֵ�kZ�Ʊ�k^<x�{���������c���<��Y�e��_S#��9H��JY����������_G���ֵ�kZ5�kǏ5��턐�0�����$����n{o)��Gg��!$�~8�_^�Z���>�������kF��x��ƾ�;��.�&��ˤ�$Dd}g4�א�ɳ�y!	$�I'�<q�����ƽ������������hֵ�<x�ׯ<���*�#�Ni��g4�,7��DG5ԉ6�$ɐ��5�h|�x�gt�3]���S�d0|�BH�@:Q�*@U��b~�N&��DM�O�oQ7�r�"	�ɴ֕�}�H`���� �AE��m)�9<r"qrwz�,��&�$�zө��DI��O[:�e�N��d$H�"H�'Z�H��hE��x(��~i�٥����_�6�7dK�-��5���W��;{�e뵜^�F���}Jhݗ
��T�����q�81�1�)�^����^�T�}7o���^�3���8�|�ݏ�a�?w2x�>�B��o֞~!g�����e��Ҁ��!�d-��v,[�9�\B�����Bh�����a��:sl<D����R�=�0yO5��w��7���|��mi�2���觩Q��Q!�?b�k���x�^���7�O�����Ԧ���u�ȧp =�h�x7'ywa�����@�~��󈎒;���dBB7����w���(F\����40�=�`$0�*:]�`"�������U��~��y������e���������x�ְ�oliÓ�cz|'|��� ��ƖE�;���kގ��[��;���d�a������0C� ��}li�%��K�ݾ�����v.@�P�ˎn�m�Т�o��~ x���ˀ�̯������ǝ.�^��syS�Ҁc�%�p8�i��{ծ�w��������,*�O(�������6���`0s��\�ܷ0�^���[$_���i�v��g������̜��|��xo���	��0���{h� ��qpmtn����qcg�ش�}���q4Gw��B2S��E�o��M]�{m^�P���gC�B>�4�cQ��9ʝr/U7je,qq|/^ok5>�z��BW=S�����\�ӭ흏�����ΰ�>s�n�эc�fq�1�0���sv������.u�'^�����^�!�dw/	����A�K|}~���c��|�3��G���^N�G��{�Q�]�;V����H��e�|�~x/����Y���U;�=>�����܈�E���6�I�N�#��?��ڲ��qy�&&�����\C� 0mc�D���Fv��_-Kp��x{�����5d����~8}�K��!��}4Á`'���&�����#����]5�����T����7��4v� "�s�o1k@w�?��J�~��/ɍ�f� �cZ�W��{h�� {l:`8S�no�T?��-�xE���\�ƾ�<��U��uܾ��>�\�*�tVv�]��)8�������/t�0H�PdXJ?|��i4P
z-��l�_oSv���j���{�v�˸ƶ��ڪ��L����ɽ@'�~w�Q(Ŏ~���]|�˴�>�.Ui�v�#p����Q-�ܰ~z�����{���-�:>g��	^��u��Q��P���o]D�$�R������)�����e7���_Ů3'�?ƕ���+���=<.1ݛցXoi����j�cW\�o&_��2�rG�޻eM�y,)�H$�76P��^�i��B���"�h(�hl�	5V�xȤD����m�x�C�+'�VCw�#�h�������N���/�k��ާ���qf6b����â�eR,�W�$�B�h��h�ߤ�d�dHF��x�|B>Lpc�0c��βL�ɜ7���=�>���N�:i�6a�T�ٟ�N{�=�S���,Z�@�'���
�
y��.y6�N�����j�� uQ����dl$+�"��)? ���U0�`#����`zy�&��G~S�+^lf����IƷ����q��Yz	U��K#?�Έ���ԃ��G��Vz��2��!V����l������[�-���l`�W�u�vc�r�`	Y~��,~_���mg�5m��Y��9w��o�}��Z���tٯ�n��XH	L��T7�3���e�����3�4�\nA�vZ����&	�9�y����a qZIa"�ۺ�P�5���\8��IY��O^fq���	���=�<��`�0�j�[������v���q�T�^�!�MƖ���wg*�q��m�)C��rD���%��_���6@���&M̧c�\��[�e����t1<H�$8>��|�/�{��� ~�|I�����<�V�Će�6�3\
�L��Pj�+�W�����d���{�a����Ӑ��{��G���!��|�!����]UNu���Ճn��T�o��4����!W�@w�iU�t���r�ʯ�a;O��.����8�:�ʃW/?��ޏ;n����';- /1tY�r�w��8rU8��ż�瓄�J��I�3OWΰ�ra�cӃ�1��0��0H|y+[�2�?�zp�ώ��6=�L�d�N��Ylv�q"�9��33r�L�(���� ����/I頝)���U�`'��/���^��}���<`�w���֠(�&��wz�������ljoT�xoS�f���Ǽ�2p�Ϛ]~A{�O'$�����	��涘�h*!�ӎ8+�� �{-�W�4� Ènl`;j=�D/5c�C_����j~��蛘q��y��GP�5<?z�xP$�R�3Լ>�O�������dǇ-��4
{`"Ё$�uD�
�q�_Y<<���,1h)�x^�7��i�~���X���_�@\t?�eO`%�*ed���uU��uz�� G~|̒<q�|�:�:�>�c�$��߿~}�w</�KL���������m_MN�����4À�i�q�|�0���"�"b�P�D3v�������� �Ǟ��fL���rU�u�ҍ�^��{F8�D��+�ZS�j
O��s�QM�0Al�>�0���(�l�U��P��h����k&��>0������^t�k8��~��@�u��w��e�>�;��p���ٳ���	�PL�2��.�"c�S���B��"M�:��%&��.�Һm�3q���sk�mν*��O�������)5άl��su�|��e`���n�i��$��[�0c���0�<��z�ߞ����<a��~�~	���^���t�1oML	np/%0�1>osn4����y-�P8:��h�ɘ5�k	f��p�����&>���Z���'��\��\��{'���<��r_�����fk��W��j�h]�n0���"y� ����p�m�y5R�\����O�������y���n�hߘ��P1*�����礶�]U�y��g��e�%"�����䉦D$�~ӑO~��7�|��>v���g����,׊o�>�N��I���%���-��4Tc0�;/M�v@��yԷ�M�7�{�Aa���4��!C��Mo{�y�|��7O��1}����f��@^/�?o�� 5��6��G����1�V#H$����~sp�o���J���c�{��Tz[��l8�S�V�0~���F�f�̀���'C��rz/���~�Ӟ>��W��r'���{�}ćS�R3�p��Eڜ΃��]�Ԟ��!�;��憬���B�A����Y�Wdך��`���V��5����S�rc�������<����<�ϙdJ������ps��n�Z7�ML�)��giV_^{y_��j��K�^LL%]�s:�]N��&q���_k`n�s��˶�sor�Uf�e��������8�8Ŝ޺����>N������K�W��;���-e�syˆ�wwJjg^ܟ;��������w�j�W[y�i?�G����?S������J_g����������������Tl�65\u�=��0.�8=�p�&��󷸽���<���Aސ��y�M�b���Ϫ���ٛ�[��y'�u|��%�����4[o�E��c��g<C��lfRhw��,�`��%mq9�����q�WxzK���T� m>�z��ƐUJ������7�N���n6Y%�'�J1�]RK,�K�����O01�*@��������+�l���@Fql�^���`|��m��ζ��PL�s E?K�ou������>���>�n��=�P�� �ٿ�ԞL��}��&�m�Ǧ�,X	�{�+�u�s�ok�K	��2Y�nX�tɵ�u�����j��YU#��9�j`�잀i`�~a�dW��Ż���=�C�Vw_����fjx"�����>�2�qM^��WQ��I[�zӀ|�\=7��}!I�%�ސ q��}��a��?�����o���E�Ev(�������5�nB�b�L�Tj6u Z֞G���O'<i��*��6F��<��K/ȡ!�2IQ���D�z����v�$*�]���� c�	�J��
淫���1=�:@����C�aOGV��o���Џ�9#,Sa��@[M�6|A�BY3u�7SN���9���U�ZU�4�������]�w�Jv�����$��]�D��}�:xX3���x| �)=����/�$��M� ^r�tݯ�q�����0�[�{Z<_X�-�������b����7d��_#�՜T� �w8�X�v�S�[{�c��7�Ԟ�ttx.�S�N��q�y���	���IB��4��_K����t�����S�����v�9�q0��1^��V��V8|s���H�M� ��MsJ76Ҭ[�����ڽ�48s�z�Y���7��;��ǳ����ĵ4ۦ9pҹ���[�Yo-���	�쌾Զ���q�=���b�?y陎�B�����6x��q��͌b*B}O/':�0��������1�:����1e��`�34;P�>?�0?޿N;m������SY6�2�(�^��Xp,��E���w�E�.��txaؽv`�>�4�b{�:2Qi���������^���o�D�"	l�l�����ϒE)�[����Ϭe&n
�����Xۮs��,h#>�� n@�.���hp�U��Vx`a8�[Ý�9�OH��
�6�k�!ٝ�=n�����韯�����n��k?d:��lSw�mS^��ʖq;n��g6�����ͤ��ӣV`���"^��8���k�o�<ʾM2r}o��"��ݜ��̝w&E���۸4�̇��_<�s���=�����!�ǌ�x��81�#�o��z���>��$��ך���uOj�r� ~`\�"A�֦��@9��}�f���o�總^m_䫀�ـ1����Sx`���0(��p�֠��p��;�N��q���1�����Y��T�n��Y�)p,'hΰ�_��z�Ҡ�C�k��ϐS���$�|���D��?w�j&C�6���n~��.ʜ	a��1p��{�-�n�R<�CA�QQ'�s�x�H��ȓ�x�zw�g՜wp�<W���7�
y`@�y���H>O`��~i/���u{���8.��*(TLU��G����>@��_�Z�Z����U�@����AtTB��b���>[���Z_�~�y��=�%�K�� �����x�H��s�C�����k�p =7!P�K -��4淂z�8�+nn����)w�{q�����?N@=z}�&a�z xo8p�q��dy��Y����Y՘��\�Ǣ�E��Fn�0��'��`�>�z��l}�t�s@��q<ȃ�<ܩ��t��a�8[����ĸ������w�w^�=���8��ޞ~O��n�� ��c0ʵ{~��dVc��qv�H�v��_+����2h�1�}v�� �D���կ���Η�0�?W�ԭ{�:�Ǜ}��%�v쳺�,Z3�v�a��k����_b�~}�!�u���Y�Pw7|ߝrs��1����ǌ��38�Ȍ#	$�#�u~���ϿA���t{�gz��Q�=% o���u�0�`a�SG>���		�2��-n�1n�嫀��#<
�$���fׇE���ߗ��k�s^m�n��W� �����5;�lWp �?3Up�ze�N8��@}ǣ�Z���;�n�������׋�>ߞҊ�Sz���w��[f��s����7��?�����������7��'y�i�7z|.�zN��P�-�m�r��O��-T�w7\�;-��ɴT�ȿ��� �O��'��B�����"|t�g�����/�o�Xv�=��;���)��-��\����1UH��Ő���@>'밊K�l^�\�r������R;u%�^K���V.�O>*���`+Ă^ְ�I�@i��j���x3>������Y�bD�����`A~�d� ����C��� �+���}���|��+��%���{�fލ����<Cci�t׵{ϭ~?���n��R� ��P�v��?n����(~���4���*O�Cn#�ƣ�L��5l h^�D�i���sG��K�:Y��eё���3��9�]�{^�Sn�^���)���
��(��^�|� 2���̛;�_��F��ӻZRM��aɵ˔�=$ĐI��A�	�",�0�<�__[��Z��O2nj\�fsĲv�kk��u��	�����S�������N�$�	�~ ~�#�88��<<x!��Ǌ�U�X�@�	$@6����{�����L����ݺP)zqɡ���w�o�b)�L��2��y��rWCp�{Cߺ�����-�#X �|/��B�
�`C���hN(������VGw��[��`�շgN��a�CBқ����or~'_y�����fB�i�=N"���k*<7C�W�lӜ{:��q��ɇHY:��r7��_��q���¼(�-}jOl�^����'�gnNDFZ<xPhY��c�O�~"_��̊o�����k�~�����涸ܑ|;!�;KV���D �������n�E�L�%���0�q��=P�J�'<��6d���}k+b����=e�~�ު
ߑ��+#����S���ނ�8���t ����5�{v��b�X��,��ޮeZN����[xQp�������8�q��-�Sf��P�7��J�\/K�[Ŷ�@���q����� ����
�4��mߘ�����Ǔ��Rtl�K��Nf�*\�N���C�|iڱ�t
���d�ȟ4��^��Y�;�L=�"w�h� p�������:���$���
pS�Y�	+K3��Lܱ������lvtr�tр�� Y�&l4�"5��f�n�����Y{�XS4�u�Ek&r/y���>�`�է��N�qØ�l��"�:��W����8<��&���Κr!��{�[�5ُ�p�t��M�Uǋ� RJݰ㨯w��H��yYz6���HH0a��/wkZ�'_�D�/�,��bǗ��i��Ն�b�bd���E�m�}r
&���<��Mv�W&t.��h�ǭ���������e���cpL�{C%��a��{�v$�A����Y����:j.ar�>t+���������{:�3���«��^I����uaO�eUY7�m`2m@��ƒ*kikx�Zѥ8��Ԃ�ձ��9�^�,��5�\Siz]���1ɱp�:��h����-r:��Ê���˅K�B�n��dΔӦ�sK�����{�V�l��{cS�h��o{~��ānS��Q�T���FӺ��2����p�w�g��8]�|gq�׹(|�׶-#s��-U�kma�
����RM)d&S׊o
��(���Oe/��/���!�1�z�2 ��=��)g��m�bc�X�x�Ĺ`��Аl�WiB�,�
�,�{D"��:�dw��ƛ�Y�i:ղȳ��^�Ȋ�_�b<j�����l�g�ʓ2ĒEA���!����TV	(]��@�u3Y�n��]�YVK��vVH��mh1�qbg�?}f���k�_��v9���S��G�����=�ם��D/�]n�<a��؏q�lYM�Sxr�T��'�&g(�:9ۉJx��,P�{��w%�ڿ�4�޽�j*s-��Z}QG�Y}��dV�g��e����;7W4��N����ЖvL��β{�V4�GT��ViXp���sc�j�K���uS5��Y��Yɢ��Js[�n�΂�٥�v�x{wd�{Vn޻CFc���:�tu3~��*�K��`VZx�6'e8��pR�F>c�R
���ݻ�r�]�v��YS3&`wbLr��"*���o[*����V���c�F����>[6C봻	��k���Vsc|��l1\�Lw��+|+DK'�G�S9{c.V�ubn���wpM�IU���<�`�R��������[�Ք�;Έk��{��2F��_
^س˦�1��YS���~�KU��Օ��)�9v��Ю���{o��E}�"Yy5�L�J�z�{�.�鎓�`f��ү>���A��*\�
(�xP�Q6X�R����+hD��3BFr�pD)t�Sֱ�B�H�DĈ(���5L#@傩�KϮ�
vo���H'L�S<�$t2���HH��L�'�i�V,�1̌�� ���2��f�V.�Fq+F��h5��c)$|YF"FGF�ۢ��iX@��)�H�FD�~�ə���O��=���r��D�̬��
&o��˟>��X��ǭ�fI�2�<c������k�Z���������־�kZ��Ǎ}z巒����6���vz^^i��曮��0��sy�s0�1��8㯯�O�k�ZƵ�������}__Z��Ǎ����1|&$��*�D�km_��'L�>V���Fޭ�i����fL�΃8������^��5�k____Z�>����x������'s+�i��Q6�O�Kr:��2��$�E��u���������ZƵ�kZ�־�������������޲ �o��Bm�_�d�����fۉ��M���N"*$B��Dy��R��C�a&�9�'L����vT����mw���:l�999��m���TB�g<r/5iͧ<���h��lm�h�~��ք|�#��m�myX=�sM���*q~c�A���$�|"�'��$&�IB�MJB�����I��l���LH6�{ӄ9�&�m4�_i��i���c�@TA�@'� 	�6P-y{l�E��S�4�V�����\��'9MN0�C�-�F�U�K�Y�w6^��5n��gv�ݨ�K�v�#��a�WF&U�]�!��T�a$M�A�8mH���%�%��vdP�\��L��9�M�һ>�5�ǃ�&A^<xǌx�9AF{��e-SZ�9��;����EL��LՏ�"<�ת$>b��?A(��,?�]���́f��_b��c��ն�鲯�6�w�`7{<� �3�	����?]y���g6�VϿ�Ff��=��Ũ,k�+��A����x�6�4�<�'XW�D��gl� ���0�����5��"q�8Pl(d��b"v.2�(��G�=�D��?W���IB!x@q�V~�~b���W��{�����>��7��ף�/[sZ�FE麱���pX��NKy���� 3@O�;��9��\3?�P'��x3K �̴�r-��mp2������q����xoL ��`�����Ɛ��s�������<��F/ϡ���I:����}�	�Ǧ�pV5[I�p�~�`5�k�i��v�z������r��C3���;�nŀ���}���4?������ւ�Q+�)�hC���� w���>��i	�b'~w3����L��-�,0��=^7�|�N��}^x�-��N��{g�!>��ks
��^�����qsزH�_et���<TǄc�\_�+�9�`j�s�g�,ϿG��c@a�\Cvt��Ԥ_���⦆��m��:���}x�m+��v���u���$%�)�e�%��_#r>�h��:��Ŏ�,)�ΐ�B.��R��#=�;W>ي�NPXk+�y�:*ڼ��I�3�w�9{���[����x�ȃ#��≏����<q�' "�H!"�w�_g}{���}g�X~xu<��J������S����N��#����4�`}�[������U�!2a=�xvOV�'\�x5w�-�*M�����S�������<1��xn�gמ}���=4�{�]:�f5V�n��q�y6�v���]��)����Z��w=j�ŽE.�a�p��M0�p��귩O\��a��p�r�<@o�g�[��Ý�sBKzF[����[��zv�J1�Om�4�C��hi��u�\�p>�a�/�#��!%�ټׇP>�}�O�ϥŁ��nOE�^��a��}�WS_���b}3�ͳ�\�]��0��H��:\���C�uϪM������X�Ǳ��B�U�%���������l��p�CW��@�x�E� 3?��H����7C�@fk���u��&d�wj������K	�d7y�=���1�`�"X$K@D�Bh_�o�"��~������}�y5��K�2ڹf��)��p��n�����{= Y�C�a�VRy�=���]��`�̘;��u�;�<���u��g�C�>��kW��^���O��P�C?F8L��pg�ѳ�V�}�o�r���L`Oj��p߶�Ö���wTڿ��ƃA٥f�\O���y7k�6���s�D�-x3�{[O���ά�]��)u�H�ynv�׫9+��}:� �h��F�P,��� ��zx��+��������q�<xp���" x��$�\�<��P�{^_��b5�#���T|��.�+�C�����D���h��T���!ڹ_.'��,��)g�o%'��E?��6?/��e�TR�r<���^g3���~�{+u�a�r��OF��q���dg�	�a�	�c(X�m!��|s~	�fND��%�����/��)�}ת��P�����v|�U����b���������q�)Tҗ���ݮZe��D�DLG�����:�޸q�[$\&���� �f�M�Wg�\O��xQ��������͌�G���}�8ޏ;�` �6j1�)��+5��^m�n���
V�e�Z�4���m�����<��0�䁡��?y�� ��|�}O����*�E����9���'�}jESSJ��WW�����}n��;X��Mq��0��w�u^�-�7��*��:�5�6�����k��`5�pΡ��q���z����	�����
���*8����b[��5�ǖ�ނ�_L�\��U����^��-E�X#ʪFP��F8`ζ��~d����{�q���ݘ�]9*�[qZ���GՕ��{��h2*��"�k���iS���_t#uN�on4aɝ!�vZ�9���b��%�Ky=���0f�۲�2�t�t��Τʪ��ﺬ�/:���iڤ�����$E��� @�1���Y$�1��ǌx�G�������x޿P��� φK<���������>�(�w{�(��xxX��8��F��G8X`(��K��0>Ö�w+���l����B� s���*���1HU�\��fv���.v��޲� �'�=L���4-�!0 x3i�\n���sL;�#G�ND��f��}����V��j��Xa�?�P�ʅ/~Qk��2�>,P4��6U�y��y�L2aVউRvVen�pI�0J�a���p:-�c�qb5�>��
=���z^i��c+�xUm}�p�=#ñ�5�:���1�>�6^���� oL�P�x��|��0@�*xψ�������ݘ+��ԕ�����+;�/6��;�z�x|'�XX8�� �������/�֥������s�y��}�
D[	�k�א����>_m����흮d񔪽l(¸��Ĝp,������B�������([�?+8p�r��:=�ܽ��m�U{�C�]�"i��oP�x��y��$C�~��_�P�����W���J{�-s,�yV^*���T%��۷�E�y�����Ė�����T��1UWnv߹[�I�F��gۓյ=G�T$��*���lSeFQ~mGE�yhAm�*�S���rN�.�PH���Џ�b�3GRzm�7��W����:�-�w:�2����~���i�m�Q��T~o��fNs'8p����Ƿ�����*c�<x�
q�<x
�"�x�xxx]���n�՛���� �T��z��������v���7�����d[xG>��h�W�r���5=�B�<%1�[�l�s�M���@pƸ�[�ֹA@��vǺj1,9?�j�}���;D[0����t�f������;�?9lV��;��<4�m *�:��H�s�b��K���������"OV�C���t��,2_r�㷷�W��|������a>���plv����t��Tg��l��<'#��U�-7.մ�0��A��4!~������0��������8�������.D�n�8� 9�����zDfYgfwr�Ŀ�I�ӌ ;�8M�i�SW��7>`�>
}q�p���"XN?�#Q��ne6�c��{߾V~ i�>����'�XsKek��8gtަ͘	�Eǃ[�r��y�/`+����G���c�7�����KG����5���b�c�Zhߕy�(�{�_E�M��V(՟+���~�^ذ  �@\G�8����;sS��7��*� 8���<�	�s���򡸑����L^�1���`N<K�:���\_lW�Bw�.�]�F�-�I6�Ed/Տ�X�2�2A�G�ψ�����↵����r]���M�I�0�h�Mh�M'`&�}R,�u�d��Y�g�]=�B�Y�v�\ա�Ee��`���n�m���[fA��]������;��;͝w3�\3?�폯G1����x�q�<D�I	 VEYG�|�}�}��h� |���D=�d[��ڨ��M��w��Hi�Q�&���
��ux��-�r�ӪmT^\mD]goZ�<u�zp�θ�O�]��\���dOO��61�Ms$���\��=}�l <�彞a����jڋ����p�a�c�v"y�A]�����Z�1�fCs�6��o(������h7�y��8��l��&����,�1����������얐Vi��NV���<[Æ���\&���\����]����1��ln`m[K`���5�խU�y0�ɇ�:c���p/LV��ދ�n�G���p���{��\m��4j���_�|���߾�yc�JG��q�Ϋ�i$�p���+(Q���W�s���mGs�PXH�Cgo�I�Du�+������.<��7�8,Za̺�27��3y0��������*�5�,��84�y�c���q�����ޝ���	^�����/գ���wS~ C���'3�	��Ǻ;���L6�{23�7�o�q�V{)�M#�L:l�{�`�G���@�w��P��vT&݌*q�W[�W�y���j�a�Ꮭ��{����j�Q&�n1j����;��f����� ���Iҕ�� �\�'N��w+�y���w�����w0��[+���A��d����^Ad��D���~� LxǏ^D@�x�Dq�<9T���y[���� F���\G?���z= �@��J�^��(����j�7�!�L�0Wpx�$�ř��降y[����4>t��U��H���7��yw��2�m�v�n�<u���^�
���SV@߭�C7v\��@L��t�5x����xmr�:\Ȯt�)6?���i�&�2I�O���k��m\W���5�U ]����3��kzvw�wv�7n��l驍%�0D�M5�����}����
�a�1�/�����ؗd
�
h��������x�1FV^�oR�T�ɶ� S��wZ*)��  ���Ý3���4�F��(a�Y��on'��o�������{(��x��ˤ�+��Έ~B�6�cʫ��d"�����s��B|$c�tz�_�\��K��ё>��z�o�!��(@�h�n�g"kzyrG���K�	��Z��`
<,[��+�y�w�m��<�)��]s
#����7�������n�E��~日U�I�<W��ݢ#�]�z���ޙ�*t{֥޵������yp<�/�����'�_�����ehjV�o�\ �&2����.�h���u�lD�����Z�lm虚T��*�O�!�82pW�Y<H��Ry���DbjS�Kw�;(@�ٍ�fcd���:L;'t���|�{�j� ���zx�� �<cǈ.<c�=� ��n�����<Z����z�;@ז ���<y��Z�ƪ�O��rz���z��E��;T�elj6��N1�����f���[����*��ii���G�i����k��i ވz}'��Wv;S�������dX	�!JiW��_��+�����(�[k�j�7HC�~_�G��ɝ���5�z�ż��d�y�a�i���=��^z
.|6�[� g�>��PBG��$�>��Ȼ6�
ɘ�7z�4�1޷wQᘺ'e��[��|�=0_����Fj���7]��ԥߩa��<���}��`鷟e۟{Ւ=�q\�A���a�/����1jƧ��z��e�C�p���D�|a����_=/��Y5�v�O�)�y�ۭ�@������."����mr�֝���f=���_��g��_��e���~ ~�R��=��3�k)궘�Oe�j��{f������!����~��M��L��X��p��X	it?���:����z�����a�)�n���x����i���-�V��*�q9�ao	G���o�@`��_��T�G�}����#�2c��Ǟ�����粲V���`���-��6�;��սt4(�N��Ni��h������7si��N� UN�� I9G����Ѹ6h��L��$mN��g9�5�Ⱥﳺ�rҮ{�S����u3e�E�Vm�I`��i� E2"�9Qğrs��g	��d��?c��Tǌx�1�<q�<@@ޱ��[��w��{�h�#���FIz�����
�<�s[�d�ߕ��q�[��s	���{ǌz�3Ty���5��f���t����q}�%�!�->���
r ֏k��qlC�cbJ��]�#�&|y^A�����������`��,Xϑ����~R|�`p��K�1�
v�s�i��9~����x6��wr�A��]��a[W���u1�լ�����8a-��2�!�����0ގ�8�5n�n���X�����8���oJ1e���zF�0��^�c��)��5 �;_�y�aɷ�G��lդmnr`V�t��<!�>c�6�瑴i�o�h��.�����V����\��8Cr�X��.���Ev�TJ^�����u����~��a@���I?e��CΉ/E�W�n} [y����m��-Uᐹ�$VFs�
�;*��w��Z�'CMt3�E����u�p�$����V�08���<?���{�o���k���EnG�|�h{g�u��T�ʋ��7�V�W��Ͼr��:���,��XI�G�z7Ft����A�� K�ؓ!�v����׹&�l�~�W����K��ҥ,,�#�6{�w�
_^��e�wcq��E5�B�-LAXC#	���h�!�<��� �~�	NN��q�6�_\�t��u��k�5jѫV�\�w��r��p��{� ��N��z�8[ǣ�2�T�=��o[��޾^��y��|�'���ƼPx�c<Qq�<q�<�@�A�p��b��;��V0�%����T;�5xcf�]��7��،i�-�}m��Y��򺦼�����k�y��z]��C�׊3�= KTx	�RO�7ō�ك\]\&�3���s0LT�╯o,����?\}-_?9���^� �0�Ǿ���؈v{� ���y<�]og+����[�S35�/�ѕ>�lc�<sT��z�5�<ʅ��*���Mtۮ�]��i~��eo��Q1�ژ�v���}<X����� c�P���ٹ�n2��u
���h��_a�@�ꋗ��z�38�⢄ S�T����2����=��K7l#��س߶�i�G�W�տ���W�)�䁾�1x�L=���PU�����{���滘�%9���z�s�cԮ�������nS��vFyo�ҷ�da#���� ��=V/�M��!������=�4����ݻg�5�*�w�NZ���1�<�/��V����|u jzw�x`[Ç=1����`�̛�ս���CE��0NL0���ݮF�y��t��}�ߐ����3��� u���I�g˛�!�M���mq"���R�c��rfü+�h���u�%�.���t��ڴ�p��o:�1kk��Z&H�7vhH-K�����+%���h6L"�pF�`��8��B�n�H�"�9Ԃ A;�r����:��B�+r���LW_oKwZ�:+�^D�KJn�-7�����5�P�Zy]יe\�VǌKp�<:�h�@��}.�;�Uu�`��ծ3�۽���T��'!��V��d�K�F�v�
�d��'f�5�����P��q��gy�-s8�᧚����j�W+�L��ty�C�Z�!w�gb5�!�N/dۢFYх�[ԧ�����C�\8H%�b)7�fy�d����sU3U�sa�3Y�TnK���ttHЕf��e^ꛆm����V�74cvk��嵽�Z]�V-t�d�������;�QuX�5H��ef\|�u����xz[r�:�9!�l3�8ŧt�Tĵ�c��}�5ίfh}��]~8Nm�w�s�y,��x_m�
uo�k<����˗����"%����U u�7V�C8�Rt��_Z����9��2*�|�j'O��ŹƜ13�?q�I��Ƴgk��{͉�ܢUAC�W���;��� ��1Ծ���}���ZV�Fm�T^���N��m��[Z,5m[n7<�JS8	t��'}Z�`�Ԫb��w+o���)�������,�@�w�4V+����������3��{1��+�&kV|����=�S1���_��:�l�P��9>eotsP�Y�ӗk�j���^��w�TXGN���D|�m��D����ͥ��VSb���s�)F�7�Vm��ۨ�Պ>��C���έ4��M�]oo:��[A�ݻ%�2���"�ޣl�X��<+37\v��fF���d;�`]����L�B�r}�Tm��8Ԃ��6�	[(&�h�r7�+�0�F���1�G��W�����T;J��c���^�X���\�K�]�I�f��;�ԾוT�U�;��8ā�o��_J޼��m�)�֭CN}����tV�M�4�}��1Ru*C����:8�{xh�Yc{�ii}I6��$�X��؎��+���k��TMɎ�K��ϭ���ڽ�VAS����q�t���д>���b�
�T��ꂷ���a=d!}rk�������.�7��o�(:���R�6�m����� �=�����Wշ�A��x�Y@A���ߩ�6��-�$!b�79�T�����'4�&�C�8�x����ֽ5�q�kZֽ�}}}}}x������d����$��#ֹ	x�y�b$+�uԜTN�d�'��ں�y}߷���^�ֵָ�k^�5���������_^�|�*!�����&�Y�#�dӫ|Y8����!��[�DW6���ˮ���o��_^�ֵָ�k^��5�}~=�����׺O�Dy�F�?9̉��w��#i�'l�TC�j��dL��=Ye��������	�w����c�O�����~5�q�kZֽ��kZ��u�__�}͘������:�&%�AO�B(�擎%��,�-��1<���Q`�A:��� �)���=rzwktm2%)+�A8�<�qtHJ���OM!L�q�G��x��޴�B �B-:�s��}r��s�uK�طF�zMV����x�i��g&��d������0�R��x�ڶ�*�E
��"�2��)2h�$!y�['9�e����MTZ����Hmg:�?p��]f������S����֞%^�}�׉Ɔ��;U�Vo��@�� ������y�����+������r"�����k��߂�W��b���nO7���� ���;bO��zOT0�n�}f��;�[ŇK�@gǗq�,�����E�P62;�U2��S�r�g��o��۹}�n	�a�ߘi�&1x�?ާ�^/�P������p/�=��Kך�-�_��ؾY\[����P����k��ÿ���/8~�?_�0���B ����4��t��;k�7wF���"7��)�\g5�o-��w��M�`$�� '��_�����y�;-}�����^uipR� C�O|� �)�s��(�Vc7�ܮu��$���L"�	w��εF,7��ۇE��<h�NVE5gO���(����v�PN�����u<ʹ��^Y5O|� �~�(_r@�D_�>A~Y�@C�0�~��/:���!-�B髲H�a�Yѯ7�{l���幤���_:+�χ޿�����e��+�5>z�ឹ���1�M4u�m_EE������ϣ�����.�g��j%�mB�p�h�Кa��->�,4�r���n�ț���ZZx�/6EdF���$��O�<�iۀ��m��k���h�!gn}�����h"��/>�ӑNlR**9�N�>q��d�n>7�+4�刹�q���/���z�
�'4y�Y��l��;D�7�im��ݧ���|����G��ǈ�<cǈ���q���"�� ���յkﳰo7��q�)�'ʽ�8�h?����uY��f��	���QL��斸5z�}��9�v����#����/D^i�_��Kk&@oN���`����r�����@Z$����BϞ������\J��](�(H:/%?~�槺Q�_���Bm�&�y����ǟS��������k�xIS�l���o3���[�:<-��[����'�V~eHߏ�����5u��no<eܝfz���̘�ک��Y[�7��w�Xw��:�0 J�h���g�%�pX�z�W<��ٮsܧ�~;}c���vӍ�ז�Q��������9ĐsW�����O���!����W�W��p6�擄�g���z�s7k���	��Ȼz��x�uwW�+�l{m���'����P�J��M�_���6��K��v�w٦��5�L�33>�dT�xH��z��S�������l1�4���۵��SD>��'7�6{k��)V��A���!V}����~fn��Ӟ�׋����ǰ6�;}�ߴ�	VB�V|������0��W�\��չ2!����dC�kGpv�M�>uM�^%oz-����B�:�"��ʣ���p]��Bt��^Vǽ��o}�Ӷ�́�EMQ���)J9��㻪H����t�=�t��
Z�3�83v��ufl�z��M�E7v>�U���w�ƛ�&��1�D'�4�P��U0��iUD���3&�0�݇:����>���<x��R<x��<x��A��� =7[�_*�^oX�;/�XW���?�H��C�����0i�p9��.i=�\n��Q,=���r~�nz��'�vVoQ#�7���_�@ǖ[�=x���
�ƶC��D<��^O��[�v�k]�N��F0�p7�®\K��n�`'�o̙�����3��1�� ��e��|�z+y+Z��Sw=0#-��V/_���a�@��S{6��z-�?�/5F�5��lc����U���C��~�~������?1G�s����>[�0-���˵4K���	�^Շ�r���,|�pL�|3V����s��E�Z���cH��c�ݝ�zMZ���@~��(�T���/�v�Hi/� �e������~����y��ڷ�m��r�]	���Ժ�-m~�oG�������q�⛻�=y�!��X(�<�zv��~ �C�}�G�G�W�O}��X;��[�a}V�\�U�υu�L��Q�����U�!_����׈Qω
�,����@��w���>�o��ְ��C��s<���M+y�m�0V�(,�x9���(��7��-6�eLV}w^�c
�-˻��)?�׳��;fӛ�;w(��=��Q�nr� �Z�U�$y�;��Wc��_3��vޯ���Λ����˻O�&�7�]�Ρ�.I���(�1--O�۫�d�ǧ ���|��T�x�q�<q�<q��<q��<���|�~�C�3�}��z��
K��"��6{�'%���'�z���"��о���w������A�x5��e��=����ٟ��Lx�n�`.��7���u��X�G�8��s>��7O#�o�o�����9����Z^�}o���O�mO�yO�ފ[�����)�e����eN���N#�����(;~Q��|ny�����!��]����}]��V��Xr�3���`>,~��$�x1�>C�xq/�vL�ub�tɜ3>��Ӿ�_�������V�x�/_``r�iTx�+<���T�7��I�?b�|ﹷ|�Ufc�_+p;���ldz¦���gE�i�j,"y��m +`��O�����?sv�7Rm�w�=~���跖L��^��TPk&<�L ����V5p�͓�q��o���_���
@K [�}�?�'K1C�!��#��~ B� �o�j#ǥ�3"�=�
��Ζ �!�� w���=�9��Q`~S��b�/߈�=,��~,b����m�uۍ^��y���+Qޒm@J۬<���������fC���b���t뵮��c������my�]}��y7��w�����YhG�ulA��ĉ̛M	�&w峭���ݐ�Q�hrtK0nw�3��ק�(����������y��� \N.�W�=�������9�#״��S������ϻ�xW�g���D����T!�u�	���8�o	llm���_�4z�H�x]��0�k�?I�`/�&��srq�m��O�D������^t����a<�dLX,�1��q\�����N`/A���\V8�U���T��\Ɩ�:V���<o�ڸDx �)�̼ʅ�����8���GD0�Z�sO���my����/.�`��s�]�} �/�q�����A� 2`W<�����f�����'�깺�����m�W�RU��7�|�vl{�w�v~!��^	I~��~��������z����ަ�Ϯ���K���a |��|��a�p����~=<�a�l���u�2Hvx���3x �lU�3	#�.x�O�ywfp�'��UG�G���;�B�^�>��M���<y���3*����8J��j��T��3Y��/�ߏj��}�o��w�oUy���x>Nb���D+�qP�a�$�i��Y�q�������x�1���ߤI�p`��0��v-��|���˼��F��&l������V��=��)�H���l��V��o{�D�����0J�@���i�SV��l�=<Y�v�ӽ���}����P�%�e��-��������Y�N,���Nw�93?������R<x��F<x��Aq�Q�{׾{w�Ϸϼ���G���?��1�X}x��Ӌ�����W��fe7RG<S�w��P���Q-��`�������n�:�������_Z��|@����1��z�VoTx��w`�P �7� 㽝#�E�?'h��ʰ��|�9UO�+_��'�6Ʊ�v����=����܌~���d;��㶩.}� �)��$gy���"9�C�ks$�H���*�8�u0�=zG��]c��6��+k|��b�Z�L�^�1�|��A3g�"�Y�q��� _K^3�oP�j��f��>O^=w�z�N��>Gg-�<���XH��V*;[��w����y��{��Z/l�o�	�����[��
�n�s����f��dCZ��m��mn���˘�A&A��������)��O���>j�X.k�;y����WU���ֺ�>�t���?�Æm�a���m��@���ư�2*x��Cǭ�xox �{S�6�d�N��w�9G�ϖ������ X��L!Ǥhqm�8f��p΍����ݗ,!��
�#sݰAtĻ7�W��-��Ng�N?k�M2��{�,t�hj��4/��wWU�|� �fS񪺶b�ҽط�aތ[۲��ʧ&q��z��v�����m�Ot��;9�|T	��]��x�R�E
t[IB�m"AD�'�:4�~l��~"~8���X��H��I���� ���V��w]���m�������bDpܘCZz�K�9޷M�]�	|�l���A�՘�-�r��{<��.s�D����D�<�� 
e��2y�s�͚����ʹ�k�����;j|.��a �`�fZ���r�G�8���m\l5����������Ⱦ>�C|cH�N�ֿ�2pvK=�g��-�hTr�$I�
��~>����(����1�e��^����0HF�V��nQ�n�Kl��J�z�P6#|��zw���1`��9���]��;y���>�y>�4��\�Z�]\���A�z�#C9��m�Zq�����'��h>z��\}A�)�gŗ�[���K��r�]=���mqDu����i;�{�;2 ϧ�Oo���>9H$�"�0�|�h|e�u��	b(tJ�a��V�Ah}ؾΒO��>w�9�|���S\�P� ƞXs�VE7�+,#�}.�ɵs�.�UP~s���#s��ALO7ԉU	���ݥ��|�6'��@23e��;��@p!e�ߖ��8��c<v2����ڥ��uixO���~�s��.Gp�C�ڬ <\3�[׽����;�drA޲��6@}Yn�J=Q�*z�-������Ƽr����~ƄχC���������e��tD�M����3����ק*�:�e:yN�y�g���@g��;ޥ�4T��pn_=|aN��&�sY?��?��x"G�x�<q�)<q���Mَ�+��8_�X
gk��:< s�qu1�#��%�����a˿q��G^�_n�n��)񑖔@l�o0��޿*���<��5��T��'=E>E�v�w攜���~}�߾���+��Ϟ��2y����z{��g��^���iHu��6J�z]E¸�ʊ�7���7�4cZm����V�/tZ�2�m+y��h#9�qE�K�M~l�q�:���}wy��{����x����ڔ��1���x���݂pl[x�ۍn`5(�z�~w�ɝ�T�Q^l�W�ǯ��=.!�/�>����o�Dς���d�� ���tUϯ���צ6ŷ��.�����ޯ���P�0|��'ͭ!����~ǉxi �����?��_|���쾞�__�&5���av1�j�Y=h���^����[G�ӏ���0g�q� Gyq����Ap� JZl�t,���,d4��8��-�K��e�<�%�0�&@�����o�(��g�Y��5q�lh^��4��c��v��� Kapw;yn�d�Y\��q/}��D��'����C��ㅞ�!�5�/N���{�<�#WJ%�~f�V�9r2ؘ�w)3{Q>.|A�1�9v �b?C��D�w|>�H"�uut�_*�]�G��J2:����!���0�IE�����aZ��m��NB���ݯ���}T����X��cǎ<�8�� z�*X~��+�G��[x���������	��L������r2e�D����c����2���GW�}�MOʧ�*x�����gs��U�T�"f~[��ӄoHI��^#Ӌ��t�ެ��O���U�J/I�3���@�@?~W�2-�g�'�[���̱�`*��krO�[.�U������A�𜘨|�z�C��v���	�M6⣅�AM	oz��&͇#�v9��� r	�z_>����� Yg� YA&i��o�� �-o$��n�&� �S��͵��D�؞����b@�|�+�C���_�7Lqփw���L-���Ƃo`��2��Ő���`��=Mm�$w�(�>5��p\BVyiG;%�:��ל��o�������n�#>�ܔ��,�5�����uja7%�1q���1�Z��� f]耆y�s��l�z����z�]� �4{��= �{���Y��ٜkg�_��/ϑ/Qm#���C�P�r�[�ߘa8��-�[Q��l�!.횉����j�Ǫ�S�xF�><����|�3j~�E�'�7��y����ҽ^�$�(��z1�{�;\�oDV;<en��9N���/��0e1ݶU2 ����$B�P7�M��s�gNsM��!%D���Ġ*���+3dZs�G]bf���G'\![<���9ok,�3�i�L���R���ww���_/}��~��>������8�<x��P�~u~�Ͽ>��~�y�7�>���� ,��~R(�,"I��N`̩�!����2c-��i�%T]Օ�K8���a�O@��ֻ7>�U c�L|Lw0���E�Lg�6�%,�_�H�_�����#�����l�SH���;�f �\�d3�h��p5��h��Ttz|\	q��R[��Ԉ�i�n��h����H	�?z �f��n�O���=	��L��m
��}���	����a�^[��B�pnos\<��
��a��Y�@3�=�c�Nt��Ֆ�����gv���H��I�F[�]�+���ſ���A����zRՙhK"��]�gIv^l��:���O[p�t4w?Cf��x�1B������||���4���m�s�P%_���:fD���;#y��-�F�����Lb3\U�7:�=.�.{P���6?-?18jx����gt�	dŒ�8� L�0�o�lQ~lOz�(PF3�i���N��Nj�`ToM�J@~��y�6{�uj}��3�����)��c�XSo���\g1�x5�xxx �q����Sa�^L �//�ke�;�u�tP���.BQ,u!8����{��i�o0E;7Q98�z�d�[vv�wڄ�����^l�f�J&��]ԭ{	�;S�yc9�N:Ͷw.r}��d�) �n�@��ʢ�m�ꋕ *�j�k%/���֜�<~�[;[nu�(���(Z��&��h�]�&�+��C���M����,
�E����{1��/$�bs�á{sD��������uN��v�л�j��o-5{|J=D4�c�����d�/��X+�t��;�� �����q�j��]m�#�b��J�;�͖o1]�"���mX͛|�����t�1�ν�ec3qCÅ���Ž��*���Y�;�}��h����aR�<�+*R;tF�c�B��$/C05��|���]g37x���#ܷh뵤/ge�[��X�=c�4���T�T'pS�d�	ք���s4�>��ͦ兵9dō�X�WW;mo�iU�8s[(:����f������s6�8�z��/*F�^wѕ��£��}�3�������(M��a�jv�=�k.,��IΤZ(�Js�%K�����E���焮�b�v8pF�E�0�F�6�	���c�PA�1�f�N��
��nc���fco,�E�M3P�y�gv����/HP&+m�Y���R��xѥ��^�ʑ2��M�W���Fgׇ��T"dIء,�S�]S�����U�V��M5��2D�u R��/�.RI�5Fr�����,����l�r�����#�`s:�r"_,������&�㦖�ȦpَL}�M���Ѿ�+�pk%������0y%�B�{XsZ�b����Oƨ�Ȗ����
��a���n��Vfc��T�H�;�X�
&]�T8u�)'0V�>���ƻ���s}�KGkCY)󓩮	�K�;��bY���Z�x_-(U[�w�.�b��t�(�3;l*��z+�G����X�3����s��fki#���.��)����GMuз	�zȉ�9��D���#�("��n\W3o��ƟWF]-w��)w�;����.�i����Jګi�`,/��Y5��K
���������d��ͭ쓏��CQ��GG�RiN��p�CW���4k��U�"��S�e:Q���B�1�(��1�δ��O�f���5���ь�����#YH��s��Wݐ�B禖�g���Zr�Of7an��)�l���7�C�y�w.�"����=l�]�m�F�^drWfl|���L�[:�$���`�kr�m%J0Q���GR�y���0(Kb��$�LûƁ0���P�Ӏ�N��XeIQF�%JIBLR�I���	�@�YpU�m��b7��Ke��J��Y�M�BH�m"d��>AE2�Z���N�,�K	�, �%1I�T�00�!���N4�R"[*������!�M�h��9�҂���5)��so8�;��*	lU�dH����-E�$��>C���y���8�k��m|k�k�kZֵ�cZ�_������{U���R�@��	�z���y�sLP�����H�		:��ǧ�___�kZ׍kZֽ5�kZ�뮺���]�dTK�THH"I��^S��DNi�B(JC��L}j	 �����^����ZּkZֵ�k�k���]}z�xN���\�'���9�2A=maKhTTDXXHP���D~��x�|}~>>���ֵ�ֵ�zkZ�Z����_^��@��&�cm���ɑ"��D!|�uu����$ ��HBPAa�iu2������Fؓ��Je���N�BS�L���'� ���A��z��MaQ�,�ӉrH�>&S��,��@��P<����*�Q,,���	H��"�K`U ��%�&�ifRu5"�$Z)<[�U���!�����zڑ�����H*U���k�FA0�jsh�-ƃ�$������ͤ�2��5�;Ȓ��ַ�-��n�:YA��.p����=���s[��&=N�p�n���J�XL�(��(�dq0� >F$���Ik�7p͚d�f�~���!<q�Ǐx�<q� uѽC�39y������)CA�P��06�%{����%�!���g�!�3Ռh��/�U�;��noT��IyV�x�r�-�W�L8?�dN���y����6��"?�[i���R�=���Ν0�a\�Z��u*��Ý}��̢��m,�X)�=���3�kj.=��Hʈ	�s�B��P��d�UxNo+[ڜ-t��bY�E;�rP2AF�޾q-ޔ�9���Ǜ�@59����zw/6L����
��4�2#Z�����/��<��ߢb��0���2LG��jӳ����`�g�Ϧڪ"۔@�V"=��'sN�c�uO^>+���7��h��r��}��y��\�e���?D?
������A-x�,���,�\����\�q����9���Eq��{Z������H0��3����Зn|��6[�)�C?����)4����^�+�6MF	p��5�!�WA6�te!�͢ޝ��3И`c>qb'���%����h�0fY%t�p���4
��|7�]���z
�޴`�h>x��]���@^����]zQ��w��o��C4<�XE\��#����=-E;�o*�K2=�C�z6����7]�6�{�n�J�fu�{��>�6!�!,Ҙ��_)��3z�z]�����oo �S('�g>����3�cڹ�s���wY�źw������ǃ<q�Ǐx�x�ǀd��u�xoT�gç���9��zG}	�|t�&p�������k��r���f��:�.���Ce/E�����5�/^s�1.7�{bt�ϼ��ijh�
���ü!�CvX�����7�Ra�$�ehaUz�q<����D�S��٫�=�݂M�����X�~���a��r�`!�-�~Š�--�����Uݐ��_���B�A��-L�#iA������c�������tXp�o`^�s,�=���ݎ��%>���涱���h���(�V$k@��o4�郢^D�K����������t��L��FBQk�ߙ������WT�Ewt���|�.�b��x w�Ä���8�Ny�o�H������xD���"9�9l�,�Z �����5e��z�u�BpĖN���l�l��7���hj��_�.��^1!���ߖ��I�����c s�F�n�nw�ę���ְ��«x�����:5�5��<�y������%~������5��!+r�6�ڜ$��=�E�#���f�Y׌kv�C�=-��h���/l�V\�hM�Y6I!Ԃ�ﳥ��:�d�#����R<�mgCv�_M5���S�z#������Yv6"�r��yu�y/y���&y��~���\xǏy<q�1��{�77��{�O{��
A�w�W���ь#�8|vA�^�%�N�;2���	���ܱ�h\�/�u�����}U38�5���'Ľ$�S�^�yj����csP�m��yGr��;�/��x6D��2J!�����M�<�3�X5Ls;F�/%�vf#'�r>�~�	�@�6��{���D���������D�����wy�����yw��V�7{��m$�d�A�!"?	�����oߝ�����/`T�����Lp0i�l�}l�y�ۚڱ�a�={��Rz��~)�����ң�ʄ��?f�M�w���\:�Ʌ���0ca��sw*Ƙ�������z��u�ع�MC�S���<�ݽ0vf���5�K{_�2��Fmgs��z���iqV�l�A�˻�r�"o�?؂7����➲2�i
r���f�[Á|-L�ǹ9#�ɮa���/�v�xR¿|A � ����E�ǚ��=�o��[�Kt������c@���r@~�x�N����fMz���UA����ޏ�Z�Z�#\��މ՜�n�}k��lv<ȶ��oh$���&�5bf-��vmT��s1��gҙ���E}�&3���҄�5� �T��8��7�,�h�"8�8U�}x9oh�ٷ�rH� �y�|���8�cǎ<��;;�����}���ӆ��_�8W��D ��D�S�}'�@L����5�
N�pu�����kM��U{��V���D��}�Ƙz�;O��~a�*5���=k�p��`p+��8wD����$�I�y��^�K�m(��ɑxo�ٯ9����'���ᱮ+ѩ�\*�\��8������[�[�4w�����R�p�=��{������Ib��~aY#=��|G�U�~�%v3�i�T�҈�մ�r�{i�r�M�5�L��:p$�e��[�^z��kd!�����#�狙fT�:��q��%���*��:\V(�z/���_�U8կm�6�L���o_-���Ń����s�"]�O���{Y�`���X�R�Mi2���S�aE�4�=�.I�~�������	�q�aq~4�Z�藗~XI�����V�6/�,q��𓏀���ܯh!���v<�yぁz�8p���%�s��o�Eg��p�F1�&����j�^5��An6�}����p?�{U�GfP%pB�|*r���~S�KP�����;s.��J��hm�֗�m���A�Txn����;�//U�	G�,�KE�N�4�z�q�g&����LBO�aDI� K��(�>�!TIi�Qč��w7��p_>�^��釛��(��_E7{^�/:�^��˅��Ņ�N�x�hJ��L� -ĐQ�J�d2''$ɓt��7�����\xG�xG�<������W�v��߳��i�C�^���3���	�Ŏ�C���)�FL!���TO'��H�ۋ�FWoW���H���1�=�����[	�[�������{d]����J4�6��Uډ�]L���1ۏw$��G4V�8䫑��c׭����VV�=�{{�9�`Y�-A�S<;=�w�m4w�^�����z E��='|}4���O�Ҙ+�+��⛋�j_�"��훡��o'ꪃ��h`q�����؏O����T��arUW�J�{[xZ��&İ�w�Ox���1/���^c>?JxM���Z�+�*삅^m��nXu�0c�u��:�7��t3b��à7�א��"7F==�N�H�'��<`��댧)���Y.�G�}d�����<��0h�-��2���o��Z�)�F9��Kq6�D�����~[B<?�KM��U�{���j��WH%��~i	��m�fy�#
[�>��L�5Wy߷�#?���o�uH!�=��w1"W�U���[}U?rƮZ��t�J�_�����9�������A�6n��@s�ǋg��*+�H�k)������,�w��;���H�D��oL��^O� �utr̈`oy�8u_pBt/gi��C�E�u�y��)2~~8�q�<q�x�Ǆx�Ǌ�{��Y��Lx����8���pd�������F;U���N���Y�V��_����(x������E�T8Zc��3q~g�>*+���^�۟&��O��l�z^���7��n��.B��y�#M
N����!�W��3B�ǉ�d~�2���,!7uJ������n���=tη���{���Ж9`>c;��'��~���p�}�oo�<�[��;x�^��:�D�"�~c�Б٤�_6�xi��L�/��뻳{G^y�!�8,��g|Ǚ���>��Š�����wHU�o�hn�Z��Ӂ�]�;�)3M�m������~��N����'r���a��zu�V>{�1��Hȱ2���j;c3U����i�v(~��`B���O�@Q�X]����'2[m5�w	������Wk�����v�q��孝�Sۼ
{������i`�өm��W��7k���y����r~]±Rknw��=���x)��w����W=�*r��#3�wk�d�b��Ok��9.^��qD򹅀�w��Ay��oq����䭂�P��~��Kd�O����3"Y�Jj�i�. �l�m�]�3��-���*�u�W��)�Y&��Й�=~�/3���?��<�?�l�Y˺O@o��@0��R���6�R[܌Y}v���a�X�}|�}U�RZ/����B	�	z@C6Y�3ty���чX���P3Q�g�6��e���tSq���%�3���9aC�M��,�g��ޡ�t��Lh��/Z�ss �l{cM�g�kym檾�q�/ލ����X_/����_���d��������>��)M�*tK	4VE�?f��.6+�2t���Jd�H�س����f���@W���j?/��{�Y�����{�k%����5��I�y��1����|Zu����FT�Xo�Ip��)���sH���R1v���59��E�VI��bXHǯ7�4Y�
�C�� ��F���.n���u!h0s\���5��k{�gH��C��fM�츟O��,ZZ��[�V�l�J��Ӹ��.���G�C��e\p	���ۻ_� 8yt]��|81[�u�=o�-����v�U��%{����
z���	��|��!0��d<?�\��ޡr���
׆�yq4U;S\�Y9��I�!���RM�_]�'>5V8�ِ�B���k�`�/D�n�����(Є�;L2�l@$9��!!�$�I� p48�SƴWD1M�tg��<o��a�ݏ�{�N�gY�:v^mM ��p���=�m!��ĸ���'��>O�||�q������y�5����&{Rp���=�QFi�~r,��9�����ź��� ��qM�薀ۆ��Yw���#�� �O�P%�m��G�-�)��b��
t>M���l�uߪ��s!*�n��^��Ц$��qsl��6Y`4E�����������Εt�{k�H�)��-�O�"�)�륨��!ޓǭ��[��0�o���T!Os�����������F������ݡ�]ا��?�CH��s^Ϝ{d���w�)P*(�0*S��ͽ*���G[���/���� *���C��~^��krr�5ϩ����QU�܅���EY+�pցG���r��N�7��ý4`9r1�C��Dq�*�y�\f�g��~��ֳ��nU^���D�nxa����q�8��C�ߥOoy�	2O��|9�I��ё����q;��%���`K� �Z|?5�L�I=_�Q~�����,pͪ�
��H�P,��zy�\[G��r+�����Gs�}צ���;�5�:ū|�D@a~�]�c6F.r*���:C8gʺ���c9�hoe��K�(�N�6VU�ٽӳ��յz�P����.��v�lu��)D���>���+r3n��� H$�k�3Ʒ� ho&��.��E�s@YJ�8E�(c��=[�RaN�M��ڷq�Ցe+��E�P��1��q���iJu�4�j܊&bn0�%�1�����^^^g���yyyy�͟w�g����M�@Cy"K!��w���H}h��o>�fW&�Ro՝e�1T6V�P��/1j6��#5�g�~95�����*3��#�G���Z'��hW�P1���0j`�����we��dVar:F7������x�ƴJ��=g~�TVoŔ}L���
��U5N����VS�t������N�3�ha�U�g�<׉9����
i�f�yީ�ޘ��
�%-��&�$��Zs�/:y���g�����0N���X ��lF%;zC��)D�M�،�5����Ǐ��^��F�aX��S:\���:u����lr�[r���^�˪�τ@���9<��FQu���n�nˈ��.Xw��1`����L�Ks	�WW�����|m���4�ZzK�,��kJ�f=���O�3�ߵ����Ѷ�3�U�����y�o����*�?+�]�ėX�Щ�?�;���ڢ����N*�m��)�]<��QT���C�6Q �}a��Cl_��5t�����|ё7��ۤ�3���������U���>$gc��ֽ;"���Pҥ/���!nެ� p�/~�,O�H�}lB̹~6芬�f�6���zz ;��N��t�=��" wc�kg\|�_
858�5�X1f;Y��2菽��/�����������=����}���~ Ȅ�����1�eX���h(X�y�3?��[��E�=oF�go;L�&���5I�O�"�
z/\��8��8�B�&��)���4��7�k]��Q�h�W�V��l��&<��R��E��0ƾq3�տ7u�|�1o��z��0����_kUI{�����d�'���ޤ��)�L�n��,':9�k�?'T�697*���g^#Y7��<
I~٤W A9���$
$�0n��j�oK���&F�7��F��fi�{kz���q����Ưw\�/A�͵�Ѱ��^�m���i{>W�_��w�yѽ6��?����7!��"&�B�+�n.��Z��v���`A��4�\o��E��U��.'8A��6:�՝��~@�o[��M7��^ƍ`��3�yBӻy�ӡ�,ldS<p���i�ǆr���K��7�g�؅ݪ���w]����3�>7`��y [i�Ϊ����X$����B7�N��@|�q������~��CD���͏��oEW�&�L�ø��ع8����e�����������}�m�ҶvI�_K9;|g���GSV�љ�VZ̩Ч�8��);ŕ(�w���!ڎR2W"��ͬlvSz�%M�zx6漨̣�-�j��uq�NU������>N!���y{�0_�&w��9�[��*��w:ujvH��c�C�=�����ëj�:��������Vq7�%e�-f��Q86���W,��H�NجjfXv#��s�q��S�m�],�
/kN:��r5rmڨ�v�*���eLY�a����Φ�0���tɴT�R��]JFn�.���i�.P�����3S3���e���{}��gו�T
�1�Cfl'�,�9�w�)���.x�>}ae#LE|Eu[wt@OJ�pi��.R}Y�Is�sZ�IlB떯chi�R�!��.�l��,�)���J������Ƞ���&GohcC��k���k�Wg2@\��Ž׫���[�]n�����<�ơ
*�ps�ۮ�+������+��y׭��T�r�^�-�,�N��c�Eڳ���[y��]������"d��V_o4��73�~n��g|HT�>�U��l8�_���{�S����s|L	��U��U��S���D�msC�a�S�%�A'16�/0N��>�q%�ᢺ�b6��
	3��L���aBZZ`Ãx��HqE�A}����.�q�v��b��:�;ʯP��w$5�����k���ܭs,\���r�p�8��É}Z��i��4cٓ��>���� K�l�N��k.�]�f������v@h�ԡo��6�r(]fVK�%�Y�t�����8�5k��1�(������<�Nf�3��d�JI2�	,�$�&���2�v�]��\����<���������^����1�F�_]B#\8MZx�Zw-��Ix��ru���	co��R��+އ�i���6om��Ӷ�l��fխ�����'k��t��q/\Į:&��Vl�yr఑�W\48��榟���>�{����ɱ��n�o\�5ax�hJ����e-��(0�4�G�*bg��_E�
�ٸ���z��K��Ta�Ɋ�wX��n!�/Ϳ\�]
aP�e�ps/�_jH�QRux�R�T��;׃tj�|�Q��>yؚY��:�}����F��^�LJ�xv�j�7D7pY�_9�	�a"y�T"�[.I�=i&H��Q@$*
Y	��ח�׷�����kZ�kZצ��6�����oo��{�_����h�6�W��V,)a	�
�!y�D)
�����ח��������kZ�kZצ��5�{{^�����
�D��.��$	���*>2Z�"*ER�ۯ/o���־��ֵ�u�kZ�kZ�Z믮����!p��d X	�D)P��*�'6̋�`�!�2x��k�k�kZ�Zֵ�Ƶ�x�]}~;_�-�V���|\,�h��P��(B�,����B�^�	iI
G4�/v�D�!�i'S!(BBBC�x�^ĈBm�!!j�A"8�aJIK�$�"-��� $D��0���ؓsY�ų$����TXKĳ�B���"'��%�"&j��L�܄R"�t���g�$�IHu�,!H�����I��K	<L��O�9"��>�ܒ�B;��<I$��=�wrP�������Ge�]�ʏ3�(�M�N��������jH�c쥆�!]�����{��|G�����z=q������򸮫�I�-�����C&�Ɋ�3�A�����Y#��"�`����V	M]���h���zl}��^@����F}��X@�I-���7�{�NA ���j��Z�_���l��ua���Ų݂|��U
Ƀ�>bÿ-(��'�~a�O�.���sa[Y�;8P/m�>�Ť�~��W��_��6�%�ַy��r�D�3�mn:S�w_~�����H|S,�����G�NCE�`���1tq�B�w�]��sz}��ӵ��`�E���p0���xV�k��}q���x�Ը,7U�+�n�����������[9�*<�Q���7_S�ll�螽Oso�Z2�s{L��J����.!��ms�\c�5�u�\齻w���عv��l�%��b���C{�޿}kH�X@�!~w����|� &�4�T��[��Qi�~!=ŧ8�~VU�OI�-Pf`sXN�x�l[&���<�Y�+�c��mGb<�v���{�6���(afZ�*�u"Fo��_��; ٰ��0F*$A���X�Wl]���fiQg��t�-\�nm̾���(5[m���oqZ}��2�������nڱ@��>�/yyy///|ޏG��57�M�1��t���(����?��RK՞�i�� �DS�O��ź7x�������J�0ҳc	��`t\���F,�nL=	x�nO�}}�;�M��28�d@�QGE=�0�g��8_3�ni�U�5��dU����7���)�ël�(�n\�x��@5&�g�o��l�N8� ��NGm�nJ'�UqB��b���x�g�>����*��_���X����yn��Hl0@sę��زi�u3��(�T���f{dv	tM��1H"�m��/DѨ��Q�#U~/騊b�f$�C��ח�j������}���y�WP�I�[�P{�zR��j�|��b�I��>1��-�#`O�Xt+`P�����O�P�\o��hE��9w��Ķ�ay�d�S������<]	?N�{��^����Uγc^�C�ni��%nCk�塲��vj�3��E��f+�ʒ�lz%i�|�Z��Y��:�iS�r����B e�!q_6��5�g��ک�}g�	V��i%݋�v`�ŕ����}���5$�W��vs��干\Y��j�2�𠪥]1D�F�qF�>&��e#uLS�zpq�pq�N��u�7vL�}��y�Ӡ��f��i�`���Y���g#�С8`�F |�`�@(Dx<��S��N�q5R�n�y+:�=Њ�&9��;�د�yMyς�{0Z��&���W�3s5I&q�d^B���|�-�
��e�'��X�&Rʖ~�Y�l7����vwf~��P�}Q�=ӹ����1Μ8�=o̞�=�̉˲V�3���9�R���N�u�v2��]����s�qf��2`�ӶR�]�����Y�K��F^�3��3��|Lo��:ؘ�|ά�J��P:1�>���"z�0��
��1�'���.����l��n�_a8L��s;��p8Ʃ���>�-����e�\�gc{���:��9u��u �eG8�`�����损u������y{&�N��0ƥ�"���gΑ}�,7����qb=E�l-/���U8���B��q ?��ȹ5�V��0=_�?~��j��b�e˺�]��;������=wRܬ���@�[N���ǈ�ywJf��{�Lɜݜ�x���*n�9Ǔ�t�v�/�އ�KBu̽�';���#ǎ8��<�m�߾��ߡ�n���!]{���-�qU�=:���xع�ƱLb�Z�W{J��9ж����
��r�{��[_�܊����G5R4�o�����Ƌ��m1�4� �#�޶�|���7}Swx�U9�7-Gc�k 7�L��I/u��!e>N�p��T�m��#��F>��I֤�ja����_�y
����9RO������)�ьyk>�]�l�vgY'���v���n�@R�r�Oͽ���y�gw|��85˹������B�ܝ�²)�X�!����(����u��_�k�Xb[�T��;������-טz��zKv�V�w�u�>�`}�;�����6��34M��S�,7��n6y�-͗�K]i�[��^oƶ�}>�q� ���2n\��~���M�d�[j�b���G�:x�om�#t�{Dy�,���f�J��P[�K��X��kq�b��
�[�f.c �B�H8n�Ѧ��;����e��ׄ�كxS�7����w�Hљ2	P�Z<3V����x��8����%P�gAj���:�U�΃�M=U޿o�y��q�����z=ڼ�K�7:����``c�	|mDC�3�{g{�d6c��t�����`3���S��tPD�lؿ1�ֶ�Qq�B*�+���d���%��1���eIx��9��fq��v���{NN�2�0��i󸱯�}��{�N^�@~�z(邛ڰ�OuLh�n����?��::V,X�#W��R�j}�����s�퇪��������W5�:���;tuJ�f��}�����S�k��SC8ec�{$A�����!�9��e휜�8C�ؿ-��3�g�v��\�z_�yrݵ�މ��"�������RL�'w��w���
w��ѳOI�����n��M՟ne]oN�W�++[}~"_�ߵ#�O�c0a���]I��)�#��e�~����{�3�����n^��//�!kh� �U�'hY������ɫ�R�x�{�jڧ���t���wh�t�ε����\T�K[�U��k8ط�,�N���$;%�J�k�9b�m�������n��4�睆��JR�jl����&9�״���<�r��e��g7��냎88ノ8����ߞo�߿z��Ͻj~#l5>�3�<B@����;\�=��T4�3כ�w��n7�����ϖ���an;=ŝs�ٲ�o�-����N�7��<�c� �,�h�O����
�J��:<���,a1��'6`F`S�s��ngno-�t�0����_�n�IݿU��¼��Zrz���y�8��9�w7Wլ {�u�wԺ���*:U�W���'k6]�{�[6�6�pg�\(�(�![Z�S�?��A�lw��}�p��M���o���m�N��h����Ik���?^��֥w�䯐�%���M[Z�ꩧ�7�wJ�TJ^���vW������B`վ�O�޶����vH���BWB�t��XY��o���n�xI9���� O����E��J��Pz ���9^�1ެ�C}Ѿݢw�}�V�Mc�"����G;�d�I�u��¶�3�x�����U�aҤ���8����^\n����d��A z����S��O����e�YX��E�XCy��r��Xo��h�ۨ�u\����vB�NL}�zk�T�n[/��>F�F�B�S$a#2Ì�����nO���K@DLq��9'!��s�����q��3pe������߻�hd �E�-�w��p..��.|����~�پ�PQ�n�1/�;�]!�%��F��Z@]��ez9`�P��`�a!�*؉�'Y�Z��g *�Χ�}�CO��{~��&����|s|�FE��Q�!$�ei+����K�?Yk��d36�t-uz{�����\Jwo��W������m^�P��F̆���X�6�αf.*��j��γ�w�ϝ�Ol*�l������wE��������d1���~��ZO!	=����ñR�w��]0fmR�R=,=����������0�7=�9�!����^�|:�/�/��ճ��V"���QO_���6*.�fgw�;J�`�lЫ����^��	���>{����R�U�}g���`��Y�pm�(+^�N���ȿp�g<!� w��q�
��8�xaB�e�HD�IiW���X��o.�)a�b��a*a�aV#��c�}��R��E��C�kއ�K�0��<,� i�b���n�p|:uت�A�8l}�����q3��o ]����M�7� eg<�iӟ]i'��>�5��q��9�W�=��.̯��RK��1�����{���L<u*���g�ͣ��75}�tw-gi�B�衾(��T&"���A��KK؞އ�*��H��"w�MV�N�}�0� ^�� $��1��5犭��
���ľ^ҋ���O�"�5�ǧO2�Q�w����ɼ�_n,�w�s"qJ�f�Ε�|]�Ā��2���Qn��I�0h�=3�#�Y�P�4�ًN��Ϋ��~��3��싰��zz��Oe��hl<Q���L��}/2e��v+�
�&�C�S����[��#���?��,(D'������ǿu֐�xS�Xd�qEa����Œy����d$|��������8y�����X�Kb�z���4W��W��t���[E�k���gF��-Ts�P`���m�:�0�٭5ڏ�]���,�5����>�J��{���{�������*���gvT�U��Bܖ2L:�d�M�#`��Z��ܖ%nl��Ĭh����[�yr��A3M��vE�:�S�#k4s�};o�,ͷah�v x'%|���έ��a��Ž�;�c��+#��W����<��8��?��ן{����u�Ͼ<{<���Ǉ��7v���'ja�Ԗ�>�P�9Z�w�V���q�γ����t~s\�͖� fws�w��������]�+mn�X��2�f_�9��*�8>��~a��W@ɷ��Z�+a�"�9�O#���%P�N_��J����A���0C���۱�FC��A�t+&�=���"��(����������a�"v�*<dA��Q#��j0�tҧ�g�v���t{򧒽��a8��^�0%�4%���D;�N{z�К��@�S7S�N�e�g���~�^�Sr�!���qu��|89�3U�g�Y���!J��q�ݬ'���T�/���@���̞&5�嗕�Q3���W�����L����g�MW�"�o9����L�-�;�����~�??RUy<��Ӷ�9o�̓����������˲V��A�g��l7�����b�~��C7I�Op�n��xr�T:����:YΤ���|���d����(B+^��;�޵���=k���^El��`�A!�D���KY�1ܢ�њ�-�8PJ#��;���v9���F��.�7v�l�Z���N96﹙�N8��8���^y�~���Û����B�N��ӧ��(�ۃ��s�z�K�r�(���Ҋ9qEtF��s��t��o����s���ʀm�Dv�~y�!�,�y���=��5�11����>o+�z��Ӕ���h{����	�?��]�wKam����V��y�~q�Yv^b�Có�fJ�I��dv���u�3ýO�����iVM�	�}Nj��)���<C�O�'k�WT�i��UY�Fϲt�`Ҍ@k#�<�.�mt9�<��{��VS��V�aԩ{:x,��V�9�i�VFש��~h	��F�� ����ZF�I�pF�!��o�indf�@�P1��6<�;�׬�;�HZ!���q��TG����6B�m�'c�#�
y�0 )�<�O����Gq�w0��>kO��~��= [���U>��kG�a�
u[�E�t���1Կ��;�se��Sy2r�y6�.�c])Bŷǵ��}�:H�\��˚/rv._p�p�z*v�k�=�p;�!�m;G-;�l$���X̾���>�&'n/ek9�Zn�;tt�Ӳ��r�U��uF�F��n̻l$��3������ڭ�ҩ�H��T���F=�c"���oQ5G�Vᚩ�O����J
W�'Y�?hn¬�V�������7�
z���9���K���Rۀ3����VY��hq�nP&���+�C,����N��}��hֲ��:���}e��<���Md/���\�I�nu�;	��s"�+�-Bc�)]�/�����U���1����Ѕuڤ�n�-�=hc�d�\�%��i"���:�b���Z�wnÇ;���U�p��}ƕ��M��Fa��]��,@ʶ�Zި��Z���\9�p
�ǝ��L��q\�r$ç3��{3.�� u�������yr>ك���3�"��1I���2<��Q�z�w;���^�%5{�V�c�����V���η:_�3��r%��XH�ފX�A�\�'�-�%E�]���\vJ�ƕ�,��%�bQ^&x�����x��.�uj�f��,$U6n�ddLU)�a7|]�F�6��Jl���\.qN{��$�m�92z:�\g B�*Ԏn?QnƘ�|����fR�Z,v�ذ��`�������xI�0d;1��)"��Z���-�;\������1w�m��M��H̵u������w݈����ӓ�@w$��ຽ�u;�¥�̕ӽ��ژ-�%G���*e�ckq���i�K̂^��}s���+3l�2�N���Gk�לm��P������UM޽哛��P��8��%D������nYDU��q;��z�r���3����f�"�M{md깚1�n֎c�앨h��s��pR�l�U�|l���}Ro@�d�Xn��T'=ą��vi�[/��=�s3���A����ȷ��ھx�ұV��.au��M7�N���v��5՘!W�^8��	�D��G���^�a�k���t�mk���.��ڻ'U�X�[��t*��h�]c��亼^ҏ���.qA�i	�&	opN%�	v�_t�7��R��*=6�^th��VZ��̸�w�n�m���g.��Y�9�e��+4�Gq�23[�R:�*��Ѡ{I�������bI�gu�5��;e^e`{�l���U�/��I	j�Ք"��;4Q�˰ږ��$�T�F��8+hU�v܁T��?@�adm(��*&*�B��R �Jc.Ġ�.WiƂU�"+)2�(wP��cr���p�M�{Xg-���nv��F���lrU��w#/U�"�8�9@�(�U�[e�C@�h���A!JFkL4A �
hT�#p��?5L�/������v�	�h��	=�"���ק=>>��5���Zֵֵ�k�k^5�]}u��,��*/�˥�ie/���L!�$�'�W�ǎ�>��>>��kZֵֺ�~5�kƺ믮��� JZY>4"UH���OVi�EHXJH�H@�Ʉ=���Ƶ�Mk�Ƶ�k�kZ��Zּk�������M��QlD��aa�J ��L��f�H"�T$�HC��>����>���kZֵ�ֵ���kƺ믮�����0
�H��D|MEDB}h� �ܨE!Q#��a͡ ����"ڈDm`Z��V�� �\��&�>���'�A�"ԋI,��$-B"%
RBJD �Oˢ!=,�wbT��$!'ķ!j���j����� ���Br%ȪB)lD��q��������E�&��D�Q*��Ҁ��n$À�B%�$A���P`�к�;u͕�4�4�usy�rbfgaw�Z�D!�v�N
9l{�67�T��V�"��BCFl0ɂH�`1�!�Ɣ`�Z7�����^^C���yyy{�,a�E��wR�����ߋOG*�I��X�{l�??o�Zҟߺ�_m��e6@�d��K�Y�����,t�ˋ~��|GĢ������MK�el���x%�sQ��ړ,ޜe�<(�L+��[��]���ʽ0wg-�(���+A��Ow���M��<�M�l�R7hώ�����k' ^T?V�ى���G�
Z(þA��>�"���+j�Z���E�]V*��8w5��ﻺg��s��)�ۖ齔��)�f7CJȥ:�;W�M������Pgw�a�yxϟ��M�Nz�2"�m�vwr�a�np�;'9���U:�
=Y�1�H�f�`���nm����K0a���>0sh�R��6[��lvWC�\=������b���ޥ���t�[37O__� �h�!:w�qu��k�N.ݐ�g$��,��MĹ����u�fe_�;+>���!�K���QT�e�� ��P�H;͏Y�4�������Wq��-nA�٤V��V��a��sP{.���p-���ٛ���p�t�����C���yyyǟ�����]�IW�&Է�����WG�H��"����e^�iM2L��c�f�M���.`1f�t��������F�J�N�a��t��[�F���V�S���`Q�����8$7q���ޥ�:���!�P`�fgV\���Gc��5r�Ϛ@��|8��2�tP������W�	�>�
\���ߠf���$�[K��ѡ�?R=[V;��M��e�ì�����Cf��m��:��7���C��>ƍ�Ҁ�/an����o��?^���Hw��ba� p��u�W�dJ_�~�x���`��5�,l7����@Tv��3M��v��yZs,��H��Eyw�Ϙ�5R�=2�.��� �#=ij��/t&\�|���[˲��U7FK|*h�K	^��|�a��eR�<=�`�l�n�4N_
*��Ϯ��?S��U���X�1�:���Ν���S���W#op0d�:�ݤsي�gK�������tN��+JBm�줖�M
��%y]\�����3�q}�0s���N���>gru��)������ģ��e�w:w�y8��|��śN��q�1�q�y�g߾}�߾gȴ��w��S���첿M4=���酐#������ܑlf�I�� כ����t�.��>K��[�O[���*��qm,,D쩬����a�L��G*$��aܺ���ot��d��)�)>	���|k��Z��%���k	[�\���szvVujN��}w�W�v���=P���ә��f�.�$�E���h�����͙r���WG����.Y���,�JRVLZ���-�N�xk��p��&�ڤ&z��}�<,
�FXioe�uc�i�����7�3y=y�!g�Ж���,4Z'Dw�l�f�'iy���}m�����x*�ѥ�l��=���� [^�9|N�����	�������q��~��X��{��q��ɋ����v�!�����dTbn��3؉"5��'�����.���ga3VŊ�;�[��I�A0��ܶp�-9�����p[�R�]0o�?�grD�5|ޱ+���v�[����!4o� �mr�����L�"ƞ<��T7�٬t��]��Hi7��L�_';�I��8��8�����N����7�:�Tsi�?����i��D�yT�!�žt�`���Z�K�!��~�>g�b��U�ި؉�K����/��2r���;��f��e�D��u�"�5������e�U{[pr�̙�owg�+jq�V��;����u�wvp�&�^��}�pR$��s����Ƞ�*��-�T�B�8a��T
�ia��#�l��\�`;w:�o?�u\9g������;�Hund�q%�;�;����#ռr���������m����s��f��N�����G�5׺����a9�E4����j��ǜ�^3�
SQ9x���uwz}�d>݄�j'���C�d�Um�6�sY�3�n��\]���[*Pc���$��~f�P=�7�b�z�g�'jl��+���鳹^��r��n���솰u���m��s�.:�M8N&��4k؜�����)P�p�	�͇ 겉��E��7N^֥]�G�{�^N�ꦧ��F��餚Db�Uۀ�hT�4E�@���U�=�u��Ijիy9����4k��W@�]�;���*�f>7��g�N}u�R�#.��훅(D(�)N���
P0َa�U-1"a\�m�s�6;���w�{u�뮗]t�����eE�쯻3����Za��37�Z���{��-uO�ُM�&S�T��͚5f�|k�Ll�|�2�,��oau����
�u�{(��~𺀏�O�(��8������8�Ѷ*�g�R���п(��8WV����pg�_qOɿ�4oU�oW�r�/E�O0P���a3��guY����eB�#����a�F�TH�_u��"��@���C'��:���Mݺ\\v�ܔ+�
��&��.�y�����TlǛ��T�5r�nǴ�Vj6�:��9;���k�`�x-�U�-#�S�-����ކ��S���g��S�v��ݘ�n���nvT���_�yw�3�t����g���a?h (�ߎU�0P�Ϗ}l}!_w`o3����G�,37uvi��<y}�v}�����������t�K7+���6y�8��έ�oѿm��=ͥ�Q5@�Ywc$,��m�P�떱�����Ԛh-y�D}�7�תTD���u�mw]�W^��Ӹ��w�k�g�Z�fus�y���N�����\'�]�,t캑�a
Ty=88ノ88����/_|����s�̷�^��[���:�g�e��r!��x��=ӷ{�Ŗ���;�q��^��Θ;}1\�*Y-�����pW��O��z1�V%�w��\�~|�ڠ�W0�1�	��譸fwv����"�$�y�wyj8.�C
&7��p���%^�1�~�㭩d��y�Q��|{m
��"d�  ����̂�I���O/��:���x��f&s:ɭ�~i���s���\����owW�_%_s�?9n
2���N����vw�⼚����=���s�B�g
q�H
o�T�<����w�5�q�kgC����7��gV��2��I��K33�8-���tS	���$����l>`� �����CUp��4��Sr5��Q��}9�^�;@�k����7�S�"ԭ���e�K��L�4ɷ6�C�WS
�׶a�qgh�����V����x�w�+������?)fxq���YT�G���}�g�7��p�τ�2g�F���\����7���I�n�:��:�Gͮp�C��W`��|~>x?���?���V$�.�~B��� MO�r��Ǖ��y��z�]�����+��f��u���r���C����ڪ�^e�r� h�W�կg�gǉ��'�r4��Z�g�f`�p,r�"�T���4&���(�}���ZpWgbF|�_z�q��Y�~�W��Ά�&fj��g���ChUl�3S��z�}ߖ�N���Tf��*����:�����9�[`Z�h�4�	��W�fM��s�yԘ)Bx��N�5�c�W�����Yo>�x�ezݸ����ZhT���1��k��KǖyHػ�d���nf����N�І��v�'��\8~����/=�ϯ�T�<�d
�W�9��Y�3lU��4=v��;ט��]1������"=O*<��1����A+��3���]�<==X�b�[�U�e_B�z�v>�~��e���w�r�+j��{Uz53{cPͶ�t:�N �LМ"UL�ӛ������4��H3����Yo��vȅ'���@=BQ��k��uH��Y���d���֯��yz-��-�&g\�M��mh������8��q���ǟ�����J��I���O�5M߲�N��7'�<t��;�cVn��i�����ݚ�7p�U��Xɷ��W�{�/u �;C��S�8�.�b�j&�m����V��n�[�����a-�^ v��^�JZwYT�XA�+���!�#0>0�ajw����F<׏�.Mə�r����3�.Y�	�I��
RO�����x�`��7�ymB���TM�(8|a��|�~�caz|���cܵ�-�����dG��Y��ss�[0�Cn�tz��͠K-�����!���yo���e_5�ub�53����cM�}ff�4����Y���w�sb� ��dͳ�y4sZnoO"F���Cz�n "��;�"��{��7�5:�]3[w��Q����˷���0�<�65�Lg@�4���fCW7�_v�wT3��Oq��8����L�{Q�i˝\a۵��PrQ�Ժy���'r��"��ڴ�<�I.�Z�pi��F���X� J�с�r�$U�M2�M�aH�M���ר��M�ܮy�'�d�R�z�D'/m��z'Z�;bz��Y݇�-��a���*�tL��jeA��DB$F[p0����0���RC�R)�MD����C���yyy///�̆G
���y��\��03�&�G��3�}7}����2�x���q��x�3��".,3]�df��Y���f++�*X�nu�O���B���b��s	��K�vw���3�1Z�	#i�u|��z<���cy�Iy��'��8n�5���;�Hvi�̍&�9>�qm����>�ŷwGv�v���hM�������)2W3?6��Ɏ���ހM4zt����������Jd
�`7]��=����,΢����0l��͋#��S�����U֢�ΆQDd���]P6��^�~h���}�rs�÷%��k�#8��r��חyOm��1�<�v�y�}	�=֟\��y�5�ۯp����VC^�e���{Ӓ�fC̼�vcH*�ΰ����%�0c��~؟h�\�=�TR}wf��Ϧ���a[�}�N�q�|<}��i6�ͫ0h`�Pn3 ^�GWOp�~������TչY+��Z�[5��_��r�g�M���sW�ћ�jeA{uJ�.�	��f}�/i��/f6���&�L�1�Cq4n93����T�ֻ��^'��M"�>��
N�J\�m7aR�\�r�ǚ�[���Z���v�\���bl�|���o�u�Η��ξL�3��9����8��<pq�0:t����|&��h���7�(�{���2��p1]����"(�LwU�/����{S>�x'4߉��;soK|���f��`�������M^u^�*m���,��`Oe��b�y��&&a��4Q;B�{�%��ڷ��፽�ۥ�>�!Y���xj�d򲞡���ΪU��Y�D�)O��cs�������s"E�*Y���ۂm�φ,Mn:8�)�w���X�n�c!zۏ@;*RH�����G��v2��J�����H�`V�RI�� ���f ��XG:9����叞�}O�'˯��w!'���E0���kj��y`��{(?y��uW�E�(��{��<J��GG+��f#<+:��9[���Y�tjdʈ&=\bs���%��c�-�T#2�o;,��B�ye4�L��>�� �G���n�`����^7�>���X!>M��{M���u��Z�J�Kضe	EKҔ�;
���͎�v.�X�ܹ���M�51fZ�	��w�`I�;\�]��}�t�3-��F������z�;]j-WW]���ٶ$���*��:���m��ۦ�N9�R�pe�(�,�1r��:'��W��]�3���ƒm�ff�ө�`��vvu�E��.@Ck{J}�xqD�щ�Mmu/�_������mk�F�З]#���W�cĔ������C{�r�;�݊�k�m��se�U8���+���(�Z��V"w���I��(��tW���-�WM.����r�����VV���r��"�,Gx�P�Ȃ�ե�r��O�og �/)��m�YiZ���SD��oyP�zfk��Z�r률X=�gܑ֝)q:-o>]1�7U"�7��M�wu�mn7��}P��a��%Ά��{�L�׺����9eR��/QTՄ�s6�b�t�~��҂�Ǔ�¯+3����-�㏅P���yG�H�4��
�7��%�Yg:��RJު�T�H��h�ZtQKy�wMȞ���vR���Y�r�,H�D�@�Y�,6�g�(oo~F%|����@d*N��|/�A���P�c���WT���1G���ȷ��	�=��>�H5M{L⧓n
PРD�LS&^�K��2?�/W��ަ��N�����@�U�E�����΅f�-ㅻ�6	yǭ��j,ף�e�G��}r�����q��We�뭹r����;�*��h��O����zˮ�t�=��B�bKnZ",��Oi-��ֶŵ�"ӵ6�.�f*����jm�NdD¬�7X=9��5�sl��1Y	�F�]=F	Չ��i��Zx� ���*�i��5f��ۺq�BtWq9��D������e�w4;z��J�K����୆^N��b"��;ҹ�).��D�n�L�]w�6�S��Ji��e���a L/Mj�IL��{+v�v�US�rة q�[L�[��J�陝�KGG��&�ԴH���.�D�lf�̚�ോ"�#q�n{#�L��Ҟ��*<��*T\ s��OJ}��;���b���[[ɫ]����Qnƛ��V�A��T��~������G�*A�-�Q?�V}�j?�m��Պ��Z�Fﵴ�o7KW���ة�Ͱ���a�� ��F>[ֺ�n��rv�[��饺�ps�K=��^���1��gn!{c�dN#��%�̐��ɥ�"�$�,"Z���۫��^�ߗݯM}}xֵ�k�k]kZ׍u�^>����D�`�A�E��c�Wi�%Z�HFi2d!C0�;x��Z��׷��ֵ�~5�k�kZ�]u�__^�˒�$��zg����L���ԜL�����DOw������Z���ֵ�~5�k�kZ������������m2*�������':U�$�B9�ɤHL�7$=���u�����5�kZ�kZ�Zֵ��뮾����""Vj !��B�&$~eXH!k�rvKc��%$y��
�:��h�]��E,9-�d		 W�i�0)��i8�r�cR���̳�jZZ����g��&"O�i ��b! v�/��&�B
"/SE�����DI	�fXYX��:�D".O'yȞife�,@���$	@D����v�γˢ;���ls;a��>��I�Ɏ�$�l���Y�񾋰�SqoG�d�|>ノ88���8�����~���;��O�9 ml{=>'��#x�����۷g�M^:��`a�����M��F���%r��f����%J��
��9�wC��x!����\/<��.�# j�����Ѕ�M�dΆ�����[�$ �Ρ���4�ߵ�T� ���ܥz�7G�Y]3���K�)���e5���ц��^�&��^0qS�9�-鱞��1��a����[��͵yʲ�ym�x�z�tOE�p�*	Ļ�������F}�O-���l�&��5%^e���e �!@M�@��ie1�YL���[�D���1�2=9�OV-��nV�!���r}� ̇�يf�#zf�L%�]�]ǀ[t�a5�\*�s$�>Ͱ`�Y��6´���籱\�y�IˈQS����~��׫�g�p�]^�rA���D�jn��/�����J�v��WW���;J�[RWu޼a�w�¨&WUH�Ү��C�C���ݘ�7{dV�n������V��]+��9�z�l*�;����1���WW(��:��圳��h]�x��E$�=��/3����ǎ8���S>{�~y������ι��N������޸�%��y� �仼Iy0��͌;{�j����گp�C3@�u�-(N��������r ����&j�������[N6�Q8�\�⟻��X�k�\����F��y}�g�n
7 >7N,���t�,5�����tL�z1���`0���<�9�,#+�����r���\x�j�ZOWJ�ª�/�|����
�YxΚ����#z9��Q�ev�X�&ݽ�F�(�8�ڭ�<խ�NqE���v�����jrC���1���;����"^]�8�14t���^:��<��S�w�!�l��)a���.��#9;^֍��}���!�w d�,��v��x��2�Z�,�I��V�0 -���㑰�0�������q�������X��$s�?����#dkwh���ߩ���t-G��U̱�n�%��,��/&rr[Oh�h�e������~w!�^{��xE}~��Ꮃ��R,#s�p��w�/#�g>�f�Fo�q�Ub�w;NF��Vgp�UgY���Wљ�kC�;��|'n���H��9E�1�BQRFW�M �r6l%.��V�F��&8�A�#�����_����� G�x�x�ǈ�H�̔(a�9���~����j��������X`�j�T-�zޅ`e'����pt��v���jf3�rLO���E��H�9�#7��\7��9���dfL�c;6�s�����G�ה���V�}>өT.�ڭ���֝�=7��cI8qo��l�;3��tu�?��Vy�M�U]��=�M���MS�mBV�nKj�%yշ�.�o_�
o?�p��S���gf�˥6�[6َ͵��f�/y�rF��7Ԟ��f>n>�Z6Ð}˻�Ӄ�v]=�ջeƘ�yJ�6��9���\���\�#�^�[ղ��<uC�1t�{�z}B��=^��K�<{6KX/�xv���:^:]���4c�v���E���B�Al(�(��x�9�";b�̌�.�U�zܶ*��h�L�f]^Z޿!s�����:��D0���=�2C����Зda�/1i��Y��Fu1L;�XHx��wA6����N\�<k:���������Ϸv/�������^f��=��O����^���r�+�����qɊM����o6�T�w��w^���s�Xm� ��<<x��<x��cǎ<F@���m.���
���÷���$�Hq�&��_th��3A�2T��Ὄ��u���v�P ;Z£A�����I�o�z��^����"�^�l����\w_
��-���=x�b�.�&�Wv�[to���.�g��Ο"3\7/Rs��<<�y��U�<f���g���:NXG��d�ML��#�aʞoJ�f�C�Xf*};�9i����WM�;��q��u���q��ͣ�:�`0�P����5��5z�M�����\K��ᾭ�������=�X�(E��6�d�X�\>[���H&"�O�ؗ�sm�~���w�EU㍷�{V�5��_��f�s�=n�s��n��E�q���׏sr?&d���,�A�uL����p��5��-��m^�맜�y�5�t=D*覦��"m���L�3~@�@1c�ԫoc��>�q\�N�L���Yf�G3��ë3Ʋ��=ڟ�|�bf]��nu��(2p����j��>�ZE�ٛ�{BY����ˌ<T[}w*���߾�<x��H����	@�:��}��[�{�C�`�Y�@�qxT��ͦ���h�g�Qf�/p�i��l���Y�]��(�1��\���7��ot���^|�vSRr���Wb�^�,ޯ����`�u0�la&|���,u���w{@��Xv���4t3��a%xK����ete�8���^��&9�W��<dkSK�h�w�	3y�r��S%��m!_gn�߶�t䍭3���G����8�p���Y����	�qdǺ��1�����>��J�XZ;�+�D��K79cw]��x�� ��6E�t�b}����}�n�f}��y_�O�p���or�s���)I���E�tf���7���4����ŵ��zj�3l�j�j�>�_0�x�*�g�F7�����@����
ʪ�{O���\Y������(�Ͻ����g�`�K�찶���;�og���'hYl�p�S�������滞BQ�Q������:f�H�}+#�����R�����:,�xhcS���,;���3�V���5��nN0�D���;����y�󮷣��pq�pF������/&�t�+��m�Di�=Q��:�0[ԓI��fD��j��aŹAО��W�A�Y됶�ji�
�}�1<.w,O��=�L*�؇���Ͷ��t����`,�Om{���h�ϫ@8�>��=N[�-nF<�u������5���SКf^:�G]z����jQ��ܤ�;6u-mz�%�C�o6	��QZ��ݤk[c�<3����:�J:��1/S6�|�(�v�p��aj���<���LS�D���R
/3�ŭ��ix��y@���+E�!�����tN[�+f`��r:o2��~$�+R������L��?(�c~��BMC�?	���$��a���v�@��
��f�)w�o��Q�O��f�f�XІ��?�:�=����̀𵙆wf���ݑ�D��f��6�E���؛vW1S�Kl��(����#�-��p��R��c���1'�E�Wpm�e��ȵi&��餴�g� ��B��C��Oc�T�dd���7����k���v�7�v�����|w.V��g\8+c�å�TH�1<�
2�Q0dL(	q��$�T(4�S�䣏����yyy//!���V�#cf�L߹�!4Ai	`���07����Ý�u�+�W�[^l#3�vgr&x�s]\���כ׵�d=d�-�ю���xg� _�n� <���)\����Q��R�E�+|���Ѳ���G�V�}\�O�9l{��X���Nj�;v�,�_<n�3�Ly�茺P��o`1�\����J�5���osJ�)�@���k�R/pl�Ī̤��@�g���Hk�k�y���NЩ���UnQ���1g��6�o�w��4���y�V-
��#����sTC3����9B2��󴚋S}9�p�f��J��U]�a���6�����s��5x��h�}W�'�%��fg-��!	�������a��a�	a�<a�عWz�e:����<�e����<ק��.�e�o )�Tc�j��-�iT�|���E���V�#��d?^Ϡ� eSm	������D�<]9ެ�L��-�#`0��o!#lCvM�*�׆�z݌��<ի��E
��;�\��d��I]_�7ζ�N�U�l3�[�؋7<��gw>m>�x�8㋎88��[�sS�h�i���גt�od��I)���uWVs���;W���	8큃)_>OY�{B[���ot�+ԡ�����n��q3rg�+�0Oo�[	~�&��wMfr�C&Za����O�d��=;�S0�/[VI�J�YϷ��m����Â���{����/��̜��9j���ӱ��U�z�s�ra�x�oKrC�uzϪ�G���Ԟ���p���\�\8�Q���AG|�Y�s�3�WR¶�Ś9���� �C:�7�M�M�@U��v[T�:�f���cdp�3��c!�� f>��g(�;�T��KV�"4Fk�4i��#�C�N4o�(Aҭ��O[��Yk7�e!}Kfe�S5I��G�7J*b�&��FD��$p�H�~����1���T��L����������<����F�a򧗟���8���l*�3�QWm�q�┨ĕ[���Ox&˵�VLK���A�e��$�ӛu�R緓�i�wv^<��\�-��k*�ius�yh&A���:�7�f	؜�X���O!���<����������^���qR��<����`n��䭇{�|Qn�r����X}ggĩ[�UXR�l�=W�エ���z�4��Ɋ���]{;/w���9�z�D_l����{C�_L��)�!�v����T�@PD�H�z�����%�Ӷ�M�S�&
9����&='T�Ư:w����ZR�hf�`�f ��C{Ǎzq�'�!y��K�u�e5뛜�6`DE��%��������@J���1�5{��/o#���[3��{%���'�{.a��y��g���� �W�w?m�Jݙ��T������í�	��R��gf��L����K���o��;�j�����v�v��arȒ�n���iʜ�����p]�`���rѨ����z�r��N�5E{�Q��^���v�jP90��F��f��O���b/Xn�'AfVS֘Q̤����̗��>>P�^G���t��ˊDA�I ���?i�'^��|N�	�'�c���$��A���o���Y��cn�&Fm���z�S6�xU��nm��\F������Dw�r��E6�ڳL}��ּqq�pq���/}������ם�8�*W/,/���`_�\���CC��)OwX?�,aoz�{1���a�H1�R�{@g_�_���c:�Yb�����Xkn�2��^c���b8HI�C���/���`м��甈��W<^E�t^���wf��9I*&lIowV�[n*�w���X���?<����#yjhϻ;v_e�i8�{�.Í�����*p^o��O��l��*��u�;��m�2Vb�M#�4�L��]�`Ed��+M�r�B۹��O[��L�q8�ݻ�L
�
9i�':�u��7:o/�ތ�&����2熀��f�m�|�b�t��+g�C=o�S�"u��=�gT�zy%�]W�nݠ'�Y[��/zn�I��u��!�G���;q��wAE�c�M�ٛ��$�33h�UyR8e��ӎ�e�0	}�����xp�>�O%�QW�ٍ�1�u�k vڈ��]\�X�fT���=
��gj�[K]��ڧ~ڰ�]y}>[�@X�x�],6f
������n��)Xw��Jwx2z��!V��[]w$s#S^ӽ�M�
�d��
x�&�5�gO�c�z&�eH��Τ7�l�^LvU��A�-�e�6���$ڜ:�Y�K'ކ,%N��[x 5cI��=�u˵gK���F�Ҿ�l^@��Q��LT�<�Z]Zje�G4N���<X'�j�<�%�N�+�@���OI�u�wf�\T^'�{X�h�34uRU�q	���]�V�����'�\�h�`���re�*!X+<+�F2��ǭ��
��\. ��X��w���yZ�kt�]]gA���w|�t�d�F@ݱ�d����]��tSP�
	�{vd{7͡��󆋚�(�W*�O��z1�jqȮ�W3z���V�N{�J�5���3���w���:$��3tj���ܺ�_MϷM��FB��	�1�m�Uv�](�vfT��8��b�oq�C
� ��%*�I�vK$��ⰺb��1/�.ց�����&���C�T�Ƣ�8�To_U��&��-�}A�=�᧕{*-dŸTP�CC��A�E��Tt�D#�*�R/�v�e\��	�FϹ��}@%%ɲS��ƷF�ї�蒩(��p,�6��<����+�T��(L
ã�n��Y���s��4N�t�����"]����2͞��^�$h��$���xc$� �%ڻ1r�E$/X�;-��	q�4�$"U�-U��AR&�l%C���>��CA(p��B�b�}N�E�u[Xv4�U!�r�D௧�{��gA2��˝T�[0�A#8=�k�^��ɡ�B=���n�`ՏCЧy�\�۾m	Y�e��[��-�TfvS8LYz�=b\�e�cF�{�"�W�/�����u/-��3v�\��N��;-b�q=�.N��<��A�c�!�g�6r[�urx�<�jN�Ue�ē����,��N�W�Z��� ��.54���I�o;�����Qx�'��Tko��$�����r��]!rϹ\T4�Z"}}�uF������/�Ӹ�� �T�ɜ[�Vj\{Pt<�����Gbx��G/�-ӥf�F(N*.����T�v!c����f�b�*q$s�����g1Ů�̀��{�P=Vv�g8�Ֆs�6�*�ք|Va���+om�o˕���q�S`�B��Br���8��7�m���r�f>�KF�U�\�m�Q
\��ʑ��a��er�r�@�ח����q���[;'*���|��
X�}����nM�	�'K;3�&ЭB����,p�� deR�s�I!e�E4h�A%�;��6Ҳ������m a�FdH� ��[���e��(�&DJ��G$$�<J�h�`&4�H���i�f��#��*�23�A���M��.	���2�)t����%J�嶚��L �ؿ!lHK���.�+�6����K����MI�BDH��m�)S��H��%�B	f(_���ED���h���w5�B��R�/5�*���ǏO�����5�kZצ��ֵ��뮵��|��A�D˖�#,��DHDAȎI	$��q�Z־>�>��kZֽ5�xֵ�u�]u��}���eT��!R�XDZ�02I�2���__Xֵ�k^�ּkZֺ뮺�׾�2!+�R�'6��&�u�"I!! N���־5����kZֵ�kƵ�k���z:! I	�*)g��>��I�--FOi9"XZYD���u�2'�������t��М���K�	�ɳ=n'������*L�),�z�^�Hd���"��rC�{�=/�#�ss���b&��jX6���W5�	���s7y7����PmPe��E�V:�ʹS�M�չ��Ρ�Λ����i䚰gs`�9�Y/�W<�o%\�캜�7��#.kt	�E��p�Ti�i��y�$%��
2�H/�޿!���<�������=f)�����/8�ݸXn2H�^-�9G{�vv|����I$�ὠ�uzE�oT��
����2����`�#*��3�g*a~������\z����%�Z��w{���-��T�cw�0mq���u�Xf�{)��a�Et+x��f벎ipah��`ٽQ�J��9�j�8�7r4�S�7q�{';��XUn�{_��X��}��#l~��u?}��uc��<<���3���Gvʂ}|h8�!�u�{�5��v�[Xō󗜹U[J9l3n`"�����kD��5��.�[˙�l�ej�MNv[��4���'7�w�H�j02��F���:���e.��:�������Ѹ�R��{�����	'��~��L�H��>4��#2��-� ����
P�S*�M\x�5��||'շ��*%�*J�z}�.���"�n�^P���tw/�<p�}Q���kUA���θ�_M��iF`me�����
/��G�WNY��z��r���d��}O^�i�뷧j�^A���8'��g}	N���̡�V,Jj�O��w��� ����xSÝҕ���B�������f��{AG���]�[���zW�-��B�ܑ������^�z=�k�1��%�V���GEы�L�2ů��8U��ՙ����uN�{n���.8���"&qX���g��]�m�ͼՅ������k������6&M�9S��Z�i�G}���'���yz[6�ݞ���}�k��|ۍ���j���V�Nq��FH�����;���Ns��2i%�;��]fE���y5L8^qU1��������υ�ߣ�Q�ӽ��7"��87}�5��eW�f�S/&����ʥ2�/�}���(,�͝BT���ˏr(S�/=;����;�Ks���0=�Hג�d��]�Q�a�����2lg0L�x��Iu�c������{�"���e�ӯ��$�6me-.�R�cʹ�Ŧ�b[x��1�G�b	�u���ծ�-R���T�é<���1���wy9e���Bde��,13t�Q����t��9��Ēս���+��AV�U)wdV�)�OHmdᓻP�-���'�����G����>>��u|�ݶfS��;�W��`�"I����p^0f`1�[{Ä�Z}Φ��U��K�\ ��V�I�eAtD;w�eO�Y���!�9���`�̋ˬ;�r��S{�J"��c;��t�ffj��t��'�=�H��Y�"e�Z3:�R����Ӑ݃8g���윅�i��n��FZ�k�ǈ�hL��ܬ����R};�A?�9�d���>��v�������.�b��E��x�:;9��p�w����뺙{/��N���4�E�C�;�+蚘���"��{?/�GrC��~����>������A�u6�a������1#��;�9J9q~�q����ك3B���$Y� 줒����}�^x�U��b��s����/`�mLE��n�3E\u����� z�ޯo�݅�߮/��ț9���V�G�<��t;�ѷ	�,��}gϯ���wSl$m��m���/t'���S�99UP�P�0��U
e%�u���{�um�E�3ĸ�7�E귣1Ǣ��l��Ĩ��YMv�=[c�ؽn1�K��8��-u)!l��­�o������.^�W�����,`�+�ߞw���[η��R����·z���uA^S}�]y�K�Ȗ�6�B�����v�����	m�ng���yX`�A�>YƓ:���ں�b �������vzC� ���$�'v9Jӓ�>��(P��;���a㈎�t˩e嬆��c���Է��B#3͞����}S���nx��#j�6�/HއW�#��O������) �����z�F�l��������vg�3��}Jc��]Oy�р7�%�w�4W�
Fx��"<���R�?b��/o_��h? 0�?_�▂�?E�Y�� �����ΪZ���Cy&*�ԡ�R�Xf��ZQ��o�b�>���	$6���֑����VG�{b}�K�f�m��^u�}'����WR����z}!�>���ULK�lt��܇�ߏ�s0�x^����O{Z�
]ś1�W���RWD�e*ӷ��Rh�������(�|%�v���z�$�|�4�5�s�/y�u�BBN7T��mv�ǵ}Z��nC{� ���ŷ�g�����A䤇P�>�N�s����f�f��O%@���a���Q8�0Bӑ�m6�Ԫ�q971�/{���ns���J�U*�BJn�L��nW�o
(p�P%�[,���RG�~����~�����}�9�%r�O��~�QT�mw�3Yۇu�1�:9wv9�:D8yp�ϊ���z{Cm3k&ء�[.�ӧ��	�����O��c�,㩉����'8�u�e�Yv��a��e Ʒ4�pș�ez�C�w��#�4[�C!�;T56P͜n��a����ʹ��F��8�8��Τ��!G>ϑ��m��Y���+�b��X!v�kVծF2��)��K����u�	�Ce��&ʭ�:s�r�F<�z!X�igo0k�R�/,&�?���R�ͫW�%fҬͽ�a~KLaO����謿EV�������Kwb~����[��T	����z��!ll���
�fvgp�ϵ��-s������+�Hk��K��U�ثDb��ǝ{�KǪk�"�ٜ�7
Ǽ;�gVr�㝵0lQ�7�啯���� �=E���<~�*��ˆ��Kn�*���:�9w��VJ7M���>��@��˸�,�?q*�6�	��b}�q��s�7݀��s{q���5Dy9�۸q��y���'���yx���<|G�'֕���>��%�����;C�O��,�@���t�>��s}��a�� �h;Kߧ�S�u�� �W�P�{�Ss��x	:p�%�-�||�2�ŽW�z3�<�ҟtc�_��ɏefU^^�y~9�-j��YΙ��A��шDҺ2��U��6j�Uw���FCj=�l᝺]%�3����A��� gJ�g\�.���J�}�dA��s��w��Z�{���/Z��qS�"����\��	S?t5����u���0D#;�����������LhԾ��2*�w7���P"���6�|t���������Ʃ2�=!#����ybCf>�G������ĝ��loy�=璭�<s��Hh�9���:=�7�wd��э�CZ*�
�N{���,�P��l�&����a�j������{�;�Y}�v�o�H���|i]E��gto�Яݻ�c���ޥ���r�hV!f�k�YU#�.��e�r6Hc�����n��7�X��ݹԷ��"͙N�E����T��)�b��~���Q�[�Y�6?}O�������u;�����s�d$y����m�!��0�����v	��.�OW���+Z���Ǻy@2�+�=ޝ����w�gNK��T� ��q���E�������yUzgگ�y�]�̽�}>dP/����ql���K�b˺㸲O���o��]�t
��7���>��$>wK�6��"�;�ۨ�YZvs��0,6,~�}�3�wl"����$�8l��g*zr�o;�����C6�Z���eU��g�[�o! i`W��۷l�>�ͳ�g_W���,_�}v�s7�e�T�S��	�}�#z���]��kN��%M�Q������ (g[����Tj#��.;��",����X�o�(��	�w� U�f=b�����	^ioz\���ǖ�|3��m��?���;kL����vB�y���E;n�躮�/���q��wi�Fv�Z���Ũz��DH!��ĸ���%�m���]��zĳ\w�w����̑`J0���R�1٘�(j��)C��21��7�u�<霮e��.����>>��>#������ߋ���y�o亁��T�6�7!7j[Bl���]����z��O�#�Nh�	f%eY�L(��*�y�%�\Жt��r���-#��26�0�]�]O�/�R<��:�r%�8��[ݑ�b�വ�D����sI���j�Y�'���`�]ٺGOtO���E�p�ǻ$2�Y��i�Z�)�;^�%�OX�pu� h��,7��ϗX�8�O��-.X]M��InW�Q'�-�s�[��N���p�����<�t3kJ�8J�[kz@���{�Li���}�ջk<����0�4���DG�<ڞ��z�k���łݡ�*�� ��\�N�X��M1��D4l�=y�^�&�����&�C�<���=�I-�rk^�s���#{C#��[�p48¥@E��\7�|?J?f~i��C��Lvb��T�hvZGy�_W~��?#����EϷ\�Q���X�k�C=
���*�`dz�#��F�뾠:G�am ��y"a��b,y(���Jٝ���]�y�:]��w|��R���5�����͇ؖ%<]��2u�zs�[�*���ۦ���-� ���� >A3HBZ	�h9	aA��9M�_��>��>>������*�^�s�K�"]�;��cO���C���kA�Q��.S
�]+�MU!Og,9����{+v|I��|nEC�6�"��(uy��뭖�r��s�h�n[7�������玼�j�Ա:z��";2 C;Vw��R~�d1�3&o�Do8�>*�	����auoM:p�#��z��
��H��Ͼo6�)�'�W��w��_ �D$�@�����TW�
���'z��S)�j��U�s����:��,�Ȭ]䳞h�L�d����7+��`�}}��7��=v�`Ɔ��X��Rӽ�~�6U>�'Le�����}�
�՞��]a�<<���װ$v�i�\� XD_�k�µ�@5�]>'5��:����
�{�b�yF΋����=�`X�6N�ЃB�O�㦶#��k�q	�"�����]�,�m��^s/;�e7��ubV�ˠ)y3ȇS�Sѫ�N6��6�7ﯦ��Y��h��wIsЃ @�����1��� (�|�Ay8�:��	$��4��/kAJ]�9����mĶ#'MMJ�����ĸ
֌�b�q/��Ȭ����gS$�Ԍ@c0c����^u�b���XḎ�=���;�&��޳3m<��*6�ƬR����>z+�ޟ0�O5*?��D���)0�ې�����{t�w�q�w��0!|�0:�-�yeg-'�6Cۄ�go.9oo/��r�hFC8����g�"�z�8�}�C��}�8���s��0�n��p�`�N��!�����f��;3UN�<�R�*�<Qڵ�'�(><��;-ff_pA������{/~�7���e"�L6A�f���Y"=�6^h2Ɇ�(v E�G��J^�j�]��t�)��FA�(g���cT����C���4.Ǘ���8�:7g�޵k�sN�p�' C���U�mj'�=�w,���ݨ�l���Fjs�7�⭟�3�S��3Y�i�]n�S�['J���
j��:]v����m�;~�t!��ln��MX�Z�^ٓ�_Wv�k8L��jL\`r�0�ް�YzU��Gr!L�d;���W�h$4#窥��9:�FN����.kځ��{l9Զ���N������,w.��󄒒����c[�l��#��d�1� 9��ݍ9��a�3N8-�̂������#ܤD�_kWVY�9����"TB���x_��	��_-�vB�{u�ȳ���w�k1\��b���1!�E�D����;�zm�����oU�wX�v:�9�_;7;-`�, :h��+E1|�ѵf����U�+_.Ҍ�-c����R#d��m�N<0;9%������]��9��W�����.���L�ݬ���6�}��\-�F�+#2�*����5�[�m(�#gI������1�u�Dk3���㗐^����g�3e�x-����+����f�={���@+��v���x�l%ދt���ʙm�a.��x i��5$�ɕ���w���L���z�dR�\��^��L� �����˳��\�8��D��Qv�R��wh�qQ=7�W2�+t���tw�\��9��nJ#\�N�b�,?W�w^s3}䛲����Qt��4�ƥ�2��V��Sz�/#ޡDTV3�j�]�3���A7)�#��4�1�]�mI6SYz��`ʺ{����y�hH�E��x�Ay��"��nA�WS��zK�1�'�������ѭX��/��]ޙ4K�$�����)̀�G�d�8C���H�f�U��w��x6���.�Z0��[9��hPX��f�<��]1|5'*ﻥ˻�\�\ҋG.p��yՊ`=u,IdX���ȱ6�e������H��i���`�ϦѲ�=Q05����A �Z�(��p�v:��1:?+-�i�/뙎\�r�sX��v������3 ���ꏎ�mE�{�L�Cw�^�k�z�^��ţ�o0�M�=3��}Ĭ�2c-`�ɏ���	�6]v"���N:wb�|����5���� �{3.�ǳd�a�`�Cڂ�=�}�d�T��涭�z�����&��ۜÞf��<�X%�ro}Z���1��n75�!�eA�c��)x��bwV��7�#~ޣ�찼�ݺT�חl�w6���
�Tf�y3���Mi�G� �د7�����l.��
8��SrU��|�oQ�̴�hŭ�=�F�
��k�z��q���檖�z_J|A�����gi�Jt����g0*�BL݂�j�bˣ&ä���pwkȋ9�+���cV�ftݝ��d����<�;�[�[����IN�C�b+e�F&�
�wy��qq�g3�VQQnh��S����y4��&�b�b���f^���{�Zjۜ1Y�,q-~5�}��'��ݐ�*D�D�;Nz�u,sn�U�q�be�^ؾQ�D�qY�`��˷X7��vZ�҄oU:�Yev(A�7nƷ����"������mRUՏ�ɩ�i�ư��:iՍ����O��LcB�(oF�Y����?��چ��'s��{�z�����jv��e�v�m呑K����%�V
Z;�_:J��t��`2@"��ED�9�1d7��&$�>�x��������5�kZֽ��5�k]u�]k��0D�;����y�u9�ǊN�94.iQ�s�nix�ֵ����kZֵ�{k\kZֺ뮺ף���gS��2#!	���^m4�i�9�L�~�]yk_����5�kZֽ��5�k������������Vi��hm�щ��sI�B�6�4��˱bl�uǏ�������ֵ�k^��ֵ��뮵��I��I��,1����]%�ɨ�>�H^�Y�����0��8�N&l�b2N�Hqd�>�{��XӜ��<Ӽ�;�9��s��ђn�9���K�dx��Ah�h�'ƚ3ӎM���0��t؄��e�S B����$>�y���qx��4r&B�2q���Sӑg1����"#i=���ǀ�/J@"�$� ���N��bZ6��=U�h��c��Y׸�X��Nf��[��3����r��8ŌX�#N�����~������p.]��:�q�O���`���y��6�nVj2\o�
��T!��@ϱ�z�k^���nQ�-v�>Ŷhũ���Q}�I�d��a�ʽ�L��w�dvmy������tc{K
�hiھ��=���b��H��'lWD	��=ږ�I4@�FXE�U2������4�L�
,��a�3��	�f���&>�W����W���Tv@Z��g܍���>�{���)i�;�Eet���8���|���
�W��И�	�K^I �l�#ӹ�;9�'hn�t0#wП �Ҷ6��v1ev�I�'R�)�,�~�H��?�FѣK\��3C�f�+35
�m��B�W[�3/TJ��p�h�K�Tf��3{]��f���!c�O��>y��z�Sy���z@<}�|D0n��?�	�_��������7��WS��%&��u)z�ó�E����f>Y��U(�HO|_N���Uִ�\���7lwv��q�;WV�:�I�ť]��u��zjQ_��@> ��i%Y�n1_
T�#F��^�~wfv�{�153T�0Ӻ���7�%���Z�@&��/���/��(�/ܧ���/�&:CW�xWFjJ���_Gv[�?<�A��ͯ�w{�t�`~
� ��a��FY�:�5fQ������ l"3�/�Se��$��3������Z,	P�Mr'�d�n�#.�60"&���z|�)�����5�~��y���pf/y�7���`���
ڍy��`�˛heh'/��W�Ϸ��;/���Q�J�Mel&ʯGV���� ��(q^�_�X����}�lu�;"bc���=�l�<xDY�&G�\Fk��{�)�Ƌ�R���~�>Q����6�zc�k��GvA����^ַ<@��{b}�Dk��d�g��H�����V��չ���}(��^w*�f%�.Z=���>���YR~�6;���p�ͫ�xno�*�{�xML���6nr�x%���h�t;��뎪�>�Q�{�|�(5e��NP���MH�Y��6�Q��V��w�-��y\t�ʘ�w�d�r�>�<�v�WJ�=�h���>�2_E�&H�QSF�h�ϓ`2ɨ�d�'��ČQ#�9�>s�9�y~|��~�Uy!~Q�'$K��_]}��24�ܻ�ƛ�Tf��<R6�z�mv(����pq86�l@۞_WN��wf�R�{�^��	?�]r�g`y�Yy��N7E�
v�� ��&��w@�S�^@���9]5/(1�ƛwn/���PEf�걔�:}�a�T_)��fg˶<X�f�K)�����j���o��N&t�
0@� wu��R�.�Q��'��F����<���`$��{v���]k���;jK ��z�VGm�ݻ��cf�9��z7H5�͝x�<.�����ݵ�~�C�f���Y��H�KE����M~b"G�`���V�W�M�����:/�uU��v�6�J��e ��_����c���Ë:]����;	�hvA��U
ڎ��m^R�w��}4���6��r���W�?k��c㹐�ɴ�A�f�a��b��ѵ��m�e˴L���pGΎ]�*bD;G�e������ۼ�޼V��o-��\]}��"�SaO��_���}rIY-���-:���s�Ǘ;T���S�u���d-n�'rY�h��X����κ�Ϟ޽���מy���y$���cq�O�N@~P|;�b��]ę��6�X,ߏp�d��1� �`5OO�v�G&}����|v�m��2M�f���z�=ܨ�ķ|������Ck|�]���{�tv�+g����ɾ��s����Wإ�����ms]W}�٪% �áw�G����G5�~��tng%;���W\��t��%v��V��S����$'��e��J�� j����y�o�u[�_g�]t�`��`�������ё�3Y�ih;�Lm\xW�����,TL��vE����nqy�z[�7�	�(
F�Z 3�Sc����v{� ��6�u;(g���w�I�1���07B�C{lo��Em4pv��O�4��fr�x�
-ռkUn0qR^�o&}�m��Ɔ_��^u���6a�T.��s&!`�t��]����en��ɦ�0�{���7Ll={}��bC]j-�OgV��2�2�MNQ�3;q[��n��&�I��er�f-9.�����%��
sv�T>���gbXU�Fd���x7�����{��J������i��a\�2�\�^�g8�LyNf�u�`;3WJۣ�k/O
�Q��+Þ�W绞��/]��FQ���q��8�Z����v���F�lD`���zP[��
 |�q�-����|.Y�l�Է�b�ݖws�إu�@V��1�t=(>z�=+&;5��>��vm�E��̪�W�>��)F�E5	�!G.���� wr�]�09>;o�0ߤ^;���c=}�#� 4�FG�І��[�x��0�fz�5�Xm�5�ȋ��ۇ���7���סϪDz�����-�c��nK9����S5����īg:��ÿ�;^��g�ao������3�ٟR�cA��|�.�Q�&-
�{�v�E����ǜ�u�Xe��2o`.��\�9:����񮀫#U0z��c#�&<Dq��������L}
s�ܹ�Ȯh�"��!�7d���JX��֠�!��O ϒ�ߴ+8u�σv���oZ7�%v�5,�}�ta[Y��t��ۑ��O9w֧YVgn���.)�O43/�~Sf��v��r��j�wD}��1�X��o���=�|�����߯�|d��.��MM>�`�!�L�5��n�;��x�?y����Eo�نI��N��#���m/����{r��N�{�n/��@
$� /�V�7�߿3M�=�@��6'���]��x�2I��*���#}��6ݰ�J|�}����k�1���uz���l��v�B8ϧ�c�����
Y��y��Ǌ52%u�7A�u�=�@�y6%�7�d�oS�l5�,;���MG�cƞND���a;���������3�i���6H��'��h��|��o���� H6Ѷ��#��.�[	�S�ө�,���rgn*ڽ�-��}}81�.U�#�l&��2�pբ�F�>�K�T>_l�a{�`��Wn�q���w�FO����y�Ǯ�"v@U9D���3�N�ɼ54#��5��
��&�*�jː��;F��ӏič�Np�b5
���V���]VՄ�2�8/;�
>��"��l�-$H�}β�ls��Й$��>�r�m�v��S��c���&]���;�v�X���!d!Q�T��梂2P�$:nzR��j�-�$f0����� ��|@a�D�v��S��~�R�-�a�����½6��~��5��Z�8���z���û˭�D�����W�z��fd�qO�oy��`��z)��76�w��sN��;�ej~�:�!��}<{=��ָ~ʐ��)j2��^���7l3g���E���?�t)k�5z-�k�*հٛ�݊E�0L��
>rI�}�����>�,�D�O����C��+��&�'���}#=��<��W㛝���ޭ�'O���<�����)^{]^ꡲ;�ڽ����3Ϟ[#p@]�8��3��˓O�©��5���4VN�@�M�O������\�oF j��_��싾�si�o�fn|\D�tߤ����)7�����"����;�F|ޟB�o.v�؞m��׷�ga�wN��^��b�/LZ����d쾻O��g��A��6k�Л�ݽ�vco�8佾ۛx3�?S��9B��>�G��ώ��lF�ͩ+r��v����m�W�"���Y��v)³Qɹ�)p:{'kw/�E�ݯ��nl�����צ1��������^y���%���oM�2��N�!z������+����"b�(#��wI��a�	��滳9��]�ZDS{U�IU�̷[�b�j�V��^ϩ][�������5G\���s
S�aV�-�x�*6�2GX���I�RK�:Q�@������=�[W��>�ɪ���'?`��s�@W�����&���S��t�>�x
�?(r;20���Ub�:{��q�_O_�apQ}ݲM��LO��<�͍�o�P��������`�w�8�3W�?����'�f�T6@��K`-��Fx�74P���\��Yӫ�u�q���u=�4b=���wv���c��{�;�*�7�u���ת<Ür�s�a�z9�#�`ng+��+6�kO,r���'���`���7���B�h�^�_o���g���N�������_\M�@sMM���
��+�M���;�]�o�S/�+ ���p����poy:��m�$r3�K{�w�Ot�lrq�bJ�v��3h>&�V���9jΜ˖��o7���� .�^b�Kkg�EJدO�\l��7�1
|C��9�՝6tďL<��߷>�>	�+����XI��;���"`g���L��:�Y���(р6�L ,[�����}~8"2v�sMW<�Uw���t*ۉ�*���߳��+l��
�=�u����l%���{�� H$"�⏈�a����b!�>�k��]T�zȬ�)F^���������o����WM~=�Mx%z,v�v��۵���r��9s�ף��NY���f��rwk���7/��� ��A>u������:�Y�����<���wo*�)6�uq�n�U��W̪r� Db�'���	����<�|C���v�>�`����c�\�DGy�箊�J���r"�ݵ^���ؑ�6����[[���Ha�߫I6��y���B1.�\�BZ�y�ޙKW;��h͋��.�w�S�@Ex�H���m�x�8�ɢ�y�{�|�˗����������h=�;.R��z��kD����=zFm��fvX�仏t]�����ul�0�ɝ��=
�1# X�z�~^�RZ��K�[�:���#��������>Q�dv7s�ٙ���n9��z'�}��5��@�:�ff�!��k�kw��b�H�&���H$��4��~��I=�΀����-������o�3��p���B�����I����4��Ѯ�Y��"�5Pfg�� Bp.F�;&��k�[���j}���w���oAU��[��֌B�z�3���˕kN��a�bu��R���%m�p�R�����`�7��Zb�v	|�`�aϐxX�;�����~J|�'�Kg`��6��A�W��ohFw������z��Y��%,kv@���<��ax��~9��;��I���y�`nS��f`�Ch"M�^��W3U~ᢨqf~�_h�Ӷj���Z�z��;�3�f�e=���������޽�#��\��S�_�_�?�* ����3 R��:��	� q�TU��إ*�j���U�b�A��b�a��IV�*�����JT�J���m��)VI*IU*�*�*���d����X�m�UQR[T�Y%��QR[��m�J��VKb��PHȄ@`���H�U��%*�$R�U�E��� ��H 1P�H� !2A 0��BH��r"A 0��B H@ H 0P�� 0D��BDBH 1��A 1�� HDP 0@��BA 0@��BE 1@��B`1�� !P 0��D 0��BH ! 1��BT 1P��B H:��WE 0�� HD 0@��A ! 0@��D 0��HD �D 1P��BD 0�� H ! HA 0��BD 0�� !A 0��B 1�� ! H 1��BD 0P��B !D 1��B H 0@��B !A 1 ��BP 1P��BT !�H wT�1P � D�1R �QHU  T�1��8 � p��` �1 �@ Q �1 �@@  �@pQ2@ �B � � ���0�1@�0P�8 �D�0D��HHHH2 �@B � �1�HHH�� � T Ń �T �`���8 �A���2�HH1 � 1  ��H1D� 1��� �0�H�)RK$�*Y*U��RIb�����,�e�)ddb	1�`"q�`1��F1A�9���p0�~���(�H" 
F
$����z���}���`~������?�T��������
��?��?��~�o��rE������DW��������� ���DTW��?��>�?�/������B� 
�����I�Oǌ�L��v�� �x�h��������*�"�1@�� H
��B��� T �T"�D � H�P") H"��A � �@� ,D#1P�@@BAB,! P�$EDQ�E_�H�9 I	DP�$P��B�	H0@�	H�DB$#$" �P�AB@"�X"A(DB) H��B � �B �@��"�0��"1��P"�B��@T7��L�����'� ���*��   (�?C@���_��~�@��_�4�;�_����������?_�9؟�R���a����������DW���$�?�?jyP_�DW�����dw��y��W� ���L���<�p&�=��~�L���@�Y�������n�" ����?i�������������(~��X��_�?�;��D@i�?�?��Q_��;�ht&.����0;O��a����z�x;��_�ԑ�{{?�b����������q/��Ex������.O��o���?���O��PVI��v�$w@�v` �����������-�M����j �*��F�Q[4��D����ƕUH�%!E"�D�ڢ���T�E*��-aR!T%JF���͍T���Ͳ����KZ6�����mYV����kkP��3%�Y���@հ���IF�6��kc0���l�V�e��Za�2�J͵X�����l�R��YJ��kii��Z�Z�h���%F�Y�Z�ZUdղ�m��UE�L�j؊5Z�̙�)m��l��ZU*��4}�  g^��%���m��uv���5ٚս�ڰ�[�7��u�m��ݺVյ���:�[4�V���J����v�5��j�Z�W�+*j�v�fV�mm���cU��ZP�6Mm�   kC�hʔ�)y���n��D�ZƆG۹���e�i����I̭��;�V�����V5�j.��m�[je˄�{8'U���ej�V��*�6%�C�Z�M�&�Z�ʶ��Vͧ�   s�UD+{�E]E�I���J��iѫfS 0T�+��)�Ϋz�����ݶܓ����FJ	GVu�Bmkj�Eڳm6�ֶͶ�l��+X�w�   ;��/V��v*�6kjv�T�weWf�%��tT��R�أWnv�Uge̝i�ݩz:⪠�n��m�@n�Ʀ���U6ٚ[Z`�m�   ���.��8�cj�53cUq�RP�㫆�*\)UZ�:uT�*���EC����(�Lʨ�k.�fն�����֐��   wOUD>"�>ۏJ��+����
S����EJNpܠ �nz��*$�N�K��*�޻ݽمJ�Wt^�R���xsĩ/a��P�L֚��e���S*K�  0��V̤��}���K�)R��+ǉ��Ӝ�l5UE�^��JTHK=N�eE%�3u"EQ���P����ބ�S�w��ݻ�Q��ٙ2��-e��+��/� �|�%_<�ޤT��Gkם�d*)Ug.�R�%+uzs�V�=�M�UD����(�"�]�7x�U.�su=�%;4��{��ޥH"U�'�fk6�Si���L��U��|  �}�E
�wڞ���0��x�Y�=̂����Z�����W���7���s�������<�@B\<�K٩S��+u)Q	Kw��ՌVemKZ)�f��Vl�  ��f*JI�w�(��i+����H(�.�y�B��]�j��*Dj�z��h{��9�ׇ�)UJ�={�D�R����p銢^�9�y){H� E=��)JR   �{FRU#@24Ѧ�T�yURz@  ���R�@  O�05U$�   J~�)!��  �f���~����:�����^䛜*����>(xX���b�C�
�I�eg�U��}�}_}�可�+������]wuWw_�Www]ww�����]��J����wWwUwu��������}�?��V"��?t�� H���F�F9����w�ß��#MU;)�F�_k7 ��Tɰ6�������(,E�'�+݅�8���CŠ@���"Zb�J�
�ټ.F���f���%��V�5��d���E�X�?����1X*PV(	���^BI<�8�Gw�C{Ǘ<.p���.�[m{�$��fa��w��M�D�� ��2۸66HqJ����(����N^�蕻z��1�C�e
6!��t�G,p��ձ�u0���X$�^Q�b�ce���fk�@K�"����h5�6�̀�\SV���Or�g*�F=DVd1}��9�t���#��	Z�N]�U��f^�n���Z��f����!�W�cVv�N�'N�X��
�Gw(�خ�cooh���y���ed� ��$ݖ���/1;�u�7�cM�X(VM"-<��ȷN�f����'c��ʗgV�5Z*_�[�^���Qd�(��4֫�Gp
����ˍD!I]n�!h�7��č� Y@1�7���u�Kj�Hn�AVŸ���J��`�jr
xq\S�~)�ڍн�s/�-Uޡ+j6�Ժ�w����u��1�6�̫%yQ�g)�B�&�fܼâ*���ڄq�bLRMm���tΖ�K:6jU��Z��E�X&b�+ZN�L�ƳH0p�l��g`Y���`q����4z����b(F�Pֹ��4��kr2Z���MDO(eF�m�Ct�0FL��}�zs����I��1�6*��6JN	2X̻"����h`Z
���M��@[3s/^�+ ����/c#Si���f�U�{c>kH�ً�J�Xa9P�R�f �-7��JqVV(/4̭�r�}��;�Ġ�-��z�t�{���6Re]��֛�M9�7.U�l��ێU{�2�^��mDoC�f�Ǩ�B�QJ�aE,��+l����nԣ�����9�Q8�I�m�zkY����p=K����'B�9zk�M�6`L"����������XհR��9��M�@��
�6�W2��Z��d{35�Ձ� �[��P���JV�:]�d� ��y��� �Q�n-�@X��M�eC�j���j�=TZ�-ņ��7�\Ŋ�:�Xݚ���F��t�0�퍺��+%ۏ��t6���Ѥ]���b�%�(KO�ԡA>�D,ndZ�7t�@	;��n��ʻ�B���u-`�'X��FHl�p�PU�2���B�vM�K%m	����1Q�T�������t�j�����ߑE*	jk����^�s]�*��-n��A�F��u�[i+�Z��-�p^4�h�i��bE$t+Y2�0rbx�"[���0��%3g~P�Rj@B�M�	�Vn���-'uPEX[��S*�V���+��K#���ч���sΏ�!�b�+�RO��CB���B��OU�p���XbQ���Wq�7c/�b�f���J�'4ڲZl�8p���k6\��奯�q�C/��X�n�t��L"����[��k��'(�NYZ�+��stY�BTii͈^T�hn��(�Y��O1�B<��K�ԡ����s	��ǔ���]�F�̦�eM!Ϧ���˫1]��ݰ�Zw��"�%��
WW7��]��t@�Ҥ�`l;Ծ�z)̷��VoU�����$T�!IbLZ��(n	v�ۚ-ݼS-[��5��2P�nܦ ڐ�(�n�յk�wGk0�a���J:Ň���6�Z�1�³�MW&�f� f�tG�pMx/����p��遌���w�t�� ��6� M�R�=�0�+r��km��x�ϲ,��R=����U{1�6��bDVie� %^�m���c1]f�AƬφ�O�ր:i��Z����1��w`�-h�
]��h6�V�^�%�jR�`
�ĵ����Y��k&cCq,�����K�ĩ�FX��+,�k`��"XS>b��;L�z ���ű�b��E���YFq����fl1-�޴fP���٩-Tj���vZ���9���V	"H��ޅ|�{x�d�xk*afJ��f�݋�
�dt1��i���(��髉��k:i��n���K!ŀ��N��߅h���Seǌ2pʐ+f���X�+�S�v^-ӸJ�
]Ð��r��7f�i�y��ж+v9F�Qe��ql5s-�tkbd�B�h�����Be�n�Ȋ�B��ub��]"4H6���j���0���VZ�/&�p�:#i	�{�i-@S�%N�*��d���M�WI����j�M7� ٍ`Ԕ��tZi�*՟��V.���ly���DR`�qAkt�IR�S�[Dfܬ{h�R�\X�A�h fZ�p*��m4[�<�C2$.��l�`��c5�w�ko7*��2c@�T��!�ʕ��{��4��Y�`�@J�x�{#���|�ʷ��t�Z#��I��V#fl i��2Lݢ���{L�KV�����	(�Εr8�!�#�A��P�8�!be\�-a+y�ڰ�񷊖�b^V�4A:��w5'V�Z��eXt��P�5h(�׺�5����I��n��D-$�u���-�klS�a��-�^��ͭU sU�����R��:��cL��{i�N]?���V� ����/pֽ�6,�@�mk�v$7��oS�ߦ���zBu��j�KC�{P��(6B�n�:˶RB�n:x��UY�I
���%�[SR�Q�.:pFf� �*�ذm��&��J˲�b�a`J%�oSѺ�@�b��/��*p
�5l�S5=*�^U�4H�j6�ca�̡���D@���UXܻU��r��iZ�+	4cz��miɳu92�]�\��m��E�`Lov�j�ɵVrG4u�zSIs$�.cv"WX�Ѹ�t�we�W"�PR�Z�m[:�˵�	��X��.5�*��]��6.�F�yt�ۻDaT�� �
A��cl]�i)�nc#2ݗi_�ZH�Yօ���eށ∴�W��\����֫ǡ3(�T�t��e�CQ���Fe5.L���0��zU+��b+��N�;t��Vjbv4�J�������5-�D8���CpK[
ɛ�.'BǲvW�(�F1�m��F��5��l��e�h�&��[�7�a_�j�^X�-�N$�e��e��̭5�P$�(c*�� �̿����r�Q�N�5�k-UZ�NԎ�#U�7LZݑ p�[�Et:4&kS�n�2��V��D��
U��-�pb��t�`�Zl���L��n4�l�u6EZ/	� D,�u������hY��I��(r�Fr�͈ܣ��&m^0l�AƅI��-_D�e�'(f�TH�Փ�����vL30���5e�"��ke;���?Z�Q���ujR�o/T�ۻ�J�V*�y�-��J6�['R4�%}���5\+k3gR\�4`Tp��,��a��4�o�[��0`���
cjjE�9l��2�]<�x��n8������#¢�)���5A�&Vǥ6q�T��ऋ���th�H�Ӎf �i[n��i���Lَ�F7��t�HT�o"kE�HV� ��Mtj4�T���f��Ci�DI�V�L@
Aܧ2T�"�:c6r�!^lư%��FH۶�YS���'�P���eԺ�z�-�:2�	��Wx��V݈v'��ۤ��[q�M�92[�c�Wt6�^�բfZ��mҥ�<��٪���T���TvrըC	�W�ۇ�Y�Z��,3
	5��y�H�$�J&�Xo6h�Gp�55�M�HX�U[��ա*M���f�VGm0ա�2�#1�bV�k-E��p�6cڹ]Z�����FdaV�E�[u&L ŷ[�biyQݰ$q��YgwSiܖ]ګ�����*��I׶����������]m�&Z�Эh�Kq�����cvi"��m�1;&�;��1e���Fjf\r�F�IV�xC�+P=ܽ }�c��v0�55C7n`Q ��,�iۼ�f��ԁ����ʄ�[*���^Մ�I"�eN�1`���k�,��8��Lҳ�H�`��$�֫�]j4A`�����	�R�f�X!a�,n-�$�P�ZZ2K�E	YA@����i���6*�^�����h�
����e+cpe*��iQ7P���,�t췄m�,�����n�P����b�@`ڸ�8��{�MD~Ј�\�W���AQ��[J^���Yu�vxƚ� � ���DVd�3�p���f��J�.�+oQJD/u�����A�Z5��cw`�M�(ô�j�+��a���o06�-u�P͠�Y�(6a�@/�@�d��������m+��(Qj�k��,���<�X��h�4�YNjưk��Q�+�Tİ%D�J�����4��<�č�m�3&n8�d�(�V�.�iӵ7YKLے/�uX[�1��ā��>�%��YE���q����/U���7-cq���$�.S��*��QZ� w+ݗW��n5[3U�� �*F"P���`9�����K�B���HU�u����!3R9Su�%n-� '6n�bR1G %Õ$���Ť-ٸ[�í�.��%���\)&j�+�J9�x�TV��U/^K��Ʊ�D9��bجn�Ė�b���H�gI�w�se,BAVN�Skhf��%:��vo",�@ɸ��	�3P
3B�P��I� [o"�9����R*x������ݣ�2�����8�'А��A��eK۷>ծl����*+N�c��ʋI5n�c�	�z��WDP�+u)%e���մoXH C�hʳ(LX��c��X����[���+6����G�F���T2�T����
x��IL5%fej����VVk���֐	j����h���-�FA� `�Q�(;P�pԖW�a���Ի�7/#F�̵��h�.��ئ���˔�����˭W�-ȔW�mQaCM�B�H�A� �f���2�7.��E\�ݰP����h)")��a m��Zr*�3A%�B���w i=�HA�ॕ� zs�Y��1��t^4hY��,�4�QdM��髶ɶ�mbg-��v�_[� lѫo��m<�׉��z�f1��&�S.5��xѻmS7���ɱVÉԨ�دJ9��%��Ar�7j�`�RYƩ%YG1R�s\���v�4�GnяUn��r������ץ� �B��Z���w{���Z��`�XM]�[�>e�.�O1�ڤ��^�ҦonZ�H�Ӳ�{���HijW�Y@^�兤d'�r��i���T#PR��ۘ>���]k��6�����"-����]W�+S5��b�4̅�i,۬��X�j �L;�n�2[���n�%�ac+ijU����S��!�2m�V�һhl�9�b��-n�Zm����/ ��in�l��>TuN�h�� �D:$[HS!��H؋qPH�`�)f��Y�SK���	w��8{E=W��jc�+��#1���YD��kd��G(����E�%�Yf�f�z�Z��ݕ�䅭M���V ��T���ocm�j<��O)���b+j-��կn�慢v��4�52�e�E3�')���Y��Ǘ� �Vo.��#g[i*-� @m���Ca"�%�Ѐ3`Mu���ڳ(*ةTr��l��8�	��d�RKP�i5*�/,���e�K(	�v���SpHس��e�IED��x1<��N7u�V�ٷQ�W��FdaķsSR����A|2V��V���ѻui{����%��ӕ�nT6����Y�|��W|��7�0���f�嬥nq5,,sl\�ܗ��=m�h���6�m6�V��<���*cin����yM^BX�Y�3�{���Q�"�-&�:�?�m��s!����qڸ��Y�Y����/��D��9��N;����[����-���,��%F�-�ț�˷�6DƁ�u1�vzs@)�lEu�(�f%��M�;[�õ�[�U�)&�C���E��³�շ��+V�N��vm;Ph�)�����CM7<4��y���A��dX�c44H�zw�IE���wB��Z�L��
�u}�]֪E���-�.Z�U��y�!K ���6ZȔڻPӁ�z���2)*�����u�-��.�Rr��*aK�-z����劔j]k���ÊӨ�f@�I�Տ1�Ʃ`�j�b���q*�7guR��͢�xE ���]95^dM�ڄf�K�4-�i��B]��Rh�j�+mU�L��Ro�l�V&IqRT�[�����!c.�=@���;A�L��eցZ�n�U3h,IX�&��n�t�B憲��L���#�f3#��l)�3f���sj+�#�[7�1+X�!	�n3r��YH���,1Ed�)Y��s-'�]�-�t�]���k;��4�mkl�[��7{)��b�`�K�u[,srSw-� ��#@
��Րb�aJ�x"���飉�T��n56��{IЩ���1�ehݹ�B&	�B�G��t�A��Xɕ�����V��:J��Ze�1����xj�ś ww�I5i2�=��=��75�=YkfEx�n��U�v�ͤ�F0nVS"��C�w�f"���գ����cr���S��PJ�=%ݼ�ZƖ�5XF CH`EZs�*���`�f�%��kF���&�"(#�ko�i�UaH����Ő�f�J���q���'�4ԁ�R�+6��v��t�������TE-��Q�ڸѺ�ZE�6��Q��[������6�����.@^]Lx�1���ך�a�#.������w49ď�W�h��εc~@î�����9g�I�����1�k�:�}"��n?kOH��34y�����)�-\�l{������(g�KCB��,��c���Ыf[�m���pX֏R�ZY���r���eX���,$�KA�	��O]���G^ٔ�[�LWOe���e��7~�{D�xV���G֯N�=)�<��a���Ab87�W$�gJ�g���L2��$����V�l����݁g,Fa�W`��m̝��#�a&r.����+zb�4WaɽE
�C��I�XKڶ��"ο���G���zb��z�ݿ���xjo�fҶ«5x��'C"���{4�V#��kő�^c�b{�]��q��|���� �kRz;�t]3,�`>gr]���Z�t�C��}��u�u�Ry�	�[2ա�'}�������� ��\3�����S�T%��X�m��&�_^彲�ӯ$Y`��1_a+X�i�lF*!��ܑ/`9�T1��ɼ~�\:n�طY'��/A$s��I�=P���]%J�'x��"n_db���ُ��$�n�I�̗��{h�����sӃ��������)�{ppe�m=�S�v�wKYL�b�! �:$dxs��#���`����v7�-^L�x'\����w\�E޻����M�
 ������f���oA��XV�|F.μӍ���qn���g�z|v�N%����,L�5���(Hï�^4��MU�Y��3<���ǰ���y8��P9E'����xͅ��F+��RGB���{�8q̱c�f�Ûv��0���f��oW �P�;.i�uk2.��i�ͮ)�4���+އ��H�<�*�&��ãl�=z��{��C�.'4�У���u�ss�_rD������կ/۽�c�z�^�ἅ'�����.��j��,���]�@��sy��T��_1��T�W8�������y����'��>>���;g���-�>�ڮ�R�񾠳'�X.�����>�g��vq�k�_3���iaK3n��ʬ���8m�p�ͷ���ۀ·:X��D��c�"e���e�-;V󹬌�ţ)���������D�Qb�y69���zPw����l�=ᖬ��Np����x��QM*S�غ�q���(�T�,3���#��fP�"���4���]��nˬ�Y���' �vWm9�/%���	ô�V�|7��#��:�n���"Ls1��x��s��$90E*�a*]P�Ԩ�ݪ�I�ZkG#�7>y�U��Nn��(3�t$�ru��&����|o�lTa�{��c�MY3	D$��t�c�oNd}�w^ӧ���E�\/_3[wa�x�,w�;��陾Y�J�u[��!��W�d���T32�;�L��c��a��fum�`֨�_Gؑ�W���;��}��K��k�X�%��C ���ʂ�4wrS"����ԛ�[�i��	�D]�����|���]�SW=��Fdiwv�1Z�Dd薍I�rrX�ju�s���>����#:^�iz����흥 O�-���[d�����i�js��r�DdZ��գx�d$N�Ɖţ[�J`�-�����#�ɚ���#1��[�昡`N�Cr� ��L�ۣ��o0�o���	���L�̺6�n�e[[�عϜ���Z].��8%y��Lrغ�#t=y\����{����AU;o���Ȃ��L6���ȶ$�{��c��9=y�Ε'ՐV��å:������{�G�|<��q��ga�]�ܙ�.eur텙i�+Yނ����ueq���ھ��ˬr޼Oq+��f^���
�	ݕ�Ns%�5W��fX����(�"WR�͐��0�� u��t����
�m�	���'}{YEK�<���%�
u�B��n�o�i"#�{:k�1j=�דn6�s��}���H���B&d����H).�B����P򺺰C����˭��?/S�;�P�r��n�-82�p@N���iu%�9Vc�Δ�V�K%�Q��`a)��u]��y���~��x#՟��W�d@�s_2.��m�b���]�Y��iT��^���R��-L���ʹ+J�|��,i+��u�\e���CM%���嗺�G������������={�뺭|5zd�UM�7��DE��V�IX�r��ٷ�w>�?L��t�C����{���4R0�2���&�{��n�ڗZj<o]��J��DVT�,�!Ř�w%7LΜr��Mpk�}��j�����;fjO1l��Smo]�)�Y��H������}�����
ܖ������l\���'/�1��e��Q��z�QŌ�=�,9]gc�Ť�h���ٗq�=��w���6�?}R��~�]O�˒��P��]0l>�`�a<�uDI�)9��#���)���ވ-�@t���
U7F�6%v�*�$����sß������w!����s�}���y/lV�l$g��Utp�=�h!�T̒��a��P^?��/�i�,j.�� iWol������tB��sT债�*��� ��V)Ы �P�p��>���Nw��r?<����J�we^��+\}a�#����~y>X(�H��~������˖*pbh@��`d�[�E	jm�c��J��tpb=�[���XE�!�{����FzI�VU_-{Ս������[��m=�_cQ��[�鄸Yۊ�l�l��]���j�eHk�_1������F��u�ۓS;R`z�a+V/v9Nve�UK�5��x<��t�p��,,��r�uL)Ώn�Wg��s�v�ў�^�\<�	G��M[�}$���9(;���=*�����Z3w�c{ڨ�K�X�d��{�R��q4�-�~���NC7G8.x�
^1�}�{G�{4��ðQ�7icϰ.�˦s.��:T�L�A([�mY5t����鮬9v��R�0�W1�f�^ʐ�[�[���P�)����ؤ�{m���0����E҇ap.��^ǣ�G�����j�о��-��;���&b�k�Gr��ʚ�D�i�d�x���s��ݶ=q���)+/��r�/DZ������J����A�lL|ftZ��DlKo��^,]s�U�m�)�hՉ�ܡ�{����R�-��T734�X�UŚ�<Q4��c��K��>��ye-�l�z�B��[�0N}��Y,��x�37~�rN��1�N�"��=#�<���/�Q1�^���o0̒s�*��g3���S�oC�q�wNԈ+��T�t��T0�j^�c�ܫ�����kjX6���G�7�$�<�<�����oSf ��m���Y	�e���a�����e�6�X�ر�,j�p�:�fМ�4/�%�uι�����L��x��T�:gD����K����2�;��щ+�[�����ܔ����'�y�)�B�*�̀����!(+�r���O]��s�Îr"ʼT���R�ȝI�%�^t�5c3�QF�M�#�d�At����`�a���ϫ9�[������I@�+QˊN���zIj=�F���cw�0ӣf	Bȋ�Ⱦ�K-����/�j!���፷��8���h���2��}��[���lWZ��	�[������iR%���J�fo;�]�5S�8���{@J�ᥗ����Kq�v-q�&lC�,�P�`�ᮐ ��z�E���:P+��J����%:�mC�2�o5����r�wA�*t�YC~�-\8B��c_]nr���Q�|���Jh�����l�;��9Ǡ�Uu��<�==Oo^���9`isu��b���|�SR����
�j������r��:ˈS�����Ls/����K��G��gi]�?[���v�7�s�eZ��tC<0s���nm����!�v��q�e�'a�Sw3V��gQ":`�Z�h܈Vo��]�V1���ϱ̠��;`�bU���%�>#A`t]�x������ϩ��K'A�Ⱥ��n�9�%+����-��i�7p� �vF��GtM�G_U��@�i�i�Nr�gBI�x����.Q��4���lJ �;s��|�"b�
����40P���;��gt�98����P���h�b�KE<T2�m�mQ���Ũmy�h��w��=)�Χs�&(���L=�'��o]P��e�\l�N��5�@!�(=���������3��Q^B�v; ��+����rX3�.��|�=U��@'>$db([˽=�ǆ^�׶�r��gp4��P���d��s�D�H�7:�lly��efp�������ן�Nb�Y���$�<��Qۼ�>}����f�t������g��$~�N�NV^�
��Ӻ\�'72<�8�{��tŚ�'�P�˧�Wb�L�io�Qw5���5i�%�N9��Ԫuع�=|��ԭݘjH�d����	)�K���,�g�o��[��j�ه�V:����'��k� ���_eQzN����r�R�uZ�]{�����;:��2v\�[]m��w���;�{w<��8"�9����+FLF��N�D�'������{c��g��0g��2}{o��]>␭��^�hC����2��2w�y�4x/vu�N�:��ܕE<J?h�u�"���I���.�j.m�4[�#PR��5.�%�f�,���eʺ�K;^�n�@����rM<F����b�o0Q9t��^Ew�c�x]�đ6�mu�t4+��1g�����~F����;�e�M�#��ڐwC�	l��u��_q2�38v�CI1�u�w'1*R�b&9v$��w8���ו�0�fr~�A����uq�_��լ�x�W_�](��B�)���<��uG���6�c�f-_�VWq}o� �
/C�Ѽa�+Nog&�{�fi��H,�:h����B�c;Sq2�rk0�����N�����=}N��yA|���	!V��p�<�wx���S��N܆e��5���ݺ�L&3)��w���y���vf�3�p��p��K�=��2O���\,1��D��M��v&��@�������'g�,{|qQ�I����37��|�	�+�-Bnp���%Vj�W;4�d��.��EÓI)�PIb�<�b���YeЁ�oL�����,�#��/�t��\�=���8���X�q����8>U/4�o�[y')�ִ��ӷϡ]�)�%'R�]�;utN�,2]�`���.fXpqa6E���ʧ��E��5��eh`��@����sj�6��Nl��3�g���:��)��+4��ͣ+ɬs.� X�4�����o�+j������#)��Pؗe�_O�]���9JQ}O��1@a��Hs9-��D2�u��z�����6��y}Q�!�W�OS)��yѐ��v-�����9%e��ж�%��A`	՝`i�6���cUEN3�;��iP������hT�E&����m��J��PN���-^@��K�I��=�\ْ�[�|[�X�9a¹V��_�A�q]5��QC,��TЈ������J[R�%�����u"k����l�,@�ǌ���n����PV��,_�����r��ص�5�M����|����t oV�We�8��}z�-�:�8���핞s��3�CƐ��ǂ��!��8�ޣ��rM<l��s��`�z��x�����P�Lz�b{۾F�[�*sD�� �Z���YP|��˃���t�Os�C�@��bھy]��j��B���k���c���_*'��|go�$gj��+i4`Ng��d��7�#*�]*ͱ���#�m�G�H�1 �r�-L��nf�r╴u:F�[��V��-�؂��']̉�޼p�iuصð!�f����Jޫ鰽�[\�����cǏ��fe��3��������O���ګ�Og����f�K��aG�9�q�.��h�V�mܚ
�װfa(P}��8��n�rϖ�4�K��,o\�����^h�g�*O��`!:�g�y�����>�N��{;Hx�/�cQ�50>k�F�Pgw�·�Z�<
ody�̠ �&��Hr�}t�8^SYV6+���v���7��F�W�j�����-#��{M+�VV��:��^��[�cÔ}|a��BIښ����_E�3�gJ�@�wA;��c$��B_�@@����ҹ����bY�V�`��9B�[99�A�G�2�Ԥ�=4g�]u�H�R��bRo@���p3�7C�<o�b���4�x�-T�Oދ���#���v{N�9p��L���>�j��ڶa
(����r���� ���V%�YwG�ŀe�sr�nb}�Ei����n�V�z���R!��<ͩL�؝��wf��#��뇾�{���ZWu���2aqh~'.l�y�g��6��-�{޵�Go�Tt��D��)3�)�{�'� ^Zk�tE�e�K{�,�yn���U�3�r�I;��Z���F �ŧyY�6��k�>r��E"��}Y��,���`�[�J�F���Z��H���*�֬DeC��r�]=���^���q�w
�E���n���|%�m��i,[H�����6�k��o5Iz��K{�����j4ＫZ��E�!��F[���W+Z�7V���-�pZԽ�|�BA8w%Ƨ�$��Ɯn���I��lu�������+��p{�?E���qG�sf����3y�ʛ�D~om��H�����j��%��r>�Ժ�6��Z�aé��ݖw��W�R��+x������y�7�N�{�2�tc^��Y��`�s��g��h^�n[�/Z%u3NJ0+���k��#�w��TJ3��L��e�m����]����/^��6z�-�_]O�E������}�����}�}��G���b�AR������].4�u
���G&�X�+�b)�Z�ؠJʘ�Ø�I*�*�K���<�h�"���/8�Y��;7�f�����M�M;�w�v��K�j����3�Ѵ+�2�uq���1����}A��ي���k��ޗ����^���GN����3Q�gyRX��[���F]h��"�E�]�u��m�u�[6��ש�j�ǈV��K���wr=&�R����R�6���/��I�l(un_����|<�=WC��t��};{���v0�����oAƸw�o������/����C[���gH��m��JF�o���i;T3$e�o�^*���:���roc+�+A%FZr�j9���r��N�3�n��M0��7��p��r��-T��!�����Y6���w�O�;��hQ���5��ؼ��]��{>�a������b���Gh��ݴn<V��W�9B�kMӽ�m���f�kM�R�F�4�љ��� f�X�G�y�ת�Z~�7Gs��l����r���mm��W�)�R�ZPL՛P�̘���o]��Xy��3��W �L�:�^$y�o��s ��3X���cӯo��̩��رKz�����^������ܩi^����%+��5y�~T�a
_��*�w^�JbJb��f� 6noV1s�k7��H�.λ�D��9�`�B�mX�3�ibcO6	\���D�-����(S�jt+�o��r��by_�wh�G>a�wx�@�Ԩ�:���׈R;��s��w�.����t�0ک�DhA��v�Q"�=��LZ�O^^�^A���)�,;b�:�.�w.Ioi�b�e��ptw.c�d��FQFXl�ۿ8Z��P�I<<6b�Q�h9����J�o�`���q��6�I�]�d��YT�b�}S"����R9��Lu�[�3%��M�c�.g<��=�h��}�����:��[P�i���S"u��(���ؒy8�f%=$�XQ;�^�����[_mev�xB��c��vS�H]��<N-��+�Ex{H��R͉��a���	���vZp�^ݧ�^'�?�<|r����>A�Z>�ﳆ�i�C�0�?;���*x텵��ds�ɷ��3̃zUN�K���P��v����OR�>@���+*vuq)s� ����2���NoɼR�5�}�a�se	�ix�]^=}؇vi�/�Zi[}z�Sܽf,����m�-룭�`�3k\�r`��s�f^$���9!OSKjR��y]i��,Wo�s��!v�sьǳ�"3 )f�TZ��g��۾XVěC�z�Y�\C����|S���L�z�oS�޾逺.�\�V(��."�y�WBك t�%����Щv�X˩PW%�2�O�ʌ� �e�^�摮���w��ۨ���on)��\��p��Ƕ�uk�`��=�kB���d�AI�[�V3}'���4����J(���d���dC�{	�jx��坕{��Q�E�o{31����Ĥ��S�K��znJ�����܌Xhh��Ġ�sĚ�];�n�ddvA�]�2b��h�$�i���a�oxE�6������47i�+.��3R���ą&��=X�C���a����ܹ�a�'C]�lP��̋�f�,V�E�so�ov�ˢ鷏v}5��5��D�2A�V���{ɀŹFc.gV��l5�bnnb�T�������Y�x�9|�NރVt�m�a}�
mX���V�>�W��Qb�7K�]�,���T]����V�nQ��5�>*:�T�)&�73���Ϧ���C�p�cg;&�t�D�7#�]��J�WռiiD�~�ݗ/��:��4}2��EoN�'�5VX��ք�*ܑgTp#�z��1C��4 ���ܵ,}��U>b�fC�]X�.U�(!���<=7G'���X�X��۽����A4MM-�)��m1g:2��>��N92���広WیӬLl)�p�"��.<�n��m>{,Z�����͠��Jĳ�ror+�y�Q���辷�k|�:�i��f�R<�uDX٘Aze��۰5gB��S��Ê{f�/P.[|&���,�j���&��-	�Fk^��БԸ0͵)91יuջif��IF����;. �o#9����SU�:�����
P��0��k��la�It�g��\]�H�n�!ywt�,t��
��n,�7>��s�C��y�v��
.aЋ:����3NL��7�ߊ�F.y�ܾX�&Y��9xl�<���F�W�S��i6�"�A��K��h`�Q�5{�����1�뺼7>T�pW+�����b��.�����<���5Ю�˰bѡ������������/oU�s�_���6����p����������瑾F@e�ݓ��8��2�E
��6f����&��2��:�*�S�]�.���2�0G�Q-�`O3�k�1�8z&;���(VM$�!x{�����vW0��:m3Zw���KH���f>O���b�QNg!*��X�/�뫾�>r����Q�\�i3�Z�<vÜ�U�p������{N\�}��
�-�o�-6O>��f��gw
Z���f��w�|%��WfU�4P�bW^`��K�t���sP�O��6�НkA����MnSm^����v���0����1SI�
w�&`+Ko}���s�'A�k�=@�r�X�Q
c�N+4K�B�.�Mޘ-%a
L�����;�<f�,^v��J6^l��4�z���WgrgVf��WwDB�k��sq^��|[�s"8[�"do~>o�S.��]��$A�Z:�YS-
����� 43�eYXA��فNC����?'aa��:6%(�-*�)�W;A�̕����3
��rA15�H-q\ZYAj3M���/a>�}�9Rh�\x�=����νϻ�k�+񬫎�˴�a�[G�ɲ���Z��|�T5k[��׶;��ce�ƻ�	�7;��XD�_��hcb�ֲ:���PV��/,�����Ǡ|&����r��K,��&k)%6�{e���.[�h�g5��&��.��<Qn�c턹vr��r��h�[�ss� *�HJv����V��^g����6�g|<�i��^�fp�|�C�ѳsk��--�R����HK߂j`�q!Υ,`�@P�U>ʈe�d6������U�%�U�I��)ld�y65�wg�ʉۭ�{��y�%=��R(L�WM�3��,�E(ݍ����A뾱eXb��qGh����6�|jga��F◦B��r�*�F����/jbř�:���P������1h5�ye���T)�%��y�3x7o�W֎�ξ�"�X�B�b7N�Z��t�_l�^T]+��1=��;���<�Kz-cvk�e��;V����lL���q9�\�dK��F�8�}��.�@,�j��%�op���V�=�mFb4]�t��n1ڎ�*�!��ר>�7�-Ǜᾷƍ����]�� ���vl�穃�	7�&�c3ms�)L1��4��ᖬh��$��잠縍���je�3��`�S8��1�Ą (Q�͸���eM�P�Zav"�
y��u���*�Y����r�.w-��s*�嗋p�83+�MxmlА���v�p��D=�3����o��N<*�Wt�G��]�^'ҭ���$�(��z�*;��L[=5H��T���k�n[��֤�rd��aV�u���>٧3�Щ⊹Pt�����#�bz�Ћ�ڇ_3l纳;#�Ǖ�;��UDpئ��L��m0�&5�lW�Mu'�;��Į���=M�fI��Sx̌Pכ3r�l��V�t�Y¯e܎\��4T퓞��l0x��ʰh婧Ψ�����JT�c �Q;73��\�6;J>�ь|���m���K��Q%!\ֵ��X��^��H�#a!��\꒾3��E�k>Ëa�/E�N)]g
amkU��8��yJ�� x������Q6��ۏG�Ç�����Mf!g�	����N�,�t4RLަ5����f��JPw#pu�k���R1��\��b��<��s3�Ac�8ұ���E�Wy1�:��8Tܗ���gf[�Ąp�v������](e�D0��e���漄��{��t���ĉ�*��̽���`�ʄ��9����ՙ�_�+�^�y)�v�L��ݺڤ��$�k��ڏf �֪+y>���meɎ�Ҝ�݉V�p viX1��7��ŭ�o�ͬ�E��wgZ@�+� Y���iX0U�\�{��iWL����P���c*&�!�}��+��ᕕBM��ܜ귫�m����w1���BZ�y�����A�����C��bޙ�'�`~����$�Vn)j��ξ�ij�ݙ�Gtػh٣ˆ1�b�hP�}-8���6f`����F�3�:��f�R���dfq�W. f�EN�e���!Fn[�Ǉe[�z���m�%H�ƨ_ �q-������\YǦ�kMvu���[�R����o�Cn�nS���Ԇ��ۜ�t��h03>�[�o��I�]��`�ӽw��ݦ�,Jb�����r7C�Ӗ�hfv*_W�������D4e�:��uՅq6���"$�D�(f�E^�hFt��QxШ���)+�R5��y�R�f��ն�n�:�*E��Y�2��I��n��uܿH���=��D�>�G�,�Ë���L[���7�.�K���{H���ٗ�9�����ÙA^�%0��hdLY5t��T��f������Hfd���(�٩?0�L���<���2��8yn��D���n�!Ty'�}�(�F��.�S��{^FG+�}f\���i!!wcSAߦ���gO�=�`!�������Χ��_�����v��d��U���X����է��	P�#�B�����*�{��J��`ʶ��d> ��t�=���o�C��z/��s�Gh�v;;o����7x�7Iu7�i�y�)�W�C�krٔ�r��⬷HD��L��v%�����fP<k�-o� ҙx�<��.)x� L[|`Ne�G��y%XY���(���9@�·�.¬�NI�{p΍Hv��ЮiKb��c���T�+�E��i]N�������L�Çe�����;:s�G�r�\[�{C��X�r����O��5�\�;ğ\�����!@�Xu�����z���3{{PJ��OS�t��r����x������z<��Z=�x�06�˾oJ#�Cw��˫S��3�^C�9�׮��}�l�ih��41�i�J��f���mg^7`�tT�[]ZE�5�k�H�F���W{��fLcB
���Nr�F�h�%�%B�ֹ";��'���i;�w;�Y
5��A�DMu��.�r�.Ҡ�c��[����R� eS&�:���0�����t��:��t��]'x�+�ܝ>wI�w�*&�Ztb;.*moQ�,�4���oX����F(�m���ܽr�n־J��kYni��2��p䋼���.�S���+�I1�1���T�\��yj�6Ă�x؃���A�f��rWO�LS��q�g��B��@����p���$	#���@=�����"3����&����D�f�7u�/5��9.[����º�x�e�e��́�k���5yR�m!L4P�6�1�4e�b���gM�[��b�Q���2�〄_=]|�V�Ne���
ڪ v����J�q1gm��;�{)��ܹ�B8!y}�m�Px�U��������4&U�κ�#�7��z�"��I�k�4i�{�/��$QyeEw�J����-�9�U��u�p������kqzˍ�r5|�黪�A
�v��bE��b��ئ�ӿl>�D��&�v,���.&�y9rɷxƼB�[�?
�ᘭ��]�0�E�$8���:���nFFzoVP�.���ǺC3X��.)��=��.��;��,XhR�̢��qn��:%@o^�c38ؐ7JoD/&�
�	��f������r����i���hY]�: �Wdё�S�R�Ͱ_�w >a-��?��$kA5(���,�+�ÌJT��H�B"�W.�ˢ�.�VV�|y�)�htTZr�Dt��޼���M�Ks�d�;��LB:�a�)�W�����ڵ�����_h$�>���tyx������8׃ԱQa�מ����|}����k#K�:��N��k*fq�L9:޵`��d}�7�]X�f��B7י ��`��7ʹ��ZP{-Px���4e��f���p��x�Muhሜ}�S�׃r����T����.��]Jf+t��{M������/�{�������]���12�]�m�=Z	+�xe��i�Um��Rm�J�/nr���9O�*b�O�gHWU�D
.�\sm�B��|b�5�&���3f4�ih��_l�:k�6w��}'�}�:`�(���ի;<�Wǭ�)K.Q�����gC����C��GP��v�/$)��n�ZP{�'V0�mP��̨yFw4+��5q	��a
Г!{�q��cM&3)A��a6�X��u�i�(wvP�n���0K�pH�R8kj��Hl׽m]��cÞ���f�R�$�8�sgtNol^��G���{wt^�c�{��[��6P9�X�,�z#lᕠ��/���ݡC�b���:{B�me�G{\8| :F}{�z{�c}C(̦Jpe~���۾�Ez��Eu�9�n2k���8�!�Uuްf1�R�_VN	O����V&�Yr;�Z,5N�oy��l�ưv��ﯗ����߅��n�s�V}��'��V��+���������֐�}�n�=�ÅZ���̒kw'X�dq�[���I�IU��=���6�<��9C��O��hǓ�D�����öʻ��a���0�}��$.�R����h�t)�K��zn�Sݢ#��jpk0�	�f��6�Z��Ő,��u�o��b�����i���15I3��ze��n���T�s�5e����w��ji[	C�c�
���ڴ�_�8���L��Y����jv'���q[�W����ܦ�Ć]�)�<�����a�)3#y�n=�i��Z'V��`�ʐs��djZ-�Z�����3�T���X��:y.��e���b���3F�Y1B*|^e��n�ىn����6�к�F�2� K�M���C�+���w�a�|f�v��zq"a�~�4T����e��ʓ̉|B1g8��k�qJ��@p'���!�--Y��.��L�,W>[�����ȰM�2��m�F�s�4���;��?5{J>�7ޙ�p`u!P�w,�G=��'"m�R5t����8""�����V^�k�P\͗���83m/o�X����m��h�5��,�Ku���~(=���pY��w�Ʈ�By�{�zy�Xe�XT�zoEs�Q�T�g�N�B��j[��.�d��wI��0݋7�U��02|�%ܺN
��8������䋷ؒ+�Q9�r{��Ru�|*񒣥F-W��,��"��&~��  }3xu�klI!�Y͸���(��f̢Ӷ�c��U��dr��;���)9�݆fڬ#�Gsm,8,�m�٨�+�޷1��l[+"�� ��nE�^]�5ff��ǭ-�f��ͫm�N۬��mcN;�����m���[E���ղ�Z[k�Bis�p���y��m�f�e�a���vV���Ye�[�őm���Ͷ��5���jO{	z���F��e����8���ֵV��N�鷝�ye�!nł��Sm�m��\zv$�È";nܖed�7kks4��q{���Cd�7��<��b���C0��֭m��$}ws�^t~�+���Lt��qcص�9��鞣%�����97!�%&K�c�S�l4�$�n
u�L�y �f��_|y�����L���&v������`�H_��p�*:�J�R���gG4/��O���#�6N�ywM]v���e-�dP_w:�-j�{Q%�j��g||��V,!]oU�=���َo�i���05�A�3S&r���c�;hW���;��ǸW�<���y9�G������5�ԫ+o��˥��?yՈ=�$kͪ�c�*t�)nl�,r���z�Q{@�����Y����{_������M�?U�,6j��-������"v���$���ptC���g��9=3�[;0~���n!�c�]VOmnX�Es<�^G=���\�g�c�îK�'Tl � =�� )U�}�X��u$ ĶH�qB�Vb��<�������z�D3�|z���}>"���+xzڥ6�����֍E����}֕)-��P�U���h�C�R W�n��Nr��4��t����Yc܋�7WoU��2n��O��L?����*υxd��S����W#��H�]R�14�HW{{��)@б�&��^��
n�y����1R�	9�</��n�۾}[���J�;]e��4�-�`u<��m`ܾYI7�ﺱ����c�	���Lt�κZ�H��z�ձ���}܈�!{�p�ej��[�̥���ڕ�;	u���ԃy^�̨����xK��K�[
�����o{k�^5L�Eyv�^I�7s/�=�.��B� ��X��b,hY�Ld��x컌N�h�
M�Q��UIښ*��YY��Chq�m�C�(؀�6���|;%U��k����b2%�� ٭�iGO�<�71���-UeB���u@L���0�>Qn�����Z�
z��x�;�!�r���V;��_�Y�w��I�8�%Y�(Wi���C��4��*��N�M�T�h���N�ޢ���'���I��y�&Hs3M�@p�#@�2�����u�p<8��)K��oC��Q�9�B�|�<���:����4L�V KF���;Z��/X��zFc[�L�=F���<-�m�W޷[~@ �ׁ�w�<3�n	����v��]��_u��px��W�sn�V����ѧ�������)YT�XK�Xodin���#~^��IRO��o�P���t����,� �p�k@u�-I-^�G��.�p6��O��#���Nn�}��BWة Nc8t4F�ﱩ|��S�"�4_xT�?T=G���n�_�Z=X������`w
��JIo�=��\��˄Q��B��L��.b ��c�{�+�{t�7��,��ɘyp��aoNs�l�c��]��Wj����W��0N��vyoJq����A��U�ђ�$�x������ܣfe�{KD�F���҈s����P�8�֖��%b�W�|ɫ�6�ז�.s�9���R�,{`�~t����T�l೎������~ɂ�s5\kç��1��^ewT���Һ7�ê����詎8�EE��*�)lm�ڸk!־�X��T3�B<p����hեh����m*��\7�o���>�\/��f��ה/��O�zQe{}�����՝��u�,`3klƗL9�&����*4)z3��V3�����51��s6��z�A1�r�ʴ����@�T'�/C�ˋR�|�僒���sZ��!��'�9!�н��x"x{��-�H�Йةs��{R�mg�������^��H���Tl
��m��?6q���)�LL�/����ԏ�OZ��z���N��rl)�G0~��=�P����1��F�5��y����=�
e�m��;�v�nd�n��&��\^Sַ$G�
�ƍ ����T��/��x�]Ζ���8ڛ�v�qd�P��jW�����W9ܙ���ʊ���>U��)�����]P�4�Pͭ%-�6 |"�q[�:r�9r�|�ddh0�2�o"ݙ�6�8�7�l"� �;���иk���g�'��jL�Tc�9�jG�sS��}	�I�Q�E}�~���^�E� P�Ḃ)��V�@�&x?�ɊuMv߆��Y-�@�~\�C���˜�q�aB�U�#��v�I?r�t�-�^��<X�/�=������{C�oώ��ʦc����'r�8��]��D��F�z��U�|u�g��C;X��d1��RuuW����K��Us�x������2}�Wf�{���w��"�j�'�Z����y���yԼɞ�V��wyO��_Z���,�Bk��+ŏ˯��\�U���R��S:@�eH`�nz�������=e?'�א��5��Δ����Z�y]R��׆i��K����ub+hc׼����lD�su��~tM���g�P��Hxl��:U}�㼽��.�����=Eק7ݧ~�<�oY�A�}�Ȟ⾫Üj�̨K�4��-ꗳnh�����ln�7�"��f1�J����.y��h�XSʋ4�LF���T,u�L�>���kF��)AbՀ);*9�t���}��_��u֏�6y"�i����-���$c�ʙG(�]��.��a8�Hb�>|���J�Hu.�h�F�c��yI��p�W�BŖ���e��O��޸0gV����@ȭ�Wgi�J�9��m���F���OQs�DK�צ�{+�0�e�{ֈw]�8��x�T�#Om+k�P��)t���qS*�A��֢cp|��p��a�;��o���~t�U?H�$x��@�0�y��2�.��ٽ��(e�K��q���l�B�.�O��?F�ȫ�Fuy_u�w���=-(��ql�e�Fm��8?��B�a��:�dJ�8����:�!��b{��ϓź��z��H�ޏG��~F-L�Rч���b�r�:�W��aHͯ&_�E�F뵊�mr§dK���tvB]L4=ʼM��|=�RI���ٌ�Pnٞz��g�F�Jq�Gt�Jn޼FeD�&cOЙ3�����>���"�����h�����W�5{�`�\�s��=l��
�fウ�ZK���9��^�{bHׅ�̀�^����
>}S9I'���=���x 
Y^�^���rV>y�y�u�O�o�k�D�P5��~��2b����n�$�yãj�T3���E��	�zP����Ͻ���W�~�;��k
f��O^\�R"�KNFpTԩ^dө�E�u�g�e6J��E3�e�7��wq�F�o3�3m�t���3o����rm��Z�=���\<)%�2[c^�}{���ob�;�Mu���[V���#K������wrW>y��H�֗wCͻ���xa9�+�/�p���V]>@{qp�� ��<EO���f��w�+7ܪ��X7R?T<Wu:��aPB���OO�C����vU���'�2�Ob�q�e�Tl���LdS�w>Go���kk�p$����҉\��Hh��nZ �i����mz�=��V|(��W��I
��a��ͫ�,��Ed�.d�r\�m'��R+}3�bn��,ڋ�U	��>�~��3QҾ��K������ץ0tp�iK��']x�{�,��{:� �bx�Z ������5���1��|;���B϶��(����0��Ƿi(]�W�qT>���x�T���3<�vH&����U�+��{	G�x��c���� �DS^>>���!���MƆO��])IR��@{��4�Ćҵ�T�
��XU۾���yV[����u\>��_���y��"x��o�Z���JE
��e�1U��l5����Ihbk�(��Қ�p@�А@L��sW3� ���3孟�H`��3s��C�PХ�i{���Z�h����W+FS����:�:$�)֩1�5�j�6�y�jM�W��>úu��@��.�j���i�践���]�길�y�/:\�Zrn|tH��`��ax��΢��!����̉<9+�ի/��4yΥ�x�#|��w��{��X�η^���Nj���P�pHOm.%X�+�����n��M֦���w�S�F�͇OU�&[pp�g�H��Y��6������]�r�cT&*z���[�K�V�oMP3��+tW������[����|������e���e��<��=�X�!���:�����W{^N�b������7u݊>{֜˱ �)���HgT�.�T:�jU;w�R��lכ.���cZuB����t_�D>	f!�lӪ����n���-D����:�'��Þ�Dxf_zX���h迧c\jW��~	pa�����]�u����I�^����^�����b��Z<�E+.crF�-Ә|�{�9:g.�b���.��opV/�e1V"Q�O��S
�����a��밵p�::���sa��F澥���/݇1��}+��J�85�NydY��.4A���*b��R�0WYn޻�`=�kϧ�v*��=��Ƣ���?V��u�0�2�����^�Z:W�Y��K����#���o��ZՃTۥՒa��z��z�[��]�	�����=��Y���E���ܭ�ng��sm��R�aX�K�[���홴-򽻻FO�J�ݶ�ܯ_p��Z���F6t����ݧ�m�j]o��Iɻž�F��t۷�|���u��K� C��G��b-�S�tv�K8Kڜ|�y�OS���Y3�?.�g{���g����g�'��R�- >�>��O�g�Hڼå9ԵL��X�S��u��(F�)��۽��g���]���mԗ��{}BN�{����(;�Z'��u�}���ЏC�T��.6q�:�M���JNr����;1"+|HC��4R>���j����!t3��[�� ����s�Vljw �w��{���:/܀�*WfU3¼�[�a��Y��2�8f�;u0�զj�K�3��udjo&+���ڭ%�0r�KvW����Dd�I��	�c�E�/jV��mh�x(��+G��y~��U��O��_��#�20����9Z�=��B���A8\��y��G�kƪ���^���+n����Wf	^��p���,���ל�"#���>����z�����O��V�|���8����w��s�צ+p��	�qHbO.iт����'��w�ʚ�*V$��8E�H$Wnr�r;�}O�U�ѝȼ26�fUݧ�y��ْ�˛�g��~��i��Lj=���Or���P��:��m,�ϣ���yh�~
�=إ[��[�	������}׹�C�c��LR�y;4�ň�1Mr;-xu�(��}�3�`��ʵV�~Qv䃓7����m��m�"��Ts�������tҽ3��
�i�|�__s��.��Ou��'�{:6����R���{~�v�w(v�^3��Ȟ��ԫq����6�7�9�u�G�~k����Ȼ���}Egp��be�m=����4U��OH
���::ȥ^���S�M�㙼:�8	:�ru�)���4�.!3lz�ҬNu!��4��Z��}��f���\�W������{�jx��v⁏-=}�/���	�l�x�V\v�M�6��	�5���o^%6���
�*{Jj�j���7���U��>�j�·�������S�f����VW'R/=�wu//&x��d{ׅ��O�]�J�{~+E����|絁ץ���q�>�gl��E�9�dTVk����7�b���7�}���Z-��+�\:B]��Rˋ�V��Ү҅��åȓΜ�_`?!r�t�=�����y�c�hP�v�{ζT\R�ձU��F!:nWw,���;,��G$�q�n�pL�寴�u�6Et|�.z������To��*��&�g#nz�-w{b�:b��Wh���W�Lb�e7�1ڶ�w�Ds�\ɜr� �f����Y������4�!�����t3�I�iߩ����m�_09�C�@�{�+�͐a�X4h1��
���P�R}u;�n�Q�R�A������?�A�pQ3�?�K�~�V ��iSO>�;���Y+������.$��xkt|b� ��u�i�5����b�\3�?W�W.�\�����{�����N����=�o<U�kp��N�|�ug�_O<V��+�����MpM�޿u�t�����p�ѵ�WZ'�ߕ���6T�핏���@i�K�ݹ���q�tK�[aQ��S��<Wu;�,:��.��}>�H���WP�=��[�ۓU�n)U��zK�i��uA��r�Ȋva��;}6�;B.ҐUW+~���}��,�w*�:N^{��b�H����C�Q��I
��aζ�9P곇��b��׽�,l�	�g�K�7��/?{���m��i{JiV����h�Խ�d�v_�!A�߻�^��6'�1aՒvv��ecִj)����s'� uF�Y�-�Q�=�=_*�bf�g���mZFI�������d�&\��Y�W��C�$�
�跹9o�$:5d-|�#+w0��G� �������#�[��c9}�n�e��U�h-��kqv�����������F���U��0�p����r'�,�)���\ߑ+�z�[�{\��oF�n[ͽB5�еyܐ��8�`J�#�� N�=�� nV��(A;Ǝ�zi��HU���i�E�	<�_Zu��=����C��s�)<�!�]�.�³uu8�{�y:��N���>���4:+9Gr�9�����.\�A2�ޥ����0旰+��n�92Gn�%��k�@��Mu�p_�L��Ad���ܛҔ�L�V�}{z�`f�u�7���Lʐa�����g�d/d�N��\ Q����_h �&��ݵ-4A�ۺl�s�LǷ[����@�)�r�{�����<& j����to��>�z���Y�&���E{J��RZ�`���v�2b���o�]�]��2�q�#V�IKo��!��oY�����r<٣���$�«qs����e
�s�3-Po�U�8���
AK]�n���#���e�X�����s�M^6���\�>k�v��+fm�+��1���Y����Å�{eo�9�vtE�4p�2�����@x���+W��v5b0��&3wRxR�rn���"E�<����o�-̗�c����ը�l�N�+���DHrZ;���L7�8�Ƌ�1�BޖOz���[�#�k0*Τ�����G*�u�=���p)����Pw�����B__ϗV�5�jlG�:������XY�ΐ����lla�����)�5X�"�wjژY�A�\�T���l=Oj=��Ww�wj�+���K�����|���XC��_�>q/��t��eX.Y.;}f�x�10�_�����>��4��+s^s��j�Y�2-֦1VE0�P�k*=��ߠ�[٢=�/.Ml�#�D������9ɔ�����o��:��n:j�u��<z��ad��u��iv/�X�]�l�i�~X�KF�B^��Lz�p��g���0��ѴcZ�I�N�M��/�� �^�q��j�V�y�Ş���Ǐo���C@�)��q��Z@e.�׶�NRa�ȷ����]�fO\�廆�ב������$̋-�i<����`�=�)i�'3���9�Ԝ��e��r�Ձ�7@&Z:���%�*�h�&ڜ���#J��x�f��dٴ���z�R���ے�Z+�35�O�U[b��)����ȓ�Ӡ�7Ժ��JY�˔1(p�z�H���dPw��F!�މ16hBr�S������q���R��n�S*Pfľ9�_ʤ���V�]�W%*�[�/����fm����>�����ϯ����8��ͥf���Ks�,�f��m�ř�e�h��fv''Xrՙ����i<�����]�͵�@��h��&�flk�ܖ͖��#���8W��iq��k4�#���v���Y�����m��o'�͛6�-�9�8�Yi�'9Yy���퉦�8��SMih����a�)�e��Ղq�e��3Cm���B:$�rfE�ie��:�\DKK�H�{Z��˴�5��n"^׽���,���iD��1ge��:m��:�"�JR�v�f奅Y�9�Yi,�	Φ�i�B{im.fC�c�n���&Z��L����8��nm�^��&�p':�PI:G�X�#�$��r ��9Br�l֦ے\�3AaY	�ђ��D�E���b۴]�e�k�Q������Drm��vm1\e�C��Ԣɬ���V�H��Y؇w��y����l��M������уwFn��MQ��)X�[k�s r��Y�{�����c/ �{����xls!�{��j�)�kv�Me��ƅ�w{�e=:�����c�m���������+�{��~/.����y�⼻����Wͻ���~;�����VY������w|U�W�����/�v]羚.�V��������u�u�������>;���[��6ꆻ~5׺��#f�����w����Y�wy{�?~���|u�ۿ�����_������t����e_���2���^=���W��e���|U�eߟ5�_���yW�󭼫�`h����+#�Q�"�>k=4h�sΊ��+�t���_ߞ��W�ם�]�~����ۿ?7�_ŝ�������T]�VY�;����?u�u�>~{����������wa����;�����Q����W����$�����{�O����j�z��W۾+�_���՝���yߵ���Y|]_>����������{���^^w�?���w~��Y�_���߾��J��+;��M|@��A�y�B>,�}�W�}#��C�}�:�z}ޫ�9O1�A�n���m�W��é�߮�|]�2~�?}��1��c��H����*;}}:�w���������^W�����������_}��Wү�������;����D<M���"{��v+z��t8�x^we~��=���ߺ�:�w�|u���׭��ם�we����_�w�@���!p�"��O�*&�}}>��}����;�����wgŗ~_��W�W��a�Jy[�GTيӔ��֫�6�QqB>���7� ��$DE""�Z��N��:��ߞ��ʼ��_�y�u�W�O�|^\�u�}�_�;�����W�w}*�Y߮�������]����|����AF�Nq�k'��1����_k.���~߿~�;�݇w������ׇQ�_���w�W�t��5|��/���꿿�>_K����x��:�/������w�Yw��5ߪ�����\ �����K�)c�檓�q�|�g���W��������.Ϯ�߻+�v���W�?}��_����/�����wgDt<_`��A }�f��|���G!��TRX�W櫇�b��>��kA�A��C�QZ��*�ߨ��7���E��^][�����߾�:�,�����|w��wyV>�����X_�쟚�+˿U������u����:/���������;�ݿ��ϕ����x_���_X�"�Q���X��ڱ�h~	�1N��>}@I[��r�5e9��X���B�މ.��Yu�Ư�eM;�f����*��v�8�Ġ����ut�R�a�9Zy��	�W=9���=\L�+�K9��;��gU9��-�ԡ������0��CC<y�J7�BM�n�h����������X~���}@1\�����Y߿���W�.���z�.�un$}�ЄDxAK�D��G���ܫ���~��󿿟=���ڼ�����Օ�Up�������;��{��l��b����?n�����?>{��:�.�ۼ��W�����u�W�}���ϵ�_�W����~{���{�������w㯵���/����ۻ�"LU��Fg�쌬��vh�,B�~����V]������]��]�yyߋ�۾*�Y�u���ϗ����_���_|]Y����_��}��w���γ�����@x}�K?F���������㱷Ǵ���+73o�#D|G���E#�u�}�����������߽_�����^]���EDW��w����K���;/���_���,��{w������w>���w⳿]��⼻�[�[�����[���S��z-�E��G�G�$�B����<���޾*�?�������˯���������������������|U�=|vwm���g�=����?�"D} ��b	���Ѭ�DG��T�{	�!'1*b|2��gDD!}�,}C�M���W�e}_?=w����^wgo�Yq�����>U����wok���]�J�,�����M��������.1����!DW߇�w���1�|@W{�|�f��[�;����(H�(C�@����^��~/�|W����e�tw�߻�;����~o.��.�V_��=W���^^w�~u�U�Y�_����_��*�(�?Ϊ
�>�#�[c�����`���������j�~o��u��u�����߯���;��������]g}_[�˿����}_=����}_��}:�w����~~z�u�������}��*"�Ɏ'�����2���O!��.Ҩ�ٺ�ܷ�ÇЄD!C��}>��x��/��������W���e�����~��ʾ�|u��|ם���w^w�Ί�������t]��������__5�'��~����0f>!�g��^�N�Yͭ��DH���~������(1�����
��5S�_VW�~�>�x�LURw��u��Wŕ�YWy�u�W�}�n���.?U����W���;���=�{��R�Ӹ���o��������f=N�z�U���7����f���4z�L�B��Z����g�:��mom�;�3$�3���]P��t�ܗaBjqtՎ�VV,�I"�O;��8.�M'N�[�Xp�㶺�fn���Ļ�E�z�����.�]ԝ������y�t�,����,���b��ř!�/���kE+Wx�vM�R�e���Q\m5���}��
�ؗ����~�Ϥ�<�)����Mά#�d5��XK��:�=�p*�Z�
��K@���cX�d���|ny��r���[=��nk&��s��[iJv9|��fĪz��x8>��C~��<��\��U˦}صoW]n����G=��6}^5b�'��s�|X��1G��ܵ�5�t�4g�ֵv��j��`j�{������Y� �����ʉ���t�X����S�s�Hxl�`I�=��/T�:������g����}L��Z6�J�����OmrRÜj�*i����H�S����Yn��]�Ï�ћa�]����m���v�{ ��)�Q�k�u���1g�^n��|���#&�z�����	
_AF��S�5	�i�]NZf�y+$L�MOD�����%��}�@*�P�[��+��=�^a���{F'Q���U�v�K<(�7�z�?#�b��i���u� 	�o���Ф�菴kY^��'!��f�J����V��3uI�����AA��:z.�(�\4�k:C��3���t��lan�3�S"���c��z}<�k��rS����)��CJ�E��`��fjhۅ���P��>����z����d<}�� +� mY>7��C�sW㓓q���n��M�+�wtUckx����d�H�GN}z�8:'AWKED�xD�3�|��9Aܭ�
���7�	�|5X��E@=����o�ũ��o�(�rC>X�E�Q���DN���b[I�q�6]��*D���#���yh/s�֯��P��Wed���/+Ah[���77��i�i���N��7��)����3���]E��F��J"f�lې��}�p�X#a�!�N��E*kս����b��ז���m+7y� ���E��j�L�qi#���q��k0��r�nZ��ep����پy�y��V�b��/��y��#}�r�~��%������tB�[��ve>^:��/��	Z�\I��OV�JwZ�0�=�f��?���L]ح�F�@���ٯf��}���T�UL��S3\J�x��Tm�j�Ca�ܣrf�v�q\R(T����>x��e��'|o���~O���l��=�jN3a�6�o/)���[1Z�m�a�\�])���Wr��131�l���`]Y��{C���k�A��bx~����Q��	�Qd�||�AJf����S=ûݓ�C�s|GK:%>�^r�Z�)�̾	���/m�f������*��/�N�q��V���!�_r.SN�9�Go��v�2�B'%u��hW�	�3w�KU~iF���iͬf�HT�`sv�Wo�U�ȹm^f��u�sw��ݞ��{�K uZ4��5Oj(�6����8�=���O�?��{��	�5���=/��}�t3>���'�V�Z zio�L�h\A���1�z�pRjp*�;�9>华;��K�_��C�*r7���G��,ׁ�tvZb����ͨ�A
����ېx��5><,����G��)*C��ܨq�ZCK����ҁR)ו�aww�N�{h��SN�U�=�]�����v<�5 U�I��������׳>��l���mB}���KMg�0��B�	�叕E��<��P�03�
� ��� -��?^�.����Y���4���ޣ�p9����[�J�msW�%�/P�_��59� X�n�ػn�v<�k��0��.��tJb��6�~50�Um��g�J�[�`!(�{ܪ�CY�Μy`��*���=��>��D�=�s�ވ\-�nj]�̚ȼE�r�%�3�z��xf��K����{��&�U{�9զk���t{2�v�����z@]�c{;DY�:���Ȃ9�@=O�X�}�zk{Ż��1�x3�罐2�wr�9�]az��k�Z�f��s�o��5����,p�m������:o��v�I{/:��Tu�˄��u���S����$�{�fbSٴ8m���B�U���K}]�g.��,s^�7�I��^�*nT9���1i��FC�׸r�׽�kـ�^�ƴ?
��4f5Ы��4�pDG c���N��O}ĩ�0s>�_w��u��h躝�q�P[x$õ�������Ue���Q���xl�CO�A��mt~�ʳI�r�R���%�+��@�����j��(T��)��aB����)�Ҕ���u�.i�x 4/gi<�u��	�Ԏ{�O8�0���$��w�V��tҫ<�,�� ʮ�3i9���K(��޷1�z���G�N��]�Ƽ�Z8>��^N��ŝ�Ga�.�`=[ʇ�9ܳ�>Nz�K왷�%�S�~ب�Q�<:W���/� pC��{��I�uuf����'{ޢ����4ˋ�5�0�xW�Ϸ��^�D2S����:��/݅V����=�>�rS�z��d�����}Ë�Ò��~���%�v�*�s_�T�f��^ğs��8���-�S���;9���F�f%e0�5��^��x���'�f�o{��	�o�1i-o��B�h�w�fQ�ӀӀ�0Qc)��*N�_���u�/Ͻ�@�!��2�R��j��W<��#�`�z���93��1R���*��C$�g�2�[i�&s_����*���T��)|��R}a�b#�:��tR2N�c^����^Z�r���.� !�v$.���,W	u~pu��\�Q8'Zj�5ir����s3�W�'��^�F.��p�q]��<+���c�b�sN���(�^oh�6=��b�_1��U�.�B��#���V�u�V�Vd�����lN�د����΃�Wo�+Y���[��P#���0+�b^:���_�z�S�
�I��M��],��'�����_Z<�`�T(��q�+��(o�x��߽��Uv`s�Q�9��L�{�p���ֽ�0��;0Y�W&�f���տa�ְ|�<��	��x�1��S����������g��G�ج\j�vO'b�x�ŉ���:\������(Zsƫ[�0���弌�r6l�:ur��⧐�^�i�4oܾ�_��b�W�S�s�Hxm_�!,8*Q�W�]��f�v9Z�4�N�	丛	��A��1��=��/l:�)p{z�&ϐ0�&�Z�����5}e*(㇯]�E4�>�=z����:^�l0Ιa׏o��N�(˪C3��Y>��ug�,|���0�כ\��߾���,���󍹟E�?���yL��*���]�L\[�@+�T~��F�pE_oZ�a�U��skqI,��rI�`��1��HU�����ڧ:����h�J��::��zf$:�c�VI���{�+x`�(=�-8yW�u���?^�h���yA���Җ��M���-�ӏ���/�P�t��q��·�@ǻ+a�Q�w�0��N���X��g�wq�^+�v���}���(u�p���Ρ@k���|�.�q�j���b}��{��[�tͮ#Î��E=:e>ų�\�m+\��=ё�]a`pd� ��U�p��Z/�y+{�=]�������y��|9P���"@_w{��R�k�����G�Q�4�Z-�#^��{\�{�d/e����W�t.-4_�xp!�/���XI7ц���_U�Q�0zwQnZ�l�;����e�li1s�j�M���"1��3���a�X8ÈGE��<LY7M$��`�B�f���-�pzi����E�-���`�)kX��I��ж��1��FeuoN��js�sf���E8&X�-;{�u��.s�ǽ6D�Nx5�C���')jD�ڞ�b�ǷcY/�5�&�� ��}#�u�}Tp�)� �6 �/3,N���p�-���B����Z]#;\0,i��3�G�BY�4蓹d��������g^Ƭ���X�9>oP1.�	�Ƽ���r�nZ��X�W	�X����ǰm���s�S���O+��+\C���P���c�3.������AB����C�� ��u�yM@�,�fv��#�U{v��gޓ{�[>���_'2}�������|�����SÛ~�"���C@�Ȁ����\y1�9�_w޾�謝��]�^O�ζ?F��m����%�z�4}�|]�Ჱ��B��\�2)ه;����ͳ�"�wJ@
�+�nvB�=|�Iqq|u�#'*�Z$p��xo(��~p?��qBY�Ý�m\9�uY��o7u,+ڊ�5tV<�5�`�4�X��V�Z�ng<��Q�\�#]0gG�tr�c�B�H`e���m:~��v-|���4���k� 7�W��*� ͮ�)��i=�*����m�}��(!7Z{ΗI=����b�ZgCz�V� �����bИ�]i�����j�Gee	�~z:Ҽ��]���u��1���
���R� ~��������ʀ�$i��л�'o����C\��T��= �P��=ʋ��C�	��E(\�����>=�*�۳�O�}�����@�sɼgX�WVݢ�qx�K���ykvWe�|�[��_6��f��O=^;�<mSI��h];����}��ˤ��R�w~�����o�3u�����_����\�Wag|���ǁ�j�7�s~J�(Wi�{�7n�%Y�Q��d�~��YY���T�x9c턌�]�x�Ǽ��_��Q��W ��s��V����[�`�Wt-z'�g��lܛ������B��� �vz��VOOx�����w��,]��CD{�#۟��
�`���k	��3��^�=�9���Gs�-���怃�
F8�pt57Fv�T�c��!ТB��am-���"�׶�S�g^�^�.u;�,���{n{zf�cc���%^�y�ڪ�mm��+mXE�F��\�]��Em��ꍙ�{NxS<:\��/�c��{������H��t8]�hz'��xީ#��Uo�^����A�����Y�D�[�^s>��z�Dpoa�u�d���۞��i��`����-U���k�o�<3���{��q�]2tfGyر͚�f��zw!QT�C�je�Z?1O.���`�?c5k�w�=���xR�f����/���ܬ�唅sg�R����\�޺1�#xVu���d[�6�oF�>>�˽9华�EU�r�N�mja*܌hS]>�Wk����s���l�|����G�-+y:Pf�+��v�ғu��/V�]�s'I"Rн�)g#��8��X%v����>�&��)�Reζ��$�Hѐk�caE^y�������ٓ2Wv��&-
�������t��2�%h̷].�Mȩ��'�wS�È�aՍ�w���^=�Hj�<���t���	�u��9�_EY�d�,}c	��'g��w�:m1��W�	����(��jf:�s��=z�O,=X���Fh�p0Mz���Dv�L[�h��h�q���Z�k؉��*�n���ՙERWRJ7Y:�`�����R�c���6[}�Y�J�q�wޡ��	fqځ�8�+)Y�7p!o�eΊ��tkU���`�y�prT�\�}�y��;��7<i�oF��%��]�G{(�?.��\�E^��I�	w�Ťh=;��f�\���r13:�0xg�':r�>���a��;���vS�lV��[7s�1����9��(Һݣ+s�Dn��u9�^����{F�޸����[�r�ѩ�槍Y��x�\ڵ$g�
*l�6���G-4�(hs�4z�V2�1�3f��x,�&�Æ�;�T�1zTL�y�/��᙭�";��*;���K�>@Cy�[�j�ڮ��d�2�\�f�WW��)����L�X�Lг�Z�fCx6}|p�=�qwa�H�̍l\��^�QG��^�\�N��nxiL��psV�Uz��f���_4dз�rʎ빅'�Nq����nq��Jh����zT���6�	1^��Yb��8{z+����bҁ!��C3�zLr��4�4_)qn/��p�0q�&B���VŻ�ӽ���?k��Z����Vw_s�7����tgll���ɓ%����R���2Y�8���h�
N�/%0�1�R�V�z��y��u,	S�r=�/$���X�u����^o�iz�M�������zR�8�Ey����\WS�2[�W�@*:���6�X$n�X�ت����p��2�!wH�7n�5��}�_�� �C	�|��	���j�:�z�aB�B�s2u7e�1�͓�/�����V��
�6�:��.&���:�s��M�j��꾦��YgduV8'��c���s����=r���rr�3{^t�SU@V��
�<V�M'����S{g�t���7
��v�{,b�{���T�0�}��Z |Q;�sʉ�p�ˈ-xe�~�H=�3�]]6ƌۅ�؏�N�]��W]lL��;&"��	�>���)%N��̼Y�p���Ͷ��"�no`r���8�B�Q���s���\w =ےa��0S/N��M�5�����V��4�_0�6�{zY������-�<f��f�ϳ�;�if6�wm�Sh�ciܦX�ݺ���Ӷ�m��n�D��,ȍ�Y�nܓj�$q6-�t�A8���k7oz׶�q9�aVݹ$fGZ9�Vۓ1�Sj۽�/�80�3;Y�-�e��9$%%�^���{n̐3Rp��t�\NR�Ԅ6�9H���� p-m���)��#2d�r�bD�Vlѝ��M�l@W������+Y��B)Ȥq�[,��D�=�$lH��/m�R'8�;�{i���JE�
r�Z$�����^غr��v5������$E��AenS�n�G=l��58ㄡ)';���$�tD����B����ok�=�Ӕr;m�H����[m����-Hyj	�p;���܅���{�w��G�����Îmi�8NVl��$�mbY�u�8���8�#�g"�gB �rI�y�����ƅ�ް�wX�g;ܫ���!��:E�8��׏�g'ɍ���Vm�(L#w������G�P�$��ٺ�λ��<�������ΎB&w�컮����Y�d�؆��0�FΫ�b�zq�D��V���}����W������4����N߽�Y��j�*q��r�<�L��/��{�u9�X���H�f�۟j�g�x�e+�b埭}Ȝ��|\�H����{�e{ϫ��Uz|7�]�M�Wn��X���xŇL(��U�e�x�/��/>��)��q�T*0~�!.7+��粡;���g�k6���X�l%��S�>���h�p�^���3��������V��$��<����c��}�
���4=��+��YX�y@�}��qIݤ�.�\��ƻ�*���h��e��Z�n`X�b��:m�]�8�(��(�q�Q�U���
��LBu��}6_X}2��f��3����i��^�;�Y:�Ҟ�J�<1��U�-�[?է��w��]��g��9u͇��f`&ct�I�M��h�2��n7=y�����&4����=�������4
�&ެXwD�zW䡪���Q�`�ܯ�U|'0�s�i�b�[����p�Op�f�20TL����ח�%�ԅ�Q,'�Hv 3u9�}�U_}_Wڗ6p�����D�n�9Z��>>}�+s���="�C'�|�m�9هKq���p��Lf_�B*㺚��.��}S�J�gV���):z.����O}���\_�ڮ|�=,vO+��5kZ����j��B]^q�'W�5��8&Մ^nG>O]��N����]q��V�\=��]�K�+k;���ۇm�ɦ�綫7X}�(¥�V;PV�� �\�h�d��/{�6}�Wn��q�I�J^��'Y���eN�9Z�ܖ��K:uC��op���U�ּ��I����0�{�O�{|�[	��+�nT��յ�Gw��)�ja#�]tT�������F�tħ�q���4�C�k�ܼ
;!�i�n��c�����{��U|�,�~�k���Mx�zѓ�F��*�Z�ۉ�=�'�i��0J-j�uDK�6�dN'�}2��6�۲Ab�%)oṧnV?QꜬbKS��K��o:�D��<����[�d�R����]��/�u>�x�c�f`4śl��(,�Pvi-���d!�U��'=#��`�O��J��m��Ě��g�.���=۔��et�6���ﾈ����X�8�F�{�粡/�B�n�ʦ2T��`�®_V�;3���V֥�.-f9����F�rBN5��n)�`�2�����sx̫?]��qT$�ٷ�{2�L�]�>FW'�B�WjU]��Z��r��Op�y=נz~d7����~-f��[U����ߖp������w�cS�ڶ�ss��N� ����{��o˼��|o��a���D|4�:b�N}٤�U/g�5̽���&�Ɇײ�Up�6�!޸����]��kWAP�rS�vV������{��4�3��kؖ׆vn,X��M����&��8{��i*~�z���lΜ`"�rO�ξy��*hU^F�˵l�ۈ�x~��}�v�I��Ӱ��U���9߳�1{(bď�&N�y�ސ�(_�������Ho֜�m<��O��&������j��pK+���I\$o<q���[�u�[ ��^VS�m��o`�J�/�6�{� V��S�Aa6}���s�{�VA�>����3dWm��7n��aȝ����ԧ�o��l�߰�-Q;����LK��q����>���oM��P�OK�]���ogV0��-����F+�cK��{�s	yZs�˹u��i�<�w��,����Th}�+���u�*�Od^���R�c��LW��hD�۽Q���0�2���Y��+�����LL��8d�fT���Ӆi�%k�in����S�?6�e�BSU/�ci%�ι��7W`���_tүر�s�]*ܫ�.*��S*�эbu��cJ|��/�����U贞�|��o;÷�ޫ��2�qv�T�q��|Wf����:�u�Zb^�	�啎َ�T1A��o����9VqjI��u�!�i����{������io�����7��<��y�z���%"��8���F-6�:��Sd���"/�q%���1y�F�<y��ƕn���$��yk�����j���y"k܀��Cxf#8�'�&z̼��:
�^վ��򬩛O6�m����1v;֮A�;��"�Y9�ܻ����&�Y&J(�b�o��g�e�]-ȫDRX��F�1�}���ETDp�2q�rd�y�:v�ӆ�i��vN�9b���q��SUw��E��������A�T���������[旽KO�r���|�}Z'��{<�B���g�v��~T�ˢ��N��Z�S%�N�E]a���1@�[5��Pz�v{�	�[Ԕf*�,n���椡���!�a��Tk+�E(\r��ְ~�h5o���R��[��rF�j���wD;S(��a�yqB��(�I���`�\�xr>��~�iz{ފ�}n���FS(�QQ�V	W�P|�^��^ž*�p���}=[���{����ڮO��O�7�G���Ԙ}k�����q�e�[�VװF�۽��I��O�{ˁuY�������v3��j«R�'NUz���^��2~�ߨｹ߭cˈ��^1a��N�U�Ir�[�� e5�r1b:�^��Z�~�������<�����i�b�.�gL1�f.��^r��bp �T�s��M���)�ג�0�g�=���1��)ڔ%�7tr˷���s�MMC�E�!�|�%��.;z�1�(���s ��8��qY5�����On�#t\po������f���9{+=��Q�9��\��\i��4s:��c��}�����c�ܣ��v�і�U} }���F{�'z�e-��u���qMۓ�� V:��[��Ɋ�C���1������z;�A�N5�fNCE�U/z ��A���-�G*l�~0�����Լ��i��]^���~�b�K;�@^�~�w��H�$��8��$�<�o�ʾ�(����]i���Zc��x�N����ev�ӵ~�/�}�$6�Ҟ�I�VyZ]K�����\��~�I�L�y������m�g���T�:�wQ�J�9�K;��Ԩ�~}@\�E�0LT8�0���qӯ�ǤU�fן!qW��3��WP��8����.8�"�7[�AC�|�aݭW)T�5o?��n�����uϑ��'���:[�-)��P e��p-�ri�眫4���Ds�][l��Ɯ�&rǏvv����5\����E���/:OX��E��o_�_z���0/l�c	����D��SRVO3�3���mb��^�v���	C~�[;e�Sm��D��_�e��^��X���W5�+��ݾ�V�$'�乘�qx�S-�Q6�G�.Y�B�ܲ�C\Y�@��N$�_{ﾯ���&�O_-jL�`���1j�C����?}\j1�ک�/o�	����7��M�a�G��t�E���Y1��FJة�`�<��h�n���d�zT�Ș(��[�ZuK�Z0�q@�Rͯ�1b:�V�}6����g%d��眱��sӫ��RO}~y&y;`�T��Z����{��}կ7�H�ZϺz�?Go).�;���r��˜�GT���LtԳ�3�b�m=�RC�����%/�X1��	8֤�>��jؑ��s�#�+�ڼ�sN?Ou�'�@dۍ#U��5rC9�L�{'z�u^�Y������^Լoī�rS�+���@�3~��]�%�����ϖokZ׫�]ߡ=�-���}�s�{��uW�)x�7��k{�r��.��JzW��:�}�l~�v��=���f�����U�L6��Yʮ��[U����g���*����h��p��	h]�,����|�ў֗
�C��C0����&�E�v|}�lI�z>�=v�w�x?_`&��z�WZ+&bm��s��~յ^�ҨCG\���랤�������.F4�@Y�|��k����^�>����cw�,��m�P�2�y���0m�-��.�UjN�b�.�.�BmG�?u,>�%>�^��E����t���O�����shɳP�o:��қS��S�%�8|r��E��ri�e=ϕoiRj8���MrΞ±�>�l�9��9�]r���/oO��u~k�I��iY�5�ФH��
;���pո���/a�2ʥ:�>��Os�&v�Ӂ%�F�}��{&����u�����N��(��ɎG�J+C�3��k_f7�������OV9�k-�\�ӱ�?S(6%�Z�����[f�m���7���XX����:�n�zK�+�{�o���MT�A�ʥ� ��v���-�����.��]K�������҇O�q�ݱ��j�2�Wr�W�9k-����-�^G}�i��{);쨰g�����ޥ�3����wV���MP�V\��o0o{4׭:�n��m.��.=0��{�e�]Ҩ��L]�p+�n��>�v�SZJ������әn!,��+�x�%�6s�=�<J-��F
�}���a�g�s�U633L��E�Y|�μ����C�s�����ﾯ��9N��=��!1�;m��WX��[fwG�c/;hY3��nCc�:�cV�,9r�O�0�Y�^�{��]��[�r�/�o����3-�ֻ�.5���Wf�1��-M�� h��cu�Effv�9@#6*E�h���Sv��~PrsԽ<���y��^�G�@%�.OQ9���'%q�VD��]�OI�g0h��z֯Q�������8���4��V�%�&}4���p���z���ίM��y���c�a�F�|��HH
������QW˕�ֱ�vV��0��*1�Ɣ.9O�R�y�Ć��/]%s�'u��n5[ͻ�L�Uh�O��Q���vF�>r�M`���Ƈދm=QM>��g;�(�����V\PY#ͯ_w��Sk��SJ�_��Jy��~5����<?,ն��(ů�t��ù��`��9v7X=�&���)�7��^8��3���fǗ2�EdY	0Q��a�07%���Z8�ށ���A����p�?�^S�+`�ys7��r�R̅�O]��YNG�u��,J�����]tĖ`ȱ���F�����j�]!��ՙ���UW�V�Z��Q��������ݝ�Y7�F�R���0�L�l\�=x���s�0��7�Oƽ��y��Y���S�;�o�ڪ�^F�y�����*�Z�A,~����軇�ˏ��Tʫ�2��7��M*�y�s���_.ew�B�<1�԰ywN���[U�[�'���b:�Z�0S�������6I�ҵ����v�N������{a+¨�z�#�P��,���[p^N�=I�C��x3\���S��״]*�Oy�h=N����*9,Ѷ�^(��)�G�YQ�Y�Y��ҷ��n��7��ɺ!Q���W��d��\�|w�D�����T�{X��k����u��ո��}n�7({;��|���Vם̪�ߎ$�<�m.�T|�~�I�y���\��s�	��2�o+�X�^�msH����j��s��J��qu)�:�tA���"aW�ؽ̠�o�ڇ3ٸ\�o�;fRY	˹L��`_n��5Et���z�-k�Jx
�5P�����db�T.�-onQ��wb��On�eo�`@��/-���E�6۹���ݚ�NW��{��>O����L�vZ�e���%�_�P����V�ѡo#��VS�89Y�rg>��(��D<,\��Ђ���&���fW=��NW)��ޘ,62���O-6�F��}�f}�pP�>n���R�+�K�	v�u#7ͣ����2�Y2�b��J��Kpu��E�,����5j!)_���G"X.����l��w�-%��Y[tT�4L�*֖�)}�MgS�V����{��?�i� �'����R�/HIMݲn��c���M�w�����>���M��R��RqY����\�����c�".QN֮
�b���������O�˼p7ͅ�k�U�2r��}�:٨sPve����W�/_��S�{�jQ`pn�tp�>��4 _���K.�W ǝ-�rݑ��2�ӎ����i^��K�m9f��h�`�����r��ǽ��H�ˁcޮVq���*�@fQ�2�X=�ֵ�Jd�N训�����y���	��z�"]�^.��X|!�p#O|M����|��W<֮�Z/1��҂�M{�����:�K�Y�t��-��Q�$Ap,�[�%39&Ü+p]�vm�o�e�6
rn�z8x|ċS���v<U!&�0Yr����N��3(G�ޭ��3l��d��V�����ta���ckN5�dY��⻕�_h�j��i�69���Hg[�؆�:+ۺ���� %�t.e+<wL�5bѹ�j���T��,ݷ���֋zuZUn`�s��NF�-z��Ij�1M��V��l쫠5��'����0%BAu�������2�Y���I��Y}�!ǜf��Zl����r�U�ݚ���s�A*���٤iu!�j��eg5��J��yWm�7wf5lG�]l�4�a�=���*�b���]c���#���g�)=����7���*�s���̓���1.�u����������t���P�Kǹ�^S�b����P�,��:pz�=����Zf9yc'g9el'�|7����*_��#\�A`��쫞_cգң�=��F�{��A��7��H)�v(;/�vB���H�u�I�LkY�kn�q��NA�����p�������\i�����:�x���+)L%���v�h9����^�	T�.��Y]�gC��H2�tJjƢ���٘��������O�(����^��O&h?���6,��e�Hf�v�T��FѾͰ��6��ns]i��E<y��xR$���mv9�t��C
���:Qޚ^]�y�w,�u�n,C�웸�LT�N]rx���:�"s{����sZ�)(U.I.1�Iq��|b"�ejfd8���(E$ᵉm���gYۏ�yh�H��6��mZ��䓄�$�� ��;4 �
p�Z'f%��):���&m��"py�H�=�C�.��m*t���8�����Z��R�'H�)BE��V�g'YgH࣒�DrD��Ў���Z�\9����N��6��V(e��R��䈕��9�f,�mkl�Üs� G @�*D��zU�9��r���N@DA!f���'"I8��B��s�Ge�'ru���!�ۗ�m�n�N8�ӄ���s�f�#,��[k���)Ф9rR%be'C2A �B@�ÊNN�ܶ�՘�9"q���[nH�Y��u)��N]�`촁9(�í'�BrH�@H�K,�ì���㣀���33\����Om	Y����h�!$����}.�	�oZ�ʥ�(T�;� �}�f7Ws�nW��
/m�Z��Yᦟ>�������]���E=Q:���ZV��;�VF�f��0�*1��)C��Ԁ�빧ƶ.���:���\�XE��s�����ڙFZ,R���A�ǳ�Wf�9�{��^C�WP=�&��|��Vi���Z��m�i�����Sp��ˊ��T�T���j�COu��{��W�w��]��/`l��k��_.������������-j��ѧԽ=�d�v��jWt���i��7�]b��ں��M�c{~�v��:�N�/Km���u�7e�{%�b�A�/b��ж.mh���NS��%>ww�X�y���a���Kܖ���v���Q��-\`����t�Mq���_��+���V�=~�ү���y��V�1�ݹ!'��ފ�7�"��c7ޫ%��u����^妏��� 4��?��՞�q���W 4���e��y_�s�9������ek���t-WN��6=�	�]��T���!վ[�[���O��9u���Qf�&?&念�R\����5�u��2ۺ,,�w�j*���L�E>��c[�a�)ԣ�4�kd�oD�G���}���<8�B��@����Uq�s�Y��R����{�"վmf-�Q)�йw�	=������� /mH���ߖR��c�ȳ6ĘCn�s6�*7N[|�LCY�����x7�=��kiw�v�{��Dy������\`�oF�cnޗ䏸�����ma���S2s8� ^�&��/�����o_N(Э�+u�E�A���5�H[l��X<��i�zjd�},��b�ڬ��^�z���mL������W{����  ��~��n4�1�?wx}�K`�F�����Y髨U��w����$�)��=��~>��E����8r��
��i{z3���UN�/�r#:�ΝQۈ��}�.�s�m��w.QmL�
�Th՗Aa��s�g���[�g_az9��ڽ��?S��L�q����:QZA�XˑSv!c�i++A �/KT)Jh��x`����.�={����!��	/*e�h<6�K7V	x����ܙaAD���7�|ށ����V��%�����ɗ[�@��ü��ut{��C�-�!���O/L��A�l�4����=o E�z�8��>�;�}UU�}��f�u����,���,��������2��������*?Q|m�xHpVS�v���R�ry�kM[2:޸�O$���X0J(������1�~UeQ�����X�BJ�Bރ-���Uf=1<�T"�sl��Y����/FT���z�c��pٵ~�(.�I�bw����ڣ�>[�3�'�C˺oQ�`�S�5�]���F=�f�ۊ�,�x�5�rS��J��\������Ƶ ��ȯ��2��oЁ�ƃHr���]�G�_a�rv���6��/7*?Z,m�	֖����P�����$։8����өB��kT�U,}�����^y�~z�{��@%'�[5��&́yC����w�"L߰����|�~��m	����8�~ކ�5v��n�4N��ukHnl�\{,�W�K:�R<��V�3�Ϊ�������D��e�Q;��2���r'���8K���Ϡ�#���q*��u�P�z�+�s{���A�޶Y��1<��_��޶7�}K�xyn]�
�v�1dgz�_�|���+��94����r�ۃ��Xh>�ɜ�N,9��'��������\��_��3k�!o!���K�;bɵ�]5g�����f����oW�X�7:��ԗ0�{�
��Co[�2��F��v�˧���j,��,�/t�ٞ��[l��즟1|�L����!U4�z�o���*a*J'�6��󇂶��D��ӝ�{VU~��P殩s��v���[Sp���1��u\���O�5F3��&��u�̬�nD4��ndk��w���M9S>�:�<��yi��������7��mu������~��t�l고����F,GB��,{�X�뾮�9PJC���}�O�_!�%?�m����,��S��+�!��¾��Of����Y�VU�s���^��o`�;�~�e/zx^6ul%c��E`)��Rc{h�=���Z��|{hQ����]�f!��T5l˙��-X�tP��Y�+�(5Ia{���s���n՜��C�\|}�g�X3.��EǺ��{O׊������ۇz;���-a��O3��r-R�~��y����ݽ��v����N��r��O�s��� �9o�Ni�e�(��X��o�w�?⪪���Q����	-����~^Hg~ſ5���^����0�l�ئ�CfF
ov��^�R@p��? �9��kWy�~-�S�c؆g^�w���w�ϻ�I��Ȳr�w�_�~5�=�+[K�>���� �j#��7y���ݺJ��zE]�'}�R��s���a�;��W�cܯD=���D���sS�\g>��S�pվ掵}\U��'�;%b��c��x)��#L���^n�z���ܝ8���jzv��	�뾝����u���+����9�'�B��t'��cIM9z��ʳLb�ƻz�w3���.��/XU���|j�+�9�m$6җ��{�m�fɔVwu�s;ӝ����K�.v�L��J+F��V'��o(�5��;,\:�-�F�9���-qi�1ȷq�啓��EJب����e��=�61��^ n�,4��ttb�{���;��h/���^�^�X�9��95p���غ����1�b�C t��SΆ�Q����&h�߱��sv!��qSUڭȷB���Ѡ�jI�̩x+5!��Z�����uϛ��le@�Wb�:��Ф�u��}�G�V讫u��ܯDM�e�'�~x��e�K1�h؎��vy�O<2��h��^�W���R�l�mDKܒ�ȖX��Q���q�8��t�.���kB�/|�GԴ^l��f"�]Df1[�e_ҭ�Ra��@E���g��I�E�d�ƙ�����oW@����ye/_eE�>O�y���~<z��8͊9�_o.�P�bz�v�Oj��9�Y����=^��C�{�kY�'w���uY�ܱk�5�t {�� ��%������Y��yӏ��<��m{�Ǉ��ܩ�U�}����{�&���_�g�+�t�Ō�E(��Q�VΏ_W8 ���R������z�5��涑�u쳕\#�Z���z�c������sju->�r�~^�|��>�8����U�/k� �ӝ�7|��z놯R�,
M5=n,S�YXb�.8��#oճ:q�o�ڌ�W6\�I%�»$s$��\���f��UΕ� ]����evR�B�pi׽;V���^��^x�q����p�pY�K��%`-8Y|#���jb��2YN�W���������+p�YQ���&��Ѷz�d�]�?��{��9�y�[��ߪ����X�<��X�Ws��ČC���P�r���`�&���yK�cd����$oQ��fx*Goܧ:º�3]%��L�ߐ����&Z��(/)�q�ˮ/{��}�x���a�2�ʔl�*����V���7��^vv��V����n�x�E��-�h��WS�%u1�^wϦ�X�
`��D�:�T�����7�X��e�K1k�H���q_m�KZژ����K�F�镏�;�m�1L�{i�yL��4�g7r����GT�@��FU�%�W<�__"��NU��-ج=�)��:����O����{��w��Ζ�[�YK(rw��ųъ/Z��T5l�T����\�|;�6rr��ͣ���i���]�z��
�'��*�ϧ"��*�}t?*�wvZ��{N9O)�m�y �����Eb8^
̲�]G��fh�W�mc_.9r�`�v?��[�p[�[��(�f���'S���}�][��⣍��[m����m�N���-�PZxz�Y��Du�˭�}G$];�_EL�X���DuʦT�/g�`J���{�����g�Wk����W��<u��p��,jc�Ol\�c�C�����V�|�rN�8��$�<�m)�>Pyk�����|���ݹF�-��R�&�z�q$(
�
�\��"��np��[�c���v�!:{ŁQek�^�%c|�w�����w*��^9�Ҋ�.�k��1�u�,U�coe������r�Vn�{"^�3~��&q'�-��߱dڬ���y\�tY��Iݤ`����Ë����r��{���6�u�S)��}BrGӡo�xo�Z�Jt~+^�J�[�0k�1�������M>�Y��\���r�C�dg�[[�}ӷ��~G,��e��Sr���]^[��=��?0o�"�cIܝ��c��M�%�OƟ�[�������a��Ѫ}K���]Eu�/�5mۍ�6�.�E����_s?]GTJ߯�ϧ��-���+��'H)��	��o&=��v)^xPEg�-�|�p]f��v�q17	�L<Z3٫���D
s�K:63^�ע�u�Z}ת��Ƌ�Y�,q�sog%��-�S��d]�{tr��+�{(u��9�8]��)�n:1���$3:��n�X�}
Xz�o��9�|�W�}U�^�,a�'ܴ�E��?W�J0��\�B��-h��ܥ��7������ ��ϔ,�Z�\�ra��~�!ST�s�>�(yswW���ܦC��Q����Q��C"7�ʄ�ړ
!�r`"���/��W���Z��G���[~�Ԑ��;�2���hNG'�o���-�ds[���w�Ӌ��n��<h4�]��,���k�;���,_1/y�T��קv��.JwE|}� 3�߸�ߎD�9Z]�{i�&�K��Ԟy{y�<��s�x)���lo����7��y�iu#��:�y��Z��j�E��߾����="���2uW��mW��p�6����\��4�FΓ{U�,���8P�����վ솯�Ճ��Y�����V��٣�_F�ݭA�uыvにX1\�\^ns�^�n�ʆ_E�͇:u}#*�z���C�`�����\M�PS��F��t�@�,_r���Q�8vjC%�06]ӖZ���.7�٫2ZќM�A�@�=;N����3W�ޣْ���z������Ok1)A:P�����;�ZN����fB���|��9�}���}U�#�Uq������#<�������C�MD�nf�����q裳��~��1}�ά������-�9f��@�R�.6@�cp�9馕t��;�@��7�=.�}�N�Z�}n�������[ʖ�Xк�Qѝ=�E�kS��nF2�L��e�,��b�VU����ڹͲksמm���������{��'�a�b�@�R�Z������y�.u��ۢ�ݪQ�{�K:t�S��^i��y��ky/r[w�v�
�5R�H�ʻ��;�V��M�n��-�CLm��U�%�Ny�����k+�>�ͬ���Pz��Ze�ў�����j��/E��%��UO�y���~����f���V,�;�U��YU��6��Ƿ�!�8�,Y��O��?3�ok}�-�=Ӱ��3�׾�����z2���.ן�"[�r�~>���dU�պ��M�qT�_N,�g�9>�-s�L�oD����)5��E;�5yVv�웨ԡM���BS��v{�����X���=i��\��x%^Z֑��[wK�ݣ,bԄ}��)G�m	Y�����m:�o��`�P�*e�ϻ4�)�2���4��,W��f?E��m�&"����|y��#��k~/��|���[��Ŭtz35���_{�r��n�Fg�oo�d�An�{�
�R�һ����al����u6%V���x��oW2�Ja;};���bY`�l��!yk��y�a�Dkęj�T�b7jE���_r7�[��%9���Ǵ��0_oz�M�0��^��	���*�y�w���<�E���rʲy3۠3�.����P����:��;�-�����"�1S;�x],�N�^sn�M��/P��e��=��g�.sy75°p�Pk��Od�~ב�{t/2�b�u8M��h��s�7�:�z���b���vz����,9}�e#���<�[�k*'����4��u�7��z`�\�i��<����D�6d��㿋l�#��+
�K���/T;`0�=�-TNө���O4��֚�$Y�c�г	�N��%*!q�qfk>0�t�m�hN�7�PB愵Q%�ՙӑ�gPx�!���pa�=�Xйs��ft�=���8B'�;-����)��{}Y �����>��(:	yѕE3����4��$Y/N��^��[g�=��z[���T7�G^�c��d�x��\W=�+m�G[Qe����~w�G͝]����xJ춻|�c��0�wv֊�pA��KGnjb7i^� �����壝n��k}9�D��/UJ"
��Mwˍ`yt�DG�K6�y�\Ec����f�Q[��_Y'�oxz<�G�.��y\+K�2[�M�E��9���RSv�2�(^:�����dU-�Dg}Y��ɪ��L�wl��,��#����a^��y����sޛ�z��l���Xl>�>�SP'�Օ��/v��}m��ז�-���SNIG��b��P=�9��@]eb�yd�:�+���޴�@��H�&뷔���h#/7�sH|ʬ �0�Ӗ��]���������8�\��S�e���qܶ_�v)fnβ�_6�WK��^>&jf��}E�nYhmtK�)kS���&����|_�/zYV�uej�e��¸�Q�(�n�je۩�y[�龷�Fa�'QL,_l�Zzć��nu��j�fV �bi�5���<_�1��3�����\x�f���}���Z�"�1�*fi������W�BulX���'W�>��އA�=4�pq cL��r������J�o��ŀ��t&>�	�c��IA�56纔�z��4���\[�\���N���U�S�j�a2�a�5m���[,�2f���n�`�ϳ��B$I��H�Ͳq8�p���Y9�Z:$�����%m��98�"6���3��5�'�;8�ٸ	9͹�6�H.G:Yd��qN��rmi�?���t�K75�:���8���$�r9�vFKl"��hq[nY����hr����!%���m��b;�G�$��rvve�m�G(���$����k.D��h�C[�ΰ��Ii�$�m�G�� :t�6�I���"\�N#�s�ly�$M�ڵ�����m�Yam�	�%��q qТw$�"ppF�6s�Hs��#�	%�:s�;V�3��;;%)H	�p�"L�ӎ���6�P4"s��I�m����JG��I6��$��tt�NIe��9�� (��P |>@�z�L����x-8(�[��tN��Ƹ �5.�ޙ��ic�k#�Z�"���i��s�t(m���u9�F.�%/�����ۮ����.G��MuvJ��{��ܑ>���؛�߂/�5��ս^�B��:���锱�jW�矍?g�5^e１5^��~�o���.Ԏ�ׅIK9�ˤb��1�-���u,w�'o���.��)=f����fB��+���}�;	}�^���|��??V�Ν}�I� -��.Ff���8f���؄�Ľc���f�gWMY髨Q���p�󺘎V��v��Mo+��pkqV�n��v�Q�V�}�u�Fk���*���vG۾0},̛�%�o(�pm�1m�������h�E�2�*QQ�V]��i+A���+��ܚ�d�X��Z��y���D�+{�k���	� ~�p����]����%��vT��{ь��0�(����'3WLSDh�F�cz��kc�ب�hG-߬�v�R�I��2��:�s!C���Q�����LuA��]���C��6!�,�ztEMt�:��ix���R�딽��7N��2鍂�.�ez(����ɡ��\�-�� � ����&-}�`^�}j7�}����2*�9˅�<�K�V\���Y�s���}g��,�꯾���L�|��~.m>��4�J��o��M�����r�<>�}�����]��Z� k[�êW9����.�qi�f�kt-�4z�j��%Z�Z�h}��"[�jLg���CV��R�dnJ�0�[S��4������󇶛���vl�S�s�ӑPՁ_5r������t�J�y�XN)���+(����n8Tm6w�?��?l$jw�:˴N���rE�w���!��-�+K��>ڃ�\�?<�3^e�K���vh�s�v�sӻ/}�V5���/����Z���l�fyx�4^��2�+:�x�՚�^���݉3�O�(������3�vJ��	3ϊ�ns�;SJ�/w�0�`�T��l�~+�V����F��7BN*�Y=���$�l�EB���oN4;}��FՍp�L���b�)J�SЎ�C8f��
#X���?���̤���g� �WrH��r��P�Ò��[�4�J��ty6��k�\�R�3�зR'�K�ʭۙ���[ ��S7h�.����\[��cl�@�����s$#��\���i���nS��2g:���""2�ʍ�m�O��7L`|c�Ii����^���M	Gw27n#hxg�|:���;�%{�f��R>�H���;~Sr���]^\�)�b���{���ہmޑ7�׹�{��������V���;rj}��^��m�~wٛ�[��Ÿ�=��ʵ�.���[7�m�{G}��߻�6�F�A�op��|KԤ啋%Z�`�R��|ѱQ+EP<�������gb��Ź)v�]bS��λŦ'�ʄ\�o �l���+���K�Rz���z|9���qjPoi�WWד���{*�S�v��7nLX#�_+�ڵ(k��R�����!k�;�/���#����rq��V_NE���SӠo.�����{~�	���@��4���/b�f��b�k�ٵ\�A����'�oijn����w'�\@�{�����Hr�{�gw�yZ�IBׅ������[�כ�|���ڕ��;�����i��l����E�A/3���5ٽ|�`ڎV�HZ-� VjX��O��W�j��j�1��K>B�aTQ�{��]^��y��o`��[��4���~��Ő̏����w$�\�������{��KoR�q}�ӭ��:�����H���N�:Ğ��V��R骒TNg������Eo�^���z��5^�a��\$ͬ8�h�8�R;dW/ N��S6�T�{5�A�X��ݐ��#r�~t�о(46����5J��G�d�-���.��.���o�:q�v�5=;��Lf�G���q�)�}� &Ku{��������(��Ϲ4���뗰��O���6׏Osz�/!Ʒ�_ogV0�	=�T�Y�3V����F�t2�ނ�:K�a�\�1���N�E�1k�Qt��F�?N,���J�D�à<�e�S���m8;�ۚ���0�od�W1�}y+>�u�fxd;Z������ct�ʿ7��8�[���.9=��4�!��b-|��r�9���4�^���C�����÷���ky/rKo �l�x���>^9��0��k�]��w�`,u�R�<��=���aN�����Yv+x��.֭$���LӺ��b�߼<����N�-��ZЛ���{��Af�	�1z��`>P]��#W �)C+k)�7����>�"wQS^�s�5�q�6�ҹ�A�� �����Z����{�@��13r�1��{*�%[�h\�oOU���i�yq��]�K�~
���@�>o����r�;(W٩�[�)!U��5�]j&���wZ�������Y�R�����{a+ò�U.�ͥ�)f�U�{�5�2�>+��WA'SΝV��ſzY�� g��~���D����W�s�ܔn�V�r�w��f�>F	���.��_=��7�n�t�<��s^z��i�9k~S�T������??<������0�Oy;s�q��9�볭�2_��c)ތP"޳5D򷰝��M�Zh�v�-�v��]�Ԅ���kؖ���ŋk:�7��2�P~n8.]@�a���OO:眑�W�sx�oy	��b[^��6�:�h�=W.�5���o	E���t�H����C��k��o�Д�Y��YE�$��Ҹ��B��-�׳M��٠n�M�M,��Ʉ3j��QyB�i�;Y�X�[eV6�]+ْ󨓄�T���k��66�,�:�
ԶEo�����ӊ�m�Tw�L쭷�4U��(.���1��4p��Рy�`ǋp��u/}E���=vS���Xj�bӗ�����Ƌ�a�2ʥ�VM�o��o�U�3�h"_{�m{��#��<���ѯ����1:o�E�?BɎ]=��i�FL�
�ւ;957��18�J{�KF*,��%�^��]g���S�̚��̓��of��,Q{�}��r�_�eY���N�m�_/C}�{w��է{���iy�x_�*�6��F|�uJ�_@<�߽7⯒���gF�(	ڠ�\�py��N۞�b⛶T��uJ�|(.�M��zԺ�u~�1�G�z��^P��+�8�p��CsqM[T��+c��M���vc���1���3��b񑁑������wU�}9-������b��wP���z�Kj������}i��U����?��X��#Ǣ`
�Ct�,^�.{�@�&�گ�Imgd��1:���x<;�5��i֐Dp��2u�q�8}x�
<��h�$���`�t0�&�\Wa�:(�g,�p�T`��G���ܔwwn�
0�h]��4^�����a�T�
.���A˻Nn�v9v.���ݮ!%N�	:�sޢ:>;�O[�6/���}/��O	�����ﾈ��݄�zՃ�i"k�XH��s>�����]B��lD��S)mͱ���y��Mެ��^�W�L���5쳞�~�8����WP#��3|�.�H�I�8�/9����^���(C��:b[U᝛X�}�:�ܑ�@fZtA3��ڋ�oԽG��Tފ�-�*�-�q��1
�uC{]p�K�#�P�ed�9�G�
ܕ�W#^5i!i����/S�E�˚��\(W��V�v�T$�����yA�����iY�������s3�)ǧޤ[2OK��p6Ͼ��K�\���fNy7)>�f�D�O������-Zу�-�.Y��q�β���͝���1%��xP8�;�nS������/���Q��{��_U�1��{��Y9�+ӷ������v��طLO-�r��n�C�%�}�K�w���{OG-2zS�s.��DY�nY�=�{ʬ���p��}kx(ƃ�5��z�0d�t�fX&Ҵ��-�i<�S�43+g]򙛚���gpi�Ln˝F[��Nj���C���"^Ʒ<�=�*�*���O��bZ�BCk��+�'A�:�����Q�y�y�k�#�j��E�X�F��W)�;�.)�rB,0����j��ION[��h���v���Pu9��jA���$��ݑ�NCv���d�m���W\@��[����Y��
k��b���qVn������8��a�Y���ݷ�t~�Y���?�oJ�g��ը��\���w/�Q�nq��ӭ�ޭ>����d�߿;��7�=�����M���Q����g�/������="�3|�&���~�m�Y�������]�F_���oJ?c�of��
޵o�!��V�⯙x\Usop��OS�.�	�ޗ��:5��S��1�Wؠ}�X1\�_����+T��P��h����y�f����:�~b�\P�1�����i!ɧ�`�/���Y��8I�lո��s����|��aι�3I��3�~RiT�rt}�V�q���#L�`���}�;5WNKS��)��[R��_4!1���T�a���N_
K���'Y�6����w/%f\���<�s����q$ֱ�y�� ���vk5�!��Ss�*�Nw=��YΉ�o/ez���eu�69j��}�r��9����z�kk˽��i�|z]��u;}j�-��'���������I�//9�d�=ʞ���&a�)��E�Y1ˢ.�*V���u���2*��5�J�?YL�n���/��/���f-|�H�g�KK��p�s�ti����y�G�k��__�����&w���]O��{��9ۖ�@�k�GTD�ֈ��ʻaF������[��9���^�X�/{�U��0^7GP�ϼ^��+�~�r�Z�_V�%Wl,]�c�ڊ�9�?t�\�=�?S����K5���&ߡ�1�U�Hw�5ˏ�u������'[�z?ToԦ�z�;�B�ܭ�D�����{@�nI����<��_�`�g���,Y���_��9�S��N���y��{�ݼm�TĤ���0L�g��]�X�jV痧�����e��:P�W�'�ߛņ:����\���Cx��n���"�����eF��$��-Rb����ʊ�*���T���`ZwHW�!���rA޷����M�{�'��y�ǖ��ɧ�y����E���YD`�X��]�6���+�Y� {\��p.ї��)[�`<-!�y���f�^��Ɛ�y��C�~��?E7<cz�uF�X�;{��bͥ�Q3w˽8�W$��;l��K|3�j�b����]Qu?/V8�a�//��4�B7ܬ�k���ĕ<V6���Y��)a�`���g��Y��Z�S�w�V���k�l8�z5��e=�U�[x�hOm}�{X�F��n�㞑����\ۚ��F��[H�9{p�{n��Ƌ�ڙ|�FZļ��cu"�[ɼ���)=�y�in-P��ߓ-�W�M�}�*t�w�����<u������n���,��i}:��˂�8�L�z�-ݸ]���y�O_s1ub��xm\�qs�7\�������fȹc.]�N�w�0�U(�e��uD�"v������+Ψ��[󶚮-�a-p�����\�r�����`�LR��ٷ�3�-Ϫ�q��]�̐����;^N�����������^J�[mp�/���,JgKb���#H*��%Lܽ���k#q��8�lNx�Z�/3`ˏ�)XUZ��ݱQF;E�ӟy:'��7��r�4=����Η�^F���*7��M���W�{6U@�*�1=ȓ���j�e��[��nN���YN;A*��:�*yNz�n���oG�T�7�X
cY��v�E��	��c��I�W-u��>�;u�ːs\N�zL� �r����Mni�p�~I����Z:��i�aƚX�
˲ٝo��1��";99�sm�]��:�λ�EL�%�������A�bá�*`�t]��n3q������;͠�Ӝ�V�YX���0���`�Q^;I��S)�B��)��ԼXx���x�f@2�Xf.���иf�� ���ș��j����N>��7V�T��He���p��D<�tz�0K1c�ȋ������i��ԫ�ZL4��v�s�����1�o>�d145M/��b���g��Q��u_c����~kk�J��q�!|P�\@y��KCa{�ס��<���vaa730A�ʘ�eG���̣z��U���_X�~��Wgl��PִGe0�ӳ��ņ�8.�5�]�Nَ�r����Z���r�aVXÔ	�ݐQ���a���{v��gu-�����f����Z�jb�_dX����,J\}qj�N-�X`��1��I��q�p�C�p���u�����j�3y���#�C�/-��[S�WCI������}*�q�W'g7+�)U��)8��+����; �̩8�2��!�a�,��vdzһ}8$���/c)�i9��5ջ��#Z�Y�<��6��Y���>x��+�]�%!�*e�HN9[�x�ƅe�ә帎`/+����*���vLR���BZ�-��/cF�)�V�^��|�N�>݂�&�R��u��/�%�ȃH�T�g���j^-��7��s��s];���U!�AR4�&vN�	�r�;r���(:�j��bZE#��2�C���,�f�E�yX)E۝�EoeD�!�y�c����U�~zm�Q�_Z=k������W�W����-����~93���z˂;�0H�s�d�J}�����������7y'H�Õ�{]9$ŵ�wm�B�E��z���]f��x�	�G��q+��,F��td��tk�f��x�����KJ��X�ȷm��69:ڈ.�@JWc�:�lC8���'\R�Ι���!���x�o-����/��d��x��g^ѡ9�u4=�XÊsa�T�y��پ(u!\v�rwO���g�9f� �ƏY�rOy�ɧ�1׌ ˴짂�>���<�8�`M_gk����:�0�yLIu�哇h��X�����E�ް�炇����r)�f�m�
�=e�퇝�[-WI�-q|�/����4P���G�V�"����tȶ��t�E����{���V�˕�-�Ͼ��Ge�s�✗��q@��E9=��Z��p�Z�S�A�������'8��+ktpC�$9DwNNmZBQ��R�(.IQm��K�������Y7nd�m�3R	�H'�v!)$��DS�m�'ܢ!9E��!D8S�Jgn �
,��gHP㢑��.r��u��;m�$�! ��N!([d�nq.9�6ӂ��/1����D���)'9Yh#�)��=�Nqy���$��f�N[d��mgBq$�NN�9I��� y�rD�2�ᵢ:��A�ѵ�n�-�f��3;NBY���ٳ ���.YB�ΤJk{�q:� �r��M�G)'����fY]]X��rH���jȉ�C�r�m��>�NI��z���)@��|��u��9V��޻�q:�@v���f����H.VO/OR�K�?=JUħ�����h���_X�EZ��f_#ѿ>���q�Q�)q��B��P��q��
��r)�d�5���=ӊw�����[Y2�e,�1��q®��X�N�˞�k��W<��Q���^���lM�o��Inr����������h_\'�;S֡^����v?}�\�uT򰗅�\ͪËs�k~��{�Qr�ϪG��Yĺ�G4�Ϣ��3�����nu}�;����5�z*�8c�&�P���|�r���.����N�����ǜϣ���{�%W��Q��{/�����N�+G��k�.a��>�S��nT�/Ncp\��jzb׃ًs Wc�-���������9�u�~t����y����=�fn�Ŵ���=Gog>�U�Yu2��R�#|nLce�_�Ϙ���s�3�J�0=�(�.V��kF��qZ���t9ފ���g��Lo��R�Q���c��e�U�W��a�7��y2�V�m\�W�ј-9O���ŨRy#�A���9u�;g[p$&��^dOW�xe'�Q;�5�wc�i�c�C��U�/��u]ѐ{ԇ���sN3�t0��&�v9��]��:8���vqT
Vn�`�h_m��ց�QKe�Z����U��=J��3���Y+ ��32�_�9�Ý�����Ȥ�!K�(���w�4L�4�m��>'f��Vn�z��.�P��?O�eP,�c���2�K�bF/TTJ}[}{���p��+sW(u=�*��O�&=�z��S�e	����/� �b������NC�{��O)5f�j*���^�o��[�^I�PyS&~m�\	�N���F.l�rg����hQQ�SP��9)s7>�Rb�����A�����I���'�r`[�3��Prp�Ӛ�:z��NZ8���mVQ�g�D��\jOյ����A�asp����E_�ߦx{��<(̍�t���޴��Oz#�;q%#��U�Tg��8���o�lÿ��蛎�����S��*9�G��35֝���Ȍq�v�I���y8����\yu�fl�>��.�L�Y����w��KD\v�<��I���g�~����`F����	��-�ĳ��v�
�u�Br}���*j��ݓ�l�a���0g5�3Xיݷ�CCʯHn��w�ӣ}�����~�3%I��lj�9٭&�E���_���ʟ��{{n�E��^Z���B�Q؟�]k�cu(ٮ_�p�g7d6DZѷ���Dݢi��a�+��I��1�rV�g3/�.�U�gj"D�@VV\�Φy��,y����K�hJx��F���z��~���q��k�k����;E��>�!mzg~�zD�����m�՞u���\�sܤ&��B�]H'/���֐� W��ct!L��:J�ϕƟL�?k35λ¬��yL��GV�*�pb���s[ּ��{g�}�S�t�&k���]���V!pC�Lh��k35�X���39q39,�uM��w+�d��lw�z��y����\��.d�p�q���'�1�X�_EZ�p��S�`̐o��t�:-�9��4ߋ9M���Uqv�Ǿ����\�Ë�r5�EgX�$}d�97�qL�۩I�9FL���.N�;\69����U�m�L��׋3a�1��M{FrgӮ�T�ga�������L��2)H|V�����]}�xL÷0��y�L)�׋3��l��䫪R���z�����4z
�2~^�W��3:����T�x=�,L�o��'R��g{��l���n�Mw�qNr�{�E�4����yR�*c�v_���C;��/�յ�|�hk�	K&��Of�r8���,�w����x��iH�z�ZV�\���}l(��_��Uな��V(ks��e��8{�(Э�N�`}kBC@3y��k�'�Lb:63u!U��5�醜$��X��n��ks2N��2��O�/���+\�'�Q"���ռqQ���̬%6�ʗn�0�����M�-�g
�^�_Dڣ�~��Xev��p��~J�%moc��=�<��3���gH=��l��|X�}������އ�=��;��4 �8,��n�:����y�dǖ�~��'� 
��3<z�����/2���q�7g;��p���bk�%=jY�W9�a�}w4*ߒ+Us���f,M@X����˼��&��h-��A�xg�X7?_�1�����jvղ�O?}�b��s�4vz��"���/�w`�F�Y�[�T���g	�pC�
���Q��Oږq}����Օ�GJ�ő�Drԑ�[�H�y���s���{C��L�=�'t\z��7I�d8�!q�ģ���i������=�s�w����;K�t������野m.���%B��\�j�K�j�u�}th@���Q�qL��8s��J������D'>������0�vW>H�^��
�B������{'1��Q7F��}s�iwQ�-tk��]��Y�w�k)��xʭ0�x��^�<�H+;�|M����}��h�~U��R��)�*�Lo�hv�3���SX:!��q㳂�n�a�:}�( ֑��V�G,ܫ��Pj'���(OZ��G��*wf�B��@���+�ϲ��fܒ�tq{�T�%��C�[G�������x�S�r��s.�L�Ѵ>���V��8�C��i��*���B^D=�7�a�D.����q'�+����_�j���K�Y(s>�w��-����%p
��OE_{��)Ǫg��H�Ȯ@�H�6{=�
\ʙ
_#e׫tX!S3�f]*ǽ��Mt��vk��T|������w�O	}>/�}i�ڡ=�@-꾾3��ہ�˛���1Ň4�˃��<j*d�
@mK(r�y�u";q�H�hB�d�NZ�q���V�����z�q��'�����I��nO<�u�EG�oƈ��y�?-��z6���|e��ssj����R�տ;3%���1���!ﲻ��N�`c��Ro��gW�\Vy�` K��X�o7E4�گ�%x`㊨����p������^�������ե5���&NmÙ�ʵ^[����S?c����P+T��dï_��ǏY6f"��1����U{B���E;�g�4��O%�/K��y�1�ɡ��͊����Vn��c���'E��h�'x�cƩ�̔�Ⱥ�z/\e�@{��f�9��n�=��U�7y+��;��*�*N{ٖ?*�(���y����#yMÉ�a`�7��(o��o|�5�ԗ�_Vr����E�0i��Oi������oW��N����G7�K>=>��}>:l�����w��Z������������7^d���o�S��+�Q���Q��.�&�����ٛz`~�b&�o�"�����ҧ���
-֣�P׬^���ZE�V��=��f^�u@�`�*��\mj��L�>��\Zt3�sxG��\%��Õ�S�]M%���e��� >tc8Z���Ϡ�b��}���*�|nN6\��>c�`���9VFW����L��Y9��3�N	G���OOQ�z��nDOE�Lu�)w�ܘ�S�y�M�R��7x-=���Q=���p�s��aTOMw��~~\�Ý0f Z�3+O3Q2��"3"ڼP��W�SȯC;Yôo�N^+��tP�b��x+�fx��~��@81��oĚ�3�+{4�֞����~vj#y<&]��s�2���<f!� P@j�կ����㹞z�̊�r�פ6���	�:�O<��-���)ӘR�P:���=��O��M�S����T� $jMe{�����\o.LF�I���:�Ɂo��@ Ps瑎]Rk���}���R�Ez�кt@hdEQ0c�Ƥ�[O�o#=7�\�@�H���YX+�N�?Y�K�1��������r~�޳����V6�4��%�B/�9l]Ԥq�V�fK�1T�:x�ֹ��yg���N�Q!���T�-\��vj���[�����q���;G( �<����m���s���Rap_`[��Ώ���W�od����.����Q�	��E�}��iL.R�IC=Î����e���T�˜6�oo�p��y��E�񙮸~�;y��#��
�xG�����Ggn=G-fgޓY��5���<X��l¾�E��<�C�}'�#������s�'�"�_߸��z}v"	���3Gs��8{c%Ǳi7?E���&8Lj�3�q��Ƽ��%��Ц�؎g��L����˻';�����5��iT�+����X�}����Aʆ�י�q:
������RW�C��n��ct_΋�6t�.��+�>��u����w�R��W`h�d�;2��̎\<��7헃�+����mԯ]0���E�nX��O@�3i1�}�:[�Ѣjvpgb�̪ɝ�k����}�a�_'��u���z��4����Lp�q����|Sp^=B'�&\��S����M��H�[(g����;�vz���r�ƈ��=E������D�B����L��}�D�m2��������c�N�_�\V��ߌ<�9�X@oVN�v��sv+Mg�� �q�L>x�e�v�����ɦw#���L)mU��M�b sp
�*3�嗶���fK"Q�,6�K�݋��ul�B�[*���t�%N�Ub����<��];T�W��>	�R諷�g�R�Β�f�>��z��>�2��̓��S�&�#�L��RB�_�u)��X3���.�{�	����f|�Qw-?���A,�?w����ߩ��?q�02�
���}xfu����p���{>�� �~���`����Mb䐤�d\��k=�~�RK�V�����z.¤�Յ�4W�>��Nz�:㕗O4ݼ��P`�
@��X'��Pu#ؙ>���Jޫ�QG���|�zziQ�UqgܹFˎ�٤�+�0(\7�3��`�Q�*z�D�gq��(���z<"����6U�7S���'�u~�cM���UB:�W�u���goȍ'�,5@��!���}&�5�S���Ьq]��[���S�:M˛���qy�2��_���1�2��hK������/�9�Un��)>�wBk����N��dm�s�:x��T�ȸ�}ެ�*3������L�Rt�W��W�%ж��̿�z�u����!�z\��F{���Np�PA�B߷��\��[��^t+y^�[9={���bg����;��=E��8�Ϩ~�+�u���~u/a7YL~9�W��c�ht���'t�8�k��9`%.Й�vٚ�eB;ݺ��=�A��{/�%����]�b-!�X����,JV���F�%��h	�x��X���r�'\Pr�n���j�mV��gLͫ�\<<�����������g�Fu>qK��S���~.S�9�tTK�.;�P�g��h���� +��%Mվ��-8��=?[�O���s=	ϸ<��^�2�vW��@���i����c�
�3\���[��A՚ʠ���DICvb�ďEwt�2�W������^�u��x�H]�s���[6o/{R�@�GQ�Wxl��h��tY�LRr7̴;y���iSZ$^�{X����z6��37�Ķk��M�=FO#38
K�H��AGd�g�4e�"P�.��f��\��ߦ_c�Sk}�
�o�-O������g�{�K�����˭����zx�`���
4lP)N&�}�z �����js���U�L����dy�F�L�-�X����#����B�����18�
3�w�N��x��L���� ږP��{�[��L�F�ε�{/��o��:)�A�W���^z����~�~��^��c2��&O�P)��lc��أ����wp��]�%1��b,�����������jOc3�I�L�1pps�Q���:�ٚ� �A��Y��8�z.l����a���v��]c}��޾5��ǟ������ԙ��4l�qؼ�Wq���ċ�&Q�b.�S�bԭ�.��ϠV��p��[�S�7�^��/�mdPiS�.��/.	�f*J�����&վ\�����_����+�-tFz^W�q=�.vv�9���2��P�{���o,[�q��i�<^?o
�������*j�k2a�UF�Ǭ�69��g�^e���,�	hʹ���Ϊ/���ؓ�y42b��KՀV�H@�:��o��!�S���Z�6s�^�P�Nۨ^�+�&Rj����1���-ڪ69��Xr�b���*H��f���P6/ћ�{ޏi>���Se���LDc�q�;�f�t�������1:�i��V�hd����1wb��0k�`i�]>S��|���p}S�hϖ�;�>��R�����_!�]�:�jcUU��4�o7A֨�ը���:�_��0[J���zV48t�?8-�s]Ϙ�{zL�޿w<U�	G��H߮Nq��t�~�@;�FOf2�<j�)����K�F}e�Y�0��Σݜ��\/��,�#܏��X\�p��c2�~\�t��=E��q����r����͉��x8ַ���,�w҅��ǘ2=І�����vz��>����+� ����e�fhʙ���"o>x�*��쨪.�E��/cF�"�6��]�f�6>5N�ٻ	���C�<D�7̪�m�Gc~�`N������J/f����՜P��]�k!��I�7�D9و�I�}v+�N7)ǯʡω�nz�KA�f]owȋ����w���`�k������+��(Θ�w9��'��<t�_���P��.�՗�m\����*�zHL������E,v��VqA'���s�5�1̪�	�I�<�=:_C&��ݥ�N���6/jPzJ!a/��]�� OAp!W��KV>�x�P�I�����q4�ٛ�����sQ�`���k���̔�p�Gٮ���w^���5Jэ};�����윆�a�s��#G������s�J��6 oa"�k@�X-����f����n'XpN����k�:w��C;��=�wQ\矼j5��[��<��|8���3ZV�tg��1^���8
�o1�Mr��iNe�P��M\w8"�i�l���7(3�&(|��IĜI�.[�'b��˦�vހ.�寑
�*4mr�T���rJ�-}4��N׉��Ȼ����o�9 ]^8 ���0��������x��֍薣J�+q�xq�Nm�h)��9�5�E~J��S��k ��j]&=�:���o{h�>d�R�3s4���t��n������<.��+�*�εM*/��Χ*���V��{9i�z�H��{r3.k��d�YsO������<r�/�:f�'$Jha�Sta�vx����H!5��L�x�V��nS]��D�����Y�)g8]j���]�T�u�����8U�h�M��J���l��'�y�T��ǻ7�{9<E>��-���ܓ�7��i>�*b4���EJ�`�_i�ފ��֙u�'���kޥz��kJ�	�0e%�]&瓒�Ep�:����ݬ�k,J+��m��7���te�҆�G�7�3x:7̥�~:p��{�zi��}Q�pi�6���פ>�W����J���m���&F\�6����8Uѐev,,��;$֕����\Kpe��N���`>����"~�����;���]�
9�qw�μ���0�\8�;�.���ёp�$N�{��r�I/U|�}���BO"���xH�].��+����.���%W{�w��R��ת`�+�ؐ��c|�ɋg!O�����>~>�GxK(ZF��W�͸�]���+1��q[���Im����Fv9�܋hZ��1��ύ�ݢ�(��.���<9�Fn��K:x��1�,ɒ���8-Zx��&��b�e��%��õ�5N޽�<��H��3<���L���2�ʳ=�n���SeYų4�E}��+�!�<��s���<J��%~��Ϝ��7�Ir���4UV/%���3O��o�F��i��,Ԍ�reݾ��)tBGbu6՘_U̫�dq*��ts�gF��g�^v��-^����<sf��m#�8��"s�J�lkmm��b�^i���l��rrY��8�I�M�gi����!���ԭ�z���/l��l\�6���nN���H"õ6�9���pl]�9�N:m�s����gZ@�9"8t�f��9N$2��=�G^76��NG3N�rP���mi�Qd�n�BN���N�8聛�p��FZ��9N)Fݬ�m�֓��΋9�Nm�I�'Dy�Oh�3s�gk-e���٠�B��wgo5�4]��.2����>m:S�ϊ��������8��\��n���Á%m��g8H綐����P��X`��:;�v��i�-p��7q^V��uɡKjv�n�AZy��uC�͜�	{ .�.}}�ҽv{O�W��ZJh�'ޝ_�<���������z}�!:�q���mx�
���3� �d'p�����/-��@�(?�U���l�����[��גx�Tɘm�\	N��a
���=�]S��|�)y��n$��}�|^o.Ln�Ԙ���<�u���.�Ֆ�;q_�U����K+wIq`8u[Pedˠ��Q=7�[O�o#=7��_A�2u,I�W�W��d:Y�:t��x
vK�q^/E�|��Ҙ��Az�%Ꭰ��ǏY~3����\ �cD_[�Gپ����j'E��2ȸ��35��fv��#ߑ�&<���C�O����P���>'ُQl�Fg/8<�xd��M��Hx#��Z�گI�D~�fz���8�i2�q�o;�#�/�?E�g.��=���Y76��y1�cW\���8�c^gv����?<��Yp!ǌ[�k�{��!N�Zb�Z��|r�����\�c="{��O|�{�ϼ�'�W]������)���Lͯ\�=��1����GR�{*#�ctxS0t�(Yu3�z}3(Ƴ3�w�~�x09A6<Q4�ņ��\�#Ix�G�1�|6���d,��Vl���ױh̞��g6)���ϮOQA�����6e�:9���R��r��WD���,eU)hV�-�������|'�!���<-9�zsيg��|}5U���e�rԹ��r��\ч�q75.�W�#�}^7/Gl6�����R�=��x�3ŕފ@����f-&7��2���L����i<+c����ε�J�;���~.hl�2xs��5X�4�3��E׮&}nyf䓅n�I��[^˸�5���S}0�\]� �x��9��0�Ԩ��Y�\]�,����ݨ�Tߨɔ��.O��;\7��,�w�
�9̳�׋+o�1ړjd5�9׿������jz�t�ͯx��	��ʹ�W���zw!3�����gW8�E,�������jp�;^:f+���1G�h����aW��x�o��[�/Yڦ����f�֍�ܶ���u��am:�y#��|��Ƣ�|^�B��T�}Vt)����)�ɧ&}p�p��^��֏�,�|r}#�T�m԰ew��R=�R6C�B&ު��^H��[��o�ر4�8���SP�v�@�u6��f{��ɓ�y�LG��ј�l����+�{�|@�H��V����!O���d�m=M�����;mעG\/Y��"4L�����Ĵw��?]�:��;�c��F*63:�c�hd�Zڰ�:�PT�d*�8d�72�F���/U��ԌL:c}���U��tX��P��@�ae�7��R�9�v�L�s���"��ve�XD0\V缶���f&��Mۇh,S\r�$�3u)�|t�Kt�s�爪pJ�Ί�6'�r�r����^+�N�+��)ees��B�e<�s7��FeN���vw䏞W�[?3���:w��[#v��r����L��}ޣ�z�_����x�x��z����{��Y�[��000��ӄ�~v�39�L�9���j����=������m��c��#��ɱm*���Lz}~��:C�/ew����{��q��|�G�M{��3]��&��0�N�C��~���D_��	�d�ǁ.u�`�����ڽ�����y���V�|��P.+�̡?o?s5	ϸ<����-�eq����Q)<����5R�\Z;�O�wт����5��P��%ًs=��
k��YM���Ui�_)|�J�Ӿ�^�u�fْ�ma%_΋�<+�٠5JW�LtAUrc|�C�9����sb�To0�_�jU������6�x�1\��k��=�����(�Ӳ/�����y�b�[%� /I��Jr��3�љ����N��ۚ�o�-Mr o)�!����=�2�����Pjz�G�Ŏ�r����J7a��YQ�R�%F�29�	D�ˤ�#j�TD%V#�m��{�)�>��1�1΋3aX3�B�eD-gly���Yљ�r���,�|�@ǻ��v�ߕ}��m	v����K����Խ[�mfNB۽͂�bŶ\�^�=�=���>7�WL���u�L�h®���r����/{+�a�j���U��w��1���5��L�aHߩ�$ѵ�������n��1c�����*��3yy��a�y^{l�R�}��+I����z'���1��f�i���k|*w�ۺe�.{�>�S'ǵ؋??�eկy���'khm�L���W�^��Rs�� �p���1'�]P1�O�@g���tYG�8��1�˛��n��џ*��{S5�{��|�*7�@ۣ.������r�g羴���ʁZ��ɇ_z�vgǬ�6��B��E�jG�J��=�˧���F��3߀�i�ǲ�M�n��W��d���B��g	��α�S����g/\<�p�9DS�C�ҳ����ٯ��O�-�7:������޺��$N8fƟA��%yw�z�r��8������� ��1������k���<4���Ʌ�Z^N��^��{R��{ޣ���X3���]K
�6��_Ѯ������ar���z}�<�ޓ��,��i���O7�ݑC�I��lG�3v������/���JQV{�H��d�/�P�.A�]���N���xt��wr�s�w��٢�8v��Wn��r��c#�c� �����|�Ɵ��)�ش�����Y����+r��6+��{Tg�!]��엶a���S5=N�v��1~���ύV!S)��jT�����4�������/s�k������+�a	z���3�J�dp���t��^���ŝ1u���&7�DJZ:��ѱ*�7�jō��̜����=�#܏��<v��>�X�ffS��2b8s�-u��}Ss�Ed�r����rˉ��n7'z��s��=��v����.G�F8�A�2�ȧ�����(��כ�ѩ�`�5
`�SFCs��10z���u�������S���h�V���iy]f[���i���({�O��H���X�$�ʙ3�nb�V�<�c��ɇ��Y����*�k��7j8�J��Ԍ�غ�=�B\��I�^<*mz����w���y�\|�qz8\`�����8Q/	)XiGY��E�n���!>j�u��;�뙬�{ڋ��0T�\W�K�sϽM)��Az�^�*�q��_�����隞�Q�Q�X�g���l
Z��{8z8هs'E�k3,���35��goȌ~GhT�<!���s���D��S7��^1~���T�S�0U�l�]�Y}ywj�ĵض������D��"זV���T�"�h�=~z�J-��^�vxS���{#ݹ�P�%17g>c9^s/0�R�ɵf��k0����6ޤ&jA�隑��9�[�Q-�ˉF�u/�~���6W�F�0�{Dv�+X_>'�{?~�p�j�����0'��AН[��pl5vW���}�`EK�[����6�6��{�9ߕ=��w�Gz��[W��l^����Օ�����u�o�؎c*�[������|��ؼ��F���J��6���i���z9�,������.�z!�h�=F7E�z��7��P���� ����.��;k۲z�n��KWq��!��׳�a�Cj b�f����q�Eb8��Hz�����Z����h� ��l���1�ey�ǭM���/�� ��Owj=׾��w�K��<o9?G�wQUպ�=����tة��xo��=����!���|A者�׷֩��;w���Mz����ڋ��%�2e:F��y��ΧG���g?]�G�H�I��;k��q��KE���\���x�Zʟ��9?R���{s�5��7��Qʨ_��1O\s���������)!A��u1>w�����Xϴ����`g����A��[5�:_�J���z��o~V��vFj���;cw����.���;4��]��]��T�/�;�}X�'e� ��A^�<��Ŕ}���݆����ظ��U�
Ĳ�ݦ�;ڵ.ۜI=�:�r���ʬ�C�V�:��5�@�� �	M���m��^�\;ݡ�R�d�ϟ�	�:u
~]�S��$�5i��1YO�_�#e�_��Ԗ���=��{�j�U�lHqί܏�_���Q���n��0��҉����L��}m,�<%w�������:ή��}5��h�x
������>T,��ޠј��Y�ǔ�c��/0&�����}���F�x웍��h�<�Bv8>"ۯH�^�;y�gޏ�Q�M�����y�<�/��+�U��+l؟�ճ����_�#��'s�V?Jb+���j��)oM�We*����.���i�=�Dҿ�p�aӼ.�����>����T��}��{�
�:�곽��Nf�G9Z�2/��b{UZWw�/A��s��W�et� [6�ʎ��I\{���h�x0���1l�:�÷��P�ysh�&x���;���t��<!.��үў`J�y���q���~cXȝ%�`3^��~�.��x�
r/�i��������Jz��]�{bz�8�%V�~���X\w"��W{�Bcy�����py�^�m;+��:p���f�R~��R��*�J7�Q/I�v�N�y�S�\�۹Ae�Y�4�^e҂1XWIv��WQ������G78B�l�)Z$[�{;�+)FF.���>~>��i��p/[JJќw�}��p�0�O@�"�����%pN�2��;.�������ZW����64��ܽC4��)�i�Yb�-�6�1O��w��{\l�X^^	}w�~�����/�a\/S z��s'�s4��j��dY�L\|U\��2��2dؗ���}�).���c'�E�K�ukǌ�r7��؞��QD��;2��!��ԣ�c��o���SI��[@],�N7��0％Ϝ��E��@�5�4���.ey=Y��
�E��\��|<��z�=����!���m�1��eH���򨴀�n�p�l�'���_����58O䦚� �ꚰ�������4yS'�RjY@�M��h�/��`�n��g�%�7.SS�[�^}O��oP�V�B;��a|z'������vԯ@�i��8��������Ͼ���H�-L����Hϡ_yٙ<*����n{�{��~C����=�u+�i�Vny���3�?f��Cꔏ��x��0<�Y�1��^Tqs�b4�s���z�ܧ�q�v6
��������ސ�*�2_
����U:��øǔ;��z��ߚ�:zM[��u�X��&v�r�]؎.�T�ʘ��ژ;&��,���ݽ�.;�����G�1�������ј�~���<L�t`��D��})gz'�G�f����9JQk�� �b�O4-o:f�C�lړrbA��|2cS07@��Y:�+̍�[�yC,m*S�I;9�l�<���<���lV�D�5����\zOS�H������oV�%�����蚌|a�!\���>;���R�7:~z}��=����3�ٲ��V]�撟	�`g�na4ĵ]�̪�8�q��F����]>c2��443.wY^�۫^�E�e�����yZ9̪lQ`��v�]K
��3�q��f���*�4�u%�x�����\f�s�H߶]���f&w+MDK\����3ÿ́L���e;�MJ�q�7:�} w��>��É�*���N�p�͗��<�����Xh�-�� ��FI��w�E=j�)�pߢ�u�,1�V�Ъڜ͏=��4ٻ�Ļ=7�e?\�u�Q=5� o)_����I��e:%_�+��G��w���9��epkW�E��w�r������>6��
��J(^���j�+ �N�z�/7C��@[���-���G�sL�;;��.��S��e�6�)^��f��;���X�L��j���B�������w�߰`��$�ʙ<%��:j`פr�2n�'��l��]�h��vz�bf+���B���Y˼x�R7m͋}2�5��JǶ�s�9S6=2����`�z�"vY���'
ܚ�	�1��Ϩ�-ވ�R�@���^�>���vL�BRc,c�tk�IQ���uvv.ce�RW�{�k���V�)������i��=HZ��.}x�����u����%�+�0uŢl������i�xO8��f(z�p'�* y������Ԛ�~x����@<��؝���/w���5�+
G׋AOzX]q^1E�|��ҋ�������Tu�ʸM���ɁH�UU�;�.�q/�َ������f|O[@+��+��љ���P���g�E����˞�v�fgh��=~�h�&�Ƅ��6a��+�"�}��|O��?Y��������;��N�����n�G;�7�@��n�ۆs�:����L�5E��z8\*{p/�^����Q�J;2��_`8m�?��_��zG�ݼ�_���F
@͜��˯�Ɨ3X�H��{����(��'���^��͟uN'mP���dc��X{�d�T5�3�^�+KMǹ �o��g49�����#q[���?��aS�v��L��G/qs�xj{���[5�xS1�"����Tm�Y��tMG��z.��ԡ�
˴�t���q[ɍd�-��'f��3�_����3Q�ޟx��ᵌwS:��irh�e�6�����RKE�p2���f�s��,�8)'4���
�q'��[�Y������ �.�G^C�˕S�j�����xn(��9Lj�^[]���{V%���'���q�yѾ�Z��=d>�/gJ�o]��U����Ew�鲹��#k[]��\���wdr�ꚵ:����;�0[�.�+��;� ��FFtz��ݗr~�<��w���򢌔�e��3~�n��3덽��'�:Eb�aJ�L1�R���t#���`�ﵩ�[b�/z�*A�m�r�K��t떉G�W��#�6n��L�u��O<||_�;5��4�����fHm�BK�LS�qEd��6�RNչ"��7Zdp#��dQV������;�D��1��ų���3{��m�z��pTg q��,�{A���/C	�žP�N�;�!�Ù�\����k#��,�ǋ���8�u\�+7wO�&�k.�w&*Gն� �H}O���{'d��r��x�%\8�Pv�����dC���
��8UX�2g��4i�a>�����ޭ<���u�B-o=Y�d�u���*B���T�_=�SU�t�{�M�}�K+����f���؋�Vf5���U�-@�y#�3<xp��^�uGq֥(pA��fwF+L�Ņ�+ǕXMfTF�I.{����v(hN[��u*�8M�sh���U��H����J��jt:+	j�ʙ����0zM�����S��F�-mVJ#2���v���cw0>w8��5gd�Ϟj{����;<^t�͍��}��#�-�N���$�29���|5�q��A�iPN>���,����}:��̲Whr�Ƞi�l��ཆ̏I��J,G�Q�> �8;�a.���KZ���_KW��Z��K����a)������'k30�O��ӌ9=�ˬPG���x"F%�P4��LU��	�y�M$ee����3�٫^GS$�ʤ�[Rr������ &�g` �%�.<MK���QoLR�Z�5Jp�;�D�u$��>�i(��qg��_ k�fZ]\���W!y�ʃ`57�HL���/���m�:��$c����$�������S}L�F-O'A4��L}O��>j�!��ҽ��w�#��#��5�)���qc��QB�m+߆����T�:ib�t�rYdƝ�u��ۏ:���:��/%��9�͕]7��#�hی�*ժ�;l6Q��GA�-�zc[��{�?\o��w�/�ZM���9��]|,�7�sU2f�e	x	�g;���%7lyJ������ܓ�a`�uo�ר��vKk��6�]�lQ������fg|��\�wz�Z3�b��=�vE
!������<��5ŷ�8E�{rt�������jA4U�1�4��T��!�,�|�ʨ����_)(�u�Y��._�������������EY��.��XI@$�lt(���T�r�ܔ�{��]<��{C�c��;NN:���y�w=�9Nw��2$����3�;ΰ��C�ʐC��K�9�����_sڬ����X	Fݸ�;#�̎��|����緽���X�4{V�rrt�܆ڗ�{Ђ�����D袶�'pS�����^��t��|�aqy���egv�ͭpGYԇN�����糋���w��Μ{u�U�y[�;�N@ee�6�8�"B^�U`�ԯ��������::���:f~����Y�|�k�:�Z_���V��S���佈`z�7ӫ2q���nNVW�?��O(��o�Fq�����P���g+��a�*��A�^���g}�vbջ�}~�Jk�A�Q��}"�F�j.R^�&S�.Lo��p��B˗{0��üs�Sn}1ws.�pwxĸf�t�X@k��{@��@�Zʐw�LE)�Ƿ=�O?`�fSdQn/��gfm����Ʌf}��
[^,�W!���=��
=�\�d�x�sN0� o_�^x/3�i�5��=p�d�6�`Jt��'�Ľ=i>/|��T�
H	a�t�2�Dǲw3��xr���Z���`=C�A��)���w����=��R6�6�FoS�(���̾��	�������1�����1�O�P��f{���#_z�F}��������t��;�=(ʿ�Wh�¼vM�=M�ww�����עG\/Y���u�%Zd����uVv�3��u䏞W�z���Vٱ>�l�*��ḝ�O��2��V{�sh�*�ܱo-Ƙ�zaY{�sB�ߒ>�W�[,�0�V�{��ݧ>��<\�9�X$��[V.;�$m��Kʲ�H$�mHS�Χה2�=�5��T�7��f��;�c��V��9B��=�6��]�U�ғ`��&�O��I����{atz�=��kW�K�y�r�d���.	�jU컉���˒�Ȩ�a�σ�'d}Y= �.�N;W��'�E�U1/UZWm�@���`�:/��^33q�~n/+�y}s���O�&9,dJ�1l�:�ûg'��r�'Zθ��/�]������y��=��e�q�:<B��.4z%��5��K�����3/���x���_K�.;s���z,���?
�����[��1h�j.<�z�&w"��w��&!?�<iϵ:<�e�^�2���NǼ�5�I�b@�#^�6+ʽ�}���H�J��\\����\c>��%J�`�ulnN�n�8\�Q�!dp�</ަ ��r����t��M.��8;�>Pg��� �٥�T{�Z��w���:��Tՙ�.a��x�r7��G@�b{ O��Y�%����oϲ~�Mޚ꺚3�ם	��DzH�/��&fw����N���nj��KS�r o*Di����O������	��iE=�^�G�xa+�=�e���߬�m���*��w�O	����O#�g�r�ݽ���6��U�������~xF����<���)�S(T�����ߵ8�Ո�Mu���rL��^�u@wd�� v�F��[��-�^r"�o,*�quȄ��g;��O9Ø�{ԃ,�z���{�Խ1�rK��4]������|��e�EYg�� ��h���"�6��K��K
�X�<����:�u����b?�V��_���])�5���O���BY�i4#���#��|-�����Yp�]>�\\8u�D�o�2�6G��Lh�k�y��/�^�~���{�l�k�d���-�=����4�9��1pp_�S�$���xD�L�������{������.�^:E��A�ս���VE���}5ސ�*�k�	�z��%�*j���&G��d�X�����1�fo3a���z}~�1:�Y��~�y�1쨇�C'��lUk��Z7<H@=5�P��*$�[���M�<�-/Ųl͗E<�t������C�>����z��tt��48�/�I���q�I~��x�8�R��k٦'ʲ\��� ��1p�����{�f�����[˹k�=����:��g�i���X���,���B��m��q3X��q��j��w�p>�r7�=^�Uϒ`������_K\����3לب�U�q�O�ԩW��6��w�w�P�S��{7�Ŵ��1�������P�~��>�^\?S��:0�xs1���I�>�>�..�@dv�V���B�3)h�1�}jU�P�%L'23Iν�^3���T�d�ƺ���ߕ��Fk�?:/g�}�bz�Sޥ��GlT�n�湣��ç�ٓm��_Z��D�#x�lv��yB��!����,�B��󀘔+͍'��yI񓀁������k���ŵ^����+� �S����rC���5-MN��W�\We�YȻ�.�rw��.�tz���o��l6��T�"��!���z!�>y�	�=�&'����U�����z}�O	�v��r|kK`쬇9�늻����}�
��s��A� �=��r<¼�%﫧���Xc��g8ntY�w:��9Z�q<�]fL\	����.^h��}�;i��=HR��}2�����.�اF�P�T3GR�j�������"}^��\f(7N��閌�^%�%,����k���.;h�']��ڿ!>�͇�2V����r�VDoK��*b���ަ���H/U$�1��)�]��ّ8�i���T[�=G�<E�z�1����Y����f����Ǒ.��#�*\�qEĈ�Pg�3*���#V�pQ�ۈ5�EƇ�b4هq½�/��A�3�|O��~�f{0����^��+��~�S�}�-q��I#-�;�g=���Wg�}Z�m9��s�B�����r�=������s�'�L�N� �R�[�P> �>y��ki�q�R���� �H�m�����V���ev�v��5���]y�')Eg^��m8�r6>��ܮwE}��n�=���"�2��2���&\���{m�*��Aٕ�K��=顕���t�O=4ܿ���S����ݾ��@��r��.�!^�3_c="yM��o-:�>�-�r���O����]ʃ�O��םt��u+'���Eٖ��7IBນ�%��mV�{s�kt��g76���
1�▮�ڻ��מ��xj{���\3X�Ǩ���Ω�\�/E]$=�k3�t�C ]�'�8��
�w
�ϥ�g��_����Sq�gh<�4��ٝW�_�$�~�����w���5��Qd��2}��ܜtة�l���釕ׯ��;Zt�tߖ��yu�e���D�n��18�:�MR^��)�0g>�����t{����_7>�k\8�ڵ*���m��8a\=��N�1!�02��D�;��|��\zF�0��^�>��)7���������Ϝ�mx�\D�6 �xD]�H,vF��a�<.��vre��p���{�X�w��L�o��N�J�x�)%�!����p*q�ޯBR�A^�V>�:��Vv}w�G5���ޠ�u����`�^iE���jW#�x�G�{�9�;���!�+�ZA��an<�9ݏ3/�5�b�c����v���|�N��j�F�K:�q.5��0���9!ӷ�w��l�V��M��0m�#�_=����\O!������wU��dG�[@v)�l����Qc�I{�Bʎu	;3{��O��н��W&��>�w�����<�G;���Q���d�����5�S�bo�jr��I���/}B��ʮѳ�x��z�0���4 �c��-��H�)���K�)g_e�<��)^�i&Ls�$}��=��V1�[f�ǹ[9Q���Ѥܹ����h���}�eV�rDߥUz��Voz�}w4*ߒ>y^!l�>�1�����ݧ>�~28�k��RB�7�5࣊�x�����~�O���*�;�]��00K���t#F/[X�g�諢f}�zQ6�=���N��E�.w����9G����ݷ�9:�6w����J*}����ў����_Mߠ��,T��!ѣ�+]L�z��n.S�;>����z9�t_<*w_Q��v���i�z��K�"gTd{��V;\�o���P��~�eϺ�����Ǫ����,h�!ﭳR�:9.�Qcf�ҝ���u�*R�������f�O
�WJ���/�,l��z���C�S z�t\Ɏ�l���+�f�1�����s#T�2m �t�����f}���m�.��z_nHϼ��zo��}X9»�_�_f�` E��.���i���~�ហvN�ώ"[��i�{y��7M���bA�{;@b�ǥ�����\�]k�xg��_e<�do�*�͊��Ф���\2r�XKR��E�c1���;��fy˘u�a�3�W!y���Od	�k���53&r�¹���n�f^�GO{�,��>�	���_y��ॿx�1\��k�iYSwˣj�5~Y�Y�VG�N�c��N�� ��k���?f�	�/M~�e�(Zh�V�2@s2_�oes������O3֟${���^����S@�mߞ���<j*d�C>�&��ʢk,��녫o;�klT��=B��H���r�}JjMk+E�FS�;�%��Ѓ��a���(�$�w����.��q����1��2[��H�>Y Q���M�Zϴ�E.mHcs�&��i�����ɬb�7#��o�ƴ��Qf=F^��|��"�Q@(Xz��f~��/OТ��Hli�+���
Ļ�{'��l��+�k#��+�!�U�xd��S/}i'�AZ�=]��P�:n1�=S�n���<X��&�мi���W�_/��ϣ�O��}�-�ت�~�U��&��d�/j��������X�R*M�p�)��cC��r��\@���f���n�١���G=�[�	ۧ���mv�;Ƨ9���qA3��-伄�Y�����NK7��#��M�A����d+p��M��0`b�+�T5�͑��c��^�k:k��4�I�;�`��4��/�s���&�|��y2᥍��0��U45UyP�7G^��\h7ג�����(����6n����j1��1�<�M����7�dOY�7�����79ޏ+�So��!�<��
�͏
,���Bˡ�f׃ً�=S�ȵ��j��Ό�8O���R�!���9�u�].�#�����y͊�U�~� 7�H��5�WI^�U!Z����h���E7��y�{q�<��*}�0�.��������r�1�4t@���f�lv_�KFᨔ�;�gc=M��e���G�ެ.|��`��@�m��1gT�d�W-H��n�B}c6�\N״Y��$)}��O�p��,�}�+<�<{�kʥz'���˧�e�<]As�������kZ��Uɟy�}�%�{c�;��(lv�"V;	=�n���p���j&��t^�wV]���\�:�[#�y����i��޼������N��|��cë<��dOW��S����x�'��jLEe>w���cN�[�8�G{�=��'� r`[���P����t�D�D�9	{�bCa��U�>��V�[��?ږگzQ^.z�V�;PJ:�����>ٷҙ�HFgِR�>����r��o8��y�̫Y`e���m.�	[�#�X�Z�J�t�їʞdq�����v�c�[J��Մ�`�]�TV��Y���Ӛ�q��ʺ��Uy�*�(>��a�?o��'qyDN?0T���0����z.`y���+���Y�.3�9��6�N�fn�)ޜ���!����i����:/���p��f�߬���D`���#0D1v�������x��b���{N��z��i��W�E�o����'I3�%��LKј_�	�����J���}��0�����~�lK;��� ��Lp���;W�5��˴g71W�6�W��������44L<����̸k�1�$�����is>�c_q���<�S���������ԝ5��P{���󮖚��d�W�ע���{�mR�����M����l�%�L�y� m�cXʘ����B�Hvr���x�Pڇ^�O��*��E{��2�r;�V�Z���.)���>;�����������ϥ�ey���7�y��Վ�+"=���;s��~r*�+7C@�8���C�q���UK)��H;��1��&"��Y�o�IٸR �s8�\��g.s3�=�.8��O|Al��{��^�Y�KՖ.S�*�����£�bsH���U�n��;�"�j�i;��r��P��4����&�5d���/mG�s��jP���+���d�iT�[��sҞ<���]M���	%c�t�q�k6n^�e}�׬�4�ִF�C��x�)B�z���O?V�ta�Z�]���.��bV�t��������ze�x%z�;����@񥬩�c�쫟0����%;�׽X�:�X�����h����eۘVf<����f���5�̩?|���|*�ݾq��=�;�����G[I	}�Fg����^=��͊'>m�����)]�O��|h��������{O�#.$�pQ�����G��N��Ճ.���f�`=�0_ t7R��]�iF���ʩqꪫ�};���a�zU˹h��������j������������6��#)���o(��Ѿ�ټ�<�{�%и�d0��g���v�����{OA�f������tnN�I�WU��t|y6��+�8������ג/�� �c;F������&.���2�-1�>�F�K��leOC�~��r�VTs��}w4)���v4����AӼ.���aoO�j�/���d��yG���\������^҃�����KwuP�׉f_�zG-˂�P"���wݻ�����w��
x��o�ߖ���\���R/^\�8���	sj����LGo��X�=��= ���7#�3L�T��dH�Hl��t��7W�w��Ꭾ�tq=:����G�w��]���|����]C����i��Z�[�v�*k��wK�~�e��t�E��F{�Cx�~�3�m�}�x��2�d��Џ��ԧ����cy��Y����.%�C���Sj�� �b��o��]�LS<��uq>:Hc���^[��"�E_M)Ѳq6����f`�'	����H����Jմ^�yC@3<y�]�:z�%�~�9����.�x�ԗ�]s;#�bl�v��ǤJW9�>C��o�W�ɺ��[�e��S43�s1�k�𛻶:K�2Ra�c!j�Y�]���9H�.�!o8B���2�7nm�+0��чޮ-�^��Ǚ������蛈H�5��7�J	�5�%�i� �1ZM�fu[�|�J�oĕԉ�A9Ųn(/���eu���:���A�wn���ܟ^%7{�3+��C6�ދ���־���_�2�*��=�{w��,�\�=�L�815����6�*�������R[�%gw,s��ˍ k�F��+����ո��</,[
����1�H���d��I���s׃�yջ�2����YYgk�ń�3��u���5 ��YXYؠ+>sh+��<פ%��&�6��;��yl�
��*��;����c1��
�S)�v;=!3؏��m�w���܁�/f�2�kr�96.E�����EYg�ZY�A�X�]^�:`u�����;u䦯%�.�}\�a�{y�Hj �U�X-{� 
Y:l�`塩��j����w ;��a���v:6������[O��Ea�Ƹ��OeAr4�����o����7QdI��k�<#&H�*&���Y��ðk�T��ss��5��0�v�+�;�c\���tr@[�]� �4 {U�,��N«��S۾�a�Y� ����O����MきzY�~�̫['m��Xʂͪ��P�S���V��㥪�;z0�>���ǭ�5-�ٮ��/e�`l�AR�ms�;aU�U�8���Iت��9YB�v��ٯ�&�"���P��OI"��x��{\b�Vݛ�v��t&0�d�Z�:�s�wB���B7�����]%���}HX�kj���u�}5w�L�|�pꉏ'��`�AQ�P�H�JT�O�5NRN������
]�Ş�F�Q氈Dם��D8�w1n�enlC�N���u����9j�a������#X��҂�|�$����B����2��{�%�[F��p
oq��Y�Q��vxu�5����^C��"�XQ�*ի��靠�1��&v.�k6��jxY�k����ܰ���%�Vy�6�����Y��� [�e�����+M��"��m��kvaQ�7�>y��,a�DY[o�Vga˾��i�
����QY����gv���T��? $T�MUI�����{ے�ѵ�G��(V[� ������{�8�������S�m�>|�Ya^X\����z�	N�Yt9N��i^֝8��������)��Qg�� ���p����۰�3�4s���qt'����rHY��C��m���3�N8��;+m��d֯����,����^w��'���m���Ŷ�$��Q�j]��]�'��n�mI�y��f�u�n�N>>{Vd��m�E|^^vZtP[o��z���6��g^Yd�3|�o�@�G�QI���z�����y՝�5��WN��)@����$���J�2RTc��Ptʵzˏ:�w��	ؚ�j�+��Q�oѰ����茣�pt�(������k38�25.��o�së�,�x��"z�-��Ǡ�FÞ�-=Oޱl%®=U��˩j�A�W����S�	��7>��{ఞY����f烈	����g�)��������w�
,l��¦�y:嵐�1nbF*�qj'�Ǫ̽�S�Y�.��p���ʈo�2�L=�^<e�ď[��O
�6p�=j��zZN�Ds����2m�OgC��_�H���{���;Z����Q��x�W!z~�������5�3;ٰ�D�.&WO���`s>����k�����Ė�� 7���W�͝�+�<���7}������R�*~��b�X���a�z��Py����r�ϟ�����p�o�]�˩��.I����V�T*�*�P�yU��C1�}�¯pg��x��i�^��U�z�νZP�Y�4eo�C��7*���)�5��a�v�	f�B�n*������ɾͥ�Η��\}oƈ���Ԉ{�J��'��%_y�$z�羕�{f{??"�������U�(^R�mk�W��:�D��#��X�X��p��L.X��-�NG���/��natlQ�έ����2�C���o��b8��3,y��Z����sBK3�e:��1f��w�Ǽ�rv6�D;lb��2���w�֝���<�_��MI��fY�N�3��b��)�~�ȑ~��?u�JcG�Z���|!\���%3��?a�y�,Z��X׬�[����Ts^0�T��=�����v�l��������;B�����b�TT��&i���W�_/��ȏq>���H�n��R��5�	s�Zj�﫲��J��D%T4z=\zM�	�s��%�ߕCP�s6���dC�>���^���ݖ�K�n���G���筏Z��A?f3�T��5�l�S�W�}�����"Z��>B�<����]jpo>�f�xz�e�v�w�����	�hdz���xQ`͝���R½�>G�����z���=��Ÿ�vL)�g�y>�^�mܭ4�q'�9z+��לب�U��RQ��������ڬ��z��Ѧ�e���rc<˚�g�yi�����>\0�/��t��q:��3���ڼ��<�Y��o=�"�E��R�2.�K�F��z��k,p�y�c*�x:�0�'�����Ȋ��N�����)��ٯq��S�06v��Ȥ�!K�7'��~�18<����ޟ�=���m��L P���*zW��»!�b��NK<���@=/ksei%���v̊_u��>�aup��ˮ�M�<�lw=��~�����'�{_�䧍Јe��!|��L��=��� 權�T�x��b7����ېY��cZ4waAh?r���ᜡWu{�woj��g�eP:f����7�;=�ֵ
�,�>��}�.����G<L����͓حeX��}�O������U߅M�2C�3�x�1!�?V3�W<¼�%��řjf��nFf8�b���.Tɟ�sS�0�/4N�Gn|π��>F�`|�Q�*�W�5Xo�r��PŜnx���!��	�Ɂn��P���Pg��-Z�K�P�����l8��ª[��ت��ٹ��Ѷ}��������N��0��*^������~s�z��^dj�����M%ᮾ���3�2.4=4هު���������u�������-�E�����Y۔�q��Rc��bz�|�;;f�������l������0�5��R
×�V�y�9;�~�=o�<2s��T2���8��n��>�oi��{������݊��{�o��ڻO�$Ρ�t|�786]��Z7yz{��O��������z-���Mq�k�O�Nflw �2��׎`Lo���C�[��Cg�y�KMu+�}�1�<)�0�ȯd��믰�s��"�EU���uq,|9�ɔrM�`�ċO&��Vf�����
y�gs��f�t�%_:���u4̈́��W�%��ԟ0��w��^�,�s�zO�:���C�0��(�צ�$��;�����j4�q�n��6�.�/��Ԡ�$~*�u�zfWo��G:�
��A�S7>�ڼ��ǻ�u+=����"�#��[G`��4b�Y�5>����ψ��#�+�@���Y���M��ϥ�P������'D�҈ŞĖH��V�;�B��¤ �<K�?p�q���Qd��2,R�|nLc��M�����߱/o���G��{��A�uag�+$x\cDHs�~��_��{Jiw~W�0w���T��Q�����Z��<���wG��<���+��2�:��׋3a�4��z�&R��
i��sO>��zв��T�=���N�^�{}qZ,���l��DW!��G�h��y�<�:�z��ϧ/\'XS�X���Ⱦ�`����z�5�ɘm�����)�{ǔ�RK��<����w33��Y�����b�.���xT
�j�M�5���!����&=�H������l�I֯�r�-���JB�x�iH����Jޫ�Tz��D=������ߌ�{7r��p4N�
��v���d���[><v�^v����{OA�6a�w����:�jw�~��F��L �LVdL�˝�l^�)�Bq�����h���]��<�m�3�s�Y��,�����HP���#�ӳ��щ,+k��t�y�7���|�wq��4w��3�5���ޒ��ustR��p�9���}�<y����Ǻv%^����a��3��F��Xj���'�" ���
Z,O�[9X��s\��i;�����[s���Mr�VW9�a��]���.���va����zr�'��rP��&��Q���>�'�<}6���q��T=^ث犆KwuO�x�e�נ�!ꖫE�}��E�9�9'K9��g�-������bu,���9N�8}�p�����+�8O.�����~@m���t]���Ѥ8�!zJ1��Gz��m�0�N�g��9s�u{��;~I]{'�}{Cӟ[�L,�N��x�p�bP��Ֆ|��(˙A{��[k�R��F��l̿aiϘܾ^�3�i�\j_����w8k
�&��dX�J�Q�^����defc��A�<�SO̵������^�ukǌ�k�.y{���Vq�Pj��7�)��ٌM{;29Ku�>2i�>��g�5"��i���g�
�s�0�x�� oK^����yk�{ա�͚��c|�We�p�L�:}��3��Y����f����9�	��]Tϗ��~��^�.`��v���}g���u~6��2R��}g2k|��p����YH�veK!� �����.��"�IU�^�ݡ�^���ƭ�m��s:+���>�l�>�ԑ]��3�9�e0����ȫ">K��w$˸�5j��`뛥s~�--�yG����5��higu�uB��(�.V˳��,��d@~;"������{����4��7�yr��b�ZH
o���dZ@o�o�y*�P��[�5aG]��ivJE�M���r�|�ܚ���*B�t=��G��W�SRb����)���J�,��5{$�پ�=�K�a	��N�0c ��`�?y���D��`�=��o��9�ͺ�{!�gix��c{�=���r��wRc��f�!:��{�8.<�LI�˪<���π�=>�]K�I�9�7��آ�1�=���.vN�>��ƽg-���]�b�k�'�¦%ꤓ��W�Z��\��rE���?p*+<�?;���h.4?��(`Q��g�j{�{+�Cnz6�6}9Ժv�����;��V��.�������0nQ�a�!\������Gs��.�{�Ϭ�)�H�����s�|wGN{۱iܯ͑o���Ϛ�pJ��?r�a���hs~�9f|ס��H�袝S����q�]>c2���V���d��5�q�E�7h�p]Kކ��VVL�\�ꝣ ��5��x��yT4�g+�v�
��:��:�|7�I m���֫���w��̰m�@1�c7�R{�\���,�{��������=�/�ҕ=Vzu�0�Ɠ`n@���9���BWY�-�eL��ܝ-�R4��Ggh�̩���\0���	��Ν_��ez t����o*�r���)�1-�����OqQ:y�9��ZZ�������D��W	�ܡ.{�k7'.j�1�}n|�}�O�n��N�y��������hqPD�����ϒ�j%-z�.��7Q}�%�y��x9�*�`[�}X_n5������Wә?p�pf��?x�<�G�+G-^���7�h�8��@�ֿLҞW�OF��R��T�۞;��|v�Hq����=����*�'�x.}��
���~>��̲����n��u�7��u{�����Ϯ�*o�d�%� O�|��U��� �M���BF�Si�e�d�*��ؾ#߸`�ǎ�Tɖ����N��<SF�o�Gm|��S>US��m߲�gNH�s(/8}u�q�D�1��I��� ��u��1q�7.`�˦Z3�-^%��j���v��כ��~CЭ6nj+���-׸Z�4E�>�W��g�����򝸓ڌt6�k�{��b���.�'� �T���χ�pG�x����f��'E��2�f:߀Y�u��O�q���!N�����f� .Y:���gFt��:��-buvt�ɝt��$�5�9�b}�f�ܚ��<��������m�� 庹�q�90.9=��F[��qm]�D�/;��;zrX�үy��+�o��@��7:y�s׽� ��V1c�8 �pEt�[Kg/7j��r@~R�P�w�Щ>xG������O@�z��6a�
���Z���Ea�foۏ$�*7�=�}'��޳=q�����MPˏ�d~�Ï^Wgfɪ<�[�{���h������z��Acs��5�wm���0��X�߱�;����ۯ�X���~Z�|:+�{�.�w8ג7�Ǧs��';��&��ʃ�W��Cfu���h��TU��_�]�}�Mv����I�eTϕƗ3(�35�:�
��A�S7>���\�w��UV�;�-tt͛;���ѧ�$ ,{������"��Jb��үY��tثL�_�W�~�ќn�-V�:���ֹ��|��h<����2\�O3��E�>)��� ��g~�M��3�����f�Ƶf�mzx��m�<eW�U�b�|A�Wxs��7֢c�n�RdoCwp��Vd�qn<�����,�w�
�9̳�׋3�X@oLR�����`e/
K9�I��=Q��X�hj�1�Ur��/�M���N�ɟp���h�a6Qg�����B��%�j��!q�끡U���f�L���j�`T�Gcz��z���4Fسs�-�)����f�e�:������Xi���%���O���:)��^A+V�^7�^��;���CXz�%d�|�d�` ��y�+�u�=�5б�9ҋ.� "���iGꋜ��W/�~>2��?òk�[>�-�i��3b�6�`Jt����,A1g;��;������������������C������F�����w�0_ EwGQ��٘�ɝ��ڼ�z+��TT�uW*�V��W&���`�\RZo2|Nɳ�=����$K�v<̞���	��&O20I��O�hx.�Fz��h�ϋ���T��kӵ�<#>��2*)Սµ��רÍ��f5�d��{�d��5��C�%X�PVٱ>�l������˼}~ V��q��&�M�Sى��J~�R��~�g]�
���<��~xG�8g�^>��LRK��8�^�#v��z4�s*gd_#��dyQ��p�m�LO>��Y�A��6ǂ���~r�}\��@���J��'E��
�����J'8�[��}μ����P����{� �B��k.� �F�g��s��F�t����������u|������}ru����G�/Ebά����X�����״�E�:�>���%���U]KUz���bK�����Y�3�Ѓk�<�O��
7y�E=�@���s(�N�n��\|�����8o���&/h�o�:/��+Y�n,�6��b},ѽ���3x����o<����Z�fu vֿh�]�S��XyiqM�с/sdc���V �4z�qR����MέB�f��r�Jw���׏�2�~��;�i�\j_y�T��WTT�'A��=�z��]�}V�8��=�<6��]�Zʆ�a�5���׏��\�/pq�)5.c�ᳱQ*e��K��5JWg�n_��Ur~�2��f|:]�B�<��:��^<f��n�}q���{2�����8�V\�&ӳ>I����.�;'�����&fw���8���	�&�`_1B���,���=����@�1��q�19O¢T��]l�>=��������:_��}�k��v��=��*���\H
n�?:�&WD�b�V<P��MXQދ�<9�tg��K�צ�f�4ۛ'��<N8g�jYB�{������F�kB�m���հ:�<�˙�>�S��ȹ������'��dx�'�<>�qH�>S"��C�{"���e��Uyڜ�b���O��CD�缇�+���&>�%�[˪��,�"�`Լ��~�w%>S�����!��gN��e��z�����X7ސ�*����|*br"-б'��^ߩ�mP������{;�d����(�v��ٸZ�sjk�W�Z�g�ne9YV΃�f�XN�dU�P[�`Syn�7��L��y��XÔ��uc 'oe�=9N������1��Vf<�X�KY7�O������Í�]}����-�i�m�5�Y�srU��.WlX*�W׎�R��&.l�D/�^ӿ�wt��Gπ�V�!��7Yb��g7�s�Z����a�r���[���ɵ'_$�a}E�i�e��bqq繪�3ڻ�����}�P@�%w-�R�	%�O�p�?��I����I���u���+�%
w@XS=���Wh��ww��)-�s����k{6fvR�@F�Fد)�i%S�345���V����j�,]?�0�dI���\�>ﯞu�m�)ֳ+YD�O4.�cr]d�҆��^P�m�ޜ쪃	�]H�ő��m�6��#h	�/L�ymt���p_.̃6e��|<�������\��'fF�88����~� 9��V����2"�4CG��ۭ�*�p��
���OA+|�Qݍ����jcw�n�on�3,�P@�=d�{A�Ò��y��3����.����T�#�>4���2!�������Y�mf�Y�ye��i�j:��ipBb��d2�,�n�RZU�3�.Y\A�CP�@_E��kY�z`�I��l���܇�+n�/+�=FW��6�����X����u��Y��nK��Wٙ!w(_V!mj�r#m�p���Z��������Y�n=D
y@5����l��'ʃ���P��)��zɾ�4��+�S�}:�nᬀWtYǹ��E�K��xG>�uj,).��j��v�m]u�Z����EM})*���>�����T۬ϳ\���+x�]1��;�<���D���z'�l�ag�LxE͔P��^ӛ�d{sb��%ƛ��M���<a��)6+��)�L#�(���Ӣ_�W�m�%��}�Q]�w��1��.8S
WP�k����� �ؓ�(�Gu�GZ$�;3\��gY֏q��Y�p�@]}[d��̴��t��[s^�}ǈB�Ɉ%�ģ�I�N���gf��D��Ӆ�q�]�Pffl���`B�&�)��ЛS�J�'5Pus�cɻ�u������R���->�5b7�`e͐��e<��I��e��uYκC�(FH�B�`y���B�;:���oim���F���Si�B�39�;��T�o���K6�[��!������1-J���V�1l
e�L���J���Sc��ݕ�6�Y5cT�s7��o�8�>[8���г������	��,�*�C�LEt^�s|zv�{y��9&��9a�1�{G�"�5��,�o
Fյ�˗F*�;B�6�ɧ�
�&V�h�v�L[��:��s윲9��&���)�{�
�o��6^�[j��}�sF��ч�gy���n��|�tVVBw�۩��^^z��my��n�p��#�;��<���,��vr��,��m=���z�h�5�-��yH�;��k�;%�k����i��(rma3'�`�wz[�6�r�=���-8�l[��G�w�+m;��f�cvv��޽흹Qu9�pu��=�zЌ�3I,�0�[F[k����H��e���6�[[��qէYy�Ǒ�x�,ĝ�Y6�99����sh�.��9	-�Ml;)kCm�嗝��q@A:9e�f�:���N��m��]m�m��n\��k�:ڙ;�-�Ы�I�@Rާ�^*�gS���}����cx ��θ�siʾ�}�b苝��s3��+���r�_�����M�������ԝ�ր�v!�>����>=R�~��QZՏ\��96��
��u(S�=&���~E�q5��^���.�ü�Ꜽ�K�/��v��������0��g7y+4��g}���^6�dY��Q���s��y������W�{�G�D�#�~��{���J�=�C"V�ׅd���E�6v��z�x47�4�/\��޵�C}�Q�w� QO����|�Hon9Ni����C��tc��T��+�=�EB�ܯvfؚt3E��@s��6����5�wɖ�<-R��%;Ш�_���a���ݪ4�Q��?B������0@R�j79��Έ�X��G�ѿe�E��0��s3�oH��D���Z���z#�;�s��\H?B��Q�?oS�\,���x�SuPnYCT%\��ۖ;я���{}<z�T3]i�����P+�kZ� �b�2����.�nO��Q�1Y��"<1�"�p���m�]�T�2C�3�x�?H|*LV3�A�^�r}�ĕ"��grڙ���r���Mllthx_���-���޹~�^yKO��0k>����iۖ�[���zwzc�.�c/ˣ�,��bӕ����7�".���@���g�m��_^;k����.�;�ǚ���<��Vn�5���S��p��}����S�dVɘ�������)�r�Fao�Gm3�4jv
z�v���z/=�o-�y��R��qu�z�x������x���;�bb��7N��˦Z.;q��N��;�ݨ�7�&����T�\jLV���Ȍ0��asp��|ϤU���g���3��y���M]���2a��e��p~���W!� T��wEK��:#C�tه}�t\Gk3>"�j��O��>�o���W��5�{fv���*O���(VϮ:1a6l{��qה���z^�p�'M��w�y�A�3���Og�Y�����NG���~��`v��/��ļ�	>�s1�����*$���l>�[��נ�k�f��3���0lC˹�_7~�s.�� gsٞ^Pwp����GO;���oE9���A�0?`#�cΘ��[T�P{��*1:�i��d�{4� 0'���j+w�ϧдX�`���\Tϕ���2�k35λ® ��yL��Gl/
�f1+�`����^e�h:м���>�c��+�Jb�j�+]L�c�ʕ���н/5Rv���ӵ&��:ՙ��/���\��Z
y���8�5�0�(K����{���Bd�ܨ
�X���3%�Kqa�I�a��L\OQ}��CEܻ���׽��μ7���Ŕ��b��U�M�����!n��\2�72s��7#�.ԍ�;եΥYA{�� l�2c�;��-TUz�� �|n](.�rp�+��y�<r�o�2��.��h��E̘��ȹ�����kƏQ78�Z�h�me�á���1#����ΧG�=������x\C٩��R��������L��Xz��Wo��{e0{M)�ǵX���Q�xL�[�Vf<����fb��(W��+V���ȍE��5����A�v��+¦a��x��y�����3b�m��t�T��6ꏭ�^�y୺�����p��Ɓ(phԌ�l���q�5�#��~�z���~B�8��P�wP�]n�=`7U:�,���V���iH�z�\%oUɪ=f�1�I"��K:�9W���r���Z�g{��1�F	0��2�|Y���9`�+��{OQ�FjmQ3O��7~���;ډ���t&7���~�>0���e$k�����c���6
�C9c�~v��;������	�����]sX�9)��,��s��{���yi�=�D�EӘ������0``AZ����FGC�!�띞XY�YX�R7�T#r�2��!��{\�}�p�I����D�2�L���"w%�F�Em�/�y<޲q�V����D4WE��P8�}Mr/'I w��+������p���)B�7�m����B��+)���s�h$�,��:_墦,\j��\�k����`�o�5_=^ت*0��E9��%I���󽻧�_�U��с���\8N�#�m9��mzR��&�;��}�T#���p3�����]z�}v�^|�x�ϼN�Qw��:,��/C�G�ff�����J�d���Mڌ�ܬ�$��W���ߛ�.����
r/�i��������;@Z��.��ٯΨ���d!|���%Y]��n��<(N7�f�9����fN��_K� zyz�`+�eh����nEy�M%8���8���ۘ���0�+��X�z�4u�}0�.#ަ ��.g�<4;��K*3Y�no�C�65E�{��4�j�mӜ�Y�����&|c�8ar�c�*�9W$�j�B��ne����:��%s3��ߍR��>��K����p΄���\{Y���~�x)�?��F.9�r����B��S2�YBP��Ę���W!K�5*�&��^���tf�9�+�55X<}�N���F.���G·�d����|��|;}�%]��ީ�
;��<+��e~��D^�O�|w(ri���:Om=��v>r���̴����&A����V�֬�㍶�wk��VqΕ��N�f�0�u���h9�.����\1Q��)x0h��yӓ��c��Fʏ$�\�y��r��ҏ�3@�ۑ����NZ�OS>�<߫¦��H�-dx�s�SRkYRcaÜ��&*���>��������Gi4#���=�MEǢ=�0L�<>�R$��щ�,s�zl��ݬ�w?{7s���p��ٙ<*�Hccs�Cѕ��w���91V6#�tğ<���N�*�xn��\j����ȪpJ���z졶z�=�ů.ʣ�oÏ����Ts^��޽�n)��۩��͋�ʬ���~���z��Z̘u���e�hݞg�~�p�Iؿ�x���\���#=�L޿RW����;χ���?o\ت���%
�hi�jǪ=��pC�.48��q��뎞�w��ο.�q��&U:�L�J[����Ǹݜ��Y���,���AꚏEN8]����
S���|�郭c03��f�]>c2���V���Y=��q�E�5�ֈ��'W�Ì`)jp|H�S��џ+����>�ҋN��\�Ƀ�B����!� �v�$��eM��WwV�[���W�)�ޟcC�J��m�5xϘ�Ex���gOK�5+�*�ii�o�1�Ĵ�Z�[�D������f B�W�s��0'���B�U<�!�[GH��9x����k;��R�\��k�s�{�Jaڶ�g��E����1�c�kE�K�}(�a;u+[�-�CRC�,O�g13S�#�Ww3���)����Ӕ;,�l���u��%�j�OK^���ŝ1h�~I��QuJ^�3��lnk,pO�ޔc�C��6�
�Z�a��q�r��`����N�<i̞�hx*B��җn^qI����]�-D��R��h�������B�^�����4��{�o�g�@�j��o���%��U�ol��>���\�=�`e.����g�na\�̲���x�Ѐ}1G�o��ag_�:�S�Ǯ�	�.�LRi�/�O$�<��?6�.�t��6��#�o�g\��i�c?mГw7�x��h:�k4��Y��F����Ԙ���<�^��d1q�'�:ukv�nBs�fU��T�N���h�T�c*�鰸Ԙ�����Fz��.o��h�}"�>�����"g�r�cQ�qG��t���ع����4�)ꤗ�:�wE�G��x7M�}�߷����}S�R\��d-u3[;~D`�j�P�}^,�"�9����.�l͞g�{��F�g���ebk�����KD_k��c�}'����G��|2s��T2��� �OW_�	v�u#���wR��@�a=�~�y������C�[�n���;]wmX0�1p���ϊX
���a����msr��=����6��~�Q)��Q���X���n:��Ζ #�Ftg��y�uo�;���k���5fA˃���W�r@��ԧwd���L}���lO&��u���s��)��{44O�.�t������F٦�9����S]�{��Ei~k�����Q]�z1�L	�{�����U�T6~��t�ق�}��/u����@+ޣ�
f�%��g��O�e�fk�u�J�|����6��t�Evߪ�-sۻ)й�5+а����c�����"�!Ħ/j�*�Y��tت��K�ƌ�o�lo{�]�$���^g�cǭM�y����\��\Ɏ�7 �b��'�1�X�7Z��Gu<�k���~"i<(LS~,�|��=���{�\�;"C�Qs'�"�F����(j+T=�#gG�Z��r����s=ϧp�g!e��B��s,ì8G���je<�S�"���{�O��)����@j�pi�>��C`�����}�^?\�[���z�������%�ӿ)uy}��XZ I�)�__�fu����j��8G��8�������w��׼�b^��S$*�����j-!��^�D*]�@����t�����H|�ّ� ���B��X�Y5b�`Z{Q�+���
������e�}~*�O9�3`<V.�r�DV֮��@2�8&w.$Ru&��]�S/�E���v�Hf�c�|�᪄��Y}�٩�#�::OmgU����弟�m)Ƈ<n�ͱ�s���|I�i�Q��^��Êj������p7AH3jX3Lߪ��!��W}>F(�V�V�ȌF�D7{�1g�zkgI�헾���T�:�� w�|h�|��2�|YڈEzz�]t��S��&S�C��^g�S��I��g�P�ɡ/�BӯD�_��fޣD��;�>����c�v����.`���Y���<�g+����8N'sX�9)��R�ʎs�0��hT=�$|}��\r��x�]�^槼&��b=�N���}�Ϥ����S;"�w�=���|�P·�G2GU�{�S��7��������Wv����g	�R����
�y�'8����l�h���V 7n�z|��7�x;�G'���{=��gs��<)�:t�C���ĭu3�g_�P��/�{m�f�9�5.���1�p�n_��()W�4��N�߁.w �b��%���7��Ng�aح7��=h|��?6P��y�����\r�il�+�Ǳ�!�:9.�Qcg�O�i佣;�i/D�\��]՟X��w&1�qW��ye|�L<�kצa�3�$�.�Gg�+�~kN�X���wnlutV*���7��[҆$j<�ë�aD�U�j��|��(�v��aD����=��.q�O�z��N�6ڴ�'��]r�߰f0Р`�:�͗9�bn���h������rQ�i��UW���J�6.��.�^�"
���e��k3�OMh�N�q�p�z���ޱ��u��c�-���n�8�^W3���5J_G����9�p݄���z�U�F��+�X]�Qj�䐼�M��rx)]͟)~@����>�Aе�
�
_˭�gǸ5<d^z�=z�Q�ԥ�cüvEǟ��l�߅_���Ǻ|_*���@��/|�v(S ���4�r���AUv�E�4����N�yS'���o����h��x����8o����I*>���{��7�릁�5��~�1�������_q�T6��*#��]"D�n��a��cvK����K�A�~�*ߝ�����-����!茮�~S���Ǩ��O׃q54x\6j�SSם��E��^!����f`�h�g�\�6\�z���T�TC�s��<��8�)�d5y��}�P��l��s����P+T�5�0�=~�3��M���3�f��vg�:���f=�P��_�����^�i<���vzE�w6*�_��*]J�Nɳ��������'"�ph�P������p|z�ٛ|�1 ) ;����lC{f��;t�m���8PShaտc�ow�Y������p����Г��]5;���of#H�#:� �k{��#Î!6��A�}�z�2�̣p�ޠ�f�2V�o'��s�)R[����;)�6���c�>���+����wGNG��uö<H�?x"�٬#e�o�J����~��rӌ8���03��K���Ϲ��ιZzM��ԝ��z�F�as���t�0��:.
��W�w5��aO�ݼ�)+\昖���]29u�z+]�75�t�I���Ea�^�	���g�����|b��˚N�ǜEx���O� R���I^��2Nw?;��sZ8��Ȟ⣠\bΘ��P�&3MD��g�~�L���\иa���\ywfmy�=��~c*�x:¨���@�Sˀ�a�p.'i�"���](�{�lt�ޓ�sJ���{o���;��9.a߈�G?O��T3]i��+ލ���@�5�B(.vdW���2*	���\����g}��g�2�p�\V���r$������7�89��d�y^�������pN �@w�b��+��Py[%��	ӘS���G]C��3��i�3���镎3*H�5#�l������MF�:�!�B1s?�>�ﾏ���x����뻿��뻺뻿������]��u����ww]ww�k�������������뻺뻿�������+������z������wwu�w~Www]wv������w]��]��J������������wwu�wֻ��뻿⻻�뻿������ww]ww��(+$�k<�c�yc{0
 ��d��H���R*(�R�IH* QTU(�R�(J�QD�P�
�B�
P

�
P���!IV�*�
U"J�m�Ԣ��m�T��d���*��E�f�;�IH�
5�mf�K�*�V�ѪcFe[J�1D'\\��Z�J�T�#mK��]�-���H�m���KY��1�l��Z�*�Ѭ�Ҕ�5j����[imKImVfjk-�-�l��ٚmf�lEmkdke(��IJ���i�wv�v��ֳZQ��  }�}� �4gM �\�6� o�qv�U�s�zj��iX4�A�q��A�W����A��pi^��s� ݉ZٶXV�4�;�meV�l�  7_}A��-���f-�(����E��:�(��o���  �_^�QEQEy��PQEQE�M�P �zz����(t�N�-����u�s�v����� �l�  9_��]#���v��h��{��v�u��؇=3F�P{�:սr�eݶ���{Gg]��r3M4kgqӵAJ���p���ك[Mj�H:����il����6��Zh��U��   ��^��ݴ����ml�i�f�Ԛ�m!�ѧT/a�&R����=yB�mg��[f5�f��5���zn��v�����k�U)�zݬ*��Y��R�Kb��΍Z��   y�J���L�i"� �}��k(on��t�ν��كE��
ۭբ�u;��Ƣ���]��R�oo\/T�^���Lt���K�fݲ�jIݝ{��J��[e���RB��w���  tW�m �Դ�;���D��Ү��JSg�ǔ=VJ��+5%�)+u\�۫���jqǮ�wq�j흠����ZY6�u�R!�vҠS�i^�j�����ic*ͭd�KY�  1�_VԔ�]Ƨ�N������뵩v�}�n��Kk�wB��R�]4ۊ]N�n���Nҧ����u����]��׭L�V:�u�lwmv�*�ؽ۱��XW�݌�eV��5le��  .+����i�hvnm�4͵�����\82�J���n�:M+l��3k.惥��&��IsZ۲̪�w�ɺ�\��*���[k�zj�m���kI�ڒ�6��S�  �}�����6��4�5��e����:6��wcTQ+5����5Bq��ӊ��jWm4ݥ-]+�^�\퓵m�N��V/@�w��[k[36�i�����ޭ�j�  ��T���u=;��ըa�EQ[�\R����G�N
F�VTը�硅 {+ٜ� �G�^�{����T��h�)�IJR   j��i*U2`  "����@ 4 j���UE  �&�ʩ�  �������W_���,�X�L�Ի+g�
�/�o�=��1���c���$�5���$�		�	!I���$��B�!������kο�����g[�RS)�QQf���X�Ws��]�9�=�Q�l,�'e`ܓ��g��{,;[�E�
N&�C����{���|�T��!�6�xq�ha��%v�F�5 g]F�=��.�L�-�r���4��.��`+R+��o�Yz1����Z�J	�9+��/�F�)��%����Vm��>*Ѱv�͏t���2ÊRo���-ߋ��K��ӏ~%{u����r[W����;�u�a�D WZ�+��[+r��Kr�ۑ�����q���W���ȍ��nmS�cŝV�ޓ�b�	���9܋w&�4c���)*)�W֎e�)�S+sC��
n��iՋ:PY��A".�m��9�4�)��-�r �m�P
�\�(�Y&$c������u8�[�"Kt�O�_J��ڨc˶E����)^�2,�D����DT�>W{}�c1v�Z��n�B���r���]Z����;v�D
Ʊ��hlބ�
�#b{ւ!ܒԜ��ђ\���Vay�	��J�PkcR�9`�.+x���^����R��6�Q�C����<q���6F�Q�vዹ���O�eoV.b�����l{�h�&��vKI焗Rn(ܑ'�4�v�h\��Z�[	�ȣ��}��V�����v2��J��H���]�p��ܟ=���{����^�������f��[b47*�oP�������,JN�H5��v�;���Mw��3qЧ�)\t6U�Z�9���F_�#�I�!�����ܝ�N����Z�Ґ]7M"P��DE8�Λ��]���Ds��+Y�Y0wЮ�������wh��q>�i%٤=�K�[���BrC������D����W+.^Ʊ�����Y�(�+�$C���I�{0Û�
sI��[��QҖ���[z6n,.��F���K(RY���D���8��1N�����V�WF��+R��*�졫`�N[NF��Kq+��1'vp�H��X�R�:�4�$*w{hD����ն4A�3c�nñ��Y�x��e#T�p(���n>4�/��ɗFA2Jַ*��]Cq�H�L�4�h���tGwx$��CC���A��ؠ�ҡ&RX �����	��tE/%����;����|�Y�4I�~��T��h7T��d �E^�8%�� �]9@ �y��Aq]"�r�pcO���*7bǹÃa���JSCL��1�Îͱ�j�̵�Ӽojc��Gr���P�d,T�fļ��L�/)71-w���I������J:������d�a\I'e�֭���7�<���-b�x��ǚ���h'$ �l�7�4����0V��|��o.�.���WL�qnQ�W�fwr�A�њ_<9=UvdCu�ٖ�FqL�X�ۜ+�O�dg.� /��V��F,[m��S'{��cv�^�eBp�b��cT I��V�p�i Y�L�j��*<â#B�T�5���	ف3��;W)�:��h&ɵ@f$�@��l������.�u]�%��[�g&�<ݬi!A��֒��ṷ8�{*j���$��5�:��c��҄���t"�i��᠅��Ҿ�է�M�̸"�li;6���4�\ކx�n���Mc�{;�ۭ���=�H�%��M&�t�t��>ˈtŇ��%R�lj�0�0�NIv��,xS�q�Ӵ�a����5^᛫�I��o"��X����t]�R�,$A���t9n�gM�����Y�Ϳa}5����!�޳k�H�[W2TrT�X�bҴ�"��82����;Nl�gm70�+'�c&�G�g(�B��ڮcгz�΃���jkh[T�w.#٭��/l�6��@�������O��{ك!ށ1.��EΗv�8+di�ّ-Xe�n@n��1k8����!��`�I��YQ%{� ����&2�|�i\m��Mvo�8)�4���Y���LYP9Vڲ�:�>(��ςa�T-��N��2"����pz%�	uZc�wOJ/'�^�����=����;Ak&���9t����\�D�!F��l�.��҄
�P�.G�M�!1���v-s^���$V�dcZvE��V��͑	I�˚鼨/u�A�ւ����Q��m*�ݼC:I\7~<��$VJh�2��"	[�eZ)��(��Q��Cgj�̋�c=����d&�����q�Z�WHn�v� �w�����'�	�m�
�8�SS���B�|D���zo����k�,��g;�M���rs�
�+]�N�����ǌ7v"�1ǱVd	�KD�X�)7�u�.��
l5��d���!ˣ�Tz�t��9M��7��䜴���Ҷ!��[����q�;�M�n�=�Bl��)#��6�:�`bxV�K�a���[ �3��f.^{���]Ӕ�ou9y�K�0�}G#213J
^H�7�Q7�<	�#�;e��ى=�:��ٳ7t�7�-u}e8��E��.���D��wv��3W�3����%&t�%`hHR�ۛs����n��t ܖ�$U�8��ÉƇ\��:oM�A��b9){�xkZ��VD.h�Z\���eQͫ;J�=v�dI��4$j7�+�r�Lי��R��T-sҘy&* ebۭ5u{�V�%����.G%�E��X��_҅-Xn�[��1e�-O!�9�s�C�*j94�byDű���$��l�$�A��k;��I<#��E���!5�w��T�c�V
ח�^�WB���V�Jl���oYj��C�Mu�rv��R���fo:ac#V�̂�2:�\u|�է���d=����A���WQ0h��C0-�b���v�ƾ�ag�K��݅7��Ѩ�]٩oS¦5;왝��n��H�(0\�Edl��,���ۄ[��Z�8�ЂC��gL�wp�fp�&ۏ���p>�,�G>j�.;�I5w[�k�[�I�w(nw|rY�j"��^���"cb��hR�ғ�n�-rD��˟�	�ě���_n�L[/��Z�3��5j�0t-+�-�=����U�Ǎ8��M�V@KW�cg�����'��h�U@�T-��5&c��U`<�\�j�l��L�|�3�|�H.�ü8�9�cQ	Z�e�d���|���ڵ|�=�0Y���B�.j*v�bfhx��)o��6A���V�2=a��Ꮂ�s{;�����΄����袰�r|��xf<��6������q��D,M�Ӹ��vvn	�#_P�����J��e�7v�nE�)	�ՖL�Ɋ�Ƴ�=�dT8�O(7Jf�q��1�d�.���[����(md��4�[5�cv5�ߴ�G�K:���0-bO�;�\WA@���im[`d�'��.�t0`�Rbދ��U�y.�3^�ܙc�E�=*a0�L��{NW����i�W
<���<\��ð�1�{Ft�y-� ua#�e3<"<��MA*����EA���Oм�HU��eT�;�{�ɻ�r40x��g�љ����l��ff�IЩqi�I��;RФ�;4�A�3ru/2��$�Zs���qq�M��9��-59$�Qf��V��72�d���۷7�LV�{6�M���g��M��`�Z��X&W;��cл3.j�rd/��|:<C�������a�`�ta��B�Gwa��<ŵQů|c�K�H��%6��b8�А�YZ�@��&��K�_�;��-!�����^�Ý�o"�v��ݖ��O��k�����;%�C��щ΄�&� �T��{�
�M�z嚱@����h�[j�����C ���üP����ىd��neסhQ։�q��Q�%�.����a��0�]�9\z�x���4���uc�
yF�kRz�e�gd�!8N�IUT��\ ���om@���^�v��(Cl�k|�v��grq�w�Q�⛑���]���u�*=�ta��4�Bo�䝯7�FĮ���V��i6�����j_D4���)w_�N�&'&�ʷ��N��u�P�m�E��D�T�[E�n�e�7�q���c�+��H2v��V���2J��Ө�n�|�Y��|���%���6�@e��M*��v���<��p�c�`\ŗNB���#yB�c	mǺ�%�݌���ns�<�Q�����ᚫ���7��̇v����3�D@��e�0��д#�%}��l�{��U�At5��-��N)̄���V�ۛ�7w^/E���s^���1��i:]"���QW)��Ƅ���ؤʹ���4��h����9�w.����iWQ=����X��ΕЃ�Ӥ��f��ns�I�������ܽkS 8Mq'�Įӵ��2���:�o*4+r26L:&f�6�eܺ ؁���!��ч�zW�Pyd�y�.dYmXp���#��1f
��#H��z�i��ΪccY�m��fD.!�%�s�ٮg2;z��
n�+	�N��~F����o<�H֚��wzԏ^-��;�\Q�{~K�yv ��̑�qÇO6�)\PXr�U�t��5n�{Qf�0ؔ�I��s�{2�(�x����_b-��.s���bj��;�uS��x!P �:*���(9JM\_�����0��n�+�@i��y����hԛp��wT$MS0���o�{��
2^�4fhc�c���γNj[ӡ}�a�0��ث�VE�7D©㜎��"��Z��:t\8�(ݻ�7��ʂ�(h���3XA��vn,�w�]2�JM�{	`��q�ދ%ZKaګ���K2_�����ˢ`R�<=�D5�9O�1ɫ���T&�s��U�8�7z�a���̂�1t��­��HƱ
+��Y8+���0�y�5�0��s^g�x�ȯ��x�\7H{����9��s���
z�ZҚ�O#�{E�7��MR�5����zN�U�ц��)n�Gq�ݺ��s6�v�;^�^	>�4�ހ�ERt-h�걾a�5��uE��X�ںcu��ټ6�p^bN�l�ӹy)O�ݥ�j@v)O7��]�Җ ��à�po) �r2�>n�UOuP�Yof�"}�s��L܉SP+`�M�#�y4�:��2��:#yWPIq�:,|�I]�=�lv��8�,����c$�̻��+MnB�ѳ4Ĕ��vnde����^��}:��$���Պ��|���7��κd��+6�C^2��piW�a����|ot5wE�upH�:�����v�ļ�P��	�bj��zRHA4Mgm��)H%4[b	X�똖�cך���t�-ܳ\���T��t��ِhv��ෆ����h�c��Y���5���P���8�sS���`�~o����ށÙ��o���k#wO��Qǖ1��ʳ�aJSi��&��L�zb�w�8��#wY�4��M��������M���4����,BJ�軫V�e]L a@��,L�tX:����,DE������3q͋]#b�Dl�y�tك�;r?��I��o�\���9Avdaz%��ja`/o���TOؙ��ҰXz*���#�_+�D�Va�}�-��ZğAy���R��Z�n��e�@�4Z����~�)eZD)�j���~Eэ�i{��I�N��K1�P�Z��f�f��gm�V����ú�����\�;�oqh�c������2-�$���W�sC���;u���C������X�}ù	ņ��P����B��Jsu���Je�Pю6���f̀���[�\˯\�٘���$z��t�h��Ռ����@�]	h�v���n�$&[��)vk|;b��[�8ɧ�I�P+qEhbV�@�l%�V72���_�I�?c�a�;�kP���Mw)C�<<��̋"���CeI��2�׸.�bk�;/V�5L8v.4U�nM��`��������n����xA�˦��E\��-��N��5܁����+N��k�$�Y�X�n��JcZ���d��P1�(S�$�Z֛��s<,I���5�71�G�z���Kc�R���o,Qܹ�f��6��w7wQ�sKZG9��ep�(S�|bY1�ex��y��V���������#/����-�a#r���D�����K\vqE�����9�(�+�9AͳԲ!��ދB�z�[̌qcFLǢ]ԡV4�,;�������'T1߸-�_kz0{O�M,�Y7+K9����Kp�3��\.��T|���Y{�.����ӛ�	�[��
V�޴��;t�d'��X��pn� RL%H�F3�$%��(p��R���`
�����O*Ĺ��u�����{��l�y〆%8Iڲj�f���]Y�DП!%8�$��c���^3��t`�df�%{Z0�f&�Iu��@�L�NŇkN��HC83����fvt��
�M��q�b�Zb���Z�R��e_�%x�+;����ǰNֳ˓��M\j�g�$�Iٻ�h�2-�Np�γƕ�j3��ػo:J�,:�:��`F�Wn\�,����(������V�*kpʗ�f�p+2������&����oc�.C���
��w��R��K?�	�t��Vn���_,���P�Vr=us�P`-|��S��׈��f�u�؎�(����Ԗ��k�.*;a��;����\t��{M�� \���'؝�{�*~	����:_�è���6��#H�]��n�Lx�y�(]��4IP���ݲPxZ'-}w9`���4����)���<���E۹�d���S4��\G��>Ÿ�|��
��MřVԠ�vWb�ň�T�~H���]Ђ)��u�
�r�h$�ܛ[/Ǳ��ַ���罸w3:ݘ[N$�3sNt�X�^��#v"��A'��>k��1M��i�3V�$
G���l����v���Vl��H7�����w)t�9�d�/po}��X���`��d7���9� ���/�J�y�k~vX�W,�/wR0V��>���ֺ�Һ�۸��Ը`'k��D:�NS2� ��P���wE���$]��tLh{39�b;�w!X��Q��Jl�Q�����K��:F��A���\�Ϛ����	�;E3N��˾z��iw �����S�u+����m���ں�V��i��y$��w�-��ݲ�;i�ҚVl�~�Q}9=��ޘ�W��vg�R&�W��^VoV��f��e��:����	�r屚m�zzo����[��ކ9�8c��+>����[Ֆ�2f`���Ck;",�O.�v��v�vL���e(�goW����q.=�7Lc*����B�eU��(])��6:�BT���\噅ރkNq���Y>3�R��i�<<��u��5=�V{�����=�;ɹ+Y�{�3�\�4go_P�E:��O.�e���p`{�ca�[W�;��͖��Hlv�2���LQf�w�	Sk/��JНx��t��Ys�v��q�[`f���G�G��X�mu����������/�x�f�����Yg��K���3!���Flx��� �}��l���SWc��Gr��0�}�.�)Gv*��l:�lr�\�ю���Tg%���w��q��Ã9ݥ�G���=���Z\D`�kSS��� �$K���>�H�r����r��	s�R��� Ud�ð]�������k�{(ܝ�s2���6�v�(o9�զ�`v� =�|���7��*R�ݭa��W��a�dJ�eޭ�k+�T������)��d�ԩ 0IB�b�[{��˨1t��y�0=�٬����]0�@�%���i��U��F�l������ܜ�\�Ǔ����^̘su_a��֢lxW�'����yO{t2]�8]�h�^��Vᇳ�h�P�.,�>��&#�0��a��3��*�����r]�[�*|�WW�w`�|[�#���Iđ��;A��e:����[Q=�:��e��ŀ[�(F]9���VZug�#�e`wL28Qy���������$zP�vT����y;v�]�+a�6�n�8�ú��z>�}}�q�%�ۢlY�F�#L���>�e�*��{��LB�W��m#w�.E�Eج��Z��������N�	儣�ʒcM#�Ly�x�_Vs��\�,#�"�F��-<�,(���H;��eBG�]�g�[��8���ئ�]1�d�A /$�J/�A�+a��6iXr�L̜s�X��*5��gXz�F��4s�6\}��t�j�t}�g0�^�KKm����RJ�(en��>�tA<�:����R��|d��J�|�5�;e������.�Rw���)!�����Bs�S�T�r����B�A��u��3�c���:���·2 V��׮ח'3���>v[�>����� ו�q��k���/.Ęw�/6+�ǐ���:�
2�5��ht<h��=�sb%y��̨)9n sk#3e��멷�Ϳ�;�u�[ǔ����1��Ւ�\Em*�{EX�����d�T�9�*7L|Pcf*���2�m���|�Z��Xٯ��$.3��О�T�Ξ� �];��E¯օ�â���N؀x2�f[�h�f����u�6л�|q(�i侳.|�/4�ӷ�YV�ەjj4��y�ϓ��5M��:�Bv���+��{��)�L����v�c=���rnn䱘�������/bG*[�Q!7�2P;V�Ү�m�n�g#�.���@�����\��6�7ڲ�B��E֛�h�1�M�'�m(,f�S�l7��I=G2�B�q��͞�&qO����/�m^}��{A��f�2N�
�V�R��R�ϜTEO�9�VX��M���cG0�V�ݚ헽�9��¢��v�A�$)��Ι���c�6Z����V�y�IF+�QL��e=X��T����v���y�n��*aޢ@2����ŏ�Jmw��%�4P|<9fz]�84q7�,����p�ܶ4�Q���T%[��Mgւ�֫�Xs~F�J�Ӻ��4{٘/�.��ɑg�Jc�oy��=^�U��)yD*�9�s��7b0T5�C8�0�+2�������F�b2��e��C3�oH��f����Ŵ��C�v,m]�TR��MK�kL xo����5����	t�#��Y]k*��1*���m�+!���ԓ���k�Z�1�,�/�\T0mu�خ=�I\h�
0�q6�/��s8N(�WW�	}y�:�֤��"�v�[�����F�e�֝�5��Gaxx��9�9V;�����n�9�p�Y�@�0v����y�U�n�gRT��g�&-�A�	���"J�!{W���W��#�a�׭�s&&�%�+������h���۫�x(�\���r�����轛�IbB�;]G���Z��ˌ��ɝWx���@�Ho���xC���3��fwi�ens��,u�V�zkmW8�g>Xf����u��Lt�a�z.h��\T�7/�
ݨ�&��q�I���\����� ��E�h=3NT��pg�@O���(���̈��賤y�/>�Wͣm�,3�i껱�d�>HQ��x��.�c�����R�w0����(0�Y��N�(�l`�Y�4�T,�(ųwvv� ���ʰy��9R%�����A�^����ӻOy�y��٧-]Sx�%��#���_&E���O�8�j,v֧J���	ge��jVf�/OP)�_qa �<����Gf+:w4�<�o�g��� ��F��a�����=�-	�Iv%y_-�n�Q�/t�#ީ��vR�<3��e\�ُ*AR<DV^)�=G�\��d���_)���fǺE�3f�cz�v�(���ըa�J��Z���囐{�/wj��YER�D#g1�v�Sj�'ZfNl�U%/��=�*q�����/8Ƀ��LWV����칅m�5A�I��<v���0��>@|��a�Ó�X`�l�g:�7�^��k(凑��k�8��1s7B_5���F��iN�k.�-�����w�,Z?MZ'k'ʖ�3-Vt��ȍ�;|Y�y#Դ�~>��|�Ѕk�r�������7<�ۥ�N��HoVy�������;Fx�u���`���2�|�)U��*W|��.�1��S��fx�%�(�����*+nc�3+T�#��*SFX��]�f���ӈ�J�hXԩ��H,9VtcS�ʂ������ž�(]�X�p$ݬ�|oo�~TC�ua��˨'Z���.���6��%����ׯ:I�S��Ҩ��r����C���V�5��!�"on.�WR)�-�{]|y?��������׉l��wQ�8fG�0^2�t�t������,����o�����5nz�xGA�|qn�G�G�1w�sͶ;�W%�U�m�'S'�������Xܾ���N��vh�!�J-�Oɱ"�'�;+NMEvq{������l�g�Cxn>�m�N!2��q�|DM�U���y���*
�i�;�}v�N��w��~�N9s��QCM������R̊]I������7Y�ն7*��B�6P�g �X98=��2�WRfsn�}�����baI?Y-ލn��s��]���N�+!c�z-K��5��Np��%�M@�Z�lwjF�7��\C���a�j\`���F�h�|���q��Ov��rw����	�{�,�V��5��ǩo�*�@��a_{6��(����^'�>T��nrI��%E�n���[�y^V�\�j]:%�v|��u̕o
�&��
�e��V^��B�U�1���Χ@S��<�u-�N�wn�RgdlÛә��3w"��;+]�Ǝ�mӑVg�
���/��n|���Y�-���4I���N2���Sjw
G:<��7w3oq�q�-W��_*F9U�݄���r�o��%�)1h�1f-�m
VԚp��>V�Ԓѧ`JI�_r�6���R�-��4��rAl1蒦c�1Ws��3 �<�K�͂=��eE���Դ�� ����W��_'_T;0�'9��/-P���?X�뛠��b/mM
+m�"�)�i5.�d��/{/%r�f�炨߽��{������n�X�hms��+6�sH�&���	(��yQ�Xl�wwBf��ܼط� �;ͧ��%����I�s�k�|L0ӕ�ŋZ'l{�\��m���cD�qY�me��/%$�F��B�r�{`��ӥ#L���e@����Wv$YڌB%�!|f��Eb	��;�r��t�V�����	�Oz:��ۆ�}HV�"��U��Ά��+��7���w�9@Y��c�:?o77Jf�Ӧ�X�3{!��J�;r�"�l{�Ҏ��RŘs�j�|zp"X�?"+:�����9$��� CY�B�}�%�+�P̋� ����%�8Gz������:����\F�Wd7��[��uH�B�0�v��BP)��Z��S�;$^E]m�d�|��8��R�a5�-t�''>8�GX;�d�Y{�'Ƕ�U+���t�S���޸�޸tk��JwnBq�P��U�Z�cy�ɧ��]�q;�L�@����<&��s�:��s^5+U�{�`���y+��$#���<)9�;�띡h�]N�ph.��ogA�����uv6���6Yl=�<�I4n�H�[�έu,8�v�c��"N�ݣ�ה`��gv�&�xK�Xj���~����ק��$5\�ri�ר�*�WR�4^è�i��f�ݹ�o)���Ԕ�K��<����=aع!œ���$���-��V�7��O^��C4T� �ֱ�ԇ�ʽT[t�'�y.�P����0@]�0塳C�^(�Hm��hھn33�<-�=ه��W`G�v�+8���yw�]�ۄ�.���
ʻ����ͣ����a���a�9T�{|GG��`_#�L��I�� l���n��/�ݰ$z`x�'kc<e�����[Vb��*7uѥ��1�,�����^���;k�������Gu��7���	ŅV%S��I@e�u6o�\ٺZ��m�}3S1!�G��`�6.\N�]��7A���u�Z��2����O���l��o,�t�<aE �̅�aӸ���|9(]d�ˍ�}ۄ��<j����*(���w�E�gT7��@�n��]����d`�J�]��N�i#��͒��}��FM�Wf��oZ�LL��P�ݬ)�|�(c�c��:�]Y0]�\�[X�شz��EIr��H��[�t)D�|�Eև���k�QĀ@��"NR����a߶],T����+��+��j�4�*����B��^ӲS�}w׾'�0��������ǚ��.��㰈��&	���괻�(���� ��2���kvzNn3�C\;2�REH�9>��%���U/E�
�Kv����v��o$��(�雕���e��N�����6鬅�Y:�+�cK9GW�q�3����M͗�l�o8��ԁ'F.�f��o��{�u��[ԉ�/^>]3�%�d�P�]MJӫd��J�J7��ut���(����Z���̩������:�C�$U�}��ۡ���lDpβ����Y(��:m^؝a;fޚ:U�����[�c�Vr�u3PO�ȍ�;F�KyE�P����Y�rT�>w��%h�ˣ�-ʕ���F��DɲeH/yk�Q�&�rn�)�����������ۜ�N���T�և6�p��F��l�װ]K�g�����%��Ʋ�ݬͽ�}u5*r����آ3���{ tˎKm'�(7�B���;A�k\�P��uu��IS
�� ,��[J��ޓZ�#{
�X�ʂ���@���1_��`�N-��iSPR:�֗��ur\��f���Ϻ��Y���i�w�{m#R�9w.)q�Z�-�N5���,�H�Ԫ�qxinHG|�l���Qb���s���Df�ОQ]rfV:˔�l�6ּj�M���jU��M����J�Y���R;��	�P�W�dݺ�h��P=���-B�1Z�R}�wF�z�}�b�o�ן�ޅ%]m��J���Vju`������{,���b��CM"LXy�x�7$C��8���i�+�����ٯ>F�;�s��S�8,t�j[{vk-l��U�ƚ��(�f˼�Oc���v����
P�H�Y,���$1H��������SJ��fw�0�Y�9�n��otZ�8_f3v�~�ɓ��:tt}�A�š��[*���&Զ��6�`���" �*��㇦j�y�G�8�0�x�"GO0{�އ�qu�[�).J�d����H��2N�:N�鸐R	�\�}�!1�I6u�I%I$�!�I6CIjR�G�$Uw-J3��� �u���~��@�BC�H@�h���xZ?��/���+���\�(;d�B�r�x�������	�
��J�8�����o�����2����ao^1k;̼�/:=գ��!(+��cΔ��`y��L2�@a��o�k�a�71@�[U��a�qn�M�sd�L�- ��fi�|	K�ix3 [{)%ꘙ���йs6�@��zt���_v�Gf��
Fę/s+�,D����e��՚PX&b���z{z]W*Ӏ�ƍ��&�"���ڶ��S��۷g���9؁�^ŏcD5�W�_^��]���+s\!��z̇��*��V�ڐ����_;�L�����.�� R�]O�v�G��M2Rk��Y�%�R�e�in&k5j�[e "���]��c=�ޣ����JT�-��i��#F������X:*��i���Y\iT�mb%�EL��eJ:E�:L���Gf\w�%�":Ļ�;M�Lҷj)t�����2��
ܝ	t+-nu�R�y��tj7:Fa��}�v��_sṱ	���u��ץ(�ދޘ���]H�T�u�<�t�iq��R�����c6�m�>�����T�8*���#��S2�׽��꽵�lEv��1�g��y��X���!���_mhBu4e�%k��r
oaԅ�͉䏭���3�ދu8��p2q�k[nD�<���e�T�8ޙ]
��d7t�gtx�iG{�wt����Y��&��EAΘǙ��N�7��]�נ]N�H��0Y��]��c�w��r�94-2��;GZ�:��q[3lu�ޡl�!S�;�P���^%HQT(}��d�E_JW��Q���Z ���κ��9:ƚ��B2�` 'fլ���Y�.jOA�l��F�V1���us����W����h9h=��!��љ�y�l�(�^.��W >С^O�u,4�/�h3��^N��n�bs�"2�u���D��O
/�xܻ� ��9��غ�it��%�͠�r�YV�X������N� V|%�(f�J|�i�甭��+ �.�b4�@]0Ui=A����e�p�|X(�k�t�l�GƬ7�&�?A�r]�Ѿ����R!ϴ����ܙ/�ZWى�ý��Bs�L"�[}��0˽�bf�����6�Fq��-�g�z�.qz�H��M5��SC���n{ɴ3/���.�f%�.�@��r�q]��1ϖ�2�lΠIqǗ,��ѫjk9���3���q��l���x��ef̈́�α]0-\*-�yM�����vFwS���]Һ1�H&�*�.<���N|Z�Q7���W���{�H|m��t�呐�T��]�EB3��(1Հ(N]��R%j���.��}űUӿ=������O
5P��[9�D+���wԪ<ȸ����g�f\E^�,�Ǘ+���S��δ���B�,Gf��!�o1��.'p�(�6�^t5�E 15��б���nΪ|�x�$�ѽ���o��dd�zC�ZU`Ǌ�����wF�h�~ڣe,ӻf�ӢMv�tpk2��^��H�-9���Yc�'��.]��_F\�8�.����Nf�����ڃ�Le���84�
DL#5������c��{R��V��]�f���Y��#5p!rt���f�N�R	f�"��n���Y�b�2��n�Qb��.�TՕ�$�V^��]�u����s2z�n�4D��4�<s�a�db���0V0FV­�����n�K2����V�)�[�d�.�y�\*��p��`�r`j�#����6u]>U|��-AXF�讙 B�q��-������'kk�S̚Iͩ���u���/��a�.�Qz�C5��Xs�'!usnu^�ӱ�E4fF���t3˸�v.�2����l�3�u��W=�R/r�Z�|I�p�U�|k�Vj�T�w�dV-Ⓩ��Z;�ٗv6"2b�ڵٱ�Z+��PL��M�n���(�8�i*�b�_���Y�%��A�dW�ӎS�k)����e.����{��<[鳴9ۇk��K�xF�o����nx�P�Ls\o��fZ�� l��˖.�t;3�XI{���٫�a�N^݁Z��MW��yc��J�tb�aN:�~?Eْ��a��K�޻�]i���.i$����3,�$��JyU1"��s^񙣂�;��>gݗYƉ}�oR������w�۴�jx�?`��ۮn��x�5� P6�[��.���WpA��\k�an�i<��1��i���YmYd�n9�i��R��pqc��^������Y�+TԈ4��Ж���~~��<���ص���F���Զi����]J���L����Y�j��'e�%���Ь�p]�� �V,;�d1l	}}���vW�"����w����Y������΁��]��LV\թ�ž����/k���^lW���ۙ�(�w�A�Ŗ��l"=�dON{�a;	!:�ނ��2q�F+�9���g���
�y��*�(�U�����ē�5�췑��P��4(�M�Y���r��#[m��+��ǥcYȱ,�Z����~�.lc����E�ၪ������+V|Ĳ��)�X�Q��%��:rAE:��^��)�0�ۛ�R�k���ȫyHP�+<Q�ކu{�ҵ�����8�֑{n�f�񌲸��t���-Z�J��6�<�ٜ�P�_�N&�[�{��Ҹ��_M�;��jQZ��)p8��)j+���y�*���rf��CBN����;Ր�¦<y�k��Y㡽�&�,T�b�;zvq�:�U�"iSw�u�:3E��mPT��)k���ǵ�r
�Y{��6�7J�.R�����6κ�M�Ј�oai��\��N���گF;��J�(�v=n�4Q�4q�l�����/����!��᪵f�`͢��3�+ܮ���j&,�K�NBp8&i��A%��(a�z������e����%u�+����&6�2u���i�j9}��f݁s5���"���\��_X)K8>2ʓf�5����B��^!-le�Ȣ�;O����C���.�8�o����|ʧ�F��-�o��J��g�����Ta)k$b
!�S抹j���P!)�{��2���cX�3��|�x�jJŴ�K�1sbu'IX�l��V	�STZEoˈ[�}�5{t�������D8ZJ�MU�RT�nՃ�g	Y(���>a���"|���//$�;���v{2�.�n������S�"��B��o�]X~���y��;���VQ���b�	g�d��ǘ��'{��fj����g#|#f<C/U�F>�MR�އ:���}}�ZЀÓ���'+�Fc���s�w��:��N2j��y�E'yxs���n3qt�.�Da��(�iPɹ�яe2V�N��ж�
�WaKܙ����sQIs3`S���E��ǣi�fim�s�H�^��8�V9�4�n��^�h�C%CK���y�����7���a|�B9S�t����6�+��	���S%��e�r�0�!_nȹ�C A$�᦬Աz/hX�	
y·�j{��i��8��c$�}$a��E}�E{k�qQVz��}�i�pM�Z��8�޸�L��37<<�p�7�H���K�]��'�����:z���O2��b.���;�q]�����鏴�y �s)0SX��Ⱦ��^6o��vNg00ӪB��g�K��U�f�ݓ��]�o��.����g�$���l|I�ޘ
G�x��(G��5���68�k{i�HݧX�]\l�Wqx �R����JS�z��R��c�|�N=�
�Gf�8�-���؏�$��x���
'd��>Xߐ[n
߸)2-�i�1Z۰��6��1�@����Y	x���u4��S�-��r�r�b�<Ъ��u��<}���`��*2J��[{l`=6b��L�#h�g_�q���|	��ɖ2�(��T��Y��/K=��m�� B3��Ҷ3o��m}�&q�d���]��a�[|�!�\{,MxФ:��wl��u/3����;�n���MU�=θ&e��=`��Zr��*�(7Y�-]����K��<.��]7���8��z�̾�`�U���������Ϯ=ᘖ͕�	թY���X�Tʀ�,�����[WXN�$.���X1☀V>2gTe侰��������7�EW}�v���b�1-�e��yj=["��RH�ַn�|��L�^��gLp����M�l��w��O�Ǐu�}^-��FwV��;i��Շ�[b��N�}�E�Tc�Q�an����n��{����a.�;��4�g6���9uۮ�3�S!�+�AW}��y�Q��;AW�ce�,{���`0w<�3Zu������i<u�����u�ў��;��K_-s6�Yw,G�c��ӡ�'.���_6p
SBR�8�<ML{}���0��-��⢚���M�&PF��v��s׃����Ѥ�/ݽ�Ǎ�:��ym���s��-��P�ܦ��4��˂�#hng�$�wګk�����������@��k_VmD�]�8py�-��ڽ/��0]j�`d�X�L���'1�����,�%�g2pe�����Q�⪃�u��h*�@.�)�H�v���\�h�'\O{�G����6eē�C��G�ݱ���7LE�J[�n�k���P=mҔ�Tɉ.���HfV���9+V�ᑲ�s9���QSA��l��,�8\��7+�1gۊUi����.����(d�l�>qz<�aZ;=�����l@�L�1k�>G��SK-Cy�;۞�e�a1`D7�/�qL�3˖l|�����H�ܻr�ڽ�_M)X�w{
vg��0�D��fcX3�zs�%�hN-��NiHmT*�bXWx�]l��Ar�=W}}��)z^����읜�A�.��O(k9��]��9�wI�M��f)�E5�n��e��+��ʷf���goT6����̂��"�Sx�����ْ�(,��9Y�8~{���dlX�n��;��Ց�P�������B8M�ҳ(Nk�vTKs[���Dp���X븓j�`�4�8i8���v=׬']/�E��E�S��F�;����A�49)Z;[Z�}���SwN�cS�ݼ��nE4�-'x��c�&��7�/���Պ_- �߆8DD�v��K�%�j�c�j����q�FY��t�
��|aD)�޺N�!p�����\�\���5'Q*^�l�e.֥[x&#�f��s��^��7I�b���f�=*�p�*%�OS6泹@V+�R�kZ�[��d���+��V��_/%6`縞�XEkL�=���<��hޖ_׽�0����O����R����6n�9r�W��Zh��X\ N�Rl$YL�ӷV��6���3aZ~��#�t��b�fM��#��]��_!&���!U̻ͥ"hf����ǚRR�A����*����Z�3��Ժ�'�`�h&O���}0�m�yRk�6�y<U9/f�xٵ[ʪ�zv��9+v�4��?�3F�fL�A�u���@m�C�f�|@���Ε�3&�_<� ��{C���s1hSK'.c�����4]���RU�庋8����f�\Gw%���=�����<mx�˒μ"�L8�m�yy�
�>�����tTS�����\iAa�HE�vQ��ٙWi��b��" �ǯp�M�-r�WL}7˂�Xpl��ھ���S�s��;�6]8ͽ��Yv��÷4|��"i>k��{7�v��=�P�x�KY�.XH��$���[I���I�xa9P�7����lMJfI�\���S���	�x[:;$��;��A�d��]S|�K�w	3N4z�������g(�*���Mb�c/����M�u�ul����N�#���_0�or�=)�{�N0��7YW��Z�F���`�Xv���tS����s5�޳��Z��H��U���8h�\���r��>1����� F��=�C����S1p&'� :�����(e����_3�U�/�^�lʍ���YxrŞO]$�xWܒ��I��:�	���>�~Iբe�6t����t�t�	�CD���P��!y��R�$�$��	�����U�
v�rF���7�Ƞ��jf�W����B�f1��o9Q�F�'����4hq�s�W��~��M9�`���˖q���]�yI�����&�Y�Ri�96���� v�I񋳓b� �-��1̩;L�V0�����G�P�F]Q�h�XzN�H%ٻ̢�|o�0�ȅ����i.f��E���@ӊ#z�Z�F��Jޕ}�޻$�I���1����m��A��(�O�JY��7��{8�ݕi5!N���we�+�C+�*�=Vk��<;���3z����R8 ��b�XR��ŏ;�J�x�<�M�9��h+�^��
h�3����W�+p��Xח�Ow��]NK����ˊ���8�R%�.-�> F9V��Tf�ϼ�4�Yt?�w��԰���廝H��h�od�Lʶ�c���'4r������s�����nճ��u��D�y�W7�����{y��k��3)�o�q�i@��)f�;!wM#�`LS<��`c^/(�7YR�[�L��%���3nl! �No3���ĝ\}��Zz�"�Y9{���)�M���y��wg	�V�=9e�A����Tf��tۃ�t&�M5�}��j\�$�PV}�p�c���$o��u������>���}�|2�y��v��m����s�x��iI�7NǗ0E�WV��/�l�x��o6;c�\:w1��)�[�g�Ưͦ��;ՒMa����,U�K��Ϣ�	�[i4��;��ޖwHH�]�9֮�]$\,P���XM��\o�qG����
>�'D/I����R>���w�;��P��;D��P���r��̞�*'d�1\���J�#+����i���E��9�1��o.�\�B�~Xx9����thjU�xܷi�jML��-�:�S9m�6�㽉eO:��n�|N<�>��vg;��O��#F[��G�6;�1�!����&����ZWfo�1m��⎥��Z�p˽ŌV;��*����T��b�4�f�p��0&m�hG¯�o�6�Ʉ�7R`��AD7�����:��Y�t8��m!W�$?�O@U�1nYy�h�J��s��l-kt-s;�o�ih�|���ɾ�o+$^�:~0t��鐕�Qg�zgM���z�T;��..�(N].]/��=i��^��O�7A;�qf�'=p�S���(ya��Rƞh������������i�y���"�ڳЇ[WόFqCe�|��l�j�8�b�t�Wr�9*賬K�RN gfL�Մ5m�Oy*�d�k:�4�7�����E�I��/�oݝ)��/�ʖ�t��! ��Qb���*#Z�qL ��QUG�SEb-��T�PUZ�\`�aiaZ��J(֕3l\�e��ҭ��[Q�PAU��AҢ(�Z�[)U,���e�
5�J�Ъ5�+PmQ�EV�����UR�����l�Wb���%U�Ҷ�mFTb�TFR�m��U��ֳ-����8ak*e&1j���DD��Z%h�L�8�(�T1nA�[XUŶ�Q�US�1CF��Æb�6��1p�"¡�j\YD��nq0�2֦���E͖"�1��1D2�p�5-*ᒎ)X�Tm
*�%L&�ҫ���ЬG3�(.Z(�,���,�8�T-��l��)��FжŊ�W�O�A���(���j�{vά�����P�r�'ݽ�f�c=�C%���\z����k�k���&�戥��NU;����fj¶)���qs�Y��H?�L�qN��s���<Ed2�W\`D]��:�sɘ��;s.<7���Gl7\�Z�R7��s �ᢍ���c+��|�s��04��dF��R�^7����p�}r�;"ccƌ��I�ݐ@q|��6�l�ʃx�VL�F'�:�ZA�J����u�w�%
l���l�@W��§ٹ����ɞ�(#��ڸ	wR�Pj܋P�
�0[����c0:4ڡ�#W�_�e��k��y�|qR�\2��K;��	c�|�ʇ�j���~j3m�Æ)�U��O�����C��0��η1׵��H"^g}��zf��y�E�������[����.���r�/��q(�[��F�żOw!�>o7jz1j�3����M-�W��i������11Z�_�&/9W*Z;�����lz���{�A��&���K=J���<��VnL$ru�魚J0V\Y�^�Q���z����<���}�Od{�J�y��KY�ܮ;r�i����d�����X�v�弌Qӥ|�x��͛m�����ˬ��cjZ��C��q�NV�(i�c�$*��e�m��l���:�I�h�֦,�B�:�Z�9���^��8������^hՒI��v��l�	}	y�yGU��Ġ��uq;N6.�v�ǻϣ���ȗo]�[�1C���.��Ԩ?K���{'?��2��}��iNz,�"�xc���qI�n9q�q�q��m�9-]�
]���GNV�t����̒1[�]��1:��W�Z�K޾��B��ZV�c�
h��=3��uz��>:bQ�ob��F)6L���Q���|�]��O8��ZC��>�>��XU�*1<�,�T�$�v$]�g���V�G2W=�w�������,���+�C��F�{�đ�޴�i::��Q�����Ì6��D��B ;�����4���)�t�d%o�V3�Q�@�wc��f��&3���pX.^~;�8��%C�&�Dj�4�{m�~.U�0�����������;�h�R���
�9Ӌ|6.����o������jɜ����hF����U���ʝst^7�����';�l	�3r��}]�,�|�s��^�S�n��tjҨc�P0��]m�9�eȕՉ�o6��]�훍P&4�����=;W`Ǭ� Lkӏ��olGs���R7�����\�L_�c�a��r���gu��u:�*����N3X��Zx�?�=)���wU� :���MAޫ����E�9r#�[���)y�ʧ\sd�9����L_����|��W'�41F^]�^�c�i��C/��Y�l�|�d�=�{F���K���H��g�sw���A��-WҞ|��!��b�jmN7[ʩk��t���u�^jc&NaH����J�+C�ֱ:���Ԩ��{�4�P[Y��4�n��~ڥ��F�ľ4JK׸���9j���Xb��q����u>wW����5�:�������{�E櫊[��]�w��P� ��v���،��E�kO�W���g<	�2gBݎ8Aj.�W��6�A�s�ƨ���b{(�Uݕ��o	�Y�����Ew�׆�d�|f��m{|:�E\�����7O��)Y��ū��#3���n�.6v�5��mn��e��M�
�+K��ȩf��������]�벥7t��(G��Z�'���v�'Fd�4b��|�B�dE�8o��`�s�l*���gwF��w��':��as��:�r�\dSzGd6@�_1���Q�Y��f�V{��7n�N@L���Q�bj���k
.�9&����^�	�/��g-6Ʀ�TU�K(�m���+&j#��*.! �-��ٷݢAB������u>&�#��
�Mf�=�E�+9�~)��(���%�@��ø��&N�ilrS$���um`�GAۅ#�F񭃙jc�F�8@V�v��6�v��FưaHNK��fo4o���XQ��-<q�.�I�6w1Q9Y[5���J��1������si}�5q告�x�f���I����Rv�u�Բ��?����lƦ��4�r���5���\�n�$�Oi���T5�����p"�щ��,�c9�[)����^�Vq+����W�0����R�������^�do[HXy(��j�=Cڂ��t�JC��&DW 4��I����ż���7Xc��!�6Cz ���*F��ʒ�m�X��!z�VJ��x�'8�OJ�f���N%+
��7�ut���m���3:T/��ި���M�WF�l�u} w<����v^J�kq-��s�]��OFq��^���s�ѩ_�KM]u��Py�1�U�g9���n2��$�b]�E�@Z��f�k��˰����� K�ǰ��>����}R.I3�oU6wj�K�j��0�"c\g^2"�aE���L#}+��ڶ��Ǝ��~ܞ�q�Z��<d]��<�{x�atc"*S��Y���tvE�Ǥ���I�;պ5S��T$��2��{�ƌ�uF/$@\��VK9T���9�V,`q�yF�*
�|3�xR�sN5��-d��{ZV��{�Eű�4�a���w򘾫y/�v�a9=��P2褷�\�C�}�q�*!�j��tq��O�U��Wo�/m/;���Z���-��f�T�հ�DkC)�um`�z�q��z�N�Ԛ�=J2f�Y���"
����3ԉ��C[�����?�Po^�{u��Sw���.��T��b�ƦV%���=&�qa��f���E=��Sn�ϟ�$��R�`\�4�*��y˃f�:5\��gq���r�I�׎ܲ���-�8m�}�N�9���� ��.ǡ�v���5�Fm�q���^���������r߫f)}�Z��nFbߢ�n$.c��o���p�6hv��
:^�O����}&�T^[��8�^r��tn56-�{��Gwss;]y&�75O{|ax�p�u����4b������\�^�y
�Ʌ.T��[�E.5;�v�b�-��L=���'�m�}�gp�=�nU����rX�n3�ю+2�s2�p�[y���)�8|�;�ꖚ1�k���H��Je��B��M��u�_J�8�����˸S}}Pw9W|��-]�c����^fpwO)�`��J�/5\R{��]�tF2!�p�%��۵9�'���<�c^Ҹ����&#�ձKS�{��n��R�F�����1w��?^��Y��F�,�ya��(�7����Yw�R�sn�w7w-�s��P�U�Zi����-4��Iێ��g�e��z���_vBHt��t=�)�L��{�~\tC��w'v_u�/�L_3��YM��ٽ��i�.�K=[Z�)FT�&�QZ[S���'n���.����	�k����puƸ�dEE�8_��eR��aTE�ʌO4ĳ��jI�击/
z��j��\�Fz���`W�1��T�*Qȃy���Egc^�Q�7J�޾v�.M8��WڋH<��6��]�!���{��)��i�=��ų��l�oU��Om�-��bs�E���PٶE5J*�˺�)-�a�Nb+f�{�5TJU�o89�e�����-��Ǡ�C+���M��WP�+�y�6A\\9p�5y}p^Z�/u������r�۵}S=,&s��:I��󊫇��V�f�3sb���Q~8�_���tsꁻ��4.�����-���mW��w����B��q��1Nk�E�n&jMz��-G���<�d��qn��iiƟn2�O�Y�l�����RR�F(rz���V]���N�����[|�eN}�2^����
ʵ6�q��"�j���쨖��N^�U��:yGv�s�n�te���C���<I�@�����9ܫ����k���v�AHY� �Yy)�A�R��P���Oe���鉍����Ρn{Rb+72F�Z�����;7��J���QI�'��ou����d�}6U�Z�+�_=�o�U�W��Ziֵv],�u�e����5
o�q����͊5�p�J���#�9rP�2�ؗoyw.�ͱ�^�r����G^E�u�K�~�ƺ"�V���Q3��wkf��Ki�H�q��ȴ�E��ZfT_W�,.:��]Y7��s^r۞�t�y���h�'�����=b��xpiN˪51S���2��RSYRm,�<]���k	����=�Qq-�K�����8]S즍̎5~K�Z�i��>^W�ź��U��vg*@���K���_s��f��4"1��K(�;���Y3X��o	�~ha�{��\&(V���G	�� �q�Mf��z��XS��P'9����)&���H��-��9��������;~R8�oәj0��Q7'$�b�4�:P'����"�բ��ּ����k~룈���N�^(79O���¾�MY�m��x#���'Eg>�M񎒌�u��mu�����6�[؍��MO�Eq�����]���Z�WS��!뛕�%�}�KrN�xzf�����N��4�yl���=37�|����f���gm�j��GU+>	�᏷�N.�;8��!�7��X^f�>毱�ٮ����̾�]��.MiW���ױpq(��Qʍ�oLcO�!��<�o����9[X�EFj���[J�JfKٛ��Ԣ�&.3�{�+��xa������9�y'�9�����C'�l�:�ʩi����䅔�j��]��S������m!i���z��˿)�i�c���~�ɵ}�F�v���ŋA\c�#�k�.*�����Ƹ���u��n����{��F����{����W��ʸ�q�:��t����3�؆��C���q�9h��8GYʹ��Ky3u�ᰑ�-�j����=�a��xȊ�EO��X/y.�}�)������_Q{��죶�Z�����:;��b��1��#��r�VlU��޷+��`v_P�ӺT�E��%G�ƫA�eC�v8�?k�-5�[��H1��sK�ٰ�� �ז)���Fή9��x�|Xݓ�CI��[8���!ot=j$��7|o]�*fV��Ԏ��wp��W1�������`V!��WvQ�xXU��b�f%��GyͿM��t����'R�
�آ�v�;�r�&�m�9�x��+&q=��++g�9�9]��2+��7"�PٶB ;������nz���+9�E�P��wg_D����7�- �_�M��k3�n8}H���8W�I��w|���!u�s.��&#1,zCC+�N��X2����K��
;��gr�QU@ZN+Mz���{jc�pkq ����W�=Lz��f�kIG�j��.����uÓ�2�Qe�;���{Sb��{�͍T���z�.ă��67-��}}5�#zԜ�4bkZ����r�*�sgK�Br�A��^�'�r��{�v�{�Yˆ˝/c��6+S�\-�BDNy������v\A|��[�p�t6�UZ�6�p[7��I��W���X7H8�IL��ˡ��w�u<�W���)����xZ�eO����*��a8	��!GʵT����Y�8-$1�s/�E�[u4R��D{/��K;oS<�jnYn�����������N�r��.(��`}�.��`B���ci�5�ثN�#���Y^������}�	��X $0�q������T��[�%�f�,'��U�!��&w\��Sy]=8��޷�9��;R;h5S㋭�T�؟[�	n�sMl�t�q�,{X�R���C#?h��]q�C�iV��{&��w,na+��s%�#���g)�8zz/L/hXk{�����5����Y_9�-5-X�58��*Mh�v䵗��P:��j����f�`���g�դ*C�w	wxĘ��&E�d��vh�"{5��Y�������X��(���dۘ`I�d��[0����^��\V�>]/�<�$���$�L m�����`��٤����=�8R�v��{���s��LԐ��vP;��.䧓�y�b����V��i��2���ܣL)�`=K��
�����GG7kB4�(���e�&g'9�TaOȺ>YYD���K���1���/��oo��װ��jȻ/c�֫bǇy��8��v^r�"c�3[���>���(�{Q��Ք;���AK�Σfԓq�Y�n�Z��`U�[�l�I�]��74,b�9�I�d>Q*A�K�7Քvk� #��ap�'t8i�C�28��+���ijL�.U����_+��.�y���e&j���x!b��o�2S�E�(�t����(,m��cr��5ʙ�n�(���,Q�Y�i�U���s����$aϑy����!Q�2eN܄�.͵��#�D,gev�يO��Z��V��c;��;b����_1��ϯF�*I0{�����]\#��,L��Nzgkh��fI�q�}���!�7R��*��}"�r���$�~A}m�|���5� ���;�fYW�EQ�J��g5��S�����ا�v��6�LPa]>�|��{%����w;�Ws(�ڻ�v�rמ^��u�y�e���v��zԛKĎ�GXsڱ��H�H.���w��$ �&�8��O5Dg�ެq���!�s�v�ё۴�E�̚��T�73.�F��k��t30�yηݙ�ic���f���}co�>���
�%s;Yf�9Yy-��,9hF���R�'� �%S�pzr3�݀�l<�]="�r&(�"��ȱ3Vx�F^�.����#�0�!�r<w���Dn{�#�s!
�"�8�~�]ԳK����9tI�uv��Ft0l��u�*ϲS�\͒9{]{|���q�p�ъ�z�s�����Ս5N�t��Ix��U�4�pə_@�Qv�ؖ�{4x���`��`JM^���}�;�+�r������}�����m��6+*VJ-�B֫�08K����Ub
�eA�JԬP[iQA���+X�Z�eb��Z��m�AB�V8�Fa��D�b��X��%TK`�-`6�D"�����i
�+UY+eU�0a�(UT���Yl��(-k1LbQ��+��YYKB�Kk�Щ
�±QQe�	\[RԵ��Dkd���U0R����X�j�QPPU�m`�(��
�Q������A�aL[�[j6ԩDU(ֈVL5ŭ�X-J�)R��¥FՂ�
ŌUH��a�R(�°R�Z���+YkB�J�Kh�
�m�caE"$�R�)P��V�������}�0���un���0�G9�Ղ��"m�/��̜	�M�˻u��q�N�,�f��@5%=nY�;#��̸�9\��Wr"��"�xݼ[���13V��%��e�ž��=�`�9�n[+�%�&��tic<_<1�U櫤����\c\g\c"9J��j�[�{�����a��=�c�f�VDK�av���j�Z�{�U�U���H�[�*z����MS�=�W��і�=�N���q�{��+΢�ݖ�%���dEz�&W�R��aW��bgb�5
��J�|�o5��Ji�/�[������;�|��}�(��!��c�hj��݌��_�r^��j/��p�ۉwl�@v:8ߥ�ۥ�bٚ/dƟ�syw-�s�SߊSTwyK��ޭ�,�Sf�+��DoMM[�\���iyA��y봎�)�ި[��,zC��Fcy@p4��%΍�uO�pb!�ۈR8��#y]��9��5��Le}��LX�u竷dăA�]�c����G��e�k=�p��3�ڕg�&�!�4v��}(�8
�*:����^7�����9)���b�������`m�7�dSÕ���*I�z�rW4b+!��(�MZ�Ъ�ْc��7�c� ^M��m�=�M��Ǫ��6jڌۇ#7e^E娳�E�k�Mv>�n�<�'շx�����sk�^��q��W]o:�/4�x���|��pbr�v%b�;l<M�������gj���/�<����W�D�ũkJ{�ʶc��vŖظ���V�t��1��v�:��)#T0ɡXt���tɉ�~ʥ��uE�$4�\�_�V��kW�n{eu��=��Z����flʃ��o��Z}F���QMa�J������[��%��8�T�2�v�Q�xʿ9aE�KL�����.d�WI��VVc�}u�<��ϋ��.���tr�Ց���J���׏����������3p%������\Y%�:��wKQ�O�����+{��ftB����������}K*bƾљ�t+΀�-V�[��:��*���${�D�yh���EU��lY�m�k���pl_�>�۔)�5��C_v3�U���`���Wr*ύ;ۛD�L#%��>�eq��:�k2ڊdC��:�.��^K�kc�J�Z��^Me'u��=q���*�(���Bw7��Cu EM�hN�^�ǯ.�3T'U��N(ά�Jj�}��`��X��}��h3�-$��P�%|Bd�`x��5=�u!�t4���}�T2��,��0�zɩ�k&�'c>iׁt}����=�}7d��=#��zG�Ơ\�q�:L2`m>�>$�Cl<a^�=��C�0�!�(d:�L���l�AHk��*d�5��{髆����ޏ�Sf���H�`���˂=�u&���K�$���H�|�D�pN�q'���C��P���4n��<M!4n�!�0�!��8��T�I����Y�����j2��pG��@��{DOY=JÝ�+�{�w�I&Y4w�fK�uܿ`�M��5�b��M�&��06��S���4n��<f�q1�E�KW�u�6���+����B"���`��{�OR|��h9�Ou�Ԭ;���2w�c�I�O�{�d�RL���Rx����1
����l�!Ćٟ�񬂤Ri��ld���1�#�d�B��Au7I6�Xu:�d�f�|��N2�瘞$�'��<����k��~a=`o�y�|�$�js�H����c_w�.�ϻ�}���p�t6���	�������L�Ad��!�N�u���fS��I�h���d�~w:���O'w�<@�'������毵�EO�_������W��"=�#:}�"2���bm!�=f4��o>�:����':�4ya>a��S����5�0q��XM��:���Oq�[�y��YQ:P�-��:�:?}�U1SO}��	�G{�é�'�l︑C�i'����,��z�a��y��N��5�|���J�d8��ϩ��O1���?nS\�}�Jٟ��{L��=�
�<}d�{�:�����u!˜C��&����!�4��l�q�I�=M��I�I�Xq'̬��'Y��{ﾵ��{y&�gn���f���f�36��o�k����@��8k᠝��D׏�MV���G�1�I���5�V�{Ƒ�P�į0�BH�hzj�v�L�J�hw�n�A�e�J�E{�me�1f-*�Z}l���:��<�b�fE}�m�ٺ�A1��$}���B�a��_XN2js�:��&����������R!�5;��'Y1��C�Aa��8�=Jԓ�6<�s�X���u��W���%ټ�s��<s���̛͐�O:��Hq�gT����&�y��=~Be7���q6ɳ���C�>f�;��PP��pu
���`��'�u��u��f�߻��{�qs;$����ROS�wvCV�>I����P�6��q�S�'P�N�� z���M��d�y���׽" �9�f^��qf��%$9pg��0��T��� |����O�6̡�Y'�Շ��yd5l�Rm���`q��=�gP�@��0zÉ��X�s�",G��5_dչ[�)������Nz$�>�d�RL��8�����Y�$�O�<r�̈́���t:��35C���`x�oX{1@�CG虋b">�s�h�Aqu��N��{2�C�M������C�MLwY�I�/5�*T��^���n���:��'����q���i��n�RW�ދ�cލ"��[��;�G�܎r=�}��� �!�2���=A`jw��C�� �G{�'�����i�u��7�*T��~ċ'۰4w8'Y>I��xfb<Ǣ8E��#G��z2N�ڜK��o�x]`�|�����C�0�!��8��*by�2u����+��N�*O2��i��&���2W�IݿbE���9�B�|�o����^q�;E�oU-��l\�����P�B��|=�	�Mn��<M!5��I��)�IS���'�;�6��<eC��*O;��I�sx%v�e9����\x��o���u5�ol}�AD}�^����3fi$6��<f��$ѻ��i��.甓�:�}��RM�'�`�'�4�ĝd��O;�@���O~ϟ�m_��ů]|F촅@ms�3�Gv��uYE�oc�s)�^d&�ٛm9��-Go`Zw!��m�z�Կ�����*ۭ;�wU��w�r���R䳫3goH��J̥2���\��D�ق��z��K�sKI���E�s-���4���%ٕ���N��3��I���2N8a2�9�H������l��z�f��Hx��<f�8�ɭ�<C��Au�	�N!���e��<y�|=�H��^��������4���X�>d����{��Ox��|�'�w��8a2�9�$Xz�04s�d<C�a6f��Y&!�pd�&�<aĝeM�=I����r�Y��������Y�zi4�zû�2|��n�2u��l�wx�����淒O;��:�!=Cs����L[4�|�OP�$��pd�V������־�<����w��{�\��*Oe�;7Bq'Xq8��q��c�:��l<�I��'{d��?��	Ć�cY3O�l�u�z�s�,��z����Yϔ˃ßg>����;�a���xɴ����N2s���q��2j�|I8�G���O_�M�8bRx�ɳ��!�&����\�8�2q�8��s�fUǞw�s����=��<d�:{�a=I�o6L�O���O��2n�>d�7��'gW�ԓ���������K�OY8{�Ad<C�g<�q�y}1�<��>��ߝ���|s�T'w�OP��A`���$�I8�I��,'�:��CE��O�=��Hq�4���q��<��gP�{���_7�i�q�~�|����/��^�����'~� ��C;�J��ɮb|�d�+&��IĞ�x)'m3���q�5a�N�2
u��M>�R`iy���w�=�ʤ%�<�.�r,z=�">�UD|=�&]�!��d�;���>C��$�P�k�:²|��S9�I�'���a8��fníI8��X|��2;�l��t����y����:cGN0<I�œ�Ch}��XN�g߰q3l�Ag��$:���1�d�4^�2T�&{�:²|��Fs�:��'���6��3����n�+S�$�DÃ|�F�#���3*2�.,\� ���G��ɴT�+p圃��k,��)^�z����
	�^�of�#�@/��«���8�Oq<�.���>kp�Z�؎�=-�˘/581M�Ug�jEnr�W�څ�Z��8G��FB�=�I�l0�0�N�!��M$�
CG9�T:��4w���Rh�u����7y��R��t_�E��h5��1�W�κ��|�;&Y6���4'<fM٧ē�57a�3�C^^$=a���Y8�W}���AHk�
�<JÜ�*M���w����9Ço���gd挜_fn�6A~�#����]{�G���!X$��l3Bq��ɫ4���M�x���!�w��S�0�^ӈ,��=��u�C_s��z���ɽ������b���4z$G�{�J�{�d�{�d��']�bE&�X�X$��nf��!��x�a>I��u�N ���!���Aa6���}���}O�����@���D�z>�Q==�R��l<d����RL�h�d��I2��1"����q��z��d4�j�3I8����'�u��:�{:/�u�}rj��t�\G����G�T�2�mw��|���<��N�z��Û�Y=d�{��I�~�	�)�<Ċ3��i!�S	�i����z�f~Ǖ���<TeC��{@�O��z�Ĭ�	�N!�}N3)&���'_O��8�ԟ>��ĝ`|��g5��x��{���'��=Ċ3L�y���p�|)��*�^�����=��A�a ����C�N�@�O�q��Y��'�:�O��I�Zq���M���Ԟ>����N�=I볚�Bq�����"pR����>��_D`��!���8�2|��pe$��fhm���jÌ�J���>a�N%f��2q�Y�l��>��O_�O��I��y� �{@��-��Fq��������{��'̆��d:�$��c8�>N�I8���46̤�:1a�O��3�d�'�<�d���O����|����v��d7id�i��g�#1e�>d<��D�;'T8ʲz��EԶ�@��=�f�������7ս$�_L�I�Ow�x�k��]L�C%9Y���]Cs���GS�	��OI�ڛ��3��ǌ���+|�P	�������g?��et�"<��~��q�2l=� �<a�k��!8�jw�B��
G��q�ģ$�&��T>fRO�F(u��iZ@�']��Blt�}�R9�r�G�,z>���IĘힰ��	�����6��lCi�7�bJ����|�d��N� �2z�d�I����q�}��\��>�s���o�>��N���t����6��X`q�~�>�:���1=C��.9`u��N�x$����d�(Mr�%d�+'�s�8��O}�8�;�����^����(���c�B>��GL�OY�P�%|d3�`q'��oaBu���`�3i:��3���jc��)'�4w��++	��k�ͅ�;����9���h���u����9L0��m<����N��:��!<<�!�uOhHx��4����!P�N �\�qY9���P�&T)��Z�^�B��G��yq��=�:��q�f5�u䞺M��q��gt4��q��z����C�0�!���ߩ�N �9�����u�ߔ8V��"4{�<��*����L��y4�8�r�y���:}dY>t���pN�q'���l�X�f�i�	Ě݇�x�Bh��C�a�C�o����	��Y�����f����#ޑ_Tq�����Oq�Ԭ6w�!Xxɞ���I2��o]�'_o�"�o�1�V�6����`m�����'fwb��uZwU���5z4Dp����>�x�Xz�AI*l�x�I�VCG9��N�z�����'���X��e��{�d�RL���I��S��+�>g���]���_�e����=#Ї�CP�$��!��Au�M���L�M�^��Ĝed4s�Ou��ԞO��>@�&��o?0��;��O�$�Os_A�߭��c��#�'OC�$����.N�^����q�~�����m�����ja��)�7���$F��2�l�C��u����1�~�W�%k�T�7M��0c�w����yw��o[��ݳ.�:S0�ܧėi�:I�W11ș�����.�'|��T?}�!���]�6��3	��'���i��,���x�Y:�ז�a��q2�6�ygY;��y�d�'ϩ;�"#D{@U�X[��E��[_b�No}	�|��N�Bz�}�(|�H}�bm!�=fp͆�RLg�Y8����|���J���|ì3>�)'kڨc��g��=�k~���6�_�ڕ���8{�$��'�}�I��=w�ky���o0�a	�︑C�i'����,��z�3a��>�q'YXn��d�T�n�q��5ߛ{{����<߼7��<4�|û��s�	�j�ԛ|d��q'X��nw[�N�5�k0�a	���!�4��^�2N!�{3a��$��Ň��膆����,����sB���M�i���|��2j�|a:��iԟ<a8��>�{�E!�>g������1��C�Aa���C��"D{�z0{s�S���?U#��������i�6ɽY�C��d�6yHq�fj�>��d�y��=~Be6w���M�l��"����u�*
�>=�" ��]?����<�7�'~sﳌ�I�N%&�i�5C��I�ыY9�!��8��M��ً���x��q�ٞ`���L��{���6�s�� �N!���y���s�{�{����9ǎ{%ABw����|ʓP�pq����a:��4��d�OXz��CAl�Rm���C�gP�@��0zÉ�&S�=nxl��{�}�s�w����e�M!�����,��5�w�*T�:�IR|�ɬ�q'̞9p�qi�k	�5C����`x�Ǭ*RC���|=�^/�%��\�&����G�DG���B �{�,���'P��S�b�u���%J�w�ԕ�����	�O�=t�6�&wCO�'kt:������o�����^ۦ��scHCWf���F~���0�2Y�%g�{�A~bk��3��r��[�w�3�F�W>��XZ�1d*�{�����HJ[�F&$��[�h�-�뼯z&J�z��k� �Y�6���;j+e84��t�R:%w#xo3�����G�9��]�����bL0�P6��u{�L�A`js��C�� �]�T�2g��M2N�y�IR��>�,����w8'Y>I��y��S�=^=�g{��{n|�g���;<���CP���3d�Ad�1��:���s�:��T4w�!Rxɞ�y4�e���$��'}�H��>��g��	�ٌ��׽=�骡�����~gsd:��d5O��5�0�4��i&ШxyN �J��x>d�T&��ĝI�*;��<d�ݗ�=�������z��o���zG�&S�s)<x���b���3a�C��f��4��&�u=C,�Av�m��{gX��f}�8�	�ͯh�|=��<�ۉ������?bP���/`x��'|�y�I��̓�&SS�ĊOX�i��S�4�&MS�i��,�7d��qה'�8".��=�`����쟊���2�:���;^�d�*�����2{�'���Y=I��̒z�����>p�e4s�H��>`r٦C�=f���$�}�u��,�ݓ�I�T{��7�����/ǛeI�E}}�]�?U|�}�����+G��Xvӌ�v�{���'Y>���Y:��O�ky$����a	���X|�`js�I>B��P�$�����>��h�������d�2m+�t�I�N���П$��S��'h��I��g�1�<}d��q'X����o0�Hk��C���7;�H�P�'ɞk_
��%pj����r���7S��z�F��.a�)'�uC�N�`d�'�8��(o����w�w
^��q�i���WE�F��3I�L�+��j�\��/V�W���%y�b��n9l�X�Q0/j�t�YFj���ܫ���Q�۵�l���ɛ����*g7۾�)^���5һl�eFw�^�a�x�\������)xl��j���Ɵnc&_!���q�Ɩ��*�{"r�
"���51v��B�,��AfI��is;Xr����{������M��m�7�g�Q~��W���q/��]��'y�u�0'��qG;��e�%w+�:�Q�u�ķ�K�����k��T^�����FUf.Z���oo���{t��݇q�X�i��]�}��	���1��ǻ|�eF��/s��ؖcy��"�ۗp��*1��esW6�g�B):��@�k�����^J�y�ԣ<�y�ۗv�D'NJ<;V�I\�q�焊G�jy��9^E/.wmp�Sz�����|��E�f3�ɮ�w����Y8ۡ�&<���7W=���o��阽1d쎚u����W��|�W����/B���#�J�����yjf3��s�LJh���
5Q��p�y�Cy��U��٫��5���H��V[�� �Zis���M���b���J�C	����ς�q�S�8�X.��Fe�A��g���x��s0i����@�m8�C�a������W3��ɇ��c^�����v���.�|Q
���?ZM�ڇ8��=��]��6��^�����'��@:�V�s�ծ�{9�`%�[�"H5�0�`�t�v�L��W������Z�!s"�.A����-�-ԹŐ4�uP����Jk1�\��n���0g��r;�2�S8tE���4j%FR�ŗ���pY��[�=xX�k�ٌ���:/���	,_f#Y�m�T�*ͽ��@��gW��"�o�偉�;+U6���{G���+V0:����RVU|2��|�9Br�S�����0>,b=�9�>bL�֥i�/���<#�4����/I�3\)eT$���4��]+�d��������us���[g�nӍ!��g*���k�Q1|9��:YX�8;�F.���9Y��Dv��KS�1@���L�Wk�Z֥$Je��gfR��B/ru+3T�Y���	����V$�\D����j����.=�9�j�q_]É��z�������.8=<6�f�Dm�
8��eބ���
����z�zl3^d�%��Э��D�b����F�5�&��*�׏šp�MR�/��@����^�6׎�$��fd3�]���y��0I���;��s�٘�Ty �}9��[J��~~w�s7	���$DY����)�6=�d�,cZ,�λ���I�l�a�٢�B�˃%w^�t09}s���I�.��T*a(�W�>���-�Ϻ "u�+��WD��<��v��Ut	�0;=�cKP���t��f.0��X/��!�~eST�rS�4�Q)��0��*]{N�
X��8���np�����JFi�q�#}jƞ�
;"�MH���������YUp��Tٙ�=b3ͳ���w�l�'u^A}��h���*p����or��m֞!J�-X�J�ƀ&�rRe:�R�g��`A���qOզ����rğ�zzs/L�c��Y�G��_'9�3���>|d�]��2XS�z��j�ά^p���w%�˄�p��\fy�Hf�c;�<Ϟ��5�ks/�:�>��X�t�a�"��M��+UbV-�	�'t2ɸ�R��h�iKO"���\�KJ�Q��#!�kϲ�2nT%�������Ȏ�I�zi�x^��� 9>�#�3�*���=x,K<`g�0��Sty�X�zY>�oVni��l��zsuì��x�F�B,���x����NA�Z��jD�E��;����˵�]ۼ��̻��GӔ����ci�*P�:�@�ShL��۷N�r��^��p��͠�#�-��wq���u�$;�^��x�3�0��Jvf8���v����{��+5��;�����E�lӔC�Ρ�0j�Ƿ ����n3(�zh�8Ko��]��޾�F��ʖ�Ȥ�O��UTQ&��������b�J��\ �X�+Y,F���R�U��Ym++(�
Ԩ�e�!m��ZȲV�QV����DUŸJ�lc*µF)FT*DV�UE0�((����.�-�K(Ȉ�ER�(Q���Vآ��ʬT�������� �+X)m�,@[j��RUc�0�+�Q`�mZ�ĩF"
*�1PE��k+
����#EkV"��"J�b�Ĉ�)mQ�(��,QTYm�ZT�e`��#p�cR�(�X�0�Ų
�ˌ`TAa��Y����E�DH�QH��J���b���K��"���X�jJ
2)Uh�E�b��(°���QA��e��a0ʬ���Մ��Q�aYD+�-(,Q����R�(�X
()�p�.Ƞ�(�Y�b��  *����j�<x*�.E
W9O&fa�%f�',yIi��y�9YکtAN4�mF��4��TV�7PԵ�t��N�}�}U�R��y�k�L^�>�D ?����'Yu���9���;^^�'i�<41H`YQOh��e5��EҗYmMT�}M�1Ss;(G,���*F�o�h!���!��w[T��O���]�m����x�+���F�T�o0���Ƅ7�i��]��ù9�7��s�kzP�5s8��C>䠮�����ݷ]j>%��x{r6�b9êu��$咻T}v��WCu����y��A�|L!���A�]ԕY���K5m!���L��Χ*�'6\Gu1gz�1o��Q�����W�^\��-ܩ N�J��EyKt>���L$]!�����K���0;��X>�\�e��2[ȸG�����Ȅ�ݲk�^��Vd]����I�o�Ep�0�ْ!�r�J� ;�j�Q�"�1.�㱱���{#�'�t���v$ׯ|%(�Ɨ�Y�`b��Y#�5��& �B=~8�,yl,�{!��)���p`*��${�����"����+(�!��x{-2�^d_?i�Ǧu�ܕ��J��vܧ(��̈́�Kz.%]ոvsepT#ιE^�,�kB��gc�-Ք(q�{0̩�>�*�Q�]Z�+�Z�����]ᭋ����~%�����;�K귊�U��79��v�:�e��wr��{��G��;�]��2*T�+vBu#ؠ�@�3�vQwL-�ۖ&�ρ�[g��f/X�D�qvʾ��_m�{|*}O�1٬��v%t�9Q����#�Vܡ�st},ž�֖���h���ԡ�{e*;q���o��Sӵs����Λ���}����Ԓ_��p�z�{��X#�B�Z��ty�-�{;��3�W]����\^�;o��;Z,^���f�/Spe�Y
�f�r6P|�������5Ov�t*u,?Xϵ�U������_�i�E��7J��-�2��7Z�w�N�K� 1ST���	���aÞ�w��H��R�yz�@���v��1F**�s6g��X�wa��EBw�w;B����.���������<�[΋479�Nz��b�t�)��'��E,n"X���Ld�7�/m�
X�'\W}�q�oQf���4�Rw-P^oVy��춗L��#E�bZU�4��w�e
�/�mԺq��c+�c��q>��2f�����W��Tr�No�V�=}�n��69�m��NM�{�ʕ�,x:��S+k�2N����pi�<�PԔ�j�ϸ@�> +��\�[jY����Z�y8Y�C������5e���Iݿe[w��P5�At6�n����5򮶳3��ƹ)Y�ZL��@5�9�w��| ��Y�$�*:N
����;/uj3�xSF.���jϼks�6�"1�DX-{T�y�d=Y
�_��(�e*^�B|�ݒ��o�H�a��,Q�'�dN��sJ��6'�T�l����<��ъ��9�l�*�,�;ǧݻꜦ%���zMV�pA��XzB�z�%�:�Q"���b.�۪e�uh�X.�Om�Mr1���/U�V�V��tuڀa*�;����7L�X�>����ð��n�mW>|�%�["!=Y{u/�U{%Vz�U���.?p�#��rbWA�Q���Fvi��o9��[{a�.6�x��B���@��y�� r� S���Bp��T�����ǩ����Ⱥ��gf���'}b�!}����ۃh��N���{@U�%��9�X�����z�^�F~�Cx��[�`S%7I����ޠ`F9Qq\:�)2cGs�9YĆ-ol΂8t�x����7�vr!���St��t^&Ɠ�F���R��뀎@m'G��c��z'�Cf�rWwIq�'���wK�/�f�3Om�'��v�0Zp�jE�e���1�@C1U�"��O��5;����e"��Y��՛��]��B�} /��܋��¹.���԰q�&*�rqe�9zf�)Gs��79}�Dz$�����]Enɟ�+��7v���og!�v�l{:��������]e�9��n�̵Ϟj�u�
�q�� C��d󛀶a_�U���qLo��r�@�n#������Os�Cޘm
���U�8;)�:��Hu�TN�SPh�{�����h�b*z��8o�ɝ�~N�,��z��^���?Fу~^P��PV_�b�;Ǣ��d*V��vz0<L�W0;v�*x�̘��l�%;���Yf����Fy�f�(L���l{��+�b�Ë�e�w�s=�b�0W\�,0��銅�pxT+=oe��ͦwy�=,������\#�1�֌�lEMs��pg��N
���3��Snʟ w�5TwtL	&��QT"n�v�pY�ާQ�E�ʡq��ɦb�@�d�К�|��1���L��+�@�0R�Z0!�r�q�N��W��V��PT��B�	=4�D��O�ȓ�T��uK�כ�ɻ	,z��0�z�aa�a�y��j��T�� *O��̸^FR����ݭ�����g"��IB���x9h�}��v���کg�k59䱢�V�u��f�J���S��������k*��н�:rjJ\9[�7�z��O+�ak޸Nʸ�
�Q��L�i�=�*{&E���{��zbi(ML١�3�ge�x\���
)d�;�mSmڨ��7BiZe=�扤����VdZ�Nٔ�D<����֍0�X3%{2�&�|)id�*�m�z�5�K�|ӧ���)��L���lu�m0��ޙ��g�v�0�2Ói��r��k��~�k�� �R<�c�bg���]�Gd���]�~:��_U�Uħ1�0n,
�:o�YB�2�z�E�VQ٧Z*�[�c�C `෕\a���͘N{g=��G��Rf}k��ɹ*'�+E�g�yc��n��n@Q����B9eG/t�{Q�֭�z�G{���m��p�-�̥�����>�>WWr.�����*aɌ���u'Ulp�d���s^��s!>������/�Lׄ.�'��A]~HT�nۮ1q;�x{e�a<���X�oL���Ƞུ
u���{:]V��e�B�%��]�N� ��˩<��/oW�y�=�5�H��Uv����t���[�_�����+T�ٖEZ��4�&�=3��x���^;g݀k� �Hv�v��3�Y���b&>ŀ`�Y�(��XS�mf-����݊M���]�Ѯ�QvI:Њh]F��p�׹y�x�6S��
S]�sQ�O�	�����=����Wf�:�g\��a�[F�2�ˑ�d��R`V_{��DD����z�_�}�*0F�@1�+�Pw�X6�U��Q�Ky	l�EX&�m�����j�*]^��`��ḩp�4ƴ�A��t��Cν&5]8n��酻�ΙX_3�sH�螭�d�w�	K�z߆��ZL�40������t_���9�*M��o7p�r�k͊�F�����=�U���i�<�G��5x��H2*r�Ɨt١��\g`4%d�j�mâ,0eP3:G�;��m�d�a�������<��`�wg�?f1�s��K%�#E��l�8##���Q����7��m����MC�{uy��;C�lS�Kg!�`�C7C��=�z�,�C/�����w���R_�X3���s�ߋ�8�cz���+uB�r��=ө�SB�׵�x �oQo�]^
�A��u6=���F��=d(6����N��wf
Żv��ҭb>�OR=ɱ,f�o��!��s�7%v-���4*��z��������\x?.2����#�Qj�u�sf��1��૬' �;�J�q@-�y�5f{�j1l�TH�YwE���ޒ�f�Wvw��m
2����������Ҟ��KG��׮�b��ٙڧ6�3��'KعV[Zz����d�m֮_{�v�kP��$΃=PGͫ{=�����g24&\�h�5-�Ө*�Ҥ6۾:�����Xz݋�S�r��b��aK���⽚[,k�g-��47#��T碦��4W�ޗ� �Rss��hV{1!{B���NJSe�|��Rc\Wu�`�����pWN_a�y�����ɪF�~���!5*�4!�Z�PD�n�ӏ�Nc��q>�L�XF�jWg'���Z�1WL��cz*)��J�Up�.%WܪA�zsf��������Z�V���f�	@�lowS�S�!^;�+ȩ��>�MOdTS~4�X���2��D�{��)`�eQUg��v�ђhP!��D]:�z�� `
]�R3N4��߁��}��<=ǯ��0O�u����`�|.����6C������T��r�vY����0pW�f�(	Mc�����*m��j��CZ����sr��H��������3t��Ys2��sWD%�P,a҂�U
Jqt�߉�r�UA�~�{���|5؂�&Ld�I�]P�+s�^U�$�vt�����P�Np57 �ySJs#�4��<�ޤf�+UZ��+��\���T5�8Miĺjٸ' g�ǟ;�:����ݗh���O�s�J���,X��-�<����J�G�5楖��]W
'qB�����=�4���� ���q����*��//11��h.�0nZ E���N�A�ܫ1܎��IL��6}������6���]y��0[�˞�XQ�Z�;�Za��t�����m�l�[rbۍ��N�sE��6n-Cv7��I�ͣ�=Qyv�{�Qfi�Zj�n�{iƸ�;E�4�p<ͼV�nyѻ-�h�5�L[��C����S�T�J�;N.�=�o�Պ���crz\W�O*�3�N��C��ȇ��i�p�����}WBp����k�h�`�q��� ,p��=���Q��r5�1�9Xѧ��!�wkC˳X��Y��P�q�Qؙ^i�r�gБ2*�pA;���K�D�U���Uf����f��Z�4،�/l��̨�H{<���k��yB_��f#���v+�����[s�i�Cy���ӕ���u��4)��T����*U1վf�,�6��]g|�ȱ��gI�fm\͏8:�oYb�-�)��qdX9�xA3M*�_��T'	�1� '���y�$J��E��1A{1�����ӥ1��OM9{�f���\�J��
z+X�|7�G�4�L@��:mX��;�����;$�Ji]�iꙩ�S�5��֥
+�(�c�=:/y��Z_[[���ޝr�˵}I���4j:q����T���S�}_}�U}{5��r���vL���ьJo��Pĭ�f�SrC��pW� c�g�����N�)�O]t��%����?&6��o;��b�e(F�d;0u�J�\�b�O���0�y^tq9��a�0��AKԖ�e�~4�j.1VӮgpD���-�{(M碯F��o/H��F�KÖ�߁�R�m҂�V`����dZ�z�+�T��<�3����=�J�D�l�.�0��0��Y'��!��v�sa��'��F�eD�1A�r}�7C��q�L�W")��Z4��C:�̄ri�=IB(�в�]�K,�Q&�#vr�REn+s'�[��-W��c�����po���	�cw�1�B�0�r���*[yQ�9�'��)⫅&_/�׫DN	���*0�!�Rrۋ�=�k�1���io����8�����<'B��y�O�����9�����}�|O |������-C�#{�O�e�5�Y����*���PR鮥�Sڪx��^^H�k�@P�R�h��Kc�L��۴�^��i
Q�L���2���}��\T�a�v��KN�ݧOQK�{ʎW\�d �Q�},�L�\7B!<�ФNӔ\�.��B)��ē�jK;Rf[���mH5�t�h.p0�lF�޿��vo�WޏG�ށw���ڕ��Of��ct���**N�=�;Ю��]�K���L9�a�+���u��ӯTb��wppi�C\KͥΘ�Vf�**J�ĺ	��]���y�{ ��������(�]q��,����r��+��t��el˔��Y��ӭԍ4�u�"#�36��z���<�񄋄Y^H�>&2�w�aA޶����-����Iח0,�r�]t��j��)νh�c�5uTK��Q����k&P��ʔ��x�}n��X�ud����9��o���mĢ�m�=y��֋3�w!L�]�Cr���V��kI�Pz�j0fוz�רdU�v�M[�|�N9�Vl!�\\i��Y&�_@�6ߜ�x��,PÕX�*Y�c7{<�
s5�F扝�C��zEוA�F�A`:u��sN#�y���/|Ryc�~b|v���K���YD*��P-!Od��Fߝa��T�>C���aoV���fd�^�x�gg٭T{W���8�gD�B2�N�FF����D9�@�߽�O}��p� e^��(�o�N���wU��l�n�j2�f��M3a�����u�י�.�z�̤�����:�EDDUnu��4nԴ�����+�Q]&�|�|1]aN�y�K�z�\��a�쾤�V8w[��'Q��q�x:�����Wd���%E�};�a�	���%C��A���&��6[�@�2W]��\Ѭʖ�`芬m��Kgoyއ7��	���&����nM�8l �F���;k�˸�hP9v-m�#�#�EÊ�0o3<u�b(j��O�v�&�s�e,*��1���p�10��� ��m-TU^�oJ�=��u�n:�Z�q�	4�i�+
J���5�$o�K	M���yp�u��˚M%u�)�d:�cmw� ��C�q�{*�pn3vҽ����P�ܝ�J���ps���B���+˕����Y���W�C�3}yB{�wB�|w�%�+T孡g��xun���й�y?�c�㷆�j���:�jU�)�f�i���ܟў�a滉�C+X˧K.�4Ȇ��=�A�O�{o;�0��,nm�3;�"�c�z0v�ޅ��3N+Ȁ��jyܥ�4��,Z���x�k1v�r4.*��Uwɺi.��]�E_�[6N���qg�a�è�֦�SEZU�L�332�������B�����\X����M��ތ���D���̩��<��}o�%�65�&%[�p����ݾͳ��,����T�R�\�ُ�{8>�â2�tq���0�VF��܂Lo���i�<#y-A���T0�w|�)|��v���[Gv�w��ˊ�{.;^�ۦ���cP���z�O8�Y�t,.Vimdo�q��U����{��vgY��J�kͤ��B&�\T1o�C�2I�vgL����nV����/A��� I�-m��零`���/��4k�!oil�n�U��m�X���O��,e�͏�]�C-v��A��]¸��Ks%B5��}�N_ҹS��:㱋$zWC��������(6+-�������WN�2���|��#T�Χ��6m�[J�w,��C/���v(���r�R�W�2aYS빁~ vs{S~JȯN���|y�=�����U��/��- �u˳{T��ݛ�-
�򯈀�g������UW.���z�wWћ��,��M��0�œDf���nMO��	�xĦ>��!�h�9vN���<Z�V���Yb=�_V������v�yvG�Kʾ�7m�:_vJ���{�Z���Wq[+z#Dk�ku���"�=S���m�7�(QG��8�W?z{r����A�����Cp� g<۹R�*��̥l�5ٕ˨h��<.>8c̺,.B���\1�4Q��γ����YPLyd)��<��.A���JX{��~�9�"��PD1h("��UE�l��U�L0ª"J����`�kZ�V(�m�� �+F��TX,R)b��5)Z�mU#m�%b��b���U�L4QE���"ե��*
E��"��Z���E��"�*��Ra!DV"�1"�eb"*�J*(�11p�1#"�"����dUE�RPdY"�*��E�0U��X�,U�(�6�(����X��`�ڱET@U`(,UYP�@Hb�U�(�F6��QV��V
,Q����"�X�DTX���**�Y�(�-����U1R(�"�J�UPE
GB�D�Eb��
 ���R,�`�X�EX�QDb�",k*
�F@F1"�b�Q �X
*�0U�p�AAdQe�b�-�����1bőH��E��*��<����ώ42��㝍a������t�e��W��z�{�Z���
7�C]'yFBC6�m��B��n�dU����z=��A��UP�uP@�u���g�W��Ӵ<6�MBPo��gE��6(\�FLV��z������Ud/� ���5ᗩ���8E��!4-n[tB{�w�n���:s���尷���{�r,w��Z+����2�����nA��u@�Ë�û�";��M�@]%u������,bE�j�"x���9��eu���gRNL; �skd�k5�[2tVpiܰ�T�ڷ������g24&\�oN��u�i�]�NÝ�wg�w����YD���zT�u�fy���e�s�g-��479�K�
.s����g���N�a�HTt��B��rR�/m��,r��h��+�u2v�0u�sDV���\���4�lK����1w�`�"y�R���㏽N�] �V�͆9��z(����z(L�'���ʗ�;Q�]R\*�1u�Ϣ�s�0��7��/L\����[�����t]uwnr+�p E"��dӦ����\S,Y�ݓ.�v���V�C�Ģ"g������i�F,#I��q. Q�T�%-9�|n���H� o�%��:{tQ�ջ�n*�]]�N�.��":��t��TX�ή\z��5ѥjV}sfEI�뺖�yv�Q#{FgE���J�(tW�������;s�n%�D{ވ��^���s�Y�S.�D;�j]��� R}�m�8�ϩ�s�^�Rr�a��y8�v��:����:�4��/��l��t��������shM�3It�9�lF9���)OV)���s���jJ���n�h����V\̷��o�y⪫��_���gC��<������kƖ7죾\�u��Elu����o�=�z�ڼ����+Z���s�$^�vL�r�گ0��5Ǐ���v/"�^�[��
d{X���	��O��s9}�r�K���,��3�b��t+(��\���Q����������Mn(\,�`k�l{��7k��!�.U�������cyX6k5]'��r��!d�w�Y �Tz{s���vM����ӹ�}�Ù��؍�oF��{|*n-��P�oU<�N|�����_��;�F��N��]*LW�Mr�@�i��a7�Ǵ�Y8x���9��q�8��溕*P~�����|� vxH�񩦦��?i�qLoNC�4k��"�(>.URF�os !%������w���d��2ڥ���<bz�z���_s��:`8#j�/_��K^͓)ܗ���r��qfnHg�cis��$5+5�Eקz�+�����,�{�#+�\��e;�ݒ$���v(͚��������͝K����G�M�8:W�<���x���zL�V��3\n�9�r�G%�/�����$�;N9�F��d0�aL��JC���~�c0_���<����9��yBY<���A/�,�NW�@oo��
���A�R�T�c���k�a<��Ϗz���2�OT��M����ͤ6-j,^z��ȉ`*"��+�@Ai��Y3}�U���e;g����J��[�/������6�����V���Sȴ�"@��zfQ��L����M�
H=���p�|GUk���e��R�t�/�B2�-�=��f.V�mm�`����/,]3v��I��!-��R'�𱃟ּuS�ȵy]q��0.s"q�-�̹��Ox5
]�U�Rۻ����0Y��GÆ����/�|6�-Ei�����Y�Y���}�S"�ȊR��h�:����{��&x(��aؤ3j�#I�B�V:���e����������e8*r S��Ɇ�DT=:b��Z4���d��������$�j؃�^)7m=�}�|�()�(���%z��+���J9ݬ���ʞABm�b���F��=�B'��^�~��`���8�̧�V:��i��<f��f d�x� ]\;b_I/���(-0܆�d&���XJ�,jw���ꪫ�~�+v�$�Gѕ�EF�2ak�	j����`�i�~�hs:��Q����q�)y���Y�%��{n���/����W��u���a3"��=S9��|p^�t.,�	����I�t�^�b�o�����G���
����^�'=�=��E*�aZ�j�����+��W%�Ht6��@u|�'O���:�D=4WR��	\ft�逹�(�q��Nc0�baQRtdC�����:��M���.��s��Ȣ��'}�r�S5�*Zxf���\�o�fa��TT�#���0�-�n�Y4�{��Yy������g+C܍�=��'Q�Lk��=΀�*5�`�0A=���q��Q:�`�/ܷ�w��aV@w�;�\3�ßl����:-���n�#*5�j�f�܊{���<����4F��dp{3���P�k5��@�EJ��`ۮyV)�uλ�ën��2^f���H1P�Fv�e+�	�o��T�5ժ*kI�Pz��U:�t���>��+Ges��r��q�]� :��]m0��;�]&��s��sQ�O�a�h���e�L1���d���qC&#�+���q�5A]���vqu*a;��`���k�����ޮg��^!����oON{M���r��	v�����{<۱[�(�d�����w[�30y�S=�hm�1���($�5/~���Θ7�N{:NJ�pK��'���UB��@�|�,��MO��cE��b�1B-ԣ]/���ΆTq��`I��ȺfPr�"����s`u�.酽P�[ŝ��<��[7�`�E�kqҙ����ʼ�<}B�߂�^�a��DN��B���Ug��wVGO>[{b�O?lԇ�Y�2���n�AX4����SP����১j�_[�^I{��w��;F=U���wVi���}z�L:#�ł?$*�n9�����ԬΗ�җN�f����ؗ�G�"�UM��������˃�B�c6��v�q]2a��j+'�.S�u=[����\�R�o���H���p�|V��s]Qc�I�B����}k�U=nR>�ӳ�P���=^^gå��ڷ����vy���|�91���:늺�C΃��es!��{�V�Ɏ��;�fHN\�Z'��yS���'�:,k�g-��E�75���t�����Z���7�z��Np=k�>+]֞��^T8見Tx����������*�[\��]GL5�3$��|�a���ӫ��Sp�>w�������ĬW6�'M�0�)lW��I��)[���/jޜ�T::|�O�;����m��?za�����B���O��+$�d�6^�1�Tk�����q����Mk���N�W�t�Q�S^�^t�bZU�i��ز�A�6�V�U�1Li����r�w�0۴�W��0.�2����TSeT����\J�3�(7G#��vƇ�#�Q�N��b�(8��/=n�ed3�*<�B�K��7K���|�xc�	��1��ֶ�x߲�yS[H���f�/����2&����K�8_���Dx��8��n���W�yv��;���h({���w��0�4678k��#ԪXc�)�%r-��.�sۘ7��{&���f��xk�ۮ��C����j�\�v]��s�a�����bv��S�q�o����=�]٧`V�Uz�Eo/�d�\V7�O�33_�*�X���p�3�yi�e�����I4��&��&rQ���+ㆡ��|8ސj�c��@�[^K"(�z��Nړ�_���:���A��t���=��Ζ*P�;�@�c<�YR��t�`��Vn���/���I�|,a7��ᒯ���sr\FWel���_8⺚.v��Τ�}Sn��7�� @n�-9���\ڛ�էr���1B'V�=�in�M�|Il'y:U��c����⋶��U�Aw}G�TɅ�K��;h[��=3�UW�U��}N6�����0_��2ݸݜ��4Q�sf�ס��b���>�C�{���rRu���d�U�����>�RFGKe�#;�ލ��oo���I�>z'fm�y�8#p�zz�pb�?^EEE����&��yU!��v�q�v�<,{J�p$�*ᑓPE&m\��o
�Sx(�~ް��&�����������O9��zU������*�����<��O��i���ԑ�ò;�c�/,pi��q�N��[ӷhç�~S�rW 7�T��k�ޥ[.��x8�Be&C���~���(K�<��!6��Mze�q���͑L�7�����q���1�2`E���2߾T�c��3��'�N�'�(g�յ���c�S�ej{��>>���K !^,� �� ha�d�m��q��͙�O`ߥ'~�S�3|��~��X#�a�Kmd�*nH�b�0Ȑ�uۥQ8Y�h���:O�m�F�V��L��q�����|j���~�*��K��ם���}%���]���ј��>&��������f�R�����q��/z��x{dڍ{m�y� ">��=љ3%����8$Q���Ø���V�<6��a��û	4���j����M�sR��ip��q�FDj���k�PJ�K��ڞ;�G���M%ڞk��.O��
8��|)ZPc����Z��N�-^W���+� �\8��g:��8QK�%l��{�}�}_a�Ys3�
%�ƌ��B(Ϋ�BW��^;�>&���p��}��͚���/d����Syf�90�JS��n7��]��(s95&�$���Rq&��rXc�j��	�� ���d�W")��5�L8RWC���b��Ύ(�ο�.���{v|�2�AʌSa�"���̕�lt�;�..M�h7����ϟ��_�w/bD{�c0e�~���EJu��[��/��]T��;����Ϧ,�i�c���{��v^��ȫħ�c�}�x����܎� F��U�L���1���X	ϴ�g&�mqӆ\v;�����4�\d��Jk"� T_Sr�v{�n�S�3݂��Χ%���y�9v�9�M5�վU�ct�9�ATQ[Y�g��X{�x+�3	���fPI.�o�]� ˈ���Ƅ6:���)�Vs�9�U��/ʊ��duR�dB�n5�����m��v%S�*��E��8]G��$Ԙ4`���x���	[{�;�5hw��E	�����lJN��4�$N�Q�g��[��O3>����L�5�6�k����7��3{Pfh}���]ו�u��;�z�L�\�\����f�f��cS��W���k�?=ofcqA�+ofn1�s�l1g��)�r��q\����k�`��2�7U��iZ7`aRNS���.у�5���k��ϲL��y:�w��o��Su�Z�L�GN�ɱ��U�>]�Y�4��AQ��ς��5��Ƀ�V#�޿���Y���X��JO"�N�	�)��NT�_��A��"7��ᮭP5�8, �h�����d��0��c���j�1��f�[�"�%�\q�xff,�m���/ڬZL�/w���3�b��j��|w�]K�_�h��& u��T!�dBX��[9F��5L`~1�E^��%�)Լ����]�+
�YL:���T�B��0��ۇDXb�B�z�!؈�Y�5�|/�w�w�I�M���bZ�!�uy����PΊ b�cd�dh�>�lu@]
��9�=�����Dp��E�H��˔0�fs7=A)z��l޻��[���p̲�c���NT����v��p�������MA���g�ub�<H��
���[�͛�>�'c´ú�3sE�b��4�i�=OT�7�.����v�y�B�FZ&�b���ya�0��|�ф�t�)�=���ly#x-��ʐ.(qb�霴K�떑�=�72t���g3[!�}�����{Sϒ��3-w�9ܾ��=��%̙��j�=ӾN����V��o�l�Z"ݐ����u�y�XM��+,�0��+��8���wc�Y1�վ�fpk��T!���?v-���Ыtݬ��f���j)n@q��9;h;�N�N��m[��ylwg�̍	�71��[Y�^#'��>}Zr�V���b���s6g���A����*�������r���B�3�(�V�{�7��P���r�BD�줧�x�;Xd7�:��O��p��� c��usỖ#����4b�a���3m]�cՕ���O,B�vV�k��6�y�&���˒���a���k��tc&`\7NfP��z�/uj3�xSb�:����1u|���՜���jŹ�0�=l���_<�C����B�4��&ΐe+<L&b�Ov�����M�ɹ>�'���<�lV��)v� S�����S�ȯzS�BM+w������/C=S�z�F���.��o9�g��:}����6ª�$L�^V�['Z7����a��t%���v����p�<ܱ/`
s�F��B�%qYbt�^v :K9݇6�
Q�V�ڜ�e�9�R
�m�fJ���/)d�R��%�Ս��v���Pʵ5-�&+�� fJ�w����K�g8�I� ޾Eu�I��^�T�;x����L�
]�N��4��H�}!�oU�a�M`�2,|FN�r��y�ԝv�%�S�d��M�x�ނzP��yr�n�o�N4j*�G\m*�N�� o�������1�B�!��3^��`5�r��`��|�����>�	�����+[V2^+���e�r��b��Y�L�N�9Ob����2'T���a�XR9�h0q�J9��eJr�wvńgk��<�$��0.q'�Ѽ������9]�T8m-�2aj���4�V���~�=G�����1���/~�&-sL=B��2�I�ƻ)g�O�v�@�(e�Mr��-b��G�e�t�I��Pwm��p�9�|v�df^"��Y	#�Ρ�0�g�.����]^����yf��M�ܤ�&d��6�����-���L��[P-��8��p��[9ַlKgi�81O z���R̹M���βt�y��^WfJl�)}I��]�\V,T�x�*�o]%�֢����.cD;X�_gE��ru����F�W/O��*��48ӫf⾡���z]+�K� ���wv�D�z�Wx�h���z��4w�d-t�)�#�t�l-�׺ 	��J��@��/�Z�i���9�{FoY�*����}*�t���F��4l;�8�	�Υ��|�A?�Y/+5Z9ۥ*�0�NrW՜9
s&�ż4�E���] ��fR��;��F�Y�s�DOPڵ�jө��d3ٝ�J��},h��5j+��os�۱�ZWD�j��&-|���Z2�ԇ;Z#�T�� �Ҝx��3��ص����螵9�z��wY��|�� J���G���:�A]nT�+b`%6��I{u,����(��T���$C!�|�]u�=;l[�~g�E�դv�={(2��>�;�O��Wt�
E���X��ws����
�$��`�n�����h��^V*�jK|f)��G��,c��Zkŉ1���~.�s*���&�/k%�nk3WO��Եv+�4��v�bT2�;9�ݛ��YȞ@��s����'���;���f>�/�7�ֹwJJ�+j�k��g9�oG7s$5��͚��}�/���b�"�c+�Y�:�S�1�/l�-2�i�R�d��}���M1������+]s��ำ.�U�Ŝ��)�AЅ4D�]���S���Gq�&�M��̬��p����E+�GF���� >�e�k��)�3I˛Iq���6W'�iǗ+4�����y�m�7to��plf����p6m���-��`@��S��oć*Fm�y�m��D!� B��aTEY"$�PF
��b��PH����� �#A����Xň��E"!_S��ȰQA������%�`��PX�b(��H,QH���b��#H�*ň�R,R��1�0Q`��#mH�%A���**��Vł�Q��UDk!DX�*"1VE�,V �"���ʱTAV)�H��$U���łȤc#Q1j�FA�Y(�b"�UR8�UE�$++F(�QH�
*��EdAEY�X�bʁQE������LZ�Tb�`� Ŋ,UQ`���� �R,UQUIAAE�����X���DQb,����,QQ"�	X���b��b�������J"1cTUD�
��FEY
����E��qIT`���QU���U`�d��(� � ��H�V1D@QE#=�kx�n���q�_6;U�\k:ةD»��jJ���Č�G}����Qή�W3�x%���� ћ=`��R��.��"#�
%����!��?��kX�Ǯ���y?�ʵ$�|�����K��܍6n9�OK=a�Z�j��/����e8��-����o]K9�U�:���TV�^�9��s��f��$GG��N��	�q���+ㆡ^��1��A�Z%��<x��)v�ݞᗝ��i0�� ���։�j�f��q�-靛��_�X0]#��xR��"-.��"l��;��R�^��{j{@Cj?x��YIN�\8�X�,��b�7cz��1�Yƨ_(N�Qjs�[���c�]��"1J��z��,9���؍WX3'a��]>�gg��)�w=�}�r!���İ{�ǔ�S�R���C�t��Utn�^~��r����1�G61
�z�7���
H8לhs�
l'YhI�����		^��6�+��of�>��u��-�T���7��~�cF�3p��*�U83��yؙU柇eS���H�jY�`�
WV�7��8.*��\s�UC�/6�9ҭ�^v<D�(]rR��Oñ�f^P����G�+�۶�F���[Y�UG:h�u
��u��W�t�u$񑵒n�K�ނ����[����E_+�h>���6�T6�Z��:u�y��1i��<�{����j��G6�ڄ��T[{t��й�KWI�$E	���f�nt�U�UV%ޞr4(�]�gB��/C->Y]GZz�ن�?�|*Pg��M�Ά/;	W�8e�� �A���p������<�@��X����9�� B�"�����-�w]\��ѼҺ�����~:y�_9�ϔ�W��^Jk�Z��6%R�S����LW����z y�6�V#b�1}~��\u?���唽Q�`]�~�P��4���YG���|�9W�P��*v)t��$�á#�m�|)L�r"l`�Nv��1Vӣ�7�<�v��� ���j�3W��Ԉ���4�0�˙�J�Y'�,p�7hEx��`fK�S�l捗�v�B�F�M=�\@��
 �"1��c��	��T�,��Pf�~)��N���=ױ�ܮ�/$ܿf�6�	�� fKW")��5�L8RR'+��������j�T6AJkDIC�Q�o��"���̕�lt��5�p�N�\�������싮�n1X�F'�k{��ee�J
C�b��3ce����a.d~���^3��Z����"w-�=�{}ܬqH1�6�>�&xI}����]e��o�'��f�U���+V�n�Eoj�֫�د��׺��M��f��铗��=�Lc^W(^�.�c�w�ޞ������faneQ��줈˨F������g^�q�c{F��ZJ����0Y�=��k�S����Z< u���U[��R��U����Ӝ���W�^�ח���,x1°L���X�)����@�}�Wm��Z���$\q�y�G,��8��Úoj2#Z�ʢ���baQRtd3�3�u7)��ó�8z���H�^�~���Q�Tf_��N[�F�/�iᚢ��g:c�EY�b���*uR�\�w@�-����B�VM]Ts�m���L=ȍ���`�u���=����:�x
y1VhN~�j��[���ۺ��ʔ�JUĎ��}���86zU�w��o��Q��ɍ��v앦�>Emfاp��c4\��,��4�ʌ�
�5� ���A��`���0���5�vV1Wk=u��"��a��i�4ɶ��ܥK�l��p?��U�]U�uT�[p�[˯n���;�s��
r��V�l�O`\JQp��o�p�0,(2�v�7�e.V�=��eG@2�k*X��I�]�8E�U�Q�P�U��Q]��[ �X�a虃6�M\�rr�i�ں�ed�nv����`���S��c#f��3��!{�ś��o�ѠP�x��A��b6Hw5o-�rb��졉��.�R�'
�[
׋�8���S�����/L�;"[��V����`��R'-+���JJw����4�^��V1�<�YFb�<=�Sm@Q	
{ �������R.a� ��s|q�����v�A,�9<�m�C�}Z0�!��q�
�AJ�ZP��0v�Iy���S��ݰ�pF`:Y�^X�����/Ƽ~X��PNج~��MBK�w����=�rޯ��>����E�^�mޚ�U'{���[�2���h� �V���Kc��o9��qf����֐�{��g����`�}��6
حnH��b���.5�u��Z�;��9쑆��2=�b���y����^wG�>�I�� �w��*l�A�s�u���y}='`��V�������C���1�Lm��;�S��a�og�!�������Ɏɼ��T�5�+i��OPz����b(�E@�.f��&2�b��`§kg\O�7hb�a>��@e�]��D�V�*��GM��H����)���w��a����r�QGT]�8�e�&̹���~������TY���NEU1��j�#Q�`)�k`B
� ����~Jr[d�.��F�zM���ͣ�"B͒��/U�e��{�\k
f���u1��y�X�_K�w0[�Re�(.�_6a�ZH��Iܮ�ѾXN�U��+jͭ�:�w-������(��w��]�\�Ȼ�]�Q��ξ��&v���}�d�Xڊq\l^���ֹU��1�ш��d��t�T)����:���\*�٫�W+��^��42�/0�L�Nsf�Z�E�[�YY�s�!^T8P����t��TS�o�><�:]��I�<��fPݜ�s��&�:E0�����j�&� p0��"�WT��]�}�.�{po�
Hwi��n���RUN�ƺѠ,n��B�y͐�%�&��$���`3�4����zG{��c�1)��Fuw�]x���"�Im}�O
�;�Y��3����2J���"ǆ�P_���2��Lg��vϚ�w�Y�4��e왙�Օc�PJw�s��JY�p�8*�g&Ju;6�`�,�W�6�F|Q��ug�I�!������9�O��������^������W�:]{������chJ����Jn��f�#c2� ����.�:�8���9�/�� �ۍ��7\8�őa�t�[t3k���Ҙ��S�ƽתB�^/Rz>O�.�d2�.�/3��Xs6�[���ݜ���\���-Əw�4ef(�)�a�;,9���C�b��ǽ�9z�{}��Іr�ݢqq=�ܚ"λ;�������~��0�S��SZ�A�}�2���c����/�ђ ���H�3��dj����!�$õ�F���6�͠A}H����4�޷���]I��3l%FV䲞R��T���>7K�tn�^~��r��T���;o�����6�^U��f�d>����В����`�<���Ɏ��-f$��tsx�%���t����6&�83ާd,wV�g�,f������H�.tU{;/\7}�s�*��'2�B�/5wz�l�c�bU	�8���i�v|�3ab��%������C�cN�r��hQq���9z6�,���r�1����L���,B�~���YX�2cm�6,�V.]S~��}}s����I�Hvf��ʹ����x�� A��	�]1�qSï��l)�7$4,q1P�O	����K�3������U��Ms�q���tz6X/�z��틧�X *r3��6�+��A��GV��z`���^U�t�wU��;�IX�����?_\=��f���[$��$q-�>���0s�׎�u�j�3$4���''�c�zN�5Z.߂'A��Ddn�̻���e�>FR�o�|8kJ
ʲ���U�<�4T�]WzK:����h��ƽ��lcvÈiy�j�=a74s�c{	�;n�R��/\O|��׉켧(%��A� ��^�����<J�667uj�I'��,�t�����+�CJ���Y��ǭfB�r_7�&gq�%���gv])2-
hڝ������w��U�p~�-E?�p+U?pP �Dc���<���&D�K�Hf�Ѿ3H?q��6�r���|�SY�T�j��	��l��&Z�������z��`�ɞ���?\��Bg�T���V�e��(d�\�ɂ�C�En+�ٮo|%�m0�����V��c�+�g���A��A��cy_�#{�3Ꭿn�/�:*S�\.�|�`�a:���9C�r|@���G�f�Q|����.u�.O�\J���o�x8W��Z< ���
��*2��e�cCm�ݨ׉�Ӣ��O��f�k�8F�b�Ɉ��VSYA���V{t糲�T���]@[s&P�	m�1�I�F�Oz�!���!'FC�u�WWN1Z+��t-wwf�2cT
��f��N[�V�8�|:�R����/�U'f�!p�2k��m���M����j�-�n��}3q��{�l1p{m��9J���yT�����^o�緈�nN��7`�d�V)�S�AJ����}���86Sz�6��E*��E�v���#	���BE������'��Z����ܫJ�*��1�9ښ*l���YL%U�sI��-�%��5�t�6H۲޾W;vfjwܫl�>w�UB붌	��}]r;X���G�G0��1��Ol
ʹҍam۬��e�fe�}���`,��v~�QZ��˘��ʐfCM�0R|GF�؝Q0vj�`�L��D>tSx���b��}\�d[��'��:���4.y	�o�ϕ/v���p;�-�栍1���j�[�JuE\!�jA\�jcU�n���*;<�����m�����<�?z�n�(��޵}���40�G����/�'��ͥі�w��O�-r���7�D����Y�m�:��|�X�ւY�#\̡�H���dk�ǆëh;������<���:A�Աz������Y���)}�u{!����>и�cf(u��[��$��M��������HuKo��ed����ץ,l�R�]]]q�~xoOY��V�652g���x���j�����}�tڞ4ؘ1Kks�/4q�3�s^[s�:��HS5B�^�+u����)0��~�k�X�Go�����<��ݓ"�|"�*+��1W9(>N�a�p�`�V��^W�Or8Ǧ�-�ƙ(�	��%R��b�O�Y�� �Lf�.R�9�geY액વ:9����'@�?&�%J��ky�`r�ԣ|��wO��Eƣ����Ah�R9v2Q��J���w'f�=���fjR���4`Z�K}[Տt����l���YT�?.����]V�/��t0�g��R�p3:�rcmj��.���j��3Ln�3�.{�\��..���s�����w���F�yGPU�+�J���9J�H0�>��Y8�|r�x��]�n�$����bpa��Z�hns�
9�H���Β��Wx�7Xd7�^y׮���M�qat�QHh����7���E�1M0��USb��G�Q�`)�kx��	��O���;�s K�f��k�Xb9]-q^��2f�t�T �1�QLe��r�޷xeE_YCb��Z{��g>��l�%�P?��짎_<��A��,P���7Ęc;�hq\��zk�&1��k�qW↸��z�d)��/8S\����b� p>R@��4�o+c�/���
a����u�v��q�8���T�ߵ֍e�4�]!q���q���Ⱥ��{{�kZ����x��"=���R0v5����Գ��kY��V���~ω�q����C�}���8�r4Xf�+.fY �6�~[����q���(�O�318=��[GT�\Ϳ��)=�좴��({�͎�im�y̨Q>��q���(���0ڋ�$�Xg�:3.ފ�1W�\��5d�2'�Ҋ�퍦K�6�ޮ�;��dX�n���G�g��/�u��U�F��!��ԭ�������ېmxt�rTj�u^�_������zm{���~c�g	Q��&%t%h������T�?"<k�h�9��'��5���z�	��@��މ�j�f��8ŷ�96!@9=�`�zҦ�A��4}s�����+���W��8�Fօ�Pg�[2����:7��YZ��ko�;3oj�Fnu��3_��so*���O��Y�+	����<V�n#z7f�H.s����0�	A�ɞ7N���Eu�o$��>U(Y�R��{��r�@�i���&��{m[֖�\jtp�㰱�.���wCy��l_�8ױ��/ U�x{�[T��od�+=J�k����i�x�hҍ���T����ձ�h�i������m��K�e��.���q��_��&����37��KU)�,W�e�}�4���rfs]�#՛[3x�Ô��9z��P]F#]�c^d��,B�C��4\h]�&�yb�w�%J�yR��\��Y�|���~���B��b�[�S��q�b��=�����N��̺�\-���	��cCS{\�v������Z�ڎ���YG$(;��u�V��wJ�Ha����x{h��h*cü���{w/�2,��*J!T�r�G<� DŜn��L���Ԍ���0����He�t��`3�_�+]�n=K��XhX��aʹ�HѼ_X��g�E��T�Q���t�%�ee���ne|ʯ=�zr��������.��94�;o9W%�4s�
��X���,nk���J���@��JT�̶�˺�z��w��ڱ8m3��:i����:>O���!1�q����i_o����frQ�2l�8�@eL���҇{��f�ח��:��Daw����1��;G�2c�HK�9�غo��ۺu%Y��R0_Ƣ2���6�rբ
�F���	��q�
�2��o)u1��x��tV �yYOh��|F�|̜)��|	O4An:h#׸�:;����ylQ�'(��k-�Į�6{��M�@@��r �/��Dj�f�pY��ށ�λ���8{��'�/���RBz[��m�X&���-uBG=Oq�P�Ԕ+1Q:]�K�����bWq͹'C5w�����1)-�.�z�xz�\��vJ��͓�3��:������߲��7z�Mr1~�5����V]���ώe��':�pGpP��C�R�XwX�I���HL�w�
l4��W ��VP����1+˽��4(�|��렛��'��<���z&E�v�W��u.�׎����(��|�$R�͸�C��mT��5�0Dzٷn<���Zo��ܓ\��/F�ՠ�y�v��6&���l���Ta�����VB��r�W�hy��6��!%�qs3�4Ħ/�\6n�Շ��I�ɗCR�/��D6r�%"�Q����}�2uZTs���Pit,��{���KR�L�-�C�}Q���z�I��;%-&�X�M�iP���寃z;0�1��Ϭ)�n�]�f_5S��s4��9�x�c�7z����J����E\tL.�R�f���]`�ֺ��4U֧ܰ�::�C��� VOvl�V�����)[�����{t@�J-�%���f걹�fh����TO�|�^��2�	=Rұ��{Bk�U���v��Hh��1Z��A���ոT+0n/I�I]w�n�{��۞Έ�_m{����~��uɜgJ{)�<X������h��f�Ż���3�\X#�΍�N�����]��#+)��	wm#c�����j�>�!�îm[`��[�Guub�&�u"�q>ೖf,`e��g��!���/�:	>jۀe�����B���aǛR"�Y�:Pr��˳�%�g��r�ty����-���DW�Al��xA}6�*ãK��d�fvVU`��l���X飢ҵ9V��$�TP
���0bF�����H�h���
E�

��@QTX*�H��U�Db�V+����U*}�*!�b�"�Up�Q��1QQ,Qb�DV,�EF �h�0�QU1`"�Q-
*��**��d�(��E+AkEAX�A�1X��

��TET`�DEU*�"�AE�6�EF��(֨*�E�"TEH��U���A@F*�DbT(�Qb"�őER��(TX�b�DD�A�V#F$�E((*0DX���Y
���b��("*%�"*�(� �EEbE�+��(��bFH�LYU�U`�*Ŋb�*���PUFATE�((����U���D�%J"*��X� ��(+[_��G����9��g�7���`1������sCo��\�7^jR����]���
�kFeo`c+/�qh�Rg�VG}�ʯ����v��1�*�� 1lҩ��Q�?i��v|W�ګ��Jk�\]�ˬ��ۛu:��El{9V�4<E����o���ب1}~��\u=0{z�"�Fps2d�O#�.R������g�r�ҽ�H��:\N��}CıyE��׎�\�nnz�hx����}Ș[�t㧆���`�R# [t�LS$��1�|.��0����p|��^E�'�\龨^��;�|&�ȵ���Wڢԁ})�q���3O���de
���w�a�i�U@Q	8�c�P���2`0�j��J���d�ٓ�D=����\K��k���5v��l�:నb��B��U�~:J2c6��,����5��\��K0m4bl�+ޗd�.��ȭ���v�0�2Ñg��e�~�+8w�U��3��E[+5���Y�&o�hݔv�8rztʸ�10uc�+>k�U8����c�r1&T�)���>���.�0�l����J��|;à�#�h+b�Ʉ��V}Me�4�b��F�^���C�f��.L9K��4F���lx�j��~�콼�jg0�&%�zz�k�ܑ�Rg�:Q�;�2��Ǥ5;�$�p�mq�+��H_�ؗ�n�K��Ĳ�$��q���f�N��GS3v�#����T��߾��y���`�QY }�����n��Oj3Z��S����z2�~�{i�y�{�9��	����w�����qK{�l51��Zxj�y����*���[p�y�{3ם���Q���W�
�B�1f�8����)a�m�������:�yN��
�T^s�sX�|�n�~��t)��u]L�:�������	|fNk�.���U9�RE�_�#ry@�B)�NF��Rc^\�-ԩ2[&�)>
������;5e�Odc����z����au^��u�*�[��%���}�����S'�n�ىc.`t7�u=���Ȳ���$1�1ѩC4�+�j�Q�2�1.��xff,��M۴6�Vݶ�"w�&�R:݃�^V��b�x�3h׆m ���p���֣b��,\���4�ə����ae��÷������^j"�Ł'�"�Y�/�
{ �W#z�up׽|P1�'�y7ڎ,p!�z��d:�]�z�1�N�Ha�^C'�$���ꅌ�=㑝�mRv�o����Y��޺����y�h+�8���2��.0xk��8�fb�=t���zT���c%��F��n�)jv�:�l�8�^^����aI�4v�n�n��W�};rMp���a��+M%S��ZMʅ*�2�kV�ퟪ��[���#�!ч�K#C�r'A��Hx���5ז"y��e�׊��xf���J�=�KN�yo�*pM ����2Ol<NSӵN�WK��gM�*��Y�q�1��5W�/5��G�إ��4���#ڰy�HU��rW7}}�x�B_-��ȱsih��c���d���{��zj1=�����"Uj��wc;���U���y\;���G����������,����v!��f��3':���A��A�*w,u;�ͫ{=�-��v�.]��Y|v��y<+�u�u�:5Uj�_l>'"�&2�b��[
],�Iͨ�����;�\���;׏QcT�3��tY������	6�+�S���e��!�W
�
�nY�ނ⯮��~�c��k����b��TY���Ḻ��*�5���]ΔY+/���1�TNS��^i�bվUa��u�'�U��p�9� �v�eE1��Wf����7��l7;��XA�t��u�Gp{ҥ��j��e<���W�
��΅
�
�i��u^�/�JktwI��i�q�@��C��6�
YK�ss��Ӡv��Y��ְT�kk]�JrV={�
T:����Q7י�Hjl������:|5v��W������$��ѧ��jW)F�^��Ң@��hN���ǚ�͈�U��Y�ʯ�7+�މ*FY���Z�.<z�d˯>�@���U��Z�	�HfG@9�Ӝ����ދ EbG��k�����s��8N���2������
6j�%���ҢU��u���;#<��wLv�g�P��0����\c�ڪ��u�P�sS�Ve���;��fE�����N�h�uLg�e�0q�X!��w��jZ�C=�<2�e����8���j%�0$�S�uQ�(��8Ld��1+�)�8b���[�u�L!wF�f�����}&_[���;l�ւ���*� W�k�ע:]W�:����m�,_�%���T��: ��d��RT����2�/l���߹�.;[2ݸݖ�F�X�,3��ٱX����퍻N����f�N��� ��r��2�+�w8�Xs7���HV���};��-�	�o�>{�.�OڇE�lf��x�S�R���������Ac�CIQ]�����= ����|��0���t5��Mp����� c���%Q��z��#ïI��](��O7��9{�ǫ�\�u�#�G�8n������;�{X�Ym�GQ�6v��t�H��T�֏���L�&�;�=�Z%LԹEYx��Q��r�g\6�K�L&Z����}.�<�I�V����5��Gf$`�Ks	Że/����o�����?�L;�og=�)���rƍ*�@���������+�y��iR|^�qr��n)�ʨy'%�e�IyU�н���J�]y��u�L���u�6���w�d�m�g����-r�.1��(.9z��8�N5��5�H�W/Y����):�sDh���'k�*U���|e���+_���.��|7=�����!�(��މ�� �e��� Zb&*M��W���C�w���~�چyo_I�d����W�E+�����^�p]P���<�m�+��Pe�*��ſi��ˆ�3�p��l�oS[Yt�U�w���r��Ǵ�:^G��/��$q-�>�(1�cH�<�Suv�7u�1���*zqD�P�1��u"2�Od�2L8F�e���MK6�M�9�/����i�ȽB�V^3㨭��V�p������F[yf#Rfޫ|:3-^,>ŋ�I2>�kE�`�z�x!�D�u,*�S���X�Y�"�L�M%Gf���9���u��t�Xu��x<z\3���.���]F�J��� ��Ip�y���k��y��g�Xa�*OY.���^�澭:��S�5��JXyw�R�`Zr�Nv�a����rVwPK+��"7���Z�2�f�0��"o��///z{���A�p��t3��:�7*،�%1�,a
�)W��uV���S��Q�/����;�H!����4�5����"7�c>���;:*S�W8n�݆���785է3r�r����}�l�|t]{�q)��8�=kx�k�8���P4j7�Vh��Q<4 �Pw����_N�Nw%C�|;<��#A[���3-��\�{ys��;�('mHJS/i���M'��[�[ �5����u�6�Hإ�O"�w�wFm��U\�+���P�������We�Σ3U��A�����T��/HKrf��LӰ{�<*�e�vt��>�+��*a��#�l�9N��H Z��L؜�%�Y�N�[���	f���:DՕĎ�K�(��9��anJKd��6��b�Y�fý��|$���6k;��
K,�&�=+��|*�Ƽ�Bn�<�eMcI�IWF�:��,�\�d[��&ȸG��A��2!7Tߜ����n,�{h��m������,�|Sٻo�)���0�6�`�^�Z�/j�Gָ�=d%�
u������N���������eH��'j|���}л���q��]���e�.mý�s�z\T��g>�����E8ݼRVSp��rOWCƧ~�������[@?������J�;�p�5b��.��6I���p��4�9f߰I!I�5��o��ZO*���}f�3XL@���V�*�6�]�A략t�=&�^��.���1og=F��9vƌ��6#5W�E��2����y�e�����G:f���n�N�z��!آ>5u3����n�WY��%d�G��O����6���r�;!�C�aѦ笍�m���`�q��
#�VS(e�fN������3Y�b�m_.t�gR�'�A�|"�Ķr'�=;S�]�k-^�eRw������T���i�2`��5��B=�,y!V�B`��{�}	�R|��|�o�l-��'�j��Nl:.�KT]P ��w�/�]���nA��ӻy�=�>z��V��$_w��F�;~�ӝ�5����JM{%�5���H91���N���06���n>���e,�ϒt;�����4�F��91�:]\*WA�T��vzn�����}}�,~��#��ІK��2=n���Y��fvoN������G�QE6gR�B֮dB��]%�i�ҹ��0/<�G�F�z�'�z�[�}zI/�A�#�c r(v��C:S�\b}�[�8����� �������q
��������e*G��}�6x�N�y���7���[,k��r�.�479�N
�Cn�B�����2ȝ���.���>�s�R��`�c��q\4A���y�,E�1M0��U1�-]��xd�3�N�r&���f$[�f��É5�+�.��F-[�V�WX�}�]�әP�lu2_
�yc0�[�����7�_W\��.aы��|���ߜ�짏Ϧ,����q��@����j�30��=`�^��ς��L�y��KB�&U���@�|t� v%�!b��ZL��2��e�^�Ͱ�=���G�H�N4�a��SUN���iHf_l[�ZK�X�����q<�HD\��|+��kõ���7��|uvyV��W��裷��h�ߩ�w���S��H��Q+.fY��~r�d�z�7�	�+cY�ٙ�-�eZ}��REwb�VyrKa���ר:�&�����:+�ٿ: j�hϊ�r�~j>�nO6���H��p1��A�uh�t� �ƞ	mT��>�1e�3�aT��9d�:l��#�^���b�'=�w�j>�˓�]��e6+=;����F�<wVAX��jN��f�d����I�٩�S4T�c�
fy.�!Oq]��k��t���]S��Ns�Jh�n��TxR�#6-Fh�g;�{����{{bt��)��q1�<.�!FDmh|�3ݭ�����uö�a]���+�^N�����݆��O1��5�����<nP�<ewظG�̠e�z�GMR�z�s�l^���t��������ݜOo���I�/lr�2F�\�R|�Pug!��B'W2̕��3��]KV�̊�����j������J�f�>���u�����z��6�]A��°Ś�Rٱ�_�5�F}�����[�ȍqLoK`�F�5J���p�^��	�)�T2��LZ���
�1�v̋�P�NJ
�0��[��{՜�Q�d1p��L�Pj�ޕ9��6����W4�vSX���.��
�����i����V�:cZ�}9E�1��w�x^�:*Pf/C�J�L������>PveV��j�i͗��T	�:Wa�;��r�QdXW\�,0���
�z�ɗHgd��sg�u5M.z��$Ш!�w[ɺ�6%R�S�Ǭ9�x�m�X�Ш1}~����U�r��%+�
��G�sŬ��M��-��4L�ޜ���Y�Ieʂ;�9�w�Z+jgn��2Nj��X�,���]��r��I���[S��,AS�#w��o:��/[��+��֋���u�����#ɘy�)m��R
��Nq,Y�������9�:���&�R{�B2�-�=��\���N]	�&����csT�)�|B�{���K��(uS��+��7��.��[t�M2L8F�e�2����v��)�wO`��T�������â�����QN�@Wک��
 -*�����;��
�K����n�|]�g�g�JS�0^m7�ݪ����&f�i@�[��)��e�۠+��Z���4�qJ1`��L<
�uuRnE[�t�Leʃ��ÀA� w[��6����e�^��w4[��B��4гXާ3#{k�X�:K4B���V��_);ٴ�Y6:��wYg4�.d~�j�s�����r�%9�t�e��Me���(��u湩\eEj�є� /'��Uq�52�s�0�������:���0k�d7\ճ�5��qa��T���j��qj��73��o-�G��ڌ֭��!�Ҏb��bkI�mtbzg;C��Fs������N��t8m��]d^7��΢�:����Vy�����߲����cZyJLŶt߸���a77��B�����a�2o���4�n�u�C�1n^p�D�x�˼\!�v�}���2ŽV��u��b�4�}$�����*��Ų�ħI޺^nl&,=Ԏ^�d�2^0�����h<윂��#��m��.Jb#=Tk6*�E���⢇�;s�Sk:���1�La}��(��jd]\Iaٔu��xf�c0��k ���7|���)����\o�nQ�Ɲ��i�@�^�D(x(8S9��lFC�����ڻ]G�*�ddɲ�v�hQ�ۤ^뵲��T�eIWݷc,+&��zj��d����'>���v��5,�+;i�_A�CIQ9n7k)��R�Cs���2a��WV�I-R�2�Re l2m�9�!�M�z`�[�:�k�m�t]p��t�͑v��R����}��1K%!|x>̲�"01������:L{vP�(�&���C]��Q�S��`�S�6V���\o#r�"vv��Q�y���vnt���m�K��85�vM�[$�y�p��6�B4S1�:O2uƙx��k�=���V���俲�0��L@����9�'�rR��;�Z�Uk;f��h5�;1\X���B�v)��i��B1�!a����i>;�D�Xge�m�R�]�ӓD��Aoo4;�n���vR�|h�%�ոV�NQLڇh�j��֎co��l63g�^k�E�	�P�t���+1���"���3��KA�2+�o\�R���a]��#�x�/\V���G+W�O=Q��ܯ���o�¹��Ѩ��~ȶ�$!�2�����w��N�m���u�o`�2㔞^)���F��L�樕��H>l��,r��E�0�tjef�tq<����ג���Ҙ�Υ˳4��ׇ�ЮN�{�Y�pD��^S�`�٫aM���냱��\2��^R�vK*V�F1e�@�J�NW�sBIV�/U����K�s���P�6��lSz�g�F�*zyiL	:����
2������9|���lGf���R�ܽ@N\6X�/zkɶ��hk೩���r7W`���Y��|�W<�]��5����X�=]k���u�R�{� ���^V�ք�E�T7��`n���n!2��sh�Y�4��j��e&Bwc����J.]ҁjX��ɸ�n[��z�][�8Q�U����0�+��N-<�R�'{&i���\��(����0a�A��k⣽4 �z��w����F_J�1G�v_IG9|�(IL���e�댨3Y:�YAs����J�`隌�՝� �[�H�Y�Mɕ���r� �u�t��4�i&	9l�Tg7z��X
��Sr�6X���W�߂7����z��M��4N�=��i�1���K���n��kz�n��E[��^=�,C4-O���$�}�n ��
��:���vZXQDV
"#0EXTR"*���b�ET@R,�Dm�UX����"�p�UX+�B���"(,Y
��EE"�+
����a��
�b�G�H��`"
"�PE"*�	�X�,�"�*�d�am����*2"�EV,TQV�*�b��#,AŲb؊������b�QT�(#�*p�UQ*Q�F������lZ��
�����Eҕ**�c��hQfDj�1`��$��(-k!cETkUFa(+C�*�\��0 �����R���)PF
-�aq�E"�"�H�֨5v�ØR*.�������ݦ�����:J�9Pl�����Vf+\�j�w�Rj�j�OhY#
k�Qʹ3�{�#ޫ�u��g�2j�4~�7rPWSӶ뮔|K���ۚ�<�����z�`Rv��f��pw6����RS��v�1�-�%̩�H*DՕĎ�K�(��a�b4}a�ݹ��z�;�g�ݫ����R����l�PٖEXRYf�ԧ��]�ԋ]�p?w�DP���v�3��5@J�����9�j�9��^o"�^�,�us̈M�7���M���,��e�QGԇ8��j.�g�mH@��;�p�5b���Tjo��M�cmpܷ3M�xx��'ϗ��S|5�-'�١�}�b>�^�& u��]EPl�]�S5����׻�_!Ģ���-iʥk���7���DR�����pyC��g����Y�n���G9ے7�F7DX@)0�u�>�t�ޭ�bmρV��K��݈=��
	�]f�f��wWK�f�K�g�B2�N�dh�>�l9�@ΘSR;6�.P�:�;Sؽ����~��i���W91�U;b�kښ��߶'=;V'g+����yUf�^Ags�%�w@Q8{2M�Z3���w4Xn(O̥�т�9Ҏ$���
+�x�om̔�G�2�$�
��:)zX[9�Mr��h�Xt�,q���^[@�0v�F�'b�2��J�K���A�u0������Vtc���8u˭��#}�˯&6�8�d3Z-�9X�gr��=ө�RB=Z��0]2�L+6a,���YJ�w~�!���0�XpKr��;���L<�{���wrq��n��qݹM�t��U�"�{C�95��A���Τ� �;��=��\�e5��G?1�[�m��q�̍�&;=:]Z�p�Q���s*�ξ��<#a73z�/d���KՉn���)�������c\�9ltY��������m�+��Nߏ�&�f��9�Ы�I��q��J�c���N�� �����`¢�K�EU1��SI�b6C׹��M$e�(=ላ���A^m��V�U��1�эq^��2fs�e}`Һ�6Tʙ=#J��ʖ�v��Z\*ãY�J:9��nl�Sʭ��X�hWC�g�����EE'�,P�5i�$����י2�w�J3�->�@�KhZ����LLˬ���&��:���c6�^}�n�S��P�w��1eT�ߵ֍e�5�.^H܋�%R�^Ϋ��A���{�q����^}���@��9�*i���t��k^�(��uo3eeIV�b��u���u�ϭpSt���+�z�gQD¢D̗VZ9ٹ��}�Y'VnYi�W$��#�����ʤ=���)�%[g��I�Y/��y��D<}פtd��]2@`�"�_���&���]�{H�\��2��R^lz߀['��FUSܯ+�@Je�G7r4\@fׅ�������ð�SPl}cpmE`u<O��^�+;�z�{yU�$�o�k�6L(���������Un�Ky:���S.y.�� �t�F�p9�a�:�:�	��@h��;T��>�5��.�}�2e��(��9Н ���ꠠb�t+,�Le���(��́��o�d{qVa��j��6�_vzT2��l"�5��w����9�Y�OVo�����Wb�r�8����S(ޝ֚}S�@��,�|#r�����-b���C���o%�/�*������kD(m�<�d��T��vÕK'��;r=�Y87���}aIe�&0��~���֎�����[��|���Vf�=!��]�8��[�>�a�-Uک��ò̌=�����}��w�[E�꧌Z�ES��p^�F"d-ꂴSެ��Xb.�nm�e�t�aVU�E�K���mgM/�vd��ɍh�Ȍ%��u:z��w�2��ᒇ"�V�fs"��햻t+����u�X�N��J�+�\0'�;zH5�|�>�I�g��}|:?o�Sj�~b���jI�*@�z�Y�N�n�%:���NP�r�F��e5��t��/����s�2��z�NX��Aō{��}�N池e����^0T��)�*U1��`>2��o���p�vj �p�W��Hپ��r�7��
���2 t< �tiT���*���~�t|�R�u���k3����#G�]���y���^�}t�{��Ny�&꩷b�!�,\*eb���,�V2�6r����Ԫ3��b�B2�C��f-��k�H�R��J�|:�r��_�M�B�`І��:���Z����IxeH��ۧ�i�a�Ys2Ù����u��V��m�ㄊ�o՗�ӻ°ޫ�4��j)ꀭT�� DF(8ǘ��	o��ޏ�$k�>�ں���n��r��:	�B�V1�WJ��l����Ol���t��0����ˎW"��Xƴi��P΢�,��[-jN��2�g�B��2����:�iP����>�Pi��{�&޴��P�oue�pt�1#/{cz.��+�ys[f��o&J�*�eM�9�TAJ�ή$��[�η��[Qj�Z���1�ZU�g'hD�sw�_����It7�e٤�����[���k\75;����S{�iT���"u�B K3���|���:����⬬n�8���B��h��7�K�'V�Q��ye_���Y6�ܮ��_R�;Jw�멌q�ϱ�[�8Nd?u��zv�zi0�6�dB�y<�1��ӑ�	�v���E�X5�"
cѢ+f^{v{�\�����b��VSYA>^��/x���#��-���"5�|�`��fڦ�ν��ow��'�w
���~�z"�f��@�pU9���L99l51��Zx	��禭t]Vo6��g���x���q\7h�5�SJ���ed^i�,L���ݛG"1��}Y�w�����q\�����LF��@�2�_F�p���k��Yعu��Si�[�Xu�YWy9���LY޶��_�%�<9���el�"�Ie�_R��)jݬ��a;;����1`ƈ�i̠�k*Xw�X�<�X�Q�L7�p�k�hL�B{��OV:�'W��[��RB;�*+�٨�]l��a�Ԅw�Q����qqʮpH��<y���Cw�vI-�l�2�3~���t�Z�rG�k�5����p���{���۹Ms�j3�I�7��s�X����~/�ߝ�in�a�zn=�~�\̸o/	�+�u������C��}t}7�S�e@�7�7�O�59\˙}.��K:ho��\�80���Ծ��S)>72�)�F��W��)�=�ဪ�ћ)락���H_�kb8d���Z��4��ȻcE���EmŁ'�"r���y�lDֆ��gK�fEJ��X���~tE�J�fC���aoV�厸'K#'t�D�yY�y_o_:���&(<����O%�#E��`��@Ο)��Yw��,�2^�6��o�T���X��X4�`�����:L��������}�;6� �̒�5ۜ���%���U �����]�]b��X�G^HU�)���vZt��z�;;�sW��$��4�=h��Υ��x����n_;�ͦ�l���}����z��Q�oB�V)�ׅ)���.>~j�4!���h�*����A�����A��K�Br�����m���M��O��t�Ȱ���l���ݐ�dh>O����R��,�?��!��ū:��[oBw�w;B���Kv�s\W���1�g���C6�����	5+���N��4���|�n"X���NKse�aK���5đ��`�Qf���4�S��Y�S �͢�[������:�0�1�;�e@i^����Մ�D�[����+�~�l�9�=��P�=�P�y�J��.҉�n��ģ���(vg�<���N%�\ڔ��bBa+k�K�J�4Xor��D������������:q7MX�S�ĺJ�f�Q��b�OC��V��o�}β$ExT��Cy���5�>Tt��~��xc��g֗
��]gr���暁ӛ=��L^��z6kqZC���oK��lX�ꬎ�
S��Z��f|�xe�)�.V�u�"i�0��Ӯ/ed,7bn��7uGz&�`�}lN�0c��tڜu�u4����#�|t`kݰ��y��흋�9T�����,1���c"%r.��b���i3r�@�-ǵ�����}�1U���*ԓ�_kܡu">;WU�3[B_�+yd���TX��:��v�F�Օ�xNYs �;��4�K���(*�9T����	��a_H��]��w�s�[{g�}�O7����KF}yj�������C���[� )���N5S��vN�{��YYu��"�r������z�iq����c�4��J�1�����b�7B��[	���{������\r��F,s����c9]f���p|�7(X���p�zU�ٙJ���#Ľv�����Y�4ӵ�a��Z�X��49f���dxw�j����d�"\\�Lj��7dK`>��Gҗ[o�ں�B�/�,U�y��PRP{���ˀ}a|iRrk��`N�`��u8�����<7�2��1Gի��Et��O\q��()�x���F�n�y��7��/:��YyQ}0�K�����s[;F;V'b�+vL���sP��i��a7�=�����wC^�鰡�Z1t"�L�a��ZM�'��LK`;��\���t�:U��q,f��4i�7)�U$NOݸ�E�{��{��q	�{��-Z2��*a^�A\���z���b�����f�j�����,0��}��=�V(]TK���^�5��|a7�Y��^���!�1K��9�����9`'�~J�o�º���i����N͔S��b]!ٴǙ�]&��O3f���u�v���/=n�N C�"�����xA6�*�]�UU���=l��J�!�������o6�����#���5�-E����C�
��<JT����3s�L���OH�'J�ӧ�i�[��u���YKʳ�7��*�}K�	�=*�n�\K�鶍�$��o��H,�K�h�E��q�Y���,oES�H���=�L���y�J��a�o[PS63���P�2~.
�fL۹|!�sgwa�)��/��ɜ}1^�D�̿,w��Zy�z���`�[ϔ���n0�%�K���K�KJ�'��j#WM��J�`�{yʚ�J�jG`��,���:gP=2�����X��8k��e��a�VE��Z�*�S�� G\��H�g.�<�V'��L١�1�vY��.raF{��!��v�&��ns����P V�#v�*fǙ��X��� �'��u"5�����*�a�X��پ����U����p�!b�ck�]�*Q+����p)��L��lt罴��`߹�po��=�aɊ���F�ѦY��^���2a+��2P��U~;����\��;���|<�Uħ��8���E���d2�k�}6ST�^��kB~O�]r����?�'Yu�)� �=��}]�bڠs{��o]���*'�+G�:���jB���	�7 T�ɍ�"�m�1�I�F�Oz�mmy����j�Ƚ[�����
���?9�\�Y�y��Ng��-�p�4 r	���I����8�f��q�)oV{�1�=Vf��EIC":��.�ɭ;�v˽]�de"�3dk��n�nE^�:�S�'��v��i��#A��P�4�х��X���Ur��Ss�[S{��ֺ�~�-*xk�//��+8W�e�8�����|C���2�Y�Mn2�]F�g҅l��=�E�W5*u��{&���|^
V�3g5����JU�"����W�'9j=�z���?����r��gmI����8n�K�-��r�g6^N{]1pw��o�������̲)I��p�����Q.}�`a�>��>��$+�M��)�Y�;6������\�d[��%���5O�����JK#��=�y[����3ԩp�4Ϛ�p:{5Z0fה=�Q��n�����Ԑګ�z�:�4�]Sճ,�W�	���7���40�8��׆k	�-
p�m�2���D'{��!�Ct�� }(�qo����
ס��o�C���H���u��|��V��d�Mt١��_�3�-�Kdj�m�"�H���C��;��l\����Q}��W�}\����F�.�^�/�+آ�k�ȸ�d��a�#C�wc����YۨQ������N�V\R�{��/@�=��5,l��꺸�]���\������8�0�nvmL�{SH9WA�D���<�h���Kz[_npE�&�-u�~HU�� 5uSw��w��)}�� Zܳ�E�u*�T�Ŷ�l=���UH��!@9�܃���N�a�;��
"6g֪�Ƴ����Yhs#�+�6���K�C���q�n���u�cD��ݡޒ���PqN���;\)sH��0��0�δ��Lp�{ٳ��^�{�O�K1��W�]�MX�IQ����[�Du���s�FF�KV�t�aAҵ˵m��Ķ� �}�\�O�E�q��՘��&[�
�� s�L޲ַ�*-kv��%��q�*���d�y���	��z�
��H7zû��GM�3+P�pcһ�WuK�9���h��W��u8y�����4�Y<�l��J�Tu\yA��N���A�i�n��{��Xn��^��Cm�`P��Pc7��7/oxѳ$N���n�Տ�jk�Æ���4)>`�@^��M��9)�l�ʽ�F)���B`P,X���0w3�E��A�w��A�3}<8�r�.%@xW�.^��=3N���7��̌$���[�z���,�Ӷs7fvh�*�]��L[�|����]XM��wI:g�G��4�eC�6u6ߴ��~ǁ15A˩�y�WP���"=���Ka62�u���zuU^�5��Ҍx�""�+t[۲�6��dS�¤�U���X՝|�C��������6*a���:&u��sg�;����s��noT��C�v��H�X�ʾ���T�`��nU�+@�졉C��dN6-nw]���Ef��j�r�F�F�1:dk;a�iW�����X]tlRYWuy�$��3�un���Z����A���ߛ���R�򫝇j��-�G��/��g&MF���!�b���K��Hx�T*cZJ:�WH��O,ַ��a�(���E�#�Yu�c�F��eN��O0�P�n�?��8��0� �v@�#��k��=p�U��,C4��z��S	5�q�����z9�=�3�{�4���%�V�ȁ� �n�(]�S�Wfnh��K��^큜�	�IT���f)�y�`
�X����M�����ܢ�����\�=�bBR��v=�B�^��l��|��A�G�7�ա�r�盃d�e�U�a��R�&7E��h�p膬	L��f�zy�$A��sg+�����+���_��uTzuD'I��-���,�H����̫�ڧ��gF̬�R{7{O��N \f�M���V;ܭZ㣌ZYj{��j�J��;Fin顠�%�i�$����fQZ�(R�Ν�X�:���l�j�5�+Z�����r�L�^��u��/�>�h����Gh^~x��eC+<a	�`lj�f
���}�Ìⷴ��W��ɼM��nS��a�-���W��v9�W*�me:�Z�����.��6�ř��}��.b��	N����L�ݗ�O�l����^m�z9=�U���Ś;~L'� U�M����ӏWo��4W�W��R#�S�τ�}���g���k�M�{���,�'w&��%�W����6�J�8�D쫲�O��}gȫ�Rڋ%eb�U~j��X�%j���͎-�Z���*��b�DX+X"�(UX�,Q0�m��b��ET��R�F"���.FE�1r�QAV",X,�X�Ͳ#	��QI�PTY*�UPP\1AF�nR��ȪL��B���ܰ�, ڕ���1d��U����VDAk#J+b+Vֲ�խ�UQd�ڱj�EdE�\8X��T��ȹaR�UA�TQDf��(�D�"�Qb֢$U$Z«�e���PPcp�"�kB�*
�E�
�W6��"�0�DZ�-�j&.0*��6��b���ֱX���Tj�%-P��-(��+!R(
6֪5�V)*V
ڈ�m��jD�[h��m���m�p�Z,U����ۊQV(،F��X��c�.���9�I�M�B��ⴴR�3:�q�t��m:��d�q�r
/z���:6_gۨ�;-�a���R]\ؖ3l7���T�2։�s]?�ګ�G�r�������^Y���V�Z>���ZI�=K;k�6�����c�<�dh0�91�@��p�Q���̓�+����}�غ������A��7����l�F��g6X�r,�PܿVoK���YC/
g��mov�\�jC&7S��p!�Y8�yL8R�)1�+��>���6�B��\D���b�zzI0�&��ԒѷO���k(��ł����K��&<+�R��{���i�TV7���Z�tˀ�7��Y�r�EW"�Uq�ʤN�r���P�%��M���P��rJjpB�c�!5�;��`�)�6�����>,_dE�9z�fw�:�;�;�4	2(�w:"��*�X+y#�q��iuY��t��=Xdx��':ږƪ���gAE����q��q������wLv�*�����2L[ly�vx��k��xzc*�ƺ���P%R�`�r4\n�1+.f\t�Xq��eY}��n����sv5i��R���7ݶ��:�׶�T��.s���nV�^� �m����� �۫K����O�s������l0wE�`Nf��}yZ2������un���R��G�牻|2HJJ��ӡ:���qk�ۺ�<�-��Xo�	��B��S^��n��U�:���EV� ��p��âLJ��q=�����G��s��n媖7�����U�����ސiv1z�@��kx[��o��u�X�����Bn�f���&3��ٸ�B�`5(�˞�XQ�����oes�b3�����]ݫ]�d
ۑ��i��[W�r��^��{C�E�����/�7(_³�W����tw��J5�1�-�ӹ��3���ލ�����I�1lr��U�z�"��в/�*��d�K��������~�>��������ǅ�i�po���6�f3��wqz����N��������7l¾�og#\S��3��C:os�κ_cP��V�O�Y!�[F�[�ML��P�LFJ
�����2�1�s(��]�G�Bn{���&tVV^&4z��x�C���W�~�5��R��{X����69{/;�U�E>|,��k�P�� gv��nX�A�Rϕ*���0]/)�x��[n�e�^�!�����C�V�u��]��C@�%�Yc�ڨ�<�	y�����r>7��&�.mH��w�0���j*�.Iٌ}*if�p�;Q���⣷�/�ښ�ȍ�F�5�*�Y� �N�M;�vH�G6�y�Noe��ut�;�j�b��;��ofk� j�&f������hS�l]:ޒ�, �AdX�s C�	��U0����J�/̐�{�U��m�.'kF1(�0�����lE�y��GI�m�X��.L_l�V�-s�}��A~5��q��ެ�:����P��ȷp�LS1lv�4���V'w�<]�H�R�'Z0P��9ڋ�*�tc���.ظJ�C�~n��5��)9���r�{�E�FxLd�����h�p�m�J��0X�>���@V�p�}�w���w���R���l�-��
�3�(��]�C7+��0[5U^,�P{
�ƨ'[�����wӫ��tY���x��M�9^ztŃh���FT���V�e�OxW�^.�b�n�qI�w��R��Q�*\ ���nenS=�q�E�>�/з4вՍ�.�F�U��x���]T��=6��.�tK�;A�"����b��*f�b�;�ag_�'�A��3THg�]��f?t�"����+)�*-U��C _�x.SPr52�tBs�*��|;��ˬ��ؚt�/AIj�pzKF�X|n"�N����ɈY��uoC]�iF���w�˩vW�U����5X���P��eN�tk�T�R&w;&*�+���:��yM�GI��Y��l��Vr�1,�7��90v�Y��˻?nM����۰�a��u��z���h{�=�Қ�02���b��N�Q�n��Oj3����o�L��ojW�=�L��P��EIѐ��s�]\-˼���U9��*aɌ�m���֚[��V��C���qOz��1�"�������䠮�>F��v�u���a�K��>T����@���^{_�^��9I�q\��9����`�s*G	B�F�b?MΓʅ�qO߳�����i�Yy�r���L\A޶��F!��u���.`Yn�H[��of�n`ݴ1��H.*8)U=
����N��;5b0;��,S�f�u��2a����\fΛ�^J^d�hvh{s�M�����TT֓�Ѓ٪�3n��y�E[-x{�r��	wk�p��sQQ���W�(O|ߜ�b�`�CdX��0v��f���:�˚&v�zG�A�T�b���=�i�k��������ZtrS�G�c2%��K��*��U,3*�)솪Fk�,0eP7^?	�,>���1��Df����U���e�7��F'sRd�������N�,��NV��)N:WCe�P�r���;�e�5�H��y�9�9N��"�+W�;A���r�p���h���P�Xp���L��,���q�-HhfCRQxV�0#M<模����r1ׯ;�;G�W»>����Q5��\K%�#E��ls�03��Y� 낻3nN�'���.r�S>kZ��W;C` ���Kg!�{��lmz(tcy�խ�/j[˟?�=<^����,�Mxc�v%�-���ح�op�?s~2\��v��(�M�z���э]M��������V�:����v�\��M�1���'v3u�TO�.����d�@]%u�{zL~Y���@hC/�bnu��_VQ�W���gRj�CW��k�ޝ�G�$铢�[4�X0�\`>m[��ylwc9���y�u�ti�Q�j�VxΔkmp>���5[�7�̳+e��['��D�kg5�{8�X�.�0������*N*!���W鏽8[E�3�!\���t+$�%)����*X�&5�p�\V-��d�-򞢞(���ư:������/��*�4���Ŕ*���#j�*��s�vb���w�ޥ�gslA�����2�N���E1�UK��:�JJ�Pq�ߥu�y�x͂@��yYwUr����(X���nlҘح�ۮ�4˾}F/C8\<�p���{��Cy3��طWn�eMR���k�Y.����&u:nS���m��zeN�ҫ�����w�v7:��zt��o0�3��'�����v��(�E�Z���"c�"�S}2}N��Ȩ�2�ҙb�V�K����X�;�u�|�����������`p�lI�g��mN:ҩ�j��xof.���Ze���v������f���5a�a�~�HD\��r�vI��1��~��ۡ����n{���0�YǓ��*ԓ���k��$'�*W����z��3'�����,��*��l��$��W��[�׵�K�Q~ə���5؂��p�#��U���z=< �W�޾�XH�6#Lɔ�:rK�^8b�W��3v�>�Z&�U�;���F��z�'X�g/��~���~�Ei�7�vl�fͺ��,A��퐣6�73gwr���|�3�иQ��43ˌ��n7g"�Ző`�ޓ[��F���1V��/.���j�*w9��E�{�LЛ�s��g���`�>�-����Cy{�`�Kf3�]�G+����f8�ި�g�>�r��+�ӷ���;Y�=����f�EO��1E��X��Yo1��;�6a�rΝ8ZJ��v��a�ڻ�IVM>{�y�u��x��YJ�𗛶�%�hמwR',���}������+c��Dx	Z�hβr����d�&k�u��������^�˂s9)��.�F��j�Nʈ���vR���>��B�0~ŏ����xc���a�&��"�N8�3e9cF�wG7"(���y�.���x����bg�~�<`G��BE�*�����}2�B2\p< �`�}��f	�Q1�ݐŪ�S*�R���;�`��	u�PV]b�^��`��Տ����A�ϖF�V�;�}�E?
�RʥJ�Z�`��0��ƅ���\yr{�1:SFn�z�k�ŭE�ȷ|�2"X
�Ȱ.
��a�&*Hgp�r���)��<����Mn��������79�+��Z��E<�@�2$
��zd�8�T�*o�
H=��W__^uk�����Y�u� ]�qʡq��̻�b2ީ���K�{��n�_�0WBi�[��+��1�X��׎��uyh�͔�J�C�����:���«6&���$�ec$�fR�H��[�������E��0�y�
��z����ߩ;")H�Z ��F[yf#Rf(�2�ؤ3j�#`��/�+��W�k/%�к�i�y���8K�傂N��m��t�`;�.�̖s):��Z���AlG`��β^`�	�Z'�:W�7uI�
�g\� ���Ó3.;o�pI�ef����Q�ޫX��컾��Op����i�p ����C8A�o��Lݜ
�fJ�����Ρc����S���j�C�ۋ`ˆ��>�DLܪO²�ZOH޳���s��R��X�<1��)W��w	A�ܮ.�}\(Z��BϚ��K�4l�26zj��mk�� �ӹ�㤠rtB��͍�c8�%������i¸�-�wW�s�[�;��'��%<C�Q�=����\�x �����9�4�s�=�:�uJ�sp�����Ɯ:��0o��q�
�Қ�]d�n@�b��N�)t�P?.3Ӓ��fI0��{j��-�q �7J9�A��M�.}�-T�,ߛ�.�Y��l�W�.k��^������T�f�C�iᚢ��s�5���^+���J
��jaߝ�\j�o>�r��#���P���͌��i�9��8��,������i��XBҸp��Q���{({�5Μ����z�4���(g�>��V>[�)\��0��Y9�+T�ys-���V�w-�4F���#��>��b+�¡ߦ5� ������,u�*�9���}�#�#�Z�?n�fp���	�/r2���W��Ôz�
Vf�����-nfوjo8�&����Q��^{�;��j�CC��F���To��BFn��:��j�>�ַ0E���_eA4��vQ[%�-�9iq��"U�wz�W.�E�%�j�\j	y��x��O}�vY�2$!=M���T�xk������ڐ��uCoT+CV2�\s+s}�2�:�+Łi��ER�u'��O��	����׍�k�Ť���ª�,G�%�:��.nrNy�jV��^	����Pk��e����ϸ��o�C��~33(�����:k��*�"�O�N���X�2��/i���^�,0b%P3����XY�n��ۚ�i��v}���,��[�_�w)ue^s�`,�6Z�7ϰ����_�>$n�;Ooi�鷷W\zi��+.��n�cF�qQ5Qs'�V���M:�߰E��t�^��6�5�gk:]�Uf�A�9�5;�b_ش8F]P��I	�btrގr�^�'���r\Bt���h0�o�l[�-�6��g�� �6��ci	Yƹ�bثjO�i܄32���3��yd.�U�q�m4|�/�&�����j)�R�by��ut\���R��;��og��7T3�'�LvD�uj���=�V�f;*eN��JlJ�9Y���ep��S5w�я���7���Q��Wm�Y�t1��fҭ��rbۜ(��9�6ΫX��z����.�l��
��*pO���0�8�7����.J!w&��T�-5�8�[J���5rb�I�SCentA�̙:5+>�8O����)�A�v�r5�{4�,k��9l:,���:,�ܓ���J�1���I�Dg}A#��!Q��Ю�pH_�x5,r��h��qX:��s��]���u�R�"���Q�AF)����4ڻ�U�i��ز�T溛N?tLR/�7r��ڪ���l��v�oD�^2f��2�N���E1���1U���]gr���3,��I���ꏋ��=O����[�YL����靧MOdEE1�T��vTtp�+�koq���U���kDW!j��j�&� p0���#��f�|�M7���E��u���S��9/��E�����y͐�%�:�Q"���}un�R��M���?{�fЦ�n�"�L0��ʵ$�|�����ں��n�����M�1�NRһ�U�&f��X~0vFoN��[�U{��'[���Sd���W)`�]�6�K���m�	���������Aj�?�zA����������r�mG���e�5�/`G!*�)��zy=��e�oX&��v�j�������<
�m�n�! ��rV.d����3��0�hRW9P�͓�Mu�Ⱥ��2�l�+`T'sk��ݼ�#[ݻ�.$���K�FWv��V���F���k�xNfg ��<�S��v�Wuq�L������l=K]=\�7n��Fey�y�W�E�[9�#A�E��U���V�=^oafF�\<0�	��F1	��s �C�����m_vz�#ʙ���:���fd��/0�	Z��N��*�;�U�w�h�<��:�\�r
����f� ������o\���Z>OA�{"B�bu�F�W��!������P�O^s9�g+޼v�b���K�n�n�؉t�8Gݝ#;	%Y��Ys/t}3N��s��O'9�>�.��n.��<�� 6,8p+�F75��lֲ]D�9j�htew`eM�P�en�����:7n�VēM��C����Yނ�S�:���b�Fdx�
�fDo2�͡��6=��]$I�M���#�̱�L9�I7
W�����G����ww-�d�YZ,ص�a�h���V���r]L�w�x�6o.=���8wP�<C��{/Xb���:��2b\`a�g��OX�BZ�7L|��wTe��sg���h�Q�s�['"��G�(v>GGh}̽��NMs�J���Բ�Nf��KF*�����3�_�f��Sh+f���.�q��6v|��=�^B�����x�˵i�]=Ye�LpR�!+*��(9�ڽo0�&A[},"��"��ܢ��r���wX����MA=�r����F�z<�́�#־�X�g�Y[��r�2���z�e"@��wR���u�X��+�b�c8��A�T
����VKS6�Vi2�����\�%�R sj��4M.ќ����:S�6\�])��lT�x�΃DTZ�d/�,;!��/u3]��h.����a��/�y0�}"՜5WJ6�uG�j�F�.���$d�޹c�3�V�k^M��v�"��+�n��W�hL��q���z.�R�޺R�{�|� d�B��}���U���*!8�p�N���[�����R�Ib�z�Џl\{�U�̭�t��.��ڹ�-�(�fIA�͜ϭ����ɐ��v�Rȝ��(;5��t��{{�vOMp�٢�t)!���@�툤	�WV]q� �>ۖƺv
@� F�J����ť�s���H�o>�R�8���o.�d��uI�w�VJ&��i���KQc�KJ��W�}@���V(s�3J�k$�:79��pU�Y���:�凌�#yp���=�����3o��,y;��wMU-~J��+��p>������j6!)+��hknѝ�DƋ��j�I����ohPE;wJR����,0�&\�,U�nP�>�h��֚��NhzX�vrO;�[
a$�껌b�2�MKfʙ��fR�mt�L�; �> Q5@ EQ}R�ja�L-���e-Yi�,*)*
VT�6ֈQ[E(���
%���)qF�m�cJ��D*Rҫ"�k
�i+���1I�Ve�p��Re�EűU��d�)���EX��V�E
Ռ"5%aZ*�V�ԣ-�m)[*m+�C	0�
���1Q����QAe�P±pȰ�2��Im*(T�[C)q,��PX����Zص�`��P\6�kaR��(�m�KQ�-���D�0b��RڣV�L��-��KDk���sp��bUj�6�VƱfZ���%��jV�6��F���c)KJ5ikQm�D�sJņ����0�Ԡ��D��T�����IX6��E0�ҋ1l��*)U��U}�־���{����K��q�
�{����|zJ�/a�Y"�2�nw9r������	��xe�r�t��ԝ�VM��^v��ՋH@�,��9	�����a�3�b�|���т��x_�1+>�W_�w����<��iA��^��9�ǚ�̝�7\9��X�>ޓa��}L�m�C�Cu�ܳ9�d�U����'��u;��,9����WX3%C{|��Rb���YC=EV����q�����)�ԕ���P��>=T��UWF�1N��1���c�|��^���u��ׅ��3���+hnjX����X}Lpg�BO�y�-�[�og\K�y,U�g����N!�r����6$��芃}OկBC��*�o
������Y3g������k��M��U���ǃ�T&P�JC�T���eSV���/<�������Ir�����ݫ�"�)-�Y]F5���o�����J��|�T���f�l����V��\�:��|qh�f�>O5�mj,^[�S�, �AdXu��Ah�S8�@Vےf��΅��6\GpU����H���+���^Ms�q���<�@�2$�!��Q3���@j�4���"ԫ�Bv�p�d]vE���QB6^��6�����؆ϝ!3
��w�z�g��=G�����:�\-|};�,��FN��8s��s~� ۝�ţ��p���n"��F�){a�I$4t�?gS�[�V���S'�6�V#t+F+�Գ�Vm*u� ]��a\��p�b�պ*/��Oc�YϧE�sUXj��d���&���q�%:,`�k�U:ȵy]q�ް߇�M����5XhڞZ��p�{��# }ʾ�5�&x,���QK$�K5�e���f�E��u��^l����3o��iv����5OH�. :�Dco,ÄjL�࢖K�(؈�c�P�vQ��hol�Ǫ�곕-��^?m(+ۉ�!��U"=:b��kF�yPΣ�B�U:v���hvER/'�*M��d�}�r�&
����su�qϼ�F��\ssm<�o]�+o��\��fd-�w(e�%����<Up��u�TrLȼ7OT�|�U�;Z�dx�/oN1<	=Yx��C�ֳJ�5��O�_- <<#��'Y>���G����7砜i�;���RZ7��^(��
A�β=�{�ۊ�}�=� ��z���)��Uo�4��=r�\s��kj2#Z�ʷ��7U�mEpތ�����:���긼M{���	^�w�m�����)��K
	�*���p��ת��p�ڬ�y��Cg"��v%b�wRm�iWݷ�6�Dt�*�&�xu<#e���Ld�����Pwcr������T
�\���2��J�13j�ý�w!z�j��O�Kԧ�ц�;��|#���A�k�ղ���x�o�f��Ep�L�G�u��G���Ɲ�~I>�[��ݯ[2�a��Bu���=����'^?��9G(��J���WozaHv�&&0e�v�:��H���k��1�o��Qn�,��qZ�*�Kh	N��J�t������z�M&����Ƽ���;6��kx�m�<�p���	�	�yA=B�Swꜫk��7Ck��M���*^�P|֓��=��e�N��j��x1+[�t�d�:^9\�p�,GK�������Y�-L�:C/b߆�ZL�40�o�Xf�f��=��R��h�a1��������F�@}(�qp��[9i�㞻cAT`�SZ`nn{�
�b�TȈ��Ł'���߇P�CU#�,0}*��q�8ԫ<�$��Z�h��T&�J�\�����uyd�ğc�:()
xel�h�����S�������r�Dp�)���+c�(e�f�V�3gDTk���(�����Q�I�m�}Lh�h�@ls��9���o�3W���k��Ȭ!^U*�G�R�q:틗e���Kon��[��J{�����ʮ[̸���ݜS�`���{hJO�ͭ׮󐕎.*i�W|�V�u1L��w�jv�X���ωKէ)j뺓�ΛS�f�h�߯�aڰ��#��+�T �/�u��X�-vf��Lgf���)0��|�o�l[�/�H��n��=d(3i�*4P��*o�':���,���\󩦼�<�uyd.�U��c����s�j����7�a�[���i[v��QKr�u���A�*w,�q��O'S�c�!���b�&;"t�QJ��׆�3���V��b����O�ʳ��c���s`�v�r5�{4�e�s��ۃ�z�y57;���!=��p��m!\�)�ns��rR�/m��,r�q<0E�(��3{��pJ|��t؎�_���|�A�yM0��U1�֮�1Uf�f�B|�n��;�)�
~3�lά��=�{+�m���a#G\W��0�2�t�lvz���4�Y��\��:n sÝ�꩑�{V7�j�[��B��b�-�,���Q�yСI�k����{j�݁d���N-0y�d���u���__�����"ϭZ�$I E_&xmN:�L׼�k�վ�P�u�ܒL��î�B٤k��T��Y�f8�n�#��>�]wt��Q7�2�гƴ�-G.��mHw��n㎘ ��Qj�����*�6&1���sP� ]�U�슯�����A���{���j���d4�N\O�zP�m)՜�M>��'~Ld]�t��0n�f����sd8Ȗ�Hb�OFߝfr}���#>�Y#E#~��<��p=E��_Wc�ڪ�>�v�%R�a�������d����>l���ŷw�=�Q��ܺCn �0�wF9ڪ^�Q5�W�G7��CQ�礩R8�8l�}[���xM�L���*�x��B�/Á�7�]�Y�-Ox��9N���j���N
�`=pN�1�+�>��O}�mނ:�w�^�� k/���k=!>�Y�S.{O���R�^xǶ{@Cf�d{����>kE��zL[t3��H�݉}pe̱E��U�ݼ���GX������d2�b���W��uZ`�̋�3��yz��1g���]�ZڜHXq{��K>f��R������UѸ�����R�n<,{q����3�M�x��Nor5��״:l95�R�����8$'�'��م�ҭ��aPP��IU�Ü�ԭ7;�쾖4if��Uw���Rc�4�����֧��*���*�*��Wϻ��{N�����8�#R*���ǢPy���[vr\"�5�Xv윹��+���)y,�L���p���e̫��x'�������D�6���N[Y�umweD_F�́��]��d�^-!���������v㓄G��XnAa����z��ս�]ru\����D�lUu��˼k$�;�U	�8��Y)&��L�.�.���ʽ�M!F��Ǖ�����r|�2�˨�]���k�!@��:����\�Y;��go�+��a�'+�<�c��y��-�+��S�� B�Y��"'�s]��KQ1�ևsn��Pt�xf�DкޔOR� �l�Kmd�Z�0�E�.k��F��)z������b@~�w*d���D1��:�t��0{ye#W��y�:����Qw��Z�B埤��#�§g��]:��$���%/˅,�Jf�rk�d:��1����R%����m6nh�������4�)wu0Ld�~��<8c��V^+���ϲ��y.��8]�W�`**|@u]�AN�DF:���{�pװJSך�7��"K]b�K�x�c�ss�ٱa���$pbk�J����!N�%����Ph�p�u���
+իw������$4����i�\��ʃ��Á�*��Km��w4_�W
�>�U����,�����o۵{DX�Y�齶���ި=Ż�Cs7h�f�{+��͝�	O
K�����.�����o8ʷ���xq�GDL��u�X]����΋F_d9U�%��{V���Y8�
ӷ��R2�`9[�e����y�L�;cn�����dW^H��YTφ;ۺugu?�U�{��]Q�a/��t��ޮ�N˙4dxOw�vKgC�z����T���`@ϭ敍@��p��°p��:�X�Z�@b���󛚀�J�.������g�c�D��Y���w{A�k�u�W)�|���0dy�0��)CS�x�2�!�o�h!���s=~�T�}�<�UL����S���4י'ӧW���ң2ʭLF[�F�/�J�b�g+��9�\���0}���.�P�,�D�':p�4����P��;�	���_��u�������[�K�c.��Qʇʴ�5�U:��D��{�u�K�7D�>Õ����<�R��	e�X�ц�dt�9��c��",��n`4�T�$xM6��I���������VR0y�륻W�L^�熷[��F����cϼ9��,4>و���Ƹ��-���]Z�"kF �괁����M���g,;���Q�
�VJ�,�N�&O��Q�C/)̠X��M��x8W*{e:)�������52`�smu�Q���&}����kOy%�|5Е���:>�5�H�a*#�9بMML9���T�]�+[�iT��S/���B0W�]�j���ild�p��7֘�F���]���"*ށ���e���v��(��C ��h��p'��t��F0:�x>Ӕ�z�sn<f^��+����##C���3�����?C���{H�y���E�J�!��+��؞��-�������y��eu��X�Od?w�c��9� �A�����cv�]�2ېg;竹V/v��������5#�V\��[xw/�p�`��.L��׌h���ڷ��KMI[;2��^zt�0�ݻ�^ʤ�~�`���t�"X��
�C�@jWv������h�j��/�p�>{��N�II��T[ܽ��R������,�(6�z�k�j��d�WN\�<U@��p�[�ov�ep���#����YyA��VX�w�㼴j�פ�s�v;�P��*A/Զٝ��[�#|ڶ;"�7q��[�&9{=�����N�N�%*���j��\#�r�lr�+.�[h�og=�+٧͖4g���'HZK���fy�~��P�½[�=]�Ô0m�_rjp?w����B����x�,���>��e]� ��)��^��M�Ca���e�cfw>�Ƙ<��D���yO��^�E�g<ÞZ����[ǻ�V5�q
�v+�{0����&m��u+/:�:0�t����˝��E��R��Rw��\�F������`6u����ɓ��`�"��c��`£r�L̡���b]%\)U��ł������7Ǟrz�R6/`��\�3��9uq^�f�^��2��b�o�JZ�a>��}�^�KoTi��kRޫ*����yn�eg��P A���f\�;������z���gy�$b'kt����([�a�Z���Z�	�H����g���xV�>��I
Hwi���iu�TT_T�߱��X:E��v��on]� ��@�Y<S�svE��|¿T��1O(�u�cj	���Qp�y*���e&��ٰo*��@W��ħ�L��eU�y�M'+�]��"�mo���(5fE�~(n��W�7mY��7�q�H�[UM����92tVU���[A�oP�/>����^*�����$��Go�#7�����M^	b�Q��Z�za����ksf��Fi��k���f��^&{$��[�Wfy�
�؛R����x��<r��C���ua�쩏+gPݛv˅�y�m讑G��䗤P1���l��r[��nVJ�Bwg�Ƀc�z���׏	�SLM��u:�ݦ�c8z�E�4w�C�N�I �=T��)�y%:ɾ)�$-b{��5�� �Q�n��o_w*����Ww���M�wҟd�u�D�'�&�㖡l���q{#��s�C��ܶ����\��X�k�����s���nbZ7~�B��ޭ�95�y�U�{z��{�i�dG�4�x#=�r�� �5�;W۝ﶮD�E�w�+xǖ����6��m��� g��>��H��U�{&on�ދ7�q�īת���-�.:�:�m�9-,T����n�r��ǻT5݅���N�5]-sm��"�Eu�۱Q[�e;���4F�~���*�:��ˁ���Dn7t�>��i��)P���E�� �y�E�8o��a�X��z32{6�/�Ҙ$�R�n�\�V+s�Q̇\���Sv>c���YKu0v
�~�k�E]����+֎mye�K�w)��V���!�$9�j���ј���X���-ŕ�K�v��u�;���Te�}�1�#��^vR���>��;q������7EN�t����@e[S� jμ.��*z��n�(��ω��4;0�'4c�	�y{�f[�L�u�}���m9Q�x�n�X�i=Z�����j�qTp̓j����-���4��B��F�9��1u���fIgqxz�Qu	͍��uw���ѹ>�V3T��Z���ɝ�o7��q=���m0+��F67���:H�tS��H�l�F�(�-QI�7A�����[��7�����Fu^���\JA?�(B5����m�-��Ւ� ��Fp2����sJ#u�f����l��Vc면�D|���Yl��׎�ʹl���!Q�̣�rbO�N}VB6��T`ͷ���No������J����G�9X]�=�eȩvw�g��0���8��3���|r�M��[05�bKa�l�.��WD��w��nb5v�,='2�q�-91m pN���7�.��s[-]��_-=�r�ZCx�@��y���+7*�����������8#��t�⫐�w}�
�ǣIU��
J�-[\�P``���}���]��Z-�n�w�D��7@
;��LU�Z�E�ޕ�Oo^��)\�-`���T���!��lυ\7yF�&,Ys����te�+�̗����:�Q��ox�Y~|���g=0ݜ�@F�(Z�X��4l�r�i@�o6R���՝r}uĎ�l���s*���e�YaN�N	9Z�~gw���+�T�4*���wٛ��U���S�ݕ������-|�V��1l����l��Wa��l���m`��A�� ��j�Y	��5.��<+xH��W��Z�fvr��e��e��Qݼ�����=]�Y�"���lW,�c��=�K�23zi^��U+x�>X~��N\����ّ�񀩺��%���Z"Vڠ%���}z��v%�[�dl�x)�!�+��(�OV��T�}2�M�L!�ޠ�~!b�1�y�T^�)ye�ի4�2w]is��}��8�K[ևwG���t��qr%�.-��+�zbL1�2{H(Lm�Cue"-�h#i���۫�k�(Җ�N�6�:D6�o	�v
T�LӷҬ�m-��@�O�1�4�u�KW�J��4�᧫��JP�35^Զkr�K�[K%���F3�Gn_���Wu��]Kϫ��=�Gn��F�T�n�A:j�Z�EWb�<WaӖػcC(G�d��[��ںv�$Kȫpv���f���á�E�-�!nZ���>��@���ۏoz��y��X{!tc\r�GvI`]��q;�*�sv !qVG�i?]�J[��6�æ�G�E3BZM�L�Dڝ�4��N��gJ��-���]��K�w�%Q�ZԬD���Q��D��B��0�AC	������J��[EbԭT�E
�[[1K�,�
 ���-�P������-h��jUIm*D��-�e�B�me��c%��Z+�)�U�*���
1Fg82�5W6S��FՋn)�
�J"
�sh(�*Ƞ���"-s��	���p�Җ�jkWQB�
kD
6�5R�AV(��[\�
⥵��*����	0�h�kYF-���KB��[h�J�j2ڊV���F�-��3J*,p�mb�[TTQb�ZU��ʍ[q��X��PA�E(�V\�[s��p"j�**�ʥF�R֪��A��QU���)ijզnZ(��jؖ(��6��b��.��|�f�M��t }Y���WՈ{�k�6���\A���[����\�[M�pP嬛�\�q���s����'�l����5��zMtcrİ�8ܷ�f)eA�K��EGpS)�)�ʎ/�o&k�D�m���������,Е�!^�Mo�����/M��wEͣ�M^hx�LFsq~�A�heC�4�̡r{Վm��Q(���Nz�T�����Ayj���Lt%�A�{��jP��w{�ՑUW�N����Ƣ����S��x�ܐn� �̞��N�pۈջp��0�:j��@vrM)�����)�ڛO�2"7������ծE�^s�[��E�����W�͂�1��w��I�a,w	��j�!�URE[)��=��/uU�%7|UR�ݳ�'
�kkC&?F�
�����\t����mbP�SjT�CQB�����I�s��ii��W�Q|oǺ��O�~��z��v�|u��.���S��pa}��Eԟ���CuQR��Zr&�g\gU��P���+�W�,��Ԭ[�wI����3u��N�;��2����+�����>��y@�;���C%��Q&l��rt���N����J���h|e�d_^5˄����Eb�^�H���w�G�;�ܢx{�/L��N�3���O���u�s�R���by�>[�ǆ�˱ۯ�at!�6}�8����6>��M�ʉ�}���P亂繪1Mq-�+�D"49Zz&TE���	|��VZ�#�[>�~��䏪��=����&�rK�7��]j�Z�+�tY;K_Z��A��ʈ���{���p���ߠ+���{!ǀ_g_0�B�*�[�>�9e�+&q<޵	�m�n�˕��}3��n4�^o-7dnG[��6)m�%��J�u�q� F������CJd� ������څ"i�ի�J[�Ob�j�z$��L�:�Qu�E�x�tO*�ե�*��u^#1��S������n�[����݋�Fۃ.-�y�.c��7�p�緳[RVG���S<��F?,0���ǋ%j~�m���<J:⾺$
�ٜ-��2�f.��1����Z)Z�����7`�h�Vz�N�yiR���e������Ng�j]�<����o�u����N�=D�.Y4�k��,LR�4���,jv��p:3�]q�E�(��QʍƦ�'�����m���q#{�ۄr{��,��qwC���\��b��ޮ����o0�u���PSQx��Y��)C��Fy�z�9�k����
��cOLC���6w�S�s���kFq�����ۜ>��_;�O�ރ�"���|��X6����sZ,��8�4�\g_�.��轞�13�.{"_Q\�h(����cU��7-ڹ�Z����|�\.�4�{t�����(��<�p��\�A�j������W�:4���j���h�K\��+f��a����:{���9��`$t+��떣R����~l�2�m�_Of�`��Ub�U�(�ex�1Z	�Xw�)To;p[z��7��{T��-i>i����@ʯw	��_E�9Q||F'��j�At�u���=uZ/�݂k�/3Q�v�{p�^�Nw:Ӿ� A�@|��γ̽�w���¾:R+H���2ڕ{��M%h\��͙��7fߩa���ŶU��p<ی�5j�Qe�5��9}��I�+泻��6��ha��!tM��]-v��ܜ��(�� a����څ`=�n[�
�Y/�l��0��:3��v�o6l�8�[#|�ʆ��4Adtq�C�R9��GU��zj��=Vr�^>���@�)�rǠ�C��D5�.���q��v-������ϗ��`����W���=��jxo%�}������w���\���˙$�������y/��Rʼ���S����=�Gvs�OT�k�\�3G^�����4�7��͓��j.;ʹUF&���M���Y�)���]�_�|���͑�#kzOt�1Z��Ag?u�\� ��SQ�(������Kot�YHR���mª�1F6��7�-���ٜ�s���m�T�+���ahy�5�7oaM�P}җ�YC�J�s��qw=ֶf7-�s�Ī/W'���.>���<�
$F�������]^p=noD���`�=����/�z�.��k.5NV�x�q���՛��%o�.�w�����n{|o"�*
��a&�8*-���۵}H�S��hnYê�w7FV��Z�2B��`/���]��/b��ܳ+���5�P��v�q:��+\�7�L7����gX��d�;����b�tu�KD#�|^��ysν���-F�_.�s�T��@j�w1�5������\BdEE�8L�!�z�f&wbo*8un��ʳ]���&��\�D��.⡻*�< ��E�9aS|���B鹅�P����W�r:tOVT�Y���^��r�m�Y5�Y�����
k]��N1mAY3^-�F�Qi��ٷ
Ÿ�����A����r�/2u$*��Sʋ�W2�*1@��n.9c��;�t��˨�Æ�ż�� �/�AW�#����٥��5Ɣ�%�G^HJm�tvF9�q(O�I��v�����j[����!ՙ�)�3�ÝZi3a�p�Sjk�X� V�0��n�5�tլ�A��1H�^�E����X�� �#�\����.<c,Yu;o�T�b�3VjmB�y�X��G2jl�L�w�r�ɽ1hk�f�5��(��50(.�3��r�`eG�V�(��R��D�j�:���S�L�1n,2龖�+c:��S/b,r��fN�+���4�<�X�N-Ѵ�����w/�ˏ6zt���-Q˅�$�6p�{ݯ�]�`�R0�b�rU�Ɇ��dC/t�5�V�q�ٵ1��T$���WL�:�k�57X�F'�X��p�ʹ꾕�C��g(v[��/����	ꗨa��}W����ھ�_^�x���}�;p�כּ��Xr���w,A��z�ڕ:R�+*/�������QΣľ�Z��-o.JP)m8�1�*�!���^�YQʯY���.��eAAY�ٸ�_U��:�^%Gԟ�.�DW����*�B�c�Z�u-=�c�n4��,�J;	�l�2c��[#+��pim����c=�y�1��4uz�f<[�go�p�Щ0���{Փ�{�c�*Ԓ,aq7�l����|VL�'[֢�"ᱍ=Zh>�m,�:����=� ��]3/-���7ܔ��]�cW�E��%d�ے���<�ɾ�ح6�n�{��\@����z�٥�޼�5E��Xٌ���j�Ct�6�f=W�Y6󘕸�Zo8�����q��;[�[̅Aw]��D�����{G����f�-�]�Y.�s5�O���]�U�D��h��a�ߓ7W`^�M����V�M)n��\��HX׀חY��𫪀떆����S��H�X�'�U}�U�alĻ^������==ޣ�J5H򚌃��y�y����=w���x<�;��e���(���'�)�U.�����+S�;��{|��*��5�'��Z�U%˝��Hr!J0�+��V}s�U�]q-�i�o2�OrN�v����%�۩���=�]��������v�f��|����m2�-71׏S�4���p�5
���->��k�k%��4��<�G{������Վ����	����ݨ�a�3��D�f0C��W�z��N8�u��=������DW�aE�v\�^����f�a��b�M��Nf.�?	�:/g�=��4A��7B� +��Oo�t�4jc������dw�x�J��rjo[�>>�anc��[gb?]*��ں��kaf����;������8����������.��2�5�Ř�M.�kƧa�d��ழ�U[f���^�TO��F��>mQv"�k�����r���e�df�WU�9���^,��Я5����&Ɉ�c�;����yD�Xz��_kB�E��!~��ʖp�>��/b%��3��o��%�xic���;N�>��q���oT�ʔn�ich��#�ك*�=0��r�w["�Ȯ�C6񺧁���~��L�Qe\�ޗ��ݳ�a]n%p0�0!-�w��!����DGGT8��"���h�;��s92Ѝ���x��w�di��X�hey�ڶ�e�nx���w����T������t�����9����{���4�᥆����V���"�i��η9�TǊVU�?��o:@�On�K�������Wd�t5�\W���\���N�
�~��k�6�읝9�ٚ��6I3=Xi�e��~�Ž�Kj��asX��8��y�ٝ �pG�i(f�5�e]�F�@����n��ێ�y����:����[��<�J �4���`Q�I���\��3�um�g^�왫��C��5�n���s޶�O Kw��X�ԝr�F�9��K�I���4��������}Ӵbk[�<�T�h��L�]�s����-�6q������B���ޥ�%�+�<�=�rhI��b"��"�����[�C9�םm�p��*���劽LH�M������'�����*o1.��^���������c$�+�����|�6�zf����{w����櫥�[޼
]LO]��S���{̽�� ��"�F�-i����T^����7�xU���밎�m+��Q4r���۸�l��Lp��]�VTE���f&uҰ�	��+��-"y�kr�0�C\������.⡻��/�O��Y�R����}��M�繷��,��ܗ{ٷ�t5�ܫ�`"D>�G��H="4�f�O{�w��o�w6�8�L�AnkѼT\$[C)�l�A��9�50k��S-#�Y��,+���O�G��e*�e�Q�6�Y��,��^�8��I˺*��Һ�Y�&6�~���c�z���+����u�]@��\z��1��7�{#�9����t�wK��9:��\����2;�o%��;��mJٳ�79��L��(�,�]�g2�cq@��n9��e�vUr�kޞŤk�(����ҫ8�ב�̶��lF�*�\x����o��$]��No~�37��^�Oj�aF~�9�{J�[�3�77��H�w�4�py �͎}�����F+�ɤj��ԕ[:%jw�u����o�����m����օ�����:��׎rca歋-�q�}���y�M=�e�ȩޙ�p���-SQ�n9������KLQ���A䅔떫�J�8��Co^e*����O:j�3��Ux+H�%�'|}.�����\*5��2߹�K�lݘ�ý�����`,˘���3�2��mʎ	ozee�W\K�p:x���j�'{�
q㉿�tnZi��o7��^K��T6vY��OW��U}!I���$����$��IKH@�~�$�	'���$�0$�	'���IO���$�IO���$�@�$�H@�XB�p	!I�$ I?`$�	'���$�@�$��B��$ I<�$ I?��
�2��"F� ,~f�����9�>�^���SZU$��f�E*���)���1
��E[2����i��BZi��m�ҭ���Ui��J��U�*i��eeP���X֢��c[iF��ee��ٰ�e��ڶl�
�ET���m����n��Z�l�j���-���j��[�ݚ6Ͷ����1[4�����Q�UD6}���f
�mL2�l�l��2���Q�ʖ֪l�SXi��mUM�����-��i{hEP�-f��R�Jlmld	���6U*��Z����X��e��  k�J�k�sN�΀k����[S*k��*t)��\�	��J&�[�Q]5+�}��#B�u�uMwn�����uS0eSw[P:��T�QȤ�k6V���j�Vn�π   㼽��;Y̺�eKl��VP���E�\�ڶ�n5��T�.�;]w"������+L��[�����n%P���o z(P�B�w�mY[�V[V��K��f���   ��B�
(y��(z Р
(]O8:zB�
�/xP
(P <<�(�
(P�<�xP�CC@�e��JBHmu�C��]7w\����n�N���w�G:��M������kkG�  �<-I����H�6��mv��qڮZ�˺:�,Rkvj+;��EUV�;��)J���
U:,]�nJP�D�v��R�:nUq�N�@�Y��JԬ�ǀ  ����֫u���J�:ݶe����p�4�m���cKgN��˅��e�΃n͹������8j���]�:��*�m����f�ջ����і�����  �JU�Z��,�E*V�r��"c��������۵l���eu��Q����h�+�q"�� ]�wUGTt�!�]�֍XV�U5�jօ&CO   mxAzk@�8 �� ٔP;I�Z�S�㠧A;�q�UMu���3�[����Vf�YX�e��hJR�  �h4 �` �\��P�� �gE 's�Z�r�l� �0)�wc��p4�����smL�)e������Җ�^   &�ۻc��U���@�]խ��T���w\pA��qE 3p ;����Gh7[�2-�[lV�>۰Qd����f�  u���Mm�T[AT���Lt������U:�S��R�"����WF��]0%(���`u)J�V	���K�wM�m�� ��eIJ@  Oi�$�(L ���)���b�R  4 E?��   j��Ji��ɠ  $�DM�JI�a�:����(���:U=����	s:��h��M[��dǯ��*�f7�����������BH@�h�		��$�Ԅ��$��B�	��?F���/3��茤��ӃNiB�Տn�	x�y���$�	C�����N8�z/��,���ԟ�V�72 ���On��5��yS��1Q����͹�-<j)���m��lk�k+��Nn�� V%y
�TS,�\����K�&/��Mښh�b=��5�I��R�iU�.��v�9j��&������	��M`ӂ�p`�  vn��MZ��hd������(�qʍ�(�(+�b���3��˅a���UKoz,V$��Nf�a'�D��X̊�y�/lL�"h(��l�|�x&sO���R�Kc�hjP֣lh�V�솳`F���BX��!�����{L�7.�4�w.�F"����AL�_K٧m[s6����csQ �aeІ,yR±���Lm�b���O^]14��S
d�˅��*����4�Sp��Zh��",!8�<��i�"
�{��j�����E2�����S-<H��".ث�J��]DQ$f�H2�Ugo牻�X�j�Bi)�ا���%
wJ��2���di��n�6�P��-�֛�M��� ;���-��=D�0��$�R�.V(�-Q2��k]e��h,��nY�tTȖ+BU�b����*'S��1��_"�jՍ���aҚ�[nk�܃E�q��Z6�D[7�Uf�H�\r[�ײ��}�(o��D�AC7m�/Z��j�`b�@(�y��8�zn�a�6X���lݴU<w%�}�3I�z�.|��TWWjԄ;�w]av��t��0<��m1���� 4R[�T5b���lMa�R��̥5jJg-e`бk��E-и2H;�$�,�|=����-�'	=�'��sF�0��3v��/`�n�E������sV/pe�Q��)�i�ܲ��t㍨w,E��D��z%í��_�T!ᰍ���.��T��h�Ź*�ُS�L����i���d���L���`t¼H\k]�U�yy�.�E������)�f%���Bf�"ͬ��X/hku��EXU6��֭P}�uӉZ ���"����LT�R�bbCQ��E	�T6`��.����Fb�:��`[B��Xa�4V����P5h���+P�,���]<�0ѻ���T�^�ժ�oR�HeK�(`�E�%t������&Җԙl�am��odYl��;MU��E�^� hZ��e	*���T��²�zvó,n����t��0m��J��`:x��.�Tr�P�3bk�T7J��V��`�\c3rm^[��lVv�c�iKa�5�߯C�D;��f[FMF%YF���(��cu����3�$�
�{��,C�D;;ˁ�hYM�Uؤ.`&�bx�`���͇0e�[����5�/#�7eef��E˶"8���a�9Z����n��X��}��Sձ�p@��oF^��̺p��5��j��f��Q��bl�`���un-d᫚�2Un[L����[���ZA(�����A�;�,��{�b�N�6��&{m�.i,aqŔܖ��5��w��{{Oa!GhRÔl9���6­'(�R*���7�Qv6��Lؕ+f��N4�U����wbŨ�r�T�e�e��e-:W[�ee�J�`��͘Ԩ,�Ƞ��Ş�b��kW���^\��o�&,JI^�PpV�cKFD;�e1���X��)�@�R�|���;"�|�ѽQ;ב7y���ާs.�$1Z��V�ژ*�,�e�{P����F� 5�a|�?j��{'��8���]7�!LG��ȵ���eؔ�f�3�,�	挐]���#0���"��)��w2�����kYcU:��e���*5hSV��J�p����8ʛ�r�����v�lm)V�h<��L��E� ��s0�c@B�L�X�����jh��ذ5�e�2Jq�n�V�^@�R��[F�U����w+*��v2�+��R�j�ؔ��)m$*,��ܗ�(��J�u�A'�S����9tE�JTm��@j�����؄�4! �wjfЙr��J�0�1#2�
k�Xja�Ӄb;`� ,e���k5�LQXJ7��P�N$�'��n�b44��W�l�J"%���O;��Cb����N�j[�����V�V��F� ("�����0e'�z�mз`�h�sGe��;��^��T(�1�e�A�Yu�ԡF��ש:���ڪ,����x��@!3�7�.^eںV�^|"��2��ʻswr���\����æ��Q#[մ�՟�3+3
�-��*��e��`�WO%1�J�ӟhPG���m� ������ʽ�e�,��:�Jqm�-��J�M�Ir���3a�jJ��!\w2��Hӈ��������Y�i�P]7�V.��{����InNds�H��ma$�������B���"%��*�����:�{hA����`؅m�ҧ�S���a/e���h暇3��<%���:C;��^=��+�� �r���Sy���ͻ��3�W[�ڲ4�!;
V��4)f�˔[5t����m�u}�0��C̭/����%�ew�1�jskMb9wJ�o�x��a0�k]�:������:l�]�w5d�6ͬ�V渋��T�����1�3�F� ���Wr�4�7�6�d�%@m#Dv&��������9�'S6�.ǜ���������:s\a�yp�mӬ�%#K]�Ik׋!W�W��uO ��d��FT�"��rG��]�8uʈ�^�AK ~ŸiX[�E��B��Ya��*Y�WX�%��i�Ԃ��.Fb�m]ml��#�J�N��a蹎����{l��������rR�Q=�d��Q Ę^�����zM�x�[�4&Cd.��yqS5���z���8/�B��,�4�^)��²��I䐽�ܣ)нz�{�ݕ���N>3��(�YC� !!z��G|2��1흠�o�h���3�����9#�Z��w&��5`ɟ]X��Y�nHQu�{4S1-+��KZ���o+ �nb�[i��ISP��fk3��RƉ���h�4GIP)��׍]-����+-��I�[�L9��n�d�V�ׯ$Ќ6+5��ƕ��z��ј"�#kc�[�k-�ң��f�Q���P%�Z5�n��1]�3j�Xئ�"0R2�aִ��/Y��"�*�]=XoKwhØVL�?	<����r�*6E����TE2U'Z�l�4D��s�%�JB��oNV�	��X4�+N7Z)�����>8Z$L!�r��#X��B֚�Rܵ�3����t�a�I�f!4�ѩp�/k-�6��j�Y/&�ը�\4?��g ��W�#�Qu��,�ZEn��5��sw�H[��h��{Rh���)�&� ��Q`L9F���Ę�hWb�`}�la�r��.En�t��$x4��A���H�86�{r$�!��������H>��G���^�Ӏ��:�1� ����I��dz��Mn�u0�a+l�#��`n�`Q�Z�	�$\쩕���H�B������y���O�v�>ҝx�ѱ�r���c�*��T/[�ԡV� +ǲ�K׀[�)A�4�[�ڕ���~�&։�p���АB�{�נJ�
Кm}5����5�.�2]^�m[�"V�Ǻ�WoLl7��U-w��^Ll�B2bi-�V���'sKX~W��|������D\����Qdj�$�Alځ!�܃�i|Sz �N����pX����fdv�Yq�iȭ�PB�]�h����݌��p��Gk�7�W4A^ж�'e�F�&�mQ��]��E"��eG���`�{�$�����"��ɚF�Ռ��^�FIYhG�/�JJ��٠�!��*Dm
�DY�.�����N�7v"��&���zRn�&GtN�.I��ͤiJW��(� ҆4�^��<�oAV�O���sp�j�}��љ�hV��8db��p)m�" iQ���D�u�im
������d-�9( +0�J�Q�ل�j�n���9�#$/:�n� �Y���$��S+jZ�nʹ��N�ٚm����Ƶ�(�-C���J�#8�E=͆�L9���U��@�/.��iAGM���gt#�ll����sM&+3�M�"�jfXk~�L-ǹuJ�����;�$�ׄ��)��q��a�t�J���qmsa�T��pj�Wq����hKB�ܔ$d��XR[G#ܻ��92��J�R�����Շ�\�|"�C���yx����8�دr�:��ʒ�ҫ�� C��**8�K4B2�Y6n��E�2h��׹A�6�m4KF̹���"�b�noq�(H�r�0\���6�~����y���%��QEIN���nk�T.��sn`���v�ƨ!)�`a�n5�����AJ�5V����F켏4��[ZRn���6i���0�1���2�ɒ�@+N���Fm���2T`c��SPZ��8�Vn��%շL7��*=�f��x�F 7(`Cuj�R��^���U�o�M�5قM���!�@1�l�`$����<�+�˞9�D���sig>�(f�FUF&4+^GB�^��RS*�ɋ4H���ކ���ZWB�7y���5��@��P8,I�SqZ:��q�x�C��żf��=հH�襛��OJ�v�;R��Z+Cǈ:�/5����R��j�j�k�ƕ蠔E�bH&`y��l�N��9������<tBD<��|y"�f��,�$q��#����p�� ��[	+��-Z���f:r�UJ�AZ��ճWA"E�nۓ��N�lƶV��nA��]�wK����bl�#�F�];#ʻ�) �3M�r�H!��e|j�lcD8Mn#�	:�=bo�7��k�99�-t�@�K{Xn���WT��Djm�`nD��ȆD[VM^b��	j�D�0KO3uȍ8&����r��N��\d��M��,��ԣ�4����B4��a��D^��nlhG[>Ԟf�A�CtnE%J͖����Ѻ�)D�7�4׀�8A�H����� ը1K6���.Zt���m��K�ԁ�X�)��d��@�N�t�xڥZ��jU�jf
9��Uu�e�?;��̆RF��\�*��o�}����q���2�-�.���=j���i�kYG���:����o+[J�#���H�]6	��VjX�7p��Y*�[��"`A��YF�e�t��7X�c����&��ы�0����~Bo���=�fm��*Z�5�)n��m]�֠v������X� ˓D�_�u�d��nӰ�(��d�ce'�m�eR {^u3Ş�,nj-<�f�G
'h<L�Ȉ�L�n��ɹ�������n�kU����oE$�W��+[�V�,^T�hɩ��]��W����-�8j�����ZJ��A��\Z���X+M�3\�H��J�?�-�K:A2t���b1�91-��t���Q��c�X!݂#Kh[�*-��f1)��{wj�5�6��-�W���cq"N���=�nְa5f7u����{n���5bK2
����qV�;�mݐ����x-n#4e�٨e���4���!q#���ԝLyZ�{r��х\����'u�ݭ�LN=ص՗o&��Q����
֡V�b���n�F.Q������Aˠ��1���-貎�D�hj1;q^B��i�K��8��BZOhf��LJ�lDV��I�AM��[,#oi�٫pk7��*��6Ƭ��+B�0��X��6�jl��$�f���3����)�ֈa9硬�ܹ��T��N	���e��V��=���(����O Z7�w�?f��Y�I�nЍ�@VIx��(�v�QtM��W�`��W�ukTPł`�UM��9)�2:�~�0u�4MXٔ��%� B�4toaL��WBւ��U�����[E�f��b5���G�}��Z[$�zGd!�܏0�Gf��h.��!N�d^V����һ8���T���P��v��1�n9B�0���V]J�ku����d'�"�a�Ӱ^c��^+n�<xS�kw"�\��M�"�����P�D,�E&ɰ�jb�E���Vb���)L��Tč��zZ�X&Cp�j��@���*Kmԣel:nں"�X�՛a���l�{I�>�s
�[l���>a��bS?MW2�;��R�Gb��X�bmm��)��
T��^B��;6!� �^��29F֟{5���:��)�e5��Q����U�bLr?�8l�����Iwb7"T�͎���ʍ\�h�'ldW����
vձ�y����-JH�fXZ)L2��n嫶�[F���5�[O*�|![�����Ø���G[��f;��B��t�i�*BMZ�k,f�Kv4��U�(�/�XIu��Rr��(nʂɒ���R�HŊ����J�5x�ԙ��	uu,��)�t�+,20\fA��fJ#,�� ,TD4�C!��6����!Ue�7J����/^Q�6�V����JTj�[H^e\��P�ɘ�PZJ��,��.�VH5�v��P�4��qY�X��F��-d��jR��kt,���p���	c�[��Ϯ9���R�!B��7(f��|Z�)b���س�d95�4��̫!nm\ˉJ�V�a�W�Ar�,ǡ�vQ�[��q��E�!v�\y��d�������5�֝���]��Aڮ�6��1>�k����[EM����w+�Ҭ1��c��m,�Φss���٦W��>�;ʨ�Ȭ������c����m+79XKý����W9D�OPbNkW5 �����$��NZe.1^d��f�=�=Y�1�Rܓv����p�d���!�%�g�^iU&��n���@s�9���2��w\�9r}49�SEC���t����xi�A�'m�t�P�v73&.�"��j��Y��+��[j�����d�X����!�Y�أ�d`�FX��d$N��ek��`ͣk�otF�>�/p�Jƶ��y��2e�N��E�̐�|�W o3��Κ��جKEÈ��ݖ���Z�a��k���C����q���Ou6�����=7[[M .�[O+.;
s��5e�gWJUֳ�G@��i\��|M�Uj��mY��yѯ��P���Թݫ��]��֚]E�B_fB�gR���������8�v����ˢ�$���|��V��uL�i��:v=8��<VL��m�R�m��WӋtD��bń1.���	#Y{}jڑrե�m �'�2$���Q�&;ּ<8f�!s��S��O(n��D��z�MԌ_.���ɸ�o\�ٻ�U��R%l����l�vv�!0���6��Z`j��B��㠊�����t��M�L���wĥ@⣦�訶��������ץd�N�R9x�fmf��I�,Y\�b���T���r��a�s�z�s��MӃ��	�ہj���q��_V�sJK[�^������̦�G��&@v�S�5z�9�v�0szk;��+�feoAA�iB�üi�n%�0{��!�p�*�f�c�	<��.�푡������ǌ�s��wn�]�T�rr�����T�C�R����#������3����s3O+�.�`�yb7���HF�/��+�g�����X��/����w`��I��Mw5��820�$|��Y|7�{o�nd)����c�b�.�|xnvNA����;"���Tyy�n[�Wi�ۯ�V�����r`��XǺ£C"}*�*��8��V�sNU�.Z15�ٝ�:b��(.�<��%�����m�u7��Gv�p� q"����d��|-����u)m�縅8. V��q��{y���[����h�Ήnٽ��4b,RPD�U�T�t�o�eV���dn�u;*>�NΕؕ�W`�ʟ��/����b+���0��'�uej|�1�#k�ɠ<&^��MV����wϵ��	�w�ZR|<�h�Eovd~��U� j��,�'�¾��i��q��)2C��[��M�wY��_ٚ�v�+�`��[�����u�Q:�#�Y�3��|��+�T�>F���8����F�Ҟ�gvq��]2Jw�h�a��h�fm�o�G�ޱ��v�-����$��,�!]R��n��a��fq��� �Zw�݆78C�!2����꾤�n�k@���}�'D�Cb1��*H��Ѭ�EF=Y15z5D"�S�IBV2��k��K����,��c.rz6�	��)6¸e�\h�y��m��ŋS�h�ܝj�]C�I8��XT"�9}�F�V�x���q�Q:xn�8dUӰ����C4o�h�4I�[��}���u��&�1"p�(�)�@M��H��%��:1������a�%kyPm��ou>�EU���õgQ�u'�ŀ!���W���}	��-��]�wv&���o7n z�����(;ٓVC=Zg}�A�����ͬ���e�e&#�r��*}�%ǮJ3�[׻���ݡ;qR�p7��E�_��#���p�ݳa��^�u�A�h��������{����^a-O%.�<k����G���X�]����Tbg��+�,��-�-��n�y;���g��{(�A��	�6��l۳̭A���E{�p7Ԙ_:����W�lŞC�Mk�i��"��{UŎ��/�_ޤ��]ݗo�ˮ,1]!f���|&�p_���xhr��QttQ�/#�믺a"�����:�e��+�'Q$Hz.�z�w�iG���B7�%|�1Ҧ^&+$}�"��;]��|{Zo��g�^�٥�"�]e_��3<l}�</�V�uȨ�	������V@��]���k����~9s@[c�چ:��A2}Z�&�QQ���j���UƵ�o�̞��E��@M.��8�H-�e�HcTu���;����\��H9�&\-�qi=`�Yg^��7"�h����e�
ga�X�z�C��߼�k7�؂G���k��IB�(Y�9���}��"�βs�5g+��-��b�@;w.�|6�a���Dx)h������"��X2��y�uo�8;i휵��V��j'�b���T�k�,����Rk#�E�R�<9�oL���uȝ��P���1�P\��Z�s��s6�v+��7�G@'���Z�AM*�#�WU��f)�Z��WA��0�{Ϧ2n�j�����,>a�d������Uӝ��S��-Jvz�̙�,O�ԝ����MA�Pv.���.�G\EX贾��eki����{�\�h����^�s Y�ܭ�7�-�0�$mWp�#Ԃ��G�,��+�+@������A��Ԅ�Iޜ��ps,N)\��0��JM�jgJ��=�c%:�h��V6Z�t���~��1K�t��*&��Ր��	��]�V�f��L�(�%����Dv�ˁs���5�S�oZ��|q��氞i�WB]�|)ܭ�8�[f�\��jy,V�&U��'�U�1�r�����G���IؘU&���}����;�H��dvd�a���9H�e�ע�n8���_<Sy%cdu�4���U�����#!N��N��&V�K��zة�^"�0.�v��g3:��n��4$r�r�y��q�s�^�����^]���@$>�pý��C��)�����O�$��Z'Bd�mN����eE��'p6���}���e\����a�.��=n���,f�APNS�oy�*�Z�{�2n���g&i|ҫa#mwb���7ݦaH�ě���u1*7j���}��.ӊY>�=��v�
�O�o��yֈ�)�6pǔ��Z�e�v�	�Edx��=���R-*m[W�$�TV�,D,e���I	)��WK�����B�}��O�M>u�X�v'��%5�Z��Ǜs4]ʓK\Yo7H��纇�>��t?]/�q�ﮡ�C,w��:�D��ۚr�%k���|e��B�F��|� �gW#â�s��(.B	��%��b��m�u�K��8o��+]V���D������$���e�.P<M�l�˾�.T�[v���E���J�b1-�&��G��^Hb�iV�P������Q������<�bm��!>��6��_3<O�U��!�3i���Ra͑{ː���g��מ���L��"�$`k�I��Yӆ�q�FS=��,��y1��=����(%�X��=+n{N򢐍YU��W���R�2�[�������M1P_����E�F#��V4�����+�F:'[r�6�[�蚢�	��k�ih�r��w(��ܦ�YƉ����Ho�n�:��ϷN���Ѳ��`w���	Ub�=���1�*���.�;���ۡ�z�t���	pQkw|�d��
��㼏R�?0"�u�}�]�TuKf����Զ������Jt쮾܈i\*�gY[Z��[�����50�[��%�v�ۗLR��~�edH��l��*ה�2sg��8�m��y"s���j�4��ʯ-sY#Py�p
��F���"�4��t�b��7b��5ecpv���t�j�2�t���]0u9�N�s�p������%��E����4��=(;��5vC�M�p(��|��u�"��ί�,���R�`�Wq�����C��<��y��\,��<I>��W�T�T�+K�+)�1!�vZs��S5h=�( y����M���N�#��.�|x��6�����A��r��:�0� �QNߠ���Ȍq���$b�;���e}T��ZhHu��|�"�-I�W[n��C~Wv(WV���H!b�{�׍Sz覾�����w�5�i�w�_S���;OW#������ݗ8��{51e2��y�3L5�u��3k����4�������KhooR-�;v��C*5�_.G�}GPV�^f�γ��M��x��u��w=G\�D郝�l�DHhC��j�*�"�Z�\O�G�$�(��]8���C����98�W�mXXd����7UEݹ}}�Z��OWa'�_��/��gcɧT�*�<x�(��EAocF�)�G(+���b�S����ad�j�@Ϋyv���4%��b�h�ڕ���TL���o��4
�i�SL��]b�T�sj�An3�P�0�D�+H唇8Lsz��6�-�n�����7��5ζ��W��/PT�jlv�B�P�*�����^�Q�!_R�k)�燕ϗ����ӧs�D&0�#�FV.d'(u%��۸*f�(*ul�R��D}]�͞��{k�����~��a[@YV4�\���{N���u1�c=GxN�<�GVQ��=�V2#�9ff��z2iv��R�h�۵5h1g���Hc�i�3<i�����$5�p���&�V��ˊ0W��"njq��'�{/R�]��j㽱k�S ���p�ڌY�r��l�V��tɭ1iX��%[����k����.�WZ�;㏪��I��Pݨv�y}��U�-�K����zz7���k�u¥s���HF�Z��cjry�U�w<Y�C��X_|�Z6��y�x��od�p�G���n�>�gh�tܢ-�(57R��n���s��������ziw���֒93yL��d����,��L��t�],o
]Kp����|��RӸ(�}����tlz��3�m��ݸ����v� '$pc.��"-Q�4�}��Ll���7�;}�Yf�O2sV���Of��M�>'�7ơ-x��V՞�z���u���2n�f�ܵ58��nm�O#u���Г8=���:Ý4Y���:�3D�:s&lww@��}�[�Nt��P�Ԣ��n���;ll�R���Z���)>A4�s99�o��,}]�oV`��ޛ<V�PoF�~��Az�%����wRD��b���<�i��mc<4���m[��L����� Zi�]M@+�Z��_]m����|���r��]%}iw1�Ǘ� [ه��j�����S�
��/^.-�*�����7������('��t`�w��bbjWR��Dnw"u�����A��]>��S�4�cZ�-�u�2�k6ۈM]f}�S�*����-'Ճ7�c���6Z ��k��"�`u����M>ؑ��;���A�_c�n����{zE��T���w�s�}�98��&�!����xi���q7�E���Ҍ�E��B��VM�7�w��Y�K �����F7}\��T���.6�m�Ø�Ƭ*_
���Nݼ
�w�t��%X�uk��1��A�����0J�u�S�B���˺�떽Z[(�ԙǙ���� ��ܥػ�����u��Rt:|��i9@���9���:�b���u���ƺ��p*n�;�j���s���n%�%n츯]���Y����C&i����
�]��]�v��� �^�-[$)r*��R6�������Ę����xtZqk<M�|�eY�{;��o�sb�0�.(m7�G�� !�����1��h��4��Fv����	���wd�u[o��ܽ�f�_UtS0����A�6�7`�jv�}�r�J��]�,�Þ�mX�_n�i�f�Җf�%m-E=�C�Et��4+҃$j{�����M�bR�]�;��*z%�v���;@�k�'�p�D#ʖJ6���4��l�S�n�$��J��'^X��x�YF��b�$G˼� I�J� ���y� c�-!
�+ݳ������h�F�jZf��n��ݡ��6�ܨݎi��R/���+{��2f�C$���s`��|j�lS��e^�G	�����)�[q��W,����% �uf5ҍ4!���e�}���UU�ދ+.+B�q(΂���YO1����5n�x�~X�;x:u/q<�`Ŷ�l#μ����*��z;3��wZOy*�P׹�^w�៬�$:��*��\�#N�ݰ�r�}c��Rb�w9��N#dއ 3c�Rh���Em��jͬBB�M���w �Z��#J� O0����}/��H/yk��Z���z6�;\�ʒ�p�>�ՠ՗����������c���&��7e��{��B�#ص�+E�]]����TÏ�/�<��1��4������)�7J觷��h=�W�9��Nz��죴����jJ�?fu�ʸ�Ъ����ҷ�j;d����Gѯ]��d�.�e\�����e�ogJ�R��벩�����5hJd׈cSp���M�7�{w��A���B���]��_;�/>�nX�/<��؆yiE��"d�Q��t]
>�<��ɾ�k�h����Y+��EJ�>�]u���r��H�'�\�{P�U����kq�2]y��'���F�p!�7�Cb��W�\��)r8��ő��c_m"�����v=�^�f]h�2�����-�ZAYo9M���Ͷڅ��(���n{�>�������}��A! ���@�$��~�7�8=P+������N ��(����{��~N�v��\K�}�Yku�0��S�;'x�wZtរi��'Il��Ŝ�5�7n�$�:Qxl^n�v��QWԷ�R�!M֜ȴvJ�
Xt���n��r�.m��U'�H��-��{����tn��z���4 ܝs+epJ�r�g�YLU�䫎'��[�S��֊xLW��]j]��^bi5c���/mf��5�Ua͏�+�|:mԙ��o�R�˝�{���L��`�S6�+<���F3v�l����ak&���,-P�_U^��Y�����S�'���U�c7�#� id"�5#�i�ٺ|��6���9{�ߣ�R��9�SWKH=�M˫�KҊ�8�x�2���b�%51W]\��(�ڵ%�{Z�m��`7$zv�0 șRۚɗ�.��=
��_)�Z����z��.e�3(����iX��|m�	�������7hv��o�����X�у��Έ�9|��/��W�v�'I��h�Ұe۞�Dv��i���6�.w��G	yK����<40ƕ	�ٗ{�x'ۆ�
*P"G�`��l!s5Lgۯ	v/a46�h�yr�k�<�ڎz���b�j�n��W4�95�{�bw���Mn`��~�Iw<Y��(��}���k�;y8%�/�#/y���^��TY�Tf��.5W�oAR�N��}��r$k�ST�-EҞQz���;c��m�w�M{�2o��B���@�p�U�1}|͛���)9�ؠ��c�tG�]�ǥ�y���Yj��I�N!V��8�8[ҝC�%�$�,��gEX�����v<>�:.�{T"8��(]豸A�`{~�qhG�`�b�M�+5�������V(�Z�<�A2�V��l6�^���C�c����[�{cZ� �[t�YvtW[��^:!4����Ӹi
�q� ��:���N��vm\�3(xNvF7�<�<�^Zt�R��=䦺ۡۉ��"�ÿ��Kx}��=M�vi�+�rhq�PK#"��˽z�q�e�;�������&s��f�X4e��@z��2��!f�Im::�]7��o�CL3�����m��K)��z!.3O�bq��[�gW��k�X�;��0QA�<P*K9X�3]���佚y��|�L~�E"��혴����c{���	��XН|x ��q+�͜�K9�jy�fe�'B��B� ���'��za�����7���yfP6�7�R�f����J{��=�R��WY�$+l��J���*YOa���ɡ��,���mi�8��Nyq�F�����UJm�om��K�y�in�Nqnۂ�U�J�7gFc��]{{b=��M�, �����t�B����gd�1�ԝ�[��:x;��]Ѵ@S��j)�����J7Y:sr���J���Ijv���f���.ǵ�ÝV��!Q���r���Tr:Y�8���
8�8�{��J�(��	�y���v�;�o"�/EzRnĭKk$8���n��`���ȯ���N;�ûS�Pڢ!��k����	�ͽt��-�����&k�E.����N�qF��%}ѡ3��ե��3��s�gU��b48���e��ޫa��wz��Pv��wk�H{����FWp�7����5o;?S�M��R��D�ˀw`w��6���j/�v7�nrM�[���-c����$;�Y�J�&{����f��Jr�Wb���\hvA4����Eˊb�m�7�_`g�]��&I���7>9�9�h�r,�t�t��%hC��GM��Ķ..��^<2c�K��'�S��[XZ��{��}6�*�ǵ�I������`qy���\�4�8E4\�K�b'ͪ���,���څ�����	��ތ��z��9n��c��}�&{�Q��W@n�W[��ưS�o�v��:PYW`�����}:S�h�t�F���Nj��=u�
o���b�E3�η�<8k�0AC���ms��^Y�}-��+����Ѓn�rT����n�ƺ�H�\���h���̓�]#"Z����T.���#+%�����G�j������7�Y���WqU��ǎ_E��o{Q��X���h���T����)�w�����;��8Z����6s���e�#1.��CWm�D&��q��X;]AE i��J�f�r����VxA�rԋwi�)��g{���-�%q��)kJ
0/��_e�"��'
��_<jP�X�Ţ��=���׻N�|rKc8��o�ws����$�;*Z)��ݙH����;o�՞P��[!��ū<%�#ܫ/�Q�����j-h V���4>����l�F?p����_YE�FQ���u��uB/g�b9��'wx1�2�7�T���c���{i�k�G��n��q���ݻQ -����3�e�U����vsE/��'�� �����zK��!;F]6�O�Ã2��ngm8�8�]�#Yu2��:x��:R�Y��3��р�{��k�i8�.�������;�j��4E�rޞ7��j�ZDL0R�0�ד��C��{&�����}Q�6
/Nr��-byC ����R�<����Q��ati�5ݽ�-_Gx48<90
��c++,k�sيN���1S�n�G�o���xf�M�iG��=�<�=���O�vвO_X�ӠnT� �]��q����:�q�O����k����˫0��V��.g�h��+�?��)L�w��n8,�;�'��m)�e�"�+|:�=���wr�����r)�Hz��q%��x���js�9ހ8�EĵY	�u.����oX�=Yg�S�'yŗ�;Go*�>VP�GZ��݃5�%i��Ǟd��h����5Ӝ�U��\]��3�*�gd=�{q��6�4�]���1G�m#�+;�rb��Ś�B"�����cC�ޗ��DQ�%�ؘ%C���ݜ��{����;�Y���(�L��鏸Yad�vY[��o��H���.�a�[��}X���_Wr�E��w8� �9vy���Y5
��N��T����䳚�n8M�x��#�AY�2�{����V�����+M~��H�N��kD��W�҆M���{���(ޖE������y�L������� �6<n����t5�l�-�$��^��qTިW�e]��w���ǆ����q����8s�+{(��S*�dn��~uxCۭ�T�W$4J+7���qg:�J��eX��m*2L`b�f�eY�J��Sb��O�b�/�D��b��wC�M�L�Ҭ���}�s����r�=9�	d�H�H�e2���q-�5��	H��;���l���7��������F֟N�GR����gx=��xkz�޾^NDH�C�L�Q>ۀ��ԇx.A&���
��Ւ�j�r3��;�����z?���"�M%rD�����e�vz��O��ký$H7��0��(Ѿ6�'5U�#�yǴoV���0�RD���.34�R���g��P����}\��(�����t��y�(�g|wF�t�8Z@a��\X4�oƺ;��1wq�8�ð�	��s�5�-�،}�b할cէ �|�|�܅�D����y��5%��k����ڗ��lSxЦy���;|�R�U���r'�p���w�c��U4���V�H��cD�W|5�tm�=��.�%��q���
�u���kF8sL뭦"����­�0��:�9�2�bo��ġ�慺]��z�w�7sx�_"*~�g`|��9n�t���RT�b��J��fq���7I��r��hb&�J[�/��IN�R�E΃k�_Dfe�N�)i�^u�҃�T�:B���uϢ��}[��5�UԴ�g]���ːmoF�K�gZ5�#��8L�u	����5�[&sV'8�Q��:$�n��|:V�i=��'����W��m��o�3s���֝��~)�r�ے��WTaNy�޿_1u��&vb`��m�7n���K��i���i���(�Hgb���-0��{�(|h�Yӳ<�(�݆��]e+��L�OV,p.���Ϙ��s�O�փg���Uh+�}��u���M��-���o�`Dnw[\4إ��rCgu��&�E�c���T�oR�uN^ScC-2M�L�<}�xL�����s�W���'�G!AS��ų� Ri�Y����L��Y�.n� -�١ǲN�ti��<;}��הS���maO5�u=�ƁG���{?k��˨�h�h_t�a~az)=xx.���5�K5�}RIO�vVw.��y�ggs���Be�kwn66�|�6s�n]*�v��q�V��|b��mȂ���D�7ޗ��{�� ������m��r�Ve��M�GCսv�{��L�L�s�23}c�X�d���z�7�W'A��Yd��:oI�s1�⩭m����v��8�;�M^%}���GCg����	Sy�̨o�+�v��\�����-tΈV��]O=�1e�x뻠�et�R����gP^��|kxv�H'20c�\����&���l�J�.�N��ָU
�mZ�ݤ�3Vz��`8�������a��@7�)����]�I�BOg�V��H�78K���v��-���Vڃ�iW"hqR6q]�Q��J�L8�wx��[��_.e1].�:.lawm��ͩI�V�$���=��_s�P�hu\Om㞌��$j�: ���]���Ռw�Ι�&p��^+�tkJ���zv�V
��R[�`G,���J42� �1�Q����p��'=f���T1ZĎ�����<h�l�q����R�u��jCqp{�����e�0W���,��J%�&���w7f5�r��%zh�@�U�g/�-)�/MI0Q,�}.���YC��wY�	�e13;�r
y��Yz����2W'�ku$�Ʌ��	&�o%C�@��H]�?m#�ܒ� DIy5�ȴc�m�jZa���I�2���}Oj�0�/���W]� �ݴ�R���O^'�Ŧ���I��7u�h��%��Iȕ՛����]�PX͢��ŀ���` ����FDxIt�Ӽơ���j��Z?uNi�e��Kŷ�|�x0���)־o��{bY��!N�Kq ��i���������Ԕ�h�ӄˁ�Ը�̕t��Q�K.vCx��9	���&qF^��h�	�ޫ�f�0,��3��9�_;�|�R����➜ Y�eFL�`9��G{<|�{r��(Z]�7_^��ErEdc/)�\k0F:���!<�'�����9�x\>�#;+�]�9:v�y�<�=��7�1|�9�k�'��>{<&>�d�C�T��2a�3Ny��c����Y�R'Z�E�p���J�ə�vzG��|�l ��?m�a����̍�T���L�P/�������z������J;~s�^���97z�X�<�
(-���mY�r���;-̱��ʹ��<< D��"
�B!.�Į������k��V[ִ�]>��WU�O=B���u�"}wR���U{�u<8��qPu�&>`�|6��&&���v���H۵G$�WF�1�0=ڰ�u�ۥ�����ϪR�p/GVL���\���jZ]y/!�� Ă�p�Q��ifF��(�p\����H��z������E�˺�Y������vn��h�F[��ĳ'`僧`;'bO|���2��o�3�su�����n�1���C��_>�%@��	q��pL�t�<U�5�Y���,P���WJ9�`+��V��3I�����f�4c"'B=�8ް�*�	?��|
�>��1��03&WT�j/)���+�2��M�ӹde�������m*�����7ʧp_�ͺQj���]^<d�� ̵p�+��Rs��-�ff�V��/d����O�t��lq���Nzq�!�=��N{�s�"��J���j�4�<��B�w5v똲�����F���u�Vf�K6�m�ø8J�Zj��Tx�o��o�ǒ�ϥ��(f��H(Җճ},�	r赋�DE�ӹ���VЕ����)��A-5$�Xk#Q�:b���nov�$��5rv`���=q�r\��@X�� �������=�;����8D�Mʣ�p�
�Z#~!���Í��2�`y3H�|Oz�!ȝ�%N9�o�Ԯ5��Xz�͜���5f��u>�:����{:w��_&��TE3z�β��������g��7!��_F�|}�ׯi-�zޯ����v�JB����L`�R7ʆ3���\�����y�ݔ@iSwҎ�˯WA�m�F�Q0�	#Ќ�qp��lf��;O6F�-�x&q&kp�$V٥qn�.��V0�n��IDD:��վhj;m���fqp[O��L�x���t=��1J�����uhm�4���"Zàź���y)	�W:5+Gj��֦����,m[�Z!2�M��W�^����/�آ�8r�z9v��RE���Ӑl�����f�j�D�c�̴pv=Ǩ�ս:�/�p����<�ŭ��G|r��Tw�Ỷ(2%��]�{PJ�E���M�|J���Kh9��u�.� �˭NY�Hc��]
W������G\t�qAN\�Fe@ �=N�W�ɂ�E彪q�i�K��3�ՙX��	˗C���y�C2��ej�:iV��.�Il
�F���5�D�P���<����(���?��J*��no �G�Nق�z�������!�@z>ӳ��_[ekJ���c����v�=!���)}Ba�K���4#Ϋc�����+�d�Q�����+z���2����۵H��,QX��7w����ӯΎ_��k�)4�R������˭���NN��;�g��U�c�n�-]�a�-���qM;�O��3��UN�� 2��*[�޻{�T�nvMݨ����
�ȗ4��.a�bٞ
������"�H�i����O�����I7Nq���w�[�Q�||S�=A�#pݦ̾ν�i��-��h	���oF'�%ϊO�΅��{�� Π�=Ɲ� ��dgD�W�S!\��s�Wn������Wo\^�u��:���ջ�f�'7De�O���(HF���(�>J�Vf+چ^������8��a���
m�	�QlX���N��+*X���K�Y����;�j��L^�~��W 4��d�y���̥������Պ`��A���O@&K��:�lw2�q�8L�gS�����J4.���a�ô���r��Db��]v�\dʽ�b�3���x�K��r��%a�Ү(Zj.
����gt�ݴ\��q�P߬�:�O�vQS�,�r=�yPf��)��&c�ݨ2��jer�q�:�'���+:�];����;� ����U�����Z2�d����B�0�����YXQEZ����U*Ԣ�mJ�B�Z���EEEAE��E�5)JX��c-�X�֊�*�acF���Z[F%J�bQX�J����QDQ��k0�(�Q��Tj[e�l��""��֊""(�ƶ0jUh�e-��b�[R��-�RW1F(�KB�������E�
�UJѴ���Х�l�[,Ie�[U�EJU��-�����Т��Uil��ղR�E����0b��Z�-�U+Vң�r�mQcm�F�n&*c*�)l[j��P��T��\J"�,2�Q�QVcJ�b�E+FҠ�֫Xf���6��A1UQ-�JU�Ҩ��ic+
�U*TY�Z���-%J�hT�eQQ`�*#1PD��T�V5��,k�"���жYP������N���ώ�z�S�E��Rי͘�R�s�I��/��!��������&��#4챓�.V;��J3�C����w.V�\z��3�;݁���^�*�GhP���q��CT;��ˏP���WHl.��#��/� ν�*z��B�����\���Pp��{i��r��cq���tS�M5�ob�d��h�젮B�P(F�N���Jb��>Z�I�ԃUpvՏx��|����q�K�y�&9��ܑ1��Caʲ���{T/%��*�3�Nd-2:uN����#n�����y윈�=/2�Z5���n\_����3�1raǫ�U0�󽽆�-V��R�2/b�5�����/�"��Q��AA1R�V�o���!9�s�yۊ�֮%TQ�m-ְ�%��$�!���x�ʛ=)��5q�w������;G���9!	N�Z�I���lO_���I�Ī�G��^��mi��2p��w{��L��Uh�X��.�p�M�-y`��V,)9���{�/u�a�Ԯqn��	���k����'���nYA��]{�*� h�<� E�t=ஏua���ɝ̤��8��-�˭Y��
��w��%y]t�!��tȜAx��l�=��˺�x2Tu������P]廜J��x{��M�<zc����g<^�l.[w#�}�Fi��g��P� �=�ٺ'�{-=�r�{�<�9m�#�Ep�9URJ��
Tt@~���6�C����茍�}C�h����޲�O`9�.["�䆼�'y�"Q�l~ɠ��p��Stl��D5 �X�l6k"��ߦ�Q���,89���7~ίDe�Rǩ^9�]3�è}�E�GXS�"�:��z;b�U]'��C4��'�t񱑭w�譟�X��U?82�%�xʴ�:��ei�Z�+
�UJ��+�{���2r��t�7du¡�$��Q(@�*�0D�1�&+���~�=i[�f���L�/���dj��ai�U��8�p��W��������EDlة"��]3�-գ�Y��-����:&�>�}��G&z�C��+��<%ӊ3�YR6B�g���!\X�1P�Gu���W�-¬�}�T�; ��3䎹��'jT8���YQI�D8�v��R[��lݽ�X����-�T)��`fR����#Fˁ�gvC�hi�+���	��ddP��r�����u��	TOg	��v`�݁"���p��7����x�؈u;�6O0B���xg��7���C�Z�Y�[=����۩OL:�I:���J�wa��C֨J ~I_އ۞��s��=�	~a�eĚ2�i���]H6�i���Q[��]�jYe�	���%f9�oK�SNX��{r#*P��>�:��BK'n���^>�z�}^�����$��Z@A^��;O���{u ��$FMC��XG5oRa���ވ��4����H��}��}KEa4��f�*�����һ[{{j��Z7����<�l��^�B����(�@��&�p>0L���Y� wJ�$8s��љ�P��U�X�s���ECY!�x�+��A������Vx21��gJg��m�{8��)%��"[K>�+��]/�"(�}���.�g|�^ȣ�fⶸ�-�w��)�v��vٳ�����-c=�jv(�GEԁk)$d� �Q�~�]����M�o'/������׺Tv'��Kʘ���K+�����Wb�f<���F��d�ט��B�#��o�ῷ�qB��Q߇�
ָ=�>^�P���9�+C����S�b^Y��E�	\���!�{^drv�`d���1ѕ������>�*
W��P u4������y}�6��W���d�N{f܃᪌m�.d'*�t�T���W`�]>^dUr�yw�P�Z�/לwn��:����{����\�!�q	r��;U��+�j	��*�D�7$O��N��k��EÌ���J����;��.�1�[х�\bC��p��w:�+�?C����B�����Ӓr�Ϸ�{��c^��;��MN��m�'r���7,J���J��+*?�`�S��&v79Si�1L*qBP�����Sŉ��N`��u�k��Tk�*��	��x���	L�a~�N��xf�6&�
�Ky-A��B�n��W�/ =�<�N�\>c�x?����}Z�l�u�w>��Vl����fAξ�5�`�S�",h�C��X#�7Bʨx0ͯx�����<-5�y[=}��`���NJ`et*�����w����`�!:���1dc�V3�Z��,d�� u�a蜂��za��"���[��b�(	�̸���quGo�N�λ:��g)�a#�X�^�:B�G	nlh�� �LEG$�l�1 >0,��۞5��I��8^�z4m���+^��iޯi�e"�Irō����u��٢j�v�y�ع�弄*:�e1��3B�Z��������*߽+t��Ya7ʶ'�����j�IU�[�l�a�A����<-�C+���[��A��4�m�714�ʧs�3�*��L�l�Ç��Gv�泰�b8�����{D�:�χ&�MG7�T3tZ���#���)o �y·�%p>���O߯�͏�`�y��,�\&�5B�\ŵ�&$��kH[�VO��&�Ɲ��1ݹxsL$V�ޣ��;�D�/^^-ɜp雕G�N�nnT�-�����x:��xk6�v������k��k�!HT�E�:�!Iަ �*-U��ڭ����D�]E������|FӅ��e���{�8�Ă��2i���S�1�)w��w�݇qh�<MX9���OÆ�g9s5+6V�?f�|RSx&�L|C`�?W=�0F>�|��T�x��h�*�7��Ç[�;���w���:�엒��T�`(OWA�����=��BSc���`2CEɵ'z��?s��N5�~o=�9^0F����C���@�x:P����J���]ny�![��[�D>nQ1�׮,+��,��jt�H{�-��4<to���A������Zvy���]t&Ek���Yq�7�B���ǕJ����#�E���yg�VO*��nߟ�}^�:9��W�Y��v�G�Ϫ:��G �;S$ÏR��P�G\�N2�d8y�Ub����Q�|�Vz������FLT�c����#��NlC�}J�F5��:"���l�$#��}�xn�b�43)����6��kY����HU�&@	�~�ԫ�E����+i��N����~W�뗧/�}9Z�J��q�(j��J����vɇ���#Y$�f���e�&nC��|�{Vˋ�����;���7t�E�s�(*Dy%W[V-ߟ�gJy,�ݘ��H�7��PV@��qx�);��]FܼHi� +��I��
�0lO[XRs�/��r�?yM6�uk�6i�^wMM1���`߷�6��jO��z��mN
u�-H��%W��s��C0�5w1K��*���(C���-��Mx,��e3��~�
�֠4P�i%H��FK���{��-0ot��cM`�rz��N!ڻ�m���}C�h�gb�pr:����u6��u֫naҝ8]�#�_�U���Au|���\>a�*�cc<��]��l������C=\s�K�'z]�OgfΏlP(2:� ��h�:��Gb�S=�+ً�E� �7��@���T;p��A�{�D�~9ipp��]ZzrQ��V��G��T��û��0+]�T��]*�]w�=������)r�:�zN�X;^ζ�"�Q�����RJ��ܱy]ħ3C�ث�q�"�!��v
Uϼ��ˀ���[���|q��]��x�Ú߶�8Fc�A�P��B�s�Z�����t]՚n�Tj��<
Pĉ�W���_
��uw��d]Q�/z���h+����B�I�Цo LX�S��ܭ�z�@XJΊ'EZܝZ'S.��<Խu� �����e�lଡN���q�P�rg�C3Q�b6Ud�qDN�
����fj�Y�0��L!YyV.]:�6��9�&2$NC $uϬk'jmK����0�pby�̼ɻȘ��d|��fY	e_d�Z�箝�+Ҩ�2�n�1;:"Ս�]��b��h�>LN��u�T5`����P{(�CN��\X�<U^�C2zFǠ��#"�ʶ�`lBz�7��0�;e��TF��$��Z@@������ݯC���l�Y�u�i�z�|CR���V@J��W��S6�L`�#�"�= �dVM��g P�F���v�	]-�^n�PWTmH~٨�7�F���Ak��!�A�(�5^��ɩ�3� WIb�瑳�W�n7�����{9��Rb�T1��r�TS���@�}5�pf4\N`���(�.�ƘB��)ɨb����Ә}�] f:BB�{��\]�ι�g�h���S�����ֽ�P��W��ٳ��	�׵�m`n��+����ծ�gWA�[Y��x�S�ӑm�d��~�+��t��ԅ<R�\x8w&���C�a�oR؊*uvD�;�ⅽ?E�����R���ߘ�bd0�N�W�j�m����
�����R��G.���[��+����2�kl]�Y�n�n&�Gݣ/�[�����raWs�v�oU잗�pV,�X	�^̳HEm�c����y�ұUw��N�}��)o.O��$ڻ���������T��	~Z�xp��\ٔ���E1�U
�W3y}y�L�O��B�;���o�D��6Tsd��YIOE+p}Рp���.�<����K˚�M@~��dINplڐF�1����Bt���z��îw6�n�H��1y�e�&����{�X���ע�Ղ���u�]��gc���'@�9��Af_:锛�m ����80Prpz_ۙ�좨GV.�I��p���'�8
��M�ZD��/^4�����,n�qB�>!}W� <�yB��|���������Kx,^C��B�w)]���k���͑�YOd����N+�E7���`����kW��"���{ĺ�yD�TGT���b�99�6p+��T��a�}�4��	�'��w�e�W8�&���P�2�s�:)�Ǧꈝ�b!��5��\]�aû�}��{���5\i�R
Gt�)��iIKq�4a�ƍ:��^^���qw��oN��'i��6�u*����ʄ�M�N��`�KRb���Wul�mp�㮊[��]0*7� ���9�O�#e�P��x��	���Ӭ�RM��P|1�z�%"}ᮆ_Q� ��ň�)37E��*�L��]#���+��8pO�ǘ}�5�U�J� �gՒ��.Xި�#iײ�+hw��K����i����=�Qb�'h���S'caQ�x[���c�9�M���J�����;^�j�bP���ܪ�Va�L���v��'�=����~>�w*�C�+�{Og��ճ*��ȸ�rq\	T�0;�|߯*���6r�+6Wg7���w]��7�k���u���rw��Ȣ�L�s���z�c�H����#7>#�j�RJÙ�X�"�,!�s�\���
|F*�.��E��p}/F��T:'�'8!�*�3�o��OWXH`�R"�V�z���:�ur�aa�?.��������1�"3w��0oEA���m������IV�.K�C����_�w̄�$}���ޞ��χw��3̉�|�
��XU�)}��<y`��Pu��a�:�O��G�;J\Tn$s�ϥ,%eO����)W��
�F^�m;�xIL^y�YV!�2e�:'g�CU)���+!Y������r6�J��)e�A�u� �]�y�-%�B�
s�,t���AM�u�w���'+C�
u
�5d�ڹ�d����z��B��:�k��±��+)@��ԟ=�J��H�u�7�,�;���j�ËG0ĝG��4�G9�.F�wCa�+����<�TPN(4�#�B��:3���e��,gW���ld�
rG�)ų^��ܸ�,�m3�1raǳ�� �KTK��o��r��=Ws&ƅ�7�)�����JLT�|v	�,G����}s��V˭���{���K�^�\Ш:`�I�g��Fe�A֬N����R<}��x�:��\�\�s��.�2�
��$ҟo��
6'���A��ʃ�M�=2���樎pn��y��!P�����LP5#�zo��"�lT�Ub��Np��X'���������L��юv鹋�g`���yF��G�@�ujE#�0���iwj�7��adRL���lֈ�� ��Q»�v����F��[;S�����+�ך�nxy��IiW��!��6+44�.��1T9 l��!�ʱ���5ae�������3e2n������(���K1F3L��,�ǓKy˗sz��Q�ғѽ�U�	�m٨[ܝ2-XR�|��k��'={Huc��{�� z޲_3��BF�:uP���.-��*Fvc�m�I�Ű.̓P?A�Ӥ����{�q��tm/r<�^Pp�����q^o,r�q<Z#Y�+��3ʕ�yw���?8,&�@�}N��n�X��o�PAt|Ͻ��a�*����S����|J%�j��;����uk`k��髓z�F�j u��]/wF�j:N{�����-r�U~Iį�w���'���踮Șe4t�׬�a������0
�]lK�����c�x�� Zl��J�vЗ�ĺAq��q���c<��wp�X�z��RK88e�b�v_v�z���v�]Z�����0��g��^.����*��A�k(�7��>|�FV3ën�:����NU���4\17�e1�:Ͳ����eOo�� �����,��,r^�A�3�^���,˗]j�w7���xZ3�s��[�ھ�j�VjfZn�����zZ)*&)�$�xZ����$pYX�r28mӍ�B�A��ZN�X�y��Um,���`����Jժ�ж�Ј.]�]���/�K�
2[�p��w�������Ɨu��$v��X��
"�O�N�8����nX��$��C�3!GG��u���9e���6ڰ?u1�� �����@�a��e�I^�M�LU����tf\�I���΋�&=Ս�ke�{��=�s}�:'d��%T�7�	_u=�w�g�b���>�)axM�;@��a��]3�j7#h:��J��$�HNoZ�Ԋ���/7V.S53�5i	V��yӆ^�Iɓ��j+���ܭ֑����m��\�H+Ԋ8�we������L����Ǟ/��vm���TƂ�cmas8R�ՔI�V)�u���!�V	�M����z�.�)e�3~�;h��M'e�F�QB�zuKh/���g����(����)���
�������K���s٫׏�����|�Ӗ���^����7'���4��8'��7sJպ]d:gcd�e�q��4xkK]�U�}��g�����W=�J��փ%� ;H�'o��_vN��w�gJV�?w������l>�!|C@)��OT<N`m��Ҷ���]�`�j^��ݸ#!�[;F��u����:��oU�mIgu�;I�.��ˊ�j<':��N7�WV�D��]Nv�<�s�E#�
^'ȫ&��O�Q��{Hf<���:,�v<��1���m,�Q�Q�|;x(�s;�ըBJ�m/L���m���;/S4n���<���U�zM�v�q ��F����]7R �},��vBt\�UK�4,	��դ;[
�䕞%[6L\���9�}�������V*9V�ڪ,T��,PX�e��X#E�Ե*)R����)L�3-H������m���RR��*R�TV6�f3��-#j��ʢ�KAk+J؈�̦�l��"���+XV4�0��C�ȋ����1b��U���R�S��-Ab�b�UP�1�Jւ�e0�bŖ����	mJ*8�1m��YUR��dĪ#mUm��QR��aiTKe���c
��-�f4*++QJ�E����Ebe����b��ڃ%�Aj�cQ-�V�kdQUc����E��mEUX�DDH�����
�VJ0��TX��"��QDUX�-�[h�$AEQ�m�*ȰUF
��+lkU(
1V*�jYm"��k-��F*����X�ԕ#V�UAETU�le[mP�F-��D�+-�ԫ"�mBѢ�TF�caZ�X����D�e��Җ�b��UhQ�kQ���Vэj"������n������Ɛ�ۍ�����{��/�����QW�O����-��u͸�v�=���='B�ݖ��ڷS���������f4G�|��cHpC!�|bB
k6������$+Wb�������$"�\�]J偵]z�w�P@����[g����)-�}ipC�ui�g	(�z�f�.��������mr��Xr;d �uN������Uт/Ԫ�������k�ˢ�	`�P�Q��^NH룮S��/Ob�uN:��9X×~�����i�A�������6�1x���^����jC�&��}�5��P��o�#eVxK� -�gZ�1���'IŪA��aѳ*E`�] �d��9띀UVCJ�Ϙ�Nԡ����y'4���8k��^��[{^����`�B7�-�S+�<9�����O{e�*[�֛��՝M��xF䌊ʃ���`�<�P�v$�p�� ^2��OV�C3��4[��X��Z�Ӭ��0�@��#��9��ʯED��i'f��  UC�?;+����&Σeٳ��O�uv�F���XS\��1s~j�0T�l��L/�+���ɗD�s
�/�m��%i�e��2�L����u��Ep�5:�B
�=n\͎akG(���^'��`9�GV�j��.Ή���2�^���}�����N�	<�dsB��YY�9�C��]�,�.錏�N!�d��iA8k�ڧ��^�{�(�5pvA5͍�0�����������RC�S��s���5e 
�L��;I��F쿡�WЅ�
�������U�)�	�X������ʅ���Z��!4�����c,�.�D�R?-�u�x�Y�}p�8���l��j-M;m���
%�F
Ǹo=�w�Ɵ��k:�Tq�>��(�4�����r���R}�V']�lQ[
��>wO�k�Ī�0��LZ�7���e`Oy��ȍ����fC��-_�t66�踜U�9�T���O�8P8�Jd�>0eF���x8cX��;�}��[����e���W��n�,d���f:-b�ܸ'<���\_3�^Ǭ���ռ%�ˡ�(���8���a�h���m�.d�7�H�J�"C�r�����G���Tҕ���D]T"\�H�u&��=x)�;kδ,�d��|�T�Du�X3����7x����\QT C�#LB�d2P��Q�l��h�z�lOE�l�n���O�����i%�ι��0Y٥\��.7���e5��<��
�~`[���E��"#����W��7K{�Y�e:��6�L1^�v�Js�x3D�Xz�v!ۇ�h�kX��{�djS�q,$���n���T;	9�D��V��(�����T�g�Bj](��?)wJ�?�U~�xp a�P�R���*�8��b�s3d�����ܪ�ͦ.v���#��H��j ���WXC��`��dcjL�C7ޏ^�Q��u�=��ؤF�eX��$U7!�:07V�WN(���WӰ*�P�f��*��s���L�giE�*pC�S����ަ!o�C��j$	�L=��7}�_"���?Dd��1ꤞ���gvs�Ӟ:B�YT����8Hw�P{�m��i�u-��ú�z��gUʺ�W����X���m;��>�2�Y%����8�,d�l��{�x�g,_z��S��*Ӫ��_��g���ĻIgZ��>��S�1�1M��K�pq�g`u��x�zw/F ����r�K��Y(�J]o��o�u������YF��;[���HU�#=�L|.��eW��d}���p$m!Ne(�nk�2���'��OةL��_rQ�'�q��^���u�)�}'����*,*��v1�z�`��7Qr6���*����ΌV�SdB�#����27�ܖA��N$]u���A�`c;C�_iv����r�By%�p��7�} z��I�v�]Wj�;�$mY}��ѯ�3����U��~��tay����AT&Z<n	C��Z�\��V�\::����w���uu��S�7B�| ;�>���s}���t���K�ш:�ʖ'����~���624z��Ywb�e>p|�����
��sсiݧ��{N����2��~����%�8��rd#頙�.,
q\!L���K�R��G�r������%,B%�={�51k�^ˇ����R���G��t�������>+���*�Q�L�5����%xًj`��8�m�w��S24,��'.�@{�-����]tFLT�̚�ofa����L���B�Y��h(>�Y	N\����áJ��g�7�B���ǈF�P!8!�Q�d˖�s�J��4�|��Vb���8Ϭ�K���xFkӓ�ܸ�,�a�v�'0����\(rvu{�;z��"<dɃ�M3|�X�Ǐ�m�&*[�q�3��x��73���qf����<!��VDQ�V�"�a�̌2�Y@�\T_A�m;�F�@B9�@3o\����u+#tE�:��;�C\)�w��BM7[����
6'��Z��~^��j����2��'��������sFU h��qv�%@{NS@��˹i�8l�{��<��{1���f����YN�IR��ȳp���ī��3}4�`�1yod$N�.7t�}x��o���N��'L���ȬE.�a�J�}u���2T/:"�� d��n*Y�����l��وu�J���c��I�=U�ԑN��9Ä�
�4��o�g�rg�)��������a�#n�����+�8�ɨ69��!�8����t1{M�����D؜4��e��6k�S���^.ߕ�C�7Ddl`}C�h�l�U$��k����dgf+�wq�C����J�>$Ld�44�\!C��Q��Uc���f��F��e=7��z+�vϊ|�8'xG�/s�ճ���W�퐂��6j��M^ݑ��KN����̱U&���rZ(��Ѓ�xs��x-�XY��~��7�J��e��v$����m8R�R٪�r2�;Z��Sw�/��퐮�!8G��J)J��c˔b`�s��g��ý^�o#a���y��|%�C���b������ˬ�v("����z/�\�\OS�($#/d�@z���a�	=�}���VN�Ǉ�A�󏕟/v��Y��>q�_���-�9�?22B�+���@�U��.u�\����BG\����'eb2�����o%�����&���&�a>+�v�L�1��6@�0S���� Į��Ź�8�TͲ�
�08��z�l�mTP*21��F�*}(.سz�{��,�ϔ�d�N��-ÛY;*�w'�j����Q��y�.1�B�࿕��c�� ��\$[ƥeb�0ב�D�"�yz_p��<���[�:"����!��b0Tp(d;�¢��2��	�6��Q��&[x��U�:"vX���;�&pE�g`3>�T@\��I'f��  C�?z:�d����Ǎ��J��/�n]�DSunb+� �B�.m���S��2�l"��(e�'ll�}�s�_bC�RɨnlnQ�,uD:Z�"�d��SG�D�ͣ�p^U�W�z����G0ϩ%�pU�v`�q�x�Du��xz�k���^(?^Ӣ�Ѹ8x�YfHLm���+��ڬ���8Df����dti��E�Bc(A�Q�8�p���4�ڤ��9\Y���N�/Np#������(ԟR��'ll�Rܠ石d�ADnM�n4ɣw�q@˃s�3�D�v?�?l�J�o�_�����Q��D�7چ;T�WT��Q+ؠ���b�:�j �6����.x�tw�qVl��P:�!�
P{&�O�ƈA�\}�BsP��^d�g���W1�s+��	��k��4��2�F�1�b̥��q��p�5���9kk
]SP�MY��l��ݾ�G��.o�72W�'yx��{n/r�o&����krY�o�wNo�y-�>�4BݗhΝҶ��<%L�i����Mk��+B�n'#�{Q��6���}���e�A��^	���ڰ�(��p}֗m	���������b�/_���||\�mH j�x��:Qn\�ږ ��Y�'W6��v`Q,m�XWH� ϥG��mV�.�i��o��xԷ� ����{Ky;��RMnv%S�"���,'�B�U�1��y�[�\�j��VO�h�zǇ�>8�c�:�����E�l���3x���a3���pB���Su�L���eFW�}�ygo\D&�C��O`=R�r8�;��@�� ���H�
Ѩ���Y8��$FK���x�a����^4纽C{N�߄�R��b�}]���0���6ӊ*D륋7�\�UZW�9����uG��$`�MǦ#�EV�bćs|�P�,��WM��⒆��Fߑ�.^�az�:!�W��^W]b��64MB���TX��u���;y���ۗ�Ɵ�(Wp$T�#��%�0�li�V6/����PB(d�,Y��6wr-�Sn��K�WZt_Y�lLL�ty0��O��V�Ҷ��R���E=��`�\�'����� A���=#� �U\�찼��:�^FNʰի�j�M��F i��V���%�v��B~���ϸ��Ss�����𻫾֦j�Θ���)׈�f6h�"�ע&-��L�?��f�-�n+��7'۹��A>��2����{����ò���*��U�TxS$���8O�5ء�5�Z8��]s��@޽����c3����eܻ�8��s'#~B�]ן2�f���t��,���x�Xbmd,�2�tco&�@�b:��QN�1 �QP�C����ꕏ���e���-�d��=ꛜ�?j#G�?�/�:囚�6���B���}��8#��\ackS1���h������Y9 �S��U��
&#n�@�q�&z��<PG�b�{��P��5��OA����Sw{jB�@�b_��B>�L�>x-����.�.K�G�r���^�a�������Y���s���V��ê�]
����)|��mE�@�W	�)�3��O,?2t���t�B�����]�li�aX��,���Ժ�
\`CM_��;}&�h9���#�d��,�>u%U�յc�7P�ҕ`�v�͛ڡ~�pc�iE{��Wl�����T~M�m���#������c㙼9�'@J���c8Nv�8���$*�� �e	�3�!�t�:�Ћ����TLhS�S��{�1��肋�C���@o��v��Jx���7�ˢ�V�#�y����`�Jv+�x  ���z�<ɻ��~�24���V�����UY�Wk�y�����	G���x����2�/�ޡ�g5��U0|�Ĉ�x�{i�fo*W1��6����ox��U}	����%�oU�zH�������P�$���jŻ��A͝)�^��ڞY������D���@��%368T ��$�u����bz������p�WtN1bwi�r��PWV���S�9=�����i:m1@Ԙ��q[S��`Z��=�̘]o�m{�=2�ب=u�u\�sh�v鹋3�
�	׭�(=��{�*�^�]x�Rz�G�'4+ŭ�HDm�7����^�O�>� ��Q��C�茍�}C�h"f��\9}T����(�.�`v��|�MP���"b�%�e���a����H��z�wkR��K��}�v+��O���������%C�w8�l������d���ݪAOP*~�0u�A��=R=��8����T`o_u��ѭ�ɯi��z��x!QH)���C�����5���JŘ�3���ZM!_���M�(�y�+'��1'=�ta���'���|¡�N��k��z`���b~v��̻�+�{/��v2<������E/�z�Q8RyK�zn%�Q0w��:%'w��;oո��Byà��	s�N�M8����`��S�|��(��]e��-nh�E�W��	F��I��	����G���pҁ�p-�����{�o��p�5������Sl?��4�h}�N��+�B���6s�甂�&v�]���O��E>d��������w��>��*c8�*�9�L�2�����p眺��������!��z�l�d�a�
�Ϩ9b���ԟ~�@QN�|�׈I�>O3����a�o��m������u���5�S�� ��h�1����\n���q�|�e1���e��j�H~���~k+?!��V�mJ�o�ӈu@�.�8�gW�v�Cԕ�w�M (��{�|q~g3�Y�O3XB�����Ǯ=�f�J�s|n�^91��_�r�����6�SL:g�UR
q�u� ���gh ���ÙH,�^a�>B����0����C�yd��JśN>M��C�I�Xn�ǻ��� #�l$�����y��z0�>���ÈVauE��l8¡���Y�J���
����S��Ri%Cyd��ܚ�!Xx���Z'�s)?*O�$�TX!��P:=��-���%������^f��1 �������Xx����i��J����H�~eM"����B�c-�9�+&�q�Cg� �œ�gY�PPS�L��6�@�4�0/6�����0g��k+/�Y�*����X|�I�Y?2��W�Me;�a? Q4g�Vm ����!��z�T>�݁������4�`cR�氬*~C�bM���a�E�@�&�́�=1����Uw��b���y�錘����I�� bM�l�>d�;�<��aY�NwXy�2�T�>�UH)��d�u�8��w��!_PY��o��� ���ئ�P�� >B<z6�{����sy������<Oǻ�3�%b�<�i!�I��f�d����0���1���1��^QO�Ri�aP�4s�N�k�I6�m�O�P1<`S�Co&7�����X�9�y|"<�8��˪O�~�C�ֵ>I�?%E��Y1=d��<�� �@��������d�VqRVh��d�*u�����
���9�Vu�i�RI��vg9�ߏ�Ә��;�G�j�F;>�¡��p��;�b�z`�w�$��9E��9�|5���"�&�9�7��Jn�VU���뚫�����;̜W8+��X	W�Ɉ��d]hV-w{Xd���K�khj�X,Y�E;�Q�)� s�u�H�M��J=��I��;�X��G��٪��y��x(+��p_+��F)��]f��{�;)e�lFF�֖h�!����:��*��t�E9�!�4���ˣjme]e$��j�l�ᰲ�JݘT�{"�y.Q�lAE���V�sV��D0*W[�7�3w�L��v|�*Vހ4�,����+^����-S]"5�MA�����\?:皻��2�y��8��"[GzAwW�����c:����	},Y����0�Z�S:�.�vrK#q�M
�θ�!��n�<��l��R1�d��30sv��~M��c:����)e�JɊ��C���*
=����.Ȕ�b$�����v�mڌ��Bɔ��r�{�B�-�B!�+9Lg(�Ҏ*V�QY�9�+7a�T:-��-��p���X1�V�S1��f���D�9�nVƀ�a��)L�{٤���S�6�]�f�|��Z,wT�х�h�H�>�Cy4r�)��w�W^|wz8�HMTC��Hs>�+�������f(�[i���=)s���-�������Z}��������ޛ���[��n͗�(aZ8i���}�iVk�c�/vTv�e��гf�+2�Ɓ�{}*.�������B�ݯ=49�eXK&z�o#�P�[x�����"�PQ�h�q�7V�*�]�v� ��s �5pࠚY���L�Q]T���p�����y���!��
f7?�'���#o���g� ��oBl����8d8��W�_F�P|~SQ���������h�ɲu�%�o3Q(�z�~nɤ,r s��\r���f��r�N�8�	�S�p��(S��A���z��C ��Z0��<"<]���*�]��O>-�0�Y4c�U�M��fY
��[�s;Zr�'`Y��+ݝ�Pf��ҥ!u1q�<-��|�vg]�TU�4
�}���5n���v�J���I�w��Ih���g"I|���7Q�T�s�^L�5u�Q�¦��Y�ŉ�tkQ�X�Շ�;.�xHQr�[�V�V�6;0��nC�6���!Vd�q}�:�6Rns�L���n�p�"��=�pn�k�j�#)m�Q�x�wɔ��$�+���oC���$�Mމ�i��b�L������Dl�1"��z�i�1u�� �x�J�I3j�m��?M7�c�x�aȕ�z��7�i�z�H�9@^-=�֌�Գ��7s(t�%]��7v��L�X3��L'Zeľ�ɝcF��
��`\��$�������O�w:��=�������R)�A�"�D�X��QX�"��E��(Ԩ��*#QEV��1*B���!Z(�mQVT����Tb���Db��kUDdb�V��R(�EKE�eB�U+TF[U�EDEPbZ��QTPQF*+*�X���E�������"Q��
��,m���j�b�b���kD-�V��m��h��Q�� ��DEX�V*"�DA�DDE��[mk,DAb��"+�TPT+cҨ��-*�
-��**�QQX�
F#J�����ň��D��DX���6�H�(�`�ʱ��l� �Kh�h�X�Q��R�TUbZ�+TD�UTTD�Q�F)"�cZ�R�EOi�V ��h�S-L�DDX�X��(X�� �A��+E`�,X�A�UTƱTV

�#�#EH��a�2*��UV&�Z�毞|�{��x���{j��s�q�+z���$S�2L�<�Eo�v�9$��]�0�Uw�t�)&*[����E�$�p�x{�M�������!���i��&�SN}�v��R~Ca��ь�9�B��ܟ0��'��Xi�g̕����Ф��)8���=��;�*"���Ʋ��|�}6s[�9��ߺ��������=�6ΰ�=C��㙄|���f�;CI�a��8�2b�}��T�v�޹��m�2{��=ݚa��f�7�{��,�%O=��D@��W��ɪ��}�mg��<�����qiR���&tw�<�Af��{�q<C��������m>Of��H?Y+\�<a������3��LI滆�a�=Փɻ��!Xm��?{��?���5�=�@��T:{�'�������^�?Ou��
�h}���̇��ԅa�s�C����@��a�q'I����tCI�&�f��
�
�~��R��O�G�����{뽸��D���SÐ�Y�n��Vz�+�Y1OS�l�0�I�+&��M[:Ɍ>C�8�i�>�xɤ�6�_�'N�&ӌ���!�c���}d�~՜��ޘ0ڗ�WL:�ǪX<V?MH���0�OU� �s���x�Vc'�`m���<��X�Ĭ�N��1����Xq�"��0Ć���{̛z�Ɉ���!ĕ��&vI�3�ԫ���Qw�� �x�W�[��+1�~�~�,�'�������9�T����dՆr���,���m!��g���h~B��&옛a�b����m �d�|���-W��7����7�������u��Y1'{��Xm�Mv��I�+!�wX�(�T��p�?n�g;a�_=�)�
�Hh�kR~e�!Y���0��>C�Iئ~���ڠ�,�|G����щ8��v�=B�P��6�a�1'y���<J�+';�@Qd�T�����T=fJ�l�Ɍ8��I��浩�J�����4�	t����O5�XbN�����8 Lxt�T1=d���>La�
�ɴ��c>d�S;a���ӝ�ؓ�e@�����
��� sv����p�mE'=�����bx�X���ΦXn��6��)������#r�m)rG��Iw-������Fσ��'�M�~r�p�~M��XZ�{M�ey��{O�T���������9��U윅]!�!�<�s#-�!���P��0�U8tKr�P[�6p�+�͋�VU�t�_�{�xxT��'m���A�a��=̝aR�73�&������j�����l�xJ�gY7��Ϩa�
ͦ�k!��Y�^��J��~�@�x�͸�\���	� Db�?i����T��n��U^��S�C�@��c6���=B��Ձ�Xx�CS��H:�l�Ym:�=�Ru
��ɉ�iXc
��>��J�a����M��a�	�U�W�>�#�SsV���B_��������AAE�:ŏ��
�����~e�!_5����'�s,�nɌ���6{�4�ALd����� ���ɴ�����H�IY�eb��������~�������z�����=E%I�*w߲fퟙ1��¤��~�,�J�����F2~q:�Y�kY?!������~7a��W�&�}ÞR?2W��7�)4�=�hI�#��T����ۭ��wg.����߁�i凪�H[`|ײ����4����y�봬��Hm���� �a�7;�QeaR�׽¤��4Ɍ75ܚE�+���ٴ������t�������V���7�f��O��������z��CI��Uԩ�
�Ag\~偞��8s��u<Hn�>Ь����3I<a�����S�6�P���f�c&r�5I��n���b��9s�>�ߺs�_��@Qa�7��|�a�w���P+����w-`_��>d�

/g7�m<@�7���yd�����0�X}��Cy|=̀��Lqr�1��� ����{X������WSy�z`ǅ�
���/��0�v�n��J�χ����&��&����>C�u�q���LM�����u�l��ݜd���N�x�z�N�D�O��1N}seD}�ح=�d�|���{��b�Wt�XT�)�0��4�&�A}3��Ğ�*����,8�y�H~���2��b�z����1:Ͽ^����SÝ��,�	����>��__�vO�����S˕��@�x��c?e�"����:�CĜB�L7�p���8¾k0��{� ����x����P����Y�;� �HW[��&�Z�1�a�* Q�����U�d�_)ٮ�Mq�X��~�|��������l��mwV�r3�UDd�|�HWM4u�ʜ��P�Gr�-]�%,T�����Z{ݾ�f�d�ob�R�p�� Z��3i��I^�I���X���6o���ç�>���Msـ@��O�����~��5w����������AO�|�ß��:�C���rb��1��܇ۤ�
���&�a���u
��]°��P+y�j
$�-d��q���_&��O�+?i����I��Yо���x���1�RN�P�s):�'/wH,�N8��d:�H)�o��>|`��d��rk�k�=����ց���}�Ri ����Y���'_s&�>e�~d��{��M%��]	���
���:=�3��O�Sv2z� l@�'��x��$�'���R��3��6�k�2|�b������{�RO�>3��0I|g�����w��������B����֥g�13T8���=�d4�: l���RW��L�y�1�+��2)?!Y�g(o}���s��l������ì�6�U��˛��?}���A���`>����f�AgɉZy�2��1~�i ��=���C��$�Y��M��=�'P�����f�ϰ���1'P���gۿg����c����CL?}E���a�C�Me�<��Vu����k8���
������/hi&0�<�M�C��i''��i:�H)�œ��*����Q���$�=��>�f��}������ĆZ��{�N*J�Y����bx�J�g��2z�l��wu�I�wu�?e�d��ֲM'��8�CٺI�=d��]�+0��ϲO�G�G�i�����}s&�D�_�l|ɤ�N�f%@�N*~q �C�O?}������:镞!���,��J�a���Că�>�+"ΰ�?\�k(z��'Xzn�H(z�����ca�Q�|w3���@ ���Vw��o�!Xm��3L����J�d��`T�8���4ξ$�<��M�AgɌ';���a���~�IR
i��w
͡�4�2~�s��B9�����z��}�{.}�D{ x�����+;矵&��k!���I�=?SL6��w���4�Rw-O�$�?2T�ϰ4��SL���&��,�e�=��l=a���{�׿p��7+���A�u��s����ǛyQ�- ~���l�gg����Fe�9���[���:���+N�9R��~Ҏ��Wd��޷�R]Ų�{�"�ݔy���Ĺ�^�lk����y�g;�❻����=ؖlr��_���xY8�[,M$�	�&�x,��+Rx���0���.����=�m1��d1!�{<�g%@S~�I�T�)+=g�1���γ�`x��'S��n������{��*t�o�(�y-P�Y���{����p�I�
�Cg9�����>C����<Mj�Sz����2y�Pĕ=@�N?�3&��Cfu�qP�m7퓎�Y�1��Y��8Ԭ�7���W���������ߞ�S�=COu���"��+=>�I��~I]'���p<@QCѾa�1'�+�;�d���C�w8�l�����t1�d�����1H)����g]��?��}�ɜ;��C\�_Dt�Q������a����u
�AG�2f��>C}���X��99�<H}i4�|�/,�@Qg�����h����m���'�]0��Cĝ���r�S�YV�������W�ǔ{� d�(�0*|ó�4�hw,���+�!Xm�2�9��s�Ag�]���O�����ȧ̟�`�C��h��I��9�/,6���xk�*i�T��U�Ĝ�y�F��k�����(��=06%zjèi��[g���a�'���:�?[8���H
)�O�w��I>B��ya�2��>N�f�̞'ڰ9�f��J�ɬ��(>@�9���Rﮭ��C��9��8���:�7>
!�5�����c1�E���g���N��1�i�Xq�"�0���z��J�;�2M�(��h������>g�s+:��kV�Ӈ�w�[���v�`�ZL
��(��M��&��J�a�������{����$S�]�6���Ɍ<Շ5H,��a�>B�����l:�C�ug��L�d�Y��4���u.~��5��y�y��t�7}�����L@Q{=��m?j��y9�u
�l.����`m�T4�|�]����%M��*
/�N&$ĕe��ɮR��</u�|�2�S��R~t��Qa����8c����?}]�r��4��t7M$��l�ڇ9a�C�g��C��?*J����H�~eM"��5���VLe�A��Y6Ì*>�T��γ�((
)�&��N T�B�;�?�r�]O�V�ײ�9"��V�7�eBM+�]s������O`�X'�n���=�b��T_m=A�gM�H�ef�Wt���ݮ��3�����&y^&y�{�K<��
�!���<7��bM\�s�<#8��$S��8�$���-B������x��Dݾne�u���q״�C�?U�?�6�Փ��c+%zɼ�ϳ)���ϰ:��A凗����B�y>�݁���������R���C|kX݃c Dy�s��Z7O���y�������y�տ~�hi%_���P�p�v�m��4βy��]0�+4���;@�VJ�gܳJ�8�мɤ�<q!�e���L�w���}r<"=�1��[�9l7K�w����b��Ш�[E1���6�!�f���X��)�Hj�z���g�i�N�������4�l/(��Ri�aP�5��;�
�$�{�AAE��S���߸��~w�������k��@�O�k,;��YHVM��d���e!�kS�8��TY�Փ�O\a�38�H>�7�������l�J�*J�{a��u�:��*�{`	�y��Mt�N��ɫ��z��g���ܻ��&0�
��rA�!��?r�H
)�=��+��
������O�Y!Sf���~d�;�0�����}�Ф�g�0�VT�ힲtσ��&��쒦j�{���3c��gz�Mef�~�h
,���l��?!�v�;���"�;�$7hi�ݺq<d����RiۤCf���m�2{��=ݚa��f�6y���8���D|8�U"��q�+l1L׿gI�U ����'�,��Oi��
��L�;�e �_��P�x��*)?r�&�z�Ci�3�����y�0S�H{hy9�*g�����~�`Dx\xL3�E�oGϕN��|�����q
���t���u�Cϩ;�X�C��i�{�? T�C짟y������<���Rz��zs3�8�M%G��O�4�ҿ@�:G�a_`s�S��WZID�:���~��M{�n��V~T��J�&�S��y�M$�
ɿ;�Vβc���N �C�O�׌�@QN�|�_�'C�ɴ�'�;H{��>a]�x��>��9۪ߔvG}�.��ۚ�n~��ɦq��C��仢�S�ϰ�O�� ��,�a�Y�j����͞wh
,o����N��1�����E>�x�I�����H}�T���s���/s�h�<�
���uhtڡ��j^f�O���E��)���^��2f�X'�-�b]�x������n����4[I�'}����Œ��]��'e�OZΪ�g3�*��(
��V  _M�7�d��(�l�`�$?ʯ��<&h�o8rM���zaF��*����&��,>aY�~���0��2xk������9�T����sV�B� �p��6����)�&���E�옛a�b���������	��`��w�LZ���>��L�cH~��{�C�m��Ɉy��iaS]��ɴ�B��P+0��iR~լ
�&v�H((�2|e�I��$���B��B���W3�?v��=���=p�'g�1��qĝK�T���?8���
�~�����<a�1'���P6��VNw6��Ɍ���pRi'P�l�d���̘É�k̛I��?X�����6�r�a
�d��z`!l�8� V=���q�P<�SL>a_�<Nk���|�^�滐��)>C���lI겠o�����j�|���4�W|��(���C;���3�����+;=�Q1�!PQ�:n� �Xbk���!�Cf{����&2yj���� l=��Y�M�p�|³I�a��Y���I��U ���:����q��q�}��V��g�����	� Da�0i!�@��a�x���?!Qq�R��1f�a�6�udߚȳi��ߵ�N�Y�Y1<��,1�N�Ϙi%B�����M��a����ys��������~zt6�쵁Y�Ϝ�H((���̆Ө'��7�ݓ�/i
�P�ۤ�e���1��~q&�{��H)�����`�B�]��M��w����G(J�+?~��j�����ߛ��y��_�:~Q�ꌝ��X��*}�G�Ka�U5�]�����M��잗���t*�A����[��R��1�F���Q�"���+je��/|N�f>�W��U�kU�Qѵ�F�L|������w/F ���4ɺ�u��
d��q��_��|Ml��W�Ȩ0r�R�z�
2����Lz���"��j�b��P[��W�VԮ8`��a�����Y��C�0�w��nOy �q�y�V�o]��o]c�7�M�juo��4^������+"��T��tu�������{vP�/c��7�	��P���f��|�ڎF�	�7�6g�� �Yi�P�ؿc�FA���(ñ�^�]*>��x����>��Y�e�ʌז�$��#(=���`����R��\IQr4�����|F� u�>���-T9���Y�{a=�����d�E:�����p��:P�L���
.�;(+|�������V����w/b�ƫr�G�aJ�ѩ���]H�l�sr��c��Wy�>���Ml"�.B}��nPf���opyUdI��~��;m�ߺ\{�z�An��<�z*
��8���X*�*;���],1Yy7lM8����{*č�r���#�Ņ~A܇ָR�뼼��L��/<q���]�]ح���N���O�H5WV�!��\����êWn;f��g�JO�;��֣ʕނZdt��T�w�,�@���v�'�?���u�u��]9����D� ԥ�V��c��$�}2`�|в��Γ��>��\6��1Z	X�5�dc}�i�B�q���!�{哎o��Rtݡ0���ή������T�L�HH�;$2a�u�!�1<[&�<P6�|��g7 Ī�&�ƻ�&p�\|���-��TI;��p۫N��_��t�ٹ ��.��YP�E��U_}��Q�����Q3��=�,@	���dEw�:���\=mX�W���Z�]��Ǝb}��T��­�f 1^����D'Qr=��d�p"g �֋K�W���H�[��c�c6ʃ�M�{� ǈ�T;)�7�6I�>?����Ω%��9~�<`���22(�}s-�h�0��nb�l���Q��y5F��=����'[���e���s��9���m���Q��p��Qp���y��ds�}�5�u�Z��l1�Cfh��آ����iV|����#b��*�����>��yˎwt��O3S&�ڱQ�!q���V�z<o=>*�3	�����MT(�۟lE����s�3u=��)�)��
U'�}	�󫋱p_vd����[�|@��+f�D�6����-��nw�6�EZ�Q{/�U�EϺ;&�wD���jD$7}Ñ�!\*R�vKV��R����'��ζj���j�@n��g�+�O>���(w���{<�#G�}����䲊v����-,��f���୬�Զ��h�׀���D��H��k`�d��Ώ��}����c�j�5v�-��}�vX��6�Fs�s�Q16�N�WRXg3��-�����gaoj�Y$��f����:�ʪ����;�c��#"P�}���<!߅"�6n�� �nr
������#�G&{�J�����n����N5-A�����ï=A�Wg[5��/=�'�+��E`^9�
}RƪV��ʟ-�x�7
nV��;s���g?�>	�x0<��$"��E�딅��kp���,�mƨ�Q�9TN)�2k����`�hlPRLFx#A���@�y2�Z�v����6�19�s"��zTp��]혆d��l�(,�&pE��;f�И�U�];�r������S�l5~H��(�62�ʱ�Mչ����1su��j�;����7����\����/���]</�ٱJNhW��W��=�>|t\P����>^%�r�R��L�,:�UK{C0{�}X,���< tѻ.n7�%:����.�8ͽ�t�&��k��~���jp���Ҁ�[~�X�Ǿ�����$~F�+��+�����2�s��'݉P����������6w�E�"ٸ������\Q�4���m`q1VEw����DKg���`_Th'm�>~�~�bm��C�Bc2��N�����1c�bvo�*��(@k����F�'����,yj�!d*��I�_6;�ޑ�w���.-�1!ܨ)��ɖ�gW ����Y����aǦ!v����ii�#���-S��c� ���ʹ�`�iT|0�FV�$w�����a�:�3�)�g25b�����.1t�g`�5iJa���de?�X��w�
R�f[�X����S�)��2�xL� =���d���u�ΰEg���vb�82��5�Э��x��!ګ̀��%l���g�8�ncM��7ݣ���
*`c��6�����+���긂-�QU
[�ٵ#T�m.�ٛO-rJQ��4)9�fG\�*a*�(@؞��9�3 "%G�R���z)ǯ+ރ��OQ�rܹy����Li+��&v/ؙʛN��aS���@��4�+�d(��aZ35C���x!GQޅoJS�\�K�F��xWg����®�?�^�KÀ2����Na
��b��"3����`utu��s�ϩ���ɑ�K�"5Z4�jlt��ֆ��ys=���,/��B��Bʨt0�6�ƪ��`y�MZ���;��7d���X7LL���QW��i�UšV��w��b��DB��(E)�੿G�#�E?�!�×fm\�_x.x��o�&��ٽ��mm�v�<g��Hh��3���E�u��Uks�ɜ
�9�D6�����B����gbr����Y�c<1px|��� �~*'L�|��BI�q,��m�c�o�n�zLp�/^tq�3p'��u�_��y�r��k���R�c�',�{����R5D�_1r�ݑ,F����,�#a~k8xN�/`�6 "v9���'����k�	�"��L�7-��&b[�]�)�wkMX���E6�[/�ݘ�(� ��-��pk4��-��*���{}�$4�gb�x�DOax�����ꝭW�K��]ek�ϳ�8��Uq����A���{q�l�RwU�s�B$��y�ld������d���w]Z��K7Iu�������7F�zzc�Nxb����j�C�q����s��P�.��A�[���{�u�,���o�����\��8��m�G^\u{b�r��͒�}�z��t����>��A�ت�!j��ѥ#:�/�O����F]��-^6��:�K@�d�.�3rγ��[�
��m��(�S_$y�:�B��,�̫�)�����-�hY�{E5@b��ty���d�f��s��*�௵��ci=�a��E��Cl��I�PC�*s�vkbј�m��Zn��Oj�ք$�QM�����	HB�Yvo�0����:�w?����$���r<�zʖ����8����A�� ��]�^o��Vq�6�F]�o+�x�&Е��tΰ/���Aw&�lf���&8]�@�\����17�@9;���f��� ���L
��-�40�"z���u�H�r��L�([�=�%A�xXu~��:C�ne��Qݛ{:�&��ړ��<Suuj[���x塝N,���2`A�g;hR�>(l��w���ZI[G���:��nU9CL+[�RA�Y:�;��#��ݱ��î�O)U�^�:��:��L��y�ކ��h���������?�C�;�ˉ��R�C��*H�����aS�}˧��,�|!�4�EC�to�ss/l�"��p�*�&3%���iUy	�f�k��Ź�ux�~X�"$�8w�r����c�z���[�r��>�"��,�K���u!��׼���\ѳ��e^eDO�.�M����ν켌��ǝ�4�^2�w�XB�=�_Z_U7s�o:;|�Ҩ�[��
�~�2p$�s�Ps���f(���ղ](��e���8�J.�W]
�7.v(�$�X"������9�$��s^�):��3Ax��9��ur}B��y�e��$Ḥ̂x�h����J��og�P���iL<�)?��GpC�� Wx' �
pSLЭo	�@{��Qޓ�݈��N-��n;�mvM�D�oZW\ ��z�k5��W�LT��w��A<��z�S���դl��wiN7��w�_� AAQEPU���("��U���0�YR�YQTTQ����QX9h��VcUm�UUF�QPc�Z(VX�b#hX��Q
#TX�mEW)QF9J#�"�X�"2*#"*�"���b
��
���"���*���(��"��eAQPĢ*�F#EQU"%�D������"���*�1Ʊ�(ZV����"�T�lb"1���TQ�*�Kh��J�B�E��kEQX�������Z�*�*X��AYm�Y��h�cV
(V��HұX�ւDF#mKZ�R��V9j*0`�QTciJ�E��UUT`�Q-��UX�Qb�T���1UE�ڶ���U)m"
����,EYUV�mQ�!mh��(��T�b�m�*��~��<���|��������9�JJm�#-P&��hQ�M;*�$]i\`Z�5�[嵡9�(�%�J�A@��P�%����xL�hpL9����HW1r�hs.-TVÎ�Q��;�;�qצ���Q	no�Nv$�y������H
F�B*L���z��J��J����'Y��5�.�Ձa>T�X�v�� �V/��m���Ꚁ���/�wy�)��J���?�A}~t���j
�7*�x��nmu���?b;V;:�z�I�߹Vô�ـ�4e�vV�_�z�לx�qc�/��m�F�̺(�a�O�(g�*X�ݧ�v���7}��������O�|f����Ū`z�����������9FD�t�u�)D9 oS�(�Xzb'���w�p�w8��=w#�)�(��CX껙��}�����`�G��V�����٠�;��q�A�5i ��t�G��_�A��zpNx>Z
7"g��%��C�-��k	o}�	`�P۸{'����d-�R9��z_��B>��T��q\!_��Ɏʄ�^��综�Xz yհG���.����{���=��3O�#�P���80���һY�t�X�����%�,Z���p��K��[Η��衃�-��EGq^�}�5�;�J��h�i� ��!嚙��0I��dn����n� Ю��c7��w@�ec.�_F5岍�������;C�:�3U���7��6 ��#��b6�5�b�v��U���[�`��A܂.�p�r9���{xx��$FAGG�hx��~u+Mp������>��{3�}q����em� �!���i��A��<|�(�S�Zdt��T����"k�Ɉ���N-���b��ղ��:�%�5�X��pz�7t%{��q��Q���|FM�Yz\{5��/����J�:��T0�)f*S��`�����(o����*E�RJ�FQ.;�C�6f�z��AU�zS�����
�U�����}O�=�,χ
��{@MOY�_�GRw��׼��j?p�F�pؓ�����_5���O�SM�#�!vK �,t�b���W3v�Q�v��9s��f��I���nE��]��nsFф#L�1����PqR��yB�w�&�o�ԉJr�b���z�*AcE7f�ʤm�C�6F��X���}�i�g��cQ2��tntи�~]CINy�N���پf%Dh�j�F�t�χP����w"#]R���rȉ��RS�>���ɣ�Z5�+pi�QN\��a$����:+̐�O��"�Ak熑>S!�hv�uf���,㋃�i��u���v�xP�~a���-�LM�����E[��Ӧ@��of,��yfφ�'e˒���i�`��� <=F�v��M�[�R`lB�ԅ8���^�x��_3	�����cV��|3����>��.�;c�89���u�@��J�����#�*+�V@a�9��M����_fd`�X&V�P��l�8+B㷺�O����
�
�T�W�wF��J��ʐ(��ЯQբ�O���<�9ԫJy��4�%��ry��4{�6���
8�Z��8���Sq�!������pxB�)�b��<[�ɵ!E�k!���.�VPL��9�0إY9��6�=
栬Fʬ�N(��
��#d+�3�f�*�U��s�jҭMGL����ԅ��L�*�s��N��R���eE/�P��iVZ�3�m�0��o1p����)p�P��R6�swўNΈ�=��@�&"����p(d8��3���1]�i�މ�7@�/���Χ8OW�̑�6	�V!3�,sgb��LEC��v�m`{�e���Uw`$|�xkI���N��s�^���|��Ur #
��~M��˂��d̓E6�������k2�}����*��X��}I��4�W��:��W�=���d��O��ᘝM�FWg�Ǥ�B��p��Uw�/��G0'qd�;ƛܗ�sl�� �n��ˇ�����;���"P��;->y�����	��Zӈ��[0�O��w\@>�fx�3b���c����=㐡�Z��q])�T����ؽ<�DW�� � �.�m"�-��In�hݘ8T�߼L\T!�1w�-� ��_=�b���U�H��8e����x�1�ȶ_��,���/c"[)�}T���o�[�iYxƄ+��g80������ƬQO�	�3g�U�E�Ő�۶�n������_+���#���.�.�r|3�\�CW���T�wΔ���ѐaʱoٙIP��~��茾��LZK�.hV��7}W:X���r��L)��2��ON��l�~�b���V���f#���.��9´N#�v�u
ќ~�w��\{��9�0�U�\�R˜U�6���YY��<��~�&�l]�|a@/��T)nplڑi̪�Ǔ�9��B8r�����s!�P\��x�:'V�XWL� ��2MJ������c79�N���ܺ��9̧~}�{K�V	�1N��D(WQ��1M(�p��Q�~���d_*��XV���- �g(*�?߬K=�n�ر���.���~��x4ҭ�-B#���ݯw.�vF���.���mོ���T�(:,�i�k~#y�՞�o$�u�+J��><�݄�uq]\E�ҫ�����b�����6Lt}�y���qP7g}ʜc]�T�$n(_�>���)�m��tB�R�ci�Ĝ[<���T��q�����Q�������b��"8�ٍ"C���s��TC�����o�Mв��x�����<ϧڴ7�^�K�,�d5l"�����L��W���3��*�a�u�SN
�F.hdQ@��)H�Ӌޒ��
�Yz���a���/����z�*����r��O%��s������UC��1����sw�GTR��e�P�ޤ"��f6lCb{\T��Χe��c-�?�;uk{�����3˥xQ�3c#�S�FE9c:�P��^>K�aNo�Zy�
��#c2YQ#��wͶ�?����%��;�gm����ǫ�$�oÕl;�T�ň�95H3*6�(8���n'3^���J	�2R�x-�7��hϭ����{�Y�Q7�W�މwӛY �ٽjJ^iZS>�XOp?fx*�j���lϝ�:U��~]Cl�;��B��4��{k5G����o�_������I�"Ա��!���+O5�CwH��C�l���o7S���k/�Z\;������
]1�?�u���e<(�u��wT���;^E��O�@�(V��Y��ю7��p�KNa�E���&��C_���9>��4�����|�b[��[�2�k��f^����O�!�iP�+a���x��Ζ�5�n��s)oEN�3��a;����P螕ޜ�\8j#mWJ|���:{���(#9dY��=���`�OU���?Rն�G[d[��� ���R�Ɗq\!
��gz�&#��mh�#,0�T�
�G���>2\�����}��{�*t�i��z*'2<���x��V�4A9�;Հ��Z��xJ����5�=`�K��<�,+A܉P����io]�ۢ��t�S�P�C0�9b�}]�4<tl
,���
�Y�\���P�g
sЈ�����&a��m�F�F��X�rc�Q@���V�*.�.kݵ�aֹ��.6x��ܢ��Gl�{�DYe�|����%./�Y8!�YS$Ï)����`�SB��T���57po����!�V(�Ѵ��j��`���x�NlG10u��
����IU��<�Ϧuo�����%� �g����V�i܃��T<Wپ��w��(p�[�I������/��g$O]W[R/��ύ]g�}\q,��̱u�-��\���.���O)S�
B�<l	�"��:�+I3x��*�7��v���cJ���[x ���W��/H�cTIE�wh��-8�
��:��ܗ�>t�����x�֭֋����*>��ؼ�}�^���W��9U���i���� r�^��qc���U��OR<�r�!��.2��U�x�^X*z�U�
���{�/A�ۦ�-��hz㻭<�J�r����u�z�ܲ����{�k��s!�8d�s�u(@���7�[�N����?2�Ɍ	��O���.�ګ	N���
�"Ү�GF�R��\�U���>�B�S���\���c�0uTh���QӰC�CR�c����;�Ϧ�I��pjǩ{�ƶLOie��U�&�x;�����t":
tf�=��{c�V)����g����G�0'δV��{��̛:�����S�'V��?p����%�*JԬ,���#�B�1xR6��E���r�6�MvgR�B*%D��]�� 瞇��U��V/���-(��#2wU����֡�5�����U8�c�E.�J����)s�0�H���U��]{D�{C�I1b�x͏%�w=\4*���̨P��hX��Y.�Q��,26B�g��ҠH�]V5�0�ѵ�*\y_
٤����Ю#�#��͹�Tyv݇T����bc=�c�Q�L�
�.��R���1�R'ˉ!�ǂ��K���?3b��_ܴ�pmT�%�+<x���_AžL(���L7Mr�+"��7g�Fh�ƞ�+h��\$!��"�E������mt&����*Ld
߉�g�s��N�ߔ�1@����{���`�H3���iNZ�����H!V��Ō��FҀF��`��&������{Cb���b(#E�7�UV�{C;��	�[��r�8TT^:Q��<U^�C2}�6O0B�L��n� ȷ'��]a*��	����.�N�u�@@�{�ʝ���^���-�x9��T�:�&7�1���HN]�:_�uL`�!&Eئ@��\ᜁ^sA��|iՔ=㐡��s���f�������j�ӓT�7�.��ޠ.0�/�H��|I9��m#v\<*�o�.'MVDiu���p&r3[��.,�$C2:>\rʊsP^p"b���Mk�0�?Y�=^�D��8"~ϛ�;!=�0��ҽ�"�yň0a�29_���l�r/dU�1X3��(��*!a�7�x��z�!G�-�,Ӄ|�Q��@#K:� 陼՝���wI�k*κ�L�������9Ω�=x��b�oC�YX��`v���ӻ5��+æ]�#G�L[`���xD�@׼�+^C^dwL�3s˻�P�Z�EeN�K�ܼ��`���'~�Rd�R�B�(�{}�"�cKN,a;��x$��7R�pfw�۷�Q^�\�*��ع�G�=Ǖ7V��;�1�7g*�A��Ŝ�
���xx
���r`̼��(WY�P��Z�p{fR��2��0tl�<vV.�Z3��б���:��A��7swTk�U��a1Ľ�YZ�(�-��P8@R�،��� [>�P��x@:�R>��7}�OS]r#N;ץ̂��=-�2�D������f`@�2MJ�̔��&緞'�^����rv*(�R���Fq�pg�}�h���p��>t B�#LB��6�0�8�Y���+/,rU��豶�)�s�.,�yS������8&}00��%��so��El^^@��.b#?�yB�:>�C��}to�ҫV����@�������ؼ�.��9���s�pkn=.�>H}�ˬ!��mв������x���ր�>�Z�ҚC�>�-G:�,���Q�u`Ϋ�L>���"!T�Γ���ฮ�i�o9�=�m�� Կ���FU����P5�@u�
���?	�,I<����u��̬X�R����<AJ�T
zO9��j2���T����X�C<�����c�>Rn[�=�-C�kn��bp+�Q���<��z��8x�-�Vz-I��4��y���|��� �e�֝@�:��s�z���m�n��t����i�/*_���Ǌ�.�x؋�%�t՛J�+�:���f�4t\fP������Zy�bY��`�5��g�}���Ir��D(��u�1�G�ZϢ*we�y/�#sE� V���8v[X=X��D�F�#�w*߽+t��Yc��x���/F ��q��UA����*�쌙{��+��3T��a�O�(�E�#o�M�F�q�4ώNAܥx���Yu�w(O��e��W��}�<X�F3n�*����۔��ӊ�.�h�f�:�n�$@b�=�'cG�V>*$����~����П
�z����vz^��Ϊ��?nTt�T�'a������A�ޜ�x>%"6�t���C�le�zU�yS����*�ʋz�z/d��ϩ�کm�nlK�VB>�	�R� �ǐ��6�U��rW�&�k��1U] P=]��a?N��wK���=��z�An��<��Ʊ�Oli�2�jJ"k��~��~60_S �4,���C�P65�B�cO-�v�S5�a�W���M�npΐ�m8 ��ԗ�)Aa4��hJ�uCUp�l{Ŋ��UU���+��4�m$j��x�Wt]e���X��t��%���R�4���-v�ș��V�P�������v��u�]��V���Cˬ�[��Nޱ�Q�=�sr�Ϡ���n�!`�����a�-YU�7 �'`-U�����O;;,󲂇Pm���E������`��`
�ލ�n7.��=;�nK�Z얾5�5wȖ������8:e��:j�L+v"H5@j�&�J��'�6z�9\o�j�i��"�+<�ܽi\"��^QoG�:7��R�G������L���A=����y��|�JZ�'}�{�_h� >��9V>N�A��Nu�&�t	c�j��_!�i8���c,=S7w������e�t�i=�M�]�3N���A2������Ӌ�U��SE�&�nk����b�8+������]f>�H�4����Z&��R�WX	�u�֤�����M*{veM�L�>���q���;�X�d�'���ݢ�z��͐f9�ʵ��=r}�B��|����KΈ1��8"�q%w6d�5�r��.� Շ�в}�Lz>�j�u�GE���P��{u�_d��v��Gq,e�Nv�� -�5���z����.�¥tg Q0ob�@6O]��s�#��3(��Qm�(��U�G������D*��\;l��'l���q\��R����]Sh���)9:Pp�������u�l\=eק&s��</�d����q��94/1�:�l9%��3�r��շ�>%Ϋ�_40*��wQ(\�?,|�\��q�g����>���V�������/d��b�Nj<9c�ù3�ׯu=�����f��?K�q���$[G�ö�=�;��R�#ql}�
b�|��E�%�h]����\*�웇�ڒ8r�\(��a{p����\�esVC,�=�{w�bq\�� V�)$�B�,��W$����HiKN&��T����G��s�@	�Om�f�e3��n�݊[|���1K���lbco�l�����LԷ���4��&�| `����O��C�+-y�j�����R.Jt����X�r�wȎ�f�|��nf�H�ӄ![ݺ:H�R�YZ5,o�t��g�c4k�S�V�}�nޗfĥs����}Z�' ��6e���ϡPN���_4�YR��hR荝ˁK&�����^F<;���;dͺ����5[���N�V�/�:{�]w�rW��-�����?p|U���Tca�(]����rы<���^{<�,�Ev>�m�d���l]�@, ����+�0f�*�򊝷j�c��[��lî�U�ˌȀ�N�;7���-�eo�U5�CX5���7���xy���x�]�	囡>����xN'�m�ЩS�Ov��*,�56K硪f�M9����m�h���Va�P���o���;a[ʹ�z�K�v)��ÆL�ZA��F���~��.-����Q��[�1Q�7
cYk[KDUKJ������b�(�l�U�-eAVEU�ت��Ŷ��X��b�A�J�*�Ķ�F1UUE�(���hډmb�DcmF#YUUT��E�",PV"���lc�AZѪ�"�P���kTQ�FQb"	��#�T��(�ьc-(U��iQkR�UP�J�#X2ЩiYZ�b�0�rܥA�TAUb�m�����,LeA�(�AT�QkQ+V
�Lj����b0R3*4�",FAUQ�b�+j��
%B���DQAAm��m,�QF"��DF�m�U��qR�**�k���mFڈ*,FE���-Y��UX�*R�F1TJ�hQEbV�m�T�Q�lEU�"	iX�QTUAkm�V�-��-J�R�ETC����������<��U���y��)'��>u���9��x���g �jt\@�Թ��T"��65���WFa�U}�}N'1�Jܡ��k�7�^�5�iE���B�#�E�����^&k�5��2��dg=�_��u.C�@��Ֆ�O5�М��Ub1�v�,	0�Ԫ�s�����d�;��fn�'r��5���h8ȉ���+��rDsq����*6C��R�f%�U�t�\�ĸHq$��M�)�^���@��Z�x���>�y�3� :�k�Ԟ�Ww�O��	5�R��T����O���s�O�SM�>u�U[kқx�\񧃹T��JX�7�H��*����<E�,:�U�
��󨗼s
B����v�T�;<����jX�Y�u�r�<�;�gjE#�0�Z7P��Y� v.�M�ʌ׋S4R���+b&��N����>��4E��Dñ�|�J�:6�خ�۫��H��ܡ�(�f�9;!�"�jAU�����Wf���Fnv-8��X�㚳��8��T�o.Ďz�vl���\jX����m�����N)�8W@�L�Px<�K�ƍ�{��'�Y	�B��r
�iu�T�N�'v�C�#
ˮ+����U�zwP�Z~��fn�$	��и�ѣ9�Y�����i�T�7N��%jO���;t3��9i�S�J����f<�/�;ɟmǏN��p���o��������%f"�rLwf�O�{��2��N:�dN���Vd�7/�]��U("��8���H�*O��a`��ہ���"�[�Ú�rf�JGj��{Þ��຅3�EД�@T�Ѹ�b�g����	��ۇ��&M&Y�Û�0�X^:�T�E�Q�)l
��+�TF�ԃz��6�(ǮVQ�k\��6�b�aڌ�'���_�C��!b6Ud�qDN�
�Xdl�b��*E5(�Ij���*"��|�b����ryN\�윆}��^�r�C������1�텴6�gku4��b���ʂ�i)4m8�CL�6z9;:!쌊((��4j�z8�x���ܱ �K���U��	|�2�.K�1�#`G1A`��I�;zM�s+����o�Z}�p�늈��$�����ʝ��ʵ�{H�^ J�wb{2�ժǣ�a�f��_����r"���)z��tM+3����x.5vP��^閍�����Ym�*!P�WG͐21F��¦	���-ӂ���0p����գP״
��Rs�WA�b���)�/��.�P�8=��e.I+�M$�LNHb�ȑR��:�ݹCtt�}*?z���#ɩ�LJ����j�g�-��~�wվm��v��� ������{8<���D�ڂ#&��{�k�n!��� ҳ� x�m�a��zd��EG�d�o(;><���D,����#/<Δ/C����#�P�����:�窶����qb�g�������"�E�>�6~�<��e�g�7d��A9�">�-�m`o龕�[UV��W�����՝�⮝>�`�\e��s����7�:s���WN���O[�
=�mf����e`Oy�ұUr���׫F�#��+&+�v�Wܢ)]�%Ժ_�u%5�yj5�·)p{d�SC�9´9�x��!�&n�f��!��]0ɜK��D�����8��4��o�~�0g�(,����b
h�W4��dR���X=��IS�T���m�Ẽ��(�8%��^D���-�����J�9[�v�R���y��L!x�(�ƣ��v�%ά���Y3�c9S~N��w���5�����|�)�7���`i��xք�j��2y��t�O�����^������&\���t+/���Ρ�6c���� ï�P�E.8{*	�/����s��<�t��)U�gO�vV�s&1�g�pj�<2�&l�%���J���Q����7w�w�<�)i������:S�����Pk�;�dM�0�1���z@����eQ;�˴���L\����]Z����pD.�v����r�r��L�3B��7�Fٟ��$����/st��r��~
Ѩ��PY8�Dd�(���nlG�)1ˁfQ��!=+��W=s�Rr:�*0�8�WN(��yM8*��y�I�O� ����הY+5L����Y.=0�TD��(�^�[�UEo������)'���;�i����9�/��U���C S�[���5��,EBN�'a����L	����n� .E&W{��xd�H/w����F�]���.X���d������7��S�c��Z�k���'*b�w�hlG�`���[�~%�zV�jc�2L ��Vð�;0�T,�e�5��h����J���/�[��+���[�����4�m�71�tC�*61���1G@z�����\����*"}f�������ub�5ͻLt���O�$����.~���M!l� }�1SDN�h
�<���z�g�}u#Oq>?CJ�n��{E�A�3��m�]��`c���Ψr�Y�'a�<��R�F��N�Q�Qb�;(/�
Bd��d�<���F�y��Y%ɞޅ�v���F��]� [��"� ��0�Wy$
��j���DU�C�,>�Oҷ]3b��g�.����2&�h�ګ�41^�c��:���iSy��8� z��)od�+ݴ3b������Z��tv������vPlE��}�3�A���@�_�OOX��Db�29:�K�R�H��e�̮�k9u ���|�,���*�!�^J����o���_̄��O��{�Tp���q�p�f��77��3��ƞ���'���C�I�
�(8ppu{
��>�f�{BAJ��(r����Y�A5n���W��u�)ө{To��GH2�2lQdX�
7d70 at�N�i���Yr&1	��l�[���q�a��=��F�܏dGAbw+ŤS5η��b��O*��~1��fS�f�1�ܸ~�N��8����ܑ�d����o����}����7ʅ0/J�AAɊ���"��"��M�Vv�'&+z(�n�f��RXARJ�F	1x!���m�;�F�@B��9��
�S1�uio˺i5kRhGU�@�@���$n�8:�Q�=7��S�����j~�l1���JT�e��%��}��*�n?0ؠjLp�U{��4�`Z�v������1�35~�(���Z�tB�����[�X�ݢ��:P�WeV�WRV #ӆ���t��Uic.+eڢ�o�ne>�5�f��Cܚ�鯘��k�*r{oe��ռR%ΚΝ�uf���v��O8�j����%!�Z�s�}��"<.���%Z�_�n��(�)�nqُ��; �PQG޷,���#��V�����i	�6��79r�E��K*: 1���m8���z����FL�u�H'#���B��+�=��S����{�߫��t�d�q��\[��xl���o�c���n��v{]�J�3��0�t�ǫ�]Mޅ,y^9�[>8~���ζQ��+��FBe���p_WfK�<��a�a����3�r�*�>"z+�V Y��~��92�@��#(����*JԬ ����xW�Y�5�*����ԅ4*W
�������pf�����Ҁ��`�p������I5�>��8q�1~��>Z{9�R:t
`PI�p�Q3�,-�\�j7*�ˊ��[�V`�y�_9�?>(	}~#-�㧱}.�Q��,26B�L�ٱ�vs���IF�X`��oЫ tR�S�; ������>��d�M�pb�VTQl�G;���9
�T�u�&�lz��VM� �(���r/FӀvwd:��9\��&kp{CB�Az)H>�uge/{�Zk��풁ӯ�dTrJ+B.�j�:��Ef�6�OCr6��S�s��hd�v-�y��9��3��xNϛ����N�[z�s��l�)�=��G���]ӫ;A���4U.qhR����zg��hW�5uJ��G�����J^���{�ɼMC������2 o���/qc��U~وfz��<�cw��s��&uz�b�#�{r�@����]t�!�����V�J���x.gk�QZ��ML��0��،gH}L\ߚ��$sd]�`�$ҳ<P��NhW����I[���-��ڊau�V�ܣ_TC���E6@�>��O���n�����%�pU�vNx/b�@똇�j�}���Tʫ�0&�2C���W*)�Ay���<Ϧ����S�/����淞�7�JIg���G��y�e
!��~pWy��r/dQ��qU�9�3!�]�z��RK''�2(ԟV��'l-�
/��(9ѓ���FE�b��b�P��`C,�y�U^v����h�]*;���1j|ކ;��k���g2����S�\^@d����,jbR��v��Y���%5�:�CÅi��L]F��
�������*����1�a6�CW2�h���k��v�:��Й�����Ew���P8@G��UX��ŻG�v��l��V�Ug�o��k���C���5k����l=z;m]`͝�Nodk��7vȜ2y��)9�뫳;��3j�Kܩ��	��Q{xen�k��t��d�ޮ�B�8`��f�M�����c��[+��K{Lo��}?��Q����蹽U��n�'�sf܃��m�.d7*��Ιy��4�XR�`U����p�}-C��b�T��o�}e��QJus#���ɝ�N��9��\Q�b�}r�nS����'0@��Ⱥ��+��eLw�)o��nA��"����?n����t\9���4�.�q��v�� 0�|���)p��a����ߏ�jѳ�.z �����}������vP�=]k�]	�Nh�x?��g���9M͈�E)[\d����ҭ^���ܸ��O+��T��~�F <��fµૐ\;��Z��S�:_dN+W^g�$�L�
����v�=0�b*���f#=�PΜQ�q{,U�S�ȹ{����v�#����8e�]zk�HP(�-͍P� �x�	:����5�L�ʔ�1�&V�r�*�nnL:�c��l��m;��?aY]W����Aw�.]{�I�٣����h]�__.bUV����A}x"ו`�t��\,E�:�����^3y`���:Q׶������r�b^�P�m�rkmʎ�m���t�����mHW��{A�C�5={��!��J�B_-���,�Hp]�hQ��
]/����3�8�YՈ3�4:�F.��7�o��{�`�(�*ܫ��a��A!r~����y��J��y����UB^x[��xS%Rñ�>��g�*P��nb�X"�bb3�,�k�h����p�{�t-�yޔ̪0�U����V+�Q��T+������S�w�I$8SU.lulB���b���Py;��=R�><�!gr,�t}����[��p�)=��(�Ă�ۉP��B���K�k"ݧa�<��SʨtOZv���B�\�7�q�-�sUg�I����.��р��E�����}����	�nn_��h�����y��w���Ξ�mb�vL� Q����g����U�!)�t�_Ӗ>��ly��z��5+/�7�ќ��B��K��hzR�d��J���֊����c�w���w�H�(��W�LY�s����
Bt�^���Q�!�D\�:c�(O(f8L^�l��Q�#S�u�T�����Ca�+����Ǌ4��	�����Qb�.V:���,wN�s�L!V�߭��Λ0)iwk����GG�|%7t'�������Y����)�l��>n0���������G-4\�M�[���a`�Cܙ2��9k[0���.��d�f���蜰�K�]��:n� �Sx���3ܹ�1��g�w(���Sr�Z���`y����A���̙z�Z���Τ����u�a��]w#~55��Ez\x�F�Pl�}�Z�7���?�x��Ԭ4vH� �.&n$�N���4��x!b��%W#��>9��<>f���]J�P��b�L9�D�d�՘�19w�U,G@�
��I���N�(؞�������>V'�)Zl1�<|���6gK���ޚ�c:")�7�X��R@��w��Z��S�A���Q/x����wֻR�
K��<�h����-��<V�ةۺ�;�-`Tݱ�lbʤ�u7�T�=5���b3e�>Wy9�q�����-��>NGs�5B�t�]��8�1w(�Q�!Ըnhi�FA�*�'�!D"H*���l�Eo{]�k���թ[��&xKX9��^g��'��Z+��^*{�M�����)G��T��F�Z�JomEA�J��N�`��.PʥQ�,��$(.V6md�v���Ճ�)
���	�w�,9���!xs�)p]B���J\�y�F�q�Ψ��)���ç�<��xܨ���6�| R�x#��(޶%� �ტ8QT:����NDC�j}f:ָG���i:ov�x���-lI���lm�XMN�c3�c2�MςB�K�3f�r�KW��Wg ŮC���
��7J��[�U.���}���6��^N�t��)S�/^u�[����ǣB� 5u8f)v�&��+Ms��r��EZ��Ή�v��<s�	{呤���D�j�����E!�jͣggw�.%�����e��Zq�ݝ�(⓱�d�we�5����2�/sK�CB��9GtR���z��_LVy���x��n�t�z���q�2�s�F��v���Ve�!�w�kI��}=ӝmv�����=���Z��3��Y !<�N���^p]�(V��nY/;(s�ӱ�N�{�ѣ8)�vxczt��F�^J�/x�)�����cg��nͯs�oi�~*cx#��s���O��kߔ������r��M�b�7Z<y�0�h
��A�!�]�}JUк1d;A;���k�9���z�T�K��U�2B�2ccl&�q�و�������S��I���(��v�.ќu"A��Ib�;�
�G�F���{VkЦ J�'�xrN�+k��K�,��o���T%u�ڗA]@!����$v�܅��eAN�f��L��xm*��`�9��:��]�v'Dڒ����n��$^�h�C��}� s�W�_C���l)fU���5ӗ��ێ��x�����8�3��PG���b�pɝ�o[:]���
�4��K(��C¸��5��n��1��8p;\��6P��삝��2��F�k���Q
V�sA�ᗔ ��-{�;T�vS�z�v�dS7�e�ek�)C�(�8��}�Q�:�nM@2��p�2=��Y��DFC�}�onu�͐a&wn�+4�[���S�X�;D��X!�=�Y�sb�5Y#.8 ٳd�϶���e�4*�ō�%�;ޤ��U�7ׂ�,h�X��6�#"�J���\x6����_h���i�#/i����۽��Uz���˛�S�D����WûS�H��E���M���lc�-c6�挏4�K|oje=���,I�d �,���O� lϹG�d��26��-v����.�ψ꯼����N[��Cׇz^�S]g!C��(5��e4q�D�C��j���P�w1����])効�]�b�Pu��Ȏ�B���Ô�V�U	�3/v�Raj�K� nX��G����Y��/(7�"Q�.�.�S)��Ec*ڗ&�r��2��<1� x���8Cn��| n��p���s�v�~�0��7���"���gAl]LM˓+�a�`١�{��^SA=��\k%�<��fCҷ���w(gy%�<�
�9{���������=Y���Z�U��UT�� �,QEQV(��,F%�\lU2�%�b�U�1A�meQ�QdQU[b!EAj(�Dcm`�j��QE*-�DQH�ʮ[\�1mm.Y�I��AYF���Q`����)EĶѣ"��A�H��-K,A�Z�5VZ��T`�TR�Q�\K���,m,D1���"9lTc"V����E���K҂���R�dDQ3.e�K*,TV((������j[,�kEELmJ)Z�����E��1`��VDP�*���-b�ւ��b��R"�)U�����8�V(1b�5P��-UEF&R�EQ���ATm�X�1+QШ��q(��UDEQD(�2�V1UU}��o���y���w$��K��n=�F_و�V�TY�L���l]�q*�����W�D�S]�8�V�d֕D�Ϫ�D��9urVW��𼮇r��qOb��q�"�(��($�B�]���"u�NLv�*��p�
���/f�GE�Md'���Qɞ��F�Fʬ�N(�v K*F���O%��F_�[/��:��R�<i8���%ι˝�U�r�uϬk'*mK�
���p�:�8R��mq{���`!P}�,1:v�IC��YX�)�����3͞�NΈ����Z\�W,KW1'J�Pؘ���*9��p�@�
:���*���X �:*��|����w�b�9�`�X�\r8"��;f�И�� 3��Iٮ����P��ʝ���^��xGL�>�u�^�sS�g����U�P���j�0T�͑v����ns�͊��(�,/�+��oS������f���ܣt�-Z�"�l��G1Wg6�+�=g� u�����b��T���ȸj����T12C���W�<���D-���)~�����왽��(��95����F��}��1�� T(�������pH����]y�[�!�YڴDF�ڕ��4#��;Aoڗ.k.�Wn��|��ǵf�h@k�h�Vk�B��b<ݒ�/��r�������!�7���9衷�jt�8�Kllw{8rK[m�C��q*����잖Q=��%n�9zogBU:��r�LJ���������E�)�쓆�	��(�0�FRNN�
lA��WyCw�ͨ�j�u�3w\�j��ޫ�=���^
Ŝ�N*�o��ʰOA�~ɭ�m��{@-��dN���A$9ǊRp���Y����LO҅u_���xp�t�=�){\BѨ9��}$���ty�B�;���o�Z (:��6\'U�)�f:2���\W�:��u��of�m9���@��n!��� �GJs�ٵ#T�m�s!y�Qnr[:e��Alu����|W^gG!iT�����-�Tע�Ղ�^7��Zr�pK�;FUw�0��҉�?{;�+n��P��V����Ul��x8J��)˞�qP7g}ʜ;KI9��M���Y{�/��U������ �ΔyB�K����<]��գg,N׆�������J���:���d`����*�s@>�u�0�ct,�x0,��L�̩�G\����uR��(�cLB2﫠���;�F #�8�WN(*�P�����"!�}�/1�˕�'��ZYs�Hޞ�V:Ù�t��/V�����`�cΖ�
j�0,)]D�������G8�p�]�>�:%T���S;�S�J0�]Ԝ{#���GaO�O�A��Ef��fz�%}�y�Ae-X�U���70U��A	��(S��'�����g�EP�,B���b��Tw��;�&z��^e��y�;s���I�A�L�af�u���C!��,EA	36!��Q�b�n�=7�����4��8���#����lX�g�FPB(d�,t�(�FS�'�O�����=K
O�����~���^�x�;>�H��ߑ���4��LR]�ޭk/tGT1k�Ʊ�Nȟ�ܪ�Vgǅ2UR�x-�7� �z,4�hU)��Đ3g�ژ�{@#�Mÿr�|�Κ3~���]�}���V+�Q��P�}�����zBe��������^b�`��{+��K5T)��r46�T���M�\�)��De��&Q]F��M�X0G��;��"��O�*�.��n�vxz1N�U��ޜb�c�N,���V��=T��U���>d�t��	�s�0�;+ϝa�#�2-�"�j��L�kKZ�57�"��>��R��N+�+C�`�T�
=]������*�����_Y870��_5Z���gp$Ϻra�C�b8.9V���C3��հkzZ%�Űe�>�v̜7}i�b`��٨��R��N�Kc%J�d*z�|��&�luGR�D.�ъuޢ!�ֳ/u����v���Je����e_8�x�,S�M`yTlv���(p'��y�6fYθ��g�*�f��T�+�����R=�C:�����Y��:ms�8�
�=�(Y���z=�d3#VR�B^^EװR��i���,���y�ڶN�7̕�6�BkQ�*n7��r6�P�u�Wn;f����ʥE�ϖ�*""Ɔd�d<%c�cqEK�ux�FW9�d�
rFe8�kӂz�%��/�3�1ra��;/")v�|�&��L\<�2`�ha�ʕ�1�|�W �{>ׁ���x�sb"��gr^���5��#h� �R�A�0p$�����[���A�M�)ϱza��j��ہe�
�{�����!y����řC�@
�fA-S�o	�E�r,vT9X���:ЗQf�OK�g� �,��1
�e+��c��b�� G�P��]/,:�X��Ns��Z^>W��ĠWUi�{F8Aۦ�,6v�8�1<7���w��G2�]gñ�Y}'|���]\���9��y`���}m{�Ռ=Aͥ�7@N�����6f���xk�e\r�ɘ�`�h,�����m������ۜ�/'�>p��d�s�T�*wQ��ɳ���oȊ�g���nh(��xt�t�_R�we�EMI��y���@мcP�.\x6p.,P�m�!�U�Ƹf�z�g(�ԬF���!��}����T��w�9��ү|�O��Y��>FA���B(��)�FF�gb�jMߪ��?':��������k<��T"��
������Nǔ�s�]ŷ:�9h]�v�S̗Bo{`A����<��~pe���Z\C� e;U�#cv�wu���%=8�R��wKZ݅�����
�*R|�#�k���-BU.P���y��[ܤa^��e��R��]~��c��ث<�uO�t�$$���Q#��Д\�U��ă��\E�_K6�8����{W���P��+TOR�N(��
���u燳�?I�_P+�
"�n*A�J�
z{d��&6.�9���>�m�<<Uy�wS����CԶla9H>��,1:�k��<��J���O�9����&���1��}��ǏX�3st�P�n*���*� r��
Uc©�\��\_	���C3�l3�)p��o+��ۢ+�:�d��wBV�� fz* .@g�I;5Ā��=��i�Ui����"c���|��Vc;؀2ѹ}^���͘�x-λ�0�Im��E�P"��F����B��<C���/ìBfw]��j�pG˓M^�V��^���1X�E�.S���{�3�`��J.ָ��]l��yF�h6�S�Jc*!u� ���z�Wk�n�y{� %\�¦.Z��;͑n��̊ɷ8g v)n����yq�<I���5��쌉��w(���k��-�21Wf��/��{�1yyB����;��xc�
�#v\8*�[��� �W��v:�sP�z�s>�CiP8d��>O��z���(z���䆋�}��S��P�Q����ΤuO�j��i�ڡQ9�H�.�q	���L���:k`�m�Qxh#)$d� �@MsD�U�d7_U�QI
�®���a�°R�j��)r�-F�u
��q��	.G���:-K{���P��n�v2��N:͜�IM@�u�$C��Eu̾�#�R.9j/%�d��iKb��D�,��z����^�N�]g���J�U��vʁ��:�T'{�o
�Q)����������>�>�z�Ks�6���n*s!��*X�Ιx"GD�-]d#��6����Sgr&�0+�gFՖ���S^��V
Aq���VN	�L�J�S'ƹ����uiNITCzH}��h�#�.��vzat��bR;��`����������x9�c饣�h�Z�\˾I��7Ʋx�snNr7V�����JZ<(��$B��ޞ=�{/���+A�wк�0�X�{��G$=�ګr�	�a+g9@���.0��"8ő�!X�@�!A#�a[[�8*� ��M��������=�)�J�ss�e�7S��`�U���)���EY� �R�{*�N9b�9W�2OwZ�jJ�x�u[�QY�c!?R��X~utZ��Bt�}��U��~J�7RT�X�:��Q�pL)�ʏd�q<�0�3*�WA�nCj �l�3`+�F
��_N��IUgOUT'MjI�ı�2�>�I�.
�=0�����X�~��#��'2⯦w�[t���ODd��1���B������:�J�nwD� D�������������"��b���J�����������K����q�K�+k�~²��^xz��.����b����tF��M53'/Ueyޣ4m+��� ��"ו`��oݮ"��gjc�5MH�W>w�y�/A���^,��ш,;(?�ʢ.���d<)��,;p�TP-��{��,QC�:�͛/4p�*���T����9s΅��ҙ����}��Ͳ�*��|'?4,�ER���g&X;��t��m��룏h��b�Η�O�^	����F4$X����-E�H����<��0�AF���ΏrJ����r�b�Gvq83G�n ,{��]%0$غ�����op+�쬷�ձ�ۭ��
"wN\��-ԣ��\w�f��}�}���R>S�7k�X{�\�N�x{ம��q���b]����L�,���j�����������jN�c#\=6�4%��⨈k(�a��VF�s�:m�q��4^dn���߉Y���ɢM'	Îev�(�����u_t��AG	��2�V��1k�^�ַ��m�w�]4�I��W>�Eմ�!�vצN��w�x3����MV��r��'r�U	�����K�wj2*�w);W�0�j�v�n,�K��VuЕo����B*Bp��j,c��mS�|�հ)?H3��Lv��)f:}�Sͻ�:�?Oye*��4q�ۢ�<��:��@)��{v��C$�8����pKdv�	�\�ܗ~�R�j���r�O;����UϦk-g�2��;J�z!z��_v��V�4������cP���%Vq�k(������G�Ҭ⇗���}S��cUOg=Ƨ�7�ذM�O;�;�Jr��<���� �`���V*|�봤`^��4hb#ǫ�ξ�Jtj~�<Eo$�=Y��J$�v�p�Y-��4�1e��+��	W��̕s�J�N�Sϕ�
Vf-���o'�R�.��2�e*I��D�{h%�Q�d�w���@Y��H!W�V���2�䱮�N���z[�1}�M�u�	\a�}L�_�.1}f�uQ��t��
5Q��]�׳D[٭P�O>1b�k��R]�qR����υ�ׁha��AhE����uf�l��\|�:��59�O}Ϧ�*/O���	|r���A����]|/��E�^Xә^�2� wU���س�{g�>�.B�����ys����ނ]�ނ�u�j�Wi���������~{%\.�	��%G�`�A�ۺ�5�S�n5�q|�
�Ɨ�ڻ����p�P��N8$��b��ќ�g\�HF^X�,�;�V�'���j��ܟ,F�ni@d��ј�ӣ�W3Ӵ���X�&�̡RQ�{V��/ԭw�ю�o�Bج��Ru֔Kf��{�����:�6��A�K�msX��2��j�c�:.K�D*��{Q5�v�����pd�$�h�L�amBl�������j�W&��v�;�;|��"��,{�Oٚ�u��	uB;Q^���*�:������C�f0iՔ�R
��Gh1��xwy�+�Ɔ��&���R��l����R�Mͼ\N�x߲ʛy�7�W���R�\�m�A�4q��imjg�P�wRXẃ[�3����	�<�
!"�F���YB�s����3^�J�J���/D5�	���"G1bhsd�3�~�����Y;|�!݋��)�T}��ۤ��݌JL^sh��*���6z�8�|�LY��X����̡v��7G�HW���#���<�\���T�7[��؅GVM؎cz:a�B����ЯaA�X�Q�3=�1Vg,[�Wk���ezt*��c�U݈�^��#s��~�H�
_�:H���J#�էSSS~דit�R��e�Vmd�C��'��_�n.�ë\x㒛���j����e��my����R��n��������c.��,8mn��b���'��h�+]��!M�b���.��5� ��UV�80s���F؃�o�Yz;����תܾH�Y�<���*�c�k@INd�#ʅ�r�n�F�����Nn������R]�3A`�wڲ�9t���H/lx�����l�gcl���4
˳\;�X�VC����%g�]b�-�'�姂a�i�}ݹƆ!�v$��N5�g���[<N+6�;p���L<o�8�Y��i�=4�
���X�޾C$c/��b��K�F*��hH�n3�R}s(X8s2e�ކ*���]}���go[+���շSM��`����KN����b�Z�}��Ӽ��N�����B����ٚ�Z��VQ'��+ w�Ή]��W��3�ü��r���7$AL9�s!xnp3Ԏ4�<���gu�����Ay�K�o�I
�Q��:�v<[�y�r�2�g9%�7�Q]FYi,�ڐ]s�7	JlF��w+wj�Ѳ�Z��Q``G����3dhTr�wkz����GzFs�{�\�h� RG@��i��	ZAʖ]��I>]���|����ZB5r]�[	�Z��l�;@������Tg2:��c.dl��^gj�K�uwN�#�一\�iue�[�O�[�Ȍ��\X�@�\�5e����̒m�c���4��a��\��j�?]n��*ּ���+{�����sa���D��q��U��o��M�-bW��L��3Ǥ��Κ��:����f�Q�ګj��f�3;��t�&�׳��ݺ$	���˙�)��/k�~sS+��%�nԗC
5
(ֶ��?,�ul
u}��9���.�G�N+� UJ��7ܭ���Fp�Z[���p��ˠ=VM�)C���>��C�a$D sMfh͓5��0o*�E��l�nq��m��l���;�0ܘ�5��dq�r�2QŊ��Ш�*�{tb'[�rg.���K�Զv|FQٽx����%pH6�OvD]�F�*�����{-��^Y�5���ݛ��CL�:�r�ڃ��s<�z�a�D�����җf�����<@}Mi�Ӿb���X�_��T����j��0e��}S�N�hܩڅ�8�z�����y�ە�"�zx��������O��9tʉ��ǀ��띸�2���j4Qi�<Z�ojӡz�L�:��ι��A��r�$�\d6b�\�|��cz���s2ko*9H�����c��c�VL�m%^���F�~/����utٙ��Z�l�����k)����d��)�(i�zZ�&�(���Y��D��̋A��>"1p�eк�8�����-��J�}V�M��K5�Z�M']�/���6F�,���Vi3g5�F&�v���#�#k���Ҭ�j�&M�!X7�T}:?~߲QEX ����Q*QEA�/���1T[j�nY@V,DPTUU���EQ�P�����A��U�Z �iDX*��[QDU�
8�墂 �7-q���1A�8�E`��F���Pe���aZ�QUL�j���J\���(��TiE�.er�-���U��e��W-�ZQ�h��Q\�2�UFf\Q1��
�DR�3ڶ�Zұr�Kk)�3�.0��ʙ����X�F�6��9Z(cQ�`�[�nYQU���*�,AL�
ˍ�r�R�#YR��UD�DEDEJ�\-Tƍ��
Ҵ`�B�qȢ+mT)h*�U�ж�b���Tr�e�*���lU-*��Tm�j�ƶR��4�q�1L���*�UEr��4�ʢ,`��Z�U�j�9ZX�XĩX,QKj�T�b��ʸ��T*�>nJ��SW����ɝ�t)��J��B�\����W�cQ�7��x�����V�ɮ�ܼ�n�\"�T��)�����]��"���k�X��E��Qמ��tI��*��K�y�X��c'h����SЛjå���N�IMx�]���%v�9ǳy�U_(��M�,�����q��18�ڷp�Sq3�}��VFd��z�pFD�y��"\��JDq��2e�i<�k�e>V��>͘o$������N<��`n�*�74�TF�D�ec�/U���M먊g8Fׂ�7*��u�z�I��h��{����\J�U~}	��E�n���\pEPw���u���ucm<�B*Ey8t@�wꭘ�NC1�K��9�z��;����#�>����ë��
(���7���0&�k�UZ�����p���8%��w�A2;��=J��=���.ٍu��'��N�1�:Vz�*ۓ������o1/T�)�N�xV	xO�mC����)I�t�㝜�u��疤�l�Ę�'�+���g�������$2����A���v	� ��V�`d�D/�X��e���g��+jgGxV]sV�����R+�u��.FGc�j#(FFf�����-tΠ���=m��*�Ƴ3��f]��-�G�)�Ì�'3(-��jf��l�D�6h�|"olԽ�y[�j��M랳����n�)%�KR���Dr�B�t�kz�y�ڣבO������=�zc�}0ot��V>�b�k�dr׽��c����Z�?YU�XW{��\�=��ڵ�O��M�׊c���#�R*q涶y ���Nq��¬�K��1ֲ'r�γ�8�;@���	�����0�jj9�Q��>�af,���9��JozK��%Gb�V#�h/��{8g��'<�
�3���Ha��L,v�C�`B�N�q�J�Q{��燨�f~��NWכ�ɾ�UrVT�����{�Gͳ.�t���ヅ��Q�r�����ϘuUr���wS����bw%b4
nk�`%�5b0*�����g�tY��w�Ze(�N�q�g���3X�%<���W�͇�X��v#����Rwq�B2���.�h�vV��(���s��RSP�
̣�ҍ����Grz�6��wm�!�Ft+�9�:��"�]W��E��s����tvؓ��)�+o,[H��;�X:�U�n�t,f��ts�m��']v�I��7y�@�} �u\-x2Uۦ�ڎm�Ո����d[C��5��o1V���;"��s��r.�Ol��X!��mmΩ2����<�vKb������nE �5�N��Vܝ�Y���TDz"�J�t�nd���x����!1e��49�Uy����[�̡v�r��{�Ou���(ATյOk�t���tRcy��|"��lЗ�h��Y�IkAVJ[Oa\�e���>K��y״y���#f���
�Fq����Q���'���*�<7Lf44�F���O7^�"�8��ݴ�s��l�A��k������;@�0�5����gD`�4Y��8S��K�>���M�����ʺ�D\�1WxI}�s��q��u\	�rq�}wxˊ�]��]�*�_9�`�o����*����>����7�R����Y�7�}����pfLʜ1��
U8|Mx��bSG�X�2��xTVi/��+��$ق{'��I��Ὀ�J���	RN	�ɾG��{zp�M�}4�У�m3��n{CN�M��l1L�r�S�/[V�kq�+�.��p��*8(]c���]D��Vb�e��k6��`��{O�ڻ��C޴���il2������c�z��hEZQCX���O@�g�V��o�v���N䅈�@C�m�T�C��v.�޻̉�����_2��v��볺U�q�Ǝ0tf r"�;s��F볯��WK�: j M���O������}kb�Gf�\{�W*1δ���h\��U��P��ln���jr��BuȊ˭�UBB�~2;j��A20o"�PUș�� ���Zv��7(�rV���l�#8��S(L�����b��6O�F��8��ch�obj&�;��߫2�N{�G)�2�GcA&0�h)�DO_:��f��ND�ze%��Kv���Ŗ����]\ӨP���_x�Dv\=]�b��/Gi�ȰP\V[�*M��o��#/&���~����ꪷ���࡞u�ۇC!k1�;�-�f�������I�x&�ш�=w���ը���Ď�N�:)�w�B�G����L���Y�v��7G)
��#{��Nc*gm���x�=�ԉI�A��FS귏�7�X�v���0�he ړY�Lˤ�q��v�U���٧�18��9�%w]]eQo��C#��WmS���16yh�OW�&��qtG�Q��e_�n�D�ܭ�&�'�.ơ��v�q�׳YV�"�nk�X��E��*;\޳�Lj	�9��1�fÎ��(>8��5Cm�t���В��u�V�3��y�T��'X��D�`"x���M��v����E����q� ̊�Ou�$�%}X��@-�G��2�a�k�r)�O>�-U�^��u;���Ӵ�Jl�	ν��F�EªQڏ��U�On`uzj��U�8,Y��`�I�W�䐱75���	�f���A�e2�z:71-qذ�.�JH����E���R[m+f�����T��N����n丌�6�V���v`[��+��t�{�N�k���Y�o}S�u�z��]�p�ֺ�\�zx}ۉ� �`�R@�CC�6�F�������k�k��ǅ I<�uu����g27t�עU�n�m��EHN,���x%\�;����cpK���3� `���t�f9��:�G7��.EPs��\�;WOu!�U�n�����|U:G��/y�D'~8ev͓S�M-ʫ|u�Q֐BX7�H���m�����5�*��l��{��3x�M�N4�[i��QS��%�!�!bhk���CY;��³.����!b�L�Orz�#����G1�J�i��<�h>U�6a����W��h��+d�Q��~Ͱ��3{��|���&��s@k��QS����-3u���/^�Y�:J�8�}���bb�j�m�Z���٢lRB`8��n4}3;��'z�^V����:�k�R!N<��k�K�D;	^g�ݱ{���v���S�Q�TqF3AA��dk-6���m" .�W/�Et)�|��[ل�I�ГLs��OB(%��.n���\��j��TV�[�"����i���OU�<�@����b�Uh��!Ef̼�b��m�3��HU��Y P7��o9Ȳ,���A!w"*�f�K.V�V���=i���t(�[H�>� ���Wk�e�ےw9�U��h�R�1.��ջ��W��T���ʍ5�GW} bZC����s�QE|	_k�߾������fX]+ .q�1+�l����X繜y�+�;����n�wk�GN䅈�!75��ggP<��i��p��IŰ+���aH�׸q� �`�V��e\�r�U����"B:�j�7��Փ:�	�r��;������f2��G6�9�!��V����3/'B/dW����D.�}{v����q��ևA�{gu���n��6�'c�CH�v���*�dL�Z�Y�-�;J���w;��r��H.���{�#	�-E��q@45�3Yo+2/d�m�V�.�-A
;�q�g��6v�8)���$Ƒ�T�這�?_#ʈΟ��Li�(�G-�Q� �)oR�G���(d�gD�Mא�%�Y�j�H1j�]bz���T�R�.&�P�xO�J�DC� ݓ��@7�f�S�Y}	�yo��}E�ۋ�I�#{�z]0*'-*z�#�X8Z��/P����	�����R�_e]۬ʻ�7\����-��2S��{F�W
�q�m�[޶�Qbi%�]�Mzwv�rp��(^{�5���N�&IȽ��^zy����[����X	E�}�WYH����1��W]�-gs���OU�z�����s�1��E�	��/�U������A�@��as��9\�-�S:_Ӌ=����h�q���R��	��v�'ѯ-=R�\��iB����Ro[V�k߼"�W�ew������ճ���-8&������v�*A�^���WqS�{�w���bL��%3ekmt!�s s#=��(͛+U��ړ)��w3��/n�og����Wvʷ��4�YV�|0�UB;V��Y��^p�3e;>k3��IY�К�ˊ������dDM���L=G7NS��@k�fq�*jP!3a k놘����b���{k(YRT�C}��I���䖆�N4�͑?��g7 ;�k"��+�A�aV5H.
pfR�h��{w;L�������K�ZF	��\���il���rд�Y|9)��ɜL��u�p,yAS���U��o��uPh�*�q�o�GZ���6�+�{��#	�#��E"�[�1o{''�v6�b��X��C�1@�TF2��l�&w�DBb�1by�w�c]���yȣw�i�����B�It�Sgn�#�����I�y1n/����q9ޝW�gTy�j�3�.q��X��.����!�����&^�;Γ��JW7VK�t*��1g��}�=k.OC(^�B`fi�s�rit!L��P&�g��٢ˊ8�:��zWu�����#�V��vr���Z�*�oۃ�P{�o��꾮��J������8Щ᷼2�+7�nw(�|���K�C��x� �"����t��h�'��^w��9��]j��=7�˾>���,>�p�!�����n{'gf�c�c�}�o�}��p:t��"������l�-x����T�����a�j�޵F�w&e��;L�i�Q����J����Tz-�ұ_V���N�����4�!D�0�1Qug���ݤ�s��z0��K�90o���j}�7��N�+��Z����pf�۷]��v<Ex��
	�һUn�N9Մ#��S�Q
�s�rM}�:���)\>�[���ö��t��kog��p�>fJY1�����V��9��̻����0.���;U�J%:k��sR�&{/���uf>X��9$,F�M��,����ׅ� �W�uc\�Vnߣq`ď�t�:�J����}i䂊�@'���U�S�iI�&�l
7 �s�1��)��#ݵ��C���W�.�a�F�'�9��g��CP�km�gT����&w�Wsc[]����O^cT�����I9$c\D�X+2���*�SgD���ie��6���F����c1bk\EPg�;��ک:痗���i[/x#�v�G��ϻ)RLd֏s���*���=���>�.~�^0�ٸM&�8�w^�QZvp��Tw#��K�'��8�n�n ���z��J��Hf�:��vJ+��1�T9��T�vl�/�z��l�D=͝zk�L�+�3�`���	�J�z.qR����[�՚u�Sc׉���oM�bd4z�wb����i,���N�o&�Y��#�U�
*��9��ֳNg�MO�q3�.}�㠏ɣ�Rˆ��T���q3��Bg��	D���e�<5`��h��n�����g*�7D�]e::^xq:�Ų�ff���uD��c���#w���E��8>��]+w���Q��SDn�i
4��.u"�w��]zrOz��M�]���;=}l}|��2vIm�<wӬ]��IE�ԭT�N)��.
=xsr!Ӯ�:sydpƶ�;#�p������I{8F=��3^�Y�v^�Ǧ@��zJ��nxo��������:-�[^Eu|/�P�u��a�T��-צ?{��pz'~���S���!ɬxx÷v��Sn��*�%�^��M;��ծ�O[ ���S��"����5����w5M�K���8�LH�[�Fk_���)���}�z�I>�O�jZ/e�;��9�Vy[�nvp�CP���o�/��7�}qSZ�/�r3f�vrP]��n[�M��iO��Ҿ^P�{�egՄ4�Y`o^̾!�
��e��5'2 ;f�E�:E������:�I�-� D�=�I�ѝ(˨E��|�b�c�Y�r�(;�u/R�����u���gZ����`�Z�Iީ��(� ���,�&����ӊe����J7&���4����uj$^q�t-��f{�F��j�X�k��&B��KB���>�W�vZ\�K�)�I��� ��^L�O>EL�E��Y�����,�/{���ry�vJz������s1�.���*R�<�����L���Y����}�z�z|G'����pc1/��Sy�����=Ha��aJ?nؼ{8s��5H�z[F�85\;	���+���}e>s�{.�-�B�T)��>u�$߸P{-r�.��W�l+�̏Of��J��!Pk�q�e�}�aFf_o��aEd&�f�\��-���<�i.�j�]yN��`���^�o9K�)SC.C�N>E�߳�4zw?wV�A��B��Ҿ�󲣗&���ӄ{���ɗ��� �zװm�O!����A| �L����Fn��c/����S����; }�x�E�{(t�i*�*�P\���D�f��%b&��ӔpNd����&p�{ȗ�ڳ�:��Y����v��`ٔ[xɺocw�5f�-Fy�x�=�y����i��*FjWw�3�K��%��UW%�_J�����<��`G�p�;�X�1�	���c^�i�㗻&�㽍��z��g|��0��_�'�{�F��۠j�쿼�����6��R؈VV�ZV�m�jx�Q����(��TYR���D�EJ��q1��mF���Z��
�YQV[dPV-��+�QX��
QAѵh��s.Lmh"*�
V�b�2c+e®2�Q-1��R���TX�2�,E���T(�%j��j�ѢƖ�V�R�6�-��r�[�U���s��
��˄X���D�Z��9�-��YU��ڥ�̳�f̡SV�ʩk�b6��F��ʍ("(�-�,EKhTZ�ڃKR�W)�����+Z#[�VX �K��jڕ�X�m����iiT��V�b��e-Le2Yb�m�`�V�0�e�%S��mX*Ҵ�"-�)[JT��Q���Z�T�K-@O���_o�~כ���'9Aw��_C�v�h ��-�5��\5��Y(#��F[����4�u�p^�ے8�9qT�P�L�:�U7�����yc+��xrh�o�ǜ������{�o�sc�yj�w�Bϭ�����<�m�דD<�'�ǬNY��ʨEl^0������;E�V���8�-(�yu�;���X�^f>A�f�{��l2��s���_��WH=�b	�m(�ҷQ���[�0{-'��V�._p�M������Kj_�3���x\�XfE*���;v�ii�7I�9�Mc�=�����;��3�81�﷤�ԧgH+�ʳ�}�i����5�^���˿B�-�������8~㛣�%{�����o�ȣ����g!n�,����X���ǚ:W8�Qe��M��́Ր/��3UB78��n��*�V��g&�eeq����K�W�����6YQ���{�-��˿��ХL(TI
.�bi����j���@��hM����F���������J���iԱt�H�*\�G)�[8���W)�֌��g(�b�A6�!�q�c�c�]��\$a�f'W���T'-�~ΏV�=-VљdrU�u����܌�bP;��ت�N�j.E*�^���\�S@l��hT��f�ѱ&q�J��`�����N��by�
cL�Zʹ-̪M��ip���{,:��-��Y%��y�}	�-E��s����fkm��:��q:�{��Kk�ҫ��n�>�����1S^|"���OJ��唵Ø�}���ٻ�]�#�M�d�^��>��B�tC�ٮ���ʬ�	��ЅEnA��cz:k��n���-�����V�%F�]t#Mi�j!�]j;���f�����=+���*�^��� ժ��ـ�m,j�SDѻW@�eW��f盽��c�
����ӕ`V�s�r�E;��+b�:�K�Y���N,�9v�Z}4��ң��ub�Q���v�=���mM=�������-���|�HK��p�d���`�YwV�g�r��ݬ�Psh��Y	���+��Wb�D���q���m��T���MSv	�l��P�ej�\T�1�RµH��ܳ��'FM�Z��\{E}SrR��TLf��pL�Y�Λ���81�-S\J��*ĤyJ?��ݛ�9�-��-^��V���S�9{,D\��B��)������S�J82%p��J"�:�5�f{ޕ�gϕ��9�3k��*��ן)!I5����k4�Cs@=������UTv���+1��CDUS���r�7*���nƳ�BʑC�������op�"}Q7�J�Ooe�s���5=��1،��O'�gX����p�s����tob�`��&���i�R��K!U�}��������\�1��\���14�$��n ե�y �t�p�r��xN�!;���F���k�UyƟj��ޭwQ�D�e���jh������8=�$��.�|��	�y�9��\��"�Ük>��Ǖ�WwE�G)
[@�y���Un���_���H��f�}r�F8�Ϗ�箖\�/�p���D+mR3�������b��y��¾ɓf˹Xu�l��I�]��l�/�%CŞ��E�&�	�^ݻǂ�[����\���K7;Y���*V]�N�2�a �Kus��9|4�����]�&��v��r�q��=�*��}�\�H;k��<+ke��ɦ�`N/u�NJ�$U���헡hs8�t ��ҍ͋y��k���y�����ps��5M�(�W�cݨOWP�\�z���ʕ��kE��y���J�1��]���N�z�vf��㮖F���D�8,O[>��A��犛�|�M��^˒s$�E���s9%)��4\.��J�x��|PO}��}�[Ȧ��n��m]�Û���;v!ܣ��9hゅג���F�;��2,�n��էK�����ؾu���fw��e؅ u�q�|2n�3�$�'b�ѱkx:���]^�u;;�9g�䐱	�y��gq7SB63��Ջ�z����-�"}�FcgwJ����|�^�i�R#�av�
�t�&�"�70�5{W�����L����ͻX�����"�V��et�� �zcM����*.�~[/gU�`y2�;խB2�0Z�<=e��r�"�����v>�n�׵v櫗�L��q㖨t�3��]�eG?��-���z���ũ�8F���#�c���"��R�+5n���\�u�	ع(��\z�vF�+���'bj���X���d��N�y0�T*���c7�#����5��*�ff��
̠-��t�m�֝�7�=����������)�B�LY�,Mq@45�ayWwj}��4]��w�w����jĽ�U���%դ����|"�s����l��gA��{;��o�xg��vE��챠aL�X�]N�xrh�w5�4*d�
)y����$�}E��>V��|�g�[B����/��O�&����8j���w!R����h�A��*���EΖ�Z��|�cs��UnwR���w�r�c��͊E������\�A��A4/��L>��ud�vrA���ǯ"<Y�=�֜M8�>��αL�3Ɓ}v�o'3���c�İ{(i~��q}�qMcq�+����Bh����m�95�Mau�� ���O/)̄�ُe�uLYD���"ⲻC����l
�=�/�{�q,	��lg����i��`֤��Oz�s=�l�CW�dV��{��t/Q��<1D����Mv�إ���JryD�X���:����NY�$�ǃ�.>��p"�;En��Zα����ܻ��wk�8��-��~�Ҷ��Ȯ����[���E ز'H�u3e곍����؝��)9�v�eW[\�j���09��������6[vwJ���o��Ե�zb�V���q���6�o:�?"�8x��w Cڱm�ˡ���M�Ln<ˮ�ގ4��FF$�U���r¾q�Sg�Mob��%72�Z����^�#�N��bkÛ�^Uș��&1��!���:-�Vn��S�,��pr7�A0p5&��C���7�,�� ^�vp�F�r�2z��S�.�;t���4c1Sy&�C��c�t���3���ʫm�,K>�xn�>(U��؈]N�o�����JTd�����D����hϺ]�~�0y��NYn��HaЬA��M��Y�f���w��y�PeV̓&l�e���md��u�/�u�L��݅��Q�^�K�n)����,�za��trϷc���@`�_$�5�F�MW��l��F9��Z5�,|Qm	|�aj�;��f�Ѵ18u�c�,� ��:�-P�6�fu*�9���%uo6�Jg�U��h�q!88F83R���VU��{���X�/�vf>ff�-�{�(��7sʿiO�]ࣣ�v�,ZQ9�@6��ѹr��T'վP�^�O!��CP.[S�{�a��#�*�O^ӽ (5�u��N�Xx.ƻ6�jå����$�~�==��RQ����ڨGv�4����_��:��8���<M�ރ��sj"o3���y,-�^N8"�
��΁�β[k��s	�m�t�A�3Xsn�#'�#Jṧ� �5C�x%P�[O8委Ԛ�fa���X��3��N�xֺ��U���ߝ,�����4�ED=}j�hs�8w$�<�ќ���ks}��c�#y¯s�����ʷ��3(n�~�ts#S83�U<�L��
T�P�oY�䋠P����!7Ppv�Ȼ�ww��/P:~�q�X�ϾZ\��d���}S9M)�gr����=-�����!gd�$��1L�3��]��Ȯ���!Vr�Ytb��%�(�Z����hե��#�U����8�V�֓��k��+0�ӂ��W���`�����#,���0��U�\V�M+��r�'=i%�|N�j"f��n�ũ�YT}���B���v��o:6�V�����V$���4>��5����<���ݖ�nRUc0�{�g5lB��`c1P�u)o�Ms2��c���-�nen��a�Q#WCyW�
=ҥ������,>V�.��j�5p�f(��<��Y�g!��ğ �/�'/���a���s�i�'^}��W�Z;�����uN�w��2���v�8�f��Vg�5��EN<�������E�N�ݧ���}Q\�.#A�Ѡ�%r���v�ye'�+^�s�Kg���W5��9)��q����d�_QA22�u,�b���O�.�G5�w<N8�5n�ܡ�<�R\pDJ�"Q��8%�	��ٲ�5,2]M��<M�N1���^RWV��?e������WOB��ygl����K�{��RffC�E�hmS	r����T��+�.kE���׀^�^���E���0�����͆���w��[G�5`���m'����ޭ�i���4�w$6̻���4-_���H���I�+뽾b��`����,�N�V#@���`+�֪���A�SO�ql
�&�aH��g1���Y�@J����7��զ���O�3tpB�:�	���H3V�mع]�<c̡=�P��w��L4������Ss��Eȯ*�C��x(\��>�[G�F	o�\��^UҾs�r�7�CH�v��^��F�&k-efP��t�c1�R���܃�����)�;b8=F�	0s�ŉ�q�׳9n��(�5NNw��
;�r�m1��`�R;)�I���fh>U�q����r��.�4��ʻ�*䝻�y����B�t|�i�C[��'��tοF��z�wtcq�Bw6����)Q�,�hVo����O&�P3�X�i��x͹�ʽҷ�(�z��<'��2k�~:��\�)��%˱���Q��)����B���w���x���K]֛˞4#
w��2�uz��۝��	���ܶos4j{E����,���+�w���6:,7s���m��:�y����?w	���ס�eNJ۝-���;�0�r��b�żƦ%��z���7�F�͂��s����'�s���w��Yf��Z�0�̥�q��׵4D,x�)�i�3B[Sk<U���{����z�g�������֚��WB�'
�F��*� ẜg0Ќ̻Y�q|���O�uwG�d6�]�]1v0q!�^H&�k�,�@�v0W�t\:u�e�q����8�w0����Ui�����=O��x-��� j"_��#s����ү�ݖ�[�rӬ7��(��߳B{�\P!c4EMᬁ�d�D�{^�mD[��O{#SMT����T^\�����P!"�B�s�� ߎ)"���޻���72�:�,z6�Xmڡ<�0�����r3ʣY��� 
2v�&�i��><9eh��ycJ�
p���zd�V@��Η1�!G+��z�sY�T��޹y\�B��4'/���vֺ}�x+��;��jM����G*w��ÂV�	!���BF���b�
�2�Tz�囹�`õj��1�1�{[���6�p���+NKg'^��A9x�)j�m���|l�pN���x7��(�v��\�EV�ٷ��A���OgRԧv��_���k5T��gg ����ɦwLO[YM�K���Y�����*����'p�g]8�Xb8G��8a���0�������eN(�����K�F�@=-ʣ�;t5$��uX33����5	n�(��˩�uyK��)��x>�4�Մ���M%���(��5��A�y`	wu�dt89�<�F��
n�[�#��r�f�tk�e�z�	��`-�GVK���8"�c���p�]��b�3x'Pu�^���#��sCeAV��ݧH��3Q�7*Dp�n�y:� 'FCr��L���-C�}ȿ��ȵ�E1n�f��o����<n=o�ަk� ��{єi.i�<%.��|s5K�^d��˨Xy��T�8.xX�V	�s[���R8NE�U�(�V*�����*���|r���;]�JWU�rF(�}+w�:5��b�۞[�ͯꟚ�qk/	�����+d{~BPw.0	D=ׁ��vOv�*v�_tPu)dX��1*�zƃt���^%6��Zm�Ĉ�v�Y�x��3�r���x⾣6�=P2�lW�N��GFf�[=ٽ�ʆoup����++�6ʤ���.��3�_��`W}q��U#|��kh�|�Л���,;�qhW�ލ�3�%h�غ��cy{�D��\��U-��2����ϟ�n]��im�5Z�dWbi�{e��fX6�-�k�
�ΐ�9�N�����Eol뙖����@8qt�����0(��X�	�zȩ0��*'mv�_&ҥ��0�f��_POID�l9�'w�Ī	[���&o���Α���>�D2ۊv�O q�>���{��H`� �/��w)ٗ:sHCj���ٵ��v��u\c=��ho@sldz^ۤ1h�T:�����.��͘)4��`�ٮ�k�y�/��,�c�%�Z��>	)G���&�p)o9sϘ�{l��$9�u��8ۘP\��6�!����vc۾��� h�t��7n�1��p��������FRY��P�8���0[|�,��紭���(�VI��a�O������W�L�zM���6]�t|�i:fjl5�,f��-� mޤ֨osm���U�l����<*�s��ǻ)�N�=�	��j���y�:�W�����+{���
ڲus��H���~�T/荪��֬6��AbR�h­-���m�Em(��"��)KE+-F}L2�e�Q���eĲc[h���l��Jb�Q��m,�R��V�-+hUE3*!�c��(��%*��ƴiR�-[A`����FDe(�`�*�akJ,Am�Ud�2�UV6�#l�U���pʍ�T*ZU�U�iF�QQA&%d�#Z���*�QP�0�h-
�j�TZ�%2�V�*�V�����
`�B��ZQ�k+iij�T�ԕ��+#iRڲ��KG��iYUZ�*�s.TB�Ԩ�E�4mj��\K�h����QIX��-�m��Q���*�b�l�R�VEh�0�
��k��La���mD���[�b�J%��*Ҷ�X�J�F��b2�Rڡ[mEm��,�YJXQ�$j��T1��`��j յ���Tb�V,�b�[B���(�J��.��o5.����dr5�j�n��rr��U�׹���<V����A.�/$O��\�m��ұU%�$�I'y)�A)�ضh*������!1mA�&2��Ҩ}��=��*���9��ɻ�v��Urށ�H{���5��s{r��c³R��6DK��w
̡v���ϲP�lg��	��j��uU�|�8�˽����h�W5�qZ㦥�݉ˢ�t�cB;4�j�5�����x�����W���0�Wz�w�ʣ۱JV��N���S*�Bnm�pB�:�E�y�5O,y�w��1����o�P��&���o<.���O�ok��ЯW&"��������Ӥ�jf�d<��i�6uD�u`�gH��������m_�-v�L��Tr]s�͚���:cu���ȕ��OOk)�v,N5�-�ؙ�Ez��5��א�x-���2�a�E�5�����3���`ԑ���4��e����dGx�L�4������c�E�(X���A*g[��׆���o����D�n�h��T
���g9���7��P�]0=��Q�y��rj�I'�x����1�v��&��ˬ,vĞ9�n���t�3�����pDv��G�LZ�8��|ѥ~�����5|0�UQگ�t�fvc���{��&{/�N��O�5cYɵ03����,����H�NrW��j���� n�"�Оo����0$s��#G(hI;Sqw �֭�Fءrqkpe#����	�<�
�������hْef����ת!hZ�֪�.�g�����;�!su�y�8���k�HS�x��u(��7�g�*�2*~⟟'i�6PycUM0��g9�����X��1y�\��^�Ϧwq�2���-��h�U��N��tT�R�[�����tC|6h����F8ٿK̷��/��%Ѷ�r ot�ɻ�A�a򷫩�94Z����??Y
t�ᾅz�R�p��}}�z�ˮ� �i�C1���7C�n{U���|c�-�͠8=M"�`mosŰE�:���&�i�|*�bK��&��:w�Ê���'v��i	}���6О��v�C������6y�-*N��Lz�"j��Y�=N����`\����ns ��nj�ID��S��1ه�JTߥ�ҕ].�.�����N��0��r�CNpy�*\��h���pۡWZ�6����Ҙz���J:�K����s"�zo�3����_J3s7��K��M��l�ph=����ʎDJ�x������\�tw�aJ��x^s��6��;�@�ٮqȉq�]�Q���n�ONλY��pyV?]^�^��s�n��ܟ6̻��W�Ƅ���WXQ�]��r�b��,	}G;�^�u���z�<���hM�=���{�����-W^�W[ƃt��L-G1�ݥ�u*�[g]TO8l��뼫/A��]!�K��@�2��0�>������Q�"�㷰sz9R�޾��Ua'u�EȠ�gq��v�}�W��X��x�^�<��e�J�F.do Ȅ�s&���Lkɚ�X+1T��]*0p���S�-
ǧw:��s�B�$��R8��a��[ƅ]��֚�oe#�1pض|�aN�K.������%	6v?t�^%T�kM)��8����%`�CB��5%(�JŞ�����x{���m�DE�m#��w�0^�bvRm�i��r�����y�	1g��5�qA��#�r�?�Wv6ؖa-�1�^ҭ�u�-�8)�D���S��U��HV����GJ�7�r�;�r�Ivn��\(al�,d.�E�ɬۛ��/{��Vr�u�D=��>r����7a����;�+ټ�����DK�8��:ˮ[��ݼ�+6+�^�pjvU�YH���xZs;6U�'�[����&�ں�+��Ӌ7{C͊E�����֍hyV���\.�՞��S+i�<�Il,x�)')�i��αL�W9w��s�qo7+՛ӷ�leԚ"�$����a�l��Ҝ%��S���a��v�k���B*�E`M��u{�����]�k�8��-��Tc�4a�XZ��{��D��R��:���B;E��(H�z��d-���WAb���26!�#7xh���ȉ�y����y�I+q��Ն�Iږ�R�ʏ��� .ߥM;�������=L%R�m��y��L҉�u�,Bt��몁6B��0��3��/���t�0���W��i(n/�]k�����:��2BY/8q�e���מk���\��DK�MUxF�-�;�t>�"��s��u^jZ#x9�X�km:��,f�4�5�5l�����d�W����|�oE*���>�]��y3����P(��{�n;�}]Qj���g�A�̳sj��گXi�ک���v&�7"��5ȑTT�-�m�������d��k�
��e��ad&-�"h:�A����(�W��x�y�S~���֮���Q�l�n�#��v1"h����8�r��R�Q���&^�C�k"gwVe]�"��C�24��
�t�f�ܻ7�j��[�gS�������mcJ>̞�Yj����&��@Ϟ�z��)l��x"XϗS����jٜ	����3BWu����m'�GO]��Y�Ђ�J/�X0�^�a^r׼��� �w���.şjlZ#؆;B��q�A
���o(ۚ5�(�^�m�{*q�^�k�_���k:SC���m�v�dC�&���{cb�8s�X|�C�!�f��wi�҂>m�Ѻ��n��Lf딤M轖�|yg0YyԹ�-��������Y���G�P���O$����N�~A�v����0i���>�Q�K"u���>�g�=l���.�O[m[��g{�d]�%�;�����䔦������TpDJ�x�/�	����j:�ȳ՜u�+�]e�lRsr��n×��кk�c��.��<֋+U��Ao�{�pU�}Ȕ`����Lk��1;��S	�`%��C�}*�d�k�٭#1pb��Ɍ9�~;��v��>���HI��~t@բ"��=���ĵ����-�"c;�l���Y�@J�֙���E
5<�*R�>��ځ�y�IM��EB}���p:dv�soaՍ��Գp;������.����+j5C���.A�4@��`��Dr����#lbۦp �9�ްX�VNl��z&k-`����Ҩ���t;�;gtiU.��Ww�/)�p�%�z�6� ��<�΅���I���t��j�s�����['��Vn�]��?	�{��d�%��x��v�����`3��d���j6nkˤ:+�5vf&:� .H�ڨeK���</u�:�Ryd���Pf�E���!5��`�|"{�k�ݷ��+�k5��TV���A][T��V��
���7�&��O�Uq�C��P3���8��DN9�ؑ�qͽ�(aA�X�]O���M�/d�y!M����\1To��+��²�Ϗ���1���Ѝ�v,�Gj�E 3HȚ��jG'��qi�SW�\���Ь߫)\n��<���n��u��C'��M�����˥[ފ./JPrU���nv�A� �9;��s�(S�ν|%�6�k�����Ol����p��QجR8���d�FM�d�^pBP=�:����,�Qŵn��R�|�'8-��#�fs0눷o9��b��{��uOu���}rCl˰!t��
�,��g�����j�kb�9�u=��k Yz�u��^���!b4-���p��9�7��Gh瑔d�9j����K�h	Gc�y�Y�'���}�`i���X�1��
v%e��c���~q��5�Uz�t�5�������D>��OnZ��y�i�m�oKW�|���}�����7G�;���I��~���pu��f�W�sY�O5t��zR# Gj#7gt�]zU�6�J��T��Q�M�w����j2)�:d�~�rq�����z�H0vNó��ƕ\��'S��*�@i䂋�^U
��� ֩�n�X#E���'��eT �)ǢS=�S�"!;�ŉ�sr+ʣ\D�X+2b{�ȥ�����2��]��%
��o0��ő�X��+�k�]8��[}�P�+;�2ج�k�]d��t�d�I�����C����c��}���#��LfaSv�������-�䱮�GCr
�vj:�Ž�����[fX�#hk����u~���7Hf47٨6�%�%@���ZBe�-n��u<��f���ד�ӮԾ�����й��.�mn�=
�[L��,���-8�[9;�{�EE�NK�~���Y�D�*á�b��s�f$*;�����̣��\EqX��{=����Mwp��uJ�v�5���g>��W(�ˀ=J�_)�+�hޝ��pm����9�n�u�]�Q�Fe@� �.պ��x��h�)S.�-���Iى%wl%w�K�3���{Ե��oO�H'z	G�����C}	v�Tp���B/��18p��G��'���G�ܕ�X�9�~�ӯlA��6\��/�Sgr%�98�=��E�7�+���Z��!�ZY��TE�����&�9_I�����2�a��͛+U�q���2���G+����'7"���b�\!���,�����tQp��d�:��jx'F����]nD��d�d&uϬo��g�|T�>	�]���t,}����)E�eCU06�n��y�#FO@cgvB�d�����,=��AHq1�s��ޔ3�k ù\�\L�������p�.�"N���(O0B�L�������DE�؜ĺ�������$� H��LVJ4����|\��C6e�p<.�Sj�uh\�OHr�����j��GR>�9ԕZ��O�ia�6͊U'4ƝYC�2��SP�axy�����7o�����zSOc�P%��>��[��sS��B�a�z(���+�,S��׮N����@�^��5F`W�M8�����]���z
ESŚN\�c��Oؤ���p-.���+�J�;�U��]Ҿ%e>�5a�������Ѽ���4�:���4]{i��=�-ӂ���0p�q�x�AT�[g�C�v4d���;��Q��Ð�z)MC�&+}��u�k�� �9�b�2%�I�﷬���YݽE��J* [�< �0�������"�Efⓩ��qF��K�d�q٦.z�j�s�o ��N�_�;l8�a�0�1�����wC=�]���k����9N�Br-��ח��:#/�v}J�1j7���83��0:|�e<X����R��So�����3�w�����yw��X�Zև�b��2��.��tZ�sݴ����ϛv�OT��k;���Թ��ү�n.���v�侠��~w=FLtػ0���f�/��6�dU���2�2�q8�Dpj"�OG<Ĕ�As�t�T��Alu�.�*���H{Ga�
z��ԯ`bl^���n�D��-p��.�X7��1L*qZ��F��~�@�G9�����ZK�`��FɎ�:��9s�.,�ݓ�T�'�ٝ�$n(Zg����W�?N'���s��F�u	z�M�*���:�Gb< s������%{����n�^!�6� [�q��	ҵ6�Ӊ�u�[�|���a4 f*�� �MN�6��<��! {��<���y%�0��G�$���l*�g����<�.`J��P�Q�QV�a kZY �7�_r�w�s�kb�̟Ҭfo�e�/�������buj`殷q��ܘpRn;L����1�4�%�7M畏N%������t�!�~�ɼ�HW,�Z�Ik��bnNz��-�O�I"^ũ0���]�JYN��r�vAҟ$�z����/;��S�-��Pe��sr}���Lc�{�6KD�V}�˦��Є!#5K1��"�@�G۵�HŢ���]��'��9��=�����j�H�%VR��=L�=�<�G�U�=�e)��^�
q���+�u��՚FU��[��gR�`R{S�j!���ձ�^�t���=W�c��{C��1�y�}&E��]FlCw��v
��Q�˷·T�����N� 3�Vi�%�B-����`�˵��o�5Y��aL_{��P
ᙳm�܏'�}�橃�������KU��{�Je�t����"���QLcOw�|ū�����.�|��%��I�T���an�#�� �Z���:�n3���/۾7�W�<�~M[���u~i�Ue�C��.���ǆ�e�n���'^�K�+�"��5�u��47�gzй�o������>�G�K=B����[Z�\�<�}�*>��,M*��f��gyw	NN�#���(9f>�΋�}�$��@���Fs�_BD�����}#9CD��Of��]_�����hf�@���c-�it~9�=@���-`�a)��ϊ~���ͨ�Ķ��{���h�Ҟ�^Λ�SG��^:rՆ���Qy�2�kH�ݽ��o�{� MZ�\��M2�µK,�K�BB(uNǝ��M�7����u9+Ǝß�3V@��v����r���Ŷitt�7Y����FA��9��[���fwY���0���4(ȈN�wt[�a:���S:����_�q<հ4q¯*�P�Ln�mҰ.+ށ�U$y��m�Z{EDqEZ�af�G����⣂��C�x\M1�k��ɇw���R�Y&MGǹ�b��We�,V-�\�d�[��#��R�X�R�0n��r�;�?v�	�z���W���\2��h�݌(f򺃟Xc�����{z(��`z�;5A�N�K�ڔwy�DE:�Gk��kwhi��=��vs�y�7����boY�6;�w%y���d�cEN;����ٌ��ؽ�6�*��	��,ͧ۔�+�gj.r]Ʈ���H��P��vN��u`F�$��6��Lk�6�&�.����(����#���7� ������;�D��H�@�'���ph�Oj�k�r;�wv_t�:.���&��B��(���e�R��-#eE+m�[i�bZ�,*SX���P*�V�JZD��dYm*�V��ڵ�*,�b��*Q��m+m���eh�Um,�i�eD(��mjUQT�(�ic��UB֒��,����F�kPe�����kkm�!�S-X(���,,�Q�mT����.3-�
1���!RT���Z�eQ"�+�F��6�ص
��D�e�"�r�J�+��G�
��ZYP����YYQUKmJ2V���Z6"61�kd��e�VTX����k�P��al+D�G,�+m-��-�V�
�֕+*�m$���TVѵ*J��[,ETkb!
¢��ذX��&(��QE���(�V([Pc-
1DA	Z�XԪ��-�ʭ��ZZF�W(a��3�n�<��f���_3�j�ZҾ߸�ջJn#Ux�8��Ue>�΋��	�g8per�Y`�y�ng�^<�+t�m�3z����;�Y� �R�#�\`�r����Ys��<�oyT��k�]�վ��&W&���r@��XC�*�>3k�3���G�b�~��'�M�w5��p���k2��S��� =�8�WN(�St���DB�y�EO�������]�X��I/���7a��R�ᣕ�v�E����kЁ��To|�$�a���<���/zh�
eΦUK�R�&���QL.ڭ�0MB�o"������"��E��`c׹��<�8�e)�{L���x�Q�3c!��9A���\�{�!A��ž1�F�;D3芊Vԥ�Gً^�[��Ny=ڵy���z��n��lXS��Q�VI���a�T�ni�C-��� �hO)��������K��9kwM�����J���J��79���fH�bn+�o��sw�	]�V�ϫMa+�/�<Afٔ�1��r�oe(�'z��3�X�˹�yOw��Ǌby��ۭ�2�,���T�|TI�B���?3�ut%P���Ь����М8o�����ʣ�V�V!�o�Ow2rHw�����y�֛֭{d�
gJ��j�X�*s����Q��*10��"�������J[=9f��E����4��8�*���2����'g'\j=p�gA�C�w�b��H��jƲ0��.�h�^�Pֻ�vXz5N���=iڊ"�
&#�W.L}��u;�9n"�Bzi��w��I:���0��*�W�/mT�n�s����B>�Lʗ�q\!^t���:���׮u����a�� W�S��9b���BS���oH�Mӹ���ؘ��9�Bz7vQz�>�s w�"lG1\x�W��{
��>f���	]���5�ء��'%k��;̲�!�W�u�)x>���g�@�)?:����h�7=r6
�P�g�����j0��6�^�{T,d�1�R��y8!��:�<dYU1|�,�Y�Y�"��w��4$�.�$�bbϪ:�%��u�1�L8�Q���}�Q�WȊ�2�u��m�ʨV�y��Ɋ����5ň��e��`-��T0!���������qSCrs������z*���7��A��@C�C��)B��d� �Ns��ǆ{��ǯ�Da����)0:C���]���$��\�'�)��:�m�:w��ZS�P��<6��8E�o�<��#IS������ތ澚�b���՚H|�����|�����ON��:�'^F�d���Ĥx�Xo��áT������Xu��L���ڳ���`YEc��g�v鏠����:��໲��b���Ȟ6)� ���q/x��X���/x����}����-�r{w�W&k��nYA樏�������i	H�/����4����ۈQ�������4ˏf0'����T2���������f%N�ѰԪF�s�Ua�+�+h��`�����p��GN�QQHS����خ�k�IU&v0'v%�8j��E�B+�2�N�F�o>Qib���8�t":
^m�Wj<ac�R�z�'}p���G�}Z[������w����O��Z\C�ZzvE)���T���Bw�U�4�My���k��5h�˂�8�-r�:�}�(t;^��T�w	L�1�rQ.���K�'z��[�^�\��t+�x=���π���z��*��\#j�s��ҍY��ވ\ܪ���̫��w5��.�Q�� �a���g���D]�U�,��i���iBA��Β����z��e#�}cY;SaK�VP]����>�Βۀ�o�&Q��q�ξs�_;��常�	`93�"Rx1N��,�6Lі6���V:��
1�])�k�x�b�or66f_N�yGM�\=0�I�.V�YJr�(�آ{�^i�����0_ܸh7���+r�4qK6x�;N���Ww5����{�*�\*�(/��}��4a�ݐ�Ɔ�"��������
C��U�nvM��ݤ;��k���Bj��T�O�;|r��M�����u��R�`�p��͝�3f 9n��}�kG6��D4�$���H�����le;�~ꈦ���UD�;)@woaj+�R�y���3�cI	C"�3�ia�6͊RsA�ƝYC�3-1��1��KJ��&��z�"�P0�/�m"��{�>In�R7e�­�[�FY���y+���
[!�#���!sQ��&+�zs\�:����C��ކۉ�p6�WQ��}�m0���0�#�i��AȽ��T�>�6~u�	���>�� ��NpuoE��=inɩQL�aE�0� ��� ���9k�����OK���á��tMr���H�l<ثٱ]@�U�z���>���ت�Z��͚�P�S&�����W[L���f�{����ҩ4<8V�a�^�P�F��P���x�]B�<����W�f�>"�>�c�Σ���z]�\��gޜ��}a"A�E��K���q��Y�h+�^�sC�o�F���1���H�z'3�iW[�R\����	�w��챴�F�]e՜���ۤ�k~*����x� 21|0Io:�C��(�,�-_u�V'�{	��}/�temXJ�Q��@��E.�b��"�{U
[�[q�N�w��Z�uB�.�]ԇyFu9���,L�K�D����:¿
f`eG�*P�<'�]ל2��α���r{�����s� DtV�ɝ��&r�Ӡb��G?��P��1��$��[��y�r�bC��FWGE��p\�K���:9S��ftbFⅦ}0�<�Z���y�V	wH C�Q�
�����ѿJ���U�\�2)���20D��V�f��W�,���/n=.��Ho�X#�7Bʇ���x���ր�>ϵht��2o^d�vxKz�E�
� @I�m]x*|��2��ӂ���:N�������0_��z�1�gy��ﾌ�HC���(	�s..у���Q��5�n}-�8�u3����bS���E@���&�� )ň�I�d� ��")V�>�ǘ|(���=��_u�,�/Z���kվ�FE9c7�B�N��Td��E��DTv#g��/:36]���C,T�s�:�\�/,n��EWDouԅ��0��P.]�+��sT���#}Y�&�f�n��*^��<�t�˟�_x��7�]�{��<UŊdW�o�!��8�|�z�#�Nb�)�a�nvr�A��D���@��^L]��p춰z��K־%�4��lX�ݎΣ��9�9Vô��܍��P�n�"eu8�1k愪;�2e����L��X#��A��DG�^������"n ޽����7��u�:ˤ�r����f}f���~��U�fٟ;Lt��(G\��0����8�������I�D���=�'c<�=R�R�^��:�f��T�t+a��+�P��{�UY���0wj�g�ʎ���}��8>u��yI�=��:����i�����[�ns/��^>��Z�Qa�z�R���.������ȷ7/�AY�h̩qDlm�����'1ޖ�6"�(�C=�UvC�KER��CM��O��t��K�q��&n��=�iz*��洢$Δx~Ha��`�a� k<hXb�.C�P65�^[}�b���/jޡ&ŵ��wt�W[�/�^J�Bt�O����i���,��Nƪ�h����`*&d�|�`]K{P�R���u��<L��.x�J('2�:��Mz��L:�:�'f
�
�u�*�����	��[�v&�����B���0qK��&tom�m��nk�.M�U���c�%�
�	���ܐ�"���˙����+�Ab�ό4�i�F4�^���+��]q�xL &s�grif��,���Y�_> u9h���E��ǒ=]}%K���Y�T�'..Y8"�L�L_�ÏPUS
9�9��ɺ-�	
���i'v��U��h8#&*S��`���x�	͈>�+"(� Ll8�HU�QWs[�s�Ƙ�X����Y�J*4_Z�oi܍���us��(�Jf2lB� 5�=����X��w�zk\
�P&ަ��������>
����δ�*�e;�D�ѽO2�3��2�f�8�V�:���>K��x�^X*x�\��u��^&:��"���^kA.d�L���B�f�c:��YF�絜�hD������i	�#l׼`��u
���/����&o�H���*́������.�����y�N���پf%Dh�j�5r�5��sY�N`�i �q�2ͨrvC�D"�B�v607gb����Fnv�Y	X�l4�JT類Bmb��L�0n}�G�#�B
^��+�":�9�U�'�;��.��шK%������}�a]����2��h�eZ\�|��k�vGAS�"��`(T�ö���O8et� �V����Bҽ^�ȯX���u�k"�Ա`��`.��vr\�ٳ�uYJ�
�G�����$6N����If�+Db�xzJ�
��<���8;��1�qoI���8[�vL-Ǵ�b=���r�˷	]��bAI��A)�e�-�=)E! �Ut`��\A�A�����I�]�����o/��3?뙇�X~�Y�T�E�t
[�N+�.�"�6n������M�
J�V�Ɍ}[��e=�j3���CYɞ��F���U���pUr�f��E組�T��A_8�2h4�����E(s�&2&NCJ���Y��*�.��>��8���v���v��L����'�q��V' ����2}\��bvtE��6(*�X�=`Uɹ��6m��<j����?�_?	[G_)�<��X)|y��L��s�@�Si�jqE#� ˸����$�f��C�?'i�rס� ymx���P��F�#�j-���N�7��u!s~�S*H���
`�M,3���惡��Ӫ���U�U��-ԣ���E�����
c�����Ԛ/�H��|�ϒ[�Z7eԕdc�qԓ��ս*���L�!����[*)�A81G��׵����y�(:^׷�2��`3_�������"�\���,�Z�+F������|v��s@��f������!h�X�䦒�sp�+�����6��GxF&�i��+��x��[�f���b��{M�w���J^�ㅨ��a��U��ޭ�˓__-�]H�@�q˚�׉�<���[CD#8�(�}���u3y.�������(�)�X�������sFD}J[�-E����Ô������^P#���5���٢�'yfclT�܁���L3��LZ�ކ:UYXOy�ҙ̧8���"� �x��R�����'�Ho�Wi�۫��S���X��Z�\ٺ|n4F
�p�����U{esl��"��z���3�{��v�g�+e�� �;���~bx2_���,0���:7B��I�mnhBP=��IRr5�F�2
t���z���c�+��
p��q=Lg����a��iF��H��z�.u�#��VL�^&r�Ӡb�T�΄PX��̲D�v��wCqlQ��+}#��NÍ.�I��p�dn��*p�lΌH�P�Qwi��$���yޡ�l��	�x{���]� {*,E�{;z��C4���R�Y�]��s�,f��!��[$E�F���,a�[t,����6��>X\����z�
xaU���I�.Q~��^׭<���Ni�$\���*�H�r��9N��w�+-�v�L�yHfK����{�ĲͱT�I�*Y�������H�E}YB�ty�KR7�1�=4VR'31s��N�Fm!���0u�X�R����ѭr�a�ƶLU1͜l+�
0yM�u};=S4�(��T��yk�Y��湞�ap=���	�1��Bćsu�hs..у��RO%��s̛�^��!#����'�g�U�O	nlP���x�&�C�%
^�DR�#��泗c��0j�8��.��u,���[}��l^+>�2�Y%��b#i׈o�l��E�5��ÝGy9����x^t����`X�X��X&]���Ҷ��tpsc�l;J��ȉ�"3"��U�cr�;{G�Gw��C�SUB_p�Y�2R�x,��E�E��#O����P�}/n+��d��X�z�>��ߵ�u8��t����Y���Ͳ���e|��P�-'�rG-����[)��r]R�R
,��������=R�R�WQr4�f��_U{Uu4vnf ����IA��
�cFϏ�����-�v�F��T0�WzpN������W]}*M�g��.�=]ND��TM*F
���k�7Z`׋��?e=��o��m��엤$�	'���$��@�$��!$ I,	!I��IO�H@��	!I��IO��$ I?�H@����$��$�	'?���$�B����$��$�	&�IO�!$ I?�	!I��IO��$ I=�$ I?��d�Me��4�kf�A@��̟\�{��QB))@�!E*�DU*T
D*�P��R�DTJ�UUJ
	T�B**�*
P�
B��"�E�Q�D�T�G���RB�F�U
��UR�QA}���$@J*Q		֊��E �U$D +Z�*�ԡV���N��UJU(%UR*��l�UB���
R��R����
$D� *��R��B*�T�$��IJBR"��   ���3`]�9�Ѧ���3��a]��\��]�ݲ�����: )��q�u��8��4Ѫ#�ZGS�]ڍv�iN�8�U5�])��T��YB�I��T��  ��Ӷ�Bt�mv4k�S:WB�·\-�tҚ��.�K�m@d��]]ڤ��h��uv����I�V:����B�b���6k�I$�`�PRIEI�  ��jڔ���]�ë��1�1A���uɻ�t8�]�W9������)B�M�QEQE���(��F�(��.z(���.�PQEP�THTN��٪��  �E 
(�ܫqE)"�(���(��M+��9Ѣlu8�NGS*ʪQ���\�TUhs��ճ�Ƥi��2UEP����RD��Ux  8z�Z��r�Zڅ6� �5m�D.��A]�U����(�L����f�(�ݖ�� �:���4T�� E%Q���x  6�QOTi���Ӝ��,�ʘ�snS�N�6C���2l�\�E]�t�b�J�*l��3AZ��i]�;�����H�  ������t���r�m��F��iI����v��2�R�l)J�k[CFJ�eYZv�Z��f�wk�[n�v�I�Ͳ�ܴ�&�.�U�EKlK��!P����'x  -��[�4��kN�[v��*5n��Ew!ٺ�6��j����.�D�Ԛ��e�n��ݖ9\���p]�v��tkYpf�
t�P�m(�JED�S�  9OZ�ڻm����]�@����7A�]�\ꫝ�����0u4t���7m`��5ѧm7R�l:N�n�[[e���wZQ��mҖ]�`V�J�UIE�S�  ܽ��v[]�f��*T�cU��8�v�+X�@*��m΅��펁������kvw
ˮ��N��"�)�*릻�h����@eIT& CA��$�%z�  j�b&�U@ O��Tz@ "�#  �1�JSM ��U�"ٔ��bfv�I\�(��f�E�L%��^wח�u��W��7��"�
�* (������Q���+
�
)���Ӈ���;��Z˽u�u��)Я��.�]`�)6T�VAGU��ĳ.\E���is5MT�3%[��*��ݨ�5��Ќn!��Q�hY(�6J-�f�Ђ8�Mȃ�%C�F������t��ęF� L1,�5��������,ʊ�	�^aJՌ$�Sf(l�J��4
����0e!a�u
�7"����5�p�X����Z�v�C�x,*ۓi�t>��ʷ-��X�Ж�)�`e�Ы�fZ�̲F6�H�q��ݍ�V�b���Ӎ�ǁ�uX���6+n�ݼ�1ԏ��l-3�N��sP�u�T�)R��X)��n���tI�$��kihB��:����.�ٌ�Z"n��o�� ��CKA�4�*'�Z5�k0?�Wm���a��;�*�����ل��CHU�k��b�n#����0Vܒg�37�yb�]It�Tn�Ԓ� S!F!R�*��ou+v�^;�� (k�*��HCZ��n����B�v��٩������74/+Et-+�]��<W��nQٯ^Tc[���1����C�X�,�QZ
�*�TD
�wb��=׍��s^-M�2�������fxsQt2b�ce*�ۢ�؛,�aV����iݭK�Sp�f$�Y0V`:�K�[r��ӂE�	H	`�h7@hJŝt��NԨ샎�	�z/i�st�lX���Y���z3�ƭ[D1y�bɊ�r��T�,h�Y'*�Qz��[@��1���*b7Gu�*�b4f�#[X>�6� �u�'t��vK��z��PU��kX�Y�5��5�Y��X�F),�&�2��duCN���E
x�w)�YJ�5"S���Q��qLF��W���"��`�X��Z�B�
Z6�@1@^6�C��pp����*;��Q����Ub`�/#�ي�1�˴���I!/1A1��74��@R.��Pr\�̭�T0�5$�1�[ie�tM+x�6jV���n��X�Icl����5�3%�S�����C,Y�aU}0�"i�z+G#kv�e�؞YgsENZ��K�{CӦ6�s��"��-�E�n=�Ԭ� "�9�Cm���*/Tlb�����>]X1p�M.��)'F���U�QY���w�[ڽt[�;����t2������D��m+4��( R���z+��
��1�h&U��o�!KRX)B��֍��@n���!fT��w���-�Ł�ޥ�˩N�Se4��]Z��\�r��)%����tR�X��f<�	�\ww�����˕�59�YRt��x�b�i���[�F�y�m���):��6�Fc2�:,jZ�����@ԃ2��IP̊�&�`�EeA�HV캶�6�֧yZi&�e�-����I�r�[��2⛘�]���yɓe��c��N�8�-m9��
k4�
���\�V�ۅ0���P3�^֧ǚt,Ƕ5e�6�,2�03L���W5X71l�X��Gk@�TՍ�*5���h7�� E,B��L��	K ���9�c�9-��V��,c-e%�&����R6Ŋ`%)�d�J�9��`�G�*Eck2l�iVJ�7f%f̻��KCX��Տ4�t4ܦoYt�5M dʱ.�(7��Z�J��z��[F��Z/1���s� q�����ԃ��++2}�$Ғe�"&�&ۂ��r�8��S[��j�(����)f�b�w"����(�y�e3��5��d�l*V���_�Ҿ�}��ډ��ZI��ifT��8d!���
 5��v�[�D�	�րN�{�^%<:�{V��.�٨�لJcgB�X@�׎�|6�BPw���|.�#T��Ԗ����V�1�VfY4s/@��+v�&��CF��R�)�z�[ �C7f����0r��6j�$[zN���u�'p� kQ�X�IQň��H�h�G�E��T�<Ssa�,6
2
�H��9N�����ձ1M�X��.�Һ��2��*����Q�饁-GX��B=@]\7A�kv�� v��n�G�dtc���$-����So0��ۖ�Y��Ǣ#����aQi��%"vn
��,-ǡ
wo(Y��XRVn�����U�ʹ�n`ue�y�@4����[V4�4a� �t���Lo�@��n��P�:J�i�sX�cn�RԄ��hQ�n��r���iKh1�r����<08��x�c�%�3
��R��lm<j��RI��mhdU�f��K�
y��+�yt2�4��t到TU�[%*u�SOn���������3HqJ�⡕b*bU�����1�EE���X��h$YZ;��h=���p�{�uf�h-��fn�t[0�u����j����Z�뽆e7� �@.�	Tz��u<�Y�G-�,��
1����Y�y���V�CV���N0v|�y�v�VEṩ7�䕕�SJ���vU��Poy�;�r\5jD�֭u�Z*�ҭ��=�#���v�&Rx�`2��U��Ϙx�{/h���bvvn����+r���edgZ(�oj<����C�Uѵ��n袬w�6�zs6���2U�s���P�oS�E憩,�BQx�Z�Fc&T�,��L�-#"��i��;Vt�3��,Դ��NM%J
s5)%e�ֵ�Ӓ���̩33b��,�T���:��=��k,��U<Cn�i�2��DZ̧Z�E����A�`a��/$��j�����+���K18�!\w[��V���$	���8l]��dir
9Ȍ��4YRQl�qD�bn���{��f�ӭB4X�)�lݼղh�i�([�(Q����9l��y�������[�+�7x5҈p�� �g^��t�J��x�Ӵ�a�I�r����lNƄL��1�����X9�\�+@���+��k�'(�n:٪��2k;h��˺�-�A��6�X��6�Y$�D���cɚ�e
g^2��?j�ݥb{��@yX�=K(K�%�iK�l�dU�2(�Yug) ���,6VYwH�%��8ڦ��*����L��T�F]���X)��[�$B5r�<eh�g
���d�o��2ھ���K�F�I�Kf6�a��y3)D��ÕE���áB��Ȱ��.փF���r*�J�^�1�c11�q�Ҡdى�Vr��G"�Ovf�h�L�n��E����c� �Q�4��.��
�i��i�Tf��[+*PemMû%)-��Hի�A"B�ؙ����Y�-Т&�e��Մm�7w���8�V-��o !��,5PVŒ�E�7����ZQ�������f�
�XdRƍ^�b�����-
���3F��au�L��j��+i�����u��F�:��nD�����<�[8��t�T�А
;��-�d��%mV�$	jI��x�����N�L�	է"u����,�?���h,+*�
�c[%⣢�
mV��!0�m���dy��!ͭx��/-ցA)-R��(6�*���2m&�h1l,ݚt�h	/-�B7zQ�q�	��	�P�N�6����x%�&��Ԋ�{v��KU��Bw'�������n6�=ON�6R�0+Wf�@��ksJI�V��*�02��Z��)eff�M^�JH�� ���g.��ؔ��%�bY�I� �δ�+{�j=R��b�t.ͥ�M=4w.���\���ˍY�ue��,x�I����.8��v3mDJ��qܬC4�YO.�Lq
�@Ja��s
��rKa�Lж'V�`��m�bػ۠�N��Q�׆I��Z� �
�I]ی#���a\�iV�(ll���I�B�V`�v���,&���K0
�(�5�չ�/���L��eጲ��4��VQ/b,��3.��B�Ç-]6�=�U԰��{k0"(`Li[&;����{�bI�2"�)Y3t鋩eĞ��t*1Q�0G��5r��Y�BęHk�t�`{�>#H�!�����H��w��n��3���J�K��U��lQ�6�@)Ģ�jV�Yc(��𫬻Ʋ�H�e�t��d6mH�h�cc)L{	Ǜ&Rx�����L��(��6b��{X)��YgF�lP�m-�n�`Ɏ�M�sU%�33�F�Ȱ�fL+5hLH|(4.�9��y[��bw�&I�P�-[MW�.�Q�j�M�Ii�p���d-n;�R���uS' �ܼ��W�I%e)�-������5a͢�ٴÔ��e��S�ܴ]fK�n�0�![`ƒ:��S�%��N�Fe[�;��j�rU��ڼ���,�Z��6f�u�mꨜ�	P˹/#�IV^[�H���O��2���Y������n���2)EE���Yjh�4��ږ���Gp�&��k*
۹yIk���L�yP)�Ƈ��H�X�4D^���Fݳ���CE��P뼥B'�e )�B�Ժt%�ǅ"�-�Q���Ѵ�ԫ��V[!V9�=2�[���pQL^��R�(K� �B����Щcw&��
j��"�ɰe��DR�RXL�b���5�S�یAZݗoуj���&6]�`f��:��vm-y�����o�-�VZ��ib�W�m���[8�<pm�C�ve����i�a�2P#�R���X��K�ޖE����
v�`����fb#鵕�%n]�xơ�lԺ�ji2aʻz�p�	�@�q�֫^e���ǋ^������cq� R^�m^ֶv���{�J^����j�hP�m4�(�́���Ǩe�xCSEM)���qR�ڽ*
u��ر���j�
�[@F�/F��y�� 7r�$�č��(�N��`���ͷ6БX�J�T&h���&^RqS�O&�0����]O�̷w"�SKE�L�N�FZ�����4�I�۱����Ia��l	�Z"�0�6��Ɓ��X~�u]���4��]�M&���qMu��ј�K�f�sc{4�]e�t1�cJ�C(��Bb�h_��(&4���rV1Ǥ�8]RYgGQ�ӎ��)	���\l�:�yI��
6��4h�J�M�@$���-R�] �e�pM�F���!`R������*S���*a8M`$�r�N�<��Sj��2�~QJ/Y��:Pr�^}���{'ٮ�6��a:p^����8ԳRѩ��Rf�&��2���5�=��{���m�Y�%�i`�YN��[ײ�DáX&Q�j�:�,�{���rP��6Ff��Y�����-5{��5���wpV�k"m�c#�A��Z(��=*�E� ��(Ӗ�i�M���E���k.�� ����Ǖ!6C;Q�⊪�iهE�-`���+ocY�W.�MC�^�5�T١�R���3>W�F��w
��20�W��W�n�%�M�d	�j��҂�̶��ͩ�-|�%+��r�bn�P|[p���i�#SƬ�;Ńo��78nl�mH%ὍՒ5�r�/�c��f�d���f}u��$�#%��cõ��ܫ�ղ1�F3q�W�CEۤ�⌙wOr^n��u��I@�N� ����L�0��n�PSш�4��ܭ��qK͢��L�koZ[U��H�S4j��Á�J�ܕ�m���!%�yH*µ^3%�����0��Rt�m5��h�l�lJ�fV�b�u�(	{W�z�r��J�����N�ܱ[0�5�Λ4,`A��]4E���J���i�yJbKl��j�.��ޓ{+�Ǜ�;u-�z!pe��l0�C���4�y�lBF!¨�|ݛ��	���T^�u�U��Jg#x�/j��cl;f��rօ�ա�� $�3���j&�ۻ�L=֖Moh��U�����HEHւ-=��R���jS��)M/F��А5�cfh�6�#�Vp!R�P��e�Y�A+I�T[V�O2�ud"�n���i�qe�� J�B�5ma��4uSv��&���4a�U��E�[P*)��ت�$I���5��C#�(��F�۔l<U����Nn�ں
�LT���1��J71�g0��dwh�j"Ř�lV���z��T�շ��*��	�e�P)������)��.��C6:���^�FF@ރh�Х�E�=;�j�"Ea�*�T����sUXI�A1�$��>��e�KY5���Hl6$t�jy4�jn��4��'[Oc���l[�yGZV�մk+��WI50��t�7Anˌ�^,sF��&�ïm�,:��,/\DK4�\��k4�+iL�)^&Q7P��j�Yhgف�Ԁ�m�;PՙXJ(�0%��i�F��c)�t��;�7XU�K���3Tf���Ro"��*�F��Tr��N�����@�Y[��C�ҵ\�jA/ �Uj��Ce����)�ָp&�d��f�$P6f��TZZK��E ��"�X#Z��v�X���dno)A��(伽�
�!�i�ԡ��(�*2F��ǥ�_J�腴�K������Գ��X��{!!�Rډ�ӡ�X۱���GC�����&AC��[[yJ���.m*��T�-n��,�5��,vS��ݙ��"��03�ڠ�d�č��cPJ���j�$V�DwE����T/f���=�Pn �0��ӄ9���y�/!׹��(�[����*�-�Ycvna�FsvU���/bi,Ӎ�F�76F��fi�Մ�+F������fe�HU췗	��m�Q�[*�Ѹ�Gv)T�NՐ&ն7j`���e���;GU'MB����j���
��И[z�a��y�lZ�\��v87v�L��WwӯA]'m��Yl����Q�8<��qճ�)K3.���B��'u��v;�X���vdm���+�J�|�jxbR�����'L���q��;j��\�`�p�\љ�3{�k;�)Ы��7�t�C׼��z�6{f�l�M��u�{��9R��r�8�{��妒���ȓ�]iÝ����Y�Kξ�]]i��ۙ��T������p��!��i���|ci��ƫ;;rS�O0����ʑ�zzhܗx�%`��3�Ĺ&�3�q��4�ۧ����D<o;�&�d�Rޮ����*���k9��,���@17*�r+:�t>�w��ѻ6Ҵ-Y�Ѿ�I+�
͕��72�O��WxGjqgP5�))Y�o�T�zS�"1��dW�Jt���׬M�KTR�fi ��0�Ib��O�N�B_N���
���4�;�6ۮg�8���}��Ya��}l����3���+*�4(�*����oy�\N�xv�T��/YVu�����tٜV赆F6�'5
7��u��Cʖ��>_�7~P���m
�{��L��܁=�\ݣ����vlp��9 �7L���)��p��x�$u��-�2jD@j�82�g`õ�h��f`P_k�N�ܘ��B�S��]d����m�®���vb�u{�5���C�R�9���4��i[ݠ�(���N����r�n}��h	3��Z@�v�a�D�WںRu���p�Y;2t����f�N��j��̜��qfD� ���;k�fp.������tL-�^J�ں�R���on�u��P��֭:pc��;��p��u��3��\�0���Wg�'��l����X����e��K��&�t<�Δ��x�����뎻#�d�t��`X^]`>b�;Rܝ�u�wCd�݌�`���I���,jV�5Y�ʊ�Gq]H:V`��G�,c��t�Q�b�X�]�_e�6!�?Ao$��GG�fc�8����U-`ݪ����j厏EYf�e-��}�1e�,0m���*Y��v�Ew�w�+�R���W��ޕnr�_;-�M삓ǵ��{���.Z�W�6JE��%�(Qj�X���[I�6�X�� ,����)%�yWS8�`AL���z���ʰ���#D����޼�#��:��g;����5�h/���u|�b�f#�kS{K�b;z�>�$�$�lK:�H�U���ӣ���m_]��m1\�KV��]��5L��	�W��CmV���'�q��mc_)��6�,��
Gm�~��&^Q!ޛ�ɥKލ��&�D`��|�^M �9(��8���8\oj��
<n��Ε2*(rx[�)��	I������Vsx���צ=�[�@70['��K��._uȑ7Nu���s���N̮��q�͑��ۅRVOp&�wn��D֞���%D��+rV��l<�S�.��&{�����c�8�(־���tXp�B�JE���,�V�ݬ��sk7�f��q�(	�p�{�ku��6��yȐ���-<�nV
ᝡ��0e@:��j���L�@8:�Zם������y����7��d`S9��R"�V��<�t̳;���!hu;�yqɩ�Z�"E	��.��{B�x�{2,v��� uG;��lA���!:VZ������ʾ[۴��C�2$>u�8w*�5ݡ������j��Uu��3�M�R2�*Y��׸b`V���Z��� ���R[-⥝Ñ���8s�ϝ^�ɰ�ڑ�U��^��Dd�fkآ�z���p	�q�����f�#AK4���(!�}٪�9���	�N�WX��n�+��_2�ٛ,J�A�zz��RR�D�nHz�i��j�q��tb��L"w*�#�̾ls�*�ϱ�}kk:N�		.$��.=��h�%8݀p^��tSv�ݥ�H�K��t�A�����������9D��}2�B�̾� DKS{�����4N
w@���-'07h<ޮ})Z��|�\��棼�}I[g;ywK�Z紦S�y��k��S/� �]��Z}C)sP�bI�f���V[�:�o�8@PQR��a��3���ͻD,B�ޭP���f��o��J�k9r����r���j��8�l������ѝSp���X�"�T�HwTxWl��t��&��{�"s����8�^«qrk��Z�q�ݠ·�7����E��m���I�su��C[��>َ��l�.<�L��̍��^�)f�#��L�� MG��Շ�]���#��c(�{���r��P���4n9mk�`-�1�2P�}�f�	ܒW5�B鼈�ڊ�k��P��<.�ն2(�!��s�_�.���9��w�X����f��ۘv�\�:*�޼�,=�&1r��B��v(�Gvv'�4���-��X%����q����V�ޝ�¨s�*�i=��r�s���#E(���ƪ�f�,�[�hql�Jť^I�5�+v��z;����ʲd��R�U�(��4*�0�tl�fm��m.�ǻt�rP�}{�d�뷎=�1��d#h���O��f���pC���8]����=�5�'�Y�ԣ��0֌��i��.��V�/Y�{{�z�4��ӈ��-Vʜ�#W!�^��O�VU���Q��.:OB�ܩZ�˞��!�U�wYc[;d�"����o��w�ϮҺw���f�l��lڱ� [;���#BX����1�^2M����D`�>���x:�R����v����c[���Ν2O��B��C�(�k�]�xU�4rW*�����E�����x!����O�l̑�ǐI�BG�v5� �fY���S�U��M�=��z&�%p��Up�h��K���ewt*�$fiy(A779���5v�u=u..�U��]W���~L�0�l7v�}1�&� E�މSS'.�T,f8s�)M����2����,3�.�A1u�t���p�Eo<�\����e�|�]vZK4御ՙ\o�KL!� �glfj��5�l0�&��/杝ܒ�ٌYLj.�*���pa�f��;����j]pdLk�Vb5��ɤ��rcq����xfL��}6qyr(c��Z�!cŶ�ZY��WI���6t湉�N�*�6���/�3��[� 0��.�%���#Wwemd�N�|�S�qb��L��xP���2ga���'Y��-'���,Nł-��E��P� �,�c�K��Y.j	��V&um�N���|��g*Ir�����x`��@R�y�5��0�P�v���떵3�/�Ow+z奘�"��=�>q1%�gq����-r��F,{�<�����gڤK.� kM�ضM�_=;��,с��9��2�M�w����c��F�hK�t��wB�vH�}����7�Y�AD�w��-��ΖK�/��H���I,�v�x(�w]����ɏ����c{�`B�G';'�s"��ھ����
���[��6n�I�1v��:VE;�H7�i>%��w�H����cŮ���m�tl%�k�R���n�g^ҧ ���;�RP^^��^3�v�>���ғbԳɭ�v���Wb�������z���eR%�Ӿ�YEuIf���▌�Pl�;r�u��nhG��P�֪KX���Տ��:٢��`�ۡ[��[=aOku�$��C����bc�in%W�u�,S����S�ٮ��v0MM��u���J&�iq#��3�q�)�P �x-����˩ѫ�7c��V��Ni��4�9ʔ�:���i���ŉVs����d)��_[�|��/�6���Y�YA(�����\���n�fMrf���2����ǯ^!ʏtɏ�S�j$l��ރ�w1\Z�d��͍���`9u�
�(�9L����÷�t ��g:�~WEn�T���I�ٔ���!�f��EG��9�j����ͭ����s�+5O�T¾������Ĩx���z�������*
�N� ��b�d�4�x 4kϮѼ����d��X���wXh��G��`�<ʷ�eSN*�Y}2�6���:�&e���Mn������j�r}Wt��.6x�;4�S]Q,��`���y\��@E����W��=
����F��{Q�g�h��(g��HcH��l:᷼�a��U힥��\/�#��oT{5=�f)}���GV2M��P��2�qE���F��k���t��s���Վ���9}6�"3��a=�V���h�x��7v��!�� I����(�$��<t Y�z���q`� �v� ލ�XR�o���)xS�]�e�'6n�]!��7�)�h�R�N���'Q�fgQ����h��o�ݗ�[��^k����ݕ�>Y8�qeގQ������0����gJ���ҕ
�]��ʺT���2�Pl=B��u�@2���=x���������"��3`	I⥚Ks;V�2�v_)�\3U�<Ί�]m�w 1Q�%��|�}�8Fr�0lǤ�{�js'F�brb��m�݃!��n�IL�N��WWTgg�G�.�s2�D��y�ꇪ����D*�X����BN���x�e*�Yz�{>��������r��%��Gb�l�
���	v���#ѠN)�X�N�H�&Mf;L��n�:^T�Ut�-D�3y=L�xh>}qf2����kt��uKq������h��8�S4*�f���`�{�jv��۽91|���,ءZ�}�����2U�R���	yi9כ�P��MZի��3i��kL���I��s4wn�D٪:W�u#�M�E�8m��`��0`�p�/���.��̻�),m�T�N{]+L�z�)1u�%mm�x�QB��;��_
⹜0s[�D���Z� �1v�m"��{�ݝ���f�ol��RNwgnD�1�(�-��,zx���]`�����N����,�̃h�a�7Xy�M//]a��.��u�di�5
���/`��������Z�"��.�l���+�|iG�+�R�+�@��AlZ�=��|��#A=Y�y;/���!ې�ٗ�և-t��Bȍ�u/�_(��H��O�"�*\��`����8^ʗ�����`��\s��[��@��2�<�Ͼxq0a�ױ��Mm����K;����S=[6�ޖ�;�u��N����S�u3sO ��Q=�����8�n��mq`�C��pm���ܼr�X�}RR�9�jwC�Y�b��6��(v�Ѫ9���}m��u� �DG�eؑ,t��T�4�'Vp�2خ|��X�*��::<�G�U�ђu���2�R�orC������j��璯�_u%s����vc
mF���#6������VЫ�-T.R�Mv���^	��&v$&T���iܘ�î%�r�N&��j3Q��{VhoF�5���k���ή0�^['���&�b���)���/fa�Q��jh�ۻ��7�}Y$�3��Y��׵��p�g ��S�1v�k�cx�n����[�o����m��nv%b�����:��@�'�u]��hF�Z�<�V�[у2Eل���ӄ55����f�Ŏ�)�.��|��8�L���8��pa�Yw�&vt} �QsB��N�9[/C������\;&(B�ƺʱo�ٍ��:�d����3Lp��X�
�G�`һ:z4��].��t�ݽt�o>yJ���~}��殬f_f�h����y@�����c���m�T�ͣJ���ƅL��)	3uV��j\���uH�@�CV>��B����7]�A�a^E#"(e�F�����$�:+��Ch�:���t�B���X&n��/�b�ǁ��	��+��-ѹ���k�-��t�J���� �n�X�!���\�������n�gv*�-Н(��z��e59󽷂���켽�(R�>�����N�wZ��@R��u��m(S�C�L���tU�VvYw3ܕ���q�8��]��*�PX2���t�۹Ư	[�/�\|��� _H(PJ���ց��-���U�Xfq2V��V�̳M��@�ٸ�';�]��L���0r�M��ES�b�5�״��Xd�
�o+8�Z�����%��>S�2�u��cl��:�.�t�6:�v���mԬ�NN�I�ؚ�s㎇k���Bf�=��>���ʋv��O�j0H�0�ȑO'`��3 �7�S+GQb�ڠPq��!���]G��3ˆ��� A�6���re�vޭ�%�"Lf܍B��<�S�]�o�5��&)���})�Rԝ�4:be�|�X�<iլ�B���Yh�ij��yv2�k�Q��jw�S��8s�aё��uN���˾˧;���n��]5bPל���[�*��pm���ɕ6�&[M�ZC]����+�B�Գ�������̸���)wWL�]�.����6ڑ��tON�T��S��uo>;{�b d>�a�O�8�ZZk����1�#B�[� x��0z����-\jR�v�V�:&b�0d+qi�U�u�&E��C劋�SGڷa3�IC�V��������ڣn�oZR�����o������� �]��s���O ��M
̤cg
�b;t6��Y��,�؅�ڦ�w�˗�����;N=���U꾶��(Nf��4�&&�ޮdu���Z�$�܎4�3�*��0�tg�������\x������g�����Z��*�k���zn�2C�o8	4i�N��Y�����6���G����p扼��W�>ڳ���x��m=�#Nq��n���N��V� .��yo��vn�S�[ó���݅N��e&�V��8�{Vq<���/gw���w�>������>}��G��!km�t'v��m]�of�"ĊUe�QV��ۆ%m,��j�ʛ��"����Cw��:�4�9X�w�Nu.6.W�HJ.�l��2v�m�s�+6	[@�Ӏݮk&U�j)���Q��x!��k~������p���1NZ�q���6�5vQ�`ѧq�o_4;	�56�9zgX�d���"�+��v�����;�9B�U�h�b�%'6�%};# ��V����&�[�8��<,��{�f���}��أ����t�7�&������Ĥ.��.2���&-VI5hT:ĭ�b��p!��M
�x����;'L�]g>;Yb*qoZ��F��5�۶&���n���f��H;*rpT-��	�Q�6�W*�(=��x�Q$-��R-��y�������:��/.�<hm����f�R��/����}oz-�+jꔟU�G�l�ϗN��N#o]ݗ����r�ޗ2V��*i���̛�ڡ}�T��V�YŰ�:!���U4���m]�n�M��7��r�ˏ�Y�6�ͭH΋6P��;i����yR�M��IGD���a��.�њ/�[F�Sѻ��=t��2kF����4��qޚ��.g*�dg�oE}ui�77T����Wv����С[:iӏ[�]o�RV��G˳TquM��W>t�a��aܔ�U�5�բ�r�_�K��ݑ�En��Y��8��[p���c[Zu.�N��%��T+��T�3�M��GWu1}@��ɧ�tлݍ�:�<�M`��S\�[����쌺8�����g3P&�(���e�;K�>qc��j J�Y�7{�uV!�����qG�v�X�R���.��W.!��y�MǦ�YaT%*��dh��7�aX�u���{�^s*��f�9:7h�?^���uk
�p�֚ޥt���.fRD\�5�q;����k��Z�s�X�L�#u��-W(*qou�f�pZ�Tk�%9�P�q�"�Tی�'b�uY���kA��Sf�n%}u���Ĕ݁�z��o
lD���hq��KǶEoRҜ�V���A7J@^
V����&���P���E�7:⺰�y�wƞ:J�XY8P���k:�m�$bw1��^t��8Ӿ��(��/4Ax�ˊ�6Q�m��GX{]������Ѽ�wL��n��c$�܎J��G���=T;b>4%�Q#���iM|4��dΡF���(ۙ���Я��dXЍG�#��Rtr����h�uP�o�RHl���Ȧb�w��L�ٵ��W{a|z�V:�4�txG�T��Zu�Л\à��
^u�΂�7��!}zĹܣ�g�y���ŷg���u��m	Ţ]�}l�k)��W�L{)mc�g^i\5N�w-�iݒc�9��JLc�]>�Iz BT�|�Jp�Lr�j�$��p�μ�;)c�׻�/���{R���֬�f��'���.+���(�X�m��[��p\B�L	mpT͜V�f��wm�ʀ��S��[ ����ӚU;�%��w���o4�n+��,7�8p�:63xWe�.2�۽"]�P&��Ʉv�"��ڏ��3�GO�Vq�]����v<N��1�J�R�=Ƿ4�%0�I
FGZ��:��/��<d�n5hb����m��M�!;�����	f��6�m���q.����h��x���6+��w��b���'r�����JF�m���N���Rv�	�Q#��
��GsQ/R�dţQ�����1��c�VX�����5�C�6�؉(��QQ��7��-����ԏ
n�`��%�4�q�ռb,���ߦm�ʂ�Ky����dhBN`.����c.���y`��DZ	�������Yf��F)�{`�q+��-�AS#.Du,/�m��*�30R.�s��|��X��h����[
�;��i��YlI�:�H�CV��vGn<�=ԝn�C���h����^Ӥi�J��ѐ�R����J���BƝ��g*>�B���Qq��r�C7k�����л���Z�m���򇩐��#(�j�csj���
� ���Ы!lv�w��Iu}R�6%�o8� }2��e+��6i�	f�-c�[H��Q7��;�1d��oV�%z�A�AV������9�J�Y��A�޼be�c�0�<+�ڠ�P��[��0]����� b�n�"�y�7����m5��(jbBU�2�{lAx��`�Ս�z0h�S�r����y.[���Z��+�4��ĭ�F0�=�������h�
��.����ʇ#4CL��m���u��I�9���aQR��G�t����1����e�V����\?O��a�|�fdsv�Fjc!��"�H��x�7��ӣ�J�l�@�)+B�P��
�������6��8�ZUu���3RX-�Wr�x��{��!+�k�-<hiy|t�[J����bT�K��:��MwdLХt��ف�t���@-.MH�R�%p���d���6���Zgy�)�Ca�;Յ.p
m椋ųU��i.����2������������W9�o]�5�8�\v� 3�XAk�G�����v�]��%F�����ү�2��w�CӬ\ںd��P��!ʜy�k�-�eEj]�E��鈬�)j&�u_�Y�:�U�00���zj�w���ݬT�lIggo,��S��>aw�i�ճ�
<6��Kv���Q<i�ww�"�Wpt��J��ux��W�����#�3�u�<�wyS���1�h�̩�4�-��6z��+�G�4��ۍ^L6`(�uc�5}�E�o;�beA�Y�`c�侽���Է����AhV��/�me��]w4��Ƕ�[:jT�[���W e���x�-�t쾅<8B궟�cF��)�񣣀b�j�
7�����i�ٸØ���f��j{N�ّ���`s���
X��O]�t�p��{T����:i�ԎV�Y۷oW*s0�4��of���[\��!�"�Z�7���f>U�z�F�ޥ-��1�e�.Iy�2`�Ym�0%�����ˬ���*ƈ���6Q��b0Ư�).������}���V7P�Z�i�M�ӴC��hL��Vս�3"h�Нb����nl�y.���[�R�Cۉ���
��W�U��b��tbӣ+I����d�SI7���jZ���Ⱥ�ұ�}��'!n�vXK��e�>�.r��P쒦Ճ�XW>�m�ʙ�� �V���l�0!�B}��n^����LY�%��
f�T7��𾉚��s9Q�ɀ�/5�m�����ToT�A�s�Z��v=z�#��_h ��nN��ÝY�4Zf�p��릳��;���M6�h�<�or�A��%f�*�.���)s;=��V�]��\{qܥ���/"W�	�%�9R%�Y��h���]�f��_9��,,8x1Gf����QϴV҇ggHU�8St���V'����S�=������Q�n�|�}��Z3����w[x�-�F[y��:�-#�� ��E#��=wl��ڵ52Xވq���o:ٜ�7:kg
��F�󳘾+���7݉���ڼ��7Y�ls�x�ɇ��*	���C�-Ml���F%�c��@�R2�fV�]����u
�H|^�խ��<������j�:�Ow]f�ô�����w����[V2��c�S���y�^}׽PH������%upBX#-R[@ ���iq����E(չ�rƾ�l���{76jl���U�l�V���ς[T�Z&�M�Ƨ͙�3���y�wu��s�͠N%�X�����{W¸PS���h{3���XpW^�څ�д�r������Wq����ǂ�E�9u^�۵��/�q�Ѵqۮ6��H�gU���8͡"ۛ&G�|���>O+Lt.��J90��ߢ̻�i1��0�T�I��;Q+Wk;����](ti��4Z��Kc�ʄ=��2Uհ�{9�쓮�A���t?-8)�@	�F��d\c�ϤnO�5{�x��^BFc*i] v5�b�}�o5�
}� �0�V]�u���[X�G�!Ԛ\$S �X3��]�z� �q%A��}3P�����)�u��ӳL��2�H<�3j��f���䡑�Tٛ7痖�0�C9	��h&��%�wثo�p�˧)xݥ�u��);�S5*:(�ۛY�K9O�ɄWI� ��Q[���K�՘-��o@��\bb��rN(c�WqA+�7Sw!d��ȝ'F�ުYoP�Tn��_��X�R�x��ON8v� �6.�Gs;��wl�;�]\�*[l�Ԕv����'O;�]I�B�-܆52�}�嘧>[2At���X��o*�
�o#��)�i�݅�;7CoV��$��zh����\��OP�P��������=e5�r��r�pi�\(`�wR�ջPu�k�鱷��>}��\6��[v>��]��Bz�;��\�X��Vfީ}��ʞ�tr��ڜ�R��]�<{���꣆�� �0o��@�2eKjw4�=e>}|�@��nW�����i��t,��0)��fXԞlH�Ao�������6T�� 
Ğ��Ϳ��}ɭ��r�l���Iep!a�}��I���C��ji!ᡡ��9 �����`t�G�(�&�&#W�����I�3
]�	 �n�*�%˰�빗�#⸬�P�"����HvSWww-1,�-���F��k��郄)�r�]u�)�c��r�1|�Ō��f���ٺO�{�D�c��)�'$�u����[��*ގu����L�BhLɶU�[�䩭i�u��.�&�����:��Nݡ��s�'u:�:#_L�wk��܅ЫtWFe}i����grC:�l�m��/�g�c�ӵ}`1@E}��K�����n������*u]e�c%���}����zK!��� �_We�\��1;8� ���$�W0���s�ݾ��xB�퇖��w&�puC��_�0u����Ϡ��:$�!<nM�P5\h�����;�C\螗v%���/""�rt'����AGgo���� � ]@U�&�Hq�.�<�J�}֬mB�b���M��m�x�7�R�IO��K����Q{̲��(*�ӭs���ұ8sM[�4N�U�}/�B��1� �|� 0ݥ��7��-3�dIR8��t���A�.��k������'m��a�R�N�B;����+���a��X�un�n�8��z����e�kmgF�J��c��}����Y&3{@�9.�G�V�xt`7�*��u�d�:�uY�J�1Ό��P�hx�v��3U��7�;���s�
{q�7�]e�mc{\f���%l�u��5��@�-�U�L�&�96E����Դ��b7�kxw�Q�M���:],���,�V]ҮG�t{�=�C�l�}ټ��Y��ϊhPn�
�a܍VX�bdӽ"�¥K�n���V�t�k:]=�aެ::О�+C����@�]�4���y�L�5]F�}�IEғZ����2�m�� �`�4]s�Ja��������s��]���3��8��̝`%38o\�׭v�3�*�,�p�/v��u3�9��N�2�oNv�{�*�h���SK����^��,��jGI"V��򥾦���`۬ݰr�z�5�μ��J�9)��>�}}-����["a��F��n�{j�˹���7�o%�}����uvc�Bf�i#�i��X@�8�X�	;�g(�(ū6���z���:�\���.X$��&����V�U&���gPH�	�*P뺽Ȅ��F,���1s� D�v9�A���f��d���v��d��]�	uꓸ��Ք���v���9���4��e��/TO���Ifv�Ҭ۷y��6�����˚��S�;��(^3S3����A�:���qkQ�#z���k��n�y2RV��Ϙ��d\r'���E ��ۘ!�<����ޫi_p_�cvb�G͘��M��X�,�L�/>o:�Yf��["�p�̩oe�R�;+M��h$�s��q�F�%]�ʕa`���&/3)ǣK��;�k�ac�Ej �R:���O���h��-�z��*th��KF7�\�U�*��|��E��C�����J�M�G���qA�
2SF��`�bW��Zj�O+�b��9r�[�:"���Ȭ��V���ODh�'>�����e���Z���Q�tq�k�J�}���9(e�q%-�;�s)[���&k5g�,"$��;-`�SU+4;S���z��	�Dr��\-�`��^j�1
�YW�Ә�i�J��{Q�Yi��&v��\t�EJG�F6�3�we�	2�F�����rg�ְ���뚙�Sv'�9�̱p�ɗ���Zqw�ז�:f�[�y�	n_-0u�ʎ٩΀oUl��9�2��X�#p[��gus�ۅ�v��R����P��Of�)��V�S��3:�3F)��V�U:���/�CYRiW��e�kh�#������P%/�Q3=�Wy�v��Ǡh_���,3��N�ے�3j�u�v&�[䨫4ͽУX�fqZ�.�v��Gka<:r�6��px��ټ��9҆����;U����[��Z]${�;4A�=.؎�$n�y4R����7���ַ'\�������\��-�PΛ��+JU��J�2����ňȔ;0Q��	 �7c3Me��jj±�V�9/pm�)�r�M���@�����M�gF�����ҀsW���zC5��Ÿ����o�����=��*?v���ά<;0��Rqe��Od{�(����p�*�f��n�U#'DE��Ȁ4�Hњe�'-����ܱ�w��|���/k��Yf��U]�:΀aӱI�y�PV��4��v���2���T��������u����jIW�ƫ+Q�s�c�x�y�S�FkO���\uA�<�v���x7���}�LC�\���V���vf�$3wj}y��%1.<po���ٚe�VdN�j�6�P����0�j�����ZB�r~O%�3��Qo �R����.֬{��k:��/7�ƃ=ٳMC�WU�B��t�.;Kmq�cVJX2�!�W��2�ä7E�0��^�L�4.��;;�qӉ��n���UX�8�:+��ظ����(\Ox��CM�R�N�X&�-L�S�3n�� �z:oun(%b�İ𵖗4@T�C�}0-����[�Že�A՝�>ת4�s�`�����;�T��o�vS���_s����х�Wh��qwED�����9Uź�g:S]����Ե���z�����u�K�Z�-�8�c�d
B��u��
�y���&�g%,a��w�3���p:.*໐��OLm<45c&Qt0�9��:���v�X=c���F��5@7Q�M�}�,�6��*ت>Z�h�Y�k�c���NS;K��nc���pݼ\h��&'ˢxD�-s�'vc�v����\��ՈaR��sBq4l��4���!d�"<�*�eu`�C�p�Fk�;{�N��V�yt�u��<�S���;�w(j�qd���w���Xi>�kVpx��Ժ��@��֫��,����ן{��Z�==�����30�)���
2��"0�23q��	�� �H�3+3
j32B� �k&����ȥ#,�&"jb*���p���£0��p��,����� �#&	�2̙���1�����3"f�*h�,�"�Ɉ�*b(�"�fb,�2"�&���*)"�����̌�b
�2J)�(���23%Ȉ�Ȫ���0��"�"�3 ��#12*�2)��H���*��"���2��"&"rƈjg0hƊ�(����s2���r�`�
�j�
*���+����������(�&� ����(2�j�,H�)�����,��&�$�
�0ʢ�2rh�̲jH���r*��,���0ƩJ�Ȃ��*`��0��*��*��"2̲��&��s2�+#(�H�+2L��b�!��*���"�(�si�f3
ƚ���*f�* �312��1�2"u��|��uI|m:,�>���bv���Z�>���q̔���N9��t���b�+TkZ���N�Z��;ݝ�{6S�s�c�v��U��ӆ�vW�tTX�T��N�avZ7�=�4����W;���wV�6�(��+��M�F��1 �V �/}��!zS1a`A[͙�����5[�ꭏц��q�g�Tǫ�M'	�~�*I�E������ۚ�uC���v·�RV���)�8!�GG��q����`��=��F�f2�XLb�����U�C5�s�ʅO2E��zm���X��k���r�g��������+�o������A��CK�F�t�B�j��)�^�dR���� uu!zV��+q�3�ʾw�|�A=��D�S
 B�_Q��9$u@��\��� [Sq�t23T.ޚZ�34�����',L>5ƙb�Uc9
v�t`���:���W蚭[0{�s8���w��͂k�\qNeA��,��dF�R�Md��]Ez�F�1WF��`�y�}���'��:�`��9��i����裡��`�����*F�gL�9P��L6+.eFMn����ϭ�������;`����)�n�j�c�(�R�|�%v9j�^k)l����]yy��{R���t~D!i����w�:�\i�,���>�ҝ72��K�3:m!`��{��χ-�.��u/3�\�U�]ڕ"���#hz�ua��Z��qp��N�	[��O��
*�X'piJsq�xWjK��,��;�֙��b�J����b�TM��g|��\�9�~�Dɉ%L�kR�OngS������^�Yz'"9���s�eM�0m@q�,;'*'����I���a9힁3���̫��/ʥ��S,v9�3��w�]w��bo��nx���Qb��,@��'��Ó�c*U/�o��,�8�:���f�Kkh���u�~��AVSVj���RMS�y�Se�	�+=V�7�F�<�:����c٧����JXa�vw��I�"2^��(%C�FkTΌ�uX�U��Ԉ�ȁ��!7a�4�tr����a=����ozEV�����կ&�p�]W~�!�2�^$r�ƍu,�*_>=�_�:���a�k��U�8T�����۷�ī��
��(�����Zd)����Uc�R���Mv]I��ՉZQ��&�q҃�qZ�p�{��N��� B�68	e������"��yؚ�>jY^�D9X$#�gWy��3^׈�<�o�6��e%7i�֎rs_9 ռ�n=�nȁ�b���"&Pƒl��AsU�$�Wu�s|77��[w��z�Uⳣ��iv<�Xk�Uۼw#h�Epdv-�f81��,�T�������C�����I�-�������[h_��"��f�e��_S�g�f��H��"&�-#�o��iJ��-m�r�ӓ\t8�6��F5ֻ���f8 ��V�6�kY�r&YbAx9MSTz^�i�՜�5��B$P�+�A�V5vֳ"�Γ�������`���|�z7;z��6�5��V4�ͣHhȽ�	H׬�Ŏ�����&�����O��=���dV�m{ob�s�:!v��5�]鍀�N	T�xSMWC��9�7����4��ة�Ԛ@)z� U{z �ʅ��P�{�a{��Kʗ\���لmc��[t�#���v�~�= V\#��%�}��7�A�Q�*d�Gpq;��d)������ɧ�k��M��B'�;Q��V��/%�:�YA�yC���Z=�hl�4po ����Ss�7rp�}�z�|r��*��6�'x�]�C(*�6Lg��qKA����i�^X��`WD�R�સ��R�r�@ke��)�+�k5ٝ×��o�3`�=Kk��uh���Z������J����^zx������U�v��Տ�ݩ pc�b�����������i�x�}]Ո��yu��=��t�`�4tg�[���J��o .�'�4�r�(���3�?x��oK����qk�E�Dgps�Dˣ���Uol��w
D1톞p��i
�p�J_gET��e4�o�+�ͬ��ݝn�G`I����N��e��V|�m|+�VPb���eg^+Y}ן;={^�vg��.�+h�Y[�N���#�p�2�|Ѩo����q�<
�u|����K�K�R��d�ި��m>q���n˳c�u�-�ё�,E<ډ����t�T=`�k��C��x�J�,fi�݆ �q��u�]ci��F38�iM=@���4-���m�ÔjBFn-i�)Ί�hd��U���+�R�Z��B������-���Z�����Ƶ�g���Gy�.� �;o��rej֭�j�7�6����.p;U[N;T�rr����D��V�}���Qj`�+��A��L�K�&v�0X�b���6�s�*���>�N1< ��)�I�*=μ�Ȗ{D��ڸ쉞{1+y����ݏ4Z�a�� �H���P���(��'GH���#�L�����v�F�h�t܈��p��ެ�\`ǌu��75�cʼ�F���غ
�캲� we(�ZDۭn����4j�!�/��&�v�Zb��24�B�gH�o�=+o�Z�y����wvos��ၭ��4��_�[���s������wrK��oՓ�p��u���ǈ9a��:Բ��F��Y~z0�l@>��gG�_�^���P��k��,�>VJ��ؖ����k!c���`�]�d�³X��=]��8�qr��g��X�}3//��Џ�w�=E�;{H/�
g��3�o����z{��{&��4sGqm��q��en}�[�:�-	Z�KE'\�<1�C�18��W-��a�������^��Ġ����ۼۮ��wd0\9�*bx����M�D̖�\v��%�u@�u��,6TK��sá7M�lH5���g,�Bj���t�m����u��>���G����%%17?77��x�
��p�7�T�<��*3�Mӄ�"�.�A_��Ө��%�ڙ�S$v8P�i\nF�'1�G4\! �sتeCd������@l�S�u*O2E��zr"�l1l�����g��mnM�$o��U���;���[9R���O���f�I���ʃƋj�Gt�=��{���w�z�=a>ǷY?n4q]t�s	�X��48�ѝ������pt�����^ )����֑Θ���92ټ������ӵ0%�vz��.�u��7{��K�+��R\V����-��	-���������z0�V�:��We��[\������"�ue���c�nV}W�T9��/��#�����K�}2 ��']Vvq�[������E���>�U��&9�L�n�����#�XtGTu­[�!˓�l�Sg_F�f<� ���b�{i��4<'N�*Ƿ��v�F2T͇Gz��1��c]t��C�ض��P�Ჸй�x#�<r��G�V�e[�@���P���oG{b�P�x�����Û4M�M�t
b�k�u�\��&'g��7�W9��(!Õ�J�]=Z�C�v�͔�ۃ%)�����(c>�V�d�X�]V8�MK�^�ڛX}ǹ�)7����S�5��|ꗤǵ9�u�gY�2� ��eF�tM��@*b�.����]��tj��#�b����n���Bey�A���Y�s���S���bHU�G_;�7�ⶹmϖ��u<��p@E���3���n#����e��n�\c�\tJ��+�5\6�wu^��.4p������C3xˊ�VX� GY`t_+�Q������J�O2�N=C(�k�M��SO��sG��e����Ѽ���|��9�W+iM���K�*�7
�]=��s�]6mG����˴�[i�ƕ��B��ݝHN=ˣsQ5݉��9�#�#;>;��5�1C0���E�Ժ�t�
�w���uh`r(��OqWQ=
��q��M>U;�R:3�걙�}R"l� W�*Bn4���tr�����"%�J���=gz���Q�7;jt��4�T(�To;��d۩���*A��*����l�ܳ:3:���]g[�a3~/���CBx�pp!30�i�Pz8�.9Fp�r.�	����4��R����w`MP~��\d�Zn�t/��n!�%�C� U� �ꁐ6ut�V��&6��N����Z`ֻ�:�*	����t��O�t Y���@n�e�Sv&h_BĜMv�l7��"+H~=�FT}7� j؆���6��;C����"�XϡЌ��W?V��M�}ʦ�\�/\�:�\��p�3�}���ֳ"���=q ��L9�.7�{;�g=��Uf�u��esMz�!��cCQ�Yt��-���d�F�d��pT
.�l�o{���(�:�����X�Bo<�S��{��t��|p,GML+7l���w7.�����d�rMGR N�ȍs��u��s���Ύ�B��u��d��٪ym#X���'/w)�j6�,\�Ľ/�ہ��:�br�e��������=h�wwd�3���^�Ǯ�<�9ę4�ٔ��ܛKr�4����O�`�2���H$
�F]�M�%W+�Ͱ��7>��|�N����}���>ƨ��*6Yƫ(��䮮�E�?m]C�F�iP��bj �@����u�ɬyS'�� ҂��c�H�g�)�*xa;���AXa@�q�FQ��N�_�g4��c$��<��yǫF$�rR'q��]:�|s��	W,	�Hڈx���=���y��`�ռ��V6���s�cy�ʺHF�����s"oM)O�N6��>��ֻ�����I+m�\���}�ũf��9cuN�A�o�:\���q���]u��)�G(��j��N��ι��'v��{ܧ+wm/��MD'<�l���5!��T��;��r(��^%g�O\W�.Ύ�.3UX�r����4j�A���Ƅ�*�C�^UH��g8���ӹ�Vt綂,��%�8��/�s��۝�,ECͨ����.�ĳp�H��j{�,s��r� �4�����E#�saԮ��~<��#�%C�B&����(8�:�C�C��v��gl�{�`r�9D*���$Z[��zk��c֯�80�z=`7�4�!rmmD2�2�'y�]���U�ï7�oA���^N(u$��}����U�suش-���b�vB�yx�H���2�:Npu�C;�p)ewC�-�l��w86.��J3���:YI��_Q�d��.����tj�چ|i��Pܥ['�R��"+l>8��B�ɟV�}h[�#������fǰ��A��s�!9����gdwh8�JG���'U_ܭ�4t�{��cx_�S�g�G
	.�V��ܝ��c�C���ۙ��C�UxK g1,hrN\��j:j����3Cl6�8N-W�l��4�7�㯏f��gۧ���7R6����*��H�����D�;��^���A�Y'�z����/%�5�j��z�z�F<A�`<m�,���vGyf���>�] ��ʆfףL��!���d#Ni�S������\DŌ��#�B������*{��57�}��� �"�'g��C�м�,�Q����Dd�,\B��wi�su�3^��kp�Q��KjGiz�`�c{��c�f�\�ɸr}@���-��*y�C�n��"}8r���T���J�7���:�Ùa��SA��6�6놨�]ƙ��(h�s<'}J��y�J�ާ��*�*r�h,�V`�S{9�
�U�ͩa�~�u�~��7M�9F�}S�T�b�H4�����Y�+�O6�>�@n����Ⱥ�b�H�J�:���|�%��C����A�hL��f֙[��W؇s�۵��uj��p�+[��e�/v�9;�VR;�%]N�iZ�S�;�.����Zƫ9�ϵvh������)���-�{C۱�����A~vد��P�6}|�.�����-�/g�a�p�{'	Ӷ�a�R3��n.��̒\Yt������K��S>J�pC�����������}�>W�h�M&o{����*������0�.���d�=���T͏�k��Y��=Èb�����NC}��󵴤WY�Ҵ(Aٞ	���<�+��<Cj�Gl�*��}q�cϫ;* �*�<O�����Bc���z���T����: 77��:�Z늸��<B�F5�M_l/�ӎ�h�SLϸ_W/����wx莖�j\�"K%�㪃�q&G���&33XS�u7��b�b�K�f�)}�����������M��o10�"�*VEA��\Vޥw����5�A@~�j�,E�x'�,��C^��2*#��'�����e��s����Ǩ��mn��+4`58��U�
c�=Xl5k���+��Uo��\s� �@��96�-@�X�4]8�� ���Gsq7δ̡Z`�PXu��+���:Z��U���lvqY��wZ�s0
:���6��ůws���H��W6�:��ƶ�ietbaGה���cb���NA���t�1��z����tѡ|L�|�DZ�|Apn 1\EP���ٮ���^�Ͼ	���&l�A�m�y��3���_Vñ���m��ΘnK�n�Q���}Xj�.%\J��`o���:�}�Vc�t�J�q���*���r/��ذ붖�Ti�1�5��ޝ�௾�5
�fQ��]T.5���*�ӛ�U˽���i3�Kn��o�PU���)�/Q��5���9lԒ��N�e�ҸX'���jy�H�:��L.T�<��.��fwNWn.n��8�?e�W@s#Ejk�:6Î��c�7���,@��ebɃ%ֱ�fꑷ}���J2�!	Ekok�Y��;����ٰ�H�>Nfr͘�Y�z� �I��q�����J��=������,Y���ܩ��ժf��|�@N㺜�������EP�:IY̓�t�wSH���L���Ye��$�c��(�r-�Vvl��;[Q�T���/�����˾ST��P����s�f�cb��&�(�X�7pc:8�
�7��Ѷ*��ك{!<��(wZ���u{��2�����%/�1ʰ��Am�4jJm��7�)R����
�]�qf&z�X0�U��	io+�]�[�J��y���1�6��}&�;ك���ݨF`�q4y��u>�K:��7Y�P�<+.3�'���N:�ʑ�8-v9�$gݲwmr���ז��b�w[[�+��
6]<6��=��7�&��;K4y�y�`x{��͌┴v��v��r����N�D�n�6 �r�e���@�]E�(��7�ḓ��L;�V�<��]u�<ޓ,NQ��.�ImtOr����U�.��&��fRy��V����*�/�t�s{EK��L����YYO�OM*�:^_��k�>��$6e�#დ��������͊�C8R�x��Ļ�ܭ;h��QF��"�P��T�­b�aD�0uլ���nq<4]�Bs�W�ȼ)��Q<M_d�u_KN(I|C��4��Z�!ã9uӸ���b�Q[�`vR��u �mt�y�<�]��܏5�������m�ߝH8�;��Sub�V����Vw�=����ZS�帄�N�M��m]w-�[m��]�m8�U��W;�`v���E�[ڸ������K�T������} ��B�J;Ӥ�;u�Q^�]
�ˈV�TX%]���Cye����Ef�ָT;X��s���a��Y�;k�m0�샃�,z���ϙĒGT��x�Vk���y�����t/�I��Ӓ���i�PAc�M��x!�[�6�m�Ʒ���:�n�ش$h*)����lN��+��{���5��[�x��A6����\0K���N��Fvݢ�ӝ�^b-QE]ٙ��َEA1Se�SMY������%RQU5��Dfe%KD51$�3Fa�4�XEED��cM5QALD�T�Q5DS1LQfeUfEUT�Y�e�A�fefaD�AM0U%T���UEMIL�DEELFF4EL4RSD5EQNfQUM4�I5�嘹0��A3E2Q5EQf3MTUSQUSQf8�SEUe�Qe�D1!�5DVYTUSEQ9�4�-dS��E���AfeEPQREQT�a�LX�L��Y�eQ0E�QQ5UDQD�4���SPQQA�dDIEa4FY1UYDQAT�AQCQ3EE6f5��f!�Y�fYY�D�Qa�D�9UEfy���~�����M�G���5Y�Wf��k�Wn�'���a�I�:<v�ݏu�R���5�4�m�+I��+����:��*��4��^�o/D�)o�\�"�1�X%#�M��4�ܦV닗�&��#=���,k,�7��X�Zu�g!:�49��7̪B����)9ta�Ų�;�wp�8��MF`-0uΣ��������X��0����Gc%�ѯ$!l9~�s���U�����S�
�V�	��
�򥺻�D��ܞe/b�\��;V3�̩�8���*j�	��d�3U#�h|��!7�)a����&����<�\4�����.��2)˒j��IƢ��^w�ʨ�_Z�nwtѢ).��{10"��x��p�WK`��A�t��p!S���gU��q�\r(��Yv7"�R�6ل���]{�9j�[0��:�֮���z'Iod�!
j7Y�yNƋ�[���7��U�ˊ [Sxl:�j�\�"��f�^�U�;�q� i���tޙ�S�z���q��ט����[�����[�*�4�UTW�����������ށ�˿��#��M�d6w�GcTfM2�����C�G����H���sl�3�������x�j@4�j%I�� �����悪X��r��Q[���+����L��6�1qK)<���Sv#�j{Ӕd졥Z��'I�;+@��.rZ������s��inoX�qv�K���F��� ��Xn��.�����fEs�'�1
=�ۜ����[��F�j�v�v'xh�<�̤P��}��H�Ya�v���̒c��52�f�%`�ǽ[/R#�	�8����C.�:�R�Ж�t���pJX�)����]���>����vW*�a7�Rk�@sJ� ϵ;�yP�V)���^�e,+�s��c[ԯ]��I<x���R�W�"7#���֗ ��R��L�1��7�A����0C�ݍ5a��0�=;��󫠬�~�������@��9�Y��q�FQ��N�XL���\�q�w���}
rc$��R'.��WJ�_f�XX&4:���1}2��D3fiu��|/�fH��9�Q<�_�ގ){����7!����h�\���m00�@�1��y��4L�y��nmGE9�݊��*-���뺦,$cp�\��\Vu�+�}R�{��7�dk��!Kr 6�\9A+�Uc���
e��=s������A��\�N���J�=��Jӯ�nQ��J����W��[q�k��j�e�5�WCW�z��gm�;9'ڑR�g�	�o6�2��G��չ-,�l��T�:*�g�Wv:�yCm1�t�c�X��1R�vPܜ�>���d˫�뉖!��Ĥ3k�soO+�Ѭvq����9�Y	G��5�X��-���C}H8ju	�Uè`��U 0�����a����e�u�� ���D�qϝ��=�7�I:7��mD��\zI�Y�ue�v���n��@�pf8	�+���,0(���#�ci��F3 ��m����K������%�瞜]Xa��EJ7��DvP5� 3��**,vJT��m�uV��֚ڧ䆣��ut���]��e�9(�jKj�E�T7�t=7P|���
&(X��1��r�֌�͂7H���(p�$ Ӫ�.�Rt�{��(:�Jr�y�Z��}�`��y��[y�f�}6�fO�%�xJ M^�?	Cț!��y=M��A&1-q(/\����/���Za����Q�N?9�i�Tn�I�iP���B������D��_���O1�"���"�#\"'���u���K�4z:bpƸ*N�L�yK6���e�O��Jƺ1,Q~�7���حׅ�P��ݔL�c��
5��.݉��⃩�SyQt�Wz������k�).ZsX�h���a�4� ���%�MK��R���g0\��T����`�����͡P�w���^��U��u�������'&7f�ֱc.�e�e>rާ�;!��;�$Kr�sr>YW�k�F��Un�{ͪVk�'����W�H!���*��&�}d�|g�P'�ʞ �=��s�f�Ҟ'��E���6᫠�絺�~���;\�t�VyhJԯ%���a���9B<�G=M�C����b�8��"���(��4��XX۴:\�e����a�8O>���ӫ�ܨi1�U�=Ho�U�s3~R�d��=��\.tѾ�LH60�  �%���\�C���`�|خ4;�F���T��ʗZm���A�s2gG,ܓn6��m*�ζ�c['�����I(9`h��xd
��1��t��C]��u{X���67Z=]r'���q�qɑ#�fTp��m+I���5*O2E��zr�l1qCn^�M6��ʣ��C��L������ҙ�Z�v���&5$�J�U/��w&��[@ߣ�;[VJ���8�ٰdz�Ά\�/v&�>W}t.!S�c"�*�t@nnIB�\QT�Y��-D���sV���8k�]-)��:F�`�9�&5ƙb��V3�v�tnL�%���{b�7K�H�`d���`�e][��.��wFj0H ��п�5 �r��2V�oX7��CU�-�=7���+9-C���oQ��K; L�+uL����j7uc�U��DE��V%7o��.R�3zEc�pf��e-�c�����@t[����Ţߪ�yت�ڿy]a}������o�!��K�M�R��!��7ã�>�m��P!^��Y�S�8�k��I���0	�qp/,M�=J��g��S�w�)��+��ɣS�Fhz��8+Ӓ����Co�5�s80��E��J��b��i�Ȥ�`[�*���`���(u�W9����PXu���k�+ݠY�'��$#������]�gG��
e�j@�n�x�Rv7n��,)ux��ʀ��=V��v�V��fimp����j }�:�y�Cs�,k8�X��Qb�Ӭ�9	�q��L�:�� �]����s��P>j�K�P��;u(@�^ B��]j<
8�x+,uƷx�Zp.5��
Cr�O*�Î�x���]p����Fn�u�2�@����+�^0��Mt���M���812��L��ܵ�;ԯ.��o����I0�b�C�gFS��r�@n��E�D���	�tQ�1s�own:��]/�R�,�N������9rMx.�P.r��Fm�����B*_l� ��1g�|Y�ؾ��U�L����[r��4&1Z�Lv3w���H�\�c�&(;��MuG��vX3��}��uwt��!G
�K'V�'d	HeFNp*�6�k)����V��w|w>|6ۼ�k�ܭ.ɉ>:/�}���;V�q/s`Ѷy�2u�nc�f��2ġ���(:���R�ƅ����_v>��f�7Gt�]����0��:���'�z'Iwh�!W��:|�y>�{��3�.���{�{RJx�U89�1~2����;C��	�K�q� [�ŝ��\ͫZkyb��3i�窆�)3]�V��>� ݎ�j�2 �f�+뇜�Q�����ޭںqeY�v*xߑ�Cq�Gh�aY�*���s�x��|��[�#���)��y����"C�}����O39���t1���^�õ|��|_W�׌V<@	Ǘ�P�P���1x��p9�<��|��r,/t����5c�;z�Rv��Q���ѐ���	��Qv1�Cx�B�J����s�k�&j9�	jA:8a�+��3r�{41��zI.ɭ�َ,�k�"6ad��)4�X��[�q�%0iLAM�G�u򽝘;�d��PhIUR����NN�+�+O�6��2�էx4_&DT�=õ��x^�mW�Fe>��[N=^wWW:r��`��6��r�>r����S �M�"�8�]�Mh�W���u���ͬ52v%�)��R��.��-�4
�{�b�-Ǔ`�Ic���!*1
�N�k�޻�=��R�\�v��U_|���S3�o���U���h+�^�s��i^0���:�S�o�1�T��v�����1���9!�J����T�w&]ʾ�]m|�6����Ҕ�d�t��1�k�@���bp5]�t�;�'���� ���=�c�!
��dvӮ꘸����q�\l�6�Q�	]�3؏,�m�!.΋�A��Q�P�^�a+�Uc��)��[=ES�$!@�S�5�[�s�����h��/�kG,�5�Ջ�-��d���J���4'�W��K�5+%�_�k�O ��c�\)�{1~���9f�T�qz[s�4���MC{wŰ�/jz��<o��fg�νc
&V�@oO����F�+;�E#�saԮ��g���y����FU�X���J�T�?}N�obg�����0��^;��\����1C�$ji��oE�6��$�G��c�B�é�a��S5%�Ƀ���WB�N����m�̃6R��Q�����(
�Ơ��v
`�$0��1�r����R�.l+��d���=W�#�/CE��.}�3�$S�0�����h�F�nl�r�Լ~��ݓ�1����r�@k�
�J���}WH��&.�w���f���5��U�=7X�=�=n�iu�\��#�vEѤkg��S�5������ݫ%��?�����������J<��ˢ�W�FС��!G�����)���.��_9�t�	g�	|�W*W�{�f:����}�6}�C	��v���$߆�
�� �!DW���FU<
7��|5,�ǵ��\��1��!h�>Y��w>�+Wړ���`�C�K>�b�Qr��i2W��K��z"�?w=+���DX6o�)�weѵ\�R�åo[c�����຦���(jt�S��f�_��%�F�!]YB��0�h��{�}a��v��i���'��=���L�,�[n�=.#[��mƳ�ug���x�����i�ٖ�{��j���;301=���H�r�f��\4��n�cn�j�u�i��}�^:d�W�ۛ��#֚���[[�k�T���-g�
C9zYc��-�c_A�<:!7M�dFA��}�[���.
qev
�R�����5�~��|�owXd����0`YD�J{tߦf�w��]����N��r��	��t�:"Ivd�$��GT8P��F=w��,��k*YK��g�u�x�d���z�3'���#{k���V<���|����q���������}u�A��_n�烺L���N�_m�T��pL�ױ�z�l�)i�zU��"�<��/jֆ�2�����qNe�wW[�}�E~����ɜ�<�͵�+�������|2O��`%~sP�:y�.u=2M6���GR��yY�{��g(1�X�w�X�R�GQ�>�EKBa�]���mT��ONB���Õ���|����9���F,����D������1��'D��Icz6h�l�rZ�^LMoE9T�NQڜ���l�	�%��c�#���R�1Y/>㪪+�`���X���S{;�)�!��dk��ס���电b�bb�y��j���U�V����nܚOZ�}�����&�q��k3�hp��^���+�8��y���E�|��f'Z�瞙�b~����V�C���c��in���S
�rEo[?<�:ꮚ���m!���%����j A~�@I�^�~)M��Pt��v0Q�,W2bQ};ۜ�!y���MH��Pd���/�{M�5۩4�����NG:�2Ǝ�=�F�F�A_X�5�9wGEd �N�8|�Rɇ��+�X�q̱׎��E�;»�0���X���[��{uھ���^�t��
]�Υ/>�[�įK|�!�tv�r�B�R�ɐ�긎�;�:�Bno�+��g�&�%˔��ǹ����.et05I��ĵS}Y�v�����c��/�NH�Q�:}�c��
�[F	=�ﾯ���g[�=��̜��U1Vhe�T��aP'�i��ue�e��kw��V�����j����ʅE�ܭ�����渨��qZ�pyк5��I֮�U�9��yPhX����K6��V;OiAŷLF��r��j3���3�)�c9r{$FE�D((����+EN���rwlT�f�Rtr�	�!cyuB�.I��=��r�c9U8�o�Y���������U>�*@8},�����1�3e����*��B�5
�^>471�~��B�g����G{5g.KϾl�Frt�؝x��v���8g�#oD�-�#��+��{�͍ŝ�#�(p4��
u��-t��Z��C}�ٯ,����T�K�5��2��s�V��U�+� .7��$FQ��C:���k������m�f8 �<�i��>���ݫ3���nk��v0����F+ו3(@Q�����j���Y�jt�"�x#p�LB��l�:M��O�u
���f*�tmT�ܘ(�^�ny���
U��>IJH]�vcz��ѡu�k���W\�	I�k���٣�IG^���fh-�'g�Jl��H���3��
��e.X|��������[+/�W*j�3;����q+�!�uպ�v����p�P��Q:�ݠs,v�3VKVԏ�V�������7�.��dK-WD�uQ�:EAX��t�(���6M�v�[�x�c�����@�,�kR�b��T��\4;V�@��=�Q�ϵ��cӲ�+�ෆ�����A2mL��q�]c�������U�X��I�5Kѕ�ܕe
zw��o�BQ�ĺ˴�@���o<WX-W.
B�9c� >ɫ4�#���!�������;�T��u�j�+���O8�S1���y��:vj����[L3��'��;r��Keer�ʼ]�ƺw7�4�hn�:L#	*��Z�Tp�5"5��
k:�o,M�&e@�� (z;<rm�+/*�yͅC*_i��o]��N��em'�ͬցp�&�s�GX72���g[<c*(%��҄�Ytj2@��!y�c�D�\$����u��H;Fl���-�)�ܻ���i�oX��qȍ�}R����@m�X�������Ƒb�^LZ��tq��/�š�˵�k0�NA*��}��ůe�a*���gu�Q;/%.���E��*8��"�k���+5sz��k�vx�D�c��X���vr���/ih��)���l��Jo�\���j�r�:a����.���K�Rӏ'��\q%������{b��չΖ�S����)ma�׊���C�����͓-��àeE��t3K%H[#�D��wܩLg.��צ'������A�zԭ�7�A��2Q��[R�֞V��}�s��c]/��,�6tO�9x�k⁮��u�z���y��6ÚրJ-s�!s-�Hg3����^��Ey)����`�B�7)����1�ʾ.Y�B�k���e������w��'i����@���7�K2�bw΢�B9e�t�#\�M�ź�������Ud�0��K�W_%�e	�%�G����k�#��og1�Ws��gV8�
�R¢�c����Z_Lp\s-�`Ռ���zY�Z
d iI���$��u�n�T�k�
����/uv������^�2�Xg+�&���,.��s[����-�/�w��m�r��M)�������c�@�J�w��!�6��[�Y�U��uV�Y��\�w�1�\�,-���L'ڸV�]��J��i�="ǎ��`Ʀa��E x;�iM��vM��7W�a�_5�,1K^�V4P�$v���~F�ʛ\9����Z�` v������κ�[|��ެ�Gݣ�=X#n�:�o1u_k ��l0{x��ϱ)���FT��Č�٤[W8���Rǻ��� �{)9�,�� ��x�Z�{:�#���yQ�d���E�.���y]ҋ�����t�%ɉ/q�qY�AJ,�]�mmE��.<��*��<7d���͙�~y^w皢�J������j h������,����&b!����\"���01�������(J��(�b*�,*������ �*������������)�H3&
 �ʢ*�$2
��%�%)��,�"��*��0��`���"��)�*
��,�*H�h�%�
r��!��2�(���̡*��j��,�3,�	�*����b		��'3 �i��30�0���*b*`�̪�lȈk3#'*���k#*��22Ȋ��j�̌�1��2	��2�J#!�� �2���������232�')"����"!�,�(����I�0�(��
�����&��,J)2ʨ*(�rH)"Y�i��h)�**�)��#,2̱f����"�""���������*��2��j�3�"����)"���,��,b�"	(�
)��(PGf�۵�X�yצ���n˴�,=��&��v��b�T�i��Pn5Y�h#�-��׀5vFN��B�f������F�f�Cz�
%ݓRk��(�3U@W��ˁqε��j�]1�i���vƄ��o�=[4�b����s�m�@y>~ N��k�Ek�&j9�	jps�P�bG��iOu����1}��c�)�#�,܅���C���*�&�dnlA��WS��>L9҉�Svm��[�!�ᾬl��d���J�c���v����������;Y��.�����ɾH0���G+=�s��.?<J����
�4:�SԖQ:t�ݮ��r��Sj6��;^���ͽ����s :�4�S퓍ӈt��ʻJ��0x\Fl�\���UiƘ�iL�VzUX}���*�}��N��b�$cp�u�(ͣsL��	J�WY��=l����Ǖn<˖b�c� �K	\V9)��g����bMH`�og8������v�u�k���g=F��4
;�X�[2���7ԃ����hO���c�w�[�ܞ��]�F���޲%c�i���~� v�����cL��`�AL�V`��(vc���[C׆f
�ï2�"��(�����ej�����w���@C�9 �Q�f�q����` �k9����ޤ�py�����S�u��"�/�&��y�'69��T2.��Ƈu�2�f���p�c봸n��oވ���A�Z�Ck����´�%����0�����>Xo��Go��k:vD�X}����y?f)�gƯ�L���-o�0t�F[M���9D** ��s�ۉ��}����7c��f�@ݭ�#C��M��H�R�R��z��Y�2��9m��¨]���C����e?��}�v�����lJ��C�ꡋ�9AԞ2
S�\�]��(*z���:�D��S��홳a܃}wU'ɒ��P9�cC�p�s�1�3�wos.y*�&�a&6P��[t��&s֬X�nch�����	"q�*��W
�o�[�Z�� X���oF�m�
c'�Z0JY��w>�+V��zŻ�7�mc޽���\��e�9�c���"��hɇGǳ���um��.9W�]SI�J)	,��Rt���T}���*Vk�������%l�4i]YB�ٍ��W2�mN�gcA�0Y���qr�:�q�xX�9�E�{��5�����oy�wLֹ�3�~s<"W��c6H�����7�9�=PT�6)�{�3Iw:s5�Ո)uuۺ��T�b-�ROz�̹X��Vk�1����W�,־3j��������@��1W,zF��m�����ݺ"�\7��NdB�l�oa ofZ�]M�鱕��S��}D+�#��{��X�n�w������8�H��s��GL�ŕ4��n�cn�j�]ƙ���t�w0�NO2���R�X8��eSqJ���P;�	f�L�*�f԰ٸ�u�엿Ug5E/g��%-r.�t\{;�B��v:�*HV�M�>C�U*�T��G�W�m)��c���M���3:q��8t\s�$�@N�Ǒ��*K�$�-����
B̖�ͥT�k̩x^�c�����}p�Oh�tϻ��<�z�վ$J;��m�lB.�2U�eti
�>������m
�h8��c/'Qۅ�ءp'jxZb`3O$�J�T!�P(�8�'�Rz��r�ѕ�����J�2�y�OV
��Z^��%]�и�N� �)��V�,h��=��M��y��׆�A@b�� 
j{ �u1�g0L�e��UX��J]h��͗��reN�g�PϑC��5��O=&�U�W�X �]�#����>'�}e�]v�ez�%�'�c��SD����2�����P���%,��Y�3��V����Fu��tڸ}z<e���GƱ{)S��i���it�E�{J9�*���c��n�XL��X�zAۇi�M�5���YX6kc�E+L�w_�z���`�}��Q�KA��!/�t�XS�82���bŇ�v�@�ڽ�R���9k	�2V�*^�o��T��DG���X�6�d��'��p%o
�Z��0-N&�]H}���x8Ӕ�ˉ���W�V:J�{/��[�]�P~{U��)�`���lm�xRuƠ>��.�	GԪƝ���Cc�f���Ӫj��~��n�Mh�Ի� k�:��>N���o-	�u�gY�2��e��θ���
������$�'��[��?Y�����L�<�:A��1�py��)&}[�Rt6��E�cٞi�˃�,[9)�
]U���-0f5֣q�Q�p+,wIW�y�������OL>:2)�m�W�e�u�X� GnJ�T��|�=i�P�5�dsֶ�ڊ��t��~�E
�������Wj����(�K�4�"��x�N������Ӥ��LM�IMJ��:�Ժ��9rM�
 �U�ͲTu�h�	Vp�uK+���4�w;�c1"�H��N���͗�hcBx�0!t9�P)ă�܆�4�r�,ݬ;j�*��g�w(��Di��\FN������~g�#oD�-M�՛�����e��G�x��ӥ9�T���b�*gWƳ�`��3T�k)(q��ed$gtt\<?s�f������=�`&Y��g�k�����]�Q]��<���<�s~�a;�U�\�N���%N�.�V>��{x�7"�ԍ�]jtB�W���=�y�[z);��"����b�Ԁ�mY��{�uxE��.�,���X��nˑVy�5k{{FW.8����t x�,w(��Q��:Y�P}�l���=+;�U���ow��<�֟\���g"�X�t#.Q���7��"��Xo��w j�3ʸ��{�ڡͬة�!�vY=��"bp�V������(܂��V�s�S����zc����e:�M�K�o7�+�2��!U)lU�S�b<mQ�*�mm�D���.��d��}(�=���SMV�((k��͢�9�럀gz �ʅ����AYǒ��v �ȭ���PҰN�� ���6�g^Lh�/{*���.�P�X�)��9K��w�_IɈ�a��������.[�!��W�4$��Z�y묪X�����śdq0����g�Ob��F�8Ƚ�>�n���(M�E�{Z
�q{��~��"��*�X1��y`�l(������`�t��{ӌŇ��o#՛z6�a�O=���JU>�8ۈu�[���C�$�tm֒5\�y�Eɝ7o���N��|t�(0|�D���١��JWh��*�y	�`-�P ��	��.��v��87���-v�Sq^$G�<���-�:yI.�wj��I��X��i�����k���y�8D�4j�B: ۾�*�����./ж1� >S�@�F5閊ȉUa�:b���oE:	�7�\h)mI&��s;��8�7+�ڠ�btc� ׺XJ�UX�Br�e��V[�$�:/`O� |��n�2�׭��F��j�k
F�G}�X��rٜ>h���A����vv��*^��T1b�&A���I���b�1R�T�{����T��s�#zX��Rv�l�擓�|�8��&gb[�㋤�,�=wa>/��_u�@��%E�k�	/^�[�����R�vD�ط)���B%��q��},�&k�(�^�W�����-��5wוS�t�t^�.�ؙ��c��)�E�H�Q	�n�`������z/]f;Q�sN(��B8{��==��z/�-)��|��y��$�\�`�1M��w���������/��Ζ��R��I�K��^�^���{�@5�grݫ�~�X�G����C���$<�q�Sï���A��������u	��M��ryfb��N���{���g�8}���T+���]Mڌ��������/]b|�I���>�ɚНB{���GҞ����r|������<����ey=����:����C�ԝ}�r]��>?}��s�3GՋ��NQ�u2ݏU�Q�U�3;���x�ӄ=U����|oN��E��>�7��7�V%Pz��K�v�k�uN�����`C#ݽ\������7'dw%٫2������(Kbv��݌��*�q����/�>����2�����{�
�Z�y�.���=#��ݨ�������25!����5'/��НB{��=��/��<���y>ǟ���c����=Ò�y#�~�����(F�9�[���Ǽ�ďG�@����~�ڴO��C��:�y��L�Hx}��MN�鹈y)�zg4S俠�_�X;���>G~b;��T@ߍ���WahY���C�����a�y@��7-�!�x�7.��|�Н�s�'�쎣����&F�:<�`u:���7�<���`y/S�}p�t�UG�����?{�=#�z�}�1Oe������ђ��߳P��b�y�/P����=�}���<�e=��|���ԇ���MN��?{�?zs�u5��߳c�x����{ޡ�����>�~:��-�����4�a�����y��{>�@nM�%�kz�9'��s�#����N��S��B�ztO�m6�Rܸ��k5��C��R���nW�?G3zN��]]����nRu-/���P���}�V����n@��>�7&�r���{��{���5�caf���w��˾�#�=��ރs����=�@nMK��o_J��q��i:�+�kx���'�X�C�pv��j�?G��z��7&�1���1�ک����,�o��s�z#�7K�{��Ӹ-�J})��td�K��=�sHnMC�}�#�h�=�{nW����AԼ��c���x�f="!@�9Ms�\���wo�%^@�=����'ѹO���C�9<��b{)���>�}���y����r~�����hw��Zp�ў�=�#�\�G���w�qϳ얔f�~���y;�;���rG�ǘ{;���G���w>Kۿ9ӹ^��{��?@�7�'����y��iwn�Z�����_��(��&����W�m� ,�����=�k-�]Cv!�J�Ɗ�r�ٚw�]�EA�%��uoVM�[��)�n�!N��U5�u`�����%n�+�
�P������3�dB��OvYP�t�w{8I��˻ݺ( ��[�#����� >��t��������qZo1=�����;�����;����>��C���7>K�<���y.�u��^��}s����;Q�=�Ǽ�����$W��o�Y���rZ/c��h��z�A�q�ϱ=��䧽aHw&��;��@�;��Jy!Ә���>AJnNC�J��G��*B"���W^k�z/�v�}���+������C����%���g4@}=gz9H�'a���I��S�_���7<��iOgw��>C���8D|==�=�"m�J�u'���zG�}-�yђ�C�����#�����:�;>�C���n?9�)�'�ۜ�����X�O �S������M���{�x1qٓX���k�u�FΥ�u	��$�jd>����s�����:\��߹��]Hw���	�9G�֔����j�`|�"4D1���"�3�"i��˟�}���k<:�=Iܟ�Sܯ��7.��<��K�ԝ�9-[�4-���s�GS߼��&F�:��������Ϫ��}.�]�2���q�����IS���:���|��r]����F�����5// {}ǐ���]�d%׆�д�擸܎���i}�(�荺Y�ࡷl�U����sAhߡ�jO���hOe7��O��rw.O���r�k��ewђ��#��ZC���]�d��=o����v������������V��+���GSÞ�}�`�C����S��=�Z��^�֓�z�`=:��K��w�)�h5����>�%�x/�DC�����,��6�?�w���k\ПI�s��H��������[���Ի���H�'���h:��u���Oe��&��^G��y�nXDNA����-������Ms"|b{��99@��Y�����v=�1*��+8U�+�R��4�)"*�⫔n�9�aD����teZ5����z.��R12���Y�f�73yb�u��I��!H��S,ξ�o-��A�N�fj�$�G���UU}�Ut��&ٹ���=䏣�?C>��z>�z��i{��G�}Δ��sO �S�>:�ܚ�"�{+ܟG�sA��G���W�eJ
���_}%�=�)?nsC�w�~��G_�����8'����>}���~Ò}���}�rM����{)����:�N���w��;����9&�ȷ�H�Z<�A�nW���=��3s�����/m�1��>���`B=Qz��9���P����������ݹ]��=���{y��;�O�9�K��G�a�y.O��o��5.LS�����!�:k6���ɬ7��{�Z<�Oײ9�A���`j�?[��xp�Iӭ��G�{<Ǔ������ϒ�o�tH�'o9�{�<ǣ��^3|�'���7ڏZ[G�2j\�����\����z�пKGA�h9}A۞�<�~⟺�Mǰw��C�u���S��gprS��Gޏ���3~uu���ڥ[S�{ez���·��G������|�K������@}�I�pZ����U	ԛ� ���Jy�0����De�`��}���:G�c�"0����w/7��~�俎u�C�r�k�iun�|�w!�y�g� >���O#���]i<�w�?���;���.s<������9��׼�9߇��{�y���u)����r}��ܜ�����J�^��˒9~w֗�y�!�}և�C�q��hN�>�����!��E��-oןm��T�q٧�E�`��u�y��1�#���<��ԧ�nNK����Cp���4d/%��u���-����/:�;��p���By����G,8�c����\�'�⟤=��G��K�X���y)�]���Oѩ�Wq��<��ԧ^�iyj��9.h����כ�K�a���
>?���� �K^���5�.��>��u.�6K캋kˏ���7)�����d��U�p���W��	3	otG�\�vw}�5�:�fEǄ�D�k!��.�1��G�]�%����5L�.z8���֫s��}p=9ʄ����U]��L�w�=Cё��~���	�>���kHy)���������O'�~���x~�y'�ty�S܎���u#�g����>��P�G�=+�/����=U�t;js&��-�}�I�<������ɖ�:<ރ�&�P}��!���sT�/��R�N���y�#�9'���]��������\��lI�_ɴ.�sO׽m����K��x}�j�ut����'a���=���~���z����>��������dz��%�}����~�/��0�I�w�����=����o�|��vp�>��Na�|�#������p���������<�I�{)�ޗ���;��>��O"�&���zeϣDz��z �U��I��_Ww�y��������k�s��7/��}�5�7�7��'$�=�9қ���9�r~�����}��w?�u�{��D)ϷƸ͊���7����3���#�s�4�C�9	���iy}>BjC�y�����~�rn9#��М�v����=�};��s�>��7����y����\��ոC`��f�C���#�w�B��s�ϴ\��9�&���'�c��w�O���������<����nGWi���w/|�}{��G��`ʍ�sA��&���X���]��� yϵ�{.O!���R�˽��w=���/����'P��S�X���s�xp�Aֳq�c��Cǽ<������#�%�j��{��y��9#�:oޗ��G�td�Ó�{w�%�ݻ�\л���}��{��]��59ԛ�$vb"�z>�������I߶Vg����5Jy!���=�@����!��!�ߜ�ܯRvs�z^����-����K����ٯ�$>��惟b�����)'���_��}�=�<�����3S�8ʦ�urW����ʥ�YOm+�sY+���ͷMX��MCI�#�Mi�V�F�v~i�*"{=<�9�^(�!�l��T��}�f�SR�"[�P[ųԉ
��z�}��;�W(E9�PW�w�K�c#.��;�H-3�݄Uiݳu�[EP�׀P�n<��a�9��4��q�j�3���熶� �\��^�Aj`�{5]K�N!�J}�D���� y;��D�$l�Ca�C0֩A��K0����gm���t� �h���#�ٷ�Q��3`}�Pg1n��iD�ֵ��&D�Mx}��fAL,zE������+b�'�5�l��~]Y*�ރp�\꽫;:�	d��J������[���dqyx������`ʱ�{�����N>�!|v�%��=K6����-ۮrN�d�7�����k��ҝ�z�� �뺖�n]��;m�����6�jh�l�۴�P�R��,��p�kP�v�{�n���-��S75�(`�Aαws�N��Q�'�_JZ-����]f�3�C��7+�<wC!CR۔�K5�U��`�|�EW�1�`9�=�Sж����m˥ u�h�[�%�ڔ✖�7+�6��E���z�Y=&��A�f��"}+m�60aX5���Q6��g�ee�톍]0���E�v�Yâ��Cw@�NL��$Ԫ�Ph�U	SK꓍�>�'[��k!�;�؇�w� �W��eC��5�M8��6�Eʇ����j��J���\������٦��ݺކ�G��ҳ٫E'qڋ�dtuY�49���+�+8�	�Ή�.[��6�U73f����2N����O���Y٧R�9pΩ�G����nc4)��(U1�r�C�e��Z�T���y^wf�L7�*����wr*K*���[�����A���D��*�R�l�DT3p��Ǎ�
b�a�ME��G{�В��1����b~�q�@iОj���=��U�E۔9�=YP���WT�a�!��X'�'�1U�q��J��*�!�3��v���w���݂$�u��c��w_}�+@��g*v�7#�c'n��X3�#� ּ%�n���û��3���1S�c�y����d���i%Yɧ��z����Ji�8�kc.v{�������j)͊�$�,�1{ڵ��栰G��dt��u']�/���/	j��r����h����I��m�=��:a�B�����g8�e�t�uGt
?t�f�WF�<�z���n���N��]W�Rɕ� ����LŻǦ�yK/�.�,�Y�%��`��m�:[ĐZʱ���VC(̲+��uv��WSh��2��u�jiu��4�Ľ���L��#�@.����ͫ\k��r.���J��o-S4��EWZ	�9]V��}k�p��wm��R[	IKry��AAE1�eUDMUEMIQ%QKUQT�LMTDQEc34DMK5%DAPQ��9DdUIFF1CUE$�Q6fM�8PQ���L���TYdPVX9��U��d�ĕA4TQLDM10�T�VT�XSY��AUUQe�DT�DUTQQ��LMQT4�DD5U!M��E�aASDD�IU4RAPSQPTDQQEUTLPY�M	ESEMDQM15AE�5QLD�5DT�ESE�%MTUT��DUQQTEQCA�SIEQSM4�DLQQUD�U@L�EMTTED�IIITQAQT�D�QDO�����~�
�~�i�ۆ�{YSP�kB�\r��2< .���_����j����9��ƅ���M�X,Y󏪕Q��~�{���y��(N���O���'��w���C�����/'�<L�9'�w���Ԟo�t�ܕ�~��������R�~�4�@}��y����S�W���=�q?D`���T�!��)��(N�s���ť<�w^a伃���y.O�w����o}�����|��9�z��ԅ�o�<��ky�|��V��Uj�ފG���ǧދ}�~��z�5��M��O��hӸ9�1iΏ�~���'_�7'!���!�iu���%y|�w�t�s����c�Kx���4}� ���=�菝O��5&���f�'P���yJy/��=���}w�<����Ó�'��e�u)׸nZF��������o����7޷��?�iy�|�$rC��~�s�V�>ޗ�25!��4�5'/��kBu	�w�k �S�{u���K��;�ܟ��:��w<�ǹ��o7ÿ7�}租w�~�?K���䴿Z����7.��t���C��:����25!���~���~����S��9��%����r~�'ȿxtw���y�}����ٮ���9&���~��FK�~��9-��x�7.�;�;G�'s�'�쎣�b�&F�=<�`uzDB�F�G����� �3'vK�1vw�=���ܾN�8u�쟡��;�䴚���eya�}�����1}�4�@rO����H����7�y�{z5�1�"�D7�hG�p�V|g�>���׼w)�����A��W|�A�ϰ��?KC��{<�w&�a�����>�����r^:އ�N^���W��#ѱ��~<�럧��}cy�����7':�K��=K�~�kr���~s�N��]]����n��'r��}=�`�@rO���ZO�;�ې:�D1�b����
�oo~�Sԑ������x6��w��-�;�Y�Iʇv�Bo���6��J�c���#Ůk.E"C�¾�Z8+e�W���Yw=����[Ϛ�Vmf>C7�t�,Q�Bt����;�ц�t���v�����J /�u����O��v�u�Z_�œ��z#ނs;�,�|2��z�z8y�_y�w)��9�r~��=�þhɩr-�ҽɸ�9��䯑�:ރ�F�?`w-����	����������KĲ��YG'Vot��o����E��{#�q��=���������:S�N�{�$�\�a���Crj��>�H�Z;3�'��|�u��y��>�=��Eo�ÏH��VVN}\b����ӂ{Ԝ?oG�=�w�I�rS��y�{���4��}<���'r<���r}�f���;����(��81���۬��SZ�V~%���Y����z��{�EH���!���x�p���Y���;|�����?`����{7�:w+ԝ��ޗ��|�$�\��<�䴻�o��s����V8's��6�\��""��O�8���^��yy)��(N��{'o��NO.���$(�ϒ����	�<�<����z7ξ�z����q�.�|��N�N�wݻ*�L�ޑ=}�=����?h��z����N��'�r=����rn>�������y)�Y��?K����nNC��~�������ؓ�֨JWVL��������U/����z��X�zއ��{���9�����}#ԝ�'�n<��x�pny'�������1�N�5�j뫿�]�?}�浱�>�C���#�">%������^C�u��rG#z��:�=~�C���n?�)�'�ٜ������'��<��X���'��Ͼ*������;y��8������ƅ�u	���r�~�䴾}�d�@}���瘭v��/���C��Z{�Ԝ���ҝB{2�`K��y�2Í"�}ڣo��"4{��#�^O��<����+�������q�4��IѼC����B���:\���{�/�djC����!�9�����K����z��pϟ�C�b�~��*�/MU�R`���Q�;�tf�a������L��z�e��� Kr��)dS�I8}ԟ䏤�\�muD�$*D��[f�v�_u�7yr <�r��V�,l���ծ�',��宆8Upɕ�P�9�l���}�G��]y�����������~��P{)�_�Iܹ?���y&�������{����o��_7�ټP�]�G�Dj���`��H��7���n�FSYC�}�οqz�#R��G%5����'���y�Py�송�˓���h=?a��Wp}.��>{֐�{~>�G���ǣ�(��D���wls߾����G�N߽'��:������=�@�u=Ϧ���~�볝��K���:��K��w�)�h5�ޏG��W�����c������mM����w�p�I�p�|�Н������>��������.����y?����]w��Oe��'�;���{G�{�D:��[����U�5S�]�o�;���Z��sչɸ�9�^�9'�߻ҟ@���t��=���Crj\��޽��'���h:�G�FS�E{�N7nB����_�~_�k��4�����PA��~�C��ɸ܎�߱I�ܹ�e>h?�}��,���A�yt�Z����c:�쩿��[G�-}U�I�����z.�oh3���Ԩ\��Z���f�ZEs��#Y��[���0�U��%���+��ڛoF�����}Y��[V�1Y͝��T���W;�9��]���u�������An�4�,u�*l�B�Lgw�>�8�.���{O�]~��YG�1U�Q��oX4�� tIucw��jw:�n����n��i �
����ۘ�S{��`NV(l�y�0��u�N�5����m��&�s�\	���K��1�(<��{���w�G���i�y۵�acSr#|��ވ�Dj�KSbn����[�iO=s8��*������O���}��:�Ľ�ߗ���q��̭B�7�E����L��:�
����k��Y�,�a�W����8�9�9���FEG<r���5)�'/s�+���\����m�&o�fS���'U�S�,෾Wܢ*�M�[�t�X1	���++�ͦGeDV�-�����5�#�)w���3M�F���y�����נ�{<<�ߩ~��kWy�3�l�W�f%}֖�Zצy3�j��`�7��|#�Ŭ������j��$�ޔ�x��Gz����=�F�un�ޚ��ܰ�E�s5͙�Ynj����/��x��E��^�
^kmTE��r%��x]�� {x�,�/=��;�i���s��tN;�%�򉴙�iQU��>q��l5��v���چnd�!����-㌘�� �:�f�4D�q�g�:.ٛ��GX�곕�w��eE�Aw��eݛ��6U�)�sS8>��w
9����A�ďo�������^Ȳᮂ'gv��+�%�;K^�ܴ�r냏b7O�����S�UU�}�}�ȏ�O<Λ�9�~�]j��ˇSj�fҺ=|�"�F�Er
���s�7o7��|6fy8��]�ᣩ6CEF՛%Y�EW��'�B�g�kY�odU�8��C�-���ѡ���F�����&>��╝�Wf��+���j�X��9�����;<��{&�sz��.���:�n�B�A��������^(q�u8)9-]F����$�ھ���oY�gF���Ejۘ��q�s���JC�No�9Y��vҷ$ʙ�ϢT���yZ���m}s�'z�Dgx{(uKz�:��ԡ��ushK{#"�b������ySX����:ROx�z�D�j{2j8�˃腼����v_@:��uAq�G��{}=�]���fWDw�y9]Њ,��[k���d��^\a�Z=�]iξ����Beޭ�.�jl3��d�H�^W�w���4����|�*6�MLÆ��nvx>�����ƅfWr��Ŝ�$�f��i�wN2rLf*I�`o>��݊���;D|ʎ���n���Y}�G�WK�j�X.N˳F��tΒf���99۳Z���_��z=����V��n�}�rw�8��k�u�4��7�o���zOtqH��U�k���ҟ_��3a�6��P���5lqx�/z1��k7k��U�jk+5�@���ń��I�ڵ��צ��<���);*��u.3m��0��g.;ȔL��?F�9��W�h߲��j�jJ�s��kY�]=*����BX�ګQ�����6���M!u����ʛFc������4ͮ�=;֜���Vk���ZJ��W��W��Q�#���.K�AM�{>��K+9*��fM���i�E��57y��}��P�BL�ڜ�dqx��J�M�:���o\�_���>�)�����z��Җ�K�״�b�5�3:�R���?y��1c���u�A��@�ͽ�Z�g9�4�/��$B�x��*��`��Lgd��{�F^ܹG�,7�T���p��ь�3F�Kcrt��{�-@&OC]s�F眝�0G�U��kq��k��Bs��hn�G�c}�"������3L�����]�r\b��X�Pik����B��yXP�`M"�a����-J������Z��T��DDG��|�%:�H<�o?t�+�9B!-��L
~(Y��[����I�'����̓��1�ќ��m��%�v�7�_�(�*�#��0�F=�S����9�7�c[�^rc��B�/��δ�����ޞ�^}(��Ppæ$7�����' ��}��:�\:�9��iSͷ�᥀�p��P����4�K���ȳI�AkXQح�˫}kGbXb���v3��	���$�g��]@��G�]��\��U
h�̥�M~��F��~�~3Ƀ]���~��1��ZǍƺ�h���˳`e��z���خ��E洦�l�;��n�T������ڹ�P}O:A@=�}���Xݽa�͉���1��iQT���Um�ܖ�������@F�x$��ec���G]뉨j�����;�*+y_�|�-��M����5���(��{�r�V
Zz0=�U�	��w�wr��q�C����D<�q���+V�ƴ�:7pǼ�2�o�:9.�qͤ���q����:O6��	K�ms:�HǏ���9jgR�t��렻�������F��n�X�����e��W3iH���Ui#Q��7��}�d��êu��n+) �q��*R�}�P�ӫn$�;�WL�X���}R}T��)7׎9J�ɞ�o��֍����0��k:&)m]0���S��-Q�T�"M�޹뭚�t��-؆����+b�צ%mɪ���\.�=�o��fl���:Ju��3���AU���} mj�u���Mu�|��ӕ�bo]�9�c3�ׂz�<��F��t�IQC29�ړ���m]mk���gY�wl%�'=�3�y�r2����}z!!�׻+�s3�4t����f W7k����xK#�W)cj��
����pÞ:eq6k���=���.-��a�
�1ߌ��Q܍��)�֏.Rz*�E�w�u;�~נ�;'�<��g8�]ꗀr�z�;tǾ	N�W��n���!m).�)7�����cJ�[��Dn�e+v6���M�γ��C�v��]K=ZY�q�[�QuM�����F��i��Dg���|&�z�GL��ȭ�j�o
�7��]��{ȭ ʛ9��������fڄ�;��e[�E��7�vk_t�l���/fr�Xj�Kk)�	��{�5�qX�����Cś�䷧~��ѫ�8��	�t�9`�����f��V(7�'^���R�|�Um��Q5FЯ6��Ez;�8���^h�̈p�y�"��w���v��lk�nю�M��Ԭ��z���c}���6D�֣J�&�5ܽG���E��V
�gj��|�h��;y�)���4��sуy��=Hfu�k�U#7���Z���R@Lj��|�݀i��<����ok���J��5�P�Xܱiuqq�Wܥ(�Éd	i�1[ѱ��]�������uݵ@��*&�nĞ:G.��V�Z �{
jk9|f����ܼP�}x/���a���{1�����=Οm���)w��5���gfMߪejЎ�S��-nn�2­9�7V� uY���4y��r`Bǯ�#����L�ض��t�#��MV�^J�c �O�Z5�u;�VwmX1�<Qݓ�]̢��͉��յ#�����1�a�^�\��kN���1��];M]�`Jy����W�P�<�yڞ�a��GHD5��T@��Fqe�nӸ�F�L�a�7X�:��U��U<{K*�lt:�W$iN^��fC��u�D������/?)��'>�4uy�������<�Zg��c9�1���`�;/���27+�q���\�/^� Ν�I�W��f�~ž����N&5��]���d�<�z��ә��PGzIR��c6�������ю�Fi;�o4�s�s�ٹ]�]*T�J|�`�N��)em�J���-��q�Q��7/��ݳCww�o��f�,��s�㯛x���m�V���5u
<�>ת���mŽ�6b���y�ά3]�����Wkc�܋��@9�<ڑ#+(&���[�i�9;�)qp�����o�e�:�W�˕6�&�"���;<Ve�>;]�eU���/��yBzތ\�9�����F��B%Tv&e��EH@�	���-�������ʈ���J�"Hl|w9�[�1M�]"L��C���Y�r��y�K�7�]�M��5��z��d�XW`�,%Jv
�o�\#�B����D��d*:�yrE+�\���D(G2{$n�ᲭT��}|z��;�,O�����I-ʗWY��hU|��V��&R�hF�d<�Po=�M4��1�F�B�Vi��oH�:t��y��s�IR8��7��9�J�J�;٦�*���#�1�Ըv[�.ݬxܗ˥K�p�bl�Hl�	��6�*i`/��͐�9��r)�T7�m���*�c�K��֩�Es��A�:9�d�k����zj�������C�2G\��;"�9p�ڸ�h6�v�K%p5�)�Sr�u�ӳģ�볓������v�b����8f=6q�+��u�yV
�51�i�9r���v�I��S"K��N^*���n��I��{�����6:�Yy�M8�ne��������=�ʀ��ʕuǘ�� {�'j��ɚ���&�3�����&���way��r6�������yϦK�bWѹl��u���B�Nβ:'l�/2)Gv�4�[�#����&fՙ�2R���Y�c���Sm�]@�(��#ݠ20��Xpf`���
�f�ڶ�E�x�p6����k;&���O�-w	m��J��,掤38��k>BE8a��$�w�JɆ�_�oq��kaǮf�n�r��D�}ok��e�Ӛ�V�ϭ�B�d�7E���[Ue�q�jww��W+�#}ûZ�%GtF���;�Dn����p͚J�P7F�u �Ӄ�Z,�tr&�.��us�)�y8� ���"��t��A=Z���_=ˡP��;o�o|��t����d�XF��5uKuus*
�=�F1wW׈c�qj�ia�j����r�4��ˮ���rWqkY��n�{�M٨Y����U{��̖𣏕=ҖMX�)��c=a���5���Vv��]k�ϟb���	Z ���;s�0L���.�ss��<�u��5S�8I��sj�HD*펏�-|�h���n�,h�N���h�G\��.\�\.��R��΂8Yi�����еQ��R��*>ё����A�2�SpE�E��Cn�)��yw��d�A��-u:�Ճ��N�Ce�.qJ���>��^2znw�s��ݬ�^k�{4�+2Q7�f��t�GŻ�:�}9�鵛v�Cc�va��i\�n+j�6.��-�=�y��fn�l��5��;���"�sV�.�����lF�Ӗ9
��m����[|�۰q�d����Y�ގx>�{���V%O�٩�L�w���� �2�m��]�q:�����������Ի��'sj�m\����Z,|�.ź-ot�鈮����@��sY�����"��� ��%SQ$SE�eIAUID3QMD�STd�IHDSA�U��M%%URS0L5E4!TTM)TUETRQa�)JP�EITE5R1%4DQAID�UDAM�CT�A�U-4TEPU4�DT�LUPC5CfVFfDQL�Vf1TEU5U�EVfAUD�D�QAADU14RMTR5TQLJ��I��UR�QTQKS4R4UQPINf5�Q4$IBDUQ�1IIKPIUTUE%%SCSD�`�1U$T�3P�KQE)TD4EIFFUU (P�*����Vn�1�׶�N�c¨c�5*4�tU�!ڰiW��� ŝG����賃E˺�qBm~�����J�è<�8�_U}��z�W�����ڿQS���w����b�|4uD,�fq#"�܉���XmR�s��.$�s=����٩��5e,ji��Z�EY���/;�Kh�5���Tlt��*�c!v�&��5��=�Nh�3{��D�Z�	�U�=���m���Ɉn�X��y����V�4����VV�)/�f@t�;#�[&!u'p�q�#�栩	J����U��'xzP1�:�=2ǒ��ˌ�g��mx8>�a�'8ũ�50{��__�2��rZ2int^=ꅍV�3,�q0_���r�ה���f�>�mfלⳎ2�V��	�)�,/��sxK�+�t$�������W�Mun��x���H�Մ��E�C�]{S�*���k�T�17��Dvi]�'Wv%�W3�H�yso�{~����=L��� �0}Gk�ynQ��Κ�@]��or�Y[�k�A�#x!�W4niysO�\�j���Zi(��;�8�b�J���O���R����,u�V>TWf;*�pȖ����Q��(Ȗ�G��hT�vr�p����έ̠��!!fH��S�����@��w��t�����W��;ð��׵�6�t�8���sWV�괎ð���$jb���	}���y��4������W�F���s�v[ƌ�lɩ�<�Xb��z/�^�f��US����}�-ʾfQf���\�Z��t����O�>�=\!���u�=;��SԺ��Zͨ4șX�-|�5 �8!^ُ��>%�0���/�w]�m�!
�69��kqC��w6��ѡ�D.�*'N�Q�V�I�wꮒ���|F�;��wZ{���#�5�i���`|�BB�3̾��n&)m]3���,3.�5�nh���c~��ZW�Q��re	<)����FY�X8�m"���nws}SY��Ƭ}��U���q�pV�:-�N6��oQ��F�<���VV�m�̗�fV�]�U�rS��C��1%�-z�b���Q5Aץl�RZ�'5��\:Q��!�i��'�n?A�«p-7BR�DU4i���V�l��d�~c�G�=�H��y��V\@�[�z��}��C���]0e�yd�G��cGgu�T��
��}��	�J�*)��a J�#ވɚI�<�`�8����/�h��8��]�f#c����{�56�:�rp�,�ǡ.�L5���M��{���u�\��Pɱ�d�˞j��5�N2:ˇ��EDj�g����6���4|���j��V�*/{���I�{��q��e'��׀�c�z�͠�/oҬbb1=�ڃ������o�6��l�h#�I�BO4�=٨���#�:�ۺ�J핡�}�ը�q��k�q�\V;����w^x�w<�����k�[�t��g�r�c��;<j�(1|�^��AT�ᶥ�KS}	f����u�3���]���;����|��a�&-&k�ңfz�d���V�����<�}X��΀I'�g�ItEw��z"/��=������)��?l<���:���>���;��ɲB�ueƵ��������*������7*kTl�KC�e�c{p l�!�ǆy�j5<�q�7#������2�M��ӗv΃�9�'3���v��,�M��Dz���Y�n2�j
_B�k���׃sl`��W8�)���+�1��'cT��R�
`j����{3�{�Ց{�o�bg⺪癩�y�a����CX! ���i5n��T�o3�jq�M.�YvP���eBƥ�����x!(7�xyߢ�7{'f�;�9-����>/+y���f�������aeR��{�ػ��|��V�fP~��8j�����o�����>��Y�t<A6V4L;x�:9Ϊ�(K]9��B�=!(s�Og�g}�]�"gf��1�������y�CpG�p|�P���v�}�%��;^��vf���ƍ-���y�8�=�(�d��g�^rc�x:/���#r�PY��X{ͯyZ������ϱk�p��f|���la�׀�s�xv&�q�Ef�d��\��^\�X��N����q��Fb��n��Y�ҹv��o��\�d����Y;�.�V(6�WU^;�N_W�J���:E��=&�T�ٗ��)|�U؎�:3���F\�Yo�q|���Gϣ�g��m��*����?\,']�|�N�Zo�}���O[�3fC�C�Y���V'd�jf]�8ފ�O���q[xjfSRS]&d�]�uQ3r�������ֽ�����W7�~���L�X��k�iu�hש��fs0�����Ԩ�I��l�x��tk����E�� �mI�<,= �gM�8�$�^�sZ�`��/������m�nSDO��W�ˉSjȗ;$��'t���g��,�m[��{t�p��x��p�z0msDH�=�"��>��g����kW����7Ow$�B��an��:v6�����ƗpF�%�O���a�8x����u>�O��MK*,K\1#/�n2��Sn�P��r��x�Rx +w��j��@>f��b�Y��K:�+|Ԃ����k�=M���~:`R�^���W`����z�Fn����he@}�-�m�G!�D%���
}5�8��>�[9i�w9�̓]o���#:�m@Ps�t���8�d�*�!R�����oʻp-8��eR�B�S���;u���&�vi��m.>�� P9+�Yb��E�ҋ���~�r��U�����o4-w!u��b��y[�#��Ģ�[[w�_L6>�ݰ�TT���NU�(� � ̀�ŧ�eNa�hRTs��S�=���y�{V��O�w��k^-{��0y�r�����c/���]g��+�q�E+M��(�Î���eFM�f�5C3��$�gx�ms��}�'�V,�K������q���N}�J�K���v�{���goR�%^������y��/5
�3X:�3���S�v��;u��u��V���9���=���7�����{��eiv:[oDˇI����ba�ݎ{��/�V�[����r%k�5~���Db��Q�3��|�z9y�j;�#���Y��IW����V���h���襦K:�k��7�eY�\�j����D��F��TV�Otܑx�S\���g_X��%��{�B�v��՗��4���N�"�F��2���v��U9ɾ�Iqٙ��n��p�����Ѩdiշ&���]+X�U��|��V���\��kgKTu�x�*b��=])�ݳ�y���Ᵹb���<���bj�������Žۥ��,̧�A�սB�w-�Wٽ.�m�s.:=W)ǥ��њ:������N���%2[ٷa�r��F	"�
컸1.fs��gӼ��zf�Ԟ��J��O�}qm�Rۀ��9�o|Wf��+T6�c�����K�i�O7B�P[��{��V���K�NWk���.1����x;�J��9�v�AU��.��ڳ����o�uY��oi��y�!NLgfK͙Z�t#yT@t9)������Oxa�n�8��&�7�uux[飏*k\c
s$�&�!G{*���j���ŭ�	��O��]1;��sά�=����s@2�z�����`�udT��&�����}�����y�}`�:� ⷹo9�}fx����}���r��HgA˥pu�Y��/fU�����3W Ƕ�i�m�3�)�V{���L�c�PrcŠ��N�'�y�Nƾ&䌎s�V�a��\Z����/�7եP��޺�:���c�n�^�un���0v�E�:�T�QݯV�����%OAf����Ren�p�(Ӷ��
ſfs�{]��-�3��sf�;���),_<����y�39q=�� VL+qt_Z��<9#v7���νJl;�'ѥ��4jvV��N�}q����EqР��ir�;���~�{�O�[]sp��A����]�
����C�g��R5���9�Q0��F����5}�!���Sj棺�\��E����Yd7Ʈ娾}��Z�\��oG.�M����!�҆.��JJwJgxw\��j)��{����V���E���NgsᣫЛ!�)^�W�R�t�o�����Q���u�WL�Yq��<�>ok���J�Z�
���ʥ�����鷑���/�\�{qT�����v���M9�������&�;χ�=�Ĝ��y���X7^\LRڋ�U/$j���R��k{`���&.ҭmF�j�4��:�����
�<���[�is������o)�(�O��em+�8}C��q!p�`�:��j��T��d-���d�>�٪�{K����<��dW<sQ�%��u
��[1K�o� ʱ�o��ngͨ�̸9,mY��p��H�]F`�y��j��n΅5n��.�E=��Rn4=�#'��0�Ú��9"�s��0�#{T��4�#�U�/1](��a�]�*�\���˭`��u�8�m�ڹ�:8����>�܊t����&cT31�3��Ȯx�;.�����N�9�xy���x8cFd�M=f�\#*YI�F�0�{NL6�4�inU�-<�=��=i��ZW�γ:n�=s64u���GRE�+�vg�1h�y�����yO�Y���-�᫃�o�w����<��IX����OB�����?@�Luڵ��ע�UG�����́~Y����������o��Sۆ��Ks�n�a�ˀ�[(�v���s��n��7�������5�*����ɥ����Z�/���;�6�kcw�Y�蚏�F�"��z�F���TV�=7y�������V�[Ev4�c�C㝖�^�Im�]U���N����Rp�ڕ���d�kk:�"�n�P�{uӫ����
�����|��}x�tb�5���x�w ��9բNaܑ.v��=i�%������\JI�ں�
\�˨*FZ�Ք��Vb���Y\2ڥ�'T}���k:!�����Y�k�Y.���]\V�Yh�Ո��h
�4���:��C����<�:����;9����+�y������{uY�YR۞DՉ�O4縪�L^�/��NY�fmt�v�AI�o����h�{s�/�0�ީ``��w+�M�〬exr���m�oQ�s^�2R�;E>�<,U�=[kg�Ǻ�6���\*�����~V��)���rS��B�����6`N��C���7�sӯ](��D1x�^}��}�
��R�U�X=�w�����\{���9�L�
��:�xn!y�0�fZ�!�%��uӶ_CT'w{�pw�/*��j`3��Vm@q�����4��^mH������w��u;Շ
y�����8��؆sa�^����N�e9���fo#{J���q��C���[i�ŧ�nݝ|Mo�Y[zz�W�aΆ�.V�<���	�A�[�;���pվ����]��[��>ܯC�L�^`����ͭ�����[��"{o���暶����d��)�=�;t[�-oL�D&��Ɓټ㛯 �[-�GU9s���:5�+N����+1����E]��MV�ln��VP�����<�]�V�^w%}3�DUd%7��4R4v��,��NM�<��u@��|�PF޽o���f��m�DM��Y���K{��2�]���|�bV�or��>�g;9��ݝ����oM�'��ޛJ�R�#QcB��PGha��'q�svu��[�-��"7�wo�#|����y��Zr���u�,-�{MֆB7��&��X�i���.H2U7���8��[iղ�'��;��b�
���4�io<����S�#��X��Iu��b�?g%���m���h��:�hv�p�*�KA���j4�&m��M�f5�D6iŎ��U4�f-o{3�k=��}8b�n�_�P;9ZY�P�lY��w�z��u+&��(l��]\/��C!#V�ǖ;.멛�	e� �B\v�Z�Md��o`;PV��79�'0e͸���R��Hݩ��ˬ�7�6*S��֊w-77vl�;�X���������0ٔ\�yQ_�bא�j�<oQbt�3);��M��խޣ0V02�N7A�M��֭�Vۮ��ۦ�����m'��3��,�\.������[x�eZϧe�ͥb�EYQ�:�R͡Lt����6JU�d�S�����똟3�w"Pj��ɝ�h��P8�3X+lm�]K��0�e�(���-��f���V�{T�­�D��!Ƙ�2uiX�i-wN��38������^�w�<��$'��t1[X��o'����:;��d�HJm:�/�����/uvs�I��v�����c��L=�qF�9/��[i�S��G[ya@ݣ�oA� �m�M\%��(<�����4+� ��ѽce]+�v���;��gz�;�-�0�Gic�<����š��^�H�T�t���]�p���鬵 �Sp=�e)�7�+�^S��r�.)�Yٽ2��H���"K}��ͣ�:'$#6��bV;䳞�Ҳ[k)XG�k��vZw�;���Q�Wm�	�n�|�x�72k��f"�:P�T&�d���>׃�,RtUN��|�;�J�a\������曶�e*��K�YT-����ŐtU,�uw�nd��ܡV(�N�e�%\Գ�h�;jZ��Q��rǨ��q�[�FA�.N=g��Nœ����X�*�w��2p�Zj�vBʩ��]/k�7p�K�kK��6�S���`�v�j���=��Q88]�k�w`��U)��9�(nv��~��h�:n�RђP�[Z�$b�^
�jmb��1ָ�<1�U�Ys^m�*\LTѽs&�|)p�4��:]�*��7f'{�3���F�0n�6��GH{x�b�e�$mv���i��۝n�,�4{�a�WQ���¾p���brfo:�S�К:D��G��'nC��Kj *���JH�$����&)��"*H���Z�"H�a��i�' ��(2ĩ*����"������*�������*B���&��R�b�)����*�j�JbH,�3&����B�j�"����
����`ư�)�""��fc,"���b�X�3S��Jb(a�E4f�ETj2���5T�%Y-	QY����Q��b�������-fT�������������"����B��*&��#(���*)���3**
��j��*����2��,�"��j$�"�"�((�)����&���2
�)�,Y� U
��V�����w�[O��Ы�9���NG�YAd��N�:��tN�9�*�RGJɅ��퍹^%���v�p�c���]�`����a��^��/�j�uw�kW?[o����2�r\��u����Y��=�*m���Ք{�OwJ��[+{��^���.�7ں�E6D�\�����M%����U��������s�Ն���(����pj�|4u,D*r�t��V�F=�!�����MW�gA���uy��[�f��X�i���`}%F�&}ḷ7kw��ܬZ�\�W�T��bf�դ_LU��g�҇�Q��q	�$Q�("�{9*�n�ʑ[ wvߦ�3��Eod����Br>��oVp�nky.t-EI�~:EwH8�"b���S��Ƽ	�j���y'\t��G�=X�h�[ӊl79�^��5a�W����k5r+�� Wz�>,��5�N�zR�o*�lt8}����#"�c�2_h3���*"i]\��ЊVS�e�/� V��Tu��BR��t���ًmn{4�O�7	a Bt��e���H=�!�o��)�x\��u1���ʏ/ɼ�n�=�s9k�s��r����J�9xh���s`��]�X2\��:7�OS�v5G��5�)��I�X��1�U�=X�֫i�X�����hK�b�抩
�>�wr;d��<��g�T_z��xK#��;�?l�-��Fq�=PnGpB槚Qs\W#�wGEbq;c*#9aב�f�mTRv��;�g��k����\�p���D����Q++n%X�b�o]{��ⱷO{���#W�ho��	3��ۜ�q��<\��� �Z��,O!�,?p?������l��Z�\����5��v��藻*�$ѫ�Dk;��=�u<�P�A��̧ݩ�N�
�/���U��s���YM�!u����ɥ�6���]���U�t�k��&�e��j�T�'po\>:�d4Td՘����@2֍J�S�G��E�m�'�����oI�ra�Z4:��	Kː���v�_$6�(cob�c˓Ko�N`�ʁ����X��C���3|�-<��ޥ~$[0��#F7X5�d�g�i��R�o7"��FS�U�b֝	)`NfTж��\wq�Ӹj뽗��*b��w_}�8�Φ�H��b��S�H4�ї!�o��_J�o��f)���[3��Z=�%>ڲz�v�Y|�C9�����̾��[�!v��@�"��{*>����9W�X=��I�'��-}x..��
�g<�<��g�4�>K�7"��w��wj<��9\���ߠ,�]A�s���5�����-���v��kqKImr:�c��w�����Ppc9���ٳ0z��ޏ>u˄�i�����B�e�Mne�պNk�f9��@bb㝃��z!��٨�;׌{e��C,�c����#
�6[_\��%e���UfVv�i��np�\�j�'�)~�6�w�}/�U?R�_N6u�o*i�8|��M�6�4�7���{b��'v%���b��z�����s�)�B�_��z�����;G�6��I�� >�1�v�gzoԺ�N%�~�u��Һ���D2�
^o�wV���[����5~�7��L�j7��Jh�Ԏ��t��YS�J7�&��x��#�����=���M����03phnTck���f�Ɠ�Ӫ���{��vlJ[q2q�g���^�Ѱ�	����}�f�&O����2�'v�nY��:3��\{AP]�v2����X(�<�y��Z�j9%PU7p9�&�V穢$.��a�Ppo e^cGb�[�|���'&���r���{֒5m ��x'�F���ٕ:�"���f�b���q׎K���J�Z馕�s~y��ĩ���[��v�Z��6ލ�J�����iԍ`=�Ⱦ��w��˅y]F���^�q�JGV?5�5�;]~Lhu$,v@o���ˉ�[Qt��eq��Q]��|ٞ��tnv��9������BD)׈���vt��H��o)���M>��Y��By�ݹ�v�C��)C��F	�MI��N�\1V'����S�̖vej���C����Bt���5�t�G'��y�ޠV:���[N����Tnɘ����3���h}Q}�����-vBa��SQ
h��w�����ٖ�Û�Y�ʂ��Q4��`e}�c-罤��"�N���$�c�����W ����"�ǆ�:�&����C�+W��:�1�5�;n b��s�S^fݮ�v޵���O�c�]������N�۱>i��<I���r���ˑ��룑�ʾ��ޥR��j'u5���e��6��ʂ�^�fyp�f	�W�q�2�o��T3��T�w���3�I�sa�^��Κx���2�'*�澋��0��n�����[T{�h����o����L�\����3������x�ŭ�pV�R��n�-�ے�e0\9յ��(�9��x%�����@�?����������>��V-����Ϻ݌�+�����e��Tڸ���<���;�&EJz�T�V�5����Χ��=K�Kdp���n�1|�/��~!�P��,�Qy2�.G1PȚ����|��}����X�T�D��+�umɾu��K6�lgB��u�L��䕼ՋO7ԭ��髮�VW��67��+�)���6��}��?_{���cўkJ�>�.)�$�s�d�UkR~�u��8I��J�L�8�P����9^*� ��nb,rk;G@;��a�����[��ȗ�Mh��sۗ)���c��RU�wWYe�zc��̧��fh_w0��33�C�jFu;�v��`�7 M��)���2U��ݴO5��ow�~����_Woc��ژ�90����q���8�	#��;{����5���W^Kɑ{7�ex�Jx�g;�c8�3%���w�����xJ�=����}]1;5ӊjHJî�o��<��Yx��%��9����l��^us�_oT[`B8��}���F�٥|�%:���'��9��F8u�E+%���� �r���Ek�g�쾰sj!�پ����fv�W���QK�bś5����ɜ2��ϩ�����\@	q�=XM�]�Q����,�\�����v2�1����^Dl�w�4���8���I�7S/�����v��:��ص�c���`)����z�����]�PnG���o�u�{
'��R���?C�~�oݯa�5鴺��^]�NV}Z�ͧM�Mp���/��������=a��g�
�WQ�E�����k�W�,�ES�wJj�]�ǹu�`���pD�XeC��&b�9b¥hә(��/�ͧS�sk�es��)�kj:�q!��_:�Ρ,| ���V��#�^!���k�t���4i1���׎.��%�8�q�����bZ����C�R
��de�����SQϻЛ}E�6m�2�a�ڴ&+n���Yk�{���߾�&�=�%N�:U��>��w�-���,ܸ��1q*_	��_��#��ɽ2R�rO�����c�47	��;niFT�B�f3}�e�	�;3�Ю����mr�bA�PK�n̦��<<��Y�\,�0�B�Z��&� f�m��Ƿ1GO��[7/��Z9Ra��c����n&+j/�=)q^H��i�|�ݭ���!sJ�f��9B!-�S�6�����:�b�n�o6���Zm���A�s�9��nv:d�~u���M^���v)��|���}�|�˟�o|�� z�#:V��v�9����t�`� 6ź]�WfV3{���N&hGz��飗G�y�f�ΩZ�+ķ/Q�0$�v��6V@�uj�Q�V��5��먐�;�Z����4�t�����f�i+g����o�8\Sc��6H?N�x닳2�Uj3�2��Ŕy�v�
֒��R�#ܐ��҆;T�Q��z8�F"�^1�����`�Ԫá\ɘ��r��2�޹XP����JCe[��P�K�{�6kd�]��35�%�v)^Ul�6�����
sH��i�O<)Νii��\���3�z����L(:�gq�z��N0�
.NI��G��ti��j{��y�!͋Y����c�o��,�
K�ۼ�aqъ��J��F_���&z��?K��N�+�ܩ�~�N]�B_+�F������h=<�
M��%ʒ{��,@��B���,}h�z3�fD�ss�ӈ�XХ�ӝς�岧G,���V螘/8�T���sY��/�&��V��K�]Bjޕ�^�������44_B��]�Y�>ح^Y��9��C���e.;39����!<J�6>�~N����t�4��6ʳ���k���E=vw���YΞ��E��A�ꩈ=+\�c�^LN��� B�b:|��BUYڐ��w�4(�ήh��yQ��V�3� ���{s%9���� �P���DD�J�� �Vrҳ�Qǆs&U��]?v��AZ�dVg����4E[���DifQ��"
�60^MAW���@�����[� E�8���YK���R��[�y�f�*���'
г�Ӝ�݋�K�}���>�P�'<�Tm������qP���·�tl,����Jo��l
c}�S=��:��c!��H�d������0��R��h&�mY�#X�B$P�+�eaWmk2*9Γ� �9���	�k0n!f�C[-��f�|���^&�}Vm!~�j����HX���14]Vr�+O�{Ş��6_t�޽���@WH#��לԮjt��pX6xU�j�ACZ��B����t�άpEjL�qs��vEp
\F� �VF����\�3QΰKS�Nט�9d���},�Y8��;��s�\���}z)��z�X���b9���փ'$��3�a��<��j��t��r�jo�o�>>����1�Y�P(�E�V.g4ȴ�6Mk�9F�5�eR�Ƿo+#����;����zp.;w�4�Q�#no��=��
�������u趧���t�+1�*�#rlW��β�sziG� ���>��Y� g�Ƴ\R*�UX{Qzj�N��f.;<J&]���?��]e_1FC��Mo'|m�C���u7���
&*��c�H8�:*�yL���m�7-������><$�>~ލ l+�n�^�k���� �ϲo��'�W����X�>�����d8.����S�Q���ݽx]CrDd\d�	Q�+QGnG����_u^�{�n����K�f,З-�V��$6cx��p�2��z矂,s�����މ�=�j�/c�/���;�ٽIX�:��8g�|�o��U��	�z�B��P�]n��Ϥ~��0�#��"�ޤ�#[�|A���4X�r�κ����{�0t'I
�����.�C���+^�>7;R6�L}�U��=�8o۝;4'y��U����nX頙|��rZ����%7�9o+�vhg�"5�]���~&���)�cU���n��DF�"*�oROEv��SF���)�ځ�}22N��P|�z�
�5�P�3�]���)-)k�{J�!�F�٘��ک~��R�����t��n+��P������{�O�8�kd��.6x�ı���W:󚎚��X�����d�=��;sN����)j�4�}��b�H���Pڡg��?��8D��X"�V�4=�fS;�3�j��_wp����G�2P�ګaኈ���#L�)b�V�{FL�8���ϔ�0���];Z��2���u�Xߕ�M`D��Kj�����L1ZO�lGdv��h�ف�"��
����8❽7U,ޜH%��a�2,�f��-\YY�o0r�S�U�5:��6�+6�ɭ��tv�9\1�$��{�nm�}ֳg��б\���|4�H�7�H�&����[���|*��q)@����.*O.k��ǕB��u�
�Pt��-`��g�|��+o�ڨ�8���,gm�R��Z��kS�m�F�)c�$���.��7���<�fT#%1C_1��Oq���n���҈�����^o*�����f�i�-��A����C:�n�t�Ղ�دxVBM�[,��-�&�X�����"Uŧ��j�a�y7�t�@*��
7u��Y�#�`� l��T��݃A�م҂V�X۬�}k9�^�01���ŵ��QOF�y�Ajک�y�e^1F�Ec]A�u�����{��0sh�7}Ή�.��(�f���2�,&*�[�ƫ����i�ћ�@��x4��)�{ר�=w��K�����o.J�h�`��5���9�a�z=��u]w%Pl\�4�����;1�:��[�B��c�9+,h�S8[Dp�T��̽��/WS*mD�	��|e`������Ӡ�[���)�ƥC4GyX*�C��]�a���ͧ�����ʹ�z��Zﱴ��7;@�L�|k��U=�w�G&S�n��Լ��\�K�D���	�u,.<T_G�h�}�V,t���i	S�����#Y71&6���%�s��Vp]�Y[����nu��i���ݹ�\��%'u�Q��'�y__-�4�]*�,��2ڽ�P�E���^���7��hm���a@6���pn��61�3\�Ev�Ք���kU�b� SOo�Z�<��֚�ģW�äTe�1�Uo��W�h�ZNf�xRJ]pؾ���.7�
�͙ �W�'�Gq����8P�N���Efn�&Wd�(]�Dc�pAR��ԯ�%%�j��=��4J!'�n�V��Z�W�^�l5l��}N��6(;��"���x-���\;��7�H��9Wj.�ڶ�o��j%G����s(�v�����yiP}��vg̜�'���e�k9DT�5���m+ͮk�KZ�V�j�Z)d1��h�剩#������2�i�4�+7c����:�FyQ*��)�g;@[��v��i.{�n5�n�I�z^�bU5W���=����J�e��J�?E�6R��O��	Rv�q��9��o�ZӠ�v�:E��WI��Ӗ:پ �V�eq�S�\���]��|s�&D�،V>�E#���x ��%�j�YWc]J��ۺ&-#2�W�,	z{�}���{����r�x�L �[�bD��gȣ!ݼ!=HMŊ>�-�,��t���G��R;{y��$�]����1*�j����$ʒ��)��*�,��'"��2����f$(2h0��$)�����)������2�,�s*(�JB�Ƃ��(h��(h�����(K+1�bh�0�����j$�����&�iB�,f*j������*�0ȡ�3��(��
j�*���#�� (�!2�h"h�)0�"&&�
b����i��(��X�i��C�2p �#
��[1ɬ�&ZJ2p����("J(�
(r\�Z)�K2����������̂h��2C#����,�&�&�(2ʲ2��o���<8tn�K�@�#f ���2�8�����xt_W:㷐�v�=��4+]c�d��V��U��Ea}`ѽ�����z��zֻ���r�ܫ|=�h��U����+�_f��*V�m_��$*{1&�󸼰ų�����"Bb��½E�8Pr��q�<��)�c�g]m�;Ѫ� �sJM'�jr;KiV�6�z��γ�Ɨ<(�X�L��X�+��K>}�D���&�L�Я޹�ʔ��UJܒ0�n�n�:�4����3���P;�`�:��^��:Iqy�� j:XH�S��B�n�7�N��j�����1çPW
7�[wm47{EX�R��
��)�JJbo%�M� �9�d 5S��mf�ӽ/8(�;�1�#Nq����7��+���(p�XҸ���'60h�����n�
	7QoC�'���Y�y�F����P�t���RÕ3a�A���5/���	��ۇ�����l�K��x\%0Y�����,��(J�ĪTX�������9w�7Ѵc���+�//!=F�)_]�v�x B��sprH�)��O���+�~� 4�CWc�a�ϰ,*�j���]
�Ӵ�Sx�ah̉���:WVv�����w��#C�� 羼��n&�pFAu�5U�dRP{ۜ�nt��%����l4���y��F�ُ08Lj�z��wC��콘z^��r[�זj�k�K�������F�L��!�'�7���B�V2�H�DI���v�u¶D���ŵ�:享u�.�9��0�+'9NF�.�a2Y�%@�ba�s������7�4t�ܨ�%�:�ۤ#��>q_�^y��լ���^%i�W�Yއ	�a���켤��zD���ݿ�L|�6+]g��\.�g�����x�n;�[��ayC2l����T�{kX/�m�����
�+i�p��B�n��P��(q.�g-ם����{��J��-d��ⷮ+��^��s�346Q<_�c(���f���+1X�۱uڻFj��K̎�q�X�9�1��X��,T[��9���%��2�
�42��+�%'\�������"��	����oV����E�����s���{�*��;[zI�S#�����]i83�,\�V�P��!��+������zl;���M��h�$�_k�k@�K�3mO�N��ŉ��s�d�ƅ*�|i��|5���,ջ�Ǥ&?0MX4 �E�ݻv��|�nđ�)L�W��A�5w��3H�:V(�^M�mY5m���I��B������%u�F�[����D�k���L�]-?�c�Y��59��(�X�܅[`V�c�|���*��2WiRQ*s�����/�9=8��k2�(�f��RM@�P�q�u{�	I(;�44?��0�q��2%�`��a��m`���!�0���m��R����j
�����R� �cwr\Ɩ���o�R�b����t2�?i�g/ѓ�i�B�R*�\n����@���_\ӫeξ1z�_�w]��&����*�_���.pa�B,_��;o<��	�����@{�["�'�z�Ky��VLH�/ǧ��Ȩ6�n0����mx��L�w[�x�kY�r&A�n�S�`6^洪mEH"���#��-����̦gJ�s�y��|�����T>�3���F�V�[z�9oNsp���Mg�H�
"�{c��T��c����F��2��=�@�<�����_.��q�x����u=ʵ�ߓP/u��6���Z�O��l0(kM�w{Q���cQ���/4?s�:j:� ϒvF���Y�g=ΰKS�gG_�
�nb��.��g�,��3�c��P�i��7iPD�!2{��u�'q�'�87&E��I�F4���eT�	������bv�����Y�[��ɿjy{����ú�ROQݝ\_*0���S$(t�>ڜ�ρ%&��Wfܥҡ{Z���s϶�s��4�6�x�*x��*��K�&����t�������;�\�t�)�;�S�	ۍ�������ͳ��6��Х�٧Ѝ6S��>琇��<��u���܂�i~�Xxr�+'p�j�*���Ffs�/
7�_��^�	t���<{}Ԭo=�R�ct��>������.�5 >�e &2y8F��R*q��"0Q.^��y��eNX�p�1V�쎘n��v�~�qF7⳯�+�R�y�F�[W9_�<����yŹ�_J� ��D'<9��QY�tĘR�F_*�^���]���HC&��i2�F�C}}�o���s���'ɚo����p�N��aJ�T���0�i��Eu]�Ǳ��Ꙟ��'ȗ8�\�s�e��4�6�j!-�㋤�"�	u/[/1=W�s�!ή��1��7�������#�cj������v�^Q�brS;.�,ZI���?Mf�;pn��d��H^�s����K2��V��0-�LP׼�9�U�*pD���c�e����+P��o����Wa��>N�N��ˢ۵jqWEFFS����vV*&���̑�2�*��\�.�Q�{�sqz����iR��]�	K������	��˅����:��訴b�Vv�0s8�B��4��7�a:�
�]��V��N�*`I��4�fʗ���˻�ŀ�$����rg���BuP�&�Iҁ�]T|��/�)Ĳ�MX�W�v�ع�Ζg�z��ʩ>|NB� ��)�I�*9ל�,��L����iHvS�\9]�=q�ǳra�͋!d.��^��9>p.3�Q���/ŌD��T��+K�IF�Qz�ꎰ��5d�h�+t�OlL���]jYC��["ut.���&{�M�p�;�۞��>�!���k��jlE�r�?��"b�Dix�ѐ�GI���{�f'�*5����M��dpC/&%)�/_T��`�<��Nz��p�2.^�/�y��KF�����R��qM���%���u���ٷ[�\�5'Y��>Z(�X�vL(�~��u/!ݭ��,�u`=��mL���4�m�U���:�4�x�0\�oD\�q/c��ݎ�,�$�.��r`��.#Mq��P1K��D��+��n�7.X�x.�	LZ��3����v���z �\lW��f��S���JJbn2Z4�R��Od�:Y&���_�p)�0�ј&�T.�1(̽� S�_^(�}mBB��.��S��������)��S�5iI�RYw�G<��'^Ll̔��9I{ӈz�k��Fn��4nS����åJG��*.kPC������Q�d41�A�wZ�WPGl��� �a>�V�Ƭ���Y�/����Qᡆ��i�y;�~�n��Bd���)\�sjb�8z6�7d�J˨q^< ���n���v�t3���W3���Z�s������8�Ҵ(Aٞ��f�I���ʃƼ[W�u`0$-�ʱ��B�'9e��_&؜��'C���{<a�	WUT���p�	9����#��g����ת<��C����S�vH�|9�L`�9�c���A
�uX�9 :$��:��,��몽֐���MWv�dVN79@>��"l�K6J��¯x� ��;fSF���n��~�� ��T5n��S���瞏MZ̎��.r�^����Z�$���)���v�b�F�)�D򺐻"���j�Y��\-�p�g��7�
8��X�n�B��yJ���FF�w 
���JUo���j���c>�V�dǎ����p�%�
�%��}�tsj��q�@޿*��I�dsyz'���k�*l��:�E�vNG�A�\��t��{�*�u���!�sܖ��3�#ұu��P]l�}R��N��Q����iU�)4s�B��Y6'2��R��Af4ѫp-��8ؠ�K�)n��E�%�Z{h'�!�s9�w���z0;���������\��tD�qWP�!�ıl�2�8�Qb��f��s�hn���*����(�	øUwI.�������u�Po���E�
�bJ��c��P�kd�0���;jis�fr��c��O�G�!�ruFL;�P2-s�%=*l1���$e'˪]T��l�OA�vzI_T�3�N��>�L�wi��XO��P׻�L�ۏ������Ϳh֣� .�b6�h�r���u
�O+�tg�̈́�.�p��1A��Yq]��y�/ ��.8�UØ��ߋ�1�<J�����mu^���0M��1\��N&.��ևVA����F��ؒ�O;+��k0V*��(P��&��Ge�7	�h�u� 
].#�Q<�:8�T��.��Js_H%q��또{
�Jo[��UO[*�����EN��=Pmt߰��]F�6#D�ڐ�ו{s_�NtpIv0�>�DHVy%I}e/ �F�� ³�P|}���Q��Ȩ�:OX>��8��V-�fe�Y�I#�OV�[)g&gswb�O��v�����Y�x �{6ۢc�afJBS��Ǫ_-���[��~����:�nE�7v��V�;�ɾ�do/�p�4��ѩ�����Rx�U7��vcsX��[��\c�����O��<�F��y�\�G�4�[�D;9�C̖�ݚ��Yy��}��ñO7b�5!�;0�{8��'�?��X��8Q��{YW��0D"��5�l�l�w��v��˾�� 3��5�r5�5��8fv���?c8��L�L$�{|}Faۦ �>�q��$u�X}C���� *��s���rI�/��#)��{��
��c"{OIB������Y�V���3~FQ�憄�i�]U�x�g!i�΀���j�]���qz\�L6�������/K�1q�+\�3V�+Y�=Iө������(�u/��ڿ0�������ҟ>���@{g�������cM��i���b�\sĶ�ځ����u��]C��5�0������ܧ����Wu���ɗ�c�٢>�in@���by�	1����U�|R��=@nq�FVu��	����VL��Rݞ���;K!"A�#8mRsB�H�d�2�J�����@���.��l���
<q�P��J|�	f��\��.u�w9��Ѐ�\��6%��X�}W�x�uF��.x�ժ�xM*
V�0U���
U=�v��F7�۫v��/s�r ��v�ouf|ʷMb3:�K[X6��e��`���y,nm��iO)d�V:h�AÁ<��?T5���SJo+�k�T������p�]x�>�M�]��#�9�F�P�W����,6�x�peq����G�A�K�Vw�*�
�,�ݝ��̺퇵�$�\�Ӌ�?>�E�0�:���
/i��Ln'ئ2��Gyl�Ga�n�-���E!�^4Mz	���':�p#���Y�0
�/���t���)����0,pm�W[}�$�B�Y�F����(s����'UZ'",W�s��1Y9��'r�GՃq7�ޛ+��.�B[H����g�Pb3��.�p���^sQ�PY��m瘕{~	�΍j]��>�L4}�c���,H`��6���<��^�oy�}�p��cI��OVu*�o�4��O��#��>��Ȳ_���U1�&X_l���,��P��Fs���o���8�<��C�ݣ&����`�di�x�f�����>������>��6�Ѥ/&�Q�N2���qa��1<�$)�}�.��QxMd�,�,o5��e�1�c��£C�F��Rz�V�u�^���@㢁�0���OY\���vr�lΛ���7sm47���*����Mj�J3:�p��٦��\�7�W_P|�#�z�nWj�f��35"��Fs�}�g����0�c5ÎH������:���{�z���g�a�ku���odr1�3��.xAGD���j���A�V�Q��$��k�ѭ��@��:��L���SA�m�SJ�c���/��<0\�y��
����9o�Ԗ�G\f�"�w�Fr��T���a#~�u�p9�M�F���Z����{��sd�>�خ>傈��ow^֤��X�����M'�7X�v#�g�[�Q<Y��h��T��}>��Qᡋ�s����ls�����N�:8��&D��*4E���ͭ� �����RÑS6�4�]Q�]w���BK�W��$��e3�]1AxN��'0Y�y&Vr��ڸ�66`�[X8��MB��lb��6�[������&���ݱ�!W��-͜�:����5+z���w˲�'ۧvˢ�\`Q79Ƃ	��:�hF���];W��b����{�S8�ϫyz�)gi��>۪�w0DŔ�d7��w�20��2��rV��c[����+U%qA���P7L�1���/@�Y5���ATcd{]3Ԯޙ�>tI>eu�X{/m,�K���@��P���m���fg!�곕Û��G�t)�hB����ld�k\O��y�ZpX��S�|/��^��il2gW,ڽ:uJ��,�@����Ra�\�q�vn"�����	L;�l;�D�0�I���Vރ��vR�D��RN���=�lM���S�
ai22����i����Y�]L=麱��ɉa��q�KًI���^Ӱ&f� ���W��[���b��O���+]�*��b��Y��Rb�(Ft������V��},#x̽��X�����J9d��]���r���n��:��L�\��sr�m��� ��\��7�Oq3��uCfQ��V�E{}�Ŷ�q�L�7��9�f@A���h:�Cm����b
��Er��9��IU/�c��<��R�*�9w���P�A

�yp�P��3?n�?{x��y�Bu�3+/7���E�Zmu,\Cq���3Z���,�Ms�>"U��	Z��r���tnȮ��MSǶ��[���A0Dī/`K>��D9�c��F���4���Q� ]���PKM�d���$�P���F��)��1��q�`op�*uݛD��.j1�M ol�H��os�����X/����W�ٿQ��02��x\(��j[�X�u^qt��1���1� y��Qb����Ȧ%qˋt��u�H��A7����
噀�C�yS��>=f��Ӣ4;ah���7�vR뵽M-#!ỳ��7hB�|k��[�J���I�-��s�����ڳ|�]��-�˩���1�÷���:�(�m����u����V�e��Q��,��ʸ�o5�# W<�<;mwK}�Jd���H�(^�WQ:1oM�����t0���'P��XF������N��3��5���!6�TOs�����M�h��$�\�>ެ�N�I�z,�3OM냱8�8�"��h�WB�5t0X��Y�� 4)��m��F��7n����v	uV��54MCDL�o�]�%E�
��M.��ev�W��*r`v�����""�oqJ/Ď�fUhuܡ�'(!�l �p ��
I�B,�.oY�En�@k.֗���8��i�:2�	�D�͕���@��]��������h�JWV��4]�O��9|x�	��{u�����M���X�W�X�7m�[Y/j���g��Qe�� ��re�%��t�.��������ʭC��t!<�o���nd-���!`�l���J��}�3�=���̧�ԙ�L�K}t�E5�g`������z"���Y��[-��D���0ܻ���\�yآ�,�	#��'v���|����U���kQ�wW�  @�#�<"��),�ʃ"�(��� ���)��&��,�*��"
�
����r�

hh)*��g1ɉ�����**����,2r30rrr+ Ȧ���"�"�i�������""(j�2�����"�(
��$Ȣ��J(�ɳ ����j�2��*��'
���30ɡ������h��)
(���i*����[1J0�)�0�+,!Ȧ�#,"�3,��2r2��&�3$�,�3�J"�3��3�K0)*��')��#$�h0�2̬iɠ2l���0�C&�2ɠ2L�������0s0�&���̱l2�	0���J�r0��12�!���(rJp�pA	#�`�#�{�P���r֥	�/S�>�ͨ�(c�Vu5}W�(���f��$�/p��Z�m��D��ZS_K�/`��Sc�-��$�����m���5{MO�睈�9u�z<fM{Ux��o�MZ�	�̡�OJs<�i�1}��,Tr���5<*�}�8Ӏ�V^��!�f���O�T�c}ֶ.�yOH�� ��51����%���:����2�Wmj �����/,2vG|�@�������3��Q�^��u�gY�2��L`�q�8�}��s��Os�jk,�>�ֶ���ei��cYd��1Bb+�=3�N����d�snm���wR�P�}�1h~,k9�CK��+�ѕ�y�q�u��VX���x.#��9̋86�����+�퓏�]p܀摛�:�,M#�%7��Z�'��ƃ�s!��8�$�w�k��4���
�k�"X[Q�e�걙�}R"�"zҤ$YQ[�����7S�ukغ\�� 'p���َ�I49�(yTgC��g7q_���_^�_�'����=��i�1��d�g�ٍ��}��@�)x�B�5
�po�R�ҭx6T���8�4Nt�L��iT"�5P­V���N�ۆx�+*LLlj�n�"�%iZ�Ν�M��&m�2��#m\�uf���`B��X�!�컍#�o��[T*�qEJ.�Io,�{��H˗���fT���pT��=憄�^�y��vIԚ �lz��{Y��n���d�Zn�t.�H�	o$�#���Y*Q<�qE�:k��6��X����{U� Oj�`�^�^�>��e��_S�g!� Fi�U)����j([�{�f�:x/츅��c�w�{�;��lf0t�׻��:W�\��FI�Mv��}8���9:\#@��e�L�����m}q�0�o!�e�_z��=���E>ͷ����0�B�U���`��t{ʦ��$p؃o���L<5����@ �:̛�)�^�A}w�=�\n�&x�3ڪ c\���]M�j�����/
���i���ocŞ�<y>�	��}E���č��U
�`>��
����k�&s���8ftv vx;�/���t����fB)Y��bhsu2�ۂ�����P��U�B�]h2v��V��;B����-�d����*�~�eeޱ�P#��z�m��,�7�3Qi��fI��Lq��ګ�&��l��j��v����K^X��� 8��]�,�~�>ʀr�D� ��m���Z�
���f��î�7;��$����{6��uhn:��h�q���7�_�t5���G��<^NX�y���!����i�Ц�S�nt�G�#�Z��e>���lgMaep�,eؕ��]$�����gycdy���~���*��H�l����4o��qK��Dtk����M��f�v�c%x]�6��ըSj{��e�Ԃ�젵���E��#��I����a���l�6�E��X��Z�Qt�s�!�΋�a��X�<XK���D�;E(�����υ��1r������n�K[b�o=�\��h��.(��z̳��e�/'����x�E�t�$��]�D#��{�DKӻ�3r]��ʖ�U�#Q/�U*���ܐ�w��(/�jy��3;:�˧cK��Tl�j�?z=�a��@oB���}�_�݆��R��E��w�^��V��#�*�gBj��O`�p�.��B],�=���B�a� n���4��S,`s:���)��R]�4�+Q�[n�
L�8�G��гrgը_Z�5L��� y�Z%oO1�r��$;��ذ,[���8�A�THb�����g��Jp������2��O@��2�Q٦�ϓ>����hm#k�.ྪ�3Ҕ� 9'�u�5�T%�W�a����zp���0F^�gE�s�}f��^L�Py5�Z�%�!���LZ�\��w
�]�3ݸ����V���-�+��+���Q�K��%c�Վ6:7.�u���WO��7��ys�wr�,J۸��ã������#s��v�<,Sd���c�����N����q��'<���:@�H�|*@P���F��E{t���M�Z���I-��+�I��)��V��`�<��r�xc���=+U+4�C�?�o�aP��,���^=ؖp쳆E�[FL*>=��m�r4朥��/z��%��fR��7�U���KD���T�|���ʃ��׊�������V(�z��tϬ���Tea}�D��к���yq=�Ɠ��3�mԇ�����c{��s�:�d3�)�\`k���l륕�����N6��Lc�"����)��*h1���q��C�����:ݮy��/L�5��V�]Ot�8^M��?B�iv_���t_W37�,6K���θ\Bn�7ϥ8������{`^.��Չ)M�`�c.�B�&�%6 ��ue%16ZR�_RX��V<�gz�eڌ��%�ʒy?>��|tXh��i}�C]u��hmqF�r�3��}3_:�z`��R�p��Z6�7d�Jງ��"�c����4e<F�U��Y~�usv��Mv�}� ������k��kN�z.[u@�X��S�{�u3���8�EE`e�m��x�d�Tt�Ǯ+�\s��;s�p<*8j5}�3��S]��kt7U���(T�
Fsej��f�r�fd��-�.��F�Pp3K�Q���lP�;S�����&]����������>��t���7�wD]
�V=�����,*��
;�3��Bt@nF8�lWhrD*K{��f&����K�@��d�c�윃	��L��f��;@:$�,,���ҺkY�V�H�k��#�_/R���a·>۪�f!t~˙w-��Lo1P�I�z�������&��sv5�I!�>!����,�N-Gr5�}=FG3 ���2�м��4��|�,�ȹ>�����t]n�8hq���rh��
���A�����s>x����P�/�M�i��;|�S�&Qz���wF}Ҁ3	<�5���δ��#W��z�A
�L�6�#3�C�s�B>��%�]1}3�n9H�ԏ��n��:�3^�<&T�
���n��1�N%���D۟(�a���}RƲ���i��eo,����\b����lobF�j��X�r5�B�a�:�Q�Q�x+,uƷx2C�]'{ �U'Rv�¦��\�y�Rׁ֩װ�J�1�Q�`1�,���f�zr`W�q�#��K���*������i�A��������zt7��$�C3�5�p�y·���l�}mM�)vQ�E�Y��6:�#V��;:a��+�z��7{����4u����r�u⴮���]8����\ޔ��*N�wr9H��:��wݷ��-���Į,T[t�h�r��j3�:�tdS��f��mH��E�3.��qY;��ƻ�5����J�n*�)�r%�9�(yTc�8��T�l�^��Vj�[b��4��/E�b����FN���͗�hd4'�CC���U��2�<~�M]����+��3��TX-Ma��t,+U�m�%�� Gj�Q����zk�۞�7��)�� 
]=��-V�=,E����a?(ܼB�v+��k�v�=�ɪ�����c(�PZF@s���{�@�Cc�\�L]�zY�:
:����ܰ����Xϸ�F[���GX����e	'
�0)������df�)5��&���t�p�]B��'5���U���){h*cC3��׬�Ŏ����K�r�\�xhs�(�dԚ�(��2����T��X�1�"�"��ʴ6����\p�{{�ڎ�=ʷ���ҍ;�{{&ӻ�T���\U��(����a�}0/�ѳ��{S���/�h�S��b�����N��] �oWM��#aR�u�f��g-�����f�]*Nrօt_b��FX�G+⡾�{}7KYɬ"���.s��_���Dy�]�C���6�P�*��ގ�}��˥�e�^�(�1^I6�����s�Q��_z���f�!����e]B ;9��RjKPS ksbcӵ���3ҹ>Uf�d����+�4$��Z�y�W*�3��xH�3��NH��+(5��>jo&�A��xP��E��ւ�\^�s��i�~XJ�����bf����U��Uny=�6�kqJC��S��oV�p�O�o��]��ziJ}�q��@{�?���%u�Z��_H��V�EN���3Q
e"�UX}�t�!^��dv�:�1Aq��p=�4��^JdBr��cG���(o8��TbtF9bGK	\V9���l���5!�ՙ������O��8��b����sY��5���2�b��_��fo'��}H8ju��*�j�Kb���WY;tqu&���^��i�
�^ߏs��Hv�o���f%`���b���A��lmu��YXV���މ�3	�2������H�e�G��ӿtc> ���*���E����ot�|�	���V1l-�[���ބ�mO��s�V2`9�P��-��кt��n��w��N��]�W��Z���b+t.���-�7�Lɭj���m���)
��f,Vf�޻��^0� �|^�6�=�s��gs�������c�:nU�S�p�ɖ1�W�;���۶c<�EK6�Hld�����,F�LH�8���p:Gz���v�,�u4V��T7v��u4�#q2��sr[���m]�����2�Um{�����;y��u�@ ��^.pb�T@_+���萔�⨋�����{�ܷs�-=饩�\\�u�6�(�����T��	���s�2m�{�E�$��L�7�si��B{�ֺ�T#X\�;&y����^�a���IР9>b�	#���;R睆*��>�.�H��#z�Gk�3Cm�<4Sl��թ:������H^�=g��.�dN�t@��g�y&N�gǡ�V��m���*���j^�H n j�.��?x����W��,�?1�3~3�X��Y�Y��WؐC4Պ*��L(1��4�#9t\����og��)�c����`����;\�t�k��������Ql�FL39M�V��X�\z��ݽ�bcQ�y�S,1eM7w��ۮ���wb�s�r�c6�]~�g ����i�,���Ǩ�"���^VS���n=gD�M:�`�bԽ-�v�1�o�nD�]d�QIn�S��s�r�-	�q������{�m��
��īeJ��
�id\+������t�-;:D�I<Ιݹ�wX� ��pKU->�S��]��Q��{s3~R�f��y�u��T��9om��j�N=��<�P��0��=�Ǯ�C��tlW	J!ܠ�5T�J�gweb���ͼe�ΑILq%%�����a�N��ʒkȺ`GgDI>��_wJmW��J�]�vu�:�*�#Jnl`��ڎ~Z6�+I��s
�O2E�m=93a�x��Ù���:��͍�A�Ub�6X���v���.�O���C�0��<jj�87�b�@剾���emiqPl%yV>��e!z{nn�+(����c�nP�uAo��sʅq���.����Y=cQ�ón*�]s�Ȋ [S�4>��`�]��&<%�6Uc,��L�{]CMu�L�����P����zM�b��i�{H2`����n	P��8bU�&=�]��a}L(!5�v�䲹[���X"F׃�Ɓ�86*�Q�s��r�PX/q����ǮR^��H�O�̠��4:/;��9X�/�h{l��8ӂ�%ayyHn�x ���t�Hr��Edףi�M:��c�1Zx7j�DLYC��R���s�9�3X�ݨQ�mRT�Z�#o�R��Q�{���g�H2�㸺Z�]�M{3�AB;v�S-;�������*{�7������V��c�"�����@[���9�].3�T�N��[��v�W���T�
N���6�n#�i��#V+v~��|���ewP1T���z�~m��T�Q��V봺��'��o��^hx�tsyz'���tL���ɍf�9�ET5:�.�Q�IVN\�@>��
���q�,k,�6�H�W*zf4��TS���y�,��ˬ4n��9p����l䦼(ivz���h��<�+J�¢���>�����u��w�}<Zpud�~W�4��S����;rUQ���c�W5�[4����I�Cq�"�[t�h�K�$ׂڌ���걜�����t�Ɵjܰ�܍8@qک��0���:9d���1��ʒc���\nC��gN^�mۺgg�����4�w8���c��V�#7:�f8&W��3�	�U��B�9�P7A̬2j���h�ݡ�j�aT��6S=r�D�V.#L4r���i��]g�#~z'Iw��ZJ�n�;vEi T�Q�@_V��B|1gj@ڶ���K�0O��
�V�B�d�R1�a��}N�	�5�ͻ�ƽ�V��պ���*V��[eQ�Vj:�˚['�>smA;|���1��u��C ȵh�1h������T������5��%�:���i8"�>�g�8�[�;�íM����q�����㋵��߻eeo=�}&�N�kUsFg!�\�w%�3�g}�&�:�E*�uˈ�\�s;���j�
3(����8'�,��Jm>�i�0�yM�w�.�z8��mRJaM��fp�$�0�[;�U��!7�ō��0�-j5}1\��+7%�Cq
2*:�mc�*�É3�a��Θ'pf�oyY���@5�|+�U����`��c��.�W^L����x @7wƈ��,}�u��C��zAk�ž�y��OL�w��iZ���A�:�Fv[bO����^�Ĺ� "M�&���-.�!�y��.�.��pX�P� ��&�W�C5�h�A�Z�t�L�T�=�b����Mne6�.*��y:R\�AY����}��S�`ʱp�Ϡ�m�vw���L,���/�s�m&�0<t��@S/8i�'�ל(I�1����Ɋ����y�J��|���k�{��e�#^���N����}�ޞ�����M�N�ǚ���C�G'��9�ux~��k��J��Kŵl�s(,��y��M�sx� ��-��9����錨0劗:����J��!:�w�`g�4CpdڻTs	Ww6�ʝ��֒+ T�Vv����Z��ƟCF�JІ��C�<E��,<�+�r��k��u[�*�*�|����>���@�Á��!�]�syn��ZG^��(L�j�l�4B�&��'�8�i�6�C�\nV�C��hr�7�v��j-��R��7�%�\��]]����]�R[:,�kOXӝu�k��H#Y}׸j�ؐ�ăE�������+���z� 귽,�=������,�*��EL#��{l��\�$_m�D�����d��cq�@����w����/5t��=��ƍ`0�{��p��!�.�^αݥ(gI\C}��h�Z�;0nAZ5n���-]�ZOxQ	Fp��;�!�WZ���t5V��d�bbuj���=�)4�.�zm �	U��Jw�vp�����Y���!u�n�S���
����vY�R�W*��Y��,��_!��7B�^l�-(�.���tė)��nlXqr�[�JJZ�Z��$-s:��4�e�3>�Ү�G]7-L7��X/�oR��sf������uBX1�X�i��Ƹbu���n�>�3hvYη�䴁䍡yL�Y��>�7z�n�^Jj����+�)���� ���Ŗ'>�޽��P�B}�y;U�h��:�؝k�J!�X�M���Ҍ�jӻ�D"creֽRe�Vu5��mu�Ķ�����d�\L�/=�2��7�Hz�lqu
��.V����]���4�?KFf#YY�e�A�da4�S@�a��KfN�K�fa��a�����eX�fFQ�T�SA��dACT�4ДPe�IC��QI�乘DENfQ�fd�e9d��S��6`�%�T�U99Q8TE%�M��da$A�X�YY9���4�&FY��fY�Udaf,VY����Y%TđNa�YRSUTR�XfeaRUQ�dDd�YY����IEfafefdVA�	�`&AUf&AE.E��Y&EI��EXM9E�FY�ѐ�Qd�fA��FE9��T��Y�1EY4�e��fd�����LS��XYfcYe�PffY-.FFVb��e��dPd�Yd�E�a9�VM�&Y&AYe�����bQ�FT&UFa�8Pf`�QEVc�CFICFS7V��po'<\y��R�}��fܫ�ܐs��+dsE�.+h�A��Kz���'Y{;9�v�)�s��!��h�W}�7+�UV[: <V}(��Aiγ�j���������ӻƍw ��jxk��:k�y��Y���3�s�R�o�(���"E@�+Ǫ��$F4��w�kg{���횃t˿:�@�*B1Э�/�S��̖�����ꑱ&\�{oF�;�rA�e:�T�����T��`dj��r.�g:�R�Ж�LH���s5���Yכ���Q�c�,Z)�������OBM��ƪ9J���R��Q����{6bD1}ػ3n�OCK8���q�"^��h�9n:�D��C���bBd�y�YO*����s�m����W��(�����U�`�=I�nz��]?�=�5Pg1F�<��H�U��@u��%�M*�e'ׂ9V�V"���W8�����4������y��w��c'��_�m9:���l�^�ǽ9Ň��Fz���,:#��F�U�&�u�9諐q.U*��g��#�f )� W��F��-T�{��B��}���$�x.1�n �w�;aOt�r]����ip�ؚ+���X�a9��x˛؃��]T{0iSSL�_Sù�w�]�}+a�\�/jC�A]��⽧
�� �6dr�]���gx��'�*�/�̳'˻&^)Պ�g!9��{/(�:4��لJ
ۖ�al:�Ž��u�*Pz�	\{j���l�t���Uc��)�6v�Qn��#E�)�(m4�1l�so���A^��U\���v{�¸�N�^9l��O�5���x�D��H+o����ٓu���@�U`�����WV= ���/��^_�d�k}r����O7դi.:���,�u��d��`��oD��0���/��>Z`	Gv.l=��i�^ҽj�h}O�b�b�G�<�yd���*۶c<�EK6�L������{�v���4�%�t�ɋՅ�k7�&�l`�� ����.M3�L��NnKy�mU�fp>�k�)e�KsNP�."��:������`���$1P�T1p�(:���R��fv��*���w7��~��֚�}���ڔ�&ء��*=UY�FV�7yu=�/y��î�A?���(�Z=9���i���c/(Eڑ���ɡ��At�!vl�O�U�ˎp�=^�g�tX"��h{o�S<B��:���K�4t���]O"krѬ�<N�4�ڛv��s1��ߺ�����am���U�a��U�Τ��7��������=�,���n�l,�Y��$75�j�q��+��v���/9�9�.�ŵ:����1k�J��T�b�[ka;�ʘE��gj֓ �K1F=���č��Gi��}V]��h����&{E��?�+�<��o���4�G���n�gG$,8S1�����
m;��3H>�,��M��B��on�YQ����b:�R�ɷ\�(\)�e�{��[��mƸs�5�x9�x��nr[��C����/�<+M���]�
�Q癿)��c7ͻ�q��C��ۮv-+�����:\>'�֥�gϝ>0S��]�����
�U���)a�]O���ќ�w�Qާywݡ�]M�lH4�<�2���\'�!ܠ�5M��g��!y\z�aR�Ƨۊ�E��:��a�p��p�7�y��>~|5o���������Shh�Vq��=p��P>i�ؽ�gm/}O'�b�������v֫��M��\B+��"�{i��m)7�Xо��7\��\�7��hh�n�X�X�:�t-v�;3�S�y&W*c;_�;ƗB|�N������]��u=�W�j�����>�^mWI��^o W]���k
	/�NV�m�tHh�f���Si���P��K]�9S�s���-��Ź/)v�X�b��������Ne<�[�)�������ۄ�+\oF�v�n�I�fq*p�޾ƪq��ɯ�',�
�&gK��͚i�EU�{������u����'SD	��u��\QS�g��mN@��6c ��	��L�%^�rOC�WYm=Ϻqmaq��V�6k�΢���0R��0��� 9�eA�X����)�˖է������`��$Z'UVF��U!��"F׃�ƅκ�~��Gs]pk%A*�t'=��Sp_]�*�!��tt�g1Pkڝ�0��ꫩ� ��M�����v�o�,��v�N�9uv�+�[��a��g�9�I�Q��%-�q���`�0��1~��ǻ�=���$�F��������ε^&m�=V�"5���GT�&=��v�ǖ���`���<��i	���F���ߍ���*��9���Z��/>���u����	�.ym۝q]�fV��k�,J�sH�����ų��
]X������?��³}&�4�n���S�y�C0�o��~��]�\^� 5\7=�#7N���:����_#VXQj0	���d��s��j�d��Uq�Ř]M��}H9������}]�g�&^W�Q,�U�I�]Ǯ��Mسn��h���w�O+�_N�{������s����entN�\��0x*�F��)گxk���E��B�h��p�D&���"�=���|�同��{+��R�Wu2��ԕ���Y��a��2��t)d�E���9��͙��.��5��+�Fb�xus�+ר�ޟM�"SҧG(N�7�c��9RMu
�q��%{r�l�$ϻ�ӎ�3����1^�1B�Ԥf�'Ql�ʂ�mhO��B�&&V��:����Ia��mQ��FW~�l�=�r.{�L4r�'B�p���p�
F7�7CSf�m>}�[[Dd���@��|��cgWNQ�M��Z"��E2��䰭�g��j>�Kn��4�H��"|(-"�pmA��q�U��@c3X�P�W;���t�8b�]�;Ϙ�[,d:�媺���u�e���p�7Pm�*���^p�oc@�q���L�=����C�浘9�y<����h��1��^؇o�#r�iY�D�EM�ꉍ�G���i[�u�7���x˲�ʣ��R��X�?��X�6%����tԇӎ�̗u�5�����t���v�$n��O�~ ����dV��{��wʯ�yc�3)����Y*E�^)`�\G:�T���ne�Mwu2�����e:7�1�ey ���@>=��yyv���&	Q��݇ډ�.�e�R�\��fW�q����,l���w�b��3��r�GZ++=�w�x(�6-�ݣWU�|v��_1�e^�;n�}ť�����;���[D��q�f��7����\�����j��ǻ��3��I��.[�!�w_�Unz��]5�k��g1X�Z�;�e{�#ܸgTap�Э*o80w��B}�U����ϸ���S��"��+K���q�MR�G�����S��!�	�%�S�#���)u�;�O�i�W��+�'��Ʌo��}im��@�~��0� dq�g�H��Ua�:b���l��0�.1�t��V�Zv	޻o�7�diY/�S�Ԫ
�N��r����*�r8S�.l�<������(
��Y�H�v�/,#�L`�1n��*"�aH�Y�k؝X�c����G��A�1��r�vb�����]\���V��)è`���4�!�`��"_��n��=�=�!ʙ�i�e�L�-�{jGe�~i�MC[w�"I�Y�z$��t��/�g�M�)�A������&9+�#n�Jw�'�,�2И}@��kr���ni�R0/(�@���cۡz��l�[�M)���'U�A.���-���\��.�ZEKl��ѹ�V�}k���fe�s��{��g��@|2C �~՗��;*��j�;4��}N��>#)Y:7L�
�����J�Qc.�K����sWD�r%rh�P:�zy�>ޠ��
��Q���
Y*�Nq��p,WjГ�kv�v�(S
3v:#7��ܸ�ݠ�'��]R�,<(��v�T_�wR�D��US-n���Q�:�\yR�*��/Ǧ±�\U��ٿUΆ# Bۺ�4!2]	@	�b�]�@YĵM
#�X�5�q$?-�)��)Q��
%V�9���i32�	�v�ok�C{b�����/sV��p�3�
YbH{����Dds���"�pȞ.'Uc=��cvf��n�X7�_8�w}������4������q�z���~�n�5��x��^��F�GA|��D��%�V/�3+\�sh���)�����m���#F��c(XY|�s� �>d[>��7}���L	�\X�3�ڙ�6�C���`����9�ݙ��ֻ�;��-�`�@�~�"i�
�tn�P7غ��s�f��\4܆��\31p��m��cy��݃��׺_�x`��ZS�O��N�騌4�r�����)a�N��f��o�7=K�gc�5�N�b�M�����j��@��r�6+���PQ��T�z�d���<�4X�	2�m���v��Tz��w1A�F�2ʲX5�˸��e�����a#�? M�-e�J���W˧��)u�2;bUoP��\���Ƌ�J�lm�yn�W����u�#E�u��	q��#%�ҕkLBH��]�w��{S���bZ���K�A烘�Od�:y�$�� �O3� T���S>I��͍���d$�.���L��
�|�76y9�=��F�ei0P]C�<�Q����)��y�[�s<0�˟"]u0�W�\�g�k8����b|5�w���<�#P�R{U,�Ok�5S�������5u�<���o�����ܕ�����ba�
ﮂ�T�t�3�)�j�sg��!G�0]��Z.����;e9K�}��'�K���XTO�9q�0�O�VY,_iCֶZ�J�ɕe�W6���2Awe25�	�ź��-X�����-�u�|����y�س�����+�� \�
�ndc&�V̪���:^��Y�8��z�qP�i��=��9�6�z�c(=��&}����*{S��6�Uu!��u^���}�h1�=����Y�q��+�ߣf��|��s AE�RO 
��Z�~�l��\�-ܭ�����8_.�uѶ��bÈ�ن�MJ2��9]é4���^����4����x��2}p#$��\.�Ӛ��+�����qvdy���z�Hm:�V������jqZ��d��>�����4bE.���������ٛ��-[v�Lb�y�W�^R	����P�S[��3�:K�����m���B��=H�ɼ�]���)z�x%�Uef��6�����*�sP��_e��,6r�hm��meG:śܦ�Gmf��n��jfM�*���C(��K8װ�i�:�Q�]�֡v*|EUd�{nmB�:�u�S��aqў�{[%d���sH���u�2*��*��������X����A*�
k�SP�%7*l=��P�n��.P�_g����(�K���JttSǻ˽6�	�7_T��<�iR!�=�S����Y1éʒhs�P2xYt��]��-Jz�6ed�H�H��S�{�Ǻ��N���͗�hcBx�OL]=9�k���#Cw5����åa�3�3���*%��za���J֪��,	s[���:�����Rݜ���9X@7
@���L2���:�dK���m{�uxT�:�F�M*r������P��ˊ�uu�9�t B�@KD��c���εu��"�Nͦ��b೔s���(���Tq���bg���}�K6���:(� �VF�=UpK�����3�z5xڕx;1@m4aX��D�<}��{2�y\W`S���5S�T|�;�u���<�k�Fލ<]*�S�m���BRtP��u�y��5�;Byk�Y���Ι�ǋo3Pan�X|�����;R���}�X6ۖo9r�}�MY�y�k3��Y/>/L�ry��(:�,'e�J�9��~�浘9
��U5%��1C��Dw,�rU��I3ڲE�Hrc�С�e�)�n�I�F�d�)`j���C.�9ֺ��C\S���ȸ�Q���[�QJ��
���7��pJ��5����u�m�R�, u:;�y��U�{�t�X1@�=�&k�`�� ���d*���vcgc*�����ip�����ER�w��>����s
�|�Q�瀢��"o�K;^^���Yw�2�u�"M�ruR画ZHfU�Vn�p%��>Ҹ��pWx�(g�Z7ؐSB�-r�������=y�츊X��%5<(�A�:�q;��3a�a��d���N�g�-:#���7!��S-���#�[�]�r����E�U�	\m00�@����]*�>r� �-����d��T�+�S+�e����&/�U�Mb2*]�TF'@W��k����U�G
t��5��W��g-�\j����&�9ue}��=��f����vz�Ή�fn2|��D��n�ei���:��Z�Q۝��1K�j����Ԧ�ٴbуev�
(���@7�]r���>�5e�U���)J��7=�}Z�՚�Ћ(PW�dPlV��}f�&p{�IX�h���^�>B�EP��[�>�PP�-PH|�V�RU�l��qr��Ls�*豻<��9��b��a��W5�-d3E� �_C��%�����@uj��<��Iٲ�I��:k�<iܰMD��fL�:$ѥ�����%넾�t�j����kŁJ��n�n\�0N�՜^�eJd���� ]"��g��Q�$7h?��i[���]�o)�d!r<�nZ�k��֒��]t����s��(fJ���+||��u�e��!&�8#�=�P]���62"
��WV*z�L}�Y�NU2é;���>Z��ҸO��:�^ok���E�����u��4�Lβ.��}��b0�������s���V�.<��(�ywh#{%˥��
�����e�Ȣz�3��때tê�m���V���a�q�v�tb_�A�B���ң;�Y$�]{��6�B.�ՅSɱ�3"�W�q�*3�%�������k�Д�K�����#���t�Ah$u����,qd�;����$V����
�v�{5e����1�X�V�4�u��k�Ǜ����j;T�㶠����m��L���ZK4���q��-�}��T���(8� �[7u��	s8T��V����ttcPAd��]�v�|�^��x��'iSuLiu���v�1��<�ç+n̩B��;х���Of�B�\��Z�nNcm.���n��퐵��y�Y�����^3e��VV�lP�Z%e�\%3N��i���T�ǫ�fW>��Fv�γ��jMm�ԙ�{��o��kK� ���XAO�m��E:Ʊ���[t��#	H�M�e��C���j���y�u@@b��F]~�ˬ�x~o�/!t�0E���w3��eSQ|�gw1��'��Nb��<�C��x�s���ز'ce��XMH��S�֛���9�	/r�w�g�T+�/O�m��ӝ1<\L+��k.b4S�C�͜0ʊ­���_�z����x8�mj�!��>6��6%�ǝuʑ=���ɁȐ6��]������[�_f�e�B��DKTX����]��nT�Z�J�37���5>�
[�\֮|��YnF��)����Z
�5(ᶒ㗔����dl��`�u���[�þ��q`*��zWv)R*�J�b�6v�X���v.�2��9��V��ģ�3�V�ҐYw8Ӄ%u��̾�}O;@V0kT	ܡ��gN'e��(e��Y��Ho'�P�!c�wb�zb��Yx�d;ӝY���a�"�lY[b7p��Jܷը��'3ͺPA�3����� ��3ݹu�sV��=���(����K��;�6\�/��t�~Ed�Y9e�fe�dd�A�YFfQXd9�5�e�FY��d�YXd�NFE�S��4XNDF�AI���dfN&Q�ӑ���1VM%U�&YaQFIfY����&fQfY5QVK�FFYa����deFFY8AMY��d%��9dDVKA�UUfM�-34D�%Aff4fb�e�X�.f9�S�fe�YbQ��f1P�dY�M!Y6b�dd�MQFfM1d6a��91Y��4�VLA�QCKfU�.AY.fE�Y	�2��Xa%�NKQ�eTPd�McC���.fT!�DNY5M��P�Rѓ��Ed�FfP9EY���CfFY@YeFALCMa�$f&BPTA�a5�eU�Y�f1YET9aY�EeLEH��T1Q6a�bd��T,UE(��D
��7:�G�m[�sz�y]a�VvV#c�YĮ���R9��� �K����Ji�ܭ4�=�9�J�K���O�H�g׽�6t���/�}rl�^Bxp�$�UH�0VLw�f��n�}�)��^#e���]���ls:��{8)bl��7�|qt�%�z$��{L�"�g�M�"���ZQw�+Q4�h�́"\��B�n�2�4�xDוm�1��EK7�`7g(�@��̻�ю�Jv��z�C}�r�D;�|B��%Ք�yl��W+$K�V�T���eNnKc�oB�������ы�Ϋ;�x�ͺ'B�0<�n����zj�n��$1I�C9,�����¶{)�ps'ԑ�J�������ɇ�gjP`�Ŵ��(t���UR���;�v��{�[���)Ø��M����JAx�����V�%��I�C��mN�H���=�������j?:����btt��c<�>�f��"xh��ڼ#���Z?py/�¼���/����*M#L�,@�n��������x:����xU��i�����ٙ}�[�&��kF���%rUc<D��(q}u�{�m����hשJKN�:�^���b�dюࣻD��i�+�S�~zn���[W�J�iN2��3&�=�ti�>��Ƨ�Q��]�.�[N�v�
sk���s��o,f�/rk��W'O&U���ŗ�1bPWT��wVz��l�p��:��ks��_ ��J�	V;�Z�'QΎ뮇��`Z9 ܠ,�,q:�S>�p��|s[���dqO���\�ot�q�]^
�fy,��2���K���>fP���]A_k!��Z��)����a�%1{�լ��;��.��6�����8J2�W	�U�
t7K���^����s�]OF��>ji��}������}�g�:��zU��!�U2!r�G=�����wG��QE�:��u�i��N��HY�]SB=Ji���C��|��q�tD��C!s+Sf��]�/p�{u�UH�(1B�m+��l�sc�&���Z�[��w;�@��cj*�7؏��2�7���J��pJ��QŎ���N��LLwt�yѥ�[���`u3��AM\��Oo�{
���唀�=�7A��7��Q8z��.ֵ9ύ�V8@����܌$v���q.������:F�+�������t�@�y"�G��,���C��kn��r���?wO�y������o;];W�X ���kH\�c�s�:��) �+$}!�N��>;i�d�Ռ�̨z��[�����}�c��V��;�>�ێ�勡���y��7�������ϝ1�7=:p����ʏ���b���}y��E�uJ�g=�Z����l��+b�������ZP\ήI��3%�e5�6ٛ������#}WǓ��Y��!v���kҼ��9�fkm	�!/ibR�k�W���>�;�N�p)1��ɣ/g�Ui�{��u��pМ�yM!��Sf�[�ci{ ��o'wWf�eaC�,]��/+���ab�V��� AE�m'�w�޶k�����u����s%cy���
����9V
�L�]��B�^�� k�:��1I��L��/��s� |����e�~}\fu*`�2�D:&��>P[���;R��]���{�a��gT�[畷�:�L�;�����lt��C(� q�aUyW�Pm�x�{��O/N���� �B2��E����x.#��=Kkh���z2Ǔ�?=��2l�`�86�ǋ ����;v�Tz�'�JJ49�P�n���$����Y�@㚁3��Ow���,�G諐>���"&"�2zҤ&�|�ҩ���B3�cB�*I�=��Mp�n���U�*V���;��p�T��F���B���Ya޸�#��ʣ���7�EZd��̏�r�O�{W׻��=�W]>6���ν�Q3��_R�[-)S�K��'n�b�GV�p�q	��%�iDgL�y�97z���vv�5�z�!� o�u�ԒG[K���#zs��w#�*)�/z'�n�~K�۴z�����K��e��m���W��(u\���(��EܡQ-U��0��:\t�j�v�r�ls���=YA��%?=� �P`�<=���Yڮ�v���<�{�
����	�i��_@���;tY��+U��{q].���t Y��@n2H��H����;[@���5N�h��J4:�rc�K3��_e��w���L���0C�R�n.Hށr�H�3i[CMզz_F���m�?,�~�z�2�K�@�������-q[�Q�%k�`h�RX��q�JysӮ�ݡ勦C�C��d��fN�ɔ��1��*5�r��>�YZ�ՙԖ=����E����C�le,^�U�����$��rʖ 0V�$E楡�\�����C��d���-)`����Y)/CV%h��ӵƀ�!�����~;Hڋ�ܝ�Ԕ9V5�:9���b����Q�s2y��z��=%�'7Ѳ�6����7VF�Ũ�e��q�FQ�����i���I�k�8���Z/�N=Y���d�B]Z�Z}����֕u؂���5�I,��p��N],�\����[����U��؂�Aj�0�Ek���?o�����c�{su�#��_5�2
�Ѓ�zC
O�����5n�1>��;�r�b��E���Ŵd��+=�;��:�S� ~�I��q����[��~Ʒ���\xEz5�CO\�u�6��S��WZ�³ի��rW��d�@�1��L�VJ����[o�:��sxL��Yc�hG+d��c0���ȥ5����̆-9c� �K	\V9�����bsv�w��]��C8���1&�!��T�빬G(��Y�q9���[3]���yc���9{�f9�������h'P�%Ҫ@V��3L�꙾s�M�dcr�o�ގ�D���&�X5����:3���T<ډ���.�ĳoD��0���g��Uo>�)����)纓C)+�j�#L_�1��e�0���C	�T�����B.ʒ�N��	��w{��c�J�<w^����슘�t߆R���E\�R7ԩ�T������{�����������VM�E�ϭ�F"8=�S����`X�l{>VJ��:�����]�Z�/�^�z3�t☱��j0*�q�p��Y9��٥��ڗF�
�'w��xK�eP6�B�~�|a9��^��jڦ�Ռd�L2sW����f.�[���\�|��_P�����!դ���=��ܑ��	��#��.�o3������ˆ�W2������\mh�����ux��ћ\�����Tj&-��'C�|q���o�)h���l����jl/_��%V�9�'�Hi���^P�^{�4�uJs��W}vK��l��3��198G0�>�f��C"xh�9ߎ؋ ��G�5Ɣ"5����N�� ԝc�����������G���hɯgǨ:�����1�L;��$�%N��^+��_kݗ�5ك)}��B��qA����뙤C�H��J��V=˗��s�5\�#	eޜ�+	��@Ld�,Z��mL��t��X1��9G#�j���cylʺ���1�3U�Z���W+LfP���]A_k!�9�mL�����Y�=�e�ƪuhɝ��\6��n��u�i���CF_���2�%���a�j3�@�/���w�/#L�ri���+��,4n%�y�9�Л���:bAQ�����c/��!sr��ҫ�]��eB|T7���./:�xg������.���)���m��zI�]0,t�<	Ph�;�sO��P�{E��|�� �z�W�����0hu����ZѴY��`%�����N���Ym�Ouߑ�����ܒ
'3E�920�8,:;�=��/�I]	��̼��Ц���SX��3��C�R�ޫ['X���N��޵*d���]�a�Һ�cJV�"�]ʘx�nF��s6h������q�{*����%T���ܐ۔aC���H�����(<'̱��.�������O Xր���� >��~����d^���A�E5p.u=9�a��bu�G�)��st�YXJ��M��Ϧ�Cj�mJ͠�m�@��	����F��S�K�}��{��8<�U�����a�/@�|��=�ہ0��4��ߍ����O����#]	���v*P��)�"�T�du==��K(_�xJ 8�T;s#7UX���\$m@r�И�X[)�5p�rjێ�5���Ӻ�C]=FEG9�L�7��uYއ	\�y\�C�)��N����Ѕ�WTi~ōUEo[4�p�|�_9�K �O leD�.��kݵή������;�c��X**&�a3�ںB�^��9[�<w��N4���3C�nW�v�K����vɛ��/��#`�6�Wo�)ΘYei0fi�������x(�Ѩ�<5�1TX���4�s�hw5S'/̪A�-Ƽ(iug�v��(=�w�j�,�5�<3g�z�h�e��N"��f��'W�oi��}�Зm�7NBl��s+�uncze��F����sd��8�ۢ��Ȁ�ݚ�L
����Ұ�'y�W\��5�C��C�T�{Ω��Z݀P
v\ܹEщ��3�$���o.#����ef7���"���P���fxʊu�X�뱔}Mv��������X�OU<�yFx�+���������n�}Iȥ�0��_=�5C��OԒ����OX'ֵ�´�8��b"��w��s࡯w'�h�;�#VLpX��g�ѐ�WfnMϝ�8S�F=�,�u$h�RT�JFp�-C����Y��7�����֮mN�o��.� *��gU��V�}�x싃��pL5�7B��9|�֭�)�aqs�p�y�%�� U�c�a�@�8�dKeF�R<'&y+*u�A�nl\�O���؅��q����t Y��@n�Q1F�Qγ�6qCM�uv�ɾS���4���{��ƪ��6������bdEl��C�lKUu#����u�^d�u���\�c��'tD�t��A�U䁫gY���t��X���38�U����kv�o�O:X*�N'�1C�z�!)����-���E�/���U 0���@�hN�z�峝�4sh����α�\N1V2u��b�̍��W��yu�Q4��m�1�٣��כ>>�-t��6P��s�*:Ӌ���knx{����$kc|f�p6܅�+�LK��˗���ݤ��j��:��q���tau�U��ylE�]�*�U�W={L2�(�v����]g <�և�<����Z�9�sJ23���+�`a�ɜ�X%�����"^��J��.�u�{% BŽ�v�׏s1=��0n����=%	u���փ'���gGXq;���,a;�����1�]�����#L&����,�7�3^���g4Ⱦs'i�n^#�d�^f))f�s�}S{�T&�l�4��x��� �)��~��D>���0cY�������..g&E${;Ȭ�7X�bn�]��rWL	���#Y�WR���LB�#�Ɋ�o��˛����Uw�k�[��
H����qYׁ[�ƥR���܆P���a!7b�o���J�{���mL��Y]L[-�����0��*c�v�aH�(�s@���S�Le[�}s�R�L�*��\)��P�R 5\�4'�W!*��亩�:�� ���%�<{V����p�A.���N%u�ߔ��F{zX�y�P�����x�m���0���3�]}O=W�Q�|uۣ=EH�yc��[���ߊ�C�|�;�b�U��u/qƄ��L��]��5{Q��җ�!5մ�W�e�f7�M)O�������g�`��.��6:)T[�l{�����
���7�1V����_>�j&)靳�rR���~��쨠�K�Vw�*�z����-nX�:x#-���H�Cɞ�����K��ڲ.�g����{
�*,vJ�Lb�U1����V�,e7v�&Y�UC�5�r�j�D�C���e�ZU�O�Gz�Q�g�1)Q����c���.��(�D�Z��¿h����9�\HC���`�\��j-L�<X��5�1��hw�T�WhD��<�:x�t�ll��&؛ O��L_��p�辅x�F_��U�NCn�a\v,��M��ζ1®�"��Rk�z�B�Q�"���u!�#u��n�ұ5���G6s]�jf�(/}<7fh,���:�34��ݜ2.5�O�W	���T+ʙ������ԇ?��4�6d��gC�f0V��<2�6�yR�\<�VKFr�x�Fg�~TϥE�����K�e#{��s,�� '%�b��3~S>��Hzw��5oz��1nW�waw��4�e03�]�q�GL�(s�U��d?������
�Ȋ�+����+��* �����ED��* ������ED����+�b* �������ED؊�+�* ��ED��* ��������D��* ��Q�ED�ED���
�2��ϣ�H5�� ���9�>�;��O��R*�*�(�����I��T�D�J� 
�����B�$�UQ��
�J�B���R$D�J��)�B�PQJ�Di�AQI"�HKL�T$H T*��T�""(J���@���P5B�TH����T�3N���A UB�AI!*���	U*��LT�T�$*�$�U=��H���*�UJ���UT�R!"UPWYU R�x  ���H+h���U(������ 
V�a�CY�a@
�0���fJU����T���Sl�*BJEMf�  a�@IE@�-@4U�ڡ�R�[X(M�F�� � ]�kJƬUhf���Ws��)(JR�5E)H@<  �4)�5��j��a 1��
4� ���SQ�4��hV�V�Kc�����B��əmm��:�i�)H�T��Tѥ7�  ���	��TaL�ڰ��C��ۅ С�CB���
$(�
ݲ�(P�CCC@ G� P (P�Cu 
 �P�B�r;�
(P�B��\
 ��'HU"�Ak"�"M�  3�����k[e��-�*U-,�l
u*m���h���:�hsJ�@V:����4.�h��n�!��5I�J�RT�+L�J�x   �ͦ/X遳��R�q��6n�mS��:d�d`�Z�`�݇U*�1l 6�s��SK�@�%�5۹��-���SE��"�mt	$�D(�x  ��[5���dom�N�K�5f���wn�ږ��� 6�*���m4�
m[5`ڭ�+kl�Sl5�h�V���M)Mh֦UB
 ��$YUV�  =�����ʖk�ѻ0�P6څ���\1Z���T�jV���]�CK`mF]n�k��Y�Z�:u�N��mn��aF� �Gl���R�<  �q�W��j�MbT��N��l�k:Ӷ�3C��[�4M6���C��4a��	u�6��6멑���]RXT�BE�(��Qo  ��=NԶ�n�@SS;�'ka,ki���@᥍ �4h�`(,�m�-#h-�EfLV�T���*Pa2 S�0�� h���a4��M0O��D@  D��
�� h �I6U(��M��}K������e��9�;-%n[�s�jIJi��eX竇s�01b�р6�U��꯾���I�}���H@�y!����$ I?�H@�bB���BC����_���?�Un��fG�f�赉���ɦn"����-�?�}��ރ��cKkB��`�!� L�7�+Y,�k34�,�p�6&m�͍V��f
�s2�R�b߬Y�\zN)hZ�����T�#�h){VS�e���#���28�J��GJ��PE�����}�޻�-��ݝI��� 4)
���\ku��������0
`�U|���`��ó>Ct�S�!H���N#�An<f\w`Xj��Щ�?�9�40�)V.��Mc��<��(�̡" �9%ȺKd�V�w�֬�X�0�ĩ�&�� ݷ@�]��-�ݧ߷)l�E`&A��a��<�b�h��(��]���xn�Z`q�d��72�)�%J}b���
2�ZL,��xn��{u;	P�9@^ҼE]@�+"�q�'#ת�R�C��#�u��Y���r��[V���l�C/h9vc��
�X���,f=v4�ٺ[�R�� �]�8���4NFE���,�:��ڕ
���,��F
W���d'/M�״h�Y�����`;
����ׯJ6o^�J'-cg��k�YͽHl�����Q��ʖS_=z��oLq;���)�k���H���*9�*� mi�\L�zJ�N��b���Ւ�Xh�W���Ѳ����J8ܸ���pȪ�J��vmh�!��&��b�9A-�6��
L��˺��^LW`!Uf`�E���{m�WF�yO�.��a��@��E�I
��E���f����m�VRW�h�Ȧ�^�e�s ڐl,�I�+cZz�>�l]XU��~c�N
m�BXڽ��L������/t��c���&ɍ�n��L��n5�ci+1�+��5�Cj����R��#0ӧ�K���*M�C6��ݘ%�yP��e$ks+4 �\�'Jf����#M;קv�3ae1gRBñ��[�21f��Ų��X�l���Op�x�F�a�M�J�iɫ6�0C���iv�"۲Ke9��vM�J'�j-� �E�O�D�n�wRGO��ݭ��n��+n@��)I�X�2�R���N��sv�=G]�%Ԛ[B���0�^��YM��T&��f��56�y��[��a,3\�d!
���p�4��%Lf��`+$[����a���\�CX̖%l/H�i���Ŵ�0�l�)������Q��o.��wr����TW	իpǱ��Dۓb��L�wY.赈#�\��a7wd��)r+`�ߔC���G`�&j�d-Y!E;r��.RZ�1�<Ԍ��H�w���5n�3j���eX��]b�Iu	CN�V�*���7���% �eI����5 �,��ջ�Ӭ�v:��/+(�yg��v�D�n�h�I؝�;�8-
�y�]e�'�o0�b�Ö����A�U&�7�m������iц#j���X�w���V3p����lx�Lka�)�Z�t�M��ѽtH���^�"���$]�b/6�E�e���i�-b���n�L�Eplc��1�{��,�E���.�2I{R�3����$�d��W�5ú���e?��k����Qq0�m�Q^�-:z����u�j��:���餣����Ɩ	36�Cq)W������4^ђi��%�n�5�����k{�mGy�k)CYfXc+ �r�|m-:�Q5�`��T�2RH�C5c�A�,Y��so6�EEY����퍡�&G%:�1��G1lucN�IV��Ջ+�P�c���]��`����l��Fb͎Aw,F ���@l�1�#`7R�V
օhr�Q"��,�ԩ[v/.f��+F���s�u�
hT�XV"�X����Ơ��7c���rPv(<6�F���EmhCÙ��U��˔�T��.�ϝ���Z��q���.q�H�@�L�RѨ�ܥY��p�<��U2�z-kp�u4l�C��M�m��Ta3� @��K�m<�hH�6Ň��
��ZD�����,���8E<���5n����n[ ��u"eV��Ym�QYD.,U����Qȝձ�`N��n�ѥm�//f�� ���Ap�*���BWe�Xۤ�eA�PAaPë�n%Ԙ�BZ�\Xz%]�!�W��e$��76�R
 m[�M��*�(J6���oRց+h�Q���oie�A�v����2T�ZۼIT���b��\7E3���4�ȡn��a����T�3{`씴(攨����a
�]�7V�\�X���лð�� D��OY8Â��ԑ���fh*�Ε��m7j�v�[�u/�3��P�n��ul�ܰ�՘��5�������t�:S)Y���ʚ۫�l�Tʼq�ҬA�T�DDU"n���fL���m���v�E��Hl��ut�ih�����ۤ�EY(M:��	CQ�r������'mn�;7Y��Ӹ�(ֻ# YL֊�>-�-�uo��60@�Wf��ԡ�r<&�;X�e�Է���͊�͊�P%�*��?K,ѱ������&K�	͡�����۩1	��U��i���ӳZ��ϔ�W߶�F]A�q�N�Ƞ�U	O��ݡV�;S[V��%��sSkv�Z�K:X㸤��G�`�^�3T�ѻv*A��a�JVo2H�٭Љmf�mQb�
֍O��Wu�AX"Y,�+�r�hk��c9�*�-
9i��ɟn�YF)��t�-��r��P�i*�&$r����V\$�Wx��V���nP)+�d�z�5Gtӳ���	\�T$GM��t�D��b�%e"ΖBK����d�e�ݨ�kRR�ְ\#��`��[����fJ�1��iR%�,f�0�@V���F�x�u0���J�R؏0k�!��8�"�&Y�3v=�sme���%�bhB���X!�-��k/ �,r� ��CB�佰4 �7+ь�z������'�n�
&u�׮n�%�ĥ��\�(\�q�V� �M�Cd%Z�!fa�h9���Qc��i�*�3��xB��c�C5=�Yln��n$5���kU��[-8+Z��͡�8�Uy����T��PܻX��!TN1��!:H�-���c#wun7�6VBo5)�i�s\�ƭ��2���Վ�b��;�[�[�P�ɵ�c��-��ö�⠈��af��WL{#X��-敹/T�C�XNL��aV�/Q!-q`�nl��ѱ ��Z=�tr�9��ǚ���Y�i�ݓF^X���MeX!]-�7q�P:T�
XOh��HK�܎�ʺB���-��өn�wfG6�`���iR:Q����7*5� b��cu�	�Ǻ��W�4*�U��=@fM�!�D���PZ@�10�
�wn`a�W�xaxp�/��3���)�@��U��{aSQ�ud�#�7i���6����]+�5������D�n�P���9H��4�U�����3.����r�C3d.���	F���X��qY��am�%#�/:�1B��y�u������ii�j�@��oc��/���H\�l`���I*ϯ�͍�D�+�"�K&M{[�A�du�u�k��tI���Ĭ:���bGa&1���u/rd�9������GpL��M�Ee-�J^�ڲ�8B�j�M�v�[��lƙ�EnF����'>�s\��ҳsU٠N�1a�� MS-�P�f�zk9�:��*ə%�WPb���h��"Y�[j�u��V�(iSe���Uǚ��It�6&�vP �FS%5�oB�%e����1����k(C�a��&�ۘSx�٫�K�3ڲ*P7>aD��^�)�N��]��Hv��Jk��Ai��u�}z��֪�[� ��.-���@T�4Lv�dhၺU�H�P;x��{����Hq��p_���X�n��su��9QY�҉� l��!��ϖr�D�� 7e<2���#Sck2��e+�ٴQkd��R�[ut04M�-m�\F��C�J�dgDׅQ��/N��
Q�o�C�e���cS��f,��BH���r$�}�h-v)�������(f�8h�;�X���$�>nDޕDeee�k��MZS"��n�M��_T�ؘ-M,��A-fY2��xp�L����M˦Pe��o114VP.ZVa��G�e_�^�0⸝;��i��ƶ`��i\�"[GS��4+C�-2���o5�pUH��K�Z�t��%t��tS��W)j��^R9��.-ەiӸ�i����]�l�s�/iPXj�̸�[�����Ђ�K��b�y`�̼)ň�/Y�M[*��#��Xt�/qV�kU��![i8@�x�AC؀�N㨕96�젝�[�����/�`�F��ӊ=cʏ,F^mB�5�h��3)L�AS�P RgEX�d��Ub��ꥳk��#�M��p�w������=kk�y�Cn&vY�K��uc^ef!��9��Z)B��'�Э���ٗy�n��8��C�.�l��M�n�4�1弩�Ed�-��b���]╺�kh��)�8˨.�L�4ݓQۥ�V �wC1붶����Zu2�e^⦴fe��Q�XB�iR*��Ѭ0�Ī�Y���6\�m妪LFb��K���]	�5a'e��ݺ�1R�qM&WbZb�j6M��l�W��*š��l�;[a�$Mj���ot� VMWA�^ָÀ֭��׹��Էq�b��Fز]��,E5��v�ū%in�ӱ��d�g�lA� �vta7G-XCbrB+F��J�L�ZM�d��AB��pա�))��2�A7X��u�^m<Z�#=�bQ%d|Ȱ��	�u(wsb��+1��JE>�6���,ِR!��z6��^��r�vC�,2�u�#^ؔք@�����2�e#zf�n%rnC���dV�ToU�f���o�X�LA2F��a��#�5m��\;F"�š�*k�Z������z����[�%�7Z�����c�zE3V,�Dd�&�Z���C�	�\2�ej�E<8���(D1c��,ʍT���6� *�w@mj,;����2��o":�&��MA���[oh�-֭8����9Y�[̛z�~�h�VE�-e�)�t��F��R��S	ưdǨ�ɻ6�Y2�
��t$`%]��X�ի�:v��**���I(�:̛x��B����yN�8��VA��d2ԛV�ш�1J"ܺ�ِ�%E�骕�2���`�X��5i�2 ŷ$x�4	�|	k0� ݊����W��%Vޜ��ŗe҃�8_l��R������u�>�l�P�Y�Dc�z12�u�fٲ&�ih�%��c�Y�� �!6�]kxP��:���ㄗA�T;6`�i��A�Y�#h����*a5h��
WG�y�h��*�m�t�pYF���l��5%�ƑX͆��m*�.P�GhI��M]2��{&K�lB+Q�b��nEnLh57E@pἽ��6M��r=��n��`9Y0�ֲc�P��*x+���j� (4 �W�((���Ց���/]��2�X�Q�dX��i�H,��*fj"�
���6'F��yC��"m�i��j�$�h���@�L+kn���p�dLX�
ܪ�.FY�n��y��׹)[���W��ǡ��[&��pQ�.�e25�Tְ��Nf��-��M�Bi��M୛�a��vA���ZP�P�q2T۰���^)�����f�b�4�	�n�h�W��;���$Z�cB��l�BV�+"�@�)LB�f�4L!��]�(��yi/T���]��"��[*l��j�e�ˍ;����Z�ml
n�ZʓI�j�PZ�tY�n�oQf�{kW� $�1�3j�Ni{s-P�@]�rk�[2\��
6�k�;V��+ ��Zȭ�E��+��[�O�зk�mn����)��Mn�{���k��j"�[e�B��^,i�nSF�cջ4iec��4��� /)�̆P�T��Ѽ�-sA�t��؉ݩr�i�ӷ�R-k�MP��m�R���Ԏ��∀�2TZ.�:�]C�lR6wq�P�.�J�zf�j1�&�w2PI0P1�t�F2�T��8����C]e���
�U��n����B����Ty	�2�ԭ�T͖�'�e��h��Vz�ͬ�S*�j�Gj�%�F&�rd�D%[X2�,�B�$��pf�����fG��5�,hc�1�,��=A�凵��0KY��ݖ�s5hˈcű���<���VVQ̃Y�:@�Eiֈ{�3���e#��k/kl�oA{P�ov��(�Wwr�sf��-f��"U�"N�k4n��!�8�D'�����a^E����*�V1�a�ю��ӣSr:`E�0�m�u���ϥ�wuA��W2�b 0����Sj�"@Bĩ��"�B�������m�t��2Z�d��j�Ԏ71͔n�P��ȁNӗc%Ū!Yp�%J��g73�h�;�/,�:����l��$�XOl]�a�Y���-�H�%y�l��72�w�lnRf���c2���VabVρ��4c&V�d�-d@V���.����O��o$�Z�ߑ�"U�޷7	�B���d[�t"ٲ�:	�6��۷cM-nb�b�9{)�p �F����q+L�1n���{�-�E����v����Ն�de�������	*��6���ʴ�Z�k!.���-J5! #�F�̂�"�a:RYuxtVՍS�0hRB#uoA���yz�!B]�ľ׸'Yқ�Q+IU�YJ��)��@}����r�f�5J���CW"Q�-���#�l���k��z�
[�k�9.��h�3Z��|�li����r�(�`�����Ȯ�P����ׯ��]�L]B闭�(wG�,T.<]SX��o��4��&]��q�xz�y%_�B�B�ru���Vy�����[�Ԫ�Z�D��ĥRө# u��@�Wٹc&��l����3k�8'��u�P7�,�oI��ڬ�\�I�=G�s�
�\O>U��0e2�Vr���g0��˅��C|��-�ܸ��5f�cZ���-��jQf��Wj2}2��5T�{��ċ�E^T8#k�U�D�y`s칯ffGU��rt$���ױ�eӶ/�2�z��:�:��Z�ٶ��On�Kؕ�'�q���U���m��͑�,31���IRKF��ߝ<�S���Ww�,K����ܑ�R�;��p�9
�-��3>1���-�΄֍��� l�%˺}�nӐ�ż���@���mVV-��܅9c��<�]HK�[y򙧾���`��i�J���׷m�Zckq��f�������<޻ոu��bw<���o^�G��9��K���IQ�)�'�[���D4}�f�d,�Ǔq����Q�������~���qLn0�P�<�SNI�0��md��ԕ��_P��e�^�mΣ��%�K蘶�^�\;:i�v(�����t�sQd���R��ð��Y.���z:���7�?i���Zë�;/y��6��Pr�7 ��1����.0�YW�nF]=Ql\�el��>ћ�����']p{�ޘ�?e��x
B�9y�N�V��m�
��w��¡9�WC�q�Mg$$�ݠe��kT*����!uP��+��7�1�#J�N�xU'�75e��p��FMz3#�L���t�r{:���Ǳ1-vL����`BF�b�!N���%Or�Vi�n���
�P�|��$Ǖ���U�B)�᳀K�[�y۴�A���*�.eIX?#�	S^�XVmb���l����hq�8ܒ=��(d��$cR߹�8�D��^��5�����t���b6��)������l�H��S�k%sҸ�涃���b"s�lK+��:U����H0���3"��]YV6܌ڗ1�4^N��)ܣ���8N��Z�K=t��"�3�k���7����[��:��-v���P.Ӓ��ӯy�x<�?������[���u��:G�-�a1y���j�MC��Q"�z^��:�+*ƣ[�ƻ�\Ϻ�����0reh�����Y(ahŴ�bC��W+�f��c�}\)܉�r�U��fR9�%�%s{�_q��Y�0�&:+�1syjqP���{@����7<T�GJ���qN����t����r���o���]N�oGF��&����:�׻�Imm���:�G���j�Z��_ ]o�e�� m�]:*�,ooE`C�Om�T�f ��-=':Y�r�uh��D��*WzH���Ž�K�7[��ˬ!qEr J�Z���&@�9����i<�˧ J��״�fڱ6���:�eb
��)��tD�iv�����c��W�����K7R�l�I��r#*&
G�K����]����ol�a�e��Φ�� =\�gl�e�)�>̝��9��[����B��<��k����2R���x�`1���*��aL��Sq:�X���w�O��ʵT���N��|vR�t�4�x��D��Ԫ�)C�4�d��.g'5��D7��-�Ų�s���,��H�mt�Ȇv�q�I��&����$��A��1[GRL�vn�:�+��껧��1�pT���>�ٛ�a�sI��o7�q���)\����2��]��q셜�4�w��n���e�=�������7�S|b�X��@M��6.��r;hǂ��0��$d�:-�:-��gm���9VC�@պ�ۖ��o��͔�2�����L��輫5��iM�G"��9mc�g\KmC@�rxq�t��rm�p��8�w[;�=rgWN{L�3^w&��Ffl}��_p�I��%=�����O1���j�Qe.���;��A�gp�ri�QZN�(
�\a�s#�ܛ5;*��ucxg\�Rsќ��{���	.��t)s���9�F�����	G�ԗU�u�A�>�Y:���s��_�F������f���R��2���I�}.�6:J0�c9���Ь�⬆�3������� ճ�Ђ���ֶ@{N	�b��xjֳ �,�t= *.r��N��_Z��t �R�D���e��}(��.eC)��ג=�R��9�һSgk�$E��|ڍd̛o ]B3�$ǅ�[�8Փ[�5�p�����©E�!彙�ʎ�#�����]�m���8E��f�I�3-X׮`�;������<��4x�O��+d��o=��y{�vRZ���GM�I��B�e���[�a�G���їO�E�@��Bm墩�֞�m���҄j��yV�����>���S�\�+.d�;�tǗ>N��y�'u�dN���ƪxwvZ��*�iެS��e\"��n��}���x=�N|�����0�I���bǶ*��j.��^W{꘩���b�� �i\F	!♌�n�yI�s���ŗ�dY�y'D�1w1���3A	�:�*4�@�efI�+5�݁A̫碲b��ҙT)J�1]���7h���kf��t�7zGRw���-�qx�Z���тz�1v$@4�e`�/�ޭ�=\�̒��ړ�V ��r��]�Z)��Zy�]�R�R]���z��\�IT��g<Y��hE�U֡f]h��s)��6��g>ܭU%v�!VJ{�Y��LU��i��[���J�ݾ����M\�.��d�'L
vИ�X%WdS�5��L����o	[�'���G�5knvD��I����}��I��T�v:�J���Rՠ[�g�l���`�\(�l�%X������vk��sd��u>,1�YW,V�}�9�Ռe��Y�7O ������t�$��t�}Z�V�.ę����Ս|�5��N�;A��]����!��7��dWHP�^.bH���yS���ˏR�d!����T <�չ�0����z�ŉ9���j5���n����":�V��Kv�j]��hv-t�E����Po��T[��`fL�����*�h��ܣʮn:0�9L�4����Z��ExQ��ᙽ���E�nFb�;��<x�JN��2:S{Nt4ai������+e.�;����ī\���sf�,����i=�j]�ՂsS/w�~�^��JY}W�_u�(T+huh��KtIݍۡ��&p�A�a�V�+W\�K[�8�1s�.Vn �=`k�f+')��rmD���#
�|��;�I]�4�����?��ͨ�WX��j�Sȓ��^Z[�`�VQG����
�0���u`�F$�x:D��[�����P���:�z�6��L�܅0����[-P.��]9��\����A��b���}B�����ݷ����3RaQ�
�f�0V�8�g\���UʮTwi٨�I�݁�X 0Y���%�I3_���Gp�����3H}Hd�͓�^��7@����8k�*H~�E0h	;ڦJ�ko�j�叙��S���gE��q^o|D�T��{�PJ�e���%��*J=��&��Jb���]�Q;�蚾૬������PiJ[��+�,��H"��ޤ9o���t�,��V��"�dT���:[|z�I�'�5p��h�q��:�Y@���x�����=}}�1`�P!�ޥ���`r�^W�y:��BἬS����RCs&)��nqz�W�[�N�����Ԋ�Z�xw���O�OϪח�>:�wwoEx2��8& !<���L�b^��䛌a�Vk��)��(Z$]�b��U�Bȶ���썉wb�M_^� \���,�*΍��報�w]ܐ�xp3�����F�-r�����Ҷ�0Y�VG�Y�h����]w &i೙��[C������0�I��4���K'&A��������ƈU�:��PXMJZ_o��qx�m�/��+}��%gC���Ȼ�
�k���nuA@��X��2�WѬ������:Tnk��3���
v�}�[���k��x��'js�9��ưg)���'H��͋T��-��_7K��]]�tUok�P4�9��0��S�����,Um�k����&"֍�F���Q�6�tM_ ��k�N�W&�;��Gh͋��zrv��~Z������@s�J��n�N�՟No��z�LU�w��ͭv'S
�6E��a�v�ݲ��s+~�c��%�)�v��\�hW**3���n�G2��h�;e�2�8�L3��<p�ڽ�:�jsrq�X��4�`gږU���a,C)^�w��7O�f��q��ɲ�j3l��0zھh�������w�>$w���B�8�R��Kd�����lQۨ&7j�eN��&����r��K]񣘊����j����4��l6r`��Nl�z�.���*���Ve�˖�'g2�o�f=F�X��D�Ͷe�a��4��r��m<����L�4���{�ۡG�+�5������vǿ+˵۠k��! ԋ���G�3�$V�9�b��g������?[y(j��n���:�f�&)nr�%�(s�!��� KR*�fͺ)�9P�^��݂u��n�M4Co��[��[t�yY��p1,
�cp�hm�Q�U����tVq��/ Ωt/�Y�8ek�\�Е� _	���&�}t�t&.�J��K{���U��d���UϏD�ֽ��YVw����T\9i�F,�K&���#��_-�0rx�Sn;���eK�ɏ,�q+ =�)i)�Oi:$��`����t`K�E�V�(a��;����L�C*��v�,��}g����gA͹Qmv\*��k!CB�B��ao,�̿�\�ܤ4+���8�u�dڎ��Bɶ���Z;Q����)����B���Q�o[ۧ+� �F�'ۮ���9SZ�J��1�Ξ�������.��u���eX�j��p���[����L�-��� w(V�>�,C<D� ���K,C��K��5�V4�c��[CL�5ɼ����ǲ�s39)�l��|8=ښw���2fuW������A3v� ���Cǰ�w�֖c�Kc�6M���}Ƅ��y����)�i�O�X>;+��Y����U���(�X3�}H!)��ʹV\:�֟o2B7s�nZ�`�',7�U�^��+��k�i�a�gGw)w�Wc��.�ޭ��������
��	� ���;gM��"q��I��OH̓僬`����Vv��e5���C:2aw��y.�6���u�Q�*,�,�����Y�g�5���R����V�]W/�FX���E|�E�b�`�ϹaFsS�e��7��;r믲r��������q��/���l��[�� �?mh:�Ӎ�qh�����:�X�_+z�!������o��3�6W�G�����D��EBj�R��V.��x%��p� ț�
yY7,,v�s{���PC�ad��<��/���q8����ٵ�4��z��;nj����Iumr�ΝAbH�ͮ�6�(n$���;�_d�
u�7�����M�f�ŝy7Oj:��2�H
U��@��M{���w�N%+�9B]K����Y���;��Ɋic��;�<*YU6q��;n%kf1o�n�`[�f�ی�\9��40=����|�)AŊt��T�H����r��6��˄m�#���S�8e9(��E��1��%ڻ�iA���{��5%�`Q$�Pޮ��굒jĠ}a0R��VĻH��e�<��`io:�*¶�1�:�$�ѵ]4
|퓸Zu>F��E�XM̓���V��2nX��6��ֹ�D���:���F,�z��+L�� Փ ,�WT�z>���|j�wn��犆ם��}ZOV;5�]O�eě뵺3:-
xV����:��cS�ސ��7��ʴ�J��b�im��+�Ğ5�"�K�՘�x�8���	jj�{Yݚ;)"�:�����`$'K�uA�7+\ٝ���;P���;�]u\��ۧ���n�!8������w�qj㋚�^dǝY��%�;:�:�QgN��J}Ql�&�VS�k����)����C�\����d��.Q�Y���ة�fڠhݺ��sw(���V�Ԓ<1�p�U��AWj�fL�u�E����q���:f�H>��:
⾺j����/�^��M\E�!�n�sEL�
�WG�<�T:��1E�5��-���N�C� �K�Q���ve�"��rs����R��._8�}@MԠ����u�я��rS��9zpFN�`���F���T2���[����NH@y�����ye����w|�jou��E� ��T)�h���n���1�N�xm�v{��y�l��0b�s��Z(��:Rɵ9��:�':�r���"ztGO�;A9xH	��Wv����"��Bބ�:�7�D
��@�};#�!Tz�S:m�ܤ�鯞�VZ\�3�up�������k�(�.˽����S��w�Zo��9�G׮u���������&�i�B%ʻ@���ם٪�1'`�����K����s�-�ˏX*��vu%C�[�D:)B�P�b�(�IRħU�KW�R6���joe.KbT�z�s��:��9%��)�bE�wbI%���Kq.X��]�rQ��z�R�^�T�R[�j%�A3{��������G�� IO����׺(�G�|;q?=�g9{��k��Z#_\��3.�Q̕w,�e�p`����e�圳^��Bu �NKr��(�c:���]dx�|A,;��	��xL݇"�]Ƣ�O]˰5�íͿ�:'�P�{��pSDKj���w]�練g��p��N�9H�RS������[�B��t:q��ʱ��c[�7n�ph^������c���c岎��F���ï�C�<���5�Q�H
"�.S���r�l₝�[[���vk_bEb�$M���B̼=϶�q�95���+ذ����.=-CqJ��o)t�P#ɇ�w�/�e,��VG	H����ehRK��e�;OD��hA]�+��rZ14mmHeqW�0|:I��u`���Aᮩ�'ׅ�]���ڇoy1���;P�bKi���XN�}G"�ػ�����M��+|!ۡ������x�D��[\���xM]�%��%dqng%2�z&�{.,��Ûe��]��L��n��V�,���ai]r��]E�%���d��՘.���4e.\��\���4K�~��{�y��kQ+.�2eq�%�B�S�^��w,w	eI�՚��(�����gos�R��-�u�к�j���̢�J:`7�+�wK�hٿ�`g"{�}�ތ�����c�anfl���_ gR���Nw���}ԃ��\���� �z3Y.�Wnԏf�:�bݦ��!M*1�B���/��v����"F��.t��FY�ktk\#�L�e��,ӓ�}Ӛ٪�Cr�`��*�M�d��]��:�*����T�C���A]e���C�k4`�ooZsPM�NΒR��k�c�Dk\��}V��@?�>�J����=�y�ɵ;q*��H�t��bí��/��t��pw̢�2�p�Һ7��"'�wV3�M�\V+"�uu��o@�H���Lp��,s�[�]\2�M�.�t��r�q�}�1�D�y�0�,�ק �����Z;�r���i�oy������l��łt6��jo7v�쪅�x���Ӗ�Ξʕ� Z(�f=�cS��}�����Ї��،��h&n�GBB��<�c�F�k��.��f��;]�{��K�wQ ����ne�P��?83�[��))@1rQ��B-rYc)n�����@ۋyer5#�''�D��Fn�9Hf��5��27(�7���fc�,q�*7å]m�m��u��EDr��}��X���\b��=�2.,vTF����}5gt�sh)x.��S�:�yJ�<�oonڭ��5<����c�JYڕZ|���%t�ʂ,��t��8��o]��2�jƑ��3���ك*TwU��&�����MZ�Z�V8���yX2Γ�IY� V��)��
���;�RL[g::R����h���^dU(1�D�i��;n����b�x�F�\�N⻫v�$pH#s\���b;x^�u�.ٕ����es�>��H]���[t����ޗy���_�Ғ�<r����ZQ8�k��%i���������V�Y�,jt)�Ս�f��Ocf��}܆����[�0]c�*m��(=N_89�e.�6�f��u�(L\�R���y�oJ+�[ui9kc8��3z�Q�\2C���mD x�I�;��Q
�4dm2t�}R�J����b�b����)+��Իu�Xl8�:y͞�Qse.��K[[�1{W�w�����{-ٚ8j�M	vS���D5Cll\�k%l�jJuC�2�����;\�⫵��Ų�J�Ht��z���C4��։�#
��N���p��7D5uЎ�ohӌA�������^v<j����AmmA���NrN�oZ������H�E3��y�E��o��vWJȈ4yk�t�L��D�%bf���e��pΩy�Y�nm���#_[�9��EsQ���g�!YK��=��W�9�X������ܾ�-�W�l/�vR��"��a�u/���^��t1���MWI`���e���kY��죪T2�V$�1�~}�&�����Q��+GK���h�Ҹ%]�sJK3H5��ǷZ�U�nm'B��E�1�̔��9���ҥ�0�u�m�\o:�d����,Q��A��<��[q��y�LPw%��cՕʍ�X�E2�Yܘ���h7y}82�t�����۳9�z�=�!Mm�nպĨ�n�@j��"6=%-��;s:螜�'���x�ŋ���|�pç�,���.��]s��aJ����.���V�h5$��#�Zku)���(c�1X���_e���2���WwΟrsx�L�y�6�9�L��H �����s�A�V�u�2���L��.wƵ���Aa��*���]��7Q7��M�G!�K�n��1΄
�|����\uwػ"�ڐN3z�GM��4�:�TU�6�0�G�S���v��a��s�O6��5z������9(��]+���<|����CX�ź�ۂ���n��[y�vVB�A�\`��թ�";�6�G�O`�/o${�(��.���*�S��u�j�6�,ťz�}��p)��ӻ�'
�n��ȁO	�\��7��\�ˣ!�k[��gK8n>���AB���C������|v������sGP��펷��J�I2;TێT�U4%H^L�����u2��m\ζܽ�\��A5.�u�zeы�x���e������w�H�;�C�<�k!��J)^˸9�M��f�g�Z�K���Y{��
<�l;�L�̿��[����(�c>�Iv�}6���3�L�9[���VSڻ]dVr�g��w��0�)]�@p#��'�Y{�ʭ�P��h�/^-���Qe���ٴ+}8�Z`��X��,"�6�b)����u��h�S�HB6�m�V�i+m�L.���p"�_'u��uݴ��}a_""� ��-xط0�e4F�R���9_�b�>K;�������8"�7K��l���9ˎ�7�`�z�W�,0\%}ۭ;� q?��nn��D�7!�-�̔��;�8�]m�jկ��p�m�Cx�X{�w���R�8�L��Vh��w%v�#�uA޽,iT�Ѐ��A]E�Tڝ����ͻ��+�-�i�1Wy"�Zu9#�ݮ��LA}[�HAy`[O1�R��C(ܝQ�y�����Ȋ09g]k[X\����w��M�U��q����Z'rݱ��vw^1wVл">!���� ���Ve17�E٫	0fe������k�ծ�j�Ig6��*�|P���Ge���Z72��ו��)l�W�b���lL�;� ��a��6�d��Y���ƶ��!T���ݚ�CT\u�p`�µ"x{a��{����.c�ۉ�2�6_[ڹf��l6�卑mu���FJ���reKAAv����Y�3�-6Rm�D�Fr4��,��l�d@�c�M�f]��YQ'`Q���C�r��GJ�({�Jl�ۗ]��N�����2�<p6���*�PV�$S�j����V�G��Jd��%�|�ӂ��Kߛs�8��<�U�:���]��=����z*f�2�#��C1���]�xq�˜)������HJ,���Y�²�]����(f%�6nV�T�S����s���jf�	L-f���kwt�W[Epeg)J��`Jū��R�[Lq�ǹj\�ޯ�#2�iK+R�d_=��k�ZM��VX-�L�3�r�#��ShI�7�!�ȉ�X�	a�Օ��@�̲����[k�a�<�,��j�Z;krYL��b�u�J�<v.��|�h�3(�h����卺���pR3���n�R��Sq�R�FK`>�
n5r!&1�����u����h_fp�����Rϒ�w�|;yҌ�mJoэOi�Ш�W[�FoL�J�Ew������Tۻ�ɧ�X���q��G2\�#�Q�q5[gv�\�yȝp�S�� �`޷@��H
j�����]u7��Է�oQ�W���f�7��v_L`�sue˾��l���RN��<#��'sn�i���jU.� ]��Nʨ��l�}�,	`��m����"�����;���˱��Bk������[�J�U��9�S��vz��Ծ��4�k�� ��X��e�S��}vɦF����Z�${�ws�b�Cԙz�ݡc(S0�ˠ�L)\�3;2�z�J��#G�Zu}l�wN�ի�o٢�4�e.��FN[45|�q'*��mmc&����E;*�Ew���/{���k[���0��#]�uuݸu�I�S91��0ob��u�`��nnj;NP8['\y�p9��ʱ�xQp|�c��T��FnWBJ��oI�p
(eʵ�h�ή��S�ޜ#6��5��vơF�vD8�p^�H�:j��:�����Ŋ���BW���Nn�Y�B��%�W1�p���!��ˡ�6���vÁ`تo!K2��:"��F	J><�X�0d+X� �A8By�aב*�5P�]wY��e����v�An��J�h�L�趙��u�e�`�-Ȑ�95u�k6m	LZ�+��X:dH�vd]��
�>���v^-�Z�u��� �\�ۙ��z�b�C&��pU�bpxU�Q7] ��\jo9��C���:�I��x�qD.�E�:�4�q�����{ s��29զ��]"u!ʕkY��5�k�Ro�_v�m�YNoN;
r�6��M )E]ó��7��t���x��D���8-{"\26�2k!9���|��U�Zw�U�\���^wQ�R�᎒��3M9d��pF^�BA��j/��:Φ*<�1�'z�y9��N��B�Î�����D��3�;��w�]+�,G7��>�2 n��:�C�}u�<��
�c$�8��2��&�A���ۤ���U����)#�e5A�}�XW%3�3���z%�燋�yQF�R�œ�H�Gx��2��rX��& �]�[�P�v�_��WN��}�y�+z7+�#��d�)`�����.�k�;���I���3l'@�AVAMQ�+o�������i�h���򼠖�V�V/�!|W�@�yy�+BOE�C�!�%+�Ĺ(����]Ն��N��c���S���th�:�|�['K�'uuya̮Stl9q�bV�/Lp짴��mfD�&�=�%��� ��c"�
лic��y;�q�+F��/,�c��3�x�������w��f�`!����)p��HDU�ov);�5����"/tv���)��4�N�������}���m�]�ks��u�����7�P�}N�NhJ94�K g��oKW:����XM7�q5��3f�h�^�Z�r2�p�%%G�)��t#bZ��,�q�GR�/:� iB���ocƍlur�V��l��h��c�p���8�ug��F]�\�)w��]7Fo�|2�{Q�1��%��`�ݛ3�ή�9����<�I= j� F�	ҧ;�@*��6�k�t����D���3ݘ�s��q��s��!���]y�r�Z$q�yy�������w�E�1"�ɱq����Bqes���I̥�36.[6n!��ACsx����[��Bb6��%���4��6@n.�o��ڃ;5�ӆ���}]-W0�]��oq���w����˙MVͧ�l��d����:nsy�����FT�O&�%�^��e@_%>��X�!\���)���\�8_�K.0�2m�1��&��]$Z�d]nV�ƦdU�S�͘>�)v�L�B��N�4I��.@��R��ȏt�H�vRȽ���Ѕu)�����p籍G�/k�9��{���vW6�U��7)����4� =�aU�F@�u�kerS�+ǵ��7e_Ɔ5�e&P���
V/;���N\�����EwGY�tSb�b�w��\���G�pŖ�+x�]i���u�#��v��}�^>`�MK7I�m8�͢+_uh=�.���'R��fgn��{���2���,�}D^�G[ܪK�M��� �����D�VGa[�J�Qq��E�@ާF��S�0T�YN�]t��gtt��^Q��X�h3��6�0=N!��YԱWd����� h<�N z�7�cޭv��ڊ��%�|.]�LnsS.��œ�-��i��ԒT��յ�,|����a�P:K�W-��uV�.U�tӫ4�iB���)A�pNvv����b��Rz%jǘ:}�]Xp��X��D�[p���-�4S;{>��u�4w�dd�=�Rǘ�X��ŝ���	:�H]^3��7��N�'��(��	�rCV�v2��s��-�H*����۸V�:�j�˝�x�gh^�9|�<��x6+��I,��ȩ��eu`��W��7�_WPFt}y6#,U��0,���Q����Kv_^	8b�A�K���K�W�V���׼��m��1�2��95�*F�!'WI���)��a^��M�hAS�K�j�k�ܨ�{0Gh.21��v�:xԳP^��E�]�2Q�v�v6r����������� 8�5�kS���Wc�Z�z]�h�]�*�bnwq��B]�2���;�D��*N�7.�I�c��	�;/��Z���j���Y/e`����:[��j�'�v�>ؗ^�t�G�m`\�}
`�8�NjҲ�C֖�a�B%t���fF�
,c�I��p�P���ܠᾗ��PH`U�WK*�ּ68�W��2�ݒ�镪]M7f �Y�=34ܮ�Jc|�a�ڳU����{o9+gV��x��ЮB�Z����9S9��8�r*���8�����S�-�č�q�\V��
e����y���y���zv��ɻ���;�<�
��u��Q�L��3��V����L۾�ʥ\�e_Q���jjU7�m�钞���·�������h��(t| FWGnJ�
ڗ�:�����P,�=����}�2�ֱK2�_=�Q��;N#�u�+W�IΎ��L���>���{z�kE�$���˸��Ɯ_L��.dP��Z�M��U�8lT0I�U�����9�G($uݖ+�/��)����;�N
"�n��^ �n.-��$)-�ե�)ޝ��.
0�s*��t�c7��D{���W��.F5��n�U�Ȭ5�%bң=��yٗR�U�V��u����e����tP�ո�=��B����+w�y��`�;l��:�&87�hͣe!Ԁ���\��Чh+�fG�Je�b3c�����ūw1j��N��q1�܌/ඣ��geguv��[x/�Z-D����u:u�}��� ԕ����xUB��3izĖ�ЎE�<�ʏ�BA�)1e!�(Aޗ�V��#
�6���;VKZ�t�2n����wf_{���#Sl�L&7m�Wc������'�C{e��;)s9VYݲP��wv���M������ѵ�L+��v��sɓ�.�\��NY�&�����Ҳ1+�#9�>}.�Vc�UmwP���"*��q9�aE����(Wq�1p�8c�BhZ�PN$�X��B�A0�>j�cШ�m�J�JT�Z�%B�+ ���I(֚�ĩU�l�%f�R(�+Pr��Ĵ��m�X��L\��Q�Q*
J0X,� �*�����1�CI&2�UY*�$�VAeI��.V�,X

�	Y��(��k�p���-V�QAeB�҂*���B��m���Y*���!�ə`�UI+$P2�UDeM7)Z�a*Y�q&2��-�CL����T"!X�1.4� �(ʒ��YP�m��2�U�HYi*c%k&1a�%`6���T����J���E4�q��aP�)+P���b�"b�2�Y/:ax^a7� W��gf-�3Z�mv 6�лG��p��̼�J�>�Jށ�gE�LYۍ<�����x3�[+���ı%�̚���&3��.��c9�����>�3���)����c��,��N�5�����n��xύ�)��*�9Q�	����)b��������������K�O���N5��5�сM����Br�y{������d8:�*�ko:۞�X�\�A]�m��C�����`N'�Y<��_Vd�7�U��2��ڕ�i�ŕ��VS{Qv$-Ll�EB�S�S*֛���w3�Me$�r�~s�I�[�C�;��v�"�hJ�H�Oh�MHڊ�[�9Er��ފ�^����qlsޥ�yߡ�ɶ�[6��q�Tw�e�v���l�i�B�~U�(;���c��U9����n!�Ց�"��Y>�5gj�SJ�xR<T8����T]bkO��_B��UD��V)���Vl��oq-��+�vl����{~�4+7�r�tU���u!ƾ�k)w�#����*]/C�x
�)hT��J��E#O:�����eq#d�"u��3�u�M�ukk�fZ���h��k}|�	dN+����Y�/���E���JA	��M�`w7z ��f5a��(��~��B���P���5����<��;�gH��]�f�������T'�M&4:����}>��=�hY�{�j �B�lV�8�,�Q=<ĺ�R�7/B�&ae���������W�4�w�eX�[��j[�z+�XL�s�K�n79N�f��P"�UgS��7u��-�D�0v�M��L⃒�W���ڙ��!�d��J(�f��:�����h���S�9�F���u�7��M�KHe��ç,�[��3��ry��8����ڮ�0�w�v�R����臍t8��L��C굗릳����ZÊ��f�)�3�elg;/6�Q[�U��ro\�V�y9P��.O.�:in���׈uT#kn�,\N[�+�=���ӭ�y��d�R�1<�6����.��Z�\cZ���$GBq#Wsn�[z�Ķ+N[.د_5Q)��ڻ*��~M���s�~��5�L�N�V�|���9v��x�5R�&
5g%u���<�a��!eX�9�AJ�:��13}��XUms��#�
�}�6�]�x�k������I�!�ïn�Β���&��:訷$�����>�,U��ؤ�ur�ͣ��L(H펀��D_5����嚡h�nM=ͩ�Q&m-T�:�S�<5�+w�q�p4%Xz�"���0���+������k���H_�M���ڕ�/ڷ�|2����eE��o�K���WƁ�ھ��:r��*�ܽ;Uӻ��Yx�8�B��oО¬x'Ԑ�^-����
I`�	�}�{�$\�&�z�0�r�{�QMڙ��>�R�<"i1��������2�z�3����~�KJ�U��Ř쫟Fĭ`�E7�9�+���9q�m�wob��8����X�s^E`ٵ�ϱ9��\q�����A-1ixn���{|��dӈӄLk����\Ϊj�DVc��zL�-��Q�q'@�Z�(و�u5�V�t�uל룛��*�=.��rWV����b��4�+�|ϥ���y��ܭ=���^"G\���-�Oy��H+M'1��'a(=����3*��GS:�
���iڙ*F;�r[�ݞ|�@0����c��+�[�=#yC��ީ7�	��w��t����<!�dL\��nK�A��޵��!y��'���yɴ�Y�k��˽̋�n�������NN�[������Ut�7�Բ����G��x���1��L�$������z�oH�Z�[)yW]N���k�ֆ����b����5:�r� z��'�:�{�^Ѿh�6f��}X�FO*�R�����)>D�:�Y���msW+��b:��uW�����'���J�y�-U��[N2�+&T�c���[U��<Oh��~�qL9c��)쀫�_5��\n僒�\�0���G��̃
��~P��ݻ�mqBU�t��PW��sv&�\!ּ%r��9���������[Tr�U�jUx-��$�5u���E���,�算����=���1��٤Q�&�Nf7of�KTUZ��x�T�N�&oW�Y������w�W�T[x�bܗ\|4�Ε����
1N-�b�W1��+t��8�m�s�*u�z���V�Xk��r
��������M��W�k��0��`�b����^�Wgr]�W�zkpSO��Z���ҷg��H��՟xϗf��@쮛f'�И0��Դy�vj[S���eI������u���Nr+�ٟ�1�QP�]υ3�]���ݎ�	E��5y�Z���$�s�;�4Ӝ��������z���}�>�m��=�?%��A\��ٴ~.)�����'Qn���>�!��6T�[Y�u�wBr��5M�'o慫�{��S����;����p:���u�F�yOf��V6�O%��UE��Q�4�m
���l�5�+�ށ�]	�5�9��.��K�V�MJ3�7����c�k��LJ��'��gH���7�+�/��g=X��l���"���7���:��U��9������H�F�%�4���M\�>����5��s6���ΥqG���^�9�2�c4@�k��{%˭8q8]s�����$�H��iu�ڮ�׳V�@C�;;�F���q�完3qϞ��Z��*�O+=YM�حGS<��P��,���zn�:��x��~�!O>|��~]p�mAo�#���/��B��ժ<b�H�c�~w�폵�����0�,
�lյq��o�"/ۈ{�U穭گo���X֌�=�Ex�ɹ�G�����-{+8��\�`���0���� �6�^����q�#P�U��3������
��Hk��Gub\swWu���t��>�r��z��܊镭v����y���\z���z�CO�O8�:��a�pZ�PW�as�}7�DNc�r|����X�HVN�}���ލ��ͱL�ѡ���غ�*i�x.�	�vkf;e�=�F�x1�r��}9��{	�Ȯ����x����JpZ��ב)t�;EU'�Ζշ��%7s�P�1I��}PNR�[�*�:�6���V���D���kɍ�|�|�hܨ���#U�?u>���_����K��'�dS���%�vz�+xNF'�*���=N��8m�,5[s"��cV&��8�<��&u�٧��Ui�1��i���r=Yݹ	�9�\籮˝�}�r�@�~#c���3y}*��u:�Ϋ<qw�K5s�Φ�	�[�����|��k{�:i�Z��7�3{ �o��=K���V1{4u"M��5pp��\����̣ ��w(\ YI�V��U�I�ꔫ%�g}m��ifpbs���ǭ�]���9�˼�t��,oh��$fH�������a�p�8���+��)N�].�ﯲ��f�1�=u��2���J6�8���ם��?{�{�O�A��\|f�4g�M��Ն�a����Ɠ8�����ֱrw�Oz[��x���B6�m�@ÎL�M_.imr�*�RN�2y�G)U��Ci�Ȧ���̾Z�82��Bz_:SFl�fY��)�dZ!��;����s�ݔ�<��Y2˺�W*b�j�\���zs��.
��
���T|*�����r�q'_�U]=��K/�Z�FO��mew���t&v�}v;�]�T�Te�I��;�3��CV'z�|�|6a⹯7,��@֪0�W9ai�q#�65��;�l�g,��]��y��=�n!=�^ǂ}I�c�z/ʚ<_JYis��g&��z�����糪�Sf��u'�M&8-���q�uʰ
�'����~Z���/%�C�U:�~��ۜ������ަs�6��=��4v��R�Ҧٴheޕ
V�sg-k(����O/���ޛ���l���0�bt˥��z� #���kaf�'ȱE7���X��@��� .^eV����p9�KE&��B.vu]tu2^�v�5]N뻡�36���N��ߨ�_�_��η5͍ص��b{_���iBUSJ�'v�^^����X�\w]m�!�L���Ϊ�v�M��c�f1GL��܎.�Z4l��,p��Ä��>~;�<�~�z�.�c��MqԶeu!}����� ����7�V\C�1Ҙ������y��ܭl�	�'{�ʙ�qv0sq��\�Q�qZ��Z؍q���O���l�̰�r	�ʽ51y�ƗOL]j�t����%xyV�ʈք�O.�*�kwvUfv��Óp*9շ��wna�l�k3xOZ�V'Y<�9J��o*!��6�~]nY�9�EC��볽�"F9j=q�U#i\B��:����G-P�8z��3M�p����N\]�yH���8��&0�l)슈*�T_5��;ל����eS��1���ڦ���C�|/bv�EF��P��{S\ܞ�C��>��
�c��j��I��Uc-種��Ү7X��p��1o�sW�k�����O��%�EԲ2�
�ʊf�{F�s쾷C7�4�s��Q-TS:�$:FEzww�<|ҾO`7��\Dt��R^���|��ٛJ���JGʎ���vA�~�NF��nj����J7��1mY�7,���6�;�2W�ۭ���`Vm]@}�~��:�S������ߗ���3�[ʕt�ƫ�_(�(2��
��0��yA���s���U{�6c:��=��z��g��R����?Z�ykc�V�S��ߊ��ġ��J��c*5J���u�G�=�r>��	���Q2��NR�u��+���	Ҳtkw��D�w�|�8�A�k�iӛ�p/��/�	�Wr�mj��]�s�ED���v���'ͪ|cb1C������)t))���u�9���K�W��4��Pv[��hV�r��j!����}o!0ɨ�g�����|`aP+{8�я\^jb|��I�d[@��EAo�����HZ�.Ll���^�d
�:����s��.c�,�R��n�]��Uܭ-�-�=���g���턋q&�>�ح'��m�(����>U�X��Ӟu)iK�7a4T6u�|U��L����/R��7�'ma�x��;�u�jd�O;q⾫|�ϰ:�G�;���QN�A\�z_�^�Xr>�j��'�O�A�y	����AM�Zx��+c�k�.�����g�>��1�ŝ�ܾo�ve�7�z��B�?f�S]
�V�m�6��Z@8�n�N�+���O+=Y�ok�v$-�LuR* o�A�
�ir�Ր2�?[N�r���[�C��|�7oQ�SY�sJvU�����9�{g���z�Y���sިZ7��P;*г���V�R�غ/M/gz�����}�T��d}v;���Y��s����F��ϡ+v<��9��]�\o>����a��Y�\U��ס8���wWv����s�[�&��O�'��ٌ�Lhev�Gvy1{5��-�Y���?r���Χj�6o�!<"�6&_T���wã7�26�&�j�άv,+cVNĩ�1.��;s��,baY��ӕ9�gҥ[M����� Zݺ#��0W[���<��ձ���{&-F*a�Wum�b��ͪ��=E�P��L}��箂G�:�Բ ꍫvTO@�1ň�9|	{�urҨ7�G&`X=���6���{-�����n�f�"���$D���XC����� e1+C6�sl�O��8��d���,WBA�{�l��=X�Q_Bv��m.j��j�oQ7��y���.�p�`��n_i���v�.��bD���;�DZ��D����i��8�p��������S�H��r�t0�ޕ�ې);�B�N!P��D��r�f�.8�\f��n�X�4�h�8�ܚ(�'�'���0��+�S#h�Y���,�)��)�-���v���K��!Ȩ+N�5tt�)!�̭��e�zt�s���P��J�OpE��#�����WÐ���ȏ�����R뙗W
�.W#� .�A�HW4�4;���º=�}�k��MO�f[�n�B� :wG]g,ɮ�=�S9kz�q�f�Ú.v�S� ciG�Ϙ0����[�[c-!-lB�PN���|��g-�,'cq�԰�9PpG���+��)�u۰_/V:pgbtNE1��r[Y< �-�0�-�&�J�y�$���q���r��OS;C%0�JGr������_W�{؛�K� �k���f��Y⒈QsWv��
�wUkJͮ�:��ޔ��Xr���Մ� y/�Y��ۨ���]
��Ŧ�$O$^Mw$o�k����X4�nIؓ���ʽU�0:�Q��p��Ժ�]u�S��`�{]�&p����Ǳ`�C/N.�a�^,熏*![/~���}7�ͨ�q��ا��[�]u��������v&<��R�yP�����t��Ч)���t�m�E�q͝Sa�fY�I@\_�:�ֳn�-�+���[�o++��\�(q����o r�!�]΅�h�CR�+o��f	��YE��K�c"H�^�����+����i�F����U����K�1��p�N�s2��f�h����n�N�|��줻�8�(���
�! �8h����U	�V���侗��3��`�e���CMA/x�z��Eel�Q4-����u&�b8�!uu�� 3C��G��%�;�ή�6��o,���!}ae��l��k9�&���]W@�mv��ȕ
(��׹��`��K�����wk��f�7(+&f�2�ϸ��$��B�x��Շz�Y�nˮ/��C�Zޚvb�89��B����1�w�}�2+ם�0���Y��j�Ѯ���c�p;�3�=����tu��w��3��$Z�M��6,�ͮ͜�Q��7(Z�I%," x>��q��ѹ;1jY:�k�ʗ�5�i������:�T�f#�o���f�q,k���]#�q����Tj1 �(RI##�=�0 B� ��Z�����[4ܰR����+��YPFJ�Fbb�2�ưP�1��T(ʂ�j��l�F�RT%�H)+XP*Me&ZH�UYuq�UEVE3,U�$RQ+	�b�m��1�J��
�e�J�l$��8������YH�*H�*�E��Qj%a1�(E �l�Lf:@Y�11	��$"�cf%d�@�D`�em�*$��%il%d����6�H�(�(����Ah���!Pm���T*)QchUUE����Vj�V"(�Y1���GZ������H��f8ԋAT�!���̸�B��	U�����"�R3)�*J*�PUB�H)RUHV���<(���<�����IH2Ƥ��ؠ�\��<'Gf�b"$܅o4�΍wh�^�]���uM
�U��Ϝ}0��5a>������U��� '�2��n+ъ�wOhAu�鮙���yܹXf�
����3���Y�̪�ɜPr[�����Y,���$nn]^P\��-ڙp�V����9�G7�eU��Zӭt�,���y2{l�>v�p���x��t�-���xsl8�G�o��Ѭ�By@���s��V�NW&�y�SY�o��z-a����ѡ��*bk�!��<��o+�Zwy֩�ֲ�ryqOCKv�o�C��f�ZS3�[펼�:�jt�Ua�pK�\�FO>Eo�<��Ք�׊���Y�R�H*Y��gwQ���*=y����TSq�j�ա�K Z7�j�����#��0��.�K����������3܊�^r��3d\b.@I��Y��ٗ�nu�ቺ{�*�BUzy�`�]Ys�� %��*�+��x�m�{�Kj^fs��c�X(N"�"�Y4�;q�Y��{�V����fԝJ��='F.˺˥S�17��+��<�0���m�YC��*����h��.M��L���2��{�����$6�eqz����ʝ'L�i������7=����{0�\�Crʋ��V
��0%��ӽV �I�\�h��Y��|�?)�7��5ʦ}G��l�Y�c}Ru{r���gy���s�)g��=����qdq͆�#���Se���+%z��w9�\���9z����d��g����k%�C��J�b]G)N7/d�Y�������+��m�1�˩}^'i[��yX6b���ĩڡ�$0���r;���KL8�-];�p���uӗ�s:���Z����I��M:�N�Pg�r�[�MeFCBqC����F�h��s��n'z��0��M��˶�������j�-��hTj�0��R�y�m�.��;E-{1`N��9��]�"�*�[Un1׵�LF�'ʛ��<�O������v@[�z!���R�Hf���qhώe)�FU�*5�>\�\E,V�c��G[�$nf�d!r^�-T��Z�e!ܛ�s:��|��K�Ɵ
�t�7�pweqwKV��$�VpѸ�"�]�k|:�a���)���]��E�-Kfu��9��˰�pY�#\��W����ì/���e�V}-���9��<��T�H8�ī6�w|4�z��9���O ����W��5�Ӿ��yu�ѣ��:�}b��*��x�)�5����+��v�1w�*�;��=�qo�ó��B������5�׸��׊�HZ9��uL�T��(��CV�QfIW]��*�ozb�*�KCθ|1�OQ�ThI�lM&�:I�0�v��_*ފ��Y���UKͨJ7��mQ�啝B(�V�+�#ĩ��wM�qW4t%;ao����w�ϫ5T�4^��Ơ�A�,Gs���D�ƒU��۔X�گF
��0�>[~���)�x)�7f璖�٥<�5�6_�r5�&)1¢esOc+t��XɌO4*ؐ�� �fs[nf�;�v�S�9�A��*"e�A9J����m��"��-Y���������Q.c�N�'Nn��,a�t��x���a�k��--��6�u��pD�F.M����EFǻڨC��m\z��\�/-֢7���\~'N;x�ϟ:G�S���u����Ӟ�;7�8�e���t��|���f�z�|��(���Μw"�2��l�i쭙� ����C����ӏ�
2��9ׯ��Uf*Ťϱ9ڧQ�&*1C�n��B6o}C[n�H��=�oL�bK��]�S�<�U��ʫOMj���W[B�T9{1$¶���v�X��}��~[���U���"�z]�(��^LF�'ʛ��T5[Y�}�@�M�ٮ��^Km�"��O��R1�ZŬٲ�nm2a$ud�"-k��!��<�X��|`�!��I��h�
o�.���D��ډ�����~y9Q���y~��Dٗ���C�����`��T4�ռ�PF�\������϶�y/sĽM�DحGm1Ե\��y�:�h�����9ҵ�}A��;�QΓϥjޯ-9��ݤ����s�3�i�o���}�E0�*�e*��P���>�k����v��=I�4i&D�C[i��s��#��З{P�PW��I��]�(���.������^:y�+�6�b���^�g-�u��YJ���u�*+/cRη�>؛��(��2`#P�TTb�p����\�������V�ܕ���U�Պ�Q�ڤ��ɽ�NS�kN�������Ιv����]�B����j��JV����g?F;�=X8-��*��P]{ɖ��,�b�Q鮖��bs��:[�i�*{�i1 ��t;���(��;���7��o78�ݝpz�6�Χp�S�s����I�/�=.���31�y�"�{|��M�\��Y;���\�;s�����B�ov�$]>��B�>-��z���E`�m�3��ڥ�7����2��d�o-�k���8ӆ�Xt�'\�]Y�^�ɜQ����ᰭ3*[�Z�)�����*5���G[:��7ƥ�G�yP��=��R�~��<�(b�S>�����L�j���	���
޳�6͍��5p�'e�Jt����*5�0�����SY����ZÊ����0���ѫ�R�Ƶ��y���(�;�ʣT�{Z�\�K���ݸ}�xI��/�^��+�o�֕����|�S^+bY�=igmc��-�9��>�uj���RaA�Wuc��ċUԩ�d����yQ;3�ik��n��J����c���.�H�W�;S��t�8k'>�i!�}/J��V -��6i�bO�_L�v�ݶ���Ѝ�sYQ���ru<딪�O+ͧ�)����-ѨTof�;���L��~׬��cH(Z�����W�T\�^�Z�Wfx�q*�w^�ܵ�]��n��1=��;�8�ߗL([
v�49��}��9�Y������Z�l��]CѸ��ݻGV4%Xz9�௮T������;쩔��y�7�!oVj�y��"����ʌ|�e�|}S��ک�Jޤ�m��gj�~-�j�NsE��{
��p�$8�yd��V��{7����D�%��ő�a��gU{�6Y��U�_+��[��i�"��L��3��w
걓�Y�ʹؕ��ř���K��˖��jy��i���-1�u/�	�Nv��`ًXL�o�lF��L:#.73m�QŲ�}
a;�p�1��/��&u@٥���ڧ�u�ڢ��.��F�ז�!D��l'��KT�`�>��hm���	L�.��Il�6��T�������>S�u�	%���<-� ����u��Gc���U���*�>W6V���Xioh�Eq۵�z�.�O�~�����ū�~��zS�t&'9���k��^R:�θ����ƙ����O#w;r�{M{\�LW�����٤�eDsÛ�lh�t�]Y���z���7����_ю��2u!*��OUw�v�����s�:��y���k��ۇ4Fd��8��*�9Z�\��|૽Ij�sm������OZݸ��>�g٫@���������욅:� F4Y۬(��J�5b����g�ꨄm+SYPO[�B�T�ݦ��)���Z�j���=��zZ�G��a�y�	�[��	��⧠��MΙ��wf.觊���-:��m۴m�*��5ԻodK�����V
���E�y~�՚�%��%���j�T�Ċ��}��5��:��a'Xx*u�����n���U��h���[���N�Y�n�f�cm�t��ҕ��.�஠:���G�;˛��)�r���S�i�L��⮿uz�ݛʲ��7R��:�x�w���g���6��daN��{R��K�J���Y�s^>Β�ԋ������B�h�Iˢ��\�hX�cWx6��m��r����%��G=>[W�YZ���[��ES˴B�Vqib�ӛ���uBxbb�*3:o������M�]��yZ��{7���3+{g�-7�S�t�Jw�x;a�8TL��')[��D���L�͉���u�%���^l|Cu��st�X�\>��B��)�R�w)�wN��^<����mS�!1��tгF�����Ϊ����@Z܇u�:�U�˜���Tdl�F�u�́o-�=�s��m������Bc���,*����۩Վ�^N�j/,h���;�^��h:�]�)�e�<�g�/k�+9}�{~+��h7"�Icկ{k��b��������}�mY���(�4g�:���]�
�r�yzxL���ſR�-���}����=�t�6�t
�����qx-�o]5@ۖ����U�}�-�»Ux��}�#I�Yن�p��J��_.�����Io ���)tţޡ����҈�]�y���:����ty9pc�ݘ�[4gz�d"�K��+��N�˝rs-���4P�E�)�+9}������4��hWE4���Z�Sʌ|�g���+�!h�/�����sv�$s��G�j!Oex�����:9����9ߌ���d��}3�xVʨ|�v����O�s����&�=���^��"�ek]��C]�/"b{h���K5o<�q���X�[8ʱ�*�	מ�uC������헪l6��ޕ����r�9�t��_V�(�R�E��a��Y�][��k�\O9�T�Lݫ��;+��}/5TNuWJ|n�U��&8TA��·7�ۯzi�N*Ƭk�^�8���r͸.���gS��R��ΨO��Lpꍊj�22��Z]y���u�n�~�>ǅ׵d�bT�1/�O��1%U��
��n�ps1.��.
���T���W�"�}1o	��z6�W�7�=ẙ�}M����w9�r��Oπ�~^딖z�'�Es�M�h^=�)�Χ���+q�V��MG���wG!=�{/��x�C�#�˧�+��p*��0WB�Lg{I��r���е��Im�^H�01u1ԙ�Qe�J|X�y�C:��֧B�-9ݗI�0#�W���)�ơ�r�.�����bC#�\u���2cV�vR���舗$fG^��z~w�V�R��yټ��Ր�X͵��R�^bt���'sp&�����=)��[B����)�͕<�f�Fod����ƽ�UP뉑O��Z�[��Uj1V��Ԃ��{�o�F~�P ��� ��\�ά��j�֩�M�^z(�wyV������������T�Լ���ߵ:~���x�]�e�kn�W��W��d�R�1<�{����f.~0o�+���'����N�q��c��P��Lu�Ur�G-O	�����w&�eY��ͷ�;{�;p�*aB�=����e�Ӎ��jW<��ʭ�������G�ޥ�q�ᒛ����hJ�B�=���Z�%uq�ta��gs�3\�+�}1��%��|�|6|����g�~�۹9ӄ �G��()N��]L>�����vj9��W��Od^l��4�;��*�0�^Rʵ�e�^q��nQ�&��Ҿ���� �t�{W��z� ��H�mZͧb}z��]b��N�������/�9B���K���ҰN�R��.�|r��1�J漲/2�]yD���m�� �``͍�&�+�����S���	��俒&j�U�ج�n<c/S	D�#Aټ�X��}����5��-��Q�(�P��c�/��h�n��o9���Y�ّ�p����.���g,!B��hZh,s�*f���M�+.������g=�#K+��[O�j뷓�����|���ؗsgT��
�˶@��k(7���u'���u�4�U�k�2�{N�o{���ug(r�m݄%�CQV�!&��ݽ�q3�Yu.��*9��lVvT���D�#l��+�X^�p=�޳Wr�r�p�=y
�`r�����d��s�"�C��q�JS���Aa���s�[٨c�E��K:��Eݳf�ꐤO��WVR�EPZv�}�ԸV��Ǎ4L���^\,b�5�K��R����g��i Q��|2*&�o&�cuEDr���8����mc� ����Ә{��%�*�$U���L֤��2��p�]��Zx��o1����(�����՝��յ�Nn]���8:7ӱ�W}� �K+q��{��h:�wAV�B��1.���I�`��~z!t9����72�Cۺ,�ow�,?�O���5$D�� 4�w`X5W�Nã��r���z;��di���M�J�:ԟu	4*��7M�{.�����o9Ǣ�@��!<��ھ����[|�����֏Sx�u�D�2Bf^8_��V�*�\��s���8�a5�)�)t������Yַ�1 �}��sv�z��!aV$K5Rh=�٘��Tx^*�A����WP�\$�.�4ګ�N}�v��h�Jv�N�9٢�_�꧝%& $X��rN�����&u�peJ��r�B�x���S`Z����*�%tȻqj���;��	 �f�.
� ��.b�C��6;װ��X�ڵmc��`֪�?�+��qq�jV��}ʊ`l�B������85�9��I�����Uc��;Gs�_;�d���-�;���U�1C��vnG{R��WY��|8����<�R9��|�t��:��흴'���S_	-np�(.��Q�GM\��V�9���]I�0��\���Z�5��X�������Wmm���� |Y�e�Ú�l�zWM�y�h����ь5@�\P]���i�5�G0I}��4n`\-�Vʫ!o1��d��-�|`�!ܗq;;j�TmJQk��}к�d�̔��<��/�7�1�4��� E ��y�7��\0E v.Ë;��%7������q���׼$G6ձ�W֮��ި�̨��y�[�P�X��tC�o�9RN�S8W� Z��c{i����n=X�j�z��ˍ�9p���ãiu�ߟ����}�������¤XE��%cl�Y�D����(���q�`E%aQ�C-	��MX�a"�YXi�U���V"�Ĩb�r�*�3"�f!�E�Q2¤�V!F["���-H���J���:d+ �Z�a��e���V+�YV"#SE#l�-J,uu��V+[dF(E4�b�&2Q Y�+U�"�"$�2��1%Hb(��������*�c�Q�,"��Y�(�T-��"�u�"��R1E��Q"�� ,��M5�[%�"�`(��ZTƲ"��e�����-��*T�

�,"�Kb�dXUm�UEX���%b 	�P�%r�E��"�UTR"���Qﶟ(��z�5;�!ڮ,m���Vѵ"����Օ���;(�A;:��X�5���˽�y��9�s��b��Ww�G��3��;N:� +;����U�PN�ʹ��}�<Sf^,Ʃz{}�Ų��蔭�h^}�뗹+�����WU��Ř��\�bQ8)T�m�����Z*^��S���X1׵/�	�W�5͍�Z�}Q��΋���Y�Ҽ�n!D�Ɛ���4�^B8D�>��ױ:��On����m�:�f'o3yV�Ӆ�L�(9-�Bc<�n4��m�du�lϷ�+�ͥ*���Y��_<��r���*���Q��b��Ш�^��BX1s�׋q�{��]{���������3򔭝��\dƤ&!Sy~OV]����MWvN�ֻ�r_�&6yZf�g���r�н�zv��-~�d���J�g;���4j���I�84��W��j�!�]��ͻ��/:d�!׳#n1�5W.Rz��U�_��z��B�Fo��a������Nlp�в�[�Sڙ��Y�!c���:ک�T��g���:?^]k��G�<{R���-#EsǊ4�l����)T�kO+}E�v ���]��ӴRp���G�96�0��ո�Nr�PK�݃5{�|�uj���W����YM�S�'�Z�OmFj��#���M��M�|�~r�������y����]�G7ɆߏWA��t��N@��G�es�����V�����r���\>1�w\�<6�gk�ρ@��}��/'�s�7^�p��?.����y=�<j�-bm����@�(W�lO�Mk`��p���ua���w�}um߱9��U9Ϝ7�z����;95<vnh������y��x\�{WY�][��n
��,�C�.��j9o?M�R��f��ቧ�]���o0�p[�M�� pP�{<о3�:���}N�
�6m�v�Lp��}D�)�m��;6��r��,e��
Ե:��"�Q�'���t��°1�`N��<B����sw=����\���=Y��i3��S��u->򫕽0#�򮞹5�S�:��y�C��Nu��Y�U���P}��u4��&�=�[���O,~�ivd��h�{�ef��I23�$�ǹal�<g/S�l�%uՄ��:�NJ�YWwn�38�]��;������w'�+�5I�_%�'#y(�Q���Y��pB�5Ύ�67�+�@3X�M��dN�����"�(0Z:���UU��GӶӚ���Uߤ+7��kgU���p�v1�@����}�������FV]1��=�1��5��B��u�}�5sO;7��ڄ��2�!~��e|��-�����W^-���#[�-o7yU���f�4�+Y�,K�ۙ��y^8�Ӹ��Q�s�����au�7�z���L�����{�iԝ{�Β��f����sU�|�w�<�|�dS{Qv"��*�w�����$к[ιR}C��L�ӝ6��k�9ߌ����}^��m�~}X�2��\{F�U�U
{*ᖚ�����\�=�:���9�B��o"���j���R�gQ�.�<���_]���J]ɅNl�ڭ�ɡ����D�>o�Q���c�1JQ�ڨ��\�IU�Q���y�/�Ƴ�y�>���]NuqO�'���Ȥ�
��O_T �[TeK`Y��4����..�b���~�o�oc��4��>��,������<���H��d����㯢�6�>ڹ]�1�k��t�j5�b&C��o�<�}çk��
�M���lk��K���w��������\��y�,��lC��meR����;�t��R�7��u���d04Li�)��X�m��['���c'Q�&6%O1.�Jt���G��Տkw���+�����_�?*�z���x�Ճ鶀�]�)���ͻ�YP';zzA�73ю!����|�9k	�&�EfUz�'k)�r�TA�s��i:��~S[^�|*5C��S\��F����s�����q�[�5Ӑ�TOm�N����ίj;-��}ׯ����Z����Ϲ���poE�s��R/Ǖ+�[U�k��Ԅ�o/�jj�7ϳ���ؑꪱ��ɗwz��y����h��YG�˵NV������N�ELNK�}ֹ-���^���!�H��f��]\�d�R�#��9%b��x�I�~��]w����c����P�����^�J��5M��kU��^�Yv���W��%���w]�k�Q��)�7�d�4��o�	�U���ƺ��C��ꏎ����2	Ҭˬ��Ԟ5cm�&�Z�a��4LrW+��ZV�v�L|��q�M&����%\�3+{�Q���K��(F�"�j�舉Q7'7���k�X����i�	��q\�*z�
���L�s���H��S�?W��/NN`�n�&��#���Еa�P��:`�Y|�l;�n�8�T#+)�Ԯ�t�Vj���\�#~|6^+��nYI���#:��n�m&�+�9�f�6���ۂ��f���Q�/x����mط�*�n6�qg&�_iqm*j��^��*k/ &Ys�^�}�}xX���q;ڔ]�32ˎ��Ց���J�v�N�SB�]�U�@��-�{0,ɕ��5
3[�-��9�p��4�d��d�u��"�i������m��[[>Q/�O#�9��K�:�!��L��.���۔\=���Z���f*�ZN8��n��18��S<��끷v@r{���j�]��B�ɹN�n)˜�OMF�Ҙ�hw�C{[�붎R5���Q�O]D���q��圫�P�U![�%���Iͥ�ς)D�BUv)�����-Y��bcrP�W ���5��u��q��5��{�k�u�5�A�C���,��+,�����]&9�p,ZĵI�k�e�H���ف"k�(�V�}�G�=�jSi�:��+l�}Ȼ�)�0o+�)�U��Q�2cR
[���˟D�ݣ�@�^�D�~�1�l���5٣>	oe�o>�nr��dH�i���"�P�$j�n�:Mk>���>�%���������0j���8�Z{�����kեuֿ=���yP�vJO���o�cg�w/)��G\^�2���:����fYʽsʹj�jyP�<��q]���v����ZٶB5jܨ��m5��)ÞȨ;h_%v�E<U��!n��ž�7t�ᖶ��w;=kE7٫���A	�RG#qU1~��ty}��Ӗ�]����oJk٪�q�9��ƙ���ƷH�{�r/�әBΪ��և]+�&뤬T��т�w�f�#�L#`l�Q���+ms3�X���~iR��r\�n6P�U�V`�ӞA�g�ͦnFk��"�ݙ�޾yC9�P����l˙�8óⓣ��޸k�3^�̀�<F�ļ��WY���F�V�]���o�5,g�g��2g�;e��h���eՌ� :���|	�A�	���Y۠3�
f��gk��ǯ�k�	}�|��.���.G�[z�q�{��؏Fmfu5"*�*���&��� H���SyU�+���un�x\���_{�����u�,O4���(f�K�b��1!3~u��72K{GD��{yz5e@���M��g���{^�oo��\��>��K1(W.]�1^f�ÅrI��΢j���Gp�*V��X��nY�0�L娬>y��%0n1HeMT��R�����I��K���{�E���t'�^k��Z�8O���U���5p
���*��W���]@.kmcL{�"@�r2�?}�x�T��I8�"���ߧ�0��]�nOZ0�]�ȼ���B�y��!�x�
��W��
�V�q��E��9����\�R�m�&��W�Co5m�載Sz����k��F2���)"�)V/��F���]'L�K�΍�jY�P�ˉ��k��#���^�'>�����g���h�/NzۯW���T���QjL��&"&�W+{��V2�U��8${*x0����n5Ϟ�Ȁ�ۦ�R8�a<�!��
A{�I+��r��ؘ���®���)�᮵{C]�AX��Lbt������;��w���z�Z�NM�W����k�M,d��f�%8+!N�B}�Y0p��,to]��J�tRg��6��s0p�.]JYIh��1�7�.ɗ��-տ�SOA�����q}�����t����iݴ`O�7��
��6K�?�G���ε���V����T�Bw0��D�gd�7�*�Q
z���++���,F\FJ^�eD�{�g{.y�� �N�p����#^���g�%����5�ŁG��(xm�2�K��}{�:v�cTǫ6X؊Ɇ*#��
q��ױ�jUH�a�Xz�BzkmN��#����2z��6���x��6�~ڍ׃�ka���~D�c�yX!>�#J5�6���wġ�y�����tG
���=���v�e��$z����GLu/�擜u���7c��ֲ�Z�$7�������:1 �Uqj�l�<��j׷=���m&+G���rri�?j6{�+{���b��o�j�-�LSr��Oȓ��qj���b�	�a+�����̗�R��^�v([�(?9Ǳ�����j��#֥y����a�Ed������&V��pxml�n�6�� �8 ���L\vJ�#a�؉�*p�l���z�.�Q��K����s�<��c���5}03���M�q�Q�C���ED-�"9�Ƚ,D�0�+��0�z�5Bwc��!P�tݮ�c
�0k�޽��� ��NE{X�wQ��u�̦�H��5�	i�U���A�=/H8(�K� V��,��w�(�+��T�^ǵ"�>��B�?�S�o���s��ne+�#��~��=�����Jy�������sj�\QZb��0��sQ�PD�B0��p��6v;�����ƻ��58����]h���A��pu�K�X��͋���b�pO&�O��\�5f.�{zy +��k[��
cx��1=f�NRq�݉I-����c|)֞ٜ8'@]��=���ϐJlS?y}=��0��]�~��vx�F�J�
���D\I�ɱȣd�mMot����T�F���Û�a��<"��c9:cT��8�DZ�(ï�8�{b|4� �c"畴��Ÿҝ34KF8v\eB�Q���cx�-���0T&�؁nd.%��Pj�� W�D�^Fg9ɾ���� /h<3'	c�Ni�Mf�+�K���'	�xo-vHk2�E7�Q~]�.SR�;�+G��և�\Ub�|jF���:����cU:�%Z�^�X��s[7�qm�;��mv����8���h�:뼨!\T��b���Q�,>9=��V���ZZC���7�_��֝�i�D̘��UC�ZvJ a�b����_P�uׅ%�i��O9֤N��\7(��pu��l����	r�k�l+����u�]�CX�(#z�#���Κ5'1�{mg2�z�`v����V���6:ɵ�r��N���~�ca9�~L��,U��]�t�[O����:'�27*n:Һ�4Z�G��#Y&s��t�H��{xM��Ģ��D0�=#��v��F�:#�UO<���J�����W��ݜ��5�l%�~�R��,��T���bʘGV9�;IDS,Vvӽ���ig+� z��"�e�
I�Sc)��3��2��P�f,<E4Y���1��¦�Z�S�B�_N��ZE��q�����ٔ��㌢o��N7yN��Z�9��M>�5ժ-z���xn��ǹ{T��v���`�"϶�UZ�q!�K#Ѱ�)2�P����3Y.�
���=�ԪWv3�� �96�����ҿ㣬j�[�9�o}H_�ȧ����(>�^��R��wÆ�3�S�gm�b�����i⧈Eٛ㢈�W:���R����P�P�qJP`�����;��6`q��+��t)�u]K�.[\�D
5`�-yU�9l��T��>��N��r��)I�~v�e�s�e䬧���Ҳ�1w�b�62��Cb���t[��q[Ҵ���C�8=�x�A�e��	m�Ȓ�c��c7 @���t^_�T�c�ևe=C`5��4,u�j��&��������C��vn�<Hx����ѷ��˫nZ�������]���A�X�v9����n�b�F3�Yg2*mC��X�� �U�9�{A6��V�ԃ�o�LΡ�A����Q��,��v��B�Ы����V�m�&e�f��,��^|��`�`dT�g�E��`�7&q��Z �/Zܡ��.£S�]�w0Z�����D*X���B:��RR.�v��NM�]���N�HV:���wV]̬|������u�C��U)Y6��5싒���_,M�%ʘ����4.�fm��m=�{�S�'[#��y�j�ܱ��WH�+C��9oU����vn������=�o�E42��Wh���0���F!�@�p-����Qƌw�"���[�t��򡂥��a���k�\�,�i�vv�l��2�@#g->G������e�l_L�xAN�^��.��Z�V<�k�v���,]t:�Ӎ,�y/�doM���ArV�Q%up�M�00rګ{ݖ��߮��`�08�㔄u=��x�'��}.HKc'��yggb�Kt��k)��>��z��Qw]�I[Q>Ђ�ik��WˍrÓ{��_+�c`k��9��b�`+�]�q�r�s�gt�a^�7�9]�7��]MJ��{j�6�X�+��h�z�^��h�C�]������g0�,V�x�.x�mv&���V�J�]�]���[����!xD!gg&o8�1��<�M	_t+���ޭ�،-\\f�헲�	!��U�����DxgJ�������y*2��y���m���;�U
�6�H�9��.��ip�^�g\w������(�:T��XB�O2��i�e�l+�[+s4:�o,*����530�l�|�%Nn��J�.{�u����=]\���TtV���IS����7��t8�1�[�$-�Vf�3r�Y��c�؁�J�3�i��W���"G��R�7�&���қ6w��C��w%R�v)�1���;�V�r�uWF�qtZ��v�k����pmp]�h49���n.�/�v9�E4V�)�/�P��;��r�u��]�U�dI��]���|;k.��G����rzMfn�^�v�EtJ�Abm[�ϕ�5_nMo�oe�e\U.}��e2�D�qn9�5,"�,�[�ߧ�sSǃ��q��'=�Oq�]{C����`9L�Y_�^�4Vfغjn,�*�;㻈�7�b�n���Q�Iv��Y��wN�w��#5�9bT�N%.k��o�]�}�(Q�JF�����n�L��,|�T�.HE�sW4��V�<����l���
��`���5��GV-�9o��CO19��>n
�&�/{���9v��\��Ը��V��s9]Cg�66wp�w�3tj7��(	Ԓ�  "< z<���b�т��>�&0D�5iE�1�b�)*Tr����(*�f�� (�� �"AdIXV*��a�1`�I�F#YR[�+	�Cƈ ��
��E"�E`�1�Ƞ�(i%@�VZ����"�,Qj�d*c��`"�m�%�(�R"ńb��+�UT`�TV�X��+H"(�� +l�VR
1�CV���,PX�R�dmAb����H��,F��(����*�I\E*)R����Vc����Xc
��hJ���(*�UcY-�H�"[H�VT�
�QDQ�dFҮ[*�(c(��b��ň�V)QkUB3-Dt�$ȶ��QA~X������ר���ͻC��� K�	#�e�tF��Q`�.}1�:�e.�2eNH��N�Jn�gk.͹R�B�_�����V*]�5�l�!�&_�l���r��<l����"���y�t��|ks�eG����/�N�����u/9�{���"�^K�U��Z��x����WF��d�e�,�����*�a�m��8鞮N:���r瑕�j�F;�J����-��+�YY&E�=5*l�4�f�ms�}�̱u�s!:NGR�������LRtx���:�ۆ5p�v����.%�u�oTγ>�0�vtvD���5��yS�LHL�:�b��I,1���M "�n]]�W��zքL�����=�Ξ���.kK�2�{��.�ʼ�C7F.�ࡆ���Q8��r���K�$��L�hic�	_nY�0�gEn/���ε"{��*�.=ǫ(�^�'�[����u3�R�+׮�(�G��\��mX�5K��a��}�yJN&G��h�z�����~w8ɸ�t���p�l���1:���9:!| �t?@��ܱ}�pOk�Ҍ� U�:Ѣ���i������ռh\.޹���zp�ڮ�k.��z�tf���p���ڷ�ۘ�vKPDyR�7gf��Nu8�f��?^�g���K*pk@Lg���iu�J�r���u-´�7j�θ�E9]���WdQ-�@rcr�{��ڨ����B~V�k}�l��{�@(�%ȣ�U�l���ox[u6YC�������{����%>�n�J��@��j-O�l�1��T�H��J�!m�F��='�mOz��O"�d�K��N�e�e��>�u�qS8S$G#Ѫ�ՎV�y�-��AQe,����*��ɮ�$T-w`���9�H㫭2�����O�XS�~�>z�s��!�����W8$'�exO���G��
�|��ҹ��>��ǉ���qWz����q����c���uɕ&C�BwzZ>�-�ø�e���)M�U�SՄ��Y\N"�_\��9���Mr����h��xߑx���F��x=~g�%q��B�;W���U;Sp��{]��������C�Y����a��난u j8�H�T�DC)�%��d5�0YV��y��E��i�ys�f�O��L �;j���=*X�9=���C�,.:�_n��x�+�!3�͝�E�VIy�'ke�9'�1���ɣ�k�o{�J�|���M��}�>�e�K�xq:J^Z.�$�	^80WJje�,G�W�(Re4����]	�)8��s��`��F�j�[<��1n�Y���J��.��V�}�* r3fv�ܒ�$ݚ��{��^����Vk��s��͔�^�4�j`�VmE}�2)�Γ�K����y�q��<���![l�\l�_<��6���X����̍I����6�-���?������sxn2����>���򜚇�h������bgn����(`�LE��2+{D��WA����V�"�+�4�Ƕ1H��]���gg&-�%dߝO�5��z�c&����o��I�:����[��X�� ��L_�%y���lR�7��l�(�����߹h�C��ŭ�JY5]G8��6�s��Ѓ'�2�B�O	r����X4�T;)�.�;�r)8F��\����V"�E�+�΂�&Q��ju)�W��ԡ, ��v��~���k:��� ��P��+v3�hgԳ\ּ>���|�����OR�Y>eN3�����*O[���}���_P{�^Q��Q;�;1b��߳�i+��}tΓ�d�AH�!��0��=H)�'���O�b����� ]P�<C��a=v��PSúރl���3.'��$���0�
#�G\Ǭz!�" ���ɵa��T��Gs9��߽����_R,�'�!�J��������i�I��X{�
IY�6k�|�� ��|��?0�c�AO�L�IR|͸�|����xs_h����Vb%C��c7w��:W����w���۷����~�N'x�C��wx`~k'����V��Èi�5"�?YY�:§�X|�Ou
��<��uS�
�RT����0*�>�ig��gs"�@���N��Rʷ�=�ڛQ7ڻ�F�}�h��@gC/�=�'��x{CXq�:���H)�O�v�_P��C�������$���+��P{a�~Ͳc+'����m'P�}s'��L�%C��_}󥠓�f�C�>���M��Ř��*�ik=ټF�����u�L�9��w���������@��ѣ����L�_n�kzض��[�?�{<��'��O�H�-����=��Xkw�u_B���dKB�#�1Wr_u�#%іLb㷧TFU�����G�6f��9����&�c6�>d���Ѣ'̩��I㉈�z�&�>���)�q%~d��ԅH/��n���� ���v��P6}�봇ևHc�~�+���j��/(Y�;~�k��VoЄG��eI�,Ӥ��a�8Η1`u�8¦��EI�����}`VNy�<I^� n�	�+>I럩��Vu8����
%O~N�H<|<�f�~��;�>z�Η'e����U1Sl������u;�=Oj��0�J���c���'Xq���s���0:�M�<�Sl\IX�7�I���T�a�c����<�a��B��)$�{�k�ݻ�Kw��=���!=IӔ<a�6����3�9�'������zɉP���'T�2��ְ�&���l���k�'�0�&��@0z#{sbw蘼�ZA?^�b��D�"#iP���'Y<Mˤ�����*l?Xu+�m����9��4�8Ρ�w�bAd�-�d��+<�2u�2}�釾o!�:��d�Y��|H,z 2�>�Kʅ���6��LV���p�H)ǧ�M~����q!��<t��Xk�l4�d�*��t�ΰĝ|>�M�+Xu��T�6�jxg0�E�
�A߰����>���h��)7�<���C"���}���+>I�:ol���J���'���
OM������H{LN�T��q״:H-f��S�Z��h(J�Y��y�$�:�M��z�!�*�"��6�K�?Mh�����;��>C��J��(�������jLea�
�xw��:�a��;O�!���~q�}�*g��O�������C\�u+��LCԝ�N>� ���nJ�T�j��8�N2��@�`���6�ͤ��ܟ�c�`<�1E�1?wY%t��T79��&�4�ɹ�2i=ObO���d�O�g��<��I����gS�$O���O��X��Md�f������ޱ"$D�M���'��3�{�i�W�<9O_�
���O�?:M$Ü���O�1C��Ƥ<�?'����x��X5�i&Ь�eO7dӤ��a�=�>�v�2U��I��+~�P����rj�OV�~�T�W1����-EWy�(���o9�+��zk�; �����$�ql��r����WW*i TQ�:�/[��_ɳ���z��!���2��ԲoB�D��2�up�vNN6'(���ur����Jc&r�|;�!�ma�?��I�6��kH�eH�\��4�W����~B��<��u��B��J�Sğ9�Af�q"�����NC���z�R~g���G�4�2�+���.�_��{�1�8���6����T8�5f�
~a����Hc�Xu�b����v�Βq
Ϛ�r�d�+��k�>�@�'�+=;�>C���
�g�d�!"ǽ�T!q@End}؎�:������R(q�3��֠)�f˙:�yd�WxyC�'r���WI�Z�>����H)��Î�u�d��a] (���Nw<`u����s�<G�ǈ�g}���5]ԓ�\ZC���\�����#P�H�pl���"�m���$ĕ�q��7��؂�a�����xe�!S�������J���C��Ă��!^$���`|s�i1���R��9���[�S2�[�u����"Dz1Gk����u���X~v���d�ِ1��q�'����a�.��1=LI��x�"�ʑ���b$�_dRq
���ݞ��HT8���7�^;s�7���>��?$�ީ��ȤS�'!�;�I�&���Oký�;gP�i�ƥ���(q*{��+6�S�<;��O���0:�Y<eb�%OfY8�'�V~k�5���;����ޛ����C~�1�`���L�"$�syP��g�7�I�>a�0�;�PR(~g����@�����y�'�\Cٮ�4�Rs)<��jWi��7�LĂ�����VtO'SHgH����;�{FE�"$D}||�E��5i��Xi+'YY�C�T�6�}��4��������%IY�/p���7�f�>q1���q
�2g���wm�����ښ��9������<Gg|���Ă��&>$���&�l���'�̸��RZl�E6��k��:�6�d�3"�Ƨ��;��6��Y�����I�1�a���/@�؛��6�2�����R�uWd^2��Ld�*I^�^��q
�C�}�~|���q?yCL���`oۈ)��'];�'P*�E�t��Y7��阇SL���AAC�({��g2_�!��� %*�*Ǜ�v6)��6]��3������#ײ$}M��qR�'K�����4�x/#b8j1t����s��s��.�,�v[��S&GY|;q�
��v�m��K��-��@1��
,�n��W+s_Dze;1R�ض#�Q�ΧWh�W���G��x���V�9���z��G�&��O�11d�~��&2�|Iwː:ԟ!Y�ֿkiN2��5��$�~�SL?!���3�1�i�I��&�R(u4~�fՀ���ﾭ��΁�e}@���_}��=""l�m+���`B��P�{���� �����֤��bC���a���sy%t����s�B�:�ƽ�H>RVN2����i=Oc=g�N���yAJyٕa��=�E�W�k�}�DX�ԕ%N���<d�
E��O��'�&'����J�N����߯���Ϳ�4�t�S���H�'���L@�Rz�5�`cR�&���-�����Q5Y��[��"�@`+�����=g���6��V���Xi:����x�"��7��i��T8������1&Я>��>w�B�����4����;s��S�G�	,���^��X�J����aI��@�*t�3n�5%�\g�q4ɿ)�I��k��1 ���8�!��1�ܡ�L�eb���M0<jN!^���H�z��~��O�J�+�{�_�3�R�	ү�������4��'̝����T?0돥��R(_l��V�a�c1�!��u>ֲ�>I̦�P�6� ����뤜}f2y�1>d�:�C=�wP:؈� ����l�#^�5���?Om���ϻ����kyg��RVOϟSL�ʟ�i1�,<CL�'�3�ߚ�h~IRfY�L�,=��O�S��q�۴$�
�Jß�$8Ϗ�i����CUk��x��@�zoU�e����4��t����v^`:�Xo\ϟ�8�Ok'�������a��t��B�g5��m�Z�g���P�'�*��t��:��'�:AH�M�.�,�eC��Ǻ��?k9����9��o���z>�@Ğ2�<I�R���&�ԟ��CӼ�i"��o;��H)�f�N3`q�P1�q&�}�`q�AAC|��6���bA��8��m��{tr߼��|�~����~���߼��z�ɶV/��`zԟ�i���O�^��a����B����'P���CT?0��;0*
E;i�u��>N_�M3�3�O'���� �ĝ����}��O���i<�*��wCޫ�39�w�%]
�:{y�;L����]�J2;����W�\�n�xvT�rg�� ��}E�P^5��8�w����6�5�GI�����A=��Ԣ0K<7Rr^[n��:�ܻ9I9�#�yʻ��T^�B��P��%�ޏG����OV�����'��
!��5'��c2��'a����M�:�����l5�n���i*M��gY�O�S��;�)*�����Y6�$�l�m�|f�(���_���<��g���?k3}�����Y<eO̝�~��*N!S��?jO�|H(}�M>�q��ɖb
E�'�����8�{M�P���a�X{�'�b����:��/���Ͱ+S���z�ߏ�ϱ��_8g�y�����?0�1
�����§Sxf�l5"�w?jT�'YP��~�}t��8��c��߮��JΤ���{5@��x�O�S��
u���i'�ی��Z�;ο�3�:��n�W�=P���C�;���w�=M��c1p�§Xc1��f��u�'̬�Zֶ��8Ԟ��
��H�q4�����1��Èi��4�u<�ԚC�*���������n�s���������PXvv�3��S��4ٶq퇧w����AC��/2~�&3H=�0�I��c1��Y?8��~׈x��P.��0���OR������ϯ��6�k|�-��~~�]}���2xʚM'�O�����<ͳ�J�RW��2�gY(��y�i���Xl�p��<@�:�Nfi?2kۤ��w�T�q����wV��x�����F$��~s^��fh�;��>�oW��8xDp#�=�2���1'Kg�`q�)���4��Vk�u��u
��<q�T�bp��0+PXw��l�M2��wRm��!���(i���>�{���mD�������wU|.�bAk����<�8�9�PR)�=�~O_
q��a���n l���Ak=C����R0�q%C��bMϨbxì�8���V�d�+���i�%`i�-��um�M�W}i�׊���= ���y��l4§��zw3i1
��>q<���6��T75�C��Ag���?3��++<C9O�����?>e�-'� q*�'_�5��?G,"k>��B��z,B�q�����`~jO>�"��0��9��@�TRWú�zͲzʟ�ӛ�D�&�����>v�*a���&���u������d��8͟�q�m*�����N�_����*V�u�Y���Y6͵��N�h|�H2��ěÞ����x�G�6 �����%-��]R�q��S����P��ڧט�L�-�����垼�aQ����9������u�����lI��ۼ�;��Ԇ�p���., s�m��_UW�T}x���|��?'������I_̝}t�<�I���7;�8�OR
~Iܣ�'�1`~k�,�?&��s��z�Ơ����d����f��z�q
���L8§S��ow�����5s��������O���2���Y?'On��%z�����!�q'�9a��
IY�7�a�ﴂ�����?0�c�AO�s�%I�6��Xv�Z�!��}���˩җ��s|�����<J���c:vɉ���q=�0:�N�ܺb�IXk��CL��6s�J�0�
��a�ٴ�B���k���C�*y�a�>:`T��_SH}�� W�T��s�*��_�;���~�ا���C9�ړĮ�;2�I��8�q'�TjN>?Oi���d��~P���:�<9CC��I�~�] ~J��;�m�Y=eM�w�=I�N�P�x/s�ٳ�N��}�{�����>t�2T8Η�4���O�"��T���x�ba���4�2}���S�J����^����~M���<H)�<�v��P����b=��"�D��c����/�߱��{�+��P��a�+&�Rw��۴�4�q��Łְ�
����&�j{�E��"��b��W��=�XN!Y�O\�OMP4�Vu6r��a�@ Dwի���묕Dv}���'�O$���6�����z� ��O�������)�(T�|�f?�w i:Ì��
�0:�OǞ{��.$�y��O���Xq������>���k_p�7ݿ��sS+~��<B��:v����P�M���q�Y�\H��u��}�d4��VV|��7�I\H/�9��.�8�q��I�5&��~׌� �Y.�fF�=�5��"�Jv%�Y��잢�t���ΐ>J���e�'YY<M~�J�I�:�M���WL�%C����T�ggP���lAH�u���WI��w�:��>�t�r��B#�!�z�_����x�,խ"�����=H)���_�1�)5<����M3~ݰ8�Z�S��eC����&3�1'_�f��:��ܩ�m&0:���a��Yn����|?+�
�����vض�z�"sf�˶Ib�ϝ4���.z�|{#m�Gv�;�˵�*��w#�(.�t4��9C�q@M��6�ٌ7Ũ��2�qݎ�H���=��r:v��޽��`"-��
�"�Ռ��-m�qQXaZ�߽�DGL�]u�o�w�G�$�'5�i8�gR~sٽ��C�+.}��甂��B��<N�@��1:�Rc1�G�:H-f��S�Z�AAC�P�1<��AJ�>�쿧�O迅�.��ו�vT�"�z��P��'��/�+&�߰]$�+?5&��jLea�
�w_��u
�=���z�P��SH~a�����H��z�T�?Y1:�YY����,�������1�efoK�+w�s�ě�O�=;�Aaơ��a���$��Oό1��0<��X�������%qiP}���l�ed޼ɤ�<I�>C��d�O�g��<����=�G��7�?�T[���z��`��d����x��g�O�u�����;�i�W�<�a�󤂂�S~t�H/����O�1C��Ƥ<�?'�o��5��{�AM��1�!���4�_LODԥ܆��Hb)�a�8��0?5����4�M���ϵ��^2�Y�P��C�+��o�I��a�{�|���|����=I�yˉ����s(bx�Rh�*J��|*�&�o�%���=���٭d���C�)1���o���AO�q<�]�����S��f����6v�Βq
Ϛ�r�d�+��k�>�@�'�+=��!���\�>SI<��z���5}i�}���<x��'y�i"����|���
z�Y��>C<�q+�<�P�>I̤�<�y���í~a��4�S���;a������WH
(z���;�0:�"8A��g�;�vn*oFk�ߡ##ӌ�=�x�'I1'�9f�18�6�z�bJ�8͜�ړb
E�N3l�8��ܢ��*u���>��W�o�>$��1�O�ɧ�r���=���ͤ�>��D��4c��)�߲J�!���P�ֲ{�a��
b��f@Ƨ��N��m�ְs�'��1���H)�T��2N3H|��}}Y�H#�z�>e}1?�X�7��=�[���1� 8�wM3�O��_'3"�O�>N�C����bI���S�����;�Ӷu&�j_�������R�i8����S�?&!����I�+�<D-��W�q����s��
�ȕ]�s�޷Biq�X��9�e��(T�F�-��9��I:��{Q2"s�C�=�O�.�U()�}�w�����.�+,Z:��1.��b"/hg�=}����Im6E��.�n��e#)bp�7&$js�!.jd�F'���W���@�M���<����y��'�Ğ!Y�_�VN2���̢���bN�ua�:N�V~9��M��8��
��C�q������)�q���W���4�Rs)<���J� �����r��#6�u��3SB=���G��>�
���t�:@QC��xe�`u�&����VN��C�T�4�z}��d�u�i���C�J���>K�=d�"�o�f�>q1��זvG�aJ������|��#�"�=��߷�AC����O�;H(?o	��1�4��*u����\`q�-7?QM����q4�d�3"�Ƨ�ӻ�=Cl����|p�9�緺�������Oq4��w����)��lְ�'YP�%s=͠m'��;��'�ϩ
�hc=I�ڰ>��R)�N�w����C_��N�k&���t�C��y�����y�����%�[9����" ��G=S�{D��$E��8�g��^�;��q�zLףg̕�(Ȟ2x��X�oz_��-���z˿Z8��r	�7
������U�\;1��W�Nnh�񾾼2���T�E{�Z&�5P�gdU�[;1h�^�$���SPEa}]�zi�^�j*G=��ufÏ^�P� _n�*9K&��������ռh\B��p���Nv��8y������J��/��$T�R �����tc/U"k�K����F��gq�w��������d��3��83K�4|3��=S8Sș�֪�c*��E��S7O(\�����]ҁ-^n�Z9 ��
��D�!n��9m�r�E�ތֵ	wΠ��R��reeA�
��y}uӦlR)���/�����*N��}z�x��S�P��;S���@k!�
ٺ+qWBZg~���]��֡���vF���#��S�*�F�L�f��}��Q�5-#�1-8�_h_n8�4僖1*u&�an.��h1[�T�aw4t�]��՘�5�����V,��I77+iR��!�Z(V%O�|Vҫ���,�ܮWaT�v�Ֆ/)l�Ȓn�^J��a�[#6���&��op-�%	�m�o7i�Wrn��8r�_)u�f"N�om���5��:����%�1ʷ,��5�k��e�ڏ'X:mf��y�0�����\�er��=KkAc��KꋀJRެ%�$�u�ؘ�"����q���/wf��\Ť,��ns;�אS"9�k�WX��P�7O6;���/���ͮR���Vk)��9-nd���*Xb��;L�����ȴgK��D�m0�V�gɬp�r�<Bl���eqD;6��FR냍 r2��r��x�;��tݕ�X���`G'_c��y���͊(&5�9n��0]K��u��0�R�w3��aG�R��{+aۮm��u�7�����vhwiJɯ���\���bqjz��]�\�v�2C�k�W=؈�a\�!d�NE�H`����XpJsF;�ѳ�n����s��,l�G8-Ԩ͏x_jU��M*7R�N��͓5KS'D��N�MZ{�oe:��L�K�������x��1�Pd�kyLq�(�h�냉����͍�
V�-Ϸ�<M��9�$�f����/+XٶmL}�>�s� X����Bn�[��W���ҹX	�d\�g5�oep�w,;�f��+�0*��I�YU��c��5�F��U𚭫��f�����u�v�[|�z�����	R�����W*(�ř}� ��V��%�6��C��z�E�TڴՇ9�s�!vsc�3���U�=�	�ZݮPQ�N�v��]�s�C�t�w�R���]h��H�tk/i��7R���t��9�Y�{�j6���)R��X�0��N�D��z��N����j`:�5�]���z�r���۬W��!��60�9z������č�=Xی�ݨ�Q��y`����*=e
Vw-��ƺb(�vw];�a���x
�Rq�*򶱌#��C��&n`n�c|��+�ƆS��=���gYHv��Zy}u:u�bz�Ҋj6��ki�lq�:)v��̝.�o�9�<z�<�W��^���5D�i���6�d�m�q1�bk2��y��D��:�x��,�i)j� qM��tq�S��l)]��奭T۱؎�p����!��m�ss�����a���dtV�����R5��D�·�J�*I��;X�d���dH!]�"�:�H
�J� � ��wkQ���QTPR+�V�)����X�
(("(*���UX�Ȣ�\�AX"�[PKn��AX��JȤPPDE�H"EY��E,`�r�mq)�Q�b��(��A���0b@�F"j�b�(�QH�����ȍB�,�+3Y��,Y-b2��A@���EAc1�EUeXQF((bTm*:��PFEb�D��+�E,��X��*[Q�E�D�.Z*��* �Q�1`��VE*T���QUQm�E��WM����.Z������j*[(�h� �Ԩ��Q*QQX�UTU��Q�0H�X,W8� ����԰TU��c�"#U�TTF*��SL�(�(�P���FG���݇��jIK���J�y��\ep�Ơ�}�oe�R
���\k3�b;a\�gu��p��ΡG ��[+{�G�=ھ�ۅ���ݺ����A�H�=�9I�WZ."eV\Q���<��rB��܉w���ܱ��\ڕ�Z��'Fy11A -�Uע�*p2n1O����.�;H��cn8ks���O
��/zr�m�a�3�.�JYS�vl��6�M\��KXbb�;u���9d�'(Fac���9�7���>�6����f��%p�^@�[����Bb�w��1~&�Y�~��dF����B�a��N�)�P��䂰5p�g�̸Vս�G�yH��^��B[��Q����u���A׻j�,�����^��������sg��P؞�`���24����
�u�G�����A�I��0؍�%
�H�qId+66����TByRL ��v�����B�!I�p�)�,t
@y��6�sUe��,��{�F(2!ƞ'�^�T�ǳP�,�L6@Vwꟑ�L���S��Mlw��(̍��ʻDHkgD�De0뮬!jD��R���<�gg&.VK��z�����F �gL�ܸ!:��+��J����wA����"b��,q��`����AWb�е,v��m��9�m�[�{�Z�� g��
H�\"ch=�<IT��5���7YI_2�}s�Ӵy�`�Sv��� �N���ĿDG��#j.�,N�#|e]ƌ���a �@�S�/ݒ�7����ٱ+�T�%glL<ז*kvw��"�`$l�j�T/#�ʊ��9P�(��Mq�Q�C��.A��w����n̰��m�^萙���ykAҖ����Ŏ��uEMVq�a���W���>ޤ�V��3�z��a.���\%y[��\�A�K)�g¥Y�p�����N\��9�=&���|+j�7sqj|�ɭ��s�ց�{�e![�RKl�2=�:������b�U\"����g|�PRa�=��֢j/�������_���i���'c�q&�a��#*��L`�Y��T-�vw��ʤ��M�U���Ŭ����Rb�pR�)ݱ�����z����ٍ����K�I2�6�T�����Y�M�u��
,�:ᙈA��B��\��I��k�瘬�o6b��O�^7ٙ�뛨;>�д?�:���+<�L\��c+�1a�	C�����w}��G�Ny?&a��j�n{_��|&�����\�k�_�ǎ[��ۣ��}���+Q/5���XM@ |,����RҾ�@��K����Auw]��WH�W���1�:���1���}w�u+�6�Q{�r�u�����$�j8�Y���������	k�8��I�s\�Мƫ���j`%���I�荔�7�n]���ѕ9's+��H�~R¥:��&0ɰ5'{&*���ULp�s�p�[�eF¨oC���^�ra�Q��b�#B�"��sA�BQnf!�.�װ@�6s�g��	��ޗ'd%\�MV��+���iC�V�x1Hp�O���U�E����xÛ���ݑ��p� qlIٖ8t�Sgo3�s� ���S�"f�u�.�'3D��m���y�C���J�6��u"4?$F�<�xO�+����5c�YY���g�Kb�|��.�,��!/on*��8g�<>�]y���@�ܪ���V��-7��	<DQ��#'�)�*�f��u��a����'11®�<6@������gs�4ŏ|��2�R���Dl��LwK2��W֍oLé��j�\�o��+-�+�fw>ނ��1�8���Y�eTr�u*1Q�,-<�R��]����3$�+�2�-v���f�쓳���A��A.[�sͫI� p�� ��S*����DsU�����|^T�˽ ��w�N}��WlN�e�V9	a*�w�J�]��]++qb��Y{�(8�Ս�c$��� ֍GB��o���B5t��}��o�`i��3��p�cx6����>���k�>�0_��-���v�����ݼU�]zp0�ʓ��B���c�����5d{:��Q��z댕�m�-l�+w<��(צ+����;PB�$${�UE��}�3����[5~�N�0{C��K�F�nleF�oL1��*I/�\7:�P��B�xT+w�����
2DUin�w�B82�����
��+��Fsŏj�w�&)R��hܾ8�^����%�W�{�){�cÂ����j߆K��fb��Qԩ�iր��<1M�p��/e���sb����j�+g��ǘg�3j���D�
���<�=+� ���`͗f�\���׋9%��v�I:8}�*�^'�\�/�^����ug�>O��RU:��O��\�g�<1?k�pB�����4�@��¦v��6�ʋ���WJQJ��8�J�F��s�w����ul�/�"����X4s\�{��������XAz"���Z7�p��t�'j��(/w(F.�Q�5�����rM���ޡ��%�5��nP�������b�Z��N��]�ó�W/Cn'���O�p�s�����|̊�ϻ[{���{\����dU�h.�+Ao��](����m���<;ǟQ��:����NN���|�X�/{Št~��h/ ��yx��sν�):�;W1|}ziL��a5@h��"�(;�mk]r��
�
F$d[�1��Y5
��Tr��V�k�����!d�9�N�r�m�s�ssf��&"�=Q ��!c�G��Ѫ�5���C�u�u�'6�H9��,��Z�y���y]&�ԅ~�gi�	���ͯu�L�o'܌��F��O�C���+cC��ny���9��}ۗ,]Wv�#eZ�e5�C�X�S63��j�m`\�o�_A)�M+��٥�"��Y7���~!��{�ʓ�&0��\��_sق|�&��=�Z����	�8��x���
b�qZ_DC��]�}�����LW��Jn��P�o�P�᷵3_B��9�*����;FxmE��G9�7��מ�^m^[6ϕ�o�AB�n����ԍ��Ǫ�>�MB`�@�>�X�)oD~U���J�u h���y])v����:�U�o�n��;��0�0���/v�eN<��}YPfu�u�gYwu��3�r��=���u��Y2T�&$���|�n�\�IZ"������+bu���Y]L��k:;�b6w� F(E��g#�B�a��B�VۦmDe�g:^pRx_S�wI�8����Eǀa�n�WP�r>/�����Dn�>B��Y������Qw���kq:���}�@6l(��K|>uゼv�����^��~����"嚲H�YZ�(��d�q
��8�k���8d�5U:)��B�΍��@l��\�S���{�����a(^���hD�d��G*�^Cڇ^
����S�7鞻�\���O5��j2خ׉
�O0BjpL�R���
D��R�O.��gd�4$��)q1�_3w9�B��"p� r��nm�A�3(1�鋎(3Z�lЉxoL���\���շ4\>�!W����/.���2�H�\�1f��xў�Ƹ��FM�R���9(���t��^הDTrʑ��"�Z�t��)a��t>��Y~�s2��
`�ֻO5Q7Vr���4����n <銇�Mrʑ_��`��98P릕�
�N�fQ$�	�Kky�s�5��~S��@���#尚܍f3���QYHEǜ�XNL��˻w�K���Zj��Y����<#G��A�>���u��̈�5��pb:Mɪ��G�|��t�qu�vt�"����&����r@2fvk�J��U�* �y��,�
P�]���OCIKB�&M���t��d��e��\�ɲ��mcCd�
	��X�u/0�L��D0/�(}�v���#���v@�~x��������>������l~�$�L��F%�;���n��U��xS����;c��sqs���T�����U����v�D8jJ1^fҮˋ���&�0��q�{QQ�3MG`�!���
�^�ޫ�u��88�Yl`8H���<y�����E7��TF�t�Vm�VLn�9�B=}�0�lu����a�	��xT=�)��%d�:+����Vbú�8l;�Uk��<�UY+[GMov�F'1��G��]�$W�LĆ~~�Qhg��ab��_���3�m�,��b�������)�lZ���[��9:�1���M�T���q��mj�.r�k]�ܣ�vLUo��!s"��sA�BQv��Av(��Yѕ�X�hN��r�2J	ĝ��s��
�l��!���0立�m�_dU��Mvm�]t6Mv`�dW<r�������z
�zZ�j�)�.L��劯��]������	�oJ]g�J�����"4:�H�y�����]�,W����X�f��Y��tH,�r-�K���Sh)��ٔ�{s9Uī��㒘}�(�^�4=�>�J2p� ��z�~|N浏b���|�W}��a=X"�Pb�3�J�B��]�9��D��V�w��TpT�.�����L���r_ls�U}�Yom]�{�x�U|x[(���'�on)�f�P��a~Ah�\��a�w:S&�S���Ro�{�1=܅����b�t��g�ٳ�[9�1mm1lō]|7�V��R3M,��C�S8_�g�c�u����ϸD�K2-^�����zf��[]vU��������pC�9��7�x\5�έ�ޟk�i�~U�Z<%)A���h:�R.k_I�V�����v@�i�Y�ل��ڔ#	�ZL�e���Trڅ~�OI7c�<i���ܺ����ϻ+cE�T�B�NR���;��k�[Q�2p��YC�ĺ�k��皮�+lߚ9�V�zlsYHw��[>V��'�a�H,=i��O�l�'Z�̍h��o�vu�5�N�]/zb����DM�w��@q�;'���!���#dM[����L�Tΐ��J`a�A�҄�c9:�g�X��LR�s�1�eK�b��ں5m'4�4��>���1��=9�x=0�0u�,� ���^Ҫ�c�B�\OF�X�J�J�e��B��bY��9��y�1A�M}.��̍#k+��w�V<�0[�Yw��[A�y���KQ3Ak�U,�}{Hf��Y��;z콳T�ޏ���$yY���޾}�W\��n�e\ڕvﻡ����Zk!��G;LG���&�c���5�g'Y�ʺ���ʘ�2��ˏn	��w�sS�PFQ~�ʊ�]�$�,{�zfX�q3�hc��
M����.t!�Sr�썥�����ϟ�C����=.گ1L��e��hX�r�w�mR=DѶ�s����5^��@�x��nL�>�U^u�%3q�C5	�߮�l�k� }����;����/a�
cA*U6f�3�F�����j����L����츚��'&8xV�n�s
{�6
�p�x*��������z`X�<.��
� c�m1�Rɥs�+��p;}[ƃn�C��OsR�u��c���7�8�<LE�=Q#"NQ��׭O�{eь�(�E���'M!`�c]�䀣��j4vK����xzUcz��\{&��=�f|��E��ǓPAN������y��s�k��g��:�1Qfତ/�j��k��7�a�KE�&�WWy�;_A���<�s�Ϟ���R��Q�)Iѐ���JU �u��G��º��U����W6���y�N��r��B�xB�0�X� CH�����p��YD`�I�hY�Ǣ���F(v�:U��4��{f�F�;+��'��A�ȭ����0u�W�����Τ\��2���t��w���Ø�d�a�0V����#��ꯝ#�9識Z� �'�Qs*�zU�C���e3��-�ôf1P�JSw�=�2��7���f�_�9��b�w)~]\��,B�s�m4:{DeCj�y�� OK���r�yݫ:���J.��B�J���Q���ͨ�y\.���pS�J%�=��:�ԅ�׋�� ��n���N�z�w���h�k����г�������F��a�F�#P�ƥ-�e­�E�{@&l(��|]!�gD1s�rV����A�OS��J�[��Ŷj��T���.ai�&��'.r}��k�O2t2d!�΍�s.��<�TM�X�nh4ZR����ѥ��Qʩ�jx+�LSr�~�S�1)�Go�sn�g��v��Y�PW��a'V�y֦8>BX�G)ד˰����\!P�-���J��g��tCֵ�z��^��>,�9��f2P%��k]�`0��i%7�vT�!�eN��:��!I咩�˕��E����p��2�������S`F�imb��Չ�S�zH.7����%i��#��MoU���:�\���=�P�ي.���p���@�닱sӶōx�*U�t���U���dxY��]q��]6��f�&S.r=��c�9�GlKGNl߀���%w�i�H{3�F��+[��4���Yu/)�
xN�OHq�O�ݱ�y,i�Yjj���G����1�\&b2�L��r^��1éR��D��k�l?��qR�Dg.ʖ8�(t�O2�$�"�����ѣ�q�aS�<·��,�x���)����z�_v�r�vi���Z�kc��1wE�<������:�c&,,���i=º����H���oA۪�B����\oYs��.F$v,��%�Ͳ�`�Z�E��ҏd�+�;�7]�#�̼�in���7�������f�J��2�^`��<u��\jrʏ�J�X��eR���6�92�NǷj�ާ�h������kQ��]A��x0��8�]f�Xr_-"�9.&9�ػ��s����]V��:�5u��;�v茮��t�Z�L��:U����T�V[cU!�\v���3����m���}�u"�=�@�=�X3]�W��e�e���'�2�rˆ�MrY����h�d:i*���g7��FD��v��u��+�NZ�PϺ:
����c�Z�|��Hr�Zj�e�w��a ����R�ˬ<���g�n��Nsv���J�43�Ƿ������wfK�b�R�)�kE���H^�!�ά¶[9Y��:�"V�%3q1*T]R�����qn�,��k�p�|�l�P��`/�����Z����;�o�g�BZ���3��w���J�Ý2�,��!�r�Y�Fۖ�doei��y���}�rBu@&�3�=ofv7n�1��`��/N���g@�If��4�Ń��=[�ּ�\}�kh�xR�����|ewq�ad�W�\ �9��/jI�k�6C�ֆ��v.�Ayp�����<��ո��cEA��y�e� ̝W�A����%;N�u�A]Ͷ/���S�7W�M�]�dZ�T�P���yɭ�B��g:�G25X��4��Q�\�V37:��=�|*^�H(��a`�<}�3GI+���:»�;\�G5�9SvkZIZ��E�Ƒ��|��p>�oTuw�T�0�&����e�)w,�	(�vDy�s-6�L��Ià���:�cU3-7}|��u�4�d3WB�!z�LKt�5Kb�����m��h�Ӎ����D�t�
�<�_:/<����O���goϖoa���k�4z�^_�瓬�Ih����b��A���=Դ#����D�|iMx�Q�Wh)�&��mR2�P��ۢ�t�q�ҷ��h���NJ�v�t��ڂ���̜�J+�Gp���s,����ۋt��_]��w�d���i���6�i�ɳ�^s�p���.���}����樣��AB��k,Y�,DձA�b1�X��5F*��
�
��UUb�jь��5X�[EX�"+�����b�����F
�V1AEQT"1TVDT�m)�b���4�(�dDU�UEPF*�Z���TYEb���1bȪ��Db�
����*+�̱c,Ƣ���XZ�+R(,QUU*+R����ƐTAU���Ne
0PX*�
,��1��"�)U�����UA�Q�fe
�,Tu���AF
�A��(1"5���b*$F,�k*0QQEA1,`�U�J"(,��((��UUD][����{aDX�ª�n�lF,���dV*�*�SJ�k(�Xb���E�E�b+UQb�[[H��uh�D��2D`�ȵ�b0�`�b�T6��J(�Z��CD}@
�Y���v��i�1n�fɖ﵂p��p�9U�$�,T�o#+������ǫ]��nw2R��C@�=0Pʤ����9����{�_r�g��LvΉ�QQ�*Fnz�0T%���)a��@���\�+L �ڗ���S�����T��{
�Y^�XK��hW	^V�g&��X���M��o;��<�R�-Y��2�,W��X5ƪ���ъ����#�e�'1�}QhN�~S��i�lR�ޅ�&�w4��^�M����y3�4p���a�|PK�0�=�qb5�������S�V���3�̺0z�2�=������D�Ɩ�>1���t��X���35C�2NR�U�7�5��5�"%%�a �*츹Y\M�d��O&q�҉�qQO����r�}�O�T�-\�����
�9�r�[q�
�y�Z�Y���	)Z�U�P"X�\�ޭ�{���|'��BFCuNJ�}�}s��\;��
�Xv���6��bW�fZ�m�uh��K
�����9�.c��NcU�ܑQj`%�/q�^�!�ֳ� t�ӷTf��1������X��a������2lN�L(��"r��VxT�뫩K�^I�f&���fc9T�5:l��|�ʏR(m��:�΀��e�=���@�8�Cs�:�\�O�L:���<}�����K�;�q�
�t��*�6th�4��(�,����[��a(�����#W���쾏vUL1t�_}�������d.�~ՒV�Qxqt�g��xW��<+�惲���TC;˝�TI�ѵ��y����$�mQf�XW'n�����4��<����\�-S��s����#,
!:��b9���' � C��H���b�w��>���Us����=x�l�+c���_wc���8����W��\�(z�@�=H��"4I��W�g��h�1�R�*	��f�����:-%����⭭����4�O�;R)m�T�;�#79�Jp��B�-H¯f#'g�"��e3�����B�͙�kh�Î�4㮛q-ck�t �Z� ժc�i_��u������_oK2��W��F����YZ�B�����p�6��d؍fG��R
� �f9o���u~Ua����͜��>1싳ϸ�����%-��Qq�Mp>�9��L�P����Ὂ�m�WSo�pm�3��"���b��j��r��N����=�p�1�F��[�nOcw�6�e����������9��q7�� ���>eb�K��x[sR�VB�o�I�����z�G���Y���o����6�C��םM�x��Q�� ���\��qC�ۙ'WZ�k)�y�ڥgS���n$0i�v�㱪����_}�X��R|���;�zz!l������I��U�p��en-�}ϰ�Ȳ@�gl>lN�Na�[s�}B�9�&�и�鎄}���I1m]��s�e��.Ws���!!nӔG*J�;��qn�� P��w���f�&���#9�ǵV;����H8��y��m!�}R����b��u�F���8O���αW��5������iy�g�(��}�3'o�j�)9]��� �/���OtG���ɬ(=6LP�e
w�s6:�hq���Al��SX��3n�71�B�*I�X�O��c|3�^�FYg�>S���S-�d��]� &s�qP�Ԡ(���=�x:�ץ�I{P���Kp�[�Uf��[�H�{��W
�I���گ*�[7�3I�߯��6kѮA1^���~ݓ���F�>���u��+mg�ˁx�X߅SȻ����{nD�u��<�˨J�̽��3���S��yi$l�j*���T�L9����[œ��|�r�η۔3%�J��:'�[�P[\�����U�Y�f�_*��\�'�xoMsz��ZEw������2u.�T@Ix>�Kn��Қ�]c�]bq�kg;,%\i���Q�Yo�箺#Ղ_;�������sK���7��sr��FTM�>/��������!M��Ϟ��yn'�uZ�{Ys�LP��m-��F2���-6cn��������Sy��̺^�5\�<���E�]��0L4Q�K_n�M+>���x�7kJ�@����
�MnF<����r��N[�5�V2�;��{�e ������H����JI��䫥
���PW�S��[>x�ڕ��唤��LM0�s�Qur�:��JOۛ�ַ�0�n|�.c����C���g�mAo&1{W�wV���)����8���oq���E.�����L��M�[��D�����L;��׋�r��\|���E\a��V P�<J���QRމOʼl@��h�>on����F"�V�ֈ���
�ڳ��//v�I�s���D��'T�t���#���[��ѿ*T�i� ��&����������<�{w��n VQ�}Ϸ��A�/#�U]^uεV�N���.r|��&82t�S��!
�Ll���=�D�W#�a
�\�CmnB�6˹��6���L^����]զUmA��@R�4ѧhY4Sm�gbS��Yٶ��@�I���=���m��M��g�(�:�;�g���zQ�N�����o�Cʛ[D�W[q�����[�qZ����Q�t+�JQ�B42|�ܪ�nr����$�d�u:vͻ�W4ŷ:�6�S�V�NUG�S��!��8&rP���)ǹ��a�X���![�\�+�0��Iw3�5��Kx2�O��)�*�
*� Ӧ.8���Ogd�v���-$w���e�ދq��^/��c5[A4j*9KA���:�]v�y)p\w~g8$"/z��K�7���1�{:$TBYDEz9�H��DA�rփ�KpR�Y��r��pNkgS��`Y���B�Fxm9�c�Ue{a;�!\3�+v2�Ȅ��V�9�3����m�s8u�B��������v��Rkr7"���E�:������!��%���K�P�5X.&e�c,��*�Ei�Q���p�PRa���̈Iٳ���6��{�wu�F���V��D\����Ed�=�L`�Y��-���	Z#���3����Po��<+�7�"9��w��@#J�..VW~�rY]�e*��D���.ŝ��ۈ�*����r��|���u���u�Fs�!��a��w��=\$̼E����2��޾hg�mp��8-�h�Ү7�z���9�<G;��\s ��5i/y��ٰ�C������)��P�ٽ��X�+ev�ڑM��1�Q7�:�������;���&O脄获�F
��[ �,j2ۇf�e�c^p��Vu>�:M���Y�9�'T�?y�Ob���e��<�2�rTp��xs�����uӫ�K�F\��7΋��X��<yo_��s�N����5\n[���K���ݲ����#M_f��k�=*���1���Ep�U��ϖq�s�l�&��N�L-������,�R]6����+��h�zxW�F�E�3£\�a�1�Q7�AA�+me��@DW��h��H۪u���nE�Ҫ�έ���E��}�]N��7�4٧�:��tX��6�!�1��k�9>����xQ%w^/��V��Orp^S�M��"�B��<��W�^�+�CL^z�rDh��<���P�aku	�UuD���n�n͆�v�Ѐ�ڦȸ����q�on*��:a�"�����#�1�����R�zU��(mdq}11��"��d����W�د���;�@h�Qјj{�1����/�{�+xb����i����ړ/��+���N�]{f�l�r�#��%f�T��ɴ%N�H1��D�X{X������FM�{a�m�S;��v�"�k�tl��]��q39�N���ط6V늉��X1�N(�j�}�[�i�cw�B0,��]r+ӓ���q��N������ūЦi�������VT�oS}���]��*��GyJ�%b�W�BW	�DW_�eNu7�S~�6��;3j6�d�T�2��=Y"��t�����)+6`q��:�c��y�گ1�̀�%U��}�jWQQk%az��.����
r����f�
!�]QM�T�K����_V�yЅiRlc����oJ�C�J�[�c��A
4���9U	4I��Q�O:�8�F�gg�"�e���+��1�ٮV�!�ڻ����@���U��ګ��[����EB�{zH�P�aF:��iB��q���38x{T�G;�*���������J��W�P�T]ed�Y��xa<*d��y�X�BR��g�Q�mx���ݛ2m�o]�[B�{� ��5d�.S꛲|�
zj5u���tѪ{Z�*^f�u�P�+Cy1Aۘ���:ʎ��䚋,{�%�3�hc�������'�z�'����,����T&wX���jH�q�\B�����1#�sX�x��2�,�CM,]��5	�C�^S0(�V:y4���r7�fj*J/�p�[ՙ�=/��;�v&�7�fr�����u9-C7�Üf-��K�ռ:���'ӿU}PS����rP�yD�uGK5.�TPbᜣ|��n��jR�r���&�auS
�1�Vf�1Z�i�s��^�;&j6|�����]l.#z�}-�"H���!���[}��j|.��([�!��(pqY9gbg% ��LDu��j��艽�O����5��"��r.����?3�jȋ�~S^u�B�&(Z [ݦ"z�2md� �&E��3��Ѽ�����{���=����/�
�6�l�6�t�^ƝNT:��j�<�_�]��Udv'���f-)�����E��WI�[R5d3Z7�	��9��u3���9+&Z|��rr��W�%.�{%+,{�w���C�xW�Έie`��PG\b�:��;<��A�&D:ǽs�j[�n������T�VP��%=�Ϟ)A�6�u�9e)::5��FF�t��kv���[�[����q%�d߱O�E� �:V�!���Kޜ�N}�<�f���+c������Ls��ڻ�0�V�x����_�Pꋖ!�Gx� h�M9{OsԽ��a�rl�0����0vJ�x'v�.��=�g�'�6�r@Qf�"��I��pؔ���FT�71N��BoWr���)qN�!|���p<uT��w7���U��yHd}�мz��%���4/i%��\������Ka@��b�WR�J��{��f�ն�
�F���x=h�>V6J*���p�f��%d���uS\6�x��C>��:]ܡqn:�%+n$b������m��˩ᡅXz�B�/v�Y3�$ulcprF�����+1�]��pS��?���T��(Ohp�JQ<C�=�â=gwCӪf����z�.�N����oU���eyמ��i�������{� ���=��Zl�\۴�U���V����e��8s�׆P������UH�u���YD��R�\��ig����]]�!ￍ�߁�2^U_��4�3�h��8&k�H}�IAX�{���e�4Mp���'}\��Y�-��$s���S�˙�TA������o��f2P%��/j�ʹT��W�9�Q�`W�<��վ����"6��:x㪁4k��Z4��<��[}۵��w�Yk9�m��44��6����{:$R�dV�$&g�"��{j��^�]A��t��q)�X����$k�\t;�����%a��Nu:bk�j4��"4[���
�{��!2{&�R��нL֒�g�PR�,I�ك�φ��.k{=���k�<cG�ل�o;Ki��ƥ��+��ʰ�o��T�z��9��*���.\,�soU͎�Y�S�'jd�71���vG�y��^9�z�K�z��]C���*����S��il�R?D�vVE��b/pu��f��8'�qj|�Yq�cx�L�ģu۷�*��ؽ��v�C362&g��CQj6���-�a�҂ܺ��	�U�)᲎�����7�,GQ�3c��I��$��2���ҭ��Nu��q���d:�d6d:|��u����S��f;
�ȋNK1P� �]�W<N�^T.*'f���b弩H=�1|c8�Z%��}D`��[�%F��`�0��Ex��'_��Ml��d�ފr��
�p�j{]��T����ʧ�bECuNJ��FO
A��HJ�"j�c�}z�^���Xۨ�:�ͦ�W�H��T��ZL�"3���S�i#-���33*�R蚼�sK3K�:*���#��C�p��(el�.N�CaT�f6P;�Tt���i$w�$���cj�:��+�T^F��n�xVJ5�q����~�G���⌰j�{�7Oz���`g�d:�y�&U6�8�n�؊5��3ƞ�ݿ���{��K�p��ly޴FT�[��e3�\�֛ʂ �V^Lct�Tŕ�:���'��֙�SLU�Uj�5GG4tZf���,�U�qQ'�����joD��U�I!ӱ�bķP0�^�I������yw�]Zʰ;J�cL3h�����a���Js�SEv�f��K9Qt��	gDʺ�jŞ!a��ټ���es8��Z%6��9��r�<�#˂PNݛ��j�9]׷�'�m�E���^�7�uE���+�mT�z�Y}1��4|���^�j��N�nH_g؛I�)=�:O�X�W��4^�VBTG�V�]>{�oVAbL��l�==V�c���
v��'���9�VDݹ�贛�����U؝gN��^���Ú*Ҋ��
 �GdR�,e����=�2ǃ�-��.S�R�Iz�}t{"3^v�`ZX))���t�O�c��;̦��u�'{q+�#�%�q��St�ı�ĝ+�w7��(���#�.L.+�2Y�u�F>Yg1]ve�5ѱ����ʵ*o���ȔbRp�r�b�����Y(|�V�w[�Y�K��x�4�G��)�u��SW5˹a���	��{m�A�WMt��tKwD����m�n^ȇ%�S��]��]nU�}fl������	<����Eݢ0����s�s���]G1T˫�n�x|�f^\�ϺML��W��2�J�X��n��C-7z3�.՞�M�w5�{E���5�kص�]�������,��do_ۥov�q���1)!�q�4Y9��,:�.n�.���Õps�����u�D}�l�f+�u�DlT�|��dqķ�w�0��bk�_٤(k��5�'�Մ�{�w,��ޫ�R�XD�BC���Jp̼Pe�
ehR1��fa�B�ݮX6�_W5������7�*VNϸNQ ��㣢��7���Jj��1q��ZC:u܄�vۚ+];�ã��m�'F�ά����^�fh3������IS���&����s�ys�&��E��i�@�g��D�	(�!}n���fecʺ�
�6&�iw;�����8��$�G)����[�HoH"��,�+���4;Pא���,l4���*�xlgV/�F�	yk�E�����=;,uq��K�i��G�淆�y�A�2��9-eb)��4�����E��o�I�C��S�pC�7\��J�v>�u�Y7w\ShGt��EY͝fS�j������6K䝔��̣ў A.Wu�9T385Mww����<�Q�p��heom֚hV�uE�� ��+yӥ&���WRM�5�g_���B�#*d^�T��N�n2_@/��Q�|a<�*��k �h{�lY�u�c��:xfD���k0�1;��lܨ/��>�q�l�}���/���)=��E�e��4��Ҥ�[���hb�rql꘧7l�E�j��
�$=" ��=  QeY�����Uc,@D�
�X|�bj"E"8�����qi]Z��Fm�-�+F,dD̦(��+1�F,q*��h��Z�ZQ0�%�ADejDT�ը��"�������,,D4�b,b.�SMb��"F�TL���f5���ܥQY���Z ��DE����Rc�V�m�,b+DQ������""�MR��5���J���UT
ъEU`�����`��0Q2�X�*V�RҪ�Eb �X"��R�V*��Q-q��":�DT��EV0[J���PDc������U���V#wqMڲ(,��(�",���V*���ݪ�*�TQQ������0�QET`�F1f�EQE�EX�,��Z
0b(��Cv���(+b�'߳��~׿g�k�g��.�Z����g)%����n�3V�h����(���Ӓ]κ�����^e�x=�Q�خ_��rp�we�p���ǿ>�N�E�`# F>F���4O��8_������\�G*��UJ�gRօ)����
�ر �U�����%zɳP:��"4>H�W�O]A�Ӽmq�F���vNȂ��9�e
Zb�Kcj�#������%���5�p� E鷸jO)�`���U=;Y�/�����sAҊ��|-���!���UV�s$*-���hv{:}P.��S�y(8��#�����|�!^�!��ŕ��j�g�c˓���D�t����J��"��j������������<0vq��`�^&
��Ɋ!R���Kn��>f��u������iGC���Ά.����������08�#>H�:��@�E��)�s�#;[����=UT�=�ՑN��r�
r���M���x�<�Uuī��e\sҗ����ݬM z�+�mθjz���0��~��V�����;PB�$$m¼�8*v6L���Z����pe$i��nXXa�¯��h��*ImUB��n�a�-k%�$���K�Bwj;�Y�<���l4�vi�Μ���XZ����Gb���y�Jf=�ptK��i^��n��s�\��U���j�H�o(���:f��>��ׯ5��پQ^f^n�{Pr6V&�I������F�
]!b������kΪޙC�RC�P�,�96CJ�1�����5Y��/��oxa��i$�B�\Q�t%_�߳o�LS�s�d-�B�WYY&^S�	�S%U��U`�[�l�+�О�6��5)`T\GVV�9�n�nመ�N	g�Ւ��@�MM�>u=z�]em��;Ε��3uy��-ؼ/�6X�����YQ��I;X�K2&r��6`�tfb櫺�j*�Y;��Ŧ6Z>��Q�����|Y�{ʢ�\�zQ%�ɋX�p��s�J.�Su/�%|�� T՝���~�s�f�g�f|��[#�1Pf��]���ؼĩ�2l�0�U�K���W�R�e�L�b�vb���o�3[H�b#��Oj�-�u+�d��싺#���=x��\ә#���Ӄp�qy1B��K�ԩ�ɺ�J�.������s���T�S��b�5Rk�l�=��sTf�d4�Fٮ���:����}��`E�}�c9-������i�3�V�Ɍ�+��ɑ����`��9��')��N?`�j�q����p-���3-]��^��I����N;�c�K�t����.���9fOY�kЊ}��8�D͎+܄"R��7X�E�9�Y�n�3.;ą�1w����V�T-��Pc�t��so:����s@	����7�}轋�<�g����0F�U^�r��<��L����ތ��PG^*#��%o��aW��K�zwi>�����<������f�*x0�
�y-,�a�7s����`�8�|�T����b�N�r9���6�u�=�~�>Va�+J�0�aZΞ���10,�U�2���=E���W{�2��t���Ψ�OV\�;y���Je�cyN����Ry\0�zk�~s�˱|�Rn����F��%cd�+�bɱ�n����u�TA�Q���fdH�{�r<�&��pS�u h�[Yr.�r=cG�X�G����&z%���4�].rQ������{>{���*u������:�;F��tr�5��2�&���t�>p��)u�=��_s��j��/�\�:�]1�b�:�73�u� 7rI�<N����Mj��K��E����=:M#��
Ñ�tk�A�3�ȍ�*v�/k7~;	;E�`6q;~s�L���v^�a��S�7=w=��f���}npLײ����� ���s�4W���8��;���v	��^v���B�!
���ܳ��]��}��C��\@��w�qǲ�$F�x��ݸl�U�f��B���Kjr"�(H:ҙ;c�,���;b�/�^�>���Z��}��rgmvۺ��ט��N�=T��-���z���uh��Dwe����j��t?����l=��i����Lh�1���TԻ���y�-������nlD��<��q�$�˅4B�솫Bh�*9KD��y���q��!@m���X/&X� ��Mq�Q�B3糢EBYDG;��I/�u�Z���h�4,TL��kU�݈tu�(+\��J�0��p��7�LKٍ'�̈���K}���u	�e.���l�'�ȃX���%��J�Z;<��}Ď;֤S�^MnF�.��p�\�ME�o-ƫ�;���Z�y�ֈ�5X.f{
5�6��(B�d��(,�Soy_`:S�-�e���q=ّ�Q���t�S6�)�����E\eTs�Q�F���A�s��Y4�{"�<17Lj���(#j�F�%��a �*�.VWq�XzM^�=<�Ъ�=�!���u
���X��}D`��[ �RU�l�U�1!�HB(%�dU�q�dd_a�S�j�p���r4��6�mK���̽��bCs.J���M_+�P��ݭH~��N]�^� �Zgn��
��P5F���nm�b�L�t6w�G:�u�mKc՜�@���� 촻Z�R��s:����g-V�%���ܫK�ҝ�o���w<����y�5�t���L�v7}�DD��f��3�X��`�f,+�	c��m �z�E�^T�8���fH�Ԯ&�[w��qZq��D��<̓��?��Dtj
!\/x�Z�l)0مb+%��pվ�͵�s �[��p|L��Z�I^���5�*U�����2��j�^2�_K1a����UQQv(���'�ULq�U�痗\͓Lt+���,Uͫ@ܶեy�F"F��̖z����t|%T*��F�^O�D��NE���eb�&:�m:g"ss9:�ܹp�$�a��ؿ!qTw���<�'X���4VژjxU���-_w�<������FW�^�>��Ɔ�R�~�S6=q�5޼�,֟s!��{� �M�o,�>��
z���W_��Z���t�d�H�W-���q������X�?t����Vezy�b�xU����t�S#J�e��^F���$��XNGB
R�S�^�򮽑z�^���:4m�T�*;�}�Vx�DZ���p�J���cJOw�S�k�>�Ȿ��FT٢{m�S]f{�Lg*�^���n��;k�c�ak'^gX՘YS���W����x�5�&p̙��c���Ev_�F��ϮOы�I�+*�w��l�`9����s��]�E(��Y��J�K��_5�V����iy�zc{&,~�t���������R���08��&,@�L������Mm$���:���=�]���eĩ�
6�9JN�'D+7 �Z��͜It����]%ܹ\�ȁ���a���C�#�_�#Jޛ��C����-�v�_eЦ�o}�</�����&�43�^.}�*԰��',�/�����_"r�{&s�=q;��v>�����qL�8��FO
�p�I�V�pT�c�1�P���H�4Ndhڤ��*��v�c�z����||�-"�y{����1a�\��0~��#:��Tm�q��3uaT��Q���j*c���2�R��gI����Y�a�Fa��<x\�yH��[B��W!Qp��ة�J�Hw��[+����1%�R�OY%�P5K��A�������z����5��T״��3
�����bC\�q�$�楓"]�J�w�3n��ܶ�{0h&*�N�E��w�O�U��Tt�-�q�2��y��I�S��k
A���(��Q�cٸ7w
��*G��xc�ٞ���w�#1�JyAf^C�)�H��;C�[*��]ל���Nq�l�g/Ew��O(f^:u�+MÂ�91�5��ݨ���q���a��>7��;��v�7]N뻙��)��=m��q`2~�p���K��b�8Gj���'��_c~O틼O{�.��m�7�V�kGr�O�.�[U�J��y"6�W��c,�vi����~�b&WMb��I�c���l�-��ׯدޘ�ە��`��㘨
�7�손t���^Ĳ���0�r�����:� �r�e�*d�6�e�U�kj4J���e�43��ӡ3�/f߶Z��T{��o+�:�E<��9���U��+�<�ӑntECKoC�#{�m<�bm��&Gg؎v�{�r����)/;��3ѕ<�BB����m���8cTω��w�G-�\����&�l`��0�k�Z�؈�&���֎ãpԶD���2܊m�h�ĳ�/4:?PG�gL;Fa���*�ܪ�*:z������f3
ދ�!�6)����h
�2�S+z�� hθ}dkn�{ag��b<zU�`w�;&��6;O�o�܊Qװ�HtviNj��!���q]1����<� �1meȶ�܏X�¨��B��/���Y�� 3&rꊏ�Ob��
���K�G2_C����� ���vzT�M�4k���1r��C���ŏ����q<�v��M�S���0�OTwFs?�(�u��*HA����=p����a�=�`��1��r�.��v����$9A�ܾ�t�����t��ĭ������Z�Q�Tvוzr��T�i� ��$LR�O�;��1@2|�$��
IwsJ]�{f����pW��'װ�t�Q��T��:ڀ)��H�4^�D�oq�P�a(�U<�&�Vp`��	e�������[���*��~����������\4��Ow�wneb��@�7��?#s=w>������4M��3^�C��Ppv '���I�9	]��,G��Z���9$�hIY.O����^J++�4A��	|�OJ��՜=�g������ z��z&����;'�͈�\��$u�!e���QM빓��C�k��Ȋ}Ś�յ��@>�a�Ge�=�+�e�r�U�ժ��sm���\�F�|�)\�ʬE��*��t�9�a��ӝF����i9��S:�δ��+G�����KC�Q,>b�.�T2�Z$P��Mڟ#̫���9�ӝv�����8���VgQ肶�C343�3�P�:��ڤ"��U������[B�H�#��kA������5�%�xS���R�WyQR�;�mNNp;�;���BS�m޾°}���]�յm�eS�bgɿK���`����Wȝ��]��x�V��YȞ�����`>�����^��d��Mw}�<����Z׎��߮��W]�d7��vx�EA-�s3a�~�ȫʨ�LVp���-����(5��T-�vBv�\�v-N+���b��4��������ؗ�N=��9E��7���\�7�-�u��06��l�*��E\31)��g0��������Q}�_���R�}��%jf���銈�'O2��lH�꜔n��`}n�	ĎN٩���/W�E �ň[�:��PṛH;ޯl��1j�Gi���C6�y��ȗ��J��d<s@�M�\�`p0�"�.W6��8^�\-�,��9ŅR�]�]�󛗼ުP׵+��1��ʦ�h~Y%z�/#]**o��fQ��P{�·�/��c�gh����TCآr �w����R���U���~*��?rj���W\ќS�!��L�]�*��d]0c�$uߜ�	�*6����b�꼌�K�y�Է��G1M�B	3Pu�ۻb��5�)�T='Xu��F���RM�"��׻"�2�j㸔���R������j��.����(@�N�8#ˬ��x;����R�zel��إ�=Xw^>=��8m���
'�����e�Y�u�np�b���&���ݔ�H����c4쓙�G�]���e<O�����;��Z�Iu���VV���xa銍(�l���e||��ڊ��{;Zj��1�o���w�5�
zx������Y�cl�b���LFLl�HT['RuS#Qr�ӝ����������v��U�h٬�:�f��tҿ�V���ו\3-m�2��˭"��.�H��p<�Z���xG_�����Y6#vb�_+�80Gg{���L���r�eZ����__E�]F6��Q���PbYA��+o�IY08���S:.J��A.W6�ཌ�q��B���<Ϻ�ɎQ����(F��lh�S�S���rG27�1h�K�X��Y���voi���͢l��]Jϫ�l�o�i�K{lX���6:�[]��_^��RG"ʘ]x�5O�EZ�g�銝��g�e�t����¤���,�DI���"^��<�Fq̡���+ѓ£�zl�@�i�<�xJ�ᮍ^��X����#r2�5+{(��ԙ�<=��߀O�E�X���.��v����¦
��b"��I��C��N�
���k5q8*��$��s��X�;Mj/.��CF$v�����Ԭ�܎��㼛m85p����o]�|�Ѧ�bw5f���ˁz����*��n����ۙ
HXD���어kpݻ����-�o��K�o��A6�Z�f�(�]��/*vT�1�`�V1pZ ���N�N��Ef�=%�:$ʕ5-�뢂�j�|����f[\�{[ 4�Q#��6��Y�Y}%�tz�D�˰��Ϊ
�N����֫ e %����"��GK]
su��]Ņ j�v�h��Ddx�7Ǹ��an�ζ.��,@kX�+��v9��(d�3�U�W
�d���q�9Kڎh��B�g�+jP����y`L�78f������e؛ײ����+R
E�ioj�Y�ւw��:�.���:�e�{���-��4G��Թ�ou'VS�W�&�r�S����Wsgt�����	gxJ)��<�xse��ռ�f��J�:�r��^���~��n���U�5�vn7����=*�I��{w)�SA�����[gA��^0�vj�6�Us9��4M��Ғ�m���L밡g��T����B��뜎
Q�����V������ ���ڝ.�,��lμy��H��}]�u�':�a��*�,^�'U��fU�|/~��t�H�2�5�7x�7+�����oڂvo�P�2��V���G~k��hiX��PC9X-*���&&��9�ܷ���R�/]�a�]3xG��w�Kxb�Uc���^��7w�h��0�: �ơ쇟 u�<s:Y;��S	ʅ)�.r��>�;�Z8������P&Բ����񽝇�f�i�Ji�I�;7�$���p�#��'�ZC����,����a)�Vb�S[<o�݌Ej��v5��jh�_3���0�.t�h���V��d�Ajp�S��� k7���mr���g�t�%]�	m����� �v���PsS3�����&k��G�ez<[&�T7]�S��]�2��8���,yo!C%�i|lh���L���G��q�b�����*�9��'0���<SO��B��<d[ڔ�P+�7GP���	O#�S��%ŧ+��t!f��j�ә�nY]���b&�T��hjc�8��v�����&��(�E�l�g�w;���E���q�!�B�)�V�	#�1���el�[G 
�	�'�����X��ۦ��9�r���4Z�n�kx"�[�7�zµ\�)k ��B�̔�3%Z�ѽ��ZQ� ��7-�Z�8\�1-����iV�G�^֔���S�����Ď�z�L���}w�i�O���u��`G��c1c����6ԣ�:�E��q���j�B�y\N�[q���+���s.�����KP�>��-�gK�黱s1v9�IbK=�4x�� �� b��V,TEG~�:B��,AC�QQAA~l�EQV,X�F*�&�r�+EҢ*��Qcb*��F+A��EP������X�TQUPD�k*��"8�TWM`��xb(�X����(�,��4F1X���2 ��+��H�Q5m��X��*+�f#�R0E��4QA��w�F!l�XiPR�"m�+q��Q��"1b��իEy�DF(��X�1��Lb��b��h�TEX,�Q�Duh�E��b�*�&��".�X����A`����ݔX�(�o2آZV*�Y4��Z1H�f�Z��)7h(�;�EVT ��"E���Xi1R#m]�X1UV()��&��L������Q�^ZӨ�Ƒ�N��{�����$���ɘ2���'6.�`f�i�}��類ܦ�T�<û۵�"�)�2\�M����H-���hb�F�N����f�ሚN�sT�[=D1q{��N��U�uHc����8j\#ô�1�vcc�b��1!3�nw�"`��F$�4=�E?-�t*խ��Wu`T�d������.j4�¾�j]�r���&��I���;�Y9���mn��P�i1��a��چ.�^�:8�ɝ��ٟ+�L���T���=�9��lgͻ�y\�a���Ӏ��ځ;fy�
��V:���W�R���6������+�TN�io�]��T.˱V�l��
��2GeÚ�g����U9~��ޓʼfr��&Z�p�y��d|�����k�l��:Sɜ��b/��Ă2L$�s���X�r'"r^sG`��� ��Tc/]"j<����C����o��M�ڑ�!�Ѽe>̬�)�y�'/Il�>g���詜<����r��<�Ӟ�:"�����*#=�@L�6��9���b"i���py��\L����	��ʞ�P��%=�Ϟ)�΅
B���ީ��Z�zpsՊ��=�`,��*eߴG�IR�(d����z�p����[SEU�u����ʁ�xt#Z��W>�����Yù����%���ܼm�=2�b� �����]�ɭ����c�o��g��r��s��|�{���eق⡷˸�h�s�d���	i��0�0:W=�'��*�}�*��Z�J�v�B���V�7�eh�[/���PSɇh�"cmusp�TJz��#��!<)��s���1pL���%��E�A�<�f�F7�Fl6����=�a��Q��ϛ�f����""T�oE��y�|��h�8�Q�&+6��s99�y��ں��n����haTF�$�f1���7B��o^��TF��ܛ'���ju��ry��T�i�Ҩ��
���t��5��K�)��撱��Dp���VI시�Xy�G�6C�t�Q��-��:ڀ'�(�[�5�PS�sm�{��,1Ĳj��P�t1>�զه�QZZ�F��g��g�d��9cǒF��%�>�������Sra����I�{]Fi�d�m�	��C�r�k[D��:���7�B��C�"P�5 *O.��#;$�hIY6�}�),5���}��ߋ�h�ZyY{0��� �h捫 �8 ��L_�:��76"Esʜ7�$�˅4B�z�.���`vfߟqq�J�P��nmڽ�GZ�8G-�,�ƞ���|�eZ� |F*���iR����_H4ou�H�:�m:Tމ`K2��
b}���P��]x2[�k�]7�q����.�WM�7н��R�Ճ�ɻ���.>X(�Cϧd�]/��h�q�W��F���q�Q�� 3>{:$%rDs��y�Ñx�z'��6�\V�&�\��ڱE銈����]�Nya�':���1*U�`�QOoqbWۑ��k*Ep���T�d<���[VkG<�v��s��X��=�?i[]Ow1u�zy +������7��-�G
��j�\L�aC,�/fP�GI�>�ڀٓ�V~9�|��3��x}��A��q�.���V�뒃��v+)%������wt.go�ȩ�	��v�V�P���D����q3��8�D&K1�f_=�����nW������ܰ��.!�ٓ�E��V�7�B�,G\>�0T6�؁EI]d��=����%�H���ֳuDPl�$5��c�J��͸W/LT%#O3���=�t����I�p�v��Yՙ�Sɚ��H_��`�~1c����s"6�w�^�I�s��q5�"U��Q r�Ѱ�3����﫢Yn��i1y{�A�r\�:SPxS�/AB�gYu3L���G^8k��9u�]Ҭ�����;ԕ]���q5���Np�v���92�NTS�r� I����������c;��f�V�jcSɋN���.�l���g����+Ft�Te.��v%�35�Ϟ�y�ɏ5(P�+����|g��C��b6mLo�9����Ŧ)uSyd���5�QP���^��i��#�[��{&u��tmH��oK��	E۪�`:CNN�ު�U�/.Z�ϛ��U7=�R츟�����qy(`~!	�˸�P��d],��"a�:��;6���c0M��x��]h3O7=�s�ab	3��T�xA3^�p���b�F3�t�q���z�.\{�AB�m�t՗�;����Ƌ5'��w
}�\hK6�Ya5�y{x�Cl�&���5ժ-z�����Z+�$1�Ϣ��e�}>�Uj��x��m�b�O�vy�zp��*Ї_O��l�5�pƳ�וuȨ������3��)<�mmaF9�����h�:���,;�W�78����1֦)�3�5�A��B�h���ِ�wR$H��U״��똱��.������)+6`q�F|��v�5ծ�%��imr�(Ր�Z.���W�mB�/3�3�S�4\�����Rv��;�:�R�Z��;�5���ٶ',Q�Ǟ�(���%.K.�i6�-xmQ��)��6�gF�L�]-�ҩ�CC��η�71��|x�ظ��!���ϟ�lchA���f)s;B��M!
�7wݗ�b߅�Xt�y.�Za耚����b����2�6ɸ1�#rP�������7d��/��s�I�My�'SqOf����L{B�i!#�UB�A�8M>��
�!�*Z~�����۟ �sY��s2�b�Vb"��u���p���t*��ل�%a�O/�X��Ų̜���Ҡ�����а��W:��N�3���V;�Ϣ�+��z��V�5�/Y��..�:ʛrtt�,��gN�ncB0u�,t�����1�&��3�Cqw�U�5��B�j��yѳ�^��i�X]����:ʎ�OnI�,{��6����_rSִ �3�hg��t��8vkO��Єf��.,̾Sp�Q��Z��/����Jnow8�$�<M@�KxJ*ܳ����x��=�{a��;��1v���,�޷w؜s���ܻ���ٯk�Oa�u,Eʤ�x:+A�ݫ�_/�> �3�ו���;{�\-<"��M�j�Cې9]�M?	��#g���le�� ���4`��IȊ%�́9��h���5{�6���=
�L�;i��AZ��c{�)=7i��/��vb��-QG�
|��۰:�U!��s�)8Ә���y���gT�;ܽ/SM�\GaȆt�Fݮ�����Xh��ἣ:�nh��u*d����p7�������ƳU�U5�\�R��9��$��V�F,Ftˈ�0����J�m��j�!mmF���]'L�U3iU*ƩX���ggg�m��}A3�7��qS8Sɂ9�U^�k����^��:#k�̻fD������������$T-.�6��9�V��X=qG�f򧃸(HU)�ߛ�=Sh�B���́{}�sg����������LP�*�V��EĞ�ɼS�f{+J�ܽ�Q�J�PW���i�������^)��@�&1l�R���*�a1eeq89��t���n�
٩�N>hn��pF�jw��"�o��mՏp�}ф��z�V�^��X˸����M)�"��_��D��i�9���R���m��ӹ����n�4����#ZGP����fwa���!��<�=բa����r��T�~Oh~/	02�ν�ڋ�v��C=\T���_�H;�����K˜��(<�#հ����1]J��w��Vm��"�82&�ṷ�����6�s�Ub�⭹��.&�V��B�+d8y-#BD�o.�k��.�Q��{#�q��ϗi�nL�8��fH�r�q
@�m.ue�V`۵�P�;+Z�K��U��ɹ7;��X�� ���J
�G�.�q'
qv�VK%�u C.Z��k��Qj�q�6�]�ߕ�R�]*��A�!R�C��'��]WS��(��fW�q���^�����,X���a!��2��uݶ��-��:*#dK�� :O.��FvIВ�oΧݗ:a
����ʻ���HBcqOv���r�ϲP%�B,ֻ'�͈�\�Ƹ�;.!M�$�Uc�]�wk�KbAO.;.c(Ք��b��5m�n%�:$g��"�ӏ+�+l6������2�ޮ,�+���pTg�Ӌ(.���ڂ�&aa�L�&�m����n��v��ۓ��4�k*Dhf��g9,Y\K�K5��g�1{�38�x�K�b��y�x�d���G���ˌ�1�}^����nj�z�1�j��}������1S-bZU�X��c��;*c�r�2"��n81%C��VS3a�� ��辸�D�X���g��T5p�4!Q�X��z%��펹��(#j�F�rY�f�z0q���ǃ�KXR�Uu�yd.F�SEu#�b��uj�J��ZaX��YU�[��L��v$�{n����m��i�r:�E� si$Wq\�3����+����r�-�g�V�Lud˧���ȳˮn�io9p�/�,��PtQ����R�p��J�Luj�\��b�eq7�0�ˌ�\j"��$cx���b:����x}j���ޠ�5k"��vbs�����f�e��p%��g[�Y�x�mB�I��x*�K�r/9S�ݐ�"�����]Y��C�T���|��d��(�\4e�>u3g��*�A;=y����n��b�q�$k�ْ)�8�-��ي��C���X��}U�v}�?5�kqԴ���A©��2l��d�V��LɎ�n�ӒamEB����-����{�b�V��Q�Q�z��4%~�U�x�E4�@n﯎MV8�:W�mH2�r�+R�Rl���q�Ə���K/��jd].
�GVǡU�o\4�@NG."�ߪ�4j�~5���D� �9[|
#GZ�q[��P�:s��ON6��Z���1!��!�I+!��b�y����5���X߼D�~<NJ���	���@�[]�E�Ԇ_�~�q�u~�p��
�_�Z)�Ɓ��܋��4�-��T��.}�[�n�/T�Rc�p�Oa���WOp1�j�U�k�[r�"t��^�-�y4��1YAq�0>�/m����5U��t�g>����m�#�l[�-n<�@P��౐�����p��$u��kH���]���#�೤)a�X���.�âX^Gb���+�D�8ΟW��l�[X���rƆ�T�ҿ�ZХ��G^tt�`k������ߔ��\Xw�����:+f�[9Q�S��V+%W�@TnE��!�N��ʷ��̄�UG;�Tcu�X�.��r�+��c}JJ�فƺ����/�7�UR^v�:J|�����F\�*�j��rڅq��r�j�vƂ��8^�l���In�*̼�/uŐr4ZCld3A�<�b�*.��s��z4��ZHxc�!DlY��7Sۭz�p�}��S�+��!#nUGhv}.��g���+�hhr�R�ef��/��W�S!�ߟI1m]®��U�����}ӓa>��K1���q�a��}�\Ӟ֐�c_�nY8��t��<=���	�J��Z7����nѮ�|����	�3�{�}׷u�"���
�:cCშ��c�����1�N�sT� �y�0�v����B�~�b��ǘ?�B�B_0h
�6cc�b��1!3n������=�����]�u]��H�����T��	��<��7q��`qy�z�eJ:��O"�$�oSX�ЬN����'@�c���\3Orܳ��]�dy�Y��=Du�����Ӗ��|�$jtm^XPv�:�'�]����~�7��q�]�ȵ}��B�A���\5�WIYU�O�|�p�����ڼZ���Lxcʛ}�:l�O܌|y���V���@�ˉ��|4?��\%nY쨰V�d�{g�cj���0�Ρ.�Y]���ZGuL�t�I΃(�t?&���u�ڸo��K�]7M5�o��Sɭ�i��v麭�s��w�������8�^�$���5�G�Be�S��*%��N��Pp�@ν�"z�2md��_b������0{�q�_TfN��)�Prq�w��w���g�)|�3]f��0ݗF3T�P�b�U�kj4[쮓%ϳ���*1ݵm���Ѭ����ί+�L�o"`�GTϳ\�6�"��[�k��V���t��V�,���{=���W̍�r��o�L��c�T���Oe	
����؅��Ռ���m[�{J���/�cj%u�.#�ړ�#X��^R�j��_��M�)�E� ���՗�t=���̎��7F���y��L�:
y0���"co˨��T���-�m}B��M}�ͫ̔$�_��]]۷#�ov�Aq=̎1��%�Ӽw�m�XojU�)@�,��8�xq=s���aY٤������0m�)�,�u�}��
�=�J�g�uh��������� 
��0������:�m{��X5�)x�g�SL�3�!�����S#����t�O)�b�\��겸�����B�b�h�҅,����^mN��4��S҆lvi\�ϗ�HTn��t���q���F�q�|�K^�p�����k3{�
�I�[y�m`��u�����y(Z�^��gP�B�&�]�.$�;qM���vme���4N�F�d�����&^��2�7�:R9Z̎�þGkA˺��Q�o��[�HaJ�fL5�9�ť�s�i+�.�z�+Gi��Ζheh����CΟ
�T�j���af*O�,l�)��d�Y��ّ�=��}�l6��7!�����lw�C`��%���_L�w��=��w^;5�e<�����6�;R��EPO�֊ӣXJ��W+2����:�����[{HfD�����r��ʍ��R�Vf���X�OB_>|r�m֎��4��/
u��BC�Zr�A�ts�̙ʹ�c6���
�����y ���L}.;ǚ{��"k;GmhνQ�D����Η�����E����)8Z����o)	�ׇZ��j*�J�����f���C�����ܫyW��4�{f+��Y���wD�@����8r��d��s���.�����j�kP�L�\�������&�^_l��l���wV�Ζi��g%�8F�����4��|�e�Qۂb���g����j{�qG�̂6�P���a�q�W\㒦�C9�NB��Zf��iE�/�I���b��\��<SE�?������r"A�*&���X���(K��H�×�#��ƣ�ˢi�kߟ�z���^�s�zN���fp��A�j-��vַ{Mn������x�����} ��+���2�Ozq橩-5@Ǣ�`��z�^��=�@t��6�T��i����qY:��j[V�.� ]�A�V;*�O�#4*V��Ԏ�9��XD��U9Z0rܥV_l�f\�׋{�cLC�7i� ��İ�Tt��=rz�O��ι�����
�w"l������u��e��+�;�^TCCu��x�YO9�p�q^
�VY뵐�:��d���nm��L��x�@�#\���=������M��$5�T�zt��X~M�]�;�����J�JunG+{'u���}���f�W+�#�¶���ﲹ�ͣj5���p�1FV���-��n����ͧJ0��[�L2K��H�+�X����|�'��R�˟kh:�z����[{������I|��u�EƍK�Hpլ��%�$���z��f�wi�!�ʼ휎�x�)�Np�;�������Z[��Em����QR
h�l�*��U�*VO��E�+��X,X��N5��dR*�X �Y
��qA`�

EH�f�!�PSV�,���&2Vڠ�Y�e�
9d��X;��VA �Hc�i���E��DTD�F"��
V�Y(1�m��**�HbT��@�+��X
AQ՚pAdDq��+DA\����J��P*1��Ҥ��(�,�Ub�Y����
$L�c"
(1EAA4�a��F��,]2�:��T��ACB���s�#��3�5��H�젚Σ�cF�����;��i��*2A�x+{�E̲o J�-(�L{I����)���i>����Wl���K�Wc��:���=�@ю����m�!L�t@�(��=@ �R�	�1]X��(�YdÂlm�'QY��D�m!t�4rs�J�P���Oy�!�2��N<]#J{���A���_Y�ȸ�1r�гCk�����W3~T�i� �UҔ����Y�%=�H�x�Ytǰh�*nnJ�\�ݿ	A��X>9�:�׷�SEc�L+իPԀb��N�n��U�.'& �ktI��&4C��J�I���G���_#E��n���J3�6�(Q�!�6O�CUH��[`;���1^n@�7T��=U~;I��F���1hԄ�S�U�Nw�b&�T��"J!H�=\�P�]����)�%d�:�v\L���`ۚ9;�㐫�Է�77ń4A�� ��L_�5������H�yS��đ�N66�V悼�g��}usB�{��U�F�Q�Zl �g`1J��l�r�e��swerB\�U|�c��!m̋���.uȨ�ڱ^�������L�<:��&L:�ͩyT��8bn.P���r�`(tn��*P�]!�CE__A�ŭzz�{�J�I��}l��>���̻q��o�HN[&r2!�E�;wt���}���6�</�g[7�;����ep���}�P+,ʱZ�r=�Z�<gDM5 �q�-]�9���0v�����'��%���+�c96�RŐ����S�Z9�x'��Ͷ)�l�2/�۴H~cɻ����k1�|�z{�<�I-����>���Y�Qs��-xܳ3P�=+�lC�gDuFO��AeLpn=+�"�j7��k�f�w�t���e��-?N2r��Q�*�*����V�b���D'lu��v/�q\��NK1�m�K�[&b][��Z���;t�ܤNA]�-4�c���4�K����ۺa��	���]�n���^�����%��W��;�]�}�a�6)WKqxj�U`��m��pА��9+ $kѓtb�=�:���s=�����e�a�+Yp�S)N��qյ���Ft�ݠ�r`�&//q���eIr���ǆ��vuN6����Zg��=�{n�7=��N�b�L6b����Im0���h�,����7q����Tq9��,܁%����\�Ȣ�k���Д[��`:G4��7�aI����u�!�����-��ױ�Z{��#����Ҟ�v�ɘ��t�jn�_6n���_S�)*��ˠ�7��;/P�+�43(�b&K/d=��t=�෗1�˜�k+�2�×43I�5�Y�sH7k,ru_su����z��x��k2�X
�y���C4�r}"���ɪ�s��ŕ�]��<B�,�S	�*K ��#9S�AepLf��ժ;�![�)��L���7=�G1��
I���ۻb��5��3��L�q|M����W5�kg"���#C�2G�:�b�9|q�l�!^b���{���rP��/�;�S<߳�v��>���5��
�E"�n�èfyz�*_��Z*9��>�Y䲽
�Z�p��ꩆ{�C��o�ևg���g6f�8ca�v�ǘ+/��ı�RVe{kӭ��(�����>],<ȵzs�荽3��^s8#E#t������|�� �n�`�[u�1�5��Pgj���/һoFD7Ԥ���5c��c6Y���l^����v�&,`<mqsȫ��y�[0�U=7�P�YN��hQew;˷9�9$k{�#g)���7D+7�QוuDi���	��C��_�4��sE���s�E��N�Z�|�'l�FgK�r��
v��~$$YS���B>�W9xuڮ2�!���<ɬfs�ws^�$s�M���MdW$�Z�&��q�v����B)ԕż��7"e�J�z�0�mR�l[��L�sg&�����j��4� �+�n�R囍�C��ť�O��[�h��<�%�=J��7�k栰�;���+��x�3y�+���)��󘸁�7��>�"ڪ���g�zHB�xT+�}zH
�0�_�sʲke��Ko�o^�Ǝ�1�X���f�:L���]�w�'ԩ\��o�(W�^�sG��˥�}�3Wd��y]��O��a�Lhb�Q��T�Ny;���>���(��c�C��H��}�i�8���/t߮(�ɨ���d³�����	��:ʎ�}yٝ�9���uA��sCzԓcG�s2�����V#��k��|�a�J���nxnz]��/�2]n��a�s��%ʐcզ٬�:�%��������,u�ʼ+ntk왭�44Am���K�^Cyx�ѳ���B���IH��T�O.}�Q5��%��PZ�c�4�U��(��R�dx��&֠���-ր��[x��������*�~�������sS�˭wѹФrֹN�l�w�+��v��J�*ϐ��8������˱�{��ѡ'V4�{VuW,8�|��[v4�r�9��5sU"if1���C[Q�i_\Oh�U7��Z���� �J���
Ƽ)�Ww��/�$�QqJ��'�]\!�q�={�͒5�A��N�w/�1^�V6z�j�ݩ�g��e5]�i�8Պ冷j\aLӛ�ؓZl�Z�����q�|�@��Zձwch�{]J�3%�����Ճ�̵=����>�垩�-�����f�XmE�ٵ�nq���n�s�- -!Z�ў]�l�26���90�����2���℅�Ŋ0\��5L���K'g���K��R����Ԟ��
�*�Jz��Y+��X�lJF��hŜ��p�q�f�4�KޜN}�Sɇp��&.[r��]��k�P2��z*��z��o�雲_��1�(uE��{��D�!���	���G�QY9w�[��`�w���7T�N}zL_���n	��ٳGDVm!qNcEG'\�Cڻw�G܎\�bc:��"�J0��gVr����Xz�B��l���ǓpO���B����"r��T�$��C�g9�Uol��|��g��L�x�,ya��:�`�q[f��b��{k�y-�'��bΐ��-,�f�V��NL �p+�W��Ss��R�Z��0�+N�b�.�8Ѵ���n��Rb'O�uH��[`;(�܁�n>����fBk���L~�w5
ɗJb0��K!�?u��q�Ş��`d,�yb��Q��\r&[@ լ�[
'��pz�ʀ�4p�+�W��������w����D��x3��t>��G�R\�{~�M돋��R��M��;6eM3yu�a.0�mr��!
���W[ܗS��~tgQ)9;Une���lwY~��;��e0��"��"X�r�y<�"�D�������orHx�@��os�zbFfU߶no��CD�J Le:b�E��`D�6"EG<����F�r;T��#�ID_w��/��d5V�����-e�7�@;(2j8�(� 2P��kȭ���<Z�����/nH�eH̿E��W=�?�ゐ�ʇ���`=|-w\�������W�9��Yz���q�:�R�*�sz��W��ɴ���,B�1�GV'1�ۗԭ:��w��_uOju*�n-O�k.3b���e�6�V}�݈��<+B!�j�*���P�����z̜p��G!o�Xx_T��WfD\7��vAb:�&�L�Om���]�+5��g��3c	�Qh���}
�B�X���X�N��)�/��B4�|pb��^Z�-����kJ�m��J_�0&��>j�\k���_��񨅢X���Fo7/:�Q�2�&�>^�����D��o5⪼8l$Y�4�V�o�^�;�]*��U�m%����2
� bݍ�:�Z4�孯Ζ�a���Y��V*�W�=���t�O�]3u��O]�V�)����!��d'r9�V�ά��ULhj���c�/�Ν��Df�WOO[]PYg�1�\o�˹���gNC7�4+l��/��N�Q�������͉�9+<�5��s!��՞�(p��m ���XKH�̫.�Q�W���1n�G�#>̑V��Ie�� �0�.���qSa�3��هC�����m�$v��:ʓ��Ra���	���1H�������C�I�d>�stR�&���_����[�u��dl�(V��/ Д]�:��(�CNO���^�<�
[7`U�jz�8G$�����,&�>��+�)
�Ie�r�N�E�`G+��:�	��)���̀"�$*qi�鞻cnn{=G1��B	8y�v���e`��8��'-�]�9�޸�u���,��u"4:�Dh��<�b�z��0�*�{LW��1 �]ΧTd���K���̭΢��M������mm�7��zYEq��f3��CLp���ʕ�Q6�	8Ωm�})�*�d�u��Ο-7�0�I�	�v�W\��������/��K���b�2�ߣƫ�tv���"bK2��W֣�<;8�TNTw��+�����~4�m�ˠ_E��6>ל�|q-��KM���n^�Cv�Vr�G4Z�#�b;�;u������gfn���!X.�F.�P1��	kko>���<����}F���$=�'����V6/���N%[��v�'��K����hAS�2wU�iQ��1aiA�NPb�Wm��E�n2��܌�k'{��'Q��[3䍺��Q�x�"��W�گ1\��_�S�~�r�>�E
�M��S��*l�v��Y1_�Ur����y�����랺�G��3�R���θg������S˾��akh�ʩz����Ҵߥ��3ЧjWd���U
�g�EO�EZ�����⌺���Mt��Q��[�gn!J�>��S�"&ڻ���9�3�zHB�xT+wפ���{�S�苽�κ��pe�/
F3JY8�')�px{Uc�4�\��o�� 5J��9{!�����3�y���0��a�%���2�����F��1Ӊ� �m���4{�j�_fob���櫂�z�b�/t߮���<;�aY��r�v�Pw
bBe@wpъ��p���-�I�����^�g�Xw����<ߩ���ku��2�[���<���]+\9*�sN#]E\�p�I<��5)h9bv�L=DѶ���!�^�{�B&z
�e�4�m�f���}eد-��]];�9|]������R#�J�{i�!��C�w���>V	�����|l�7Y���*#-�K���#����(8��-�� ׀,����n�9gx��������"*�R%Զ�X�R�콝�Ta�>p\���H�:��͏]�v
�aqވ�6��!��W�𫔖V:���
ti�vY�I���,�/�[<&ki;T�Eu�d�C�����
��)�;���8�]��JKZ딽��xP�Ɋn@�q��OR�J��7T�o�8���GH�Ju�N�ral�s�>��Վwsf��I��EɄ�=���0�l�1��^Fٌ��B
U�}��w�%�j[י?k��+i�V�q�
�x<�b�=��w����[��%����Ħ�ԬĽK8o2�W�vBp6u�w2�W��
�=��m�ɂR\�})��-��v�����g3��w�0[�8�o��꜀�^������0�y�ܵ��Gl�����έ��*I��|��{Q��KҬ����Kޜ���E<�w�f1�����s�Wn��ub���(xO^�[ͩ/bW]L� �p��K�u��s����̋U���Ǒ�A�& �J7V���s:����å`EA4;�����mBY���9��pS��Tlh�2�Pͮ컄r�r^�iI�c��q⻧��uoI�,�#�b��)��͖Z;���G%�!��B��܉�c.�9xpN���p8��@�=\%��:�	��Y�VÝ�ڴ(�>�3�m�w����!;�)ݷy#Ō�0�:�z�M����ʷo�F)U#�ha`���ȾY��B����y�:ų�"���Ʌ�B��j���C������O�}%��^�-7(���6�^����t����F���wq�s�
�8Q�5Ø�1^�J��6`��k�O��g���U�+��@l�A�����[�����{�N��a�V�饚�O�G*�^{ζ�p�I1�܁�oꟑ���M{e�� ���iq��5޽}]��Z�5H:��EAc��@kѱ�����Z����N��j���[���t� v��++�ƈ3� ��t��q�^�`Cf�HS�v�+���5���:�&���$,fHW�� f�B�EV��ĥ
xx��x�:��J�SY4V�2�\wN	�W2/2�Y.s؃W�
C�k>����`e�v�1�رJ�����$��nwƽ5Rʯc�'z$+W��u�DŐ�İ�W����y�'�"�+�u���[q#[ʡ���"�pO&���&�#q�oW�a�G�h���WX��3{IUӇr��:�4.��]�r!t�_*��h�u��|�^���.K�ơ�n
�a�LL����ni�k�df�Tpݔ�'��]Y�S96�IoM�bT-�
��&EE�V<�N��oU���9�j=#��:��q����0�/�q�ޫ���VFơvYu��4�"���{����U`��ی����<ʻE�d�Y}@�.��kV��,���s5�#9Ӣ�)��&���m����s֑yP=��k�{�c᧟,{"ɑ��y�+~X.�J��'B�n�yZ��*�t�y�F�#��qT��*���- ��Q�\j]��ɵ�d2�&Z�&���-��ɴ�h��EM:�8�ebU��S��A��C(і�wZ�:z]Ө�<��%�ُ^i�� �\�+�`/�����ފbbVЧ�{E���!���gE�(�<�rMi
5���&�U�3쭻��̗[9g�s�������{��J\��a�Y��ݔ
���1���Q¨�,�w.��[��Y8仺L���EQ_TcmZ�0�/�9C��M��l����+jǍv����4[�a�����2�������h�r5ӛ���cXWV�Y�}ն^��_*ĸg,�`��U�����1%�P�LN�6�J���Q;CD�`|m ��8�ҠW6/�rp�R`�/�}�X�.�����#;�u!�������9�Im.p��n�!�+5����d!g�����1�,�g�S�_v�7�B��j���'OY���⦣q�e�MR)���QU��at��V�Խ��Wf�K�3|�C�lv�F�̮�׷�0���2�(����ER��K�^.�����]�r�v�=�R��]o`��|��uˬPz�j����7|F�{]8�׉��L��<� ݰ�#�{���\8M_e:D*�.�"�w�]X4�k�ͼfViK��x5:�ݷ�o�w���;�jV�e�g�ҭt:���}���+�m��B=,t��7�՛8�Cp�	|	ۑ�/����tkGwK\N�V��!�7�Z��q��7���u�36n�ͩ��-�G%�oܠ�uqP�t���()Zt�¨|���u���j��Ku���Y��@���Q�%�XV/�?�x�v���G�/	�3c[��m��)�x!q L����(��Ӽ�z�fM�F.��&ɶ�u��^j7�#}��{"�7qj}fT;³��i�C�S��
��as���F�uqɇɦ�t=}�v�廌:����pi��j���	�̣�P[�)�}����,4u)du�G�5�a�J��kyi.W���NZ �}����g=�{V�w�6�)-љO�K���ޫQ�|5Л�9���u��wX�O����k���0j�s�n�U�������ANߓ��i�R�Eu֖�]�'���ړ�$��n�\�J��ܫx-�ob��s3;���O�]�7s֋A��֌�w��vi���279ܷ[q���
y��3F�D$JI%^���,M�*,+R���)uf+d�Z�����AQY-�"J�2�P5VX��1̰X��"���P�ʊWYcR��ZŁm\A������LM2�2(�fXc(�Ŋ��@��lu�bE�VQY�Z��#P�"�L*��R,�]R��S��[Z*����e(�#D`�K�RWH`�IZ�A��`��"��P�YZ��Z�V1YVV(eh�Z�"���Q*Q�Ci*(�,��!��&2��)ZE6����J��D�1�1�ܠc1�U�r�31SAeL���k�eAt�
*�"����bA����_a�W	do�"r�o�tC&w�I����#��ќ�����{h��x$�i�� 3)��2}�ӭ0":��o�e�[z�oJ���-qT�W��
����p�P[�u:��ّ޳q���*�����^P}Ky�IX��U�L͆M��2�2�9�*�V�b���'lu��aB&x��֬:Y��gv�H�Ԕb��@#J�,������eB�^��
��f�]�xVՆ=���$���v���5e���RU����31TB=��������C��i�Mf�"T��jTt)S��Q��9Cl�]#JG!��lH�7T䬀|����H_���vb�\8m�Y��t����Jw����,���c�;Xf��ۙu�:���>~~�|�ClL��Z��Q�!rX�wh�p�}fxe{gYw:��U0ً�s8'Y$���"n*�8kCv�=/FT�y3��17۝�1�Gdû�f1K����E
�s�X�Q}�!��I�z��-	���>���33����U�e�G�G#.��Ə���e�r�NN��4ޕǵ���9��&�� C��$uښc�ĭ��Y.}���K<(�c��$�	t�����w�=|j�6j�-<�:�x���r.e�^ܿ;�$��RޣX)̨9ŻB�܋���˻�6�&�NK��\��:�i��Ц&ɢk\�����Ý+u���R��3(��u^NY�$�+�$��3٦��hui�c*��3��v�<��F��9�l~�"kʨ*��F�\�$�<��)g�,��^b�i��dk@�-1���]��邖lz�Bp�'�\ܴOm�d�rI���W\���Ep�t;�O[�B�[�v��Ȼ/�HҮ:b3Kd��W-�iևg�Ϸ�'�G��1F�*�~���Z����WuNv-�k
]!ĩ�$�Gb1�k��tv�|�J�a�Z�
��xd@��5��=�'�cq̭Zc3��@��ݘ���L�]�@�{*���iQ��u�(0��k'a���W\�޵�\��A�9�)+=��T#>H�1c�l�<�ɟ0�mB�/	�5�r{"���U�KiY��)[/ҧ�)I܄�f�D"��#
�dߌpH�]Js׺�#���s:����^~G5M����Ҵܷ��)ڂi!#��T+3�	�*}�#�3X��d�V��Ρ��:}S�W�a@��oϤ����l38�P�=$!Q�¡'Z��*���̦��(�Wd�wXPC���3J���r��t}���>>}����W��$��j�\����rjӍ��rLl��g%�$*^r�����w�*��W�2r��x9�PR����N��Z��i��c����kk�1�,|Oc��꾑�[A�]�b�W�'j�|T^{׫�I@*��$�Ns-й���V����S�D3х���i�ݒ��
����	(E�A�tƆ#I�u*c�!;�&�ch�WD���H�i�~�}E�sT�O�57d�Z	)�]d�l�m��2�1�Bw5N�{Ԃ���왙��uqv�ܓa�pؙ�8_�r�];%+�;5�>��J�3՝j�Ο���m�6c�2�j���Q�aej�L`���
�L�Br�
�����|e�4]91K6��>�
�Σ�IL��*�u^�p4�I=��b/bgC+��=KH����w�v��X0(c>�\x��o©�]�g՜��m��<X�UA���0��=>wͶ����^��̋���y���P�^LP�@����Lu*d�%�u����\vJ�i��W�������}�cY�d�M|�Rf�Q�cO֦ U���_�R&�f2�P���y�qh䀣���E�et��[R5183�xMIί+�T��`�F�UW�ZY��˛�L����/�Ӟ�:"��/ۮ��W̍�r��|���Is���tw��^f��%f����J��Q��I9Q��fd�]B�!Mq6P�b�u���͖nD_������CQ�pfZ+�r�ΘŽr��V��P��,���.P�)��<�θ�Y6ZS{A����zWR;�0����\p��s�j�zpgr���E�����8`#~�O=����T�a����츎[jN��<0�����͖��ك{��+z���Xp�����uҴ�u�Z%�N'>��O&�0��]%T�p����VX��xb~s[f���d�o P�#0��,C�w�� h�p���M�tS�kݦ�:�kC��Gܺ>S\w��4��Q���F̓K0J�%�p�\6�zͤ.�Ɗ�ru�J���Kh�������u^�+6�C�N�z�haW����/v�Y�y6O���� �;k�`S��.U�֣��ɕ��Y��U��o$��!U>\N�|�>Y�^�ݣ�QX̔%�$� �!v�U]-%+k��eC�LgS��s��j n䓁OQU=�}��g
��O.��I���י���<3�B�DЉ����2��[`;(����?"&;�oх�*~7v�'���5�;��(`�'���FR��(�JD��D��]����":�2�����>��������0���|��gL1Fv��nm�c�� ��L\q�^�b�����u}�m�1�Q�*�TU\]%o'��2��g�rWj*����ّ���0f���Ŋ�S�*���vF����\q%�E�E>iMJO7��odxާ�M��i9�T� ��57#���9�(u&���ɒ�-뺾�\û[D��D�r��Ԥ;;��pR��j���#ny2:��[*��u�&2�YA���b�A�Z��%��=
V�K�Tl�B3��ٯ5�+��d]�)�&���Z�|�wvk��*BjӽƶO�C.g���>ڞPmy�'_��>�'2��=�b�v�J%��44�Ǝ�j��h.N�ԱT&�no��U�#��x=�����}�RImr�M�]g:��\�،o*.ˤ�ٗ�<�C1�-�A�*�w͋�|��Fo	�B�+<�9j���w�{��n�j7��ɋu�h��'q�l9�2�R�Ȣ��_5��]O�-�&4Ћmok��}�����7n�E\	S*yO`�����w��Ƿ]gJ��d44��s��#x����|2|�\�rʱ�TF
���v'�{ȟ%m|���x�s0�5=Jm^4��k���J^�Lj{FQGGAm+��j,+�/
nX����Ƕ�OdJ�u�$���b�w���k�$ia��ó���\2>�W�6s���e7t �Q�+v�ʋ&����K�/��O��y*�O_9�s.u,���jQn�ӽh�ܬ�L��B�\�}5v�H6hq���t#h���j>)L=��R|B�G�\����*�������7���LpQ���NN
��q����q���}��/y28���j�;s��#Y� ��pz�>����2�����oDV���k�ؕ1/޶5�`k�v�܏���}�L:�@X��:�|J�9x�"�F-&c�E�r(e&�(���ⅽ.	��(S	�;Gָu�#��룕j�2���LQ�;�i��}ued8�N*:���Ǌ��b�o�Lu�6:���Ok��1�9>�S���\�_Fv���L)lbx�gJ�ӱ`�C�ٴ��H� ��s3y��
_O7���*�X�5�V�&6��˽��~�k�7��N*5�cht#9��ͷ4g�:��Q��'�F��j֧uR2����cy�"�
h��vg<��ʄm+sYD���W%Y<�#��y�H7�D����V���ͷZ;����.[�nË��̽��kBBt�:�@6���y���ˍ�U,\�*�e&{;����Փ-b�(�ˢ���W7b�g.�w�uwk��"C�Q ����S�D�!�J$���9�w�UaË�Vsuv'�׊�W�q��R
��*ؾJ/�q\�<P�������oս�Cη�kżv�"��BU�T��,=�7�3��{�V��Jx���e�c鈭�\�����[�[V��U�	OT�u�Qn��>ĕ���T���|��Vj�Nc�����U{�=��Qq�Cn�U�{��*@|�Tu!پ*��hw��~�Sw�ށ�^�f�O`~�t{����O2�kDVt�~�+���n�걓���W1��ҕA�g��=�ŵ���{��Υ�>��
���fr��8֛X�T+u��`=�dW�m�(�1�'�#��~s��X1֢��+ N^,���NU�|:`�:rC��:�ل�Oj�{�n+ء�wN�7O��r�>��2���&�j�g+ԓU�VeTZD�b�-�z:���=���A{[
�r9�kǻ!2�;��u�`�Wl�� �v�c����^�0w65�IR��-��ۍ��9�9p��/k{��uf���4�K8C�}]ǷE��oٷJ�p��W�gb���|��Tmȡ{@]q�����Ȧx�v,��"��*�z�_a4�+2�E��g�)��hW�V1p��z��seҕ���ƻ�2\F,՛݀���-+�-��'�;��+u��匢#<R���q<�çf�}9�q��(6� ���m��':�����y5��6���j��/��ŕ�����in���׈uR6��@Cե纴C��HeN`{$�v����*��W�<�6��o:
����1�ȨB�iCV�����Į}ϖO-V)rqr�G-U���hyɼ�)�Gݞ�x.�.��oM��l�	��l8�W���].��-�Z7�ꝲVS��V5�N^�^�V`�}n���	]������\�֯Vj�D��wS=2�D��ז]���mV=׫/�h�ѷʎy�e{Z��+���:����u-u���f�ESn9j~��N^��F<I[U�C�ԇf��3�s{^���sj��9e*-h7y�'d�
��!�:��e�{�ԷJ���,�w2����:j�����Z�"�r���B�"�n�#��M\�� I,�;�[ݕ7XΩ�����oG�Ѿ��z���)�W^������c����o1�Z���i[c��CS��Q)�nr:��&"�	]��k0P6�|B�L��O����%'Q|G?EX�Y�૟lJ�b_"�9�t�-1�og���o�6�Yms��;�r��漬1o	�b�v%O�r���9>�U���vˑksB�����'^�;V�=Y���>�%����" ���w���	i�S^�j��ͯ���C#��l~Y�o/��s���Y�qmFp�E���+,�|����=����[����U�$u�
2��~Ɠ��u��P*	��/���W�
��OUs�6��1��L�$�f��R�ҫ"��s��u��kQ\�0�s�И\�\RĚ��}�mYժ��u�	�1V�%'��.�Of���n���U�R��|�.����[����k���i��\��Tͥp�����'���{9jy^zv}Y��:.'�1;3.�-M���Y@�DV�qJVzwW:�	#B�tLJw���L���Kd�ܡm�r�Y�Qᅨ���u�)\���#���z�6:��N�ܚ
��kU��ξ[tl�hJܠ�v.x����Ρ[>�	��*VhU�ٻ�+����#��S*B��
�e�Yx��- ��#:������/��|2[v�E\@ЕW�W�ܶá�C����"��X�
ŷ�Z����ע{5��i�ɶ��rʿ]�K���~��k}�3@A{��q����]�#7��s]y��)�]�f����[CV^8u�����#������l󊵐��J���n�:��6m�G'fi���d�@Y��!�s�0 Nsgmd�ޫ8�hU��*u�;�U)���`%%��C�"�+��r�[�f����fzhx�^֟-V���~N� �V���Ú�R����MӅ`g��P��~��W*Խ��}���t3�}I1�-�UuF��b���;G�k�ֈ��9�Pr�w�2ca.́.6���Z;C�P��Y�ޗ��v}\�ɷ��ÿ5�u��$�	'���$���$�	'��IKH@��B����$��H@��B���IO��$ I?�BH@�rB��$�	%�$ I<�$�	'�!$ I?�	!I��IO�BH@��B����$���$��b��L��<S� �� � ���{ϻ �������H(TH��8R�L�Rܳ�	RER�R[�;�{��4{IQ��v˩p۩��Z�h0��t�l���e���-�m�ٕ��q���/Q{h��lSl��Mxܗl�ٵ��E5S..�4SF[kkj��\��l�lɣM1Fr�UhdT�&q�'L����<H�    ��))� 2h &�4� )�)J��      ��L� �LL&4��)� ��S@      )�%J�� �4�#  	��J&A444�45&��&�ړwWO
�ê�4ED��Q(sDi�A�����E@*!��"RDȓ������?\$?���A,�J�>4d�DH�D�O���X~��}��,�A ˊ9ܨQ��P��7ю|����ơ�#;�/�[�
$7C��O�Eۘ�k�!���:�V/�A[4yzhu��Y6(�<�V`#n�vrِ|�^'c]�6���ܷV%۰4�v5cv��(���t*��hjT���u��*�+�[��c���p]a1lW2!%e�����L����mF�f�W��*, �G5�ϴ������O�a��XKq���k��yOw�`��wv;�؃#��"�@���
�s$z.H��jӇ�aM�Gf�e(�/]H��4[�˛�n�Y�ʘ\��W���,lv�!\u��l8�6i+��lg�I��l1TfU�4�*U�xʽ�6�l�+��ʤ�K�ׄ� �-t��R-`Ș
�������X�nl�@*�E��W�dXͳSl�-;6(2���`�yZ�Qf���;�s7f��[-V�R�����.�b��ͦ�2�@�ؖ�9�Br\H^��*\���ے��_̄V��*����8�ᗛ�!h��*��٦����W���A#�K��o30L��㵊�5���nPb�H�̲~A��Z�j�
�Ç*E�5�Cr�%�ڳWzr��kR�
�D�Y1�2+&�ߴIp��[�e��T:�Ɲw����CdP�5y2���$�-XX�u��<o]rή����xx2ãԴ4�����Mձ��MkY�tiG.���jr��Ǧ
x��|NK��� ��Xg���&�S*#"�61�9��)I�+*$-Y�2��nވh�ZO"��$1�t+W$39sH��%V�em�v
r������D�K9n���-���4V�˓/6��^G1X��v�c�(�V�W�6Xi��lU��z�b9���^⊥D���[��D��U���2����а��u����sseCI�{�pL�$ɹ/�^�w�fP�����`�ǭ����CS��e�A!˦j�;շLC�J�"��__,F� a[���]*B�~�����{iG��+��Ǝ�j���p�Z��Bv؎7����)}��o��Ģ��*Y���0a!�{�˛��C��j@��\�gi)�l�ԕo�4��E��.�&�J�UϺ.lJg0e��y�r��s�nH�0u�|�r`ի���r�K(J�#���5����5��{�ޤM���Гt�:S0a5&���d����4�הa$^io��c�尲]a�����"�m��D��b�Tc�o;/���N�C��vy��Nu;����>�GN��|A��ٵ��N���3�Rn��s��+L�QU� ��,^u���򖬧�×4��"�֌��\򙳒X��z�1Iܻ�bo#�ە��C�je��Q;�K5���*qU�t]�5�L+���A�\+�t�e��[h�r�ZSi���$\�,�����4oq4�\�}�w
9H�V;/>�sri|�O��I����m-�@\{�B>ۑ�[����L�*���2�3]g��o���U�v�K[Sh�TAI0PeYS�	 ��B��%iD�+Ma�-1�	�H ��29H� �n����˾��r%��2&�&-� ��aj��
��������R
,��zy��q7^��I6q)I.�w2ԑ�<� �*�1�0�Z��@C����n�s¢��=�b6�iރ:�-��=��Ѩ����������Jr0s
��y�  � �       Q��պ=f��;-5��I�Y�kM68�E��Ċ��6=��(�s�ΗL��V����2�К3:$���L�CN�6T��\&/���c	�ͽ��ڧ�����X_8v������i�>cg�\�m�㓴R�cT�3Q��t�j[��n5��#+o�y�5����lou���,Ҭj�U�K'X�G^��t���F�dSY�R��諚UF-��v���HΫ��p�9k"?nq���u��L�1FI�%q�6h�g���ٹ\�;)��7݆��z�ؐ���m�uT�4�d���@:O9���_~�_l�ɜ��O�_Z��S<;I�q��;E�r�ٔ~M��u��=��.�z��N���\]�ӓ8�cm������ե�Yz�����#��V�7��F��9�h;\�C��:�қT\�ug��Fdg�n��" ��f(/pLWq!5��F'A
������PC{��$��9�l-�2�f�}���]��8�S��G����]��[7�S)�X�(Q�5,���L�pX�`T�RoBjڢP�~���}��u���Ŵi����Ra���S۩W{H���eJ�Z��yv�V�i[/yQ£iT�p�@ahV��u6dv���\�����{���`�[���$�6�t��҄�K��h{��3���=@Q���C�c
�����?>%��{*d��P�����&�!\:g[�i�]9��x:��똴�P��1�	��_�n�����E�[��Z�c�
!f�t�y3��a����p��k[T�5R�&p��/���Mk�q���#���\T�e�b�yf���_�:��Gi���cr��6�JB�<�j8�����}��p�?#N�4ѕ{]F#�<�rK��tÛ>���TU�����P�ᵗ�;V��d���B�n˒��u,�ʼ�g�>YH�f�є,�`m��&ٸe�k�mCN%���2Ҿ��خ�X���6����h �H��n�lE5���]̓G)H�e�%`j-��v�+zN��6*o��Ը>M�sEcUjv2t�T&�f��&e�֥zMA}��{&d7��8��]m�7L"�wϰ[f������BY��$=��W����a�dl׶�F��3U)X<ox<v�����2e��1+���c`��ic���A��]��圙�raU�Wq�Ɔ"(d!P[�|�q������,<[r���Um��)��c6�lTLVmF�6����8�a �	�ޅĪ"M5�@�a�V�3��Q?;��|e
���!^�)�6)ɛD�+.;2��2Xw8nj�y�
��a���a��� *��B2�=�!T�5������;��-�f��ā�H�hФ**��m�!�c�d�T��鱹�0�zȣ�����ӈb*�]B�䶰�2B2]���#,����=w��"?\�pe�贤�8̳q���4-�/�r&v���F��Բ���bz��h�k1-S�:{�ZC��ڶ��^d��-���W�:��@�y�k�M=���W�Ԩ�-��ی�0�j��n�����J1�$�{�G�|�r�4D�wW>�?8��?~A׭�d��R=�X>��}@Uwo���iګj�ˬC'l�O��ҋێa����~u���ܭ�X�Zk����|��vw�E��O'�hԮ�P����kC+\�%cA�&=�7��V\6�����+���j�����M�Z�rRL,BF������v�f�[j�o��cV�w
�u��y�|񪴮�쯝6�ךӦ�k���Rƶ�D��t�B=m-�ѫ��ΐ6��NПJ�4��4�:��=��J��A���l�1�%]mާ7{�헧9��{�'9�/o)�n��>�cU���^����>M:O�#~�֝�ݡ�i�8���^v�� ��v�[�Zk��s�:��ZW��w���[�xrt�]�#IS�z�x��MZM�l�MF�Ω�m����'�P�P��b}�+orQ�Y�7���Z�4�5��
OΕ�C^\�kI�Đ�D��(y���$��ظ��F7�Cu#Q���&���öa�vǮ&ˏ9Վ�+-i����]-EHj�[���_��T�۰t� U��z{�����'�ԋ�9�.gl�xSPl��kǗ��i�(~�Ji+Q_X3ʀ~��̜jWAI�j�n�v�"�K�P��7��;n�Y|�sj��h�%a3�J��Q���ŏ�!����mc��!��G�I'��-yZ��T�#^+����o�K���벴�f3�Te�C� s��Z�4E�3TF�T�[���I� {�	i��Z���`y�?���{���QZ�wձo������y��㪀�4�2D�j;��>y�F���1�kP���7gIS�Fz���i�:լhOtjȱ^��q��;�ɍ�kz�w���9�>?&��?u��<;����A���^��H-K����k���l�m̼��.���o�7B���ˏ��-�.���.���&�e��l��z�3�;�<<�S�f�a�u^�l�V-�η����������?�߹���h?T
<�8ʛ��͌h*Y�49V�Y;�mjZ�0��c5�5H�vm����+�nL�9�s'k���Xe���D���^��-�BѸU��E-�X�.喁�KT&^6f1X،�.�V����+-am)�DK\�RK��\��ݑ��.�Q�*�̩j�5�+ٞoz|-5-���2�U��C�.d>�o��f������V����h��3��f��4�����7X��H^.����	�U)PU�r�;�����E�*G��ɁH��h����:t,V8�+Gɂ�$ןA�WH�[�|��1Y���Q;=<�,oY����Nſ)=��7^���{����{ѸڏG��}���Р�ND���ϼ�;fLYPS���lTwMq��_����/�WlVh{Ӫۻwx�5��;��o��8����eu�.壧���۞�}l��jdVab��8~��p#k�0߁�̻��w��*�W�gj^�ج������>�N##Cs?y���z��W���a4�^Y~Ϻ&���X[;F���OY^<4�-����m
ڪ{Y?�t��l�e!:����}�-&:���Sj�Gʋy�t�eFc��?b��7W����El�^L�X)
��?&�
� �yw�r7J�?�9�uMr����a�~�5����]_�S�$����{�};���&�.=.��b�8�Ľ��e�S��t��hQ�/�A�zز0��h���-~�A���ߣM�<$%���k6D�k��צF�٪.�鰟5�($r�����1���w�T>����߅���̤���`���\�k�����c=]?R^|��F��;��d�Q�x���������(�5�,D/�\K�οH.�f��hlb�w(͈�Gg}�2"��g�����Vޜ=��=���=7B.N
�L����Z�HIi4=O�_����6*`V�3����d��oZ��=�A���^����.�{������Æ
�����r۳�7iѦ*��`�k }Ǒ�ʸ��Yd�g�F,w_�����~�)^;}�H�-M�Ab���+i�Y(c��p�z�y_}�2�f�+I�0T����e�&0���C-Y�5�r�m���Vό�ma����,@�R]�B���E���Q/���)��坧��yyG$K��ԯ��҉ �	�ʨ���j��*$�b[�P[�H�,̙
\c�bAU���)�0Lj	mF���Id�v��qV5v�܂8�̖\��m��$-"[!��J���J�j�-��V�V�ZT�_����^��e��H�w�r)�o!X��1`RS�_�M�2_��uC�S�l�W�/1�}$c����c���EuO���}P�&Z�cִ��~�5���_�}w����꺱���u�xк"�_M)Q>�MM@��{�yj�h
�D�y�w]Z�S]]v�8"o��[͔ך�c�d�{Z��	��z�Y��,9x����pSKu�w�P�W����%_�R�f�"�1�A~�t��'ӉJ{�tq0-�T�T*�nے�?⼦K�2ݷ\1�^]��xto0�����=����!��zx)�I�I���0�^�۾Dg�Fe�i��L����m��i2���Caù�gW���;��o��`���=QWˬ�F��Ǻ����<���V��4�k./ ���G�)3"q�&g��_!�����f�ڤ��ydS�eʼ����}��{-
�Zqk������0�C��l�ؘǷJ�Y��N��&���Md�,y����+K�5�q���x�����N�������Ĵ�IȌ4f�1i{3}�	����}ix����' �ȜN6������+���Z�y-������C�����2����lЭǩ�a��~n���͜�G�>��r�4�2�s���\���'`�x�ډ���y4�QfZ;�3�Q����x��/����*C��t���{�<a�w۴�U=�/s���}8ҷr�n��p����P�p�=��YY`�R����-o�Y�|Fn��5��f��
�B�]ԚPCɳt`���X*�V�Y:d����+�V���s]h���1�L�!���׎�n=��)�m��/�Jc��}��k��j��Y��C\�aE���f�6.n�S��(���3\ye�*q<������
ki�g'E}p(��tQ�$⨤��Nm%�{l��i�ej�[&0ĸ�4h�
��H./C5��[�'{�/&t�����N��*߾#�"�a���*҉�d���ݒ��j�cJb]!l[�-����LU���j"� &0�����,�DRd�EK����e��q�A�B��՗vH0#�L?"�����5��6�׵	,>�f�I���g�'�Z8�xg����;�+4�VY���>�|ޫ�=fyR~��,ZfH�<�|�{m��2��Y�:mi@#��ܬ��y��z����k��Qm��~JZ�j�9��H�J>�k�odx�2Q6U�ا]m�׹�X����ՀS�%������oMF�/q��P`ݩ��m.'���ܿ;��o��"�gi�y������Fx�ZJGv*y[M��=wxLbmZ����/J����.&kҎM�[��R����[�Z��S��T(�͟���O�_̓���9m
K���3��m�x��:f4*�5onVп/9���^L�[�f���C.s+l��aN�j1{��q�qﾇWW�9�ݪ"a�j�H�~�]��/G�y���䃺'B�4�Q�>N�cq<�j�*�y>=DK.�'�In�(��^n7�h�v���[�s�YA��Ǒ�������Q���(-��[��^mo��%����BK&+苐F�`ZQ�=�33NyDe-3���<r���Ս?!M��7���o1���ג�m�Fŏ\.���N{˃yH�6߼���k�cHJF�D�d���3q����O������m��v�����z������fmk��I|��Q��������ٻ�z�ڵ�+���Nf0X$$��s��Tz����\�o<�V��@u���4���eŮ�7�n�P���ޞ��V�����񣛸8BuNv���Ew*m���5�{���\ϟ��e��'����Tͪ�Jej���s�f��k2o���hP@5��L1���T�*e@@�,��7���8@��*^*cAK��r����!�--2���*"�"�*9�J�Lc�3������I����z�;�Qc��ŝ9��TǗ;{�=k�����.PnڝxV<F�Vd�jR\�nsVe�ݭ�-6��cT)������5%�b02.2T(�k1�c�`�&!���/'�5<)$�9%�nh� -'Y�yz�@����R�V��S�@+iԥN�d�<h���H./~����g����_`Y�ZSe��z�%�r��3o]�.��.F��m������Am��u���#r��!n3``�Ww�DjJ��5�G,�kuF]��t��j�-㼳�44<�k�w}��<j�+���7.��
n�t��`�"�⦗����V�R�[�
DRռ��1R�R�T�".�WX�k����q�ٸ��\n��p��<��cm�u�i��|)mz�F�Q���~�����N~"�pu�3afVU�Eh�q���ԧ7䐆���ޕ��Y�x��+��v�do�<�Y�ݚ啔i�K�[���p�݄!5��|
0q����^�tswX�������2�;.�u�#g^8��^X�O��NEu�I�����������g��x�#-$��Jl��i�{I�v.�5������j��8�U7<��䇉���7���O��;KU�	�W����r�\���:`je�'�e���F��x/M����7�Q��v�n�1�fh�E��s�s��)x?��ܿ~ِ�
��]��|9�Q|�����\�|d3bb��\���&�%a�5v�
[�bۗA���wX����Q��s��u����e�ʣ۴Z3$�6�.l>>�'Ek}�ׁ<4|_Z5��j�L�y��q���8���U7�CR��4�[v�8-Zo������_��t*ƶ~
�o�G]{~ �d��%��A��]qJ��W뭖m`5��纘�E�>W[�ǹ���O��z�ME駸�ː�
�.1��7�>��]c�M��u�M7�׊)�a�[S����_��~�LH}\�u��h�/2�Ӧy�9�9�Rr5	Xy�����l�b��}���������v���K�`v���,����<��IhpR�˞8����Dz?���rel�xzL󫷚0-(=��5e�|L=xy+άY⯶+ =�:��
��/����B+ſ6}�Y�����%�[~P���E�EfW���ߪ��
?�^%��!��% ��W��"��W[���;�A���c�})u��/8:�am�&*u˰��z��h����Ƭs��/��F�U���{2d�ęvj�|�x������nG�w� R��������;n)�z#+z]�n�=�V��p
�u)PL'q��	Ff�Qzo#)��:)b6�j��9��.�5�P��JձZ�e�j�H��	@,Ah�J��l	"��-4�
"%�dE��A�(�����߄�5�_\ffW'[�|�>�&�����%��e\��)|ìK�q�����O�(��a��kw����GV{�i����U��I��i�h{��e{�gjm즬/�OK�3�bh�Y�ױ#J�׬j��G��C�f��i�S9VՕ������3�<ޓ�oH�e���qɨ���5�>�S5%g��ݫxٝ�����*m�u�=c��ڗ]"q����s���hZpxw��i������d̮��ѕ HX��3rc�����1:e�{:���$i��+�V��m��^Cj
3���b¥zW3P5�#!�����fUT��{޺`ZP${�_V�����qiE$jr'��589
��sq1k9�8�uWy����.���y]~tn�qe��y����i]}�i��c�Q����T�SYt�q��[H~f�b�S$�6�u��"����!��u;gS�� ��6��}m��Ө�m��t�f�j���&)Q��ڟ�����4s�v�$W^�jY��m�5�m]p�0W�Z�HW���ɉL@��5��t�j�v���~Ex����v����_�j-�s���ޙ�ֹ�������Ew�<�e`+�>8��,O����3P���X<.��'+����q=��n��]�z1h�z����;���Q
b�ФpH'&�c���y��Oc�^㣛���X1fkO(;�e�]��7XI�Y�sս@����r�)��wZط���eN7����M��E��ѕxã�ѫ���TߟD,����_��k���iU���{~:�Q�.��� �E��b��ЯE@�޼a�=9_Z��i��E���Y��&�ЌN��j�4��Y�\�	�u�R�a%����
?7t���2�u�.7(G��$3��D�R�.m&�c�%+f\M�&��$\�5��^��E3���&���y� *��6�40�([xk�i��^6>��}���a��C� ���q�l��$dX-EI*+IBl.E��K1d��D�R� �[i&f{Ϸ�{����w�U�\���}W��滱I��g�2�~�ڥx͘�3���[��X���M�_�gy5��^;��6q��u���ci��H���NW�\ϻ�q�k�z�Ý�2O��B	W-�ʲӁ*����ݜ�~�h�)%�Oр(QxoY5��ޣvp�P��S(zH��$��gg�r��2�#��П��Q$��D!��<���7�o8��fs�/{۔{���P=��ҁU6>�c�L�@��t� ��:%�n���5?}�d������k���眹�������>�n&ۿ5D�a���Ѩ19"�1�����R�.k���]ݴK�_\�b3e�v0ҭ5�5ŕ ���x��̟�:o�ҬqF�N?u��ʿw�֫�����̇��(��~^����j�Ig����U2�Nr�~�Ȫ�����{�_�7�`���~�Xr��(*��c�
0XB�5}�F�Z���r�5Ƒ$A]:�f��^\���-ؾ�E�P���U�z�n����|w2�
��_��J��6J'���{��68����>������S��h[8�+��TmE05���^Xn`��`4,�j��=Wj�ڝ�{=z��6��+~ݚe����M�ێ��Q7u=�L�1\�%�j��s��;�OX�N�͙1r!�8���W���B��~�RM;���^ݺH��O��jv��{�yP��^;����l6&�O]�����f����!��By�:NAi�h|nq�+��J��������B��|n��Ўc�0�X,>u�Yf��o0������>�y��&�r�o�[�~�7�?OO^�����qe��4�l*u��
�m��!�Kx�D��\+:���e�WXD��T J���DN_K|��=�/x��P(Cˤ�(��&�_;��iݦ��+x�Oi}[4�Q�x������=�p4��fJ7#����U>�n�;Ǔ�Rm[[!��&��L����7RF�f���,HSteH��UM
2l�9���X/#�T�,jH��,c$B4Dc�������JD˅X������=��4�7��1��{O�n��	�g�B�U
B�[��z�߃mz<��V�p���Ee������x�zuI���0땥�O(�Y��!����l��W��L�F���f;�3[z 6�Q굪0�6�-x��رE۳y��)��̢�2{5��Y"�ȷ�#Z�~I%�t����{���X�ޕ^��i�UnD��)�J�?=Xjٯ[�Jz
�F����;�+&��/%C�(u�8/��_�9r��MmMݖ��Zt�5���ns�Pg�@'��q���G�3N�wK��YG؋zl���s(z�7=!�^�Ϯ�Y�i+q�Tr���zM;y��ViǶ��"�i�i��9˛C��V�~�>��nݦ i�z�>\�!0�
8�̻��Ǎa=�>��Ͻ��J����L6ԭ?^�U�l��nk�:A��i���_}P�]|���WT!IE4O���}W���A��^h��^Z��)͋W'�	¯ګ�B�T�Yٗ�V���w���#�-���������Ihј|��Z
����|{��M�t�cK���������8�o���j[7�d�I�K�;���`P]=w��iuKr-�`�Y#J�No��
^��?U�o�Y��n�'����#�?s=x�����j�-�
�f:�B�N���!|��{j[�
��ln��.D�2<���N�\k�g�:q�B!�#J�MM�;w����֙~�Ӄ��p��p��HQ\�n����83f[Y0%�%`��/Ty�ĵF��(�G"+���'��ؠ����2�0>�nJm[�l�nۼ��O��y���}�&�3���؀ۡ���n��$�&�K9ȭ��寯��sw7��jW �S��Yq,�7J�m販k�poq7�dk�Z�z�̠�3��)E�wur�/+��h�����ܱ5$���n�a�Fs�1����,p�Y$�뚗F��Ak��ړ0)MM��vXNC�A3 *��H6�45 l��VH�+Z�P[X�̷��xx�UuQk�Ulh��AF�TH�i�E��Q$�F�K���˼�_�E�"�߱��nr*���k�|_uO��X��c�������-,ś��#7}w�&��mC*'�+��zR�t�(�=jW��'Je�K+�䜿{tV���+J�6kJ���`Z�	U׺��sʕ4�4`���zv�/iP��=�SP��瞋��ע�F�,]��O?a��N���=0x����肗��-V�N!�l���0eF��B��Ne��6�i�>�z!��T.D�(��HWz�\h�1��& pfJ�x������E1�J��>�Ϸ��U0�"�����Z�+�fEWؐ��W�%5C<4��-:LȚSu/4p,y�k��U"wʺ����P�HP�vޞ9<�!tɧ^x-ͮL��Ku�E�g�m���x��2��/8MCQ9��n��?g��&���/:�+���~�{�F�;U�;L��I��R��K��AS�x3��,/{К�.*$ʞ	�N�������k`6�"��Eu2�#<>0OmȄ)��̬W�����傄���u�P~Tg�(o��,4�8�S޼�>��Or��F����%Z���4~�[~ֆl����k��k����"|�C�㭓�I��ԧ�Y��n�
��,���U�ν�>��8T�C~o�G��x��Ʋ⟏�E`��*��wVc-/NAm��t�.����G����&��i���c������Wh�Y])�q8�o%��p��ʵ�
h|G7�O��^�w1bkO�޿�~� _�Ի�{�d5�:�c���_ߩ�w����"����ˈk#���N��x�b�E	���!�&媚[w��Lcs���-�N ܐmL�U���8��g*wwiT��\R���:�#��r5�.�U�t�n<��L<�ij9N�Ƙr��nH�Z��0�AΈd��dQFKcr��f�75�SSf���c	�l&`@ vn-��a�,��*	�ۙ{w��_Y����ƿ7}z�PV�4�m[V"IR�U��mcH��Ր�� �-��0��|Q}DJC����������ѷ?W��?^����-�~�E�~됊�u��:����0~��y��l�V�����ٽ}�]զQ��·˱yl�O(R'q�~�1xz�g��V>�7�ް6`���R�u~4�BC�;�g��u��j��ʼ�7�Q�ODxM��5��=O<P��,dP-5-\���4ԷhYCZ6l�j��+M��N-��ca�n��-y��зB���My���W����w]�|����VvwJ~r'
��찎����P�݊����^����[���:����c�=̅"R�~X��\��y����	�d�޷�q��Ѹˎ���XΩ�LUQ��X��ɼ7�i�k�.�Lw������i��G�_8Z����R��Ɔ�]��F��h�mbS6����U�s�}�/9�liMa��Gj��^q+���y�4=�X���%we���������FH������Q�V���*�����Vk ��߻��%
m�i��_;}J��r�{]�ǩ[J>s7�3���Z�%�D�������6��>E��J�V�8��J�Zc\���5��'Ɋ�M�(�U��`���W���Y�p�ί@ˑ?s~�e���A�N�G���j��Zq��Lk�9�m'�=6��C�TkW���u}�|J>k6�������aB�|�Y���k�^4z�t8��[A�����6��4�)��ʯ1��*�T4�Q�Ӵ4vW�>�����2�W����W��(��.>ԡ�1+F��j��D8��X֟�iX�j��i��hr����Bvq]�]Km4�(A���Ū�i:�ƻ�ݵġN�[�>���ȴ[A�L��_%i#�m�������d=��z������s��3�s�0/We(y�in��)�՘����iS�������^��|�Ƽ�tm��ַk|��[]J#_^߹��֡��+@��?j��Q���@-��w+�c�4���xѾ{�Ƭ}�|�R��l��$^�܅��>ܬ���}��ݷf����5�X�U�=�|�4�J�7!�˂�ӂ|�'�"W#_%j���G�R����e8�������bs^���)m����&�%
Q�<�wvy��V5Ѫ�����Э�e2�4����'����))I$$�I@P@+(s�����B��( (��HF�(`h֥��je����0�����'�iQ�K�	���T�EPP�U@T�$��1�SZ	��#GV8]��A���M(�a�b� $6�b���Jq����=�l�P����B��z�xJ��7��9����gj�׿8��
*T6h�m��c� �|f�z�.t��`����A�E��I�S�:?�üMJ@�?���C�������u�7���^j2�/ P@2���}*�a���T1i��c�R	w�����B�L���+)��R��n�m�����q��\��]��59�;�Qщl�J��g���^�.�sfH����J�R�1iP�[���Q8]��`l=@��j�R�$�hq.׀6�q0�ǉ�P�R������,����%���h`{^gحo��������!�A �p�c�P8�M��H�9sCwҥ�����(Tt�Q�Cϰ�_2�=�&K'����wd�m
�{��<�M�5@7Y3.�.���{l�6r
��� ��:�B�iA0�
(aW��>��T!�K\S��%�Tp��\�͆E��&����smTQ �\��	�I�����LQE �E�A��D�t�Ç�et�`^���@ �������G�5�J	�����VLjqdP@3j�A�x"qS�D	�Oq�͈�7�ۅ�bz~����D�G@8����
���C��aA���'��[�ӜOb{k�����d}�yE@:N����'RO$)B���~d�Ԣ��~�d���} �8�����r� jm����dGcT����R�����o_���9��ަ�}g��&����S��8��� ���K���GBJ��r��dC�������LM�u(c�zqȰ�+@���;v��@D�������	�<�3{�I�z ���M��j���Y�h.LB���T;�[jH�P���"s�j#�����ܑN$�M��