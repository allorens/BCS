BZh91AY&SY#�2��I߀`q���"� ����bF��          ��>�2�[m4-��D"�QV�J��@��H2(�)Eh
�wiKkmU�X�@��f�E��SJѳJPUP�p�*v74�їm��b��j�F���V����՚V���Gl��Z6e5���mBfe�l��(�CE�J�-�[d�+cUB�j�A�捩m�m�3�;��5Z�e�� �.̌l�I�7Z�ld$ikb��V��L�J�Z�Shڭ�Z[4LV�He�m��mjR���*�[e�)�0:���Y�6     ;��}�mܻuш)s��n�N��v�������̽��N�ִ�۪����꫌�v�m�k����vUm�7+�]��m����6k-#mlXj�  ͞{ �T�W�M=�M�P�4�GXt
�����/_q֚[�>�r�_9��W����\�z�J�w�� �*�cuz�s��hi�7��ZJ�2m�K*�-Dle��  ;�u���V��l�AF�oz_{ת Mx���F��������@����}}|�uK;�χU}������{|�} 
(��|�ϡR�}Ǣ�4l��C�vX�iV�  ��z�n��_q���h
����O}��O�����j}��/���B��UZ���}R�hh-���|_kz�)R����֕=O�������)O�}�O�Um�}>��U�b�[	[R�-����   X��}}���W��W�@
��}J^��w����(���}����@�O^�}4��|���������M>�.}7���X����g� w���˟�k-�V54�6d�0���(  ��C�bx0i@�Mw�ϳ��LP�=�J z���k�(w����sӪ/w:��^r4()o����P���q����p�U]=�ڈ�l�j�Q��m�o�  n`=m�!N�u�������^���mr� �Nh�k���� {�z 5��mƍP���
.zG�z얫3Q�+hƖ��%V�o�  רhӟF�h��{X� z7�@��p
7q���q�Ѡ.�p���� �^uց��Ҷԭ�-���fM��|  �5����_^t@3��� ��鮎����84=�{\Z�3�����g�x� ;�0:��Q�s\�QYQZ��-6l�m>  ׀��p� �N� �4�
(�Ӂ� 󕞀�s;@ ��W (;�������       S eJ��  �  �{M�)*��h�#&@4�M2bhE?&!)T� �@  j��	JR�3@M20�d���MUT4�@    (���&�4������2=MI���~?��K��~���u� �����֒�Vn���{��������� U�|�z�ß�@U��"��Er� ���A?�����j��@`��U�ި�
�X>��0�
��������o�a�c:���ΰk&�k&��L�&�k&�k�k:�1�ɬ�끌�ɬ:ΰL����ɬɬɬ�k2k�k�k&�k:�1�ɬ�����ɭ0k�ɬ��ɬƱ2k�k�k&�k�k:�:ɬɬ������0k&��ɬ�&�k��L:���������냌βk:ɬβk��L:ì�ɬ�ì�k�����������ɬ�ΰc�k������&���&�k�k�k��&6�c�k&��:ɬ��ɬ���:ɬ�ì�:ˬ�c 8�&�	�̂k :���Ȧ��� �� �
��&�)��k �ʦ�)��k(�ȸ���Ȧ���"k ��&����k��!�2)�
k ���k�Ȧ�������"c �������k ��&�	��k�(k ��&�	�(k �Ȧ����
���k ��&����ʆ�	��k"����k��&�	��k ������k(��&���"k ������"k(�ʆ��ʳ ����"�:�&������k"��&���
k(��&��&���L�k
�&�)��k*�&���(k
�2���k ������k(��&�	��
c(�������(��&����M��k"��.�#���(:ʦ������"�":����ʁ0�ʁ�
���
L*��� �Ȯ�(�¦��� �:�.����0�����*:ʎ�#��":��:⃌ ���� �:ʎ�#� ��
k 0����&0��c
����.��� �
��.��&��� � :��+��:�&0��0#���*����#� � � ��� ��Ȏ� k
�ʓ���*�"���� ����������� :����� ��.��*�#��ɬ����k&������8ΰ�.�k�k�k:�ì:ì:�ư��ì�ì�ì�ì:ɬ�3��.��&����&��&�k��&��&��&��ɬ�ɬ:ɬ�ɬ3k&����!���1�:ˬ�ìˬɌk&0�&��.�k��TN��&����:�ɬ:ì:ɬ�ɣ.������Ƴ12��k.���ˬ���k)2k&�k&�k�k�k�$����ɬ��Lk�k�k�k:ɬ�0k&�k&��ìɬ�L����ìɬɬ��2k�k&�k&����U���#�3����*��,/7[�o��>�ļŖ��/N���-ѷ[j�ŷo8^/��+e��-na�?�C�]�TH$হS�Me�`ӡpl��;{�q;�ʋ^' suee��H:�7*=h�4 m:� h[@k[�V�ZS�/G|�Bz����ӣ�"MC);NāV^\��m䢫$��W��C����� Ǡh;6�n9��û��q�I��ڂbj�2f�C5P��#Eܛ5��i�[�{vf��e��	��d2�I��j�4B�&�ٙ2²Ƽ�l ���wB�s]�2��,Ù�9Wt��A�o��P5�;�\�E�*�*F��v6�1�i8���%��g���yV���o��f����D�a�sol ��F}jIL��[�n�ʊ�b �Z�'yfhM�����+*���v
`f���P�qm�]Z/�4��<�MZ�r�4��NP��귒��bF�ٓhQN��c�uhku��<���6#��v��˫��Š�����)Y!�d�YLj��5�<��I�����I+I!�͕4�-�Va���8�4���Z��L�ko;,��{k��!hIe�v�Kf���q�Sv:��*:��-P-Ӭ� �#�Rii��;b�@r�lD�FH,��:u0�̨ʼ%æ	M�x�h }�l@r�aU�D��,�&�m &*�]�W�X��^T�Ié�֯u�mK:qý�[�^P�-��t�-�j�o�Zܼ�f\L�{[�	2���h���y���K�m��J1剅�/ :��$�� C�\�Gmp�6�����L'a4X�X�N&�,�q먨#����=gf?�.fZ�Q��[̔�{�Őo.�a��f��ԧ����!�V�c66�oh9�]M�Y�����Z+tPKNj�՗�Z�oL������<�ۻ6�)�~��x��YȠ&�U�'G���Z����N�Z���援5|r��*� �-��aZD�Z'-U�����I�4y<6���e�mm+ܬl�RJt+�BT8��tCw�Hc�Ku��ז���ǵ�+i�yE��]kj�X�*������e���uYL��1�m���C�'UVU���^Lɹ�W�L�*��lIna�:*�= �X�ѷ.�9D@E@Dx����M���`�)��Wz�ٷ�R}<��PC�f��
004��VV8����j�-�Ev��?5�)At�yx&Jݺ�'Nf����IU���V^D�:i�FFn� ��c��a�3l��X-��˃+XJ����� zm3�y��e��ov��X�U���'S{j�8̻���B���F]�(J�� Z�z�N%+0V;�٢�J�o-�9+/^�V1�0p���1�mZt�^�lv	
�+wzweAZ[*�ژ�D���]�i�-jHi�Q�n�$����Z��f�b��q���ӂ��s0��v�M�Ow.�j͈m��b�ߍ���StK�G)֍�9K��:�h�Y�6H$N���T�،7�lG��4�o��������L�;fZ���.��Fu���B-�("�Ҍ<ÓPH��Q�Wr�1��)��Q��D���.�L�r�p���i�������-�;e\�*l���%d�
��aն�6906Ϫah�kj81+�dŊ*�OjVˬ�;V��i�d�8�b�I�(=lHowW=��LՁ���I�01+�nG,�2P4�]��TĜöiW�ċ*5�g�� �-jD7VɳKhH�$�8�iɎ�4�$��b�i[�`�����F0�ꎊ�ӌ4M�ظ[�m�-_i�-�	hٙXoz�n�oX<C+z��/ZR+��0�o�&��f��N�x�Bu�^��$p]�W`�m��38�Xf�ͣI��|[���p�<��7/5�i�e�`��KMM"##�ósj�(k��q���R�d5���Y��d5�+���[��VA��X����r�R�w~�ƨ^�d�W� b�qT�,+���Q5J<	��G�����F�$��[�g�5J�.�aŷ�J�EB�6]*ra.�eÔ���2���u�x�ĭ57n	q`'��);}x�z,�B'l��n��������a	w��omR�ڽ�9�݅PÈJxKb���y��ʘklm��%\h"�5,�u1����	f�N���Q�̐�K�5�k�Cg>�W�9n�`�[�̟cT���'z��W�m��򽷵t72F�kZ1EA����55of��N�V@��֡�]��{��&n�yOU==g��u�9�8��\9�"g8��v뺖+	���0:;�/K�R��ʴcO�K3P˼���w>:�t���b�uj�Ó#�#hKB�F�������3iT]��*�ʙX�LE����[5�sD���2j�q�Xc���&�mZw�s{7*l���Y���s ܅;���Y�$�ܩ�1�A��0�7���ۡR�9+nGw��r�kRӬ���,���"����p�٥��+F��������n���z&#q�VR�6�̗z��{Oh4d�]�HKk�����u��жn�����ۧ��vH�w�iRY�� ���	%��R�^�yaY[	+A8�e��nO�����2#ûnL��$�(�aK��l��9qR�Vr���/���;Y���[vh�)`�=�V�o"#��l��ʳ�*=�fLN̤��P4�M�c0�

um%�r@�E0ۉS�x۰%Y�U��kwQ�&�5��n���e,t�/%����N7+.&:ٺl�-аh��o�oK�53N䱖H��!Zl*ƨ7�{h_�֕�Em�٧U*hH�ݲ���B���YF=7��:�C��$Ɯ����.�v�S`EKƭ�c��\�c\GM�n��Pkr�j������7����-�thӈ�rF0X�B[c��p�h�ˊ��XփGz���l˅°]n}u�������x�Ua���m�6^�E7�)�ބ��qL{kݼU��O"ܢ�@ֵ���sl*���6���P�v���Y�C
_�6TNG�Y�-w$�+"�ӥm*h�[{Gn�5j"E�1��T33~ؒ�"�yJd��U��+�u0���u��]Df��GZ�M8ef�j��=�)ڣ� �HM��0b�U�ȕc�c7(	�26n����O����Za�͡m���Uzd������ۑ}���I<���[��p�ff�,Mpm�-.;RO,S�����(J݁Ȏ�r��:��Y�kT���ia��-E��^���!��q\"X��ݰ�ZXtk��w�0����V�l��f4N��w��+ ��n��L��0]�����Y;����:���s]i̅LwL\w���ձV�aJ�+�ia-�a˧+OQ�v�r���u*B�;*�r����(Ө#{,Ŏd�l���PV���.b4I-�L���&��N���Y� ��jla�j٢'\�.�ur;([�&T2���S!3�9�<�wsU,��سT����9J�U��!�Mgkz�;��֊2��o)�UzQIvVl�f�L��jlT���n���x�I����e!�B��r����b�E]��DcI!'5%�	c�^%7�ӗ����;J�7]a=O2�v�Z�.�坍&�)�rQĳIeM�sq%�Vf�t�J�bu�"�%��ok5�ߵIm꧒��謷��Ǖ�sM24;�v�b"�gK���I��kH��W��g@ٸ�RL�XnS�:Y���H)��$�d�
:�b�	:��Ul�Onê�f
w�o��;(n�"z݋�WR`؝��������ݸ��4S��o,0�u���;F��I�V�p�D�����$S�L57\��F�F�i�m��T��s_+�Ȳ��i�.�Y���DB��.�̇X�@���hb���V/m���ܸ.��P�5���˳��S/{���dU�SEoR���L��*n�5W�w��5:\^�x�6,�n��$[Ŗ�:��b�I+�+2V�bWͯ����U,��˴��*�,q�]a�iOZV�ܗbQ���m�	�Yd��NՍ�KG_k�e�jT�v�`�rl���{U�>�0�c(-v� ٽ�]�j���x0ō���Wv�YwD/��2��9*�Uc��Q�7-ּaV��˻�ݴ ��cR��tֲn�\J��O׿4Q�lw�MF��l*m$ly#9B�Oo.e��E
���/"r@�z�<�]ؓ.����6Ȏ^�+�%bd%�pc+BuT�Ϯ^f�ϴ�/U��e:ךdM�.�Pdi9���2Ȅ�Y�w��vyt�,�:'�iႁv*m���o��f�̸6��Cdf,�z�ʐnm��Z��� s6�e�ǈM	05�&�'�F�6��E-��2��l�6� 6e:�8��Tu�/%䥡Y����kQV�]�0�f�B�nL����ͺ��(�z)Ǹ+�%��M��l�f����ۼ�zp�d&-|Û��Գʙ�U���ڭP�K/2L�!��uU�l�� ��vR�W�8���^�ksĉ,T�r�(L��t`��$�n���L�[��)KPݷ�3P˳PP;�W��T�Cé,��d��%�.��˫ȝ��r���2%F������-&����yõ4i-ںGFq�T�3LfdK�^	��%"�{t2�z�4�����8!8`F]�ס
�%e7	cmfn\��rORg,��f����-���-�6QVd��1m�J;;�����h��w�3Y:NX{r���X�7Xظ�.����̭ �!���i�wN!};��Jp=+(����w+0J��Ωiւr�M���Aػ��`juH�h�!�R��k�*F�V3�1H��Ck��m�t�͙�R�f��!��u[����"���|N�&N0-��Q7V%��lH�f�7�j���8�� ��U`�c����ڑJ	+����ţ�Z���$�̷m�լJj��V�n���N
�L��=�V4�4ؼ��FV�F��s)��1G+��aŊL&��	A�9��koO3��o��C�Sĩ��j!V�7����@��{5;]��&�r����]e0�t0�{F^I�&��2ӲCYzp�{M�Ϯ[F�hI�p9�ʙ0a�5-��a�[b����͚K���Ly�QwL�']2��xI��Sf��x�ز]�l�:̨��K��r:��`�/s^act��iI�2�B��znY�P5GB�gO�Rҕ�&��D����,�Ѵ���Am6�^V6���v�8��(�-���rZMYw(V�� n<C6�-]mWShn�����KB�[Vp�Q��VGpL�,a�ǂ��opBdH6�cq��F�z#��M�O~Ѹ5,vu#]�[��P����wtq=ޥmM���/7ab�K#*FtV���5B�����æI*0y���`����N#�sr3���� c�p�����X�6F�W�n���jjc#�·f�a\.7T��5gdb�m-�d��+ky������Z��`c��{z���*|�Tz�l,�Q��^	t+pE4C��:v�C.��^��%��%#��cd�a�&ļ�\�%��n��LfTje��9w $�TlL��v��H60�ԸSܖ�) A)�3EZ����X����q˻{�ZѴn�S�H���$&�J���[�[��;�N���¥�ƗGeU��u!ۨJ��np�$:��Ӂ �ϱ<�//{��ҕd5�V�2;�a��-C���1�:�Y���U*���na:p�yH�#,n-�)Ӷ&n<�̒$��*͛�Ƭ�䷷,H�Χ���PP9��r609�R��$�fRI�h5ǵ)�@�Ei4�O0�Q��X�C#�d��7D��G�.��:�7&f]|�3��(��6��ݑ���6�g��j}3�z
e+e,YZ��Ć���(]R�q� T́���E,�E�f�c/��ܣEY�V���,̲%7ebkv�#m(��j,�Zܰ�nrZ۶t�ԬɂD�՛��pJ���Z��j�5 ���tNs8	�e+�m�X��#ԩ
'v�dj�zv�[݋.Qݒ��&�1LxrL�E3��X��C�ǉԕN]�	���d>��*��[6��=,�����(������$Y�x<DM櫡�4�E�%:D��]xG�g� =�/j^g�'H�g�V��4P  E�<>�b�F˩d��i�}��Z�6 rB�;�]bBȳzy�%��dAl��ei���Z�ۉ���|Ɯ�P��������͵#�kD��ͷ��ZNWU��K��|�m�xukdrKR"�L�����W�kv֠�	�]�m�V�f��T����I����U+Md�/� �/�M���� �$T�κ�=���6N �\�#�^L��T�1�P�h�����w��6j���T�z*QL|54u�1]L�X�N��L�)$bl)Z�E�i*���.*�%ԥ�m���{�pK�Ccv�c��9��@Z7��,o(��ђ^�%��fAkK��Z,&�Й�1+m$" ��1��&��n���9WQ#'>f�l������hQ�`L����t�	2�`� ��HS��b��|�D������\���M-'��C��%Y�Ih7�Ŕ=�x�/��ߎ�lr�
���.G>�~�`���`@�m�D���	6K����H��@`<�����U��V���ȓQ�K(XmEp�$Tp���b �(�1�မ醨p�$R���3�Pm�^6M�`���l�&�P�k�Ϭ�'�P�R�>����"��m��b���~���j�e��Nj���7gȜ3���*^�{�3��pUc�l���$Xj (�۴q����!�m��a;؇><�cV錺���e>���!N��i�d�&��)�ItS< �|e�E���� �dgb�xG����uqg�Ԅ����}�B��E�������ϳ�����]�'Ӟ~O��~�t�Z����+��2A�H�L��w3�m<���4�=ά1�C��KXh�i�uyJ��2,�Y#��>���&e�몣�Ȁw�*m$��u^�K�]�n�_7W��q��S%_W:%��4٭�Vm�9�ҚG����6�2��1gQ}��<�q����7g6�i.[�J(�� ~�g�sJ�-�8l�W~�[�s,��ɰ���.ѓpL�F��<�E6SJ1�Yu۬�|�]r��	�KWj�eV.�Њ͎�Gc��; �ŋ�fN8j�wt��D��^n��%U��P���I�4�*ޟ��]�3�1WeY�{��e��C+�n�I�m�1^dy���KT�X���ӑ��Xc�N�X�fYU��8�#�3z�a�mFNfgC$��؃��pE�b�W���^+|{�M�m,Lv�'A�ikB��,�� �C�<e���UM=6�X��mb� SQ�[��^	c�NKk�\qk�:�卥�ln%��]��b��.w>O7b;��.�89H,�-)oGR��q�w]��s����N7{g�8��AܭYled˅��4����](�I:M�L���N9��Wu�5mpu���n��2�YWG�Л&�(/.���X�:��ʝ�ެM��˫LY��wt��5����/0�����Hwo�V���U�ǖ�-��E��B�:uZ���:���5���z�^N+�T�EMԞ`��3���a�;�q�W!n�%��5���6�躹0c�c��{wu���G�̖�l�F��3.��c��WP�6�[yP�-Ý۷�"k�z��X��WF�E,�s�;��,I�����eθ]��S��E�����PmH��.��A\��f.�G�(��Y5��j?s���lR�5jSx�]c�j)A>݄��j��n����諭����aa[�m��^>���S����w��΁��n4���y.�x�ɧ�uV�j�%�޷J�v��U0��y�qz�i��NML�\��7��#{9�(lՙ���""[pS�Mi'*g SC:�4[ҹ��%��;��q�噭�u+(�Q:�$ ;�ˉ���w����'=$]���3Cs�gZ�6{��]�pw��{�������{��rɸn4D`Q.i���#3�\��U��f��Vx�W�0b��Kۗ�77-�L����)�"��}���pnX�̫�F;ǧ2���B��ӭ3:�<�+��9���;�(��g��r�:p��u+{�4��������v���x���Ӧ��s�'(���3�辷�xtҩ�ӧ�/�_|�dE�-���<��aaܩ�^V_\�ېܵ%�y����i̩SUms���C@'*��Kl�tBpAc+4�-��۸.W.�x�|`���94JP+G*^%��3u���8a�[ײJ�L�od�>��p	S��Y��[G'#w�	չ}	��x�z�N�E�m�g^mFX�0�W(JO(���>X*l7�K�<���I��[{��k%�x�i��09�ӂtwj��' �)�r]B��չ�Ά����C*�]��]�oG[�%fT|iEZ��Nˁk�h�hݛ%��{��*�*'o��
��/>z2t�Tw@�b::���2tm\�^�_���5Q�(Ԫ��$�w��ؖƭh�m]�=a6	!�6i���,�󘲺��cJ'*������o;: �gT��"�T<��[�0d�hlpj�g��h���5�^��	و"Z�ԇ[t��\�"	-�ΰ�3�@E�KJv�tm���aᶄ�մ��w˹A�&�T��w��yZ*��+�ϝ�`�7����G��4fS���M��/̾�%������$�s�:��F�7�21�u�����B���{����=,C֯p3��)wpN�^U�1.c���E�\<��[��V���^�����j�r剄���h��)x�R�4ر�Q˭���j���ܹ��M��2�X���`��m�虆T��Wv���$�g��##8S��r2�X�o
�tX�}2��M�(����i�W1w��ah�+5
����.�ѐ�	h�r���x*l��F�� ��
b'�ʥ�!F�������E{\-ܩ���n��L!Bؤ���J'�%�%�_g;��Z�`kt�j��v����y�Yeҽ\�Z��S�\�.�k�|���d�'uv��5��֜	�s�W*t�Yu��W1E�E�*m�N�#�;
KC7n���f��B��;5C��WGc�����}���w�C-�.��yd��T�\ ���𱐑�����C::��a��a�;�� �t�7�b)ϐY��ibg;:� :�ݺ�]O;{)S��@���<�Э�<�3��ٜ	�z����T��Gi�;j��%�mS�5]�j��9:��-i�o�t|���nV��1��&`�
��i^s��3�5��3`�ti����փj�8n� ����{%��O}t�*�o5Ac����C��U���.iC>�q26U&���wD_A�@y�@�,ړ����N>W�r��$[��8!b�^���LCnT	nm	���}���7Ҋu�jm�\���(��Ab0�l����r��p<�ŀ�7r�Mr����G�֜�i!yWO�Vʵ���
�u �b��L��fJ�m=y���];�#���c�#�,�����T�3�h��7r�\ѽ��ss!��9��g��v�|Ӛjdmڥg]y����
�)
VG'�Hi<��N�����F8��Q���I���4OVD*pn�ŀ;�1Z�+"�R��/��vE/-Lf�2�n���w�rzƩ)�����֓�P%��ǶV	��p�8����s.��R{������/Y�Ќ��.n��{��Vڂ�aa�Yr�q;��5��uSK`�vuS+Y�|L�`tJ6[(�퍅�-8��n�ܰ�gv)�HS9��<���V�Bݹp�2�v;�ފ gA6��o@�]�¤�n�8]MSr�W3�J���b�+s����_9�4*���r��ּ7���ͱ�}�ݙV�������7i�ꂸ�ywW�x����)�6��ñ보5o69�I9[��\ }|UXU�OM�wy��N�P����aʕ�*:�4R���/��+�ln��;�R���y:ʚ��ˉ�$ػ�B���k,M��=+n�.��
óU�kx��iU�������9�g���`ɴ�K��Eu����M��|�l�ofTܥEfIp�Yv9���`E��l�Dۆi�F�NW	�߅;컽��՚
1p�*�	e��F���;ՇXw133����|Ou�4b�V��]^��,�m]p]�M�Ib=`��W��w:*��`8MfR���m�Ȉ���j�Xm������^5�w�6Ù�&0n�j﯑���7t�Pu�*&��<.h��+yCw��Q<uT��:S-l�iqɽ�@�`t>}�V�l�&�ċ�̓�t)��oM�R"z[U��_h�S���) "�B���0�ޡ�����f��^�md\E�����䳬ea�D�hNklEs��d���B>i/JV3Wu]դ�[�34!5Q��&ݙ�dj�E�HA��m�̔e��i^fF��]����3�����_1rJ����nv#�o�Ʈ�����^���(,�����b]�9ǂ�
U�v���-��N��m����\�zCYh8��4h�'�Ǯ�0jlf��36��.ZmLB�Qf�ͼn��r��PSb�o9����^�_�U���>|�B�;���l<�-Pɕ6���ʺd��f-ۇ��w�,�|�5�܆>�`�};��wH#�Uf�	\a��7�����k�،�����֟-�ܗ��G�L���ک���;��2�֫t���K	�D9�
dj���c�o�v���Jj�{�HlY]�G�0+V���D�U�XU�e�f�f�+8d	�V ��E����`��S��j��y���y&�-���	�	$r��
��y�:r�.�O�W��Х�a4�(�gR���[ю�`�\XFb�!��;�^ ��O�����/n52lH��2֊|���ef%�n>6�f�z�C\(��5��r�[��R��1��J&�X�p/��a����#,�v���ጌ�B^��s)X�R�EfL7XCQ�|	�[��q�.F�f�͙YIl��uZ�uX��o
��]�le��T�@��|��� ��D���w%�Q�V v%�R�@`8m�ݷ���fj�gMJZ�����!�\w�O�1�÷�{X�TnՀ�����cs�<�	���`��>����p�k��>����@k����h��^�)��i"%gH�)��/��W6]m
i��U�\�<�;�7��x��;�b�+���.��5�VXӰ�Щ�m)�җv�Q����sﺌ��ө��4Ε,f�������b�o�=/*ͱD�����x�G1�v���)h�|B��g����/���`PW��V�\�ZZ߶�5&>¨�,�۷� Z��6���C+��h�U1uB�RNT]�y3�p%.��e�5��n��am����ip9�p-�>�	a�p�V��εn�Č��$�!ԋz��!�<�]Es^ȶV�s:�Ք&fa҆�-�;�i[}P�ǳC\���+(��5��^+f�����h\!����Ƃ�zp�m1@X����Yu�Uby��Igr2����֧Wc����vl�gV�Q�Xd������.�e�&��8�"���G�����o�3�(�D�z5:�}8MuBE�	�u�צ͟���܉�(��9鶃�T���^�Y�uʉ.�,�gjz%�b�֯��wBp���0���\M��£��n4�(�����ej�o�W�'��)�=o8�cw�MԦ��{�͊ł6�]ا9n⛶����7%;[���X2%kW}��4,�T���� �<�B�
h�Q�cU� �2A�:P>�Fd�-�E:v���qn����RW�j��MN�N�A�+���O@����z�U2� j϶]m=�������3Yʵ�96k��71j�e��n�Pl�t<(C�f�1N��J��ڻ�؎��K���2�,ԝ)n*Z�\�d���a�R���e���F����Z/���qd&�]�`�}m��e�HWT�%�}��_J��4�1�# ����eҗ��u3T��1����J�o��@>W�vFX9]��hǕӭ_fzӔ`'�+��W�g2t��Y�L#Df��w.R5*���b�H}�l1սY�m9^Q'l�H@��V�i�/�b��n����^��L�B㠷�b�p|8����3g:u)Ք�Sqy��D4���۱�&�nR2
Z5�N�'Po������wڅܣP�;���b��h��>��o��K�7�t!�gt[Ó�}M=v;F.�`���p3r��T��M�8?�iv�����^�֌��.�kCNZ�����Up�J�V�Y/=�"�>&���Hޗ\j�`6_)^Av�ڨc��͈��n�ʛ��Y�{�	��`$�9��@�Ou�����Svg=
s���T>��̶h��k���.W�����%���:��h^�|�J�˧rM`�^}�8��!%"tf�p˧l9����M�]������HT�;Z�\�s��ʶ�Nh�2�aj�*٪�/mP1{������U�5�
�j�P����'�����>���^?;�#�,��BR��f��Q�u�D����8hfTt�LF-=�3��[�I�����l�����v��Kj�l	�Y��ʷ&lz)��.)��u����ĝ
��MJ����HK[3�Զ�^��1��T��r ��|6�돎B��J�y�Wř�ӏ'q%�gm�+X⤱��݅s���n�7.F���3��.>�l1/m�<Z>Gk��PS%�2^�C��R���(�0�ƥ�v���\�ZmB�-e�4��V���� }���bƫoP���ƛKq�ڱ�����N�ˬ{W���C&�ξ�3fX�RC��}�v�' ��gs�HP.!*GQ�ʼ������H���aY�@�4+���x��i�2��R�+�M
����u̵Sc,ܭ
�nl����`��������� h�W*Ӗ3#W��g#������`�{k�Ҵ$��<�M.u)�W_^h���\>|s꧃�@���OXa��}z��]���]��H���3�=�ߙ�y����3�^��#�H-L�?\C�Ԭӏ�z����Ϟ���o~jmK�v�1h�g�G7uvL��$;e����tK1=o�|O��|ۚ����.H{����=��~�|�O��~�$9	�Td=�l>�����.I����`�~g!L�����$�����2���]����S��Ġ>�>���P�~q��]�����7�!jqY��@��g�:��@#��pB>�~��X�_�x�G��������ӹ����y�s���|��vr���9���n�If/.N��{�=A��@AG�?i�w�� E��:�?z��� ������Ǟ~������s�g�k��G��&�d�;EJMaz1�xv��a��NeҺ�F�yZ5�d�����s&}��U�:��E�mg�1\�ǲ�_ �iU��Í��e��_G��AIB�[�u����a�S��'�ѵk�m�=�ċ�}�]��7j_��O��d�أ钝��TB�0_l�7�U���!��<��z�2�c2/� �Z��R[�Q�}	��q�cL�S;�)�֬�V��n�C}�[ ��S��[ͣ�R�7�]�T�����Oc�^�v�e�y�	�1���ێ��ѥ�БHB���Bޫ��[tS�ۚ�O����3�m6� �ˤ�r���&7��#��[j��)j���	|�I3a4�Hmrm��LQ�
j\6+�ȴԥ�6�l:ӵV�C풭�R�h���C�ײ��J�o��Y��p�=�w��[�.@�/����3��e�wzt^k<��#�G&��}zF���-B�rc ���l܆l^;��aY��m5[O/
��$�ܬ��t���U��tv�Xi2�ּ�f��6oq���(PI;S�]n�}�ZΜ��}(��r�.l�4Y�Dm�p�t�:�ƒr�t=���;'P���#(�Xԍ]�鋍@��5�H=��MI�(`����ˑ�w�񠫶|v�ͽ��x�Jc	�u��~>�o����ׯ����]z��ׯ_o^�ׯ^�z������ׯ^�z����ׯ^�z����=�z�z��^�z����ׯ^=z��׏^�z����׮�z��ׯ��Y�ׯ^�z���z��^�z������3�^�z��ׯ^���z�ׯ^�z�����z�����~�\~�_�ׯ_O^�z���z��ׯ^�^��O��ǯ_���ׯ^�}�z��_/���=�}{�Ef�`�0XLZ��듛�A�w)�[O��OU��Q��)S�������7�%�J
��ǲ�@ ]T{4a;C}�txU֮�ԓH�N^��$��Y���K3g1vT6���Ly��dT����S�c�$����|a��]��^�C�	��w[62QcX�I�̙ ��Ds:B�u��W���<�U�2�C��BS[@�����:Ab�N��sQ������P&.ˎvY}�3�A�	����г�J�3�p[�V{�T�هh�]ۆ�55���� ����[�M��9iL��Ù�-��]��}�x�J�Wu;�F�]GD��ʩ���[��t;�Wq��bn�`Cv�Byٙ�%a��f�C|���B;ՙͬ�X�6�9ͼ�[�/����:j(+��hwX�(�"O��x�6���p!���:nr9��%]W��mܰ���*_A��jb�FK�U��S١]�̨z�{0Π�Α㧜��]7%+�lw`<*]9v��͓ٸ`M�]�bZ��.�e��u�SX���xw����n\�Z��"Nۚ��>;�VYY���ȃ�k/hǊ��8��z0,6�5y\���;S=��N��n�q�N�Ђ�fr�U�ڤ�҆�]A�	�ƫO>�{_�q���eV}>_?��ߏ��׮=z��ׯ_o^�u�ׯ^�z��ׯ��^�u�ׯǯ\}�z�ǯ^�z������ׯ^�z=z��ׯ^�~�g�^�z����׮=z��ׯ��^�x��ׯ^=z��ׯ�z��ׯ�z���z=z��ׯ^��q�ׯ]z��ׯ_o\z�ׯ^�_����������ׯ_�^���ׯ^=z�������}<}�޳��}>�O������>ύm�	�w݌���@tٱXf�X�8�(uh�]�B��P�8��fR�v�TR^��s�{���k �����ыU��PV�P")G�:1��T��t^��C.�Z)��GIT��,�:G�+e���XnM願&�6���~���LtUm�Q����C-f��k��<[����no�i�:!nVST�H�[�h-%d��
Tnn\�[5��3	�뜜��ד���Y;hs��P����|e�]����x��rHv}e��u���Y�7�WM�p_ԩ'E�V�(W_̺�ڹ]�uI��e��sB3]��VFsZ6����������E�����=�k�]��'�x��Q��u��F�e#}�*��6�eP��_}J��vKF#�`4,�����[4:����E,�.�	d�N	c,�1q�1H�7���b%��5-�����g�Wt�gu��|Y���s�T��c��u�jSM7%��}3#8�����ui�f��X/w#v����.�un�ٝ�d脤�?�W�����,�p����Z�5��hZ���`�]r�옞7S+�����.�
�x��+��ͩd%�89����H�;+ �X�\(3J��+6��#��ou%��Y��0q�͔qZG��pQ��xOum+i��pi���g���q������z�z=z��ׯ^�~�g�^�z����׮=z��ׯ_o^�u�ׯ^�}=z��ǣ�^�z����׮=z��ׯ_�^�ׯ^�z������ׯ^�ׯ^��z�z����׮��z��ׯ_�^�=z�ǯ^�z������ׯ^�}�z�ׯ^�u������~�_��_�^�z���z��ׯ_L����Ǐ������ׯ^���ׯ^����O^��f�,� ��� ��E:�Ran�=�i=�Y#�,���<�L�팎+2�W}���.5��q�#-�(^V�-ls%��u龓'l[�i�WBV���*��Ʌ^՝yb��M��|u���}�P���5�������@o:�*�o��k ����6��ʧo��S��um��w�@su�{���۫���W����zeh��
�9`�0t�a�b�m�Av�'V��
��q�uM���$���4+=22i���_n�y���ƾ31�����Zb�*Q��ø~�teՍ���Ϙݼf�Wx/�J���9�,Nq��L��#��u��e$X�$|.��b4��Т!�ꂹ.Ⱥw}��[δQ�=�[3#�|��7@�N���S͵ɪ���e@�#eJ4^�Է��_|1@��q�x�&7��_7o������|�L}RH٧���t����� <Zm����j�i����5;����ﻌ�� ����;��]/+��(n���1&��һl%#/v�,� �4��X���Y���]����[{0��Q���Wpմ{�҃�H�Dw"eZ�I����#Y���kjq���JV��%��{싲}r���+ u�L|>��%�2K�Ԙ�7��:�c����^22�8�3�l��;�N:R�+�.��Q���}���C��B�u��D�UH��zyi5W#Ì���t����^���<)��i���)��+w�
�:�|v�A��4(�y���;"�����[�L��f�k+� ,1i�pz����繏��Ifar���f6�LMTj�����}7o�/�)�+ݗ��O�y�]�� f�[W� �sPE;$�H%s��y2;�"�%��(؎�q}�e��2���T�Ο+�Eܔ�i�X�<P��2��x���EQ8�=2���'�BIw1�,5G��\�F�+���VMò��bol�����]�G�L٭��4bw��!���xM$mH�U ��|�mf�>LD�I��,u�i�bJ��Z�'�A�J@�p�('��#�6���C��վ�ydU��.��g�	�}1���:��$W>�J��m- e��f'� v���UP���aZ�ʧں�i0��w��>�q�
��ȡ@IA�����n:�5�v��vK:�Q_l��a?>�t3��	�%����Zb(���b��@c���������9�ڥV���}�G�$�;��"t�C3 5,
�FR�{��X�n[*��}\��F�B[̔n����V�b�s�`4k�Cm�)[�2�һ�M���e�}���;�U��S~Ͱ�w'�y�5�JI@2s�\&e���`��U6'Y�a����G�%�������<��k&C��SB6�I^�&
�<0�s��fMi�ېc
�����Իx1� �G��喇zGo����*�Dz���+B��UoA]>�7�/�nڧq�P�Hh��i�<������;j�n�׌sw70Sԓ%�G���!�:=��_.T��#���b�˅�r��wJ�����x/�4��0���>e�3��U4��{��`��G�RZQ2���
t�r�V�ٰT	����.�(��B�w*Z��ח�mt�[���y����
	tcu��fWMA�u�֜j�0r�>iGօ?�@��'���{((K�d���٬�{�i�r�TX_sL��Ԫ'1fZ.ַF�����{�����Z޽-��2��f�}7C�,p+�F�gb���_&$��Q�� Ķo։�b���2Y�H|�����N|x��v�O�E�͓O�ٔ�a��3�����9�G�Q2�5�4��YZ�/������+P�N��I)����}��k�H��!l��c_���f�N[�������X"Qsu�(e�+�۹ٸ؅�p��Z�s���XӶt��Dݗzq����6uK0�|A��1<n�`�a�q>g�7��R���i��tjg���q!�:a|�Q�Ӝ��ڒoT��|��$�ϓI�Gf7��>YI6����㝲�F�����-�ȘpS��X���
=��XdX�>�p��v��̧�\*8�cF�J�+'`C-cȒ)���c$�}0֩��_��x
�mf��Ï�@�_V<-��VV^� �״hfĐ��C�a���[���S{7�X�],�FЄ��� �K,�A[	okG{/i�Vйtv�8jj(��׭t�ܞ�u�L�;Gd����y@�����3w*���E�9��V�鴃�MLL���gjR-<_bN836U��mf�O\T���s>�u�Yd�C��w������r4ӝ�����c��v�MV��{�����hf��Y�-�4������oh]�=��-��E��PH�h�0�m��
���h㋪7e7N�2E�<�p�u�D&v=��4F�e�KJx�8����G���M�]b�=��p]@*������*�X�.�RM��U�]�������#L�t�A7o�"�1��Τ���m��յ�#:닷�Cw�Dw���Z#�}���U>��e�3t�uRɳ�SE��;��@�d��=URjC�%[tfuJ
� W�;�8�ܫ�3��gD�!��$��uQ>�9������$Fh�:4�v���9�dW��^��lm���ӎ��K9]����=2F́�Pf0g'Y�>x/�o���ZJ� �n9Ta]G3L���5��v�-Ӯ�E�D�ξf�l� ��9L��gH�M�����骮��롭�~,�y�!g�U��Jء"}�e�;��z��k�QV��m���4�{��Hm�7$�3����,�X:�ۅ$�̖f�A��k�jVr�s�sgSa�����t �>ʇ��Yƅ;ᆵ���w3��`�3~��B�����i�N��Jz�n�#g)�8鬣���h$Q�Uy%�^.�[36�B�TP9�jجU�ug!:'l�����\[ֺ��9G���cF��<��lq��H��W��l.��i���%�r�C[�8b85/�ӯ,��b�K���9�W����݃J�Zq�p{}�-;l|}���6,9.I/��(�E�2����N4����̡�)�a4�.�1�Y�hNĮŉe�s+]^���A�S,-�*>tZK/�'N�ʹ�-7�u]�FV��Ŏ �&*�1��x̘we�t������@���)G|;�̀�%�t,R.t�;QD�J�g��].��L+�0�k�0�*���]�2(�n0v�Gs멅Ӣ�>���{6u1V��M��]g|�kAF�J�u^W��㆟f=�^�7Hܑ�0��v�ᝧ]:��v�UYX����61b�qɼ�q8,��5N�M�Cx��]�G10�Vj�nt�Py��0m��#(�u��e�H��3_�!�+�{�!L3S	̇�r'�e�XY�WEW�󭥜��74��r�e�2)�{%�8fS�%ա�"�==����pC/�`-��ѱ6*�b��50�f�w7/.9w��n��E�n+YR%lr�1R�y��L�a,Ƭs�]�t������L�S�gk��7�2�!�*�%,˃Q�)�i��*�bCh�l��5�+�m������6`Z�0�P��d{}w��EJԎ82�l������Ar�穷���7g	ج�IB2Z�����~=��S�*p!0�1FԆ��j����ܬ�=d����cU�]ɩeʺK��{�9�|(����T�l�ڈ�(�	D).�KAR��mJz�tXLoJ�r�P��c��O�����(]�H�K�����m����!���-|�b@�#p���U��-���'Z��1.�����w.�6MI�v��{g�����f���㐑��¦�;,F��p�(V_hӔ��_�2��2�����5^ե1�l�Յ�S��>�Fv.�޸NmI}�D�X��4e!�]��ǩ��8�k�$�K:e7��Q�G��i�v7�)����i�M�:��p{�h�͋~�{�R��Zo�s��*��C�1�W����()H�]$�ᕳi�M����7W/<����ٸr���e�3��ԄI4�-r�N����%iY�j6��8�y�LW���*���#l�r���7&NsVh�PĆ[�f��Q�b������/����o^|gw-g��/�_E6����*W3�[0���k��tP�ڹ��M�N����픲��v� ĳf�V���vS�Vu�'��"���r*^3����yQܔs
j>*������
�˔�a�1>Hg}��k���:
��h���$�Z�2����Nu<��T�ۋ���2-}6�6%4�9��`nЫۓR�Δ��p�8lv�'Xe�!;���\or�s{��s�l��� ���N��nP�suͽ�X\��p,����Cd5�g`� �s�K�4WR���G�����;���z]�%��.nm�����uަ��p� Dԍ�3w7'fB��1	�N;jR����79R����Y�)jn���������ls�N��m�%$��[��km��Ȩ8��%L�ΰ�G��}�XRh:4�N�{L�����R��-ˀU�u��HF���.��图�nw���s�~t�������J������_�����/������?i���.fi��7oԪ@O�4DAH"1&��$Xi0�m&�rB!��K��2�4Î
&�"�e���N��H��i�"L�A_''�'�ƃ"4�e��n �%&�b�!�#���C!1J4�N!L/����A>�K(�d�� �LP�IE	���Z����XH('�(-2jI�RF��7!aL)� !�	0�i�\A��b�_'�3��O»Zъ��k�!��=��K�s7[IWCr�+,L6Oh� Z����ܗҜ�����k$�\.ʤ��4��K�ސ1�����c9Y�(޽4�y�����Ձջj�ݽ%3v�@1Ik[s��O#/��8)ʄ#��uoP�sʽ	=��}u˕�j&��6�m���:�J�m����]�̶���YG�^,��:Ĭ�km���]���;�_\"�̗��)�b�t��U�t����{Yg;o!�a�ΥX����QQ�4$1YT�GIB9��Ԓ�N��^f��/z]mF�J%�kwrb4�i�5�Ľ��$�͔�l]}ԑd�'��P���{�Œ�i�u_j7����թ���X3>|]_a����T�o�U�����b�^DX4E�(���i�t�Gnd�	d������8kbg8. � 7[[\�&k�SΈǹ=���g���jT:	x���[ˁ��$�k���"Wt��n��2l<g)%[�P,ٜ֍mY���Ï�ɚz����z�i� 8齧���
B�^>���tN�>�H$��\��g�V����J1����}�C�=7P[��gY�pn)x�}�x�T���Z$�O���*R��h4��a%0P�@ԑ�
6�)�����4�1~d�H D�d��Rt��I�E��H�T-�a�]|hDb*B�i�`�I$��i�e1N$#���e��P�"%S!�l���\(I.D���	!��A�H_F�pB�P����N$D��-��DI6Ij4��F�L8SBIO�$0��Ȕ �1��LH�i����hH*J�,QM���،5 ��DF�nd����IH�*0L �>E&�JA��N$�2,��mc%6X�H�(jQ�����rK��2�r�0��i��re@Ъ1~d��cq!!)����"? 1�>FLi��eO�?2�aDQ���$�#���n&�r#���B�?2�;�A��U%A�Qg�vs���;���u��׏<x�z�׬Ώ���2�BQ@S�dQFC�QT4�ұ4QN��hκ��Ǐ<z?�fp~���)ZO���v;�70� ��X@r�l�)ʃ��AHShc8�ׯ��>>����3��{�kc$���J¬��'s+�4,3w�ͫd0� '3!"i0[0��l"F�1����2T̳
���I�y���,fd�A<�G&�f$W2���7p�(b�vlȆ�C
#c�;A��UR�͍��#��l�aQ2�0HV�l�Y�p��30��br�3p�!�̐�)�ʶΉlz�1��Adb[�nd���9a�f�ZE��L���ȧ/�m�㸘Qn�dz���"�冱��x�����\M�L�ʈ���d��p+h�1������sc,����+,ۑ�,�,���M.e�û��P��ː����C"�}����噺����A%IM���ѹ���h��ȹ�9aE�����NLA�q��02�&G,�3"�9��!��i<�	)6����E��%2M�' 9�0�nPl��2>�� w�>e��F(���a�l�`�>��̆$�	���*	��*��S"{��>��_q6z��S���|6��ǝ���w�7��1u�;<wM4d	E
�����)�,@�26Iq�L���d�\_4�M@�D�����iA��g��L�n3r�\9r���<4��3b��Ý���*�@��L��M��b�,�ߝ ��Ek��"�f���n�����T��ͭݛ�n' �&��*`L��W������?��=��)�M������yUy�-{�ۮ�x{�7[^���W��S߷ޏ�}=��R�7vonD���/y8q =���7ݕVw(zo����L�&P�r�=�n���q�0���]�DΛ���^�1T����q{UN�xVY�t6=F�>�7��:�O��O�<)��[��2q���Ӎq��F�י�Hk}/} �x\a�ߪ��Ϝڸ|���wW�����)��@���/uL��\����o���`����y���/I��-��<�+�:�x��^-w�:}�Vd��s�`2+��S֕S��|g����W��0=1�^��X����RǍ�oO��O���y��c=���4�!N�h��_��sզ�=����3��р<q٫�Qd��ϭ+}Y�f�tQ*ßy7F�#=��Z���µ=t�1^�8O����m�2��=�;��a0�;�͵v..�<o���:Is��n.�	��4l���5�.�ĥ��yrg�Uk���1�[fߪ|�N]/AOd���(.ϯy���{-�u�X��D��4!���������H!u�꬯$z��R���נ�I����_����=�j�L���6t�P�q���9�c�6j��=���>�<�:�g$'�*���~r��Ol����e��u�����񿾯�)�z{��_>V�����M�e{;կ�������>uy�ݡ���Z\����/���3�"��KE_�8���r�<�b���0U�{��!֜@"�YIxt5�v��T��N9�5S�G��GnI�(A�k<��޻�5��_Ssh�� |x�Ǧxo���SvAw��ݢt��t��s�,ɺ��2A7u@q��M^5�ɍ��{S��O�W�������WQ���}�~^<�܍G-��>e1�w�=B�����-��ӻ��g2���q� �abbw����!Щ�vm���Kݽ��J� oNbc�\ݳ��XT�ވ\��Y�wC�m�[��.}��WX�1t��Dd�m���x[��)��0L�/V��;� �=��D��2�Sd�����EX\ٹ���o}]��x����M�s/ǉ5���4�a���9�FrA�x��l��7�E�\6�zn���$�����$r�q�]q���>�b�K�JS�~��l��ޯ�	��]��&�9�Z,�GI���1��3��z
��x��YA}r�8�V��.[����*k�%�3jP:TP�#<+����;���a�K�p�����|���os;ӟ^i.e�����k�U�S����]}>��i;�X~wBD�L�>�mz�=�&��Vt̯�ގ��Ua�je����>�K�Μg�U��p���9�@޸����0�4��l^���e{��WS���ǝ�׎I؃�s|�oɀ�u��cj�����}ᖼ���w&�b��fߚ:u����Ӝ$Ѿiஔ＝�Z�qs��W8{�vŴ]tʹ��}�NlZݣ8�P�tvTŶ�|3��`�/0_N��9��:t����H7�n��wڱ\ �:�)�[�(i�����Q�����q�]��RE�J�W�]����-D��<�9Z��P66B�]�Ơ����@|*�W<x��㕣�^�\�5����}ن\����/��5��|��U4������G���2Mx�������ǆ�c�BJ�b���x�S�[ծ���Y�`v|��GnS���o��p��<���1��{���zߪ��13��[��/$���BMߺ��e��$�7��@��F�v�5����EǷ[�a���37ҩQ�:�Z�.�
� �@|�׶�g���W�<���c�u]�[��mb�5��S�|3ٽ K=�w�L�X���mcp�3��SS��g����c��0����ȝk%���}���&��9תv��{�{�����9}y~D�Lj��>�W�i*�nwo?U
�ɥ��JV*����]{�+�����PU���
M�9�߻�ߑ~�;��3/�v)�%=>_U�6+��=�)��S���n�T����_'a��m�f��8��#�E1y��v�A)�rv�[�T�>��O]�]�I68/f�.k�|t\�o�2�3�­���z��ï���S���oNMH^��̒ec��a�z��y(*�߹UN�����$!�w�+����n}l��*�*�ɫ�O�\�?fg*.er�W�|�z���ߺ൝2w�ZΛNfT�9�f{c��i���P��G�^�~������FUb�j���R���y���9J{�_H��Ns�M�Am�>ޡw�����=�,�F�z������Ʉx����M�}����/�Mox��נW���2�Kc����v>Pk�|I�O>��Ï0�����;xf���ԍ9Y�υ[�X�7�Q�yL��UB����~�Y~1��������&*E_���56F��ٷy�''R�]ݕ�<~���>��^�yi������$�>���bU�}Cg_��=1-)Y�g*똥t����[�S����VP����`{�������޳}۬[u���ㆳ�t�e���=�t�{���[��g5�>���W}5��,��Օ�
�Χ��ji�K���[���u�uV����0{!�w�ީ����F�&��j������Xu����[Z��]�Wx�n��|��@6��c��v��N(�th�.��t-��S�u)�0�3��0G�q;sV���nb3~".՜�f�u4]��fU�={ �ye�ly�5���%��h�IֽϾ�]��7~�%��g�g�w�
�׾m��'�?�=�!g���;�����7����<�L��2y�|$��>~}>��積f�נd�7����#W�o�<y�-������Q辶���;���1���h=�l��=�7��=�}���~�-�:��S�齚e䛒�*�����j�����-vn?�z�Ֆ-˥��O��^��G���\�=��Wޏ��ow���59�5�S�A��!HU��CY^�)C�}'[�ƽ��x��	_���V̦���6��^ڡJ�~ÌBրL�҂m�����}b��vٝY�_�w��߫��K��g=Fs�2��{�o:�V���j�����&��Vo��{Y�A� 
�N�/;���]dO#r���%�z�s�t.�<K���M�aW��2�h�냒��A�v��F�ۖ�w%P�׃U@_k�3�r�s�F��]]r��a���<׷�1.�>o̆�u�u�Ć�͙W�6�Aa.��x820���jv�`r��P'w�:�sN���6%X���W��ש���V�	ȝHQ�2X�5F&w��|}~}E�Tg�ܺ�X���)Cܱ�j�{���OBv�{l>�*���{�.�Ш`�0m�l��GE�{����2v��H&����47�7�ص��y�Ic:		cUmG�EfP�;m�5#�8���=��-�|w;��j�ɋ�7ӽ^Ng���/+l��'�Y~�{+����:q�W��ov�����xk��L�c욺{����A�.vD�NbwZ=w����q���u�:Es�VB�sݧϱ�H��mo-uyAm�Ψ�9�V�ۡ0�/]�Y��F5��Zc���[�{�w��1mfP�}�����u	7�̮��U~��/^���~�m{�/}�܆�����+/��sѡ�?����I�T���y����=<yy�g�Sg��g�;��A} WV8[�(�r���T/�GlP�S�jB�̆�W]�`'k7���!�~Z�2;�S�0T�e�����;G���n��
k2�pF���з-�o{m��tTj�aܿ��;*s��* M�sܑQf���s��N؛�oA���OjmG��#[��ﾮ+�TC}߯���������ʶ�m��F�Bl���B�������cz�i	��W]�U*t����ھ�fJ��{Ƈ?Yۢ������%2�E ��뾅O��ߧ;�Y\[;��)�:���c~��/`mۜ�@�,n�6���Y�CY���8�Uw8,���Ά�������ѓy���/}I7��AL�x����Mc�z0�\���7�ީ��\	���ދ7��zu�{j@�������Gq�cM����&FvEF�7�No����v���{��W�Y�m{�M>r�@3�դ���i��N\��Iݝx�m�'{�zI��Ả�_��|	��Ǧ5�~�1�[�o��,M�ྮ~�������i�,���K;F{O��]�w?}_K[T���,�?{g��ݖ�]�m!�5~�W�;��r��+ٓ)�#M�'���{��2ݓ�x��8�+tn�5Q��7��G9\��]R��n�L��� _Ty�����2/4L���1!�\ �u��0��Q�׻�nѣY�Ơy6ev����\>�tyDI�h���\�{5���0���R)�J�>������o*������PG��>�O�U�j�P����~���jO;������6��P�N�p�7�1�����d�~����=�;���4�kj&<w����L��UF���E��7�φ�N�q��(���v�FwP&<��K������i�*q��ޟv��H�s^^��i��y�󌭚���9���sd�,���Vlۏ�SW�� �Yş�4|����{����J�v����ܯJ�f>��������m�[�L�&�G<�2�Ե�Ӿ�|��§�]#�<���u�\�0�g�;��FH�~i�b(ә����'��{y�U���^�Q�ݫ8O{`�II#�K��ͻ��;��
��;��o�{m7Ԟ�|�,���AA"�t�8����Wp�\�C,��wrx�:�U>�*����/R>�麼�	��<�CSv*e��o}�6P��֔�$g`�`��F���y��j���gq��3��}�\(��'VZ��d���`����R�a��˛� 1��Pu����� E��v+U���q
�:�=�cWVn:t�z�}�j7+����҈AQ-�q������xԙ�뻍��ȣ:\�a鉘�m���$�O���ijY�f#�٫�ʳ�B��ץ�Sj� � �^������1�u�Dn�sg"Mt�1w4/|�����/��l�*�����}�k��\-5t��@m�@�3ۤ��ͮ����0��xb��|�* �s��)��S��/|�юT�'M�k��{��3�����/ٕ�0���>rr��S����w��+v86���m�\]+Ϟ�=�̚.q�J������Rd���}�6<}��>O�,�BkG�ߢ�eO%���(�^N�`V��}��;H�wY~�+���t���� �$�ߒvt�󽅐}Vn�3��_�d!*�6W��c]N^�3�~am[�[�[9T^�����Cۘ�o��������7k�ގ�Wo ���|���.$�3����xx��0!+��zɍC�ȿƐ��ڱX
,�h��W�wb���t[2��F�A[���F�qB���!��2�׮<��腲��p����L�a��(;���鋅0r��6���y��֎{QG:�aV�9q���6������q���k�K�����ɺ>��9:���4��p݇J�b�D�;L���$�v)ٛ#6#LJ�/f��ze�ː;�ii��16�%&�+��q7(�{9�Qw�5�󔪌�(m�Bɧ\�
԰U��r�dckmZh�ndַ=���s`7��6�,��47�M;U'ٙ))��62�`Cu@�b�O��j�����Tۤ�_dJ��d�Tu�3��`�]����HC�r�^�Z��bhJ�Ӊ#ͽN�u#є��XԞR̃{�7���~�&��S��m׊��K��3zN����N�����!���Qɜ�h����ڛDk��e��e�:��9nӒ�5�X�n�G����&�c�V�`l -���|>�k9�����5��*[q��"r�"��N�ǚ*�m�7��#�TȻ%ژ�&cH*T�
��ӏc�5��&^�{-�]a�gN7��bM�!��61�V�����	оuq˭+(�`��Ӗ���E�z�c���SL����Gua�����Ѭe��C7Vu�*֍P��R! (�d6�1�H_1���}=:�B�̉n����o�_��ǲe���|r�i.�٦4����2�Nc��wd�"����`ޫ�(Jخ�Q[�Z��z�
����`勬Hh�Sr��{Iس���ά��;qu�d��%�j���a�܏�w@����})��/.����*��m4pb���@+�0�jC�Ty$�֑8\�D�f�/k6C;7^Φ1�n���h������뺋���N�@���3�t`��9��%)t����ҹlK cI�2\�c���(�7:n�ౚ4y�Wd�,�u�h[RF���S4
��1BBh�����U�[wO8<�(��:ۭ]�cns]�f���wK��<��V�W�%㲪d��\�w6�`s@V��p$)jcws�K����b�md{o�j��MҶ����!r9�/wpR���9 �XLX��^�yr,რ����W^׸ĘP����.w�!�X�Lu�]�b��ʻ��`��-���������]���Ϊ�z�=�D:8)՚>�9u��Qc��#5�g5q���;���\�ƅپK��<j�B��\�.@�o{҆B6�r��}Zػ�B`96BK@v˅'�BTY�Μ.M#8�m)�����qFs���!hN0��Ψ{Sm��E��r�ԩ��>��@ ʃ ����3���M"��W0�9;l�ǬI+j@k3������<~?���3�����M��((��Z)���,���`Ȥ�)�1�M��g||}<x����|||q�]g�yyNa����M6G�ݘ�8Y���م�����sg]x��x�������������'���n��m�}37��$�9cN�s$6��f��9 ddX�4�9���7_v�QC��9f`�9®`RQ��Mll��VMY�I��lFm���m����A��ffPbYdd8YQIXITY���,+H��Ƭ��`V�e�TQaef��d�bO�O�=bc�0����̽�]��ن0��r�2L�*��,�4�c7�2��ss/d`P�sk"�7-0��2*�s~g-� )r��ZU�A���C��In�Pifn��Dۅ��[��h"�h� ��(�_�ʺvYQ����o/b�˷�d!+Ii���BFM�����tft7kH�y���z�~��>g9﷯��a������>�^�ҕZ�<����n�@spaI�~^�����8��7@�7�lw��.��fg�쇨�>�ަ-��0���;0g2������x��"<,aSe���Bx�	>DAkWf4�v�hx{Xw�fv��������L�l�-��<Z�;GaT�R2�mq�og���笽O:���@�����˘z/M�>�����𦘸��&�x��o�%>��,�ɠ��[��pPj�Vۦi <���O/õ�1P숋�<���yRY���f���g�������t���r�p�ٙ!Rt�|[�����s�b�Z��9ճ-���1k�j����<��3[XU�@��*�v�J�|Po_�p��n@��n��v��M's�yO���[J@�p.�T�>�k� �CG���<b��6�pDB�vW����c(].�C e��,j��������Ux^ׅ���	�cd�j*�F�Bew{Ί��v�opjaǀO����o��=<�;N�U\෸�9���8�\�s�/ə�k۫��H�1��7�dz�C �</�4c4��r�E�ɤWt�|�LX�(�����ڡˆf��B�Z�X�1XϬ�s������$O^�xtӬt��k9i��W]�U�)�T�+n�m�6��F����+Rg9�۳4[�Y��ڜ�iNO�2�D(C�S�Y%�@���+1}��hs��cU���鿾��|~#����2����#��z�Qy)��H=1������[#�"`w*�~]���$��1D�|�����L��N�z������l�x�5q��=�?��X�G�5�ְ�IՄG��@�.Z�&��%�vih�ͅxy��n)I�.,	��dC� �FW�i�/�>��@8��֭}/�8������ssJe�pK=�H�cU>0�	�ios!���m͐
q���׶�uɠ-��P�,IaZ�oq�
��*��2P c3�3�;��?)LS�sYؕm�8�$v��kzۋ��3�a�.6u����;�H���%��!�)wWɂ~��^c�jDҜ��Ր������׶��{�s���tyT�e��h�m�?|/:~'�n����P�!����	b�=�K�2g�>c�6����^y���{�g�4�Y��+�!���_�n�L���,1�f�US���7�Ӽ|�1�4�%zZ��7��0����N�Z�\l��21n�����
h��A���a:�ƌ3�g�l�H	ߝ47���^�����ߧªv.lr�o*Խ��zK�t��L���l�1okYyO�\�NU��MCLC�l[W�?`���+Ԟ����D��̀r��źe=��X}�.�!���bՌZ̪��'P���Y�����f��9j�C�nA��w��p.��v��U�R�[��K��q囨�=�7�h�K�ML�r��	���m��o�%Ӛ��'b?�������>��#$bH8S�9�{^�ԮPTG�E��!CQ�^@AXi3����ɧ�t6 oa�����%���L���R}��}�/l%[�-����(�NfȂ�Ľ@
ڈ`��;"��{o@�@G��2׉��&����X@�� $�`���]|���,�������܎��%�����۝{󾷭�4�2���cL9��@V0�CNtx3js�U\�����M�9��m�s{Rx�\��EP�P�e|6���uˈj�@aE����E�y�͍
}�Y�3�^�[,��P�U���)����_Ԁ���Ҡ�(�d͗�����~�`���y| CH�Z�=-8��x���dSz��q��Ϸ�ݼ0Y���Ka����ϭ�j��@�؇F�����d{sڟ�U[l�{r�)�\��P=�-sb�uH\m��P�O���),�@�]��'{{e��9z-����$R���p?g�l��_�z.�S���Ld��Ԩe�= Q�����{h
.T,�;}�ۀ�Ý�x`�>Șւ�`�hx�~S����7���g��?N/��q��Y#���Sډ�E��xގjF9�{y���Ԭ�����8�'��1�V'�K����z���~j�����6�AV�-��X��3������x��W�8;+�ɽ�O[2�Seؙ��u�I��:��ԺNR�[S��ә�>�[�� Q.T�Ӯ�}��GE�ҳ������3i_c�8���+��|[��)�qLOC|{�Z0k��,t\8V���y�����y��k�w8nMt�>� � ۛ�+����[3z-T����oC?�)�}uQ��a���R�.ti5Gf�;��)ȝt5�8�wj�����߁���6�K �ޖ_��-_��+xS�����R��jؚ�(��̄���Q bȱ��2����(t]�D����S0m6�捬چ���v�/3
������Sıc��=U�O9��)�`�����,j�
���%t+����j!���e g̆m�h<�+1+6O�΍�!���As�-B�j�R��h��t�.%@���;�xv���׾X�o���ں�A4;��Lą5��"��0-l���.m�V����4�c��(��oaULK�(��K+P*3&^C��wj؈	��򜅝ٓ6節����2�A�<��s�*���J���7��n����
h�{h�l�gJ���K�DI�(ʇ`���h����C�o���{�qv/)��}m�Z��={�bU�^��_C�~�v����v˴���tC���oM�4 �<���9�Xs#q���}�!W�~��/k�Ǝ���v]f*�e-���t̋n�a{����>�N��l���X�2=7�&���0�*lѬ}�ĐV0ˬފr��D�}gY�1�b�2����HB��73�W|�;߹�������~v����_�3L�2~"t��6o���j���$��
�C�"|Dm�;ѳ�����B���6���c�QV�Y�j[�P9�:���02�0NlLh-{`��}�QN_���Κn�]͖�ܪ)��R�s�1��wmx�-ɴ�hV��;Q1��W�)ڋ�y�[��Z<����zy�l.e�Za�O���Η�ƽt!@�C�J/���n�cfN��ސ�ƾ��&'��M���a�v��'��������8_�桹�s��VSô3��\��4�ߕ{�P<�^.�sR"���\w�C�*��ӹJ��^�ֶ�=�vB5Jj���QX�v�^̿D�a�(��^n� ^������k��չ���o�{ob9�<�*�{NW�㜁>�5����*�y�7�<�/;-<!� e5f.��=,}������
��wѯ�X�?r�AP��r�z���QL2Q�bh�ﻑ!���b�F[��/ 7z�R���4�c�m��計�W�<1�J���|��>+��[���P�X �����T�r���82j�ɶ�ʦ�+k¨b����g�1�/<�_�М��O�ua3����c����_ �m�w�&�4u�R���tX�U�щ�8.��^7��4n�1�X�Y<8�%��5r��V!�i3!��Gd�7S�L���y�P
����=6��H�j�
ۖ�ȲP{�ߩ�|a�6�{�w/>���p�翰7Y���L��R�F��"�k�Nc݂�Xk�W�!��w9�d1�8�#��������ccTb��߃@��qGs��R�=T&J�h^V�W������~ꬎ��\�~f�|�.�>����2Li��{j/���������g���{�<�)֠���b���=L̎�5*I��B��{ݎ9�����7Pù�v4c����75c�'�0��~k���Z���m�|=��_Pg�݊�ʐ5����a��!��l�M,�8^�in7F�]�7����7"rs��32����]��&���d�Ǖ��_lc��y�A�n���E.�ƾ��T��7��z�~�t=N�/zEP�<�/�Y�~���n L�H쇷�wy����ٛ�Af[͉c��]�8f�^N}�-^�LPǤ���"w`��6g��B�H|�&���SAr�OH6L]l����`�������Hu�1���3�������aB�=�q"'m���j�S��6I��xg���Џ��;�|�8�/0���`�e��ۦ�z� w��W5HӉ�3*�盖��ư��N�U7�(�r�wR��<�[�����F�u�Dye#QE���f�Ug�w)F�Z��-5�}��T�g��W����||"Ҳ�m��u,�`4�����7�;1lr��r�o0�m�c�j:���C{(�i|������ĤA%��vw�o0��h�IP�L�v̹�ȹ�4ߖiaaO;��<z��M�5M	�Þ]��� k@|�O�?O��{��~ow��W\����܍<���fjʍ���^x��b�C_��ê����C�K�ّ1�S�[����d�z%�  ��qm��U�� VA�9��#7P�"Z�˧!�yMÉ0����(lW�%)z�x�Ν�=|��fd
B#r�C��^��)V�1�eE�-�WB�ƪ��Y1�YبjcXm�,F����'�/9}9�+��~V���涭�Ly�����PَE�	l�|�x���Y�_ὠS"^4}���0���|��1�ƧL����z_�=�i6&�]hw׷��j�I��gV���ѻZ�b�/�(W{&EA{"A���k�OiUM^��]Y ����F���.��V̩�B ���[�t�3�쨦\��J}�H��mɜ>�*l��y�4T&�xb�)�}���v��}K?��k��VSp�J�>Ӵ�P0[���I�.�n=c6���pm7����d��I������&`>4s�Q���0$�M���g��K�̊ln�gn"����]誗����t�xrC:3�z���8'������[œD�+R�ָ��"�68�v5I�4��q[=�t�靽xl�'��I�Sa��s:�C n�7�k-�p`��<��z�H�>�2���a�q��h�Ne�H{Xy��`nxucs���fV�%��!8w}�Y�lz�j8��y0���s�e��|���)�]Y��,��|2�w�u��.�T��h��XO��Q��S伲��[Ȩ5h&v./�x	�v�b�A��$�/� ;����F2Ŵ'�=.G�:�p���j�k������5�FKy�魰�r��a�Iy��|�	t&�&y�����DCvtm/0������]���u���7-@��A��*y���P�l
.w8^�lږ���<�z�9\|���
�!
c��z���7���/�w����8Ǿo�h���,�;�����Z�u:�rf�Jg�uG]���be�"G��ß�C�P(ME�Ōq=7!�� ���� �\����p��Gt��=,���t@�}yM��fQ���l���Mkڠ�sT��i���f�V��A0c���%�6>��h}�/�d	/�v��nb�]��*4mw�C3��{n}�??Ҏq-uɼ���)�R�r��a��bYm��zٽ�^��*L����(@����%Qd��Cs�Z=
#9M3x�C�ffJ�rR A��P&����	Gz��cY�����ep`\����H�7��-�΂K������L	�%������?/�����$y��0�f=���7,]��ͼC�P�̲�e>l`ި��1��t�֪�Uу��k6����@�����n���Qy�@�^5���β�	Q��O�fm��k+H*/�z�\UC��$nf�rU�v�iKo1^,1��t9��>l@��=
��.�bF�1*%�TSY�8�E�ۙKk��qJ8�kA8��^K��F�и�]��*W8�1���_��ɵ�'�s�P��i/�6Z̲0�f���X��g@�M~�)��z>{�(n|geu��� {
V"�[\�;�b���G辪�/fV�}���|�-�(YIT�A��~���C�>L-c +ڇ�'���鷲�[fԉi���Q#��v��F[q92wT���-1̻c(��Fs���~Lh,2?u
>���
U��"��x�j&|��MZ�9�4��ь���m�kb�A�3�4�;���ȃ�Rio@�0�����z�!4�B��g�[^���|Bͥ�U�oO��:�u����HZ�C��C�Ӯ�ī�m�¿c(�\��}��hj̀�ǙNk�>1��C��6����OHʂ0j���(40Ν��#.Q�e�M�;��)���ɺ�B����#1zfT��7gP�����������>ע�L�
�G�~*��7I���i"�����nc�~�IN�%�y���Uy�-xuҲ�V�����4�׏���K�5�t�K�DM��5:=���rNc�M�)xX��X�t'Ϥ���ߝ���s�;���'��ɒ$����%Lߗ��B���!�^f��D��(kk��xo���x���/s;��s�T�q��svW?#�=�f�h��m���&ou�P�;礆�$�d���?�(Gp��d�P��m�o�Y6%'w�/?l�x��͏���CVS��Qm�ʒ�*���4Z_{�A�o��0�z�Մki2��yׁ��
���b�(Ĳea,�m����v��z|\2P�T.��ɁU`��'W�;��P���2¼����teo��$�_�#7>Pu�4粦q��e]�v�Ӈ�� �➚��˵��4g&�p�
QtT&&�*�b��-D8N��~��>\���y���TYgz}�����Ļ��� RS��9=���N��5���6�~����C�NPۓ�bZ��>=��P��|���g�߮
|�~��e��u(}~G2�sY�f�rᙑy�s~g�;������^����̲`���w��{��N��>�OKfNDw1N@��*2O?K�M�K����9���u�oM��T)"�PG���B��47���l+����Ϛ5�H�t����r��eVjͷ,�'\��Ǘ��r]I��� �f�v��G��l���ٗ���v	Ȍ���"����	|Ջ�j��A�<2+��K��T&�n�=�̿�[�����K���sM�8�� �L��]0��U�3����wZ�X�3R���isL_4�<�B=�NH<q$�C�֕1.cv�?;��ms��n��@Aǔ��גC�d	_���*��9~K�������:�`4�@�t&��-)L�=Β�В�@{bS�֬��_tEF��剢��,�-�l��>�%I[=�I@��z��=��ʣɾ|Zǆ�YDl�	>����%������[g-Wh]z�jޚE�t��H ݴO�v9��\�9��ͻ���yZq[��[gc��X�Rb/,�}MC5Ϥ+��荘Fo<��;.kW�l�2�!�F��Ob�[;�2�f�8��{��Ph�H�-�k`�:W%�q[��
��Ϗ��} �5I
s����oS�˪�_������j��؞Atf��&dB����voZ�	��t��v�#&sV�9!U�t1�H.��C42�/1�%ǝ7��J��J�lcZ*��0.r��;�t���%�4e<�x�[��Y�rvN6�Ԇ�㦗u�(]֓��T���c��*�TSF
���/o\pAo���^˼�v���q�w� K'O��WS�K�����-yT:���뷈ϸ�wʌ@��W%ٝ��$��B8�,
�(R-�D&��3��ｙ%`��T��{�!��-uY!5X@؞[ms}�WyM[�p1�
"ٛ�wVc�[ejő�����{��D�="�+ \�|��ٮ8�rwm����&Mb9���q}��лv���N�t7)�҆[�z�����J͙B�qV1�}���|��&������w=��g�-Υ(�(�K|eio�b�ҩof�\�P�bN�sL#�%�gC������s���T�Oo����k���oQT�W���Hw��
�d�3 �Z�(��b�4�Kz�ͬCyNژ��ј;+�ZXcL���T��X�1��`�4�i��XK7A�q`e�k�٠��:�96��H�w�*M+���5��m
P,��O�Z�,r�㜜.�+۳W/��r�y���h�ׯu؁�L�Ri6T�P�t�c/�����C7�
�F�\�L֗Z)�r�˒�]�������uD�M�r�fe�4w��YD��Fj=������%����Wk@�k{f�XrѼ�uNl��3p�\�G*ۈi�V AlU�7;g�aL�c��F�w��f�;�f��鎌�{�����5�]��n����αt+�ec�m�M�������W�Aw�3��� KG^�Jq&����Y��ٱt�-�RZ�2�h�{o�ѳ�-@�H�N����.��f��# ��U��4[F��n���V��aU�-�"�r�ܢ���I2ʍd�kr���Eʬ�32����׏_���Ǐ���3���Ȼ��ya���n�;�Y��9�z�E������2��2�j-�c�l����vЌ�q�_o������������q�={FNDFf^�V����EF�N��A[e�=n��=n�9n`V̈́�:��~>�o����|z��8����Q�G�f�-��1�e�-ֹ��ɖᱣE9�Q���2)v�:y� �72=�;a:FEi�U����[�Mi��V�e���0�������NA��E$�Q�Y�F8f9dFa�faC���XE�m��U��	���d��Pd�{���B��"2�,�2rm�#HH˚�W�3�9/�t��s-֌�2bk2�"��2�#$٪�r�f	�����ٝ�7 �(��a1U%!nr6L�7w3K17#2]#$��4�L��̳,�}�374�\ၷA��HD��"�(����#$��6�q�I(6L1-���ݯ�����y��tw�U�u;��+2�%Q칙Ϩ_ܮ@gۼ�7K�CF���ܷ�f��M�pa�0�Q��b>Q���.�)�?�b8���A	L�R�n/��AIC��M��A) -�
P��3�A���-�E�b�/�d~�~!��B<�z�=��zfת:����0��fSI�D@������Y�2O�ҙ��g���:u�ׯ�Y�՝�]g�	!��<���Dm#���&#z�7b�a��g�����&/^��l��)�_��K��r����#+m��˹Yzq�4[�0mkw>w��]�4(��C�P��21P֐�r�{z�L4�fB����ʘ�̔�hn-�8�>��^4(I�q_%�(^_�Ϛ�H�Y`�i��t(�}Ê��2{ީ�d�l"ڥ�p���"�H	G��Wq6Ҟ�˿*��恐�D�\[rz����9rS=��m�ђ`/Ywd�$↨L��8��b�CX�7��ͪ$Cμ��υSKm�vf\C�>8��1-T⚩šj]���C�0�i0!�B�w�Sp�L÷���9�Oߌ]N~�t�����7Wx�2��X_V�y2���e7Z�޷��X)�*��l/z�
��7;���2�	BH4�k��h�6n�Y��?��]���E�x3N�&���Ly�1I��f���r�psx	ڽ�O�D�^����8�v�����W�l��!?/?<>9��������l����w�ժo0�iZ	�?�Z�1ڱc��+1;�N�h���m�L�L�ј�
.�Cm�Z�}�����B>���ͪ�[�g]ϟ�Kݧ��c5���w���Cv^�D�Z��r\)*��6�C���giUu��>��>?>?|�y������a�{�����%��#O�|�����׭fP�Y9/B��4����8��?o�L�;�(m�y��fm)�z�L��\��O����g2b���˽���t�尣����K*+��Wc�bihk�\�z�û�Kqv3	������&kC"2+���`,.�/p�/��WZ�h"�T�y�²|R02�qq^&�sH�d��0�>�֗ki��Da�[��:d�u5�b�P�&#�7X�شhUS��e�󟾂_���>{���b�]��-ֹMIٷ��h����9�/Bf4'�ye1����EXԌ읭�
��%ݸ�l�!�� ��vi�1����kg��l��,�g��d<��`ᵯ��5�z�QD�î܊	��`��ދ�&D�f/�����z���B3���y�
ˣ�������}[����x*���vT�e��<�i����ht�@��������7���3p���h}gg����F^E�˫͕{�8b�[���;>����.Bƺݛ�{�@-�nF��5�3m	��|y���TK/����"m�G�O����vaj�B&e�Ü/���	a��j4�(��궶�u�.��35�ư���!�@gS��7խ�[՚F\Q�!q��v��E��3�b}'N>�s�݊�B�<GwQR�lkh2h�ЅbN����@�!�r�R+���YŤʼ`�;g��Ѭ&#���E�1�[��2x�+��_��.�xA��RiT+���)uUp�#IT_!ë����U�#`62�����w�S��)���DBl��kq
�*�y�w6j�(�mC����F��v�����)��(Y�� �����᱑��л�g�8� �t1zge]Қ<�8%Kۃ6rb��h�ތǠ�m�>�?�J��-jju�t�
u����w�f�!��q�_J`]�*ª�s��l�%����.n>@f(k��n�@|�Kf��'�8%职��6�:����It����&��U����f�î���mBW����ܵm,��e�H�[m�`0_t���R���<^��)> ڔ��FM��m��Pך�Q�ָ�2�����0oP�g���?4��L쪌�z��%W'Cv���g�&1�ef��������_��Ѱ2A_�W��ό�]'��`\� �f��Q�j��s!�������L1�A�9�sbcA~gg�~�����
���8�B0U{�R��>�:�82�{���ޭ�S]��
̰g��'�44��\zUi{�d�jn�چ���;�=9l-U*V�ːdݚ��`���1u��yF.y/`���J��\/�"��9OX�zl��#���c�T!� �a� ��KS�\��Fi��T��ɫ��P�Wԗ���x�F˾Ais���l�MܼEM��@�"��~\��_�ƒ�`��k[��e��ڽ��:}[�/:��5�z�S�ɪ�0ݭ�y�5ߓ��	ɇJI�硏��l����-�^��N�<��E�۫���-�9G������v��͐�v�A��Q���i�I��p���ސn�Lx���������=-���J�~�pCzl��M�圢ZIG�L����{����=w۔��*�ZlK��PMfO+�[�tzn�	v܏�$>���ͪ^��p)�h�|�\z�K3篕�B�u��O�����]����^��k�j�v�."9�",�4[O��U�+۲c�7C�؍�sx�� &z�\���M� �\K-VbY6�+nۖC��mMC�O��r���iJT*2�����꺎6 ��grƝ^��vդu��c����\O��P�� ��{��~�m-}�Jg42܇dh4y��5����~���w8��+P�:nᣮ�d�l���b��i���ʌ��~Ó@/�Z�J(���V��GK�Y��k�Zg-���l���6؋y�İ��}wUR��(1F�&�������y�=i�Uv��L˨s���k�Y�"N}Qom����̄٦����7/.w�2-l�]
��'��\�( ���a#������t_l+b��~����J{��S��ig��Q��׵��*?RXC��>�y��j������J���ۜ�Rg��%��=(�O�E��>lu��6��i�}Mޝa"�"�%�`H��K�j�ҝќ�x��&ģ&'��D�ڕ΁%����A^��m�#�Y��샪'����^���P{S�uMz�D���3�P���\9o�Lg�a#%�����,h����whw��3��	�*+��`�lqz���צ��<�/�Y����%�sS��?��躌
�*�E�~�Y�M(F�Y�`4Q�Z�ƣ�zN�`X��I���SM��׶��'v*5�9����"�5�0mffk������;y�[�?��f+>hjQ������}��~�����!�����J�!^��)��^�0�5��[�|��2��kNd)�|�fdSG��▼��ǅ۷;�g�/u>�/1��zdO�= �I��SBz/.�i��5��"&T�	�n]���bN���o�����^�j��N$P�ͯb�F3H*�vI��ƿV����g����z$�v�~��?,�]+'ON�3G�G�}��oE�A)�}d��W��S�cKk�|.���u�l#���(�D?3���.�矑 w�ϗ�6�s��8��QE��=��.�	�y�l���|���w߯x~Q_��$0+�`0`L�JAR�E���~y�w���|3�<����ŵӏ�Z�h�ds(zFm��D��Ӑ�>�7*R;�{Q�/&VnZ{Rf�����Ј�p(K�;zEE0�	�mK6Pi��fjU"nt.m�b��𾾛��]+S!�����)��a:�������.1�s�M#�������;o��{:^9n#.l܌&.�Sybن��^*�ӷ�K��5�S�[b��7?J�}m�0w*��&�.�c��ImP�}Ц`�۸0����U�;���FEȝ�koPdɽ=��ºg�t����0�]�(���}�I�1L�����o�.��|V,�+� u�t-�g�6U�^Ow���aЗ!�:�-�FCΙM�=�%���>������7У���E]�o5;�"u�%n�:CCBn���>���hȗ�\������,�9�a�Uk5D�׹n��T{	�T�˜��f��&!���6fT�A��o�*Czx���0�)�����RN���'~��n�؇~�I��zx��ɍ���c�<&���H�I�:�z�m��%,W�Ux=�4|CP�v�����w&�q賵9���3}�� 5��HU���v�o��޴���5p���զE7�����ζr��fQ��[V�l���b�:�Nv_a!�zv�J���|����8P���h���z� �y���(bK@����?=����ҹN>r�77�Lأ�������\�ó����N3�;��u�n,�C*�u���c9}d����oAj�L�d�	3>�=_g@N�F�#��߲���ڛgrb��=t����AaY�/��-b�1�O�~�^�hY�A���ؿ&�a��k�;��fkN/j�"�'�'9�1c���;����)�c�6� ��Sl�FO>��&�ɭ=�]�-h�֗/�&pZ�E��~b�;�<#�]��ܟIbޖE�m���\S�Mp�}��;fצP++�.f!�q�[$3���=����⚤TSt��`���58��hȸ� �&����
Z��YW+�j�{�B����+�,|D�%G�(�Aʋ�qʵ�j���*S@�}׋ �����'�Q,��U��*�`ŵ��˞�
�X���O��������+�P%�RmzFh� ��	�)��I'�}	��7u�fv�R��q8���'}�&.�7%�v�EqA_d��D�}ס���lNu��$�aa*���M6��j71��햏jh8Ѕ��Nb�����z�c��o"փY�M}��Î.���,�89YaTC�Mc$I��O�^]>��� �(@H����v:�x��B��y���$q��R�͹Jz���4�^�:�����s�S���7�>�߼�ۇ~v�3������2��� �J	���?Z�V�qmr��'��	��W4_t���JP�]��}m���sپu�H��]��Rځ2u��Li��/C�����6�����]#�����.�����s'g��}�M1�C0���`�������t��ۛR�w��h;�y��`m�;��L֟)�g�&5k��-��d��	��o��7-��c�|��_���gx���àq����:�~�Ţ��v�o�XD�j9�ma�&���u"�y����i�`v4
;?�8Ϡ�7����_�c�i��~c�z��iߣϝE��p!����&���U\k��)Q䅓�?H�x�H�C�����v��,&w@�H1��c�:�è�u�3���&$e��)�Vo��w�-�؊&�˴*ɖx C@W�.Q�͇s+�7{(nc&��V�.Օ���Jqn\D��6\Q�������J8�`��V{���"��+���y� �����E�=V��,�|Y��t��؛�K��,�����[9Mԕ��&]sw�;/�v����t�ܤ�Vn��2Hx>���JhvF7�ז���m����� 2���F7�N*n^����Q����.������1pN����U����_���z��Nٗ��0�׾����0���H"�
�
W<�g���9�3�iȾ{��O�v��Q�#�H�N6�$�-D	�A �E�	���Y��Ϝ�q����Jm����k��)��+�dDHB
𠧸�5W<sE\My��=�\ˢ婛޺)��F�6�@����c6(1k/lЖU6��'F)�xk~��-Z".�qaP�A�w������e��qR�&��;�տ{�.|O)��*�e��tk���k���[�,��a�א�M48����*]����6�XO�A.)̚Z����-aF�8��̤��`��R��mWU�ơ�'%����l#
�O��'�l'���C6Z��b7���nؗ��Ol��Cb�)>oyHց�F�e��y�v�a����̷�,c�����Z��X��K%���D�ԭ�B}]|�قn�beW�D�L�5�c�[O:ȹd&a������n��~i����8�KV����L�����`s>����+cݝ����(,���qѮ\�zn�����s�����4�'�F�g�����6�5�=;>�&z��{���[����맧�nr�F3`43��\j1���"L�݂��8�iƅгZ�[����+7C�]C���%T��ش>��ؕ/#�ӏ*�*]K�V�X\l�Y�EtM��,V��p���'zZ�y��I��E�֎�S��/��\���ײ�z'+jm)Yئ����.����w��|:}�]�Ϲ�{Ͽʈ~ \QHeP�Dh��>~/|�Y��>}��oϿ���ɞ�_�~D,$N?��$b�"DV�WG�mv*37x+m���<��/wB��G�Z�ۂjp�/" �|����&!�H:s
�������i=�يߡ��&3c�T�7�P�щܘ-,��b)�=�臭k6(͚L�Df	N��c)�'B%�cx!�|�og���]���6>�4�1W!����>|��nl�iwKlx"�.��+8ˑ1�y�^��5x]�=^�f�r��0gśɓ�z*7�_ûHz/�e{�:5WT�0i�#�ޖ^�����e���E53�
�X�P�&Us�&��Tj�F���ۘH ���J~�ڮ���F� ��39OR�����.�G���m�9����,f�� ��[����Y��0w:ߏ!�#d����mߩ���|���T��|l���S�;�Jj��h�w��c~A����M��6D�L��)�&�+�j�g̓��L��bB�[���T�5����; ����އ��v|d �w���FV��#��<��)G�
G,m�=[���j|��xx�׎��l�"�4*���{mm`s�Z������\.�5nXOk��'�y*딛D��u��'n���Tw5w+b[V��*Q��}yN�� +z��e:/:J�m�0� �Ug0�q�������cNW_^RL*O�T�}2�I4��er9���0�(�6��V�B�M�P���w�m.��$������һu�'�gLuEdں�qR���Ǳ��v���̴�\eM�� �Onցη[4  ^ӌK�V�����.�-љ��{e9�MS=S�E�=���e�Ԓ�VŶ4d7�{&�9��X�EwYCs[O#���߳6�VLe�9��f���y�)�������B�m,C'.�@����̫\DU��:����Fq��J�mu݀xs2�.���sM�Ǧ�n'�W�IG��p���X����ۜ�f>絕��[<���ӟd�S;�Fw!�p8�T
Gw;���9^�����b���X�s|�U
�l(1wq�������G^gia�nB'V�����H27k7�'��n�urL�3@/+``V�T�w`�e��cr�뤫��=�CrH�7�:�s�n�˥6���k�G{��;vk��L��)Ҋ
=�WI�k�w,�(���Q;�	r���f�7k���th�O�eLq58��=�]xi�W�R�1��������R�"���KdO�s�M��*_k�mӅr���$��Ȫ�ue�xa1���,��n�I���uk�e߁]��]hI��چ�4�lDU��_;�3��"�pH{Ȅ��^�����ɦ�*��+����Ԍ5���Չ8=��oI������hx�o���ۡϛ\9�Ju��\b[��hEԦ�
��s+N\7b�8d��dSC}t��QE��-�n�lH��FU��C�]�iVwnȆ��W��e�gl�qZn-�\�p�.�d\��l�V�����k�ޢ�3ӵ���Ɯ]�ʚ��̼oj�q�*�h��3i_B�j��d������-���Yy����y/�����q�_>h#�Q��.��s�X��ѧmY�ٕ�OiA(Jj�@��$$����m���=8Sv�qS[=]�����E��imŮ����]��T^��nH�Fl�&�q�Zs��,˒�����2�t|o�G���d�C5V��N��:h���	γ��aԶ�04�ϴ��Qje�����͡M5Jξ�Q�"���<���ڹDM%��>̭<��N���q�rN���:k��:�LE��W/���e���2���	��.&�m� �w^��4����:��6������o �*��ng</���%�ض��ف��gr�.�e�+F@��â]�]�\w\���u�y::�%>^�m��d��;�z��]IR?��f�(��%���ff�ESDQ�٨nb�nfF�nD�%Q������N�����}��o�������q�>yDO|�2M�,�4��6�

��e�smu��+33"�3L�ru�^>?o�����>>>8�Y���<����̱�p��l6�؈�"�33s
'$�mn�r3�+gY�]||}?o����|||q����xG�a9�l�eA��f�Y���g�C��ܨb��#c-���!&�JȒg�spr�f��Vջ���a;�&�̷��f�FI��3�f������̃`����9e��fY;���Pm�T�`n���Y;[fa�m����囸�����I�feE�QfXd��m�o�6L97A�D�\�!��2ܭ�*��pl�����p�,�j�r��(����1�`�k�5\��r
n`l�:�N�S�}��a32S,��w'm��$��&��s4'�LBUǯK,���&\�(����tz�ѥ\������1��7-ס����8��Ւ�n@�L�*.wMn�@����V �Q���^��K��o�{mO�mO��ɟ��i0�t�n.�a6-^�n>�+\P�ܴC垺wzI�X��Qz�xM��[y�K��#*��q~��
K���&[����C{n���3�jZ|�v1�+�b#薱�ٜ�F:�q���2&��<\X�!t�$B���2;���`���(��}.-%��k���vm�q~n`�a�iz��OC�)��, F�*b;�=�8:ݜ4�Xy����F:�Ͻ�`�;/ʾ� �O������	���Xzs����s&��ıd#cX��|ō��/Ӌ�Bz��w�@��e]�X-��|�����fB=_�H6#�a�ϯ��>ZŜ��W*�Y0~7E��KC�\�����2���i�,��>�l��h��W�����c]T;Fdp5�ܶi,��͇7�n��W�{v����z�O}F�Y�=��ko���P*j1d\cn@>�-]Л!��^���aY�[�z~5q�V���`�����L�i�L�?�:�����اLK`�J)�d��s���uEnk��j�*�Z�7�Wf4��m	;��<\��1���j�$3���cL�*�.̡��߸�=ˈn�A�9(N9>��%��Fv�,v؏�{���nr�����7Y��$���s�%*��������2d	�"��`ʣ�` �y��,sɕ���sG��O�0�E�g�&Ψ�/�
wzzzc�4�kdi[.L"?~��jM�ó_�s���P��2ĕcm�b�bڈy��2�B�����x%z�W�^�W�����2ƆP�����s9a��)��UL��(��	ec
^M2b��.F2�e�f�>4�Z�.�wS�B��*��� sz���v�)0�9亿8���k��m�|�qv���$M,PzW1͋k�A8��g�����.8Bm�\����T�
�3��n�ډ��q�^wbU`mut��۽)��s/��׎u�y8�v��Dq(�D1�Jy�xj����>!vW_5���i��q]��Lz[,_{��]x�f0kNv菈�`9�^�{�yN���f�[V��V)��
P*9��N�P/c,s��Ƃ�_�p��W�~��x��&'�5K�sO��MY��Rn���q�?�j��w���Eŕ�/|T�Owӑ��O_sFD�,��I�~X��q�o�������{+'�yd��T�����[��_S�>�a�JR�����ls6W��a�t6
��jA_�N������vO0�����hg"=��&[��l��4Mo�ǉ��aa��%od��{v�v3=+�Ʌ�(]�{��|#}�W4��xؾ����������M����C�!�B�@&J�R4����lքGs�׆_�u^�	0�|�mBXi"C�H4!d�����KO�!��ٸ����
0�y�c�#ZƧ��#}�EL矇�m#�ŭ��7.����Ƈ��Y�9ؙ8�>a���0%�*+�P�Y>l8�������[;����"�'H�1��A5�o��J��<��ˋK	(ޕ|��~���g�vs]3X��\����zY	�i�}����;0�6�*Y�b���U�[�;6�x�/p)�lK�/��ձ�&h�΄�z�ՓlڟRvO\�fפbm�M�0��`�=Tv=c����B��k�z��Ļ��Q�L.|��/4��X��t��[���;T�kv�n�(��ju0(Hºz\V(��Xᑉw�����K���	���蕏~��{њ�Ӓ�ó�q�K;��v$�g��=�S�#1�������T;Spl��qGs��Ɏ����o0�`�(N��o<~QOZ廯�x^!��5�ܮL����l0���02��;�w�"5��v�,��\%�wﳫ�C���b)>n%CZi���;,��b����6j1����C���gi�0n�F����W?z>�<x�1M�A�J*��ݏe;�敪[w�� wP1�/m��8��o7�6v�3F�h|���.͝�uژb���#ch��c2��w��
p�V�V1� t���@���� 
PqDx3 ��Xc�ehko�<4'��v�ZR$wT�s�cH��F��Gs�,K�w�}a�tE��k�UG#�Sơ
^WsD�	t�VH��j�ݰ��p'*&K���ϳҵ��v�;��{�UR8�3ԜV���E����.�f
6�ySɿ��Y9|�_�=/��T�4mw���Y;�>�́�ڵ��G	Y0E�
�.5��kŏ���]�,m�~��_A�-�F���"`�o!M���I�i���\k��@�$N���5��� u�UǒW|��v���y�B�}:����'�~ash��b�ƽf�/����"�~�j��<��]o��5`�R@Jj	$���d�;z���}0���.ޟ"�O��-@�SBz�]�Sö��P����궆ʔh�_er�<��"��g������E�����N���f*���~� N0�KZ�5��csk��m[���aC�;�b2=Kո��wÝ|��0xz���;��HM���q�-�,�P�^�É��#�ހ�H�n ��%���X$�}�C(x�7�c���5���F��dtͩ���ݒ��z��9��S�t��5�^ڮne���#0e��촨7�M�V�.�`} �&��]�cmqY&�%S�i�k�NX\�I�b�Bm��q�O�.='WXt��������V�qv���o7�����=�����#$0��
��#�J*�H���D#0VچＰ����Cw�\�<�C|lO�OR���H�d����	����g1W-�oz*�cū�+�l�c�s����P� ��qw�N����v]M��6�ZDW����+Yk�]�9Y�qi��B�c��l�A�=�)>�#ɠ0i�6�����W]�L��1b����i]��=ƪ���^=&�U��?2�#�@`o��qI��:`��9E2��J}�H千s?I9St6�}wf�!��;�喽K�eϘ�a2s�m&�	���_<�7Z���e٘���侺�3ǯ���=,Ǯ�=q?h~ o-�<��3,��qpM)��7\0�>�r�[%t��R׫�ҘH[��Ϯ�!ųC(���ܧ�شhS�Z�"��œ�w7������%��f�]�nq����Ak�Z����lh`� ����ʄ�+Q޶eI�s�js�7������c���i��e�P� ����8��Ƙ��i�$�ob�/z+Ej�}�J��� S���ڄ��������zΦ��w<{3��x�I�B�[��Y͇�nǾ>_e�i�S���	�$q�w�Nk.�Fh
|�hŠ��l$M&��n,sh��>����zv{k�������;�5JӢ�z�x�sJK"��}aF�����xU1��3���]�^�"�A�\!�_|G��"j����ߗ�n���Dya�
����H��Q��\�o1	���i������y�'e\6�4:�~s_~�)��_@���y�B��o؎ �6�1���t8����6���>��6�B�R+lHH�?��멄k���:�jb�1o�m~���N����:�s��*j[n��)㺻5��g���$H�횁��z�;Kd���!3���w(�!�4�6�NT��eq\g[�Pн�`0j��+��i5"m�c@�b��y��w��e�����U���<^~�����b�/�IU���Y�E5��-�VbU{ѩF0�7g�ݱv7v�ٛS���	q����t$c�~ngl׫�Z��hs�a��f�Tȼz�lNf�h��kXvu�s����3�I�]�mV���T6�r���Z�,��c�k]��8�]0K�R��u:x�N_�.m{�72+N�-h8�^	NC�Sᑍ4ύ%G��D&ڰ ����9�.U���&P2pV�yV:uo^��u�+_��l�,L���C�lzmN�C����
�j#ig�z�woV���89F�u�����;e#�����;��B�`|&�+�x���`�tˡئ[�+�}���(f_w=Fۥz�]JS3�v_j8�Iw0F�D�n޹f��<����K~4J0{Lz����)W������ꪯ꾿�� 0 C�!@����$S �U{���0�m�$f8�H!|@=�P?���;��:�F�=��e��P�v�E�6��x���ε��x�qEQ�ţ�ӽ!@�4�nնr���Vt�i�g��d2�
�nZ���E���9sJ_j~^��1�^:<�.m��0�!��?HI�E�@b��]��
���I��:�8�̱6��ת�W�9|u󳧐j~'��a?G�T+yA��(��1c���z��I����{(d�2��9�Dn5=�扪���D��~"����?<�X}�yus)]��I���tC���\��N�/�N[�M���!3ö ��b�a�W<�� f;6Q͒��D�yE,���5h&�ô;8-��"G��G<=�aLp�Iy`��r�����~�̟D|��a��m�.+�c��N�p��P�m,�ҕ���S	�vmS�:�
��,z)�UγիRw`!Ϝx�k~��/���E0=�W�i���b����&S�6�!��(����:�t�e]Q��˼�l���>?���Si��)H��}U@}
�l ��f%�m����	��o]Π
,��>ԣ�>��g ��ļ����V��2��;ͫ�ܙ���Z�h��q����[�Xt*�WS�b��=��<�!5mW%ѵ{S�Gw׹��l6�.�;T�s2M�ons��V�"�^;�����,0��,"g��sϼ�tZ�l��xb��F;�\�W"]�\U&���l�����0	��p	1�%��q��
x�wQ�6`K-J�X�Mel�H���OA�q�%���m��ڝaGnۛ7y���� ��*��Wgik�0���B������'%��bS���
��9�O�;u�x�)�L���?s)f��v꾘�:�	(��+wT5��� ��dN�/���}�L�ē���k�i��p��W΄���v֨7.�o@��R��8�s�=y��|�劃��K�Fnp��t$e�j��,��m	x\���ns�ʑM^�ޘn��ɭ%�c�����1Umw��c`��+l�q�[<|l[����I<w�F�Ug��MƸ�Ξc�8���S���ׁ͑�Z���8�cV���|>	��}����ߟ�ɯT0��zO"4ȥ���m�Ve��n-���-�zC�I�i��^�vK�"q���F|��������#k\6C$�%��`��*�B �=��^������<�Gʆs%z�D� j�x�N�u�ߚ�W5����Q 'pk^�����W��s7�mL��o3�Q��,_���>�jk��[����o5�7�@�����ԟ��ӏxNO^�/'��b+h��N�<����VP�c �Ԑ}�B��d�XYGztr�3��+V��-t�������|�@!�2ZDJC��~�~>���*���$>����g�ȳ>��8�mх����>tވOk�_|ќ��Y&�C��]~��������-��� q��WXAU���7�� j�d��X7��u�$)ۮɒ��s��"��{��N7�vɷ���0�j�!uO�`��<#����2r}1�-�F�~���}�
�����b�� ��N�қ�V4��(q��c�N��u�332!�j���w*�Vj�a���Y1 �h���J�p�~K�������E�
�[q��ok����a�_B�i�߶1�o��4߿q�؅^m�<��>֮�º��f�X&�K�Tͅ���X���۳�N1j�R$wJ�ہ#^I`��+�-뛑P�o���jǒ�s�ج���f�}���[u��E��1Aנfy=�=6ȹ�Z��tj��gڡ%A����4�ٿVLv�H��b��N`���e�C5��2�H�4�^T	\�[7���!���=^���ٖ����)�=�&B�0gϲȎ}���l���a�f8���M���`G��MK(c����ϕsv��-۽�8��ݗ$�[���-T�\o������=���r�@�-����e��ˢ65������,�}��mMA�w<�n��3��λuH��}m)��p��y��.b����}�s7����|?EC�V 2��7�<�=��˽r�S);��r��[y��G�K�K���-B�~���F�n���Bn��[:�#��qq~͌O^J9��2�RXHZ�}\�]��Ş���y���\V嵜]DeGC���5B�7�^2����#|H7���衸�z/��q��	��� <Q45��4�]�oHxή��� �W*w(C�G0���������c��U� ~�9c�8�T'�c���Kq��^Z8(�3�ZzI��]z���<���AXV�!����,M�+���lݦ�QMr���Fn��Gi���~l�/�r�.���Й�D��_���ߕ}��]�|��/�\f~첽<D�j��iӶ����8ʹ'�� >�3�~a��I@��\���q'���x��U)W݊a�j�I��fƱ���!��b��Kh)�~�dM����Ð��V����rX�R!�*k�N� ����I������@��X��ZD⹈~i��.���������{�������	j�C�KV8��U���)�1p(�K->S��U�cm̺ I�����`@Vgg��BR�/R0]���玕g�/^�o���径-�����4gN��q$����s����b"�r]u�3 ���B�S`�?s��̚���0mZ�Jڴr�8a�N)L�]�P|��N�mR1`ʠEt����G�s ���K�1�U�.X6���0�L��t�N�/0�9�urД�K]a<5��E�:�QXau�ݦ�]і�H�N���Ikdj_���U��0�o���'x��u�,I���3;����<���(Z�z�p�Fo̫�]yk�[�܏�]a��h�<�����g-��7`oa Ru����U\�ܤ��\�n�f�7�PV���@�r]N�`X�47g6^)��Rt���&�ýX��(1���''<=r����V���֧98����l��X�
bA��]��]S뤹���-��s�=��հV�LΌf]��
�!I�:��x�,@L|�ى�[��D��7t0��cӷh�9�U�K|���� ޽�ٯ���b���\;�c�ee�U=�d�mk��G��YYM��6K��f��\���jwMBr�(�[��nCuuӟ-뎺�:��%wcP��D}�Z�l0vH���w�&^fp�Q
n7 0Νw[��f]��hi�{q�ysΓ��hU�=wI�X��c�G3S�9Z)�)^���
#)�b`��?u@��0s�0�Xmfۧ�X�B���+h�I�h�@�v�4� ������M9	�:�n��ʏ�\j�ȡ�-��Bx�3,od	��)��ld�S��x�Q#�^�ɿ7lvs:9��)Nゝ�{:D��M�nK�QrǛk(�.��T����.�N��1�8��W:a�>B
�VV,W.ڑ���;i������	�e��bc��:��p���9��C�*�*o_K�8��S��7����t�{U��0��ޢ�+�����ĥuV̸S�K��w��$�i�{��%�y6��im>Q�A�­Z�,l���pA�ip.��I�t1��J<v,�۩5k���M��=���%Օl�m�G��,<�������G��Ք��CR�m���㏨_"��ٯx>��Y�@}��y�4���;�9+��u8�u���Kz0s�vM�	�5��Z/Y�nܕ�s�*j;��ݔ�e$X��t�2��
Y���΃��+$�a�]E-e v!7J9[���^����mm��Q�܌!���h�ܨ����ǖ�Mn�6����@���12��Zo]�p�`}.�i옑�bV7"��z��f�wevfE��F�YB��h�}"��\;$|��H�v����l��̗d�"�����ܭ�=2�Rf��w��ß�vDFv�/���NҗցnD�
�aZ�7q}X�E��#�����H��a1���d�ne��Ng���E��I�3g$��/�A��M���M�eQ�-��u�����o��������?Y��H�Ny�F�%:n&��E�a�swNA���N�i14S6���k8��������}����|q����L�c7 ��sj�# �3i�2�*�0�7M���*r���d���u�]|x��}?o�����ώ3�1]�$�3�5�l2J���2�����>ၸcQ\�L7
��pƫ&��	� Ͱ�*r͍��(��%���̍�٬2�-���g�T̊���f6�T��[&Uj�� ��߿V�\�s7]�-��"I��#1)����3,�h���*4�O��q�2b
�����EF`eY��a�Y�V�5&NFXm�m�NI�نf0EAUF�m��%Q��]�(��#����s�sw2��w
�ɲ1$�s0�0���3KH������Ȱ���,���"��j"7=�D�QE3�ƨl���>}-�Si�7���nQ8�����c�D�1�diF�!�d�^�OkL��6Z$n�d��.M�Jx9�t�X���qVĪ_.%��XbEv�,Y��bQܱ�ւ%��^�����-�c&�r"ZHBS!��@ș���L��l���(4\pH�3!�� �
T��
%�_?�LD����O����uapaH`P��}���6Q���8�s(��"�0aj1��H$������o�	Q���p@m��j��-úfS���"��)��E���Z.\]�7'���E�`��2a�\�@�Nz�H7?a�f��Utba�A�fr�InM/�����ڍ��JFw��8
�X5��z5�L
�σ��o�l��}�����g��j������OeR6�>D#:����F9����s8��v���&h4;��kUt6��M���m�M�s�Ie�+ڧ��w�؋.�O'��:�6��z�Q�4�}�"���>W�s+55��E�,��Z���}2�E-�j�aEx��层�e`�������NJs�hd�dO�E�^zG�;�I�]��Ѧi�ke�օB��g��3�yz0��4�J�;��v�v��xd�<9����g��<��_��
�x�͟��{>�l�U���ۣ��<��z<��C�Wlvfl��	�>#��^���21H�ZPz��&\�L=� xd�[Y��P�tσc��/F"�C	�؇l4�.�,�e��r��EE���&�z1��`���T�w���C���)X�cpY����+s-����\�'wzh7���n��@�}�����d�|Z��.ƖíL7��Z���g,t՛��
4Hs��dيG�丱�r�KW{Z\�W��/������
C+�	B��s�}��r�6�ܫ��a�m���K���K����eO���\g�3�eᦚ[�s�͖��hx���c<=���O�H��m�f���Pn�����"]�Lr˄噻�����-T�s����C1~��֪s�N/�
tG����
·�q�ͯ�7�K]WN���r�a�	m�ƕZa�^�����(7E�|oK%"��L��	:���A�Yxd�36v�]���v�� �ꖏ^nP��q��s����G�����������=��c������ r����g��Yz�#�b���M���{m[�*��m4	hbښ���[pm��]�qz�}b�-#�uV��L�w��`��v�C��������*���j���+���v=S�{a�G��܎��e7� ��~�8����2{R<��%N���X1�79-�kÒ:��[O�`Ge�@��F��)�oo��M�o��xbZ�ۙW7�a��H�\��=���$v�p�{yܩ���ѽDS�k�$~�QJ���-��L��{ ����1-5Ѽ��vO��L�#�a���Cte��b�^=��Jň�9���F@]ś����e�V�/z��&S1�֌*�f���ir;����}��q+JDYW���W2��s�y��xn��Le/s�7r�u�A+9��ϳ�	�/�]����wfCX�
�O#�s�9��o��_=���~��S�0�2�3���o x3�`�+�{J�>��v�T��#�D�������/����\]�}ꯃ[��\�C�_�?\��{�PbN"�]g�~���y��N��`Z2�=Ǹ�X�F,k�u	6�eN�z�Z����H���Z���s�FA�,����S�AM~D,Q9Eo�-�B�~���1��,�e> c�Nu�gӔ7���&9�T��1Bc��;6�p������/�c�������)6�A��g}�2��V _�[hg������r�9�|�D�%RZ�E4yTFXU��eMA���(a7�?�za�u��c�WϬ��72g!���;��>��!�H������ݦsݐ�,ٸ|/�����s��1����EK���
�����CJ��q�sb�����fȖ�1p��*u�I�����j
�C_�l���[��ږ�Io-����Z��t5�=�s�e�jU"j�m�_��� ��t�>�����^�#��֬�g��Wk���mD�{h��Ly켧�7#��S���-��a^݋e5���M�'�Lѝv/6fn�[�x�����X��L�%x����X��T�tnK��v(����$��V�s1���947ye	��K{�>[+�puc`���Z�	I�����4lZ�8.��L�Y/kNO�Jx�Un�ؘ%�g�w���d9`�	����0��>Ws��7j���k�4	3����t��)��"o�V%�7��r
��z�'Y��,�M��a�p���c`���u{ �f4b��}~��4��Q~��~ԧ���5��ه���$@j��N{CRB��2�!$��߄{�Ϟ1�#e31���sͺk���0�wT����5{;��pª�et(���{zSm�j�>,����Ҿ�?�1�� +�y/"�>��3�vR�۳y�*淲	/^�;�d��E,�3��Ŷ�6����������Y�ϟ��S��J��y/���1��^��P�5���h��;�
��`����[R��q@�d�Qvn,�E3�g�(�K+��SwUUݍ�7��c�^���2K{R-��L�dX.`��^�9���6�I�\�p�JJ��1�v��ИH�־��I�K�EFO'��[,�{y��'�>͋��W�b�6�5.`�䉚����=y�Q��,(z_�&CS�g�e�w_v���B+�{�n_��<Ou�(�ZQV��c>�O�<�L~�����dE �:G�E���2:��<BsĲ��ր���_�n�
J��D��Q�N �v���82 X���)t����_t�vFN7U��>��	 �'gv��������V7*h���r�71�쎳4<�ne����{����4����aa�q������i?4F6���y?u��) �-�!l"����i��Q�r�?(u/�� �=�Yw���]�J3�9�â�P��9ӛ�'g.u�[�����,�t��YC�Fc�@������~�DkH���B�_����{�"�̰ulzOSI3h�R�ڜTK+�)�z��4q��	WK�k׎ܑ b��~iw�ó�ׅ͘:���������?	�Ϲ��7ʭ�ݦ[���[a*Ɩ��@S:��eGkf�LC�vnhuT�_
,y6A�澤9�|Dݓ�ۜj�����v��=�a���؋b㕌{����ꢝ�ͦ�fD˞��hghVړ�8c�uW4��H����Ƽ��"�>9��K]�L?��0�^"����[f}^?�ȄƆ@�x�H/mm ����Ѻ���A��;�+�O�1I�(��e�9��h&us��t�B~h�,�b:��=�2��f�SN���ץᔀ(�oZ*Dh%W'�̺���z*1���p"6Rk�_mZ�lf��3QDZ�C<"A�D���!����~�ǀ`�F��[N��0 ,j��D��h���u�6�ӎf+9�zJCG���o���d~Q��q@��dʷ�,ء�O0�v�:ׂN� ���uC+;��+��x��u�z��y%v+%9�\�#%��N�������'�\���Vf�FD��M���|��?��BUHP�ϟ���~���Ҽ��n_3����z^za3��?��:%��JF[�b�7�w�Z�2�̘�����zN��e��#=P{���f�ngr�8���%���4��E�i�?'�d��273]�oU���A4���机5���C��"���r������(�����N(a�*<�k��uӈ:�M�>}�/C�H�1E˼�P�5�s���E��8�0�-d�Ug�J��m2���]�)y~��$mx7U@�7����|T��Qs	���A?Y.rb�'�=5��)�u�>��x�S�ZDL[-��m��h�������0�-�rȪh5��M5U�.a]#��V(`�D�E}���1<�X���~�b�=S�a�L�@�2�⑔ͯDĵ�j�|�B��V��`ɞ�N�� 	���(�5�P�c'�0��iCwt+v�C�x^0ix^��hfov�-~�(��n��hUS����pڢa�X܉�s��(
��K���J�F|�*tp�E���FC�v�R~�R)���z�:Y�H���>s�0{��o12Tg�-y���ޓ�zXrmM�ʄK����L�����i����*��y�<�HL��ҳ����Jq�����s/1�'K������\Q}ئ�[�P+��ڀ�ډ�����ˏQ�c�kf��Ubsv��#�z�tp���dY�P��? �Ra����(w���}�IN�1��xv���*��	��T/o��4���P��HU���7jT#�Mv�]�4h�&W��2}��l�!�1)֯l@�b�����H��H�7�Fh�-%�[��[(^&�a�΋�CsE<2i�.�P3��s�_�tFy����۰Y����L�=���^������䎡/���q�ϖ�KO��3�����w�H�k���;��j�O�HBA�[�����z�����[<1�n���4�]��0&��c�8�Q����0�Xrޘo�y6}u�g�NCۉf��l}U	a6u��>����y���7ε��6K��>�0;	8�="��Α���L���*� �$��������4f�!�[*�������N���q=��y��
��z&9�9�.0�1�^�fҶ�*tE����Y�0�I����>@v�GBOBFz5�0�f��Y��8ݬ�^B)���nM=^ͽ�~����U�q7�Ǎ9���">lw���>�v ��.��2FC���?��~KVxS�i.�Ϫ�$\Hv��k�We��:���Ew�{hFj�D����[����p�/�)pIP:�*�u��Y�Y��wz �0��޽r�R�YJ��O)�j#��0L�/�sӆѺݬY9ư.��1"P�a����1�k���a�s���P�������f���{z�4�3p�����w���	x��3-
5Hn~�\����ީ�Q�����!�q�-k��ߔT8��"=^���u~X����S�[�����+n��V�ͻ��S��3��ycGk�?�~�6�R&�j�aMCLC�T;hkk�����[������j�8ԁ�Ol:���F�&<��1I�z�f��b���z.�T���a:�~��5��l�h��c���8\Ir������'�e'ԣ˸�k׫]����y��������qi�>��~�~�i�2��5�Ֆ���َ>QeE���7�L��p�m��+�x��7������Ч�i<��i5��Mg=W�,_����kn��t9s�kQ��Z�׌]�n/͜
��
ߡ,阬$�=>i�8��w��K:��
�b���W�+a�]���q�Z�����`s=�L��.'��;�8|vvQ�`z��\���Wʻ��C�m��^?K�����pm�?s�8���'�74�܃e�X#=N���i-��s��y#�����/%�j�?r`,˩e�c�CCqͱ��Z�w(aPo�������A�e����Ʒg*ۖ��=W
0qF̥�S����� ��x\s3R2�-��k7�]Lh�D0k�����J�'*4��߆B~˃d@A	!>�P�1�ϫ��-��%�<��@Td��%%4�	�o� +��2ϬFO7�a*�X�FA�8	��#�[Axq��:s-ax�x��v�R�-�z�I����Mx���H3,�<E��i{ӯriYn���oN��ε3ط����`���j�?�/�Ƭ��Ȃ³��L3�Y� ��s�傍���ǽ�=�rvl5;�����Ԓc�Y��>�?�0ʯ�<����~�qQU8��~M�YU�j��}mw���H�%��j0��GLGG;�D{�]���Wj�ݕ�;�oYt¹�\��C�nAc��ۭ�As�Kh(;��"lh�8pmv�C~(�\*9[fִ�:v3�zqRE1��i�5�Vi�)d����|Տ�J֑>���z�m��mL�F{c�ͻ� ��>~�oCU(�\��)��0��Y�e��c{]�bʶ\J�`��[��0i�!����O6�(�h���&;��m�"��8�X�j��<�	�W!�I����{ژޮ�Z��y�Q�0(^4Rz�8�P.�e����rt�����;��!'�xoQ�_���C��u'�W���QB��ǰP�¼�Y7Mc�}$�/���3�vj�SM]�2���	#I��O*���_�7��:o����j�-�<tyХ�X7��Q���k/���zo�~^������^�oΟ�����c!Zf��eJV�EV�4�o���O]&'@SM�)M��k���ŵs>4IS���sY/t�h���o�e�&r5�5qΠ�!�)>5��@2�9�Ҡ;G�E��o������`�v�6!�m^�2��L��<6ϩNo��3�P�T�rG2�06�|TcsQ~v��y�i����]�VCo8��xL&"9��/�_`R%�U��`1��Tsr�t��\X��-����bm��--I5��b�ϛ�ZzD�~�����tE��QC9�9B"�?V Y �g�G�+�����.���pND;N�
�?����_G�<�[����^���}ݗ����7�̻�,�(R�[I��R�z��C�W{4t'i�����_��TG�>os>��I�mi��3��F)Cl[׷��*����~U��t
"m���0���ͺ9S�iylC��_m��]J[�qg�vl2e{wN��g�|H��|~�#/�1���Iz��z�ޝs����AҼ����m�;��bKu��t���x�hrt7��i�J�C������9����+0q��Y-Z3fђ�B��m��,i���tk]����A^�m����i�\ۼy��Q�hf����mgRU;w!x���9!j5R:m}�n�mpx��cŵ�f����u���s.��W�4[�یiS/L�y�^�Ĩ��5�O��v<�>�P�FK�f�����Q�ԁ=��}�ϐ|��	�=�@ZǤ�U�LD�"3n�������@3�nR&�PGC	�	�4����.���Ź�&���6��ӹ��WixB�fٓE`��n^�����'�ܙ���3�۾��AX,)��}:�_������S7M����"c*6��Hm�+�!����|��7��q?��*�I�����3+��p���T�V�-Zv�Lӂ��R�-���e�ݶQ�Y��U��Ҁ�J�Ac��"�8���e����趱vbm�;r�>ء�@����}��%�BNL�f�sjhJU�[s_>���d=��t���4�e(�x�Nm�����:�X�dhH�o.�Qm�g-���/�;��w������P����waL����Jܙ��=�2�<�Jz���.�[��<;�Yf$�60e���Ef��q:�("	5+#�N��^����7��un�u��9�
j������P�=#���nn[��ݞS�X����Sw�V�����V-N��y�
=Ͷ.���Ѵ�'2_m���G����
�l��$���:����{Z�肞�V�&�bE��i1N���ۮ�rS���yw���e�q�p��Ⱥ���yQi7�s�ب�"��K#�e��i���_�W�U��^I�x)�${E���#��:z�3%c`�Jep�dr�*�*b��p�����-uaxu���$�H��f�!��h�'P��ws�/n��M��x�X��x��Rļ8�"蓊KT¡Y���y�ѓIB��K/���5Y�I����i �⠩Ӭh�Y�O��袍����t��
dV��-�o#�ٱ]Y��v��報��i�3E�sS���������c{,puw�8.Dl*��h���N��˭U1!�:W*����+S��2�7�EǺ�>�� �̧�Qwc_hL��WՌw>0l��1%!��ُ��di�ڛ�Y,��k7B�q�'v���o.�aG7$��(�Eؙ���jeYQ���oj�Ɨ����/Ĳ�fJ�웪cp�,���v�q�A��	h�Z��Zk���+L�AY{���BB����9��Cw�[�ON��(����+_;�آ'�k���#�kH���gA%�@[
n��x�4��*�%�X�6q��+yӣ����oS)Q��_�~?���ęM���i�ET_s��,�L���(�s
�ȫq�������_o�����ώ3��ɢ��0+)*��,��3l�h�����(�<3*y�U<�u��}>�O�����>>3��g��X�MM�eSTď7�%)M��-�B-�,Xm��S�a�L㯏������}����3��<�)��2�c2��c��T�LD�ƪ32�*1�BZTs2�,��'*"�1�ޘ�z��DV1�%��dAQ�L�f�daQ14�[iUQnK��l�VTF�DQ5QEù������dDf9���o��f1ɡʐ��)6,�b�+3�O8�͌C�͹lY��U���e<�n%e���An&iL�9EI��De�XETQ�9����͘eM���F�e9E��9dcD��Y�e�VfVYE�cM9��ME%Q1鲠����*�d�(�2"� ��D�I�h�\s����zAǻ��;�2w#��+M�Εb��:Ne�E�]�,o�UU�ZG����C1�) �;����?�Y������G� ���V���	O�迁����>0��L����7�$EbC�L6��o��G���93����h��]S�(�C|�-\�Juoܧ9j�P�u�;��CKa� 6�s-��VP�Jr^XkR�f��nD����(	�N�\���uԻ(ZGE] Pg�}� 2Oآ����Sm�Un�_F8��ʠ~������y�1��R�.���c5��[�x�.�@����Q�G�PgP��鴬U�l�S�9�VNS�?���q[r2��;���is�9>d펳�	�/�3FRU�o�����0���K$sJ둅�k�1��!�:^(n�Nh���L!�ʅ�B]�vM=��U�)�����8an��5��z�3bV��R��_{��S(�`#�[��ki��d��+�5K��0m��+����+�K��Uoދv�E��$�d�Ǵ,h��|w�F0�B��Nz(�/���-�"Kc�Zܲ����C���2�N�'��>�c�N5k�4#�`�'���/��]�=�z'[����S?un~^�/dg'Bt�u�p��s���נ�&���y����	�</���r��V%�#ī$�#��Y��o/��*�@h��s\+�3zuۚ������t��˻�r��J/0���������¼�0�{�p3{�`8N`&I�\����[�f��~N,��PƯ��$ִ�h.Y��Z�6B���O)['�3�~��0��6\տ[��R1���P�0ރo@���@�1����	���}t�WF��n=��)}�����n~	��'���C�P	Y,�l�O����=[}Co�х��N�����=1Ngb�lE1��5�Ԙ�s�:�~�D�˄��x�I4���p���0S��=�ےe���f���7�u��ͪ'��!�Ȑ#!(�3M���T��B��ڭ`��_�uYf^��c���=D7g�k���;�*nJ�|s^��G��B"��=AA%�RK�Q�����\��dz��(�9��s�wReu�g,vN����%�3@�?9OJ�5�%�ܝ�����A�KT6��W�	��1����i?`��/�`���.�$v���*/�)t�{��;sdQ����9� �[H�%��9f�Ż�M
��1�	�b���<��n(���Y�����6��F���4_�[\������pef5�qI�?L�v9=GTT4N^�?;�����o)��N�����X���G�ߝ��ӷEQ:�`|*d����T�Nw{��9��Q�'12�Y��\H��?�3�s��(��̍���҃4K�u�KF���X�6�5I��]oG�,��R@Bn"B��њE<�_;���z�G�=���a�������D"� ]��R�~�s���YQ��蓊AE����,����DZ�.~%W�����	�1E���a�]6�ԿK0u�~�M a2��ci�l�����_v�,�N7�b�7X]:���O`����}�XS��(�}M02n.�5�T#���HD�W.���"�	pM)�䌖+<�y���mnf�c�͡�k�~��������oㄞ�DF'7�lY4+qO��������	Ia<����f�U��d�e��Q-+#F!>l`���ЅTqz�˽Bz�{N)�'�1�G�D�45�fK`i��g��)�K�ȃ�>Lia{�|����:on�S����o,\o�6#�j'�c��ҽ��>���	����FP�	�(������$�^yTG�� ��.��ݴa��mS�A�67e���r���Qt�f�#TX
-%�Ј�`EzT�q�?[l����-���\��f�ntZ�&$Kh2k�ː�1i�������j	H�6��D�П<:a���$5�0���&��ѣi=�2-?!U�,��5[u�,t]��"�s�n]�����$ڗh8��아�.o%�9��6���z�V����2X�w}�*�3$���c�͒,	�X���k;7��|K)��4;�\1��R�7���O`��6#{�B^]���yN���Cw�"�'*
��Q��&[�F�0:]��|���|���������c�0�2�y����5wq܈~7i[W����#L�W��i��dhZ�E�	����hr��z���c������hnum���]u�5�>�1��S7��4ف����*U[^�b�F �X�:wU�S���lރֹ�{�t˾k�ʙaL��%����_t7:[ ��Ig�:�0v�Z^�e��u�D�^t�{=ږNHp�E���y��i�B &Z����ab��������h�Ǹm)���Q����	T��ě��k���6Cό��w{jI���YnV�}*�hn���I���o��\oH~1��z�{b��ZQ�QR���	P�Ǡm�TJ��T�W]�����Z؍r�P���vۥ<ޛ���J�N����s#g!�*1���m��Y��9����Mb�<F��_�Hپ��QK#��;�B��Q>��Q�v8>L��Q���P@v����~��pLp,/t�yg���I|yh����9�}6z_}�PodKa�m���E���3Lx��cik���6�8����>;����Z���*��TP���x5����HkN����������t��EG�f��f�mZ3b��է�����'l� �?wRn'��G���7�G}�ϋu2��������o��l8fX�O/���ӄ,�T�T��:�Q\���yB�\��Y}��������Ha�w��o �3�lGX�h[|?Z���Y��§����[�p��Z�D�,*��z�}�z��0\E��*�2d
W��/�}9�6|`[cW�b��,L����Ƽ�Ț�9��2q����b���G���yJ���7����K�fl6�l�ن�W7@-��
�.�\�{��g���F�k�d�Sע-��6ϘP`����%Ai1m��}��.�L�(A���O���N�ĩ5���Q?x��ݱ!݈��p�1޼Q�e���(kq,���D�z����d#>��c>��j�����`�bzhΨf��x�θv�O��I_�6o�� ���n�m�0��ζZ���i��de��072�>߂[T�em
�d< ����;�X7��\Vuf���3ӂ�3SdU
C[�&|6Aۖp���=	�=�QI���E6�oXT�8�^DC��<���-{��y�T���mb#"m�4���8t�Z�O	��"����a��vv]��U�<`Y���2�͗��uzS?0�R���b����h�C4bS�^؁Θ�^���J�3{�V�bŞ��x�&Z���"�˵;d2l&���_T=j�Y��*�I��ke��E� mq�|M���)⸋�2��<G�$�ؽ=��^Ŋ��L�B����{�A��lyڷ�<]����ˬ
���X�zba�V9<�u�K��n��@�|G�|A�|�	ii)nz>����y�}>��܈o��/���Juϒ�0�O̚}]��|�wL-~��_�mB8�������
:9�7z~��l�ݣ��[a���翸߆Кy�Z�qI�H���}Uՠ4�l<3�o[q8ɬd�Y�3�X�D߯�� �X_�缨E<�yR�]�0���빶{aAu,�)^9���o���ٳ�zq�ƭ}>Ў-��,�6�[3�3{�
�,Wo���䢆=��T+�\�\v�5��&���T9j �8`����
���Aȝ���g�|�<�F����-��2� �(f��}��I���'
��=�Ug�\�l�����d�|#�C�\V������w��j����9�S����搳��A�8㝤86�G2񈦂��.�wd3ap��,�v{��/�U��(P�őߤ77�秶�O����,��q��T��:k�_O��t��z@	�TUhY�jg;�<��_�N�Ev�~c����Ժ.�r��/�]�k#̓@�^��ŕ�񒺌��9��2��a۲�,�Yז�Y�}KM�|��y5�9�X�	�5����� U�!ϲ��J�eϠ��$�fⵛ*/�k�we�t�n9c3�������Y��f�v�r�:�-�����
f���1�pa�1�]���9͏���z7�'��� �CN$�S�v�r`}:і�oL"�i�E�6(1���m������5Y1��X�*��_�����&�$�^��g;��E�,;�X��s��9��x�f3��6/��v5'#f�.���]����vF�5��A�wd�)r̠
�nm~��S�*|�U0��o�Cìƹ�;q�!���@;u�Ԅ1[}�a����Րx/����sa���jlFu���#O��Ž�����7Cw�g2b=]��:h���vZ��.y�e��RH7�����CCe�Rf�P}1�3fo?=T�ԖQn��j?�K+�H�W�+�t�^�ƥ�Q�6�B����oL�����6�aiY��hx��Y��v������Ԥ��(��ⷳ����͟>˾8^���o���"oT�psb�Q���Å�p�P�����
gU�T ��7�j�g)��@l�?]��ⴂ_���*1��K�)��oHĕ�g���i��+�P�8i�I�(C-ض�r�{|��j�����7�.Q������5~j��jNM^�S��F�
��~��Q��bk�V[�x&���T7�I�J�F�e[A�D�25��rj}�V�?Uz�Q�xc��vV�Sd�;����B������kl�� @�:�@�2�w8h��Ʉ��mn=Vn��C��s"������9^y��Q{7�e��˵�����`��4u0�~�|��DS�	������:��V:�۠��N�eq�-������f��Y 'Ȋ�>��^��D{AP!��\�̜֜�8"&Jr�n�(��Q�?P<]�q���m�H� %6����B~�1��ӓH�Sj��&�m����+kԘ;ml騹Y1�nei�:.�NP��}7�L0�Ъ��ⳣOc�d�{���(�.A�S�`:J�@�"SEd&�'(V:��l�����[ܢ �)�)����ڄ8����mx�z�m̆.ꉶ#�t�l�ޱm�ܛsF-��#�MU��(�hw��(��Ҹn��!�{t��U�M
�:79�k"�f��-�Ʃ�{��A,�`S���up�+�jk�v&eo�{�����>cNt1W�#ݛ&�<�L(���ؕ[uZ�m	��Ơ\[L�{cKq�dmĪ����"x�˕��!6��`�9�&�?(\�}�gy���6�Y0�T|d$��at�H3\?y�۬���8�7�rgΌ��3� ;®�sE�,Q����f��mɫE+��0%��ܰq�����ȁ�s���PF�| �t��o�tꜚ}Lۧ���N�]l�j��1���j55���7�®n�;Wu:��w3x�k�f��(��/�=�1	��N�kȷ�S�����c��8�����\���_d��e	��ٜ^c�u,ld@$��Wj��#o�޺���Ca~��Z7?��t8ўuwm��c�:��kP�=�����V̀��B|�>�
��6�ߌ���y�7F�U%%$'s
��%�ls9�F��Rzu�j�|�]�5>�0�З��o]��h�s�k�d��f8g��w?���(����{Ӿ"�;�.T���HZ�__R��0{���GD�t�"�>�U0����>6⁸����rz�'Ɔ�E�A����v�w�\0�~�U��Z��Zm�h�R��.7�V;6Q�ey��`7@-��H��Mˌ�2
e�wS*c"�v<v�w�r��%�}���$��YV��mQ��s�qlz�}�v����hrtٻ��ɋ]-���53e��p��7P^�;6�xT�[c�ߕJTC�H�����%��D����M��gi���G{'��M��>)gZ���O�<�x��8��V4����.��o�cȌ��'�s5��-���:
�I�^��Sg�v,�g�_7��*�~��,��h�e�^&V���k�[Y��Գ�r���JӇ3:��SK7��[��gžS,J��ԓJT(_WR����Y:R�t]h��1����^38U�2�|?�#ow���9E����t�(�M׉o3� F�Sp�������,nF��昄_SnÛS�+\U� ׹�c׻�2籈ͧ86�����������s\�4?4�<�W-��뵃��΍mg]���J1��;�7B���Bbr���7��i�K��f��B�9Ge��҃=������d�W��C6%�`r1`�'��t��f�ڌ3Q����ۑ��r��s���FO?��t^0Zg����wO$����v��0|������g��.p.�Bs��0����:��.xd�w$N�>K��F5C�T�
���乓�_Nk�TMA.�d�ǵcE0���!�4:�����VS���a-�c�Zm��]t^��:kށ:��^�dy�99��<�r�|�a��f��s|���r���R�B^�O���-R�O�N5'�A���S�b����kK�@��q�y�~K�B�Cy���6��#'&����r!ٴ7S�S��"��Uǉ�#uތ�i��o����mt�	��t���9��A9��9��]
cx��X�*�y�R��r�y��Y�b�a׸'W=gGT��l�%�P�܍ז���dٺf6��b��e�4q���U�n�:�_$p�C����ݷ�h��õ\��Pv���􆞍0I�b��-���ǂb�VT�Q�!���I�KW�!��ъc8�F�ʹBNv�[㭧�1-#��-�َ>ŵ�85����#��p��8����zw���԰�U�GV��XQ��݇�7,F�Ѧ`���_�X��2=�Y�TYb�}��r�e�J8(i�9��רI׶x�c�x,���H2��h_C�L$/7x�#ƛ��W���z���Z�6v�S�{���e�/�c�:hք1�y�� �̳ܫ�ցَ��;��EE�f�=��Oz^�]o,7a�s{�lTբv�x�w��չl.Ѣ*��U*��1�rg��U�}�!�c.b�n��U��t��4���v����<V ���ȁn�	i��=��������d�вku��jN�({c�uk�z��rIh4o���|�l�W��ȭa���a8�����G�3��k�>��67v[f��3L�!n#�ú�T:��D��a;������N]̗"ܓdcn�1�j��o��N��B����};�U�Y�cʹ�����P��*����(3����un�`�?��M�Ka<c��ה���4�<H��+(]e�~�lqV+�I���yҎ���h�].�s!���O]��<���Դ��J�����@bkd�n���dS���$�X�/���ݴ��77{�΃WV&�[/kTqa�-4;ۙ+��6S�0ɤ���GP:v��F6�ut7q�����e�N�݈p���c6���d��p&��p��)�BRw�h������Y9�.u��5y��-]�!w@�Vhh�4<w��p
��˔s0E� RHK�2d�gw��3rL֞�8(�@�y4�S0G�R�ND�+�����o-D�J#5�Y�,I���;;jw�d(�U�n�8\ڦ+���a���'N���f�Ϯ���y�]�
0-�x������RϞ�C|x�p�8:�!vS�Am��|��9�Yc���j;{��ff*����O�3[^U��0j4V�A�-vn.�b�)�Jw^L���nWJ�s���ۺPZ�W�(c'G�k�r�s��<ζ��a3�u�h︑Kp�8m5��wn�z#mF��C�O�[2�n�$�I���3��&�"rl�;�,�լ��7{�k�l��C��f ��+��`�Y�N���^p48ZɊ%�O�N��G�i��V7��H�Z�N�4����S;n��IAqd_��16fF��TFa�C��Vn�2���556e�A8����}>�O���|�>>��w��L2�+(*����l���fS�1����bj�fFFUf9�����2��q�Ǐ<~�������ϧ�|���*i������"��X@ELN�VM�i�EA��cRm����E�㯏<x�}?���3�힝�
���1�!�(����b��*��1�B¢݌50�2Ȫ*���jp2�-�,(�r�,Z���7Mk,���*�cs�i��PO3���3**����"��fA|�b�a��0��
�Ȫ��l�3+c+,"��I�3 �b�2�q��̊��b30+g"���p��&()�K�9'�e�5^�LUz��`��5��j����Ɗ"�**rp�,�((�(��"��3ʛ,
��r����#��b��b ������""�"(�h��"�c,�)�h���į[�QTa`UVaf$ES��g>�ې��!�AL3Q��b2P�Ip��7!G'�/u#sq��C�ˋ0P�yЪ3���6�N�[�Jp��8�˳
�����'`R.A�� 9�a6,K*�����Xq$ȥ>�A�0�-���I#aD`H����0Z��ʎH�%����\L�!m�? آY��0��3请�MCdb��&����6~*(џ118�$
�J�'�!����V�{�	����ϋ2c�T��>�M���)�{���m�lW]��:��0�;"������[�0w�xכ��*���O}��?ϸ�P�+�N��s��w�
�j����L��;o9f�l8Dc1U!�q��M�o�:1��$�Kw�ry99�V�	Q���M��]p:g�z���pՎXît���f�'��`,�}Sۏ�>^�����GM7�%y��s ���[��P�N��P��c���n��D�j�P�}^�n�^������ C����֬�K?�P؃>��3�?���-T����!�54��Ly���Ŕ7+9�29���b|C�/�Y�,ˑۚ���������63pxrR�b�2:D�)Lf�F�,�[�=�L�^��r�B���`�9YN���-�r�m�g $?�<��>�	�u��w�a(�����VӈG���^Yc��ة�ؼ��E�_����}C��O���>6Rg���N��X�C�^�aC�q{�)�)�H���h��֬��߆~|��k�����C�"{�!�F�6z�1ON��uP��<����˯V�4��]c������bZda�B�w=n�Ǘ9��|~�n�{���	w1�hARv��AL��W�u���e�V�侦�2��5��m^���dr��gMŘ�����$�`�>��`0�_S�O):�1�=�c�z�qq^&�s	,���a�鵹��u?�^ճ���1�ˬC�n���8����.}hЪ�<\W�l�zGs�J�8員Us�-Z�G3�2�����ݤ0���ۘ�&�d�S<��T��g�"šn�ەX��8ө�u����L�f� �Xj끷��r�Պ�����͹~2L��-�Kܹ�`����6ϯp�����vPE��(��s�@eVwWv�P��Rd^Wa�W��g�@���%�9��6Kt���xҲ���y���N
'f��q��ob��q�V�=1����4���8�:�|w��v���G�4k�s��k����r���q��T�Y�i0�_��T�]�Xұ��AU�6q莣.�KwK�C)��/�7U�T�	�ø��lk
a�|�Vp;�E�n�@��fs5������Ԁ�5?q�WНV�"�!�T�W����T�M%��"����j�9��5��E$��ң7ێ�o�ˮ�S�@�b��QU��A�zZYω{�n����w0�H�Y�]��httœS_\�n�!�t��lؓ;uJ�������6H���s��͎��kh�۹���At4z�ù�nBXL��y�3�:!���b���+))J�NI7j�S�L^2���S�l��e��~�$;��Z�^�}��~���J����_W>flS����M�a�����_�#H�ݰE���g�<�=�m�[z��Z����uls��=�Y���L?�d����@�q�J�\����϶8n[�]���^|J�l���rg��pUmv�츋���"�7Âz@�[�1�)Dy��Y��x&�T�7^dlJ�L��rçVҽ�66C��u�}�<�vҍ��Rڴ��od�9rY�y�MS�N����y�!��<�-W^b�ꎃ�U�txQ���z����ƧAƲ,�j�ﮞ]+�qn���<�n��u,�J7z`,2͓_����P��^��<a`Տh�^���Z�Z���/Y88oS�.�_��"z��k��[���q��mG��bp�N�RU�Z�/n9��aMMl�S����]}�1�z��F�>����;�ەx�g$K\��u�Y�Ǿ�G��<�9��׃<a�hd�{���=��=RMKT��63�5�*O�Q�m=��u�e��G��U�.$<oKZS���do�e�Ɔ*�6����pL���ʜ��ʸ�_nl��+���C}��~�B�Q\������*����6��������n�]�3S�FO��l�g�q��36K��b���6�nD��(s��0F��0��r���4eenq+�Yq��G�z�+��嘭�3	�quѩ-�2�1dQ�<�絼�ՙ9W�_XYrU?R�ì4 ��qu��f�i�����I����.�n����yc*�D��i�#��2�u��E�ȟm؜�� �D�/�S--ڋ7S��գ\cf�f1��'��i�=՘#�D�����h�Kf�"�@��v��<9uv����3�{�Β6��Q�u�"�;gK��=1	�Ь�����B�]��]b�oz�5��A�.ձ�dS���wmvd��7�7en�9{�9V�0*��� m��kl=��r�*�j.����]�v���!k�gwWN�y���fN[�
�j��`���-���V���:�W�%�"
D\Zw�YU[��	�,Ki�PbC���%A$33�fj>ߍLȫ�=t�%��۔�Y:0X���ﰉ�]��K�ȭ]Qv�N�Ŋ�	^����1���ݏ�]�P׵�'}��اu<T�|5FW��k���m&EʇØUcoi�<�q��D)�q�i�NY����$��0�N#ʺ�|���g8��MA8��2~���M����/�*�hP��2@<��	_�0��;���+�w�δ����e�}�@q�f{�L.�mR\���fM�;j�.�U�t7snz^�M�fj@ϸ�
��֦ա�`5��H�@��E^=o���׋T�q�V��
y��7���s��Rs7��!��;;3:վ��"���`�K+����Q:R�l"<��U��_&\���ޏ����$U�m��:PbR��M9*�������J=��wd�̱S(�в�G27eV�ف9�F�j̊��g/>ϵ�PJ�@_�,C�4�k��deQ��ͳ���tQ����yThj�J�ӈ�c��*g	w*Ry2A��+��T�ld�h��f�K���3��j^�N�(K]t���0o�����"کr���c���>k�ڸ�\�Ұ�?'�Q�Yt��϶0f���z�+[��32��I�mj̉��K[���T%ӄ[ÈV�ۖ���w�%��-Y��V�[���t#��(��1��839sN�����GWu>�F`��x9�`�"�NO5�¤wQ�`��[�˭9�O����-�60��ܝn���}oz���d�
:g���I�(���-ʃ
f�dĭ��`����nX��m�0��ˮ{bљ�\o)hwmL΅��1Ǣ�0�-�U.L@�vf{>�W�wk��ۭ����@�o�W��ݝOE8�����GL��x�wdo+�ǘ1�o3��KbN.��R:SMn��CP�уq����v��q�ɂ�`?o6,���L�1����{�g;7��FRZ7�:3�6[��h�ؔl�����lN�Cۖ��F���n�C͵�|x�wё��Q�4�"����8�:���ױz{��}��W
���oYw�������1G��k�Z�Z&�N�z�U�{��C�o	lE8i�v+N�[���׃�m.�g-�L/3检����B���������=�2o��7�=S�dX�v�|�9Ü摶0#^����x��ڇ�fL��ǆ���l�6�Hȉ�t/��϶g���D�B�ǻ�fY:��{ܽc�բ�����˟k'���W��al��v�TD\,�x��tQ����rhiƳ.�6Z�]ߛ�O��.1W�Z�a�1v�T�VK��
a� 3�����s�Y���6����fN+w�e����zgג6��,3C�N�/��ɬ��<�����Im�+�Y��Lz���x�d3�����C2�f��ݜ���eh�p�����l�$���&v�wy;TD4g"i��w��f�8���H	ϣ�,^���Էݡ��2�m.�2z�.R0S��w�Y����t��b�u�tN��p�˩�����yS:~̋!�A8��r3sg�nͽ��Bз�cb�	�~ukN���w�J���Q� �m�A�G��:�+ul�]�����;ҥ̱��-������[��f줰$	����y�]�*��6�݃]S�\�Or%K_\�{��|�a4Y��F�:˾Γ�TI���qaBӵw�xp�Y{�w�~ �r�w��Gua�+�V㳪qފ���_��W�A���[�n3����yǅ�ϔ��2�r6���*y'x������xb�u׃.~�c��~Y:�}X��wF�h�^��TY|Y>l*����^��q�8�r}���6���١S����0G����'g�ґ�-V��M��+���f\1��H�ʙ��Og���PkÙ�b?����W��w�E�6���A�VW�\�MFP��ڀ��Y���#7�&��W�=��Qrg���S���yEo;�d�����sиb獆���_+�K�Z��1�/s�;�*a	�"�H&*q[)�6����ӱR%K��$��hf7s��z��j*t��{C�u��M�j��ڀmI��9�8Y�睚Q����٘X� ϓ��[�ʯ�-�,���Y����<�����K6F�J��J3��cy�6�b�Q�����S�#��7b��]I��k�g%L:퉷�2�kݮ�t����H^'�dݮ꽽ئ���;��24C���W�_L~�(��ڞ��j��n����楷���j7�M����D���?}1�@,I��k|6�+h:���*(��07���7��C*����*p-}��GBY^.�xi� �opg�g�̑�z���[A,|���^�Qr��VTE-�j�����=3-=m86V�3k����sau]F�)��0�H�7��:�̪��3�LN�w/'&�}�5�΀E{�q���~ܐ
����"�t�u�QvIQS-��v�	f����F*��z}�T�����5d��CFz���mn���C��r۸أ�)�R"�OV(>�]7õ�I̳ݠ�V�1��[:�A�O=P��dñޘ��*žYѦ��3������Q�]N�9ûo��y�,v ��0;��"�[��ړ�i��?L?vk��:���_4�?U�@�@���B����{��p��Fy\O _>슩��^z�_V�7Y�Y�R���N����a�ǃ=,�Ce��<H����?įʹm�����eo
�E�g�&��(�F��)MK��+��J�[
�5�\��4���m��qL�e�=�l_+hq��P�]&�]�:T�o��}��63��ع.�.+ǝ����������=�t�Ys+߾ld㙨��(YT#M:�M�C��s������칒n��p;xD���i�m\�͛�I�l��ޣ���}"����f�U��ʧ�[��A-V0O�3:R����(�fi�s�:����Y1�/ǜ��4��X�`����%��5�i0��S!wj��|�M� ��4�Dr�=<FV@�`Y̜.��/lv_�F�x�t�I)a�0FL�L����gz޺�uW�v2��i�wlg[��-�i�������q��K=E0�����J��[�	@d����-��t�-�ƚ%�mf4�^kS|�{�+��"��<�tQ�~�)=yn�G�\�ps��]a�{���t3�:��zFB�F.�ut�T�{��=}Z��u�⽙�rg��5ă�(��O��.��F;Wx돽b�\S��CL۰�zm*��|�"]F^N�B�c@U�W��%-S���:Wj��b���yi
4��[�l����x�ֺŦ�:ic�0����ʉ�{:�J��f�ޝ�N����դ���U� }����Lk5`�����#���f�q7�0�b�Z�7ki�\�ʠ�����5���fͰ[ُ]��N�]��^�[׷jG��W1�or0���V4\@֭�V���s�'-������j�]���2�NAz8#���\�����J��c�HA��� �r6����(�
D�j_j��Ŭ���d�vͽ5"g�쾙��c�B��L	�0>V����k�;��{Q������Ai��#�����un��u�Ѵ�5���Ky�C{6D��|��B���,�Ysh7�������Nȯ��P�ݍ���S�W�>;ֺ;���P�4V5�l=�@��G[�d���A"a���`̖����Nʽ����]GX����2Pu��me�0�|4���j���!���؋[��7�
jL�;��Y\Ol8*�h&��n���NɴJ�Z�g-�i�:�=����w����x+dr��Z��."хy�D�3�k �gf� ubs_;x#��v$��@�8hhm�z�<����a�B�j�i�-�S��8���p7����
�iiɹm��D[��4����}�R�O�f��76�5��l2i�C{tE�k�������7�ڤGb�f���K�mG������9[����;��xv&kq�}�N�ҝ@��_j[)�ݩb�#��F�7�c��T�f99�P��Nՙ}�=]2�K��<�M�\]���.�J]���R�+,�{�OvD�pv�S�Bv^Fܜ�m]���*o|h��rt�N�#\0�@e#� v|iaIUҹ1��|+B0�5[�5t������!w���B����:sL�J��أn��B�2�eM��k��h��C���w;cp���S��ݣfg6�:�̦�^��g2��{��a�1a�i��\NF�Z'�i^��;�Ѵ%w� �G7o6lW� ?���L^wp�m�ʒi�8����1�9}�-�`����)CB^Ҭr�;'[��e(�U��E��N\X�*���c�#���sk��Z�`Uڢ����g��b�).�dhe>ʺ�{�~\*+2v�y]N�����:��TYJ�u0��;�[Վ����\��X�����*E:�t왵�u�Q�17�ꔄ����|�Á��z^%B0���u��Ƹ[p�GD��IΪ]f^V��Z��N�TK:gN;fŮ��1m�	-.9��w}H1xl+�d���:���A�9j��5>�Cf�\��5<�F'&(⻕4E��ѷ7��8����v�$�S��Q�G�MTLL{�&")�k�bAPDIdQQIe�QI8��Ǐ</�������g��ET�PSy�ndђe���U3DEY��TQPfe�3���<x����>>3>>��;�ST�-U8�ULVf��Udd�Uf`P�`{pr���EQ����<x����=|f|}3��DT��E^f��S1CCM�����k2Ƞ��$("j���Ă��9��efaEMe�َEAD���%�Lfb�IMT�TAAD�MdQFf9�SED4a�Y�e�M6LfLIAf9%86YeUK�ƶX��"��2�30��������b���*����Ȫi��9:N�V�b��
Y�aYW\͓$������B �+*�j��bj��"h����4�f49P�MD9�Yd�c$��eɉ�iL�=|�C���=�ݭ�܆�fc��j���.�	�=�q��k[1ge�w��z�-����Jt�G�$/��R��1��bj3s�0��`Fly���,��z-�u;�����u�5�i��<�₏�JAƫ��r���4��e��y�'|�4a���Y9�+GmV�����ڰo�g�sB��Ű덖G�B��q��s�o�w�&H��UX��9���Pfl< ���^*����s�ϔd�tc�_����o�fh����2��n����b��g��r}�X�)�y�
����3������߱�H����K�&���q�m�������hG�a�y�8a��i�n�t�l���R�����J�f�������D�����yF�	s��u�,'�Q^Սh�E��3��p�H{����p��6������ψ������,�mm�W���m3n��zf�.����6�ש���M[�=��(Y��zr|��+�*�g��Av�iu����k���,��h�q^���s����6�r��V�SU�-N�x -���4PrMc�+�O�Ц$E7���\�*�B���ɬd�#\j��r�AY�Ɏ���-7�9H�m�vUb�2֙2�s'��#���������P����a����)���P*��	VMu[�1������2�܌U�W��P�4r��,����Iuo��Hj�k�div}}��j��������� 3��W��$g[��=6)̮��k��4w0[��5B3���{s�V9�n;��+[�s[����9���8�m�^�>#�z�k�Nٯ_\��*p]ʭӀ���bl�؟8�5�t?s޵��6�纓�V��V	����ݧ9w�Gf���9�v ���y=����:�3��ޥ��,�P���j��C��l��K�mx��%��s!��v�tN�M�玉�G='�-�;r�!����3T�h���6q�ՊջT>�ܻ���9@y����Pq��f�.��9C`?��w�YUfCp���pԿ�=�Ahϋӭv��b��BP�괖��r���������l�g��;�S7�+!JWT�ٹ�U�A:�Ѐ�Y����c�jf�"A�^`n��8��Y����������E�1g°���ަOfn��y�>@�IӷFQ�6���{M�A;���@
��� ̘���Wr<�sh�C��{>�^Û}�-s?�|��ySv�M�[	R���X�ܪ�v�(F��4�$
mْ|��$Ӛ����$��:�op�����[�R��1@x�F^�;d4u���Ɣsdq��5*�V@�����$�N+��l�!�cݼ\�lv���|:2�
���dU�nT�IUZxY���N�-��X]���8�v�[mX�=i�2��"[�<�O�oO��e{R��&���d(tt�ｼ���|5b�H�n�zf���Я�{%0�7B[��3Fa޹��0�]W��7�v��#���sjG��
�!nz�W	]:4	�L�f]E��=��hd_rc+v�)���ݍ����lxK\�0L�t��U�mPz%_H���c��݃�v��۷'��-�b�2��	���^Z'r1>�]�d9A��Cw��^��9]��)%�I~P��'q�����i��P�ne�m�"
3�Оz�3�VWf��;�^'�qD]�z|��ok�T�#K�CF �t0m��6��)�w�
�HZf�<sf+n8��jm�u�Uz�`ճ��W\�n4�8�a�O�,}�e�f��/�b*�}�JIpu�n�f�mn�WIbs_ed_<]�㬵�qc�4�4O��{�}�u�N����$��ng]򥽧&-Hy�fs�J�8�}�����fl�c��L6[��6&
��r3�PW�Q5*";it\摽��v�s&|<�g��Hqg��"x0mǡ ���B.0�*%�OL��2����kP:�|�P����\�i9��KB�n�WsD�*�l��={���oyX���+P�#e��Ii]�au��l��%MWw{-�����*mu�Y��~���~�q5̊[fz3�>_��ߪ|��}�lI^!l�'��-�wlO�¤��p��s�+2ԡ��"vi�_��8�tR*{��R�yP��uCw����G>�3��f��]V�m+��N��]-wڸ~7(�Gi� T!Z��xt\�׵�ps2�-��8�]���=^��1�h�PzL�}��4/XT�e�ެ����S��-�Of�B���i��[cT������Mu`��h����@ ����V�۾�9W[�ګ���L�7�a�[z4S��;���/�W]B�\���y�$��w677/�����������X_{�
�� ��}��hi��`��#�B�OE^��ie��Ev�ck;�'�wV%y�˚OwQ=`��v�r9�S�n0N��f�S��kFɛ�/���
a�GzE��RQ]�Gu-V$��2�U�.3�����U�HwZ�F��!��:�>ק��&�q�EpC*�g��C3-�u�\�mlM #("]Vz�,�"q	�f�|��hN�s��D �Y����f�Cd���od�C��s�{Ly����q�G��>�qhc�OӺ�H䱃���3=]"�϶L>]��[Ƴ��eA�p�Z[��Sw!D\	�5|�\�p�v��6X_�������5��o����{��>��˧�;h~�]�,�>��y�@XMNB�`���h�vc����b��&�i�;&1����˵�s�f�<�p��t�)��_��q����p{��#6�i<��k;H4(��_X�^�6=��Y�#�P;��k������{\�����2�(��wT�,��,��H �A"��~<-��V����]+F����v�h5�c̫];_�ݺ�йjV�R����|�꾺�.�~myz"�	]����a��p<�4Q�ޙD��f�B:���_���z�vx��:��G�.�%SoJb�{v����!�D��s4��$;WL DDy���`c�v F�0��6����f-w�q�����Mm6�;��W�n��L��Ji�R��S�{ht%�_�+Y-�0ݪfBU-���YR{�v�'u�Kq��\v������$S�V� �m���]g-S����m۰�c�w�*���5�T���@�/�J~s�}??R����޷���������������G�����е��מ���U�=].��sG8�Ӛ��Σ���ϡ���{T�v ��'.�:ۓ����Ț��J�I��0n�Xe�]{Sf��2��Y�/�����n��3��Jsj�O���H'o��}���a'�!�e�q0�r��~���9��Nz��t�"��!8�߬��sͱ�7a�#:����	(��'��-��s+����|��] ��jO��\!��w�;��ـ����Z�Wj�mM��vT���c�-�
+�{.�"ޢ���H~��'j�A�ۋ��_�E�2�8�i&�f|�e�T���$�C����[�(}�z���>e�9f��u���d�St�p��=�_y[�!���|7�^�L���y�w�9s�.����?Ӽ�?P[0C����2�U����]�X�aT�k3j��w'T��a������'�Q���{�o��z��"�{��<����9<�*�nz�M٥`����Sӵ�T�E�e,�ߖ\�}h���[r����U*�dV�B(d�b�m��V}��}��RZs�C��}��Mu	]��_x+t�'Ժ�\���o91�4�Ef��w�d��i��Oo�>�)�\����S]�mM�w��vۮ�k;w�Ͷ�C��%o�l�Cj��&"��=~���d6Vk"*��t�Ǻ��yy�\�+�'v�����B�>��j]��h�X���l͘���˷��\w��{�� �#&�oc���Y�n��Z����X���^�B����oGי����Eq��w��P�u�T�*�ɲ�;�%�V�r��\��������G�������l�1�Ū���lE�c+v�؝��F�`lq	kl*�y[�ԍ��v�đ/��Z�*�hV�-��1r��܂���x�u��SҪMn��f��LOsDC�Lv���P}��9Kh%]���Tvr�sq���Z�w6�!��ٗ��nT��(О�1�U�����T�p�`�3�k���+�ۦ�~�Ԁ��0�7&fb%��j9	���*hڑ+��բ���;�?O{L���G�n<*��!���o���W��/+��7��$�o�=���oc�6�2^C�w�������ܕ��jmBn��[&+hW`�^�7�{�MP������̶�w᭗��g?vI�y�q���@<[ym��f[@�}��:b
�i���h�\��[�<j�6�玀�Zѱ]t.��W��u�^o)�ڇy�d�����گY�`����VSKX_.�}s1�[�GSKW���g�Peın�!lp���?ag��x��>��\���W�5�7Z(���s����2n��F�k��.�u
��Z��,%�.Z(@��=�u�+��~��g�y��P�����u��)b���fc;�'���;z�"�V��yI��T�u��8�-~�k��g�,�_�{$"�Y���e.ؖ����y�۠�է���j�|U�P�.2{5�Hk��n5D�Qw�x��/T׉����{��5��RF���Z��_*z�*���5���|!�Jyh���s�hɭ��n���^�#��!�*�4�v m�M�an��V�׃w-OA5��4��Ƭ-�^����bIm��	P7k����[�3�u-��.�ˡ�t^�����qrcV�d�Fr˗���b�-��K��o󛱛[�4�
�>��`�`�X]�=1���h�]
���=j�b�M�Twf�����kV嗀�}�m��1����U�w�EKoS�O`��俼��O�K܃r�ې7������V���_��G�����5-ǫo�2�Q�y�:
�q�9]CIɦ��ްxZ=��7�b��'�ʲk�Ɓ���wP����p4?��&f�ꓘ�����Ns����0�,w�U,ue�"�;WǮEqn�=�k{��G���<5���Ɗ��
�_Uo˷����4MAP5)�����$
�7ޯ�����h��Ygb�߇d���k�	-��ȁ��Y:3k�ey��}��'QȗA57f��홺�9���g��ֈp��#�mӠ�D1T��.���v��q�D=N�����4f�im��6�=��s䟳�k_��U6��t'��[R�8��n�#d"��x�#�%���[�4�-��g��obWu��CZ����/=���Kkĭ���@l�����w3=߷狾��'�2�D+Y+�EY�u>�����Z��*�!��1'�@�gv��^�Y�ɞTYoHu�$�����^g��\�{�Mr�/x�P�5 �+�O����ƥ�f���^�#���R�vy��� �;5DI�{}��A�{�Qa�੗�[^�ŏ�yݽ�Gُ��|&�2]��K��$��sa���Έ\��t��8��\ؚb��$t�az�Y��su8�ﻇur�
#F�O�ce�-b�2`�'S��}�-��0�ɋf��9"lIG�����9|�;�Uim�m����8Xu��ָ�B��Eι�n��4�7F�K��ל<=��u>9�q��oL4��8�tuTFڠ��ާ����lQ��ۡ��6���V�-_A|�Kxȥ]Nw#����w��M$�n�����>�Q���{�m��C�hpA�6����f�`ժ���Օ{�4d��L�͍�����K��J�:�WE�W��[_-��ܷS���X@#�y�}tCˇP�X���!�n\N�+9e��� � �o��u[�f�7y�.mX,]�-�t&
�\ݻ{�L���yµ����CL��ٛ��f��1�Wd��r��e�ze&93"���3(���J-V^.�{���E��ι}\�/D��nʴ����c΄	��9���S�{�nf�B����(T�P��"z� `��j^�=���+��&n9�,E��J#�������ց�n�}�;�>g[綇j�һϮ��^�-�2���� ��r�uϥJ��yu��@H0Z���-��	��e��Փ+e)�g����ݹ��[��>��:�e���\nS��#@e˱uՋNo˨�L[�9&��q�("폇b�7P2�Q���^C�չ*�k�d
n���4�hUi�s��!v6_Ҁ�t	'C����0��H�d�@��5A9��h��i֗a%�t��D�nU�}��!ٸ\��ELD�D�^)%�/�0��q����t�rH���G;ʾ,�A�	ayɤ�J�i��7Wy�vl"�T�2�Π�H�ە�6O`�l�x+y>�ZUJ*�CU����=�����͘ڋo��P����f�RlL���+�c�2aTXF^�L����Zf(h4��ƗAU�]|.�ӫ�jf9_u�xYDf��A.������j��l���"�rVΉ{�)�g]�b5�p��pk搔^ˣ��N���^�z�ɼ�f�(Z��:^�p���I^�V�֝�R;3Q��'u�Ջ$��$��-�.�4R���ƄEQ˃��t� �V_%��a��̽��x�h��ھ�N��nln�]
��nz��y���!1A�0�x�v�n��e�75`͟Y��Rv�M͗p�"���"��o�b���B����|��"�/�Į��V�g$�w��)oDc2�y����}ieTo��-he`���"	�*����Ý�W��]nm���@�+;�ੋs.jf��-��'��Z���*�)���[y�`�RSWS�	K���;P�B��7z�1)�׌k������Ҏ�W]�]_d8�8n��&�f���8�(o�� �(�QQEVK�T�DT�A���0�2��%�2ju����Ǐ���?������~σ�dq-��&��1s0�hh��*�2"02�$0�q��Ǐ<}�>����^�fcE%&f	HQT�M5EF`dٍdeY9#��3�8����Ǐo����3������S`)S%ȥ�p�` ��k&s2�!��ș�� ���� �Xl�FAAETUFALAE�����RPS���-EA�@e�e`d��%6Xda�dRU%PŹ���	�*�70��1r2ʛ10"��2p$2ȉ�y�G��.�E,IPPĵO�1jm���"��UAT��6�4D��M	�Pd�dEE_3tƳ2� �����(�
Z�����lX�AY�|;�A�������6��o!b�_&
-t��a% �9M��B�q�M��m9/��F�DE��)٨W��軋��{sI�ı�ެ���B�f�v���TwY4���PR��
��\b2L-��!0�!D0I��E��p2�N0�&A�!�)(����)i��Ï��zܽه4�x!8rD@Ye1�Bo!��C)�����h|p����g��q�j�wH)gW��V�Y�[q�b���Dv&��ލ�ս�L�Uj^�Z^�+�l��uÊ�);3�:�9� 6?'�<x��/�8p�E�M\s/4��Yc�b�wmW�(匳�5ejm���5hȋ��'�s�z)0���] EzN�5�Յ]U��\Z��-5���*�w<h�ɭ�v��s��*S�G��G�1�W�eD�>�lG)��/u�� ��d�����Ъ��c�sܐ����ݴ��8 ,7g=k 5���l��Q�Ooְ�8~MCBl5��cX_�2�\6��é/��K�����öP��깬�{�#�$f@/N���^2��(��lG��"zo(s���a���;3zn��0cF�#x,���GKk_G�E�l���J�fAS^�R�{>���W^�P���b�L:�݈��ש��$O'ʂ���U���;Rqp!%潴�R� i�!�$^��Cb��Pq�A�^�|hej�r�Ӝ�nTi@�#��-m�+'�ӷ��������<d�T�1��;{bA_3���J3�.��9 �}���l^��2v�9��]N��B��H	\K�o�l�+���_>3꣹Pb��|�x^Z]�I?������C��;�Uk{G{�@*Μ�m�����k��?ގ7ʶ�NeP*r3%�f�:P*%�7	��olPrOly�U�7�l�Hj������v��}4mm#�wh[���L�beMd.��jq6ܻ�.��`��9L���'6�(����T8�D�۠��)e�=�)�X[ow��գ]pP7eos��n$r<���	r�\Acn���"q2~9��o6�0ko(A�)��0x���w�C�}go����s�F:x_26sUp�#���E�#y�6%{�׊goO{[5�3�`�@|��-�7�G��nC{��VO{5��)�3��*��,'�+{����n/�;H��s�kz�~�w�Ì}v-��W����{L����unP��7�0ߚ���*�]s�b��)�Q��7�.|���w�5v�{�B�Q���n�M��y��sM�nG�N�jRy���OF�_:���Ƅ$����,��;���%���TC����yH�㱆Xq�����<����ͷ�	A���x̎��I�Z���
�����f���KBo5�m�����\gB�+����6����ޝ�9Gp��MT-���{B��x�*bo��c7�5b��vV�#�Uy��d�!u��=���S1�_2��n�|Mj<�S�u]�ŖM��虹.x�]m~�%���f��X�v`��w��C�a�1�T�}����䕼�0�YUUa�UX�'����jm[�t��U]o�RVW�c���CGq����V׭JUj𪩻8�ot��6��#{�2��[�wCsxgm.���{Xkk+��o������͕|�U~�[*�M#8���B��{�=������Ȳ�7zF���lr�3A;a�.�W��ә����_�����t%#������gQ���)&��� ĭQ��AȺ"��,�*'w��u8�$:	�s8�4F��u��!��-)-Y(퓭�me�<����=�pB�������N���@�����uj��|�9�Ẃ�Z+�;�؄d70Z*m��'y[�Y��X�WiwH��n�.��>��Ȳg�m���Ͳ��l�{�]c��ѐ`
G}9���/l��CW��Qǝm�ic��Kgdu�]�Ā�:|!�����雾�U~��?-3��짃 } 7|��W�9㺯�F֭9�mky������S5n��g��$�ջ��
p��O=ύ����}>�oվ �Mi�W����[Օl��M�؆�N�\�����z^�y�PWn#�]����!Gp/����v�K-��7-g���{ym}��Aۥ�-+��˙�YL��+���=��Ye�����fSgU����c���m^Jt>�OG���?j;�ꍹ������0u�1���^Ti�DSKeTK���-
����m�[{��6x�v!᳑�~�"��r���Ŗ��F;-��Q�|�84�6�Q�ؤ7�{.J��NNV�h��$
�s5m�:w�2��x��H*[x��4�����š}Z̽Swe�\��`Ay�k�!���a�&u��]�Y��,i��V"�*abL5�b��C!��=֨j<r�^���N1	RX\���Tp(:\&J��0�.-Q��f�no�e���9i&
����DA~4�6���E���t�D)%�E$������!��U�'U���z� 6�Xz�˙�n�A��i!�}�(����83�ϽrJã��09�4��R��]��I;b�qǷ缌<�cm-�ț�s� �G%�3�.�GO��J���Ց)�6K�իL��s�{�f�O�|�kx@�6�*��V���5�����.�����:Eַ�k���qJ�a�ղ��-�£��.���U^�l�m���ؾ�@'�^I\�m��v\�Y^�#��NK,"�'X�޴�V-�ݥ}�Dob���lCI�3hl�r��¶��bl�VN�D��j���5M?��zC���fv}1}S�<���]k��t)42��zi��˜2�5�g������Zme�Du�*Kg+���3:-%C_ YƝ؜��Dj��w��	�0P�8d]���C�������=$o���8�<�w{�����ڐ<�_5p::"��Ѹ�&c�)��h����a)Py�~x�
����Z��jO[��Cъ�6��c����j�aWZ��t.�:�C(�2%�YV�NVV�q�ﾪZ�����g�ˎ�mDQ��s��q�̫�9m*�J��ǱIm�H�Yf6�HmK��b�%���6)x�|�\�iܵmLel�+N^�zjҁv�7����k�N���Sۿj㔆D�����n��ϛU>��s5G�Vg�l��G=�s͒�~L��M�a�H=�K�W�L�[0a��EQ�R�5V�,Гבp[?��jD�G�5.�{������wlj�er���б76�E�n���M��ݳ�5��&y�g<��剽�tU�U��oѦ�\�F���*�;��6]��E�^՚9ʼIwY��H�>�����aV�FnWQ������Y�j��!��|r[#a���KeufGZ���ۍ���8����4�Uvn]iF�scs:}|�wJ޾t��?h�b�i�4S�������a��)3�JWu��y�1YE�	f��;[�Y �І��a_��Ϋ��. Z$�dA�|"�ޜ�2Z�%؛P�d=[���0�ʁ%�nKũp��K�\)��>k1���LN7ls^�M:�v�/���}��x�Mt�Hc��R�wO�q�\u#*�z��	I*��F�-L�9�%�
�7��j����p���Xv9{;"
�nD5;t�Vf��z�,.�Y}�;��@��t�q�'����hv(�v#^�R�K�;��ݱG��8���Z�$���ϒ�x�w��z�����k���p�6��8��.�3ӆ��p�����-��9^��7ރ<��Tzuee���Cf�1sv\��Pk�j���wP���}X2#֮��K	�Zm�:U����Z�UU����Z�5�C�H[�mbN]n���d�o���%v9��/�xN�`>����>0	�u�^���o�{���� �w@�g�9�K�bb��\m�@�;q���_"|6�R�*ayL����ִ��ƛ8�F�_B����^�9>&��%���|��D}�}�Z�e�g۪��v�2�A)WJ�����V(�2����k�y�1�P���G���|�M�ͺ=|���Q1����K#� '�H����GMvӧ+_Mf43�n��D�#�fP�'%zs[�pbm�g�����Sr��-p�������V�u��8��O��#-&���]B��USb�:��]!���q{:�/��i9�>��8�k��x)W�u9�����;QO� L��x�|=�>@@����#�Ա58�j|�v,��-l��*�+v��c3L�	�I+tN�k��>51����]K���g%>�,ucT���R�e�.:���/I,ʂ�<��!�ez5o?�J,�1U1يn�&+>���3O8)�$�K��%,��G�VOs;�e�>���F�_���h��h�76c���5):���S�vՄ�֝�3�>����BKve�4�d⾨��Օt}�DF��b+(��i6�� o�G�ЎJ���jF��cs��r@m��¤@�3o�J���#�k��d�������b���C������Km����|�����o�y�Ŀ~3�wG�	y��p`�2��R�k��ֱ��5��%>����T�{��m�p�;����rX�qut�t���װd�<.S���½�T�-6�9ڱ��]ݸ ��m�+Vv<ɚ)�1�Ύ�.��ŕP�Ỡ�y��*�7P#Λ�^�5*���˴�A�L47j���|�Zٰ�(��L'�2�����B\�p!}�
�������M��p��w[�"ʛ٘�Ȁڇ3����ms�o~�Q���>�i���.�l����L���5�E���Q霧���=��}��x��I�S���v�.��-�|��m���n���)�"n�H�u>�ajy<�`OC����SQ�|
Z�>S=A~Aw��<�;W��1��{���ԍ�"IM3���uh>��V���D5�X�49^��w6@j����ҹIEa�~9�T���%�%�#�^���n���v���f��3!���M�f��m�1s�{|���<<3H���X�WJG��T^�*�{�2kƦ��T7�Z��+�x[����էr���@��Y�������mQ7�\k9�|=[!�����MN孖�Wa��&l/^1U�C�QJ��ʧ��`�(��լ�ж�Rs���^����M{�r�y��V#a�e�]�*�g'kJ�W��'ю�]b�ƯU�w�Ɠ�%�|9�z^/VF�-�0*�ayf�qܮ�.�]�����P�}�JW7X%vz�yNR{y�>�+z��������빳Q(zSshLl
M�.sky:��j�8��f^��W999�m5J�}�kW�q��J��ǟ:q����(ƜEB�zX���%��3wD�n�ƨ�`��89Jm�)��8h�uoܟ��T=��V�թͻ܅����ގ�����an���5�ė{��Z����֤3럵�[p��8���6��h1����Au\ج:���S[�۽=Vŭ�ُ��x;�h$o�JWR˭vŞx�:�fc����F���K�J���a:����~6xv��N�X�;_�Ө�'�Z�V��;�%��V	��̧�`b/�5U��I�H�!<�P��0+.��N�fs����u�����2=�E�]N��M$�Ef3xz8e�8�򊓷����H8p
�2ڠښ���y��X�-ox��7]���^BY�S��@r �dP|��\Ż+����[.V["�Ve��Z�&驦�'�Yi��=��A8(j�U#h��^�W�ֹ��/��#wyB����%�@fV��z�dX���v�N��\�
�
���sV\Y}WD�ٙ�n��2�րB�!�(��s\21�qU�ל5����������HWK���8�&Ҷ�Ĵ���P�X�\c;t�`+��������G���l�Z2��r=f���8�G/��#�:���J�mu��GV�ݛs.���ohF�r�ɐ� 8�=ٕ%�Y#��� �:�>��[Q��D��V� �\N���{m��ֻ�y �{&�}�_b��P�3�y��[�Cz�N��TֺɄv���wvb�<R�	�0�,5ج��"T�l�P-�����kA}:B�C�\�5Cf�;F�ₘ���`�3U�%�k�uhQ9��Q��.9�c�1�3YxvW�d;t'S�P���)ѵJ>��
�)�L^�q,�Է�
슱o;@�r8�/s��{ ���]�����+oo��8]�Rb�����:�޿'Me�����g��C��V-����2oyH�]�pNs��U��������fK�<�����oጻ�Ѧ-:V�43;D�v��۳-��Լ�t�nξ��ݬ�wcӔ�1�5�ž4���pQ}�Q/���d��F*ؗH'9\�I�ӯpǷ%� ��{F�t3���!�r��Vˡ�cB��`L��0�љ����\Ƒ%;�j:�0-�
&pv�6��z�V9S6���2��vͻ�0�CWj����5�.ZxP����/e �g48�����t�S9Ju{��[E.��E�w��h������u��E���@��>J����8v&�%֜�ps���n��j�3TI�2�̘؛ox۫_%���6o��֘��<��	��crLBv@�b@�Q@��Z0��(���L5�jY�[��
�{̚^|�Fn�|A|��Y�S=�C��N|���qp��y�^��v_L���1��z��c寻�N�{����
�	Q��ۏ�q�۲��1���#~J�c�Ш;�P%ۖ���Z<��;'F�X\�Z���J�	�K�U��]`��u�A��'_ׅN�k���y�r����4����WVES�,;����6u,rp</�M�e.��-��c�<�f����H%�����
��geZ�%�0ZZ�v�:���<����L�*�g�D�,��ᛳ6|������+(�}k�2b.WH�Ie��/B��sKJE�J�����C��-Ǻc#�T�vVeq��-e�����uY�9fe�w��xE$�[7��ʤ��õ�'V�$�K��ؗs�4���f�ߞ���8Qlj�M�L"i/Xd:XVfTE-D��${g}=x��Ǐ����=>=��
<�-��B���0��
�2�$�����h�a35�||x��Ǐ����|x��Q�I�;$AU��QPl��QC���ٙ:3��><x�������><zy'�BUR�$A�ni[V����,�[;l��l��[��d!�8���6����9��r���7t�ih����QCldf�� rL�`��	��L����t�����W�ˁE��9�i�d.fffE&Hc^`m�Q.]�\�����x�NÑ\�����	�p���)�Q3 IdPPd[���?l�(�cfr2
+$�1*��Z
h�*`�l;<��$���]U�&�j3vu�+6l$V�j�����Nֶkv<L�����F����u�]Z�f�co���bnƴN�C34�Fq�����q]����{f�f��x{�]A����k��"�.�SU�
9�7�ތ8��OKt%�R�7�Q���6Iݑi+	��%N7sbO�3]�I>��z�8�LT�[�/+u��R9��5��1M�\����:{�*���O?Yp�WsG��N�ޮr���Ϋ�'�_���빺�[��z�H���>��Z�'�$:O����:��������(����T�X"�k���lM�y����ȥ��l�9���r�i�nx\�X�3:�nۢ�f�[���
;�@��H�G{6=�����ZMR�S��nK^Xh�-�=<����ꩯ�yN�^/'�C>�^l�\c�˃Mí]�R\a4��ыa�NW��wa��2�qBG;m1�6Y���3B�`���~!�ޑʽbҐ->�A0�Ƅk�vb�I޳|�<�Bc,��^�Z�?T��uYם� o�W93h"ˡ��s�&��͸u����A�yS۝Z���jD;F=��I|�f��++%hv�i��0�I�]�hY�ECbxk�ޟ����M�rG �w��n2=�ػ�2�&&}�\�e�@�9#I�i��9]W7�]6���������s��f�B&��\�ɑ3l5.��s�rg��A��7c1||����M��+��*x̻��W>f�EO���5-nU0���\��s�#T�O������i�T0�t��k�fW��Sͬ�\��c �sqs�ƭ��.g=F!f�BWu^�9
���fJ��ۊ�쮪��K7٘2k��Բ�kr:y��	��*�UND�L�u��W*��oLfd�|�nr�\��"�Xqih�nY�Vt�Pi0ՕF�����J�Oe�`�L憶j�N�AvO\Z3�̙{�ZTd��U��]�zs:l����ݴ9 yVx
M��<��}}@48�X���+�o7�MT�)�,c�����X^x��H�oλ�~����!_�s#ts���/Vt��n�âun��R�^.�&rm=4�M�E���֌b� J:��;HvN�0�˵(�i��f�G�	-r%�3}K�Gn�����]�J0;��y.�m̓� E���c�><1��|n�E�s�7�}330@�Ab�|��
#�㴩�E:��V��7�zx2[i��ETlBB���.]���[�Vǯ:gO �:��ue�F|��d�m�}�����m���}��{��p�L:ʈ�w4��d׶,��0;3x��ٱ�p��"�j!"b/�$=��ۚ�F���tY]�{xΓ��ڗ'�~��2͙�ڌ�\DQ�]�����<�}"�6/��F��Cc�m ��!'/��n��n���zd�<���f_��B�",���sf%ozש�<;��?�l��0n�F`�4�A�u=��b��Eh���IF]�<q�&b��늦q�����D��v�i�R6[�bOJ2�c�o�I/S�}y>�ȅ�ۡu���N'/ �����Ս����Ɗ���gd���	 	  ;U�w~n5!�j@<����+�1L"M,��)�)��`��c�b.z��ok�P=��7U��U���p=�)j�S䨰L�6{!ޚ�\Fx�Y�uZF��=0�"'�-��	W�)�Ro�_nN�.JR-����9N{�+�������AÙ�����L��v�����#�������
�!��d�3Ӑ̤���f=�b{�M^�V������7���c����X��S⯣(c��|3L��s��]�a�3�� ZY�֣}^�!Ň�wZU�J�/�n��
��N=�B�|�s5���ʄ)c@:z[P�t�V�O��[ε��_Pl3c:����/�Q��|}N��lV�v�z+�l��r8��<���U=yܚ���s�e��z<zlT��K�6iD��|�%ܬ�ЧZ�q�OBZ�����[ULT���vqwԲg`Λ�b��c�+�Œ����Q�����O	��2�]W����<��y�̗yW��7*�ʦ�Lp^�36Or�|�!�U��j��:����[�'�1%Jiv烥*yߩp�ˣ����U�g�z|���s��p�e�s��z��,ѵ?g����ʏ�����4�`�W>l+)p��T_���{,�f�S�A!��s5菻����~k�R�Q�C[%C���cl����vW`�S�Νs,X<�]�U���`�6mˇf�o4.�����.����J##��z�.wfA5U��t%�n4f��;�Ͼ��0��9���W`�gKm��窟x�B�8U3\
"K��۪7y����wG�2 jT��"n��U�|�E��u��&6a��֡Rǻ�م�C{�M��K:�ᙟ<����f�;r��J���iȷ���]�=��cxBC��sZ�cڗ{���i��69��jn"W�������962g)�!��%o"��}y�z}�T�WrAX�>��Q8�0$��^n��̚f�M�5y�5�v��K/�.���qYB�&�#Vπڊڛٛ��]YL�Nn��N��7E�i��.��<�l��=A��%�|�5 6�x.X��v!����y���4�w��
�4ӭ��+T{vV�1Z���z��ʽ7j�]SeFv�t��c�=�%�O����o� ��4t�s��'B��u�,���t�&��'6٨c+�R���f{3e�f{M��+o�$��!2�U|��9X�ֽ�e��#�岝�<�r�z9Ce]����M�D��i`�&��t��l>9�� �)�"�c�ەz�w�5l	tla#���W�g==��sO�{�E�~�u6������6��m��v/E��Q���d-k����`�6�dH������6��*/[:zX+���јU�i������ǯ�2�N�<��,��@yޮ�ӳE>�`���^p����wM�q��N9���?7L2h��l�eZz7"r�Di�PC�v��>��09Uy��������46U
cMWI���e������mM���!Y�}�`ʦ�2��)u6��Y���ghT6 ab�vЏoS�M�^|�]^lPmLMmP�=Z�U<-V=�d����7����v�/��p9�~*���ݳ>Qt��[�&&v��@Ga����	��6�qc�Cm5S3C��n#�mڻ��u5:uO���<�W~·��e���]�g����YmԭC5Ԫ�4�#�kV��Ak��ܢVn�t���*�,���4�������/z�N�eb>s*@<;%b��!�Ŝ���zF��؈o�cc;=�^f�J�'�]='�8C��#�}�h��.�:�K�Z铐g��7�HB�(,�03Z��-�T�7]�Ǽ7���+�#��T}������&؟9�ׯ;א���s�	"�p�ca"��?�H,�3۱V�q��#�-�.�D_�j=~m���ڪ�}z!f�n'�?=���n�Z�Ci�$]z���>�����᲎���;<��g�e-ܐ91P��c/��,����I�|��#*:j뭉��꓇r��8bg�j�WqVwO���C����7�&�^e��,�m%��78C���*ɪq�Is�\{�-#{�}GY�[ea虉۱���֚jݐ��UoO�<�4J�] N�h��Ӯ������L���b�@|��dX?�]���oI�YGx���:�m��n�n�m�L���F��ހ�}\���3�&�5Y���X���6Q�135y�ŸM�6ϭW���=϶v�-x�,3Vy�l�c���[�A�j�/Ҷ�:���ʓr��b�#.��k7t��&e2����㟓�d�+,�m�Z"W[2u�D_l�)��i��J4:��$��j���H9��hEV��a�9HpJ�KO�l׻ds����cLc�_&R.�ܾL�t:W�7��J�Ȗe�
x�P�y�t�z(Fڬ|5v�Jl����r��~�<g�����L�-�R�h]�P�N�S���v�H�}5ln�ـ���|��ڵB}�7����cCy])d�sq5�R,�0���r[T��xE�⻎���)��6]c�y��}���n��#r� 9fU�w��U���i\�3��	귽6�{����2v�v�3�Mڢ��LDL�L�EǰW2���=-[���8���n����8]3g�����lqVU.��h]d��oq�����ʬ�����ˬu߫�����ٙ���6Q����Wg�m��+� ��|��(�v�h�x=���h�wG���"��=T��Ry&|�&��\_p��ގ/�2�P�'7_�Y��m�>��L+ޙ3�1���)oO�Ʉ�u,�4'}7����Kt�gv��a�i2 s �6�ϷǨ9&@u.c�ga��w���wa���}�W���\�@��Ѻꓗ���z�I�׼F�E��u(#jy����;����lwM�.����D�&�.��l0�	���f���P�(goΤBض�S��ؠ�YΫ�m����X>'Q@�o+�oZ�k�.5��{9o����ƨ�^G��o_�X�1p��nj�OsSS!�#���m�����j�֎僵�^}�OT{zC�����NKy�F�{Q���ߍܙ�EV��E��� moo���c=����l6��bCp�,��7���d�^a��˫�0�na��H$X��%����n쓈��vr'��$����{���|�Y1v�{�y!��#=m��>JeP&ѩ}|����eyOr8gG�2R�&/���V]��#�����C�s����S���,����[u�,2���۩m��t�����R��4��+w�	��c���A��ʅ��mJ����52�wlj n�.gCPf	��dm3�
�5圉�l��J�R�G!Nh+2��c��-�5�mn�Ǝ��[r�t�]����`
��'�P]��	K�9�ie"k۲�!SN%�ח���!�����c}�T�E��.��W774��{\��Z�G�'�aO]��wB��n�=�-{=F�#T�#��� �y�͛�D^��KiV���&m�t0TdJ��,�9�ȟ:��i��%u���&��ޕN����r����7�a�_�\�틌Z����!g_�&}}��u�����&�e�y�Z���'��������%�i�o�SQ��+�����hފgNI%��=�'�1�z�g:7]{;ﷺ����+D7^����.6<))pn��+n�^H��:��N=gI���;���@�*}�7��$2��Bޘ����x��m��㱍���o�	|+,v��9�G�Ƭ���3��-p`1��uT�͐"�����(0l��n��-�Z�a�O���i���D*��zi���6�` 6�[t�[�Mw�k���m^�T\V1l^j��y��cx�ֆs�w\4�Q�� % P��"��dMu��cz�G��������#��"�T�Me��dٖ�h>���ǡ_LM�`��Sp�NT&�j����[����(�����46�ߖ}�w=w�wׯ��������_٘�ꂀ*�����_��?�@Ds��4���	��}����\!�HBa	T� F�HB!�$��b`BU&�dR�A�i�a@BU�!�J	�@�S7D41C7tCET31wD4y 	�{Bq�@!�
�!�B�!  B�!
�B�!"�n" �J���B��@��J���@ ! B!( @�� � �J � �J��*J !�B(!(�B�!�B�! �B�!�B�B������B!J$! ���B�B$! �!"�B�@$! ���J�$��H@�!(�!
�B	@$! ��(C@�$!(��BP��BH! 0� ����4�@�2�H!(?�����0�G�AI� �PER`�C�7�,���|����~��G��P;����O��������?��������Q U��������� �~�
 ����P~�����i���?��� 
���X~����H�?��O��o������g���������QP(T��H��JQ%�I%	T�D�E �H%	T� �I%R dRXT�  R%HT�����IH��IP��`$XY��a�e�`�f��` Y	BE�A��e`HV@�a%IE�A��ddX�dIT�d$Y`E��hE���d �e$FU�`Y�hF`Fd$bEQDF�
DB�?�@�J��R�J" R�R	H�H	B�4R!H%**�!J�2��B�@�B�ʄB�����Ha`���?П��(�*%"-""%�@���w����������>���
��������O���1�@���?��'��@P^��C���x�� TW�* 
�؇�a��?@@?!��}���*�����8��оh``�3�='�t�><�p U�D?��g�@p|J�����?���9���?��I���?�|A@}������*��~}��'�?za��`|O������.�Ϡx�~��?g�W�{)�����8����~/��;��� */�<`����������/>����1ޟ�����)�� �����0(���1 �>\�V��Q%$�"�*UQUJ�RUBJH�BD(PIUR��U*�T)E%TP�*T�(*%TE�Ul�Ԩ�AEUA%*��l���**����ZB)��R��D���P�R*�T���UI�DR��{��)J�T�!J�D�D������ EEBREH)
�R�J��T�֔��(�m�!IkU	��$�X�m��*�]� �^�m��V��XN̗m"��+Mm���v��T��Үڕ�f�)SR����%k.�\[TҊ֚5���dUYk��]*��mV��[��)E�Q�5K��  \��CB�
(hntp�E
(hh��S��C��B�
9�����K��9n�ۭI[UP[fY��v��wt��M�Im�fڪ�m���v�u��ڒ���]d�$�UK�AQ����  ��-k5�b���Umkvrv�����eM��n'l�P,�V�[[K(mZ[5l�T6���ڭ�����ʭ���N�tj��jCSkvd�f�(��JD�REGx  s�{uș�Y&eRUjʪ�UT�vR�&��6�̬5��6�*�P-�@�Z��U����ښ�iB���P�JR(�0^  ��j��j5PbSkD���Y`bF�)�fڕX�k@�klR
V���5����-���h)(`�JPEEJ)D��   [�֘-j�J�*��#eEV��LP���V4�D݇"�!]��6ʕf]���P�����j���ER�I*��)R��"��   cĂ�\`�  l` h� �&� �S*��Ұ4�5��  �`  &�%@ Y%
T��@�
�AQp  p  �  �0 ���  Ƙ  4�� 5�  �� �� �Y� ��j�)QR%JUJIUx  0�t( �+  P  �3@ dX h�@ڣ  4�Х 6  m��  �f%T�E�R*IERJK�  �� J�`( �`  -#��	����f� S4X( �V � ̬� dX �"m���� "�ф���� 1�L&��	�)� ��F�  j��2�TmL� ���M C5=�����ߌ���;K���Bܐ!]g��,�i�P��b�/%3mQW��� >��}����� ""��U�`����""���EU������~?x�A�Mnft�=w|wy-�ǖ2*��:4r��ڒTi��`��t7��w+T��Y0����6���ʒ� 5�z���YT@���n�Mbb�ҦʬX)GPY�]bf�f��Q+�7�l�a$ic*��׀��e
@'��Y���,�S�E��.i�ɟګj�K�]Y�Y&L@�;E;�[HJ����M̷� #��b�6��l\'m�V*��IXD�jR��R�v��&�M(�kÔa����NZр܅!�Q'6X&̕����K7�V�(e�:��m\�ъ�T���͹���K��G9��w�kV|�Z�m��o5�(�6���>ɍ�/fV!0��f2C�)&`����w1��4�F)j	����0��[f`U�e�[unVLF��v/h�cS.���ѩ�Ү�ǘn��R]a��6S�EAN�K�2�!@n!�h!��x��M�%�n`�(�Z�48c��-�5`�0b?��LHn��x�e�;��2
����5fPgU����2�ݨ�R�̂=�7/l{W72�X�2�؊���5��;e��.dPX��g于ٷ���Y��ʰ�*m��[F����Lq^�=��`�a�S.�m���fퟐ���rS�)���*�9��MNb���ɭ�����R��I�D!���vtiz�]�Oc��!�(Sղ��мU�NHء���� t�MBخ�!s5��6��Aۣ�+{u�B�Ӵ�ҙN�j��v�̧F
Z�v>{��QїtO�Ē������R�7g,��R��ѡ�e�a"'P�q�(\�6K� bR�@6+i���W�%f]�ioҕ��"�߃�����Ydl#���t�=OI	bT�;���Ԥ.�נ��Ef�J��4�IV6Jӳ�4�t�l]��b�QJ�!Vfn@��Ae/.^jl����U��հ6��(VP�d�D.c��'m�]��'1�J��p��ޑI"��/+i��\��W�U�ȑ�/u�I)�@�W�;��=�72��A��R����E
��:7��m4�pۙy4�du�W�l^���P���l�R#�6�
������.����+�ӕ���Mhl�4Ę"�·���c��*�%���nx�j9��4�k8ZR��*��h�՛ێ��(uV�T4�ٷHP,]����l�Z�j�b�l�$4��K1坏^LZ�Ӊ��3�=f�Sf7����^Tz�z:ʈ��Z�ݡE�c.�B������f �"�<� Z3kU�9 ݺ;n�*�C�%LD��/%*.:�Y�ۧ4z{yb&�fln=C��IN�{�LnADҭ�FE��\�����Ù�� ��Qg(�X�M�+m(�=fSNf��p֚v$�8�e$]�xd�X��j�D����9���ۊ�iǹ���*R��oU=4 l��Q�sb�qb�7r��*m���F(�O�ˢ(�jӧM<q�NX�p��Z���%ZG�mZ�g!�VL��b���/��;�Zg*\��"���-�YyK�Y��&*�'wgwmX����O �[�fӲ��JP9f�!��6,̉f���ષn�$��(SV�i��L�yz��-��мXR�~gV�_^�G"31T������Y�ZR���?m�]�f�T��d�K��׆�� V2sn������
0�J��Y�/]�9J5�d�ov��"�r�݊a���A�w/ND�z2���sҏQ)��k���a �S+nV-�Ft�V�CuyjN�遾s���qR��۰�i��S��eʴ^[���+Hl��?��9[�<�4`�{�:�&�Q���{t�nB+8���2��V����j��VEq9Z���HK&ڼ*�j�j!�+t.*���t��0,��)��f�Z4����1 f-�n���Bl�Xj�7`�Z��UM���İT$�Q���h��&'��d���MWO��gL�i�D	gַ�裶��S��יl`4��ى��m*e��W�㧩-��ZN�̹a*f���qiV��LV�:��cV�q� �.d�qRͻma�*G&��62���ˣ�y)mbEa�~i�%����2i��y!PeF&�P���ԑ�"�kU�*��%�i�9��k��������M33nQvv���r�V6�[Cq��d[Ch�{fk�4�6�;�7Z�V�X�ՕN�Ek%KLM�`ԭL�j�*��H�7�1�f046
��qռWR��t�D�@�w�)�5��P������L��F��9M*tj��5�aU-<U���w[gc5�����	6& �5�b����[��)M�l�b����Ck(�����`v���U�Ty�7E]��~[F��qE��ּC�4�q��U��v��-�Z,`�f�G+Z�A2�A[OC��+!�)���,�t͠,��Puv���6����;v��DTT�9c f�n�'�2X�j,`3�wZ[��h��䶦�}�vkrS[&+�I�����ث�T���2�׃K�c��2򞽨H�d�7I1a��F��:)hWr��`%#7��Y�އ��-�hLS�)-��Y���=@�T/+M�JhH�]n[�\&\�lFn���6�X1*���w�/����Zx�)���˙�v��������?3��l
���M�5a�-����.=ȭ�z%�"�+�F��K��U�iXO5m�4�Y=�;y���?n�ȣ@:�a�2��)��kUz?��j�q�բ��S_�s!��Z@t�F�2�YG���a
߭К���	6���%5���2#xFAac
����ty��r�I��Z�*VХu/lT-M��&���>x�h�oI��
Z)�1�RV٤���x�;��bYq�yw�QM�k��
!,M�0��G�TkZ)^�2f�Or(5�R��Zp't�Toh�����(��=��!yV�wQZ��鲭�o*i��va�d�7Mah84�� ��`f��rk4�*v,�L��[��i�E�L1/�a��B��q���*��hh`Yc,,��4�%Q8رJ�L�{�=���dk���I*�]�P���hn�ֳ��F��w�1�{�h&ٍҤ�;�Ze4�;�����͟c�+!��1ͥ��sx�t�ne�S)��/Iݔ�B��2�Qll�.ٛ��P�`F��
�]�n�Y��wf�;��[�cJRW����mK4>mю5��0�nae�tH�4B�t�|^jfqJ�&4��'u���[��*��gv�M����*
.V��o*[7��w\2����YKZ��
 )���܃r*���۸�#1�@�ŕ`Ә0DN@�6��^��B����,��sw~.����v	�su�#��`�l�t��LV�;K&�f��ӯE��%+�+U�n���f���M�m�q̬�!���
f�[?)<�����=j� ��`�Bw*�*x��j,��.v!;�`�+S���k3b�
e֥R��/\U�.�h���P�yt�-�`��ͬ&��nT�$f`����N�xXSw^M4Vd�וv�c����q��R͂�+�C���Q��X�4�oc�`�ua^V�e��Z[f�Gr�{�:�/1LCez��sv`6\4�۹`g�E���^�i��͢��0��t�0 |S��6)T�,T�˔���I��e�P�n��]��^bڑ�i\��I3@R�zE�ι��"�S��c*�ڏ([5�Aa�MF)��wtQ�%�GE#w�+��nT�ձ*d��b��L�L�؂Y݁�B��yN�ڇd�m��kB��YnӸ�я&���
I��F�M:�n�LL	"�E�h��0�3ê�N�%��ld�� :ؗ<pX��<0���$^�[�`��؇H�.l�!P��*�r�R��v�&va[���"�2��h'�
����V��5j�e ��S16�$n�o*&ا<�Ѓ]"�5���,��&eL �4ֺKU�BK$34�%F�^т�qK��N���ɰ��Ų��Fc�ɺ~�[�H+X",R�;������i&����];9J9��,;B�2���ǚ�nk���y>nCZ����[N�HQ[�al���dֈЩ��0�zm]�5%�V�6PۑP@�$�=�N�U��3,�YF��;Q��sF��mF�6��/�*ͫj�
�E�,&�% �&����
	0��Q����7�ԉ�#u��N]�����ME�U7%d��P
�,w��Z�EŢ�)ʑ�bYK�V70�#�{)�q��&"�)e0�&����s^�Y4��<b�& ���b �4e#�1�[��M@V\[�cw,OݩX�n�Q`��a���	�"��ޛ��M��Ӫ�!�2�3h�����0(Z�i��) ]�&�ɶtjd�ΡS�s%��SJtl]C�TM��η+5Ӭ�u���VV�.���1i�D,��J��t˺5 ��D��R�p�Z@;Q��Zj]��Z$��ˤ�X6�R����Xi��n���[N$�,��ӭi	Ֆ��+@PL��%Y�pU��+���(u��t_���3t�R-S)��B�A���4�M0Q(�A�7%X���f^l���JPQthd;4�jmM���6�n�v��V�v^��rF^�jL���ݚ��wOs�	)�Lh5,HYy�Ղ1�L��N��P{AY��n= uz
�R�n�v�e ��̖tNu����Ӂ��hTf�ٮ�w^-��Z�|��i��o"�V��t�qeԧw�ѻr�M�"j��Cٌ)��Mj6��b�?ag,껈;O:%f-���6�5�Ԭ��B��(�Y�v��\*��M���eM�D���u�o>�͈�OI�S����pX�-D�e��fMj3
�iՀ:*%���A�m�D\�l�hU�����a�� !$֦$�)h/Fe0��akrV5�6�Ҳ�`�a�W�n5A�Z�i�iΝӕ��-�$���L�
��i<�!�Ѳ�f�b��V��^�V��/D�	�1��M�R��z<�4J�dHỬW�>f����H7I��)�րc�v�a�w m���qQɆ\6w�j�
4\��Hn��Է[B�9�uC�J��p^l�9+V[�,�n$j�[.���!��f��%qJrQ�W����Q���ot�%�����`��^ǥݛ�^0����n7�rn(V"�*��b���;��ڇю�b��,�Sk@V�2T@k���T�z� T�T�, JK�Ӗ^.�0�FFr�%)i;H��%ۤZ{w�ѫ����j`�e]�X���B�EW�AM�HT���7󺊃�D�����*�nX���֒�ee��Ve�Q�6�h�E*)U�լ��aR�r�i!�Ĩ��	"�a��_��������S�ƃI�" �v�a�b�fQ��BѲ�*�!8)�(����x�n��4˼0j�!�ynTk[Ae������8�ǖ�	QD�M�K�h�����ն�*yw�Hn�����/@�٠�A.ҽB�ͺ;�'ʯcu�n�+*A�R�I�U���Ƭ1�I�c��:��bU6�+�H)	X��+fn3�'$U�����ch�����7�'� v�Ԕ�*�ͭ�R¨d"��=��a�k4����j}��*[�e�D]e�J���F�xuM
w��2^M�r�
������]H��^�uo>�\ڇLN="`�J��-�5�U��^ZLF]����ܭX�E8v4�3R�,�!��
h�x�LL��Oln�0����%�o>ql˭ں�6�էFX�K�Z�n�J0�^cE�n�)N�X~�y�M�ܖ���5rM�H��6l$kUX�ܴ��Y*m�f1jS����"SC]�P�eK��"{*-� �`�|o��mP
5��Փ,[Ӯ�0��N<u�d�P��6�WP$\t��ʃ,i1;cEX�.�G�>&���u�S��j�2�v�֮^�It�����daS�+P�Ĝ���V�:
� ��n�Ӹ��a��^�%����Tr����bRKӶ���M2�֤�^j����3�e�AnL��7�Mot�.��,07!ɍ�����a�ԭ����3%A�)v�w�����u�K�
֋Y�@ŦjB�z���La��H`'���(Jf�@��oY��¶&�+^���<u(\B�M��M2I�	4����Z�Bý���׌�0P�K>�z�b�ڽo�d�J�Y]1m�/pZ4�'
���Kp����g�ob��5�����RQ��юl�(<U�c.��
8��Gq<C[K �O���E���b�t��;R��� �f���u�` �>�:F"�Ў���=n�<��\,٤9/X8(&�d����xD�`��u��������+6�B]:ZE GPz��$�ӛi[DMKn�@ҵt�	vrf��A�b1S�R��Y�׀���<��";y4��;�L�)�(���M��[��!�`Sj��8�C��%��5�Z� L,YA8�[V$���)��-����j��L�Ad.�=y�(9g(<���0��M���S^P4D�U��J��;;$vE֍8�p�M�v��[/�[Ëwq�o]f�ɛ17p��e
OZ���lK�@���ZR ������ڀ���%n1S�w�d�E�ֽV�Yc*}��GK�WX0F���X����P�+��^�l�!Ř��f|��f��pCMb����S�˹�q����r�n��R��3�B%[��c�w;�u i֨�n�=��tE�0�P�#z��Y�IPS8.�&��6���r*����o]�d��ױ���������I^AV+�Ά�K�Y����8��u#��lq)5��#kZ��K��+�(�1��ؐvw�Sh�B���b�#Āq��ڬ�%u�B�	7�Gֶ�S��J���6�V0����^��e�hX�.�s@�kgf(ED^7����� ��Վ�>�{�&H�ї�a��e�������/���rU�Of,�\����ݺ��DⰊY%�I�ĉ������Je&F�s�'+ښy18�UyA���7ӻz���1�����;h�i���TB���j9}���Ǔ��]ǐ�NR�o��*f\pv8��תZ�ޭ��@��I��|��w!�����e�(
s��sص)HKK�\m���������O�J�
�
y��S|���n�� �t�o ��2]e���3VӮU�-
8��JỨ <��\YI3�
P�h��)�1+�1)5��B�-"f�/%s{�t7����\�9U�v��.�V���+�kۄm0n1ky��`���\TCk�ăK�Ҹ*ƞ^YާO�1ݱ��m�h
�m�ԣ�P���C�5-�����<���Z�omx�[=a�^���$�3+�B�e�
j�.����u�xѵ ����9]r��(������0z.v�u����� 1<u��1c;y�l�* ��$�(�Iy���V8Z�U��7�)V�/sAe˾jX�x�6���o����e��痗3�-_9����*��)�:��{zehq��t*1֙���z���0\��u��D'�7[�]$��^�N�v��v�aj��[�/�d��4�Ί�6guel�C��v����L�.�9Lr�$���}xD7���s-�G�*﹣ñw<''��X'?���������+T��a�T�M:wӂ%QL5��7�:��Kq�%�6ު�y�d�KB���I���g��f�J5�ևADM�߸1`E�6�)�L��JG�k�ݬ
ׅ᫠�Rà��e��G����B���m�r��W�Y�FdИ�Fm�Y-�:d��t*,�]m���ڲ5۔�N�2�]+Ej���M�ۧ�3&��r����n�hY[D�5�۬����cz�A��k�7 f5�IL>�w�^���]2;��,�^-� \�L�*�̴aY[y �ħ�T�x2��9��(u����n+K���g.�]|�]�7W�������t;呪������ɝ�7���z�<l��0*�82pR`W�!�fPů���d���X_Wf���j����s����
����maN����N�vA����X��"��R�+r�b�զ<�ͽ�#�1�^�x~2�����.�WE�%D!��_ZZ�jQ�c��s/Ĳ�́ 	���t1���ނM�XɈ-iB�^r��ovi��m�Ɗ�h ���[f�f������~T����:����Ѩ��a��o��*��J!=�41�a�y�(@�+�.}��X�#m�\����[D���	�2t4�V!t%eΥN�t�us�t�KS2�y���Wj���g�0���+2cW�B&ެK��YQsK'Wn���������nk�!`�D�UDl]��&�7%�֐�U��������u�q�q�a4_Y�hc����C�����ּ���b�p�b�=�RwF�^]vgg']������0%����!g�v�޻��'+M�  ޽ʓ%�tu}��ʸ�Dtz[Kg!k�P�Ԇ�'w6�N�)��[�$�<��:7�6˭{��ݐ#%um�C6��#F�/&W>G��J)��ٸ	��p�Uڅ�Y�\{��e�\͊�d�ݍ��+½�h�4��O8�y�L⮹R-�2�Ro�_Up�R�oPS���_q��	��S����L����W�wB�ѵ�sb��Er|_-)�|�T���9���p;����$�s����dQ�!wg4����c�Z� Ή1a|z����	�-��u�mip�+�"V\s��s����o4bB��]׷�ȭ{Y�=RT}��.v��vnj�!��N��xA�ޑ��%kLP̑1XX�ڡ̾GV�,N�Ĩ�N�b�c���~����)kŰf��U3;O(ҹ��R�}�j-�A(��v�TY/K�k��6Ђ�#v�-��N�	w�9=ا5՗9M�.� ��u~�|#�,�n��1Rk��2��������&M��H��Z5r淰>�3�]pH���g �|�Z�;��6�|E�L��Y���No�7���/t����K�tB�
X��{ݫ�S�]&v<�t��rӴ�J��r;36��(o��=5K=��+e�AP%��P>��v����[�x��QҮgo[�o�lb5�vk/
j���ގWf�2\�tF��^�V�.�����3!{�[Ɗ�.�끏��L���G.����&�>(V��0�q���ۧ�o�RW/88����T��w��}
M�{��M;A�}�֜��kw!�YE�Od��j�7�M�3m�]�U$_r���7��*�j���X�Y�ͩ��+Yث�5����� ���;Z���D$-��nW-�Z��rNA�{z�Yv�Fo[�Zu}�L334�B%�<[�.��΢#Y��1^P�z���c���d!�U�8Pm�y&^QsbV���V�kU���C�R4��
q�}]��� ���<���8E�,^���}��	� ����/�&V�ѡO\X���IL��n*u�)QZoAJ/���|���6��X@]�!�k��iTQ�o��=��Y����ُ�Y�8�zyj!#$���w���#q8L�m�Uî]?�����'}��x�>�R�A���,����S�T�M�QP\x��p=诬@�X�(u�i�T����_)r�R��.9LP�T�/� =}C4ގ���b�©��:!,KA?���� ��P�kBe��T0N��m�QW=m�wN����#X���?�̥������h����ݚ!�A�Yz�Q�W��(�Ű�z��QB�Qbqd9�z�dtK0��[y�֝�䁊k຃�]����&ݥ��<�Ҁ��z���Hh�۰�r�Kp�}qn`K.����S\*�i���f�v	�G[D����H��/4�U|��Yr�ܹ�X׳��� ���Vv䣹"�{����Ю��y�kӖ^u�q��%�-�cq�+{�\���f�|���/9�8��J;�	{YȎӽy͂�v�YE���y:w��9(�g������J$e�vq��	��d�cɻf6���&�Kh���O@b5�W3�����m�]�
�;��)�� r傸iْ�(���l��	�Ӽ��ԗj�S2M��ɏ�.�w-����P95�Bof][��F+���<�3M�V))�V2b�v�`Ku�d2NL1Kq̖���!;��YI�8�GL���3K�;�;b�Y�΅\����$�M2;d`�߱�os:���x���X���uV��4������k�q�޽���+	��r�K��c���rr��2!|�� �3���z�j�S]ϒ���N2�G�FN��WX�s���c!�@s��$�E�er[���=�D�ǵ�nk��¢p��d��sԪ�fR�N���-v
��P'LkA�1hOB�����U	XXws�N[�|��,�w6��*ŵ�ǧV���KCi��]9o1�#�U�\�����6�1�.AYH.����"S�cwc�v��k��)=�k�\�B�61JHq�k*���yr5ȓ�.rٷ�Y�� ��b��շ��	��$�lkZ֜йa��T�Z��@�/2;7����#3��Ӎ��T�*+�&V&���)�od�M���k_Q�ua�z;���\��G-u9�E(˨q9԰l�Vtr�\
����|^e�(�u���N3���k�%�J�[�`P�:����%m���"pt�ԘX|6፞fS�PC���[BwX2s2%���]�32�뇘��p�04\#n�qĢ�H�ݛ��3F�����b� վ�5*Wv��֍p��)e�N=Tu���I�J=/8�jۼ�د
�n�-�mї��X�ʎ���8: �sOw7f�	�}ӞR<4�txn��mh/l:����=���e�{cy�m<xe51M.Ege�s�]�����v������*���s{�m2iBp������n۩q�����+r!\�w:�G.�x�+0�!t�Ա�˶\�0_ַ��`(fv��XFkF��*`��wQ��.c���PM���78��1�������l�&��/b4�!�)У�U��
�ݫCj ���������!m���-�6�J��{���R�2�'#�-�Xw}S{7��;^������WX�����z��sM.��rc��h"�N�dKv_oj��)�_u()|�wʗ=X�S���P���:���:�c�ݵ�h���(������#�e�51J��e՚b����a�3/��</�D��S:r�����n��o���4��^ui׆M�o2�r�y�3c���|�F)�}iY���T�V��4�C�@I������'b�֎�]V7s��V��*OtIxV�v@��/�\r�t �/ ժ�5r�am<�-�y�O+n�k��� ����jF��V�3uxe������:�]����Lܽ��a|؊�f�����O1�%R��w�x�-;jb��������e�m;���Kw���ע�5�&����5�m:��7K�%'BJl�_Az��C*��f�T�`V����3)��g0A�`U��V[t��A1y&ِ�P��mݢk����͔�gee��8$��xa�
�\N�aܻL_iy�������.�͏�fh�DV�@�.�{m�,l�jmӔ�[ǌ��\������.�"p�	]��z��=���K|�^̈F�q=����f��
�	QS�v��X,Rz���S]�k%�[lʶ�H/a[��0����Ȕzw`�{���#��LF�B: j�7��y��'}[�û��f�l-|���c�����k�eގ��W���T�%dqCX�+�0I��Q��uK���y
���_9U�m�u�E�xz�;�F���,��_�cUG�ZT���"��
xd#7zuś��:2���a0<*ԃ�2L=��jef�ի���p���٤�s;���?���zt]�c�`⹫�^i�vB�n��GC1�kݧ��[��ky�ґjrl���e ��˃(j��iT2�Ŧ�B]��Y�yJN�q"����e�ީ�03{rs,ժ�Z����PTtv��
<WR����W]��{`\�m��>�@�@��G6�A.W*�]03�q����}Y�^�UJBU�Z�:�'��5[��R��uI��|&X�#9�+��M=
���>�����EV	:J]pu(��K���d��٢�ⰴ���
���;G[Y��4�g;������o-�h�3@�xp&'ϧ-�
��lM��v���&d���9)��aa9	$�n�B�Q�wP�B�\�;N�Z�aJ����R�^��+<�.�m�|��(ع�g@:��T�;g2��4gy�"�ww�G�\+ MK�0�K�f�{r�K��+=�w{�7�%��n�N�����YeKU5�83���2r�]�S!3cB�����x�E�H\������ub�c([I��;&��V+T
N��u)Yš@�ﺯ*ۥ�k�u�13�ue�����+���4I��.�ge�c��6�>=�"��!�e"����^��N�����"���	�I��pCq=�}׍�C�ц�7��O^-ڷ�SU��W�5�Fooq�&�uW5J]`��-�*�H%�6�Nd�D
�Rvn@a�K�`]B�2�^�6�
�����n���wvNW�PW��m4$z�h�B���n���y]����{��]wMnn��0���hM�Բ����ta��\�0n��хd�nu	s������>9� ���^��t�Mk��ڂ�9��,n-)	IB�F�z{nw �9��j�*rR�L�E�I��7j!��k�Z��n���hA<�얨ܴ�xaVջE�VXD_vV3@� J�z��S��,���٩�Sͣ��/���[!dW�ܭa�Ud�L'v0����V������Xn	ʕB@�xx,��y�����;+�Ŏn��*Ɔ|��{����.ȼpD:R�IwMz*veAe� ���݆�vjҞA%Ո֢H�gGK�Y	E�)���m�O�go�4�v������tu�[��_:w��f,}9u�����z��p�_<h��k�ŝ;0\i���|�T�N�/(�%�+?[���P��tyQt[����Q����duܸJ����6�z	���5�:�Z�X/V!�_|6�=49�-�f�ɣȱr���ȳ�ݽI�Tvm��e��}�i�=�k����zͪ��N=9��b�2�+�\"8{GVW�+�y�4jw�/ԧƆ[�XD�<�s�\�h�C'����_=��Sl�W��㿉2V�r�+fe�:����orܖB�{D����.I����t�M;���M�]������R]�K*���"f�9��
�ٕe��)�ew�K��k�x��7�T�Q;B�X�):�n��ֲ���V�8�yښ�$xJ���#��^�0��|)�[�,���r�VdJ��׸��sj:�o.-Qbv��B3�
�$�O�.5�@lճC΢�i�=}lr}�J��P�vb9��c�'wTj-)���f3�7��(��ǆ�wGU��F�Uj�v�z�L(����J�!12w`qk=փQ*��Zs{kq�@GNr{�U�M'�l�9��o;���>�ƌ��Z��V�\l���o8J�Ó#��gt0:��Iuu7N\z����(��o(yȩ�q��V��j)��,��㛱�;���׿[�w>�}�|��Ͽ}������ܪ���m\1q�4ˎ�v/W7[b/%��8��y+
Z� �W��g֜��kk^v���)vQ��1>�y|Nu�$�Q���ͭ��&Rf�wIˮW%2���3���r����mԵcE�M����\s8X�ڷ��C�nSn����o*�k���b���v�[oe<tI������Ղ�&�Z��%��ۙ����}���%IۭN\��J��c%|̹��U��T��[��j���pbs����3�u�p��b��[#��ŷ1����6�VV<y��t�y���]>L��fw$G2�;xl�z��_R�QYwR�v��L�����^k�\�I�x򖄮�L�o8P���]	����������ҟP�ұ<�lc'��T3�o&�)ꆷ[�;��z�֝]н�����]��궱�H;Pվ��}l%ӆ^��;;3BXm_9}�3����N�|8�$S8��0���¶��oۆ&)��K� �Xj��E:�.Ԙ������X�4X��G��v���0�X�vNn��Cfl����y�GN��[l1�b���M�|,2�u�$�^q�|\��KN��X)U��bx!˗Q��f�{[�;g��c�#O�y&�&h*WZY�ЇW��9b��X��s`��:.�B�:���F����t�`�跛�w�EQ5(���a�u�%>�{W��$@��ܖ6��	�,�NԲ�֦%l=�b�ɻ��hS�IN�@��hG�c���-�AV�q�}{�Wrê���CG;�C������V�������v��FQz!�����5�д�]J��G�5]��x�5)ܱEf�*�=NToXm����u�Q`E٠2՜���k8r�H�;V���b�k�;��֝{�:���PBV�`��+u��:_lYu��6h �a�֣k��Sy1ҭ\Wk*��<�X}�U��ͻT�oqJ�p5yɻ���h��0q�|%���z�+�;��XdF�������q��HV��M*��}�Q����պ��������X�Ty�;��W�:=k�\�{Kû������X�磫.u3�k�!k�J���s�2f���ө[˨�M����;���^�xZ���ƒ�-<~�M]"*�%۹OR+6���P�)f������*㩝Z��5�{�<%tcu	L$;o��'�-Οf>�2�sX�]�'&Yj펢���zڦ��^K��>�N��L�v_+�;`�,�j���w����1v:',��MT�a��<�\�)a�	���M3k�F�W"�t��2s\K{�ZrvV�A�t�L؈�u��
���tVuO�Dn�p�AM� b'g�ZsP��X�Oe�r���1:6�\�D�jQ�mn��eL�P�])��zu7	ڍt���7lX�͎5�Bt��}��م�_ҕ�u��w���v�9�iNc�o����ҟk��TJ����L��n�5Ӌ.S)m��S8���м�ihg&�i7ר�7�V%��o�:|���"j!�hό�}�sM�U\�5�.���2l�sE��&�E=�W*e[<�k��S�VW�`���Ma�ߴ؊��n]�xE��Fx�)�l�:&G�6�	L���'��n�����vU�h*�)�1^T)l�:����۳W&�<r�#�6/�2�LO�]��5�ob�?&mۚ5fZ.�A�bs8F'b�����:�.y{.PD ��_^m �C���,Z�TSoe�S]���WBt�EGyEk{K��w,��J���t[C����4�b���aa�\s7.��ծlh�M���`>��F�3+���%�@EX�x����;7AÕ��s�{g$��.F]6Ν$ͮ=x�9�\{m�\B�[���n��A�	��j�mԫ-E���(h6�ٹ��ZV��a���q�dV:��{o�6YEP�A��ƍ�r���Y�������|z+8�x���W�Q��uyNżx����9��e��:s��{�;� ΤOWj��:�s��as��Qr��S[�i;v��1�Y��{�6k�6�V�/F�;��=���wkY}�KL�����35g�ϷP}[�K��jUy�;+8�䱇�_Y�H�(��(+nW/�1�b�;�r����ϣ&��%�'Ҹ���D�,�|&V�+сS��W�:�N�E�:�H�plkpdm��KX�)�[�n��\#�e�Գv�q�R����E���jYu���LK6g.�o�|7"���/*ܥعqA��.���;������32��zU��n�a� n����={ �G	��yR����=�.j���[2�f#o�#tuv���쳦��XZ�Vm��7]����i�4�"�/'0x���x9Å���f^F8e&�Aa��k5U�^k����َ	�Z�5����5�1�}pֶ�y�PΔ�3��9Ե�tT����ҕ������̷;�\�+-1Zy\i��K�b�[[��+�Z(�rNc��y+�O*�{(b��6�y�+�=?r������e���)D�pЯ��^c�`�;�r��82\����x@��+6�xm(�]�%��LZ��j�"1�R��J<+�m�4�b�����%o:.Q䚰�B��X�B���V�
ؔ�>�	G6�j�!5Ρ\����܆�*S���� �;�h���/��Wd��w�z�͑l��B�"�їXT!�6~n�g!��q���+k)m��փ�A�6��{[aj��D�6VY���=v��ͰkR�.v���u�@����OX����.�����)�]Z�i�ޜ��>�ԫR�>���%��U�ͽ}W>_l%�<��1��ijgb�2EP�'-rU���v=n�An�m�H��-��t?\�������yQY��޲��@������[���={�1�˅Y��imUS����E�^dϚ��E�ޑ�&�P��Zͫ�K��df|���U�t!��C{Y�hu=;���A�J��*�,��h��YßlY4�Γ&�훬Q���h:���ګ�q��t�]¶m����O�lgX����9�M]kwShWsb5h����!ǯ�E�ær�����t}.�{��.���^]Ѿ9��Mz��]�i����Rħv�hn��I�Y�;I!�}�c��wָ�\38��J��@�u*�o5	n�F
oǀ�@췗����WY���I�*i����!K���9�%�&ծ5o)΄�F���-$��MT�a"]�MO�8��V�+�-Ic�����ȜΖ��%\Z�tos�7Xt�R��n����A��j�����`���Tf�Y�-h����Z�ҥN�]�o�=V����OP��pk���wSi<�¡���A܈���b��v�V�}����姝L\��b�[{���ފ=N,�MЛ2�� S��y�d��I3�5;���z+�	*�����P���'rh�w���A�U��>�Isܝ}}�f��*$�1�mmj5�e(-2l�S޷8��m�����(=/��¶ٵu��0�Ŵ�iP��\1����8�X��޶�]�/h7����v�J�N��k:y��4u��n��������z��m�Ibf�۔����QopΜ���lX�Z]nfŚҙ�>����Z�-�<ܫ��rP���]�ϒ{MLD���W����d�k�8��+gq �o\`Z���c�@��W`�5��H�[ڣ�ׁq�j�\;xnf0e�ڀ3���br�����k8:6esWJ���\/Ry��>.�ilgv�W7g8Ta��趴s�Y��}�]2R[�R���DRT2��h��aٵ@f�Ăl��
9� �ہ�_}Eݦx)u�2�ͺ�Q:s����ֲ|@���X��JAX�{[�Zd[ޖ���k�n]2品�� ���E/�.�b���WD����������f�W�k�U B�T�J����V��f^��|��_$5I3�i]���Gw��W��8{��׺�t8Djۤ0N!_R�����O���{%�Ѕ�ޖ*<�n��1�d���5�(2��H�{���*�[����'��iD���v�nY�{n�\��L'
�aT���G��5�/-�۔��"6��g*��
������rږ&[�X���zs;,7�j��y"x�Co]2S�w���Z9gC�-���gӞ�#P���fSȺ�e
ٚ w�(h�e���je�Q��v�L|��;ڝ�5
j�Yݍ4��d��m�̮�,�^5�mW;�U"�9��p�lD��Mj��gti��\�Wٵ�up���#�N��#3��&kw�ɴN�*�M�:7���)m�e��j�C���� .9m荭�@!�R¢�c�u͇/�|3�ȣ��!�����0�������T?i�x���N���-�o�v��)q��t�'�Q�޳�5�G,�,�W�����;��z˱��	h+W6�ٵF�wC��Q�R�6i�n[�Z9T`�k��1��2�㖦o"��W|�x5n�Τ��L�-��Bf�f�^J�e�nnu5Jb"ɮ+9����3vK�srQxGV���f��zk�{�Q�u+I����7�޳W6�9+���C�S"5�Ø�7o��v��7IV����r���/8*͕�������.���������7;Lĝs�x˾���T���.Qչ�iw�7|:^��ͮ�ܵ�u��t��
�	;e�3z�'��Ͷ4PYF�l�KZ��r���$e�hWW)i����3]�Y찆�v��}ɞ�:�f�d�s�;���g$-��:Ů�Ue�AJ�+nw^6����_<��N��#�֖ZGk{q[�+R���|�|�)�*Z��90�vq�J�H��̥r��uj�osV�2����Nn�����d��}je:Яk��XJ����B7�#*n��x�h�24��fu�\`S���
�h���N�*q�$��ؖ6i^_n�:\e]�6���a;��g�ڂ�m@f̲�˵'3&R�|7��D����'�]+��JN��C�+������X��r����6P[q�qX�#t���P3���=+)ڥ�rs~���]_E:�2����Ӧ��w�š.c�����nn�������j�6I�rA�^eDX6��6�Eu��z�WG��"�Z��`@f��},��/iԡ�*\"߳(��0Y�:\��i�A<Iveu�}��ܧ�R:6�O��[���5s��\�;�IqM��B�\�N�[��v��G�S�WWֽ��E���q�8�ӳ���q�WN_HY���B�h 345�:����\h\�]��Vڊ�C�U�B}���pj���d�>��@��.��"�����{��n�n�#u�ik$��Z�e�kwWAY�ÉvX�utFrm*&!��+Aek���c%p�0:8�[[�b�mKdJ�a�����뫩bڡHv�pwv2�Y�T���&T"p��֍���s�z���V�A��b�Ӊ\���5ɰ��F��P�4���J�i1���W�a��^�f�֕]ת�Ɩw>��6�&�o�֋=����l���`85yݐDDbsB����Y���̜H�"�,���
��q�eP�+2�.�t�<��j������q�z�b�w��Q�WxpC�VL��G����v�-��Z��[��4���  �C)X_=������Y!�p�pU��l��B�F���ˎ�dU٭��`��o�esv���[݉Գu"w�)�]L%ʶ��a8����(���Ж-S흮�����s�d�e�M���n��I�8���x7I-���h���=FN��;���WB(����)Sn�]E�S{�������g%�I<��Wl��E�B;̗�gM�Y�"��3.��g9���A҃�-���u�!Ȭm�hg9O(�\qr꺔UE��͂��,W�1VK��δQ��Q1y��9���-bԈ�O[�+՞����w|V
���ń*�lɸsp��Grv�8�.�m/�`V6��W����eAX�F� �+<'u�L�Hv�(�����x�ej�1Q���ېew�
&�5�]��U�
��h���ϝi2R��R�n�T5�@$k��ۦ��FY�ټI
#ӴG�!��ǝ�=ձ�Cx�¸����"ʙ-V�]ވo�b���:;����Rf	5�B���D7Nc���q��Z����N��Ha.��MA0�8��R�1���[d�6n��I���|��w�s'=��A�o�dsA[�j�7l4(�òAo;i������c;돁˺G�L���n��`K;�M��+k�(6N\��ց�oo$��M�J�AOP�ڀ�7��7�	���Țc�[�;��Wv���Q���N�幘��*��U��K�UL�$e��Ƅ�����慛��a�T���Z0p�Ipvs���_Aԫ&D�� �4d�e���_T�m�>\�(ᾳFCg �$�v��wc5l��zlt;&9�uj�n���X��m���^�en^NBI��{}��+�p���`��0;�ڝ��g��v�K�_G.e�링�6�rکA���iF-l�g�؜�:�V.��1O5�DN�*�n�'(�5���:��h���X�O������,��R�3�'}�yRNZUݷZ�<Қ�gG��]O���ՐSΖ3���җ*G)m޶T�j�^+j���W͆XWK�:n逶:���J�7yx�ƅIK�цby����hV�²��K	Zz��l5�;OD��!gQOC�Wd��u���7yЭ��D�5�S�X�K*��.��� �զ��`��tީ5����k,�H2���V1�T��U���ա��f�.���˘Nv�j�U+zec��ŵ#]��i h�N�n��tC'v2�=x�7�0 �|>}����9��w��rhZn�gBir+hl���3��J
G�Xn�;4#�Gl�k�d�rޓo3S���T�-�(`�רo(�w�:4�Ψ%A��9%�D�����۔�]�[��t��&:+G)�!gT��]n6��:�Jy0$��\�Pa%R�ޤ�ʘ[�eY�{G>����[�t�тY����No�S't�n!Y�|�D̋&�vU�uC@�>��T�T�Xٔ5iZ�J���YH�׎=
P'Z�<�b�f�o'$���s�WN�5v��2��!������ϝ��`���ȹ�v��.�:^�5���K-��q�Y�e�����@s��,�*�H+y�JΠJ�W]HK��j����aK��I�!Nq�sHeY�J8pMK�T��q_w}����r�]]�XSuIt{�]��íƞ��@��+#��+ aV)������Pve�׀�r��Ԡ�y�\���S1�7��̖�Y��&����{b��NT�a�-��ks����]Ψ��5�>��nJ��s����i
�t)G0ո��D�\/q$���5��ԫ7]b���}X}���n�u�`��Y��s6Zhѕ�(hK],�(v���t�fM���-�y�
Y�.�P�%س\��^W*�WMf�ub��Ϯ����D�-}iȸ����Y�;E�7L���^���@r;���]5�IIM�bj�"h(䦀�ht�*Wl%&�IT�T!@P�	�AI�4Q�t�E+A@�4�d+s�ZF�B�JS@�]LE#HP��,MIIl�\%�B�mA%Rkƀ�j��:A�)�P��h1RU5�AE�4����h-:�,s��C����˓���A�9�-�i#m����0����s�w0��y-��9�s�S;	lEK<#�!4UV$�Q�C��F�������.d��;cN��!����5�u�i4�!��F�j�%���jb^A�����:-�����w���w������s�_:=��-&�.�c����l�˨�W��zZꎤu�Egv��Ӌ�Չ1�s�UT[��1���R��Շmv�%�`�׶�P��MG>���.Q.��������+jw��ۣ���l��%^���[�������f���D���v����{��k��}�W�wn�gս����l �����w�O°@ǅ�o�uQ_�U�R��������.R^��$~�P�^�:�{��x��ǔ ��D9mx�CuNРh�{_y���y%3���{|������o�Y����23��L�`�Ez�M<s<��F�Դ���+�=�j��o���ѳo�
˾@W�V.M. J͞���|:W������0w�w���<;S737x��>����b�^u<�8|��hxS��`:��q��
ꀾ��ޟ=�eٯ{�j���e��c>�p@�^oW�3���8j�]C����g*X �������R��Z�d�褡�齮ע �w�L���iq��Ez{%�i�t�mL'ծ��n��)>�,�A@��jP�����#k��|g˹�Y`&�H��;Q���z�v��I3q}ao��7��*stcǧ�ʭ�Q�)bx)u�p�+[���uC�⸤��ˏi""o0XX��z�w0w#�g�9�.��7�}c讳C�X;猅��/!�*��rc�KT�#Nw7+�8�x��zV�Y�5��N�s]�f�ț5:�g~y��j�U�>�:-ز`�p(�z�b勶�v��`=ɪ=����z�='6�{��w��(�l��([��Hױ0��Ů��׆��c�ؖ`jw�o���}�7C�>m�^��7TMh��[��`��zwC��BGq�w4�'R�S�v�����T����aC�:Y֝=�y�9*ù"퇓���cPe�rlf=��;�~�1����c���u��˘R����Ax���j�*yw-Jj�G�A���d�z=����Wު��Z'ּ��ހ9�t@�@v�-p���A��6���[l��@���=��Z��ѫ�5�|b@c�L2C�f3Ψ��}o��-�y�&뭡�u/9z1b�����t�$61�	�4vbh���PP�x��}���míwADU�N����QV����<�'�;~zq!^5j���y`)� ^��J�D������+-�j+!����.��-OD�y��'�,u�oھp�V{���#���� 0N��>���I9o�����"oz����Y� ���{U�+gݙ;o,��!!��Q����ٞ�y�eJ�#�e�U��v���%:F+����,�Ŷ��PX�25��MG���]38N�����u�r.��ي�N�2��yDkFHn����:��� �d9�,�塾9�p5˖�VV�e�5Q�sR'�����&}C�i^�E�[�kJ>@K2��*�䭕V��Jb�xm1�ǶP�&m����S�8Nd�|y�k�D���_X�,#O�{���z�Y�Z�9�r�*A���#g�Ť���|��+ԇ�?q���� M������̃��ԃ�V�}���.�iP�G3cxHfOr�CG�-�iv�_ڐ鼉H{S�b��D���YA,`�����M��M�eפk��m(y{���/�ʼD�o�Y�>Լ,K�/a�*
��r�D�5��@�PqѬ���е]ﳙ�MW^/�T��j�w�o���5ʯ���έ���6�JE��;�%�3t�L�ƫG�8�J$���x�����}{X븺����6�-f��/l|SN�ٛ����%�Xu���n���Y@wh�� �g���]u�n�!D�@})�3��=�F��mLgiHN��T�X6�C�t��=F���zHQ�:�wVuݢ��M��.,Qr���0l3k��5V��Rg�Y0o��5[ގ�Ҽ��aw��a��R��}�oۣ�f_���|Q�fض�� A�$���s
�Gqv��[WO�������\ws�R�1ЛG1P���M��N;�v�v>|�oIA��u��S��WM��:��go!�ه{���|�w���$w�4����)KC͘O�l�^�k˱y��Uhg�RWV>����	�7��b��]���񙞛g�q���ͽ���z��a��O,E՞���W��׃�{���=�V߇���=�ݖ��B=��O��^���~`�ok�'���N�b���rE;�51�m~QeXb"��0\�k�S6j,�w�^t�������+x�3`/���JnKf�o��v�7
7�fXgi�ب�A��1��]�Q 
7+��Z:�Y�P���w_R�����m4�ڡ��3F�w���0�Ap����ʱ{�(�p�hm{p]Hع]�r`f���~�o��?y<>�*����0�+r��ύ�XH���q�jڂ(�EZ%m��q$Nڙ�حG��8�Z^��Hpɇ�=�=�X.SR�5>><h�����I�^���52g���:崌�|�Գʺ���|s��ƏC�jwbr����F��`d��Ӻt�!��)��������X��c��֓r�ϭyʄ#�&׈|�l�inQ�|U�v+���t���5��N�Z��,|�>/�]�8u�\�,��]�8d\ձ`��4K�ݓ���jG��SoFa��ʔ�讅N�u����q�Ӳ��.��e:��ų5d�V%���_.�����2m����]��}(obʹ���=9��z	����tc�gZ����|��]���ж��w�D
��;_��ͷ2g�M�!�`����[J�C^�3�6;S�.ƙ� ��x$P`]�A���b��׶{�h?]�o�a������%Z��2|e�|C^��N��k��WT���mn�����{�.�1f�[�l�m��i
���>J47P���#�:�,�	��1U����IUv��א�:�2Q��T����©C�]�auS�R����O�L�]��u	O^+f�4j$ضT}�G����oH?W*��F�:�*�ܔW�-�ds�x��a�2�Վ���MӾݴ�0�I���A�W�v��yj�3�6�T�6 ^�~g���+�ǅ��v�᛽�y�WN䅫X�s��}	��:����a�,�5�0QS8���ơ���k�j^kW���X3�/g�'Gijr���,��[K��b�]���νo{Y�=����)�l���k�w��Y���:�QEaiŔ�/������<'�²�� +�x�O�7�<����G�)+3]�V����8)�9گ��0 ֻ�B��p\[��X~�r阅�q�Zxq�۷�pX��y{�ye�D:̋Bw3,')���#�OC�h\	�qf����@aoj$,�����5JorM]N;P����3d ��R�om��������i푨�r�{~^czU�F�u��
������4<)����^h�~Ǉ\A��3��ɖ+���x_١|��C�����U�<1�}'��j�\>��e8]y������0�H�2��	�8A���i�;f	d`�<��5�o�������n���]�Z\}85ݣu��d#�+!�O�]`�
D��e[NY�����h;.�I@{�:�'}M��罢�^���\��q	�a��:-휲���Z*ϧ�)�]��i4.�,6���������@u���MW �<����S}�~�hy���heq��Yv���Hr������z���AW���q�<�p��y�[��Q�w�鿽��B�(L�b��9E��w���(:���+���)U
�؛��;��7�=�'ؾ�U���K/��\[��ԉ0Ӂۭp�Uo����DJ�<|�Z���~)X�����TvR�Uc��z�ܟ+2<�-�N�N�EC�j�hMJY�֪��k�\�#�A�@�{��&��k�s;���݇8R��o�R�K���yZ�5��k��>�d[m+�9�˝��*s��VHz�\U
��vVd�P��R��]���#��jViHiע�B��KV�_%���u�#Z�z���D����u�s>����釨���>�ʭ�K$�jwV�*���ֺM�(A�����:{��ye:ePd���f&��ա��t�`�5���K�`@�|���oa�)�9�ݙu���V6�P�<�V���O�e{����=���^޾�����{yu��&	�g�7	�W�\����n�|bKȿP��3������U�/,l��wk�%8��Qho�S�z8%���X�ʿ/�����mf= *�Vr���:/�}��fvJ�~�7��'��"í�8i� 6̯��-䭳�q
�Ằ�ү�$Z�ݾ�M*��ˡ��F!��׋G)�
v��nC���= ��D�4l�/���6�x+ܭ/QfC�[�f�ת˃�P��vs��Z0R���ڵX��yv����8�H���v�~���įL�K���R
�$<Q���T�8�[A�U&3_#s0��<W��=9�*���SN$���Sɋ�5D�~�V��b�ըX��ؒ�2�^�Fw0kW��m��<ć�V��e���U�)}(���<�Ǯ�}�Vz�t�ʗ�d��B�?��Y��X� Q2�wY��/)��Պ�dA@�ҕ߾�x}��t��rp���v�{ڮ��vq�:_n*�ٶ����o��X����X������;�ڹc��e���,���\���ޭ�\��]�B,G��"z�f"��s܅5]˵,Ƶf������2�=���C甯���5�~���� w-�\ �>N���\[���\D0Sl��;e�j�j�Nd�fl�	��q�W�l��c�:���Ǝ��T��<�MԴ�<�^�ձ<+m@|�o�uץRX<W��h��l��43��f��J�
:Ia����97Dy�y�$�;kM ��ۻ�b��C��PΪ8���ޒ���� ,�sܪa*��zb���n�%��kI�Oq����aTUG<~���G�b�
v]6�Z�K��M1�s���ho���@�����?F����ʫ�U�=r�"8�C�V�1i�:������jCM?%���������5�7۵R����8Z_�K	��Y9���\`���>�v=|q�}��?%[|�z���~Ӌ^k�N���pm\z����@/�Փ���DZ�D`�b���svT
W뻖A��׍��q�<�����{ϘB�6>�C5M>u����j1�%$��f�(e��ý�0(m�V��@�	W���W��Q��n�]��J��b��R��f1��n���1U�X�t��|�Ï�ɚ��Q*�{x�:s�w��C�=��r�f��Ql�@�(�S1��_w�0�[�,�Պԓp�Бu7�J�|sP��3*Z�vV4=�����^�^vW{�z=SVK����ő���QyD�U��笁[u���agD&�rυs�Hp�U���*�=�-�4�������{�G��h�����u��6���A8�+�*��e��Y�!>�m�=7t�˘��&�Z���	%0�m��צ��i%eK���H��B�U}��W��k؝�4��_4���⭲���^0v�Һ��{:�G����lq}������e������M+�m�y���y<�'�h6��P���8iTHmLc���ky�P��>^�[�����3n;�ܥ�iC=']o�2�|��X�a��5�d�{_]!�R��b�Lm�P���H����r+/|Ч ���]�*�b��hn����
!��c�'�|���ի�Z^�£�ݽ�z�.�u�LUm�2�����+zk��z�5y]u�������4��{s���<&K�¶���#w���]ľ�e}�9�G:�x����|6#��tl�AJ�%G$9V��F��B��ciy}���:U���J�@/��[�S9t�Vޢb�g��{n�t*��L���k9�c;tk���;�4����:;1'�%u�3s���+��)��y���9[h�}����R.Ky�e�U7���1BDo{��f��5Õ�����*�jƻ*��"�T��Wݙάzv��Z�lZ00����wq�T�Q��ӳ{tt���J�6ZOy�׫��0�D/T'�-�9�j�t0A����Xew���h1���]y�i�7�pOS"�Kڎ�§���{�M�G
w���o�_f�]x_����.6��Zaw��?�z5�C�}w}����(
��J:���p�O��f�
�V.j��	�YI��l�U}8�6��-�:�'s�=�a؞��o�6rR_0���yc84~u��)e�����[s�X�aV++4���fD��m
g]���'��܂2���ê��3S��=C4���g��Z|ٽ���z���5���mw�=��� p���u(�:���2��%�fZ���a�������1^��^`�P�-*ݶr�g#k�%��<xU��=%m��KcVon����zs��+2����c'����Hp��>5H�t���r�L��D�r�ب�x�3�7V�j� ���w�>���xNש��,l������63�x`��!*PG�γY��)�w]˪���r���=X���R�_e��k�C��]>��%��E��9Xt�D��4 t��t(�Əa㹽A�۫�R]@p��u��E���$'��dA۸���9���kk���h���{�T%m��R�}u*uvo9k���(\��:M�{�!��Vb�=����ہwtX�֭m�&�P5�W�鲕M�tKH���w�9��9@�n�F� 6�uR�n��^k�M�����9���7:��
gOY�:E�{U�u�s���`�L��������@����_t��&6Y�Guَ��D���G��{�o��a�ɔիq�)���(�e�y3��oQn���]��uvM����p�����yݚ+:>)Z}�t�[2�n��lI���:�ݛ"��L�y�ܕ9][��.���4��ʯS�F4b�,�a��)gTwS)l�BM�N�����:��w������fۧ��9K+�u�m��W\!*����
�9`�0��w-T�5���dC\��p
䨖�D�b �.��V�ּ*Wu�#8��$���!؆�%w�����|h�m�ƶ�۷b�Ŷ��܍�I3�}q=!�Z9�z4���ʁ�z��rʺ�Í(��T��iЭ�Z�ќ9e�˘��<�e�V;!1��>Д������o�>�v�q�i�pb(d�lm��fC�0jnec�ǵ����m�+5�[Uř]&�����hK��t��P�eٝ�`��\x�|'T�H�{X�w����\z�`���qta�� h�o���U��F�m]�L�;�U��Yt�uB�B���E����>�V�Į	$��7�����>Y�zwnV|��ޗ�+	�|�h������nt'�+Вk/����ѓ����2���78�-��a�O)�ST�2���$�r*Avb��f�{�՘�ŵz��z�Zti�${�P��n�o .�9�Ñ*vtu�����3ϥ�[&��&�Yj���Ya���;���LB��%3_x]ݤy���Ե��2GFQ��]���RX*��h7ܒZj�m-��C��*ֳh
H�qԯ��t�/�5�V`�S�B�Z�׃5���H��9Ʈ���D�U�O;����Y9���U1�I���S�7ifcN��̗w+_'��̑7'-U����S�eH�9���2��r�f;���uv�r�HS�X��F`�i�r��ν��m�zw�ŉ�R,��R���e��^Ar���U	�v��vܙ�<;[[Y���cy���N/�5Ǵ��ڵ�����ڻV�d���s������L�b����:�SM��qL�v{�8YzJe��.�����i���U�/u�Y��1O+:���n�TC�]+�\`6gV��Pܥ�fcM�ʱN]J=t:J	������Q�� ��,Z�����YZ�E8����]wcr7\M6oE��ݦ���'7��޴��&�bw�|�����uf,�D���5�K��r*m�zi����od#�����g~I�H��Um��Si1!��O4P:Ӊ�PD�MP�����j4O*8ZX�����i��h)-PV��Mr�<�4E�4P�J��d�M�#�3�"t��&���\$�r�r�i�1�"65N��5m�Z3RSF*UUSF$sE$Z4�e�d�Q�4i�F���M�DZ��T�iӈ4r���Ƃ-1Ql��jڍ�Z4�5��Ӌs\��LQ������g����A��[m�նv6�T61��TU$N'�+E�X2Pm�������[b65i�!�-��DV�m�ch��75hh4��C\����AT������%[.��� RH�I�$���C[yr��}����8��B��}EI�`3Q[��b��R��{A��0�Uc�t{IwMΘA�������L}Φs����u�]����G����	Tt�\\C��y�^�+A�=G��w�i-w�>ϐw�4�xyP}�G�z���_�}��[����ѣ���<����?���AvO��@�z�z\׌R��oL���|��4>���]�~ﯲ�R�����O.�P����'#K��T�|��z�����N��4���#�<�q�}������$�r +���%�گ?�5��d��ʾ�=��u�����=�_�xu��pS��%���z����_a���)�.���߾����~��k�YA����=���9~�ޞq��%�=s$�!I�]�p{������c�Á��(ؑt�����r{����<�u>C����� ��<���|�H|���w��r������w.�?���=BR��<��:??u��G�y����ާfd���=�|����#�*�	�<�o��]-4|��ʐ���_d�/q�������|�!)�'p�̾�����κB!��<�K��/W�
�y�羃�C����|���'f`��n�P�d����ًv�_34��5ɣ�x�����A�=>��O�t����u�:��@Pz�~�RhA�%�>p�{�A�������%>y���iuC���:�B�����[*9f�)'fb.���n���MO�K�Hk����O �ܟ��r}a�����#�X:������Q�BW���PS�̼�����? �˨;�4%'�o�y���h���Ɵ�O<<��t'vS�jm�c��E���ﯿ����]K����t%���}�'������9�a�ܟ<�����~G����)����<���O��z������'�rwP|>jvf.�������)�u	Vi������BPy�ﮟ���:{<�p��e��p��h�~���^�?%�z?d�i~\�z9���k�c�=�9�u�>���ǨJ~ϯx:�/s��S��q�m~�t�)��ُo���"�����!��h=�����P4���->��9%�y�;���h��箃��+�=u��?!���z���:�������=þm���N���<��[;��Eɪ�䆹�<�0�[U�r���@Uj�^�st�j�vG2�r�_[���T+YS�U 	���u�mj�]�\�E�-;}���sN�ɝzPX�F����P{eܰ�GI�+;7�ufwN]7�=�c���������n��|��ԇ ����X��J����z�.���^BW�z��ޏ��O�k��n�����������B��}�A���}p����q�G�9!��κ��fw�t��v3z��BQ�^�2��[;hz����:����Op���M��g��O�|��z>`9+�_x~��/o��O�~����g���>K���^�󴮻���=s7W�'M"������ߖǚ:���s�^�����z{�p�K������C�J;������;}n���k�y'��xz���<��7��K�ܺ}����nC�篾�uκ��`\�coN�4;y;0|{�������u��|�{��S��y����t=?z�u	��Ǯ�	^�+GQ�>�����O.���?e��=BR}��[a�ٱ٩���m�6q3S�\Q�{���<{��Op�<~��GP}�_#��ϼ=BP|�~��Bu�i��ﾗ��pNA�=�:O��9�O�tiuZCBWS��c�|�\���f��7;C����s<C �=:.���+6�~������߼�J���O����%�y�_$�S��<��4rPh�{���}BS�z?y��9����é4���!��3C�>A�9|�^��K�_��5��r-ٳ(n�U�y��޼u���C�j�o2��^��9�?\��}���%?���\>Z ���:���h���ur_q�?^|�������ﾞ���<��y�KOS2v�o,�y\ѩ�̒�W�ٵ��A�q�<{�����=�è����]zy��|����e���I���#��CO����w~�ט���뮏r��y<���@QC�����}BWP�kזO.�r<����<�����<~w��S�|���}�Y:����<��9	z�'u=C��y?GPy�GȤ�%p{���&�����K߭�'y�C��<�]C�~�[�bE�,���`�/�`��5mK�y�����I�u��&�>�����}�I�=�oQ�%?��>��|��J:�y=A�:��w�'/�h+���!��q`�ƚ?}�|	�r���\��έ_��!��v�tqslon��GE����������G��_����U��Y_{�J��P�a�P^��w��j�_�����Z�L뙻��^�-�r�����������b^���X��獛+�_ns¨s�2ov��R 1UZ=���w&�_~���r��z�������S��y�6_�ʓ��\���/���uz��y'ˑ����;�����O�p�����hy��[���m��/q�NM�w��f�n����OPcI��:����<��cK��p��:��pk��~�Γ�����<��_��Rvy��(�/����q
�k��z��w{��~�r���kBꇴ�_Z�t�f����/�o���]�/'���*B �ϼ;��P��>߿�uw��@h����!���?`�|޸��g�=t��Pz���>��9*p��7 Ѡ��t������x�p8+�k��G|ۛ;���	A�;��6���>>�S�]��!�����`>^]A�����]N�}���*��>��W�|�#�>I�_<�u�?G$���~ǨJz�|�ǐ�����|&����m����ә���+���t�pr|�/\à��������Q�9^��%z=`�'Uy�����i5��O����: �}���Hi���y�����pz��G���RU�p��fj�Ý�r�f~����޽C�y��ѽ��:�?��y̜�{���Y���� �u' >Ɵa�I�����z����:���1�=A����~|������އ����>Ď��P��5�)�'V�h�N�O���P�{����wR>��~y��w|��}���Cݥ��:��n���.����7P�HDq��������Z��@v��RZ~��٣�۳x>t�[fyv�>2{k9�ٛ�J�Ϝ��M`�!��/�y'*~A��8w�h>C�G���}��%���}#�������A��]�����;��:t���Q����.��������ޑ���;���^��5
�C���>Ǩ�O�b䆃�#����?��z���{6?OP~�@w���5C��>G�9���Bui4�w�;_P�C���Q�케��|:�K�����<����`�`�G�ț��#�n����boz���=ǝc�w~�ӡ�������NU߬!���O�׹��}����?��r���P��G�{���N��s��W�}>s�Gpyu"U�F�O߹��Z;&�؅&:�RK�&�z�ae�r�;c�y���ce��Xa6����5�KyN_��C3�z��P�oס��rN��_R�c��ϸoV�g/�[Jr��"�A>�B.\�a��.wW�ňY����!���B:λ�{!G�����n'�l�Q����׋����C���^K�uO��C����:��%������_�����8[���3�n׉��1��,��y��&Ψ��'��>�r�����c��=��<��2e�"�Z&40}�Y����H��7���\�K�1�3��%�U�0�̺A�(U/j�- ;��[�]�+֑������c��+N�t��{'f�L�v�5��|B�w�~h�U�6|W�-�O2<�F�el����k�,�='w14�)�V�*�����}^�0=���\}���뺉�V
�˗��fo70CA��|2:}K�1���/�	�Dc��bhW��0A��-Q�כ��ȓ�<(�(�l�|{e_�s^N��g���V�`w���p���^�e�:�-8�w�����K�_njkh�c���f�j��^�ف
�n������P�+����0��"y�o���E���M���p{��sݸ�%e�Y��˵��1� �u�~6P�϶]wg�羻���� f}&zs7tX(-}���<v^Z��q���ۮؘ�u�Z��E/�1�t=��]��9����Uثt�Nn
[C��ʀV�X���w)=��K�[�P�u�A��/�����ެ��Y����ڛ��U�KM�x�=s����<�J�=[W��(c;Sms6Sz��r���p��L�J8$�Ƥ�m=��R��J�ve>��o\���ݙЪ��-�yt�[����^#離=�jwu��KNV��+��K���� ��>��������-Q�C�`V
�Z�6<�����x쯽�Ƅ�����Ӝ6[Ɛ۠��<���>���*k8�О�#]V��{l	��	Սh$ן3D9�gB�����շn�x�I�L�0;o���5\ zwǞ���'�c�����hX2E�O�M4�V	��
K;�[SG�Z}3�H�&ڤ|tT�φ�Ǯ[�ثeԦ�ݤxZ���/��W�7,-/��؇��x"�X�QLo?
�q�[3n��P���{��An��;j���Qǖ4�a�M�Ҥ=�z4���\H�!��4}���w��v�R�7tE�8$f ؝(׫��������>�dBy* ]j�;N��mj�)���ܵݱX�n�Y�Օ8�l�ܶ��5�UL5!䁁,���˼e�ƽ�t]N�F�,��Tk6E��mW�����V:G��� � (d�:E��Å�&�@��k�;��y��KD��X�x+�Ā���q�;���f�ȶ[�~TTI5�!�Ŕ�a�Eg
�����&�lt�a��ZI��42���\��)|9�/���m4PB�]��:�k6cw��\��r�IlWlg!�,y�ܫ2�F��;>+� �X��~�����ꢻ5��U�/9`)��યy������	�t����}�"�a9�Hx:���<d�gNJX�߭}�-X��6��Gp��¬�1��ޝ� �G�����J��zD��ya�4�>B��Y֍-f�J��\y9a�:�*YҞ��"�F9g��T�45CF4����zl�0V��3���c�7Mn�B����.w9�=G5�Vc�Q~�b������%s��2)��w�?G�@,���R���7v��c��L�nm���/�<�Dc\B�oL��f�C�fu
� )�.Y�So��T�(vÝ]=�7���8���*��3�<2Ү�\7غ�xX�+Q߉����p�c��GQ'*�)0_+�n��ߜ[�l��IS��씾�rT��=�}�$��+������̩��k�U��۪������������GҘK��/�_u)(��W��һ�<Ը�V��Z����؋�-�MnO�J�E�(wl"�<[�2�4^�}���e�E�`(�W��n�-��e�AH��H���+��Kzλ���S��O��r�^ �)�E��]7��%ea|r�R+��.�c�����i3��#���ǝ��]geD�"��=�7�'�7F�ъ&�A�Em�f��ħApw�3��M�$���p! o����<�;�е;i�q|��Q�����wMp�V�1�`>ԥ���Ȍ�mT�����K.2��U{�q���ۖ�ݔi߂x.�VЇ��=@O.q�>߅y��`Ӫ}�U]���5=d�����Ef�-�\���/��h�ǚa ����|�3.��+¼2����n+��������qxy�������ѷ�c���E���FAz|Q�IZxQ��X�K���ȩt�����L���/h[8��EH!��y��^d���P/I�k��I+Dj2��\j�V��}�����H��x@��ݏ]Wj��5/�Exh[-�xZ.ܶr��#���n�i�_�f�T)��t�w(����zJ��� o���%������S�o��7=��h�κ�8�PH=���]��3Nl���YA"q#Mc�zh ����F��w�	��v���"�'g���|�����M��S�|�jmZ��Ap���{7ɉ����#./�C�>F�!�mϳ+����}G1x^˺����k�z�׵c�P͔ۢc�7j�oC;כ��]_ws��0��V��G�%�ҧ�Hc�IJ����C�ڝ`�ʻ��.�˙����jy�o�Qמ=L��]SU>b�:S�}kh�1�S�Q�T���_:!�j���t�V� ��\'�L}�!Ԓ̭#��!Y[Y��֦�wy֌���6��X�iZ3{X|�PB;>O���T�
��Q�|4�Ə'�=!�/�,ٟN��1PPm�	����c͓$Vߑ��O@�V̀R^	�_���V����W�b��B��=�5o0��xf�yxPޞ�en'�o��L JU��a�a�֚�OG�r�y�j�K��/�5uFU�6��L��nQ�T�v3a��~����oe����|G*F�[�n�*��\5�s�����{fM��at7�Z̆'�\�Vca�%�Ј�`�\�L� c��{M\�{o	��Kl�>�|��%��l�٪\�q��w3�wm,�#C2A�Y���ꦅI���dׅ�z��<&�E���j�P��I��i�]1[4��o`ʮ�����@%\6�_p�JC����x��kZYZ������P*�Ы۽����s�n��
[�����uQ�
��^�,#Sޠo[����9y̏bj��'� ��]cB�t0A�"�+ڦq�{�n�lm4�E���Pb�[�Ӯ��3o;�ݫd�x���0�;�^��p�s��F8RxF*m'��vݧ}������"�O��uQ���*	Lymjk{(Bit4El�e�*����/C^_S�3���I��I<V뻨n8s����ӑ�dy����7���gx��a π��=9ڊǅ:�,?�' �6z���c�{�~37}c?[���CI����7N�+�wI�j��ٟ+E�V냇�xJ�|�(��.�S��51� �!�6mߺ֒o�2,��=�o6�ͫ�S�E���Z��(p��Y��A]矧�'<Ỻ����t�~_�]e?y{i�ϲw�D�c�&e��Z�Í�X}Z7��!C�lc=��
/ZkF�©K!��_�;f	f*�ױdƊf��p� ٱ}PVyoӷ��W^oxf��Εҭ,??��391ПY�*a�T6���CT�T΂����7>��woڽ`��v�Q%�)��轧��#]V��
|t�f
*�W��2��VwqZ�*}+��QiT(�˹�f�`3\ Zwǟ}X�R~V8O�vϊ��1>�mhtl��21%,&�+d�`"r�(��ԗ��06�s�[=K�j�W�d��+U	\4�����[/�D�",x.(]w����
��KJ��{f��"���{�h���]C�{��[V3�%�v�%oJ˵�y�z�҈���D��7���J���:���;ؿ\�]ɾ��1���Z�z�E��]#���ώ��G��4�3�K|:_G�����6���S��s:�u �g;Qg=�ط%_�'�}U[�%��$_�	Z2�m��i��em�[�u����>�ƃ�&<Ȝ���ô�~�>{�.�*����_ɦ�v���P�(ש���J>SO����dA��t@������1ڈ__����%@n�(�S������0�e��b[D��Nʥ@��&cY��l}0�Dl�XQ���af���>G���h����n�s����'�ݚ�^��
��*��Ä�4bզa�21�OS�K�m�e0��jQ�n+�]-W��倧J�xEd�a��J������.�f���-̨���K��	��͝9:�7�_eT�c�=��F��y��;�۽���| ��x_��׀��|=v�� ��#����GY���ݝ����)�; �>�=�X9�_ܼ�Ϧb��.[���3�[c�-�{^���5�������r���X��Gu�ҭ,�S<�uX�z�O�X+;��"+���(~Ѹqb����g��O;�m��_3
��(�9�O��.^}QE���؇��)S,/�s��X�ۈ0߬��[�t�StdnB\���'1�O�u���;>�24��f��׵vh�۪$��v�SH����,�lK�}��Ɇ�gQ�d|�ԼJ�x��cB��AKȹ*B�r�
C�ǹ}�MJ#�Ln��olc������p	��q��F��4����nZ p��Y[g�J�[�
&г^s��kZt.	ܠ����`���Y'gr�=[���b�t�Z��}���?�*�,N��)恎\5��v�&��֙ݧc�|�+��;�k]�����5N��V�V�]g�mfK���YYE�Zv��Y��K@Kկ�.HWn���y ��m�q�{�J郵V3��^�:�v�q�U7c���T�I;+EF;f�So,�mu%�'U
�w�k��^.�
P���x�:6�<�ǃV��ݲ�蕣��2Rj�̻�(�b��γն���--��,�F�L�g��Q��<��:��=�Oh�8(��=�3(aLd��R�P�����1�Ռ���V�ʽx`�\';y���n�!Sa�5��W��=�tmz뻭#�+��i˒�역fФV�40%	� n��d�75LLZM�	��-��'A���J�|������!m��1�Y+z���S�U������p��$30��h5�ud�uV�{���필 ��3|h����T^ݾ�q�eU��+��+C�!GEZ̮)Q㴊�˴�[Ϣ�+�����г���Ʒ��;���U��(>W§m*�h�=�p񏾃cT��ef�!APN�J��߆|,�<�3�u��׆��q��+�jV�ήCqR�)�n�";���[[j�}eV4م_ҙ�&��pQ�9�}� �
���V�hD�R�Ts0�P�J)�y�cS�Ecx�J����Y�V)|z�����A�U���ݠM���Z�%�Yc4��pW��*��f�EL@��N��픶5¢w+oGn�3S�ɽs4�C�(.Q��H<Y�R���Cnro�#�h���n�YV���^e��a[R=:��SK7����9��ރ��c�(5�S�������/D�ƻ(l�co7
�OH�1�]�]^nfc����op�F4���=���$.��W<c���4�B�U���V}r��ۮ�5�:Bs��\5����ng�݄�M�]�����p��9�d�闲�uJ��7n�z���Cf]v<.����z�w{����n�FX������N�[�zv�W	B�,`���z�gW�6�hx�w\�uZgȹ�(u�]pV%����6�un�����f���y��v�J��H����&��y4��8�J�u'e�c��P-��j�j�s�װ��oq�z*!���i�t�{��Bo�.�Jq*I�Uwi ��t^��촥���rr%��r��JJ�ѵ%��ws�ȝd���G�ȗ��G;�!��υ��|@E������4�UA�rLM\�MbK��8�"���5MThj��i�Zh�-<�E��ӫgF�766�Q1E��Z�UUC�mlQ�9rڵsb�����t�Mi�'Y�6��$�q`�1*4�լP@Si6��劶ճ������`�9�Ik�U�����mȒ9��٤���E%EEm���*Ջj����R:uN+j*�q�p�0T�ns�RL����m���si���ZF����F��s̓G#��IE%Vى"�l��U[i�J�Zc�5G�X�3�h����h��E1QVΎFfNZ(��\�.hֶ��c���4���779����mÜ��9�#s�A"R ���;Cw�w5X�'�Ӗmr��1w%��. �w�|v��Y	��-n[�u���#�[Bj����?{����S7XY+:p|̌�W=�����puƧQ���Ǆ�J�:�p�]c�<-v�ew
�&�z2���}u�*V��N���c�ۋ}���R$�1�f9M�q�&]� �
�j(��
��n,����U��kՖ�3/�l�/[��ǡ w'���8Ԫ��l��y��xLr{7��8s_=�qu7�Wzw� +<e�v'����b�k�0h��{O�(����Z��i�|�
���5*�p�-{K�����>�{*]u��GO4r�_���i~����G��z��++׵B��Y4Z���Oo@��lv.��6��e*��@����BY�SP�f������9s|%��ꡑ��y3�����_Z��I�:A�_/aˠx[:<+��C�ր�ֽ��黇�N����ˏ(^ݹ��{��an��s+Xo���C���vv��+(i�N�y{u��'�r�K��wJ�b7B����5>'�rQP{M����m�v�iU�-���K9U��EUZ��#����4Vy�_�q�b���7L�33ˮ�	�Z���l8�n�{����T���:�9�_���Ly(;N)xd�ܮW�lT�6�� ��$tj^܀�b���f��V����l�g>�2��в�w9�I�!�zwh;z��]nh�1�\W�m�
��׻#�IҲ���F�<ܺ���y&'�f�����-�pJmv��kɷ62.;���*\@�������x�����宫��VT`�! z0��\�r��n쐨�4��H-�|.U���+��嵧��D�8<��įv�
���^g^�IRzϟ���U�	 �O���ۂ�CY]g
vxO�ʘu|����d�rpk��Q��l�17a�Nl��t_oL�<��,;H��䫴����ߌ��{g���s�����Ԝ���ysg'l&Z����T��^�`����m�k���vRQy�]W��uf	� Y����F��Z\5u��0�
����&�޾3���bs�O��[w+7Ƴ�[�＂�<?��%�qߚjY��7xO�䱭�+�0������5c<v]��zߜy�&Ox	=�t��yc[~�=�mV�]ϣd��F�!��`����u*H2c�vn�]xy�+&��J��;e����<!���@U���T���<���p������v;3v�N�t�v��=�
����hDW�s��&п���X��T>��]�C����w<$���	��#�.w���BAzg��e[5c9kF���ܑ��6X��;{�
ÅcRe#7�$� hwf������\���D��գ��=R��Y�V���ufs7�IH�d
uL��M��kv']R�������37�#bS�h��λW�+��'`s���Ʃ���-���f�K�@c�~zrߣ�i��k�<�'�T��T�^)	NVĠX+��iw}�*��Z���%%\7�����h]b�g\�1����Y#�<Z���m��� ��������i��v�� �r�sM�+���y�=o�ם�:�1Z=�c�o�:���Uk���߷�?�MOu��5�o���Qs��~�����������;�����5�5>8�2Q����ǅ?��N���Ҽ3�˪��60�b��R�ų*���p��i��vE���0h��V����XV]U���p�v�*����'d���	�.�ͱne�]x<�J�Y��cd
�ہk�lں���쮨VŅ�<�Wrzf� ��= R�o�o���zh�[��!/�_Ϻ�×��a�t���f�����q&��1�j`���>;���Z�<wpELtW�/o6�c�_`V�*R�����Q|�߷���S~W�:WKKΠe�+�b\�+T1�T5�����h�ܹVn���K��/Z���fjK����~^��n�锵D=|�	\��)0�01��n�`"��;Θ�skK�e$���l]̢-]	̒6���v���'y;�n1�>Mv�aܷiŢ�+a����R����o*ls8�v�%k���nJ���������	࿫�o{�ЬZW�kx�3�?3.�EAv Mf���߭-�:}Ҩ�i�x������`�W����F:��c�E^ϧ�h�}�~�V�0;m�5\ _=�F'v�Qn_��YDj(�Nl4n�lT�E�z�VF��Wk+�|�֪c�5H�	0f�#�T��A�i�}l����ޓ���i���R��l�k��V�������uƺ�Vv��1��u��B��X���緛k!x��V?�<�]:���X�z��z�C���e�/Yl�V��:%�5�6��ק�� �I�ј,bt�^���'����Eܟp�;j�ܽw��6��v�R�My�nQڨ��Q�<��g��e��{�ؐ�*B�,�Mm3*}�%jXL�=�X�w�bnT���6���v��C��	�]���V��J���2�Wlk(6ow��"3&����п�aw��8���k�fC]���^rv2�G7t��Zr�ֆw{��ը6���6�D�*�q�y��9Y?hGL�GM���"�߽�Ť�[�چ��+{;���1秭Xޗ�ҭͮ�"���-���2�D�T������`��.�׊]��o�ܫ�F���yͽ��*ȫ���Eg
L�)�Pᐎ����n��V��d#�\�±�חNIIGjj��I���yL9ǫ�O������5m��y��fi�j�-�q�L/�`�2+�$��ߴ̲w�[)�3��ؕ�,%tG:>@m���}]C�Ts��Q�3��Y��k��X���O���: ��7^��C���JyX����,K����`���¥����S!�y�c��ҭ,�Y�a�U��-�.�ütX֍A��^+�Et�gM����rB	�d���q��2��T��2�/i�$^g?x���W��dZV��0�d�'&��2tS@�tVE��]����58�I��x�߭*��%�}L�8�Q�| �?�m����4t{�K�Y�_��׏���k�����<f�Tz���w{�����l�'Rl��߽�4;��~���tc���]Y�o�z���u��\z�$���pj﫺��ђ��c����~��k�m��*I����N=\�.��C����*a}��}�=������9A/i�A��ahܽƆ:�,�Cc�zY�1�!E���(԰�2��u���wM�L'�T��4pu����W��ym���yV�2�=����,Ю�>ņ��D��5�˚˨��XfQ���=
n�@B�;:�e� gק0��%��b�z��U��o$E����r���
m>��!��<y�u'�ʕ�P&��gu�4�a`�S������Ɓ���ih��g����w�f�����l=��W�U�y��K�r�i"��C1�򻦉7���㆏�Z�4��:A�W��2�.�7p�#K�K"61!:r�[����ϴ�ypB���>�]'��m��;xv����>��,s�!�},L�҇�y�/��>��X�A�оo�0�����Bx�6@U��<i᷅A�>���jo��Rt(�M��)]Y]�F�x�j�wlyQ	�11B�|���t�����:�7~�ݾǖ'��Kv:U�x�):�U���ݥg���Pah�V�O�^�ִχ3ܰ�y�&�:�4[V�\�^�+��僅ûU�S�}=�`��Q� C�E���VF[j�3yܬ���:�����C�a�戫�\���_�0��ɲLy�&�&����r� ˊ�׷�FϪyry�p���۔���T��b�V�{�O6bQ����+�~�۷-����O�^�kW�\U�g��O=�ʦ��CF���^m{s��V��*��{��^=���<H�.�\7���:���gyw�m�?����i
�Zo��[wY2��xv����>�gf��l�avJ3%�5��Ziq�8����t�I�Mn��8K<%��Ṛ��b��:c}t;������S=��z��n��x�;���-P�.���}6�Z0�]��:�������jPkf=�.�J���9t4VTh����o31�3��R�r���=uI��.�Hw���u�㫗a�;�t[ ��I�e�+��)6N�lz���|�,���!PO�����1�K��p�T�\��W������A����F^3 cm7+Iӄ�[���Q&{��w��Y$l���l�5���p�1�ܥ؎ά����,�c���K��a6�k�!��
Cv		�a�M4ɑ@`� v���\K�Ր�*ӛ��Λ�H�-=K��T��]�t�ٗHxU{������Ъ��rHѵc� ���<������
��cj]OX��ɤ,��(�kwrʡ��)�p�n�]�=u5C|<w�ȇ���<�Tzr9��;����v3�*��3$e�~R�����]BL�[�Q���l�m��'�X%<-�-��/aO��
M�F�Ex�:Y-i�!ۧ��7��km��J������ O�N���@ZE�}���:�ǅ:�,:��f�J�r��Ol�_��Icb���}��y���r�}mY�� �̠�h���=��@a���E+w:�T�_c���Y�R��,��=�޳;([�<�c��JwKr���`R�*�ڍ�}�ά���Uh[u�|���;+�x�>�H�H�dL^s�.�ӧ�e���Q%��{��+w����D�re6:��s$�{�Wh9t��{��
�"�(��xeN3����{J/j��ۋ�/ fw��ff�L�4�mff;�\4�w�TrӺ�������X�zՃdہq����WP���@�̖���~��Mq� K��
�_��g�����l��yk�gλ����hL"x���i�SJ �o��e�W�Y�k�)A�u\�4����
������`>@�����Q�r5�s�*S�R~}��f����Ul۽a�Yq=>��LV�4� �QPP:1�Cc����!��=��5ce'�Q]-C����9��FRP�i���N�ns��V�6;L�u�F|vEB���[���0�S4�=��^2M*��6��U�OV���ºϸ{�O7��c6cc�oi��n�x�����G�ӥxi���+���:$G��ZI�[��(��<�N;�i��*7��iÔ�ύN�$�_]`O�I��T��8��mfvm7r�|.�X���ka+Ä�ۡfU�fH˼�'��ǖ8a��������4�P�BѦѧ�3����ݿCǃ���h+�P��Z%�+&>	U�h��>ҍz�-�OLV�EC��ܐ���{��^��ɵKv�;9�3V�����k 5+����X��]zub�إ��+gf��v�}N���^�����;(���������	T;-%�*�3z�e=�Q��<��r,6�����,|�J�6�w着���r�5��`��j�\�����E_���sȄ8m��U������ɮu���N^�0�p;v;�:�9���궥���G�x���Z2}I��n�s��18X�V.�8T���������^@�Z d6��]&"�<��2�׸�ҏ�uٮ���C�qu���$�蓱��}n�[����O:�;=��	����e��O6t��]������5���9r�x{����|���ϸ���|#���x	^��a�=w� ���X*��ե�-}�Z��]��<pH���מ)���pu	[|�lB������ʽ�����[f��E=����n_^�C��致�`�G�ߪ'g�֓�Q}��;�Ş=c��xH&FG�z�7�*KQ:�a1W��mܑ��kv$S)��v���4����}���Ԇ2J�Jh���j�۱�䐓�0'Z�5[6�z���x�$��z�� ^�b��&��W�wؖ���vg�Ç-OU8U�MK�ī��i����u��\ky���\�|jɛ�[�����<�-��#i�I��'i:q�l�IT���Y�;��<{�h��/7��N�Eud.��,��Օ���m;M��Q�=r�#q�����]��Vs���^��	ἶ��d�D�/)�"�Ű.<��:|o�X�-Ч�o�v�@o��>��B�|��{�o5M*ר�6T�z"�o͓>���k��vԳ\�<�S�r���?��L�т*����Ud"B�GNL;���<���.%�
/%�[��m*I��g�
��Μ0�9��V
��ж9�\1�Nx�u��}��'~�˸=X��%Z��鮔��L��h�s���n�W5Y����ѩ�F�R��}�CH&d˶��<p�
S�0�}O�h�F���Y!y�wwk��z����*���J�����X]�mR���5!���'�ajT�a��K �{*�Q�������5hg�u�L���K0{����6��.�u�-�?x�do<�>�^ɗ�E�0X�V�A��_��LJF]���{A����*AS�q<1f��v�'xۍ���=]�k��`�Sb��]��v�p���^3� +�%���f(4y��m�휭��'0�Ϝ��s7L����\S�\d�V�"'0͕L��sg���{r �s�K�N��3!�wI�_vY��m�=�I�2��������+��z��k�*���MT���~u�&�S�"�9m4̣����*�A��,�㷙�]}�.�6�ӎ�(��Ƭ���b43y���Gi�Jr�X$&7ol�(�Y�tMh�֝d�`�jU�3�����kq]`��$tN����+r�h�s�������{�6�Ӵ�g]�ňZ
D�/xS.�7�����y|cx)��$8@l%Gu],�z�:�ۻf���t���A�����a�=���VEH��>��/m�$��ʐp�/�X��q�{������#�vnAz͇��=w-y�5��B�uH;*�r��Ge`#�o`����L�n$hm�O������ĸk�������,�0��hY�2�TWCa�`h��+#�]bJQ"��i�PC�c+�n��b�o �����S�:�[�ԍZD��&n-�F�!ʝ��i��ɻ�=�(f%�M,�M��"&�����[u"T�o�]M����_^�\��}ڸof��桷yXGb��jF��VP)�f�u��d�i*iX���в6<�9�	���ł���Rh���II��o}ݘVж�w��V9��1���6�$z�g̜5k�r
���ё�j�e�,{:�5|EB}��S�ν�)��rø��ת�@��#ʲf_�s�bC!�.9Ϥ*��&^3�Ƀ����KX`��6)�e'Z�s+��w
H���[7�U6�6����`#q�<czh�"�!sB���s+w���/�0��b�e����*feZ#���(;�n�6:�W7uz/�6�\��+@�`U�&����|j�5��2ƴ�! �<mH��<��̌ ,c�̈J��b��h=�r�N�W����[b���v�|a�������9&kej�b�6�2TҤ��,X�w�ؾm�ɹ��U��xU�MLq�A��Q\�J���kp�!�K*]��F�XH\m�����i\��;�����7b��A�?wu�ӭ�U��b��u���7�d=Yڸ���}s;�4�,}+bY��P�&�����;�a���ު��<��ȝ^���Q�D�:_:��e�jm6�*s;���|1͠��,��A1m�GS������ ���"��\�S�}�w�"6p���ZBTtbn�L��]���Wn�iz=�zJ�q��U��
m�����z��/�'5�]H�r̻ �7��-GX��"�{�ڃ
�ޘ}T��1��T�I��i.�C�4���3쒮��ü��غ曎{�)�=�}���ĭ5�^���2�����b��y�tN[7��J'�S��� )\]��E��V���W(�vR�x%�7�������A�rY�ɤ�²�w͎�>��yV�m�ޚ�CtYj�j�r��<��&��u����tw��0���%� 1a;7M�]˸�݃�M�"�ɗ�I~&�@�	��h��9sY��Sͪ"�b剶�EMjܮf�6M5Mrq:+E%$E��[��k��'0j�����79�M%X�NN����q�%[�j�DG6J&���U4E\٦gF���9�0T55G#3Ujg�ˑ����.U��i�mO3�kF(��b�4kQEEI8�lΦ���h���G��m�*�b*
������F$���(��Z�cMEs9
�v�h1�9�����q4ۛ�\�E	TkA�#DAM71����MSlh���AI[�uF��V�kA�LI�i(h��
�9�4[���1����h���֪*�A��b��&��ѹ��EA�ڞcS6�F�14UEۆ�ȝ`���V�m�N��h��5؇@$@�|*��
��k��=��ޠ5h��:s֢�����- �	�y�p��F�}	�o�	���Z�H%何�,��ylbӖ��~�����5�ʔ���;$�q��$Sl�6�l���4�w�
 v�5�����~T��p�����-�b�uj�W�p�SE��EA}�S���TC�S��!�U��C~A��굅��v-�P8�����!֏ϼ|���Զ�}��������./����qש���b��������=�4�>h���f}9�]`�-��m�a:y3YZ��NL;i YL�ʼ�D
�g#��_9�<�y>u_��
���L�yuѤ;��c����a��
��3��(䔥�f��.��^pw��v	��cNϽ��n�ù����KN���vU���D��	�[%d�SyY����֩�y�,`���q�W:�qUX&	�k��|�V]c��gxmA�/7t�C���7�������?����Y�s�n��;=+j�pn��F9`����*�
��?{~�y;��Xɪf����2�A��;oZ��V5\�	�y�T�w���צҺ�:WtΪ=����U3�(W�Sl��hi4�'h�$�@�:�|w-hV�� Zİ�5����N���H��u��(�e�a���s�]�7�n�����[���"7�+���3ދ����3�Gx�QCv$�{�i'�TG�̹�����E�#.�hwS�k�i\����00�<�g5-�9��U����n�f�f���vw���V���v�e39����P���JX¶w�t4槍�,S���?EW���q���(��|�U.V1w����]0z�e�����0�$�2�ؽ�d,<x�Ԩ[��O�.ڢ����]Y����;p;�o�Q�Pp��͓����EiWY��)ڿ�~���V =�@�s.�cQ�^�[�8����;)�/T�����{�)�j�XY�;�<�0��(&r"��J �Նf���j�e���k"�,�d����1I<��0{|Û!�8%��㋴�%��i�`W�'U����Vq��n���-WH��z��~�%p���n�PZi�L�lJ䢎BW�Y���*�[T�i�#g�Z[�H��h�j��hb��BjI	/���+ nJ;�Z��9����5��[��)ԗ,o"�A-;���w�뗦�i�Nݫ��$P��u��E˧0�҉� u]������CN�2L03OR�n�NK�ͧ��C���{.��Q�I��_f�1�~�J+���}bF���-��ﭥ��+�BmD;0
C'c��:6�uY��x�e���H�O�LmN�{��3z�8�.��9��y�N�')]�ǲ�)�l12�?�R�^[�� ��>ڜ�囪)�q�oY&���Na�V�M�U�%RbX�Pn�Us˜'���;=#�����W�M���U�9�XJ�B�s~Ye\�6k����8l�6��IjO+��{j��ר8��m�3��ժ�ʦuZ�|޼^�Ƃ^,�}�zNt�b_og�l����yi��΋y'��ʓGB��/���-%13Zl��4��1�S13l�Z�b������[E.>a��{6H��vw{�+��D�b�X�%���S,F"�z��l�g���_��N/���K�,�%�N���.-+���t��Yb��z"���k�qD;��y]����'�eC�^ܵV*����r�+bcSVm�^Hmw�Y��>S���ў��&��m<B`�ܰ���E��-e�Kak��-:�����UO�^�<h�zX��]������e��օ���^.o�����V��+)��e�L^\;�ےǕ�G�J���!�g���JW�;V��6nY�7q��XGv�Fr[�;.ɥn')�Q��]^�oy��o%,*��:�� ��M���{,�;U]�/.�͏-��u�_\	]þ�uy�2�5���OM���[�J���+���ό�6��DzwVƈ~���N�d��N\}^}��iK$ۢ�n�h2�(�M�ш�5?i��\u왛���G�1\}��ߘ��s�[�*�jf�[[S�&�ήs�WC��-�J$���k�ҷ��#�SXe��8�2�u)c>�&�\�)��Z���ຳ� �zj��z{܏˦C_��ԺmW,*z�d�[������Bk5�#v��FS��fvó�V��ڿk����4?)�7�1�?����i�z�ǳ=t ��A��v�s��q]9۶(�0sI]�M�P{؊4��52�"h۪.Qc�UD�4(s�L�Jq.�7+Z�^�b',��V1{x��AH)�[*��Y^1M��[C���r�>��;ݙ�u�b��8���y�>�Ƒ�ɍ!����{�F�6�q�:v9]X���#R8�H[�P]wE��8P�����Z5�އ�9uiԛg��k+"�=;s��ԝuzl���_�2�1�6i�&)]w�l�&�V�{"fD�5��/4W�7i�S�Ly������n[;���g�pE�Q-��d��&i"��QBX��@��共f��=�h�x��^�dCY��T{v�ט�,�Xd����ګ�xMMD���jH;��L~|7Õσ����o˿X�����t��7��b�x��Խ;���Ww���6��\Z>}�V-]K����12u��n[So�N���W�8������U�V���.��+�S���ח��g����q{�WOSm[R�x�gyt���������PF��t�|�z<��y�������ڧ�l)]2·.Vd�6r��`ݦ9K�,�u�1`Ɇ���^{�ڠ~�R���}9Aj��[WXP[�Y�A��\o���smz.P���Y7����r�o�q���ϝ�.�ߛ1jV��v�W�\�&�}3���*��-�s	���
rZ|�}�U��_����`�1�C�S���*�("�T޷�[5��8��7�V�)�h*g'v���MEc�o��m�L���/���B�GA�x��<���ʻR�7�h홏9$�y�W(�Q���4�0�2��� ���}��E�T��La�7y�����	[:RVl��6]��ђ��}��ܙ}cr�6jڧ:��e�g"AQ��E��R���,��W�V=g�I�����������<�2�K��2.n��}<;�pj�na��U���*�ϕ؏I�|�#8��������̞���X���5s��5�����%��6ϊ��l�˦~v1��PW�*~do-����lBͬ�sP۲�BR,�Z����˙x�ynt�yNT�A���d�[����[�K���3���|�����(�e��S���徝7Y&��5�I���ꅸ��=Wfj�b���V)a%�H�w�m�h�Yi���PZ׼*�O�X�fZ�ϩ�����*/��2	ޙ'��a�M�T�秩P��x��,�����p]@�CJhgm����Re����ԙ��;2�e�bj����k!,���Ѵ����3���ʱ�u1+{5���"M����y�Y��+D�1���V�
נߦI��$"�X��,F���Cw���d롣�e��z�2U����@ҥ�v�gk;I	���j�#�5�r�7�+0΀���� �W�)��]w��6�ԁ
���C{z`���E&���/w���9|qq���-�[vV�O5�]x�:%��`B�L2�AS݆nw�'#}�]��4>��ڡfh-4�`ϰ%{Z��6�m%gvj��g�_?Uy�v��{���C����#��`��i�9���kw��5�̈�MF��{�(oZ��x{e��n:��J��M:]j�~~�����<�c�lϴ�,�ս*R���=�)�+"ʈ���4i��:��X���f��,
ݭI�����Tʓ�,[=D6�{NJ|�)����	��"Wzs�J�V>��Iz�����*$�Ӂ�R!�dq��k�8���n��թ�B��Y�N�$,d�i!6ʙ��tC��a&擆��U�9��tҪ�hC��Nl�M{���+"Y$)�U(צ�[��&�̳R�����0��RP-Ri�Ml]��J)�ǛF�x;�n����z�R�0[���lo�ν#�V��uF��m�u�[	�hrU��t�n�"�Շ���w��5�5j��ˑ������(Y��k�����Ũ^w�����2�����F�r;n�^!�%��Qz�'st�m�	��>�v*/_�7sؽ�.z�=���*��*;4�f��*-�]�r5���ӓ�OT��o'��~<�JĻ�<,jR��S��{�[`z�p�-;�#��g�o�����׷A��b�^ڧԲ������w*�����Z�w��=�r��{,�~�8qv��K�v�ǖ*6�+�x���c�^s�=�UG�������.NJ��	�<a��������u���|PS7�!�S� ���z��~��Xۚ)�e�4c�TS+��0.�N}[�Z�c:ř�t�3��խ[�)d��f)����U�ð=�{ᣪ.s���Ն�.�ޞ�K:k��C�W��(���y����w��F��ZvUl�ϯ�Y��0'^Y��t�v<��N�wU?T|;w����4����g,�F7'�u�w��t���q�_�,G�(����:�6��q�'�w��V⭍
��ekX(���u���v�S��Uy* ��D�d쫚[��o_P�%b+�gu>���4;Gi[NS-��u�"�ñ9۾8���w��U}U�w�W&�)�/}*J�6`�3ۓ>v�r�c�z}<J�ϑc���g\�/r��Sg��)��u��������X�eT���2�,r���"�0�~�t-�s�|9gP[*�V��Lw��43A����P�Y[��̻R|L����=6tY3Ԏ�S�Cn���3��-��|�X�(ǿB�eu�;��mH��ܦ'��=��?{�*i6!�ډ�݀o�P�d�- J�"��5�sѡ��}J>����ΐ����_\�ٚ�#�m�7�ʜڣM���V������S�h��ܬ�L����Z7^Q�(gd�������[}�)dNT���A++n��^��jT)c����������'��i�#t.����j�[�.�t��j>ϗy@i�9��	%C�q�8�ys���X���{�Ӭ�7I��Dש�C�d[�-��+��9M�o�D�߱�@�Ĝ�vi�б�{}V��o��	��������3���Y��2�Y�@l:&��Yu�
�j�E�R�+��rg��/S���K�1D��^ok�ғԳq�wә�˫q+F��`�jԬ�(���Ϟ���zI溧��a}�K)�6�W-V�3����瑱q�f	��m�4��=�7���sW�+�mZ�y��崧�N���=sk,aK��{˝^1��^�a8T�3Aj�0e�WLQ[��)e`c1q �K[F��KaZs7�god�g��X���?,�m>}��Esoӯ���z��'�Ν:�t����6�[��J�t�q�{��;Z�^K�y����WF���+�wN&۽X�T�L�~]>;���t����`������d�� U�]a"h��f��`�R:�ǸeRb|Tʓl쏴�U���O�2�j�Yp����h��CN���Q����.�h�c*�CI��ve6׊z����o��+�
�6X��5}䫵|燷���|�P�1����Q�DE�����9��^5n��fn}I�4툳k)��۲�Bvʱ��8�@��k�D�i�b�%
h��Q�M0�)�I�j�4�Q�e&�|����ն%c��[:�f��D�F/�ͱ���x^��t�hf��HE�6�d����^_`�+/�'�7M`,ҫ��Dbw�$�OG@nKY9�F�����u)t��"�1�W�ms�w�^{}lu�V�f��Hb��pm�x���Q�ؒt��}���5V����٧r��]�N��Z����>V��������A�@�й�`V-�1������������u�X@�Α�'����LҘ���-�)p��ᗢ�H���<e�Ϯ�e�r�[ܓ;)��y�ܪ��Yb�r���{��N�
\�=��WO��b�Q�`��N��:�8H���1E��p�=��nuCSGWR8�U�,��wk빱�ۚ��sYZ��CP��]���Y�t�������/+c��Op�j:!�7{�Tg�v����]Ϧ*3�����2�,��.�����FH���+'�r��[i��J�J�r�N��8��i�|Ju�[����Jm;�#a�y�#\b��N���K�7[�3mV��͠~aT�ޱ]F�◦��wr�$�c�@��j;$Ճ)(���f�V
���
�cx�u�&�<i�#������73�(���q�(��
�e�N��˫�Z�oP]*4����b��82�n3f�\� ��|喛�컥CF_s��s_�O:
|�l�4�`N�㹠p�t�p[@�-�b&��}1����e���چ@o��|�bࡨq��E1�"՞�F�/
V�]h
z����!�u�C����3),Vy&�ʼ�9���ċ�2���73P�j�I�R���9�����V�s/�;q���X���㘕^���M��
��/:oft�K�]�
"XDf�P�hN�@��@�j�f[��}Ȃ��۬�	�]Y�0��{�S��v�q̮�M`�E`�J`�j�_�E�`N�<P�B�ⅷ��k竻���T�)ݎ7���Y'yAكj=�n[lՋi+���򧷏�z�	y����H5��Ȭ�\��oX=�
�@5�و�<jK5��Ӽ�r�
h�ZF��J}V��Zk����S7qI�
v滹S�]��0V�d��-O�E�v4������JU;��ݜ��O���dԣ���+X�
�gV3�r��w�.v����p\�j�Ů!�u���t�u��j�5������v��g,HJj�r�N�t˦��
�W%�	{ڎL�� hN][���o���vKԱ�o�-]օ��}�=z;k�ĩN����-ey�/�U�9�{&�_��\�fEt)��5��5|@®A��qE�*�����̎l^ز[�Y�>����䌬ĲoiLݳਚ�!��D���q��9w���bw+��p��l�J>z���Z�!�0-��v�9\��{ٛ�gk��}���N���=F�}����X��������M��wN䬐�g�a����b�;�kzB"�뻵䀘���5KC^��/&�*��c,��*vY�A:�iӏk4��oo:�_T�x)�	�>�ULDEld�"��50QZs͢*���m���6
������*��DDRr�PM$lj9h�l0E�r�s'#Eh��UTT�-��"5�hkmT��r�\���+��.l<�4I;��&� �3�4�TA\�s���,Ub�X�i�rq76��v�.ULTD�hܵTUED�m���P�lf���6�ي嚢(�0UEU5�ᢊ�Ͷ���Ƶ�8rq1�Y��F#X9<ی\�3�TQ��W,0�lfHbi�r.&�8�i�b9�I�DS\�1ET4S͊.l�TEZ�TG,D��nLF��*��$�MQN�m�5��sj�n�vQTM�G-W-%5\�s	���� &�b��`֊��H*��T(P *·m���K��B����:Н�܇��/���ܰ��^Ȍ��WU�7�C��{[Y�wk-�꼨�'e�E��Ҝ��U��WҒ�{{�J̉��O�Ia��)���J��L���h�9��R��ߍB��>(I<c�ꒅ/l�@=S��o�p*���]��p������fZ��i���z�R��P>R1��!ާ<�S�NT�`גS�5�R���o�7���ڞ���Sh����Z��My��M-�d��j�B���G���7i^ҲE/,�9J.�B���>�j}e�㪶�2���i�f���д��y�r�z�˙��O#}һ}��`ӈ�ٗXN/Ic��͢�P;� ��Pݫ�J[�V�����X�V0;�w�Y�����߂A��l�v�i���3rJ���2̢�9�3���&��<��v�'�U�޺
q����ة�̄�geY}0�e�^kY��`���ri�o9�Uvq��5�+.��w�ʻ=H�x^'�Q�vv.�nגm�L��T}8/SȗK��j��S���|B*Qp��':^���Ms:��r+[��>�'�k�������ݞ����F�J>T.dў����+jl��҇kGi�ՉZդ�2��)+7-,7����=�S���V��@�	�s����g%��
1��DGy���ai5��2��x��wﮧ-�əWބ��D�����fX�R�U����
{b�b�.ZLH�I^<�lJl1L�؛��q]3���9��Z�<�1��)Tq#�&�3�a�)�|U�!��;�$�'�h;qe]ò�3u� ۶�x	[�g���M�LJ�^}�t_���������*��K�� �	�h��Wp���&��lWݐe��IY�"�a�}�eq��C[�d^���%�}����P�N���]�O������T�����ӆH�E���It���x_P\O:+��0��C)W��&��e�'"�k�Q-4%^��y��Oq+���Ao�V���~��SO�o˩{i�,�:�_��75׵ۦw��3ݜ����{ǆҖ��z�U@�q�8���]K���M��.[�֚AOn/!�bw���mo���ף����bCO������$��W[�BӄK�߃�u~-�?Y��|���(��D����y�|7�eۢn(;���q�sk�ՈLӡ���w�O���g\k-�'_*�C���d�������������z8�C�!nq���MvJ��<ڼYT����qu�.��-��QGk���[��������v�}��8�^�f��Ju����,�a��j�;�G�r��!��{t`��l����b��n�(�4����F[WV�n�JY,i?@����=����G��?{7^�h���ZM\�ņw`�y�2�"!���J�0�C�L*E�,�2�'͒1Ҧg�7-!�:��(�Y؜�-�1��v��ި�ʱ5[�J<}\�eW����q���m�嵂\��}<M/A���g�(���3x�'5l�L�Ұ��fY��"8����wӊ��+9�,"ڧ~��Nf֝b��iɂ�U���k�y��v�!�{)L���+�;���WFI�Ur���/L&��)�Cn���[�E�S6ƙ[8�^tHؽ��(���FL'.��*�B�a��s���)�ш�R.bI/	5�] ��U�4�����nz27ȣΊ�\�%�ʐ�=0z�?{Z��@%)��le�8�� /�cr�,x@zX����TmTɫ�U���o*,Ɉ[���)]��wx��������J���48[rM�&���n�T�Q==���6�緌Q��|r+Qr�6�:���|��|��D7|"�D�d�������R��j�L#����B���ɺ�G,�욻SW>��"ϊH�����1a�*!lfW>+�ϳ=��S�җ����k���\Z>}�V)u�j�T}����u^�@�N�O���vV���~�׵���Zگr��U{,�s�4;D{���w0'�M�R�o�yjo�~3��*���~�����䯚�-�ÀwOlP�e�M����3z	��o��2ԛL���,+r�f#F��N4�M����3�t�%h�QE�KSN#O�=Aj�a�-��8�ݤ ��׸xJ��xjE7<z��.t�r��$\�Ӭr��Ӹ����}Zkh�kE��8�ɱ��ݵ���i�%�e-zsd㙔��P�����b�lkb��B��XswW��e�M�啡�������Kc�����3ʰP�]���ͫ�߯�����'ֶ'0�+v���s^X�U&%��Pi�7�}E���Z����ُ���x����kӛ+ �W�࣋�G�ŖD�%S��:��kPh�mp��""�b���7���d��]Můz���w��\�m��i\*��rq[D���vu���n�H%l��Ok;C�U�˧*�i�h������}_}؈�'`���b�:�T�n�ʆ��-�u+��4��0�=Y`�Y��o�nښ������u��b���G�PEl-gTP�-m;&�&2*aZݕ�q�V�'�ƙ���O�?=�:z�t[���:OT�	�e9j�;�1ìM�*g�:�}�y0�G�7��R�>ar�>�3J�Vh෩o�N)�l�sD��3�PO������e�|���p���e�T5ػ�V��닽d�	K��m'�c�(QM��V��츦9�Ǽ���9������u)�uK5\\���}��mIi�j���H��y!�w�J��ir�A鹧/����q��7|=EhL�����]K��I��_N�q^K�ǼX���0��_	�� �.C����ET���.߈^�]S���);i�N�q;�a��MĒI3V�b{����	+���ؕ��u����Dzu�Kk����n�����+J��͡N���e��9y�mM�j9"Z �����mퟺ�e�J�s.<S`̊���ݧ��w�q74�����y�mv��b1�t���w���`u��"_j6r����w-J;�4�wW~�8A�%���o{ޖ�±��b3���6ir��C�t�KmycA��=��X��Q3�q)����1��t��{r��+��H5��[��<�uu�x�v�j��pj��Y7�/n��M$��vU��wj�,�tZ�ѮM�}���&���ܔ�5��2��A-yj:��ga���u�l�L����Z�r�CC*��J��F5$�de�����9[Lv��-9�AĴ�5���0���I�����{=r,�iE��m7-����$o���u���n����y��&�ى��BTSiT.L ����rԜAۂ�fе���3B��uD��|�� Ε*�Y^1L�����J5�[o�N9~~��aə����%0x�y�eR���o�����������dd�7�e0;��K7�j8���s{�6-){J篝�EF��^c�O�f��*-4�ë��	��l�a+��)l�����-+}̥���k�f��g-SZN�͠���b�c��*�p�'�]'9�
�-�m=�񰬋��NZj`����u�V�c^)���)�;3��t��L8D�]-�����]�&����:޻���7��9l'l��$O5۾T�}�j����+�`�R�i3��N�)�Uk��*q,XW��ɱ���:�T=\���ql��E͖�-�-b�b��O���YY����z{��/R�Nq�`>!Or��/LuY�.���^�>�آӪG���t��)]x�[J+n�fm]92���4+8�Ƙ��0���Ƭ��Ʀk�Ϋse��t�
܄�A��b�n�h-1V�$�Z����|�D�Q
)�	���Z��Xh�l�ĴW�I�ٖW�e��P�?[��>�,�R��z�n:�YZ��w��q���2�4���r���:mxm�A�ے���h��g��.��k]���s;"w�j�O$�ٹ^D��~���9�QJM��L;i l���(v�h�[R�= 0�����8UV���i��sK̲�h�N�K;aB\�\�D���l�6t�&c��5�u��/m)T��>�W.3�RW�ǲ��.B�ʺְ��!ĥ���rT܆�vG;�m�'h��S8�Hf�k\��3�o�`X둊��k؛[]˒-m.=BWR����	���էj.�M��U_Sj��#۝�Q����ןV�,`rM3�O�Ĭd�T]�l�����h�1m[�ݴԃ�޸�^��g5��+ak��)�SiT�f�sy�}������)����8���!���5m;��	k%襣�^���a�El��i�[BJ���%�J�j�2�~*���n��z�u�!־�М`���G7`J��$Ţ�!|�h�r�f�WK(�Z�������oV/8⥞0q�w*..�l��Ƚo�l�*��-w˖P�r,����Ln�TSD����H��ͅ�g�M>�X����Z%�[�4�y�JP��,i��Fܞv��'����sZ���[,�6ѵ�rVꍬ��Bg��=�\~�����\9|f�����;i��l)Z²̬�4�fc��DT$�(ӕ���+���X�k�4SN#/�]bM�����{�f�n�h������3�l*+{w�(6`5�;Su)hZ�V]}j�.��rP�ܩ���*`�+U׍�h�4ʝ;r��BhT��u�'J�y˦�؈����&��pb�v���>=��Yٕ�p���W!�rL��,�[x��e�}_U,�­�$��̘&��͜��;K�,p:9����*�y��-c\��E�/�����M�yt��nX���Uh�8q�k!����uG�6��׶��]K���2�,�6�R&�6�RǸ*R��Pi�ܖ�4b7�w:w^2{Zt���lFv��`8��d+�8�dĕC��gX%�Q��Qz�Q�g7V�*��)�q�5}5}���~��wyW=.���ח8�o^�oTi!�*NȲ6�Y�\4��9Wt��PY�(ԧ�V��SK�"l/\Si�
kvȓrԝD�6����{ʖ��Y�t�2!5�	�Yf��R�SG�R��oI��8�K��SR�h�on��\�F�\/#g6ch����b�!v�.f�Bܡ� �P�<�A�DY�{��>�}�~z��ƴ��e*f;4�־P/ͪ��-wʈ�^�mO#�a��~ʝ���ŝ��&�XL�r�K�\�5,�p��隬�'��+�e��G�M��y��<"2^ꝯCuzT�j,��NÙ:c�i=����A��c�����:(I���*���^}ל��QWZ��R�U�i����X&�b���A�����Ë�/g�����h��j�1�>�=F���8zW˼د �1NPaW&��5��{y�p�IPvمUυ����[�-jq5�Yh���{��=ds�)غ�pf`�Ҿ�Hϻō�{��[g�bWg,8�H^�]S��,�;У������{��N������O��崧�CH�w7�k_��ٞ��n���M�0�o�C��C��>��[�)c�ڛd�l�h2�+H՚�S�V�䬲�{&W�.߈�Ɵ�c����I��*���1��{N��Ά6��'�4�	���D�F*��J��wu��̦X�T%H�[Rn^�)]ʤ�壷���}�+�����O�f�8����M�Ш��)�e�g��Ѵ���1���2m���v�F�r����Օ��aE�8ki���Dbk[��N&|�t���t!�A�E��v�c^��ڥ�9X-��7X�^e
�3�d�����\��*��ٱ��%���2
���J��UVfĦ��A5�D5+��n��|8��T��Y�Q�/z��']���U������Ak���˭�~�e�˾�j���> m}N���W�v�*��B�����)m%�����;k�G��x��=WMtW��E=%˃��"NY�5Qu)�[�.�V��ڼ�lG���_��Y�V�g�7B����X�j��u�J֞�t����"�0�C!��tCT[WN����/�1Yv.�3�U�΋4�:K���2k_)N�ݕ��-��0�G�+c�9�ݽ��KV( �`ӌ�/��o�=����v�o�>a�o��Z�4k<�J�#���6�^΢η�9��ml��P�Oz�0^sr��H.ͫ^�8D�Z�7H��]8r��ҭ�3e.5�a�Ƨ(���A�(n��8 �-�/�m��(<|z��wY�\�5Ҭ��V�M�3�Al�;��EO7�LgdL�h[����3�y���]"0n�ȭ�6:�srC�^0{�<�Ԉ!k��'R�-d�7Ԙ�얛)[Zj·�b��x��K6ܫ�b"G����w^���U����FN�C���d��B��h�J�X�l��54ǷQ^*©f��!yگ��n��+�����Lg-IA�ȱ����FG�Ѩ�À�]�O_r'RT+ t���/\��+(flG�.0�b]�m,"�|f���V����Ύ�9�[��l^�g��t�j�EiB����z��xл���/���,��}c�K44�Ef]� ��Ff����E��%
���˹��K�F�__3-a�����Z9t�ȅ`�Q!���N��ٔF�3�Zy\POo��EC%r{Fn �]��'�t��a��Ѵ���Y���*�����t�9r�π�����U��ߺO;6\^غ��V [f���T�n�˧WK)W���7�6��N��y(S�oZ�o���dʻzEсzn���)��ed���U!]V����uɈ:�����Nm9TΓ^�@Y����_lT�;eA�]�g�wJ��y�{������z���/I�(P�+s�U��+/EB+bn�s���+�'K��9���U���fn��%�m��,c5�@������U�R�q�l�
��;����'a����͚,LDO���6��ו­���yr�ߔLv�7��In��Ed��y��*V�����/�Ρ��8c����s)E\��Ճs���O5�+DP*�f�]%���\͎�P꡸�p=�Q_�7)ش�`�)r\�V�C�:�ݾ+)eaGne?���vBu�ַU�]�R{�Vֈ�MȮ�mwK��<Yx�A8���&��pk̙��v�:!�)��Cn�>��]����\˵��l�v�X�����y��a�WD���sP�\� �YK#�PM ��n�^]�{Kn�z��|�8Fu`=/6�nf�ȣ����`nl��%�D�H��779������U$SMEET1s��NG&� ���H�����L�la��������5���N��F�*$�6yb�Qh5��U5L�576��nlp����T�U�TG6��3QE1LEEE6�+Nym\�E�p�L\ےi���1���f
��lj("����*��II��u��m�UE5MPV�b����(��ks���)��*fj**�lŬE5UZ515A$�D5QVآ����������AUTU�\�tDM1�V�(�������"��ֈ&(���Uɣr�Pr�'Q$IE%Er1H��Z1�lj*�*֢�c��������$EDT���X(�AQ$�ƵQLsNFH()�#���cKAT�DUEUETA?A 9Mc}!��ѣv]Z�*-56��%������iK�]>�Zy�t�5�6�U��C���I棝�pMF�2q��w����f�g�Gv
����U�T�Q�~y�%�kiT�h�s�^n}^����9l�z�x��K�Vviz�Q�!iP�΋,��Y
h�J5�哮'���?Znp��9Q��z('���Rt�V*8#�f�b�����"�]�"4;eO�a|��#bT���w2�%�$ܳ�J��|�e.�N'� �O��bE3{׽�Z����_sS��dg���p�{.+]�����y���>�}�-_�,�؃/�Ft�S�J�ԧ����^Il�[[C��\t�����ћ^t3��l���`�\e�L�u�M"��H����9�/+�Kغ*��%h���k�%��������jE�'ܳe��l�˕���Q��ͮJ��{��ßv�m�ٙk,��v��������l+ZS^���v�{�I�n��8��j�/�6"W6��1�0NXQMU��,��2u�����c���y<����s3,}|��N��G����\�3�c�yi�8]���@jn��K�y���7~��_rƅ��-P�ˈaS�GNb���7���uxG-�6`�8���t��C�L�O6�*�|�)�X4�v��V�L����i����U��e��w����9L�:Vm��3<�K"�dƱ�h��YU����7����IMi��rBr���E%�J����� X�4
���n��&���og#v�[U��M�V=b�&�Z�L�nL�i�h��ٖ��OZR������<5q��ˬ��A^9��ԽMK1�[�h<^�cIb��$���~���T�.�ۘ���sI��U��v �(h�m�nB���{���5G�.u�X��.�X�sT*(�-d��M���,�Ʀ3Uk`�����ϥ_�{��+�h����6�Y��n�2u	m�av{Z�7	m��L�J񈭤-��@�zanW���j�5~r��.���qMN��.��3'.7W���}�@��D����FvM]���Y�~gGȻ�]�=ӏ;���yWL~����/-]��]��{.-�����b���)��<c}�~�-��w���K�S;-*R�%;�K� ��\�:���A�YW��k��أ��2�iz2����fQ:P>|9��Cہy20�wU�����_N5��O)i48N����Y--�<:�7��<�J�+��ew9��opY�Ҭ� ]���H��𖻧򾪨�Go\�>�&~�b�W�{��jKO�V-p�f�DO�^��Dn�X��v<�t���P��7Ո���x�z�kZ�VT<��w��ػ�k��}K��{4V+�4H���)�]�ס\z�M=�}O�w��;^]�>�7�7��.T�^�7�i�Vr��&� �܊a8�>���W��*�٦ݣma���κ0I٭LJ[��K%�V�1�i�4Ɗ`��g����d��]�W�]Jy�������9m��(��e)��c�V�U��+p<f�Iڮ�3��ָ-��{NW�-ئk[�ju"i�ne,{��*��@б����\o%�ד�9���:kg���O����it�o�w�5=���������N�Y�6��a�Nի�*{��}�2���葾�F�G?xߋ�1Q��-�[�^�D�Y�$�Ƶ[bH!�e�|\N�K��P�]ϨtU����k^����2*=u�����)%��mefG�;~�'m`#�5����>kg}.\ޫ�֮e�bn�r#<*�nW�8g���`S`�v��:*b��/Bms��#kM,��s��gY���W��i�v�7�ިm�3$�wf��+��YSA�[a��	7,ԝCN؆�k��-�4�'��S��m�cX��ԥr��9�k�\�{�����Ef�f8��&��j�y����a�CY1��|v�H�����Xu��6�n>!�؂�o�ҵ�^^MY�fŎ,�d�%d�M,ח��UȝV/�8��N�5��N2l���pWx}^��q�<��V-]�0����X�������2v�b"�	Vn
8O�ڷ5e��C/sU���������R���K)���by�st�9"����E;�"q>��ѯ����Į�r�=�k-�G�����gU�jk9�D�����b��6,&��"��"�4�1�
�M9j����n�͝NMB��3�	]1ZQ�/z�UiZ�5[F�A�%�t�	����?zECdO��Ϸ��~^�7��3�����^6{q]�ӮJ8� �.��ǭs8��P������c)�a ��W�O���� hb��j!�>�v�ܪx+)h�Npچ�0��������Fwwxoe��f1�j�r�g��͚ŋ��빫�m��Z��X���OZ��ܛ/x�|j=�8�sjvILt������Uf΃[����c���Ն�d�͓݆�L�g���5�趕�����f�ï2^�F,�0�FD#2ו�v*dk�*�4u]5��Na�V��+ٷ)�k#�!m��,sY,%�i6���>���Uf��·��Ԩw�A�rU�%�ef֝%U��ܳ9�fJ�I�3��4�B�%��Г-�bnZ5�W�5b�9Q����Ot��'���W�*{�:�L�^QM�U�!��;�$ނƠ4�NA`�Sgp�u9�'֖c݀K6�*��,��Se�4��Sm:��p���G"��O~����K�ٴ���M|v�$Ym�S-u0g^��!77y+`��)�YoJ��9굒͇fbf;5��3m�4Y��4�����C'v'��ن��[2��|{H.�w��Ԥ���үl�Ms:w4�N�]8=�y"��m�e��n��q^���g����Գ|�^�)i���ؒp5K���U��w�y�U�}����7fgD���2\�\^%"�n�Y���7G3��9��'5�ޘ��xn�C�l���Ur��7]�w�%�S�&����#Kȇ1�kF#2bKQR+a�SkH�����"Tmdԥ��n��Z����J��d��b0/�{�w"�J����賱�\�nMvG��m��R�o�yk]YP�/*����3������o�ݷ��O"b��ռ֥-2Ic�O*6�M=����mOA������#MA�׾|�>�ؒh��$	j�b2�CL���Xh�`*�֭׫�$��M��/E�FU�$��5�����b�	��SA-I-pv}���ks�7�4ooN��e[BCj�WJ�^h���t� �}��7�ِ#�zg�t���]��^���k�8ˤ4��>�Wa9M�*U-���37��b�3�j��Na�x[L��fX�UȳPcS�:��-�u�xD�Jְ�Qn!t�n����Z�6bN'��V�U��s~�؇�g�d��N���\Q��z��e0cq�N ���Y��j7PRVʦu��]+vA��P�Sy��M�ʷB*>#d�t>�s��
��hP�"W+�3.K���]*y�I��WfS�݂����h�۴�QTRWeN���ڳ,&g7S��؍t�Z����T]���f��-V:u��43�!rn��� l�Dx2WWr��E�7�3�*'�#��T6c
ڵ��3��%'�Î����g	ҟ�U�O��OFF�ߊ���!�.^���Rh�]��Ӕ56���,�������*X�hdi�r�J��3HkY�C�ͪ�����Q��R�ņ��f��b��x��rkz9c�^U��j}=j�Slbr�T�)��-�	n�bo��^�������]��q��ȗ�'�q�����bڥԼ��;ծy����KZ�%e��.6 �vC3��X�1�W�=Y7Qj�FYk3�W^�-evN���1���)g5\��a9���m\��������>�j�i��M��<�>�/�Z��zwf�}��Ǔ���9��-��^�"v���OOo[��{_2e\�&�r��[�ґ9��mά��*�W=�r��2��WW\�O	��`L�,�Gp�k,�(���i*f�c�v~]f�o�R:��V���h�E�Ý��v&�\.*��O��L�/F�O���Q��f�^-�|�9z���Lܼ���"@0��a;W;t���BCe��_�ھ��q���nk�Z27��&��Z N'Ì��B�u:qq�X����܊����}�.q����>��Ǿ`�CI)EY�V�R&���;��[��)��� ���鞪4����2�,m4	mW�ꪳ�Әd�L���j��"� z�F�r��eg�����.�T�2�a��;a����*�;wNT{s�8��E��S��VHjw�.�҅�K�+q�3�ܐCC"�|��k�9w^r���j|�׼H��ǹ��y��f½{�eE
c�%[C4�A�a��xI�N�heM{˞t�2���&Y�ڣ~�s��s�'�KY*c�H�ԩ�cܑ'V�ب���wx��H�F�>�?v�)��Ǘ��`6�`)H��mQj�����k];޴;�C�k�&��؇-�Sr}WjZ�d�,qe�ٲ�3��Ե��y,���S,7OX���nL�;� �V��M,5b��WT;մ矫��O��%�����$7�<CN���]��)�M�Խ��W�Wa�g�u[�m�R�Q,��F�	��,�VmT�w�rC�l��X��v��Q�[��=�Y�z�Q����c�/X۔�J�ꋪY�����M%�:sS��@e!�U��ش��`὾o�v#ŌN��,�S���:��Y������@����~�%pqTqv���YW�T~J��5�'7�;A�����������=�����'#}ӱ+�+��傼�w/�#aV67J��V����2�O�6r�e���Bܝ>.j�JZ�J�B�SF�:�έ�60X�j��y���.�s��^[ ����Iu����=�����TS�Z=;��5��J�ߠ�.�7�����E���>=ֽP�Z���XbS�W���4u]Y�k�n'ur�>_nf��S��8Hv�I��D2�1-�*��&|��r�S����(c�'��Zs	ת����TΫJz:��!�FY��k���[�ҧ8TѻP�)a��I��ןj5j��֫(?�vW��Ɲj�|\�����!>n��۹[�!+�k+2��6�,�T�g�W�}�W�J��9
	�^˴훗��gc*:{v�:O#=�F)^��m=��s�+��<7+@X�e�4Vc��]��]�K{#�kws�F�.�X�Ŏխ���Y{(�J�+�ut)ڦOBz�&�Z�ޗ5���˗d:�Q��e�X�YJ�I�\�
�
�j���N���-�U�W�%��}W��m
�����lܭr�r.<f�gy�x��0�/a~M;��؊h�wky��a�u�pʽq5�L�]M�z27�~)v����ϗ{*q>�?9b��^"��Q���պ2X��^"ĭw��2i������n��|z���p1��Mh��*�QGm��[��L}�fZ�̊V���]�A��P�^^�Kqm����XZ�[\3m���V��͜U�iy��m���T`�-��O� ������1�4,�jY�
�,�{kYZ�+vY��Y�ʆX�����{1+���8��L�ېjv�3Ai�'�R��·-�,@+J-ݩ��1U�i5V'[,q���"��F#O�\�>�Fpz�5��*:<��1�{��>���{Ҩ`94S��,nZ1�A-+I��;YI�4�ySYY��3��0��~l�y��>�{������씌�uT���}�|T�Wp�Ǝ�Ĥ9����-��b��t��x���Zף%h]�pf��)gZ[2���d�Z�S.��v�Iy7��C��U���SL�B�MՙyN���[��)jF��%(f�N��\�������+Uku�a����@/k5����:���Q�T��ޡ*$N �Ō��tn��N�L��:�@.ژ�(r�K�]'EVÎ� ̾x��|� ���Vn�:�[�@�|�Κn�ࡠ�aq�'%о\�K�3�+��k5� ����%:�L@.��{������*vf�^:��5�'�僎w5�.�C��J�)�끮z޸��഼��V֌�ó�v����Q�l�݁T<4qw�]J�F�Z����2�ɺ&b��ܙ�I�w��[Х��e�F�w��.jKl���㦝BB!
�ձ�F�j�"����͗h�k�a�N'�h�T�)�Hb�}�V5.�EBE^nFӥsaX�/w���u�n^(S���O�I�;��5��*zVL�8(́*��ҽ:ԝe�r�����|J��՝�~��n�B��U�1��:�n(6t�h�toE+��@36�x%�c�0�VȻ��K�Q8WwN��� '�eum����4�'.�=�h� s�T� <j��,�����	����]N�u�,u:��|�ը)��V��o~�S�ªtvp�ǩT��C�_*D�v�M �d^���|��V��Ǆ��)	�O/o�r��b�)<'Y��V�kᘆ����h3�[��o�qmb�[��6{Yrԧ���7D=�;���n\��(f�x�%�u>�,i��eL���ӥ<Vfmݱ���5��I����V8����Ϧ7���c�O���#wj$)p�^�������6�����M�2m:��ͬ��˫k����f���m���4t%`��N����s�����w�=@t�G[�aSx�_[0�k����A�ᫀG{�7O���oI�q��v�_��]s ��������A���]唛(�:m�:֤+u.��0��2K�8�w�ݬ!#x����I.�k4�T�y�lncעw����]�4S��ȳ�l��#��O��lu��2V�c5�Uv85�����ix{lA.+�Vg*�aG��R㇗�����֐2��b��w1�=qZES6��N���CD��{�|��Ύ8��["�#��]�d����ĸvf^=M�d=��f�z]dIo$*�ƨC�$k�[��ŏYY}O��3��It�;��[A$p5��Z�5b�й)�)$*@R��;6ui��m+;�yS���G�J��ݢ���u�B�S�cH!�~�v�k��t�i�5�,�J�gK��H�_ow4�ώ2��%�!3M�>�[�r��X�X8%�!<SJvw�V֮�%��)���.�[x;- :Ur� $�8R�;��Ea�#L��>8f�!vw�}c�J�Wv�I�)�qQ=Y�W^>�}����9dR��#��SsÈ�g]Nuv�.eul����v��������)�"�&��X&�pREM!��AE	%DD:�UD1	V��f�b��gUTQ@A%QTSIZ�Ulb""j��EQU4U	4j��UBSN�MTMV�&�*j��b�Y$���
�F	֚�6�[h&Z�i��� ��b��8��*�*�($��CN���ҕE5Th4PD�SI�5�IEUkQ$F�TES��T5F؉�4 �PR�4���f����j *��H��(��)�V&��ZCc����Pب�1�KC�4[�(�T�b)""
((�*�)"�:M�U���*����J����JZ��UQZ4QM$E1S1CI��Z���4bh����������j���߯����u�(��3k7�K`�]��\ާ�Gkݗy�^�Y�ŭ�<賝����K	2����6Q��	Z��+4��]���[��&}i��X�I�QjM��I�>z�en��V����/(��L�l4�8�*�Ա��2��PcN���/#g��~�9m��T:��}t�md�����$o���m��o�J�uu��2��F���$n��N;-�[nƮS�ˊ*�Y�Cn����Z�$&y	ýd���GM5J1Le����,5nP�unsҬCY����e��*�\b�8:��6dB��3��Y���ֆF�1m��eex KU���^soc�>�P���\&���T���X^��,�rn�9e�:�+C�.Pֻ�WW�eX½f.m'�L3e#��n"�,֎TS+����d�9z�N0�,"/q�9�Z��y��X�z��>����x��yǴ��l�W��OC�(���^�מ<�3첡�o�5Իi�-k�+g/<�dF<�4ZyHVȄi�l�E�Ҕ���՗;�w]�T���C��c����&�{X��`h�	`�{t����8��z�U���w���vv9o<�ۉ�{�Q\;,s�Ad��7������:����σ��KQS<d`V��:}��]�p60�K)�b�aWv��*�Ա7:t_��x�i�&�+��M��Q��B��T�9fYe=�&r��W��)!9jl�#ZqX��h2�b��E0f�F�H���e�Yʹ��$���Mypt�I���b�U��y��]���5v��<��Z���i��h�׽�+a�}=���~5����6���ݱ�P�^� ږ��M)�9�B�DJ}疒ۇ�s�Ι���F �-J9	��t����T�����푂Yuu7>n�;�u5Nz�qU��9u��q����9�,�)�a�Ϡ���#�ٲYf˭���A"��9Z�b�ε�J��YhF�^#g���*5�j��k�b�t� �{o��-�Df0e�Y���V���� \ ��"���D�V�s�:���WfT=(���sܳ#!�ңpe�\3 ����#��Q�k0���v%�.UR+�C�S)�u}��#Һ��0���T��k��d�T���::����
ͬ�aB�}����14)���m�r���b����w��= ȿ5Lq�<DE'��;U�E�v���q��'g���-`�<�B�rĝ1oe�ѣ��ct[���d�K��k�'M�����ۥ�>.��J}/����H��EG\���Ʀ�!��!sܾ]9�@����"~��/�ٛ"��*�-��s*�8\'���%�S��3P�-5m~]��b�C��FT�x��J�G?Te�^��hwLw�F�-����'�V�k���N���������&���e��{�L'7{6�ޞ��lIze�E�L�2�,�U��+ȋ��ol�w�t��4�Ku����f�w�H���/9��*��[��U$h�{�Q����)��3��tcc_pi/á�Ꟛ��5�S:��������u1"�Y��l��Id����'����j��S�[/5�Y�i���~�P�ِ��11.���s���ôetf���m�Ǎ/�,�2�8��xU�4I���]5P'��N�1H'���)��{�r�v����
�6_���3<N(ys�q3M�ݾ�ey��X��Ԕ���?.�V������O^�+�_r;F���������y̳B�49�[����u�w.��63�JR�D
Kd�"k�YW�RHY�q+\zL[8�XD�T����-ʺ��d��:Q^����!�a*.*��l�,���n
b%	����i/sn��c��vED�#�ضe��	�Pרc���O;5uA��C�{;�����U�ھ0W�K���v��u�e�Y5<�WS�hL�n���� ��ޗ..9�F��w�1t$��M�m���X;gn���O=;�\���XI��&3(٨&�y�;8G3����z�T�莐�`�t���/b����LoT���MI�|�a�����ջ-��[]��V�A��v]C�+�R�0��]Y{�ٙ��z4�1b� q�\1�G`�q�r�z���t��k���ܪq�u�^R���;��[\�Z�=Q��:*Ye5������>f���;5=.����#|f-�U�Q�4#0�n0듕@q�'��sQ�<�g��h�e�a��N��X:u�y�ɑ	񑙎I�=Q�4���:I�w�퉗�-��%�Y�xe7L�O�)��%��vд��e£l�j�l��>(I�;��T� �5���~�21C��Ek7L�8��}8��E�-���s�h�ږ�rb�|��e�F ���Lh��̦����Dp���{��O}x��c�2gr�$��3����4=��hN�,wV3����k���&�e����CSrǝ�1F)ep�w��y�P��s�1��x]���0���I�卙���}�.�/����#�e�ƛK.�ȟ��Ν���Q�?{�u/��u��[N�K���]3+�r�2�cK�F�� ^-��´�&�P��&s���w�ݒwV7�iT]�_,*�;���-��f�Y�;��Ʒj�	Rt�oj�{�{���͛�����9�,�q�7�w��~�Ѽ�/�3 72݂Z�Jz��B��9���7WW`��Urh�-��q��:n�������ֿ=�x/���$S�t�CS���2�P��Nx[j�dn��u��\�B�5��;�Gp'=]\���6i=�sm����6E�ĥL��*US@n���ͭ}�NY�o�b;-���h?��:Q��ꇚ��ù��y�m6��7_,Z&8'��ͷy{�Η~k��y�}[8�WRA���!���L���=!=�xH+��^(p����Owʴ�t9�i�s>��
ŰPx^rZ�u�F�<�!B��)nt��U�H�n�%Q̈�ݽ5V_ Ѽ+��:ʙ 4J���"3-������P�i�W<�ƽ1��9������(��wγ����S�hDf�;�\�Ҷ2F`\7o��K�y�pNt[�Cg(<���j;�V8�4�3tM���nR�]�c�mxE:}����k� K`X:B�۳U:�m���k-��hKuy����7r�~"�LͿZ.�>�<��D�G=��~쟶������V���2A����,��5�޴�ŧGj���݆�1
�&m>fufnu�D9�W!`�-Zw��MN���c����+�2�����`�d�|�aw�G-̣c)L��G�t�� ����.e�_h s��N�«1��Y!�K���៾Y��-Y�U2�#3]��)oUk�>FP��c�!��f5H��֗���⠥f/��+?�F<��A����}w�8��=�޶{ޔ6+;&�+˲����=���Mo�>ru�w~����gב[�s��N
�b�|��r�w,{g��g-���l��j6����ݮǇ�X�]�b��c̲�-s�ʯ�hb����m�N�7��4���/M�={�,�W�ͦu�t_^���K�,�m�L��1���S+:5�s9B��1���8��|�7=.���e�z0o$�^��Is�@/uy;���M�+�-g~jO�-���y0�lI�AP��OE�D��Q�5�B�H�WGh�6i��ʄ�l���K�ڰ�/H����K~��W��}�>�A��m�ǿbn��it������6ܵ9��ˆn�;�C�F˾���ܴAA�h���%9�e�k��7r���Ѻ6�l��j��3,�E5�y[D��sl����/Z�F;�k:Ȁ�����v�,��N�NA 35Զ���N�P�X ������fU�F��7�:jv
d[�q:9I$�h�4�;����#<����c6E푱?(26ߨ���7*C0Eȍ�WiU�<;Y�6�����h4���gF4���x�vҔ��hic��K��������;&	���!����T���G?(�ܬ�������/�"3-�P�nf�7���=��;�Sgl�2+�k�^eՎ�.a�L�^�/�=�(�x��::���UQN�&�7�f���s.�-Զe
�Q�te7.�vS��z��G$G���1qќi$�V����x������5�������5�'�8n-����p����a:~�*]���HR-aC�������ݾ��z*[r�s�:��	f��'%?O���	с����^6)�D�q�P(������N��'���6ۼu���f�l�m\�Uy=�xk�ܔ�񦺹�U<35��-	ʻ���.m��ozȤ�e�����u�X�Q ���cbU�]t�o���K�
�t��S���z{I�w���v��̨ze�'~�����)b�X붭~蛧�K��*�՝[U��k��1�5�t˾�E�S~=�܂�2٬{kH�ppW��S�6ѳ�&�]L��Y�S
�*: oz�1CaT��ں��_J�2�3E3.�M��0B�`Q�Yݙ��R��!�d��^�ޣ�:l�m]�T����	�j/j��T���ϱX�E
_vɰ�����b�>�m��m���=��K���2��������}�u�e[��ݗ�W��pPe���K䝫kVA�6���g ƃ	��y��v:�Wzf��a	���U�q
�!������T�#�Gu�e�}�����!	1 P�43M��S��f)5Q�(��w��!�k��Mq	�^ʰ��V=�sGh�A�$(��"j�i�I��~r-Զj瞡J!;���kg���H<�d�"k�YEeBM�{%��q�L;'Nl����S���_^�zy�EHAk�*8��"�*.)���b1JX��kv8��Dfe��ʉ��F�m��-�J�޼�z�`�t�0a�e4�=Ry���REd�nE����3ԅ��V+�
�[�ʚ�p��z�Lh�ɋt��[�G���n��~��w�Z�ѵg[���g ����6,�Os���\t��k�����k˲��לZL�:�;;�6�u�w엍�a��� Ҍd�lQϻo	�N��	�D�2��7f���uEZ'5[���t����Qql�F�EK-����v��ӱ�o�&��κٷ��Uswa�wov��Q#�ɗrmD��Q��<�^�s�"��U�K*����fд����T��/D1gʼ�3������gC��6��ټ�ʼCu�V�7ԁr�U���xS�7.���0�a��X�����ms��L�3�[*:=nr�w�l)��R�9ڍ�okR��n�6��ǳ*Z��d³�+<����ץ����N��:Ji���wX�U�O��.4K.�Oֆ	�������z2�5����.���Z�gC��ZT���"9�'ss�ݞ*'x;�Qve4R��Dp���p^������*�̇��T���!\s�
�����+g�3�Ѯ1�����|j46��I���w��(6�T9���� �c\N���)�C�*ه��N�>6g�v{�u���_6���[\�.���$�n�]�hpn�xHn�� ߦ[�Y�O�q���QfهO�ں����8[�G�^eL
n��D��о�%������y��l���S�Eĵ��N�2�P����Y�S<�2�Sų�K�F�9<�̧)`��P[~��}zc6k��D!��<���Ŵ�w���h����
[�Xh��W>h�[,��B�E��7E�l-����sq"ϐ!MХ�m̓s�6�蜧Kh��{�%�}Q��,	��N:Euw}�� �b:�S�#�i˼�gg�Nc��u�;��:ʙ�S��lXPx^rZ�u�Q���v����D;�PR�6z�M���^�5� ]���}p�evv�1��>S��V>va�w���m	O�⁡>5
�*`�t��{�ӹ�9�;��
�1������6�.� �O��4��sk��{R�R�;7��5�T��we�7����g���NX%��n�ح:o�������5�S4���V�`wD]��~�1�9錣WC�����6h�f��N�x����� ���D'��2�����-�Hau?K��x����v¯YMv����Qr�+�ht�3a٢,r�~�en�ivS������K���eAᒯO��~�wԢqk��Q&Ց�9�F�T�ʏNP��]N�E�3���2]�lt4�Ϥ_���"�q���y�ڈU�t���6SĶG>������eh��CWii��-�PɊ�
�Y�Ə��Fw��fI;Sx�wO]�hR�i�3�\c�
�(�9)�=�ﱹ�)=l��-��V�[F�u�˿=���)�f���V;��~�|2�%���hOMy�w��N���w�=���m%]x�0)�eeER��{��(����w�Z���wq�ǰN��c̲�-뜖U};B�C�*ه�ɤ�����c[��:s��ќѲ��*K��آ�@!}�c`�O�fYPѱ��{����ó��du�k�o*������u6�労K������������:�Z�������z�Vϒ��R{����n��ؒ���ݝx$]��8��J�]��ZU�J]�S��ՂJѠ�u"��/lmm��q��"�$�rvN}�. &��k,��Z��=ך�սߦ��R�� C�]��NF��&�a��Ǜ�����Q.��8��Ƃn�9��%����c�����.�#�${Q� �/��f�X� ����pU�j�N��*C��vsr��7Yάѻ[�ҖY�Z��tB��[	bf���.�a�N��4��&R��c����.wt���|H������^�u/T;2i�6���Q��
�e>iDMm#C\t�ݭՋ9�
U�*PUIq��Sl=}M>���~�WMFGN�V���E�:1U>|����|Ui�G+ٻC)�N�򥷪�%5����%M>�fn�up:�,���gi��|^e^����Z>����no������03nlK
� qو�;�^I�C)���LyLw���`γ��lf�[���v�Ahj�3|���z�Wj��[��+HXGI��z�1+9P��&�v���ⵥq�`.��Z�p������uԖ��%���=̍U�n9��sS�XM�@��g����Қ.]�6�]v�]�>�jf�51��݄��g`�/�W!�@��S�{�����cvV��t�9=��﷐�U�^�k�y2e������-��/�p�ít�^���\e^v�a�a��,Ďooe�ls�C�l�]��%]u=XQ��40�^c!�)s�͚iRź�v2���3U┩bw\{�P��l�t�Eu lm� @V1L���ef��h5�}x�;2Q�{&em��@K���k;9��}�Ĳ�f��V�*�cZ�tТ&�f땲̥�X��'.jy��F�/	5�C�\JK����Ö��޺Ɉy'�5�U��8���ӥ��u(��2�9����{�Ў;�� �\�H�ң�L�[iR
�!��
�ӧ[4/��ׁ�$� ��ǽ�T=I������7Nsm�6���6�n�͜�����Y��m��2�eL�5�kX])�	����)�g:��Z�!M\�G )�N+E@/sh%WY�n��dy:,��N����\�9���WA���|�)2ҭ�{�X�5�����5���Չ�>�{�]f���r'zHZ&٧f��	�Ǖ(ﮁ�i��5��i�p��}>�$�}�n�HV#����e�{C��+k8��ߑ3m�D��91�fR1�7]r�/j}َ�eͼV��2���
�78��b��"�t��5`��R%%v���`!qH]�����bMK��OrԬ2��GH�z��^�"��2�����R���e�!Y��|!8��x�+�5L)��2�(n)E�N��͗��h�2�c��D���JZ8R=*��)|UJCV;��l�K�t��M��q����*Z����u+�ۈ:���mw{�GV���ooK��z���5E1-�MT&�Z-5ISL�PD�N�J� ֝i�LAA%IICQ5TER4P�b��bj�*��)�WE!���4�����$*���J"J *�"Z��4�)�"t������)��h�JJ("�JB"�)i"�5T1QM	��iH�Ĕ�iIT.��-�`��bh�������f�hj�kl�IUD��L�%4��,�S-KM,AERR����5M%1)�@��DT�h�!TU���k1JP�DK�D�*)*��4�!IL@UL�U&�AT)AE%R;clЕKM!M[#�������{�}�gdC�S�Wl�2Mn��0ue�X���UAu�]��l�=��L)}�lf�Ōu�;��+M�]\7d�>;�h���N�1�o�DgCS\B*5tt)��и3ԺF�e�i�i��w���ƪ�yԶX�gڝ�ud󹾙�x��Y���_��f��{lMӺ-tv����;��
��u�w��mcWc)-�ᡗ6��C��u�3r�	yj0x)��Nf�V�=��)�9�P�̆:��lv�To��.�m�lbs��y�ΕL×��� ��6K#>��	�5�F�6U����x���;NIp�ݴ^[��K�.��ex!�Exr�)�ļ���-�Df[�ʲ�/������ab��nA�H<�q�̺���e�;�J�C�O���=��.�����پ{�M&�"����R�������.3<�:��s��)�Z��@z�����(]]G�2�N��q�nRMB�-�'�m�'�f&�2�������?(ƁL�(w�[fS.���vxȹHΊ��^V:�����Q�#!?:FGSw(xȞy�K��h;^�hni���7�w��9�eC��$��7Lqq�ݴ�9��^Oh�ލq	��Mus��wE�vE������/��Ӣ���6x$��ֆ(�{�Ү�x;�Dz�~[ۓt�]_�f�tg�c���:L�ُt�+��)�n/�L�s(����iҜ�����ZD̕�Üoaqj�5#�{�
O��t�.e\᜺��8�i3�z���8�nMᎌ�ײ`m2�T���縼� ���eb��YU��u�"��� El��U��\g5w�S�wE�zn���ٕ^��8���1�n:]� ����)�:y��y6wg8����5�6)�|�Χycjs��wSQ������׼�A-W�z�v#��e~�jmD�������k���C��m��뫜2�n�jD��4��{j��gV��ob�38�+�'L�h��rq���w��s���\G�bϰG!�l�O�]=���y��w�������T�\��fZ�(R��_�m�cHw����5�'={*�zm�]x�$�tJZ���k�AK5�doa��MK��1�uL��H��N�n%��R�yj0x)��D^��������BY�2�(�u�#��>b�o�]]\�c$ �:QM�	߶.D=���R*����r"Fe�mf���m��2�Cv��$?t>�@�<c��M�yD(V!�^`�!�[p5��'qa�'���Gh�}sb��	�n�*h[]��E�_�@���.���)�$])V��s#�t)c�/��*��ݢ�<�wYٻ=����L��̸{E������󴓊�SF��K����#z?No����A��Q�׼qd��pSˇY]�q1<=t;C���ٮ��T��]�F�8�O(�e��\�jUۍ��qĹ����ȂɍC�A���X��=I���1n0z"�zq�]^�c�3+/���ٷd��0c9.�x�<2����� ��FrE{s�ߞ�10��\�0��N<�]ո!�]V7N�5�u;�p�gy�����g��h�e��9���l��t׶y��&A�-���g��L����6d*{�3:9��]��k.��zU ��n��:�_�c5�K+��p"��CQa����,5�@����޻�{dfc���x����~�2b�qx]t�s��!=�UŽ�\���̣C��l38+�����|f7]m��D�{�3�-��)��Ȱ��� .͔�F�A��ތW����3\N^�O8+͝��	�%�+g�j3�Ѯ1��H�޳M)��3�S"M�����d����q�h��3���ݧ��}ig�+<��J����Z� �1�u�遽}Y=l�lU�Oi;��}��w���q�pHM� 72݂}f�=5�bq�^�:}�{
2����Ȗּ|��]d���j��څt_�v�.o�e�E)�t��Z��zYe�(k-u���jLݨ�ӓ���N�`밒��9��Y�=[y ��!mfX�u�2�r�w��\��R��O��{Y��V�}�-�F�oqt���#�w�yd�noT��~AwM]\ް[R��}5�d�7����g>�zD�Ma��M[f�Ao���U�ƇԒ���~�|?8��N
{���vں���٤�~�!�l]A�[0��+�5߷�֩�饭�#p��t��&9��^��dK���U�Ф������Q���~&V���M���/����[��'t�Ȁ��%ށ~#�d'2ճ�����[2<ʏѸ'��2n�}<&���������^;��SLÙ�<�@���|ճ����\�d�����
�T��H�yKu^aA�:������1��x0.� �ж:úۋN�����1�M�R^�u�)��Mu`|���u�eK[�R��M]ۈwX&�ᡚV�H���n�>l��r�k52y�GrBS�v��]�m�M����x����}�"�>^@t��n]l)�z�x�ͣ���0)����sB[���]�]��fS3o���Tt�S<�Fu�sTFI�ڥ3�s,��z�g�\g�l�� c��񳙌�)��j�h�)�L���1Be����!��9�3�+33t��*��L}��h���ȷ�}q�8)�G�"rS�i���F3���L�Yh���>6V� A���n�<�&�	m !�v� K���5�z�/����(((;�u��U�m��N��f��oH0��^'3w���۫;�_l"S��n��rwg>�לw-+W9��>ΩB����릹6�������Y�&ow*/a��wzs���F\�64X�eK�=�=5�N
f���	�eZ�l�G��ݝ�]�f7��2����g`�zc�'t_Lm�e��k��T�Ӵ+;���e��-��f^����A����Ӽ�S�6q�V���E��{D���!����b�����S.u�_��9��v
��˭����c:"�b�j���epG[����JyΘm2�w�^cn��E@j:YD�5�UZI޷~�ҦUqa��I�m�%�3hS�-�B�H�WGh�6i���@�4�E��[����؅Wy����pr�.��3n�7��G��/ۚk�+fQ�̻g�C����P�©c��k~e�u�ց��<��ra�7�]҈@$��
m�%9�WN?=�I�������n��s��nVIn���!�[�u�=�����P�Y��.F�w::�%����[��-^�R�5ו���~n�T�gE�p��.��̺�_��lC��,�i1/!l���ۗ�\�v5w�љ�����k�[�������7fT<�)��K�N���
�LY����~|/zj^N�Q�}��*ލ:�\�nj���G���S�k)J��M��!��;Ӗf���l�m�Xƴ%]6��	6SnD�M|��O\�{{���l�ɓ;o:Jm���H�::�
�R�:�[�g <쉧#Z��ۣv���ۣ�_!;N���R>��/�Ց�e��w�lX���[����ӈtf��wU�R���B�d�66+�8V��0���R��Y��>�8!��ќ6��X�&���=]�_�[2��~��G.S/��dU
��}̼�Ui�w�j/��f�_�����d�y���ᨼ��TƟ��b@O(��`ou�*�i`�9ܾG	3��t���!��ӃC:c�Ѱݚ�9���vލq���lҶ-n��0���?C�Z�aa7���fzf[&��p�F�k���L�2�2YX�k�W�"L�hpT��ǘ엹6N��Ѱ`��n�w�=��d�!M��P���'�d�b-�z2�>��J�!�;g")n�@�ײ�W�|Q�����ܱ�9�g=�LH=FZ/�cK$>���&p-pt�5�۸	���g&�pu5�a��b�*)�G����;��[��\�6��{��u��:	8��}98��L۽����6�8��9��s�.S�ku�^F�[8��k�ڙ���{+��f�5d�OkL�L�-�6����B�O��U���GN�;ca����:�Vl��"�f1O����޵��2�F$�оKgr*	S/�͝����2��`�k���iܫ`�{� =���C���q�Ҏ�T'��~�@n,�a���rc��ش�Ft��K.����S�yI'N��(m�X]BP��|Fsw��Ȫ&K���li9W��`pf�0�̮K��1���ٗH�wY��-l��J]���y�G�e[���;W�=
���-�e��	֚9�mm�z�3.��`�J+��l[H��Cj�rl�G�Z�9�͒�D�V첯B�$[wC��_�^1��L�yt�HW���j��.�~5�b���ӭѣ t1�9���\&�4�A��x �]�˨qK�!�kM]?FP�u� ��)����Z
�`]eI��*7�=��82�'�����m��5��:��B��Uuf��b7;v{t���3Y�h�R����e��,��x��g$V(�~p���	��E����S� fh�#�V;��Ȧb��L�'����i��6⥖\e�Z�Ӱ'������g�۸ mZ3���S��^�L�
�R���L��Q��>����L����2YFʝ 1�\�8j:�p�$�6��l��U�s��g��FS�/�g�#��"雦C���6�y���/wr3)_S��sf�:�\d�c�t'xcu��eD�{m1�3��u�X�z�E>Oi�l(ӷ���_�LԢ7ܝpE����n�;�P�@{sl��ٴ�
p���"޶. ����}~u�7Y�tG�=g�=X�w�س�Ց���In�+ށr�!S��	��gC��A�3�C�˳�^��N/�̂<Y1��twW<�v��oV�5���M�sRM�� L��xO�:�W���9�{>tSF�w�l*��:���<C�zG�T0kn��s���dNN��o����7T߅����KK?U�@g���߀������{[��ys�� ����p�ߑ늸���R�1��[�Y�O�q�z�9ʾ������9ݮbnh�Sˮlh��2*x�ʎ~�����^�ݗ��-Ҋ�mw�N�2��y��!,X�%��	�m�U�O`�gA�NWW>��2�X�Cm�HyT�S�؉�q��s����;��{٫���3�B=~ȗDS6��*�j�Ex�#�#=��.�}�3u(.��{"
�k�v�TM^,�|�9�l���L�ܳA��5	�������uEu$���u���UE��s_=��ư��;���U�p��O�پ�n�[�Pw�CZ[����g�p��\��@�r�V;/�mo-��*>��>&����BƸ4q��:�i�CJ��#1�~��z�{�����9H�սR%�7f�XW<��.�wU�̶��R��Peэ�X�熊~׌���D��]J���o��v�S7�J�4��f�x�>�M�zvf�aʈ�	�墮k����W�aR�]"��ĭ�-���.���	];��٩j���6u�ڳo�N�ܖ]8�������>�]��I����V%��Es���2��j&����y����c���O��遭jk{^��ԝ�s�{�2�K`�"�,�ЖT�TP��.�B��~�!��<�z��|T����*����5=.�抂�^��~��F�B|�p�&�_����n,f]2��꾷�Q���k�{��4�9���c�m��ϴ���cŌ�8��N�۝Φz�j{�E�,�T�]�5aꉎ+&�8�ņ�]�pt E�d����	�X�����)��+z�^�`@5+�`I�C�f���m־�T�����^=�wG@,��+뜖T�Ӵ(��n�pzcaSu���r��r��_7���Ჺq����}{m�^�d�7�-��	��n�WQ��5�Oi�c�#xS5��xh	�5uv�l.s��ۢ��+������w�`�m��M�*y�eo�{q\�6�����`q�:T��3f����ں�3f�8��w�⭞�n/o-m��Q�w��y"�T����w��=�G�����E�D"1�t��\��Ɲ�~~�]w�*�fN�0>R��W�n�j��;i)(�<*�j���]���42���l��%ofɁ��ho.��Zw5�W$�Q�Y�vCU�V�S��Ԉ$5L��$8� ��܋m6w_PS�a�>��v��w%u�J*�n���V�I`X�{9s0��;�����7�6n&�C��u�3s�w�(����e�k�k�n\��%8��{�ލ��~a�;�s��O~��)�� %�u��0����#�gd�Y&��Vv^�8y��It���$����v�|}n�U.�K+p�a �"�LK�A��b��/���V)��c�����ݖF��Od��)�ַ*!@{f�/ß�⚤�rP�+)���n������2ٜ3��O����g�a�htSr�i�e;��+*{���$b��w;v����͓!���T��k��ꃂ}�3��`��^;B�S(�jn+��ƵT�h�e]b*3���X�|�\���P:D��b��U�`V9��(�-�����	�n��i���p�՛�v��w��xؤ�_:�ʇ<]�ئn��6�e�n2�-����ލq�s�e@�L�kFQ�{߰�6](������.꧇�+x/,�<�~��0d2��}��>�K�g���ڟ�UƸ�S���22����S������^0&�̨ze�'�dƍ���{�T����(h��t�h͈���VL��pAl�K�ob�{�Q*�ub����/��;�
��64c�S�i'{�z���][�jhw�S�trL8l�H��H�p<�a*�O)��qG�o����e�	㠁}�VP_n�F���S߲�}��#3��9i���V�WE���:��0�}R�U��B2%��v�b	p&e�h֗��pN�'��Fŝ�v��@�{��º��`�j�ҥd��T��R[���\��˶��r�s��(*�rU��h{���Cn*�����Ju��ޠ�+��Q7�-��}Dg^Nޮw��8LZݚ�\��nLj����E�*a��"�{�H�r�V�(�����c@�R�g+��0�Y�"��>�_�����5]č��F\�m�=���yvә�#�����;iιׁ��f���/��.^�-J�:��Ҳ��tB��X�Ǘ��Y2��;�ץc�E3 �`j� 3�mfh�][���K>o7���-�Ջ��sI��5�6�gw}����	i�3hb��s5���P3N�b�9��,��� MKs	�8sz%Qz� <мK�y�~q$=�O�f�_�j�[��J�B����]Y�����T���o��_%�z{��'b��ې��;M��1J$ݴ�¡�]��\[r4����9H��넃�wAۮ�{���u.+*�M�ގ��0�uҗ]���+6�����q}����\)1/�Z���b����,׊�n'��]^����TL)[Z�N����4++i�aw�\p��yX��"G��������E9�) lV�;]�y:Ҵ��3L,6�qF�X�,�:��x�4:��ȨA�tn�W[�H`Yc�w�x��M�8;��:q��.��]�9�-*ÑVj'�8�0�.1K C1ق��h��W��[�O��"t�Q��£�J\T���%i��\�k-�EG��;���j��J�*��>r
H��n��'.���T������Tf����Si2������.�b�tw;n����3�+�:�cB��oY|H�\R����΅�%���b:�i�__v�jQ�@�c^W�±X�m����H�E�M}�)c.�5�:Q�w�ޥ�p��j���ؙ1^G�����[��we�@��2���E�-}rV���%��6����/ V��D�61�8.r�Y�'�Df��nk���y�s�gۀv��(!XF�9b]#�G��72��5��m��6���@0k����m�kN�M�{Eؽ�z�	,���Ӌ �sq౱�Σ�л�(�u�"2,��]����>��[��oL�	�ӫ����yk�D��
"H������j����hJ"X"�(�J��A�hh�*�")bh�����S1A�	E)HPTKBR-��&��(����)5�!b�)(��vD�S� ��h]��#BR�PUV�T�)I�4�UL��4-	B�kEi��14�Q2USB�l���)i(h���E�**JH��(�*��"P��P��Z����"bJ�4-4-R�JRh�Ĝ����K�9�',�C��AJS@SUIM5SIH[Pi)�CmQ	E��P�����ӭU���4�)�!�G!䜓M|����qE�r�F�n�tڤ���&�≒e�n��/*[���L�n�ivt�}8�X�ֻ[y�\����ǡ��m�!qN7�֎M��Y�8X�[�Z9�'qS���[���bB(�mx�m�e���4�/��Vf5�dst��m2_'��X�փ��������)�%p�����㵵8֛Ɖz�{�P���s,ܘ#�d`	��S��F�BZY�>��q�֤9�a_�j��+�C����:z;J�zh.c}Q��Զoi�u����h(��w��;߫��Mq	�H��WR�Rh��n��I=�r�lf�>&�B��
�r-Զk.����m�ut��풿��_�bf�̭�&�;p)�l��4V�APH�ßs��A��̺�����;��!;�E5�'h��\��.��F�٪���$�o�L뎸�-�%�[��.�A�#P�qo��t�^�L�IRxy�f63_$"%;���!�16�Μح�\&�e�{e�hS.��D���!%ۨ��+:s�ތ�ܚ9
`�]e3L�%�o�:�	�OI~=B��Q���v��7����[ꨎ�u��P���X��#n*Ye\�(�H�Qϻo	�af{�S������֪��7_�[�s�<�$d��9� �<��].ή���l��zx����X2�&|,c\��w�U��g`t5����Z��f-�Y���+'��ڬ��>�[s������e]�y�,!ϐ��k�Y*��NT�Yق��X�e)S.ޛ6H-�i�gt��p�@��ȝ����yw��L�,z�(����#n*Ye�Xe]�Ӝ�V�c��Bx�=Z6y���Ϸ�O:1�{���/|�w�����s��)��q�70u��l�('D��͕��-'͒ˁUSό��p~�/5��V�c>FP����~��ꂃ=�z���ޜ�m�Y<H�P������NF:~ȍ����7Z|�zcEgfSF<݂�N?@�5��@�ɻ��r�����L�/�'���p�\s�A�t'|8����tk�ona;N���z�h��sF�8�v��״�Xr�CW,y��������=��7;���J����M��ٻϥk���p)�uN9\v�L�R�1���n�fa>\F n��t�b�ȼ�ջ1��y�a����ʻ���7+��kЮ��\�\���
>����+i��ju1��iͿ��6ۋ"�/�a�c�l¯�g��v��t��>�70�]�n��D?uD�Q�}M4٦��K���n��T�-P�B��tE{{e���A[��텠ut��K��f2���{�%�̶��5J�|��N�5uK�f�Z�pg~�a�O��f�I>����oX��]i�����í��ǺwCvx,��Q��w��𗴲iV��fZ9!=}F\r�Q�
i�*��:�i�<,=t�5/���X�(�� m䙭9yzkc��xWB�u�3r�
S��B~#��	��/k]Z�H5P���qzL�u�?�싧�Z�����-�^����3��ض
�ds��l�i�۰�u���ޜ��䐢���vU4>2�QLo�G!LYS$���0Fe�^���m�;d��<9��'�e&jE2�����um�LẸ=3�å^�wZ'��][=�9���#�5�(�]���R9��~xcbX��K�����Dۻ��.�J��ޚ�h�r�Z`��Y�m
�cVu�z�d9��9p,"�,M	eLȞ�����4(��Lˣ)߰�9\���6K^ne��G=Q%�h�O�y8��p�l��"%�'�&��#[��Ɖ����
�P�q�m�Kᕅ��Y�����)��8,���6�6~}����q�8)�G�"[%;ƚ�ny���6y��Wt]��$�s?B4�b�vM<�Yrw��p-���W^��	�"pb�ԟ!T�Z'��������~j3X�ǖ�;���κ燦��8���'t[t����YX��ɯ#�Č���?�OU-|��4�k���+;���Q3�v�=z!�J����:*Le�׀u�u���k91S��Hw��ݾ��;j�:��N����C�tr����X��\��%�iMU$����h�d����ҫr1yo!V5��
��w����=�.�%M�R�q���/����{�[�|���\ën%���כ�:�Q���v~�7Y��,�,��p�lB|�]]�۶���ۢ�b�{�ق�`,�<h�9o�����z�s��n�i�w�j�M��T5z�8�^��Tͦv��n�j��j��ua]4�sV�&��O6u"iސ��w[M3��1�=!>����GD"1�1M��- ��q�g-
tw��v��+�n/pl�Ф&�R��a�|�	y�<�d�-�C'N�Uٜ�岥���k��iDm��,�����g
eo��`:ʙ�/0zM��:TE fE��]�`Y�M�e-�}S�9�кI˲K�}�_�T����V�!�E0�dd�q�O����P�F6��f[<2�wa���p�s�
]X���2q�L��8��T�����y�\�-���,L��I����p��؅�������W�b��v,�stM5��}����Y��w\�-�!�m)���������b�����1S�Pٱ.WÀ?�}�$^��<���dG��,w �(��<'��%��84iZ��ްI�շnJQ�;�*aX���_����v�z�2�t7c�z�t�����m��޹ݛ\�Ƞ�M��[�"|�aqˣt�;̟L�A;=&�*��h{�N\X}����D��v�/�Z��!%{��_�����|��\��W= ȶ��#n*Ye\�^����8���n�jq=����V�	�=r-���4��a�E����dÇ���#n6[��s�S^Oh<��Mq9.�˺����;���d��6u�fc������e���^��M� ����V6�;m�`����ʫ�ސ9���fpVF�l���T�c��9�.4w����v	Ǧc�1�keF(U��~综��;� �z뜦6������qK�S�6s���G��E��d�`_]�Y=z�(�#���$:�~����y��`Y�Ά��TV�~�m]|��ip$mq<a�TĊj��M�3�{:�7^�Ku�xߞ<���E����K<eZ_���ԁ�k���R���oܷz��Q���*�l��������-�6�#Hw��(+r�o�B&Ŧ���{��Q��y�8�<=6��Ǿa�e,��#�Sč���n��~��]ҿD���&��wr5MZ츛��5Q���c3~�n"k�YW�RH�M�o�C�����"� �ã]����%��j�i "���J�U9���g8�y�*[C�j���B���L9��Ӗ�g5P�՟�A6�*��{��ִ��ߓZiu^����G�o��<��N�y�u#���񷃝AnfN�uٸl+ �S���9�m��X�Qc��F�ٵ;�w{7��~�P��4�S\";-�Y5�,��WZA�Y�nao�w�No�zv�p�uu�3'���3��w<+��!�昇t;Gc8Np^�s!�h[]��V�@�1FX��YSKF���n����T�z�&�B��*d�*7�=���-�{���_�e>��嗖@{��<s�ms�#����7*aҺh@w��!��R�i�x�FrE6(둷���/��=K[������}��כ�?.S\,r��fS���L�p��}3<F[EK,����Z�w<���A�fk�G(�3GM5�s�ї���Ff8Sr�w�z����}eP4�t�9ؗ��ggd��U�w��QG��h�}��NKk���;@��e�X���fc���x������u^8�;�m�k^:F����.��|t�����ѐ�����5�NE{~؆N��ܳ�݈F�w�1\����h�Nh���$�7<�Ys;�t�����2��w��>tShN�,q[:/Ѣ뢺�8��͆��]t�ܭ=(Ƹ�2H�FZ7��Q���c�����i��b0'�e���v��}�Ӈ(��+��>\#[�٦F��w�Wg�;>z<�nѲ�J��),���[i�6`i
��fe<�
Xr��������d���鑸n��7Q�	�k���Z�nE.��4Fa��ɢ�\�S�&�[n�2��J�)�n[Ζ>E>ܬ&,
�M�R��s�%���:�6mk�ϕ����ѯ��ʋ��CS,ǔ�@� ��v	k5)�f�X����0���[3�8� ��w�f>֮��}�x��WO>�+���A}>Z�(R��J-'�A����ړ{�7����F�[�#Z���Ч�_���'�X}zefS�;0���,a������6j��W��Q:��-�='����K�)�{i���Eyd���h�Sm͕ob��o1��cz����h4��
�A�u�3s
S��GXO��q�1]I�� ^H��9��z�p��V;�``��T��d��Ϯ� >��<�
��fk��zOm�^���uq��r�W� `+*Z�Ki��A�˫ƙ 43J��{ �ؗ���"�*�xuy�xN��	��l��86���Wf[C�)�L��-(��h�u�6��FdV3]d�~njΞ���35����<��'�3R�2��ws=�N�ԯ�����t�6Dt�oN�np����0�}|����Ӑ%�v�Z	&���G�(Wr�~"��fߛL����¼\�ḄL/ݹ�iWC4�^�Z���ٜP���y�=��&��q��Z}�:�'wG]�$�*����]j��;9�c;9&vwA�W/ ݊Wu<d�u�k,����� �x�6]�W1��&s�?]�����]TO��6��2^<���N�xaI�͉��V������ݑRa�j{����'�ۖ�4ܨs238����	����������Աް_���k�]�TÜ��H)��^��,&���L�{fFTlW�;&�+̻*05qw��^�FW�%��\���y�&]�t���=�v��F\j�Z���)�w&�w�=���Ǎ'7�UϯmݻR�y�F���r�ݯ *�忼=����(���F6G{;�ه���T�4T�lNy�N��=t_^ٷ�IzY�߿l�xCS6����]��s-��H�2����9��^؄�M�uvn0�ʖ�%����r�C\4L\+�:�nm���|�$iލ����u޷��5�WǢ�D��
{�.���ྻ�)�֏6�]�cY6{4v͚l�r�������m�f��cHyf���\A~�3ε����諱�{w�ƺI����������A�2hR'�Хܨ��m�w�:�D'�n�FFc�%�.�ӛ��6l����T�y����C��uu�P�3�,� J�Yi�r���M?9&.��8̠t��_O`��<~��~]�-�aW����.�}�5���R�p�u�u��̌{�odm��w���dd-��z�o{,�uN��ǜi%W�J�n�� �P�O�u�(Ư����f8����^��9��f-��9��P	w��Q��.�E�vIp�����׻+�^���Y[��	�H̃St��x�
����M��#�r%�q��`s��<2�-��ʽk�_�uθ6����e�:�U�5����f�װ�)ݽ95���r9���=ϑ��ңpe�����=�m�g�pHtj�[)�yGm�=��;�z�S����ú#i��>�@~֨8!����vD��yĥ�x��8���t��lT5�C���L됹w=Q����0L2�s��}�h[�#nូ���*j�V�MoS�6���ڍG[_�C��=��p��]�دt�>S����ֵ��!��.N�Ns!z@�C��c�D�w�5�ΌDps��05tC���$�Et@�i��y�=��(��U:e�z�g{pئm�����S�6���㌧���a�陡��\65A�F���e���J��e�+XV���Z��x�a�u�����g���(���pߨ4�K~�I�e�@�]�t[t����E�����jlP�Eh�����a�0G>��4'������Vu~�Ub�@��~͎i�ۤ��-G�u��/�ss�w�?o+�b�Dl�,Jq����L�P�t커��qk��9�o_N؛�f\�V��:9j�ȼ�?{��л�g=j�q�6M�t-��O��+��݊\��6t�pf��n�j�7�t�e��$/̧'�w�����B����X�ּ����e���x��{vp��B�WJ�k��C�n֙B�LZ
-�m�F���q�4or�*)5��n��Z;"�����B��l�ѫ���]O~1����s�P��N�v��2���OoRT�YW�����]�9�9}���R��dd���)w��} ��̗G�mș���רO>�w�F��Ŵ�{�\e�#��Y>��eM��m�F�m��*�;���e����-���=.�}=S`�~B�0�2�!ႎ���9�w��Z�e�F��l+�J޾�5�4�%��d�%�G�,w�#0o�C��2�;׹4w
`�����%F�Ǳ�pe�O}�n�evΩ��Pp��S�4�0�:��E�L[9��M���"��^�򎽓���O��A�͉i��lJ�Z��X���|��	/��h��'���6/ǣ�����̳��3<A���X��W�s36��5���ǮC_{6L	��t��><�4%:1øÿo2����%�y<3��豔.��>�e��jov�
ٛ�.�yP��pw`�mP��WJ6��t�ͥwd�)4�)q�sp'b�5sn�7�QzS�YI�[ԃ=���fӛV��ea���"C%�����۰�9�u��Z-�a=��d*�1���n��?\ğ4�gy��\�V�u�� �dW�U����5���1��|.F��м����
2W]!h�F��`��K����a�tz�2���8E�߷���T��5u,��ndY����uHȡ.�G���`k��,��t%�)\�֪p��kB�G'i�@�v�E�kC�S'ց��!Y���^:v4c4Y����]�[�>��5��i�D�+X�,3N�L��d}��&I�ݏNL�6'��d�zs(��116ú]�{�p����������\;T����X��qŖU*�AL]кW��˭rSJ��Z��c0��V�vǑ�۵�Ɉ�k-�o^����6입�{V��+qX�W:��ot�$K���Sm$j��ʝ"Q�\{�λ�a�t�+5C�������˚j�!��s5\)�6�]Ԣ���墕.�s&&q+m�� �6�T.��y�4�r��o�7a�k���%n���w�dQ,Uu�;UՕ.�ͮ�� H�i2=��Уz�6��D��&��U��"�E3��n�ţ9sx�8��MguG9Y6ul��D�VV#N;�[Fa�륗Yz�:�dp�;~��q�=4�J��������Q��<���ÖK��-N��盖���?a�E,��Bg���$��m�lZ��f�qq�W+���Q��r�T�3���6�	�|EI�o(�/n��d�qI{s2^4�Yg��;xgu!t�sI�����u�@殩Affj��tw=���_:B�	���;wu�NQ�K�஗`��m^���Ȩ�K�]�����6�,[���Է.���(��ծ�G�"�� �t�|z�����w/~}a���wK=�C�@��x?�<��]�'B�'kj�ɶmWWr�EC��U��l!mr�'�;��sv��_Z���M����W>���v�7���ºud4�76�'��S���WK8Na��L1�d�i��]W�6M˛}���E��zk���:��*v%��unmj��`��)Y�vh�ŹRa�_-�G�u�8p֪�m����-�������5���૨mr�u�wD�WM/r7K]^�7�꜒���5��7p��n��Zq����\^8QC:�D=Z�svV,��k�TU�bTj��-��*r��n��n����+C�����C��պ��lj�,�MfW[f�sP���ȿ��"9�J�F�A;����%�2��CFlWSH�|���V8�SO�ݛ!Z�nk�DRĜb��|����fa6{Uۺ-�ݽ�N�r«/����'��wN�C"�̗����q��v 7!U���C�yqV_4�e�F_a].Vm�W�����G�v+v*=�䓀�s:�!���qUns�7w�=�9��׻�=?a()i�o�/'UH[:J
"J��DAM1�N!�
X��s4����PR4r4EJPX��U�������kA�I�����1kDCM�P���"�Z� 
h&hi"
SZ֓N��[gF(�#�qM4-$��6"k��%4�14�Q�ZB��PUD�R6�����v�U��Z(i�������9�T4�S�iC�)t��cr�k��QL@BSKQ��*b)��l�BҤT��F�JRr,'%9r�4�4<٦&�C�J� �f����Bh�i*�" �h)4hy��T�O!sD�IIAB���[Ji��)ZMv�H[#��M>���z����sǁ��������%u ���iI��f���u��|�^�����Fl�yԂ[�Մ�W]����W�C"�$�FH��?�g�m�?�{_��1*��7笸I��|��Jf8=6F�L����ȋi���FpDa�����rm�h�)Վ���^�SQs�M�?lEhN��n�ۊ���ʷA��v�F�H����g�G3�M�*0W(c��{�FJ{�\N^����F���_�q	��. 'o4����qR�Ʈ��j2�L�����o����b�\N���^WrӒ��f{7n�o�ug;��0����N�&̬��:����o�CS,ǔ��Lf o�-�:����Yv��'���9Z`��ȍ�`'<va��{WW`��<F�+����O���|>[��by���x����qyU	��·��-��YcX�®!9�z�Yk����9]\����'MЌ�c&��z���&v[��!��tJw[�"��)g�TqP�"]M��4Sj�E2��ː��]ϓygy�4rιs�p��ܨ���hR���	�������{� �����ח.T'��z,��g��w�c:����=t�������1� �����9 �4²;�#_X�<J\u�F���Zxq�0�V�oX�T2S�dJ�֜�0�3o0��`���߲��C��I��2�N�mԠ���r-��nr���Z��-��DwP�cUr"�uC�[Cv�ݎ<���!�D@ͩq��5��#�`��P�v�T�gKY.��)��v���۲�kѪ���(���v]�3ϕ�,y�rώ��L���SA�UU�u�S��DB�8�2������^��H:�����u�t��JxS80��,զ#k�scf���ө��u��D�NH��xn�<2�$�z\f�^G*w�"����N�OG,��H���nH�D���X���!��[4��R�Ӑ1���	&���z��{�K�y.�>	�bU��=rŲoLv>v�y�W=!M�O9�qQϗ�n�ד���D�O����#oVhS(nL��S�8Oj�ި�j�h�媫_��#(Sw�X>��-?>��B�,n(��W����T�Q�i�$�l�w�h��(��z�l�lVvM<W���Wx�� ��h�et�=�<�)�t5pq[�i��5�Y&!"9�C����;֞��{�:�Y�\�����G�N��Lg;������¹�,Ӝ��\�ej6F�(wΦه��}�N��s��t�m�t���K�]�ru�x7;��곛�+8P��|.A|�2�.#:-���v!>Sj����ܮ��l���N�Y�H�Y�p�G���1�k�&��6$����"��Ү���a;��Vt�]�
�ռ����O]�2gm�����1�0'��&p��R�O�+$n�'�����{�b>��V �v���_r��:�w���br�N�iZ����'�[0��[.�Dۧ�3n�սL�� �jk��ѨC�ٰ��f�8{�0����;��XxH�;ءM�]qʄ�˼��u��4�����n �At�+6��5�Qyȭ���FhǼ-Ӻ-tv��+�n��m�M*�t)w[s0�-�w���J.�Aꍫ�Ow5��@[�O3l��U��}�S�sF��e�'�����P��緄C�gV���B�1�V��E��1���)6-��
�Y��	�I"�vIp�ݴ^[��K�.��djY�Co(��1����|�� �"�LK�0;*ú"�|�˄�M2Pg�v�q��Ec������}x�m��Q(��~b��Fy9̱2%F��p�fX�<%��q��f7;Ŧ� �ӳ�s��b]i�P;�7.�e;�+��� :#�{-}!�Z����b������u�|y����L��9�O3�f᭻�^'L��]N��:�MS��T��ɷZ��ELٗ�\���Z��ԭ&�6�w��sב�����^6{�C*<�x6+�8��F�v��*2�Y�:��w[u�T�R�t����ۺ���bH���
����O`��L��%���2&A��P̙Ϩ��k7$	dhů#�r��4z��3<��g3}���d�����j!Բ������W�yE4Ȩ����׌܆�\����z�-����Pt���N'3n�'#NtPk�͞�^mQ�##��ٴ�W=����xҀo��/>E༳.O#F<�^$^P���^54��<Х���Z�e^�����dkl�w�t�޴���	������;�t�V��N�B��7,�#GC���,_�ʷ��U���>?)����M�w�4��)���2vʇ�M��ʪ�Շ�lr꽶�Y8AWF=t��!=�'�3��9QZ!���,�]�m��:6�e���#Y�㘙�7D��5v*m��ڂ)�F ��98��ͻ�F�O^��Cj;2e�*+{���ꑽ�ȇRٱ+�>r�ї����Vi�����1�7�H_�Y	O��g�/5jrTb~�mX�����������V׶V>s��t��B�.���:��e�:��Lt��qf�K��A�Fɳ���Z��;ߩA���ȉj�TB�E��i�'<�:�򺺹�>�3�LJZ:r��ێ/��=w�i�-	QqW���dD����[��By���m���L�<�M�����ޮ�R���*B�`�������'8/�Z�e�u�8j{P'���,�;�	�dz�8�ton;������ܬx��4R��H�J�
��(d�.WU�W�@����1��)�%��;����'�Q���}��k�bb��#\^�L�Ce�vZы����Y7B�կy�f%+�=��]l]Ӄ'Z}[�	����6/@B�tƎ��ǖes*C�3rh�(0.��d�(o|g?v)��$e��Vb�U�'�b2��=L�tE�tŻ�e�m4��w�/����Yq�62e8����m��3q�G6tݶx�bf�s��\/Ô�l(���,�X��Qqs3�o�w���u��ŕM5���W1�e'�;`�ݞ|y�b�ߒ��C�r\9��K���w��(��4����&߄����N�W�2YU���m@�l�\%����Ff8=7l��������[�����ݜ՗�z�?Vj^��s�dvK���ǜ���	�b+��Y��n͍[�q��`}����1ۡ�3`h�a�l��ʌ� ��^�FJ{��s�
�� �V����	�܍ӕ��z��:�Wю7�I��i�����CSrǝ�~�cBzƸ�	�fs�%E0�6�^�{K��2ý�lÜ�ܮwyczk�v��.i�����1�򐾘� ������L�[�T"sx��6;�u%�#}q	�[lç�]=`�j�#q��y���|{��\�*��ݜ��5gQ������N��$���� Z��+/�Wgt�Z<�A��m�'���}a
����>�´,�C�nc�z�>^�ǫ1oG�5��	W)Qp��v9ͷ�^Vj��Ac�঍�����߰Xy{}�t�&a�ȓ��i��2t��8WWn'�@q$��_�^~��s�q-n��T�Mb
q	�����^�U�/��s��_n�4�f��� �39��u/�?ݮi������f�U)S=t�u�6��*Ф�Cz����ws�Y%>�<$N[�*���&W�����R��3rХ;�T'�:�!9� ��K"6�f�/2��)u�˹Z���1�=�f��e�|���-������9 �4$�92��z����xb�wY�OZͰ�KVοT)���ݒB��l�]�m*�E1����ZS�}�h��z�i�c�ӑ��	�X���bP��Y\�7E;�ʘ<{��3髃���Ѱ����3���;��|��Ύj/'g$S`\7o��I<'��q��l9K�m�Dۻ����!�FlTr��՚���w�]�壥9���t�My!��N@�X:F�^��^c/���J΂�<
�ՇN��{��]UX�`?r�������E�d������~)��}�?j&؉r�<��,XfL���1�ܴ�Ɗ]3���C&(w� �}1��A3�ܤ���T�ް�{���-V)�=y���:�֗M�)8.�s,��U��*^V밙!�2�VR���(���kA��2_hW`t�(L�M'�dV0�������'>`c�+�<Za��;Q1��ws��S��1�նk Y�_oK�o �ܺ��fA���Q�uP�1/�4d�';\Gx�w��g�<�z��ݲaEgd��.ʌK������ey+��-�g�T�3��s�5��@O�bpSfþ-��j%s�����ξ�g]s��v	ǣ�'tgN5K������|��B����,�x�o������Z��3s��wz�����2�ʋ�Jn���UWn��^ѲB�Yp��L��1�y�5L��#:)�s9B�!>j����7���ܜ^m2�ci����k�Ȃ4�l���)ӃN�սL�� �j��</TK��k��7d=�s��	;*��J;�"W@�|��e2&�}��(��f��;�Ɛ��!<���p4�^�ua��s�ӆ����oMi�wE���P����ĺ�ؚU�o�a�0���g���9wtl�u�w�1����5я�{����h:6�d>.����[>@J2��&�t�./3.:j�Q�:��n 9~��V/�":�%���D���=)@�]rߕѩx���TK_<����νU��͜�9�ww*�LKς���"3-������1ƻ�8=۝�i�Szs��*]U؜�oS��Z�Pp��Q�0d0�"*��m����Ƭ�Xj|�	<��n�'��/����û.�2ԏ����'X`�VoHr�^t���9vp�o8wa�$=|��I)R�zul��ml���������٩�{�~�v�U.fiL���r��=��ңpe�����=�^� %�v̈�ѳ.[��L�:F_U�/D@�a��w];�+��� :#6*S�3_H~��8!�g��JCɪv�3�g�=Z;�hKu2��jn�/�/�b����w�== ؘFkEK,�5�`F7E�hn�s�n4�)jY��X�GK����l�tLL����kl�.Lw{��4?ph_Lqʶ�nb������[;�oԷ���CI�3�K���w;zy������06�tˇ�=bK�an ]�Z��;U�W�zu�H���)�2YX�k[-�y3��.6S�ٕ.���|��''˃@kȠ@�<ma�&��W'�[�����R�dSFB{���c^��B�'|����;���)��Jhh�Y��-�_"����G��G�r4jY!�E���m2�'�q8�����U��R��:ko������k:0.!m���2�,�b����,�@$FE�1�u�?l_s��ʵ�e�y�&�S��9��3A���9�r�#q���FZ��G�ƈ#�Š�:2��K;4i=�P�:�GvhV��������T���X��OU�Dݦ��(���pN�k�bΚ��.�C��|ʍ����.Ҏ�Г�p�k��nM���F�w:�Um��+[�Ά޵�sGaBPpgs��s��*]���נ7���<��T��4�H����eXO^�]X�ۼ��m��Р�}��m�N-n��u���_��om��oU��K �*�}��t
o�,��Wd���10��-�A��.�])�a�:�7��x̿M��p߲7�!�Z����,��ݖU���lkI|�M�\֧��<�*�"u�'�[�:��gHZ��;��9�9�G���$dܳ'u�@�m����j�_4q�E����e�0*n˨uq
C�7&�B��*M�iQ�1��9��{��֜�7�cy�=���O��z�q����iv[E.��:ч�R�kVs�*�Kt�x�$�Pp���6��{&&r�'���9�Ż�7�w���."O�[�)��m��ޛ��If��<�Rەs���Ӱ%�`魞|ybhJzdMT���i�L���!��P��Ʒc�N�S����������2YW�'�W�-'%�	*�����v�K����A��E��oiҭ�G%3�o�LP�E��s�dv���s��ǜV�`����USo�%�z����B�����e�P5e�2�� �ѝ�|������ހ����Ӵ���Aub]c�M[ś�1��H�H��'+��B=]p��;g
�H�1�v���e���q�<P��J�ks���M�5�N|4�3r	AvvЭ�NM�rԿ|�l�֫U/��|��`�P ���_*2S�5��k�y�1>��R�(ؓP{M}1́w��L�n{:5�tn���i��r���rǝ�~�c̧����+�����]�E�w��0���I�͘�[�u������vΐԳR$���p����`�W&�;�����aw��O�F!W�U�t�؞��lأ�e�t��z�|~�j�mo^̪�b�-�Tlu:�2�b���Eĵ���S*k^Y�Bs��U�*m
{�t�d[L��˹Ŝ�k9�������'sQf��)N�#d[�zR�y�G
�%�;�L��4�$�g�#8Ҕ����/`�p�J��2A��8w8��a�Y�Jw��O�v�瞊�iة|���'7��f͝~��H2�c:���	n�TʸG ���!0a���3z튓WiU��3�� ��IS� ���9��t�ʣ�:�:;"1����������e##)��
������L�+aX�0��xe�=A�"���l��yWt��33y��o{����T�`DW ""�¨"+��_� DE�PDW��_� DE������DW ""��PDW��""��"+�@_� ��� ���UE}��"��b��L��GAq� 2�� � ���{ϻ ����6~Ey�^{UC{��q�<�ضiZ�oP�%ق�((@i�*(��    ��CI*�L� �1�`�F�S�i��J  �     s �	������`���`5< ��4Ʀ�4#10 bO�%(�i�т1@4i�&M�$� Bd�LSѣSQ�4z�5Q�Ǐ-U�K
����B9  �P�~$@T,,������?�������c�1�"�*��
�o�@2H��eU@���J��2g�����Y��C����S\c:J���x|\A	c�{<�P���b�b�(�_4�2�"�*9v�+VhYEKq[�R����P��
�%��JÛ���Rݺ�N�bc&�xF�[e\/1���v1Z!�nj�un�,�'"��������-59�%d�J����F�ob庭��Q�͢�
�wM�&1�%�T�<�E��U�����&�T�u�n����W-1j��w��hP�[uNj����������y� ��vҪh�f���N�tC7L�
V6��h�/�z���W�У[-��$M9� ���	����Rx�7��=A���X�,�5�s Z%���(T�J�R�j�Z�}�Ss�͠�������:E=���m$�,��w4��ԡ�	�ƭG��V�5�ev�^�c�T�u臰��bk��:�Yb1�>LMf��I]��3Ze��	f�M)�/:q,��`�4�-&�a�A n�HIo]!:�yWj��=���n��/�BA(�����pdw��3�#bg��x�}nnS2/R�:Bn	�Q�`��\e�e���Ct��Kw�i��A�$�ٛ��VRns'Ph�CY�
F
L���ֻ��=_<z�7��_��|s�([T������0R z�3��Ȣ����o��G)h۪�ꯕ�,��-%�L���z���¨I�@ĉ�����󀔓���� ��* 0�� ��X�(��H��Ē~k��r$=k��M� C�6�h�F[r*�.RbV'VpS-+\z�����)&�, i1r��#B� 8��VQ��.$�	���[��H�0Яq(�L���$S%��43Q�D��C&�ЁA�=BR6� uN�� B�`�B�µ(�kB��<�E�$���,�2%m4�%;��;܂_���J͜|Ŋ�1��x�@�7M��Rj6�p�|��0�p�^�{ԗ=�|~���T�Kb�E��k���U;�1V{���U^۬�XXW4L��Veuf髌�Zַ�EE��ML�;���t��f���A���Fg���sxd���޹�ݨ)]t孑�7Ǌ���OLWo�x!��D0j���Msb�Ql��8㭻P&��hO�ݰ��Y��7��(#��!�ׂ�q��hk�̷�Dy����m�/
�N��I�N�s����s�A&����ʝ§U:����Եm���x޽)� 9��?=����[A��H�f~	2�:ܸuC����/��ۻ@I������Ңm��
۔YS�<��~k���o*��jY�9�3��ㄓMQ�B牬3����/m������Ѕl�c���͢ܙ尔�9��};�B%�6��<#,K"as��oQM"
T� ���I4���  Ȩ�J�VпᆨJ��B�� ��R]璣�K�%����f�ړ}O���V�v��2�7N�끉�3f�������X(�\ۣ���FyqFłM� ��Lr6k��4�ǲ(ߊ�����Zj%��ry0d��ՖdR4k�U���.��g�[$�#o���~6Pm�V)m���E�+|�̜�|���2��*<�B�__h��gT._�����P�T���7�rE�
�:u��66'x�K3z���䛿IN���I��0ۧ.Y1���qs�[TiiԮ������@'zSV�z/NF�6m^���g����<S5��@�t�Y�I��g��x@��=*0؊@���c�Va�c�0�"I����فW�ÌɱB%�l�-H֮ۚq�kzc�1C�U- <i�jpY]�75��g|9n��hK�h���Ζ��Sz$g�'.���J�T2����u�U�P0ƃ��v]>L�_6��,��x`��"60�O^������X�9M
B�_T��* !���P.O&u�*�w����0aNHB:�k [>dqv C3J3��|[6�h��H��R$!�(H�G���n�.��(���[�M�\�H,���X\����U.C���jӆʔ��E6$��wwyW��� i�9�O8Nfh�����Ժ2��� K�f�֙�4��!PICh�v�A$e��.d�M�xmNX�E�kL�	&$�N&���@1�����8����������9Gh� �*-�P�PI��6����xg�I�CL���%�TCyQ�1��-F�D*8�ih�Y�*	#���2��H��Cx���P*$�{qB�%�h��Z&�m}��ƹcl���ks�v� 9}u��)�����/
�B�c�B��#�n���۬5|��U���֘��{���JOL�,�޸wh&nDV)0������ؓKj���dl<�3ʭ= e�^1�̘�x"<�i���g���C%��5�1�r�vF�����ʎ�Y*�(�A��̫����g(�o3��jV�ؒow�����W���r��%�J�X%'�xS�)B��|9��" �H)�o�g��x3�+�����k��^�wy}2!c��~�6P��R�V�^�}�8�7�Nj۟RA��d�s�	[WC.�u�-!� ��.��4 ���f�җx|��a+��ɷw����>a�ƌ�7����3���p����vl����1I�H�Y1E�I1&Vu�"�7@Oc�.4�vl�eQŢ�3�f����]��Ɛ��FY���5Gy��b}�XX:;hԉ{�B�B�HK�ʩN8�6f���I�]�&�2��E�jٓ�-�9XJ�r��w�N]\b�E��.3))9댱�A�U�Y��b���K����v�7<�'��)[E�s���of�� gX��v��^_��|�tխ]��+-���އz��Zg�n�*�9�rte�c��yxLD�rn�a���88�n�����Lvf�D�U����p�s�dt���~F؞�zѲM;w��}�P�`����4^6bW���K�ebzjj�K��ěޓ6�
z�����!�d���@��ȶ�[��cEEI�r�bТ1'��,�եj@��"3i�� &��$+v��nS�UPܹf|�b��[V��" x�P�V�"+Nn�dr�����%�D�>s�8%��Zܞ�,;��.��!\e�C\r��ܤ��*7��L՚���LD�k���4�`���	�A0�]��{vt�=f#K���|2�)����l�K�Z�:�W^>����ނ��%D��Z<�*��SUw/��x�J�k{Ud�'S������;S�އt;&��mdVk�F�0 ��������w��j�	��nH4br�"��eYL6�*Kt�%i[.��Uo u�� Bh��U;�˫��'��uO��̀y[w yʵ�+��^c���s�T�Z�3Rr�`�gK�Q)�͛���pSЧpZ;�L1����u(������U:���@B�{�S�o���E���B����d˫���f��-�ͭņ��&.��8��ތ<�*��Mt�ۺQCr�#e:�m/�]�4Ȋ�|$�sT-,h��"�)r�z��c}�`��u��\_`�؆���5�7z�;v�'m���2o#19�v��s%d�F� B=x�g�k��4}B|U�j�ۧ7՝�Ὄf�u�3��L���NT���<5k.+6���j�c]�4�&R���ކ�S�]-�/�/�����(na̍�6.����m'BV�B�F����݈͐��\�_.�M���BV#1Ld"�X�S؅�K�j��bHv��+k����5q=�N���������e���[��ܒr�nOj��Y�Vde���l�m՜C����d�B$�͔�����8��]�S��
j|�3(��٠ +u�}	����8�nOl�E�N��Du0��$�]9#<��2&���u1�P��:,���SwJWZ:sd�Y�1<�L�|X����i���\��eX-���*���]R������
��S6�48uA�o#�fGE����v���b��z�s��n�,���9�ݡ�26���]��l�)�t⺮������}{��^�^��@/a�2I$�{��DP����<��N�"��T}a&�TƲ)�놅bzr��Ⱦ���,�z�,̆�2gb���8D=1O�~6F�v����'T�A=�8@�k:�:�9c�nf���`/^X^p��͜�.� 2דx���N���	e��s�nY�"(}�����/_k?@ǵTP��hȔ�;�����:�:��/��>I��G����g��.�q|%�b"�������wFH;�m�4_��{F?)���MS�U���AU����0<���i8��g�1V� ����E	���2��Ց�K��>�ݐd!�/$�k���_�g�o��s0�]8�L��!C��1��x�6��\q���(>]���q2���_�����~�����Zg����ð#B"���;S,���N8�O�v��/����P�uge�)��ux�x�{�K�5�{���=�m��3�s:�C��@�ӯ��2?Oy�馍�,H~ģl'�� ���g�DP���i2��/;Zk���p�Mˏ���삨`0r��������~&��f B-���^�X`.9}���d��J�$=�1�%��(��%Rk�{�i`����E[���<��u��/C�����@u���w���s8�6:��<�����Tϙ��ھ�����Oz{�=�R[�Ӂ�e�~�EQ��Q�sA��*�W���}�"�/��c4lߪ}My�~���rN0lq/nɋ�dp-����-�mxq�1���P�< ԏ���'���4����̿c��"�wa�\5����[�v�a4!�QZ�y���Qgي�p�Z�\_f������`������=N}}�UE��v�R@�e�����ن�B!|��g�ֹ��B@}a�B�������]��BB�P�