BZh91AY&SY����/ߔpy����߰����  a5>:,    �р4   �` @2�`  �vﷀ�JQT � 
������*�"�AA ΅J��M"�B�@v �                c�   xˠ=����(ؑ�v�7��h�냬�X�3)��p�:�L�$��=��r'���hd<�r�*�]ݚ��<���+OAЦ]9{�uE<@ ��  U^�l�����5�{�8tG��o5=���ҫ���5��m�.�0p�v�t���[��{�ڴ�Ν
j{�z���u�ӝ�`��Y�Q绅�ʹ�Y�l �E�v    q^�͇l����ws3��TW�;3`i@T�6�e<��}d���	�>�ݺݺN�Vס���\�t�xR�F�   PCE\������SF��rh��=VzC]ux���	ޜw\����]��eǒ�(U�FM�
��U$;    r�Ӯ�;g��U��͏C����Ͼǔ=�.Wx ����{;n�3�p\ƫV{���ǥ��J����P�       �     @  d [ ��O	�UJRP�&�!���  S�$T�0F Fb` �i���$!R���d0�d b2h T��iJ�B4`2a db`R@����&��S�1�M4�FdT�	��R���4�  LF�M�>G��Ϫ~��b�5[a���|��>��>k����$QP�z��K��G� @8T�Q ��?�T ~�ZJ��{�������m������>hCs�* K�0��k�����* pT�eO��`�8�
�̧�����
�ߟ�~?eƾ�O��͹V��l��3O���5�3�m�i\�k�ZzKO`��	�rrx����=�g�f%�G��b{��$��%%��1-57
#ĔL��&A�N�L��}�zb,����Y�nr:YA�]�*"�J=E���$�uTF����_Ϣ�7�"(�F�"G�b0�9�(�\',��$�1"p�� �qW�������g���4G�3ǉ�I!��a\�DD�}%��M�>���"DM��5ȔF�'��b|P�"c�DE�?�B'�'
5�����~GcI)��a̉��+*%�D~މ�����D��Q�p�n!ؔOk��	b;�8@��!�-��Gaϣ����Jn'�&�BxZ���Y��$�Dؖ�J%�Jae1$��H"S�(��N�s�qᭉ��b|QOЉ�Q9��(k���f%��D��DZ���Y��/�����܉D��L,�$���D�bQ3��(����;=	���gވ��E'��_D������'�3�5�*cL#ō\L�_��&�eȍ�gM/�=c1eD#1ed#хt&���,��4�<Da0?;3�����)��C�G�B[�(���,��W�tO譎H�� ����1����dE�Ǆ�&tN}3��bdG���33)���1��x~f0����K�F�Z�γ2i�="�;3)��#�F��oDD�	�;�n��±+�=1���}������\�d	p'@�;2N̓�$�JK�q������?p��{η��o+n#ͷ�����}����[��}���m�=~�s�^����7�ᾝ�0���z���qՔI~�{���g/�G5s:6޽M�}��oѽ��\�����7���1����׵���7ͬ΍���ͺ���Ëb�s�s�̑�Q�*��)�#S�������Q�ǔ�Gz#Oy�|FP��Q��<�$<t�l�_@M}�!!6�;��%�*��)�;�t���N�����A%��#�v$s�w�oڑ���Iȍq�\RG�_2G������1G��f�*�n K���Mv#���#����+�A�7&������L"e1E��/�79��\o7�s>�s�����-�b>F2#���r���CP�7�Y%,DSBU$l�)������H��HG�8NH;�䤡�LDı:؉�$�"�X��^�~N�)/�������t����a�x�I��`��N%�4t���8�(���=	�i	�'�"t�|G�(���D�HD��$���J&�BP���a����"��O"&�	�X�I����ĒT$"e�")���'��NL$zN$�a!(nM#���"y#�%�>B08��!1!9##k�>F8�M$h�����F�Oԉ�$��H�H'	���;�H��)�i�50��L䏨�H�CpG		zh��"E�g�		�m�#�F�g���ˈ�NM;�#��,�HLOn��I拓Q/�		yDp�#����"\'3$�$}�D|%�e�X����S�	��#�3M���� ~4�G"��l�gBa)��q��<;	�#�1�`>�8M�Lb�b�ď�لӪ4J��c�q��0�Z���w�+��G��� ���qcq�>�(�H����~��3	�,_�CSU������{Ǔ�A�Iva��jͿI�y%+��	�h��K��d�@�\'y%!#G�\DȍB9	��腮-K�طW'};�%�UJ��O3�u���L�ǅc��u�ݵӫ��ó	��ٳ�0�肍!$�f=�X��22<M��jfh�"0��L";	���L.��!a<SA5�n>A3fa0� ��d�"ƞ)��F&a�}S�i�ُ�F&a�L"1	�LƐ9"-LOɄ�"9���`�d�I�"�a,@�L�&|�L"Z�H�Ő5&�zcDo�	�c�`����	�!�!�#�P��L".�'�&c1���p��s#���K�bH����f$F�-����#1ǆ�0��L"8�5�AUX��0��0�Z�H��ǈ��L-���L"ut�%�1$GȞ����6bDc�2ُ9 ��G�ɱ��G!6�!��Os1�z55s��b��*����1��P4�k���P���=6Q"DF�d�	#0�śbi1_�6#�I��(f� G!0{f'��f4�I�8I�J�Da��b8�6�c�%��c� I��8ȢI����{�"�L<u	�Ic�e�2H�<W���"3$��L�I�D��'���}9�z4�g�(b8���8o��D�f'L�%<]�bK�!bN�W$�e;0kQ��y�i�;mt�3�L㳅FƝѬe�g��̋γ܌�c=�����Ǹ�#<����3���NLK��18D9T�z�öO�a�c���I�N���b���e�C�0�3��q��ͲjbD���<^�g����1��d�1t�����Ʊ�ى������M��'���4�I��{	Oaބ��0ɊOL]Ǫn>݄��^܇~��D}�_:g<{w���_���,#(H�����3�7��|.������.�k���o�'<ή�k���8q�X~b�ۣ���m<�p����EF�n2/p�8�T{�V_3���N�n�8���;�.�^���m<�pˢ�=Pk�{#1{�^��nq��������]l{����b�
� [8�'��^�g�3���A{�<^����l0zu�5�p}[^���xx�j1��~�z"(��Dr<�8Q�О����I)��a̉��+*&�F�7�G혛��D�_D��q8Q7��J'��ҍ�� �"C�?%�B#��'}|�J%7��Ј�ǆ�'��bQ+j'�[�(��)�i�b~��D�Jv%9�Ҏ~�<5�??,O�)�<�J'7�}w�ĢSq(���Q<x�������Ji[Q>܉D��L.�����Q)ؔL�'J9�8�E��Bl�4G���#ı��Ity��bd߸Y�^���McJ��"<X���#��>��u��Gb0��3TB3VB=i}	��#�"	0?;3ꙏ��g�}L����h�,Kv%8��®�=�[턪��2 nr1�~�"<3n5ؔLˉ�G�2�:D&�LN��舓�@��������#qfD&t'���3&��	��;3)�T,}q�@����|�D����
Ĭml\�dF"�h�l��t�:q�S���Ӎ�����cs���G��ok:ox۵���I�m�ھ�w�n{��h�r6��~m�cs�׸g��=��:7ѥ=O[m޽�������z�]��*��.b��2�8XSL�)��k{�$8���q=�p{��vo��B�O���@�|�?�����U�i������p>Di>&,U��fY�:�;�]��ADm��i��aHE]8��QH!HB��zq�����vg���9��F�n��dtc�k�׹?ğ�b�+�t~Z�����}hKZ�!@�D�n��E�"��s��1�-b^[V��W�%�U�q(x�����`����<����d�}2s�F��-֥mT�@:=�2��I�D�}r�aҟ�e����	u�J[�Vr>�0%+k�Wk�RԴ5�`�L}浍S�%+~�Ik}��ZҔ) �������j�ˊ吝]�9��s^b��)�jR�ܥ k�u歫bߝw��4j��H|zfg�s�c���Wߟ��o�y-u-KϊK�~R҆�}�w�4֭�#���C�`5�t���ա	y"֏๧_s��q��W�
8�;>���x}ɭ���S�!��F�����O5|������9Լ?�Z�~SZ�-��"6iiS�w�͏:�VIܩ���1o�B����-+ʜk�c1�hĥMJ�K^����Լ���?1�zg��cP��)X��jܟ���_��� }�{���uMQ� Xl�$�N�%:p��Ǥ.�SX:�^u<��խ�),JV��Վ�:�!�)�3cZ���='%���A�{���lҬuo%iS�5�\�4g�^\z�vq�9�ٗ_r�3���yICZ�p���R�p<p�$�5ј|a�gN�S�K�\���%�L�<���<�#X%L�L��cvuk�]S�c�@BG_H�C��L!�&�8C�s78V<��>8u��g�h�C��9�:���6L���::�f
`��5��P�)�S��%��	b�ܶ�B���%�5)�_��d]d�X���#]S���>���<-���.�N���7:�^j��!%=-���gOrľ��l҇��m�||Q.ǳ��|g�n��a��4��������df�.䆗'~.	a�|a�.�C~�\8}d����&�w#;���ݚP� 9�x�;٥���P3JqE�f����Ǎf'�ve[�A�[\s����㦖-����8t�v4��'���ʗ�sIx�sS+~��ƈ����o���G9����66e��9_�;?��C�ߚ�^~}B{���8�S�ƒ�Ç���-�[�vO!)̜<�T�f�� �7����6ix��ɸ�s}�4��t���|*S�џ4����y�Ҷ�x�2�ܚAӣ4�9:��
�:a������/9���gwR��s�k0����2s2l�x6J�����i���?�OvC�c]_>D��^&�<At��3\y=$׳��|4���c��S�m2�/
�0٥�l��Cg-�ss"N\��Mkd6x����y���v��͜4��r�Ž��&a ^��c�gM��<1A_rS+����ɥ���&��A��(�ɥH3f����/G�rCK3��f�(����6�x٤��!�x��&�6a*R��&��3��}�J��9�J.�۳.�0b�~*n	Q,͚����ril2�m+ Վ��ml��r�[W^�[��J��4��dS�Oyk�[�nC��嘍k͌g����x��X��(y/'QLkT�)�BAÆ~�f6Q�w��Ό��40Bă�u�מ��Z,TT��>��]tJ̘�[�ӭKî����Mo������7ȗW�BT[Ƶ陔��^�'�s����g���zl��lû�1m�|Ǘ�82��k��800�y?����w��N�\l��H��妒����)hٚ@�)�H�!5ۼ��rM�.���d���C�}���}���]l�B�޻�{5���3ˏ��P����x�N�n�1_�{�s�e~r\���~ɘ��j���l��O�t�H�᤮��g��{��x�O:a߹)��΄��g�����<p]���w�0��t��|=��e:R�׽۞��:-p[)��mr)(B���T�ցE�-B���n�孼�W��,�;��:xÓҔ�-�����g����3�Scg�K�C<�HN�����档�d�ȶ�*qbL�e�2��쌢�4�̌��)N�ȇ���w�}���X���y�9�"E|�zIuҔ���!{3.��ԭ˸��ْߝnl�C��ǣ���2fzpbӻ2�"����g�h\ϐ�6�0:�P��6C�v�3�0K�&p=�IS�8}��gc[P��MKΥ$��˚6p��T��!J���'2M��bǔ�#g��}�b��ˎ��}2)j<����R��!�R�%=�ey,Z�-��G��3��@��$<��S��F�?G-םB}�z�7Sե�j�frgǆku�,����/#J�n�]��o_s��uݩ�_���j�����#��<���T�X��d�q�:�-�� EM�c�B�֢ji�sȦ;�������##5o�RuhBֵ!�BV��K�C��6��(�'&�'�����[]o��8EL�'�5���i*Cn�?L:q��c��Og�y�c4�(���G�Y��T)�	jЇ<�>����u�#�:�L��wvq���rPż��� "9����:/	 C/S����ӣ)����K�H��uK@�����=�=$-�d���T�S[w0/�͗�����sϛ.N>�)���J� ;)��������L����o��w'OO��u��ɤ�ܲ���kJ�i�[���p4j'ܺ��M�{�i3�0���	ӹe�������y�t��l%F]�����W���ǅ3��0ؗD��{\��n~�����;�3'/�3[>90�g��qm����7�./8CZ�Lc�cGW�4���;ڝS_s��,�X�zYc[{���l���n�8l�\�㳆����0ï&�-O����S�/?!D��y��j��=���;�ǝ���{8䌡;<Q�s�)���SIsy(l}i��6��ݵ���x}�9薥�@��r`c�R�����)B:��Kܨ���=���qϱ̫��y��6ѓ3jy�{�~�_s�J�S�ub��=��)k��9ʝ�!/�j�ֵ#R����S���=�k�Q�+��u����ϵ���?>��~H5KyS�Bݛ����}˟M-�FNN�n�J���j���~u�?:�-����ű��G��j�B�w��E��o9����}Mu�Xʙ��N�:��H�jS���g\u,b��][+9�����)o���%����J��J����,yu����۟���|��O�y��8����<;>Ӕ�0wp����Ek��_��?V�^�#��!@jG ~���v�f�]j�Gn��G��#�pF���w�������JZ�=�-���}��̔�����JC�= M�Cc�@<���C�8��x�oj)�9��.IԤF��e�&���%�&Ќ`^<N%7�P��dg���5m9)܀[F%uʶ�㶃Nݴdi{+v������#m!��8����|8�7�܂!�L�{r{�H��;��h���k*��m���Sќ�"�%L�"�T�n�J��f�P-���"��mI�p���7B1����41Fȩ��YE�J��TѦ�$/[lM�L�Ц�i��)��hl4U@�m�41�I�Md�
���%@� Bq���STHviSJ�(��'5�&��K �5412��%Dė*�$Z�Z�B��u��� y�	UJ[�������f�ٽD�U��F�`f]S��}<w�嵫�{ҸN�'���dx����ZW-�!kk��[@�&��g&.b�eL1ܹ�����^�Ч~�^��:�6��঄y��N�*p��y |��,�:�u�:�@��Δ��E��4�1dx�3|M�<$� ��MF�`4JomJklN`ޢ��J��:��"[�Hӡ���L�&�Ch�$�M"��"YW@�M%l:��mcKZ���9�6ū�hˉu�+��o h��CRqN[^Z���5uHq��.Bm�
��}���y��;7��w��Z��?k}��
���������(���;�#�C��������?��}�I���H�Q_U�u~�C�����2���
��0������VUyU�iV�W[U|�J��ʪ�������Ȫ��J�]|���Ȫ��*���UmU�j��U|�jʪ����ȫ��*�U*�J����0���*�⴪���G�DA|G�Dt}0DV@aR@,`�B�(L �!E%	�S`�2G%
a���J%�J��JVeB�H�}^���"> �>>њ��TUUU�U^EUUU�U�ZU\XUQVWʶ��+J��[UmU�*�*ҪⲪ�����*Ҫ�ª��*�⴪�+J�⴬���J���U�UŅUU�Z��[UUՕUUEUUEUUEUW���D����
�%R�� 8�2�h�Ҏ$ ���C$��*J�a41-�M��uYUWUiUqV�WU�iU\V��UuUueUU�1ZUՕUqZU_*ڪ�V�[U|������U�ZU\XUUXUUTUV�Y|���ª�����mYUWQV��VUUUaUW�iUqaUW�Up>���D�}�s�S�a`14&���������)u��Q }����">�������ϕWʶ��+J�⴪�����
���XUU�UUTUUTUUy�U\y�UWVUU�iYUWQUWVUU�iV�WUyaUUaU�WȪ��"�������a[��EUUUmU��V�iUqU�WQ��ʕ��� �JD��J2��L�B��"j�J@�R�JiR JAu9"����B�@@.�� �5�.�r�1MK��I��@RPR�I�:�>G���ؠ* C�����?��@;��1�����G�6�{m������)DR�Љ�":G�DI�&��"p�xOH�!" �"I�%"X�"x���h�i�p�h��p�H�'��`� DI,DDNM$ �DJ�$��H�"`�%�eQ|�"'����& ��"'�H�D�<%�YB"Q�"I �!���	X�&	YƜq�p�rG�DI�&��"p�xOH�X��A<@A��2���Py��nj?BۦK�)�rDӵD8���0�
�v7B*�v�-�7ӊ7��MX!	�j��5�Qf��]�c�?=Y��qH�b��H�U�;h4V�UcH��+L ��[�]4�jĊ�`��V܎ЍE\#WC��u���M;cr�٫���V�	h����UHX&�@�G%Պ4��KG���DT
7#���EcUUB!�iQ,�:�q�B�D2��1�m��H�`8�@�iP���b�؛"8��dM��R�����T���**���ET���.��sC�J�ZI�[cqO�q���R�!Se�A==IuFtet�)dv�H���QM9--��f�-v����	S��[�+R��r�jR�Z���B��2Z�?G���<+i�(Y"�YC`챫*�n7
+�t**uD��b�##���X���>Ř*�:��ju��A#�AFHۉ�
!�C�El�5�Qf�Ƭ�W��V����R(72KB�mS
�v���@�X䍳L5uc)�TVyˈr8���jR&ģ�ѫ@N�q�;el������f�
84Ĝ�"龼0tz���X6�`ܖ�T�mU�i�Z�B�U��`��+dv��'\��Z��+ch�����j���*�|չ��Ѵ�%-N3RD�Ũ�ѫ)l,dM�h����)loQ̔UR�M15]��H��ԩGFX�v�,��H�N+l��GT�KZ���ldRJꖷJ�M474E\��"X�+��@�Lc�)UP�c�L�R��h�ԓ�-X��;"�-���Z%�E��t��;��%��O�		cjʝ��H�u4UU 뤨e�1�H�u%NF��U��8���V+��A9+��m
�D�haC��#,�2�j�_\��VW��1YV�de����nBUj�N�X6�-R�4�l�QR��H[b!K��v��e�UeJ�k�M���l��PB�)+��^�UC�%�8,jWp-�f�$�5-� �d��Z@���&)%T� ����T��=\�Ti:�&䔪T�Cm�5D�i�+SVj���X�oD���c�&�h���:�m�;'�1y�&]�+��[%R�7mj�z�'!D�cm8j7TvJ�CQ9b	"��(��X)E(8V�D�5�Z�������,���m�ț)GYn7��dv9SqX
RA�!%m�K4�tR��(�ș�4Z��H��#�����P��u���5-�J�ӅoTC�4�
J��-zl�6�
+$p�����Ȇ���jJ�h���K
�n*�ad �#��X�r��UZT���R�ψ������B����i#���V�:�I�7���^���Y)eU��uQ3��:�QU"�J����E!$�Tq7Z��llqR��%� *�%�iF�+UV���U7"i�QZ���T`:�Q�ۢ��&R���:Ȃ�,Q�V�����4Ai�-ڦ7&�l��[L�	[qW�T�
)���k�q��P�%tE%N��H)X�H�"��I*L�7^����YETb�:�cѪ�
�Gdj��IdMW��-�W	@�Gk�!�슫�*�Y �+b�jB;\�e��4'(���d��k�$h���Z����Z�P�
$[I��PZ�*jm�m�-q�+�,T �jꨪ�=I5a4�U2+h�6�h�68Э�NH�u�5d#��Z�@��Z����a?VD%G�_����AȈ2�U,,m8�`���AV�#L������r=ZA6�:DA,N�`%q�+V1*YVX��E)e% 	i�P�"����'��@Ӎ�%��4�҅i��ME��T��&)��f��G	�]$���"���e�:��
��z��R6�au��9#m4;!���Z���&���(�\�ZJ�����B@��9�F�J*JڎUT�T�p�Uښ�Q5#b*$uUal�W$�+$T��퐱�Jh�8��;d�7]2�Œf2<�m�N0R�!I	Gli��wU�e�F6���j�*��R������0RX�j��H�5"R �vZ�p�4�Yd-�ȡBH탱Vj�	U�Q@���X��ՁAUm�R�.��u���5��ݗ¶�����4(�jW�Qdl�2h���+��7q���7��*�VSN
*ۉ�l�N�QE[�$dN�M�'+�RTIilc��!-$��2V�P�*,Q7"����!2��{���-T�f���DU2$�׫X�M��Ek��Ѳэ��
��KEf��V�k�i�TL�u�QA&�R��Y(�er:+Q"�M8�;)MɕLnB�b�j�p���Nڬ!H⨱ȣQD!�+R�Z�UR��Aت�D�lQFZUm��鲀��dtI���Ў���I%- R�M6(Ac�B�!j��dCM��]	�4Ǫ���"��cznB�R���I%���]lYQ��F166ܬP�@Ke��m
�dT�AJ�i]� �i�Z��,ldu�Y�NH&�!Q�Kd&��`ݍ 뵍�w����_s��}�x����*�wv����YU_ڰ��Ȫ�������VUW��*��*�wv�>��eUjª�"�V���1��YkE�����~D�,�4�8�0�����"!|e$d ��KYQ�Q28�%q�(�b�[N�L��U�IZWP�qAH�ݤ��`�XJ&���%@��akU�[�+r2M;�d���X�U�Ei%c��H� �v�	�f�4��mj��;%j�e`�K#��!*���Y
"��FՀ���(Yu�В��u��"m�j��+�*m���.��SQ·U�=5YZ�Ƃ�X��r�D�V�n;ب:NG+aa�Z2�pL��Vԅ����n���j��`*�%�ƜJ��t��F��-:@�dq�Q6��i,�����N:B���lA*V��TTjJ9� �Q�)"�B�A4�msR��6�멦6�q��N�Z�RA�(�ڲ�ED��5�[$�֥n$�ڲYu!m��S�v�%c�-�6�l���+����l	��u��*�&	��!�!�Ӄ�"��A�DՕ�J*=1n�e��cQ�T�.�� �I4��UV����)�͵����ռ�����&�ʻΗ6A˾�����n�����3w.až���"��:)#�Z�ɗy)[L��5ʞ��L�u�G1m�>����a#���Pf�J�&�wU�nnn���6M�h2;���?��c���Q��T:�U�r����6�,�k�Y�͜v8�mb6Z�xf�Yt�Qbg6�cSJ-�F����`;m��Z#��d��Yi+,`�&���
�͝U��{g	��/F����EDzfp����!F�a�(҄�?��0DN8a�d:p�͚(z��%TO���BoM��6��c13�F��ƨ�{j���v���`6��ci��
T�xh�ǥKB�խ�����04�f��h�����i�Aʨ뗩�|�����oZ��D[E\E#t�F׶�e��L�bڵ4�Aj�h�GL���Ͼ�"�8|�8�O�u��S�P�'	��'A�{��@5&A12��Ѽ�� #�{�G�tɎe�J�.ǽ�6&h��Ǭ,�E���H��%H�ӣ�W�$sQ��h¼�llcb���#f����{�$ɭV��5�u��Gb�o��]�C�G[kze*ё4p�^��xb��6�n��T�4]ר.�$m�������G$��X�l��l�u�^#;��m��q�^S�"p�&@�q�Q�V�0D�GTce�6�m:qm��r��EP=*��@BIEؖ���"@s�^��rY�#O,vd����9�h�F�mp��6�R4X6m���h��b��t�k��i�.-.{˼��[���.��˺�I[��oe�#¤yx�k��O��,�Q��!���GQHj�ٍ�k����0�e�8~0DN��H� �
;�^�����9&�����&��z�����vu=�2�` 	�w݊{�#��nm�d�z�P�n�'<����b��n���.��}Q��n�������v�Y�ޝ�j��=~���oI�����3���פft�wۖ��p��7���4�ny���]�������س.�3}���O_.��m3���7.u�!��ͭ����i��.*�IUt:��;!KH�w�V��#hz��{�e�)ֈ�I���)1�W��{�h
�u�R).��f��{�喤�w&���k��E��,��5�Y��� ��5��3�L⥵ѡ�+E�=�֢�:��E#gL$�94	bچ".�մ0,:�Q`Λ(�G�4�&��p�iq�aG{��"F�o��29$y4k� ioOJ&DR6l���UEa�R1tj׸�v��x�H�yu?�!�C�KH�<.[m��/<�J�Z,,P�]����ޥ���N����qJn�w[M���E�cm����7"������7�m8up�.�6@ҳ��6Ò�E|wq���<i�(J�8L)�<�E<�:�H̃)�I�UM�+i
i1�r ��6E�N�WVFf.���`����^��!�,�H�m�����(�M]�&!�\�Ԙ�\}�e�*�}��nm��/1�n�]S76�����kH�C9�H���K�/����-7~�ix�.��>r�ٛll�8�R"T4A��H���)ma�0Ã<aFl�D�`��'	��'A�na����e�^ۤ%6���dL���UQ��@m���I�h��j�,�
���a��]�p�b,�rg�ydN]U^�ɹ�&�ͨV�R�D8un�c�kz��e�E�Эy��nR�R�R5�٪o!T��F##}n�YC�F���e#J�KP�h�L(� ���ѴCI7}�� h�<YG
8��D�8M4� �
�5YJ2�2o��l	jM@#q���<9r=p��	����uX�W� ;ܜ|��;9��8�,3t���a�\�Nl׍&*�����=J��2�;JƱd�5��VQ�D���G�y�w�Np��wwow����73�:#�q5�3o#���aE������E*cj�T:=�y�u�A�m����Oi�������ͧ���b�e�TJ���}�1W�+"6��]�C9)�����1�TP���co6b������U:�U��������ccl�{�]ѻ�7d��%�C
oiEž��Q��k��E�l�<�-T�.�Xmh�Q��h�j���{��`�[�ֵ�u!�w�3C3om�:����. �4D���ݑ�	���@A�x�(K4D�8NM�4Zn�%TTht t�+u�g9�<.����=��6h>�s���Km�n`�.ݮk�����^h�h�1��E
	���ǍyXE����E#h��ڥ��3��L�co2bu�L�_k�`�Mp/h���ʲLCG�Y�Kc�4�8�pi��B����2�X7��qh�b��y�*O��Z8�/2mK/2ٶ���Z�:[V���r�Z��[6��6��eųi��E�%�����8�x��5%�����̈��G��E�1�>����,gőY��0���o�������O̩G��L�L�i�Z�ZRZ�ZR[��ٴml�y:��e---�mlی�---)-�r�[M-4�F�ͣiih�8ͥ��SV������N�l�-M���;Le,��6��3Kf��f��ikgn3��ZZ��ٴ��Z�)���KG��R��y�-��m�M-�&���[L����2�Q-"Zb%�E�GR&.LE����E�Qi�[���Lul��T�4�O=�皥�����s-��V��6��g�f��̖����V�dql�&��b�1�.Iųo#+H�m3C0g��2�j���s�e�^�����[����~�H��6t�����8�Ng����"������*��^Yf)�Y���a�G|8,��{������w�]���3�;}���ӳ|��9}�Z�\۾�1���..\O��˙k�y������Ý�s=��|x��0��{7��e�@�gmBo1v����^��Y��G�r=7�5Yq�_y�2�Qs��#}�Y�6r�k����QW�|��SV�x�\������>����nfrV���3���9�'�s�?���߿O�U�U��D|}�wwWww~���~�߿~WQV������wwWww�߷������߿:��UO�㻺���~�Uޮ��ﶪ�ֵ��0Ǐ<�<��8����D�8M4��i��!����@�^���fU�%fgQh�J�Q���mQ�A�S�Gn�~$����q��ܝ��:��5�l��}C�'V:]'��'�V�`�$�d�I.`xA�C�ن$v��'����FFE��]i���,����F�8����n/��ݠl3��A��=D<xs8�1�!�GRn9LHMmDj�
1C�\D:n#Jj�ɤP�q��
؊��̔�4���"C"
g�C4|v��#��]sH�m�!�[�����aц�+g����Z!�f�YI���4�>|��)���Ǟu�^qJ3�N��F�㏮3�˧y��7e;���j��#r�����@��K�z*K�I�U,*�ln#`Ģ�lbP�!Fʤ|��7߷$����v[e\�r9�m*C��C]e��nA�B�I��[kcs����z�h%9 ۊ,W�]1Ľ1��D5�.����71Z��b:���V��.����R��*u�]��c���7�a�}�3A�I�A�	�&�ˆ{����%���R�la�6�4w�F��Q��Hz|LCbS���X4�3����:��|�8�N���?���8NM?	'i���D!Ƞ�GE���Y�,���f�mm�m��M��8�4�$�� ÷��z�5�nժ
�ћ��wϊ������t�Q��o9��G����f*�����=}^c6�{k,��ͩ�����5ɩ��2P*�|{�X���w�_6��*�\��ڶm�t���V���^fw{�ڌu�
�Y��
�������0�٣��+K�%&1��h��$���yL:M>�'��a�!�vm`��v�|;�w�.�ӺiB#�����E�8;��24�-$���鍚Z,4u1x�R|����W+H��9��ZXaA猡�����F8n�,zb�v�n�=�G ݗ�<��n\�$0tA���Q�l<M
x��#��!����>��R�����UB�.�[-�HM��'�Q����"I���x�+��Hu���C�q��Jd���rh6^p���(�4�
?����"'	�i�����WI������r����3!$$�� ă�T"
�@�q�F� ݂ �L��F���m�&�$���e�_�/�Ye�#�	�(����qkK��a�L��u��t�D������ˈa�`z�;��D�C�',��,��H�v�p�8$��D;$��޸ �_n)*�G>rq���MkZԃy55����2Ht�g�d�}�c���x٤hC�����	N�؃�GPu�S��pFI(�Aϵ�:Wxi�����gJ���G���L6dč�N�G�n��vNX4�7LY/	��I�Q�n4�K[�8�)�)N��y��:wR0���
�L̈�E�rD�M����O��rR�>�[������h��)� ��1@�� �P���} ��qL����GC��;$� lBv��!�H����<i:b��0��a,n����X;KFU�`$:$�;!�/1���K$�o�y�2P����n�UT�v�r7���u(��)�I2���&��u G{f�;��bvC���m噣iJC�F�DQ:q���;`�%��p����F�U�6_Izyq�b��:��F#�o��%S����bF�X<$��l���I �%4B<���azUH���e(�BQ�<p�?��m<��)���)JyJS��y󬻢I$cs�ׅpBŒKHkh��ݴ�M������Y�$G�5�؎������͏\1_HN�}�e��1F(��a㭌�)\-���4%T��tC�wU�G���h\> �Ɂ��p��j	B8�IӆӴ��&��dQ�B�-]�hg��O��iҌ$� ��:�lA��'c&�,Di0�4�����
����Tn��[^��F� ��H�m�*qG	!� tK�x%؇�]�C�8	M�]���4o�p��pa��y杞��4�$���!�S��c�p�h�M8���??8�)�)N��y�[β���SsR$i5�NAE�L܇��̝R��h�{\�M��M����ת_w(ɝ��.�0��^�[�9����{�ٛW+�L9�z�{ο{'_e��O�u���=i9Ӿ�V{ޗ�ӕzZ�D��A������{8g{]]�{�L�C�$���ryy% ��5�7�]{q?����BNϡ#� ��ΰ[k�Zޑ��C�z��$���s��޶�4�&�:Hhߊ��,3e$��
��09�4�"�F�@�l��5G��w��8$7ަ�ܐ�X�GG/��SI�AG�DF0��μ�]��wN���ٰ�߰4��Jlư��h��yR0cF����2HqTA�dN�Ej%�!�3H�Zf�<&��������(�������0v|��{��T�Ӿ���<܈��V-�Jn��b"6�T�������t�Hf�H���C᠃�KPA��n���L6e�uM8�������<�:l�ќ83����MݎG1Q1۶�Ӑ~�ʄ��@�����q�I�̀�L2�~U*�E�J�h�k�cc��H���6]�:F���Dlڹr��A�+k��'	���8N�4�i�H��!�ha����Q5�S��ET���`��E�bR-R�0�"),a�zIA�}�=t{5e�h��Z���#�N �h����-̝�1d<�n��x{��y"�*+P6��`��������h�&�������N����k��oX�ϛGiM-O���R��]R<�:�Q�ϱ�\Ă1�� �U�)��F�̫�BF�i��B]�b�7"��%P��sZ_n�9$����Æ*ٟuH�"/�qao�����{֗����]���wc�M0Da��ɼ&��N�9�h��׸w7$핱���4��V�}��o��։�Y%�D���#�dC>�=��yE�@��P�h���U'glv��E�����P8�!��#�Z]>QuD`B�"�7
G�nJ[6�ų`�Ba��	$�#!#l��Dh�ͽ�6�.��Ɖz{0��J]�F�vvh������"'���A��H4���"oPH�n���1�bM	wH�R,�I��or6��Z6��7�e����
h��QJ�N��#e/�:��i�pdF���zU��5�wr��[8��H�(���l�Ŵ0cB$��˧�O����p7x�Ӑt0-T$��к�X5����a�����</I�5X���w��h���h�ڀ��ӱ�)��u%*3��i3���ϖ*�#RFh5h�u80�Sh�*�ȉ5�D(��y0<4��r@rc�0r�>��L����e�-���^Oj���q
b8QP�~�����~��?���+�ųimf[6��eo3im3KkS,�E�im/R٥�֙��fE�%����ˋg��KH�E�Ix�b�&�ɋDKH�E�(�u6�m�mm4���h�l���iԥ2��e�-����~[/�eh�Z�ZRZRٵ3�'�������[V��6���J��ÇOc(e'����9����>��|C�,�<8?m��߉�E�ɴ�m1���eim6��--<�mjjѧ�Y-l�il�[��ٴ�Z|�m=%�Դ�:���-Ki��t��%��M%��%�KDO%�E�F�&.I�)h�nIi��e-8E�:�Y[*s2Ry��3י��R�je�H�m-��[+N-�KVd����2�Yql�1�i-"Y�%�I��dZ������FH�9��ŷ�ekC�����_��{�_o��X�ܻ۱^�Ϡ�sur{k���s&�},Xh��F�q�����.�f��p|o�y���_�9��o�m��lߡ�/��Ϲ'�$q�o���k:���ml��1�ݜ�l~�(/s�:���1�9�ϋ���Гqs��껳��W�[��8C$�im�nO�~vv���\�<�'�=��ϟӞ���ط�������e�S�o^����o�K�K�~�g�q���+d�����O�~��~㻷~���0(柕�w/�b�LY*&@��b�ӆV�ӵ��/��mx����2��?��}����?���O�߿~���߿5UO�������ʴ�����~���UW�ﻻ�����*Ҫ����߿UU~Ͼ�����߼�J���~������9y��y��[�R�R��G�B��q
�b[�mE���Zq[@�[p����bՈq�#����vD��bl�KJ�M����q���R'D��fdln�J룖A6ț�[rZ�&�m���:�BWGj�J�q�X�**Ied+%����FG1HH�:�h�)�V�Q���j�2��Z���m q�����+�6���W#��*`A����H"�B�j�]d���V(��FJ�!��RZއR1��U���T��Kf��(��En�KD$
���=K+$��[k���VR�KkTr�#�PJ�N��A�S����Ȧ�518����i��,MB)X�D-Ӫ�T+��N֤�Yt�M8�T�Ye�jX����F"�#tiG�����!�"CH�+�oM@TW[j]G^�`WZ�q��U�B��2B7,U���
��Tr��

6E.�1B�-f�E5���n��nT�PK$�P�EՎ�8��C�V66D�A�˩buʤ�v�W#N�%�¶Z�R8�5v�c�$Б�Ǿ)=��ٿs��oߏ~/4�.���>��I�w�y�2<���'8�x`�2��Q�{|{�Y���H;.�G/h�o�1�ٗZ�zu��ә��E=&�-�9������۪/k���j�8�j������F?l�l�=�|�����f��K$8fru�.mw�\���a��9'���]n�kc�è�aֺm1+TP:rQ{')�;фƜM2�@Y�*[
�P�FD�)��>@�r����v�2�kVf������lM��"� ����R#MyP�d��p�&�ɓv�l��"��ŮKcl�s�Qb<h�5$��t���&;�'���!+�u�8���ns~!c����[�!�)��wN.�0�Y8Z8���:�x����0��c��$�I0�sZCL���?4��[�R�M8�OƐ/5%~�����<W�vYe�Y$�u>���RA m������h�1��F��ʑgȈ�CD[L��rN��uv�*��w�D���gB�5	1)��n�H�y���hjD���Doٳ�&�g`��v�o�Q�Ȏ�E|GV��`�
pL)��C���#F3φ��F���m���A����{����2۬�ְ�񶎀��,yL�r�]�vP��Z"[���8��-1!�ޕEQ�̜p�Ѳb�b;�c/.&�n�=&.j��Ǔ|��I����:t���G��8"&���i���G��L��.z���� #L�-R:�ګ�1��`n�&��T���M�D��)@:t�#��}拪�c�I\Z��E/"�Ǩ5 �Hb�n��=�p9�|��n�0�bx�}d7 7ч���^�V����gn�H���u*sf�<;=w�/2���Lۈ5��Z4��i��޵i�Ӡ)9��'[�&v�W�|ma�����h��KK�h`iR>DER,����w�;)`�z�q�e����!GU@������.��2�[ɤs�E9��)Z�!��7�LAc	���2��1��#�Q�ұ��1�e�Ϳ4���8�)�"h�q�~8�`�8����ww�X�^}q�q�`5�A�n�A�ꐒh,3� �b1�����ta�ҴqQf�|�����ڤ@����#��'�q�UZ��c�tc�e��]���hgEȔim2��s��m/:  �I/�n��g��-Ù6c�NH6w���ݓ#�^NSmI�6�D�0w%{1p]�N޶�va�l�4[c�my���D�^�b`�7g%� ے�M&�lA� x��p����d�0�����$��:�����vz`���M�����D���y��N�X�š�L?b2�&���)q��i���~qkS�R�SǞG\[X@��K7���m<�Ǒ�"�N�����U钫��՚��p�3�X8�>=^Ã�1�4%��߾��7�[�[���ǟo3�Q|���1G-��^�{���9�ʸŕ�*�}�)�ލ�SV3=�{�.�3g�|���m�F{~���ɨ��}[&��u���;פ�����^1�{�xs�6�֯
�ݼù��|�$RC9�H�����e��LNM�3pȪ��HHz����3
�8S�N#d���rBg�.I�ާ�x�;H#RE!��"%	��ܰ�FҲG1u;��̝8���Z:I4� `���rG)X��I��-4q��|;oL�Z1|���rۡ��Z�L	�1�ќcM��°f��91�+���:���å$bh���f�#Vp�d�cH���a�0s�Q��,�ִV]}7������I����7���4{J�������Dq���KA���%�r�6z^F&�o�EZL��w��Sn��>~~qkS�R�Sǜ�G�9"F��-�N����Y��/H���n8�8�<�(�"_��`���y�*A���M���.���$�z0���Z�>�C(n�滹�lTjS����h���X���d_�4��K)�MD��0�}��|��='�]���zɝ$q�!��(��7e"��Fn(�CKc}��Pf��P�R��9&&�)�����Cd�1�#� � ����⠟��o�KF��h:0�=�R�<��ۉkC�IE.�a�=G���Cbc!���#�o6�k~|���<�)�:�WP��Qs�����K�����fYd@q�2Ȣ�3G[��<bDf�|�eF�D��pn�l�$�iQ��"8��0if���ѢZ"�$�FE\wIav:+gssD�	.��c� � 﫳}7�G25���d�|؆�Cx�7z���v�d�_*_,�0a�|Ź�kD9�]#.0rc���$%�ѡ���o��SZU{,�\!6L1zI�$�0��NP�PaH������f5i�CKb�����vKk�H�v��4kQ������'���]:zH�9%44hc�,��hc�\븨��� ��h�jmm�����-jyJS�x�6Jl��d]Į�*f]2;�:,������c�1&�������~����=1zci1�DN3b�L�YIX��`۠��sPv\Nψ��7-�\�Qe���|��$�����.��4�n�z��+tƘ0������TQ�E�ڤ{r����q����m;�OY�G
zۉ5g��Z��� ��a��)$�d��՛``�슂��7`ö��&t�&���\$�b	 �4�۾$;������9�� �2%�",F�J��	�`Pp��m�ߛR�-�ŭO)JuOy[����a���1nM�	5"�+S��1�4%�,߾��oЈ�>�������U<�M�|{�7��,��i�[}��y�	���xl�Ǔ�u�f.d}=1�4�5<��Mxy�6m�,��6�ܭYU��힓X�\����T}�8���S{�.���A*Scn2�J�R-�#FՈ�]R(È���qhj+"[޷AAcJD����@�1E�����������u(����F��Ѻ�m,Ez>T��F���G:�'���rѭ��"�St�G�O$h�1R97{�Ob#-^i
Z���%9 �F:M�s*�$�#ܓt�I�lA�!#
Q��=�hj��GB]�Ǒ�6&yI��C_[�eU�u���K�#�Sln"�P��,hw���404���E�KJ� P4S*�
M�"�E���ͩ��ߜZ��T�����'.���q�n�&&%
�m�r"��8�8�0��"]��#c"]���U���ѳ
a�2�rah�440�̩ ���Pe&4B*^a�Ql���#㧑A� p`��H�}cE��3�wH�7���c�K�4e|:AI��2��M��lvH[�0I�F�p�,a�N/���}޵������aR�A�H�& ��j��MN�d8���N���n&���5��DǍh��C"�A.A�I��)��Z;R]�����i#Q�QhCP��E��Ã,��"ä0���8߈���Q�z�ͥ�ͥ�2[�c,�E�k��ڴ��ٴ�f^d���Z�_�ˮ3�|�KĒ��Y.I�E��R�h�e-1��-�q���|���2�Zu�E������&-L�L�L�R-)l��Ϳ[�?�ߖ֞g���(���Ζ�%�ͥ���"���i����-�V��%���eirJ[5$�Z8����k�Ks2ZqO7�KK̙����5iiij[]K[9|�Qe�ii��in-�KJKKGϒ�c��z0�?�ð��?�C>(�����/J/H��(��EI$��)h�m-KFRӄ�-�V�Js2���>G�f�ՙo��ZE�k��ڵ��f�ՙ.IIije}�.-�#��/[1^U�Q�G���UxQzP�kF��⏏_�}ujٽ���%��&W�/.������*��+��s{�{�/x�ˬ�8r[�(�#�3��l�L�is�^���3=����z��ߙ�^���6����s��o�Cų.�1�����t������&�S�u����Y.�{�����ߔ�f��ų���u�O:9~�7g�.�鬮Ȟ=]l��g*�S3ee��꛹�ي��Ny��}C��/�ٹ1Sz��*>��L�Ƒ�	�n�����Ҫ������ﻻ������Ҫ�¿�w������߭U�W�
����������߭U�W�
����Dy�y��y��|�����:t�ӁÃ6h�m�i�8�0��{m�T�����_�F���%�tj�v�M�6vp=6����(�v��N�8���1�A�W<N�D��F�]��Y��*82�-��'���,����חк����3��aXX�$��E]TV�$6��4<�MC!�Z!���Da�k��Xt��a�;�n��h�0�(� �͎�vNS�!��:/J4��I�G����|b0�BY�����m�Ab�E���H���
Z7�(��#h�� �
k�p���a�@R�!�c(�g�0��S��qkS�R�SǞGq��
	���P�r8��	!$$��4�8�>"+"�h��O�*��ymM�I�]�ؓ��p�M�O�Ҽ���
��|c�E{VG�9Z�u�����k!�8�h(k�4h� �u��-����h�O��CM|E�
�|� �3̠a��˧x�H�.�rth��(����iQJ|��8�)���!	$n/���"
��QGȺ��&���0w٩>�q�sa�P�CH�΢�)��8|W�����G��&��>g9h�s3�s��r��}�Ƒ�m��~pO�����4N8�J���jL��VۗO��Y�{ʖr>H��F6{W	!$$�� y��z�..�׊���{��������3�t�}�3���{:���8��L����8�$�u�6;�
�︻ʦy��\�g������Aݜ��c�f�\��!:I��K_=���߮e�oz��2e��˼Ww�]��|��+�ؽ�6:�������Ν�]V��4J�Q���E*UFA�>' � bc-[8�+�����}�։6O$;H8#�������*�m�lg���"#�Y�(�P81��ch�D�3�DCdE���(a�8hm�'�ʒS�C"]g{h��Du<|$���R�H�S.��e��0acS:6�t�t�Xp<���>8��m��Q�e��J�B=�ˆHfH�������])���R/�6���٥���Mщ�;MٸbF!D4u�������ַ��:��<���OC��  oICR!όi��d�g��#"#(dDhf}���4a�q]����	��@�Y�*
�=�=�%>3333�ea�2f�%��5���a�i��y�:��0��J��T���,��E`�f7J�"!�援iZC1������T��]#��i|���J��wm�P�,���9J"���5�:D`�`X�D4m��6�&������GlE�s���[��b5��j��"1""���Y<Q�y���V��jS�x�����bV@V�6�3�Zm��m�4-^�n9#!ت�-��Hc]CF�ImVdڈ�H�hh��H43k�|��Z4����j�9h�(e���ݞT��ȕ�����z��U�YY�V\5����H4{Z^G��G�#[9�+A�u�ҋGl4u�u�r�H���4ae�,^8�������	9�8N`܍)����:xi��2˵zD�ڽ>��3O�fhc����K�EL0e��K��u�ۏ>�����{mc2ˌ�֝in<���ZԵ)�<y�u�c?g�
�\�@�ơ���$ҕ���HI	" �|D��,r�FDb�8F�O��fc�
+s�t� ��o�|��9�?+no�ͪ��Ss#��,������h����"ZC3cX�4EGv7H�./3������cC<5��a�qDoF�ªQDb�!q�ؕ���'�Tϥo�˙W��x=���W��AT��,�:�F"�8�fU��.!�09v���4�!Vqt�K�<����W:Tm���C�E�4��\[�ZԵ��<y�u��Y1���(�ne�h2�ӻ"���U��$���"�˯s~�~��r�樬�2桭���}�L�Vo���]��r�I���s�55�_o9�p���s�r1��mE\^V����YU�7~I�e��5��V�3U�n�<<]�ŵ�i7�鎽��[��\i_9=~���{>͛��$�-�fe�V^
<�#�h�qQi��E�K�Yke�`lc@Ԉ��ꢩ���csd0������(�jim�C8DF�շ�b�j֗���Z:p�]�"�S:��is����#���:���|��Ip�64R�h��z `�cEA�7�W��H���G�0=���o;6S�R�h�".&{�0��>��><˸Z��rS�I[qmw�G�"&�ѱ��!�|�p���ќ祱[�8}��L�q�\q�Zu���V��kS�x�����������\:J�
ʡ�%EA|u��m�ޖ̘Z������D�I��M���'H�È���F�wtK�+�o��]QV誩m���qF�(R��6�B��*]6�����"(�p��hg �R;�[hҝ���CU�f�DRl�q����f�ˠ��S�֙����,�<�˼�.6d&�-����EF��E�8��]���5�ޛ�4������
 A��(T��49��C2�@�.�Z�6Ls�g̆ϟ#�o6�R�q��:��KZ�SǞG^�d���朘k���,P!.��i��i��о�ln��\G|��Ov`��h��k��Y~�d�#���-��Ј��"/yQ`�T�F���X�MQ��
�L}��;�1Y�X�e��4�����}�Q�n�Lr3"��4��*Z(o�[zp�)mK���c�DO��
������}��C�#vAϾ��lh9���ܼ���ld�U�8�v:����t�G�fS�7��B�Ix��Q����R8ۭ���>q��:��KZ�t�╠߽�,��[�'���L�J�e*2���HI	" ��Ph�Ͷ����h �"�,�������炜�w����d-u|ޚK͟�b��u1�l����?a�����E�)2#�yq[-x���c-F!���z,4�p#��l�
�wn�L���ѳf��G��*���{�GUg=��(mE�ZوсiTy�h�hѫ�#m�0�c6ky&��v��tj���i7c��a��>!g�X?��0vz6Y	�Ų���S6ե��ͯ3��lĴ�Y��-�q�KKu�IiKek̖�8�ɞIfx��IdY1d^$�H��-"ZGYŢ�ri���+��q�L�%�ӈ�[��['����)H�3�-���JE�-�"�Ih��jf��^g���-�m���f��ͧ��ii�����Y�Z-6���y�E���#�iĴvKg�8͹�-8�O6�?%��C�|;>'�4|O������x�L��̙�ٴ_$ͭ�왴�������Ru-8�?&�Ѵ�Ԗ��-6��:�4���Q�-��-"*I��KF��/�|2���6|E��/��]�8W�y�/2y6�bZ[+Զm�6����%�-��2-�m'd�$�x��IdZDY�"�&,�H��g����2����w��|�����̿���\��9N���z;-���\Ͼ���ӣͳ=�{[=;!����=��4=���˛�.�=$��1���g{7�oi�^��^ƻ���{k���g�s��S�b6����Jgr&/q���9��Ȏ��
�s��Ȫ��f��em�SFA�t���=o���[�����6������{�{�������U�Y�ۏ)k��c���s��o7{���ݽ[�6��7�vg�z��H,�5 iإ����T��"���d�٫OmN*��coy�=ƿ���w�~R�j��������wwwg~�J���VV�z�����ݝ��*���Y[��������ߩU�W�����ް����m��y��[�ZԷ���ĸ����0|�q��c�In����U2(ԵW!ȓ4 W8�X�@��U
	�F�ҍ�W�R��R�[NT�V4)��v@�bR�]�ED55�Zu�U��i�#��ƅl+���m�MǭV �u;������)mV6��n���۶�#�rZ�oB�n��j��#�6܎}U�\�\DQ��jd� ��*���X��!�W�� ���N���i�J*�R�;y`�#�J�R5J��ҎH7A	-��h8�TPv�����PsR���V���E���`ݔr��F
W-,��hH���Q�mtn�厪�a�Ubv��&��nEI�hR�	�ڊJ�VE5lNT16�R�GK`c��Tݮ�WX�n��$���RM�"�]��F;#4�Z�U1���Ym�Z��R4X�:Z��k��vJ��� l��!$58��!c����P�"�+�I��
���+�V�DTA(�-r7cQ��$t�Bl�S��i��i��о����d�r��ϻͿ����;��_:�����9�qe.y��2�m���7��c��&��+.�K�י�_bys�;���<�������Vȭ��m.�y����y���s�sP$`qɉ���R�����|^�7��7�!��Q�k��aR���sPҩY�\FL �sf�sz���HI�4p>�-�4x�,F���N��!JѲ͔f#�7F�C�l��-��k4khY���ː��>��)�`d��b��|��D0�c(f#TyQa����R�.�o�t����!�9�������l�|l(g�����hߠ��e�{Ky��\��r���u�>��y�8y"-���ZBT���3[1aG����v���:�ᖑ��m�����V�ֵ-kuӮ����g{
�iH���M��pSx�4��'��I	!$D�Da�O�΁�ц
���x3H:��5��k}�p��yN��6�̠�E�Q|�:���ZE"�37��6Yh��G���}�쐷99=|�9}x��K�^K��O���Kww3hV�۩��GDN�Yh���l�(�;�:g�������0��H�:�4"(��su�q�%Ą��k�!�-��|ۍ���έխjZ��a�c4\z�$=!ɚ7��5���z���!$$��gWJ㑒E��d�fʢVѠ��>�b*цѨ�{zK�.�m�y4Xѣ�8a�Ʉ�m�䳨�6��!��W>x[r��D�����nH�enI���j^���l$l�`D`;wU�m|,1�1bሴp��
�X��c���[�c$�����m�v�K��U��#�
��k@�0V��p�4qX��w�PΖagŝy�~ukZ�����Q��u�E|4 Ŗt��ۍ$kx����M��$��:���+>�nlm��Z���1o#H�W��I ���KH�l�G�h�3AC>H����o��b�t�D{�MlX�v\��b�4��>��'=�mױX|u~���vIw����4����c����Bv��k�Ob���6��^��7m�\6ѵ,-x�����>4�6ڛq��|�_�Z֥�n�u�q��Q�M�����#u��A�.�B�i��*|y��m�ޓB{\��ُ�q��*�o�둛ܛ�j]���<Lv�ٚȍ���Ms�X�r��z^����9N�������+Kx93�\�h���������̃ʻ]&�3�[ݪ�g;���������f��X�ۓ��'*��n�"�7+�o�^C1p�_%>oA��8�f,��]��*��4�lh"<R#�|���{Ͷ6�g}��4t�j�,:舫כ�Lɹ>lr�Xe�^o��E#��V^��[G�~q_,[C,��Q�a�0�l+{��vS2��B�W#�+Kg���6*��iq�dY9�8#e�v ���1�!�i����Ð�^>�çm��~mOϖ��ZԵ��N�����jTN�4��!R4��\$���"���~�,G(�1���'�$�#�-�i@�Ψ�ϑE}�E#�a���74�������6��x�8R�R��:h�+ï9r~��^�ȉ1���7���O��F���=��%�d$��C? R|�����+.��>��|�E��Zl>c��`�!R-5�t�Ґ43\���Z1�0����G[[o6�?:��ֵ-kuӮ���}ֳF�޷��H�	�b��i��i��лώ0�*ab�f8z������w���6�63�4b�E�͢���,�p��?o�B�c=XO�Q#k���G�#�^:b61��*�r5���kyR�kWXji�sG���m��XPhe4�Y�F64i3KQx�!٢�ش���s�����G�HJ�l��Z�-���{:a����H<�Q~c64��hF���1qx�Ph�m�ͭ����~ukZ��:���hp�j���* S̨�����DA�EDs�L]
F���]9E���}���^7;P��I/	��&���t�5���F�2�������m��{�0Ƣ=���f# A���u{�ym1�~�QU	!J}\��o�m5��t�t��=I&��#M�V�xΰ�c�Dxy�6��ͽ��6DZ���W��r7	�g^7�G"�i����ukZ��:��Q�}�{5-5[5��}�z��:�E�����i�KC�����M���hO�ow�y|�7^��M�r��x��|��ō�~�����|����L>TM�a�l�v�|���8G���^XA]���ْ���:\;�s�������w9��a���hcY�)����(�I�����i��@�unw';�z�{��~�b�U���=���7�_�-s�=���pwv�gQf�-??'Ǌx����BDw���0�q��n��wŉ������R7�6w��[��Q4��3�{�nn�v�l����jkkeZ9��9���R(�<��>{����C��u���3�����J1�N��٤Z��P����)�5OV�*��#v��D[1t��(gW���7�{HԈ���)>i�o�>[o�[�κ��KZ�6lf�h�)�l�-���Ț�m�0lEfg7p�BH�1��>�	`@c>�xqf�"�F�{�e��ۚ�߲yg9���
�>у:@��7�ܟ/���D{ț�\PS�Hn�WU���F��ህZ�0�-@����}�yr��̆dO
�y��0m�����^vNX7"ꦶ�Mu�t�rs�ɂh��<�i,�<�#T&�
gi��qY�u�XY�V�>0�e�Ĳ�� ��B"&��P�$�bh��	�"&����d� � ��$�BX�%��0LD���8N��8N8N4�,�4�I$D�(HDE���&�	�x�J D�DK4D4�H,O��i�p�'�ĖP�$�T�(�����Ylqh�Z�-l�R�R<�:��yky�����%���'��&xOH� � �~	?����̶WS��_w�y���	�xM�[ᆙ/����sr�9읛a�z��mLu�ʯI;�������2��u����o���#,;qE��*�[�c��8g\۵��jzٛ]�ݮ�>&7��8�����3��{F�B�&m՜���r�^�����{.��un_��9�lS������C�d_�r\��o�������Mu���<��=֭�Z��Q��?^M���L��?�{��}�mI���}��dO��y��of��~�U�+w���wwwvw�Ԫ�U�Zn����������UWʶ�M�������ݿ�J��V�i��ۼ���^y��6��un���K<tٳc6CG��w$$���"����l1������J��2!|�e�~,\��օє�FZ>>4�T����Z�D���'��R6u0����9n�'aEI3-:�UU��Š=�hP�b��O��f��8�l�2��lv%�6�!�F�bc8�/#H�9��]�N-�he�7Q�h����4q0�=��e.,E|{ç�ee�4��ֵ:�]Z֥�N��:ˎ�r��7��n1��13B=I�^�Zm��m�с��z�NLE"��~;�Fq�jC�ŔkS|^���7�N\�I�㹎Ƣ��Y�n:<NLZ^8��c�Щ�mq<�`�(g�q�^ØV�s��a�1�O��>6_�f�EaC=�|�FȃC!���N���n���Xsd⯇��țC��WY����֛�G��5k�h�/
����ɘD�h��{]�Dj2�9�h�������ͭoο:�ֵ-ju�Q�\Y~�m�����Aף.�F�,n�b>�m��m�4.��f>��d~��| .߱���ق����n����d��_]N�v�2�C�����$�G����/g�g��
y{�{w�G`|�V!<P�62��L��3��d��L{�S�J��n��T{��g:gw�l���m�{޵���ɭ����7�a`�Z8�R)���ȧ��#b��A�K��O�l���:��3@�|�(������yٸ��Dp���yY�Ue'|���q������3c-}��G���sKe{���F�W�"�jB�x�gJ^���{��^��[�Zz��Y�ffX��Y���G��W2�3�^6��4;��^�M�G�[�P@��X,83d-���mjS�κ��KZ�u�u���<��a#��ۤ*��C��$���"�"�.4u��ʶ	I���ރw�#~u�a��!�F͓̰e:ω$p��|���v!��u��6*����o{Fܐ��Q��R׾m�x�Y�yח����y����U��u��6L��n�n�*�0P�k���#�Pl��|Jmr�k�!�,���ux�㦕�{�Ű��:q���h���#rG������:Q�ŝyn��V��kS�����X�S'z)R��,�A4���m�"!~�N�_�h'b�r''�a����I;>eܦ�)���e����U���Φ�H�xа폳�*8��~���uZ��U�o5z��b��ϐ͔������,��1X���N󝦰�ڴB-T`2��v:�leT+�ѣF��g�Z�e,08Éi���/N�6�<��4�~R�~qխjZ�뮣�����CzH�NW^�$$�����j6��-�((�X�Y�r߇<�uW���]�mM�2\*�
��U��H�E��Z���;q�#c��fo]�	�x�6�U�(���n�:�Q^��5���BScF��kmÌ�ӽi�w:�O4k[xih �GV�����e�ٲ��,꟝~qխjZ�뮣�����Zj�y��j�W>t*}�I�����s[d\޵�rBHIn�\�kW��3��N�_i�mI�}���;����+g�s�W��ǯ�v�zs/�/�u������[��x�6.{+v��2K]��e*���ɽP��p��6�3ޕg9�=}�9W�Y��Nm��ڮJuform�,��h�hރ
���j�t��/��iK������4����A���'J�O#�ƪp>]P8�o:M����>��J�*�T���#���OX@�Z"8�����TR�y�щ��v.�0�=HJC�2ˬ��ck�mT]:�
:�(��d��3GFR��6ی�����Q�_�Ӯ6���_�ukZ��:��.+�cQ��������/�BHI��KJ����a��ÙJF�xz[n�Y{�'�|��hk>37Ϥ��*����C�'���"4��׼+�w��X~Ɩ"Ϊ0�˅��H�Џ.҆,
1~?��)��~�6��y����ᷦc���n���r^׵����qp�Tl��7�٨|Qhh�\l��1f��#��Ti�KB���F�ؙ���ca��jE2��~q�V�_�ukZ��:��.Ę���a��3��$���"�R��6P4�����mA�u�t�;�L��af!�-�Z�nuy`[Z�i���|x�p�����!�I�w2�0�و��g���5,G�Eٴf���{A,\"�È�Xl_wc��!�N�'|�qX�ʰ���m��lh�-�6�����4xg&��ukbfQ�]|Ӯ6��:�Z֥�N������~G��H 7����j�$$���V�8x�>��#gA�R�v�lI�d��}#z-#�r��j��>��YV=kD:�3����?v2G$roͶ�l��;���#���>P�|��Fw����ª>\XPA�2Ǳ3ȣGƁ
1,٭�QW����:̼�Ķ�������f9���7��zI$���#E[�F�#��fi��ԇd0��af�H��Yg�DJ��D DKN4��0L(��� � �p�QBX�%��0LD�8�D���4M�DN4M<H�$	b��&� �%�"x���%	�F	��(����DM4�
 DK��8L�'�,�(II���QEy�_���kl���kt믝qũ�:ʊZ�Z��ַ���)�q>S/�� � �~(�{}��:*ۮ|&|k*�s�h��	��z�~����Q�g��̍�yqYų��"g��E���Q��m6��3�^�	ͷ��=�,�����N�{�o;Xqm��me�q���{�&*����}Oެ�w����P��q��I��rCfEUغ��>���Ҡ�a�}o���c~�N���ٝ�z��r�Ƕ63zb3o2�as}���:{ܳӛ�Ͻ%��QI����|j��hɲ^�Y�+�fcsR��әT�E5u��������=v�;i����ʪ�V�i�����������UU�iV��������~�UqZU����������ߡU\V�[����a��^y��q���[�Z����=�2Pn��;����[� r�B��J�;Im��I�!\�Uk�B��H��A�,t!%����uM�+B�$��2Z܌�p+F��9������ӭX�����F�V@���X臤E�cP#�BU��-ӭER���4;Z&���l�v�c��(ʌ�Q�'���k%�V(V�$�OE`M��*�P(H��hz��h�Glc��ת�e�C �E��((��[-,j
���Ѻ
ʡkԢ�����R�R�	����J�Uu��WVGmvUl�ɪ���,#lV�VHARʫ�.,ő�k��X��Z��e�І+"q0�CSVE-�2�!D1�!%+�*Ԓi��(�nF꨺N��!EPjI�m��i�T46�V��&��a#t�" �v8���$ �WU���[jt����5[jjDY(�B+d#�"����ЭҎ&Gmq�eU�*����4X�ن]Q�Tʬ&���QZ��%D�曕[ER�l�1[�F�P"MWr\.��)�NBHI	"!y�v�!�[�`��[^��ڛ��9�js�oe��x�跛�;==���Oj�6��N��L���o[[�,̽7���9��QV�1`���+b�U��w��Ƅ�V��<��z-�w˪�۱��!2�<�/V#��{^�pX@�is���-0�Z��"E��j/5�~��,"����=�]����31ݎ]d<��C8*ƋGQ��ӣ8��CM?c8u]\O��|P�d���0��Gϓ���Swx����{ۭi�r\*���{����#��<�2��ui��M�Pk�
(e��i����_��:��kS�:���Ү��l�.9%�>�i��Jc7pjS/D-��x={2BHI"�-�������"׍`���CG!�ҡ��e�F[d�:zF���L7M>��D�v�>�;����ٟ|��tr}h�Z���a�5�)�����L�m���P��f�&��UJ�m�}~@����H�_4>��ِ��
��$D|E����a�uw��-�Z8ʝi����_��Z��:p�͐ѼH��*8	�E�nBHI�[�n29�1l�-��9#�4��s���,�]9���ŜDF�h�9��ϝo���\������{�Y|�r��G�����RCH�>>;h�#o�����<Sp}DT�kۡ��Xe����}���X�Mh���o]鏂h��f�G؎᳌m�9O��Gmm:ҝZ�~[�-jZ��Σ���7�����ynlyP���-��Ty�̄��DB���B����Dp!�Y����f���Ĭ����jEIV؛��=ߴ��Jj��N��5�9!�y�� �1�F����q��To�MGUE#����K�k�f��/\5��p0ę߇���,65�!�z9�m��Z�F!2�%`ϒ����c4�F��1hz1x�兔��� ͐�4�^[��yŭKZ�y�u��j1?�i�0�]ݙ7n4I5�MܵJ�v���m�ޓV�o����X��7*3Y�ѯ�7~�k"�s3"&z�!���{�_WL�T�[�34��+�W����g3w����ٓ9��«z{�g�z%��ɵ��R{��͹�� v���J^�,G{֯f��\Q5���Xڻi�0��\�z�u*�Z�:ѳ�gy�cŭ�p����N2�i!��t�4�4x�a�͢�������:�\c��I���H�a�k�͑@��G�[7_h�m���L[����8��3��iKFzwYmݽkSU,�&�)�k}�\�U��͚��2�֔��[��yn�KZ�8pf�hm�M2���{b�df�2��Upz�SIU�T$���"&��-Z��`2%����U�p�ip��5*�)k��ϵo�GZ�ķ�8�Б����%_�bo��E�p�#d:��.��CZ^Gt�lfՆ�գ~�����r���`�H�Q��d��h�8�;D��|C]h��j�����M�"�ȵ�q��UBt:l�Yk�6�C�8�^�e��H�
׾�A��h�������Z��:���./���s�Q�L-�9	!$$��q��VF��Tꪑ��#�CGLDa�H���|k����5�4@g��ô�$��k@?��}�}��r^W�s��Z+�N-&���:<LM����=��*���GC��ș��hi���z�Z/r8F9#>Q�ae&�\�$���ՄB浺u^ZE+�ƍ)eo4�N�<�V���Ե�מGYq��fbBg)�r�j��NkP�BH�mb>�垒b͜$(��ǯ�F�8�����P�fE�{�G\�mh�{��
���fa��1���"8���C�_[��()w���N�Q�h�5s����[i�iB4Eť��;pn�<�7�I��>u�z�x-@��a����'���J�l��O4�~u�o-ũkS�<����/�;��֊@�J�af9Mj���:��8�
�4���mg�BHI	"!�{�>w��C��[z+ܾ^����������ٷC1\9�|w9=9�'�"�s0��Ovw��}rv�l�����F�w���Ҵ�����U�:�4�jq����wx�oyD�r��fO�b;Hüm�t��������;��^�\�̘�x��gE���i:�q������҇�ї��ѵ�ADQ2��>{F�˝�C��'��o㑍�&�
c����]�Xlx��1�Ͼcm���;���dR��V�J���-k�:F�i@�
m���K��&��ń5l�Y�����n�*��f��Z�F-���C@x`�i��G{��ܕ)�?�#H����SN����ykuKY�g��2�rH�HS)�ats{���DCH��ym��a�����oKF�ު������]F�|�p��F�B���E�6�&ݡ:�hH���SG��/�)�s(22#^J��UF��-C:�F_����m��=#�]~��Y���d���/Y.���ѷ�6�c֑�"�>°yi1~h���$fL啚_�-1ޙ̿�mit�iw�#+�}��?9�c�Q�/��K|�ո�M���h�"%����i"�"%���'��xO	�,�A�A<$�!LBP�"xD�1��4N���<'	�p��Ɖ�� DK<%	B&� �$�BxLD�D�0Kı,��,��""=�H�$�'��0D�8L�(J0�$J(�J(�LQH����-n�[�M<i���4�H�D�-k[ϖ�o�2��(��'���>����=��艝���ں�&3���3���K�������n���s._sl�M�?5}����a/Z��Ǽ���o}k�c�g{8�:���ܾ��"��o���nX�T�TN������_no�)�81����8���vd�=���}�ݑ�9a�N�_6C0Ûo;3p�9���g��^����y���Qc�Q���z��*��xZ���fq��g{��~�Ъ�+J�����wwww��
�⴪�����wwww~�Ъ��*��ݿ�����ߑUWVU[��q�y�I�i�[�[�[�Z����4܋�!$$����p���"͞M��qU>�1�h����Ӂ�tD4��&�dG�ȏ���6�ŞF�C:�徍ʕ�]c��'ywd�#�o�#�t5�U��_#H֖�����yE10h����8D|Q�ut>,���U�9�ʪ�g�{&/�]�i��^G����N4��~u�o-n�kS�<�3����7֔8&�j7d���]n	�+�{�֞a��f'���%��3ѽV�9\SO]�W����ho��tG썦fDeD�{WK�� ��U~�s` ���){e�R
j�5�rFj6ͱ9o�Ѝ#���<��h)n��nB�:��IC�=���5�q{�F��h�5�>���'��]�2���x�^�3	�yUɣN>�Gn���|�I�i�O-�張���N���յ5⨭��3-UA@���ݤ@Ȩ���6�m6��}���^*a����f������˴zȳ'���r����\���*������x�N�b�[;���w��yM�S{|7����q3e�]�eƻ��AQ>�0���O/2���[Y��f`����r��˾q{.�0�os|�r���uǑ�=�3i��N�iz�tb�8�����A�d9�G���>o\>ǵl�'�&�M�9)���'_z�F68�D|��ci� ������wrI��,u�K�F�v��k��>�}�Ԯpl��[Aa��üm���ɵ\ C�c.|��Y*�*�[F�F���	��l,0�>g�y���<�V���T��ל�=��z����Lʻ ٕ;����1�ɖ�Ӑ�BH�Pw��>m�-YћF�����/��7!q�y��7��R4�á�6��Ȋ��t\@_�Ni�ҥK��A�a��fi�G��W�F�|��h�4<�cV�!�}���#a�mY�m�#�UX�GA����D<�zL8S�?a��Z���Q�jN4�����V�4t����i�H�LWtJ9��I	!$F2�h��#J�Q\{��d�td.�s.��SM�{�["���>I���mb<Y�DѠ�����ka�RO���l��S`�\����_�[of���pi�q.W�l�2�)�R>"8��o��vt����i>�܄>��e2�"�>�y|E�kh�Z9A�O7���x���_���▵:���<���^�%QT�[���Dg��aJ��G�1�K��7H�
�!/a��i_����]�yI$jjjfPՄ>�����Xqq)���֊��3�:q���>ƽø��֤n�j
[2|��[�~�>��RH��l�Ʊ)�&�ώ��WM��F��4��:�q���k�X|㖱yG�W�>#�o����F��QC,�oe)����_���▵:���<���X�қ�����1�m���4��/hEAy)"�q��m�ޗ����9
��<t�����qs<x�۬����1�{2��Ǐz�t"	$��w���K�Z���4Ut�ۜ[�__N޼���;!$��F\�ɽ����#��F[�����q�y5�kOH�x�/�v{f�{Y�����q%+sy5]�ٜ� �����4�]�����/��U���$��+w�F�m`B���Iԍ���<f�ކ=�c|F�h�`3ӣg{8:�u��E:|DX��&�F��4�m3i��UQ�S_fU�R�/2�~6�<����������${Yŵ�XB��>��)�T������Z���p�n�}Q�BU7(���HI	"<R<�8{Aͻa�N�G�U����$I&y�+���g�H��Q�5�Q��>]Y������/�4U��5�r8��C��Cx�l8H�il��t6�1ȅUC���ߪ�zz̪w��D�f�6��و���T�B��ȝ*O��ٓ�Юj�Q�&?S16���/�-�!C(�o�)J[�~[�Z�Z���#��N=�ǥ�F:k�U��Vw���=X� �����$$���"�˪�����"1Dqk��ц�#+F][����1z£tɵW*�ZS��4QK����W��u�<ٳ3o3.��J{�D6��}������#��Z4w�$�0)�Ͼ�B|w��p=��\��e������cy������z-���x[��>g�ƞmז▷��8��מG��j���)�fF�(�T\����Dl���k��mJ�q���6��/������{cM|�_y����1��,՘B�N�Yo4g��*G)GC����4��>*F#>8X|hm�ي*'b�	>,�A�[
|��P��"��EU*Na�4y�1Xoʹױ6}�kdTh�o�[6�Z>]���&N�˪k�m�N�믔�|�DO��& �"X���p�����(�>A��%�"QB%�D��4LN4N�0�$ND��O"$��""u��&� �@�B"x�!�D�,K�b(�(�D��G���& �"X�&�'	�xK�8�(�D�$�DA(�LQH�R�����mou�a��p�H�$�b"&��R���Ÿ�+eYe�P�p�1�������s���L�}�]�s\��������Y�[�t{՚�����5A^[����$�{y#��9�/D����$��?��-�_zw~h��o�ǚ���o(����]q�j���w�������*i����y���0Ӟ�2��l����d_�8�9~���/��K���u=���.���٬�|{SO�y=���s�ٜΙ+�D�m�l�Gm���پ��cǡye��ٍ�8���,�v]�^I<���vGWG�_M���C�O��9��ެ�+;��=�ۘ�O���gb�̪�����{p��C[c�1�~�oEC�MNo1S6��d)�d���lo	�q���z�z���'.�(�O��s�������������������ߑUWVU[�����߿"�����wv��������U^aU����q�qGqg~1K[�Z�Z���#�4�T�Ǿ�3�����z�":�	idFR� ��W��4��H��EcN2�J�T���lR�F��V�j���U�UM��$A+��M6��P�-R�
��[*��B�H���G[A4��D�l�W��,��t4h��(�U�C�;�Ui((���!���J�
�i�P�u�X�F��T�
)%u�A�('*$n�D��һe�N�TQ8�TEZ��v�MMQ=:����b�� *���E"#d��$���h���ǥkv�K]l���2��#CNGZ�6����#�mA�JhvhLdz 	ʜN!�JU�c��Ɓ�讻.��YrV�T�]h���a��P��zQ8��TTm7�,m�cN�Uv���]j��*풵U���U8�\m�:J*�[v(�h���M�"a-z�є��5H����$�\m��:J4أ�XESN���eE�J�4��I�E4�ڊ�����JކЊ��V�D�TnZ�%dv��6���N���J�����q��M��ү{����X�{�>s|������qe��k�œko�����$��������}��5��:��Q�y�v]��&B���}�Gk�Y�U�H���V3�;w��}�E��Nw�|Ym���wa9Ï�V�.����[�F��M+�׵u� ������o�<�V�]|��K"-��}]h�4=�n����Z�p�}n}3�L�\˹̸fY7�x��*�\��ӎ�i9��`;<�M��χ�h�Va���8�6Q��"4݈-�K��_0+����H8Y�J�a�6�.��k���2�1�h��:aG �6A�p�e,��S��Z��֧^yq�5��a6+�%�'-��rԸ�c�<q�Rk
*:�ӂSv7�8�Z։*��SF����4q��UBA�����k��|M��G��"��˪��!�^=7$&�Xb�p�|�y�����6A�/��Q��V�Y�aT���"i����֙��uh4f�y��$�0��&9��ӎ��g�s�������m?4�n������>Z���#�4�Չ�h�970oj�|7�3�ͬ󸢊M�|�&28�#H�e���6�)XQ���ke�1qip�Dx�M��k��p_-��E%v��˺�0c�V�xC1[�wqUE0q�t�}E&q�q�r�mɠ/B)a�+Dx*�{)h8y��{M���h�5��}�Ȃ����T�A(�0��4��"����֥��:���&=��v}����7��m��q>r���� @�EjҖۨۏ�����"��/(�hz���������	�cCO1�C26|���⺍�l�n���3�gƎ�_Q��>+V�^=y�-�iY�c�UB6�R��H�A�i��m�����"$���L8��ْ��k�E�q��Pcl4@=��1�:�N��ַ�����<h��g᲋��jeJ��$d#����lC[�WYvg�@���mῲ��8e�~�sw=dX���^ә����&�������'�6`�^�y�yk�%�TO���v�҈�N�i�u�����'�o^|&=�.��w�-�ۼ�],�L�5=���[�I�OW����ٿ�F?{��o�w�i��F��#T�c������ �=�nţx���Ѵ����oH�Ú�����|/�ߥ�T��*uTϺ1�����0�:��G�ܔ|ìh�E>�؋9\�q�Hۙ���η�")U��|h؆�� �s���a�ܜW��;	��7Y�7��L�y��#������1���jg9��7�?:i�um)��������֥��:���=}��E̔Ǖ�oj�$�[�M����ccch�Q��T�KG�A��F5��||xx��6l#��W�Ӓ�FJ�P��iN}z_��<m��z-i��\Ul�6	�u�GQt�|��8m���|}��<�er���Y#�uk���J�:�]Fβ>�A2%Fi�-���U冖������Y&�H���NXb10іQ��|��Z��ַ��-ũמG�i���������w7�D	1jWF���~�4��Ϊ��J~�t6Xy}��P|�������~4�Yh������~�yޥj�/N��.��WZ�_#J�����e��c~|��n�Pq� u3E�]����BmA�o�ه䀞n�I)�um�6qM��Gi�����iX�0�5��~�>m)�������ַ��-ũמG�iﯰ�-U�R-��z�����y�,�Cm�+e�*Gh8���5�9"ר����N�l��Z,��JG�p��í-�9"�T:G��Ma��?1��"&+O=������^�s:�(Q�1�V?,ic�m5���`
���P��壟)E}"A1�:�&d�o|�|Ӎ)������֥��:����A����*&��sOHp��@��-��ݝ��&��;\N�=~��ӳ����yp�g�nEf�پos����U�V�Vc��Ou��t�S�������cy�'���#��g���l�)T�޽���y�3���Wy������fa���@s��n�g^���eE�te���l�m�E�3��ki|b���8Bua��U�2�~6M�MP�����YN<�K|c��,vfQ}P�4�,�(p,��V�ڭ�X0�4Yg�)D=��8)8�#�0�9U(�4꩐�-l��.,E�(4�-�����6��4Q�m�ŭo-j[�S�<�:�v�2�"�3;�(��������� ���^]׺��J��շ�R�@v�S�����V/�1=�)-MgRބ�V��=܋D0xp���zI���:�#�b��"/�6�1��W�0���N�+%7rɍb;��p4���rl�ӊ�w��x	_-��ښ�kf"�H����4`7�iuo�����l��ͼ���q�G�CH<""p�H�"H��4D����xOH� � ���H�%�%�BP�4Mb4�D�8N��N���O"$��""%�!�'�(DO	'	"&	�X�%��@�'	$�����D�D}�=�&��<%�dp�I"H�Q" �h'�"H"X�B`�'��qƜq��p�H�"H��4D�)�:�O�����K,��,�H?��#;���frk�>�����x2��k#��-i�����h����{�^�r���38\��[�\�gx��X7�fOq�(��n�l��;�Ǐ�ua��f�D�3��9�y���o��y8��5�;�{���%ϧU`5�(�ⷯU��#���Yw��K�Un��[{헒\O6�׳q�3pV^Ǟ���������}'��E��Ss��J���ܾ��{�*��«wwo��������
��ݿ�;�����ª��*�wv�:;�����ª���wwo��8��i�m��Է��-����#ˊ)O1�Bk��+��_IlaX�z#����o[rN�����r�U���Q�gQ;�>F������E�!�qM�S~��"nKR��b�j�[K~�Н�o/	�:ON��i8Lx��_$O]6}�ܶ�c�c��Qh�Ώ�E��4s���iq��G4�Km�Kq�KykR�-N�tGG&���/-iȲ�2|ꪠ��_WFѵ����66���5�r�=D�Ύ�$ӥ*s��!$���ibڇ�R��<�H���1��-w��C�����m9K���Ќ��~����e��卺!,h�gǺ�����l�li�ܔ��u���a�c5�c���Xl�Hӭ<�ͺ��~R�ZԷ�S�<�:�$���q�ȖL��'���Wu��m���_� ����yt�F���c��>���{��^7�>�=�:z.;�$��fy���rb`��M��1y2f��ݚ�y˓}�[��cT�{tL	���<��5��o����o�[��I�/������^�mZwo�yN��E=�-ə��(�w�殖�^�뮊y<�&yyF�y@j���Y�x�3���Pmq��F��^��ҋ���&Y3ʏ�o��:��G����a��
ǃ{�$:�fאÔ�&�R���Ce%���Ԫ}��¤�ʫ�M�hƝ���5T[vAǚ^��ď0���9����]�~��u<FQn4�N��������o��N�elE��y��s��&�T�y�RɅgi��bh�4�DZѠ��F��Vum2ҥA��s>ܯ]�8���7���+�|P�L�-�oQE�/T�ehi�Hz-�#ȳ��~kiٌj.����+N��ʳ3�"ɐ�WN�GC=KH�GJ{P�Z�{\9�b;�a��C}?B��M�|�i#Kk/?"�����Ϳ<��T��m-N��<�K��9��'�9%	�keBe3�� .k�����v�:�5h�biԄ ���;�\/�m'GUWD�&��'F��EC,j�>>GG#cf"��.0�{0�;ǟd{�wo��+P��u�����K�#�\F`�aĵ�-='�l�m��<;��q��&�ik�c�;
{k��ԸO�cܧU-�_�pX����B����H�;��a�>:�8���u��n-N�kR�Z����WSZ�>>�K^F<~`c!�cF#88aJ-YJ���-���z��vfz��h��!������ݹp�4�"�&6��\a�|�4�|Q��4�kM�k��3��}��o�ǎ�kWw�Q�K��U���4�ѝF�A�%�s��~�l���4m�D�8%֩lGS`�܀7N
�Σ���64���a3(�F�6x��uJZ���'�G\i���=�s��E}RȘhE�%��(=��  �n-���R�m���\����z��H��9���o��p@9�����P9�������Q��ɼ������p�|��u����nGqs:g7�˒s��;�Lv��Bb�7�y�g^Lz�'gt�{پ�7�����^K�NЧM�C=�Vrs�cq�e�`Ü��֐֒��$}�YT*>[�ߛ�6��p�K���]�ԏ�T�ڦ��j8�&�>6v�'�����"��6:�G��0ѣF/�m��ل]:�E"� �6��=CV\���{���V��f����iԘ���4{�g4�F�Y3/a��?�GZE?��iM���8�ꔵ-����5&��u��d�;,�w���6To:  �������N����)��og��ܻC-���©l������,5��uV~qlln�7��E6���3�E�#
�[j�Z2�����]��}�!�Qeh�����l�&]�0"��m�K�^׆,�a��0�RCe[>�8��]:�����^���N���l��
���u�u֖��o�~q�N�KR�yo:���o=��kX��\�ki�.v7�ѐ����[���ci�E~�UF�=E�!ỏI�vwvFYo���)6�5���i����DY��
qdof�ag^0��:��=��:\ɷ��Ž���z����k`t�H�څH�,����+6���ѵx|#o=m��(���F�Ʌ���f#A�"ѱ�p�qlt�H�֜i�ߖ��zJZ�&��]]B�ڈ�kf�t���ZԗC�e��m�Ȱڰ���pĸ�����WW�0s��*j��nђ[��"�F�qiis�i��n5�aH��6yDlkH�D5��R-yC�݋���;ٲT���7�6Cu���5�q:a�x��mF�4������t�{���'o�����>䡊$������aAP?����������� �l�4]�`a(��*�
�������I�mɧ[��� �<���;0DDLPL!C0��LL3���1�$43L�10L�B��10��0̎�0�L4L3�0��&	�Hf	�a	!�$�b 	 �"  ���Y"�"$�b"Xb"H"&&"&"`������� 
"$�"b"H���5 鈉�� �"$�$��""a�"b"b"H�$��"!f"$�"H"�(f	�&H""H��%��""H��Y�"H��""$�"Yb�"$��"""b""X��""$�������"$�"H�Y"""H�$��"H�b""X��"$���$��"���	!b&%��b"X��"H��"%������"%��"��%��$� ���"�"X�$��b"X�� ��%�"X��"%�"H!L� �"�""%���%��b""X� �!`�"B%��bX�� �� �bX���"$������$��""H�]8AD�DLDI��1LDL1ID�D�D�HA,D�B�DA110!L ����"H$�!d��"$�"H�$��%� ��$�"!e�H��f
 �&"	����	��"ab	�������!`�"�"H�	!`�H���$����&"&"	���S$�� �	"b ��$�"HX ��&"!�!f"	����`��" I�b��H�(	��$�Xd�HBHd�$Y@��`d`eHR�� e`e`2� e`e dH�� `�`B�� �dHB@��`dH
���a:$�b���	�02$!@�00�� �ʐ0�& ��0$���2���#��L!��2�) @�00�*@�2�*0$(@ʄ @�$�@�$ @�$"�0�*!�1@C@C��0,
@�@Ȱ0��@Ȑ2,�(@���
@�02����	Ȱ2�2!"��+ ���2
�B���"�*�! ��@J��) �*�) 2�8DAD�@B�@J$ �A� �	�1#
B�2!�0�0�2�
@�°�0ʐ��0�Ȑ��ʐ�������B�0�020��	��2����2$000$2��� C+
H���� CCC*C
C B�$2�0���C+��20��8�Cɘ82C�C$1����1����DQ@2C��2C3
A����2C�2B�0C0�1C0�2��2�1��3���C$0C$1C,2�),3�C$1��2B�C$1C,1��2����2����2C,2��2��C,1���C���	������������),1X�2����
A��2��A$@�A$�IA$���,�L�@30D�DIA0D�	$A$A$�I �$�LA0D$�D@K@m��`�		 �	 �H � �X	 �	 �&�	 �&`(H&��&�`�`(�`�`�&�`���BB!	�%�"	��&��"	�b	�H	� &�& $�� ��!�H�� ���� `�& ��`H��"`�&�f d�`
`BH`B�&` d�� I��H	 Y d���HkZ�q�H $��H d��� d�d��H&	 Y �	 d�d��$���H `	 d���`f`Y���6�ȶ�L`a���f ��"`f ��`"	��	��&���" 	�`��f�f � " �&��f	�`I�a���$ �|O����w��x����?��P�Q@*�@j!7�=����������u����~��;�$85�������&���?����?��퉋����W�AL?W��v���G���?A?�����k�y��g5�������з�����g���> ���������~��	�x�S�������	@T ���`?��O���o���h������(I���\'������?������
���@��O�������>��4?o���$;7�~<
l0ƙ~i���ɉ��I���
�����������}�A�|����ڢ ?���O���pb}8� �[U��M  ����0J�z0 H�J(L�$Hk���H�����¥E_���4������,�� ��c���#0a `H;0P�`T�"
 @�"A��~�}L=�����/� |��ϼ���>|�x �?��o������?�?k���VT ����������<s��t�8����=���o��C̓9���>��8����;�$���>O��|�����{�߰���}C��@�~腻_����zg����;�9��Ǆ!>#�U@��C�(
���؁+�_�����X�v�n������wN���wXW�u?j#PQ��sꨏ�~��|O�  @1'����7Gpp`���q,L#�	��¦���p���5LVR���%��q��?�< ������_G��x�|�_��P�~�q���K�� ~��@�?���.<�>�Gп���HhW�~���_1������?g��x7��H�a���o�������P >G�g⃟�'��+��@A�>������3���OO�? ���zK~�H}<��P���DD~;�����F�������]$���~ t�ǯD�G	��vu�;����@�҇��X�NI�/�����: ��`�#�?���}I�=t��A��l��������/ ?��$	"����������C���n;���r���~Hl�����|^��!��c�q����g̏�34�0���������)�(�l�