BZh91AY&SY֨k���߀`q����� ����b!�    `                                      1�QT��  �@       T  �       �          �� 3s� ) �I�U$��U H(P����DHJ�E
��D�H�((!AAU)R��E�
�@j�R��D�RU�*s��n
��J�����nER��	�Uw[�(��"����L��C����A�1�  � ��� TE{��|�_6��g@�yUsХP��y�E�W-AO=�=��AV�R�:�8�����ٽ� x   � �2DUAJ*�
R�J*%/ C� ݀rv r��9*E�!ϰ�@1 ��` zw(` d9 �{D�    �@���� �}�ϔ�� ��z w�y������ s�I� ���ް bJ����z� �P��P �_
��RPIT3a)'�!�� �`y��`�c�` y�y*�x��c�����x�� ��RI��q��{< 4  �J�p>@C  zX d9 n��@�� 8�*p��@�@� �2 >�4
  �*AE�HP��H�$ � $<�7`:��wX u�)*X��� ����� 9¤\:P�����  � /��@��������K���@d� �s� �8� H����Tw`� i@  >�
PP�P��@!TI*��& �� hn`�p$ -���t$��� ��A��9 r� @QA�>� ������qR��: w`r� �7`�r*���� d�d �� ��     �@
R�&��`L��h���~	����h�  42   ��eT�j�!�!� �a� y)����&��40�!�&RJ�2�h��i��M4h D����FѤm*7�='����6�'�S��C���~��m��o��T�7K^����m��^�9���*�����Ȋ(��Q@T�Q_� E��ȸ$?��������̟����~}?�
�����$�OX E�_�(6^�@PPW_����� ���*�Y� ���b�]�����'��A?{D���TL �H�T#�D� A��D� T�D�P�z�z��D�N�N�S�@���:����:�M0�P���X�u�b'X��q��db�� q�b	�
u��bX�=b%0C��:����,�T�z��@� 0�:���������:�z�� �:�z�z�r�z�z��,�:�#�W�W��W�W�D��������W���:���F0^�^�^�^�^����l�^�[1^�^�^�^�^�^��:�z�z�z�p�z�z�z�z�z�z�,G� ��� 0�z��� !LPC�C�,@z�D:�P:�D:�P0�D:�:�:�P:�:�P���A���T��A�Ql����D��D��T���i�=b��`�`�b�b�b�``�`�`(�*���u� u��u� u��u�(u��u��u��q���f���|ݾ�+�ڛ��hD��K&����S���v�S��e�o	�����0�o��ގ;�wb�;ۛ���ǏgXnH�dY��]���͝q�F*ѯVRF/��8��p��Y4�]hc^隬�2����:�\�&'R�+�P����L�a1v�R�
�b[-\�n����E�� jq��`�k�ܸ�c�:<O��њ]�K���[�jȻ�ĕ�i�?�sw<��Ďsz�x�}١�чⳕ͙MW��j��D^�d�=�8�{y�d�!�6�Ѵ�I :,X�M�<@<͘�9o.�8u��+�F�Ǯ:����C�sX�C�%���4��<Tr|�����6�4`�l]�[�����m�.D�^i�|��yw{Y�������ou;t�.��7���O���+�kqy�n�wVi���ʵv���E���*_���8.��n" ����Ь_(���o��0f��3��l��>�'�ʑ[X���Btw"c ;�J�f��0g9>E��l���b�d���Ȟ�Օ]����d:q�3L�};.��s1��.<�w^�2߻�wv�"�&���L�L�:/ �k�7I x�[�$�ɖ��Ծꬰc���ˆw�F���-a%bhi[1nr\p�N=�٪-����+$�i��a�D��c��d�;F�$z]��[C��Z*R��bٶ�͜Ev�Q���Y���3z*��Z�
�\�0'.�*����Z�N�ɻ�:�gY]�7%Ҳ�Ͱ��vT�n-9��v�	;.ǻ�7h+.!C,38�|�a]��(	�+�b������]��k���k�6u�xA1���sHO9��oKEU�^�*W���4�Mმ��d[��L�f��Ɉ��um�v#˧��N���Kf+�sHt��t���׊3�:�� �ʃ�7�ѭ��D��@%{�j��u�\J�y�� ��i6�$�A�����BMչ.��8�#Ѐ���,�{�{4�.�w�Ն�C�^�E|��n�@}p�Q��eN��n�����R\���jO���h+8F�2u��=��\���e�B0�+��mS�y��[Ǵd��q�Lыg�'d��f:�{�`���9��oh��B2��L��(�03�ŀ�I�Ug>"mC�ǭ�`�u6�h�;�aEk�wJk��D˗O䓼�Aچ\�/�%F�(��ܰmn��\۸�a= ����Go<]�ܹÛ,�T	x~}�2��&�x���j��a{��9�%<�V��!���֮�^Hh�LǸu
qE Rز��n�цs��`3V�o�q [j�.L庬.�%������ag-�<����bl5ٲl�Ӵ�7sM��3TV(���Q�����^�7�]7:�f;0+�$���s�$�ܻ��"�!���Dqc�,�Z�b�sm�, F5$v��P6I���퇆-u�[�^X�S��2
n7����<���Ujp�1wl4�l!���R�۝Q�gD�ͷ����lA����i֎-մ.p���T�,��;l�2��� �`��v��M�AT���7�i-r׻�ã�,UZ�q�yi�xP�c�w$���e��>�V���3��ط7E\p�G�t�u�S������!Wo1M�η5h��lz��vv����A�(�vMks�M/�7{U($��[倅z�z����]1k�j =�Y�ε�B���#2'�`�%0o7"TӚ"����Bq��]�
wn��u���&�t-|�ms���#���ۼl�����a�k���:�A&���rݔ*�b����~f�7����@g<.m���p6X���a�5���RR>�7;ݯ՝�K"�T��S��^�:�ҏe���uK96՜雥ct��"�V�yb{w�G�G�kxg|J�^X��8N���J��a�Q
�gbl�Vj[�M;�{q�h�>���nT���`��e��������z7vaod�~J`�s�<mؖ'N�'�SS���^�ۓ��+dC�������k}����|l���-�a��Y7o'�C�sB����Ȗ	bkT]��7a$`ʷy��S�s��Ë%e- ����[L�8��ep�G��E ���>ܲ}�t�SR.i}X�F9��w��y��W�șh�2-�;��׎Ww(+ȁ۳�jх&��7f����k	8<��k��-��K�۽f.�j\�廑�-C�`~��)q�s�"3��qlI�ql뷞]�qB���D�(�E��Q��E�Z[NT����M�i��k-4��A�o�ô߂�'#������g6úM�D�nv4�}����/NټY52�40v������+ٽ���c&r�.�o���W�A�:4vH�ujJnn���wI"hJ;P�ҡgS�����;-������Ϻ�wa��n=�x�I���gc�Awv�]�tӝ���:<Z�g'�v��in
:'�{:�`Q�fw-�oY�;���ѐ�y!\ͦH���^ �U��̪��TNd�ۜ.ɔ0��t��*�V�L)gd�)�s��� �`՗�8�	��#�3��K�O5m �%.��w>Za_(��j	Ǥ�|�lǵ��)6/ZJխ�$u�;��;.h�� �|�׽zg.���q &���lcQݽ�gwF�-�U��'���w�X�A��v_����N-Z�ir�Vnʳ��xu�݌77�1��=���ӄ3���y�zҋ�qr�>�g9Z�G]^F)�::N�o��;ɶND>;��h���ǡ���~6�u��g/9�˱邞����$į�$�N.��;ݢ<X��7�F����y���M���G*�'�u���w�35=�r��wXYÍ�Ci�DШр	1 9�乳�^�8ʧ��L�N$j9�L\w�B��.����q�n���4PM���V.�転�˱�ӕ�'v��qe�t�_�M�ǥ��\5jW��-[�����n#�ˤ���g�A�>ǡȇ� �H�zh�s#��>9;�Ve�u��jSU�U��ܖ���Y��hh�w`F�J:9��sw� �C��o�t���4��PVҦ�\0M9&8�����<��j��P1��gl)�;yI+�v�'JzZ����\=�8�H�$y�h�@�Yki�=��[+�h�;�L%��0�7;�W�Ǌ���˷��[9�i�.�5�I��u "�uoL�{��z�'������ ���N��k�v<{󁳏Iw�8c�϶%`sy���S���td���:�C%�M`Î�Wy���y�{�w�ْ��`����X�	U��vgN�֦����I��0�:�ar`�	`��	�8���gS�E�5C�8ɲ$"�U��i�zE�4�Aݏ@(68Gg��u����eb5b4J�Q�v����o+�o3˅ �ܓ�1e�8�\Taݖ�q�:�P��퀱�sv�&��V�%'���~���Kv��uȩYZ���u8�����d��ˮ��aR�Qi��i��{�W;=�,�'fۍ�&�*�"� �����(��w�7~OJO��Q,�u��a,�g�����Uym�������:t�7�rł�t�|6�6qWyq��K��8���x�q���p,�mi�K��\����FLiЖ�؎X������������+��֢ZO&7��Le�eX��\ئ	IB!��w\eaT<���k��$�"�2f��]��wƅی��uu�
*j�bW8�+]���V#5�ol������<���ܸ[�������үu�����ߓѯ�I;��8-]3�'vB���7y���Vj �ݝ0v�_��g*�ǆ�֍yė�_��{z��)�����p;�Z�ȷ�^8�׼�;�X�fy���e�m��7��j�t<��9��:�[���Ց}��z�0�0L�����C.���j��Xf�Sr���a�P;k2uos�00�c��x�\�L�Z�zx�]�u����[�[#4��ܹh�X�,�9�ܹ�os����o]�:���Zsp�ȽX�rǅ9t$�%X��u���!��z6��sh�&鳻��;�������U�-g�}L�̊�8q��+7n1:�Vltvu��uo	�qЎS���o%��f�j��r5w)�n�)+7$�{��X�>�;�o	�*�ǋ:ɺ���8�>�jk�f���wr���
"^Wsn��7c�N#Tܪ�V�5ガ}+��:���ʋ#*��9�{�4,:��!�.i3���3e��ޘ�f�Ȃ;�`�)wR^�T�5�5�l�5�z�Ó4nnط�}��%w���Fw ��8t����pMv��C����sX��օi��fV�
x���G�z>�7,�K�n����O53lU�\w�}.s@��� d5�8_A!�w"�5ы����	�Hz���9
d�œ&k�jUӐ�/v���5z����uXN� *K��N�9^���8pp���X��N�Ͷ�Z f�LCyw6��K�M�Jk�޼�{i����y���~s����+i*N="���Af�rb�<�;~=]�GX�k�4w"9$.��'�i�;����o��p��p�5:���f�ܼw�6�ҍ�"e��t�����4��M%�3����F.�'�y�욳K*r�4�7s\�jɷ�؜M仏	pv�����l�ݸq��U{pq�v��b��ِ�t������`�ԋ��7��[���_\��Ō�<
d��&��t�w�۷�ݬ�\;�O-~ˬ�y�d�[���7z�"t�;8y��e��3f^ލ.� �>Os��^��.������x���˱��֟��N��j�{vQ�sYX�0���K5�=
d궘�C�𷰴86�0i;�w��1�}ҏ�Q ��j��:�}ǖ!��ǧLf���SX���:�I�t���Ђ�5":�^�lp\]�"����u	�ʈ:�oոۂ�]XЦ+;�>�Q�G���)Tobj齥O��%���ݲt�h�O�	j��� L�NY�+Μu�s���=��xM��0��:��9���m{��s���Pi��
\a��n�gL7b�gE����x��`�3q�B\KW1��L�3�ZwR@ua��8^�"���S|�@%�g*���5r���8�v9�8��/ط�kZ�ٮ=T�C����gw�î3ڷ�ݬ���>s�gl����9�F�o;&�v�	��Z��(^�A�}��=��kz83�#8E�n���䝻wW%��gf�Z��V�y+�r�9/Y�j;3{f���W�mX49z��D�؃�!x0G�w��혦��ټ��q#dߎ.�,z)�r�,�Ǎ��7�C���ۆ�>A3���zg�Vn�N�I������h(�f�n��̊��no��﹟O�m\��4>�u��P����ẅǓ <%tn��� 4�6���(��� ����2z��h�z��G4�Z�q���H��3m��u�(�-ð�ۖ��f�h�e�Ż�1�(s&�O��3��~�4��K�-<�]�yꘙ�M�n�:׼0A8�2}��y���q�mS%-/_X�:q4U��:B�_��=������U�p�M�d`�����pE8]K7�=���oC;�$�r�͂=�lE�ZB��:�o�i�O)� �y��
����}3vSV:�t�f����+�n�Jѽ�1c�
'���C5��%��<{4�ke���v�t�Ư���<:�_̍�ݽ���u�<r���ڹn9���f�Y�rhP�jC�Ѣ![�k��!5~@���Tk����{yd�C�M\FBI �k�}���4<���M����f0�����E�cV�Z�*@�qt�q�L�gA-�z(!��n�F���;��Z]z���8VR6�x��^1�J�9
+
�I�͘ฆ����N�Ә8&�ܻB��y3��N��Z���!�#�B��ͤv^C��C�V���u� �w���Zh����]c�^�q�u$�<b[��.ó�,�����_�����tn��c��V�E1�lZ�݊�����1^�ND2�h�7��"��S�n7�gê&f���.���,{���P�ջ�"�z�w�]c\z8b���ػ���)�$R`'��(U�T�nnl���
BWR�,��$iwN+�p\:�޳C�{6�@}��9�V�}��>B�ƙfF�!*͘�Fn���!�r��!9!�f����'���E�x�rb(��×,R���X;��MQ��׳�q�F�>�	�N��l�)w�E�s�>�}��7Vk&� �WR����oe��H�&o,�w���cVc��|�Gס�܆j��^ћ��.�F���:�O;�paa�z���a��N �@-r��2���!ڣÐ�;`#_�(��N阴EE��[�t#��[A[�\F��Y��$��ٺ���5����U�G�����{������Ds����4�1`}wA�6�f�e.��oBF8C�<\����e���n;���r?g�u`���{�3&H��!�����N�=�������Ƽ��OC=�LM�vI	��YW�a~(YF!����}){�4��6��f0�o�{���y2:3�3���v�ۨ�s��(×q[>��U���=N-����&�ݛ���Y��!��G�G��1A���f�rֿn5ӆv�D�����ߐ�=��˝�-k����/]�+[��m�Bg|J�y�o����������~��~�����L��j���D�d	�Aj"��(H�"PA �� � ���Cm��������0i0l�0.2�N��M�0aL �*(�"���-@N�e�����`2�i�Q$@@	�Y �DBA@Q�IID�dTAQ$Qd Yapl�\� P$@�TIP�Ed	6 $1�ƓP�P��U*$� 2"��Ȃ�)" T**-@@���*��"(� � �����$�Qj"��"� * *�	�v�Lc�������`������W�Lp�I_�Om:�����o���	O�NayN{A�8 Z�X�� L�7`d�K�C���>M���|N���Z~�o��|� �y#��@��0����66��B,C %����6��_7���.����HC������,��cĞ���y��=��������.�  �i�W��S�� 
/�����|=��~7�-�VV?��f�Δn
t�1����� w�|<���:�O�ݡ�E����u�Ӽ׷����F0��5�Ϋ
s
(7��Y��_N�����,�r��BE$o�s����t�t���N����W1�^P�y��ٛ�� d��}���H ͉��ϕ���N{|ñ��Y�w�|uu�07�|�.����ɲ	��n��L��G��#���<����-���s�윝�8c���s�;��`�d��Lxs��K���7�L���oo���B惣�̵g�w����'����X��]�)ɼ��y�f[��go�����"}Y�=ޛ�s�qcC}��=�{������w�����̼�f��h��0/�o���]V-s�`��}�v	����3�z#�67��>���q�N%��?guo=k��3Ȥ��/Y�`�7�=љ�qx {�=� ��n{j�`3�x�s}����CYء8i��v(��י>���-ʱ��;��4��qˬ;-����ɷ�F��{�+����e+Q��f������j]��7̍�b;���'PK~�w��ҡ�m,�",]c��>���T30�`�FK�lG��a����E��-��(2M��=�!͂����v�@̩��n{�!X^���=�>^��C��!���sђ����7mY�R�F���3ޚ����w��&]����wSg.{�f��ioNP��;f<A;p�>{�>�1�]=]k����<'��V���$:5�u���כ5�n��������M�:��%p��S��>o}-��Ͷ�b:�f�Ș�����]/�h���~��b��,���v<�	i�z�+'X��"/|��Z<���3|x륇=�k�Cn���}�^��h~!C���N�7�(#�������x�W��r:����DX�!���z{�X�y��'Ry_b�KJ\%P��}��!��d�QG��zs����|��\1q���LK=���{�}�T��m��mOK��A����mK5�^��L�2n�~��^�%�5hk�;�˵�#�����x�<}�3�c��%yn����/�{}�3��	3��;��.<%���zA#���ya��OINȇ��ݻ!��1T�&F�q�=��o8��3R�ݝ��w�@x��
��ZQ��P@�ֶKZY����np:�)�5�*)���#)�V^�©�ʻ��W��ZVz������y�;@�n3;��7|r��g��ʝ�݇��?4��'�Nw65�9�8H�o��1�^�D�F:��;G��Ʊ}�v��w�0՞�G��1v��X�'�7�3�OhO���k���Y�F��gM�:)V,Ө;��3�x�������آ��ލ?��>�q]��{7�Af��\RQ�o�i���Ӂ�V|gn��^=呩�|X09�HS�G�z��9�a~�+�:�g�}�<;��x�`N�e��s�H_tk{���;�'����J��j�g�/{�t,�q��xq���I��{�R_�<�!*~�E�]����1�7��s�w��(�R�������~�=K������+l�Zm�o!Y���0<��;����ݻ{4��{(�`g����\���7W�������_z/O]T�|)΄-$�f�,����A�z�]�:9�W	���m�\*6k���QZ��
��y����`��˰�"�5Tc�{^]��m�w	9r��=����&`;/�8ۇ�7���l����iok��c?/?gs��:c�$�8w��瀘�7�l�|���l����`�%�pp�^���5�Tv>Y������W�7�y��3|Z��|��Y���лh^3��-�7��x�@{xd=ɗٲe�~���4����7�ۧ֌��}���wf��{+���8������Y��3��Տ�%����tz!�J��ӋeSq����_�^���#a��x�S��qקzp�O\:�{1v��.@X@<���W�{���뽅��q�y�7���y�N��bs�kz8�!�ŋ�*W�Ow���L�8�r����:���s�X��{�F/��o\Z�EV%	�K�	����K�h5A4�MN�[��"�ѿ�A�+Wbʤ��Ʉ���>�5��ALIgp]jcc���
�S�k�,{��27��F�E��3=��i��t�����}��w�o��_�E�WIVY���E�E�N���,|�=7a��N���3b�1��S )�2�|��Ҝ���*���{5���xm&2�m��=�^�u^����#�l��W���J��s�,����bV\���ڪs3,@��ޛ���szvq�g{.��/jؗ�2�y��C<��4k��r:/-�5�^�W�u<&r���Vg�=ᾚ1�h\�w^���=�nn;V���t����9^�[:`f緽@Y��n�u-�[���J��S�E�Q9���M�����M��h�D�ǚ��:W��grx�׽t�9�F�Ν�EZ����N���%&^��=0[v�2���X��~�k_���`�S��u͇�H�#���Q/e{�ߛLQ͍�����7���Z5\��4X�̇۽�g�+�	*�`"�PN��C�=�ȧވ-��k}���`�-ܳ����=!�[��on{�-�������x�f�������;p�g�iݚ���ĵB;͖�v��!X=�w��S���Xx����d�+7GT�ʉ���>1�W�Y�"q�v~�9���������0�$�{Yz����ujcv]+�s��Kq��|'k�6�p�/�<��Ow��l>�ɞ��w��[��Be�������|�������<q���k^�7ڦ�e2�~&�'�0z�=��&�j]4��=z�^���k��J��8����(b�x;;ݚ��A�2�c<��s5��sq����ޜ�WǕ�ko��CR����c�Ϳ{����F�J���c�;ڻ�Y/P�xIǉ%�0���v�*��}'�����5���/<�E��߮�̭�w�V��-0�Ā�N���=�Z}���W���
���ɫo����<�w���p����8����s`��^oU:N$U��>�G=�q\��6o�f����5W2l����G�z`�yz��G,Pwv�����_B�����Qn-��rSl�N�=`{��̐���Y{r���'ջ���.(�h�|�r�k�\���q�R<BH9�i���� V#b݅y�������_�Ná{��]��5�l{��a�1�W������;{�r��d�O���O�Ó��4��ٞ�Z2?+G�=�[���3����g��{'-�9�7��� �n# �t��*7|^�������OG>�06�٢|�o���{ܐ2R^���]|�<�� _(Ova��~|��6`�o�緘��	���s��m�$��+>�t���]�>�zL���B��Q��n6��}��;=�Y�ׯ��y�$��n8�͢�;�
�Q3}��ۚ�_�oڋ'����1�1���<�l�j\<Kǎ3�kU�Z�ol�{�&�h��)��I�q�rStwfɓ�ˀ�����2��<_>��B�t�Q��OY���N�{����{}�;FK����ǀ��u.-,xQ�������9Gf��d�LDN��sۋ9�K�B���v�u����W����(�W�:s�TyuN�>�q����w����Y纻p<x�ʑ湰 ��� �Vz��esm|R��WۡL֏�жd�C�3]�'>4r�<��m�����gzCN�5^]��n��{�&�O#��*�Y6�w���B�͢��p�NW��/�{��meԋy돵M�{�T�o�r�ʺ �.��^�/��={/o:�儐����w��%�� ���}���?�����<@�\��>�����i�+X6ˆ����Z<V�t��z��_ �{M�Qk���L{��Y�?2�4��z0w��&~�������#�ͼ���S==��8�� ��h�.�pI{u-׳'��z�8�����c�c����=V�ױ_s��r���h�����]�����X�r#�U����(�ǻ�z.ǝ�fIk�Ц��ӝ>���Gn{a�c�ޔ��cB�rD�0���4���_j7ŹG��3��?gvn��_�T�OuǶ�N�h>+;(o�Ɇ���,3�>g|��6/L��n���ܗ�~��� �`��%�ůs�;Y�$cqW�U1������o����XZ{p/{������}������/oQ���5�ҕlM��n�U���ڬzn�Ѯ�9�oqx{�F������i����'{���N�ަ��wb�Y��^N��v�g��'�oI3���4M�q�ye�h�$,�8�ݝF�h-\�D�x�s=2K�� �Ƕo�Jv�Wod���7׻=-]�oway<=�o�f�/����Y�=��M�n����O}"ݏG���N���G�Ox���w#ݤ,�U�ÅC�D�/{���S�V�L�c�����W�gv�_��V�hs����������[�9��Z~�r�Χ��s�=쉏	��[�i�/uRW�z�ܐq�����A|��Z�~/@����0�Ɨ�hXwf�׾���{�Wv�����x��{�p#�����6�{�)�ق�z=g���=$tP�z���%����Sun0g{���ϻ۵��ݝ���u'�|�W��.x8�Ѹw�� ���L��N��3t���5�yE���\㾝|B_E��������l:q�>:��)���Vw��򘼼��!]RF�]�0�[�y�s�<x�2�b�5NjihL����ni�J�}�c��J�.��7�c�}�ݫ*�>Y�I�ԍ֔>D'��_#�g{�{/����;�?Y���g�`�F���k��M��]�!���7�M��:��v�o{�ɗ"}8����]й5�Ρ�M�
��;w��aW��P����=�`e����G�������c�X�we�02���3��g�,=gM��y��R-�������Sƥ �|H��Ɣǈi4rhmJ��+e���y�"$�y�:�9��߁:�CLH�еf{z������{_{}��
�1d�/,��4gY���g׾!���r� �G�c��'����R�1a����������:W��I����V;�#����I�Ye2������z����8n����i�@u^E�^>X�<�h݈U�=�N���[�<�w���˧I;ѩ�F����N/O{\h�*��6=��K��=�++���;Ozo�{=��.�K3�28ǊN�#=s����ܻ˴{[�9����׼^�2&y�����]ס��}�U>����/�����݇�熷�]��<5�\F_s�ˋ޵�������u���h5w�oyK����(������S�{�Vm�B���Þ}���^�t���{�os]:q�۠� %{5���^4h{�9����g�f�L�w�gv�W��F�ׁO_@�N>�f�r�����:״i�M�P�75�|w�Π�3F�Pe8�����ݫy��==�3{�Ǉ+�d�W�ov=���B�l�x�;���>�}�����d�|��'p�Ap5cI�^���n���v�����@����7��z��	:��O4.y��.G��9���t!����ط�x^ۢpE"������-���6M�4�����ݳ�9�S���N�5�Lx_\K��IG�������]�_��Z��󊧓���	7��C���1��p\I�"��F�v�q�3��	�q��1�N��}��nQ�#��z����B{�/i|^�8w���t�nq}[���/�=�{�-��P=�x�I�����۽=���y_�!sռ^Uъ˴W�t�hDohGy�띰\}=��9��>��f��ڨ��X��K�D��z/eoG\`�Wq��>�z�%;�N��;ֽLz�}��i�m�n��ɓ~�22�Y���Os�T��V�IW@�B{#���7F����gw�OL�o���8,�p#�L� ����S�~���\;±�� �V��>�a�.���,s���[��	�'/��yj�һ�˨C�{����fM{��_��{��ove�ecݜ�o�y�V׽D�)|�;���_z�|I֬ᅦ��������g�YK�2Y�P#/�"p��o-?E���LK�q�xjI
wRv����xG��B�!��u�/sX�_r�^����f����&���^���:����-�E�UzW�`����0z�3��Z�L��=����sq���=Ҍ�@>�z��S�t��sj���_���n���J{�9�~��Y �3�������׶uΦ���cڭ�%� μ���S��/��76.�{�2���_�5�������t�Ƀp�7��1T�މ���`��-#�n��vW�X3���Z<qR���'w���O���^���;�ӂE�)���Vm�b^�L�t�-�:����c�a��M�d�]��ɾع�����a�B��D�V�"����=�.�q�[�ĺ@�ox�3��en���$_��ˈ�S�����������I�p���������j���hr��;�J:&��p��j�T���y�Y�u������_i�x�1m%^���6�f������jk�z������O��v�n����ô��/��/n�����H4����;��<s���ԩ��]駻7T��W��^Z���ٛ��:���^�|w�����z�?d���}۾�\k�������P�t���>RoP�~ۻ���9����{�Onld����+7��Vg�'=�c	�sb���:p5X����۸-ַ����@�e6�=���=�X����1�ݷ��{W`�����U+V��V�5�s[�g��?����(��H��������\�+�E_���͘Ƈ��L~���O��v��~������"�a�Hb��О�H�K��)��kv10`�6��Fv�k��� �.�
��,����pf�O���컘�7%�k+\Qj�[��FV\�[H�鑌u-#�.�T0�mp�0��G�a��:�s�9�tD�E�9|f�2��f�	Z�m�%���5s������j�C��\�oM�vmZ��6]uݤu�%��r�\���#-�
Ŗ6�r�3pµŚZ�o<�֊�m��u�E�Ɲ��(�s�X�:�6@�g�wi�n�ت�����\�c�����z��ᶛ-�
�K�9���;�ϤɃe��.�!��w/d��u[�'�Xu�*:9�G�k���]�ٰ�tκ�'=Ms<��>�q�s�:�Ķ4�Ok�ѳ��*0��VR]lfk+�J�3P�0!/mb���v�Y�Wb�ۊ8�z4��=Y
֞S4�ic�^wj�n3[��L���G�.��Nm[8�!-��v:� �V}K�띹�`���{O/j�A��+IY���@*���9��k��3VC�i��c�c5Ϯͺ��\qɱļ���+���=���۲B��gӞ�[���t���z^�\�q��n��ɻ'k��e�^���XB5ʱ)��(���fa13V�:T�7m�+:�ˬъ�J1̘�[��n���$�2p��$�O<���x��'K5��e6l�D�ە"���2�ce�`�.�V�����h�u.ׯJ�e��M�ޞ6���[���c�Ʊ܃�U�c�#�=���&��M뱙#J��.ɮS=M��ʉ�g�������1��y���6�71�eA��^8�(�m�-�C��Ѻf����Չ� �cJ˳��68��|���;�4�B��ԛ�0.���՛pi
���˭e#��Ik�6m���kZ�{B��g�R���e�	,f���� ���>72n���q��n��c���J�������On/Sl��,����-S%���Z�Y��c#���V�5�\��v�wW,�qN؜�Z_f5�Ч\X���	���R:�1b-�LS[�x���⹵v�c=]�^�ܜ���*m�Zؚۭ9���m�';��g87b;<�B�`c�ks/�9_>�����;v�d��@�iZWsA�5�UʻcRҜm���}X^��]vl�sɭz�1��[����qv4r��	��'1�v�\	�c��s��=kK0�H9�P�=sW���e���!҇<d��W]W*v���u��쵀�.�WNp�v�H�xb6�7V��C�7nż�DKY��6,���]��nl�^�*��{u���El����e�Z5�i�R�o	M�a�j�gS�1B�'� ev�9��M��@�:ۈ�Qm��ܺ0����7�R����5�4je�!��gZ����XX#[��$�g/��2�:���ѕ��m�MZ��W���0�8SfM0�xW4F�\]����X�֧�i-;�j'z8廔I�1�����=]�>�20a�muY{d�m�2�Z�V]�(U�`�Y+d�9l {q&+���7��/$MWu ���8S�kO[�>7a�Zu-�)�γ�ڟ]�-�[f��N�#�k�z�R����k����q�]��5ъi��C�a4�&ń���5�9��zDq�����Tն.n���x��݃�2����p�v!�m��:y��F�Qe�.2�N�K ;9K�{:F�tRl�<��[gs�n���dښK��]� �u�X�&b�����!Ʈv,\�.Z�;n�c�����;i[j��a��0m����3\l�!��1��F:\���[�.��7-g;uA��]Wh�ْ�fA���;n�44��l��p���sH&3�Fa�u�s�25]�����Hĵnu,� ��k������R"��l�4L,Ck�	Uҽ4��h[h�@�n��śW�n�n�9�r�̷��m0n{��uïn������ɗ��dh��D���N�5U���OgJ��\6U�m3HƦ��B֬n�	�������-(,��˅���ie�&�ΉtE@4e���iL;i9�x�v�zЙ냷��5���,�`�E�&��lE�ݫJ�V�g�m ��`�۫����c"�m%���	hk��eHJ�i!��P�	�-���6��˓EY[�70Km\�CTk���m9���<3�7v�dJ˲�O$t{�v��J'4�:��9;�Xz�>;U�M�.���Fd܆�ʆ
�2���3�;S��v��M��Ġ����ĸ��v�n9�.5rī�v���>�����4sv���+#����Iyԋkc��5F�FK6�id&�@h�mY��m�z]��i���#沢��ܻ�.����Ge�]uk�K8�cu#s]���f��q�5����۴`zkJnǇ
7�R�t8�;hCgQ�D�2�
59��0*qN�)�
:�n3]1m�%�,�ԘЎ���=�b��� d�O1��k7;&���uN.xrs�^ӝ��u����m�%Uh�z��T��e���d�&.Hᵕ�Xt�AC����N*nuηh
�W:�`�)�VU����d̷n8���㰓�� J���4r���;`���ۨ�WŇ�� �vst����d'KחF��L�#�j�b;s����EFq�:�N��-��-X����f���!]�`��lF���ڻ �cm�-�8!�k�r�Q�jŊjg�+E^�,sm���
�v�p/��x�9�6��=n�&@��-n�vSG;�sg����Q��": �Х
���78��=Kvܰ��팇S����Y��[c�;��Q[����'m,�"�(ˤ���f��J)������M���ľ�y(�n��x��7.��G4$Z�H�%��{g6��1�	�cdy���+.�����Wqc��2m�^��k%��x+[��e�Y4��Hۉ{1���۩6h�X��˜���RQ�G ��-�h��l3X���`,�͐��Vʖ5��)�w��e� �qi���M3@S��#�v�6��SgA9X"ٖ���mI��C;��:���V��$�]��{S�֣�Jx�i$}��Fx����\��P�����j&�$���i�Je[��j�n!�� �)c�4�iu)U&Ϩ�N��^v5�y�n�5ԙfiŃ���16�֣7g�q�Zqmm���>�&��f�K&uwng:̌�	�i
�E��2�SVGe�����fZes��,l-�7cZX�2�,�*�Y�'8b����ܛ�C��	��j�+�h�"�E=�x�j��;�ֻ��w��p)����sƻ��H��ޥ hL�U���̅��Ks�b�U\vM�	�[��i�6��6I��b�tM��I���#��ɳ�7>v�K�s�K��/j��]gw$�ۭ��1V���u�-l�MT�9јLL�X�6�H9{8�1��3��S�9�JU�a۫�j���E�����݇�w�F�Z�lp��-��5;�vt��K�ѵgv��޶���9|��'T\k=�L,�A��N룷�K]k#rJ9e�f�Zm
����� \=�C�s��e��Y5Z�i��E�۸���%x7l�mb��&��[�Ģ�S�M���q���F���6�N�n�̖����y�P�s������9���z���;]�C���:�
XiN.ݑ�Q�C3n��9"���BӲ�5����:�V朖wq��e/Z�&��M��bn�W6�gL�=��uly�N/u�;T+�6������j����mM�a�ٴ�]�`�=�y�w-C�xv�Uҏ>�^��Ol��غ�%m�P���S�6:祑�g)�pe4��n�sݗx���n��)���nm�lKkL�ꝲ.E��GB�[���b�+t���eA�dSp����h
�EGFӋ֗ s���'�:γ��1�Y�̖(�2��-�0b�K���t���iH饎�r�]��u�n���ky�Ip���lic�		X֙�G]�4v�ƗB�eINE���F�{a���"
FO�vێ,����h���8j��m8�7
�ѼOO���f�����@�d����n5�#ے3̜�ٚvw��s�pحu�WU�Ў9��-\�s�BpM͹whZ�ƚ���%8�t�\l�:��#XX�Q��1m�;�uB"�Y��XD`���QnKq��m���j�غ���x�tm������v�R��F�p;���@V�B�n�c�d���'s �s��V�yˏ:�>�we`�Ѻ���N4Pm�8Dqty�-��m7�\t%\b`,J+l*h���#�mb�]Ŕ��BY[���Z�L���.�+p�kwl��f5ua��^G���rQɩ�L��X����,`n2C�{&���m)GUf�4�z3�e1�77���5�`��%4�j�ia+�i,�6ޣB�c���==��m i�@��uz�V�7N�'&1���{Vt4vʈ��2���)m�4.��C��^`�ʷd�$�a�{<	��I�m��0ڻ[nr[W���д��ǍMF�A�u�v3w5+K�Ops�\�uv�gh��#U�/%ՀKZ��u�u;[)i5��-�5!l+,ݙ�ՙΜ-.�O6��;aF��ͽu�uPvm�^"��\f�>}��jp�qڗ�q�a`��9%��KY^l��a��9E{\�.��$o9��k��ԙ���`Xyqۘ<�������nݚ۪��̞�L���h��踂iz���.Mķ�	� lm\fW��V��%���6�Fb�<�'�����4�"W"��(Y�N�\���q�Pu�9�w�8~�3��K�!Ij����v$~�\��p�*��$��tX\t��rbL.q�$P_y�u��"�4�'$"rӅ*Qr�@J�*� fG(>[*6�gN�ΈeEd�s�p�S��N��q��r'��
�;���!P�}�*��H����ʯD���nw�� ��	D,�+IkD�:��OP)��-�G��U�Vj��B�9ܜ�}��@`(��t	�6�����^���^����Rr5�r/$á�#��>�y\�8Q��
��Prny'
v�:��r�i3���*�C+,*�I�&%�'��0P�I������R.i�(�3��\�	�W��	��=���7^��I�2r��J!S�f���<��=(HU���-A5"T"f%#�3"��_%�݇;��c�s�U2�H�J,�-��ܚ�^���:ːs���"��Iǈ�E�ON��S�ގyŕt�\�Ȭ�Qrsɺ��y��r�?	#���~��?'���m�v�����]l"C��oi���i��WWs����n��غ�Bn�s"�]�3�������b�	f��nz�9�<���Yr3uyK������c��+nH�}q	�uǞxG[�ٰ�;Tl��
��N��2�+��:��"d	:�g$e��r��=�����]�t������e3�F4�,�����m��`�fss[2�n[Τ6m�ҨƐz�%ˈk{YC ;=����5�E!�䧹�{It�6;�6�,YCv�c�BZ&�.%n���u��^�8�Vy�bi��bMe���XitL9�YT]�ݜ��{{E�g!�g����u��кUbj��$�q,j�ӂ1q̴��%u؁-��PfVU���,�qESu�XX/,��5���ՖmW��x*V334�ir���-%/�=�`C�f�\�=�����X�ugX�<5u��xڡH��&
���M�tf��R�n��Ic:U+�+���Fk5������A��;����I��=�f6�$X�6s�mc`�hJ^�E��,�۝s�҇*�N��B��:�x��!�ݱ�`Z�M7B[��M�Q3�l�n��s�tU��{'e8h��<�e+�����yh6���7iƶ�%� -�l����r��{l;�W#���y��k��s�oj{�Lg�sh��M�t�l ��{cq��lѰM\bh�7�&�l�����
��caG=�D� �%|7����#�'�y)�+m����4j�\�5؉������2ظm,�t\X��ųV<[,Ί��4vf��Z��4d�4IyF.�\���;��c=.�;��Mղ�1(ԥf)�]�8�t@�i)�a��PC����ǜh�K�4��"l텉v�sGCa����B�|5���Kcj32�5+c�t`��7F6[�W��,hNj㞺��֍+��JLhQJ����/B1�\r�Uq7]�,P7f!IB�5[ay��m��X�e�`qhV6���JIaa�S��F��)B�"ְ��Z�-�b�Q+�֤��e�9�<Òn�K�w����Q�����ff9ҝ,�ؖ����*PKZ5��Q'���㻚wp�q#�xᤖ���֔����ьHYG�ʹ�V�*	-���P����f���7������H����1���V��䋷�0'n��y��f}v����-3�ǋw�͋㜜�}�� �	�>�A �f�P	�d�Z�I�6��� U�>�H;�E�,��ۈ��+�|D�:�fs"��i{ �|f/b'��Z�zHw�q�y;9fE��g��-���N�e�L�u�qA �����1��S1�|VT<����:��5���� e��ਹ���û�����LרG�oe��Ҷ+m50KϾ���%֗[d���Mk�b՚�ݛ�����r� Ō\������G߅K�ܷ]{ϣ���x�+�c�A ��x�o���9f�@ g%��f�cW�Sd��XT�y��|H�/����Y����~G�yպ�����zy�#�O�ތ~��yi�����ڊ�4�t�U�q����]��M�r(�5Y�O��,۪ "<����;�p!��Y��lw;��i�p,S'mE-�@!]�ǁ�5+9��8d�G��1#6�������t��|��C�7
���Ô��EnK��'���L	�4�Ցo�c	P�
��,k���M��J� }�񿵰��A��}} �Y
	�k6^	n�DL�����@|��)��;1J�4����˱5�.c1u�`cb����v-c�>O��%��㵏�N���A{/�I��YR2ciF���z�J	�ܖ�|%��d�M�7A�|���$��j����}Uܴx�srb,Ci���Uj�@&��`$�+����˾ ��� �fg�~�ӆ�����$9��ی��9����K+�2��V���-c��)Ӵ<�ˆuP�֏�?i��Î]b��S��3fy��i6K'�7& �����t�ض
$�~����؆���k����|	Ml��$	a�Pe`�gl÷W�>"ɗ�ǔ�G
���
��	%Q��gb#<O�Y��I �d��H�j��@;r�;��Ӊ��4��חnS,J�[c�k2=���<F9."�7t��\��������X�E�;��u�L �7�'�Z��T\�Z���Hݹp�cHZJo/;
-
�<�ٍ���M͓a��S<�%n�A$���@n��:(��9{jj���=б/�&x�S �m���N�ˀ�����،j���H#v� F�V��5����;y��h���A�Y���P�mU@�>�6ڀH$[r��9�����B�Yle&�L��޼�g�B�6�X�����,�;J��zt�cd�n��ӊYiW����fL�9hc
�ȣq&�k�>{�7��d��a����?x��nZ<a��L���x�g.$�؀H'!��|Hŷ- �̛�|���(�A"E�e��l[ �v"����\�	<�Z����EpƷ]=�������O�.ڱ���{���r	 �ۖ�o2���U��nϦ�{��gg�XAa��fߙ�*���F����s�>]`��/~0�um�G�gT�C�E=G��rlϙ�����x׋�}�1$7��J�:���a��BA#a�֙�$jk����5%�?�h|m���-�KZ�o�c ��=6d��>"�%�I��}&��:pe�Q��3j���g�1q�[D���
|?Oc�$����h�9�$Փt٪	'�2���I�و���H�!�A֘�6�<�fTdN�1>��暧�[|}�<�����4���.�ц�ޣ')ݱ��s/�{O�ήC���d��;��A�� �J�����lA6��]]�*Ef�%���-�u�HPm��oC�Ӕ��^�g�� Z�k/\��lű6���J�v-��ӟ��7�w^:y��:�z���1f�8m uV�N�5���/= l�]�Lޙ��;K�u��S'��^W��n��!wYbi�-r����8�"٥t^c��x�wS1��S����m���o�l���*�p�wA���9�{q�y�s!�r���=uh����I���NX��vE�l㚢��A/'.� $�������-�b�ɽl
�� ����ϰ^�_���A,)~��,�LC�7�UbֶB'�y/$r�b���m�S��Z6��t�l(3�:ł)�:`��zhǷ�I �l�HU�ȼ-�_0�9��x�������X3C��_5�)����y�t�@ �d8�O��و<vi���wt��gj�`;�q,4�C�>н�s៧�C7��ԛ �j�	̋Y��\���������|�����Q,�C���&� 9:��0v���k20]�n���,�������d��w�qv�	$�ܼAȦ����y|{�OG0 ~��uu{"݊�&�r` �J7a��c�5q�i~��QN1����~�R׿X��)=ӑm�p~$�����^��ځ�MZf3K��	�w& �FE>���RZ��"ְ�w�|�θ�0J�X���} 6r���y��PҪ��[��$��n�b7�l�9�H>�� ��,�>/�O+_f#hH-5p �	��� �3n^_[g����p��X��87���F��'�U��jd����S�`��5�g�� ט�����UHLѻE~|��Z�ڞ1�>]B�7=�r��R��Hۃ�mhY�%�.���b��t�|�U?��p>�[/ �;�).s.]j��W��>���d��$��cx�y�c+$c}Q,+A�����B��� �����Jdd�e���[m�#=yr��,���̚���L"	ܴx�}�̵O�ΏJ[K��n:��H�i�4���<�� ��`ҵ�;;�'�ٛ��~�xz�r�S�'�'�͙��`�o�ME6� ��5�4�w٣0H.R`噂fR�|����uCy[�ב��#U\4	ojh���C ��ۭT���a�DXL�9����P�߬�O�@��BP�0���­PO��,�h�N��ꪗ��us:���]0$���1v96�K�r����W$#���K�dԹQ���ߩ�~ħ�Y���*�1$��^�IF��A�t�v��m�>і�
	 �Ur�L���)���߹�tk-�36~'޶$j���I{P#�;�/f\��!N� `��L�o�?�� ���`Ĕ���3��D�d�$|sr�A>��l��G�T���ݞ���M|�n�� �	�ڈ'�V�zi�\�ĭ��N�uo�'(�ra𛽯=��sS݅�K���=�Oߴ�;����������(L�xz�g�)���{ء,�yM9=s�d��H0���~��u{�YN�C��<�M\� ��@�I�Z��Ձ�بgq5���p\941�;RZ�4�%�I�+%�6Z�6��l.�m�bR�	����� ��8�L���>']�TE8��a����X�	$�m���X�,�A�B��&�3,��
a�H�ۃ�@�v�^��룗�Q�ڷ�}LeB����2n\xA$뫸b�����E<��D��z$c���>�_�-6a7�L�t��G����Ȍ:�jk7��6Z�|Hv5�ܵ�^�a����޳&e�/�6�$���-D�b	"�-�x���k����DI�m� 9�}�rhnn��i�|�d3�1�Pmg˗w��Ԩ}?I�2R�����=��/g��+�bo�yd�vRn��?���cIa�K��龱\�[0&60$p����5u�����V�v9^� H��S�:��[\�#�q�s��S�.��il,��ZGY�m��ZGP�5������1s�dv��$�����k���B����ws�ś7�x��[��8"��z7X � �w`�b��u�b���ԖQU��X&�����0��^.��/r�d���� ��u������%��q6��v�����ؗu�m�4
J�����|�3 �X�d)��A�&]f�x��F����laf�SQ	:�$[�Z�N4�Ó��u����N*G����0��ڠ�gc\G��L1 �TA�:K7�vF<T+��|E\k� �/s��$����ʩ�I�Wj	 ���>1�bb,ɛS`dܷ��*I�$�pHaU�`H��x$wr����9�� (�96k�C��`,_��;0�����.�o�7p~��`�f��`���Y?{M"YMhŢD6����%�0�[�Ia��[pm0�f�mVkp0��#���g�8E���"�<kIw. sr�1�^l��m��ϒ.����"�x3�왘8fI� �<�M�.����Ӫ6Ϛ��L虽�o�(9NjN��6���.C��E�jܝ�|����J"���2tۇŕ���"��Ә��U�l�̼�eR��F]�� �ܘ	��g���t׉��̕��D�wf*�v"�<N$c� �m��NUmcA�O�9�/ ���>�I1i	��Y���0Q-��ϲq6N<��$]<�@���  g���S��Z ���0 �x�I�3�̂۶�H:��a�����4�� ��q<��wm׈�m�5>M��{�{��o��{M6�a2n�ᎅ[�,��YS@N�Jm0�Q�8�R�z�������39-��u��NU�A��@ǧ��3okHc:�;� ��M�<UT6yÄY���� ��Ly�L�ʜn�=��A>��&�}���A�����4��~|�-�ݚI%�
S��G> k��L��v���v��Ϝ8nݿۘ�z���
'!~���w�&�ð��:�=�v���C��K���Җ�<��oZ��xI0���~�^�c�$KU�w�;����翇^A{ۣ���7�^���Nݝn;%���H���Tj�z{i�%�<���{���Xtu��C/V��2j�O�t+� ��
N0<���ד<FA�r�t��Ɨ0x��SW|<�Y���#Se������X�Sl
�������_������	*��MæW��V*�w��wE� �Czq>�?\>=���Jg�;��l�m};<�yi�^�sq��%�"�p�����]�;׾}��~C�}��F����l���x�G�����'d����y� �Oŭ�o�Tg �ڳQ.C��ܠ���4i�.���؝�h�v��yOS�Y/������>����?}�y)FbqwY��k�.Pr��ر�]���;V"�3��>E@_D�یi�.'��Ƚ�ުz��o��Yx��?g�S�A��y�]S�G+;}}s`�X1p>��av��Z5�`x��s��������yO�����I(�1�7�۫}�}�Ā̘G_v�YO��I�����P��_,G������f�q�ܙ�|�k�7q�5k˝x@��<�|���� �׎�C��3*���z[���wh�������&tZ%�S���sx�b��cV5�3����75�Q}^qsހ�;�7������uO��͌s�84����L2TM�a2� ��h|m*��Hw{:����M�ϥ��
�|��HH�u�I�U�;���3��3��xNOA��Aoe�>D�R@�p���.�]�D��o4�&�"'�Q�A�
�rB�8��:�-�JN��P8��M �m�`aW(/^{��3�[�r���1'	�^|��'��/{���>�8^�}:BG �\�(�L)�����o�~o"#%�j�qTDqP ��Iz[{ST��Jާ[hq�!u3Āvxa����mQ��9j�.l9����Ś�z����䔝5p�bw�=6c[��5g�BľYs4"@�a)H��ɕ� K� @��Y� fxw�h�����D�+%����mzb�"R����j���R%�𤅭�F�'�k!^O&e5���T��^��֛3'c�:U�N�#��@�/j�y�ؓ���<��<��=�Lt�!�`[�)��g�Lw��鯗���~_��!!!�ގΚ�c�[c��{F��0s�:!��NII�,%��8�$Ĥ���6{�xN�"N����C͔^w�Hw��N󈯞"9���~d�Q	=��NU����yUۙ��w���؀9'���,3:ED<��qF{���v��9��*	L�����j!��� � t�t"$ �J�L������0��(蛈>���{bn�� ��1�۰�E�
b�J �J9����d�Pj%E�5����F����&�����WE$B�*�-ɷ�O�b/~�?�����;�����nZ)ER�U	7��� �x������M��p�T+[���3�� ��7�c��Hb�
 �w�cB}�͹8m3i�Ei$�$-ܸL�vgv��y�Mk�ãU5�j�k,�0!v�6W#�coaQYeXb̉m.P��G��"61��'�1j�h���>�ߘr��
!P�=�!��Avu��% 3��;3^KC��N�G��v!�4%�R�J��ֹ��j"
gG[Z����E�y2��X绌E$s �&���^���m�!��ۇX��I��%o\ǲ5�rD�$���b.`TM1�m��3��~��_n�h�*9��#�oj[|��,���l�	�TN�7���*��I�sX���@��Hɚ�=�Lk�����=@6�E$mo���f-@�* "<������|���ffg,�4�1�|�n���:��;��oa���rv/`TZ�Q7�߸rF�I�J�s��"9IPJ������±�b������Y8�>R��۝g�P���,�V冶U��Y�V&�acC��/`n��\�����[V����esyǂA,ʞ �(�=��P�@DO�]QZ���t�	E� ~�y��� 0���}nC$\���\�9�oLd�:��s�����<��p0�a�o��\\��;�{^�����_�}ݽ��H݄��E����A��U��n��Ϥ뇷v��Kv��͈��|��~�}�j�D|ʉl����RE$��o��	R��
�T+����2D*�7��d���h7eu� 4�V��" }�@@�@�=�y|�dMZ�Z�i'�yR7���T/�[�E����+��g�;��Q3���}D)�D(�A5����d��QJ�k�Ȇ�ҒT�M���W��Y�_X�Hq��l�kZ�/{ؽ�&��4�1����XE$RC����RD�5�=�jռ�^_6�^�����Oo>�"�@:��B����\��[�mн�-{U7��H𢏇F�G��\3<�k�K�lxa�S�B{���4A*PA*�S����f)#�F���E���V;~��k z-A-�����5�9��kZז����q�x��o�b�f-*)"k���5��!�_7�;*b��x�,�%��5F��j!�ҒA*'y��QI1���s���������Z�����\�.�?߷��P"wCN�ǿ��1����*S��t0/z{��{4h�sOy������������ �	"@_y���T���͘&��\i,�^3�:<P�悃���=�O>3����-4�m�v��&����%�fͽI�pL����.�2�r��㤒�d/YQ ��������K]m��f	��B�[',���m@c�K&���c�4�(�Md�&���ZQd���c�Be�+*y-��Ŋa^��]֏=@�.�޳b�
�����p&{nBO68�hq��u�kz0ћӇ,l�fV�^�������˜2�؜�Nk�#�F�E$5�[P�0�)�H��g��3��9"T���N�E(s�Y==�xm��Q-D(�C���m_����D�QE�Y��brZ%���QL�P��b���f�ϞpI~�����%Ad9[QC1
�@*4C�׳��I$Z���j�_�߃����Dy;�i��V�z��o��Ĩ_ܷ d"f-*-@��湌!"aQ
aP|�m"������+.���Ex$���j!����TN�^�C$B�[Ǝ�34�w`��πr$��>|�jF���3�c�Wl��T
�P�9oD1�2���{��r2H��TZ׳�cy�~{ض�r� �F����Ȇ �{�	�sv�^�ꩽ��A9*&��c"��RD}X�1y�	R���sX��v&���s}D3�
�@*5g��E$R@�[�/0j'��o]?>���__)`�W�-6�[-]�7!֖�e��q���s�:e��9�d0P��?�����5�m+j����|Ĩr���d������q޽la�j&X�E$�m�s7�d�<2�_781FY������sMG�Aʝ ��ﱁ���Sǝ���贖-{X�Ƅ�7 ���b����,g�^!ũk(���5��5R�(�{�.���=!�[9f�%&�5k���og���f�o:�x��m+�9�u��x�-{�V����3Eg�x{���&`S�Q�o�02X��TZ�m�����P
�D1��6��|M���b.BG��4�%-t
dvT��Q�iތ&eE(���7\�qx������^�ε͗������u�RGp
��7��dŨE�����b�3�V���Z�-%x��o��J���n;{�4{;�T\��,�}w�Ø�B�Q
�A)��=� �eA*TR���������֔��J������d2!{f����C��N�πr$�Έ>�R��Z���f"���Mr��r��+X�א#D���s��r**	=���HcQ
�C���!G�id$o0���]�K&,X��d��3�����M���:��k��q���΋k��w���W�Jokx;Ԩ��u����R��&��c0J��TB�]彚C0���չy�Ml��h����@�Z�G�m�k��1�� �J7û�/V�^ז�T��7��%C׬n��\�
�V��y=k6�v���æ6�Q
�S
�Q\�{�A2J�S*)!�W�He�>�<�n�~\�t6���[�", �U�d�tİgf0���G����G� ���Qj�{4d��� G� 2�X�*`7?M@��a�3y�a���U�Y9���M�c��o���͕m��O9��ݙ��v�c�T��ӈ0�,W$kU&�.-��h��[�Ϋ���G��P���H�;��Y�Ir���$�>h�D�<��',i�@���/�&s�VL�d�9��
�*�I�o����D�m
�>廪C0��� ��=�c������5�sF�'�մ_jA�_<�"�&}�9�Zͪt�z�[#�:bT;���E���>X��1�s��I�z�S�W>�$�w�b	�T�TRCܯf�ɚRE$����C,B��opݭ�~G��s�z���q
�Ⱦ8�/'MÖ��/Ge���E�[nMl�#���s��o���:�pZHs;�1���)!�W3FH��C��'u��PrĨ>׳X�똥`�[`*�e�QA$s����[��t]�^fj�]�je�6;��T*�6�	��k�{��^IW>J��ICjߥH	/$�E��2s6�3�[�en�]�I�E�zJ�iԱ -����ĐJk_�Y�Ce�����]y�	/-ފ0����V>J&k%<�`��¼*�y�z����:f���I�$($�	ec��	/���x����̌=�f`��{��K�v��h$�;��8����mo�]���Ӻ�sgM$�`�.�;��>���DI��|"�<��[�� ����LWP@�S���3)�f�^v@$�G�i�WELѱ2�c�dy ���2I!կ���/$��vS̭S��e����%͗����<��. ����eܢ�tu��ӻvdm��������۬��Qp] �8����cܩI$���%�	$����y��&8	�q�6oNO?�P	,�~�L���,��Ν̴��N���H�9�E�|vm�F�E�?g����K+�eHI�K�)�	E%�g:��Ꝭ��=�R���;,�fj�]��(�Iy t�̥��3;��=�:UU�
���Kg[�JI$�y��y��|ZA��H%�~'���?�?��������0����y��)u�J�<��Z���$����RH
�
W:bX�tB�RQ�O2�H%X�2O�/a��ư���*|�),�ׂI���L�{�nrw�)���%��DK����!����xlB2ŷ��P����MS�pgu1K_5^ºhW�$�ԝ�17�ڊ�Ot����O.�,��`sQ��H^M[�ۮ�v��`3cn91�F9��K���8�s�T�Lܔ�[v�g��\|�+�ƣe�8�a��r�@qs�6D`vD�K۫V'���۫q�N���i{���O=�ֱ)Ɏx��-k �kpp��mgE/3Ze���1��u��B	H��t��[��4t�K��Q!0c����7CN�p-�땱��뤶bY��#we�r�uA�v����^@n����q����g��f�Z��Ҵ."���Y�׶}�>�c����Z�L����x��ׂM���L��P�@�`��#k}y7k��H����+�v.�&!�\:E��mk��,����J�7O���	�$�9��>H�7J�E������g��I?�hg��r\�t�e�ʭx8R�ceP`$�䳢���R�#����K� �Gsϥ���"Fs=���G41%>��~��'8J苔�H�6�+��A$7:(�3䗪s�Mj��T��`�&��y��ޚѳ~N�]�p�Y�\_���R�>^*�y�RܕU�[�/j\섍�SĄ�KobL�)-��)DqՏ��Lb�� ���%�@P�ϲ!��9�g�PD̶�f.���&(��+�
ֻ0!�אC���y�~����]��-�3$:�bI-�Z)=���x�y�P	%��&e�%9�)Ӳ,LJi�y�$���a����N�RK�	���'��{��/ ŶӇ�(%q��l�Y'�`*�ޖ����tS8�w���kѬ~�_�f�CMGԸ�as��NEC�	y,�y1)�s�L�$�is����F�#6kz�D�+,]�X�>��Y*gw|L�i�{��<��($	X���|��i9oo��(-��0_�|�s�D�	+��P�tΙ̱7�n9�ۨ��݋�O���BPI�OtI�$�ITw=m�qT��cA"�O�3껖:�.�;���T�e�d2$���̡�j���ϝ�Br�/ʩ%䗶��Q$�W�"Uz��UC5q=T1��ty�CX̵�#b][!l^�����Ƣk�őE�A�_��3�%�1f���%�/2�y#�Q�N?B2I%Q��)K���٨���w�<ę�PJ���HIVHR����(U���D��GH�|MVEK��
W�%{'_�I4�ϒ�:4k�y�����Lfh�>�6�����KU^f�ӿD�^I �Ⱦy��I"==�񵟄ôC�w��ם��e#i�G=����d?��P\���gg�������{�Y��\K~|}9g����Ϥ�R�1��;��S�32^�<�J��y��NO�<�JV�i��a~v)�j�l�k�<Ϲ/�PI��dHt��%���) ���AnZ�=̲�J���� �ɡ��wbt�e��/�e$�]�� ��W11�Բ7�!�ٲ�������<�)$�nd	�gF��T�;$�jl�d�a��Z|Gkɏf��-�����f�n8,@���9b�v.]f��b����$�v<�@$����q<ۢ9�렱���*��ZR%%ќ���>�7�L��ĂYX�ٓ��[��~@O�=�d��$Jb��R%.��(��ػ���V��^V�RQꑊ�1!��A
i=u<�$����K;W���l}�搒Iy,�ǂI���"D��p��O:%1w	2�V�����z�T&��4�;o"RH�y�"g�ҷ����.�.�s��"gkhB��̹�J�8h�Y96�	� �0����m�Fcd59� �0���.�_� �����i�*Y��Te|j��y��3T��kv�jǛڪ�5դ��ǄJO侕��N:�7:�o�/*xǙ	 ��́ Ky�$�[zX�<5_�;����0��qE�q����x����'�u�y�܎��x���B�e^&�/��C����w\�K����@%�3"|e �KeoCJQ#)ݥ�!5�	EG<)%w�"@��.G; �v.]f��.�j�d����)���p�fs��@D��m􉐒	 :u�T��[2�$�tp[�D?kܤ��K�wb\3iyK_f'�PI$}S��>dJ	ck��q�2�a%��ͽ�2�Iӯҧ�\Juىr�$M���Ց2p�\`Ig���2�A$:u�T�J	=�=V�6�mv�I �n0ϥ �Ԕ��bSp�+�,�� 2I/$|�y��af�W^fo=Dq��I$*r��f��������5����v�i�<x��Μ�r�Ât�΋�;n�2ox�eL��;�ݷ���.ݰ�i�9%�?���p��Zϋ����{��vM�V����5���٣�<���Y���x�d~�X��W�y��=�۾x���!�{/�&r[��r08�����Ceo��x��q�Y�w��p�{�+D;�F��x��o�kl��b{�{��o���(�v/*Z�놠C�^�D�ðRӁ
vǁ\�lvh�{�-u�>�j�\���uU,�;���_ۥd��ܛEy�Qój�;Ү�x���!4���ˎm�(�#{ֽ�>��eZ}ɽ��;�yI������z�x�G�|����+}���c7
�wC���罴g����:����C\�y���､nZBs ���ޙL��Հw����C��݄�$𝉹�y�;��{�)q�M���+v��ޛ�;��^��u�Q�>|d�I�����\���=S7�^��!|�nnY*���٬ɁSֹ��P׋�Mr��}�p���ܵX���HX/6Ј�!���c�ǉ�p�~9.��>>�����Ż9�����̬��|5��>�����Rţ�r�����(�����v�yӝ�c��FX�^�*	,r���n�j#���Vj�}����{�Y'�^������u}�y��p/#�������^c}����.���Ռ;�k���ĩ�9{��tJ`Ӵ����sb�	�]�`λ��ޣ�+\�p�|��������TW^����%�5���k��3��ڵ�?@r�_���x/�/��x^��Ł?��1��K�ɪ�\��4������g��O���㡶"�{x_;)�m�(��O����?8�~�BX��Y��Jz\��~ۄ|�*y˔e�<���S��D���u�P�"�A����9q�Q��ia!\�n�U޺��H����9fQ�=�$\I"�n��S%����$�Ċ�;_OwUАΔr�ۄ��-Yr���Yk9���k"H,Ǜ�$�nz�uR�"Wt�P���J,�62��U��Y�"T�`�O�T$�ĐKLY�e%t��O��S�2I$�.�w��{�Qr ��*�"9+��V��;�����".\��!;���НR�4�M
H� D�!���=�YW�s,Vh����e�D�2P�Gt�H�\*�}\:As��S��Q�	���%�G+Jؚ��s�~NeW@�����b�I�G:S˴�z5�!�N���'PNr(5PNih�XRT���2ު�ܐ�r���x�u�� L��N�<�F��*�A&l��@X'Ed��ƴ���3(y:�>|�9m��S���X�FS��̣��������۳&���4Ml�GMl�.�:֚.vc{%-�b4зR�	Zb֨ش=P�v�Z���!{[{<���g�䲷`s���\m������nx�͸Xi��؋iz�J�oM���nzT`�v-�nevܻW#�3+����,,�5f�θ�e�����&������fN��h�(WnZ���۔�T�l�pS��[ul�� +����.���]�a緕��M^�9�i3r����L��4����kۢ5��"nsH�����Xs��<�%ˎ8�Ŵ��GH�y��6�h���KX�=�Z�k]L�9�bNi�����tY��<s�C�Px�8pa�ZFd`���t��VT"��m$����q&�Ǟ܈���ز��W��CN��s�H�����7.2���ݭَ�i��M5�f�1֖zx���谝��t�1��Tvfp��Y�x������X���'1v�*�-���P%�in
�������R�.���;o^&7�y:8NX3�uy����є6��]�
�=��<��	ճ��tvg!^�Xѕ���k[]�^) �^9Jհ�.x�ɫ��魝N���U�+�Y1g$�E	�-�ҫ�e�&�l'9棜�Ա$�Nt ������M��:��A�]eV5�ɇ��X�����&�d̠�j���u8љ��siM�+���l�hn{e�r��v��;T&���jg
WR]yc��y���A(�.N��.�1l�ݥ�R��6emt���Dɵ �z]�FXJ�1��\�w[��9�$�g7In�[yD�<��m#6cY[�dͽ���f.B^p4�ه���u�c�S9�uƸ�i{�v֭]���fN�^��;g]���S2�vk��Ͷb��,��ɍ�%�1C�R���Om�7i�ɵ�6�)s���n�ƺ�`X2�ԝ'q&��y���;�l�5A�]�����5�&�'f��{�H\��%���+H>+^0m��gb��������R�^�ܦܹ�k����g�ި�����J5!ئm5qt�l��X)��-E%v-",�ɰO�m���6�5�p�kb�ݵ�Lպv5�a��6��;���/6�n���s4s���CLK�Ў�7���{c��W14��8痩��f�o7:kZ��S�X�ҷT^KY����k�|Hr��4��%�*y"}ӏ��A$���I���En0�B]EE�I��T��eWN�J��kIp���p�t��WY�"R	cLo��ӜkS��y>^(�:q�T�����}�y�	G=�on@�a�u�"RwC��H:t&MUAv�\�$A#�x�)x �W����f���!$C�_�!%�Kzu�ϛ׃c	�݉p�Y����w�6��ՋY��1<��)z�Y�+^g� �G�l�e�y�CU;�n�K�[aH	-�iN�1.Y�`�
��u�ȔI4�:^zb%v�Mۄ�k׹R�H�{6�D��K˛'�eG�V����~��z�<~|�v�l�����,�[���g7l�`�+�kf�6Lj�ϟ_��B��S���q�d2I/$r��	2C�'�I�әu�GT���h�i$�K6u�	H_���2�m�t��5ݠ�WO�W�����)�@�WL+{�a�̲�a�Y��i���B|_��o^^���<�m�|>Wxwf���L���,'<��^<��1�X�21C��.G�������$��f�ǝy��	%�<|�J(�I��Ɲ����R���dg�N�%ޞ���y��K�7���e�^I��HO�(�3CⰒ	]<��(��c�)��2�k��샖b�v���Z��ͭP��I���ϥ�Kz#�	$�ٷ�V{:�C;ssVQ3��^e!v1��ؗŚ^|׷�����_7���/_�Q�'�k_1jjU�~IZ�!"N�?�D��^��RvŹ��R�A4*gv�~&�^*=v\�h���5���a����[Dz6y����k��8g^f֪x���H�!�T��$�ӏ�����������2ɗx{�PH�u�q�),�!��bΊ]��z晖I&���nvE���n��ǃ�$͇����d}.q���W)�a�|Sn2���� �*S3ys�:d�ڪ�|��
PH��l��%��7���z��F�u��ٻ9I='��3-�%�=Κ4O7�����҄�٭{CaJ�Ņ�ۯf|���>�~�7nd���sT3����� {����~��%-�#��Wy3$u��)*��`3��gpP.�ҕ�k�	�˪q����D�s̩I$������^Kc�ϽL�{C��C�0��i0Ѭ
$0D21�)�T�I5�m���s� ��S�e$�Z�(�J�7����x=���౛���w	�7 �69��6n��oO+��ͷn.�	�����>}�\�wb\3nrU��$����$2^I �	tv�ϒݗ�����"��I�$���Q8�Ts9b�0a"K��h;䗮��v����i%����D�)tv<�QA)�:hn�+2M	G%D�v%��pR�	��e%_����漉I$�ӑ���m���I{��%JH$N�k̀�UJ,�s:�A�U �O���MĒI�ֈ��$�Iќ�#��%�1���+L���C8��1��X��ɹ-�8m;zf����^������Ue�g_?byk*i08�Rx,��F?)�׻��� �s��%�T��kA������D��O��y��I��ؓ1Լ��O>ܶY9v�BK�/$���H�䗖�t�����:�[���D5T�I$�nw,�-ǌdL)շt����N������g��@��U�,��&e�B��Ar�;1Y��ms 2A_��ܗ�J^I$��t���y��}���s��/$K�s̥���d�b���dY��.{�)A|����`�Y���C%�H'��	���헑2�K^�SXn�Zϙw�E��Ujė�$,�t��p��=2�%$�GՑ� �����������W�^I��^D���]�Ҽgҗ��G$�b�H	��ӯѽՓ��&����I �n�y�H�;#$I2�:�+���%Ś�O�2���C30�e�L���$�[eyW��v[L)R�L�MWq�JrRJ���@��"	��Wm?J������ɺ��TN�sU���`|[ԯ��៽G�����g*򚅬ƻ��i���Ҋ��b�8Ӓ�QtA�Ѯٺ�w�1��TI�r3JQ�Ɔ�04�d�{�x8A��I�����nː�;2�7]=�<6�S���`����mhf44�R�+�ƉSm0 ��7g^F��N:$x� l�t��Y޲[����`��������r���K��-��&��1`�xݰ��jb;J�t�s��G�4���v����+�-t!FU��/$���:�e�oeڴosȓ]��nF6�װު�\�z��N:ݛ�@��h���_M69��۠�d]0ke�/�����%�[�J�y�}z�y��D��ęHJݧ�D�i[�=B7"�i�x����^YѲ&R��z�C�b���]Z�5�XUb�ed�Fi��L�����2I-ڎ�) ���4�U5���K8k�.Yݘ'�4�:� �	V�tK$&�eN+�<�OKĿL�{>(���?J�W��:NS8E�aB�*���u�效YW�[��>2JH�zHH�c{]�&A[�7Ē��(��%g�b
F$�b�Jk�5St��$I Wk�SN���������\�$�^���R��I(�יM�[�\552�2�>$��wL�v%�1oϛ�#�c���fS��Ena��j݇�5���#[��������.������� ��I��[��ϒ%(�גf�E_7r�+r��"Q%/v�d"i�Ap����8dYቩ�}�Dz�*��iM8m�pfm+�Hs]�&��nC�7Y�}�y�f���'�,�c�2h9���e�ZD�0Q�r�qf�n�L�U���u�A_�@$P�G�7MřI ���J�$�D��k�$�=SM���ȧ}��Kò��.�vb������Q���3쇑)y$���h�*����g��-�� �I%��%+��d�N�C8tY����n���ؙ�Ȏ���ao �@,�n�e%�O{� H@$�Z��\,w&��x$�S�ҥ-�)�',�	r�Ț�U�O"Uy&I��$&��C�}�T��h$��?L�	�OY��G_��*Er�Z(W�~��k4��:A�8�&�0�0����\���E��v��I�)��J]�K�8�� �	�׃!$C�6Dϒ�}ۏB�ѫ��Dϒ>E?g<�UTIfA��!ٝ���x$�[e%�o���c��M�mx��RK�=޼��� tF���Og�Q/�!�[���i_�������gb��%���%$�[��8��	$#ӲhŖ='a�C귾�iF�C+qR ��:�zww q�z�g|�-�#�(��մpE�e
�PK1��Oa�Գi�
���4A>�����{�Ig��ћ/"Q%/���"R�/\����`ʪ�]��<�,�kw�Έ� �7U/2��A$:�8̄�K���)m�0	}�%���y����lht��b�jzK�$'Ȥ��ؐ�v42ރ�]�J�-�|�&��T�y�$���ҥ+��A~{����Ⱦ�u��hlCC1p5ʴK���j�����kneKpLَF��H���?�k���.X.�K.��Ґ	 �sl�)$C��H�]59R㚑�/Ͷ�%3\��D��|�� � �jN�f!ܔ�SF�J2���-2q��$�K-�Tϒ ӏ҉$6���kXw5��\��]���\��;j��O��!�$���ȟ2I$��S��"�]T�ܤJ櫎�BQ^H�n�)/?�k��Ν9w.̙��~�u��>�|�>ET����)�3%t���A$�����i�����B,��S�ʩ蚐�&qY��C��}��Z����9�v�y?cw]�i���J�Yj��ʫ,��r��f:������H�/>5TW�_��ě|?c���9vL���/�]K�K��q�V����&LBG2�^fl��S)$��m�b��	lv<�P�(��]��F��&j�X�iQ���nU�r�b�R�ˮ���N,L��n�(;�,�Rf��%�ѲPI�Vt1��I���! "kc�_e��桵;��S(���k�i�IVH[L�9L�,
�%�r�)�f�)�.���Y*����J���{i�e�+� ̂W�/�	,���-F?\KN��)> �YN�dC�*O�f��
�I"�8�% �,&5�wbN�:;t��Y-{,L���]ӯ>��QY�s�C;`�UI>5w#���y䊍��I�WQn�� ���g�$�	{qG%Ut��e�I�������: ��3�/id��%�5F@8�;kBe�wZ��o�,I3�gG��]��L���鴄s��\����fA��7�
x;;���� �A��)���y�r�x�|�9T#ŉ{q�}3���W��2{��BJE����!p��w��4�8I��X�qJ� ���eI�qu�p��Gcv�v��Ά�#�u�h��u����VM=I�^ء���� 5F�\Gf;r�g�J9��L5a� 	��hu���j��*�[�o=U�9��U9&@
+�{!n���=�x��&�"EɈM��m��XNP[����]�ָٽ��.z����:y5�0]P��f^�ȩ�l��w�f���l�<����.�q���e��t�	×d����n���Ig��kԢRJ���	dK�eOơ�gChI�U��>����(;�,�RM/ $}ЮTJSq/5yEF�Q÷:�����	 �g^I�$��x�2RA ��Ćn�:�[����S:N�8b傡U�n^e ��U�!���+���\V .�oZ|��)y.�יE��x�2�@E�����ȇbR�M:kK�h�Ӛܺ I$[�e 	$���IRt�������r�ϳ-"o#�Ǫd*fYà�vKcOo�	Ib]Kv����{�	/-�Ǚ	��%���	���k�iffK0�k����E��ם�c
iLd�M�[�%���@�ٍ�[iD��������&tggN�~�J�y�Q)-ƍQ)$��Z�X��ٮF2��rI�%�	E$�ͻ�	R��!8r�3UP]��e�	{�-�Sm�ף�d�y�֠�?��r�}����`li}.�ä\����N��wP��[�F��3�o�]�`�؅��&�N����1?x�=���޿җ�^I}��|�	 :Z��|��J+��޴Fb���[c�×`�w)&��%��2RK�T�����/]ZE$�_ֺ��|�$�5A2��k�iH@$�P]n\L�˖
��	G\�L=̇{�� 	F���I ��KnKO�K� ��z�����֨{��X$��D�$JJ�^.K"�JJu�蔑��x-c+"'%���^fg��2I �-�l�I%䷶�e5!��I	`NCEXe�D<s�g!Ng��-�M�qH���DMR��QH�B.�v��8"Igr���I�s��<�	u-ؐ�A#���>	D�[��D�#���}(���n�iI
��%t�;r�Jdv��Iuݛ�"�+�fcƅ)$�]��% ��S̢��/�}����M��rR���Bp��0f��������H�e<�R�D߄y���x�����8t�˗I������N�x�?S�]��N�J�'���P�&_b$�ewuT�S��n�F�h�0�G�c]�Y��h�~$��¼p)�e�vs/n$�OZ�M�p2$��w��4'��9/#�g�|����D@��v���xW3��NDa�Y8�\��Vl�i~�E��}SZ�u��x{��p3�9�[�g�tt��)ٝL��էs���tw���vyg�$Qi�(�,[�.=�W���޳nZ1	j7k�x��;�xt��b�!�ol$2�J=�l|��Y{�B3��~��T��������on���e�o{W�A��q�۩�}���{^-U{yy�����g�2���!$�Z�3�3��4<x|�dFz�����䧜�<��� ���g�N��E.�8S��;&k��x�^g�|=,���%^����E�*,����:��Ã]�c ��r��iܱo:�K5�}�]��y�:����&�-�W9bw�5z�'�yQ+�� G(��g/'�F?I��;
��_�Uo}�s�ڵ�W�e5��^�}�Y�|���+ޏ�x�g��:��}��hs7Y��[�c����T��-������T�����@��o��ڏ�Z�o��1����}HGR5b����w�����|����4��E;��	ݶ�r���g�Hh�<����Cu�>���y��yjy�p���>�w�zt�����ѩ�Q�+=�����뒜P]Gs�)�����n�
�<�b���A��0�ΊA��	�k����2��	�ID���@�Ra�%y�9N�-sf#����)x���i�K�S15�<JsX�7�R�B,�z�	��HE�Eh9�Abm�e��9�.���O*�Յ��"����t3"(��G��41MRWw'PH�����Z���$����j_'"����Ђ�V���E&VI��y�}@��\�R./�Ȩ9S|���u..�ϛ��F����e�]nTR�)"Uwqs�r�D#0�T�����t���f3t���"�(2.Չp��$����S���T�,��b$\-Mde	��T�X^fOSҒ�*
��$醔ˤ!$Fr�C�Jz��&'""�Qf:��g%I�S�1�w]E�8V��0��q����I&O�B�*�
�������H$�ӯ��d$�W���)y��9f�r�4��ѯ1N	��4�L:̿Hf@$o7B2����e$�.8���Y!��Z/|�2^��S������:g�kJ~��I �����e.�*�zM��*BE"��SȔW�Kr���l��/q��3t��N����v%G'TN��Q��tvf4����3K��ͱv1�}�0����,�v%.�h���2A"NvSȔJIvTq��SZ�+{~�lz׹G�7Hgt�K#��JV�oȐ��UT��?O��r�e�wa63��ad�U�O JI#�]eoQz]dagh�š-��%�'�'�'65��IvVĂ����'[e��GP���T��H�ݧ�J+�%�]"D���I��\�&�'��`��i�̮h����"�KUt��I/.�7�n$L��Cfߥ���b��kw�:��/Wn.��qD�����/�ys=�d���T��'�P!
{>�(���a��9S6P���C�|7��k���k��뢪|�� ��|�
�s�})}���;]�$��9?>D�$�U8�D�M�5s��J��I�[wkL��I-��(����R���]��Vy�������<��Mw3j�	�V]	�����q�؁��.lj4-sн���s���&�"�p�
��@��A*��e�f���RM=e�.&__$ʞ�����J�D�(��G�w ��)D�э�,�	 ��Y�T��:��I�Z�$�K��D�I%�~�!$�hn5��sc�]��U�p�w(:oUPJ:6$�I%Ӎ��2%5f�<Hi����z}��+�:�D�(����RK�U�'Ƀ�b�%.ݗw͆��	���r����M��U	���O>ʐ�(%�<�ԙf
df�I/+��)�юɈw.]��5U�mFd��3y���y�{KZ���^��R&|�	!Rג��I�'�D�=�\3VE���XVyc;KUͳ�u���������{ac׎���m<2J�{�$e�]�+�\X�Y�2�Y4��S��+��"��Y�L�:������������������;��0H(�� �� !"!sɛ^ם��}�.;pN�w�5n]�z�;�kp���He�a����Y��F�9bm�*��BXU�B�A�Z�i�A�:�ݱo;x	��lA%5�F8I�]aP&Ѽ[t��n�������*�Y����λm"�6�lN����4.Y��e�BB�Vݘ�SX*0�Y�[�m�s�"F����Ȑ	%�n7mɠ�d��D��M��c[F��BUv�JE]�K���*�cjE�.� �h�;�}����d�8b���ܺ�2�^J�^ĺI$��d���7��-#��+1�j�"Q%{]����fH����vp��-"i(z�(�����q9��LDa�I+v��&RA-��e"�m3��s����%!>g;(�.��v%*��t˥�fo$y�})$�M�����z�d�Is����I;��"R�L��\�;�UPI�5�k6��s��O��LK��I.��I$�����y��6I�]�A�u�!2tC�p��5E%����K�$�s"A���y\*h$��&X�I��eR��>��;*�	s3�����	j��2�%����ӹ�R(B����{i6]����ňw.]��6w���] ��F�u�R$^��2�S,����"�����0K���JC/K�r���iy	vED�A&�C�s�)1ҋ�q�;0�ޜ�_�&��׆n][����K��<l����Q�|��y��R�q���#����M��.�G�\��vi� ��x{�=�YD� II	�^����#�:�)$��~�L�&z��=�y�^]��K�D���w���*�P��2�&��f}tK �s��|x~	��;ek^I%���(��[`�cP���I�bR�M:_��(o<1f�c���I$j�})$�C#`D�Kگa�Nc�dWL`U�f]��@�t�+��>,�PevKG?j��	k�Ȑ髞U��l���I(뗒d$�]g�QI-vޖ����ҭ����Ҩ�(#�_��p�'p:s�:C�
�&w:k���CE&ݒ0�ipc6���~~��E���8vr���<	я�'� Z�,L���_�c����,���I��ц|%!�Z�.�˦d�T{Lc��Ǌ�����t�)�[�"RA$9�:Z|�	I�Q�s�)�.��|�ޗ�$���iyK�*$�	$��t1��Kއ/AV��F��Y�Eѹ�������4��)�rN��IzZ�?�r��?~��G�}��9y﯁L]�O���=�1Ů[���O�� H�Ȫ�  H�H �9����UT���2eO�K�l�X��$#���bX�MB�%��h�~ʶn���I%�7e �̋k��e$��k�!�rޞr�$�+$L���",��Cyؔ�SF����($z/^@��ß��5;dn��	 *7�L�$���(��K�tƼ�T�ۚ�O1�)�@��h���wr���.���!D���Nt�u�ܯ77�X����6��������џ��<]�W���obA��1�|�����	 ��I":�*�VNȑ(�$�>>�&}U��'�g�)�K�5��Y�w�՝C#�O�+�/$���PI ��k�$��6gl)1��=Ä�;��`b�ܹt���T�m�dy�	$�GcϤ�^K�p����H��j{���"W�9�T��	$�;^�iz�y���Birz�#'b���|�52�ϒA#���sʙ%�� �y�%�n�Bx��������W�f���)Eon��M"9�u��s�x���w,�� �r�nY��Z�5�7��5��d��^EL�iAv�1Wv��� ȫ"HH��� "�������}�!%�����K\��T��y�I%O�@�ON�K�E3]Ғ��*|�I%Q��%���ΑhLh�a���'�5h����9d%f�K����Cu�tf@��%E!p��\ff���z7�.���"�7p�y晐� �H�^��RI ��&|�����=���2�aRH$�~�y�9��j!y��`ʨ����%:�J� �`u8su�(H$�I���BH${#�L��KgEV�|#�{�D��S �����9
�V��2�H��"L��dyޑM��ۜ#7X�$�I=v<�($�쎑2�f�}�fL�˦L�UAv�\�[��7m��;�O"_����J�zD�D�6u�We����j[Ƃ4}��$Q7/w��b���g�;�������^I%Sͱ,�r������AgMV� �g�e$�W�� �dl���H�<�c����2�=�9"޳(3��g;���G��.�n�\8�3|0�=������y�؏n*/b�$�щ�L�����ڹ4g��R@FDD$IA�G����yyrֱ{��n7nV��z��4ce�8:��޺��")t��5n��sH�4�*f��p��܎���1��b'5��Ѵ�<Ml+�O�F[���"lЅu�eu��0�b�2�E���z�6󻢝��O=6w<���=�A��nl�7Xg�v��km8L(���e���\��$�a�a�c��nR�	����D����n)[��9NA���ƞS�gr�e�n3d���У�H�����~��p���59/"R	 �tl��+�_�c/��"zS՛	[�?z��H�L��3�R��O�;����%䵴�JVC���)�Iz�:Dϒ$����D�S�����hMc�E����GZA)ܸeUA'��A$��ȟ2I���]5SC^.)��H$����A2]8�(�v:0���v.9T���|��rH�A�E�ũ/���|d��ɷ�R�I�;^�8�j%�v���m$��dO�.�d�m�3;�%ܳ5ݫ�k�M�޷c��j�
jl�r;Y�䗦#$L�%����R�)-�ǟJm曅MyZ�{���W�,GVa��	n:�t�����\Ym��*�b�7����$�;N1p�?���,�ؓ($��N7D�2J�����=/$�4s�ʌj-�6Λ�2�ə-�~�Md��E��(1r�D璊�y�����ޗ-�#�����^wr�:_tb���٪���Y���c�O�q�o{�	צ�ȷ��PNqQl��ۛ8Φ7#C���g%��W�o���9k�ݾ|"�0���2��Ȥ�;���Y����un≔��]?c̢��b$��Ά�4�^i9^X��,K�D�^����2I��x$�K`����qo$�-�0d��o��^��K�1�R��(�!;���$��b���f�ɢ�$�mƘ�I$�U9�3�IywlQ�̚��S>��פ�h׹D�Pk���8^uި��z�e�V�*^_Ƿq�r6]ܝ��U��
@Iy$��y�W�D�m<�J33l=��w��+?��v�[�(F�I�9����(eq��P定�GhJq`E�=���v0\Z���s�s>d�I#S|�g����y����C�O�0�$�A,�Ǒ)^iy�I�_ɥ�y"�7>�A*��Yُp���AT��Y�`����e�DI��P��Z^+�c[�$��BB)k�%.SP�J*5�JA$�s�甒H�k�zs��F�(D��i��^��ax��ǻ������k�j�U�D9�s��G7^=�TQ�vۘ��6֬� f�1,bc��Ǝ빫n�Cz��~
?"�ȡ �"2
��Ȣ��3[*�'��y����Iw�:�JA1���w)�tY�j���3�U�K��a=��ӿ�?�����BI%�Ҥ��UV��^w5$�l�Ȕ�D�n�,�N��*�I��e��]��l�5ITסq��Q��2I%\��D��Cr�J+z�I7�'�?'�_3Kꆖ�N�2Z�t5��,T�e�օ�1`�M]�j$Bhb����\W�u��V���I$��NHi%$��?J&�.l}Mw��{_y�&��d����)G�+[	3�D��f��ӭr���!��mT��3<�(�y\�A2���S��Wst��2��1S�׽)xDM��9A���?�z��H�B7�I;:r��<����L��峭2�+r�HIVT��MŁA���*�QQ�:wm�>mS�?�	g���-$I���N��%� �M������~f����8I����&%�^�ܣ���L���,���6�zE����F�%m6�Ԯn�fڲ]�/��y20�S,��=m���V���<y�m�s��3\�(�"��"H �,������(�����UEU���9�k���O�ئA�$��	���e�$��q��n���K�i�R@$���T��D�_<�J�z֝�Z��@�kr����$�8�خ�C�4"���h��j�]hK�iE���|�d��7��p�H���$�����I-��of�jػ��N��2\��*|��5��'b�����f�̤�]@tGBvn�Rcw3�/��2	t[l)	 �;��M�f�t�j�ݽ�y��g�[d��$����v�"I8H���擅$���P��`�+�}�+�3%я��RA*��>��	w	�_���$z.�bب;�Ϸ8$N�5�3�Gb���$]ӯr�`�Y���K�:�*|��t�HmH�MB��EF��K� �.���"a�VkFw��d��or�$�*��z��m(������a���8i��ӧ�8p�ӗ.]Q�J��mg�4_��;�|���)�=�:��@n���]=_6`��ߝ���<	�]�NL�KW���i����x��{��݅xh���<>Qe��z�ڽ�E6ͣs�ݏd�α)؈�v�EŞ�r���� c�\��KxM7:2%�\w)v�pz篹{7��W�YT;�}��_{S�ܘ��=G��U�6�[���){}�w����s����m|��M�^L���ϜǦ9'�����G����<3<�󹾾9Poz��8�{V����c�� ��g?>�/g�Ө�)j=��٣�.:;�^[��hz��x[����%�ӹ6/�{{���T��D�C����])�no��Ta�<���t>ި���{�@U��ܳ���d`@G� ��Rkk٫l?8D+.wY�֞xe;����_n��A�S��TBw�S%�6U��!{o�2�v��#G���W>��	��e��y����1S��1�����*��R����&n�T����@��@;�L/9���y^�(_3ݏz�(K��ӛ�������]����Rn�7սd�S���scy�{"���f>�O.RiT����9�5�q��"þN�TP;_c᝜B����~yzƳ���%����g�
��{�{tw	��2)SK�ޗƥ����NdH]����6z���e�����|l��p9�=}7w�Mctc�4�zrC�B�En�Zǉc�	���=]l�^De՘Lw+��6�K�9�F|5��.ℜ�c���d��E��u����ၥ
x��'�$��:�!v���7@KJ}�?ǣ�҂��+�ӔQ�+
�Y|�r9Ts�R�b((��,��,��@օA+Mwun���IU����.ロ)
�%lr��t�x�,�P�.$�eC��)����L�����
J��.���ʎ��΅�5J/�7t�{��\�Oy��8���6��&�$�"*�R� ��3�)�]H.���ă����Q�T�"Y�Q�ne\�JvaU+��F��AȹV�3��@zkI
�3lX�iec����DV�R�p�s�	�F���aTR�9J
��� ����sI%�iENX��"*�Q�(H���'=�6UB��70��m%�=i*�AIЊ.�%���%����~JK44]����;n�����v�n��=v���Uq���N�̽���]G\���˞��sݶ'�ݎ�ɺyI�ע����rͺ���r�{e�g�7�Y�d9���^�ѷ���ݵ���ܸ���r�fO���yK�53eҬ<�ۙk�u��n��.��35j+A�V!�]ۂ+pֻ
��Y��v19� �'���,� �O9㛻4Ak`э�bY��EЯ�˪:�ԕ�F��9��kz�l+GX�t��aD��,�TfZe��!mL��G5aM5�eo5Զ��9.	F��]��זrN������c�9p��,�.%etf5p�]����EY��p�H����V4��й��fc�FB��M���lD�����J�v�v�{Kɐ�@{N��`�.�K�ACL��Ҏ��c�b�1��Rʋ0��#1u��4e�����u�ͅ��(r�zL���\@�MB����fyC1<��7ld�մİ�X�Ʌ岔�ll����ѧe�o򌷈Lm�8{�s�6gT��'3$�M].�Wl�#���1�J��,t���.;X�P�8ps�\
�������C#�*+Ќ�i]	H�3ڕ��F�v�^˳��R��ngQe�-sD��[+�]i+u!W.%�1\�t��S�X���ge�dIF5����;]��kv�S˹�EF�ZhƱѵ�jج�+v�T�SQ���J�3]�e&��%SMP�=�b�+:�mˏ(hK"�P�hۨ�b�7#�n�� ��s��/P�,��o":��m���p�h���k�Ű�Յ����&)�K����j��ѷR�nr�Uݣ�!62��'P���y�+����Dn�F�5�
�G�l$��/�}��7�|t��HNBI������Q&��ۋ���u|��N����Ѯ�����Ÿ�&�ڞ��z���v�\����s��V���s6�5��m�^j{����w=�c~�ˀ����v��0�0y�~?���^��Y�!�t�[��)��s �^��b�cO&	\�����幫Ӟ�=9b�t\aV�F�tG���k����^F��n�[�5.�&��Vj�k����"��j֪�Bf[�*��7u�i��fl6�<l"�қB�KF�����Du�%5i`�U�]k.&td�"�x�h����\i�ze��Gh�+y5����bDt�2���L\ᖒ�m͔X�m�i1�����������+�Bhƹ�Kʼ���I$\��K��S㵬����D�H%Q��%#�$�S7�ܸeSI:��)-w�k���sQ���1��LR^Iysμ�!$��5A$�BB��˺�6.y�kV���-��I�;9(���N�̠	�%�/�	%Ouq�b#Y�<vF�H�ܞy�	�}3)��+p��D�pɪ�.�W$l#���g0�	�ǙD�$�Oq�I�$������NU7Gfj3y��q�JY����3�K�<��W�����2�:Ή��mǑj��t��I/*{�3�E$����ғ�G�a��E��lѸ�wc���=���K���Ʊ�u��/��&b[����"ɖ��r70�!��K�S��)$��:\�3&JA��͘N���H䍿l	�̹�wtID�1�3�K�{�4��vj(<�k�6e'�tV{��w;{�OyN�$�ov�:\�e��f�ǎ����v�gr|C����s3��6f��������Q���	��	 �H���o?-�5T�Kß>��2A%�3�yI��41��f��ܖ�J@`�ز�����*�'����\_2'АJ��O@�W4�YP��~U�E�hΑ J(�����z�ͷE�;8("��6�ml��9��/%5��	���(�I.ǞI���mʠ��^ٯ$���$ϥ$�]��.���*֜��2IU��y�R��d�w	�����%��Fdy"P�v^@I$�c�)�𥥹ju��#�i�����e&��8�xyWs{�L�t��c�Yh��M�t(�8:f�G��þw	�_��tpK2���W�y�����I$/�yL��geXk���L�)���*�RKe���%�ْ�$͈$�MB�K�r�"<�w�r�2��;����z�($��B���`37����z�>�W�Yǣ&��ս�sҐ	ˌb��tIL���,d�K���I ���ބ�̓�9�UHf�hߕCBn�V����g�|6��kn�b]=�'ܳ$����$K�r�|gbl��mnٶk��O��B@DD��E>��=������_�JD��~Pf�H'����p�UW�y����\k̝wFT���ؖD�^�y���I�����J"����O<�
R�F�79I��hs��K�I���n΅M��R@\���I��������M"��N県p�ݙ����4p�xu�պW�=�� ��f��ռ��n��ڋk�ߵ�C3yزNl�Y��2��Um:�	H�1-���d$��*��$E�S1&RA#�ӊe!xl��'pI'���)�T�����
!�s&^1"I^�y�2L��]9g�[�gd:3VnGEö���+�6�ޙ)2L؂A�t�*��޹H�I�q�@R�%��̍�;33I$�ƍPN$��G��4ܝp\�NR�M�:ӕ����v#4$��k�2�H�:v0�$�FtI#�PM����k����y�� M�!������~R��y�]No�w�\��_K��w�� ѷ��~[e��5�Y<�g��íퟂ� H�(H��0�;j�RX��������R��hR���U�����[o�:0Iy��T�I$�r8ȔI��x2��
�ڔ^_k?{f�k���v��X�&j6緩�,�K7`kq�n';B��<�������ջ`a_'��<�^1O� �	t��;���;1&R���~s-�fh�`*��S(�$zu�ϥ,�]�37��vb�UR�y��M�.��4�m�<�I .v4�2�I��L������MQ�ٰh	I�Z����$����Kr��O��3�	�A*k������qV�6�v|�	%sѦeK��9�&RW�%&I7�r5
�)z�7�-6�GW0�&��׶�b��A%�ؓ!$�]�Sۘ�.�"���Id�q�I9q��8g��)���>	%~d{i�ЕF�T�L)֤�%{�"L�I ��މ3��	/.Ɏ3)�C�xxW3cC���.�[	����t�wu���e;��i�-�z20�A�G%����9÷7*�7Q�VPn�ƭ>�rݕb�5z�{��	E|O�VDd�E$ddC���ު���+Z��ȍ4t�X6gr�aqv��s��nH��\[���T�ԯ[C��m�Z�FZ�q6�,	.ً�ˋ��C)�Q �����H��J9�4n-�کǶ��ˢ���Y�`#���'hv.Q��#��;�a*��R&��Й�r�����&�!Y��֔�;#.����ewPԍʳ��.����T�;Q�]\WM���6/��q�Ϝi��<�툦�2嗙\��2�\��֒�S����d�g��%�.~���x��IC3{r��ϒ<^��9W�����(���7�L�$��$�F3733'wrX��<��,����q,�=z#��8w��%��!$K�vLq�U���މ�e�8l�֊��O-�1�3>���v�) ��̮���PI% @��gD�:RI\,v�@e�7�[�J�ܙ��L �ϲ��?��D���L?�fq,�i��I���2��2AmGH1f1q6�Ɖ�0�M�
Rމ	2K%�.�|&�R�d	D��NtH2ِ�Ic3'Y�`$�m?J&G�Kv���Ey$�t���gq��2�Hk,NW�c)E��h�Y�Hdː#n]vZ=D�3���D�îY�9.�S����	N�Rw[�H$���ޑ$�-����ç'��۷t���5��`�j ��d�g�ݥ5�ey"=y��Py�Z몌<`=G��x�C���z`�Z�ڧ�5�<�wA��?k^���n�{������Om*���| ^���	L} �E�D�B@ E$��E�Y��W���
��*����D�|H�Ϡ@'�禃oonVCem:�Y�����,	i���B�9� �{ Nu[fŽ��꬟H>���NE����;�b�#����Y|D^��D��L�I����F�OKQ�=(�fB���*�0)��d��ɍ!�3:%�	�}�-&�$�'�N�up�)��X��5�Tω$\k�	��l�T�g�L44�o���������e4���ule���o�KJ�m-��[W�-��:�+�H����-�E�e�p5/Y2�G6�$x�v�tϋDLV����]g��&|q����5$��g�3'䳆N��<�`�僠e쨎���A��� �y�:gĂ�6��z�d_T��	(�H3;�d3�u�s�dH'Ă<l��N�PǪ:�Ɯ��wL��cb�y����gw�
��3�z��s��>jS˥��P���l�<u��1<R�S�X�Lԣv�>HH�"Ă���+���"���y�$���`@��>�$X����ݓ;;"���*��ܵ�̗����,3m�	$k���'Ė��[XӲRM:얃'���`�$������Q��f(^w��&]���ċ�}0H:��I ��lW_�����|�e�ǲX�^�,)Ե��.l�M%Ε�*����F4��.��O�^���m-љ~��i�"��؟?�1��bJ��9�ץ,Q�o+n4A���ǠS��+�]<�5]s2AS���A9j�c\�"I���A�{fAs	�d)w�^k�a�0�3��'e+�f,��k��-��P�y������"Cmt�Ї�=$f`������]�Y����#��&�I��w'�9�� S��#o���0;a:���Y΋�?ye�ǁI9#w�#�{�eX=��)�-Ր m7&r����}�^��/ps��^�@���T�W���T�@� �$�$�a	��g�5���rH|��7Ν3��	hF'7�	�1ൻ��Zԡ�x'�ļ�l��$��7�>��q9[uK��\� q�朂Y2wd����:���=��LFmP��]�aͺ��n	N,�����̜3�-�7�y��D�	�� P�ܳ��k�d�M4�L�yD�y�38NR	�A�q ��	4�&�v}ƽ��$�Hӹ2y"y�`G�O�%�jm�V��0h���%�^r��H��fO���x$��[]���}Z����I7/{2���?�7F���ೳM��T��i]�!u�'�G��/7dI��n�O��v��Y(�z�9��Dى�&�?���fwp鑉��Hϒ�ؒ��Sr��9p	�Mt���G5�%��c�(�����/3B��P�)�\A�B<�힌A:ޘ��,�+'k[����SRN��))Y[���M�X�5Pm�uY3<��6�P�|�ǈ��G�F���M��w�:h�	�0����$�� !�9�q�1�����߉�qx�T&�8]��{/8npnM�(t�aP�nHLt��x&��h�6���%kU�!��v�B����*ڳ	e�;y%CZM�773�'9x�&���{n�T�-�Q��L��.�+���6�tm5���j�0Y���2ܚ8����skJͻ��4sv-����w]>�z�@\6��e�up�Цn����Ԏ�gxӀ�y�ґ���
K:�v]\k�˓V#
��
�Z��cqbA��+��E��Ē�c��|׏ �I�~ɟ|�]�Ѯ������1�%x�}���Tb�e��2pΜ�z��.fI�"�d��W7`Is_@�I��2H+{i7R1�N��Vjȋ�����p��Ȕ���I ��� ��M[�7M�[[dkv@�rIf'�z�A>���%�^r��I����9X��x���� �#��e랸kn��'č��ܐ�ùd�[gjd�	)�g�dUj��Б>����}���> ���0�l���i�;͵���x�A&�@�q;�7F�"�6�3aa��.�����T&���|����;�I��/;��|�ddĂI�>�~ِve^�D�=�8��z��7Dlω��=-��3�!U��gJ���%�����H�Vzc�����wA���Ov�P����ߪ[���rC�Y�V*X�g�bêL��|@�Ā $ !��s�2|���&df>c�'׻�%F�s:�kO�1X��H�t]�i��ۙ$��$y;k��i�{�.NTOp��k�:d�I���@��v���8%�;d���0���lTO�� �b�r$�v;`{�ܪ�`��KuVH�P8�0K\"���ȓ:�r$�� ܾ�w�?M׉~y��o�~� �v��t�1Ӌ�{�����ř�K7K���%䋰�Xl39�9t�S�헆�n{�p(h���L�wvft��5T�� �s�$�H��&7�D,d-�e\� �۞�	 ^a�S.�;;9)ɻ��N�/Mz��6o�Zq�;�O��rd��ͦ<O�D)�k,��|N<�-n�3�+9'y�{9��ݹM�>c���o_8p�ç.]���I�W���5��Kۤn.~Я�Y]R��AOk7���٢E��8z�w�����Μ�f��}���.i�ny�s�}�A]9ݨT�d�+!�K
�=N;���n����X2���K�� {G4���O�87ݹ�"\�y�C^:=�:?{�z�Uꮿc="�j�`^�����3�rz��=�s��,؛[oC�yxό���U��k�k����j-�w�~O"׮��㋽���}����l���q�-OS�� ��w�g��U.��մg�\?���_�{ͦ�s˯t疉�����-��Z%�Bl�M���Id̧˻�ӘP3h�����cڿL3Oo5��sԖ�|O�-C�|o }��pQ�`��ק��m0��ay_,�{�V̼�y�s�l�==�z�Rz�<E�;�igg{v�*l'{}=�&{svE�</���랞��;�Y�s~ٜ�(&#�<��<�z�=� ���^^�D^yJ�t��j�h�@;���o۱Q��8e�+qR�5���%�g�m�呴��:�x%_�9==�~��~Ký�]�
5�m�3ò��i^��i	佨tr�T�����y���ץ�{v�N�&<��W����އnq�'	��{�qg���qbԼ2/.U��C��"V��!6o��6��Zrٻ��΃�5\���r�X��?�߳�M���ʂ��}j�d����m�#F{v%7ݽbQ\���.��l�����{����z���{\���S�}�e~L瓋��W�o]�̥�c�)g"9�=ts��M�M��2L����#����,�X��(���EĬ+d�a��8��:���t����t��I�U���r�ar����^�s�+Xe�����"G�<����%��Aމ\��2d_W�ݚ�B�����W]�#Ͻ��r�瓔-X�U�t99�J�X�*nbXA�'�'W�Hq��I j�i���Y�r���d��.e���%�r2��QD�e}�ty��
��eU�/[���b<�o(2��
���)ΥUq6T\���(�!K����klx���jV�^!�XV*��ۙ���������
${�:l�����N��Y�\�UUrD1z�+S"u���z<
�:��#��"R΂�A�_�o�Ȇ�ߵ�e{�	������L|�1�E��!� �?VԚ�=i���G���|�I�[�O��|�-ð�=�@�6�R$�6	��;&frB	�v�E�	u�|k�fV�h��H�홒@&�T|;_:d�E�)����&L\p��n=l.r�os�u��+�]�Ix��=�R��?�����g���~�-�s$�]�}��� ��)�`a����N���\*�~%�A��v)�:r�A���@'��U�0݇����w�I>�m��Ι#zJ��\�m��o���נ�y��9)ə/+6<ē���$��g5YU��ݠj���A#}qj�rE��p�`����i�E��9>=j����oL�nG8��~�;�Q1V��y����S;��3�8������ ~�<�V�8d���S*��bI�z\l
wg��j�y$���$a�M&�������|5۩@%��k���!� 媇�]s �|~�Ȇ]��`�L����~G�M�����mw��<��".0�z��M�T�3�N�ru�v�2v^{7���W�J����W\58@�ߏ��>�^gdS;�?w�Z�o@r�$�{ ��}���q̥.�-��HWْ/Lܙ݋�˧�$�=G��vү��m��X�O�6�D��۝Ğ1C�� #[���>���o:)�:r�M5;3�A �g<J����b�l�0�B�I���H-�� g���Kw�ܻ�����6���7,N'X�z#r'�K��@$�v�WQ<��!ۢ4��J�����0S �g@�I�Wjm�]��lH[7� ���= �u��`d�1b0��p_���ʬ�=J+��[����S�s{Ϗb�m�y�P�0���0%�Yz����"j޻]���?�n5�ks�~V���%���|�o�i>��R�B�Y�ta�vk%���M�3�{j&��m^��hLv�c�v�|��e�[�NN9�4�a��!���msv휀�/Oy��2-��[S���nyz빎���Ns��7��1�vz��l��wZM<��a��gmjvi鋮`�ˋ���t�y��Qx.��:ܵ���L�V��-�j6:�Mo�׳+�ձhx��\���7p'k�v��������Ʊ�]s��&��3WpV��2p�w�����:d����˹� ��@��I�l���Kjf�Za����|�� ��@�y@��;"�؆E�@$r&<�l�ݻN�P��H$���H|��0�{#�dsA�R�B�ۑ!�S��OB���@ �}�O�c�c*��Z�ߦ]d�oI$��؀Aor[� �g�Gi�[Βw��P������I{{��������z	>$b��uwD��C�f�|�Iv���=����v'�氂�ב>/QT��G��g��>+�>�H-��T��BWlU������Tpn�Bct]�pۛu��cVEúS[v���� �Kv�%��L�rK�ޯ����{�K�'��1�3�t업�6�r�q$�|����bQ,]2Z.���|@Uվnv~�U�C����g1w�@�J6�Rg��ʲT���#��`�A ���Y��������[9�{�"�$�Cp�ٓN!��d��@{G��牟��	�6����>�d��6��w�>�wX9�NȦv!�zq�����Zk�$�&�E���^�"�n��ٛ�&�yk������ȓ\��V��	�ӗ�'Ķ�l� ��v36���	���w���`:p�Ŧe�vd�O�Fs�a-͛ǡy�'E4 CV�D�H=��=�k����N�;�NX3��vs���]��;B��觬tj,������/[�H��|�o�v�Jˆ l�ȒG��ODx��v��x:�Xfd7Bo =U�ω�ĥM��ȆrK�2r'����\��SN����|CUnD���zy�)nx�5���}��ؼ�Ȼ;VV�@�O���A!�G�L��Jv��h�>[�
�]���~�ќ����aK7�_X���_�h��m�`�t�a\环�s��{�Ӣ��2������P�v�A������y�$>ߢ|H$�ӑ2��N�gD2/#�<5&�x� ��!�'��EtI�VOD~H�6���j�'�K[e���"A ^D"�8L���.�D���=��̭�i��U�9��?L	��OG�	-�����.S�a�t�t���'d�"�M��ֺ�6;5������6%�����-�z�����`3�fb��^7f@$�\��$���E`��j����p�4�gLߩ	�ݭ�Af��_�݂vdĭ�c�h�J�5:��uս	���ȀI#���x�lX7{��T��7u�	\I;&��D3�\+�jgc�'����b	=7k&��l�mdL�OQ �Ftz<GKo(�$c5��YȻ;@��Y7:�%\��>���|H'e��x�[��x� �Ӧ<�i�w3%�ݥ�9Fff�%w�{a����~��m^�^7��|}���s��/_M����޽�=������Ͻ�{�� ���� �!'E��,�Ń�(�c�z����eU��b�ʘ�I7:�`�[7�sU�|���<���$ˊ��M�P�������RR��b�3\�tYy#�[V��`Y�?��~Ue@xD�nm�A ����c�VےӰf�5�����ȋ���8fdZdK�T��i���s	8�cĂ|ݽ� �ۛM���
���"	,��w`��Hx��\C��� �r��-y*���ѰH$l��yI>/��
�q�bf��"�.W�d�<��wl���Q-�� ��^ȐH+���q��rO	����c|�v��6dC"�v�T�+�I �
��oM����M�����CWfD�I>+s����fE�g
�x=o��f%��d�?`l�~�Ec(�� �0z��~�%�?�v��B��ˠ�ٻ��Q�t]"��_`�e�Ƽ�<��L ����fy�����4�vZ�\P�v�g BŽ)�6��Z9�д�$�gZ�qJu��{>ס�1��ی]v鹷T�8�quF7�r��u���6��ݻ,�F�`��Rb%��,4�W]����t��w5����%$4�4�5ʻ$ں1�3sŎ�K0�Ŗ6�"73��,��Nɸn�
FHLӕ��z�ڱ�urٳQmx�^�W87.z���;Zֺ����{s�8A4�:	&Sxo�tɜ��9��Ai�ȐI�[: ͓�$if�ӓ���S�Az���	-t9g�O[�'��iY;Ͱ��i	n�ْA �gG�5����tLܛ'C�	L����f)�1�bɯ$SgG���,�w Śu���`�$��Κ���v�fY����]�L�ͳǈ�B�(rL��ĂI'��� �η�����M��@�K4z݉ rfxK"�N�xΈuv��ӑs�$eGVT̒	�"�>A�Z9
�"�b��}����C��=U��"��;tS�Mi�����!�Ƭ6,�dم�&8�#�׿�J��'C�sU����I~́ ���0=_gJ����u3�d���x���✲g�^d����7�ֻb[�Ъ��Um��{v�6�M�zȤ	˖:�=��F�ö�>ѩ�|���{��	@7Q�DM�e#�{�3<lp'ĂC�lA>d��>P�$i�@44���ˮ;�"���y�9t�$޽D|e��$��M"�y߶fsI$��ǣ��9A/b/&�fp��j�~�����k��A��� �A�V��$�}���~�\��{Y��!��!��dI������i�bWl1 �-��%8�}��P6-h��� ��ۊ �sgt�<�r�������$���D���E�ڗM1ΰ�f�z�m]lXu7]���3H��9������+�S��b:�<O�:�PA��oL���U��O���*N;^�$Luht�`ř��*��0x�^L(C���3{6"�A� �)ڹ@$9�z@�L7OH�XWR�>݌�}@���L���ĝ�2�k��� ����xkƪ�S��&�b7g�������
#F��7td��֚Y\�������ݨI���t�k�Av�� ��$<�y�|v#�xEf}c��;�PH:���$�Y�w`�0N�y�����ڕZ�6�Yu�`A!_v̂E�����wS	,�cQ�(���PMp~�I����I0j�x��	'ƣv!���b�-(�RY�A� �n��O�5��0a���5O� ���~�}ɵ���x�H"���nй�t��b��-�Ĺ\j��C	������ś�����n�xĮ�b	OnD�|I=�j�f;X��cg($���2��Үt�`��p�E�� �݂K[We˭�A���7�=;� ���x��j�\��u$���gI0fL��3�}�$OFdA$�4��D����|r�w1f�ĂI;��e���3�R/D���{�53�`e��$�I��x�s�uy�����.1?�҆{u7�r&���ז�O�*>>� �sigM�}�����a�r��E�⇸|x��]�~~$�ن�i�I�cpX��!5�jx�{�fv��߳�s��&%�w-B�c�ǈ�_ty��>o?*�}w��p'��fI�'���x�� ����)��֒J	?�;�Ń8ww��cx��du\�u6���öy�kn��oRZ���߯g��E�9tX.�K�d� ��؂I s���o�h����Ȫ�}�� A�1ŵ�d���y���0�X��{�*:�q��A#�z y��A�1�*�$�v�ɤ�7�;2L\4O���$�ήᏉ�3c��3ٯ}��99�:��g+�E�,��h����DG8��Ӧ��A��H#q�H�n� �Z�zqt	m�s��)9� ���� ���N䔋ăآTZ��$��(v>_0���0��� �7j�Ij�蓞����x��nǯ^>xݻv�ܾ�͚1�j��o�#s߰�A<��Og��7����.wj���Eo���-�ɦZ����j��-�[�^h��\]���=��`�\~m�6n��{ ��s����K|'��a�1�xvw/�=�:Ϻ��~�h����~~�=�^ܱޛ������۞���*��;�v��fIj���

&d�ؙ#�	G,�Y��@!�<K���1���>��IƯ�6a�����/�)�̀��WK�c�\�s�����zR��}�����b=���&jŜ��1�D����;¬��Ò�f�4}|m��k���5直�)\�N㷻Y�b�l.�����P�K;$��C�6���T�o�ť�������������׊�w׏fz��9�}<��K����o��z����d:��*G���Ň{-�s�}�ݭ�_I%����p�=��|�>����y��ՋN�a�gn��Y3���G�,��E�僻��}����jIp}KZ7m�Rwrl��+W���<�����z������4���v;zj}Ay3Fs��y��=�]���	���$�����y�m$�B�������w��j�����G&��ME8I^��b���X�:��˨v��<��Z�<x}��5�t�7�_M�J����󃷽Qc֣��Xݢa����v8�{:r~����j|���y�4�X�����'ފ7���kP�彳X�}Ў��� �E��Էq�����M��u��/�#�����f�1}BQ㻯ẗ�c4h ��@�IG�=z�����7��ŗ��|
��#l��O�]^nXJ빁	F�0� ��M��Y�K�y.m;�z��C�eOu�*�놆R�]$NQnl2H��C�uJq	l��u�/��(�]���l�VRW�!Jr,ĕ�0�@�7���Fv�f��=�uJ���ED^)��n�
#I(�"��T�z����X���R=i�'>����9E�AEp�GW2������k�	��� ꕜ�v�z,�4����U�pL��#�k���=�ʢλ��fV�d=�S�!I=ڙ�iBA�"�KF9�św$�O�̫24z�#2�W��Q�D����ty��oq
�ގW"�=��(*�M�y�����Ew$)������"׸�\��{�<�Ȫa$#�Vߩ�?��,�>����\��:ݳmd=��Dn[�poA�]��Ŏ�R�h�f06�^�u�n���n�&e�d֪�Iv�&��Ԭ;:j8Nyvn,�37���Μ�tȏ`w\�q��s��(�36�3X�J�in���-�l�Y��Ð%�:�lB��eMu�b8��lE%�ڪ�r�R��Qζ<��Mׇ�hm��tVl�l�R0�\�\���5�Z:=�%�j�5�Ĩ�'�*nD�E��m�^��d�fٹ�Wk�i�Ba�X�۞/ll�f3a[�v���dy��ۅ�m�Hv��R�sخh�
���G<P�YE�;\̉SYW����m{<�Ź�:���G�=�d�cfeW��5���C�˜4'��[Z�[�]z��8��[��<��r]u�p����af�ܬ����hHL��v"�\�=��&n��t�jC�X���}v;c�Z��Fh�����ı����fX�u��0���Lۉ�Ii�rY��p�L�k,�k�xmó{6�[�5��n��;�^;Xfϛ�|�n��`+ln]m�k,�:��,���6��Im��қ����j:b6��c��^�;n��(]r1�cM�v��Wd��FW��Zpۓ�f�Y����I�f�Z��p]�Kq�:��S"l�����s��Sjԝ��K�2�s��fF�)�F��9M�w�0C�fa���L��B2�B]�-��hSnY�5�ᅛb"X�۶�i#��B��,&ڬe@����J��9�q��2�3�+m"Y*�]k��`��n���kQЊ�[eE;VN��GU����y�{�p�3�Ig���
Gi����Լ�%6̥ek��]f�{N�P�$n����Adݨ�|���q�ny�c������l��{���m�c*ݹ�Ν��mvaN�@J�^�Eؼ��F�GV�es3�\d/�J�F	4N�(�ݙ�#Ϣׅ�g/X����!GC���k�ֺ{f��ʽsi���{�Hs�ڇFx<��.f�%�93�k�ySN�g����c�F�qS��Q6�<�zm�^ܭal+�]h��n;<e�R]u5�3j����=���T�Wp/D�������h2��XY�Yb-��i���Mtc�J���7{��_C��ZU�'��\�����Z�s�f��ٌx+y�	�,�2�5`D]�^�ֻv�L�/pճ��r�g�m�x��P�	$i��q̙�\Yn�'��iݝl���������C1p�|?<q��	>agCWoL�n�{�<0_C�_�B����07�v�ȗ��%k���������I�j� ?���G�D�wV����L[�N�]��o�L��ё�$��uԍ	h͍L�KMl�@��Պ��n��54�����I�����[�"�C<^�T�WtH��ӝԭmh�s��׈�B6r�1t\"��f��ٹ�	�'�2 ��I?NX��$�4ݪ<Ak�ْH��x�8��g��Șs1��*jfr�vlۘ8�k��nxܥ�^�w6M�E1d$�˗Z�2>N�ud�x�%��,����$�f�	l��\]�Xc��g�eШ�vfH�郐�\b�0�Q p�p6�l��yti�'��nJ��=��3pxW��o��X���ww�����!��P�r�{��Qܞ�Q���DU��s�"��~ ��S�� �[﷦A �z~���.w��9�� �.L�o"��(U�2g�_�����x�˝@�cI'���r�@$�5�tω�'{nw�%���w!�LJޝ:�vu^�3z�$�|Hyq���˺j3��FK=�|hn���-�JCqg.�r��>��z���̻��o#��n�̒	=}����B�P	��x@̓o7���&?]�\��<�Yʑ��hz��F�+�hJ�h��#5t$2frȱm��b�D38b��uNL���c�$l6��c�S٪��I�� �j'��8ggE�M2b�� ���w&���6�%�"�$ݷ�A�m���@���=*k�N��Us��b�;�@�N�fl$���m��w=Û�i��35mI�U�h衔%yP�w7#=�_n�)-����d���,���@hh�x!ػ3�Y|�"l��>�����}@�I���@^K�m�.!cX��ܖ
dK�\�������mM�tA$�׈G�i��VboiଛD�{.������!�g+��w�'�Dv�R��	qq�}0��	%�;�|e�X�/۾����a2��&؀��ۭqK�\p]v5�]<�;��Q7+�wo���~v���ne�c2��I<��A ��tIlj��z�C3ų�� nݛ'�>'�鮽r�	�?�f��dWL�|���,�-�%�\u����H&��HU�� �~��ǻ΅�\s\���r�S�����>9jfodI���wD�ڪz��$n��	��&�D� �.b�$ʊffm��j�$u�|H*�z$H;=�=40;"(�^g�R����	�L���Ɉ���妹i�4�͛X.Á<��اZt`�9��ҩ�9��;B��x�
s�X���u�<>��>Z�Q�o��.�����L���vU	�����&*hnu�=4����=��2'�:"Оνq,ޯ��̰=��@�gYnl���>T�/-aϭp�ͻ6�k�E��i_ϡ����i����Ī�bc�.����[�97M�69TaP�
/�˜�R�8dYpwN�;�|크,k2�`b6�Ѭ�G_FL�H=Y���6Ҧ��=���Վ\��33��i��ج�IY� ��g��3n��[�_�/)ܞ�$�����v��Ȼ�wd�d�Ȝ�F��׋w���z.�G���svǣܟ��'Z��;e�ES�P$vG\��0NXv�(;�C��<�Q���n��5E��^m�ɒA'��= ��ƃ�X���ɺ��ff3����h��KY�;�L�h�2儴����Ƚ�z�L=�v�y������� ��h���mk1�ԉ�ż
,C~M�����;K,�I���%���!A�j�0ٙ]2�b#\e*.s�Ɓ��U_6����2�[(��6��q�f:���x�ym���ٺ�hܲ�=׍�
y����h��l�y�#����h�5�H6`j;3#t�Q#M/ku���)j�]k�㞦<��GP�\c��Zٌ��iɖ�X������Gq5��Nŋn�s�nd�q�7h4��8N.�6���vUKx��w��}��(9g���n�A7䁼΁�^<Z���k}Y�Ätn����+�Aڼ�אO�H.�,�<��4��ջ�7��Ѥ�ʼ�F��h��(Ķl���Г3Vi#j�X2�.K�.���A�><Z��)�r���.ݯ���(���L�x�kA>پ�wH���C$�*��&^�)2�ec4{n�	>$jkƃ�A|��Ch�SKN��2��|�!�M�V�8� ��zc����}��ȏ�K=�A�/*ן�'{�Ϥ�*X��ܚX�M�L�s�ˍ���'cv���y�D	WgP��S���>~��y�!ۇ�P�H4[:�Mf�L���|�UZ����cq����Z	�/�]1d��pX)�޻��'ޜ��(䨘1�i3��I^@s
ڐ9t�Mճ�_@�߶\z�8��]��6́�6��R�2�wZ`�xܻއ���c�񿡧��,c]P�����������r�H��>��,Y�W8ݖ�4A�pH�;�.Y�y��c�@$��tI$�z���k���Ηl΂��v�Q�I]"EI� �X�rY�;L���|�,�cR��o�I=W2O�'��ng�w#���DC?($F�s�A;g	�2��}TH$�ȍ��S�Ve�b�I"o��A&��]]60+�z��]����2.�r�<Lܬ/)q[t�-��t]�s���9�5�P�eh�Ek���w<�Ⱥt�7q�Q0�ױ� �I>�� �a:3��y���A"�#�A7�k�HA��H+��	���8sOea�wA��#�|H$���-V�r6u5;�4�t�t̑.��`�y��o�'ֱ_G���������ZL���Ue��D�"b�v�Ӌ�V�Lɗ%��S�_�Q�^�$�z�ǐ��4},��h|�����)&�=�����R	��t� �}_DM�D�!ӂ圇�4���V��y�+��;vtI Od�A��4љ���;7�MA� �X�p]�u2D��|$���y��q��5�"���}�9S��"֜q���Q�Q\4�oSɝ�L�S:�,K� 
��g�x]vK�\i����{]@ufֳB鄔,��׿��H�fg��"+2d�	7ӑĐ6WZ�j{�+ �K-ȉ���A&�rK��^w.:wN�$�3bc�[W�}����$��9O��y)��S�y.�Dn���P$ �� ׋v��>$�\��"Ob�3j%�g��E`�I읏G��j� �%ٙ S��`bGtU�WM�[P�{��A�$��I#;:����Xfe𛺹i�d�3B���9vh9�����(7�{��y���/�+�ĿM�ߛiM��_�+��L,(��ڡ}�r���_����w� �w�	��N�r���bH3Y�D���e�k��;��GJ�PA�n�L��z�̂��~>��LXg��m��YQt�X���l������f��L�!�0gA��'0��'r��]Ǫ2H%]�I;��2����1�ؑ�>dz=2��DORn$'N��� ����� ���D'�&�쮈���k����S$`f����u�l���W���N�Ӧ�qL�o��A>$沵�eg����y"rZ�A ����>�X���Iv� ��U@���� �ԠA�ͨ�I9��{V�c��â�K�](;��K�1I'L၉�깟	&�=C�'w��&�A>����EOtG����1G"�\@��BE�f2�CF�������{����-3,v��m�ټG(KuN:�k9��A�}'�-�d=��ڮ�Ѭ�?�E��+�$���a��h��]i6�B$Յ�e�=;�hC��A۔Knn0Y�Y�6(��h����ۊ��̌��
t����5��l�q�@ȷk�d�c�6ݮ�N�:���4�y̴Z��ůdiEB]ɬk�7h�5�^3i��i�e��ͣw8�B�H�9fqvh)1�-�vɽ��ٷ:�Q U!��x�۰J�tq\g��+���NFf�<n�\��Z�;����h�s���-��WC@dB��F�%ӂ圇���a������I$��Dl�{p-����l� ������<��0r`d�=��t,�c�,CVYX��}=�S O��t@&Qq{]�/ۿ����z��M��p[I���}�� �n;�A7��n��g��%O�eZ�I�ܩ�_�ȃm� AS�ߞ'�2�in�������S�$��O�yځ> ���\�r�m��"���ə�_�pn6"�w���AU�I�+�����ͪ��:����ݓ �z3`@3䶝��i��kf\S��P4W��rj�n77�^ [�A����t\�J������8r�d�����
%�;{�\ÛA'��=�M7f�S޿�f�	��� �GGlA��H���r]3��1��>>�ȾF����f5��L#�3��8�BrK`���M�c�_f�N���A����9���z��m���ڲr��궦��Ȋ��P�����I\n��HM?�<H��h��[���0.#�d�9,��r��'��#��7��F��l���h�v/b��~"N�a�N������L�L��ݝf:��:򺭂#c�H�w��>��,x�'Ƴ� ��뒿8w.Ιӳ@�<�f��veD��NKۦ��`O��b#!��I�ީ����~~�Elvm��f�p����XCS��S��㬷69X����:LJ��V$ �I����	&�gC����2y�N����+�m{��2���v]�`�t�ę�y�i9�(��k�q�bt �O��@�Fv�L�aޥ���gOP��u��K�%�94bV� ���������C�lcwC�o>nݻv�Z���'m���y#߳P�2��mƱ�C}V!݉��
]�d�����;׶��%X�X}��^z=6o�y���\�nK�P�������]<HY���� ��D�����=ޞ]������y�O��Q��&���o� ��8��뛄N\�r�Q�Lyq�إ#)���;��N���y�<t�i�N-�;_���_邗���,:=l�vht�b��gy�٫��z���@=����M�w�#�?$Aj���<��m�z�מ�X=���͎�}������]g�wv������t��uv�YP,,X�K��j����w.��gc��@�6i��\��;��$zL��
��O~~:9�H��9�:����ry�^��A�Iy+����l^� W�s���Gb�&�ˀ�#��E�^�}�9�?n��5����՚��ҝ���<#h�����`�ѾFe��}�p�\ӯ��ӑw��_@#8F�^�3r�<�d��Z�������g<��W.B�h���2�m��K�u+��uK��"_S�.~��y�}$
�O?g���@�)�4����]�}�,��p�b�-�Q[Ŵ���p�k
ŏP{���8�����T���k�\�qD��>�U�Y�pY�wG��c��؁��M�!�����Y�'n����g����;z-
��ۉǺ�ob����]�^w��m��{���w|���V���z�J9��Т'���g���a��g��{�]�m�o(}�Fۙ�0�'����b7X4��	$�v`��5�,2�`����O���_��9:I�V�\�Ђ
�9G	��%L�(�T����eU�=�Z""\��^Op,PB"�U"(������T���䓒;K�ׯU��Z5j �h!�+�ҵ���A<�8�TQy��<���Qn�̝J���D�ewS��;�r�H���L�g=H�g�';���wir��'d�Q7�\(Q
��D_���:�Np�s
�����=xU�p� ��\����ʈ�D����U+�;rN�s©��"��A���� 
��P���KH�Rتp�'�����
!_lS'wa���;#�N`�(���)[ݧ<�^����h�/\�y�9ȏ��]#�,�H �����24J�Ve��@��NdYy8�UjU9�\���(�s���=Y|�ȎA|ʋ������wwNQ�$�_t=��t���D=J���΁�t���y��j�I.��^�xT�O���٪$���L��TG����f$̙l�Ιj�4[k| �'���ܨ�	��j6��ws�	�p��V�0�&vwgt�j����_��ޭ��+pOk\���$���I�����_P�i2"�i�l6�< ,9���[��� c�r�^U�ɣn�p�D	S�>���~Rld��;7q�S0������Ǥ�}Xb�=Y��j	����A�^q��!pH3��9�rf��i�m��C	�nuL��ns�񪳥b��k��;nB��\�t�A�;f{�ndIjΏA��/�7fQiKeJ{{�$�m�x��'��\�L�=Q����1#�\vV�2�j$��Pkވ �����b�ƬA��\�'��x�?M��.z���eĪx�|����[��ɓ�&��C��4m������CE�x��K2Uu.*���9"/���ۉ'`�B<F&Iِ"dn؂	��"�i�P�Q��Du�T�$���A��2�5���߶=M�_6͵�dI[�lG-�P(�RǇ��6�aJ���=2gt�7}�?���ז��n��}2	I�Ȃ'�-�~ G��h�Pb�3����tω!�y�U1N��@놌GƟ��ֳ���� '����} �z~0	�u�˕-��Q�5�]��`D��"�;W��z�i�� R��8��ħ���n;G�˕7&��]�%�;f{��r�z��*�^.�	'�Z�x�ὝSUs�Yv?
1��{�=PO���9.�9y����A&���A�Ύ�ٮ����h�Έ��~{>�ݝS'�j:;wr
�P�w���es=�r���NS�{�Yuo�P�m�>݃h���u,��/x�Q4=���c�����'���?܁���^��[�}����KjKʏk����{�Yy��'0e�4�SJ�����\Isl�t���H���� Ll[��ce�.�E��ݍ8�I���Dj�,��Ѹ��!+l�ۘ��Ā��T3�HL\�3&�b��j;g����1��HKf��غv��FZ��1C�^�f����aƕhj�݁GB]Ѣ�(xݎ��n�g�����U��t0���e�\/F���Fhkt�TI��"����B����CI��;$G�����|k�������x�i�=�-O� �m���%�3ʘo�;��R��>vN��͍�-�=[�mɘ$�E>��v�TzP4c1n�t��d�L�׳v̜��t�;4�̖�D�eD�	���[u���o��<	�w:�Ey!7�pk�HA�-C��ǫ8�v <B�/�H�k�A ��ʙ'��Fp�4>eyJc���w���셕�v$:L����MȒ)�bUU�ۣ��<��}9yS$����9�>��Ku�Hg�Hwt����ܳ��.Q|at�L5��ZX�l^n%��H���� �s��9�18��f��$�O>s��!���w*ʢ��6p��|0I#+v�o�\����X�2T�@A�����l$�ѕ"��A.��TD�a9ُ;Vp�v�b�D����6f-M��ա����,�9�n1G�3���SxL���vr��82+:�x!~A�2�H'�: �@6.�os!zh�3:���3:,� Zf�fA �љ|I~瀛6��gD�� �o3jD�A�΁jvٓ�v.�;�M2{���6.7���$ſdH��y���|��A s��/��ܫA0�w3�{��:@��";[6 �H5��!�nK�:� �ʝ��I띏@'b�� mڴ<���r]�.�r&ϲ�f�>5�q�|��v!����B�8�ϧ��������2wb{��UȒA��� ��1M�4��W*;]��Y~�g�	��؂��yd�$��1r�.������ �����ľ�ǖ?\dp$�@윈$�t��H5��}��Q�Ә���A��0��� j�t[V/�ޜ��l����
/(͗i�,� ��ӓTUͫ�a�����%�����>g,�#5$͕#F�{_�vb-�[w��/a�^���Ӱ#�t��DΪa�I��p�-3�|�r_m]�IS��y#�m}1�G���1B|lLȲ�����d坋�L�٥�K���"GveD��7��v�W�V���H$t�قNoeD�u��#���a��� x�%���X[ ���8�{)BV�f��)�H�c1��%�yN~}�|�� �	�ۊɸ�J�t�ȟn�ܿ�+sWՙ�}�ٗ$T��y@$o���ؗ)������I��,Y0�W�����*i��$�ovT�>=��^W�v3OP�.pr���^d��i�w�1��D��� ��583����)�vT��(d�3�$U_�?cQ��֪� ��Mf	�_T���'��Ǧ�G��3�]'�燇�l�YV�WM�W���2{�z���Eq����a�,�y�۩Y<ee@{_�}�q�z��3܋.���ќa���5��D�)a��K�dE���I��y�x��Y-�^$,���̩��(�O@��}P_�ϯ~co��\��P*ӽ�i$��e����g��Cv���Ʈ����ߟ~���m[���*;ȃ^Ag>T	 �OD�����~1����kĒ*��d}y�=�B3�d�w�m���YN-��0˯�Y�x�9��>��=�|�[��`�^���6	��`awb�3$�T��UȒMd�A$j'�ٝ���z��dIܞ�|��y�r��t�&'�B��j���tX�_;f�Ot�@$�\�d�c�cz ͜H;�"D�D���;�ށTZ�^	��[���Ec>�QܰH����I �vD�F�W(�a��ZƘ�Wu]1t��1�ؚ��0�����:y�v��hl��c��.�曻�����@'U���=��~[ᇳV23�
tX�i��=����-�V:hU�En������$tԗQ�.&�;F��&VKҰ�i�:�lFͽ'km�ͣS�I�GU��nk$�`�s�܉� a9�[6�&C�)�q��Ⱥ�����ӻ�{;f���/j8狉Ni�Ľ�vzcv�c�ڶ٥�+���;�$���W*r�`���ɝn�r��x�n���y\s�d��ts�v.y^.�Q�M���.�#�q���]6.�w,�=R�6�&�.脖�Fͫa�gE�2����dI�́Ă}���<^��W>��͇#o�"+Ē�?d���u�̃�����5P5�ffyfv����i{��	�9�"�W�l��75�"o�nz�O���s������z=�K��������vݯK�]�|m��C���W(��.]��d9Q=�u9�5���0��.	=������A>���|�7)&�����*���w$���)gg�𷱈$���5@��5�GL�A>'��P�@��ٓ���s͜g׾�"V9gE�?��%J1)i����vc���}\h�F�Y�xt�<۟�Τ���:��⧮ q�\1� �ot��S�ڴ�i�5�7��d@>'��K�ܩ��]�'p���fI�y��5����xݗ��!�2c������M�P���y~��[��+��j^ 5�޻5I�;����[/�=�ք�^�䂋������`�q�bH�;"N���`�v��� �賳��#1<[GWND�I=�1-�0UJ�6	�U�A#��fA7�k������y��j���=frv�=�mA'z7"L�"�qWf�yb��m�o ��b��dt�T�$�M���m�Ӱ��[�}EV��輑 �z��n�O_6���3`��ѯз3k�+��ػh�,E�"K"��h�Kw��]���J̀�ă=� :�&�z �ә"���ED.c����m�D�"<G"[���v �s&��$��v���V,�bIیؐI ��D7�9 V1˟a[���/�^�,1��;�@�>�Li$��ǂA��ak;�����C�T2K&-�6�y˙V�q��e3���iیE֍�e�1�Ǔz������p6�k۵���8.��8ݷ���޺XH$MFd��|�c����Y�N�wd4��Q=s�4SfW]�Ɗ��ؒA ���	��_%�����Z�q��FD�܄l�A'�����R��Eq�q��Bܛ��>$���W��X�F���8vf�-����q�c�Oimi��vٹ��˭��[�9w�Ō\�8ggN�]۸ET��$�؂GJ�B6�m��c^�0=tL��|w'^ �Mٖ��I;;�P1*��t�56:���zb'�n�<I�W� ����d�5�н�!$g�`AÖ�W�5lA$��� c��yt���ǹH;�� -���3��r.]�;�@�Ϻwj^\��a�!��'��nG����^�����%c���ꋦh��`�w4���´[��wgD7������e��qU�_4��f	��,����Y=�F9���ֲ{�H�\җ�}���H%�E�tzʍ4ėr�wd4ώ≆$����O��쾡��"F6��dԯT_��]4r��r
�:�L�4�	���`�Z5�{c�U[Q��9��tS�Gf�f�,1vbį:��Z��$��;�Y�"�g@`|nOD�yleU�v���� �n(&� �r�2wd]�dGEt��$�wvn����w< �|N�=���'�G���-"++�x�:`��0����]gw�1<�`����$^ˑ�'�9.��Ŋ�#�߈����$�HI��)ș�5�)ቍ���G���M��7�l���I�~�k���i"=s��r.�ٙ�"Zg'6�A$��F@�w��77�F7ޅ�7�>$������c9�z��v�۷s\�ɛ��~�sG�O���K��w=�NM�}{R�!}=yũ63�웾�7��ܙf5��խ>��>��t�w\�<_A|���[��w�x���"��;7���̀�&m���ı���_����oN䩙�M�/S�u���x4_����P�/wzz�Rg���[>�*��9����u:sj�eü�O{�f�я��=��7&-�������� �U��0�yL�����I�aq��M�x����E����{���@gf��9�Ah���µ�U�y��:k���F#^pd��J��"`ee���6_��l�{_ ���w_V/����,�c�0]��1=�6��+4�Y,��0o4�{��ާ��V�����F��9F�oK�+�چ2sw���˳���=�R���\^�m5N��^|���3�g�6���Ck���S�}.x��#�>wø=�v��z�/u���a[�On=v����9x�盳��5�y3�0=���oe�Vv�s��A~����uZ�x/���^o4gy����ss�v<ְaG|6�k����
/�lql��3��+>~��*�X�{f҉�u�8tn�qxdw��/?f��AE?"�A=���ٳܷ�g*�x��k���L�S<�ዜ����y}8gmt۳Ӷ�и�SE{}�d/^;sg���ϐ��|�6�v�1<p%�ӽî��Ξ�5�x8�de12wk�4�y�������E�D�~Nv�9�dEȗj[����c�#v��sft�����x�q����7���	��8�`����㹧r����@)�04�q�<Q�F�ܙ�@h�XYI��L�f�
�N�*s3����Hze�%��;�HBØV�\��������#�^�#�NG�8�g.<ª/D0�J��K��X]�].jEEQt�xU:�����8NHUN���u�*Xz�X(JD �3T28z��B�Y��tYE���.URsy�̞��Ђ�@���n0ml�m����֞�Pt�}�J�Μ��!z1,��P�Mu��G�t=��s��.S��]͐Q�A*��*�9zcw)ɡTN���w���R�@��%�]�oy��x��'�I�k�dL��dPPz���A�C��i�FHqT�T*���w��EQRX�Fd�ȫ����5m<�(��2��e��;o8�E{�S��*˙�W*�J.Uf�"�ag�*Q���}�(�쨎}�Յ�	��|��yn�g�ź��<q�M����}Z�gSͶ��LkYet�3hiu�^��i�H˕���|bݮ��g\�:S,Y�U��ہܡӴˬ;��]���e�`�c۵��w>�Y"k��=f(ܼv��{l[4\!���{*Y�mڎ�"f{������u�j՜er�qs֒�ڻ,Z�Y۲E���<�t�燎3\N�e�g�F�n��3��Y��i��Vm��IfJ2�4��R[SY�^wN�v����=X�a5��Q!��نm,K�p��9���n0d�s!�z��qÁ�{�z�X�5A��ۑs��u�F4����Bc���]5�R�ί�a{���s�۬ԉ�`�m���*.æ�]s��xƎ�^���f��'d��eN���mf���Zc�y���m69˕e�x��a�=�C���[���F��ȱ��Xb;����Keϭ�v]������=J�rsCL����^eu�_a]�����C�҂X�j��m�+��]��v�s
"]�a�%�Y�q*����J��N��m.���[s��ؗ^���GՊ��^nj=d4����-#88��1�99�ݹ��H6
:����^nt`��S.�͙J`*����b�Kps���\M�ێ�m�a:�\�M�sn�ݳ��.�y��\��p��q�0q�����m^f6]�@dhuFX\%8A��ю����Vۡ+U�b�3Raѣ5M�W�-$��ΑF��͌�`�xq�u���%�l���"�V���YT��f6�ز-��4���q����K`���Fke�j;JuYX)���8�ur�k�Ur�[���Q%]��1��s������<�.����f��� sm�5���Y7G!�Mt%�fl�8nw,��J�.�n�P�ݽJݻAWl�Hβu��I��.�RN�`s�]-���z#\�GP�%p�,��v5�k�5��ݍ�n�����^��s�k'�{y۱3&�㓍R���������H�+&��+�Wf���v�a[�JӓTq*�u�v�#ٕt[)ѳ�����v��-��\�ȹ3�`#��,��p�
��k[�	a��]fwO1��4��6v5{�6�ۿn��|M����҆�<�M���D�9��6��w#��� =B:�������^���Cv��n{m(\�z��X�j�E:��"L]���]���RN�f�t��T_G���oc�k_��WOMgݏ}Kh$�����a/<H��=�} �g%�xx$z�4��o#zd�|o��9���2
���{� �	=uIpt��wt��]�����>'�.6U>�g�5=��d�s�zf��$���FX[�K����@��r�8ZN���C����G��%�[f��(N���G<�L��	#>C��): ���F6@N������H�ْI7�0 }�o�c�v�]~���~z��Mj��*V�*k,�6�aoXʑUh���4���,k5
[�����V�h�Q���ƀ �|v-���z����Ve ��r$_LE[�� �I݂����Tff�n�}���94:�Oh�/E�����������{�'Ǡje>~�/
��\X�_n���;/��m���y܉��.md�Uy1Ă�LA3佲�� �|�۰ʻa��=o���`���R0� i���Y��$��T{���Hۺ����Z�\@ ���	Q	htΒwt�;N�����.J��wY���#O��I=Z�Ē;��N�^��k���� �i��\3;��1+6"!�չV=Џ���H�ˈ$2�@ ���'�媩�=O��'��ȷSS�.�p,n���v03&�fFX�3����v	�ECwm���S�'B��I��Y� ;��}�1�'Q�Fe�{�]wI�����������a����쭙�D���ago4@$���PH':;&I�v&�:�-W�ѐ}���.Œw`�4���lI<��I T=��p��������E��ȕhM�l�f�/ys�r�띷��|o=)��0��ihNgor�h��p�
B/�F���P���˘Q�U"���|f�I>���/&����'��a�A�9�ߥ�u�N�3j��I��3�H�~�-��ʫ�Cd������Ӻ)��.�=SO����vv�ֹ����PI W�;^g������~�l�5C�_��Eܻ���lk\����g�U�ٸ)�ͪe�sX`�����~��	-� �t��|J�^�2��}���f�ib�'A[E(�>$vB�$S�(ϙ7"�v ���@�x�f�Վ��rTV1$Ϲ� �I�~�����>�P�W��hz����vL�-2"�zd�I�|�h���~��gj�H'�7�Y�u���
�A�"���b� �)����7��Ҿ���9�q �M���ǉ�>�l���T�f�e�l��w�-��=P�0*�Z��0��o*�{��w��~��#��Xf�e7���V���$��"25�(�9"�RS;Cvǹ�"&�fA#.o�������G�A�[�ŉl�Υ֯ 싺�� m�$v�C:k=����Ϸ���|UfWf����7k`��ڞȎ�'Y]�iNv���N������?���N��gnᵷS �H4���y�9�'���B��3}�>'�^>�C�e�bAm��S�]���A��5}��}���"#$�v �u�9@$�f�f�K�FЩ����'ٱ�LF3�Ίv(.��$t+�� A>=�3@�}����1uv�|w_�EH�l���4��;�d΋��&�m�{�5K�y�|�^H��A'!n($�k�l���g����So�^��V�;2L��3�1MCA��ȟg��s(��$�H��$.ʈ'��5Z��H�n��}=G�Y�r5�Б��[�@�
쌿b>�I?_1*�6{�.0N^��{�'�gދ�7���1�}�ݶ�}��n?T���i�$f��ꖋ�����ѥ �WD%��N�����)㋍�{#�F��qfJg˽��GnV��<9�S��;��D� ���{m���u��Jᮬ�n{y�Zg��]�N:�k��v�6��k P��ڔ�2-HV0m��+7;R�f�7BR���,��;�̌�
�P<=��/�ƪ�d��7:AN\c��SbS��t��r<h0Ɲ٩;Sn^��0Oiy4��ܥ��p3l��:��k=��t��$|��4��'�~,a��u	&�v�'Č}�&�'Nf̍'t�gD7��6�M�X��IÂ��5�ˡ@Y���������H9
�$c�lψ���A�#��mlVL��`7�h$�r��d��|H2��O��+Z��������"�����ٟ3�0�4�sL�aUⶹ�c�F
�ʻ`��.����5�$�{:6AY:y�`C��ކ�X�T Hz�KK��N��pZf;+dG��̘�KI�Q�Y ������>$�nt;K�n�����	P�Ç�5�k�3�^{���l9��٨�ڹ��V�n6tU���Aْd��X7p9������'�s��=ٍ�+i@$/�:D�E�b�O��YC��p ۞�ɠ��8�Ț��W���p�(�7�s����p��*�Zf�=3��݆�ĭ�����;���̇ym���U�s(4,��׏z���!efU��>$.�D������<Z����4�xY|�eA��ݜ��9.�r'�=`Έ�A̧ن�iɖ�+z��
�sb@'�v�D>Q����I.�;�H1+:��w�Q	����>�|M_D�5�2L��U�ۇ����{2OK��� �'v,�&@+6��|	=
�<�դ�5�Lo^D��F_D�����I!����(y����$Iı��s�G0a.�&�:�FG>24�9�ay�8��<�}�R���t���+g���C� ���P+ޑP�7E��[Mtω���'�ҏ�0�)6�X����o}��?�����N�X$�Af$f��DyJU�A��J:�fFS5OMl�a���1�'�qL��E [� $�R���H���n�Wϳ��J,���O,�qmK$"R��#��/`�uY�ypЫU����{g���S�M���{���7L�V0u8�-4�@�Mv����>PuJvwE'�9�u5�4����|�H9�Qē�S���NF?
]$eOS�EQ���7�]�gi�s�9�잉,�1���	�'�	���������:.�XP��'Y��@&�<C�v��4{KK��d�.`7=~������3�5�z8f��	'w�&|b9t�m��Eu�z&Tm�^��G�;�:�pUTt�L�YU��j��b$?��9��;�rd�w۹n����3��f=���]:ggrX4�<n� r
���Ƞ|��y��ΩGQ��� 8l �ӓ y7Ɉg)?��e���[���Az�h������I#��A>nt �ͽ�GY6��:��2��.g�ͧ7�o�i�v�W�_��5��b��v�ow�O�gu"�I����{ꬕ�6����Ӷ�$J�Ƃr�ڔ�΂N�c:�SH$�������U/X�N��3�;2<I&��"�:��fPW�|����_z�bX̑ƏR��D�Ai�V�F»@#iB�tP/=���g착��ئv��/89�=�� #�/^��x��&~ٖ��ce���w+"�.�0ڃ��va2s�z	Ŷa�^��7ŷ�d�!]�3$�oz"4�m���<��wxOv[A!�i�������S>��ٟ��M9l[���K`$���$nt�]<k�t��;;���A�uN��PƏS�KvnĂA'�e��i��k�<�B�Q3��p���ݫ��3��Ό2wyq�ăF3��u�e�o�@��ݲ+ԅ�Lz=�+��=:�%9�8����@pG��iͻ���{�.Ԍ��5�`�]BN�׊*���Lf�E�|�
+�}������.��y�Ge!�w�G��犸R��U�
f�W>��MŹ����m���:x��:{��@��K<nKA5F�a,b�̺nEf�h��ǹB�жUӺ�{�x%���`Q�ܝ�/I0q�VQ�����v�n3��b��n��q/=g�e������ɋR�$���,7<ˀiv2��Ԭ,4
�UM+�]em��"����V�!Ƥ�ԁ�%����k�����S�f���9�6�F[�+\��Z��;YJZ���g���\��M�T| ?�/� �|H���Zr� �r.z�vD�k�b�0���%��|`�t �VT�^ݝ�w��m��I͘��u=s@$Ʀ�=%�A��M<"�s�0g.�L�n��/��2 o����g�X�xs]p�A���� '��i�������S1��9Qm<�Q$�׀>��m��^�詙��|Y�x�x�n؃|�n��w,�ܤZd7UI���K�A�E��H�=���ƂF'�h �=��u@2�����噌���z�`��+۱�`��-����:dxR��`��6f���﯂%��m�!��� d��9�O��jd~��pM�L?d;� �/��	���S�:r	�k��� �͸/^�B}�IC2qL�_�Z^P���\:�_Mś�ﺝ�v>'ܑ�}g��(�Y�_���5���&z�l�Ed���2�̥�@%���-���ʉ�Mp}�E��讃�&_x�bX�೴ό�h�ٵI���t�y��V뷁'� �O�#{��A��I��0w�U��q���8ՃΡn����S=w�$��ҵ[z6���i�l���)��U�vw^g.
��l�ț�@�Ɍ������2�Z,��i&r��I"��l��j�'��
i������1c�A��
kt��U��]]��ԭ{8�@8D.��t�S�I��E�])�~<
�ʉ�E�LP/Xȡ����ؚu�';��|H�����'�,��%t㊞J���`1���ڙ$	�� ��5���+�&n�`&v�N��IӠ��gc��rHH�o���N9n�M���<c�}��G�����1`�iMXm/e��!Ӿ[7� ����g��n��#��X�h�Y���t�ow�M�8�M�B��	�=Է;Ĝ}���~zxa{}�����$�Vk�a��7�����{���-��O�c���Bx���K�2oz{}���w�gH���jsz��zȋ�t�f>�n��f����.ѯ�K�L��ͧ��i�AV���u������[�5�A��h��"�^bQ�v"P{J{�b�����mH���y�nO^��|��9����>���ܽ؆����D/_����-��<Z��`1���R�og��_��}�ܻo�{�k��Y��8ۗ���5�����/leg���G��|�lޯ:_S_ywy,�z����=�$k�F��O�b�"+�*_�͘&Q�/P]p��3��;�>��@=�קn���%c���8��8/�3��������>����u�Ԍ�ّ����z4vT�'�J醿v\�{��	���}��h��W�.�)wq�e���*�Þ؆�-��ޗJ41���;�{�~,e"[�Nb��x��/f.Xx�l�k3n&�[���B݀�=�C͗Wb[wҳ�#�rx]i� �ٗ����^����^��.B��5o�����B��)�6�Z"^��4� �J���r�Yל͊�1vv�PL�EO��]�+�w|�p��C��K���/��v
�2�gh�n�^��n���xE���u�C�5.$�{&��|+�l����$�P��:q�Kې��Q��2E�g�ÜH��m*L����q�Ȏ*�K9IU�Ri���9�*��Qr>�N����ET�H*���DU�$�S�!��LTɼ����"(�����E� �yX*)  FɊ�HS(��Ȩ鲋:p��(��$�L�,��LNG3
*��V簫�Pr��NQUW��Er ��2���{�ˑ��S�AU���2�7R��!Z�NTU�\��e�Z�(��DU[2��3Ҫ�DEQÕR�v;��՗U�W�{���t�L3"�D��q�m��*�v!�*���HrB�'J*/w&�������E�EOR��[�3֩E�.g<�Z��C�N�D��
�9���F	t˓�q��L�ղ���
恋��}.��S^���@����Uq�S��s�XLǶl �-B���p���M�H(�|��I�{��eL�I�� �Y�3x$����pl�M��x������s�^;-\�;4K)+�&d1�$zC��8wa2�� ��y 3�f�b��۷�\�d�+�Ȝͨ��D��r�Y�'e����0�'p��"|@�A�l�F��%�%%k3��I��\�R�
_ɻb�3���9pWp���	7�O$�l�r�]ι��3�x@k~��H5�QO:��'vd���'�U@bV��7f��+&=^$V�D@'�����X���S����dr��I��K3���=9H�Y����ii�Υ-5��)�l|I�ڈ����>����9E;:���쨹8�;����� j:"<j[qG�$n�T���]�
ɥ*%M���M��.\q���#��[9��V�;�O�M��)�����ljyxKS�ݝ�.��6Ecm�ϻA �>Dd���"O����	��M�L��wTI����v��K���A�W�	'v��K��F����}~1Qn+�.������h��ç��%�v^8�W0�������ߦ&�M6���=ߖ�'�ԯ 1$�ʉ�f��ڳw�<��a����<	LW&ww>`��ӻ><g1i��-�Z�	$���x�3�*d�6����t�cu�8d�س	4��3~bF�eD��*2p����.����ؠw{*d��ZIr�%K3��];O�r��<����#�A$�^��$ H7�',t�
�NG���[+�{<'f`�&gA��#f�A$���SN�WC9g|���ۙO!n��H&�����.ɵ��&�|�m=&�(KŽ��wa��5|�����o�ެY�^N�t�5�+5Ai#n4!,��(D:ٖ ǽbg��4�ig��,>����_��7Y��-�k���ӷN���z�Y�\ag׳��<��n��7P���N�#�ND��f9�;��v78���i]�]�\�����|��o�{=�*�yy�����жx}s�э�l5��륬�����l&d�H�5ֆ���e�7f���K��s��5�6v]&c��sUI6�f���r�vRs����3V2�&�D����WP��C:��QqS탖�_o9�	�h8◢���#��Q�B\iص�=}��u@�	�������x��[�Q$��}�"�N�~��gb�q�N�*<H$UfT��2��.C�p�݄�]VN����❫��eN&]� �};�3 �M�K�<A;�yF�B��F���c3���p���l�L�����<��	I;G���Ψ ��ə$�}��y�N�;8f৙=�k2ޞ�on�p����y�}���A-֪��zړn�t�OEL�'�	�@�L��R����l���
��>n�M��i��3q{3�O��ہ���=L����\�nA��_%���v�^mm��2Y������2��K�leF^���������d�2������ܙ�w:�G�WZ�K�E�l@06��fH ͷ��A`N��E�CG6�'ޝz��y������N��]<4	nuj�>er�������7[��ñ�C�S�4�q=o#7%�(���r���[�6%Z�I�ǌ����YI=<�D?��d�#Vij\ӖH�2��n��p�݄�O��l��M�>'��:Q���s�js�@$�S�� �2ww>`���Y%�,�w�-x	�3�Ăwi��$��闘c�x�'����6���;$���3��Q�ָ��y1'p:��	X�MP�`��Qq �Gm=� ���w�F�ܠ5�fw�X]c���#�2鞳��5���Z��ɥ�3sC��Lr��^���Y��LY��ܸ�YMЁ'3zfLm�5b.T,��^r @ ��;7e�S�`��w!�L����R���\�4��O���^DwtLωg%����r���p|��00��r�]��\�sA&ozbA$��������D���c���ٶ�0�N��(7�Z<O�7N�6P�H��_#n����K�/}�k�:���k(�&���HY
����>$OV�	7zbI�\�D��A�;�N-�ޛ��5�T�!��1k��H'2�d�B ���������KSf��`��S���p���d
�x!��5��+nȾ̀KCL(�$�oLH���~�<�s��厕ehwt�׋���8.C�)��\^<\ny:ϑ��`R{K�T��\l�Y�������et���3|GndĂ|	����Ş�s�d�g+�:����yD���p�Rb���1Q�{jz�]��tĒ}�q �8zR��^9��A"�>J,�ӧS	�ٛ��^�`A� �x�[�fh�h�Nk;�N����[�c�q��%�<��v��vή�Kz�H$z݉7�H�����kޘ�Z��h�>����w�FR�z��e"�����hԤ9�ׇuuY�C��۳��Sߧ{I�D��7��[s�71�V�T���_��$�s�D��A�;�va2<T�DO56G�=�����&�[�5��H$�u� @ �sY
�����0ƛܞݙ	i�1�&�ф��"�h-���nl��5�R�4N,	��;7�g)oDfd�Ǟ�=O��������2�Ún�A��@�U4ܜ���'I<Ϗ\�ǐ�r��AOt�H �o{�������0[z�[�ݻM��{r�u�r�Z���=�1I4���%D�K$��7�v�$O��|5���PȝI��:t��aU]3s\ϵ�m�3�>[v �O����$��ٞviP3��t@F�q���%�K�7��7�Q&���ݱԏ*�#��	�@'���H�홓�W>c��ތ%�K���Y-SF;f�R-�4����>�}��q77���[�1��b;�.����i\�I����(�{�N1�
�{e�a(%�`2�X@/)<q���iC��Ή-�Ds���`�'m%s���6cn,�&�t����t�]-d�`��h�C�1T�6�w���j�,�綺���N��g�Ht�:�YKm��,�ݸ6��)0�R���\h��$���ن�݌�7
���C%�&$%u�X�L��6�V+a�Zq��{l��W�s��	l�v��i�v v�{I�ƍ��B�ʚ�A��k����a��~���}O��1�;�vaT�DAƦ��>$�ى2Ӗ�4�(s78�m���+�(k��ق,�%N��oƲhƻtn>��������}|0g�Ȏ�ڙ>9�ƻc��[�̚nA�g,�t^d��y�A �^LI$����ؖ�g�g���x���1$��W����Ô���=�1����۱�	.��`�ܙ�	���>C
�ي���$Dk���q'�&��Ô�s�* ���]ݩ�f�ob�ۈ�gwf�N�tg�:�X��ήvL�ɘ��'6���˷e�MǠS��׵՛m���܊���~�ﱒ��(��ζ�$��ى�I�>t@2�1��S�����r�`M9���tΓ�gf�&��#��힦���ñ�$�z�7=�1�g6p�`}��?-�0)�|Ut�R��������1�Sj�c�QZ��샶�Y��c��E2LO\SG"H$foL�1��잁 ��&q��F���OF��w`œ����d�$�}	0�a�V�ηd*�'�ۻ��G�{"=!�茸��2t��NKĞɗ[q�3�մ�-�&#"H ��؏	�O\� 3�MX'��S3�|���8�9z0�"��
ݗ�S���u-��N	�3�I7q�#Ď��n��Z���1�]�z�[�d�b]�fmX7E����X�Z6��%6��-�m6���c�|��}kf��;�ú�f�A!��t�$��v8�o�d�_
h�x�ْA �F�>b0/1�d�!� �^y��:0ى{�ތ�ʎ��&�:=��� BjR�F��c��N�$S���t��;!2
����W�3;�ߒ���2=�
X;�Gx�X
��e܂�u1��#����e��C=��<ت��75��Pќ�Y�q��nю��-3�H$�GCǗ�[�A5:Ò�ݘ�N�����|��q�7Y�x�w��A ���BoF���C����]'��o�8�,��7b������ؐKr/F���j+��A/�p �n�j<H$n�l�5�$^�ix��עy,�f���7bKE%��de"���e�n:���(��]"��'=K�]���y�ބEB��NoFD���wwP����ZzN;v(�"�\-E�9vp�	�oMԉ6ժCU�5��ހ|m��wF����f�K�1��ӯ ��p^cl��i�����7ӱ �`fĚf�.:���gO��s�uy�ĂFoT̂i�by��vNX����a�y�tP����*v<�O��rdO��n��y�h��R		���'2-P�T��WF�C�{}'�����w���Z`��-�[��$\��F�>�yG�Ѫ	�zㆵ��wf,]�������A漈�-��m��#'@�4����=�S�"
n�|h�Bb�1�"��vD&�:/�@0�XSٔ��{L��a��i���v;��~?E��vgo%���Q*	9�9�H'�����z��[6�7��9@�ꮜ��/��^ӎ�z��.�;!��wdA0(�lO3�$�;6vd�y�\AM381��疂}����yݜ�$³�����E�~���!께���r�	'�'�A�v���^c���h;J�`E�E{"�A ���	 �9��(x4�OR�옒}L`C��軳��J��I�^C �u��S���m��y���������uR?��
+_�E������J*?�� ���,X��3��#� �`�E�PX1Q`�E�X1QcF�1c0Qc0F�TP(`
A�(!��b�``(`�bj��� � �"�(�!!(�!
�(����F�&; 8FL�
�"�b����*�*�b�*�b��� A��"�(!!b*-X/� ���b����
,��b����
-�oʋ���b"���
,��`����,�J�
,��`��� �(�����b�چ�l��`
���
,��`��� �(�`�����b����*,��b���+*,��`��\��@ƠQ���ª� �+ ( $��l+�����~�`}�������S�j�?�����������?�PbU}�����?�z~��(����o��ު�
��������A�
 p����E�D�����~Ȩ(���9��V�d�]���A����&�~�~A��$���U*�
H�� `��"1�(�"0"��+*,�`"� ���� �� ���+ ��(,B*,X��X��B*,U��`����b��"}R��ߐQ(~���l}��� 
,��� ��
����[��w���� {�����
>��7�����~���_���l��lO���������s��|AEh�}�~����ޙ�(��
�����������˖@q��6�DW�@)?��u��?�[�PP�+锹����E��,
���}����O����~��(��OĪ[�3�>����P��� >O�h@�Ъ
+�g�C�(���� �B��0'�o����I�P~���}����&�����L��N��R����������|N���~�UW�>��l��
���^�n���!�'��(+$�k'su��(�0
 ��d��C�|��P@ 
   P@        �   (     @ P
 � �@ѠR���QJP RJ )@� 
�R�a�P))@� �$�(4	IBUBUE( (��                                              A�^٠�@dh�+- K �:.g@'N� �Pdi@� 02u��@�Q!I�x  �<@FN�;\ d�dvӌ��<$J��P]8 ��7,�o0^`�4U)s�@�"Q! �           ��()��@`4��r�9�\��;�� p �0n`=�0y��B���  #� : (Y�^{�
G���U�4�x   �y���9rv St A�y�<�@N� s����yJ�CA:�� ui�$P
�o   �        �����b$�� �h8 Y:�iZq5\�i����:�� �P�'tj�M�5ڠEE(��  ;�x��;kswbT�� \.ڥ�.��һXkss�K,q:��p =ǽ�/1��,��jks+�0��P�� Qx   x         �,�B�e��й����ͩJ� ΍���vm$qwj�\�k����:8 �vղ��V�s\�@R��  4�3�hl���b�� ��.ù��v����uA;.[��� ��;ۗ�k/;R�[Mq5�Q;�`CZ� /  �        �
�&���˭�'R���!�t38 fq�6g]mj�v��l)R� 2U,�!]9ڕ����(�  ^f�^1��� p����Zq�����g ��# �uUR��bhS�S�4�� �Oɦ)IU4��$� �OA  Ob�@���2`&5Oz��*R�  $ҁM�*B ���ʹ�Ww�Dd�
aM'Y�u��k5A���?�!!I����䄄	&�!!�RBB��䄄	'��$ I @$$a��W��M�-���Y��,�:����"��S&�so53{9*�J�Tv(�b<{1PB(�:��5X*����`��[;�X�^ѱ�@�o\meYA�䑐�ܛM�C�Y�<���.��b�mˈ㧺6{�j���1���n�N¯cTFg,���fs�ƛ,95����L�
��+'C��!k:�TkS2T�M���Φ���eК�v7�E����F�Ї#��9P�R-�퇦���
al��I->l:N Q����-��T��������y�pf��n@�A�ɻ[�`�l�� �qQ��MZ�h��vD���]4��\���9�w<չrF���9�ՠD�j�k6��	Xr�dqR��]�w�c	��H���)��3��4,�7�&sD�Q&WMǍԶM5]6j�!,����Ob��b̷�`��͹����ɔ��L�kk {��f�ey����[1���Q��<B.�b혙���c��eɶ�����^�٣u�I�����-������y��0ok"��9j^i;���D.�r����7yn�I����v��r�k�S�b�WU���A���s]���˅�Rq�<�i�q�s�^�ik�z���æmlR����GC��������Q��P�F���SS{7�ͱY��q>�x\���h*��:�3s��H3Y��F䝳,��v*��.n���Յ�w~�zngns�'a�>#;�<-��Ж���8鹺�]�w��=�W<���z�y��6h=����.��,\9+�����!B>a�휲���t�Q�e��k
cm۰9���Q'Yc*P��ɻ�KF���,���)�W���ϝv�Θ��^x�֛��z���]�.Y;4�KQ�pf6�Ddk�@�w�u�ي��+:9۰�l���s^V�[��^l�x�i-n�,9��x8�d�Z��bU|���%��E7f�&e{��QJ�2�>��ۖ���s�%��$$���Ywӏ��ǭ�1���'t.X��;�f��������n�g0oj�3j���0��� ذ�˵6FL/+S�G�J=�t@my׃�r�%�Zu���͝��l)��yob0�oX�vqܼ�Ԁ�P��К���"�m:�D�d�Uz�t53�1Y�t��O�wv\�,�X����S�th�A���
h%N��\��d���]�~3�'�I����~�پ'"���~m{v9b]�U�9�����}����^�^�,��`����5�Ո:q�374$~��w�ӳ4m-	,�[`��j�#��P���~y5��݇��A�y-[Q{l�o���JՅ{un��]�A�"�Ltگl��y��p� ,)sb+�I���w�]���֠��1��7�>R����Y&s��k�h.>z%�q���7U�jƯ[�U��X��Ҟ��tj��-u�� s ��
;)Na�˷fi����o�D��.��L�\j��Cl�ضk&��b�\@-��S�,6z��n�������9��}7NѪ�r����Y���|7xrq0t�ձW�3BR�8� �"`�ظ�.8«���ͽ��J�r�v��>�>��o"��!-�P3��]��ݺg2�=#��d��Ow��:N2 ��)�g���#���n�2���s�i������lGB4K�F^CUkX
�rB���ZY��J������t{�]�8�v��0=	8zp���k���E򐶓�ѳ-b���:x��/%@���x�0�;��&�L�QC�&˅H8bǱ�o��Xz N��D ��\�H���ve�6R�n�<�k���";s�:�(�_i�qWI�,���lܝ��[ݽr}�D�������P3�r�6�¸�p枏fw ��è�9!�.4�۫{�s�����m�$�\��\��nn'��,��<死���� ̎AV�anL��1f٪N�}p\���Ǵ ]�[��TO�s�{�����խC�G+�eܠ��G�UW.Wv-��i��X7P�C��v�`�x�a��7:w�3� ����m���Q�.}LY�l��<)���A���I=g�g#�"XKP�h�q��g�`aA�,�aj��sD�qa��g6o}�p������7G-�"x�]�,�+� �+k��v|;{e��eE�eQ�F��U�w-x�p\4��R�/GI�꣒D�sX/E�'�:x��T�	��۔����iK�uO���P3w�wn��T�Ͷ�Uvws����ڮd�U3W��ɷV����=Hxo[Ɗ�1,��P�8ٝ�NwGK��Hw�dY�i���#|�o7F�Qm�©�;�����،x�{���i¥�e�iС��Y�h�E��Ep+�t�>f���75�!�V�݂rw뗖�4�͝�r�5��T��i�J��͢n�7�B�א�ABy�{�����:+�f6ysQ�F����Cu�*1v&�ر<��#
*$�ӆ����V�Ϸ�����k[��xFN�0r7+���4o�5�Qa	7A&��X���0�A���Z.@zۑ�&Q��Ԯ�UT'�+h������&�v�&B�vj&��[#]����Ț�j�{�fT0�וWvSH�A��Gon41�YD.I��� �6s�<�N�����N�ڛ @����������&{�͙�=b{ϯB��1��췷2�k��m�,��yT�F댟k�V�{��U�-�J1w��w��E�����jy�fsܸ ���<�B|���N�U[�U�w�iڮ^*��`�i�f�*h����-�սq�	�v��Z2tJ�N1�,?>��Q�J�ӵ���%wo6p٣xO=��C���8F�ͧ��/b �]8�!&(�>Rk0�Q�B�;�G[�%�e)0D"�QL�An=kz�J��i���L&%��x�׶�k�oQ�е���ג���僴��$�%���i5�k�2b����gj�c�G��'�b�Y�����F�a��E7���!	��%�
r��T��ݠ��H�.}�N:&�6��,=G`=���Z)]Z���ѽ��<uq]+�d�H��<3h�ym���/ew�4x��4�Y�"؂!�=:�(�׫���Yi�u��6�Tˮ ���6Ė4��7�kW�g�UE�V<ǚ������l���k7T���wk�8b/(�8ӷ��`�Iض�.���Bk���=Ώ 2l�g%�9�u�pL=��d죠k:�V�A<� �K�K������V��0�I��\2c�qoon����ު9��{x#�_�;���0�ǵr#VLՎM�e�L+i����wh��\f�8c,ѹ$Y܄�"��᧵��qHs-�sez�[��xR��g��1�n�+�������c���9����}p�CNa����R�BI��L��Y�j�F>5^��N>�<�n�Wi����Uu;́D�ý���/j9;n��ٷKZ���'Cco%�7�Q�Q�wpY����x�DpAu�U� �x!�֭I�}c\��&��^�1��(�t�F�`�9��)[���:`r㩋��&�ww1��%*gf��sH$���\��j*dq�Y�gn�Z�
+W:	[�sit�|.�v��뻱b�k�p�a����X�|z)5��!o�����oV�a.�Ɵd|{1��!D�_w�k�֨�R �̛�mis���#����Uغ��w�R�N��[�iZޤa�x��hw;��+n�1iVM�B�,��]}���7�ʒ��޶������b�V�&u��7U�x'�v'�����&���b+8bk~�cK�r�2)�n��69���B]�j�I�.��ɊYm�#6ÓGp����R�q��Em�յ�^�1�^�zsצ���� <[u"�穌�����k{��e�N5M�q��V���n�X$}�k����U�$c\-�s`zj騬#)��b+:��\5�g��-�g;'�j�f�w63x��ðC�����	!(љ�}"�*
�e��Ъ�.�ىbE���.�'3Oikͻ�%����r-��7Qw��f�՗"��]�78"8n�;�m�[�Z%�Gq:�Q�d{׵��Tb�<�㇊��u���g
bbMi=$S�T�#c��ڥ�܂������t���.l���{H�v|^�����۹��oڏ�U����1]o���&��%3���pr�fL�!|��p���4TVv�y�Cx�U��)��Q9'ôFov����Hwz@���zU2dhwd�wv�n�kw�5t=��kX�x�jpf�ٚ�N����!�xWn��]�ڭ/9v�׾�:u`ͮuKôFj�G��\�_����q"��qUO�L�j7gjP� ���m 7�ɝ{�3���/6d���B�%�1=��%��D��`7r�nĭ���a����d��t�hK5�0���e�p��^[�o5ٺ��KVp�{F�٣���%��m�\�ɽvܦ�Ҽ{�Y:�𗳐�L+b˗�L ZZ��]�}��h�a-@-,�-���M��c�i�~�3 i#���,b8�`�s��6����Y٦�	�N�	��މV(0�nU�����[�	R�֔Z*�0��r�u���!��]�s�����N̆uf��H0�#1J��s� \V��䳎2�� 5�������ל08~#`n]yZqMAÀ3K�h��	U1Yͅs[��J�u ���/W«LQ�FM�׎��	��B��4K�s�hB�f)4��~4'a]i�4a�s�
Y^��s�a�D��#X��zx5'A/Zyɕ۸�á��O:��ۢ�����y�.i���� �:\��8|�a����r���L�K�]qU�%uå�D8;r-�V`�y�Z���u�h�XxtL�x��S֟��sR:�)�^v�[�LO��X��h/'��F)zLgj�dWxכ����靈.�LIԜ��M>�D��w=�H����������v��/�lӀ.r��U�� �ab�
jB8-Zm�q�E��e���
�a���7�w�k��=�a�{ֆbj�w� �\&n�Kq*��=;g!u\��M!�	��§%���z���7Zgv�h���A��%8�hj:��\z��ѓ `w9<2�r�.\�99�)�E4������2q�]l|�B;EKqnNv�TK����1��'9�6��q1]!�ż��{�@S	#[�CS]�%���-#�]��qK�����ga)�vd-<�������d��2#9� ]�	p�NC���X�-=]:.�8��J�wje���Y�l�R7���Us�t��u�`* �j���N^n�`��2���ڠ�D 3]��GTR�\*Y�f��.�X|�v��l-�v���rW"���K�<%yĤ�w07�a�E��7��
�K�d����(8Cn-�����!N�����8�V�Όu�r��qp<�M̪�n��a�2t�[ӛ��-�RѼ��q#�����a6v�GD9k�!��(�m51� ur�>ݭAE�|jB����n�(C9�v^�ޗ��&<k�C��L��ƅ�Z�Η�F��D��%�Ւ�7��8�6p����)�w�wI�71廼����.l�;��;p�7wQ��t>�-��%ҎF��]��G���b��A����$j-\/�@�3�M�ˮ�<�'=�șs|js\�I���&�`�s �p���u+�GNW�A��w(T� H��k�ɧ^�.���Y��:y�6_�ˉ��=�\3S����&�{��3��0E�v=ش�¡�v ����u�[���-{M�a�
��w9�fw-�;":�v֭C�|xkۧ�5����f��t�d�p�6���X��MJ�&Z�CB�ǭeӐ��h��{XG;y�����kD��`�5��e<{�w�׸G�>y2�=�;�DvT,7��LE������n���d��q<����1@Z@ٱ�c�54����ݗ�A�nߩ�.����x7W-v�.]��`�7ۛ��0�㐄���_'�<�̎=��J���i$q�о07���9�9V������	�:MJ����Ĩ��h�ξ�Xw�%��P^��o�N�8�}�n���/��L�0��0O�r���ŧGj{��w��ܿn� �*�asv�~%-�����T-Pɗ7�=ק�壌O9��ս��>-��yZxҹA}f�0��/uR�Z�,aY0��a����H=j�L�y���B�ai�H�rq��*�*.�p
"�ɻ��n$��I�h��݆�ass_o��mK8R���Wc�a|�v�t'p�XUP���x��<���r��n�nY���j{�tg6 o�s14l�[,����Y�3����v-�7�n7~6����ӗGEC����;y^\��F-�Yr��.����E��ͪ���Œ0��;��I��q�Ü{�;ޜ�����:�m�C�j������6��I����-QrBw&\m��:t!�;�v�yk[����7zH�M�+����4�oF���0o�6���k<V��v����Mx&���,D5���г\��<F߬�٣(7
;ʽ�� ^:z��zH'�գ����k��=�t�|^W]\�cm��Ժݛ4���3!�$��I%I$"��`IP�,	"��RI$!�I� �P�! ��`(I XB,� ��,d�(J�H$�!$�	B��a H�	VI
B,�!�("�H! YE�
@ �� ��H�B@R�%BB@�)��R�� T�E�,	�J�`�H)��d	! T�IP���$$�` d�����B� BA`@� E$�
� 
�T���*H(I"�HI H,!$�R�RB ��� 
 HT!X��$I$R@	T��I @$$]$$ IY�ش���JT������C盚�C�s�^��?[-)f��iX����:�&����9kg;l�{��_;:�ô�3�}�6vgI�3�{dU��P_*x�������,��YsT���wϻR}2���j��en�����XK;/�}i�7�kNqo'9�.������/��Dh3�p�o���{wO��۶�Cb���T�獼��]����˵s�@v������8=-�(Z��w}�M���:<w܇�>��>^�� a���xņ��_6a��]ˋi��p��s���E�,~����J��5����NtFvk�=q����^d╎�Bj��\���G�1A��p<�L���/�ջ<-���I�>����hX;A�՜⼞�<]C{�ׯ��\���w�5痑����M��J��<U�?�:"];�E|�S���MX �ﯗ):��������3�][� �=�k�F��܀�.QAѾ�ܞ��]/x���U�&�1x�Od���nz�_c���ѥk�!��jt]�e��|����'ܴ{�{P/�/ry�g\}�jA���f���H���2���-��wo�:X�
7V�1OM��F|2����|9�ΓĈ�BP��Y�2�6fXڍ��U��k莫�ڜ�̓�����!
0q]����Q9�z������!}h��������*`/���}���U�֟=]�����̤񭫥�!�ȳ�����$ח�t��Ph������Z����K���}��-������u��n�"+w�N5�i��DӇ[t�wlPC�t6���!����J���*�^����;\]3X20T�,���V��m����=��$����_c��,7پ�7]�w���#�*���j�<]�#���Wܲ���p�[Ձ
!���S	J��][f���s�Cᮈ�e菝ީ��t���wG�����v�a�BV�T����:�]f�N�gt�S^�.)���烾	���f����4��Y������)�|�]Ч��qP����5�����h�L]
��_b|�ֆU#�������7{|����rB֖�����]
�g:=�:M���ܒxqO=�����߬���0u����Yŉ�7-���z���rvs�ƞٝt��r��r����"�B�|��=�I�;��Ʋ,����=�:��x�3��}7ޙS��:�w�	���>�O[z"��6�R�i�]��n��e�سm-�����ޖf�y�>8��0�{��Y�u����q�jw��\ש�A��zw*��dr]�@��-,ݳk&�#Y�i>��8��w�ˍ��m1H���	��vK76�;��NvB7n<}�U����>w6w:�/����T0��iZ-��H�%���k|��fE�x�=mq0����Vns��{�2����A���T%�n�y�a��{B�{$�M�]�%4xz�fᰵ�g���S�'��q��~���k8���<�x���׷-�_n��=�&��zz\�&�)�׽�	$2-bU��\�^m�ie��pT
���9�L�;jՒw���_4|�\�K��7anZ�(
���M�w��Ej�D�L�e�F�������Ky�����m��0�L
z1�E&ȡ�=¼EB�$��f�3����V{:y�:AK�ն4�C�1�v+���zR�ܫ���-�άI��=�0���vN<",�=�nw���)�Ӓ#����u _kR��:E�pĪ�����Qwu�;E���V�����.��b,�{��G\;�/{}��5��}���M���l�������w�s�K�>�Ǹ##�LH��B�y�슽�u�e2���H��=��Ŭ�Ȼy{�-�D�<�}�{ot!z�4�A�'�.K��pe��e�i�o8�u��O+6���@^�����رLR�Y��<�E���9�?4���Z�˝w9S5p��7�N��� &ʆ��������kۯ������rK��20ǅ�۫����0���������~;~j
/������t��۴o2q��|�.��t��ZOp로|��p=��v�����MK}m�֟gl�\�=�dI<�/yg�c�C{\�rq��d�T^���n��9]��rn�z�����,�v\۽O�x秸1�v���T�ݍn���^��\�570�O�?y�¼�ֵ������c]���pSt���4�ѥb�W��������mH^K��9��ю���4�慚�!_�d�@R�9��U3�-��G��Ѭ�Ε{a��<±�g{G�����<tJ���+�wI�B�U�SO2鯪�E�r��H�/��4w�����so�|.gVp�W$NF`�j�E����,��WNj>R����eK�o�ϴ�L�Mqd����>}�G���w{yʟw\(����9�HFn2??8�N���R�V���{�8
�e��f����>��ؚ{�|(�wPcqyE�����.���{z7�Λ�P�xz��頳1��7F������@�L+�L�W-7���w������j�b���a��"Ѽ�ZB��y�`���y��DB�������Շ}�I �[����la7��~��������/��р��"m������y.-����� �|f�]a�z�^�WUg��gw�ۤ����ˣL�<L�G,�X�u�A�Y��_J��"�y��͛�������k*z�v]�2/���γ��ĩ��?2+�_��'	� �띂�ꍏ@:{��7�T؍�|�z�����Wб֬Q+u�84G+�v����@CTc�4$�|����{�$���}ډ�W���4��u٤<;^"�=��q�����4�_��v�ܩ�|>�q5�g#�����9�Wy�Y�n	Lv_+�ޭ�D2`=�YWל�	�Gۮn&A��zG��t�wgY��,>�x˓�;o=mޓ��פ��?h�i�O�=�յ�.��㠽��Ɏ,�q1�8ڑ�F��h)�"�fm޽�G�+��ulV�����Þ�q��5f�1wz%��1n���>�/�{mb�v�m��E��Ya���c�;��#f�Ol}�%��U�����9���E���&�6��n�u"x�l���/��{W)���no�{_1�x�+������E�9ԥQ���u����_\�������ߥs[˝�<��u�;�`�����[���Hɪ�h�r��[rn�:���3WNs,Z��C|�c��!�>�n�w���(k;�w����^讲��Z=5g<~�@�hzO�{�)b����$�$;�}���;��2�Z��K���.N�Y�w��%�{GjW"x��׎�܁���.���Z�L�� >3x��l:���$B���1�w��t��>��X��"b���9��h�/��G-8����8�u_��=}dy1t�1�ؖ��Nzږ�Uu�Ug,��C#�OJ6z��8I'z$�2;���q�:T#K�"Z�R�ы
�u%G��N��
s67�Ii'|w<u?AW���N�^��y!�Sj���������<%�6�S�v���-�G{��}^�v�y�ڈ�֌�y�K�Z�Aw5أn����y�_��9No+��t��wz1 䙰���)��4}��G^ۜ��E��_bv*�v�4�|j�6���~qo��!�8��f���i�V���W���o�e9����WpCW7z����mvS�ng��[zK�9��ڽ��q��Uݴ���ي<W�u2-�,hP���s�������9�R�"��4/�>�Z}Z�j>kA� r��}����ӋZ��o�M�;ۼb�؞�#8���o�܉���E��}si�y�6��b�.7��M��-Y��]f��j3;��Grs������n&��z��]�N)��?}'�#x͔�����i�0yX���kƢ���Uʫ�,�|�>�����=��	nt��"��{��7����v�����wM�͉>�^�>�	SYh����hT3����y�^^���ezw�O&�J��2�c�OgzM�pCC@��c�u���B�T6�+��gLU�gsa�n���k7�>�OsYGF�z�ރ�ׅ�OCu��I�I(5��=;܆�!�v�rb����!��\k�B�f�f,���.�WC�Wz�ݻR�kܽ�3��h^�.��AЙP��٥,���f��׋�!:C���N?�-�>E�S�r���~�Xק�
�qc�}���[oO^<����V��Ƙ	6��s�<�֞Z��"����:{��Wz�=�=΢�]��VL�<�U=���-�������޽�o��ON�C6ʐ��f�3*T\�~-s���n�7�\��WV+�L��ȭ�d��y=���T{s��9��9�g�N5A~���fš��oo�����K�ॆ���W?w\�̸}��n���˃�3V�,K��-��	�V2V��S+Y�e7��W*�����g<I�G'Z���$�[���h�����t���NwN\�� �W	)rs
�u�h�("����؎���mD�\�q���]/��t�4D�kd�M@L��.�H�VF�"ή�y���j�&���]����7ؽ�6��SF׹���zSxR��=%�X5w��'Ԫ����(�~HLGw�좼~�Y��w�!'��ř�Å��brVN�wͼ~�{y���WL�������>��y�����xw Q'v���=I�������������\y��~�or�v�x��{�9_��׾�u�5��F;�ȳ�� '?x��<{��G�~���T��-�ѯ��}�s�Sc�p���ԣf&��ŗ]RNR�� o�(���y>ʾ����$���1Y���q�݋��q��<;5i��O{�sV���z)q�x˄�x�n���2E|{_p�az7�^p1>������o���P�e�3�s��nF�{;�7;.�����grg.{��L����c��7iY�����Gcr�X�z]���S��C0���aŗ."ȁj�]"G����$�>�ί{���o� 8p������3��im��/I�O�1m�W��\=8[[�쁱�{�z�0g1�����0%K��l��a»b�w{��k0|@U���j��l'�OG�s������s׍��+���7.�9�f���1i�Vq��E�f����=��47��	�Ǎ�ؖ1��}��Ɇ=�;���Χ�yLr�pMZV�nvo���\���$��y���Q�튶�U\�w��0��v6���c!��.�W-xUmy{@��>Y�{v8��V�w��[lj�\��O�խ�C�[o��j�����{�j�w6�*}8����PW��O���54����ל�z�p��/�Y`�\g�˶�ГװZ�m�>W��#�Ōu+��K�qX�Z� Z��ў���u�{���3���B&�`�V��ޘE��mL޽B�;�P��%����ȁi@��\�ӆa���x{�ǝ�ِz}|
	D��FÖ|s|j��x}1,������L����l/����;�ꢡ��EL�6�X��SB+��־)t����ޭ�o8��g}���9��$3�UX���/{�8�;$YB��2ԅ;�2-X� �΁L����hLs��K"�f�J|}Ӝ/�oy�����B6v�'
�L�U1dY�t�#C�]8n��=4*�_�0���'H}�ǒ���զRZ�=��S�uo��w�K��J�ɧCͯ�|���v��S �_g�=c�D�ܐ�X9���/p�җJ�x{���������p�Ȏ�v�n<7�XC�%�6�'��Z�\�m��f��Flyƛ���E��M�j�X�;䧯7�,|���R�|wܞ���xb��F�{c/���;��-j�	�i�^B0]o	���C�����4h�!�c��"�7H�{�g��l�=�dc��=ެ�W�71{��b��".	�wn�k}p���� ��<}�r�����Nҟ���׎yL�ޘ�b��	�{����1�zQ�*�V�
|B���a�5V;[��Cm@�s��:J��a���i/��*N��HY��r���#����������YuǏ:w�jβ0��o�<k��$����C��Z�,��>F���Sq���%��p���\�C<w�{���[rOc�Nb>YN�Oޟ-�H�v��W��T�gfӷ�ݰ��7Է�}����{A��1�N�c�h<�"9�=�2�T��R�پ l��I�,[��am�V��_v�.$07NOx	�6L}݌�o�.1�.��2;������7�m�c�����]\����"�r���Ho{C��/}$SN`�xa/p����ڦ�'�"�\��H�=��q;���v��<�w���	���I����#��K����C̟/8��xU��<h�m��f������^�	�-��3Ôs9�5U�}�ȩy�>��f����;���_R�x��K8;��ۡ4x爝.ܛ�e���rt;�����"�����V�~����(p8z�Y�0���g[i~"�t���Xz\��/dT�U��7�(5���n�ւ(XSx����9��1�{9*����q^�b�9{IO=L����-�2:�.�,[�<��f���]���Fq�d��W/��ߓ��~��|ѡqO
��o������ӳ�����v�V;j�`Z��w�����Y�{b廞穝�w_W,�J^�n����/��9�{}���݈�*T���n�=�c���rY�ý��_�Z��6}����� �·�O�Ε�'���4L��>��<�t�[�)�_�a�pwN���]��������$I$���qq��9ƭ:��\�Ƃn�HW����x�7W������d{���t\�qmqM��譄}(��LODj��׮�J�s{%��h[Z+1��ӎ|S��m�>o4�Z��q�o=5j�Z��Ѫ=�Ok�9�eB��1���M���Du�k��h���+�CpF�����^�۬��Rz���k�=eę%Ӯ{��;=c�K��q�0\�v{mm�
/8��2&�-����cӻ.m��lvw=Bi\��mݦ���ګ�uA�k�����r;�l�^љ����wE����E�v�!�yle��=`�k��,��|t���㭯x�q�b�H���k���0ɧn��#��*�P�F�r��X�n3��tm�3�^����Aot�7/)�&�q�*����{��\��҈>y����|�fŊ��\Nw���k���ԏq�Ň��)�ol�9m�:a���ƣ�ؽ�E��	����e8# '^����W��q���q�+�s�5��X8u��\���m��ӻ����Q��=�m�Ạˎ��Ү�f쳕;:;���.�����75��lj�lI��5Y^�ێ+��wj�8c�
{���w]��7�f7k�}��c�_=��c��=�n9�����N��^��V瓷:u��5�}���}uø�ݔ��r��6�<�3��c���L\ci8Rp�r>n����O�h1����1Y_3��)�+b�o\���*�ݬ:�[�:�9��Oc�+́��q�3�lV��m����X�.9����[���rw]��d훎
�x��;����J�Y�L������s��+���7�N���ڜc���\ݸ��sH^ޣ\��q�䃊� )�������Iv��tu;�m-�vq�m�{��f���9\�lj���q�\k���ۏ&]:n���`����[ݶ�^;n7jA������rK��tX���ԢK�^�X��ΏjIuv�8t�mխ�Ďy{)m��ЧX�C;q��띷od!zN�^Twl^4<���v9w�&�:�W3����u�K\v��{f��u�xM���=1�g\�b��#vK��t��Ǉ4���^��.��GW�2�<:7\�W�Y������8�M����Y7�v�8�Q��j�����9ݕ��	���_Z!=��ku�cX�f�;�kqc��'��� ��pn�㛡x{�},���:�m��{��{1K{e{;���n�A�Ώkh�ܶz�	ّ7�G��t����WӼ�\�n��=��]pn���#������0>2d���[tt�v�#^�f�˞=����2;v���>w8�]�y�Wgu�\�n��=/mU�з:�� ����4k�mXy�7j�ͷl����)�H�{uO���8�I�:�E����=��Iݲ���V+�v%0H����'�;�6�����뇂���1�k��ضyx[�u��pf�\�m�jp�4-�FV0��LFn���v�ޞ�f�����ݹy�=�f�w�7`��P<�gl�c�����!47��r�:�r+yp�#rۮ5l�nͲ�p�zݑ������g��^�Ԃ��XNh'�pk�+Wg�K��޻�qy:�:�\]���f�����@�]��f�{��qm�kxۮ���tN�:Cs�i�g��]xLe�v���ƹR��ȹ9�+�N��y�\��O#%rM����<��e����Vݛ]���R^ۮ:�{6�k[��`x�F�Έ�v�;m�Ek��u�1�������ܼ����c��o8��&��x�J5�<l�3�����{;v W��h�谞3��z����v����K�;<�r�cg��&r�p�4Tmۄ�Pႌ�L�4��E��x�gղ��;��s�m��xX��Z�w-�Ɇ�mBc/�H�k�=��g��Pip+ls�hk�ұ,�g�q�n��9�J:���M J���C�ȯC)Vݘ*Ԩmwkj5����׎Y(��.wZ�,Z�rt�1\���q�%#��6���P�-{�Dd����b����������կdT�Wf3�hs��u�=�;:�`vw�뜏h������+0��u�3�v��fvʝ3�^�ݯBR�{x:��H�v���LDy�۱���Z�9��"���q�c��jk5���
;�Ӝ�nٍ�ptqf�]����i��GKdݵۜ��Y�ˑ��:IS�m��ŀN�!�Vn� �g�`���v�<�<���v�}g�T�Z9WF9:�Oh ]=��ۜE�]�pl�=)gՎF7g�s���l:�+����ǵ������'��軜g�H�� �w�*��8�ٷDN}���y�n7X�[z��k��<�	]� ���p�],�,���ٞ�d�:�s���buתw��T0��;����ۀݷF��f+�θC#E���^ٞ����
z����-Z�OF����շ���"�f;u��==r�v9m��{uN�q�=�-w\��&KY�Ap;r�np'�M��R��j�Ëv�p,I�\g��On�HcC�v�8�ܛ]lTX�s�;�]�a�p�Qf�s�xRT�+�77��Ku����g��nl��ՏZH����s��.�5yE��aS�������l:7��s;��V�<X탌�5n�\��N/]۝��x�mc$A�{q��E�����yre4��FR�s��[v�b�d���>��׆=���e����'L��ܬ$y�+=e�mq�{6�커9�Ku��c��x&n�]v�Od��֞�󋷜g��p��:��t6�k���7d�׊3[<�Ӝu���-����u�`��t�{;��5:�f����Fr�"t8�K��hEۮGYX�h�oq�Mɷllѕy)q����6X�܆�Hn�Q�]��lֺ3t<X�\��\sÓmx���ɝ�vRy2�)�G���=�������F�X}�5�w,���f�d��%�r���|��kH'����.�VK�u���9=i�!��|�yx�V�kX�vY�yƮSǖ�8�!�@�(�kk���
n��v�:�F��7O#��ě�9��B,��7e���r�iȄ����g�9U�nI�.p5be8[�ۣL�юT������1� ��>w=s^��[M��8�r;�������û7�g8���\n;Y�]��mn.����w0=^�(�\��۞�7�<Ly-�;۷\��Z�{d�����j#�%��ruv�������[q���!0���&�={nj��q�ꌧa����F̽y鎧V+�-n{�n��&b�>����>u��후�n�v7{t�����^Ռ���9c]b16��m��η+�۹�9�v㐫�c��sڛE�Ly:-I���n, Ê�t<f�G"ăûS웞7Q�.�v�9JG#��T��m�F�x��U��\�Ѫ:8d�ss�X�{�*�fJ�v�ص���v4��L5��v�s�ϣ��{�/KLA�ְ{sra{2�az�a1I�n5��"�����lHv�nh͹=g�il���o�qt�����h뺯J:뛱�����\[�x7n��w/\��v�q�k�{j�Yx��_[�/,������9ե�6n�Ԋq\�v泞|�ۤ��҆:v�9�gh��;��ƛ�ϵ�ޮ7s;j�Ԝm����-��v�^ݺ���׳H��И�pGm��'��]�Iz�r�F�;b���wq:�3��U���q��,]=�ے�]���<�k�r�v)�^ �NӍ�豊h릛�kRɴ'.�u�콻b��p��k�nsvuӫ�ٻ\�ۙ��m���@u��=Z�v��<Im�+ �M��^��m�Q ]Ԋq*m�m���������dn���]V�9ƪ���lex�;�훷Zŵ��pc�\��o���.ʮ���p�:�+�f�:AzⓌ����hɸ�r̠^[Y��}�<v�����,Rf�r���u�zN.Z�!E�����6e��r�|c��#p\��a;`�퓙�(X��\Wn�!���v�z���[��ډ��y�h�nt��M7/��ݮ�o\�l�t{��n��;kc����a�ݳ�O>ڧm���	ۆ��R�dc��6ɺ�]6s�lut0��u�{[�[����G��f-�k7\a�u�ms�,�va{���Զu;c���;�+�WDc{NuΰN2�WNvCp�[iv����^��m۝���㫭��^Y����N���j�؂S�N/Q�\3���e8��&}���Eb7��/q��;P',u͘��۶w.ݣ�� �ω�]�Վ���l睵�G�W�$1Y��d��<�F��m�z��nں�0F��q�����b, ��NH7Wnۚ6�C9i=m��Iܑ��sm{B��Kk8�ac�znݳ��M��n6��{�vx�{��Svq�2q�p=�*�kE��ӻr��gb|`H�͙%�!�.lݻ3on�Mv�l-�w9��ѳ��=�g���e�n��&��ʝ�W� sÕ��]l���T�g�vW��n��qA�Ey�	rkԆڸ��E �Y��1��Ng����v�,�+��籭G\�M��i�sໝ�]��Vg����=m�Dt�ӑ�c6�\��ӹݚ,e��ήr%䳱�L��<qt��n���{vW��LtG9���n���zw[=i�ku�&�8���=`Q�zL\p�������u�ƈ+	�{m�^.�mj�qq���]�ݹ������p*X�b��^�k*��z�)��^.ٺݔ˦���v-�u��:3�{\����W�ƌh����Y�lrۦ���gFz�rz�{��ƴw&�6�1��Q1r��\v�qs�Aŵ]u�յV���U�n���A8��8��Adʲ|�b�&�h�b��,����TŢ��YY*�#P�C�*�mAU1d��h��UQl�[AjE"5����`��
���L8fb��PF�J�H� ��KiTkV�V���W	U��mAAŘf�H��VE��GX����J��)��Q����Š����fqE"�R�UQj��mA"b���m%fV)�Z��B����J�I�mqef�dF,Qam�E�"�*T���(���E*L2"�Ha��
�m�ȥE+!R,U&-&���h��j-IQ�m�E�� �aq��0�H(*Ņ�T�[h��Ԕn1�$��֍�m�(�F2�ÉmA����-H��1AAX��,\V���$�ɵ.nlGm�.���xl�]u�4�nζ�#TO\�y�c�!�:�۝�d�ζ��ʜ�2�����t���ig`{]ns��M�{n2+ϳ!uv�Ckv�d�`�휝Ş�Y�5�������x�+�s�b9::�;m�G��_8��:�ʬ=gV��p9���������˻v�����A�\g�F{��=�%ڋ��<y��6��9c8���{Gl�G�^˔B�퇏@��͸����O����o&+D=9�Ƿ��60�c�=��Y�A��v��܌��-nM�]��{r�.��=���v^%%������n�����C&�\�'���`ۗ�a���m��su�sv-g�ec�k��u��m��u�vn�26Ԯ����0۹
�y�u��+��YW�$�r���G/:]p6yCu6��i��"imn�&��k<e����#���p��/�3�Œ��3̇A�&UR��Okv8�ֺwb����p�'��f�
�T��y��u��v˰I]��^����A&te���1�sF��I۞r�Ool���e5�;]q�t������`"e��u�;�ۇ9�=���n,BX���\��8|�u�k�睷H��ĲGZ�V�<�Om���u"v�gb���jǧ��;6���=`��&���;q�	�4�.8K��8��"p6�V�t�q�27�cg�ˇ���o��#��o����Ӳ���{{�ŀ:W���G�g;�e}�m�v)�%�F�a걺�!�vx󮘧[�Y��x�p�-ۇvī��4c��z�e>i��T�=t��Bm�k��L�n{��
T�uɜ��:z�ŝKl�>�q@���:��]7l� �U[�!�,rq���n,[�wS�^ϭ�.n6Q�y�Vu�${x�5�t]6h�^mr��a:�:2v�m�v���^N����s��vq2��mFn�ע���w��^(𻰇��n^�l�� yr����|m��v@�.�7��v����ls����q��.��<> �v^7.Dv{d�ϸ��y�۽qy�6�0c<�*'q��N�Ȼg{����=�x�q˄\��q�nݹ|睻�;<#�p�w��9˞�r�����q� �w@�	�q��(s���>r��S�����Ɏ���������3n�|;.���wK��I?n�C��l�D�~w���Aa���z�(�F:���'z�Òr�8$��^��$��8D���=�KԪhZ�����ȓa�TZ��������I�� @�k��3���5W< W���ٽ�F����SdW��J�x*�Nm��׽�H�@�ʆ	�fu����k}�u�ǅ�ۓe�+1�;L�Z�W`�9��G�3��b��}�<��*��I�c�	>�gXp�][�X�� �ES=���FwKgz�#��˽Wk�j��mX��E��WQM S�Rg�y:����@�#���j��O=�z��d�A�c�#��d���sP����׌_ԅ�{��o���'S����S�W�~=�w՞�Lvy�_>$�4��s[��E}��������;�{�����$ij�ݻRx�A#/�$}��'�yۮ����"�}�� <c��:��-c�ߐ�C��i��.l���w�W�cͦ�N޹ _�ge�0?��,���7Vy��J�_���p����?��d�����u]d��z���<0D�*�����DR�v��}��,����+XWo�}=�I>��]�gY�>x��5ߠ�rם�ݱ;q��H$�����&���n��2�����v���ֿ>�����g"���s�~'��ݖ�A��B���~��5��=�|F��]�`�i�&�I�)3={�'��n����P�-�H#�ݗ`�?wN�� �=��X��,�;1�c
�Ri"��E�{kv9ӽ,�A���CW�U��g��BT���+�l��>���4p��:��z�.?]9�2yYr��~�퉫�d�]]9.�]^yj��w�{/O�=3rł~�N��rH���%��h�\�UsYϱ�U�I{�}�޻�}��#{�Ϲ=� $c���&��|�ɪ-Su~Nzi�o���tϽ���&N˿����������w�Qn/onM�H^�[	2A�{/�K��e����V��E�t�H�/]���.���o��u�}I��c���t���	�}�f|uyVG����V7'�{��<5�[n�-5L&]�;���d�ܯٓ�:��z��7� �����>�����m�z�>��~��
OAi"۠�2z������Iڳ��Oȓ���;�'����� �k���>J�(:3V���������޸3�?�� �0�����ܕ�;,��k�e�bq]�˲��Ou+Y�E�۝�h��R���fP��wT�PtD�v�̏1#����Q��KSw�f�Mܞ$	�m��Xǒ?ju�I"�P���^���=~��_�},�o�9u������xT����p��'D�h��%�T�������ӯF�8�aI�k�s���������rK[��]�$�}�Ȅ�z����y=�1��o���� ]�����E�Q�&�1�z_Ǭ��W��y2���t�A?o�XD'���d�jar�G}��`������"Ӧ�eݝ�;"���	�ex�������H$�y�@�}^λ��/J��E�A�`��n�]I�����I�k�$\���$�wO[���GN⶟CV7��@�ji�Vm�#;���s�ś�?xz���O����d�w����y��*�n��E^�N��D�rhٛ��:`���f�4R�҂��K}���q�GC�p�,�v�ز����\e���gC�h�TɲA�T���80:����z�.�Ÿ�8��z������<p��.�w皶�K%�ڣ�<0zf�=\u�1�m�G����Vb�#cV�����C��6N�c��V��';�Ѐ�
a���"�"p�\t;l�%�)���Ǧ㱉捜�z�����ٽ&�nr����uPyMġ�npîaMr��Ν��[���5��c���]u�������wO$�֍a}�~�{>�k� ���Oy����8P���w��\oџ���}�~� l�۲h>E��4�T�]��W�H#ǳ�d�����r$��ݷ`������,�eJm��}���x�ΚU!I�~�g�w��IVyFA���'��8A��m�=�z�/ I^�Zt�n���l�j��+�K�:�� ��I'<�-��뜍^�|��Vu�&^)?�M7B�3��z��w����_��y���.t�� ��]�	`��N7l���o�}�P@�)-8��籺��m��3�℘��!1���j�����o��孅Ɓa�"�p�y�����,�k9�73�Fji_ޞ�b�Ww��~\ǂ>eTLzs��t���?smS�WBMd)�mP>#p�R�&�Ϭ����;�+y:�~�U �̧{Vz��D�`��&V^����� �=��]�I39���%�!�g�`�A�=g�4�T�]Γ�d�f�؁.���z���/*�٤�H�N�� �fs��1�e�(ѣI����b�/vש��~*wt�I�&z�ψ?}����>���y���8+����uPD�I���@��ݐGWAm����'�������A&v���?u{�w���V�w�?�}�]�qqbx�qHE�Y�v�O7<vy6���n����zz�>������q�库>}�vA{�������=I��@���>x+۽w�$Oy��|���b	����0??Pw���f����,�fmi��O�^�]�A�+��/�n�W��9B�A6@�>�7^�]���.���:�f�=�8�+S�N�\��!j���4{��R��d�-�����i�����4�ñn�o�b�	�j%����ٸ~�i
����o���'OH3�zD>�{%�)��~I�L�m������k�tl��*�'��#+�˲A f����8�����>��񒐪T�P{���<����yW����?z�	"��'�~�ge�'�^�v�"�������[�#�l$�Sp]xSq�A<�����o��޹Zݴ �]�~�ߜ���m0�����3�D~��ݖ,�H{�����㏱mIX��G�}u��c�e���U�e�������X�U=����؁���ܻ��K�w����|gնed~�J��@U⵴9�,U(��=��v@$���K `�}�j �	�^=������^��d�?�9@�A6P��nW"ԯ�
)^1����~x�৵�b\:�״�x���J�ގ�x:��t委A�mG�M��ܕ��yH�w�O*S�T��S���9'�W���fj�_���х6��G�`�����]݂E3�u��aS*�u~~�7�I�����;[>�� ���e�=[�K�A��s垕��pz�V�z;4�J�&i�H��G�۵Zb|�`��s�ד��r��v@�+q��������ES)/w]�I����8t�M$�������N�`��{�febzA%:,ܳ���?<�^�]��n�VOO�~l���������z�_���� �,����H�-Ц�/�vA5��~$���I��j7;F�G���,���8�����n%�bM��o[��e���|�{,�}�f	[�/�_�����	��w��@4lPA6P�[���u��T��n��vzY?� $z��vr-{���eW����yv�u���f���m���N�*�߹�P�T�������S>�c���ι^�0_[�o����5iI���cs�,5����0�=��8�s��u���G�v]�z�cGk����s���M5�;x{'P{n�:�Nr��6��`w�[c���9�^��6�5���Rܷ6�%�v��í��k�=6��On�n�����Y���^v�'�v���y��O��n�9�&�)�j��c��#sǡ����rnL=�	4��Ok���i�C�5�Q;N흴Qˁ��]a��tXˮ� &�d�b��<�~)�n�iV~�՝w`�K�;��G�}�`ϥ���w�zi$���#Hr �|�(��RP��v7�7�k�UW#�w��$m՘Oď^�n�'�逐�ӱ���{���1��tC�z�B$�^�X�	����䳝/'�%��A �[��>��]�%�ο*%E��;;�^�3���o� #��l 3�{ߘ�Y��yS���U��4���b�*��̛��@>��Auv�:vA �o�d�};���P�o�|0<��S�q���x���Yn�{i��v�	pw�iRm4�=��/
&��=ڄ�I���� �wzY�s���}�.W������>+H1��*jJ����Wco�Oj����G�߶����-�˽����xǺA{Ғڛ	�����"���2z�&��ra��G���+9S�~Dg����d�OI9�t$v�L�&�K�	'칽w�$Ww����Vc��P�{ޮ���A��6�UH���7�������$�l�{�{i���=���,�}[ނ��@��ĚtC%�ٕ]J������oX�r�lY��O���,���l{{�T�+4h%Nλ$K$??&J�æi� Y�������z[��/ߒ�V~��}+{�d�O��]@ue��bn6G�����wό[S�qrw	u��@v���Qg�wZ�E=���[�=��<�*�"�x�n�~>����I�\�xw�����5��A��Ww��$Z�$O�+�M�T*{jx;��ђW��ɂ�ewzY$��5�0 �`ܞ����� ��k"�M$��՞��%�]@O�_B;�z�M]���G��էFR�4\&�|"�B���/��9�Bپ�¾���±S���̽;�o��8�~XY����GEK��h�!�5v��8����#w���[��g(s��l���Jj{鮟�f��k�5�!�l��E����ȼ�rҶ5���/�5������N����ۦz�Ԡ������r�O��(��Dս=잽�ߟnHɩ!�؍���S�rΙ���{�u�?]��ͼp��͹���a�K�/,�{|��0=X�}�9;�/s3�v�{�
���j�0��q�IݳiwY�^�p�����n5q��0@ꂗ�i��Q r�B����RbйU�i�7Tdp���zNP�["���i�������Dfy��͗�k�7
D�9�w9U4�!���L��u.���!Ki�1�֨e+�ܼSv>�
�K=��>�\WgOn���x��9� ,/�I��I�o������kn_{����,��=��O,��j�;�w��Z�i���Q��˱�;_oQ���V3�����j8x���K�	R9�;����0眳�{��z�^nv/,5`�E;IP���C��)����2빃�U���p��2'e7g��v�HҮ��-=}�}k�f�U�_�?^!��rַ�c[��w^՗C��=���[�u��j� AF�x�PwӵR
k*ՠ\U|!�����=^�OK&[���/Y�v��;�#�1;��>@N���y���7;��矴Wi�Ub�QX��*T�mPmP��X�B���������ZX�A�C�mqje��aU�,m����VE �ZR�U�*����F.�-h���2a�2��[[�TkQ�jZت���
�eIR��űbR�b�#kIiJ��������k�-1��ZɆ`Cc%`�U�-��+l�\RT�T��V,+WEb"��k.�ʪ�ekXTZ�1h�H�F)��UZ����m��0��k��"LZ��R��k��6��V4���cF¢�elUK�1V��h�
�����A�R�R��Ķ

J�--��jV�ҋ[YiB�QV)Qp�	AR�F���k�J�hԢ�FE��*���E�5(�E��
"�6�1mB�R��P�Z��X8��o}�����[PH/��DCȃ���U"��ew�׽℻���'�ۛ���_����}'s2��Vvl)�">��ƚN�
6��"�Qd�v���$�����<����{��}/�A6�A=:�vc\��{�����q���!g�y؁|���:iLX1�Tn7�E�T�������?�x��̛���g]�H$��H'�GN�]�/��+F�s��H/}u
�8�����H�����ܰU��}�bw�z���>'�~%��$�N�]�vfj�x��
ٷ�sR$2U�e"�J׵$��~�$Uf=�ɕ�����P�O�6�v
��?R4�I*�����u3��M��7?~����$^]��:��gJ�-�1��;T��n*�8�D��G1w�͔f#�m�Λw`���6cn�����wf��)]�DX:��':���\|	4������e�N�I@gl��6��,�/�]>�V�s͂I�~���>6=�"�xOW���b�?*k�>=��X�&L<<�$M�Svk@y�]=�\lZ��F�t }��&�ʒo<f�O� �����$���]�g�L�E�J,��gT �N�|ڈR����B("iMIY/y���;����Wd����/�~���	C��N�jn�Pߖ��YZ�MU�]��d�g�ޗ�?��^�/����?�tλ=�뿉�.�D���L�i���}4yq��}wb�$D��X�� ��vrh׽CI�|�wvHO��}��n�2��]�۲;9��e���U�FO��r���{��?��|��:�#�0�ǜ�Z��Ս{*YK��pmǵ*2U�\��%��yΕ8h�]?f���8��'�u~M{}���V�˰�r{W9a뤛�M^�9���srI��\��G��m�v�g'7�����Hv68�K�6�qB��qok��e����sz��ѡ����	��j��=�a3�6��;/g��8�@�e����n��9;`��dA{]rj2���[t��k=�8�I���.�7���'/���;��{�o� ��b퍍z\]G5���Oi;9L�M��8	�iܮ퍺���nɜgi�5ܗD|��y�%q�B�c����J�{L��dLQN�W�J�E�QdS�R_��Y�df�,�#gU�0�Eb�;ݍ���߼��=��`=��|@(a�o���@y�!�/������'I��>o��~#g;���{=���=����j�,�XAR	�Tу]�������$�Īț7R{;�q��A���/�A ��f|����A��j�ϳv�q�ת��"N������$}Y�f|I�K���u�Y$����g"H,,
�F�J��|�'�u���Oo>��/5T	�����>8>^���f���?�?}�-�\�=nm=X�q�U��vS� ��5��������W��-:t�T��{n�Eo;�O��������%�n�uI`A��q��*�MQ�������Ñf���Z�z�Q��ylͣ�7 uo����k�3_ �>� ����3Z��>��g7��_t�>�C��2���A�5���A�u���yp*��l��믑*�F�R����$����IZ�=D{[���l�	o7-�|�y�:PQ�UI�o<���~�Q^ -� ���|�V���	^o�c��� �c�^3	z[�Ъ ���������<�T��=��u �{�|; ��x0|����+��:���|ߝm��p�L(GIn3Y=���Z����5��
�uf�e�����~vݿnt�b���~0�_��?	�{���,Il����8~����HO�Z�iӤJ�v��ݒCCÅg�����t�����$��K��훾��9�Q��(|J��STj�i@T������A>#��]��E1��uk���2�:g8���&:}���nn8�N�y�(�7����*�	w�A���ۇ7���.&�Y��u��~y�۲A��z_���pؾ @�F�,������Ӑ��ٗd�?
��]�I ���۷�q�Z��"��.�$]�Y�0��)�T��M��I���ܯ��gu�Y$���� ;�_|M,����j^�-�JӺV���2`��Vꂞ�hvnl�\vwl�U�&�N��}�_�t
DU�;۷vA ��z'�o}V`<�SE��d��������l�a�d���
!�w�8�"J�_E��.\�ͻ��o?jH)?x��T�����t��Cl�R
�{���$�����y�R��wox\���K�����Eׁ\�U:�ç>��>��vA�a #(�YY+���h�d�IP�J����߻����9q�z�y�aF�罣i8�d�������5&���V�^��:4P2 �B?�w���,��W���nv����D|@߳���*Aw���T؁R,ӳ��a�~����5[n���/ĦfU��}T�k(U���zNы�~������Az���yC�!���w [ �xL��=���Us������>��d�T=�}��!ĕ���}K�q*�r��70�
������$�T�
�߷ϴpg=���{���|�Ĩ�o��q�Xk�]��<���O�?�y�|,��]yx/���T�T)�n�:^� ��`�O�s��=�"�\��<knۧg�VhL������)sL�˛{��c���8�++%ed����F�0��*IXY߷�na��8c_��~�?C�(��{Gr!Y++%eu�皓ba������.s������? �#�{S����wW�o�S}�R�!Z0+M{�sp*l@���o��8�� ��l�0k�cX�?ҽ���8��?_����m2�)$o?��0��%��;�{P�AH(�����}u���|m�V��]{��l1H)��|��Ă�t~�1�78�L�5i�Og�sG?w�����^��@�7++%{ϳ�d�%B��)���8Ì*A@�;�h�MW���2a����;��� �~D��E���4�~���6��������m �s�}����q���!� ���k��SbJ�Yb}���C��%ed�X���}��q"?	�Z�z�v�g��Th�ο�-ʷ��B��a�%wb �<�YI�/�h�����'��������V�'�;�_
�9�:���QtiSTApv��۴Æ���s��vE+��Y�OEٷn6�͊
���+���>���n}�y���i��הN�"Ǜ��������v�����Ga{{`[��e�q&y�i��%f{�X`��_>ۥݻ��7K��;@�9��z� ���Z��V��e�at �rn6m��nG����c�T��w	�[�����͑���v�������=r�i���σͻ�	�>oF�K��&�l��w���:�Ur��?���a_߻���0�RX�a����9�J2����F�8����ߍm�ƿ{��P7�A��a�����
ٮG/��nnWsn�T�O���G82V;�~��u�n��g�u�~�4|Ʉ*J�V�w��a��T�&��}���������2�x�ߧ�~=��U�t��2 zb���i�.m΍�p���sP��HR�7�{�7��*Ak����.}�?a�������,@��s��3�����o���6����z_��2g6�N���?����] ��nQ��Sw�f��>ID*J�a�����3����@���}���Xkƽ�������r�_>��t��ua���5$��ݶ�[�s�����p8�}�oF�
AH/w�y�;�ps��[��a�+�k�0�
��w�Ѵ�B�Q� �����6�@��߻��5�}���}����k.���{CV�z:��kU�t�wmrm�'���3�/�V�w�����_� �����y+�_wA��F���}�|
BҐ�`V��k��T��7��ޏ����?�xO���P�8�YFJ�C}����q%aNd�K�?2�SŻ�pa^�����0�K�8h�w���w���e:�!��o��[ĭ���".s�Y�?W��~C��Mk�[tw_'��N{7���Ór`�Y0�ӻ���G�*�I�Fg��+��ҦF~���ppg+*�S}�}���X5�`׻�?�a�A�!c��q�|��\���a��<�>{��~tt\g8�ͻ�P>�5�H,���_w?�l0�IP�+k�ט߳�l�7����� �����h�AH,�eu����x�߰S9Zfg-��$���~���{ٗ%?A�|	.���v��B���}�ہSh*a���6���~����;H�C%B�����C�%aL���y�9˗4����a�Ϲ�����(!Xs��pg���><b���vuIP3ϻ�@���Z��]{������l=��ڇ3�~ғ�߷?8�_"���"�!Q����KV��
λm�jIM]��U4p�99�/����L~�crc8���������R(�]}��ѸɄ*J�V��=�q��5�j]~�����M���{GpB�Xʐ]~�?�&�aw�v�W9��2\�@�V��ClH{�=�g����[��}�*AH-5��p*n T��Ow~��q �����>޳����xʙu�{�Ad#�~e�.�j���Ì80�>�~�la����X{����3��P(�XL������> �Ĺ����3s�-a5[�����{ꔈ�މu.�[�>��p�P+O�ݫ4��1�3C�")�s�߷�u�J��X�y��ځ��e!ia����C���v쫌�����p*lI���h�s��c>L�u���:Ό� �ﳽd�IP�+���ۇq�aF%}�h�Mc��w��d�eH.w��Rl���eɜ4��K�@���}��G�!K@�{�h�
B��s�]l��
�=�����+*{��ڇ9�D���@�G��=��o���v����͇�6�&�Ϸ5Z7h��/�]s����e�{!
gu��q�jw��~�,S��G��ow�a_�����$�B��V�}�Gq���*��}�h����,��o��01���ځ��JB����O�� �*���i���b�:��#&;﹣��@���)�����"���|Ʉ,IP�+��}�m�VaRT���q �ped����w��97�9W]>��2 B?���j�R3[0���7��� �F�-�o��/G���&�I��3�5_�S��|>@�D
����چ��J��P��{�H,8s?�?c��\Z������G7հ��Ε�J���#��B�����q�H){�Ѵ	R���皁���)�ٽ���𨇗A_��´[4�x+o&`"��<��>�	���'=�'��T^���.�'�����)|���Y���	o9���똿Ą�� ���o�jy�����j�90g&m�
��5��O�*Ae+��<Ѱd������Y��)���~�6��
°�*o�{�I�
�ded�+���jM�?w]�o:�`/���@&�D�t�Ȣ[$4��.�nٺތ����Z���]�N_Ͻ����\<t�@�V�{��px��H(����!m!Z���}�7��
�����]׽����z���wP�8�R
߽�h�IXSx=����npf�77p��w���a%�&;��~���Xw[��Cl�2�T����@�J��R���j�H4�.;h۷�}Y���~y��:~��4X�K3���q�߷�i�@��d���y�ĕ
��׳�g�p��绯݇taXV%M����$����VW��y�6&)�xi���ܹ�0a�� m+��{@��z��|k�����-������R�������7*X�YD�sڇ������	�3��f�*C�s�h����3���5L4�70�¼����la��T��߿s�83������m���a*����8�ȕ�cX����@�)����{���8�VI�����*?�8���۵"�O��u&�7V�5�te��b���9ݏd�4��W�TxJ9W��Q�.���=��>�C�z{n]�%`kx�P��w�t�sK�^-]Μ��'�^SxOo�Ӂ�n�ؚ�Y�{�\R{�O3���38ԕ�!���<_G��_�wd#�5���X�Un��n���} ���@���2��;؉/�m
(���=����:���U�z��"߿C#n;g�?�j��!�g�:�n��l���|��H�ͅh�=&$�����h��6ы�Wssm�5OGV��==%�;R������k����{�P��Y��n��?[�\�l{��H��T��v@G�_{n;�Am^#���+�0����s�]]�ũ*�l^�aVg9+�<Y/W��m��އ�'������0M�؄���jz*]uӗ�{�	�x�g���Z{6��hz���b�|������ސ���B���}dX�F������9=�֨_t&�-�(�S�'�;����w����~K�t����}f�� �.��w5�=]Կf������~�u��m��5����u�>>��c$�p�Ԥ��/{"�P��w;�.���Ycg�<���]Af����M:}�N}
j��4�!�=/&W���\�T��+~��W�{td�u˜-������{�]cà��Zh�)�]���dՅ��g�C��2Z,�O[~��1t��� }���/hF=Y�3Iˇ�6Ja��?��^aw�]�/|rJ����%j�
�Z6�j��"Ae����"�Z QZ���ʕ
�$(��\�V�-e��V�
$����R�"�j4�cF�0�bŘaP��kh�Y���fT�j)U����1JTU���VV�p�
��c��-mKhV�j�-��+��pJȦ*WE0����
��m�F�`[Q�h�(��1��F�b2��������0+mbі�UVZ�Qn(`p0QeR���Z��
�[FJ[YXYm�j��\V[kEeJ"���#ZԬ*6��PZхA��ZŶ�V���V�Kk�QEPQp�b��XQ�l1KW�06�UjV���ËQ�������,��V,Z[X)jR�Jȱ`��X����µ1�)���J�ZEmZ�b���5���V�Q��
��ae����eV-T��\e��d�sۄ�ys�r.-]\���t���v1	W�e̹�ݒ��M�����!Mճ^�cn;E���ٔ�q�;s�h�Ƌ�V��yB�E������k*���ۊ�k�iM�7��M0swY;m��z�#Üy㮘y��.��vL>��_i����1�h�u糷Zֺ�9�n�����H��y�����H����plî���v�0��⺷�n��ۀ���a�+�i����ZkXTJk8{Y,�`���4�֗Z�ڷf�ۗrt��2`�W ��˷8��!�玌SNq�,ִ݃���v�K���;=[S9�1�����eA<��n���ع�	�rwm��q�\WQt�c:�<���[5�\����gy,]�ng랷@K��˃��m�Hx���:�%�rq�Wvr��8^^7h�<\Ė�w��Hq�きk:)���sc���4����8����N��=�f��k�����mحt󶴰�����vگ]8�ŋ>:�O<q��݄,�n�r98�T�\�_=��SѺ�5��ѻ=�b��C��.���p\=���iȕ�u3p>�V68������f#�+�%���y��-d�y��cm�qŉ ���'�������h�G��<v�k�t�7�kNN�p��2]ڭ����;��t�u���4���q�e�n�m&o��%�Y��'xԜlb�>ܛc#�׃��^K�p��tz2&�ع{;�t;��A��a}*��x�ۙ�Z�����o��v��x#����t�[Rj����a��<���<�nG3�ǝ=��ےZTɮ�-�kmg��+������e-�G��F���THt�[�e3Mݣq؋���Xgl��wc��v��
{�Z�5j��xP���m�Rd���ɂ�z������i9ړQ�Z��zf3s��9�V@6���d��]�iϴ�|�W��3��sНm�`��ۭ�Qƫ�-�p�0uDf�kV煄�Z�'��	�N�o����g_�r�Dݽq1��Gk!ڑ��$ι�$���p��u��K�ݷ�#�����Z���v��B�uv�p�թ�n����ު��pC��q��m���j뻭Qn�w;��YiDq�n��v/c����]>�f\�Ş�VM���i�\l��<t���j�tS��K�vf�Y;h6���h��9;yWQ�ی�vN[���a����ȕ���3�!�`s��	3�s�oo.0"��;�	����=��W=���yj�90g&m�*�&9��G��2VX�^��T6���~�$��oO��v�I������$��H,�eo��T�y��g9�n��\��Aa�k��>x��Rw5p�-�k�e��Jނ��#�H���u�������=�m �2�+�C�L���oA�>�=�{�'K����.nn�Xla_k��P*M�Rw�=�m ���q��u�\k����X5 �o��P7R)Kv���Ç�N{�h&4Sl:5U�`�������so��u��ܾ��+,+���tld�IP�%a����+T������o��o�sS��4�FVJ��|��I�0���i���nZ�˝@�J�}���px����A g{����_�y�8{�n��r������op*m�X���{P�Ag*!���q$�?oG{���������������0ُ�Oeg� �":*�5vf�%��d�1��&�_�߸�~���c.OC�0�}����AIb��s���q�������H,��mW��oq�Q����-��)�?{��P���Zg�z�k��r`�L۸7c_w�8�*Ag폛�_��m��ڗ�~���¤�;��pLS�:�^�������}�f�QXfY����@���҂���s돞R�d���]����s���O�6�z�u����bJ��w���ĂÌ*K������8�d���c�w���{��za��y�6&1�}�9�[p��es�h����4�jB���{F�)
�yΟ��>]{�޳�
��*e���ڇ�J�P��;�C�+9����qK������Ϲ�����~���|�(T�B��~��8�2XʁA*>�=�@�J��X����P=����G=ۛ���Xg���Co�S��@���lҪ�� ߫n#��YY+,d���y�`Ʉ3���~���)�����m�XV�IS��}��8!Y(��Y]���T�o]ϿuG��w��5���7�-����h:�q�{v��&�e��o2�#��˶-٭�����c��5���=0�Xk|��<`Q�h}�{F�H[)
����{�nM�T�4g����9{�gS?���g+(�P�w���!ĕ��֭��[S-.MCl9W�����T��T����3{�o�5���{���ǪJ�N��{g�R�w<��l�.�魹Grg¿{�>t�EU����Y5T��p*lc_��N VPd�����s�@�m%B�+ٻ������{��tw�sw������	����������O��W�>�2���<���(���ъw0�Wb�N]Al<5��?f�_s���s�������aXV����Ѵ���ed�+�w��bm���U4�-W�MX� �B?
���%*kx�[������=���H<)
�l�}�@�n T��YS]���8�I�{���Ϝc>uΐ�I�����l��x����q] _��!�A�����I�{ʿZ�o��� �D �=�@���Z��w��077H6�H/����|0��}��ǟ�[5���������e�9V:��豌�+��v�q�����4��,�f��,p������~#�������YY+,d���3Hn$���{��6Ì+���g��8�o���8�������߾�d�&�.����Wj���$���P�AH~Ͻ����ַ���y��-�+`����j�h �����3���*�����{���g���m��k�p�As��|�i*%B��=���8�FT����Sfu�9���w�������Xk����ٺA�������jynu��Ss���I_�"/�>s��#;�p��k�h����J����&��hQ%B�+Ϲ�na���*J'��}��|_����z�-�fDMab;1`c�_��U|礻�W�ߊ�twE�$�P(�Y��y߶�Ϲ��^�.����
g����>��sZ�� ଟ̬�2�����I�����}�g-���es��������<`Q�-�����!u��|ǽ���9�<`V�{����
�Ybs�9�C���YY*C��}��pIO�ҥ�_�@k�~�D�E4�e���:�r������+6����F�v��l��{/���??w\72�9Ź��+��ϴID*J�a�����2VT
	P/y��g|Ϟ������{�`y�>�{�1H6R�߹��H/1�|W��b��q���=�}�H,�d��>�>��x�������߳���B��T����s�na��aXTs�����B�VVM~���8�h��׽�k��Rn&.����Ǘ�r�f6����=��Ă���}ϻ��!iHT���x��6x�����O�*eO��}�q�d���
{��q	+7���P�!R+����~Jg��z���Y�q�>Ib%�5���g,eH(�>��q�X���5����)�ԅa����Cony�����9Ƀ93n�T���H)�2W^�y�c&�7\���?�����ξ��Ă�Rr'���Gq
�YH�=����#��W���L���ݲ̞}^ �3��y��nz�rr�q�o��T����<sӎ�^y���Y{�ٹk%Heo�t6uއ����~}>��7k6t�f�b�з���]{��E�s��k���n�1յ�Ϲ�2���C\��a�FN91xō���n�����i��l����Lc��[F�m�v���k/T�`�;�vq�����j���z5���=:ӌ��:N�%�*�7+��:-uk�MpS7\Sc�Z���t�ړ!�/k�`\k��v�v{�*�ssd�Zz	]
�nY�N�v��5U���\��m�gmζv&�g��~}����k�z�������v+�}惏�h��{F�H[HV�+��<�
��Ll�}ۿ���e�=�oP�<2VQ��P����C�JÔ�~K��&m��-Π��0�}�����	*#���&��s�3��e���sG��J2�Q*�߻�@���Z������P71H4�.;���sy��=���P�An}Ҧ3qq��5i����$��2W���h�d�IP�J�9�g�1���c�k��=�m��aP=�����NFVJ�;��RlL ]��ݦ:�(����X_�?@ޣn�ߍ*���Q@{vH<�+Fo?{\�
�*Q�"=�������3����W��=���}DAB�{Z�tq ��o'�����ٓMÉ����FH)��s����d����Φ�6���}�hJ��RϽ�jH;�-����ǀ�>�+Žq�Qt)�����R<�ѷn'��M����]{GoiW6(�r�__������g����*y&�����ȁYc%eJ���4m�X��RV;�sۇpaX{{���x�a������h�NA
�FVK^{��T��߳�d�\\̮vq�X{���<`V�=�r�޺�;6	0��l�?b�����4[�nB܃G
"�{�^[�eH�w�j�5����0,�t�ӎi��/�$��޻���H[HV�+g=�sp*AM�e��9��q�+,*����[�i��|oyޏ��%a���Ɍ73k��\��+�s?jI�
��Xs������~�q�k��m����N�~�Xk�y���P*A�HV�9�Co#���L?"f�h%p������v��;x��J���82VQ����0�T*J���=�m� �}�w�6��z�\�n��~eH.��;ԛ���y[��Q�*g;*Aa���h>0+R	 nw�Ax��}��ۻ����Qd�5����
�YS���jg#%ed����Ad|����V�gg������]�i^�ѳ�k�	�{,'��$u���f��@e�������a\Vd���� ����A�T*Aa���u�q��@���m�X���s�����~�Aw9�|b�iHZXw��<��LmL�q\�ͻ�P3�{�O��R3���>���1�O����B�*%aO}�{p�0�(¤�>�{�H,�Y>�^�9������=�?	�1󿽋��\�L���=���0+R
y�{F�R�����^q=�'����\̈́�wZ�e�{}��
���v�a�+��qH��.��S�T1�M�ؼ������ �o��'�*a������pd���
����q$�(k��	Ф���_����~��: �=�����i'*J�a���r3����P,�=�l�"Vk�y�w���<?c�f�dJB�w���ǌ
�=�`��%�s\��;�~ލ��e+(�^~�y�c&P��S�/_�P����߾����aXX w��m'+%eH/;��Rn&P1�#���y)?v];����d��4js�8�3�b;:;�G��7��g�;�C{o������v©��P<����wAǌ
Ԃ���w�7�H[HT�ӝ�y�M�
���w���{��� ��w~��C��%e*!�=�h�IXSy��p��&��pa_�c��n0�J!R~�k_?�����=�3��2�Q*y��F�8%`XԂ��5	e!OO��~��߄]�|0��<+=�/���L۸7k?w�8�@� ��;�2��
����o��1��߱�a���°�
��~����$���ed����w��i�1��1�&�(U� ��~�� ���<X�k�HRZ���h�����[���nbH,�w��ڇ�a�>�����u˃Y�uU{�U	�Z���q��)�o#�v��W�MMP��y{:��]qHN{��3��/2?o{�Y���u�ܟc���O��*����q$�9~簎����k������}����%�V��jdϏ����r~@�%@��}���
5�F��=�@�A�!m����>s��ݖ+�;��w*��$AN��̺��o>4Â0ݫs�v�\s0�ng���yz����G�*��%���4�<�n#�@��%H.�c�ѶL�D�
���������+�w����C�����8��
�YY(����5&����Q�
=�qs�@�V�������!���~�~L�3��g���!m!Z��׻�nM�
�@��w�sڇ�d����������o����|���+�̘2ja�
����A��T*J!X{�9�g+*�g��{�Ѱ���?������V�\��jH;)l=�sڇFsϽL�2�-�G7P0�I�y�h�}�gGg�}�o���:�̕�2W�k<�
�P�J��wp�F�T�&�}�h�M��_3�j��,�Y++߱�ړbew�˓�ٓ:6�Ĭ;�sP�AHp���{F�R�?v��}�g�:�`V��~��a6 T������3������mB>G�b�����ZT��	�_dߝ^�yŲ�D0�������r�Y��%>�l�{O?Ʒ0�ܞ�]G�2��*��#Wu2uڬ�����}�_$�qp��Z6�q;n�B�۶k�t���G7g��n-O-�ֵ�wt�ټIXNۡ�c<А,2<r�]��`nYڑ�n{
;�Gm��'��WOnC�lk��;t�=�ḋw]�d��=cVz�V�&Rt΋"ۉ�a��	�ǋ9��,�Mٍ�Wyu��ϴ�iz�l���|e�|9p�����g�WH�}e��v�Gcu�kS��ȫp�b�S�<�pqt��=m��{hCg#��,�ș;1�9�����ݞ��s׻0�+��ϴe%�T�
����tq�d�ʁD���q�X?Wgj�Y��4�����]!�)�?ۙ�Ci�4~<�)�q���]��r$�;�h�AH,��_p�ui�}��']}��G�&P�*Aa���چ�paR
J������8�H,�kϻ��γ�w>ž�o��5'(o�x)��-�s�@�V��
B��o��o��H)}��q�]f��Ͽ@�|�R�VT��9���q���T(��}�h�V�W��Tp�WMÉ���������o��`��B��5�h�8�P(�{�Ѵ	X�
5�_�|���b'�;���||_���|q���3�}L�2���Gp0�}�s�8�@����2W>�h�&P���Cx���{���?~u�C䕇�s���°�*���Ѵ�������z��� m�5�&7�~�\*��Bh6�ܗ+��2��c���Eڶ�ڮ���v�%��6����=�p���m�dύ�y+߷�h8�Z��h�}��!m!Z��+�쿀d|	_�w��� ��|EM�3�%e*s���!�%aNc���q�4��gpXn0���}���(�|@D}�ߊ�<z\�����=�Z�>�u������s����}�M�rN��S��v�7O�*��@�{ý�3�8n��W�N^_�7d�ʕm�����}�_%�Ea�{����JʁR�_�����8�Ĭ
5�Z��ځR�!{���8��~�����i���8x��]Ql�]@�q'=�sG��++%s���F�0�IP�+~�ﶝ�w������a���P9�}�I�+%ed��{���77�˼U닆ֹؤ�'�~�L�*�<MUW���x�>	 9��F�)
�Z0+f~���
�@�P+(��9�C�u�����{[������,�D@}��a�tO˩ X&�F��{?;��O��K��{Bu���U��zt���<� ~'�/�g}㞷�w���zl2ÉQ�Ɲ�H��m<�	��{M�K��X���V��_"�u�Pc��E�U@��:d����wm�>=��^��/�Rd��y�{e ]oh��E@T*Tڎ�o�:k��eq�<���L�=զ|#�/�,���Y�j�W�Z���J�M*%)��Om�� �~�Yd̮c��rQ;��n�j>�¼y�^g�w������Z�E�PE��ʡ�9���UW�o75���y[�0/�]|�ba��:�M�D�/x\�i�d3�NW�۬�����.mqh��C��{.�)��;��y-x��m���/��vo���LWe�QX�{��6��Ce���޸w.rl�n!���^�E��/�pxsuy.�Q$���8�������5��O����J걨)��|	����žn�^���������}�Y�o���9�������c��d:��<�ǧ�{EP���+ȑ�`�{�UN�Ne0��>ˣ����۞B�Pg"=������v��R	�y���� ��G-�<o��t{w�ߣJ?+�E���d���X/�{�>�~'wqz��o}x�a�^Cc[�m��������N��د�)�ݑq?Q��x%��]���#�:���	��˲���њv��F<�Jo�Q{���;�\�_U�C��w�K7�!��.`����	�j9,��P�䧗�~~�%���DlB}�����Ì{<8#�sEnv�&���{b���si7���3��{��|�0���[��!�[���X}��g��y�Zܠ�ksG��bB��޹J��rUW\ׇs����4��P�ҒJ���'BmY��m���^�te��>�.>po%�w*{���;��M�K5��^���.�<��ckO��\{�v��U�oQ��A��B��y��i�����Sh~0У��������k�ET0��Z�JZ���-����V�1hŮ,�(�#�a��bʈ¥Z�-��RW��m��ʶ��"���"��k��F�+��m�ea�h�Y��T*Pb�Eml�TQ��+qq���m�k*V�km��cZ�qp8ţDU�m��KjU-���QR�V�R��TV���U�����E)eER�KJ��j�*&�0��V����U05EE��*R��Җ�[T�)�U�R#$J��V�j%�cF�J,E1lL1eU"0Um���ѩF��V8��X�Jؠ����lU�UG	m��QAUW1m�(T�J���[V-j%���²��KkkVPZ���iK)R�lD0�X����%h6Ո֑��*��[h�*1ũ�)QF�Q��"Qi`��[�W�m���7	�U_� @o�����:���=����7��2�&SR�+�s	�����	B~;J�B̛�	��X}����}=�@=j���bd�3I�؀�Otw��e_�9���PE��� {ѿ�-��؋���T�h埑�f��4f�v��Aً>YvWFT
h�d��-��V�]�5�'�y�@��6��=�n~#�;/� �H�v�Ʈ1{SV�W�`�H���`�W�ň(�LS�� ���x��0���,�	$vOe���v�_Ē:uY�^�F���0��b�N�,���y���A�����${`���خ^)�i#�/�`�}ݾ�v�����(4�*ו�^��͒g H5�o�Y$��{}w�$`�}(�%��)��p~_��x�	�s�?�Oٵk�G���m܂�:�t��M��&������US�"u��KV��-���N� ͩ��ﾃA7^��?�Y��p�`����y��}�6�5��U������d���]�A&j������r�&���İ�J�(��������Ԇ����Z��`�9kr��{��;��j���fL��$��o��A'鯱@�{g�(|��_�� ��(�Q87�IXؐ�����U��~ݓz~�y�dFw��`���k�����4�z�e�����b
�:%%N�� \m�T}���s����]�Q�����Ӵa�GB�w�
�[��[�,��Io<h�����5��H����8�ު�c��/3��^�|�)�*�b��_9� �~����$g��X�������G��@�H����;����]�C��8��ٓH�Yt9윥D]��X�hb�����,��Ÿ��옥d���"n�{��wϯ��=��}����}~�v��m�7>���5� ��v�7�=>�M�W8t[n.y̋�73<�2��J�up�N��vΕ�˚y�[�^;�"Ïn�7u��3��S��]LF�.;x��{Y������X��"��ձ��s��\�nv���2�m��]Z�OA�l�\N��5��I�nv�[��\�:�ۉ�>����]u��v�x��w;ۛ�s�np��ڠW5�i�v�v9-hw�@<���z�n8S��a�ιԉ �7��~{�8������}����?G;%?{e���f�X�Ϟoh����Iw����qd6���龱g����~B�k����el�H�M,�p�O�_�������wy���5�8hl�=����2�]�9�>C0�����wj�����e����`����/�.�H��%���)(�w��pgysx�I�+ �I�{b�>�������ݛ>K1��+4������6���I�{}�2X׵ZK�0�P'�U#����d��oo�����'}��}]��C����N�����b.�3a�4Q�.�ۮŴ�V��~����톱�]�X��2 �K �H�����V�����ȳ�`�u_K�3�,��%@���_�M���\��7tz��Kz)6W�Z�,]mǈ4g���6^w�vK{n�*��ՏI��zz�������N^e�c!�z����M�ş��}�_+�[?2H$۝vA���`����nb=K7����&�|�ջ=������d�Iښo���=�ߕ�I$��nu�$��벘<w$�*��r���M,��k/��3�]O���tH5��qV|�J���=�ۿ���bQ �]:%%�z�~$��np�L�%��]�s�=vOĚ�}�A�#�����{uvv�WQ�plI�
+@�b���9�u�<\�
���UU|�b��=Y�vI>�g��H$W>���\E'(6���oĀw{=,�����QA�LP���������_IRoĒ7{=w�$�o�l�](+����;w���
��H��R(&��=.��O��v�	�����~���m@��j��Y�ȷ����A�q'�����)����~� �_��3v��J>�4_|q)��W�(,��U���=3��1�$ ?o������統To�l�3�Qr_&MR!�>3'z��ִ︡}�y,I"��I��%
����U���:����c��*e�gqu�� ��m�f���1�o�A�3_7}{v?��B��M������.#����}~Ye7n�z�σ���{�/�x7�˝js�۬8��tV���ߏeI���Wu���E��ϐ?���\'��e_�e�$�o{j|O�\�T��lۻ  f�Oչ�����g�$�}�#�o��M<T.�ڐ�JO
9gC$�TPt�;�^��	���;��'�Խ�j�tM�ۜ ����T �H�뿉T3�-"�d�Y��l��f{j9Y&W��m��K�z� ��;Sz�F��vL��Yt���ni�{`ܖ���ZL��	��GYQK���u{�==�^��.`~;uxX��\o��+�%����3|�Ƈ������9�g>!$&�s����_�R�j��O;���wz�K>�&��gw>]���H'Ăn���'}��`���/���~ǎ�	�)?�U�Q@�(v%*�7`�[�����t/�\j�^u�p�u�?ߝ�w�����4�T7��ۨ	 �z�m�g�@'}��}9f��o���nWT �O�o�_�s�Ly0�n���>�]�I�Q���n]6���O��/������Ǟ��ke�>9{���b5����1�`��ޖ	$��{v��k:볷ܴ�~����$ﯽ,���S��t�!�+���jWҸp!of�I=�ޖI ޮ�oU���WC���I�vJ~$q-%h�$�����]���A�]������������y�zY ��w�_��vG\G�{F���9��ۢaTr.-N+�N�u��;Z=�N��&G\�.�5��^�#݂����s�#�O
�HJ��������1��`\c��0�S7rs��������v�u�c*荒�^�a�ns�`n؇��n�n��ʎ���X��{��孶x�����{n�iu>9��cpn�� �C���v����<���[| ����.Gtpq�s���f�m��Y�y�ۣv�qs���d�}�H��ʌAծ�L<[�n]���+�e��u��)y����aDX�+�����Ԝ�x�s��n���7Q�1��;ZS.xN�����m����8Ѫ����WwK�w��,�H&���+�!'���z�����!P:w*��i��7��f�z�V��J�7%��� ��������n��e�����Z����;>4Ǔ7T薔�wO]�O���c$�u{}P�rd�� �{�޻��z�T���������۷}�=�P��{�z�|	3k�,H7�ڡ$�u�ϭ����/l�O�d���b�̖�Y�����̂2��מ�έo|1ge�%Oo�� ����GW_���F�ʋ;{7Z^v)�
	WԊn�f��2[���glN8ݸȳYqic���\�`~�����Ν�rc� �]���� �W_��㸢����7�;��餑5{`dI��*I:B�^�V�?�|�u^i�C�w��<y2���^ÝSz�P���j�Ċ�g��m����U�`��r�i��{����q�{ض򧘃O����Ŵ_m� ��1�s^F)����AOg��{����B^���9|
���j��4�T �]40~>���?A�ާ���5���_Ă'/j�����	p�/S-�UH��vO_no�"k��#_}��z���~ɽ��9X���7�d�2������v�ő�?��K�R?��1�����G[������U�1x)���6J� �-��D�m�i�=�&�{gVݺ<:��Ӂ5&�����x�f�t���3���9[}vA ����s޿����mu��H���^�]�S�O�V�R,�]�4�V�_�ʺ��H&�߮�$���]�g��.P��Uu��^8.LP%"1o�_h�A����Iz����u��^���ټ����:^���\�E�����;�P��:d��@��P\�s��Lj��xx�ʱ��� >=������A5������u�,��_]g;̒8O��� �k:�~5�ޖHWs���^�H�~��w`�cH0��	���Jo�ző[�"�!OǨ����'����$3}�O�Ws���l�\X����[0����X��h�ɋ;����ͫ<x=�js��;r�`m�4�pv��OIDU
�9���,�H3;ޖ?�xg���nꚦ֖��ys.�?O{�w�/җ�D�M�T�'Ƨ��;s<|.]u��A���]�O�Ws�;����r���'�^x��4uE"͙�I��MweBA$�<��R�A�W�n�$��������ꄘI�**���=y~���OR{'��/o�B��~�Ʀ�Nd��(����P;�c�쿠i��)rT8�GP�yY�&��Ε^ÐB���Zdk��t�ʪ=��2�ɫ��G��^O�Z_��!!㓾����w�����棒�ɶ"��� ��][�=�Ik�+P���,�O���_@	�T��ŕ^P�{����1�xy�ӱsg����6��w`���<�>؎�y�Щ	]w��OT���[ ��0�O��=vtwy]���W�H�}?PbƲx**�B�U�7�,���k���3�_Ē�H�z���AUS��Ke���5�׾@�TѣA�Yo�/��zŒJ��K�_z�y�va$�5��	�=b�`�8��T�B��w�]�#��yD/�X��`�O�O]�D�w���럭Q�� �[�2$�$�T�*�3�:��~ww�����^�;�b�(A=']�O�7�v�и��3����e�P)Urd헗v�d~U2��Lo�u���a�������T�6v.q��F*��ƙMl�[�Y�ok�y�F,�ت����;��6���'�����(�-Nd�@�l�;�t^��g���-��^LU��5�W782�6�M���\+�;)JK��>#x��ǂ��f����<�P�p�=��Ǚ��"yKю�G��(���Ӿ�2e������M0 ��5ã7�Ǳ����d�/Nbt^�;r��w��u`�U�5��x��W ��kW�T�~�v�.tk#H�J4۬��n�n]�{�|�J����(=�����Df�<��c��DM=���ϼO��z+�'��N�`��YwZ�����_{�Y�d��g��iM��՘2�'���֞J�T�z#������!�(Ĉ���`��^X4录̷�Ч�� �/KO.[��gW8��g��{�U�u�/}��@���LЫ���6z1{=���X��1<Yd=;�B�n�e��}���{<º:M�v��0��9�fu�vŏ�v���m�>�U�^���A�p�m�tg�38$<�~��n��ೱ����,��ڤ�nQ,�a�.�	�.wt;�S]H������X����
��i�ڡ��������v>nn6��a����x��	x�'y����}��Q�l�7�x�)LZ�|��E�m����f�������r���^��g��܃6�rʍW��!7d���������[i�Ep%�)R-�qE���X�j����UYl�(�*%K�pX%��*�DbUJ�mX�U����Kca��"��ZYF�eJ �X�-UP���"���jQ��-*Ĭ�R�V[�0ի�-V���ձEZ�F�5YD[m`����ʉkF�T���`����EU�T`��TG	��Qc�*V�1q�+QA�Kh���)p�jU-P-����(��*T[j�mm����Vʴ��[ZS�U�(� �Uc1U���`�ѭDX�J��R���b��`ť���*����A�Z��������RږʍJ�c�*�ڔ��l�`ŅJ�F8�$���hD��1��-m[V+J�A�5"�b�
�DQ���5��a�	R�b1����-��Glm���}�����F�db{c�2�f���/n�l�Ǟ7<�9�����o1��n+��q�����PEٳōs���n�nA��sx��9�ƻV��u:��Γ�c���������h[��s��k� �xݜ�{
�kz�&�S۲��7h�9u��&ݠy�Pn^�Q�v��,�7.���n�ڢ��(�g��L����b+� ���r��"���m˭e��f����u����ײqg=7�ö��W����?>O�t��8XIӋ�<�����|t����gm���nC\>z��.�x6����W��.�7]-��y�f�[΄&�E�1�lj+���6לm8�zJ�q�[X�3����<�9ss۶�q6�kpq��a.m9� �g���K��6uV�1�=v���룱؎S]��Wc��1qd�籎=t\
n��K\q���n=�����X�̘�h,/M<9�Wo<�B��ێd���������N�nL=���<�b63�9�ى�x�݃�vu�]�ݗ�[յu��{>��.���(�X9s݂۫��H�=��=��n��v]�N��-ݚ{|;�g�D�u��vvr+����\E�NJʜ<P�ǘ�����:Q�c�X�n�:Ghu����7b��z+b��B�c��Zg���)���]pO?!.<9;ls�2ey�ۀn�=��mCv�p�˼�N�:϶^��^�a��K��lv�/-��{�uٌ!�m@Α�;I݊�yɺwtO=#u����*���;F=k-������hwlW1rv��p�`�ʶ������t�hy�zZK��p�v���C�\��p�'��u۱$��6P�=i{^q�;W<��1ۉ�L�ۦ7;�N�����ʮ!�Ҷm���q�8�v�:��J��R�o����>,��s��{bۡ��=vGn7/m]��î���9	։�g<�������v��;��u$�l=��:;`���pݹ�UY!��ѱ������\�]q��I���]O!O%��=��w���?�Sͻ�Y��kOqUt�g[��⣱����wm]o��m��̭�v���{h䰢루�ݳ��V�7��N���k��g���3��tg�v0��*[��;���i�0��i7%�mhz8̃I����b�Ξ�m��S]cs*Ʒ=��l�z��L��v:"}�d�Gh��ϸ���3®��6��ln�}�k
幮�qݶ����k�y!�J��U��p5���V����7����o~������QH�J��6���	������j%=��
��A���m���D�堁�O}};�`����Z�s ��ޝw`	f����9N��EM�Iz`t���)Qh:5,�V�� ��zX$d$qf�Yp�ܷ�I��݂A"f��d�C]�:�DҠ�CYo�2�wjq�^��D6�]��$N�z�H5���ӫ�s�%���L�̻��YG%H�*[����u�����̺b���� {�]�'�@����f��Fb��+Ik�%������d�L�m[�a[+�q�\yΎ:HK\�n$NZ�͹V�7��
��I�g�.���g��>�S6�"���'�T�7ʍI�v	$N�z쐯91��4�4.��m@ET�Ԯ������:�͂��3�k���T����6h~�z���P��d�̱Ny�!���䷭"���t�����h���ʜ��"?� ��5�{Y$�����$���&q��p?r����.�s�&�QL���%�&ZS��O]�H��ꄂA�g8:��*1��+�v�I��X�H���,1cY�UE �Գ~۲�q��q��d����$+/`���o��o�e`9�B�8k߫�v/!� ��:D�2�O�Lꀂk:zV����m�Qv�&\�ذ	�ʀ�{�������`�z�:�|E:��	��:�L0j���.j��.ӻtl�=�r������w����7��B�M��5��'���뿈s��.��ļm�%a��f]�H5�ʄ�a8YQ���u��h�ΪV=����N���O�$>����v�.�{����m^�~�����0�4.�;���C�u����ip~m�����zWߎq�s���n��vm��`��{���k¼E7F�g���ֽ�b;��}�Z�37UH����.�R�������.�^p'�+߲�����`����/��%�L�����ӻ�Jo�����z�$�Z�  >���0���5_ə?k?`�V����n�An��o�m���g{�bV���� �(�z\�m�	��z��y<����=@�)�AB���/��s�2�=��Bώvu��"�]�a����}��f��E��T$^u�Ő	��ozY��v쵞����z�.m�З��]��x"`MU"�7/y��#޳��b�{C�$��L��f����p�Gvi!����P�0��,�LUPD���BI{��d�|h��mc9��$��ނ��v?[�65��$���M����6���d�BOĀ�w�,�e`�s��]'S�V<�Ah0K���]�ѫ�3٬pGw�f��x'ҷ�T{���"|r�ڳ[jCeC�wwh��3{��J �"�}��������	�MT�o�Kt�Ig;�4O����]��^X���7y!$����$���S���}�[�O�nD�4���*���%sڶ�/lt�lLW��nw����g	qc�u[���m�I�F���@$���,�� ���>F?{7���/��]�H���S��&�BS�_,�4-"���tx�{������`�O���T���~���˫:��|�!H��"�^r��D(����BA$��q)��� ���H/�����	�E�d���>�g,~F��[^�n�zY �C�0�^�@bB�OXy���.�&�y���i"�D��s��ω��#x�U�ϓ\n��=�����/|�	?
�z@}����5�M��FDw�����N��m8�H�T�x�!�l����A��)�7��ܩ�;H�o��ҕ���e1+ʲ������/�w��wϸ߇+�kH;d�D`J���;kM7��]P���)�e�^���+�7]�h؄��(�t�Av^�� [�n�7n��Gl.'�F%�d$�jӹ��Nn�������9s�gs���Jzk(Û�;q=��i�ط;=�ge{s��uu=�h����6/\wd˹-5���mju�0vD���\�Gml8�Xϰ�gfv�)=���&��c��>�s��\���D�F��3e�޵�g]\�ێS����_���K���K�;0�~��Am��{�,v���˻ �����6�s-��&�=�By�{�p�t��1�l預A���I?W�� I7)b:E�=u=��=����:F�_:�����v����e�X$��	5�� +0��QR&��}"�>���&u="��	��w��/�ҡ��#%�>3�=�X��4J���$�Y��ӕ٨�m�X_ߗ�ـ�������><�6�y玾	�A�)�e� �8/��n�t���;��|�v|�s�(�v������� XJ�t�3\����>?W��v�x�ګ�p~�Xݑ�@{���pAK�~	���\��DD�hut�H�:�\�p�+�=XdUw9���.��|.{s��yl�4��uw@	���*�zw���QP���|�|�z���!Ewmyp$ǿgSa 3ܟh�p�?(�Po�N�"�PM3/����ޯ0�>��\�W[;��{"!���m� �gShU�#�5�H�L ��A^�; �����I�~i� ��8�a����.�f�o��d��J���Be`�_����z�@ ����o�p�����P	uf6� ;��@�'}����b���Ͻ���>}/��V�$74Ӻ۱Ų������	��cs��X��v�7���ݿ�;����pR���� ��y��@N��ᇺ��k0c��"���9��.f�%@���Y�b�7a[�u�����z1 y��;�4� �ӯw"�^ɭ�����$�Q<����%:,��enS�h��l�>V�s'������o=�̟�+f�2��A�~���!���'�1���@(�~���z ;����7�İ�{d�T�������,�y-��far�EUL����齗߾I��g�~�{ �j"2����5���+}u�X����� &���CH�o�Z������]Z������L8 5aD%�S	O�O/��7�|�dݣS˸�}�l��d�:l" ;m����(�//R�0�o�P{`�EZ����{r�nn����N&�b��0��'E<�$ϨѠMC<����""{?�  ;m�k��[�W�c��nH H��M���E�X���(�)6�����f���m��e 9��"��z!�!p�3�TToM�h%*(�m�:�4��6 |���'�0�q  D�:q�Y�ʹUJ�K�QMD�9fQ����+Κ�^b;:7B#��4Ȁ��������$�Ύ�m��N��c�=�l;2i����yv�ΟQ���ցgh\xTV�"��#��{t��޻�(N����-3�r�=�~ �\$���U�N�?��D�T�
R�y�o��gy���Qsz&�����p�H}��DD{��j��]�6yEo�����V眽a���g��ݹ�iOz�ۣřx�r.�r�|������J_��)��ND��6  Ns��{e���{�St�+�w�F�y��@{1z!A1�
��Rm��j�+�[������K���������o� %.���Ԓk,��Џ0~�eA$&!J������ e��iP�MEW���w@��y���9�P��[�l�~�+�/��M7:�D&$>�4� ��9h�H�����:^�Z�a_%��%��<�-�!A5 �:��D|�-��.���NtԻ�F�@|���gkR$��w-��?r���V���,�y��'�.�xK�͉F��[��ק����ܛNV%ѵ�o�M�RU���Նf˾�s��|e���̭ͮJoڮ��f�q�V����Vܞ�u����Ԝ�DlQ�)�;i�qsv�X��f���y���(�]�!�[��z�n3�]����o�n���2�3�z�wGo=�Fu�g`nSnZ��^�W�k�L���v{r�.���A[�����lgvƻj�vfѤ8�]v0v�m��gmi���G�3DgU;�{�����)=�+S����N^�ѓ��W�ŝɪC��n�\�i9܄v���-T���ğ߿$�B��*��n�1�����A;��Dj�NOk�p������@$vv��dF�DE%'T��6����V+g�f@I�z9����� m���-�$DV��
4��Ezu�>����ڥ�}AP��{�@|�-���
����)Zz������@|�f�j��'z[r	��**�J���m���;��K^{rg�n<� D�M���n�]������Kn��HF���Qm*R�ܖӐ"=����b��[���w��0'2[jH ��6�{��eL�/��믞pK���&��׵j���Q���qa7 v6�l�ә�q�ǌk���}���d���2��D9�ۓ�׽�0����og������9�Do%����Q|�|V�Җ��2~o�����~�O��:���f)j�3~���5�C�#\Ϝ6�+j��=<������V*�4)�bO�ۛ����/� ��~�t�������g�g�a~��D���!��������Dy�s����Y���W���P.paб,Z)�熂#۝�C@��^��*):��q�H��]���Bg�vM��a&�W�kԽ�0_�gz����/;��A��m� 9����L��%m��h"G8�?�?c��N�D s@Xٮ�m�� �f��G�y���T��wv�>�o� >^����㵺���{��W�*� ��4Y@�H�p�4�K�Wa�s��QgtL�\s��ݾ���qe&)|�sz����� ��v�XO����f��������l @/gsq�
uI�@�f��r�2�������$�mz,���� "��m
E%��-�{��	 蓺�S
��NZ/���q����4�[������	��{o3�:x�%���v�PgUg!w ��	K�h1}>5�4(VH�+1���I{�@��P��]K�˙J�O�	� ��:)[΢�ե糘=�2������rT���Ѽ���=�Oґ�p��+}�a�����?Q�ѝ����\=,��Hd8�Z��M���{|7֑[[�Ű���Y}�'� �	�yxߺ��4+�K;5xt����u�yH��&�x����8����x�^�P��d�"}M�M(���s�32^Wj���{N�� �>�H:N�>!,��{�� O���G�s��81G������y`�?sh�ͧt�O6]9GX�:w_o�YyJod��f��gw�`�;�bX;�ɯa���C����O_������3G��M�%���KHv��@�s��{p���/v3�ϧzP�x�V֜�ܛ!g���\��6B���#��8�[�b\���:�/kҙѱ������O/��n�KV�{l���#���fr-�����}&�|�a�22��N!�uq���4�{zrG�a7�R��c�x�q\�w&��/L9��v��%vTgn�X�g���Œk�vW��?sF{r�����xzg���.us��Xra=�W�V)��ݙ��蝶�]���6�i,=��}�c�M�����]�ﳸ읲��˶u⟦߭��Gu��5Y���`�t������Y�U�Pqԫ��������452:2�Z�1J���B�_v3{zu�Y��z�0�e�I���咞j�<���U�h��Z�`�E��(TQE�FQŖH��DŢ%��F����m%B�IQpˆ�kKD��,+l�,QA������Z5X�EV�Ֆ�cK
��QE�QJ[*%��0�W����+Z�*4�"���a*#UeJ(�cj�F*��b�µ"�*1A�1�
������a�
�Q���,D�m!b�*ł+mQ`�����)Um�R)EAb��TE[eX"
+h,hZ��E�\b�,�XQ�֬�EX,P��[T��E�1eQ\-���-��ְD���(�H�"��Fز��U�1Qp�`�T0�eaX*#RȉiUiF�TT��D6�b�E"0Q�i��l�Q@J�6��b ��
��QUUaX�+?/�J�߲"? �߹���~;[�^�Fh:�J�#VIs�Q]��i�f���5�~i���s\��|V��i���n�$�=�d���&�W�)M�x�s ��z �;]�*�=A7��4�H��n�g:o�諮����������Mr���Ƚ2�#�l'\=�Z��mV��Nvc��7��ߞ�T����E+���z8�V�j��Vs��N˽���k���@|L�mP9Q�Q2T�"b[�/q�`��t�~�N:�u�ݽ�ȁ37����i�?���y_���/;_��?h�&�L�I�iF�j�D�:�?�"oz��:�XD���� ��o7Ds�6�R�Fj�|T���N_�v��6V_��v�]�F����@7��I��{���rl�"x�au��#8\��4��/��2�x�=�W�v�����pף	�rg.'���뫑5��y��ν�=�����+�Fa���=_��x��%�V" o~��I$�=��5�s�簾��k���Nc�� ���a7�#��u{���/�4i}A�KG�����9�U��v����qې�tv-8�A�q�saB&v*���D��r�[�H����8O�=����^����m;�d��4��]K	$,��m���!�B�)w��$�C�kU����/ڤ 	�~q�]��wh�E��ZΨ��s>z����.J�*h�b[A{��`�A�}͒I�$dQ�z��n/$�A?u��H��]���'�G����L�h�l��˳{T���AۗM0�e�]�	%W��~!�Ē�]]���3�F~��������Ղ +���S�6N"����7�~p� K�w]����O�=u�T�d��9]W<�/��7q���`w{6gr�#�3�]��N�R�R!uI�c76/)�X3�\dͱ^V�6t?�������yAPm+�=*n8c��=p�;�]�_#:W�\���]��a:e��v���8�݌���صɚA��p2�#��G�]rf�����ڹ�0�slv���u��s�˝���&ˎ��Uϧ�.��u�V֠g�N�瞓En�\+�;d��:��v�Mh��x�`C�a� �c��Է9�[`�8+S��z��8;d�,����N�R��i�y�^�7�*8��0]�f��Ҥ����p�J�=V,-��`��
�w�02\=��S�����@)�� S.$U��M�M�Sh�c����{�{��Iݔ� �wuݠG��^����d�ӯzp���W�$�w�l��!�F�.��$$�;���2I=��� ?��Զ�� ����� ����4�#�0��Y�H�]���Y�}����/�@�s�`� ^�w�4 D�:�-zyp�^Q�{2�_^}M,D�e�H����l s�4ˉ�v�R���Ahswwh �{���'9�hMS�����	��&��a�٢��=`�3��f�qh��&���
4]	5D�HT��}�|
	���
��n�]�����{�H s��0���T��y�]� {\�!�lj=Q?T�3!.S���j����2x���N��{tYoVW7n�/@������uǾؠ��#g��1yNף�m߸dc˺�q�4Ȗ�O#v�e�y�La�/������Ȁ���1� D���@�����;���k٤A����S��@�n$U��M��y� �A;�^��AO�j��._έ� {�jH�]7�q�d�eJ	>�Uk��!R�^�*/� {�{��" �ߜ?� .{�w� RoF�� ��ͩ�L����`��/�ס�s��Y셦��J���/�ڹ~M��h A�{���z��\�oXv�犖6h��!T|�,�A��ޭ��x�m�C׭c��݇	v����}�!�vӒ ���N6�� ':��7oz��Gf�w:TSۄ�c��H'�l1@������-y�n- �u���O0��� ���"�{�v�.w%}Ә�Į��XJ��U5H:4)����>�l{{�� 	*_Q��RZ�.���W}�3K����E}�AF��A�c\�#2�!�P���ͮ���W�O_yM����*w[���U}�f���=8�|�ݛ�? ���M����������)��"��I�M���O�&:�s��+t��z��޻����L�\��IԮ<.�)����Q+]�����y����nwT��������6=�����>�����n� }.xI�y���c��ݫ�wZp���6L\���o�\����ϙHC���L��Îu�{��R�$TR	�?|��� ݾ�N����l��g�w��A�L.��v�_$�{�ل�$���i���c3�.�ğ�����ν�V���E�ل�����!��z"AFu(���S�uO�F�!T�*%1��n�X|$�nz�$��w����礝d���o�� ^_Sh��5����D��>ʘ����>�S9���}nۋ K;=,�H���Q��P��k4��'Bg�G��TK��nm�u1��߇���w��d��l�T���c����vF��N�FL��.�{/�U�4;z�'���#P����2o���M�K��� �˯F�^-λ�t��� �{:���{{N"��u惖E��翼�����Xጻ�K6��@㵺��v����l�<l�k�du�{o��ߞ��&��n�>ཽ�0 S�~p��.c�'9��q��O��݄A�/oi��2���-XN��0���L���ߓ�������������	 �κl
I���{����ܛ�Ud����E2���[X��$%�8"I$�_���D#z�%#a"~��<$ N��0,1@�
�
Uh�{��/g��b�{ѭ >
{������� v�]�]����� ����U�#�5"�R���>�i��Dnns�g���6�Ouv�\��� ��m� 
�s��3�t�|�g~ͨ���|h���87l�E�V�2�:m3٣d�J��egG�Q��k��W���.�9w{�'��&�o[d�����fj��^��hqy� �x};��ι�����\1��-�xMs����ɱ2{<��g�m�X�l��9��dm���F�yyA7�u�N}���m�.��M�\h���=0Ǔr(F����9B��ix�G �ku���ф���������Lg��&���=��^6z�a�)��I;�ֻt4��}���v2�=�mӌ����.�M�s��.��.5g����Yv8��jx�ol[Շ�0���'l�r���u+EВdp��K���ǛLb�\��\���W�� '�_� ۝wi����L�g[U[��:m |Nl���BzF�3T"���]�]�����k�}C��:�]	?͕6@~�����PHᮑ�����Wo�%;�<b�
��3a{�ۑ �;���"TNnx��+.�}��D��m�$D^�sw�	SP���H*S1Qr���wm_\�y��}<܈���� #ם^�r���^1$����i ;�!S@Ԩ)�{�wX z���V�?J����2������ =y��
�>>ޒ����IP��a���Be�F(�jϫ\v����g{kt������;���~q�6s��HN�mη ���ŀ�^��8ho�+��\�ec'.y� �n�N���3�*��Rm#*��C@�s�}����,lܱ�n��oJ���Z��~�x���A����G��WA��yd*�xoqp7Ì��B��N��]wz�8xoOx�����A��L�iV�o�h�O9<�
��6q2L��G�|�b ݯ4�@|ߢ�}�n1A���q�y���}鈾Dܪ����t����x�^���v��"�W1�>�{]81b���]7�I{=���<y�0�4���ٿd�'��Lܹ���[���z�E���{��" ��鰇�\�L���l�4SI�dH�P\c����n9���c)�;A������?]����q����^{:�� ��g�Ґ ���������K��7��sz��:܂u���U"%T�$%�A޼���vG2�D� y�x� H���"�6� j�Ƭ��=���E}2_�%J�R�2���� |Z����ƿ�b���Ư/yw���wC���,ByY�4�����%��m��V�ս�@�s��ۿJWT�)--�Kt�}�a��� ��Վ��\Pc(�b�Vjz�w��V���n;�D0�}կ������|�R�����<yhw6��^6(�"�����\.I�����
^����8h�GW]6���w�����[����M�R5�+�*��5��N�q�=s��ۓ�뷧ڽ��=F�5��ۿg�\:�����w� >���0�}wa٧f���f�3��M� u�M�����AR�����;��n,6��e�GF�z;=gmz!��+�� ޾���Isߢ�x��'׵;䐕��9T�R���7״�" �����A[y���t��`|�Ve7��������|I�4�2�0B�v���f��VJ�~�n�^���븋�e_S�w���P!I!�ϲ��bcxH&z��-x���N�-�Z]���Go�@?n�"姩���k����!����%%�ތ��?n]aQ�wwM����D�TH⽯�+[��b���&���F��پp�@-;����FW��ґ�:[�"7:T�e|)(3��޶�B`m�q7ase�W�L�ꍮ�w:�������Q��/�m㦘 ��;� H���g��q$�������� ]��N�+�Q��H���9f�:l ɜ��똺�m�L [�@|e{���Ӵ�l5��N���#'�g�@TʢH)���m��D6��� =5�9t��Dt��h~���"Rڞ��U\x6�*��Nͥ]{V�}���u ��7�m{���$�Oݵg��J*��q�%Y;٘�Ě��a��fW�h	�y�W�g�+s]�7�ח������D0=�M�%[y۞�E42���rq���S�����.��2�����:�in���5n�������m˵]S�����Gڻ���&w���b��A"cݿ{|�x��N#ϲǻ(y4��ٻI�(�跟�M�3TQ�PwS\z��i�#yZ4PjW>v#�a�K����˓��H����~�gY󊼮go���z��!9��xO`k=���G�*�=}�p@O1}��4Y�绱״{U@O{�PP���n{������u�Ҫ��zmD]�E�=+�zKk�ҩG��d��n���{�]�鐡S�qӞ캽�#�+u���\����ӽ&�;��c���5E����r�<棊�;�ΘP�E�����t.�V}�������	:.g����8�qt����83��$��}��rFT8'-Pr��c�z>n��0�Ʊ9��!6݃ʚ���U}��.�cקL�P�]�u�BQq'4K�����B
X��׹�ע�w��XO��a��#�\��p5�|��������Y���u�p�#U���d�"]�xC˼�q�hL,������8��ǔs
���[帧v֎3�rk��s�b�^'Fj�4�d�9`�f���T��]�@;��gZ5��֨ϖM��~�y���Ν�[�`�e!'�z��،{�Ĺ{WO`�N�t51���ۋ^�i��q�������F�C<:�9����N�lM_wbU_}�y��nǽ�X�yk�9y^���>�l���݄��{2�c#�U]y�����l�i%U}Ww͵��h��iAb�JR��0���� �8j��Y1h�R�",X����mDL2��ŀ�R�Im�+b�(!�Q�UHa*(�Lb���b �)iq�W
��+qV�f1Q�qJ��#-�6چ0����`Ab�%A\Qf\
-�b0�-�0�q�6�[p�)���X��*a�#ZV�8�H,1f0(U+X+�7
�0QJ�J%�+����"!X�F�X�H�U�
,TUAE��	F�*�-m��+B�J�VT�0J�0X(,b"���ckl��Z��Q���-�6ʪ��X�J�eQPTE�DTiQ@b,���5�l+-��mTE"
�تDdQED*T��ږ�ڪ%�d"�UH,F*���UEU��)R�UDTH��UEU���Z���*ѱ*PR�AAJ�bR�� �,Т��V[
��آ�}�?�F�ஂ쫸�@)d�fʞ6���6��'7;Wp��qk̥�Ϙz��{��=�<bL��]ۇ�X����m���V���mp]sV2����cZ�S�Vٻe�j40u�Q��nػ��-x]�x��a�۞ͽ�C�x�vv{]�;�77����K�NNq����Nݱ�bw<�#t.�ɫ��v�9��������|:5+�ț1��n��K���cn��;���fxI����VhkA��kr�m��5��u�um&���7/\#�b�
y=͟:w;��Vׇ���nޱ�n�]m�7cˌ�${���w�m�s�>�����m����;`��Y�ۣpd-�Ny��n��;�Dr���-�5�ە�72tM��;]k�k�8��%��!x;kr�	�lN68m:�zO,C֮{����{v�f���¾�嶇�Uc�'˫c�o��B�C9q�h��nS��;#����Kȹ��RS��v��A�<:^�p[�:-��3�uю��vMv��u�T�8m[��v#�Ǿ.��\U[�����j�d0���h���[[q����wL��Y7;�mO>n��$;M�H�D&1q]��xU��q�95�mg�]&�P!^�eD� &����D jV�\v���m��)�l/%�]:�7�DG<q�'�����43�ɛb�rV�r��ؼ�vu�n�c��=��.=�f.���[�%S���P钼<I����7�v��0u��8�ˢܼF�N����{c���;#t��S��lm6u���2��2�<x��ݵ����U�nI<�n��퍪޺�e�f�ɶ7	r=��u����[�8�ۊ�m�Z۳Z��d���+�)�c�:ZWz�Gon�q�����s�Y˪�n���u\wmڸ�g�qwn���9�a���s�a^���l���ד����J���=���x�V����sr��U��l1��D�=�ƋZ+#\���7
OX��� �֭^D�N[�粉��[X��%ۘ�gnS��s-�ܜ�;0<��V���X�������uۉ�z��ݠnYN����,�I1�q����K���yxC�ٓ�-�$�ϔ7.n��ƥJ��yaݹ�w]�#�ۃ�;��nb�U9�dZJ�鵉�\��u��u��l֤<��m��m���<6dǙ��N6";`�R���.���b㎎���9.�rq�[%�M}����рy�Q���۵` w��� ��<�Yҽ^�ޕ
s�7�.� ����
�8|�EJ�L;'/�m�#�n�y���� 
y�0	�t���̩�{=��o'��%x͔�e҉���,��Sh�"{n� ���h񘊗=<�3$���I��/}�/�t���6)�
�Z���<㵅���3���ә~p�H5�sr/oX���$��ꘕW����1M��?�S����o;���W�����Τ�_�0��Λ�<4�޽���h��/�B��XD���th�Gt�@�7��-�D�'Y���i�c.�|���s��;��
ig�i�;�m9��>��w�gе�e\^�}��ޯj D�M� ���9H �*���y�[�A����������gk�ē���y����wf�L����_�t�7H�M<�2����<�����y��� �@Oe[ .y�wa�z׵��Y��U�	�B��ȈR��T���%��� ��w7��k&���یH ��y/�+��fbH^�Ґ��$�����SȔ�T�sv�#�o�r|��ل�IVߪܡ�u�,�gBH��
Qq�"
&j$�W�Ggmݥ` V��0읧����Q�����l��f�H��*X	�qٜA�k0�n˝�t�7n3��jnyu�l읇�����+�	�4�l��v��@�M6���Vc�� /ټ�X g_�4���y_��"_�������'6"<��?IQ
i6K�����u�Eo{1��~4"~��� Y�M�� ��㧓���3;=7��@��"&�"�R��C���� �u��R��w����<�v\R��wI:����A]��{��i�������H��{pl��	� s�S.�����=����3�yn��G{{�� 	�t��/��3=G�XUM$û	ns��'�\�� fw;�H fߜ4]�~��Q7n5�dPovkw�]�z�P��)T@�76� 
�no�UU�-�� =]{w`�+�)� 
�h�6]c�~�=җ{gKI�Z4#O{.���ez��ɮحu�݉������l'��n��RP��Q:E��n";��4AWu[r�7��Z��������*�m]���<��%2i���	W��MA����͙3^cw�� 
�k�J
�疉�����<]/�f$��4�[��$:�	ߟ]��I|��������=�T��^��;"7�Y�m� ⻦��A;���B�5
�S�r��.=����$��c荤J�ڶ0ٽw�WO��qV���މ[�1>�T����#�o��l��X9K��/�[w�L�XK���m��x;쪕���"��մ��@,�O2�\�1�D��%���/]6  ���via�ή�MR�w`*��c��}t���]���w7�$/������%���r��<��/[��Zr٣e�1&�n��v�*a�)���{Ծ���"��wkm��A]�M& �7������g K{vE|��*����p=F�P�iR�Ggc{���B����v�1�{ܤ>�ۯDC��7��-m�������ze��4��>�M"�I'f�S����o;V�Dw����_k��bj}ݼDr�.�D4�y�I ��0<l7�t�t.�N������WE�٦.ٛ� n��a�Dk����F>���w����Do�V�6��,TMDTD�*G��]����^`�ӧ�r*d;ʖ����o�0��޻��粮�'5<��W�ľ��rX�����`�%��"-aʇ3�͛P�\;|�p���y�Uj��^Y��<3��ld����(����M���4�
R�,�<-G$�sg����'�v��O�y��
8�ۮ9+�{m����:m�O��y��\x���tb�����q�.3��kpik�{V�n�;��T�crU=�[]��Km���.��9-Ɲ��@��}�M秩gnx����$[69���\e:�۵��պVv�);�m�Y2�Ϊ<�OF�`��'>��T.ݔ�u��f@W���h���{��Bq�jx��(uV�?����{ແ7%܎3���}�!w�~�ª,6^�w��h�{o޼���_]z+��>�olS��s)�C��w]��;P�G�%!J�1�~� E�����o�q����M���� A�W�!�U�wTN��v�Ȯ�uv��B��
&��f�)dv_7�X �W��<�&�r��V��fF�g{ٙ�H$v��	o��h��4�p�����;�yD���ω���	$����@"{r���GM�� �wل�x�B鰘%��М��]��A{t�)�^���S����|��� k�l @"{n�Qt�:<�g�Lo���2a����)�pq��n^ N�N�	�G�ڽq��Ro�\���@�Df�8��ޞ� D{\ Ou��
�H��_E�ͧ��^]�� �k�o����>��UD���?��6 ���t�ȧ�-Տ��,�t!���R�/��y�i$R͎�I�>��kȎ���O_{�.�����` ����g��G�5�"������9�r��y��Y���`|=�N"H��L�}���^U�$�`"�)|ڠ�T@�3�o�`DOm�`���]�>�x ������q(Y:AI��[��m�<�w�n4�H�����I�Y&�U�{ٞ�*�9ƎRʉ S-���s�Tz��T�`�
p�
��0@ ���X��{Խ/:=�{3�Y�� +6鿂"
�޻����v�/���A����Ǵ80-��U���\�e�q�S� �u%�`����-�/������Hg��J�♜�T |}u�` woI0�6ts}��wh0�T�Lr�{)
i�!�!N��S��I!c��yl"nl�zb"!���8`vw7h V��/*��<�+��^����e��z�@ ����"��;�d�¯=���.�cc�ĵS{�z�����L����c#��.3)�<pjš���i���8���/5/����Gm��En]7�@�
�7����Gg�~�)
U9h��nn[�K9g� ��즘 ��ݤ gM��
c����]	�jX	 �'�B��m�aڵ��ff"I���`5�ѱt=�=���cg_y�CV���� ����خ�ՙ/��J�Sf�L���e�-�mգKv��M�R�{u�<�[]��[����w��uˊ ��
��l>^o;���Vu[q����4���D�m6����	͈�8��2T���ӌ��rM�Y�{�(g�j0 f�m ^Ͳ!��޿{�4'�9U�!8�W@T�ª�T�����Շ�|�7� �!� v�l{��,�y�w`����j�����E��6Zp��9���̸Ӛ���7� {��� ��{�L�z��/^�yM��7w���z8��\�EԠ���Lx�*'i��G�c�_���?P�o��
���9ϗd�Zh�X���Wp���~$�)T@噹-�!���nrf�k���j�g�>�y�v=�6ܐ|�+�m���̹5~�X��H�SD�"�@������ys���5����q��������������[r��O�;3n�XG���C� +���h�rfy�e�ꗻ�v �t�jI�q&��ҢUBK���R�>��;�׉���XG�f�4����ے{��f��~���]�����j�J�����Ԁ^ʹ� �]fop�2���{:鿂 >+�m�!?�L@�+F$�-�{�?O�=���U�Ay�^aU�[���63^��<��@n� �t���">��&��Im^�9#�����F���9��Y3�T�
�3�D�ٶ�{w�����~�.M��CbWqA.܏<��Ț���`����>�yR�-g�&�#�a���bˣ6pQ��K:}!~E`�.0~��Z��*��ۑ[��Z���횹�i�عJGtX*`��������km��ruۓ�ɷ��<���\�o�5Ɓ�>���sc1v�t�\���	���m�u��۷L�s����L�!�}$���6c�=��y�� ;T�vW��.A[������ε�<k�E����)���]s���i���t�ǚ�};V�즓�9,ɭ]�@�:n�N�.D�]���Qv����iu��n������/���QL;�W�? ��fۓ��޻�]9S4D�\eױP^�v$��f����+�&C�)J�3�:��F�V���3)׳� �v�� ۯ{3I.�A1�j�HU������ӈ��F��)�J����'	�~�؟�B�ȟ��+m�|�6ܐ =���ē�m�htR,��=�c�]>� q�?�� ��uݠ I|�}�bi��滧��&�4���9�D��Yz~;�hđŭ�{�~�D��ݺ������6�N׸�����x` ��Dκl�//O���{����@� ������	�+@���\�nz^�ۗp�m�]tnuMnu��������&c$�|y-�c�w`'�~qa#��<�����O=�M�_v�{3 I	�R��j�R*���SBH�J/�J�x��k�UYe���#=��[_Ab�z�L7,�m���׎7�U�Z������#�S�O��%*��S��F���_Ua\^l����@������|;���ʻԇ���-�l��14�h�λq`���� })L����9�]�Dκl	�{� 
Ѡ�
a��M��S��ߘȜ� ���� <���f��x��I	ӽ�N=�#o�A0�PG6S�S  6{]����l��ے��$�g]݀�Cκl" +�m�\l[�&z͏nw�$¦�*�(�d6[Of�!�Оԯ�b�­�=�v�:�S��~~?���n��n*��� mך��n�1ǥi�k")II�^�]��{ΜC��q}Q�$��RI-���M0A���W)ͳ��~�{����~q�Ev�x�a ���\����3JyUe�J���C�EDMD��f��@v�4ȀZ�����kK��=�;�hCY��`�NcЗ*%{~�hz��ܻ�+�6w{rv'/mw���.u�)�ؖ��=.�4iK���X�5���w�ٓΊ{aG�~{p{W���ltQwn��#��d�gj�ɰ�䓻��>���TC{b���!�76��ֱw�<�e����_!8K�q�9Xa�|79�0V����8���X�*��������t�u��g���f���X���sS!�����r�X(:4-��.-�9iZA^�u,��g���:���O���7��0�3����/zg����Z��5�Ǐ��0/L@zߥ�K��h����f��\9����2�ҙd���.Ջ�{� �0��k(�^��i��	�v��Q�D����,����v�Ύ򍘮�������7r��t�����P����&j���������;���Co1�#�v��ٽ�p��t�[���]B�Y����;�e�mm�o�Gw�٧@y�Qݯ�:˵l�O�,O�����]��!��Dy�)@e���[�;s؍���s�G�{��ʩ��l���ԈK;J��J7T�Tsu&{h���$�&ʫ�cu��xu�E�pg��1sL��134˩L޹(���� �M�����G�h�Ԁ�_^f��_��۽�L�U=��:J�ݷt��'�
3HD��_m�7��G�ķPD�;[����e�s��K[4y:F����n^�Q5uں��x�J�M��`����~���_L�p�h)����t�*�w�T�r#s����,�����>�Y|)z;^ȵ�zL0��Ee�(�����ʐ�*����JDE�%h��F"��+-+++T�Imb�TX�KiXV�%b�QU�԰QF�U�KaU��������*jJ�F(�m�ch%aF�-*���(�T���"�1-�E`ƲTQb*��`�Ym�
��T�%d+iR�""[)R����Z+��"��j�%k�"�E���iF����Tmb"#Ņ���eV*�H�RQR�UdUQH�Kk*VT���"��ёT���eA�R�R��++X��DeE��� ���X��b"
P���"0TjJ���F,��TX(1�QZ�Z�#�(��B�jB�(�eU�*�AkP�*,-��EX�*����[H��+��B���DBU��[�{Λ�+�鿂W�a:��b�%�_��+�]=���W� }�^�a}Y���v���>��x8zyE��5~���u�AS
EJi�D���� >޾w���W+k�k7OHz�������ۧ%��{3X��)J޸�{4��F������`��I�m���q�^ݲq�0�$kp��\B�DR%LU R��{���|{t�� �z���q;u����L +މ�Ng��v%��$1$qk��r�?_��20<Fo�T$���{%������v;��]Ln��&z=�y*��1<� ���f���g�x��ٷ�Հ��l����fn*��n�+�鰀޾�������D��MD����鞪Ptu�Wy� כM� ;����>s�]R�]����������\�W��Y�e�:f=�������n��淘���n^���{�>ap��$�t�6�s���Kѻ6|.9؈㯺�J����)��f߳�Շ���:��7;�t�Y�UU����Wϼ�ou�v !�:q���U�eoX��ab�-��	$K.�Ǝ���
�ٹv1�Ar�b:K�kY7WN]]������"%Q50�R��r
��i0 7;��$�/��<%��jcA�irT� ;�����%;�aMi��\�TԒA��UWEsg�^�%������f�*� ��[E�ꛚ�� �Y�T��U
j�S��u��`ݺ�@ �z�U�48~͆ 
�{.��>:�_[y��h�Y�Jn��;k�6ny�mm/MJ�u�x�� |OeӪk��Ma옋H*ﵸ�R�?0l��F�j݅��VM��/}�`Y����5��1�D��wv���"!�}t�Q�Ճ�|��y~����D�{l½��w�}�<nu��y�x]){{�kH��n7�tHT�������}_7'�9�i�4�<�>�������l7^:�M˛�<<m���c:�v�^��܈Y�JW(6�y��[��7&}n9��v�e���A��ѥw��	�s���ձg����[�u���M�]V�8[c�f{g��cs���زEnNɌ��\vաݠ�6{g���Z��lq�i���\S�مv��{�aF.���8��q��:.�����u��,\�1�+��]լ�쑸��s�����k�.6�^ۮ��w��1[< Iݰ�;�����\�@�8���`�=��� }~q��=�^���N�{�w` �s�o�O�l���Ha8�S��T������=�s}��� �^��q�&���"�	Q��.�]_����,�$l�`���
W��M� DN��`
�K���{�b/�s�l "o������
Ć$����Y��ӟ��?a�ע��_�0{�n�a�L�WEI��Bl[����Yh�L#�ez@ ���j̮ˊ靌�f����4@�t�@]��w>��q��G׀�j��0C���ɡK�A��ی�.�m��@��u� H&%
�kt�Q��!M*S%�#w�M� 	κl� ��ۻA3鸰��ٯ��'�鰁 �7�l�*��� �MTc:�6�Z]�^�wǩ!7��t���x��䲬2Ń��?����p�WF�>���E�� /Fk���.�$ec���#�e_L�֒�1S�s�x{�����ۻ�!~�^����+u%U�y"�*��L�Vl����� /��ݑ���g��(sY�ѿ 'rm��v���=؋��AQT�
Sy��:3������nu�1 n�kv��"���d�����~��k����Y{*�Ҫ�UT)�<����m�y��]3uj����R�c�n�]�� ������-��PC���60����URU_"�&�y�v�!�t�'�w˧�{�l���7��+v���~c��Ʋg�L�ws���nvs�`��8��gI���Dz�VI��ݾ�����y���F�����r�� y�3���5���U�� ��s�� y�M���8_��RJ�����A#��X�G��ޫ ��� �{�S�V�$w���
��n��Y��ӂ���]��~lP������Aya{��{�L ��Tr��n��E�fz+�aY��G|e�]�_�:鰜�J�UX��'pj���丄wX���0��]�n,Ϳ8h"����9#�oF�+($���y�O��I*�*�(J�W�s� ��+r��ﰃ��|�P�ۗq�t߈��g]6{��3�g������X�\)��qF::{k�6���&O`�xɺ��E�b�C$�������k��uQ�������Cݛ��u�h�K��c��qO{2��!�M������i"46M���p��g��5�z�';_Y }�~���?� ߋ��r����Q�ֻ�=�@�b#Bń�Z3r[r	 �t�`�7*�����9U����� Hzu��h�ΛmH}*��� J�T(ds�o���=���n{�Ǽ�A�>� ���� n�]��'yy�w*S b�;eEE)�lDt����b��d��4w����	pɯ۽wWw+n�x�^�zSΦL�8�N��5�}y�|,�"�ǂW
�UH��M8h<�q�'�$���>�~ֺ�^6�^�|� ��Ԑ�]ݾ����&u6Mn�z��d6�q@w+��pQ���rcg��i�m�Y�9�M��B���:�I*�&�l1��Ξ��U�nb n�]�@z6��x���/�LwF�d�=���O��E:�PĒ9���˻V�����y٘WC�����U�["��n�A��t�ƿ<����銉"`TDǟ�3rq� f�;V ^2��ٙ���� ��D?�����
E��:���H��B���g%f�~׮P{���@󳛿�@/���w�+츈�Y�m�*�(�LDҡG��Y�lD-��	�C-�9�gl��D�]N�m$����v�Y|�����q* �OeS���x��r��e^�8�:��ko1{�P�W�x��=��,��6OFo���w#9�ݧsY�=�Ӈ�N�Q!}X<�h���v�<\f�=&
v.�}�wW6Q�+D�vϛl7j�{��L,L�E\�mf�Cr�m����ۡ��N�������W=���|����k|@��&;pn��ԨPO��p��lr=�-��vg�D���)=hMv$�U	����K�٩�5�����F�ZM�Piz����3o"�y}V�[!tr�<��($v<�v��t]f�Wapz��y4�q=mo�������T�	D�� ���^�sqh���o���R$�G���Av�u�$�p;lU4�b��m�i��Ϻ7ٗ�y^�� ���H ����2 ~�[���8#"��4��'��J����{�.�X|@�r�� ���u�0�M�p���{���H/�9�iS���E2YB�f��̣�B_+��U������
3�ߘ z�)�N��\_����۰��\Π&*�&=,]z�a�=��裷���]ϽS���� !v�y�����_�WO��*H[A$J!B��ID��iknQv�3�Ӆ7T�+���pe��s�������IJ�G�n��� @��<�$v�Cisn���7���]�}�N|��l���v��T�U [-՛)��h����u�a���L'MS�T�������{�uE~��ާ��0��G�2�ϐ�oڀ.H"x�u�q��q��y�<�7ɲ�>���*Ob�mT���u�V  #5��DD{���|��ىns{*�����,�
U}D̡7��L> �S��/����,�:�S�}|�DB�y�}�^`.��m*ET��3���G��dć�n_֢"�ny��7u�mØp�:'2��כ'7pq�B�sA�F�~�� ���!������	?|� ?ޫ�v>�� �nVn)6���DUJ��ݚ�9训uƶ��<
&y㳎��t�Eu���k�5�<5%�QI�4�;DL����H����4�n>�@������(�)�Ř!7d"�Jf�]��O��a�b��o��153�
�'i�F�=��0 ��y�Av>븋@��y�՘�^ЁS��K����U2j�L�Vm)���4���� S��g���M�����Gr�ٛ�G>��wG���Q1#�����}A�hMݩ�]�G&w[�7���G�F�1�=�nZ=�u�r@>̯?��}�v�����E&[K{3n�cϩ��r+i"{����>g>��"��q��3��c;�5 e��a��N:�"�UIB�2�w��I���Ϟ3��M䁧�N��8 ���7@'�m���9	�k�����-q�\^���6{�E�!d�>�v�s���[9��	�M�w��o��ߺ�<�;��6�+��;sqa}�ߢ6�TNF�{)���l" ���]�!��'B�<���o�~��?	e^^�D v��� ��y�� k��[UW޾���QI� �N�
ѝ��တ �z�� >A+�.7�AO]dj �^�ݠ��~����&&��������=�U�_ƽ���D 6��l }�o��+���f��E�Y�D�l�m���<6�!����c�>ɫR�1'\��=8E�P�|6���̓9�8�����m��U�r�z�8�ۼb��~ү��x�5y��w�Or�l̨��T)�Bmϱ�� {t�dN�WCܽ�]������\g[|A$�_�d��z��RP��<r���^{{sx��܌���ۻNۥ��{b�o(�&���J���i��T� ��-�=�q�q�~~�@*�8h0#ٗ��efuݠ .3m��T3�Ȩ�*`TH,����-)�5�n;�}*ȷ����@8I�G��H_�2@y5֮���숿�+�������j� ��n�" 燦�v�ޮ���/�� Wmӈkʢ5Ej�ēJP�>�x���X,��+��:  U�~p���ݾ�s������1�/ǹ�5%vȪ�"���$�pµ�6 ���vS�{�9�}�~3=- �Ev�6�����,ҝTKz{�w�Z�ԛ}��N��V{��M�=�=�3.�Nf�����ws��kh�����J�N�|t�K��0����v\��Hq�e�m�F/)7��w�3�{I󮝙)!E�d[@����nM�)>��VM$ҭ����6i��K���|�v�z�M6�oڭz�V���,�	+El��G��3B��U��>�}�V�7�t4��J�]���"!���6Lv�&�K���05u�krv?�H����k��Z���w<�2 �5�s�:z�滹N��X������x���lgy����p��ıa�b�s�&�H�V���՛�X�zo�1���������p��絥/��DǸ�Z��6�V����.�ƚeR���Ѷ1��<���껞�;���{�ON�Ԇ��|<S��A鰏<}�ܽw|3�_Z�=3���@��$,R|t����4�-��Ns��=�5���Z7�NU7d{?i��!����s�|E��ל����RRg�x�V�r��G)3]��N�oey�ٲ��ޔ����_勫 �u���_��K0-�L��\��UeR���T�bN�N��Z�d���,~��OHwě�N�M��B^C@�]�b�l`����86�Z������Hoy�[��gY������A�6�'9_�Ղ=������"�z��x<�gv���s.Kbۡa�$��6���cu���P�ȤFERU�J�+X،��Ic-KIEb��*�-�E��j)m*�,X�X�b�,-�-�XVB�"�B��* �
�VT*��
(�*�J"��T�ȤPDU�"$PRV�"���"�[k�Q���b*��QR�D��H�A�X�����Q"��,+�#mQb�V1	m*J����$PXE�("
����X��*�
�*����X��*b�TX���aQU`�J�X�J&0c
(*�F�[l\2QF
�X�H�0�V�X�QAa-�J�0E�)*,QH"��X*�($TE���)XUT&-�X�Ř�m����KJj(5�����p�X��皙�j;���!e�:<��y�.���Z�m<%϶��7k��&ۮ��ۜoS�R�E�]=9z�Ɠ���㔹�|'E�����o]n#��v�����f��f��ʽŀ��ۃk<��nh6s&޺�v����U��j�b\�ܙ�i�sI�h{�9w�NV�<櫋=���9���܆��V�CT�ol�n�`���Od�����'`��u�.9էr�����آ]���	��g�^VÈ�;���F3a�ƕq��6s�A����\n�ܩYn��\H��ܫ��[vvb)ܾ8鷌�6���r��"�{w�j���{�۵��N� s<c�:PTv؞x��fKn�tc��{;O��a�4%��t��Z���)��l��n���D�k�0G
���̻�M���t^: ��ǳ�i�o���S�X�z<g v��X�t�y���g ������`���� ]V{=�b��8�7:�ܜ���/gs��&z��2�ݸٸ�6�������7hNrf���7�[y]j4(țq�ɀd@Ͳn�u'uы��g2QX!!q���öt���v<��A����q�,�g�;���cx�5��r7P��n۞�׺l��kr�g�Rۦ�g�n(��ìv� ���{ES�;�v�iD-5�)��nݛI�]�Mh6���x��'n�(8��t�7a�]췯	زJ�zM�e2�d��=�-�,�h�[;:�2n��MC��ݎZ��]��X��Tv�
.׮q�s훩x��68&�^:m����n�qq�r=nz{�7��˃^ܻk<&��iNB�����Z�lrWh�vފo=��^N�nո�z�v�2�=@vC���c�c��<y9���`��i�1�����u�;y1�}�;��e HC�n�u��{��S]+��U&������J�m�y���&y��3۵����aqpϡ��)�V�7S��
�:�g��sV��^Lc�r��N�Ru�í��I;v�nv���:���n{>�=�G{0糦�ezM�i����	scn��j�w@v�R+��7n��w��2Ѷ�tp�؞1ń�[�dܻ�·�ۗ���#�Iͺ�r��o�r`ݲT�\uѸ����ݒ�s�M�n�)��z}n���=�JnI�ݸ�q� M�yѷ�H-dyŹ9ݘk<�8���:2�չr�Ӻ��1���ݡi,��fw<�i�,�So��Ϯԇ�^�z� ����"ڛU�Qы-��:ܐ >+z鴀�Qi�TR*�St���t��`Ē��R���}�- __�0f��݀	�z���ڝnF(g}�QJT�Q"�F=�ϙ ���v ��|"����>�!�U�ך�������� ���B����w8;>Ƕxɟ�~�V- ��븋H�����z�^�w�ϒJLʻ	/��|pi|�t�V��k{`ޜ��q~U��{ �=��w_7h ΜmIݹ^�W����-�q�7zЦ��q�q�;u���n����iֶAr��?�?S�ڮ-��7�����>����v ��V1��zsv�7>/�'���|�|݁;��$�A2�b�/�Wia9��||�@�]�����4��b���`(��\Z/[p�(�.�a֋��S٣��S/��98���L�N�i\b�;_�w+S �}wh^vSa�4Fؕ=��Ywo*��0r��	U&�%-�u��v ��y� DW�C��G{�w��.�컰E�my���-�T��D�e�Wy����x ���XA}�����˧5��$�ӛQ�ov�"ԑ��� �*��񝎛��.�Ӟ'�oq[�`%>w�v� ��� ���A*�=��������=��b�j7]��kUg@\�ź�l��s��+���'q1�����ߟ��r$�:G�w}`�"����D	����꽥Oֹ|<�̲K �_�Sd�*�8���`C4�a�+�I��g��󫞮�� �O7<�!���m$I��$�O�w�y%��	��e�")��>�l U��LD):g�n��!���ǟM��؞m�S�Q�q��Z=��_B�̝�«J�N��w����и_{�j�����9.N��z���׳�/3_�#�y�^a@|Wm�i �T[���ATL�
[;���wwc61r���y�N��A�w^�h"
ܿ8` ��뼽�s��1� ���l���)�P�(&S�Ƿ^�����X��3|�nr7�>��� En�8�in�7a+5������5AUR��"��N��:�9q�o=[���z�}�;���ۤ���zt*TQD+����M�"�.��#�{�[�[�(Eg]7�A�	W�*�%E��j�.+N�ݙ� �h�N(~��`Vm��@n�;��JEB3g4ei~��y��2UP4CN���6�Ԓ^�{o>�J	[2���7�E\�"#~yt��{.�H���:U�a�
_�W};�2��V�'5ס�7�.� C�mZs�ԇ��H�}g�a�Ҝ��wM��o�c��	N�����˲FFq8e�w�������e��~I]=�##��b\���tOe�L�r�Y94�$}��K t���T��
[F�]�� v�d�yn��g{��������I�����+��fTS#���L�,Q*I�'fc'd3��L�u���b����.�C�����I�v۰�mY�#WB�%
B��Y��N4����X <�C8;(��s$�k��5$ >��˻	����TR#����:l�=������a��}�~"8��ۘI&o���	��U�ʝ�k��B҃�
bI*b%����Y
��R�I$�y�㒽ޒǻ�t��N�ٛ�wi <��IXb�$�j�S	_������#ޏ��W���{�����;+�� �]�mK�٨*����٭�	_j�DhEU}��6�}��E^���{
ba������='Dg���� nW�@�Ev]85�O�����ŝ����reNy't�K7O,.qG�uX���m����f����Dë9NF�Vn��<<�4nʸ�B�~ �uf����
 rl�9�;7-�q[[��V��ݧ[֝�`6)�3����Q�K���{lh<�d�'g[�\ �;nmֹa�g������۷�q��g�:��r��͆�9��fw]0�6��ې��@�W s���=nբ��ngvy������[`}��޼���>v�O������[l�=6^M�E۵��8V��BѸ��n��䮸\ym�$R�L���!ե˟p�P5l�]� �ͣ�����GG*�
��"���3r�����W�U�~p�?�ޝ�>��S_,������r�H�Dw�*&�fSa��M0�)�l»���?>�׿X|��8 �v]6|'��
3���y�y��$�5��)$�L�L��M�����.�`�	m��ܝ���_���@;)��+��ި\Po�LL�HD��^�݉�o�v�������  �ۯC���]�uzc��D�d��>+��RTn���MDL)&�4�+�û{�\���/np��ez�"�.�A����y�HN���'���FYD�h�A]]�C����x u�v;v`A�C⽼[W/���W����hQ�MW�BK;�u6���� �7w��"��W�3_m��t�@�*z&��L,�X V���}��&B���xo{sϺ��ݠ~6ow{�u��o#���7����������Á�`ʁ�
�=��F�(z{ݷS$��u^�9�;�H:����,�oswk܀ 
ܿ8`n�7`�*�rɚMQ-��9Q��Q3)��/r�`�H37�݀ �_)�Q��=9ί���V��h"#;o��(��@�P
b�HƟ����һ:*���d���ޱpd����fbH$s}�%`燪�{�=�K^�ڻ	)G
���,��]�w��Ă"����8�qckv2N�9��AWn��}�q���Ó�v�7��_�X�3��Hs��c��ל���d���2�G9g���`�cgu�>�{���ɛgr7���
��F��w`�_�?�́�>�}�A����3�.�$���f���$�����.�U~�m"|�����0H ;��wh κl" ��vI�v/ɪ�DǷBq+	����v�"�ݺ�DC@��9WU���UB3����3=����^om��ܯ^O��m<�{����ٕ��;�2�򗷞E3gP�{l]�+�%z����
��A���� ���@ ���l�'�"0p-#M�.���VR[4���Q��Z��V ���h]�O�Ng��2j�L M�˻y�R+�MH�376� 
��dn:�I��w�ᠯfsv�@���@�ϩ�|��5�}�3�H�pi$n�F�@A/	7,6[n��X�0�������;\����g��x��f�>9�n�X ��� /�+���$�f�Ϡ����'��$�������2âY:�K��C���v���*�{[�`�	���0>���?�W�&��6�{��'����� P)M���� ]�z��F�K��U�=nX���l$I_^�U�K�3�=f�b�t��m�׈����^p�� ��ט  �����?Ͷw���������~���LA�8op�Q�S��oG��@��P��"i/�H��
�b)�*�e��,j�YS�Ά�w��k��ږB0N|�����6زv�V�I/��ϝ�&�.I��[�`	K����M��ϛ��ֽF�ti0{2�.��3�=�p��ݚ�zn�f�����*`㳸��^���D�$�$׆g�lx�H:��^�vm�@{��" f���#�9{��{۴�!�>�m +�Q;�$���d{{[�`�r�q:}�~���]��z�� �y�y� �=�wh�=/3Vg�bAוJ���_g
�-�D6^������#s��� A��M����""�=�m����9��Ep�h�b�\�����^v%���#��� 3=�w  F�N����ۃ&�� �^U�Hy�1��%�%�tjϮ��qO��K9�m�6�Iv�y� {��@ �ΝnJIh��k��*������~V(�w�2,U|0���ݼ�.F����r��^�T��Y������s���Qt�!�!<���%vr���rZn�CO!I�
���0IN��������[�la�D�^sq�|:��9���x���_H��>�/;�=m�tݫc1��rsv%�)�<���noah��TTn���c�ۜ=%;��8{u�G�8�3���������g��
��S�<�懫���v�������;����;���k�R�٘��M`�.ɕz��xV;gXt�<GZS]>�/t`���J�=;���ݸѠzxpk�d's�,�w��m������*dO���� ���s���Ӿ����zc�]vSa�o7~Z�ʸ��LL�O�%��C�8}����<�ɵb�$��z�O��g4P	xfgw�&Dڰټ��I}B��k� ��"������;�  'u[��)E�E>w�� 3=�݁����Ct��5T�$�4�Y'_����xVq%�U�c� �kX� ����!��t��{���}�	!��)M�����AC��?�+�I�d�GI�`}ٛ�v�ft�jH>�z�� �R7�c,��_&T���u�	����Y�YC�M��nNѵ� �TE�����1*"I�z�~{w`��+�H ��k�[�m�jo4�U^ܻ� 7:u�J0O���Q!Sh]��=P��g����x䳐F��^S:vR�e�����h6��6�½+v>�@��0�OYQM^[b� o��Cݚ$�Ƨ"{S�����ʯkq�}�լ` S��"#����k�۽�>��U��S�L��m� �O���#�帱i�۱�Ӭ�`"�u7���jMQ���Z3;�~��`m�T�"z��F��>�8`$�Y�v��vk�ǟ g]��?j��Rź�(n�L2v���P���Ց�}em��e�b3�ަƀ ��N""Vo]�O�ꞏk�V�2<�ݜ�I��S�����V�=�.1v��)�Ӹ��Q��m���HExP4�1�	�g[R  �{M0A����}X�������GwmPU��mv�(U(��5�F����$,+�����t���  ��� ]�wh�ݨ���y�eM��G�0O�#��!Sh]��-�4� ��v� J�l�F{��ͧ˃W�v�8��;������]��ݾsQ1��FG�7R>�1��k}w;�����]��������;ג3q��OU��EirG����>ɦj�'G�l/���9�.x}�d�t�u���7Z�(�ic���|p����4]� �Զ��[�ۓ�;�'+�����������U\�ΜD��w�t�Di��/��,>^Ξ<<&��v��`���v�x�^���3w��i8�2�y�Y�v��_!�l勇;]���o���k���ՈYd�O�L�zۓ���-���s)�����J3��ws�5��Z=q�����v�$�����|J~�A�k�V'7RfoOg3�a��� ��Oh���{P�k)�>R��ɔI�e�V�e	v��
V���~M���/ҡI y5�FH^,^�u���%�h��{mD=%ܓ}��O�;�>���۵������f���S$��yY�X�i5��A�~��s3�Pڷ�)yU�[��ED��A͈�.�J���L�]�@�j��R��)�b�=5�Ժ�g�����t�}�d9v�s���ւ�Q��dh���ώ:� s�䅃�؊��{�b�\�=B�|,��jE%����q���r�R�_�̇�#�pҲE�@~d@�S��v�E[^��>O�� @JИ�C��!]�`�Àk:n]����G���w����{����s�`��=����Ɇ-8�4on�Mt�qG������i�#�������}��ܼ�ju��6TΓ��޾^B�Ttj�i��d�����" 4�QH(
1DX,�aR�
�p�	RaTeJ-� ¤P�@�d��$X*VȌSd�%b���"$�X�K�`R,��VE"���R,��[J�U�b3	Ra
��R��0�1EYDAE��aHT�e�a�`k��V�b)�C	QAQ��"��H�+����QU����*���ZS�B*�n1(�E"���8l�E0±Œ��%)V,�
��-A@U1i�B�Ȋ�DU�F�Q"�e�0��(�bŊL!QUb�	�
�" �,���Ʉ-��V�"�1@S	A�V��,+Z�FKl0���U	�b�¥���Vbب��
�H#E$PX4h-k
�ER*ȶث�VR�m�X~��ޯ@@"��� �7��v�^��%8�4��囹-�Fg雚{n�`�����w` �Λf���=������%��U�IHI�|� ��U[�M�=�@ ��93�3�[��c�� �/��{��� ��m�^�v_��ef��WEI|�L��I6(�L"���S�y�s��DW\h^�u�r���>�{�ƒI��DKۮL �7���� 3:�������tdE<���y� �}�wi����$A�2��kD޶����ў��^�rL�s����Λa$���s7�r����$�^�T�ED�Jj)�w{.���#sf�C����Z�q����݁���C�ң�����6o�z�z�.#�=8�u�Qv�	��v��ft߈�]}P��u嘷v����' zA��ˎLZ(?_�W�����T�o��;R_�W��a�~�!����Mܣ����"��峼�����g���O�V<�	N(M)%zZ7r[r]yO��]Q��? +�ۻ������  ���©��f)<L��r�J� ��T�F�\���a�$$6�:�ͳ)�V�	�<b'�ݵ$B�$��+g��λ���ft@ +�<᠌q�o��z���]݀F�η ���*)D�RI3NA]{M0%���=��]��m���� ���l ���w.�r�I�x����s~Vw���5R�P(��맙 ��즙 �V{�]e�<��ٳ�� @$WvS`qɅJU)�SQ.5�7���������@ }���$�&��6D����.�#^8}g6�#�Y-�R���*dM�_]z	k�w��aJ#rn댈��� ���DDf{y���ۨ���o�����FLS���vv�}��pؖ��.�nW�V����˕�v��ܰ'�4a٧��3��nP1�����|Ϗ}P�gqi \�f���6^0Wڭ0X�A�W�l���'a����t냆5݋2ub��ګd���p�r�8�������q>fq7s�p��[���[q���ۇ�&�H8�h��A(Ů��d��ʞۮ�[paܗܒ�M��Y��<t�"l1d�۷7�qu۝��6���\1m�K�e�\�f���#�gg�IUvk�wl�cm�4�v��t��{Y�7X�@�����it�S`�54�Ҙ�I �2���Y���)�A���� @}�������n"׃�Ko� @Μo�	�B���IQS���:�Ղ;�b��}=�J@ =�XȈ��c�"�{�����i|�W*��H�l�Vm*�>�m$�׼�X z�r�6�$������jH1�]�r��N�P(����Φ�{t9�����󘈁n��@ >3�u�������)O�;�!�� ��JU*���mm�ݑ����r=��xzCu@3�M�I&����$�3�u�.��[ۍ��{:3j����H��u�g���xX���[���ό���d�$ݶ&�"+9F(��J
�~�.�m�Dgu� �3�w��򉮓7&5�~�$���v����	WA&�%:{-� ̷yя<�U�:�%�S��ݙG�֍�0o��pۛ��Ԛ�wQ|)�!�P�e�庈;Dn�H�z��[����\]�^�ُI'vm��E����� ]��fJ��È�N��IMQ%U�W���ľ@�;�"�}RO��u��8-��vζ�>�eiT��"�d��xJ�g�/�����Ĝ%N��@����=��lڂ�f<�����D`�gf`I|��� �ȅ�@�fz�����7���}۞���f +������:ܐ q��B����������Ɔ�p���y-�陘t����L��.c	����H6�z�m�>��k�?ym���"7vw�A���r�
��t�e��ywv��9��U+���Dg�((�7����	��WD�W����%wum��"PS�����MȦ��⽷����VY����L[>�rhi����m|�K��ģ��(׶38P�����uE�v3W%+�3��h���oy52�ʬp! }Vom�[�ngz�=��+���*���I>[�{h�	/��>�i}B|�h(�EJ
r����33�f�v���3D��g|�R yu�k�6w�3�8�����|�U�~�?c��W��*�mT7�U�����;��!��	�X`�H���d�w��K�H]�\���Q�~ !APt@����]�հ`�d���q�Lzs��ΎM'x��??;�7��v6��>9t�>D�%��� �޻3��#���{�� I�}�d�|���L�:������\�����LԸ�>����B��+x�y�Y�9#�C*0O}L%I� 9u�b�;���$�}����~eQ�I�{�dozzY!�#�0��t[f��p_�A�Y�,���vjx	 ��~$�oO]�H�k�ު�7k�n�%j�O��y�,���ݖ�ط�ٕ��Q�^�xy`�24>�[��H�e�[�qw�����dX�C_Vu4�=�0F��>J�g�4'ޮ�����H�=vO��}��
�|��diVa��W���wOO|I ����M����u2늢*H��z�1�۰aU��;Z��n�>�G�u�@W'��d�(��rf����������_��	����P���Q����=�.�?7�~�$Mc�?�
�Z0�����Ru�`xm�U{��H=��K�A�k� ~2�}Q`�'�=�	B�6�`,Z����)���{�_���v]ʝw��	������H>�r"D���B��6�9u��:UE]�By��I �{j	���]rK4�{^9��ӷ�,>��L]$PN�l݀o���D���]v�b�W��d���������e��>�������8�^�����gٝҚ�+��}�W�\c���L�3�KI�M/�D�K�g�
2�S��;�;�C��}w�����:Q��'Y�(l�a��	�wE�v^�Nn�i����S�ۮl�'R��ɺ�c!��wJd��F��wn^V�X)�ͫ��ԡ�9�Q�3�k7kt#������g7oO��:����6�+�����LKu���[��&v�1u������h��q;Q�\Qv��gV8�7f���omW�e ��x4pi�V �k� ��
�sX)Lܼ��aB�N��-�#�{[�re�8�nj��a�4*����y��Ai�$�T�v~$�n��'^��	�}�f�w�n� �o�[]��( ���
o��m��~7�Α˷��| ��| _����{�#��6UU�� �<Ƥ~�T�E"Z"���@'�W~��g�M�p]�U�������A'�n��E{��B�jXdЦi�]���v��S"�x��S�~>��� �+7:�	�޺��k�l�k���A��P���%[�DR���&�m�	k{��혪T�$W��Vg�W�۲@$��]��j�]3-�Y�Ѫ@��m7IEUp�ssg���AwY����k[�t�v�Ŷ�m~�~�G�ZH&)�w��r#�$�om�d�!���`�-����o�?L��%I���I�$�S�n��dn��N�w��E烙�;��+�ѳ&��[~�Z��Ƅ�(�U�z��h��8V1���v���T��(�t����[�Or��|��$��ޱ`������N���uD��b�J��Jλ$���z_��I�����1��/ӠO�=�vH'��޻3�G�UMJ��=�κe���{���H���vI?��V���j	W���"�����B��Uw����� ��w���=��@��m�?��O��s����w��|�A�t���m�[q����O=)��Q��N����˳y�$<��#8y����6��͞I/7�/�I&���b]�]5�V�+(���FN��DB�����I��
$�P�^��o(�n���`�H�{ޱdVu��X�9)U����~���ʴ��!�P	Q7;�~$g��$��b�U��ۖ��1�f�m�_u4w�� KX��J�fu�y���n�#��^�h���pE�����pr�"�����=wf띯���x���zX �k:��xGmSE�C)���q�����=3�������	���@��e��?'[r{;Ȃ2�8���B��@84��L05��x�;�N�%��y�o �k�`�vK"�k/{7PC>n/�E+�R������ƚ�v��\��\e��c�//�|�:������B��U����7�P�$�==�vv{��A��鳀$�{�	� |
P�)
5M�`g�pV5<����ed�I��{�fH������lUk}u�2"5�e��j�
��9�"I����� �ɣ� ��G�/�|	�z{�vBƦ�E4�UIJ}/��Vף�8��!�rS��7.�'}=��|T��B*^���e3����شMx^��eTB�ᛢY�h8�p��d�v	�_C�%�z3Wy����cT�as�.��T�%VG�J�$�`EsjW�|3׿~���Oj�\�`g���6{��O�{��޳�O֛�-�U���2F�귊�m6��I�GX�m�wѸƺ�YQ�~~v�����lvM���	������z���ܕډ9��.�����,P�5,2hS4����{��>k²���`��d��^��'�T��|,+8Ӳ�Ƿ�-�J�c:TSdWmt������k��M�;��M�`Gfg�Y�zX'��Ds�)�6U�7��<.?^T}�q9�t�0 �U�͏������߫c�& &�����.��@�H�������v9T�͛�>��|G����� ��cZ��BB��RBB��HH@��HH@�Y!!I��BB����$���$��$$ I?���$�䐐�$��B�����	'd��	%�$��BB����HH@�����$�Y!!I��IO�H@�����$�$$ I?�b��L���ך �� � ���{ϻ ������� @��)T@�x P�/��L��F�Hh���H�e���Q���Ux��{ۧŏI�	 �}��ր���ǰz�=z�Ǖ
��F���Dy���Ȫٽ�T�u�E\�G�ܥ;��67w�:4���    ��JR�dڃA�LL�FC1�J�@      '��U*0C0ba0 O2�LML�   d   �� R��d���4�	�� �M�`@�)�Sjz�S�hlj�jNޞ�zj��\V?�IG�*��?���"�@
*�O؊*+aex~���3�?:?����A� j�B���F� �Dd�s��5\/n������~�WJ|l��9F6u���>9,�E��7�ĩ��y���{iܛ1�U=�t#�Z�C82ْ��b��C�ס�����eCr�X���xBoI�3N8�[��$��Z�"��J�r�����7#GR��k�p̣8�p�%�M݉�N���9�4䳴�q�BV��y2`����!8Y,�%*���XŔ��Q��4N�6B,�H�[XE��5��5��]��V`�u�fJ��;��5>̬���mh�P�T#��m������*3�v�$yz%�I���0��֕�ҥ)��r��7�-�"}"v��G]�n�;ŁK�t�*�	��T(�æ��Ղ�H��Y��ׯLV7lDX̋zk%�c3q`����B��]]cl3VN���4�뿑6�
@��D���cu��YDc���R��IP�xY��h��K�[7)��0��J����o,Y��+V6D,J,A��qj��^ːT���y���7�(�V�:�^&�EPd�f��ng�@�j�݀Hm��Ȋ�J�n�?f� �5t�!�]K������ɺ!K��g�F��m[���֌T]��b��Q�B�m��y/&V ta��Z�!�tf,�N�1m�ܶh]X2��AD/jS"2�
�K~��SS7�䕗F?ے݌��0��[diW������+�;y��F-` �ӛ�哆UQDʼ�*Ed��hg�oV����Z�
�-yy\z�ݺ��.nCE�C3l�NQ�1l�������V�[m�*�	w�M/���F7F���$�,��c�A2l�96� ��h�'�U2���ӋmcL�֪�7�\��j��n���w)gKurF��
&�L��qT��\��v�J�Tj4bkFwv�]���-�HV+У{>�pD�
a$Ōu�������?�~�#�o&��^�ߤ���ry��E�����2 ���(T�
H�H*�H*(���ǉ���ǲ�,r���TV�HZ��
 o�Y=���5������us�����Rf�O���E�n����0��@�O��2��f�Ӹ6�aڸT�0N��x�%���\�<U��I�h��|�e�n��-�Lc������e趫�����Rܙ.����R�sѰ�i��R�#����-�qu�-*.���ͥ/5�P�a`��.�Ӱ�}R��MiR'�B�)��-�T��%�%f��T�rKpP�cm�K0_��BΛ�;�	X	���m*C>�}�ċ����U ȓY�F�:%�Xgb�JZ2X�i��*�^^w��ɺ����΁�	޴�gq��U#2t0i�s�,�	HL���n���ӓ� -���i�U�!�n�&]@��O��7f�Q�dN`o����.��Y� n�y�V>+'u>T���$�ګ,��S%��A<��PR�zE�I]��/D����,��;@ӕ����dA�(��C me�z6����+z���2�B�ZNR����d���gi��k��v�[/s�����I���RJ
�X�L��6.�-9Kf��gbD��Ӥ�y����������Z�/j��FLvE�u@8ҿ����i�U��49�g�rh�9T�HgT'b���yo3f��99zQ</3�3(Ý�m�Ve�**sE������[���#쥻j!���.����D����&Z=�L|�/�F*�=#Ѯ�Q��w�.�1M�U��g�eY9]������U��X�R6�Be���1mvC&"�W ����Ե�<�*�ԈQ��������S.���q����58�ĳͪ��%]�
�A��8���Ɯ�k���7�v
��%a$��c�j�����f yK�`]<��2�=���6�7
�\k�O��Ps.�#jL޶2i��w�їQ�Y��߭�����'؇N2\dJ�md�j��z���h6�(5�6bU�c1�K*Y�[H��B�M�nۜ��Y^9����B8�5�$��&�U��$+<���z��*_��^�,TT���9��v�p��pm�M�Gv�܇c�
T�����Nnh�%�y:;��3����pA���XĬ� Z�,d�e�mv�����&���J��ý���zR㋏8�뭵�5�O�%q`�/ha�v)�`��
�/R{p[�ǰ���P�kbϢk#^�`��{u���v��w��À睕Zn��'��z�����!��t]�#��LEȃtix�ܙ��'Win��2vwl�bĹ�M����9Lnʬ�t�;�G�mm���C����\๱V��S^ffS$�KI��B(�w�瞆��<i]-c;e��QۺX��Bk��;�b箽�;A@�k���8jRX�F�e�%���sa���<+�lY���P��[;�&�V��-/&kN�j�&g=+�cb�k��e�lt�7^Ŷ3�-p"��!R�B�Kn���ѳj[h�i����7��&��@l�e��V�.�UUUUU@�֪���Zs3Y�u���g�lwY0�l���v8����w=w �k�)�-���J5ۃ��Z
��[b H�&���� RE�b �l@��(�F�P ��b M�b�� o�R��.�u�tT[r�k�u.�>�g�L�b���.т󎈐��tR�H�Au��'�f#,/B3D��m�-�JM��Y�vX�J]iGC��dN�@��������CJ����V��9��+!�E���B�Gkm�hK(Mn`С��)�K�����S�'U�8�by�w&��gU�	�)NEfX%zu�X�Z°Z4%��3;-��G��l��D�)��,A�L� �����;@�ku'�Skϙ�v9��p��Gw�ZBd)䬇bѢ�Yע,1��ʳ��tĬ^�է��v���Uw�D�2X��	���܊)a]|���L~�fo��(��TD��g�U��fϤ�>���"l�l��]����G�����#wQ>{�����*=6�>�$��^�$Qx���D LZ�D8݆z��W���ļ�
��׽��swn�{|��b�T�bF���Z)g��jwp�"�:e@=���@	��i�j�`c}Zj&ت�{\�yË]�������j	2K.I!�o2'ZEQɰ�T�Ǉ��^��ʱX�Pb�j��Z�A�T!��*¡�#�U�mAuf�\oN�{]D�tg[
L��Sq�x��Ƴg��$�>��wP�т^ ��!;�e++��b��
V XB��gcRXX��gV�X7dQ�$�4}G�⌙|����j=�_2׳�v����D��*�N�Ъ�mYh�zU���Z0@�ǹ�n�q���Uwmwo�;�Ab�&�c�q��Ϙ>��{����F3sZ���j��l�k�1�#��~}E���/,r]��s)B�p��]���Z�Lb� �+�2ʱx�{QF-7Z*������N�Y��ni{���x/�N�(�v�h��K<%/,�� ���J1]����xX$����'{,J��D$�rci�����+�ȍ�\)p���l�э�J��D��ˆ����(B�Em��-vgs�z�����9�����eH6Mj%e��5�X'~�
�)�=֗�v��.@+�S��'.���.�81tAJ��¬K�Y���>�8:�
]����S��e}#U��iJ��b-���e�K��gǫ�
��ls��}vx�N��m>�����RS/%K�v]�>Y��vl�F���Ѷ��WQv�Obw��V�	Qodk-��=n���LDt�� i�
h@")(��� x%%�/'{�����bL@ j��+�pO[�c�%aZ>����Q��|:�0����"n�"YN?3��۬h��[[0��X�>[\�&�D{k��h�>�zz(�>C+�h�7��0hë��_Ӓ2�$����4�h����o�i��E�YV-�Q�0�GY-E�謭�T��禆R�Be����]o,��ZN����>C��Sp��a�(�⦴&^&���0Q��nZ%����6�n� �s����T*�I��z�,�j��<`�V��Z�߽3M&)�bȢn/�z"�so�0D��O���eM)�|tND�����੘{ڊ^�h@�>"��#Wf���GЄ�*�m�Ͼ����L��.㊸����DY��&�T��³[9J�^�"HA�>UdU�E�������;���
��e��ܒ���w��3�P����xw:��y[/Q?��,{�T k�!;?^'t�^�=r��
�bk{m]��\|Xi�`�t���\��‟p�ǳ�h�����&����"�oj���G=�¦��=�%b ӫU��	P{�GDb06Q������2>��X��˵�杌���z��ei��$2{�p��P*Ⱥu�TfzD&���+@��M.*(U�5�!5��[j3�o����G!�t��	��k�ʐ|��GcT�5�w���1��6��a��W�"c�(�l2;Ʋ���%���F���}c��޺��3�Η�<;�N�x��S7�w�x���V���ن��wî��Wl=�� �w����r[�,c� ` �o!V��z���P��z5H�+s�`������O����I�4I	-T��DYL��I U�*�9~)�ڹ�CB�q�۱m�@=v88��'p�zM���4�,vl�ո�uøȶ�#�,�N�v�xz�\��e���&�.�&B�
K�ዮ�hḼfkInob m�z�e{��A�s�{eņ2���G�m`� �{�Qפ}� p�N�.�Ń<L{v�xb�:�])��
�w�i_~��b�{`7>-*�ҘG؅��q�E�+���S��w�Sr6�ӝ�".�B[�O�Yb]o]�0G}����e栮RH����i��ȉ�y�2��Q�'�OE���8F�_��(��#�{L����U�U��[�k�X�PQ�0��2�ngV���o{ƅPf_���'i�\Q��
a6�w�;��/��RH-�L� �0��*yצn�hjF6� xB�/\Y�Yf��c��X���rR0�q�� ��
m�ڻ�,�f�`��z%�%+$̳�vT��ran!���S�U���V�\L��xF�qm���72��6�#2�������P����"*�~q�юFa�Vk1�M������zwh[���9z
?Q	�
W��ÌBc��T�G��DOirvy�v�=�+���xK�~��˼��a�ۊ��pf2ڟA��*L�[�[�@_U�۵x�NRۊ�g���sSxa��s⪤��<㋤i�%�ڇ97a�-p�s���B!I��Q���=x�f Lf$�&��IOVP���zA� @w����ʅ�bW5��wT�%^����]\�]��Ҹ܇/�����  Q��'������ ���9�TE^8΅X�ͥ�[ﶨ+��F������ �m��t�k �h��UqS["�bG��xXW��̉	���#�^=���89��!=��V�̬��Vg[�XՔ(˷���PIv8P� �������1���l�Y��6��o17��Sd߶��[ ZT�*�U	Di�$h) (�e��*7bI��#��( %R��%�yhʤ����X k��@���0�"�f����`���7m�9�%@B(��:+m�i{��3�`	X'� 7����6@�[�8�� � �E����\A�*`�jg�1H�}��`k�YB"H�h�#�'�Ϣ������u�C6r? ������7�k�q�8�b(�Q�i�6�k��{޸뾻6�)J�m���L�{��qc���77a�E��U+⣵�*����}����xx��R�^�13���96�Gif�vwT�Dj3e��㹺޻vq-�t�	b�?m8�B�t��q��q���r�\��7Z.y|=�{�gRƱ��~T�v$H0،E��{�, �[f�+7�GuSyծ���$g�̑��3���Ȣ?$_�G0�w`ڍ���L����7A�s��P�:���.�����[��"�"�5a�I���&�A1�2X����Gjv ��~��@����F]���=�P�n�3Z�0�:S`*#c�\�%D\JAأw����>n��=I�����+�CJ���r �4E2���pDT+V�㭭�����ED�֤�=p>c�+�רL���+lBV�mG��7+��g��}���bQS+b���#rS{6�T���xq��	dq�Z.�C7�,�Gn�3z�S�o&a�wxyu}�<�(Fm���g.	[�R=�f��.9j�Ļ@�X�T�a֍���M�q_qw'!҃v��v��U��h��xh򇝋��"�m�<���^���
��1�oq	a����c璞xs5�����)J�]S)0@P���V*m�b�
���:0�ϑ��<< q��ʹ���^R r�S5��ׯ�ʴ���J�Xj�.��@������'l��n���[j���$��O=��<��sn=�����B�,���ژ�.�T�:/�1���QX�l��@���o,�Bi	\��V�lț9��Z����CE���0���t�\�m����2TE�&J��ϟi߶��=<���R��{��=��4L;g��RA$n,��Q�M�R+^X�������㾐�1X�?Tz�o��9W�#"�"!������9�>�x8T��*��C��z�J:��ͤ���2�n>���k�Q�ζ�c�!��9��l<Qsc�� �m�2� �m���)5�f�r��ş��&&g9h��TU�N�^�]��x P�*Q��!E�L����m��^���Ť� �P�0�VwČ��a2#�'�Ql��Y1�3<GB4�}P��W@�zn���BӇ�X�u��Y������މ����Ϧ�dv}LLB�T��u�S�{M6(�k����%�c�&�� =qr��RH��5P���ˆ�}�m���F��16$Ut��F��c&A]��-�hr�տ���@�Joӳ��2�Q}���_�:be���ᨆ�C���ljA�5�n��E,���^�>ݽ�o>%T�����Y �Q���S�#���:��䩕��fQ��1%E✤�P#�j7\�U����	Q�C(�BC7ke������0Krq����W��)�d�ݚ5P�fz�G�������X0[j{���W��!+�Tݻ����&�8�}��Ն�.��]����X�8�ַv^�W��M�h.�&h�n�*P���NX����*��.�L�9��Mw��ԣ��Ѐ�؝�3.��{�Nb�@�A>�y8��|7h�<���Q�`U;5��O���<v���{�=�"۰{�O�_l�w�QE5"�� !�/��W;����)G�L��9uv� V�4�]�ϔ(��b�OR91���C����1������U�B�\���~�Z4��DY͠i�"c�ѕ��L-b�O��'�kI�6B�]i��V�������)QH@A��S�1�e�腛���bSl�2�!چڌ������%oT�籓Ga���~�W�s���Lo5�#��=���ܻ�1;j5�uW��x�8������B��"~R�!���f+�X.��gʧ���Y|�!�K'�Gޏ��3�n�+K��r�Q����d(MN�d���ĉm|�q�
�١DP�fOw�vQ�q_{1�b*�C�$	�JG^���o�v��kw�o<���9d��+�q���D�`1�V���P�P���h��#\\�
kkpv���n`�E��&.qY�����UFRDF���yV1�%f�"e�M��*e��������z�9�mI�J.5��ٳ��A���!|�,*g���':�rP��`?n�����3�iu5�X�$O5ܱ�Ղ����1�[�WV�8EM�1$	Ho��"f�4 h�i��p����Hƾ���2q��u���������,>"jw�R����{�IIo]g+`Y�=��ۑT�Xi-�t.X��:���wL�]*�v��m�핿me�K�nsy�C[�nH�@C�v:h�n�]��:���@=�	�32�Q�D�n���3��9��'a=�o:�f�����ؠ�1�j�IЛbX�`��{90nx�a�8��s��979y��D�v�<�pٝ���s��pv�vp��M���YhMM��'m۵6IX
�9v�ueri��t�|:e�c��N�|��mt�`��T�.��yf-uP^l�+�yɛ���ΊA5�����R�ħGNsruvs�����M��=���Ռ�	<X�v�y�3US�}Y⋌�f�>�f��Lb:�Mŋk�u�����x70Y��ݢ�pۋ�z� �;��o�$p51�gH�4��s�+�6C��F߸�u\�Tf�<�YJncP��/���W�/���30u_?�?�AY��'��P���ڏ��4���{IK}=�S�s��3?�u�j�&L}�0z`���1�"�M}y���T��[N��H�5񝍑�7����&��w� �x^)A�����S1`��܍�&O�����%*� ܧ��+ Rw�۸V*t����"(�ф�tu�^�9kz��<�e��0�h�n��s�r^�fmU���H.��#�O��fE�2���7�8��ݗQK�92{w��{��xxt��Ϥ|�Pg����g�Q�����/�B��Hl��b_k�(�T^�u��^x���!;� �I�b���\ґUT�K��$�i�Ϲ��y3��ݙx����R�����L8���L��ce���+��yM� �;�dE��u�jl�<�Z(8
6�V�� :?���8	�2s]��/F��kz�0���6Z�f&�o��Tž�nL�#��ʯ#�T�4Wl�R�����0
$K����dN�ʒp�~�Uz���qxca�ę��we��X�)Æ�Mw^�8(F;a��ʠ�~>��dP�b�z:�5?�0���e�v�U�gVa@bLm�ˠ�,�P五dܼK%�+l�H�΀� �@�L`G���J�y��'9T]m�p�y����M�]�b�
$��L�PRd��B�J �!6$��(��B �rq�e����c��y|n�.e�A��%����7��I��10bH�
����7ܲ����V��JZ�ZG��f�^vϳ�x�u#��I>c�-�6�n�n��*�,�n�^&�,��W��ϐ\0�t��5��{�u�oi���E�u5�j]�t%�p!K4f6�%DsWd���v��W���?L�{�¢�*�_7�ZI�Q-ɒ���'	���s�]zW`-�0r ��E/z�V�vв.�-�t���)_��R�j�C7��P�_z; Y��)�~Y�JO�'�����f�Y�^�EM�>WP[���z�]�٧�w/�����}s^s�k���.�Akfo(�%uy��AH{�wyS��W3W�UB������bHT�j
�!~}k�PּǛr�b�RFՊ"ZZ�qRӋZdX�]L���Bl��e_	=��skI�Z鳺��y1i����$�q�2�e�$�ܧ쳧��Y$TzWs�N99��t�+������,ʆ��j��s���\�Q7���c.�oN�b�K��x- \�cI�\%1�U"h�f�L�(8��ٹ0V�n�_��PM�Q�l�I����q�\\գ�;��w�ޚ"�\�^9c��FW�*�xlkm��ĞF��*��:E;wq{!��닛����朋d=�1nð3nᜰm5����9\ݾ���v��-��S�Y���
cl܊4u@%Tw���N�{r!��<��$jL6�D4��1�TM��8�d^M���;� ;�8Gnt��m���6��/����h�ˎM%�̎`:�
<����Hx�����)�n�+��	�]��2�P���B\�O@XG=.���m<��#�۶�%緞ٻE�c��d}��#���3���	l��3`ׄ+���4^$P��8�U��3��1��ݡ�4Y���G"(	D��o�}��ެ�T�ov&eW0[!C����X��)�m���t�yr�ה�e���
@����^��>�o�&�8ᑎF��3;��5}�J
Ys��2G=2��pR8o
��"-[��B��&c{�Nr�����U��/B��7Wa��\���3Փ��%I���
��z���[ƥ �7�+b��^����G��@T1S��o��}ï3� >E���؆˅�������	�)�;��Z�i0�#���4�4E�BH��u4�H�0[�D���=yD�IH��:��U�l��昿x���h<�}Aybݍ�@�_C>gE�AJ���_v�'�����T��dg9n�f���H7\6�4'O<l��[Ai��9V����Ӽ�vo�T�$OwK�^
wF0�&�ӗew?2n)�b�|�VQ쭖&�$e����O7�3�����o��5��{�'�jV���Lo�����j�6�c���r�R̅ ��ˣJ���>�=������S������f;9ӔZ)(a����A��ci契q�N�'�i�#T�-Y�mE��ή�H��*��F����LbڮSR�;�{�{�1q"���:�9��pOA�檾��-VU�0�r+M�����m�(f��W3�vK�g]��J[{i	����g
��;�`�Y`���ݹ"�oo4댧�/	�t0�+ݖ�OtATE6���@�pbA��DM'BAQ�Q�`���	E �Ҿ[벘��j�C4(�[j>����6d$i���-��즛\|iŲ��.�8b��v�MӤQs/R��tH���N�;���\�Q�D�!F���Me�m��@�6�˂� �\��DY��\5�����4�����4aեz�J(�i�m�u��jf�ǭڡ��{D٭�` ��7Bzouѩ�d|V�Gf^�Aψ�� ��d�O�{T���*�@$�˝�{Ʉi�i�U�m�-ʇ��S�ę[��d�&ȓ�")	5j!HI��y��zVc�,�"��<��X#d� 
�-����[�@��<ug=��e��4y�4��������5����Y�Q���\�E���]�X�F�Y��{��Й��9�:�;�@��X&"�]�@��"�`�;���y���f���v�	�tvl�������њ
�u�P��L��L���0���*��Ycab��͉l |ܫ�H�J̽]h�V�����n�Atض%��k��y�Qչ����$�d�E<!J�5�}�q�� p��Z!J��:Е��٣��h��{Ƭ��lX`��YXS��-'28I�w#�G��ڀ�/mKuXS![�d+��]���ɱfU�͵�E�aX@@$]�fi� �ke`�Y�kː����^�o��I���'�D�ݕ�P�mZ�uWL*�=��X �
%�~�-޻~�9�]��8R舓�"5d�RTh�m���i�,��XU�L���k�t�W����
v�X���6����k�䖕>'��=���I�*T�I$��Q[J<�`E�{ҝ�Wv�}!&_R��\���:�_3���s/������ФDBёU.X�.���!��<c|r�94��N�h������i6�?�um����Mé���?J�C�,u�mzu�i�g:�f�ձ���PӘR��tƍ��E���-�߳��`�EP��U��֌�Kc���%�Ӯ��?��A�O�
?^6��X;~g�����(��(�������w�H;�m�5c��/�Fy�00�d��Š����U�l�t�p>�0�r�����[ȃ��y,��lN/������!,a��B���p���$Sl�+�H�k{~�4�	�p����Q^.@��3��uE�����A��Ӫ\9}�7�������g�=KM>J8��hEq��e�Rr�r���͌���Fy՞@S�?_}y���x=ĘNk�?���j�V⇙�������AEz�f�����N8Mup�bC�ҎOB=�<�W����[����\O*R��Rp�z��
�������W!���HF�6lN�	��)��*�.
^��2�[��&mR�I|�C���D�M�1���(?�+�`��<OM��N���;���I�����~G������p:��z�X˿�8ޙ���bs;��~��y�qҖ���������o<t��4>	TR�^�5I�PQZ_�>ձ�}�m�s��/��N/0lrOw�B9�G���,�����>������w�����Mlh��9��������fn�ӯ�%�Wu̦�=4
!ѳ˘d:H�N��V���|��n0H������:Pz����::�y ��h��Ґ2���ˌ3-.�C[�ϕ��)Ȅ��?"��ߊ;�t�]��BA+��p