BZh91AY&SY����ߔpy����߰����  aR^|(    P@��)��� P���IH�x�� �%B��)E )D�@T���Q@P�BT�IW� t  �@ 	RAJp}�p(;uK  ����(�n7JWǦ����}�w�מwov�st{�EsG�y4�޽�w��{������5�u  x�'8h���_}�R�8���P��C��t�ؠ��+����}��� o`�}>�� ހ�*( ��{������ w��{+�oPN;���Wtܽsݸyh����Iޠm�5\���Fq��G^��z�^�-����vꫝ��k9�)ު��`=���u^g��� /= �K9��Ǩ�5OG.�Y.��Aw��^�K_wݤ��<�s��g��A]ꞻ��{ ���r㻜ֻ�t�ށ����ג�{�/3�����z��vw{�zkѺg&���� @  � wp*������;i֫�{�gP8��=��Wv<�g����=opn��֜ x�oL�uNq�׫��^V���oo�׾]���7���w���nm�n;�i� 0  ��7OzSop�n8���={��� ����{oy�{�׳{4]�x�l��k� ��;��<��Ǽ��]�������X�o,�������n�/6r5�m{՝�:�                       �( $  �=	�IR��A�Fb  `��j~�D��(�0i�&  �224�M����T�� �      I��L�J�@Ɉ4��40�2@MTDhLMLe4bS�)���P��L���‪��i��*�L=@�0�  ��# hy��O��p���t�sVrqqWn��ㆹ�]�t�k���v:�������R��~��6ëc��6����o���3a�u�t����O���������u<\����
��n�fl-����[n�K�W�'\l͇�gj��hۼ��*��3�c�c���|�{|���?��Gw��p�L��c�fK�c�1���<����wQ�#m���T�F�������D_j:�6�#z�����"�����u���"�����q� c:;\ec,C�L��c�Dmڈ��h��T�����Dm��#Quii�����]E"8�Ti�|�DD�E����6�DI]Z:�O�"��=K���ݫ�����">�H�����]DDD�D[H�uG���.=�""7+�DD��DCoT���Qy�Tq���|�Dz�m֓�6��Gw*�S����Z����#i�um�R-���F�"!��ڑ~DF�H��4�"���z�Du����6�""�D�墑�F�Fԏ"+�"=G�D[q#�֋�E#h���q����r�W��H�D�z�"+qp��<�������#���z��ֈ�4��8�t���z���DZ)Q�Dm<�6R�Z#H��O8�G^�)�"";u���-nE#�����U�R"'��"6��Q8�W�Oj=DDEu�DG����Q��u�DF��U"4���u�O-5P��"�Di�������u����"4�yDDD�DF�#�DW�"9=F��}�6���Qn���b"6����֍"5ʈ�"/�DDwh�H����<����DG��u��8�DF��DO.+��ۈ�Q�O#���"��ґ�<��EDDDG;QKD_�zDF�͢"#��DCi��H���z��e�c)&`�1ұc޸ڢ"!�#�ׯb"#�N.���h�#Q�R#��V��"O"""'��B=F��DG���DF�Q�+����Di��TDG���F�"">�U""=�iE�DDw�uh�#q��)�Q/h����!�^�DC��#��G"#H���)��N&i��x�E$g#GJM�y%w���I�V�N$Q|�I�S�Y��sN�2F�0c;�e$�Ȟ�"""���=MTH�"�_4��Y�uuh���'��'j,���5Q�"-%uh��W�K����WQ�{Q�"5UH���E�"=���Dm;ZDz�%�GQO#��hO�>Dl�DG�BJ�h�����Ԯ���9T���!ʨ�""r�8����Dq�N#jD{�}���#H�ڎ���1�)��Tn\���Ria�C�$�:=H�t��i3Ftf5�	�>2�HǊ�,bmi��4c f���te�MI ��b��7����_:A�ɤ���.��2���qH�/�tc&1�S0��шc��iM!�}U�1�� �1���z�E�N����Ȥ���^�uj}Yݨ�+ϑ�|ӜF�F��bc4f�1��,���@��cVP��GiC�3Fh�h��V2�ۅC ��L�(ҡtc(v�e���c4Ĭ���Lc�Q>aC�1��Bc�X�2Z���t��U���$|��DF�ʤD��✄Z:��1��c4�Ic)�Y�Q�������+�{Q��t�a�F�QFp���c�Ld�ԣ�+ڈ����D_j:�6�G���ZDO#�DG~��G��H����%���"#o�uKF�DF�*�������G��ҩ�E{Q��:���h��5\R"&1�1�o�=F��m����)�D�$f9LcƖш`�`Ʒ�����*�OV�#Q8��U""'*#H�u��D�qjF��Q7_"#i����8�V�G�����<��ꈏQ*�">GQ^iڈ���R""r�4���DG:��+֚DZn�"6�yբ"�u�S��H���h��#��Du��U֑ڎ���j�#H�&��ר���z������j-u���DDq�T��|��"9u��[�D_���gV��FtM!�gF1��f,0�Lfp���K�c����$���;I�f񌡕*>�H�%,b/eE�2(��f����4�"�t�Ti�4��ڄE%�ֈ�z�Q�r��JR�0C���J:���=X�
[��Fi�V�d�i1�#�TR=F��|��">O">DO���"=}��DDD}*-O.�""7U󨏞��DDm��}]c�P�eB��'��n�ަY:A&!�A�B�Ac%��،ek-��$P3
����t�#4�5�,�b������0�X��1ꈉ�""j�NDZy�Ȉ�]k�d�T:9H�]�FY��r��aјa�YCU�@�o�4�����h���ғͩ��"���km��-.���J�$�4���&����6��K�ǩ�¸�1�UR�(��b0d��:ImYd�}L�ǩ��$��cզ���$c��Ι��3��c&Q���3%2�Hǉ�3���1��5_" t��`�3M(�#�2�ܪDK�����Z"]|����f2��3a2��L�FJPY�TDDu�)��ڈ�����"-�Di�""=�DF����b"#o�R#H�j�""8�����GZ"#�����Q~G#qm�������4���GȊvZ"7Dz҉�F�>��#k��ȋDu��4�E�DDD_V�Di�G>{�i�Qh�"#{Z""q��F֎�-ʥ�D|�;h�i�#���|ߑ��&�6���kڴiW_4�=Dʡ�cGa`�2K�!����R/uDoȎ"8��T#H��F��k������qh����#��iq:�|�H��h���j""���c���GH��1��3�0Oc/�1�|�m�Duv:�׫����o�D[���^����4�b=q�oc�R#nŤq��W�kUh�=��}�E4��]z��m��Dm�|�Ƒjj��Gb��s�/L�����"N�t�le�^�0ޝH��U�C(0�ʣ�Yl���:2��K�h�t�I11yE>�n=k��m������F�t�:n�f��%":_ ]Hbn�:�GF��Iʈ�y8�D�z�v)qq�D��"���d��0�Ғ t�tL���C�e�i�]>m�ԤDq�"4�+Ȏ>G�G=G6�)�򶵖TD{�=#h�ԕH�&���_"ϭE@�J�0\a��DAD��(�G�1�S/#�i1�)I�"6����=r�寈��"'k�����D��6��*���Qtz��(��hgF3���3%6�jNTin�h��r�=Zy+�֓u�Di9]t��""}Q�Ge!�p�SI1�S �̅#IV�C�k�3�#�&2JISHc4c O_ܬ�2��ʀEp��D/����y��;,fO�"+��L�K��t�_鉚Yj!E���w)X�ױ�ߦ�J=�3K��B����]T&�}=^�=���[�Ά��^×�{��a�,;�su\r���p��G��i�����*�����>jw=��k��g0y��̥�n��fRwU�qh����{��c��)��ʜ��~܍1'�;�^�&7{�=�v.�&��U��C��S��P����r�y޹�ϻ��Z����y�ݗs=��y��w�u䖙盧JW�߳�f��،n]�U���Q3�]R�}��ۭf;R����:����_TEق�����f��Jke�u�=�`�7���=��W~�?z��G�my��g����񞝻��|7�w%���=�Ŷ�uI�\;��J��Ȭ����v�1g�뙣K�߾���a���v�65�7<����V���Ǒ����_}���.�d�5߯���^����Οl������u�Q�]���L�n�(�˙�e�;sk��ewzujk��+�m��n�6f�.nk0<�;ٟnC)�Űf���n}�����5�=o>�Wͬ�m)�ƽrn�&���L=�Y\���S4k�ü�
��ƻ֮�n~Ǚ�_�o���$��;�{��MN�5�;�§��\���ӽֳ�1�P������o�{���5��0rn��h{�M�iyҝ3�ŏs:\]P�fsLȞ�ZX��q�MM]��z�r}�ۇ��g �t���=���a�w�M���s�y�0��@�.�~Y=���#�g�2d���{���_OnϷ2��q�~�M�nf{�2}��������쟦B��+����������O[<�e�	���xܯ�=��/|wYs�S>��l�]>e��%���z�.�Ԣe\��u8��`듴Krŉ&�6qN��o���j����'��db]9��I4&��R�{�=�W����ih�Oj��F�]�oW��ި��ڒ�����/��ۘ�,'n|���k�?�y?�)Y�9Nw?�~���z�=vZ����ϻ���E����k÷uY�d۞���ӿt������9�Ǉ������/�0�Y��;���.�R�"�s=�Q�1)f^��L��
F�z.���x�e�d����3��n����qB}>Ҙ���Z~�\����O�M�?&z��L�w3��;�U�8�1�#�h�k�~��u�5��s���;7{]����/{���gS���ʱy�r�9�Trbt�3=�\�]���f����b���t3����~��'I?��~��In�oL�7nN������=��6W��Ð�%2]�qˏ��9��{��ٚ�ˈ{�S樬�^sن���A��<+^n�z��Um�33s�vo{:e�ٛ��-�r~��q��D>�}پ �!J)5�ȷa��ߍ_��<�����1,��˅}���uw2j}Qkt��,/�ٿs�e��w��������HS;g��ý'd�ϵ����w��g�bq��S������݂��f�g����w��t������̽�=��4�������	 �2�^�?�����\����Y\���>����{��w�7�O�5X�����pN�Sk/]a���2�{����Z�V�'�}�^���~�?^=b�Q��m��]e��_��g�C��RYu�٨�doЛf�������@_?HJ���>�d���q1���	��٘ʶ�s&fOn͑���|}��&�%�N�z���{���N��ݵ鳧s�v��q��i���O�{wq���>mMjC��n.��̵ek�Yu���2N�f����ߝ�H'H����Zh���,���}?k,z�+�M�;�ڤZ'c�[;+^cYs5�`���ͮ��o�=C'�=���t�ر_a��(�jz���%�x��{{O��K.vt����I�j.�m��$%��B̟���Dgvߒj�Y�����fe���=�z�Rz:=����h;��}пo�^ߤ*뻙�ʯr ����p�1A}����vۙ�ݭ��r]�,�<��S�xCS:�����l�ۺSR�������Tj&5�~���_J{��s���c���˩��*�{Ќ�Q��^w��]˖���Ig~��̈́�^^���O�+Oϳ��_+���������讞��O1��3[�Q5�n<��ʝ#׉�߼�2��k��X�zsw4����2��t��<��`훹��&>������I%�yai�o�]��{373�FWӟ�Z����۟{�PɤMӞ����ޓG�^�Y}uζ�٘��v���8w��:���o}��w���:���ܙ��������_d�z��r,�~�������H��=�Ǯӧw��k^��e��i�6���Yܽ��_�]��p��ȼL3������s�Y������������Ђ�m��m�|=�ҫ���ww17�&�nfά�vw�{�n�:�^b��f����w��uf}M��R��3��Q=�Q*;Q��c��9N����N��>���ޫ�[|E�����Ε��fU��yUTIW[j:�}O�}7f���%ܡ�>�XI͖ݓ1y��}�c_8Q��g��žR��4��pZ:.g������<{���ed����M룆�$��K}�`��L�Ǐs�����vɊ߷E<m�YW��M��F	����]���6c�>�����2���g{��O�O�ό��ǅ:w��;;���dG�31^���<�QF�
�5SW
'�&oo;"��3i�O�}���n�y���CDm�I&�x*��(�ݓ���oE;ۻ�9!���Y�<ws:�j�nv	��{��엧�o
��}�E��h�=fY^<�l�����������G;�����ۙ�\;H�J���aC�9�If�RSk{����t<���&k����g^-��t&aHw�3��s��K�s}崳����ܯ'��O�D���kk���L�[ߏ��;���=ޔ�ۇt�yc�y�y�%�0Z��v"�*+uKP�t�5*�����\ww��xn����.�4{V�﫴q垾�|����޽�ænm�o�+�,��ٞ5g��m�]���]b�����+����,��d���0~�;���vBR�/uvL�Ǜ(�=�_f���)��I����y�uw�d5g���&I���g����z�r����$��l���c�=�������M˹�o��-V��Z�X�N���Z�W_7�I���-���2��<P��T�ٻ�پ��fvw�o�!�w.l�*:�9�j"�iw���kF��h��:gǻѶ̛4����͛g`�ʮ>e�X��_�}�gs�e�Y�|s^�����5����3왓�7}>��i�+�=s
f'zN�ݖ^ߧ��~?{C��_�uZ�k���k3����Զ����-0���~ɽ�~�g��&p��}��C�_S�i.��.zE\�7���9ܸf����jl1w���S��ӣS.�|�����;VD��ӫ(��l뜔Nd�1b��.l�dE����f�ę����Wj*s� ��SK�_�=����g��y�K�<�2E�w ���v~��o��;�
��)��}3�{���^or�k�~��M�gg����;r����W��q�;�G$��W1� �=A�ǕoY�9W���ɢ���t��	<������ǖ��[���$�������aqc~/{��0��Ͻ$�C>}ǝ[���g�c�<��C�ÍRc�������g݇��Ӽ:L�J�����V�wQ.jmUM�iBד����\���S�Nio{���c�K2��Ӥ;=���W�Y_ƟU���W�g�����O�r�f��ow-mv�3+o��ާ��u�ǻ�C��?ޒ�}�={����I���ۮ,F{!�z�C�b�O������~��37�\jY�����U�n���i�9�w=�~�|�aI~ܳߏ۾������=}+]ݿ<�S�����l����i�خ��Y�M����wl�g�_���7��L1`ϛﻖ������|8;�iq���;��D
gr�S,w6~�'fٛ3��R�=�{�ܛZ��c��Y7��gZ����wZ꾫���ߺS~��^�Z��#׺�J��ʥ���퟉�L��k߳v�	ܞ��0;,����a�{����ǈ�x��׏��N}�f���Ewb�;[�=Uֱ���9��6�Wς�N�3s"��>�l�}��t���\���h�S
�!�8o�.���BD~����7��������u�>6u��^�'�:y�������f������/~���lfl8ֺ�Ҷ�[��V�	��e�պ0��6�.�Xh]KM�԰���b>��muS.�^�@���r�`�2��r�]J�+e��ⲗ��8��-��ך�34��t�C�,��k1P�v�Ƅ�:��<g�JX-MD5B͠ܐvv��;`���8���M,ƥ���+?�fh�T���TT4�����p��]-�a�����&H̲���[,��Tv�T�Ŗ�v�L)IB�ʼ��8�.�m6�ip7�qt��;cCc���w�oSicX7Fˮ�j�P�5�Z��M�ץ�0��q=��l���l��b���[wSm���m�Ԍ8�L�h��g��OKp묪X�L,Ԏ�m��*iCY0���e���5�`YHf[����][��_���(���iw3����5�i�i.Im,�c�*j.)�R0�3/.l�0�m)Iv�X[�쇬=zZPx�]M�U��v�iRb��A&��X�ٖ��� ��f�v�kc� 
�����*(�,�	�(8���(V�E����R[4��ôH��K.��]H&u2Cs�Z[)Zٓ�s�^u��=���2�6�
0ؿn�������
��)�\B�\�[�u�]��������nn�7b�A-��	K,4T�u�]�.��;}|w�`�{|D�t�[�M���;eҗT5�Y�T��j���V*�]�Q�1T��V�v̈́�4&h�J��t-�$��4],Y�k�������J�"��4���?��k�h^�"�S�����]�j��@�p�:�k���F�c(�a��v$�Y}3qu�TE���8A�e�Aפ0���.�d��:�ca�F�`~/���1�����t�kˬ�15��N&�V	1íJ�%�"KJ�k��v��{˽2��2D������5�����; �g�~Y�hYs��bm��Բ���e"@�EM͚���1�bM�R��Sh9V�sqi+sS�f�kj�r�s���`�n��y��2G�c]+2�L�s�&�Ъ��[��j��KU`��-p/�Y���3��A����C4e��!pU�,�M��ֵm1�k[��m�nz��o"aJ䖕0u")������N���D���{�/�E�v��u�(P�)H��a�/s1\,���٘�U9��p�e�w숉�-�)Z�j9 ��s��ٞ�>-�٢��lu�Z,L�p�s��ɫMu��./��5$�F`�F֥+Z��im��[3lZi�],)�IwVJ�Vb�Mض%���<��hEc�Z�8��c��ku�Z�w������&���.񡬴�vi��+V@fq��X�5���eT�+D,�:4Uk���V
v%�o��|��n�K51	!vLR	mU4+���Z��7��ƍLB\Z��|�E�}��qxH>�ݺ��>�������Ԏ}uͳ<|<|<���N��cxm��k�}-?�z;����o=��q�z8�b����sa��d�a[ZF̭���.9�z���=������m��i��6��i��o[M��m��o��M�-�m��m��m��m���m���x�m��m6ܶ�oicp�m�����m�m��7������m�cm��m�m��1��m�RI$���)�R�x�Uyᶭ�w�p�8�ۍb���b��l�mAM�ۋ� Q��I��/l	Ya���~�=�y�m�m�ձ���m�m�m��ۖ�n��m���m��ۦ�t�o��-�ݶܶ�e��}m�m�M����t�o�m&��m����m���m��>����o��M�-�ݶ�}m�m�m����m�pj�G�Hm��B2�!&2V��ߞ��6�}m�m�m�ަ�m��u��m�nm��m��z�m��7��[n�m��m��z�m��-�o�rۈ��p�m�m6�m�m�m�uUO���o��m�nm��m�$�$�I'��^
�<y+Ǟ*��耤�[$���0���ل�-��8����Q����$w����)%I�f�E	*���&����XUAAAb�,*VDaĺk�X���d�O̕ (�X���O��ohٛ�J�ç����?��ο��k�=(������󔈈DDDDDR�Du[�u�#�E�#�]B��#�8�O�>B#�DDDDDi���":�"#��4�"�E#����먈�H�DDE�")i�>G]E����-HZ��Dq�Di�Z"6���M4�""6�"#h�G��Q�ֈ�ִ!H�-R"#H[��p�G���ޢ"�[�:�V��"#��]u�]u�\DY�DDG�E"#OQ#���Du��4�ͩi"�q�^�"#�0��\��� �c�*�"�HS4��hҕ�읕��Gd[����0h��5�k��٪�Kv� ��f�ZƎԊ�m%�Ƞo�[�e|&LL~>g�a�Wƨ�II$`Ț���\)�(��f0�]�h�W�&Z4&Z�:�&�Sr6�(�(c����޵��B|��zWx4�-�K�>�ހY�U�uaZ���,T�=�kk��ٝ$��L[#Z�K�n2X(��"ؙR���	�6���eT���Ymv؍��q�6��lܠ�v0���+�SRcR���Xp�#wf�(�*(	n)AWS+�3Ch�������s!
�&��c����bjͳ���%�&#�n��r�ݠ�ٚ^q�]lV�:�Xd���$,�s7��-kP9�YDV�W�
� ԢA��[�k��}0���=f�))q�^,&��#�����q�,��@AP�ERh�L�ɐ��Ph:�:4*����z�)�����1���-�q0�����+m�Ҭ5Ԗh���-�mq2�˳ָK������V�cV["8�<�7��#�	f�p��GE�s�2�6���ȥ��إ���5��v��n*@�����&|4fL�r!Ԣ���
�e�oe�����?
���җv�ݜQ���x�ŮZ��,�U�QF��쵠xb|(F�xeփ�.���k.��(���p����?6�owi���s� �{��efI$���{�����ٙ�̬�$�w��oz�<<�Þ|�c1q����DG��m�O^��˿�~}]�j�ԺjeQ��zYP�>׉��� 8�G�P�+h�ƻk�6�[�̄��q�H\�ە���u���}�\�/d�f�D0,j�!�~x�-%��:&�nm�%vŻ�W�{T�Y�ـ�7����+j �V�H���� ^%ƓX\+I6����D��i\��g����xϖ��Ї�=?(9�n��-�S	5Ӵy᳇OC�����Z��ѡ6`�x��9\��zYF��	��
$,ء�MB�,���N;󅙭a��92p��蟵�A76e)����Hm�i�]4�k%�Y�1�r���sjo�y
��:%�+��H�t�Ԥ���1���q��D#���GQ�d:Q%i���S��I$qp�X~0��#��S�Ψ"����͔�̊r0��r?������h�7\U
���Uhgf�肙в�nȚ �MEK�(\� ��2lG����4����W4��Ǎ��L�<��]�5��tH"RJ����Aժ�(�&�QT%��򉯗yZ.��H��'Ū�<���K�]:l�9z�����1%	�a�2�3Fi�>DB:�>Du�|��zѣG�E
�3-�ֲ�*���T���BhFk���&�yfcf�$&�M}��ʹ�H��j3�b�I0�"s\�vP��	�G��LFgz}�:�"�e�WS��� �� ���A���--J�d�� �"�z��N�
"�S�p��-),7�Η��,�29\&o9Ț�ϳ�+�TUb�Պs齎U�Go���CG��~8o�e��P�p�����
Ç'�(�Ժh�4��8��D#���GQG�)�QUV���/X�� ��T�B�
fM0b�I��$¡���#x�p���'�����㔦�[�˚�JK�*F��D�\�	��GZbjV��Ľ/ʮ�p5H�����h7���
��ڝX���,����L<�z�58{s�33�!t��D�P֥P#;�&9VI�.2V�a��#��"	�0�<0��<Oݻ�e����=��vz��p[�`jJa�f�6t��采Q�1�1����DDq!%��3M2�_}k�v�9�H>t�}�������&/�Ϗb2t����%����6�2�*Qy�l�5��h�s �`4�@KM��
V�\k�E��Ik1�&4�qcMkiH�)�rZ�x�uP�l��*��#�lr7]M��qD��m6����W
�4`����3���96!��5����~�7��Z~<Z5�dM�WU]>c�WN�qR�g��Mщ6aӧz�����pԝL)����Z崻7����HG��&��x!��n�P��V�f��_�����rN�xT.i=#W8�o9ըK�>���CDr(�W��X)��A��"�M��t?.ɇ`�����G��e�E4�U����X�q�"�Q�#���#��֞�O���U�<��%N����I%@�1���U��ht��|��g�)?u1b����'
�+R��˪���TKVb�d0�����{��х�%/��SF����0)���Ge7} (��x��>�X�-O�~M�MU_���=p��ʚw�uX���8�Y�HeɊƭC����=<��iMc=2"������Ȃ'®3y�$ �	4��\��"-?j��Q�:֕�Dv�����>��i֚F،q�ȈG]G�3F1���@#�Q\)�"�	E:�UA�0r&��ꛊ)iUva�
���\��B����=0K���M2�ML:R��BM(�y�h���$�9���zbbP��X�0\�m+y� p��Y]#�u�mWg�kV�\"�*L�H����g�HiBɵT�*R�������of�<)ͯL4jw��$!��7�K��mL4"y��7"����6Y�g�n�����p�N�	&�Gh@A%��Q��DDS���GQ�G��m�OU_{�(��h�� �O���|!"� 틁(�%�*��x�{a�1���#+Z��ƽ\y����6Z�sb�X�n�S��*wK���p?N��8�ǖ�zR�	2S�3�-��p�<����HV n��ZSx��0��/�O�5=7?&䒜<6ady㻘e�6�f_�����y�t��>T�.I� f���4�0�t��h��I!Gk��r�<�e��?=�t�OX��1���u�ζ�B�������I �D��˳ٛ�������d���G�XI�R�1&۬�䶠��_��!�.��-��Y�-�hD�V5�%��]IN�����c{jV��R5%Q��R�l�0J��� I�.�nS����V�r5(*��kG^��4I���s�4�`���a'��+"fg9ѝ#���ؼQЂ�uMD*M��a �t$�ӊ �m�<m�<����Ot3�	6!�����m=ٰ���Mh�4sd�=�K�� >�h�ʎ�Ә`p��Hh�!�m�0���F�]d�e�yZ�
���)Z�rX��#a3|��_6��D�gi�������a���GN���쭔�OR&�oF:��GX㏘����|�јif� EP���1ȉI$	��,�فӾ�h<�S�y�}�qٜ���"%�(AuU�+��4�KE�{G�d���$����Á���y�^S���(�4�9���uؒb`�(�P�JҀ�p0�� 2P���qwU��f��E��"��H���	�=���/��P�h�L*S�~�}�y83�=�N����u]<6د5������߬��h�����G����O�8g�/�ʊ±��.��V/�b��]U1x��F/m0�1x��ڱX�����Z���M[��)��{~~k_U�W��k�����c�^1x�ⱋ��k�1�b��V+�^1Ʊ��/k^#�/��8�in���m"������/H�F/�X�"�XűZr꘭�x���U+�c�U�t�ұ^��b��ʬ^طU��Y���^�b��c�1�b�bب����k�/�b�c�����b���������Ɩ��l]+J�.Պ�z�4�W��bدT[▯0�V+j�R�WUL]+��L^+n��b����5X�b��+J�.4�X���1��~jѦ1�b�X����X���+*��|�5�^��.ؼV+m��+��u���)�χ��^�ah�vR��S��_-zV*ؾ1{b�H�8�VUb���8]�����Л�c��iu���k���j��8������] b�ͼ�.���|��ў��B{�s�y��9��5#D
��j��b��7���:�v��N]M�IDw�HOe�Վ"=#�}^w$� � ��0Z�(��ӑ�晃�B�q�eIզ�%�69��[��oviƦť>��y>���음��dX�g�Ŀ�9����{�LG��y�;�;z�6�����wW���z}�������g�뻮���z����ffw��f}���燧�i��G]|�":�Q�#�㯝c�-��6sLÒ����P@�2� zXCbB���wϷ�2�)���B`!&��$����L�Ce�`l���D@�z�$q̀Qs���q#�޿����'�j������RH*�,�(R����C�:$�M�um�$��C%��Ʒ7���0ӽ�r�l����4����}�2���8P�rn�Q�p �s��ؾ(���I�O�%M�)�[	�$�Tzx'{f��s�ND�J Y�"h#�'�pd(��ѐ6~�{�	$S�!�� ����|�<��T�ã<�LE;� T�'�x�r����~�|5 ���� Ȉ��8�@��0�O��4y2A�M!?F\)>lI� ��l��ғ���S�T��,�=~|���믑�\[��뎾q����m6��Ge!44E'�L�*$?O�$�&���Ե)�Q49���C���6C�[tgc��k�O��,'�0��&�DCܢ$.K�BK���;c((�]`[LJ�i��˳�0��ͯ{��e�0����D���Mw�������h�:W���h�!�C=�LI>�Ρm�Qt�2��um�Z�<O?-��盒��gғ��	����Ƴ5��2O���(�P�9�4l@���CYVuC�x���(A^~[?@�}]�!=I��C��~��[h�IRO��P��'�,)�A a@	������$I�@�$=6RhM���9��[�5	Ĕ`H �8	�@�(~`$؝0�S�'�+�<�Oκ����]~cպ��G|�ly��m���\_u������pXew�ņ�FNE+ʭ|�%�`���cX�S�1����Q�{���e&G1ՍA�q����^ݏ�2�s,�ҥ�;pȖ�ƪö�cYl,n4u�շ�7'���5�0t�,%%���ل���t��tv63t��=�zԬ��U�ko������t�J�^�\�h� �$���L�-���	e�vѶ��Z�L-3[�6�ڡ�*zY��~��&�BM��MC_��!�z'�N�t��r'�鮘G�e���74fi�C���,C��m����q��������E��s��c��<ń��P�c$��۲�=WP��B����$�g�{�N9��!��6vJK@���M�R	��=�ee��h��
� ���?	ȓ�2��e<�K>��M�$�Ųh�@
&C^l^#n5��6���pdĔ`dOBCP	��x�11�hO/�����O'��H	[!$��_G�Დ��*�gk���Ck�m3�����tm;��tm�[�(t��=�o����b�$�KO�t0�0�P`z g���'D�������m��S��hٱ'��'�l��|xzl�t�����X�1պ��G|�ly��6a�����gqf�z�*I��G�J�	� В�C 4%@�L;OԿ�\�̝׵���O�@uOD�l��C�P�1���IFz	4%x4�x=0?}��\�kG��(2F$�x `������):&��d��D@�z!��Kd/���#9H|z_�*��U-'�t\���0�?��B�.I��I�$,d(�$؈ z~C�?2f�.�WWj�������Vi�I��q�;�5��;ۈ�Q�5.�i�6lֲ���0�݇���	蜭�P�	a�96�ގ��?~{�9�3�<���{i�n[��ܚ�:��Cg|2 c ���ߗ$�T�q6&���x'D���akϚϫ�4T76��y➴�<���V�P�y���kYgq�>~cu�1�un��GQ�_:�)Km��|rz*{�~�(�2O��@=�����LC~�H���v�|���'��ܡ=tM�	���-��M���a4&��MP��$,
$���f���tIc2 ���M�60�d�I������2��d���,8XqvR`�3�]$k�)�m5��E���X��Uʦ᫽���5
pO�M���n���>��o�䞉Y(2Oz���Nz6O(�)D�~V�Cq!��y8 ��B��lL�n"0���z_D˃f���"�0)K	ȅ�T<-�Գp�g�ۢv��Ҍ����By=���ۢ~�$��M�R?Y)�&P�S�/�Pҏ�Y�_?��α�N����]i��Gξu�R��m6�n�\Y��1���ᣈPe ��	EA�'K�z!���>��'��;kcd��H�	����l�`|0
$8!��d<���@�ֻ����V&�Km�ʬ��Q��6l��\��p^�'��z4�H'Cb�LE�M�Ŧ������짉_i3�f\̧N��O�x|;�`�`2��2i�D�0�!?�<pIb�l �:h�'���:��=5l�d�/��
l�P5��c'"m!���n���$���i�3�p4C��%Ğ�Z���؆~�4h���R�C�B�6r�g<��؇ ����և��Ć���M��;��W�<ҟ�?-8��κ��#�1�#���ζƔ���޶�������<˙��!��ّ����=/�F��{��,F2�WO����̦K6���Y�ņ��YYG��̪A������X��wܾ�Ȟ��aEw��Љm\�����Ҷ`��u۷f���2�a��F�+D��p9Af�		+q �d�.�Ŧe�Mt�����#�KJ��.ϙ��i�ߌ��M����|�V���9ߵm��z�����X���UA�"��&�6m(�<�񘙆��N��%C���$������2t@�@�����o��UH�Ɖ\: �@� �.s��!�6�D7Ŧ	�&��n��GW	��l�AMD���܄�:���e��7 G���?tH�:2M��gt�0�M	:"&�N���E��M�td�<��Io��4J�Q	�A�dI�|�_]>R��JL��H��J����K�--��\�jI'~��jz[Hw�ض����vr��u)��I�`}���\�'��)N5���������#���1��1�#���ζƔ����X�9Y������ A���OC�n~,�Š�&����1!�J!�:3�>�"��Ab��?'�hd��l��O�q
��I�N�lѵ�C�fC\Zz$?#����mJ�����l(� ���l����;�蜣�۬ܐ��9�ӱ�(vCE���qF� �!(a�������	���N'2 FGN�ѥ���B�������W-�:��.���2�{���+Q�!�(Ȍ�9�2Қ4 ��O�RNt��<�6$9��֢a��H|R�D��N!Sq�Ɂ蓢� $=�VJ'�
�0@��S���8'�E�Zaؐ� tC�
c/������-�)�|+�#������#��1�Di�����_:�R���h����n71�w�E�~82j!ц��O�C��ڷ-��t�X�C�t&�Cڴ>��t��ð4�R�K�``�F	��'bz~)�"nC��0X�<)I����L�C�&�C�����?�?L��X��z�c7���B����7��C%l�j�H�!�
_aa407)񣆀Ao�@��XlN�j����D�j0�q?	8��)��h�����PN��=���4 �z0�a�L�"Dᩒk�?:�D����^2`h��I��>T�Է������D
0�C$�����RpNS�?#�G��G_��"1�<h�4�N�$B �'J:ItJɽ�A��T�}3zfd&�炊0���=	zs�Jg�w�1����KUZ��l��ha�L4zXQ:$�0>C�"l���O6��6 `$��#�O��-2<el-H�h~M܉<a���,���h�M	�)A'ų�0<�$:l���~�&\�j��0<=Qn�0��z&�Cc������N`$�hN���A�������;0�C��W#&��؁���&�N���N9�kR��vj��x hv�HLt`Y9O�!�4 Ob`ɀ�l�x'����fbSG��b��Ԟ�ac,��x"�N���I�8�d|x�pV[�~b�"���ű�b��c�[����צ��V-���/��#��zE�lk�|ƱX�����/��k�^ޱ�b��8���^�Ʊ������^)�^1xb��������"��5�u�������K�/���c��±��>z�Um������g��?���ڥ=>2�G�O���������ϗ�c�/⽪�5��/���+�/�z�^��b���]b��cV���3��x�{Vն>jؼV4�+JaX��ů�z���1x��z�Ÿ�Q�b���^���-L^)lF�[u~��1�Vظ�WlZ��1z[�c�1�E�WΦ���\E���~f���lk�c{��-��V��V+l|�+�[�b��~S����4�W[_�j~U?/o��׊�b�^��Ei�5��F/����~�~���[��)��k�\�����
Re{����әcn�#�Ox���;��挾��eWѺ�U���T�P�%ל.��GN^>=mUS���������Tܕi��R����vF-X'61�6aKI�c�z`�?��]����O���ŏf
Wʘ���8&H�����x�5��b�i�>�:��ی�v�+j5�x��DP��y�}՗|<���+eU+���o���	WT�st���a�a�g|�#�G[�5��g2�Ko.4E�ph�eǊ��LK=y<V7�s�:<�^f��nnm�P�`�x���V}����X-VV^7nf
��..)�ܰ�*<l��s�7%M�4Z�9�8�f�#��u>�nׯM�7SPn����p���IǮ
�/��uz��@l��-%�}��6-z�8��,��%#�1R;���&�����&D��{v=�*ǝ�;�ν�NX������q���P��$B�BϏ�]ښڦ������|E{8�{�Aؾ|�\�d���������{�H�"�q��`,,�ڒ�ۛ��\ض��L�^��+Ĩ����p[��jS]�F�Y-p�\o2� �`����ы��b]^i�o�zx�oDB3����Mfe�uL*�&,��i���e����%�h����)l�t$��k�.���P�[�ְ3EY�kv6�S�k��th�+ei�{��➳G��SR��Qꕇ^Óf�:�Z�641	M֚ռ&�*̚c��[O5�����2�D�g��Bbmm�1���vg��V����݋r�v]`�����̬�k�=�����=�~����~��s35&fd�������ff{���$̒wy�}����O���GGX�1���E����Җ��m���լ�����GKF���ΕA(��B�f�\�^f"f��XlZ�V�(Z6�0K�u��h늯�OX�e��O6�P�])��F���jMmv�%�\�P�b,2&�&����W�J���e�Y,�]}�]4�x���КqmD��%��U���d���ng����_�)�"��6��⍹oA{���62}�o�a�f�l������r��5d�[��Y���0���0a0DJ3ak߶&����� �p�x@ʂ��!�M����4Q�A��Q�O;����!����#D>��ZOp����-���ɱ>OA�D7V�ؚM�(0H�L����nnSfd���L�`�'��h"$���&�6vY8!����'���s8�K2�.,m�L��٘S355�f�����>A�4zz>�RXȉ�ta�4|~���,��6|Pɩ�D���h�-�yMy��y�UݭN��c���1���]b�|�liK[m6a�~���s�08'O��2hd�68�D4v@��N������-½��Cf�:��,&	��y&��DK߻�sAFyJ`����2�R���i0��!��o����{�6�"���C�AN���$�g&�-=�ѱ'Y)���!�lIA<$�G&C�0�I��/=���ֵ�^� X�3o\b��qd�	K�Z���	�@L,	Fg9��rL����! Z&QD�9;�4DVӧ��#,���?%̺?A�M�r$��q(lI��ٹN�'�,?L)#?"2@���\������*��1C�_�i��R)���~u���b#1���u�4��ن�6f�5�:v(�A&�<���Cލ�����0pϽ^Hzu(�f�&��~btOf4h�(PC�=��PF��k'�Z�f��>�|$� �;���D`��|t�Լ�뙚<l'@9ؿ_�q�ɒ�1&ӆ;�xܻ�OR������1aUU1J���:���\��K,�T|XzD�0`�wOp˘*Қ<Mw�G� � "!��L�)�Jh�_7`��Dʺ���|>:vOq}�gJn #��OFv0��뚊����@ ��A��Rdp�G �I�Da��<||i��1��q�u�u󭱥-m�Sf���5� o,����Cc&�No�*(�A&	��agOl���{^�~��qM+����<l�|X��0�)�p��3K�Hl߯��8"Dʀ�2�Eo�Pq6�$rE*g% ��y��Sþ��:�<�������`�099�.R�y6|~����� �6j`d,B��dU_���T�C�lgƊhO|���� �%�Ώ���R����1���O��N{C��2�i�O��C�!��A �������ڶN���FC6-<
SbSk��������θ��b#c�u󭱥-m����﫩U�]j�QҢ�����(��";%���{�meCyu�7��Lxq�D������6 ��> ����P��0��q"�Z���/�����5]�kn.�R�a��:%�ۯ-�n��.�J:DL�G��m����M�R�R:�~��BY���U����)$��
X"�D�SV���yx>�9l�f`!���5;3ɣ{�ꥻ��s&��k�s6���6PA�)˱�����~<&�_��&�W���qWuV��-��sJ�F����'�{�}V�whtk�;��4��������w�Y�C��Sg�>0( ���[j�O�ne�!�Ƙvq`fb�Z�ֵ4I��~��J_������ g��>��Oy����u����O���>[���G�\q��b#c�:���Җ��[o��(�z�mjT1
HbE<��)A)�FS�O6pC�3���f\�i���;���ڨ��xy<��(!���NjyO�4h���ж�P�G��#OU攩���𪀢���a��#��eiu�O@�q��m2~���(������w�:X]R���Ҋ���ɘ�t�7��b�|i�I`�
�I�.�J�`|4�� �D����?t6t� �@�9�mqZ���wwJ-�]�\m֖�ۯ�cq�"1��q�F0��[cJZ�6Sg��ގo�!�?mt�=��ѩ!aZ�*��5|�HK!�Ć�90�?}�mf�`�wU��l��C���!$�# ��($WW.��<�gN��ώ�9�6��6!$iL]A�lv�42K����ִ"�n�N>!4	����>_]�'�܅Q��/���JC�d�D�]W㵿OC`��Y�����`���x�g�!�*���p0цL]�7=�>��Ea�}f��C��񅐪0�DY^>���=u���c�:���Dc�b1�_:�Z��km<��[��O�X(�A�Mm�)S�>�MS#���I��q�����Aw�T�o�Uf}3,�.ֵEk�ԸU��]f��	��i�@����`$���!�����*1�Ĺ�LF�d!+<s�{i:��a�C'�~��YF�k;=�y8$%�=ϳ��勨(k�Z��L����
y�@�k��͟�?N���<��0��ci��}$���>'��1!#x�V-,��G�������b#�F1�#F�mZ��km�-�7�����Z�m�Oo�_cC3T���]�l�Td7*(��Y$G�Y4˚K���y��J��0^�D؉���ۛl�	�`]t������0�1��ѻ�6��+Pv؛�,V�l���1[���e���L�B��1@�pHJ��ҝ�.0��l��4�hZ��[*Z�m5��qH��*�Q3QT�a�������h�.�rt?}�%Ktmxs	A���Zto�H�_8t$Y�=h��.'ʁ��ƴ��l�'ц��͇��
z0�;�5i�x�G�������p�g�F~����O�('���I&��<���K�i����ߍ�=���D�O����<��Ёa� ���3۬�x��0r��p�a*ܳ:Nl�Xϐ����DD�6z4$���xR�(�K�xϛ]��8�<E>~z�8��u�1�X�:�c�6�-km���''�n��j�۪8�QH�jS����3���%ߜ<��1���p��`�z0@�1�O3a.�X��ާ%R��jڞ"z7;�a�a��à��@���tQ^؄C0$���ύ4Q�w
p(',��������Y��e�0�������հ+l��b[���=��%���3�$��:%�#�S�bS�g��K
xl0��(�J3���s��G	�u!���MѴ�ٱ"�>�.LЩ�ԧ�<�p��zk��֘�?/�����i��^1lb��ⱎ5��b�V�[^1x�l{��u�k�Zi�.��X�㭱�b�.*8�\u�cK���/�qx�ⱋ���ck�X���/�V+u�k���U�J���F��[^1x���cwX�|^cXŽW�b����==/�螏���ھ�F��EV�uk�q��c��x�E⸬{u��b�?/���1���/���1~�_�W��/�b��ⱋƘ�4ŵ����x�vű�Ҵ�+
b�ǭcK�b�im1x�5�-�x�,��=X���c裡�Gҗ�0�q�[_U�.�|b�X�q�j�x�S�ǭc�^1|W�W֑���TW�~G���L�c�/�F��^+�X�|��|b��)�DWU���^�n��~iv��S����_����Uz�E�]i|b�X�A��Ax�#�	��j.MC���fE� �H��u��)�~�/�F-���ϧ~zۣ���7�lQ���M�3�:^FZ�G�j`]zAl�P��1cb��3�v'�1��`�rg_�l����5߅���G~r|+d�SXw%�F��1 -O�sY���%�+�*Tc|�U�"fX᢯�Y+y��'��J��/��~th�{����6ߛn����=�O��:m��n}��~�{5��=�N�Y�}��_)�z�����":�1���6���ֳf�l;�E"	���9�6�����iGgC`����o�j8۰.��A>�D�0��>c�k���L52�d$#�Qc��g7E�ı2à���i�dh@�,V���8ШĮ��ȗ�ѱ�4�ϒ�|��90�8	��C�xt�b���O����O�2RH~N���т}E�9=6'��R���e�"l�~��5&���6�4"&d���?|p�:Mwm���|��P0>_4�l|��m�~b#�cF1�#FѷZZ��km���ֵ1���pQA�����w�2R�iCZ�~3��o���a���w�p��0DG���e�|��UR|�,@�̲$K��c1�I��3*S���0�`p�٩�""@=J0�� �#	�$�FS�OG�Ј�K(h2v��pDDD���n��æ�tDOi��l2��afť/��؈��~a��vl��"vl��舉����������v;K�T=�B��K�,f+���o�̧�x�|�X��#�cc�u�Dc�q��lX�şu}��L�q�
UKo
�"��L�`N$fv)������-�{�!Uհ��X]���<LQ�DD���T�i�-��i�l��x�	}�3{]Ak�y��ޗW���D�hj$�Xޥ�bٮ-��`�SP�-�v2�b��v�� 1�s^�\# -$�o~@�!B�Xc8���֔�6�1�dUm�TTr�/mHN�ܫV.�����qL��Ҙ"&�l�������Z�WV���((B����JϏ�Q��A�@�!,Iw��g��Ac/�:!G�Q�����AԒ<Qޝ�}4{�Z]�a�Ј��#��詉o���r���ςh��}0b�f�6����|�>>,Xa����B_Ͽ~U��el��8�,�Mm�\#���i,!�)o���jY�7�٠d�,>��V��-�=|���:��#��c�Du���m�KZ�mm�u��w�TA��O8��g�`��N}���p�%!��ORf�΂tE�o$�v���X��?��ANO*_>a�qpe_(���j"����S:��O�QSb j~���^�8�PC�uN'ɅҦ�����k�qi��B�&4cVa�2�3�B|+�G�-���a�ϯ�4 �y���X9�tfپC�@�k���ÓݛT�W���S������Wv�9�+ƓN�-Dc�":�1��":�c�6���f͔��V{�6��M�vf�ࢂ7��Q�bVsƖ^A�jT�bR��$@�4L������y<�=��w��H��]L4:�DܟH/��4��є E�A4a�Ӣ����"bbZ��@�MW]/]��h��%g���|�����B"X0����g�~����^����wϚu������d���a�w�|��)�506J�ߚ~Ex�1"��:�F�y~{�W��K�nS�d���Z{ӧ➟c�~c��#�cF���6l��ء��Fe���(��@�%�ϥTL�p��0e�/�Iػ���8a�H�g�$�����eI���T�#�e��>c4�?y�R���������?x}�`��J��������B��"��G{�!�H����^]���>c1��_���)���ѣ�MϏ�y�Է2n���b"�ؔ��#M((�Hv����N�ҍ�����f���+v|���SM?-�_���c�:���1�mm��m���Չ{��Y��?ҋ,ġ,\�4��=�1�\CX��{��b�)D�@	�I����,�ԍe�Bn� �ZZ�
� �F-�^יJ'�KN�X6V���MY}g��k��f����ű��ìɩw ��V�Ԭ]VUٕ-1f���۱��p�39H� HBMd����3u2��uc�	rb�,3���k*���2����?0�ل�,�|p5�m�OsO�|�� �CI'����:P�������4t�]�)�Q��>#����,P�,�ԢJ���IA�)��M���|0��;V����&x�,��r�
(A������)*������)�?"=�(���teP�-ol���,KN�뎰�Y�\�������F�(�+�\}��"P�L�􍥃;A�������G_��1��#FѶ�Z��km�W�;EڮԢ53&�PD>���3�Sӆ���'A0�f�a᳂ tJs��t�DC��l<ѓ�p�����Kt�N��H�zy4" Ξ�������N��X~0٩��1�ܿCȧ��`{�m�<>6rdN͈�3�p^�|k-`��Q�iR�.���T���R��� ���{䷌ҍ=���B"ΐIe}�I$B#Sc4R�'��`�M�j�W���Y�E��4���>�:A'H~|��b#�c��GQ�F�ik[m���#O.����I��?ti��ò�5-�{�6�R"�
���9�R�=�5�σg��f��>�o��ˆ�&��(�v���=>,6gJ!��?�P�,���)�X7J�A·9�Z`���PV��}|-�a�^�ҏq ͓IB�y��>*��t����va�����<(yh��Q�D�*����f�b��2;���6!�Ό蟊,O�7yH�������2���|t�"5oX�_��Du�b1�b:���6�KZ�mm�U��.���e�fY�������ޟ%��8p��4!�BaÅ�S��8`���@�m
�Q��+$�-B��g�Bm-�ű^����er��e��aes�D�����0�9���%L�L�)v����0M&@�z�h���C��3��Tx�φtC��Q��Z��Y��\O��h�a��\6t�N|}��q�zpC`�f'�����4!�æ��H=�q(��R�E �Q`�9��?%�
BK4�9��݌��N�u�""�DE�#���">G��ڐ���=DqƟ"�h��6�Q�]u�8����""6�����Ǩ�"""""#H�#��#�_)�]q�DDz����H��F��m�8㨎6���!�DD|�Du#H�����DE�M-�����=B8�����V��kDR8�T�S�1�0Ӧ1LZ:�\i�"6�hB6���c�8��뮱�1�1�""#����"#�m�8���8�[��)��>c��ǆ`��iC$GF�t)���"d���R�Vr�"r�K�fj2ͪW�����!]��Ҋ��1���C��u�Sql���ŃL	b9x�gd�|�-�u�l�O�M�D���nL��2��Lƈ�	��c1�u�-����Ų<�x�{3ޏ�H����� ^8�Ck�Ym��W��d�f�6�	�%�B��V���"��;rL���k`���fH��}��! �v��qֻJ���}��W����)�o��n�Ed+4b�(�j����ω~:zy�"�̱�Ou�&�{.�R�k[�8$��b�Nc�y�Q��N��z����f!�5�'��{�0�yC�w6��\z����a��&�aWE:����]6G�E�!EA��q܊�8��r
h�Vs�GN�R�Z�4�1��F��Q�m��l�fV�s����k5�a��Zj�����el�g���8��U��l�T���2����i��~̍>3=Q��]��n�m��ko^g���ƨ�y)fU�mY��Kxw�d�q�xV�+��,F8�#�j�6\�+���Ȏ��1�!�U����i`�f2˞а��ɥ�6�:ۭ-ua)hn6ˮ�]�@�W���BR��$v�m�.�b���NB�[E��eҳS�݀#���mafQ�С6N/%�Q:�V���B�B�]n�#q���l�3@!J��{��cn-�.����][;\@^lGZ3fl᱘(������5Фm̶m--�.LU�{��D�(�EQ�*V��RBWѧ.a�+c1�gBj4��p�昗B�XvM�qm��z��$�+|�ʢŕ�nT.7o�)��d$�*��������Y}y8������>ww~�{��m���mϝ�߽��6�}m������l����u�1��1��"1Lmm��m����U�\`=~�Jm��vy�(�#������IR�5�����Č/�ԁf}F��&�%�ѥ�!���(jȗ4��cCcM*\�͓bݣ��Z�R �9�׳L�\�����݂Ɯ�1AZu�i �y7�$+&��|I�lM]	��n�
�X�Y�"k����ϩ��Q�~��<Y�^!#�,��	H�yY,���n�**��(�x����|+��g<YӠ���mr鉙�4T{�)��_)�M��X�
p��nro��$LI>���5��ǉ9��X"�?{2��}��~&�*��;2������=���������)��SC���a�M����f��wͱۚ��6��a_ڴ�2�V-N��0w�TAR)�)H:_=��c�I��I���4ῴ���ua�������b:�1�1Dc�6م)M�)�a�oS�j���EC�0��,���Jl�D���H�RUx�g4���������gD ��=߃n̞�a�zto&��7mTZh�Ybn�$��Z,t>O B�,0t��eQ7�rp��J!�>@�B���wB>00D4l�:�Vk5JmP��1��Ѥee�WJT-��^���>77.���h�ᩢ�!�&��^��{����W10\��>���DC�z|���|�j�U|q�Z�~Z��4���1�X�b#�1�F1��m��)�e6g���|��\U�������C���D�.a������8"G�:Sg�kS�0frhMh>rI�����׌�L���>����cg4y��(�}�֯�J�X�V7D�L\A��׭s��R���mCǨ��~w�Ƨ�9'~�56lI�ϧ!�ň�!i��t�7�d�w"'5&t�P�A��!�x������ݔD�2o����Ld����X�oi��S���@|��
>QG�`�>0����Q�F1�c��cF�ikY�e6>��,P*,����O6�(��P�����rK���?Js�#~56g����C����,-�����Y=��l���]0]jZj��8v!QD��.ż�ƹ��)��
,�P���=NV�ٳ�K5O�Ӑ��gK��Ѹ^�O����,6'��S:�S�Te�cD�=8`�==�-�<:rJy�o��{I�9�����e���0DC�K3��Г۰���ฎrH(d��Ϗ�4���Dc�:��1�m������-�Э���X�ۏVK��4)k1̃U\w+�phP�k�f�R�ˠ����ǜ�z;P���̅�P����L9)�x���Q�a�DB�e	3qfzsr�jt'*DmeQ4��fecCvl�U�@�����;!]�lڬ�3Bˠ�����y�$�U�(ج�V]nU��6��cU-.16���^�!�Fa��F~�
$0���;�{󚪬>��r���}FB��߇[sf�8QD:��p��ӡ�z���âF
!��6aMH}��ݔ�sĶ�+m�k��
pD$DI<'�" ��J+�tRUUT���F��r�,�i������	���C^���_��1.��bX�)rka4z	�h�ęa3M�`��MÆ��6l>}���w[eRIl��[S8���	I| թ}
g�1�Y�&|3�N����1�u�ch�m-jl�M�����5�EC��5u	A�H��Bj:I���TD��u���C���V�Ї�)�,;=���[j����S�=���w4|X��F+��ċ0��!=��(͍�ʈ�"H�pD2��<�1?}d����4��׊�-�ɬrF��+�TXF�ηSr�B����Uٹ�(���\>��>>:`�;����/�G�g���;�S�p��lC������	������n�4�b:��Dc�:��1�m������s�z�?�2�I�IX)��(#"$��iK�"& ���=�0�=-(SI1%g�Q�A�e�x���cb�Q�>�_�GO1��(A�S���*�g�4-�Js��J�M�f�B[H���|��tf��x��(�&�%)����V����l�dp��b�	����?�3�3��i�q��g�2xh�������A�O�I/��5CA�
�2h�� �������1���c�1��1�mm��m�������JAٳ����~�zS��WF���U���!/�U���Ӧ�!.m�i�2�T�_4�F`��.���#~�?�F������Ģ �&�v�M���{��ܞ3�Ҟ�}&._<h��Q��(v�[Ĵ̶���p���{nM���'��Ι<=x��)k��g��ԥ����Q�,,ߣ�;⡎&3��$���,tO}ݷs�����DG���"1��"#�Ѷ�Z��km�<��w��D��;����Vĭ�+�]7�yJE`���Қ^��5���r�ɗknM؅
�|l�(���oj�zτ�ƥ���q��(� y�w;��ޔ��x���]���(*�m��XCMq�
�[mB�Gf�Rk�:i��B��՚<����$!)�=�Kl��ϱ��Y�jbWR:���:笉s���R��2�����s��� }$=�ʘ��s�g�%@��I����[��៌TM�aD2��h�U�I1�*��3E�Qa�SE���K����8"�Ou�fe�w���e��O��F;J��F�z��=R���#����<P�
!�╦T��u�I����v��\������X��KI�������:���DƱ��7��8��LF8㮣�F1�Dc�6�KZ�mm�x���T���8$�1F'b���4ѴXV�!1Ă�Tc��9�EA7�ɗ:3�?~_�D4 �Mw�J��c�]�O
a�y�nhN?��B��h�a�5���<8$�.>�8h?!�%.�=�_C1�'��'�GN��nh�|h��`"�����qѐ V�������&6I��D���_OϾ����t����OӦ�n|S��[�.am�<2lDD0J|d��}�;��١�J=�V�������ӧ�<{��ۍ�������#M�DF�DGȈ�#h�T����F�G�)�Di�q��)��"=DDDGȈӈ�DDDDDDF��:�#h���=DDuDDz�GQ��D>Du�Qm)B"��-DR#���)�""Ѧ���������#m������J!H�=ih����Hc�b��mLb�Ƒ��Du��P�z��Q�"#�:�=G]u�m�1lDi��"#�m�#���8�[��jB#��m�1��c����|O�ߴ��7��w���TP_kk��
2t�?I��"��c`�����c]�H�����;+�WH����~cg۟7ޣ�Xi����TL���2�Ap(�M��|Þ־�m�x��6JR�c)������؁�0�6�EOv�}���z��|t����~�ag7�Q6�c�Tdc��V�Fԃ^ߺ�7eO
���6���4��LB�E�60��]�~sʦ���~w�_Z5�z/�����9^�պ����wWB�ݸ��۶�~n=�w~�{��m�ow�Ƕ����zm�m�����J,�c���F1��b1���ch�֖����^kj�QJ6l ���?�w�A8P,��g���u���h؈��=��6o���Ե�,ٟ.��N�!�8na��^<:k�r��6pC�L���[��г����[*mq��Ŝ<z���w{zܵ]���qn�i�D`�/��o��\��F�g�4�s��	�T�OxQўB�+���{����0b}4*�C��\<6����6~6i���?:�1��b1���cg�f�)Jl�M���rI4���,HH�L�3�sW�g<i���SC�Jt��m�����ҝ����sƊ9P�rZ�������A#-�����c3u�+�Jc�F�Nk>0j{/c��`u��==>8~�i���������msG����F	,����6y�R2J~��o�/�:o��B2xt����
 ��i4�MW�TY�Po{>�94"	���ׯ��g�Q��x~�A���پhSfΔ�a��i�X�b#��:�1��=6~6h�͔��e�M�nf5�!��\A�����D��l(2�Gc��cP�8�Jm��e�V��d�M�At��`Тq-Ɩ�v���S�)i3��H\)u-�º��6h�hc��BҎv��]��Z�f}�e�Yd�=�\Y��a\킌z���k�.�f�b�S��zzp��|Ƙ �hp߿]���k��;N�<4
:6u>2zaOD�!ӑ��՞}f8��>�<ᣜ��	�!��Oc�Fˣg�_���.e�{��t�%�@�i"
ޝ=Ȉ�ĩ��.O$�>0e�{�ޛs�g���xhЈw��>L~�w�K��+z�e[]+b%]Riu&��UT��f�24�!#���%��,�p�͜8}ގ�s1��ǟ�������zۯ�8���Dcc�F1�m�KZ�mm��z��b&�ࢂ!ɿ5mП�Ɇ=2`����}���Ge���ϋ�bOz�����>&�ګ�B!O�JI�ϊ(����@�sD4�tf�ڞ�Q�K���t'��ç�4%'�U؉*%MDԨ���V0P��0��k��s�����2SB	�K����-�zl�v��D��L:R�)G����AF��t�,_.�{U��<u�Q���������X�1��#�ޭk[m��}k[�V��E�ZoҘ�"�[�r�QA݇N2l�׆56o8'��)EWӇN�x'�3F��0�4�A��V��������<=<;D3kD�цK�C���˕׻����y̩RL�%��=�F*!(��\�T̑1�o$���c�,:�j�%��E�*��k��9"?r*7��x0���&��Κ+�$�a�J2!����q3��b�#���׻-���S�����ݯ�ɔ�X1Ht�΋��w��-��YƘ���Gq�GX��:�1�F16�kZ�m���hUǽ(��z'L;<��W���b=����!P YL)J>{�.f�O���-B��	{�iz6�m��Z�ZnL/��z3�n��w���)��5)��J�p�7���h�Cg�Q����Ò���Y��NM�f	�a�EW��B�O�W'��b��rF�	�C=�śD4+䬣�WݚAR[�У���agO��2�i��:|k�?1b#��1�|�զ�k,Q?��#����K*�o���=�z�K��&���f��A0�-�6��7��`5)<RZz�Z�#�P�9K`+C����hG�.��.�A�U��Ц��Ju"�T"k�L[fM��-�kr���Ax(��f�n�N�-�q�p�H�$*(�M�z7���>�[N���i��KQjZ���7���k�8"���7f����-���|������� ��$����A��2�hm3��6�Z]y�DA$��n��͉���ϴ͆�;6'L<�зC��sƥ��a��t0C��d	����d�����5�V�J<Q�PU�����b1��H�G�������I">#N2�Ha�mDLLz��I&C4��1b#��1�|�խk6lه:���EA���� QD�(��+�B�d�*#��V�a�9J>�%�p�"�AÞ ���M�������<�>���N������E�I͚���s��a�&��(��~0D�D��}���a��q{�	�K6�.	6e��8������އ'4x|��Ȟ���TMp�ڮ9��ݏ����HH��$�K2&i�O�C4N�><5ĵ�6l���|l��6�����q��c�c�c�E)Jlٳv�Mɘg������/�O�ꪾM"R���M �3��y��3�㊱�D| ��&�L�	*��Gy���v�%�+u�-+���s��RS5����<>x��|?bQ@Ϛ&�x�4H�0(ߐ�B��'�h��H���V�K�/jD�SOL:o+f�i���}>�|�S��1��~u����X�1��#�ޭk[m��s�J�����=���J�cP3,���x(�JR̙���[�d<:}���xH@��4�a~V�|�b���v&�g?�q�mh=����Ͳ��,��:�����j���?Ξ������G e!*,�X�IfqXrL߭(Ԥ�����$��9�2c�ǎ':MY~��W�����Ȃ`�#�L(�9џiB�	|o$���맘aV��\Z����(8u�ˋ�xC�,&�|t����篑�"#��4���"8����4����"#嶈�G��ӏ�#�8�"-O�G��#�������R""""""#�먍�>G^���6���H�ڛD|�뎣���qM��E""#�DF�DE�h����F��)DDDDDi��z��#KZ<�E8����"-�=R")b>c�4��ژ��#�>B�DF�"6�]u�G]c��1����)�i#�Ȏ���qh���"ԄE6����F1֘c�#|�ʧw�.6R+k �q�yl�[�jcņ#�"��+�.��ֲ���Ż�d���e5ݎ�=��H��W'm�fR��q�c�=��R��]�U��3�n��O'1V)��ל�lD��D;��x'���s೻�x�&r��R�̓5�b�O�)��cEF��}N�����̂pM6�W&{W����U߉}]twL�b��م�nE���4!�:��8Hf�NJ@t��Z�j��n9�T]m�~����#�9�������!�F��MSX�rŹbY0n���n
ٓ7ҪD�,x��֎wjF��\�.�mm���E���꙲��c�ە���\<��Wj�������w��
����1�2b��;�.�Ǘ0ג��&��n`�=���Na2
��Nw�k��nc��ÞN+޹*krHfa�غ;z}��ϵ�����=����7&(0M�ؤ�Ӓ�=xU���wnl�TdUJ���(5�i0N����h�;�=dP�S�p����(��2vN�뫫��妬|����;���uU��L��s�m�]�w��߷|���ʯ��ot�����cS�
ʲr̡6ʞ��k�<�p�#}4�[nvoU׫��ʾ��уkTj���Z�-���d�\�51V�A��Wj\�j �I]#r��*((1��f+�l��v6��R�.��.���K�cam�Ie�]�eSD��b-߱�e/�鬌�F�+���6��fku�J�bU��ݶ�\��ȸ9�Ĭ,�U!@�&͵�������d�m�%\4�J�\u,,�ٸɖ��g���n,1�� %=kf������C]	��0�VK<,՘�ey۫�.�V�j��&k�vp)X��Q�46KK�CC��ct�&����!�4�%I3�'��X�[m�{����{�{�~^���x�wǯ���o�m��=����{�<c�n��b8�F1�1�b?/��M4�X�b����	,d�݈-��f�k�1���hZh+
�Қ�4qQ*�5uem�9�pLBR���bkm,b��#��d�%yWT{B�wh�MTM�Ev�����k���S\%%�fE�%tdv&�(��p@���X\�˭��t�Z�,��"MIx�e���eW���U����}ƽϥ?��-�~,,�O�]�z�ڵ�ɺY�"���}��r�i�9J��x�9�nBU3�	��U|3CL�����l8nhÚȉ���r��J���f6�f�I7�tI�>��V�s.)��>�����Z]�
���^���{�kLd���^7*��%W5ŗ9��^n�a��ZWJ]R����Ql��:_HtB�e�.��>�_r!D"&G�c�Ru�m�q�1b#��1�|�խkm��J�/��M&�r��f.0�b�^b(�N���ԓ��<=���O=������ᐁ�B��GIN
8}~;i���OU('|s��FO!�h�=�@cUr�ҪJ:y�rx$���:i�sޝJ&NP#v�TT��$���q��V�eB� ;�#��M҅�I��@Y�'�3ԏI�G�����e���'O�=6>��`ih�8h�6||���q�1b#��1�,�DAN�$�[欢J����X&�'���S��#�'툇L�'�%+�ȕq���d�b�y��Y�ߠ�/�C�W,�����O �5����!H`�&X�]��QDID��X�z2���(\�"!Oɂ~���>: W�Y��Pa�B�,��P��*'Ǉ���g�=����͜��b8�H	Q�҈߄��Rt3L>~m��F#��#��1�b6h�)M�6d�e�J��]��D*�іIQr�������K0DɜF2�B�)'��	,AE��������m�\��5�����m�bY�(�|G/��*�74Xxn	���r�-�xx�8a�x��Se��k���٣_x+�m���̣��C����ǡz��.cWá��K8ç��'L�.	MW�k\�=������S��%<8τ#�F:�(�یS�ͺ뭢8��:�cc�c��z��m�X��˼<j�ՠ�*���RG�L�1J�d��^FB�2cC�?���
[�d}aMsn�M4.s�X�n4Y ��m�iɖ��ٙ�ι�,W�U����d�M��7=��v/d��tH���I�PB����3o<#���3
�]?_v[-�a������i����������l���&1c5eDq��Y��q¦����p���C	�﫚��u̙��<��ն�P���óF5(���N���20����_~��J|z~7<I�̽��G�hW�MK8)����S^X9��KL��u[���{<�=Ki��l��6la��&�o�͍f��M�k���v�̈ �9)�th�s\�~�D�> s�~��*����gy�J�$�������g�1�F1�#�ޭk[m���U�n�
����E������Hh�N�gC�ĹT�;0�a��
�)4w䙥��T!"9f'I��l�E�F��w��6'��m)h�Kݒ��y�zp��g��ϔBB۬��pm1Em/*�bf����fj���9�:�K�)OӳFhG��&Ք({a�h�eM��R�y����М��á��ܶ}��-�������[�#lc�q�6�����#�����)M�l�OHz>3Z�HMwJ�!N�:M?�=�'�>���Z��i}���?;�V���Q���:��^aO'������4~8~���)�
2y-W�%�w��Ѫ�mD�cQ�T][�܁V���l��lŝ
�zxl�J'�5�ckKXl؛)O�"�) z!P#ө�類�SВu 4mO�S(f�|a%�]0E4�z���==�艚�8�j*���П<@�	:R��y���*��M�1#�1G]Dq�c�|�|�խm�ٲ�i!1"�Af2H�ڪ	δ�'��>S"�"jc܃�@���i ��݄�#g��D��)�BGBUl���"*�˼*�o��:r��kX�)��{��у/�A���Ai|Q���A�4���۞�<;>6k4[�у$/u%�=^�D������QTm�p��L��$U$��ǈ8�ޥ�;��H��Y㥘x�L0cmu�1�F1�F޴����,Q~c=����6&�t�_Ԗi�/�5��ɳ�Uʆ��@Bn�0o5�����.�oNEZj�;��Yr���*�j�Ֆ
ZHw$�k���%,������n��^�Ʉ^��\�D����)�
髤*b�9F$6�\����{UPK�7iW6���1��[ax�6֗Z٫�2P�R��:ܶ��Mg3�����?>t��XoU+��#�LΈ�Æ�Jhfq�܄:�
E$�?��~?N�e(ǯ�~\����5'�p�PفA0<������+�L�殦����<O��,���������̵�D7�btD8y�b�������M_��}]��eV��m�1�,h�Y[��(���S�~�4G�F�@Q!DR$w�#�ǥ]�zyV�'�Y'O�0e�`�t�����#���oZZ�i�l�|GXL�1�ј"6���&�8d���A?o�=�5��n���A�%1$|����I�.L��:"��-�Ƃ��u]���9����1�g�g���o�3��8��l�~9��c�!���]���J�Amƫ	�4muˣs1��&�6�(�6iF'ǟ-��zm9��b�g��iTq-4���)��!�~0$��B,���zGg��<��Vەe?@�m�<R�y���|��X�8��DG�DF��Diգ�#H���u)�"�Ï�>GZ""">D|�QH��DG���D"""""""#�DF�u��"6��DE�=m�G]q��E"�B���������DD|��F޴��DDDDDz���oP��Z���-�=z�DCN=R""�p���1�m�b:��H␍""#�G�u�]m�u�i�S�D|��"#H�#���|����||�-HDSh�Q��E:c0����8��ɘ�����i���OUBi>�[�)�ZD�N>s��6�ݝE떵86l���n�X�m��/2z�ł��l�u�]�~Zߤ7��:�y�7&o�M��Sq���ץ�z�ƚm{�O�e�W}�>�γ�x�s{{�,�6�(a�Q(:E'TW��0�c�>A�ܔT8�~�.ٺ�g����m�6���S���L�m��w|z������ܒI�������̉$�NN��Ϸ��cq�q��u�c�clmz���M����ꪪ�w�m�m�<�h3G�����->�t:�Ý�vDO
=���j;O8���,�-"�H��ZhW:���⥟%ݮ��B\J�i�] ���pd�yDv�LӺȈE[����4�Hv\P�q�]$�E��w�jrD��z�q�&:r����G$�8f�g���Zd��D�J1+ذR,��P��Q�>;ϐ3��uq�b=G]Dq�#�?4aJl�bt�u���_3%O]!%n�����k�
��|x>=%<��o��6���J�ƹTlN��~��:��Wi���@�K*4n�ƈ�!�p��5>�ۜ�"�$/ˉ�U6E�*0�K�ϑ�V�B&�	ٳ񣆃aL��	��Q��>Ac�%dQV�њ϶�8}�S�A���anv��|�i�L��\9�`���^ZxߊZ����Y�=F=G�Gq��=G]Dq��cch�ф'�=,���}}���
�4��m+�1-c��Zᦪ���J��R���=�[���!(sf�e�A�UV'"�X�RR&��[����\��za.�u5��sR����M���8҈�ԧ�um� $-���c�98�)A���2Z1GD�mV���*������s�A��iVK�&�=0�Қn��	^�YmZ�/�]�[X��S��dǣ<���ݖa�Ç�2zw���%y]�U�%�(0�b��逍��f;��+�.[m�'Og��~�<+�E�+���>Z
*�J(=X��1a�Riz˶m���!C�D*��Zy�=����֣O|٥�[�=o���*fV���Y�<i�a�e#��8��#���oZZ�i�<!��_�SQd�5�PK;$�v{�͙�_KJ�6^�av{�UԪź�?4��4�i��o�}U=�1\8;g�O�����pᾌQ :|�}�֑�3�/�Ed�L�43�Pc0�q���K,�.�[�j��^ذ�D(�g�z�K$�)#�Q��H��r�d���cq��O
h��3d��Ļ��]�K���F&(v��^��lm�|���q�#�u�G�c��m�K[m6�[mڡ�WR�j�	��'�
��gJ���nftq?~[R�Qbp)Æ��3����V�5��xy��xt(����G�P����
>)^���>O�&�Z��� ���É|�N��0����tu�1��gߋ8�b�YFKN�m��TU'�6=�צkW_M2ĳ�Ƌ��a�4R��e��O��L���hv�N�����d��p��D�ᣇ�8��z����"1Ƙ��٣
Sf'��S�/*�;�����m�2�
	�b��G�!>O���~V��-w�NM6R�٦�c�4�" [�>�A
#�7�.d�_4>e���֫���iX�<�'�����oTy爯�X��=,��<����4�m��a�O��f��O����+������x`��^劍�.|�ğ馘a�e�F31�Ƙ�6�����Su�֕�޷G_R��O���Oa�i����]��%f3(��e
W� �&Zˁփ6F��$�Z��B�����ib�^o�������F�XLd��[Yua�vƶ�큹��m�;e�j���;g]|���/y�>*ى���X���*X�u]��H噖��k(V�9g��)��y\,b0$�Ya�D<�[��e!Z2���G
hgߟ�̮n���N�����f͟;���a�r� �9����b^���4���C�-$����$�}���d��^�5l�R�B*�!� ݮT�r(��uj�ή�ۦDg�ब٣�Ow�w�Ř�U�A|��D`�s���q����8��F1�6��aJl�g鹏�C�]\�v���/����0��*�D������(�nfL*�af�oa�y�V����q�1L�0�s��ѽ��0f 頸|uxٙJp��8A��&�HR�J���7Y�1�u�cf��G]����u�	m�t�zh����S'���߫����ǝE�B���:��*��#oJ}J����~�--w����b�O%<m�:�8����u�G�<x�Ft�H �'N��ک�TMU��Yi$��D@�AL���xB��o�=:&Ǔ�F:70���ӻ�5:�(,$}~̸g�J3�Oc��cg��߯OXxey�S[�}My�n�L�.��k����k�����ً��kn:�N����RM����FQ
\%	��O�O��g�~)�春j�3��Ϛt��o��P���CI����oe>Q��u�~�0�� �y(��s�-=�>$ �
�:��b4����":��b�?0ن��b�lĨ����H8U�9�Tr�<������vn�"R�N��~UJ�g��r��L�R��M�Si����#-#����ci�:xp��Lf���'}�G�0�n�Y��
1��:h;M���&پ�y&�z|�=��Mf�k�ҺV�x�FpV]���ђ}0���ю7�+o��]���8h~^���	�u�M�Ʀ�M���mUi����{<;�h&Jw�n�C�'��h���X�~i�F)�DDB8��DGDiR>iDGȈ��M"-8������"��Z���Du�GQ��DG���8DDB"8��DZ#�|�":��Gm�!�-8��Q��"#M4�>DF��"#h����6�m")��DE�M�"#OV�>DE����Ӭ|�c�8�8�#H���z�]u�]|�1�c�1����Di�>GD:�:�Ţ�>SHҐ��|�QGȊDG��u(�?/r�r��c���*�U�|��c]썪���K���&{#̘����S.6A�p)dw1ܖMs5�9s�eOm��ǫ��E��f6������s���|"NX��9K̈#��p^ن���Ű��}}-r(+qI�ۻ�bd�d���\��	kW<�r��6���O���H0D̲;`[r�gل�?u��v]��k���tx��Mշ��l�&�ҽ�7b��M��U�X9x�d<�T�-!����m��s����{��ó�	n9re��]��䃁���1����cg���_�G��z�P�/Vǯ3�-�𞴦�*3k���ka,�4z@��ڊ�rkPg�_�S�o]\m��E1�<aۚ����)�W*�RfzÐ୘�-�g�\��<f떷��=ط.4V�E;خ����ՀH��*̌u��E�b�+(����2��Ӧ~�F�>h�8Kqݗ3�<n��&�� 3�;��;s闻�_�����.�y�����y���\�{n�g��
%��q������;�"��zt-O_��{61������2[�L�9�8G[��-&��F�h�.F1s��9���ـ��P��;X���n�]����+�b CJm%�Xe��Fm�J�ճCe
mh,��Զ7!�t�ֈ�v��ƳK6�SJ��Л])�M3s��̭L�g&�j2�lc5#�1\`/�oye�������Ky�uuf��!�qe��u��a�aLm��me�f9�3�ckd�D�}F])4i��X҄7�6Ի�/Z1�z����m�cq�@o+!"��{����m���Ǖ�����xm��{����{���3��I;��2�������"8���#��8���Ŷ����X�����1b+��kT�'�5-��
��/k.%[�e��ĺ���"72�[4���l͕�j����.��͚��YkfV�ZU�:�m�pp��鐽[eW4���2%��mT���Y�R�Q��%[s5���uڎ�q�	;b�ȉ�G-�� �=,�1�r�q�;8�Z��_K���d�cf�櫗l�N��?�}?"�N΅<�S�ف�^�U5SU1'�f%�������`[�`�sÂ�:6���6��^�����)�ξ-�O7�L���6H<o4���]�Zx�Q@�c�؍���m��X����6$���=�4\pg����<U�(�˶�n���=�E�@�[Kev��i ����.P�(��=�d�x��>|㈍#��8���?0ن�d��MiUhE1SF��b�f�FY�oM�G����z����͹[Vէ����N襺6a��6���D�L"����BI�/b�|||di��:w�}�q֩�V���NMM�֐(L�f2�-�����Y陘"�:~;�, çy�"�ze.�z�����D�(�źcn��qt�ֶ�4��R1�:��>|�"��QDGQ�b�R���OO'7�T=�tj{��������˧1ל?p�h���q~b�$��;����xuɗ2���Cä '�st'Y���Tl14p�lZ�;K��2�+����KM�y>?><;�w�Á��Q0���Q%�bh�/��a��t�����dDv� O�d�'a�姦�&I�&9�pUk~�R�8p��O���L\K�|�F��Fa��ae�xd�QDGQ�b�R���OWN%�N��� Z��? 	������gX꼼�PA^r��M���#�B�&�C��h������ҫj�DX�J&I��/�߄N�a�B�g;�{l�L=��Q�
oϖ�<�h��+�~������G\�����p��E�FO���
^�x8�0٬��.�.rs��t�� Ƅ��yq#d�g�ҏ\i����>q��u�G�<x�D"�(���S�J�ꭊ�h4�zl���/E)��]y��')�nT�;]�9UVZ�4�ݘ۬Q>$����1��LL	�)�S
>}���LG.��%��DL��P��չ�ln�Y�GMD��k�F[�4��e����][kc�m��]��M��v�̰���S*��s>�#�b
�u����Q�/Q���.���[�h
dC4�3��O0|�D$�bY,�:�/(��f�p����@�)zx}��ƫ��բ�kU~2x�����N�>I�òtlD&Q�J<s���J
5���-��Y��a��TY�rh�t��?��'������
A��LK��aMHj�Y�X�q,Ւ���_婮�Q^v�	��1�_�Dȏ$��s�$�J,f���`�@�u�Du�-�)�޴���X'��*���6��bqe6	�t~�HiG%IQ�,�x��3�ҡ�f�9���\/�I�e>��G�Уq.�w�#bd�$ӥ�jIO0�CM�:�CO
}8׷�0�oF{ou�ce�)�n�������}�d|(��RrE�_<_ �e�ŏ��6�{ʽ�[�����������J���O��Z����_�5}��ۊg���q�G>q��u�|���1�[jSսi��*��4��Ca�'����f$*Uuݪ��3K�y/�yh��,n[nu_�����5�Q�/�ژQ1�J�#�a!����L��x�:�H4a%]�-U)��
��%۟g����u�s��m�b:V�R�o�r;(U��B��	Y!uDO�B�f�D�3���G�R�Ş<YrvR�E�%�sMQ�R�3�:ϭ����UQ+����o�䫼�8zҲm$2N�t�,���u�|���?1�mJz��=xCĐ�J�M��6*�s��&t��<֭֝.���Ä��a"Q��9F��cJ�%e/�jkc�6[[u�S��!l&�ڊU�O��6�؞:l��t�こ�<�L��f�⺜98P�ʢ9\4���:L��H�ə���Dv(Y:;5>=0����-��'��c�94y�Οh�8Y�ym��SG���Z�˹�C���EgL!�����W�.|Q&0��,�ᐎ���F1�mJz��=��b>8�g$�����M�f�8b
Ej-�G��5�X�531��=/�R�a���0k�_���޴�5��ۘ0�V2��ce�.Kfl�$Q���f�� T�⣤EN(��@��.�g�P� lgYf�&ű�2A)H���N�������_U)	Æ�����0Y�e��[���)���5نCe�5��er\6&�4x|�4l"lL�!�@¡B��J#䣤�I���h��9��2~ߖ�-k��l����#C	$U|�y҂���B¹�I
Q����,�), �k�FR�=<2}᨜��҇
�sϜ����:`�:"Oƍ������K�Rُ]m1�>q��u�|��h�<A��
$��ᰢĒ�q$�!�>�������8Qa��b�����%�u0T�O��/����9�3����M�p�tᆻ��i��S�݉�R�p�%#xh޼���������`�k��
x)��-�]^Z�!.�9���a��B��l,)U��5y#��Kb7���h,�|�\��%(�X�
�)P��a�ӧ��{�(�4l磇F3
�(�i_��N�Q{�I$GL<3���E"1�cc��E�E)DF��Q�DDz��8��|�R#�����D"""")�i��DGQ��GQ�"#��H���GQ��u�>q�^�8�>)B"��"��"#�QDDi��E""DDF���m��DR-HB"�F�Z"#H|���#�p�G���ޣ�1�c�c�aDDDGQN��]u�_:�1Lc������Di�#�q:����q�[�)�4�H���4��c$f0ad�]L���wg=)��o\�>a��dD595�6H`�q��mLlU|�kQ�����i��47{�y�[��޸��o�U����[�vuP�z�z��b�K! q���^���}�ϧf(|/��%��ooٸ���z_��%�A1#����w9>������2g����y�q���>�}�2;O�x���ġ�����IpHR.BF�j���щY6���樉sp�	pX���@,ZQ���s
�'�f�k���V5��w�o{Nh`�~y<M j���RGY�=���ݛ��������d���x�̒I������y���RI$���f�{����cu�8�Z:�>DDux���EI%t����I @b9������,�/��Y���>����76xh~)�O	LN��T�U�W��+��>���ݲuedn��B�ڋ��r
�t������`���IÜ��^$�Ƿ�Q10D���)���P�<��t}�o��m03�~�1H�Rg9xa�\��
yv%�����r�l|@�TtFmV���4����F1�8��G]GȈ��1�mJz�����g�j\�UP��!��N5-3S�Ä��ӆ�8�����{�b�m���eu��:jl@��Ķ[@�6)v�H:��oTyS��~s.`����"�L�[
0K�)V����n.E���� 'G�����q�e̷2ܟ�t��l����f�:S[\=�-�'a��''J<�A'�/���~���*QU	.|3uQ���FQFqUT��w�"#�X�8��"��Q�"""1�mJm�M=}}�0���%���h�Wp��b����f&]{��4�sXi���	���Y�nƚϖZ�Ri����x*9�x�je�.s2+�C@���ju�e��U�K�n�VXR�KN,��m�hG�&h�HڃMQTr颪�B���9Z�$2:�ʽ@�X�
�m��0,(Q�2**'9�֭�K�6�l�me�=�j2��	qz,�G,�+�Pi�9� �K��{1ep��1�4�=4P�NMY�J�a�A��,>凹�}d�s��l>>�a҂noP~2r�_��_M�U(��	C"�A�4�(� ��\J"�I<�A�9f��p�1�~�(����0��$1�2T��.dИf�d3�4YY��U��/FR�Y�!�	ӄ晳���A�E��)��FHΌg���E����DDDcYM�a�����"���2������Pd��[�ό�~W!g�C��r�m�M���OJ�"�"�,GӅ��_ۘR�;߱L˃χG�<�M��͐�>�o��N���*%��!�.��i����<t���J(����3�,�̺�PKpi���Ąmk.4�\��~��&�`��?8_�Bi��Ta������z�mNWΥ�J�`���}��V�/9�B��4���s

�i�GȎ8�����Q�""�ǧ��	�Fjp{o��q��P���煣�����"
p1r���\�i4��ZP2�6�=Q
	�|`�ʢfQARtD����uG���/'�/}�ͭEjJ�D4�T�%M2���6����i�G��[>:y4n�|��7�Jwo֗A߼[�uUת�����J(�ũg��|�ś�D}����x��a�3��I�j].������L���&H�9а�_vb&y$�b�����Ǒq�E#���DDDcX&�a�_�n�]1��A�"@PFQ�P�a��mK�4xs{:xD��
��Ҍ,�yA0����m���ߍҹ-�MnYm(�M.�\�g�`�\m����?'����.�g�P��P��ϏAe�l�J���j~�·�:c����gӦ�a,�\/[����D��E\�V{^�s
$�g�$Z\�ϑ���,���Iz�*�S>7�:@`i��K����5��Y`�4��i�Y����Q�#���c��֞��~�RA�"$��tlu8(Y��-��-�����b���'���h��UB\��ً��р��XK�p��Z��h�8��k2%nK����Ѕ&�n�\v�ŸM+�sB41KK �i�&^� J�0�
�k����$bݜ�� �(�b�F�0Us���~H��b$��6w���?r�xYx�y(7�A�A	��[J�x�S~��)��p��=��&�g>��xSg��<���)�$�80O�⎏���E���߼�#����кY�H�=~*`������Bb�u�[��Q��mU�P�5*�9����i�T/�JQ��r&�qp���KB:t��θ��u����DDc,f�4jc��lmt1��{NᲷ�$��|�e��9�ၹ��J<#p�ҕ�]9Vt�I��9���ѹ}$����Va�Q\�􈯐�G�0���vgÄ����z]m�S���d�}yD��m"ܔ�JT���%a�v�Wv��v��"fc�2�2L(�!�E��n+�(xZ(>+��E�O
pᆏŝ2����eǣ��4{奶�$��v�o��z���8��"�Q�#���c��֞�s��y�ߕ����U��t��S5,��-QQDK�]^�UM=0������ۣ�Pѽ����j���PI$t�{�*���P�&��'ON0��u>�kݧ�u���B�B���|Em�.��n�e��	��#5�7T��`M�ںR9�2�=��/�\2jQ��BM�V�������\Z���"�>?�a�����	�����g�q�}Ne�k�:����=F+������7w�>�TLI ���
������'�u�X��㏘�G]GȎ�!�,�GJ$��ө"*d�	@ЪfW10��7�T=�o�ܩ�:ps�oM��C'5��ʎ�6y>QF?�S���jϏδ2��S��Qq�ːX��gQs�.�n�5t�ٲl�ϧN�&���ٹ<M��F*>|��:z3"����||l���i>;ޖ���>�k�-�y�N�o�`̙���pO��M���>�t"#��T"��F(�n&�����0���x�O�o��u�iK+�U*��lٛ?�{�����;��+���.W(��M$dd����7�#��(��Ȍ$8XC$Bh��"h��������D�dM�m�4E��E�4YȚ-�h�mdB-�""�&�"��Y",���h��[E�M�4Y��km4[DDD"h�&����mE�DH�������&���&�"-��dDM���r�8Ț",����",���,��D�D��m��F�"r�D�km"""�$M-�h�mm��h����[kB"E�YE�"�DYD�m"",����m"!D�[kD�d[D����"Ȉ�dH����6g,��h����"��H�-��""-�""kmdM-����B-��Bh�h[D[k""h�mE�"[i�"Ȉ�����H�$H���m�-��""DE�""D��D�DE�4D[D�m�"-�""�m͢,��-�"h�m���h�"E�-�E�""Ȉ��e��m�""�m4�D�d��E�%��i%��4��i�4�m"E��	�i�ie�I��I��$H��h�,�&�$H��-�%�$Ki%�ikI�K$�K$�$�h�-�H��i�h�I��-�H�HIf��"[I�KI�K,�"[KiKiKk4I���%�iċ4I-����M"Y"��M--�I-��Y�Y"D�"Id��d�4��%��5�i%�$I-"E�K$�%�H�Kih�H�H�$��"�	%�$K$�%��$K$�$��$��4H�H�HI"M,�D�ZD�ȒY�Y,��ZZ$�Ihܬ�&�в�IdIm-$��H��%��[Im�$��E�$Y���ĲM"[H��i���4��"[H�f��"[H�-���Yf�d�$K$%��$��%��[H�Y��H�HKi4�[H�Nx�奒ibD�Y"B[Y�D�BD��!,�f�,�H�H�Kimf�4�D�L�&�I��K"K%�KXZIdId֑f�$�$���m%�ȴ�[I&�XY&�HH�I%��Ĵ�Y5�kY�m"D���Ki-��KIE�Y�,�"�"��I����$����4��%��&�D��I-$��Y���E��Z�ZH��dZZ�"�	i%���i4�i	%�ii!�<lr��$KKi%���6�^�l�5����6[,�l�5�6[-��t��[�����6�-�6�X�f�ɛ[&�l�[-�l�ml���a��,LhA�m���!f�[f����Μfܶ�Y� ��	�M�����&��p�B#hABlBm���,�!��s6� �h[�$�Z8�	�8��CMB��6�BB�k!!d&� �����Zm�4�d�kF�Y#YMh�im��JI��Zh�Mi�Mi�d��h�Mi�h��I�2ɤ�5���kM&����Zi4�I��F�Z2F��5�Ŧ���D�k&��F�k#!4��M4&�BkM&�2ɦ�ɤ�5��M4Mm&��&�i���FD�Md�5�D�kD�M�e��4��i4Mm5��M[FD�M4��D�M4�MYm5��h�ɢkD�M4e�M5��5�M4Mm4Mdd&�4�[M4��I�ki��,�&��&��4Md�4FY4Mi���h�&�5�$��D��D�5��Mm4FY4�ɦ�&��i�M4�ѓMbh�i���ki�M[M�dMbh�&�M4�M4��B2&��i�4�D��D�&�2&��i�ki�i5�����i��ki��i������dMm4�M5�M4Mm4&�2i�5��MdК&��i���i��4�Y5��4Md�#,�i�k&��Md�M4�#"k"4[D�mE�D�E�&�h�[DɔSE��-�h�[D�m14YE�ME�i��Ț"-��"-1h��,��E�4[D���$DX����,���dH�-DB��DD�"DE�DM[-D�h�Ж�ȄH����Z""�[DD�dH�DH�Y��D�!"�h�km!dH�DH�Kb�"BБdH��Бd$Y	��B�BȑkbE��k-�Ј�H�H��--(H�$Z�YB�H��-"E��dD��ȑm�d-m��B��[�D��"h�DDYm�,�"!h���B�Z"D��D�[iD�D�E�E��БhH�km4H���Ț-�D�e��8�8&��D�4M[i��"h�"-��<lp�D��h�m��D�dM,��ȑ�ȶ�h���""�"�[E�Y�dH���M�dM�m[kdDD[D�h�-�-���m-�dE��$D[DE�"ȶ���D�hH�$Y�-�E�M�"h0@dA {�k�<gۿ�ɹ�q��v8g}���n��d���kY��Q��3�F^�Ǐû����|�?O��3���۱��N[����{;�o����n����~v�����z;|���x����ٝ��)���sм���s�{|=.Ǉ�s������M�O7������<���|o㷟���������?x��#�oːٛ�n"�\������ѿq��1���7ߵ�6ys�������z���u|�i���v�hٛ�g�~~��J����չ�-���3������v�M���W��,,?��{HIe	��;������ϳٻ9���9ۮt�g:����{��o���8�6fۏG.q�;f:Lc�33m�n�g�B��ٛţ68Y��l��M��� 3����B�ǿ��B�������u<�3��}OCuo%��3cP��l�BFlP��(I�����`������wɦ�gc;����f�ҷ�v����C�C�:8��~�_�}X����C��z��6fÌ�no���ӷǳ��۹��g��|۹��u���nӦ<:��f�m��7���׺�:7��?�<=;�?7�{��|%�v�ǭ�a�6��A�����S�x����?#����~�����6�Xm����6f���o�mm�����t|�y�\x<~�>m�;�nx���ɳ�f>���l�:�q�<[�9ާB�,��͇F�O���l�6`R!��D�6O�B�C�nB�<�s����0LCFI��ɸbC�O�[����q��o_����>��f�^�v���~_��Ϲ�s׽L~_ONX�����#��z���79m�g��|��{��{�g���7����o�&�{��oﾖ��|�l�Λ6f�ό�[g��m�m���o�l͇i�����������c>o<�?I�zv�<������z��we4��)'ǯ��:�*UӍ�n�y7ѹ�菎�&�������wLz;���ó;<���n�����v����ަ�o.�����y�Ϳ����y�ަ�7���wn����ݖ�lS���C������x?�����G�z�-� ���s��/Vݩ�����n����~� zN3�q��~O���/��k���׾u����ޟ�8�r4��坿���]��B@.��t